`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveA6kkXSsx2qXJpReDQz+KrdGJ2yXs9bHoO7w0vdjaWr/
hD73oiUl1F/HTCKYjCOtPkBNz1i9Lg2JsYONXFM4MRQj9YIYFnSxqUDJpSnsI0EW
ynneQQgnrhpS7dFimQgX0Jyg3eyJ9saG0vkyPNYvxhJyDwIAwb882JwiT8F3TqcH
PJpevoGPypX0QyO2a5asIEKgw/fOerhuPEx243+8pHA0OUHiTDvjy5EmAKZL6iCx
aYVQuIOqj7BLp8QYiXGeSWNOBhhpz00UQsQ8V0/0MD98f797cfJS8QmFlXNQZ4si
Ei8hl9Kznd6n0s46bX4MYsvoADoM61rsxDy7SGqBVHXCsuOV71ilqomNEoxenZgg
rI9SLtX92qNl+SLOCru4QIfHNxd6U9yStdpuVuRhobfWlxKKJm4ubGabJnrCHIF0
S+6T11YFk0lyBBVDU1D0oT1+eEXVC8focs3gG1k46NfulsD2u+dKEz5hDwKzySnE
dzdaN6zneONVZ3fb8TaWlDGSXyRanRq1rpoburs6qOwbumZe4XNrM+NnmQm8T06q
n6DMb0kdAyo8Bwj9OfyBXg==
`protect END_PROTECTED
