`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJaFW93puFVqIYfnx7jsjeEFHjBDuLMa+zX9Bdff0zvw
yuisUgK6M+eDaI24NLuDQhNcyP6QOx5Aq7R30AChHhusPDG0xNJP2HCuf/DSBeuw
2u9GfZxxuTu9gyWx/4JDcZOli7NlMmpZmjLG+SLjNz+0cfUO2bEJPCPTIbDgy1FE
91Ec9LF8Jo8+taXxIJHix3d3tT4Gsl/RfJ9Zqv/f9iwgc6f2mGDZJZQwTkt6X3No
jQcESzTcpi5uN7t3W5lbBZO94E2I6el/JfSMKdLobh/gIxobQ++NKutPMeG7k9VF
OEX4Li5inrfyJqLyZOZ1Efd558cEFeKKPDfI6LrrgIiIQNy4IzmkjuCXQ6h4LeYV
aCb+QSzODfmmw6lejkVCzJNlql6KtCdvpjKaL2rxf2wCnIYonHIR7+9sAzln0gzC
4VQN0ZGKf+5JB8OWkmQGphNObQFIbrSY6dcSiXsjJ30=
`protect END_PROTECTED
