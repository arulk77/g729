`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFSa4qu025EbTaoqKNeoKst4cQmn9QZHksaG31SqU114
VpSc8D3F35O/ooow46X4zQUiLnTSF/yz2lraAIxj/oswO5MwAzkZTnDM/czyj6jk
X4DhQEisW4GqxtFb2mCbm1ma4Z84r88ieAXlCCY1s9rYB41aJdaLgcr+S1rqfn6R
vnmh9+T66vkfxR8n353j6JGlXD1a6eC6Zkb2INOn8oXB07p1i+CohlX2aF+ZADyQ
o1FObVLxDtTQgVNIZNNKhSD8bCLTMTt6y+cGQF/vBu5luXm5GuWOsOHxK+jBAzx8
GNp48tssXClhfFGKrotm2tBwPd8U2yDtpjsBQ4W4Lisw2A9o5K8lzpadpbZS5Roq
1sGzTFTDFSuVunY1Lcv6JvR+o4pOLJzNqO4Wv6ig/FqSXJfA6CdBPcDdApEJwi6q
a2YF+BPRr+o+lD2Nn5KIj1Tb8QBY2dkPX+Xt1tSPLWTDvpMGFu8y6oUEYr4t2jb3
1s8vviqTWzQxhf/KCrNGbk++pc+85uZWSdniGvCVwUmVXBv/3f5Gn99L/VjKdfK6
`protect END_PROTECTED
