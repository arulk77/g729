`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C3pT4YqF4TsAgAfP0frN6INkHSrjKJBrRN2lK3XCEEt2
eaDi04ZhBsR8RgLC5KRBs0YG5WwzBOqmgZcCFe3dJJ2947lT+2M8CJBgqfM1HPOo
GcyJe+X04BwXmFvxUQgvoBPvmpNMZNO1+0zABHnUM5Kbn6i6KvuHfjXME/Gcw4g0
JffIyiUSESjJ3xK+e+k62gLspdtzWJj2WuKJYHu+5sXEmlVddGLSEfAuFewiJl8B
m2WoT/EGOfENCFdPjrPf3TW0Xm0UKF9cJiUT6ypIkyJqbvn11snjn03D05X+Dm2I
Em27CcnMcBgkNztlYWBjs8be0awx+B4YJ29hf9ucw6KPMXj+G3x2N5kuKKOsjw+u
BXeIwf/8PD7p8Wb3XoWuJ4NBwzaMeMokvgoogCA7CXeQPSA7Uo6JYfjNkIqWIkR7
Pe/AMlLRc+adbvAIcvXABZY3GjmFPzDsi8WPa13a91ti3p6ac3bwojKOiJRre9zB
D5HPVsCh+hNu82p7nlzHlvrOajtYRj0P18zbn5v1KvMIxhY1X/WP5j3g8zE+eWdH
IP9Et8RvCVjXggujF0D2B4HNZWWNTn2p4W0WAdDA8bVazEG6Ujh56yWeh8DbCNTj
auoGAWEHCn3tfDkhuIAjo+EAlCzbwDx7MBN9hRj1f533ZBbLA9uA8s79fCOQr5Ht
Jw5z34xG/ACL8nIRRQ0ZyaWOVY8rjEtpzi1Nb6NNRbFqjrEIkQ5UQ8ywBSCU7q9U
FSeEy7+QEV7vQwapJ5NUXUwWqhkCSDSAPprEH5aAMhV96vQuTBm4PG4jv0z8VhNv
5K5GFkWgerQaXhd/J0vZL502ftCQ3dXCChY7jWfVv3K/J0syKCyx5P70IEA9LZsx
Wh95cCqbkWLvvuC5KnAVn0eju4p1tvR2BX77WTqy5BSCI5fWKbGbm+x+fkIdyXpK
xa4jeO3RpVshOggYJ7fy7dAF7aZjAmZaaCiN7NHUAqk0+kbr9ATzVSpBFjZUL38R
t6n2nVOMSFQw7i8dlxpSJ1RZhlMeD4HxgI42A1wPReI/QNo8QvKGOQDk/7KXmEu+
xVnR/AXVKzFN9DGliS4lY17behid8o4lfowX/7aK5zsp0B6WONicO9gRAw8fhZmB
ceO4JMLofeqxQsSVKh67LnqVj4RoNIBOWJ+quP8b1/VTNUu9CLIV7hKT5O//zfSa
siO0DyqAdTbFE+Y3TqlqYDfIGgm1JujcNpz8igIxey05M+HPSSEaeXobN1XgS0GG
Mik+sCnC2zdYzj67pPl0NW0TiqqZjIPk/beN+f+2ABYWzfYN0yfNsxvpslXbhB8m
`protect END_PROTECTED
