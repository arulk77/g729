`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
WtahYbPN1+BDOXTiX23QDnkCmaaz4w1gzjMz2HuliRiAW5DE1HMb6d4jtFSIg6Le
fpj22OJCaPLWuPHil4mQqczBsrW73XrrLVVyldlWb3N0C+jzPHtu3Q7f6XfRRO7p
S19FQ4bTxGn6Zvfjxc98njGqY5boc2Codypv3yWEGEZP4DZezgtU24SoHTejgqF8
zWHXZwoxsa4vd76rab5nMumu0ZMRNeXMT75gTaiF0+cVqf7e5YImw+ewdVyxQQp5
50I97oSAFtJwdM3Gh0GhKWVdQY9kE2rvo70X/82aQUwzceOgQowPvNPKq5r5w2Ta
h3/M73wIq5IcvGjXlHaGznBXDrHAVk/K7iJ0k5PSz4Y=
`protect END_PROTECTED
