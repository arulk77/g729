`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHXiEqka8kfpws8Vc3TN8DVjGJ6SMlkft3uqVAAgFNmq
WTYi7Ua7oZvHyudQXG0Kga2yJTxpp2+inSBv1UpaCY+jk4R7pKeT1f1bpIHbgrDM
ftdUtt3q51ZZvlIukwR/bs6H46Ndb6qboKReHlqDXP3G+16DdEgZwTE03dVLpQMd
qRqsKVXKuSSU6A//R3UEzC+SKLU86YF+MlFKqxS4I2TPc99JZFMlnBVmpR49MQPl
MmCk/rE/csJiQ7pd8D1CvdHlfDDyfF8Wu0u72fGqJTRDL8xs7m9TUd40WVcfVoYT
qKJ3pQ2f2KJ16w0eOj3qzA==
`protect END_PROTECTED
