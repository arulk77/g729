`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
fZHSJlnpFP09p4Ry0twVB5da9lbo5Cdq7sSP2narkIF+nJoC39DIeC+00oC7nIJC
+UbBrfER4EcLqx/undS0LjTiNeRomoLDDP4ZD+QpmAMCU/yN+mDf7deMcso5yh9e
BxTHijnZPZSnqHyeL75cZE+Tsr/XEHDMcyVNjmC6H6v0fLgaTdxgFRqQ2ap+z9zO
`protect END_PROTECTED
