`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI9aZr7Xv88anYEQpvRyZtbR2voW7T8fiSg7Ez+/fXT5
VnYECkhczFa7A3vFEkxx9HwVSrxd2nxr58Y2dMLs1EVvda83/1k2HtfZu5BpBJXe
SS8oDXYGqgyeuIjD63Ya0lLfrlushD/TgCsdG1kTRZPxhMGC7qy1np9xhkV+HDec
K17G5GRFM5i9d7RQAvZ6tNRJLI1HFLLq36yS7uhUjW85XRINshP6xfe+8E/DBohw
AlvxUDrQdqDtQ3lkoqwUWdT6RjaUiliYPjn6ZRMNWZJQ3JqqJ184jE+wn+C1K+7C
Cy03B0GHKKcnIRdkBOIm9lDPaKCxpv5KD+i3c1xkE228O3g98TaXO4uUSWOLMRwx
hD1C6aHsxR7sJZucf5QAYcV6feFOx9sDSFfHSfRCnRI8vjH7ud56wGSnfrxfQr8a
denvapi5Vj1t0So/s9b1Xi8GdiQidy8WhrJA82Ox7gkenBCMDAg+Q5MlVuCtSmlk
`protect END_PROTECTED
