`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pvbjr4149dxGRwC/XJov1wDDplAeOHOo+nzxoKd+lPOsXNw/G/0UDJuplFJJUQaL
AArUs9IjhkqmdaF8feBTTXekjaq8aUqZZkqQJ3dL5QTVDqBisUmsWjUa++kYg6Th
Bxi7w93/rHVKSSDh7yeIC4sIdSIrOO26c86t2JydXkk=
`protect END_PROTECTED
