`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
if7OW3neLerq5QTb0GME9weXK6UH94woshqgNNlX1Qs9Q6EmCdx9N9o6c3g7wHr5
RogVcin1k1YsdbO8LBGj97TBq/GdMyMu5ieBEOWkf0d5/bjCasnj1W4TyjEpDBsY
YSvMBETsu+rVRz3W0F8mkoMdD4uBiFVVI1/V97a00eMw8d4FGby+Wzo4L2K74E1D
sJwd3AIgixo6b8wl73hC/IOwJ8YmO84Ylyl6UrZVAFFsw7EZFlkigm3Sl9tFNdQn
`protect END_PROTECTED
