`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIJ1Pzh20yVyKY8CxO16IhBLHFZsIZuVORyii9U2r7uX
NwRZ7GNEq6aHvQhBwRzY3B/Hx+hMDAz5y4+gpBKi1OxpE3iIzS0SxEprBTc7LKjK
JDW8u1bREx+z89TzpBCGqa5yjp9oj92py1GVIGUo86bitKooD3+nsBKt7hKSN6Fh
C+iS//KSAHhyVNSLOL+nd26qF1qklUJB6hiiQ9XgB8SjOdo4MT2fCzd3eOAOWCDy
3ngiLcMkYn4Aq2LmQGUL3EZivXZ8eCiLFLosu72m+4XXVQGvd7nvSm84qkwpG1Ck
GTAnKu4TEdKbCJLWRh4b/DeprB0FFgvbhg3iI4pYR8rLc+NKdcFQKgXLZ0qfZglh
+8TOlHceQbXEB7rAYqUaE5YbFwR23usmtq+jzH+8Q9ekK9tSifb0IuWM2L0+4YHI
7feEMyIcg010IV1SjBcfIgAR6gFwo7e/M+sKwbsgifWDkwpWOYn9WMguf4eivGhL
1fb9tqrdUa0lEP2CXfh4y8d3ISIVZh9ggSVMfFThElo=
`protect END_PROTECTED
