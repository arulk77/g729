`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNDL2JjtGFEXSQIUSp3ZbNGJede3BvvPqK/yn8bmEwsp
iyj4HFqgJC1l6Jq/C/VMCugcvtlfuKbuhFqy7wWZqu66bLp8XUu92RYZ79nfrhDB
ev6WRnK3o/klrbKv399E/ZlHvD1lkErqJf+knJ/uL4mVNVSBzyHg54CFLiE3p3nt
V3d227vh3TPvTMvanK9zXjK5/2ntqTNzEr4IXvf4bKr52SFO16kTUYkRDG0HdXHY
v3+RXHhNS3e0sJw2W7lXowtJItRjzyMKV7VmQRYtLUSxwtiIozw3Dwq0urnbx4Vw
Uq6nyjceEzUyVLdIVH99ax34c5kuKhlVDvVQ14Ob657/Bbz3+eUwiMQsEo29mTLn
nSvZUsmSQJ/hXXiK3uJ8GiQcFRJpZIRW1Qu8GmoDh5kClWeEGIEnvjJ+dur6cNhT
`protect END_PROTECTED
