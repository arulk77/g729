`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKq+oyGTisv7gTDjRNcFdoLsQQPPuiIrqBYzyhzq9vZ1
GDmxlgnXSqSi/eISjhyyfsPt+lRLRQx6QpO7jUSIdEV/sY192ipMa76T5Rdm7MyA
los7QpR/empyaUNOZzP8lW0D84Wrgm6d93hLCB8jrHRFJX3VjFkSNe+sZTMpj7iR
D9vVDlyfNFwVtSXX3X1pvTWLdIs+/7viGtW5oJsXUce0ApPivsRQ5bzuKppSeKz/
D9mbDulF3bDwaT8j+9loFyxnhziYp6P3yXiVb8Ku8f/RdbK6aOgUO5AGuJCbzHcP
bfGwXF85vLNqdVpl5ziHXpHGub+nM5FA6eJvwp0ZTrH6J0ANQt5glFsZHyBM3yib
`protect END_PROTECTED
