`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePslb2MPTNWQkMQpauXoZGpuJMgyXf0Ts+dogOoEcX72
Yac/7O/DoQvGYPQqJpN51FI45dk94THvmz5cjrpzIZM+qCRRWPciY1tTMV2/4VTq
DmEtx4hg3uYGExv4E99BcW6ZJW7maGzWw8nCk7N+hEo9jDd8GuaoGibPKK8YKz/l
AqSIrOnjvGSh+PshIb6kleYNqDsGRUydRD7YXFN23/pHPYzPw6xeLyNppcZcYMVV
bKUoWj7dK35vxUW3k27eYnh77VofRNApI57FtJ2nLyKuWdxwfAEVUhU/ljCI9Xb1
yFTv20vaE6FqRNagv1AxS+UpIviawZhuYINsVIPx8mSdn09oSMzxRsCsq7UNytuQ
/ybAcc/rhs6DL2n9L1P7zyiI9mtc0nDSWPDKaAK5cHwp1W+2su9urtOWAlP0/lWx
LSvQhy2v4W6vCpGB2cFAiaGVISKm3314TKsqpybYLZxtvCxFi5HQeMe3tE+H9ZjP
D3WK2/IZQLSM0a9dg95Pre9bxkZUsVLoYMPM4geOr1kxDfzoZNC8QghWcFm4rszJ
QytBNVsu9Lq8XAD0cwDfeqspC6iuPLYdCA6YxNEx2gk398Kn4D+clxuqZi2jevDl
`protect END_PROTECTED
