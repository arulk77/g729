`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBKnefVbV2s2d3fLmWlFiuBjrAzkrSNlWcZH2nprDXIh
sqYKzoQFufVlTS8Rre43LQcWlXGekvWUhhsb3TMPlyVGEfwCGtfywgOddBzjbm4F
pIahxcZQFqHje2cI8AELVoprxOwozt4O6hd9O5ozc3nJk5u/2Zo6e3g1F4zb/vdu
Dnh8HGG393gSgRrBzPHjNGX4YB1+f2NXucR8IgarSIeU4iP09FffxNqeKl3np6JA
2vGOZ5ZgHJc/T27yNduJSUPHOMALrf+Ce4LlmHR0detmHzE84W7tZujdleiI+fHL
Bid+/rI6t37sU0Geu8UahxY3xhx3el2lBo3ILNVSi0cNQEKv3TfdR0IWNT1Amwab
`protect END_PROTECTED
