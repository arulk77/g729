`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGefuF6qq30Zq0kns4p+JTJnm0wz7DeG0fVRx1SS6aHW
j9dTMK7Z2maFJ7SaKr7qp1Kv5vnN0+TfuHuvcmt9nbbo3smGWDfCHT0OlKrqdAy8
2Are/eJvYwIZx7OLz486oC9IkLKoRqrAS1O/nxYK9RZsArJphBoArzFZsyeROdCE
8of/9dIWRnmOdeixPEVK+zaVKozn6cBo72FpO823K6fya2TN40njlGIzGOoEjNQ1
BpL0cjLZ/b4d9jnFJ0ayEzEeWs5lW724JRx5xAbX9t7nZeRZW5NE+BXnNl522BGq
8QQHw+frU5V+6j6Fxh7ISFTeuJUySjdszn7TtUKqajkcb/2NUEWjYiJ7mtnj8W55
B9gD4IknJBp5GB+JzeTISL0QopZfRe1XiiwJa/Pn0rzqoToBWGBBW8vi2m6+CqW2
z/dRAM0FpTk7H4lGoofiPTGCEumnj9ijPuMcvm3N85DaHDwc1uQcAHNwj1p+f8E+
`protect END_PROTECTED
