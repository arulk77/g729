`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGUWh1gySWstJj5B33KX8DUNH1Cr1w5/Hx4My9rM1P0f
fQg+AbW9klULd4OTUUROS+Qcf5cuVRfjCqW0x0U1C30Sj62A1xlinMMwoGhUBRNc
P7w3HM+qkTWRFLlefUh5p2/jYh+HOaOIYPiLOln67MjQQ8d3hQqFXNFa0x1ciTj6
qK8xwUNabeKmM45QnwowtHlxRWEDipQGKY16blLt1lfEupMZDCJd+bkhxm5TOpV2
LsMvGdwfyqROQ9snMBmTA9FecPRl9EsftUPsFiBVzMxpGOdCOA5ia5FWwi+j1z8g
IdEZGpi3/Qa5+Dx8N4kTc1qTn2A8/ctXgMWJ5yGAFBpV6lIfSimq8vpNdfc9Ibuq
wPiE2TpcTQ1d/GxVQnmRxm/0lMEPdxzM5bYZpuxSTSeodpZfDkEU6F93Q3WMBhCu
won44tCg99GbkSDpxMGDn51v4nVDRauXKz7i1DqC4hzDZqMQEC3OVt+G9p0FNDeN
whUJqlIGys7uoNo8RsHuRwsHFTBJ6/+XBjrXdF4Ah+WUzvle7ci+E7KZ0T6ID277
4j816cCR1w7C8daLjYvCo0ugylUkD68QrLOXz7xxxwAOiPdU7W9lrNqucpguCpGo
HNvMYjJsRMQhbRJeeX5x22aEZjbT/ra+E+wv6dM8Js6OuB0EmpggxzqIMBr1LaFT
U9Z4lABacL9p2It3aZ5sh4wL1VxLeccSDqdnEq2HmWZiqCVtieFBipb1mlRGNCAf
3X/ihymkno0235Vs9tcPy5bB+1SQ/hfMO2ABg+oRwDNyii7RIgEcH2fakyZD5/6c
uX8rJHREpkUxKJGaTBUl5OVZs7oqaeurNvAivpldoLY=
`protect END_PROTECTED
