`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aaHqfCING4uwCXLTJ239ySBn9a/uMkPH2qi0ELvNR9O3
AW+00BGBZtq0xZwwKmw61GeShtOVAdB0UWgfYOYt5uRBmX8L03C7NSQw0ng6cr8O
s3n6PdcKg3Gn8/NGIbMvwKzMFPIfxMwGXyuXB56R3Gw/KswR5pn0X12gu2DFM/wh
AUy264Of5p9UY7qYathoSqSzWVBbf5YuJHqAc1Ld4S+42nRNzzed+nnVdeyfj2lv
VsXUFd9Wpcxrom1KghAFCU2gbQoFyMfxdSMNAj9M8gIKIYkrXgQVT2mtLs3Jt4bN
vR2OFrgAyYikt320QmGIRKu3QBbCFhao6qRGkAoM7Fb6872I2nwMoIi6wZxHwNzS
fmLuW9Za6JrichUJtFbYOfVRjP+agH4WcV5QTJTteEgBB+HrI43+pd+DrZKs6gS9
TnNwn9NXTc12EKKs11C3gkRx1QVx8M0Cg5BxhLItX9SsmiMijE3XjL5cShoYTT++
o3Y8AdJGx5EFPvoPAhDFn2Ps0v/wmg+d7eUNbmZEpLoCvKgqsQel/BG/7h3iCcgt
9Ua9a1IGB16QqLFkjNolsed9Fk1l4v9TCzVLGPdqgWiH5WNbGpQo3WlDDEVClLSa
nD8Hb1iRdQGqkyIPI1TV2QJUKP2xmzQxnTr5GtzkhICllmdEUvy0IrqFbngHqauf
uKfvG19YjwHEayEKJD+TLXr5LXEzE8eIinl0wgfMpcbo4HBtNo7cCRxWD9uiwK85
9yrzFoOrz3tYrIoHWu9m+A+FA+/ChFnLPop5LMhbYQbZW/y4TbgeqFt71/UiXUM/
WwbfxrrxWMsDLzySQl0H459sN4hHGfP8n99PKKXd8h6kDI9g/GFPD8jG36G6aAVj
ro2nyrsYNFqZLvcfrPxKVfpmhN/vr/llSb+bSwJSbhLNN3jGO7+Jat8DBQ1B835a
q5glEQfUti1H9JJZ8AdCH9suJ3hmDHAfIzPqIgcO9IjHaGDHZvjNlkO97Pcv39Q8
tHHmfi3O1IXZhytT/XXNFtbH90994g5OgkQLAztR2Wbnqjbe/Z+/qIypi2xsAq5j
EeoM8R2TyffCAOmuoZmzx5g0IMqlVa7vbLCkEQ4vHUvcejPHNFoUsAjWlIyFeL/S
m8xFhc0N0JDhZ/Eni3RPGJXoUPEdkuZbxj+m0DbkZDk8jo5tGYNVVXjbQeq6MWmx
Ce9iqI5sVUxzIAyAbCNxSMcpmkPEiI+BDw4DQOD30/BEShwqtjUKOD0FjU6w/2Ry
md9i+Ix5rYEmb6kdaPQtvUutw3aPQLnS0Lg53pX0sbhBY8z2tKPzKOOWWlp4dGpn
EGGH6LfE6U9En7lzRLBIMYjd/Mqa1XZJQf4nOYGaGRDdh+lc2zPJdpuQZkk1ogk5
yOx7vOv4uH1NlPmtV+MOgrEQe4qgeTntbO0Gea+3+5fKWaxu2P8o7PbqQSVAr2iu
MbJrqDXjE88lKQPCl9pSvZyC4ZH0i1p7+jMRpb9UK7p97Mmb5ucmFJikHn6jEVWD
eI1qgHVxaTHVNccvRcje5Wo5A4yO3JY2vqxhm8gVJVVGMxJ3KW7nMurOoct6Bp28
F7CWaMK2I93M6RsZCE4NC7dwxh1SAr2JNphhj6R/6TH/WWov7R6erp0PEymendGE
Z2UQF9XevvUUeXM9OxQP0UJ60chWTlBV7KZIPqIHAoQ7GJJQ2rcdilV7L88BxfrS
e+9y60NEJc5yPOdRhGw7t8l2GSlHyCy5kzIUwtM8tyVtrGymeVH6Vwi0OlGK5yIv
zzzJ8A2zufzSImn/cqmvzYnlElEr9CIFyvDXNZwKRZVOOMM70+GeZFfGx0QyG5vc
3k0gOAgB6iU2bNf5jcVRdTYN13WfUapJ5WEvm/dunvv/gavG8gFPpsyWYcnD0YZs
RpGolDKPSzcLzVmpc8jD8sHZRM+ED9GK3Ox/qS62X5UnHMsXFyC6hWzEwDBZ1yts
RuEzkDgczIxC759WNAVEqfMavk36zVyhk3JlMH1OFs5aVwqjYgIhDlIHUj0RMEMW
u3omqN5kNQGUaLW6KCzkgBJxmg1yG2dovAVa602quU3iku2oQyNdW7nLff/BO0o7
Yd30+m/0Q2nBOzO8pLSq9vWV7u28fXR5skyhEXH0WNPJenM+C36tkEXtoSrD1nL4
wWV3YRh/SxnfFAvtJuiL2ZpqYxsCK2DDtNUqSkHBgfdgi4S8Lzrhq2EK6y6ghXQ8
c6xlVmxPpddbxlN3qSelwpdpv0mtKucBh6L7UjYQCwuTW81LXciwzbJODaCxMbG3
/fwEOlPwJWyxWH4AfWYabPy8s1dsrDZNyRT2/7bPbsgd17tGTwq9MEMi3pZZKMDf
XxWXqtPgFaG4irShzXEpCWbanf2bsMTZ3Ma7R4W8kyrUMJyDte77e1GLXYi2+Y/N
wXvaJRX5xqdf0tesFdMUYghmCHs81pVcgKMsAwYfmwFe1+FQB7AicbgKmxAbxGJK
iUBGrsvMfInpdB6+KDxscSEUv7j2yLGzyxYP0me9CdvZzKf1pkamykX0Fpvm2s+B
z+n/FuA7fZHNjNdjJhRHE3ggcKXcGIi4LsMWcFs+7iZwFkHLuxtDuhRNLdFk5PCv
vo1QY4JQX5CLLNN15TWS+ZJp4De+J3dbAyL9w7AJKe2CPUfpfg6SV2dhLRIkYKyy
5mun/QeA60C0d+36yijIInQieVihkbI/bqPd8dPrT0xydaD0+ZSO4aoEoaVMGku/
TfjZeOik4jRBmrsF9wJamPRHadLhu2Chp7VFUqscEFCdcxy8eEy2EjbgCmxHmX18
DeWX72nqvV4auxN15IKcCtqn5IEdwhL0RqwtOtDKjElcUkPvBNHppXDdk1XlP6p7
rYdf5L3clmvbowSTiEBP6/LT9ki+dPrJLYNE+QzrlNOP9GAnr//6XwhpybEGoe74
vY3+CwfATbyMPgWtZy7Y74bjbXnDtxIER4LoI1GPpp8MMyHdIDSLQamq/Mca23xL
zTFJSejSWgBOVM3jEZsDSlnZEYVW3gl/nM0ajHTXcbntJWEC5F+Yq29E5d/lWvrq
Gys+aTB3OkD0XxuXBxHYV648U2HNjYva17TMdPJvpB2rgtwKmtheEWaArgsDHW4/
RUTbeottNCM6wTVIuI/5RC2wJ/vGW4kOW3ZfeiOxkoPN7YK+of7BjGZtDdEegqNQ
1XktryZ+ajBL3VW73SU/bwJVkxGqgH5F/2NVaPON0k4GSOgq7AkIS9fYqR60P5D+
TRFunveO5YFJQMHQlZV+0m9+mrwNlW9Es1I89+UGVDkZsolHgq/sFwefhTGA+78C
SJ5YOktTw687eJ+wLaMWXBBdjkHseKo4xbo4hxm6kR/Jb70P3QwKEp6eXr76cFGL
p78X+D8fKrhHjn25YH+bcx+w54lsVZPjD43PzPnrZK5ySJdl5V9u0J1xnkN2hPO6
3LRm7IFiH9ugi0ty/hNaItU3PgtPd+ZhTzHTWgVp+s9tPGijwaqXX1HtDaVQPekh
bQJ7uVgah5fGX2UXYQmrNEYez2GYsPa9u4xbKZzEzSM+86UaUSrURgFAQFj4+Nx/
1H7XMoNZg/bnyko2/AyhUcfuSPzlUx1mc/O6MkPQXiFosJZeJq/2LTBDkiEkMcPv
Io9L1LdL0kzdU2/N4GqX1YHeiwYIW5IAMKn6NecpC8uZnp71dwDBse+oHo6S6Esw
KD13Ux31ZxHakzeyPA/uuFWdZ6Uf8x5TBW1Qaee7IC/gOqCzKkBLqJYUrvGbIGx8
mg6UeaYcvu0TVojAqinNJdLZul/D8xG2f/KlorEVXbzMehuw+dquqo06iAbwDjrr
jA5igudbOO0f+j739148UPuYRhvRmQ9Oi9ABya9yo446mg4MCEgN5FMPbL3d25AU
krTZIl/p1+eGfOfWBcBq3QebtR+Kq4+ebZS3360QNCh3evYmB7X+5QHmERK693L3
nog9mvR4WSqYPensrqBlEU0ygresUFoJRVEOa6tqIwd+/PMRFWWotxEaNed4U1kr
kyzngmkYNotgKvKVCwXibkHqHbh02pFZTObJYiLesU5BkSAikq5SUdv0mRdF2ucw
qTyniBvdDTu3XvfCk+xr4uaAAXjy8AvUyvvlrUu9arerNXn/0yUksJgOiPQCOl18
qGcNRM2/ut5V/qUanfvOc4YqKZqeNsS+HjzqZW/oOYMGv9XaGIrcFWEbk8/I3KIj
y+7FX6EwZeH3NPqVf3uBOG+KvkBmHgTrdwbFEV85U0fRXsBOBDgfWxxe0wmMwbSr
Yi4YUMKsYSy0KtrrPL7MSPdylqJOutA2yz0R1FnumjsbBzGD2T4/NnZdedJM28rz
dM+rGaS0spAO1ilgtOE1kU+iBa8l9UhIX31pohLjKSCvb0N4BAVCaw2ZC6I9TLnq
32VgGT0ShZOjoTO2iFM92yA7wMJZ3Mi6i6G0o+fGhfQ1pA4chiqPlx/W7tpT9W/M
493l2O6u3QInZzK/Fng4fD0Vq0Fb0B3ykhgZwxIzPQidcwADavKoIQfP/NLlP+qS
QX0HGJ4rNoK/l3ud2yVv3MCGwbGOze6YyuKAbHTkJ58fkkSQvc8rsg6WaOWWf9mr
ly5RcoO+ChgNbugaLZwGYb56A9rnRJDCWSRzZ3El6WUuzY6w+yqLNImGacAGIiJP
M5TH7FQ7i4AKMHFANqenUCHgxsrxgzQY6KlQdb1xeVJbTep/19XVwb4SSwJFidww
YQMRz+Kk/wN8No0M7Z1cY4WbDQsobVuSvDs4bre+//Y/mwIaSWeIpzRDMQgoyRln
qGe9xkM6b5KB5CAaQlgqKmwxaAzrpvawJCMtJTV3WeUKVIPmr0ErSFkinqdX7ByU
e0WrhTsQneyRSVbqUKq3UBW5fQKeohe9LeRrwo430LvbcBLu9ytSgJW5c8OrkO8I
mfXp4s8FwCnEKCOK3w9ublGI0nkSvXRhfr22AE0AdezrGcc0yc3CHpMnWYzdTluq
bvr3j5EwoJFg+zg+BQqLOyUGVjedW5j5RcvGl67YlShpvNc98yqgTF5teBOfkXak
omCiSH7chHpiu0W4D5YY5lXcp0CzPf4kIL7LfxuUyYALhXAHe9cC6okvJsEVMPfQ
kZqBAgBZUYya6ZmHtYbW2ZNK+cL0mbkr0BdvrtvNOQqFW51OlWjCe7sqfiggeDV+
+DwY/zLLL1GHcW75GaUnQu2WV7sCcS7fWeQsVe85Vfes4MrGhlWTodEZ6yxk4kMc
vtOxaPDECFweCYiyUshD9r/RkucifJQVhLqY90e1vGE9f7aNp8mQaIhUb6pSMfzW
gPDDnhDkBPRFPWJdAfJWAy8hvkeMAX9uONqxONHEoDA3+b8rlpIWTwTlEjhrz4kx
usFKKiIl6p7JyIpoga3mmNLl+Ta90G9pcdh79iF+JXQSKEYI4XdEJmAoUeVtLYKe
DCXAKu23BgQFNLREeARHPIWxjUpVNGID7sY3t1fGdmvZSNOBC5LbLqw1RpLxM46h
zVnZB+ts0xt4V5spJbnDFHM2FDFG4uzzmHXA9Lv44J+ai+cxCnbtQu/MCcB81160
xyePd/58oW499Lbj5T6k2Dd3M5on0zm3Us0TN79Po1n/KBQzwtT4WlpgHbFVVVLL
kPLxpfZtPO2l/yXEEBZE284vOcDxpoj52TGUoQQTzYf5mhNeqa3Ve0iGqZXL72p6
DXxNCVmmYTgo9YrJoz7+swTXIqybOsmNdWZ803D3FB4ecm9Z0IHhMWTQgDlb6az9
bGWEbYOYI7CH+7xiFEB5AIOBxy4YxIbA3arypt2ixFYW1bZxdJPXXajHR5VLjazR
wDDl+64KtQ3nJcJemzyTLIppHiHByrSIbSWUq8FPwbxdL9zHQxCSOTxZGJg4gZQ7
ruMTWCV8+9BQToUmfUkM0O2M6bpNkCB35c2OSbZy1IHJTYf7HJsdRZcA7mmajWyL
iO5fZi1niUy0tIczTxYij5vbBF1GA6fRHAOJpKyjAlD3ViwBRplbDbcFMCORyvV2
l2hdcA9SF2PgS/OOXvdYXnUIevU+iuAxkenECISJ9x3Y6E1wFOsnUy0sBonqey9J
1F6IdYnTe09tJd8xJ7UjtGasRNp2VYVfMEyDo5Ese5FowDjU2RIG/Lr4qFM3GO5j
9U6nfutboOLOI42cqlYEyHxuBCsOr53vsArFjm5prHevFj6V+na8Qzt8m683ctL0
Fx5/ohVTNzzS6iN+RbhJzkXDo/tehzN5h1ViRhueme1DYrOX3+SGgT00ID1iXUDQ
f7otHL4h8UQlJqYpopi8qz85zk0rCiWcX5cbMgKdp5nukWBxZGjdSL08Ec0CEO+L
Uy1I1twYxXeiwVoXFLPoPREgVbRKuVL2NqYAN015ujjT3T5140Xw+xH90OYogSX6
XEmo52x1hR2u0KXz6zToZpEIn0J6ZYfMQsX55kDLnUH9ZueF7M2m3uLorlW1qkn+
yYqNmz2vrStxPhtaBSBSyzLwkF4a9QtZnuFQ8RBQ5a/ecCNLx+gFEJjnX12ghe5v
AS9GIAeM5kD7ssSsSwBkhqoLsftlHyTDIAIdPNaztzEndQrmr754ovS9rNNvd37f
i7Ool/8uK1Hcgx1zAx+o0gmeolw2Aip69ccQMAXKL8bgr2zhS0BbaBUHO0d4H5l7
22tytALjglEGmd6tPKq2lORzeIyTyWeKE7X+Hr2ZvJS7KXkwcbrhQy9bb52UKGo5
5wdrUEDOnvXvxk2zqujhtsT+xjZY8RhSEuehPtA2FITrSdGO9RCM0q3aP+2J8edl
rAGTb6lUwRYbbXJenI+c5LMmgJepyajf4x+17HsJNtC45oXv612YEzkCNwaCzb+p
uqoIGvrT2Ohno/1ZmkPhihbrUg95g5FUmxor5kDbyUOjFqh8pQ9Qa3vjPUqYlVIT
XDIhWQQPWQ6/b5oIofHw8bwZu/0p2y/cIcC3B/I3wzlne9AH4/EuqpiG759DWuWV
y78cEAiCMAFSYQqfA+destW7n9yLghPJdpDjhQ1dcGqKTZYZTCHbqTlPvKz6J6s5
RLccXhm5kJuoPX2RCQE+MWejOL0P3kJ9C/O8NXYH4z3/2FAAGaqRvRHCYWj4OdDN
D6whzEA4tU7aVPUfHBvdn79EVgA4SWfxrJtSXZzrOX4Bnv9YwcLgDd9tVu8zoYZM
gGBTPTA+0SFLqd3jaakPoGpGHiKmPJ5gKXkC9xu6lgFrwxhsDoAsHnqk+conlPbF
cUpywEDioxOIHfrI47dSHfnepquO1haGrKpeQHKgrhBPuyqSpK0Ac8u9xAukz817
d9+Qru9zm4bZFnlLwLN22oTHf+k4WjGxACd31aXEFhHkitCQRv95nBGpvYNcsfQM
/Ks26sZXyDd/X8Rq2TObl40zIHhXdDnt+pEwvqc5/hW/v9xgd2HBu58ir9VqJ8Hb
b+c4sCqHXh6BSLdEFBirjYYCBd0CeG8uett51NSoMAHiI2hPPVMrpF5w03sEfcny
zdS8QTWctGSdrevhnt4LCjz9gZPsxt9roLSQeZnl/2Vb7hcZRB4tUyDDG4fm9fvH
OczQ1wCzQi8bV7gwJ0X9D/pGQAm2oj2M2ZP0wMrQgouKjlHiN+0FYqZ5ihddRMFZ
c5ViLiooFYVTcqQN/cvjapCeqg/f7agfvBl/eLRHorXZer2uZt8Wo5kuoEXAvLKl
C90ZDjxnFmcRH+x8NlM9KdLCY49g+t/9yQHilx7wFUmSPo8dDZskN/7ahXURm2KS
eWunxvh8V8hHTSZnITT3IEvX2Ab4sbkJUSm8W927OcwJPq85rQ7D288Gkh/es2cg
F56rFNIezsD5LhATJSxu4fEZ9p5872VS6eYYUN6VcIB4GR6YXmkwMoLeKEiy2G2R
bU+iJCappiCuVQDRbV7oMbHvYOE//hOV0OgdzSmMVId4uq0nG/FRtSr5eqbTwsjO
d9OXRVut5agZQtrIjKaisnVHRvZfmPRGFIGAUlpq7vOWxe7/SrU5aZxm2K+Yoyfh
/bz1CTr1uLbA4yHmQLctCpSnzXoJIoFggLH3YaI121uHQDmC99e2QG69z7S+2pgB
Se6kFpdNhA6gyFq3kHvsi/Ms68TbKW6A4EmHDQZ1c3V+57b2jGICV/Jbmn/lHjSP
EPecF8m7Yq07ELhbudrBeBvY+8O1e9yT1lioD5xVvzOBSefV1Dj/b5vUArtjlveY
eTc+ABXK7EuHDcxkMIiVBM329To7UcANtSivIjuwO6yGGNwLMw6ac3SoPRsm+PrN
dne7qvKeIbYYs75fB1Fw4ZgrL0Ukk+8P21NmRcmCJQ9EyT22xcdniOzLf2f1EKRi
/MgbTkjOV1iYD4B7KQWZguXLeiUSYVOuWG9dZVJP413+4XCv0AHPUA3RTwf3ELL1
cTXg7Y2IpWosWuRmOrJnNlsCUB2/R+c/7R12uEQZ+9jtBKzKKfpzXl2xqRwNuDbc
0PwR2axBZPdgvm20KqSwl/aQy7m6LQomS99raWb/IPAoZj08uOA0qReVE7wdRueg
dZMkEBMXx/ho035DdNtarYc7pWp8Q/nO8aTTK3PlGtn33JJbxjqkCQlbFPahbYdl
91YgCpnGRiW89478w1SKUnfCAcln34PHO0DzgsiqQIG8daGJM64yzz7APPQruDwI
DYf1XKmYon4+cQvT6wUbOyxfpvdn6cFXAePzQlGru0FJENdAnzhaHAl9grVgvmlT
0UqPTfJCruoF1K05K7M8gx3TqPLH4yBrld8C6Fw7zNvrnSL+vxdW/Nha3HJQK00o
3VS0uFvm62bOxTaGzkwpZng+A0F5+7sxxH9O0fKLW++mmXErbDcedoWIvC48Dm6T
Vcfp14cxUYp3ewZd86yXf/x/ONZDHo5yCGX+GMfakn35TkRDRojP34KYA7kwoFK7
RAf3//lvaiXXETbYiwBr1IhC/S9JUdRDcyCUE3hdC9fGmJ8Tl/tyb4x+OlP5JW6l
Mod1xBT3EiPBDfzLXL+vV6UYSDjlcDRg1FcrSVntVNPUE1kzvI0TGDLMAk1RYRQR
9Gzf4RWVWHysQhuMWzmZQara32kVPOJ0bEZQ7Lit/T74I7/SEPF3nkwbugxRHYNS
Ko0UKXmSvh6RcN+p1FRk0To5gfceW2adVqCvN98PSdlOOCi0b5hvbm9VD2D84t5w
Y5v0eq+9HEyAnORzxw22yM+IbYcHcHihoiw3IcAKvk46/jhiBGU7/ahZQaEIr5Ee
JIennQiTswHRfkXqGT22MJcZAqhy24GDI2BLUnHUeAB4vHFn0/gGV085uFrclgNm
dOdHH7VekubS1M8mHjDTdPDknYAgxskCkOI2+NI4OQ3h+09+tf0AqM/pyrMUB3E7
vUKRTEByFPvjEGAUuLwMAQiGZlrUCwjs7eEjyy6yGJ4JsCH/G9zbVzLziq/7CLY/
0OW7Zi/cNB6iLfiz5VR9rV6kMfDr0uBpufZqZXnhWghnl37aHszHJmXW/SnuqUZX
q7ZdRYBI7yDfyx3jjLyQik8m6iD/f0glO9iVvhbX38w0Dso2OQs1rOUojONCQWg4
KLrfKoSWX5Z3p7zgnoiZhMIK80XgLu9/8sYLzYaq/jRk2/uJBHQDNc7+TcdWRh7J
cdlYL7dkzav4ZbcCy8QizizuEzHjpTZo3op+lBbMiiFpXcJDmb1RE/ipM89AC4Ix
AWnzkr9RHERcI5GT/da1h7AWdIED3e0wsmmmtwUtxXWKt2Zc/k75iOa5CkJeC4P6
2Iu6s5SwvAvYIxfkr11dBxJfsTI8pkP/bT8GHJcU5GfJuP7Hdey8ANJ6KBKoFSX6
7G1N+lj7nP5PCP71Kz2/IMeLrOqymc7q+c5c0BNNsSfSeCke2O/+W6FvmzdpiNis
QZ78XGVG1gYQIP8NzukxECJw69q6E95sg7xtrHbPqF9B/nk4QQfkllnafobrJgGy
yKqMhXWiIEv/mTkp73ybwCsMJdHFd6qgHT7ln4zbbVxj+xoRinZGlivTd6FWNzBw
agzICqPi9eqWLA90Ehu9pyKYhLY8sELzG42XPS9c1z2jzkDuNdyzLK8u74GRTOuO
0ozfpdvtUdN0FANaYIH9c1DKm2J72exzEjunMAPLoBDNL8ylbR8laRPWfxoercfO
0vDgC2Z+/04QeLOnx/0Oqm/C8r+YmC56jqAhCR6A2ZX4Oe7z1dXDWffhn8lfJlcQ
puxHrwSqdKAQhSH/UZBdsg9Ijc7GcC1GzusL9q4TBa6Qcb9fMaobpT9k9tukDwtZ
kX44b+ah0xf745BuYCB3ETB93Tb3xzk/z/3vXORgQdwVhXCsoKAMtGSGYNw4Ny82
TeZMu5emXRlCTwxYf7ICF5DbTZWLsOA3eCXNlTCq9jKWI48sugrWSvqloks9LH0o
IJ+hnDG2mKzv60VPsBYY27+5Lvpl0fK/Pf7nC0Uen5/n7tOjTS/h/YfQ5nWMi1ph
NufF26nXeHLNqvUHdk2zjQnmcLOLe4jYcMlNoz19ayorg6mCl99MKjtXg6np+X5p
1S9R3vdwslyCdwUCiVoqSqCKhiIJvzixk0VbASxs1jr0S+8NICl0q+qDO5+wQLjW
8oSTn8n5cbe7fIO0e9k8Oa0iHOJHreHNr3txiqDCGDQXYkm7GSD4oxVcKp0IEfGk
FG3ZQtQBTV4x13eBsrHoxH1upkNt1vuH0Iu4+hU3f6Sts6+fMftBBFNTd+V6FRr3
8HqO8EG8Wo3rOcpQUWgh+JFJ685fvwiJwIKIhVNEXQR+If+nN/wBcnE36r+26ZQO
EgssKvzb/jAxMw63GCuuKFzM1tuV7dj0nlquIrR13fsYnc7y8ncGSWEVDQctCNmb
AQMtM4vBYLkPHiLsTbCJfiQ4IWIR3AnpODDOh9euulnuhH56bQeHryv/4BUtCCST
VLhXvbeiBpZ3rdQd0yTaOZW2gLUhHTRgUO4gY06cK60hcg9h0fKYQLA50uO7N5p3
ECya2lXpDfVKJVxO5mRKJTR+Q3Dykm74ow3iH0JZ2XMEQrnglmBRvmsekl05zTg/
MJeEQObQrC6Aqgv04JWYX0GiccFIr3oAC+1e7V0TW2r2jRLL/kgaiRk+owcAJ3hM
OpaMSf+9L6gYiKYxpU2/cSqz3aV1o5TrMUnOJy5mjw1KP9Nxeeyreii4Do7WQpeF
ANYOScV9nqRf+hNODB3icmbJCjPJ5S32ZyZx6UO3kQNNlNE9CupIQlS82gH1Zj5O
x1PfeNq07Z4Oa8IrFK5FqN35gq/NuiyTxP4biZ0C0r1EB5RPvM3JDNikd5Lwn6yw
YM2itaYUD17DWaAyGhG9wPQVVV97GmCWxPhSZNDA8u61bCaxAfgn/giJ+p4lbhqP
P6OtzDziWYIMtyJSoWL/FBVmm61ZUB1fH/+AEJY2DBIz+4DvquOaS6AMDIxwuCBA
IG3WAJVauXgnbFAdL3+P5zx/+Az8VC1eCBRQvagIYObxW2UJMMwyyIS2PnW1mK7E
B9v/uLHiTBnV2S88u4VV5aCGUH9HsKIcfC2IYDI1kuUtIq26YtsYxXU63I4EUC3p
Slf7sdeaQEZVCQBxQVwHpRrsYteuRxhsOTiaNwccNyB+e3dG3lWf5iiSRFbpkwhH
snndbEKxxTUuqqKHc6KYP1f8UZxcMPmwnB8divgQik6/nQ8X+Ij/E+j61bN1qx5J
k171hSosmJUoWFBeH+tp+hz6YsbqM60xzMPVKSfml98buk7k9QYTDuLV68T41mPB
BRXqvW7jHeudaYBqQm8xQVc7RPIYNpd0h6DsXhxjwsH2xQC1cocxAdIKpqTxMuSD
+FAt2oViQ0lZgGkoX3WlwN+MNsYGHk6PHaH9OTUICS3XJkD7rX6znq5NNfeKnhNn
4pBbQTtx0Thtw+mfIZUfnlRLJB9JUXQDZo+ZClIt0tk8pUGZWnfw9jci6uirPz2M
WJ9/E4sAujdfOGFHh/ftjCTzRI2sqv++5oSEJk+ExvroWXio+ToCM9cW0HApaO0g
uN4Z32wTfNlWyDAjeb0F+cfJlqC3EOTbumK2o93mSdBoD5QuTmjbbHLnrEsm4LHn
Qgr56cyuJdnF7uAZBB/6j4YoUBVNiurrL60anPOupa8U2xYQ/ywAu9wJ1GByBZl2
3gn1c5gWOgAGtC122aiQxfuVldhtmk85CmGrOUCjJOwSpjShw2887TWgG9jR1fnc
ILSJnOG0VBdx0iFlzTtX+FJRp0sUx+dzPejBT+gSPn+uffXSCJfhfylcISnpCmJ2
7pHOaA8cHDLsCKeCtpa4vgcilQz6oDgd495Q7k2f8c5HKvySDCBMqY2rbYAV5CzT
WVNz8Pc5EzTpskOQmGrZpmKx7lu29VOZu/A7G7ayFCI+FkYkflX8o1wHD9popOrP
YfKWrOAdZbgjTjqHpCh7mEUiHJRh6eSgML3PrUbc6Mdhm63ZzBwMCK7HNgnjuufg
hf9yDo8a+dgClgrZluJizPnI0TbEiKaLhPijNX/hL6iBKFjwjx51X08CN6tqFnjA
evEYfQovxT0jam24ATMR+LbkrZmbHQat5YN9hmsPf51dJOJgK3+y+JN/z46wIOQ+
CkEJ4hka+NtM31bu90ALiA8+18w2+xaXD9IZcLatzjJS0Qe+rxMLf1fFnB5uXt5y
4RZEUhPtD7SOwFRAVq2C++s0IuSBR4aga/cLFBArgV+9/0UP8kIPb4Kfq9DBT+SA
u+GOxhzVmF0f9q52OUUekfDsctb1yDQkZ49Y7iKB5M134TkTsJx9Q2gUT56DlnHj
e+RSuwnlV3C6AmfpiDNJQLbB+jvUbRxMhDf6PqP3fLsEbNWvrY1amOmSwoYeleAc
SLbER72XjmJDyrn+Rml8c/lD3b7YFqGO/psYE/pneZAbS/yKbqblofucphidxyL0
dHbq/I29bOkU+86zMGXl/fWxc59XWwsmoFf+rNQYo5PfN+sn5huHKQYMa+FGpIL4
vOfulzFgHcb7mix1f4sxvgSiA+83gwFLGHTX0jhLMUHhiYYv7g83PlSs9jXSnBjy
nji5532IQBPaTLbvTs53hFL/4/ZCAssWIsQTpsYzfVD4co8Re57i14Id4ToS/blv
ycbq5xCAiz/Z03WDBmaU1Y79QJhUIl11KcyzKXHd6uryFXwgI4RIIrzqWZDqXL/U
1A5MiUXFSFYD2vrB35sLlC3FPpKovP2gXE3oLyMLaPQvSmw5ZNpdOjtFsHahDVOn
i86blij0Qh9eqmY3vVNoC2MaQ+Q5tlxMA16qpXEBN5haFAhTluwBdtjwqICi/ms8
6cK1f++TmARbMXLTicTFpv+IBi50zxmLbgWz91LI+xR+Qip1UJFPgWYR72OzHkmK
STsvVXEar+lIO7Hwh+q+MZw6kGX69eIkRLzqymgzNcFXP3lwgbvbdqxpDt4oVQcP
05gOh2GfmqDwpASgCk3GcFn5MGo/33yzkSUIG0+VRR5bAT41oUMqylqgLrp2zP/S
HQykOc6okEAgJhgZTb8RAZq3nYqaCpI5oo55CMvcfW3C9xdtbh/DUoPWbzksPx1X
w2R7U9zIYew9QQlSFVZ2FeO9PTNMYS1F56mqgE1oEY4qaVHEDgFZxNK7mjsP9Hu2
X0E2iIpOHcOgBnqPBFULI8vUpovXwEfOZoXxuNU2nRXbrn/dR+dNZ3OxfGR0gzjG
RvbG8/emSftIOc0IlLbM0PlHNy+afpv+QccxaNim+/Cz061hfmXDLGmjrx2mUe2t
CdmiHFYhH5pIRmWc7dwu7nUOXqU8qFuJ7J4p0dHZaFXMAObVPAWkR73nSMEmhvMy
g145Z2oHgOA60pOlvd5embmpm74eZ/J06jAz1VxA3rCaTK1v+g8/k7WMmeIx92y5
0Rq+k6QHqoQC1i1d7coYE/BlcANN8u9J0Ocu+Gzz/KcnOAkK6d+rXCl/7ytRadPi
6ktl3lkR6K2FpF3Y5Wae/uJls0iQwB4syt8J4ME0UAsfIDmUS+5JJk2QMxp3TdJi
bT1WPnPNrOioFpuhW63Ig95u4J65airmzx6E5355tBzrPYrLJ/ynGCbqtJtPqjKZ
XFNNFdcSBet64obWMaxHzMfKZiCQ+19cBmPVeoCK2xbmnHw1Fkxuc9OGP2wNSM8e
+VhD3Sdb9HaloMTspHhn93nPMfimFajIzknDvM74FMQpggyZO1Xdw84N0jcONfaH
0gBjdbTqh+yQvZK/YZVh4xmRjFXnX4twTJlfePcuAqNtW0x2BABEDKvvbevXAa/l
HDVJsGtopG+vzUxAHEHaYNQraxXewgFmEKsn9YUA0MJ13Kzk5EMKDF5+pl/96Gqk
2sTNc9/jz6JY8MG3R3Gygig84ZrapapktepfBbVHdEHRw5YTuCxaKPZKTO/FTTeu
atHWMC0bOPWNuiKuXPj1fwkj9FnzuwXEQKbfUiUun7VBokhKy42Jf/WErSCbJXgO
FyntzwCnl1/2LmqtloQnUs1mqMklc6R3siVjSctIZdOUvxuIzAUHgDBm9soWXC+t
B5LSvUIroUinZdHxYh2HABv0WmodhtgDX5f791BuTuc5GfIvk/NLsbtb6aMrpoRM
ONp2/U5iSwa6b55lb5s2OvS/QuvfepY+SKRI+dxwcGvRuSgKQ24aYSLJfZbhSoJ+
l3aBKnVzP9chbfCxkss7pwm/XNDyVxT/lgpH9hgDC3V42cA7lXHLsyiL465C7NC6
vwv/MNpp9kUZC0iSlrI8Qxt8bLsV9F3TqgIV7MSc5gqiHUozvpMXrafF691It1MN
SoVcda1KPAmsjq72Vfu8gz82XE8xwx495kXHQmayPvLzFw3vQXvwOrRtMlqAUI2L
aQtdYwKHKBHo6bGyW/UjiiD2RMD81+8O9awSxfYShaYj0GFpx8zI4w+S+moAMFB6
/JlCkOJystObl2MNAg8TyVmv/Akk2QXAb/xNR1mFIhWDpy/Mj4Wu+qbZqLBR48AJ
TFOT+BqdzJB9sEgEvVKb4gSaN1IrF0ppH14SHfoIld58SVkeDTTQzq9CWasOaPLR
ynPHHmCVcyyYvIhJd3+lsmtcHyV6X/WSg6AYv2DtBaIVxvlMIRcuygTvHRv5EdFY
c6TSi5MOSUuseRCMEA/ll6nsIBTD0fR1G76WMtLpXLwHHiVKZEhDWrentCzyP0TH
jkOmDE3l3E+GF4LUVNHLDYpGCmvRaR8OIl+TUE+1tukssSa91Gqm5P4bu+Tjm7DV
AGKe1vH2EH+AErm4yvkSeGz/hBMMMToo92ERAWsj9LqJurUnRpG1Te5DagCrFwQ0
ExQL9+5XBObQHELUXBEP4SvJvHzMlCZ1pCAQ2jwqNZpMk4GfpZpqS7IpOLf61P/Y
CXnG5wdmRB4OewqgTzqF1CusWlJVaehNk1tEc4IgJxln+P3lLHetq6HFCep9Vfwy
iDV76qkc4tD09z9lIilOL+k0aEa/HM+mcqBX5BMrVw6iLHuna4Gabp2k4kdJIrL0
+XRq7LsXgy1z+aBEAn3KTqNLs96WBo++PfIXPl5pVmVh2MoFnlBY96NWLuVxTpZ1
9RKgx6PfAF8knGMWqIqm3pWRMlTwntEZlOgxZSNVYcOcr45iEKram1jbbJLLaTTf
2NePnrestab3xSqlibicDFzreHscYU7tTS1MEzCJxHL6/7jWHPWwA7E1ZPvE3cpC
CvFYCFYXbcwDt/OHfebi37c4BYFICsyEMmYa5igyJTJ41DtupUkC64JEHrEieECT
LOFsTFX/sEHkPBHSkSFGHk0l8/stJXthvvZ/smK7+p5seg7eZSLKV2wSguU9OX+4
PBeWV4QgRme6tvx0CZHVyHTnaYbVkiqHfi1QyCtD73lDdBK1eNzPJA35Q9tzacQq
NSIktw+ryfLdvL+ObNrYxDbsPv95NXSpUZQZqv7yXOEk33UZtZ+DiFf3ITr3PoVD
hRmMjeAyG7/atjLVW3IuDXxKzG9XfOL97Gov+Ro7oBOhWYz9NPY+LMkd7VR6dfJb
44Ug25Ml9fc3fWczVihPwCxBVZw0kMj5Nobh5tSk/WSkg/CEO2bNj5nHVEThH8+c
0v99BBBaNFFVru6XIcWP00BIMVpkdFrgpjAEN9J3MbsqZgKpy0fwnPK27te5oWmn
J5UAY4Gsbt8u0VkLfsAaxc8cXDbZTgCcQ4vIxDsErNnEKBN/3XM2n52RQ/yvV7Br
o02NqVt0m9KUphDfU1K+Szgzuenpm7ZjC9tApZvq2HF89ZcrS2fAEftZvJz9m69I
IAjJXOSq06W8QuUOAK2D9YiEE9hlR6pLPgpCraipLnRBeTOvUkA4pNbln2NCLifr
MUkPC4Txbc2f9YKZZUkZ9V3ys3O7ot+wVi8CfwrpCkq/rQhsT1x6MH+3gyl/3/Xj
HC31VGreQXNxlPoSi39TliiFJAB57yjyVRcATblOb/2ftK23rfeGtuEqrr2mC0aF
pJ1kTWbX5UA6l66tF/qsHotMJ88QVfd9CWx3e1BxgOwhXDuDa7W/+D+Wm+OdIKp1
eIVrEnwTLqrqNFGY9DOHIDvlHyc7RAC1NCteIKLiWuciabcK6MDNo/8yb6MYQHik
d3gZgTBn0XKLNy6QtVrA4K+nQ28i+Wafmp8FEPqDdRiVis/jzXEqcKe2kXswOTHJ
K2eH/enApqPQpQodrduMCE3pt06dtVIomd+etIJ/crq5qqhYzTxPKRX+UnFksUUD
j9lTUJXFnX2aGK56aCCNtG+dgWVLOciBjozAyEc1UQKgp4AN7MsI/WYiaxrjynCa
2ujabYfqFcqF79haKfzb7IzRy6gRjabBHk8/M+V7QCFNOYkJNl6l3tUhLMNDxn9i
9+IhNM5acW/f/E3mN3uJcfL4jkIZ+U77U78KBW0NYz7XNOG3aN91ITbxVYgri68b
7NL05jDl6yu67iAoRbyB8PSlyYKldGcJG05D0ypS3xqfmvEgAEpwXxbGLQlJo/E1
iY/w571zfYErPnepAiC7LbTYg+lfYJXZY/Ud0Ihh2wK1scS6VcawDh2Y82S/YdlE
AN4ep1F6PACiRUZi0BqL4TDbIhXOy6GXljTW9UyHOqBqVVbV2a+GqnHx9HIQR5Rb
Z4KF65mT5Yo+kxHjbB2Tukcl2KEJdUeqApEcc2Q0hj1D/jWwER8JMLSAqEEs4YHj
LnyRlYkTXXZUqIyjMIS14983lwxzuxyG4A6CsPpWdA2WvJjAPg23nkbQYSNib7tz
WLEE6ggT02kiBY2IRiDGnGRX1sEkFWEThFTRJW+MBMjxuAJDMjOY5m3e2KNGEzDJ
K/gq6w3RI9vhSV9rY+cvEBj3dpCEq6u+Bo79CCLEI5bUiWIPxmg44qPA8KngqU+7
cUXTMI1g6M7LAU7ThLKoq91crGliLesYTTFK+Jj36MOEWWYUpTBpu1wgyoUOpybI
TT1qd1iFfGaFjTT27gYQzqpzOMe2MUXAyP7jLwVycdEAnnO4jXRmEcgzI6/0D9DK
8ttAgQu2VEpDVWhfyd2CvXEeXbx3iUamHoU8KY/MopmCqZbnvebsOxuN7MKzoVC3
gQCNdIGMrrJ5wEiVhbj1rlBVm4ech4VTX7oWrrjaAFh61cREX0UEG7L8tJfUqtXs
VhvI31mVHOCtZ7tDxu4FSoJwTobNMCD5s24Qte07DeeQvO66QJbjcnvdHMTr3tbT
Urcid/hQRtOJMLV3VZuGjjPtE1pm+2/dVcSCazS/sNhlwKW06K0Y3z5XVsZOhaJl
hKFss1qdS0H1r2QUvL9ERP3n61lMCLvRNty6Utfh01hMj0MZM4gtaeIMGL1x1uFY
mT5WQoBY+7pa5OL5YvzCgmi4YVZ8r7IOhk7fflWDN/pb5GeVgyPZDl3iwij80knS
ceiP41Z3lSY3u7LZnAPzJVQIkHAn9hq/Hi575YyzVrF+erFTsZq4bAzNoulkG7oq
eLdqxw5XEFpaxpUSYafw+HhSkUpOmEbHEQZaiksaobswNpDZj6YKFB0uE2TJBmbh
vDA1spngQ/9TsdbzRpRzscghJ45PSsFWeLAYhw5H0mkGxr80765s7ibyyP0iR0+2
Bm6H6NVDaaVhKxdFcf1gfduoBiuWBtY27aPEjHy3EF+D9Am63E3/vPia8jGMWSZ6
133vJy2lVtV1h70P7gUi2kNfvM6xjDuylSLipbtO5Hv98EP1XyxHv4LAr0K+GZQ3
ShKU7QPjnxnxgkg0ngbsxSRVB/sT7z7fBjPkb466JqsSWWLi9atnmg4B/eihyghz
WagaHTsONeJ1yTHbiyya9UtY+02oW+N7++r/zFyHflilPb+dmcF2FhOrZB9qlAjM
RqNWO+0Z8/9UrBQ2cxLYJh412G+gaCdzy3vF6t4QDkmdc//jTWHHHErqtr6yXckD
IkU54WknHnpoCTrRXUwxBS0yVFAwIv1deZfjPIwk1lUKOPsWpgQ+qObPTGO8sdiY
xNRYuFwxwqCz9B05C/kXxe51EMcDd+5GO9pHwFz8MPSv+RJCSK8B4F/+Iwz6vLb8
+N1KNvsQZNLg0VejKa6iz8HCx6wPpJSYPlhFgl51aev8iozNBOt3FxGAnOgtcDbO
Bj/1m+j11rOoX8TVpjvYZpt5Y2mf5uBL4LhGOKE3br6jD8HVLykHsst4I2KiAaBQ
FamK//P3jC6prfPpr6dEJiZJiO8Btn6plemP+KG3394ZRlV32QQqfrt21MGRpwdj
+5iZlSddWcxIemWKkZ+xP72kwe39NOk9rks9tC4wdQxaoB2GX7Znf+tBfBZkpw0q
Z/66u/YxGIyrudqLY1Pq1ToG830eNTt4ze3w5+z74WUV3wWuFt7sfb/NLXBaPBT1
7DjNZ3SA/krKi/RwYjWLNpKRcUfuRjywk12s7q3eSC6Z5sb/evpeE37OQchVejBG
05H3iuCRJNQ3NziKR05TpikVNbq+HRdLtLeg7ES98sjOaynaEpjLHZ/q7HW2Q1gS
Rw/UCXY1aCtC4DNIgBvkbLTJGDU+Iw8zgoE6E8QJhPfiwMk5WvJgI4wAqM8doN/m
Jd4lpKrOZxQOTgB7bPy9dzKR301SJQeBpwe9xyE+Zfsdly/fkEKS8DeUxr/bpdI7
HEpdyibMrsAA0RClGmDEe3OIE4fV452LoYxFYWZn5iNk20UqiJ4StuBnPr66LHX/
4CEfI/obMSniRJDb5mKHbyRuPqSdDFfQ79K+A+GgUMMLLsPs0EbpHGYr2lvFcyGO
4V1LKNM2JyoV3+W6wEkq6IEFBRlGj/HQ+LuWK/Ftcq9A1YHdOBuFlzMMoiaZy7w1
YDqJr09UcpUZRKmEZVZ9vru2NoKDvhPfdQsRUW3MrQBUEhLZhHbPow4WCUCdo1vd
+YrdPsyAqmpg15j8TSsgLjuknEbacG4n7ttaW+u2Z/DH5oXFpCEGYyGmnyoYZZgw
Al9hFZ5HyUCIPWC2Jo1d4MoHk6gRgCIrdHrOehk+HB1spZxkpB4QJ9A20/6SOD20
AK9mzXc0408Cy2xM1bRzt3RiKMOrJy2WR7C3yIw5sXfux2CbHJKm71gGQeEt7yBz
Gaj/thHHR0u3+iXAZu/G+cuw7PH0TczosJVOyihZK3h662OLGNvnOudr9Z0Qi5XD
hTfF8hyKoRvCkhnlzoow4pZLEOWlGQ1jAbOKk1f4kuvozsOiS3Qx4Y1pD0BIlVG9
RanynnHa8/l9QGE1T/gTzUMzlWFdnYxFSqr/MfIW99oOwg+xeTcLkn+MXXx4SVRI
r+K7Yi7Cp5Xs9gOma5aJb2qWEY9Pz/X+BkxOWzRA6U25DVKzqcXVp7kaftr4n8v3
NksTGuRQgSn9HnMa2OR7fnxu5BRWpQoDe2MlH5mP1dCa2CCAbpB5rR5NHa7vWpLN
KAEwT5mpcFPj8UOvMIOAdslxLvi7lQQjev93cipd5eKpn6X5M2xsoHqH8oNh+4wf
GY4JpvlDuV329gRwK6vwIoNqOhpN78MjxY6OFn3JUhNHSNaOY9fFH0DkTmjr+TFY
CpbVoMdyhzYx5hY7X9kQcIysXV/hb+EDWGek0yA/SHusBnOszk7tqKTidQz6Zduk
xBpop0XfzJXHzI3KVwR3bmyAmEsaLGRmltJH76iwkICXG4Iaomfa6Y9sQB67UneJ
kBvj2jsj77GEBbtkxiFW2i4dwKC+RKHDQqW0z9uiy1qICv/+o5qUxPoD6o1xFs+5
2Xu/5kRBFlsvOIvljcUpNnd7sfP+wrZXGiXU98P1U3myHmWMDjcUaAuj/SrLL2My
AvfLuKo4jMaJ/94amKlErjwQDApgBgHwXbm8SaJ1CxNjMdbVCJyj+YyAfU9X0fgG
27waowWw8SMRUOMV9wdM5UV7CLDuIC+6DteUfINY4zq9Untcrg+bDsRWtGq9dICS
/8VYg9s+p6Wba+oPUnTWqjdWap7Kf3/A5wQfDaeloBHiDNsZhLzvQTt0w5ou/Eg3
h+7WdSp7qtXQ647SnRu9Wc537NpuVdQOY/IZ8JT6bhdQAb1GscuKW2MLWusuSS4F
QnYP1jr3douTi51cZTfDOuo22XhehWMvo7uP84my8G9dSGXhVVz4GoCOrmJYGNX7
Nj98kI8QhkqPeVdqD8RhM7BV56AKH/0i85hQLuIpiBCs+9aE+mWeoMrJp8AxjRyj
MpzWtds8ZyLc6IYn56oLG+rtnFu8PitVfyFAAhhXcSOI/GUf6MkXHO+i6ZPB7dHz
lRjtSH1JoyI0FoYYoaUOaKD4uqQ3Fuv4VOP2nLK84JrCHlPHZQuUwdPUYOA6B3wQ
b27UxhdjnyTyl0ml3j9Waon+m1ooG2kVvcU0P1HSc2unzOxmeB0Xob9z8HL0wWBn
Q3yEWGojs4MKTT9ItGBt4j83pIsL4m/rD9FBKGgHZ0Uj8lY43wmmp/bOsNb2VtQl
vumjht3Bu6oDUuS4P0I68/WXqtZ0ldeqZFZaul1diIkaCI5jlyfynK7vtRJu2Tc9
4QXV5K5Mq0Ji6ZsSmbsdhJb6QgQxGnCLUJn+ViZAbPLHnZMnTy7JpHSv647PlNx4
aMe8FS9JNBX3TgNhSq/MfT9JqEFv9P8P1sdHnrSfNL3pNAR0g1+D/p2qZAeyWk3W
p8Fonc9W/Xrv/jSED8eAEA==
`protect END_PROTECTED
