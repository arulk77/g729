`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK8MKyj+LWN+3z8sfjDj95j+5Q+FWHOFmfFUURk3wrnz
TQo0cbHyHKFk05AwIvfo/yz7addMVvDg9qo91xSBvrzdthNSBl/8N+vI2kILJh3V
KnutXfQQjJ8OEUje6KdZdHPkCbFC0frNWie7FlNpp8wndX9rdx4QTmuJk0dYGpXa
gcbAw83lCy/SfSlrVKdLE6mP3ruhDuV+WrrEv5gbbTp/SGJSM7wjK8OZEmlzYB7h
3ZUvG+rHLxg/f0SlA+chNUMIm53pmcegRqPV/Gl9PmcCSlgP+LvRBNvSX/aIQAGf
zLYnVWXZPP/k89DtmvwCpr3eKmgbFTqwGGXvU2+MPq3ZCKTsDf8h04U4eQfuKD6l
p7COHStUYL4g9ytaczQVCDt1WedMCuj3SBjFrE+b2VYz5CCLtnvS1D2Tv9kLuhMt
UULW/6MVLeUwlk05s5xOTA==
`protect END_PROTECTED
