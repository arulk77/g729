`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
XXQHxaGvAIS0H8aeAYMU9Qmb5Eo7FemW2tRvnrpPodTnwQL9JWWhscsK/W1ULNC3
yv6inFosUqwCuQ+Tm6t2ptT7Unm+gOnYXIY+Cm5Sfef8AIG3exftZFYD4F/VCMxV
AY0Eka89xjT/KgLa7n1eBwu4vVzkONnwAOlKcjzl9oc6kDNFXpk9h1/kHdHXBU/E
`protect END_PROTECTED
