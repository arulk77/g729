`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKzggBWSxrmv2RBGEfLKNo4JcPSn/2pSzUCEDRbHpYqj
NvuQCVUA3E91f1mLQcwGF0exsjzCTH2VOCnCRe+iU7H64d3j/5iMKeYS0PT86dyj
H8c+WjyCecvGBxPZPvglOxEknyqALm7mN3XuwQH+NmGAnyyb5/VmgGMGMBkJGbh2
Ve3p6uSMi9L2E6EXrgMImFBUNr0GWnggYvAq/ep+5kUuaTs9WBMh+kUt+94U0QQV
33r8NfGMLtKlWrdosqn8pOOF4gFsHKKyD0oxtRh2ijuk9s7gNnYqay4gWhAMD1OS
/AQz7uodKaoMz4/nyHGC3//13M3V0SCUq1DgAHfPgqgPiaeu5ummyBmf1QqLfSV4
9nosEjelIk4wedg9EHIzI4gamudpHubVH+mBwnvm6mXGN786aOK+ghS6HdZmXrx1
KrC92sei0ulo3lbSrJU021qDhS7yBd52X0D+zGXMybdkvMqUUv65qTiGHz2Eu+1u
TLJzdo9MO/BY5LoE83bfEadhyXfGJNKOeAm5x+xzVgY0OM799M/yN0ULuK1zdsNt
`protect END_PROTECTED
