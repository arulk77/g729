`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNeblrSs8ySWPz8IHO9lEErx0Q20lClhNmnZgbab/EL/
yJVj9LQe/CVgiOixs6drzvVJ76bxyOA8dFTng8nx/EFbvahoAeOUwvz83Udql/YP
kN3pfqF03BnN3dv+5s8/9FWUCnOLMzKEr7z2NaMvek3QSRt6l33UlPTBr8UW5G3L
BGnmYJeWT/YSw2VAQgk1kdi7IUngEYOCGfWlfkK6fFJ2iPZlzV42oQC28JIxnzxs
`protect END_PROTECTED
