`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePNdKkbWXmLBItyj1iRtA+Z29S30jW+/8QR/E70ktXxi
4P0i35qSA/dbGrVs8g2JMUYcPti4EpG7MEN1zFQOIePbtVE7FB2AdlnyNF7opr4F
4FnRBemTpWoi4WDuTTywfY+JauV/IOobY12a1s0DTYtl6ydFIJ6tJAOHMtcOwXjR
bvTJ6/Wz4fU71okGCYevaw==
`protect END_PROTECTED
