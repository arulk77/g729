`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
LHgk99xVuUNemSxvNoiAbebSBjdLnEcc6CaCfg/oPVokeqkvq7xMlLnG/5JnDVUG
KcAQl/KBQjYJNrDgUCd4xdDXG6P4tcB7YTLcErXIk5pugbpW5PQHwm+YGOOI8jW7
8qUZifw1ofDoFysdsPqzjaZk5iGGMwnbm+uZFx71Z/ad8G+enlLoAEmPkFD83C5T
`protect END_PROTECTED
