`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePiU8UB3BZXgz3Pk+TRtrIiRK2nFGPIPY2kClGxrZ0ej
OIcpbCpXtYv8VG0Hll4pJBbPZ02iBFagKIyTTkbw4ZA+gZv+O39PxJQQvSCKs8S0
hUNlurJvNIsrxru6NRM7AuLqfl8WhRn/Vak91i3S/JW6suWiKW6QZVFrkibG7WSh
HGmyuI+w01bNr/LN1EsizQ==
`protect END_PROTECTED
