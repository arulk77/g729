`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2EBoZu9tBf8wFLCnm6xiM47jcfMNPVJMTqgkCkAEvvxsymshIxk4CBze9/9E6GyC
kRlmjNzn5RXNQHzIkE+pp2ZlUE8BdKcFLVANsWO9DiXM/19kwx0ZbjprBHz8bixm
qJKnhFgLvmW5oL2Z7NSbT6FVaerRc+WBhu4X3fV7Dq6k682752y62ZaA34O3fwi1
+YlNatml9URyxeuS2iFOxd8cL/KDY/P1UDzqTVLW5sERkrofq3dsF25oqI/9bxRA
`protect END_PROTECTED
