`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4310+pVe6CsGe/ogWmSHXwADGidCm83bnEXRHcytznnz
xSCpXztuPVJiHd7RY/yczriy/KR+qNKiOYHfxn7GU5VV0QQJkEMZRJ/ttjI4WdVU
XH9HqbgPYBh6HgNLYp3lZl306xf7IAxuS7QErEODVkg4Tf/HiKJGeFHuGmX7O4jK
JTkg8amtVIA7kAVpTs3+QaJa3iT65LasCYds2R83b8+vXdKFWtiqwBn1A0NkiiFg
Va2bKUS+0m5spzfOz2Rb6EOb06HPxACgBFycq42JkWSmccCKn7yQgqpMwcGCVukc
KuSxAwdBFRKSuIhddXcRWw==
`protect END_PROTECTED
