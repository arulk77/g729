`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47SQw5q+/GfWuhBFkIKLUiSv0m5tdQSOGTsVU7EbN3lb
QqjRZ7K8I1YNXEhIj42VZvJEEoK1rMA/LNNR815d/NI46IbjGpOVPNVdbfAwRru9
VLb4/WDe6BI4z4E38ESpim3LxLn3ert4xT0eVjgRNv9JZTKPT14sNlU4uzGVRCJg
AuQt0LCYAOhW5P6beAzz3kLLI7rCZIF7rEQPQl8ie6EK17PeBgeKA3TNUdCNigBl
Hcg5LsvuA9BClwQb6EUWNKBrpuQC4r9wL97AfR49VigK3hRvNHaJW+3GZWrrz8Hw
KO/ZhByzRdvXYe843HVfEQ==
`protect END_PROTECTED
