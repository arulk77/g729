`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
WMYlcA3qzk1rdGOqyiYA3XfnmECxe9qryh8Z486ecBl9AOTK+AWbFWWDH/9ThHWd
YeHFVP01B4X4Ys7+yd61xJz9GYUC3JumOhLdtMqz6yuJceJHBhqFQynNxcCDpmm4
Zu0233tYaF5WmRzaLb4n8nkIUeYUtUmkYARRe35GksciE99yayDSJRnqg9zR54L1
A1OTbmS8TzmiWJnvkvy5ppZpmGXTQ9LosTUmomohJkuQB6FpPK7wGlhH/nhLlE08
053iPp9zdW3UxDEbSAc/j7Spf8lx3OLAzSP6X2N/BxcSYs56TkFTHC3QjrbBQc06
f+HHasut4PJgRYnkG9YTKeJKqXyM3rk8ax++ixCt/w9OCdePVK4xpTkDMHc0PK/9
2pFQ1Zal+6lPAQLkA6KMar6uFrMeo+bqEGYqtmGsT/8=
`protect END_PROTECTED
