`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73CyHk9U+fMI2fkRjXdCcRGmUdb8rAuyPkVRUAJjtKmoFg
pczzqyUcgJPEa6LSYmn5xxAtMHkDMfeId7tsnxXgThj7rOrfr7X0mLA5YhwUpNum
nzyAVrT4ScPPHqJUUnsMapR7MRZvQnHxTBmhcxcBvbQPlVZ9dC9jIoHfaJwlVisZ
a2blrGkNE+PK+JZGbwDINw+CPknSefxPy6Y6/C5K8dRxH88H5Nw0fTfsEWTMTZQw
+MVFRE21QSSapcphC/4Eoro9l7BbuxLP+zREWryYIPVbbOi6ycJivd00lYcDJr/R
xcKOhkWoEcqe/5oMW0mVtMNzeH7T13N522whAFhOKK9A3icxPRyHCeyMH6iUU77F
TqI/THYPs1cLnfj2NgoJwV8wlj4k7v9CI4sFrjHzUEyn/Hz2QctBcCY3NEqUp3ZB
hDdjQHY584ivQifOuUs/d0JD8WqCjwMkSDGI3ELISYT3qbs8hcYZgDNJbvbsq704
3G4vm43DeaZMnPNY+RJcH/GbnwBu85lzE8dq3MJJF4emOJNYd6FvmU+RKEFdA7E2
h3oINfpu3KhZOPiqbsP3na24OMMM0mWlpXWQ8a/wmn+luUUSQkcELZEffm8b7Ds8
LEZUo0/L+1fbIzClux38lvoNhswBeTp5nZOgXeCcItCOfp7Lg7BHisQwTECmhjfy
I0Gj8+UpLDYTWXcHz2SYsFSyApjhlKaK4CMkszpaf0M5OsMJVv9Wynp4ix6Xh90a
0N1KL6oKg4uvRcnvEL/VB/p6HXZG82zIX878lzzl7TWgM+G6pEg8sLsawwWG7Dfc
b022xfonm8g8GksHZLC673oJT/gY0+OtAZ2tDNE70GECkkMmCLPhDS33LbBvIaPG
kG1ZyvHCLyWnB1je0hS3hFdnAIu22iEM5WKz1PJFVU5387A7mkOf2xlVzKaxh4o6
9G1Yc7HyQQPCUbN16PqlCrMmaOrAB9vBGC8G+6oS6AKD3pku1aXCgsffYWzQFlw2
+fOxK/bUdYVjBt6vejVoY7hGNOY7VGYyQ1yk4exDLYgtGhbP0cJTscaM6qYkCUPl
mCkAtOMkNkDZkvi+cICkVSnHlMFVU9HxMGAP6DsAK1TIu9uczv5nbYk/38aukFRw
FSdF1vCGlEgUwh3ZJaosVkmxidzPfBMKfLs+quUWR1HjKBol71xZ14J8a0jVact7
3bsEWzvt1lwOuSXYtWsmMIHYC+Fr94aFu7U0QRjQzAK8UN/c5oKUP8CNdVL/v20B
5VyfVY+VyVUWfi679/ZQeJIiScXp5jk4TevW5CctBp/478eJYJqhJzrxWhLyj8lz
cD8zAZtzgeWP/3N00OxAtTV0k0DffJ67s6+jEHy3C/e9+XyIKyq5gfJQwCyTmEwB
x7A1KqJSKjXflq3OKGOlOSEfD6rI+0Ms9mvpLUr6gWKGd9SM9yc2FwMwsPzrnwz0
F29VZ+82E8VJcmPRRnP7M8axdIiyQ2MWU8+zxveXwubLS4I+t6n8budzBc5MDXuh
CXi2U54Pr9cpkZ3cmWYPoldGOtcU/FeJEGLMqDf/srFFr3O4VswdJ4JdkI4Dhg+9
ibx4/DjMdzz5UN0f144ml5Q6Hl9yEK5KpCL0m4lZQvTVm4W/ajJxIUbPsMA6lj1X
xJ8n92+dGvkF73uULc7lPBgTd6CRE2gJHp5Qa8OZ+Q6AEFbEeEtfc5JrdTMc5UFJ
m5wVBc6og/R+kSZY6S62qCFBpHRxYR0jwxwYdKmd2kZ0+FuZhGy3/QFhnv7qyrVC
PSXbtjm+PD0DctfJZHRM2iA9NK+6ss+6ruzdSs0n8bgDt06OaxTx9Z5dgqaZnPit
UvhDY/A4+U4fwocLnfzR9Bsr+/zm4j4U3wvW1MH7erECScZvzwHOv6Y7f+w2M/i8
1PnGjqNah2jT26f7jhP3BUAcSJmrnmyK6hjdDkjGuSzxpPAbV7dFUOh44gpFKVWx
DTAectCaQL2JbcIEXW7nwr6lwBJdG0E/Uc1NkOrTqF7g7ERy5OHFJ154F9RctjQ/
gHj1NaXTvkL/OwfyWbOsaxpD0fJM6NQSVG2gQyWdldpLbTsvTGrIbTBER93uGwKx
2Ei+Hppkzr1eGxI/nINQ2noEIaKG0izUEWz21zzLtYDeefqXzmOeO8y7D/8n3Q4d
mk8h9W6IYaOgeVjRqBtVN8LeNXoJONZtg3mtpIgfkku7W2AwnwVYHOO9IW5/XZUL
jkz2Oiy+RUeWLtyNthZPR9JGnMIn04Lf9sZTJAYHg3UNBag/DwMyCQ6w40JQcYeZ
1OptSpuRLJqSUFCpoxXiaMND3SYVEio8MojSET1HD4AjKaa/j/yAX447RTpRnhCp
WLxKlQhTHQRTS+6OqWmOLqzgxg7hggeStQnngPz/CRAPHg6iBT2y7zXF060rrW1u
ql2k1K8L30deZTEmCPMBVOsXgX88i+2NMUUJKQzFpm51AHxEjYw7dFQ8dPxODgSU
wri4qhUk8mfNLFdtot+yDwCh77fugnDAQdGnAfssc6qqQZlt82QtiPLC8iLbvG0c
hPy+69DsjVpsvvX50HlPLJJNCg9g5K5KhfivHirbndm4M/mpbr6KRsgbXTx+kJnI
IhPriphdn8t8DOcZ3IkyR2NX+QtF+21nnFuGZBdXcbJhEr4LPjAk2hxGcZw3peI4
FyjVqCj1dsYAVdrV582UVeoMQYp/X5YPsum9gYno5BsMPJ2q3r8x/nZUFGLpdC5S
U72EnK//3NtgQR9C+b0hXehXQi8JHqGAyM1J3exq6kXosCniVu/NubQviB67EFxa
qCwuij0PWUj9twvWIk+4rwcTmpBh9uDXEwtNNOjiSKthQAeT6oXt3y+ixF5oTW8i
LzpfSfj2WEhO8Aanwy0Cj6YIZMEA6gDKTuM3RPhY/MMkIguWqycRQGd7tAdjaXgn
N6lOgewJQERAsjvu+wXPq/UGq/HMxAG0h0U333Yy8we/gjuJx0EfIFH6LajPDNGs
S+yYI2shbkCJIVMTXCSDc9YFvJFw5unPAh2fKIfy9tRD++5DY+anWdmU+uZSWm+p
2lXxVaXvWFytAP2PSkC4WildrGlmSe2QbXYBHNvAhkmKcxZkxQHA9VsSUXTS0ita
BHjLQqayR+lKZ3LWzCALPmw8hS8j2g6UonPkOKLCh/2CPgb4tlV7klKcXoGuGOVz
dJ6Fe9r23oeUH9LnUp/7zy3RnejT5Hd39hSiFX291EQ8YcsA6ARV1rIBcReZpGPr
sKtXwFReHa59m2qvrVOsWRb3DFLrlg/Qhj2CfYW0O9Ir2hTAd5KrSKfBst4szz1u
NQRlHSeSKE0znuIsTZJmkJwfKpT0ayCfGJXmjRIxsocehT5ajlRtJy4jsa6+JKvs
Y0wi3EvVVejDQRNRYQOFO8HJBc3eMevyBk6A4j3+aoSqZRq00ICTkAgIZlM/rQ8l
pEOSyozj+DeGXc2ZdYsBmI0PUUFAAKXUfe20mVS5uvbozYzjUSu9HDtYdKgtRjvo
akj/ZLilaKFlqYh3NXIKjiBX12GN7rYELl9EKJW+QKjkRtEGLOixygr4RwBAgEjS
tQ49qnTCjTAHZJQWXGvnsydAgimQw+gT9/S20DcrQf9zKY1+QBbXc93Mk5CgsH7O
5HjCksJmbqPdwReK8ALEjPo5Wlya/GoPVwWAasHA1Lf3bAIg/ECRlipuRiA+/WWE
h67itcE2ssywyCX67r+F/u1nCn46ZHncmtGLAdjMomndiRHfgLnzujjl10cx0OO8
jDZD2Moe+2kn24Q/BEA1Ku3GChbqQw6XQ1w72raCHfuLPZ9n97kK6L9AkSAjovo4
`protect END_PROTECTED
