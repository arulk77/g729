`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+BO5h+6pwoA/pZQ5OYiaD7fKOeSTqhNqzZKgl4+FcwB
AsYUKCx+fLFGdlc9jkZa3ys2PRqJ/xWciLrq5Z/WBp7oxG2FuZaNk4zb0WaC20nn
vQso7vuDQtWNwz1H3rQPJVLBAsLYU6XE1EIhoj6fheGEX7SmBr7guVNtFlOnbWE5
sQMKuzWEo41MUCXz5KwrVWdeO9wFjyhttazk45dFED4X6vwcViy69uYfMDQ6Rx1V
vpU/2W2gguXj1a7pWztv+9FZ6ReI+mTri2SzBjEqnW2SVUFg6M4WQB5F0+07G2ag
vqBLPjtJ8DBMfB+RX12kaQ==
`protect END_PROTECTED
