`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mi12azJ2vIvFycJHBsk7nRs67kdvyosoXu1CytalQq9+jtkmiygRYphJ+vZmtFNO
4IV3Qjy3iPJyw8mhXygHs+paH2jz2ARpxb9R/PQN3x8gq/RC6jprroxLwdN7ZWST
WHW83KVw5iMitJb+kTMmsSblmkUahCuojawMt+Ef7s4=
`protect END_PROTECTED
