`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGzD8vvzIMsovOxOl3hqgiQnP6ayKNY9SW6NZxXYeB9i
kpkWkv27D6Ke5/KBHXK2hDgkJByZsl65YwpK//T5q/ZC/2n5lsniL5bz48jKl/8+
tNC5eC4dDg9e8ja1IkQhLAVP6x1IHTPY6CfGZxGNkeoQmPgAQcac4+A8635STNJN
7rOgqLMsE5r5CrG1+nVLTu8mXDeqWgx4dJO1ZhLCYPnNb8hHu9isWKF8T2/vdXBi
`protect END_PROTECTED
