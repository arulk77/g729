`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJiDj4BudJb35poj+1IhaT5+WzcSmdVamlkztWsfbV0y
e+tjKcWB+zIyV2BZENRxSygT9rp2M+mOKT+nGfpneNbLX0kq1c2B1ijnTHMUUDJ5
WJ0mirrSNRs0GLCimiE/xM6bFuWRM1MHQzVM/fdTWjezHde7O4yGPT7GFLMcbjvk
KXbqZzkfhlbxWFGj4XBUKsuS97VH2+l0+mqPAJTEIPeK/abk3jUW9tK5JNfR8zdX
4adTzfUvHIbwtLacmzLp4N8TRQX6OHijsGmjHfSfj8S4oxKKNE8qPIoC+RQKoIRD
/PZgOS0hSXtDXyJigOTDIGUmEWYJ4IKC/GY600n6QRV80f9OK7S6HzMO8ntLuh6B
2PBBbAqvFMmDyEUW1n6OYuu9u2I+8x68socEB/vehIu8Hi0LIvv6lKCIMm21k/5e
+xUsPgS64zHgr7JQYCi8EwpkrcU0NXYhagfnJkDsW/9lmV8HkEazSbypJsfCiu74
WOt95HuAVr6PiwSpU952sLR/rhWn6i2ssec/ak9ItMs=
`protect END_PROTECTED
