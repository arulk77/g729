`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44PY4nKrFyMw+DCnwptYIJ8QdwGEIPtvgI6p8G/gg9mt
ZSHQ8TdTzkoau6udzGK3mn9CeAmLXzwPGB2GD7oLkVpPoq/bzVGMP7+vd9YDU1Up
8OvnE8b6NToL5Aepb4IHkPpv0N1b7EM6TfwBXEYs64ujaJJt3eIOBn1sL7uH8RCV
UEdSggAP8oMYROedbejSV8yWtbKl/EU3yF07Ij5PiGZbFuV8GzyEhB3WwHaztn3W
HVhOqJGHYqUtVcqi9T2EkbYuUASyMs3yzR3Fzcig7r4=
`protect END_PROTECTED
