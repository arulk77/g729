`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEvyTQ/n0JIuj9dUn9Ag6OVOKjRWW0/N/l6Ia8x3+UQ7
4MfQmTDlX3knZmdrHke3/Wo9s+38lmmZs+qTcMdE1VKXlkCK8tGcw61dZ6D6xyZI
0/sD307Bn/qQ+8AmgpXOZKN+U9mt93a7hFTYPG3CnfK1ISw91HtCafYYKJTQ8bJY
oT/s+sTEDXGJ485gzZIdQQ==
`protect END_PROTECTED
