`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40NuLOYfgjCLGZQfQwBDo+DMVwFfcGOuFLRLcHmr4/1a
Q0Z7vWVx6Lhxg/z0x5ltKIWJpvmEhg9pqKDvDv98YDSbonl3vubyP8dGrMJJWZRb
ljs0SVYUG46vBTQ2fRbvKGDUR5N0j7LwyokOz/L5VnKIFkMTjyWlnIZjz67sg8Np
a5gfoqvyma33A2Dbk2OgpXCokwoweuAaQNEqTjpYwkeWea+RG+hV3aQ/fUSJMdgt
pDCukXDkU5wLj3mH3YNUIfBAkmSpOBTnkRJuB34TITc=
`protect END_PROTECTED
