`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
6oIfdjGtrAcoTkCQY8enO+AcZoYQdagMMJshro9YUuE5TIYm781m6BYfhZmOIvkC
5mA2L4VlcThBbOVBdpjC/L0B5zCr/3uXPkGACqc7BYZRjUBc7EqTliAzKkIjTrUw
o6ZYcZW373RcJaGPxdAYVk3Yxeo0LSzH34JGxQx6GzMPyJSp7j6ZxCznOgh8gbBV
cWsKLveq5gfGfwLWwbC+dvLri+QQ4IoQovebp6IIk/UmKQzaGGpgWNSQtiM3Td7K
JIh8HuqiL92FNPk8BRHEQ5LP1UOoZj5yz37EXwxQN28yALICnIu6Wl/uOBDIMNEV
aBsCSJV9lk0KLtsJVUnxNCAbV+EUPz7Bhk1nwfqNffgvSndoaCmWCnZeUNhapghY
tI8O+6zIY9LUCfboJYkSSva9PKqcMqHtfOaPVpIc5mAl0TNRLXI5Ig71lRMLMV4H
FS9e0Js2RU2G/tkZp04bkwjqaq4/yQdQTtN+3DH+bumbCROp7Iq1ClPop4OduNcT
Nry4St+ZMORXll/5Q7WR0WscwBZl1HBwPyYCF9R8ej9EV3Nuj9UWwmy7mRo1npPP
mwhlSr6alOGu5aiZw0cs5xgbAH1c1SQuyu1QTPKk6s8Dv9W385E45d2cnxytlNBG
cBz1C96uLxZyYDO+NdL1V0ajE2I5QwGn6KcCZm2SEaG0fh2kR2yvPbSxLDyOjIE5
6ay2xSg7Bzd/NIJYt4GUuoUD+zIvH6yP0TDOHo8NPUsyUkKqBLSUR9kL5EYnJ1ob
g3ipuWd+4IDUF33LRpq5v3/Y0DKoSho7Xw7YhKNePFdy8SlxCdBnIfu0MWIgYKgx
9f71pWLxyEY/0IMnu10+ZTj/06j3LtyiGc3k6sZno3Sd0MKr3R3UXEPtTt6UDK86
67P8wA8k2k8GrCg9o5ezvHFqy9g2B9RjMQukJCKkUsSZCvILbluI+BxElNA8TjMP
308MiMYKTTuiHBWAJ7gZ2i3XZyQjPudsUsbWjxPwenUMGNIzxXpA6CcRBZxPG5uS
M6B2YiT5RETL+HBFiaJeHbsivqPyPb85YjXNvjy6gunhS/7ef2HrERp2/CD4Di3i
15l/kjCqeDwILa47jmqQWMSs3qWQ803JygW6PizNBcxs2vub9AUvnmVEmNijTAOA
x9EzmTOCUxaJ+pfbuRc3gFZlkUfra4sakJtre+Y9ZWY=
`protect END_PROTECTED
