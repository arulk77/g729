`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
CvBGf/VRNMnz6w/YAELUfp0afDqVviWxIn+4TZdlxqPJ+b56Jo0MVEhnd2HDrPnw
6/UiuOlhAmFZc/GLR2BFK18HThqHzQB4fPegcaj2l3UNuMq3UfS9eUDz7IPWV8C1
NsOdGxVlKNMEs2RD+s7eZMS4TLybDpdZ1e8l/AyALEc=
`protect END_PROTECTED
