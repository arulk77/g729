`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
DqBsUz/qnp5FdJunYOYiVzFRhLBQweScULgjQz8SSRNdrGSjfq6EZcNsic9hjuVG
o7/GpSQhKfphOkxv1HG1TLvnyxwSFMWw0NXozUa5VPJQiT/yJ7qlAUA/zVz2kbs9
NREqH/M57rREFxCkdUkKuN9fOMsu9VHlTJmCyO6Mnq+5o1GNuQ4NpjxIc0hVbyBs
vBR8tgzTuA/QzImUS/f/mG3ZzUsd3g/sBWX28/Ad0X8PfQyF/cYpnhPoaAJ59kn3
nWBbgsgkvE2eF3Bkd3c1PjM3OFBL9SRCneO7rKGXEzM=
`protect END_PROTECTED
