`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
dOzHKtH7yHl8v5JX4DkKAkaQgHkISc973nbv7jAGdX2AWyDTYRojtG2hFSAdstqy
vlgl1FDxPTm1/7+vnm1Szoy+mszOiqHYXzoZTmmAlKRhqhjefukipO4GLK1LaDz5
sT44FkRnkuCclWEjDAWhdUVcSpwphkqNZ6YJmVeJ3ph9YLvP8holRoYPeLQ+uKwA
uXLczhOq8EfwpswA+TtRbSrhQQ8I9bmA22zGiTVs9/U9ylB1vHjF+w5PErLWzt5/
TxPGzZd9q82MN/KJukUVDZjxiwDxNaY+qdf1+RlpgUf60i6A/83s8XbfI4zUz7n7
i/LI57xwQQWaRd/n3gh2dvUIORvbA5YmmVjzIHCJzRkWXuOSOTjAvFMSX+ENRB5C
M7UO/nEvtRZ+VS7BQJOfE15gJRA2oWhkGC+bsCXeW8c=
`protect END_PROTECTED
