`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
o+4BhrxkTh4YgF8QzpEJjAa32TCL5lJjiVzONZd+3mis4+IxTTfU4VH+lIlAMP2r
pvZxKmHq7ZyW1rB/zUYJedxEuHFrr1XAg0rwDfqnc9gLb95CtuOBJ3CWhx6KvDy2
SYlPyhaaZEm+m8v6iOdHiEXRI9A3X/3zMmLDTFKuaR26qBx0WrofbtMCYz1HFfz9
htEGWaRo4Ctar5Z9TbpbP1B8ENqChaFce/qI40cPJfj+ozZpbuT9K8V6oCGS45RV
kweHLhyasmOKcPQFcKBDE2UpA4tzCZAzV5LjFl+VeYfI8HnwVEqlsVITDTFtH8pU
2HBzJlr8A+CJ/5emtvhbDzDshCJRtoLjl1iNrdO1gVA=
`protect END_PROTECTED
