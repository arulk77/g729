`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP3MNBdAx5oel2RkSws0/tTv6vgm7t1rcL6GXIjbCMLr
Tixwrch0vqRo9OtJkypq08OMnC8uqYgPXytxCso8Zp2bbh9ClY4I8JvW35BufjxM
51lq4yRF4K9cFQw+l6jjHbZuA/l8w71IrzFLc/0MCuxFPZ4t9bwrm/MUCmNZqMg3
oW+88taxPnkWcUpKjFWKZQ==
`protect END_PROTECTED
