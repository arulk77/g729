`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePSBkxQIitcmvrYWDQrcr22HvbVLH08V66mcxUtRFZWy
eBNLndNmJC9bCvDZCL6TKtdCKQY6wveO2qcEZcBDsoA6Mm+fhXKqKx1reSSFMNxT
33knOSHXDgXVfC6YLkJW0rYRWDd8ixJ+L+LiDVpxScKDo77X+KUWEU6bSJKuOHcl
1kkeuP3EYTVi847tycuvFOC/HZWN4JlFfkgN4Nqd73WMFHDlQsLoRJMmhINGpRCs
TrwMq7pEWyXXXoD4lP28mgQ8wXKeIeFjrCmK5uoXKhrQoL61g0P+65oXp5y6L5tr
xEjw24WveqJZD+fiDs6Fr0yj3rC7RbK2fCd3cq7o0NeEPo37GIIivk3hcR9dKa4u
5Ty23NiGaYPzNqysuE3tOoezkO/yA9fAXukGBmPUbAg0B+ispyESaOLaVzBpST1Y
svFaEsyNvw1YpV3Za5fZn6SG2qXTe0D9tl5V6ColaqmeCda5MV/bg7HF0CbyjI4m
U0haAgchQEW7E0wMEd77gpG9/iaBQ54iQFh+py91IbGB0U8hJ5ovQsUBPWOeEvL4
`protect END_PROTECTED
