`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SeLJPrkqI39W40lA+maupwA57gECcoHMgeQWM1zvy0By
ikqZdG55gSLfC7U5t4UuFXPRvJx4DxFYw+n58QsAlOiMXeQLKyR3xhg15aLxpLML
5KzKp/+hjF55AduhJON3e7iUWj1DVAQtz0favLrqc6Vn9jr1V1O8uO1as36Vzv/2
e0JhweRdqMR23XhpGCNk6a4AmVyL9N2Mv7s4VAbMdCVou/EsiWzbWschB0gL75cE
EO35J4+qPpX+PzM1DPR2yW4YPPLg+omXRcprHnBFmHCZ/v718tEcNkZXM4evPK72
G5Wj2rI22ChF6ynKm8ZZ/p7kMUa/YJoKs76Ua3a4L72G3NSssg7Yeh5x7sid22pw
HHiCx+2kItIvJlYhNIV44ZrKccDCnX7vfFG6AahxxC+8rMbh0/IJnmcb8lE1Q0w0
9pibwswQDdHVmWAlm5tNH4/MQQx2fGSQvIaD+7vTcWJaxLZIBXa3igM+24LZKg26
EnRhk+RwetyRcfEQQv8aTEm7RSp9d+CdSWhUqE5RZ+2t4LTmOPVpRHBZmiQ+SFTI
nkZwrv1kehl4kmLgs/uGtga31ahjBqXPufV+N8mlGSCTnyCCErW5ZvffjgNTHY+P
y37Z0giruf//NeV+uY9aa9t03KDZwW9ZbP7s1cjrlyhkL7alIuvodojjm8oYVh+B
2O8M/Jjgggnyi4bG4gxEpSlQe8iyZHVqd7kot3eHpQwAwdFj4a1vMcdOUV1fn/EN
sieTWFE+jDYhxN2wsbEK3rL6XsHU8AASyLWhyQ0U5BYaRVi42xcv10rKBrftZPrr
NXsZPuy7pnZZU7jYzZ9M4OvJ/CGLuv3m4V17UK5OWsHSxvXpWUUB7JIjRhv14XAR
AeR6Kw3U6/f4y6uwMRbIhFofrg2rvHXTZznYabTHYCYs7CSuaSdPiOuLT6vOlYU9
K4Gd7HjWiwAYI3Fd3Pp6/i8icSGxdJfgfrm7q3lhyCxXcfG9Jq2BUzqvVeWlkZyG
HRSlC0Vsm9VieGZcRlbwv+8B+KDq2UTefkVQiDJ9VZ974+E7f9TVYbKX7YFKEWG4
R2bHHXSOnsErkDkTp+7nJXxP7jWjpf830oMCxpCKDn1hkPYrBScRu9HscTuAi6/A
dJyZzbfQLvnbZtXcncQ+QghUy1sfc2ifS2n9l22t05pZnMtPqYS2zDxpNKLC0Y//
ilUS+Sc7JjfDuyQ2G4YJR4xkolO0PQjMYfQ9RK4hc/9oGALi7Gc45jYHNDT5N5GD
aadAGEbSZyx4R+T8ftSxIMBmGvKGT0NGZIYsSBZjIZ1f6acGJ51FyFcw/ulXLTHP
bGUHTXRF/JwbdxA8MZyB7D3raDfl1xgNa8BLZ1JHEobDSa3L9hKcua9Kani+lkCj
5SBBWzFLGjQ0qLNKQwfpjvuL2kfu3DJ8QTJCY3ggOMJoZJpRefOu2WTV1prgLxFB
gcEFGdpbNIQvsFyz5jne6tFam9kD/B0XgQcwDlybPwC5gPJdf2mUzlEOBI1+4sfV
nBnqszFoj/DLFz9yzd9AoAdj4IBF0cnDCfaHeJRkQdeFpRl1gaiLT1ZdTsd0ET0X
T+SOxj+OdN/u5Cfzv1voMCTwb94LQiTt2nNFH7+YuJCmdm4gjx+yu8esnej0RgO1
s7y3AAZyXrDnnnjCk+wFj0tATNXWR36SVHRvFqy6WAUmh2e0Xs4znz3Jmx7sTkSp
7/HjMOzxSVBZ8hobw4bKgETPQ8prc5ZCtW2XNpeTqNvBUetCfrN2nISH/er/Wqr4
lUjZ/vUe9BpkqBz+TNnYpkr3YApSlK1xuLG5lGspPIoZPJtxXkEZ34QhaF57e60n
hNl2VKUhoT0g1dxxY5hVFH/fZQnHXTSWkh+3SoGKc4unFA756bLS12nhJNp+8/oT
XbEQTZwwi9qAP6TbXwemIgWrlRibZBrSLBa/zkOuNQD9r1++ChvGKeXIyK1WV1hV
GbD3penoAFmK3becd4e402SNBwzqCWkqysmEAH9sPueH34rmfiJac7JlzKyeOFdm
pCO/O/qO0ih+0brX6N0PhKavWyjTuntjwxB42ceSnC76eDt4Lau5Ym8rok8u5b1o
KgJxXnzUz8CF2TyALiXlysMO98WiMa1rbQ7sZHQS+TOl8bYzO8cXktJ4OFTdxA9N
6CIxp8xvhtjwNAevfdyii069tk3iQDGfRFvj80BD1vIjoewwMSEBGQEvXwNm5T1s
ruyu0x1ye9+iCi/SVknKIe6MN3Ryzj2R3g6RG8+qvNkxAiD09yU0PCBuEOuaSB9r
Rn4+Z4GJfDPDwvq/k3FsHkdu+DurD7QDRnjp2l52MzWWnO1u9Y9rAYFyyoMyGgIv
9Pb7AMU3HlIzQ0SKCSCYZyqYBj8zz9DfcXTr6OO+RXLBOasNriHPRq/d1dDNAeHu
SAAxqWBJx5CbnslSbUk0DygIwAY6HzdLxU9wBU+hCokvIHyoOCL5tGv4rsTBczcN
mJbzU1Exoji0MotZ4I1OIiVDZv892DxIx9DuGt+1ycJzzMSeP7q5Nai9z/dsxhXv
k6ihhOputek+a2Oqk1nZ3ujJZc4PY37mR/iog4YBdCNbCO2ZVEW4v5y6vye2bYmi
t1OLqasdaompBje0mZCjYKbwZ7J8YuTsKBu/w/LPCyO+H+t0h+PWlf5ZcNf7IEjE
2p4LVSQ/zzAseEmkfuLPH/9uQZR07uqmizIbAf67rXWJIuUtmaZHsd4cL4E1Q3Dk
vViBQzxqZ6z0alTVe6/qcp6WrYHOLQLpDryHhamBtr4VuvjYcxkz8uKBTdGcQgjT
1+tJm67xgS0QrEjP1CeKG981EZYmSlrQCklzwVd0XmL0nZUmQ2GfzHTDInjmJvyR
vM1tdoqtRVEFrqpM91qTRIWhmKf9YqjuRST48iZRmO/2ib5hDTCLo+lcWbDg0fC7
DlC37P4BziaEo9MbzL1SBeTG0EhHHNd0NbtHb5TmUAAv1VWT0ao70ISwULDmvofv
ItG5GaoiQqiD648/WnJfbreGTZytBCuLjFZpJLa51w4tH7pozPeny58creqrb9Qp
BeD4AQxWyDNcgNbuQhxoG9IPAInibKN5V1bXJZnM+HZWxHrVZ1ygjRb2glF6p0w0
jGAs34ez1dWblouaSR1SVMcnn9GiP04E2rMOD1VutdywLVHRGcAp2hrbLnY1QW5V
xGg9NI3fFRJAJjKc4nMkWms/dLknYDgLmjyv7zrPlHocMwUvxfi2yziajNMHK3oL
OX0Zm3RKbWDkesgYFe4eareIYLsstZKK5oqj7l9BmlavfA6ZrBq6PMbci6W85rJm
HPiiOWydqPyQzrN8/dDz/bC3ry3mE3nzMn/SbsWC5PaUfIyCIWe0yyr8WN9O2Znd
4Ry358ZT6q5YR94I/i7bWRwifa6rgd8ADvTEMaQvMjjiU24LxByMyjUCJubXpLNK
xr433pVU4MzjY8SIrDKbyLyvT0Puq1ZkGznfRvP3Dn3KJc6S2msoS4ZrvyQZ4bGv
xLHhCigg2WCOVCv2p9g0C2IhhjIKVVejBAZsIGzlbvkISP1+IG2qwUvsrItAeq4n
ZjGKABPQ/h1U45UrsnrdS9vz4+T6t4fZRxy29lmpC5xUcSMTwTY7vWp3asGvs7pY
8ADjzNcV/RojKnDmcU+FzCLysGjU2X7wdQw0aQHtk9ii9KaH+KZ2E7OvuOnGkHoY
kiSBYVQdtv1WrwRHYExPesYHYAqxWA+QLYNXBdR+3XS9J2f7PuaAFtSCy2XeDhTH
Qce3icI2kwdizEsXusgco4MaXoyMaGL1EZ324w3QccPrX63kkUnidTNVOJLrfQkh
DtgKerbuh5XWcSW9BzpsDBMAE1SInw/tGijmdfUpgTadCBujVuGQciaNXIXbcDbW
Kbl+PLtBsqHob5Rq0QYt5IKgx5wuz4SdAeCivoQRgZdNT0lJmohF0W7b7BqjIdEg
QQpnXjvmUmwFpI9OiZG94fnml9ZidTQj0hQZhUrNOol5ZTRyrs8SgkhCDliz7jry
LP15CNBzQUSOuBiplq0F3ATJVnJD7jwYiPUX0kk3HkGtUDI6TKjYha2MeH//LksY
G5pMmlG6pHnFt5FVDUHs4bH2OCNloxQwUvQICw2VzIYcaSrk/DykBWBKaa83p/Mz
qzVKjXiFy6mCm/B3xoTXWATidzfZv26XG0V4/TPJQryrStjxMdphd5vNrahIcT7Q
cM5pa1+2TqVE/o+MGiCaqEnkdlVopxnI3Xyty+dLITP1EtiWSvVzdkPqCCXEJxXG
nFQyMkobMiGmbcdnrg/URrg5Pf3L7iVryDMgJgc+xJCx+BWLpeAO/dtFLQxJW9yN
u15nWDMTAOXsDHA85+Y3JI4SnXMyWq0ojctidaWRCzZ+nvizG61+av/H8rOwmJGx
ucLMRaAvCmlMrDcG97r6TXngqKP+P1HfT/SaQyzLBf2ks1aR7qpbdp8/J+EPJB2G
7ZmszmLKMa6sr0KvNJjxWb7quWfgfY8MJF8YHW0yKq5N8oMD0vDl9L9ICqWHSc9t
8Cfq+3wZb8zrTj/0JY6JI9CYZLsEkycxbm4UMkXK0hd4iwML3k6UCwXmkXW4W4T0
E/nsfLo8rqnwMbKstILHXNj7rAMekGkApuXQruKN10KhcfW+ZccAkWUaj4+2DLHJ
ZhY/tYKSdbs0ltnywcKm8tNhC1WT6S2FCVyke5W4hcZP3bgeoKJXb8h0n0HZvpK+
GZ6mMvEXQVu+xg8OcdbiW94PsxO8k/z605OQO0nx1rWJ8O0uMSXjPsArAdryB24u
DhHR2y+hfjqgZbWLZTYHnlOp6Q8Oe651iAGtWtgDDVW1KteNiScHy/9mesDGKZKZ
y3bjKXne2N/zcsaV9q+zNvmcXlYme5QsWVeLApQsLltr1hNtpPENrPD5fjvgu271
9cxbzC7xgvbo9IcRgqt5HWfUQ8h5JvzTPoeaYftUzJcJL+V5TiR8CHGtmXhA8yWU
TCCpzTxMxamql/zOEP6f7SDTdn/VBCJw9/dSuFf9kcR6+sB88/5yGqoTWF0lJESz
bn2faXI+VvCrbDszBu33zZ61LyKd+JsC4mcFQkTpgOx5nOC5I8pmivqbXdN5hUKQ
cB5QE0hLAZWzTWFxbNblldmYGN4htXmvB9chgUdQkZWH/ozQhDoAoNSzbpSoley+
mW+yB63aq7u7UROP3rWg/6kVtRUEPtb9Td573/wUpfOxG1FZjA8l70cmJqvL8od/
bJ/HX1BR9h/NOdQ8fGIFHs+25FQnf1EowI4T3fdR6t+PmY40Ht9Hrjtr7H1CsP5S
QVfKWekQYq0N/ymv+Dcs5ssxDnfBphrYrxbFd718aUKzl/Ezyg5ajFMY90nzzkmZ
ZuYV1oGpHSXLD+ZAob7ndHxvcndSugTZ8M3yuGuXTWmqmeW+Gq7lwHLR79ssmG20
wAO+t+4sQX8Ut78duQHrh+SSFwWJ139a5seZeVZeATZnVNkZFl62aeZdLDfl2RsU
PIFPzrUOHTh58X7TTeEDzQEOjjcXrffR8feC5HW6yPINjBhMYdFAxE9mEPFRotpF
klqHwZcl3Yv0VTtNB400wR+OA8a8C/s1veJDuHH1oRIkKqNF9E2RPEq/B79Sx+kb
DnVgUPPzapKffaXWp/H5ouJD2r4DTTZzkWYN+mDqHKMcQJC5CyMwfYDcX94DbP5s
qbHut1ElBM8TXLS97SYR/vIQaOZBQlWqzxt/LHStYmeawFA7dJznk+36825hoAa4
/92f+O6TP1YwSx55USb60uCJ2EWgDPluNDANbN1xWujSvrqQXS9q5rxr3g7Xfnyg
Je6q8idu2BwkCp7X8+HXTzFAeBKF2CZE2tgekgf49mx0iQHrcnk5sfcoXePqRpwc
BDKYXQF4wh0B5xJOe4AnMxui09DNjJJ+L6mon0sdcRoO6nEvbjPW7bqzJcX6/ShF
YaRp1GrwtdevCApRdVTQP+ysOjYqWxZFfjTgbJKjb47Dj2MzlQuJl5Z6QNToyHgB
RFKNX/v+eBU4EBMKuFl8TVFoEi1gukAOFg6X7g2hleJ9gnw6BbDTJBfDLcJOmdpv
ttKx1asHFRbZAskLbYhZ6sW4j25IRNWKMThORT/m//vXF9vNOcgVBy276ENaeabV
aCBqpjY3sDVWambS3ZfXKKJCS1xdfZeE5Hf7BS2QG3mUjGogibhXeVmqhngbkb2p
ji6lmDTfQd+e7I9E5TEVveD/w5pBNLWTBEq8+2Kwh5R+gnj4BluxNggrnmbmXnjo
cWAYn23j8wbD0EL/y25SaTwivEItSWNYCs/jWUAfwnTUnY50+kRfaMpYVel8izcj
gvkSsLE1Agj/EOdofmnYDIzVHy+Vl8h0SuLEcJpS33tNYL6CaTFwDPGBRWsSUFL0
5xlSTyCV5yyebQlH87HVHZQ0u+vxYn98tPlviP4Iwp88OVAqkcOxyDTnTgVcjtog
itSRFPPvHifJUDcS701bKKQyTnk782zoUX5cLkKoSTcu9UosV9rTexmLyWzQw/EH
JfDZwxg5qrcNm9JMN4CU+lQeHVR6RUTcYL8W5F4icVH2xqiZ9fAHvSKF+YpPtt+G
ocPQNJK8Uf9hRmtDFJRIbHaSF1BBp6OdANciZHDAx6JNlz5G+4M3emCYFQWjOcoy
A0vFOMnAFKsIpVRnhV9ZrmR3o9J6WDgsH2jXNgSswGjaaHx+tHxtrFjsopzouKDc
P7L9HrnJDzgbGslUoKasHMOPWiumPNI0wWcEAYjmvED1LVwXnMXySnBEmDMnW8id
k16g/BMja5r2Oo7H3AtsSCVrjvDQsyhOJfhxyfXQSzSfJHfQ3V0nkqQqXTuHFWVy
2OEaK98YBSMLdcA2IMU5FU7ztkQbU6wHm5hCxWAtLkWl3Jvb3VVDy6n1IeQ/s84q
8PAKKVNDi8fzG78Ip3ssS7fjKmGwkwsTRog2lxrSpw8+i0Y6ScUHi9ZxDVGmiCV8
qpL0mtrpU1PUhmn9Jwn4mcYwR9XimbHsiV9QLAYNEZvIo1n3ruhnhhfqawTAz3GT
rgs9rW/1AVm9xQYk/m9CD9atXAEIQEnEWf9TQXg2CSAxkrOsd/yaq49G3H8GzZUi
t8eWxEyYWV83uUpqzMsxe0Isq+6HHM1B24YUH0kK4vJYNSe7Xe/WQ/1vKY0ABHgr
mUFrATnQljYycgyqaUQReZntfujQCL/MC1489RElwizLq3rkrBw+Buer95DgVFru
5iV3H6Lk+JoRduZx2H2pqQ9A65CV6Y/itw8NfYU9oKq5Ufq924lqDV0F9SCtadpD
+/UX+abGjx8SpZCpNWZv3tNCVmHfmJIp4tgGlPEweXPShqjyO+UEaaZWzoHMHexC
y9aLY31qRJ03caolO6Z+VmbavGzdzcbu8b6v24pMg53vZBPCxHUNvteGJmh16uA4
PGE95F3b2HeyV6jeFYNpvxmYnqVYYDjW/fTZsRKawLkMR5Ap8/uwTE9zlYtCV3x4
rtV9jysW/1LMg+8X0KMPTsCJTzwldVD2r9Mi65HVMAWnkFxYKIvgU3k6mIx6vUg1
1sPgE+gW08AMtrlEUhVnoBvBOPUpiOurmtcYozVlHOtLpnv/9HHbNNDihBkkSKmu
bvDLdU/DfEbpRoNuaxk65EMk/pIiDrhUSrK6YZ5QosMCPjpypNLf/bKWVTyqG+1h
VRuOGENvYVVqlyMwwe/G90atsUF7mNkjMicjGG5niJpDly+MPu4sGsH1dl8lzmUt
W6c/hGIs78NjJ1+nWV6EhVwN/WqCYWhQiKaVQIAZ1AQH4bg3aTBw2CGGKz355K2t
Gyuuu1vyitnaA0UTUNKEZBpHty0kwvrGSYXnhl2fYVoAWu6HTNxYGFYYj847sesO
G5kGOXuHqSf0/QYXVTZ045VyCmknhTYGnybmOwCp4mfkdBUG4IpwCAXq3bNcQkLd
w3lneqyFijo4MyJsF3chLuWyXNq3GldCR1i9eD4LHdmOjy1V7W8PcbvL1RP3HSEz
kJCM2AYM78FABbDYF92GOK14wfmBMG0cLtJcxOXSADdu+36S95V/+cmIjk3E2Pg3
lQMVJhF4ogihOMtraUdYwsDKbZpRfM/jXbOD1NKii6rp3YnGt6UqVtBWUpv9tZjS
Sy+NKtoW0EN1mjJlQDcNjQ==
`protect END_PROTECTED
