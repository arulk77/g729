`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAHvqucvL0qEy4JH07ZsMo0mgAI9Z7Wl96fWn/vY/KSV
su2HEcvnYZXuNjLib7Jb2tpmueShza48kYCE1562MYP33vxh7FZMNyjaDt17LKm5
OMv8CvHr7xgtKb2GzqdHHwIv2ZH+aDtlbxBFYKkb2Txs/2YgmOJL1aD4SZc4fcOP
PRAMWgns9BOOMVkiDMZFDzFIh3/n8kULXp+kh8/iNSWrzWxsGTg0fEcDRbiXtL6i
e8m0tSR2Qw76Aw6sowFVpef2TwbXRTts55kjVC7GR7LcbNOnVnIeieYLOwLLoexm
z976Moja5PgfZ/XUYN6jYTzRm5ncYqibKrbMpV1TMBHiujNvyuf9kmZPsrjvkC1m
tgHinKLsKKbC2CidFa8U89dHw5IVRzV2Uxs9vgyxfGCQPxoPj9GjjbntDA+lO/cf
ksC52z9CltIJYcqxfCxrTS8QyqO+KvQ05UQ02C+RjdO3NZWOI3ck+Z40K8xgBv5v
J4DG48cTV12g3+oj5pvNeqv8ys0oEwFxa1+TCb2zes/BlSR2zYzHSDi3kyttqZ6N
0kQwwuB1pPQccAHFZxlP+uNNcxMKucTYYkD0GlSiQBrGJxFtsqpcEP/rLdXLJ2df
ZkQkOIR4We26YAyWcRIjnosRTBNmN1xBKxPQBPxEDS8ALHZsT02LhtxcOm5oIYeL
Z5HpDGvIRIVqiU/N4nHn5Nq0K6eRPgHfKDGmVz8x27BSx3WSMFjGCnC1+LIN0Aou
n/gOl9pm2yEWnY2lfUXBVBqBJenstUNQBFmAC7A9E2l8uggSUAeWZreFyT1JXzGy
CSToTg8vxMP0bCK3UiZs2dozs6g5fDNR3ApiSP/IJABTJ+Cu8WaU3Am7IsEzuaFF
xp3hQnz4a+oNa8q3/SNWqMvUW0IHVmQ8UNpBUlUOqcnLZsn02N9rWOIcCJehFSIZ
2wGCH6RNWOQ/OaG6EUUdoBlBsH28I6ZGBFPXE+fvrUZyED9lqKRqMD7gpOnSzDGW
MuzfjcvDWCQDKAjfhfQbTKkJue8AKjjdT/kuruZBLN4j4yOiUDNQt+NHGmjFFr9t
8jCa4okrXgFPpYp+LnvwnAH0MtZOmjrOl21BfQv4rBqcgLhB4Ew2zvSI/oJmrX6z
SISAR3RCbr31N5Mf46C+93F9Y2vjylMo60mJKr1Lv/AqHSks2Ov4FzkQOnrGTmVj
eZjtJ/a04KcTuDsqctpOcmupQb9BQFhlIuiT6g/6+rwxsHG88pxyTieEC5gNhB6n
5im1wLheC0CANDdi+f3LnYQkXkDmfGh931aWD2cTz2QrKvxCZFvNm6CsQ19/GYpE
HQ/3d6vdks3oi5x2v1umtBHBiZ5lGYKVZUuQKEi9jjkCLEu8JPkV1vslubp5Pa1a
fOgX2oVMdqkBgGHyzxkFXrUUTKVaVaDAiRItnmjUYMt9UhFFQI5eK/EOODBG37wI
9MCOL9RMabQ0yrG+r/KRP7mYBmOAMWNz9Qs5cel4e7Ah6mTWrQdgxVYLR4d06hhc
D95gJb5riV5hYlDJXZD380MKgLf8RMF+AQO/L3pEQ0UJUQZHLe7LZyG8nuxAFImX
nLxoI215dPhvuzw0UlajvDCRST6xCnhea1xHyERG2O6WaZSnDqQUfbKV5cqmi9J1
xiAE7cOjFpIGKtv8UJdKT/XSuCgKO9phT3fTGwuMPDRC1VDOj8kGkzV+H+luFyky
Spu1NmoYC4u76+Gg8UjA8izo8GSXQ55FwsGhq8yYAQv4XIuZq32ITafMvysF7ljM
hPyhLWUJlvx24+/Foseq0rgEyohL/46X84N6MAa0MkkDLZTaYMqBzIp6bGZY84He
VDc0qZ/ucka0KLt/D6z0tunwAbXLbwy24Q2w3jKX+gmUrR/Hs/8PjQN/FGF3+ouv
Zj2GiDuhV3Vf6inluuprTAwIRlRVKKrKgSUVvexi9DMkDvfSh30MDxwoJVtGQHcn
5pZ1cC2viJiO5nimjlZnKNE9JQy9Bzk0V+dcmLAKiDN84FQUBN+bIGrWGJ0VIeRB
Kn0l/p3Brjuk1HpPxQ1jCAow02okPhim4/nuZ1dfxhyNBUf/b/ZSQwJGcyYCnWoP
QNrgxlXoZIXBVMctt8g98Yz8J7ts1K/XQVyPCxw7skYsmNC/1XKVTB+UykyjJfhy
Sr8VDTAR135z4NIY/Y/ecBNjVpym+zdUqGFZnJ4iwdhx175sQm9QR3lCpmUHw1fG
YOy/L1bY251g7a/302wdNT13JM/LAy36quDgr5AbDmECZmRlZHErJqUSasOWE6F+
u4QhpwL6YYCZegeV9hXxtc9dWCnu7ciI5SVDx2geqv+2m1zZRq1+Y4p8cd9vAc/P
XFGfmEUZn1HO+T8uAZiYbv3u++LREmCiFQtWM7f0pWAGB1M75UwFIIs10M4skV45
yYq+SsmqOsAQJhxFmPfxbaDgoteoo1V4shePWTfVzoYWATtEWJ3RCK4Q9rMJ2gN2
D9cLIUHTIw0qaPY0gmdBBtopYEM++zl9NFoglhtHlbgO3ZsEp2OzPxqxuUcgW8cc
2v1hZPULJar2OcIO6jxfjJyKqF+LSJ7cqGyZpBPd29d8MckyMy8mwk7KJ2cZ0kiP
s4lkEoddoaYOj1dc4i+yWw+Jy8izDFaHCu7M8y+A+GlqN7WFPNHjOAkLhtQkr8eH
Nha0OZfhGRaX9rgjfLfAecx0LG56m/z/y8EPeuj9Z25GekDtISfCgPbD1Lp+zFCP
+HhCroUhsW4GITUFqkxZU2LQMYiK64qJy0dCTZ/Exe+fRJzgcEroeNBtqFBKM+ER
auFvq9+enfIWq2V7FajwDb1//kPazE4oA//mms1xCk0tS7AVdjiobo+k+13QRdei
/LviGE2yOurzHatZh5ZtoaZTfYadOjxrWQxzJpm1twRZ4UNcc+suFEFDIzP/FnpG
qovxd4bMU7sVwPgbtVkv7qwSACSlA4Nb2Sm+KxGAmxgKSe51MAx+ruRsWoC4h5Tu
pXMbO77R0jj7lA6gVy7llw6RkgUf82jaGNcJZVjV5zlmSmqVTSl9eUbriRr9rscB
TPWdg14vMnUxaw3qzUG1uGOe7P4xOaA+xYHyO8Sf7482fTQNTjr8cyc55eYOk7ao
H5vpqmekCXd9Rz+dHYfDYpq/0LXDBbFg/rYf/ZrPO0ibvGNYq5Nb4e40tfclr0DO
qiekVLXAm/1NAit7b5+s/JPcwNZkixR/eEptjAHRBEn54/fg85I1Ol5SZfUn+wuB
slas+LcraRPxjbfq8qiplIM3nj0JaRyFXG5VSmDpNd6yc5Q69MXjm4pdarzd7HPA
GY2FrmdEFUepwdGaz0SOa1/F7qWIT1pPvxb06BU04Z4zHj3Dt4cyHNEedqt0RK/6
/cpKKvOpHZp7VetpEDv0M2Vu7Xt2URkGKY0Ifd7ksMY9LEjqsAaMIgO+2C19zJij
bvbXqFiESqa0/6HoykmjjiAlBw3FOYE1d0uA4W46KwP3QD4UQO6Sah0zU2a5wx7y
SCMiurEaoioIsx7MZSnPaXXyTBSsfHtYD6JwKe7AlhWRokkHm7uQj9UU0qX9GYhg
RwIRSNVEbfsy3/wVhEIWgGKG6gxVadrtSDLWsMRTE6SeN+NPzfS7IiPEU+dl7fNV
ianeKfgIzoIOdbObXc5wiUCzjbHnlOAoiaypeNdCdfDCXE1ZZv9prns3TKuWmFK0
`protect END_PROTECTED
