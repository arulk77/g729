`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGb/Y+NZf0/1OxFc6Trc1Pd3QSreB0BZIBSMMsdJ1/Va
ySmDOL7UPCyg7NW86cGajht7VHLsT03mf36QVXbu4MYewWdatnGfKBAHZ1u/paCh
5UXOb3pwFsrl5ql3XZ806ip42QhP3Ca2Bp8BSsi0ik0QEpgNPIpP80/ZyAUR1+OU
QvCER8EKv7MBqxbAM3VRgBlSqdO281XR/ocU7UVb0fr8tEMoGto0POPCJOJ5fG4p
5NlIL6PJQF/LGCe9OZZGcxUCnQ+KhmmSOB72Yb1AzdBbRJmiX1vuqZvTPPRmG5Bb
15kCm01kR3BXfWcAJp1A6anbcMAV96OSvzKdbOW2Ped/oiqcdtjblcGip1hwrWR/
chqQyLSgkg1eWyfxzpDZ0CWdn2TlAMFE5lCz1/FUELlwpzUZuz0PxhecNGdq2S0j
/izpsKlDQYqfXL1YdcR7uc1fcyoDIVEsET8nXAOH50rfg1C8ubIbQP1p4nJv7Y+M
SF5Mx5ixVdsTDQ8VYrFgTVLPbTrOcZsgtRg/DdxN3B89rcOWXkbdf1FPifVawQ3d
`protect END_PROTECTED
