`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SVQTUz2seQEHfJl+/1AfbiXU/u9mcEVAlEw0UPU7wZMV
jhzGiI3yMoU+GU/IIlV+N7AVpZRwjbRYLhGIDMv4gYGA0nJguFP/Tesm5vK22BmQ
t0h1i1Qd3N9R+TrBumGRuW/0x6X5gRb34DYLDB3lxMzZh7WcXKYHNawNVzV7pMpv
7RRqwvbVnWzuZ8cejFtxotMVKu30iuTv62EDc0ZmInx3klMbvXD2E8OmqIWl9+PF
VVB1pbP64eimeGU2CJRlDfYYZOZ665QeBFyqnJQ3yUbju3pIKir00u84I01Dfuxe
ynqIisxeo/72zYTNkEp2kCaUKvXjpX8ioTquC5P9AEd/I4dB33WgS8Bpt2UhuO2P
FJvDYQMnxupbnVSmcLcANwt9rBMCzTKD4+rl31HAzDlTIZk2kISJLNS5N9tX6PYW
F+UIrBJL2TJLxb/Ivs1QKiDVkMxdJvg5cf8I9V+coCcD/u+RGIPHFrF2E4xJA7jz
FemZbkkNlj2+ogS9OHTDdyOTJlizuaxgBHa/P5uq6BYAL4HftCnohyZ95vFbcjbw
LmHx5A+eN6YPI6EXcqk4UvUsOgxMg8m6OswKWdXhN8eGcKOZUZNDnBZFZ53ozcHE
VQ1BcJbMxFheySpSnAOwBO0eX+OGiKA2Skzx9OgI6KT7dwfQw7GUb4XPl3girgzB
PizkVJ4N+DEfbVRHkgSWwUge/4JKeyWNz9qoVknoon1kwcAwkjA79GrzuPK+jgz5
kbjdV5qxHtEW2zr2SRnGszXYh8SIyJUSlfabVxT4KvNI1WSoTXchNB1K49PKjjKJ
GKvHVCMMAVbbMWtA8pP08xYYIYvNlRF8/4mcij6HSWkxnt51D3LsElAl75u9NpkE
IHIXOKuFhgu/I6cMzvFkrDlLLZTJaf+JuN+CGGdaMl2k6kr2Uq8XCuMwRwSvj9yk
Ta1xaR3jANjU9IKFMozu6x7TYvtQ4ClzoronofgPy/OnRRViQ7R3Jd7LIY1yliW9
XvC4wHzaX7H7d3ZIYx7go4FWSQJQLB5vGXL3j+D7bg7F1J3RexaRpqQGxnhnCFpU
NMu3gPjHifd4VXdSjnnwzUKzNit4OLh0rrNBpS6juMs8fM9Svzuw3Uhd/EnqoMdG
ZR20BVDAFzhSbdxi/pKUjS3Bg4BeixC6+aEw4G0LzJpkeP1UrYXZIbGJiY7rTBEN
ULkXQshXRYAzxlhIDDpq3usM63MdAmDRt1LKmlEa9JFxhJkGo8Y2NNAyeMCUzwn+
Uvnr1zsiwVFCcHRZrrBIgmIuKnR6Mg3tl77605SLBHRfx3a2vvUI/IHdhF1fu0G5
rqFXhribZUC/8Lhs5Vo8mcoMx4KfqrjL4k0o5EqG/imiaZzYbifalUjC0eUwvU/d
SYT+6Y3jTBUhWIAqSbAA7v8A20GNrK36wOrxi7NF7PqKxil2RPzVjXFlT87uFBXl
rqnR2KfIXLLO2dQRTtkDry280gAhdAp3+7NpGxFiwUd0OKnr+2kVhV6RZNBr6QsX
jBP4YIpAxMTXhrEqR15FnFwqSKXKqAZLAMFnLMkD4pdYr92jGqec3pd2frapQS+w
aCYHfRdrmrXqOdckrsIwKEJSI/uASQI+3XRofZRjtp4sjsylaASP9k92h1Tn/Uwq
ALmSCAz+yNW0GOB/N2rj3o47dSNShbDEAtlj9TBUW/4MJ2Vta5O4CXlHxffRL3J/
zlsdrRUI9DpLva7Vp3QzpJoD4L8ds/mKJYR7WTpht80irquO7xNzQN2tidBM3EH8
s/jSd4nQ+3yK7U4kmpYUwN8Tn6yVMXpb9WdBTnOC3qz3YY8sHPVLHZrMID33cl8h
v3jyEeNPz2dTqrrLoCWeBfU2pVHc6SXWJMyPEpaeLxWyfJZfkSKJjmCtWiLjcvCc
fXUecg8oSbI/5SwWMYhdaZOsjzxGj4Pl+gGBlZMgK/HZh/eYCDTmJFZ1OrC9ul/J
7nqrxSnS27HpgWE1qbueZ6XVk5rbZ6uV1Rxk9X96k6rSPjBuH6B7YMQnS8aLpFcB
7MY/liLF2zYBcp0GJWm3jgdSc2zlriEAPLckbW6EpkEW/J65QOVEckry6VPmp1cr
xZdaFSdVJb2/NUQaunH7AFDlpGzEeZ4jdN0sXOss636sWoryFHZ8+FLUu7NbD5Ag
vARdcE/VP3M4phaanFM5YZgDxr6p9v1QAyv0V2rQKi3D8XKTm+qwuDb6uwzdkwtE
MWVbnHxotC9dk5CWdi9lLusgAWyTfdJ3wflf2d7rW728qHaTv5erX1EGq3d0Y7RP
JxHQ7DpbmJG2bXNPD/u5rcRORGYTAakbecefN0RQCTsTMJeGtjqJj3Yyki96+Vh9
ePwo/MzPUfMppIoIvzIfBn656881fAgYubKFvNe7XqBDPX2z/803mz7YUtIUbmXI
sFNgRSCSoqOvAK2GSen5fZq5fLxHU0YMzeVePe3/ebPpk2eJlawDeks1NoPP/xIZ
4qWXw0vsQVm+Xo7e22ZDrsMEUiWycXQC0jTDyh6lqthTlNfyonRg7pVSGCH0TC/o
v5BskyrRsXnjY/sjRcXaNYri4NGIMtR6nDR07XCHu6FUUAuTJonudM/GHwue+pHY
mGrW0QV/ZpqSoh76hc4r/lJJuqpI6hLktJackwazVSdZzPDHckjxh6ymn/g5Yx2A
A7R2Pxu+cHq+vppE0w2odm1oDK1ChNAN4mJpGL3f7a80mxa89jM68B/JBDndmcaX
aWiMs6KlP0BCqMnxUpm6iWP4PQc1iDAtbkl4snMzfbBLTEtfZNiSvVBjrckAss5k
xW0RZW63Kx/ouNowM2qe1v2ApHGkwQVL0m8VXHeE/UCLHDgFocHTkk1cuTKTfF+P
OiV5MRbqYSUbW2Xl2/COolKMbHBG62RmEYWyY95OGKBXRzdhodZCCRPtXaDQKinc
wkyJWfP57fY+cT/9e4rqHF1036Th1LHvh5wWdvctLRavMsK2X+kBClti7+P2yQjV
ECSdTQpIELeOTl2wn2fx5u36b/Y0DP+F8x7wliK6hBHK8bpLjTKjMv49AVhAp1S2
GQi7Cy0dxpbyBrZfEEhfzijDbzVpEta4iumcH99eeJ7If3sE/B/UzEmq06p9AJFM
Et+NKPHGlJ9RWheJZv/ANETF/UpTpuJ4cIrUsY5c6e9wF8lpSZgF37YKdfy/uhpG
CHNoAuNHIuMEvhcUovRcRk8O+YDrxlS/lA6Xp6g3ZE1oIifpghnHV4xdHIbn6knO
u2FHACPwbLXi0PXHQRybV/ARa8H0rpllMwWOypkjBhkgFuRNrt6Q/Ofjwa4r9k/2
PsQROoQofgkxXGLocqRc8Thg0I/8GoN8RtHjh2wwsoxk9ZeNiRqroUN92G1fJ+vI
dV3CafvA3Ipg/Rzu/r/WCYUugR1zZcyXIgNfJsljsUV/wMCJ0VLJt+qv/28tR/rD
T9xPo0uvyb4bPeuyRf24xgrnRaq35Jj/CSkNvnyQeTuosk+aupTvG26V24kBvHAQ
7UxfYdfDZszM1IAauOKq5A==
`protect END_PROTECTED
