`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aXMZrX1lnzxK33aYc3KUzpXTyTbRiCxKYC5b+VDe4Q60
zaLW4SMs4JpnNHeRjsieO4TloOoUa85qWONRxUpTwH9eVeLA2ItYVmKQXUhmNawB
ygqquKyBWEwko6jT265YtYWCGsFRmcOhjrYbFjRIFc58X31Bit7Yhg7B7ER41wdM
KAyk2rHVEyf1tVfhnyHNA8tUY1rM67hXyr53KJcY7TQoCngBBUr8bXsylWvhPw5s
T6CpRx9Z9voKz8qJjR1dgIHR0gXcEyArleJnbpALpxMkiyQfzWFlWT4U7LzUbbct
xY5g7ICy8EaAbn9LzEqEmo+NsOTLjLnbFlpI6QwDxAX+t1iUuLAAJ8yzLZL7Wj0m
sAYlbfNwl5tgr+v6j4STDJpsPK9HH+efBOggXwDvMYhDu6SNacWDEy+diKL2M8Fl
rIPnBJOzUVVYoBoeqXQTDmvNzz/z400R+I4dOZTU0mUX8NaHlpnimjgs35LcEYrR
mW32pA+snEky1jXMZ1W366S96Q1rBUTNN65T3bfzhF7PVnanrCHvJwViQGMIBNzU
KE98XL+Vy6ESq3DdzGoZpN8VYp+fUDVqtTYJGlh/tI/wTZei2kXMSKmNqZau3iqD
hK1PXDEFL0+tUDD0VDkWQfcU/dOBYfmw0B2oOOPbKuZOq4VqEWRELlkuyjoFSKd2
H1EpAmYS+lPSJyIovrUSs0JFmNdNFiu2qCT+VQvWFwySX47l7dAjKtu9Ug3UQS3K
hI2e50s/nN8McB86MaOAq/HJu+hF2FUdeahuAfri1+5CQqa+G+5z+//k5bYiAqNE
M+by1WERmJovO65hbpclPDMyR5ZoC5kIYI0Sh1Y3LXTKXrDV/AAsnZ6iu/GS/g7+
aKQwsiW5mfcHCYpTw18HSsWaD1pUgpcVszLCMH1MfSnCG5Q1BRvqWNCgc91Um85F
rDlJMt9AsP8gHjyC1ltnJDknug25nRENDSyHx6A3vqeIdw40C+px5aDeKRzRvR1V
vCHsaNGx9UK4p5te+0lWlDkayGR0+kfSv5adOSMGXrfUN5AkFfmnYC4CuDvgrvNE
GAkJ/ihbII24l7bqO+V8XvI0Q2bBFbik3fvIHJ4RoChYGav1bFvP8mkqgPg/xeyH
VQg9BfHIXAwkmQlDNnb43Xi0otzd7/hVk7cAJ0gB/+4jp5sRNpPJnRJoZonqTQ2+
zOf5aUywFMMZj05cQTG5OA==
`protect END_PROTECTED
