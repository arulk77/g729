`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKSUe99B9DUvBOdRyhlBOQ3Uxc4ZbDfw3+y16S9WqUde
vdfNx0WtRfn4ziR2+GrFDhQK3vDmpy95hcQhlBpdW0TWLHfpO8ATA5W+f9X9ov2F
sbn2LiUcDc25mbgBl+gd5+jKuGqEgUQakHBwjU3vCj5qLzPG/uLMMEAvlqqcm0nf
aUseU2K14XcTGU64mbeKwmrO7O6f3Li1cOtlwhQBGOfapwRT7S5p4IX9K+AW/Y1L
ZJfmYzCHNlZQZs+pXNE4e5bunxnjFB51IUV3j4ADOc+aCj2fSc8Z99N0TA2cw9m4
xpJ9hhuwUbxfYviwe0KuAvUMlfiwj9sgHt3ybh4awtYOEg3EHYtjTRgeLdfdyEMn
HlOvmGNjilSBCuTrqTOOzI1ErMm4S7d8S2SvXKEfZabAbJe2QX/ONSXxrRvKlOFf
RaQAHGOczJJBEAQt+rqPdvN+8vJfrfXOsXx0qOYxjEjfapOwsm0fMLAiwO3Y+dLY
6ADBkoo4Q9GyXjQetCnzVrvqoA2cWDZUGijlRwoCWCBlTMb5s/x1Rf9l9/6UGrJ+
XvBs9hDf0/8Qj1VgxJkpQQ==
`protect END_PROTECTED
