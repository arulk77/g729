`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD4x9UGWCF7eM0BqnKcI0stPT9fTxMuthq0JQwIrFqCt
8G+yx39G4ahfXsJXkhTMn+pUx+RmNwaarjIfZ7gH8jXB0IAYrj4nR6LAFJNhmItg
Rnp92OqTJ7M4axm5xZMi8H7lnpA4a7+OLZvSOm9QBR5ldmc236aOLcVAAoUNdXSY
y5tHADO+QJblqq3Wv5eLzqdJqGiPu7lengpylOtvZLIfLGybupCXRNtcTcXE24cJ
+O0TBiLl+9oqMEelvc9Qz1FTpNqtz7jKPW/JNL0Un6vAYYwccTdEiqlfXBbI1PWW
eabLusNh8H+wL2RmJT2RE+71DSFvlJ55HvpOwly1tpX2tMNQx5My8p+KQrXn5aZR
2p4YCfpXUuLme6SpEZVnHPTZNwkVsm7vRsu2jPg9Y5ToNUHPrSBuSGuiVR3moH7H
jaXrM1KPD8wDD/aTuuVtiXGrGyqaL4MXWE1vmLti06y2U3tqTIcVi29vQEKjz9TT
`protect END_PROTECTED
