`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
MJNTEskNbylQfnHSNFSY5S5byHMNURMj84FsvaLsoCUyGiK6fT/i7DgTtKKKCgTw
u0FA8/Yqd8cbUIijnEtNHpk83zWKS7uHcXHowznnbNTWS5lWDkUoVhip+zmKp527
FFVmHqpPADhTxgtz0D5AfwUDq/VJdJwhPYjT4Y4ZmcKG7O2mEEKx9YeuFbgoO2t2
GmogobgqLlyfIQ37qyQj6jTnIwgyNcaIwJ05akvHB1KjMXioBLAWVSaZuNMhUE7v
hTyN22Hjy7CrLeQFf2SDyUJ5KIGGpqw+K4Jyhgrm3h+xhJ5+E0xHAluIA5TgJe34
jbc7+LNxMIsXrFUEA9PAyjdrgumTpoLvamth7tHckBE=
`protect END_PROTECTED
