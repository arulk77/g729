`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4x4uHFJvk0bY4R7aDn+MmP5i/KaEq9nKI8n7S+9jB5Rp
78F/vXkWSyNcMiKa/OfQMAKViklZgUM/vJWoKtVZxneKZiX2YMOXCUEwfBlJrmQW
magiBSzylUKe0/hFxu7e4T35p4mfl8iSFVhd04xetoTGDrjEXa8iEHnKiH3wsdC2
JCyskmGh3YDSl7S7ElAlT6EY7wYzyRUX3nQDnrUhQCOGtoOjk6XqPZJVR0eHkseh
irqBEUfzrNlOTq3Z04RTsAdfdG5j64VzD0x5Xp41gRP6uH6gZ+dm9w+aYabBBZoq
P3o59tP7tLgjE/tvyLzIrVY8/KrYKmaMrVNtMt9fp2mGcCTZJK8o1lQYye/Nj+s5
4LW3QnmD8rMDARcL7sjy/Q==
`protect END_PROTECTED
