`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDi4tmvScuiCGKT9lfk1NWX+5DiUP9yBEfp7f7DGZShZ
3wfmfIuuhtIxRFfDeUBLojdHNGcrxxytDF8hFTV/pHq50UrrCEqdZFkLBjTeP4nn
lALH1ARc2uy6dPgYQKvMi4UJq/P6L7bR7k0pf8gkq0bSr7PSThMGJet58F+fZ89i
20isE950l8ZnOIrjXPAPdXtU2RvPN7PUOTrGvrsDHp5ZrGiN5LV4BQ0lnvZ8d8HL
`protect END_PROTECTED
