`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCPwkYPzo3KOI0mC/Qw05BZ14dLh/dZJzNV0+CV0U66k
R/eo7s4Iv5B9xzUs+29fKnp0YbYLSd+4n+0m2frxFQH0VSu9zMQ7Y6az+I7oadXO
64Szipax1x5hJQ/RCdtWGqIeUZpZhyg5nkq6NYgFPQ8=
`protect END_PROTECTED
