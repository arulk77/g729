`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
J5VmRJdDYhLU/oaRbU4HViIG7u+Q77GzYji47i8aqOrmZmXGHK55xG+cNUTrAqlu
dzlz1sxHnrEKa359l7+zcIgImu377PuKlZg/XF8qsu5ca4sWbKtxnoCyiB5amlLf
/+RTePAwHKE1X243PB83irxEWnfcp/AENTC1aujAzKDdgTa6CYy4nLSsdZA9O3A1
MTXLG5ykGu6tj3PWj4lLAlSs4ZssqyfeVc6RQGr8oBa9lj1Y5bGjWa0Ksd2yzr+I
it3mgwoLvhu9wsAYZIxF0T5tfb82eGKreuzTioKk5y8/NNYz4ep94Lq6uooT9RmM
`protect END_PROTECTED
