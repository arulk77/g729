`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3ON6twM0bRyFDJLDX3TyekmynVzN8y0Pp0v8wIpPvNEX3DXJLgjRpxpsRUh/goMF
G97sXXxI5Fo4nfflQbpg/eF45y9CKOzN2dtrbPZrdRLFEkf9NiTMTZTFiQh2G787
vc76FotoIBP3JVHUjPHREqAErbITNR0FmKZeoXK8VDDb4tjn0sqv7bCnc9OwGVPT
hnklB6BHa4dSYga0qNa47g==
`protect END_PROTECTED
