`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xxUsdyS6ijaH8cUdkqf6tzGfZD2oNzVzo9LeG2HxsCI
0Su0Jj73tcN2T+VE83QdbIJ67Rx20lEZ3m4LYZhTSLuvwMdOReKoKihrpHFOk/gJ
zlq16EdXuSUsq704t78gd2Vem6E8keGWOZBldyNcQ790th8Vl1Wb1G/lS23puUy8
k0nZJX/XRk5nqi5s9YlYIdLxndNYvfJvzeaYMHOhph3YltojbugTun3Y5QGmx4YH
d+KT1Q0wsv165dYCyv0trygGt4L9TEi2L+QVyPVBqyF9T61Y2i0RBTr3YK5Qnv9m
9BuFCfD7SisOA6FFrdNZ9Q==
`protect END_PROTECTED
