`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
YJiM3GJmDrQGQ1uMxQzLVFGvMuP3EQfzS1deXHUMBjlAPcY59djLGhn043hQyntj
iGtjy8qE+PlM0h5NPOZqiyJc2h/nlASF6jLvHXvn0n9xxi+GCa4kj31yZGfq6lem
CPFs6WcIkraU0lw0neVBkKF1Rtg4xu4k+dCnc6Oc/gNh/IVIM5gmI2CX5HqMEgvT
0YbGvLlZ5Q1sVL7Uf/4aiF7ahW3dGqik0IP/lAuDD1k7o68p9aZZh8uzBXCweN0h
ZEGUBBDhZZg0JrDQKhhTusrvt/hIqYX+4moBt/TURx3fZrHGZ8BvNVo3PtM1PvZd
`protect END_PROTECTED
