`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aZe10oKFBNXwezn5j2abHqkuW7SPrNdBrJw9W7EAMsUC
mFTC6pkSYiNHIGBzGVMOqnYLgeIDszLE3Hs7MPDSxBVH8wDyFpAN4RWlhx8caZXS
a52HhPq3isQqOKDbvFmrhG5g5bUdXlEdhlqWUNAtNJIozYpBB+vhU4V0CFWlH82m
yJlZGI1FfY5Fj552/fLtGVACHFF5r/jKMo+s/edQ48HgLX0OxzFbi4CleJarBQjU
TcxycSDueajePKObmjmrd0V8GagdyZadezXOq9DpsQ9sirLLS0bqg2vTIBaveLA/
WQRTOr43EJIxisMrluD4sLauAyYT6L+bAsI7+iHHYju0tpw8ZXlE7BBlZ7tc4ciV
iE4alRI6eI0qladKeWQn0DsKpEhO6imG3gjCujXTS6PPf4vxUOzeozLpBF+kte8G
GEUdWDDX9Lxt1/XFYzeGhyldgyl2Bz36mBkXY6WTp+Z19V8W3Wzlyrk2tM6EKxiC
AhVeoCOQmdOHJCLeAfZPX7MZJK11bRb1Bb9BV4CHG61pD452PFH75xtcmg+MjpgX
fqgvhtglUWnvvyZsqsOELYEKV9bG3sXsL17Wids76b96bNfw8LSZ/5CCVdyU5dM/
NmUdQzL17oeeZtGcyCoiPLDw6FoMlEaV2c4UqEkprnzWYZ9gdj8jvL8JL02jZl4k
J1xh/HVyZY4IqCJnVB4LYbUmWkbsGjK5T7NzYzPQEJDsJtd8wqlCICdz92UFJXEp
ogOZAJFG3lpxUU5plaTAaHTSi5nmCLQFxiqGHCkPVSBtw5ivVDl5VAHUAgubFfBa
aD/R1RQDiGMyRR1zQUVmOTWQZbsGmYJc1hm7lVX+1x+eddTxhVlWyamkuo4GoY+6
bgUcNcR6ro12H9r537vbqJ+zJeMuByQXoD/lPn4geFqafq8/Ii61+xgoKqA34kjx
NZ6XFH9Sy1LqDjwHqgPOTPqEdskusDnHMyjMu/Le1eGWgGZzQd26w6PE4RDVAhEA
P67w1PO/OKdoWgaAFJUND98pD6oZ3DjQ8qDh8EJEnfmRywpb3O21I4cUvbSm840z
UEWlUlhnuSAp8B4yqqQ6UiAxjTknhrB5HkRzd3fKt10uo3GMbTviFY1lWmQqn/Xy
/p9s/V1SrQX4YMpfDp2bf7XTAzYdjsWiDgx3P0VOgiU4lvrjt5YX4aYsPpGD15Ht
o3Uks4GR87vi/5X55b0c5NGS3x6FXxfxEzQyL3U8JIuvSZdyZUVJsrK+GzxWDHHK
I37IGgo9diKcNoABwxoRKOfjNkAiPHsGGu1vWDtSRpalODKDAESj0jZ1Ynssabxi
y6VcPvoYsj80OZxmiWa5QSyh0Bdig76R5z7Kin8fVoJelgsJtF43ZgVIydus2KSj
etlharY3AsnGGZYLi8VJLA3uFvcPMuUx6Z1ZoTVTfl8KKGDHDZQodI4u0MWWGwtN
/q/ImJYsrY4paw1a/TMOMRrkSIf8rPY/ZoQ1PQtbWLUucuJgqKFlmF2qb1zSIgNt
NoAi899sA/98RsqVAgZ4+MuK8XHB0vNqcGrntSZZyNgPX5yxkpmn3Kl/P8DUORKT
WDEtlLK6VsTfaqLgUMQXLS/SrGggqX9AkJsq0gn+WIM6lqN/bxZ8WfO6kZZIljhK
pdtH3xjxLo9h8m8GabKCY1xXcgjBvnTIBdP+Sq8uWxGqlHpYDras74iloIA4o7YO
z6HvDygP4ooaVvYYWiL5zBqrBGKH9I2v3jJiBxBmsh0I5IGrQiDt3qbRONDPRg4b
n8w7NwgjBaFjzjTrCFzrAmkLDr4Ph+d6BPo9orG7wUXmAUwFktzwj7bCK6Nco9ga
q2Fc9gulVgV5V5K2zvvETr2OUPWaauEY4i2ImFpQjDtOWraGIkB7xfVrFTxFCL2O
KBUJn4CuG3BDjwFjUqiKagflVokWb8YxlEDa5SXpaRUf0OYrIGTVPUe3P2ryw6mW
b/cUDqB0ao3XC+NMKss/qMisbj/hNp+xCSbAYof8/Sg0sXpye8Rp0YF9wnEougR1
NQVsKGPz87ZIT0i1iqxFpo8AUvpTSlTFiPnyBDbRdtoAD5XGHLgjS06HuTV8DUDE
eeqTcADOCN/SKMNOq4jiJwUBTiBkgNu2bRrnKtzk5b1As0Wi2AdVFLI+7sHHN/uG
GA/8DayfFZIWiY0iqfBIce0oZBpmTaXCtD0OdiE72JyAcsHPIiXlu3LF5OZoXxrN
7ifXGFB+53I/8uqlufWW3ln0mkTUgYwDi/orz1pa+ho6yNDMHDMBTrI6W1BrO3DA
QP+SF5/PGNsmUnZY4apJn//xl2dIEkjQLFOId+mrI15i1RxrOX1wFD+4Na0uNx6O
vYsTCq6E/aYfOPxPq5NE5MqLupYA1sh57OwebWksSeGitNRjLvTqOBH6y/Al3qf7
4sylGQPB/Ee+E2uaexdMqRIxzfGZqnYKD+5Lqdz4LHiyWMZVwLA70buRjabbjuky
FT+TpVfv6JbT4AZb6HyPQhd3KkikL1OgrJHhrwwD7vOe8qV0Hqr1Ps7gA6AXHna+
Gy6E0qQ8weAhA6BvJwpzDlNIHJqQZl2hQJp7snw3qxL5qFsVH4o1vlD/zKH27N0l
SB/ahZOohH1Ay6wRuFp5G/2fugi42hb/aFwJsjRL4ubZqjsSUqvP5q68psz0yjp7
X+unhUm1K+jrlTFjRSKSvOoBsJud2+0ygnAx/3iq2gY6Poz9D8yA5cdCnx5wkQS0
oIOrBcv1OLyU0tDZ8ZLb+t35D64GgroPEf6PIY2qz6f4efgm4gmxpgq/MQnqjUX7
YCmyYo/W2g/OHDQxFZYHEUils1vhjLHYrV0WIctKcWnRRkZihogu+os6wITaSJ1g
aAEDaaNjI248A4gscdEOiMrDYm89/ZCAoDTdLAgmoqNzt6D9w486dR4XWcaoS4gL
fiDH3RzzyTkPsE2rCEHpQQ4H5JaN46CDRasc2CmMt3iVLsymzNY60GLy2vjhwvIp
2c7VCwtyvQR3aTbiSwOaQ7ulelVk7k53KQ0LqM3+FqtqjyhRhICszbWk23uvX4SI
4pAL1Cw3psqSMHrLN3nlMw0Gvlcgq2Xs18SLQvlNiy6YOnSKOdy6t6EbuA5cwxn3
4MMRmg8DyBKALPFCIbdrmG2UAU11KxxwO86Ge41XyjllsW3E6bok3sO06eHNgiFU
s+ngKFuvxKjvLQd2bSgIoJ7O2lRzjSEeyuxdv7al8qvl+W+7b5yufleTUjG45Eh2
Hp4xj4WBvSuNX0feWaulazBU4wF+izt1tzRwjCs0ojtRrJGqFTBPPKXm1JRStqn6
i+uFYAvKb45YCXE0tNXO6fWM6XyxS/Fo0rrUHAhb2wv+TqcWu2UIJlZjqxPBK1z9
w7eBaNJY+6ZqmNF3xG6Xb8Q5Foc+3nxwAjlFtHDzRJokRJnm8sU3AKx9qFRcbJlf
6WzIsQPkXtx12adMjBbkmmegDEUT3AuD8UK87znbCwYxwOdPRSipKn3BIQvuuqwm
MGrwTOh8fSKnkVp6uHJKM0kLoKfLbgeSGQ8x+LLDnWFi9pN/HGU7m4dwb1prbUnc
sMysFSl5yP005nwGlMnYdRgokit3CAKmU3cCSGH3omLw3gteGYZxCb0g+YLGx8CE
ed6U2aZG4pp7SBeudvMWkq5pm56loLZ1K9W1kkN0RhgNIvjSDJy2MaoeI9Y+hZch
SCweAjIqa+DOh/tckAvI036rp43qenhQf7Q0oYB+/QZ4TBvrf9tp0xNm2Fn2JLMd
qJYHL5Vsb8l/cyr9IsXAqaWzPqYV6HBnigmw9btUNQxFdwtY/NES2XfRI34Vh2U+
UPp8A+Gj55KogReQl5z9KImx/5jVASYvTNaCm/KqLYUZKoPja3CvRCvHRTbjRwS6
67wcdmJLF9RqWryDbVEvt7nflXXtrnPWX0xReCwgeTlFGI71temPSWPw1iSDpB3P
3ikyJPi6Vj8oCZ8LP8e8878FZk3SUi8bL1bRDqDAdnr2Albjf+cywPUMSCdzRq6j
LSupzCKGy1NmAOKB46WPdbUAGNnzg8BTdSN98OHislSPPPxyBWYgoEfkQb+AQj0I
FseIxr08RFY6nYMFADmndEDQIwY308ZAb4oh0GajI4mmX4gx+rf61S4md9vqi+tb
jAz+z7EIvKeKRB24Dk2fexJ7QArHFZ133XOtI6/rtbvLLspWbjyVi0WlNZDZMWsM
vEDlxT657kWsoVj/3rHgSWMvUX0CwfVd10FWqxRrnQNcp0bNFdvx0aNKFERVSNsY
PEDFGSgei7SXmzbD7OIYGCux1D7Olnw5t3nm1/80Vn60x0AZDAzdudcN+PU6BSDB
Xf7KTzfahiH4ZVAVSuwCicCp6aONdmoAmOW4TRQfQnUjdTLt3rJdM0uHzzAMnYYA
FjT4vNMaxYgUPWth6iGzNVJuX4BR2qb2MoVB0mb5+1pPy1hGuqBTR32Pn0JHRBjE
fhzfNj0QsE4QuiLOEubcKujWQuS3XeSIlxQ0YBitelkH24nYX5mmmjh22THYq79u
gUmAAN4h4YAsMK7VsdXSK+ZJDrDWYK1ook34WmAbYiNDSTx+zb8tYgWzeJZt67+V
KkD1oHENIQcSnjgVF1v2Q3EftMFYM6+s12O4hneBYxi/Zw6Xkt+GDH1srI1f6Lqs
2EUoed2m/rlCZB3p6db6dxxXKiQ+4YYxuaFL4iJhVN/MSvSbhgLbkwGFH1hzOl2y
XDDSJv7LVcb7Vf2rz/W4qneJwgxCUSaaaDLWgUUNERVOI9Eu+uv7wGMV+sOge9Ij
GOZQGd5BPp5yK/tux1oJWDNrnBoz4Weg034bErp7m8xZ0QBZZfgV02jwobiytLCM
I62IXpS0Ps8n3/iy5Ovp8OF6Tya34ey4Ff3NgDNEQFZ6F4m44eq4sLx/a1FvjVL3
tGd+VIyckcjHh8qyvQwWYUiMETxgNviyWHmyz+VwDUqtDZZOz5ICacfjmw10okZU
0jeAlWp+oduAXGChJfrmlntieDBh/a91u4T1Wrioy71sE/j2Scm8uOV1NC/4nJEf
F8hmBAMam9kJ4cK8zdUW6pXUVinmv3aZNVi1fFoB7IuPj9rfNYwOuYO7cs5VgIqL
lobZ+OEccItNd6hQW2CjYkuTbcMH4rilrZRF9AepaiQYfgTKstnMOB/4kA7+fHn8
xtzqqyT6Bbkrp26Iv6ejwh4DuAwwIJTGPfnoO8cHHq/JFZy9gYqE/uDphXcCSx4I
q7LzTYomdY96wJDU7A2G1hs/yqksvtLw5YrChaglEos1F/wV3xPxlGRhZut/R1Tr
WTHreEzP96Hqfm/AsonSW54zm3cshE5oeDYnXqzmqU9Q05eX+W1zvxskDklBDsXM
WkGxVRXOEYGjwPXp4RM+DDGQdWtajyxcPSoo2X5lw9+gJVWjdGRuh11+4ysaNG2K
1BnYhWuPC8ToC+AVccl2Faz4uEjxb+UOlZO1gcxqnSc+BK8736Jqgod7txxdYxC8
u9gQPXa6lckK2Az6hx8vI3ks4OoLjdoevB6KjEegMqarXn6LsSoG2mk15lSXtQDK
yqQ6JZ5ARy8EZnZ0qYkbChgx1c+xFoPebFXzWBN6AD26a/Jr7B5mBH5KtitDYnfU
1k+IDO3lvck9ppaCe4QlW+bghJrG8ZRgIgIMQblmksseTwBBAe9DCz+U2YrEKfru
x6+/TG4a1ANNkYEw7iU2JjNuX5ZxlY/kQLF99E7mGkHMH7dAeVq6o0krMFyq/i4M
ALhewf2e7ggI7jz4rTd+51l4Rr1CUKakeKzaA75Q1HFh3RZE5n/kuz7vt1AdImlf
In/w9CgdOaOJRhQyRmsIQjPW1BP+eZ6V52ztxqICO4z3kLRXOIkFt/ybKgwtUaFA
8TdhqH/4XNxof8DlElm2zmHFWN2SH2Rc9oaFZch+cQ9enYCvu8EiNMB6sQGgszqV
fJ5UlxIQZy/FRr+vbqsj+97dTPB733AgOCIR2NvpEFp7+T8I+FO3LFciF5PNBEZm
/2CWR8y1bjTQM9pgOb/3YDN+ztGQqryQjDXrFBGJk08=
`protect END_PROTECTED
