`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
AILFoMUiDgZshy0SffwaVwXMf5+GdvIcBRfS/9HfrrEceHR8sCCDwm0I/Gf0nAAC
p9GNQEGPBFmJjCWklfN22XJM0yAYXYZ3aHl7+5kM+CJvzGDXpor8B3gUb9NKQY6o
n/QSbXwc9qsiUsjdTfr20dQjr/5xm54xPzcPnioGVLzLBkqOxORIvakzYpWl5hDq
zE25BzI6nhbmi0rJBaerdws8rO3Kt//hY9D6V0PaMyW/MboU8gzW5jckQRF1Kt5g
C3rBSs1CeHslThGGws1RVm5dCIa7NSmW/k/8GuU7YyY=
`protect END_PROTECTED
