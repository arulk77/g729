`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL81GBO8I0QlF7JZdy+JfZsOxoCdF2y2uwLV68eVDoyBdH
qMAf4qO9gvb+vB5IEH/PZDhgm4x/ngAKu3eYdwGNW5kihi31LqPL22zMJSDKh7yI
luS/xIQCvF+zz3mVS8MCatoUaL+dz/ZP4pEUIXKzoaLH2JkikxboLtknB9I/HA3B
vgpcMdczx841atrtW1ic7FpWpCRm+EXAgZf9aaaRsr9BY+W9QYvL5swvgtRTi4b/
50gWR40LPVIpZodVNe1gX7TJjKU3gZZ1gt9rK3C03+UakduduiGWTiQOjmAuqJgW
mEl3CWb8xaQ9HrT9YuTcZNIdZca5otkGiSb2Gml+QGztxhXZbP78as04IsaYc1IL
dXb1rB0rNqgl0HgSe5mnGBohggFM3CMEPCJ/PWT4NvHtrku8OjPqQ9blJtn5Tt5w
hcxRTTxG6Yf50qjVhn6IuRzxNmL4zO+dZPRYQ6VuXLIfZ0/pFIiVqjkEXPqd2nYM
UitK5FzjgcFqDWk2G9ubbyb0abbSEE3RWlVtpgTciYbKd/3zeSb0rCK/NGUvcyc9
PNMYm/iRN7sIgg++aOXVhkQQoK4dGIEKssOKLX57SdLvNkNdk7dw7vZLPXy2jLOK
D/bxGxn2ZqlJLTghYUgk4yBNtVyVKB2tZW54cK1JFCCLJclp9doRIC25Kwpsl3dp
WEzECLLuRUKs25PflziBZDVeZQWOip3ndEOplOV2G1Iv3/fNfbnWket+S7ObR4AM
vzsvJl3GRmckgw/1q8hdlBa30hlGOHsH6DtEB5mGGj8gCyJfNS6WBd0fI+r273I8
1hl0VaUItfx4wphjATRVjlXV23NW7+41jV2o3kgOFPBRupm3HBkJY+JIQQRwAzlJ
DJKwQMIp3uEuBwa/bO+iqXF6ndFL4Kl8NfFCERiUdR6+ViqZtdImiqWdQGJvAZ37
bgAEYGCVLLrikogJEn1Y1bakyp9KIF5zeEFIvfi4SGB88TnerB73MfR3webXfaDz
QxcTH8txZhhUL3wK8/1td7NijKevqz94Ph3WuYLJ4mfiLREMDQsJTNvGy9sWytvh
NSKSoaObsqkAXlcR33uztzfpjhOpMALIGm2l8bXtXvPeOd020uxyVBStIsA2ab5x
wwSctNVtXtzb9PSzGYAcQSHDq+wHS1rb98yQQajUMOmsiz/xbbHCeMUwUi8QQu5J
Kp/zrt8Ydhewr8qjHz7ZasQRz0maJXq2D8y7WVehJg2zHcmhaokQa/Jv6SCw5A+e
PpGw7wAgNqgwxoi88EgBwCBvR68EIzpdbziMYEPGgdci9kZ7Act4NBF9GYQV+lez
y1KdB2J+8cs7zsYw8YjVgIAjHXGS1nQO9MF8YsrLbRBcUg2bmp4X7IqUaZaWGY9/
x/CToVdb1yRZ2s3Ytk+IIYrpBjjWJuIjVkSzs3OP1y6r4F5Yk4aCX87DEvImggJG
/J2jCzZIRd76ugZD1mLqYosv33IEAkWhjrs2PuyW2SpWs0LT1sJiz/9++Q3nnlPW
tgxZ7l+RrDA6CUNtt3yp4qRCCNUYgt7nknHIQztpYByFWD+JT22u2p+N5FCLT9Y+
GwFmYMef4HRsx/+NY5VzNsoX1NacVYfgOavFfKhWeNQ+ra+CMkd9bp7ByAZT4n33
R8J9CAR2dTkr7LBqD5Rawm7FuRkmjA7C8aMjGqoOc2XbaEJM3cy6kVjLHPQRa1ed
HrswZLEwY/CnD6Ga3tg0uUoxNSy9d6u3jvzWV2ZhXhffrViPq+Vvv9Yjf9GBde7j
JYpEGinqB383j7E4Rt4JKiz6crez64WrHtrpD7SNgUAaKyDbV0snM7jUV9YNaArB
A3oSfj6xNLpM3OSk8GjKIw90VJQu3xqETni2HRh/UZAMSglW+zbYMNLOpmbnzDvI
/DV7sarUDOUhDWQsSIazKv2+0nqL5oh92dtnvqO9ZoM=
`protect END_PROTECTED
