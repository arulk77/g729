`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHRE+cPvPH6JASqS6VKuAL8IhKJe4JGVHOBv1FFtGgLg
bYhkyrzQy3H7g1a5SCZIdLvh45cc2qXPYR022uufJuwQchc2dDeOinQ8Y9TAd/rl
cY4EcwxNx/TijQL649/5cTAXjuGN51nX1Tv8s3vY3MunDiOKXxqinimB2I7RbMEe
dZFon77j5AxmFfIurgcBS7y6v6bE2p5aI61udcNB9jOsRn/Kq2P3FzAOM/2tS3EN
794JxtFZaKeDwzvh4FLM+4NcAAo+pkqQQ2nXn31EnmulW5fOysgc5CIR/eIxzl7a
5e23y4M4UMeb7jzlOiHJSfE8Ada+liLKhLbVwDYiofVBApCVj8qRrnXO03QlswZX
aYjuNb9S8H0rGpY1n4Ccwjv4N7sUoLZN/dm4v8th/oTqDlJtXCoI7thzC+SRmJL1
9hiHgaLVcHdGHy/dOHaZVURqFwBy6f7zrJMooDWi/E9nJN5tLLJ4OtfcghlLfzVa
DQ5w9Hgvn/VnGyg6ryfHHwLiVLcpbxv26HqgGb9w6CQq0xZYhfgyM68k6PAuz69W
/Oz7g4a91Go1n8sMNiGGn2FRnloqmQc+gKjVsQHeaYGKE75hus5mVJxzaPOryImT
PRyL09NKGtlkQpKLRlNceYOKEZClfC5ScT0NDWhZJgjntC23xdWM8PSK8KFVVDnL
+nNBo2TUU+o9qPKXEwmSq8QnInTqXVno9z3RfNIcgck=
`protect END_PROTECTED
