`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL8w6aWZGuFf899LgAPYdODeCxy58Dx6MA3wGBYbyMOGs5
/1qpLZU7tl66Hwahkjmk0V2/vLzBeg68kQG88DfI6d51g0XiV5cncaimj7M45ep4
o5pxftmycQo4KjZpN3TXe4RKIVc4Mbxqb/tYhOsrUJWo0gPh+uRXTvIAFiPICRFH
vXCltr4oega0u2r7z7wFiymanhYcbWMMTxGSJCCANYwiWck20QuVfDFw6Mxm51bA
35KcJJIBFC45VRuenEtmW3AsuZUEKAF1ne1pZZHOX++HxJfsvcv24gT6YNtiwbBG
ol7H0Jp5Ag4VL9QLvOm9PFIpMY4FMmm3Kni9/91M8vPTR7JNUQcGkpFPu+uJThTf
WFsTPolQxSGUK+GWeUhnDqpMvcpmTxu2kDBCZz9Fh4u3clfEW0QMdrmTylUnmRry
`protect END_PROTECTED
