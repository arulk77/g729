`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu441Z3gDY+EPG6Sve8N1IPgyGm6wa+luZqciGDfhq771F
10DI9Cv/lymTxNt3NkJhe4EqmYW9D9JBqxaxs4b/khyFrtQbLfNqRd00nOcpBiFk
jaUNuupi0q35PB9xXXA0F3v+Qe7Q6C1ph7LXoXcUO5g9sK1Wgaygds7Zouyq3dnY
1VD0PIseqPs5FxD2jL6AQw==
`protect END_PROTECTED
