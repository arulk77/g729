`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveO9sgUqSX6Emke2Ox9+hkt3suvNUewOn29xgOkMb0Xat
GFrnCr15H4GA8BzaNFk3NPHZiZFngtXMRFvN42AtrOtTkCxHSosq4UiyzPOcRdIv
VZy7+76/LtEp3TK+iq71HBGvPh7UjcX5STz2ABDOjxev5GsC4zvHSt3Yiwxit73m
ezRd1YXGf+m6OLosWlzlCCwl7eEt9wHoG1VJsmeUY/TzCk60imb/AMugo3MCr1AD
RIy+jFOuf+qeNPIr9RJuylR3/PjVksobhi1lW+/X75INjO3w6ashnuQ+Ogrh/Cyp
JH/EfckOPsshQePpq0Z270lk09ctgD4LrZycr0B0Nj9R9rYJkP1DFGaDK5YTnGGv
3ZaVi6HyuPBT6LlSIC/BEb0bFLcyNqcRJpkGrQGBofxEUtHxmnWdoD2MP63U8ZQJ
2PSwhTKwmAOb2QJ2qLZctbf0Na5SLfwyfk8LTUJ1/6NSvN/3hhWjKIm1GKRzlRrA
B9mXZyb8HG+arpKuteBU33UT0Krupq/Vo+Dt+9CdxuNl/xQAocTZhob6gB1qFaO0
5P9u8XTMwXjidHno8I+d6AuHVwDDEB9CVoxh3q0G8+novgskplWXsWRWjZfHmVBK
c1wk5h8LkUm7bFzaNrUb3AIhYeA2xtPvz+vzJiVcJT5z/VdmyEzPSht/FXq6xqb0
`protect END_PROTECTED
