`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu458tgfWpNXTAvA4J7KjT/j7aEVD7Qac8u03T4kbsZ3CV
pUszpvCEMixKDOev1SZG9lwiA7tO+5okzfUKwcE0dR7soFacA4ARWIB5s26BlheA
QJNjLlsm1nyjOK+pDJqlt2PLWtGqms7UYSre4dBZfiJjmyNqWOEGQtnh0LWm55gI
eCm6Kvx5+Eowg1XsJMY1bjFy2WLeQVN5zfxSc3pvhhTL/2Fi4DpAejubH6KTYsQK
HIk903Q9zOd6muo5p5WfdN8FBO0EZ9S8+ctxxKmiflwVwkfaW80qftLIMF3byUPS
sAfqjVCDRLs/arjEUPtHxKTFw3xR6LMep9lmT9NkNIP/HhapAjPFqGZWXY4cHWQQ
3g/laIDa4hyRIYZlwbDoY34SF5qH0OzaDmGScrgu5UCxLd+k4H0ESZ3CEngvt+b1
CN01/4OG6HKzolwrQLiqiwMppzCBvj2r/m8KfV7MHg6GC8e8pM/AYmpPAwuDrrEE
asRmoclfCamS+J+uD7nZOM2um22k5Q0+a9hSyPehCYYNhMw3tLNbYKo5Ssy2u0vG
oLVZHf+cCRNBqb4jeugYedNWziiBZnzzKFI2qYkrgPY/9ASgvD+YGaHCjEv3T0ty
fGmgNil5IyZQS4dc90swh6FawQFJ4j5TtmjtUOBrbTs4B5GLK9QzRV17M7jGGlRv
qAgKk57u7wOaT2zIO7RMOQq5dUOX2l2kQqw9g5RDCgqte6mfjidi3odCbm5GzU13
KBZb6goptliOLq3vGNzOEY59Z7VWZduxOrf4tZRNcgUcWdPoiaOKunpevWZdHdot
Jtt8/glGhmDduR5/JC5IrQ6FkR2DtkbI6Hn0eyLNBaDINWsmcthpqSkGZhLkU5+P
N6IBwZbfp4u+C1RGuKxPgU8yuKmzr1hc7Q+jcgj2G9wAu87sGHgmD2/z2+S9Dmwp
oPUkuibKpM0+BtLqYdExB4zsdG8DQsKwOPSkkJmGegOawUdV1JDqMJ/tFwU+Qrnu
VBZuBKGJ861hsbnd5PLGdZBS4zyYGyUUI/woLIyNZq/Ixwraor02C/Ndvq9TEJez
GTkAfgo8bwYzKLg6PInoHffQthj2y+Nw4gF48zhiT8MZ7k9+1NaKYIdBNf0OHQ53
nPGVR2WHIsEnn8Xkq3zVIeWgwjTqCdrhQ/VQbXvasSWtTN2dIEsoFaYrjT/xmpEE
vQDxEQE/4L6SLlHURxcPCChKLiC4nX5JnoUfB4YVKeHZB21syqQ7HlP0W3yuWW/g
IyjSz8qY7B4dhJAddHHArugUBf2HcG5ILqYRbJmlNFtXhX4Y0LcQdOI1aibEnASu
ilUKpqFP0CfNChVDp45aIWNJ+3kT9B5OTTXlxN9GhoV8bMZ/q+kZJAkHe1G7WQ7/
s0+B6tz/f7F4NdusLdr5/TT6lCJwlRxN6HxQBn8JiZVE/LjW93YbpkEPqdavrUyK
peSKeANxzoC8w6p9P4jmSr1h3O1anOyoNV0qQyIoRCzn4MiEEz44y0qBiFvJfrKN
o/Aegvwww9y7C/rETY+FC0Kui2qZ6/wFfC0bcDHFNWJ5mI8CYYxyh4TH2oUpmWvO
JAhU7tCRbq/Hqm/IFoGD4qpzOBWpF2O+mc44QIjCosA+w3aH16nGzorK8U50bVpC
OoYzlK9A1c26tNU24lnGU8QaJkSG0efjfxD3hba5lzLwMVsdtIcGGpbjGKoPYp/N
6XTA28lddZYuyLvWINJGUNSsbqRx3OED9+0GDd3WUENU67UDC9rp/+MjAnyPhLFq
V7MUwiNTl5zzZHZVpA9R6OEDNyoDfOOxtWwZOr5m9R4tcRB50WySIA3X9ZCMbuBH
oD70YmbDl/7nOX1bX8h9tguU/GrG1z3MFg1S9v3egMNJ9bA+fv2XcSNy0oRbzGoG
UYSnmRc0nvw4L8zntGImE6g5ccUVL/IBmzP/DBXv/crpB8Atct+ww3O5mWuYSee8
N6hdW6m9jCH/ZKln+K7DAh/gD45XeBhaiv8g3bBdnJO8P0U/JD1k75i2kjlNDO0N
MhWTP11Z76xmaTxozkrAp73uYp14ADdS45e4Ush0HMe51F0sVGVDaevCrmepx+mF
HBiWyFCq4hV6QwV8eMb2S55jdy7K2L5T7KluYbl3IIEtVOxLaT6MXVzyybULmZIv
4uDpboVDUUyawkhPuQDnhyikvlaFrXWcNmZt8Z4Lc7lcPle8w/jPcbsYV98D3pZ5
M75YX175yXncpxJGLoiEOILWqMbdM5M9r2ViTnUzvJ3Hlor2GYfLsJPdrZY/c4e9
5eYVR5GfL2ZnSokWNTHsLP+Pw6OB21PcY9PwTkXJKa0Vnd3Srk7XKhiCl1/zf8Qv
doe8SQUPbmm88syUhVgT0+R4uTXf6AINJCZBHCq/n4vW1SIAfhX3SuqiUAXw6Kss
sdsNy6mEc69cPJMLdfm7j/Xq4JuyCx3lWIbkhsaAee3hViyVmaZ8g/+8bxxhJIPC
4Whh0rPkQImbEzIGoi5MEQ5AxQ5qQKRo1XkHh+nkjKiwTSq6G4vF3ZbaFPmrU4XR
j7kKDauRVFSz3nCClsUJSdnv8sJh8AdmQxWvqJzU4VE=
`protect END_PROTECTED
