`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
MCRrl0S30CrTZdmk/JXB2kzrHM55LxO786iG5IP9R9D4LOTtgQ4U1lojLOLlPlkc
Sp9Ct7KSfdQB6Oqr5u1zXbcrswGdt4v5+0+AxpoFKfI0wb7SODrtWgjMgZ1NELfJ
2dSRk7Qg+aYAE3dTI+v6+NnraGuTqgdvu6/gV9sInxcnPTFCDt6xTY8Kc7lusaRb
GBknvxinfoMTKNItozzOWxPyauyTw1YMeqUggCBhTh+W9uUjNAot7Km3aoTDFVRc
OksSPwtPXb5gAhPAG9uJNeNC/jw/WR2sKYSaCFeaXWQ=
`protect END_PROTECTED
