`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42XXGO+hii/shHKWApj9GpbF+5+cjtP8N9qI1UEf1AMe
EdoXN0yRc6M1SJmO3Nj9+MrG0La0P9PeNyi5JeBy/Oi62HsQZaO38W1aszXNaU4k
TIitSP+o0L93XsnfYhc70f+xC0CJBpnrrufTsjiLTZA=
`protect END_PROTECTED
