`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SWamU7ZKLlGhSvyz8VUtJGWJ9dxNspo4BApk7O6yNH4t
taonmwKMtZHoigd5Ll9g52KklWiW1PdYCA9LeCEoi/1I+hcqeTxOsM7l1ZJ1lUcB
LCpNZ6p30oMMPyjzTafVIMWrS3IlLMWcExMXGWz9dd1N1rtTB6vKqLADnE5b5eCg
PDKmRFSkqIpbJx2wPMYPW5PzeEWdmYwAEvzH016ioJws2J3TnDwZZeuI23k6pm77
TWFNFWP3to82paQUtzfEq/YuUkNzIldaEJB4aquc6EoXHhGj48ouXXMuaVeTP878
E1tSvYR9eustF1yum8tE+9tQ442yvLxH0cCOoFZ3WI61/aF2K/vCrkDlJ57Q70Af
d5act+SXW1llUmZRMfzsSWwKXP+ghnPyMmcVkUXdJEIlchXLWcVkAsBv/LnOmHdP
4j7FpSDovgPqoO9rdH1tUuM+x2GN0j3xEc4otNCKLjRYp6+ATwEmYNG/xPcgjs0j
oAcCEYPTeSVcLSnGIbUgTQ4hCqGQpI5uTyaq8nVH5QZTCaFQZNMMZgiG0rJuKW2R
KOoY5qn5ehxzlkli4NR8GdGLWXV+YzIYcjR4fpdhs4XcaEFJScfWN6U8UXJceoyK
GE+nPNyP2VN8fp6K6nhUeVc58ALLII4m2M+/P7g/hEyY75n62+KtsBP66Aty2dDM
Uky2VHIYFc0sOCRhUV57wxlSNWn75y38dh+6cJffX7zl5QuQ3CC3BbLtvh0C5Snr
T5X3oXREDQtLpyQhQNDQMCmIXq337Y5zsiz+fsmhAKEE4OHDAJz5b41Xr+A5hJb9
/xNWT5gQyxzgtsNtsVmu9dV3017uleBZzaS+nUfOaaQAyZDCsGpq4wMuCaOypIcW
pU7X02YBo+Mxgdmc675XfBt+sWQWd+OWBYh4zEgt78kj+6fVGlPw2uiygq7TwZZt
AVB2RP9LWoQBmJulYEjRANzHVaSMBdlCuIYmthB3+Pdps6JMdhW7388s/7Be6OJw
Wtb1gK1P/XRv5WH4UgIKHk3eSxFO49qb4YkzEZ8QHPzSCcLH3vuRl59f7fudcyFH
3jA57sAvk8JgFXjqxDja6rL3UzTSb8fYXaAFmHh8cRJqhJj1yqOLImafr5DD6CLC
2wiE6G3Oz+XP0wMDttg4dZhHamJBaui1+YL2mAiCA/uLbskPzRjscSL5MIK5DAz3
5Gdno+3ZZzQ5c2fbaWAOOSgL3fzLVwtddJTkUmoa1GXum9+vUoC0um+pbUSxjA6k
holAfZ13wqhyCD8qllndmIIzIeEZgxydTd24pv6JXsjdizULcu+LUeYJMwB2y6Xr
Zs4E3JFBaigQxfIuxsS+hiyGDnC4deWj+tOmmCrglNh1r49Slrk6CDpr40l55j5B
QKI4GpKw5Hg0NlG/4HPDEQiRZsBxMcT7DiKKa7v2kulMwbQ9tqqsOg4J9RNaapSR
p0G5IejDjmCzkRRZ/bCEnQGtRYfLb8ICfiKnpKuJZ+ZmIi8K4lyLW2DS6/p4jSne
1IOmv8nKJ5hAo+uGCCxpAyQTcF4htNukW3/zX3N2ZKZv2Be99mc40wAKynS23vRD
IKRi9Z9ic1Jb5rA3xgQtKHRPgKSskgf/wQWq8fIX5YzMZ/JzPuvQwmZ8Gs2Nw10Y
wOsvg137lG+wT9i+JrUTfMzGgqt3p85EqJH8EJlXW1XNqvidTw7bmSUBlcyHTZty
kC/0PFfviSLifxAJSCFALACOLHK2mEOz/WoPEcMg9yLnyVUrHWL6f0IacyYMfhr3
8ES/L0deFMxKCj3sB23bn4bpgoTXXo0v2XvCvp321KnoRDdbXnGlu9K3w7tuCuAa
YJVYqWD2R5rjwTGZal0BR3C2vFDVD5uIiGIiUPIgHC8w66rMqnbtGmT4d9MXAYnd
5AMeG0gjBYzHxaVgF7xaJra/7oEVFcvXdEYQfz6q5aK/hIRadsazNiYr6+FcJR+z
oI3ByW0W5Iq1+s5TAHUhF58/oN9Jl/b+02Z25dIBEqEpsjnpwbKIQbs6qv0XHaSR
Llse+bmoJYNcFecbhHpkLE2BagH9WtTh/7g25GF8Pr3e4ZvAj7Ts+JqdzJNwnTZ9
PVNskD7dlqM/3csA1Mb1VUXon+J9HFgBlwWWEZs1HEzcVAl1hxX+4onBzOu3yP0+
0F3BG9JdBgA39MSR3FN5UNsRcvmXfN6OmgVL+sKQ+oPj43FEt2WMYOqF4F9UZyM+
UDiHzYdgO3GVcyxGAyhTLJHozL8wwe75yUlmHIv51v2oYdDz4ytCMlY9StKeihVk
hTSu6YPTYOXjdPiN/Ohl824Fx6Gc6Mns2j6EQ+l3vBmwuXF9ZFG4Tjm958iHWQ9o
IDJnj6YxLMICt7oMnf42BcLsETIMzW93YlWSJGbb3qeUBW1RNMixDgoJKwbPcdm9
qVGoTD7tcsAEOBauP0eiNhhWGId8B80Z/qj0hEZwMB6xj2czipKJRj0a8ggj9jkJ
uFo2aWiFHQQSHGlES7PppU/AHLYPbqEKWN8NZ+Wf+L8GojWmrwEgoZwF5C1tFQAn
cKYCcCFZpnKfV/TgtPID3+mWgpWSOB/p5iIeLdkv3e+t8b4/8cc9IK2b+NfvKEbs
ynGk7GccrQ1yC0cvzopq4GYW5K8RpPyYWe2VF+EynHqmfzDGIaQPI3or8pCndXoq
7XZu5YhR2OFKOgUHioCxNf1VgbxDnbbg6TDaSK7Gclr6HxUfKSirZQCXi5YoC6nu
0nvysHCedN/V6pHmv+4bZQFqUYELX79Xn2W9cj2UCOYQQW/sXGfnkgHJ//UzrHDD
wlCAGNl7b1B6B9DyDVWwqqUpwJhuh8GPdu+tuulsd1xkJsyabHhxDvt/Vr8NAf6c
q9RcHvPWg1nINUVRM1eAG8X/XTuy4p/s/TrpvZD5hOvpSZWTzlM+ZeVcGfiptA5f
opxtLo0578oJniGsxyC6faNCwK9GFwQe8kP6dkyjspQxgT874q8zPFW4LP2hYFb8
`protect END_PROTECTED
