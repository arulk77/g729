`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCY3rwU1WIgPzr1Fqs6/EKvgX+30iWk5l+jt+nlWFE/2
bVVhUF8258qybPHW9GJRpIKoq2bVSg1QalGtlQhVZFEaNLMWHir5E0B+bqx8WLps
EP+lrV/bCE6mJdnS7vgNoZ6j0ECP25OPl2yWwOwhWI9FxHXb8VSB486filTvessf
1TRez52/VlDYrzH6UPvOUpESWwK9O90VrUcFapi4YUQzb2qHvQNYVj6Ni2YxkLFl
77xlCAhcwrAZKANyoBIzhpFX9qBGDuQIZH0+RjdVVzLHHnVBY+c3dNZgmX3Gfhc5
t9CAJvHcEkx1sjw29umNGjU/TH0l7cLyu1X5CKUy03uYWbCfqqLGHS1M9aFXzoDx
AUO2DOSyAF9177jSygCd5ifHmqNNOQUF843B88j0SP+6CUtc46PRv4mlmqJIZoE7
gMBDY0B7QkKtBBUjd4OfHfWGoVmn7eSGEVdMbdiK1ETObWWhATCIu2jSNJO3TO86
D75sB+3KpV9AUKMdItY5xkENzFSsEVA4qaCfFIZAmWOkgjrwLD0///+6jJWArMNx
IZqwHX4U6z+dtviwNRmOgvqMsSObOxkPlV77VcGzWMep+MwoHsfTM8kvj8n4b7Hf
tchqUsEOxgYYwk/DRJ1isnVAw/FSZ9CZ24sXdsQgKVCgtAFwGMdF6n0rlvjiAphJ
rbxv0dqe618/WB1GUQmy3EfHWnBruKcozNvbOe0PUMVhR7meZGAMo7s1FkkTz9/O
SCjipaG2HQNXVT3REt3Dg56+/ZaFGtxsth74oMyOT2YRfGpMoBS7A0ffPw1Wz8GA
Dx8YEmh1Nu6Alfx2OaJ8tjAQ0zfxp1CB5s4PPSqm6Co=
`protect END_PROTECTED
