`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAOZQp2hCq9McJftrXbRm2bOAkLMNXE07lsHuh/aNo/F
GocmKBhVpryKhdqPGfzh99UXaaWCfQGTCiCBI9mHNbbc/ZkAna2FBuc1P0En+fzX
AmYdJbYnW49M7CxQO7Qb5nnCD83tZnODICnUl4DMYZWM8FLq7SrLbGKZF/zqozmv
+HWMlXBxm2urBCJlTOGfbqizUZ9WSg9uX6Lc4DilyHq8ZVHosHROt49uOyFjFN8L
JsyhVaKGS3qQP9tVXyTEP1KGPJzUdpkstlA5op/iKpv2S00pRZbiIW428/J1o4/s
7A76wN+jH5dQPJngie5ttA==
`protect END_PROTECTED
