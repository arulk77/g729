`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1ae3wX14jgwCXQLznGvhmRMFXVfcfsiv5KJp+w8uuG/WH
OPw/j1ktu4eD9yGUmr+hRTKOaNg1qwd+CY1yw/+9PgE4GNomsEgnpj5NK59YJ9i+
Pnqc29ExwGzJAt/y45pzJVRzK/asB9rk8RWr7jlxQ52BpBb1LGkWxrE1rpV5CS9Z
cbj7D3ieIfRfG2gmGZSJ9ESFFrxmY9DqT+or4+53OvEBjIDP6lzw1uRv756HCIfS
`protect END_PROTECTED
