`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
BRLRVOeHshyC5Dd0PeMDgisbrfHCHIkDquNL7hXSb5PsoxoEG4aCv6tcmQ0l0hC9
CQE8sXfcC3PSXmvnqHFtuhSjpFOPLWLRuYp6ZhJp3ZqgV+qHofwtUsqv2+Sj41Dt
KzimQWXonphfJtGSDVhP4+y6R9Esg6aWOezD1uzTOdYgbRUCk/Jkm74LmNiGqjj8
GGummrcWR8BjkGOwq4N2bbtJQIUliCMWdQQ5qpIwyfTwfjfUxAx4WXxEzpdvqHoN
omieeb0HFFBRDwC/afAMacVaIN/6gFOzBk2yAwlO0+OSXUSVGZ6KjZDu/QjOogBw
Cv9vdXE9THBgMjzFTgG95OiX4fxKfEksl/nnAHwk2RI=
`protect END_PROTECTED
