`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD5sXR7Faj8SXQOPpkjJvbc95CGQLGOAt6Pf0+cB8TD8
c7ECY+iTC/D7zbSqpJN1OaU0H05ZvsqPpw2Vca736EDLIBAc5Qlkr0C9J2L2SPOw
CBMqKF17hHkwEgCfvWP7I0T9Q/z0mceznmb1DpbbF/LXJgaDClHrf7/J42rRs7f5
+nuPFaX9MgxAFOSONLxi+iYP+PsLUHx+eUYxexl9B49m5zx4iogY7PZ5l2xVWT1h
nBr4GHVFnwciUn8nabPcGHzGJZvKBaAg3JMtkrSuxdOHQ+10wYOXHuU25ZTYqO0h
XzskIKqw4gOdPWvtGSCU5YY3sAWmfJCVpxm0CUj1gsOHbwXLO9Bjh10kN6KKAS5h
8OufaAcwgfSB0uiLhkrJZs7FCrgc/Wg1qAleoHcbiZGw0OpRZqYJ5V8pTcPql28N
aqtlrhu74blyxbrXbeyUhRvVhZHu7zWZtkdMN3043uXeZOL5gk5u+pIRu7Dy52Or
c989xnbKIaq4528ZsCgznUbjIEVu9aJIY9jLsDCKKzlF/veDjAPhNgPUBM9MhPRC
`protect END_PROTECTED
