`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ev3uNhgnRfo5AzKtMQQiAQGd1fhD42DhxRtP3hu2nbxwrpYmCbhVsX/zMch/00pE
0qVWqzhwyqx9EQpoZsfqxbs1e7z+aa8T/WZm98qFPXeYVQ+DGZEmbH+5V5r/8Kdj
40H0Q/4KOTAEhKRUcIyYeRTIZFxB211QBD1fQlM+PeVW0YEGAsRlDsRX2sXBDskj
4dAdAalcYVDHe9c0AbV8gUfHhvxxcKTAm+DDOLgaiTOpnfUARlvzVb1qFFxtXYi/
uEMs1WG11YsaL8iMrhPHniwN5Xk2xyCpBaWJdpUzjfo=
`protect END_PROTECTED
