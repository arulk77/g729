`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKeaNhi+QW2vSH36NAo4qtpBRP98Ckd5BRXdpyuNnuGR
kIKZSuHtrZ56j+2/WLTi/vyPEnyHzg24hD5UHdNXIeqANyD2lDhE4tauAWdxdBhS
Z/RyVFnrdfqMcyZsqhyLU6xypjyAJ3XpKADKJfebuXBDpg2XRaZ5r3fMEfuc8J8g
J0P/1B35nJVzpyCfOfoh4lrtDJ9oMz+usyIm7u9go6VFLSF50mrUjyO1D4/3geEm
BCBuJrBVdWWscZyEgHyyAMgo5n0ThabT61juL6EWPGv7DRGJ+b29wEE9NuHXUuIK
ybL3jkw/AgAENA3pkW46Yw7bxNnItFFdTiXn8yI5eI0IQtlkwSwdvLV2vsrKx2ar
Q60EETxULkh4refXgOYToXMdtFpd23Dlej2/n9yw7AOtuUUR+/rre2AViwA7hnKe
0dqfWHv1eIcimgreEstiDG3iTue9IXKd2ampX4GU0r35oxcuVmQO6QSyHoN3iRYP
jeeIzgrAXlHoZU5leuaeSFxZUu/Ts91iiF/AlKuWzFIDD24S5cSRKTVpYbYeeKdl
v67uPHGJCyUiY7a+ZkNpOLiPd9YizKyDNmWVvfBhRLexbkQb7uVuqGywsbM0wzCL
3t9PiBmDNV/GIglgO8ixKQ==
`protect END_PROTECTED
