`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
52Zv0zYHVcDNOhmH4izDa2pNQZ0zCJQ8HJadoLWiOULTT5CCSCI7mju1qlk+Bro+
xP+Hv5lSVcRr3fKb2MltklbXHNhH5BL1OUGTiaTxJTkRq5XLILnBOMSRa4BCRnUo
nQcHMyfecETQt7ElU6Eqi/Hdx+k+VCbe+Dt5Ix2pfOF+H0dz1sH0WtRtai+y6YAv
`protect END_PROTECTED
