`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePEOeys/8TVcsklfjYYer71Yqd+hbs2m5cFnpPRUibXN
3yktsvWPG/xQWju5qtosRI+8VtqRuxCaxCnMPNBbNSiU3soraFBkMPQnVBg8uehs
Kom0SUgLThVM6SnyxnhJgkFzlKAy4Kz7hQSfbZba8kAWufN5SEQts4byWcE8j9gw
MNhF7i+plJOP6hGCbxb8satA5UADWYVFOVk1CYx8M52zvsIKaiSQpxyC1CDPR8N1
bH0/Foz/IJRVmDjgHQzrrG9IeIVw8q8Ftc5UN94Wx6vT4SAcl32gLPwZEisXWU4/
IIDpMFSFRt4cZU+UPaLicFOMR87/Vt/aC4smmGUcj2otUNFK+yUN0/sgIzIlqCjm
IhVRWv5px4Z2OgqARZiJo0kUkbJN1Z8+0v4phoYyjI+7PqdKw7781A/7r9g327Ub
QS5OkMQzDvc8fO6Dy3hypIxyA7Oe/snvSi3GSibphWrOsUV0Fg40/xS0lir2Jigi
`protect END_PROTECTED
