`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
LY7i9OM+cE60vsptvSNq+YlVZH41H/f5i6aISMs8GzCskXZ3XE+IVW0svDrniHy6
6eqY1m9tlxKsDDeWBncQh34v06DuuEvYdUMbW+rb6Itrg/bDy5p03ndUtDONBEl9
fHsSiMG3Lxsz+DJF3yxkEnf0WrMrWMvvmzdFXq1VfjUqHL7Nyfxwrs2RpGHCYznx
kByLD6mhGnBs6w9KJNaARe72UlqQRkKVMCL9vKc4Qus=
`protect END_PROTECTED
