`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QrWOSRKCfEUd32Yc5WHKz84YwOewGkm0+egr/1HVEnDKRUfKOUoTcpgedvzGrHZX
ByMbb8jgN+ydHAJlDVLdA3GadX9wfILrYfEWXehIKF/Y6+qIYn/wnphCnRZU8xv3
8+td/6MaxKZfssPI2BnJm5yBXcgmyQPPZ1eKf6mYvefAPDvbOo8JL0QjKFX/UFv3
VRnoWi8gDo4zV5acvPfywGc2cwlasWLTfTsFJiPy0QxTHVndywwwJiPSsL0OLR20
rJp0NrDLeP7uIN7woCifLM+9l+/G5uw0XdkN0FJk6ck=
`protect END_PROTECTED
