`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4ytKwThV/y7hCU8eUJFbaxWgqjIx3atUYMokRfkaf2uS
RO00nhFNu8gs9ctNjYaXGdvGmCyB5fVp2okWEcvmeEXxOn0mt0B2F/GVENamQQka
UKb2PrkNyqriSSaIyjWYyI1ERkw++4BWFoDL7nC/LPakt1YEgIiDiFknmZi/ufuc
xL0OcnK4SfZlwbI+3HJ++BOsizt6fHQFOX8/6ujjbpgT5D7WH8bz7nzk2MR7lFyz
yZ28l2zh9rUaLuNw7FMncuyw5ciuGc7nZdEvMzyiLYgbtruytHq78qqiJ2npLhA/
bdGm5p3w5I92eDLTVggceHcp+glJ7b8576ysCY/GwLDc0IC2vVKGqGJ9a1vO9MV4
dVIRiORp7JYtrKZWBtcA0A==
`protect END_PROTECTED
