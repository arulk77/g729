`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aQZ5cXnG7hIkCC2Af3psCu+FoeX6E/o0ygavpMu5TIGF
84+uQvfAObYRdJuACq+QFvWAIh4V1cStts953e2KdZxNe3Ezaaml05wbiENIbBUK
vnNSHcKpM4AHx4YPf8oXEZbUtN+Vfz9+RggFl28D7uP7CxsL2Fyo+9juKwSxDVc+
dAIh/9ewU2/j4xkTQ5eXgnxqb33a6BEBtaBXggizbpa1o/S4Z8ws5sS+NzPkC1lA
`protect END_PROTECTED
