`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBSmYEopXBMWvHnq7o4MHlAsB8K13KApG+vKp6FCARYY
RGaAWisQ77AI9UIopdlnT7VW7JkgflFziPQR+hzktOAEZP2mbVImEBjaRhiXMUuQ
iVF83hZdjX3OZkAMz0U0CzEuFt9BwnwHCfKY7WmUi58O89NxHyJmjkYoMQAsJ007
qfm2uOK7Ruy9B1Ma0JTbaeVXkWKWAZkmG/rqwrffslmxBpD3r5gFZBYleRiwgc2p
ZmnXo86YOEEF1qSpDRH/2WNY/i7zN2N3Cpz+o1VjfCP5sbRG1SDxNmv5ZmAeZKg2
gZXhKlhsbVgrpULaZ8go9iNXwP7MFw2+HF8QGstjF9p4wyqz2h89wOheSq/r74RB
ne8ArlmDdSAGfU/WBhCUy/rTj7+4+viadBXrcplIAt3HGCyikSkEYbAHtNWTzo/o
NcHe9dr8c/DJUt1yESxTXw+02IFzpScYbR4akDgJyVs5peg3u4xVR9vN34LS9ALK
6bJDEThAnyvcHe7fCygabMbYhwE1TA8InPfUK1gdXoIbrp8jSbTua1UMEAqlS1IT
GyKjo1zAlwUBNjUM4OGqanSAadKJA2ZZKj3QaHjqzxkDFHzYITFGoA6XuwPVBw8q
xruZkZLMp7AWjBm9mf81+/ZBwsnrlA03lhzd3o9PPfoRdUVsMJyKBeLpX75Q1trn
`protect END_PROTECTED
