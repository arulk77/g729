`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFRjFSiDrhu5MVk8uCcEfDXiVcj7O7rC1WmL+4R0KPrR
0sIfxPIhfBhX3jxq3evzGk8Bo7BIS+c+umIV4LXnf1vchEeq57OxCyamKyGLMdDy
dPTFIJ0K5ETlEoKUve7FJby/Zi0GXWjAxHsCjZT3UYBPD/XusIR5rGZl4V6R1Q8r
yDm1oy45S4rlaQyYAfyt3rIHRM5MAV8r42EJEwisOS5dOmuVSxwbaP1/LaEleTjl
FRpB0SwSYJ91QFSVxPfjnuANG7Pnc1MQbvSPHvEcWoEvcdF2Xsrxyvud6td6gndy
9cct05e8hDvWW1GCI4TF6w==
`protect END_PROTECTED
