`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHf++UtJ/8NMbNqqvtf/i5SZ+68bBT9MEdWOXq4fxRyH
sLeUTp1iHeqSrayFUidSHPV4cB/CLx7D9NWiBzgtgTd1HiWWZYInDLAbCjg4KZHv
E0VH7i68MyXFu4ye1FoINn2T/GGb9Y8C/ora8r+u2lFBDi+wXsjdbPsbkdK2syMn
ugZq1HLCWKyHxnNkde5LbTgR1yaL2d5oNXSdADIPfA0AJ9EVnIT0mrQE3yvTXmDT
YBNtR8ENe4i8HUXL1bKQE0HDjjni2wc93S+g1ifJO0UAlhdYC3SPN4U6eTxPmEOd
s7f+UgkKXvXL/ODh+8R9Of0p5CL4FWUMi+wSzqbDvmVy7MIwYBK6+kFuX3M6u+vA
5qHNCuqjO3HB1f1CnOSX/SpJvhVVJ7kcj+kRNrDC2Cj8GwZTO9lFL3DroSlJ2I1I
w9OqmiodMbFyU1WTPzFABXVnn8K2xN7RoVKaJLusXaY9zGZ8rzlKho+AvAYNjywS
fW8SYO5kOJP9w0ONfCryZcIIczJlUcgJ5OkyZg0V5mqYijMT3LnOMIieqMSzHpfA
UpHdZwufH6Kb12hTGb5pNOH74x4i3T6VUHoBlY75wzMpX/MxEPr8u0wChEfTRcyp
RhOyDHeWYS+d+GTMkEt3cqJ9fF0FWUKEsrXSkbcYbI2PlE/6+SDDm1UUJAW1qWVs
37xjuP2SYFUHUxE2Qh8HjHns2jSDsI2aiXWm1ykCli05zRomH9d1740DwEwo1fvO
UCz9azdIROB42diOoGXMtOg0VbdQuFrpWBrbnxSWWwvcba3gS5ti17wVcjY4eb4P
wxEZP1XOVg71jzyDtX9PCpptTBV/ll8V9eog2IIf9a8=
`protect END_PROTECTED
