`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJxot5vckwHAjoYZ8fR1S3TCYra+lxuLC+fG5v6Ldqsx
IaOvtb0b0QIDPZNZROVamg5RWkQMYVeebBI1Ow81obwgl57hGCIjtwR85WEYePwA
LdzQFXITm5H2Jmcaltg2vHyleXhU3dw6ADd33fkezg709s4twDiIRX6cSAgvxG6H
MrIxxmk02QkjsW700Bkaut6MbwMjaQlw4nX1y3CBMaK/rQuY/Klyueb/QpkrGklA
OfSu/tBxipdu4VtS8JGgmECqWfLuvwqGmw5b8MY8PwaP29NbmOdsg2uXBUK9WxO4
TGPkmKGOS6VBdbXyJgEtHw6X8PcaqEulM8XRsVROA6qtDgeBTXBmb+K1QZLhEC0Z
wdNPdO9W6LF9ocfm5sfujpZuQrf5ckZKoHTTDji6ONH0+3jhQD/AqJ0GsfrWcmfg
wdFi1TT9qcxOhvh34MreS47y1NgtqDtIUHZdHwj2O3EMaSl4GMNwmtAxckZB+q4j
O/mURFrBje+jXkMk2wsu6ey8vgM6p0tlPWfDcS2z3igfTywON3N0jauVma+MGAel
`protect END_PROTECTED
