`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGekD3KT6mT7wkU1ruDEUhqy3+ZLL32vQKNlvOlUbV79
0Aa3P73v1Xb7ZpDT+ccdRIlzLGOGImHVqxp906d6fEiPRm8gl2lCPX9nMY+H7LYr
KXg7aC8pBD/ILUM7BWlx0AAuH4uKXAfTduKKAM1HrHefF1QToQ2Xj8Ehohiq45/Z
zAAh1B7kfayO2oLY9PxpYadzNM1I9IaqZzVnUF28PD3aMhA2H6mtQJ9+j7tyAS1U
/q1r+nzG//Wsplm/bCFPSlqh5PBhGK6owhtNCKSZT7SrSdIq4RPIv9FFwCvl7V32
Xrt0RdzHFxuItal/ZCU8rzRWp+v4/OQerInKOO2GP4qwAYs4YGtvpAY1QFe+q3FM
MiX0/PC9bBqHuoi/qtBozpsfW6KWnsVs0Tz2AvU4YPrUtduxl0TpqBWkTAReAgmS
SyCCQhvAIBJMhtZXV9jJMd3dIH81IAQFiUqJZ9djp83ojg5xuM483NmbkmTxKw/o
QYadz8axtA4uNc8TKBNUFbLRlcPU9Owdij8jW/SXrY9YIa5D/4L3DwE1WLEgevXV
`protect END_PROTECTED
