`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAeEb9D0iiRG7WT3U5C/WVfT2zPKdzFS6miC62oysDeki
CEw4FYL80u0i7b0Mn1f5xOlbro8PwZ2ujJg2AzMr2SNH9mLcGuN/70TVksQ0b9Ws
OGY/oDRqjJZPTdVHJOWlJ/HV8e8EWNtF8Z2VI5gwqG598lX1uN2iBbhNridUJYUj
uWNKz2PzErnR1vFjcYsMsHQTTCcpPI/C9M1dLv8sKwinbvH0reIuQMDPcbFOGZLy
4+bTZmyK1fQ98RfoE4yhPq8MjV1qHtpD9zGzgQxieVIjFGLc71UOt6ucDtOTsaw3
YS6/q8S6nOnP+I/7rlBR6zFbnZI81JD3on1HKjc3yZRsMitZjU3Y1JB+oxSOoavt
zNirb52qgAsz3UoVnL26gRaT6HTPjriyO04f1yFaSmrIU0CtM2f2HICC9QI6HE/R
UC8AkVwIu7Ka3/OMdBFzXszJmEjEGp4IQ9GKyFJJrValuJzcmw0pV93RBw1mf7iG
/HJMcW7mXNJsdW5zsREbRmGktcjjFYQC7CUXk6hEmcuDkdG+toj0m/zwsXg6uNve
ewO3owvQ986hb0xUtiVtCrEE1ecP3aDHHCyH5u++NJxhOeH+Z0ZoOlFY8yLxG0Ya
9nQcfEZni4fQaMamSn/i8H9t0FpKwh1up9PQso6Sa9FDGjUd2KOhMv3fLhuSNWi6
1eJwOCVXeZYoY+Hd+IJ+gFerIwyUxj/287D0cfmVq3ZpmMlVLQkwqy0FTnDaG2rJ
uX3vJfr5diXiyJ51dql1dBTfYv80EEOShhyIh5X0yZzdyQIaQw8hZs//FWyv76oy
yFx0Qw6vdldySa9juOXo1wFBb7oTgoUiELKU6RbujwwIpmhT2prKsD+LIJIlyM4B
HH6lJ+4GZuOWiRdyUSWs4aeUPJWNMudctLdVkhUOBKbgW7cj/pty3FYeHARYBiFi
gpVJ7dwapAnSeK7UMcqZWJLBQOSxZWviDvtX9lH2tuY754ldUmfbPMSsd4cO5UzS
7njOQ4X3f0WaT1s7O/cXGyDUQZA0efcD+F/cdMIYYJicrtOe4DQJIiFKTHM7Z7MF
Tzc2LM0nXmSzcTgQj3+dP9vuCq1pE3y+D5w1QCFTV+Zw3J7d+PKdEFYTqi/Qr2c7
EeKx4jNfDsCEzdRO99nljLZllyG6ADRS5wU15+6HcKPG/L3W0dfGnaGIxf2qF++B
DIAJf4FJIE2NS9jJ7rhcmo0k+1CQdIoQ6D/wasJNt01bqr1P8gBgO+dNtcGG1ypQ
1ZG9Q04+Qe2mEYapECleO70W9qZJLI14aHk15sDuj96OcABtrTT5fDZdMxnuIobh
40u5IRand9IPIfjK7R7kndDO2NsnnKs4KTwK9oaRSZ7f4007aP0+WR01mLnZvsYf
rhOHhZYFfMp0qMaLLyntQYc9AcRuysKeWjSjn06f7HGHv2lDJgoINuaiQ35BFa8J
A4vzBvmlsiNf7vmnl6x1iCBk25PD5Av1pyA7v5EUp8B2kWYufG282yic+jY99lDB
bjtV7258lVtFAf/iOS54g18AIU1xucqhpapNXm1+Q2DVzvph+DvyJynv7/72zOs+
AiSlyuxiJQxMNh78SQ6zdlcLC0uKgcP4atqPmXOv3zGmj1xi3wB2uiFQ7qCpJ2EE
+YCPauXYTcZeOxil8iIh/i//gYZW5nfDh/0S686GOIf7ytloDvmyzlvOek6bTXFy
RYE3NGTF3GsvN4OWYWy1LRcXbfXUuo00HCwxeS/QCv35/ySgqgqnsXKqhCYdaKwh
bfBu38vDyqb+kquH38XiGosd0k5ORuPTvaNn6zNb1+Kt8Cp6AXKOu0GS83UXBhzs
mdFbKVogjVTDHWGGQ7u3HbT5u7T48dpXNwU310/qA7O3hIzg+pKGpQX1xh6EI36e
aWgCCk0LE+dqxgAW5CTcaSXC11i5HQ0jTnuXeyFuikqb3DpRZ4FWgKIOPSctqYJ9
tZiqkcAQASLRTFdylNiMmCBtMNM5O9SVN46ldBKXe9e3dTroCIyTqbX+Ke/t2t0s
gmuXcbQgcIFanAX7WV09dhwTOEfy0wIbeIqwgzC8qQPS2Jl2TPIUHTalMbEIok5q
YAeE/nBCKvQ0jyBPdbcTbigqcOxN7wRxuKJv6fuFKaA9S8+fsnHLU9qwSsXhg7Ss
Ps99uTTX2RpP4WGtjyQ4z9ZoMot+/rZhBcvojfPNJPvH4Jn2NNNexXh4bpC5TW5l
l5gTab0jdVglLQds7Nn5FNgTfQXnxYaLnsT1HeKpAvc5d/q4NWH7RHjc2LH1b9/P
ia/USbnaQhJzSYz9t34Q9enSfIQcpui/Gz69e2zFuFw8k8aPxXPc+ogvMkQ4nFRy
JLfgYunHr4nMwEL3xNCxmVRdO2xO9DR5Bm5BKNZBFRtg2eUkToJkLWOxZ1y6TiiJ
6BgZON3olxH1ImiX43n8Tgwbl74gT34pv9HAU4DwNZLFCW5K8iv4prU4SPubn+G9
5O/DZZzNsI/79hy9MGFNe3RYbOMttqLz0TcJ/tcwDsTiL/H9uQoxuyGJ1vy+2DfG
cVDTWIGsXnsl3aLCeW8DpjMjL9nJiuVMRyoebyrWCYloWP11YFcgXpat1L6o/4As
3Tn3u9qy0hVqz55/JBsrDzg+/hYMpkdIclSLR8tpAxh+4DLu95gvSUsNKLeKgxj3
nOAEaYgdEdSgezAlt9/otUXcXpW3lVlas/ehjE7OwZqET+D9RnJT4S1QbmAt30+C
uv6PCPaZP/k0EkWLvDytg65QV0+XRZ0eeboJiT4PYWJyKj2vAs+lt8jtP8z6H1JC
gUlvX3dgIjcpK7A6RRoRr0GaAIjiDV5Bfr6tjY6RuJkudBiE5WPfPPAI2jMNiavZ
TrbOtx9daHY15A9GKjIj1AKryr/4d2VhhuZUHvzyxBAzzhCb20SiZgH98mDKbBgc
S0FG6YUsSqf81ksP9ozgHnOgt6IxnxemXDH/c+XdIbEsH89ywHYEDBSAAIvpOFg/
Jz0z7pFjEC+H5xMWvH6NKohXl8b5jdS5SAbCy5MRU4B/gwtfFOve55j2d1NQsNyn
GVB+0vyiiTyGLPMwFP2B4lFYHzMaYttF8BEZyksJwxwqEhRvrqyI4U8CO6Wq7hG9
Gsk6XoIv57Nice/htdQRFtrF7WYZsZkh9HDZXtQZc/RGN5aDjxBcDcEI8mnDfKcQ
QTzdEmBf95FqXvusaNyGj7ao7xQT7GeIXszssm/xSw0fSZUQpL98gmiaVvWSa3iE
Wj46FpLN83tJHjCYU63uDUv3EVHIh3R22Y7CnrfGQcW74cMttvHlVvMPak07YVJ5
/Are0HIF0PQPgxmIefqGUv6HJXWkumpwvKnQCvYQuBMsXAfg4kv/yMeal+jHkb/S
ssJTti5PzOhU/0LyVvGIVsFuDZPi9f45MGYleBazJfegfugDOXP21jMg2yTy+r6Z
O98My+JhafKXVJHo4jif4dPDtdo2yTHmyPkrbwE4sSp/Ku/B1Nq/xLST+V6yc8jQ
W0GbQZxg6YWQ4gFDRcOSE8K5igxEAkXnCg8Ou6qQDV47un/43ukAdpMMWTx9RCRS
sSSjGEZFu4SIRLGyEzFWUXJAwGPwCIt0XJiPiV4VIXA/MwDG4TsiluR7fAb3Z8oH
czusqboQFV4AiornWJ4shQprdBlffh0JIqGO4VqkiI6cXQpoywcwNOecgCu/BM55
C7d1Im6u5WUfYcqvfE2xwIIEZPiltejil5QBcv4O2K86McAeNw4041HyAw6P3YRN
9udeoYwFNL0fstDLmg/w0urt301eqFB69Sm2YYc97odPXkkxzvuiqpe4KCAkWgZl
1HI1wPpUs4wvY+POsGV11u1qlgAiAJq8gFuGnx+UoZO6RlAQ/rGpqFAgT8zuhlZ1
fXWAKN3GL/xq6OhO6YNIoWmp2wgctoVQ7zMIMBFfS4YAYZo1VLIQOCeVl2Ms8lpL
J8NYpOZwzZPbZ27lHrza3ar9oRzTXdc2KT1IPEE2660JD6aWj5QsK7oyF9OccMpK
vbV4ySfpKRB0Ww8kJK0hYeIS2PNx6KVm/jLehkEgWjPW5WeOPT8tZZ48JbnMdPSP
rwK3lwt4n2MkWyUOf2DQlRtD9qzreZjqYGCOKAnn7KTAYmP0O70JK/sMt3SzN4h+
CCflhIxKBOtq/EhQm6ZTdLe3/QVu0Zo7kr4B+Ts89l7HtIcaLUy0qaUZwxugkyzu
H2auas9k3GKJCDHbr3fJt5sjg3Im5fkceJ1J4v5y1oI54ok+LcNnIiM5gOoJQQHx
Uk1Pe3eERrNf9rTeKoPPz6Rrl+/Rch+EPIEWhtxNhqQP+cTzb7MknsmB//qKjH6j
bgg51AxW6WA4/5J+tUBxGQ41clZ0JjA0oKEpAQzlWZC0ExP6a/QVql4HQPAIsHsI
f9Qg67GtB7UYXJYIhlqWX7loug4DdTj+Kovdx0lAIE/sr7/NLVF4sznL9g0WgZ0n
cIDupBOo6RyKuBys0ey2edlD7SPkPie3Ycb0B85Rd9KE0UnFnO5uk7sIwNUStIH1
CfunBDQ5t18zCn8Anj+xz13GlyHXQgS3IIuaqugnnuu/tPPXFDKFzeViKTaz4qmZ
nn8CR9atJpss6Ufy/ZtC9RFT9MxdV9UHb/0feWctdHr/sdNGaNY5jBvBoBcdjQB5
n1FUFt5TYMz4I4K4eonDl+XUUkZ5UxMFL1vGpC4hktwGs0uLnLpnhyvV9kdASl8e
0nKCdsTf4F9Z0fusAPxjdXRbdy4bs0OpnUkVHkRtL006f71SGIE9CVQmzVmtQVrB
kjcw6QSnw0lIN+61c+F5EhVrsTCKkQsWBlEcKvQkUAoRnGo5berylPwpVjCAH3Pu
PdShdyPJ+bekAvCNHZ8e2Aq4o1zNRc2DFxI+OJGJMLZchteuIHIJCWv+HpHJNiYx
gbtWVHrUiqdEvBvziIkv2oxYidq3N/v6LGSsH2+sjgN55H3gNZpKtJkqeRN0wHFi
xDLJa4KM7aGn4AGQWxgGfSRr4pGvseNNOWyGHerqCXZN4EOZJ9oy6kd2u5+ff6tl
iJI0U2pXIN10mFE/rOISdA/YlYAGFAqTwpALskTjQYoCzDNpPpLFcm1x5k3/hSAm
nYB++35I8aqbfrJsFo/DRKRjzZvnI3/aRoDanlwT8ZLz0+WDqe+EoruXBAtr1ult
sS1wjmZmCePADR1mykOjq5rlPUHnCyQrJ+XmSb+P6ljXbzI7ffrPXKW+r96cF5Ey
VLT1cBFfInMTI89uLU95y3I79JBSUz8jLG5C/s+cDUcjVzZaE0lM7OF9cPY6kb0k
5bJ2FrxbdPAtgQnmytJ/Is23051t87sLoJlglhMkLkxUpfFiIC/F7aoEsQp7b1iL
ysgOM37HnRgRPYxcva5Hg6sMLpsltXD3wdQI/9CqPCdl04jYjwzvHiIOMBnLjLgl
sewkBSEZI7PW6nL+TopaELH1xRYph3F6wFSd6z0SanIGp8jStsJIhPU9w5aiudZQ
NTEGSatly5hqdSTxoIn4jJ/6znVkDHFFV03aLFqobfU=
`protect END_PROTECTED
