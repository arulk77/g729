`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
SNvz8HrX5+iYiYsqZYVmhWhzXGffQUcr0KcLV1Pu0ouLPHk8kKZfendsDWfQn3//
hokl82uT0NMM3GJQbY4ZkP9m5+DODkEwn1Y9lZn0SvIMOR1yZdmgMea1CPq8+7hi
sWC5OFL8MkEAkUoZXqvhnWpY+R2rB0WCdfYEl+S4BPqhrjsyKUR2jfzQT1G+xAeK
GDhiaHkD3G36rScCViGyAAALKdSlqe9qC/VHUWnoKc8=
`protect END_PROTECTED
