`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOAQ0GMC7Y2edHr2q/igK0dzNiVv7h7lT5KLPgLY0SGP
xi4ve7OGCzJAUKAz4xD4dhDXW9BsTOmN+0w92pHOcwVwqSPS4fWri/7CWMrRAGWz
1tgB16cs9tHOPjxrij3N0tqMHfAvNut+5exwt53wecSiI8U/Ey4iqUSYmFySETYn
/+pMY80j1JBJ1HM53gDzLmcNVGUeEjtKESvRoCWHzFX0zx1ZFcPu6XH/Zp2Asfvu
`protect END_PROTECTED
