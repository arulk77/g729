`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4843ZI6oUCcS7BtLW+J1YTHZJz9Ba5ZnSE+ZNK/cO2kU
XKA1jSA1YriqW3Fjoqj8RisgB7RN10wTJgZDt2GIi7THY8RJm/gObqKhBCRx4c8F
e3MmQMuOezCCaVqWv/KYEv8TuxlOrY93/BbV2zUo53y5iYPs+iuPiQysoiXTp4Xc
jwPu6vdhKGDeHSV7CS1dvm3PmCjYXi/kpiUrgN6YOJbv/nrYyOQLXTnl8Sa0F05O
66IW17iT+3JN6rCQmENKkQbLhrVv+irgjEJM0V0rE4prCzNJItGVWgUWumhyzSV+
mL63U0jFAmNW6US+2I2ZkiM4RefLh4CMHdFCJ0xCjUKw+a529/bxOyAKOGZV2P6B
iI/b1dGMQ5faQF1SVKENuw==
`protect END_PROTECTED
