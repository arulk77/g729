`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
wdKtYET92IAX2YgPYYR4YR+QI1Q6Xv9ECmK2OkqvCShaBRLC5XUTTyAsb45qzoLl
ruculr2y7VdiEB2d2SN64a+CBYOz/LkyauiyTVZv1i0VmZdOMsp1wnqNIhwiFM36
6WdV0m7ihDAzQfRpbSHLKxm59WOd8DvLDQxwgO1VJQKcZpL1nG5QTwq4MLVMxKAl
iN6MXYGHUb/wPRa3bl/9QrWUgahU/2Xpi/empSScKBBK0uy2QCVmo0ysirVqcvXo
siUW1dSDOJkENqu6yHus/HwCv/tC4+BnN2unJv1nZmr15tNExYdfaFcCzZQvMKAm
l3EjzQoybriYRl7U5fQjWZ7yMmjUUqzNTSD/W71/otO/nwz9B6A9b1ZexlbvUMZR
ADvsiBkLZUrhnRUVpH9vECePQ8RL4NsLYtTJt5FKVfyQYrj4VRJOzseJBL1pIsNv
DSb4z7Pl+aDy2g9JoTqRvPKa0g7BQFB1yPachHmSJeg9fdo3xsB3qwG3AIf44PgV
+WApEucT1eabaWrERtGnMDN+KZuSxKdOpNAcErJzheEG/IK2TsHc37ic5yKt2uQU
K/YapI87sEYVR+QiNFpfNS0OjTvB8Gi5t6yGksNXU0Z5UyLLftSNWTjqN0VrEoyV
DuHeWhjjQewQLprYVbmussIyGq9iGyP4FMOaHLmYKmYz9xUa0G8VQUQDb1MVlbcG
IMIDr3hZuD1J9QRrG5RuDs02toOfDCMTFMjfBOUoJF0ENWmXu3pVnIDPQf+2Mfk5
capmFvIKUZrG/B8dQLIcPEPDLhQ4f+c85LvYTBbcgSpAoEUt1MZ1XI8lqKdkQoSr
fk+Xmc5dEYeogQMkDOpFpKvEcnvc1DCtcQNy6QN8MSyor/uCL5AbLvr1J4aIeE1D
RYBwlk1SMCXkOEQoWAR36ovnaMLbbOpwTIbWQxPWXXTaEo6UEuWepD2gvYYnTMBh
hj0tbjsTpBAbSJLzz9Wy19/kfpHfmr8UuKW161nxDoGybJsVgY7aGHLBEhTLtrWW
Rs3PIWW5UXoCpBZuMjBS2EWJxIdD89FNzHQLKVj98uPnrH4XpQiQbuAHfMj/0Pcq
rMgs7IZNHTPNa99KghJEx8Ymyg3JSsVIjjjTtvKWdZBwQhVcrWGMBgox9OBEyLfA
yPDThWLgUNQV0WalVGC5yZoryf/OmZmRPC+vtxnb5c4kazfGQARo+Dwfva7Bh/7s
hD+DS8mPqyJDnJ/zJwsoBMZ5/3pZs8epPz+akZNOO3MkOn4DTkA9DHzA5N8wSNmL
GLsntTB5f7+gcRQl02KUyoIkDL+JkOlskYcde9hTeIblfu3/z6+fhHp7wPdMTBXt
x05NvWhZ9UKlyshXojDQH+so0Bm35W0Pg2++Y6ApEeO00/BlHvMKoRGBKbVFy7RY
nnTIvf74V/tyTv/FOJPwq/zTAv50bHlCTORrLbtfktVFQiwkicCaLuUSY9TDQdpJ
xjI+ob5SjGMDBZ2ChujlpDJvTNKCbV1lLU7hQqypHDWfnGugBrWpOfAw+YI1SQHJ
CMxJ5CUWtuxSXrhx93C8h0lMHV/v1cY3M2xkC5cXLMaLIDBTntnfTP4GqtKUThCa
cv30BuerRKR7LGtQnpAKvZNVxOECdlOziN6VLHf+Bfs7UJh1sb08refiVFYQRZ3K
K9TtMqC7yXEf7MK4B8pJmDiIAihxDWd2IdX4Rq1pG4q7+J5vjztsdo85f/Rjmcip
xycZPNNJ3279FSL7yUcKfRTo2AHXfV68WzcUB35QiHKG9dCaGUaa2uf78C9YbnU0
taLtRNXh0BYawH9LmN2+EaAy00C7MYzh4TiGr+HXijcnhycSMprQKA9Qx5J+ZDEa
StmTBgRA5Yiaco4tFvuwmuwqgMdT/Asf0faILAQVcXpP8k3sxaR4Ib9LljmTnzxk
BUYBjw/oOSUxEjOzL589j33MaQEGSAZPzASZ8sRh3JGUBAMzLX2XOH/JV2BugUX0
KZR7xKyH73FCaLlOYF9YPZ+bZeeK3OHn6McRIA0LW7G/Gk73QXIii87YrCxIwbP+
JiHHmLMMlIhOTsbz0CfW84I1wa0nvzLwNQjoRt7mhwUTrBe+ALbBafVEtRL/QAih
dPGA7+QB2eyo84Rc1IMuZfnqWzcKFBM+PVVBuqc+ul5l4YpAe0o37cBS3ewgMUtt
gMQ/f61Fdj1dC0mlLeQsoip5UT7/KacI7zDye8BkCYe+VZSVp5/WnBIFvuFMg3sv
3s+1NED0OYZ7bv46NxDXnV+fe1cyBywzb634L7EOsRGKtsKPQfUAHRhzryCIZI0x
VTqSgbMrjScaxcjDbjpQoT9715E3dfdbKTcryHPN3WY9BcsMpgbqaTBmqu7MjZkD
LrurvVx5oxYr6wldM30Q9Vjfmh1Y6Oa4w8AM7AF/Vi2fKcOyBen7PSpJlA48OzYU
MXvsUwBd6tPWuJ7tu3okgApFuW9DAODwe7ACmwGT4OaCsvLYmR6ktHDPRznjXnCP
a6/0w+P6T15cosVMji1aGSCXzNxh1wO5kw8lwMkjdzyM4AghB78j42HQNvpkW9Ie
10K1tBXbBEFj+PlEKQIyFiqjyUh3TZTOgtj2vvp/BxxXHDHAW2Grh4onFq1rB39X
j2oW970f2jutamEobd4rat3J4Unh4CzRZHMDjRvNOaG93CsdWlBXAAaTyYYQ4XYn
R/Jt4ldKXNuBvGuLDn2Rn8e6f6af3K5ZbuS2PRkY5blm43yJbCu41adxuHdl5fkh
8g+C/iQwIgFntyhieRd2NKo9Wy79U6ocET3imVMZpASn5qHEazcUolbx580U1+lL
luecw4Zsh7OlMOooIy8nOx582jjm2wMFqmPSIEbgmSj3zWuhqU/FeIExiERkkpts
iS2Lm/8xRbvlxkwx6ObnLT+XUP2sWbYJe54E680O3Ir6X+WMy9z22YpInbWmUQd2
4je6ZndxU7geOHDm6MUZVEHmOh0TQ6OXUiwEgrXFdt/ZCW3lkQbJ7mr3OIQ/V4IW
dORqgeA3750MNCFnXxm2UoDjzsdqZqJO6r9aoLj3tI24HZHck2pl7MFazZtRf1MG
0v1CFZ5cvUq0otgP6xXqnh7+pQ0Wb93oeyDyADboFiPGg41DtQn1keT8zb468/qG
+KciJw4DDANjd3yM0bJejyXN1FuGkWSwDEtKCBRPF0yhFJcqlamZGbCvsnZMBirs
M4nIaBxbeFDgpVDEvrLq9Ae8U3s4oAtOF4CNWpbP7nXyPbJUMnEzKX0C5TwtX7C6
AxKxDeDf8jL1hShAT9/fFh2FFz3VH969qrCouYcDEK1Q34d9+uyGkwhzSA6sefGF
p7I3/gcyBL+rU1V8mNiUZWM7nzrprANIMwfxdVtURCqfeuQRSaj3ZQMzoNYXKOTl
aZvInb2WxSt0RDDB/THW/ToUbfkYaUUXNM2ik5Ryq4zQOFfLG4SvIkZtNszi5Hgr
LF9xn8usx6F11wqyU7QVIZ5LWoRgSqxy11QeNz5l7QTYywWxYILAOZDSY2e79Zht
xGJP6PsELOPZ7EXdv5TaUY7PDBPYtlX+tD9XgkhNn+BUqp77u1NfrSvnSdUlSZVi
HMTapEUCMPp0XYxeRV49sYievFZHo5imLIbU4Y9JqUBiJiO3TYfDkh+63siJvxp+
JFmSrDtzesAoz7uMVOZhb2TYSAwlIo1gTvPZxbQYs2rBmdG7dPf7E0xn8ItMvS0R
mkBHhnkt4Z6FY1XlyqiCkXjWmUDXCtwGsk2iZBCif3XWj6tY6s0X1Rn9jkUoVq8r
fGRNgjwhQZkRmnXQZcj6JSbjeoUoz/Taupr9MoGBotASKTvYYfm972Djqv5T/Weq
gsugKBnq8iMpvKDE6Nxr5CjXaj4XLmCPsQq/iWlX7lCnw7NbM2UrNeXkATzUqN8Q
MB/AMv7/w1ihCPzK186cLwoFBaeU1ThhnjaYz+gin5gXE9LAouiSOUajbfU+L68y
Yl9catJuR+Rg6cjI0Z5dJgGXrI2ldLzeUUE0CNtquBabnEKtcCwTgMsTbXEEVOl9
TgyxV8imtNXe15cO5bNB5Y6vdAJN7jyzmyUiqlp2t1oH0O8GFEWv6a/C5CesMWvG
2FTxUnJYgiTYidHS+QM5b+cOsjwagU14uu058IPvUHIeWT+VNmd/+fjjJXlnGyAB
8BX8+pnAAxO7h8IzUbTpffnNovsRbioSYQNIhP62CZbwxViVCTJYN3M7xM51X72I
2Z4Yb0AxDc9/KqumpkCa0tMfol8IQsyoiJ8iD+N4cM1i7AIJiw3aDCEYBB9n3i/j
X0FpBYA1S2FZ8lcbRCCmVoo6UWIFEeAaxo+xaxAM60f5OIX/VcuR7vzVlPRMXi9N
qg0Nzsg2k1JUdFMZqTAHUadQ+VUBS8bDAgrgX6Mm+W3vnhmAXhDKDcziaJVhK8i+
bRzGeF5lPcRlIY2SXFkMGFwJF1pR5S7N51QJF4iQzxeYMCmSLqMJmoN51dv50EeU
25i5kRDovqG4WX+7ABVBFIMqTfyZgMEWSMF0PdfMslRTZvflLla117Gm+cwXsTTv
PIQKwIoFh00AFf6Tv9kcJjxnnd8jvT7fqx+tJEMeJeXDGCzLUKDvz7jeRGTZdQUg
RZ4ksOZNkrfIEy5uwjGpMq+oNF08zpgrlFw/vau1k86ra8bAimHULSXt3cDyYD7V
ZBFk1i7t1SIeu8hvIs8FQMhPS5qAYuk11HOXEQ2FibwElRvi21T+tod2xIf7R5vC
8zOSzncsYyssynV/go7ASymZ3jntrfeCp41PmwHg+KfgFH8w8a+lz4aZgPYQ4iVO
sa5WpCLeWhDjOefKAjqNmDd8tXi0z9rf1uow0LAzDOaZnOAgxmQpl6+aQZLBzGo4
HhKwJwhe1MkQKVIuXFpkObDMhTIsyHOQT3GccqGuUt7BPmygtZ2pxDQQDdyrMGKI
oXav2LnDRhGw1bTMJwPZt/YTHc8wgZp1XI9BlhDW5mjTNIkq7F+tquVDOhv8/Aqx
zcM+ShGD3tVnyQ9aaod15iG0u/YKPBqgUg3rWMP8rr8Kk4oDQlud6+zDCyYgLvo3
FY9UNHyhhqpYHjs9VS0ovdJTpb2/z/bp7hNSV+QJa81saPakJk5bxcnt/1y8MuoF
irGATzo6wAwmO62XeBtfuQP8AZGjfZYxCWI9ov5uh4t2LQjGNIeHd32yS52q+tUP
E0IcoO0YuCbpJNu61NqE1Nk4I6rYt1YS9zDFwZoBlHmaKyIALTg4vlQk3amLr42b
9oTnRmV7Gy14ODFP3E8dO0fuusI0S1cjiC9c+aCrzJfFOWknx0s29WhMNUrdhQ4W
kOCkNqpj24T0JEMCfMJ+dsxlF9ZndVEH1ka9eGfIhttDY3S13sKtMZghDQ0uwDC8
rdYu6zed2CO3SiTzaTldWo4Tm17oTrBftxupDtF9LkztTwS4l67SKw1c5e9d3/x+
4fzmai321tnbnUBPu03lDVkM/yGthKR9aZq2FosJJWgmrcBUvtPkXlHIZPnyeesa
PSRJFGGAqXnn5ZoxIvzb7ElV/1P4jQnBoEiaCcSblHS2bLBPcGeNKLAOqIRO7oAn
5u6SIKL3JPzVkKvvMDS6H0Q9MhTqXg2W5dF+McWomMHDFV6KZkKLictC/qN5ZM6M
Oh7OLv3M2ek7kf9ijQnGrE69So1L8aYyorbOUlpYamYgFfk4hRGPYLrAhMrMIdvP
vwRDI4fcTR90nzVl+8h3ZZUmyptIaEBues+zkLXZSJxO/4+zTKgKpxqMnexWIzQb
B85OExI0FNhLZM5Dnrwjnym+95D+XvdG8Fg8RQs4b6ePfziFAS4wSF6po84PUGwK
GplT5zh1/OFZRCRAU6WjSL7rZzMcppIVXV1s3/DD8PeKApldJJhQq5Ban/0XD9Gu
s5h/46y7e2b/rEZxKY80jUKL7lGcI3l9ZHChq/y9Oy028vN3IGCescCPAUEAmcad
PYiPTO9oTLjJsaXhbFUeWZyIh9n5HHQ8vtNICZf074Hhepl7nA/X+Bm/1pDHLrim
wbwnJ6Ky4oYnbV3hsFLrpHMIAkEMofxM8ONmB2o6yBf0Npt6rcJHAuv66yJTh0Y/
ijxiEY2SgByTJm0XtLRayL80qi9iETeU0D2kxsV+TV7VYKN7X24ta7jI8WxRlb42
rCagnxio6p51JsFOxm1Grl9P2ZBVmu75zt5Ih9xX7qKtjqlYZigkpwCHJXskWqRP
bvjkuDjYdwVqsewJOSxj5t7eIXrOqraxpQIW87obCJ+mKrbN3Jnot800tA19tDdL
OkBpYQVmhBwZthG+vN8VVrn0Bc+LgSqCNNNVtRuJjLZgXEWoj4jDa7WN4Oof0gI9
FdL2azAB09Ercn+ckoYsdfdvwZ9QUigKRSHZGyh57QyY7wst9Guy6KCy06MBvUXc
RW4rF+NTLd/RzqnJwsQhbCG9HxBt/RtrNKaaQho3NYSoCpPoWe62J391NEZF4ol/
70qR9kVZ8oH3njncI6V/etmovxsQdMCm2YL3Yd+c45qItapbBNm1NLcpJCY/NOvG
xi6qvlj/kSBqaUDpRkd4inkDI0pDX0p584llvNn+7VwYEXsFJ4mrUvjD89qdE870
0OSeItAss4yoLVSvKhRMgkD//P5NwruJDMzUqvgLSc+Yln1k9UPI3KseByJDX2AM
AD2IGWvQfEMOEOX2eYmqi3yvyQaMCPBuqBgYKe/SPETcwNxE7EKfawdBBFhqzU2t
UrK2HMKfmWa+J7ik7fry8NybGQ8oL8XkKVpgTLWYRy8QMmAuyiHVa1JXh74oV6Sj
HvslWbdtdS3tGrN+w+CELogupWcIE+P7MVeVrvW5hEDH1cSE9Co+1sWWYjow1zAt
Ty5jvdpPof92P6D2T+bUaQS0wmtVHRCSKlJdncNL7ubhptwMXoc39Gu/43fucet6
MUzZ6FS0M966Nqvjh+/3HAWzvCAm1MYYxbKSJe4qTsphPwsmYSS+8SG2TAlzLbqE
9Rsn8CQ2KE9s/lP9m95XNjvEv9W76zkPU3ZLM7oY+bnJgPcEQmOkVcscn+jxtaaP
Gpiqnt/I7HyimQwYXzAC7QJjTQW10m9keOcSUNZnWv+TKoeHNneTeTBTth8s8hR8
qohwdp0xrj/OB4MiQ7bvGGbcDTKep5EHzra5nly/Et2Wycl8xxBLVlGKWgfFv4MM
5XH7B/q/Yvn+vwE4eRyapRLolwsedzgBtFaPEHSnmZFQOaopZ8jLFlHzo9aEzhcg
AnVgwPjIAjMrrScnJ8MvNiTwHEmRz8IKBL4c5fwxkbye1OVOASs0pql3BlZBokYo
qipqi/7RTUOstUb3LBN7vWCMMooWWg2ZCLcoTgad5bCNkmPE3fPVkdU7+w3EDKLZ
zbhTgYms/haJlcMc8KXyf22l7DHBQMRti1NAZ1zN1KRrzbHOie635P/cB7q79stH
9GPRAJ9k/Z056Lk4FcPpvIbFm/jHWfT95Z9e6AmXMYqHWyvufUpx81dgQ0gsonuZ
s9EWgMFhrYH2i96RNew7w4I81JRCrNfeHj+Xa7wEb3D5VNT3Y+F68mjXzyP+HPaN
1SvDJa00yC97TO77JTjBRR9uGlN2FRZpjaA3Jd3eIj1EDOrThYqdyjvw8RisZtgq
7HhYwEqTFv+t+Evu3GkvxGJwllGxtXWgEWv99fTFq2vovkZSWT3/qo+fPBi5k5lt
ZYiTt/fSh0cfHkCTigRsoLbYlbUO6uon8avS0Qk11vNXlhz/5LMbfLuTrqgkflD8
ujo4+8teQtcEAfy6sO0KSGPa6WA7rHRT6qu008SDtF2Aiz002NLsxIEUwcvtwTab
HKeaYW11CQahWoedK9h8Nlf42eNTx5xnkZZp5BJF0tKX4cu8TCZ37LrlwabNVIum
3HUAvq2RtqEgEeIxgxo0FhsCtMdhOZUDNqZC6mOMFgwz7pMS6CI8BNIzf+AQjYJu
3HGAwfq2aoyFbVnQgC7ev2bdfr9ACyz2Zwrksui9O4QkQPRzzITuNsGzV/7BY9R3
HA8BEs8bNLDWUnaEjYQlQ4kJ4AFfzpK59e6sJnR0B3X9sJVUV9wNSsEK7tHcXIAY
8+8xo2wOh7taPMoIGdX3A2OeNVX4fIFxqU0LT5a51kjHbvJcXYhv2cOxjIZdKXPp
X4DV47GnXB55hypJlASo0b5swbsNfDiMIMULa9OAi3DArVX/wlhY8FUMg9LjG/cb
ioHsitzvt3IRYBtpP9udScIh4If8kLvQyT4v68GihJ+ny4QzGN22GPBBL2SqebK/
B1kkMuxye1kpJvT3pWEaWLGRlwWTzRrR9dWB1TaTL7krmRmkTAM1RzDJ5qW8DwZa
cdil0CPUxIEt2iFLUGe7uw61n0SP+1VNwhhVjA0VLUauy6zCpls6DyzS5E+hkcBO
+ear8PYFdVPmSGOcLjkqy4A+3wKGYkGOF5I7I0S2JZzldbiDxAEzw+he4tUINtKq
1QhjGf4PAJeMuhl7QF7k31qHBhPjcdrS+qPqkE5w3Yao6z/HTH5j1BlLDMo25ox0
V41f1rhRvnOqqTHaMdLt9/sgoGMsjJb13rB4prj2FQadpcz9eoMzuAFNJ58oZIR5
dBYVaBp1eQjdb2Uhi4ZsQHt098IlyhGmUo1EeedH2rgWOQbs6chntawQctXY7cPC
oYxEkX5JEhuQCVUo0IJA/JQ3/hc4qkw1jYNtYCMrNy5RtGsc3tCGxigVP2olNzn6
u/oUleH5i4zugjmF1B7X1huxXDYnsTYyZVcRTYk7PAEbuXLH0vzLEUlngxWF+5Gn
CLau2nOoKOjCeQvmbRAaJX/VEh0zvCV51JOnxS/N1HKTz3r63XARn/Gi5AT077Sr
cTIoZGtr0AUXccXDIJCzJ18nA987wczBURPqvpGCtZiEsVAHv5jPoTQFqUfC0Kce
PBER9NFO7cQppcIEqm8qR0ywHLJ7HbLFWWps36GetzyakroGtlhBeW/cd3fKGMb/
J3Xdx7mis+pW2YHx9JD0zMA8RQ18zRCGOv6f1lT7zLsvtYyuKqx4pXfXeOI91RGZ
pMuK4z3RofzdgvLuLOpuPN6SWIFDaabUBpjkbJmrzQkdTs8Q10H22Zndi2vquHag
uq4+acyHs2Vfyst+VFCDIy6ERcUtXRZ+WtZwBNIsACQ5ekAOmbD2jd8VX+HsTVgE
qfBRiQd8P1y8x8poF+V8j0VsA4ZC9BtLv990UjgvJfnn5ad8RIUVG0Gie6YW3LHc
ASsYvC6Oac3st8PDCDULBoDPOiKoy8E5ZYxkO4hYZy3nP5/uhTqjSbxEtJV8qjPS
dEnkNyafVqrcWg+LfOnafsZNNzf1oGryGZyNh9m5LsSWDWD6TDxonYoV6jXgE6PX
DfI+D+l7f/LqqjloLm+2XhS+thRB8rZdam4DT8cNbUZxIHrZsFRobb0LaDODcvX1
jmHq/E1bgCVa99xBpAuWLt/AgYBHC3pHK7b/fW7lSw1tDACQc5bDRNmpvnxA23hj
YxAyT5cMXfGqZT08DaSVzerDQ2X3x2/MioymyZ6sYZajV8kdfTGBDZn+W3WQOIMW
YifNFN8+hgS3TfH+SBYDRPgKvvL92hjeNliAYu7/Nf6MSkiY7OMM6nSdWMw0JoAI
w9V9eCEfAzJtlv+ci/SxWDSoPjz3zmXItaZhgLj0jHZaG+UR0HgrCy9YJPu5u2eD
+j3cclsL1dRBVXYIHM7OFurbc7uTr4W5Q6zATGTI3OJl3I2Z0jKyZEC7pWG928H4
vSx3NeU06nseqDaFbzIgVXt+G0A9ZwbR/yJJwLqNmZ1Xsq/uyi3ZHUAbvHICAnvc
P+h7WSGPWu9CeyaGNNwk3jj4sHti9Zd8AMRku0cGd+SgoMwJsPY3xjhQPSL0NfpT
8o8KWCezqyJBT5jFCvTGY6YdFYfnLly2AdkjSB/d7Gsy7pXwFMOku+b3HKHMz30x
YPiWyoxsytmSzqL9jTb41s4+Jg817EerIzQETDDzjP4C4SmqfxC6Mr35XXNSznOz
ZxaqrDJW9Ij/UnJDI8TRE8118xK+sx5O6tfvxNsl+TWFH+7YltCqf3uw1wdoMgcs
nhYCvgibLV66/j5N5R1ErSGCMJyWzCcOmcWMU8Qzw6WJwsNKDn9xql67YsHMs3i8
qYj7x91J0MGVXYaUYPN0CU38uWnqzLfzVPezu0BiSCZlrUhevGak8RmBYKXlc07t
uSKw8NE8xomJoKJL6uSSi/VHfL7M2YaITemSo50AL638PoB2lW5MmUtKZJBEqLNs
pfDxQvemXaPjyHq3ncV5karsSY2w5ResHmK0WVO6kW/VEKAmExVyxvN9N4e+7MvD
fmtPWAM3qOA7AbDwQECPKWdAlJZWhy0wlxdwLkK0XFcZBhO/RsH5Tm1fc3Ao1TBQ
9M0/67gKmn0rErx2Uq+Mcxwcoasdb+/ZOQ0XpnZTrrY7pXGWwr9skqIBQPgTX47T
zfAZjhM9PYS9xcwp6E8+r08kbqN80SXpYI1lLScQDJp0XFDlKAhUsIGSJfApNU7w
BGtEqTNp4u0X1NDgfuceit2OfCykSDxXBmXCOg7yG3V3hK1rSeg9nHsxlRJjgVCm
J/L9NOE7UX6pgQ0156IJTLDTDFKHHIb68RqIF3p+27SMLWkG719TbibP+Zlq1V7V
BSZ9lI4ELvXOoSuHkxiLhkBm7U2P1IgvkaHcOkf//cs4BzYwYudqcsXynWH3bQG0
ByvgPvmgP9lC7wSDQV39WKuiWMABx+wnTlNVWx3H3AMlTSK27V7lUv3ECOd2kx1z
zxhg+tlJYXtUFpjzARbsaAOSgpBBDisC8lmbJw02kM9KizsPlinLhVXdzylaXYYM
RDfRVoB18H0I0wzVTvA4YKV9rw6eXgJw9RgUdvwxqJMJCwG1omZrwkpINYws8YVO
FwtJJyBW/gFV3DOeDkNAnEJ+lBtRtT1ycOEm+Lftd8ykfub9jKg3QF5EFes3YQsd
Gy+hze17q2ZXCvk4z/lVGWPplGwAC9S3f9otSC3vEeYMO5BzpNcBja9lifhSg38X
cVTS++2rfp/eO/uIzYq9en5JIflVlE/Yypvr46QOpzFVaCc0poEZVsnrMv1B+w4N
SsyWxFAz9DAe+l3MOtZRricK1mDkf66KNDvBA37gW6t0h/VGhfjp/IivlytoVqX1
3tyJiEUAt8TY7sR1ffhp97Z1z50ziMflggQdpgzKVAB6Ou4vhwP352wmbetNeaPt
tHvTwMOa60EyWwxRZOJes+SaMDCuZn+2XgcbXHt3jEP/OTJYgnUJZl930gCF1mGv
Tibj1smpMaEZh7DSKv6LUupU5a+oMne6YweIboLpyHfjRV36Hc/PlnoJHF1g6FHt
zQvPX+wBkRHdwd/cEp3jUGwB+g+0hGJOHRdiLzTSVNFCeEDemXnJ4Rwsj0op+npj
P9CP1cdB6q5aI9A3IHYwARIWiLXvUolrds2XAUIegXuaa4IGYb2KUQgQVRxJlDtJ
pEAUCP7RLhKAiZh03AKtc6dJevSOrta8nat2rxEYT/BdYnoKc5D3s4RUPp00GTpS
LvXSFTuD+dZh8a5wEw+40Apkdko5Hc+vnBFYTOaQwRm0cbzf5plVOaHd7njgUkjW
ZRd0vfgdtvXbfKG7VpJgLxnqZ/xyc+1iY9v4q3yYh0743Es5PABCxnuHICWXX7+8
DQxNGENYoocsKdbwYy/1KEh59y5rp9aC/9K43mOmC85CiHLStwhcPRiLg7y8g2J0
xRvC3MUGsmB5QJXHk80npBXfO6uPSjbkSs0FVyUC57d/zrNqIyBDl85zh9mDKs7Z
AoJX+2ocZ3GFH2c/dw/etMuolkzGItMNYHIQndKC1EAQZt99UmPKvSpydbgBFWgj
g2dW4wMUcqeyq08vnpsyUpwmogoPh4E0mJuwJn+ccr8a1wDaad8QYe1Lb0UhsBgs
BS/rNONXdPW8OPekcNJQpLAUMOSL+RZvPNPZ00m6poUxeI0+CoPUOfIukUOUgchc
ZHFObeGMRomMjV8nAeDtiXmmoI/bBIlDywQQhoOeR8FLwkvr0OvVfIgW8NvIoqwM
TO5wfBLMVJ/y4XMHjBiq8YapSdVu3FBxlvpcSahrDYs5OoGMTgT6kQ5/ScUOfxiM
7zVBBCtVbmCz4uh0BxDy5GAJRYgmuH/M8Tu7WQLBjvjatUsBRNz2dJixy934rpN2
gag+QDvGQ4expYpBSkMvrH1Wz3m+6JZiY94zcTeNt/J0lQOhV8DIUNXlPJuYIscu
On2whDqcKV55CrlgDgf0y0h+bXHuB7canejyq/c+Cv10tHF7yRLDisANtELkt63g
i8s8drajfMhHeWxLS9BWD+kq//jaKWjfp5DLvdwQZ/6jzaX7M+1t6/1OirDZHrpr
DlIbGcrrkG3BfIwA0VYJv6Nsoiv8iGtgqXJK7KMimGDlvMnWAbRZWo0sR19dh+Tm
l8JNZvnZ9lQL16F7LoSQRQan2eEAw59fQs3ZpHGyJPSO2+tct65nGheDVnhgbvPM
nH3TFShZHitgJA34uU/RrRQ/R0b1oD49IHL/19yQrSlSDeyeu9lS/8zAcvnE93Ae
bpx8TCSxjdiIcqKGgVMIuy9787QgcRvgwA5JpRgLNYuCq+Bc2367ar08tS95aXbi
JKl2+PSyRYvDLkV7RSwrl4LsTmGVMT6CQVGmfxMd6+4FMPmr/ArEEVcAbZbzqySB
XTLVxdUGnpxmVooCv+iR1Cryvm1KOby5NYLw+Ey8HN4nY2zjlHGFb1/NR1Z/Hc91
kRDcQtQmvz1Wf6df7EN5FQmOBL0W0hEr5QfrS9mKe3HdZ6kY0tW5J3f33puYVjcZ
DARmY58iaWRRexAyNW+ZhNtBQZWllpRarFTTUfI/WgzSKZSuAad8tZT217YGv/RL
3hbyqSprBgJI7whKIPUEGBkluo8b0WA49dR8B76RoX8Y8zfgPpf6UTU0/PLsQsFM
SFvETiCVSFzj36Yg4C8CQrUxvw+y/9FgmjBeT6OXMTGFmh8bzExItUqVuIN5JPRN
W09YPRmVI+3mGTOVOGZaIS0XcK6WhabpyP4J0SPdUtBUla2PCQIkuy8qT6HShFM5
ST+Rl+0YOFxMedNNghCh/OI7fTkJ71jchTMKG0e5nb+5CNOorP+gGg+X3nxQ/Kcd
ykk1J/HSgiiJolA90TcXVnhGrqvnLzAZYPmGTVjXQfOwvrW+r/emktpWjY+K9Bc7
Dlw9M3W7xtoC/Knn7Xd7x9ztzdJY8cBopjdwROcwdfwWQz5xv/j/Lp+qKEP1y1pW
kbgjOn+Qg8ef5Hf5TrZpmdLu4/S+5Ar6pBh0+YIISMl/b5CGesgblZsB4ZnXO3xc
UScwPtjgy1LvQfYL+luTLtetijpSKbMIgS6med1OOu4sOdvX9XkW766rCMUtdcGi
UuMIpQ5ybfSy94cHGvK09HEAI60zRXkG+4ClOdZ02qkqZQ4UarywTJ4fsjaJhkNA
OFNRgiC6caBHrp1b2QGWZofPNQlZPrgBlfmxKclxJ3DKHGE2STx26fZ63Lh5dqJ+
5TpPh+Jm6Ffp1Wk28qLof6cNruBRJFtI3KCtC18PAY2qxFiIB+79I5zTTZEBFuBO
MMCyqHMDCD/dnA8zH9mEOYPX9sCuwLSoF826YQK7xMxpwe6wRNGQL3HKOZ1yG25Q
5nHJxr3X//9szCY95mgFKyWG1H23uVJ7r513Q7tjyG6j7TvI1/wcg4c9vcRaLnI3
b35rwE3aAELenlchELAyx5lj7ZRK+KFWY87zjotjgiY3p6uP1/D5ZHYM1UlztcGs
/nKbn1upDDgiWgA/vEbpQhaSgeyOIbxHgjV3THpzg+9RCVroVYHFBWugPmqVcQja
A8xwQ+OMdjvmWc/lM/PV3EPkQxaVmlVsi0mOCxbVHz0BIWaTKdOT69JrENVmOIsz
+Nn5OfVT5Y/0IrFVn8xemCWN2ciR1CzeYtV3B5gsXwIrZKso8h1lqU7Gy9bldmdG
FTPFuH1P7o35rOBT4gnsLcG4ssSjSZLb3TstFfiZ2xGqtZFmEzgjdEakw0pxu/td
r0fCkh8mBCk3qoL5XA+yrf6N4QPdBauCL5kNJ8vhHq0O0xbxEYpE7tsSb6kbROuW
+wX7PgMx6t4VsnG6pV3gvpTKmnfcOZO/Fw2kN1WgdeKHyqnwKYrMt5aOf028RM4B
eLRyjxwpgg0JGZueIAmcKTS/p3nIJVyI99G0DGP/x64MEZ3SkKIr1HKMoudevlE5
TuGoaRG4JSKipiv/RjtQ1Cfs7UUNqpY69xjOlKMNz6ZIFwN3ZZ3g5vptlGMxqjBQ
DluhDXU372G3zYK/dqKZ4f6P9MUaPsHs4Tb41fIh4ShrhgJdISZ3dRc3gDvLdeFQ
6hyqr/ZXwWURBf8vNfud6rdgUdn0p5ZMf7irlem7NST/tzBjtCZ01uWdEG6ZbTV2
5EjnmY7CyEgVZua+uZH/tcM8nsPDYSDb9vayvndPkkL5TQW04xAp/q3FReT40gQd
aujx3bIBR4D0gCHSP3MWlJ0zfSxNGnFXpKRAGXF54sgQW6NFV4y0iVpcCElKgZu/
4LpdwK1TiUVgOaA7WoEFX+yA7OcXcUfo4pjSd5Ikpjz58sdGUnqHALHAOPWR/uU3
12zlaoGJLaCkOfsmPctlwa2Ok+nU1ko+hQSTTH+FwgeilNiOnL0j0vMovi4M0Pks
38juxScL4HCZdKML8YUm+irmxugC9lho+Tm+WcxiwVyWhZIo0ts4SLTxgzWPj+iB
Ocw9B+gDQP4LL+T7wHIjnV5N0aQqtYBZmZvS2AZAKO+TFWduSxPd0sfqkvZXoP8t
zjCU24GFJ7ZKSoI/iKD9VSOBZ+NEcAK08hpEav3bOjRXR8+c4lAemX8w+25w20eS
gcnaYFnvazQf+gDcNx4MG+Tks8aGTBW+aSRb4HH8m6AcS8cTcoKBzDa5p36TFEZr
q/YWn82hy2IYy/Ib2sioIlbb7jXrQw6O4lj0p3uIC/hdlegDwJ6mAWY1+DZX88eM
z8Qpd3pjmin9jAbJY7CobOEg2amtZisZPX3y35k9lqQ2EAU2j6EZ+zeNlrJfrnH9
S38rwf9dvn0eGavKISqIEk/8/KYe5+0/MXVseEOST/yG7tbi9T07MtqeutYURnmT
aMvFutHaTpxgUPKp9CvYPyURMlL/gHpZdwqvqTc0jkr1VdmhNNlQ7m89CjqkU+fL
RCg0E6PSDGYKqZXNiH710BmQbfk5K/8fC3wHVMg6HrhpmA6cm9aF3LTHbluFm8Um
2jpVlnx2y64hzfxBTmoySRMJaNuXsNDpTFnFLS2JWWrQK2itKvcWpPWwvtuddC+R
8J1/hiFHMLrBpLoZKydGgk/cftDvA0b2uZ/eLqoyxHPHyoqmUntmq6y5k5CNkc7M
nG4gS7wRZVsrFbmAOSW2rJcauMkCHTpKGdNlrWrfPSKQk8qGr1D/KueqaoykJ4u7
7NbZJf+BPaEzUxw0rECsUjq4ts1r9F1rDOs09QdTEIjCJchFuQdP2XGNy3TsLqVJ
abZLs1WFb0KGtjO0xlCh7FpsN7bcuk03LqV5iBnIVQnRFGvbbLw/rfqDFgGkpAlu
1RwYWr1kgqvu9Xvop/97+Rwi2HBTOBETzFyAPf2JcEnan1NOW4bkx8psDOkfoPJ9
BMVHpGygylrXDGTHofpHK1mKFPpt7klShFgvW0W1gWPdvGqTi4Et+8aLlo9yyHwi
iBo6IklM8TcWqWiGJ9Upt0pLnqeAbrv+zPSF+tVmuAPexWm9HIZ3sEt/kMJsCEaJ
vucHUR3D4BFXiCk9PymcwyatiZCBor0jVa7hYzEJnXaN8XEFEnUsFr1+lXCdkqPM
nmwydDXxmnB8x3VxFyd3g2uUEXSeaQHQ6OD/n1o1D5FeYbI5U4ZWwNgr5qNn1gWy
WhLdORynJallU8bflSVyrn7YM9F/yomAo9g2R13BFPP2PTRpfj/WVKXcimMfe+NO
vd66pCwBXqIrAM98i4oIBDkz2+vSt2A7B/M6BVxJyUlOv04DPStLevyiPoYUj0X0
5eh1WNZ2oTKX1+GvphS3DEKUFE1xHELzIfgckFEdiSk7+uWwFJlOzGpHDgPtqJXw
pzDOVhKDeuJ3N1zVueRH35x5FPU/Ndu+3RlaiI89wW1GdkQxbDrsZF/noPhVYr4+
49Lpu9O/TsLwmtJV0qRgmUmD0ffdHipht50fVHiaJ/D/ffR8lLsOOtZk8fqnVYg2
ArCFlB+SFzHRD7IB8Ihu5yzhDG5/yMsFvoQHCWSLDazDfX3gUYoPpKYe814JwPRg
TEYkhsVwqSCkhezRSmLIwaSfWo9+bETC2f2tyo6iLgRSqu4PDUiKh3xIk9+BkXvA
42susvcPoGRYXX/NeOXl/aMvwNYm1NNLakNbtE3KwMgmn7m79eyg9Sug4V0Uc//1
8T0lTQv6T6zLw8IFxNx5RKZ/DxcSbMAfNEaIPzGWosqAgBSaFDs6k1TGHbos4seW
x2C8KmVqnTNKOOiGs9p3COy3ChurU5NW/aYIsDMUhzXe6wx6GhukRgsvF7M4O7jw
2HofwKG1rguRUwF/exvpZcIvsKffuBTpe/6j14I00A5oTADbXXE3gBIvuXDjWtuF
vaE7H6VwTB5xZgkGSlZJ/GaB3AiN+QSgbVisUTPhTjzFT+xPgKXJM3ijHV9VdHPe
pJajvoEFIfM8j4B78HP3xFcOdmcRQTeSNrm9L5EzqbjkvMuh1JHvRUNlxbKlPHmV
PW4jPFQNQrgqUpSOShYY6hOfLGHWaKkvJBrmb7vV/WMlAHMYQf8+8XglS5MhIoXg
mZrundSWy23Hb4so05oW73PXkCp8eu6o1bEVSZkwM9nLUlN8O8EJHLrEZuwyZqht
hk3gV6JOij9xp8XFobP3y3i6j+NqhZSbFHBW5kw8xbYwB36JV4fpH+9+VOzqsGTg
D4VPUveWnprPrsk3us3zepT/KXkj7cKBbZHRZXnaacmoQkxUKakLA+6fSH5wulpO
sq4J4gm1rb17BYbSwfskDYWu+4v4w7wKB6Ls8VXOoR3ONC9pw+HsV6z6pVFQ7ATA
Q6PfbB43OpKllFBr6O2KxrMtpMQ6ZOYWHmU1D6+mMOKdzflZ8Uvagss+LaS/at1f
dxKsX2FTPC52VLhW8RHpwYNaqTyjlM3hUmhxVLw6g8tCHKa1Gfj+sTMNaFhnlQTl
Bh1VFOIJd86U7LOLTG2qbKXxAkhHeuSfMYCF8xpcOs3EBsKbbUkODmilBZ9qlzOM
BwJl6laDeGT3T2EQPVi2XOb2TeHsq5PMS6TJEqvw6emL5RWQ+UBrLtzVg0UCnT7r
8imMAaBbICb7vPBPwoH47eh72TSCeauyDysKl7uJxjUOrDQ5n+zVv5Bxjh6l5G8/
zgxFKrIy4TjgZFeoy6dsIBf/lby7+1auZuJtSZVMTn9QMYeDk4gGllKT+/YBFjEh
ta9qolK2Md4kdDpR9AyJPztohZsvakG5pie6QGJXZKI7B+EjWJrjmyNk2xVO2oFq
VTyTxEpRVv0eWpizgfj8KWbbgK73iWld16/Vkd2KfRgNFVjn4laO+DYZHNGLexvl
0JNIA30y+cdulwiJe187JP24Oqnr2LvLQx9aRDML4u72Xs2lP+0+ae1HGSn29oHR
RHed0rgDZ8arArRpXq4VzVWJeyBlesj1Hl6tIEU0U427qx6de3CkJt71uZO0Syo4
2noY9Sgqo/JcTq3khQpBcikLthCu1QdcX60dtkSVjEG7A9ITWUiC9sP2GxrbRivF
cVHhmcexOcMp7odm1wnwLi1+Zd3eCXisBarCeE74R1SIvPer95nDWip+i8z5j+yf
1XIIDOUXDpNa0hM0DA13bh/GFG8LK4TsLThXy2oIe/3WfUqtBDAz+z49V+xGbfTE
LeEHjDA4MZYvIXf0kJSgVS5lh6n3E09t+c/LGuUZqzm1vZU0Ru9IQRv+7a35VTeG
5HMOOCSEg/3x+d+O9l340IRoJsamyAF5MMyx0YpdGg1zHX8J3APlqzGhHk6Ujtvy
MzUDo4TVLxkBW+gYpclvMcutqlQRFTNpS27UNpoMe7XH3zfh/oZVBZDeTncSYzUN
MTYhDK6nKb1bjBpodj2tYBMzStP4YEoszwI/kASq2UTsTHZjLAYjhHUvSBQUUwJR
ntRhcTwQt3Bd8Cy3LSsvVqzzeHrhu3Ii/0fzdabpX/XKF+nW/O0vtWuH+rz/mZGB
5qjzQs6C4VJ/EBurSIrczZ07T70fyzLHkT+iL6h3tUCsOo2stSDjD3t6dfYa+ej/
RRAeR7woVoc9b9i8DrkMbSFKWklIHB95O6TDO+BjUOBxtDP5MqRpMIIizQl9mvK+
86Iuf+GvAxQgXJ2ZgqauZnx11XS/x+bRwGoIUsgeptQ8JfiZMVQWacbimCkQZjc8
1Oyi/lpEPZrahSmFF8XITiWBdz/1/VCee5kJ1yygiWOYyRTHDvGpfOpjaILcfWrS
fMcXQZhZ3rt9eTH259dGyb+z8r4iCqY05ZHJitpQ5HHY0yaJ6mWLeqp8XuITAwlH
az1Crg9Ixp2Z17EI2AUdPtq1+/MxydYnlzgsz48WluRd/cizLLor/UeVKMVe58UT
7/fra1nTGnPgtuZxSl/rFNPc+kyiDHJDNJ6x8x7RvriokSCQn8rtO+dyAPaYS4z0
5JiWd4QrQjcDdYKCOb3I9eCXx1XSs13ouqq/eAGhGZ8vdeKSFD0upv5oOP+v5XjN
Ead1PzWgdpSCpeSfozExTO3xXjBAECInJmoxfP6ZbvzQSTrvkHVmYtcCiOv6K+Em
IIzfE/8PpMTYU/cwDCNPUf5Y91UwoUg4P0XVLYa5mi7fzWwQE3q0dBL3w82ike7W
hOo1aXBo1lxdF9esufGBMXnSA8NzAaQY/clFxBsRs/ySIi4JvpBR4eqCAD94yo1K
rdKZfgJwaEaS+/JiL9rho/zzz12V1mNYSibal4BmObQ0ntbgEoYkDvwPlY6HBuXz
3uu0ArQ3Ux7kWdtsNI/+uMrqE1LTNvzbOQs9IfdXAeEQBM21laf6q/idK2U44Szz
Jwpo5+kUg3Hsgpku6R0TvuwQ99SgnyAOl6xaj7dzoe6OMu5REbHafucCxBU+DlDx
z6l3mD8Ll0i8f1w5hFQjqJ9Iif2nfo5eYXIh8O1w3wbsp1uuCbVHj/EKMoxDcu8G
+BcDjcH/itN6S++Bv+k68w97FtJ4nvHt5dYBjzNZ5ZcEE148CSgrp2goG/9mZUca
09PZRb1rUpPDH9D8RKv+7WF4PHkj8QM7SOGfB94arSg3ZVW5WeUWqTKodf0Wiex5
7P6U6G1P2njo807j5+X6lWBiTwRC3pT2hFfeYfLCQ/fFTHdAgTeep8CP3xFBC51m
SxQOKokrE76/tw8ysIJuDb0L6RR+36FQUbYxqpfkdfcyMk8I4p8oSvE6gjeJi5aH
4y3oO+b2p+AKk1S192yrjo0U+mD56G8C1oziuwMbibaVpoagm5Yv/2cQX4x7IFFf
RfWybR4/R5JwQmX0JFCAnIubs4lhGJ/6fZDQRjwwyv6imdmUWX2h7GIwSrN1CxnQ
hI+RJiADUIvqia82aGX0Q95E358iRYi1SeD6bAvatL6uVeiyxF6FxB7aHhLjCF2B
x6sGvSlWbtL0CgBICS7b6F85zMHkHwUf2BJ+nBlEE+8PwCvTt2IN1sqAEH+m6xhj
o9QJrZEW2eHiWKArYx0MjUeCURCHnpokUTtKFv6bKb8vzfXv05KXm33o4iz0YnJ8
ZxDbFA1/khYJVzcJ3lbNtV+233QP4UPW5EDgYN5ao5o9XfvSdeDbAFRJHa3unTbQ
06FmImElI127MVn47834Gz7dmsxj90laiPfOPUqFmcgybI435h8fnr6fL4n6sa5/
82WRXPSiP7IGOZIbphyToeXnsy5kmFLPPEZ+XCIegAv+q6HLkhBbzVRgiy9IKPba
HY6ukzpXMHZN6A1JBX0d1PbebW0Yf7Odln10JqlV0Bg4hliGcxZPhDAa4WDsl0/d
oYIfawNVG8V4f2km7HIkR1gQZkXWkHNGJiVXGyIROUHkf26cLIdRnr46cSKWR8e/
oRKa4UY+rJC3WPwbsw3Okoh9v3kDv7nPYjW4jK4qJtwTKCzvk/2TZIK0jYZqcp7w
f5MX8aGRqNbTLs4ZTQPHNiKtDpmr7Y6ntl0tFPAIRlUcfpDUDXPo7uohkMUYBXi3
n71LomPushVN0tRRl0Xo5nhI8AhgfRTZv0zocILbXJhC3ubnsCKlR7xrWDIlXMRt
Yhm80UXWvoC1udLkWcAAg0B1WQwSurUerx5cOurDr0B4EvdIcvZPyvQkqRSHL6kW
Cl1YttO+Aew99aeTr1wx9yrcUSMKCi/Oo6kuR/EGuggv4DDp6vMbGFa2IVEdO+OI
2WZTGDUdVEue4ltc7/5oq2ipb1oGVCv8QuMlLkyRocq6eF54NhNoV32NxMWOUwpF
OfFcVKamFvKBpX+Y9hYvw+ND3Bozqepki7AeDtYp6GzdkY1oLPswo8XNtcBgIla4
NDKRrOZlStX+twTxzdnUIPs605ktE8jiBhqakLUEs/sbAfG9ddR8bD3lJy/uVToE
t7AORF2GFGxKWNURXEYcrhOmBlS0z/TEsaYwzScW0g2agxcRF9WvowTisxwWWzw1
d3PQGSLJ+NjNFqvc1bJocBYVIklRnvpEG6WWZCDmWoGlUg+pDVEa9ZFIQm3jDsET
/6bUAMzp1fEvsmSL6fh6hE40IehUoK09VPYVBrKTypKmVveK+HQ3NAGywKL0g2lu
jk3uQyTQmxsEwe9XJekQqglvOi6bxhs9Sa7Kgdz04Zxu6Mg6WBVi+a+NZgfgsdZs
ePNJVQwOQXssGdESBb7OwoJ0Dh4n8QGnDe7xxCpaSf+3x6hKve796Xy+B5TQZPRc
VLPAPswiDjmtYEQ6kAqSoTLEtZ1c45/HihW6vrJ+qsn4DmHg6HBwYshDNDBXQNPf
8/J2vtm/wLadN1+y7dtBGdwXyGe3Vb4qF7Gq4syY1S4S5XZAgvukZwcoMBIcBMLH
0aTSzuXCxEeZ5a/dlIWWlyMo4RfumrxNvOKew7T6763tfa0Vt4gOydcMNZX8s6gh
rOJ1ev9SIeDdJUzVYLlxI2M83WQk0s/NxM0uvfDnDyDmT+Wr0PMR+oMR8CtTb17m
zziL77LiHfF2TlISltkosOF3RUCxvcgQ2EfBYey9GzrbDBh1UTdd3UiqQoYcqXuw
QBLnBBTtYvZJq/GyY8IhfwiqJ1EwXlcGeDwohnA1xHvrLqFHtstKUoN9ke2mHiJY
CcjvcJCvY8OpEbswA+lMCnsrIJd4pslcr2FzHomZWgoR/mQPZ8PbHT25OoklvxMk
8GlZhpv4KFDRKFlLoxjC5lhWokcXfdBXF4TIyLhhLt/9rNLDfVV5016Z2UlPYtm6
niZ//MKFXf0chdKh3tOh7H/bdJgzsiVI6poUcDNk3/lF/AIV/ZGHE/L404qH9prQ
JkmkB7C/kwJzW3LXVO7bhltLwmtV9nwA6XJlGLcv3AJdzpPk0m28lGRGkV0TyIEv
1zGVeX4UapxP+aIaHM1yxlTYJU4QC3mKLrLzL8vHfFOBpj/X6aa9IUhVACyPOnjL
aR7bnr/Lab/yGQXbd/iPbDpfjfCDR5H3vQw4iq618uPDxWd3WKdqS+G0jc293rL7
WCBt5LO0nhbyW+hc+XsmYxS0QlIr4KblqO7WWVR/MftAHzJj2NP4M/QotF3/PJ8d
RVtSQEvkokOs53UzPaDzbAPo5lRfV8E3RCbQ9L+15FYeNCJPHMNs4BEgYFPJ+ODd
ifSQWlfJ3foIkQbggFzxJiZjNSfNOMsTA9RuR8c+WJ7kwpkkml1uUH410UiYBzH7
pxXU5/5p0uqOAZSoE+cDKry7SdXOyVEsvskvh46dtrVybG6Jj/TLbcFuuj4EGqVG
v0in7E2QceEkmAQxhmcoOX5rxW0hGFSoE9w1o+gWoccsM275QlJBS5NorMqWixpD
4M2cpyLb5kR7/gA5hOiJRp+DoVRsNxxxQoc/2qPs/u/WKCrfRBBRolN+LpMoJAjl
0zphfYJSNHTJzFkWcU9RvXTKyi9ciOQBoPcn2sDVGXcGc9iRjeIMn+hxixoveZEO
k33gTsAb/fwg/dG2W6WJHyIsemvcInCpqKLSK/FOHGsYvaoZGxfjTeOfjArlbvQT
MeqpaPAhTeWDvu3funpEJQR6V2tIcWVnwG5WOtLNmDAV4GdZQ9PrFAJbXuVcRcML
YSo9prZUcMAQ6mdZUiYrinJgEisEO0TZuPkV+1CoR724ewMNruTzSYsVU8nw8suj
bT6UZ/97ikFuq3gYDBV1lU8wH36Q9X+vrKljikayALA9c2FcEs4NyKADvUk5NcvZ
bYmX/oAbvGVO34olDmnjn2aROkcoZzVrQBrai9zH8lsw4tlVEms1uD07FDjEJpLT
hxda+mCiboCNB5IkwfrhwL++Y0wp+NL3+cn1xHkdPMZNtn0Qhwmhx71PX+NpZvA9
vnM/qeCtaJvy9Vzb1fidDUi0DntJh+m5oTpo54zu9ZwsFwSWvtgC+IZOa6jwVc0a
ksGq0LAyHknBWg9fDk+qlHXT4xJ2l+ly2+h0KhuTjsEHQgLjAJUh2ikPBFRirnSZ
5nV3bkMxA++FA2wUjH+cl+rarL2hq+6KggAozSTImgOX0fl+qXGAAL8MSWzMNxhM
xupRAticcnq5JKispbEAmFUqb4xeZNm/8yfdX9RV3X+RrEurt/26d1w9yqee2xQs
G1A1uCVRINk6G+KEynatsYsBU8o1OSJ0px0OVwKh0f2CzuLV91NzOLhWur04nVAK
3VAdT5jzmP2PxkAPOrA0/zy2IoAb+heKafeddz7KqTadruJLIk8qmwRUJmHK+0An
5YCWSlAWpmEqqjlTA824nx/Q/ZKScbN6zFvh+6yVnLtBno1DAA4W+1B+Jq4b5Lw1
D6wk/rZkwYZjNzQ6HoX4lxeX8zG+QDx2qu6/8E/1NFjYcXurPIKHYDH91l4Z3bO+
OLI5RJQOET94Y0a00SQUjSKUHZ1vk4lm0OKiLyFpNfaoxtV1T1pDTs4T9/k46wVS
qF1ZX1VJab2tr4txl/oB2wCBfvbPpL2rUAzoy5f8cHPf3pcJPd5EO9qVKo3fXccT
eloux23fy2pvag73xmwSAy3M61plylcoFkZ6LoChYM1XgHvZf22DFqE3utFk+BsR
D61IwXTWlK8c8iQXAtbQh+8I6Ac2gPwCCZjR1dFghekwnYXtPtHewQeQvEUrNSbY
jkLJnU3RCtGa1wNcO8jZ03+CQIFr3dR/B2lcvOd449ub3iBqY+3O5mniRvibXLHH
dbx1LRKsW9MBVWu+QM2QXfpGn7DW9BmY6gZUBT0JuB5sQ4LC/YSnCYEJXUGpJkgf
u4tL8O7V1542WI5vBwO6/g/rPabL0zXFqM43T0QBtqcvLWn6kTJuWzHOUiDNerL0
qCK4aaDAmKa3FxOkTduS55YXKCH+MDfbJSphm4JnEY9vBWJaNYOphRyXTRWMfybR
ELqAvZ4B8XDfe9TZ9TQrKrjgp60K0ycolFvw9Acj9SERRP2nvsp8bOFBqvRJ7TbW
7F5UrmrjHqJxDk9ryTCIsXj1+QBN07RaYgJKJL1s802VEdkqrqh33Gd9hbKcYdVa
yT2TnK+nFpU/cHqnaMxXf7EP0QM9lhVTsBhLiIuPWHOwNrkp1vZcy9MPOq97JAzk
NWw6+CxAOVqFCuo+qdSNLoZ/JyTIczhDyJbnq06TWMMEYAlxx+IxfyvITn59BJ0E
VB0d/hwuiMZy2r9GP4BGQbmHerR0RDcV2LWpngbsnVlPzrfhwL+YJPUWMYQT9h/V
oyUa4tId1+DxauG6hDpo/rmclPdgzSaQGW/tKpAG02yZ3b+sS6dQ9J/MoOA9sdsY
ICcMLNsUXrKUbGEYepYHWkWW330aF3PhwS43wzfAgNLG4aSEbi6jEmogtiavdK0q
JHz9JwfsifEHhqHwta2I7IBXke0vNmsP3ZXCIoE8zM70hSaWs2/0uSacOKB4D89T
eqQF5XmyrvF9s9V++fECvi4JlfbLz0JwyBq5egwp/gT+diJbmn4tl50yR76S2lnN
V9ZrY/QgbbcBGA0EJeHUBB1iqaHIsZHSxCASQx8Ltk24pqHUWUsqOjUh1dy+nLLw
/BtgxK0k41lggWaC1auRKgggsPA5TqBVOcBVP03bEgA2Mt597y8LTQddc64Tch8X
14oMxvOTUL7Z415+ggcvSItYMEa62tQr04sYRHf3EHbQ166wGulCvznUXUATlYxR
U8RKGnFeSJZFYAGuUx5hUgiEb5MA/bbAhvEfb7pc7yWc/srkcBZhq7wLJFAJVA7j
MkoXKu8PP9B8GcwRxw0VpZt0BnkGdsK9xKNOnV9yrF60hYEDlcIFBtZFnUNtL5wx
CgnkcNZSfFukHrAqnMnvynEg/NZ3zkimS3KFXpjYGVALgVVxT1bYR8rfxSJUJ42j
VJArA3GhtClH3y03VW4NVQF/oUcORhMWRHVF+IHJxvhI2DnjvP4zufhDgBbMiijj
l9atr4pImBGvYy9h2B9UHpvDSXEBZgHfuznS5nJLHDJ52zxlDAU0DZ4M7Ecf9m8x
N1wZAOuZwWFPx3zsTa8vCAkwIkXannithnKIa0dj/hQBPa1kCY6vLx1C+xImj3ns
s/2eHQWg1HAtbkU6Uc6fBLr9r6z8bsGOKTjlXpaVliCE/uC9EBKiOh6unvIMrJrb
cOnDl8Yqazr1EhUCRYVRMeayQ0oj0a5usZB5AqBo+77cR9o7pdT3sqdh4st4hDNn
66AnTtOIB26BizZnHdZzV+A22n5OVa7nahkHcjZSHw0MXtm1XWL5fQLTxbGnz2oB
d7fhuN3c1vI51U+GouZ6KHqXJAgD0D0FfkTMXA0jNzrKKWOU5COYg3BWDWHbEPQ2
fgD+zVBGW3fN3WVoZTlJILsPAbF2bXHWPyWh6vlkUDvARePvTfv+asURFXT/SwnW
sGa1BjWgprZ4mmnmRbOtu0dBf7VNAi8xx8JAQ50h7FJ+Nju9v/ehkshU9u6Tn/Jr
f6VK6WW6g0aXrv5tl460GSrIdyTpHUl9gTgIk1UYdapI4ZK1DliORkc3o4uys9y6
J9K7aLmjeImbFKs5futmLOBPK218x9SHKMsnJaMzjmqcBv0DfHWLuxnm5INs+G4H
5/tpgPUwSjznmK7xC6EV+AVgy2M45w8H36pFf5U4UROXMVANNcM4moIWiRjqAfMc
y+QzoJgnMwxypqk7bWWIUOKiu3iLzs8GCncAKyIfM7Fubh/SXe/O/FAlhLPnlJI1
wIKKhVVMVvbrF5rvkXGaoguUcIWqJnkD4Jv9oZAU92w6lpeAeAxqsZgfA55Fj3EE
8MnsreojhaZpYqugwmKQvaZgDPTUobbA0TBiQKCFYhTQb7ZW73xMqIGVgQKhSjkE
tvGYNEJ9PVq3dxlmObnOEy8MzOlL5X0iQJYVwezSGbDS9I8G4Iwy1th+7VebNj00
LhHSeBhuLMK6e5c8VLMKsHp/PYnvy2g2fnUediF6I76CBTNBcehC8tCkio+lSECj
wKXR0kn3hHkrQ1TeNVQs9W7kLiE+8tQY/usLck+ZKZZh6xVGFIjQgV4I6oDoXWe/
7Lif29VyyWJEApYnQot0j0ZJFmPAr9+pMPQ8Xvk75D8pd/jeUhLPTajCSR2yzT+D
Xwsp5thWMbQGbCyD37njR+7a8hWwk68u4F1Z7yyi4jeBrXkBSqdJ5TC6+CM9JOpy
4dVm1JcfJE9SHAGgIa0YuDzpZ2+HCYdhQq0Nfqayk1M763uWCFGmSQDJ+8dE+9rU
e6g5HovK4M+GFeuSNmAofb0XDwoiyTomtEQq3EVxFdTghtbysTBlmz//vHhICy1L
AS8s5JaHfyNcjsBfMMHHXgPoNfr7+kCwLH9wiTdxYOli8SuU/fjU8j1Dl0TPhEdG
E3telYE4Yab38Y3dyxKdi5WKxVRsAXBEiCaNTIb7AUMk8KOyQJqCwErFUR+7Vws5
+NEI2Fi95D5IFnIsmaguGGGReRi1iBFsGid7ko2e/yU5IMqFKq/rT42up/gU66yy
yyKp78eJxcc/n/+dk5N5SsPH9J2M/1cJTTpB4/YT5kEaMiIK7qRuznAa8dk6mTz3
JnPB7PW0NTYKFywqFs1F/vWsQ4HIpAOjKClmF7vrS17aO2l2AQ4bIfqR3sMY9FxT
Iw9YsuO+aoPQ5G7jlnuJUbYaWp2K+PVU6YnDLR6eEGT7Yd8GqevTdXG6aUv1nDur
GTI4nXRpayAL2VqVzkrzND3GivP3Uy3eRZ/nsklJP+UsGq0qgGPSY9WM1PyVjBn9
82a4IVXdv1pVPB+uXV8Hoz6q519F8/SQZWTY9/Z+zU6ym4OKeXwdxQaKBJkB7N5m
IP0nlDwHUSr1J+sgUPQaa9ZfIWCQOYH2PsiFx31AF/8gJsNn4PzU6wLzSuDy/EKz
3oFYdTJ7ixACQi9gGVYcoF66hykA/Bibk8Au8KQ9Wffv5ZsvC7wlhlnL60ZRO7+9
s7vvW2Y750yRCHwglzDC8YGphuMGr3FlJaeA+bRLYYkJoZIvld7Hw+kOLAIfLQB/
Vr59HGXrGEubPAJWjhMmXA+zLFBi9BPLFDvVzD9XhXOf+PDcPs1mNo+lHEta4YRm
hZ+ETZ2IWpNe1ws7OaPUe0dYkvvLgcQqKvmTULYcJNoHi9LVjaX8rEaEHrO3ZxPe
q8wRHL6DYR8RxoaNyg8owxJ1hrb8IQDcPcojdf4fckzEAk6mNTRjBVmBGzLRer/V
AMF9s33gn6UADD+raCS07nDvQxZqQCCieGheVODO09djNg989fREkWsUQ3TUWlcb
tpFfhzZMHuRFKojH19qsOxMr1GGX/2LDxhQaF/vLtXSKGnz+Yc0bxNamJTbsBO03
Ho2YfAXT02NwO2Vr5cWxNtRfLZMIE9jRIFoDPbDDnUIrefcw4PDdbus5JjbYbLqg
K9zyCmq5Drlu4wnR8o2Mw6QIfe2ALRfu+Wf8yApx/ApJEyISKy1EYUxG/9OMIPiB
vQ52m8VxRuY/9SBLHHvUS11BqgcQ3/zKE/98QZvCtNuumeY9Ruq6lg4quNZr0oRy
pdOT531PA/0j1Zh11NWvuxNpuFXtF+jrzw8RFK0aPbi+3DTBeyJipV3RcTVlSQ5o
42lB0oGF8KPTNBTNMOf0AsAoooCelNJ4xQx0VnnHALcd52dL3sPis5xdfLo3pQYN
9avAttAJJ976rlwI1qruFkg3pvYSmjF3IOFnn5fMmakv2SIpEsLOsuiVAPAb2Uxk
c744PtsFEGwNNgUhqmZkBmhauHhQv2Y7PMDsYCcj8bFe2WIk8bqlRnSoJbMyXzgq
Y0+zzUpNNK54PDWLXvxJSyzKvF+TJaRX8CjAIHflJr9gZMfn1GIepwKKXhMCw93g
Rbg/k9YP10IEN7UlQaoKfcETNr+ibEJDHepcl2QeqNrtT6EFtpB2NkvuL5Uwj4tc
Xya2Hb6dLv7uWNLk9YGlie505/yZga8BRMBw3fNNdGfw5/xizBPSZ3iR4UpglWnW
cH3GQV7AOrBf7ttqOMpBwmvdKQ8ViixzZCGpQMQTvhQq4tnQM8pCvHj9bsG/M6z4
i3fMmWLeLG2MdhsQu3t5Joe3QcCFG6OeOXG0fnIA4pMxuPndT9/orCbjOQrkplA/
iuO0+X2kjedSk+tySzMGztZtSJnRLiOCtIuhinWonlm/yi4szKzXm0k7ctP8/2YB
98OkRQ5wsxLGrLwcvYL+dfFTbWdUs6hwH8qk1voL8UxlnP7a8iHew/6Kx9nhdCjH
mvkG0esNdXxjsQckWlrTPzWoL/KWmHbLdkGdVTpfpku4uF8nD/naHe4jmkIkutV7
Pwfa4ESAyZX6ZeAy2MDkpSiMhaZhcSFjOV6s0Akadew7qn4hH312bzjJZWk+4iw7
PVieuMuJ5icA3AlyO3R7V2AKSUT3921fuaNbIhnuyGzxddwveoWWbZlcTUWnmmoF
DvoUXCfvG6O8k6l+Rqu9UMIYOwSxZRUcx/zVYbarHQtyoe3+yjsPgUoPXAkLUUJf
osP7hhwTwTrNlXDXERxsWVafgevunppy7AJT9C11nBEykGonyPK6b7aAZRnQYF4G
VsyUw2gMu+L+CVIOT73nrbwUMYqZZYtzIQg9DywmdfQQvnj3FTYVHxwqwjP39fw/
7Pjhix3uLIC1MUUG6Imfz72fbPv3hBxz4rqjFWW2wU+9gvyDHT2nB+4nwr777MlX
IBn2TDiJa6dfqcsSTH2DlEKN24mYMIWXg7RO639Gb39MCZY6kHFDKPLAhNhZwoOG
fnrPp1tanogNDTm51CPVobG93RtVfK1u/8cEGwOiuScd7pS+yPsqS5DKrI9on1yf
ZYO1/GH/oirnsQ9DeJKS8rHWK3s4kHIxHFZGs9l+5hFika+PouX4g/kz7pEg7nyt
8y2tbCztmhTVlCV5b/s3zEq0tkQ3Vt4uWwf58r9jSCltDPSTLVeJjtnnx6o9qXb2
FO8xj286m9iET2u3GWSmyI5wvpqyNkoyRDpSvshyYs44E+T1u61PYUsV2rRtENIi
XRrymKshVwVDt8MV0sR6pj0CcsuUiV1dLnObUCXyrOYIhopva0HOsnoO4WFVl88b
n5Peo6X3aQZo9Ojz7eD5tlePrBQONix7N6yMDhvZ9fEmvSViWWpJIw+ZsXfMA0Rh
ULZZWrAQ1dnN0ihiq50d6oMwjX5nPx6CzOG8xVKJCRl5KczWHfr7Mhk8o80DQLKx
xEfjkyE6tBkDyFWBZ3kMggRFjFZuHPoRjJCLA0wjbEUrn2U63Je9ciEfx52Jq3mb
smn+fnvO7WmlLHIub7jBo+5ckBe19JCTf/6ZKv43vxjsyZ5CWP5ul5wXNmE+bXBC
dsK7Iul5DvIdNQl+AU4+KiEc2TNdIG/c2/Saw5ZkLDdxlYk2iqo+37L7YI0mxgwl
kAyMioy3+dnGY/1WirosDngJaAKrurYCOVIW9kXs3io9ku08QHgbfgFKGVh3nqBF
h1LyaZJbtz/RPnMuTghqlxmRig+YefC3ENXt22a4Y6polpyC+tQ04LxAFGX7aLSj
UYp17m0UpcBFSzCPKGDVnFHhziX+H8PHVN9OBNz6zoXfu3aGmTWjIB4jPFBTbRjB
w9Ur9/aN8JQH3J6jEVR9s3oREKGiTQqF2A0ZmUEynpAFoQJpeAnYAT6btItLSfAy
8QVcahZKI8sBOzKn7YeM29D85wifNIed6btZU/Ug07MeN6QeqboysG9PtukBqWWe
HVgsYYprMQkl1UgbpKiB1IXRXF2OBu0+SyMIG6Z0R2+ZfB7dZA32+ND01U1FFMxm
KI8ebdak/RvJnLtDOo4q/LjFkc50QbWCj+au7cLNGgmyRVuyTt28Z/JjL5ZM7sh8
VgYZM2w65Co2r649UXJLK+3TaLfPCxmv/pt3vv7lL8HtFndGvjIzR1MBX9/jVHPr
+dqGRJ+7CU1gyrpo2+QKAer9DfRyTLabingBBpKdCszDOPjHJXOrMAPJ4h38Pv6Y
8BWvN2aFABWhP8cQWMeqkjyA5cexU2Lgg/9TqyYAETNQXOidhUHbvwSBd4OWUarv
vjtHwud6p3zzlyWQY5ths1pDZamltzdvC6rB59hoNmBmPQdmTFuYUE5EpkJoB4y4
KSN8Ji7YIPDEqI3+bgYRxl+fTQtZtUo7oDwsYFEpQd6x3VgAT5utBWH55Uw0mSjm
ZbOBvMzK2fm5ky9X/tNVGPY9t2zHaVIHmjNpBuX7ObjwabnkbYX3WDxVLWpiw7us
OWGBhKLVgoXuzM/qysyZCeJ2Z39P1PMWISbE7h3ilKIUmfIn2nFb74tBzlRkxnXr
8T8J+qbVPMPbdcbr/V8KFcAOEoAJ3uszgVFlCzT+aVCZYJpMm4HTRvmskKVc0Aqk
TJyH4opXmlwPAy5/jZtN2kjjIVx8h9Rk56+R3hb+q8G/OljTACU2Z2+oBhjqhwgk
qS4z67RohZKpcgQnG3PL3+x5hiVKSzjAIA2b99nzjpe+nPV2jdzRXOYhfK6yUrUH
AV4+gnFN8dxgS5GceyfdCFPMpA3y7oI9X/YL0VZH9alXSFFCQvmBrB16ggYdW+sK
KMuFRJDIdl4FicUks7D1URvgeFdLqmtwmIEIF+4QyaFX+Jy+LCs2ZGNPpHB9JLtM
8vbBzLxxK5IKNixt0kFfi9Pa0sNeP4rTFp4XkW4FjqoxovyJIT3Hx8zDwtOQ3aWf
Imt6gow4aoF6ptXYA6b4yQtr0jZkAFsL2bJxWdh3zfm7NH6OcrNV/LfDSenQTTQr
er67vcIhN/MlX5B7aIcuCe5fO8v1C8nI5rRb8w6/BiO8iyl9spqLaMRY4wSguJ7K
edt2ejUDbkmhgnpuXxRcMRlyTy0ySYfEc6Qvp0iV2ngJgUC4f1BPOYvPp9vpneJw
FQZtD/qZ3LVi+9e/epXmU0cVHAEuVgm4I18MAz8WYvc3SCvx3sXWwvEBb9PhX5C2
HHnoDRklMX0sRxj8Q4wLdm3U5AlcKUFWmc0JKvftuWIb/FgbxnbhSbpDzbPS6URP
Ou31NnRqYuf9OBKGdt7j+2mnNTzwJ1ZVDxd3zglLiykO6enu03AibzKX/yFslk8d
3sVl/eJ1U235RBDxy+vdENsWNy3o15PLQeIR+WzbvFLDVyhTKAKMruURlRGu4H7A
3GgUotaTPYW/iUH1HiHlxgxq/0hEeKIihVOkVnsgpd2qSLR7obcdtryVQj4brcg/
wTZJDVToZYDX7Az8PJ2P5QhQa/qHal9N6qBpvigTQ5quZ+fn5B+J1BVN53SU1EN6
pE2NDb1XEFlkl1nL6yNKBAFXhj1MoK3AH4VlwK3UBGXxbece8vSe7bzbVf1Q0K9r
OuLG1Xw7IQ2sf3TJMeP5AHJRjYREtbJN5sO8RyDZ71KFsgp5AtQbFM4jVpvGPusT
v8Obi4IBFNE4PqvwsCn0Ql7bqza2qE56of8N3aLw/x5fffZgpLjKF8WOGjUjfW8E
q79qddaWY2cf5yi/vqHdtginJVh3Bwraawso2MfBjn+zHAtgPJj4frNyux9r9foh
xbtMz5i/Vm499rxL1BEE583bxO+Kh35ifMVu2wm0OwdZoRa0i/upC0db9DimhTPD
H5/G5mSc18D8VRV8pgkT46EKzCj7JvTicm15Zo4lSnWIDr5eKFTeWuHZBsyUkPPr
nHRzLzHGgIkt2N9rLof2zBHTSUD+oPDBlyF6T3+OTDsTd+jrnYZVFfteq1id/CUm
cobWncGhqcWJk4PchJcH3QPA247QUnzVf2dBM0ZJfFfxJZSKCpfrrN0SgdzQZu21
4aeEOITmWFDP0Dw7NUD966PHoWK3a8L6OpnaJelblbLz05q2iqbjrW0Knlcu4VG7
7tFsxN5nqd60VJesBirFCyyx5CFlIwAWnWHT/sFOl0J0woHciUSxUVuZOczqZcTF
Gk5Oc2UY/KGmLtm0XuH1q5zjEufsAs1xf9f82rgKjhzuMynEhRK2Naen9vZfX5p+
G4OD4+v+fnkEyrKRMufqPVR2DUD6wMls8NYYl1wmqxWGxFJusX8OgObUDvCmviaM
g8e0afWOp0Uik5z9HGfmVNDhoFdRqkGW1qFM+nB4+cn7LkzHx4MWeREVKWe7nxSC
8WT91jIb0YvUrQ/TZFkzKDvWOq8kQzgGnapuLjlNyE+Cb08I+0DlYn7WG3+NQMMH
+1iuiipBbz0G3v4n7Uq0G4/ooLKrZ7cm2q3gewnawsp09glj22pNg9W5W4rmD5XT
ON3QOV0dRO8ALecXkhfnbpbKG3S1G/yEA7G310+saJdFOv0Ce81YuFfYN55HImU9
2rQRX4sOG1x7jKyqxvFAL4cT/3MZvFM4p2xFHWSeil6YgTNEVjOT1wDXGtvk+Kbq
d3dGGwLAnAWL2olxxdXGxf28Y4h8Xlw2zoQKGSx6gQQPOFb/gK2KvN+GD/GV8kz/
CDq89gR0AKydtVEUixnjKr4oMN3itL4iX1bnPz2j2o/hDxtag1Titn2mBHT5RHPG
QuJcc5fYbqrEou6g79GaExGB8WsQ8W5hHhG71AiINkNM6M9r+RC8Hvnk3D0wgM9S
AH4Mt0+JcOcWWodYF6h8ut/Ih9OVNHwCmcJqYbHUla+NRT/ckhTJ9Is+0jRGKDms
wVH7N1tFDZHnSBwm7KC+0qj4fqOEoc0BWxRx+fRL4tMyXC7uux5PVKxh7Nd6LD6s
iIZIHl5WNHOSpTMWqixXcRGnvlKtU0YJ2VhlomK0BFOSDL2mL4Df1eWRp00iAF5K
9sDAQpzU8VrK+Lhd9PqJGsxrkVikUsCLTmp8DigufNgJIv+ruclS9bSPKp+U1Xd/
IJQVvN9TrzW4FXUwiTSPG9hGBjCKQUT4uE+tWOt3zgMJnN9UpxPwQaHrA+CCcmrE
v31ormT0Kkh4HvTq1eSJBSWnJaGn07ZcRZyEImYGv71TkK5DfrblE5/rKym2ePx7
ZqyOXOcCie4+fhMsVhPFpIXHMSw+lT77jIt0wg6jj2rT2nmR/n5j5wO61fpMxlWs
MjeMHBtI8uPIs3EhIDlIz/UyC4Zyk/yiP1XPHF6Ar8Q4/GOjgnaAJ5p4t6cOal7J
mF3GnbYnxj2eRJGCrmKzjOZd8qSJqK0T7naFL1PKYHGY9jl/3G/8ULjpqdnXZwKD
NhxpjKEx46Yh8EgoCY2pCY58WdPWWIz6ooGtJLhtZZgQf0DEn3DY/5ZinG7Mw3ti
MiQp+ssmJ9eExKoAY0ps4yWvX6fbPRIHT5J3+mtfSuEBOgPacLLLyf/700ssytmQ
4RllFC+eLJwbvi9VhETMMi+84YKmZW7BA2eEt+jQ47GnmKm6a3mhCCpijC0aWk5Q
E5unmbPShv3FHtweRErQWQU2wUWRjNBHT7Q0ZHNSiS1W2PyJN7GTnjAie9iGoUKJ
BDrQFa43VhUmzSo9hAEIV/FnXqXFCaFbxdZN9ZzquMUwirAzABUlMcixu5Nk89eJ
uzt8De6ZGRq7oio02r8ue6MYOS61J+YJsT/D8sDIY0d4aLQbIYmef9MyAZA6V7b8
NP7bQZn5/w2deKwojEsVKTeUZ6yrmFccmH27Cg/7RIZtLyqRWtcW6z0KSnN4OAFH
/T3HrQGQR716cBx6g88QqBNBCcfeG4eH2egNnqHAVCMi7I1Foj1ySxlzTMuD34FM
o/R3XvxRwrQvnnw0PvgJMo2VEDiXS8m0/Vn1kv5YeuqA4X+cQTWCVfGeddugwGbq
V2lKlNujy8R+mt+Uuh7zHHmwjYbOckFiV6HvfkqS8h/H2n/WKLZakNyjHZk2degS
6kd9AljxEejddFvre0TBDG+hBVN7l+egwrc+pxXhrWn0HzJ6nJCJU9lFIvn3wKkf
WIp5mEuW1It87OBarzz2EVQyTN5bCfUnaqVtqWbDfHr4j8pLR4Yt1SgibiV74buk
OHhgqLjzOyIStQRmrFGVb8bjesPw2xZsRzxXhbF1ZF8hJkJq+JInxFQnh9EUYNSr
7GZcIjTinKPEKzzPSZmsn+/7nZyJtVVsOUY6d28z1ZWo5PdcYp2SGjmbCkwk7N99
mHuEbPlxI8PPrPnb6XqQTwUgiqKjBe50AXRYwu3CacPkmdNrmAvODnUG5DOzLY1z
naldhZUQpRV/7jL+/hG0pkcaCgOW2ztJbO9F6ogr0xZ5HbCS7ZTW/UkBQJauG9gu
5PdjJBPYLHffvrqNt35fdxb1qS5PpCDDWBF15nb8VEmIa7+r+ab6/yr30NhLUHen
ZyHRvBid4r9bZlGtTY009FjtN4GoC3nSKFIa9Kl47r+GSTH7NalsaJ4I+3bv2ZUW
piUPfz6QGcbqL/nAl24hTdFSWGV++s47mgTymUsP+1ptwKaXZ9NQb+KZffN4IoMK
5BAHqycuetEcIPdlKEjU0bdzW9Ku+XuQ9yRIaNK7XPTtaRHj9puWFSGlpNS/ZIiS
ZBtI27k+t+HTuDDhf6vcWQPbGy/chpFZyLCmhZIEv7sedD4OTkBrwGxd1d9VdLXj
wz0ARnmZ3W1fxkiCvXNCuqS3vaa6yvQsMtptIHllsdDYgdDdptFc7frMEaKH4+mQ
I1GMEoYYmbQ1nUWnUrqPbnAcyqqeGJ5IS+b1gmQaar1ohmFFLplVnEAdWhgskkvl
iLmFztzCec0TDXtLLFpPW2ZQ4YJI8donjXbbvOK/1Qy5UnleT5GrAh9dbdpfnb/U
nSR78SrEZOHfiR1rc2wpeeavvyLz711rj6Q/y7zT9hno4510RTNkR4w3MN/b2JOw
fvWNDShPxOlBVqKKL9rXY4yLANPQN7XLu/DG8JXbypYF+pIF+Mk3mlwsOF3rzSEl
ULttru3YZ+sKGm1qfDNEnoJJ4VQv7tiZqTn5zb22lM5m9azgdMclvk4R623kNVfv
DPyhJ/PtJJgghhL8THnmJjhuG83irKD4Dwa7TRTVuzYHNdnSiM2mNV1gqK5iSyaq
s+/rEf9BwKRv+oV14m8uJHD+HC0MgP5/dLKt6DCVxxSJ1BhE9emsQNLBF6eJsdyZ
hEdpsU7YAB1P4y3vGwTV9f9yMffSQRZL70n8e6Ij8RNx5kF+BsVR/Q+L7+oCrriw
0hBfeW93cmXaV9iQCCZglfmnIMOORQbs+0BsS1SNfFEiDT0AMraUqr3HRQ9RhA8e
AoG8WUWUh0Zha5sKpInpy2eNLhNR08/Cnjmka1p8DUSY+1cSFiCMTrtEcIrmDBBX
rnvtMzPu/+vIpNJtZJ851N4Aoc02jtptd/3u9lK9kEO8e1B5qP1M45j9xOwjAoDA
Ik2748UuZqOb2CbSUd9fSNGOpDJckW0yLvLWqzqOKfHOy2/+EwGSDz3V1mCA/QG2
RLUL0bCnc8Fkz9898JmPJ5jOohLpXKGahMIDQrCzrJKSCz13ZDp1kKg1OaVjP3k2
je+yiY1KUM83Y9FsIhGypxm6zCN8Oz36GNN1fbWxTbSEp8WLaWlbw7odicQdd1FB
AggEfjoXSMthiWvDqjSbyAFxyQgh640LT4tyPhFzsS6ChnFZEv02s2ks+vvykHtU
rBb9PZwZPiUTgUlgGPagQo2WO4GArf65UbOSRj/g2989SqmQDYtbe2HQ8X6TlWh4
n+prSWNfyO3yDC3aIQX3hN0qKgA8gEZtHUVznPrBs+B+UXVupnHEWfQdbenikYTR
qq0XaHGlGp3fmC48W5J8bCBTxu7TFtt44RHi3AfqdfxE/jwZuzPjyPuz07CWF+dr
6ZWtQdzNpp2kK+9J2imeFlHFXarfQ+AjLYkUeWryJZo/SRuFWl14C7ggci9iy84D
pskqYliV4JfujE/m+b/Xr0SyJp4cmQ2SX8knuGUJ8jCFc3qJ6aVznmj8H3NAORKt
RV2ogn1YwJuM5oQyIdr/qVbPTUWX7Zmif+vMCYdHKoQ+cCkahRWArJXOvIxFw6HB
N+llEmrv+5RCOZ4mk5Jp7TQhv9LtFQPT1vn2RWBm8RtNaL8sCjCjV+thyFCyr/9V
EG5dDfuE7meoXMbXv5220xCHfy2ebU4pPeDgouVRuozzXEt4H8dBIYrNQttYJkYp
86S+z55hExpePDrBXjFzG1oirirCZSPhGT4lPKBzeimXPner/hESEuTt7iQ0VMFG
W2jxLA+MT29FBPLUcz5J2nZwO8Hs8Dh7WIBoSmsHJiALpJU5h5bQy0q1wTgszMWe
dIZEKerGpJ7xxHF9PJwSJVPQR78C88IpDb+AoJWl/vCHt3hoaNnoEJ2xCPYLTk2S
eyJyXlxYkZ9hxhU60dgrbYwlzQv7oaeBJ1jP1LW8RwBi/KXWcQmLVn5yxaLJqqdy
DX/vqJbS6KYyx0wtivr8pZsUxTCJGhlUz2nDXJtlF11VIKn4dZlsT4LYG3kHqZuO
0TB1smFr6+yw2L8WjXPaekMyDVZiMaVqwiED4zpSgjfiqJTuKsZq8o4TLixamWEU
pcL8m32aw/ILoBLKHEAQuEZuNbWMMmyp9+s4EZvSjCA1qIFfTfoBU8saQmarRnZH
uYuJ3ALinPEa7kZ6ZwQ6s8kJURgVcTAP5QeesJA4bzqJk763yAWFcSyeEae48pT9
fYXEgLQewpx2SxFusD4Z8a3VfXyD+p5f33p6/YZq7tXHumphXkf6T0DrWKyIvdF3
M+ZLn5zFY/Vs2/TAy7T+dPcSI94Tf/smljzAi/Obhmp2Z9DSxkAm2Y/frbwUKIoh
05eU4R67n8iDsBhdoAyGJAhlJffFFDIHoTbaZ8alMZXqgeUrIiPg84RNOOwg6VTV
9xGc6EMR/Ogatr6wqpj9P0hiHmHG41S6JJ3NfeG/vCtXscwTgi7j1k125Nyfar8Z
fzoW/BACzIXtkxXLv3a9pq/6fqZdb9Y8CdDMtjx26neXq6wzxbRN2dCHB2ZTJ34X
Wb29iN2+9kCUWQn0Luxm4uoedbmfT6uT9QSCS0bNH4qJuSAJJ9jg9OJSLxci0tAn
v0hT7VV2xxkrCNFZGJKxDoLe/+U7LjNefcjM20Bqq44TZBmT91Drd2xTW7+0QmrS
GoYpuE50KtvaZuiDIupIrFXNDRqoOHp+pQ+xwavTqBpKgGtVWGJg/w3tRw8YfW6/
ti5703SQd1DF8mQe3n7/r2TB28L21xNXpxwJzTCNRdzslp39m65mIeEH3Y5b9LdW
87f9MA252IiAJJ1iGLDY2eltwUlcWanXAs0YMYsx3XWen4AvWz91Jdvq12d6/akL
m7mNKz0u6Ro4Y5X4FmeWL4Zau8xCCcidIfPq+g5PLvSICNr+JwDkzBJ3G7sfKt9c
/eX+oFZk7IrRre7OM2FzaCxVl4Fdp4ASl2JSN0F8xYcJflnYzWEhbeChjuRMhW7O
7FFT0QVWUC44FykKV/Bct5qw5hPqzQPNPra8anWWNDexczRhMeR1MRrlc3PWKoX4
OWy5Sc6PkKysXAvIIpx5EMDTSbO8r4HoVpzZMflPI6YYlia0SEYwOoKxERY/cPN7
czPlKPEEw7VFHvNz4pUCr1GOXwSXiBOdum9TgrW4zVgPh9bobOOVl7JZH5Pt5aOx
0IK2ZEESEEZ5186MSx8Mn8zVqUM3fQS5kTW2X7FGTTUnjEUbBqSSZ4xSa/vgXvbh
NHAu++cP1I96Ep+4CbMe5hOTxoEzBoaiLQFRvbgj97Jk9tcpXsdEfJnzpjCLH3GH
oCiv+rwytnABkk62J6b1ODcKwbsqkbn/IAO23yqEkpr7GRgtOvwFGAZgIA3CbpvL
w7JoFeH7DMEtnUkWpHetKIsepI/bC6WEqdAuwpKqu+Nny+Zi0PVx3cLfM7lcttsk
BG52O9FHi1c+sIbIzPqNA2KQ1vfPeTWyaVmhsGOCK5diZ5OFudAH9aBvgJhsa81t
Vz9risVudrvp5HPy8I55bQ/+zNw2xQjRCEjWBrIzAbg5iLtnSJrj3gMsw170wd6+
lvlV5UKm2UDke/84bYsZM35kJyLm/IsySqcZRoer2SxpPspz+eGzQCW4XtY66cXO
oXIgYDRTXCY20xaWL43fkWmUDtsck4oDS6Uh5X53HHLV6/fNFxRQnww9k3OvdGzf
4ENaxAOMM2opPitjms+aiG6md9pnA79HAkjotTNfYwSl6DD95PsCDSBWt4fv1iZa
kzpsMSZR+E1zn/yhhb9FNqCKRkTkDz48RpeDQu6VDcZZfG+I8xVXbU205v57+7k9
XNHx4znV0J5NCa1BzZSWROQuAY5mAHjvGQfqdy7RrTE3gFhJQVGa+waAAW7N/YJd
iOv5V7MiEOyAfQ2kbxNs1SGU1MU4bajEMSDFlPLNEqLgQefJ8x+luINcD1yN/89y
PHNNZsTqjwt/r7ym9uUn4MkqVNQk34xkKkcbN6NuXeqLJXXUA3CEEPlfBuVIOiLP
y5eTaKEfD2/82uaq+uhWCl5Mw1bzWQbjsjAuX7IvJu6f7yJbVm8Nohg0FoaVUcvG
yGXiE+70Th6G4dZkvqOtMBZc2ihrwxBvNM8hyTF5RD34qechlBglCytqozVcK0x6
/veHEmhHYpOgx+1mUiLa2xV0n1l0WK62ZaFLLimMT9V+1bKrPZokHOhGS03O9L5k
Fy2pNf9ooL/b76g5L52jTzGDmdqxk1MPyMm1N9TYBTK0MgBpJ1/tkqvkWrpInOcW
j57qtJqmILoZWHq9VeXV3Fjd/NrCckt8etPdfdnlSat2Xl3rHfMbCTxKP7OVJal7
dt+bT44lSZX/o4OUu/334/tCMN7sfAIPyQvMwL7LDETLIFeSIlFh3amySzBQFd8J
tvBqGr7v+TccZgDDS0Kg6YBW68DTsJRPcA7E9jTzCm+ReBcm1cGUJgrckXryF6yX
EY4US/ix42euvfA/HewbqIIGeG3W6d4wkScFsEqrJb5blK7Jh+63CS1/lVE8WCUD
xwsn0KwboKvNmIjb2dP8iHgSh94ksokcwq9KIR3hjmgbQxWbuJIEP3a9wUn7N4UM
opFnofIS7fR/yOHt9MRk0IEz26umALUKZO96SAkEliMvn1UJG4nf7hkuPUEGGdod
o6jAglW+soi++OTkzzPN/FJ0anIMsNVCR1cnvYf/Z2G9O7SDX9iEPvYKl0+jVoQV
dqofhL719CcdGcsYo/OBe/93m4mOCF/6RIbPOPHnvpuvxFyg3D5oIRblxTXr8WRy
O24vDQElpCIzp5qR5OxASkosAKErCl6rF4RAQPOyDgLNKklblAZrSd9AfZap1+ub
fuNEL65zVPtZnbRQeyDbjM43CnxdqWKJTVsFT6SKBREKtvWrDSxcP+YoGpg5cxLE
3+qTE86jeQPF9fdENzfZQvWmIEfDtsvGAP47LVVume42mxUbEC+3C4pnGg9iz0Q5
sAV7EArxcDAC6P8h+rQeU/9eTLli3b5EU97nzYa8EPaDEQcz9D9P+rlT0hHdCWFC
4sih2zqONV8wf6nCNmVD9e8t84rWi0bYPHASymXKX7uD78FSS3nq3WPsu95L6WXP
1kkD1epDDfCRqpk04l4OuOwphO8cTUM4JID5Y8Bj1uoTjQ1iYfSd+Usf6fReFKLh
pRHJMKKAVEX8j6RIeXX/pWFvlS/NdzpgyzqXGs+WVs5HsTIJiPPZOr22rUVN3W8e
kXTrLPpqv/0CVAK+ZlngTE382b3iv6MMgJi9wkYppj948Z4wVizImPFrgnJG7zie
xFKy/aegheXkqD6QLWvXH0uU+1imeyuPok4qCITKH+G/8pPivN7p4++yEk63+JuN
9tBl4rK4vp6GuJmT7IwwQOgwdjb+7F1l84XNMswComsFoi4y88XE+Dy6ywPYLqG0
L+g3xyh/0DoTR9mn5ByuIgX7vFA7WBrYOG/xspcVE2NpNgmauLWb2BpdXTD/lA+i
QkFLQFVIueuYYVrT0hS9fVQHd+h1Teb0FHP7dX6y3bz4rl8XKARRnjrr4+o8jDx+
r4UZ1PukwWny1fntN2RT3AiKMCLFuCYFXiPPNX8lFjq1+cQxTAFGH1yeYt9+PxOo
7IuF9GBME94TqgMsWaZgATbBq1gDXRSqVIbW8qoDtdpdLQkZ+xtJQt47EYkgH0VK
9r5QxoLRqYOD/86rFVuHtLel2SadH39C2w09bGIga/VFeLJDm1OYbr7z8Drr+Jc0
757KuhNQ+LBUuQxE27FP9c3Jc78B+bl9yLeYXU2lsWCwNtQCpfNqYPI2KWEsCf3o
bzH8mcODnDFhpnQ3cJqNywukFUK2Z8uZSQc47xCAzMZwDBwnR6EGNmFIWC+Lc6F0
8Mc/TdT7cocfo95bXixFfaErEkbrwSVFAoIxrtQOt2hS8MT4b/E501EEU8+Erwbh
zceMoTGUvefYVtp2R7ho8mpYrfTMmKpSZ3Gd1I+LFDEbucku4SdcP5ivW64lKHYc
X8RvXeiFza+bZINEfNhqE6L0N28pWKsFbj1fW8BuF0oXWeNa8T1K4s+N8YycKezi
dAqNKDbYb1quk46VoqMvL/7vBKA/OAJdD+4KY0mWTMjOIuL6WiaGqzR4uDpsvKOQ
SvN4R2LGxHFi/SVKlZuvgInumKt4eLs4A+FmqriqHxIA26elOrms2Oc7nXANQyQd
OK3SGCQkaMbGRtV2W+CFYcDVYIQH+lLaWfMeNN8arkWv7MwtL1wHzCouHxhJkHXK
l1/Y6swU5d00pNEg3LurWy3gA5vAo13h40FJK+RZx/q1OWsZsejzuzAS15jlLy69
vHaHZx7Ch+9FXWuJRaoElUefRdzG7/a5/jAiFHa0UOXF+t4/nMB2ivaG5uSiUdvH
s4vChWIqK+U/l1XHxrM5YGKOgp+0oYOtU7d21zRMy/bjjuWqapnLMm39XALH76HZ
1Hzsul+9LmLtdo9SJPMBhw5qdq/evwQVxkIQynFevElsISP3IvO/EfYDAq9KrJvX
awsEGJywd2o+MJOE42/Tyam14pdDQvTnh6coxKOOxsVVE/21viwzVh3dRd569Lfu
jrCghc8w6z1cNtoOIZ2Ay1yu8gN7ACMfdDWg2YTx92Pf3UVJgWlCR1BCpm5qO8SU
YjluS67i71UvqJPm9Gx7M5FS7ZfcEEyumwc3ZMgnOvAlsXD4og9SrXdE2mJ52ogk
0UNKzImV90qXNQAaRkpEyVZUgr8a8yKK6zsNa032ynj3TWOad+i6yworuU/+EEMD
VhF5zsAOqpmtYPcCbLaLdtzR1PwKpYmkFCFwVxrAGcKJ313SZDKH62ktheh04peY
j783LNIuAy1gpyCdct1OsZzNdTliBugfmMyFjULH4NgEsqyc3LaFsDW2tam2H6bN
WEaI0F06f5o/B6IBaZ/FlBJSzXGJeUR0OWC+7vFN3htDF/39Plb2hDv6oR/+ms6c
71te5PiyAMcMKtwtkj2BRWTZ/PaG2eVYMopdqntDRB3i+6jYQGyUv06QRsWgaGxx
CaX4n8ISL7PtpTokK5HNrpc5kq75cwOnBd/6mBGrAHmTq3ITal5hWGeE/uvBGEag
QjYTv4vbPqR1kkFqOYBMMihkkw0bmS0PQUi96X9XGBcMmZsv1W2g4Lp55bWo0hOm
JPaBxKhdO7eat/L/F0eQmN0icAPpDIceDhXk0NqSmThJq/YabkVO+CtZAEZIrIMx
2HUC43//c+vefj1TMfkWiuPFwzQ169gQf6YKelETw8XkRZkGczskLv+50CaEk1yz
JgoJZ10oAUPBbIkkwVHb5RLB8YPTKJOA8SsgnCNOhrVrf9ghRcycj/Js5LcGWkLf
Fh8M0OSm4S5OYBlVED8qf3Fnefhbumm3F22G7zEUErIrXu5aUKw3JCR55F4wlb8W
uj75LQTlOa3byh0gl6nKbZsH8n2w8Y/RA7IgOUC3qa+V4V1oYrF1fXJ8PbjHQanD
cSPgpBE3eafJjTSKJcA/C9ZLOCV0PBM2NDf14LE92IhAETspDn2Cd+phWj9tBrSd
hNaXstPwt3jQ9nIpsIgyh55+VPC6tto2Rie021HwEY2AQOzJxrd4rGd3Mrlt7iLK
movJGV4yeOobKfq3XSZEGKK7DXNmAC2u8hxUohotrCuA5k6HfTg38uvBO0n30jsj
k5XkOFTvYEO6+74TkNqxz2I4n3cwgeVEgE7Hy6wBlrUR5lYNicPvRfyAefD0SlgJ
30TrDrGAY/K3C1krvLMYa3zRA2KfQeH1vlH5Unw7ybxZ4PgsVa6QjmkqY0dLLuC6
+TECbXw0CRSVs+6sZxELJyf+tXgyMUi+MDc6htDRk4MUmrCQTrDFnb3HL80j6JtU
Yd2/zEzasC975PKuKUberfSe7lNU1ec6s/keWpdR7oDJvSm+tTnYyzW9QkW6d6jG
suQaDk43FOta0pf9V0hyU02gjPolRICMWxtI1aZhsgOQUx3/pN0sPMjGpqH1/kL/
8Zjj/m4GYMQ8yYOdq/JZcMx5Vw2ycLUJELpfx6ZLICwTuIi7UhkEGlrNWQA70TWR
LV0PrK9Gc9mQblfs+BEhxCdzAA/pZgMclR7kF8eHeWFDQnyL4aWR272vdO1nfSqv
7pHb9sYHmJmgPgcTYxPvaT4LFcFs9wZLLy/51zPI0E66p541ts9GQN4v5On0H/zu
MqpAjTkrrlsrj/liMaF4dYBhxmKdRNVlWNutSa/iSvVIidLLrBscNd+q9Ph9bleD
AUISb5k0tD3mnxBvhzS9mC2+cRd+hM/embc6QLfoM/sFCIt7/C2bVRiwLEihUi58
gzCRlvmHYGJJwqgSDdCiglhhFj8fk4XnGeNiSuEEOAWZxIrDcRKUPRM5b1nzKyHt
/E+5X3b+EB1J07ZpTrDhLFv+YH5SVLkLgykWPoFSA2hNJfKh8QcNaOKRnhE663n3
1Ob3NUsMXqVO2ID0RrfOrhImA7qdctLKKTnekCWrNTLn4VzzFvO8vyNVf6q+h7xD
rllv+3vFZovHRkUJKw2B6DOvmHj6Ydl8xX/sNDgzLBBoNyR+lzMaxmkaevpHpmBH
VuGV9BZNxAtZkW11aj8MvWhgquIJyPcu/L/DrLCD2SmL+3AGj1T+JvbUFb0W12eT
LQARY0vJ2irgiefSUCV5o2fwjuGRz7KRVjmN9F6Z9VUGXWb9q3f8dLGq0fK8IDPT
RWic2plXrXrF5Jwk2Tq0vqCNE4ibaCcw800+2DXZ9NQbzLi5h7hJ/i1e+El4OKZG
wQiHy6GrwWPpVF/vH03tyalD2zI/9J8Ir7wnApF8LTvm3CXi054wjPEhvhGBkLa7
3hzOC+Z4WVh+tNJ24iDvwIS5XEGB/te+c5/uYJlRhrJRzlLYNZCAuHb5JMptiN5j
UKYQodx0mAP4odDONKnavNLOv0Uo+QtNH/N2ptrKVfCCzhir/Sp3+DfOIsPjwAvn
QAtZRIiOLXpkiNoZTriYN2aYKRDUz4jbKwrPvYFBeIeCDfmRrxe+2eunTIYnREBY
RFzjcCuDWll+uklN3V3Ik/4GK/4M9a47TUUIi9bpJd04K8/bI4+8Mz2qnlApnpCZ
7dgtczvTWqy8tbH+e8ELIEHaX8SqDsKOVAoL/Knj4O0UJFwbaiCo+y8qVdq2DaPI
98qVz9im7+MTM38u67iKqi16uE1AkDt1vXrGGO5irgoBZDTXDizTrrx0hA6fS/OH
Y4+/FyfH0AgCxXiU2Lb4YcK+eu2xzXxgrAUEOuT2kCFNKGZVC60PYe8C36TjMDjj
JwmfokCkiPbuJKvmJKcxBc65VWNJs+nEy7XjpC7v3qH4xFuv/SYMWm21S09uIywR
+/In0hNCSi0PYP/EVe3Zh2h/Ke1XsHAITrIodYNEpRfyxD3m4MgH1Qk1lVMQLNIC
GCp0U+KADaCybB43lMFR8dWAW7Z237L/5Q60K8U0qe3yL+KPrTPvUGHQSK4Ki2nI
EuAqiQGfKGX65Ik/sbTeFFFK3AUlIAYcRFVGIw+c00g+vx/i0X6EK94utgsFl2d4
GEwm7Qq3LwCY2BMRBxZBv8DKwV0wJhK1+g/3hBn/MGVEQb7/HZM4VU9T0EyShPYU
pWaRK8tdauvcd6TPYfqCFlLw9s9GbXaqKMh01xQNSreZdS9aKZA8VaoxHf+SuCMB
gtQSvL1U87UgO/rgvC5e4lNlR/szNCUdMfcLBOSe4eAbbUQu6OxgO/riijOSZ9W1
lOF4/RbWW0p/Cyr5jjrCEJvS7fYJSNJS9W7grQWbfuTQpItgeKchTuzfQ/jBxLY5
RHHpY6Xs5rEiCojEHZLnGt9nVDr0/xTG0JB6Vyk04m7nwTveR999+3a8xD/UhGrv
mSDbRt7r0GCXd9Nfu/2KrY1fgyU7E6XdN/kxFpv2IUbrVBy8hukKq1ajdC2Xu/43
Ubq3VMClPsziu5YTrvs4xL6iKf/AOyJgMh4cL2albA1hdBa0AN397SuI2Lp42TVJ
qpatVKhh9aCmUSgYY0Hms2gk2xFgFtMGpTvAqJyWZj6NpRYY9kM/8f/ifp6VK8EL
rx/rtccBHcpYwGiZ7ve9PkneV2KU60LGd+gG+Ss9fSzV3AvU791oJ291lTONsRnq
xzf0j0djYAiZD0Fe/DIqlqQn2Z4FS2ENHVP7KW026USTeZ5C0bH3rPpbjbD+SesO
RrrVsvhwySFo0xbM5uA4F5iTbCwsZzZkn67TEuEJ4kO8MODXI+mRRi9qnw++qAH7
Exca1c8IH54koe2zztB4tRT4a+HyGlmyFZF+0v4jlcKkf1jep7CDyfNAp6U3EQYk
1b6lddTXZuNpcgwNUyH77ZAXKmKtCvVhTdG6yiT/dmng3S1v33jxygvY9oWlEHlO
TrZNN8Q7ow4tqK1i+6G7hj8+O7hC6UGJFkpvukxoRnJrxXJDSVCGUq+9T/nCa8tQ
EzDdef6eUlu8YpTFiY4vhQvTboaXnEX6qUbBM1PnWe1xwvSJ8M3JUcnGhn9wfIQG
Umb16GF2WDOAarQ5VAm1sB8CncoiftsoO/i9svg/4cWZXLjXNwbQ939qu4DTvOUt
h7BORRg/XcCI9s2oC6JLMB6MaY2oMjsjbFtQ6eFBFLe+isUqGJhtdx7h42kUP9sh
2buJFjcQoWamWOXa/T+jLJ1SvJWOZ4ORDTW2tqFlfBCqzqHyP2TepwGHpSwjiNFu
RN6GVAzkq+2Hhul53LpBJ80TX1EBu442g4zIm9wYvbc88x0+Un063+HdhMPKwvSt
OtDRBFaEpUxF6xWs257FDmRj4mwJoFUdINm9sAGPHCBFTrT6EK7Lj+6PbBNHXrA9
i+5kcVQ6aqsSk0MqZ/1Vrw8OT2I7SWyuRv/sRyw5U6YX56wZ7Fnwmn8ERjHdh/O6
4yMYGw/da6Mzc87XnyHawA/7DgIqcjtvPhi1vId6uuKX6kLXTaUOjnZRt5htygJq
u2ZquJpn8MXIa/CI627d2NMD08COviuNCiGT65FjhyT/Py8r4Kpq8iYIQbmdUkQR
DpCmNcoL5BscvCI2s6PF6b6xqQLW0I6tM6LjtyxBCWIsPfnI7RG0crNeBTX0bHtr
XDocdwF+gyDdstfXb4+YGEDtN+WwMCyQoxrVIoNLPIKtN+WDhazNHNOHRDZMD7Yp
GFNYl+nYLttnnk6jn71j6k6heEEXufTv/TPMIWrY7D2bZJkx/tam6mMCyCkllS+s
dSAx50acIz7H0d8cQv5YyEP4ysGGni7Qu/J2fOJBVzsEYrQ5dID8eP63UXzk/9R8
n9BT+08nsBuiM4BCSQgIziKyPl0naCGySXm2iGiPMf1bViwDx5lxJ1PyCYpFN57h
KNCOnRziUrC5IaU/nTJ+i5iLx7/+9waUaLMSlJbIbTEUDVn75/6kcUrK4uwLpX+r
XvrtlwhSxmqLS+avOdHCPNGhh0vB6InMzHjljv31wMXIHLFQHLas/zBYXjKIfnCa
AiO7Zwcbr8sshHWfISfy8FsXdLUyarWOqeshRuTvNmFa5uP3vkCjPziNqnwcoqTR
HRzft4klVh4dszxKZtBCCKA9H1seDqSGYObK1WgxrwekAiLv1DXBRbBSV5L1VFmC
QwB0Uaw/hHQNVGRirlk9IZti19z0u0gSDPT90gT6zHw8YUVZRf6UMh2YPiAaRH5I
I9mFKuw4eIjQpP2D8d6xassVJJXdDMInC61Q7ospBxyLHmjh5PjCtPRXEObcoiC1
cqbdouChteadFZwH0ZKO3n/ZXnObwLm2O04eUU5ba39jzT8E9tCqay0K+Iqa1J+V
tZ2h7F3e22ljHoIoGVnjZTzrJ5NSZJPKTKPMtJ79EvOjIPJjDVcg4PufH2PKTqoI
WWs0F5elHC/OVaiNr1y0Qtbdqj+pUHm9r5Q5MHNRrufH3v08vobFqtBCg3GZzpn2
Xq93OpoLSgpW+TbbwWRw4MWOhUa+Wx0beJrxGPZl4FPms1i/NUOCMm2x69B4S9J1
fa1+JwToac6XfvkZQ9j7+9g5HD/ePyknad2gb+SM3WNqTyzewVnnz8kJTTr6pEuF
er+ZHSe5W302iUId4YvxLu+7UYevtOnCE6D2tYxySjd9GH39zVEhwRgTNxp3f+1b
j+JuBfUclge9dVTrFQG6Z0CmoyCCCDgbysfNuEcA0Bzi+KlzbqJ8GvNpKMkGH1Dn
AedaghiH0SIhhVRqNSyZ+odCmOueubkAZ6WlTgvrlko4CpK3e+Mtrg2xsfVS4F/s
pWihfjw01t0o0X2TZc2U4Sz40i3TcEoP8jchK5UWFXO1ZJXfftyQqJScSyHdFbFr
2GWz/iULK2UgO4r5x7MvEYPxG4ty/1XtnlLH0soGVLgsNgpKl0Ua708lexQ3Ce4i
UZR3Ur581bLK6EqdQm1LAbgvToUDUOzfJ7v2glci6QPYgcwGrTHapSdfL+6CAVQT
6xbL7XruNB3lrBX6qNH6sEUWCVrfHNO4LCd7IxcYCluYaJ23943HtE5weyy8V2Ic
oOJLj6hUiG7yx0PKFx5lWu15YdcpXY2mPu0wqzEkPsyiTFjBlQAPreSCDCNZ2XCM
2yVsLkTXrXwL4aarG7qGTuiTsA3gL7zFUHuZqC0LMsTNgtJDf6ztmN9sNuaeZZTR
Ej8Eg6IKWfnJ5+8PGtE5BK/3OrdDGe3sp0IWT6pABM7QY3KbXTvDPX7EnbTpPIuL
rmR3hkUDBhgJT/IG3QzkmkLVxtnKZrhdeDlijvVN1/qOrYul3gWPpXvMFvhURdnL
cH86Kxsq2RQme0y5hFBCRYsS2vsi8To15eUKbQa0vDi45a3pXMAp/nXx0juwlDoZ
cN+cv0GwsoqOHvGliekKXlg/fZfrCmTuOf0O0pTgdL3ECuKrTDj9z5/mlC1Qgce4
5HsW/aBV7naE3EAyCijWaBegllA00x75SGkpsL4dfqJsJK/Uja3Y+MR3hC9wIcLZ
fhc8T4MBaynvQ/2i82XyEvDGzHYVQJDUhVrJsrP33GvzVKMdbAkthQfV1qXiDbON
nIZ3RC/y8ajLaJ2EML8Mnvi3BKsCOAxRzq8laWEETcfD77geGmIC/lSb/44BCioH
WQi4VNsLVeo3s09+fUQKVOBLxGCKyWMPw0ccfFEE5X/wNWNojE7OZZPc81nOhtM8
nWJCVkJtU8ij6B/dBwjO4JqX8SvPclHunz5lc6uF4W5aBuqDxpP7GirRJOXfJsbJ
Gu/CERlg3tH2UIrxsMXGyWryajETKhGbj8VMtR235IkAlMS1PWYlk3Q/MlfmRVW6
9KOYgaLaH1CnCjp0HJAVzVSp4nOUiJEWlyjCTx40JWqCELQC3uZxCysY48QKdHxC
kX79XGfKkbsA/pGblJRhHVfLW4lrtYta0wj0e8vP9aWR72bofyq0379EFlej1ghx
cxfFhkOu4l3veQl4bKoWnFu3pQ9EP4I3rmzb4Iu+SeGND9IfhdjyA6Lkj2gZ+gVi
8K/Gg85HXF5E2VLb8CRZvJAdk7o8Otzl8qUlWhzHjVAxSwFVKUeZFhaSauAY4Arx
XDoUVytUldxsFz6TxLXgi5vuD91hQ6ovuawhXVG//J9hTc070tvsCPCpXAL3Mgzu
IyU62qjtM7yqwPLyDBdE+2xxcyC2CvHJERqbvlV2JmS/K4TxeSmPNJ5kcuzWloVj
hZVGt8QyTJFbeVARyurpd+ninTOsfzPNiBuEgPlrVEPTP19eL8V9kCfkR7a25kzg
5ZKYnaqpUXBgpeMk7wKB09UlaLx2DYfW9bMQzW52JD3oEwU7A5sOKHEE2DZXDAxa
6WOq1bBU5HB491Gv/XbYQ5uyguZAf9Pp+VmKxmMzPe1w4V7xDglfgGs4vJlGEqrm
0yveIb7p+X/WMWeoVZXuMfp30G/y3mKVwG79rb/mfmBp2H6FV6G2CXdAEYCX+39d
BQJh+KSg/kkw1AgOzjpuktqSaiRcmT/BbBZi0dqmqe4qwBNweAD6hE/fvE26DYLV
BxdGg2Ocuus1K8KcwX5zqQjO7Kja4jCUiPB60V8bfVU5kuCQn/AYV9HOwF20CdqE
1DhJzE9PxpzRtE6qHrTwsTul1pbiYrRWirAQ8W9+V+mz6Y+OsuY8UI130NsUg5Oi
UsR0vpAv6ERBTR968ouNCSrjZuC1kWpC55+g9zf4FeTTUZrlFS9jPVQcf0eF9W0b
dBcBo2TGzYe1tMArhmCmDgz+KN5h/KEhJGF1VQRkxY8qwJol1reAZX0WgjIRBmoJ
korgz988wetqNWNj3Fy5poq0EGk7812Y5bRyXUz+rQk3q0PkWIFrYbWVRfABnxd4
uSkRb/eaanujNe6dCmF/hvtdMS9tLwIVEp/3sGX1ENA4Gy7XNEGpTZ6xkq5ScCUD
gw90zl9qZCCNYCIdQuFchohjb68n8VhRcu+9Rxjw7iK3o9na5yNz973IV/VgDFH+
s9RfdmVQX2wDAcARdLsYcs/tj9VK1G7L1SPDlZtp6Uwr1nEp/H/yx80bVmINobq/
/Ghanve2QkClWNJtCk2x0TH6oz4vWuadFjbIedjdMaDA3q7vqxXgpH6ZtY/k2Qfd
o1TablkhbDBaFOvwWLoq7pPmZQza2mrEaiCk5Cj8pXFLQbTvpHUE63aLX5FkCMLg
kqJqUa7PZoVetc/snS1cKqhql9SiL8Z14RDs81J+ye60z/H5I4hUR0+/i/nHTuMm
+bMO02ntjTOUQjIskcm6Y0NkHYBeMDWg7PVMdacZp6def+sMhlhwGSCx3IQeFm7L
qKkcNsOTn1H4KfDIUJ/lx2vsR8T2rO6PJC92RHUFf3ZXVQQtfIR5SyM5m4BGAXbK
72hv0W0QwoBNslXbbfqsn+I0/shoToXgOLXVPibggEt6G4ypSU5bV1qlu9svWzId
7HSSVLZqrjdKGRbs9Zh8DMVnqNT5/M+B0nO0xye7mQKXLih7tnIkUODnJeJTSyFa
E1cF/jUulWjT0Cf0dZrpSROUfEJ+2vznSZiwY7w4nhUShTNfqSBs1GiXC8NpMJpY
8NA671m1yng4fVhnmvArqaOVwLb7pmCPpzK75OHDiPk2p9yIbECvrSlnDCXWR6ka
NhQwDBNJX31QuBIJT8mJSomdfr5ZPtNipwzbUsdykbPT04IBoK0W8refI4j1tsYs
4FWBiBqvMipdIjIlTNDnNsc8robwjMHafIFpIP7sGkrMdiQ79AqHLRvTaR25DWVs
aa2xFdsNfCsJ++YINR/EONSFxigjIYj2Gl6f0qJotdfcE7Ui/1aQNDAJiypeXkyZ
jWCmx2ZDfsm+qemNTs8GdVZQUukr/y0HfxdoIQp49vokD5SEwX77jMSA11CfWcxX
gW4ZyAhCvRoCeMi5fbcZzJoiuyucsPcSIeE81gpsGTZXm7Opdz5nG/8mA9FyAiFR
GNb+odVvvdMVqSCyarkzQAA6RcLS17XCSdJ/mqI8iHLC1b0Hc8c/F9HqvwiF1eAh
5ZnEak61FM4IvXSTIjXJSZDSrkPE297W9CgPf+m6XFwPMBKrf0VAkzzQeh7ZvLb5
RIXxXt5sCr4hGRpdA2hqY42Pcv8o0cafXih6V6N9Ua5wKq0rpROCVNBrOjCxsB06
S9O9Tk5zbKz2q71Lj6G/DW1rz0/9IKAGwCQCGaAD3D6UTg81qeJWqHkYU+RveWuu
+XLozl8mNKiOPw25vx1/XluYpsOts+933rhEP27wGl5UhmGAOcWNx538rRpTk1OW
etF6T4n8Y8YezTnlwTqeaQFappQ8MUcHbEMwegQ1MdhIWZs1NzbOHH2YVBfnHQ1G
C5RVLBNaAYSXxxgQFJMeKhegf0II9QiLBpe7rcAxJuVOte7ai2t3Wc/QZI8UVcpz
nW/bfdAm41KXUKIDkY1PANo0VInIeD/2wjYlHTiyWHrZJGqHnr1Nx9B1IXH1//eo
pj2YG+Qqt6WIy9jm0T8sZm8EDoYwafq/3LlQfLIBUnNtit21h2/cCdCa1WWPj/7Z
HsZSAtKuRfQvcpYFHPvVGyjJRFrp39Qmkzg7MCGyWZN3vObo0EY1FoZm+AekJXDu
uriXno34goC875WlaPH3Ygc+pqFU8dW40AvAMmaPNU+yPiFDyMTYXYezX4SOOCsE
SRF4IPnLzEunILys3wDYzL0PT8Q33vCzSD1bE8iFikUjVVNNsIlwJmeynL8FNeTy
9o/+zjQ66vtl618Jkk2pIsV6E3Zi3p4h8YSDPdE7i8iX/xjsvChpI1w1l1FAC8wx
tEVrceVVrnSDJpkfQWbr7XeAfGHpKCFqbyiiliE6SoZmvrKmW9Q6lsr5hbPjUOjQ
AmTJGExCVBm+0p+nRhibP9pgGpL83ekWtmBL/eaYjoV1sIwuHEsM51nSx5P05DU4
7wvL1mVW/sYgHRB4M93jjOOVhYIJg2P6ptOC/yh5XviaJfBKof3W5EMrnO3hWUxL
H6uOhJyucegLHst6teH6yc40dmLC6vG0ihWx/1EEhJ1S2jHwvhddfWYwxYs72Dy8
h98Tvu7m6gz/VsiIlIhIdUdqD7k4o1kLcO5tbHjUN09eCa8f3YfLZiVz7e78UciV
5Gi/CXe2oIRXk5/hRhqYXQ9FCk5/V2raZ4pBJ3Hzp+m6JxtoMlpg9Pajl5+WRk6a
5vkK7kazF2r0r0Ca1XP4gJDeEr+9e04R2Lwlvc+Hrwi0o2ll5lE8YVO1+qCo6j6X
AKouv8aoXGieLWm1/nCSOusTiU+aMeqkEkwrhmauBFa6dABii0uaMEGTUM/qCPsD
c3kN8hQKoDzl/5q35nQWQiNgpAuXM1jyiye53ULT/wOPPT8V4bfVen+ldswY86iD
rvAuskhiHNbEWdSYMPVxVNxGtz9CdqUGUtptXxTu6RwLfVd/pAinwRScU3viv4ee
m1EWRE/R5NG0u7wYOeBgGH8fFHDhWYYncBJ78oZGoR6M3tpEnlA6RACSQCp6GrDn
QmVM06VdbX459eh0xagXtFlYF6xRlFkqnhe7v+0W2HfRk/wPgMj9aTs1y2qBsqjp
vsUyCicDpUJbjp/abhKo/H3nsDzSyUZYrB0e3p3uonJ8ut5AvZUkEXMCZ5eo2dux
nS3FAcgdiUftj4AYZsBgfE/qQLtidG0Cknds+BW1icHqr4ekwEW+Xqo5YHKFyW6S
FIEIY2aceM/ocxIhQzQPI80KVksAy50H8RMcrezdYNbQ5iYe0cN46GsZb3hQ9TeJ
6a+Td5NXgJZxsnZoLvNfAEFLLhQWuJ3xl9q0HDMERwZ8WFlVQh6vPOKnXy60RWLy
hYKv0Bq+ndmiL7QEfFV2/gzwDUAjaJg7pvtz7x+9ddwb0mRpa6IjEP12tRVFRt1f
HqYm/JOg6KLhbZ3upGECshDD3P6WDAS1UT47vNDV9zZBGRxIw57nKxtlRoJGBupd
dmjbwB/dpeEFGbF1dmLCOLl0YrZOaVLdNmbSE4HjpMOFYwfQhKZafBMovVJyV8Ld
tnA9hNR470C2/XBDlCJKgCf9UUcHFWq9nOX4mvmUYag8ez+0Ug6uoWnRdbWKbqIl
VbAjOWey9jmBsSh91GuF0/USwyemfcSDFmeOlqkTE+/GV8fiQ8mHpkhRKYFrAvfU
vl3LiBb+jC1qhXCQS/CPC/GIQrK/ETYaaWED8cL4g2GcMc+c3xqzJJCadQS6EMHo
TujaTqFqBxOZd8+5B8YvPtBiV32GCgcCd7gK3EjU6jTIVtsyb+Pv0e92csKKI2x9
1TXsnjg9OyMrevRBPqffd33bff4UpvGh8QpGmC7E7+wqVpDv5EgqiLf4Nx6pUP1d
qw+wkJbMZmqdE9f2hnMqx9l1/6TA7JylX1/CW7Y704iPVQWD5H2BknanhnSFBtXK
YdFMvQwsfharB6LshpKsyiIgjTXyCUoQpqgPMQ7jGDFFBQpTtXBbfUUKPOK1UB5r
4ryCL51bx4tGAWGnJJkjBrIX92HAQHa8dJvxGGthenPAjdNWQQkrtJDettov+Siq
4vYiTqK6e/vQLwIZNhz2wYN9Fphgpaf+tFgd7aAaZ/uMqTdBgzIK9ZNHs7daSVBQ
ESNSiUfYYq4xghGqTose/2s1MY2Lq2oIB28XqWIINeTxN0rnlfKAeLvvW7is+UDn
bUgaODKLKTCJRkjFxla8d8iZ17TufA4lbzf1ePF3dGmKFJQWA6FmW+R2Et24BWWj
kKMKZOLJj0OuGjfQuAwrl0y1qFmupLyof5qrpEemgKTuPddHdyzScaIbnp4AV4TK
qaqikvHhFDZbmDkEVsKXKBDFxW6Yjc4e9OHxRVSzn5Dv5U+6OfW/PliMcTkXF5H8
WCFyEptXu12nMEbP1rlDwjH+jqTkfCmOdrqsGuMXVdokybabSu5sgXdiUE2k46Mc
O0SQkf5jO89JExYmHvd7dzWc5+/VBM1N+ezbWXoe29xtwhNgexGUuF8W0TLpjt8H
mJ3exl/zc7w7gPP3Z07xK3LdoezbqZHr1sccm+42dc/53g6/kUgQReN+ylpMFhnd
AiferAgfiVFONxcqvDSBBFotqZpovTBSHQZC/qso094I7I3uAUBkcFXDI7+d8p/M
sgjwfkjLudBnEjaojLVF81npwV3b4krUs8DRI+kwhkQ4ZzgVdTxKA9fVoo2U+osT
zFw1VsBvbIx+ZBMDgnINAU/3voYGVbA+PRb0LKmQI7Ptlw7+diuPX7Z4dR4HX+xk
n7a7KMBBZwET6cy7It+oesVF0z9iLmyhQxIMFqBgExw6UV7NvO6tMaNUKZqa2CH0
ReoBGPGQRM/APNi9cKJGKo5Y5FVoTWO3FxATN8hSwRGFaxR0umbddKfNpkOj9uF8
WqtJCd6V53ehd0Iz5j8qVblDo1BFAYwp6ZvCF6Pumq70LdtsHZFku1BXeVNRBY6o
MGxkSBstrShhSsPNXrsyMTTJT5ykRDOipy++kz5HTpFcxz497dJvokNXfYA/xQ3e
Uo+Ftop9bhNxRUgKUFJoaYdKAlgef7gXsMz+WLOXyMjeRt6FhG6RFoKhEzUtVrCt
7n8JrJukthRkgoMfRU+2aJ/oXTbCIbSNHILeaAzOpLBYcKdEcxtqyBPZz8FobFBX
W6pN8DIXuPSfL6H2b3RSgaQecbATUjkTOF5cnXUVmUDqT2OWyP+zpBjXbIbFL1Np
UkM/S3Svf8+33TllBzHafIOdDD2yquibdX+VMdAD6hWfXLGxJGNmvUy0+9PTodD+
f3aizYYPZAHIesn2RGii3vykXt/9g440wGR/b+dFh0Ki/D2YJLwYIhnS0B0Wuyz3
WncI8ZxCwyYmrNaPPcjNFRIxyVA3fxXFxYVvYMQtGlah8wyyVkKekPXSl2hFCwvh
YggRz+rbo7r+/HpH0+O7IIE5qf9sqFrxuvdfuc4oNY2VZHyB1Zyh2eH1Ox+bZu/I
/aCMPBYnndkuFiCMUQ26k9gy8nzbe7Hz4Lz4+NG/XaF0ja7X44wNnmfcNUC6+/rG
YubkTVjrXZ2u6Ktw0GHJH2fIi+P2etD1rAJRp3g6Va6yxYw2lsTqBHBkPxctKRsN
RzVFDRRHVol1XY2s0T3EYAd46I6Q6jCnOZIb1fiL49sAnUPuSvRJdvynf4xJP8T1
KFvG7lWjvZhwfkTGdmk/txLVsg1qcLIAUW/OazJPKe4jJRFjDQExfYwDiA+HmhAD
w99ggpElJYyphMHlN6ZJh5aa4bLTZsg1jgWawa3xwWkXDaeK0sSAmiw7MoI4pNuM
h1OpYjWt+5hbVXb5LTZcE7BCJRw8K95sanI26C0Ar6AMSsrPCqoO+Fxx21zD+ek8
VUtvKGOZmuKztiATlNNIW/sVRKjpHJJIFmzZ2BgaIofYSzSV7ZThchcLtA3IclrL
jGlWOgbz9kqtoujUeGfwoh8C8GHt5qCE2ETPEEnK9roSr5nBfDkGZSBe/vJqTEjY
ElDkvR+sWkdrnpNknt7EbjZ5tEKNXOgjdlb3dt/t+TSEw7Y0n/NuWidzuJiOnoQA
btxgeSpAZuFnvBdcwSddEcPsIq5dT+ee9jyhQM6N96nEdrQt2R2QvyL+o9qdzm+d
ni/JVpkozIMPnWNnSVGqqjeYRIafdHkHDOqAksZj7vFu2CIS6CktKDHICbP3WGfA
Xd4Oi2DqTE0bbCuKJxrK9UyU8gFNRfo22ymxmGhtKYvu7YEPc4GsWkfDwGiZm2r/
VhNBOpAuSy/Ku9aCPgxcBvwq0mNfUkEFKnfJCNQPI4tpiSZ9BIHnV+EK9hLH+uqy
trWglpz0UWojEjwa9QEuLES7Dt/IvgmMQIgj7wLPJD8j37sAzL3BPLM7/gwsGulu
70lesyxYf9rDGYKoJM20qM00jPf7X6IcLGcmR7KVkZWGQBZXc5UeqvPu8NwvMZHN
QahwMnen/NNWvzOXlVV7iw8CaG8sHSib87xqUfU8gT8T1QLBGlksmP+shUNv0p8e
9sUqL6h6fI00UlsGMXuQGNQqjaWOLrAWVfUPVj7915dd1u9M3j63lT0B0iCVuWLs
rgYH0hUANo6UR7NG5f5tGCzsNaWVGEdGs1c8uBdBEirvvW4j43Po9EQIS61GQQ6t
hLfYxPJzkkeFh+RosWA6gS5HTR0C7bBkKNTm6d9l89+2+CIERQOdnuLUG6I4pEJu
iP67h5VfJF2OU7a5Y+QBftjGx4XIDnkEtdMwifjDmzNiao8PjIfLmhoyGDx/u8VO
V2QsOnr4RboZ4R0aAbeZMJ74NWuQcqPpvxH+vPwfZr2JgPXKCZxldn9HG8lSm/Dg
+hQYRNYSgSaxq+IHdtszB68U3h9j2fYj/RYOS82h7+vXQKTie0EuASRDP9VNjYyu
8AkAA0QoTVCl6Td8DuF9FpToot8q9scj0n9J3ige1N9f7LoXWYy9hJCGLXGYsKWd
LItXl8522p6RrV7BXNHpGQ/loFUONYepBUKdmDdj2r1el42TGm8Ovvg8m81pcROJ
nXEmhzl9AkDFpObnCLKXHfEml4n0CiypcTs+IP0kduIb0AvgXK/QtHHoQOtGzx5b
k+MPpeTFnMWewZpqPlvC9bzsa+Vnq8uL7W0E2wBmyDRpmfn0B8h8It1xQEYsnUli
zuu6VmqMpYxn6qmf2ADF0bRgiaFF7oxn0AdmtWgRiRq1/nCzOYiST8mQdO+hT8zN
Y3qMTUx78vgoeWCVStugQ7eCFbcQV7BFt1bHC8MWf5ebGGNLx6oL3WeHYWZJFNvs
yXYoZdn048xexjfofzAudTZU+I2nfG9rdbtZXiORq2SYa0PqnqoIMqPGSc/QA4kT
07ESR5NsPpxAxm5TKTrXAD5Es6UE/9MYVUqpF5Ne5T67QcwoozXx9WVtPKsTQ5sX
2Fn1IlAmdnEiPPCLXlG9tpVnxXOzhNkcfxnlRpVAFQkblIyw7yr1rWvQtkx+Yyeg
EHoZmO7gPEwtKL5U9x7m054/Fy1ljNKrKhK3dTCqz9lFq51Ejfl+rq91JzXpSoLu
oZH3R+B1u0IV1W0pFXudsusCKR5UpX+RnOssq4IJSekobIlhnAH/ga4WTaLnYwdQ
2+Pwh682QC+S+whvE/3XjFfsJE1IsdmGeXtlXBCfvgBL8fmOYkhYSL5oqV0269qC
JchCukVukSMG4VHe3jeE/Vr5/GMfa2f15WuafswC92H0Nf0vO+OPOFHDvQXqlNk3
dcAHROsMMvj4Lou2C6w7INie2H3VhLmAINLppY/O3SKd5nncXaEMQEpRwnV77JPo
YPi0X6/28144iUz6p4PZiJ+ERnFGhDEQAGfMylavVG5BDycq6iw3TBqgY7nxl/sI
G0StRk825yxy8i78F7XDJBS8xdOw7PNK3s9QOnBUMfT8NVbUfjddfMjryfk7Ygj7
NUbiRf6xRZlRswSCJVJIEFQsof7It47ssRnGcB/yle/6Nc3a2uhKfYWLiovCSX/m
YbNltRzRfgfSnoORMwaYWOaH/yO0+p+fvPjMPUuXSkJSDpz5VwCUJcNx/WX7cDnf
+FWhkqWO0ROwezmkaOCvDxiHnelP2xqsTfeqbRdd3mVBPlXZct3y/NiZy3D/EIfL
9Lb6MLxpETyhron/lA+u0KE/J/FPCadWc3m1IDLOaXqT0nJslrxeGf2taYZGjDwb
zmN7GDWIj1NjD+u3dqL1nU8IE2XEekcnPKr/gMmVdBZshon2jiViMfg+i64h8ygU
jt2YG1mFzVKanrFzZBOs5shC/UZL1vgkGkdZDC3JGjB1QZc8N8fCWZDMsu6TWq4B
zJhx/VMHce2Rsha0ILi8xDiPAJJCcJyYuhq7JbLkYOfDiN9Y/cQvntOT16JhGKSl
ke1rzf9txUDk85QfR6N1DAHi7qXZJ3K9LubAIfXY/TIppKMdre1sMpOcH4JRwyGR
gGqCscCfQX3kX0WK8QyyP0OiN/YQ39YDxY+7oZTu407nYq7YobpbV8tUKL3mehF8
Kc15LAeADqigNTol9r7ht95zGrSWv0JILuKgynIJbR8H1dRq0ixbWfw5/hPp9m5n
nq7oE5Ku/5YNM/QWM947NSrHKdhbOixa1AzO4x3hdUta+fSX595+7O01vO68Tls2
hDg5cJQzZHMxxwyPBxdKPIW25POZv4DPod4Gu7SM5a/A+vo9jWxcQK4B1cYr2QNX
GHDChqKmI92Y+QVVNpkkWZchyDJrS30HPxfp4667fTNMWpzfwYzqSOMC61BJaFt2
03ZSNlwJJk/GHarkrtl79vSo6irHoO7pRC+GSmGnEdvCJVosIygtFiERmqefxbYC
Rms0nMTHjPNWpPu3zobeDXeX+NyYdHaWEDbxbMukOaZBhfNWse+2A75Sp/Q0bXQm
2rkBB8/6G/pgPsFsmAcEQhdOmuVCiofMnEehhkqriLVGSWA5Y/N/0JKPpDX+xSQM
r2phfacsLxmKgwPZDWcnUODE8pgA8FQgo1A3f3M4wxIBVYgTO6hsRWfdEK3jXYBn
czHa0ol8QyiJaBQOktzIqK8G4r+2pGgd0dadwszrju+/fqcW+Qh7MnQ/pOpXrDGS
f3840xYHrTm7wq1u7sKPgyLUggOUfqpWMy/afKJ9YwrUN4Ik2WJma6NGDrak1sOe
ZhmEUw9ObzpOjSkreFTsmfMqf7TbaUpSQ71iN7ami8Qa9YFOvs4OKFDbDDBt2kyW
mItyM1tMgsoXxnRyzm+zvQJA1WVfU+lPPdurr2EhUhBpGlrMwLS2yFdtn6EhBuCr
I3sYwCU2ZlJ4sZrD7jL2Le4XWmg+9PEjw6SYR9Ut9Bizlw+tz4nhq+wjqjLMeNCQ
21O0aNxg+ofxk6z34wmrE2Cx0B540OfyZRg213mBmdoFp4cGBBqdf3NDIOHaOL5q
n2Oitx4PTSV00qyOWcnzarleMFw43ZyyxRBeveIDz4bb/dqb1n+sJSFqdSloGwCL
/dYSVWgWTXanbRJzXQa+HB/azCFjQFdgD1FD+kUS1e2JxDvzO5EsQX3qtnU0Y9u6
GwpElUtE+ao6bR0E5rfRwaUz6QII4FP5qF3kw2xdrTxl5BRA9GeasM7z/7zDx9y0
pE14TlN28zCsrhc0MpAwTOakwD8mrmVpsoolPWscZAtnGowuPVpA9CevRx83Wqjy
ICkF/VQxi+ORsKI0T93W0PTGmvS9d4hTvWD+xC2hsXYLALsYu85Pp8ccA8en+lqc
ZmLYAYBsitSyrwoJBxbJTzCthbmH4uWJpBoRmG21xsKFU5jXyJxXfKPAQmt7EuPB
NMB2BArpYaELSCVHt6jYST8r1SodFFrheG8lEgesATjxWYgHe1ujAFucsSvQRDeQ
Pa+k5eTzg5xLtoo7h7Ik77PrbByu9S4WaJAffvxwyo41wu/VPgAdKLodgZsFZ5ai
PgT7SHJwkwNhoNE8b4hn64KL/3b7CjN3X9Bp1LULuQVoev3A7jTC81VguXb+2tCM
M773SORRgsdQNYGmxaZpy6j8aVOu5i4oUbtl23T6aA0BOLd7gB5t/YtbYr3ci6Sr
+xiB11k31aHaXNVi6BTF95XyHqZNRqD8YyB3iNrmN8hCS2KgE0kbBpqkKpvkJdyO
tS2+aIQYAS3UEGjLIXwSKvKoOSFDfUGSyhI+0LlH9p27lFh+OoIPSClxLhdc8Qq5
Q0fGTKmVK+ah2sQRjtRt1ZEtDttlIhIPhJ97tCgwg53NP+xzwMhE3i/bkNSlp53W
yfvz3mmLPSqdvTuhkkjIzy65RY901r1Yo9lTB+zwZBvtLYX7L70rh5BmmrakcSEE
eCyRlmBgY6pC9vcHxbSVxPEinNUGNIcb79ZDH7yXHRkeWx7oOTfbwEvUam6mfZw7
QTHZejP+4KPZSc48aJeXrNjdMIU+3sbu5ZjHkDgEc1XmgGXF78Y6hQDd8XOxbFek
oewNGRePILmGRiD7sfuDbyIQ3eQ6lxEuP8oWSZOBt9oxL5ouzDMgrUP/gro8KgRL
b+zSpziN1FE7Ya7eU7dXfGomzLSly0VL3QeT0brebVrNIV/llhAsQ5opK5OBaqmK
YVr8N07tSg+lWSYqr51NX4xkJm2BCtnAR1Zg9KynReRz2dMCU/+2svgGGGK0cH62
Hyo9TWO67EPCDJFUECgQii3LtGhMjbkjcbOO+JcPEXARijdKTAtNKQOsRovmtUQM
GXZ4jmr5DPZtYoliXD6O4TVUrqQYtWnS04G5GfiZBD1gLA/RDhNFJ+QhpFrPDnD8
SMlA2a9ZAPZExHGId/D43D9K3pGEVlFlXTk9oaFF1jbXSP2G8yaUOqKtEult4vl+
WBTp/H8mW6ow9NkYQD9wjCvEYfFrt9GDItQJr1RcBzw1V2GdytvJ923eAnmABam1
ZATWh/OA1E3Fvb8h0SKtLSAzuqFcAqiV+xU/ORBkZdpuKDfPxWB8ZEK/6YZSJHhQ
p2K3fUSPu01p7mGulCik6O1h/hkrca5NGObzw7H1FFIuW1RcBHelJ/ryRGhYgpI9
L3ioE6tghaG3oS2xI1F1pZhBvnGLs9uqZT3OQe4bYuyx7d6X94+4YafZZ2qh3MY+
1S1oXp+66agmWp4/jqUyEqQ752zkdq+DGuWvP9/m5RVUJkaomJR3hEyHz/b0dLLX
14DVhptHz0FzrSZBdQMlHmUD9g70v1leJTWlJcvnNL31S+GxKj/uls5exVbglU78
f5Maz3APzGLbgDMhVpbkVe9JIWuesayBaKml75GjmnRU8WQmLraqa+NAP1LfwMuy
CAn2N/7VI6HBCU+H2HiK8uWeSBRqDbA6tKt/w6bbUwTDNC0DvSc8Wga3UVYAgDsC
1ac2EytyiM7gvEeSR5qDK+sZ17DZpltRP2XoeDJhCRrHe7yaT+TaUsAvd8jSiZLU
jJyraCPn5lHgj0kBPu/WtpxW6UpggZ0vTezBFyZ5B25P/VV+2BKebcOoQc6QbHaW
OmTIuU6kTy5ZXqnh7IQQDi/sHa/eK6kHOL0rAMK6WOE4hxW+t+6N8urYLzscb3TX
ewz6ErgmQ+5RSRCDoPFWjz6qaMELOB/VYI+1XJ0A1IQlRNcpF3Zp+hztcPanHU0w
9pknEC5IefDUkOy3guKT+JF0Mz2Q8Wl2IyHvySbI1ebbzYQx2Fh51pWbj+ISf58N
i4JyhEuRqIhcwIDLKWxvoiuMP0Zvbt3Sgn1HWV+cwuNODecbGhASWtAt+//4runQ
Gfdsq2/CkVcdcxULtoRomeYc8Il9zJkan0V1iF3GjwKV0DuWjdFyXMlZKPKUnZ3r
IDzWdnZiJc81aO1wxii9p1YxUYoRcDSW1xKWVtYxF+h6GQWJXSDo3DUIbkivHTOb
4QhDAJ1VJ6zZYvkh6MYNrNq1Nrdvrl2YHNVH+Et+Nr0St0ZP86gmJyaV+w/bErHU
dQ8HOdUzg8ipE0WEE51Eoaa07BFImxm8fPPODFdPrZ6GmLboyAxumQXJqsNQt1jP
vBvNQPAN+7o7IlviFa9qe6Vst57Z9RHqVk9Dov/7YElXRCqf3gqsvBIFMXhhTMqh
tZn1ht6mLPAZ6BJvlntKKLsJEszjqRNGy1D2s9K4TiyDKUPx7Ig002+8xAtBRKfb
PinsiYw8a68sUhWorJgbI4mGoujQKT/7QtfiyeaaaEsLZub0QkR/FNM+nwOJOV2R
AIINBpCVjYw7JbRpB9g6qFhlgjY0IY5lTGg24O1ingA7wZSLIRR5uH1GSxDTEYc/
pogV/Y9ukWyn8u8BQqvJmytaRrWaxBcnVYyLDgQvMwtpEQ09/Osu9NwTWxw+BGTk
zGUkbu5iFdueKiEnlqrF8QH8JZT7GVXNHOMpiLbB9IvZsvJRpt/6NjACeiXIiL1k
gd7qdMutyTwbI09ZqOzPNgwzlDgjzDOUTlS2KQzWab/2YG0myMolHVvlztNHO44z
sWLAXANRC6BVKy9wf1wzb/SL8/H8X5oiUEYZcNnEZnaFCR0NU/h4PwB6eITT3rqv
WZg+xhOixlFZZKqd6j6IkeJezz/adUO2r5caLmBMf9bkNISbhI1mXXa1ICZoPOzZ
I27c8Bf3Rt2jbG1RBBiRK9u9Yjzl10Ky0neE2a/NyftGZSVdv/FGnQzME13NrJNY
IGspVB0aPDOp5fY2XncmqheUWBuHt8CBohOMh2219QQxzpupTfEEi1QKZ7ergDEt
YtLcV78PuXMWnvcBMkIQOPdN7EiIQ+Dk6XycHCMWslVXLp4pmboKkuPynNqz5fOi
WOq6Zr+L98TCTs3psMaZOFnwn2mVIv4K4kuI6fivuD5bOgd55JHuQof+CRVFA95i
soo9Ewv6sg6ZYDqPvlm87oxqy64FZ+3G2hrra5SlYJ1alnXKq2U3cPMcZPXS6jr6
D/OfZZaWoR3bEfdD/PGWec06r7e8gEh6OgYWCcqiPVSbjNgd2t966LZ6vwTDXE65
iJp5CiUUwITOqu7kwg2XLFKOUFIKsvSKysMWKsC41oF564xjm6ETHmQSuoaDN3hp
rV6X8GSpQPb0zcwBXulO9SzSuDz7+fOGhrdsN/Zjn8HIy0DJijiIDaW0y7ZycUHC
xOwcYLtFTDbIn+HeMqQ9TIdUINYSeobKQDSmV0u+Nkpp20LyDCLXmd3+NJNyd9bC
bDZbwK7GbUODzLZ2mMkvv1G6KfNW5akVXZL1pwcZ5jXAls+6IaU8UKWl8Iw3pUgR
ktSxBF+wN4vi5W7ojp6BVbG+K/5fD81NWoVds8WG7qnrD1RfPidfmk9paKlYAU85
kg7kV48anO2Umufdu7vB/uJRfMmJ26xX1WcVLnjX5O8AhdoHanUDLEi9yGMWmYlO
QQJ5rekGmZL2c8rxY6M1wBPDFcr8yyCLPxYAJ/bLOBSbkknvyHXLl5Jfmb1La/+x
0hpP8u3vWHp3HBvRQItX0mrfwT7cecQoJUxozjazdRSpLq+MSkQ755DXWqkquvD3
FuayWROQ8qHAX71KkcD80PhGRtBxqZ8LC51E1MHW156VFZPtavLI6PCLGCiVL0xY
hJhYl0Ikk+YVdSe+y+1qAB2JsLgtWBzlGABOTq24uz45YZBPUHiRdOfBUXUTm9g9
NYsUrZt57idSfExqZLkOUpMl+Xao7N4qzKHrDi0/6iiL8FjEI3JnEKrZhlGNC/iQ
Gwa/gcTvEHz7sSlkZrQIEE2jJWWENQYpEtORzrGTXX6FyC/PHJJcNrfQe1KO10Hu
Qawpv6NzYrm0GelApoE50CDyqRnDOecmMdySdnSfu6Lf21Lf/knCU+2SSgInOGax
TP2uanxRo3JLbe6VuzyUOiRq6PSZlfc5MMhJ5i3PNiNQRewIDdXNISEH/VCOb9il
5/2Ent7K0l2UIBcHE4bIXVrQSs6gj6sZyojgY6SGcCzokTXkiTLgSg0XcdE74YTW
4vqNEwVENq1airhRF+AG+NpHQvW5nLyK26HdZRJEy29/Lf6IazOlVqM88O8gwCwS
/kPCn5U/MzEj1VnRbbHBau3/VEAoCUOLcRd0/RTSGGpE9dsqqFm4FppD+lmiREO1
2J9GAsxcT7TSyAJP1suub00JSo3E5EDxzBXfm9iSHkaOhwq7M2b5lFP0aMZLQtcb
TkCe5G1YszUbpXziPmciB67/lj4uAH2PbgUXnnVCQ5rt17RsvLRhPy3JYlpRDRov
54gFHVsjfDkTitB7fPGvU/mFw7wbHvzYyH9rQsk9uhH5kbEJUU0Ex17JDBExcO9f
ae48tIe9kDteJecCuNiB1z061hGwe1sX6HmumRbL5N2LLe/lGacK/rd0SUkBErTO
01mdhQ9wLYtaTvt2Ya4vsDryK8Ov2EKQjPtmCflUdK4m2wOuM/1P1mpzsoIdpjnn
DmuGqRkb25Tl5EVxz8Rk62PEtHGHUoMph2C76BqSy608DoyTOTRzQmE5HzLy2oOl
s3nDBmrbw+Nm7cA8T9PMM6AMiGMzf7dO6O6nmwPynKiGoaqQqcZsGLdEIkSHDJ43
vxLwj7CkaP0Ly+Cen656KwAw1inbHIpj9iNJdjoa0LckWxJhMU1lq4QTW+ZD3H3s
YT+ubsVpcBGcSS3JnCqiHNj/+7Z3f9bjIZuTjRZKJI11W9cpEYBMS7mmuqJqGpqc
EQPmb4vp37xx4V5lybzEDCzEAS9jSKj3rOxa0Xc/nXpdqFZCWmM5pxUovkxNehr+
eX7WEwADmxYVQegl14BV08LCTSSx7YX2aCZbcZjWlXxSWtqXi40pqwkL+QeU7z+R
BLlJUjxnmymGPn4MtwLjkzagt4QcCz2fycSiyAgpKq060TzZCIhXe7YQaY7Ivq48
oUQdwARhJrP1TqqEQbB/uAV6fZKWcNkw/lH/veOIIKiYqJvRa2jdLo2+9J6n0/s1
KyhXDswyEDsuBxu3lA+h02H+seapMOWT3fmnmfQfwRpMj/c51iw/F6lLr6QIwwkg
eQsbP3/kGwNThJ/3FjXA/QHISsdlipi4qTbvYGd3hME9qYMxS6+1vv04zq7HKdTU
CDYCQou0NeLtzuGgbLfVkGDKTcW43kVrU6I94vKf0JnqvCPJlufzSM9f4cdXcJE4
UY3Acm81A6pI2YMkYie38nEyANgh/3E+uDaET+kg6xkhCOqrzXrC76BBUTSANa30
JwodqjXEfSamcGyHqhkD10LZVD7w+OeN1FQgbe6funsdGWhdNI7SsRIsjGz+vpl3
2V/Fb7+pu2KxBJrZ/tNJ1td6vpv6QJseKspBoCDbOcAygOWNyObc9fehKJ7BGpQb
AfzD/N9wGj8Iq3M5AFnBn9maz5ddaHQryhp5sq0TQyj1sEPLyUwNax8e2wmmzwI0
vKOI3ezSzW0GtxI8Io+5NgyxWhAxtdfwTtx/Rhe9SZo9XmnRo3biRJdxjqPh3ZxR
IaCXEOfXXey/uV47heElp8fZsTVgmjepbDnsiiZbIy2Jf14u6+lCEfH5Gv3xmQiF
6K4v9FfgH8hEawvD1eUDJsSM/qnLKBJPAhuoBSGBUze6Mv8+/G3ffYIJk55TBMD+
amDQxEHbf4gFJbDUbN1G3W6KnEUFH3l8Ct7gR/5vu1mN13eclgQ219eZuAFGNPDp
EiNAYeuwP+ADQBt/DQkKtNuh6W7gQtUv/KggNR5FPmogwUE+VBi1Dl9WdYRI4UFh
uDOtTr01wCO+5fd/hxjLb16cg/o829F6aMHdzIdf4EEHLnXzq0Mr0Xsp1K9kdkko
ZahseUtiXRHPDJdmBYGnShmXm3qIIF8vZW8YHiGUoQM+lQySUGT3Lx0yUk1kXEq/
DspMiWLzdCQ8N3zrz2OJ+0E32Lc3Xm73/nncfIP9K05fFd3uP/3Ps2t4boBY+6Fm
Xw64M3/ve8r9DucybGzdtp37+wlgydR1KS9QcfAUXai3Ea4nOa/b6+mJ2b3CRk0i
pYp7f3Y5Rj4cSthQ9bcjJ70IrgL/7ob6Zx0cUerZTvVcVVH5RgYezo0/dNNia1E4
na6tjy0Koj394n2P8htq9IUlkgBb8LXhh/9/oIokkOwFzRU2iZw20nZtvduVGpBi
QCM8O8lyCECsNBji+6aDcqI4DaOEMrCoOm7ZIz10iDdBdENoEZWxZBjxt3+Ag2lt
vtysQA0rBQH+8MhoB8Y+kScWi/wr7G0phO3PJMC2INgm/EmbW8/Z6yePhgiSb1Ca
G73goiaxRQngMbNbbt2U03PjWPxkCwMkkdNwWeFW0coz+qHRiAWsHFh49wYCTiva
q4HQGFIDnoq9GL43UrtHMYdDG0v5BbnSOMh+zAkocjV9uweO8/RkNPS3JGqvhCNM
dBaqZoCY7Oymp4yQMFyx1ErimAeTkaKym1kYgSE1Pyr8vHlIzeeTpQp5GjqUXpdb
mo266COUI1u5kfz/TUHZsOS8P0vNMww/Mi+4KIGC2u7bcRO/EIZ0vYmMPB9SJyrD
cI3jXJ4xPVlbvou9jkqgXNX9dxXoFXafS/r7jPN8KTinRvoOeYNvyZ2De9qfGK69
ZasZt33PEhKo5smOdOZhwjIeYpCkhC5jrmeN6wQAN1AR92+9RstKdwXgx0Ab+Jxw
ml0Lw4tG6fbbb4Jja0mOVtBhdpNlNQ5vDC87ZUUf0cqPzWEIUXzsnc/5ElXnLyKD
J+c4s8m9g7/rjMW5Zar9e7HyVyzamKpPvyKalUBjrhihxeuyKcl3G/VzKFVWh2m/
gXWHtVufprSJ1SQbwEVJD2jhfrR6wbMzjCtTHjOtwiGuVEGv/KDZf1cJcBGqLWky
RXR/u2/4awF1ZlJQf2rKpF9zfRisTPICsbrBxSN6ZVE3pmqG2YxM//luLQUKrq9F
ioinCz6fez/NLTXE+KxcvOZshbxo0kz64GYeuZnhsWdcGN/vJev2F+mrFtuyOvrt
wSVAQnl/iNugVkqDX+GxboXdy+UuN1ZyX4eAxrP5WyNcl53GNxXD80ZGCWA1teWD
5tUOeAkJX2QbBk3GqCSiGd+Pauw6Gj7nWbSWK1JRyjSFVoKkx7+YVkge1p5KwP0c
YuXqkCQfQnIpTQQWcrhbEnZ3arFMQvlnmvTWY4N9s99E/0sEgN+sX7UuLxIZ0Fy9
5W5AJ6CNZuSwDp/H6HLpoG3a54t+tTHZI2exGGT91tZnKMfrj+P1LuvrAbPb/THr
R5LRu/spfoIXESQtjiwbRq1rYemrOdhfBx0bAizDZNzCjhzWRi6xptEHN0CAsxlz
Jd9p69QS3pei7mN1UXRU3rEpmTKeTX4hLUFIGa7pYR1mcpq9tIcpgAAm7rkVkGTu
zlESuHtTFJQBJHMC7PxbqA9ssK7gZz20FuUcCNlqhBE5UrtDu/8bUoA5saDasZVj
N5csHHdbBwzyxEjEzrgJ+Z0qlfudi2McFVwmDTUYKTKzFA7Q1V0xoTZuAqyz8OhT
GxP9hzPL4egcJJCvVnoHNOF4+/h2e4/SfMFACQxt1U3BcRnBFBD0M0TZYORwlLpr
agyj4HeMbou0pJpwFZdhziz13lO0TR9H659JKMtaORT6i4bXl6jxKm23WcBgeH0a
xTmS0VtAa5+C2GF/kULngj7W74BdrbxENblS8t5wAvuPFPiHz9i4dJslPizoVPCy
No4+3tygyaz2/J9tbMvm3/GVzxlJa4vkst31gnG3tNJW65iwQ4UbjytSdQE3EoKx
gMBbXIIWI8NiHgC7u4ya3nxBixJax6ssv0jnXNFWltBrK49uoXLPJkGw8mHWzqP1
oXfTEuB7f6nWPoiwFxE3/oa6aAWaaPLeWgJwSR3I6zRtF+WcE7tg6knhIF3SVL9Y
kMZJuZxbt6geGiMerc3eTJ9Ybecb0cMym+oTIdVr2v9NXrXmACkpdq1yeRFIJegV
f0FHoQBN4xJxZ/woVaHvun5jKwiYOK7x3s0LjDPWezeYSmUe7KvmVJMX0R5HAp2+
S1OE/gSeBr7da/KTGuJr660HGJ9MPIkPtInJO0Gazf+OxrvcWJ6lzt3kOCwAkLz4
46ENZZBNLOVSu6VZHNKKhmxsLhdGmmDSkVN2dDeXHUWZE1jOOeIfOn697fdetZSi
MaQXBMD3aivTsAvxCVixw+OT1a3Bzlx6GWCIqnC/3ttQuiialoAzO+G1qv+QpSG2
KvHNgPpf+T/maFwHB5PhXJPXXCp+CYUcd0Zq711prT9V6YTX3V24MNJnRYXSfmwn
o7kwLIjbpfkWjW1OlXWktHTLUxS8Aox4wZZyEFvHtn9khBjLboDGMUqM4oQbFAoy
Feso+8+mZyMDjmm79QjtAlfTuEvZvL8/jaap/Au6+XdAKi0zElYWP81QQ4nFg8/a
fU0qtNTE83S7kr4L08+n+SqFwd61aDvCXYLBlB0x7HdWbhJdzonrPTXEAN7LHWA4
ZY68FDcsjhwLuLB4XGs7n/JGmHYwht+Zt4KWrK/vCQ1uhRm77g4e4EJIqqVkDVnC
9qi0uFbaRbp6LtfkPY7iLxeFvDkwSEK234CEbOMnWTU+EU4ZjBJdIUa+R6dzZbyF
3c+Elz/TGH0kbM77kxbu5FNuc4nc9WDj6DJK09YL/GIfU7n0wj5fqnmuHRcrBix/
uBQIy4WkkdOug4HXcK3/8oHz6IGAaWKFlWEW3YJeVXEqQj3DcHKrJ2awGiasxbv6
caKKj4ZTC9NEaJiUAmv8mN3gvOUkQn1fw09wq9AfzQylmY5MxsSCadzKe1L7Ja5k
oE0j/KxCEiERuWHDybD9F4mlXQG3WxpJObdQstpTH2Q+yeiGJbYhBPShTm57GcTY
OkgyLHomoGr4oslhc/wcIMd0bRc/JCz+B4U3NCzNjVIPINPcrIs+MMOylJhNEpRr
Sw/nua0/harh3zLPQbutRwiqcnWkyik1XNAgHcNmdvAtCOOMk9xPYRmcie5OaWg+
I/j3Yv8kQvlWrkz+Kchriza9/8rV5pXwhTEEs3PZN/fYf/IXcb38oalyMEpVhB9I
ygluL684idLac3pfO6ZqSUXNsMMkk1Daze5NsYn8QXCApTahmT44VrAhYlLB8qBe
3sz+gAjodSXa7nGhZe2I69zBRLmxefwGRwVsf6PhAM3rS/lcUCM0zu8uj5xT3u0Q
4F3qbTk5opy8s41/rLXDKer5gHstkoqJBZduS6swLp0SDoyphrkQ2BtOVo1jICh2
HsOQYy+icYShlZ4albj15H7fXbQhjWShKD+hht7fmRzY4nCkQ4+rwDjLqpyhYAwf
oDF99m8gWonNjoFXdAxz5WCljziVzsrEN1NwkPxoFoY0V4eTpxrJQ7rO5Lb3JQG1
rIf9czCnUCnKsNj9iYc+tmFOq20f15lklVU0cF3mG9EaBNZODnOBbY9k135GzYdL
91sV8kUKPLLgzsyDr42+tW/YiYWWh7AuSEz0xuICYfb4AZkzUF2h5NmTpN4giMil
6eWktLkiJYbIDeWbV8fdv5083R+1g/4kIZwDFQsVTYNgfOyWG7kgBGMes9P6DCEA
lZ/pLSIoFOTNwFk3lJOAUvm9A2Yo0Pu2Yd7fIDp5i2/C7jRR5b+xibDSHjde3gv4
7oR0bqFiPYRxobxJMn/y6VxAcIHVd+KdA02lngWXBYbrGk66ByW83xOdBVa8kDQv
4NR9yRg6woOhlCGMR6UPpDeM6wFYieIGifXePOEwKBDZ+MWJNEZxq9vWRNQN2R9e
U2caaCSSJtDxlfBS3bGp1aWwZiXaF5EbvB/B8Tn7CDkgsb9FFdD5JHrhqrx29Iwc
4yeq7/jktj+Dj4rPIkzhErYH1x08VhsSodyyTZHshKnT6ig93ia0TUgnVF6RtDM2
olk/F/S5TNiRup+docwOmT9I29S/FUmxuojNfHzWL6khYf5iqP+Xc1fezJZjbAMx
ITrttjvEZJlsiHgF7PdY2ujKr+BFqq0lwz1tkclKba+yrb7sIeOmtk4DpMBoQ+ca
kPOpMXvcDkYPG5B5FWLB81IWJnVar1bBRUbMUPt4YXMxr5b8DZqk6To5zGD+zeVc
gzjnBjV0ULvw9EC5DpLAzb0vSgx43gi48pY3fluZVKuH0SpmEPrEt7aou5FGh7vu
iJK662HN3V11z23nq7Wi8vim+zm0gXqPnyfuFckN8+AsCQDNih+81qDBRjtwulSJ
StQHsU6bLXz9gsPzTqaqUUyJcuso0Mb5kkZFJ+myUZ897MPYit9cSXDuVTN8OK1H
19u/EehDzNCryw65xDfhS4yONrZHO/Y7NosXM0uhl05CYJuxbz3r7Zcnp4x7aEQQ
IxXRh1x60C9JmqQZcSmtD58MWpgbWFVB+rwK0MXqpDHS3VZ7dpjzzy5cuCjAG2Uy
s9Ghms/7SrlfXOv4ScJmx15kCx/lGkZbZncsSN6Bw2OhAgQdaOfQMC3oHD23aMht
kGHp4ZNZgSR7qb+t2Ar4Tm2AzLjJt2Ps4IAdAHx8XEomcxq0ykAyayfbKDhaG0Z6
ANzTs+M4g3+VxkoYEtCr1jKtBrB3bAAA4w2ii+wIC/eSZGnZDWJfLHGJA/qwMZU2
gFt81qpFjG7W3in2wk4OZO1ZIVK/O+sIn1k5N4CRVSV4fB7wJ2qZaq/C6GoH2hpI
BfKMF8bfrZ9UgitHQQPYvKF2n+s5S9FttUfDy2JPSezZuY1tny/vvUg+YHki5KSk
39hk0/NrdPZnmKudS8KmzuZEmnqqI63V5iXQnEhrcSmkp1If+Q+4EpR7Tf4nK+Ut
6c3Mnen6N8N6jXOLgKsWzkC9BDOFGXCFJtO4fpMWUE4Lv0Sj3sahDGeedbAdjefa
xcyivoc+N2Kde11NqpiOm5mXcR/nbd37wUL75vOzk8BCSF5PlFr2LzrSgQ9eNu2j
Uf+jqoPEEPzXxs00Mx/9UI3oKQPpsSadIeVoWKQgcLmxU56bXRRMATjO/C/TjeAf
BvY8Rtnqn3ZDbgb/8UzQoSSDqS70vbnQYHqEE4b1sTzPFnJMu80JftkHagBqySLe
EnokE7lQ3N8oCkfmDG0sywVVptgvSd/t5WMrtPqhZzPBiQZKzyEKOzi/lIdwiPxN
+2te7NWqYWlVk5D0nh1YM0wZ2WIIkGDGBCaC3D41/fexhsdRStC/s0X+H1ICom5j
9xVJJyOq0WWwVbCQSB2EgfwKYK9ftq3SVnTWEd2ziO0u+6VDitk+nlguRkpxM0wV
rca5lDs7/3tKCwSbdumK+aNxq2iyyGgrt9cG7XHo0DZ41f1KOS1aqURlwpMTT859
q3pyQffS3Z0Y64xoPt0/Rl0nlEl6Zm09LFHoMq36YNyEmrR1XDHErfrOqNR9pVVX
/U2pLcYlITbLaSnz2RC7+aByUqI+f3flxWbNbvoSCvJ7TU7GNZcvO4wpxm5jsgTF
2Xv91rrw/awQTCDXuRiz/B1Bmx3Ce0p6dmz9da27YPJ7rc5Eqom/O++FtVF16rbH
r/3lwQP8+ugqNC29siq3Oum22KHT0SuV7+kuyizFkjZptTIVIlrKVF2u/U9FesE4
UT86yHW5ypAukSLmNA1GTFevEpAk9Fwz/m04khvieuySNU297J9VzhOG7/nnYd6A
xlpSUz70FhkHw2efq3y01o7BrL45lvl1lNKqbtSZ2McmQBREiEpKo8MpJXSa/L/e
0QjpcmcRokgb0PDgdsAu/OUkJ9HG1y8rvkwOYjjWVmmWE7B3uOB8F7JvHU22kLPH
gsOnJLe3x2o+rUOzar50P5LcnVzpySw9/8wtW5oJ0KJJtUS+1EBXizUFMlo+0btI
TkD2clvfhRmFmQNlnA6tVbcB0fbfJnd2+G2/WuhmhShCCDWvKz8Ycq0ZnN360xBB
aZ5VtIczZe0RoaBNt3Sewq6KYwSHMXagnJy0L/W98t6KpmR2sdoUHlZK+kdQRGKh
G/qkugonrivBo9KPXKUOB7aHITi8SgK+uARVqMr6egvj4xDHDo1iQnUtKsNhLTva
nwAG2cg3xLXTScCxkiX/i7Lcy7+vYS/TB8o85At8ATNbjnUdOKh1W6boktTkVTK9
ps3qy2qgNShbAzBfP0UiI1BGo1kzVhjeRrjgXDRJtQqtL+gFv0uhR1i54YvcB4qS
G5giDBb0evrv12/1XeUQKwe3eDEuH8nLNUMuXKudAvvppXNuYuiVjOG7T3RcoZuh
UR2BXeUUlDF+N3OD0RSUW5cimdUG2h3llDBBBD9C4fqEfEyviPlLwOsWIqKxWUia
FOJAwfRv3BqBSbPRvTLIvCtSxlYxrXTFz5PpTTXgMu8aGKyQmUd1yoPn0yaVnz2c
F+eBSuG13zW/jEYI3khWPbz3WNYEGg1IyPZMyNbqSdqZpywSs7HsTBqpRECKUtF5
2U5xmWjs33lFRmlT5t2jp6mLJsf0seFjGTYS0sNEIZSAVcUTGQZS6EyUAemna0fq
FZPIjmUs5YqM5z9XjXZfojjAC8xRd49ouZuGrmWT1JYmjjG7mwyt0SdUz9ysnUiB
3mTAqKFBqONr4L8mTNMkZucs8uVvQ/AprngGceYt8dD77rSfEOf6GNP7m3dQbv/X
aBijPe3HPxdtK9cGeyxNE1Y6GB9mtDwgFQ+GbqJjzF2Fkxr31j9ZKm4mBTd21Qt6
Cbu4VsFQQ/5IAzYu+H2vCSa2fYltumWiNH3yufTjzYI94W0ceU2PvwQmXummdLq0
73R+Y7UWGSvMY+LCNDm92jMC0FAKmg74Jv3GSckPzLaJmP6p+pIvXBVQ5x+D76Xl
USyr2yLJ6SR6KTtJh2XtsPXNxoXxvovE1OAoTP3dvVtz9hyWRQf9P7xFvETchzsM
v8UsFId7Xf9Ot/9SNdkpwe/wN5sK0ANfAKPeeWMovg/GixA/Nh5DoFsaJxWR33cE
4Cz8VatVl0Xh08XQXXSKF2qw23pS5nzjumAoLa8CFQvxxSBHGzd1SXwrZA2g+imz
VGE8OYZAQDt9kxPG5QocN6sLQLngqjwTU7rTuOwN5/uf1hdi/OJJOcrGjSMNfYh8
H9I96MtoswiSEf2Eb6yigd8zwiGclgvt2xw7i0Z1jE7pU8By4Scp4BvLCDt94VDK
aKsL9XVIa/lPRQeJVcx4s3FAHYzahyg2Z5WOZP7gUtVVJJK4kKyqIvBuDnQwPBc3
BXRy8r2r0ZjsQ81G5HdXpwu+UwIbdET025J2ISunKTvWUTu9HknbEGS7gf78AQEP
Usi2XJN7NUadQilRF9kp96Wz/LvDPMuaJK2bhky9EQ0fR04k+PK7RPXQdsSahMoO
Auts26CRIj7qTZFUbdcRxRWQ0popbX0AIIVt1QwS/hxQX+PEjjHH6PxBFVlru0UF
jWO92AcJviSUZDK475y3tjaPcsZuCxHPKLy4Y23mxEhe+13ew2sUVH03AODMd1on
Al338NlUduxdu9Qbh/GCQVGVO/ztxPKv9lMX0o1i+ShEXpwz09tPmQeh/043R9Ja
7koShYX2f0Z2a0I6svZmovWfJXYXeKiE5uhXKgx8nJMqK4R1RKxy2Kzpztpa0wC/
bZ2WJEFFsWE/vdUj58M3uVyDgrIsB9ASqy66tlxgToXI4wP/ok77S0YwlfvuO2eq
M1P+jfUVHzE+QNw8wCeNT4/OcaNwmfJghd2cPHHksIksNaHpHXIVeqBJgbgRn4IE
JhgGbf39MB6Igpc0eiPr3/Q7MYTodWrLL+tkHnoBqSPlF8ZJxKOtSGw4N85PNTp7
TaRvKYHAHdXRb/Sk1YNoS7HPRr5D+e8rNoGi9c1hQd7j1JkHSNMJJeqLtS/3wIrc
KBJqbfXne/tUojPpE6kCZAK3Y8f31XuByMK39vvTWX8QKVxwAL0iijGSoYq67jKx
dG+izrNZfJArnC8eTg+V8YAdI13LFjNFCuCTIGZuppyT/d2zMhxtsBADVtVMP5Rs
sH3rxLNjHOSQEYmY3dTj3OX3JDksYI8oYHhr3l4LncTunmtj7Y5h2y+yLRcZJHon
dWkJKQ+6mra9G6UeJqOFJXa4Sr+qC7MPO4454gEkU19qsfoD7KUpMoB93cqBCfiO
OE8qBqZY7r8ExCON+l6YaJXG3r8ECnK8DnXi5GPZbLf3j2jYE7lUAY+yc/Bl4t5b
6ryX2+fcRHLKdgh5pf+m2Yh90xZCGhOdVVF31MIIk8xyz4YH88iNqXkznumuBYsS
kw4J1vs6usnxGBE5TmZfokqphCiAicxkUw41mXL8ViE9OsxB5sNCkPzen5y44nYC
KfO1HCtqqm1VgrKfQcrItCXEguxNfmbTJfWxNCE35m+DDbg0npck7vqEQZ0ULNp9
F4sXAwbiJn2tjZA2pKq6jtVQFvuadhkLBqxgaePdnpOIRkw7GYvZcFRmn53d6Vq2
MgEppiQ41BHMLOBZ1p3s8o/z/W5cp4sCJWpIlCv+88TIK0TtRkkld8qB4h4X9+jj
3OD7H8rTPBN8WRaZ115lblAWPejpvidIf5YuTYHmXVIbhibpVa9HOm8TSYzLIZOy
giQULGdmHtfV9+oRXVJ/K6BallMu2yY+T89M2YIriosfX4OhKXemxVmtyT0oWrVN
intwQZLVRbsFANhOqJV7164l6qmqqefqayD6c/+0wybfuaanbxzGKyJ5FnCVB37F
ss1g8uc+Nb6XJBQEQWxd9S6s/anY6ZZzDGrlE7JfYfIKAAS2j4C2JP+StatB2It8
F4Kd4vnWN55vhsJeflQDBJPp7big7OgTWL8TtRkteILLm5aNVM1aHSwlA/k/IitX
PaRuueIeYGi3k7IobKLzp5om61d8i6sPE9KMvXhyAE+WyL1QETb4glgISpG26FNj
llWiHlM/I0wBd5yZMmLnWipNgiRWs4/VcH/RNcgXRqiJlk487pcCQTeBc4eO6khr
Hx5mKsHrzVWSL+D9jTlRBbMzie/JVu4HLcykL/YEbOSRv82DuzaFeJyZXpe+wq25
KPzmno/fUk/VHL5AliTrBpgJ55UOCdieX+ZUDyaecgr9jSoEaAZ9e28JoXeGO6g9
+vpibeZxmc2OVOFhogdHg7LeNpepKb0napT8rsCeQsi4tJqi516S5DPBa8p7leyY
Iw61nCXdfAscz67xqC5oysDardYZBUGD4rbWN7C213fJjPuQ1oQMczyM35lhlbeD
I6XR9OEqg8WMgqbdID6rqmtJfkGwtcxDQf2GEuPhhw0qmPJMnKjCI5wnT/0eaPQT
O4DiTAzi7b5R29n74bMC4MfObkoCN39sSGA6fMPkkTuez3ZzVx1wKJBxw56yDnNz
q+lI4utsxYVR2dcP4nUDbwhPFdbRg5GAPumX/62HGE2G8TBPyD2W1geZxyoLAhHf
Pttsk0D7ykmpeIye9xrbLY4/dHmLUT+qqLbblHr8byMI/J+ajYmxwQmnum1mzsVm
T+4I1ETiZUNIZejFV+cyadELrjiU+xx6qjGTI4pusehOgHSfZN1NT/UQKUCamWes
YEvrW/wRylQ0NW7/bdpaXejBjS6FKhIwxpuFD/WiSC4YgRy712Ad7DgBTz5KZUgO
GtTALsgJj8ybLg5+AGtDj2FLvgnAvghXe3opQb0APvsTOYIgt1q2WDvQLdg/Q5uO
qPxNJHwOTPyxOl0AKofsP77Nn74v419RRfiBMcbxW44JWuT7HlpUBNArxiFNtuNL
HF40XMdGNoJdo7k496FKYoIACRjygaDu0PIOoNBhbb5AUsfuU7O+TNgHCToZuuu6
BB3MrfEXBIb3H3YrMbDBm/NnmI1BQa5O4c1yEzP9YoSLTZ3ud9HGS8Wao2wqpJLo
eDexDtAS08XbzhjkUhgkrX1wtpqaNXyangzPtR3Iq1Sxym8hgsrhlgho5/3CIW4Y
9MyCRosJIKUx3xoYJnaTQoFoeX8YqrtNjomMOj9NC8HMvHLruBGN0KODIrxGbriP
MkKrbldM9pAm/kkqFYHqwvf+ljwb/PVpsGNbTV/YRxRBq+MV0FVm3eHFV1B0kRSA
TsupN9puSh1tx9vZ/AtN1HEwAPU2Ce8gr0PirPYTFrqgwvdBxdq/idx4kvp/ckLg
6BQst8yM0jUqZSyXR0ascmPbbJMZjkMrqzKgmfEScLX2fzv16z5HgW+epQ0B3bac
qS01dkf06UV27u43KfAoujEZDstehnhQAWGA9Tt0uiCk1e7SlENtl8yDBLc4yQpu
UMVOurh7nrZKqnNs/KTBWB/AQ34mOUnVgnPmosF7nVeFkwMRxnEyTPdgTeOS5B3X
p/IK5BBqQ9Bf+7NA70DXAxbGxgltvLb18bD6C8fz1ci1EnGVq67Z5x27m1wagjrk
Gb48m9dgKyg8/R3jMiUKCoXb4xb+Bm1LUfDiX1SXpq8d+cCO7v8YVh07DQ+ddXTS
4XCEEhI62wppUlwUZQ6wbOlPBpnwIkpX/sQxeJljnZsvTdEHYtycDaLnG8kmV/rd
o/ss80BFZhUx1+pIPwlWCfSXBf/2fgNIyqbtyK/bHaMJpWFEJP3LMjggs+i5UKFP
zBPMXcUPmj/5DOtKINnFmuqndEU+flP+NmXzPA9x1kQIsLfFuKPegCviRNfcB+Wf
kDh9tO3wsCggDP8brTYK3g1N/daAzztzywSk8s+15bgX/fSplKd93OrVkInCMGPi
WK89vioU/2EEGgwHPa1Fio/z3QVHEl2Zx5gvz+7hYZo4fZfhX6fWZFdTvRkVc50O
Hn3QmpcdK/Gk+MSzVeqxH7vHMdx62rYHBbnXJZOJKrY/CN6eCRl+rJVd6eMZmP81
6ICLb2QF2RsaGep1CzMM1MbEHxAlIOTxuZtotb3HqXuwDuwWWxV3fYH6JDQWbGne
qJYJz43zLF1jHb11IvMMZeY1uxwsT/tuz2TEiGUQiBZ52fsbIol5s547Q6e9TAJf
7MF+Yamluu3LZE6yHSSJRuF1U5b8tdx02xgx2zTE188/fNFhqtBxwfD2NfVU75hC
KB1emWiC8cje7LGybsuMcGFCfrdj8rIzNdowXNx06mYbrRfcsFn58bzegT0tCxzK
YMIGNbbjVE88uNidrKVR8Jj3TvmHjaQ1lV83Pz3B1tZDgbikTJ9ZepZWYN16TAZR
cAwznaT20FHrixca/5daB6w11WyXjfqcioQ6bGT3DTUe4Iv353wXUWb/DQvzr+rV
WwhtdmfjN3OVDnBuc1zQ6npMAvkEQZNhaY2Obpc3doBEKgbM5cMC1qpfnAznM5+N
PkXosLDlkKORwDMp6a5//uzUY64ugMk4Ce7ljSYGY6UW57XKqMSLIvGZ23AEoCGB
tw7J9JcCgLiLHLa/T8arm0A1seL9eC5PZ4fsuLv3oPBdOl0tB5fgusraGa/yhwzC
XnDPEpWy/56awiDP/UQH7ZNc80UwIekbRTZQL4HXww9651vnMyBAKyxCEcz1CtfS
Lv7qdxMUXppQfekYwyczANGNEvI0FghFARiDCrWYYbarykRvsnqW1bpF5Uv4l6Qz
Rzbo01wWI9kFsVyXXQqIkn3yQx/VCEQ+sVajoPVMRlvlGr4emS+e2JgB9wCyGlDD
W1L1BtZFXfRfjocvIoOvAO3AVeY4eIZkJJ54gtXyLeMwULhsXfYJsHdxdI0N9ibF
SRfJqFq+Q6ZenV9UxZEf3ErzMhpMRxGR5WW+dEJw6G/2xNfxyl+DpMzQwGsv8QSP
QEQs+hhpu1tYOYq+arm09kck4LTABio2Yb/EgyUTixL5ehgkK7AAmaVoav2yeejO
/iR6zjFerHYRPYumERrVPNXJ0FZnceIR/Agfn0SrNQVFgDRwH3/PThNEmPRkUSaM
tC7i2Qy2k+AnFbiSXIJlfT3bf2k50ym39JZAZ+ro4RJV/875KAHGWbfHeJMLDtUG
Ijmry9SVBuJD3elmIoY8VFQaXDelDSCSxkVJNrcAb/bWRGPAcH1tiBFz9jZb2h0R
qp+gCW6tRcQsbu94GpcLuaIZgygedKSSmUA7pnWFJ6VNhkz4lrYbd+eiEKrDdnNV
3JuCaAcnYzKXH0LvdJnNhFu/y2oHnblJnMkOe997mgqDb/fpMfpS9yWldVlKQlpe
rXg24VYbsNrTl4VyZtRLMeokBiaSN49yZ/a+okKk+Zs1zdG7OqURjkRSem+waV6S
hSkX8Mw0jQsdsgSSyGRT7ulPlAehFFriOhExtHpi3dpGWme/ZtUvYEO0YPyohldG
TvfZ/61YkdvP4QpxK/bKg4PBBWWv7dGHyw2KTU85d+kDFJsmnel6fDRHCMVs4eT4
5pvFp+tRq/5XSR/1kcBqRSncCPmkBjjrUAcg3WyqRnwgEGidTpB4Gd8yo3X5ZRnG
jWPDqEKxzyDGhsQsU/rnMu48oDopMb4miB9RlalPCY19GnCbhNJgEk4wGKvT2gFZ
gwVMrsFDMUi/EqrzozOYw/tuWLGbkXiw5GIWzSSWx2/ontthy/OvtK8qZrOUGjTY
Q0KkRZ59OtFE4Q1K5MaGMgqlZxMRL9kLDUDLJ2U11T2A1SOrMMAXV/ZxTzCAFg/o
5NMqppdzcuulibqzWJ7JCxdJkfXHf2Kfpb0RqL1k/tUGVsB/6bq/ZEqF5zpPswqb
KqkEbj/e5hE2/T5Q5UQ7M0EfBWd9oz23bjawFpy2SyGkQELlKORSSg3TEiCtwXwZ
BOWDutUH8m4C9IgSI9DiJ6q1p4CNJsyk9sn/FEcAeY9P9LknB/dma0rEmgA0ApjF
AiQSY20iwHcH/9xb2L3yjGI+9d8llpW9hi8eM2ir78lULW/F4nyXZ10ypcibBlMu
bxzHlAghteNUF/HrmVW+j+gwOXj/PpzBnyzI2Zh2JfavNsg+/K0JjLaQQYaiSgXs
MdKYWvWS5y0LiaqKZnKvbOQqo5mrfJlRm+4ZbTFwFCySfAt/lO/iSd8O/XHoK9Vq
R3o87YZiJGs6bdk6bvF4vta0a72GBhOBx4wyIDLJN2yufwfBwUmEpi9DU3ZZchpA
8RtIUgOzqwxV3Q2C/QKNYMnBs+k0UxzQ/D8ilQ/8o05GRDrcFpPpcTTraRTBtABS
n4GnUgqPpUOghfx9jw+fh5Jw8rYazgorqWVdCS+9yvmRlPd6nTkkpV+Rpwc+DJsF
RvEG2fOMZB48B35dw2OjyYCxzdCt5hAKrXsiAYnFnXjQWR15slz6qYuGgrNxy1LY
CBplcy6E2M2UtOMQ3eQ46ude0cAJIVtycbXZa214kY5n4TACnWmSvPqP/tWAbpCf
i99XxeK7U0T83drMFS3gS0lwWRCDrj4UEGceUHJrhTFdqg7yIUiwcfuz4pc1Arsl
91/ED873TBOuSzfclQ2E9eQWeArXrdL6jdy3d33QnlH0BPOm7ovyWFA06bqioed4
XYbjw9gs4TFqU64zDqBnJoQpQGr9KA2xLtxJN54vbohx8JyswD/NbodjlPRI8TGO
2p5pYKTQDIEqXPkp2k+5om4I6HZOtDM7nxXtHoDLIQbN7CCIe/RHX+kYm9nJ7jAb
5zkrKRuUIZGUWqmMDJgu8yBcmIWQt+JKWeOoPtcKFQqYCAgCcTvk3X5TGU3cLnXN
PBEgrWvOQ3ZQPhZabQLOzkaixgsLkqy+SwjQImiraS17+8zTgEkvITfTNPB81ocJ
GIM+DMa747xQmF4z64vKi9FYQUvWhqwM+TS+nJYTwlPJUupuu7RIOEbfGGRRVxTO
N33WM32YKCs6Y3lusPag2VrSCbuHS+Nv8mKU3Pt2F8cfPd2jOL2KmEYFKZhMIKjW
Qv+J1BNAjVav68tQyFvyJcmCssBr5csOk8vGngPE49g3xbLra6A3kwfWamb+2xYp
7iT4Rnm6Ft1o/i6KSC0O6cyNwtycrSXYMZKDcXt2hL3jAkqMs291JmefhGV2/juN
RJewwqhULDOMQk1OVsm9tjwP42axBOHMkiKXg+xZjqlWJEJ+DQbpQJAYQb3T2FY2
+ztdrLwbcF/yVBu4c9jz3q7n9gOyTU/vM6xcdDYGO4PjUYp5yBTIIbWb7dV7mQGu
kyiy1wvhtmLrl64CxalwVrOE9GdYXdVY32o334JDBF6yjqJ79mE0ykVrjhTlagOK
oVlMHs5Q+BF6PMj92qYZbvSWZg0JXUpyy2Lxbx11prVLzzjhVSt3B6fmNu5sralh
B5amYgN2/E6Cfq14QkwFQQ98aQxpKg573HN6Gj38dPXP8psn1EKYm0JhdwtlNOql
tJiG5Nkk64Pfp3lWm9NgAQC83BG5bfLKoLIpVnWhCp34tCG2ljX0G0GUUA6VmqXa
LNWwd+OfJAWwUKUTaOuQxm9ITCXX7iiqC/lX1rs+IDNpzNoYMHL9udkJZ8lfQees
GrRH26c6JGP4cLv1P6q8e4IPIa3VpPbUzi2D13osBMpRy2WqLFSVdclDUYAs9IrY
MgyQ4RP8IaU92l9mofw2r+z07+wBz/ZqBN0qQgmnGCodRrTibrVEL5CXAOG+4xEL
UilZ4oPPnFiU6IM68TEGMeGZdGpOQp6sAWBnnds43z2tY6NWclPsZ6TQyGiAy2Q7
c7PwGvaoKtlbYDRB3fQNw9enHZYHGG1ALNBVD4PCdJsvvJZET5ptgOq3xnAzSpNU
sy7sMiXdeqIoH6pM9HKmwNi5QcasUbF0WiFdRjJcxLKv4YfbNr0IS7gBfmJdBXP2
Gt7hRLHyL88920656kEqu5J17B7Dh5Nr6i1VwZ5nbjxlhDXZuxtOjV1GGFFSYkyd
/2CF5zVd1y8aP03qSQLPHFJQ5bi4W90iuQf/62MLLhmBo3YO3bLrzzPgTpg0tuRi
UXBW7JYiAIzuSSTsVVuv9/XTUvFvdXQwzGQjyZZcvnXPWQ+x1SoE2p4MNP6L/xHs
i1uHWvCrDpAC/5CYZ5bXDopHZJ6jSQHF7gmRSpVBFAMHFFnvg8CiKRcYKLvNN5UL
Vtu16IiWCd4oWzxHWbSbfJ1TakWctXJS3xeYMaMIgIMOAAHsAqmUpiYNS2MTnxpM
l/pPH2sRDjB7tlDZm2+/MMCeDmf8kqmlKfzgiJ1AyPz4dIvoTC9WVLu6+7bHdHtH
kLKJql1IxDFPZZnde0XCTazoosYGR4Ww6HH88W8ek6KgFIN+r5TRxIcY3QKkJG8V
X+GbOImG157dtk74D7h/XaRwMn6gxugFB+8HeuTUGlPlens5GIXYD2wdhVOd/IKZ
8cHfiuDYv6UnT4UoYWlaA2DqQ28aJrXBE0zsZexMwXkOtvO0GM2fKkNNkx3svanL
uLDPX7SCHnETN85A0hSu0dLz8rTzDBelnQuBLUalP6yaBARIpFH72VtMsxDBQEyt
LyoAozfHA3mv3az+mTHMXnwe/6+ysgimdgkv4P/Xan+YB7kvE5hhvpTG88C2uQfE
RuyZIiXk/oBpLLRals/MD7FMuSUNXm8S1oP8nc8K2GQBhg8Bb/2x21LJkvoiox11
owRaP22PD3+f6MF51KowhcEBO6yfIKQqgaaTVXWWbhT25aamAyAYxZ7c0s38dDAI
0OMz2ZbmYnaITJeoIjPgLPBgOh67HBIs2NEx81FzLMRFSCbV4/wgRwGgUfGzu7j5
jVKf4GW9txtyHPqWDMq7mYPLxyuFM8Kg2vBfDh59HDTnWNnhz/cNkIpHccV/VhuZ
9drBvzOF1sMup5DZluyUBZeqdo+9Hl5v4gWL6JswQShcGuH5qO4DT/sj1WddgZha
8XZ9jGG8fYvcmzpRjlYQjcHsroewANPo3n8JWCM0bWjKpYw/IvfSFpJqmwtR0PZ5
vg8eqJ8b8I+xDhxrSmo9nCiItZWibQWp2hR6hZf4kQTCt+cPGC05gmMB6kp7i2ei
SwnVcVfTFxK63jzT0GTJJhg5k819jFVewgGQhgZaAacZiSW+/eBW9cH4a6djcqZH
lXdhk5pNnZPte5Wak2Fd6us6kbZpvD18YHfmvE+miuvQUdR67wxtO4T+xT2i3REm
BJ61riyuAJnvSenNSU3Rnq7racafjco18TPOSx7T3rAYhQTvKGx2+Lww83t7w+Ie
TLYY7B4xrS3uaHvvGaV2iOBeGWSEz17A5CEzO09b/GlUKU9lrnYxN1l81GmLDMNF
HEZkaZ0aK49PCw1fB8K+DHBCDXDYUNAlmyis2mzWko/dApJ/3nTi26hEd2e4eMbE
4nQfJTbxNzAiorLmW20U8Cmmc7GwvhTtstSLT60UjDi4zarqo98mw10w5ctRyES5
L0RrLms3J/3fr3scEoNP5LVTAls/fbd7HMDA/N0nf51jCNUTIKXNo3B67YoVHDfw
rliPz9Fb9zrpRhq4XrIs4LnYkF7FhVGJq7FgragOPs1KY0ehE/I9Yp0XzDn1P3BQ
+QSWpI81CjZ7EMfVTev4CGy/zwpbkT2IQCzi2PrMM+Cg6Y0Mr8FhOx0FGMxNFj/V
PWgDYmCncFlTlVLHxRQ3mDWkD5EnpUCWSHkHkO1Z2oDgzxlSxiqpQVAAjREAFTCs
51X6qI16JoCyHLgVfAjKa5DAzxsTQb/Ha2+nxNyoKQysu8AWgISNkB0CL6hXthOk
JRv7t1mUdnBAobGx9dN5eKlQWlbasOjPCXlm59gNA2MfmN+dueKqnoZWLQOymo/R
FPY+fAn8OSothWGV1Iz8mFnqk0m7SZrxjRERVTUHQlQ1afCdP/wbIZPSwT9x21F3
x9L7OZD9iwHjWQhtgc+hCh5EGEHpM3f1Rtz5CQHrYrJMejmphu9n8JkqFPV3o/gM
WckLxS6Q5Jd4IEaUfq8VXYZ+rCaRrByTIASF4T1QLwUsuIUll+IEkqCMLwEAZy1I
M763MU35pk4pPUc3MOOEoH5UAsvptKfGAKetEW8CmIOTt06LhlH9i9R+Gnu9Xgjq
H5ecSr0+Yo3uQF7rxzqx4y+9bg47SikiK0Z6eINW32dWmMP5wQrZIlSnCTvySMVi
89cxKS4Eru6dIqRNLDx2FY3MBV/SnSMwX/XnbWOjkXftTm7Zn6XoaPc/uSy1ER1Q
tHGsoK5shfaU2qgb2uxmARXXVug0xX4lt5s5gfMaZX7SAx+l8Hmx5aSlKPNdQv1A
b3VNOUc/4uUn/emlIY8bppc7L2f29cs4L6w+Qzn4tjA6vp3t6CscWGkGMEZnMEpZ
ox6kbDRibw9EjE8WP/QCgeLKQd7pbhFYSQQ87qA5XfRmqq2vvIGuB9vzmG7pgv+k
zh1x/2fQHRipwh/sar0xcTwqyFLBTkTe79LMU3uKShtnQiWm9mdmGX/V3uElcSd7
xzGZXp0ISVaoIhiQA50qp/AYcfproOJFRlCZEHkvOJvm3ICSiAg/loVBgPNzgRmz
Xnhx2Qwc2PBYz3cPBRe0I05pTey6SFqr/6YDUWx694D88kQdsflYhOVPgY1EZ9ZT
YhMwWSZLniWxy/NmQwyLEH3E4Y8OArmcUmiSqvCBHes6ZLczsF6z5WJInmUgmAZG
yDgbersBwh92l/PsFV4HQc/Thm20GDVPGIfnOwElRQ9Rl768Wk4Fmixx9ox9CIqF
db644fyl4w2TyTw7q/yBgwF4GiXAgYoohW1O4SRzLAjBHrzCq++FdnApVOphP8D/
8U/J69m1jcNv3dA9XmgiZrkFuTqK+iAb4zs0OjMCziHIg5I8H9LcoGfROTM5zL50
yeUBwJsTrhJqcBQKl+p03XdhsHRh2BiNnyjX7gpT0Nv+qL1KidNnPBIlhRVflimA
anAIQhYiCd8aaWnygdrOY87MTlnGDFUjBHlXwwtQqazspbnXzoOX2yRz58iQUdOg
wgjXk1JulHr6nbiQ2RFaBP1f+Wnnl8T9ihr/KrwB4XhsR3p5CtN82dg5zk5KikgF
D/qmI8J5Sgv7TnQX+UzUd4Slp4N3e1Z9JbGTz5tel4kCP3Fw9PNk7711TVYxR23t
p4yeDl6WOZ33LkDl6y10/eJP5B7mvM8VXA/ckH4CqQfTANLH6yIwCIMjaQYdd6Jm
F2EihKcCuRkgb2a7q3udhjC/rYIugRjDJ9A/E5O1JDRsPJPKIr7nxFsjwHN/IgQ2
2NGFKo/Px+/sXegZjD9wK2+a389p/yXqDg6iuTm6izTzXuUZ9AYLSPiO9X2fi2UQ
DCtSZFqkzWO6AKgkeF1amrQMHVjIANtxvtrHQMetel6UsSBcYAEc7zR4mGUD2flC
Hs1uXBd4LG6ObJ+pGhJjcxrRmBZTbsyOYFcfuD0+rXgBPoh6wf06RCFz5qpPBHdM
WG9nhRXS5deQrxn8eYNpvLh+RLp/hsQVFB5tWinethvnVik+gvRaGt8Gdvahq+6R
3GYsoh6fL8F+YRE/r+sxiFa7GIockYAdQPeVNYBbQJ56VNs75nNdEjhk6eBvu0U5
RROGRseQ6HZRnq68SuQXucrAf9oVdkXY5nYyNr3QTK4NvKtQi2SSzU5P9ybsCoST
YAo/GbunqrfO4RAvE8SE+OqNhxVXO7+i6jo9Ao8fjUEkPqFLagNxAf4mKS/ejfu1
mt2FI1L10sMh0vJSPyVU/L+Tyat//cDWVqTD76c8YAoECpXCCKJg+VkwNBwzk6Qp
GO/u8R1bYTNlu3BYU/RVghEu03/vPhYBXyGhE58lI1ZdM+V43zdGRGlanph6t4q7
LKYpuKi5qRymmfl3pzxpsDBz0BgZ9Tf38/TzNv0OobMdwFWhcG7ERTYCtflb4z7W
9sszfNzL0tGNEotpQLphqV7PygB5n2TpoLBByLBTLN2dW7KZzMrJ8KPcTXSMBXai
H8VZY0uAHprn1uDr+PB1NVmRopH1WH7mdlAWnwbcq/HuFW+/sX2ZfM/Hy1cqvxQ3
ydvKLmfe6F578hhrG2HyhO4/ycUmmt52r34vwXgybagveNHVwc8Efsa6zbp5OKrA
lVEnamDdOnHz1JsrDOy49OiEX42AwzuMr0xSLERX8gXBqhEZipmcfrxwiR0CzWbV
mAszDSdSxsGWB+KMq+70C9gyFid30cNJXX8F8+hWDAi4aQ8ojPDD5eCMHWqA6is+
LDfy5cIpmkcmaPp/mVZZ7SHoxpY95NNyFxfNel4lWqeiFU66lPb7ddS0EAGyLWYv
Ik00qNl+u0v5pLOU6+UnqCa9OVdMT6n/w6PwzKGH/zY4mztlfE7cDdjz8gq26ZS0
QXy/QZ614igFvlDjup4rKcwmX6jkaxVucNKM5jSCYquBd3pF2zmoemLwWHbdvHMh
NzZxp+0CuN7SGZhjMZ+uWAeCHkuXb2D44Ggiw2vDad1FfIIrQRGC8iYsn8ugCyMN
8c+igtuN3hNns59Fzfy2rZ0mtY5viUKyCemOoZGZCCVxErrbVuoplfzjKIa6v7Wm
K2AGbRLRToN35PqbqdrD6bvWJ6/L3hK8QzDjeEcvYgTFaPn1MVxvugzoF3ekzW6F
gY7sZS8urz3QGCozLuZ1q9x6BR1lrn6JmLXaL2+R6Lcif+xVXpuq4czJHTnbKKJL
en1ScECxnpnQGKYx+DyMPuacFcpatLtPE59rakb+Kv120jTlyPeqKo5Jgfb7NEzQ
Cr3MygQ1OxYmMyjnGOEC8lAmZC1pZw2c49odzvSh9LmPUGejVHSkHp51rJvqbFUU
2aG+HJqfPN6i4b4MwA3EeByIw555fXeJ5tYXuVdTtaZqrRVubf+JdcNljAWI91+6
ct7WbmqaYQyBuJrissfeHimSiqsa/BMUzriHqoEs4Xbt8HHi4x8qt3jDMcl7DBHw
/1gplrpTW6J3iy87hkZBjmTCNo+PRh/s5tfhuIp31rBAoIydn+0sYBjIpRoOSyvH
1yXXUZx98eyPPA6t3ItSACqoA7nEQ47lydsg01Z1tbuF+5yo4jzFF8q5U2tJSIa6
YvI0mLmP7GfLz/ii//s5USN7a7oG0vXuVxgg/t/ZEyRveABir+nKuA+4Pw3vlUx8
mwbDz8fLCA9zuxBtNP9cSZ/T6oI/SuZRQAyncod3hRYUouClNNyCsOHgA2GB+j7e
ChhGW5lHYq6jMZNrIQWD07T50nSyis7IT1fdzWCzHhwUFv8NjuLpv8S/3/fUcuSi
vyVGJDr2b3G8e/pt21EULeI1iivIhy4e3jBDZf4N6T4vBHtjZA0vVmOAPtXDdGch
t0xuh+xbD6PkfapRucAx/1ngy03QnnbbVnp86/S2G+LMVhJLFw7MLskv6r/Roh/J
2sbkRoYNIlcVp1rYeLGFvIaxpuzApJvtnJQ69mbHEUwJjyTdQJUJwuMS0El1rF1g
p9ukBEbk8V7BaCo3dBQCgkIe8HMQWZ6XF6IZjc4PvU6qdTyTs0yPI1/bHKXtkoRD
57BcqHAH/0xMueugmKNoSjBAZ015nHMVcDLY0N3J0YP+cIcK3SIHlmEj9TMMdzOe
wi1Qphm+x6xVMmizXdp8PNkfxok2xFaH9pQuCII27O4/aFS0nkDx4vAA4H8Kdw5Z
WRwYv3FC/CPgiBGsuukEWyA0KUZZB7P/HyD9U55kEtf2MpW33taACp/5Yj8k0tRE
SDTGSX4Ei4MpBAXBobUKkTEd3qKZq8YMj0eQeiokzNU1CgXv6uWIrnbAijUJa9tk
5mNKvkPef1ZwiQCZV40wn7RS6HPWA4BgkK67WLTtdvSeYUJCnhTqZer2/E+IL1Tk
SddzjJEO+F3eM2F7o+lUjlh1v6gyofMWH0Ynxi6osqksJsaRo4P59z0tfJwhiR94
EDrs4aQYml/7Sca/X7wSsPA8ENRPdY5bT2Txlmmb44kDrDH9ZbqSmQ/I/YaxC0lx
S7+vOx3US17nnsjMyYa6IJ3Wa2E/bO492ijGr3a5ePg+NoapeMMyMFe5rFZp59ru
zpyz94S5y+d5xap1bwGF0QAt7APeJLIRe09ZWu2ueIkwjcEmrjRc9XSjvwp39ff1
srZA3Hqm6mO0NVPlBmU+NM75lzMOXVWmBmaYjEkIeIsuPagNmtUiw+Rl2ZpT1lVm
eD7N/OUOMOQGVCA5PK6v07OznCAsQbNqIUqlRaG0ydm9VM3DzR9ffSfWE4VWYdpz
nB7PX9AhoAwNXXbZmibZsgkWnE2OALijeBR4m7++46swQFCpc3OmkvOgPGwo1JT6
10pMZjKLVOIXxcMApQ69mRt03lCh2MP1WiWIEfaOiXoUL6nF/s7gduc9/TMH/D/6
nfPVHj/mWPvgzCyGh8untogxXb1hwD58Nrr6suYjuDTseoYb+aKGsGea/4MtpFWc
xYqqAiyZdPmBpL/P4OM7vKMtY2OXtr7QZoGzUasKJ4LQGFyesuoUFeKLgLDFEJdp
W7o0qN9s+NCRmWxGbVvC+RhmNcK/htxCAVYE70Zmz/bZ+hr46/Og/RdJ06GyU1R8
lObKPJaXK8flYRIO8Pishw6hQU7hNNAbj6Lko6IzLYemmOt4L2fwqTwktYjKXAsW
ILS/b8NIAxLiJ0KFN/ncyOXVgmI6/c95ReRRM5Cn7fLjffq4oW1YgTR+ynNootXA
purp1mUjpKQnyriQUHA0B302ktHdBDnzg8k/DebCX/E/MdQeo8rw1WIUDpgA0ZVZ
nTv69+5sSwPCu0FPPQyM6WGQPuoufeM82+EdAkFpUMa56eQ4sSOndeZU0wK55NGO
GXFvoiY74l8D5hBz3nf69Mw+P6hPN24vtj3tRRPysBvnLHArWIwAmZq58fFmxGw8
MGLHgSjlzw85Z70QytxaD+V4vuVBbPadLX9w3S//C7qQRff0TE131cuZRCtvvhpB
18RawZgkWAz0S1C9lbd6FbIZHmS1zXyG/ZfHyxEvjPbErqVRxHuMMBbFTo5QmM+L
/2joS0Hk46jcOZqux+tbkwMwoSMfZTyu/W4T8QqlMoAz5EP6lfqJY8KJh4gLxKXf
udOKjRiYqe6YvVTV4FgUW8rP6MAOvtx/yz4g2fVgtTKaaUgu69hGYQslALIqMqEW
gRkJ7a6EKXoHN0v12u6H34K2aRYJ4VKMf1g7uEJUjCpXQPvAeA/zj94qGfG7AL8O
t6VdSyPbtCi1gZv79pIFIooVLj8ecBkw9Iv4PB5d5quOaabyw3y/JFFvGjPR+xZW
fdmufBOGg/XtDKIJc+zz7/ITfJmo4Vv5f9huI27JBnIq0HVzkHzeJvOeCMF8YBzN
Iyi+vhSU3teShdCKukx+o/eWovcSgiNaIJjn2eAUH9bUnceHtibS9BQesWH/1Z52
4ymEjYNdm3PJi1ZM+vRi+lSPDXaRmVRCPVX9yd5784p6W/h2JurJMcZJ+R6PMuJM
pWViCDt1Kl6CbED24xBl9NMI6MChUUTMl9uUwCSCpyoaJytiDifbdZ8RFOYFHZ0R
D0FDggu1ZJq0Xpw40Zdcw2rNYiwGaTEEySWK2ryUT8ICrF3JqmSgo9fbRAT+U6aO
F2pFTSDZ6VP+cJbhgoeM5H0nJe3D3WVN0pYwpKDg0SmLvUpXNwMklrOfXQq7ertW
RRTdCXZUNuzAe8h50Rz+FcLvTiNjm3RImlXQ29+dq+eAY6TNbuMAwLtENdU6Yirv
znxHG/m/14CyqoM1NGSHZiQvPNcOXewZMwikbWJFUxcmZtOPwrzYEXYZhSGMpvQW
XtCeM8OD3qUzlTDHjmXrHSUDD3XKiFZdCM3eGishbVWm4RTGTcBGi1Rpj9oTEUM0
6IDJSbw1nF4Gb6mMjx/542lPdEOxDdvWjuVSJr7PIXbo1cwlMfHtWUGB7MT5TkdC
sENrQykwdEvjxfC+8Xkf8E/Mlz97jizxQwGNTyTz2Y5ThGC2k9y1ldkYOcLXvoV7
Un2BpQUwz0+d8YuFYJRa4HTcIQzCSCyQCUipyleHWEtfNdSablb+xSKdCvDIWL45
cCBGhjuewGiK0tPAWSjJcdqwiTwKUKCMQVRv/FadSM6SUve08ox4L2U8jvnR8wS0
F1AELp1Y2yPW0EY3TGEUz/4gTgpYr+b5l/XW/m8RdtbmrdKr8lO5O28srJZFL91M
2YNAxMGGCGuZrJjJo3wk6/I1WhUTu3LDT8Y86oyYyZZerzVW69c17qYhKX7QqZUD
EOwkKuTWCwmF578qiQctq9yql2HcpLmho4UOxWOA/f2V8QPW6QX1N3+56H2b/mCe
VeOkdA0So4MsETDZaYgPnxaFsyZyHZ5WlPXwIqPS9PbibX40+AuJfUIgqKgB4Mwe
h31E2JcXnFTHKJNm+86VW7lvVdlFFDKKDsutWuUXwE3eDhoz428iNR5ALjoYuM/O
TKiVxppsqiOv2BloddYMwdYIg7KgYvbTCTA8v6e5x4umKwdNHyexHQKBLixMYkPS
gVinEyVPTXNlO4Brey6IWkm5T7Z279v1+KROOdDwX5wB7lzem3ueV8Gg2r8XKbHf
QtQHCV0L0LEZa4fziRE8/wdd2siwtInr9/g0gPHDRJubW+UGEUTKr9BOMQivHnVq
Z9cTggUrzeLaOdeqSZcNaZxtciDbbS5+ZqzNH+L10XWcl1G7Gs7Ik045OhPWwQht
SW6YEJwbGH3j+WAi56LpX2aGioBjax2slI7v/tzgi91tXIorLiIHdWxJ/smAWXct
F6qEq60//RNx/80UMcxPDJbgIxHaRlbL4oREr9ALnxvUR8RNzEZg3DNKbKKMj38T
mMHYWZ9+5zD5sntdYm9T19rUpPnJxDWUXX89arYGGZWuuYXhILrHKLsd+Q84oGKX
16p9ZtzELj13RuBgP1MYfeqpCfwT1xJA390VoCSQyWHTZJePJ+XIg4PxEJmnm20h
JiDh5a8z9YUU+VbchF/jbzAgw5XMN5HmdRLrrRMlgCG/iWeM/F3QVqPNkOeVb3IF
XQyqvL3G1VrDvdQnwxWpc4If9Gn2xMpgphGNS58eoamQWPJ5pbo6Q564GXg6df9v
P+0dg02Vy4A9f+fCjQQ7sFB4oLso/9W8ADKg50xkngnB2HVefEye3QRq5IFJTk1N
AnqljD4MJ3N/bzWaSgL/9nz7xrA2NHlSbCWI7cXIuwGZmYFmGfWE7e5G7vpCcl2h
TZEdyLDIfv38GeZ176qUOJ55YbzD+ISUvRvD3RXlAcciuaeNCYCQ237YURgtqgPi
R+QaK2VUEDRjIqbFo9Wr9S4zSlW7vLW8zH1OGCe8XDFbWvN3sFdIOZjBc2qxJ47f
xST7p8oAwLurqx0fz+3FmHcUZikkiSIiq1ACYcb5v+8LmuMhzYK1n+EaPk7emssd
bjd1PBHeuiUI0x2geNut85ENyOO3SawBDcwBqCnT8Fll8JKqSK8nBqGuq/k2PFeQ
Oxwka4ixbcDBE74rjAkSN0CSs6yfdtbwPu06AlhR94R54u4GPT9G5LaZ79YMTP1l
pgTzeDcuKUFSRpLDOha8HXzS6J6mW3ihdVugM8uAIE9M2YncqFxyfbBzN7dJewGJ
7zL3zqchrofDo3Dvx2aM5cNL+V1AbJuACjg6uYhTAPZKOu3SyJ6+ioWYhkF1QJRX
M2LB5e1jn/Z73qYsLiUoQWOI5XDPX9LoREIZPh77CcroK1uy+WBhblz1e0vkf5lt
SOBi7d/12jpBjOqKGWYcYfChMw+vTftimoSjsTf6wa6vVAjXbdE78BySZxBBtaap
had0F+F2EW6YlLdZC2nnogh3uTe9v+sHhhMepe0rtQIlFHlMwubMqrfZBDNEAudX
pjAL6F2dVjGhImG8cpPZ8nzFK03ahV1+MpQyXzUf2180XMb50whcTtifwqV9bLrI
cPiXF9DlKNjQGFmER2He6G54sOt9lPhv7Nhv7S6bkHABJ8macMXZPc/EUC/83BFT
/LNziImgAf4HwFM3VwIZDL9qL8oR1zhjFcHc+VuwSCYGYtb1Mhlf7mGopCUVUOeE
Aqb8QRYoY7lPx7FHiBhPqX2AFpZElnZ2804/hvZy9Jfy9uDwJIMz22VxWOrpx+xB
9OVliraGA+sAC4X57quPMUdBiELGz4uU7QeW6cZzckWzPP38z0zPZU6K1hU6PUQt
JQAClfXf0rrUEkrizZ8RXAdhxK5dLunlppoH1klZa2MLqJQBiIWesM99db59D8CX
cnl+/LLdyOPzy52mzGCGOgcY87ZyRkmIGGUB/UtGQ5votduaQCDxeTxvuT3MXzJ0
MK+Z6fe8nwNFmJ0WaRJq9fxA6tbLwi3JUNOGqgD0boaqLF1RjS3quENk6xCFOvcT
UdSCVkGvt0f8pFWZrgh7W2Fvix6U0D9zjvzV66V4wXKk2Ep91fpQI5poIgpMMNlW
hzbfY2Zv74GGcK8o5einMTE/ahuVseEsPgnFqZz18vu5ZMj9wjUZQjg8uRenu8Vl
Lo8PmVgRGbfWZYOtvBIyFHOC11EmsqXFI/AVk0rhppmN2SEVLPswjyLWb/VJaPf5
e3hJT82ToXZgjh0Gh6YtBnLFhQIU4ma0QDh0ZPUJBvLLg4OzLPwGEuiLymnSFUJk
OfQ5w4EsRwH5OJJzm0ALcm2get2JaLC1cT20UGSL8EGANHw5EmKfP9VF4ZvMtg1K
uc14oN4HjTK7bnz+OhI5Ma0Hh70/9tNWjJvqu8vDCcZ3uYzxFLcYZfP2mFXjyaPO
PRLeHxUKApJf5ujk0Efa65MGpY1cAwKNSYdtCTFaHSYOR1qeHQZDxiUOOjhkJ8hV
Gmo+uL0jVMBS5EjetFk5J/ZwlVTBg0Y9mynvaucgNVRUz/Xj89i5spJJj6Gt7a6g
SKfHt3XdBtKZ5CnHNj87FHYPTTTXlH9IdV/21hetrYvHljUOEiaTG0DLnNeJjWBe
Xl43r/V+wRLx5lA8h8YvH8aB/05D761F6vUF+LokdLqGJFCodSTj53Lv70AuQXHl
FY7L0ur+zDpqCck+Y6SgupAOxy+kO10tlEqR5ehy2CvDo3M91eGSOOMNDGjQsa/R
nu4vBDV7uR0b3ceB1cp2oyEJ7TITTe+g/7nx6oxOdromVGtZSyZU7oNtQNiFTkHp
hpWqpiupzsQIEdQ8xhwF4vqShq34a9VGNw7fS8LGKKjSqPBr6zANCfACb5SDF/9D
Bj1P7VwlhFxULLXMB3Y8BzkxrtrJS2oCy2ILxd5RP/nxDZQ25YqWDiaAlcu/aqvw
ya+LkZH/sB97ftUpvd5avBCGLM7CCwcMfHtY+JFFWsu9EOzc4r0/JEU9QziJm4ds
thfQ7ta9EePv6SXAdGl3IFmRKycRn67EwuAyDEZah1OHKL0VXGbaaoldcDzUNB90
Q4uylg1ipDp2x0Rvx/HEmv2Hfbey0ctvIaBV33t3H8wt79eMp7DsegNvNqEzVw09
k9d+gPSLUCrrGm9wdUYButPKcnmSIwOgRVVhaxZjnXTPza+gQsRtfpAMJWrzxTsC
qv0LYhec0NW+w/mfAxVubdTq48RRb3V+LWHB83zOJFJfIPPwx1YDH5o7L3+bpYM8
kt7h/zwop/rmtrYKgPP7/tUafhaeTOvKncwYHAmCu0CZqIEA36qDF7eV/S3RM/x5
LRkBRmpVHzrvI3dSxq6b5lKhxzpIc0SpEcvs8j2jrAMIqy0bI3nndjJEA+nQwsq7
g6tpfe91NmIxbeJm001Uu7rQepSudaoTePt5tgbcAuklTDQQSCHBrF+VupvPaPyk
NVYFuA5vmozlhkmChQiB9ZuLzHHf8lxXQabvBaMpUcmfrVz5oECaYlx3Fm6XJ0tn
rNKNbUbYijGN8qfU13XxQwXN6mXPqPvINrDEtnIsk+sKWU6guIda8P1nV2137MJM
YYeizUz5XpPAy8oz27UVufZZcilSgyNglnS9PcQMr0XenZLt5P6OY2WB3w9b0aQP
w4cshaGNfccy/CM9zyelhOFMa/heqI8cLmEPf1ABDLITIHdUC2v9L6o9hsUX0piy
LLdzab2L4+LkUaf4iyMzNdPvz2GAPOIa/xtofjZlvbqcGbLbXZtjKwP7Xis0pVjX
ad+LZ+ow7Ma1XjWJclmrgtB1EaMhOXgvf4tZyAJocJd3jB1OE0lgIwINNjiJPoxa
p5HPRdVHhdRhD0kd6KhfLtOgpBu4zJ7m99wEvc7Of15LaeGd3ZJk+taY08AnEAhn
Ccmxu3dDE0eKQcf1ZkZwjPi5FQZffSkP0w72f3sRqd28AbNsJyPSp4AMa7J7XFYt
q2jeTt+n71Jzn0MBCi7ig1xcpnhKAOjC57M7wuvNI4qC/hoOEU6XpBiTkYuSnFpY
4FpqL5eUXzRY+6jpAFBAnCd33REvJnEG2E32fI/NW7qfflSMMZajeTCzTgWjkH1F
zaZMjCHDAeopbShb8mAYY8I/DSFuRDoQ5naAi4/6TvKx27Ii01jqxzruyo0OZhYo
QLlLV2hkXfPiPHu4KEvtA4Em3ZfPxsK77qHcvISZ6XZRsvMVAPMJZMiKMcpqL98H
I982X04rP5F3ujr13/JCexes2UfrKoRLy5cOO3w6kJZNVAiaaWvR34sCrtS71Io2
SlMq3Rv5Bjd1t1uH9D7yyRn1wlcGzACLh/hzXh//zIG6jSi7A/jm51y/nLWForyO
/nMiAPTDWuDrnXaNtgaY3hugTonLddVxYYS6M7T6ej+ym8NFsSUPoKiMemgfzwHy
ujtXB0G5KhFfcvxd+q64/gYtIf3JyP/p2PYZ55BRwLLhscjb3LeNDEy4JeSV8iwD
8XW7mfWUtNObJu/8XhMbAftI/3llBrUTI7C0+GZYSJKyvwuMiuH1KsgrbFbkspfr
UJMThhErG6X4ubkiRJqnhtgHmXn/WLcJToYvUqcrbyVuXbd7Xxjbe5S6ZtmNYu2r
2vTvYptN9xJmclGr0zTcKah5u6QyWckb5bDDOKRVOXMu5KcnyXEbLhKLRBvGY6+N
kKoia1IlbnPnBPgBCofZUXVetVtH8OPHOn9qXlU7fzHhBJjyr6R83Oq/QBm60mEp
ls58hdLqMM7EVzmDU86EUFqthENLM3qKL4WJhNLYuG61/LgJHEQdJbx33N7LfyB6
0yIePzxP/tVzhZYmlAZLoC5Z4ow/XdXQ4PFh4NQVSNtOwnYupR7qlAursf2Z2kdq
x7VzOX8xfaHMf+G7rbk4I5Be8ydzJEkxBaPqR7vst9hmj2CBGBUVjQUHveVuD1Cj
5ZwRmM4Mlo/PEnKP/qFvZzA02zjWQQgzDrUV9nBb05T3GAMc3tqIH7ycqTsXZDDI
cg7Sovk4vdIbmyCqWKXCtJ+NoT3QgNSM52SpFllzeB1mkcqpnaviLB1mrq6ATaUc
cCLyUDf3sUNdj5jAuTQyEZBvJc33xhZgMxIRkGLpycKracjDHfYm8tt6HYplc8sA
44tvtHJrjuytodubKbf5ECq6WRElJz4nTGwtMO511wbXX6Kgs7JV2Yp5I8yy+Oe7
/D4uLV8f6N8As4m9XGDRhCIpgUPl7Qr7lVkBYp/y5e4CvDWU4yVwLkQZ/eK+GxCq
zNuduCZ3qMy2EYwUi9SEt029QzWjH6AiIu2NRTFuwObK+Zmj7X7hdiWFNSj49mgX
uBRiLo3tH9cL+Klr7rcYUIkdi8s8OSAUyUuh430eNEcT+VIZVN4mreyHxbqskdq+
IyFBm8fFy8x3UEunD/ZuPPeoh6z496EN83mIAgWxednQ2a13ysygkFAlqhK4oJTe
NIE4wH0rgnNW8vsXxEZAPMBQuyAgT2yPtJgZmCrGb6C3cEQBHVXwm8F1EbFSHSY4
t/7Rjvx9uAVn//RU9ufNSJqVDz/oyVH6JPIL0ZDSRlMq35B2qahh+2SuFKDReHhC
czO1fbC0zVPxAKp0awMrkyLMJtdfsWR6x+gw+W067YORZ7k5kD/jk5LIUDw1Vmrm
oQa6Mcmx4Yd4sVyl1oKQYhXb9jzDPEa+1u2WbUJajFZqPxAHp+/VcO0/67tmgaNz
/zNrbPHSEwmHxyz4Ugn3G8ERKF6OqNNcB3VjUWbBVaiIuTBt/lJ0/nuIC8U04ENt
XXXqa2bIoRWOOYaRE6A6Bhd7mKkQnmCY94z+PJoTIcnfrMyz1eIy01PV6a8LZOHz
12fVBr0cIorjjz+NWUF0M9+wcgBvTuOyfsAfN8JJO1dkqKQ2pV8rjyccMz74f5lh
wCMYBM5CaL8Gg1mjdzgs12dX5nJcW5qs8ulM3fuDTaLeJy4+wR/pEJ6G1hkIuZEf
GJIiyhcrpTXEvnnr5I5+adMYpxt2oBcgStm4vH7hI8q4z62Vs6Luazb44gSJ/D1I
3cUFUYf+Gr3Nf/MaWXtanbEVH6A/MgXHHhRY+4rs5pYMyC1OT1i2zBuRmts8oRQM
Aa8ke0gKeT1c+Vpfv2+Eq1A/KhM3NbwcoOgCnIFMf5AMjbkXAYtPLwBNfy31ypSD
VHHs4y9yELOwynu1rdRejgSeKFMgG9CW3Gyk3TZ1TBx4u9yEFIWvgMz3lNox73dm
L2bHJcy7Dm/EjxiGgeln944IPmFdo0aKrcnphOV+yxS8TmOndnZCcdO+D4E4KxPx
uCdjaHZd7lw4V/yllDm84HmwY/vjWo+cuhyd//0IzRJB3G9BE7Eka4O5t4UZgwvc
+3TIKNAvSv/f/lQTDK4nCEyUAaZM77wCVHyJs20ODN0F+I8rbdJFPPf8b2zsQ6KZ
5uEh/A5uVk0KvcO4hDqbPDREVzqSYtCQF8XPU/+nGZUJRv6AzNskedGR7NQepGQy
ib4eLRMy1SqkAEVkbLZtRJKNTSpYrfvF7F9l5BmE4z0l6PCsct8O4G/Glo8or03G
eOQk8Qya4F4Ztcc+XC6mZeoT5IcSxXjNXQ5TyjK5DoaSAsJDbcw+7f6PVB3f8brg
PUzB7TjdhDCpI1je2dEdXJqc8t5dRPRytA5Zm679hHHAaYUMif4mpeQ/hVUYdHjL
bj8fdDor1cnXGcg/wWQljNKfRnjc+zjNavIZAkjbOPh06wW02e1yXJfeXaSY3udr
i1K7FIW3mELRJ7NKp7n+F0tz4xHUPu3pGUAiiy1ygNs70ZEY80clPHGFpuAluiti
WZibDY6s1ZFY5mCMjeotS/OyeHc5zjGWCLdU5k5ZBv3xGC74Kc0UHM3ejDl6dYGi
p0W5u54TSO6VdAzfgCMs8wlPaOstFw4mcrBlxaDYfhj36CBeFJfryK+Z34+lrhjZ
LihFOMYnoqwL2BeMNeyYMERoAKECDRuo8swBLbQV+6ScKR6UcfagAPiiNLoHpdO4
aHl6ciP+FfrhlUxQDm97cGnNqab6HjPsxqcx8Hsx/rcfJAEjY1fQCVW2pW7B0DXN
tEE9ewyCYZ7NUryGpl4hKbQ9GiPcqSwfejmk0ZcsyvVBP+sJNhCxunnbPMCC14Ah
2pDfwT6As7kfsSYHkW6bSEpHo93W0kuqzaEPoQKrvZjj5OLbnLRCWKMgbqsl7Chy
Pylq7dX/hy8KbttWqPeVEx5qq+PuDs6Dl6hy+ffbiIxN/tpozH2FRpWW8lCpqrF3
YhWfjiic3/HAQJLUApWBpq1FaTpwJUdzHOo1IDpW+F6fsMYcwnlRY+HfmPbLEdXP
32F4Xd2ldSPb2shqEX9+FRa1DyqXdR3Ru1mN+SUUwEkpuD9Xev+pUxyDZqRcl9Az
ROWDC5yRr3XGNfv7oScfu0rzgLNF62CvOYHDb6ognvsrRR8nDjpJoo1V8J2EUXuX
U2/e29kQ0NytQk0jBPf+Z3iH9U3ufC/xI5Y4+CkrymGR9nHmC1raUIYPzsYURJS+
mhUIJGyukS/PImARmdee1kPhl3rgBA0aBYcyg/b+yTwE8czWvVM8qt6bajUVz9qR
552XbSnlW/xUFyVhI0S1RrzASHS9XlLyYelqoWcuGmowpPMYBdTB8Nv/+S4ZlU65
XPXYdBYtQuxouVodPyDsGxH6QnNrrR8Nbksm/AIyKLwoVQjqXczsLaAMN3BOIBs4
chmIt06UxinpZcJD/g8ttHwhnVJt7ifobUwmA+vfafNQ/LUKFO6qg3xij+Nmtgml
aj+igM7b/ie8aIaA4mpSRbdJ9c7pbTKd9oRv3l3A0+y3n0FzSMEUPNlZKJrcAWBQ
JeAN7Iocs7/WyKap8vDPk8EFidEV+qL8EQ9jgUuW9u3PgIhLBR7GLxpeQwU1IkKn
kYm356iomiW5YtWwsWg4ZzqRUASg+BVgSwCh7llA15wJOo1PH3dd5y6IfGvXgaYA
q1zqIA4EPFWrf5W30so16WSa49TINgLzQ0+amb+MNTOK2CPeX5Ewn73meAcUkahw
6zZNLbX+P6LHF8fFVp5ztAvLaT7cp6KV8zJ+m8SxL/OJgyjz9j6Fixt/CdUC4NmY
zyX+SSVbaH/EQxdRDkqqOu7vJLQB4V2ofM+2PckYVATmUy4Zcnjb1vpB1YK54Cwv
bWSHVvndmVDvIPD2JjB6t11umBV8plikwF+4p+RLy5Mip3d3E/V6xM0jL4adl6pv
kTY3ERaSlBGA74ulY9+2XA72Rczd4eccRJwU0XRtIcZzIDp1a1Lf0kk1hVKEGzkj
HL4LDNlEyL1/leGZKQRuWVWmHGF6q2V5WO2rs8Uw2EYcDKjFRDJTqsAQduUOEoh4
VhJ7Vda0LZfQC5sxoF9TB3MvcIk6rD9mVWFjFyEMKdmQiHnkzX+cwgQ+jngOPVzU
kMbZV8/QP9G6sZa2vpqQxkYRZGAqlO9EH5rLsPzw7MAEWRDpM7aXjnUL+frsRjLu
GNXEjQp+426OUjjkiJnG9M6vzokhHUWPMzhB9sd7fBfxUuTnNTkQwdMCN+/FQDVq
Zk4YtcXWwGY2aBVPrM/QfNiH1UEhiWI2cfI/Xc2kO7gGPbRXVMUFyutXz/YdQw23
ccxouU6+wFnte9v8u5YZytB7Jsjs8C5tNUKTys2ZG6c9zolpAdk4svX7XtRACsGD
IDndcB+08Unc18uGnMV1krGwRBPx3/OZjSj5rViOfNwFbpqapFPoMOqBfCuV6j/I
nGWuK2sEkiCe8SzoF4wbVW+IaXNrQvo2QRVfHcAyR2mF07CVsWSAc82vwakLe3ps
iPhwchJZCTpI2OMa3S1/C+KuIwOcR2SqcRnNzASFwG5bOS0sFawGmHT4uMNMqLzH
1ckakSPPZyJwdeVhXlsVr4tEX3jzNisd3cYXH0YBYP5X7/CtBlzzeJq68RKdQcfM
znREgP2ub/SaWUyXGG44fYNJljc9vOpWBlsDmcsPV4U5v0jg6vhkAbCdgB2JyaJc
kzVnUVbLbM9juBfRCjc3bqO40AAPtypqXua7IsYor4HTlLXeg+zvdAqTNkdCWS6y
ktxtZymLb6QSnmw5VvhmW0tZ4h9dOL+yhkxN7LabWm8UJvk2UFjtyznWcezLB8yN
fzCH+iMBpZmjNfFFunhHpmz15NAvPnsg1JepqhSLz0EJJ9Kwt71GsG3Z+efshe97
KQSv8GQcaQiTcCWunBYXVOcyN/zX9ZyIz9Nw9zC1NYT8plt7QW0K7JuVnPntFMr5
C8iit8n95w1OOT9bM/VdlclEkF+xAyO/Aq6QE70g0vbQ1lnGbtNS1lPaILtxGK6D
poWaZk3PzbJ4DtyRYjtiuyCSRZnSq0ayJP6JmU2O/sJD35IDzf0bR/sLYsPMUiZq
xb6ZFraS2IDjpAq9tNv0OWfudSFBmF2UfEgAZUh2Q0jVFm1K86qmuBThlG7U0rYI
sFpAFDW8TU5Di6LqYNw8j3Wyo93RXiw7KskBAT3ekk9y2+EGGi/hHoiwp85EA1Gk
hjD90kBI8UjY+ndSiUGlyOihTot398FJ67SQ0A1jP67EWzOndLZiaQ/67SMHCAJI
DL11gTaZOrakYykWbVL7zGjlGpjO2iMmwEN7t0dJ+hKhx1JIqr3yU/s4VBQoPvIP
UgUOX+dLgYhbywshTmlQpTsUgeRSj6JsEmHiJbi0uKgV8XU1g2s0Y74UpytCx3+J
ueb3J8LTyF1RK6XRTai3ELnMK4yF7z7DNz7WkTXtc//F+K2rR+nnXiv4LpJAkM16
APPfqjak+wmlnJoQ1T0XtPCfEbENLj42JpknpeJlT/N/yWELej3PiFr0bko761hq
tjOKFyr8yiWB48JtE/CMn+xO4EhR1rd0c6g3ch1mj6IPkPRp6WJ0OTjfx/5PQb+e
BpZUxSYzZmXXXovM6jZTwLHl/+kogczPHD8nkiwNdkxHOTLEcC4zKO59pv6mqEH2
SVhvE9IWuTEU68YY1N2aiIW0wgK6+EwbUbDUuPdAeWXJ0uaVF+7AoYonR5yquWs9
PN12TfWGxHQBaoZUmgThRbWZvMim0PFGESU42GXK4xHTb2S89NYztCR1/dKQtibN
cabzWW4oiPfkvn4X2nDb59IFkDLwYL7E2T06CTfxt44TIaK7Uj41T4AWfavQsZfF
JT4BnGnVnG88NjFM/XpANli2TVWJvoOZbbgmWe+DZMzaxj+2qZm/mMLofsXN9h6R
UiUvX+REcGlCOxRCnS0nGqRacwJkwJ3PuQZ1dGCyvikkUGeAgCozl4D5yKqTvsLn
BjEpquj8QoVCGUVbnTdvpfy1oURzGmTDMKINzIjIDCFufWKB0cb2xbbm+ta12Pzs
ZCFQZk3unxiI9A59QDGU5L9L7WV55AtGRcEL5YBcA213IdIhr2+ajCY5BNMrH8q6
VZyasAvct98G86lcw1vKEAtEqrLnC95pKDTDg525vJ+HtVEDBzbgStVnn51AWkNB
GPD9UeRM0uZagBpfo17zBCI6bXJJlxwZ/DlWSQkXZgcbXE9P4DL78DDB2iC+cVKC
GPDJdG3v92WVAeYQyx03X+cZE4JCrs9S3RYSwrdJFQBiu/qDsv89hrFwwmaYx9+U
MZhNSWhT2PylzklQWvLcnvVpFoAuQkT4mDdAqNgPRhb9FqN66Hhm+S6bZtwpmMdg
l5ZptxQvZnTH+y8Qdva+/aFEHc5axeq7ibpt9HeH1OQQuBLrMkjNVSIxLI3xopUl
S77vX7lGmMS9dLJZ203aIsTUjrIUbYgKAfYZdIMFyqwE9Bu2K67AWWpkRPT6dL6O
+Lo4Znx9Yup/jmfVypj1vtrkmoRj5GGt0FqQnMmq5fqzW8L+tl+jk+ZPULmBaVRM
BZj6irrqmf8EsbskLEYOgsGieae9K4tZu2qkzQqG2q3G4brTKkDt4HacyUU/Oleo
lpDl4lK5iaMZGdnAcwp3/5aRl1ChxbVi3N1QTOJoCK1PJodJyLCpG1aEq1zFwuir
ehy9Vs/P4MQxFEbdy6LkL2t9iiePHO7/XCiKjRzxPXZ0KjePkt6UYQQGokqOpDoe
/Q7Bg+NVEgZUEbduYfvPSzq3iodxQvTgZroSssIWb2DQeFh4f9Fk7uh5P2K2EDZs
mEQZO1mwpn6X787dGR1l9iu0Pa9WX8SGGeSElWV32QOFY2i+Ylkhvdav5zsJown2
7dfIC4KlpBQywDFREfFyJLVyFKlR/YvzNAwdW1QJo8J2vIGw1eFO3f9HZE5RiHdh
sGKNNUkEueuymFYB7mGn/1QocfNDygvWe8ECe2/KTeVNt2SftwoE25ghUcrb9JFe
Qpg3Mi+QM9FJstQXS5Nnd0pc2UWVYN4XcG45EyVQOXaU7mx/fgxTz1rLcbNgUzYA
/0O0J75f/1gxrRanBOAKVA05zYXoMk54qSDLK3QV9G/sE2rtKQ5oBf4TbaUOIjM+
tzO1Nc8PC+bNO9nBi//i3bshxY8xP53GmP/Oe2TD7FH2peQVLc7BenSKh9AlJVkg
6ERCrIuGFnhHVcqypbdX8+Kf2jTd26Shobvbj/EuBY8v8CitbouYCkjMeWTmF1tr
MMFpT6RAE0OESlMTyycQDUgOAxWKGSC2ERz9vV9P5a6HikQKNT47KF/flYq0V4Dc
FtWdYXd/1GefRx3om6W+tEDRjxOKWIV8rZ+c4lkuhEGmKZHO+1qbMr3nElyRiyQR
q9OfXSw2S2UOlqAozj4hNXqLVCsXku2NGET9T1pD0Drf+eRmetJHcOUemVyrB0lE
olTgxEWmS5cb+BFHYbOX22p2cuDnzLG1VmEA2VzzkVbEQXU3k5rrN0i6NzDgziLq
zaih85fMlYa66Xn1o0sb7mnHkxZCerXa+Jp0FA6kgXhV7qyFbP6MsNv21lDiax9G
PCPjBLr/YNgKjmDBl/T/E+QYeOP5T6TaQ/BkUzacCVaPV91jLk1BfVws28IOnkli
H0rfLmjdnspm8aeuYECKPHYbuRtmDFJe9cQ5poOVmpKT9k22Hz2sZU54Lz5mlAsW
wBbDcbgahsjjOnGs9EptzIM9IxXjFisjQ9+DLoEmq1MuU2K0HVGp/ZURWC/6ycZS
0spJioPdKarPY/YH66BjCr6XAppa54PDF14J4kj7vaHjRgmFJH8SsZecnN2RCNvB
vYx6AFEEqxgJ01StmVabdIUtEv6866GUpvm4SJ2v9r9P4fnE30KKyIb5d2QfIMKr
XEyw8M3GCQCQ6qQsKFnN1FfKIZ7F7exVUDkjSzSVgw9PPHcZMl1Y81nMWhN87erK
e1BqIujb9q/3ryYbW75dyWPncrp8wNbYzew+sV4KCxYtAGlUzFyUJIdSgdE8xTMB
Qk/oESuYZ2903kpnF4tEfmgSAYouxNpLUlwpMVabrfY6eMa27Tx4cFCVJ3qhWdFm
9S0MSbDbNQHjgQAUKozFK0txuXkN7xqTjXDjojKSjlr4DzISGr2A9mpJkN6CiDGc
QR4XdPleMEE6kwU/sc/JrAcPrJ6nvdVRQ0xhCxnD2zFpqWBFC5JUQNR0+Pguud41
+i78yrvUtl/L3b+Hcvn7id3vm2vaA2tvXsetjjjg6w1EtFaytfTYj9bANoB9CTMz
5kugaA97EJcNkluBCk4d5kyvG3roIrBHNRH7tboBfTVqtOEIlSDeWhuOv2/vwtOj
QAV8bCauDe3b8Z1iF3HkpUJuHh4P1s3FD7uPUzuUftRFqrbzVk91qeEADomhH3Ui
Qc7NUU61X8gJ6n3Hza8frbaQDq7SWDOjd62Licb/sMI3pkgWYV14kkfOj0mKP63r
pyUQzOK9zEX2b8AznUn0bcrvidve/YMALhB1oJxpvwgsNu/n9r7C8u3sUUQGUYYu
Jc5KiAvuBtvjg5BvXX9jIMYxzHQg1crX/6nxPMT7To8foSaJ+MSeSuNa2WolgLUK
BIk2HrFlx3fO2WbrYG7sNAsGUAE2iSC4+25S22POwI37EeJVlKXJP+Za+IKnweL8
n6Ek9tcZONnegDJRy+d8jMhVEIUyKfLc/qy4FiAel8EdF3GdTDStuxsTSjwxvzwo
SkA81fIE3Iapz9y6oFufO/FtrBqQuKV9y1sonfu0lKNY5K6ncNS0nVN605KPtBIn
T+u3rSZPWIzGJqitTI+Eia23FKXjtAQgnIRj6sgb2GaiASdnYi7JrvrelMU+RubU
zII8OZ92Or5C0fYwIYnXs+f2KpB1xgOZ0CWEQaRNxS8cP3AQBpdH9nNzYBlmcjU2
M+MyF0kV0TAJuZ675SutEc8s/JyvmecXH4n1+u9sdAC+vbEjx6Uo5vWEXBaGdWiC
2BiKgPIKlq2zedQwePByzYAYer4i8kd78SpG/bP6zYWSjnq9PrQXtCO+LwZRNq2V
Y3/XLYnW+C0p30rrFbaeXqg4mYJMgwkDxaaUUecObZXE3BJOuA9lHNxrbK+8+od7
Gp75ioODr8UXwAGCMLjbuLE7oExbROQJAduPh9A4NiMPNsD7shbHVPkXjIsbmqkq
Yq6gJexk/iD1339TEGx0d4IVcloaruPlXc+Wammf57nycoWAIOV4GuQob3rVa2ZK
veUdI5Wwg6Iz7BT+xRZ7TFVgsYswD7VwJikLFlcJIBxyv8GJI8pxjA6gDbsrEUqZ
qkF6f9WO3Cq6W4kbF2THIDywU5BQBg3ebPEHQEf7erFUMJwt2J3MKS+R4KSEjOyx
bY/Go2sgPejn0n6gmto0jXl8HGsoi2s2bnVss3I7HBT4nTCBhWMomYhiakyCrKlu
lzrlWwpm4HFilLqu+OnYduhRLdsBf0il5rPTLxdLHHi7wEw1Mu+volpqiKypMdw+
ORiNA5s1hxlKBVJhPpwIOjXsSIcWkvoPBF+89AW2EgC0lH9OjLjuIulf8jF7t//C
hf1/J6l1FJjQrK6XzlhVheELdhhbNlpirM7q7QQXlpVrJ9m2nmXUIrDn/78oFjju
l2jiM0JDyC4ExHB0yEucExgtl+Rx9LZsCHdSX34uklld/R0tmWlFzskoE2GqT24f
TQrCZ9l/yWpld6CdjAXIsFDXUreKXRyCskoeVpq6zLMWMcpLMxNCCqOeCVysT0q2
mD9rIQHgalQsK4apXv9VyESLSdS3ieP7ia0XZWY2E+EWd4PrNC18u7gf2cpaKZyp
VHeCCN2DdIByBxsNc8gnhNV/GfzXk91SaXjS9ePCvnyFvawkp5mQojtB1+au8qEd
ZzICeB92mYxLrzj5H0+SnZweA6x2AjFdraleu4qbe2RJjrsKPPiVt3ttGLVeQnXh
D9hIZVIlXLmESnaLJTL4+AQAezjBdV8WA+Y2hSiTO2bJi954KtjjcSGkEi6ywpNf
Scnu9214hVkYP4Mg/34M+PNgarme451/W2TqO40hzawiMEeXe08wUUHYuTvueHQo
2i5wQ9SznJEY+WZuAYI20G1oam9JFy+VT3D/6WAUG/nfWrTzEIzjifWUJP2kmhMJ
3Lg7IZxIZBmV0FzrB01PCNDA9rFRPX19EQtZIP4RalQ2omi1pd5pnxWlQOGbM1IM
Dcan4980aNu1Kt34xQz8FmtMAd0RxtLz32SyWkMPBx5qpq1CrPUDuOwDHtgMVL00
gCwAOn3OG9wE0VuNqqtcclYgXWHn+ooymjKuAs+8PIDWo/OZmrnrjrzEs0Mmx5Fm
FORmeiPK5ikCkA0apGlvHWrSSnLXf54oIM2aVVVtI5uqTkDrZSPWID82S2h+Q5SP
hF3mm7s4YI2/N81cV5V06SmWUDoZSmc2boQsXCWF9HgVgFTZFD5AVUJQEWhNJLa6
XoxHzrjW08+dKlfJiRGrKPcp9ke9GlwXF/mbUvA4vLBUKgEMRD7jU4qp1OI24L1/
TdnLM3+S5Z7DwVf9m3WHwL55oq3xJ7uxuBnu30uyeWhHXk+ZmxVesM5Wjn/1C3io
GiQ+sDL5kLCXfE9uwI370/4HbMsDJDxQ6kAUBFM8s7vu1cRaSUc7ccLNimxNVxa7
iAOuJd2H327kWo+5Q4kaSCyrVs5OcNUvxl5lOKRQtSXoeSNnQ6BMQ4mRL5YTInE7
LowrTU0m2Y1OAfHjlGnXgPvF2lVT7xpjolOQhGYEV9ZTopZQTHK+Sn0GoRG4b8PU
mXKCN19RYy1r7m8hYpRxClWlK1cL5nx/RVDob/GbUmhXE/sK6fbaJNCSOD3yQBAz
HzEEI5AxF4peSG3XL0gB/grFRAiTkh3eafWKM5fuTE1vdzewP6Tveh/kuq1OKSy1
lnduHAA8LJ8jzI/VcPkYCz4e/5CuD97Z/V7o42hh580+0Mkp7Mc1TXdRYcjaanJC
JOQfDEwS+T/JqIDQiRmYtjQ+5g0IbcRPGWo70eF4gnfnePreaPAo2bKXTnHV8ejA
bDxmgnyK74aur6WbzyTjXLQiDVhXtbu87pmiricjX8XnLmKEfaXBsa6hYcPycKQL
3lzelX/bW5Zwc0BOWNQdME7J9pFSjgwh5BJaKUdIPegEz8Y0hWiG2E4OX8TJ2g/Z
a6xjwVppmBvKJu+MzeNVzdkuAEYh1XPQGT1MkZZhVo43h1/RW2We+/Ye2ktVheQS
6qAvoIMfbyEdQ+IVY9fV1STG28oCEMrnXlVQCWm0Sn/xOTx/+Ugg3Al2k/qOxN1o
nK0kKLzPLjn9Ox3Dfg2HMPJf/OzRWwVp1dVGLtIoRBqer/Kza02SpEet3hurIOh7
qnSh7MZmgueos+9Gls2VXK6Y16s83yDLugj/1XLIIPxb880d7sHAlgYfAC+3sf5l
1aFnAkeJTHgh26ReffFY1BRxOOi7z3DZXBwgfYmDVIq0vhknznv5TP7p+aT8xuRM
yHJtniMtlVRPvFmyyXSvw7u3SMnhIGEA7t8QIZiszFf4bwvDkkfAQMjg56A4Ef6z
4CN4e18OMEEwsGIEpIP3DIxMQZq93759xoIghLmoqz7EECWdJ/NxP+Dosor3TaRE
EO81+p8FA3wx8cwDDqAyNykRtFtMxkUPs/AeNIYBCEWzersSSPhUKVrE9cireoNy
K4UtQEbidbXKFAP74INBoqhTV183H+MckzL2zei9Zwe+sEfr3vabg4Tqc5Sd0vMr
2DxEmwcbC443Eca9VF2MqoB72D4Ctr+uHCqqwIrnOw2FSbhUarVi+4lkZMFxm1Z5
jwqIWx/EhNNaetXQmFfUHTkd+2K9uTiY6FMNMkPlrUPu7Jzd1EfD8HDMzQUtlNH0
IZ0liu+c49tbHozvA0K3QjlEKguBuMteZ4dVXTtlW93+rN+azvJ45S7Tgw3oIxHE
KYKS8gPQ+iE1qBgtg1Nsw2WZch5X1tMR88n5tXUw+JtH1dZXvZXGYC98TGe0sCPp
8G/d0MuS93HoS3IkWZZto67JfKRuI0i2HiimUi+JIhF5AGpOeNGEusVVzjnXN7v+
NljgWRAF4DMhePdKJI9m0GToSRotqeFNPVKJigDxagz20/Riez4Ml8aATkAVk2HE
DQOPa3nPkHGnqvwRbBAeruXOex10ClcH/VF79UUnsmzz6GpGIqIzRqkCY6hjfyCB
BH68lIBZS4iAVEUzVC3GY0igMOWJB6a2xoGGHb+NfA6GvJSigxzgsWG+2HFv4+Uw
SditeojbKZxs6F8WKeG608tfD0NVydG63tBSmpbEk3RVGvdcbTqEVrsvDuGA0cGq
W5laOTIy83TPhUa9vqoFYiumpsvyrw58V7N10Cl3YE3iDeRIcXJ1cs6vBXmJJTNX
T3HkZ7/EZSNyO0MokCWdnpLz71WWJl4n4TXUq+FNeHhMIwbrPzRnGWnprZteil8t
/vaveLqXjaN/rmULylcoC5sjy4N88rJlBiAHfiPKTnRxxhsft6up1ZJVdmlA4hLg
XNuoq//WViSKdJffTU56UUK73mASv9EY6FqdPDFCsKH5h18CzTOj7KHaqHTlMjU9
kzL43mL35ZjDIUWUa4wXrYbGkCoF2feRiJiGoWoYucI2LgWj3HuXD+3tZJbl/waB
7dkpOxZIPpxIplA3rCxKnZI4b4vWU/F9M6/4la/opoTIbOJ/ZCmQExAPh20Xhdt4
GLh2HDAcikRNeKpwLYmNhKGqQjo6YZAofU/Ys+3t1OakrqbmqjgiBcdN4R/TFzRj
SVr8XrE1n+PfuiolYHNiJSVBFh37eGzNtcupoYvtlSwTdP9cbLvu2pKToL6+buG3
/QzZ1DIt7AmtR6L8DaJU4/EdDRvQ2scgoCVnCg6GsKNBCOML2OcnB6t9OYLPMlif
h45Iy9QVj7hBypvjNP3MueDupV9juL5qSvx8lGQOnto0iWEwXtU3wnccqWuYJm1h
pPlHOL5dvY4l5A5YKgxZGVYrTdlzzCnbTXqQPw8JHxccqM9Jtbw6rxLYlMbNF0L7
FSFOvEfMVZsYToU0F1oBn2NJsjkc/MSYenYKiR/GtH8fpLW/tHm3yAam5da04laM
XseL9civVi1wArc674WvuMJieUl56LaUyLEQw3wgxUxujuVZdx+NLVuqgM0n9Ov7
vvGQ0vB9eG0UBgOf/S09OUFIe/or0H9jwBIHW9ldQYOxgWhoGH3Gob2sP3WCnNFu
ybi3rwOzOty+eHeUc9o931jUqKkROnZKxBxBohcwXC3qKp5rBMZXbtXMPGoWjM+B
GOOCBBVrx6NaDxD2cT0/vyw5MWBnFxjYr6hYLKgfEp4cvfYlDpeJten+EXFVqZ+B
pj0VFjLrJcfqsP9rsHy1N3BaKN9pAz/ZNXHI7AzHYy2i2Uzuh8AlpEjxm5gEBEJD
3SQNfiUBVECmb3LNgp/BtCCSvOWO5m6T99w4RNsEs6w0eO37PAQY1xpN4CndcKvP
vDdzgwdzKBOhgA85ntBz2dp6ZVdT3jVgE8DNz3oCACBS+n+nYvZz4eUAyFLeg8mH
QSeRozSZHE//oGiUZnc6wvYgkdyBysEjzKvGNdgxwyvchRThKntCNmCRr9dDMR9l
D9kA43Zvy44O9wV81V4IvNbi503/vVAV3zAjx2LlYkalz/riyI1fvb1jXuqdNnMx
g7ovkmdi0t+hdYnLyDZEeNYApw0t9DsaK5S9KtA30HNY1ECrRodN81B5hOqREEDY
WTwY7p5ZVFmgOEddKn3LvEucADH8r/ARDEmCpYcn9Cfa4YIQ99Z6cr8VWWQbRBJ0
G0ZMLaRhVOaaaeyiJWi+Ls/EE4PXLpJ00oHHtzd3u5lvKfwkOJqZQre/T8cRWvSp
PuPzzSB5CXT/r6D/1dKNBC4kwyuOrJtePcRe4mkwfzK0ndZpDVjGVJEPGxCmA1iA
ocA4ghXE3MShizTMlb+kpi9WugYD1D1K9Ij0fHS4TGMkCGxoaH3KAzUP/DB7VKIB
b8Pv6fv6nR27QbU2om8jctWyzhiysUXSgl93ejgntrbWZ/E6AglA310UZ316Qcgl
q0BP3d7PqCV/V44cs+wxhMhfeIM8Vr5JdpzKwuPVEXFWW751KHUVG920iC/A0B9f
2u4bMsYK93OZtiCfoVEKi+3j2lzsnH5Pgelll3Yfk+FpUNXqHSYGgt1B1ucMgGaG
2mcJW6RzlqsxWxl0zz3Q4goXdxE9ehIsnt50f+irrlIqcjpKfVGb7pWn8ksb6OMF
Qt2RQQKlJfArndrgaMmIrofoP50GO9qM5CxL1ppDbjTJh/xE9Co8LQfRXIfA9EPY
yINAw4SZh5ISeSso+dFf3efRNqC+ERChgmP5lzRs5ER0xrYfn+vwpYctQsegTkx2
WjQJp5XRuuv7vk4aZlwAotzuRhCQsyrZg/I4++k70orvOGFQQbH/hcOqUfmC4wpC
AP2MeuhfJWVYndVNvZrLTyNmjCEXCe/xLxvQGMzwcW4zvBjTC0H4S0oaQKb66MCI
iv7Iyie1eW3ljCLxckDWsU5VIdSbG2psmArU5x/9ErEv51flahiNBL1OVZF9eItx
dfOhYdemlnV3zzPjjKI1npLB6nrp9/2JNkic/x/8A5rK8iA9t3ycfJrhR9IHL6pk
061gt2TW/1cajBnXuMoxnnbHY9DSKTydev/4Wb2fDHCWyN1mXhxDuToly0dHxbXK
qAD9WjyDjL0ioTz5A3w/nuzztC1SO8pfq/cGNH4NHuBIA82Re1KumYvmjrgfCKxK
hoE5i4TxsLh7nkk/LfrT+hzKi/48dH/TTRkDZzdY7F2yD3G5MOpSgdVVIO1hpQLO
/ghDqAw1LAAtOMqdOWaTQMGX6LDty5HLa2DYk9MCWCINwydOMuKm+DmQuqoozcWP
DC72es5wedehXQAKFPG6U7Vyd374f9PThMkpb/qcHoRnbITBWM7xf1xFhXsUJJ51
a8ycNCzhk/TZ/29sSFtu4iYl0Zbvo3gWiGWhLxwyFjy5Xm0f07rF9Z3AdOQ4k2HG
gDqZJWcr/7UD7hTkxsoiQKGTSA4MsBPLZc5H7bDhL5mW5v/SXMecOlXFWz1aUQCm
ZxmzFvOtvcbmtuFi06xsu1P04itkRhLZukaxrLYQ58cGDheSqJfv7Vom+1UERZP2
7GxNz/uv01cB/u95YOHDTgm3HVg5eIzZelT7xxPvkIQYPylmEocnBGWlsQUeA93M
MSE7JDvSZt+A0+KNkkPwS+/MBFQChodFKe67nEWB8Wf1PoW2ePr4Htx/Nu1c3FkG
RgJyFsmJ95UVB5ZW0g0b07A1hmySHK2CUi1zuHt9UCGelTp+38YFWaZ0nRK4/jna
EERAtpwlsdV8y8HIwAXh7BeJdqWmx0+aTQa5QNoUbIO4TLnxTDVw2P74bHwAoGCV
aUqHgzRMqyYGugv/RMjbhEVh8GCoPxzhYhTbwnqxDMxrOPzLxNyJuGDmiyhLLI6A
XC+B+DZ2xk8C1JVnDJZkPWGemAiQU8HrAWNXjj+VogjbaY4tRwc3OwITLhIyg7fp
TVTivpqABEOGyczgTMDyN72Ga2piAtkPdeP/yAtTHNrt9XLYRcdZDVJBTMO+1W0V
ARS6GcAYvqcDhLR1XYDUHGkDp2K2eBvhZI9BCKe2/sAtbqOQACzbgY5i+s/BXiSw
+Uf3RIvQW3/fe9cDWIGR35ayy3MbK4lZZWn2tx/txPAmH9rmY/bm4KaNqDm54OjT
oBhp4z8Bl7QmchtKpDHz9GB2vg1uf2as/wpKd0+Jl3V9xNyX2R/Ry3MG60GCK7CI
1C11k9U+D2+38dJjwZBpzlVvtKRz/5jtX/lkAaMgBWkwCF8TxVFdWtMqZvtccBvi
tMQitBNrUT4z8jyfeCGkY0alE1cYbeQEvM5D6EzrPVhBqgA0q/ePuVo9pBLkNncU
DqH6D4TlmVotZzvQvLdjl5mIaIS0w1w6JuztP56j7+u6xrLRSF+hJuptDn6Ii3ix
0WLP6s4sw0rglkKF0xEQQCLWcwvMG9t5UzLfr34+txJx0Zb9ieNosW0SVX2y3v9a
iGQXBsU+rEXZckMYmnFawnlXDxfQekg97lvE84a/CjZmVI0r7OhSUE9xXgoON7vP
076HDWwv1giJd+iWz63ndFyfkUAynI/TO7V+JKlksuN9o4XbZCzYfj27fzYyR2XD
rgRpPWCPiSxJcJObUPEkUpo3kFqEssXE+TVzc812/2cQNGTBNw5OnWWj7WiGe6Rc
YIAp/XZt0VtBKGouULn/zbUawSBLgxSc4VBoDngou+/ZWlB6MgD/oN7bBrzpWOG8
cpz2dYJEWIAPCZRGMm157OrykBsjXV/cwtQ0CXM68mZcmlzxSQOJgPeBqJ/kbuCD
/PkF816yhLJE6+LgQZseX9arhRXb3UM2GNc/+9z9KwbFlBqRR4rUEqDLUz+Km840
g6vA7DrlRlEPhgE+MYboHS7BL89t5NxQeYzNjMmjmoQrytd+fRwHZCd7zKX4s8b3
vb95z/WguoztfyoGyPnJhmOoT/3j7ee4oDFkY0Z5CJ3VcJCKu/hPwaP9USIBp9MG
kduJhsOUm/iXH71iAeh1nkg+g8GIBDwwUswA8/ehMzBUWYgxeTsV+iAw61Kh4G15
76HItYEOuxdGOXY5kpK1l0ECfGPykhvGvHAJcLHwoR+G2FZPVZ84laFbic8N96/0
MMzQOOwTWnnz6n8zSjvElUT1ovXYPtGIrn5vPeWkwglFZ99NXV2gv8bGt7+P/ovN
Ao3fpkFm8Eofx0TvNu2BL6/pnsgukZUDzOsPnygYNhk59pZzQl5wqTTDpUWJHYA+
rL73VlDH4Cl6wYcUFTEn0xtPcjpkcH7/ozqF1EtR3pbkMIpQn+xJFrLUeQsxVGMx
+nskGfa6H33CoF/qD6AFX4OP3fM4592kWGyJZHuRcaXIDw2UB4SelG7/ZOBnhDR1
cKGEdQkiUsbO/At+tAULjHyLS9i2hOSDwqMedN20u8zDYj6Tn5TDYGNKanzqh1du
ejQmPw/EwnXmyP9EOWe/BWFLJsuyz2ocn1VyYk76frmDfmhIZkBpEwpS7kLYmzOR
dEcHDVQYG4xSKSfBJoYIE/B7gqLE/5Ibu0RRyHdMpg8SRwdbF5sCwa9CF0s8KcU+
JGcqsTfE2VUpWRq00FXNhaRcB4tjrL/rZjwvD2U3qLfCN0H5M2XJbjH8EMgnsWsi
smV3Dp87DKv/fKEec0/IL8El7S39mEQIxy5QGdfPXLgHW2Q+EPRIprmjWzAeMHNr
jkqAwYZr6nWPAgaV7tImtASGYiIdgwMe+kiQpOcybRzK/ZvePWsrIreQsFxmm88/
RqySgD3ZD+III2M36llZ9ocvxaj222iZIodYr611qjwomuEKhiyjkxHFEM5hCnGp
x7jNYtQCLVqAGfHWAAdVh2lXAUAhz1EcrfjMSX0wmAMbw2mcS8l4H1SBqmru0nlQ
sEJ9qkrZb6H+dNKICuSS3dSeeLmSjzB+z9cTaOWqURqsfrM6p5ntBh3AcCni9Onm
84jFXzUOFtysfFgtliUzL/1L1IYOGhvbWr53btzYrS7m9IAcusFMljIu+tfkRzMX
ZviK997sC/NFcvBieOZiOgLcBl6hmbKUAYRmk+H5l6WqKctYVlviGkl63abqSZUi
ZpjD+3hAomYC7Liqiu872hp+P2XV4QyNO4s+Njt7YutOdqkPVrUbYDH7YE2xgQRV
vG+/V1qNRV5RVx35h3tzGdtR3OuwMVc82g4X2JpCq9Y9vtl8SIcJAvbeWNtdE9cK
c+xUG6W9GZGcEENQdBTPzRtvCIbVhFVBJx7FCvKsrJ1H2OuMtPZLBNlCRHFKrJvi
siQkNuGrts+NMTTqZHNsXXhUJgblcCKx9KOcMQMzmXDlZCFnzteUdbK12zrK6onC
c6qp2FLmb8LOcn5pHU1it3a+evx/fOL9Zsyl2Z/QC1fKTx3bs3cAY+1kOQnMq6u2
jaG1cOrXEBEuTE4bSBfdq70Z7UcDSnFNwThqNVPmyBwKS8ISXesLWZ+MNCXCTtKU
Sns0QKVia+XJOAJ9EhrX3xKFUxKZvVAdkwhoMswrrEEz588yGrFYOeMtL+j3y+qe
WK2vdNf+ZyMxNezg45arTVGobmC/vo63+oIlqgRHgu+ZGvHIVmrjiO1vnnhqYZqK
zxvP5XrzMDYZVmXWE8ejSfnk0vUHIhn/d49PbWx5+B5JRZIHjpJB0xUwDaQ0F/1t
j5K0JU7ERpffLdhIA08BrE9CgkmKZuMQ6hXJcSLu3WFXF1ZWuQ0iXhcFx5fWEnFE
M/k45lNjunBe+zAEJvfUYNlPEWkrXWHNiuqPfkkB8iHGay7TMMs2wAFaS1ykAIwd
CLRaqb4lKJl+ZewBuWDpS45h06DmZLGwd5rdIwTHl+T0Q0nw0CYld9+EvmlHZL7W
ZsAWseoQDYNZdpnVdPM7MOvg07DWb+M/anvQTF1c+xHFXgYMeonfs4UT2iHttDJv
is5AvZ6eruFAcsL+7xxaz8tY1u05/dieFrBisTCojbmIgWuiD1mpoxXFKpXZDez8
x2NKyaIdZ4ttggdjFdEqpr+9zSrSU/oM56xfQG/3ycpZjz3G05nGY8dATdFkqXlW
pfG5DjxgPWZIwbBEUPenkBJUFnMlQs4uHNWMLAIwPgHGp5i7x7beyipOi74LDJxW
4i90GkF2VZYeQBx4QmS+XwRrFqSyE3KHmgO9LGVqrc7OfHSog8rriJP1JdQfM8AO
vKAY+4ziCvb4A9O926nXlbwqMar43eNx2s2Rq0N3UugXo+e/bZzkYbf3jhY/A/B1
3BE44GQUA0EzY/sn1m6O5uqv2FoqYjoshsPPt+KeqFao+8kHISdZXfWQ4k95TKDa
c5QEQq1+VAtFt1qjixNJjVOazERVUKGBIt2jwpfXTyseGD25+2OQnSoATMv20I/a
kz5gTSNn0XJPPmD3KjX6aPZp2Nlj+rj0D1ueEWCBrcQSo9LpeaKfapjytR5h+FtY
q7z8GLDJ/6xELHPD4Qu8NdQ7oPZWknKAz+9iLTdqDNAz0Klxgp5ThUmuN74HIIDL
vY14l2r4BtTiDyWmb76olRhy4z9WEY/kDs4jEsHWm89cJzvUsIYW9P6LeuT+soGV
LcHsXkNpJf3zENSr12+4cClyHnQNMrFGogV2/Ypw0ABgNPiUsEGp4hLRfeWhUEch
7tHlm06VGm1Xf92SwWRcwlNZZflnZUnygR4/9NPfiKB9P8SZ2XmEanLGdwXhno+X
6/pRcz1Y/yCqw6Wk4vYC6wHOtJ2qnqYBzDQTcfqfcr9tn2z2VVgBWGAKkJDBp4sS
EPX+6aJMQS5iFSGtmpGab76V5/V+Sbe7bY1roRp1d0MMrOJa3p79OSwNwTEwJ/pY
sqVqOn7auZXlk3O5yntyCUr8ZOdLMeZ4Gl6q1GsrrT+zZ0mcwNDR0DdIu4hlZDQa
8sF1sNYCtqiNsN/4MAqUeEcC7Cfwb7PuumgoCE15kgKOuYO0dmYHaw8u0sI7DAA8
XC6cj97s1kPJqb7X/pAUJOQL4Js8D9WzZUSxIk6LiVmQauXXyG8GGpdlfsSB1GxU
Ps1xFtRwEON2lAPfXVkXqB6Z38opxDNrl8LF36UgK/6GCtmg7FDh+Vq2kLjR/Lvn
r4xkYfh9JMOdCDhuBTTkIunC1uFMtICmPEJRqxDciX/TRJtVeLdrnXKzPXnafRdv
evTPAjngzVjY0kDoDbLz/153hHthjQkEv3IqjOWzu6kgq6Lt47vYAT9vDSIIl6Gb
+QyS02XOECph8rfMoN9ZaeHoDfYggB9ALXr4KJcnRORW2V6RhNlkraJ7IsPsBgn2
1/uY3r6eAndUupoQbDJz22ngQvSvVaxRLDduMTs8mbi98rJZTy8R+BVsQE/LRls4
28iqOqm/T6EuNhQKTUKK+D7imDQsdA5he7lDoCNYfkBywGwOO1zpflK+UJ+vLv6l
ywz/XFujPwJOqaQf7L0eyH64aVTF0QhqbtNxoZzkIu4tUEKM6+aSxIQNF0A2Wyqf
yOdyfih1k7/0dIjvjUbfokSDFQH2dSjuQj/z0dh9goSFk1LTa19fyYvj68cD8W15
KnscsVbZI9OXLaUplenlhQT4D+NhqYJXUIZPBsf69HRp4ztwhMVxY4Gl/s+kaSIO
qoOsV13LBQH7prYYU+eqXob3ovX5qa1St1b52apPFwgwlhwAsHP3gYXxuKcmXAaz
r8obImRS3vzuAx6w1R4J8ZmwZ+PRfXd/fitF2aiKYG62wJ310Rn+y3jYTLYuKPMP
cy58audqVV27Vc2+54FASz4K25ipXbv/Yip0m+KfJATTyb+wlTDBcPwRM/dAqqRo
+bynLF7VqQlO8bhz4lG8s9WbZL/HVXMYeuOOP4AmtWOpS/0mbGRM5e0hMELs6vs0
aMfTjTtNH0qNGrlYl5YwpQXlmx+ZT0pCU7555BYhXc97lp5VU4rl+NDJXoNCwpkz
e1GOvWTooPGFyPHQJMFOTUE0Ecf/mqEIYxYs++mgTl0EDFsyuSiW1z2ZFX6cgJDi
05KuS/nw+0q8qk8lQLvHpOfAvDH1ZmUDZqJUKJ5rh8MWE8SdCSG1KOondemo1EVC
n2wKxTtP23QSvKMAEVYCFTC1s8+sVA9nwQ5IBtBgI445a6ATA2Om2OKXi7fe76Ea
pDUTw4B0NR+fx8/aY5VlXwVamRnpubpfnddq4Y9CldZNIKUFBVf6hQOVJzn5UgFO
lQdTQdpoDlYqDsoLkY76x+0LTD3ekGgTQn4W4u9M6ILHr9fU41bcNfGK5tDxG/HX
it1H0IuecS3/2Z5+WW+m5xKRMs6x8GCiSowrC13KSyFghPM8k4HDEGlK7BaO4LXk
LBCwscpe9Atn4CwCmH8ROdJx8QjPXi1TYt3/Rww96Vnja/n1iYdnXNSWY0Xotifg
+fvyDlzA2vGwAVfeHXbx6Qte2zDHtlTL1IKpBlRDkHE42NYb51w8sGkp3dz2x8XU
yiPJM+CyZAUA3D5ryyqe2koAVLcsUSEE6drV4IxfR0J2WdOEHedFbczFAbl/0VxY
4zMeXd1bV0mt1xGqLCKPd2IpyZYGm6flgUsxCZdTTIiDQQ8td/D8g9oSO5YiWNGo
Laj9f1fJgvdrFumhR7HEUKlFYJIvef3Ih/Z5nPiyT4b4BgltCiNg56pFxlV7lTlL
OAEkVU1EknDtDxFuqBa8nNybsnVFzAC0uf7pLOuPaXxl7GZ9JahajXWjBd1M5d9Y
MeshCWYAarhW8nPthCqgub3JSBVcWn9xM49lumlcK1mCyDSFJVuGCbQD+9Or2K15
h0wI78InBlYZn6yFtfWz0w1fGjp30q4X4byqAGzD/lomt04pPljCjm+LqyR5mVGQ
7PhxE2cgUOzQypOCLZ9/6ocxL9Vw7dE9DU/apuuoMWbkPl9u7uflqEwrn+HRuLMr
h1d5Wwdru+aSgJyrlfJBYOwTNS40HFa2Qwe8YgHNnuxlwDSJRjPJZ/Yrgqu97FKK
853x9OGI2WFPuGI2beCoZ/vqdN7S21R8/h/lhKrfGgu3/Q26RqCfVa5X2Kz2wxDy
7V43ebJ+xctVUJAvnf8c7SBtuSPx835z38ztTRkxlgXpLI9J6rH8nZF4uoQmOmOl
AKSr2w8VKVgtjqYPf96DieWAbgLUVMtPp2FEG64ZrmUmceJtaR5MvKMRsyn0q4AI
ZNy9pyBTUAQh3mJ/D8iJOXkNQpKxrl2Eajye5dEdSmXc13pUmwtpygfKJr/muFH8
H4adiGOjWpEF/iU7EUIRCrUrkH31NTWiPgEn2SmsmtnlgBnFCBxv4cmSyBChtl5g
qlBsluH74Fk38AcZswuLDng8slMoZBhlEAt5MK1dHo/ShAJb+7MyHrM8TSUhCdzR
RpaPKsVvIciY6HdZiukusCWIft0+u61yUyDCaymvb5xeOyw46jFHMRD2oiY57H2Q
pIG+MtK/gBFsnBwl5OHiIFB5BcHHGacEEpMHOu1EBl02+WML7Tmhhn5ezC1RLLX2
SftntbRv++AnpHcLzUFNj+sZrh6HGCG5HpMdXESmYdfHYVYwxy0QSkbgfpWcaoQU
a/ofx9aNJzQa9YHsBM/pRak/rmFhMOuhhvd8d+Y3tIrmkzFLl+XkHVc+herIQ0Kf
JxP7Uqp1gsQp9TV0FTsZ6r31wJ/5z42MQQreLBadw9VBtOtzLDT03D01m9YasAKC
kISNxBU7Tp9rKlCdqBiVq7z7LI/Mwq+AS7UwJRktLdai6BmKam9PVK6MvBjMbqtW
F8pyum7I/+B4qdD/cQBX3h6l5l5GUrsFFtf5C5xSCaErFja/4eswgaqryAgHX0Pr
TbXOShQXCd62deSJRId39BwWHhIh3FYba1fKppP0mxoN7aR+JzkBW7gWNZ+tit+y
JVgp5selPkzzoot5zwCETLhg6JCzrtndIl+CNmLgWrwCnP0Ho07S83lKfBWsGxST
0+MkTgUhydYvxhQYe/NGFwCqbt5sJ4bNuCZRE7UrihUqGbxyYdxCpkE5atwgrVsN
gHWe2GSa4sg//fhPH8h4zZVU+ZBeHvTQPCukwfbpqfPrLx/oMd5y/G1L1aJQx9x3
DaTBF8zCkrGYm9W7Aqa6eXQwtI9dp4X3fiiLy5gGL/p/kqsSKnZcmJUHC0haWUJ5
8ruPnrwztvMShV/ftr87Y2XxUDuthVWJHEPD3cHSbQnyeLqOOkmBNTlIXhm2LbL7
z85lGX+477b+TE250kIU2yO0rAgNDY18+y91G53Q4duDgQ0W7rU5x8bs5Nlh/KTJ
gRtHvytIT9riflH8D+g+WEe9JWenIWqA8OIAEtMBk9fVRh7A3EwaTrzdaPIve3x4
BuGyJJCwFjgKNZduxg60gzzm83GRC4FJjSl4Q4XvaTQD0+zpzPqlRnV2jCi4f7rJ
zUugnmtAA42hnAaQzK+JKnb9zmBwfUoC9bXiqTyaGkR2tjGY2lSOOUE5h1ChgczH
pEM1wBBI3Jr3dL1b/wSLHSV+9Z4cKs48vN/T6L6rrHpxYOSJXbOsshMiuTOebInh
XD8E1fsBh9R1mdGAWy3zq39FpqUvHFx+3qLzAr69mXBld3TQec11VKCuJXtCxxBh
XGTpZOUw/gZTqN9nlxyyZv9eAghjOHDBpr+NmGcL4kmIF4DxcQnEcgJnXYZyfFl0
A7BYkpY1oXkl4s9EaG4Pr8ilgmvKhccsff7o2ZjTgqWVMu5N3LFBw0JGaJ2Fc9Mb
pGJuR8wwkCOmP4cXjqjt4kQd6GtjVQUCsUJ5o+SSkIUoBrzL9NM3RXujtHkGisQ+
nQVdD+HnGwqb5g/V/r7q8k//mPaY2sRH8WIm13F+AYjyNPwaFLnpL4hlxQ9G+41P
gJQXQWb0oC9fawc6i/gQHFSHMQuj3O4xUPwODLYCmHkVOsfVYBRd/C/OHWhcTxCH
tybCRF7rYWsOwqnIXm67+YyOj1ePPusgGhWgF9PWuseaOgMoPsWTxtCo0xQRHtr9
GmJS+C++QK9Nx+J6v95yxeovJhju3YJs+35ZHz39Wo7YlbV7hEIuOAAfGmwATQk8
uLX8cxF3RKVkUSgKxNUlrB2s6uaVgcvYt278acy2blBauqWSDtF84zl9MOZj38hP
mRAkrxoKKI7ScTdCjmWyFYjUhIc02fEkCwT1v/T16YVj9eLZpZH5uRN5X2SqocU1
hx/xPs8XvJR4Y5Xw4lCGz1xraBcFKKI79aIM4263P4FF4vdR3VV2OmLrKvGoBCZO
vUie02ZvG/dgzgH+GC+x1h4E5XbM9w1kcrypCkNwknCQzg0MnyDY9QJJUVPAEzex
H/L9omy28a/7q9iIYYIWvnsSx0O315osnu4qEBZOR+MeFAaBrWTaeBB4LEobtxX9
O2QhSvbwuUoG5qE/TKHdNzaq/V2G6WXAOXvCp5GokfzGs/nDn991GrFoaqf+3xu4
JdO5kSLPruHxA0sHqRpSeQMcZbn2wSpr6FlZoNWhplNnQVQoRcqvPVOk1btovR6G
hqA15f9+UBr3d6FkwBA8UcoeNKVWGagvvK+m7IFVcIEuxrkSiQ8YIxpSQ0sgowue
iBBKQ38TvfOMZtmLV3rdF+qxuZdD20jwxt8oaPG7cpnmi6zVpwKob7YcTLLpD+N5
1dHYwsd2S7vUjwWE/SXFEEJYtFv0l2Upa8UOU9Vfqn1QsZogWB7nfjyMxVAYR5pL
1j2vZvpCjrNDrv1vOo3VmZ+/At5b2YhUEr1Onp/BJJXGWQVjk3ee0u5l/JZbGTHd
81ntNT1THHkRD6cQK66hj+oVdqjMmyqn5/9vJIJyBJtYteVmtYJnTH1/HsW0GdDy
H0W7kLGj63ItuqqcdZlsIZ0ssH/gjSygYaRNM55mRIl5oyGOsZ+uvco2IPOVo6zP
irYL2aLuJbaIcPR0dAbyc9f5ppbCfrqd7MLmeEZWP0Exd7Ps4Ci5w0pGBJdbhlVS
kOS68peDBsYijFUMLslURALkYWT9cIHUSUivfoViVpiClDJUVW5sXR1FJgq0RTS3
RUCsityV22Tx61h+6pwQd7CZapkTQEnm6ANgi4UdruQyopU9OJOzcDyIR6sbgtsd
1OHaYQuEubzUmAJL0rluWspI/XSAIzL+PlYwfYZTsy8c+XKarqLEESqkqOLImRaj
M0Cbi72R8VigmRiYu/oP4uZLYp7uxK5awrPH3HIp1t2XqpB2KznmCuxRc4MZMvYd
l+ASIz+l3c2wfwi4vY6fJ77WbRrJUExzo1OcTLlKw+G74oqPrV06xIxcEgGY5PS0
Pz8Hkgm2W7uy1sGFPgqXSCbQcIBt86RiuXJg95D4lO5UNiPQBAEHXWyagyPQ+uBJ
CqdE478p+cQhtqM5Xt4fhM7gq6j7PlElbp0ffUR2B3TTo+kThwRaLZ1udlhg1Bsc
X0xwD6wwZezH6uEYlsIGQM4tR0plC/6VrYB8IjM5VAOpncbdOFPdWxP5SMG3pWmn
sOMtCwJ705OIpAaYLQk7GVShHtVA4OtnxtVeLGoP91WEJ4Yt4l3rjOcfdgmI/uVm
SYM90neP/ENHNgp48kInsBsG0bb7rkqWJy9GEqKoerSudhJfQbhKhdQUPbftBx0/
gZtUOXgaqzOGJ+04BH7J0At/KXJ/1EGr5bIoF7udmNh3CSk/MA/BXDqSBX+1z0PM
6Aloie7r0eMwmIcTm5Ip5Do3bh7tpqidbz9L+mJYUbVYTxcv8L1NCHpuIEZ+djJT
P/2+r9oDNGshtmlOTwz5pRYxcFuy5mrOSfqfP1j/9UmVHTJDHeB3+tsPbRkrud4j
YwFTmHnsbMjbgqLCfDVjhVvtoWSOcairjsBd9PZVF9S1JO5lEQhBsVUtJaXvaIXU
lg87WNj8btxnjHbiUApOJP1KlCQLnrZMouP6EoejTbVdr5qA8liRUWOgOLiLARxd
71N8N3UtukpV0AJm7h2s6r4C8DZxlVGqnz6MBVLYPx7pO+B2iUZAJYFrcpfkBgly
teBSMaiiTHGEOk/jHK+J8X0P/X322bM+C0s7uM/LlAlNRNBgkycp5sKihmbh2dS8
oovTXlHpHDvPFKUCqzHuMx/DOEWMWJAo9O5bne8IjL1pOJHhHmXDBD4p0uL9c4rQ
rQi4yxiFzvGSbqAC2/7NqFkVxOS1iR57Kq1s1HDiJPym6fPICMmW4V62uWf3/DQt
/YCMravY5OG+VNxTcxHIedix0NMR1sWYCs4ShwgtSE9aqqhj66/5iM2f6vPHzYTV
o8PNZrX4Sf5HWFmk9gj0DuMOX5Ma3G9tzecheZJ9Ovi/l4AHu6NyDU3LGIE/MSE9
rqbRNF/bUHAJovdtf7nZyRkB0whf+n2K8tTjbR1XlMWJJXFbr0HEM5iffNWeR+zO
zxCSAJ0SUrbtBdiO21GM8tD10CVThFEFsWsQ5NgmEm77HdRZR65yWsl2Xj59GTM8
nx45cpIQjtgLIRipg7/sqTEFfw5uSATy76rITlkqakywwbiWHCUHpnQGDnngKSHI
eP5FAlyeIoe1bEnLM5JKL2TmdjoX1wIYNDLnFwMDTgcFgY3QqNoTk4GjV6pPlIjZ
TstE8S2myAPh+z6E9VjG4GzJ5blaQKmDk1ph/tYqlZJqxldin2mdVHCaPFL8HQEl
hKeTWSrH6QZ1UQMYTvFqf4xOlw8rhkYz0oehwvLqxv0niLIQuDqvURobEqokhqO5
mxeEUkm70ctZoIC68kQWXxcvjfkejibjAuu8ra1E42Drwr1IRspUE+VXDA29UTvz
15xAmrDklyLiXkXfSsKnm9kr3wVdFgDYyCKJtFaTqT4y1g/okUfILQuY4Qq0+1UF
FUSJdY6DtVYGTB6asypPVpRAc2q8Gl/525LopqdZJ8qzPFGxHNmaeGer1EvuMWyT
E4jz9aUbnwem3gGwplhdKeSB6aoXGeRuqEJLTdBmSCPcaTjlE/mtqG65KydZYt07
mBfxOnnU4rSkbZiCTvQ+pK+9J+P4ZBSWj85BjflMHOFo5P2W89+h5/qUdXbcCtBP
r1SeCvOCLy65ka/pyzU0aLgjxanVytTdDB0kKAu9hgNJHsjYHYZTh+/h9p0/j6bf
+weSOWqsjIwhIIJS6Ns8FiLuA5SD9u52IfAqZjz1GN8rDH4l/6PcdvDgrs+e9VVZ
lq5sz0uwDR1mD4DAih1bWzxiV6uiwLrByA4VRTyXdi/Oret7uQJZ+8o3fHoXhjpG
AiUTV4S06SaSRzSBDBWyBU2EVj0UyF838FYFaJvSIskoqCr/qnnA2YbLcmdvbbMA
4iP7HLhoHKCGjid7AMoVipqRDTyzvGKbAuHbcORN549LJaIGu3TfuVTScm6tXuSX
Vr7002GzTSlNJ17wap+yUkiEyVwfql/UlIg59CudvsUii4/1Of6IZH4KbzR012nI
47y+zuJFlMB2r5IF1Dbsak2Na7YHNqOoE1YEzq/D3pi4zauFT9b1RjZChUxr8cow
tMTxn+qgz4HSQX1wZpqJVFITSow0vNY7e0mmePXI83Rta9VYH6syNcpk2JkXyA9r
Glx5y4IVkBh0uFZ4MCIRHmARI1ZZsnSkDI4Veg6TD5DMZ6eTLKUu2jjhLmX2N4+0
fe1ZaSnk+1Vh6cZXevjh/UqiiLhaExlptRf18Cw/1CD2S1WuvLmc7k+Lxydxcjd3
nU8G4F9g7vaSwYCEmzxKUe1Ek4Mu72wHbe42SOY2H96iMVmXy+vH6k7/uWeAsIPq
8G2uv7kT0FIf+2YwpNHpuxCKaOR+HYKF7L7B+Ynwka5CDd3bCCHmU2S01SEL6W8v
xr+H5oLjkT8bfFV5+IjfG8KwPKumYx6VI3gU9nimSQ+RM7hFTDX4vzMePyPJXVKY
tEUlhuqLr7daXE5GJLbMFxcNAE/46LODGoNmzti3MR8Hz/6OWNr8bHicjRaaNlmi
usCENTVZFYcUhWwa6ZPrlW0DPnN165ZjE8iGNdpSvhSDB72XEI5Iyv3STr8tA+NM
wLiRyrThdwBryrlsiaRscKV1jL/mfO7CpW/h7NhmE0khxy8v/PGwYumgUKJO/gOy
7bJe/jBwMxYDNQxxq/bo7rIvabq3RZYaeHZRy99i7xHHB3MHlWR9JxuzFzLi0QOH
pjQY55efapC6kSJYBHTw4Au1cw1ElhYMWOJLCsrXM0PlVhYTaFNrAyQX+A7/19Pq
XM8KhZhdh6zzrIpMZFD/giQMmczvM1XTCVdJ6oHg0vPndX1S5Owmxmp8mAU1JOPz
1Tf5gJkfcAqd/N2ftNQdz7aOyFSfqhSTLDRVRbiM++lxwb/yRSY3T39KI/N+iUQu
09lJDVSWV4Tltg9/o9E4qRNoHbbSzgBxTbPxpm2iwbZAtRaGwyGmTD1pBFHEh4Qg
lVSprZOwdCmHUvrN4DboMInfdZBATn1JB73D9k4WtO7iBRQYCZCvo3D8udFxcDh+
wz8/1bhjGIWccP2eOpXLBi2FKBCu02PsMFdboFFHEzHqfxC+2zNJHnrrYVnOvi5b
xdrtALJA9uhZucQEtKNksyzUBJAOe8UBpMhZyNKLQzcNEeEnZnFV2V8CPHj1hURx
ONEr9j26M1A+MYb9xRCmi9omKqKCVCjQhqN7gnYEUcwSt9U79HyfLD27e/72RPen
pO8eI597ZSBOivseLZfeIqWf/DvbIHedpddXG/RCdmJKndvw8mUSrj2qTsY7WNIG
WSWBjjJA9YMJAuPSU8oDaaoyEqlWVAFcWz1B5rSPloeWK7PE53K+gL3wBnCaDv22
tWLT9EuL1yh1x3mYEANSs1/QeyQ093ZMgijcnKBzPwgAp5FjO6Jy/3naErmTtrI+
U86jawsXcglMPJeIqBHq2igIZm8aZ1fclHkCCRRTQxsXp0Oax14BJZrbj2Z16Zdn
433TZ0NVcy2gMRSRUXQdtCcoxi9f73zPS2OyKiDzRSkYFsmbTd8+v8vcoX59r5HH
4fFfdg3zqgfOeg/nJh//SCCVBY0XiRgXtx4/HpWQg95qzniLJxC4jASKiyl6246b
vPIcn/u3Sz4y1k64XxiHBInumJmw8lEiYs+ihEdEDQ+jM/ydzzz0ACLbdoFUYbUU
gs5V0a2Q5kNl8Z7n4ovQkitDHysSc0OBN0Q5EuQaul6Sri4CE83zzfCWVZ/gx12k
oMRLVZBzhXl1F+RL2nKLWjvTwWvYWiHAfo6MLs2E2QrxuIsVvL1DRBMqyoQcWnJv
nDMnOqyi3csXBbQpBgN+FkN6vljG3L2I31QMxCDVtXKhmLgkYGMtqP/VZ+3wsVT5
eo5ED117X2VPIzyNRR+mhanSjyihKAsIkVLpKWbqVONzI535HzYWns135qOm5fbd
hjNarz+Jn4WI7SYwE2J5dIKAnvU9gJQKPQcJPK+ich5u+K32UOt6AQ9aPo/YNo3J
eDUXSvoQsJzASkaCTuHGvminhUUaOhnV7BcghKCbbutjRSrVkGgUzmv9yTtT/akm
4e+A+ObhMnKrtSlFWHq55OLhXYdAUzXTkq5i6/v/l5FgqLeQJTInrWSjdGXae/WX
PhUaBcD8pST+MxRMVPGsnDpChwKuv420fTjh07V5QjYoAdv12pSuhqNCETT7CB5r
RQ8gs2YvygRjdPOOR+ddLuU8z/EHzoAA9bpoPaMKrKGxxQH1FzdlBD3DBvNtKFlo
UsKhHFOaIn2Zsx5QxKc4o+4yhDmj0FH1RaEUTgj234DZS1ZI/C+XcnVlF3Bmy4Um
Y7WkS1ihGr0lPquEvKcRm47QrUGh+maXV5rIM4i6sqn++G8Ew/Ss0ub0/YatAyVV
o1wO3eWo/WXOarvdrY38Gbnxs5zN+f3iPV8gjhuXAv9/cAVlJwNxVy0Y4OXn1C2R
YD9XedwmuM6cL9pXo64Wg+DzanBXoobhZpAwgI4eZBROsQ7TP9VL8v9x1ZbOKily
yn4hZInqXYxBgqLEdrZv771yzjH6RT4rS14OR78MgTvpGZi0ja9AXzqhsrRmb2i8
J8UPmn4eVmJ+aW5CNyWxf7RbdXrCbYKhoOEWkCe6iHkHSh9EFnUwib+5Vnsi8lG/
AzTaS0RzoW0cCXwp4W+ZiJniLh2pjAnZPKd23Ao6yFDYbjeFw2SwKTlRrwYNvBhX
/Y6Acv04HCsL2jr91rnIdqwHm4LfNE81t1VSrKtynYOh99RjsblNYlVL8ghEgE4f
Dzi2e0Cs4ipaWUxLC1BO1u+DnLYaGr/evyxfKXuxG/n2RzgOv4857vuiJeZ0m9/C
YqwQ+vkfoNGYjwocND+uVMGVOomuH0jApa8+Qj3WQSuKIBovpkSBNCbQdso5HWhG
Xn97c7X+d4miqoqYyhLBe96oDt93hQ5vuTyyQVayhYhRcXVWdjV2Birb3oDWa4V2
KBChEFcxgXZySUpV8WxuqjOuPQqDCbb1dsPvKE6ihAr5qgzGNkSaxkkWjzw4ljbz
VHhYtc8mrgZCJnla0nOR8d2W6hQreDZEbtEhDItBMl2zbQ3a8KC9R9367rmhMtv/
F06kUZiJTYjPnd0S3iXzT4abn5vpGRFSvDG6VDux2uFvHGJZwrpBghtk92xYDywG
V8aywkoqUxyBJlKNFNngdXk0x3GrfQzTKJGT7EE410jUuenWaRvB5Aoe9gGqhSxe
f5wPXN/mcWrN9KaZl+o30A==
`protect END_PROTECTED
