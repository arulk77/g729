`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
wX0M7bP4AH9bR2CpyH6o6ABXxp6V/BTrDrrJDIoOUUNtS1KlaVFkVLi7GyvqDp81
0/fANrl4adWj2/xGgou6ucylEXYfMPWD67N/GWL7dpORrJi/rK35ZN2eJHnhj5eg
1+L4oUEIPxfxDdn5oxtpi+GKUZV99mvFpuxnQ++p88kipQNYYghjyZx4rKbzNSig
OTYq4TLwCRaDg2m/WnTtRuV4GOjSv70qIqzZ+G7QJzo=
`protect END_PROTECTED
