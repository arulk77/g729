`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCWbPX53GN//26xZpXrOjrV++22+tywMnytxOZgtQYdJ
Lhc/UkyORv0t+klmt5RsN2WKTj0+QRC/5ty4CSUckVelITsjkUXaMzLqfXvhT7Qb
H5xnXzstXM7bBKQRo12oGCI4Qeq3An1C+0wta4iC+8EoWtzM6yG3mdYqs/fD6pM9
wif9hFHm4Tpa0a8Lzpt0ISzPlmkv4eKBCyyDenHzt5LWDcS0aqrURwhlQeL4AFND
79oppnrJKHBH6Eol8AasjmhMOk+J06o8pb5hxhX8ocfadGNnJHe4M9yofcNwm5/s
2KgQsbFX+78Ouabww/PDHL58M08Qyz+8SjdwLRAsRmmUK5SvAp7ZRAWu6CS/Ps+K
iUndqPNVwcPb0EW+/7sZZPQvnEdM2o99s28a7slcNSuaj/X5Zy/Kik3IZXTxrGlC
`protect END_PROTECTED
