`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xsDyVH6c1jfNEBGvg2kY0oa8EIZIAmLR+eXZWTPKS1M
o5wQGbrEeDXZw9gSaqbXHItqsPPn5XBSvIFOuLTVfp2h1kYLb4Tfz2ZZwhsquRCn
S7st+bOXVJag+FMKcllut4boIASBSEQRsFYJsgl5a4aHuAQUumdiDhbm9Racc4W7
Izdmm7VV7QJ3BKbUN20sHyhTAOuTNeS8BoBEtrIkBg3qZpcJGTG3nCQJzUbkSP2B
gFZLTFKTpXRTuVQmZCV43IHSmTbJxX5f4s3j7JSxfXKiN99LXJ/DdQ+6uJ9qTz6x
4yLFChvoZdksxa2F4R1S0MVmcs+/QqmEJFMO15IAEAlWL0iYEyspU9X+mlxxOEZQ
PMENZaYPVVud0WUVJUUACQ==
`protect END_PROTECTED
