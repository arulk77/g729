`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
whfZdEhQhIVICrvn0VMg7s242bG1rLB3tJ7XYGIS0ye5zQUgmHeyyaq2TYShdprY
IIYursOHQhovGdFKrJ472IxHCj5ngOCdX9GQ/5oJ5XTcvCI3NoGkO8/KSVOv4s2I
1LOWxcz22ZYAY9Nl+ZK4embYE6zGD/z1VBrKzj27/+6D2VJq1+zLwKu/EjDFooYk
mbkBsV+gnpjNvNOnbeIAPCvOKhj6JdNiGP1mX/Lvh2aUovnCICMRYS/UuU87f/1O
aXUToPzolLI4GrYDzpu6SSwrap92FH590vThDeqaghwpzUeKfBcRDG7BKOFFYaXp
N+siCgCUWyhl0+zHQ8HKyc45gPmyql3RINbPpA4CskBWD+pjsSa5bZn3R3cGpNFD
`protect END_PROTECTED
