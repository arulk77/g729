`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49gBFo81A6HjBC5kxR2enk8vDMFMFRXtjWJcb5isH2ua
lgRzcIBKtl8JdRL9XDQaqD4jspfdSkl3QJF/yduwCMOaj7UxnAESiocoBpfgKqRj
Mj6YwMGyz0CcSZkw+BGLqW+m3At1yBiZQhv4JP2bAOtp3K9Ne8MXIknEPEm8Rp60
D9JzatM7xwRcPbsMKN+PMD0aHJKm3lJa4+rTb6KaCUHyN0vrIOVf1y5w5hLhl5uB
j36oXfrUtMrlVn/BWtS2d6PCt0iXX3XoinJ9yLaPoq6SsmsGZskuJQH6DQ11iPFc
yB6j5OheZ1Om7m/fXE+mlSdlEaS7ZiOHeHEHJetuyjQNE3gTj27rU3yuB1b3BBQl
Sg8RlrIDJYyIPrEmTtjykDAl/AFzoKyqIcwlutglpVa7HQmByU4tuoy3Bd9XL5/C
OkFCy7E8DCUsiNLwR5nAHvICdNmqqU/i+NHF18yu/Tq0MgE0Sfe9ZCJeSCPpKVrE
/mYAbFuQToYjANwNQFxuyPFb6C9iRrWwLFu25+XSWOZCJedrNJgtm8IXLzO2hdJy
MfCmAmfzjNQlEZympJ6hNmIZ5UJdUca97mitTbzIPIA0oWAFJLjBiYGqIE33mH9s
Co4CijyirCPEeG47FSfoha84s3/ofyzzOWWN+UGbJiN1ZmUoeLNpH9eybcHJHllm
aDd07wDLeIKeen3ZkS0xjhZL1f/sUOjLUCheVf0cMBJAjERvk9wJRwv2Nla0b/B5
su6q66iaBJudNHQYET9PBumLuwRjt4LG3ZsC4UMAW5SqNbeK50Q2+mGJ9mnBKUk1
B+ymL8FgHZ2YcIP7Y2cADZJ/f11QOREQM146ViWOOySZ8lxEAyCISsiy5WAomJpo
gqCQmFeygUTWSnvv6nl/Vbid8SoBehomMnx746bbReq1svnNdgB69JQchCiAKrC1
a4Zn4oLAfCGGndds9NCgGg4VOARNWCDuR/pdVvgLYSJe6YsFnAgvodcxH1M+URAZ
akqrTuG4wuqUzGcKG8jAwzBCbI6WpknlMqzK7suqvKLLVZlUrOIMdpl9gP3OPfmO
E0Hi0jM+Kjfttb9Pr+U4GSbHeg3xNPFnuCn8dHjrNZ81hgOqQlYFYZQxGzJfBbNe
H/QqqXlJzzPOapHAD3ev7YTAYcJnWFOAopRhvPnCUuKk/gg7wY8Fc4TLiLnQS3y9
JtgTeAvZH2Ux9qiC0vY4EO2b5RHgz+oRmQNiro7L9r9I+qLiA0D1L9xHKzNJBVPm
PqXGCUjb/HAQaOicAOom5x5UsVZgeS/w/oUAfQklaBtQoDXxKQ86kMWA17jvqPzo
xZQMWjLilBM2S4+caDnCvM/aN8prsZ1rgwiU9BARhNMiL9SDAm3gTJLoZxGVo9EU
2RNMeJFf4kXlXfaZH2QYA4sc45jZIyFPW79JNFJLjfgy7UbAvGD6rKK15A8WIroG
2lDM7BEBU4p+9qG/vYxRNim53LHse3sfGAZC9I3FSa8fIiT5UGcxfABnra2YndwC
m7pYNdznzS9eGjHCVaQ9MSgo2u1bDob0eaHKX0nR9QnwrZqH1njtDz1o46QSGXoS
hNdRIW9LY4fVAVUygR6vKGungYIMWCss7/kG+q2VHYTo+D2aZCo8dtJHR598lejs
ILpvIeqd/5doMF6ZSxNUo2H1KkKuZ5W7DfBRS310hUelqKR1BqHdaUkVFNwB9Cjg
zUXlfuC8jfsm1+39GWQBGFaiNHXfvb3fbU+t7ei+Gm4THDamGvk9Ruo4iogXE5VI
QXzw3dOrk+MZR6vhvm18eJ23SZTUe9B1aOmcTdVEv8RwP9/KT/oYG/zx7EyPT91p
wqIXM/Je/yslYGIRKaJARggkBf6CjbbwiLzIh7a6GfiefoXcOLimIJ0ylE0VXfw5
udYgkda/ubjJ/bfAwtD8Ztqsk9GKVIc9lbHt03xJZoWsv5C5apN2eh9uf1jvRAcl
qgonaogUWK3FjW3yWoVKKFo/YK2vtThdShyCnwT2znblGHoOJpQMh4Je4mzamgdC
mz0AgCKLXwpl5FY0L1jAfbQOh5w1Vn2jZhhEO7DSy9yxkGlo6BSteOVxoXHAw2Y/
hH4+vJWKuUznWUgu5lsmIJaUr/UKpwfxCE7FymyxIcfW5Th0jLHtVHnRLXjpQ0NR
TUunnylVELF8IQy1Df9xmm9vgoZcmwNBO1YSXStPRyg0+6VKTLN6sL2YM0KOQJaC
S/6vW2roqq1en45e26CzewMhZgvNV++cM4nlJUQ11BjP1VDe0MJCRc6Vdyh60bxx
bBHMRMQ96sxMrNP7uT+UrltI1jFYIeVZvuyl0CjsMK3SgDHA69aGvUc6t/VUXvnN
GbzqidZx79IWGy70dhb8D1YNjXbCGIwLNiGMl1HasaIyxEfHHbh6ZNSPuSZo48tP
cOMfHv9x4Idg8+MosqzPxu++hhye+jOa9ns5Tfxn6991zxgCV0SeuOZu3bKAzhvE
zgdNlka0AUKltLZn3dJxh1EtOTeEALgS0KFmRT13TRfMSFK3Dfj8GGEHF/dNNoTG
mD+BQPzFtbowDud+2BnLThSKXJpY1knobegSmu9h0uvPty4b8GU0Kat019r7gh92
4EtD02+8gE8M1S4X2+kP60OglSWfQlDxfUbb85Z//eqzzr7Mq0+yMDQqI/s02rBV
iRA9TMY1X5y5yb7BgSLEptc8OCNFZSZvn/BJ8VBMR69gmcUdYeWgzNuitt6wnKjE
3/DwWFY2KAGE8jUxi0QJKOEmez9kSoPt85E/tLqnSkLxigzxsVv01JRsQ/qephRX
6avA5Zgj2hBZkImQBNdcrok26bejUas+Ljj39g47t03v5S8HNvt8Apv4IyCkFkCf
tyTYFJiZqwC5wu4l9Xi3DMiGmL4qAFXgdOJgfRrrnGnFs4ldR4EfaoiHbQVsIAm+
rzjg3k2+JfYfM8Zkyc65sKCYGKoVc2ynR0X/gtEFu+PBmX92a0XNIQN6D0cDM1ic
6Ul/6xZo3A8oKEvrfR5DLD4NpKBxFwKCpS9iwKRag35APHuxE/oNZjsidHup6W6i
qoF3G61WR++LucF3PCK2iehXITZ/N7wVXMyOkw8MYzFeaKy8hssdMYWrVR3mWhaY
0XMukweJ6Y0YzLYE1Ss1dveHqBhYKRO5y0+Dzje1mCByzYKLdaLT/PIiPiJq+kR+
YCd9gZfDajDV/ZWNQAiXWmQ06X2/LyurufpWGZEA8qqoncNUnsQsuvczL7iwT5SB
3K4vF2Gs3Y7Mo4yB38l0zs4I/CDrgPnMWAM3IsKouUgChHBaiz80qbFK7KM8vDcv
z9bylqmFnqmwnwlluZovu8jR6xcB/jl1jsFIhM6YrHfytI4POUJH5UB244U/AaTX
hSTz/7s3SKPNMPEHnqk+B0XYTejKl/vW+EY7VapJmWg6IQFgCsezH1rWmyga7Yj8
SjdECBh+jvSH8/KbMmNQjtiF8qHg3I/nFGdADnBBWZkI1IrkpJv/zXoPQ+oZgsq0
t7nOBQVjkycdp70DXCvKZrd6GBetIVaMXGlKjtQA/VAmyz8LzxyuuWJCPPngW7ZY
VLbBfyzpMaOmxfKzH4ogBVUMuIZa8sUezUpMS84NcuswzNF/MXXSUSXNYKGEpZd3
h+uH+IQSNPkjt2erI32NH8abVq2ORrABpD3spiVkOPuj229S3jHTSzj5Z7DYLUKQ
HnDY3QRxfCV3khDG3KIP511cNeyvDw2WsB52ekt8IV4AFBuZ1r9iiggIaGpKsvC9
bbfNoGzP8WC54NlfR/6Fatdqqupj69woVJvIfkwR7M1rfKVJQmBES772OJ9hdrHx
SamfIXGBu1CsKF1R/8sAQ29mAK6MA6PeT3mmqBfQekRhFjorlRRUp+Y8BSLWluF8
lwwWukY1qmuw5kj+Y9vRuWyf04hUExuwNJ+B2nbYesstr5GTmSwaAVh18+tCV/OC
Mz+fwd2vn2dqrH/g8MPAuCK+z9ez9gvY0U0xrs2adMIbFfvR7rKq7lDvm6wJslox
uld3FYcIwRkJaff00DJlwDund+Cd1bqNUPhMN00Hg41k0zshHD8OrPKtuhjgvFKO
rcWcL+8Vl1PyMOITKjXXkY3A7P+CSpSsiweiH82PAKka4clMopZKZEc1epzJSkuq
gcA0OlXEW2JscZ7ngjEGIkbQZkxuXoehfYm4xtIipDSdStE7Mv7og7azKo6TQkmw
U2M8uyC3yG7r+p8cbIEf3lySaf6SBh2cqgo79UAfvh+cYWlbDABy+ZeUTHPN68Nt
+wvLdTPk2HTL34gglUEtToHJz269O/Tp5F3rqI7MZMqccWhpOwA82j7rarkYmJFh
4jUDfmWpNS7BJc+HY1Yx2HkLrZ4eNheJLva7ONpmTQ25JdFVEu0ozcloATNAginD
SpxUmHY/l/jsjlSgYGGnsL09BJ49BuQJodM1XsfZanfQRIK1zHG1R716n/4dxs2N
m13IGqWvucjIMH/nfeoEuOgi4uugvg93mds/FLCTrsQZKiQr1Qvkc6VdHNJWPb5H
qwNBR7ln6G7kVtfvRN+3mFrQEjMAqNTguex4ubu6uEpHWmsBPZZI2qnN9jnVgJfe
lf5OYpysdPyyyrid9CmzbOORBgJA3U9kkv+VtNNbbZOkcPKbSP6LSiB3DYWXXtME
6z9pPPKXGVXdBHfYR8WZdm6gRnprqdrZxpAqsKJ7H/uQd/yzAEF1XurENX5Ux54Q
uP/NT+fqlI9t4ESma7EOqgvrjTxLic1Tu+5PldsCF3Amt6NC1t2PWwe2LeNj+Rni
rw5m3HgTtcGCStP8ugmt/Lqy3cbLXcAgHBmVt+153EPsWgLJdeGUMK8B94auonwF
l1MjvGz7wJOQSM/iqYRXYdLj7VBnh+Rw8t1mdRL2yzwm914uNXPIhELjEWAF3O0N
h8D961td3x2wrvYItYemqy6VZtyLLtePnGh0/3SHIMXAuLcYbbqy36uBCGE1qD2R
OiUT4EQeuPTQSm7Mv7rLtIZ07+V+k97mbK3CI8407g+hAdLos/osspovomzKj0zw
T4clIoBrIiQsaKjAVE6Is5aYpn+JSjgtemZZyopYKC8PifTWC0KVhXVlhwLXbf2X
024/oGWSBfVGGWLFOtlkvxW4fgzmMVCk4p77rqGRybjKLpF4liVYZOic53+HUqgS
GBcokPeFkJmyhuyqpd0tKuOypKv9xdqMyt1YA1vpXuI5hM0YqtR/qSrFj+7B723r
xsbniocF0IVgFhoHYpApGOnAKvyhID9U+8sKAEJYdeCdsgWybmemJPq4wJhQa+nj
ra2CH7O1XtujmArv3WX8b7vKc6i6JtNBxsLig6LmtDCKFqln2XsQ7dXB3dYkmlxv
4qm3jRn6Sef16waNhiPfP33G+kmkmDHkVPEJ21FlLRlgOWkdxNJD01iQpklFvJF1
YoC7D0o5odjBZQt5WOLB5Pi0FrH1G1w42QIgPTYPkXxH9gDipeUnS9SqN7SGEGLt
OtnTdHglq7AJElR5TtNWpToyH6a2uVqfVyW4utuDYfHPfXyUrbdKrIWEPUIQZ7EZ
zromPCP2EHETLmgV1K3n/tOveiHr2jtlWG5Clk/hcRJ+J7EYX9awFKeO0a4Tf7l0
6SYmPH2Okfr178QiK+9ahZyw28u7in55as77Tl8ZketUayDDxLNK1wiQ7MeXnarS
Dq1w5VRXeGFMKP8SYQS3GRjSRCrSFe+sdUiBt6xBe/Arf7rDuJRdGxMDyXXshpaY
PU8GuSipwGGljDl113WZl1vAw5hY/ChrKWJGDTuO83V1IJ5rXc5nwve7vzVT22iZ
Qmi4o5kZH1pqui1lX2dRkTyRrJqWGz+JCUgQfnE80FMXM8L1nmHdlCVMbreITqzH
Zzu6nuF33P8PPtLiaaYrFwfCWq4GfPFTehY1R8Hg0hiCgwUWxQIbZPlYt3WvNDdB
iDJC9gyp+Vgh70DMQvFnnlJfiG6IVXBM5kg1/j4sEvx5qsZh0GRdRb2pBHCHFyZB
Gd0ZMQRj/YxW03x8SbTNhP3KFZczWiTdq0lbo7/hmJM9hM7pvBMIDhUFBhsyYxe8
7ZiOyQup/u2rbBWhPQAYbRxPd2Yvdqil2EJgWMBTR/SsmTONMwBqkk1eTAykNFlZ
s/tw/T1P+aFZdPz19COvgjaM8H0mGkVNgqqef01EslCs24iZJIzm7phgOd977QUZ
NP5PTefl9uR+SzbT4ywkD9SBpyKKbvWcxHL/iv0e9/URNa20db8vdHb9+/qtioLI
u2aOYJB8gY7FpvyT/rz3z0NpP0i2g6uBjpNXB74hqRgES+kMDiSnX3nu+ukBDFaP
6fZBVarCb5eWTylVNF1GgMuTsgmRd8daAJzmo0dbwM2/GMpsHE2VS8mT3QClOxfY
J8Tv6NALzPJnE9tL4rD75UDuXIz2JGwbGlqThNaJnXIFRuThSuBFPFyR+J4YwmWc
OieSw/ukkN+DTZ17mCnQCwPgJc9r7OYCZ25uScb8t9xDe+F2wiGqpGEZzw1qruBx
mCkVUhUq0xzuVnimiwEjKVMTGWZQXZGhfDZUkLdByVwGKb9S4zEoXNAQlbPvlz6t
HUH9YO3JPhaQg9/iGxQlkKeL8vFANs5a7f2azInKKn5TTONXYeSmtQNO4lPn6Gzp
/U/g78Mbz02i33jLrJyHVfoBwYEYWMvyYzeBQ9g5P7me851LjAJxufODRGmoxFns
lxwwxkIor1nTdqDjJwiSJmLMd6LAMqfDh4KeTflPc8T5VKrEgK5HvUH8BS0BIwBu
avrLxF/eEiej1kzwPWbwLQ4nL2H5v85ZF/v8JdneAoBk/c+ZNrX2pCPTigobugGG
UkVMZsTNxGcJtyK9+XP9rvbzvAnwwwOIj47ffJqvBfXcreNPy4MtyOS/7y2Yb0eU
jTionYrpWxr5lD/3PBTXPUMrE8CF7kPDqNCoBLYOhQ+vsvLLqC0q2GkYa3/H8PiF
gNUYLBREOk5q609k9ff1IqjV7f+z9zmH5a2moq4OWhHhygfDH4C9Jgo3Wx5Fkexm
h1VZCUQjgpSHOB8GFylZ7kEF+h5wtsFH8/oueZdcMJRi3mizfmr0MUhwrYKn3kC1
wmvePpdnhrQtvDsgzWlyqPZoB02vlsjvBWTYgKa9pa1u/TupMDwSnSvModz0z+ui
9JtIPSv+nkmeK8TsqvRT5ZM26loiC4IUojiH4sT9gYUBMLngGaViURH1VSmyRuYF
5MP0GQJC06BDlKTOeJxV2bnNsrZpYO+aOoCCnIg+NHmUEoEK9sWmGPJJ8V/F2KQQ
4cVJVKz0orz/AxMKk1urFMCQ2bO2EcMAk1bFCBq8kmIbByqVyYeIZnTcppux6311
vpHxzwyZc57suxRoOJ8BbPMwpBg55wyaFAvt3OP1VqCwym/9Bfz4+KIOSpXrOSQT
XNqX+gjVf5PF90hb5KZwJWsl4MHOLGpHcyDCWFnEnGquPrhO/123FKZwvRDQi3Z5
fiARNCxgCbaQtMKehezuLfAAeiaQr+bFI5jFYXCPub4HcJ769CKHl/AH/lujLQnJ
EQf58pHSP1WiAYX7ub57e6frjCY1K3wYwrO9yFxSDJshQmUIUxahwOIOtfmPZqSc
YUJClyE5wh5n/rQbIbahiahBTK+t5hG9LqOyTCBfPrxp4koXaXIboqFtxK2D+taV
AIMTe/LRZRDfxq5zMLlBgyI69hH5iGH9Kt3+a5u02EDsjUgrpACJ/BIVuED2KHSl
HUve7T37ez3yUuXnPLVFny9zc+R3RMqgZam49Wvzyc48wn6GYp6rOIOc3df1GxlB
AVa5ZGI6X/MGrFUIbkygYiQMzCEESdyFzCfIJPBVbJzWRJ4LuOqAFJvyBC+8+4JE
36Fp36jPNCYQM9y+TLjcRv7IEgI1CosXjU/W3hOxlnTYGE4Nam1591Yqex7+vegZ
Woy+Mx3mP0ekdS35XSAWAUK5tA9Vje81xEeeusrPoRPx5DRsRHIIJhPP9H9vG5X7
azGRFjAzg9WmJZ45h8kt7tJ7NfCpixQ83mV1NtaJGk/X0j1SSDgwR4mTzQ4grIS9
blGkdQI04e5RUsCA0zDR3dXvkNwBpI1YqdMke11abTc2NwN/iA7x0VmQmbXm3qUA
VpC+YGE013jRzA6cbt6+DBZc9oYISrklofw9wCZLLmk=
`protect END_PROTECTED
