`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2EBoZu9tBf8wFLCnm6xiM/75x2RF86ClEnn6A528RFw+5tj8Wcr3IYpKtUtFilBc
6113ki1OowL27C3AsCD/9B2w8g3i51GQBvlSl0NVop7GfX0irMSmxKD1ervF+mOh
8TJ8u6V1sjX139zH3SxzJ0pmqQMpIEmpPZn/VpnXjxpp/FkCr/p1pOql+RYzuXfp
yLaTRBxGBzCuOsSCa9lIODYiwbtbU0WMRr8sa6ljB+V1mNhNm8SQ1qz1ZJLN2DSr
`protect END_PROTECTED
