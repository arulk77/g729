`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCUviSIkHb0mqToVUXjSC0HxVEwKDN9i//7S2IogC9DO
w8yYgQuBYcfdfwzY5QWkB7qcs5UxOYt69616x3psuvUFM6fFReik8ZcDsZMJK4VW
1O6QYJXerZCyt0TMFQxRcGSjqexUtpKbAr9sje902pA6j12l9gml68lTFyPOn0MK
b5EnUJxklHXzf6elWSC2+TO2vpJGrUA7w5gsyiWV8x+Ce+PVwRMyoOLvuHCIivYX
E/OFwVAhONQELTrkK75Xcm3YMX0N0zD3yrkHKR822xsAsrQdpSiUL5Wsq5lC20rm
ouOf7mqvnUP8t/Yt+bptzQ9LMAhhGMxIVU0DcwZokevdN5KeqCiSIgonyKCW27Hr
zuF63T6BIGW9M4UwvmTZIQb+5hqlxnvfOvwMgCCQMW6urwrm7KPlU8yJbXYBgokJ
s1blyliFRfsdn49XczBDVIE9K1JN1BItEifOh5LtGdBaICBtTlT1nI5teLH+ib9s
TSjBgnBBTxl4KHuKMTnVscmx5QMDAVbjkH3dzw8b7lptDGbNXnuuC5Yz7+0o8hDv
dpzlqO/MsvjYc0CLnqzsXQp+GtQ6QcJraonHP+eFiU/PS0AezK84uIrFzkZ711ci
W1LiyY6r/lvj5atyjOSv/k+xenvpArfwEiO7AOkllTXK13m1T9XAFPX+7d0VqOPI
4HflfPnOWHnE2xm2knxmXcELk/lG8+Fm94BGdfFANRabaB38Rcta4+bFBvVN9MiF
NKNE7J5BWaf526S4mUwQjylRB/osKJitBwTB+ej0KSdq9MYe/84GYr8b7A7f7qiF
dDL/OeLF63dPfQj+UHHa7Lo/oPMl2jybj6qxj/wBWZM0EUfLv30NkKxquDyuG4TG
OK05DwiUACX9ABJajT2wHpwAnqYJJY/17P6ztUxbU01weJNPSlq0DAv6Rkujg0ZI
`protect END_PROTECTED
