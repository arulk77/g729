`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN8adBSE8DZ1RzmW7Pgklj7Aa4HlsXdxPDz5AALhYadYk
s6cGpIvkWH/+VOWvhAXJbHO9350JCj4WUqq/qViXzxv5mUp9iAqDZOULuy/+gEsq
g0ifZal4DjSb8wnJTwbN11y6PPYE59L0r948A4qCX+aOX1ARGsYT9gE35bdXvbO3
gEKrxwEZTEZB8UdNfZ4Q/n5LVB+a7LtD1cxec7zJ/P0exvnMraWyJMIzJipeLhzZ
QUF9nT/yBNwUDDFUh5jFcNWwan1gOR7Gq/emkEgGmVpX8DtdL7CyqbCLyMebqeyn
riFJPktczEQcXmjkDOGZX8awgDLBmonXd9QAzRFDzzaSXnb/iRiEc2D14S5XR5Rc
b/kQHMliybbzWH+eIitetfV1tuCuztvmft5345oyz3wmDgXuqCCT5DQQvOBALtZQ
UQqsavY3xCXRRKeDWEFVpntY/iSRFbQlVo5NK6ED9t3QLKV0xGenCwWFmaQysQzW
ShPAUJQbh70Zl1We67x3F8EMau8+dB5KGKXDjFUW3Vb2P/l4u8/Ef8lGlqqksVDY
64iQqX7oG7ws1mnokwzQ2tyoO5Aga+CyAHaR00VPVYy0n/ru2ZeTTnk/I0k6Ui1x
XCF5sNSDfaJ99DBDUJj0/OX1ZOzS8wGRcYOwHSnb01tw619RSOmGTrNzvX8ysB1z
88xOES2dYyJAvF63F7wz6XFjdpl1GB4ESAt/Wzpj8Qd6ZKiPrvGb11HdHuPQNwns
ZpQStKulpEWnj1FyJgQjgpKjdnC9C+AHSi+VBzPKnIuPW8tPupSIIc7XsyNJk+UP
NgFN+X3sJkxWXNkWBMmMahTuZEl8Lzh6CYXQ22xWlUKecmicFg3Zw/K35K11Zo0Q
hQ3DjAQLup3PF8CbLnuHRuZc2CaRTNNjJ/qGi3deeeusbgyEPgyDU5nRym0mI7RL
AKnAu/pfpRlWtyxL7gUtavTqwbybDSEheo7msly0c/ZuMue6XriiupeKAificwoQ
2iu7MEkT5A7AqJ9GKFP6kQMvDfIoKKPqO1ISWJA4NP8diWh8DhYDimyKOriNM913
hnb/TLK1DHrsC4elHU04pbcpJfERLljXAqOJmlLwNcf4bTUwrsr5t9yA1TW06dKe
gcKiLe/OxFFgT7WGA+6nIhnfESeZ8wUuzRDzVLsNzH6/PQpcgcwvtk7SjocMfx+N
Js0Wq52ElZIBz8MyVH9RMhedNknJJ2yNk8vj/J6jPisEZje2MbWURioqj95uq+YD
J852HoQyZE5+KoFAR3VOD5hKoBJIY36Qh0I/CJRVO/cjIO2pD7lDJB8SZRVQr7y2
UeXoOnG58H0Qr3VIG1F8/IUqsw7cI85M9rPFBwFTyFT1L+z3kAqeTZZh4VAkJbN2
qCJjft+H+p94N273XvR8FH8Qa88Ku87/IHTrN+g/6lvG1h926IwlLExd6NdIpaJJ
lJTWZ7g4jHCM2p6Iml0P7i+mnAg0ZICnPKVxnHWbuf4poeC0R9XZ8NyW0p0W6ozK
CuzpUavjQ27aw2QOTtUM/mcaikdhBRT2UJNZ9ZDrrXKEdgx11i1n1Aj0WMCAQMPK
3c2ubgEwDdUrspn8o6VrrJ0Ssn2ZXK58KhxQsuMzfyQlRo9qjWQ8n+7FoMM/O06G
5+f4W0tc/iLx8YY2KHk5zrs8Gv+KPYIxyzfpnXXQH23JCF5QwjH5WRNF2qs3kGRT
nbqMgsA/nH2YuKfjsAnH2t8lSl/6dq2QljPChOvbUJCFxs8shQdXRGHgMiZIOU8X
vLOJh0aThyYxoJl1BuDmMcfAXGE4Pv4917Sd5p7REc4C5VZWDJdK1ZHNLstlGSiS
J3WnGKOiZQWJEvuV7x34rRQqBfrFzbfvI0bQctAh9tbne9xu78XgAs7xCvhfUEmp
WbqeDT5k5BgaDNoycFHAtfSbmYjOPlZgT5pj6XEcq5RomebqVgAiaIXAKAz4Befd
tpQCouAcfXRXPwkNzULV0UGZkkHhGQW1TjKqZLOSJnzn/gGodN6RUXQjpZochoJC
GcKPbgVZPWQL0tTHP1Vk862zqfswqtnUR79Im5Nd9WxKED3FoZ9EfWyBU83I3wWU
S9RedOHpRr/iOFDhx8KxnoEKmdDg1rZfStTpZybB8ymWTTBO9FFhK+smyb60aeeG
PXckIwfcPSdBpPpDesYEiIzklwnk/PclDm/ZyRYYP+ROsMfM9QvCD2Uib7njIhoD
enB+mQtq8R2bz55Css8HPTzTjG8m3kgYp7XBVm67R38UWcDi6sQcPU34HmqPHBKr
kY/bwlrGDLrzwxISOvBsJY0iC3Znk8cpK9i1quh6KWLHqLDBkH+XxtAuc17Vqnjj
COpwlNWVPEtck6vILjimXgO0LJaMA0oEscQcoLUTocDorLLAHHkJC1GXaAxGy39P
3zZMq6GtfG49jNLT5PWuh3/LZiRW8GeMU1k+gh7DqS+gAdKO2GALnIQ/LaCK15Ue
vv1VSSnF/S8bD/ud8oHmJ+tQurSV75fdJktii+HxGWfQ7HvDz+ODQXeJdZEQJ77b
32f3E/KRlaVjZNCCy2wLNSMF11bM2KGW+ZUnxgtkEo4Jt9Od460NXKpwDZR/osg0
Q4uItlQeCnHJmML1MX5z0oY+5Uin2Cj4ZO8HlttOQjK5UTilPtOdlfADh/+Jk0Kq
kGC4aF66YnlzdoRagdGU54wfIChif4AZRrwlIWrHaD4xpm4RUOlOkLsDIaDBEQf8
76lAHA9EfKsWUwdhOxCQsNQB3dlegljHwfU4zGAqT/yPMqaEmC8+qnxCnwrsUF5Q
/QsH6P0oUU/bpbutITlbwJCdMlLdpRQ8jbUpyf/5Z6L4fiOQuoXFejB+ExYDwQrQ
+m+wa0MIn8NfFJD9DgoRa6N1KU1+1+2LAGNcbGD1ZCDg76l5ZMmEX1MZ4NJu8l9v
zqU+BUq+Up22FKQyhijvbIRUHYT/HUXs4lfaknjzmKZnyS0XBhkJLA1eDzBKz1VS
N2b47UzwfRadEdpWgDOiL9dBqhvqFSjQLlnhRYWSdGFI9tBLj8ziHk3K0Hn+rYW/
e0yExOyDfk22qVlLhRsXG3Pg8BUHbdnc8KYPnWH1BeNZQ7HnSp54RPM413sTGtop
im24Hsl8olLPy/Ka3WVjZPzhGNgACsPHzlvB0VnSQ/ZJsg/AEmp2vEal+pYdXu/r
5ilLWje1hlMqSxkHp6CShqfFqepv7vWYEmT/G5fARx8n22SIg0cTf+iz7e34zHBO
DBMPFvUj5wiMVQzSeSLWU5Cn6A2LYOnBPut0Wn7SFIWKu2mIV2eiB3oDkr9GnotS
R/tOVyb29AEdTfH30Dh8wmCucm7HSbWsJQ8lWJVIiKEJW9sEjOAODi8ptenrpRSB
XMXqkmJASOJihAnEAo+LpVMpBl+RIr889nK9sGq+1HUe6q3y5dLEZOdG6dndqqov
FCK8nxxbZdHHV4EV4ofNWNDquPMm1cwPOcW19CXjz2Fjmvdwr6GV/+2C7y7/0Y/q
LOcFtxZQK6A+XLv4DCb904ixf7G4GaSWQfKx/GioBqsxWgVobuTflXdiLNfMSkak
ZFVMWlaS0ldIiuxl8qcmR9+rGcChvjU7kIkv3HhSz/1aoHp8wv0R2OBz0qmAeI/e
LEKV7N5qt4uNozRYGKBHMLOzPeJdUTvGyhVR3iGjWmt68Og+UQGI6RP04MA9VBxg
XwSGG8CPaQGbzfe4H92rt5RrDqLrZvgE6HW9fQWAmueERHft16AfnE+mNSg7pGBg
e0Z0kyymBt/xpKcCrPTnPiu2OSN9TgNyHTK5Te9O6To9/J0Z/NODVpqbRCsJIsAV
lVjX+NbulAABWYp22agtf0soWVwTkkv4Mqy4vpAKPKAREb04ShSg8wImPg18peBq
1c0WqPnIlM3X5WIGEzfo1mKyHSmldWUqBQnRFEjHJgPSgnA68/FOwZJG3VRE4JsN
cjBrxt9J6OWysn1QyStWrpcyqlZJ5B85sK0nXQbU76HSYDW6BMGiGRREoaafZ6rU
8ntUQGdJYnAA2WyT2WFYWtYYPzNmeom6fEJD4neTSNJJWiTtZCnbGi+eEworuoXo
ET28YGZKN17RQJH2GDStyw/6mcb2pZhwT5nrwLMp5fCjo28/FZXg/9srLepxTrqi
2i+6o2jIHo0oNFLnr00GzLb7aLuNkn+x+jtcaAbc9yog+oR3av/GvCSeGScJf5y7
0hvSEqpDykxWBbayXGqduLf2KrbtDyGxvwTAirzckco2wyOE7wtp/z6SqVAzqKTi
HQx28g+LgYgr9R5U0SedA9b09/q0hPCOinBYRnZAZIofEPSTOETKoAdVyhVcAZe2
bcHvkfqaT54Fvc9HS8t7EDtSgnrHQJyp3PKYeWAC1arX1dY/7L2PEHrDNiqmgO9r
YjhtF1uXgTCjY1a4D2tqpfe868i+AdPA/1VmNaPIT88nkyt9nMfugRfTRnooelkT
CZbQEQIxr5b8pDJ4zojam+jXb3pcbfhZ9IBXJGZEBnDigacNdujA/jWz4/3KdPnp
ijnHAjoISHvaE/BNV9YxYkz0qfJtRdA2imRlIU98srr4Z5i92ivBWw06wr2SpPwj
9Y1nEWF2vaz7wshN2uavHnImuCs7WbutAZybadujNxLaj38HeWrPLKsuvgqBIvTu
5cUlQZSjcLBOx885MehHP0/kzJ9BCO+8pisuDvygSTcVn1jkdsRkpsQfGX/xYhY/
iw+pQxhwxJzX8W3YLa4QJ2c2GVY9ddnRCrF5WBocBdbO1p+cx2HTlVEDwQsLcRca
MGCelnd9ptoh6bPxIZMx5APyiiSRm5leMwyYUwsqVOnVUk0fpavHxl7NTNBeQxHf
2IAv8/HbyLEVjoBzc5RXjmmli5+5FDg4hEMJ3nzH6e64b2ljqd4v0Jz3OzqpDdJ3
HBl+7CeXZStndZKZO91nH3eU6ugp0nqQUdX0CLU7v3a0XKSz7h2EOejo96fVcHi9
jkY48j+Z7wHI3l7Hv1uYBI3Dql9mzk0Q3lU2ZoDR8Oa+2v+5ENErYzImIUWIf9D5
d0aDQaGgoFpjQOiDiuPbdk7nTisLueUHd12pTEToAyPvq4J43fU+t0/lWQZOWkVY
IGKIejreiipoIiA0U84ygTiPl4jX4LPyM/nt9dtLxsnu4DD26RUSA52ZseYD0xCW
y/ahW2w6Q0HL6mIuu7o61oE6Wz0oBit497SVqosuQsNyQKM+raDfiPkTwpQ0va+R
eSw0aFrIlFXp0ZXLr372cOPeAqUdolQGbcJ32BIjBhUJ4A430RY+r1IT2cTkkJOx
2tGRbZ+T/tRGsFcdTFbwK97SSqYN2eM5R7mBfq44mO3khZYZtMreaFqCRT89Vcpd
S38eoIC/VnRSLItjDypMRhOPMSojtpP18JuZ6pFGO2KLoPtKY1g5c6rhGDVeaVAd
Eu2K6zIIkhrm2uN8tDJ0dwKtEipjeODNGyDoeWwHzou9rsWOMl0G7ayyIIzNw0jY
G4fYMeU855SLxkOeJgVAObKGyTQDnFUvVlGDNRiDSxotrBiDn/A4QycGXSIY5LCl
bf3OATzaoLJ2Z6u+TNKpN7nWyzeIegloffsWZjAcSkAhk6F2iTlzq+CbWoQuV9LA
tZuuzlkGDaW26RZJZRCwkN9YXftFfRFks1PyJAygbzypzyc3uRJSU+E8mx25Goud
vBWhmYCDBwfwtZVQJ71c5LkiXcoXQiB66HdkekDuSGUbr81Y2SxTD+MaEOm3WUDn
c3AKT5ordk1TcdUYZ2LWtKnebDE6cM07GZH/SguuuIDSS7N9tYoaPV41liERtoqx
C61lHYQiR9Qr77Y7Wt0aoxyBz4Ml/5GlqSJNK4KlpF2dxyLuzv4BjkHGdl4eY2O5
AF5ZnQX4AfojvPGfT8+Pg1J6ZNXABSpkuZLpjeeKncd8AhagSTZ2leBevW3li7Nb
cImDOn09UAwWIojShnLgumu00ZIrL8KsXp+mBX5JGdMNHSjapFJbSF6zjewGb/cK
D+k8oc3Xg2vDRtqkHRX7zEe6UlItwfrNDV0ggitUFPZRf/+dtkp7JqQKq4WuGWgI
4tx6oq/BJQC2PA4S7aVgg7m28Oe7qZiXsffCblzJfosH3bqTi4/TwrWt4KUjdIHa
9FqIr/UVt1VzNc89RnTgSs3xzq1L2KTJRg5QuTHnXxEgBDaBovmikb6NBAiuVWVt
VcWpEww9bavtGbKQEqQLKCl3EsOoUyWu/YWVt0db8cijgIwfPAP/3EBasScjrMBX
mrlMIb20Dpvnaf9Hh3JDJsLSZqGDlGOitg4tGSEi5f/CA7XgzXvr81otheCkykkr
uy/G/IhsogNVJUUZsB8shtHnUaPmMQndOp6GjI6BUqa+l8dgVq+O6Xlf82gKngBL
+fXEymC9XgQUWLx3dlWH8LF7tRKc261SyduYCGW4oZI+OjnVRsJP3zXlaW/zEN6k
DaxIDzdifeL8lzznK/hsIw0bBBFi5lMZhJnQsLByBe0B++IQ71cHpbushn6H35gx
BF0ZBZJjwsgjGm5H5Qfk7gKCkBsWt7euwIZMdNQWfWNHQl5VBWwLziagEg/PqIOr
Zl/2CP8I+rka+59Ru1Fu33prlcT8m6Mg1A588sZ6/mf3dMO6ym2V+82AvbofDdGw
OtGgPQGCYR/VtupDYLRxRluhHUQ7pMPslz1Dgd46UDTJH/V50kXhgVdYWOWGtQ9P
8O198A8r59Fxo94O1o0fGW+0o0G1sqZOFgLsKRvWMv5Nrp75hMWp1k961V7HSsYV
Tfu68Www69M61pmi+R/t7Ehq11cH5yPJA2VGobZIdA6ipycwTGwvz56wFm9RY7Kt
qivLAkg+PoQm6Sdg46jPwfboKz4P3QzTYa+QvuBGLojbAkcy2M4i4aYGqO94obGf
CPEu4OrCyvITAJzcFshuBezVrFZnZ149clmeEBqkOPx7egan9NdDbXI21XD2Capf
IK2xVSRJ5z1hEnvJMAtLNIrJBtqHRwA1Ij90O6KcVmGXHG0KowmgSPuSIZM0T1gb
yaietfIqkVxmhOpXS5ZwVHapVCmRRXkpS9C6R7OyOBatVcZTVpugcGPaI1G2WK3H
Vl70LfesxgI2xEEnc+QhX81vYP84g1m6pZBay3zk+qBj81e1c3yRw1cHitQPIA9N
IOIYUreuhXd7RceAfxbSoLNHFb655nIsvYPWmjiEJm4AvLFxI15rvSYpi1EtbxTO
DE3Tc0ads7K8mw6gQZK6za+2hxX33BBtL2XEGtPl8JU3PLszxnlaSMLqFUlFsCz5
En4jVlg1KJzN6J65GKkxnipup7P+d4KhrCdIlehb2Pri2CBTmfsCvLbyE3D+vTkz
V5OtE+u/B17cGNB1D+nvF03ymm0dUT/0BB1hh+oBiWbYqYl1Z+4lEshrSWaf62vp
YBqKUXfqofX9O2uFUwTMUkeIf18+w4Ge9wCf/vRJRzhjZYbJwp1q5XZKRs8Rj09M
fE18o9+GRQ46sTDFrOVleQn7lz8FgG60k7opnJd4CF+SHDfFjDbfGbICp9InKrAy
2KymxVJ4sRNt7nUusM2DWs8tJJSidGmUlvwvn+335fO/j86fUhqOfML0Hs7OlhyI
C6CR4JSrk8aR/VTnlCiK43vSWx1ek2vCIADY6ZAMfyK5SSD9JK2a2oXLoZDdNEQ3
p2hl4BJE29H94Oc4/XZ/8GqPg88ROA8KkQCplyLeNWe3abSURR1D9z4DI0gtxExm
PtvM4P/VP5iTbtNGT+/I2EqRorlwZ4Hi5yPEk6+WQ0mAmeupatGTPtM3PKvtaPOD
QVLHxij5AEHC5XC99MLVINmsCU6RsN5ju4kK5iW6OWrJgI0Jbxn24VNgd21B9CLl
V8fPvVx7qsXLKovSjnbi2To9uOgiv7wFptqiWVXPwxslvGzzAtnoHTn2HtnzfVzj
lEO1dBVHty/E2giZg0+dCGsv8OeFj9N8TKiOpLfXHM2DhFzR5bjNv5GijxCTPFFW
2VaP+AbF4sWMJtIGK2tkXxePwK6ovkYHk3bltD7IOBKZwh1mjqvdFyXZW3gpDySO
oVWKKEkW+zKt+Gat7jBKI/2do+fyiLELp3AucIoW4zcoX7jS3GRbo8J2cyh0LRlt
Zriatpqln1A3BSYAPjG77mS6Baog1V10sKEjqXJOJG5A/T1RWud7vogd38DDaC8s
5SVPgwFwXPywJzbBwe8PHlsfSxicRz+sLCJx/f+xktDwQCWl/S1TVuNOY1Cydair
J5iRZ3XvAm9CyUIr3dvShPwMm//VJab2ETNzwfVqOrg+jj1yfFbLRj1/4UdSzMt8
ylq9quzmuG9kQvUVWb7n0TUiS8g0nkrf6yT3QZ5aihL8X5begczL3vCZ8qXy/sxV
g2usue2wF7A6Xdk5ClX9l/ODogpC6273feLk6WSyWYYgEOg7+Sbw7Md3cA4uKlXQ
LdyJlQ+kql45b6qNOBwYWZqP0yIsWbRFg5Nne4kR81tu0fONpAP92rc6WYFXWhQ1
n+2i0gWC2jWRFwCocL/FzfX2A/gz380+bzilV0DbONYgVZnqJVkadT5g6YrvcAJH
HsvPM5iUnlPNiIEPqE1/jSOBTrGAw4hoILK95MjrZHGaAzJQAYTg/+6V968BCCII
N1dR9s8LuKTiP7o0m+Hm/AcuJneWxf+J8Yb73xYmqP15DFvPzzgqBR0chTB1AA1s
1UY4xfjhYSDXDQton67XA9d1Iey0/nQil2D1047ngtDdGxl+TNAEC3K0hYRwwyEf
pDdteQYTN542BL3qPAeehwDm4ivm7IyRlMIcPo7NURdTAeTK7Oa+InaCvLW2qZ+M
pv4FdP5n5GLcFyBoGO+vvR/JOLo2DeGc4Wm/w/Dmq9jhILjZJUy+2UEOqXrmiFd5
tsM4PKADfi9b85RbM//vhRyoYMuHnkf92ZuWMethEeoZ+RewXZPbkYRechQNM1xn
l7sx9WYQikjdMNFXJpUiAfbeFUhs5aFLL5j5LRNlTtdH1yLMkmjLgL6FmYxqqTPr
3iv1aH3d/aY6IlB2OmqEBAM5CAOFClEG+/Ax6r+lEGsZHv58gBRmdFb/oqIOEYsy
BEMK97NNV3JhRJyabY4BOkA5of+u48rawseigb+66cQ69lxC2ytx3xuEvD6r6NIc
XoCmr00a1roBf1Ge9Xf3ktbrR1jarBXPVI+6QEUqAnghiW7HkluOjc6y5nGVMJYf
Mpt/cko71Zu6ngwm1oFgeiw6FBtFZft1cKoC4nqVGxfhhaIqeRb9ZRvfytr8AzL/
20oX/qq+2YnzmmSrARz6o4unbyu8IzdUV4L4JPyul1VikkdeAOs5bPI/ik/n/tnQ
lhc4VIkng5Ko8zen3BbpUx7dQYyQLdEhgJhQeLb5kkIadAQ4Iq7zTuYCl4/xGlU0
wAC33L52aeb+hJUlgngIcv3RO/BJdJP8IIu91x2rnyfE4ls/Uarx7Mpu2mLlaTBJ
ZzXOOIYEsu551TmKRB2eubqRm/0WntYrGMdwu0ci78dRK6WrCfHZi0KBafj3uHRY
7hAiiO3spY10iOdMbdeCscROKHxTJ5KUQsoTlX+L+pVwpqKHn1YeqMtP0ouTfhJW
5BhELNTUzyQp96Q4CIQDtqifkjagsYOAmvzhHvvgOrKp53NL5RCP7uCUMsmLEa04
AyFnBulWbYilMEwc2SSLt+pK+X6+DPP3EFTeSHfBy6DAADj65gHK0UWvNNjjZLpe
BmrO/AfUCz97IzM5HuCRzaSEhoj2NG3NlBP52OlLiSUewTu4xnFRfsKCzqWQbNh5
dL1m9QId8c+X4UT20UYUgTHLX7WBm6RghytkNfhXcbx8VY2/G8HwVOHd8CsiGzr2
oJ9hTq+qIB2uMOKLuzZEplCp9o3pTNw2AgY1zySvHtUmWK9M0S6EcM5KWwp//yME
lG9qJze11sT6vDJBe1kDOmk4GyxDy9s4P9b6KJBcRhmgS96fJX4KIrRIoXBKjDsQ
/eu2UMS8A5PNLXDRIY8mgDaI5moG22C0APl5ux6kpgKVR6aIzEiM52PFFEU8+X4M
I/k909llOGQuJm0HNVNzopg53zUlFxJ3wb7HVkaLRknPK9Z5quvV19COaVTcFpee
seFuZCnYRlR9M5VmtJh/9wwiuAqPET8wBhKwh+r/eQZFfPFhS3pYSHaUM3mtsmxw
gzBXh4gotTyovLZ2h32+bcUPDQIQqqzyHh0ftQNR2LpYUv+hCiWuxqj1UbuozZaR
fRGJzoRUl/pZaZcJJBFDPUDBMRPDPLy/9TjfgV4DB5LrxIt8VV3pFIm2BCDo07C5
OGzldZutSR6pER/qPjj4lpqNLOT1512utw0xXzRbQRHkhIo4LsFTCPLTedEkoCX5
P97tPL+Yq1d4gvgChBEjgDtqS+OzbdJ4uCYOP0xn935CSp7mjk2VsD0Qgu2tjE7F
vtQzAn/z1Z9zYpCNPrOJ0QL/I9oLDtDP3uK5s0qJsNwIuH+kP0psh1xL3tewxFtJ
VT6sVTHEUSMl3WzmJsJc7+ov1SaVApGtKgKPtB7uBQa5IYu2p9TR2eTqz4503mQ8
zfqB+MMLUfDVlNaFwRTezk1TwweRcWPDEkPyzL/iOd1LDXIWTYRdclEW1dCeykgi
ib4UfDvgPZD3fvJ9hjm0cu4U5Zkxz33peicNhr8BeMo8oln8IuH0K4wJqPaIZg3p
kpyaExKFOzodBTEkq2CCjlR8AE55TUHPhWMYejrVyMyNr8vJvmGSNgf3Yuh/Gvrb
odVs3aL1luVSo+EDeetpTo3LZvtJs0fnMJXo7C5qQl4/15lu8vivzXoEEr0SPOAi
UMv0ED+yWuJTF99AI2T7RTtIdQ6tHycK8C1ylo5pL2su9a9TcC/RjzSjqH3ErKdv
O8SVDDelPHJwv240QG1HxfTLT4GD/VfP8v5mopAMhDtVemjV4xCpjWeOYHuUKBEe
ZI/PRMLgqcUJKfvElHRHVCImJa81OGm8O68gwoK9wyGvuMpa5NcbpOWJQb2TCao3
Ag9jLlNgCtyxx/FMQjtKfBIn64z7FvCv1lpzhLj/Iks2cnGuwBXM0qiqkKWYlne4
GmCFXjnuuq8oH0aAf/9XLS/aw653XvXjOrV5yxr6hcKdV5UG0Ba0CMaE7yQNAADq
eZnOrwuLEpC7GirN3BzTgY/2L0G+Zkg0dFm55TbOsOUK9wt00BaHkkLD6syrSsfX
sV0jI7zFfKHWOqMEoMB6A1vtdX9obQ5l4NQxQvqhA9nxP7cLNi5TuSgsAa+R6MAN
/x2+ZTPPwlB07ij2sPIpMv1uULEhxOcAazJxSGfS2jOZ97l1aVoqmTppMofNzcdH
c9rIuYs9Ibw9n6zGpBo8VjQhwD1K4lZVHNkhh7hMuEYq2DSuR8JMgFN7uwMeYsMr
xhI7ob2JXiSWwvBX0CdRNUypcI5yOrIdCeTGheyXFYXW8N1uTTfTNvwldm5qcRJF
Bz/poAZY1uLlMcGrz2s6lhfhN928ZYXv8G2r5Rg/FTU6nxa1nSD/X1SAJ1Va/ye2
8+SOK0/9HGF9XuHrBd38jZHI4zxhc/v7Y0WX5KWB5gyProQzIfEBYn86zi3DSGyM
Fs0px4sJiXgLjpBnrhZER9XEvAXdcouAHdYeLCi2LP1KQHo+Ubi/OhMdyVhv0HrH
ahGg1YdS56Fi8ZkVspWsooiKHtXpW941X2JUVLlZKtC7mjYJdLxuxHN0C9fRIvYZ
8raocaT61eYYBnNYMXl+n5zfQCo2PiEr0NMUw8KQ7qtDPHrbB7mDzTPaNQU/ul6U
9h6Kg70WUsjye1KRKi/tguhUYrOrFJ47cnC77etVh1pneL7+oW+qZDMsw38hjBvg
5oxELSRoauHx1fMOHeSZRkgqNEmkoki2ceQPGC5RTQsNgGN2HlwjnOHjr5EXcOOI
f8zgvEOOdkNNguPtx+jcCWZ/PNkZpx7TVZ5wU3c9aZdujPvA2gxT8b++93aLulyu
tjiWTrjcxZQaAixj7Rll7fX6FZOoJR3jcEEWENBMsNHRlF37oswFZ/Djs+N5LfV3
UQ6/ZX4pjE9RuQZ4o5Rbq3ECmFkhtmrszMCBL2mOfyXZj1Mok0ksRxKQTmIUcoVM
mgTQ6MDOzJv/SUgEZJu29aNRYL4/aRT0yLWo6cvrRRJw19T/+cYr4RLdty2nSVEV
F7hjL+STRkVUUHFXAm39FGR1TPmoUwhoR/2RFTI4ljcen/YAEZoZeN1PlY/uatP+
iF/nIKo3xmJbyM73KZcvL/mDYOjxeyg+PMpwjMVeM5vNKxvSOJXIqT3vKoAUHsvN
+b4T77FuXd2axN9X8h+LNeYZJjCSIzhBpZ9CMz7jWO0UlRPj6qJziWTK8WzQRS11
S4yegTFXVU2Wn8sG147TefTDg9igjgsacmvWfzkKMh4e6UDcGfIpgFmN1H0sh6j1
Umok2V85Z40Qjrv88iT6qk+GwcnjgAG47q1aAZY/Ci+ODYXCkii7wsK5RFJO3Ha0
LwJp74XDPs+F/4qLxn6t3lV3DyJAtKU8DbrxZmIOQzx4y+IeACWkxNW/6cOh3LDn
6Je4zIQwdQsBInX0+Wwk2cZTv8EkhWGsxOOBIy+c6hJmQRPkX/asr/hodCTMtot0
Vt8Qnmlwkuu7kDhMSSELS0lPbhep196Lm/3ls8r/NtPSsmET0bD7CmbulQWUOCuS
jdXLHRNc9wJRzObLDREyYud+JblPzmo+XIMa+iJPYcI3CJmHTL07KdAFRwC/ioYF
Tmk7NDCiFDgQ0VrSj5iyBXV9JUjoFs6SMKLXbkAaysXYDJYaIgY0VXacd5Ny7WEB
vS0o1lbr2BP7B6vC3VPaUx1462ccMzEhnTH5WOUlPpEqkD5OGx3cnYfP4kj8YMR3
R/A2RQzFyNlMRN2HKvplt8NCKWaipRJIqasqta1q5hmLxS8eCjHzHTbZqOj6Tejw
RMXzwO8oPPsKzMuirxdIVuK+yKIRwR40/2r4//2VGfPhf6uE/flfdNGfPJgVBzVc
W3dalVuOtBlfCvdywRoGjexd4S2z8uJxpwt2zubnYnPjSj73ZDTQwvBJPi58hXix
skSwWoNPkd76CdV2oV30JiJ62n2UAQ4O0EhdMXhcRKgLsoDMSskPLp4jxqkZJIv8
a8Hp/icNy4TgTBzyWC28xOGVS/7VQuIwaHYwkplkB3/DcZRNWv/F2pg7+J6nJWaw
bF/Mvj1Q82OcXB8uO3Z1PgE9H7NsDPL6mfMXrmYtlUYaf13vWPqbGgjgED1CF5dw
sSZadOUdC6GPp1+jrZd8KTMJ+GPT81RhiX5TBv8L21548lMrce+Vr7j7sCgr1U0x
5aVmankWvhvgAGj+gIakUB/y0KZqHSdOYCETMZIEe/Qci+5VFjc2dl8GeL51IenO
f9DB3KigqCss1jUqwhutsWmJgesQNu1Shda+TzCT0ae9R3R8WV3kYwP9jNu/0kmX
7+u0CawToZVzh5wJBhQmjKrssafIIfYplREEOqZk+p3ENYStnIDMPqwUmBwHMTAb
CSSqLOiNlzthUoZnm5yJJWz8qGsBp2rto2aAo3Cqyov46Dccb3uq+/aaSv33gQU/
g46dAhWITjafDXl3lv4kwS1Iu1DygENkJGIF0mtMRPqG7h4r4Fy/+aRySNuu0cI5
aTtg2XGxiAdf/td6rUyweO9ePaO/FDk7tQOxkpfzo+HNaRHcHxB9lTFgoLnf/LAB
RobtcMvLdsgedc5Cduq9Iv6GiIJdrzDLOjBxdMMEHgLuBILP4RfDTAZx1iE1h8tO
ZV70TBtMmHJCbBty59ipwWJPUClM/2QTCpiVg/cBDyk3YbJeryvRfQ4XIthn36If
fOgk35O02XA1s+id4xMXPNMB1K9gKz6PWLI6JX3J5gHPUN7/f5E5p0YVNh5l06cJ
hoFiToEEQU+S9oncHhEgnCQG2zUSHw/1Bn/Yq0ZOlK+ND3Qs9oKql4j2sIhlvgar
1Zp2MhsZ3GuY8nGwnK+fTlgYonlpoYvIsEyocTGey/Mmd2VMI3+rTbilI/WTQtXD
ce68tdgSZzW1vkYbqrGFcQ4kFU8kwhkqw5p+niqg6S4OMGIePJcVpVb8hE0D7sfV
z11d4Rfr6FHi5dolDSgH/r4JDCLXFzmMCjZFeRUMa75sDhCh9qcGjojZUAqSQDPr
vp01Q2i8nJAY7Hk16y16f+404sxfAmLNUiBhnK9aWbM2EIcKX8C0Z9wwEvfMzA4H
bVAnUZrPBRRJpEqEAh3OXzV4miNPEU7zp0fC7ipAdRkoX+QeMGepf61uXpNZq8u6
L2w2+ZV0KD7bGKiZK7EQWLOYuRIVLgc5TnIRtHmEqLljMH1++/nLO+M77K7abfyM
+WMUgUhftzl7qb61QKY9sypbFPmhQiCuHHcq11JMFevVHe6ArGR7l59MdmyXWc5j
CoBAE+TD8HbAODyIezF5UWvavaKVHhtEIjZSyOknXS57uoI05MSXCvkpFGfFhSlC
s05urYFENDytNSlTkaY9pYe3pwMuNAmN5X3p3rIiNonEGt2CjD+weqL1C4ZI2Ed0
eB6ZhTGA7H++BCM4eBJKEPnf+baHPnuMEFhNMz1dRnLLtaymYeT2JSm6yYmPaACZ
curJ/cqsQqaBfYEdESLSQmXrIdWhbtvmpG8u1JiOccE7+tmGzOgF0RnIVZV8eqpP
Gb66xqyl+t+ERx3sSu7lNZoSvL3AKgpLgcBFX3BHqlaYdAYtkJYO6dzKgewZPoZM
6uUWSvV+5GdBvekFqTH5tWTI0YrXTxtjqg6eCWmYdIuT8oZ6BjqGrfLGh8kQhYyD
vnqt9/kDpfilnmRfNHYgYsLJaLjhc67UC4bxryj2nlKNQaxUWAGFqM3jK/6HQbzJ
769Oc3/jyXmp4kJsGH8br1yNqZo0p58+lfadO8TAvt2mCn3bgcOGuqV9xo4/QPDj
+qVEIPPFNrclLOFwndAWYDRLF5RqlVyuoOOMkhBUDM6FyxrMoaMF6eofTKmN1aKZ
+R0je5TyWdpn7997L3zHOz+YwYU17tKx+KO2Bjr5NmhYNyG0xjd7vnaE7dA87ZQf
whqGjQ8e09fez2wJBVACQU51yYEJFxl5iJe/0/WaeIEAtbLUumYTQSxyfVnQRfWG
7FiNd/ISBGocbMQBUIEa7rh3F4P0m9RbpqtL6rB6qop3CR1wY60JhCWKeF7cUNxU
Y0SDFXwCqAbPTv9Glkehlpqy7dIRwexdd0hxRucyRAJ1ErNOxPjRbb9g1BEIfiaU
6nPeqRzNjFGCEIJD1guqbGl2Y6HcKN1dxNe0DhP2dyLNLENS+MfOoT7PYvc7Q9zG
+OeStkyrSjDEkFxIDX7rXr96YbRE+Mr4Zfmj9x1+w92uYfmc4D70dewamEKym8Oy
8oqVzfIlVJHzxOtnsk8LSaTVBasSOm24CyQlISXwSsgfbForkBKY5Rc8A2DfaskG
utjei3Y54sbCdBUAFCNYKPiZps/XlwMn+bZsDSiYAreGeusjraWFcfCTwEXAkCqV
+m7Yv+jNh4Oh3Qj7HsJ6Rq9EoIBwuJKdXX8hCYmuIk0DCBZ+pxcBrUAYdQ8O9kZQ
1OGRvr7XIDyFdiqdSsue02zVtzEpd/feDDcv2SnHnsOgixSbgXH51bQbRXn0axUd
eljWqnXJnvlHeL7lkshk+qk/RlsVkci7kSgoUbzEob4aGmqKoBa+RyURQ+jWlGCM
uvlo8tJKV9eaHmFQ156aLswTa/O7Q7Cp5Xk2l3nsNX3vGZiELVH6WE+MZmTs5PPS
1cMQVeQpebi6DAUFwrj1L5vIPh6BukfpI/xxjpBpi2ujJVsYFMwNMrwkYMtyYcOQ
gvY4dC2CEfT1JqfvYJrEYbxQdkr7qnHMZ4D2KwKlSqk8ceYbWiCa0810gmE0mGO3
unkrM34WRy+p/IGNWkx8S6fl9iH7EH/04WwQe4oasV+VDEQ1HCEvCgVpFw0DTrzq
o5oZgJleWrfmyczPLcBx0ykeI6/3Zd7kePgLdofOEjI8h6ocHxaxKbSxhv15/mL9
3tlntp1GgfHasVpMG3Ry5hTAy+J1lEbo5MGoabVWgOCKWUERanEyA85ZDjeH7R/9
xaciKwWtXU5EdhUrqyFFPZHZIJWfRBhsQRvs2zBfQjeWsACbN83jOSxnpq1SbLzR
sWJxIFB4tHws5sVZGPx5kLUMjZR4Bk6qV4XKja1+tLjod79ABkpekkmzNop2KsAc
n8ZiTWWu5RH1Hc9D2YBWbDSjs/a+5PwI9gJI2V25uSQQhn0RqAMl8wPvGfUtxYw+
ViVpS2dUVKv3H1RYW0Qu7/9E6mbqAIQcYLA8S8PBktBHDWksQfI8SKvnWBd8BlxM
m7iPrlMjfb2OJbYrwl4KpAk2+iidz0MZpdM4cBNnD4GXow/NNeWh5FJ6ftYvanMJ
LFuL5UgwiN19g/lctLCYTs0cdBFzNN82j8KqK/v+qydO6ROZHdh+o5AE96pJDPxB
lMrzo9fDppV2fVy8K/+ZUYPE9dOdQTuWEcHOzmWgL3qg2iXwilDW0zgvExa1MNuy
CT+Xlaj8vun+H4j/eCmZfADtYu7JXPCtdcsrwOOUNCacMeq/rclQ/xrEdJF0jebM
3azpBG9OhGjeMAxkkxD5XXPoU4NU9gi3hDpxk+5tBLxsiurAWpiSxg1nlfRkxCzO
n0qaLL09jb2NOzKTnRwRpZ2qMctyrznjoQUL7gLb3h9rk79dYqQC7Yu2RUSRc+2z
Sxye+yC9/V7svd3/ecTrcdIOV/e/j5CzU4MSwlxLbNktJ12uYIi/mXO/gpYhGqzf
cL1urYpdkvhDv7AWfLfpz7VuDs2g46GkeVkK0X9EP2ijRg3aqZLyvy0a7ErpaQ1n
WwIsCIWhT+h9zo3CFA+N5tYEY/ZlXX2ls6XtdMaXjarC2sP51Bw/iig8q4LnJr5X
33euv8eHp4CXxxjpkwjWywCTmh4i6aG4rerCEt3u6sSMDdYrctx+u5dGgIzR2dnF
2cCrn5mmm5I826mLEu99ZQrEOkhY1y1l1UY7t556Dwr4D+6H8MiuxZ8DYfEOD+zl
YiV0na4TWhUl1FAV9C7xSx/kPHKaLnP65x+gKiGMR80rRPcganVpVXw+Aw+D2zzN
5AbYFboNB27NKf3lvGmL2rm1Y2WiUDxj+VLfT03DyW5N3lyNoaEQFnnWOUrzawef
p8uEWGuZan/IXIqcGEU13TGdzGMPjwKfRNm6El4/7Z2OeaRaxTUeFl0do5xUiBxQ
/hJLw/iXKFTjaWRLPUniY8a031FvWPfzoN5fyhZpeJOzhXJBSbGf4val33t+squz
0wVmD0jAL69Cu8sufdR6+55Hs4J/ijJrnEUuxlUZsSykv0L/4jQW1VTup9iSHa1a
DRtxUC+9/XghHOj0xf1MWtA62VmEHrD9/cx1GyjyUWpoxRWZcpwsgQPUjH8vUxCO
7t8X3xb4wz8ETFcdM9AMqBO2EoCbaZEPtbL38lCFL89qlgCJjxRonlWpng2XwaYL
lGvZIJTGYwahL1nUaWxI4aONjHbBijJNJ+T3wNhWROpNf9nO5XpLwok3wIrkuq/D
Y2kDUnuW/LJiZah9+Ztmpi0yNpPGq87A7oJmOt2QGAiyipvtW9ILG1w6PSDqnXFe
xj2Y8TxNwn3ZydCUSAZ8lvF6bpW3l37W0Cj+XeJYKvh9wRtYlvydko5hAVDktt+K
MQJhiZpvr2icQaQZxL1G0nsXsk36ICaSHuxd7AOES9ibreGk4PbI0amVAdT/I0WR
d+FKCNdryFkdqdQEi64Pr04XA+33Y9Nt9PPBoFfMDlVWcnXFXozRbjjx2aG64bkW
Eiq+1SQo5PIGthhd7/2QAwOEkhyK+73Tt66xjOdyNBx94X7rjsy2G+/6PBvmNFwR
L8t7Uk+PvIPaKdE009I3N56jDNpxiUoz22CTwbIQogzhOBjnYyQ6g73SL+p+YImO
p9CDjlBAmj2crT2eKI5as8IRxnplPRFyBxneF4rpWxDkAVJqDtX0JIpcpZX8zxe8
Ed8i4r+P8ElDq+7jZ/1qyuH6KEgswats0hGfuCZUXEvr2n8DLesmbn8qHQ7Kdt/d
EaZVOcrQpZlQIhXn08fam+lebhHDeAX+79paaDZiXkobh4rEw4JRy4pNyH/7A249
KRfkk3f0CbBtNYrZBr12jrxDAETzWRVpFR20bUeAD9rkQd4UCG55doG8X0cZAYhs
R1tVNY9kkMq1WQjxoo7ksqJ4QvL8hshslB0PiQrgTM9+4LoUTNKXOzXtE7hgttlg
oyBejak9rf383kfPiIRoqBUIUcDw/neHaIoAEM8TpQYHuOlpfaZRF8yb00ZIM8Ey
OrUe59oVV9rdMwjTK1zLoZwxnToK/brIh/B4r52LU8D5lqI1DV3/1Y05l3hulDJF
HeyzVBNJi/hy1U0MPFo0vm3RxuADekNuD+nbzlwKkqXGDsixekm1azAP48Khxgkk
hdiuyR6wTjOHOfZSYN2zOeceLA+eCEUpSuqFYUqs8+z6nvf6rIKzVGvWvlS9Tuyo
hrHgmcuXRXrDMH4N3OasfUwrpc+leQylJ76BJtS4PS5PwPjRKoqifAM3Q+SK4aF/
wJgJIgIjm+bPCpj70EGg0IpWL/X+6OKZAeO17bXnfUYOYk1l3fMrWFDhvjwX0qZ/
vMSmwnnkv/Lxq4/VRiHMVeFSqys6LE0WOneHP39wqB8sN7HQkfQ+mUFRyyQVBi69
4UzCU0KjugGaoyqZ1bzUcSG0rIXIZemLPTl43BnlxGppSoZRmC7jGPImMpSk8WNW
3JeBDcr0aoQKM8yiojnQd673lkl84einVRq7ufz3+41d9u7+1UzfItb4U+gHumgm
Viiyx/cwWsmhT2vSZBS8dE+DtNcLWlJIUef8N+4Cnqao/gDRHYjTOm/fxeYKQhGl
G+z1CjlxwmXchud2SgoT4+ihZCtkYlAc5EIUllcsAxZ9bGPgEfEiZQ9NG8K9KavC
PVN7H0Rn0LVVZCBLblW/34x2K3JCVEwXN3B+WYtcphflg31jdh33DrLEKc5yFPMz
llpXXTBAVxNHZRI0fsP7iJRxgyhQGu0nEY6ZMpAIBSYCYJUXGtwxbYcSxk7mVcLM
zS9Xb737Yy8CyWYkdzfW5LEBlGTNdbvFa+62Jv8bTJN63zTfk1pKT2t8HKejKj//
NijCTKcTb3IqPCDgGdlmEz+CtXSujrIdygFYO5JeTHmK7O/2HX1675g26Nmsslej
ctVSpsXOC30g9MCNllXe82GqOf7jcXXK+1k2jI5PavR4JTm9Qj1wve0qkCwWHLOK
eGJBsJvdq8cxlc1rgzw6napYck7Fz8CL//7+CyOJBFGaGkolyWKcF0+kmsaZoj7v
37h6xDq8Euwuj6Nd8DNRYe+501C7AG4L64fSvKdvoKsbBb3pyK15w2OgL3Ii1deu
DL1iHuQG2abmeLuuQFmvLbBcIwqdgrRfHRg0uDa3HXigvfeESN54prGjTCFoU5Ev
QocM/V1UJ9mN8IVw11eEDVfI7MmiWjLT2ca9JH27KqbKkEGMGpNkw5fNUdZVTwcY
+bj9XqcHNNwAWarnz65ZOMTo3NQcd/ydjaMR8TAAWK+XfJjxYXKUdFOhS7LppySY
u5GRC51FvryQsOxsc67QZn5KmRnRA4tzpCF1wMPincTh+K0/p8prJCALcTGtoXNu
LSR68pXMsOT2gqM2SuH1oRqEnCuBmvyCv3PETNAjQoICyN7YEqcWo6EguDLBDvsf
DufRQbd6VmNISCp/gwGtzY9uFs0sKzX07tEf5GTRT7eLnte2mXuFoRdjuajHqoOz
gvnj2TLrQ9LzI8B8B8OB8KYmBMTmlfbleRCRIs57cgfGtGM6KVP8D5yI8+Wj5vJq
dH99xq/F3r47CsXhW5WMBI/65jFVPUbfJfPF9tOAYMFGY8J1/m+yCWUyzIOfKce5
rrhCRs+ismMaS2vO3U0QOxahHILj0NLah1L6nbQW6MfGPCBQMD0ivaM29HfLFPIk
zVYBCkQyyoMEdqD4JYUv3uD5mB3KWmlS+38OLg0Lk6dmpHO532q1uDQ74CmHzgNR
AarRA0jb31wRV3+qMtmA0MCVWMfTSj29dmQQxbEMh0ru/IdzbRQvUWQRcyC9esPO
TnEt05kZdR/cTKXhD3XLxoCmAVVhQ/5lBAS+IYHX+ifDlFotTOWRxj8MrZwEJuvm
H2JkRC3pykT8w34FySYSpOwf6UGqMBDmzJjoRAqu+i2j+wfKUoNHs+vRTKnRs2Kj
vTgcFfKGp3ldOZyXLnuHtvdlEob9WGKvCSIDlBoWw0Pm9Hnjv6OfZwC98npzj2X6
SHg5eTIgCvrmLPDcPM6HIeDCnXF52cmLp6xFi75c2fGAq/KYnooUyuuxB9aRohPv
79+3A5eirb5ROmXxCINnzMwevGNGLQ1nJ3JPqG7tWdjkg7S4o3a7aQoU5npVFERQ
7W6FVBXm+LlveVxwLvKW3mfN+QbajGORFWQteBTHJ9xsyCr9NRliao26auhl0JA3
6eiXYDgLwt8GJi7iFNTcVr1Y7FImf7IG60j3DxVwFwwYYrsSvntD4tcbEl1bwOre
DF7Vb3bHK145Blbi91Uj54tQkqAvZsMWcmKyfONWCXhXxI36d/l0Djdt6LSTtwmD
Z613PqB6yjoa7T5LqQbPcKkqW5iM5i4orIWItarSmEd+HtP5CUrJ7lGkUaX2Hewq
lXIpzBU3xoWf57kaLCo5J2wBfSSt+lgggI15ycI3dXD8xw+5NXPCB+NhKKDNTZrt
4X7kiUvfvlr8CFPQF6cbMlIui1bikiThJ2W+HdKk2eqIPVPebF7iYqG+eQTXFYRO
kEiVYybq8Y1118ZszPu1uXjZs5342FdI9ea7Kvnm3DPaesZfID0jeOrbEnbdBGU1
hOwJidAMBUaN9tp+6QhbJwPBChVe0k3lB9J4d4lKOLQHVHixRFFkwDU5ocz4baUP
2HLmmx85ZseJIECWfnS5JXelghEeF3LPltfFr0ZKNEA74bl7F+OZPURG+e1A6OUf
a6tziExMr3cexFdjqypScMDVIwLpV5AgB1ZZuoXu/lEJwmLWU28MicisppHqsmW8
wE+GHbbjN2gwlvYzzitAmfBXlQEG6YxYGDbR+C9tFGs/RZVruxLs1PvjpAJQ6qMw
YJ0xtfn7wdRMf1UoG4edItdsKYL9wGXO6QIdA3diMoeXrvXLI/Oe/BuJkpgn+A8A
33GQFzr3enYfF1SshSL8B7+cC/nL8mWe5fblcbVelQ2c+AzjCum2yIZi22+kOhVW
snH7tCxzu9sizT64O+kXYQBfrcaG0wA+VGm1bmSEpE/vtQLCy7mBcpWzf3fI1+Wf
D7Ng1NHEr/VEsb/Jtd8DF/66t1tfj3V/SDu/x8onIcRfqfnFVhljFjbVN+inXNhe
Soyl8jNeO3HANlAPOtkldl6/3KiOYIy/3Ea0tWzwiY1tSW9TFe9HZ31IfLA8blh6
gACEzdAm8ScpKaLin4gGcg4zz6VfkFhdCtD34HrFJ+FQ2aBq/cO6lUQHIFWSHI6E
qZxYfSdmf3tNAYXgqh1mD9qc1pg2/6QA917Aib/wGbrG20eNAEnKQRNybdyIhRN9
WNr4JyZw3mikxTJ9tWzf+G9e52T/+/4p/L6dl09Va2F2dQ+HTSCINVDrRaq4S/t5
IhrZ1RVd9c1dzyTTJa65D2lwAIXhnXAsr/t9My6lsLsgSepp7gb501lqUsZMCLJy
wq85vu18TjTFA1N4iftg5L7lqmQY3TWhKC+xIGI6mUFYTks9T2NRCkzYEbfTiszq
MbnC/CgBDVBa6wHSaBNWMYckxYaKzl+IbB8CzLlyedJYOBNucIY6/uS3u5WMAQ9s
tpbuXLVDel4fOe6u90cr7oFEwsmWhTCpVaUe4SH56NbFPg7LugNrwf4JrLdJuiAO
AR+TORcIx6g0WawIPUiRnbIeBIKXDPOmjtYmsBzSg+iop3c+RB7pUW98ABoJy3di
DuTF6+aB2e4q/bXgpuiRxKEsVn4/xRkLJdKbYR73x5VQtqWVSuo0gZNQ826C++Sh
t+5qfl5dDpRUUYqXZoUuk9z0ovp9L9jQkWx3Q4MNpm8LEFI+Gik2dS7pUJysw3A6
DsHC6YouoAceaxFjegB9U2+m7++43egnmEUmYRKZhxndyrP3ZJISrXXWH3HASjzm
Z8+a1bPlP51If1tzfOf2rplRowmzNKIchHBYnxN9kZunjGNW7ThGOZv5/sQ6YChm
fejsLgd+gMx5m0v8yr5d1TiJMYvXUPaZeK4e6dq9RxsNle6LNhM2tF1HD52iP2sI
fn6uDEr19Umi8aWXl5Gn+Cj4E1rP/5LTur0/qfjaDcmWbIe+NOtVOfga8xwL+Y/h
49vgkcfijJFbewEZT7iWOAbPY6bQmMuc/sTxzSmZ7LX6arR2oidHe65aaGmOipO/
xxNUqS9mmN6cXY9y4d4FAiDHjY+1b003JS36jI3RnHeydTsYpMvcd7e+HD7Itkzb
xl9maNKfAGz70UZ3dqcQt5Pk9C9QrnrN2OsE/DEldcxOQ1mNL5SuE3Y7xInNFSFg
jNnNi9h9rN2sv6NmiUM+9JpaHEGVtPBZjAcZdQh5JywjaQfmqof2gkOjP4XAC5yh
FagCCCof5jlBxDKT9PDsy7ya8skUf95K1tRA7Qnc9Df67IlIVpgDVIrr1DMgLVgZ
EDdLsNwn4NcwI1LcZ5qWTJsJNLIAfrDQuyWlHv0dygr8DnwFnB6GEEENPUQpXpBx
aO13pG+9WSsL+MhOfcqqC/UyQ4gpj9NGyGMPzws1/2nbPp1eeLb0M7U7uzCCxXLf
K5lu7ad5tHOAo7jY9vLhOCFANwQz6xjuqpi+5e2t9NgnLJTuQ0XWKBVaRwcmwx8v
eiTaPJkqT/i43AmLXa4LFRDPRdZaFACCqfvYCGiCN7gPgQRTQwcI00VORSVn4Kir
mjMuLf5bSFnHgHtqI/J2NSC2qZGnV0lTSx9w4YkBH2M7uydCADXitJtcpRtdyqCF
mbxsWMvQIa97V4Gc8JD13lbo3kSUZt3qQnL3G2j6pGJBXSD3gtXFFr2Kfih6ebDu
et1c/uJXAXsfFrhOtkcIe8NItQAclbh/keyhzjjTiPk/zUnmIzdzajerEZX8u6xW
bXUBFwO4qXBo0wa2qiZlARTcynxFKDTSzm4APPcNvfc3cXgrjh0hmR5pIlnRzuBq
MpawsL8tWd2IpspY9bdHxRossfONvikbn4HFLQ27onh6PV5n21Giz9pMo8Fj71Lm
OhTrqs85QIzEt9IfDhEp9sFoVhETaplG/OCoyh6npRsd9wDGCs5dGUcIL1C6SLnp
sHDCffeZIXKARAHueTfZUt1C5reXlMSlm0zXdtbFx97V0f7t7pOOE9OK6hYovj42
/cs1oVHWo09rIJd/zpME5LFKKvj4XKRLcIaFxqTaL49H358OIaQvSFT8/uic700l
i4dPtqlbbxLPKhgUWAVdDZ76eU0mRZmrohnrPitSky4ODoAx4J1L1hq6oF4iLzxG
3aJRp7pa06C7CmhZfTxtu3t4b7yybAYSEF0Dgi2XHR7dKTj0Z87aFAQoSQ6LzXdN
sD3CVAMRa30SU2Psd28Nl/NQRboYhVfcOvuc1rJszArQr36XTvqsMU43Xvecz/x/
O3ZkadaITV7fgfdGJ7Z/PoaMF7RACxKzRdWb088OH9gCSCULucsgFwpx56foirce
u+Q6oz+zSXhgnVfgHThVcGQMDHaFT8zvn0rX+26adNK86cqN/eISWJZ/lshlpVRy
7fMd2ymDuDcGf0Gp+cdlZdt8xxaIVfnpZ/LUKf9FKl7SYBrsRg911ihDf9l5Z6Oa
ECDl3O7JHWBI4PFsnItMutcW0yEbacZWOqXsQWqhNDQRlxsumo/Ezt9vHxaCHASg
2fJeawyZcSChqG3rbhC+s1slBli8/F2bfVlJVzUBj9LYI6NSr5VbRaH1fiRusPDa
Vrh/idSO0VG+LRX60LXGuPAz/EBNdhtnSUCq1Kr95vR+Xu7PTGBwSoVQnqgL+d+r
AD0238QO+hGbUgo9xK8l0BoTUznBhzItOpZ8MpkEJYgiDFVk4Lp/CBtF9tEkChTH
GRvacQw+gQ5ShYVhsi8ZJhP6INgBESwXf5ZiZ11rvGgFL+nUmvm8CW5X3LGinhQq
XmFYq8rrKe1aVPiaIXRwrYmfC7ghsR8HxMNbe6rKZrYkAz/vBjuqYLgaJ+asi+ME
rLhv0Jv+n50dSw8XcC6xw1wuxqvBId/NGmZmEtA4wPxC4XUbfBes/aDoteaq8mq6
0WaJOBVgIjPc84uaJMB8yRTO0zWLucECpqaZuiWTT4M7dydVGHtzTuQy0wEeYrDj
9lD8QsE0wYUZaIGL4ASPbF33HjTOrVAG5t+4cH7Yzwjcoy8HHF+LC/HKMmXFiPJ9
rvJsKuUp31CdoF+k9ADoSSfzUsWcqxyTH6O9F/AxvsB8H4q/AjtMeVW9qxQptP24
m3YOwaWDX7R2pp/4NAZXhdqe/aa3Wx0e8ErGCJOFpQ3ADTsLdNHYuTtjwNjJ3XnW
Sd+axrFXMDkHhvnrq4QlUMtwBm/QbRSx+oI8grXGxWkYvXv2xUX5Rxd9r1JoiWtw
C7/rBRKZHCnPsNVUQQweHR/H/bcD0TcW2d68OurBmR+gE20Clo8MnAihuAJ84p1D
SvnYwZLvdemiyGdR0+NUivsEDEH5YByw+Yh2RqE4prLN25kbW7Ar4XQ9BTkLPgbQ
JBqwU0md2pQA9A+uTZJNfJRivjZvW7oe8GWuQzW0cKjwD1ejTGeP7Zn++QX4FJTP
AuIpp8MceJhZv9G+zmlruidnxjjk7KslpelUHaGAOUNSoyvOuUHCjII7vswNJ9oo
xY8YI4Qd43j5w5HoMv35cxI+KmbkIztYJK76PBAlj6qK6cFvfxCCOaO1OKQHHazK
nLhMSKuvQMiUr0AyASbIu7c3XtTx3bpY4DqP3vxnqbChW5UExbzL+kLRUVeF58G1
Pmnv48ArphnfvjXgGMSn3836skku6LGUOxQQgysYAzHreHGU0Mcuz0XmnIGKni3R
heb/BJRXfGl4PMWEnV9qsYYAfD742KYSLUjP/3+9ZpxIxD3CYXoqV4e9LcB2Zfza
j9g9nD+QUy3eZYY2oeo2ivIhqqjedOkOi6C3+4yxSPR8jnPvM0zuO9eTbuvT8C3A
NtVKolHZoIneLq9NgIqdWAXT7kV8Lpoj56PMuWB5AnZ6xErKP3IWje0VS1xFPeZz
hKrCCtzIhQx3Qj0cdO3LTbs1fG4+OnQeON2jz3CbK8NYglVizfO6aaVMDNgdZtHO
J9r198NoDqyeQpfgQKz+9tR5zlHqzYMdOUvIa/fO9Kq+eLiEIB1iSarQx5mDC5pg
JCIfBItXmgmHI55hc34vCMOYY9xgSIr9YxdOk/fHRo+rS0uDdt9fIdmqQ9bPVFaT
9269ExTy6EJiPtyZSGqukwlBKOblmHfhBrMnfhXhosbU3EqG1V+sH61u3KGCwodq
JWsVPL61U8sMk3HQ+kZeK4/nrEoGWSu6Ho53NHj4LmbT/kCy9CvzXW11iBBmugOb
21mw2rxKsrD1xDghIKsyefMk30/LCksOvIcEzUyYvytIntNEb9rzrc6O6wh4FzIy
n33JJVxpJqKvCEwG7B2ixCT/cGVBlTR7h5GBPB5xiapItIx9c2ArvAxgwcTp3GFI
M9K4GL82B9rjcThurIXSY5kUNrToceZmwHQGCa/r6phbjfaCzNRd1FelBrcJpVMS
KXdv57PsnNQHj+wRaKdfnoTPaon3Gdshp4PHrCUV4h1lXS8t6ra24118sPd+hVJk
tnex2kO8BraA56K1TfKVwbaTM7K2EhOWUdDnfpM1pOxnZFftb2fdmsUKxqN1v3Q6
eep8E5IzrjiYzlCENySegR0FdSZ/+V/CnwMfsYr88613/p7OgZg2qhfo620Dbtsp
5F2aJxgghQ2zxvDoFwM1JKnsn0aFhcSldU+K/pRRqmtkAvAogfkhCWMsTrVoOhSB
uFADj5MCNloTVLj86xnKti8dd/jAYZZkGIZOKbDRdjSI3ZGwkpGaKyROgnQtbY5X
WIjjQElPg1mkUBazvRoX3j/UUdnU4R9IrEZ4QkTgjTEF9X24SLcqGPArK8R2iOic
EZKpRYETqg12YHnjPxsoKmC+MtLb4lysRYEKSfnFDUikbn0kIBGwlGaI8LEMgYAR
aJl2yRMAZwR1HazfoGafSwx7/e8RYVM5BV6lvTTiv8QnW8hgvjl5/EObTeDM234s
yXA8AHuGLbJ4KH/NlV6YBTzS+yOYXXFLCcJGpfJmwMm0IrDBDk7zB/hziSuNubLg
zFp/vLfx3E8yTDiV0c9mGbi23fEa12TYk9fZzVYcL8olkqsu30LbbxirJ0UMu3AE
LEMLJ7vso5k0K+hHIu2+UAANAKTrbPCw/t4TQoqVtLCra7SWZP7IDc7EvamduBvP
qaG+tEpgRLOsiMLohWPSKJKXJbpZTbyQ08/LEVCmgPTMJk9jkymvNio3D500dlU9
edXl+qlz4ZQqzDZ8xp2SKL1IbrGH0cHRjj2DbJM9gCPjoAD/Vx7WBKYoyFwZyS0e
Dkl+YoujtGw2lP8B42V8NYxn8ityrud9T3/CXP1pFbQj0A707KM5SQbP5flgAdZ/
MwkMAMzLWiKf8RQv40G9dlz3rfDOb1mAItJGc3MJcM6Ibf1BL9kSH0gifdnHzC3F
DX1Jg1NVRW1D03H73w4xJLxd132kFJLHf9MRXIrLOLpsrbbBbZ9yn4IFFG5oPuV1
ChZKXXju1j5R+6fueoB89C21uzT6unOLdpvb7fcnOu9+dpZqyMnbN2OzHDJtMIY8
FVhltpR3ydkh4kMBPBqjeLaXJQ+qECpPQgAsuwYMSN+kNcWQ7B6CMer8d4viw1WO
p2kEQL0yFFp+SOomqiUDH9BsUS8ohow1jWmRxfSvmBOz0WocEmqkzshX7nGE2JUb
D5DrBSxri7Xcw7Dfw3WmXhxNEGoo8nWuPibSU+8wUQnr0YpMQ6eksqllcZWHdX2P
gO/gAu6d+cnuOX1xaFVRA/lqxMCzOf8+/5orco3xbx8K3BEzPfkQGBzqwHo9Nlux
QbP0tG2ogfpiHiDtPSW8dXo+oLi2OBqgo1Xe55e++wyoOge9TlPM2pjZWgjttew/
zrACFlnYnULfulbU4cn/2upYuyd73BGAaV7/VzwGtyhRO3Nf+HGNE9gxpKgM2Fp8
Yf1iIcR65GY7pyd53oHY23BBa/7J0Kci+igFdUzmZLJoJupex6m9iZW4nJGAX8gI
dpSqbLFKwCgev9mQWmHjWgrtW43DVtkmSjSAI5ABsGdI7+/sg32kiR9dIpagn90R
PvXDOkGhc7/rbPgC8fK4Lo8j777PVKbuMXE6CLjnv1qiVHA1bpKSsPB5+fk6DjvQ
QyZCsXJuTPnnHW7+pc2+aMwCWrN0Ma/l5LxMwGa7IwQtsR4AATUUBbl2b1dF0w5d
xK+CFTvXjqiK44l58w89iOhzGZpylensCcQfko2g0+WkVFVJFw9NFCNNa3MGT6GI
tbJQDS8u0Mlk4T3JCy6k3kAbgDTzKsqNqJtQIqPc/1+pKCJUyax1ofJPE5dDFhSN
Z29hhy9eC6pKFcIm6DM48tevFexdF3N5Tpn1gBZHjkyoPWZtbSFAcLUiCj9mmo71
wrBaOHp7GPYp0WkqlY9hO//dvSC+/6gWsWTlTVfhkTf8SntbW/+0+zh1V1ra0xVy
uyQL9Ca4dYbXPrbFnI1p241aO/uPi9DIM8hAUFFkAk5MuX0Qnc07yB4agEVJA4jx
2U4Xasw3GZqxBbPTL/RjtTpa5RnCfWCmOTHKbaKju0Gl0sbb5N2t2gKVCuJ86j8P
93jIqdriN6iyOxPvxxNJGfMs/k5/81iwgQtiYnsTtxd3uVJqdccF0LEpm3dWdM8l
iq2Ka8fe/hveeBezyltzqaYRiwmoTPcL3zlUp9G4Ok4wwOpzZi1f7F3UdgMG3ti5
zbh/0vF/wbjEdYa4j2QP5RVdML2NCJp1kRcJg/GdxhIdW0mnBHorZwUc9xoZC1Ej
cylgJzI/9DClF5LHxpXUubUvdRIkxV0IY+FxbjCvDB1S1VjY6XSnDIj61DvVtE84
DHeoNIxm5ib4Oo5zq+Q0t7YDHfCgy6YVTJNHJiaYArGOF91JtxQEVQ9SQM+uYEMf
9geLoYoJP3Rl74SGM3oMErcf/3rLQCH7GZ9ieZ26IFm5VwjT1FRVdUfnmu9Rdh7k
B58QoQE1yfbvK62VK6rSiSgwz6Iqq5LhN6Fpd2AzEcWKZZUwgnuryUQOEaar6z02
syi3IAC6UKfSSmblNulU7JNT9gXMU7HWvD1BF60xGCtsjXGe/j3MAkniGZBEGLIu
6ZjJMYr248zenk41ZFgTJ/zk2EQnrJL2LigK8HgqJPjlLPF0wgrT6ISbLgcEL2Oz
1SxTLOjOR7J9O0op8kHT3gufV3z8uWm0R1TjZrORBiEUj98OTTosNYTeEK+3N07y
fEVi+PDbq4Mk6PCZnLvG0kNLe/GeR5mAax5F3VXKjkTr9iHenhIcIU59n9GhZQx0
rPqQOqvFxa5IdtQlq+VriQESp//gsJ8+LEBiCTGTWYRvNcUzkxP/b7E5qbZbET8F
2gFByZtZRXPQgtlrpN26BitXpxpQtkhAEsaQqDhcH4mA/h56da1UPB34TT0Nlcce
QdiZAQnGd4av82Mr7Dx/6ea3EESFJoy31YBQ89zA8TcdogvnSsqOS1hlvdpxRzCI
ZyP7QNyaxhEQjVII4CKCMMyKiplc1wZfwU7FsSBaYXYAD8PeuERuA7DDb7MzNLD3
gZR9utpJZ28SDEEl0Slbv134VEWuFuVpKvt7RyscQRMKgq1gFNB2Vev8FQRbpJmM
kYQkbLxeDXQ3yDBi3aQiixDtRS9omERJm0qazDFtXa00mjy4Pm1GHWlCZIsCvClO
`protect END_PROTECTED
