`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJHzwWBZk+RmgodMXd+G5NT5Ryt9TA6vD7yIahrSsbVe
Wv6J73pkqO5+EhWgOFNIPhKgOrAFIP4aXD/pIsfn3OFAcanufcM9QOkPTQkvMDUy
BcJLZY06J7MHSuC3IfliRvbTTUG5f9MUOz3g5gDkgECxtg36t8GSYHr6TlL1TJq8
rjfjc6kTLkp6KYdH5pmnXoH5ql19kQjYONgIa1EGWuLgyjgT+iUrOs4jl/cvRfu5
2x2akqAC87p6Vphrep5Cbg==
`protect END_PROTECTED
