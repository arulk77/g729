`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJssgWqcVifnNR5O5JNKUN9b+UpvDpa4mYbYFSlA3dif
4jLS6L+YRq4IJgWKh3VTHDgSud3h7fMF5s0p67ilZmC00cRP2Xpx11Vh2qpP4qrU
XIHiZmiUQlEjZ66thHLyHcGWADeDGWD+jY50LlKTq+S5+pWhfMlLJ91BPONvVb/L
s86NSWMAGsHNuRTXYA7Uyg==
`protect END_PROTECTED
