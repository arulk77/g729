`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
KnZguEr081OCiLHu++Al6hGcu5gHjJ8L8zjm89RBT9wQZkA1QkBB2SNapfJtiIUu
LSWoJxOjorbtppM8dlX6wT59wOVdr745CtHfUzffzsfhC+2jEFe/6J6QnJwnotrQ
xHulN+j2thZQPuyiKulNaVRTLins/k4ut/LED3vhbgrSxlTF6ikSV3ryj+tBPSTB
PnDg6VTdgeAkh5M8AQXLusnBcpDVn5KTHTN2R8LVRtWtghz0FpdKdAgTx4WbIXpm
JJkiOjotwnNckNCsG+jCFF8RNT1pQJdpQdxeD+dU55JbNHZ7Q8zh6jDihTmlRr4t
TxPq977QO6AnRt5pBV79PAPLXX3WNvvjAtu9LO4rdH6145plyz+NQwqEpoCOzQUo
TWk39CeeyIKnIr+CCCJkbw==
`protect END_PROTECTED
