`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
vQ23N4UIBEie5tV/1fim0uPYsgt0HWfCBlyJmxTVqiEQSmtvnZOSkmmGQpXH5yrP
sTVBG4cjuKVC7v1QVfh4pLVEYO/orZ0mrYc4lPkAFlzKw2DgCBOfLPEgQQTt1Mrt
WjtSoebaX0lyP4Ye3a9SsYrQ3CyOXDD3xmfA1AE0ec9bFu1ruAQarl/93CS89GPU
V0Io4wSCR6SPfecs71lzEj2VDEvmZNOBBfabuobZAE5hkx9OOzssl10Kthm9qKlB
AYezrKfuiKMRqAxoRTaLp/uDTQdBFxTKzFWkI2RU5VdzwNDZq0PAnACtxtdApy39
voI9aLK5ZJ0Qan3kdhpLJn8JOluN0dlKyylOaSVf7It17n6qmQoFObKOO+Sg/w/v
qZNkYXrt86Qdm7P3lgkAuu2AjDnWwSywzZZlUB6xVLioYLZzo9sJc2lsvu2HNASE
qzUrH+e/K8MvAlgqcMk25eq08YaXtVfZSzRM/iv1XoM9GODri/cD4Bu8d//qQ5Ie
RV/+lTUMG/xSBq6HlwsR16Rjqn08vAa9PrgBdPtPAvxquQ/4GNXlj4k7gudaCDf1
VF2uzUXYgZDczOaUj/zth+VWirKo93D5CesKH7A8QoUdd4x+cxqxoNxbw4cNBfTc
eHg4IUiz46aV4oIgTbnmSbs+levDoMT74Q8UmBwl97WQC+EFF5nSiKhYKKDojCIL
4Dr3Y2FaKaieK96Xs7O169WeED2CLi6hf4TfeTKiOdHS3tj7WEIvVDRZbJlIGIc4
Zpqv+5vQgtJPun73mbvvJur5kX6QBMXz6r1BakkQuEsAMAjgrI1M5rIxCwKRz863
smYEQWfObhuNWd90jqykfIEM07fvogMVssJslhBonKs=
`protect END_PROTECTED
