`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCTsWKp2BgQaxUBLj7/lICv5vvUHVvYTg5/kWdLejjev
Cl46WRHkdLtoT2Nhb83i3IrtqsebANyiw3K62ZzZqh8syL4/FgFBHxYxI5SDrW5L
sACC0dznzDicYgeuXq8xScweGuKFXBngVP57Xa4zw70IP5+Ojx4Jdz19Ed6qv5iN
xPsvCmZOyeMpQuTSNKWWwQ==
`protect END_PROTECTED
