`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM+qygZskkyVRkKdN8qHeKcYUT0YVkDYssLiS0ltbh1m
lH5XhPHBvQRqtNsoegkWGp1YUBRZ9yrpjmC/pueex7xExhx6UVSarc6J9ZXg2S2A
FkcaUD+lWnc30sWIcAG0BkLoY+98282JbXigIyiLbipzCMpbjvOcGRluyWX5AT5V
KiRSyMBDaYfkXRBJlnIwN9NkgQbbTfquBNrSUlGn+lCyOl3xYMPuQj4yuK+o60GM
CY8e+1MPqKZW1Ih2s+kCdveYJIrvUKDKnPSAvFGIrLdGN7YSnHV2F4uI5oKvyJ8Z
GQywPsjD9lliMYKIz1p4mw==
`protect END_PROTECTED
