`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
7RWERbz/SCu29vx1yp3KRKl3Jfs/UNumapSJSIFc25X0YU6pxSyKgD319HG2Q2YW
TGgn/74hrtqBvMusHoTETfhik285yWcgysk7PQun9N59nVFA0MplZcWS9UCUKrSJ
XfdPImHeLtr14wIvGcyxuPPUCO381yEPTSCFWCDkxGNBEptKgltHTWWnQYczYbu/
`protect END_PROTECTED
