`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
zp2SaK/+ayEJntKe4llSJkb4gnbchqdHtgvSPyidsdB554CB2n5zZMW4RRC7+hmv
pxv6+Gq1aeM3FyS/ThoLDe+Iz23EA629yzSAxF9ErC2D71gk0TRB0zYAtgLzSnky
VYAtWl/7y1D9f1cbd2fUP3f0aHU5a5AhixMyM7vmtmZGIjaF/K5I6c9LG3C1qqdN
6UCYDh4VIUW8qNqg/WPoSoHkJ83yEQbLE2k1TiqDpmZKD7fq8yT0BWZiJUsoXHTL
a5/heuh6WNzRc/GEDIFQ6Gr5Jmxoa5trWC57Sgso9L66yaLBmTn37XWQyLvK839v
VsUKWNC7V3k5yaCsRvhvO/aZNVCs06ZhEAqtEfhF9rg=
`protect END_PROTECTED
