`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveITzGy2xhSxgZSjebiCZQshFYXizmZ6GqcdnhQ8tcD4I
SjnF5z49Fr648Em7+GU2pFSMBBh5FimUCIXUNdm24D7PR/sIzYmAAQ7kYybwIX2t
x7RJKZ+gl6RqfePsskliG4NK9BV/gK4xgUmgEy1IoQjpN7i43q8FMBqEYXHWXaCK
`protect END_PROTECTED
