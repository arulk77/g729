`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHYwffwpWEbelO4HQXgYhSyDG8EbhY+yfZD2rjmdpH3r
gRK4iluHCjOzE3S2TYBpTnnV5E6Bld9kVRb0e1VJ8CGAprob6O7q0MmAuSUzzzNL
nmenxV9JaZdJk2ELtF0nhxE7ZWMHw5KMa+vloHB+Q2BI3/JXI9VskCjHtnOO7mZv
F9vLteTq8eRxfqrXXQAuVh2EL9kzEwwov7iXOvB/pUapk3UTNaT3SO1kgmOb+qhD
sWONOcfj2lvtPTKi2DvzwXbh9YbpwNDJvdncWrRdROGXIXMF/tEl+87bzSAsnF3L
VXsJ3r/fF6t9w8gO1nOHbdFgBAZlJZiC3kCHvfBTye6vJjUYpSFvhHfDUglrJHX9
kGfOIPRY6aXuK5F/i9boF/My9r4/EQJOfomSZufFKPHVo3awIAMhn820WuWxjbPJ
J0YJGIOpm7uKHsXAlYcP0uCSV+YPejsvxKB5rRyydcrMttg/Y2s6ynFLYYDJZt6A
OGWl97FAn8u839rvzjSLfgITt1oReyl6AEnhbomXVAS/Qa4gd9Acbf13PSlfsaXj
2OY6f7H8PU62EljEUbnGknuba8twOXOfjaLaS9O9Ld0S3qE5kmRZPESNvrxpTgMs
C+K84OnRtgKC6sYUZHJM+kRgXiVPZY4rtkJIl2Etg4tfVs3yHd9xZb0fzof8wTyz
SIAnyWD6KgyHBgVsg2gUbJvzEbKwz6ml/ehSXTK9Vnw1Z0O1J1mHykQrMULDkKOc
Qbn88W2yjeQovON6BFN66ntKZ/aocIzJq3M/omeiLrPd8B6aXGJEZgcscbRinqnX
riNmbKyUVkVMzf2lL6V6CgNPFLv1IfENmB+65dLBoqU4Z8N/9qrxtlZWGpOiyhl3
LMxdZuVSXsuyqc9ePl/hbfmnpxh/HIopk/QsshLlUbc=
`protect END_PROTECTED
