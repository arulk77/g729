`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
waJG2il4PrbpZZvqKHCsM7oySsouNKPStPWlQFxWRphYr3yPL8g+ouAEC4RgqOjv
rcZnGPASZYW4i29OGbTJL2zzcSxIxexoJfsRerts45zQxRU44o1I7GbRkFSMikrJ
8TBVwSZaWMRIp3IMA+Am8hHNaPyzW0/rq0JXiBLa2QfHAgNsDq48s9n5hTo1njRB
r83UxdXxj127VlUFy4Hzt7yTJrmwqGMymqRXckmqbO0y0lL4Pj4lnz2nZuQpy/Yi
TaN5btXWPJs/efYcsBRIzfRd1Y/0zoUuwcIhxJAovuM=
`protect END_PROTECTED
