`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
K2QT2l11f7Ht2wI8IJY0Rl0NJnmhNIaxl15csQfG6QwrzUwYXsCmQF6bwwZtxRQA
MWjDeDPiSd3TyPUiSZaQRYmsxlPauflgoM94vS+VIxGHA8zvPbIUBrzx7wKSFugJ
V5rev/QdH3Y8YnElorBaZsGotd2lyOKNocvJs2HOYTcdidmjcEt6sM+uJiYsmZzd
BQ2qj8mSObfkcrUJNdKa+pmiZIalQROilmVHKiONgqXHuCqxW8F7B5TA/QYkSqFc
26vOX94arGq8l9QaPpcXb33ttWuACOKJRkf7A5witZfPyCGC6NRaT7ayk6r4Yp7c
fht+uXUndco+vVAebPmwxSyXfjT9Sb+XIEL23DFQEx3eLQcyzPdAGZkRebWHqAF8
r89ttvjgG4Jsb987F09maGpFF4qdtGqM+mDrtonby3HZCZmvqZ8HEHfVz8fMj1Jq
3EeDfaxTHkjk8JJMinJdQTRdZMBAIbB4Mx1gRzGugTLcpu/q3UX7D2vN9oJa05UJ
vXIa8o8G7vwc3PwG9IcK8l8k6DJXrW1xHHFScaexa0SyCeoAk2SysuBUCXKR/r36
PQu4epdbTQEVJ65YWLRTJw67vC+J5954sNLojnon3DtRTPGgxlAfdc05bW3dMpew
`protect END_PROTECTED
