`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4w0NhAvtVltlTNxBqKe/hTZyITjoud/LclvpQrblWSWu
9JadSTeEcFja8+7vYxLRc7MTm8jf7++LiS50FMRecH7FhDlbzqp0QvPOoV0PGwEX
P2DuXDU6DwmETI5Tv9zdLKU4MmxEzdo9tjFdQPGxoOj3OUyr8URBXkbAXHTYLDu+
vRKJ8i1sBeEEOIXl0kL4d2eVOVpazEG7roO9Wb3bgWavobsdpxSa1TAwtKhB7IYQ
FE9KSJkGlTkEo7KeZlUIjInhsl2Mn46zJJBOXooOxnyZpMUMgiB1O/+i2+MEJNSI
/BuIctJV+GZcyXFAZ0aqlA==
`protect END_PROTECTED
