`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Mrb9mb6P/W4vjTruQh1/crtu8UCVWj3+ZWzFVoxzzXGdi9lXhPShjosB1v0NKybW
uin/narweepkowfOPrNqH++kUyJnpm3hvEm6BPgyuXNmCSvTlRW4BowztvbfJZSH
LmTQhoeCytwVz4PUEm9RdSg44Jz40EpwkgW8JXhD1OdHHVs/1VmWY7OIdKlwftzn
jBfQm6wqw9e2MzzfpvSVe6QV6/8EUmN/94EOW8nJenkcX5skQL23/eIpShR7niAa
MJxfVqRpv475Iq6sjfwjBd18IIDd0yQ9FnblqoXvwmY=
`protect END_PROTECTED
