`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48UmFlyEkYcUZ42aWjdWsk3xe/x7pJZbrCauAMJtkuXt
C95Fl4ykChz0Y1aVH9iJkpbKWggySN1KX8tmyPD/aqmdY26mic6jdHuEmSZiQ5iW
AlSmXmkTdLDaTS7qWs09sG+mWXOR9Hd2+zwD9bd1mZ/tLbqEfgZplX+jUHIELZ4M
GogGEnLgSqmrMEwFowdyEnNx3UGkvOGK4AWD9NzU5hvgxRdgzkQierU/wNcvljP0
NLfRcMlyytk06Li+tdYrxwqaacj4WLLliInaFttevts=
`protect END_PROTECTED
