`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHWRgQMjjFdZ3hsZaY4hGkEuuSNABmtuIV4ehmxitiGX
XI7N7Wc0RlIchTIUFu445wpChcC9D/fXfqFV6GiSqZMP1kw1ogkTGIJhJDm17EQi
ELPqS+PvBV1123MQ1ZwunkOW/KRirxx187b2/zsqgJQLcDjXUvaaI09hU7h2NTve
8Z+JrPIXEZGqp4j57HMyzg==
`protect END_PROTECTED
