`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C/etkn6OWovS1ja2eWImINqV4BU2kz3sC3FKmNQudZ92
ul3hXRCrWy5gLXBZmhcYBUadD6NWLrmCnKfeJV13B4rL5QoSyFq0vZ1KG3sJoG24
wQ1mUGt+dUAV3gsGojc6M6SUWbwDI8xeuFWUbopdLwUvCnCoFiXJXWgQc8C9ANxM
0hEa8JNgjvI8GZHvXF1fa2cUC2vrm1CgvyBy7oQYgkkksCgjPiNypXnvF8wcOaap
hZpthV7ZCW8/P3JmGpKtKK1vj9Fx2S21dNTGnFif3KB9+PVZGC2b2xY3dPvaSeXK
sYwMw6Iza3IuxYoOB8TFtH+MEvYh/6Qz+qJplzFU2GH/PWDcBHRCLxW8JEkCEN+1
ufL5lUUCW5ExbvLCGrobrDEbAcKpHtM8kpmhAgCawSMx4Krvq0KKRDZuPPyPQHfZ
T89FHRqwuek0o/kiB9b3ApkEzZmnj8xqYLBpekGMvxlzkVd/KJE+y1GZle2X8BA7
lQJXpc9/STBCNw4BURxfnlptzcYlvk3TL2c6izq+akk=
`protect END_PROTECTED
