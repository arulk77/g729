`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aQ5hzSd8rkASjMaYSoD+E1G4WCu8FJLvbcWvSfjyftx8
MLC7kgjJVY85R6fbL9ago7KPoKl6zURI1THWJol6XXe6FHjl6y9rOI+o5AD7ecrI
LsXp5kBlWdIyDuCXIV7ghOP3+tXV6WhrQSCgZXzsTcZ/jSie/85ysCT/TffQgPbF
R2O5b6QIDKkk9aSL/CnFGJY215REApF5OXYVHOLMcok1rjFQXn8q9JV048uafmUp
XHUCootY1ox4bMm/a5unCTTXMSGR8xD1mzlOesoV1FbGn+i2rxPVoxiERMEsgxz2
gYT7TuMcvNlmVI93i1JaQ9sQLa+ri0/6FHQVcj8nWkJ0LWaxlQHoMpD+3bLovKeO
J9uossSUHGhhhBbegIAfmTDYd1ZCe5G36rsMVbbVVvLuhppOn5tHO/O/s3YgsxlI
nBBqM6KUGP2QJMt0YlEL9HOUL4edrC5q46ssJ/IOxAWJqOPyNGyemNlaCK2lxU1a
cmKKVQ81bM2+/AmwZvzyDavi6s+mLOqKXeAwNrpl24IXwJrspxQ8QzfiV9DYUWCJ
oNnf7mg8iuterBPHSN5RQOGrTU5AXD3IMH52IVsFiyqMAIkjZz3EitsQCN3994hy
nuEBQ6YGcXRTm6dUElbLqkNj5qGnCg1zcugrhDtwDeATLeE5EfhClZNE+xBgQaAh
EHncm1lDdxgigiGnX/KeheNHFjwJ5YSaPuBX4F9gYXh7wNJRjGStxCEv3JVG8C72
K0Ies5946aev03lkIfydksT34T7d3kVn3ADZ/PYqCo6TPWSZK2euNhxbg7W1AvoO
uwnN7MCkLbcd+zM+k7PMwPg6Wo8znZWmqK7wpbs9xUsinvj+y3/XS88Ju1cPjXGL
GPhupq8Aa4Ybpr8tSHgd4AJ7RjptO0E7kUPGch1nfTfBxZxDntWDkpwyqoXGXrhZ
DY4m397OH5v5rF0QCZNyd+9Rg69D+eYfXfmvRrjhiV55fzg0lgEKr7rJEOUhjsyV
CGbSISJnHFb9WNDYNhZD2Px/DkwhljJanoFALL/rBufqPlKyXon8roV+1eBAq4sM
+J1IoVKt0wyodreGJ4b4729oqd3/XYrET3PJMme31JockeezoN+a4LZEKo8wZBLV
DxQX3pnV8iAZQSmTbECgDRIb9kEZ/aTfZJtOj8IMWwYoFYiKu4adVFEGmDm4VnzN
5/x6/CPiqMOrvY3vSPR216yeP2ZVWcURaUg1q1RnwcU1aNmOsL6Xr8VYs7sxZxHh
MUAPg4neuaHLA/A0HyzI7xOOS98+YWrphwKv7h9nDez6yXlKtxAtKPwnJBD/1Mt3
hBP0MXQ0AcaWeka2AVEAg0k5X8JD8qBp7fa+bBlaNkQgu4LKq/p74D50jw8VmRwp
mfmBj7RrBfm4qwB/QdKAnjcQQFpPcmMMz6GJ/95f7Zf0ooYWWAecdZihNOuaRctJ
n2FztT9fZ6Gyaoxwuw0OChX97mkU5BFSdyNCkBBfldjV8jxBKxb00v2sMR7izNh2
CjjbSBLMBg03GwY4jO4qND0kNfa8wZgJnQEFrmHQdPHbjx3YuCPcmWhDUQsnmcWI
fnCH5Kmiiw2EyfJX/CmU2pznb3lkRSQdCgjau4q6suJK93o4uAkkMOTkfXE1So9R
lwiIOdyV2T0Nkm99SX7CEWTKwehs1zW4gO7LNJXrlst96eN9uBFGcza3/fHdyAxG
nFAXUFc4BC1Q0MHeeub9hsdeFskH89gIK6mXNwSvoPFWxJ2I6fQJ4yFN7AdydqAX
4auwP8lpvDe85jdEs3EHUf99VKoRlqIsPq8FuZ4JWtTt+sg92VtjtPeOta9KlTgM
HLzbC02mUt8F6CCZD6zvb9t1dblSp6uOkGD+wjKIWaKP8ghEd0GDTu3yRaa56stL
iajS5fRN58NpPvf0pAEdjzOb6VsOCbP7DQ/zWoxf5qWsiX0FNLWPaWzkntR79HoL
Y8jbpqQtiV74uvgN+DsySD2nLB6f0EUjTYnTf87HT1JXan3O6Gej3aQ7r5Bg4pT5
yKK0FUxFYKmfrBVIqaM64YwEaPdHh/6CDvfbYcCEHn4UtTItk856FmyfakjJzBc5
LzxND4Ul87FxwIsENK0ch7tKrguCv1KPkc1OrGMpQEKRx/IaB6l9xuLXAvehazVW
dU0iz5XA3erDei0rtQvfIrat88NC9RvBm+OzPD/aAcdbsbMgG+m8KsQAZ4xE055H
6tT88namMm/HiC7lXwVdSFQyp0kS8hErxRKusXitb4B7J07WzNhw04420WIF6HoU
1BSZrdmOwej3pyx4L4/Xlhq3sgx7WU24cZ6VLuAj6knuwpEU2hTibTr4PNNfzrGw
9ZNOjs4yu/hFTX/mqAvuoiwR+s1SrgqAq6EK+Mta09NZSqstEUIbrjm2YQGRLp5C
IiBepbQMhEWFJjLSu6u8Vu8ESg0xbsRnP1uc1inrnRembvXb3qyivxRnGG8aKeUq
P1jNzfstbmq/omx+7612zHEC3vKMkdWGPh9boirHPvlB2fYKWyLdOfnuWSOqK0J1
rV9Gjx3ZjDoaZ5ToKeZTh1Xz541j914UtqEO+9tDgfsauLz4ZwvKR/VdEo83KMHi
1rClGRriE+49NHN6mRuroNyLLhfTHk1jkFgSehUOgcAApj7iZ1IS5MnYmCzp6sBp
2pPEwSb+uxrs6YrO7TayO4VASQ1A1ujHUAqSd66RyujMpIbmD1IjbIZEY8bsJgty
WkzhdM2SYffXb2IQ02r6FvxwdI1ZylHABSEnJQnStmll8Fb1KlLqEfPsO6SizBKz
4erFNKzHiTjdsVm/pAyv0BtEkeF4pzOIEJ+lvOWJVcLC4N+32YR5xlOsymkVAkz0
4fOtPTM759AmphII5TbyCxAck5B/3M8S4vRZIyJoweihhpobZmxjzzxW6u5VDOeE
NPa0Ew2QpZrIUAvNzr/w4TCd/MC9zo8N85rR7vQFM9igyV/03l9MRHCSjKJzTxMN
MGHQEno0LvNu0T/Lm/Jw8hC8EZbU9rhp0tmTtymxhIw4WNaZ9pn7HW4kfAnwKz3x
x/K+ShooYoYjJqIolp6PDSuyTONtdjcmSl6VyQReWjwYSte/lLZpmpv0BgY1Q6hn
1CQXAGU4wlZsfT9dWqzK65GZa+gopepTp0AKFIUxx9Js0+msfBTnayTQneZOWHye
C9PvDHwP5XMMvls+oLNt+aAoo2xi9WflIOamQ9A0WfgYJ3ZROGBBsYyIfhOq9oxB
K/CXsqsMd+MbsK1TAz2YDwzKmP9Q55GQbGd+AiFQCknQ6rHQO/1qCEln8VsBUS/0
TY6/XqW+xfqrQcDsoZJhdnw5L/dMFsMxKy+8OHa0pVaD/govfER/4JfJhrvjvbdk
xO1NA6IFFXkid3RTtl4+U4NFbYWapGf1bnkiA2EmYjQ67FaKedhriEqxFDU/exGf
wZraeAh/TAoX6CQve0SLFrsOymTP5hKBn/YqD7FIYx4SxImlEoEwDt367pp/nvDz
0Z+HN8jwyOosxgKvbzwJfp8Rf1oO/eTa7G/Pj9s27l+YjnNO921Ah1aeX1gLUn6f
51pfmxscv8QoxWtD7bDu1LPN1u6DA0R4OK9aUm4JD4YARCIXvn6uuLdqzK0sde8i
SMkDH7o8TbzAheLzQ3wF0sfOEm7J4CyGuYfr/OzxeHAAFGKmOqNN9PcQp6YBYvWj
fULZzVOR2NZzR1wlOdUNwPRKqsLWv674/dcW8h1T02wXo3Uj0oyn3EwGHB3KA6Zx
R5OImi3yGRdDPuZnQwwGHsYacJE46cQ0SEWU5uBY/Et/5KSKfckowqPwRzU9Zx1E
7GBrhraiSFtApie/lfb0FtO1wp1hVI0lHqImYPseVc+609WirHfBHNoD1JyuCR9C
FnwZTXt/zbMRzvuJBKzpzwz8ORMSNGQdWRqD9/PZeaO72pFdz9CG+0JZXJBR/A6s
3x2aOEW0QdonB0b1iL1A7HkZYq2tWm7g42JOyrImHldtmKt5h62J09IB+Er544gm
SOwPE8ZetopXKBjYL7GIujq6d8DAh2SH83pbXUdrA6E5D6GewsExNhr5GZNOZQpR
QjChdm800tC65NZxIFcBQ/z5J0Gb2IGo7yMqjg+bE3ztt8xxfJkFZRXapADP39JU
SNbNhTLXlCsb8Wb22vl8wb7brw6nfHJw7kEnORNkFDwlzDGEcLeyIPJa6aToMcl9
FzBVZcl+UHXWEi11nNgcU0o2sTNTrulkXQ5fq9itHfqa3YUXmne3sEvxmShy+ivU
sHMYA00xEN/XsRT8Dh38BCtmKRcELwPf4xP6O9OU5oIIhwoZ2clCF+E5mXycqdn2
c/EhfolfGzAiKIRXboUuf9XrjOcGnRBddP6S5IR2PC0/sX3WbPYO1fe9WGvRTtea
W38x6wKyDLeRb0rq0VWdR6mOB9Kp8tY7r7T+ug3ZXDqdmIIfcRJi0t1rbB/uB26K
plqud3sXKgnoY30bXCJffcckeRdGtVXUnkE++Ia8n3quefI/UKpeZMTvuOtHDNOe
+wjByEc8o+SM/BRmp4VDvOFiCv68xQIQXxn/zU+WEoMLrxHaV41YFeF781bGayjI
onEaQr38DlZo4XGik8vbQWZTJqUiu53BlHuFMbt+Cu7Uf9wYoHNOjLJDO4ovyMMv
GVSUZlwiN61d4nzcrqZhX6bAmWTicr8lxDymWOy9qM53UqqDRIi6Jiy9bxV0nvrg
TxL/+FiUBR+DxTxaWhYAFPc+Yt8s9GjkKlLA1XrIOnT9V5Mnh1gz/TWS4L4046IX
l+BBZakIE1mLoknHuoK2T6cDTAKKcqsLrQXduyjkEltn6C/LHMwI+bGzHKFEaXbc
WuMGFkXakjpP06JvV1oVABb0buiQ4LO4q8xwBt/fRp6pxV7KlnCxWeWCxjFqjOzl
eVIQCgkvLpd1OBWTG772aHfVMJT+qKx+2MRHvdh9kTuedDv3wcCSShSRht88ucFm
0P693vpE9wJNP04u3Aq24zgLZ2rvdHJprEMakr2ID99uYmXizMeSCtqi7S5+banf
I1mkHDH0FfJZFyZ4k4IMiDIAPcpu/KE8++9aJSf7cR17w0mME6rXs4LBtBjk7j7a
DAf7rygLxnAv7g695rPQV+hJtVEZVvd5UjkPRazdl6vb7jZGoy+E5JVhLCIESrNa
K92CYL4+j9IpxZZE2XB1KW8vEZTFjbIReJU8jE+3Hpb3JLO7DWX15YQxf9XZu8WD
h9HsZMHc8raQaWu4Yy8eNRKmCrc0EsNan+WvaYmcZghNr84HNkji13MgPiLZqTdd
bFbgKvATzigTUWZvokIz4Uv65KusNShN47kJeXFe04uEVmGZRxKeviWuxF0cm4O1
CumXWG5cPpvziu955l+VEYRjIbKOy51ciX2AHLYvzzQzlN/q0MaKOwlS5RZAwCxX
SXybrwrufTLcNALOSj0UkMeavsQOZJVJWRbwMr7lbzOiQVqy9LcGsBch67RdQ2hy
gzToaqFK2+EYTlJ54dS4nNNApjvQ7ZMFS2WC7T6WZOe6nZXWVVGg5GvVKAbW/yCR
reMObenDyXM8j6S5/riQKwwpL7N7kxbaS8DdLCoyNjlb5egK/Q9JXURkHBA0MOKj
ApNTRU0CChPGWKsZV7hfz5bhBW+c/lrLihtBQF7DqjL2FgY1+Ie1accR5L/Y8sy+
ROeyXadmNxzF49yb4+0PIhGFKuq1uIL6qlGIYitjc0zCeF99Kql6XKZ0Cazg7V5c
1TtgPK5p4N7P+V1jmD6sc4a51NSct9ZKyPZH7PpNulHf60lvi4PsnF4FLLL0e8gm
81lIA8sB96VgcQOGStqFGb26kIVacr3M7WCO68S7z+hQGg8G3TwFXxJ3gPHFKiiZ
S9lhwm9ptbOTlt+55CTwUDbK4MAfv2SnEs0bmWsGtSEHxFX32kIIPsh0Hv52CTmW
nmxtJysysgEU9oafhjw8w4FgBDoDGLQGVGwbPdHrVIFczS4+V+JAXLJxsEbvG+n7
bSE5Sj/5+omOJ+NtPKFw99Ju66mA7rTrtSb6p1En07gmJ/IO8FosepJEx1GIzXs2
MJMnZ77e14GOkSRHhA35k5gOZuTsu4LWWSkxiduZ/zET8ra7bQyj35oM8t9+uBFr
OYIT3yjZCFQTarsdWfecIJy9isK/h0JhWppSUkusD3WEqnppPULghy3lcBgNP92M
XdboILdtyjvxmCus968z1YESV7p3ai8P/qz6i1KMUw6jBGddJVx0IsYGRt2m50Cm
aynJFNFhy7gg3pfKqX6Bw+POvgnXKnl0cE+2qugQUBdb9mK4fupu576O1JXx3NUE
HPVpmcR7USoKl2QW7aQrGL5EFkz/b48nn2dEdT0bVLQV0ruflwQWeESsKy70v3eb
EgHgJl3FqqwpeIN/q9we0vsfypP0MnMfCzRk5sff9frjZ8VRu0FQQUOMoiTrDxlE
bX9gH1roAFiXGJ6ob5O0+aawFx0cDvO7U+JnQeLA2ir9MQjasmWUCBS6Y6UXMoZT
5kHPBXhs8UQDgTzsS9STYdjPjaKWVffMVcMPSw5LC2VJilmDvR3LdsO4D6E05ePC
P01OVIyS8e+y59EWy+Hp+IlrlNvnGP1xzqxjpYsDj1bLXA4OMLQTbCf+JQVGuonZ
h0bNWEvzv1dbdfxgzZvq8V0uyLy/xsdX+EHPtuTKKHf5iOkZlG9fpG0sWHMWgle3
rShkFET5kuf8CzGatz3fccJ/dWcrFNWoqTxadv1JmTWmeKiDQngsYAV1jY+UfSr6
wEX89dKH/nOlhknJARTxnTgUYhVp724mYCvH7MJ2nWAIW/rTZPhTRao1hG3tyrqD
Mmz+feZn9SCe6RrtzaxwXev6wPaEPmnOecTYBKpRvTX6bUIkVnE4YAiZptq4CASY
Dh6Lwyd96SwzpPPGyU04HlFobGCMTMbcpE2mGFKehND7T0YhsHMqFlIBWvjOEBta
0PlQyXGs1KieS1Tg+VrbbmJ9lum6KizSS4NOa5xci45cI/DFku2sjl4eHeeQaMfP
rvko+5RWvYTSzsnWeCwKEMNKZDGT/FUQNkTuCrDQ50skH8VOmqlXyyvPikI7O4fk
rKD8VqBN0+bX8qCGyDPpKOOoh522HfCHK5AmnHk3fQOvJ3lbMZGJTL3xStYp2QVs
yCj2KK2j1QvUNGKcZmvE4fN7zRd8MsNISZXLKBaNBuqVTIYI13AmVN9s8qWpNG5l
G9GyyVDcjM5m08bbgF9oN2rUoKkhX8OOXn9eo7jEDeTz1RKxHTQxSIykN7hHy4Ie
JvZwYLHGs/m00Yp1is1BDQ5bLM15JFlytGnL3TEn9wRzad9QL3Kgnc2yMFrwV+4z
GVPGRsrVGBOVVTN0MZne9J+3LWUuQKByHAinZdSxM0DbEM9TKA3hrx8QBA0+iJlm
P+QnsfkE8rHqWoPte3W9AWZXS5nsWIb+Z2sA91HHYrMcRDNbnJHMLl1a3/a62U4K
4VtdbfSfFIK1JNI9IrxuRhyqJk7pDLgNMpngcT5iw9n6at101AriHmTmv1wDl3Z6
xzs52Iokp2v6iC2AXejSAVBfNcVAF/ZwwXwT1rRtjmGBJYypSSZ8ye+fm1aqbKKv
Nhg6lZjHdJ+8CELS5gCK29Vsrn3q4kDjNDOQLKuVwq26agmHa/wWi5Ju3570Ehtz
50uZEUV4vkBdEHc26Rh0gihX+6DDwbbDvLicWtrWK7E3YTkzolE23+5EOqhzGPGI
a0dK76p8yNhUF4V9Sv5N3I0VpaO0op7kgSMxpwhSL/jGDi78ZEoWTbODeigP4VNS
H5CVizReDmdTPuBNHa4JrkLmKsDPcfe1rqAJXnYhFIxau/GjZTnexvjf8ljbqSom
q9XD/U+1GC9/0tDtevQSnT4X6yVjUCnDbXK4Xr3zPNK5yZXutitCw8WL1h/6PtLK
YNjd4HtPC0FwHRpIpeh4IBSaX+ZaxdX/z4aFt3zW59usxwWdC+aeDEnUReQupXpH
75+vfdRv0ZCaG9fDkJaIcdgPhZW4lwOhS4an/ZlM2ebAmOEc0jh9ybozfZmAzbiu
VxSwgb/OgbMAGfdXh0zMNv7Zb+zA+tHYuo3DjwC8iR937bN1b0BiiaoCtw34LV+W
wjomecGezlJPrwRXaK4JzfxcWeTUzN9RLX/7aR/F+AxoUVzzblWVrPaebqSzzsFh
3dbCqk9a//kC5Ef06qwG5sIvnQ1F36sanr0CpthEwkX5uUZle4vCcDTkO6ioZIwE
OUZ7Gvm5+XRuN+nPXq9m1/Qe0dygNbLFXFqGJXHrCicm467V6QcQGVCWSKb+PQPc
F8qQO1TCJ0uhkAaX43FU2YKKLKEjYgVSj67Jz9lDyxQtvvL3kqTKpCzk341VclA0
iXZOY0T1wiAVItLZL3NDwF5xbUpe6WhGENsAAhtqXL+WoItIzVod8z+E0w2WJ3Pe
h0RHGrEg1+JLswk+dzfWFI+eKy4C7b4u6ECOl1V8vfxBa+HtugNtqXddkY87nND3
hrgerssIE7ipSwfG5WtpaPVFJroyMkDOtbR61JcQhRJ7B8TBR6NvmEyIqgvLmmtT
QrLtI7YSHWidwtvMhBzenYWUbPw5SCBN9J++Rl66C7jRYIAr6QoT+F23u9k3oPDb
ltOospwDi9HdF7yy03uQi2WJK0EXPfMEC4ulvR3Oc1vqpotcyxV6eaYIlvKreFaL
fFACnuJ4ZS/frHyA1LxYMIYTQSQTCimQuaOqDJVqsQG4MenFEYduBAXdevGzZMZF
CMD1s+LN/boN8LeNgsXUtvbXPt/b8KJf1vl/ZwMP3jugX6T3jCEqg+bf4fH8AMbS
1A03vDKiOzHlQS1UbMAGKNOu3Zi4Q/87SlgMbJ2x4gEFuX8tIl8aqgedGza2RHZO
5ArLNHOi6Pe9hQWGT7cLfbd1gW6VJVndbWi0HsZzyfeJcBSRmMKP8Bk9qAujBcH0
JrTQtcFq4Xk/OJ2UK+Ppgw2D/kDaWKgoT5rAracgoZV2WYuHtBAYwgacMU0c8lRd
iCXZySHORfuM/2lJ2SKAPHiRotWDghDj2JOAfd0sWjS5yx/tk/IHJu1Q52srjHM2
Q8JWsdEbPcWIMlk6H3eqsqansaT9fksEZmbP+NSJW7URdWVHubxQDCgn11G06BMj
6GD/1I70Nc6JMoeMzwIpy2RjeNVuqaHv8R1QcXSU0TntiMhuGoI0h0PWRw9hzJ3y
i9T9CbnaMPCIno5MQ+iCU3np5JbUb4wAeQ/ZwYqLh7thdzFkPvdebO7msOvCYPHx
pwRHKB5VMlVQCB0r58XDZMt/EfsM48FtFGQFUgVemK+sOKV1a5gdB5XzrSaPipsF
1oMEAxEDR82lFDmlAqEZOV075hVLN5TI1HKPNgmRllNTXn52OZDTQXbGwf1ZJJgu
crYmzT7hR8eDLtTSRSQBONXTo4iCEOO15UW8SX7gt1v5CNO4jp5K7YpwybaRMuKM
WrQqIxO6+A0+TkY87twnMRxBqNvT6OP8TrY2Yz9njuZafrEKWUwQqYs9eslSXJ6j
fGPdBaa9aBfeRZik3Uu5tq++1Ab0iniQUfAEzNOiQfOzI3Ya3DMBfWk41LQbhOSw
iGrk5H5IyzFm8HVS2TDsQsDI7TdWr5tCSkFVBhF9bKfx3zfooQmXVGV7NYgqS5F9
g37HSGfeKhNL+SCfT+91EkhPViUOz10AhWvdSPZvp+Sk0ZD5oS0Z9AqX8lSaDA3S
5TRhELJ2qSumrxVaofrG9K/AMaiCGX453N7dEhDCrBHJTOhLEjXfjN8oOEqGfBsd
BKOCOtN5s/4K/hlkBsxeAO9wKN6poYSqEODWM1C7Ai9kTybYIoGcQISPgRcxiQDo
5UHNQrzQIKEYyLK/QYkmzmTHOXxqD1V4yN12SJTdXFTWA74iL0NxASCFSF66qp93
VWRENOOsa2Gj/L8lizSHMs5Qmc7gtHGiJ9aKv46zwB2264wZhJCGt4ijf1ZcHeeK
MgMb8stCVk9lPf4mtBkJYYtmV+iLvNNswN+Mkrdt78oqOWwDtRu05E0rarhOHDak
aDAOQt6eNUQH7XJvAp3ZhrD+GftzmDpTTyfrDsdAnOR6d8+j2LWL8GQAXRniQP9a
UPKHjULQ3r+8A06BxMIISIbplbX7Og3G07W3E6x+GurNWK2wMzdtlXSlJTLpZy5R
jR2Duy9i26zxgFRyLKqmMLHGALbFK/GPJhsdvk1qHuxvj9gtrR6c2UL3LIUgDZIZ
ujJOXGoT2iQmKvH1V3A1sHbr4yDqK95bm8UZHmDuRsz2c4axyCkf+w88eYw2FROz
9JywAhLLEL/Vyq8KPWy/Zem/RgyNRD+W8pxZbiQHFYdu7bfpU2kZuJ44rC3LDK9q
D3t1HCT7g9HyvQYPN70fVKRIZyWfIajKGxIGQjjBiQG7DDInXcEj3qaogvGiYpzu
HmWRsccAGBmvu/ma/nyv2G0wG+Nob2lzwtb6JxWCJB+XJBl8VFBlr1Gu16xZbsMw
x0IBxqtN4MfALZdxrkMtWCk9QybDkN6/KR/0cyU3x3mveigOl3/vs1ARk0vY6A6b
9bXIXMSai0Xc9jQ10TYUnBLELfc4qQkPb4OOTPBXW/A0dG+ySyAOcJDejyVNE1ul
DbqPOnblpAtt9e+kx2pfBiKJbijkFg/rwP06/8DkVqsY+Yhsv3Ny4a1h+pGat8IE
ho/P+dYMqC3N5fIEpTw7aJ6o42Eeb5g4TrXRj2A0JTX/UCHJreJUPqNRWT0D3Mja
qi2iqqeL/dXriz833utSlGT11kR9qeFHM79NJLLzrF4SXpmwvSI9qtwRcEYtly65
MI5ceoDjC8Vd0L9Ak6gmUEutLRN38U0f4Qw5JEt7ssk/6GwjJ7PfMXXIS8/4pIFK
IlSZSdkpOFNuz8i+pCTAbXVj3CCLkx8wMdVm1KmS0PCjG/Vjwt+MJ8JT0v69ctHQ
y6aoyiUxrY2O4lh6NoHjJInx6BYPKZyFn/Mj4WaDZFaZfSUwUIhNaWrwumRtR+Q/
g+xTeJSaMQKSALLb+SJ3tiB7Mb/82jAGZwepLS5p8uuzu8TniBisnnMjYuzJnkFg
fNz5GeWEsgVTWAbRNcPceUC064IApZZhfzcP4HSOMiBBemQtscpnGkRWJWFX+G11
FlBNwUpWGGNoD0MOzJ4KYHWjMeUia0VDimQPL5LC6dZ6wFO2jbzAP+szZ/LHQF4A
uv9eTrwVjcN74O5j8t2gqpD3klii5XztZyNn9B+DzXTU0hF1Ev1rmBYVHSp4KpYI
+GCvtp1pNVIhnmrEmfm0GHPFu7Shd17nT6AQJ8gzdpbY4Tkc4Qs3DGj9qjmzBnGM
xSzofrXb5knRszRmcaVuEts1IF3pEupAxZM7yw3iwJm56P39fFI7SZ2kKo6EO+Qw
1vvdUYeG8+zDAVN4xwTpVfJGJKKkQc7zMqjmUKbrpHtFs+jrC2FIx4mzdSr+Sl43
wFHVPIseG3FaC1jBWVqDmQSDPYbFRPrqe3/bLbVP+NdRANgR81xxCdAvWJ5bgRJH
GgFKvnBuBEgCnVlwl9NXFTKY+APsXgwVGbBKdVFTN32c14J13HSsGbc8hPNQTuaw
DUAS8Di/HBX6hWn/HB/xLoD2HbakCYr+76n1pbhffi1AVUZEkk3COBovce2O2eaY
CKS0na9FW7aQBPyTtPxhRCcmX7mnIOvnZXLCZIxQZ3B1oUpJQwWhBPnk2tMH/BL1
S1xtv84FtBm+FDXwEmZ6MnqHx8yQ5RVYiLdr8795YRwulrhPI/qAu55YQxnaaWvg
LSpuL0/Ots6BJPxVozkrjxVzzS5doEUdXKoz6nvRTHtikeNTAldJD72O49JvEN90
KP50rSvdoYgUqT+1Pr1tbhouVG3YEj1S2smUhVcSAyg6rX2ZwqIlnLcjUNfgh89W
N1bCP/46D4zsS/h2id2pRNJmHJTMU+RjTZHY1gefLpjeAP7E8mO0BM+PDl5Pu2NQ
rHMg2pMWadqpkcBTkmNLF5PPjfyXssDeUzZRBN7LSqhtsXEJ5oppmjtZ5ZDI/Eo0
bQje1Z2lI5bh/jYKyo1eqosIsBczz0v+cMIge3FgeMfYuPf6MB/VpaFqt8oLYt/3
mT/jsBksRLgdXcU0HQSozKx9SdG2sErM5vhcLn5CI1hu0Gtpp8rO4bUKsduphAOt
u7gU5CG7xIG4rXaoFqQoB+h2ggVlUmTI/KGkRRmWyby+0rxCa9ZVzFO0Iw5DDVVl
ozles6443bUfpWqIJ7pi8OUzYaf6y7Kc7TEFUQ01R6EZUfu7k2G7hxuXXnb9gWkQ
rTnyz7XQwdWeS3w9GamETapsi+KU5wGKUa76lhACqtRKdK8/vWNMDUQXtzU6bJF7
ax9jdJcZB+lx3A/CMQFhaKVYggxTAGx5ZyZNKaCdjAk52pX+qdpVPI9I5193b4EV
aPp4cpZ73THSXVyYQZ1GmlRBvISnPT/RFUrs3/JJzAN1FmP+PiKgCT8CyJ90ZTYR
4qddTN/BPIMFoHtlX9k07xOmFmAjHt6+SOqCTo8ad1U7zMMNOlK0FT970dOLjAs7
7Lo4r8J/4lH+sn7OWR6++GcQBPsSZ8Gxnh1XkZD1CvOyXTDJeKbI04cgyrh9J5jB
FEeuhiROvR94pE4tvAFgNaj62r0wba3vUVrWUoTtT/HmCt+1rXiSIKdOqVgR6sRO
YCTrThD+q42M/rAITSzbL6QQbTUsoG69UGJy0qibbDOoLRQLK9wBBIcJlCRVM7xv
G31E4Xkv6re19366uyf5mzvVJNRv+/qAyxFO2cA1tGYZrrzx7MpkdFz0GiJpIsOo
CKNbnfazDfTt0PRb2HVY9MWYmWFaPEpo84QyRH6YEeo0ruD1gkLNsODVf/GrQlKu
8x5NRM94Mzxcgqf5AkP0MDxO+XtjHJVw6NtEk7OifECcSbKh6b/kskAvdlC9o+od
8iOn7htmkm95coNUfETzcQ4z6PfWHPFqsfO73VKYEhXFBx9M+aQm+aT/nMAnnom7
g7hVrli4xZ2REUceKvLIVcfMMkZw92VFQJJxzDY6aoiVgv2tSUFPGx9BL+Oxr9cf
xoAUaOT2FL7l/GvKn2fswgPGh3RBquB+zp/UvBWI5VnUAdUvpBB+aUjKvkLdEP5r
OlhpY7mvQpm23Huv46n2jD8sS8D4es8CTWMrd/iT63zgy7PArwfDDyFPq3/GNeIr
03NYRbEXovn9cuNjBtuX/KBzkz/3W9dUXzJN65SaSET+zd+VxB/5mDIK8OYVekgR
F4X9eiaIjhHva2ZPrRwHW2Dp7T1i8DW+oAGgxdtBRFLkvgmvKiCA/8Ta0CM8Ay9K
nn1pGH6jAcQ92nfNKA6Qv+s2cmr5crv4b56qKqeQExxjji1mzeX08gl9reYxZWdt
CRjyitDszz6BwCQbWUVyrYrYACgLWGqMFSy9TvhJodTQYDFRE93pYJt/1dXBnIrZ
alwxn80jcWzvnyodwzXw3xAoiwklyBJVy3+xI/hoZYVxgBaigkOjM5eHKl+ECL66
R6K+hJYbPXjRm8BV6ly98V5RKqPWM4QVeY7omVzN4g7hsArF/c6pZ4R1CA6X1vhJ
6OqyAMjnpeXAolA3oRTe6dUMqjw0RhBr0LBnxOiA6r7ieYTCX0/hB7NXfxImbPU4
K7A70KbKeQD5JNZDxzvTB1w2YHmpuh6tfUaohupT1+LB9vM9j/0fhmAz/08YDc1R
Gv/RSM/WtdVsPNkZtWp6nE/3QmLqVN29M+WnAljg0jjebIPPRWRUJLc3dn5ZjeFl
c6fw5tdtF8I2Ums+jpk9VJEPH16Ch9ISAt5Ql6a3+O876kX6IsgPKUtryMlGe/Ij
+9kP18GhNdqvqbj/o9aVWQKD2Ds4s4Cad1+rwEGLPUFizjVVaKXxBVgB8Jd4K9hh
e+OOHq3K7nqw4xmGgox5anmp1rkqM4KLBOOezoXjmqSRckB0cM4YobA7JyulMMWN
mZjZsmihrzpRixHg4PFQYMxOQc5B6l88GXyyZ0IPyMDmLnefQ7RaWsgm8dI/TjgQ
3bqNlUcrHEe6iVp9SumBGKvth8G3epvnxSPG1Xym9e6oLGc5zeaJwyPjmtvz5XGx
SajHpSROpM35zZr6l7xFixeZZp15vqZkBVEhXAO3SbWvWMacsprK2HuhVykBKm7X
/9CpAxrht9aTlMA1tZoKPyJ2YtK8wGs+uVAqlCj33QFuF54yuUTFOlrvpZ9snY2B
B04WJjpKABthBvZxMvmV7sFGdb28isHqvTtqvNPDDgsBYymQkGTl+uWHRJJaIzx0
5WSZ+Eb/8LZtXxoP+i8afifcY7dgZuGFBv796QZdLX+l/q5cUQ33L4a4oCD0o7rZ
xc2nPefu3Io/oOOt5KnufHf9Mgoxv13/7153YeUrNc0QusRGwvFXf92oTqI4E4if
KC0sEqpRf+GNioQjiTNG7eezTgcBHfGZWxOUan1W2AgNsAtSyqKRk9u5yNgx7fGD
FAymNTQeMDkdJux7vT/MGbjhdd4cY0Y6BUK8pxq2oslwGbvzaBvXeVBnAYt57Rv6
ZTWBk6uHecCVSi7zvy0VODOIM0tA1GI7E3Dc0Cjka6ni9FOkNkU6S0YxwXDgC8Ru
Mh1RQUy4bIARz8UaO2FcTJLJrBsrGOPJewg/idBnQSn9zwk61e2IusCxI7pSe0Iy
MidJz7HP/NFK7NIXVnvotO7NcS426cPUlZr/UboWBwwu0p7iL8iGefUkZm5YusWk
1Ab2J0jlLSc8Cd49P2+/QdTwFQ/wbXkc142zZKMg+9kpT/zdo1JF+mNkhEOd+/Mx
aZn7BE4+6tjeOfQ+mxKSaLn6B4xeM113jqnAihJo4YYgfyLxaPKeK2nE71syzf23
eMQ/bQrkoSINvboQWCTdzbux8B24JybJDzVwZnAe86DcD2KepzfwXqe3Wqwy54Ge
InW1khW9VaFsKw00mMqyUuDi8PrLliyRWoAA1sr1EuJAKdzyxreO+VeeqaFu4GNT
ufAQV1nBVf5C+4IHHWJZytBRgmFxSr7A+QNltzoPM6pjmjXpFWP+5wUhU82Ti+de
q7lesJQRI7eyO7m9Dyi6EpcTmGXuXvb9h6IjXOgX064FQqQuWwavrQCwKJ91XPS2
ofrufpvmNjssqqIaCkMPZQiZ+E6uctnyh+JLlKiKgpL03f4eJC0Jwhk40X2JdRBx
ae6dVb34jR9z/Q+C/Hs9AdpvAvIdmT2FO8ZXcbwZlCVZD86uQXHL0XntEOGHZA48
UTTsJO3XV9xuVJSijd6d3Bh/12WEYPD+gJIERiVpV4/jp2MlbfkrZe3N/XO7bIIf
5jF2Ouoiml3OSNdiShwziFd0z/5gOdi9MejoOso+t2l1Hysqi4MX0awa5gsd1W0y
V5D9P/imDRhsSYAM4MFOc2XnQt5QQYExJq10C3qKlHlehgwzgKIvIop2iUFDHPSA
101IWVdjDEWIeKwpS43jsgkJzMs1JaRUB8O3DFK7XmGqZddq3a37rezZJA2LLby+
7TFICAC55P9h1Fkje1vgrOZ8we6yvJ6T4zrghDqC1vEItxjlaiLzO/9NU/kDqldn
iZuFqAiYkExcgN2GyZaf1g0We7s9RhY3RE+QqiYbTZNNF6mdt/RjtQe/GTXqWnVQ
lljX8919Jlmw8CF7ST1joUkc7JxblBN4dC4vMYJn9AtdeeS4jI7p9wbQM/TcCGsn
jMrpuZEKmvBosgD0YU/Y5RcUvZIdvf3+5WFnljcjXspL4NeRUd84sXHu46xnBQHo
xMAIWIek63bo59Jv1ezXfTprxb5IkNBLZl+L6/tOFXK9YLzzO2+QS5w3Azfmc2ae
tN1AdrXbApBAC40N7vgrVo+4PwZh3m6yi9YReQzA8iIQ3uUtPNwjtEQwnvTOoBKv
WIKuimlg8DmIdueOtyAAQCD7lBQlrwa7Ir2DqIZIRifZcerw075ZYXrs9vQEjSzR
0RMBFEZRJLJ9YzUUTttqFsGkMnM4pOl/Bcc7j6JfnN/O/aclKn7HyrZf1DnGBo3R
1rBNFqVsob2l6vtNvRIVEIw5bTaTmC0RuSBxCktGFLd/Xa2CEtoALCO/HRDc19Ky
SJvcX36+P73x9pyKuBeCCpnwrvMkKeH5mIwwUwaaphCHpNPFkWETDv7Uur5SCFU+
0N1gFXzpBF5Dwr0XojG4tKQNIZ+TgVJMMTYq/G340HV2VkvW/oX0l95f3R2aVKfD
yO3md7opRWEUIRo8La61N1bTJEbo0KA+IMEkrO8V8wixXOdZKRFi84r34WMRIFIY
nBKMM9GGCp0yzWlHStGgAIbKrIHlHcpsTZKOZaoScjqPHsaBi1Fmuq6PM06w1jq2
ayCEj7wLOBdqvvjfWWatcGmIYEQC+z8mKeqDmISzXIRlc1bLsFA5dQ31c/SEfA1D
p1UHWpc9vGLosKnXPOD6IK4LIcDJpfH2U2oCC3RT7xniB0EymC2yK4HSqrQ2dmfp
/h3Ehj7UGihYgat080B58RdF2GwiliOfHIDd5BqN2syxSkzLMgZy3etlFmA00Zvt
OKK4oy6vXa2OxEz4d1Rcs6x34wTGQyCtKhYMWQoUx46YUQPmmGptp9tyGjrpkkkT
/BtpWpwcwea9+uqw16n3Vg/V3+OafSiUHrEz6PZ4ij4xZ7K4yr4Q1GeLLUDwIym+
Qk0qO/d+1j7b/hD9ak2YcnT0caza3T0z9ivpl4YLFms0MuKtvDm8EXxGG3JB2fgM
+xzD3Fz9u5jj/7wuTX6jKESo1poIWjIygnEpRKvAv9tIA/qpdb5AeO6bOXLWJDKo
2VwfJ1EaJm5s1Z24DUo2DFrn5Vn/yfjXIHs/5XXT2sEMDdIkU+zzBKZBbe4NsD7J
IF76JPXlQZ5yeoILK0x6yzt9RjUsFKgMp8XYsl5Eli7hoYzTRxXvf5h6IrDb/1Ut
JSSGL46VxZajktJy6Ga4hg0vKnKoK/gupLx3BSD/EKDYx5UGk147+S5DtLFbvRYC
dYovELjoSnYZxcMxyQWm5yIrTy2XEcdUBQiGr1G2TGfo1YmQOwUKe9SFWjomLu9A
/7s9g+0sbT72zZxfiMlbNe9k7vosOXynGy260JwjeZSU7WmgJf5uD25XSN+YBoim
w86VjLyibQh1h4VZjNm8C/niLY3IfQ4Jf09YgvCWmhsKQxpLFAbzAe025Dwg9Tw2
yRUTltQwOOtEi9NbhBadY/+9RtUBvCR4w82bOQeMIpKwMuNaaBD0RMgKah/WNnNx
7wP395KYMnLSJdIRYRoHrs+MGQLdllG4S3EWk9/FUxXZNm1QOLZWUm8F5bzISH0r
qzV6P/OI7U+cM/oooDP0eQgnNsbR2oiz5ZsphNKjgMrEXdUfw8eGqSmvZCIQalVa
wwonqSPyr5QS2ONPUVfTOs149u8GYRjUsXxThxnBGUHWi8MkBvrdvEvaopNbXCf7
37qPhhu8+RirvRrlYHxmpmjC4ZvT/y5uawyRmVvKpWFviaxASYtV1Ota3egzb6P2
+8/YMmB0+nqM9u3S+hI6qE/XFyCerJ+vx9F2NgKUewy3Nf7UsXnCFJxnBrVI41Ja
+6d9DOisvvYWDx2R5lo6v41vi2bm7RtXVJED8CWKtIZr7eKkr81z8PzhDAK4Dhw9
ue4iO51v7QcOaO3Uijj+DvvsUAEHq/6/X5lXgHltHCuiYQJlm7XJDmvTbCIKoMjc
68mCjijLFmNuc2dKIK/IcKiQfZ4ZByxr4VOr24LNBFgtyu+TG7Kh+zcVf0rYXuw4
TF/4udhDylZv4plhlNTycszQZ4ppDBzIpumz4UBX+I3UkNrZYrxJG8bVg9HIZK4R
g0D+NwDyOmuhfYVGOhf5v8ljhkW9zyK+wKO6JmGsbeftkWkjEASS9UulODh3JQMl
njHeoLJd08IxXGcrnp4k4Oq5RBs1HGuVvZKiYaXytPCKMuFBzovGafOBRTaXOqwU
QSBnBPPFuBmvY5e67npcWxPdAI4oBKp2Diymc/OY7F+GwwJA+A3wdJXAXWWJ6dMI
CP9/aNh8i2gwZmN3wE0E5uuINivW4bUJQ1OcEs6KG2tPL7QdXsFXqPixECpRN2qi
Ll0zhIao70rzGUDWtIhc0cTxl1MVJftPebe3FFdmqO8mZ6a/jWWrc1t7W3SxGRgk
DRjONtsXezaymLeVgWY+YsosAouNCpOkO4aN/FlELQiDYeZJbWiSidws+0uQqX4j
bIae2FhimLtmWqQ3fm5El5G/HI7DpPjEOUEFYknA+eqv47kSBQxQHB7isyNPvc78
OjI2ju5j6Sujicf1t5wSqAtGSWLZ69H/kA1HXMNWgik9ZkaDAF51dcLZAiRjY5DI
Jj1Hg52oWiiLs7rdsom6i71V+a2qwjgrNyAUF/2VjQEpUQcVf8wGlh70wfGC3RcT
xXExQfYzaVSPlx0BlT1qZycD1qUv6B9rMwY+WfyJMNyr9g+8aj3mRo1mxNkn2//A
UhA6g0Lv/lwAdLL/40wMeEQYSwE479rSqfA5UpfJnN0JI77oleT1RzQRmYdzeckS
4inqRnrcpmEE4OAJ2qIJSa0LQWrCJ++CudCLrRHhMAY4QMO8JfkElRKDw0XDJqkG
m/MgYgKqBj8tQL7u8qOFYgzldyE5F2VBoOirLXr7cPbddpPdgbK/cHPs/uKrFmMu
vTL7J/H8jWD2H8Z4SJo6kqlFUmerYUDf7Ub1zDch4NLxMTnC/JGq6A+sLTl7Fbor
2zN+wd8aL6pt54u1Egb0+cyk+fw1HKe544iesLgWrwoWeK39o7EAzCKXmS27SzX+
ETHFnXtIcq2jjFMQl2lLdP61nwSlFud+Jr1YHaEcPdpvrR3c1I+4NqffDcAcwl+S
8MkJXTKrHWR38GxpzewRMv4hXV7O07AB3OT87vm69IB2PTccM4g8EbrOs9aGtBV4
YtgXzUht00r+a7+OIyQqNYixClR8cTraI4mK1jROTQfumCe+8BofJrD5YsvYaK2C
x+ImeLMFKKl44x5zzmaM3Srs50pIYoD1ukD7E2hLybUUU7HTZrDfu9pCD4ob0V8l
iWZdLMTg1rWQ2wv0/4Ft1mgRyKsK9b5GBxaSItyVu+y8rfTj/Bl18hsuDb6yTubd
jwLOyuxefnpDCX9er2dPclpOd9gBD34yWARTl/EjRPb42Y2liiTQyY4cpQfq1f7y
6cFB/nJd66ZzEsp5dsRcrlRTpWp94Yv/gWYVLyoy+InwTEsouV0ZJpu8DZB+vzk1
XdUh9qYPc2rEW3B4ybL+x3Ng9fvB3PoBuQOXkZZfFxziXCNjE8JJm8u07G2HaWO6
qhNEW980Wq3qwEw6l0KtAEWN5ID5ur6y+EKBu+OJ9IWJHN3cxcGk7eXZZNq9jzI5
DIIEAsdloOWXTkIpJ/B9NuFiJSW77hP+dqA5hmFlvCCfM+i3KBhWDRgEuepuynfT
spL/gWO+xUEnEtooEdXtYXYBSBhYm7LYWUMMx3KGPLUyAR4uwW2xGloi0XUIfdft
zMc69kqlt5OcJn22Ig6ppqyP0cKogVMTwp7ziSQEhhuPlZzv21VQXaUoXhKC98fB
LO9HO5mOCHsoaiW+trcqFX6RH7m4hFfDR57l44ICHBz5Drl+ei+92Uc6EikJzYXl
UXlpk5F7rIPcfw/wv2N/iv2U0f82YktetzbSFFdjDo3Px6wqmZT84b8BkFAOhKtq
5apwRpl0en+Ln7S99GRHkxUG1z5QejJtfgmUHeffJvMczIpvCQpC2jLNE8Jfq7z2
/TVQm56cFXY8Y47FgFtNsSyC+//4iCmYa+BfhdJA9X9C2rs9CYbJfpO42qhmthlU
m1CTouMUbnZo5SijZyM9wd2U++v0kSz7pfodYG4PP43jJnSGhmOQj+JJ3gOhBvbQ
ClV7cnwryIHCb+GuAz4OisDau6EN7NY36WB7YGsim6d8/xb2yWTv6ZwYNe4OJRJT
/NSiw4OzuVNHyBaU3sUoaqe8Rr1iTM5gwSW1NNPiVgsWdNkqkv6+EI/mE4BbEc8e
Or/YUPap+luTVypeplKofHWwpRiyqhODsmDlPwNzX1/5Y7ZOuELu8KatJg64EtbM
aoBnUcJSe0V4EoE7kkfdrBOiJTZn5ptZmqunBo22eIxnkbCj9PSE6DYmqZesDxm2
frzRdfpLZSZbHWaLpf5yZzz14C2H05cYXTvDCokr/WXGjNym+ybwj8U6OIWbQ8UR
ISDrMgIJ1I0QqT5yfwh2sk0gUydyj9zqn/pjCRrh+AbjtTxAcQYOc8lcMOBoNXVA
Jp0oTSwESM0pmt2nrOtWzschQEuq8awMYVXIEBHbyoE7u+ld7QlKcm9ctxb/FeWt
mHfl7nriB4nrAOzKCb92HokFA6Yl1cFe7kSzVTNEZHiZVq4xaClg025ZShXgQaIP
qsSRIRWjgiDSNb/JjgUGjoqCrWMmMBuuRdhaUT/JdjuXN8TLPoScGAIVsbYGBb3K
DO51lJp3ptqJBPRLxgXTegtr8n5/uBBf72Fj0MsJaBzU8m0kC54FsZOZETR1UOk2
DrFSMP5LQ8xyxH+I9EAqVf8jhRHEQqHmlnd2cE1hKq/yOwacoF3Yf6E7VHKkUaQo
oQzQcsIfEs9keSGBcuxZIDp53kWFuoLAmbdTFBLH2UkcWoKy2cjtEN24XsVETKx5
TRA8t5OlkjUGvjBsGmiUincIJFkMUSXvF3aAZ2Pp6JPihPnU3As3oFZTv/J41SP3
Yh92SbLGUNyaqUVfE3hd+pIwoD5fJkVLGM7IsmwP6l/iMu/aQm75AW0z4r3OpE9u
/uboyZAd1amXVMouAjeT7LzHf+0AyE5guEupxQ4mxozoWHn0RqFYRuy4cCVcz/B+
YTsuIspRIRyz6//pnKlUA+HFeuQdz40gZs7AEcsv0gGXqZiWjRCBR3zSswnG0s39
MgAx9xTlVoVx/npQ78nMvwVvKhYfU18R3ol4NvF7UwQsKX2q4Ho/aFzt/geKviJE
Nz3SCEsqhmkObyRYRoQq63Kc4KuFEycMBEgRuR7amS1MZ5d24cUkb6C7HVpUxshe
u4oJM/FLCgm8Hg1Rh4m2R8bVq1WDpZ+UqdXu03AkYYF7enmRRDbwVebSHGQutcH3
xXwiw49wV9Rs9iouZr9KpvgHu9aonlxNveRkZweUUZ1k/ELxfpyAkRQNjPRXbn2k
NQz3o+3bTHUova0ktADLyl17v44t8lSxOYfZX/U7BtKm34yTjSk3CIZW87Dr4O1X
0Gabdr5Pm/7Dg64yYh89D5vOWTVgO9atFA5MNsvzu/FyLyGYYW9n3yjqvTqRsb4/
RBVTQ3SNA5tboJ3AuUnEavhwbKe4AlIOKQkPBFtN7iPdZS0OQr35vztC1b/9pWyN
3X5ERNqPCzrvk7YmSLmOTOpRLNLjn4hpawRUGAkRlj9kcrvKwTs9ieZuS03O9Wck
VZwDQS0EOwPpgCyMoKOPmAsNQz34fS9n5oCw18fjt9xXSUZSqh90CAt2Tsy3+xib
kb+VBpWC/XJAD1+IC+rIBua6fGxNtdRRnAKlO5ezU151Lp1s6w5B9r1KAht1fuZJ
VKMkKaJBEzNqf1pyTrF08jgeIHWXvhXEHYKJbWMpiuoTyjtJWjV2SBiXBc2v2yWN
Yq+wPw+KqAr8s8dtPN6nkL1GnCqJMgHQhAgXpI6h2vDwWbUYKWYmbXO66OxqKYXZ
0PDXvacgA5hL46z7fi5HlHpMXkkTn33wl+D107yZY84FF7Re6SMTfSYK2bl9csDa
9IQei0ufRpsiIsWSXOkmae2xxfDTPMvzH+jvD5PV13CO9LpogKUK2f+34ECVyB9W
M7ajrmsjKWNAiOn/VYcx8Vv8h1n3vnBxRxRyxU2zXivyqfA4xAiwdTSw3oV4t9O0
K8az+Scfs36Xw+WzDVpuzutGBocSdidORdBUcrlbIEn3YuM4YjmdTTCrYCj44H/3
0yLx+Oe6fsBxUcDwQvCEWbVfF++by0CIEalcQ7B14rv0obOTUiAbNOf7GEoV6R1p
pLlXrUyywWH41SbbcJOIZlsuwMSAnuPp1bmcLI+6OUNQKD/LaPh22rTOx8QwlSll
MSI1ejqmqdsH2GA2N7H/m0vfTLMYbpNU9Eskt2DAv+fFtfsxOMgu+Xe60DbCAqhl
/JEH1vA/mCIYe5m2BDHheXbAC70Jq/1hZIAN35e4Sq6hsXA8pOyxeiNUSDp0vHNu
PQv617zJLrneebO+quXQ0hoN3Sj5fZv3Mj1C20rndE6xK/SX/2ZLrftqdZkdTBfv
icjiCYciqNfaJSwW/g+eUd/3laTvsBSx29ZsLx8dvSWL6dKQPboLTQ64HeLfVddU
mYURrOiPgRwqLi4EtJj3VhFLHP8XP+33rjaG4Z++4VNapYK5i/gMryoigBd7rFLM
KSQUtbiE4qqvyXGgYEzLVUOC7bXaUVFCS/imzXzsFsK6xtaae5c99gPtW+HHLmwb
`protect END_PROTECTED
