`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aZTgHUHEH/QwrEXMCokkCFEx+wmx2hPR4fh5s/6tmsLF
f4GpiIcdigeiumwURE/mOnftLEXWV1oHUgpVsTjkUKC6oGCZ+9Gqk0ZHt9NPw3A0
Foo84l9L5dV/qJNr7iHzNzC8T1nFUgMxeC4XQZsb4oWLwtLdufkRb5RnQ4U+o+04
h96NVlt5nzhyHNNLPrOL2cbE4tu46j/TRuXdjzakYVdc5MGF+RNOhcH/iJlKflG6
/MW3wEx/JEw9kmPJD3sTncIX9PGjpFuPpE/F87nNNNgUfH9uOFbeCosnqrbmsGRw
G30Jo6nQfuC+tXn6kUq6a0oZvaUf9C7e03tpzBmjjrjT6Vw5K+JgWwG3A0M5kRRB
GyRrJon37gbfPk/hriPhmW1kO3jcOzv2jEzTXgbaBIRyzYRPvURrMXMxusWxcia1
Mxbv4tac/DKv9RtjOFS3EAVx/1BBgA9djpkPwqGiK7M/L4E4k58buRv9496qyR8l
0MZNCNXkIfj0gtgCvHZxCJoDOj2XDmRagDKTh4jxYVaWwWlMYk5SXVA1BD+A/3wx
jCBiK+b20A1mX/5Fh4xHaZAEagK8pOfYky83WoPtVqjY0jLz6exP7Y/8W9C8Jfoe
dTzO6+61J2skM/zXM99IpdqVglhlP6QJBTSKxYvY7LosH+eWplKIVvBf05zaDzdU
+9jr/NHz+DpkGuBMSv9dKlQFyx6XdpWtOUjNw5m2U/6H3rFLHZWkYtnNpORqxdgN
xVpZUwYmpfW/xg/dxNEug+EKoRPdtSs9I/UtWUcFPq5+M4CjmCuNLQUSZVX4zpK2
SlRoWVMQtwoZd4iTNtHrxFgLmWxmfKxD9siXEbpbziBvBgHYoOG5BRh+jXKnq5wR
05xR15tyUBXj8z0m+yWmOZQAWsVf74pIlVTSS/dbP7aa/GMLIimEsoZxx13YfnIH
Ct4cd7Ieaa0TeQF9qkfyeffjQbE+9JpqJn21cxVYkAPizqTzu6LO3csl6ytQG83n
oVfCPpEdBC0aRQriRnCy971gWq4brTQoSivdcqPD1GZnCsMZkkDAU2U/2slBEtHP
4gtuiUhvjOOpceXVxqz82W+JKO93vTgAi3hQOKEZvw5g9GaBK/qKoOWv+uu6HPXW
XwA0jzIRkaiq99orOGpz7yg5ZmTsL/0v8X6+T3R4PlhxGbbrlzzNSz9UfI/JNsAF
P9Yr8UzVYEh6RwHnsp9P6KrxrH1Qnxdn28bTWxg3bE6UobH1kVMlS0Ip0NB64kjt
B5RzgiRf5nmiQ56rIS3zBdDHMfDmICQiHX/WSOIvvzy+cVpHhzfFVPm6aIxvLs4E
5mUno+34N8khsYGJhJgSQL56+Zy6Ynwj+i7gwqd+LiBx2vKmJUJfyCLxBJfrvIvc
EwuXlqooO7wijAevC3UmlruwSmRwdhI1ZdY4bS7Ey/xjHfxw1fOEnujhWu87vbKy
YmPXXoWwGrLCn9+DXBzFCAGq3i3eq+wKyJR8qvtWy/iNWMMiwHQTvIVp/Dm+/6y1
6vgdy9oPsJYSein7DBSW0Co9dtJM07nH6EbyTPhBiXgaBxUFRTIEHWCW4+dfN7EO
tfnvQJWEhAkBgTdb179BVsUKfg/qUU95TJwFjfB6tUSBUG3Qpt7wo3jNA+pfD47W
o6s4CcEQhLFKrYgMjJDtF/fMfBqb7eqS25OFMcTNGroqDLC8foZgPZRRzQCfws3K
LecAf6mE0qF+dcaEIRyC55HRi1XOEzkQEyU9QsEnLU8ibT4NK9B3rilC08GihbEw
TMy/nqGpyDVnReiP4AqGAAf5/ZjPv1Qkfgx92DaFWwmd6J9SA02+S39PNbfKJgxQ
VvcIWidDmVHD26Lbud6HFzozOpDlgic7LITlwKKhs2/7pszJNnfr4pggrZivvnrb
hEuT90tTUCYAdEFgCMBqNN0132A4KnuTxkmlE+yC+iKQYg8GlC4/yUr5tTccX//i
KAPDFFf5s1/BJ/pIpktS+EALsvhn1yAt2RR0Kbxsw08=
`protect END_PROTECTED
