`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFFnpXvqfCsCiGGoicMkaRGYok1hjVxbTXLY8c8LtAmm
xEjLsn9EsAfgeQ38HW1ps1Rot9VyiyOFYTLsRKD03RMniwulfvsuLtcC8qwuMo2d
ZaSvQ1u4RSjTiCvwGNJ2+PkQne17QlyBgP/QLCX8NhjFgL3cDCLrIiCBreR8Jk36
w31YLSuO7xYCjHsr1+oYUIfyfDNfojwpx9AmWLcQr9KG/ubjRBIWc+Oqlcyb02KT
sSKYViDIQusGGyiKEllxQze13/xQNFl1HgvWbwQAc4yNJ0X7gFY5AyeTj5Eo6Lco
W5qPafvzYeW5g1F5MCfDQzGPwqZZr2mDUmLVvNCiR/qMRbdS9QmsHynsOmLOIIC0
`protect END_PROTECTED
