`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wKkYrFwc2MAcJKqUl8NLWGE4tD7Nfojrl5dI3iAhl4s
lrYPqB97LN1OPXbCCiuvqkRMncZBgwwFM7S0t+qT37Sdzc5t6SaNO9hwE+ym8svP
ZmUNxyezzDI3EVWh2qAbSTFcs+He3CMGTWb6wT+ZBeSqdnMdSVBi8RTRrw5YIG+v
eAJ4GeRUeNRnW7XFZFbDaR7xic6Wm1qFBkhW8LQ4PrHQ7iHTr2v8+JWbBoY4iAGC
IlbSKCQnVZBBDUgqWmHfTeiJks53c/d4A6U6/q57drFFf6l1wIpXHA5ex5rczoc6
YCE1wUldN1ZWfRSwf/yKPrmK8JDVNwcFDFVSWKlRkMdGafZcQtpWhCXOfGcUYUmS
gB+73iuKo0RVnrbIsyY2RS9Sj3WNhB/SUz9sGyK3z4lgXUUPVKqC8vtAFUtgEAPI
0UWDWdqVKI+ij6hsPKYEB332qgtsd85Br+kKEUIcVNYzS1+i1CfvF+mgKc1WUtQK
`protect END_PROTECTED
