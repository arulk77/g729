`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHysfZq3FRDG2fI+94azzrTlPcsI8K3a9m7D7/ErzyBO
fRLTwoz/Vxp7iPgrdomxBg2shiGUGtarlTyy/chIX8/3I8PpPDsAN3QKpf+j2NrX
tNzzTfXguZwtqD/Pf/pooCkvGq0lTUwJmSiU7uAffcFg/8uvTMdSShzzE3aRlZie
vwZ0DRh8yyuYuvI/A9OeK5L2w8tWUzo/4BpEdWJ2bzTyRhZaLybKY9zFJpyE9FOp
beYWl5Mif2JK6CN4t45GWJhcRIN0VFxxsgel8/UbO+71lLOumZPLyC++fHw7yyDr
iVgUA8nCtXkGyj7C8eznHrUwBua0RUZoz/GwfEaXnx2ter4aA/TbzZ+J4FlyosSk
pBWJ9tkvKUl+Mtv8oset5QMe76aVrrPNUoCBlm4uJzN4iri9aPjrOoVD6YCwZWYm
L+WAyXyE7jjJ1b98yLQaIPt6R0naJG6mqkP4WFuUgOycmwf5Aa/46nvWkHyF6iu4
m4iEXblevBzOfd/BsUbCZLdBJ6792Gf7V9Fa1T8Ek3SAAqPg9U9ScHPYqqbRfcC4
`protect END_PROTECTED
