`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAL1y+ijcMxsIwr7tcYyM6AcZ3jrcv2xP/VrAb8ZjthI
lhlti6XUkCoQyhF9ODypBnfZB/y5djz9cwJLmTrn1BpPffjvgFGagWgdVDgsCZCF
VvIyuEZUfWwvUEnebrwkUNDSTsZIkRLTyYNLfUdLgZlezlsR6DZMtiVxCC5GeJTf
ALDdWupmvYV3i/0xV9xt2EeKPYyfYY6QANrhcEiPKHJDTIBi7TX1ZUfTXfoVFsm6
PZIimYXZPSE8GP4jnS/NTGmure4n0LDqDvs+FnFFnaLUho+50UtHEVZFx3mlHNbs
ZUqOAl64ndbEjlkDkFUR6A==
`protect END_PROTECTED
