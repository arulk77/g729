`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Y3mMuYfjZm1dJ35hFMgHu0Yq7uNam4/wzzJmfpQW4gb/H6C+MRPM5K8uTWggYyo7
uReh9ep8aMwWWQuzO8WbGSyXEDR/UQiFXPPdXnsTrRm4RdiuNy4vHWCkX9CcT5nO
J7EjIOdLatO3q6RkPxd354JYfKWzJTtgXH0zhDlBey0NSGX5OUkSeZf0jBHfolfk
aA4Gi6KCP1GegDA9UBDVQekOGfyFO2BtKywaWpL8AiE=
`protect END_PROTECTED
