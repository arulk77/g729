`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveECbt6Qwnqh2KSJeuJeS7TqjcvSwUNzEOaAkvCgWEaR/
sZUQ1gNDXutfcJo59MvV9XxR9VRsUbedZprNZCjZ9maP8BeLVP3j6BOIRKw8vPUY
auYxtNvQYIrQ64iQrudIBnuGMRgMrMrniE5LvutyJJIEJwERUnAZo9RegkFBMP5Z
nGP9llQ7ouHcHqBvPvs4btSO7d5Jj9NtnxzvkgpBC81Sa3u+CsY1VVdzwTTYgKnm
`protect END_PROTECTED
