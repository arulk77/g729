`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAiu85UFRmgWwVAAb2PHFC24oZIS7BSWfz8RMndVermH
EYBtokZTOtI89UrTmC0/S1xAhJgFutV64msyMRN/rmvLtjaONw3QFnyAqJTmD4OZ
pAzyQkyFSauiCL+qU+cK16x+tSUt5tM4a38d/AwDvfO+X+ZA49nDAqgC9C/+BeMX
Nmpu3Xt+Ih29Y5bL7KTDc5zKref2qfpFOTv+5u2TxLYvSRCnOgLF3GhGpyWn3BUK
`protect END_PROTECTED
