`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN0UrRN/OF/ycOQJZfVpuJOK0G0H3NIEoJB60RAchAX4h
EoTl6Rv16qiLFrEDim/CH0Ek8hmcL6pgh7CVdanYENh4b3MBy4egNtvRPCaFP371
zD5qZ4QYpqrZoZJWfwU+UwzJBQcypx/Y0VdyPUIUz//fOY8UDit+RSHjeDkN6+uz
iajxc5DmBsqRAndMt1dlmNRFpwSBkDyGwg7LWBhaR4w43k2DYxlTrzsweJFYWkol
pjpiPACSWr6VqssrM/nuqn6aCK5cROPnxQUMlHyeKCczsseEymoBIOlUQfJBqReY
0i4O4X0q+vvcFx+yBfk4T8ggmfJG/HdYkzyKFsVF7j8MixWXz2y0vvyVcSJdjpCQ
zZi4Mee6nUffZrwWgLxF/SBEq1AwrVn9kG5C7PfSDmSuatmVBVMlRLAoQxdQQqmw
xHIGmFMfyoScUOxOCioShJxQzM2tPbsWkXVrN4jPwQHbI8njQWBmFVsdETHyLBzM
KD1BcyELo3IDGe62WZuQjTXszIHE1z+U9J4TppeGVEVOSywDpUgSaVkedbqLy+Fv
DnmOwRqxN1pFk76M+Yt8CgoG56PHSL+Cr+DRjTJxcyf8q8CpUyZ78yE8wiqncihP
m/dRzoPKDLG5PKZfd0D9rczzzcap1Q73gEpLrpt5hvGi5za7YU3JBVOkkpFddV+/
SLDwurvdm722McNNQY58+Ck+HSTZqAcFFnFuLpYsLlQ/F6/MYVPwsJvSU8AIe4BV
1Yf7I5AYEgYmEml00zVKPrZal0OjcdRjg1IGoHySovw6TpyGkFenPKis9ZZcGYOJ
7irh4GZ0Eo+GJXR4Us91CX7x3UUCI+CGqzg//NuQEJUSF9HlIgw3pmejlVBj611e
4hWK5xRYCL+i+tR8Spo2/NOXT60CbPTqf3Bihv/1Q/Lzw83SjWrJ/Sy92K1Fx7gk
eHbAAZA6TgA4niaP9TqmS0kiw1TJmUDpOl8ATF6Q58KXcYsJmb+wHREFrrtDJ3TC
N+aumRG2acp+QMnxhmjJ7JIKlLy+Wwi1PPbCTNcIMo0ZIxMz5bLMIxZHKtryoRC0
KBfKAiOZ7k5DASrM7MbQAYDzLfkIRP5FbI8XWYq2iNdqngGUb9eJ8b9oCO3d3D9q
Q6+Ff46PHnZ+3eD/bOSrmCTFe2Vy/U7t7ltYu9QFldh8m7jtUthwl8i/FPNw5YjQ
fDn+YjVNOh8za3J6XlJIC1ujrTtsjzZ9L4TNyHpxnJsDVcSM+YoabeKCGNpjXHr5
sgUXuVfNL5GOCTwjkV8XNt5tCB0G/5DIHa6hZpz0vtcjww5yBBKfib0nFH4YzzrH
yb1aWtdhTEpmkGbSIq9VS4eQT+uvvBD35bAIx4tuhrUEFuO+hqItSGorKzIWJ7Mu
ukdphiv0i9vtBXQQzSc1MftJ5vXkQaQBc/VkA647q4zLmtDBQvYRZJta1vQdNBSX
i+VJSHH/jQuq+5erthc9++2WYrak9CrOmasuF2brVe31F8lmwtQMpmxdAC5P+Jqk
an/KBn0B7wegUAeYfF7c1IgfKwjdIV4VtQSaDWlGkf/gPVIqkbxo8pqi3QN4O8iC
nhnX0i3ju75M68ecKkCGuwbBVToJTHm6jIQYubfDA9bVTjKOkEiiDzJ8XLlMu84C
9U1R2G01fRiaS6gawoPZXIkB6gvHKNH1GAlIIJo3Z4nIQ3qLugGvEBktXcwfCtDb
gc1ergazJxF0YZfc3w7mCORbNvkoKq6nSnt1YLVYdViShX+f+hYRH+6GrQmYWWvD
mVZyVyAq7MexoLVgXwFTznuVXXQtmIvR6HgFgPxTbNmk1d8KZ2buYP0PTg/DqH51
rIl3f792TXUKmFzOKyWTRUtfLyL1DO1fNb940PPU8A5uMAoLZhtcyws9enmoUXbN
H1e882yhnIr3raOABqnmWeERWx7+i1mLbX6vbPBdVgzjMoUKWy2PBFwCuGUoOhOA
/R8idqHUkOhA8c52B3CsvkGJQQqsXhb5AT69lVSOlt2n6qXiUcaN8fQ8g+yrp+rn
DvuR6B2rP+SMpjusU9pC+T+cDo1lnzn4ELzyLv24BciQfOoa5ubzx/FVGX30Ag0J
q/mK7hFxeqMaPouD0M0M2CJDE3EHmhU0+Z9auSNf0pGKv2c2h+MdMKEFtygJlyYF
6TKuzhB5TKH+w4QMG956DChESQS9OIcK3f8leHv4Hv9fJqHQgdBtPOCMvCA0Vnpy
mOq5mmpcCQqni6+FwyEyWV6tVWEWlVFss/PMU3Yu8nDhDjBEbrBEVPyin5O/43w3
LOhrp+Tt/IY9+Cr5SvCcNnCYA7JHjEJMirYXEdut0zKwJsE9VqmjRy1MFUC2OBpE
MbZ5hcraN9C1hDXJh4Bh6db+erJvQRGJfl/6zpjHZUJkGIxZB+TYSJC4QWp2vM6e
DjDjYgaGEqJn7JUO8/jqC0IXOtjt4dtN3fi5eJ7/UgSF+4/53PDXWvq1cJ7eupLY
amN2hl7K+UCpiNY2nBmuU/RSGiZt6EaTuZ9dVf0Nj6aWrTfunEH/Of0x/GWjzyI8
9h4gy7UVPbierAd4JoOmcbh1e8cJSwddkXIhCJ1xLY9FFD1vMR6S9pfnNaisgnV6
gGpRJ+G8atN4XhpIroTe383spvzUrv1Pt1T/lpPPQBxpFfDCqZklT1NXyJfLSeO8
ZCpeOn2m+aEr0zENFwlaGNSui0fWjekvyPUrR8MQApMqivjtB4ZUq5FXR4eBJIpV
S7bg4dcj7Mycsd28G6nM21m6Pn5hH82ESE6qZ5T1nfIrh+V01kj/evHMWsyMK/N8
f3IUWyN9M3mljIXuKMsW6p3eiN88ORZJ0ecbotBpCei0qrOVusTn05SAJVCOtq+y
tTPhHHKe7tZAc92fOyDjbXSASdn9u1CYQ3s6mip5mJKC0RTiABHfH07/+NWmi7Ed
EH9Q+kRnHAITijNIGCjJGk9m3ypKSX6WF6YnOI2MYx5DJY3yeJE7M1ieOgOWdNUD
F6125OuuasPv58IKCO4tzPwTB6ROFldtf+3y2jTq6oiYKQXsT6YepsQCp4ndXO3W
8+Gdv1qCSh87EbGjkjwi9F+lqDgCcA1CHt5D4MuHz2NNXmsFOBH0P+H2/g8BIYzR
UhPjzJ1LfFfjoaaz1Q04CdpAMnspITD/zh9kvTRcMD1GekCQB6PI1az3TZVfSlnd
rwWuFxjjvF2VpOuHkcpgS7YLqOKj/26NLWDXh0L3PtoJOJzNybQ25TwD2+TtTGGD
jFmAn51q55nijMp1Rokcf/o52fpie2i9FBCIa15WGdy7yMqTBvZf+wZh6qToA84t
JNmogK9a+5bQTsPoZxhZD6QbgprvkmbmPWUp1v0oQd12++3m/cyhu6li0ZymnFap
CxjSy+LFPA/n9x1v9QOo32xnzjSaGu1lktF91TeI5nZbbQjO+BjJ1jTd1vUlriMp
KTt6xnGkxzsycnVtW88l4Ur7G+8nlQcav3l8hAIRgMfyLXYE4JdpG4kgoLsWkrJj
05O9bVglF0ZZpI+eds2H7Gli31uDdkNP/fSLEQIqoFb2rQh3Lhfe+esVdlhKchgZ
gI7F/MBi4TVR5m3vOVAyZmBEIK4oJAwD/BOCvZvTdTKJ/rR9+1YgYu74VVWyfwV0
UZ+taHLlZZIUoWUy6OWyB2sjbVcB3Zu8+Dqu/SYRKXKVcH7sh3cwEKXH/uf/3njH
OyiYqBIZ+HQgAk82lxSQxed8VrlPobxMihPKIGkaJ0ppFYwhBYtTPyA7kMfrbY4c
0XgsiCbJH1JlxBzNQRL6XzLicO8geHnkJGgLhpIDQxrifJ1kZ/KSUbc/E8pg93DG
l+C5lItaC9AHcFMB/VG+txyAcpHjhj11bFRa0j/Lo3IPH2dlfWU2L+hR8oaWvcEo
TaRWKwD2cVDkn2lQYLb/lE6Du4ujWpproDB2da0ODUxKDNXwyBdiEnYLzxSqVbVW
eQ95UE6vf7dPg8a1APqVQAS20o8E6nw1o+hj7+i6DSsLcQfOClRJNM2pUa0EiMdi
DHFFmWtvb5aIrvCMu89NMWLbYkxdGiksQ0D7enf4DzEDfuEvggsnfa/35HSQHaA/
y6rIrVgh3Bv29/n5jQIrElBV4qGvZ3ZVeUBf3ZqQbXbtxGB8ZWIlgZgnyP/MW2JG
kneoTfEiQDLZGkAx1MlVC+WSDsc5c26y+ivGoazEz2OSSReItsaKWp15ukXdHzM6
rrHPRy+Uff1DQGJ1mksrWPKxTiGS+Fooj4H5cuFoj0TKs2DmgjJ84RjYR090GKIS
SSo1H65RvAzVResi5E+AJNNCwR48i/mvy0bo+YoKMKgvMb+koBmdXteIpAzO9FAy
3QUbNuy2M0YnLiQdU1e5B18NXkWeYodIEY+6SBNNHf6f7bcKAsizo5OUUf483fjp
ZMTsgUTYPJLbAzESFgBoF0irMCUic1ZUyR+xI6jHZifIJYAAmCy/tp1rBvNxyhzn
jK+AnZtAptc/8KPyOQL+e35M7OtrBsIMNwHzmOL3XCsKmZZqIccCNeu2lL4ekPzc
bVXJLBLSqhJhjS4fCriVDzPf8lWqQR1lRXCDAteITVdEEHsEBE91JQguhpkDlJ59
SuJIPD+E1seiu8IQQo/2jK+JHCfiXDhXB8AzXXkRoCY6Y29hDdFErYlHXGlzzL8v
HoXcFROvimtFGa9qUrze4o2QBAzGP0rjvLRks84buix/soObYhM+56NRNgL5cyvK
/NiE6Pl8LwfgzXrC6gQFcpfK6vM2qYkqnN2mvL5huQFfXz0RSNWXEkR6ilruxdgK
GmIl47FUfsynVnx//yFvHLVo46xJQ0ttzI3KzP8HbbQCutHLkY8+CBAK0/w7pIlT
5SgV0Oxduo3tYkon41gH4drZKlsIBXWNUvhdosAohKgOWEQsLvqNdKc3NgKVX7/b
brdNGDrogo0YbNHjhFFcGlbYfNJ5JVd2/hT3ubJzBgdSWOi7qs78CCAvcYSKEBiO
z6sxQyR1hs6zeFbXD7bMA0WWOftVx5geF5Xm8ZkXhOj02rp63noASCP2E/2Z8Djd
vXNG52/nK5qK2M3MCdqaVZOiD1JqRnJoycb8qpcep4y5t6Nw+A0hxDTEWnN63/Sz
uJUPohJW1djkPFGRtzOPFlP1rd/rDE6zm1Hkcg5UfwaqBv3nGSk+JhXFtaG42M6m
maDaezNw4bn2E4uSW4ycvLUx6LYvqjcpO8oXHEA6Xe3f6NswKUt2iGV80mnB/W9V
IlztMdCenbvNGuFsrEowkDUluQfF2tm/wftYlB8RjEo=
`protect END_PROTECTED
