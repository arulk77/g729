`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAeafyzqqNwBTBxaAPdjiEdXqLvkuVWxrda/UcfXvsnwS
7n06fGwp3kzpe8Gs7gmPz33mdI3IUsBQirdSSBL7cLyv3kV135Ykj6JWbc43TW7/
KxjEz/0qBL0XXXKUhQymHtCru9fYp913Ck0J9d2ncSV9GGGjKTbc7CYMdehhxH2L
f6HiH/nKHaCQvtEGFDVMIsWN0yb8xuyU5x+wyJSKzz1K+ZsF0fSUFpdAYz9h9vnZ
F0+tI5zfqxzmrhHnBP7ETOdqu+n5nLjRWFfcvCi5KecGpr8/eXhNfeZtDW5SvFZ4
ci4Gbcku96ybZaPKHbW2pmlyrf2EtNhlmldjmm/pajzayrvDwcMOzkW1ECq6ZTkV
xE0QNaCJN0X0MVuGXwrvEk8IJqa0+6ak6YNXApkpksgAKd/jfQFaI/v0Ev7n3V62
9ooN4PySU+xC3ZIJ573AbWktYX38uUGPNmutUIwNrZTEndyFFuxnsqrLc2dBHS6u
1SXeSq5cqZDGqzZgw7G1uCGYJOFRGkCupsgGiKiCwf+/ekfQFIpa4WMJ4wlVpZn1
mwJggmZvncwcPEDm0XkqrL7E54lM+9pYPP8EJnZiKO9oVqYwgiJqeZdFD2/DIvrc
haWT+6Nv0PHyK/OS7k4jOddpBC1du8yo2fRJsasrqZE=
`protect END_PROTECTED
