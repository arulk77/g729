`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHo6n40dYySh2qRqD5ybxrkJGFgYg5fXPmZSwxsmb1/N
LkH/kYM+TAtMf504yjA3yQWie5izNtgYdCrTW9oEjUKTvy0l5wB0K6vhsNt2htrw
7K07Rot8Ej85zuifUDG4zK5Hq/kNInOOGYnohQRqMDS21nt10JULWa/gCtzQLJm+
mGs/7Y6YVHG0wEkFmTNQrwoInwOCyplino5frfCZNLUivD8XOuQA5zpYI2PZnSfU
iQg6QR/wMAR+16P/H2Z+YJTo6RNatFYhWzwoMV3ZDSV3oWWMwtTF+1uN+Slf9gOb
nAK7dNs91r7JGwg9dg5VkSq7BnMJOX705rN16NwwGiI7twxrkmu0dPnETV/XzNWi
Pl0KnNwdwdUFlKrhuPczqYbO3cN/KUrYYPDw4ciUdoIKqLmmKvQiaBS5TDpUZ3R2
`protect END_PROTECTED
