`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIXVTRopml3pFzeFYMzzbEuBPjH6vfglmEOXy40LXnmW
EXpLFoW140EgPEoWqojbLfIedLkEe1im7jbStGDsUWogoIyUGsoY2VJb7Uu5ktVH
ZgLw8824EoH00nk5EbXIdxBetw1EB42VGryZuzxtT3dJhHo5zKuyxF6PDoGFqEhe
SXUlu34+7AFhF3jku2J3m2PZwgkdzPdo/2aWldd5cA9Es1Q7gQNHX5OxHhJlyw4A
rsIDp/D4bB98pGr2NBKkj5t5DvOtdnI1R101voHXZQFtDiQlvN5+rIxGLK5GTQcF
ajUi7oP1BrZGeXe0BxCbuQoTEdewtBsf0l58YsLjcNfH05DV7ZixvItV3w5GIuZI
zkiowWbmouI+p3+eWlak6E6eJnsNm8GpO7tvOlRIztHHhpJEUzBJqvugej1HUWDP
JIDH+wII1inlkpZAhG3kYtJ+xDevyx7y2K24Tqh3R2A6nXy1RRZkV3rGty2KN4Tr
SGikDAZU06UEH3BLHjdnYfMBYVHQ6RPeq5Az4kwK+trrSU1Lom0J8YaVrbx0XsfR
`protect END_PROTECTED
