`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKaE+KVi8szbcyX1FkqQ+RUBenjjoDnTcQgIESvvJCk1
5BL6Tal7gSxSsqS4eay3uhNpEKhnjuE0NjN0gicGqQP2R8XtdTw4J69fMAbqHzOS
BzK5OBjc0czpZ9L0nj78qog1UAvtT3wOKR30f1lAgohtUp5W3loyBqG3JIjv7Gbn
KW97wsLwjWqA2Dcz+9RJf0JHx7W5z7cEpKlLiT8k+juCf2hoqpQFC14/YP9m4o9l
HjNhyK3oTzZzjsoUl0jg1vLzRBSU4MKLbvwBu5wruiStaLa6AnZGaUePy6/XpOz9
QjNl8bMl76lTXTu5KG8Mm/qNaW/nk1Ys6GAyp+TsNXDVk4ku1NKj6TRljR/tS+yr
`protect END_PROTECTED
