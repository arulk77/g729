`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKTmGlMuB+iK5dTaj2z8MMSTTso53FDXBObf94NA/CIp
5x8k1+sfGDvdPvA1xV7o3I7QINiAP/Sm0IOylsv5ihSbbNoTKO0tgMfd0Dm2X/8v
Lhu4Uxr58REUIswE0fRnNUOcIMYlssvXRTxmYpBbyfHELhnAtwOToo9h/PzG3KkP
oaT9hHea/gWfeXyTwrBQUw==
`protect END_PROTECTED
