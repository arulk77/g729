`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
whfZdEhQhIVICrvn0VMg7oD6BCZL3IUEhQeVeA547Zdbnqs7r1C5mbSUMffX4u12
HJ6E2DHPsHBqHB5n52yHj6GTvuW5WFtCRAqMdXeHpdCcn2GxNWV14ysc9TV4Boqi
Cx5Iircaml2O14DpJ1w9zjoGvh7qcekBzKfVDJylDk1OgWh0E2igdjiCSJ2Fhg1p
CWCyxXXlbS5/2n3TcBSOCjIF3+HOuyu8FvZm/BNbZrhSZLA0SBSHa1Vg/dROdUOf
mDrFNu6jRI+JIT6qV38l6f2MdDd+0QG8U9P50pPLMHpa0f7VYq/fE0umZYfGbXAr
`protect END_PROTECTED
