`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4jUYkdt5VjR8oFbu7ZiLkuHc4iv0gDRTbwaiJYJ+7Cypb1MBsZrScXFMOIplwYMg
wypdiUj+l6KG55TN9zuZtOHCp5k863cA0Axzv/79/fYM0Q8IwRFQC9/cfLELkF7x
zX4R7cW8Dip6Eb+aDO48QOoFnNpjZtfAMSRqI5i2MKUYZbs3lniaTrT1nHDxCHmn
mtmNokMwAWPMjESff3tQ+NLxI0BBQxBBBaJNAvYJejAPBIu3kPtXbkZxTiEKrjdN
`protect END_PROTECTED
