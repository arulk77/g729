`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aRL+aDJtlMELY3KRQyeRUDZKImt85qiqZ+Ym+ysojBDQ
R9QtWlO23UaemBQoWfZsULcGNlKf4Nz0pxqRN7khlX8LMYtXqz3a4j9UVwTdweQI
ix+FmyfPCi1cw+yMjnwxWB8AqqnuJD/esQX0FoD/BwEeqWclJOpnDjnEgIgvLPMl
mtPse10jzuhnFyPLMF/4gK6SM5gm1oIcZiRivBjSvOnc/o9BDV7De1bGF+UlftVj
Gwep21e3wNIdQ7ZFzRzqFr9m7kLeTcDL80FWYSxyhSUHi5Y4RD9ca+kZ8iYfBvhJ
RXEP+8TPuyUVLBSssdpE49qRu5OHNptJ1L4LnvKACaKDho+PNmlqkg8t2vOen6mB
`protect END_PROTECTED
