`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePVq5712KOCS8MmdJoq+5jmWrDHtN7JaTzXv/aYA55av
E1u+/C/aPYgTq8PowjJSKqW3yMo/ZGpg36/A+8lxkL5u7LVouheZj5f7hXY2KEeH
W3hFwsKSvBbtfkaBu834WU/y6Stiz1XLeOaDTIzbJRpQM8EK7qO82Gj9RH68mWBM
JWLu3eyfaQS5F+B11SLGB52Tvapa+7K+97mVehak2mMPljlR85+va34cvQvFOfum
`protect END_PROTECTED
