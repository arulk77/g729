`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDrtsEePUuyr12hQSpowV8ElOXnt1kMukxOOagyy1+dL
IGLqplqeU+wD+FaMgipWbSmA9y7u99BoOyU0PADClElcm2ZjCxUXWCIubK+8Q6hl
cz4ABhabYO9AieNO1rTfM+OosFXvgt874vT/EEF+fMjmbaazemeAd6U4cqWxFh+t
XqW+2g8cJ0W+msJE26Qirw==
`protect END_PROTECTED
