`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIN+nWdaOfyY64NqTP6O4lM1pjpijmSBwKJTG8oA4Bxx
Dpat20IVS7vXL0cPzUQYFr58gi+hiznf4YiHPqmxaAYVf8I6gwdRxoRZgOhMaOPL
5p4P1i0zUO4oqzO2CGsfKW9N7XOREhndpD3sVTJ9kWtK+RZOjV24r/suiX6QVAE8
`protect END_PROTECTED
