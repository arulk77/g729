`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
J5Su2kmHO4OFvl1OdV8YsQUExsxlZurMFefJWkhkbNZ8bpl80/EplNE0HyEXHJEr
BDD9yuBxIFxrZHvSLHM7RHeqOjNBtDy7m90IrImHWp0aUR/Ni9IKHFJhameWw4lQ
omMxmCYlDion/vLxnllBuTwIw9IxV0dINswJ1M5hsPgrGISKIZ2veGgFECm+Zpq0
`protect END_PROTECTED
