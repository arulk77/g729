`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGARbhhvsrYoqOALLNhIVJ+juQV6li9I1Jq5nJiVRh2d
xh8iCRhmbl74OAq1hDrqGWNe8zr1/7Q4r6/CqNYX52TP3e6hxk/+KzZNq6UUTsm2
O3/fgPjNQSrt6BIcBE3PZ6bAyVLRkeDaz4QBIRKTXd0WriwMsMB/izyKMjsr3nxv
+QDFJVTQIDDByoaDMewPh7/dRnyv2y94MMz0XY7L4s2GEzTSv/PaWvguDHyu++Gk
GiJKX6ww4uZS+mv4vzv8/b/jTeeM0yS29G4EdlzO9R49bw5kwZOadT3i+/6VMLa+
KUBPVmRSHn9t4x7yQS2W3iUM2uUfh+qSSRCtdcRRhErdvMKISSSTw0qWhhGaC76M
UgDhsQDM4AGvqyLoUKDiTji9kPmJ+uvoYGfn6y9liQfV5ut28t9ab1uLAvPbN18x
VHj/ETTsL1QJSRdInAZPUZqzjrNy2lcX7nfctPucbqxyEh7SbaWLEqbtFv4stIeS
`protect END_PROTECTED
