`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMTYUa5MLsoE+u4voz9ukjbTFDUxwsySEzZbxZlgKcG7
T4uzmx7HnJuinohuYwdwh2tauZh1h1M62WYSZhqKsKRLrY00A9xPiIkhvJFM3zIB
bIiUnX3uerBJ0JXovJdgcQsKwH8uxK8BkDxB82Jxvijhtd6Ro9lFqKtQ/EOS4Pnf
m0MsYA8RvA2xe1hifmesjg==
`protect END_PROTECTED
