`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOtxPAZ+5PDhlq/Ri6uJYxFl23LB+MubYVkvAnQ4AUEw
hYBllTH4c0oEgGpcxs3WkNNhyb9HntwKCT/ghIPuFQpFaQXerokvJ+9hZhOKs4ko
cSnSn9R9+fzy12rlpklHfS3Tml1mIeIP/ckWlqzkdsCsWqsANnQBOJlJoCC/3ZFe
vltep26eA2y7AtDcHiDd7k1CARsJjnVqhWe4S5pWsH9SkZwk5N6uOfhuH+62bmwP
QNnQ2LWzwdUxY9Vn+7/yE4fKUcA8y1QpJt3vwHVkhOpOJQEVzV7S57Ulm7uzN17Q
GzpIow3CJ2iV21/+Z1AoM7aN7CfXaS6AMKImFS91f3iczp/lNkHc/pIZUvvQrYKp
8Fo0Wl8oc0ZwctVT06ufMY16A9RKoXEKSih68VuAZJj5TYNXucJ++4YNLgivFoTQ
YtUBwdOhLV2gsec/4Qf//yndnL7lu/vu0ZpaimzkBZmEjDBWDkHT184QxH6YBeTm
y60TQOarxFjvd9NqHaIIgCFiUiV2sDBhd/Nwj5ecvUgPhb1cz046z3uGIF2khgfC
/E3sxIVguvZyjML/sJ32QXyPg9eYOlUNjYopYrUliLQ6or/wCV3lAIfo2MISbywE
`protect END_PROTECTED
