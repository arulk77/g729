`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKb9BKRDa8KUP3Rv6KzJ4JQf/syE8RqEXCFE8+eE7zpj
SPidjDhnMenM5I50YxHkUXnSkfw4m2FmmDM3h4gNndWEEm36WzRU8f4sKdGNzunL
mUW7aweZ3eWG7y5DhfUV+h9Kh7RPaGDq2KnxqUBJuY1+SrHbQ8cCrtEVg/71at04
JZcsyRrUzgqDv4VDW4qgqTPVU5ujXaUaw/TBakKS61ptJFrR+O//YMUW94/p2H+3
boSaoB43ax6V9AdlTAgCsX4Cu34Pa0zN583XPR6w5Z+SXNlpEwUEBYzsjge93uxS
UOQLWArDZc7uhw69HVZYnsz+Sf2nOjiBf17kBrXaAvW75GRks/HtlihrlC4IZ3pL
MjD+n1zt+gsyjzntrlkdUkVAh03UN+mlxhB2EPV/xG4aylxqeLJKTyyp5TF16A7A
jsWkBvqWTNK3mjypi4MmDNSbLXWGzBfsdhtT2ircT5O6Zg1hHEpig11KjkL1Ma/s
AFTFGBOJHobE00f9jQ6w4anH7ODhlJrUX12yKnzgbNTFmXHE1sg0CM6uTzv0lqsL
`protect END_PROTECTED
