`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGe8anleqOi4etsU1ZCG6+Lc8yFUrtPY7kR5Oqgip9zm
TTWS8Oy3+e8XVmLAxeiyIcnZt28kCl7AyiICM1Z5ELaqrz3JSJn3pWqweeBerGxs
l+MuXSTgfDsCLNmkLrBpflRicIep1MsVK+AH4a1pzyz/DFjaCx+BkVc2VTpXUH+9
njmCq5atiQUvdmBsVAjXv5RDLTmn/JgtVXP6Te2x6LxAn4MQHctDr49V3Px+Rj0D
leEztK70ONvhMhGth3rMR4L4QxY8V4+v8Mq8y2rcZK5HNvJhccUhy5B+0er6rc69
7afByX25iQillcDrmji7w16+8uyb/uYjASgBB726Lm/eC4UNwZaiM3frSJ5/ggxE
Ajc8+aozcwjUi2uVR2cfj4ulLxjhlsrQzEyYb8pqbZFnWxB2ukMJFUEBVLhB4VdY
oasqJUboNbAtUgfDDoBR1zhH5S7TlTbR1ohL/ZKj9pyjanTKk1dmVcc5I7zd/kYl
r9RNN5BZRcIAwRfeZutUzh4Gt4WaXiV/BkiNNuLu5Hqm+qIeVNhh1qikjGhO0iwi
`protect END_PROTECTED
