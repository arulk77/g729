`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
iafOB+JiRx/M3UonZZwPnas+TUuxnrnlbzspTqR/1zmFElMm6yAwAYKJ5lC4lw5w
ZpYV+stfFyUE44XNZBCQaVcmdiYKb1CzZH7zSnFQENKJXmI/jaIaKEM1/kkySQBU
LjM0KXZvKGRDm0EZRwmsLfOSHqILS5FsHyfsk0wfwglgWqLT3CGeeEkDTf2uwZMJ
wHPvG+gEaQ8gdX8SE2QOKOaXufyFkiZKG1Ie04wFyoxDhAmsWIlwGPCua/uN3jqR
uzAbLQ7W9oBfGXncxzyhvHlCD4+hK4CoyJq3m1Ph7q/gFYhT0m9EK27yKBGdH/YP
6G9TVh7EfeKgVwDiR4KgCgP15xbf7Ys8YaVNs1iqhejiivpC0uoAqzn8BS+xhOel
y2RcKXb+FcX7w6G0dcRzFyaZTOGEoNXHX7uBvNwhOsI=
`protect END_PROTECTED
