`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAWfwPPOmyFTbxkC70vyp+FsXyGgHLdhao3h8z7eYQMUo
hh3v+wmnb8d8CK8ioS7v6ukgI8lGUUEDpcRVh/Xap0FY+JEzSSVrixnGFPMROZH0
uG/u6YsOOt1OjWSoVXsZHoi6toF63BW5pgrivIU7M1dZLUKp6OEDr68kCEbjYrqA
5rcTYmmoYQkfdhHFeQMX/GLDtqavtWWsUbig/1m4C8APmEPia6Dv67P0R+wVKAIP
Yozr63ahTpN6WHH2a7aXrKJYpJ/2bL1Uf/Q1dwsENkzaJ4f259pPYLwW0BW3fo+Q
04czCKrrB8OliXloQq6yt52cqz/9j+CPwL4krwMsR40QRXKNWSqbi7FqG5jgRgFf
xB++XhzJXpH5yabGRB1ZDgy3CaMX3LQj3YRhsR/rN30OfhaGKgv/Gjy1C4YUCoQd
Ekmiv1DziaR9T7Twqcfdts+9D3K/Q8tdWa3fr22F7xMpICxyvuybbc6LWwcHuRMI
lAtE1Bu9eRZgjZ+A1xhN1iYj5NzrrhW7iGzvQFSUR2r3IVJElIybB9Miw1pn1PTJ
2paIs6l9p8oHFH47tyfXgJHcvf9kXfjBlJkMTCNvi5HhJ8R0VQmUzkXJ1DtnT0QD
q4nUUhkaK7ZWju4vPmutdALlFAy2W0M2N8+vrD1nKk/nlboyJtL1YAvjBh/b+4fO
KbmCsyJqv7Z2INPe7x5VZVDK/ny3WJrWJOCY9Kmqjvtg/BRp4UfMEBT/nVBUM+ho
DWlTtx0wLskQYLxmcDuxJVF7B4oxfQHGePKnsEnEO4pow5w/rFOWbNHOTxjyWHdY
BUbjxQViswrQISodFblNh1O1rD3nI5Ewf+b9GYE+W9AKI/gA5H+JM2mNFGrksI3p
u6qrwPqJZ8uqI6NAKTySggy5f+LcHxLm7hRUQru07oFyESe0lY8I2//eOjbcgHwD
Y9Ed5UX+yYxA5vYT8CgKbFhvQ3gADA9Rc5K/ZfhFFNDnZfCA84ob95KVansfhhw5
`protect END_PROTECTED
