`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43W+3WvyvPsAMGZrISf/YFSdXdm4Lo5FsTdvt+UqWT87
OUzP5MDn7sBMRIrNbx3iYdmfzUUJMFJRxTatbKyl4341p+wGulQVPSKqNwIDO7J2
tj84/ohKlT5I40ud30V9vs2TCylQqM76Jvy41qZp3FZPG144CsI4Ma0HS1YeKF5M
u7105cUfNuAymXU1TOUWg/axQwwM+ahh93nboLZl+afq5M3ztp6i1Y9RbEGgYmuk
naSSIKzPVr7t/2cIhJgMYr0FeCanVKm9FZrxACVT+OLAAzW0GufAp/DEpBzDFyQL
nMuGBw7TbXxzUAs3Ho7q+A==
`protect END_PROTECTED
