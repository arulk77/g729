`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47o3eX+dH+un8KRqxMOtQqTF1qx7MeMTPti9Me0PQymU
AvOKHQTC8WvBpxJONCSIfS1KOrQgn5NVoZMqrPKB5kHZguYGWrPVL6vtJFXBe3dT
J0nlP/x0j4euvVkMlB3gAU6Bk9zVjmR7cOvCTWzTrgAn6c4L53+s5QpF8uELzdi5
AWPQdLipT7DYWUinP2aT938X+mKH6I+JpPfqhCTRD0WfgVY8Xi0VlTysgvyAzkpU
MiDvHhXY9BF63VvrYgeiWzrF+hM/HIP6Slm2mc79I5ZoiXUjSuTpYEosJT8Tiu+V
uTsHx7fxw1tIB+NRlf6XRuPQ3Dn7xP+tzOo2tBMB3nlMB0Oym+UW1MK2jSkDcS4z
S00ym+20BzSTJNK9ngZbEQ==
`protect END_PROTECTED
