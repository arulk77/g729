`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1adqIz0jWiVhtkbD0oAYWPLpnOmD+VeOAuDAmJtq90GIk
vc0OfwPRH1oQPNfkRIUQmcW+W0D/qiyJfjiRaknJwHeDpRMVV94B/K+L6oEUEM/a
wfxa6v0DjKZBguELASqYJHPS1QJnbz+CddVASjkMA+n4a+u5h7WZNnGPxtaNpgB8
ljgGcvR8PbU+Tg/abSWCTFfHVAI2mzi61Yb5+CxNN4G7SQ2v77lzGkFsRlvpuNXb
zq9ttVF1sYRAV4F2gKXbAAyDtNxJ2kiNH/2HgNoYLaUMtzB0v3z0h0znkQdOuveo
thHqI3i5rePj1uUDfcPP5/uRJs1I6Z3LhnZc/JA4r6qyf3JMQA7A3zj203/A5Z37
L4EBj/wgB0OcMTa2QsuRa2x0yJf2v5le3VpQO36Ov/EoiLa0IkTDolrnqKxFpChF
g8BbTpbKY54w6z+DLrfPDUIERmpTZ1g3ORAkjQeR9onJ7/yEsBtsBbpMtIRvM1Qd
9w4vXXM8/7oocPS2Xg6dklIQHjX1LrHr56Zga86A9IUCWXS6ZHa+b7O9hM44FdB0
y8IvjtY6UjIzKuTSE/uYHjWi/IwJFgRmqp2TezGCkvCJ8WdGTpQZu3JdLYXFDVoE
e708v/skvMXsqgapdv/FY5bVKfiTNm03YFa01cHBgHpSdvUUQ+WvYmbNpZYvjVOa
CrYuNdKwrEAzEhiy5HXnzLXKip6Ws7E1IGhhId5Ce0NWFQONiJKbJUPhRvl8X+7F
qS6jW3HXvCy89tfIax+Q+YdKG5zdB+dwjonnrgJiQ8/WTXQ3rcH0OlsAqqCVSgWc
oNCetpKmzYSgPm8wMfuE+mTf1yO+RUruMh32ePzN5GD5rac5vjgdLSmUne2Z8EQF
TXB1xtekBYZAWCgvo0tN2uzp7bB+7TzT61f2ohU/HEWOJ7rD5ZnNQGM8Cw+LUyVE
NIFQ05QLAZcSzwH26S/JnHSnfZT6s/KOL3gPo49Am+ilBgTbUXGKPNEQZwpyH1lj
JltXy6dZq9AY5hzTBhmaJpEmSIfXSNaMWYPaTOpUD3NDhPpzRE/QZwM7jDOSAHrq
KHqAhK9tEJRCNxAXHhMfSSqWCfgV5h5e+/fZNZJJz6tIyjzeU+9VZceO5/SckWDK
tPlKz3y+dxOJK09WrrG8WvSOOOBU+H2rV6lc9fQybVv16B+NUOPo6OHZf7Rr5pYT
LfE1l24F5fYWCrlWGuW4juftkEeHFUSUP4lqwlN7MNA1CLssDgMcGGyh8hZCk86D
c1E0HEqIEnFRjPm6N+YBO00RWBMggJYz0AydHEyrlzSSzM4I2Y0Egd1ReUE0cFLv
gHSkwsYaw1Oimd0oaI5gHviW0shgsb9HJ+B5JmCFabyl5I79UXgtwelgRROd6Q9M
iG3OUNoVyZzwgsQmyXGvPxHcUUstcm2MJBtGhZQgsubZOpcofcMuo6XCNGAP3f97
N6nrXm6tjCsvCWjlcrHWgccGXlGXnRH2rf/LfIgfrzzwMms3k342euJelC0D/1iR
AC8zZIfm26QPaadRClhAg5AbbQhzA3DQh1xn4xr3AOzehFHrG/TmYWwCkkowMlhb
DWmOxKkHOsaLOb22FjN/WJpH/pPVbhiCWRoIsmKzFjOvA4nLOx3CS1w8bv62rypo
IJnZfU7fy7qIfP3ZNBjM1Foe5BF9uAaSNec6e1m4jTfFTuwg1UCQP6i2et1/7oAX
N4oSnUzbNQnvjsNrflEZzmcuz45SH2RRowapzB/cUS8qwAZrSN/nuxWZnC263tvS
vYUe4UBHxsVhFUeJAzi1ktKUg1uneMXdG1CtFeF4g3xWNFaenHGOsRu6JtimM/x1
KfH1M/CIOKzzMxcM8ekdUl2vVDw0qco3bhms8KvcAgVmiW4lgH9Y1tOCEWL1HEXW
7UDLgxt4tr+nIyCeehOu/+Cw+bmk+kvan7tghjAxU2pkwhukm/+MmBuxA/TvE1WS
xxB60dYWPOqeB9sVtr/yjlJR9AyXb+fzdM2P1oBYbkzNpyUe8XAU3gAPKdIqSyS6
55SXxkdPKDWR9ijpYks7khm8ZNPjz1OwfC9hlObevuMdSqNCX88O2O/YK3QkfH9d
C/HH2KhcJfWd74HUJLaRKTQbAQn+nf9maDZltjfoTqRRGm58tJHGG9p3sIVTjEQM
EXfcVEGW/DDcmBdbmdyXnQo/iRJe45jXbGaPbneS3rthPjzvHcOGZMD7nU+IJv5b
mGhw7UhOFGEvpAsZ747mxlt3ZYzlO8sZBPJEtnGt/Vh6s0oXzwFYnYFAMZcKtNB9
x+J1+o/jib9oqXASzRS5HYjJayssyHfXO24KaJE5GlobsqJdK5wGzetDgkQMlUJr
Z6GMsqzBTzXCEb4o/f4PK2XAewrK+hnv4rfAmycByyFEBcrZs5Ro2goy70gXyVGk
SRMBB/ZugJEHSL7s7WwMTo7UmNWnnRYo4DSXhxhoxUwrb2c7qQJLd95RPin4nj8q
BPZuyqB5KfFySX920R7k8qIzqdf+KYyqru3XwPjdpFBRjv6090hp5EeovauzQwsu
3T86o9Y3tbJeE06Xx5MiALzOpbKLoZQCeL7bqrFbiZuZi4eWHdcXfoGtMcglPSHu
1ibYY0oT2s9uafVVNia0owlYJd1KFJvjtsU3vZf5hXJBwYCH2qS/ZZICn9mxpTrM
9pKXEzST5THEOYvqhjTI4569Uen515RFDrS+rDxPJNkCxDNP9uuMVBybI72F3Eqo
J7j0jIJJq3bH+19eYnRyQ+7x2qVZPgFkrlaTXS3+c0MB2uZt65kxDgnjn/QsE7zn
CRg+3jbjAk6+sHyB2Dg9PGtjNr20w2ZM2EDcSEsRkZhTsbwasG5yLNuaPGXrmCZO
G3t5v3GZFva9waQnYb1zX4eEBIUtX6GLEF92KBnuGweducC5KsCidg0DfTgswjg8
o2y0YbAXpsPAh+PaxqNZ/8snRWigxEXfU9RaqdHUXaBiz4Gk7MB+nvjA7DFLKjDp
Y5HXMG0h53nuHr3ccftTm4ceoZkfQZXBgw5zfjSpM+RpAx/dXx4Z29ztY5lNDWq8
XzLQCKCnJz51GJsm0lsuxpEf1oUWrNGn+bkr00uAXWybUCi1KAj+owo3SvYILZKb
jTqUq337lFES7qcLiWn5FJLKu56shHjd/SwHNJaaXFtEY2VDHXVh16WRsvrB0ss4
MtLZ+luVQ2RXiNotOcDU/bYBTjqMo6l26OzT1GWFhnwLDo8osdTUI43cL3dJqtVG
Mm8A+U9DyuhBfX9v7sJ5+i3Dk2+c9sDQgxEs1m9yy6MNzSMLLvMqTrycKm2+DMcQ
Lf8+n3lr64SfXfHHpzIAGjsdKN1DrAtli9DskdmgG6KB5SPwvRj7FQ7o4DSpJi4g
z4NfiqgwDj6YP1RqBmglGokBRbefHpQN/PR7GWLnXEe5U3+xz123S7/8ZCV87CTo
nXtuXlpioW8EmLZgMTdnRxn8ZhVof1dcCoHhY0ztWO/HttuneWRx6jzaOFLH9+xF
JEQB+BPuTwJL10tjcoIacpEkyl9dOasf0dEhAosOsHoAFOz2O2HOtEoLetQEjgxE
PO5ou/7TUxD2dFurJcNHIYIpva0jIQmlzxA/O9ilvXr+tA0iOwZ79wEuza8yi6ru
9B0xNK5tWZLeS4TpRiuA8ujCrzWUAeuLwYnkF4HgaXTi/XSC3KR2Cezy0/SUBI5O
/zWg8gOoEgbvIjGhH7Ip8XvnVdwDHko75mo3dGQQYAH9oXtMHbNgo/BLRtvxpG9k
7BTf/23sQ17lvbCBULNk6kdZ7cGgSwu+RHe/nCPHWFi+pUyUeSSO3/Jv2KzNWoH5
ishAeMisk26FhjFshlj/EV/BRflcKQsWPZR2lC4Kao4inWZeTX9piyGeeofTFGOc
Rs55v9rabMMlnVyhLJWvUKxw0q4XVwLsI5iJkla2piwkqvdbMtbwK6vWlYXW2aqb
BE7m4FHwCmLY9l3VWrMs7PxcbkkqXU1Y5ka2FK17SXKtf7xGuNilSIYUOwEDZVXs
4mpCGG10FcGvzWDE0YPxLC6lf2qtYCjkX8DDv0KVLAwbEnk5Nj80PxwhuI4AAyK8
Q0iNrthOEEsr+mXH8CBMm2o10iywi2fbY5MMKX7UI8JdqFeI2aRcgqZa2DrJS04b
kp/H8WnkoqeQiz6gR9HUd2VZwYYTjZZMZT9Njhw33R5qaBUM3MtDv3HjRoZumyCZ
5fX3NQxoTlbb5ZPfE52FhAa/HFLft/5R8h9tZXwmhIeOdcxqrwbIviyhhl+epOFW
yFZORt+iLJPWzZOfm0NBkNzhrB1dxzz579ZqwS+f847NoHPnVvLKqc+SogYMTqON
xrodS4/EH1JNtVFkAsbYayhoZMAwKMcmlM01RltTjDS/u7yz/2TJuGl+E+N2tlMq
G4HYr0WXciS5nxOZOO9qnWCdQB8j6gfNJyOvvuWW7z82s8suktjAB1kjUg6SpScZ
e9EIjXZuRQdvfbpj6snSyTtwLR1s4USV6jy/0e1lRmFxgdlsbPtuSG107pJxIxwB
SXSlVtRreiLbj7RvalfUjQC9Jv+p3R4apXQYXP2e3epzhbhGZpFZICtlM5bBMBc1
EW9pSUsQObmLckUSsv8d+Uo1kR17lAgG6zGRHsY0BW/Fkt1mQbEvk5ZXwsClH1Ta
TF7wj9R6asqiuf5Nu7lLIIewlNgexAtWp9B+b+IREVUJ+IZRQyUGfpK4xpsV5qUY
LPbrIbPcy9J/md2/iY+MAJ6GKBVk6HOUKBvUjhFmA/q0efQU9upj7Da5Tvb9/Xs4
JBoGaVwOVoYVAtJ+yzv7RIO215/d29vQ+o07ZLMkw0jgJMNhbcY1lPw5Lei4G88g
2O0+Buo55Zw5euw0RoSB8PIuhtz4TrJDw8rhtXv7DhWWZHL2ouv5MQ0CjbsOHrex
MT7fVmQK68yMz2l0Yj9AFsOReGTk6Ix2lGymxtryoFrLtvTi54pQILX01uEuMZg5
Wpg6Ruw+F+ZXSb2Qt5tZi1cirluL/dH7b5Q34QH0tSSBmZJkrf8ZanZXogH6lZ9b
j1kAb3VvZCSM4NltE0WrpuJxFAgn2zdHtfZf9OSe9h0CB4xOLj16MR8Sb7ilezey
PnO9FOZz2Fzb+3DNsEx6eIgeWZYnHIWGmC2ECpurWMFkzu0xoaiPXn4djmdKvxIU
uFYcJCcy1kKeUdXzYKPPUXbRynJ66ZUSQq9wLRe6Rvr3BPJpN5a9l5ps1b98Xzrp
3D602yhvmfHsnOl6OyhVRPrz1fNfctNtskfDyLITzOu4HNOWYvUAA2IQpZ/irDrm
yvGVMDAbI/NsH4STAzu8GjHSJntYbbVYSK4pobT6v4xOKyS0rs9rI9e5pGPgO8qF
GwtmOycv8KEDr9HALpI0alftlNezVAm4gjUVBHuvVRIMA93akMuB1Wykr2ei5WNZ
8J617fhTRnRA2fFpUxw5rs0GQGVU3rEYSpBCAAZWxpInX3oKurzlhnscHYF4tCgs
sOOc94H8m8MtOf+wVL3HDp/sKpseIJsE7wSdif+0ykwPbPZwuIj0Q3AwqqxTy3kL
Qb4gUYrxIs1v+UodPXQcqc8y/e6VvKRjNu8017FBiyiHRsHSGr5+DXV7wxh9Msul
coNYDvMA05Pt5ccpAiRttpGjPCKpgm3Po3kpAyMoxViBhlOxp4RnenU9oOrb6ToI
YFVnnarDru8WRFZjYXoV2weqyGAG3FJ1mtcUAMDgASqP/BjhQ7Cgh28rstgy7bHH
OERsQop3UHme6fAa5OdYU6lVNxNwpPEXFo60UcGzwkG6IIMSun523hHJeIK0eKJ6
fXfe6h/1mxOtDvd+Krf5Jg9WhLbe3ikc6q331J3csLtVMKmlducbDT3Zzjvd23SM
zVfUoRB1iJvzIgrX7ay+61ht4UbqO8dIc/qVjyUznhjCqXISnguIOrOrL53u46tp
88KybamgGbULpdYYVq/d/DwUQUfcJTKvL5AcYQu/VPb8CUb/4RvZFVuUt0dxfpyT
t9VR8gNjlcC3xY5VfmSCoOigE7YHLgIdcWkmWb47umKboFHdx3Xto0Lm4g+rPyIk
onIG1WhCsWY2h1vZedaSd27rpMwjd/DbVmA6hwWU60sq/eLjkGl0fgnC9vvvZV7N
wPlEsnVDIdNggxI/i6Pmu+YwWFfEf4P0oXrX1S8I+cHvL5M8VrI3dQ/orzL2ORIt
RtJFRoYW1EO2vhcY7HnE8T1Trlg7Rvr5BenQDapbZVloDdn3yfv26lkNnxFeDrkC
e0B19mm8TFXsJc7xdiaud52EKbrq8b0em+LyUVN9i+GQIFyt7nMRhJCH201+22cp
mfbQiC82T83HSe0PQ4noJdssq+OTHoXws9qLM5lkkBsEbfPf5sQGOeoQmgqcdnKC
0cRWcYPxDwmopnMz0i6UE5tEf1kXFdSQuctgN4JZDCVutpMKYwrJquDf+UvWwFxJ
kvHRcrGx0wOh9V+brCgatUtmGJjvthxktNYMrByDoUxgbjhwobSNYehTjfA6wOHM
140drPzoK5Vcq2WubXszoTxCqoP1qXXvQs4GpL02x8wI6g9jj/PfBuSkVQg431dQ
tavCqO0q2bcZ6AT+QqWRNas10s8g8QEMLQTSmxIAA+noNCdl9NFK+qxnX+wYg/9i
KSml/MFAlljS5NGpK6QXLtm/xIyEZvBsOIOn4rlKDsnSgHw+TIXYTGIlJQvuu9/6
2TyUJm2PEqWVKQ/bMtN3q4gDyC9nCDQvGXVuQWEqbFz5WaJlHR3TuFWF0SctU18X
AHrtyh/yG005XpqVPPPWh8rJ60zGPqLm8ERB6xAWfK4DkJO1n0/5WLZun8f1tVzk
g6ZfmJOPOK4DxPn4LftSXRcwK1nV5PYpTjcdJi58ZuVTOglNMvTu8l5797YUDJlk
c54JVO8scnYvApMakCrsTZj3HEb2Stk1h+jx9KRoMLSG3bSFo/2s0YCoatBeaKWF
YFaAiyeJdzzcSMhpVH8a2JkSM3T+lWE67JMfrgoGANZ+930boGW8iGmhti45rtcL
HzipauC5S4LGUKhDxaK/5ynVf7+i+qLWVlIRJtPSLTWWzq4Xm17BcXQK7ukwb3tJ
ytxX7UFm1kOz8CrsGYjjGTn4Nr4a6rWFpPbY5MV0O762oVMBiWFADSZx0rXDgRW1
XjmcQL8U8ygcE2r2GLNuOPMHnCrckUF6lHclq3SG5e2LtcJAzCH2+gqEIlh8CZAk
p7SJBUDaPRE7OUGjkt4eR6gBxQsLfMU0vKpRoGb5rjUk6sN6PjuE248ZNX7CKo92
2BaUD8jkvUoJjExgA1+Tx9MKGVPcblz2uq+BBY2aa34K36nW3OANTj5gsH+PdAV9
B9j7HpuswSYUWiK0LOZIkoNkMESCNP4+PFqUYWuuWrgPq84dBHCza3VHwDr3ZCNk
ZEOyxvKm92O9bFhON6P7pTTAJME70msTFKyBkFjB511EZ/OEfee6dDxqO989xLLg
CGMlJ0MDegaOfUmTL0pcGM5oDke5eyZuW9x6VjB1EMUwu86pnxm052YCj9bfYT8L
+38sjVx7DLL2an4qAyQWeRnvcqWzong0WIhixOXFvGSkWRhGAsxsV+FBnHs/sHRD
blZRqDweEut2aBoORsRHnLNHOw4qD6aQqEf/uFDe3v+YfJYzNKzEHQ+bHgnMkhLV
puz1/vLFNhIN/7GSBXb3k2k8rYXIhmrII8fW5vnwiXgb1Ty62CMZGJsPvjXpLxU6
LwX8UPo9aCUIn7+D5LcGfajyoANB+Zz+lZE3x6pDfdLqVnrrHEqbNwLBVCiA0++s
8Rr4+xX+4FUjJWfLV4y/x9wfUe49VKpGShnX2+nl+qicOnVhJLptwln6Tb9QY5hh
mDgJIZqWhjOrgbdq/C3uBhyq6Ty3X3xdKrqXeinQ397hgd15eUnwyxzWt9m1fInA
n2aSDGjQjDylCidrogTVB2AY/7RY+URozE6Nxt3TXFmScE+fwOQy6fGnyfPwXm+r
HmN7ijeHbpaO5bxdGm/TCyhfylO8KW7hgSWmR//7V55QOGl0vglvANrJT3+US4Jd
i/z3al5XUV5UzYoVSP+i+hOM6p5etZP+7ZUzxRgax9YA5l2b8nGln0zXpooW7Iwp
zkB5869se0DIjlO0GaHpuHqvWVaAMy7J4DkoMZ7gxpwcKhxl2WTUuUUoRheZQgQe
wuMVfqVEVdTWkEuC9LTS74zk2/pQexXh+jbNnWH0x8ZmlT2BquZ6y/dy+uMjqFtB
dPRufoR+0L3zD9eu1KvrWM8+IeLCFsySVlim0B6d/0Z7yXbp1kMJzsMnUJpcci1V
/XlMecxfCsL4YsJFgavb3HlwETlIPDyaiy0HWnHzUyZwyyUXtQ6qkkJGGYYbkL6B
LVa/RyR2p63wGc65rPTm47J9NJSf2YSY7yL7nS/t0tqrAUI01t9KVK3KB8q2ruAP
v8wiNs4VRAb0YYb0+fz/GaI6JjnYs5/dDlr3ysfSSe2O1W28AlpyOzNq4NjsQ2Hp
gZsAJTZOKvGg2nU/98y7SeIfvRrIqqrFJ+dhh7B9rMdaicvDDUoB9IQllq23DUcp
6y/leoiRKHOzRhdxz9ym9BwjTo7EkSAz4ecxp7AKFFQkJUzMWfRdHYOL1QSezsM8
PJzw8lDWYyo3BcBbed9SLcIt/a2I52q8lhCYN47WpzkHtFzSUCizDkKkt/ksUSz6
2t7JfOzB5IveU+fRj4wkHAWb+TWVdRnG5nRHofZmWMqFpnh0dlibFLghQGu49H/y
sNTn8pvQupdsPjsctFVufFiPqDhmYwTZcdCw8Aeac0YsFpmr/0yK44T7P1XIXiTZ
Y4ovLQQvPuDdGZMRHMlZzJv3pcPMV6FesY+5VnW61c2IkzEPrFUc2ENnfNN5BWIP
RBkn9oChAGXEbgybKgmCyl5b+t9XcDX3O2IsXmqZS5hbVwHkHcfWpRMPQ5PkBtgz
FjcHaAzNVxkbOlrleN3RFzz3InCSKbWTBSwT4bq/HHg49zGm+mAz6iKzsQrQKPMS
sDplqxS7teG8p5IEOG+EPPxALggDWTd36vCWgK8/nHvlJ0EEF/mhAWgII2AxLMjJ
FTVKD/VulFeiKTj7wdU9PhmMkUt8pzOc7IDjlNQIEO6TCEEX6/lTciE7yzDB7hmz
LXYLUzhKAJhlc/YnocnqOXVkBrblmpqBG19/c4es3W/p9qRSWxRtp0u7Om56blTX
kofqQfF8u3zvWpdBVLh51RcVx8rQb1R+Jo0c6D7s7vZ8Ak2w5i+FU44A76O+/jIj
XK+pIzy8ORntPMLd8k3vdfEPIjx0QQHLcTS2be0bhMTQYi67awrlDSeyUwh/K1wP
valGeo4XIL29DvF6pDZ4pBXnnJ4DhRKd4abOGsbv4gWpeWchKyJq3pVAviqlOtPy
IkVziWfHbYP4vgVrww8gZWotJMTwg+sXgUJ44mYiUVYIdHvojoVcdsRhxYblitZT
RfpXKcuTWPjqmwlke6/QcAttQlbsKJ2upBNe/OKt0SufyiPJOUJcOhHLBheAXNUp
eYbuV+JWG5t3TomYA/9JEoWoDqrWMSCQb1G8ssjPQhrIMAdh7VQsU0LCk9aGwu14
Q0RLnJxf+xH8WkKI+E8+pxl+JJgBaPNAl78isS0YDrgQAmkJSAXB8Y9R6FF+pdaO
GopvYtJ6F1Gh1gxQ5PByMxBLeT/C6OQIaGSo1bDv3zoKEINMol9qnpEXhjzevpx4
AuDRS+UYlfdRBkcYKi3T40rrCzKyO/dOlbgbRazor3frYQjYksJYZyzOf+wb5f/o
Q3RPhlMF3ChjZ94SwqQ5HvnshnIA9+faH8phDy/pI+9eHAh4Q2YiTDbWovBr9A2s
nR8XdANbr2kH/Jj8uqEcGS7LLEp3SPUvkydHN2t+8VrjZvmO0GSroOXr7lGtkgNm
2ihgvKzV/mrKj/sDt6wYSrrp5XxzHnLEd6YxNnXviFZhXAy6Ou5yL7RPE8VV7BGY
pBVSCDmpyfVPy+21Soqw2Jisf4v75Rnqm+n7PmHiZxroBg5B0WCmxSd++XMTOYkF
Mq/HxAR3nZMUri190515QQL6CnUq6eDAun/1YxfafZNze14zCobTy4YDOf1ZOa3D
GQLjwCD/hpPmktxuWPfaUZ3k8dP1F+nuqgoM23jpTNjeNqj1Mt3mmmpNLFaJVN0B
RkVpMeQd16jwMGC4+MEihocwNO2UictFtSve/pVP3Z4nrMTJkXmjfuSfMJO4r9fe
A98BiN5i0parwCWrzrD01oO9uyNXWAX7EjviguLT9As8HcYiMpZiZdmpZ4us0+1Q
yqhbd3cbGfvn5nb6Py4u4QfTpyrJZlVFNlyySz7DLjlM4S8m19o5X2zG+VS74PuA
Z408eQkJGApH3rqcUd1VyeGRCLq4tcfRkeMfuxgFf6cyQm18EFPUnonkwRs9ipbU
86HYtJDsPczORQ57EkRYyKY0s1yN9T5qjL7+afuiTLUOZNrzWZanXenHmbDv+HgM
3qwqC6P4mDDYSfS1UtgvfAANE90Favoa8xWWIkh0lFI6j0xhh8SjYwLIIsRDCeMi
ECYEqa390X7t4wCrjqxP5pLrt6iFT0iISXbi2RgHpyecTEEoJiJYXl1Pqbl0a0ft
MbLMSOaw81YivpCQ2lmfMHzE+7GU+JThYfj2GauakmpLk9eqv+ks6ON2JBrwyr//
uLlZa1m5yoBBUJ5HdUibAw9IqIQkVnq3L4pDtAQtHrBPu3j20v/0U8+bEpHX7zWc
rybOar7r6mw3xembpz71ub4xFOvj7uwecUBt/8osky711uZRZpE8a14xnXjahzPD
SESJPlZbk7uKqD0pH9iF9f/EIlbwmm8Yv7bP9sZ1kB7owlEmAwIiXpQMnr6EFz6n
o/CZWEeGfnRLm7ZKYVNDH5CrqkWq1RRPZnZqux7HLda/LQWhhwI5CTIKT4i+rckI
42g5SznO5ncctMV37Ayfz5GqTjFwDHZ5uOu0Vdlv9qY46g/tc1TZ0KodZjYOi8PY
RbtxUuvo14fOeAkJMjN5oy12/nhPAtlPqTri2D6UZ9Gd+tISMmA64cR3ZCHF6o1x
X0ZvNunM+O5ghrYfYzbrvEGFWgIQhJLHQ3fgYa5Gveqa0/Ha2V1X33COeWQUsPxv
uI4dvzb+8R62cwTqvpCIRYZyHf5F2T0zKcGZgoUC1+MiAHD9QZ4QxoqFyrXKtof/
b80z5fyUsGV7vpIm6voH1KneVIKVU6VW2KhDFjIs4r4OJJiPFCrol+NYgrEBIDym
EBt7gbyMiJIk84swKfag6ZcVU7R5cve/T9mGwyrFRNtILDCCdQANHAgiDH4XzUWk
UBtHG58iDOWiJUnA+U4RfhZ/JR8a5mMiWKMELM8+u21NwQ9abM5lz/mXcFFkTJDG
HQwaOuIjMCz5B/Fb7AGBx+DuR52uQ/IXIkIIstq+MvqTDB9PpMQVVZK/0JvQzVK/
JOYRtwmiTPJHW5b3bJ4dexC1iRco32ZwRmIH+y4AGGux4VTMcmS238590iR7/20j
+KN+yeHxL7r77IJtdaYKTdGUTSPA5DGY1BUWCJLsHpfqt/6fbhPfExHLo+MqiAwv
OP8UguXU+upjaS8YfYgoeboIdF8DHzPEaVAfmzTebzUkcI5Fi2E3Ltmx8u8VIYQ+
I0Z0m1Zzq28RIRWSRdzysC7dZT7SIk2K5kvdcsaUB8bdOtIVL5zoqhDlIEmEefJo
pk5Rxua5JK2DA6YrIlKI6+OfyDFzPhS6ecLL3H3xL09BM1C8ThI7aJhYEAz2LhWK
cHLd/lDwUeY6w3RYkPJ9eTZz6pmMgCH6WeowZwYSNknPpj3jO3g8qxaox0TZZV4t
XqGFGpb43OjgwR7Tc5CVSXPw5ebmy8oWXbM4T4zkLsIdRq24THbLwqEx6R9JP/4z
iVspBvUD/xPiB9VToQh3I94cQzXyNPWtqBV9VozspXrsz9kBrg2TecJmPzx5ugu5
sF4NHxlW0YLgTKiYf2fSdc7B2q6cZ4V/eK+j9VDRn49QlSogNsKd2m5lynvx3R+Q
/u91cGsiah9v4gCjooBs/6skGXKVivICM2SUl+B7/4wfyK+6wrAzAH4areT7qAN8
+H/ZK3htnfrvfcasQsUsH3bBA37UgTnZD6pZ7sbAvj0S40gVcRtK3FfZQKIOry2N
BtQAkA7/JpBg/igsV6l2k/f+vqTnl5RqYbGGC5JmqenL0uhCEhfQnk8sWYYc3cY4
9ka2VlyKsI9o9QCa6wstayXbtBBNr2AdqA0vjMtM5AJ2pwgaUQf1ktPYV29m37rW
C6FrGQnfNEPaM909pqObodClGgl6rFPFjuXUurolpfVAuQDe9NC5iDYP54lSpbRM
caIvvSh9mZvlRQHaqGjMuIwaejlQz7kXE1tIh2YWrEFV4KXWpe3GYyZEQMwYdKri
OTLsKzwyy2rDnLBGwy3+hrjIxjxvi6hS961m9KK1mY2qZ61Z8sGWyZIBsY41AW4U
Tl5if5cz1uTE8ZRa2ihfWlfk4aUJjurX24GqNLQdiyalQQkgx7J+hlyfyqtZSgNB
QMtAhVzOr/FmoGNP2Wutx2Sum5HZ9Hj5xDNg8fDzfgP38JgpxBt+5mwOf/CqCvq+
Nd8orpzK5LcTIaq48HqYXaAU3BMaUahAXqgSloiqBnQBuVLKmQlQjQ+stPNJn8Ev
+ORwlWXG9kVFG6BW6YCLa2/E1/EloHdvAeuKfd0Cwz4ecPECvVWKyXcVo5bRJeCm
6xmxgowPXG+Ab29HusgBef8v47RPlNC4c7I6NdUn7We5bSNlBke/i0HsXR5yECZO
ToKXs//8wdGGq1eoNTU8Wy8OC5fPELsSu6iIekwz16uutY4jMyxZt1Tyi34P6F35
f2MdZ5l4xNcMC7AnxyafkEwUM3bXnBUnFjf3AulcPS+dJNWgo+bilcR11w55XmlS
vYj1KWek6U+957c/g3RjL2YlkIIYDlJ8ifCy9GT+KOXjGH8SdPrsxQERsFPXJPAN
gn6vZDIgQLrXOJnMFGgIMYeDKoKEb02MbI6sVMunGRX8DMprVWPA06PWe2uvFz+4
bMxfBo/PhzeYF/3Iq9vWe3ay/KPp7ullQnmWJHpp2NcvgqEtX28F4QEJLKLlOEV8
CmZ/nfm4+k7KiF73RyQkFtmSNUmaZgXgPfNdnRHNLrbe7nvSVoJzI8A/2nDuji7W
VBtWevMlBGf0UErcbeFr2DACFZEOSW7OUPkFl1zjM5cHEMzjMh8SHcqwKukFb/cC
xWlsDIsqPXpqeEEPSUecgz9/WKrezrpSvpAA7r+XE2Sb04a3A7jP4JY5SQ9vCL5s
cIulOxuYn2+xI7DWQJP1zpDX8SufTL8htQy+MwRPLk8fVFfUKQCaORu3ynbJUzCv
8k/PwJF20u0iDfrI3zuoiHKlS77LnYcLdLIu4dZcyrzNtU/UcvZCfjKANLR4KvWP
/8Yt3tUKHd7It06vKF9hPCqD6w12RNsVUijt8Xy/BgPWEfmBvrr6C35dgJTtQzDf
ozrvQaSCnzVyvYAePjI4RWDVUp9VY6+rCGW8VlcjJiHWZpwMyIeLrzYbxVXVo61p
pFh/PR9xPOicJyM9eU7wyvffUAxwCOBQjIBmFSQKFHN/+5LOd7yEgiJ2Kti77YZb
TjTiGI4bCccZhND3Xw/N4NBIRJGPfG3b9L2Mt6MwZRntFnDN3iSscCKwrrX3CrSH
m+PTO+NdT3PM57/UfuHFwF8vzQJ2DU80SyPb7jAIR3CXmDiZAQPQEw7ltV4eESP+
E9BofP9SUQy7nAcfXmalr+uT6dsU+bRNl7YZKwTDG5f2Bo2xm3oycdUk+tdOGJvb
v7NHLlPQZL5XAz94hp7HXSQhC2DBNeXq5ACJ5DknGRBn4lDeESCIEWBoWCof2ldX
rMepk5wbr0/+UHG62rUno/ILhfPd1GCn8lI9cCE4DuAHs+aJN0lU5/2Hocrq35+d
FIf+u2UZIfg92BVRHZ9YI0/1bCcyH4Vo0KzkfaxLUAFAKGMz/w6IlhBksKJVDuh5
2/jjOiWaT4Hq8G4Es8+rr2oacstRRK2OzpFmJRHFad3srX3fevCpns7g1LEaN3uG
pIKvs8fv/CfG8KAPL6Svf5sdSs+BvgG7hHsp/7a/rqVZJeC875a2FSBKbO4AGQwg
5cXVau+xzcDjt/c6U7IkLXl25ZE+LTP9NDyqHzFHz84P/IGJMqEkNfCNqNoKbFNB
YN2+3AsMgkG1Wdnn9YfchcroC5HshYBr2+0sp9R62VV6l9zBK1YiP/UOlFd7c6et
vTnLZX91nsmHAmtlo504xzWMhhu4wWvrR5HPJLn1pIkPpLhDY0CSVcH/pamhlIXp
7sdx23U285kMOsoqTtgnakrAsqrsMEzYZRtg2kfNt+K1+x9a88RYM/37x6gCdqGu
+f00Bu0zLKsICjs0F6l9FH6U35Xtyid9ClwA3tkt2I9WfQeo3yBP4ZnlzUkurfnE
37Petmi3fvCl5gOn85/Ewp0Qx1Y3T3LXg90KmITi9PIu1cENc3JSMhc6ZmeD8bNP
+foVY27iACEje2Q/tU+XYA1vM0/+yBX4pz3+cI3jBhYIyToqJTAMFlF+me1ZKc7+
gbygTM36pMfFTlhiIYVsg+Z7CWw5K5p5H6tNk65jprjAKvvp9T6CRjrRwfq9auOJ
5uSkwDlq+5YZFrttwxvrOoHoiI0Wcgpcia5Byso8+RevfWNu9pX9OOYcjMALoR9J
KwQmhhPkvnuggI3Lu1nlQOcZyWJ127nWA4WMsUb6STWhBfikOp3McqxNFXhDg1fu
acCrgl9miydBdPkbzDpsFlDbnG55Zsmv50Ky+cowWKCY4wmIlc2kx9bsPTSRdtVb
P1kHXcTjigxqz/+iVx7YcC+lYh1J/DpqnRPTlMQ7ztEufyuZPM0OjAdd42En0h0k
gLXquG5JlAXEafSHQgBTCJSswPWIu6oZBZDvDVxsgFMFwBlfzhHQaXd5j9yHQkJn
rdj3tbLbYmtmaQZ0o60WDR3jRW34t8tthggg1wR0TucyDwsguixzUrGNAQjcKqWT
u9pBiJhmoINv0eGQzYxVyaT7HF+lkAag2afftgVGUYRUXUm7AN4GMS9ijv0Ap2LQ
uxDexH7v081kAB/q5qN5UOva3K9NaOEkg85fymhl+FSW1wjzdIUyD3P9FGislP0i
FFK/XvOYRCpSCXmX08wYSbIhjiFsLudG8mNibZ3zvNMBUlvmOqdoayC7N9pVOsLz
OoDF6P1ep9XuK5IM2oRDwapajNO5pNND5DaIsSJBsedNdFe9tFjbdRr5EQ8nSQH9
fohckEg9Ou7csvKRIvtYa2JAe8QdB4QbO+C1c1RAgxJUYOZ6TBls0dF4RHjS4DuB
Jwv5HQtBtDsm8WSkYU6wGHGaO1iNPiUKp0unk2MCGq7IZPXVAs6ARxKFM7G40WAy
V2gBdpCZHA5YPFO2R6YB9qqbjh/PaIdSbY1iXI2pMFfGX4VKuGAFt7N940YMXX7c
JggyW7FzjlRCsOgfPrxFojfdpDGJcAQpvBTW1+vV83IIPV0dPNkCpDIvQYA40bMR
UQQEbnFuJocHF32+1ftCm6GDJRnL5tHoLBJqnEiNL7VihZzu2H4xqYCSewmuIU3L
ruytFOFdGkdjB9bMlXc6zyoLbBMNc3UvepMw9vJibrwsqVg1V2wp2hplMOhyOb1q
bz8aHN2GxTGyalBAE2xsWm9FYepZmL4u0o4CjhZfeDy5GVbXIYNbxe/xPW8UqFhF
0LlZ7PSFMWwoU0EtnGSK/j5dK2UGEG71yJcxQhDYuVePa5Mtt/1kLfJ/8ucSx9E/
0QZSHMsQ7kq07JxElkNo53xlOYOvG6t+G/uVKK/LfDRbRCQQBPpIUVJ4T52SVbPa
pIw6VJm3tdrC/cR78b95Vfxq0SxEsieDsWwICVFtq9AZReqheR0V5zqtQlP1NZ0m
3kq7SL47y7DXyPKSQLKUgRwPvE9eVCmr77w6f1OGV0vnnezIis+1LmN6LsjD1HrQ
X/K3ZbzvJ0WYoN5aIF0ApjWfVjPC4JzrJBWZ4aNDUT23rVENB3GQlllGcVWZ7iA5
XsnIqsj9YGS3foZDZ6pVVcNFwS6umTmdTsmT3O50KVXwtNqrI5snUXXy3Tsj1mO5
DGZx6G5JYpQxnpqIBS8uNyIPn89bQNd2adq6Cc8UVtWE//yfZCkyFCKBmuOR4yyh
+uhb9cAjTWey4jNBkUkBq0CNG+G0/yHUOuLBiDKdePZiobkveCieRK0UqTP5wQ0y
ewNFK/4OK57YNCaGmc63ZW+3QPIyUJ3lXi8fJjDb5kgCJ/rB+F9GsSzfQ0DDWHo+
BRIMrkRlaWcSo390VbHlo28SXdkUSHpVCpKWTnh0smmcLwSW6pokycOgj3k1vYL0
bzhNDTHhESBkk3+p3QFsbT34i7noGb9ZEb6ow8rabw8bBQdrps35FAUNZqM5OSzv
2LAT+URBQc4eGVrw3PeFrhkpEiIg5EaxYdo0EfjCoarhrAnH59DFpG85EXSVV+cl
qaXdS4Eje9/KEK6AU5ND3H3Iju1AdSubn7RRKsORKXBBe6oxiOL1UlkO37CRypNj
VhTV0RXFrcElt0z7Uiws9HSyAWhSD/UyT/HMbzEnoY4WWdPEtwfsgY0GqOuaOTAW
B4bsFy+9DJBDWK4xY9seuVKdT7k5Y3vy6q2YUmXvyUHY2r+lXeGtMKZwHaH4q3Jb
ltWJ4D07nZaqLmbTyCpj8Wjk8knvz61Jkweqm4xqigXAnN1fJkU+8VLA0v6pwDhv
zM9iJwBg7DILyN0dLTLuYIuB5MLj0Cml4ba73I1qFfu7krSyxLhywVJWLUMJSoqh
du6ZOHNvsMp2a7Vcv9qbCZM9AUh+NTrqRfY+/QOFJm0pOMwt6ni36XymJ5ZVS5KP
gtPijvaV1WIk0UEn/07OGGy4MNVTBZUNhAKNCcl86TbCW3fK5spFeHIMteCS+wU1
GF2/rNS+hcTK4DFy7ubiU6+tRl010AdGchb7fa2F02ARMusA/11fyKxIDs6dwxbS
P85dM8DZC3xNaY3pgR9X7E1YlG+khFiEqcy/iXAA3IMWTnPw6d+3Jgxt1HKERVZ8
ZDJAD925lMwS+j/mvdPVeClkVqtGzD+l1XZ/2XtKu6doOTVEINWvgroZKj1+blNx
mPztEM7TuQcIiw2E62prOPLGLJcylSVNKdxYl52vzdRPD7XeXtly5aGBrR2S9F8X
1hslRgIbmgEl5EyZSEPJWy1sM5MZ3OQk17tC5WLnJqc9L3ouoW6UFFu1yd5i3Uns
tOwN5DNtY1QjCU+aMdFtklI3s7dQmH1lMB14C+yXhyqMVny0Z+xBXZ4UOmsPuSKB
zd5vfYhR8g+WKQ43OYkNBiY0KRvTxWSj/L7dYnPNdqm6BkocIO0XbyN8XAKydxYB
OZXG6zMNM6V+uYLcx49BX7bD8L2HI21rQRRGtpro+nuYrP+mTZ/8N5kmb7YB/lgD
DDAgrL7HVkUyvE85f7r2ije71iq0t5qcYLSsnZJyUK3rgWszI7Sx8IIKtM8c/26a
jUPPvrwM3kUPbfIcBMGnfC35ctMzh5uzJIDs9kknnAeTfxKLgdr4LYO5UIM0ky1B
vKNDJfeVX2kkBk+V7FoylgjMujY+BIBJ3UH2PdoPKUyD6pkmjcrxzEC7E2BKOH1P
mgRv20ubFgxbfIwd6DPlfnPfW1OSMEivFu8SG7yM6uRSIIs0CUpi82y16ps3fXcI
0ea9GIlLZ32a8FBvb9oAt2hMlKOENC2COtPa6az41H0jhpNqDZUGQYy3T2rc4LS5
016lG9pS/WgUivEUdZGSisYMkTm8JfHjNVIgBCbWXOk0aNPLkxs/+0Cia9yuZZ0M
fbvtmyJpK90nzYBeqSI5HiCOr3X8uJRo9ZLtRr06ft8a402XhCFqYd7ibADj6nhN
yPJa4Z6nmc0bI71cOjjaP7rSTg+iQ0K+WrMMjshB0R2cAWasmmUPsfnYNNkZqo4g
zuGxucmL0AyezK3YUVs+OxMdte7O0tasWe7KvCYkY2hNS3BEhDVakEosi1KdfAQU
wfRoLCZxXSgYFjhpxQovCzr2gr+w+T6gx+v6XXJpSv4eEtMHVQO35ri6sNuIqHzL
OLkKwuRAOFM4WL/1ZqIkNpFo9GBIp2+Q8aZNwKnG6aonn+gC4MTvaOr3uCh9JDkI
ClSIi+HFEHH/f7VSCuD0349s81uoWjuu3DsQbzs/HylpsFnxtaJqGuNnSGqXDVCZ
y0w/PV4p7IH7ZkC1Mwr8atip9loUiPPl+bsnrEimC3QeD29YZrn4KKAWKTo/2GCo
Izrla/8pWB700AgEuItbFl1PxtLfA8NqPfvZqvygSjIOqcjGe2J69m7iNdzuNOgQ
iJmhkr5G+yBOdePccGdWcZPRmjOMGbaTKigBrcuCc6MZ5DdlyHqD/Ve2w7xmslHq
YsslSbx7xExy47X5lDLJngSDj41I/9Fo0Y6Xc5w1HB1sylpO1ZZxPuSC9WdK2E+X
QeAn1vcH3CXSxKvBPrylgP6zIvuoNk0nUpwBq5PVqcPj1u8OYHBShqyQvuFUbbmG
M59zOo6I6AhR+WbfyXsftZOM/LH0E5uJR397v63zKAspVptFLuwP4vR0FG4Z/d+p
Y8FMA5TvUd53LySU4tbOvWjPc6P041neMOMN2ONOyCq2MGuywQuuDVFREgAzJpmB
2J6EsMq/lVD+iArqS/0KMerMSLfeD9FLBgsOrtXd0zoafVR8m7gSWIyDQ+FH3HT4
Ga3a2TRrIUF4VyER9L1r72eIdDT0dYEErDmcPqf7LNsryw2hoP6g6M+KofUQdyRu
JvRlJmB48YBBo2SaTlNsnGVF9nmLkHbiDIlmpdBilxSiXKRlfOnnne/CAEHcdYXW
DJtd1VxAHGIoxWCWbtDGcvxfbZsYyjjR8ONwW5rN4NWnHZUFsMN28hsDqYKMHhEM
PTGhP1tCYQFyi29bfD/rTEUwoMOCEmzCFN7rWFTU4/D4uHAlxR/ep3JZEaQGAjb1
ueqhaaf8xH+ko5z/0wP8qxzS9SUPP9qVU8TFaL4LVdReUzLywAJqFov0EIA6JwSK
CJmfw0sl1CesNrqsQTA56Q4qr0K/dsA/bKaG25wAwuS8rOblDAQU01oUkPrg+ggJ
luuIUOpZga2J+KHEr70TxbNHVN2+srn0Wk9MburGRNe9M+pr4jU9etGJ1ERke4lJ
Rdeb5W/05uSLRM3GTFmAoffiAGkZ9RmAoogDAmisptCUMSBjvcnXbaImKGI2cqCw
Qvuf0i4Zy2e8bmVf/118HmKj9DLQD2HuDHVwhpUSH54D+/ZMRttJAjmH631RRtm3
tpmR1UHEVO7d5plgCr9BD0E8QefpCgsRbaZanqWiGEF+AY1MAi75p2CnDJDn3/d0
mXlL6/hQ7LLef2yd6b/EIMcOCjCtxkh7bMOD5Q5HDo+ww5tEDw1XXRuR/VqC4hHW
IDIHcsVG82ltZEgU/sfUOWxZjZ5MLblJW456tAdMrmFAtV1KtqA8kByzBT/qS88W
Rp0UmAawhfDXvpqYR069lUFdM42UanhcanwkTTRZPD5Ag1FkctB+TFjTgsZM/Yu0
EqT1XGx0iBBrwEb2cVcIZqsaRKOp6uoMyzn8w4286bAsFwn5cKBZXo5OnK7veii+
U0UZvC8u5489ODNmW5NUeiwTq+hsqJ8tnx4n5weZGVWoQX7pndEUpcW3i5VqPXTI
EwiYmOht7D5ddI68BAVuXRM1DEg5e6HKUgvlUDA2DLVHrwRpTYwGE0ecFUMm/y/k
Zp1xgemrqDSckOLu3kwBgFtqA2ZpTI672hrvxq5Du1Hcp7WafvdliIKHqL2MMT4o
GYwjQYrVtWV60zQwTXtalJe6hVeU4lv782Kya/swA0ooNlaTInc8SEpbcsa1k1+z
6d2AobWeY9JY7UkBe2jcFSHgOqjkKuXauE3IOokio07dhQ2+2B0L3NdXZlvFg/fT
sSmN5VizrQxrDH73ROC9lZaTIru/U4J9ZNpb6sYOiz402WiVfELdCBkIZKDhzSoj
fJl1xz6VJp1M5JB1gnd3nypfPYu82TlOEsXSykSw86TWQIyugR5M2/E00nOqhTDc
SAmjTmu003Bwxb0ziqGF83BpC767zdb2hpgO4Ww7kJwxrb8tyl0jYz2HlrtzWGR+
vZzu9Uhi+d7sgHBwYAknau2GueCqUE7vK6h4RWzFI0JLei6LUYpv4AxGLhsKC4YQ
dxQLehH1Vke8ZSzI5YAB0Ej7sOblack7H3dLCu0V3Ie6D8zYuzfTMZcYPKS4HtGm
Z70np6s/9ysQ+84qKVJ5lQXxKGOb3fiVsw+jQv4gK/JGpGGb6jBpzVfYvCYMB4UL
QQjIcZsqEkF5SmwMEFxwpY7d7ThCmbomkzcY42heBFD9H3FkkpdJyvVdsxzaQcK1
NCLx3DgIuVYxFuytYtwGK7mHMXkkbi0iczaQQyHyuIZPpP5x8HH279vBBlaUhGQd
AMPRdJfztn+Hp/i3mzsmYphF/PoCxq88iFtUC5+7jaYSuIQkxLLZaieR7WauzYOI
RFS710jOU7e8gCOwU/XgrNJ3zsoP0hEPIhxz5ETLD58k8wWAb6qsdACMslbk1uiE
icNLkS7G3+xkIp1h1kVE7GQ8b1JTv19lzm3vTU7KqvZBhb3lDkrFZHxmXduW6fAh
u244Xom3w3wYtj42WxCHZQN/M6FDoQK+3MkiemEg+eQiDjmcFEoI+mbJatfIVCQD
pqo5ov9c2PGZC3tPGpsz3w720svK+M6g1hBecfRX0NXw3FyBTHphyZaolrnTilnJ
lwGUnioplL84G+hRQUPwQXFaxE03lv3S8ebxQ0esL+KZ5IhlCL1MEiAFPD2CVoJS
LlQIYIslEOsIegRcURRJHDLK9dllLUcx40dgVPt+E4T2JC3aB1G7eK3ov4wlbntm
27+kBrlSoTLkM/uyjoktmj6E/hOkDNoj0T6PUMzMbZEblVtxyLNFRQWb6qakUdn2
7JKOiqiJp0b5cPxnmr8AAUZngmv5wT8Ufg8hEPndtAQaJAXLxbhHOGVlPvf4n2b7
fuRInYej6lgtFjyIUNxBCag4wH8EOQFBRu5hHUwBcdd2V4TdIcfC3D52mX31gMX8
hLdyMvtVY0+RYtBB2QXx5zILjw/p18KfjnMG2mQkhcs9fgdyFQVs4p8xHf4jbm+k
xm7JqnlFWbw8vxIRO/UrabI/7BRcT+YQTj4Tf3Aa5d2hk17vrP5+0k17q2Dd+Hhs
+Y3kkm/T1tQIs1l1ajNMuJ2nELBrZx8OA/u6NWJbjHj+Y9xvbupt501gamiUWQuY
SbCNB/U8Oo6kqDWNkjOT6pkZz5sjA1fWppqMDf8mDfl2br8WM/6zWjU2ctx7QMRc
UxwEsNW8SjrN5qloYnOn0D2bH80pfxZvsIl4fLreKsLkrhxqVNB1DHHN03D+Yzvb
FK8Hm8fZVDuX2PKdtyuq85FbcoXhBJTniqXcYwtwk9POJbTw5tNwl9kAea//S9tp
D1CuUK3dOmz1oxzrFhlWdXklQ4j70Bll6qYXoBC5q2KcJ9mHnlarqVMymaN3CgPP
1kMKlnz0xOZ+qpCMguFHcm6uXkYgBZecb6pW30Wm9tsZ4mVp5Dq2HO+LHskDEP++
NWKRfh2v7+Ew1vZcQ9CyuoN8EDVHLIGzdx35rZAApCq7iGj5DjnA8+i66EbQBPjy
7FAfytt0sacmOHH7R1snxZUE1SIYg/eiGezeO2J2DVBUkfxtyWNvEwlsbkUzN+4m
ZZU4v2UToigLK5WLONK26fqT0+tAZwizv+GxP6A5BqyaN5LEfZlTJMKFlQwnaNHz
2C5kcdaFZCuDYeCqshRvjrnyJxJjCETO9TbHi2+fMiPa24l0bIWwiqJSqC4Im2BM
D8mrcdMjIHr+ulauMIJjuMltmG8zX/JVCntlN25R7VLDg3xZOY8Bd0Xw3OtFg3u3
7rOADOOOGVuV5U+Wn6hBgjSJkZX3zFzDv2dqv8QuGGpoLk3jtFWCR30seSo7iN1p
yuIzR8w6/D/Gfk/gKneaTclZFWSfcsGPR5SHNrQ2AbtNyVtFGQejekcJxAZ13qWq
1EXa98lFB8LFxGPAJ/nBYHu770qwAWA3oNimmDIn+skhz+lUSqd+PbbAom46MvSY
j6/9AdfOlk6DczdJHOa62P1aCveWgMfqmd0UOvDRAP5XklcA0NWxVMERCzcOY+W2
5QwNr0Y7cW5P4CRWKPKukJ7XY+EK+9tZv97h5PO5quJ6Xwn9vlBQ7JhyUo49iu5t
eKVyk+L22ycLDVS2PtTQG1aPvoOEtD0JNk3QZG+ePHZmZSdApspacUJm+QErKPVY
JSJ5NBIBs7yiylZPUgKBx3dv1x8x/6Q2VLFQYRsotQMap6LiRkJ+8TJkpwAxx1zu
8V1rBVpGl/Q14y9XCcLtIbkmFjpgP5TezHLMiwLrYNCXDe1Z0s+u3gUul3yc7N/m
b3z+yQZE1YB5pON5EJDKaVxUi96H4UUvZjsX4PM/iayweBKaLp/Fc9mkBKJHQ4kj
55fkYm9EpdFsPS1zIlCOb4PTqDygfo5NRyeDEgOs1kScuskjePfe7c5TknrIJTgd
Fk+Z+zcB36VPM0X1Oj0OezoVMP6Ssu0TQ66rD5AAFqwK2gDTq6Zp+7i4Lt7V22ND
8gbBcXEfPnxLsj76LsjiB1w0xo7htRon+u5iTFEoCnLLxXTurAWbGDjgYjh/yDNE
gPeoZT1FFizChXtn5KbuAOM8dCkOzLbH6TXmSUUySyCV/lUdX1av40oZbMNgjt1s
xv8HiDEw4bNhLwN/oS6PFVWid86JWoInmhrbM7FK6r6eqG2Dq8t/pCgpSQPV+llv
mtoA6k5vDHjV5H05pYZ1Z9sGY9gSgizSDY8GIOUpu3C5Oj7L4qNewjmMP0IYIpC0
SFNsm7d9rPdEgVhWoSFRGn37IT9lDo4L29zH5ZOtzzbNtZfMucYcdxaBIoAs3s7y
snhMutzTwlZgTr2twwG8NdZFs4KoaYoUvzCUCOOOiWI78VsLGXRypudovQArisRI
vEADBD4NIxlJ8Wc9Ar5FdacX9zg8HqQSy+w1wrQ9TvzVva/NJBxwFTq0TDp1ykh9
usjtZsI9N/vKQErdQchSWB3tpS0xI00iCTPL2XjCJ4aoj0jvr2W46h4KVHbZ3btQ
LJlsNCAiPEvVqDWCn4DNdljFIQ5TZMtQ+n5WEP3CmzJWbLXBJc/HnBE5oqwhOg0K
fJuhbXPMp0tSKobQSMsPm6cqtz2/KS1ojdmx836Y4tQ7/jgbrYW2UV9NlzR5Gkle
CO4UNWk2cV5L/VofcO5rDkuhOBwX3sMjHrcpkwWojWmk0ekp17u7jT5i85VPA8GJ
47mrm5GnOqTupuIGDgIqAu+SJocfgIXlHgrapCBhpR35jU3VsNytG6+G6B2ttIUS
P5xsAAatVX+PwzSOjH8oS5atABJ526yXsEdbQwLTavyrRll+CFXjFCou5wDIRhjb
7EKcsEyVMwmLkkrzpJcOYtcpxZ0ZafIHhC/ZDY+1GWYTTR47EIPmfmYT07R4MI6p
8gDXHo6r1cHhT3pURTVPJFxiBvPdQafaI+0e53DK7Oqxk54rep2tXYjE4aET/FoM
E+MeDMoXYMR0eYO5ZYJ9E/ko2N4e8ZU77UgqsulNsWxauCZ8XUamY6QZAlXR0VZG
lHhIwxf+h6WwHEquFXM/QBjz4App70OPscx9u4T8bXM4HbUlpCRiDx82iIPGfRVT
BPzUOsJJsMKW/TX3/OnGLfJtRq6XoKFHqGkPm7QkMU0cF15YVXfnm8Gs146krJ7t
ib8ar3gmRe4htVYekVC5tjGrwh7PwopoJuG7qYyy/jeo0CAsHXXRunFEKk85HJ0G
Ja49uY82VUofukPVH+5eE0eb1xjJYdJ2ePC/sXejowzHabH7Til316kifAqgq+U/
L66O6drZcdFj6qIjwskC+NlqfSIsgXaG25qxLjU5s64M3h6BOtUI+F+PlwpWO3Bg
ttfBgWSTogUHm72RrfB4TvleXV+AJr1Kfmoxh297gzicw7APk/p1sUMrshri8Tq9
xBt/nVi+5rN9HtSomiN5xdOJWx9FJOhj5rfzYoNaZ7yVMuZXj3YH1dENErknDIvZ
iIKoLXeqXZLpMvA9KhGIowThGJqdpXeFWpx0psI0WrQgO2PuPU/3uLhYeqLY1DL5
7zRbNC15IaPJmEPSx4MuL3zqw3vOlNOpPOPCQZCXjqW32xd9VlRoo9AQx10TfOkK
biqpQcgp4vqPb7+3H8Mra/hMre9OKjbcE6lk/q3oobJ1QtkycgRg41ZkINh+Ct/x
1G8ocbozLfBJn+Ckr6l+D1x0AOxmdlN7mW/krNRuFdvC1ucHw3tTSfv2G1gzjSsq
xj5dbvcTh/OkCqwSUs2Op0yUpPlysCSXAcgwtI6LkzpBV0jlB62ei2+U+J6/rmoP
SH2Gjsxi+S09q2irLV7VkOSKvcN6oM0j9poo8EAfds9OY3bs1gNEmW2hfYvbkIuE
5sUNyKzM4875+G8Yj/GuI2+b3nFGSXTGUnary3V+0umm6xuWpMkZ2NimPhWRWPCd
wloYt01u4z+qEauzrsnKDDk7DSjauCUAK/eJ7Izt/7Z4lbvzsIyVm4vJqxRB4JV+
1dZT5Xi+48WN3AvnpCGreU6MlLkzRC1hHgtztbFj5LM7VtwiX72YhVvBxfZma7l8
SIU0YWf5FFc+bnuDlDiGROkDAyWk+ChoQmEuduL14uxLeqn+ogFFG9xzLyvBmdZQ
58qjlQbOdC8Zm0QXfqkB10I9HN7YWc1JHCgpVmXePSnpn4biWyzVmDgCOWwax5gn
S1XnemIitzkUX6YCqy1qgmt+qBFVnCOY9JLU1qvuGRzCBS//vdxgduXHWemq1uOF
OzUTiBgnu+AJDDe0do5R9XXSR9IUwok9slTpQ3i/eIbgR1+WXxurdC5O6hkczBRo
5u7lFDHOK7TKdiL0K6DTg+LCjZughhYXlUQ5a4x/OIrDResQCF9b3Z2uRnX6In6t
waWY3dXDzn5ryUQwKL+RNZStMOFhHVTIALsxFcsL1R8j3vwPzxVvDF0EgPx7GVBO
zhgk7WzcIJKPvSypV/CYtMFN/vHGRA1rw6DwffSFUO23IWv4RjerSSt7XvhbQ1b9
1S2wKfHsCgxGSKKA6yMh7JTvoeoGxmW19wDnOGqWyPl1VFRYU7+Bg4mn55+TOEWi
XKftxwSXoRL6+R5jn4n9tw/CSdyeaQGO/94Kjp1T7w830sfs46siQMBbYUtkge8t
9Rn/GFAW26Kg7/AjJIQPf5aRC+y/j0m25TlHx83RD/uc3vAx48RNh6HaJ3aB9V4P
UPj1IFJ9owaiZZqbXI8V3XnIGQHRpveF9KI4XkruyE7BU9C7KPr0fm/Xwk+8ELhd
8acnw6Vo3QSGjEs+vgfQJpdYk2kSvF6lcXuJ2gv2R0GH3zP2NZVPNRc/W+v6KMnu
ZoNci2qnn1l/yhi9ttGULuVSepeXWa20xn+u1vn/og0uQCOKp2oQJ2Txi5PAHKtK
XnHRX1GdkQ3Qdz26XVlR5oIefA2PqIsAPw5ELg1gsZF0tYzyDLYqG+/ubKP8SYZD
5S0IbzCbam7AF641f8aeP72LudCtanOM8mOCY5cFhtnjrawPy2y0A07bN0WXZIgA
57/xsd2PObIQJPe8kbuEtEHWP6V+gVhtL/iaI5rzAqV66MytL4wSSC/j1Kg2/BQB
ez4RnHEx9D1rWHUtGSB+V7HupZ5N9Zv78s/htQDWvHt2q9TGsHjFJpAC5Y0+O8aN
T64OxMNPKEJ7W0V8B2Oy5F3fKVVvrrl2/y6fuu0u3YZ+U7bjWUTfxBGPOE0OBNdw
VWEy/YPXkhijvEzqGRQmYfBOMbV7s8uYiNnaOe5j9hF29oBJECg8/9m3vB/x8cMY
V/8klGIwpta1caYxJpH7lwdRxv8gPq7lGoaM16mlvxUPmr/feYIJ330iMuiDPHRh
cDferkSyS82KxCbd3nS7AHfye2DtaQ/LAIIrDZd7FS0tOT/oX3DgYSePazMkALTz
IhE6CnFkAox8axTmiMiVhFsvSLxfbdLxAxkdjnistETJG2M+Dc6A/NR+yPt8HIDy
Z0zlowehaiQ/36V7Bp572kWXDIuYr8Yrmwb5d06r1/g8h2e5/MqERP8qdtDSqzGD
kRM9MvLdy1RO2nMoJ/iLEWXZYqIVmZEgdsCo+seo6p7WPdCWHw48NrH2s3SP5AEi
GaF745cvHaAzY8fgMXqCsArKCjpEiI6pwxFvh5Un67MPZSRd8Honx9JEtq8y2bQ6
q8byX6zVIhCEznEo8jklcuSBWLFYLjceENT1Xe89jpb3qmZp8Q5/zSrwZi+4uWJ9
Qq6d4FZS0ySGnuGEwJSdkh/tPp28CE5oZqoIHufbJ46M5O0h5q6lhJjwmDrwTdXL
aw6BpvFOPkRPeYeYjVycnJHefM4wesN+FCnkD+JLERKMAg09wRJ43tFcyhShYj70
lRq2r1769nxtIPgJeMYkbVJLzVvU5tVbt+qHU57b6ZqUEzBtwFgmxNdunySFngH3
daaiP+hsSaj4jk5q1bEHHGzDQR7Pk1tTp4RwPSiUBAr+UQ6d7bz65S6wqHvtB3rR
SvzhLyRUtys2y34FgYEg7zLf6U/s2b7Uj0M1wwKJtcRv2il6VaFOOfer84fUj54f
lqXbXuKfeuEtscHq+vP56Bluc+nOw/SMYx7i7toyVijxmJGjUHQPvIIoFTBN3AsP
cJhmAYG9RqIZSOm30KgswfqCB/nHDMpFhwp1K2btj9ryPzbSijnot2wiV0D/N4lB
8WOA0zTgrTqdFByZrmWD22srQ2siKPvtKfllnnHe2XqmEH9HLUBCEgQZzZIlk4Kt
62ePSVSsZFMmsNdbs9e58IVZPE8/Qxxf6DRu1sN7rK+NJF0mS7IDyRlWrgDQxCBx
0GF1cRhHW6DZYANb3t0Xni6ljiZOABKIOZqrwZ3l7h6Isa1xV0gpFq3AMyx3jIr8
wWHz7pbpiEcAtr0l+t28DZWam7GbC2VdBYhyZPvYic1CepYcosC5WEKds40A5MWH
9t+zVrI7IZjgpcyh2fF8g7zEAtE3jKdtgC7fsvf1oqkBQL3OAiWQIdz6RaAmxKTn
X+EdXZuECCsMGGdwIBZg0hJ3h3GEaqK7GWQPEnqntBgRM24PF+a6paY7p+UxVq8K
7vb8m13ijVotLDI+qkHSkObo1ncDJRv4DMt4VRfJCBy26j9sle6MC8/bjnOwbCkv
BEmIVrbT8dFipFJHtwkoQ00waTMVHTWPcumYl9j4ery/rvi4HgZZTLW4guW1R2n/
DLClFWt+hwG9WdqvUKvJLhudf9GZncqFqsGBTXXhCGu4sFerqO0ypMPpS6ntjlQg
2LNRtoU38NzPvZFwSnepAmqxNSshPZTOrtcfaZ/PLmedrC/ZFA8NMPG9WfimdA23
2/Mc/jVNcukqZ2/PrIUlNtglAKg+s49nH8/lEa6Md3kZMkYVX7fKAI7sJH7IAm9t
LTnjbhUBuAlBSLbXHABFveayVbUAaSXaVSKChZyCz68Buj9y7kwStuBTuANDmWz8
bK+o5wtp34vS8qxbqMN74kFBda4Oanf2DJL0WH+cgbo1Ye6Y70hTgLq3Xo4Y8XHj
Twg8FFE2mnQt6GL5hmf4PwFzbMUeotAukSKR6ziJyK5U498ZfzmltID3L3thLmc8
SvmSI1CQGhswB2ArEQhIsQLk8ZlNF780HxGMMwYLBruT+EKuBXimd6gLd+j22eps
d7vf7IVVbuA7JyYlR8hS5rGNBEL7Hbn1bhVSfzlSchakLTG4wCdoKfugFPNBXIde
HCLNfz/II9XwO4TtiMFKOjy/w8flHnh2pAYxLX3luQzrWcNV/K2+5PbUC7+K13S+
qSoatIkVNgMon685b8NVUpXQZe+c1m9/T0K3/9K5U1ZAuDk8PDYARjgd09rEjC9r
9IPvbNtRdY+fDU6F5URRFNpQoYaCQ25Aq2mhzGMC7c/B6HgmRDBgTa9rATacMbo1
MIS2eXBBeJhAexWap3ZUCX2SDsAgfh4xc5/i6Yy/nlrmKWXBKGtG/DPWWXrcp1Yk
rsmGpQSSXm1ML2JxETxaL0VK4gF5036nvYOBGKfUYyd3Z2lsZR58cZ7C8D2LTrpb
S8ZBCrRsRf6ujaQy2FsfYu+SSLi6qeFEgyWIdkzLigvX9nSg4osPB56UOuwhlUPb
OlbKTtaB+JprNIQj7e5EfEBvRhOlq6Sr5NEpqAUHahC7mTybTIwwfuIZHfN5qNCT
8L7qaxehMucYndvgcKZGVUHzr0fQFcJQhMUEA2bliJm1+1BnKrZliv5f2rJcZXeT
ZVZ1a0aOdXxnjzq34Etwo63GRZDUoPleCHg4miOGDGtEpzEDX50esTjC5FOUy3XK
+g3rN7iFw11UQsofoKV93cxJfFh+oB6x6nQ8YYwbOrc+vU1JTMti4q2IB7VuH4Dj
L31GlKuF5MlXpFLu3fuiA0QDke73o8OAyvhEtchYbDjeQ4+TJTIO5AaDltxFvHba
TAS3y5yLMvAa0t1ZGGZC0V/QW2x4e1M+zjjuBlQP8BuVyJiJGxZnfMWKb9NYIHWP
LZsrrVfcQkBSR53IUW4UOg7smhMJBWIXC4ktdMc+gKej1UagjEU/ZIC6DVElWDrr
P/p+VyEpYGpXNcn2w0c5GE/l1OAki4Nr7PO94X9GdgNNcNZ2CXYVtlsYL1eXmKju
DE+uaDhYbPY7Ul9JSQ4TS8kBbC7mwtEUvgxmNdZRNkP3Nt6ETqF2pp+1LN3xtZ2P
SXUxiolW5GgbVIns12VA0M2BX3XSCLrgp6cu28yPesF91VIKOQAND2k+At19nvTt
R5er9Q6QYxY6LHJ8rs5+5SA2fpEApqPvzcdsM/j+Lz2jcaHnGX1br3k71syIi9a2
8fSuZY5Xq91zFOp+2vDA7ZmY8jlf5emqkmXzBJfiTd9rHLLEPLui8JsqTgxzfRJf
hzWnu/zy47Bosw/lrEHdggPD3eRMUW1U2zVpGt7g2BbH3Te/QpI0pFaTuQGg7ixD
t/FFM/ulcjFtU2e5P/Jq+2t+OBIWJ0yiOhVNAZFizyJURgwx3WMHPcBzirUBBOPu
t9gAgDB+GXEsJxZPek6nTadzKI1daKsMKYY5Z9I9/RL+2bP/3/OyCNDJ9R15gHDl
z/YfnZs03sE9ca50tiy2oUou++BVDhrZKYzfcatcs2xoN+DBYsuBcvqtqbAzbzdT
qgUAFr0IY9JgWLzWEFsD+cbduZZ+zxzSwAnbHBTRvwuAUKsCLtxR5uAh4jj8lAtn
fV0B6kzs6wUFutCXIp2j44/5DbbcYxM6QZHSAR+cQva07MnwFgYcGjzFIoJfJXRt
zyK1ublywwSFjjaGHx5h6mp/XLT50UtySqezGxz06M3t/HS9HcDPyh4MpV9BVNsb
PbKCx6CyQhvmbAWEffHnz5naLbsD5GuU2wqEcK3uHspg52xbdekEwtKW1KHzF30t
XOgKkkxmWchoOq8/EdnERr1sllzmm9nghpL283GNFuGHcRrCO7ZYiv/XSialAae/
tzf/P4/uHC1Xkdnw+cv6CzgHYX+guXLYsdub8JL+9FVCbx+druaKEsmycfljsiUk
ruuDcJTER0TO9N5+ePfRmzXlhCw9ccsOlewDMWCbpw+D5juT27185K9YKzgCEylw
9IJItaZ9JOtJaQGHzw02Ah0kH+xfVEJW/u7talvmds+y6gz7lOhqgQEYSV5HjqrL
Exqn5i2W//PzZdyDVzUrxk3wzoRcRfODvw1K5PGHNDr2wxuQN4gY0EdVXnpb5NQv
5cQAovdf+cS7qCf9+q+w43L7Xa6LDnaeTZx9WmpQ5nv4rYwJr0NqiSIgzdhRG3dg
3EHSlykich+5W81ar2C8O8D6MlSMxHBlm+rvCnHwBmDblxV9dQf3JgHUIzqsH3I0
92ViXZb4AwoZ8h1Be6Wh0Bp2XRW3nhPbk2RknPVFWPfU6vb4Yf96urewtE76SQue
2imsDL3di2+BXGhe0f23u//UgbrM5p18dgo4VdjOYUIDXT53RRPXP0QIQ+i3wzsO
2N3p//5Z0o2WGGPqxWM9f2WhlTdP5REfSHZ7yf6N5QMoTZRroqMSIzZSzd5+YGMW
waaY0b66sIR60dR+T/H/qngxw3GfWefKYwNIZW3B1WrsI+bb9X2PI7CbLlpWa/W1
C2U40fyH3e1MkwT1nZAjl4Esip7/9UZZqXDPusweGGODg9G3/e/ouLkCqfWMmOz+
k/KIbjDKR8DfWXEqhm4AMBqt2xf134sFdIhFvWZrYYpAgnPb32zbqETNchIRworq
12TGZyM2IRJu2QRRBqWf+uFtjizYqtH4VHTWS/2pS6urLBGT9+A45Lz84YyWZYkd
tuNWIPwSR4tH4Y2/vOyDt9/v4Di2PXwrmN8FXzmPdpi+VEAMYzsZoNnTuOst0yDA
M2lXcAEPkizzVMf+Pde8OfN4BhEAWwYSIbzbpS01dffLi6dbheKGfGDMkrGWaSf8
OLaOn6iYsoUdrTPjOI5sae4653V0Dj/FtMdhbsZgkoufCgjRzOfrobhmefL7PR7w
w5Bn4tPNPIRJdwYGvJk1BV4e+FMCI6qtw80bHZcligT3s5e4yY7u8Hk55iTulWDE
zgSBNXv0LKpx+faEmgBNGHQeOfXl0UjYoq1IuDNO1KoqvZldZFGwkXMxXLbx9S5r
oHShsG+ZSyVO32B7dWvwpUZ4lDx1i5YnhG5ypAfDeh1K4FdA5oYv+unnYVR7aprq
zcB3TpqGngIWAHMD0kWuZ8KY++A6GFWpJEZU5RtTUvTrs3PSo/fALiWgx9Z9WUxL
ii1EQXyFv04Z4ojpaaumYu257qlcZSqW2uhTUDmy4ondChaeAN/nDYclC6yH3JMG
B/38mSReTkiQFr9lfQXo2NVwgNTVCI3Wm25I6XFvU/AHwROB58+XO2rtBNRqAktZ
T5upR9CaSGdQsAUKkBixDAfWgWGzar4k4zAqCTpntgBJ+s2WSw1kdZYKuaVFG6A7
nd7gxywvXEGOAwy5qGPmXxfCXCI+BMT3TF/X56wjJGe2jVwYgDh/O0QRjATDDLdS
oLZAklhQ/Gv03SY2eo5TnhDsozChJlnTrX2Z2LbmFf1lEWKNGVaAmFseESCbUfHv
1xh1bNVGGP3+NJSdARC9HW6C6jQCQ5MjsURZmkjdmK7O6IFHJSd9x1hJPwiHilEp
C7BC6VXWtxDf1NwjvpYWIOhEyFYFsU5jZjZ596NoVX5dI4wG5iNLdznNrRvY5GSY
Aud7JdXw1bT+UrEmz6HyJRigFv/zhYCh2YUNYWmOmLDdp702PXsCDLeElZig3An0
gRsHvyT0e33UxfychM1eqZrYdilOSA+yH6PAJfIoARzmSW10OwSz54PBXtBWvSZB
UGIp0ndxJYz2XvJrHPGorv8pWdrYiOJTJnbWjnRgcNrG7sIxQ/rYiKJG+KwW/Rh+
T2pUx9YDoupaviKEkdoWCq7I63jHZj3/HKDHNQvagRsS1xK0Yn6vMZAeiRSA0owT
QY8SXSMldtwLvcOGOYc43Nf9bwAjM21KThKm1v4qRvLwt33rNayZhV5/5XlN1jQl
ShjqATHOXjLfL38Dg6DpreRsmDIfZTURYzrEh/tu8elcpVhFE5xp0Vcp1HLJcNFg
grqOUz1lsKC3RmlBvKW+/57+ujQCX5ggyUXBlcKDWIbH45eZQeo53bqQ/gI1u42y
6JyENs0ZrfZnLf3UEQqbA21Nya/Nrtb4m6+4KUf9hh5nyjhM8VWfDhcpRxpY4GJE
qXFwoF+fDerKdZS3ClFTiQYUquo9f0bftWDEK03RXSaqVpuMnYNDmcuvL9P+hdQW
qajpzVb9uk4AYtGqMNWscmlLzLDF61Lx4oQhSfUYwBfo8msUPzeEB357/O29cjYK
yrLuVc6DjmyziSv9YQI0bA3qTP+EDMb/sty93yQ7BbtCnv72+GvMtpKoGt3X3EaE
PHPDLJYQfZZdevfXDygKPW4eo4fCIpDUmdqsMqoPmxcxctoQzKWLKm81UKrGOJp3
BQK2PsQ9ug7n0ttb3aUpBj/0E/aKHsrUZ0WpkB0cFGYC/m+WsxRt/rCSRHUhIpot
UeV9yzknWWzTWD45K1qfHreDWxWBaLzNpDXzbrAZPJGYklJ7lTZcTQy05/gKvGdC
hARZxndPn8VTRNqhf/usr1uU4q7BzM1/2EqwqsEjly7zPB2H9FRhswU4Y45vGc8+
9Sy6v3aqcCVyXsDuLoNKDCAeaBo6VTB/o1dYTvTV11Uw7tgU6uwvSM8eBvQei3gj
XagZ1jpY2ZIUXFCw/xgpU6s5F4gPpdblHRi6GD7qHLZrhkvgpqrJ0Q0lNcZQz2IL
FF0RBOLm6dD9G9amr3JABnFwvnHXkwjxXcnrEUF+rMouW3T7y1Sgp3OpUp98+xmG
hSKHKCAgwkvl8XRFqTt6RnQqrEwvAQZ+Bfy7svy7BJtY2m+fyWgAdsxP1rSUuqPa
NY+c2xmSUC0t16IuBvNJg2Mt1B5oBsnh3NRBYYaYHBgDdG+U2mr+sT5wRiEi0Ebz
Gl+1uhci6wZTE+EcnmMO+tac7d0QO2RMW8BT55qBAvcj4BBBMHsDTfrknZ5xILc9
kR2xObpnHjeKHQxDgdQusa7wvMdctYslsFqU7j3K6+odWqI/B2Zfi8F2KwObwSEE
AWetVv9FjBqpu2cPn8I6j8QTKRn1aF8mopn60Ge9KK+GvAAIO85FuiIS065gzsvV
gECplY3JXJZRirbpDRGJGJvPlnucCrrmyMxHMtGKWIP/GHPISZYawz6VHz7RJmvR
vqBN8ggCRsQU238VhYx2YgnS1e6YjBsnvqsHbKOvDvuoGBsvW4xJU/mbdd4vCIy1
hyTv3S0yPJU7dzDe8X+tqJy/z3J3JgzYtj8xBm6ha8jtuTVz+M+WUi2r/HftpbDe
AWWgmnAUNkXGIJ3j0peOabsA0d8APXWkYx0STOJ6gT6M4y8B0l0vFtRsAA9kCkgB
e9ZHcKJHS49//ESl8W1mUcQ3k7Rb8kkHJnb+SFznRqQqKsK/+2GIJAuginyc+JAh
DDZdNHcSL7UVKvwtWN2z463xiw/s2iMD/kCSGWx09bsOPq5nhGOyXUO5U2E2xuol
xPHBrx1BwNXym3BmwkSiqTiATvo4YzpgYBwTKG6XxCkmLZDqCL7dgSvP8kjpbk+9
778sWAxeLsaJL9p5fcuoZpZ0WRLEMduAQvWwuEnP9VtX1DGaZtioBYcwvlV1BXMI
DjJMZLLjw2ppxpljoYVf2lufS9L2MLoTV9lxPPyHGmZ5POJI70fBSFdLewHtzSed
pA2aYXrtz3jWGlVGkWrGuKJXFiocHUUo+307bL4nh0RGC1rp5ZXG9b/VDPvhyPXq
anEv95qxYxmkioWYVDrDu8Q1REebxD6eeTDpUNdjoSmC5N4uJyFYCdEY6x1LQ7+V
+RYMO96gS633H9/kTDlnsCqPU5gAuBg78pZNaKE3isbiL8n57uglRXfuIcW+6zfM
97+3PUZ/Sncg3ZhYXw85twMZY7pfLDD3mGo19OBW3Qtu9xodcNI7gu+B7sDfToF4
75+hvQmM2rT3uXqBWxv6lqI6J73bU67GGW5P197a00Z6bi1LEQdeji5k1g4Kh+Y6
3e8pk/UucdyAdkNDdnQ04ZsOEek3W59sYsL6dQYNv5P3k49l8R5Ltek98/kAt6DA
dn5fOpThexLLLhDNWjLSJRY+X36sM6za8z2TRyvk0Y4J3FPMGOS2qcl9w9Ou2oyh
WJSYoaaW0JpzXInwh5xsdtTJbL2T7unJE1c1vU8zseNsWI8BJTm3r5isqjgtkEa7
nQTfFOsYofBeFpc8kxd3tEECy7Jej1aOutP6pYexmR+YpIIIW13AuQmg6fvwm6Ec
CjnQGLWlyV6C1IycmyrkYEa4h+GzdNoUV0Phdc0F8HXFH6bYpUICPRnHDJGnI5Yo
yodlktXMDVOJovGttGiTE+WVdxCxLbZXV7aFm7EyId70Ilt2mKNycBJ4Xtfcy1Q1
Y4nSc3lnxyb49YCFLWlZbaSTf+WNhegREWzsiIJ6ppubfMuqJRQEHZpBJcMyOYtI
QqFSXkGs6efSu+FzkitQr8E/keaQKPvo4xlB9uZwXV9Q9rr2oFEny4PkVZjr9ce1
7lcse8h3AkErJ+7kbvduF0WB1wR0aCBI5Xg+s/tKmI5DtprK4R1cr0ylCCL3G0Xy
iwKnVYN91RvS1wbKWKxqQAsngVkAjQh1UxUJvoB+Ry6hMKOFDJesh7bp7iX5eAmx
yqrizRwmfTVjh9E/U+SYxH6Q1Heu1X6oDDBKID4f2ZXTO23Moei3lTsA/lIcEk3w
4z/eRUYCr0vGkJ3MDdOgCLB4dJ9ILA38b8Zcj9ZuRaoRWVDusqKHH9NFPhspUqmc
Dwqc3ab38+3CSMBdmtTTEBS2EbLoI3/r6GYhL7qqzMs6ZK8+zu7FAGACy7MMlpyH
zzUHrmckrZUFi/FYH72gYRK8UW+DPp9uKb3zw/1krz34zS09j3uocEwJi72puf5c
f7doxuWRu7932MTph66Y52UM9kRKZJQC5K0PqfGZuER7b1SXaJxMeZ8rxzNhhbPH
CuQdiGRRC3Pfhj8GidhqcX5M+eEPeDdsPx5A0XrfGFVRLSCWWiFVbyCJCgykzLnU
e66N68pfjmSrf7C9rn4gyGf9wIeNvkzvtUGGN06ahNeDAMDFD55tSocFeKFv7y95
kaPbZMhjvMcDXh+dNEst+dKH/TWwOJiZ5H5jzVCQtKe5p/bhQ35CjkfIVkOHYaXd
WC8RmqI8PhjFNsWnxOm5Vr2OYEHEtn5XqClVJLsphxyMDhPTivihrli43G599wkh
2B+ultfUN7/rqpqalqCyGaM/k9rxyCEAuDC+X+3MOdnJDQKDUOv1zfeKISNgggZg
darIG3/m7lTsd56m24XAZJZHBMTD2EzGhD1/ZzfVaCZFROUq42G+vCjQB8T/iJpf
Fz3nem3/U3lK7iI9C6bzNTZ3WoeXKGsXFfVZFgZjfT8UjBBUWa0AJ3zRAjhzJ9GU
9TTnOEyyLAvFaSn9g3FylA4gysGvs5cXo3YLRovDVOg6jxJh/L56DPSdRG637Ve8
rZBdx9FLcAOqedmRxvsTF06+GjmyFaHbQapf9aaL5fGsC8WZ2xsopzU6yK5x7WIX
gwdn2kHMeOGDE+C+/AF7TJHqZ25c1anh+sOSqtTVkhHFAzuF0J+8NZwBf9r3C8fi
mOiE/iu/e+hcxvfnJCmRbxMcR7Hr9fitABhYitCqHWQyQYdhVZbHNS0P8Kgy2PyW
a5L9ngX6XMYbhBPF4Oi/ytBV1t/SGRh3IguW4fqx6nPvt5rqmjMUZOQ6+Edu3uQb
HV4U/GezN7vRvRjUpiaI7p3v1P00OwDAWYXGV5dKrJw+yOT1mY1qWbGr5Ouxhts8
rg7e5jJJ8w3tv43QzrmBJjYHKzq6mypa8zqIwBfQUrWmDNaSza3dhE9KqavAZ61K
EnQd6azel78lUwLJuG1FRzLnG+O7q2zDF5wBxdoQtEtWYJvHGcWl2UZsWkZi+nUF
FdXlVzV/Xbbgsq38qZK6UVh8cp4vHMq4b4hS1M148E6g+nWtzWc9Udy3+Gjxq8Hl
tAp/3ASgfHgyoBItyrx4n0ntmHy/pggKbpsNXFvgFQOUs82wQQoxaYiWSb7QxcQj
R0+8IfkKixWyBgbIshI/tP6uUx3PPNGarUQ9ibmdqHSaNPh9vFu94Bq8uarNvvWf
sHFtOUZPfO+hKW5bhgpEFU1UVRKacxaeIxcXzw01uwis0WTawZnR/5MInhd3mxxP
HVZfwh1nVd0Cly7OSYHb6imsH69aa41Q8ltm2N3AGn+FcQxJ+38bRT0V8juVEx0J
7HPk2/12rQox+52neoVaOHKyWoId7jLiuzR/EG3b3ezsuRJqqRJKuFPkQHtqXWPN
/nu1ifVX3iLl18SV/jTdah2ZgoGjTq6f4rPohOiuPs7ngOxvqtAmaOGS7nG2bX6x
Iv1e/evYCDQGrFwJ0Z4kuLFkI7eeOAoJKfi+6dnuqSViqVyCtC/RQdA8mxdFsxUf
/ikr3xMf650ZgG7MT4vt9qc5gZai0DmRfVqgrHc3WuxWztM12soZ+DGdV8FjrXDz
nYIjANfO4ZhrvBHVL8Nv0FXmfOJfPMsVFcS7bdwYbRTlypHH+YH4yy382u2/qPlO
WlSrt2EMw+35X5+83ytVgveVESO9bnIj617Gq3CGkPfBZwaeU3nSYdBzJi/BpSD2
bg7BRCe/MQTfQ7u/YeDMFKAOMdXT3mTz21HY+WVv5h0xY77UuNHcik13cBJ2l6cl
Rktg7XEF0VrDNK+c9F9vwqy1yvBJ/5mVg2YFIyelnPkAKsYAwBXfYtfRY76mjYa9
nnlGiNOt928drT98J/kujfm7hi9QyQwFIMvY75el02dDlgHDHpHt8znQckg3W2YZ
Wv3Bempr5ipQI3pqR6+rpu8j8Eo9JjqOr1vFVqOvATnQ5+ZOjqy9av9OlOLmd2pk
fqBrr1AqIWi02m8K978vmgWgXhcCBjFj49X0wNd7fnyNzZ9v64lGtjfPIoi/mBaE
J9Pb/ZpD2yaLp1OMbc30aoLN+AeGUJfVQHMskvIhlp+EfQco5ZdUl3WfEGRk1RiT
SnsSrXbGAAf6prQOgweBTb79KcKX+06po9Hq+X43aXC9+t+7c9k2l5M7P4dp/zYe
t8+TTtqsIc6yupwR8TQQJNQb2/kYzzubNTaBEjlgacbPGDQepNJNsrvwux3LFELI
P9M3GByeTIBmHSMSGYojWncNudwcLuRUYybh9gcI6ltku2IK86rSbCWs7eCncWJ+
JJivKJqVlfY62OojEdTjQ9jutTJJDwVOrPB1LAzGoKz0n2hx6Ri/2y0qbMcAbA9v
wUGRgy+N7Za0gLQVwEHWeoFXD5esMj955rlJZGRVvbKl6ueJroRm/T7eRW43s/fK
kfmz6yFcFWpXTRdGDa/5g4g9NQ1OzREiCrPdMUEa5zkHezPNMAAPea79lQnYU7xg
NpMVD0RU73Ln4wzludXaSRxZ9UhqR5FSZJhRqi65f62oHcH+qkLBldP8nd+POEu3
y0tNbsWfG/GXGp8eqBT8BtxDAXJ5Sz5JlQdz+Okz5S77Z1x1IgMsFXCKYlRfzX9k
kF0OaCaFkdQk6+3PBb7vUzHUlgcbzk2TafLw7jphzeuZVHdETH+kFL//pA5gQ74l
gkDPZ7rICUfZ4DCrcYEY/Ao1fX3ihkF9zXHVAhFnjezdyvcB006hOaIVoNTEwzRt
0XjH/Ibi6mlNweBBvfgfvdOCQtclinc+m5g9iWDQHlFbbV/Tmw9/AglxHAjWFA//
yM26mB1CIt+kfVQa45kL6I3zjbIGq9LCUNEiMbhfiVze6I10w28RRQJky0/j237p
QrMMIvb57xddBbRDlHGl/feJmVY+OY48VnJPm3XxHQHbp5dkZFwjkCglT/FrCEtD
bzpY4lgAoD9zHhw0Gn2dVbOEwKZRlhl0oq69zoA0Pe/x27A+sT0MvKnASmLwWFc/
4Ko/vr76xtIxarK9/HiWhmMN7OvnIqLMCPjAD6JGaFssEfkZwcQSTrsCFf8CfhhA
AvvZsU5J/FXdP6NUHUcX9zqpaQQhdwSxt3jX5ReWtYC9xJ13AyQFJtYs59iSXoFp
TusluJ5SIrN0+vIUfES9MHUGGZphSVhJdt+FwuzZlmi5WRZQw87AzTYrqYGkFuMU
3HWDtmBE8fh8KNQbMYZbWJ+YfYch+az1vkDALaAJxP910ehdHOWz4hG8tOU5oEWr
nUKko6OWxioUsTLKoNXBT03KgISR8fEWQGhhySzLrI5VA+8+cc6zU2sIdVSlP4oH
3Az96t2Twgx2rdDeRESE7HD1/FeL15HvUEHPTmn4wALyl8Rk87aTD1pBMFcIc/3r
KN5BibmiG/asjYZu98MItsxD+R6oQrDLhDBvtJWG2ibCjqKlEu2mTTMpcH+1OgIj
STNZd6KE5wWWfKDasMxgQd08IGCAiKH8FwSNRBcfWu+HmjZ53iOsYTBjMQNimZIy
D7nUJmGIzt2l7b0ciOmWDwWjUob0vg+NUK+ifEklpleNhhHvNsRJ/VawCFRMCyV3
OV1RV2O+Al3SRhAFYSR7UcAT8iNfYHvaHsttuaTlaP2JhkpsNH4egQ2aNJ9aGQ4r
IZG0Eow4iXHdwbH4GMi9DeLPdjhW1xN5g2y0s6CZOp+/MdB9AEIIXZ4fg/eLtbWE
0OMeFGkZKYEU6oDytCfUFwJFkbXAsj1iy0PyP1PcM3iJVPKhmmGFV7Qk01ofPU8F
FVsaPDpRsxKi8/TqO5ldkX5ZGGqGoci3z7BrHsR0kGYlG45R6BhOW7uvqGHv9QLd
5pGDqNVkLVTN4tlot9PMlN8+4qEMmZ8LdeM2cq2poYVnJSFbxxOR5meYq/ov6BSD
eBs5/KSu3cu17cg+h+X0KWGEjW5KLxISrWLSK/aLhGt6ajo/iKZzPPoP6D0TYG2t
6fNBNZuAUmnuX28NZXWDxV33EOsrfmdju271o3bizKMhtoU5989XhByCDEaNnaRF
lDZPcEx1OecETeSfJmxvbbw9K37UgyQxWNr4nVRxWoj1gzGuuCYLyWMdnIity1qw
mzUzakELzFn3t6re0r94SjiB6WKBqqKTv5gi4hF6ocRW1yadvFp6nOF9Q6TJIs02
s2jmLAqWrwzXUVJ9KHG5RWZBoClbwn8gNjIFwmt1s4iOgHbTEuYAmEkZVyfzVNKU
nAmVEYnPxYpB0kCo/9IOQTiQ+Ryj9Md4TtFqSRBQmPTQRvM4F0F+ZU9XOlZfFPJF
bRVVk1X8/40MZgWL5yPn93t+PN5bNb7bhTTqbmiPNxk+GkDLNY9cFWJHeAioF5eY
kVeLohz+Kbus90LSFhUs8wjDTO0ZTS9Pdtx1u6ryWCu6a/rW+lBtUAEXZuqfJ12v
xv+vZGzX9I5NNZQqajYTt1I16actVeK04RH2Y4e99ErQHKglfPNGfFwlc+XKJthw
s9xUfyLZiORByeVfwawtvYSz4L7Y/nZrz/ydor/xhl59qQKQhuTmBWD382bXYaWj
mz1qEZbqti8yVx2Av2IxAD5+nVwksoHLJ+jun4ClSrne1uzim4DqBReZymwS/WXV
iGO8UT3d4bkRoTadHz6sIuoxSVJx0QvDWrtPnytMoufj+18svhcZ+mQh/Ii6i5ht
Ry9NTrR2EFSpFCW1ajHxpBrFRN5387RbkHBMUCA9TZpu2MuyaHpqMmAHah69wpnx
spIDRcfdM4300dnt/1ENCOZrijccjg0rRvh7g0mqSIdWlLVN5zaLszDs+T//d6Wz
N9ZOgDC2Bry1WstvX4g7umhrlwNlDfh4EQJk+P8cSPUDob5i60ieFrf3Cni/6a6d
aI3Nnhd2PPKIxFBmAZh70Ji3N8y70ua4aXrBa5ApoDaYNJLVDT14sw7klioI8jWy
A7+4sfi8gQ+mvu4ziaBNer9chtTmSFhjJcg/Ebg7KrH7pQSgiuGlcUcMIhBNFj/V
QAMdJXzRRd6/FCR66daZGx2mJ29qTnBdh27yRq5lobbkiLkSbcVfpgxGrH+2I3zL
3JOzn4aL/901lLq2AdYsHoBW0f9P+ZQmepSaXVMj6qrV8TNT2zHJ4w28DcvIPM+x
UGOHkzzZqhzLv8zQRBKIOkZ8Bh3ixnoV0mF7Qqb/gm6g4JYQv9Rv1Ra6OQjn2rw4
QdwCMwPtm2/R0HbOXgzH5f4XcnkxO75pKb/OQiEnRXVGrhiCrjBIZhld9qPMCPub
grvjXDcDGFxD7yl+KmqWGkeoFHD3AJDgoj+v0V9lmmFzlFZQ7hXKdH4VQ/0GP5AL
0PrFr+apIFix/DtDINtqoI+08JlMOe4/dHNUxwRUxiJ67yZPk6fzXBQ6GviiusO9
/+Csy1w+ueX6f6ZWXulhPDkDUN0RvpkAH9nBohkSyYqjGZrhNcgw2xGaStQrV1yB
Hb79ufG8m84PDE1emv9Tlgso4/Uk7lpKlDU7SYfFgxcuD1N+dc53IIg2/ao1oPNj
mvuBIdMrJlrQ+KTYHwgy5FtmnlBl5VDAz6COQB/vuOroDLbASgzcWgUWtYgqdtj8
8mmwwd3IrW8xE7wwgrTE9MljYk8AD37piGvxXXnIYaBkYq4fy/b0I/FOKQoUDzXb
x+x0K1oSpBUy2kBzhoFqITLZ+zmC5T4FxW+1D643RkKf6AhCuOS8XIqFYR0intwO
k/wJ4QqMCDtMOIPLWAUwhmMa6YkRXBoE8TZ8vEfPG1XF2d6rxI5Dz0+xi/tgL8nj
bTYQ8CK8WMs04ZqANvjd64r/W416f/PHiRlc7EkKQKIFK/s409m2XoPo7S2oNhs8
ZFGs3AFFrU83PZ6rZwHwwhtZWfBZBuYxHt8ZomutKLvVxqnD+DETfcyHyc+8XqaM
xBuyfi7LFJ49V6EHWRuUklhdS+RImBsjDuIup8QOizlHZf4mhPHvRoEROhwARcPJ
36myIG/mxeHYB2qALG2UJ5PCk4VbIuAD2N1bTGrmR/NUiZgmk02ES1TkgIjJMcNf
fR+Ln87A4mmdf9/3FWVeKIrCgXaLeA42j5v6a0Z5aeECMO74jwRy82jBTUXsiIMl
2+RJ5XdJZJGf52VTE0s7FTE6gi2xkFnea2tflk/6eVhegwyfkglR3b1xgk57HJK2
HZG3K2dhId/Ssh6XNPc+xu60+R9cujyp3paUA2l2Uz6s0ilSQTDHRUngwYkqj98Y
rJMhN99tXaz+33BM0qaGysN9cNUkcJaw+hWz8uSBpeEWeAKPfd+rRnBZfLArvApE
Xg/tqJRWPKhllwDYenHmvuPXp0Zi4nsMJKhIUAx7iTCGmCPFS/yrv/zZxXjPpR6N
5/w43rP09GhRo9D+CXKmfLOgtG1VktNQ3P5x2lfc37x0MYfHXiZt1rpm8wK6/Qte
I4pQTtQlzf3CMVS+z6TwViFoKjsiiawkl9zk4mBZ/2tzQkZI2OWMGgfqa/UKV/Mj
0zudyuCt5TQyiDYvOeS7VdXMldu5YXEqxQOpk1US1Pa8sKQVKCzJEEKqM28g5cuN
bmNXs6WdlQhk9joNOkasTjc3fe4TyxFuMpXHDoPuEuDFLpL7249+ua5MF60xWV9t
kF96apDrbTDRy0cdVpsHzZ8Vv51VkJjQk/Ygd3Nbec2Agz5xKZ630uuMXt8UZa9/
DHhifWbyg7Zmvxo65JET944TnpLvDLu72+d/wgTS1QcYb+mn63LU317PO69TuNmv
jf1hWip9LFTv84dhn8GcNOqO22I75DcELMDKsOuYhEmVl7SM6yXqzEfq2XhTIZyO
XDKpRyf0Z5UAR0ry4VvbcVrisP9oZx20GXkBidwHrCeW3ZorJbc1tcno+S6nQXjh
gX0I/dpi38tEFif4LBnwJ3N6xZHiUd2Kus2ERw9LtqyovU6w5HPpRZrwA0PZ7fO/
sQM96x0njfbfQUbiN9D5XzwjU1aaz5aNVOpACCVzLlPXi7J5jZyFPJIVHLrMEvcJ
gbP6fowdweb584xHdWhmhQkCAmy7eR+yY9d0iQx+kYJhzuiNoMEspaVfNBvIGBOY
/pU5nvN8edmvzwHJGaPJZeiHTCEk7giLMyxohlm62YNGqlojQM0um/tUVrdqtjrG
wp5g+8sEdTgy8722aQ7IZWK0RSlPG0F4LU/i2aa3UAYS2yiitYjYHMNsYHj3zRPQ
a0vrNlP90YBASo+Rbcb7Q9BbLeTrnGTAIM6AmCJ/dXGFF/LHc4S19x73KpCcp/eP
2Xb/97pURa3basNTwJB8em6/6GSkRlnPLa8So5ubm5LV5eBDjyFzva7oKR6g0Gqk
VMhNMy+7KVMlaY/X0wHZB9Fn7ony92oKnQ+wS71RsQbMsZBrUCM7hj7o96ENpzpa
cNT4Wv9llzYd5NJjLHsnkhrvVH/3urKvadhWyaAsjv5bkTwfaeOH8AuKymV5GD50
L6H9G0DQlWUz8CUhqlhhkT8I6Pxm4+ZrNfh08CAyKPWrOQbDjmK5cqXRddpwdD2S
fdIp7NM9cK1+SHj78nxZWa3J5+6eAS3p+d/tvPd8XULwssFbpooKVVt8bPsIe4sV
r3xsLhPi94OZPVz2IsJlWRIhnWGoWM491B+OqQYj9N3K/mjxARNdn0ZcV1J5OsOC
ZqkPfs61yWPQlchMowy982Vxm/betfyKxXG8kJ0IAMX/hjn7pf1kODJ+hNqEhKC1
/J4K2hiXZwLL+7+LHBr3u8rD65jtlxrJNBNG2hMjQQsW0jnOB71D5fCVCqZaQ4TU
8se1gdAiX54RY5ECpnURxzicSyuJpWN2/aezi47lCJ3k1+JbVmDsr1yVM3kGHqnh
j5Ng8hdToWPp+DjbTeYrDW4zomBGeQUCapruClfBpyDbGoFXtTHysvWawiwxyE2s
9Y6li0ykOYLcKymyRNllGeIkpLE4eu/JKlhBAWlfLbsEY3rok3JKJqt+3A87OKJ/
m2envCNs/A5qMVZC2SF5+e6GnMsUSR3ArpqqrLUCkVLsZwdUUW1GaeturY+AwvaF
HawLvjbFV56kV7SrsXcaqcZ8ZHmhsLWPHT5ehOwwVP5mYiTAtkTsWC1wRXV9q+Be
xD29/W+5VD7m+E9OEcQBw4fQCYUon0fSMPge3JXkmhVs+5XDan0hRqFbHKuarDtT
KouAbODkpmjuBIwyH3zIPmASADJxO3W9oL3VZnguRVwcQeDAcmy41fkffBT/9UvC
Vivi8fI0E9R3QnwJmnHzaf3XBkopHkj570P786+Fu0YIjAGX79W1zgllMcaTxdzi
OjZamkb8Ti38Cze331AmUfUdXF0sQ4S7PfiWa5X6bPhf/VSDxpM4N2Yr//zlK5QH
mqxvEznc1z/VOumb+/mEiQytWxy1oL7nSgr0Uq6gTKKaEINhVGrakP5Y68kDzytn
MA9GeQdPtEOAbe6VjIM56ge9X9SMZejlxaeggn1JtkgOQQhRns18W1D0o4JmaS5h
yWVjKzz4tZae3BD9VT5PPGbjIbfy9LtxBWe9vRJ8yuDaDxMPHmnBFX7anGDgmE2o
vNb13bCnWGWPf1vtl2gq34GUtDQdhfvLDTOtsFXXmoaxznP0qdxZctCFn9xub3Ew
13/aJRirlXOAdZNr21BRO/8DAJWNeqtJASqNlbqzCVuSLfbJHUVF6g+lEbs5KemT
emLK6REPZUCgTwkeNzSrjHOMFhF09s+bG0L6lIWE8aNVmMAFHqV64h++Wo0RXOGL
ldpd0Dm/wtvL3n7DocE7L6yqQzXJWXYyw0/KPTkqeJ+3WIRUosv4ly19bTPE+48X
gUKVjgjS1EFo3l2I5ja21uHiqA+TxghhjRxHa+4/6L0asHy5hdRQeuhEaDgi5pOG
P/GJ7HLENcTB83UVKPHfe4Fg3Lz5KopDAlG29yrEtn1mx5ECtp5qhQhXLzy5xebi
cLRs34zaf0EKBC0lOB4auNhgw48rsmkDVu2iM+T9HWUj7WlNxwY7FhrI3HuYWJPc
Yo/1tqkzIm1v37OJLWQC6jNVhT6ZJsnGyk3KowesaPE6vn2AuqmURZLvKILI9hQF
zPzVNYd4M17zhbT4TxLqnHGqfqs5P5QTtv+LHhJCubqnUmsPE3uSt4tPLsCTYSrA
mbWQt1Vy5HU2u9SwaNN0Ul3Zr00eI4RMMn5TtfZLSFSXgG0OURiwbLz8vZ0IRvZH
JeMhxipTgxplAadqM7tnAPqpH2CPmR0zuqQKU3rHjxdktynLH01ZOVKQZpUqX6vf
Nh30VPEYXKF22G0hL/ydJ85ac6q5vfyXNqfntBiuouwLpURKM8NYGOkyxUJi61nM
+KBYORmUL5eV6dek0Z90Mr9Piuzik8XCQjgAunwXsWVsgc7mT5NmUZQmc4r6BQZ/
z7F4qxxi7C7imn+sLPikvc5+rm1gtaGNL2Hx/AF+XFgbuCEe4I0NAyO5lFHXYjp0
iKUi1F8AV8PLbGl4+X1wRph+d3CDPPYk4WwzQ4/OPEHjd8hviT7nRmxDnWeDYrqV
z6L2isooydSCdXL9wWa5mvSMhbB4Z65Cyvx0xNX9YT/bImHpR3fWLCseWBoxZYhp
qGN1G9aSlyP8xlYnKcOXI5sHO5R5Nu2rGBl7fUyhN4oNGc8eQl1FWQUN5BUaCn28
HjgNGnnjEhtQQVfwFIl6sN9dVmEmaf88hXyQ+9xOC6vdT+WDL95lhMlF5vOpP0n8
gFCZoLZYoAZrHDbqIsfK0ggi62gMXP30qbKKJcnmNRX9R5Mpcu38GGyhuUmOTT9r
TJHlWJ7oHiBARs999nP9Rsj1jRGRX6h5oZI+cvYy2gsM6PrRXUrAnjvtI7yRqC7X
tINL8zsaScPXauha4rA6b6fcZBiscsX16Ims7HlueB9pXoXV1RhrJjPF6uSlX6HI
UnhUTAGfGt+gSywX1xzK5U+XgtWOyIfGqOPC3ICCG1Haqk0Q1cH5XrLhf9S7doiX
/XcyN4P9GaOk9HKyXRKL3EGe3zie8ptWcoeCXpdKrEFs1oXlzERsuyd92kRYEjfO
DNcOrqwV1BIak7iPFEpen+BU3ZTfbdIAhWyRjkKfwAoMmKyb2JVPbOb7xMYkNtUd
EzyB6Df8L6lYQUTFgPRlPVoCfZnCKd+m7Z0N1Sx4CM9SOI7E1hu3DchwOXPtFE/C
IoA5wCcDewSGZo3uR8kUUNRiynEyySaGv7S8+QsYq/cyt7xYJdnPqFwHgnWnv4Br
9VTKOBTXPVA7Fl3KojXqE590zD5Bw8QXCSuZ7iXv9gyecGA+jYgjv1FbCzlXodn0
jXaaRoNQ2p0B3YACDmoHv3J/wRTW1jTfI4z6FCT5uouBqZfiJNfhPNiyBSOLzGA/
SL2sNBFaNMibgyay6broB9FezcHvyNKbwWRcMflisET2AS/Uma2n3ihWah91Hnec
ZsgMi/dqH8lLaWzvRZy67NWlZgCHLQ9qVZI/3D8l9ijGwDFhuVKAC+umq2dIgv46
1nDvXrp0tIIwYQBkTAKWujWakuY6j4e34+CFCt/7o7IIGHMaLV5w/nLcCXVgoA8r
BrMHvqKAFfOmSQAsNDct2d/KNFgC3cV2rrz9nQ5eJUcoQbKRfBstc/WS3uIWyE9T
Q/UsBhXyeNr5I1bhuu/17v0nM81futvYxWhfmEp85eyIcvxybDtRd2MMdiTdLf7U
HTVHzcYivy5hpOQR4bKengo2ISQg1bSIYL8bawoBKcApIKb3kcj2SQBTHyBwQJFc
pbaimzEwXGh5YFiwW+ix+VdImzm+7SyNYeK3MgIjFjIQ8xM1TxG3pWwaEQwZBn+J
JosV1PYAanUfUDT+lrIovIhaY3nZny5jJYKGBYT0MLKSl2/8GpONBOQ8dOyS7gDM
wQMUjSfvceBBLiuUwQDJ4vOpmwK+NojWzYHXhEPCQXOFG6K+9ghyAeu4q7LQrru8
MK2kodqKUPTANnxExCM/sL0Cu8rpC0SD9zMQ7M+HSw4fhJnxt8LNfentBCYT1IO3
4yxFNJesPLKLs68PnHz/p87LU3pRXvOt+82hR2zg8ZQ/T9gDOxelmE6nNbrGemOo
14fmiWHOrVbL2OwG4T8afgmRAW154p4VBmKzBlXJAqg0myUb5UfVPk4RzMZiOPtl
+X91hme+kHvuL2a2S7Tb0aQO4UALNrXQcS0VSF0hNpRhIUNPc2vG6a0E3YraLFhS
Lp39+vitKLW1X5bb9KOMKdOE70KMZupOtWoXDttmhR9hmue1ZWrt3NFYtgB2dR8I
Wf+0iHFP0glJr3mYltev8/7Zaocy0TwWBBLdp26J5FPW1D6vegVw9CuRTYrI18Nr
k3vi40XDxy+hQvvX8oZ7cIGPj/95OvKeKzDvJAHeiV3pC6i1F+d/lySRf6h1uVeI
8x5RfhpJk1g1Wx8oX1UhEmEvmmlHJGOU2aE88fLNI43XuNMVYhicYVmim+1APRqX
nxwCw3adovfUoz6eZ4r+dM35dhO4mpA1ulyYyVPHvR8gMa05TDGFv/zWFOXCYDCa
h56lNrr632IdWfq6k8G8WPzkUIiJHZ7mj0dc2HQgQvkDlubcFvanxM+O1dSF28BK
jjSy0XTI4BeCu46AazJYgKJBlypMALNbT53dsvVWdXtHBkmzGlKReUoTuTBAB6md
jL/whvmcBVxlcjAFYjjEGGbbCD3laAT7CRRxI5eRPYi+wP1FdFooBoDmW8igHE15
o0Te0HeGtXxZBd+iEJWSE7O6rEd31T+IVF/1o6nNcRe07GMCZRssJGYAmB0QTVId
2K/sEgas/0yvfrBZ3RFzbyUXiMGiCBuR5TNuaks5hCVel6KGrIxWRmHLSC035ksb
RCFcqZc58+SS/3+sTLnStZ40EAmshArRMc2RwgKyhb150kLNmBeDcCg3iPLOxv8b
pQkB7J6/aDBH05Hqpf4F+U59GkftpEmYpaDrNF+0vvbs72gkW2A8U8Dq/6PAfMut
K2cN9l+8TF+digDyhxrjLuYMEhzIVOxpcWV6YBxnj7psF//Fn889b2P5jl4SLT4/
mJKFzv4AUP9uvX0aUmC54b8yPG6YN7Wa1OtWrJtyi2xUM7j8BHjb3qudpTuufL1g
5bnpdUTOO/MeXASP2n3Nktc/ZaptoqPPm40bXIkzWBno5QiSP6naVj3CjkXO0uU1
kbuzfP+JRmx7WUUPQWljuTaNthKuO76gG2i3Ig1+xOvUrmSHha0jA07CIabf+LDC
ZhHscoVqNkksGd04Dqcsn0OIzGj1NEPepkSuBbCQ7eriQI3ZIR8ag/9wdMN433u3
i25suihcvj1sA2mxhMRq4MAva0Y3QbJC/ds+Rpi3xfaUOwso1ewE3YhiJqL9ya1U
nBAIEoggXdfPSc0mV6FM3hpFa3Dj3+mvsciFc0ILBkx0mV2VV1+oIVZnnV72V4+I
Jhzr4tLqzsjF7tCXf7RtBpffBJGVqauaAZPIIW9riGB+hz455hUoeAqdrwLEjviz
Pqla2C8OId/vIxpeEowkPZKTM9LDzq5g1QAwrfV4N0Fta+LK2XPMoMAKitXHiVuZ
LGCN750R73r7Y3/eWB/nueziHB6AuILN8EwBmy9y8ZFDHlSCou9DcPtsdltWI6Qt
BLrM7rBy95i5CfBcVTIv8jPbVGZU6+AtufEDnnYw9TcEI57WIh5G50MYbvM+byNg
tugERvQLfIvwetgtwefeW3X5EgCwufh7qRf8UPLt64Z3mJgF/6kcjIu+TTVkvlUG
x+T7KobMr0B/gHqKcsCuGL/+X0lNVbnFgGokAFD2aOScelfqiJIU3CCvLDHD+j3+
u1PwmacdVS6Ow//BJRuaxgAHb0AmeRgKpFOf7G49/CL6bMVXgWPJ3+nRRLxsQXMV
rDKjr1rfCdufDmR16vTKvjckYjwj2j0aQJLTwU6Eh6MGJKHbGjNYRcjtG4R5+54Y
dIQfEN0b0E+H5TU9hfgePl9KIXbqD4ozq1QDqE1jDE64KcT65FN/YeD0FP3d81mx
l7ZobD3fpCsfpVOdWPuiPvYhJPAofDDOPVLjswwZOOuuQTpLGDHtfefxC6L6/5QH
I6xlVwhSlzp4YF3MUYDmNePVDY2zPqHMV6OaCiUGzwHcz8jq3/Iwl2hg2uIUaYXT
k/A5pizcA8PC+79uuFLRTk/DJQNUvhDCi43pBGkulanI/U7waCV1G7ZrdXbgb122
sVAK4XfH10qJrnG/pmQtuhVvpbWrlLKXd2nkoRpzHkUzW3Kl1NLjt+Tg0joMrOtC
W2v0XQ8VGFD7ksrPh/bmgzTss2FL0fLHmSpgxRH5OiPdlnZdTvF0e9LfJNbCjle4
GMl5sa0wQknQE89fsC7ZN3W2d6oPPAgwNnho/hJfIy2BgXhoroiJSrC3v8fhmSyd
lMqJNp8ydq/TzB5X9wvrayRI/Z8eN9KOsi1Ml3+Bo8PjBF2XWRkwI/Z12zD4dOjw
LvhnV5G0S9qQsypnYEiFw9ovS+PgrT07zRCK1nz0iZjs0LAgtEkQPcL4Vw/HXq5a
QEDW4eOJm6XJVhnCE2TzfgZhL4qrwPlr4NnT5kwnOYrR3gNL6iISvKIavAeNlqU8
e59N0U6W4bTY6FBi5zmjhzo/QBWmYfaGvWfrrRH0RAxxyLjDc8RVwXsCSo9lOsBI
zPkCo0+Sjy9D8Gw0FoTCG906qOmL8KEyQBLAoJYFMD7g64w79UY5VowLQVB7QzYC
q/CVFEtOVWjCyjX47K36pFAzCA6kL+mvHIfr9SPucPnHuOSwFYH95AWLukyeGqOI
LRj9g66kxEaemDBPoC7UHj3NzXYPOKbaFJeQmH+XIMSmQA/DUVGiQCOAx91jwD7e
TvLEISjgYt6P3WRB/g3a61Xpm2dv8upPY+wQkwIg27xYhCe0bPkH5uaEP42W1qMa
E7xF1EquiMeLS47UrYOQY+doMCsQgOOZVSeyXtJRKC66SQ7LJVHzfBZmqJiLRBN9
9tojOYfYRifw8BTR1/siduNH/yiC9XvnueHPcq4CADSqm/dDlZswkO0nhAT9FFV9
PjZ8H8dTbfxMH7kvOs0aGE5pzBW38De+Cy/zTHajCepxZCvEwBZrfMfaY2Xvi5Nq
3yPi+GNw68QykvqRtNH1HIoOHQDS/O5RK91s/Lusg+QXkeqFb3OvsVHAssTweFf+
uwORN3Z2UdQMQRA4BeOl0Pr/WXlh9AINCNUtIjyUMQK+RiZf8iqGSsb22Q3bdWkw
PAWbJd7QnGrNudjElGKoRNiRz1oe0KhnNW4NYqUM7xjT5GvK3OOHB0JzMf9zfNO5
2vuiybz9TLdfMlpidgrtcZ/yOjxw2T4o9U2Yet6II85Gf9zZ/H1qKwSa4D+lEwtF
QY8oeGufUCuulivqMOKYd+y1adwOVy1TKpP9P9fb3QsjzJoexE0266myaCW+ltee
m/kO2hWlj6B9HDZa+8fCBEMEjNDBp1LAU5yYCBNATf5XM6Ndo+ZGeP3AxwfSmm3b
KA2LXOCuiMENl0ljPJtX6uXz0hu+CgMjPsvH6lPDd/FtCmyy37Gk+TOxnaNkhuth
Ae1CNcPWItwzyRulMtAIx8k+EErsKh8C8hmRZSbkx3CrIMw89sEDHbQIjFXAB2XF
/HRbkB60j74AF28LVx6E1UrOd1q0fHOBMV/hZxAii+ETFxKs3kWABB8lTlQZeSkk
+op64vjkaNibgoqH1x/uSxOfaMTXyj+RafMCvS1HzW8fBCyXKVTtr7vw/rOYeTlz
K4Na+rz9+eumLU/2gy1YuEqBQKDrT4alA+cl7+7RMmVXdoIGML0EnOrICfRfKei7
qJVlDpBpqZ6ZORrzD7Zs7HyOwhJfoSPKlLxJnnMpyVY69XJrVO5ZH8ks/BR+H+EV
3otUkGTp8BQZGAisfmTDUPar5vUc/SaXePzxbFwhNScY/GdOr4vgFIHpyWQSfvzE
wX6QvvDkNqQOlxI/Ib3PXkuEKhCmCS8o7nmmLw40RUnGG50GHFzMnoO7CRUF9/ro
KsqlzYDGX3Yy4XoooYMTOFqnS5PraszpsBvxdmwB65ZEaH+6fnBHPHIW1DXsw53l
xiyfg82V8stA7M2+q4jVI4lWxK9YBucH8Sfse/sFa+Zc/nFulkdaGuOR5sVqO2Ms
8ChBlh90Kt0J0goGLiEmB11dxhZ2RKU/mv5sp4V1Mj+VwJkKC7XNbUJAVTKD9XHX
l6T+A3EogskI1mMaXXMCe9cELOd2qn1M7fAxiEqodRr73pnY4XKchdccXDVdMM5p
MgOcxRPuxBSsAi8t8JRq0bsIom+STCAXnA2AFqtQhfvBgz4xZSU0KrzXz1zbBchT
x7y9W3gNNydr0n2pNlyWWvGRtY1a4X/jxLbDslp9Qhvpetn8zdtkq7MZfE4B/xH1
+G2F0fQiywXnaI4qDRP3iwKEzo48qKZK0D80CKsl+qfIKxRMVdGGfuHw0I7W0EPm
lLMPjafd8i2Lb4oLwUW82asS9Wr3MGJZQfDeXDl33krAR3zoYcpcZm5FoAU9Sa/0
tfgFLKHshdAzOKJzv+C489molQ3MQLcyYakt2yZFgjHOn6X5Z2261DTEdBe4LVrl
rDkuCY+1HEW+GDL4fnkferusyhoPtl0LnYvNbugnRTwzmHNTVBVpX1BcvYa3uDvB
r278093X2hA4d5ywQiycGdNxAw5j4OVDVeOaUcgSBY4+YHb5z/3iPiFLP+dw/qpT
B1cIEds0c/OJpIVzQbAq+MUeQmLUZ2Gm1be0F+Mz9n/kfWen+Mxd1ldhyQYIg8uU
gzyYyuLcmzVb5F2FFMTen5yjtyzNGDCILU3CCc+jaL/EQV3QRpKjUBH99ro31u8r
AJvYKBHnTfPEWf2d4hhDjU8GH1rXKmreancvPcaxHf9KeusE9R/u2+8p+fmQXvIv
UZRavtVZI0DmJIXhaPIuDXQPQfiTwUDOMNjKIDOwmUKDcagfuh4qLF303TQ1KYei
EXOpQAP9n+TCvokV4oSUV6OPrXR9/UFZOgYk5HBZ285CjL5rnxifA/r+XdqkjrdI
eDLxWvfUuEgEfXf/AaHTfrSXhNLHA9G8sjzBrDp1ohsKc12oWBLw8BnF2S6md8Sn
/9cz+7XarL3oYu3iv6z9Ukg+0p4rHdlinFSV4gbM9IwnGwDKx0cvgOsqLDAFe5pp
2G1e6VAVaSLOqd8eIS8FxMNAN6Yp7BnWlUfAUH02vIMGMudnNzeyJPZxru3l9jKJ
TYYbojFQZaxWwoOhL8dEzqNMhPJ2DGlxmDGoWQ2Qzc/VfF4cBlI0TtaNa9QHSvdV
qtFKd3np+W9NpjB9V/zjF5z5CdvvgS+vf+jtpxRZR2zuaQwNsEhguDWcbMuCp26h
BlYHpAfKdLIsMc7OFAg3PVI2Kt4RtvT5vWmz2+/yWImw3sT/+jOBIqlCMLaR8jxO
cdvvt4aTZ4wJQE6mvPbdwnzk8RlyjKAB6mo5ZXd90DRU50s9GIxR3OQu21G6c/F2
mdVuyeKOK6OyIXkZCqjOJcS04v0/7NSZsVENYwJeBf/biOvpsDoZOOM3XwFPCxFJ
KrTDukPr726LarUOVYXaZOeyXIdfLKgH9uImB+pGEa0H/t9GhTanHxmHGL4/lD33
rG6cc/WIBNX7tRIVcE4LotTffZpK12avPJUB7NeyHe7HCnnxCVgKjT41GW45yz0t
SU11DRqSp7H9Rt1Pt4VvAyfCk9zkHyjV95RHm8FsU+s+GCDGlH13btdFAXRpFuH8
2ZHbSu9+zZABYnfhgNmn3GRqBE6Thx5n8zzGamQv5C7Su8ClX7NZTJvmZKWLWqS2
CThB1kgE/onKNiX5qgi9mEprTzJ/ulLp8vr73PSYwcPi99MzJ8iBXkenJeu48SQN
9C3ATyaiChwDY+AmtMov02CdDP1OGLxE6ZqwPJjbkvGC5tQlOXyguTOKyIfWsV5Z
CukqbYiAL/8hO4WpW+a8rkoVb7RP5Cn85RdWpzQQ+cFU5qEYmWQGy4DYgR8U38Le
bq07RgyJCgYf2ZGOHENqK1u3qRnZ/vc1eRqEVh5/tPFIh7MeQEDg0RhFM6ocswnB
6cuihCC52gfE8OgJzUugWtAogpcp8ouiEvrG0QRjEqxKTH4hXUefSCfWdsqePz93
QNRhYVeJXUYdF/2vop/tQmowORLwBIX6/siNh1aT/LiCgYnS/Xor7WxqxIvxM9LZ
QSzl6i+Rb9heSIsHWPPqZXK4+JnipP+T9Ll6n4h5rWbK8CqSl+IMxbnBWLuqeMq8
xhClTgar2HXWtXl14O5b++ltC6DOleD1ahOmwYcWCZXwVDQG4AoSzRF2jqnnNJML
CypAIxGVX7Ts+xV/AZMHnUz01PBnYnb4O287eB6yfCjblu5vpZa31kZRUW/d/9oA
5TTUkMQjebU0xg93bWWHLiGsBDHqRUlOQSdIyb/By53qhHmr72GsycEskl3lQkYb
gdXLEkqY0rVT7aBT//VYbfg2DeErwYgea4/Y7AYmDKwfsB7spsTVMoe/8v9cCRXd
v6lloE4YQXDiKvb4nVtSFF/eOKweoxYba+60MRxGOwlKNT1l97xK/TxER8TwPTNa
0y6aInvMD/hdlSGg4dIawaK4YaKHBgTAIDyhRDs+ItizoJ4OzICI1saprh5n5iXq
AqKB2vFfS8y+j8LqxfUqAQNPv1s9mZ021qakxZqKA5c3NqayRO65dcpkDDnFULTT
Mh1B2mWA/d6vlJ+3tLy1p2fEIeISFcfWX3vGb5A24kw1Q+x8O2tYJtGPnwyYPxDA
OLJA2xARygo8mONAlI3rm5d7F8ZMbk2VZRohrnTBfAWch0pDB9e7zdToSeM5gqOU
VejnQuW5LOzyroD1jYnGtw0p3FeIuCNG28yqF2EnyrHNpKkZvnNVjRKY+m/lz7Ol
YjDQBxc7kde/s3pjx/mQFyFc4vF9lSLfybas+nMVVvISViOeyUq6/d3lhjyfasQS
sX+4y9x0rRy3t7TLkhSyn2MxmsGZ0n24DHYuPwyJ3nolHcaBmQJNx2NFTfRFUVWd
tp7l7gA2gh5dMas7HZggiQUqEFjpAJAkT9gZeDNABqiTW1mzrZJj2+ZLaNSqtzai
RXx69Gt+KWqi269ckyd+B5gdkMah9b6Ur365rtM8izKv/I4HhIkyneVBTPlvgvid
8MRLMbdj4fxpLJfpI0wy9Cvac+b8JeR33i4fX52p98YVGCco5MYQC54GfNzduFCR
pZ8f3mEDb5BDTRBV8Mbuy07lopVJtmDSdpf3PQFmnLucYBAmrND3GHj+4iijjfkQ
dbTyxA3OcbtH3YhhaPf2FGQxjBOpURY7OJHSasVnyuAuVGO3zo1nmNqX0cCD4Uq+
/s7gOEN/Y3tiYE46dMyC0l6l0IYuJqIpouQt4RIpNstZZZSjqMJ1jeukeO4YNC4H
lPYFVNi6VIlRiZEgti/+eEDFUm6wVMXQMFYBEiDRhBbvCYnK9+QL8sDzyhvRMUvQ
DBhu/IefBajwe9/dPR8LMH2ims3OZFlO9FIg0dwcsSXXBcWUuZ5h3lJItCl3F5EX
1ez4miHQ8NNiuifC9r8xvw5LG3l7efYXgbANOc74fgigiXqFJEb/2UKBDpQI769t
JKMR8yv+8T9Hk0EY/C9TD00U91UnbAWNfRF4nVr8GaJasXqvYZ3x+5TgRE7dhYxT
KGR0LgYVmWHW4PDBbxCRMg+yiCgBaYtkXz4GU6X4z1A6WlgMFGZHqspCEISLxogA
S6mdJqY5pKGfeni89ruKfKHxXE66qhAwsZVOjCZUyA4axYqLqwVA+gl9WH5LL8x+
ZgmsC2cSFC4tWUBOFOf60wdCNgOO5R453uiqa7qOt5q8TZhIzZO7QzTLurzeYSzR
hPDfr3sDs9HzUzyhi3yaqy3PHhA6tpHhomipTwV2OeEdxsQtIIGIMA//B/l8enbh
bY8qbgNSJNLnXZjvokhsaZJJPp3iSLHrwAVBrAcfuFGkzIf6XIZx+NUhmJP68aU2
D/U+sSubPXFBRTVIg9JvsXbBbodNXVgblE+w7Af8e1nP165I9pSRNQfon3Y9AarA
cNTaLnNS3iqfRlWl8hWow+qAjQdDZi/7uJ1+DllVY5ERECqLGKdKI5rDm2FJ1rzp
Z2Wmucu2T5iTHfVW28nqIJNLAN5zlackwM/Dhv9uw800RlUxjgV60SvSpSJPHCKj
/CPsPnKM6kBnypTY+vCrQittf969MzwrCjxWZ755Rwvl+5EMz4acYvUe4R9Ag7mm
o9Ayy8/i44a3SjSVSA+ldlkrRcbUFjPmpB/3DWt+2AdRFS1aI5atXWeLQIEbMsKi
u9KOYv1w7st1jndzQJnn+S8ygjfEdTkrpZtBgq+Y+v/+3PBb8cZIJEkXITsUWWnt
EW1sX43i6QBPfaX8ikMmQ59/rSlWSD6DkVPzb1ARddlBsCKEgmfxupB/0aTgrOKi
nPrZ/K/SYz46qs/Z+wWfu0ntu1EgvLcu2261wq3jbgIrwFsD/Dm8e+1JVXeGLhjq
2NcpS0RZ1vCCM0s7juRITj4fEWYWJgFgT/6lh5sJQFgKr/Z2ODr9KqMV3GCj7kSh
q5IXS876ykDmT4fnmQ6FhvbbGx5N2bVtPaiG7mkuoz1x1BWbLiPelira0/CNizTI
SJ49ppzEnRnJX9epioixam6BfBmQn8sJhrSrq1i3CL/jS9SYgS6DpSr3kdw8BEMv
A6ee6Y0mrOCWwpRhWWbaNU/C10SFWQenLtwIqvKVDtaeD6ybH0R5vSm2CmjNfZnb
Af8791D/DsTTNqpFoQjvFhVYFZeKXJuRIUnUeSOZgMRbyiUrG0rTfzTalzTmfcIw
pOx1L1RCfCj/P5t48GVXO1KonfgkBCEhASgjZDTHDLBClaU8yEfG7LLvmEcELqn2
IzG3dr6guZ4vG3iyY0YbGDv+NeFuKau1pLRaBhi16bCZLRszxSmqVVqfqmtv8wjt
Fkxy8Hb+oSrDo4eWkwJBcwRgFwF0Nj0nfGIDo/3LXgAgQiJfebwyUsniSeySJL5G
rWflWu/nphRQBWMyGgzQOmWKZKQu6mLq6fQKLBOGpJ0tjFpfZeSiOKxzt2qQsvXG
4YShCzp3Wo2eNIPu75JmsPgZ1QKRmsGEsUxLgiXtupozGJDhR2+z+ZpNwkuPDTvA
VgXdrKZkvqv2O4Ro3k63OpJMRAMBH9idWN42xJLT/OfAoH2SiOJgIjp2vVRo5DAl
F+Tf+hRyUd2IWx3QfTLmGmGwrxWaPpCMR5NLde9BeRRiBzbAGSjGe7fUtSTvHg37
YayJaBJ7gO/rdRdcN973kCiNnqfYG3v8B3laaTGRM6zo82VBIVythqHSkU10CX4l
mo6CYGcdczr08ThCObDxleI4W4D29Jo6TGWpJdLIFO7DJr1y+FlC6hdmOSC0g9AO
OQOm2xgkkO6RpJvgZpn8lxzlv21wUTXRxUfU3roGOm7y7d8CkgfEjcyH0yGRBffC
VdnQEDMY3d2ihGZGhXA3qXwRnVZNNlO0NJ0txqu2PgP4Rl1VXv/xFK0h0x2MTX/K
0Bvw98RwRcqMj+LQujPSNz6WYJp4CxESaOrpL/0kWefqNawTy4nAPJlIyFvtP9bb
MoDiyZrrySpTGfuaEBkRx94MHO8Ody7fO/vEE83qAai7cHxLdt5A3zhBs/jOiKw0
xnxC9vSm2llu7pQrvIUZAlXqxPxrTfNmTmtiNQ7jHK47ueaDH6x8F5u8o6lLsFkK
ZQJSsmTUzd4H8t5sqqu39n2iGMGTminOtb44eQbKHjkZtAkWKykNtoRANL/qW1C9
2hpB02fPv4oW1IdFgCXynTCGMHDmN/qO2quCIW3blwxQ4g9D6eOgX94EgMaRrgMJ
XAj3SBKiWfGk77yPXqywf/QbgSmghIlWyzzykGSaB8Y4DFbNQrRfJCkxvDQS2fas
GFyHXC9g0MTjrQiTt7DmMpAlb3i5AG2ZDFohBjIRRyvo4PBrFUGwBrmnqWA5lDom
PpTPCCfxdbXetprA7gc1vkEm1ZszlIEgL84xE1ZviOm53ukbBg48vP614fk/2+s3
dkkWO+B8zOlqy4VBMSDpqEakE0FQ5N6+Z9kAY1pXRNixAVoJHRSu5sJ48zf0X97k
jfrDXUkgUinV6oGPUuvTt+uWlpI5G4gS67U/njZvhBx/2vewpBzo8Se6EyIYxC0E
SZkE4c0GqR5VdO2wt/jYqqtfpFpTI/xBhL9teXh09lrYnt7DJ3+DSkDSPf2rLCn3
H/YiWgHIdv1ICYTRFUZxj2k1G3AFrVLAAP0meKo8xjPBLe+Tf4dVRyacHsaOfRUh
5izI6G0RSks80/aZ9p57U5uyn/BrNl9T6wUEHP+t2/tEh4DxZsET42EKz5bY0ubR
Ots9JvdUjoAQ7afp1jxrAn4KFg0wMtuhwrUt/9jDO5OInDX/iDqtQBkdLXPa1XuL
UBjuIUpGqQ91koMZZCVLw1wvg6AxZnHOhVyQ6txPkQNc300+kkDBriGf2R/su6qX
8rcrfsyVYinl72G7pcGp+wK/QRISQ19S9Cvm92vQ6fduFfMeGFDctVhoRaYJpMIX
+w9fEU7o9c1KxgA2yX8xQ1tQ2oVvWTnYqI6IJA5jBOalBzyiGmQC5TM0WYDUwP77
Wqp/yZ1a121KmxF0sqjmWWshybhtrXFeChwP6yUgxNQOVDOYdSEt7VXqGYpEA4z8
QV6wFKaD2+UYZVL1YGLvSCOjhYO0omDBjJXgOOxo9k3pApfFiPBPOxZvTbkIU2Sk
xabvHK6YbAEUCvp4GNiyvZsMZaMAy2RA5SmTgvGpft64IyA43m5UTIv1xMkAVA0p
e0x2rgNYxqNqQNPeFzSixPRhIoPNT0LMhi3DK6eucCEcbs3wnjW/+mGSu5VPUgI1
xHH81ZkVMDQjIBTlMHuGlrPLgvuK1UmuJ6USGASZiYJ3Gum35BB/BXjO/j8ohBvE
Q1ikWgp1OY/G5TnuM677UoVi0YGtrGMlYCStjMhSzgRaX6QcmHQE29NUcHnXE/rj
e+xTa5Hj5rQrQylkRuSWzQKWDVOJILP29PCIkHJcpYQ5W/65QiBszXa4nG0pciqU
6futjcLRgvLhdAxvQ0amkCuwUOCWfjAqKoVuQdmrdCEPsYGiStpFSrgKdmWJeFkD
hTlkn6SVePbgGEbB4j2z/AeLoE5via6wep2ilr0OJLH29mOdxEeaW2qUwKNNAZfk
4XvP7uOkYrkGTbOpCwFsiaga7J3PXqWPjGjnV+9k7L53+pDsu5m0DgDcJq/5DqSO
a4LVB1X4lPAtOsVxLt07NGy8lYPbHWI1axepxVIiHYhESz//+sKTW2C2Lz0RaeDm
AgjfzFSSTkdSAqX0ijntAgMY4cNMrOCzaDvEkuSANfF7XTEZL/i2sL23lBFgS1w4
kKcn4EcWyhOb16nL4boEW05Ed5867wuHBUMK+/wcoSntSsrCs5J3l0UI9rr+EoIL
fJVsXNjYWrepnsM8qKPmyCKqOXy8rn+YxUo9J5yTMlNNiai3UaFxC6/r+a9+au4G
qu3VKCIjIFeINbNP4sOtcgDc+44Zlgyu+uWHWTpb/O3gH5iPHaLkzUG+GElBev7n
v7jUStjOIMZTHH8Csixp2nDgVqfa22c6PCb9GG8AApkeVJ4yxPKDvruYKqiNjrgx
aXhzyT3lNQ3EzAjeCPzsRmwMv/W8ttQaC7ZCdc5c2WI0Oaxg3ajsiOHN684eBC4q
fGhdAAP3cb0+iJO1kg/XFfK0Jq95pDXR2HK+pNy2CmhokFGEJY9gNyVh0riCaABH
hS/Q7r95gk/O24oW/kQpUIlxcdmTDQdgOtqB/QjIQ+xrd8deQNF8N1aOyNPVh6Oj
q27dXPc2kHh8igAKuSHESKB+N8zd+/IP+uuvF17wKxhUs2XLTnvtEkbXbKO2I50F
5iony3cOsePJfog5UGDDFelpGT00Jnf0ZS2fxXLNo+Md6fofJ5ZF08iUI9PVqcVs
Ee2ARDYaP1N9+pRVQRMLcHGYem6rBYNphzVCV19z96W7KC3U5bd+65WUkJqlw4Lq
uGDAPTspqlTzOeL3OYrIpjZlp28G3Psif1m43KGYfLPVQZQg0+1qnPgm86bRTD02
yf+TZXVXQb09xZSBls/skHsmNzkBUm+1mPm06ClAqC7ZoF0k6DQGHPyopUVgmKhL
87ndflLVfmDe/XN6DGPT+vPzyRmgu0U6vjh0kKPfQSvajGR5Ho9DBCDM7B5Z2x+7
jJZmEp6chpACFhOkZGTLdjB9BbcoHAec6O7igyPdFrTP7kOPqdF0CJetP18DsKKu
Y6xfUDGXe31YT2gjRVPlGhe6ULFcScnV+kQ2DrK2zfYIvduZ+mJCwELV6lMLJnAE
KbY2KHxeWG2GOe1RpyE5cC0ujP5EVl2adXp2G3DdkfoU7fDiMwcKDeZGaPq3f+zN
rac1oPPJsgRCG/nLGkdqRonIzbMJujrB2WHW0LxYWBh5B00FQARvT3YNQxvqy43I
rQ4OrVeT1OeSZA9gMqN7MS5cAkM9bVObiFCtF//WgJo2ooIiJKogVtRtqpPCwShD
g0ylFqbUFWXxhAMaLI/gB6T+m7XQYqP8J/aCz3EPGBVaSH4JUVa/LMdWbKfTbIT+
VZ/cjRH74lfuJbRyiGuU4G3Sk35cMgn7VCeEI6yB4Zo2C7xR8FhsnUUDN8je6sbQ
vgC0t1bMpSnMHHuKl3BbCHXyGo0wX9GHB14DiuNOrTIDYXAHLxtqELvB7vRSMHT6
2N0t9+d33BMyk0NBP9IZNSmlg7OlNg0nRdlG1FfHQZYxtHzbBxjfwBMQUZ9w/7bk
Csa9OqB0onDB4c+W1epxsUBl+x8YaYuQYYY4SoDcyirb2ehQDVoluyn+1t9sfBS0
/XgZ7YjsmAIMFHw4UEq0rWcW76/F4fP0tsNO5wl5ohh4Nt6eFPX4Ex1QBqBpMWip
Qfzl2ZBIpk24V4AI1XXpnHBf+dtapQvqh5VcHK+/8M0eLWtM7IGNuko/l8rUMz0H
TsNSicSadpD/w6QDjz7g/JxwKCIr6LIWIvjM+9Cyrh5M8j1eGor+t14nUO49xwIU
cpXTsTcsYWnSSL1w0rVV92bSdWyLTs6ebRdWI+latQCryA6cHPUebrczUc03QVLu
tW/rvJwsvLP8keiWbtCna1lKHJ+MbduMYlSO0ERF5AnfChzxV+jL4iFlNVX5nIIy
m/xPZ48WuGmyGMxCjNAO1OhKbr4lGjKVOkHRlkPHsKAW4/HXppoOIujCSrtnbrN6
ZhAYDAal2plwsO8ZyLQ0iucV6Q3AV+7xaQNV83cWCMGMI0ILwVY1nEosN3nmpSR6
VrMSJiqiuaVAOyIUAJSjnW/wr0TMuKYjZBvhVOBhWqk2hZKVG3vmSlPdTzyN5Be8
CVtL3IRyr5HbJuAcrIRwz5lWNqHM1krpb3+3BiSqT506oj2QmbpAJ7NvJpR2Ru7g
kDfUmg0dGMA9cfXLchX3I/D906/pTnnFR4xm0StRsd1suRWEXwlhcG0GKVuCcOh/
ELfJylcROVTl8kBJXqmmp+HqXw1kK+y2dniVoLwYKQEfCPC3UGMwf/fQRDFk0bUn
KE2sSblumn+BrcrQn8jLZYbJx+nHaSefmLSipG+p4LzFGcKd346M3XkQk8B9aMsv
3uFrx3CoyfvjTYPTGl2X4km/PxnXtgTMzCTD9yMDF8wTNfgctxjuseyD4frOJywR
irVcnLxuVvCJh5zrgzCFxh5xp3IK1rZyb/Ct8yffEOBYNmlNNl+0Ymn9wgWmQfDz
f3J4i8ay3LaMg22Kb9mKl9P3iwZcK0hepL4SUk9sOfy8STd4dM0UoziYjho1y7AE
7iiAAjl8BkvSKHYuWZSKIcOd3pFZnSlD/cLbbgPhOYix8kWCIipCrKGeeZxDrrfV
Do87XM1yIArIV8Xe6OTmqs6a5cXTLJ9YCVUjqzsa7NBR7xIU3+JBN97rZQCwHpJr
m3zWbW/nNDSX0ohRsE/JvVfkHcAxqvgLECzci6bGE6KwAAL80zWC1Ww788bjSxsS
87Day3yuRjGxYqgF4ewigWidoGHBMJQ4QWIVmehagm9s3fx8gkZqVZJpZch+RKBd
QSuZNAW5Y3avKb2zGa6Z00iOXPdTgnEE3Vm20tfC8eoBcXUD/OpfYa6xyrN84l9t
EcHe3W9xZ7jXx8+vicpjWWYn/0+7MuHPHaWi6lYb6sK8/qzFIT5BLQ+UnUGEIsWa
i+WE/3Iy1enVOrqFQj7wQiEBBdbevuBfxMEYdK0b2gNQxTDQtFa2m5YwQvUlrix7
DQzX326o6mVgE/UqTuLzL30p905jX0pfJXlBsuN5DBNj0mOPfAaqeybfLLIOcOWU
i7ks55K67RNsmk7Ri5RYb9c29DWUHaloRAufT7JACq1EooffWHm9g4vr3XuOdP4h
OsJLOkiZhLC0iiiPT1d+I5mI0AMCa3n+AYPauZ/czMSLA5E6rbWYREVFrbQP2kG4
cPa5drZPZbVVAZ11YITffx6gd67WfK5bHE3n3a8pd8zK7QnSO17IrwFBNqDveBhB
OpzfeZhu2gJu5cpTigDEAOcrzUhpndObQtBWIfQjmSDGRSHgGU1NI89UG7H1hC3A
SNw3HOjkYmfCQdFVgxiBXphl7NtRnPneQ8teYLKE1SjNAQ3vBIXe9uHWuc8iUZHV
4trMfnX3irAY76Qy9S+s5z5waNA7nmtucsmmbVvu7zwmGrC7HojNYh+YsbR3XNZ0
Ygcho+dKgIQt3gBEdt/fixvhrIQNvBdRF1MO41d5/o9D0tcUgUnEdK3+F/OgK+iq
JPj8tE6o6RbI+UmFbNckrmG1Z6VZhXNZs6LHo5CMX8WfRnbxHmydQa/V/GxEkOSv
3vEBBkuJtASMgu5WYE+Z/1GfvJlId27/QK6/Am721sTLtkgjpPw4SQSJO/2WNyi4
PTjSPgdNeUHfiEKhXFrx92qGFI8Dgi5yMSGJo64wIiFTpmkc3ifMmzvqE8dQANX7
8394wIkCvfJdehyy1JKz38SsFw5djgyJkp44IeLVyD6rXEFHrj83fBDIdn+9yVoy
SaUJo9HkZJoVQi+AELe73LoapVLWltZenSomX0W+pZGWK9HzMnQsLF0lYJDRqprZ
E1GuMrw2YwFbW63pfceJwVNZPZocYYzX4FcTPcOvVNOJvw1jk+DpndkPR/vQ4PuI
nyVDHcUbW6nfriHxd2u+tZ+uvke3aCX8xuIvWpNeGY2zyQS55JX3bN82wcnXDX4n
Ra26gT/akFBm14TsH5qiiu8eicwR5osbgCBVv1aBTmPPrMecF/T8EfOk2MO0h4hH
AnVGIPfDEVm1zTqgkaeMkH3VUCSo8Bm41lRWv2+TbrcYSY+8Hqq0XZXuRw9C6qcg
cMkMhV2ruFSVK3GjmK6nheTJHDM/oM0ZRCxrL+um69R57eWxRQ+CLfnX7ed9Mvqd
RzKpumfsJQrQxG0jt4CPY869UHcs/3Z84Oi9o5F937TkJj3PNsZguplpYbw9WbZ1
PLPsYIfpAdBn8WeAoZPXZtfEb2USqOJ+h+KRK/v+2L9yb3wgurDxGBp1ssqiPq68
iho1L2Ck8u2tgDFETuvOQZshE3lJ6By34DJiR1IMDIGhDVELAHQUomzHODAbdwzh
pA8u3oFwRt8dM4c6NIi2R9HJbUOoLuJ1sY/Sj1MPS0sF5vHuVucqQ5d4LPgyjP8l
tUbYhsXmg2iv943heSII9xL9Vy824q04ZMXfPMq0lbJrf0MWY/NElwnuzE5fA/yN
ej7Z8QSY9o5hJe/fL+42j5h1vVGLoAFgEoJ7HWEeibtnlyOzkJqpzXjXlvIWeq4Q
wF3/hYX3b5cz01t8tPFTzV99kKcLO0WNYaY2+IKGxD9qbF9fBq1KFbUobsMQBwDP
JYfsvj8BFkEihoE4b/5SkveSgWDxUNhAOK5wfKuaJrRXLlhhoEoLW4ExuWliBWwO
O8VWzaC9ZY9i1Y1Mm/imDmaXY9fl6hr23ciJIk/cuTB++4mGIU5LaQaqZYERNLGR
2BiZwKJqJcW2jaSQdtJXLcVU8A81Y0D3rQ9zkyzhW8NRLzvzwVnfj8kgRMPApqDM
JNj83tGXaU0M/3z2NIu+RtabmMDkgy0FT6+2QKlCyk2oXHy1D6yhQzfqZMA+gRL2
dxa+bfjCZsvpMrZrK2c3KkUg/HH6c2/d5KS/zWsD5hdjXshoTIv5xMBvlm1UwhgQ
wwuS19LOmKGETYCwyoEeDH0oVr2wgxHP1NUy5N/Z1JGmCLDdwHo9GEHHKx+m8bMX
+80ILB3Tb3H6DpHNKDCmW75sIUhA1ujIVGNjaKFPZxdd6Ga328z8zbLR7WxluAmj
Q4KM4E6ntNTne4nnCAGGiazQi+WpHMkFG6LC3emkAq4xGYiL6pdNlIEOI51ohntI
HE8hWRjKJUhOaoVnXmnA8Tq/pZSQqyTk989vzy5IHg8GtjRdK9yrRnyqYhCdIydr
q6yCaDDIbd4YbrUQjQyuE5eBu+UHs/K4+5MW8+KHQ/W9wkSsiGA+Wa+F++cPg66B
38NovLjIBDd7hg9jceUPfXHk97riSfeZGWWGWFQvGNIj4DKLKoU7qhV20QGz5vrO
Zy9q9mG6dEwVeaDVVRRduDrRasUlQDqQd106I9eOKaPLsW2aiU9W3Ggfe47b+jxs
8H6krVGqFLAC8RZ98aeQ2C3mvmps8ZhoabyyxsCNw7BvjrShWQAZuN9UwdUVnM95
SsD2Eu7smfzWSvd/NfN+ElOE3GDHd0B/ebvUQqw21NWIyBtLK7eePphFWFd9Zs7d
8l7PXOziDOiIUUuuRoCj0OYWUhhSvNGoBn1p2QHysYE3OvnLEm0ng41/T2zPFsI2
iLHqtOjsx/KwDGqYR1QWveO5tK1gJXeFOq4o9ujWJWNJ4lOeZWU5FKVWePwzbUcw
uMd368EBaUSzkSfYGOrS8ZhaKPuIBZVA2V+hUritu7kYT61FliP2rCr43KXv+TXg
j/rKSBkWatJGGyuA71Y20WRpUrmKmnecYK3QRjClBnEmWkCRnVLGsLbmLk6wRdwz
2w8DW5giQWJDW+ut/p8dw4UHSEqGXKEOU2H4ZiQgA2sMchecVkJR4HddJvmm1J4H
bkBHGlMBwiUC+9pSdSjuOYCgGeriaQT2wcku4whaFjhrUnW1znCzVKYhZx+wqAqd
TsqF8oFLnYvs/bdShONE/PMbkPVUFtFMatBtqvanWuSxjE7+pPPW3mqGUJTESZ9K
wAWfHoxdjITmUK9PKjynr6R7fCvq8lH4sBaEDt3nM+S974f1+dKUILeZUTXNIvEK
j6Y2T//pDsm97v+7LBlU0o/v6kqJR4oBAV4zTXUH0F84nWxDjyAHmDCWhQoXfjOF
RlkHHQVJGWsnqqMv4OwNRLq90pO90fb6xWmF2F0/pvJackPcUhP8IiXt3gAa4lzp
kwFIEO52B1WSbLy52FrMLCJvzqXFSwg35tsgaE20qPGa9VTmpdgw5LQFgJK2Q6o+
OmRXIS8d0eJsw/7rDtOQSTxh1NLTaYPSJESZk0MKus63Lx5uV0dEeR8XqiHUudMw
VcViCqwn8tE1lRsYI87BohOuqz4O5RA7WzYrWxNCc2veD6Xa7ty9UtD6Xg8nvJZb
YJTh5YuuAj6wl+wuXYSJ/eExLm6r6nWal4Qt7ymdq6QZ8WuzPgBvYAZEI75EP3nU
wsJHid+Hz9hdaI+/4cWMuKqAZUjvXD3xh7ntvW4UeXK86C8RqXymsYSBWSxIUom4
u3zDG8EqGREqqoX48XgY104XMmWiSVT7gVPq4BooIH8fiKYnHMVIteDHBK+RypLk
KXQh2OUBjStOyvHV11SEQTjmLrsYcM/uanVx1gILLPKgenOEYbeNjEnQb7LhR7mM
2ob9cH40CBFQZ3dbHT0rOWeQuktfILxyVzeeYcN+8s0PHui/z6YVv96OA2C9FNdI
MDf4Q+FB9Z8DxoAmaqUt2I2GUfslPSo7rNlHbepbser7CqZWBeJp8fZF8HLw0QCF
FvSyDoGgHPJa/Dvmgk9GgKen79YTzl0fwfOinmzxn2YDajmI7QxvoaniyxdE9PEv
4qaesB0gArqIdDhug3ejj3dGOMqBmIlyPKXBh3ycdfJHi9g5T+ocTHEdTMnrVc0o
E74bsoDFigkHtS0ThUPyFOy1xw7gAJaFcZ3DQOikQp60cw4QKQkVA4Rnc6DBlR+2
/JDoVK7XeYzM47KTUbz7jzZoyeO5xcGzMuRgyiZHVKyr/xRsXs8cNN9k58TBvoS3
xpTJnWyJHnyaJ7GJ+PezIxuk8VQbwtfmGrX96Vs+KWzsrbSuDMRqvpSixyAx9tIv
QNf9IgbybIT+QLZGILFe/y4fvw/+gtUeH55EMDyZmKOFNzc5TUv+Wa5r27SCFgOL
gzuquoM58hYaK54AYQzuCuMRt6hPR1CbO7mOf0FdOwFtCLUaiwiB5Q8WiOrfzbjy
uUhgBEI0uXi2/fKCjeDWYmD5ZxGqUml7hY+T1L8PlHV3TSLRNBE6IVPA+45TkZkB
YksSelGoZrwYJxwidp0gbB1W/TDY2Wx4cL6UBwHDAPhM7kHlA3RQ3Y3+VzKbSxId
0mWcNUZ1F4kzqw8hIpifwbi2QS78de9b/rpphqv4icUnjMJ/AqlYmyPjZqI+hdgm
+Dh4fBxGAk0sYtH3XBgLZhcVcPSfFthfI2WpYuWSl1pXdY7aTSs/Dwfk52eI1r0x
hZFn4Jni29c5q/8TC+SEsLPRq831XSQ+t/ClAv1MDPShdPeknAH2AAMFuYE6OzeJ
4/YoF+3pH9TNvXBlgRGRBY121rRZH2vdbpcKQbTjDYSTyYnFRsCSoLlebztEVy4s
znEKd8Fabfk+dxQBiqiosnHHV28jNfSfBNIgiwTDip61fIqyRtp1SpKKp1HxOhHL
BalXMnzHWlcMGAGARVxanpwrScFuvxxtCrgU2AvzS9BrmTGJxeOWxtNGLuhLrddw
kVdOUKx7JG5zXjqPtQQSskEDYaiw65COmreA4WP9v6Mxfojpj+eEEComFd70nWn0
4340AfRiuyZ17vB2B5RX5OoSvn55/vLrMSG1ACjhXAyqZyU4gKnJP7fY47/UZL4J
gxh2ynQMx9wxp8ixca3fLgGFA1Ag8Z/n1HvhPMrOYnGwlzXCyMaNhlYIKIjAfeSO
tXGoB2BZ4rCkCzazpIIWY6VWcuMkGHDWh4p0/Pq4YzSyJOWUv9yHVKLfAvL/15XG
1G89/SzkpwxphAGzdVh1CRjqjLWFO0coYFMdzXoa7OZgHLHPzUpCIodD/QmsSRBa
GjdsOMn6SjyGw7Od8eIcM/Y6wCeK+BfYu6o1IzbP6puWq95gh7rJHPBD5eHIFGg8
8v+s89cmxbT9yPta7O3ENW2+XZqYzK5qRa0RPdh1zd54T5GeMVHhn11yvVzJ56hC
HiTT9fgwoR2l17PaKwc1lRZDp8TwPF4Op7UcfQTth4hZQk05xJGn8mRBuE1cIltk
Cuz7G19vz/JauA/ilBdLMRgfto8wJdTN/BBo7IMPwq2hWyksJ7LOB7Fixa/9CqHl
mbmP6URYXg1a87yV1eb1BzrxSttbefjYrkdYSoTIJ29zCfa1TROxrcQKSLjnpei1
b+dzLEzqRo3Re3LssdbGly8ueqqLL3r9NHIyTEiO5LlvkKBSTrDG/bNxyNdrGaC0
4lOOWyZAk6zwXYwFTBLdk3rMLWW6iwfr30DrvVEo5E24/4oljJjCE9KOQl8d2lKz
hfBkCA5wdEONB6sf1i6EHTQTn/xJCb1ocMTsDCx+XVbe4ooWBQlFaT0Csu+j+fLM
h3gPfWyV1aLfBDuURdQ7FbuLNUvQqRaGukIweQAcPKD64ZRB8knvdaUDke4LHCGk
qxXWvlMV/Q6AK/v+z41EKizVwuRDYmFllQuFn6Wpm69ZxAFd4UOr9MWdjppGjiS5
e6m3Vs3IViTtGzcKMD+JN1AhhDZp3lxM21tfx7fSsICXNK88iwxc7NndXSZjdaU/
Zyt6UBPrCsmjiu3HmpR40sjIlyBdvCstU0hWErVnTqSlDgyila8FpPAmnd7Mcj+I
F485fjt2obkRSDVCX3+naRw3K4WXZC8bNjks8ZdJl7M/1sMCC6mRHMpi/4VAxfpf
RTLCKHb7gK24E99d+eqT+K0b/ujOznU29sQx0NRpzz0VLu++jtdUFByCFjmtU+GB
Hr0Hj/WrPmYttltrIEQ9O7XxjEmoSAubKJh1dKaeULmVOxyMDG0qFpr7bbEk3srQ
atPsYQpvuEHIyCfDfJztRbwPyT3VGixNDFlQh5BloT4SXtU+EB6ji+OfiLRZGTdf
+0t2WXVjQLfddO20J7ksZ1w+/3YGZFqjwdRvmOc+2NI0zA0z7jDSRNtm5H25ifxk
zHMJcVR6dKDWPzb2QJqAeylVTrp7vs0r71nbvc8FR+lQUmISfG3KrrWDmWsJCbhw
K53kw8G2gWXE6mw2lP7zkFVMsRrgBt/oIk5aRuIg8apmjhDEkEgUUP+eQOe+SpkD
9FIitTYj3856n/la6w8MRbMUGC75+PgHDUY+p/BJJep1tpNL306C5XmRI1c7+c6L
uKmGFlWyH70jndcJ6LMAV2bDts+8Lv6VjFiZp33s6Bc176+zKJjenlyZn6Es20am
7iUT9YX/piMJVUX1LpchdGbNpMnwo+6u0r0qFNQqKw1MLAXwvuEYrPBUBXg/ZSO0
6aufhK+C6q5t9hvCgo2pKUPF/UZ/hg5KbQOyUzeMtiyIOuW47NKaubwZ/bGonrqQ
eJPRkp3LD1sJj7VkAzpOe04SvR3E6DKljFiL750l0N97X+uLPXfyRyLlKzWT1bSQ
i31uS/XOwfwo+uGF8FEbAIXAY6QYYvV4C5khaQzvxyzFQ/kuugTtOQlP1e6sU6ri
2HIvP0s2yrSs6hjDGJBFKu6m9Oy+wBTorqDEnE2kn4nqrKkRPFX5abCmDoknvlOM
JK+9kdlWCZuEuvmXFgasaQ8KT4XqyBlgdnjFPYFoNbvp04N5ibgz120qWKMQ+JyO
+LY00CgDI6/2UA/Jn6YCTCgL4EWgeb5G83LMDpKvzK9E6bJ6c11rYCDrRfM2yq9n
KS5xlRwxqxioJbKQOJfrsMlD7q5XuNge9cX0AZOQRzTojGzrfuwWC8mygMpWD1lM
/FNthOleTmKDlCWKdy6Kz2TsytIrV8cuUsd4RXD2e5kVLRnnMflOyw4/8G+68IUh
9ZqYqP17oe0rx2lW8W1U2XQkkw7m61WciISmiyoH/WYanOgH2+H4f94lj9vmAgaZ
BP52bxG+15dfGwySvrYLmiLmiFWDz8PYTuiXgGnb6RRjuM27I/xefun17CHsM4W5
a3M7+tiQzShjkMnMu5+73OhrJHkJtBEh3pdl00SjngMGfYUziQ3jPSn2swPSEioB
Ztyvqt6tpjiB89S6447MQR0ubeUSKd4ZM2VvrXGL8hs1E42Y0ZWyNh9SlhFoXwc6
ySbQ0HP93qNJvUco+1q3DV5qCxZvEtXvfKPj1K9I8ZgqZVWzl141FBm8T8tprXbQ
I2XwyjR2xWMn0/TRU7u51XFizNKkvvHsh2CzTxIVp9VerNkOq3KSi4Yqc45l7vWS
e8pENWLVYrohNriWC09zKYz3jfxCRDCR2dXnUKBD3pci2nHZ6yjpx4gmhUbKAFbW
Ts1M0mdsgXu0umbit90LszyJxkOcESSaVgmyviN9aWVlyLUaM9rWLYXB3GuCF4Wo
Xsxguq/Rg+N6xevT2PVfFJ6LsK77w0xABUhvJtFzJNuqWByRaYLuKO/Byg6NHtxb
lv6ECvGDuqY+ZLu6MJZ4iokM6vq7HF8bn2PWYrYVhJ+34AoR0tIxeC2DO26ocRom
Sfu9lhM3i0s7C/KPVI2CGzJ6cjrGFgC7gOX2j3g5NAiTZSmfJz9hOSOY3tTY+SeT
gg5cwwW833nvrahd8oL3wkcKrR0Rl3l6MUUS92P0XJPzPI+rrwTaRRcc3NsvtAwd
V06uIx6+C43rtYe8geF0FLg3CLRkybSjfBxapgI8qSW1rIBj+6hPGzhAWB0Wmdyk
2cDVT5z96myYeCijvaCP0/2lCSDPOco2OVekwVapKhVIUyh6F6F2t4fPp2jBGWFb
BtFtfFb1/q+reX2Q2DsxdKsDdPjPOWm7+oPMtcwDETGSqA6uQ7UhK63bhmUthiCj
lYI3NKBV5ZLaieyE3+vvjEplN1wEvER0T7rO8ehYcp94KPjQoBRua0xR36BG2xuq
wP+fqrfcjqf4CQ75bf1r1SpmUQqwqeFeILe3iAEvD6Tz1i0s5j+66Yc8Mzlpm6nr
bRpiQU8BdJ//LRfypIoZhjC3SJ3fe+GSZCtnnsXOUez7e5HY5ziR89vKYigT2j9e
7BftptdjdfrMz9TEVv35UjyEP2SLadlq72JLg5oYGfrOhkrEoQ15HT+jit71OTAx
FmSJg+Dgr2M3juVIOpjH/ew11QaQv8qg+K7hSRK5dm8uoGV9LRCb7WDWwBQQZowK
jRKvUuP5sawq5Gj2YYekB/+PM59b1CiWbz/1hASpWIldihJm0gqxRtPpv8Cmrmr4
M1jvXzGpcBIU+DMpyzUNq6Qz4stOlyDtsdhfYedFSYOQEsnOoBFpdlSy/mH10lRT
UwmzyEzOuZGzWQ/LpyikeA2vgvbz21SISNFVS/Uv8ZD3g0tSDLUfyIvGL/uVCr/9
13gz7V/VvuFEql5hP/jTEF0gpbATppWUvkdGZR8v5m816mNy3mOVb9TTbHE2KP/+
1yWCgj+Ce06CbpeaODerRBt60SIa9GDZDndqldafRtG6nxu0NRmf42zWKDaWUmX8
3cOug1Y7Yj5PAjf1+YQtVcGiDV1t2UfpIrc1FzLdXKls0Q42PdXTi1ByF7QTdAeH
kI6oD5E/BQehGhw8U5z8kahkaY89GQggapWD2wjrKHfvH3HoLd5rsCcK5/4XVuwQ
qg9dZ/p7crPxwkHgU7hgRdZ65Tbh4ZrtGMEYFmawtiNx0xfL1JBsa5Dwq+5535Pa
B1cFhs/QkhRxEjnDrpz9ENXjmbs/sHfZDUcXCd94r7rRFegvoI+8zDxCCMS5MeUP
hjErQ8oxbZGvKwQ9FFeep2ThKnod0yhPxhrpKXsAKJ6Wq5CBUmJF9r/ngG4IAI7z
Bebb2QG4micavsQKr6NHnMO6gOkD/fbt8wtvjo2MVTW7rMHrfhtIQx6Yuqpvybz1
6llm4kjlpUTysTUTsf+46RI6ZocF8EOgPk19vHpOmS/8DaK25kTS8S3ij1iqS5am
+Qc8DLl+pbpDPfC+DbWQpfTo2tKh5oJPbFMAABbCXvTpsXlDN6ynKk+klUQBLmxl
VlTv4BI1Hzchi5gCRPkSTddKUL7iSh9VnYZTVvNWKDuHhf2EGFMzRp9Vq3+6Mot2
Cf4IdwINPbJWeSF5OutE2xtehF0AbXaJ8W3G1f3YaHCVuXlqYG56qIWbJRgKmGYA
kZBXD6g4/sR+6XorUrjDGbUX/vkggwt6dVSg5VSPlBktH3B7PMUJis7CcNJFi4cC
+478t/ez+hHW4Uk72Sg6f0WScJ/Rl6o5GHnHPEBTjGht2y/V37bbjFN91QUF4MKP
tH7rLAWprE/ajJj28jsZN+YechkTStOHC/fO/OCpeVdjOtfn8F24PZPPy6gDOHXH
0EQSTizyjDvWE28g5oTgGKvEErUHvcKH6ZLyPSbP+UEsYqu12xxbsyXYauj5bXN+
iH91+en3GxGOX+uP5otKLE6+RgTCIjh3Wt+ewbrfTKhpqFRQN4ktAIDcZ+OKVf6O
LIuxQoIBXGyGy0j9iZxTkR2lnc/AgUdK0vDxDyoKMzMEZkNvtNPUiD3RZh0UyZjt
XX/RiHOF4Fs3R8A1Lo5+1IBp0WbVhTPt2RAgO249IbrKtliEWrypLnqR4CEFuhqM
h6TUTn5ZY1yDa6ZGf0LdmDHJa51p31bjIKaNT+mleWskMl+K47CDulrOtJrDmrlH
5G0NK+jkTY/kDvR97JThh9ZHbDrJjgaVY+0CxdM7csluFSm5rK0bd2CVI6in9EYE
3egH/yMEuVTpepuEwIA34Aq46FFz3Kbzc5DLIE/x9q4NOp1NyBYq1zX2gxVBaWsy
3RXHm8rULQMnH51INwfzIOwi4JezHCJnj0fPB1RgSddYY3hVOQKVaLDHdsunHuw+
GGLy69l+qIra0gEMnLOaBP+qnf4OHtPqkzgRZRIvvRwfGTY3NVaCnWy1MNuGmNQS
no5O89m0Ec9DkAjU5sLgRV3tW8HB3G3jLSjHU9hPJNlGtP7TL/QL5cLx2nHbtb25
WMmhjKq4wIwzXW2QGOP0ikRXAJzsyBdwnQzRXZHOk0BqsUWQpdW9UvdKTFl3RFVc
ixORv12Ncjv23w06s/YZg05Pmhs/ApnmJl3OLuLSaFWatT8El4sXcX76Mla7XUPR
Y0sy3UCYWOHycrxgOjPHu0W85JVLnsNGKS8m/e18LEW8LZ0aes2u0OoIc420Hs2n
xmR9cTymrzYelQeEcbLfCgXp60Au7+k3mVTfy0BexWUYAty/NuXE6KcGVBjl+L2u
qYiSyymIoRo/POLE6b9efHAvS2R6nSKpg029Lw3/ecK31p2OX5o32u8FtN7Np3In
Gb0+52qXMYu/pcuzwd720oMka52FmrX2A9xtlb5fVamhtv34rsNMSm2RnuSobUuz
SjDSANDKVpt5nhtiLsOfev04i53osD2UCBRrGl28sgob267zv59W2wY57QUkBENx
WvHtrRqeShY2YbytIyeDIHWFmtCsQjzKuC7s0HhjC9N1bgGRl80iK8qI+3WPhEdg
or73TTa29qqAaRTlwIHU0Xz5pfTfe6iELLO9lR87yfcHsTxGyLuOk1c80KPPovNg
DDX0WI6nve8xibYsPX+zIqzORAWUbvginaVN3DZHclY3nh72uouhp7CtY4wPwOrD
9UJqYaRdM1PtfEQP9Nw5HzDdueYWVjW3134gLT5SideKweQ83k0s44MfD1fdA4XT
Wp3/hEZP4laTiIldv5zn8UNz3ALqn9s/TgnUOeSx3s25Wui6OOXvIYIkQBUt7SRf
azozF7WA1RBzi1+UP0yGxH36BeX9fpWS8uUyow7lBbzn87YrA+izkafVCLv8IbEQ
thx7CVbB8MN4JzA3OXj8xHiRgmmLC7HEGg3tpHvZxczeAu6XBRZEPDHWovnMN0fO
zbJfC9d8eo0Ue8OU+FTeOWTBcd12XhRH19opVIHTl/6Ls4y7YF0trjzoSGIO1hOB
CNEcn8H7AsebvUT4mUEpWN8rtbMK75fvbLOr5vWsl3rl6NQMKsSCTy3YWPA11Wqo
n7cNgJbZWKHM7j/tcBkX4skb9IodhDJPZ026IhXq8XunXNuA8pcp6UWwD03azH/I
BNmYN2azWKGHyNAL7unFyg98fBzZ7hq078pUMGZQLdIFg4yAtKBrBK6TgSo3saNa
RyLAi5sJHgu//RfrzzV1MmDso2PFM8g1yLXOELk0/ZBnlaRXEt1CtMIdMuKE1ao5
YNnFpyE8NBrPD8KS3DQZVDU/ITTPeHdV4vpgSwDb92hPc6OHF5LW9298EsKh/xqx
qFnbzaTG41CweU9CIR3NTV4cXHrWrkWGxUxGtvVZsB7sD6lubE8KwFOaPndrdtm6
zR/VhCuyoMVS7L4hFKSAI8JNQFtLAjW3z28179OvQbPBXaNIL4/yzpouWyQlcKeL
pi96P074x+uTd04XVochLFBdDQhgJtVQRxy7XYYv3fhLZbBKxol6EzwQ9aVwEq4u
sUJMLYdr2oastS1Tgdw6rI8Cw4hA5mVB9r82KkcJ0R3TMY9IYAUXblSBZe8l+Pv2
6mskzzbylBLTA0jgMDrC1PJ2iC1zpBKZFuSn3qxkn7kwYQ1d5JCwD+XXns2heYtk
w9/egnHqNxrQ1A0oAPWsrYeJr1ijWh2DZkRvk2AQgrZ0uKOz6xypfGVu0NPkczZf
8LUDie+Q8jOOGxbtH3dUkO2G1xCTFk0fk0VqTw1xdKzCqPE+A7IGS+cYooTPtRc5
jPncAR0HkciM+gvvfRSuu2rrSCstilJCutqLAtRRCXQ3jxiDTYMvlbAOCkWj5iq0
h5UkF3x/KOawFKo/Sl6EN7bW0DKacEX+y9WEOTQT0FUIorZ4pHISWm3ZO9gp0m/O
YRMOgHVZeLaNWsdZqGGlg2TsbXFWKqtxQaOBykkIrKHGQok/7i6p+KUvLSFL2BH/
SzPwU/hCxVqwYVCfvnvbn8wIviZoCRkgNBrGJbvQTXM0YTr0FDb1W3q1WiTi25/q
9s7U85a8iy79Vti/g8fdj1BlRTS2AbayxqX1P/D3gmvTlCODfHUdQ7/9nShik6qX
9QM3LfhM1+TWd+tUfvVVaOy0evCVwM0/16KdUbgwBXKgvrykbhUEIXVuTusuEexU
JakyJCWyPBYOVd1blEXDoJdIUSGs60d3ClLXH8aTkITnvl2YnUrWXbB9MkO42wDc
DZ1F9lwmEp+LnFOz9uds1YxQj3/0WMAXQsM5KYFu0voPy5JCPztKPS2yE9NrPVfQ
9RZGI39gAlvUBUJjETsALmPuut6tW1m5pyl63R1iFqqGOorErlUgzhs7JxrNzyOx
CtuoH23QdXYRCragIW3mpSg3FLnEClVN8SydkOynLADHr1GkBWtFBdppIvKYX9VF
c4fzVJ+5RmThi6Us6zb+m9tRo4U3WhiHPo3IUKwpEXPNLGAGPTPA98O5xnIkt4DH
XdwVKULBVhflCVCVDi8B+hZPQoNECCv8G2sldGeAacl2g8M/6Y0Z7NQPu6/a+CeX
GCVAaUmvjObpdsHoQ6Ud7nnv0lLruBINZGckTtDKzYv8sSXMq6cJo7X1sifwVUHn
FcAUrNjXPeL7IhaZqS7XId+U/g3gc9N28hVe8tRCMCQXoYsZtkHzavmQ4SckUgd9
y+oHIhhFNdGhvv03uuy+uQ730YdD4HNkyY8FvCY7FKb7yjOFfUYqWLsTsbgNldVX
V5nus4vtH+kJZTQG6j+wbbLGlNyCWhdHbcDGaxwy4YLsFY6ZL6bTwhsOp5ditZOK
9XpRiJBnLwt7f4rhaw8TtQjO78q2u+SYbBpQJ72MmypPFIGrFYJ2GxsWrP2OZpem
RWu7APGWMuF9Sbw1eiOs1sywqrzvWN96nZqKaRIQHxPgBIXI44HgJJPfI9g8fE6z
uV6tcnSB70IW2E7BxEmBLiHEF0UhKtycZZOVosB9t5xLbggBmZ1FVcJaF/wPyW93
jZbMbeFFLZLpCEqxwqAndoDo44RZY3y2Rrx/t/mvvKxR5aSIgkj/5uz5ahpmBK6L
8n2tv30sgVyun0VDcP4CZpG+5CgUxtoeJWEO1C60VV3KO5RN8B3YtRpywRqa8WCz
nKZCM0cn66TYjaFmwcU8W97lqyUwkqa5eDqrwWb39Kni84h9V7pn3a7+AkGLSiY8
p8TLvq6QlypY8iRTfH5UmEC+m6lVAldQ7i+97y18iZslvONv51EYDXI6eosI6qbB
WU/UM4MpFXnBbnfQVBY9NYugY2qQ19/wcc8EDMyNo4XgZ/MlbDOCanIE8fTxu7pu
h2TfIFEWXzn/m6Y1CC9nO5rbL8sPPOZjgBmNFcsD1C8EZmaLif9IS1fo8Gzbsjiy
ceHNnfYHbHhEqtyh6WxC4ScuIrMaYpu16/LcmrXPgBt0F5TWv4o/C3VtHmCQwEW6
iJqfN9PMhA9IJ24Al8AQssMLk7tEacxQrvJiHZKXPbzNfEclbKp7YaneZ06aR9Wq
+NjlIKIiSzep1alWdEH1G7u79NWxwLbv5vMbBG/RMVoQbgLKbAH1SiUO3384Qx0n
kM40XifYyRHbfmO3wvum5E71/d0uBML9y13438YARmK1hOIDtopAxMsLUMWEhYeV
RsERWdzh2VBiNU8XOsrlgDx7VOqIC+UBdbHt07IFf3NTcmQTmbYGD0WNTztouo/q
ZqaXGozAGdDC5xce3UgXkup9uPf+Y9DO78BxJL62toZRYeeZqniBO8u5VQxdjVsd
bVd4aCfM5R1YUF+lLAz33c73ZIJBwJVaMZnGS8u//1Fj5oVjy9zTX6nb0fTgXG8q
W6aRGuqsE9weJkBZQNfi6KeshqE7ZBNkURK2QRPsQL36+as7tCVWbpkNUK7f7QUO
fyzTsT2Wb3Tv1O87OPV0jahRDx2usJSlamg/yIr1kNC2Z7eByGB7Hos33NG0SR3/
JMxwxSCHLXnTxnlEytnRCJyPqf8FLNSbvRKRBlX0hQsXU4KTIPu70dxE5pNdmBzk
3cy5zIiv8Kgcr0Pa8UZHZqaT7JszcwmOWhRE8zQjPSxVJBnH15TMVK0YFIo+lvwk
yLL4gaV/U/QXhB0w6boCGWhKLmW7O+MHMirHlOBltt96Qk6/kwft0ZzCHXU6RhGn
wh3Ljs9g0tKYa9cqDmvIyaXMLOK/9b9yRqrwN3ShxEayuGVKNGTaNUNId95Dmly4
OlYpjonR159RNuPah6hsiHTpfAL6mDeBHtKWpHnBPpov/2YLuuLBHY7qG4FK2UxO
H4ubkBsN1rkQwURJFQmkp/T4cf9D+oz+u6stC7xtoW/h8ZFRD/65XyNLzlEcsO7G
R8NAR5h0VwM9Fj0sQD2roivsUpZAvACzbaEAtuzupmfc3IDzL9vlNPoCA0xErVh9
T95/+0Z2LrEvFecyBLVbplBNiWkNP1USneAG4cAOPzhGL8DoEuKXBYl53rZGMH9R
85i2p11cIBOChjZmT8MLP4qiXqDwP/ynpABiBVvNoOcfjpRpHn4LDSL6uyN2lgWd
0dFAXBUz3ZzbH/TOAdHHbpToReH0L3huk/R7Jf7YxLKgWUVUD8sV7MWATKs6yi7z
qfagNtJvQV9AhnRNQCGrBelUYHm/4XBQzQiQNFgo4UPfeTIQhFTmiCl5/AHdkT+D
aRi6hVsxj08t+xYLdZDPiY62YsBG3e4yIOfHhVcH2KHfDYWJDICBK/iaJiNKYbHN
KFsl5b2Wd2KGKhbbmaMed1HVvxueWlUb636eExfZExOm2wcZx2mDA3PonJ3QN6CN
fkplQxfI/zz2atFuiOABX726cPG661BCly8pAP4PK6Ff4HBR2m0UnQe2eN7uDRKE
GGE8iVWb7J6YZB/WSA7JglXrodzVg65/esKudVuPcZRkbVGeVSl8qGq5TQMxN0Om
2b0tx/yNbr2eVNxgerKSquZE9Ds/TUoXD8StoXW6mIoYhSqOhHd9h1BogXp6lecn
cqV0EsnN1HmFlApoZoR1t6P0ActtfWDrt4L2w63V3dYMLwMCtS+cJc4Bwt4pT5x9
sUy6XFiEZzjTViQ5ZpKKo1ufM0iek7A5Tznh7JhLnLt7vkWTEooYXwDMb+6kOyja
8C3UOjpTDFXy4Vr/cV/0nZVfF/GdxNwpxgEyO565kH7XyZupeFLls2h2NGCcITlK
M9LKSSq0gO5sf0NPYdz/LW8jcVlpJNoAu19o7aT3d9dqKbEFRK2LN2YT25rj1POi
Vubvh2PgBKuvAufpiHzbnvYmMYRAGJocRpiWMtZPYyOiZ4xMLBBkJMDWWmjPipUF
FDKaeyWXAavnpWqmqMP3eZeCYils9of6mramjJgDXqrvRTZQwy8voake6vTMqrP8
WPCN8dDWvMaIv0jtmpHFqU8/hffNiVz3L/P0OdV1RozqTWRWCdScvTXQjfjprWso
wbQq+8KsJHS42eZMKwhvrqezeBNgmczZg2PuTdKYXQvFPRqiPip+P7vIuW4rcfSK
jiLEHHXuostOBzSLe+2fWVaVkeXw5e+u04d5VKvHCpYlPLBo/1UudPW6bOb2CniL
sXO1otb3C3SOQ6VbsBPmLiqUp5xr0M1zbkogNuSyL6+WW3SneyWR4tmD78PliL0L
cnbYQ4YCEnxQPgRh4GBVPKLYDkgwb06vCOgvrVQE8hF6dBHtaS+cPmDt4jKT7RXa
h/J6zqMA75k3FcXDBVUzbrDQpT7FFc9BT6S2LaodmpaTs89e7feHMhETr5qiijpg
AThJolE9Cc+vbly7SGxynx+0SEUySuS2GfLODk680dnGzzUkyVgMPr4evwWuMqRi
pE2WL9aB8tEuY392M0ZKXJrD4dmiuryClbbdaiDYTpnDd5yxgk7NM1u68ZqMxgkm
EQ1YNsSZP2+oLoVZjwF88hIEjcn7I46VzSErFoz7b8mIgaaxbjnNVNWumJqO8FMS
8Ed9p+kv8/6bGcJjKH1xlE0sqoxwxU0JP5UozoXq3VnetCB7g1PTh/VSWoFcta86
UMshA/TlAkLOJW51JY88lUq6NUner6mlJSwV5pCh/UlPRl+5YMuvFsEXVINEtZ9I
kLj3/NpKDmRiXqXCNmcpHfGue65FBpnHQFV69jh0KnCHr/hQ1WSfLyyyH5hDUloE
H8/C7y5Qnfm6N+VDrv73XJj4B1isgy5iy1usYFE2l8ARVNzGnUCoIreviuWl/87K
3sWByAr1mTTlCjV+jNLVEdyTXmDPBO6WXFtt+8No99zmtZ+hXh2TmX4iEETEjAhd
mWhAwEw7EzN2DaTZ9hGjt3SRksFRYsBYzjeZORlHNNEU28ixFBnz6KxWDwft4vIj
yoFZgQ1/l9eTGktMissngox0syKTvmDD4Fz6+S7S0VQHRmzvMlE2fTzENuRd0Rvy
VbIAc3mV60dcVcX9jKGkuvJftp0jN4RiM0yFl33p5ogLoE7yGcvHXaNdht7fCzQg
Knf1a8BuxV1S875uekfeoCeMWRgQOV3SZjCHvkbOI4yTgyXk8KwLGwxN9HCz8psZ
U4U3YqGmighgxU7P51oHWKD7D3LR4Ai+d6/zvanFg70J33DIIdfz6cKRby+ulKsg
QU/UJNtF8Yz/gTKsq/hyH/aCkekNO4NfFjPedg5yVgljANl5YK4WRCgMC2xhoWya
6vZU/hZ0anlvsiLHOKjGDzwWXJaP8lGQ4oZUoUMhcYFWG98vgh5L805Iju5Bq4LJ
rHE+XaSCw5bZpiLu9AVX7TnA1B7o0h0Onlcyv8+Tx7GYfrcv/9hChbOVey8rNGEJ
V1sTW9zxPcNIQPCGdalpIuqpfTjPaW+3rBd4GCk7w7LcMtyD528XvtxKRLKG31Ic
DPs5zC8TUAiTu3x1UMs9bbfE7piK0YQqHZZa7Gmcjha/7d6gPo3mR2J+NBPsgr9H
Wp3sb9LwH9P6Rse7aGDrhjKvv/cNhEl6RYFEV4TCUsFrmLNLwNcRZiDLJ/l1gtVz
P5eqBqayfDal4x/zmulNv0BHw8/iJFfmaR4kvSMBpoiCIY1WSN01B2VCzMi6ZUKK
Mzb/zXMHsUL/aKsbEEnGxA26VhJ9QuHHkp80x/N6uxC3OGO7CvGCaMqJ8ftyzhYg
WnYkazTiiqL0H2BnqdHtaQYiG3JfPyOD017hnEsU6WWcpuo6TmM4n+nDWIeKk7Fj
t6LYWdiqEnIvNVS9cmqXmskLdFlhpUWV6zrt5RIbFurx/9JYLPYvh9dpfRvgo1k+
oyghgB2yqJkunvy0otY4zwL5BVaAWlQzJL8CwKXph0E6ShAuCo75kt5TtMjsaM4W
00orO4jydYaaOhvxs/5N7+1qg5b0K+gw45frTwvuQM/XjsfPBbrsOf+ZnC2PiMY7
vPzwlXiZrswSOcy/cgz7ZSaBC33Sw/E8HOnfezP79uw8Pk6+8tuQNKa187uLUCNV
MIJHfqSkjsfIAon1Kec2YeWIVgoxHagXCm3TPnSGyhYMvsJy/xlfDvjIGaOi1Y5t
SD3zd4+VIDn4r8LqAiJBsdxl1JdQ1x8ja7fSKnxPsCRki4MCK/4f1J54MUCaxIQ3
rusZw4Zjp1h659GJXqGjps0YOZdXtUcmOz5KrqgkZw1+hgfMoiq2mHIdjO0Hp7Ga
+RZIIR0kR+wLO7nlF0fFHOHNDzMSjxayr35Zm7UcrEOaIvlNtYx2o96vc39k7A7r
SEJDcXQUk2Y9RUFWQshSLvt4zqwZOzqJPoL2CIqpSJqbuuaWbfkbkTUO+QdrH3Ko
eb4wGRSqkVMG1Eyu9UU7pOIa8r7ML7yd3EOtEMgmMpMxlT1wKYxtpbGNBf23tqi5
P7Nukbv1PJJnTujSHF6r3NXuK+OEUWsr213EvL9VTqyEAfIQIdegTSHGoX15q5BE
TjpTtmXGMCTJIh7gDSKdtuy00tMdpb/Y90Ll7Gq5uXor3WBi9tORzwX6A8cHLQxa
imr80v3C8HreEReFDSYohusK5EX75/Ph589cQvKSOutaVFtjh3UEKd4OFk3HdPHG
7wzQFXqPplrcmNa5bPCmXEie0wCFMpSzzCWuarma61A1cAKQa8yUczztMaUJXClk
45HqsMdH5e5vrQs/tfQAfYg/Fp0G57PWPJRyRhxdZ7NI8539+rhOkI29m66rcGTJ
9tAYr8HO0sZYJ3B9oODP4DYvOqcKSdwtgl96c01VLrkiPlrrwqGFvc0MfXdGulTg
xGwXtIXezifxO0FrFRN7FL1RL3AU2a8D1YOZQ4o43lwSpf+Re5ivLF2xLXGVfhVu
2nPDUY2Jvpx32oQ63CHS4TSnn9PEzg3bYufcEl+cQqFBQGpIKAUJWotp06Klx5X6
rXE3nNhKOmBqv14jy5i0iW62dCI65IkdKjNBzFyGs8yeUNCduI/Uzoa8k8eGwCSj
vYfdbmT22Wr5KXFJhrtNtR+M5SeSu0OVTEiYP13fzfHSp26K8fNXtqJL6RRKVyhm
BFMuMkB9c4zNK/KrA6iIwhXM6GpYVuqpgLNo9cwtIIEmhZ7rLimYy7x4Cp58+tPz
l93Q4Vc7Up/3dMPoFNwk7qiLx6fxEJ0fUvPZmKvWO/KB646ebvEDRN2YwJwowwJl
JD5S30TC82BhIGl8QyDE0B4MGQOoiehkbnFdWW1eK2iybJO4nfzjK0lZy+v6ccwC
HApCUhlJCn0RCYwH2Wja8dF/xgKHz3liLeiNXQBLMQ6FVplqrWniL9NbhQxR7z3m
OgAN/GGaSS9obvrKb5bMHUokoBdh3EFbhJ8wvnikozABlCWYLEO2jfPdHUzcr1BU
E2AJ3HEG24N7NJ8NRKU6aFDbwMJuBpYWE0H+5mVnTOC0GchP42aozy8xhmZDaq+y
SZkvb0nPEOVbvN04NyKrm86VIReOc7L8Y4zaXBJrBV3gUbJvh4RTiBgaYiRxbrJV
87hAit28iPCetRnuX8I1ey+eR7ES9kiECoONcfKrtimbT+/lVShVQXr+pN9Xclwb
55zuFp1b3XDoOykbahi8Fn2PsknwUaY6gW7p3wXA31CzjQS2YFOGh5tExGo5gxLa
c29apdMFfmtPMqJpakCf+sP+Cbz7Z+GTr9VWuP5uKnA83AvlrasPjqwVvG5ku2Ow
KanTSqEConGkee7hqT1ppFAKAEGxwMuk/CF5wL42gwmpYCBmKN99Wd7jyeg8ml6H
JbewUs6zX2WAFjHD8ssj9VqAz6Y4feOQ3GrDqqL1qv/uW34NKdEiz2LUSWOEEvup
D/hruWz4M+ckulwrZUl9P3ilv0YqkkuwILqb5GEUJFlMcE0SDPCMOnmu5rrW9rZC
sTZbrH5EAgXDXobPdBKuihC4I3RZKnY9AEcZyLMp/DFnc6ebnf8UGn15Y58YswyO
OZMo84wX04SFMBqu8NXsVPFpljoD0A+czbDVofd9u+yDG6OxMFbRdkKZXsMmGMYR
hLqnzQA53q6ItjC9l8djx1Xk8jaYsQgBODKPk0CAJjDGvblBJYXCzbbBdyMT+27+
0zCyB+8UvFi7TUFvI5VULY6RDkwvR+zvNXXwZM4ibmxWzKSdi7j0GCqc5UmsVfyl
gpdJevqSW4bC55JHAiTnnwgbZStA9NHl1n7u42/ftEvrzhy78xmlHeZPFpGO/eWT
+p1Ur/GPKV4gT+qkNtJwM2Za91R5746E5KtMH2DTKKcGClPxY4fVq368YhJ16DbX
zR/l0Hjt4gIhgf8m9V44tOTtnZsWklzJ4B4ViGTpBKuqM/x8jS1peubQNDBMGi4G
VN5omTULtBmSnJWUJjbymgMc8PH3a28T+iOl0B1/3UddPQdUn5vFYD0t1AK8TL5c
BXA/7sJq2obU5oeS37jZ2/5sb6bmRMvfhxOrtQS4M9CF2KQtgHxwURobgP1IZws3
qoogJj2px6elpjNMXL7+0ggBOqunM2ea0qEoedywb8rTQJMqXI6DP5Vadx+ZleQP
I1x/TLljFzTD60SvWa3WNABVJLiwMT2iVevzP8l768X5h+uRQZiGSUldrnQAAhgO
vg0Wdgde51meMeqoWeF9uIXFG+TNw6HkyvcNVNG/gIYo7r+Yotye8e6LZlz6KL/Q
Yk2+tAkxgLOIhDjD0hVL0j65skN8tslazbY6aWy8FNDxAUJpozqGWfozS/vyMgEo
7FTKxNLhHBwUps5B8pwqQ2dZs9muftkvpCZ/A5IPK/6/EwxDoaxC6u5zyTVkEnum
g9OAEgi1yF/nr2hKrj/kki6joArNwLxv8uLrQpsEDVYrGPvjwu2cnRJoN8E4eNOl
vkZTVT5UgwBBkF6f/0UEhXWkGP76cLeE2fbP9x/FY987b4ZnTGY2xiw1wvFrzUw6
KwI26gEnRp2SEl0Uxqrc+ZRYJu0lmKU2F/adS9ZyFs9y/y/ZghocgLxfuqQRYkgQ
VtHtSIgPorgWkWW/5zHhmw85wPlzGlLbmXkefQRPgXA2/uTIwlQl5zltMcTWSotz
h3u5wXF+LwdU24HTnmhYKgL+/Zjq9qocqUqVbUFw1pFJXM/9o1j40j84yencm2TF
57jGryNxmjOv6a4+btZlrQz4PQaeCQITdj0RGvmbnxgXD7PriuLH4kzU1IJGxMAe
aNN9ytLuBOk7h3M2bHgECznkc51vMlshW4b1QJncFcT6AH1jgvVc2TA4Kc5wstVW
0O1K+16GQAHZJnhAdSVbebJZbiYxwY+qHwbZxuwfnsoqIMUdYBemvT4yW1PGAATJ
LkBjGuMMY/IJP9xhjMRPPrKBwh4wOk0chYZitn3BHwFbjMum+5uidtCUz9MVUVSR
flfREktxeA8igEWmwB9snRdd1XFKIQiY0gQOJUcekjrSZWcN70Ic3GR17dMRLRZO
9HCHhJeBZ31DEi+aKPKnudkzsGi4vNxEoOsc3Yrg+sUcne6TMuqSzd2HJ8IdQ4rl
QD2U1ixcF2bQDadID8JqXL5wibRdHz8rFQF+1M+6YRDAea9XAJbyPwBD0/LcCKRH
s9xp+5sUuX81+sQNrzsiD34yLrOhtG7rbyPtMHy5HHkUZSzhHWaFvuG6VpPY5H9y
KlWn3vosNEVqB1STXHSNUxJBbxDqieED2r1NOXAI1eAEt4TMTsZgUPVLslkVNEcM
q0tnrVBM4T+kyH8rPoH2qvziRCIeqIFNKarPoJLTRrhiX8C+oiNg9FEi4vh4JzfO
QkihPPgfX239PnV2/pS/LdbCUBbfQNXS7Cm2L42WpqUxg/braLrnSiizzYJn01RR
eM1ffbVPOckHe8oVJGby1ARqS4rX9wXoFtdglSXmFfHLKdcNpx7Ae+vEpIQyz8dl
QQfmjwlIay5AvThMPAc/zUE/Tka1cBpRQATZeCLb9RRaubQskUcS3raWSKVS1FNi
Qzxz87eP53jv73mEmSGyY41WZH2yMX1KKFaa1qQHskqS7cvTWmSsqZksbIHA8g/4
5UTrQNVPJPQ8d3hgZgW/2VYoh2+enkKWG/N2tTVz/26a3ukWnkm/rp7/E5m255++
Yk/zZgxQ9tCPoDgJMThu5KkCX0xcsDTheanPNUW//Esnf2rkYDkWxOcOTvUUn5uG
IUEKvpmZdtCI+2sxTDExJkg19yPD5jHr2Uf29JG/Yw9jwFuqrFYQjEzDE72KstWT
Cal8jNdh85BdnM1mT6O1oxOagg+/4UCG+E+CAxxAlHeqkEEqebjUQyLmD7B6+GDx
RZaS75V+F/fnyRDlr8+gfNaOYLmBsiLatMHJ0NJ9IUSKS3uLA4prhgFtatKF8u6M
ow2JAks2H2U5eNa6dV+ZEOfaoJ3mBp2lyzUNce3BQ4T9+4aWGLVasyIdGll2o3AM
Ycwp6YWKq+48Ny7GITeSgOsHqZzc7E4EYF4PodYKXQA8x/51bMw6ND6SB0yDbu7E
jftsGZSKjIGCBWoeo9KiYmTtA89EhYJJc7kLm287oOPxPC9GBnbZ/AdbKVOf6Lfz
S6fx0mjdktP9NKMnBFZtv7ttfWhhBrONT69aWxANYP1ArkG7A7xhR5iBqhL94Miz
nqPWfCQEz8yLoiu7vpqXq1ls0y85c0TW4rdlCGtnqJUmYd6eW7WHNYtX8X8Iwi9H
fZgQdSmcrGGgjKIbQUE+PFNj/khcj1BJwcwV2JyJZzb0DJiwM9CHb0QC0/di1FD5
b/vxUdtjZiDMFK1ctj8DW/CSnSFb0y5E/prBLV+xNZTaV3EyFLQv/t39+1RAOWHX
LED19ihXBN1quERlxwUYkaqBKTTggQ4c++tBbA8cWrrogOR1A9DNM6mja7Jr2lE1
btW61KlXMLN/WWZjge4juw0mSshj00b7gxx9K5eJDv76pkqYir5giFXDoKH9yl1+
Xe0RRR15TjNwPF4En7q1WpkpY5pDYIEFOJ0HUO0XHwMXSfgKdWemTeH15umEZF6L
fcryFh4fIAoRh3qKkYn5tnPZ6D5JMegGzk3IkcJtjVBkSJgyWUXGvMk/E/vxw/X5
5sD0dHuG5WupFKOaEynVY1m37HcGoE1BYiVIYZur/9UFAgl84ZE872+wBQi7FLj0
kiU7+m+rei8eAbLiLu2Xa8d+6nLL+PJh5/9+U869bALQ9gUn4vHetXruvGnUP0Ck
PoSO0HjRmTv0tzuTUJh02udXYRLlpgTTCRMa+nrIy9nkK3g4RmlTbxoU6MTb6aLL
28r5O3Vwtdh7lIbalIgI8cu9ocpOQnBL/YZMgZ6qSjAWvlmdO8K2TFuL7FdDzqx3
1fxoui8y4q3+ntcodYCAqz6t6oZfOWvNoCgCQu9CkQClaw7q3lDSMzSUlItY7iRp
yISOWLe6fqtVAF6V5RV6j8rj08mtbobymKwkMAkLZYoLOrU4bqo6TD91umm0NVlL
PsysEcvP0tlw2YWI82t10AP3Kwd04fOkm4IXUZUWj2kyflGiiT1Qxdcd1izuu0nK
QM9GxNuOcbYjXLZaCWYPle70PdNtJy5NzP+pZmrkA/nkKRb2TD8NQzex3m/qpN5L
ZCBita/G+Gkmf7nnHJ6SO2vS8h723KXPR19Dp5bcLJmXoLhfk4a3jV6BHsnJQuJz
vhzFh3qVf1BPM/tCYr+cgQ+SUWrGIxskesFWLhetfoBDWG6l1USaHlywf6hgMWM9
gkMJng3hNn/M3IaUZJmnxYpgUATOLdVhIH+FNUZ8x7M7M2mqNeoJAEYiTgc7eDsL
ygomyXqU8wLlhGjHi4TRtsVjovPdOBzlROoQB+EoEcF9Fb84NWvcygIsJMIXFADr
UQyXSd3gO5JXmurSo8LWEeszRbJpf5Ouz3UXwnRw64PpeB5Xtbxj2us46W9utjMQ
8E8etOahZBWzQ0+ib5pyT7JORA0wn6Yn7msUkIA3e6zHO5f5kiKMQq5pXd3WePQw
Vj0FbTVD3CH62ipUUKdDaDTZM3qTIEPickBbt/QvKc+s8FAwP5Fk9u8gRdOFa8+T
8YQuivTgED8O5JGi9HxnI+wIaXcAE7lYEV5uc3rHfa12O45CU1IG/K2BOIv9e0j5
IccgcP1KZLeIhUELkfrKCteO4kN/tl2V16wOX4oTqafAKP0+X1987MX7OHX3S2iJ
1/9Sx/SBpliMizPjZj4/do58TIEUn4B3R9Bpxe8CB5pxaRTi15npZFIsJsFMllWQ
8H7S4mmZJ2YZy9SI3si6IKU7MfdJtEjJf6tKa04UlSZuwwHXFGWWbrtYpxEUdQur
xkfswtLqRGfG9S7bvCziZPkyBgpIN78QJiuApqRnLzeaK5mqO/mU8ra/y9xPDu8J
36e0yrF75lABE6WrlW/ktiQEsiLk0vlHOJKeaXze5EuOr64Uu5AupiFNLiwaVe0p
lgrNRbSqCTQv5FWIV8zpihG98rfSeq59mmjZhxZGvR0Qks+Y6uHFuzE94/E22Xcb
JWdguj6B/uN9cXRlNfiRk9kyhJWjEWGRIPjMH+lo6b3am/Q5cMk73OSF0dIOZ1df
aGdk8Vy7l0sPNYqNkXcgvYd4VnqSuL3vsQyUjjPOymczS3cSpskSLHTaqJKaLzas
wMmEACJZ2tsJk6ob8J8Jwi5Yadw0igtZFRNQXtUDQwrwu7pZQrZvV9BTn+HIeXI5
Nr4j6vbvxNxDoDTCVLYSlDc0wjv+qMYGz/wJIaYz0auz50SXGaH5SoRdOmnDhM1h
jbC6K3xbH7iTgDYbf25JkmPXD20XdiVpnlYDgYYTBhkjfyapP7cwlKcTb5T1E5Pk
c+f3MO/z9zVFNa2X/5Vp4gve+xMVd6SJDMninKlfs6IRNIdUmxS25DsYa0ee8HPV
T7HUwvLeOk50A9DxbE3pdMgfGVJNf0eSBQ+LAfZzextkPr2cV4ftRJ3QL7eqT4Wq
sH6qPkR+LAhN3O0tFzOijziACsFAxvTybv3Y5w5kgjKPRUy1Zg+g7dsVUtM2rFlW
EggfA8n62VL0ei6+dGeKkDTfLYLjGjDqhvqvQBv52gHJ5TPjyFmLUN33cdTZ0+Mo
nzZf2capiNIaNFAmIh8/KmzpBUUg9Hyi5YEQLj1kwSaM6UVlVDwzOxOBG8NeTU5y
H4vnIaEevbArGeSKL9T2kY3F33Ctc9xZJQRpEY8I/COMsiapNybXbHdyHztL81Br
1wAdud6sxqn/FHW4GxeIVRCb7DLblgNYvqSj07n25MByi9YsXFm+1JPK4SbG9gXq
cDJSpoVu6R8ng9gMhzgseuGEWGbF3x6WN3WM/YAdgNMEN6Ts1vEJk9gAz23pL0Ii
c5TJ2KJ/kXTtXEvyxDwmYmno6d4Ohlg+iU0OyujdZZDAltzrXALZ4jibKG5nudNa
oTBPw2tPoAYpLjBTRO85D6ZnW+A9u7YwdLI+h8+fjAkzK1uXKNs33RXl0bJ4TpKr
ND5D1ZS8YwUR6aWmvi0tk8llC9+/gMeiDcFQs+kk+aDXf7ZT0A+4eMo9zMynQ1V3
zuIMFpOzJLeikQWmyDY9w7QKHEKwRqbPGIlPB+hNtvSj7n113mD77yyMt6WDnTyd
dKIsL4qFpy5keuizb8dM7nYYIcgbsKNE/21OrgOXYuGjj23jmR7onIm5auPytRy3
+49pLacl1qaPbZFTtwBivvecAdVbL2KARInyVsymQZ5m6Gc9vvkWcrGTwqk7T8JK
dPHiMbkFv26utXvAZGg2TC9R1i4/Wmtj/UQEvKsXNi9fodUrvlFmYjuObm8OdpGj
ian/faOfUTi1WHltPPE3Hubj7LBTnV2JJWqptLelYUTQ8l8AcuoJzYPuQRusQQIp
3GU98n398sjJyd6Rxjo+jsqHO/qYYkQjvnLFaDxMOr+Rtgo0nIBBSs3Wlfg3eTY3
nRBoFUqgEhWK4FNfng5mBQrNYr2LNGEId5eiLhYRh8L3V7BUFmAwstBLtkaz+RbC
tHq2bFB/DXkv+2GYN0oraruhF4FI8xYM9wp7DeQiQwxTwUhcxkYwiGrJtNtNArvt
hfqp2e5kisT21mlt4vFOaz5f2LB4zFKMC6QGOlbhkOvQLF9PYv0dboifiuqUOC1e
eT7Xx/UpBaNj+W6kBWslVi5d+M74lPTmI9RoFO3gxFQIZB8srtueYmgcFjMveSjP
xJY1Y1Zehv35VMHzo2v2VALuxM1uHUtb/8RY2LF+2OSg6P5+zaICmbFIdDAbaHL6
7b3ccYnLxISns+f0A6gm2hCMMJ0Y8EbKuYFQtT6EdmZJitsZ7VBW3r/ttxZyCwjm
wBi6N6l44hlGEdkuoWTgtJjqkwmjlT7Me3w1JCBsTdhZnMl1VKrYGsvd1iQLtSyt
D9r7EWGxyiQkWgajX2JdnT7O6wKwzQhiWxqGN9/hO2qNhosZw+u0zl5dVY8i4gWm
4t/cB/QSF3DOATaB5YgKB8HrFH86vUSlYwmVT2vwPxJe3GROeUElmrrCz5Jof1ME
qFuUNuS6YYY1YdjFUdN3gVTm7QHrIHjXzjTXYNyGRrOXgWHHQM7rSpzIXKyZflIw
lDL36vnA94XQS5M87OCNt8qcGUhLD59zi6eu/4yVkRkRahB0Lt4tTEoiGmrzp36i
KzSgsNqR5cLTqIiMBDkCDHfgZW4luoz8e5pgg20z1rc+lIuYDMy+KFAkRLdpaz2M
14Nj0xX+S5mPVRCHRNLgTb5g54ydohmVk/TkRnktECPnWO2nOZLBZmOrfYvuLdEQ
rXRwut7Gvx/JdmxwE6yu/gCjwN9Q+kgtVbrDy8ZqN/pwWC9KxpYCXhi5+jA7wsis
yLjR7+fj7ASeb75Ytp2XfsQnOwZbwsCC4aBBKqWNhWT672givyoJ6GVJc46bjJla
2FbrqeammrsU54en2xWWfe9djsPJ/pCLnp3Vhyh8qwMRta6w2GuRHEQVAKteR4Ni
Lotcx8tPQ97lqaKmxWtlTAU/ScxQzhMzhastv7TDzXf5/4q6Ry3PtoBCC6/6GhFh
6oBThMP2nTyeNJ8eTHCKtOU6fBN1pGIgHLcn8gx5oZqRhzPtdi5HqPud3c8wSmif
Vdpl4vUS72uzUMo6Z7nQPmBfvFxYEUbaXGp1wTD0ECj1buHkIa7EpNSL0dNRdu8+
RbzkxQwkXhkz3A/tQATVbjoB518sj8HrCmrHJYTF9JHpGDuEfVx2HrylniwElI+0
QeWBRSiJ5lJyQHGkchH3xrZFgleQYg8Lh7aZ2jdvcWIo4avTGUox2HmhbFBKnkhE
QOM7bWgQX26+EVTAjktz55F+sjJDW2QpBt49ES6DOkCuWFmEmFKyh5GlqsWMXSt/
/418zbO6sl72Zg0u7nSshD8YdQ4V10WZzaurgyXp6jHmNbkuaK+tNZFq8N2Pcr6w
tq8AojWwmpzqsdw2AF9GS145tWWXAv3BGRTi5PoXnU0zfg4TiteGqla7jAUfYv8F
6OvVFcN2rru7Y+TEDtBaZk4eMZC3YthlqvHTFz4hGEtHHK/dcqtIwvazLzxw49TS
8Z6R4sJ6ShWY1ynaZSvG0wqvG+PWqyAy8jI08NwuPV1CoAMvAVDx6sk70mLXKMew
hUFJKkhe/M6sHkIEcocR/UalSPW/wS+PtR5X6v9c5UGfCwQBnIB/iVpk4wdlqlF1
jMNhJCd1ep/7lxHl0OSojU/AhCQwfNN28ODO5Q2q76JuYPqc/LxSbD0ACG/Adwlh
2Bv07bxtZ0S+kDW7Vr7iCFCjLJbTkjZhZCA8HfaMCglfoxHYnK/HVlrxcez8Z/U5
k72wqyu4ONMPnWvNL4bwPFf41t1cbjwJ+juO3vVhOF3LOBvkd5b4B/mMqaYiANhJ
1wQj7WfxtXAiavaqVWVXdIspycXUg7PA5bgCHliqFnKdOkwE10eQjbZgze6wPpf1
fxYwjBxE/5ItnB8UBZrx4ojXMnNVOVw8QhGcXXAnWm3gGJayIuUHfTg5Tz02vIBh
CqH/pW6BafpzlWGu8kmS4QSISAHOkIVh9ogkIcKvol+BefcYNa2O7efiUawHtUgb
iGtZRD3UPwuhsGy7s1aWLmyoHR16HL++9nvkrs2ZAGSNk/VXz78jQ7rbLGBjsXNR
iBO3Oab8naZvnoXyK+om5l5TA7S0U8Rt4E10rtBStUGa51WECJev+fFVI3j/VR5E
POGyUnaWafKaRizTiMcSoLv+9ctXBUxJ6YT3x2T4x0jGpjYhTH/yoREGgwA1NWKY
TswjVBQAYSzOUAZpGNX/wrxzzpQGQQXSr4g3RUG70as5WiaBeKwtViA5G4JXIjgn
gGbQF1rdBvE1qtKmndbrMAsNPhhdbVNUJMuo3+kRbeyya6POe8S+v/NO/3R7MNnt
iuvs3X1KuNH+D1q1nu2oG0Kh9oaG0UjcyRIUOLPegCOJoBlByfCdM3Ti2HGy1/e5
6zjc+grdBupojgj2mABC9ckxTCVa7lxKgvfzfneYxUVfjJkZ5vEOFD60xmPmcqDT
ahuEYQwzRRNt0riEkifMSq5sahZ+oejrYm5cefZg8S/+7aue4fQc/uKnKtzKoMoA
NZRjQQiCFDHTG+1bPoTO8Cmb6y1MuHIxwRUeawO0RLjnjeBf1194gsg2J13N6Gdl
4Sz9bokNp5OLg0KpqfzfoVaP6XfA3z8+G8bxRGGHaa1bYQ6Krq0mNt6PHCOr68Dc
7nvcAJvZ2VFldzdT4ZTZVqXLHvfN6FyFGiGbhH+HNbsOk0+n78xFHBf06pW34DwL
+QwwtU/TjEMcGyI+ageAoWRigW/UN2WzmLb7PE6FEMK+38+xazt5JtCuQRVwNV/V
J9R+LCyRQGSzN3FDd2GQkkPgcnqWF3p/n86f95j7UPIwtFEHc35bEVITIkoIFuGJ
K3BR95bNIIj99i0b6SRk4bYDke5fz1RkY3bm/xWQKnF0dLsLP0r+aPD2wd2yI69+
3DNV2KHfm6/1Nb4AR4Drh7nQWzilMQQgkgE6+bWBt8mmc2Zo0ZPg6SnM8Mk4UKYQ
RjICR1PQeukI3JAcG9BqFhVUPYh77ZoNDX1o4LyWn96be6WCYzH+XreWu5IwXZeS
hEirEyok7RrGYDZZzu1xIdsdfwLTXnSjlmDTjzaqQPzEeEvvbfj8i42dOls5ntvw
SKugWXDxVocjd3DorVqcRfzXOVmomK+lTtaaPhLjettStWZNZ6EIk9qLBs+hgZqj
8F7xAGJi96cKObYgPtkqXNgUQ+hgBm9eiOvlErSPylAtRvlwpynJtDLVF996yEBG
VUM5uF7GA4cbkIidSXMFtT2VeABk8vnhnEym+1PfyBkavHmvRMMzzJJZC49M3zOU
LcJ3k/XICqc4KvQboxyFqm1o5rProVI0PiLYjP8/Td2sQqudQxULVUQw7ZfxQm1r
uTWB4wg5kQz8JE4TLDGkzkOidPjILnqP4xUIuaiMaYg9UJvSgyZ6P9K+2CoZTAWQ
LcGJ9k1YfhSdubbixYdxn5OZ5bmLNkdWMtadIhMHbNdzml4Sehr4v7qZlFzMDdQZ
TLNiugTx+CdUc9Maq1GxNyf5OLQ3rwqvMvnRuoEKk3TXXdvpQqbAj6xhNycHSQJg
qKwdZAwU/WHtNGJnx6j48FbpimOhAdiY88vlf08J1MGRX/zy2yEqjtDQiW+WQeMm
PzpKsKIzFI5sx6hQecYEIExmBvaiSBTpsrFSII/a3O3ldlfwFk+8NRmCIbX2ORwZ
PqcEl2yuurfP6eIQQq3mqGVBjQk1neR7yeeIbtJ0VDrsAPRf02dFFmUvlUU4Fv3T
tHkfHWddltg+UDhABld5oSWjwIw2r0rXdZv0wCBlBlLr8UbnR1xFJ2PhvFHHFGE+
AqSHUcVg9hwfzngJKRVMkeanRMVc/CrpXTjGSKiFuWsDqr6gG6oyQUClztO2C6pC
d8qtjaR9E4AB7lOiBaUGDR/sQpabfqCdj0+/CcWlLIO0/JKZZeEcTfLaes8K2+3+
WdbO44RuVAvhsZ0jMpJYroZCMhLj2xhv4jb+hp97AVYWWGM+HSjP7PD5eCSVivx1
XsADIlbfQJ7++WGBb9DABuL9/Q/Np8LT8esF3GAh0CeNUq89lbI2abMuX2DRqLmh
flFB3xubMNBEd4KmWgnNaqlAwmMC9usBDKlL/odRDgtmH0qTIYAJFX9nqzCYrgsZ
bMkDKU92kWuY68/+glXGWrhR/8nAwLQA0YOHIOIb9oNri2gZhCq9Ln2cQ2N5a+KI
sQn2s6yVIwUwuRwAaZxcl2PpK3KkyGTSExyWHhr3JynjFZYCYMJNJv6itEt3EBiS
bxlIjEMRPUrQkC/1bVVM0YUwiU5iLv59V8hcLgjAbXAL2j5NAk+mPhvmr1KCqHOG
uLDNdl2N+VBa4fseuOUwVQb7q+VQnDZXG4nTqHaos3IQNXDwCy9KZW2v+zDfuEgp
G9x/QJTWmcO/ehFo2BmT34cUhRFHjJ+WjyCZHy8VFB1JZSLgkGzYbispKdy9I9Ek
bxgTiFG2Cjd8N83akX3aXihHEoAelBAdCGUFhpf7E35AkPHFS0/T+yL8vCApDCE4
W7HcDLDtlwsYhdLWGlv3xWzutTZLS7Uzn9UphYmI6eklnU296qPRCul0A/UuBwdz
Sbvbc6q3yFUrRtIdsT8SuNCF7m28s8yKkNh5EZ1/tEmKbCHe8ODO/3b7LEERg+qz
iITdFB38C+S5RWv2lO3dfQIc5ZFcAtbTJbIX8RTc06ridAOCfayl8c89/QSRaYJC
VojjKtWbrvGS4jDSdHLLtsMiX3Sbthe6HrvlsaDi3OsGUY3JPZRXMO/bqDxFQL4J
DviFyw1NYwRaPZBrwioBnonHKF8irPYMO/nXyaK9ZqdLxC1yGjGlZ/uj513EQ6dy
W3bswMChaj8XXSYspgniZWnOXzE2BcIfskjGpqXog9PZqDyf3cUhjpktwpRp7Hb6
FHABulufD4ElN3GtEXXjXyI7dbwRpZJWqmRqrny53rpuIggfRcliuagw+6FiK3Oe
ZLz3JOg1/vhkpeN98McGudJuSR4tTdf3f8wGMkNzJNTwp+lyxzZUJdJAFx/TCi+M
7/hnsrweKsJ4pD8Johjocz9f9UpvXm3SpTVF333ugBeXuZ3v8sDtHrxDMg5wtXan
wbG/XI1gZFw+Fz5APaZ24Q5o7OFRAIru9JE4TEmXW9wCqAG4Ni77ywZ3vunB32hD
XDNJzAMGo/Q7K0cSHf7Asd+bomGj3e7StW6d5DpCxnh1RFIr2AyCSIJBSZiTaPLS
CwH0EkZXc4tFSlZWue4oFL+gb7iEOBM9/UfK1N+I+4mTAz7qzOREBe5ncg3RjTST
FzvyiOYHVu5R9XF1NlNcyszHcAjAJEd7RmMBmzNhskEbBbllWKwyh4uKNbAvvfOs
Bj4wZD1skmwpmNoCL+k2JZ+YfJwnHfqQ/6HU8iWRzzAfd/T7kSBd6nKY54jypXfE
wDmkY8k1lFSehyGlajQBYxTOCDiQ9q3y8dRASdrdXeGYYttqNM+2V2ANBE4pqisA
bmWGd7aVyFey8fUa8dQTMu1DlpKXQdFFuETkHeGYEexknDp3F5y5Kw+Cf29pbJ1K
8iP4m/bzP1WfKzXYOB6a+VKk6Hg30AHiyDqRpw7lcMNE1ZbTN8Zw533giiaSKuHG
8hZs2QmCGNZb3+Fuu4zyGeOVKGS5UD9BRB8wQxSNG1gu0FazfTobS7o5RBHV1WOX
hc424n1xRzXH5GjZYRYnNRtcpZVi2pVqvO+aJJeq8USDUGr3RQMCipRb7GLpKcDu
3fw7ha1hEIEB/wx7khHOtys4kjixQTzd8jnakbnffKaZlXsIaSuiFDNyiMhA9LDz
J7k39ZmihO7njCiN4o4KB2GztEQRarzjQLNNzHaxIN9tS+W3nX4zuVCLGqAUiA5Z
gDnWjMfgxFDQ1dTaD7BcJNh4ya6y43S99y88KOLJ2JLC5HwR8Gmj8pJNjl9E4GlP
V6EVmPiY8nmNrhn8N25IX8V3/kMEv+3R+gJ9DUqUBTss9P8fHNduQyysBhRU6T4z
xn1BzwWmipPa0wGaveT+5LFI2e3GbPuvUbNXiUfN0vVhEievIWVylaaw9+GZoCsS
3CJ/beMAGAAGov8KK2F9JgJ7vZ5xEqm1pBXjK4vcbBU1Lb+fZHJIMEAyWl2afRpF
LNb0eKbrRV5W+baQ1O/VqNI5mjyiyZUHftdPo7c8SWIcmYD879WNgnKaeoq3VXys
Yg50eJWh9viHF+cUPWMBoBb0S2ScvCEX8jmAN2W868AwKCH7igOb6MlX+qpYriKS
g9x1iuhD8HS2VOHYKeNeNCZMTVsW/vFm8HASKLJmv7dHhwZMQQXuDAxDTQeWzZS2
CZMHLYGAgJb/x/VIpDwLWGHaYuJ0CmOU36njyUJVVy6jVsbcu9CZZwJg8kl4zr+9
u6Xncv5TMgh/dvoEDgiLJqfxQct/UnGBvZ6CNhGAWOxC6QXk86z7EKalNwN9C1Hr
NYQRc3NdvYSVdOqSGH7Kbcf6TChLbmtRCDE+c2CKIU/ZdlfgjANCqaP7144BjWdu
j26kjBPl2btTzMJGqy3dmUDi9ISb5Y8Am6ECIXbPPSiH6MxmQB3HnR9E5DpYSR8o
tI9e+8b0A0dyrUjfY8Cd2vp0QBwUQwfvV0hb/l+2Ad8ph9adz4070Xga3rjMmlDX
m4OznxL7eDOOCeokR05nkzf4tLeWrt6IGDBxSJRhQ8SkidROBqzBzSGDTg3lkFRp
ByIqp5V1s1sQT0BkVhUNfSw8kz68OZUIKkeOwv+qHREg1RV+ZcGWkonzHNGBhlgg
cEeS8qzhFaeAjP9PS8N3sppHlgbSlv7znEVBGFg1BqxUQCgbwi5YQ76xBTA8oRmI
J9BY+FJLrW/9D6v/YB7mR5Z9yDyaFhedDQPlDu1RWLFFziRgKPOdng3PLybR3fWr
smZNDPMy2mk1oNvTLX2E/luGtDc3kBgukPi/caATdWg8mx2EDxYiwrsm1iJ6xFsz
OYuSAav3sGEW+XEDDZmWG6mye/ZLUxvHKwe2Oti7z5IW4Me995coy3Q5KmpzN0TD
1L1xAxU4M6DkSori179OB/ORBxzDnLVapJgcNC0Rco+osPXt4rPRNTZnCa3WpYk3
XhE25p0swITZhie/JdJdVAtByBbK3FBQTZ+yn34d5E1B8GL1wiLWfPJweCuyU4q2
D1RZ0d0ZKorLNVLygrq/XZE7NBB8Mnb8elgWXpbvswtLuiwk6+SavQm7TMkV5Ckd
/0jOgWj81Zp9QKLJWLi7PAbEvUj7fbPDx9TbGXmN3qsWlPtrb4j0pxsH8sOoqEs8
brN61w6Uog6Z87u7rPhWTHIoHlpLiMq3BYUGYjhOPJZR58DzKjHfIQz5yKaCffyz
rttV+VpwkRmGJOtcdzVypZhVSxpDCmDC2xK/7YmD4I+wUtbMXrNSYPAm006OujfQ
FpVY3A7h88psCmXOT4mngOaSRAQnQAfRZypHDqjBSWOUpC0q8o5ZcZ9iZUlIRS1a
yMBabevUJWXyl7qBC4jK7BFbfJ12x4jIl5TjQbkIX9kqgX7NwhwvZuF86AtxRZ8E
pDsjwP/kwTN6BEZRJ5+XrLcWn37MfKe626ljuIHe7nHxMfpLPwxaTeFDgNtmxQ5T
uluSsnLKmqksEWMTOXQbfAk/ruNq8hSqlzCk1Ou/m/ia3RN8lqSFjWOkAXF8TDRE
ScftMbcoiYhpeKvEoEbRGu5nA1gcS3VRxfwVBHgNhNdHwNysc7fBbsAuf0SS8gNH
ORWXL+40A+iWwuGvM/QFUgPmOnfN8RozK5NiLsofZ6JpXkGRMJ4karb7522JHJZx
WdkXDn+3JFNUO2ba6A2p4SQe17Wbgf6Xdh4Qvx8l40cSZsyp8Htu1QKvUhDyumEY
3he+OrfA0i3W+5Z+gkK7arxNtq9yzlOww553kjh14CZ2HpPqgsLorUEF22EtYi9T
UZiaF4T01jVK4Kel/22eyHtbtyE3Hg1xSExgh99M6xVqhtVzy1d4YKdsgMLLPD4m
WgNPTr6zQyOEfCQHKTxR8NGsXDPQ7b5oHZjgxs/gurqp2wB7rnpqXiO6aqtM0lBr
zFP5pJuzbgmg6B01mgjsuPipSyVs9j5lvdfPQySfB8e5NRIzlGT8nMIVvzOfpRWe
o8nZzKaqZMzDYtlslJYVxgkI1S9UL33noV4TnhZxhWnxiWAeIM3V5QGrnf6Uoxf1
UVYTdKS9xNscIBaV1Aa6L4mE/gTt+Y48z7oMeWyraads4AH9Dv2bLK/mV2Ho2YX8
YH4zQUUNZNnP6EzeHcKuC2KvjU8ORXruRTICNqfCpooxNoq5l134aYHumrBQ7cgm
pxhxUwYCKiCrVqXEpmURnKUn9ISCv8jxwZDiCIhcTsm50GM7cM+SZoo8kRHra1Ao
sH+TpuSKLfeKqv0CcBtqlzENEnSa4K5rxDyOy9nABCnXwTKzpLZB891JRgqKeLp6
FB5lfdeQdJv+AOAHbN/tMr/QqK3blikyxauhOcHKOpi2002XKRjaCcvAm5zKfj1m
A/v+lS4bSy7yUfVeLwlTbItJOEC+5SGkC00SGY6I9I0fCeXMqFzhPPldZzTfTDgN
8+ajqsL0fJLRZ+OIl3lzSei7SxXMTsxDtFSbuwZrokjAXsoT0K042FfOxFxc7G7K
Ellz/OMWg8iy958cntVP+IsHMZB0GO00e65OxamhMYkFOky3Y9cw1yGCMutcYhtv
SFW8UYf6EeJ8j42vXtv+VGuNQUlAm2i2ORrHqDxF/NEYrfbq4JMWu84OGbtc4nU8
4xIBhhbUeDeaaIe9ZU9vWoJ8qovcGGC9yADoIKO1HixHFvmAasrcxm+GjDHj8K+K
S8ztXevPBAkrsz7h7RZZ6Gc2A+bNv4gH4wVeq9B2ixb6bTOg1mN/WwI+t4GY5nbI
fu9VtOwgOksParCEefZ2NLFzgnUJv+iLwLWs93t+ptKKC1Usbfea3ubGqYk0nLdX
7rpj4VlBexJtSX8QgVw3bRSQRN6r/U6KlCrBa6Vm6wnS9L6gwqknc5JlvqDbe7Z9
Li2q3jB3BWhLQY0INFfH9WA4tHH9ANGhr6HuXF7CKhTGs0xg8O5z3CFI1KMtRy6+
ZYF4InY8+4sIKu9mpTLovLM6x+a73P/j/udglIAp8HCgNu2ZgvLBcU4+tKc/+UT0
kHdLGMvXz4wf3IgOg8NEAgVdKIfwsuQjFv0AEioAC0y16VcS8/NMihvp7ku8OsUt
FfMRooYlNznjU4OgRAeLHDW8Q1+gCohKXnt6ewHX5GW1HPvDftXvyX/l7CjJdbI/
ObIslH/YqETZzX1GiANrTqtN7BWJnjOsd6Wg0IAjk4hPBi7x2wungE5z7fSp7MPN
3BDQxiKj36r5VdxEAHbeu3JAH88N6HtNLYBovG1Xux63V4LmgZULr3es2kowA1tS
XbBS2xFQzvxu4fnWpP14kVG1n+PSZSA78ZmWTL8ycNcWkxs0rDmNdPnrFL/1VQN8
8vboqwkb3eeUUYqnedX0itC2fMj7kcN1EMvZ90dGOBX/L476GGXuIBhzPLPt7U2o
K51kqRpDCIfyDI0WrqXCtFbEr9WHMEPFWqf9w2SNYdXeC9U0LRTJ4I9wIEtDl6Q9
4ylFdKl2N342JokBq0d/OfNmGxakvSTyI4QsTJDWQQnrzkwu+r69eXrboPfyLgK+
sJlJhgC83fhk7wyX3tmuTR+4eAxMuH577C02rrbE+wM3B8XU824NEjr8odDqQrj9
i1quazQ/C7tEYDLE4I8xVGiFTVm+Gr/nBsR72rdCTzNLPRDpGTY6cnG8mHv9C+Fy
SXoJueytaCBfMnFT0yqTIVW7vwgE0CGMUC/ssobMsWwCHvlcJ15wdw7NJ3D/ijXl
EQc8KSd0eZLYQbhm94acxh0i9NQHWkddhFuuRMV+7ETNBz+PNh+MsR5a4klBAmXc
10tbIsjdchEuF+mSJeRfUOIoOAM609/S5DOBuTbzPaXQ87WbhfKokWIu4XeR2R+i
/czFJXga8X+24keze7t+OXkP5O/IvswZh0ZT+0l02CPBFY9mkyn3d7CQ99EiKsSi
ahydQ7/+rAwZrbzdxUdkNfqur3M2p4Uebr+fVWPO8UTsH9OL01cWRaSEO9hclGGS
SIbWCN10Y/Y0Rfmxl183XM7GKgeMtbF2eqXincbJLJMmmidcs12lFEsO4rDHPCV9
/HUkJpGXuj9V/WHU2GxEpnzbcrxtWjjtnxD9WOJq4q5zFDHThrbVQrWpl4yk8ru6
rdD74zqTQH1BTYZniOGf421wERRCcJuV2GEQEuELyzhe9PGZLAPY9ZdV8ZJhUQLo
dlR1yv2hTRQWTulHRepEJIFbF2kwjmaAT5qJuPEJ+fgb6LZrzwb7awHlEv+VU5nM
/5IpjrXVpn7Lfn8Tua6/zo5hhzLNhGVA/bVtpvyS4h6j4tdo1yYxPCKKc8Qjnsq6
2TpXsloBaI1I7NlCDLb2iLQosn0s3IigxP49GqR1UT8kan1RXaAgG5TiDf0RS115
yjjj6FDSnllr0iMpgUsLrxHj7jJXHkxuUxW0nK07BwvO7DDTZ0DrK8XxENb/Bl2f
BkbNSJoHS4SBEqg63qTq0W/cp3BEcIvDyGmPetSdlt2UUOCTHxx4jL4bQ5eNyx1P
HezeAb9bqZg4xmgzL+aqQLlOW9/KCN5V56vpk+1+fvbSeZCeypwQhjkzRdcwVZsS
eL6n6GNCCyFSXXATSfGO7Z4yzDKj4/Cf4O0BT0BBl4LpXqNTg15l1gbSbTJFFFmX
1tvl7wVRyoaAX0fv+t3nwo6+XB2Dye00tEUEGcCPgeo3mPDDFzBY9jJYCMx87R2P
0bZbUdwXpjLjouENDdfzqnneXbC9fDbNpeMvHjd4ti30vhwfHz5P4sM3shPmNxQD
LC93rMF84AnNkWJWO6F8vStXrWcALE6NyzlYx3wYWWUKokNXZwaEucgq9+qm5Qwn
jL+VdskWkhrap3IbnDcf8wlecZrluAaCL0CkN/3jcJvRPKeaEnwSQD1Xm955L0qY
ybSwO7sgoVSS/HhmZU3ZuaxUul7eeY11Q8RVHkFthgMOq5mErGV8O10dW4B1dqha
T9aw8xmIaOGKKqtlJwgg+rucTTng3SjZV5acXuWgukEBP8EKZxnyTJiF+cChgd9e
xkfbQ/agshWpayeSW9K7LW5cOrxRIciIUzwalYiY+YyfatECXzoG/0ghSoPvHIEj
T5ZJDJPAPWOzxrnXNrXHg0ir6fkhuqCJ8IhT7rv6+DGndk/QA67GZPSJ1+al9MTF
r//J2f4c87EJ/YJ6Jry6kYkAINcD7Jy8vEpiCKXa/17oxifP94paqtrQr+ob1ENW
pneGzkxi4tUvD8zxloOJlkMMYZf68NdtXavesOz+d3VbS8wl9f+MIeTbsXFUJP+5
2VSg6MnOSCxBcTsvfIfRCV/+hdyZkVX+9uK+FGlCb6UcAL7ZpJv3/dr3hbuSe51A
ck6auBjGVae+ammoIpEnPKPWjamM6Gy27Lx/xQsOexoZ+7aVbb7ruNEr8CTbzQbs
emmvDg+TIN7GUMYvS+5BGvfSV6Iak3SZCClOqVBHR3EK7AT+lm60rw/bUZlgSgR0
YPoWriBKRGNJ7/Wiv5m91ILJ/zsUFcZ83tDNjNBkvnGR/M5dA1EKQaQqn2NUxMJy
DHtb/6lZehOWRDo5rlLa2U3TIebQUMSxqqyUnqhBlQAf/nCSIQhHt4vWHk/9f6wn
HpLQrL9Ke1m2yRnFnAvEalAOwBzuiGCgkaAWTLPqLj6bS+CJ3yKgqRMo6kGfse+l
0CTuE2ie2lDTvKBgu6HpGm2ObDxJelx1OMW034cPUXS2jTMIndQ8hX/IpL6gaiNQ
se9zI9AqsEZEjWSvbhkj8W01+GpaRcIqWihu4c9WUCPLwRsvymC4dJ/Pgjthn2d8
QJCs40bMJ+TwJKGPj0U1Zcs9m8e/dvwbvjAlGxdqlGXKIn7ZeY1iX9vGr7l+vGNy
yLFcNBoX26sK87eKDVCYNEAyq+UeDZVw3YvN5HiOLx+aknHKcHas4U/o/Lj1fFUM
pSQB8sEUXY/MoLyHgXWMK7ExYO8Vd/c6VhsRClPv2THOIgBdnDDzZkxC9x3I/mTl
WNUEzlRsoz5ODfb7GoVuz458E7Uu6JRkZ0tU4V4icSn5FexqKJ19UBcRirQVCUGT
R9BWQ2VNnLty3TZzhLk+nMZx8cCA9zyPxMDqFfRp+yrMHFXQgQAvOhiJg63qsedi
RTDH19HsyD4+HO1XOdDI/uYoMPH1yuopKqfRzrRKsbhBVJru2dFz+0DhVe5NgETZ
dskEHKXek4X6/icFfa/j3e5mhlHYNeBY/7P2pPQtX3daZaO4QV4oAMTXou0I+wxn
oQneBx4v6sqwPmAlT5WQYVDxnqSf2IEFrw2q0UVCm99syWyt6hFaEAW5ks/C6f4F
If7KGi1fPJV4nKqLIxhw1YCzWFj+ZVTt5gVm9DAM+qYYXUexU0TmB1721sasVIC+
/znCvDwkDSQfbiA90IyR1kGWUGLueS+mj863G4tT75UBV0rLEkZXyk5q6+z9a+es
GXYbj92iXONZ0Bw0ro51d9UHtqthrRXicFpRby+ib/1ac0i4iqQUfdUQq6byZInV
vd7iJmVtnG9azRUHPrrMglpoKHGcLgHS/8VbRaUe2FVNNPsWRNE8KVRmFho36VLW
SUyrA7y4KNCNQi153p3NWYT4jEH5wIAFmnxQAKj4taIcq15T2/NKsPheLcECpGLv
tOUlZEwwurLz4UziIBr7+ZMjQDMXVL+xNV7OyqcF2TTNHXnHWFN8mJ2UcTmSXQvd
q1LsDAeZ7gHFxCuDfFHbLp0mg5rsLr9gI1MW7hkgKQbKOXC44/GdE3L9zJADYXR8
vLLaPUFZNGHXMO/0Hk55+9JS60aqLJJ3hVeTFZv455Qjc1A5K2AFtnRwgFTLVKa+
2f1Q+0z39hK0XZW9x+qQQo04QalJkm//RBoG3qz7mbDr+nyC4Peo1G5lcn4+XRT4
`protect END_PROTECTED
