`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4zMjgmrGGK8ixiYhS/WRZGplFzvLFZMdwOP31xhB+vBf7dILlI/uty7/PkQtwgYn
r5pALfg6ocAco5DM/D5EmIyomdFZzH+cBh2n4zWHdljpMQC7h40wMxuL68OSf1qd
xULFwxijuo2iM3MFMUHS1QaR5aGb3MwLEai+HgUZBJ4VhutHL21b/jqoTD/94nfZ
Jwfp/y6NItMBLbx/yH5rT3MNbfhloDK4Cg+FCtjB/BYov7UxzXNIb24rjGUCgaCz
`protect END_PROTECTED
