`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
hjxppg/aHW+jI6qJj2mBAgF7rz842uzUPhMGcEbel1kCV7i2rpgtCM5MM5J4tVUf
C2+yt/hAyetxSB4gkrppqZqb6TB6Pv8CWuVj+ZmmO9GEyJycaYbwqRoyyCMTHjq/
CdgujSwfGbj3nhTbj9Smxi7bG7QyUwwSfFqg1pFcSn7uGaNY3dxlMKc5E9y6ryko
AOoFZlmoiU0Tg15RPr+e2OkwRmHlaqRchKU0Yth/+pYRGydA0FOV3Dbh26nztDuy
bTZEf/KlJQ2D7ihRhJOVvaDgok6/8AD+3RJpywiP8Ec0M8LSOcCfiLHPZAVN3OpG
KVefFk/5xYKhb5TnqgDQ4n/Ete0DMVp4foY7n5P1VJ7Iqf0+jTvAWw00yNt8FkGb
qS8LNjng2mjENlXbk7DTQ3tnrvjsEMYjEK7gTAZsj7Jt132GDQoW/vv9LADsNpet
7vONJEerKPQJHZPy86tj/IDleoEqnhONp4UP86QL18ElmwGnux+jR8IwFBO/A6Xd
63A7OxoI5/g56lp9GCrlvBxDlpytyowVEdTNzGjdTnR3ltHQ0KNgb6ey4lGG/1s5
7FgixfIizN7Xy7NUarn99HQ59XcvyB3fwga6Dw/vhw6HiJshN4JfO2iQImVXtnls
VacYA1w3BSxmybcSMPHnmYShGUtvN665Rcj6q4D5Rnb5w/uPl0wavXUBE+adRbd1
xuZeODXF19RHHwz1tSpvNqMObv4fegiopJgjCGEr3bmNGoKc//di/VvDmZp0TdL4
m/6W2kuNJ7sjW03eBVl2/9/iUVQEIuyWgrwaTx4wnCtAmmMbTw5M/s1RVv0wAwPw
d8WQx8EmoODLRyvB4ptflTenzCplYViPQUgJ9MLp3gnLcqHNbXa++60A+39y7sIw
5XSLmSHbuh+wLMqC3+W/qURm+a5m5Pxt4PyCcTPmn2/E/blgDmjis+Ep4DnPr1CL
6jzZXpH6qvUTXEm3RLPZYVGa2tav3jkN42vO3g1BmvGMTbP1qgmlSYSTPGtbepRm
8k2eORzgB7Z5hauoyTzMBQ==
`protect END_PROTECTED
