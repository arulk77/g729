`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEfqAwspuNbf4cf2SoSRseolKrYSVlb7u+6nIYZoMBDv
T0jEk/EyfNwuFP4ZruGgpE+U75LS3JJyerJBNDWKg7DujU1zHu6MkG6p2WNTtXnx
mAYKB0Vepu+mKJVHXZqrzg4tbD2jNV+ql9wK9K/RQiWPMzqMsUmd5NCD5Za2el6H
5YQYxgIwzezwRSOP0JlHOBbCrodu8un/TTfmJzoum/rCv6LsJCEJbmJM6hZzjeez
mV0AYEzyYwKSPc8PO0dVS+/0sTSSbXCCjo+/VoxMLVdZIEGXiWpDnKWXxrDvC9Iy
o6HEVBObD1Sy+SVTNnixfOu12IQIl06HKwlGpYQ3M2gzZr2ByWvpbGoJnO2Y4/8j
UOV5phLasOVKjx5mYy/SDcUoA2ieMoEVVQOOU6lMohO3v83YUZJ4tUg8TlDPgn8t
eSneGfDGpUYyQywNEwxODogU5WeuFb/OkFCR+YvbicahUJeQ2AXycnQ3olPh6Hwi
wRuF5FMOFM5nakvqYaUEbKlD3T8iq3UR0bv2XZmiY1pjPZvQslla9ehNaocehiMa
U92hzvmt6Zxh5Me1CpU0FW34Uz5oM1R9AZ3bISSvdtUYjU0LIKCkXtqIRLO8cXlX
`protect END_PROTECTED
