`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Q4NFXO7uVTAhDxfX4uwHINee1+K+u82lJkcqhhRqNr14FZCh/tl4a9vR4NMvJBCN
1ys2DaSHHOFCG3NIm5w6bQ8dtpeF58qRlRzVkI0dTP1l/Z7Wwz3QxphrMPOM391n
t5IXxtVtqx03OiRTabV6m0PlOasu2qp53sWo6DPL8zYqWrwY6mWvn5C+5GFpn9YK
f/UxX7NQCL8HZom1ObBwzU4neEWXW4ZTJ/5S1T3FIehJj5gKL8BTd2Y2F8NJBKJH
DIcEo4SOIcGcBcWSlba2Nr1zprO+e/eIRIdt0ADHMBnuPQr6jh9X5qfxCQedVhRg
8X/GW/EUoo8CJWMQS4ZS+qjznOZRNOV8wrla8b2d68k=
`protect END_PROTECTED
