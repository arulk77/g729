`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SVE6AYfWBQ0WglgGc0KHX8U7fLARhujjWdJPHUoOEXcT
EG26GNnxDU8/4UFgB91Wp8CPd7ORAUSRIA1xFkWrctH145PxxyMKWOLRVF3ojyxC
3LM45FVvA6+fvsMy+m8GV0sTzP0sZGw81vUGwjmpET7sdLcPTU52Wy/IryQSXERB
JvfCBG5U7K0qL8oMubtFtgPho9vc5dyR8HPYcnD+E0itP2yu5JejF7AG8Ze0nvjQ
hyNUoNyZa4LxshcOg6KlJdpfggl/qlP21PGPh38jltROLjFnIn3Um+fQ4H5DCRG0
YYLZczttFtEpCOznoO1BFg==
`protect END_PROTECTED
