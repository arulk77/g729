`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
CcrdRE4Rw7OZZghkNCbrEVMkOpOuBFBOGyCRmvARqIzL1hBFeAaz/755ZYM+GGe9
wFI0q2pTReRbZEeAX++8WaKgsc/wVO6x88/j9t6I7DBm41fIEb7GGhI0MEjPyGbd
vjU27KmTYJ0g9HyBHFlphgqjYM/JY/JmaQqv11w6877u1P5jlUxrqmWYORdki7Hr
`protect END_PROTECTED
