`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ0QAkBdWh/bKRpYGK7xOZkRT2BefOgBTHib6jE+OWyM
PifyNrh0RL6Jn+ywYqq4jCWW387OH89y26N3pNB1S9IAuusO6J+9/m+TDTr89rW+
w/WOBicUPGlx15hv0lIBoK18p12sjfADaDA2/aYykSA9r5TgiVneU/Yl9DKTRz15
SM8zWjQI4zhWfReLvDW7SdTu1Csgx8PCl0fzmyJt6MW8e/YoBMz/ETHxjfCuzxlA
c8Gh7coWypPgczZWp/0eFxCT6/AJYsAQZHvn65bX8m30QX5IXqRtvI5lUoYAOIAa
jVkqZS1Y9B/eadg6PmG4XQ==
`protect END_PROTECTED
