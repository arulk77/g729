`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJvjB0+hT/JZoUO46+8n/iF701wVjN5n+vJGJvMn+0xC
e0FGbxH+gdZZBsg5sPyyc49r5k7kxHyHzYllzd9s9B5RYj99XFOtgT3HN3kN47rN
cW5YoOvxz6Ixwe1f5pfubiNpU+DH9v2I+KLw5eTBJT8EIFo01yYJSGJ5i9VC7P56
h1jjH/PwAxWRyRRS04jfQwGxQDlVyyv9IY4LZITRWcpWdoq0FpLkSHk53r6xR3+c
olYyHRTeecEUX6BP+8ErAqXqy5aXQbodK/e45olTm9Nop+YM6qaQ8hl0/YxQ/99Q
wGbeCjOrjucXzn1Wx/EFX8f8c2HX++50oiMb3oI3/CoN4INfl7Bbsbu/p66Cdjqr
2IKnPAulORa/x7iAQg7QCOiPyllGyvRDUi0Fv1rOCr4gBsqwjVHP7/CvxybLUObJ
EAbiecQwgWXhxdK1tGWjG+G/OODclbov1epA3Y5/nouCj4VAuloze5JdLC+gj+wR
76FuMAOg/wyLoRx97+EMcMK+BMfzL8XFkWJD1bqz2BkBW5pddRk8nrwfhgfgSIbj
`protect END_PROTECTED
