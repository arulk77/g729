`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wJYzGCY9LzKosuS6KB+bzGF/+uX8dGLiiLN1yezzjBY
FAdNIxkMH6B67r9Xo9Cj6wuU61xij03qM0mDNz5xmnlbnO8kIKr2n90JEvzPmKrE
eZatbnl5F5c3pLDteBrB3PBcOA10yMnl9IiGbB5BhaZoz9mv9dLvHNC8rVMqhnMU
FKborWbZfKh9LxD8XUONAa33L84SO7Fy18waMJCjPjI=
`protect END_PROTECTED
