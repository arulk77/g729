`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveENIljaGOt4M5IMr3PaiPAY8d6liti5ICEZ3Fhy4g5Ms
/hAnTt2z0OAPnjh/sPytqZqnyyMqA4f2YdyfJ2yb1vqmIRSJiDL9wglSWC1rnFnC
auo304xnYgZynrB3tTSloJ51Ot06ytxdkWpzdPr7y8IKC5IlevSxreUp6L6nULdi
UaMsYvSjPClzIrnO6hMVNkTm5mWEW/roS1iVOzZVR+cSOX1Cg3yeoE/HbZEBF0Bj
C2YkQjNag3+9W6fxPBGWrZsrdeBNMzmakbBRrwpv/NBQx8J6FkhYWbZvKQSu/Pv7
qdWdNajQsF5kuFAdEabkvBk69GEVz4DLu/N6aBvcMkI+9GmcNF5D6gqn5VKF9bkN
dwb4aZHIKLX5J2lXYqAfKnSSoPDRLuK7Wa/5HHgWITXSegkhoMQO+wSkVcUeq2aA
2Dk8wKx7IuTcvVmpSPdKOLSdfS9kAXCviW6rfnSZga0=
`protect END_PROTECTED
