`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKoFpprSEWoXEgBm9yO4KNYP7QWGlpl2dMpwD007Tm5W
EmXEOuRzrsJckJh4yCH8PxYldlZND51O1/5uGR1cMMoCzel8KJQvKpMWWJfsZg2w
VOKj6MtbK+qB2p5Ov89P9uR5cGaO2d8Tzq1pvaArYnhxij10X9sx+zTiK6RSUsWs
Bt500oQ9PyRogHx7dFoh7LWNpIoSfwjdv1adSdeTr7UbxQhoP6coaCVu+o0bpmGF
wMpB4//dOJNwiTtrk9NSR9cI0z+S31+zs3tNXb76PUOb73iNpV5SGDBLhwOCPTdi
VnvVY0t0pi/c/u9BjGz2WapxSSXdinbTBFumzdAvKGOVaGwkwQaKBu4d5hqav1L6
MjZYJHkctev5yln+ggTgSUOl/bzrKp/dl0pdc3A9yqXqkiIK/D26GFuNpzoCW1Gn
oIH7EuuYggfsKwG9f+8+Yma99g2BnXRdJnutAMb7bXHLWB84RAl5X0dqC/xVv+Uz
zpljZaUxyleQnRoCEqtL/uGz1W4vpMS+v/VY81h43jo0V6amAZwiNB2ir1dll2Us
gelTrUTWWn+wXTgw81A1MY6BOn/nOeLJrOjfA5YAAQWSEsblwOn/8Vj6H6IWutDE
RXxIBea6b1c5/ZeoFiJyQ0aWBdd9TsYKNBakx74mZM2lXviJCB/WBdh7gCFvRbae
RhUEXcT0wDP6Y9R+zOAbIXWwh7u28SP7h3I7jlvfdGBvVteO2ITSyTCnxmys4NFQ
mnWHb+hcsba0vJCMiTjSLWk2TatI204y5W/neMSSqXYUxzUnDXYhfY2bEhpQc8jZ
+wVkR4v+iXPA0Iveoi2Q6uKWSLTreFFySeIWby41Jp2frUpj5Jc942znE5IPkrIV
XbCLJGHzafpIkRzBM+G1fSe5xUtzR0wmM3bF7+DdX25qLl8eyi9PEUmtpJkfiyCt
eAjYOlFDoZDdgw3Swat3H5K4R3+8hRdIXAlvKHdaEYf/kU5TA6zOfxUf1k/rO12b
Un3Lklw0wYbMA1B2sqy3M1Cf8HOQKF2CCMVjyu6kGU1vqf/dyz9MUAKnLPYU0APH
rnk1dn+o4/ErhoUZ6FlWC6JNLtNlTEnSXm0ES+sXwDaJgq5Hrc41D8DauuC1PinJ
mBV9RuJ8+TDd/bElruemeWYMAfVATostTfPtBWUpf4K4k29/WCB0PH00Tw4AQ4Jg
dTpKwBq2xlcZ2XSqSpH73042PHW3jtkk86gcfF7GkdfXu6MiRNmaOVGrLc/1NZtS
TXfJbhOFDU9fywJy1TlpLT5yiBK0e7qIOfPd+SnajTTiJaJRV6jy9w4nLFDnaWS/
MHvRfPAVATnOkp8Xjjrdo5Da/0uz76ziocVvV5MTywnQcx8i0jiku3f6DgJMslPb
gJoLyLeewmWiQBDlT1DPE0TXyIhhsvirtaONZgQfWiKzVhrkLQazOv98HoFGhaLc
HqZ+bmM+331hrXQ41wzJQxIkDhuMh9wV49rl2zmc9Lv6XBvHpJ+ZYRDJVkONppiV
n0tnqICrIIEjBd47Y+WMnBtM4HEinPN+6iD/szmcQYnM4KzeqAJ4Ktsw4fYsJI4k
uadR4V/2aSPBd7M/jFBA7WZiLO4hDMsKCQhwGyhz79rRdVkKQO2dPIvpmbGwvuDi
eL2oHBxlWWPqb4VJetPSHntCVPCJQL1u7IhGpz/CpBTzuayJ78w41LXPOQjW/XOy
U66AOoeBwscFqlHDvxfg2daG8hBZuvhmeh2oYoUNAEIj/sA/8/JdN4ntbNSztb02
ihZv3vgQ82kkm9mmg9EOf0ROp+xHmtQ6EMnsYVPdts5QGv8WZbHuMk/ZiM6ipaKk
ZyEIsRW6b1V8rMxJ9U6zQte6hyowfJkMW/0jJ3jTX4HhcaviROQmyrX5Pr/GeHuc
JQ+/IXcReIWLjqWltoq7yUe7rh3xNUq52vFBE4UDn0YOcrQjOzDmXtH9Z4jC97Zo
ZeL1fNiub6zJYKyg93x2hgwjQd3d7wzhkT9HTyP/sYhp+Cpbdcf00a63fflNw68g
HjViyHjIAQ1Pps0sLOJpjsli29sz/4cT2XdwKHrmSeRAWOi/nve7BSXsO0gzArfY
FLt19K+8orqGPchxXLb3fdhtxvPG0C8kPUFSnpYlz3zGKGuk2+HqB2BhgBIXhm0B
ZOHnZR9svjcoWutxgstsH4jhogvIFzYtj7o/VqPLUjujbE7DszABR6hnK55OTv6s
3ESP6UudwWbJ4s3GRBta0F5dwBDtu5qA7OGu737Y9Ylfqq/CA+y6D3RwhLogxkQc
NQ7c1ZLTQ5Ond5wnXPNR6hsfkVM3T58sV7plKRzM3+5C2nPibotS1Y1s+egcTwcV
h2WtO9tw3SOvSkErGgQNlZJAOsaBQtzD8XFD7fP5k1S63dup57irJ992IN9PBIyw
SWxIejoaboTx+cKiXy8uE8OZWwV/8oqqvQQ7/nNO1ljKE6IrYccn7ma8ymnJ7HgV
Wg4fYo1RdkCBM1ao4690qBKdCiHTqup9N3fN5yf0dLDg3/Td2TWIaLK3Gh3rKUoA
UJZ7PzJVvB/9OOrfutBacGpbB2BSqeATY4T1EskXyGFOnwRuClxFuSd8roNyO59x
Gg7VutgD2mnZUBhoulE0IthUuyVc1czq6gOJIFCX719wAuzgPwkZ5OfebNOW4VwB
spy08RoKRmOmLLNR7LiCIzqExidp765161wftiBSi6pfD0xbcg9PDjXllntf9uVZ
uotF1kA9PCHtLZ/K/H6E/kLdQndWPwpuA7YEBMjY/AvRQkCougjPqY0G4Uswjm9T
fvQkhInki54YY9UskYIpQKhdpZMDOmXiSOuRVNxBOtzR6gnVeDLiGvHiWw8202Cm
pS88WPXswfB6EI0Ma1AM+rbszN4Ck+/6SODg0Lx9NCJ3q1il/VvwqsVSrMdiKiRy
t9hCaMZX8THYHAgg2y2VGVYmODu+AW3UPOriymoChIDL/Qh49o5vK9hnmJv93Msw
fGjMlmI66OKdUc/XJ9ioYtOcNgbIVFNXzCIhx+VVL6ap2e4G4Y2nUO/Pfr8nXOJK
5MkBtzc9uS+7tBYRBcLXrPO0ZZ7tXiyZmzaLMNdJkoOsjbH0hWnMroBGN7dVzFzw
GwIJ4B+wr8FHmXCQnDXzLPYkbce4I1hsuFKhEZO8etGoxSgVYm+ZmU/2O7iVgf7c
xqjfEAPM4o/1U+IGFHknL+dSTcjpEWzuJpUeAD7B4PUkS+LJ8nknW6c6BNRFPdvy
EXM0Qrpd4RwOdjP6dSat76yt4opzS9AkROEdOxVXDoRqLJrgnSg5D7MY84eRvdQM
CIQoq9jOKuit9OSUHSBVv/tRbzLgdD86kkiBBxmZ3QhA2Ah+Qllz046Z3WXgOznP
X1CBe2V3q4XiEqyyfclTVhXovBgFJfieybkvAi/QGbHe4UTny58R1BDf66kUzoxF
qM1sYATiVsIUmzrzTi0JAHowjZoegoFDKTphPa0Nc/M2BQSFbTH0yrYVVuiHhtHx
w33rFk7sxYTIPTxBkMwN4+AAmkxAqjlVeiKaiO1UaH19NH5utjwDpLx/t7MYDC53
VtbbZcr4rM6HRBZXDf3e/c7x3yUmQUM3oJUYJy/6aUKp/NjbbBVnbpmYpvxGXBCT
6jsiJk/rqf5CvK745+BAqVP46uPXL1g9zPR+N28ft1CRR03V40IjvrT24AqhRWFV
nPwR15mvFRjmzC8tDHN7PXi6ZQIi3h7lkuD/HWlGerX+j3Ijg05cPwI70CDilz/1
+qF/A7gC/7TujiT/C/RQbgxICQNhePdOEA70n0wJGL29v8GUpHVYfcEdC5ZID4UQ
cgZbhNjsIHckGkMQxyW2upjZquGH3WdhjZhimDX6+db9tKuwvhHq2pEHJh9ZzPLI
NFRmWAf4GfhaJbBM2PjCsy5zTSegVkABA1lclqZVXWZkzniy44ZCWDjRRqWi/Mjj
DlKx2mZJOixEFWLdAU+JiGo98AFIemIVgo1XMY2Lx8YNAQcNiOWf3jtdX8kK+oif
2Tb8Fgfi9M02v8w44xyMmqfxlaLfvkOnscu712UG5gY2JlGCpFqeduXjFYxDVE9e
eAx92PQIHXEBYcSZ65PVjFsVDQJtHdRUJsi0lae7xq2TYIV3Rux06KU3+kf4PGHh
K43VfU2SS6xyqiSGGAayEfzz1UMMpO6wWp4fcDwXun60nFGHvwET357Vz4OHfjqA
JojlWqcpEmczdOIyXF9QtH/l4iKwNiw4p+KqBgRLRjDztIgKFRV5E6wJoG1PvqaT
fl3Ob8Vd+0MzzyfY8LoasQCPssUgWzDBjw27O2/TS7vavKO9m2DpWbqolujSOVW/
IXg9BHm5nc532kIO35JmRHA60lGSjA4+447cbn16g8w/y0anMMl0lTT7Vpgjrddy
uwACI8tnKbb09D3CFhqYs2EsyQXubXHrAHoce3S9DeAjSg/dvT93uBjK7WWe1R1U
0rtrCujucNWAcsUOkoxVkgeVGD5Cu40vKBcCjS6q3+kWpH6euPRlXgKM7+QcR+Zd
n8ALbp+YyXp31XCLrefc6tQCP5iQib9WaAxTV8vR/JdAzspC8djqCScO2nvVntIH
BgW05YMfaros22jgo0G8n9CkTMjVhdeTSW7E08YEcmhEx4n4H+Ay8qq7OstmApEZ
VHrNOQpw8oYtKJ16f7e9488GEZMQOauoVwAeN/tZL8IgRVTIxlBN93QlVT35hjuw
iNDmLLEeV+zoeP3i28zwMv9ePocrTIimo+QS0XHmg7jY78OaCdUwNv2puNR4wSed
oPMIhOKffnP+Z9S/cn/jVPwfdoKub/mcQdtiCAy82vraW9VJHBk8R6Tp25glUP0S
2YdcpsRuDWKR1jCHH/GGX0hgTizuMEswWnyVQ0qEkK17X10D6yp/7sokEXyX6h2m
k8Spu1/QUf3hhGpSQk3O9AKBUUo56hX14fZ0s3AOabgfmo6S4US4VBenIlruQJ56
tNzRUbJhYJ076Zu7+JBjsqa3y8RWSJuUEBSV7Z901uYoaKzd4ATLbGhblM+MLxO5
860+k3H3s+fCPfKosfi5BKVhu+tEoKJ74DHvoP++iUQenmsQg4D335y2MDi72dvZ
Z6qQwBjghvnuJhokXxKqKoLANckhU8Cy/JcOucRpoJAieFNlcmGAu7kz/r0ZZ2Bp
6ljPBgZE7eFZoEVSfdNnrXGHzkyBG5xLPD7RJzX6H5EXeV+vpINCstKKNZ334fIl
pym85hZLvYwODY3PZjW3vH5ldHXZe4/qvhPk9z0dQxpW1HejIMbgrAfFZtGfH6B6
Cy21lWdDT+50BrzQ3A4aHGPPEMZPsw9d6SEORtfbTBPD3bENB5W74OJCaey/T/tG
XkehTB6D1kCKc1HbCilMAZf/3d+W7ttcW039NM63EmWYRLQLCpQzjyL02IoT/ZFN
ecjwE2kDt3icS32ygqpRywa/LRZptm8hhU26hvKZjg0Jnw86EQUXa9m2/90K+ikx
KdBvjDDuIdfuvEH+EuB3aggr2u9TPhLwcR8ni74Xfdqv052enuGBLtrEYYON+lth
c06BeOOrNWGEPOzL4okVOtZscEmrdJ+Wqm8TddH8R3AUK+cxnRljEkubX5r85apc
F7z4C0rmVwhrI+xPnzW1/bTBPSezEH3vN4TicaAxTW+J1LDsgP4CjO9eNjAQxW2L
jYnr+7e0+iPavn/ficMjT8nJecdGb3dW7qlNnLLYkOVIZxqiO+UeDFVV6fTxwbY7
UlgAWKyJwVGOMN3CuqicYUk7/ztOhITA4KgZci0B0AaHfmIpsAisQ9pGkCGRYuuX
AQdyy7mVw0oHIU+9LnsCZWpUELQ42o2cERBjbyNeJirD4gSOcTwEGj3rkRiDdi5B
OxT4jfiHVjoNqLqi5hLdqtnEPk+OMF7FjhT/utu2dKj3FjBT+A41itdfdLvyoM+Z
694XRlyg11a8Nl8qePJ99BAhQO+pCVJ98/EOA45xPenmtyG3CcOq5AcoXqhGnL1L
sQaCRF9ZjmYEV2NBfvTSJkzrMaNSB2oSMI7KsWgTM6vzfL9ct6jui6xKXfl4PlQS
kWB5iLnSuIwuYb5v5gowDURWj14agdK4NbiYn1W0UU8J6fYNVrnIswU0n4/ElQo1
4wc9P/A51DKLRVi+Xinqpc1piPf8fokWP4G/H2ttO576C3v/yqunwv80RWk01PIf
/qPk22OxxbGOxq1Q1UDt8SLkEcJ0exxicMcrtPMgUG2K34s8w6Nt7m56ecTUSWsC
9VZdf/bjPPsuHPVYFEclsgmza6YXT0ZO2KhmD8MyvLSsoqgJyJigcVA74FKLm51z
pQfmnZEMOUsXvNGu4BwA598hhmfiqv3nS2AaNw8Z1t0fVu2Q4TNTRYwPR4fuuv4e
ahybWerBaGvwmtfhc1laljliy5ueHY8JAH4yHUTiUozZQCzqeqbb9ABPeDT3R+/s
l22+zv9xCpa1WxLMV0xKPyt9NNOfp8KJvfTtJe5kqWKeTAfD4ERwdyfT1KotIdly
sfmhf2xNa2j7ik0VVm5mcx6N0NYQYT7rGqMX3f94MpDkNUN4D1FI9eYfM4NWD4mL
1uw2M/6J33g4KeVwNbDE1yEktqrPVxJ3+MLDPMen3r94rFJX7vX9v/SzOcQTYoOs
j7Z9yIsYIn5jYKYWEA4SOj4YYEtLkcCKj6+CrdqygDxZNG5T3JbQ3zv0NCcOvI0z
iY9zHUlnmyv2WhzW64OeM5lz/oHISHXHx+omMpHCsw90EtR63pYSoWz9S0KbpATV
r52ySDAuTa9vSNRY17suQ9hU0jCAHnvk6oBg55varFt0IKS8tQdC/hgoFhRCWGlN
xEZZnAB3nAG0T8TTuLSSKxcNXqYt6zwTEpUq5ElvywBTX3ms/R2DdMwLUB4TAoIR
Ip7qjR+JxP5l8DcH+++tlk64/+TpukB9mX+0ThFt6GdVQpck+hidznsBORIO4ES7
x2s15mZZsxw43dWYLpLE/Oswk3IUzY6wJkvk3Bk3rehZmyV+5azX6ti77lyrou6H
WeIdeZfvurvh6mcLmY4djfZ67Ik7AY/tT6glLrC4bFHd7nk/0RbFvNf76CV6Qo+S
jTzVtwXZL/s+OCF1R5QxnloSaGj1n24r+2npH5cf26vKX+YluJwrTvUEFvGp5Bsy
5IqyJTMkDPDU8Ji/WPPqDs5J+cf70aU4Gwo6+g/F4X1MYlak6QJ2r2vnpmX5AT/P
af9BDJBw6SlSRsf9gJhQaKEza6SkQ/OvwypgDF3Bsij9Hrt7w+eYR94pFBmm6UDT
1YAe1hfIMkiBoOlDJhZtG3hFD483NAROdA5wus75//5n++s4uHiSBdjp/1eZpERs
aeB0e2ZQEpnE3QFzqVSfOQGaUnOOk5ao9/8eMKT+JDyuRfqGMsyYLQMg9SvKmWaN
7MKPWFysPYBqbyTVT101Z8GLvtNjjU2MnugPraLPgrxrazfI+YhMXBqWjjzD9wMz
tkSEWjAAeQZzlMMKgazgEyOfJHabKdB2F/pzLKp4ZZun6IQIh4FOpnmK7QlaT286
mZglNW4JVGHhqK33SgB4MexEJo1eomJZ/rKWHkr6F4MdCPbFGiRpvTQClMh/o6Wv
jKWZ+6tL/LT+ywR4bs5YsweYWrfCUZptKZM9N9yYXgGy4M/7jEUcfHkP7CO3Gwio
SJqVYkYU1zTQb2O5WgsiBrAZPQLCqTj/n8AXdn+RNgGYBGAN/yFUT8wbeMxQDWrN
QxgNR9SrdM3PU973+HuOlSX0Ej53e/wmqCOHIdHNhcimdltIVmFuDXfT9eRsc5Hh
1cmCOx0U54jDyKFUAAgW/omYBsvFfJe7nyGyngj7+LEWQEzNC+ICgOPMl35x0RA3
b0eRS2M3fxhHmMsQbn8NEglbZm9c5jpA4Fh2OM8nW48OlGncoVeFjjXInUzCScjf
5kxYTJ4/Jbe80VHSJ8xX/henh4AbM/wkjcQg7JYehzwv+FqjWDrN80un56reW5Vl
eM9z8TvbR3D7AXn5VsXuCqxDBZHji3vKWYQJnaQRqhZ9CB2Etnrcb4U2ilxghKwf
cCs056a2p4f7SnMw39xtbUG5SfN7Cy5TQziTZaM5hLdJIj2TEpmKRv2g8KwUvFlA
AGJjfhgkJ6jVGEbwuwsSfqx3kp51LZGUcungDHh1tPjFpVC9iB/NSmzseK+KMu4c
hhXC/3rX/kEPDFjFz+GayBvu0yV7C1C26omBokusO9ELbFDLb7XKyhajxQYDZQ2i
ZWRA900uiR7ZfKePE2c/jsCy9IJWlFB7MAsnadfWgIIViLm93e+VGJxrtoTZ65PP
OuBWrU9ZuxOCc3YM6HoxFTFvZcHAxToAv2jbHbn5ajjP8kQx3gmDAaxuAVd4uvrG
26rJAj7BzOiHQLjtQ3WExbfiU2Z48sXzRtzbcTIxl7fp58wXkK3LaLR967L/HPqM
ZnHMwaTjHpxi+c1g99k8rsNsUPsEyR2VsLsNTLJeh0AmDoOFpPGWnpB2j8JwsoCI
+uTFYevSwN7wTmIiKSXrx9Oj/WURwse6e3TDe+llaE8tfX1j/PElq/h4cnmjVqfs
fDlOBg+96c9AlSAEJD1SpBGaF/+S+qK08A/vpcSTXaQA+NYznSrNJQ4vCEvgwK20
zBkhjUVzA41tZIxDv+qJkYyxPn8nT+gw4RfLJogyFkgpDG/N+3rlpEJFhvIcy75b
cknn8DPrTjQk2X+OtIOosKsG9hG1UJiL6cLvPKMAMN2pzfCrtuqYdOplQM2GYSu3
yBx1nCIfUgrTc64+aXXgAOgYKi1kveX4Pie2Y8L5B8lXiczrfbc3kq86IhhyqDn5
qVlzDQdMfEmm+HzupuTHKAwkb5SNiywOtFRhl0QBAd7v/JcJ2N++DiV7mMov2e4S
cucjow6IeZOEjM1YQ9/2Q2GIPVTay56uTcYbveUdnJIBjni8gOZZK7hVC4hepX0E
L7Y8Fv8oUTZgdpERvZ6jf4k70LqQnq7MKidaTClbSxsuef49LWxOLMhxqbQFBuXr
89wiPTdBeJZCztCj5/KE5VhfmeK+WGl3D7853q0poqarg1LlA2dnzMIBYmiMLFcD
eKhCWzsQ5T5Mjl+0tVadY3AEG7vzQIbTPnBGxi4bPeVVJZFwoVcXNUXpFMEJIMFD
z6fUDcqDEtl6jFDsuXF2ewQZNfofcmjzF1BiH/tzUSEHDfkPISTHb45TqugVhRs/
UfHzzyF+w0Ls5WWmLGPgkv/CwjpXO9uhtyZ75OQr3rT0zIxNcrB2j5ABngPEV1ex
audDo8AeDQFPtfdXZNskoZQ+euLU+G3hfft2HyNocNTshr/6ZmqT2mSdoc1mlV9r
iiIdVq+HPeIG5vrnhCIJi4O5a/3eCATPRw0tnCY55iA67ZJkxZUtbl9JnsJflP9X
cIifYLvAQHP9Th5iHkht/WXksiQ9jSRnKZfFi1IFrcRcL74OnqhggFLtf09APg86
/jRTOfNr8oIfhHIylYuDqkB588hwobs5tGsSc8po08K3BXyk6O+nuw4wacTANCiE
OVPrlVM3+3k8mDAmFYE4kbkAVFpvmOLwsl9xv7n29wuZb72OF3lc27qIgVg9Ka+l
OKo+gAldOIImOxteGT8MrNGHyG5+aY0cB5bl/9zT8TKqrRPvZhLJsp/ZFZ+tTNJu
sNfQagYrv2U3dK9bEzNhEH7yz1MJsX8fA/h9l92F9RvSpkewGgOWRj+V5OgqOX1K
4nyH4hVuF+UNXGMESAa5xnRhGQa/SYuB7GLZkEMiaLXxPAWxZ+BSEyKH6xR3U9jH
RtUTMzha9HYcrbAPh5YDpFF4Q5ytIUs3OO/M6OvRYU+A4UMigOhpKAreo9xbYLWr
8FGWG2CL7IZ0Ufi+R8BCi0hDZwSkMcXVdUTtgFUUeexRRHfsJMT+2Y0rC8atOxe4
/tSb/r9aR6JOqOjuWkDwpRMAenIhclAXIms5paV7czmuUbAUeIhyZtMeb+x353o0
Nv8a4x+pcUxjaTfpBBhINwiENr/IsoN4wjkMZb2kdltconflADDuR0FgN8/O2h5e
Lcf+HtE4u+sq2sRG51BI4jkHQyKIPCZxCIilLu+K9MXRZp8ciRQqhlOcnrNEy3kH
aYFH2zyhOChf6EVxntw4djKSfQu/pDWxLb9bJE13GJxDgyqVOb9A8DcquEmLEic5
Sigj2Gpg0bMOjxfHoM8B3IGUbqIFJiA1igk+fsHgndJ69kl5VsvPF7MWP0m/peDc
Zd1mVx27q00MyBaAgkq9vbgjQ7dfmxX7ZTqhluqRf5yXPwR41SxKcka5SE7YzQOX
uC/Mrsltp9a2uj+KLixAfti9RIxTxU9Qks3Xw99O3qN2V8dL/FKpfb+xoqcGPfRw
iZkFhyu2YErDSB04RaX+QqnbawS8btKSQ67gB9ayp4ZiOum3MrcX71urvEPyR/H1
P8h2v96dNqnUkp87aHyMa/YihlwdHWZd61ftFLsoCjziU3x/GDk/VUDUVifiBKKx
TfyMmcKMRxZftevtVVFjAMIQlXSz6ztV1EQDMc8zkgjt0EbsGQ9LDUZiIDyKnkLg
LXFmTWjVhBExZq8yQ91BHuc7nZapkJEGNYgG5ZCZjb6li8j80cOvQmzId/PqAeQT
Guo5MHmKIPNeDD9SM0kI/3k8JGCMTa4C/1dxO2Oks3RIGzZ1bLbMbItWTemCzf4H
3riFsDGQf6CPvWiyTaI+RVesXQ5BU+ZQjKyTbw6VdROV67OkRzPJCU5Vi2j8QNxl
qcylE3QLs/ZHf+IZYW5e7l7U1PZGDQaKxvqO60EZlGO4pqQv23FktS3/0HI5yBzn
omW2qM210WyMPviUEsEvPS5gol+boGgNOuvWqGGNzNKTGBZZxsnjgBui3Wp1kPSU
lBhQM/jFBjNsDT749K0VmcnRmUcjRvkRCnXYiec/upHefA97wtc29K9CUlzRTno/
`protect END_PROTECTED
