`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
S30LyB6hfKQ/SoCe6MG1w4GLRz6aTOtWZ1AGsS6RRV4ahVoRvpMVKFyOo/z+1tKb
JmkBYELHqgG7JP78Pgp1OeGKk33RqfBZ+yERDREJjj+L9jK1xpMRX+kcrghGTKAC
EkDiO98lTC55MdSWpyGvqLbqnH6IRH25aeV+EusnkWXfmOVqOkRSR01LuXP0H5ED
+JV1sDhivyYP/UWBhDbzf58R+nOZIqNtDpb0KQxCeMrx0szuFqoYcUNfBxTMu+dg
vMsMecpAUL0S61TY2GxQUbuIc5bN7zookTIowdTxxM48zkgR664AB1fTp5tDCO02
3Nc2OTbYQBOFGjWJqQd4frEkmdqneHLNftadbArJotKzNewzVcw8UNoREodty2wi
WzFIr5zuocGlePZIiHIaP8JBbdqPRlP/MTdGK8bRXAo=
`protect END_PROTECTED
