`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMm7vgRfsNkyMzz1sMLXlthNPsIhvA8r7tN8ITZ6K8qB
Ca0UbZ99BcwI8imMfxkBCdmyAk31EX7v/TdQjdeZ7X2hVLcLWZ6EKHerC1ZJdjqP
twLNdj7Okp+RpJSAHE4Hs+Vg0i90Eh25rALVBJWq7hC6qkFxnOrML+MWPXoVnnBl
fJhP6pGremhMsjZx4Z2PepNgPg7BGUS05HcxW6ggnmCrgGe1zyYeNVZKL9BqmLLs
`protect END_PROTECTED
