`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKRBPt3YVtMfc1thGcwAAfSVUt1co3NTrYnQkzgpflrc
Wc/C8doQc85md+Z9Pnm6MulwArcyx8UhFZUxDpLyKCOqqDb7LzlKmCCqE//WoGIY
GuSqoZEAUi9qdLfkcVf7PFXo7+65N1yjReicNdCHKDDHvUXoq9VLAL2alYNX3LBs
3b//Mrk2vMnIp4NWhGPBB4n/DO6tZSPXT4CWYd6EmslDyQouAlJksEvq6GzSFT7z
McvapYWGI+Gu1FS+OJn0+9zTLKMQVHEHB/LXpBdaMGEzt2kAobXQbqvklgn4ZBPr
+Al6kj2lpupsgt62vuKzV6ID8CBwgD6jEzurNxMdEAN55kHjnBBgnH6vo3En7eLk
XNAC1i/xUgcJLhewMR8JvSNed1z5RPWlQJj2WioW6L9pBTqn9fhJNrae4yr9S9jD
naMHpayQEE8mPhZ/UPIsmkMvyT0oGmpxp/W1pNOOQYIqyI8YbpMg0cLLFQqepQJ0
hTYNd4OQepwWvfcI1D+4zxkRelsTfVDCyfeGRW6bTNKaSihPkqbhUuRqzzHyv39w
OYv5NYilT6ANfreqRAG3w73tL+mkmT7gW3CnMaKebWau7Jc60u/Q+qrqRV2g4MHK
dviH74AoUepadWOekEzC4A29RKajVUAhRtOJHTTR4wBnngZr6e39MOZItxXvpu9l
x/jLsCb/NJdMCz2Ec+EqhosiXE5uP7CfbhEAEvzgncj3W3N0g4k9qeATR0sIp0Tw
t/rYHHcfXe2n4j9Gonl2pQGBlqw3AF8tXEOKtYLEUR1I0fJjcH6ks4d9ZcMM5AEB
9FECqabp102eUezmswMBNtW+C/A0hCMCegaxldSXUio=
`protect END_PROTECTED
