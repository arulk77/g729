`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
W51jmh1BsJtfS1cvfw1eafdzG51Cf0JaFEr2XFX15F6V5FxomSXvB5K+KkExR2p4
HpiG3HdOY0lFZ8ivK5SIan7emjAyRaV7wwDjTqWpFIrP0MeQcr0K3qfq1VA/mvk7
i+VBAAaRK2uZJgitJpWn8xo6lWYtVQJQ16nx8TrObqnhpJmN5vopR2vwwNQiZ8UZ
qB8NL7spp1Nk+KK3y00VjXjqjQYdVHW1ATLwnjNJsQsO7FIqDxJXe/rHOzcafpf4
/Z0jccPVR9tF/g2OT/iRCtr5kr/5xv5eMnbf4ll2TPw3NkiFaIesl416+DdoTM9h
PYsIovdZ2ZOCP12u0eO+ck18xNOb27EAPJfTqpP1/S7XwJOXXoxLcgpxG2P0d2oV
jrmKhAqP3n7l5L8veQBAX12GoYCs66rrG/XtiSiYzabybz5dJMxSP3JAVa2uc2jd
xxKuBbvCIBONwJrPyQJJ8B3lou3m3/IKdOb2PmvojJuk8Bk3/yC5iea+pIqF2d5l
u/H2Ps6A0BAWmLub5Z1Ypvu9hlG42y0RuIoODERkv1JRQCG3g/hLel+1GXgYNZXU
B9wPDybpHdj8ZEySjihDk+3Rn0v3ZpPkRPtKuThkQbVFMIakxaK89+wNObZQzXMB
E54+U+WOiEJ4degS3Z7GtNPZ00Kx1AEaMrb8hMQctHb1NAh9seVQ/Nxc7MJteapk
VFS+MEDCZ7p5QR/713MiKHCFLLyZkOO5OT0JlUOrp/hzBNT2VnoTWuXdp3Vw7y08
KUbfk09r3+inF/oXDWMSDI67/nvidYs/foZz3VVWqm2XWiY36OPmdO9sWPFlcMxn
dTXKllP+7MjSKv1+Edq+SJoxUuJewktg6hGuvNaFxA/akWXvr6eYVJ2t70AdC+OM
Ok+seRKkuznX4ZRkoEzP32nYZP6tqoPo4eT4dmposQk8b4zZPdyvLi0zrcthExX0
eOOSFtEG9OU8xDIzqRyLVtqg3lGEMhs9DkqePag5Y157Kwue3mDgFpWO9nuu98Nq
3uJJNmPsw27sJQjK9nHcOqEd74drGeNpp7/M5CFFcBSOp4ZIfgNiNYrBwV59tJIa
L9DVFHCTEyawp/xVS+hbolA4fATsa/0UPfC0m5TT+T8+KnjWGY+pA1k1bz/5uUoV
ZtVd0dwxsMVzuvG/7MDOm8FA00CBYwSkTYXWd9VAdLEhy/sQaLeWkGqNZYMFtzcW
Vs9iVoWpn9pxz8VY6mgeaa9RvzEilPrPKcbRd5x4m2t2daYKmfxIfnPMoukWhRMG
AWbmgHePuN5c6Ixx3mCsJ3LkhHvumXmssVzRUtdk1OaCJ0jU/KZ6B9t/5Wd+60Ox
DQTGE4eETKgiX5Q3CBemvgbKO2i1foEQ2wRmGvJKyGD629F2K3PysKkC8tIqHkwv
kmkKl9aP692DNTLU4j3gWyINQojYb/fYdIS35QEijG8=
`protect END_PROTECTED
