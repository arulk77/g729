`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu433yghpxdIYHO/+pKmA2TmIPiTrPswmLAjj+KEb6qmHf
bkDXJ1FdAThx5AArpMmsVdMsYen6oK+ChA5fj31ZjXKsn+wBjmr85X1u3Myozrfj
BEfZnEVS6Lh/fo/46sKz72FELu4FaDVU7n39UX5PXt76D/26p7dAZIOLhsP551tA
zr5O8yH9scIPlfhkiVkB6LUP1HAm6JdNiULIUlFWMpYJNCfUS1DA0FdOS3yVPr0E
tBmqwAZNIO5MNQvQIxw81tzzDd5YytbYME5xQvM+UiQ=
`protect END_PROTECTED
