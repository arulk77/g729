`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
lA2omtyc34Avee1JdYbva/TpaYt9bCe9TA/aQrycV1OVkklxFq3mxfZuCRzrjgue
ZmuocqE6V4jA0TpNiz23IqZQa51P6JWAfXm4qb9nUrCju1JIctGmmpj1Xmt4l4sK
`protect END_PROTECTED
