`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAIt7ff2kMOPPvKpWEQ87fpYYu3uUJNvHUWj5uuEW+S4
Ghv4V7dvpYIqvsnEqfwE2gHxLaBhxKQhyCFJ7wdzgkcAF7YRVAxqKaTSEWrkVifN
4XmbNXQwMZP8iHRh+FqviUepDxD0k7NFElOwe0lTpgsa8CJxtPDZHqMHkdfAQ9Yv
eIWMuyUCUrv8oc+bBer/zUnZgifu+cCrUgbQjeakcCsdSbrDejOwXehaEwY9da35
`protect END_PROTECTED
