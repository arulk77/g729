`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHngmEOtEKFosEIAe1lxmpec0LGvtnIORaSFihlx2LLe
ku6dZiE47vmnAZbiRD6FrZgvcVots88guz/Zxry9IzB7uqO7fUbua5SdJ5Y7jcNn
rcRADgnqqgwZZ4rcrMk7P5oD8IJepV00tDGZhHjs/3Q+W3Gfav+SBNtWOx6ZttM3
zlrwImVKtnAnhqD+jD3YdmS0mVNxpgwYzyu4eagxdGTjTJVaTlOL/G+4hYqWZ7XB
hQXOUV9qWX8uHDCWSE2Fu4GuycV5lxhZiNSd/y+gbIEnNnn8+rGz+gTYPTboO3jH
qsctHD9yjTVvDL+iRqmKW5i2LRH3XQQ5CJ8A0q2ZrKuXt/N9eDeUSdzzGCNUEa+J
OkNgpCoFo746zXUtaiMxukQhUDy5bKB4bp9S2sMrZqQosgYcANSF6kLRVdCMsGAL
i8mJhiv5bhmpKRQxdg+Tt8Pv+KNhm0n5v10XgqA7ED7/z/2wRelycY/26b4Xa7fY
QvDAyn61gAtA0duPq5rPS4gfFcWl002zxnF8+qMf9jhUi6IUgzyAr+4AG4zM921p
`protect END_PROTECTED
