`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDbpDyx2Ds+C/9xqJoyHAZnmBRXJIJpST4+FFOmt/KxF
SzyfRF+vA9Qbn6qmbyWPLicy9qachHU7wtT6Tr+Y1W9z/GiK3rs8H0wEVODso+nc
4IkgArcqFA6GhmmaVnoeuY7L2Ypx/iVe/fvdAtaTb+VFKJrDXSORA4IGiuaNu0+d
Hr45jN+6B/bEv+I9OFEkNXVzo7mY7TRetQyjqTcs3g3bR4YvQl9JBstav+DYBjjt
JNT7Y2Z66yVnOpD7WMAVa8cZYCDouWlBzjrWeyfBPzIapaltfaKCImPmbT5JeZzI
`protect END_PROTECTED
