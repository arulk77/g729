`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8Sdm9I3/7msGm6XvFHxvOXVXwKtXFYJGZdHq7hfH84TDF
jLUl8towvvGHZhXsGgXNhWyFkFMd+A5GvCUMdMtYYTf+Eh8QunhhrTbWHp0VO5YN
FWUyU13cTHdKT4uKSU+4Bd7zYw6RGMT8VeaHQZ7iHPVMVEsWRwM8jQ6PG9hzv8uA
FL3qZ4VHNYlVgAwXTcPicfzBksSG4/0AJlCmOOBOXy4paCMWWLwSYZnngyP+UIkF
jz2mVUx4u6JOFKpvrUteWoa8znPae5ltBZWNJ761c4sPagk590YlebXEzKT5cQEn
b6jv4xegJOYEXsEQNXmOKnEmN0StU1N7CAtPqpEpNkhTicZQncNJ0AbQ27afa8IE
B/8l6/af6yZs2ZmQqQ1YJJCsyVZNt4zmJi0JU8s6wc4yF5w+5Y7NxliCt+uYQTu9
cZdHGO0JcaBqDGrazo5E8WDCNADjzcA9cl0KhjbqPSdTatkze5T7CNw5A5AmCDvF
H+ncmrpI3odu88oXSSPQpVPwA/FuWN2olmuBmi8Kq0tN2qz6hGiiVhXV8cD2etag
w8Tp0f3fJDA9CxUUhIOOvAsUYq8UatWH0QseVs6SGGo4pajlRS6mokXT9I9NboQl
sU/0BqHkdpy2Bjl5LQeKe/It52MQBYEqSvOPL3CiBfqSLejz16XYogLI9Hy7qTI1
9AVOIbZEjrGOD20aw3VoVRTXZs2ZsNMxGG9OqG+hj4FyXYp4cFs1xthGGw8EbZv8
BHe6Ux30WGJwo1bVC10NirETvIgNbnpxPmtfhlqShm4FZU3quIOA2MkLK1iVYYkg
/qPn3ErZ2JIfSIR3hC7DDYjiKDfIEXC4xj47ukKELgARJfliXn5fbi7oWAOSCA3J
K7mp3Ph+yQcnvQNao5BQsclxLqG93VjrwPabBeYE+hvLoW/X7qTfACab/aL/68zr
uTclZqLckrnF53XBNc/89fsGa+PLptVcwJupXs8DB6MnI5WvwAG0hi2JZdv1zmLX
p+sfnh56x/CG0ZhrxSXCu64sw8qQ19qy/c0cxKE6cYdaU34/qBbhSoFabgpb5Ko/
sRGTykwylhz9UFl62wys2WH3ZcxyRyhBfk0nv/KV6EjjN2o2ByQLBKwL8uCCK00t
RFcvJ9G7o61AXLnlWo/OmA33Mq6LvOcyxOgle4fxoJLELRWlbKVFkVbUTOQsAgD2
0POftNAfvDI8myIJ8m9CGvbYXcFW2qgWYVmbAsa67DY4WXguLVm4aeTw22GXSXOy
l4RXkHs0FxGHGHMqRjIM7J3jJdyhxRtf/ZopNoiGWthVJPTPDfAm9DM2NIImK8US
GCAZuEjW/cY7qz0j4Kn5MhLiARXEDEi9I1cgjUEOHP32AkUBQaj0jmTRIbP5a0Pb
SDISbzYv0UBuM8ptHLS/YFg2qfMSNqcQCyO4rqGd3y9fKqIKh7M8ZcCKhHl3FiSQ
SeNtadJ2Qn/F3F+9zLmuFWXEpTWk+zsSOfxEzFja2p4Y90wqa27Erm1xw6wvZbaq
XcT7fMAWFCIqwMzxNjg6Ap1Wb9JsW4yFltT49cqj06hjoUYXDy2VqXLt1fqFf5Y5
E0aEyUD6/UHP2/4G43PWj9p8/8rduABRlOJNk6Hoi6u4a1mjhzvTET0pIf1MFHHo
xtOzipGUziUUqfndOVXKahhOY0D7Bpt3UsZnMThgxlybQua5YSI6leJyKaNzZpmi
XjeqLmUZZWu1jkUfAA0u3+zg0XPPVF+3lGHHRWDQlbN2fF+eshppYv5doqHXT8/U
vHc4Bjs/wb4uJIXLkoimTFFqnk4eq3lF8sfyda+rxySzgrV54fydACkx1jNzj+cZ
vctEkgVtGALtooaL53JNHeF+DYCrWNlUMvy3iBg67ZvVfcAQfkHCX6bp0CqaoB5p
6DAHA20ELeb7cg6rQkSQuntdJNwzHkIHU9+rJ45CsrjgGuOEXbxd46kAROMeN9oU
lpfJGLsU3JU/cyCAP+jVLA0xMuDfJJQ1GkW3b71j9lGqBi3Pa8nsaU9S1A9ANKjy
fNq+Tg4AitgCysIAy4ySPsLObrcF2i1C4LvGrUTU5uceGJ4DfMFYk1OifDw58wjq
lNbHFCo612pXttLCttvp6psU54H1nuzTd2pK6ILnssLK9qKzG2cdvHZp4PU3PqQP
5r4Z71Al3bLfnyJaG265Eztc8ZdwPE2PvhPcHgqXM4UV2I4G5pZ0xQXxJBEZxKMG
uCPA2A2BuTnXQFwB7Q9igi+4jgN871hWZ/050QQVLTqqnqcm0fAEgq8T8RQeEK5q
W8WJ9xYnZjsPKScJa8JzITLmD2C4NjD1SLN5rB5OEqE2Ga/qfTR/nODn/WNtoQ78
i+6jM/H1tN7c4YsyQE5ZtJlpu6WV66nCB/2g+gBYbDkUi4OJ7tVMl38PFvrr3c9W
2nOMePHuEMrD234VC1F1j2YVYQLgr2u1cBM6EDh8qUGX2gA0L4Mnwy6KkXY/kpUG
/TmCAhjKU89/NaZ/wcg3vE42sFAMBLTTsRxMjryBYCySjsX+HD7aGRtyvkLmzCNM
sC5pCayuZH1nE3t9oY/Q1TpM080rbepmFFdkEuvY/ArJOga4auPTgVkpdLBevcjn
1UFp4CEECmLG9i1wkNpoTfmHl9y9RuLDXxQT+UZAZMyP4CHBiHxIOC+oCXNyhyFf
FsGrkJ2gwLJnzpa9S3bdq+CY0j8qccPk3mCbmN8P539xRGEH8nhjk/kMhUA2TQJR
eN9GJgsjuAGcherOXTIe3iPTieDS+ZgbijfhIsm5VnPZBpeHi6R0nS/lLyAMu7GY
qT4E54PU89vXVT13IGUdOqb+EzFwoDMh0Pb83ESX5QfuM1OEWYXXkORm9PviHA1w
uUmq9UGLVms/OOcHeoVSRAHX2CQKwn5RXBYeq51/hgik3lm/aL6YVQ1J8ZppURxF
uOe2hc2eK5ZGavZ/o9D322HjX0ZDpiHqEtTDsdCWd01cG9ayIEoYmQmG3NtEfZvm
mXr5nmS2ZXDjP9Epy7mEbRn2DIP8lwHvpGK87tfE9WQhmgHEdy6QTitPRV6TlJ7u
Amg+N57xOz+J4mP3pw/2kopnbUqm1ANqkQtOjxuueWpq8TczptvFl9pcS2lch8Q5
oIbCwU+tgJ4SLtI4E1Rhs7O+5clo5tFP1RUPYmHdR86/c/IOxmTI5N885SQoj33R
2TGjIoE91UQgVMXuTJ5iZuUD17oJBXhQRw/fFLqOXkscDuSKmYGp4vuKPAGm6aYP
yU3IGtNgCRETvKntN7/dx2mSrji13c17OuYWlflZ1B1AFFkRyS4xXe3wanz+Lkrm
n+8brdO0rp+pYJP7juukYDfRae2NYwdEJskKnXg3gDL0Bn8VI5co+xCgL6Cmcuyc
ThwZ8alEa1q93BY2lgb5waA61eqhZaiIYDCjAQCBESMmrm2Lp7gcDhQMv6Kn9LBi
uxpotSa8LgBXLEmwweNt8JroiVwaLZ2WxVzLH8xK/UYZXTyW+rl/zAWm1Rny85kh
Kuyko6HfoT8/P2uIeq58d9AiQrWNyfWeCEwTFi70hWG2eTRc9Sy2nrhWruIY6QIk
7+WmcpXorDauCH8fqeKC4U5EzCat24d3nEeNG5oXxOTIBUwqBVRX9f5RCe5Tl0PU
/48/DFDI2OWG9dIzVuvxVf7KBaX7KBdbSx+f0DGP7TsdsSKkgdfIVW0f6kunfBHt
YHXQsYwrZWa8/Zv9swYLOfJ58uQpMyu0R+53HB3EsedB6EdG9cKrU51ZhsPHLFKC
4CXlo+/f7h2WIpxJ+nTGZlaCkW2rVAG8rlfdCy9l4tPB12jj3sYB8QqAQ4kHUx3f
35EhwW/jGuoANwwhr03w090HOiHuKwYRTZAi3TjmvDjc+DbENy7l6clxkFrf42Yt
B4PpOkI1p6vow1gec1rkG8S10DfKvK6HnAjJrpOVLMPfMFwrJ4xC7tSUkjh2QF6b
`protect END_PROTECTED
