`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ2GIBp9fSxtoljqJGwFa0BhUbM2XQC4Ap9MIPNHCEQi
ig/SwYDIaWGkqwJy47MUN1kdsCElnERHogdZePZ4uyoFs0tn6KQysiHJg1CpOw2D
bBJOXuXSD0qTgBItwn2Kr2VQjE3+9D3Ze7m/Uq7v86pH6q7ePUNeZ7J0dHa10psm
DhzLCXX7rKJSwCc4hoOIy+tSWbTbo+f6MFRGLvJj+tFnmWdb1A2u9vI0Hev9snJb
/RuFa/1pinOjjhoIddgDKbY25hOwyBykuxY/S5yCp+GlKFJK0rReEfIgv4oXQsmF
/3AI1JsFK8zC7IQZng3lIw==
`protect END_PROTECTED
