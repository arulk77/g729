`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
9Tw658i9G+JsF9Hcoq5LtrrlQsJ+8ZGey27jEz3Q60D4n4PmMwSXbDOwcaZ86Zxb
UgSLZTg2SEOdrINdbGjdgm5jBm/IEB2WSHS6zZ6aBCoUSGQD6IdqFBugP1n00CQH
OW0FwcGa2JrbTJeBQkcVXtoKEhPK5vb7LpAuxJd6SS6fh0cjszThf34f70peBpp4
HTtRxy5bxLJGqiMPiKlBkqpHoYloDVLSXlDmRyGgUR4m2FlJHJManWW7MWoXCAwr
eyYuoMQEtk4h3VrrAVGZQgTNwCIi2AgcCB4iXFPSygvvACCrzVZEmG7vfuyTqME0
orH3RZoWALZrscH8XxQFaGQU7VUTjR/aOUVXbtBHLBmsCwhVtMokn3bVI56lPSVu
IXHMHoM5UP8uheNMJRBo3Za1WGdw+W+Xh3wpPp7MfUWpz9rjqPBwizQ1DpNLMdjS
RYc32a3TnuaRS1UyIv4X5VznU9OmX1rNN2inVDlS8oE=
`protect END_PROTECTED
