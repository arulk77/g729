`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4x07N1Xb2ZsmJI5EzlBsR8rP8CLnc+QJgN+2M0zkyrOt
ismCmRJ/FmLlMA0r4lzE0P1xLe4hjZ2U/dp0Euyr6+j6pRlZDzpcUqGYa4C/aHy8
XcJKrO4uv0TPaE/sVzcW6XWcM+qxNFN5MkpZifmsj+Yxcv22V1oueJU4nnTTt41x
f5KawpjcdpmlGiukYlLwDylW+JpJL/gYj3bH3FVNcakWPhJ6iZqeNMgY8LFV26yM
jPNKIRLv/JX9LM0VWMdfsIaUVwW4yhCuCBSo60xNiKGWaq0KhmS6O5xUvcpPjdXF
QUTAwCHNHMNyxCcXhR8RQaDyjG3uqpcnqwURmcGxgsOTzmzTnxWpxO4ULmX/Gip9
ALuTLzcXKAXkcggr8xdNAdsd7hqAaEds8v6UKKRyummyW0Si2YFwuKLTMCPX6JuD
q+s0nhBp3+BKHxENYM5duw==
`protect END_PROTECTED
