`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1adFAf/O7/gTk7cFVeiipLjRfbPtRVn/azkz8D35bwTkx
++YYW7+dGv8n+t3JNKsikJjfizSlDxNl/SeXSZSY11BlwBMuDjzYiVrh0PfYnzsf
spN5IH4tOS+uiuI8npwG+PS0JG1OA3hWoyMa/rPjMa6P8MfZTg3U2sgVgl8YKux/
tPAyqJuwJroG3QJF2IaA0ALFTYVi+trd2B0ztHUprm1TZ+RGmeN+cSKOPM2Daort
oy5tdIvDuB1d/S7tVzn1+bEJCufDlT25kELRpbN3NRc9C3hh2Mn404bg3aj79kwA
2KztTNfdvsQAC5UiOqzdxR2SlPJgIhE4yC+KtZehTZhGFIb3nwkcIpj7D8B/OEyb
QTQ6xvfVyDhNjx9VJrBKJ1qmtITM1adc01ir/+WAU25WykfLTIObMA2BxLh/rjVN
ok9OIPp0HwvTjT92d7A5lFsNjmJ+SNbHB60H+kLNUqtNajcwyp7mO2eRmG2U+OVI
KVfsoiWD7Ic7643IrSIKohMSyBm1V64Gw0AUhZpI5Bg=
`protect END_PROTECTED
