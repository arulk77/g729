`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEA7cYUQqnHa1uONa5fRmkP99e8VOIpvqAYuvMihmA7e
DlTh6qK1sxTSae2wAdbIbDq15WCc4zQjdlqQ2HgoW1TscPpI/t3nWnOZS1d2LKgU
w5RyclDBYnqokh0JVH/U+LwZRte+w3J28ZQTw/+5wO0kcKNDx6NoDHMTKgRGBdj4
Vdu4kOjy1+d/sdbY1jaKAHIk1jCgUAHao+Xq8IvvKlYincRvNy/jJTz+H7YJZgMj
kYnjSPrXQElLVlvd5PjZ1CPg5lsK1zO4aAJcn1YNJohOEBXNIjk79SoSx4EgYNtd
w3j50J15WvKdULgiiMy/znOmAP91wmTDU+lgQsqJWFU/dGTA341r3LxI0iu02Lzc
0l0NwsnvUebZMehnXsEir9BChsTPg7yuJUKqFfJeKennLYKJpdeJ2u5qYnYIlK3K
oBO7HjPIVDQTLL+pYFTdv3e+Fd4goJu9JeEl9rGN7YDbCvfcw77/+Bi1tcTaSvyT
piddZ1E+DBF+U7yQn6a3B3JjsrSeXm5FUV+UeY8yInh9m25jkZUQsZtWVLc1u14p
ldoanq2S0uZfkahN0DEje776NEgK0OXZsk05jbTWSKZP/hRPJz2MJwXgnF62fCK3
cEYRPK4K1MeFZAQZ1eUWfEp0SlND/V104xgfA+uZ+IfDrkm9zsLkMKDmz+86wdWH
Wh5fmoPpmMQ+kaWCCMulU6yGfTS3sADIVXrsJwISI7rZcNBKaB5YYLexVdxV9yWn
EJdoi3JMtJDIWnXIKV3UNJ48Jii7ilMTvLHhAmiiPbdsq/qtmBK2KbxpGiS/TtrW
yC74oq7O12byBGWmEGtOkDoPaixvKV5G127JyV7o7KAXa9bhaOYEIBV7BRj9475s
OdDR6jH8QgGq5DEz2fESIxKzgbxR/2ryWErvT5B68aMNQIsHjSto7H+//i+ZGeBI
7rZNXjQVatvIKgArSYquEIio73iDQigJayUlYUp9pD9YPdTjm9svD4PAZqt0xpG2
WAppOmvAqsulTvhhgO4HhFzqawoHw7+WLzHvhG48oF+WTo8BgYBhT8eLbjFwwjsm
hXSHUY5VYHlKNMO4Bwof7rP8UzTNJY+8ajAR8K8DYEMxsL6ylNxwTYYQfZTdX5mC
3b0PBCQjkkyKgRBpuk6eaC4tR7t66I5lmohNRzUT142I3z1FFcJaHPxl2soji4K/
WmHM/2Voq3+Urp5235fyB1Cw0NLPS/cqxyS2bk4xQZ2i6+cmwS20A6vZ9x/3Z1tx
x4kvBnUYl8KNyk8V2BSHsSp2QFPuZRIpFSvIBBolN+MllzcAg1JEWhRLSIPs26ep
u2jvJNcg1Jqm5/qB0K4q/etB3QlYw2UBzOQ8KFU64SUwWPSjtm+LNJjX/rxB3O3m
ZI63agtI831CGyfov+M9lMV9OKjbOa3lfDugEzk0FRdrA4e1I1BgWmtziLmehe5j
aTwjN/FqFbDIwmYtWMSxgGFJfZfXad4nWwP6YyskiH/7467Aw0HWzPMm+1k6Tr26
9AM2FgcP94ZbMzKW+w/rsovc5vVHsktLl9IYbwMv9mu83Wx+XLbdVsn0VY+/laG3
s6K4LxKGdV5pkfX27v06pHSTUnd3sT2QFiFMcqQbBMoxciD5a3ayR2+n/1Dknuii
Xd7OMuBfRcUO3VdaVnPl17VKsNeYQYcJHpg6GDPznjQO/pEcT/zXAjCq0HXvd8Lc
P1btKPCUVp8/r0w8VxJkQNsGQl6nQy2MQY5lDKFXHIFXYeiZGAJL1efTbgRVEntg
QlJ7TgOMrH2oTXWF1YojDXqngq6lKgVVXkyjOZr+RCTBA3B1IDXO6PEP5Wp0pvGN
833IdcPmUhB7s9B/tggtdJpWAp/nUFAPGYCfcEC3ezscP4MY74Fz8xUp2GwIN/nV
RFnSaF0BebF/bY6WKBl3Lkp3jvYUMgHmNsbJ0V4n/SfTkJfCKgxqLjafc18s6skm
5cfMxLbuwoHSQTgbREyIOn1BLBvUp9BrfG2DEMPvKBka+SMpDZYgaS6Qs/FyHiaL
yfLCz9c1QnG5zz4BkxKJMnrIwXTY6nLG9TNt9Ikr7duTzhXn/bb90pFeAc/3aKBN
Qi0b392U/xmp2UB8JWvFJN59wcpOEcPcUhUhlq0jZT1SlBlRdT88iam0xp5ZCp2z
yGXNw0t+LOD2o+49yK/+rPAfS5f+NNyU6AaZocAbZk/03OxgquevLJzZWN0tW1Nj
mDCvAQ9FBx77EJAabcDyD724AVnyhM1NhBqtUDoxMW+a5mrt0/o/gfdylNZyeP7D
xgKkdZ/hKFisofwufxuSZcN0k6eYqUbj8ZjbG5Iiwxb7ENZayGYxncSH8wNTzWka
ql9H5lxyMWTEmhYR5edmy+6zlgXdgi9bspWQUX647+mibJX9G3q7YWHEsYxlNlZs
olw0kErQulghtasFywXX/CN3KBitYGNT3zEoJHe7c5RThefzXp/+zQIPKVpGb3AH
1sK+snx3He7H9ol4ErnP6uzk9OcL2COuWT1Di63dTlUJXGDnZmte+KRF3VbmHvMa
wi76BiO79V2fuaGyEdN2RzSG99EK9GRoEphOFgVId2zXfrxvx2hlMknA9tO7XeRm
mRhCRAC2EO06cTxCUEM55nL3Kf/1ZPmdgTrrsJXmB0Y5dQ5nP9dk+0YGsvf4mCYn
jxnR7V8ppQvP6IEWoGUyfHXUbo9N5gap60NfBh4qTTY9QXxFU6UWjoegv/ZGSvvS
5yd7s5iH0is8GyFOv928RnqFbpkAYzk0B3ndutbVq+h4kKxoodTQGw7ccEEmusI+
8aZ0w7N2pbYsHIXtoIsX3OA/7cgsXCf26SeCMd2oL+9644NODPWqzzio3vJbVz15
eWjKfYHdZdbbEvxiqNK5cGk1rRpQHmRqdQtzJU2moTm5y9jQIo2c4qcu4HFow4mL
PVR8bM8USdDksU1rzVaxcnPKuZJINDqTq1hI7jVHfZySt0d8inITij8BqKzERDop
v3C8DEFYG6CZHOV+8ltkSF4FCz5XSZnPks+uqCQ3xZEiQ9IVDHhwRwuge1VECTiy
pcGBc2LlhEXic3PqzD239tEmwrFNKk27CHubmq4A+a2qerRQ6KSkdm5VbVEJZiUu
OV+w4wjr6EuKOl1GIp4lABqH2tEW7miYH7EUiA4uNUORhNlpyV4Nt4DL+ERy8i5t
UFrmsjCUoPuX/bC6lXPS93fpJLrurLnipmaUyWNtn9m5gC6lAq82+WN198mlHiSz
dEoTTCb5wvaXZ4O5H36gskwW9fLLgwrUzHIV3gOUuvej2vwST1A0N81gDlIgmfIn
XWcgcI2yCJY7/IJIl7BzEH1WvrIgLqDrG69P4I58d3NgV0BZpOGSMXinLCIRansA
Wj3+oeqVMrK6C6MIgAFD00K0y38MLpLRlHO15Fk2QMa1iygWqC0+RC8c3d+Cn2C9
mT2TelXQ8U5uXWoSnuc/37XtpIy88sL7UdgVWt33R7SMKGH/pcF+HioCOJWkrcoe
DqVEh9z11HF60Oy6ICAUTWMU8SfWD6Z/IikYRoUJzLJqvnK2vZAJqADsKQ/GAhAK
5rWSnmWFfqYoH+1uOiNKhTFgzDc1koe7bLucarGbyDFIJeWNAWI8W+aCFI8U8TBj
dahOCjvOhRhFzSRjwGbQcrWrgAVWXsbwduDC8XEF7Wa9cIiB/jkAZ2PMipPcYPfD
6/LjZNR23/b9ahknpb0soELdZo3SLSIPJnflgHgCBKRQb59EwvzlCsjG1cVVJT4M
CjudAuQ53tx6EOqD9bUxt0cyF2ygfVAC6O3VJ5g+1ArmONfLyc2NjMYI96oXjSkZ
BpgaZa3hpQ0oQ6SVvfoXv4M9LdlgTGA4/SWvsNvt/Wu2kj/90YXYSMtTGu8691MZ
dQP0Ke326unOI9eR+Ql1oXbx3NkVDMX5MTUDs/1e/rFdKS3DGl057cXxxBM9tZrc
VWFmCd0WWUoYrHCQcvcfRlaHQi3LbTBme+Zt4JNWUYUM4OS4tU25Fe3GrPFBnVfg
vshulyuEvA4d3nMr3TnA4eqfcsYDzJDlRcdRhjxtdNn6c8U8dYJP2vTA9coL7HSg
+OipSIkJ3/aH6pyWVVp4/mUGrXxjaD5t30rpy8S/yvIYAYyh08xuuySJakn7VVcq
WEajhGS7OTV8Ob0IN0nGDbO1wI5u5J8VkKo7DCDEvqGP4KlOEiHS4eAoCB5i6OWa
tppf+lwtjW8scfpKTx8AmUqYfbjBwHdCSN6cXhCOkaB47jCg03v7XTUcQliO7CpH
3KW2DQolcR+fCDeaKKGmikIc36C9whZCEvaIWIvo+aLW/y3wF8PLKhxGYm3z1lw+
BJ8CRRcULR/1hgzJnVgPayc6aKHr/ipGlHvsaEMMowGuGefvL11E+wwf/wFhPgsr
TK8AUhWFmPcOm5OjQCacn0obUMDlwDmaN9KoN/oDBwGu59BZQPhTsgp0nG85tVYC
Jg63MXt3xSOCr8pDLYG3cI1upLXNTbQP0jcOiY8Yahe65+I1PqourztrEv4L6ENv
cQLoD/wrwoNrhiZ9TjPee2D0J8QiXUiGENkDUwarxxrulgnDfDrMQncBHiRb4SJO
cVOHtvBMjdfel4DfSrpA3aqOEm38gfn1GKPzXfieGc8v2QjMuD2zi3zxm7Dgj6ki
vrAaaDyLHscBo6CVxv9TJAmQ8oX67xeQeNy9PdJHrHdC/ej4IRYJYogSlR2GnWd/
hTDBxY9dI2pxRo7gs26WbLdQxrJF3jaK0bc0bDJEahi8w6BRjfCn1MjIwWSCJBUy
z5ObieEkixa1NkGTJgv6XsDB/zzhs5VbL1kJl+z44b3mBI3SyOVpxi2uy39pDOQc
hkTw+03FrvKHKM5dnqOCzkQgpciP8PlQ/7QSp1gl45SW7M90QcibgObkI/jOnJQN
fA+PQi/rg1EW0DYz/iHxDoW6lEg+pbnCv479hDOjsUPSaz4TcsYzU52NpBeeFhzp
NP6XIn22GTsAp+IDPruFeUQGuYwngDGAWxZVixwquiMN9LcLPXiQWvYl+DUlhn7V
kZRmdC/5t0EwVhaV/al2enDKavNLU51saDXRT7XNCipavH6pIFAwyTy4OCTQfvvg
KZqsn30iun6G5/iNC1BBBmFYhfkiByhIlsY0I1tN82dfYk8YkSxseEpqehXJ4SZa
j1N1hNwUduIcaX4ZQ6GcQloHrVRqRccU8CM9a0A2EfdF375PSgYTaHXn5dNVcizy
9su3bTYjVGhHlEXVMHCTETx0P5Ymb0AeK4Cv3ZktGtbJmuZKp4UYDQcJm8f6g3x5
R84WmvNmTxWUD52Aoh6+Kcq7aWvPGWjsOTLEqmXScZ58lcaIizNuL2yikyl1dMCF
tbp1lj1YVG5CFs2zqNhuPf3vCVdVjQEpCbHgN84tw2oxeNlXvFlW1Lp9wjEyQyjc
/vuDwHtUwYd8broDMstpqLxJ/T58RhsV+E/4FjpBAcLuWy2ZIIzLBAROW0gXyVCh
6Oy6lD3BCLMJ2SpyigFYFUW9lBFyArkg5urNw/ynhhbcz7K56OFQESJWl+ukcFY2
9s114/bI2chx5ceoKVYHnq1xlMKAZV94ToDJtPkTm/EfuYYHCIb02gZ1+dJCU9vU
VREthyUIpAzeenY7kU7BeLyuAMP+5KyPKoHvPYpKFgKDR+2m6X/FyL0u3ifcnTTK
Tp3PemYbx+ZdsidMh+ozzwLlTzIxHpmb2oaNZfGEpJMNICyVCWc6clFu6Vkx8P0C
2xh2qRZUZmtOCC2wcT6oQE3oJcdYBtMt7g2oNLMN49gmZ3CkSjhM3kUG27P5M2Hc
1eV649qsWNW6C76hnzrIvb5AE53EBzz08d+MxkxEIbg74W/oFb2MvCSgtATD4G4c
tFi7wXw3CwcGrSXVXDrASwHYOOMTaViwuEjtw9cNO1J7GVTtvYphm4ecvawrLz1i
fajLuPNqlABxJ33Gjo83Ru4Aj4UuTCZynp7wWh6MAeeO7fHLkj4Lw89bZHXtzNRl
7YKMV8wPCeiN4AMXJii46uoE05to2/E/oqXp1MIBi74J9W0VBeiMHg/TfBgVqB5L
Uku5v1OwxwdOe2FPc9PfIo6tSnPBq27xH1w3f7QNDmMntL9jxUX/FHDwbpLbXOxo
8AgQk1eEYZYg1k7lA/L3iAqz5lpb3L1rNvSFYBdX4uN2ZZIUe0042aYDiyj0txTa
CYGDluLVvumdPl8NMgZ858k1k5fzo2MxKXW3SCIwNmjIS+WJXxDy2uaQ28fZh9ll
MFGwL2x9gSpfH/GPm66+X+PRU+fKLmeAUS+Y3qp06KufZayENHoBNhB01xSG/REW
6HZuLvgKh3uvVS3fnlTb4fQBPXnytx76ikgaa5C7m/HDt0C4+bi+BJydajMthPi2
pODOJ7ffDuCf9JxkaqyluW3FN/D4c3x0p6/3e1vPYe9Y8xcsxA0fCnZd5RuadIlm
3kJTs6GlvlIPt2s7yByJ8SUeYBKISDTABo4BXontyzfrVd+/Bfs8pNVQpB5ZqvaJ
jGJ59nMvk/bZFrsddWZIFSr2z5bBj1I4Y/WEQDCsW0oT4b5C3SnEXnbgxelwl9QC
1Z4kvy5UEiHPy5n4L/sG6JRlsNSNwOUgwqqeBRCcPR/2LdBaRvyKt4B07KU+vG3u
aJ/iiCqH3WTkp4FKxomcvHfAmYwLaxNdI1S1N+NydJma5FDFVgDHITfBKWlaab5+
sZjhKnSz0OzS2rrK+N3aYCbN72fXBv9/yorJ9hx0V1iLZ1M5PgZHtFW6VsgbdhsI
hI7tPi8SBo0Ipa66QeHYc7znWdgm9qPwy15RQNRsYxXdo59nDVws5Dxxdd5ppWme
y0ydTOi3onI7pkcbk1YC35sLyqy3vl53mH5zoVKgtgSG7cmlQx4HTZ/Kr/UTRm9p
KZ6pJQRj7FyB5NxZitMDJFYuIlva877HmE6FHKz6RKYl5kh+2z2NvURav8vwP6Ds
YFY1W1Cxn51dH1UAEs/Ars3uhUHjjg1ASCMzFq01Mh92JJn9ZGZSLF2tvvV6nNTN
DGA5Q9IOVyQT7dKnt5XoowZB+CWGkJxEElzP7WL0Qgnlfb14ShYaCWdOPseS9K0z
B4ZSV75Un2DvHvbgBiriBcpzZjuQo9Ik20mibwUBIe3OAIScqvXn9NsWcv9SvID9
bdEO4fsLTdEk/uzvqgnI7lbhnyZXVFbjuff3c9Tj83J8x/DfqFpRgd8u1iIG9K4V
MhVpD5lOjl1UckCwpgWzwXxUOU9Wel9fy1t66rxi5DKcILDoRhHiyxSz2vKgeOuK
om29/1l7dna5Lu29hmzoOTBmZWhEIkeq0F9VLXL23QIAyacgO8zFKfmwlHytOt76
aJrDWV61d/+6WFJjIla5OeJC4kdVJnikr6Ll4ky0Of6If/Rwo/SAaZczRPG2Yylo
ENg9cZfm09gL7VSZhBcEwujb42codePnb79s3tDmyTkoj6J2njpdHGatAE8qgqMz
QGx+/tb7tfiTJRU4MVAmuAHxmpZBcF0tk5F9hSu51s7DTCBUAQmxkFxgeuRuAuRu
NQmEsKtRdzbu7beekgnf0xrYm4x5744ne02r1+/pNrX7fvFw2ERXlgkVa12lkpti
NWVWHepRFNp6jk7K1dAbeCXkPgU6tQojayWMh1pUJVbuXs9qKdbatEs8y68DJLbr
OwVAKJFRmK/arJq0YuGFXz6IOSvbDy48zUMER9b4hwcdKRE651waJ+cpiR0eyL1M
5M7f1qifhh/mfQadNkSw7ubcN0SvSNnXwbXhUvBdCtx1GygPwROcYQ2lEjbq9CJz
plxkbpwcj3ExQBQPZB5F6NZ+vzbd1GhT2jOejqZYBGuXrQOYiSMXhxFyHKqMOw37
EdMpLHiyEj5krR4pFVH9TyOZI75hVBXIxZflWRHoFNVntztmyltYpts0HXN4pgJJ
7KF742H0s7c5UgJc/wLJES5LWtv7BWVtfyCxxP57IGA10Xl4o7fUX8YfwmUaKNKr
3KSWGWiH7eI6AGXQ9DSvm0s36P01nPnXllmXG7PbBb5cmlsAxbG4cCOUiyF4xuIr
FVSFNUxIziDienstsx+wXKIKZG3LLN3jvbDu30gcjk1ANmqPB6OX8wlEwCLNuI4d
uV/ylGH4BV3HQyaOLVtuopeqNfqoeypYP1shKaJvtix4voB+mT3eY2nV5uD4oZS5
04eLA9NOtqJQ8ZxGCN81eubhKst0K/SokHAFnI0V+cg9KyUkvGIUYPdzZmBoWbrj
DjpuICubx/TXPxhGm+V0qFPcMgNlCgDTUeFchRf8n4pc7vUVY4ByDz9qtHvGJu2x
CZjeoCXy4On9lAS4j1n+4U0kuzBl5sWRW4CFUpeqpPVtwXAF+KjLeXhNMjhpvLwR
UvqHWW78S6OOLThDL8v5QWDE8Kjwv9CDUKVCzoXPt/NJbcWzaNzlubIqR6Gilkfh
jCStSYj6Zu7csYcGrJKXlzSXIjaHzint/D4CD+CfFekI/zPR8sK2p+Gd0ThaoFpG
UXpg+bOVZ4InZOaKJQfZnRuxIyQu9EsQoZWFrlS+1lLPdOOCIB//36UCI9k69OTU
6DMEDn4xrWMyVr42faRippBRLFqT1iVIYhejMDiY907b4wJvG99wIAlgzAunwfkn
8k8KWSwuBXYvMyl93957rgtFp6PjG+PWSbYAq5c1qYPQWl7YTygpYQbaHl8ZJdoO
kzhEE8JeI/hSCdvhQjzNsBoUw7NRejkqN19tGUOXWoGaQXp4T25deIfop7A0ZV3n
w4uD02ywQD8r4jpdkIZpCRjlmSASuJxH43coHxH90q7I2rg1eA/1RgjjrHIGwrTD
to/tCB8mSENiLtPstnSzkIZvLVgG/oMYmfoESYuFtpKbXEDxXiNnEg6Lm977PlXo
mClfHKTDI23fFrZ60GiDSHWOSzD//IvXCXfWaxqA8mkrieU7FXvCS2HpoctkvT3W
VGPIi2nKwTYbTE7xMB34HmJNQ6Ck/+9yj6KnmKBLw8ayG2QIEf0RjRSETI7JEcha
MbqL52N8xVz0/lgwtY3kw8WsEOdrcKqbHYXnjM+eBm39lbB5aKdMkOeesd4TEQ9Q
svUX0WNJBERSCEQmR4s5gGefj3NQX0dxjwr6CcmYtjHOXq1kk6tk5wRV+ogLA3iA
WyrCW2u1UyWUiQ2N0fyBdThxgKSbuor6kCzaiZPgQTK9s1jVy87mM4DQ+gu6X1cr
uKtiZjcNSDNuKVzY+71zkijxQS1+5G9aqw89j/irv1MwerJA6LPheOO/glDfbocC
Gl5XNUb0jhO/aLuDh1RXMugL1XBIewlNfVfyq9SmH4CE4n4/3fxiM9rU5ReH5aLJ
zryY0ojY8eJ/1XMRPPdltymyeSP2M8oV22RhC04APkm2APXjTuPvEuESaNVSNONJ
KzX+xDXP0FGC4nTUKyOkrBUjPPLA+tsJtA/RGp0YQxq2zgWqvJOcu+4wJd3UfQrT
8hWp6oYjXBaP0rkEul5DWXWjtZBwgwyXPAOTbQS9SaiKSvWGuri6EwHEYijEp1yj
/cGNp9WTq8YGKvo8orRl2pXyw6rO2uea5uLSmvUthl7/D+NJNd09EMGUF5Pr1bNl
XXh4zH4eOXTyaF2juMncZW/EYAv+E3+kceem/N4HUm0y6O3MKJkklLXBv2nDcu7X
2FyHnEq9ncYDjqCLFF1EvZWooVZxGk3AdnD94hFJhzb79HjttCxR4T07scAchtbl
CEJh+GkopJk7ZidhC99NoiDsPP5cJST8ECjG4kI6idaT7zCNS7OUOJt+dt0ndKRF
75D3cDEg3kqe+XcqNbzldus57bDjAyTSCCnNp19Yk7JvqmizPIVKNBfrmo0R7aoW
FPtB/oJFHmNpAQojdzI5mahmu3lPlk/VITiTeAocOeEtIG61BWD1iT/+/MP00I7P
ko/KGS0XS2vf/c0HA6ZV5OjsxFgwqrQGz2VunsA1Cacbb6nkvsJfdIV5yrwhs04d
WxbGWsBipLKDI66Yetx2jtbmOKkJXk8Y/KptV75VuVK95fa14zxc56OF/x34eXZH
jsGXy+/STfbezHoWPotwwCGlf8y7KDwUxdius691tzGBpu31bgx+YtTNTtXCT1+G
EsMyyAdgvryxKK/sUcZdEpewOdiADcygSCF3Vg64a3PK/BqeHLL3DUgI60Rw4Rd3
XmUGbPiV6WPBP/vpK8VT/DP6Fwjhw0hfo2IDv5ymCLFQw5UAGYc73p+GE9gVnal1
fFlWsop34tz/8gzpCy/OYpfu2NKgkAQ49lwXKq4GLaC2VKYJBvza0BS5pzgiF3C2
HZ7fatoFhQoBQg7Xv3cLblIAj/R9mafzmKg/fItU8SflTYwTG8WqTKuk86urcDaJ
moVeKVOlvGODE/mFUNfDDOclJcvw9Q/XKT0GohjJ7kXWornX35ykphcv8VTXWkYd
LgAw4fl56Q9LQFKLgA1wm3z47CGsQTFOV25pDQUCoaPT7ql9kwtEjSRoRtZgu0lU
jP4V692zXz9UaBQiY5tKHU8+g8UZiOdcqdnj3gMHL9cZIN+RFwTYh704t1g1QU7d
uSVVPWsBnG3jg8yrLtdZsBv9gy1fxhK1rsJ1xbwOUTnVhUCRshwDzRYIO74mP/n2
Gp0wHZWiDYcfJBUu9M26MsQG5OnDBXYFSMcr6oSwtcQnF+z4mOTPvyTsduwWJw51
5fF7etXrY2oHwzkvAjbV66N0u9Jd4A1X8X+EqqhjHdnXkzQKhFlxxnQVQee+ZdeG
YXdKQVeOmIh9ST3iiOQMsIAW9su8cabfoLP4DVkqeJaKxZ7VULmc32053K8Q51np
AHqYBpQr+YLUZjpIDF8xmNC7CWopP1aYGVrLKlP3aMFqO9NmBMdDTPqROunimwNF
GCoexVj6P3zAOqe4Uz9nZhaEEcXZsc9CCv6doV06HZNmcSH0Kv/eTkUWsv+7TCYy
4xRgeB3Xy6+D69t3XhA8G5J4/P2bK1YHNxmKvBdr654BxQaDuQ8kZv93GantzTGa
T7CzLsaLtyzj2gN3kE2+po3NgMtKFE/MO2kecBYd1Wo8toGSeXfbktH7+GXDG2pg
dwFp2eJVBP7HPWuePd0apf5NXYTslf0AkmR7rX/dxYdvcK5gMx19woiXATf68Hlc
pJpD7vxucNZ2StX4Gi587HiH1RVZ7hcR+3m1tq0Ig2aHgmi4+0Kcmvi3KDtSXJ4e
bKXM94roP+gWN62D2LJMopO2zBsgXm37q56OWCvMPW/9AQyJADAhWEqXWx2gpCrt
olbEwmIa2EMO/Da3GsJXmo5XAQqqvok58rTcBt5nwveQAUlruuTa1oeX0G8Urzdj
lnQTda9YtX0cq7cYBkSG5LiFL76WK09CUkC8O1YoOoyAAZ4305ZN6IwhaT0s3EHX
MaQFrMC9/18f78TExFrA3Ppn6PjcKLYbSI0qPVM+TuEbK649lsT4KMzJ58TPQhwW
z5TvIx7O/YJiuzR7LrrIncfGOJdme/0VVlrB1HyNyQqiWlupFTDhP2CRT57p0yY+
F2/m7g1S2/bU7OsXYdzXgju68U5BDSnyzRUoPBa8JHe11xvRqT2bnkGzvLleCh1X
cyrIoqZaZnKcrmznZ/T4Ut3tylwzjGFtrX62dNS0Gt9clbKizQDL1zLqf0DlRgCo
ifGj7MMdGKGszsHgLdmDEQ5mFQATLfwZekkKSBPgNHfVnFji7FsAzns6H4irH4US
x+cXikEA/+1YCrPqtxBeLgE5lqbCeJ/lSeDA3e5Om9LH+aVTiDZqB4UV4/4Ns/16
IgqJZQxLQtEgH6L3NC13/eTp67Tg/9PMwmkgWzFcNcNkN1GYL3Rc9pUqjKS/DGQz
P1i7uEJwc5BwtTd9yDcnKt7pfysSPWuh5JpYtM/5zyVs6re1VhF/MO3+KPlaZqcO
SkRYszMDB7KtmJz1T4n7ViYW150aeaio4npTWh7SGo+IZ7xGqcopO4PE97ghzmG6
AfPBI7qPom2xqYiH30PNA72z/cD4HImArW0Xpo2p9/gM3V1G4YL3IZMtI7Mkt+Zk
WgwV8mAPsy/Ml9JoQ//ynUAfJysMj8o5TLmwco8cG0dqIM1UjRubdDFyodRZ6jrD
0K1/kXbH4k3KKg+MSBzZksp4E2xuQDPsXIpriAgg+HjbbfuVk5hBoJIFvmMoca89
TaRLO9Ze446jIAwM3dXbBqTU+7JfNDQPcjsEjkAsJBEmDqK5jZZh2/bPmSUrBeFz
o4CV2WirWJGyTZLELIu3U1jXV9tOKRj2Aku73UyRnqNHrfETc/AHAph/RCdi+afW
0WAPruOIPkk96BT7dpUN20uacWn4zdHVrP7Ktb3KVCREC+5AU4XYS7tNzuMlvk76
d2TwdoospWy0v86dOW5nqEK7cuJV1oM+w5YOVqLfsCrkIg0qY+lDLQMoCKqd/RH+
wtbWgk5Z4RFBO6VvrSXg96zLjGaHkF394uIcEOpHze4AfGOTQoy6eUXFnJe2SIzh
a96RgjSadGKBsi3H6Se5h38Is6+FzLysk9ycCuIh3yiSgtEu5snUTKx72GVfT1GJ
SR1DVi6R4itBfz9zqgALz2EQLJwRDeYHHpFThKnFWS2y8ElNQWvttLs5hf+4AcJd
n1vP5sBOnk1tFEJGPqTNmbtq08hd+twJ6A89xBTTk6Ik83R3/GBvcxkhszTpzMIQ
q9GXmkPg01g0aFSmXvQCnAk4DPBJF88Q3ni1y0iISbk1SLJ/p0v+We0h7m4D2o2M
iGox2xsTVlMfjJEptt4f1HwgZ2GBVWVo4beetI5KoEhOrwsvpUy75fvvTOoyyWsG
VbvRuFMzJ/NtMhYAp7ytdQ9PYuLjZphqldynfmOEgZ4XM+KpK6xdHXWnqi+SeA2Z
IIF64msVCH2doQ1KqsxIZVelzgTQ7WGK601jSrfTLMybAYKbHJL5QZMh3BZZqSVZ
+lLUjyyxohEowkdY1c6yN9Xdn+O0pQIHDbVM9+Hq8xWBbkoplOorRSbPeGqs7Eew
0e0L9VFU2f0/mwdlAyZnTbZA+TNJZsZ9mN9zjq/ecHcSuOLxv/ZGzXCOAz7nfp50
rkgQPwy165ksZk5Zbc3gYe/lGX0kT/31bXg9s5327UeogZB1KRP6PHtweSYje17R
e02Vax3mqUt+Iqr4A5I2i/K9uPDo5IDO7cHaEVidNVpzL0j5XSrXizEhMWagZfDA
9O3cB80qqU1WNPOFXoGGVGQvzEIlSaCL6k6IluDOJ+pKBPzJ78QcYeuK/luh23GA
iB3mkP3kEZ5wxNuO4czF7nP14owo/vOgf9CGNSzOJhraG6UsOzUudD6qL8uZm2ZE
YrMq1KsTwr4X4s1H5STaKrw+fiQilsqLfX/hJxwPDZryicI7dyH8W8lPCh65HfMQ
1dqfBSZDKBTM5szncsMnm7vOr1ocG+/QAP4j18+O/j6PFkmIJFwBKx7eYN7U47rP
rySGbIzdvkxyTGOiFPTLYLk7HZc6NOmhtXmlHhLETNeNuFj+BcdIlqFhqb21lv5e
m9uBmily4aDoMt1RxaLgSluJfGJJw5sjpyJIJEM4DKs/4eLcbXfQKPJ2/CQIv3Ek
XwMJrjhSH5OLJf87zE2dxVO3LMmb4GJyF3mKf/4JHNZIJxhyDVxLLEjgsgcQnHf8
9gwD13MfoCZNIMFohxsir4yDGYixEuVAtFr+7hFJw53ne6vkHEF2qo6pFwwDzVX2
WHot80PKOtbUloRjoCrI+d1oObuT4g+A9y/Me06gFUuNWyz8yIzPuh4bDb7n43id
B1+ZTeDB6ed0SFGz/InC8an/LWBL2syHwUsKjTu3cBZJHn15s9faE0R1A8uz5/JN
UwTJYT3QrVh8EC0LsJG+UYkybPSbzse+f/Cy8+7zHli0oehtjtJ8J1xgRzmWme9b
JHDz3TVDloXBRTC+o0R9zxQO7aTHk7TF/q+e6ECnL4YRZ96zcihOsgU47aVvGHab
fXladndA3Oo4yb3xy0jMP6m06aUHy3ByIaG+xjHLXq9tWBOk9RjHnepHFIj/XNwE
YtyfeccQoCVBhDsx2hjGYzsRnZKL5rOQIzo6UHKddG/f1v14eJnq70YQcPwFMfwO
9tJ9vunE1X+/LGdcKqmzezwRR3KsJ0LCCOaXSuoBeaedbDFG9iRmNKTXwWHyViCs
/eOi2DC1K9WGqKdCpQUwhxQ/eknVHL4toNJrTPPIwZAZxqHUQbLt3TnOfoHjb++C
U5eye0ZiriZJug9TxcXQLEzFh3A6B7dv247ZfJsSiRfBFio4G/PHFeUuCTbyBbPT
vJnpMaFWvTXh+DMTULWH0sSxSJfn/KzO6pw2ub5eD0TCDVJhrP+G02sk0TYgL09t
VsZ/ruTw4hzFgdrLWt2SmM2S21sndWHBTfknPNkvd0Ls+u3a9Vc0FwgAcIloU1VD
`protect END_PROTECTED
