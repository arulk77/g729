`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C6iexkR6ixFlWqTdiMY8N/5oxR5CFNi2do+MXxznhrEC
Np76lg/V3QuT+HV7LeE/U0Qk+3O+1Ciw/WyekQkwLwlSm2skr/3a9aZzW+eyUAeN
5su1Qkhdb2L7DoN0CGOmFMmApNPpgoMTfTzuW/7M0+CzJKWP8HQ9OkZUm9JHpTVD
VTuoRjGfrU8L7KsC7hbL93FJqUh0rcnoPuuUFaYv6jsVEGZpCgvZwqzKtTl317N0
oScDpNUS/7ChopczrWNz6dERKhNH1XFGN+5Mkgvmeq49gXt0I/1xWDz923uppyN5
J51NtcQOXF7GSmJhlIcTb7B9tcJJfJpTZ5tm6o6bCbylRegdkZNiipFSKUhd2MHf
pn+SFytTBaMnuGy/Dr7e4cnIb/kUCke4CiY1AgEA9p7gLifpbdGISs9HHyNtvLML
8oJvr7vBi0jy2kF7Y8oonFD1rWQSGTWIiLSozrf3NzrklJ2pSJgbW6rg+33q5ljv
B/GFFUkcplhLkrXsSVqdopzvoiPZjhNEdi5f0u+S2pDs3BBoqLQY/ES0pDZCB40i
dA/cbySPAF2sG7T4+uD+qmRdkwb23S0PHYTObr54nQrwz45zSYHQGuqq4Xiu4M98
t4zqh8zQ3mCdfyXL6mcHaIAjw4BsM7LGja/dh/aXvrtKNk/P1eZI9kiou1ERzblH
VN6DfXaQoeQidwkA91rRHGAaDMDDG1HbfChrd2JCMqeCMeH6HTc5V+xUzPTp26wr
HLQVcQ7ipWxsRd8HlmbTGIVeeDzTHWb5nfUShI0XYJTYt0eUIzX3VQDhF612mz9F
9HoHKr3kw8keCUHVj41lWitbXob8ekWXKM2DKcRKqTFj7NIR/NktxAKNJ7ig3p2E
cJD+1XcjPAQ2P3v931iC8ldm+tEkj7Lni6QgHddzt3OranMwtgaicE8FkbpkeRaR
7To0ktaTJebFupgb5IhBQzZvbTYUAQKnNj5Vy3J+DW7eCZ6i4Xm0HmZBlc7hsGcl
RM0RHm0fhUHoM8dPrybP2A3g19MJDnKycQEvq3lvZEdh92foaxLGSh+NGLM9LGAD
5ciS7uXgLVZDxjNI6ZLUhD/wQLi+M6RA2vb5rh489XqD8PTFUf0VyTLvB8SHlITL
jVtYGiA3KTAfsO2jRzFUQMuqxKe17woF1ukMeLAlve3uzCy1ZS8koeeFF+CJAjYR
S+nl+a7o3qAiftpIn5Y7SBjrLDR9TI4DYprWqyZVopS7qpDIgOo4UZtfkLBEv624
Y5MHKNzkjE3Q0hRQMEaX5B1THhIbKzxljXqkM/aFzMig6yPz3XNb5+t0sj14Wv87
6VVqwKomV81UrcRAT81pcQPb2X3wUY8txb4cuERX5gD/ZZSEKgEYtWVg5y3KX6DD
2K5ajpAP+E389XWJBpmH2III4juzN6oLJrp9qIBge8dhvDcsf0UJiUp6rIc5azUI
5obx5fMh2njweGzcxSG+jX0YEqiOAKqtUTMD0cCs6XK8JMNYfoKQ4MsSgxHaJZ9k
qEVvd8C9RRl70iOUch0mqJmtR/wnPKN/LOwGs7UPMbzpQ3ZwZz0b08465C8/lIKH
XjJ+ad6yYK4hePPztNiX7OqAHRW0BUYupH6tpDwHV/PTT7iHJwgbfbvrw7eMxc38
g3VScXi+xvP50AzvjlBuPld/J+B5cPDOp7A9TMe7TahB5dNFLUQRwiuAtZHCi9o1
690ktH8i73h/mDEBc6uQ/w==
`protect END_PROTECTED
