`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C34GfcShWSuhR5T92e+3JUHLOl27ANRaT0m0kdVlR2Lo
mOIxtpPINntSBcatvLTqFZgtY9OSrqG6yWsOx1f3FmDwMdOxFTeRuSyxhbbBhwy2
FdSTbSWQgOOkY0zaxPXVbNCTsC/T8IRVOO0egJfS0zpT9B6RANf8fTv1Q5Q8cPOn
h81ZddSJQhfciq4CyIGdgQ4c77jHbV4ECHAhdwFUrqphIo9ZPhSakBmaOk2dF/dd
97nPuT+4qOETF5KJcQSoBVfm8xvbqpk6vLwPszJZ2pi0P3L9Px2MAGOgyZADmEMS
JpAqY1kz/uyh8uy+L1J4iEV3ckdtpDJf7/f2ULHTwXJ7pCgj+Fxj6tkK3mvbBCSS
M+VoJ9KaE3zqOkpnuUfa1dXpF4J6wMm62Fe1O5gfDxOrSpNVWAzrUaaGA1uk2kW8
w2cgYcrFN0JJdnURZj3dcAJnepI3iE9uw6bEYrksYB+p/q25I+eLussUe0o248sH
DNOEZNDDANaRnGSZNAq5r/nXdW8PnP+LK18inbjKMEQL5NDtt9YYzauDKH00aNqG
ej2rSUHcrC4YVRLcxNWYh6mqbuwXsWvVREaXfP3Jg62J07GalTxsyNOaplSIQLt2
ldbLXSWwZ2QW1hYMKuBMfls5A3+geIQPJ2X0MnH5/Cd3deren8clJx+ZMKBhC8Tg
XbvEaTANpFwwHdfDtu0907OEqbBVYRz7Ublq7K/iw+idpjgA+xpyH2nqrq+oPV/4
7Ckcuqsrbo66cSdMDtcBJeK9NvRen7T6jARkGBkuUGJyfUEe8ig8EF+OF5QfZjJL
4oxj+CgsIXJJRUD7mC691oBH9+AaAlFfQ6aqVkTxOpa8AyFzFP51obSie9e2TQZu
5mYUnbbTL6r0N1JO9gcyxO7PCcmTeqQwrAn/QbOgyfUuparwyL2iCZZoAvoK6KCL
jWYVua7jsKtKQHB20rohjdWJAcroLO2EG5vBzQOg7Dj0uMq7fMyMuP/THvad7fkV
nTGvP1nemjiFLzPfjXom18JCHc9/gZn3RYgmSwVBA8LIZD7JFQdlqXvJH0EjGAKo
SslpLwydMVLQzpo8uX4njAsgJLaitpy7KbKs/97IW3s=
`protect END_PROTECTED
