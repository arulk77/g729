`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMOB3RIbc41Oz/QsnX72m4jh3kLOESzFXURqcVmOXO6x
79PXMmpBJBRe+GV2E+ftrGNUEwNqZUl5Nc2rB2v+vAscJ6d5lTOgFTAbEs0oCEuU
S2TjcytW5X4jhODePtrWfhVSTJPyxjsleHcK2pn8XgC2rDuG91kB6RsAkKngyzzp
uA5xAY9UAPYFTE+HuVA4FYmRTmymUEUVKp1QstL4aioQWejVnm6+inJHZ/d+KYfW
eYYxhYUtlJrpO52z3x7jJtR/Ga465ZYO2ZdhN/ZzEtAHONrYwzSL5eYDm9Y9rM1r
i3B7c3hWbzzh1NANjUPv/A7fbFaQnwnKtNB+RyjP4a+FgOZqST/Nff2g2goTe3Cl
bmrBd/Z21c5pswP/KF8p/P47NzTDhgVGZVcbjVV0bHNohnvMLwq2bENW+dCu92CD
iygM1LYBTl7o5ExCqQWwD350hwruG6FMx5uETPNvNq6DeWoYxzyQRCBohvtj9GR+
`protect END_PROTECTED
