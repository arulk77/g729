`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4jUYkdt5VjR8oFbu7ZiLksxjwJ38HHIpknM26CkPJSGjtUaJeLX9yZAIk2cfyf1X
WxxBMLIID+7pF+93x8Ha0KJzpxKhO9TSpv/r3STmBSV3gf32s9ONF16fg2dPgRPV
/YIzRfSMwdwPexa/XDcB96WUuvjoIcYXHQI7Hw7zKTNaKBQytrhYY4JJfoRDGzez
QaQQbed1z1Toim+kkFA605Bxw69pdYjKbirUcQ21Mi+MBNI31KzSWYu/mOnaC9+E
H147RSOIswJLuc3rqXylhhf72pqMmyB1Elp21pdbm/1Vo2dygiWz65wa9A4Ss07r
`protect END_PROTECTED
