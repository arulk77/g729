`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
GykkTGYinxNegGztgRAJZUBDwq87lLV/Xjl6UjZ7TDpAEpADS6WW185JErvJaaio
MLNp/u9gcxg2Pj6a8RnBcKKnx24Lk9cn2KyYukikF5k+Ni65ieri6GWBHzEsVAi1
9ADkfe5zV49yac05M3QBXPngsEw0pJSqqiKlj9nHCzI=
`protect END_PROTECTED
