`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
eRGVbKx/1l8Xu897I1nTqbbmtBcLGfFc92LmdONl2rJhnr2lVxO4M48LIgNogvH1
VMIk5f1aCk7bHWbpxOslDe8YVbbf5qJ8rEZOx7sdD5LOfnSeBKsiZ56N6IncXJkD
ztLfps+3xiohkCi3lujVQ4iFIvo3ZI5tKNcDoPUY1M5r+AA+SMRQG2orASpfK3fq
0DdIEsDZ0kSQxec5lFQjHJiDqZeZ5Ic30ZGQdg1r6mbyytGn3hygO9VOKHDDRLmX
zoSPUZKoEZ6qxUc8DJ62kxTCN0VqMnFUNgflaDek9DW2h5zaqVwR5zAlSuTF5zc3
YQVWkhreTGhBspEtnGyLNC8v8lW5FGz5vjuxBF/Ny9zRXD8bs57X//CEu0VYn6he
3YzLDEGAdu8MkW8XDvelqe7Tifk0ESrIOUIhpdoX/Fk=
`protect END_PROTECTED
