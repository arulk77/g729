`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDQentok5Mypqmc5z6WaIlEMpFd9Y+IQnl4nryIAKAbo
mJftn4A0RZEDwMcaS+1S8Tg03dRgjDrW/FipseVy4gGiNiJNVLApK3u7wkH98LDA
njZqOSnrMixJIXmeU56KqmQz2QEbo9eR2y8ewX4U/Hfra6vwYLeFvJoM5b4Wbrwr
U0htPNQnXndekKpjKomYaqj+7u+Jh3gqcc+I8hmia67qgFBMjEPpg85/Fl4xND0X
`protect END_PROTECTED
