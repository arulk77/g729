`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBfXjUIVb3yWPb9vRE5ziBJeidyjfKFx7O8TEjaucddL
vCfhwW4XmHVotdK60oFQWsB8tALt69YpQaN3Dk8op3d3gjfV45aAJt2YLo6zbXAf
WsoqAUxj+3RYZmFIUCd2fMk8DwaOHxWBKSNSPhhci3/hGySKN59rw51kXRIRtIgH
GVkFbmw0e2OD/aYM9fdW+MLG5+4xaAcfkFz1nxPlRng=
`protect END_PROTECTED
