`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xt6+BQbKzcKR7YFKgnuxhvplh4k24qeeCVL5GoFUWt9
2OTbDZ9UIhE4r62SR9GzH6wrgaE6rVd/bt9Dp8IPiQdyJjFSd08YuLkAhgPG8+17
hlgp69a4YF+XcfXZ4bMwrmMUBRrwz71QgCsVfAgLvkwYUih3xoS/7MWc4o9LmiKU
XCoG08y920jdjpddFIQ2md+q0wVU4jBUfrF9C/XD59xLKtSC3bFJYALMT2HWcPla
zeeUujgeGtMMqRQiHNxtBBMxdwUk0FwQZFtWAiBn1NBKunNSDr+4nHPVuoud60UX
pAMetZurJz/g0YEqpfqLww==
`protect END_PROTECTED
