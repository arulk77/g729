`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCers+tcyvO0Na3IOlOqsk8Ug414Im+hxLLA0ejqXkVi
Kghnx1rtl4c3FuG5A7wioql+qosL7DGP2xUM2iXs3edXU2LYJT5aHTAXr2mZIgCT
aLS+M8j779ekXKxbAOdumJeQH25eFinRxWAZxclS3BUjvkTYD4Dby76tksfTnZWr
Fea4ZHthAFAY6+ad+JdvwgdKU5wGJyTXyN7ucJrmnuefkMaqBMdnmx3OSBJdsWfN
am1nX+F3HcBoB5hcoWzzSL2AMGh+Us1rtiAH7SPGDqJmpUJo5fnZGWyWQ+CSHerF
QYCYa0oFGz0L/mG4vgz+IJN25KmmsEHlEMu5aZYstiZsV/Fbz4BLHmVh243CQnis
qUt4Y2JPhWTLKNVix1LRI2lwuQCn3CtO2FlqzuruW4orkvL3KtSnqgbLaAdvNnyY
bVu5mvWoW6/NXw0vwI5d+vIkBk1P6TyNU/AdQJn634YTvDlFgi0XGAc3GFhO+p4u
Gzpi0pdk85r9qdTNLyRdS1JahEifVUdbJsvj7XVG/30o5fpL1UvTfaLfjYNS4FHA
EwICllVZAsV7U4A/uQuwTwZIYSUDaN8xvBoEiIBX+fnsdGEzZMpYrnqoTXv/YPcM
`protect END_PROTECTED
