`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCBVW+/edclGeiWyR0u4sn2HTqe/riK6hkkALdTMVxW7
6SHDDtlGbw1GQzN+rw7+5Bhv0TLL3r8aeIPAeyJBljkr6SpTys/52zLOYCv9pDyT
ofZVclYIgwQv4iglvuXUM8y7PWPBDbgnntAdxsBveIYFjH5cFYbNKWNvz1JYjdQW
m0XwJN8DbQXrfaJq98vvP9E5bKiNtnoJoeHEjfvtPDw2IfiZl9Xis9TjG2uBJLLI
43VGnjA/rWLDGMcOnLs0iK05PQeDMzNutwRMgqekjAhzHJm+P4dEE+w46x7LdIGv
qYV8zAcnJ+uZyIugFCNHSJDPLBQob3XBt4ZA8XNLwdgZOLt3f6ie1rq1+SANc9ZL
X46GjPgGI8gW8xTWUFJS5Wwg3Y8RdurqV8cnDegWspZdlBS0G2HU86YTpr2Qf+fH
6w2LTcxDWBc7Ufygz/hCUaUuHA1MIws51wMbVw226X5Z2QK15eOvW465Th9OWEGB
GaikC8o1WnMOb2HdWydAt5c2wpfzyeLRHuA3xcBg/ypN3WGr2YXnBl+YtFFdi2VX
`protect END_PROTECTED
