`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDARtCBiODgIFAUdF5C3P2wGwxk1mgFdmvj9KiMTw0YnCE
lAGQBkGh6wUuTfq6rrb1QPIo7YUN5pbWg7KkE1v4m9ViUai8bR8/XQoDe9iNU/k8
j5vsrINU0bo3luz7uBLLjxovejGprTPctRo8DeTEy3KD9gv75lN0M09kYdlW7wFG
FmwNj6yoa95JSy1dKUZbt5hy90Y5jLYD2eucE7EHOEEpTA59QHTGE3703YXvZUrc
T5Q4/P0Uz9rKV8SHYV/lVFiTllcixZHkqLFbdiAovReZFE2Zi3k6Kf0lKKZP1O/Q
`protect END_PROTECTED
