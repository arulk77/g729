`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aRUiZobP/7G3IQZAv/qr4Gf+sV80zDMtmV0KIZa1gSOo
WxwhwBe2AKEInj3fjBSZEph6mGzi5+MhrWN4jvmx2WxL/kmNojUpOxnEfQJuTLlH
h0gfVBWg9kA1lSqmG88RcV5hu5jEjX91oPA1DIPP/148xcEylM2HQ5WjyBMEFb+y
OhzvYdGsHWJVyvh1864XhHO/qN2wqDlukm/9C6v0qfQmssA3Hn8HIgZgREMp5fKC
3LTgiPlDmuRsgpQc7GQLtPSFPrhbpn9CGupNFPES0A4478u3Tfsqhdd18KN2Ae4n
LJ0hbtm6Ym1GYY/TsLEnDl9cuDbwcl3cah847Cl3850sOHcazYmTT0ZAw7KQWWBd
BY5/95c6EJBusvffh8qoqvtqvW/qTAUcSNRvd7XjZg6KURUB3P/kFyUI0Apr/xnV
25L6/UD6c2176G6vEPT+W6lOZXcjJtgNhrPx1BFN1AwoWEQTggMJ4VBQAg7duybi
z6p7BllM0f9R/dUBgiyGfpuWPKkhDo+7wJvutTdRc3+GX9eOE0C5JMGtZHyyKlds
EFb6msQzsuQGDelHRGi1VLozW7cA8aGwAPEwkNt95nkRvmCzCC1j1m2Ollybe4op
1cCzCpr1fBW+5IIVs7+mgt2hDFjy5lW9vXSctOruigBDf4xGHyp9/XNGIrjiJvk/
HwfB/33TZz/CwoagPV3M2ZN5rS/ZgjO6VHdlgZ20a1N6HL3B1ohGvguuxRLjWhGK
VDmrs24wI18Jw2YOp3UKq3jhiq9pHOqpwK4OcHWipUbtGCuFHbselO80nBTw+at7
v2yIoscc832b9f586ugnT6UnlCQxQbxayXwghHKcOjJVV4kOZ1E8/khPB7ljHiXf
LO653MjOyXwAvKMUOJtcaDtSrjqYpwm/+XQy5Ey+It54YvLvaxGjEda9q5daIPdJ
owPao6X8UsI+D6TIEawaV2nRWxjsmnrU5VLxJZZcCqxLGKvwIwevhFt0c80phNJD
kK0lK6khlonY4T69kPzQ27HfqxGfby3BKsRFwi8XoO/cOSijlO0afQCrHIwrtbTg
QNmdEl7jmot0hofjSlVsCUJlVN4MyJK7N5huaUSNp8cjGp58oIk7w+4lVsBRKz1y
qDo0kzcQSzrLxmQWpKHMFvXuFcdurj5GLwDxReOal52YVwa7TgD5YqPEaMCuT7CT
P9l2FDDTe6lg4AgNgxtkhxI00rgnlXEdZQvy6EmiFK68UkOWHv3V/A8js85H6S8m
6Tdgo6g0+h/HzPf1S3vYJdfg0l8qR2thvrA+bRX/3pTWMubajn6qF9ESz7e9D8P/
ZVUh+91dMu57/Qaqw7hr8rMWSIJI/Y9HV/zdyUu5rCbdjkF3yQpEdH/dlHQ0CiX5
akqFkAYuSPBou8QoCsU/kY4noZu3qerqbjskLrdgdOeG0nY/mJGDhduZ6eNf932d
BmHnhykp1nM/TdvDn3QruachDimN79DwYUKOCZ58UNXH5n1NvgBlYsXjdSXDxK1J
GAHv57eTpWj7qTGEEwoAI9VE8LchQKSii6YIHL+yQmRAk03kRGWY4wwD2CZkQ4Ax
yET2ibLJtkr18UpJh7+0s4ypLiAUfSFueWtsiTukrT7xQqdWaGyl0wI6tXZQ+rG6
FD8Fuk1YOZmeUGEdJmgexrm+vasgs+QISzWZZAay+rzo2KTTOoiuSB7+wBC81lyS
6xZgDlFF6aTma/IHsk7sb9oavej99hTK0OqG+OagJ+W9Wjdlss0DJKRtaqcxOsEi
BTxeSLActal/o2rEYX4E1A0FvZQYup/jqKivxqfdNBWkNDmJkvUOuHjjb9++nHGA
/IItKGDOe4uKQ4eH+54VgQWBNLMXePR3iV6iv/0RF1Uq/mY7X+Z6vdgfDL0n93yI
ThEsCFuoAYIAYVQeOv4pINHk5u01H6cedxe5g3hPwNI=
`protect END_PROTECTED
