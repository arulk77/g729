`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SX9dbmSz8G2+XUKgC8zcRiBdR7PBL76LbNH6t+fS31cW
/Jr4HtvkpMZ5Ggzygg7vmQwmavO/VgmWMKXGsmX/dZzh0mjCc2Kx5XV91ykE7Zuu
OHI+AS88xXmSIbM4Rri/psv0/3H4R+hmaIxli4BYMRFlDRVmTKEVNL5gePHRoPoQ
5soRjaTBDCLqydqCcEpQYQ7wyW+phR0xRC7S6XJCxes26eTFCQ8v4UhNtXIOBiIL
VBo2bv+7JGA7VsVqM4m3PcNnEmEErFqtavMqFZ2lBJ2NorbhFNgis8mGEiArUzEr
UnAt48XHltdcXOCW8uP2MSjFyncu57uAXTwn2vIK6094066DHGYsn4EdGGLv0iaA
TMGJiKYx5/DwN5F98QHwytd1x6MlZlgw42DTeZsOKrXo154YH9+N9QRIFKUqtNGz
Ia95kLDmdK4m21Y58SSBMgFe9JrvnjruF5piRuk2qHV2Vi3C4COq/CuAeZkJ2V+q
yQCTAQJWKD+KUUlCnGJILbs6/IUyBqV37nalbGFFHIwd6FEKsw3uqngtgZ4WgfQR
xUjuCAtUl/upF99WympvndczKN6owh3EXWKe7aJYXTrJrTZw5VCRVmKGM6TK3Jim
LEKHBZ5FKGH2Jld9eyTvrZmanPkkt7Vxh3aOemTMM3zy702oDoaV1EQNcj/HGVqm
CEzZdJZN22dCslnXdAJRXMrT+LzygnseYtohJqUk36iHc3uuAawu1opR5y4CJQam
4NrYyyKMcjEsHs9GVK7bTquz2MnI5EZny1cxPNLeo0IdkJd8KRMbbp0ePwkSJd/A
Vt4UdUovCZSWwoSRdCW0S1Cx+NsWlsAd0t1tzf2wuSYck43ZC7ebsWgTivUieyHz
JVq17SNrLMUFQ2F2u68GTqvw9F1NRGcwi2gM9JaVuluqMcN3Oy92c0ok4xI3iTmu
l/ZraIsokWN1tId0or62vT4eftQpeXVgZ90EYcDKTINQmsnjxKmVCttsZKxD0v6a
YkglPf5Vs2bRpwKJsbRvwnJGaAB8KEAOY61BLxETNSgkr1yaJBcWUpKxTKbapeWB
UqHDwrf1bAYLjpCYWkcsDmG8ml7pyfT7vCtOitlJb873caTpZAOcCu14NpAmHyPm
Pv9s0/1gZpcxfGY2VlPnad4uV/uqbLAOTsaxMyz0RbxoBhBJ6fbAGGHk/kfl6RPV
Nbj+dBf0gcdY3gDpeJRXNBBTUBchkdZO5CnxbMc0zBTQd8xHBF6F6IEsVBmneyAw
oX4qIIMNYtEXxQ0F3BGCJ44FaNAwtMdSdaA2EVFaJXg4hL1NOFNTjy7bbn2pGaTp
9Tf90Ga0EeEX0P2wYAPYczzpA21j0be+kfE2R4P4sHa6BapsC0jb6dlbkR2p7fUi
+mvKBukTn3jVhbtwj8K6mHQi54ReXI4SQvfc3RH4/Uo5E1nJI6oKWVh+T42Drm71
DAeV/fqZZQD+fkJ7XlfqB+jucP7MOkIzG5rALpE2Qbqw7XwC+mTuJkcOeg0khQSR
y5OY83ri/OUxNtdkd53Gaxs+ACbAutWJYh4x2bgB56qPVzY5MzgnowOlsJ6Q5xNM
tdRrkdH2WGtu2SkrEY2gsxnOK4pvSAiC6do1m4+N3Df3+BETVaMJucGjxV+vD/0X
DD/BCQDBi7DrC3n8S+HHKMv4OmTBNm+e5zzAc/NRNt2wgB+D3JJ1rGPnV7ZuX0fN
91qCwpDNZpx8HlvDbSxV8S1tIB318hYLu3VUoomgdECaTvq9v19zahFR809rjM5Y
A1ftw4WWW6JKASLq1polrCrGpYDghpFrxfQqNM/sSFpJmf158u9lSLUSkdsmPnYd
T6qAjdB1E26LfWA8cEBIs/uZK3ua/iq2pHIEkBuk/6KGBFBxSp65G9cXlIaVikxn
LNQYXztGN6Wz5Toqp77Jz3vfjxT8qL/feyRUTyiVj5hmz1F7cXmwFWaHSWBFkI3K
udDsUvASYAOkvo8FYc24n4eFGSOjeHR6f8CRFy3poB3Y4PFFm3diW0RFhtU+Z29w
plgrZSg1bPAY1g+oagvbA2Mx6AO5AnzaqKXnK3bLq4XcOfVgftHr6ebGKa62G6He
bVs3T8xMuHqGvojFVCd7pI51CAanv3jSrEz9dqlDzVQqtfmd9zWatKvTxHCbfeuz
7lVLPH5fJlE6S3cytJ0fjw==
`protect END_PROTECTED
