`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ2ozqHwy3cADdVQXYJkLiZ2A/iCo6ptnthKJhEied1+
RnY0XpkqPa7Npy5tG7COA4m6sT4nV9caHM2FpZ/LI/jy3HJ97m4ADEesdHVPTHTu
7S1yYE5UOSbFfJLsH0NNP5hLs1eVg8wLSCTT7cgGnLI+f7T/eE7aCvfK2RNgfquX
V986jAZuhVHxJehklBtAGg==
`protect END_PROTECTED
