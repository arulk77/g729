`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePcdqWx7ITs+ZVfafxYhaTAAjgP7ZSQUWHzGJ1/M64E5
bPJ8ONtbSaJY0+T0+/0xbmBkmHZXGjR5jq1e8fSN1CkcVsuAkuItBypp3fz33lib
kGXJ3VDyt8+KaPKjdZ/Ui1fOFbr6uV5rJhIfIQQXSgXO8xSi+O/vwhe4/Osg4pzY
A1I6dnmj9Czf+xG3TF4xSpcwJaYrnFM5R1FQZ9H9734x0VNUrO0rzAmODzuEfF3d
O22ClCNXXdFMpOqlco8dM6U1YKgkZwcBjLvWFWRl+zaEm8IL9ggQ7i8Dg4OuRDaE
LgDn5RD9UJae1R9WTRcWuJSiq7KAqvy3YkRfJINZ/WShUWMHTBRwgCUlIL2KgncM
D6UisZ3/OKGe2Th1csJLNPsAilIj2dedP+4Iss3ru6p5zVLcS7rbfJx38Stu7C6a
LnYMAbZQbhBbMnqa2qZ6q5o4UT5b9CfYMF6YPp7K6dU=
`protect END_PROTECTED
