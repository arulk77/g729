`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
l3sBjIVvTXBd93KCjhg5MQRvaq5fK2JhlNwhSwH9mxHEtwHy1qqxsQZd0Jp02OL3
sfo/MUXBAHfe/aa9Ge9jXWhZI5jeDF2ZbLfpoEZ8AvlUAaYJ2bCX77fsX3pj4GVt
uYFkO+x87Ef0OlymA/m5kEQUbqj/qtPxeabrEMuqTHjEdCt0VVqRqAsakd5U3tQV
eLHAL4WYMmE04eB1+YrHlqqjMGvcboQACu4GO/i6v+o+nXd9SCvXpXodh5/tkYcz
2j5wEFEUz/s56LdsAwe+ch01uK8xsaJgMY8LVG4LJ4MMx5AGEZsZPLTmhMpGhiV0
ylfW/Q1SusVklB/Q63fKs8JALTqeh2yPQks1cnFlCTIGl2jACuHEHN54ud6n95s+
OtnoMp0qL/nxf8WCLQR74i7DLeio7xZ+78j3pkW9tRc=
`protect END_PROTECTED
