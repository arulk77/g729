`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ya5oxmauLPBhNeyevCkYV4yDdyP8nuofduJDIzEBjQ4u64ZArcbd2isnn57WFifU
V8cM0bPx4YIO52E688QMNUvj4oj9X0gp/ckjpk4VFKQxr7Ju7WC+fcRBqJCIzTpg
p7DXsv6cMCevDdHEiu3iRmO1ypoeWrZK+Bfwqr/lC4o=
`protect END_PROTECTED
