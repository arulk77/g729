`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIHtdrlJe3GIjojQ6HWtV4CXKXkmw1cQ3RtnFLJYh5T1
WodKys+noP9ESrIn6FPj4jK0g6RBjObbWtcpuAqd+6oc8V5hEpsDYttWBQEUHXsW
96QgVEGfWeS+XtxO7UQfr/TFFLAp/+7k7GSNgWf3PxgSAYMkyGbm3Sj7dRgZN6Ge
eL0nJsU8JTkSfkMYovwlauGgaxSPjDAoDXhRQOGz7U44asHQhLzkYM4Il7ySJnY/
QuAjEApUyvv/CljuWfxTdb4MT4H/9rfg6cxPouAHx0MESoikLWHRyb/+iRhi/Lvs
Y2VjNZsB5euMq8R8fcqEYjnEjGmehmFWOquZoK2ZcLAiea1r3+85VsIFtPeAeNcO
jSgePmBwA3VMfHm7i1/MLzyd06/TrmDw1dlHTPfTN9FrhLHWgaUl4DQY75wehyLs
XqGWogU9X0SnzLtLgCFh2lHhTgeqxHn0GvYdk3JnPS/4phSk0LQB/R147gmCNWjR
JTjktSfjqhfrfc/uVok0jq4wtwX/VO2MYYxCSL6YmcseOmCxLPR05HjcWEAMRGN7
M4I+MZwRiBICXxsG/pHgAl5nLfZj+79hNh0VOgwM8Gs=
`protect END_PROTECTED
