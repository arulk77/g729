`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47rVQSyb/flA5LV6PrEyspzzKoAUXN7+GHaa/o+BHrSy
3MISrMV3cRF0Lk1eHWWXNLcowzLDX6qLeT6nTiMoW42GFvfq37Cd04aPeiZrxAQk
Zl2C/ipwZR64Fcnpednm3xNuzYiE6Kg3TwrAW18ZCskK5R8qboRoliS+7Hr3ogA3
VOGI8FXkHF5yhheJfBPQESPKIGkQOeuSu7UYAo+XZBClFycvqrZVWxnLHWjgMKjd
KxNQhwcR2XEcjgV7hXlzqEXWWyfl5c6mMJKpFIbKk1JcnsLeXZeLYbr8td1AHUlK
l6wgMhUhHVh/a3GiPpukOw==
`protect END_PROTECTED
