`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
M7DbFerZNIZiKQJxp7SY0fRK4HoOiBhw/jsAwOltdfzGzpEGXE8hyyCgM+nYQZRF
Cn19EKkeRy7fnZcuROWKLv/j0oHBSz9bWR0VQLD+ormJduagd9qnjRMH52QMQvKM
AJIETjQkZ0kgtBIOF9tT9pofnG+gfmv2jBL5Oq5gfQOOLbdZw7GkORawx6g9c62S
Kgm5607jLFXJXnCCy/kZtVwA8Qqt2X84CgqaIn0Qj1XNR6ga6Ko9ZU9nE/cuajVe
f67pwxh5FoQ06OIrvJfolZ4HVOTNw1ogZSNhu04dVyhyR99KmXPiODmhopl56dop
0zuaZLYolb4O4J+wS+s3/8x9luCOq4At2CJmkon01J4=
`protect END_PROTECTED
