`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL50bdeZhVsySYbR5Wq34GyQFM0DL/2DadNzWQiUinvh
p/yqtDwSWMRjDB/cuy6MGSQZmZoDzTaxKZG6XNyjQKaL8n1lJiy+LHFiCiSGtkle
cy+292UazoGlgFpMERj9+34jcULW/cFFyAICuX4yC0G6aDrpd5NWn6B2ZVc0//lE
HS73lOE4ErBWGCBJSf5ZaT1jBciVt+sXnz1O3fSNATgstgJFRTZ3mjF+MBqey+ib
X1w6SlH4fpD8D5b8qg7yhUP4PJN4JqkekA4gZKMU5KfJjaanF8hJyTx3EItUdJYa
Doc7iVVb0+CeKFNd3sQswbC+/OWVvOW49buLF4GaJ0/49+9YLNOOx0IbcmROXBPN
8DM8gwrzY9Pav5KUOagUhB93EQ2yL6cmkX+YGSqCUL+5joQlToKCBB1D56i5mNBm
NRoSCtortmNf2e8RpqxjL7zUh1iNinW62xnu1uK1lzB/xaW5QwfUcC9zvZ6sRjER
pg7zXpUx2tngB1PSnL73ExbgFMOP4Efm+CfU3Hl8rmtrO9JeIQLAGFbPlpf7nZpo
`protect END_PROTECTED
