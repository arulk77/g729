`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLot3F2vUBf8wJj3blqjWbVfGQ/FRGTIPR6mZy8E8pLB
RbwgxlY1cOLrLN7t4UPaJR5oHNJYc1kSRUfDEV3qS2Cee/5gHaOmbIelxB78aK+t
ydl/pTbPZXIMkthmHZWQCcmvZkBxAB2xskk0gs1SWDjP49a8m1ovKPr2uyXhcTNL
RJaqL3pKrA0CIIvfLbclzw==
`protect END_PROTECTED
