`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM/Xq3SrqSrSNb7fk4elYK1UFEB9TrQWDngh+YNiX1oE
GB98mIXEwRi8lA2VLPqPau4yKw/hTKv+gDu6QbrkUxGKNaG6g/MprKdj33OHBzju
ui9Gf31966/ZdXG/0VO7nh8qGr4GDAOP4exOiRfso3NHJ+x4SLgKEvUDyl+Q8EKJ
sWj4Aj5vVNkRhvp89ECNgpWGO0jPIztc+1MRE+t535NbD0wVpWYx5EbdEcEI/MAB
D5Djqm8r49txc0niU07XIi0ntEtOv0s9pZX5vnO6WrpH91H/v3c7vqmJqEC5VGXF
dpsAJ/ipHY9rjD3lO6GLz5zbVMJlFVvvUY9L1aiqejV48MmaG9PGR9EG0gOT5Fi3
nXFXwhiSfSzFOs709ejNAXmkrZSCVSO1Ej1UiYC0UPxDtfZD7g1z4J9nyw+Zreoq
DWJjwdRbxb7RvwvkVQNyuqC4SItvXkSvLIMhGAohdxVTDDZyua7V9s5miULa+2QI
6zgLeCjUi6T7AF7dAIxpEXGSn1pJ95x3v+jj/TgJOoyw6vPjSriBWJ9e1Rjr3ct+
H+93YKOCFDaulizqvMNI8Kpo8ERTKliGC1c0GxRziCK4LJDdkXOTVD39x0Zb/T5o
TSR+oLP7jHzDmjCn3mI+H07Yw1pJ1r+SopUtyxLGuToOVgHoQby02Nxr/sn4/X26
nMTY6DkBxShNkkuzELGoXZl8KNumuo7omYwg+FukW9fPHoZCFlOU+jzxFDA/3uY6
rNhJamgmDxdLVD4O0CbVejk3COnigi1+3RitkIMyUxoRqrhiDhPL5fmXlM9dF/YO
W7mhUcjnxzNy20q6Q9O7sQZ5SmzgcEY4KdNSZFp8nYp4c3MvsviQc/Xs+8KzOXAp
JdwE9GyT7F9qy0KS8biGbBsQZucmJraS6B2i+KVU9oM7ZaYQ0i1EnkzfAZaB+Kxl
fE0zo+t4FBoGUMB6xrT5ccSUTKX/Ut/524wCbW3wau2adu7+1jArBTaX7QqKQWj9
v3XBhqowBDciBwBK5P7KKP2375jFH5OdomFNFb/pxbY+0OO1iE1u62Q6TpDxgOqY
oBA8ZmVG5M0l+nn19yPlIYE1iIhQ4dkmQW3OqnxQPBEM2u0JdNpHt7jZyR1ESA1G
8F7Wj3BgT78R2WAtsIkCIl0ZPLvTaXagZgoKpVyQ1WyLnVzbnmGz1N08MwV8wVuv
j+JxQONPOjf/GM7RfAcdfy2LDWHCBwDGKAiZsDyFe/7OTAD4iQOXl8JjU0vcA8dX
YLfA8z+n1LwhW3aGS/1nuqdguxelee6K8gLcLKTEHmbskIgtXzvSpY55VS8rwsC4
mMNJfTwtXUSF4PRvTSY6ovWCI4tH0cx/ZSL4REcKKmvj88K2NiaKNTdFP1Q+udeo
ruhsoSOSpkftiVi/UX83ALVoxeYRog4mrNU86UZo7MUePHNe7SmG2BSzEgBPRmZF
9BF4DlJg95v/Ug7TgFhn7Ii2phoB3CmPDtCxtC31wkbXNCu9zj1s9QAtYnRpEhcz
0AeBO6JyGqxymG6XVIxs64NUm8180NXJd1VGRTzxV3tpgRbrCLSXzYqvgP0MwEhy
urGv/y4z8tIq/T88nubvn/N/FlgCauP7KoHft+NISdZ0ylApWTXqSoyTi57iCv0a
RRy0tTsRWxSk7KaCf/L/UeL4bNiSMHWp0lxhJQ7Zm6wluT0NxWL7xH2sA73NyDdO
QBoNFsn/gr3LrJg8RdvUqlkcxGPH42iFYoH+gdyTEsQ1N7j2wiIE+zBgiYIcjP0T
7NoKIdL5dhvKWEdM+aencReN9/Lyu4BOcgflxqgNtwgWyNezkYrMuhvyn6eAR5Nh
ZOgSjib2zHXKpe6uic4FV0KDwliYnggs8IYneUtTp256U/+6DV9tugi8CKlMx+7N
rzkBtVvMZ27F14bH5EsQcmn5qf08wODF7HmuMbd2ItM/pNm3BE/Mso2erAI3crTP
z2F6c5hKSqYwIikGqJ5NBrSXwdkr0ayeXhnZMQ/krKf+gmET8djASTze1+DTKAEp
qpqae3emoefUb/Y5QZ0r8NnJYGFclzVM/WdMOcUFf0PqZQ5PIXhfdhTPo+oh/NC7
31XslbjZ03JshedpWRKaQ6ATgW3CfgcYECj9HkijDgFWBrzxYFBOxAWJ9IlGYVzS
bmYk96i7AHB9WRwREJ5ojLXG5Iab8juU8u6Qn4XPrqGnE+VNdt286zzthXO1JBJh
XUexJBFxL7m0gY11YX3rPNX32oFLNqpkHEoniswgUGd9XFpj3Uhyq8wYZZixHQTG
9neqf8fn0/uq0UiOr+vh7svh7tGcmgiLy/M3s6+Kt4sdHSptO/5jD60HprADoild
Ex+0CLNgBZ+vJ2kuqs5D337HGrl6e+K9+ox+I8ujSUi5I2XMGvbaAXBYjfrK1gO7
BXswoB3NuonVB5aYWlOTKOONE2mo4nL+UUZz40+S44XWeIc1jY9z+IDiuJ5fH/om
Rk0OzBPnmcq3Wh8Qte1vUzvzAhTtYeXHAXk9Z+PviHgcqZEPhyqRKRyR2hk7wDSY
We5WavL3SXE4glr4MpKLHK1oCFhwzX2SYoVx7TK5CgjGB1fBPu2kv82hBo3SGJcT
+QQimsaneWesbGKUV1oILaNyvHe42Qekv2w9eRf8CjFjF24HaS37pMCW1HL/yxzT
e3xMGNRR+anjegvNpwjfLCynRiSv5bIDZeqq7QeamwGzUR9JrvW5EZAZAaaFbAKi
eb/oI/MGPfmg34JwjHjDLdE4OCro/ICZg/hJNE4aNRJJco0Iqi7yspI00cY25vg5
ukYPTApyjyyksQqONqKz000iw6MEuusL2OC2iNxN4OGLjGArXiZf3/bmdarKcDVX
QDtIX5ry3B47bWYzvR3Tm6u/XSdf4k7OdCpQtQHb9DOZsTr2RG5iM7RMOLxDX8zq
caR6KnP92sPe3j8LpWgEIEV0y9x2De6TCR4/d5NxXHTznmGUvm3JYQM9Sa4jPfuj
qoFFgWHGwHO96OqFWyNde0BNK7ehzFRE/uvRaKBnFooxY+m/D0L4Rus+l9xMJKy5
Mh3O5fQp2BMmM4/LoKG38DJwR1xo0TkW0kIqr/gz8HfnhiynJ6ydakT7gClAgN4N
P/Uh0ABankz2U7PcNlQwV7TIpcaeH89p3FIfahUJR59lbEqWRptORG6k8OMuTvzW
AZdmWMj2S7j4JpZafK3zMVy34Kvfov5YQ8wx/CZ655oC4Wx1hFIWhoCufEEZjnV1
jYDhBihLWukd5IpJlexDNxFkJZtfXbYw4tvlzNZpEdlLw8dZazW96GWDob/Bia4Z
MUK+IoD9ZAyOtkDyadvfgxmS6mg2/+dZ2TWYW8oqYpTdY302Yosqbi7t/J1uzVvT
t/VW0JNz1xceQRu61ZLJrtRa0L4mY/MbJcu1x08d56ys9AmGgjl0XCKa4V2WVGKy
8iM32nbWLQa9ApyZb/e0IAGAv6by5AwKCXH8zP24ObJWZfqq2cvkHCar9mbay1ox
qtZigmTyR9rish5ouK3KPriNo1uDPRIWap0taZjMCDzzZxOFRAhndIQxYGLYmgIv
rHdLhYQV3yqTKqH5feyVoaCcfPuEXVLpDZAgP0NQ4fhlZmpS8WhpZMZztQF9KVGm
hqJJOvUcNr13Xt+dxQkIR0EbV8PcLxaNMEz50pkX4VAYT13EMdwlxn2xaB5ZKFqT
EHxAv0gKN+iRA+Z9MT+77R4o4rT71KJO4NqSQ2Uk1prK6vazglyObnxajfHYzumc
3NtiHMJQs+CwtxfrSPHWNSBPOSRAx0OOCnUL+xUca3jwWNFX4JmiU7aNb6lZskSU
HWEv0Eg4LDqV3Q/UVDOdeBIb5J06KB78bB+BlN4HYqmeS9hHHG3JYCf/mU+7LezW
xw+eAtdvk2td/RX4appdHO6oTCcR7TMgR7QWYzYoh4Xa3GuGbd7Z51nc64RjeGEG
1LwoOSHN6Paqi2hPKhsES2ZfL5XdTbCcGal/YLijGjsH9KniDZ0fqRQIl65LPIvJ
dNLVKfmBU40mUgqHDFBVNUQMU0/UZDx3wGJP/tTYMiwf1K5qcbdKpO4m7VWAAMnz
0f5x2VbIHO0hD2cCBsUivUfxLl14t8hQprUeq+l0jI8KPeLC/vj87FyOr8GiKxK4
KuwH+ypdeLY1mxC9jppp705HwU9/QrXwnBtj8CAOp4rFmfcZ2m7pjH1oKH1/V1NR
y+0ABmCF5vdSkIIutK/69ZJrxvFWtahfYun+MC+ZWqp9dpC54t4x/Vz1MxQ7SJbd
2dmoFvTw8W7nNdupAAiw8utGeKqPMBpqbmsOyZSFIEmXi+KDYTjjkahpoXYNqehA
sBvjK3lkKYH//C19gUc+7BJm3ZNX7t8UwgRENe4MJoI3f6k6TlIhL4Zqp+bgo/IK
E5Zr6XQEuTDoV5qjA8MsMB6GyZ/VD/L+aije91bFSZwVBXRlY73hxzFeonDxrcjF
Q2wujXL5O09pMKe4yGvsJTqs6dxZAe9uf+Fz6tdPXW+pl3tXjULKDhPO9hc84qkB
Lxp/t5RwLWZDY8cRdMI9IqlZVW2q5Qhjf5irsNxZzANtjt6lk/it9InTaQjAj34I
spCUpzbTLvTE6kT3x1D4sOILWHzDhhyuMTFRfnQ5OgD1NDNbmV5xDzk+nrupI2Zn
btgJce7L8/Eo1HPGl8QP+IuphxTAsIyiValY1fqdPeMQaBuxphxfL0VoXmfwBQ3/
g2Q+KkSqRo6jZPa80TWe4h55oA4JiS1xHKmtZ2L648nTW1GvCnkteWjpSYOovtc7
Tixz8ONFeZJviTZNFoFfJce3xVh2AZpKyTziQ4kus4UYR+2/dEB2a4iifoUG871r
be41YM1zzF1iXuXyyBZUEyhwEmU8854PQE3fja2MGhSzmRywlNUV/pT0FXjdI12M
8eyKtsM5KAlc9815Pop8gJRqAP1lMDyh0kEmhUBRdo3rOC7+WPTiDPxunpeQXxDG
9uZDwXvpf9bpHBCGLIBsNGfkR9DLiVBcF2qlJw24hvOdVidIFEaMrHVAq5toijCH
LuELz6S7Zp0sJ92gyBMnRt9Phcy6zex1lsfIZFrTuwiTIdhrMh9FidWppYcebh24
bMU4UtMG0ePpuXz56scS4vEjT8j8DT5NiwxmacZRL3ztYqzUOyTZmjSs9q/elR6m
kmT8lWYQWEQC6gw4F7UziYG0apAVCBduP7M4j3eG2go1UnLQrNMlz69Fc5IokKB9
4jwDcpiugGN4TbKa6oRev3c/dGZ/DMd4ZogPz0WpCgWV05fAl5Et+jYs2sX0zQG7
THtOX1Q+zQ4ofsCGuoxSJfC24wHoWHJlJcBDwoND/K+9O1WcFxWZQJo0h2179l1C
FRKFkzmevUJrBsjrZjobDEK0jh10mY0YXQQSYOZUVFJQTTY4XY95otOJSrcMhOYx
gfKcGY6Ggk5LaqKdoPZ288IU2Wfc1/Y4E2qqyOmgmDfLnocX49m5DaHrKkDhSRgr
YSfkI5n4k253JOX49BBL1IH/GfneWAh6UkH3p8VKh6bhWVddqFdVEAWy8Am0i9H8
cewwZrx4a26Dg26pPPAe4Volbo1dno7U7DhW59wlFfs/S05kg/F4HzB5FSdq9GcO
KLy2oaMz5eUaIOgwv+lxCDQSCFM7HfE2oAeKjjflDkWA0B2+VN4f5gD5Yl+d/cn5
rrhcHb8bxvyGLPbG5u2kA7eD16XLCQWH9ZG3uJkPJaSpBIg/MaGB9v6T/6JM1JVI
9fT6qIYwzS4AhUBk092JE6G1Tc7PXK+hF9v9HxarcclQEMQScB3mZfCedNBGT8Yc
whgqJClCwLS/wvMRhsVJ8xo4Lq/c9E412/lWvH8rknmpEV7xUjfhd6qVwlFXqwl/
zFerTR80BaGy0vFxjAZ2sr4PrFtaR8Hd6HURvi/zljdD5WnunRlv7Tr0BOn4+Qnz
t81FnYIMnWqQ9CcXqnMugnfdn9qpXGVw2yQOugydlHjH5Yw98g1oECXLY7SfhjQU
SCFCQjIcspSbSYQS6kUvMsWiSf9T2Lyf3m9Swvv6BySof2hZWaueZN+6/E0NP6HZ
rEBYiCRFwDe7z5r5TFyquCDk0KbRwszqe0KUPs8OCQYiy7ORs2fMK7CXyfcXrIlI
P4c6xBvc7n4l0w+/DYE8HSD7o0HOlxZ8LL/Ezm+PTfWdjobPAKelAyvdSolzfYCK
LxghdbZlkM874UQCvQdvQq55RoNb3E8Ohw42RnuMEKSRWHhXW6LdUVwHCi3FncV3
ha+8i+346abtQZOtNDE7zxLBBMlSGXO8o9LuzMXoX0d6ZF7bNtinb7fOgEZuYuBV
KvdtekoiiggUkwS8RGb5bu2bQPJKR8cuupU+birR7EqoP9oFQtYEN1ou2nyACdV3
qAhF/JErs+dXu+KNPJPBjZbs/nTvjrntreJihWuoHUfV067nEvr5If59KRHzJfql
XrjexK4opLLhDal9ARf8Zgwl/jt1zQf6xr/UIz5IbrD2SDvj2W7bvkH3437arOP7
lVTgR0y3chnfm6R8GNEZgl8SNZF0N/fwutp48rnG2yFy2KQVS4eMWoCngdrR9CaY
iauhiDVdXIsxLfJuMNRJtdZAA0gqfgLxmwBpTJzU7bt9BBGAAcqTfz/tQ/zBHGeE
/iOkj1e5BJNLKvZUGnjzX98L9NZqaAQCw4F2YIO3cJ04V00t8qeFPlPURujMCJ5V
puUImjVJW0iTP8zocTMBmTjfmo9uhATs7WQk/PR/V5DkWX9JN6gSnfh6bDqw8BoY
XIHEDj3ArUvWakQT/7rwytEN7+FWQz1NocLSZZPOa/P1saZsodmLH9tQI2WtsPzs
hSCJTba8k2HSbW6dMn95e+l9VSdZKoMZoOoS6fpWBV9SR0q0EDvlObJhMZcv311/
lMA/7X6i0tMHGmSAmjb3riSifCpn9qH+E+j1m+3DGJkp9c+q+B/sJSDBosJyCAOq
Zw3+H9wxCFWOoB4C7UzDrjNatxKEI9swnMipvIAvdtWJJOhGzBYcpNk/M+MeWlf4
LhPC1jTjPCQoTJu4S6hv0y5ytUiWorD7mhotDw+BLp+Z+DGLgAvGzTVAOoi92RY2
4CzHDCgtvlIowe9KPhRLKSpgb7dAcYFTFKwgzNLtcwbJ2VTXCKRrMzmiuV/vApLp
q3tZ+znvbGSmVgRPvN8ktFWwqhLLP2xX5yYw7zwLw6XH1OzSkgVqHH2BPyJzPsqu
zdUw+BQe/57LWsDwOjTwguXUEHS+lRAUMTd1AqZQSBEF1Vd5XKtJcKo1/Zxap+7Z
QiPDSUF3TlEx8+vSY+kGuqAwwKd1I1+i41r6D9lOzS1jhG4XLL9iqAg2VDd8+ZZW
sAp/8I9v255nT7RG1Z2AycMtda65CCFzD6vxjfXnAAxvU0FTON4Pdci4JyTp2NzA
aFCDgkunat+FUuqHkZQKbQ==
`protect END_PROTECTED
