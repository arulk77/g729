`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMsNpKEJvFQFv9gfinlXHVYKopvDIlrlh2Yl4J3HTGZm
aZvWQ8+cXmaa6Jsfl0TinDYiaqepf+wGBsJev/un6fAX23BIAICOQct4PgYKDpBP
5Zd5k8kPwF2Emi1DFg1BFBZR2rqHIxhKDsFSmkYUy+CnjrPjAMJS8PNstrcwnHRn
Miu01373PFZ4lX4kwXi8Nb2DNrtUa6QTGYjWOU5w670MdnFVR5Np2eVKWrxrOm+/
6zaDSUtkJcOuG+dY4SAWH6TG9ho96c3RwYe09U0jAu++B3wo7921V22FehEIrgJO
vM4TGSaKxm4cm6kv3eZH0Q==
`protect END_PROTECTED
