`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOhWpSL1M+SL/QF2cwV64J0PY6KRlv0T5ud7pGJ1S17s
7IMZu0Bb1XEGRVf9kH/GgvvJAmiYmI7vYZ5Mlwir4YPCNP4aefY664QOziOq35gH
1ap3xR5McqTeHGEnnpB5M30dsnKl8h6DIS3zu+tZ9a4LyLz7b/HdUsgxXZvgnkMf
GQ8yn/KUKgQZXdGvuAdAR4XGRMkfKGweno6ENmYXOAHyFrkMd24jUvaf+bkfLLs7
Gqzj+VijwVOxbqyRE5+FBjIkqo1GA0evt+3JmoPxuiO8Cu5IXEGbNGS5keN2pZPw
FPcqy9KLuHJXVfYMDgFUIiJn34Jp7QUCege5UhAI/h5EExpKN9nJ7KF3UooVwRWT
tx0rGh8FMsn7mL28e/0D3pPLTt+8x9tHQk4218EqQndha5jhObZt+8ZRQ1sAuGmM
26UPD/s0gy0hoKU4pA3oQnYl3pnL8vPf8MpCIuQmSiz5GB6dxG+JUACx3OvIrMnL
hP23n01scl8X17ERJJ6WU/Gew8mAh8pelFB0lbpayHGAZp6pP/7VzIEF4ETtnRF5
1dl0PYnMQNDgGl14Xmah9+iuUIN/OppjqDRhCpIDpptVMOZrwXZI1sbLAJnw2dGA
PycsK3vO2m+glAX567u5rphKNvcoa/KxF2ONOk0x2yk2C0wWQwmLBeUhVYirTuf/
WafQoMzMMD2CmSVMM7SvUTx5NTmwKWhkteWiACmdkCcPVX34cVIVXNcUF84OKSWw
BDXCGAEanYbV106WOPFRmw==
`protect END_PROTECTED
