`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIrMyHZ1pcYwe+WiIYIfWW8Y6iZqcVTkBvl7gdXjveAn
k3bqAvKfvBwlfFgtLr293r/H5pKHZmY3ie41oYrNTfX1LiSqk/oz3D6pmvsBSY5d
onF1n1Dt0zY/9gOsg4CCBRpvbbqBKY5MBxhOom878YT4D/xbufTmM0CcgpugbZj1
dGY6ZoeD8E5WS8VlfVQC9Xv2F59KiosQ7qwDmihBAarjGHIgIDcu6Ik9Eyq2ZFKs
0LfPh9sbkNBbBqc7vNG6L0ju18B8+2MzT7g8ICLF/QmC/tfyaeEo1qWaRvMg8xTS
Y96fXKk5KyC2xLsBoc9ElV1QZy+7567nVCRdhA3+YHS344EeCertUr3UPHtXm/1c
/bNByrAorinq748Ckfv+2Pck/R9DybPxDtdWPKZ08AO1nOZzj1Q+sKUYCspmd5gX
2FNnedZrUemcGhRVF+M2hipMArLnlaa8gM2moBOP210S4L8n1169PohJQIdteEzu
bBYazcJvgsRQGWDh9JVqiEJl1qBvUxFOlEoynZfu1yJG6ABp/vKxIkx0x/2Ff3H7
XdwtMsvUulA/QBVkzSw/6qTtd0YB19EfJwwFlzYFJFvpzTv51mZnTKw69G7FmaE2
BAUVP8q8VpwJEa6ayEqig+gIXdvQ5uL5T5RN1ARQK5VhPnIqBPfssUyP0NaIenRp
`protect END_PROTECTED
