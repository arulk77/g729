`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
W9s0izKBjruQzWSMITOe4CJZvISwdL4QVF91/miPp2yY2EFplIKZkSZu1NG/WOAv
8ibQvQqyi+ecZ5AanleYZtL8mtBF6ZuPhjfdIPTGU1oqfySpoqTg9Ib6D2/jBJ1Z
kGG3YKkX874V9IsV50g1bu1TIJMGbpJGkPP+yyHaJ3LWN1fl3yNhJP6oGbH5QfTL
Jx8igAPGWaKd4HxqOkBJYWqbyVKyoU8LT35EdqtiSv22W2WiNxrv+X9LM8BVlFmH
RwVnJNZfy5qqJ4S/vyDKPb5yubxXXqOcLGCNHKYARzmv5rR37jaa9xN1XDoSUu5x
9TnY2iDD3OZcodrekbWdr+TedXfzPtAyBqf+oS6Lx+9oYcU4JGD/K31D2Smog3mS
SoJSYs9XtGhWOfGComnBj+mEMQcWirQf5Fy/N8q6E9VIemx1s5fYz4Toa7ulHlji
/nPpD81XOHEMGMceE9PfMOFPQRtj6Try/iskw7il82CtiHzohZ21G9eAEIuH6pit
NrhzS5/J813CGujgasChLOSNzdpujpUwNXnNS7u7k+c4nH6ptSbt2vtsOxiGnpR8
0C12MahOiiFY2RgYrtHCZfmzXCqC3irW6EX4jmiSjWx/3WugV4MiNhUkzafQsvym
31O12buhRBqd5NJYrauLqw==
`protect END_PROTECTED
