`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLbBYZ3PVxKnElPRGP0Q4zaicVzQsQddz8dMyyvgG6Uu
wbo7Ts4ygCxq2cj0V2sHg113L8+QK2swYqEcG5XHpDErAI8tAf7+D7PFQby4xElh
puVEQiHPwpDphu3LtMa5L09y4oRqHqjkXq/uYwJBEQ0AXjUHs/myTd1B0c7SlsNt
6W4oSvceInBkSGVxT9sEaQ==
`protect END_PROTECTED
