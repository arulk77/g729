`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAiLo6pA8OU+RYXftqCzr67LB75g7z3PAYwQ9tsdnKCM
oreLsJF0QPPzIflIqbYgZhf5Onh4OEcd4nUDQiPGFugFkDHZqkGNcItusdsgWK1W
pUm4RhDJzGwVJVApdfqKyeYuQ+tORGBt1Z9C+/meQfIGWYdEb4utXdJ8voFvYehi
/uQ+5WU+NxAHNPjYJtFnLQ==
`protect END_PROTECTED
