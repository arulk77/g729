`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOGRorLNTWH7dMyIFOiosbfKPSzVsmwLfD9ZOGAd/zCP
4nUpZ4jDwKdPVTlo4+LQaXJKyWDsrKIPtMnwUSBIUEVd4DR/zT5DCcfgFytyLdPi
Vv8LjugHs1WHMc1mfO09yR25sbmutd0E7rK1q94Kaz7XpVipmFeZP2tm9Svl1+tR
CeI6OsR4S05N4C8hBiXkGnmIU/CbBPnbsmxfdDDcidMQ1ILj0+IQZTPKfRVI0HtR
MiZ85PiI0pYYzhjLSihGKVuNFl/5ZULQ9pQP8n59hEQsFidFs8mTgxiTgL61AAv5
24F1152NHMFpFpiSSzDIVB+O0m7FjyNvfHWRC0TN/Oaw4gW0NkmgzunoYg05xsHt
9vardKheXtk8lRNaxVPn9g==
`protect END_PROTECTED
