`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLGa77G645HakQl7L9UVXaERGq5qEBZtfMEJ+Bfef5zH
Kmhh3JNTp8EEQERc74HwNK8cTM7RfpBOzkSjbzy+GcUAfh7v9DQ3LRn4PByr4CtA
eCSQc0K36X0PY9PreIsuKlsJoQeDBJxVikTrlqiWyGXIanlmZit4svO3orgno2DN
g30+wagpmdndC0DNtqmpmuoCBqnliValDJbcj79Bv8CXjRAU7OiaNQazpOmAfgst
KhnJKClK1X4kflHVP7OYKlg2ugY/c8Texrt3MFqquC2Ul50UiDz1eGhYKV9QilzH
ZXfYLNeYvcE0nPVxeqABGqxyja/6unC6iq2V+u7eMlNCqM6TaENsOfYTRwwDCWun
f86Cw5XDRbfpHPWbrFYjO1eMOz3sMnreSjDsYy1DOz9XkRIkLU+Tt6gOwGu7N4Gh
KMi7u0Qhog2Fp3IcnpxMipnl3ahg/H7RcTg65w8zmTxiKh51C5o2gI2UnDW+T3NC
GjGqKAHkyuXBfO0ef0kGq1YZVaTyw4lf1VMnvVOlXIQE0RkxL1oUOq2qW+O19E0B
BHYdZw/QCnmuHjg/ntzlfk2Ptd+A0xAwAQ3VE2vUxfU=
`protect END_PROTECTED
