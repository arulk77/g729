`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IyaNjjuMpZLgBXS0P9ar3U3z7bueFOhJibuizaAOYVh/M8xvUSA8MphXbTOOuJH8
cbSz+SxFZQXExVJfAXf1y0xoFJDyKwH6XUIT2OMYWhr267tQajWguDzB/JcpI4WD
lS0j3XmXpkhwknUYsO87g2YCSv4eoQ9eeodLsaqlSbmqbSSWwO8wAR17/331cGSn
JvwkSGP0ytHfpHd1yThWSBHNghlo5TPHiHGW/qOHvfWngFrsS7XA69PhkUuIJeI3
ZYoeSGiU9JrTuYe48FvgfaDLHuQ03W1LJqFbQe/Sy6IB7BunDm26thSdYL+vvj91
cfQJEqlRMPl1MNa7YREhHdGVT8LZ/yO3jquxC4Q3uL3LKAnE01Q1wzPOxaHLqZ6k
7uSRqHeYTiRdvnvAHFvCeE1kj/XlpJ3GhD96yiRizttEnRrv9YmO3UUh/01OpjSm
DjOCwQoIgOZbV06G75++ODrRs4abzppZGR3MYpNlIY7qjUgov44SaqZpzB8tPiP5
HQm7oZ3Y/oYbrMhBr9E99cknSbuCCfluvmBWKZ77T7QB/RA8JU1YlRJH8s4rX+yC
xBYCb+TjkqsvjbhUS6MJ2UVA0u+urxz0ob+5tuMXAyFOFgq05Wt5ZUVGXmhneHKL
jXeMAzlwYFeJvqe3P3ba2fj3SxLdxsfkDhh2S8H0SX6dCc6RRO4ggqfYyixjQNw1
rdsHSd6uX2gPOIKI2T1Bn9fyCI6J9W9wPSgXo7Vlp0Lat2qF3A56z+7q63moQl1n
FK61p5DI7t9xQXX2rBuKGkJm/KX3vXGQqRq13WbkROjYSXPdPRC1UO/5T9KZiCE0
4woTdnXWCdt8tcxUnfPDD8bwiWKZm6sU5ET37mQWGstNCDyEupQCkMubiqqjpcMF
7kJ7wHA6SpVTv7VyakKWY8s3kFtAIzP7GN+ORpJSZQuRZpqJPf8jmp2lMLTZ3SQ8
aRFy0yizhklOwWVnbJN0HcAX8F5pE9qvgnhVzeM7f20Mymhmz2cy5aCbmRGD/0t4
cGGuyQI4wq20HEB4IkleCbXL55Zz8kuNujc+wq/B1cgv8suk/PkILhEsK9ETAGmW
mVNtWS8d4AaWNyByrsT+LW71vAFsx9ubnZYvIWhbGGanIMON2D40sthKO30LMo8h
i/uPCB7Y6bphZ/HzCoc1zxLixsVikt8DlVMQ08s3wrRgd0hnyL2CGnLag+NCUqwA
NO+rcyFb92Sh2pj7BDl3pPaAG+Fxw121wV9KvqxreSQj4tFegw8ztuYiekTNRi2e
H9tdOmdH6t0FBwnbTioYnT6L4UqFjKfjRuFbV60KApCM2L20QjLgZfqZyT0jQJ9R
wQAitqiTm0K/VgPoQHTKwxyVZ2L2bpkIjw76oELuKrbgTNZUHj8s9pVIAdCDBAY8
BVl5MLdtBUTaZssOJsExh9OIfosDh3KTUbaVGjYuxwNl/exiVN+CAVIe7GZ3ezDR
3pM2NGLwUuptMmUQjz2Hm2lOPVc0/jT/IYXCEDwP1tkYxYz1NxJvNRfoSF7ZUZzS
y71FxSRzzbTFp+Nzjkg06WfYAW6uW760okn1vXkzIL01V3KRoUq/RupQiXsrJTA0
Dthk8aKqbxGOzKioOWwiczJA1hDWmA5V4Cp71J5mYSubMGcdfaNyKGHYIqZkdTaa
9eN/oPi/smxSSTq1mbU+vZho595/lMx/n4Ra+HK0iEwID+tFQHqfYC2P/iD5j3LZ
5SDwZzB8CikrZlyc2xIBevZrSsp7MkLuXNZUVKoVPbWQ5ODjCZgQfNduzqM1dE0n
M9kp+uXDYbnDjfdJbO57onANOI6zQrFOS9oI+Kdh4g6Tm4nW8i3RZla9qul/rypa
fmYndIxry8ppBVeLf8Ep9JnVjinS7ke/8k2NwXl0ptVA2m9pC/c835ciQdDLJN0R
i2mKPeAeX4NdxrVt2wqvQCIcfm/6JbXmRSiODjRseiGaG18XQcw4GN/AqvezqV2o
On+CK76uYQXH/9M1mHP62PwF1I+X0A0o0ZLF3jVVjoRI4fosCaQz0oBCBusbNSz4
0oS8tH5ce9nec8nH9JJcl5SRLhlcZtFRpUYwxaqVwg/orYsd7RohKZEbFWB7PA17
N7uVs4qgr1ysEQaKAzLeYfxVX1laqiiftlYfJzs47jRoGEqeRaJp2l4Mc20tx2H/
UTnmiAEIETAMllMRhXuJeKVsHqyyptd15OH3fAyanLBRH2EPccCb17mA4ml1XQBT
O1wYpauvrqZl4mgWtQxqTLn4M65J7T0ImqHdNQP6mBM=
`protect END_PROTECTED
