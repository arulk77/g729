`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yqWTgSwL0bV97mrBA4cKtnFYIcB2I25axLnCeCgvg+3
CrvQILO2RwyD5YT/097SW6c4q5LvGIDmAle6uF7mTpZuM4aJDh7VAIrYHJ4v13Ac
nLm2wr+h60OjfK17EU4CuAZp2nZDPGDsOzU6LHDKdioR9tudoHnQET84zNi1JMUc
eX+BTXtOSVKfjX0UaBkTfCJyZBT48IzFFKh/hae4wTTbHsyDzm2CPvrur7hp5TYV
BA39zc6h+X4G5Jd1t9FUd1gbZAEr1p1vidDmjUZjWJvYFx8fiJYCFrwq0UXHFRVE
FX2Afw2txBTxgj8wXU9794yMSkgxNYOK4ZLNRNqy2qfHrJLeJFwJAhzmx1F5p8jx
RsEzZHPi9U57yfMOJoTPhg==
`protect END_PROTECTED
