`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIqozQsNwZ/nAjed945iTd4sA85NCMosjsE4Q9f6Y3r9
H/56k15f/ggMPOtfgBZAolI8/3SetdzyGOGsOmpGNDHYyABB7+qEOOD9dyC+wRre
iA2LxWNn5Or7z4wS5UnucVFsmj7j3s3+FBPAreJAt34rqVSobgKRDsgtvPYM/BJk
CDLCX39y/r8hZqYFRIGQcQ==
`protect END_PROTECTED
