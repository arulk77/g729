`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNctHfC7jFQcbwW7AXFzrTK3o3WXJVaMRcIKw8op/nVS
NW6X3I9398DBd0ON0GMnzT4AovJWoklbxMUaQ619jXbSBJQEShsyxEb3+8ZvkYv3
KTDzoDtuxSg0LLqO7d54rAc42d4DVHIGj5z0NFcRWKIukRDGPcRPYUK/58bkNITH
pKAfKUz4TpKcHTba/hgfq7zSYmmpSxO6rNd7OspEeBdl01NWP0uxBCoGf7ByHz5U
Qb0b7lEAVvZOzxNx3ovblA==
`protect END_PROTECTED
