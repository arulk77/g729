`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJaE1wvANT1l8Q0Xr8PVdpjEKnIQySLM6Unb8Ff92FRU
TGUzB4ZA4UQeKEAkORswCAXweuuNhtws3/54WTikgT7MFwiG9bs3n9KCI8vd+255
PWxgarMdKLtC0NwR1ZU6UVIpUtAteNsD9yUHFNTjckW6IE/52Edn57hsYOMIeR42
0gB+ZX2CblwMVhSqiyoIa9huNCeYLLj/+n4o66GD7W5f18PUmWynpfvvDt8YQyFB
MW5RWls2fxfRc2g72ro6symTvYrhz7Bi2pid1h7Ifb6kERKveq8+3b0KFAhX9Vwv
3Y7ooC9reDCosW/UIEZSn1X/wZ7bhdUX7W/Ii5rGhDgz41l+da97oukjCPqPSwyZ
9weqA013hqcnM/ZwxhSeMMBtBd0KHqum7EFssLvHIkHJVJZh+28l6l7pXSLINomU
mZu4uMhG4AEGltJpwgolLlDlXbuGkYC29DjVqs+29uOET1pgZqgN66CubjxJ0U32
ESxyXEsZNMuEYsgue8FpXMdk1YuYaipz9H5IlJhbbRs+dybYTaLNxrSimuBtFtv3
`protect END_PROTECTED
