`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41Lt+Ra6iyCICwcDi+ZK/7CqtlS3ENBZVp+51DZC8Ewh
jrN3T/PoFuyibJ1C9IDeTmBsTeqXJ6W5S1AoLub1H8CvJUbN2GlLQNoyhX5WAglH
505h8pHt7vrKemL5hCftl6SPPuCzhe8rdwJuoGUct4S2HlHqHJgf/AcNutfLxt2r
THOeQNn2DpebKaX79x5oA63witN37ZzRleTEcTeIn1pmJ/9BmrlTZdxhJjmVSrOh
E82qKRLTD2eCzIVq6SHcU2nVgY0o4mwzG7FewdzoxDPHKqn/I7LPPIIYidL8kts5
nTNOVx+AVUSWK5grwcd03z0rZROkqHzdoipWc1hGbLBiik1dCKgVLkS1BHvwSj0z
oT5bmyqHc2EFUsE68pJImA==
`protect END_PROTECTED
