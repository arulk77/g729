`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SRxK8FW4lsEBXYDROhQ0uGiJd0RG5kygSK1D373JB8Su
QlNt5LPI943Fn8RQicx1totkMdWqR5I1XmABAjjgbmCa3WWzXX4il76N4LZS8Cl3
0rAdYkT9a/jtdVpBwb6IboYgKDv7EAUHeFOVGznce2Ig+Pr+XA8jL4zlCepmJFW7
xmzVdLgQLdJQhP7or6WvKQTE8ApbXI1Rm2iii1GGIiT3eof1wdTvJz770B4eQgNu
xuG6/C6oOBlZNL8qsrVMlaJdEutlXJnX+dUazZLNAhtM3wm628cWTofMr6TcBOad
CpZsXiJELtrAdVC1Bdt4Nt+gCtciT19KkyERXtvngqdOAxa4f6eCN9ZAPuPO7N1Z
+mpnKZdw9o2kSUApvaiyXDIVqTR6AYquBT1s4EdrTWZbyyNeURAzzb+HnrXxe4Ri
Q6Cr045ibjxMRyfRLGqgk1Kz36g131zJSIvp1+yXn7lGZDHnqsHM5+UHEl/mKZF7
HsjoysRE/nhRAZKQ7tGLlu+dUuH2vgpqPVdQV1zxCh4Q1ABdWfAA1qC4otQ0Gq8Y
3OZ9JCTU/6hcOENtsPKwbhoCy+t+X2vqf77+N69+Xx5GwU7OCiFcIkLn4ew+yVhd
C/Iaz879rNFvhoXMEhkA35FVRKQwErCefZbVXCCqnPm2zSY+9n2Ty27i/u/tXaxV
Z7f6xw7HcXjUvaKIVOLovnxJJ12yxYSSYsj1k6x9myygyiSk12UEKmXXwcXShyA4
4mRiVQx/qmanYalVHE85TFXflCDksbFyUr3IeQ0pB+Cmy7gw/bXS4Ml6zswxDu69
Y4msMdHU52WsR3NDl+SrEHGhDPS+oHpme4L2QZqZHWg85uYIT9pMHCyJqaKE5F3+
lAMOFWM+mzuIuHqfUIiXM7dTcQhQMRggbQ8/YFv9a89EhqWbwcOOC6Ics65UF1vH
Pisfy7qFY7CYlclcW50RMHRdKXnQY8uXhdCBKQVOZC41qxJDGNhJGbtyrwljHZiQ
1yg55hSM5tZfOyL2nxOHuynoFfY2tKVc4PXl6NYCCTTXOnm+lh6jGc0LRxPKuDUx
DKe5WVmbwg+u4bSVtU+OJa5ASbvD8L7s6vav9MxixDG4MOvcFm7OLHK5N+kpoXrP
kCqdLqADVTfsmcZ2xWd+HuTFhwn5cSP4Gb8NhqWTp74nOYxqk20B3Rq0db33wr1G
J5beSdOVIJ7C3CLiHvCpdns0Z3avigajlUVnCK/mUJKTHSBZhGBMLm+Udq+t/FB6
BldqJQC7LZQJ8mjk4F5CTAbBLrk085rvMdYRiagcFQmnPksQwDykusqwQgfPdhSG
QKrJi7iRVefKfOWKj3TV0G2s4xxmyRTmjaKFYgg1zoI0h+3nN4tbBG1MuDfwHc/B
iJH5+bdW0i1y6EFgpyaW7qElnq/FiBUy4PhIS9blKGCkP+FiE4vIf3xoPCUDIOGG
7csPn5fOe5xjekouxSgtQ/jB8RXN56FPpH2rhei4gCm3bIkZ2Wj1p75a7jp7PB2a
8mkjt7z8Fy3lmRa1iBrd5uFVJRWW0/JUrjnXc9LMET1dYi3gqu2AIfj4Yqh9UnDT
2pDouEsXZR2A9wSsj+HnkAcCzzdXrM+1kknX9tDmdy6n+V8SCMq4bpGBAJ/HgpHR
W34vDgbnVXZmr/cCirsTIvcGX7p65ZRwRNFa2HPuiTBTw2OZJgSY5J/zML1u7HbS
P4a6z+Nr9G0IEndSOaH0R/soz7sH9I5FZxST0AfzKrNe0gJlToPSBFHyB5JU6zsz
xBbOTOHKpluWtUFJN4retcmkJIkhMfAVSwacT6haBxZ0ZisiKOWv+hEB3MMWPbS0
dC4qGc5RDUiYJGKW5nWw1DEEX9w2yzXGNU+vP91HimEXyCLcXeyQ1L9jio2Qhj89
b0GLKgaOSCkIPHNiYMvxxIQQv07Wf4Dd2yAhMF76uBhCyN2bY5diQQDgFp/i0a8W
vP0peKXjh7UOHh2ijtBaukQf1xxR9hLWRF2te0NXj7JCg39RNi5T/Rd3fxfI5/p7
fFHTD8kx4GDVQ0HzFqMrqXo7R3brf+RqkrdoUDCdNMqcHnb4l0rUCyRz27LQgy64
vtKHK3jhEV5KZcyIGqfX2/LyiFfbPZJiVZTcmyWeZopceHXjbkj8MvXJEZb8oCIJ
u3YoIFSq5VV2MTXILq6tqmsY6S2s9PGib4FNUZmcsPncqvx7uF485JETU9L0JOvf
wZJv6oVLDWZX27PbRWoeeIJuxu2XN5Kxdtk2ibup0HYp24VHR8fA5bCjKIjyTzsV
90hFsYA1nHJr0RpKOnCC3arERdyBkQodRf7H8g17qwsxceZPhahDahKNgZJMxImK
8h4lpFKgoLkHXl1WtNI6CKMj9ZoG+9zjsTPYsC9PNZ3MCxz69lCLOwSKhMmBLA6o
akmRxny9V75AeTj58QnG8JkHp4t6a+o1WcNzzqKjjS6DVY5cUuJ1hSJiC0U1ruua
tvHdPwqMxOcVazvJDifj3CPQkpGmY4usL4uo/maiJRzID2iqKVZgFxc+/EifmgDT
674q5HnbQlqXgGFZO/AkFB8Blie2wpq9cMZnz1P1UsubJUPsB7yzV2C+rYCf4p3+
cYhW1ueMvgDaba7LFe/KUgVU/6XsO2+ClKcjZROk2Jtf2ehNzA+9r3MngM/LCwis
91nXtIByrMiRI4X+yktx81bSzXqIXFlCwgXUtgQOA3NkfyxQEl8rur6Z59O13JRD
Kgrwi5X4OIEVWLgIP25yKGcbfFnOQx3TeMY9h97MhapvWR4o5oQfnKxMbKawT9bP
5poMVxFzBCvkY01wcWfGp96z8X11SbaJ8QFGQbkMr84NKAyWR9ltLRkqL1RMY2rm
KsRHulxaE8YZdxx6bklNSegsbcsQw8KY/9Z3Gft4dwhlmymtCwU8FycEhSg1bRMR
VajhBSk11/ckhxtAK6fwMwrEt7IUJhwzUtvMP+Gb7nWtHx9asoQC2Vktuhh8A0Hd
3SzkFtqHSL+CgCvFBvG8XhhV91TYM8ve/Eve3bpU+E3sbvylVrhryTBibgmxI2Ot
`protect END_PROTECTED
