`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNx37r1vcToEIWQAs6YvFJJdc3vJa9JkY1geuTW96VFEH
mDt4NxqsaLsSb2K+vZSxCQ1ZwLo6GYbZmwhi5d7PFuyXjFYOjmi9qO2loYVfck+7
3kMrd9R85I3TeruVobpd4IZ4OaEarICXCgPYDbPgvCKxdaIUk+36vXTJlS9hiYhj
TKpqiZTjynrbDj8G6EV4F4AiqNehs9oeYFy4sUAvnMNLCfMBw9w7uTROJhr/1wiq
eJEG+Sx01T5Djpmmv+ebjoAPvPCV4MGOsyMxv3EDOQj6mQRKXj8IO1dhWHQ4BkN4
TaJVNiXAzIzJzU/xYGGaNXAZH2TmS6Doy6AacfjrFx6k9QNMSmmxxfMJAFEYCm9U
vk2bFeHkhZlqw30Md8d6JLwJJO5eRwUfIDOgth4jt6mXh8N+xGhZYg96FLCgOsCv
fzVpbeqyzx8ZB0w4qThacpvUU0QRLESOvT/sS6mIOIG5/LKYtRuseuae9Xqt2QoO
druiUSGK8LlApnSa2Kj3MqSHTNJ5TaJRk5aomQuSQFg+K05HRd5Wee9+lK+9onId
uplMxVj1+kp5jz94d2l3rTp69fGa5662Rv0w8+jC1UBwL0+MsViRYxnCS/SJfEov
axKr43sTaZwlmbKnS4M70hG2uW0pfRQ+C2G3FloPDqBk3HQ72WOUdbNxKzj13z1C
MdZDdGMUH9KojFRz595sA7/dWsVgabnr7AruQ7ZCBIah8ldfBNymrbIABtyu8/u7
Ji0jflNfUAEMVEK+E4SisrXbY9idkV55MN4MgauR3ZFMBPg6DOM89pENo976EC45
Yuc4WX6j2UFsh+mlpB5Hx8qfl3wnDTF95sXW/Clbjv0XREVVx7RTSKyQ2q2aLAZE
48bx7EtObBJgPKcMd7bGbErHM8sloZauF5sVJnHpt6112l3p87uHlb1rqHxl6lQB
iitEnGsGIhM8FQ3FptJ4MD20WVF6cf6mm8AtQ1Y1plqDgl/laFJ8YCPc31EZaAsi
XcaiIEIxSaf6w5rMBGddzNvSz+IJTND6tIhBUIM/pFj2IwY5zFQE7UurmUyvnjTd
IZcwRxVqSyJP51RInYWOr4hUY9Tpc/xMdVYAs7EhQhp2K2gdVPYyylosBRMtWD23
DSakKiEE/FvSxgiaGYjB0eKK2yMOfqG+pUlj7Dp6z/5TKDEeXW5v0jjGdbNn4qz/
bZBEMF4PyuxCX1D+tyRwXb8/16F3VIHsk8TK1tO0Zyd3hAOIRAC3MGbIx/UC9W2L
t3hbtPk57c6haYs8DrkzYCcxVx7hWi4a6ckalpWNb2G7aUOvMsGVrJEeJ2TeLxeh
/BLdZsu+26v6+GYHJk+WkonyY/pEzZIBlD1TkdRAZ2DOxoQfVxBP/1mHWM8/xXa8
qfJOUZ658uyfTDs++PG70HWrsE0I+br+fHHvizSki55WAH8gIJE4quksqnWL+SH8
+aOp3cxwGuF3yYIU3/UmIzNJgtB4WOW9o34OyCxO4s+gq7BfWhdkW7ZK1aLXpyJJ
XF/ah0R5HnOYYazSdATr6tWyRvXBUvvax/6yEbaBXVlGUx6JDcuGxrcF7H7JTqiw
JT9p1/ky0jgQ2bedj74JOncxfpDdTDPlfDCQBvlyOuJh6WQNapK+1XBMgNUuem5E
HcnVIzhN18GHVKXrNJ0s25EZ7S52PbPBQUrsLeprVtOYdTmNuQoeHCtRXvnvVF8t
HH3ophzbe0HVWxKxqFLtqr4EJv435t9apvdDHbX8N4SXomQw1/5nPaO7hKNuvp05
pzjfsZJRXFWQpEWB0cPlDgVvU/M/C+jjw078BBCkz2X6CXuJj1qIC5ekLnRJfsSD
6F6qDnJGiXAoYgTRJb0aJjp76HTW6DKR0I6DmUBbWushOGV0q5wSpd/M5xYCsGJB
uuUKT3FYfC5a9gXDXaE+Wx0HVBTP3dpZabAA0onMyiGf72IQxT6SlnRKqCj6o+/Y
DGqwbDNNUxqK8mZ86lxVnhSnTkNc49dsMrL3qy6j8aP1FVKiwoSgNlxGLojPdkIQ
RJM6dRIhpIvp1K7BoKokAEweEidUQ4Df1W/0tUcPrs56PCc3iqItTRk+9ildPNeL
vSzm+6GgWRnO5jeHczC/r8EfzEmbFNyhsOkRAcaU33pmh8ZIVeqgWYpI0lFW+s1F
QLVHCikuziyMu6+bo4ShpSJT2m2Zzx8j3pQKs84FXu9ncH1t9H4H8J6XCorJdYDN
fSTBGsy02CpXs7oI/iyH83t+Zg1Qb44E3X4NZB0wwRsVlWXJXBCWeOez4CvkF6pD
HKjnbXPRr1hrDHODmfMd15Je3VNCBDDSb74N0cwMsIm22bIV76YlVyEPaaYLj1qa
qYdA1+OENsupY0waE6X4cS/weXjplg5qtRiYGouxVR4UoIrBPMe69z8KekH/9B/o
m1ce04k/FszQPAu/EvxYr2WYsl0DoRv8gvxHUp921881SF8WgSqk7bzKPxLe7zBh
Slg/pbJLYqQflK6kcxxjv8C9q4/vRqP0myoZoX8jDU1dROk5GH4iG8diw5W7oLVw
qL9rkZr/lYahYsjR3+/8sysXwjTa3bAyWyQqmIEfBjo/DRgOMLsWNMraE1oTa1rF
TLZoXKzEHoi3wqXC/oKGximznVnr3ziTLd+IS/hwdqv8eGCOLdlFic+hJJTo5wrh
jD/bKNjMAQKIijKFGzksRjaz7zMN1cTfMvDtrwX/GKUm6Is5vzJFVlgvn2mqWkVX
O7V9liGWATiOiz0qP93/d4C5dpjcouWS9m0oAteVnOrNKU7PPT/x5fphm1cbczTE
`protect END_PROTECTED
