`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCtzzLVxRoE4oj4SWkmeGpTBeP1z1p0I1JZ3wu/PZMnt
vLdINdFhtzVRjhNh0N+Qd6fm3a/HrmKgxmGiw8ImP+gmT0FK/9RU4oWBOp6fBi5e
zjA933qp/r13pszz/Agb7fxmYvv1uS//5L9zEo94RGyhcdAlN5q/AYzgsb2vB0Ze
EmPy889jR5HYIU63nK17+9MECFS5Z5vkQOqkPKypm3ftzaFa+TuZV875rxaJGgvL
PhE1HkLFsOpDYfSYZq2+pjjEoVf9Ih5DxACXQaZq09MEqKKCzlyXW41SaGO4/Ff8
P5e5zGDWdTE4EE5ZsHc3jkBNRuExxmcOkiR7MXcpn0KvsLTlUDl4Y2trYGpQKiuI
SeuPnTtft5LlHmjYxPXqajpowbE2g2F3qeSz9TfA7tLzmaYZzEiB+sUf0NgSvu5C
UAgxcfeAiZMQqXK+Q3SsAw5N1tkRp0iyDM2pewvafv2ptUeh31jf75N5VltTxFsK
whWXSIH9T5GD88LEPKtZbNSJYFiN8ZTVmmT5rtwqmiKtWSjsmBdRP7UsmNGmCmaQ
bVAw82uRKs22VNbWxCI8hblgRuUiWiARDmlyRM/7ADmJDBOrnGGGZjQzq2LNvgJx
e9yCeBR8UhubCV0SNNmyB29ZhNK8QQ/2ZLWSPuG5oC183UNYtNoUImQRAZULZ/tV
GyqivkRNh+XzIN97EiNFGTldP3F1yZDOE/auzI6eSNuQXZpDFkUv/2HO6UsgJG6l
`protect END_PROTECTED
