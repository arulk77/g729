`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3ON6twM0bRyFDJLDX3TyejWf1Epm4utl/8xOJKMvO6Nm2WUVNYl8yc1OpsII65E3
9DslIW1fFkUTdJSCf6g0Og8+3h078v6mw2gXmtJ/a8oxJW6/hr3i+ITOYUJRPtpT
920QKu0gk15aGqpSYkegQbxSu6/luXlbte+8FnQE/EfvAiK6dbDMwAHZ1xTVK+AN
w3qo3+nhurb9EkgPRbobWA==
`protect END_PROTECTED
