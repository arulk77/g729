`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
LJedc2qaGPSzsleBc8MMt0f4baay23OoqrOiYh2RxHLQpgT4gx/Eff1SIu8slWgx
NIRacDyiPo4n9hwzc+xhjE7HBfOeTVplhtJoIiNnshiDbIfxGKKuXW8FHLYdvwlG
0avjpfY0dGtHPyb7CDB7dY7lTSwHDpNpZxkR1yLXtb8xEKV67/+mNkDS+1ejL1Pd
3uZRDG+Mcn7qFV0pPMU1DKlynzerMJM6iXSVqLwkL9Y=
`protect END_PROTECTED
