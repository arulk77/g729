`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
whfZdEhQhIVICrvn0VMg7i97C0YU1oBxFV9m2+yheYj7DsxyG29ThUwuOw3sQ0bT
KZJsDPokUpEiNsFt2n9gvsRQo264GUk69+mHG9ktbwRwxT+dJ2FafQufjvMDfcOR
LjqS35aiAkEHlfBzgKufqnS+t0PokI7DcVYpEJ5O2ygodDHlgq8TaGXOieOmM2hI
pzCO/V0wUWJhXJA+crVE2OItVj4DhJQTNfW4fx4gfa+WWhwRUlkhhCzffdKUBpfI
h+gzRXYBHKvCIGZfDV+g5Ee7iLr0vkRB6pes8JlY679+FEXq9v91JOiIrp2SFfjx
`protect END_PROTECTED
