`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBP0UzZLne9apBmsy6xcUZFOSWB8RBWE/mx68K2iM3qb
9LB8uCiseoSd5+I60Tm76rWBmC4gC86LhXkUIhq/6TQd3MrQbbVY/jPNtoECrcdg
r5eiG9oWt4Zv/2cgvVK8viyqiTpOT6KrFEEtCOCv64CFIssDx72mf5XX7jjHrO8Q
+3HUsJTFtMzFrzBAEknxpuCQQMJ52CreQfzUqBqWykI8P4NeGoZi8tA6cgC+e4g/
yhCkta+1PyqMZSQsTsH5ySaSz9HPGruwVqSakbw/nb5fh3KZLti61TMqK5ItPPjb
1AkfXLv6D0zn7V703zqBAnJIwa80HKKw4QejFvw308E=
`protect END_PROTECTED
