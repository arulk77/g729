`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
uXTe6H0VCzYMTmTvtbsaRRBdlWkLnY4gPPZ1C3aObPzK1nchBJI1R2USGqSnlE/U
Jtkds1DtVFSoml1vti63e7fUUBmqnP5z82coa83uSbupFv70Nf4392O6noqKlGxD
MAegAoUt3a7+GvQWHeFD6z0lxhUXvu2NCIUj0JEJ/E0Pt9nBsS8Ovhs0D+P/RCC0
0gY9UBsxyPLN/gN2IxkMFFO1hcYGHtihDh6LOJ7dWvK2EScLwHeZJ5bfvpaTBIan
2UIUVR8SURtsiLZiQfRpy3OY6PC2yOWOktpm5ypqGxgi3hGIfH3kx7+GXQDe76CK
q9jTAIcOwdRXCgU97Xk3OAlcyL8wPfhz8Z8egW09QQiPmWDpHaJicgDWTn+4ri+K
b8pAsaPEodC9kY8wFN1L8Tc6ABajPnA/Rnx0Djh+JoQ=
`protect END_PROTECTED
