`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFpRyEAV2oj2pOvY57IQhJeYDoSwrhaKmMnnmFltt0zA
Rm4ULa99BG7mA6oE5NSI9lwL9tM4C6rqk5DEGvYW4tQjGSf49zamM9MBWoVkjSqH
umT3Dfo32iXsfQeqI1WrQWI4xKXuHFx8BVShZfTHQL/SzktqPj9zE3wHmVgiP2Is
mduxkVQWC0G9Ryhm6O5IiC3sT8PhYNgD4D87EqQ47l4XAf6fwKEQOuOU1/CCuLzX
60FpofFGQWENTUtCCCRgY3cA2AciEb39MQwmLN2fHaMD2m0mjU3kqhst3WD/2/GZ
p7hiZ8yUvtWqJLRe6MXJXfUKPkqOs8zdzPI0qeVa9XRJtWDjyo1nTmbuCMYx4RoQ
dtjwoIKUz2F1nx4LhEzMS3GCuO4jO4pBKJEtSZ7cfaGfqajGGoES0Xg5GSozioHJ
dQVyWDxviI6/5hTkt4mdalaWv8HTW/yG3rZgEPJ6BWBQ9BZyz6WaG3MlGYW4CIgN
mZ+6Obf4pCunEMAxnXPtS5L8PpHl4r0eN1YtU2/voe0FK1OVWUA2EzbSIoPmA+L7
BMPht+FBH64epP63qmP5k4dOTkjL+ocMTRLq4Iy8sBHvsPwLr01fx999JYcYWoxe
PbbiJW3I8WhvJz+NoXZ/ky0OLB7sen/NBt/e8g1NHEFSzvMQ67vfhlPf2Yern7Ud
`protect END_PROTECTED
