`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKQXQXoY8O6pEYmmi0m6gEQC8i1+3EaMaTsmUdHKmBa/
0ziDvCLj/+cxk+ywwIuKiX5qTXsFm9H5IEMGquLGwZpVNAmgMI+HcIForVMgiN7u
4Q2v7Ib2mcV1mFg7ATOIcBHHYzkgaQzVaqqOiLHbA6jaMTq03nSfDioUHyQaJ5fI
OVGS7dletxsS/9owgvmQHhl39HQBWfFGbYh7O+sp6Xj81foPfLqsB1e8hg+5Z+5u
ARevUM4Vo4vzUvYH2u/e1j1343gNOuu5ugtw5Bd+u2Zsblp/KR1d2Te58C//+scA
799M4pZZrBrWiIHtZryh6PnI8ggYpWnOx0G3eHomY/n42QhpX8Scv8ViFLNRFQpO
f8Xm2dSO0W4SDOJUQWJgtRqh/ILe+NbUBAsZlrFhdk1RLt81SQW34F2+gmcQ+H8K
2XsXY7V18PcUXQQvkNVmMldQzgeRhBJKQJ9vSJHXCPmXmDmlchY6CqBQQMcn9Pw1
`protect END_PROTECTED
