`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yjToKF9OeDHq9Sld4tOkUtWuhZKJlYngm0pOhjfSTWw
kVIPzkONKLl5O6lL+aqndypckPj6zhAsDARikr/lmiZPma3LWqkUi+iYaZGBDH5b
lkiTfuzFIZf+J5S8nN/BiNSGnho7POxCwJVcU6+roSzSXBI2TO8d+ESPbBCPRoWZ
+SDqDjbIgb3XJh/1QGX7+BfW/5H5EBTQOQs1Um3b8js=
`protect END_PROTECTED
