`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJdq0M3GLFLI68sl0wk4WalBES1f/8HPXmk2udR3SC0z
cqGTSqaecYIHtFWcQ4eRms+JU5MNpS1Y9b1HM58h5i5Xwi7oG3G6TqHt2PpFkl1t
WHVmDUsQdX5xg3jwCh6VT+LRN+K6llSTVMqyMCGcb4dNpw4QeUhmZit09afxzqi6
xPlFh7Y5NVqm2LwOghfMW6LVBjsQRjmUBrlRL234iMoiAv+hTL0pYAZNsUBLRGwm
fN9uo778LDeDOOYoID8JctteQ63maSHtxXWtiJ9koEX2/ZcBy6qtuolR0IrgX1Z/
438T5rBWRZaL9ztMvEpPosJHu7/tthJ74hcLSiQQoUPjdNS7uS82WmVVzEstbND/
O3iMybaGwdBeSu7r07MtclZgy2MBw6fFDpvBn7JpL82vyziFC/unfa4tlKIFyzFo
`protect END_PROTECTED
