`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
SinINFsNSXBiw53AF8dIBn5mDXLKuhXyOs7LzcHcV8LUwVzWCr1TTYsmHi4Oyz+/
lt8AY1azyagxmbfoodIt8V7BjU4YUvGUAMWXEBS0MV26u0oeTPhQspN2AKJZo1C+
v91svHUvKXwEmcwr2O3a3tAZLNBhJ3Gfzs8RK/zCLg5ZRlXrLQxJCTSII9sLQOch
ftcjsfoBr/jBlNICYCOkWqQFq/v3G3bBG8cJbQ30dNQECQLMKrmi31KVKR4r0EPz
U7gV9WgvBupM8Cq7VScefxFcwOCAbIkBc48Mdh8x9Ly7wLESiLamO4+9/q0m4bPo
Swv5u8NEp0d5GkLSy83oMPItTH/xI0au3jTooT+teXACpHDDrQGgoXgy0n6sT/Ez
xPQb5G03uafs0dzVpNwCJvLDygjUJtySkuOLTQLeF9qzNipavDC0MM+rRXK5Qrr1
9AX9a7GOlgiYv03iGvk8qKOCnxPdj+kgf0TxljbEc31U7hWGmFcErLrdjEvbbNZT
wnfkX6PxNj8Py+gizd+VHema8rpgRyv2Odfl5BpgFloDLUP5SMSIh3gsRjyF3Kwy
mwYQcujMi5ZLU5QaD01Ndz1UdvA2FqVh6Ai/F1JJsdGHf6WNVD8MIFQL2mSc4WcX
rDE78xkBx/92DMprm+uDBuXORnDeZ2OYD6PzEN18v1ERy3vFA2ucjmMy+7ghf0WA
ftC329RtLT2EWiC8XEvIjlvE7ESeRhOq+QuDisudFXbWgcQjZ6bbr55cRlNly/dz
u3f5XXCPswWJE4tm8Z4hkiQJ8T5WOq6UaWR+wpGg9IWhLNa/OQvDRfykDNRe0gB6
Ow4fQjd3T0M0T0V8VstL3nJ7n8RnwqL/j1UDjeYwJDbGi055ZJ7yUi4xLoEQb5tT
Zu2QM8serYaN2o0IuYuBM5Dud4cLxmGElhtDHcv19xhbBsn0U//nln1HAXF+uwbM
3vUbmInfde8TE+W9c6L/bTIum5ctumvPmz7DyuP61ejGEhwovtfn4vZZdyzVuhLc
caNRrfFhF77ePDrJ4bc0o4ygd4E2NphwYzJpXfHzlvjDJJR8QAqAsH+107EQfr7f
sXvnRaYaRexB/uUr7BFEk1vebDMT4UQ98Fn+R9xotRh1wSa0iBWuLx+sgtIchzKk
fP8dcZfyyTuEWi+SzKMGN8IKZ/ZZY1XVApNTMPwBgRf/VLWtNVCpf/CFWPI9/kc4
jXLJmOeFmKYkG5TCQFTdIUXYAH2gTB4V5U3l/0RN0cYRhUV9ra4PvgBsmSDbme87
fak2Uyq9G7Bje5z2poDBeL1uPesZTltQfeFHYpV3znz6zG59QqVqp5xX5I25Kbrd
tkfrDsBVXCJMTnqh1Qj3LnJFZjEz6D5DhmPAtM7bydi5UVn03CfgdZZc2toWXBs+
iakPSIOT1Rd9zHsR/fAxFUpai1IPNL6cJSTJoM2ZfuYoMjXIBkcDu0sHvwIi/MN6
OXs6jE68CCJsHhb/8msIgigCAUfcUNZ1W5JviObLnOk0OKJOG9BfKMmU5WOFypRd
8MrNQn4npu0MgdnzvMZU8/w07xxXu6ZsfVgBpYIfdRBiqsTZjFY/oQEcD4ZVaMXq
c8ppLlTom4IIUCvjMi8eEoNnBKMZjC6N0LwZRLRLpcPscXy74u3IQQB4/EZ6lbJM
WQ0mjwfJveb+MBSry0XoA1QiKjvEynAqThHvJjg9ylLtNfYVFDPMWH7FtS1p/zck
Hor6qMMQgMDNkG0opGuoEe+UJEkbFSQ6msS7AhwivgFxlj3sFesthw6zAdg6dMnL
tv4wJGfZykHSKIi72PpnRRSGhGutsecZGULnDtnzSnUmtf6CShP5rtMzh8ND2r1y
4ThysNkwUMZa/cAXs6lL2xw+cbPc8wUERb8gL7xHeR5wRCzU35CLu7uLePKTa+eS
roKs2oUoBMOnUJZHB8TNaCvaXdtoC0sqI1nRJC2l/ufsEczWuPREXX36PMhecCaQ
vv309cKDkwK7cex+WCFkANFhGFt/3YLrx2zwzLvh7DuFq204wwAk1WdYZD0ysmw/
tIjgMeqaInEdWgKGl9ITiwvZX6DH2ognYyvDigRiD1VZb8/axnUFnR2In+U11OwV
JKdwAdd7hdwzcOypasdEtDRAgCLgjKqETFlqHzYuVSmNrldT7s0jyryRf6o2rpqL
EpxzWpGvuQCYQIg9Yeq3SslljaQ0tHH84zk63Ep1zom77QTbCvKNBIEgDG2u3hYz
vYG8VhTxfIoqHDDXOL9LwysVBcuvTv8x8dL1oHR66dhDqeO99jkFaBuXx+G1hXdo
mN2niF8h54YZ/yJv9zzycYmEsC4HCr9+e4U9hH3Nf8sT3mQKgszIA1n/gjlU+OIC
fkIYeNOi5TBYu5iIpCFLDy+VAZT4+7ssWCVExc28nbjVUyj49zgvtsWSeNAlof5D
wJHhG0m2QDjUl8kEenDyP8JaWnYKsvmiVDuPQxivKxbwpaGE1DrqrouYuWKNrsgj
zOZzqGlkootRvzRUJ17Tq8gzJ7bDJbii6tiE5vjIAi+xUgNFn+6vIQuBeHOPJseh
larEWj9VskubllPBE1Hj9SKmqYpvw8bBYEKy1SW7aTemT/Wae7swTeBajvYw4zCG
oIPgvi6UbTxH4sB3ZykQkxnDIvULsUvJ80qcFU3AyZRWJiwqF0LkMsWsW5eruwOl
B2qZzO2sy9nHal45vgJRoZOAiPXugRzmWszB6zWF065jJHwL1KUm7YD02Se8+TfR
SLNtxx1pyYxh7rHP5DVCaYO4xC2ZO8+/4NweoW3hEkYRfdaIhnHS4YzPfCpl0HyH
sbIb/hMqmdr5i9B7acCuONzPtbIwM8JFDyh9OVP7XZffF/iXf4rHj20Fa8Z4a+ym
+8B4BuaqqNxASbcBBNE4/w==
`protect END_PROTECTED
