`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
CXDo269tkFVLssJhCUcbkckc7yrjntERG86FDGxly9LOsmSLSXxEc9evwU1lQnyr
9oajgELltpVJl6QcAE+qil9iXL/dip3Cd1wjBp8l6vRY5FynimM2KFEm/42Dtuhy
rWVcbKMgwWzyfZlLMEPMKccQbAQvu46ukzsYFbeNU883VXyuAzm9mi0KMhu+OOG1
`protect END_PROTECTED
