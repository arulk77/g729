`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
leXDABmDZXJ/HGXI9vRZ4DzTGwSziGKhwnzMVPqgwH4twlOiDSo8po5uwb8Ek/hT
XVmqCjUyLupyf6S3PNo9lpnGDwUCo+r7l0UQImnNttg4jxkMsU0+eEff50w9J17a
8zoDgpuEJwor/cbnANFHpJiNbvgcxytfR7c4JVBRzFOpvK5rUZE2y8vF13OrxmRp
I6ynyS5cicikyuH75X5hkmGhvZ10v+veLiX34eSXwD5emhmmf9EGc9EfsJ3paiON
hZtwdTnMlhOC/db5NpfbzNdJR6fR51PG/Fy6T+HuiUnr3+6I8bhEMdYnbPHcTqws
3dgb1AVFQ8H1FdOHalDUj9cfHGmIX7IVbS4XWgswHnUfoNFoxjzTzVLm6UeTVRp2
7oQ7jI0fiXDE53ALYMtKhmX5Vn8UfPy6olhBOHl2TFu+5aFTCwvRMBKSBj5lxFYt
RGI9ebADo8NxSqzgMg7T9GgUyQEy7mT9oVx/IwVSHo/TqFJf8k1qYcIbs/O3Karl
V9azZ+ckLwRRDt1+in4sztwNnsnBWznSqbTfbfawdcaEFr+E8zvmqOTfoDUNMyFE
GOMJOwT6vUPz3Vj+lr4avLshPH/Zx11WcYbCLg5TyW69oTdMS7BAZtfZ8RKRMmF3
6kZJJ0T2CgTpTXXgy3xsaRRbWz/3NSvWZwL6pwKmZ8B+59KA2olshoGarkNT8ayz
9LvFGFCJHfVzGpr3ds8Bs1zmSzz/GT2OAS5e1OFAnhTRVSGaNexv3gNOfgMZC/N3
KBPWUeQmJV+gh5VnunjsxIO7PXMxiAYZ6eldwU5aFtA=
`protect END_PROTECTED
