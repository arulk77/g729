`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43eIaNc/tTOXGpMnXqzI3h5pRdn837Rrwr7Ko3x5iqnp
9DcnCqx659o5AsC1xA+/+kvcPckdPqajxVkoOg31ftcJ3ax8OHnZyo8vXZRxzr0O
9+53PkzYGbwFoGQGYeUSxMNsQstBt180KhbPp6vKDPvlLLBS5EMZwzDH3C817mEr
fVDfQL76ngRJ3T0yzVbYWjXtWDS9bOvduNpJ9YMjU3R/ILobQ7qnFh4nSkEYB7Ti
cOT9MP7dIGswe6MSqn3jZP8gggRQKfKHQpZLguOlTF6mViBA9LwuZsXHwFTB3z7+
Vd7uWPT6PtMle8YKXCO4Gw==
`protect END_PROTECTED
