`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aTep/9jaPM+ExW1NVpViGZ5dp1TiRj1h0z1wnWBB9IziZmWSMV7oyKzSsUhAsKc6
rB4LpQ1kUVs8fgqpIQVkVDrtIof/1kD4h/Yi7V9Ym53oJyWw4jbmai18ZtwodA0E
n1N+XXnB54fTWbNojvw6KdEyzioN345AldU3BvrqvtXyV3zaHH+H/LVmaSP8inL6
QtuRm2n/t7l59zfQ5p4uHpUgYT9OOQwd4ogcw14KxUiJMFHugJ1d6Cgr6Yk4rHYV
L+BIL21snJaljr8TIwgBE0NpAzwOw3eVBMv007W5QjP2JTtCx4W1crn4IbDcLHOd
deN6YqVTWKLOAoA8r08fTrqy9dO9yVzn+AB8Z+erQWPaZVzSUuHb3L9a82Kxfq+G
E23mwGt3qR4Gn9YE3RvXX3V2WuyC1Tu2qPhMyD+RA+OcNjQTEzpbWRwHu1il5Xfd
1ZQKzGRdgOvsHlry0JS3wfDH3SNr7Y4OMZb/iUiYfC1AGne9qAvOw5wnY8sZ+uM8
Vaq1FwcaFG6Mdb1TttYH27jb1E3KJkN5mGJPhgOEAuAksgJjVJrpc9sLHyw/B5QD
fmYog676rJl2nODpatESsRtbrrSd89Gst/+vVP1CAA9rLnhVuEQk3LoNip8KRIlr
qk23VDCPz8MhkKil8cseRRuhqiQ1lE1a+g+J1c58VZdU2v2WVEPARsBetknSkQSX
G02LedoMS0Vfd3o+t7ekLUJvg4xPHYFTZhJ2pacxLwe+DSp7XHzLtQ84dAFI/K25
k4+acRgGMpk9UdTSLv7D19LeJQHmnoyftqXo6m4WfugVBX6bEKBEXltjM+nlqUAz
54RmWlK5icl4BDcLdeDijU5WCj+jAz3gt0XW/4yW5OzogH2uQRU98sBoPGtWuQ+Q
7wiywbwhxufdntkg+ikuTquPmUzOZm8E8Eo7l9bxClkH/IKI7BBaqja5avhcbZy6
5/Ci6kplPcf3au7ciRynbxiNdyz2LTeZgdBARRZPJD8yS1BmOSlIPlkmgJ0dgMdq
sM8ZI4pbDLJpIxYovAdtwz5g7gw4IVfdVoi2LodKVBv74tZs1v6Rm3vFAFVEh6is
6lkIh1FKzh2Exbsp+HyZ4jq8QkCfxcs5mFU91P0HeLEjNNSJPZgGilyicZTbaJBo
RysnY0cKa9vSaGeOLnuW/yu12lx9Z0stgon3xyjIjoABYV6mwQ9RlGPwqBtdF8v2
3Tgpxy+qvT6pToGUJPamYmyRxAgkPRtdo9Y6dOqKfYXKmGxom2RZO4+wjoeObErB
0IL28TMifEW/hKC6hY8nE6ce3RWOdFma3RQyGJqxkq+t+9rxFZhsGGxM6hrE0uIL
xaJCGjSVyVySs0b08WHrlWDTaiUXpURo7/X3tYMuZm3BNlkB3WJSeC61KrzI0GQ5
XFy9DMo6ncXTXlVk6f/NkfQyp7USccxndq1niNHp0JHijc4eBhPMdrtRi7g9u9cw
OJ2weszeywvuguX8ud5ds0bERCmAV2gpLjGby6NBA45GN5S/CRs7y5MxtzzrM5IL
zPJQmaUzDTDtlTRirFM+wVJSaCCJyGikhiDFpTnEZRcf3RGueFHiAIkGu9Vg87hd
NQvVxCDwr+onshlb4mLxVhYtJSTpiALv62zf772DgPzkCMhPMLyKTVxsNED8bDDT
n2v3KM7M3lDm6YutLio1PEzyDyyVEeOxUox0Pzapaz6NP4bXsCQx9wXvzwN4XHgu
vbeUVvLRLs4YwwS5GlaZFdfWtrwKGxZl+TCIK66JxhYvTzXo5UORlI4NjeZUOKUZ
`protect END_PROTECTED
