`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNvRrAdPVQ0y72i5CgIHOLFyvHNC+0zIzG0/GQb8xbcS
yzKPGqPYk7ogaFVlVKh6cUA7BSwg/wzjcQG6IePsNzC78roXY4o/pRlzgU0TKh0H
TY0CGfrZTKY8wwOG86qLmbbd8ekGVvJl4yT27+2L8k7O5SESNGcKde9WGHxCWKX6
peAn6Ry0/204gI9k2g5Z+koE89wnOrjkB56I9mC/wLi51HAf1nRCTlQLOUF+IvBM
xRiTLOlj26bt7KF0jEsagcCYYupVEihT4Fg0Q6LOp0B6RXqoBy2Cf1Q/lrZgXYiK
tTOQ4oSHpSH/Lj9q53MqcH+03BwA4tIxksF2Ibmplvh6Vz433YmJ37oNcZULUYyi
Nmbodmzvn0DNMq/GltRs+YftvVUSJbEq6BGn/uIfsHRmzKu0smC4o0TCSwuvxYGv
56XgLkY/a/yJQmYi9vbpQ6H2SU3eUsxfhzPF9+n1GkFLZ9AQaZfsrlr216GC0HfY
2J5dWgqYlt0kOl56GvHoR1XNjmTZmqUXAzSCbcR1utINlNyW6Wjjd0mPgQ92tOZR
3UHwhczZXlKSXOjcCm7pItFEcxbMw/JkecrzFHlkbf2tgKBMXRpWb2eB+yX24zyR
27VIdN7KphIqIY/QvcfDCwF67iN1RPoZxvuujpWdysJP5s5jpZFO2OvX9yZ+B6op
fQTxTiuXcfBG2n3GQRGt/l97mQVL7M1JAYlRYiXYjksc8/lp++8Nmy548uYT9PfS
RXIPawSxTmPPciLI/tcBmaoiHx1RtMRbbsx7JhL6ISUlLBxId40t0ZRQ1xB50k/H
/vsJMUELYkaJqjxy+NLC2xNwiTObgGcocdJLNaAbDQvVqaqDjsaTjkg0EFmfLd9U
aBDjdkLG4MtjiXcz0cz+YYMXkDQds3e/nz40HiN6Htq6ajjFTrOp+ImcuTSIp10Y
W8cif37vRG6u+6Rr2dPyCcKGKcz1XJDbim50bjHIYee3fMou2GoRV1JuIjMrkmpL
JXykXb64N4gRgKssDno2P+MWJgUKOWsEk5o3m/lmyDbe3ht9Jk4fYy5w0VMZHOuT
o3DbLClZpaPvxaIqRTKz98vqaZpSKO1en7duWD2DDzQ=
`protect END_PROTECTED
