`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C4pAT1w+HBMMYj7nQ41Y8zE2oFMVhleAPSVClucketqs
PSmgXoClnf6LBclO/P4HE/p+0TxvbrgmALeNkIP+9UqYSQZnYcFRaChEH6avW3qa
WKq3HFSwu5KQw2tDPXhdKK9NrgBKTU0uZGqRr6ORYkpPW0xOuDdedmO2uh/kq6XC
1eB85VfvwprMak5g2Eex99pUiFC2jBgyyuSayO2EBmtoQZyWAytGsYfksB3w9Z38
90WPdviadn6cw/Y3VFx4U1DFdLB6DRmjdaNCv4D8JrUGf0Akw0srT6K01qZdPjn5
+nyzy+1iWLQNvH2jQe/1iwD+wm2XxxjKsIvvkDe03KnN6BYU7ndDG6fHfdSsTOXe
iJp//4nMWWVB/kCZscHKZCGLu6lfMzG/jGutdo5veggg4Zz1X1XgD2af2WNPHdrc
cT5fbdp0waV0g5gPq5Z+OA7jeVois6ZjGMwcv6F3f0/ISmKfuIuDnp9K5+I6eDgY
A8OmCMKxqFb9oif9az5wvAQwI1TisBnAWblXaSej8pSRPmE/mmdgFVEY9DEoVXU8
v+k3+y/wjuviiP+z6RZNnNDyZIZiTIpP1cQPdEu2ARVvX0zltdTb5/GfZY8SUPnS
g0YBIjRfSeYSZuImJKuEiFCrsTOwSZiDRQ5pDzYNB7aOTHWSezYKQctmsvIDYYwG
NeaSiIZ2kMEfKqxnp999PAgojQ/gF5zE+jz7Av7egmo2g8JxvbdvJhNyfrCIRjYe
fq2Jz04XF0GXYMMnBNiMymYtzpeCH9EKklNvIjwOSlFuQtcwPS6ZgtIu137g2s52
BhOTWx5HHpR5aPJw/oEfj8iSMRFNQzBVL9nOC/A7SMlPx9imePSlfzrqCVMQ+Jkd
ax2hz8SHM1TU9ZF6dpXRFsnCtG1cG7xdWk85KC2njxYg/F04CenVGnjMNrXCTy8Q
3BJRhHf36q/YCcJHcwY7qApVRV5VeTZjzbdKUWZ/FxpEbI0tR9p/ekqcKBe188pl
EPQq6ntKiGlbeHz+MkqyThuh1HxcUbiO+LccjUSRX0SLX8Rb7UR57ccMmd78CSRM
ZbJX82Ozgi263ukDfUWkpCjqJWTDNykR19gSzJHrL4HsJg7rA0GLDmd10QTQp3DL
X2EXWIaQ4gxddZFVyiBMnnb200MttZ0PmS1fn6VkLtqJtVig+WDQje1Yxbh/Z3+u
VKr5ngERSnO6xDDA1e5iHW4CTy7hAO3uasCH3BJ1Yut9V/aahHhlemo/VABixlza
GbouD8Mz+scRocEHv5BFspZr2YCtZ8G3vnXjzDKVarpdHTkAxyna2Y0GOuiTCXHN
SKImQwXJD81wTWowFkjPkg==
`protect END_PROTECTED
