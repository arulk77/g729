`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
fc0s3FUIISgqzsIPA1gu7hS1b6BZt6dqVnXmPv+QB83MC2Q3VnbNeEYWaTC/z+0L
yRM3JlbJhkETbHeZC5smg3r+qPzY/JYAcABB6j+82/fLWR5oVGA/8m1Up9wDrHGL
dFWwjmbsj8Pxe4jCJZ3biVtd0rLMK26CJTEZ7rXW2dgUG+Juv8W+bbVlcVLEzFfQ
cfLzkdbpRCemRYc2LOK5fkHdG/zl7kqFnwZHCurpI2b3ThZvSs2yasBiSuMXr7vM
WJkUIbm777k7Fy4qw7eSnKANwn1p0MOhRWxj93bawsLHJf01rXvNtV79R1D3/zkj
Gi3H5abqWJY/SgY7Ooc+oXqVsuYjnIxIWiCvLGytOY1QCB55kGoUMOigNCEokTn3
qhxFe8T3w09C8xIwGoq4G45g9O/umfInpClf27zvTkh0czfA4AzpuVrcuZpSMvwp
GE45khmupbGzSbx6VGy8gm1Udm3XWKPa52lCXk7JbHI=
`protect END_PROTECTED
