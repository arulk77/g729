`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IogVMB2523KhChFdH7TMNqbq0h4gF9C5nKiIS665CkDiHEIOhlywGeCB5Qyks1HF
fRLnyt2cv3bLqIKQN0Zlkl2AB1IUfflirgXzciJ73HXvx36T+HfMVMeJQAHoQMVh
b3xyvyKhYHEk9ECtlAieWpeIp8XYklP8AT8oMzZYZMB0sEi7VT2/Fqp8i7gJVhbe
8VKWyPHNP+GTuO1Vb94JGKS34fqNqPu1Kmh++jVfrHMgslzAX8+uuJ94IksZm5s/
6q1gtJaCMf2R5p0nJF3IIn01o/fp44JEqKJZgQXzXb8B3le82N4TmmTg1gE3UoJi
BCXDKS8s9Sw8tMpNQHuyrSRahjfG+BLOmp42/655w18uX1Q68B+e9DlEOAwzUYHj
zFuL7ajDFLWy+rhQJj2rwfH5fa6QvdvWixZvXprSarCrP0X5s1kdsQVVgADSmLY8
i71jWA8Vmxa16zh1vFgqwelBYfiUaQIlAgE2Qwdd/Ze0zfYg+y+m2isNo1edtzKL
jhUkSlXwRzBh8ji6zSYajYddz6jGqfELQFAIvHA1imLuWhu7OfPgaTXxu6S3mg1U
Xld8E+pFtBRTQ5xbyxg+gAl7/kdMc6P8PRJ7RRRAhDIJ5bJiW0a2y6j/RWj0fxyE
HZ/hGxLZk5L+l0erGYTP4xNbbjJPmayGWFFzGtk9wH6W2fsgQTRPfUNTUU3P6FFm
S43FqrNZH9kg6Fe1JXuHxVqI40gki2hWQ7h24WQzrs3R6KU5VYrYgP2ZSpe891Pr
ngqujhw2riCVMD1Pb+bmfCRTHt1r4X5xthgxxHvUl+NDAWBkjrMP9ycAlWWb/KKz
KfTHU5m4dG27yfexiZ48Zivwuu6WTFUcDsnVQ6iMVLttZuaH/CHBYtY+RQss7uMr
JU86h6OOUGpeatGAi0T/A6yS7e6mvcOYLt/rd5/HaPYy2eXa3scQPYKVbPr62I4T
p+o2fApllIvksJZJ261MlUUL+XHsQRt7775RxrJmbnFLXCkEooPr5JEVlwoKweHK
+8dFg1DgQEg3AWEm5sPJHeVGQGVZGN+P8hZK39tQwXhmAMEZH0uex+Y5tTy0UZYp
X7NB3E6c56quJqdpfQofFvMkjJ3aJbv1twEd5KxFV0w+fdBe6S0RCm0fKToqVSCw
3LdUhsZ/0R0oQLMthn/txSpB7ufgVrHud2drusimLMCBb8QC+JzqilOIXLL+lo6A
ZR8Mv4lSoVHcpMfJSgKzjxeEySBRX3C7JxvcYTmwHIkAY77Irz5rGwoqASsStque
RfLlxeEb3AcZLQitFa6V3nOms9YhayygBkz2XgpQfnLr7jQw0wcbeQs+lRpmjVLY
Bmq5JEhDHaCUkExP1YXWgQ2XqQCpf6sg2HZ/JwpJcGHxf8RKde8UflszfGVEVkAA
ZjYgl7PC79ktOb5iVdpI6Vbh2e9SM2hwB4gjEU27/hH4+3WcbjoaQA4bKlelNkvO
6nKz7wdXi1EqUg2fUi1sx5kzdHI/T+1jito+U1an8ZXQo9ZE8WYoJwV1wIB9WTMP
LiaPs935vLtlyZy36kCEUQtp2u8ZEpVgF6/YFgac5kk9QPHkGPkEvCxyJ1cfBHpR
g5b9iOUECHEBh1T2KCR1O383/tkxD/t/FEznvTG9QsmpVfjBe7GDvpT1ye6ksB47
`protect END_PROTECTED
