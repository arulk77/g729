`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePPzbTa4JtAzwRz4FoEEdiAyzE0apkBmLSDNhctoQJeh
MxpTbR5IgrLLCCoRtFU5iD5lBe0qfbBoR4bbyopfYR0TrBzyuPNhKBKSnENajZ0I
+08QTqVtT6M5+QS9C0gazKXNF5LNyi54USl5kx1Q5CA3SRnbClhdSXRE2gAQgdZ3
i12kMVV375f7CImuhQFwuOpi32pLcGQDB/HWrL89cQVXuGw4Q+7nIp1YYHdR4m1r
eHSWnrIYA4iA59/BWFwWzYSUZjSCyhb0NlLlQvIC5rT5DEKIzeOE2WcQlJJYeJXP
hPSLCZECxxjfR1F+AtuVExRLfk3lH4+x/cF6F7RT5lfOv6tZj7lxMU/ncjG1OuvN
gQBXJQdN9BJnNYGcLy6VGwRA7XurhkNFCjlH6p887oHfASys5pRa0g/sKPhNOwXl
LG0K+ZXgDwxKrfS7yqEFLqcao08skHJoIys/c0yXBYhAnJBQY27jHnZ3NBkswvhV
v4h7Ct2D/wV/m4MsTRi/YEDceFeLksB6jH1pPPe2DzGIGNLXRULduEFvHsK38UI3
wigwiFKascYgBS05t/JcQEazb8d0i3a6gu9sNnBvJSksjqkE9z5Jp5BvJg0rG+KS
xI8vY/iPVYtMFzwfQo4DAbfUnjSUYoVNaWBcV/NXyxhuGZ58TPw4jjfav1pNymlT
ea38bfSKaD8CNkyRTz3lKPhMZNYb+I47HCiHMglPyzs803zdlHo/eTOAa3+xKjIn
4Ypzj90KV3sO3G0Z27aAhmD4O/2B+8jl3oFtgxkU0+atZX7jtlWVjziOZ082iAi5
rTWHrOhOzlfYxtO7xFycS3ag8dxfYB32ghogon5/wTdJNhJCaCB2xUdmQqTJZCRT
awRz1D6OSD/dP4b6Ia2gDy6T6lEwj9ZEvFdtubAcsKbk8qAicjC/OduSs+lpkJMn
ItnwsW8otDMmuRB7jOwecwBP/Y5dCmpnvz4klNK98BQsh3LFEO5LQXnI6YHw7RUN
O/PuaClpkCKPoTW7at6Ixt3hX30g7hTaQIZrYsAJalMQlBidTTm+KgZmscT5Tgau
S9z0dXVNjdkIJt5VFShJUiUIst9uOa/ZxkzgO4BWlJtB0WNCGUkPxyx6o5mlucL4
kif2MNGMmDhXHyk3b/8p2+U29yMAgmdHPw53LQC5MmW13oPUby5TApFW66TmdrN4
PB0CoqBKummyBENZF3EH3wItlinUlUFoAsg5RiTPg6qDPJ/YAZFQDEo723WRQqrt
6DNF/xdyFZm5aFqRRhgSUCAadrKsVz88+9nh7Wxv28yEbdarJYIV8qnJipzy2x6u
rx8iRStTrarR0uf5t1UoYJCDCuSlmRDGlVBRkOgJUxLh04O5ylO8jatnFIsdGwS+
aIOhoswJ84d7EsBFydvrRPmQZkZ+L8UrUMGj3kJ6jTEVNGIWX7h6WNS0XDNav/wb
urCzYj1rYP7pbaAoyLRgyA0qOB62kgBVtJ5TdISEjJBwZSGlFQdbrK7K6B7BvAnz
z14YmNs/rQXPjNZCEvRwYz46irFIrLVKrS96aUZDnRWRXNnFRGtSaRRIDEy5F858
4GojDRTD1Jtccb0wQWToWU8t5ntt8RejsZ3G1xy7IuiUe6+EsXzBdnCmBVREKwJW
JHuXTLdiiuvA6HLj3H2ubp/nTwTtPrKTcArLyaDXo3Ip+WkMIeGRpc/mj5XErNpl
zJ9zhta58k+aCkpHA15ogu3i3qCewBoMWXTnGSN6QBCJx4T38HmGqGp3kWFGPcpU
0dvQY+ibcklK0jW5uF5a23RRT6/Lm9W5ajm0OklW0BoFz0GJmXRM+BejHn1MSYub
qDOVETp13a2Wp0SR+kdYxhLYiXr/wizgvDh5Vs0/C0hOKpoIuJ2eL7mxbl5/5WxA
KZbwqdLszmiD1mFbEzCCRZSiyKGUTljRklRfZTnE4Lx7+aow/eXcRqQlkhfYCNfw
2ch6Auye9t5M4vXcz1R7XrQpEDoK4zLHWVwBYcbfbrS8XGUKuQu0Z3WtjYDHtUrU
PemVzz7k895hGpNqhYJBmZ3cRNYrgrtQA2uGo7hp5A9Scg9XsQ0in7/EYfFC9K65
5jS34fkZIikaX3PFdyMKXrH0aYVAcR16bECi0V9bhLttKoRDaduy+jc4egkNeJ9R
r/8xhJ9+8lMYZ03VYXE1jGC/OwShNSQ+E2erwhF1X/DfpUmc/cLRbbrhkfmVtw14
TnCS7EZAZBoBCtJ6qF7gGIS962W1JxogHgnuf1U7Gol1FWJWcFYgQagQ2Pyu27Co
CeNts3goG0OQBOBMC5fdO35tvrvayveZA1KMlQuuoDDO/SgfzUcIXmwARx525dFe
RuKueenUe91bQ0cljCXv18iIsYrpXqRuQVBeO7knvOZlTDHw4AzaRsbcZZ4d4QVb
HKqa1XG++Vnb/4lg+wFjSuqvyrnfE2QfpHVeb1bh4udUXIm50T+tPHdQLOoOK7eQ
oRyBo4KQE7cgfcE2hLntClODHXy8rVlFMyJA9R9nnxYi2TO43/K3Z6zGBmSPZtVh
mhw486Hf2nM3CAx1lEqbMLPkLqZMndNWysGd9XlTX6zqj91s02MeLZHodz2cZhs8
hNXHmEBpxPjCtdu21svPnJz59f8rdlyJMItNd15raKrdQM7eJJrDwT50Bk0L+Vxr
iff6rX5TglVoMBPxs3zrET/MOZDY2y5bw9cDRmokD6xI3M7yD3s0w11z/aC0l9o0
18eeKaZ16oNpaD+XPnCbroqPEVMSRIbuQBGZ9keVpJ+McbaNgEAYbEFd4Y4Ma04F
pT3Yodpn7nFmkaVzSAUefv9uKvliZiNDDEKNPNeTlEsmPig3ozx7U9WpOh2rgdYg
7nSQ8hFmde8jdxllQrjJU+o+dXTMiSFZ0aaLDfpaZR26j/A5kJ/V8B8XSWryWpJo
sK1PEOcP3ACfsQ1QrdyjVLyZAnaKNr4h1/uvQ0Ccxj+XY2NlCF2dGFp7sa7WA3/B
ce1bdPbsnkZEh5NyqFN15gCAVoFVf0+ebYuzoLmJhUSnqQE62rMAfC5Sr68A58hJ
Pdh6sdIs5Kh4L8WFGSc5vok0jGRJ1CwWx+3C9lyunHZYOuIfmXkMumoDBDTqlmV2
m0J4dZhJZF6xe0Nmg12jSdjr0XAVeuPbVARHM0UVDgtM7+9dngqJjmk5ZwZKAM7f
F9Cvq91TBXlOym5zXaQK47xArPrZcXB1oYn0+vRlPWj/xpxXVZeqY+ZJCNJlDEMy
Jegd7bi0C7dmsQ+KEHcM3cT5JEAdJIvOeTyKuyl9QJRvGNRzvC+Gj1UIi74mgv4E
P/V38acd8+cVMUJ9Mv7NWZvnGOwF8U17hgKhealFI7HeMBsks8cYoHl5xi6i51as
VYffC0FUO2KquODSixU8Y7sV+Fd5DPMyH95TX3Ms3IQbkvY3Hd8gfrnomcRZZWjC
ERRy0yg480MLeUcCm1iZYA6I9dDQCy5i3sMIeeKrY2ZriSfnH4Q9ro9qEQXbNf8l
VdQLRqBZcvxRpeNDHOQeq7yQ/52iG7SwUDV9P8GIOQg=
`protect END_PROTECTED
