`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI2Wx7OSRCMdMQHg5Nqv3sAjZ4NagMPmFVG3U/XVlGjj
W4GHtGdZzd5MQbJ1MuYQ/YawTA1gCVAhywmnuDN+9qgm7H4NJeYUKVMyR7A8np+z
taaQn4kRuodmBnewcGIypg==
`protect END_PROTECTED
