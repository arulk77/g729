`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JKebFQ1hddqfKTEvefmayfwK8EWY2G7+gN+iamw3/EXHJ32ptu1T7H989TN6j2/d
Yqt3SrLVvcgRuQQlizoRGefA7Jt3NRafVLkuzy55L9jY6cv4wBqHGxrZIiukDHPI
A8LzqWDx+asCgtlFeUzFdmM3Y6Fyy5Al0k8CTcn6wvDLPhlYVl0cSKNypBLPmVMf
`protect END_PROTECTED
