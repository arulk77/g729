`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEc9PnVrHY6DWApVy82wpoPxP/WC3bftHoCXZ5rgQsF3
xnHLOn993t8uYxjXG2korA3jQyQJiqtsg6fJbDbx7dpUOrTQ4WE2D7Eab6QfSggM
h163aXO5+jUWye8uETSmVokTR+VE6ajIN6FRNFr8ud0g+reTTEdBnCfl+xHc69Bl
VZU5ezR5NLMjIeYSCMiWHe92mxLZYUj1WIH8tKThycNX8AGrKiOg/ELiumEjGiwd
SvCxhIY4x2EyJc/xMwVXKCt4tjI9Vzerfrgmpah7vHb5b8p6hkRHPuw0nPIHbZUk
Hd0exbRddTA9gw6ueGekcgG26epgHdq+UrjKQkWvcKcHkXuUAV2dF6WCMfzNh6ek
tvHptJd2Ta42dpZZyssbu4TXK9P5LEFLtSnepGaEYtimrbBbWvB8waVRpTBlWea4
FdbpnuS3Kobf8u0UC8Fa/oLrDbK/fmXA/lTRU1OZvGhC7A8MIy5+IskUAa16D6bS
`protect END_PROTECTED
