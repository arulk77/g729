`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SdwWJyaHCfLu7TGz2BkH26BZAhsjYtukqpy8aymDXleH
hxowuWg1nKgDNlEqWeHffw90mikso8TslVNvGKcxnhxWp6H/hzOdmKBZfjNKiiRp
sBg4CZ7I1NYV3AM8ssxy3RNM+0rdeTNIj3kZNtOYELiDkRgKRlq1D2Qd5P0+a/dI
ZRoUdQH9XW1hsXVJtsU+8AvVCEegatz7QUiOYoRzsLEJaVUVph7MrKryg0zJcvs1
AHckfEpLwUuo9KJPJEn6Lz+frWpbSJGy7C4Jo5X0LjaPeRtADdKJqgTfUco64pH/
BzcKMchYZtcvgnezkYf7NSbvOklNprKMwo7t+nvLCEYDis7qzClkm8XWTBs4YlRu
uxgl2KYCemwGmSS7o1eJLjGJPybOuFYDvMoW0F9B2sI=
`protect END_PROTECTED
