`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkbNuODd8x3Yfj1IyDJAB04+Iq20R/ZZ2nue20p7erxq3
Wsr/DFOPfP4P87K58B5pNheCDmq+qYU1n2OjvZooe8VXHzXCYXSMX44AOgod0g46
B8Wna8DUifaIo7cYEFl/WhWIqoSk5zMOq4b10uMixx/BDDfRnTULf/jY4oewW9cI
wVDbyM0m3Xk0VybO2FPy2dvY6tWTuykrFA/FpnTHT8k0ehlQtOYSdacuxvQW2GTr
LBmNyAV7izLimDk77PdKKA3EttXNRoJP0CLXkV+gjWA=
`protect END_PROTECTED
