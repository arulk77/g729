`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48kIJlUBuQqmAxXRt281Ypzwl5dLt+4ZtODQek3BFFbf
iNuSW7/K6LmyWWUJ/dolQ4In9VfHoxNLYwK7S74+6gZcEFfAYwwxsF5h1wQIfMwl
lTfW+crDIRIMGVdjSwrdNc/q4zBd6hzc5wqFw8Ps0JJl4V4AZvQUG4LEyNXObjIj
xX+l2ANWbehDaCgJvQhNdGlO1Nze4N2/NffNwhGpECY=
`protect END_PROTECTED
