`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN3Z//pzulp8W76d5WU4u7pEceGgFYvQgtPbPcqM5gTaq
YQUplYAiimZPZZX4BDms6qyEqsyqYNOeQjIhOR7xN7YsY0K+IP7J0m/ddHYfv3V4
ynIK2B0YtAJL6UCao9EXjh2nD9KPf5we+rHZmM+1zUgbz8XGwsD7dilXOH59c4o1
0ho5vZm8ImIweGFxHRYBaS74VWjSGmtfFpJRyDoPMiXnU3FC8jeDLtJyMVgUTuCo
ZlgtyMTFDUbFlc57mE6N3ixUdCKjBQbQVCdBEvhFvY/q890mauR3/c0D4vOEMlne
PVqEn7H9tek0d9N1EHsrIIlcp5JvIelGA6y2JA1H8NuyaOGYryxG7psVbi1Hj3PU
cwnhlR9c3k+TGUJkLXSPsF4QKqjKiBahjvwOM7yPBnpAYMHCvA5TP9ySlYRgv+fA
rgCkT2EeyQ1Nsc/GeV5FLA0KDtHUMIx9REh7K0RbeOKwDe+Pa2lk2CBd3yKyikbo
fQ56POtN3Rm26SLfjV/F1cfm7PUtA7RLjgdXgbRcDAm7SR77C7irBb2A/3AARgqY
A9uS7N2dl0jt8rkJGrJbSnC+66SMp/ko/V2tsf4UxLRSCe1Iqh7O4ulRCe9pZwpJ
OAstirWbjV0ZL1WCg4/cm+3Vl+ENGfAt+USkobGsm3w2VW3cDwabMXCqk0RB4aC/
eCX55NmEjgxWNFKctveHYVMsXVTRDGjiGdQumWhV2/7LFSJhibSYTz1byCXR+iLd
FEy3KCN3Ps88wGzfG/FrrQexiB0YZNUf8NLUx8DDWrptVNTz5PoAE2SOSgIJ+R73
J6/zc+5Zz2pOuyNJBigaOMQB95q9Xk4CdeCMYJYz0GSHjdqWRDUI9YDgBt+tT4kZ
x027xKD2uE6DEPeS/cHTycIhbhV/TxJr3BaQDSTV0A3lnphWDKX1/kmmrAgqpYJs
AvawyMqv3TlIryaJT+1W/nSUpo+jbCNrfVj5GVQymWtD1tdEYAlFtEfNt1AFdlKs
YuepvEXt4fdM+5YxQrgskUJlDrXr5PiwfToF57JHtX+6jDpAmcoateKiPg2hl34e
JUZQs+uw42DHxEq+TZv7kliP9MVe8ZlR900EJSnpX6A+Il+ulxEihSBTEj3DVptI
ICiA1RB6ddw66Iv8FsrwIkIcaqYBzh8T+ffACfJH8CSAj8uMTYIIP/BA5GqyrObq
yn2W2e/SXImWcIWKWrzZIq+X1lD9ezRd5cMQZPk/+J3NW3Tz5K3fNuZGel1AGmJB
A+SSrE2XaQ1QW7Sp4+7gTERxZMeY7pVm+WsZK3QL0kcDOa/cS40YMOLwIeyqNyNP
RSIIr0cv2U3m3LQYXsXF8qKPnex6xdUavDVjNPi0U87HqnoCH+m6Pa/tLdFIoqGQ
YCcn9rSpV+1OaImDoZ/H5Fe3rRNrBgyYQG5ReaCe6+c8LUhP1L6VacKujnFv/cVQ
wVzEaNe6iwo7R+L/4KHFooBaE1SZRwRk+mc24RgogJVgIMS+K7FhIdv1QVkdryp7
PlA+m3oXRz/D362079dJdSJ1Rt3lYLhNMNR3abzoN9+oI/h3dtaKFv5Zalw34yUr
rwqPrMUk9LL5uBByvG6M6eEsdaKRj6eX41GugC/BefQFU4wRUbDIioM17c3EnHrN
ngAJfUxbMpcOhaeeUr0mx4XR69p4HgtbbpzTjtB4zZD8H8pCRNdvVT5NE19y8G5b
i6MU4uq/7D3ckMhxt3YMJ4yDfeSeXOC86BWdxpPWl89hxyoNKEE1UwOWxjmSSoFg
nZpAlQQh1bmJDcWH/3+uk1Bdtc3mf3ooMJSp+9MF3ONgTDzB5R1ZfBbLjYhFmKcD
cczKEtAxNSkZvpoqHvQmRjrFn0o6S8FWf3z5b8IyFhUR+gjZPDya3J3N3QmLt0fp
yCln/Eqj0hvRG2vqE422eRcBARk4h+IDQR8KaZ37GDg=
`protect END_PROTECTED
