`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
z1k/VB06jUBveslohKXIvlr+VnQN5VuGUyR2qw1vr8vWtcwc+HS8ldc7irjCNCE9
Lj6dvc9HXASMCriff4eETMcGNcNeaH7WSqW5lpXBUEzXaYB/o3B0YB1E20YvnJqY
REVYQJJ9VvoF0GIe7DI97EDINZ5vwLRbIKpZV0muInKGn/2OlzHJt1jxh2D05BDs
mr/oeBq5rRo+24AWKmSPq6JO7FvqsChHX0YHbYdRCMC28DIxmXf6QBPaW/d0Z2zN
AiG1GhE0Um3VMkT7XryZCze8jTL8OJOerCR70mxTGnMQM08jpk4Zvjc6zbO3+Yxb
GS6beOoWajtdgXZD/H86f8cOo//D1QV20zxCyfRdBHRImPpVMvYJitq5vkWtjRXu
mSVOIiiwlf+f5BORq6AqhB6jXT+VEliWf780uQveyDfPfi4ogVMtDZrM4dsK63rM
9xhj3tLWGX/TMdPKTmmXi+VhvQ7xeOutqCInyXDc+UoYpwdJMSMNEHRk+QfESfPX
SR0s9SbsIODYgxX+Qmprr5XnR+KmTVg2Ag49SFM9fbdDX4ochu4SgskSA74r9B30
Z97JH/+sCd5dOD7WbmQ6+SlftUMWcCLm1aWimDh/xdQwnsT0z/cMFTwYmZmVfBLa
xU8zK17h/pY8C3WmQDMyejyE7HGOga++3M2cS4/tDJJa50v4/zIlGxIV6lHCk99t
90WiE8pBi/G9LnEGIBlu+fMbQgWdjHWpPBH8dUQWsTGAdngsqWn/NQmQ4dE0eLiQ
yBxS5y2zZtD6eIojOsQ3qXpMn6WZjsAw6dqCQqwn+vrBgRzB1VHeStwL/E23D/kZ
IkUEwpRYrq+bo7gYkqzTsQlskWMWWQD1JcjzPq0A5yLeb9g7M1TnaDZaUNzpxvqt
lMx5LbFjojLy2gMP4WOPgH7sdbafm/BhypEsBdUaORMxV19xW48drpST3QOWbKha
ibNZ9yM35QUkbnYm5a3AYTtH7p+WhIGd5V6i3ZeeFfdotmItS8HEM1PeZB3BgvRi
+J4HhlY85Mm8DVkxoosLMOQiUEjamc7pNIWTBmJfDPRIRUM+/+o/0f+FdQGUZpG+
nToix2fB4nelPObf0LZINEjc4Hl4zLwwo1S2/epiYi+dYCqarSmC5Zt2WEcWuNKc
UpLAQzt+OsGvclFUb/lBYP/H+n0StXl6BgD8RbTqSNnx82BrO1fm4l4G9tY21k6l
Iu6LDO7+BAGD76SlHqXvo3lWs3c6V2d6QssHZgOvkhEsnThkQ+nPJ9FNZyeeOhn8
QcV1lp7MIeopJCd5aeKC9jkCZfOZqm3QLDEFbU/r52nbRmAlyYIbjy2T8MPkkpe2
SaZM8tGP9DyXcLKW/KnrCcAb5SCyP8oqe0sO1CmfOav6zRtYXbXeadOEE+0TGMy4
VnyOHLVkaE+LElocbi3PlrFq594+Z79gLQ4tnf9MuPC3Rzf+gVsTsyM2eKKHk7wI
hSeykleiHXKli8KqHVkvWAc3YOL/WScKUq/UlfbWd+8Jmqt9YyZUCMsHIsnYWAt2
oXLddIOWwOsrqscnYPk+KjH2Vriw7oiopDxokkHllpbK41j5Af52H/7hvdtjBQOh
5IS8HgxKghgA+TJNazHhERClqNlFnIcV7Ky39c32iAPQOV98MazdMRzLd0Feqh4y
MhKFoNq4nLqs5M6ZCY/8JK3jxsDbpJnQGIWvejRsFKQBgF6Kx1JPsZpWcc4wt6Vq
FuMYLtlvorONk1d5QsUMoVTTgpWoQjlltgcwZrRtgn9GT9X1P8oEIA/IEBCWtMiU
7FCwsqlop+5VIV/VjTlXNny0nsEu21fHAHW+JgdX3GPJlTdX6Ddn1VS4lgWb2ifL
dgdxHhh50wGZsgJMGEdMX6BbGBjvAlqD9/pZ9E6XpTflZECrtx0zzs6tHS5Sm4JM
bZ3YwMwKGklm3mLl2t7OQnEyh92aEYOkMx+wmlrR4B8QpeDJRd2GP11XIj7DxhON
qAWVuPOSKEuQ7cZ4krza7T8ne9H61SBuc7SA7buG/Gy15+WZ2KyLYu0NyRRtXfZd
WKtW2Sbffv3+AN/yxCF+jPeSCd6Q6qHOA+OjK2rSK7TJXmS9Z8GXTpr97DUzewy0
kEwdBWP5tc56XmVqOk5MslFy+fkMjYJ+EDmhFEdMgj1R+yMQpT/HOarFYqa423Po
VsLVEimyrJ4SRliLT4xLS9IJqxmJqgLNsexIeykl/Z9fNBVQQD1CcyhSDoAwAQWZ
CV5zu6agQyTqst0a/mdKZTAJO91otqwuMmYpMopCWR8xdAK0pFdQfrrCxjQgLTqK
L4Q2K3wmdpkheKtEDOGSVQUFtCN1lzwETV0WTh+2FlXXnApbnHVNgSqi43h9lvVa
9O/I8Oz2YxMlS58YroVFrHcOT2HFyYr/R2dOx7IYUTso83zFiP7fzaGF3cK9+qDy
ggCIVGQQE1c52Jg1vPcJpILxZndsubbEXwqL3P9rcq0PoBNw9IyxAn2zakH4x7dO
R27PKheY0+1RVoE1EXiefR61ZyGCzcTI5n49HAY1pyJAriatlUNExCJzvF9YoYdn
13TK0J+GyfmjTiXtYtUrOmHn1/n4L1BQtcvRlE18XvQEeINIIj/fNtWkFZAVK6zW
kDIZ1b4Bpgr9kcMtzjO1E6zQHN4Z8M8l063L6NZQwMMb6U2fcdWfFrvGogKV9Rp2
LDlu+q32sFKU1jM87d9CWHgqSJjiv9N2BRrkr97lIGJ66c+eu4s8BVO7l7rLpgVp
WCy5p1u9Q+GvLBe6xelKYKsL9DVusIqivMUTXm1I1eHszMtbi9lbnIbw6KeDb2Rx
oJwg8Coc4Z2Bn4SHN1QEVFQFzkrJcN9Qk+nFflHvjZWWw8IP4vkgnRhV8Bs1Z6Yi
PSL97uQum5UTyAxW27pTb+tZ/VXO6PC2RUcZKdl/vwp/qfphwsPutEnU0YlbVm/+
ickFwWs6J2cBRpXh/uYI9JbtIk2Bd13tXhyYU4RbGEtQv9GnJUfG+9lXEHx0exXa
83h6oUJLgRMYo09YGiqBp4Y87XX7RPxCOGLbHCRlDzNZcXlxpj+GktxWMNU6EZ4s
N0dH+rZ1/hn5+3jDnDGoJ/spXvmxAFEDL2YQjOQoyaeeAUHIoATk3Qb+PRntVhr3
Ip88t33cDKysNRutDo9ZfUCPhGelYF82YRxDVkNmRPs3WuuYiVfCqm1TtDvztbPf
IjhLiN9yPNvVse/YBQRmytp7vWyEudq6gCLkjEku+ljblqTzC3mSO68u0kz46oOo
rmT3uX6J6Q32qspXfD2bJU3c0qKveCPqqgzHHY5gdRn0awAOPwTuC68Bu/LzpzNi
hX5sMxympIAlbn8SDBhoiLMPC0CeBSfVl01oLy9P7RbktqrtgMUF8crIVe3J3FV8
SdWoYEBZ89AxEuv1I4JrcDQqThNd/qKvUFNkpT+PkOdHgrKnx8VMZH2Y24q3sX0o
jh3j2JKLQG05EU7uVNSd4uq3qzHojgXCIGZlwTV6xRxmSmmuA84b0ADzD1YrFth4
byGfr8lvBk+6prJzy+ACLCN2a4+04ynccfFi7pxIoSFxrXLoZCbuXmVG5yLPAYIc
N4ThYDifiWXRFofxNHO5sdRZCUNkuPWJ1Pq+DUsbTvpl83h0j1EjJ8hpzZgAjzoA
hbJewknfHlzUGADfb/ABfp57juIvBUtRqh6oMS9n4mPI0M/JeokS/XKmYCwlXc3h
VsRX+7mIyDmENgEeStvxp+xrFNbuMlMJ+5j1JCOgpGMxHwdKrGddq/4j8W+woLc/
oeEqg+H57CwZ3ENCI166ufIAPFgS7LGR7r5s94KnX7icwdkp/VVi2rEq/35Te1+o
lbPrmsNJ8zhLApHQmIr5LCh8dtoTDGcxkHzkJON15iAkCHo4fiQFzDgl7Ikve0hu
GUQGHvxkJJJzIkNhp9JsfssfSJziAVOisYlyrik/GmhrlcdlYeYvld/UEAsdQJ9L
sfnphZTGcNpZ3ieTMuChs4eP6VgKrNhS1G3WtpK/fgtkpN4tCqSqB5vnWyCL8+AS
sMIwlMjdP5y9oLXaFl3bCMBddigGWLw4YVAVf4DbuXjaSmptc1ZxOABljt2+IsSx
yFY675iFC8tvkC1YtZTZkw==
`protect END_PROTECTED
