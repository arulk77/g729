`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCQGDEzTdN3F67jgvf+aqm3EywL0qPYXx82mUTCrvMWX
huUP3bgdw8EC95uh4Xn6N2dlJiWfExh5q0zj6ZOrq45awTeR04QduSJzno21Y9kq
tmjH147zhghizaH3H7+vJc++zuzyw07qawo57g8x30mhja7aWap3AIER0ZKZusqR
6oECbyfAHsNP7+sMlVivp7PBOZn78UMwI0iS3dNjbTCwXz87L91AUrd46n99aMXo
sNcUUHg/NpdzdEcZYW+5mHAn6qRXUYxzF1fZkWqzFqTC9gC0SIGO5ITWxoXNJKjw
vWxeP1ERO3LqF3YSScAkoASIkT9ZMGq19ACDJz56suFW2jb6Q+5zonLCU6Mx3Spv
rAKnC9a1A5ZG+593LKMXW7zBjmG7UdLfzoydtGcghUlc7J8JiRucSPPoYGUoxd2M
oJs3jgNwsE+FY8DfAfUYPyeG2y7sy3fsy2SKOPRZ2s7nHvVPtiLghO1K7CIR9+bK
znKdMmiKn2RLzO0RtuXWit8WYZFiyNqgE0qLGYmLjvqrBxmtP0w9ZwhDZuQ4Olf3
`protect END_PROTECTED
