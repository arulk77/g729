`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44PR1vHCV+EYjlkGsSsMRy0+yI1UrqcfnC1dJiBiGC27
o4k+aP8klKgotP4SBJgCRPXGFJHIz+lTUIqmPSBBj9Ez1+SRQ7/9YwiWO1Y6b5Gl
G40TJhHV6zKRrL+UxvW+V+gJrtxzeTVugq9+f8p/YyA9JxH9SSs7wAvjHCDt7xpM
lsE23GIJDWVlLxieKI6QmPrJY7I0VJApW+1BueEynbE=
`protect END_PROTECTED
