`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM6Qj2+lBcZ9g+AR15G3EECIhrGb1UbGpjZGJpMQVVlR
L0yoN4sfMNwmAVVgOgqB3hLWGKuz4QvaSPQUYB8T9nQYrEkGG6UC1d+3OXxutatx
mYbl1hHDJt0utfZ+ujO/i/7MiyzaY6XrfthtZUAUAuX3JmbSZFgDm50fntK+fa5b
IjPLF7F6jJlCSKW49UmhGWCVaRa2oCxkoOh05iSuVxPmfwA7XdIp7MywmICN8jiA
bn5ivcZzdhJxwIYrmQFgS5PxdWbYVb/nnSpE39bfz2bNKpXiGXNjV1AgfSc/WIJ9
z++OGQIA6lIwwi72CNdltSF8lO5jwxs8/HvIy5qF4AxJ03STGNRZIR4Vs8ZAFINT
fW4PXoJkez39yDKF3QuHOhG91Q657jOZ+VCn0h4K3F7ieX0QlW92Hphds4U/wIl2
ggjjDOz+z0gcmSluYTXXpORIsSXuKUwztvtz/iNjaeaAI8f/fNhptsbBjqLeUo6X
`protect END_PROTECTED
