`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JyyQs+gzcqWIVwdS/x4DEVI/t+PdwxhZFLkhkYGbwzwjyEnt09IoI4ag6fC4jUEi
J7KBOr7/NmC++GGZGtcQFgJEiSdN8WVn1a4VetOlmuMyWrvkc1zaMBhV/B+FNvxb
/DSiTDCc2h5vd1G9VewV3NeSCXY5Z8IsuSbG4JC76U/B7QHDOKZb4Pfaeke6qeMc
X6n7k/eRA3lQlQrnKJvbpXaW42iK9cHWqayDSSbKFsu+BRiSImqASsbBFjpgdhHW
`protect END_PROTECTED
