`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHNr/9amVP8qxDkGM79mrVTzwm8uPVP3FoOvML5rlHRr
naW2CaGkXBW6qBjw3jVhJ0fBv6WQQXbPZogr35LV2Fsu/E+DidzrbW3Gjjc7Ijig
CuNDyZyfkabXdEB4xyClXa6ellDX4a2wHb0OuZvn9Iu20W5kbeAv8jPz3Ax05HBP
wMRTndseVivCs/N+Tusdrw==
`protect END_PROTECTED
