`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIsiLKlaX7+jP3R82mdoGS+87VF1Q5TsjOMrAAOnDj02
aRQadLbdoxdTuKdGqLQZQxmMOO209kKIqOPTmlIdcb/p6llFS2/gQif5Udk7QPsE
wUvAZrl2+dcZztvmLABsXSvo2wCqNNXG7DGhsV56lO/dFZSEcqIYKlzNKuV831dD
jmeFNBCHMulShinIIHor6w==
`protect END_PROTECTED
