`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHZ+ngkWWcN75bck7zjwVbmfG+mrdzJ61thgaRIecs7T
1bHeI5lw2s80ASe6dQ+/WbvwpyazjI6Fk+C8t4XmcDc1WwjIj2KtbrmBwT8Shg/v
vnqD+KJ7p01QlCjdJ3Rkc59oGgneuiqpAvozCEObWVQJLCkbgkZUXV3vtZNdUimQ
H2jbLAoVuhAHKVIYLM8Z0mzpToESW7qSCHTZO2PTA+q0zObBA/dBkEiAockl+fAd
tmq9av8muh/6YK+LeiQ8Ln+Lzy6xXcmVo0GVX7Gxe7GqVNAPgBF6vmC4VQ79Txve
v2iKg8JeaqrwoOaJCucWmwI2MUB/t/T5EUjKNSNIVEKO5Mgs8Akt1LWl4Qpf1gy+
ra0dSHSIHA45NpPSQmvuX8J79z0XSmOUcGzUHKePcLWVgievUA6EJ+Lxmzzk6AIC
SOt5FyIa4Di+b749fOONgjTKuiAKSKMdgNdA+kclx8HnOZpBL7LE5ZTJb3kV6LgH
qx+4P+hfWsfD0XkWdEO5Gq8yZysyRbdVP2PEKUkg4RjjtaZAT2uc+KXWWRKP/qNI
`protect END_PROTECTED
