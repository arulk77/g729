`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKpj5/UVG4LEFiP+iccyyIfrpj1ZMW6oGYsTSZ6YbdHg
zKHghcv0WZsLvm8kL/ZQiShVThOQBzd3HImXg5BOxYTEdFJr/r8ql8nL/OIB6aGc
v0ZIciKnGzV2ugccxkshaycO4H2R/Cy4ffYl5dSZA8szpatvQtRd+ew7UWhp7P6x
GZ2CcDocHF3H25Y2Ty3/+BzkVCjpF7kCWta+Yvx+YVzpc0pONjMtEU9wk7rKBc2V
ihJK/JSr47Zl3hje7stx5i501vNyzLMZFPihgfTR0+dNwVSpS6IJZknLuFTiQHTV
GJXoLYnXDnLS7t6zMULfF7d/KaecbSnzPyhOu9SAamJ3GX/8AJHSbrQyBwbwfVUU
KWkrD/SSroj5faCvVT30tXOPq4DWBSYm0A2934zVbWPB2zRyrNj9+QpTOLtXHUjb
rI7BtMRv3NLuHqdVQ9gpZUqwRKgZ6jrL5xuCyi7N6Wmuy5rQ/7KZYDlyHF6PzGqt
`protect END_PROTECTED
