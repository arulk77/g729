`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCQTSMx4P/NHjzUtHrxatErulkNln+7WqNQS6ZMltmuj
IdLkbX4Bp2htdFHbxgSwE5LoEIwi6jfG4FFMnv8UX3iD88PVjqskwfvKaDb1Hgvg
dtD151LXAf+D7UJAUcUc07swPZMOP9uBr3f3ulcF9xymTiFLElf+cpkM8O0iwWsM
gm1Mphwpbxhh4d/tCoagj0xWH/p8Ylta1lX/w7CdikmpHHFkh5en21OGcs86xi3L
a00/uBlwhuUoC4XBQzKXx6h6kxdk3i6K6Ls5SJkeQ9PMIkUkvOe5zNZYAubPhLeN
xDSOeuacrzqSk+nPhA4akYI/LGJ7PHdXE1UBG8dQXeBIjD063lQV7WaDayNzhGEI
RTrpR7IdJq47cpfSMl/Nw92o7ZxVPNdjwAfG79Z7ybLhZSioDqO2uXFX5Zun/HAm
zaGhGMp/HsMyFad7hIxq/gGY3Kv8DfpvFytD/3Fcp/ZZqE7XXsyWgBRtlymZqPPI
`protect END_PROTECTED
