`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C+81Bx3qvjd7qZVeAgWlM2ekYqCUPAdAoLSbAs9vjuze
YnnB3PSLVU3h7+Z9dDS8vFcBrK4evOv9i22SR7qjFVSFrHTbs/3eNkpImTNkOnxk
M1Orh3MpdR/pYUbcwnRxqdJv0OcjYnGmEa6a5AjGrXMG040kpyJnzhChVghrZEhd
OQt0SfNicYzVeDYppTDQ5b6Tn/usNvlL4TYNuqUR1DYMr/lHKeJKICGZ9p9+3/5F
`protect END_PROTECTED
