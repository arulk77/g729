`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG+WphTG/ZmbBjEw/7wgIJpivEOZOtoTRH2J6YsJj9wz
nrbttEcovLqD32861SnvZSWVTQ2AoSpOV1RD8HTDfQBhCKOxpVGNXK4XaIXMBjPe
CemcZtZ5dt1GTFjvi9VtFWJMxTMj346bMfLkFL4jUwZCuUYbUP9lFBBBhS6k1vFg
YJM8tyKJG3sZEUYvE2PC02UXs3aeaMhiR184A8yRKUZ/Nj0OyqjilLr+5CHlVZfR
ZOZ/wYBfqKN7GlDkP8AQCPABzSGz9rFl6TP/AR1s9OdM/HKY1fSGIhG6kyQVysUI
Xge7GJHPg2DKD51oyu7Yv8FmgHZByXZ7Vbbf4c5lCRxQEMFIuVzlF9Qzat3yTpTc
Vyim7TDaqIweuPJYMAYNyeP07CvVjtPyWohOo5pYsdLn1Z6MQXx4L9vdS1Of8xGA
+eltavDx+WvW3SZGLuu4McX8MQ1z7YDjQvX3pNpwbBjV8httX8LCKurURXxNGehC
IbU9zngtbJ9lX55PLRSeYvfZG49LFH5EOevtde+FwwtLWrpJej8G+TjNyknXwQlx
S689CpSd/ZIkyT2fbwcutbwvD/UEmOMCj72WvsAvaOHpUMyCnl1CigYu5cS1G4i7
k946ssGy+xYSc3ymErfUarKeMvb2D0r8g2KR1c48CFZTQMlK6oFmnK0afSnqCLma
5NpNBG/DFkebhiUNXayNo1xwXWenm0xENm2GyI9PRhxg/VkqrpQiEI79xmczM95v
jqQkZV/nO1Ic0BdBN9B+6tI8GRSFKyRd9WovQEElCEadCAqn6EIij/3UoZVMkp1x
5AO+nHga/ig5r81ZEeYRryYQqypIfSYVTGLtauVOux8=
`protect END_PROTECTED
