`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN/WVlovpccnmhog/xRKnRvVJY2cSnl2ZkR+z0rgtN2HC
dTuXd9kIGds4cQ03OqgzJdxwUgslHcbknmXo1OPCsrXS486WcBzIp1fvgBHEdanp
rCjwU9EwmFbleeR8+aDe1O6cQ72y8WirNCNvTqAGibc7F/Lhh+J9WfSq87wDJqOJ
xbHhA0fU8Bzk2pCpIDyqy78s1hQpIKm5C+t4jgl7f+L4NhXXGnYyg8dcl+JCPZP/
9VczJZhxaU1ByqFfEGBkY7/1cfOcPbM1TqDG/KtsIBCt3C/MALBS93bnFgXv190j
i0fHES+NzJFGGPC7I2Np61T6uCxp9zCi1eTbunew9+magxcqfkladoXRmtDhWqP4
octR7MVL2/gqhzdQ6751CZHM+gfJaHqfrRK2R4vnEkSlhPJIXVRap232908nDfRN
5CbJglIyQ6Eg2nEaAFIa4/5+4pxG3shetzOIUlJWEfxfBIb34cigi2Ye0HL5uxwm
U2CpOcX2yWlGTm4hGhmzSnK6qrVZ8C9PBo3MViSmt/Nz+g2166ygMh/114eUrkf8
ubD+Ac7zqnfPP9dqhQOyZppCh591g+uXSTkkMyaeT4sCLy0fDR3dAq2oju0fs2Ri
QslNtQrbCAhwFqqqM5WnbDgMQZ5x/L4F2AvL41H1njf/nasRuyZ73k/U5o5D/745
MJ8WN7LcNN4wlbQn0nSXn8Qn9cVwxAPRLZyfmBXF3ihV+/H1nQE7roXshBDwiyvN
x/vSIEWqkikR6IGbaDOpzeTLqg8VlmdndYXB2GX50ci8u5mx1a5Oe5/yvxBHQPys
OqnP1enw9m/tUdqkbhIccvBk36AUHyHwvJ06De2YCdV/Jo0ZlevdJlDxBtw1lOH5
J3REKE6Bejp7Td0UGP+pL3jraYcuScLmNHnWXEc0xJO+rAqWszHAaXDZs2nS/wX3
LSAVmvojH9JkOXsIBYRtYjgN6UHNlQNq8SH4j1i4xEsiKfrrsU5JimFcywiz9wWG
mH97eXiYQOK9RdbBwlnSs4sRFh++MWrEEQ2Delh3sLqNcqtZ01Q+1yCjH6k1ljxD
R62uv7+PKEtW93xILlpQm3SkLE+3iiikox06r8P9zQ/kpjbn0KWP60njbSjmLjMN
pVJ6hmg0mVtCzjP3wqo2Ihd4rSnjVkAoq5cnqZ+79nTVPsgw5i0Tz3nFBWyNaWPc
fVTaWXV8d+pqNEQNRX+Y2XOyy/Kfdy0wY5T3JCqoz1E=
`protect END_PROTECTED
