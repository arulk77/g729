`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN6RXw7dqiJPiHbe1tG+9RXPTEHvBlr1mll3zoJTSvjyT
8uKRfMNUTvO/2A+x7yEfMMPdaG6eQCcbmtCYJ1ReWavM1sQQioir6/7PhHHHgeQu
4zZzSA4LBIx66qg5aqiaAgQLEg4MGF2BJYCUPpLufjaLQ6a1wAP+c3ddlQPU1aYp
v97ZQ+BPHYHZvLdj3lDJ2pIrJNw/W8D74kNdO5E0yDN1sr6ADu4vq2nXQ9MrNljm
mVhrwnRmxr1j/WTxuQWRLjtfpgih31RndytG1hM76iYiuuuBN3dbE59xqxqI+e7p
4pCsUQS4kfon9e4yv0K4eVGvORSXUNHve7abS3doybWWdl32sjUY1SZA5b+v57gk
jr5/pVVXKSw1EdlcJZRRR+Ewf+gFUVph282xhULW62I/mj+voEa1UuRVSad6RAtE
RxfzaYHU0uorJIH3Bw8InWSc70GDPppe4Peb/b3Cx3R/BZpYGVnM59g2ZyxpvW56
Y7WPTioQn0YTnSNlcmHf3JrbLdT7vnubx7Hx2NCfegAxhYAl+1ppJrUGLHhGib6C
+k9MPXhmwvCuXiLBZZPCmmunF8A8pGZB3+0wNrJ9eFIVh9j1k/jX8XISq7QEvamI
/1Gjt/85c+MTpz/ix+L8UtbeSJV5/WQUG+9ZvrbzX+DMGaMD9RTVZEKDyLHnYAVu
LwdacuRwgja4kUgn1nffpdLn2EdhqOwcVAMKreayNSjpafN92NMnXO0cKGrPDOSF
jsmfmBaxzcVizWXkj79QnA6AqgCd3AxOt9T6tThI95rTQb4vSmtWdNslxEGmS/7v
EYWeGPThW4GT/ZxEYW9AZRBdx+8ohfnupIq9bLs/UpEqmIdggFg22A1QZkB/kcLX
Mx0oyynaQgxQs6L//Ye9EcZ4m36guUYBNainOji4nZQPoMpuq3NIDwb6T/NtCd9t
W9CFec/jhLG23jUpwqqkr7mPryHMrdpAKlm77Z8e7qW6GmiQCHy0QFf2cB80t/gy
YKXDhvRpEz6XMh+QXVEm8ca63TjhNom0gjp7jncwVCxIdlu1ps9hL5BWb7PCa+OO
ndkDCKW5UaJVXBJGbdovCdNofYzbUtTAwVqVZcXOeotTa82+obYCI8d3t11lMyBZ
Jw2dA/jQf7RMOxffMjKht5cPKwqB3Hb6vBz++sxW6s6Adb5HqltiUJMyNjP+4VNN
bFkccPJ6C28lOt/D3IPPkH52G08gNjUlpSBo+xyrg26efJfW7nihWXtJ6gSLyW2N
FXDr+BK6b92+/1qefwiBLHJWvvVk4yxlO4+6vG8ga1T6tpj7IeMqeLKBfm9dYZ5a
s57QwlH1nolHrYNykflwSe5ZEKIVlUNcakhIJ/+ZUo5JSnEJMQcYysMHF8JP5QA6
8GYfJw7H0XEDYqXkQekkOchnHyHwfkeb5AlqGTPzp03LCn05bjQaLVoru6/Ipn0q
DeA9zEUDe1hBcqUnpTgC1Jpee2wG2jTI9Aby0nNMutWxfNbPnv6Yy5FPfTjtXnov
yNCjr0aqTjhx8Z5kGDPtrgPYJm29OEECwoPfSt0j55WGR09ag4LWECaVTRSqqtKL
V6rgo945lQXOWVksa1aSUjDhfkFq/bNZR8BYNA79rucI6JVeohXPLsIcCm2XiMQ9
C9MqQpwC/zLSpzJCUU5UHk/5WLuLb2pFp0WCgU8h9XUsN/9xmzKO0x/8VqPeg+wH
9YyISaGOMK58ghHN21+ai5MVf2R06rSUL2XMu5kU+SETp16zrqV4SeRXoIftbsop
WZhq6ABtwHcM9ZH3euet9NWSz1duMZ9vaqmEYnPO2lMMka1W9oHjRkXmueZqUpJe
ANJWL+NdxcGKrs/6Svrcw4Y4gZAzS7zlaLPWxNtBJMjy5kP3m4oc99iw2i5yJRQq
DNgmh9Rt7R45HYjjF4JZ9thm48zp88M+VaeGIRFYxjoaRcCOKuhiLCRL/x/SIhMz
WRXVIN5bGdoEx/TQgQredUghPCIR+TGOckT4k1eH3VfHT4uFI06358y3Z9FY3LFk
Qe/L6WxEbdyPsg2UQ9ri8cFE6EqGTZpS7spWxKDzXSVVMuaiTOrG+v90Y6YOwCfB
D2zZySHmW72jjysLQZGqRpoqSP2G7QWK7F+UKe7YsaRvjVx++1ewTO1J/F7Bu98Y
fWWKGlQbs9CY+sQXFO2BMekfmG6CF+hXLPc4Y1AGt9tdcSUoTcIM5XqVKmf4d8Ep
+45bNqCV3+H2ELRmMOpbZWWE2Fu96LGnk6g4lEHu5dq9ETfKzsn6KlQHp7dLI2/t
EukPExNERZnUmME8xaIaRNr4ZzSmNwu6t69zOmT+bFh7geyGrjyP0G5b89lMS6/Q
dPOvfNRiNt9mH+Fw2NzFI3ouptGhjpQHmmVRfVUEDVRcRI0/oEXsGs3E6S8BCFsp
MzB6ot8r0H/xTLxJRC3mIpikt0YQ5cfF7A6xmVuNh1Lk7peuHVd2Pq0+x40q65GQ
o7J1Ra5GQcRqymPe3GVSNQT/ZsoK4FI44Rh3tWz7w6/b4+PfVRL/N37JoG96yxfl
I8eHYKxPSnFUmllLpno6eya3rJhcFAT3RqW2GyR3yKE0eocWPeBR00hjJJAT+vvv
yP3U/CWGjdhzOoZyVMLuoRTEv3/cBl7NwH4tMrZ4F3KymYRqTu7eUdqFxkVINGB+
DrckCd9DQt8sJdfD2tIhxbqYRPdfxPIbZQCJr0ujYhy0UwRMffIUB9ZPdYPKpZdo
SQz79VLRYGiq+ZbgJGTKmmWEsBwyoUDZVb1O8A3P1dSEYU8kixAstKq/U6yewbmz
XjCc9e4FF2pHsPEbcV1VUWo3z8ZE2pl/+vD8b+h//jzyvoB7B5BznUupFJclPfHx
QPydffAyW4DPT7sPCkf7vDnvdzjnGD2ReT+ybVCqPI3KE5mlRMx+T4RGYBREchR+
SlVpcAYTXdJ/2PinXk9LI7cyAiK2lDNlGmfip9/O4bKUQzkan9/MsmuBrPauWFDt
htH3FuKRrEumnopUcX1wzB9/7vNqPm6D1OFA9bcFgbDn3/a6ClIOWQbnHnxbbUiJ
GakuVcqC1hTKExN72XJDM5lO7M2Cm9AT9IB0WOJoGyAmZMporJHFwWKTDT3VchAN
76TuOVlruHrgIbDf9t+Hr9AobQBmbth+Lvi/WwYL5reulFQRrLlwqHqYd0ekNUBS
SN9Xa+eqjNJrxxgJ0rnZn3WDVWYMHJmRxijjcVfWYLqkat4hneY3FE8gOUIDiE/2
jJN3ganMXsos9M9HzQ9qKtO4sBj8SJg2R2+JLtbISEJzLWxyi8PllO+xi7q35yFO
yiDv7cqeS/p/nmqJXZbjewcZVU5FtozOwZr6myWjcu9J7rM60ajuUWPpk1hAaNlX
m4PdG0l6F+rwY12C8R/ZIc7sX4skHbi4ceSGtt94ZQT3uMTZHYuigfieG1yLUn+G
gl3KK0vsf80YbV5nO1avdar9QejnCFDO2OUhir40SlaMPfqbZbnmt/fqjryylZU3
vkFNg4R15QapWuMAQOHb+XkSpTt4tfo39uMbglUQsEuNtfZUCi/B5m+MVFGCxzmm
vlUS0cYO5pkbPkfmoZJQzz310DE4U0lcXEYzuGU/aTiM06nqfFokNapmOGph+N6D
GHb3058lCVHUMcNDyVFg1Nv9CuCuNC7PmcGi4mZCIVWzraL1Dyw/TBDOJduSZ0Fg
k9hKagPo7FL0ZUKv4y1keW7CmE80YO1S3Fo2A6XidAi2a2wpOwUxgwAD0ZrahrPb
3nffbf8UsOY5c28i99aR21rhugRN7u9ExrEkmvBXkCxN7CfIUTn30TXiJYdy0eIG
7Fk/Wu/aUYDfLP6L7Fkr9Rh+/q2SxST3N5/hLW1fuUKVMO1Yt0/QWpJHbH/mYBG1
QZekzDPsXlu82mHuSHnpYIOwm8UoNhBnMbKLTyAIuxg=
`protect END_PROTECTED
