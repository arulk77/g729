`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/72XnQn/UfH5j0HTlB3TGQM8vR6pkAWItDTbLBTpuM7
dBvO6SxyvXRUWDX5jvaqRyG0H2xkVmRhIU/f5yjBzX7saA08PjHh3fyM+gQlF23d
d7qt7ve6V2KALIqK7Y686He9ayvY4Dg+Nxvp6RDhiJN1+xet+ZJWI1hh8ma6oXNX
4KOB/IQRNQmXwNmc4tFjct2eUZzl5yjxqrmPyQzoU/LGymu8GQEalvBGDPnj9UNL
y/iEya2ID1SCerna3Ml/iIzOcvcOGROMwg4Qw796Vb49h17hK09qHg7BZwZ+VTeC
gupt4qaJbNinLPf9pM+gqbHH+F9XSyyk3fxO2IQTpd0zGichOH/KtIkT4hkI8Hn6
txuIRHxCMVvDDcFCpW1K2Q==
`protect END_PROTECTED
