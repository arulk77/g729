`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAWXpDT++ErVo8momLVFTsklaQOLaOCtUsFtMzDPIwYeD
cwE8mEoReappRQZhOVJiMmLZtJpFh7uKB57TNFRW3tH40GB10uxPzJyfreWTADQA
wWsryQPRt+kbeIDSiM/cPH3b+QJTpjQvsgcvkqWwlvWR/WtiRPNM/3rGuc9pnOwi
MAzcPdY4qkSbIPbtYZeuHMCGieNDKZG8bdE0KtHVgxj7cIBCkAXm/yZywAsXzbqe
dPXqeDbmycPYvN1WgmDPaVEa2IkcQWIdKINCXiAzgAv3TwtdwjrOTOoVKIj3DMm+
Hove/9YMQHP6Jd6zwCX1k0LRI/xHQE8ffSBaZ0aOTjJJma4wKsqdSzuJogYakBhe
OJJ2iaFuRdn9kH2Egr1sDARZLZXy9oJyFFL4ool5RJvNGjUKI34oUEf2WI6HhClV
rU6ULsETAzR1Og9i7K/Sy90tAK6T9XFDVseUwmxrJBfDgJMDiVZw9Y11RWXYuxP/
23cBC/Wa6Spl98DCWo1CbS7PXjpQZ/YuVsvYHNE5W9JoMebMcEAzHeJi9DcMDXGF
hkvkUrPYSJ3K2nAa7OEaiMTRWTG+2PUq+lPGJ22HHBVjH6+iRQYY/mAhMt17PX0J
/PZAArLaGXwzw8Miy6hnh56w5gogBZqFOjN6MEtjMbwz2vfAewwwxP3jvWEoOQBt
GBN18WyDgzb6qFWzk+GFxXlx82m8NpN8Gfm5xHMKxVGi5kuOTfA7TjJlWpXQeQ7y
yJs39tZHCPl5ZSue/jjvCt4+CMv51W2SP35XsqpRmgI2p+IkhEgRd1EGjOAxao5G
rBF2v6S/aw6bjKkdaF+80cl0kIdNZF806Ci07qTYtvp3Vy+2MpEWo7CJt89XWF8P
erBcMRpmOxHIPPLTGd5gJv5fr71fPyJIzFnifVgRQSD/wz9EKxJHJSjmsxcXA7AO
P28pnwPSqmjrdJwiFLHJ//z+2ORlhDXVWU3CXhPoVA97Z89YScmLSO4XDCa+O2wF
AtEg/vVGg4SZH4hO1zJhNkz+THjG9AFe1rIjY48oWY/ysrtPqQoqKENuHv+tlL7y
JNxS80HPFr214jXhClp53xccJv2PcsXqcVKl01HM/knTckxo7ir0a74cnuRvNZVR
rPK7VNGagWjz5+LqNAKhEhH3eNwHMLv1j3a5iHjxk2THqsQzYm2v3evGUE3/fe2V
LHVGePope5xgiOILu3EU+FStCf3GRHlIRpj2bV4eQ/KW6pVCFS221MqEuquuqnip
YZLkUIkuaE5zm1gEbCHC1bnHFZPPJiU5A3JrG9xj0j/qgbCut4LKqzbd9b/92ISe
6ViHa1VHZyq1kXhieJoa9/ENdI2lpVPNbh/CYdx/ztJ3fWdSDqHZz1+wrRlOzIvW
rygbVP8JEJo49y0lMhMzi019IyGHiBfTrX6SwCNXdWZFNxx9LDHUTpmlzT0wkiDH
+x8fO/28yU2FPZy3RwVXA+McdsfkkHz+5VgtCnsgTSILX5rwrvOdMTrpsAXN50kL
Ba+cNtJIWWGLnzPOAOcfbqlpidlm8A0JER0RnavR3qpHyUo/4issHdjOhs/0gsTI
f8oUNAwDJkAlO8VrUpycAoxd6M9LEwodSx3+/5XYn08T7mIJJaDY/87VgJ2tVb7V
r04YLCECZNcwjbViSUQGrPxjHAOYJy+XHIX9khdqPNU=
`protect END_PROTECTED
