`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDYyTdFTNc5/Mqh2bEs3GSwSMI8J935Pe3B2uf3gekY5
larg7mngaIRpzE9fK06Jq8wioXsZnyQ0dfgZlVSD3nlfS558FJTkGUEAex/K/XMv
AXj4lsiSNGLVgZcN+UmLIDvBwaOHK4Vjaq3TunhjdTod+KLCZvxOAbOpw8FLNOgd
z2I1rlhoyzXcvTy2vOYRSMxOzqeDLkc8f99Bi0AHERnor42P7fK6F+MuSr9+Kgp+
hCBEGxcn4ZP/zpESKUubXyqfMaVzE3eEk16zLuFttlMqdDEYIgUOei5ky03+ZiK2
IdLpCQLd7fQCE2+/X29Zu6iP0Taphg3OPQHnFEZx5qNaW4sT5Z7c3+RZm9MgoMM7
vQPv+uiV9RnP5z7zt9aZlh+w3vqMB76NHbQAIuDXcMF/xC8ftSwLLHfiHsYzKE8Y
`protect END_PROTECTED
