`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aRAhenyrkWhzhh0E/yuTqygi+7f+NvAx3WnyM6BZg/xN
s4XQWl6/1e+11lxs1N/jq0+AG+/N+hcpOA+xWg4HQp9+r1efPLEfh/Ce6Q76lJkq
Y2wATD9KgJcZL8aYjqTVny29RgkpBrzdaYdV0WJ9LoJzludQ/ugyAU83l0HiLv0J
s153Xoxu9I0Qk9aFDFQ+CAKvwAht4wLvLc8OPHigOT9bAuFwT3gGw4KCdKmorgAs
OtgqdMxL7neSnY0f0YVK/uzX+b1GM/ONVd+zPxtFCAEWpDuHy6dUyg0dishPUkGZ
nAP81WKn5t8Vv0p1csdVAvKGzV6BP2MI4m4dPCiM9jjww7w7k6lgw3jbyOa87p2s
qonVUpi8g0M/DVmUYXcyinWVFo74UazPANu0QgEzsUujdoH244ZS7KtRLlQYqIMp
kHIznwr1gv9buMcX9tpyB8zb+NGBPxU1tTa7ZeB9IWUD4H0j1iJW/5qhAlS2xjGQ
XKcj36Ban16a0u5D4CkD1LJoZEeFn6L2Z8n7W9NJ1Das5NqYJlJT3xxs02ixYVMJ
0SXSCROg36MXs7vCZ15C1+NbH57uDPJNZZFzTggsVCoAF6Wvd9sCjrbFS0B52SRD
Y4v53aDfR/wNEU4GlBVxNyepQCuaUaf86PKYcvJ0sMSlFFL1KgPyhLeru55bjeUF
74p6bUtqfzNt2oJ6JZxHFS2YmaK7xkQqWdidtRzsy8X39pLxWIenZU9Mnai9pMVR
TC0GPxOLSMoEM/PqeWLjJdntd2WDFl1xuGeIy5FottceEguKUtHhCVvHxOyQVd52
6INxND6V2/7sM0m58ossVwkcxJCEBmSbFq2xZQybe4CMOZDSiC9R+bW2hHnHX7wO
UgV1oTd0acPvD5uYcYr+JB8ylQr7FzerRM9Eu8yl/joHdhknlRZChSB/lzBUpGvj
WuLWqNgFzxaE11ULZIU5ZAPpl3gnGHV0T+bq0KVzs353TMpMWD2cVCPsyS0ndoTj
wq0JpXnhZdixLYvFN0Zv78ljEcZsDHnswaNvY/4AQXvwVExVEDsq5jkXxHI2J82/
z3bOjtHpduoPlVYBIc4CrdiMIo/ov+fDLeqc3IaNFVPRON4t0jnTexAA68Br/xNG
xwFxTyAM+bWC9/uj70CAFLeVUMpH0OtPIuvtKFbEgKwhDCh0+1RxuqlKx0IqR0e7
jOLHlEaS4nWBj+5YdgCp6UslW62JPkGCzSqfrmYZ4P9R1x6fadR1b8cl0EbWd3Nf
cF+++p5M/lrfy/qcKvswjCGlesCRq1Hi+G/BCE6Dm0rpWuQYW5oVv4bhz0Hfbzox
zlNBEXKsYkZzh+6Kx6KDQzZ31E37ql92FMB+FjVv9MVWfIsENPOha7ru5F1bkirW
BA0TdrQqVtQoO3O4rc9Og+RLeEAAWTVWQuP0aV0mDaRMBHzIwA0wyH36gMRsnN/Y
Ww1Q8AVIZwG8f8pbdBuHdlFIM5rhxdxcs3AQtAeBybZhZjf77a5K00FQQhM08nDu
sg+S0lg+XGIFe00Q7aDVXynZc0oxaAK3ge7vDiiwD8l3oukp1rSsnJ1+nJ9TXR7V
lCggccp1AWQPJhkVYRDLiP0hA+qyKnSwSYqzolydccbiUSpU16j3d0z+IMFzjSzZ
4N/wxO+sHWdvDf2x9OA00GsXxTAIVUijqfBhZ1UpnB9T4OE/tXVRqNKqsC4RLxzL
M7ghsMrBLmQ15D1c6XPjBy8vSjD5yPF2fsejEjY829OuenVndRk02lDu2ChbAcaN
t3pVlpUNMDD9FREkB/KVvyRlQ5z6UjKoO6mIFqqeaa7oi8TpTkrbCZRkClayPYRB
nMxYmXmU0Ve7Yd6IiaU4Cf2yupE3G9wRLyspnZImmJmIXPxUZY1f6S03zvsPTixY
g6IprDWwACasmduZoYRbkU3wWZ4qEsZFdMVVN1/99k0vq4Oai6ifSaJhX6Af70DY
BX0qZSPAj1vCzkZz0LWhdVRc9WRXJpJCcofzdRbGCuhtE1xyruIn7DAlIxSyZKAM
bnh2f+syiXqnLJ23kFZ6qoRJVQdSXlE+vlttAOxf1DA/D0+R3NwNBtIIbnw/i3Zt
vpCeKg1UbbjOqpZKiiT9kYqoWCj5cHcT3q8W1KYkzJb1n5fIDXxRdiE+Xr8ImIod
e76McvG6R56sjAd0hBrXzMDiSpZdlhrV3ua34VN3RbV60lcgMSJzvqyhW0bLz0yz
PXwbQDxkik4nxe5sLL2RfcPor1l6LVbRbLWklXbR7vCh++ZI4rQKFaqRYX7eyDE9
e6bUfkGv/maM8IYBCIEao9k+n2Hmi/ictf3xgOOlPJwu3uTVhcOxS8noo2FWvrmS
G8Ubo0fkEd8ZGBJM5Sg+8J2Rrlm800mtYnaunTXAK/ThawWaTaaGSuPLIOIEmCoU
9K3D9DYVQSgogwKdarklwKXFFsK823CUcqpfyaCTEVyk1b9qQyQO5sGCQBSSzsj3
kx0mdongj/2NTB8IeREAkIp4zfNQqTbclua88MKi7lQkR37l9SuLDY8HYby1AMn8
4g+dEw4g05LjcWWsk8RHl7QflDK4XjA4rHUYJEXk0kDGgA1dwDJtBDq8GDboFqMD
d8pJ9RjVAIrR7pxZjX+ICCajErdBuym/lGQy47cjvvRguDcwW1vYoemXwJxRAGRl
2r8qZGN/si1HabelxuPfNYCAySdXBq8jaPWXj+mt2KGQDslnH3Dbx/ebT4UEhU4a
pdrsIBcX/ip32bYchBNPWz3kH4lrMurbE++eJcAdOegCXGceTTlWq7Rx13c21AJs
6R+ZwggCbX+fV5fpTPQksVKKB5tMg9sG6NgrONfxoOtoBzfpMe53IBYicG5WSIvS
zuPgRJl76NPvS4+r2HLw0rOMALagX+jVxgGJNlxMOa2YHf3UQXqeSaz4MclhFnrR
3UhBh/Irut3ptncznFBfOUDNJKbAz2HH6hyJZ1wtLc0MZ1cXxLEDewaT7ftEMI1h
QShI/HO6POVHEUF+kgpIOKEaUk5vzjGWb6KrxkqWJZ5R5XYLl6232VyNKPs9Eh3M
bFfFjpy51Sij1CsMR0swQiI4yu/iZ5Bakj4ygRwOd6rSm+cfyYzwlCeTKpucynRx
0r4PqNEc91i7LiBSX1XSEzQ3chZPuDcgNXSsLTpAqn6TJeHcZDh8cry1bK9iNP0j
XIPhB1AEYyJnwgP/MgbrpZp/SFPCg11yxx8P8vMLQutPBt9kojFSbZXRyQVcHkh3
fxiwU3NiBe11xoJ88qJpojty7QbBXxTqFoc1TG+diGSylWQWYDggdmHVFsoYzW6d
5M0vHIvs9RHua6BlrpECC4BnuzByL+pAC8ad1BvBx8XzpQ7leHPtXGZy9VmzThVf
8PFIxMYAnwNIFZK+ESJ/iUPt7+AyU9SJUOtJ9uL9sGm1vuSRyklEt2GJlqXFERod
eNLVJj2r6pBMoSmAHVD++23GkpanEejWSN5i/+u0klWOZxL7/QXwBSrYhlX9JmH7
6WV5sbmjw/IIRJlwIfsFuEiSs3bgt+JrUHcqcjdnuJCjL0cGodRL+WAyAwU5dool
lwli+NRVntcTMDgcYDyP43+FSBW1N+LKVWz/LkcLTMtPEO4/nHT+b0KkV6N64hnh
1s+qql1bzps9WT47j3bUv1NMEXZ/pOsTh9JB6P4XSsBTciil3Q0w4QQAmhzU+6Wj
qEBKy4baQCeemtg6DYdJ8ruxAVr0wzqimcHVfpiANjXXhMj3Bd+HEl1Tpb0swRsf
J6voUA/9Z0x62zc2TV0wvTVL6S9fSZ4hPZbj+zgYLp3SVSVVyzd/a5NSqXsf4r9v
G0jlmfQge4984KxDej5S8eWWOE+UMfmogAClREBEvJ58JeHbiXNlGM2Pj1JUhTuN
XFbmzedfqd1mtcDgO8yQVb+dfspOlBmbgKXT6SOoip99zCoNGvleG5+o3RI2TKZF
8+sPVXIiK10cNbMaLUCDYiGgoGPZXBjktEE505vJrmvCw/aRdhoTIkmq9qaZpam8
i7syveQ9CwCobBfhigO9xc34Y0X4Huq7AwcZJ6vbstHt6a7WAskauCjtw3Nj6ULC
wwqNmeFgvWudlv0HCUM6/0/HtFsDdo44VtyaLRGBfHKrtwUCIxjXWdXbSWbB/+37
9OJY6Szyd0E/fc2KG3Q9L8hsaRvM7hmwkHXdRemcthKrrAOjwD5ViB9+xBsZvC3z
4eSci2A29BygGOFLPJ0M0nlBjyE8wKW5TeeiKUfvJ5mR6S2FweLbAFALTc4m0xaH
7c8m2/Ne5WM4bL9DlES4Ola8AjIkzjmSjrzmHj1REtTAY6D+srT080CWnfe6xpzP
ZXjBL8rtGJ+JbCY7XbfiAD6qN6pRBPjPi8Vq3Y/shuBvOMWSXaxp8m1uIB/WMVZ+
ENtXRfXoD8/xvJzqxXZXPObSDGUX6hpS7Li1MfUeIapiBV6t/IP/+ZLPO8Dd+EWA
hbfqVc9w/NVGxSy0zVo1+0+5U4aYK/dF195psArPBSumna99qvV/KQatHKvF0pdg
59Pgo5FslGj4UVs78nhvwCSsfES9ndOECOOA+75eRemvCt+p4V5MLjJcO3AxUsjD
OcfAt3iDebIytnhhcQ8l8RP73nndUyKYVJdkLSa5W15t7+1a0FbLdud+iH107HZS
bT8ZWddKX2OXaCxdfXF9JIbFv+LgIexKSuc5k246RQM=
`protect END_PROTECTED
