`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
0f8NG+qbbZ9fOvrgKO3o3kKOIKQU93mMujS/RnDFxPgSdZdzrSWOZ29HFslK29eY
agpPLFmgRch4/TxOwJMBFh2cukhsXbvimPSyKh04TzfctdjjJZWxpEh7xQkLEYN6
lPkHyTBOD0f0I2yge83Y0Fc2F/ZsbweLHYB4kR/Tiih0SsPzrvt+ABPhfHHYGnEb
oUBdNMbQhyt75DOyZGL7zLRhE83zzA8vFqYNIShhuto=
`protect END_PROTECTED
