`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41f086Rl7ygDd9t/lCRD8bwDQAHr8tmEfYiHLov9/jWp
iPCO3eyAQPFPGzW02Ad1nW1auoojbgRFNcaY+JpOcYmaAgmITI3LITqrs8z4UggC
8+IBBJNWbaN0jfvyhRbiu/lOqTYCN7FM8ZDCG1ODrHygO7fQGNrbpki2wTSznMSd
QpMfahynjux0jayJjy/KI5ZDlflzuwWYfcg2N3MuNAwKZWOv0gOGVah4yR63Oy52
GsWgHn4CHW70VRBSZs0l5FuwW8bLoWhDQ15qQuNNH9G8RKsfSLCWyNBDHn6O8NFX
3Pr1FF85wpydq9JZZLyTidAr3yoMwB2bmcxOhrEj/k9yjAbC5Zwg3uOQAOcyZpvK
pFse0ka2Oxn3bEHZI1HR9w==
`protect END_PROTECTED
