`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Un4uxtKjE7EF7MO41dBSSTgDIOUntsGFcdqdDjWnK67b7b2AtTv5pXFHR6rXTZHy
ywY3gtX9GmAVMSUBBNKFAYeBlewsuMHj6ixROdQFCIBnFBtY1QyCxU96PJx148zn
0uRZbRO2DjZgrEka4ME8JsESOK1Lz8L85348B06CKGjv5+JtrLvo0YMi9i3GD2F2
b12DFWQkNO1LsGqk+Fec1BHuqrDdisK68tBGfwDnjCiSlQiuvvGWxLShULZAfis9
EHD2kqyzZ4Jbb39WNX+cDE6q9qpuPjgNLPuhsPOEu0SMBEaE7IQYsbk01Pa7VCxL
`protect END_PROTECTED
