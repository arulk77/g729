`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
gyxnv60CHScPz5rXyLyjcWhE3bpkzQfMzh1it6H+wJgzTa+IhaZlBx6hV7u/jfCp
/hY/E+ZE3VameKPsXUDCKiDlOJKrgzQ24H18AMEO2eEvpFBft54gQuBk6H0N5QAO
b13c+g5LJH1ao1qy+BMiHC/RcZXDc20F57NNvMVQ6XsAiBIEiCssMMps+FqWa1vs
ty7nDmVd/OAznkBHHq9rggf+oQXKpkcgSht8QxPfaf6cQ91HtIziOYHiBcN9kWHw
Hbjc2Vt5nbE0cibBNFf2droeX+M/oGmlgAa9dOHJPBa0w702pVX/mz0OnRKHsNZl
`protect END_PROTECTED
