`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2EBoZu9tBf8wFLCnm6xiMw8wvY5tMo0WwXJyofbBnt/d0DcH5aMaqtbrIKdefEQG
pcLSs7m2qie9ivaz0iqL7cD3ysunru+sJFicgC+lLwymQSThOgYWGaFDufj9XqZE
EQh0u8lYnFGps6Bu0XcWbJUXnkImOSkqQKvMoVq9NDTKSxnHmow7hqSC9LVZxuAQ
/ebfKz7MVMxvs1GLa61pXWhaCWjzfPVb3jofmJkkM7OhRHTvgmth4UZiHxPs2vx9
`protect END_PROTECTED
