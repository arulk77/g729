`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGi+yGfRrZD429un6mH1si09FLCkH2Hvoi6EYAvXu42X
uETgckYgceVCXS1KRceXMLQ2+QYCNiWSeZCn9jpcbmAVy7906EZoQqDrnOyGgl+6
NTzsK9GhIE5jCBpYwnLQcSRoKYfCdNE8abC5roH3X7J6aGDNyeHXo52HUgqkfDDr
cgmc5LZdriJBu51gxPPbpuKMKzIwPKionMrjXBSOdk1sQ4o04go+DGRg3d8iqVyM
Q3AIKW/0xAA8ytTCmlNXirbJBJOjxMObwex8wNb2rZLbYIRzgSMbMPfxbvNu377q
M+/okZOgFRZJQnNF5HBEkpuOT8hO7QAkEJLmJyMCxHpyWcSU2S7TZ0ehPVhMUq5I
onM7diENqeb8d7+if8y2H8fI4Q+FHfAmnJ2pwADQ29b9FwuaYt0ndw8NtO4HafMS
`protect END_PROTECTED
