`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
MU3QOAjQ2nMc7SY41Uay1Gi3XXtVrVDEKLRmQi8y3PGJfPF5iJfZRO5Z54zyDAT6
YH/IqVs/iyiFytkMTnh1ePIsGCyRYK4WX3GyTJrLD7pS3Heq7X8UkZyakTn+04TO
aCzkzQRAFEwTDa9YIrOSWiRPnm35xNeI/NJhb4mLWfiejqD4/sa+wmleM//S6Nxe
9OO/NYm2EXYYm7ljmxqIPXUmzPbETf2CD3QsYWQCzpp6cfCAomVIP4yLbleTKi7t
CVfl8hqyM+eO/4LxqkG894deX8iKgIXd5sDn3cw0FsPvmfqyerR6hV7s42SIbxiJ
BRBISuV1WDEzNtm5nfTEMWJj0BTi4DWeXoz/wsogKNLYsO2lSuQJfUbgFEetkAQ+
Pk+HMvjj9JzN4fUYOTWGaZG4mo+v1WgCunCooRcjxqmxo6OPsWtXuzv5mBcY8jNL
qKwfes6Y4b5cb02mzdriI+DzWED9RSPSQFglIiT4p9aBS1UN5z5pA9V1a9BGuc2s
HZHBtyPY/KAeiao1bZKlWOX4lYWjue2qqKtzCjo+Tq+ifDoU5agbxE4atKymL58u
Gll5TUcxY7mVGcBE6aPVZJvN6lNNx/5QSlLcePqVQ74VF8sGsaY1WaxWCIXVeAA2
N9+PmagAeOEKlmt66MfPvS+4GV+oZ9GVCXAa1S+5tprnlFlIUgQnXWFONqKCLsOq
UKR2qraPvttoxJy6SO534HvTEik3DPC/4fZn3Ra1bkhDFVpnlJuYRr66pe6YFL+A
KAab9PvPv1oD0xUuGlF/kCtew522QyCoeGojdtaqA1Mu6LD8hXVJDIWjQ2VZA97n
m0T2Pl/44KUp9Ad51+EqHf7qRgNBFW6tqNLj/2Kz2KKcl4KMEMvWU8k5qp2O+O80
G5JOtghCFxru9nE71aqptQ51sqSGmc0PjNaVnJJDB/gBG8SbS/82tvdXTsQlzxKT
2xQHShctZaO19agXdlTmC4LXA/Su22hTi3EVTH+gTw2dCdBvb3eM333+8Bw8uez0
jOrcPwI7HPOAfu/mPv1b1mhGXS05zzDw4vC76lLdCUBn/fBlMHhmR9o14dpsHXXj
O+T7GMzpgTUejYSOhW92b+ojgA4eHMpOed2etLvtEF3BVKia9NfooRbXDgPTPPFV
ankDShV4J6U/yt/j+QuHbdU9+5eXcJV7aPn4yi3lSQ0714X97nfm0fCDiHMnjZCn
QQaUyqW6hOUqIxrW9D9EK9WdoERjej6FD36ndrDlZtzCuowDA6715uyvVmAR3f5S
tMcLCqsf/CHo8rRfktXeMwvRr0gsqQ01OD57CHpFG2INu0oFOi9kISmgxmWv6OCE
qeU2I9MADw2ib9R18/qvoiRNzfS/MDzUV7GzWZ3aTGHlq70KyN8KYqAAybZuuRGZ
IISmr3hp3dUCW66d22KVF3CirnRfiwJEYUCm19FYd0t2M7DoCoYbfy0jqmDPPQm4
0rA5CIOkdDxcJZPC7Zz0jeTRPe1+mIaRwBHiAZVVw4nU+ZKDO+DRBSmAJ4oKGKgI
GAvkzDmq8BWSnitjtSJnO9uumcAdZdXaib2r6H6AXUI2Qii3dl8D9naRa1Mz8Rtu
8kxWYK3N7bX9DitsCXq+goyNgxmLsS9YQ43utuGe4JeYCa1FIOazN3VkaAadjHuS
4r2jhkVi2dXlmTO11f0igILA9eyJkaETB4tfR8oB7ZB+mhK4GXCzFTZ484d5ND9H
SPlzZu6HM3aA0MLgR7JPaZjRjbCyBCFnIf+bTB5Sg7+SgN2gUUnCOr80kfvlAtJ2
`protect END_PROTECTED
