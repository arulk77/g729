`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
D1kOeE60VfEqlhnGtvzMsZTg//68HxQESJ1+uFRcDD3e6SUHadcTTOe+cQZkwLDj
5Qr4q1WoshkJ+aE2UYdmIABEObevNB0JU2Tm1mjZXNR0Z1ULG6Cr1NDO/vqs8Yjj
j06F469Z4A6sZqx7zjwkrwViJgi7m3oFGGvTxkkHBopg2pXqcn4q+g8gKDlvCalm
iEUeFekTar71EH1jIDrRpbq6Wq9mtSc6aTXVFqP8NjmXw8P+IQcdusiEr3z6ox9Y
6mG+ARR4Ochgyi47weZakYC79nGRt8lgAAZ1TgwPI4M+YVHfIlY+8Ue2HNAnHRX3
QV0L/LlPKQn3Ugrd/nsXoCsOB2mXpaUQ9Wxtz03hIB4=
`protect END_PROTECTED
