`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu474W/z8A9NkeSULCTT2AoLhLP1rQXmeLAxD3ssWDpbCP
Nj+iSGCoLnAILlvXGi7WISat+pdw/pKpt/mr2W+rAaOhNJ5S2l85DHTJDLWv91y0
Uoby5V30MsVDw967bFe018x6j6VKIq8a6ZNYKIOFENXL/vPCsB9dXwOI8oVJIt9N
2bv2v8wzCbnYaPIjgbCdxCTPO1fjni4KFn7RD2asG7fCbGXL8Xx+L8FBuqYkUAG4
zLm79FZ9XXZGguuI1Ag2gr+Cx46yGNMCCf1F5tNDKfo=
`protect END_PROTECTED
