`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveO0Cxn+2Qp57QrEsUp39XxdCV6x0yXkcrkZWlJzn5B4a
fRcUu6CLuS/gV9aD+L/ZEsRKKfmUAyKvzxXgb+P0X3Tag/Q1xSGzf8RmP6QTZCPo
9chbz4iVfVVNECNVelIygiUUxAFrYF8JN9QooSFRmXtQ9nDcP9OACt/DxIY8SDKo
eP1gAuZSKyxEGyk9hy1R4gj24zPfZ+ErZiusvcBukIVjsky7t9z9xuMV7pVic7X1
Bv4Rg1mt82X17XEEtnVoAw==
`protect END_PROTECTED
