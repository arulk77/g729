`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/M39cq88rk3ckPqO06cNpU+1gfy0tG1QAlnu7slTY35
KnqDLpwIffjY/xc8VFdutD2xQbJ+EycvExMSoePcLrWroluVKkdU34aEummmY1GI
AkmRyBHO03cymGxk45CZFWGfPZV+DYW7XmPDfkUQeFtrvxn3mLAi6d7Eceq/Iav5
IoWXdugLjZLqwYJuMewp3Xu0TRZjTXI5o9+N0UpW1zaF/UBz5Bj5/SvEOKjXRB1s
nfk3PMeNOybX2/S87ec1fLLEZEvOg9Nn7PUURTrMUtfUiazZrzAkX8meJY+w72Qz
jC/SkO0F40imnbR9US/kHQ==
`protect END_PROTECTED
