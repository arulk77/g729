`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJfAqNC+XfSuhjabbf4bGFH8OhuUI6nerIbQqPfuLaJi
uNxz4JNUpy5eOey3yWfMWQNzmjaTSTZV4uJuDWXbkmTmFflMLd3DR19F3U5O+jJx
AzFr+00ALKR4voNkS0wQv1ursWDPtD1yqbmy7npLz1lz9kiZlB3sYAP2yA3kgWSz
j1d3EVM2vXWvB8P1koFJgBFkSuNeq0680D+erBbe3/mKfAoO7zTcqGVtjF4Pb8Ar
oV/0IEuhgSRpKIdwDUuuOdzjF+SB58xHAP2Iot6dbf6jgYp1l6Db7uU+ZaiL74c6
+OsAdQ2+LNalLftYjobaNO7pEICYm9x2ycUwzShbNKM+2+FPpWt01xv0YdPmL4oo
slP8VkKBLYg1Bw5O0HqRrLfmkhIuzZtIjYPhcs+IN4fLnfcLXf1f4x7Zpnj9T9de
BIPQ/6dFOXUePNMKc1v5jbpUPok7/WgeGSdvIrxldBJ1GWRRkiEz1LwSIGkZOYl5
JnMeZJqoMk1Lgncy8momIzW6wdJ8QMc0mSAI7yKN2A5QhIsu2mTWIGsfP12i8wmF
`protect END_PROTECTED
