`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDdDSmBhXcE/U8KHLX7v2ks1jPLKeou70UTyD22znGpj
FdHr1Jin2v0K1D40NpWGQnOdhYAGz4IA4FXccrXJASglLNA9PLR6Ffk4UjG/ZPyY
tsro8j862dDcnHK1xhj/O8QVg/j4QG1v7Yc8nktBhJjcTsOIOirQsMNwkNfLRu8I
l3XVJBNGtHWBc3UtpXD2i/ero/7zq+nF2nuy88k+DPILQ4sHxbM06J7r/sEA1ayN
2OFg+0dAU1dOcDTJ81DqhgjEPMaL1Eckm7VQrk2QpTI09F4zCQqdQ2G/GBJrzYV6
2i/MEeATgJfL/ArkbSw6B7QdtVHF3Fl4c/7zltMYcsujpgSa6YSDdsnihk5S/SjK
SkPlqqRa0/MCUm7QSR/nXE0wwBBn07SsvtVChFNxttoqj+fHHjSR1WfJ1nmnjFCg
`protect END_PROTECTED
