`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
NclMgSwWfn7kpVSHeTvjMCLs/qPndJXJ6YwW8K/l6SuCMD8Du4R7suOyK7lSO1Bq
SroH30381EusjhOwhYlvwjl3r4a2f7odF+DeKh5lZtVt5RaaJBKyipPUG2wUnRHd
w+5xuFpxRcSlg0eNl4zeWQzdglKRBE6BqUMC9H3XoEHXE5BHlR4v3AamE9UDUOyE
Sdorn6QgZPTdCYUJD0d6vMlrcW9okH+H6VRC9jGCwJAyTPDfuM/NDPPsSCdc2tgj
`protect END_PROTECTED
