`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI09t5NLy8aN+4/pPjieEVDfd5T6qY3gNbt0Txk5c/pR
5MMyXCSewsDTHKwmMVt54xV+Kc2QqeqnmlxsWLkEAqYDN7s6AmOc9Bro5OLIxj8e
sIurP3g9kWbfebjsTacEhj/upCRSwzN0CglrOSNa5cH+7ET+446iQiVoieM0M8De
tMHSuF95a1CXvNDm63segEskJ/TcJUaxfwr6xZd/GJPRl7a6YM/IRn7CiC8+4bfD
Z6RjJ1TUQakcjjplEsK2P69CVMT+JvLxL54HZFChTq7Ou7UkNXB3sVTNXrVy/IBg
zS2igCh+TOmH6HjJyHPGVvOqcuGv7tv15S+BiyX5hdcmNt5EsTl+JUYJA6UWpUQt
IKiGp8eX4ZC4eDGlwLyZNgBL/ZZTcXuoJE4tn0+KGshrcRYR5mJdzVIuucdJ8ebt
sCq5ZmcDc8CCdpDYFHPlEnWifYONxiwwXlZnI8TBs9nwlfpqTkLCFtamHNwXpXPA
EJnSLBRyrIu1+SCR6s97qBaW6iduqybI1bCzOTr0eUIXxXBmQ1PNWu4mmdoS6JIt
LHFR8A7cFJH4kTjvZHn+FGHPOi37o6mVj7d9WlU8ftaxQKpCZYxUfUcaaZfWPRxh
wuS6H9gBtmknb3xQ1rlFsKpnhQbm535DB8QTsum1OJ6lRouPc3YIl/b4Yg8HDDG3
wDneyv1Os4SNzt0Bn0bnaUEwyf6a3J72ap5OzZG4OmAc1oKbgP5B9UkbHBwbyGhE
TKfGdoLarUjElEHLdIj4ZEjrA0hxIzH0iKjVJXR/daIj5zcBwrviQh/5HNS4hqq0
7YUr1jBVanHllhnSHtgeNirSphBfEzCwExm7JOI8oqo=
`protect END_PROTECTED
