`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
tw/z8E57Y+/Wcs+YJw9SVp4Ic+/SaX6IAsa4UMVMXbtqa8iwvwZxY3kzYiY1fPhu
HIcJrEdevxnPWAP4OJS3Ctks/raiseJGXecfA95GUr02L0Q8WYOABZoMwZIZzLZC
3ZMjGMkD3FTOAeaiIaC8vGl+rUhhjARFh2L3j1M8FdSJnK0697IjmKtuFoS0gpT4
dA5mGYPfnGCFyJe80TG7qL6RZlqC2IlWmTGljBGe4r2Mb1cV0fNrYak3yp5tWI9q
fPxAplI3yHGZ5UKCZ/FHt/oADzXulr7pFfBSQZLTHm96aG9EX3eELBMl3l5iR30J
7BgjYX8uJuf2jt5CdzGSCGL93Q9oYO4BxtIHBsBLsbcfdmNPcyfYYhRMs2Zf3liS
6TPLdC0lJgzSF7m364bI1Co31/8qRQcwyiEpR9v21lQ=
`protect END_PROTECTED
