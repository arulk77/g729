`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+xXve8mWBFEmvt3T9uIv8XBzfRfmki6KNKZxugldJzh
lPCRgEh7fnT7l1ehXV5tsV7RYZOR3UvAQaIKkeCJO1dcG9cEDDRUid43kzPhT1Vh
X5Uj1OgxaIPOWLs1XGfUZYCDMjAVEMFM3dhm5YCsHQWDQQoWgQngjYdKzOIatell
kRO3MYQTdX8GbTKlSo6dXxb+bZt5SqqAaVlFSYe5g2Khj8zQDKWMm4b8oElYGKQl
nKxGG9pjYn/wp3Vo9NaTtCxxFBXoF2K7FBze5PAB99uQTpRiW9KiE5O8HpxUihc7
CYWWsOllitZGSaUw1B76kg==
`protect END_PROTECTED
