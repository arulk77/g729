`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
5MVd/WsTnrAVmwHuNI0chk7FNhXaKL4OX4zI0HwaNbXa5ddavUgmtljdMmxMDTns
NpcJq/4FOl7eGLfLsmpJ5zJyr8rav2qaaFGCgjRFjTyjzVN1Syf2G+juBgUoVa1b
Y9C0oiywbHmdtdpYA/gIv2jyfSvOz06BVOsBpKU38Yqmcyw8eGgg15XX6GnhmyGX
0vpsiWQHIaERM5xJVJbWP/QhuoDI4DXOFStBX/j4AiO30NI1hZeJt+L6N+heCE36
xMmd4A1FzorzW+g+54sqBp8ropU/Ra20939ELRt65gRDZQf47Yg7XhwKvLNv52hy
w+/vmJ1/q1uGQuATNM0nL+CCE1LZacEZI3g7fF8AM9qz9tAFt3lv6PfdHT0APdRr
uE9+UzfNGdz+Vy2tc2EUW4EuE9bPojd1tkfuO8Zvx5Nt6OQ2pLDwSnp5G1xakMYA
MGMrtpGscpZsw32OISAd5s+WzCMdmAdcgksRhZ8HURPK6Qgi6Xnk4XnQ2C9hj6GU
NkwNrH6cCbPnefQQpuwDu/J3Ti5nKAgPJdf1iARYJIO6q7a3wF8VqkC5ttHn2eNT
w+i2169ZYU9OsLqEkY2OYmUjzAhZ7F3dnbg8IzS85XZzpDRfteLbKJ1ERKG05RwF
loazimRo72wI81psstodQ5gtlDfP1gweZkYc3sc7DXVwMzH7qwCnG7FoG0fngvS8
RMJbYsO99hLj4/kONBgnxO9+67IzCMCjUPc096ZWmLDuoE/nE3EO1YFBvrbRJ5yA
TzPGo75Y0UkB0jV1a2LLoM4LVOZdL8ymgsBphJEeZv3Kpw9He/zD4vj/FP8gCiEg
9wfRVquNGJpEp8MghGlN7zTzcJbkqsiVYsJgraxtA1OeXsX3BHOf0R+zIfnnCovw
ozZyu5jsHwI9YlD1H6or6MVYeaMqLwKV5xZyblkqkYGFRnrGLOZRnGXP0xlFvqaa
PA81p53KJO0KPolU6jxk4LTys5Qdk8/r8ilxYYwqvLEe9wXC1m32PI71cImHcUbe
1JBcRxK8QVcLgrKdcj/r1juo00wvFjyezogiTORSJdI=
`protect END_PROTECTED
