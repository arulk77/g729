`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveO7JAumzQDQIOGCM7Z7DYzGu/Q4LcW0zaqOzjghtLJFj
Oi/F91OkXaI29TD0lFMSGHA2rZTzTDTKw44xGNyr25xua0y1Zsg+gnNiIx2sAcHk
b4lZ3jChn4DinKNtkT92EISVdn2fagqLuN/aDclJ/8GcO7OBZf+EpMfyimxNjE/z
uBYIBdTvmqYhSNaWL3Y9KQ==
`protect END_PROTECTED
