`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIqBK7hMqJove+aCBCL+fDfiF16cla+sPp5fqHeUf3ca
CqWwGt7LZvZH+FYQuOjtgLRBzlJGvTr4deGMTgWomBxcJ5hjbRX55xq85UrbIm0v
+yQV2qBdUtehQJm09R1oX43baAD+X/fM1WNv9jAsDGXa9XC6nsHm+UigAKp8OUfU
SAB2GK3B+NyAg6NYzaxQezdUazEzwWbSIuZXEnwrk3b9se3i/FwwSPTxA9XxUQIS
JIXlSFopKhlJ8sVwjZYBY8ztx0zFtatM2J5LMoftWEZJBe6P1fVILa/aY3QYlW1w
mIF2euL0dmWeODxMXCFKrZMeBJOyGAvA8roPV6Yzl7WmgatelG1vdg+32ctaoQ/H
`protect END_PROTECTED
