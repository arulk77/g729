`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zel+JbMVGf/fDkxntyv1PDPbTcC9tvovGUkliE8as70
cZKDY90TA0g1/7f/AwsSpg5qJeqviVXPijbdzhxHUxWQDFYa/ryqZdktOM/0Cxbp
v9gLGJ9bFlzIhewTc9o/XRTJtOMM9OZWauRUT1wJG6+tiWvUoyFq3UK02+4+zJMS
AZqdPKUiDOFy4m8SKAmTksagqsOziEVXjVuM8sls8qV/mSoELyZsu7Od0UsCqnD8
DRS7UgjA/etcuPJY3xwcIFlSBY4jPoulIg6/n39pCh/B1ux8gdn7EoqtmPuu4N0j
KKza2J3wZMziP9zzz/yXySWPNiHYfLQJL4zaw28OrV+gxQzFyLIFVO7LA2GU2Ljr
fl+Wk/EEUIJiFFl5ny82Jg==
`protect END_PROTECTED
