`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMcALYQu85+5CADmlrLKmzAdCKA9QY0YkvIlHrx35ane
DBrISKTocksAhA0Pw6TkANm5pzI5WeJzeNUNLu1LdyuNGsSNODTe0klJA7ourJ4p
8DUiTkSGc3TD49eOyXZZc8RK2+VEBOlDIfhLe6Tbd7W1v517bNJTptot5GrENs82
Jr6S4i5ggYgUDOvWuS5TjA==
`protect END_PROTECTED
