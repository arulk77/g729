`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMxyz0vL0gcdSz4YRS0qmvuNeBDG75LMmh28mFro03x7
FCBq3i1ZuCoFCLQxj1xvYLij/5Eh9b+WuzfdD4zCfb3v747pY5JPwgnijYIOhqg7
vMHOmnTThjo/kw8OmJvUPQJCi50GO50TgeA+pMJqUbcpUO+tyhDsRpwEtl+torJZ
rUE+LeFuB+XU1JTJIdW1b4Rb3thvQRT2WtKSe+OV38WCj4Ohos877VpiOloWDVOy
BpU2nj/ooWTxT+KjR8qRKuL9IykFGIc7N0IFdANcAWqiCpll6LLJpZQUMbCOE0ZA
GMcG+ncIVoDXl8m1AWDWc90xJFEcJL62qVWhxb1I7yNrh462HayGiug3y1hhYzf2
Pab4LN9WQrK6bhWXlV6WqugssFNdaQDSjmUFIohYWDk8lQ693JZonlKi7Gg6MCzE
vghO1gMQyX6SFqJ0kJj3dxznGRM/mOJcjpvXfuNeuCr1Yy0QeKC096Oih5cEsbcE
7SCvyGSjTMIve2fC0uOLinCmAD+uoyY2iBRA8tmZRRD/EXmCQXThZoTE9YxcaSqz
`protect END_PROTECTED
