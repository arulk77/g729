`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFaTEo54G9cFB8na4TQtdZn81veStPyXKcbWYx4ZbKt6
ApihmhzJim2ocGzzxrgxob5fynRdBj0wzkz8vEUcMdmmdTOwD+fR7BzBlg5lpvXY
Pj4rCBgIsq51sn7iL8pPlJXynHo4/rBelNkBltj+7NWuUVE6Fc0jUzF/y8xofVtY
hqCX0rU5a9vaeTOt8FTbiMGXQMeDL7elW5YfwQeVG9oaCopKxkFlvirxTCLgle6J
9qzzuSepaXI1O4lVvHOqfNc5j61kMa7227G0pDlBPFqsKoW7S8guvXFwaz4Vyt7I
QLuuBNJ5z/RCzEQE2rk1hyiFkULA3ULGTrWhW8h6D3x36aAC+UIihvORPIzlFpAN
/Z5FF3T40SA5s2chjgiLssls24gjRj2GpRMFJ9EIAK7Qj6L4fbC3ahwWDgLHbn1Y
4BpkbBdzgu06jB063ZJcARZI/M8w15an1mxm4dOaPTa59hMpFqWW/UrnE8x+TcS7
XKyPhz/hePWXJ19zhEH4Qp+5VRjxP9DMEEygE8Z7WvedHqKTU+LZDoAQos/eSYzE
`protect END_PROTECTED
