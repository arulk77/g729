`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFkmkmgw/EuxssTZ5H5keGY+2nTyYJYESJoP5Yi7ptNv
mFp0Hx1W/bSDMr/orsgqEeEqqpDC/szTj9pgEc3KX1qv7DKuZUdw/gZP5BJNHT5O
6ncUoBWOlwCbnoS9cNlrqzQx+a0f1bYvn8j7grQRtiR5JfhpOTJlg9QUeQB4NeyT
KRfrnwuUQaZtabICzujelpvHwoCFDYYtUVbe6xMdZUVzGC0ksIs0K7x6LGniW4bk
fZ86be0qbXpSkqaqR0W3ASjUraag3pGxAXsseDeQSDzQUUX6BCtbjZQMBdPjAuP4
FLZ1pfhraiKDSRLosG09L7L551C7CprAhy37bB37HvvcCwlOMbH/eAMApv6VtjgF
n+z+KXwLe1F9Z4J/9RZ/Bw==
`protect END_PROTECTED
