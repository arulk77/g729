`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49eN0w6M37Gj+/wphbdQi0APAz4uvsGwyKu4UeXh1PAJ
Iokl1J1kWOaqetjztRaFvM6rcp9VCsC7Eh23njOLhdYtehzdGnluoLCaLaS8l7Es
O9tmpJ03ayIbFKtbEB2z1MvDNUHDqAifBeLTYvmEUYQei3KZI3UlD0PVIWRzzm+T
Y764+xbdxgJaahhj5+DukelKF2gFo1+FGW5/b3aZA1UzCR7rQTQlC2B8PTDFAecp
Mc+KXFfOBgwXAUnGxnuy7zJXPWhVsrXpuypePAEZiBz1KeuyiDY9GT6xUNwC1chs
JnRDKqWl2gEN+RVzHBHn+KE8/hzJ0r8rkSctgvHTuOWsn/HvAYJXxzjBKfTLoP+C
T2p02L6t1zNjKnXTbVskcw==
`protect END_PROTECTED
