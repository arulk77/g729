`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aWU7Cpk9wcGUySMst+w4toqNmruEK0qOt/OzAcks0x3a
cJBwTs9nIfXcL2brxIGMHU6QuF7/8+uMRnRtrQve58TgLykzZuqd7HTqu7cTLoOw
uCkx4UWsck0f28WICPLF2V3j3w1hChgkETPTpEPJH7yUo+t55q4aQh4DBLKjMtX2
osPYyBagfmJRi48750T5WyZjh1G3G/7etWxhSW/wszd4BKFkqOVbObvTqoqE29NL
1sHcPe+xDCeP/56MqK0fWUvLDwJCYBtp7/fYKlxiTT+O9kls1rVN1of+3Xq2w1od
eDRaSA0EEvTINQKikK5lSfo3ohzoNOpf1kwtVLWk0wQDEVxNNZmGCXYis402cxIS
FRDIqQ696kEVfXADYH7kvA850U5awXA8dj95dlTfHTGN5VFYS0q2ZtGSF98UFe8G
aTMoVDIGFCOReR7DOsKNn2EPTxqglnfclAIW7UuIURR0T7jY9DDfwTLdc+H3DHm9
Efr4nB+H7TDrWZO0gicTsUxCMtlVFXmtXJyUkoMeWM5h2sFeC7RdEBeTXFm64C9y
h1HdD1L70g6HBAE58j4xwoZus5IHfWLR3GR2OxwdeOggdPQZcLOn8b63un+tV+Vq
iUE1N86+ZqeGDJXRZ3MCivLhYxju2porwAoKIp86WqopMAhuuDcwkFh4BQHarrkH
zF4JGTc41Opy4Vt3tk2k6UAPhj5dL+yYH6UksaF+RwK5rwb7M2V0ubie2VzsNp3I
/6PZ3IXkaa6CtS4UG3XewVfuyQhOg0+PPT8yur3it6uoKfTV/qibAcsQchV6p9kh
aRKdHoA0wniW5PvYf9SVT9OHFIEF14lWHhKaan3/gDIyZeTKWn9M3W0LNPdie6im
X58mwT2kgxkP8llaw/+x4JsXvJs+4nMlA2T+BwM+kzfENl925ys35Tx7OHWpfYQo
EvQouADrQL1nWEajV/6+FEG0N8Vkq6lcq7Pu/FYAJ38ra8W97H93ArxD94t4EsHl
x12BJ9nAct+5lEAo5m8JFCADGDj4T3unzX9LF/777j031QjF1Dj5v4UWDum01uX1
FcASAHhlLmUfrrAHSmEjmMivcMzSdCHDFqZP3SPmqrel6QowSOt0giy/6udnApTu
M6FtMq8c24N5vtoSp47EZUMVfPd35WADDa1FWPSpbhPqWx75xDMSYdIdTSARiPy2
XSwRGz20xMv1FradjcW7Jt5bqEtbo22Vm6mvQoXGs3eO0rXEurxm2dZfuFcyWKue
TWyDbh1LF8S99gZkU8cRhZa4PdZA0nijDeEm5e9SUzA+mh46Ha5G5Ck9zV7/3HIw
XOLAlUa3jvUO2EBFnAtuYVSS9XSyzk1vOd8mEyHdfliiuxrJIOa0h2ckCu/OjVwK
nC71ALP4eqblxJxGC+iZxpBBUwCJm8KhIvTeJXzk/9nnW0ar7H3S8tVx+7UFm7fi
mwJydqQla70A5FyY8LhkF8JGr36kOb3fYrzCmYfB8jsPnk/rwtLEA1HrRfiRFXPh
2CBbgunR0uVolyH4jwAPSkvIvyMYhdqfmoVYKveNKRbq17OVCGST5T1WZ/OBYkIq
+22jfLrWzMMckkG+TLr3s92IljCiPjGTdqpIFPQa+dZYkaR4/Uef/qBJPzO5+8hS
NCv5Bnyi8ELTE4bryvICplYYyzOu+BKnwTvpRBzDQuY6DTtAr0RkfvkbkP2jpqnq
DAFBibf0xPBJ7peL+pvl7aua+eiqUsKXE7jdq0GtAd/hJrCikT5miW1imrvtax8v
x30oRRZrQtzl3KqwFD5LUHNfIMekAnKdDx9BSuvoaGtp3K6LgBBhLmbPmaIHxSrx
Sq2J/hSr9Z1XmfpJQdX+7d2iFd9lg6dEpxURt3xnG+aLnyaeKsFGo9PBcEZUJba9
2m+PfwoaSJ3PlvRTBt7Y2UofIZwVnqiuQ4Z4unj2/r4/2hKkuwykJF3TEoMTx6CX
yXg83Ypy5RiLa9vGCh9HWggMGvyPXEXH8Yjpk4gHmkRED1slQWx72CWaD9DqpmRt
m2ET2osOR4x8JX71J2QqbrPoub3OmiemWp6Dwm92hERw0SkBH+CBNZc0HE4YqdjG
TLvfjHoZYg0wLmCST9Lomwp3aY23W4EqALYqJfEHnwklqcDorOFsfq7GpDoa+9li
clUV4ei8gnke8PP8tPgtX05Q7o/0KJJZPK+R5jekhgtrLxTYgSmExp6CfhN2MltG
7aHVOKVV9klZ8dUgKmCkcqMIzJknY9NC8KtHblERQ4n1RbDQKL2EF7rIv2HEQ6IP
uKO+XMGGk3sB2/I4nCjLb+W1b8NGDlfu8cBUfQgxC3BgKyTAVkMxAbK3U2HsY5qo
ZZPALa81ffgQDtFNzr+Dr0fLMR5XyolNSyb87YmCaPhe4Esj5lVRWbc7EZu+a1HJ
4JI5RnEMQgZdqmRKGQo7PUpoIh0OsA7FGrngdyQMdiXLqTbB3+c8t1lfSFq/DHhI
QRSQjZuXSb6GkBaNsJL8sJKvablCjhklMdIJgYPeVuncewQ3YCIfbRfQ6gTo14+K
gIRP0IRaX1gr1OzEEfkM/Bj6Xj0jCOt7+9ok28I0YBQmBCboO+RkwWDT1FFwZJ2P
Q5d0mnEtrtz2jbxkS34xtW3DRDbElisgGQialmaorxpOHvR15w8ebdPBCMGjllLn
WO2kWJi6Urvh/jRRp9dgaH9H2vT2IuAuICroWfTVXXURuxtR14JgIa/XfEFutOgl
xQiFuaNqEowCX/GRpKmQ+QSmXuR5pAJAZxeV1fLCoOWyJFoTDNfBz1v1ylG4kO7A
`protect END_PROTECTED
