`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBSDeyLCT7904j0WmaMo/Sgpr9oCjAG9VQb04MhUlZTB
TgpbcN09dNcQmp2U62puWHxm/Wx8uwU+5bS64IpCeE2saYxHVMoDuPPdkpNtEQyA
GNtD9uYKixwxDOex36rjNABDuNkM63jflSonMe1X8rE5UlV303VlyvM4COJq4D2k
ltRXDAVnJOAjIyLmhL5nRkackUr7XWwxQYhCTM7UwJNcc44yxBNYpWUThv70k3mM
7khcruSSpjUdZ/yYlLZUwBS5uQtXigxG18uEgpQYqtIq1tZBkSSHq5c0gWQW1k7h
vodSXhCF61Tt3NyI60oLYp5qMUjWdc8ni7m6/6rw4vpJHG08Vz29fizgp4BYMdPJ
beSCsNmZIEMjqgUDPFYYKw==
`protect END_PROTECTED
