`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLPznfX+0TL71e0rJjFg9dG2q5ZqwVVrAvZQdzSLq4sr
D9iaW2X4VfQMtlLMWJmY7id1VYY/YYAIg6+fjeFs9mowZgBa+1hRJbD9fcPKbWYV
Yc/OAO8Ns5ysQS7sPxWHd9++KLQqCpp7IdrN7OFfsGhyxtq73oC7jmKRbMI9Ndkn
YtbM571s+Z+fCumr12lIYpvPHLAtxbtwld3jCyJ1puM+TLvxskXzDTCmgCN234vE
jMo0kC3rJsJe0PwhPzAfgRlJ9opNzyUtbZ1suV3/HS69qElmHscbADvHqqJKgsZo
3lEeGVuYCVGzJ+UqFUcFNzMpsgvArXw4Vk9iXFXeIcRIf2QQu0vX8rKTc7YFCHGp
gPeUofE0x/Dzt31eJNzmcY7mFXYBs3ABNuxA5U9xfXiuUkRS+nwCtZvZP2Fh6Qoo
E/uXJYbB630f7AIHo4ergzhkLXOZf2DMsj0krAPuRvqElxO7ju+FJlVz1bVzLZYm
7/lcvc4TkytS4iHDcvXUtIKicL0doCmmlcCZogQkSJIvwdKGsuei8LzP4/LyNYu2
k2Js8v9HEjLdn5SjtSBEhrjctWZD0t7qfzVBd040XgV+BFzOTDTYNo1MrgyZNRFW
HQouzV5lOWL8CeHWvsjOrx5PHP9rR/7MRV350MaZ7mE+Bekusm3yAgxMFph+VSaB
`protect END_PROTECTED
