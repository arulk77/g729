`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOSOVyFqC279fB5m7UhHRBJT8ORceawQeQufkTcYMFN7
JONTB/tu2ECFJqijBHHMABWYKDZiF+2OC+GU6jLyxKG0dDW8jHBzltNJR0JLeHp2
Asmu+mvvU24VXjFQBVYe20Csbxszvkgv5WCP9v9tjSKkTBl9Eig8ZCfSphzDQGNO
7q5mShUv0J6jPsrQtwEnhlud8W1Ed/Ism/2UGZJTE4YpEYqXUpyYTeQT/p9CiDf9
z83jLaHAgM1utf6psWFWbqaO8yRm1H/rFzLcCCqiNRnrN/+zdrtziilTU/bLKlJg
f1VXq2hrSD/ykwY27H6200K38EP4rHxnJ/LO/rbmymUhqyugqzXQ/ey7UGxDoUt5
Usuaoz38JTkeNezcbJxmDyKsRtWEPc3J8sHA1ZQNEgH+A0RRzBux3Mwjok9OKeD/
Lvd//mrW8VnplFr9O3F/lTOwFMonS2StsrrtfmhuKx4ddVgKP32wQSqJvcRmG5pW
JDL0PzVP9qT9cprj0V/vfxmrFOqd5CDKe/BSbklIup9E1XL6V1quspyzsNzP1lJW
`protect END_PROTECTED
