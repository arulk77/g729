`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNTY0LDJW6/tqN2/bjaxZlTuzUgKZ2fdjCyDSKgabtRY
Jq1XNH3SNFtOEZj80GkbCs1v/dL9h/9E5v0f53axv5G2X8tTNWzKqcv7DilesyO7
avtvLKFT4+x3Q6UG3eCK82JmwqN94hErIi/AjfZrPdKr38NNoVl8DmnDufzdakYJ
diXu6aOTevZIQWzSYv6HL0IRonuDXlLcw2iqLVAeMLVwuht7kItEzXvAQamXyBIS
JyQWdeqXPYBSd/chRV168Pgd1LJ4BMb+VpTnlvCxskcfkuVZ5Pb0AunW6N0BkMPH
kpG3Gj7nyCOyPBhVp9e6f8kyJD8gDB4DDXP2GsEic1BL5iU8lweZ5cyRE8IfGD5R
8J4ywgpT5sr+nyAn00m3wmHWrPUZt6Mf/SCFvh1gLbuxl6jRdA0wFcZf6Aeghh9R
dMT14DCWi8YWwMsGcZn8ThR5HGwWmtJ2BDEFwTmjjFYfTJ5oavQmE28fab0Jtp3W
s+sVAIDldugZ1YA8z1MN+wxvLaFYlTcvt3glbUMthfdP3IJquiYUYgg0kb4VTwn0
4DhK8Opu9px0AkjMpkkmgw==
`protect END_PROTECTED
