`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73CwrSbt+ApzAfGmcN3XpjsPPVYIl4IQRbK7TY35fg0UdU
cWk4dUQ9saQWi80JTY1eXFnf9UX1UmJhGLIVTHSS/AdDzx7oUhq4V3fEK1NP2ZXI
amikLJhY1/JxhbrqrdzKnUZThkH6vwRNVTCXNJpNxwazhhoKZ9fqA9FlweelZd2G
V/n23bbMRegiRLgjpl2LBHn/2kPNgBPXPdcKRfCia+9pDk9nEAYWMF+wn5nEm76Y
rI0ozXtT2iitdfdHB7MIkUnOWXDucTs7mzYx5YxlJ8KXOCJnyTYErwidtsHEdqGl
gcbIzGQ/YmX4rjGJhkuCOlK8Q+dNugc1WFOIfAVhQ2W7Bc3xxliM/5EdjgjGi/ko
wkNWfO7q8eSW+oynHZ2Y9AgDDddHGcFL8EKTeyi7eZ8xhTGl+dqSB4fnCRcZPj96
hpSBW1AP0o6bP3ml9dE+0ynsxB5Mwlj9Qe0mPZOWTM8cEdjtSNIKW5CuwxZ+fJ4/
CHZUul2pRKxPeDHT1BXjlgfNfp/pP4eHttyBI15r6mL6cEKwIhB8DbxmNTfpCWsS
ujlgG3tD4o1kUFU5qzkHhqwPumol8Y6YJfK1if2Z/IUpdiVLLKQOkiwx/hoarigL
FLzLjKxpEWF2LnleYhMirGFpLcyuIFqpfj6822G/aGBrnd266m/mSjOXd1x9DRDQ
0NJD3gldyuay0IWCooZZM27aQkk340shslOuEgrZUEnQQ9OpMeORj9hfAeFntYK/
+oz7Bydk2pitYyoOX0Ap2Ii8POKHREnqVImfLlKz9BPBs+t3+7bSKJ8p7pKiZ6V6
WOWsYHUbtN36PsR4Mh7tukGUmNFHj894ePXUKOl9hISbeU8z7xpu5iwy23obtg1n
j6DViy6A4/lLuq5yg4A38rFmWB59XyAKw0Y+IHtak7oLl5TgEBDfRSAUk9e2wHPy
IKlD72TIsY0pPlEwGASqMwfC+qvWF9E1UwNBjzth40nmnOo1RLRzgDUVF4m/AjXP
E01FnrCvsmlWVrXI2E7QQSU/g4WeIaq0eD78RCovsoqlaFwkQxtN51hO3IImkomJ
U23v7mpRtZW6U0Sto6RhHKY/j9RfQ4SowXKPL0zCXXDBJK7T/0qlQxsH6aSPB3vR
vCRIiAUpbcZlVJ0mcE4/BWa2wFzNrqqYl8THO6ifr0WciKx6sIRKm3Joq4BOBrXs
acpo6B93BEfrUp0HUh5kY5502DC2RwEHOprkK4MiImj/QFX9n826TPE4o1Ky6p3T
6hG+nxA3xd4HoIp9U12qzWpNHpN+lOD+BekOyk4Fli0RHMTDILdAwMHa64s/V1gM
+EtcntzTssbVozEZh0Bq75J+5ou7FkbuWQ7rNZjdjGxURyShdG4xn6qKRe8Hr8PF
EyeoSBS8xK3iZC78zzVLQ05XMOgst/Vt/k/UsPoFqce3X7g3JTjAaj71ZfrrLjZ9
JZhnKi9++6m6SpKH/uAutRLhHtlQ/jrcbbmCo8OQGgRO2RvgP7+YQKpQe8+zJ6k/
x5MKYUonJih1Ri2lQP3vccLuep1yPQ5RoWvxrZEYxR5UYNGuCp5a9m+stSacfEKV
l/2jAElQZZAmAJSgUv41BPhtC+lodI04HWYG+7DMm+/FbcgGdJjGLc8+V2hy7Toj
ELkTKluZJzW/kdc6rUh5ZHWadN5I8uImUF1X2bzr0/urC/cS+uc0xzulyZLB94r6
S3cqX/unvjDzwUHwlQt+WQTpgt8pXoLkBtuMWv4ZcDD6qu+WEKosPx/Qu3x7Y0un
BrIWQb18P62xMJSrAOm8FiB6MBx+y/PlahM3sV1e3/4wxQvbeoJJRPCq4gC3E/bl
Zvf16u2j8SWdgkddVhc4WBg3yNcXN1TYy0J1rEjcOxyBEqIGyddLLevFYQMT7SSl
jPB3nLWrVtDpiZC/p7I4S9skMmA0SNNNgafEnvWhV/kHx3GOPxGje+l8YjRwrAtn
5luihoKLuyRjsAmPkkXRSenCzMb9kZOEvEL0ilRbSGktX4cXN9lvms1fCjv+Akjx
rRZ+EbQHvnH7sU9eDECWjC/WSQBDwaIDaCw0x7hl+oaym2pPCEAI27n75EM5KCvq
S24peCUaE4i5GN/IXbm64+LGynzp0LbmyfcsCH+1BA3FDhhdjmLXio2PZ2YGMi/M
X3bjB0hsnuWnwRY7u50/RRy9RW5NWCAYp/TTAkR2fhDfIJHTpX0b6DM3vGthKEQH
4NuJD8D0ZLP+UBdjwosmHk3inYYIx7ZE6vug9LdI5qMij+IWBuR7PBh9IBBZs2y/
HEupPwvqJEUx6bPs/xGbYRNkJ1TLbHMXTG1pTbDLHvyPnzUyTZ3wmuRCVpClpGtl
wB5g95EgPvhACLiQkGaggyBAI66hZopMi78RMwDejhvo8hpVFjg+ESygJcA56vzk
tVFKoa1LZrGJuufrjQVUEXgzQ+E0CtYWphCYQiXlb+aYmhaWlP3+MipS5QXJ2ao+
uApcrhOaUJeoqWcLQMs3AN+nhgJIIhZwZ0wCMvlTn1KuKTjBP6QI0qOwyI1Fai3l
J5L1qmdBVTYH7F+KMW5v6VSEdWqziuqxbbXge5u/rAkesq7uL5TIVYxGxc3KNegL
VlXg3q1jVe66FAPcfORRLhWA749AF34zBN/A5nYPufp14jcAc9KXlMrP4U0z+8Cr
McWJvnsUeQgTncZjS2bzd3GzF+zKeIuWsIRn+V+yAnchQrOGiW+XIKZCiYAx7vBx
GzozY7lL6W4mtRYIhqetC7vDs2y7U2GsF/wLi2shBSAVaeb/Jt/wwsIHkET2i8YF
tUNlMaF4DBsiNU85RarEs6gnVI5uA+eT0OqJrfSRvSjd1sHVktE//CcgMpXSfDUU
DLZgIAYTceYu3cJxTe0NjVEC2kV6rJ5e5R5hm0hKGLCIKWtyeBZiRxChpqEBdRgx
mizqyekAOeGYOPWk7yXOlvbefxN498EEIye5U7bk23GeXNCY3UFDDhE0nyHG2Cdj
CErGUNjpxl9YYzh8Hgs2rQDAtpNAXx6pwG8cg4sIIIec8iWfHmSMSY56Spg20muS
Mp05WRf7z5bhRxOWM9/dQ/x7whdI1T85YGeQDUPOpyW7DgHu1/ZAaEMw1dwiabte
neTg8JIYGKppgTiMSt0+bJcjRz15VxFube2QyMJLaz6lJt3PWSsrC3za+606bTuj
WwQUCuSX9XF0wWZD5QztbsuTtL+wqpkhy95v4I4OaLsY9JbaGS6R8eyltt1q2nu/
g30ljQ8CfaK5CTR6u48vvWafGxCmr12yku1RzOO+io8dN3ZMDRegdnrGNX7Xi0uX
uFJAfzFo6+Q2LLKJnQ0sUZgMMhH/KwDGxdamrGVnnBI8HNjR9fpZGNf7yqLBsgI6
/DeMTb685x7UmYvCNLAestHYgOf8lMcwC4hKDcZSpwMG/AX7jzKKQfZDBqWFux+/
BoQBZjmtEZ3KdtoCYEUSYMyyIh0TnBGsOb57LzcsOjQJwHgy82UDhAx6pcy7a4ZR
wDl5PzeG5yrz4wYNlH0FtUhdMjH4cXUSTuwdtACAl25elSMVH7FpTyDCOCYunzTs
TvdeKjJe4aDgeCnoAsEGIIQ3/yANfFJ197BZDhJTxz9FsyBns5tlvlqtOTXocNZm
7mmhbZ4dnBLNd/qf4x1cAc5MrCPySQbd2bdMoXyclbMElX3XxAN+xygyUG7Ogwrx
pozlOnLVciaaC6Vjc3+S2krJ1FhXH3n/H+O9ha+1XuKRAZjFDGhEbyfjTc/poer1
DPuOwA2h8GEhXe6GOPtBfofjQkjAgoNiXTWGzkOvjvo3UNK7n9rjTvUekENO/HwA
QG9IvBfAZycMwX6+kshrSRH+BjyG3Fikcjr1KITCoMWSwUdVoTuUIHNJwJf/ARYm
c76Tda/Pufrggq9Dn6hEBElbSvUstdSR1S0jV2O0bNvdlhAc8+1WI1ZM3JB1tJrQ
14oJ0lMk5D/55smafIajMoTbVDKKkKSOqOS+vwG8CtfMgrVeGHWozuIKkFUjVP1A
+ZN1kyB1yx6B9UIqpvOeEA9Y5Sd6DuAPTwRaBnMb8X5j0ck/fLCQnGwIMW6udnIS
mLEBL4X6U4HEBISZc6yn3JOA7H5y1WTx6GepFk3uEd43s1xNG2lSYHjvUK7Fvedu
eFQAbChuUOdrqBQBNcz0MIbenY+B4RsZ7W+7wefMKrJPlG57tVuOec10U1z72sX5
Cn9Lt97spi0hRFBo0K2LeejUb7p4RpAQ+BauWa5/IYUubwfI+aZlgZiE4JhBlBVk
noXS6t02oi05zY86IWMAUIWkx940B8HZWmOi7QoELOBEltEE5e2N+ywoAyzCOOAE
nG+0ZG8uihYJKrAACEXLY810CRT7jLtL0Qvq1+Um70LMk1ShJRLm9esAhg2g3UJX
hvxomDqOZ1SX2QyyWpLa+Gu8BGxZIX+PLv4j7RQoErw79ombOJbbY7TPE9yY+mUj
FkzeXA8lYoZXAAQiX3Q29CGaxYrVBEu+99Xlp+KIJzxghepe1Ok4GADQAPtorkkn
nhPrtQ5rk1Ubw11etYaNC7M2ji+bFBiIv2p78Bq77C4UI846KtsDXGdLyOCxmXYh
r5GWjzmnNZ7X6MOXGPDmOB4i9D/TcRWq6G3QK8QHYNsETo7BWSjI8VamZbIbReTZ
Gcdl+C47yaAwjnV0Chkh5IYdI9Z1guzLEC1+11z75cmas1pbGv1g5yAE/6k+Tsbg
KkTkUp5iD6M2AtJSEOqq+AoLzMq1SjLcPg02G2Fd4zsn1SwlTz+6UQH0Hx1SoKdV
c5nFBsU5nxyFJrxx7yBI96PzEZn6TSZo+zPneJFcCoicdrAYh3pt9GZt7pSaE0DY
bmLOdoyxyT85xKiJ3ruhAQEs42LEpwyU2bGlb+dOqdrf+MV8+zxKxArvuysgA4Sj
sJDCMCkKXo95mavsFAji8pgdck/vD0kK4JaP6cEahW7UKGIIBh80JS3hELCcGPoa
nQV4hpK16cvCIZ0Vh8uqDqCXBQDqAomISp9xw+IkkGFgYulHHMR9PfEQoCQBcw4l
zFfN40MnpYUwFn5RAh/Qjfcv3FzDnyxAl5ac9SxvD/ltAYAkN8+/dJpYVR8OL6a/
BP0MbxxDkDojAHp6D3jzzfhBItS8dl+I8/6KBSW96wjHw2HkZYEbF8T5bPM69wBf
N/j2wUb5PL+CH16Iy7WAwYZyQYVWVd1+1dlHrlFe4OBXr8sTqpDYeD9NPxFBcL61
3QhhYuYKYEbvQxVMqbkam7vqPZ6EsNTSTriUO7RPF9RfMAk7vjNO+ad5vN1p5OBr
M+vfKNY4VgLPsRcihq7eQKZHybuo6irxVvunl+rmma/UmoX23NNwpBsI8tVy+PUJ
CM8/gSTKswqgF0Qyw2BkNtfX0xGG2tIKC5xDrxEmdkOJHH/1/USk5t5a3NRGZdRb
TQHTXAHLNOw72StS7dNZJpaBI8jpvQh23OwAEvHU2YbmEClToZJ7T3rhpTBz+LfX
eARJg4sCx5kDA6aPKAe2iqObAOREzlt2CDtNr6DP9abo6hgOt8hMJYBhMP6UNFXS
4lsZU2Z+5UH81ov5uO++sTF4OCmmp4IGw0pMkPhXgQbiMPJxoYxt9sSHqg81YIxy
VbIJu0WQcEscGTgdU8c3C7FwlrL32O8C9Qxq2WslVe4pf18MxFDEbNBiuLIoRitu
3hoT13Q1TpRqd71YviEQ0JKaKACbM1XciRakth7OQSHTE2wMPg/UIR+Aa93w94K4
2zzcKN9fzTh/b1Hohx5KPL640qh8cnvIdN1EqgnKjh7uXbdlvYfBY0SiaM4tylzE
Po2rk+vXhMZy6iEzscvzfsUSEdikOwNATiWreemzO7Iaa48wC+Do7jRiZvAEfqV4
e6fqxV7gvco/78nD8AD9WnUBYdecd2kJlRuJKWEIh5N9wXSCaUPeLasGhL/+66Qq
n6+oML4CSGCvmH14RqvskG5gqd72dvHI1x9nMBYieHppO7v65cuNG4fAWjX4PsuR
7mbL2nAvyTewyO4vM7B8eK2QThOq1sB6fM2KvHqZ1wgd7WxKJa98gMcuEdJtq8eP
ysc/vWUvtJRxdJ75HSKKXg1kvVdSuYe+48q0xVKsVEMw0H2UZWQ/Lq4ZxjPKlVRJ
oVwRcAgRrP5REsMoOUAuDngtwBDHHsPvEm0vdsfG4lVpLB/3LkrCwbF2IFTomeNA
1VSrLDG1VFO/Zra8wNotGXLwRU9xfcPn0gFqKb369bQdpyAdm/AFTsMv3hwQrjOr
E2m3DhhlY8YgfSzs1U4LPos9cwplXsq2pMa1xmmtwkmmkixkwwYmILIUaTowxBQZ
cUF3ek26vDPXsZkmQ0xkfaqteSa/oX0qUfV+8mqBABNeo2r3LintZFNv9SfEnEP/
dv77v+SkX0vmFKXgb9FVHv3PMNDnnLyc7lhNtg4PCQ6dGXEO91Z3R8QeauJQRIZn
DKx62QiY2mDH4VMr0341dkzdpbgAlrUi7LVGlEC9rfsj7ccYrdMiOIEcggX72BSj
6+6i/3Q5ZRG9TQzmriaisyGomxqlcqsDEtgBCx3CPW+nw7YR5ihdZDIvSnX2jy2F
owDPFcrlZPcs7UiYxXLKHXy3Vfq5+g21vUYAI5xgMaxOS9x4sFyUGZSMo8eT15ay
sjCpXvvUZAkhKrZA1BgaCQYn5kb7+a1FH7AuiMTDHKgsnZOEBA5yCjoFo4xZYgSJ
jQgtohxCcMWOxQ1XTRi9+uZwMOK0tyKdMYLTMBnKbxB3gyRi8t8TKXZDMf4isGT6
CntaEKKlSW9ugNlC5xu/HgIy2Mw3FU8l5jXeKxeMpUqY5vDBL5PhvZU3sgGzHuws
Hngm8cUBtGVzVzmQzOsGUWzbRTbsIYzFZ0WjRtIp5WS59eJN7JbLtBHKexLwhfNO
cZ5z6RWrrSmX329umjhw/QRHNxH1wcLGOFWElgEtoUQ2ohNWlZVSUOgaB8gIIiVs
pvF/Ck8KUB/MVqbFz18RPLTJP/WnMKqekl9EkiQGNzcYPEuY4QFR/MGNbUJrmaeJ
h0u87yYv/19rucNNyLv4g5yTlSHHAINXIeurotOHHL/i9SWljHZJoRI1KBsPdC3j
DtJpeWNjQKEBXHGUHCLmLG3VsyVXyzKdOOnHkb8zjJmi5gXudUwSOXnKVy3aLZRY
OXAhyaDliJUzcWkAUUFF79hWUeBgW9qrrOYo1AW3nuI5V3BX6Td/T2BuQKoVWeyc
S1kMgo9tEvU1mR6yrdwnP0v4Sr7l4aliwxp6HAv5mkfaCaYJojQQEMtwsfOaLzEm
2p431HktKzGYc8SKNWZlV/xXfMe+GpTikIx1TUG4PFBM+To2KIzUeXDYVcV/61dm
Whiz1HeoqKoGEo5ndsSpD4HQVrOdk2G0Y6K3mYt2xg7eiHRhcKrWpTRmI9arPMio
u56372o8kREzqL6zg2W6iq3eJEur4ZhVKU2Fle631xG1j7uerTbYGd8G8HMKltUo
ULYEf5WxKEQ/UYE+nnzEqQTrtZSKBmuCPjGxe7lyaeCoPL4fzQqThx90VTNbK21t
uzaELThb4n1ol7CsyCFLs4Je9LihDCpuT5j7TSWgooYLzuFdvB20mcCAiplHGNHG
oJ1kfONPjTMpM3c2gKobRkLJ5aGOnKj4JjkQPR1NzEq3fy9Z+7uilYOlCwV51nWx
XyxRTwreLNnWqvHg3yS0Wmq+2nCKdLEj9PdhUJ8dyZzfaSjExLIJKSL3+EUvdSuU
udlelUxIGSxsNtX2d240xI2Q2ctCeemF9d6FEm8xvv9AbOETo9+XrBqyEPPhblSw
FgvL25VJTWWZLTSepTzr8UdPcgaVGhmtrbGBdGt3yDuk9VVaBpDlU2kIARjxXwsp
sXcxfpeIRYGRzSdaiIOeZ9JkfEm1T3iwQpnkpFKruurNivVu4rNcyyootg6InvO0
ONmZz4PXrDb3vLhJpQOvyMVvSWet+o/RRetHI7TMCT+/v4A9DtC3a+ZX0uX22T4t
mvQX7jFeUgnj/aFNbGp2/9wzgF4edpB1s+oJAJDSkrWVG/eBLRdlkskUs009449m
VAF0LZWR343F/7GWxx05TnTZXNve0SdW+2Y5zF71SMFvmGUVad01TWecGb4tH5Ne
JCi6HN9Yzd5/QpU/XyTZCAssOPbGF/mk72qv/7I7Pzs/mPAHgXTJdzDQuVnc6zS1
WcrnDkPqyTLvdUwijV8lwIdlaveiY+knf9YPPBKnCwro3PaUPaEs2RXBjNhsCpFu
8eMd8OXA0kIbq43tI5r9ISKsAwoGa48rinq/J4+JqRW0qfq2dmgoLT/pfBG0eGaf
59ipU89LhkH0v8bH27kDxCv2p3lRI46aC64LY/TAILwEwVxVNSdATOIqQdAm7Nhl
7IML8veToa4qtzUdN2MGWvUuS7qUWUfXKWs1+EiaM2ltKy12u9hyO6q+4fJsylfh
yNIyHt9VKXkaRbQ2XsQcmFLhDNHvYByx3mNb+ySorYoAcbGMILyiJcYdGPB+aIWs
NYLjVk+438soISJuH8Fcsl619g30YuWOIZv3Sp/dU3XztNYl5dcG4ez8GKbgUrdV
m1qzNbWbOvCC0d68lwHApuG9aw34zW/MetHjr/h4mvPCfrHrfe45PXTjE+jJnTk1
4+iojh6HiapbZVqVQR3NLIe7RnQ65BiCCR8N52xgdScj9UoGUbU03TAe/WSRuhTs
qlUz3UgvIJfm1bRjjAKwSf7ajv3IKLEUeWRW7wkqNqkOhBjPV9GUvhJcsoQL2aLj
GdnQaow/ZuShut+3212v4cJRlv6coujoaFCz7ChcZ4osfevxBaEx89G0pHqO3qMZ
FwTskjDy7nDe77nIN+CuNLOlXbAWx5jrEBaCOeCu9QnpswfAUFhE6hVfq57eQbyC
lbAjGn40+X5VZJsq8akDgSEdlbvVtFNqSEWJz+jgQLRSU7rTlsP/mnUlT/qdDKmA
xHGBoWiuKvGSFNpGYOivFuSXjUD2zF727lm7UbTT1BK5f3n8ue0QGL4s1Kmge46e
eOCAWOw1vMoJf0bPnEQQimDjonZsbWBaFtAKpg6uuWfzdOalRX//z/4ShjPBfcmq
htLf861C524hwF2zl3iNLexcAjYtc9/+bl19d7dqP09TWBHLUj3fOvTOok+pH458
cLyodElAMAW7zJ/SG8Or7T2Dptb6bM2V0heBHxSERkkXwKPwqrTO1wxaYKO4uiic
R7e2sLnF7Ix6zlrAdfumNr4n50M4qDFnrUGhvJqdmuTII3z44yqsWED55vt6JDsI
N0ccKjWmXPXInphdHYKgDxwaPvMlY7QhF/O9ec9QkhUy9e+IxNtezdGy+4BHr9kt
2kEn0BX57w/3u4lxWZ0hC0BEO+eCDA0+ymHNcPqUkfmjgjeDtM4lEUqLJvllzeWM
n7zSMbDgCvhCM2xtJe5FLrK4Id+d57ny5xKIViFDOYiCBq/GlsG+ettgGcwjt8Bg
MazZ1b0P6uOPydtir8W06h6hhSu9ifZuGytRA1P3nR7iEgsr+5xOlLD5I5UOz9jy
rKeHgQHKSHOHdvUMAQax1UJuMT7QVIIVNrOnD3LFyaEr9M7h3a+LC73ENLOIsy7S
W+4UxTQt2kyppDhivNA+XIgTrdQz2zyCQ0ZAO/vwS65L9hlENrS3zdlpQ/SuU1qO
EjGrRMwiPxQUndv50DdDd8htpelZqgQhkzn+uGQkR5lgiBIh95IGF1btkFzFNZrp
/UukuCVhdJOlZbCaIeou4Hk+bR6vQRDqx326ebsXuLfJZ652YFh2FIlnopPFJkf4
71aUyA8JDI1d/P+1Lvx/qDUI7F1ItIm5h0y/fFkvG0zwW/ZgMLQB9/ku3eolHJRI
sojyAWoQA1MubC49V+p3zVaVyLo2hRaLE7iCQ4dGA5BRfyeyytwLXXNnQGp6/m0z
K8iNjtbVPkB8LyAHRL0lVcqdi/6g9ApgxvZjqh6Mb+k3FGD56PcFuhla1iziN5PN
QTZt91QGETDC2peVoDKysBrz+hCxuVuDLOc5+NtwNPpNx1ksdlu+RJVqmxkXR4e3
LQbWW++0cC+zoymsrNMThVxa+l1hiscCyU5E97TWPgi55+TTDKpX0xtZAw2+a6jd
WtbAxnNgLju5s3Cd6diVfNgq49jH0hpP1ytJoRjSj0e5moppm9qcy1K8cp7MtpaX
vExJry3xQE13tZOT+tNzSdH5jdjEaTIiFZ3cikkYeE3hxyzsGYlQmqKcvtsBOPMA
jjSQsfN401GCN17cGCenQhYR+x9rlEVUd6jZsu3NTvyZLryB2rXKpKZOa6lnqu+7
I/vUwmVedM1z8N4u0ChVBvQ8P3caapZrl1Lkky6+2yCVYLMwXhXdAmhYsROgtVJ7
RogfVf7lUmnHMFw0n9is6MnzoOKdsLUXLPZD0ZROd8Ac4pDcWZO+AYmG5jskB4c6
9b61EWMR/BtIe6s4jh4A+6rfTIDQW+DXzHCvRQez1BfWsR47mkECDF/J5NICdjyO
WKEHD6mR3KxgrWBKiuClPGaxmyLYgEJi1XC/3vWh3CFQ2bbdADnQh01EM2vK0aVs
PVUs6FDw895Q3rSy0oaLdM0QyTLEvqMU3KkSeJPuI73/O+Ze2uq6cyZ/bSZaNOkE
i/jyfUUBAvKr0piVFvRx5f8oJLNMiro5HRy5BnzQVcvY7+/4OnLHwIuNUp4yfO7l
yknOlRHL77zwVtLaYCCYh6iVipKQK/EqVm3fhAgzVt82BDDQpd4rlHyAiSW/wBny
fmnxYZVAWJbS7wQO9pQR51rNREi9hm+mWEal23UgoKjIk87JT1nahHQN9WLbWYse
Emk9JgRPuuWTERLtDSZ37r6/dlWi0buVXVo1SL0fIblyNfF5BuQ2IAzIx4JedChN
gSS4+c+BcXusQxmsV8aehdSgquX7H7g7Zz9CE6PnhvkimYOnlONfVYzBqdlL3h7F
Op+XcoKflICNmxOtVKhRVP7LWJiK8ik/MF9jYbo4ivF6ZnsVpkIlPPK0B8fDkO8Q
jIr0ANG3Rh4BX4xROz9zOf+DUPygXluCydNB2EMxKmImIn2m9Vhz94JV17Lgmhe2
RuCcO8LFULQqJ2NMgOKzEtk0SuloutFMJ+AxaRJXYRtSEjYufFZakm2qeR2pOnm/
CUCmDAf5ElRL2SjF4ZuVJ6i4Ew5+KratnUHexiAHKBHcdK9oG10xxfHOLM3RPkdH
Xa3LVPz4raNPfA3n2libS+rxFOcASO+W0VG045NF3XSxdCbOoFKFo7cAqdxbGFlO
LyqtHzyLVLSZlv8CwSM92qehG1p5izHOEQAk/JdkXEPTUZk4wLWXlFxIJOhrrNAs
sHt6i7rawB/XB24zyd/TOWvKUiY4DH1+xNWT4OKmTz/wyXr8HgG/6PGNHYOL/YMX
18n748qU8nSt33SbS3cDJCSzRs0A22irL4W4Qad9UTbkxYsJOPsolv/iJkZ+2lWo
twSBGhE6JIstIWJtokwlqYFhUDeLzeAwjZtrwGmiXX33r0IL6N9OZGCkMc/0YvRB
vi0RiNG8Rjr5JMlaoNekRqpBIC9kwmmqQitlnCeJI0qWow6nHPaz8dCz//0YQdYh
nQJD2Q9RQRICyfbqSYIAqxtLxEBEJE6wjX7P/3OGxlRnrJL0CGBTNTeKCne5PNcp
4isXuBYRnwis84CWb0OKliac3PGN5jTZFLWTzk97ulFzfc+a+3mIPFLuTjydpSOk
9pUaBHJ9LBu9iInj8vyQ0p4QR2Z1rLrY4Eb7OuAmyYHJkPwJRd5kG9U+FVSCuk8C
gYKGFv0wPHY53hsmpojbyPKT2yBEmTy55HJBa2yosyKA/w2/BECLVRiNnnlKj+Nz
h+4lXPJSalAja6TiaCNn7WmGZCVMDMArrRS7yVW9CtbEOlHzd5yJ6fDxQPMyDT7V
o0lyKWTrtBoarHIbNUYlHToD3p9cJ8LpL3kMX6I2eJ8bqt0i61cp4D/2/HfoZR/I
7DEvkRSd0Yyx6n1E8isHZ2I38I4UxgSpJLi+uUsBE6h221ctKjV/B1AvbmS00hvT
UeX1HB4EUXKszi/8chnPpKcajmOVtN5U35+4ZBfs9mlsprnjdknpHgUuAFUHQULY
iInak1gV4WarhGTJoNlnbyV85e2BLVBmc2LGZE2fafucsNsmYe9WtZCA9TrvzRR4
R2a8KED22RbhiRWyCJ4wonT9CjlV1AERfALBSIxoiqAKtJFTyVTAqDefjBViqGjY
MpKtEb3OGMMS08+M51pNly6O8Fxd3k/LjtBnIxJOJmNrebcDDi7kVupUdatXRwoW
STpCArCbqYxsX52Q7kJiN6X+B4fcCihdijfVrWBFiRxIx7laiq0mFRmrK0cbmavM
rqSRwOAwyLBViio/lPGP8tzai6VcN/JbxoKV/27NEhnI4Fwr8nXJvbbxaI4xggb5
QrzZUPG0sjGge1Ahf0XPFpCZMQExB8bZAt1gJN1JhSuTXcnMtWznsdFW4vTNxujw
87hplI3To5ggMySC1UaA1bodf6pzkFikbSWjGRfzUpMrOhoBy1SJRzdnmdvl4TBN
3i9hDq1wV6ia2Z+WW9N6mKMAXjIRa5/jffZ7I4b4jUTS8C1i/Abb9bheeE8bdj3q
`protect END_PROTECTED
