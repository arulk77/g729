`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ZXukNergEtRrTZiriTtc+4MsEQXK9Gq6VK6/22IsFVv6eHD2ftxaXoat1PdoOyh6
+RsO7VX9V8YQO5a6lnREnu6P0MEKeccm+KFn9AXwWBNPQrSsVH9HZ+A/rg6ZJCJy
u308d255eOhtKomA5rKlgi70nJBTjwq5e08iL3Tw9se3LsBLhfIKyLXqa47JY21l
lkJZV+q8TVK9iwC5P1fQ/fE/INdXsD2LZ2MOcgL2ur/QlFK0qvesMZKSMg/LB5bn
NfnDVhAzo16uIsC4Kdn0jOcKW2dDrvmQJjcCGCRSJO4=
`protect END_PROTECTED
