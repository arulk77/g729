`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAbmyTft3sPP4aphjgLnEOnxCVEs1gTIdcCrndmxzVyg
RbzAIoh+C6q8Rn1uPrioAviOdu7n22m6kAH9Soieup/A2S5k9U27N5/MRPPKXxxb
/bUIe6lYwuKrSIqWnKBHoPFu2btkH/B6We4SmB1gTdO35rzPOaA73KhBn5Y0W/8L
9oLrXZXwrqDhhVlHyVhUKwzOwrYpRk5P18MYeGwfO6g13ezblI3viNUyK52WhDvp
`protect END_PROTECTED
