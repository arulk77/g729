`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIQx4ACIi3anaT11+ShW+1pILPVWuWDDW7JlnVpwzjB4
GaaYAkGuOn3GGung+iHggCP/7mqxm+NsVSQYOR+bqOvznvv6bfjSa+6t9aau30aO
U7xXZ8Hz+EAz67+Bgx/VvByeKFTXMTvEfWnC9Ncw6tbZLIym6KvxfEXErlc4g7is
SepO72ZWdTQHFvLRJcZVmA==
`protect END_PROTECTED
