`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aRrttLnQt42K5tfsZYETPjhO7eNbLsS23Xf162hL24s1
o2ZDz8iqHVbQ2XA+7H3o8Gnn20mCobMO2w0QI8DZbksa4B5/+tZanyXjw1LyI+8J
i80dpgolBeDttt7gWApUPJekfM95Uf4Df+iO9mQCjfoi0sBoFcR5r+HGOwcKRvsl
fJTkkm1+w5060eJYuXorfIvwBdHgO7PjA/vike1sJNGmk5g71jvkjULxmPwGb3k5
hHgljpkx8n/yHX7r1VUw5NU1oVfcvImV5krU7mK1cj9xdVjjrhcLHeid49oO2rhG
VAC9kO8EOgUP3IE/pcZVLv2/Dk2NXChMaQH9E94bGR2KV03bw8RpUmm0ZbozpKNm
/H2+w9WPyAxxIp5SriRl2eeGB5BgcZzvfgcuLGXOw+gNDL8mL4YUHUHEZgB3p27Z
Bnq1cGk84KZUcS6qQAxaiuWQST9FGZPe8x2oAU1EDLla/cSDl4WPRBO0cB1yuvF6
/d4Lc1jqhplidgwFwt+JbXxPvJZuvnU/BA7LjHjDsaW3JLz3EVZT32sGhILavHXe
A3sZaFdQekFwpaoQYDzGlc27pNdsKpiJRGA/3DhfD8WZFHdK0itdB9i11rthsZmJ
4XFfb+X0MiLoCXxuZbz/teNHQiYTfft7k7FrSUbvR1MpMAalppml7ncx2qDwPJy3
lQSW14vphp+0MVMlqrLIhnnry+YAlJGPZgTXMkjPj0iHu1/qYpFKkzODRoLIJOwM
BgD4To5Z5rTdrUOmfzsRTI6UJ6dbEtr/pnUSgglyQ5pqVwEQfzdn8xKf0s5KjyHH
VuMZ4+ZfQ9kisHt2braJFPQ3/Ojw7ho/aDwdhITjX3qlh12evj6iRkvfIf6Wzr/e
jYvHEtMQruyu57CIsB31/0qTcYHzcLuaxm16qar/1doYnYeI/Jt8x98JE0vksMbX
ElEgO8VvcCpR85VVkDkyBW7ZZYdzapCKXWR4NBYxDSPJR3wZHAvsGuNRcQBEdufP
37qjCpFPbA7YZR2ChuXsov5Q8TtwPxmSHHULxajyFYK+4Y3hVg3vviqq0XmXoygO
REOMSVu/S12drXGxGwKnJuS5/jxg85oYMWrm/7INv8V7DK5LVdeuCew2O5ww37Ut
+Ux8P88unYjtM9qncFrqwwBzMIY3RMjA55NJkrNhmardLWmgNa+5bcX3uGQdWuBJ
G2A9gHXjus10Ro8DcDi+c/iitdgpfYR9eUTl8IYHjTyzSzq5co0+p45V20bNuy0n
WCZLiSSRAOhFyqL0D/qrgft88GBZ5MdYD4XJGqj0xNJPP37+N6Kb6be63hnISUrt
0h8gJdKaPxDZzCYP2IOKzbDJXgRKhJLlZ3JUibCGu0z8Bzp5mjoYerlcSqA46Qfg
H0ox//hQJ7rmSokZkPH2kbujY87oZQPARIBKoNaubtprxFAhc6fekL5h4oHrKYBu
0ASw4lry2CoL+zPjm2SjJgD2jCdE6XxTiHidfcQ5vb9OVNMyQUeFZjhoKoKHXiHf
Qm3RtvA4ZnY064mRnEcbUWqK8QoPkWU27ojxJmSR4/hL742KcEOknCxdYziZsce+
ZXiywyLdUPBL5StD/OnaFZG9LtOzirYbtujJuLRmGjGB2PWcHbeCveof053Q3aY2
s6fLrA44v0Sv6IpfbDWuijDcpRmkGRlApJ5Zz6OIUuBshqcLKKMJTobysoayiLp4
28X9k2qsLL8VwC+g97PkzMRnVXW89pdhGx82eLDTHsKz5TYbit2oKt9cQIKgbcTr
1v8+XHpPozh1BYTUcqFJJ7uTIyZdzSLCSt3YgsEoD/+oGibDvWEZgYguLTnbgO3z
IMai9+QxLrazzkMqonNeZjSMqguGHFENJQmYz54bODh9P5KKD9ADRKW2pwgoMeUx
QA1jDoTdBy7/hyo+1SDJUIweS9ID/ML3BClqPhER/o6qAeiNVOVXxxNlilxMuZeB
1NcJ7K6ZkzBx4kZ2fdfNuXOdRYmNVZv8rdOumipAV8l994BTVWCT5xoCKlyz2RzJ
rgsl6a0taEKQaUiJ8HjLanadUe4o2vYhl+qFW9tG7NwnkHQkm0ZKUZFXaO2uJ8Sx
VHsAdpUQFoxm9jbZDUb94DSQSZB0iPqEH4oUrNtQ/y+AOuM6wnXcO2Jl60iA5HwJ
IGRXXdk5lhLOG25sOuHcUYqkpu7O0SSnArwdeXy7tmZ0sDOcmFAEENTudBgdlQNy
WzFkfFjo2qCpZPwCGRjBIZMWPHf1qglh6ZMC5rn9O9J/y6zbw8DL/XP4pBv7Tj9j
YixMcQ93fOa/noAPfI7cNdJsED9FKHnAeLZSSIh6IveeVDdam97k+GCL4wZMV5qP
JytOykdTo2e9KHqLE2f7YzAMuf7F2CN8YQSSjfL5h6zEm6zi1Rq5W3d6ta1Norrx
HVVWzTvHkr8QLLbllseh1yCrhV2CreblViQ1z3sE3eBIhPfd9e0xbAJuULxQZc1+
TSEirk1JL4c4s/mP8LzYjdKKEBghVtAQwQtSfaFZvf3PMAr9o7Cx7Qicqj8jjUNL
W/BftArr2m5E4uK/hMsGpgSUQFJ2FepzQt73YpziOJPd49Qx0PEBtMEK87sxN9P9
a3gEAQ9PR1qdvEOTUJHTABgdXhtRce4rE0neCUBao0XpSL55kyZVC3j+HH6dT3ZS
zZYIY/o2VChZlsIthgEZ8mUqg6VZsW9sFCM7bhbVbV9DidFws6TslUmmw/4toVzZ
SX0iZzO0xpYJMimgAR3rtZKOE2NxnvW66u3ALcsgT50FTC1xmFIl9FfUeDaZcmdh
zEkBRPChK89GsscpYrLMQJINs7uXVz5gNsl5qgisizJ4ehf50bwoDdBaYjQAyraq
MJb/5QwNlKrLFk7+ggxDQJbocVqhccJu+QeaEf050mcsyh604frjFfSfsgMnb9uq
Ub15NZ/tx0pr+d5El1f5q+ckZJkNbvawjlnbflEH2VWls7zRRD7x9Z68y8URleT6
uD4ss2HowpfaplC1vrDd5bJ6uTGwFoYJ2tCHXZyKX5sD04aDBzCslYDWrgu/gzm9
vnX+2ch6kvOrznx/V4bZKSKkU6fA1VBO1zjU3SQ7BAZ6QhyKPnhFKXD0UfjQhekm
PRmS1vo6f0eJXwR7UZGxSEUP7MoyzlWMfLBV2wMGC2isPqvvq13VduHUE/o7u+Vk
6YdV4iviSq6pp79AenTebH65/TyRnb6/+rkF/iN64/xzyyLt7H1ZWEc26AzBZ2hL
kovzfQgTSJb2oo1Lqj/rLV0AODvHjB7bjNqm28pv7u14DfOqJ/Dzic71uxKUhx8k
HERXPFEr4DXkNFPOIiPv5Wdcok4+ioe8D+ShycqWS10OnkDN04kDCN9l2fy2nx6f
3r6+r9QoEoJw+i1xn2t81gQOAs5SRy/gQoIQHFdE51DkiPapW0RRQcJ3zDoFRNY+
8/VYMcbQoeKwoyiCfHqEAiFHV0s1jyBFI/3wahJRZd6Ij67udZsjskoT1V8D3pvg
dT9BbWFWuamqU60Adot5T4rgrssjgigSWaUpJebYMeFUL+9iUvnVN+LMaRAhRtPD
srtg/l2ijXSF5obPLpE92rwTLrxuE/0ukQiZx0dAs2Pk/jy+66w7tWJGX/sLnYaB
mpqUDdJmB8eVKiYItg3QdIxElISQkz1r4rc+/TPr2KHZKGP+JYLlRb9AexhUZl62
xnv/yRYTOnaDR7THJq9pymBGqT9bqC1vqBMBwrSTocXdgAjjQZ/mo4ESY3LGlMOB
nTdAytW+5u+le6xkU98zW0cQ3g9o/D6yEJpsJa9Fijo0JDbAwQACEozJVequaF+8
32NJlHUxu5jlBHIDbozCfGuKQSRtrP2abNTTvPLiJ0X4s+zNoz7KhSCyz0qQF8xW
caaRJeMgy+rvMi9jnvtNCxQrvkuMgpXi8W4Q2o84abdcEVa30T6vRDg4XaJHkqhv
yGjBMQ2jYipcs2sh4RzvrCW7eF12+HeMgTieizL5tuCI1MGeDxz/FpXMHoAqUGl4
qG45jdjCqDV10VoTqyfmRWsxCVHhPDBzVIJomw6SLQ6+ucON3C2UHutw9hQyfTM2
6TErrylJ9jqENC9vsVy7DzEb/4fI4/21s7Zc+O7gSVTTRGnG28dhzT4mpOgy2o8E
0fQbcL/NO1n8JHfR8LlkMy1hsU9wF2upOxR7VvVIV6ZmhtnPKhUu+aJ/KfQaxpoS
JQdU+bi7z+/lmxtK7y1yUeIO7Tq9rmTRO9oXO7IUtCATN2etCzkg+RJyB/RS4E7D
Jk8Sfl2a3T5KbD/yVbJsjcBBeXfDBdlwB98riTUyj5NFvuGLLLrwYOPxTreX2Bfw
UchZt/IbUrc8W3xoSAiI7AoaFvX+g9dBMaDoXrJdz8iOOKkI+zL1kllF9hVpiScH
gGTC9CCJj9XqH/THWXNR/4Srk05shYSQ2vDDX2RMIo3ejh+JY89JsALlIYSJUxBE
XP4tKdTC5rknso2fHDDol/HxTC5chde07UsO8wiE14QQPdLqv6RRUt/HU1ade9nD
CLJfCHkrjFcgJlt3h1jgga9nsr6CrWle3XDM4P1GVmJTevwevahxftBc5zmP6q7V
a7Mk3kFPMWbqWYryAa6MIwfpOHi7FO8ZcJ4HoN6PThmaArrYbUSBgvLDZSGc5j3Q
ww3pAuzgHKO296l8JhJ4VtYMK/IPWIchatucmhIFuRPMHBwTPUBY/YJkmozBvgF7
IfMYR2Z/uwcgdEViDcbbta7eSWvZJsGMq9zqZwAxPKHJ986VKbtsna1cFrPdlfgH
ZI7fK+HrODkPCQg36nqqXRA50Z9beVS91HDU2lmEnxlyrJVLMcVAeHrJWSE+GoFu
0yovia6Rw39G0n6FhIjW2moORGcDxabv6dOrPIjAJYdufEe0TN/7/2LFLm0CPPfu
fSbk1g9nY6/H8ilBmjbrcustvoLqvT5gcAAfPqfLntnY/j23ejEksC5g7J59ZY5q
k6CUgJcug6kQk8MghPTx/KC6zPWeloCFQlm///lxj9+WX9RdXuq1weXDGhRFVyr5
R5kk3WT1pyF76JYDk04xwPoqdmRiuwNyCderVKW3gUQR78E0CnuL4jemzeFo4yjy
/gIRXacoMnDMBS11UUM5nnzvnrMOngnfa/N4Y5kaq8mgRsuPo10nWsjs56zG/bJk
9cEsKlr0wztwHg8hB54IoQ9Jdhro3Pkvbc+oOUiI8dfYFzR19LEOlM46E4In3B6t
Dh+ZrRIInbNSJmpRY8qjB5pkCgbmX1le39VAto1obCHLnPCnrQcjtWQIKkgb6TvM
qLYkeaw4bQMnMv2hl56rZ3JhYdKOgEhqGCFuvzq/8pRyWaPCTgnbkjTyggQ2cF0e
kQKdy94zm52bwFnkCNDXZCqvb5sFNS8eIjp4doIQXTbp+9rOXvR4YzDw6aGX8Hv3
CcoB7oaG2N+ZYGPTs7LDn9GmCocZi3pHDRrOX9S3y+7aGha/XNEz8pgXI5ghQpR0
fvECG7R7LNf2k4ZmB5vBgUxwMEq+Zy9rN3Nf91F06czkNbKhB9acmt1dFPYw6k93
YNTB/exkxRGEwGA00TQxNXO3QC7RPn7evG+TbxiQ2IYFTSAc7gpIobaJD3pht1w+
jr5G+k1ITzCDpfga9rYk67bg7s5ROT3DN/GqijprLxP7qO4XUh/6ISDOm78wHaPD
YGapunvHlD+ZsNJgXX+NtCwYzVzD0GD4ZaJomn4R6PLQJJqILeCTYjOpda03KcRE
i7GjpIDLbMyO5PmRVjL/bipWe/h86JMLYvp80Y/Fz00wVhnMUcJr8c7ciNScDDc7
ZOlLN9CPFBYSs3uslaHCWvwI20oyP2lHpbCwtAfurT/G8nTefQ2FNmpe1Yb3it2l
/q5bPjP9slAo3vZ5BQA03k9BppXUJz79M0VRB0u5M+2bhy3OidFJT3Bw5JyuBVjD
5lNbddKzajxIXV2hOUjZlWMWzdkhqvqcfEX3Gvorj0KmdGFz7Kj2PiUYUR1SeqV+
iQJfiDXsmVAKGG7tAH01jl2gW33YD/qhvjrRf0JSgUMqbuJx/h6so0Bo4AvVUlFW
5QWDkE6i309GBxULCbPJr0taByXZMtrADjFyuJT50JJSi/P+/l6whIGeknjC4OkE
ILwQmi7H9V7wuc1MV5zHKpclZGHjppzE7qceTN8VhVSqNZ0i7T94mqiMHAFv5krr
3wrhOxYoFM2lh4hwbBFRTAuRj8qBRvngoPxTkV2C3A8AqT8shgQc+ugDS+EjUUQ0
q+zFdMsaNifw5UckaDM3ddXEbXAHJKYTlKO32zqTIvwACvMKhHiCveZhBtb92NAp
i2D79TXpg7o/QtXtDvppC3WQob0qWaT4Y0NGnE0rIObvd38geItQNHZ8JScKaV51
FddDansLD1UzqnEn4UDTRkfiK/edp1+YWYC+a1uYiho/eMxCBnnNjmD6YSXYNdlC
tVxgAeC6uY0Xcl4y18S6kVQT3idCANcb7x1ROKjNT6NXZ50cJG1tgc4CrDBBTEf5
tz2l1rJ1DZiRuYidALNZpcbcKqhGceGMR8VX3Fly6Dlv2TlEstB5+/cYzIt6f3ZM
Wtie8quW/JYH6LQA3/+SZDXfGauGDt5cFjktDmI/mikvjcLTfWcK8Z2Edqn20tAa
h4zzYNPfB8Y5T3wse2WdUlIo5pReB7+uMfbEG82cBYof68HMvr34lkh6kjp3BOeq
kev5Q6oE9LVTrJ+FD9BSHpPhoE0BcA1RvufDRTOqLmr+prpjWN5Ci0FTi1kcHAzN
saMCElwtauGdY18p8RMMALwc0CuzTFbEAouebCTykWeKyfAe3GMtwInvcYCyoyqt
U2K8d/1wy/9guXdcPrddImgNI0kWNeyl1+Pa5qSzyoryiTqfdRzRM6TE0Vd9II9s
oBTuZ2UyYm72I/h4vDUsLZaAM55ESkoOm+liUHVa5RDEgjKT1jx/LtA/tJWxWPO8
06aoD2fhcGRxP71oV8V0sGLLTxYPGROKRLRQdqagpEQdSsef4tIhzhg/Jl5DzooN
fNM6uvdFJlPfsuZvY4iX2EDsnHKxjKq2uXgcBwoIVcejZBITeUmEFusox+d6R905
4crynGjxlCjR2eq2Eh4w4kJSejMDyVtjGNWRQjS9mGSfQUTaRu1U5L9eRUFPM0Oj
vphFZfLjCfBhpaVDSWAu6siFjcTvE9CRUxe6rB8KUZGcIPgNo+143mDQQGJ0PxZI
IU4oBkbVmyhPTO5btWHRqN74QyqlvltMnZ0fZmrD3EOJFmheRUfBELjhxL274+qy
83jerS2AKh+6Bm2Ds+B6yVDUnpx06gOvUOu0ogqzYoVDKBJ8R6mLKXMJ0HZQasYk
798Pt7+d3sSZcDkGYPYnvd3skgKSSSu1ZNgex1pYMEVzNnmLi7KPvbQDa8ulG9IV
ObXe42pzn+engxWX9H3TuEv/raPSP3GRt/9rZFCfQ2Fx7fnDAYZ/qpzt+rV76sA4
1ZrBWlcgjkpo7QhLzbu9WyeKsCq2XobSOAXnoEszEMWoyIqtFpPhcKFvHePyNxGE
HO+jBx1jNNSLPAMxXk6jEvnG09nxBnYJqjlMHDYqtw2tgMZeto/J+C2wk+Y6Jdoz
iopF7ye8XpJrtE1poa3DawWxw7OUGkdKgaKSC9p32kxrK/Wp2ePTPTfc2qabiu4X
/637xMIn7YpA2JeA/U+hu0eNEJ+a8uF1ShZFxVdtU8G9JBpbMdc4oV0iOkMyt2DI
LUhLP93c/z/or4pyGJDei+Z2Q8Sk/7L1hCYLtrWLLLuj8kTMSPeT0tK4LCSV5PKt
HQ8sHoe9LCaU93zFzrwc4NsvwZV3CdM09f5ZRiARggwV2W1Hj25UnUrvDHWYlB1X
6TswcMVHhegcOSOgjSbsDwZ/6hzCG3KqN/3JzQ2np010QElBbQ+6vR806tm9pzut
klkv/0LDrP1nSwFJC6p3GDgwAbmcvRPvIqsuEdPmpDOLJFTOv/t8dom3IbIvL1XO
FL6vqUdXTojhst+dFhyDoN+zRyCqPLRV1VNMLt8Z1pLCQImnIGG+LiGeMq/afhUi
BSDsEy2PUl9T1OWrE0tWGv6vfLVeOJPqyjmKvSutVrIzYjS5XG7S1OHHnMW5LM5Y
7h6K5048Cs0R/HQC3M5+cpurorfLTsS+looE1m50WbiJOba7C885ZmRjnWsJL0sX
WH0L77bRLrVmlyCU4UfmJGp4LX/gfXPBHvX6xhCofdpIPX4pVBdH7UhJsiKkz8DY
YcSiwk/XKafdlmPhuuGLV2MikMMx1deUxJLmy6gFkZbhZrYtZeaaddW5b8xuZAEz
/V1shNFTpjbqu3pKNrwr7nVYekZGxFa56UD5ehElTniepqupEqlxvRQnLr0B9N8l
rrTTIrqkb9xSQSZQJBts0b6dXaIiWQRrpn/8KJRUD8WZLZEUQzI0nPsuStg+kikH
TrPODBjOExxu9KDPttaBjwbp9H5ixUzEKBMqavg0RKSC5qeDxDhKKLpShLB1o8iM
Y5XIGEDNX1KaOI3ZVYyJ9biQvh1yK9UfCRicyslYz3jtYuGxmJyRJtLNGvIHE3tZ
l+97fgI1jt7xgIlX8YBSh9L0mX1OB/N1/KLrP/PuJdq7FmLrTBcBAb6Cq1J7RG/o
RZAU4jQBK/tlToy2Qib5NPIeGLUzmxLI4PFLpepSyIANVdFgBLwPpCReuOYsYVvN
4xQBSVsiK0P4Kva65LANxvIzbsce6mI9rmKE1FFAnWKuVnjXQRtQ/o8YvsWRZ9WA
YXVCAVmmClyjdlpID/2s2A4OywaYLvIPyOZQte3AP3FWczd2h+P/cgSbLnyDeHhq
KAuTvKISn5hT1BVLcMdd/DHi2XTkTru1IaTqZvYnsARsV2EaiXiMZeZyb4j5BxJQ
uoONFlQ/ELHJCA+grWtr8DOg/zU6QUyiQxFAI0wqQRxOI+R4pnbHhbLhXtu4yzKZ
igcQQl98MS7eV0Vepf/4i6g91yEF5RrKdOnBw94uzd6lQIV9zdFxY/9tTjEMy3IM
mIR1SwnVUJxxVM51IRQcv0Xf0WMtknRK+W2acSzJxtqSbs+0G9NYPGtDpE9cDCpf
hsHq40/2PCf/+gJkKe7wySxjUdgFHisvLBeOxhWRWXoDKj++Gqh6y7H9PGCcPqEJ
2frKyaKToaX7jdBG4yjctVb1DPluybMM4yCGpAxj4KUb2+PA5V4K5CYEsOuXc2Ci
XehzGYvPAZy4slmald50UywECGBInC5SUb9aSVXQQcKOuZcpaDUTEJCVZqiVTmHq
rP4f6dF5OEv0GaGr26DPSZGeV3/G1Ax7Ls+xPP+QzKqzOUOXp/j8rXJRAq9mmULw
N1uc8PLcP89XAK2fVmT9GARhiJclbk8GiVoomlYoQoAbqqT6jRbZDzLycBszxuKf
9Q1xrgyr3STxanQnLdxwPm2TFf9jU+pc2W5hqCFc4QDNUQk9Q/yocO7NXoMJOIs0
GNfb39pOU4tEgHEkTrNuF9zVpBcleDR/InAK4SXg5+ScDkfiTtGtwtQdERDY4+2n
f8vlvlqFzb+mvICyqMywJybU+TaIAVKq8sP/TBqmUUh/jWIm8OKP29heKMsTTuF2
eC1D7lahLkovU2jpRLYFSYF4nXTTdGQDRERcApD2zspMzm3tmu89E1mLAnHs0t2e
6/I0gjAJDox93uwZRjXFyyxWZPqSEum3hExl+B99VxwnQz0VDi4+Ljz6NHt8wC/j
PhjwuDbJBKRx7N/Nnhv0E1rVcCx3j4cCRkPlxR8TeCmQ0Oxx9bTdzfNyGXxrAPC+
Nzu8J8c065Hrl03AetkXnf11n7YSbYrpSlhYBeDAjC4jtFRZ473xwsneUoGdmWCN
j6QIV0hUeoBuyFlFm/PcwspT3/FfjCnjiAPw11mUsNayJ9b8sf3mzH4s1yW7K9in
Bv7tboNrqK5ooy4GJWgRoG/ED79xsNpJAi8NQtYLvZ4PLGghn0Wu9AZxcG4bObt0
AqkWjl8Ab4QOzFnKQGWm0Hg86QZdKoetlgI4aAAi1duUukLKwgOLk2qYqO1us4O8
kWprtsXWLP3eUfJi1H7SXOxAqHhWHhpxf3tSY2uQOHFs4zVGd/kWZ2K/j6HUqucq
shx47y4j9h83ZOOEiaLlVIRTUejEtrD27xZtFsU6bm0L3L2Pf3nzIw8OariMs8RY
HrFTK44T8AHtFgs/7znRtubiPT5IrD+jPZgrIsrH95pgm3kdGYDl2i7S3u43Xb79
S8hkL0817oDIUkfRTP8XKwcelEtZXv4QVyyUFGpmQ9DCddtQyAUag/H8ms9j/OEY
`protect END_PROTECTED
