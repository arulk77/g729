`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+V4j/wkeelSgXUfCJApq2K6om0UcclZ1pL5vvumRDhZ
8cli8HeSbp75T1hx36t+Y74PJOJ2kYpwZll441thlZ517boniR0A3wH+xq/EGAeI
TolBGZ1JzvwrTXFvqVFYadeDC/CCjOyilSSoHj2shaQLXLQONkxa4JhyG+cjwMf0
TcqPqFYdY/1b+Wv2Lr1cIiDiabxUKbuPn7AVy8Ms2WlZFaFxR3gYIxErl3EJBioo
VllVyMWs5cqUa2l/Z93diTC1PUMZPlvPwdFBuMEa/mM=
`protect END_PROTECTED
