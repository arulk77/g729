`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zcgSOEBhQHn0rw7kGzggnUOJj7bn0xl3T1/o38Z99S9
UR7SWJZAzrDcsRuDsiYhGX74boPbqGSpy3yAkIuqE2BzpvSBbnAa8JPle7L9NXju
HNtoo7qgyzEsrNsaIpB6LTtFlVLWy0oTqqibNBzi+MdsyUwUZqxEzvXu/5oXwEWt
8FT5rvqMODJ10vCpoNMrOnUkKPbsniVjS58RVJ/tbQcMdrupEpit2DXlkx2bWieE
pkyqhITH4SAz8e4O+umOjYp5JdtWcIoiECD9psMdbB+aq6MK7oTT1uDwVtxO9RTG
u0A2jZvCHxCiHmBm/22ANCaPRh2SolJGwGHb3Vk7OZ04rhOFPejS2BlcfZWlvqw6
eeCRg0LuZL3jao5muSithA==
`protect END_PROTECTED
