`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu485Bq2ZfbROkVpUd+EszeFDMg3jYeBW9GNbSJb+IA8V1
/vxxpSylL88GHB1LbWGgTEkRyfXmLD4Q19+lG6q8yx2Wu7KBzp9HOyDBm83JLPyG
w/9O2VQ+vuIbaAixy9AT/q7MwjRiVwYy7WFDbTVcgC5eSH7g7FdFtd61JZoN/KB0
uDZBDg8EEaUH9wZddm0wZii9dU1qutYPf7Evtn5FzO9dCCoXW+bEgJ/PgnlB/KCi
sP6XcGjh9BotIomy2XGqznWrK+xvMSTqFkyGi9sycUxYuMxxFY0ipCbrwT8pXqts
z2eKiPoTNhKtdiZCvtRtYA==
`protect END_PROTECTED
