`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
TvasTpuXIN8gcQCQKD8N7as1hbJfeLhfIwzgpLv9oVi4kC7CInZha13gmbgH2aZm
qb5RZP9n8rbJVX4N0yG3BBUdWLcbLrXxYPPrGQte1oHvK5QsMEANoxW2EZcNcw7f
L5tOjOd58cHNyY2tXua1HST7NMunrWSiU8M+ijsRr2WDpNowo+XbOqAiDMkBln3W
XK5VzC6wVJOeDoMM32pibEane5WP3ybj0cZfZ2BW5IhXuVCiXbgj1owA5YQabLCc
AHUvg8M6OapVPkFAxLCVluLjCeSNog1iTqL25lt5FLIJiayhmuYPj05I9tmFlaGB
ph1/3MBkK+kj06hq4299xYAUlJMUxNXzDRpD72Hu/Hxhfb6/ltGqr9m6FyLP7YXS
UTKZgv38BBMvz7/FU/PMlDirMltNb9tOooDQofzlrSuPzHH8AXpdrjKuvr+yJE3S
Je/ClRA5DqVkdWmtyathoqHG6TaQKVeUBry9vxESegvyCEMFuh6Vdtge7jSeKxaC
DzSOBiETmtGPbnCpOIAtDc3pWdM2NBq/58o2SYbVk3nZgHmQsmiJ+TKTXecdgwtp
9JrLzs60pXCRCoFDn+LRDqEhj6qla5hV1Kzt/iLhEVyNuMd/bDhFiZZgmKZ1JwJC
nIGFjSf/wgOmE+qnj2Kq2DRdPqJPs95vDCUXpg3ndepA3gISdDbvQ0l791CZZR0T
yRUu3+cT1Eu2Nod6qXaynN2DeEqmMyt5EKJOxBrdomcJ6ml1NqghE3KVgEJh2W76
7Y3FzIkdq7DrUm9drabOUXUCWdkNZUJaYWt++VQXJkbHlnZUlPfUJpYL9iDCbnGZ
l1Wk7AzsGE6fDA/e3GH9W6nG7NTRkWLLyBcsmRsXWp4bHdBojOl1WqKm8Qn2wDdb
IFw1crHDQmfNuk41j3MICmAL76D7oySi7snWoX7dwpnJTpbOYDhA79WzFNzrG9sk
r1lqTzJ5pleiSvZOaqphevuO3CtUAzmNUTFHIgZH0+CgH09yylnRDP2NInz+Nxxl
Xw75ZFd6c5r9D6M0FXlIov9WJD4ATdKlA4yHGIkRS7G0RWKZjXYHGMc/5ZSiKll7
ep5w2gIAxKinbVZQnkq9GPfpLHCLqMIhkowtx0CNFgeqIR9FPV6aXuiwN6NwvlRd
5SrVphfo0GTvZ+DQIylc4CbGL3y1lhPG0JuRAwtgcNx4wRMT5lP/hnFk2JbddzqV
sSN3s7hhqTFZwJAAldGx3QeDyE0kE9BPP9rANmZ+bQ9skSGAQVk99OhnImt6R1ya
HBlTWlJ2SoV6dReDVxLepn37UpROHhhusEG9H9crXbj3tLwUtLaW5CoJVl+kKD9n
UfcgLgFxQMSNkmLgRN0NOFSB9f5t/yIEVWrlC6AfP1Nu30sIJDTjwdx4wb8ftARO
93z6kX4lZQVFOxmPpPWZjZRX8qpI1CULjXf8rt5UbpUHM0EnpJ34mQ+DCD8iT23A
oXT5Rp3PDql+ubPoASZYZWMYn6tHhVgT6kDLRh7aeuF2bIvbu/BDj8RVrwJ4Kp9/
RxF3YffBv+006kGzmJqNgcA/km3c3+IFBfRm8PSfFLFYmQsDY+o+87LSAZ5VMd0e
uw1f5J5P6HcSr+ni5hM1IvSvCn5gQEHhG6Vcxj2JlDr4Ss9vqqUFNoIyl4s++0Lk
VY2/udQNIda157njNHdqKD6vL2WC1j/+aR3RM/wJ5gy8bet6vR+JiKPK/J0SZHLl
Zmo6laQCEe4SC0odfjiNNk6jDlK0bPryEO9+y4eLGw7Q8y+uH/jeoeaUgTQoeUgM
gwMOxBYiYgBH1O90rdt6ULHiZiMgiX0S9tNiKqfoz3tuIJw/PY7/CyIJid8jneqr
uLdPdG81nqe5wttSfqlfdF4PWSF0o6CzOJTb6msAteSUvdVtSsa5CVsM44XzCWpz
wvKBZXeZBzh3FVjK8lb4nv/LtZP5VS9upMUzWcmoWyBenA2sLg+k/s3hh1tMvUuE
Jk5BnOKWg6I2VS2OR6xEi7ETr2KLy2Pp2DJF7/DT+QkegY6Qi/d7eTpFXUuVLtQl
ozM5rKO8Gz1pRq6vSq5P7qAHXGCkvA7pKRb6P1Qyj8Hb8k8BCKuRHpdE1opluu1Q
xl2sxpItr1Capbph11WBrd4iRcqc636c1dWJeobMBxV5cpUYIeMOJe0RUBnGEfXY
f34gkS8XLDFSwmQYiTeygw25hBN9qGgys++mLHGx9p1NtIyFLLav9sblJ0cHnX7s
ao7Je9MK9y2DBrelfMjbpF/+4Vo3zIjkjEKTGwZXuMSgBYg2204rhqp0B5Ek78pl
aXvklNZjUHtiwgeYYFAPLtxZCCuAqRe2wbOGImuCgeHjRXwBL1LaVmne6TT0TaZJ
GDm3fck0q1US9T2FFbv7qlXcAs6T86dP1FV0ddWWO9koS9B4ZO50fsL2RPdLRbLu
w/edAcD+N0i88pUuoO2p3pHZlLCPQLVrjrrTvTY+SFJZnSK5u4k/m7EcLoMak5kl
e8tKrLTmci/QkOT9XxC66O45BNJD9GUNWlsea+ByS3jhozxVsTn0Q73X4muxf9El
l+3b4l0qRSN7a6jugZjq0GJjhj+9BB7jMNiG4N0P8BdPAbXcniyNEFSeQUisjmgO
B93e54kbgqy6y9a7Qm/1sWQpg5sWvQ4RJcUYH7+KWpaCF/GrctsefU9CSwk30F7p
ONcKeYyPlJoUTY2ssZ3WUFUqIVv8yfUj2WBPls4+rcXqjnsInJR/PS+zyoc/+pWk
exW0qt5ByupvZ47cjvSPNEEDeWRbwxmNUDXqaCcfXi7XbZV1WfNlnjJsAUvgBbnP
IDprurEdDg48txr0srQK81ENKGri1Qj5FDnejx+BEhA1MHRCAeVLaGhuGUcq7/e4
j2rYHMbaTe+8XmppnL34YCC3+PmqpMRCQ65cD9Ebv3kJSm8FrXtCwoeN7N7+9w0j
jYbBjyw5RK4Ij/h+ydBNDs7ue3+zF/epazERnJL7LmHHscM6NAl3TlZTsTTFewjl
P9pNFOxRL7Gdec+H/DL7fUD0WB8TWet47/d8xgLaRfYgRIL7fi0GfX4ALc9M0EPf
W5VXhNvl8D9YNB7o6oJ80zhnUnOb72OEV9amYnxjpxHj0DbU/W6VrX3XSZ2t1BUF
FkrZKAYDZHgacH9f/z9hjHebrFZB6dCEeIntCZtUF+aj3jOQPVukaGRG19Wlna1o
eRwdev8AVk+fEE4R7oJPOorGdZO2PgV2VmygDhv8tiVoInkmIiAhIvswgVxPVpJ5
UIgB0U8hvBwO8VeD8fOAonl8aBkkK2vmu8tM+qZ+UWhZTiahX5TgYrFR0L72VCUQ
azM429AZEAOFnNKXdL91oQ9HfqkVzmFSL2bancvIajt8PGoaHwpegX2dCQV/ZfCo
2KQZup3+Zo96GDikfJXdMnQBEgX1Ka1DCxxl4t8OqLlWp6RraQD52cjRBgyWxW/u
w4gBkJAZTVMgJdlteqh0fDbEnXAnimxmslj0XY32BZ1m+zqxgCxmmTc9TnuTuGrB
+baMuvOjf1PAEESAJ05IVhUB8hb9t8okgOwl3PRCETbv1jwjEUBs+QCd8By8oHpZ
Ho4+jw1Asx++Sjeq0V5WulwPGmGGTIGdZWKE37kJ/0TCPjI9PmQbkojwUzAAmvWw
WfV9lkrW0kryi5MI4SC4W5m/ckwRaogNNSU0ZiOQJymth8V0SPAPUfOnQx+ZZlzV
w4opC/ZpWowIDIHBiDIFzvLa3tyPISdeqLha6piyIPb7GkfmGQDt4aUXUloG/QHN
EX2jxWl0bb/z+SlrI2QeyOGzdQ+1XX0HhoLKiMhn5r/TZrYVp/wR+KbN2hyR397j
nU0gQdjM2nOTy+wISHrnQEgNfPI0vFFYKFvqIzoT3XJkE5tOmIaTXfYFem7QmA+l
2pq29Ne+/QvYknIhGEu9RFjfkEni+UZyNzcwZ3fozSji4GUUeYusmTC/rlQqnyql
jcYd6fYv/+GE+oGtDNsxOdhsyuJHmElvupfGWariNwHBMwIXs3GfokLhFdBxIU/E
a8aNf5C5Ei5Ui9rQjflriD4UPI52qyzq+WHIdFJC/dZb557mHUV1VAyQJmdXO20s
jzdSXQJUSsrcimdCdESJthFwBwJmMsW6E/ywIMDa+2CLuCxxEWGckLg8pHu+pfUs
Yj1FjmArsQ/vrnaikM6Ms5F+2ZwgLjh6oFNqzaiHZSy2YzbE+DHhgJwEksuB+qdw
VpL5WNSnNdxnKAyltmaftLv1qzA6pUBDjAmvQ5Vd2s8NbqDwUCao4EgUGWmVvYaB
/kWmmITigxG9AKsZioiIH8iny6M6TnwmvtMgjyV8pYElXpIv8613VSJn+3DN61Ny
NcrWLdsiGR+Udv5mzhLnmuNZInFWLT00DYvqZewNjfpjY+RDCjosiRBo+N6VCsBz
fBNvhk9LQ38sp2FLW3yxUninmtF73iRBPDsuLySEqR+hgRqfRaF9pgcgQNDVYw1b
79p0b7A59nO+cTYNs2BlKOP9IfZqsIOMXY9E5yjJ96cLbl0uM2nVGHIW4mGIlfb8
OflemC97+lQmx4HZYISxpB8bGKgwAg6ufuI9pkStzwbNIVOwMdNpg+58wtI7xSXz
luZV7KP1J7OjQnIUs2FH/o9iyHGnt7Yc/cjbovyyp8C44ooGAW5Bx2TcTJunqXt+
pw3Nv592Xy9+DxYS/C0h5+dZ9cxYYpRQiY4v8/Ww0sXTC4Rcm3pCmNMyZTKyms+l
6+dnr3Oh0PHuS6o4x06I/UvMbbRpvfOX5EiWIZT0OHTqSOusO2Su/Csn7Xk3mrNs
VteZPgYmvuFQwZds7TRghRtLunMA3Sh+c5CRg3puJJ2DdQrlghL4bZqP6TwgvoEv
Xj7TbuOuCL8Cdl+BFR7wMmwVLTgGlK/uUFtjN9ESHOvmjIyqQIFQTGp+XAjtcKnr
JdMOubmDuB6QylpH1JyEFTt+2XB97fdcCwRMMHLREhCUbbUWH/PNOWYu+t3DEpsT
l8auMOhzK+jeRoHzwV09ztbow0OEj+JQ//tD2UEZsVFs5DmosjtkIquKbpHrrQ+O
CcZxeoG101sCxVAYGnG5QMSNRPG6jTtG+4FzCWGtyDaPm6rjapVBBE9E3fl4BmEi
/SvDhqQ3FbMgXM4d7LMNI7zoDvPzsolFsLgNbLsnfZRI5O7j+6JQT67ClzyGg0l/
Sjv73vLH0ncPsSGo4nvnFqPu/wlwlpfs3Ry8bElxjcxlmqjhJdgthPgn0Y/XmDgs
dFkykWLl2f6KaLdbZsxu1JsW4+/kRiUGZx6cgXDNdgyud4pgF2h4PfWV12LuvbzE
QfnnMgGswARR3zO96N4qsSG0PTkQu5wtWg8Fs5RLd5CJa8VqP2jUhS+cgVWdz2Nb
b6gvmzYlAxlLEqs3+zzWozAyCngDQgcVd9yNNNCw6bZ8DleZyFLw+SELFJlrr7lf
mhuw08wv37y5R2gcop/Lu0CwS+WR7ewlj/4ll2j+n393vhTlNhIx/KJBmDLfW83o
xirhxAwCbqhNnvRiwRC9pnv9VgcOVU4VxPbwM1auUH7A7ZcD/Kfz6EsHw5wdyKuX
nmezrAxswnPQQg596rKIBFoHaNSAp4Rz5U481czGxUGRdRt2Hb00KvnSTk3xdncx
tIMBKZGEvbz9AdL2AsFFBWx3LqzpCS4mYbdg6yaHrOPCv/eRwsU0UeBq/QdkYd5F
94vo0N06pdBcG9yKw/xBRyy9dxDnfG6jz1Gl80uI7M26ZqWgCp8gE1obcGhTa9nk
77f1EEYMCCHmM+fhEXjZIg3l1stQBkyMol5Gi52tgp53KCycqSKmZeURmSmQ5DAI
Xseq2CSvQIV1HG2ukrEGIKRQaliXQxldPWANdxBas4c9c2CHUO9LBvkzlsH0aMRe
orLUH6NOsyn7A+TRHP+SAcmEUYjXvLxWEHmWe5Hf1deTJUKIEzuPoK1GWJGp0ywx
yauTxjakwKiPm4y8EAT+bA0UF81Ij93mOprPg/ZE/4/7rumU2oSTkxJIL1sn2BBt
QsUxdZkieWAG4/9n7EMGLVmHmRx9FuDr3Ke+TZD6HMsfikTPxvFosnKrB+DEGiHi
iWiaBzS7dlk2rWXTwEQXS0Hg2kHVot/Gyfyj6lhSIzSHTcfPX4J1x87IiCREXm5e
XvkL+zSLr73sxLQbmFFVOZU/yjf4p9jsm+OpaqfG9reXAUcMzOfZa4N2fPWpBzLn
C9gEjR31GURZTfmnw4gzEErEDjONX+qy41doVatpKs/T0Qu1ob4q3gGC7DSBd43h
gexjwvs3nma2wKzbAq70psxJhn+gSfsCDXx6aRWLOjFCFvVc3410lEjQpFCyehgB
ZOgFMe/TMJ8Gc2tll2Y2b9iIvzhK7O8lJidUWV/0MQJGjzZ5gBrgz5QJZEQ7aHPy
yugIKGoyCIo1JH8adQkIvPZYbvTd/6xhit+Es0Sy5h2zr7tjLqbnacDybUIyRzMC
aetO5WdWY8Diep+2pYcJ9nk8bGcpW0LwN9K+8D7wU6+fmno02csEp/tJtrHgUZv7
tYQjX19EhKcyrsoTquQCKMP/K3+ctTyWt0sDgZITfuYdp1pxhSNiXimVAuNN+SMs
nScFSTHK9AveTKZuAqCE4nQTsTNyO/sUMC+1c8WbYhGN82xOvGwUmBQV9Mhq7bki
rt9chwxoe2588O5RVxed4jGq33aEyhwXTK8fN1TBJQz3xcmlItBgkMe2ECinlmTu
IYfqq9ApC6aUwRw6NurtJRVdX0pY/b8Rh3rO0ey06en99RyXRdxjEfEiI4xzD8i4
9+AUasORAxxrCob4iqKnPPPSrufAYh6H/p2ZT+QAuW7LwodzYgM7C4EUJJUR4l61
TsuwEJxjShILobGAg9J4KGhFR2W96trv2i5RDgVjllBQB/yCPDXLpGqYjZXyR4YM
cMdsmvjXN9lEerOWBoPyi+I/58bKfHQpi2a1RfE5rxJEt25CbSAvOmGqs7s/+ql5
TdGizrdg6sHr03jlYgSn2kSgQfBWW5gFylMqwM1Qh+OY9zgi+xlwwNGdoWGGsSDG
JF+4ceCVM/D6/JYPco+gu+oyG+krrpkBl7l33aFbya8Hqbezd/aaI2u1i5IyBEws
HtGEU45Tz/ojo+25W+g2o47sfsWX4zWXtL5vd8ZPRuCNpsqJkLCmaJN5sG0lmEyv
Y0/yVWqclbYH6eFrdPsQF5zrLruopiqqAD6GevAaPy0QmYcwzKgd9aQltEIfeSKM
LScoai0GA1nSr40SVGdK8pY6J/tFGE99zj+G39Dngpzm14/7MgHAJNQyLBmCktZ9
YEvFrfkM8aThWfQEPwmT/iFv2+v284OXTWsC1p6i2ybI1hVBSJpou9n8gLgVw1oM
X0GBU0ojUfrW7OgYbJnZQgjj75TJ80zz7pD9515VzosZAO6J7GXVPJhYI0/CxFTt
3euhe8GYqryFTsK7YRq9xwJotKiOxji+dNXQC6fZlHc61ydbfLdbbXFp69hrAsqv
yuOA54aSWHPL0C0n3+3LnZd2Wga73YTtwrjp6IIKMwFicRTm5CKOe0MIzkX2Q3mW
NlPrMuts5Z49xS972MqgV4Iwjh3tYZ8fX5Y6pU6fptFp5mZx/YN9Dg6H+sVSkUdk
UFIEUiQwJS+ed2zEsEJGbMOkYiVOL/pQHS752F+sPTkiG0XzKlINwPqoojQ34ntz
qcg/6lZL/ZmUotL+x5syIqROJFc674Cl4xqeOjMKzTQgwYCoMMDT8MAOweHnirfJ
Bjk2GZBOSrw8ywIgOnkEe3A343DaoWrs8+0LOgbOq9cek1EFDWMP1VD39pDOz9p7
A9nENm5Ivqjd2hp8TLrJvvQhSiAkVJElE7v2uYDZbeCXhzZ/F/zWGrE7WslRWTSp
fZyPj7jfRXDOFgfwxin21b4mhvzncPzZDmGiTA9BLZ/LigVSSbzoYx1aOfdwQ/KG
BpZoO8yz9XgZid89vlfhFzUDZLpR/XyTICKhxt83y4IZj//xOUpl5kBfgTsHKceb
LdfFMaH/dtMQpb6xlRrbjccqUu2JKA4cd7jQc4fAhbtG4ykHN3LcrnGgKghqESUB
jXL5RP9zWKQVNj/SYE8pxaZUY8w9n7s8L915jXsTQeu8OjQUVvdQ4EQlbjXQ36ER
3DHA1GxO/x827YiXeuhHZGP9enhjcCZa30494BKs/nxkxFBT5AadG+0vjLvSefjI
UnIIPSkmhdiBVkgQX5DUTc3mzfZO3926whRxi0aKaCpfEawY0BslfQlt+9m0206G
J2t/xd3i1XIKvI3f253RCXjTJPKUvFOvRgEo46Wa+kA/JopsLGLy4QVvhwerpoc8
HAldJRmw8DGDc5QtsReCMg6DwT1ftWIdhnM5qRYqcPs28bGSWzR4PKkMhRLPQOcY
0VCFQcp/hKVqf5LyilIDClxr2wEKGOPyPgxcWSzf88imCyVmIIMx14+Ks5ZbqWCX
cXm+KIkLcLWGVs5jzlEwcIw3BaWQIV041lQqGCBiOvmej1pPqcgWcfMpZweA1q2X
cj3+DhK63YjUX34RZ9L/m6knemZJ3+Q6CVStqFWo6Uq3uvCM/wl823HVOnufTqJn
KbliU0xGu6ZOfG6dxc+/ziXZFS4DZiuudXjPXKSC7txCyTccPvRAlzmKOz7xTA1h
6icGugvbEyrPFRD0OgmJrVaTbiaGAjoPj4GZn8x98+MU2M7MdUSKuUDZhQAkLFD9
L5D+inOLQQ9FLwjwAcCRgdkQLFokeLuComfKIho3grhahVzpzm58VxBO77SQElFO
wTkwqJb7DYlfJiOaPY088hDkBfBKPTMDNF7EPch4H1DrrHGIok7KekJ1LqvBN8Pu
bqjQpm3WdrnLNH6GUMqoMkcxFh0zdEEYd6rSnbhg0822WZl5ya9TrZn/zMrW1IwL
bHqrYyvm8caHtQOTw/wGJdm7EoUbDnMPYmpuux03udJ0CLoR19WZ029uix417XYy
gxI+Pn6/0Ef1N2pyzbRiWs8itxs/lN2N24bhBv9eVAiZ62XRXRhWMGhQ8LliXG0J
THpSnId3cOPKZ4p2i2m/KE3okuh00x8uey+6OEQVKmmwmBGvrMDHc5T6pzbFZ34Z
jA52SkFnXQCw8aqjMejY/gzb3TLn7+eMnobUVTEB0GH+ApZyZ47XBNzBAcChVIvt
bqAaBP3JvFlY7v2A1Zmzg3E5l8hGP4hTHplyaERyruimC4MAf0OdNrGUt+/ZuLsS
COJylJ+OFunC+Pb9RPxedPuPnfR0gJ9fON0alkRC3MPXV8tlRDDspqn/9L6ZrBPj
QivlxLFCt6JU1eqPFVj2JW/O6FZbYiS9RgPtjHjoF6YLfdlK9aoRqisRINou4Jtp
kGCmibV/u22P+hm3IHl4If8DkbXzyJ6oBjF2fmLlKfq0rkSqrrA26lMbx6nrysaF
XG3wLm4Nz9OMdDDsDkVz+SfMVmAd/o5ePqDc+sSR3n6/WAPawgJTOpB9+IX2rK1K
eC+9emUMxEGW8AKNDBwwG9GXIYjNFMfg+AWARhtqrLE41QZ2TTdmSiv7sCSwGtAe
YSu2o89u4IjlIrJM2s1m1OhveYgnUuCHdXgsgdLe3z4eI4XZhw583YyhrifUoF1C
lzGwn7WhXzMtHcTbX7UBFWszfBQOQXqMZ82z3MJvw8fqowRdm2DcRYq2+a268udO
bzberqMwE0toIECZ+mtI60i7DE+O/lor2R2V8gaq7h46TFScQwGh6UGrOtbk8ZZG
rF6z4LS6lvy/Ud+QavLgKvVunen5K32nWElkwxT+EXZL4aA4Q7AI6lRA33GRAAwd
iWAKgHnRCCpGZTVj02MyCtlZmXzygzWNPtruRryy53yWexx6p3iyBqGy9JFqiW4q
/aWJbNjd4/91UA8cGjXKZxi3McSLHh2lKjWXdd5ZtONpeayJKwfwZMAsbJgf7km7
oV1QgxHHktNfIpWFLlsOdTQT7MBLO8x2SGjKSajXM4BNHR1aVSR7mWdF6++SJXPj
RFbgbIr4DQYC3UVTmxSaceF7NqE6VuRsnXlytmm0zvBW4lc0UTJn6gvzKf0IasPi
st/murFUw7d1diJmUo/FKb7OwHmU8W7uEeHWD5pgF0QF6Rw37NZRLIqkKj8KMwU2
LRc5nsnE0ltiKvwEreg3fjmgEq5bjo2CMOFEdQNw/yA0U1tahOXfSQ2LFDJEheux
/tnuh1r7aaGjy8qRchJmJhbSnaf1lIwOWuHpcFaQLZvKGRlkAjZ8hmiJ9YJflVRM
nbtt/NdVEuc4RZ9kZfscyGJCdQJecLUGtrKCK1SUUzuQ+jZZ21eaeFToCP+gNbOR
pDRn8gB8Xg2mvBrHfYG09BVFUzvUD65lFR5mInuWIaYBFAO0pO8nKjm7dtkN6FQN
410L6DyquxrW2Q6ceYB4mDSrUFgE/LNcygy/lHETblpNH+t16SPaAV00v3C4hrac
4ECgnjU0iLQrXzxX8gcNX7uRsCzqMc21eAbK+n3jDSYgseuJee8ftcQlY1krKQGs
EnB10V1MYMPZXcYxhOI+AssU8ie9hNO74VkUk81yc0jRUvCMvJd3mT4G4DH6hyz1
x4FFGkRBvwxLIZty3l4bwryw2lyblt9ysAsEbcTrULRjHP3Vr62Fv0U1A7v1OvK6
kuRNZY1RW+ohUdu1/mdMZyM3x7NZqEjc8OhA/4EG+I38sR8TNW5KPbU50UEDY80E
rXVV2T0bSRpZkvyXLR9wHJkUT9eYEqZczWgsyCwYaM/qrpFi0svnB/y8WLZdhRLE
pjS8kQJcOApPYpuvYOJ0M0s4tns5DTkvKCY8chS/H1eEBINWfzZS9sqVoY5L791E
dCQ5MqBln+aZKeDBkV0YHgXBib4NQtq3GCSakeDmTWwuk1s9cXfwUxmgUpyz3/LQ
MPxFZiT/6CmlLTsouavk0lF065NcNDgFDV2WmqccImWWQfQIXz9FIdtvIhFjMYMI
8AvE3+prLqMUxTAH/S5w2q5cS7fp1BCAdIEkguRrh0G9LOcYDhxZk8wsHooLfKuC
xgqYQS8PsRkAAqRJhOGkOlq6xmKBw8cndVg6nLrPVYJ7/XZTz+PwWF9Pb7wtZewg
Zu3u1AnMRJRb5+LNbVFMN/X6Vvw1CeqFTmXP7skn8pvRczsXz/UK0haCnx7CsXyy
aH4/Q5e8WS7ZUqGMygI4RSpchVjCJDSSgOQXx0sWOOmxysB6hmmm4MGNCI8M4jZ7
/HT4LZeHomu2ZTIf7gMV8INtubNROcuP9Kl5qUNQ2YxUe+qsY8YDeXtzFsGmNQJH
4YpIxuyLffMwcfHG3ikWR34HrRiuJ/txS5WcRBIxS816ZHUY6q/dYpwZdYOCPPPh
fzvjD6dXOJhnht37WNVVS1dMP6H6afV06qL9fHfEr5rC3gik9TWVQ5T3KSdYbSfE
OkRNflLrs4VzfOIx7K8XjqWlnhcQ1Aov2Fp+k7PRn5krDyuw3EBwrl8Hk2mX+wkd
0TtoXkTYymPtgdXnh5dl8R7twOcDMLuQWeLxzLlZZEzORRE6A9xwc+D+zX7Ko7tE
4M2EIfLnJrPg3+YtDLT1SmMt/lx94i2L1icNUPd3GPoOXZHepCFYJplumiC1Qvpw
eWnTaz756oqkrHRJlfieVR7xqO+KcPQ6gNL0vS0BbeFn1NPUpDsUI54UanHcLFKD
mHpFN25WcZ2IWOu7x910Z3Ll/oiG485gV0nq3+mPBWpAgC8shvjJe35/8rnvKOmY
IWFrcV1zwKTlX7LkqTHIJyP2UvOu/HfeqIKvHi8pTeAVJhKdWPMeJm8zUiY0emAb
Jk2G+FYzgHGfW1LG287OEeQyf9XPSQquYvNS4KlH2CBRVfKXHBgpxfRSU3mi55O5
QsCZPRF9vz0EqL6uNNBYbGy3tm+UqIp5b24647Pr/J5qtQdeFS5sPIkuKx2bAswB
NJ5NiPJfqA4tDiKBzMFgfyvgnyeAWRdx74X7d3ehj1qTP0CQ9qIJZUgiY9pSs/Ez
GMD1FF6JnrdTRlcAP+gInDdfQCtCaxJVa7Qep/ukTw+vi71DKsNslOacNU9HiOMO
elZ6gCAVqwS05iQUeKy6mZh1ZXEMLBZ5q7sYBk9oaXvE53s3JgsS7z5X+9Uc9Ws1
sXrez1Z/YKbbgVcq4HynaUSx9jgvhTF3uSA8tVJYYo4CrySpR657DNexHsh4m2nM
7DtzTGaFqWwgH9VcQ9q4Bu1gSYO/uwhgljouf+g0wKpqoQQIrejsoolj8KkjSBC0
b7qD9ixLZaF42PGfxyXrv9JKHU7L1B1dV1Wp4DSparrSdmnFwZLc0r8V/umNxhuj
HoYsN2nFYtkwRWXjWfaWXwu8+JpUO28Gmje8jwnxfVr+6fFcPfUOYWbBEGjtAfT3
hk7+uHoZXivkX98bD+Co4Xfj6q8gG1HONtz66feG4E2ok7uwSNpoM4BIjTGg78cg
8llSOxy8v8rpv91SMkbsZWTe6wSVigY3p2dK20HR1Tj0KrVP+l5i2frPUl6TC418
91QiNvZdqxzE2kzQRJJQi8y05zhk+Pb8RuDCNcRHZBJlnmoN9ErMm8ntUA0YazNO
WUDQh/qJ03N+koonbgEvCRpmn8meF8GQ7+5hWppcEVG7D5LWVOpCDEHn0La8qpNH
7yPVjyyME/XOb3tA3LGnTrULpqOvBY5B3lytYhGcQ+JOYrvfwl5a12ZPZZwJmMX/
igoLmogL8d5INBGQtXmyfqJwMX2jvqUALpHEq3oytKEr4ayFN04PQV7zb9n55Wtz
13UBwyLrU/1HSsq74V/nYDKWyxIOwycJ9Hc2J9IHnnVK/jDUEUuM/Gwc8GufPgB7
CLDNoysFFtPMbhtHQ3hLbbfQW0sGJ3oL/TBWG8EK/EtDPKxIJX7YzpyRPRBpjk0j
VdXB4NLVSqWoA3/TuLhJlTgjnenFsjwcuQBOGDRB7op3/NG4dvDMcI0vDl5D3BU6
7sZySyOxwVBV0PCOD75GkyW1GRSAYdAmR6M3lE2BPp5I4DOb/Wo+6tjfOAce8DxW
mDgiin6hNvIvHT9mBmHWFMuggukOlDY+k/OQF0129fCTAaU3RZiuXQ9c01QKmo19
7wfAUVUuydWbPcu9KjYvveTZyXf2wzkwBTxXQKEqOSubvpamMf/gy56KpvQ3odJW
9Sis3aLJNB6CI2wTYGLiZhN+Sn/qDqzWnFNjjrwueV/o4PldnJVV0ShV2bz8CcDQ
SWq4Y+KlpZHc/R2Xj+3FdIZt6tH/+VTl4Uou5a3SfPFLluNV618FcgT2E2JJL2Ln
PHgfWavIQkAXydezhIQW7BenenUZJiAt+8jHeQaFYLyTz1RGiPVWbUMpSkOBQdcI
1g4cMpMC0iOmuNh3qUGMItn7Hg9a6OioGfBd/jqPxAMgJgqNLYlcwHAmUynHtTE1
bpXmdEzW7Tqq7Kmkyezxy9rVuaorlyaDGC8lK1boVtb3NJfTKxrRBepisIlIKgVT
u+yFk+8LGRHH1izPRLC+dFcCUKKYMS5pDR2xs+j4qSRdpy590Yibpnmnhj5MCtqH
mtE2calRL0CrKIAaiHWCQvBEufD1ptZlWMNIgV7wkCyZomipRopQ94laGCDY+K9I
MZr6JUZmzLSIOUQSjkwrldQ7D17CkCyq99awZLEnzU2/w9sEQAXO4bIocLQ9356d
QNFYpZluKDoG5xXwbMN1jPsoRyMuhqMUcPequmbHC5MYNR36SkzpztDNEtvZ3yHn
8jG0d1kMh3t/8W7BNN06UUzzdK1sryeR2TmQq1QZ7aYczoq72GAkxNAJ0rJiPQpQ
Xft5XCrLzkPCO/rX3E0f8bDumAmc+eJyEfP1/w0e1WX95A+EPxgyIHDrOPn1MrV/
6y5lSCZsVgfmYaEp87p7KHx3hWyI6VPaZSw3EryxsmCWV6mqFJBX2NLNIaGGGpuf
zaREMAvwjdjmJxAmOEj3S0f8GUEnBlCYzTdZi+xqq8lJRmjqsCJ/Fgl6XMKgZ3p5
MkfGHzIurOf0yzIsPnp+d4tfiHbp1H9BifNpEyYUBbHLGqjhM91aHFiL/s7dVXib
eomeCleZfkhwZheeTnhFt9sx/zCDT/d5/9bSrj5bJiCCaqOtL+FhIIGw9nDxuyHi
9YcxYH8Q9lNhbrGcfRjc4o0jqw8reZFdU03hp0Ep5H9j87qiqb5Sst9MBO7chlFs
knjJd8CMIXRwEUUVFuxhjI5WaIemAvQisuNHCwKc9V72ssuztkHB+D4tDuKosVpw
YnLj8u66e7tXY0jR9Jy2A/54HU5kDfd4WbhOWa82gBJ8NycIOHQfGAv6Ei8a4a3v
kKhWyumTrIU72wFXGLLmXsC868d+wSe1Eg/Wo/gVsEwIyau1U7RBzsJpekgsvTN9
9lWMScL9YJyoJmmtpL9McK/ZkzB1jVHBaoxMToiMzIQbnTJs6uQwXVQiIoR/6YBN
1+B5WQ4d5Y0zJY6yJO0QZEqK0ld017XeIw1w/Z4qDru3VY7x6VZzHIKG1efsh5rW
3YPtd9QUmkZd/cvtaRW9X2EmeX8E5I73OZBKS6FVPhkLJepK4odGwsNKy7rPpT6f
57uTKwHov/H9TSNfI3QqsGNLsqJsVZAUhyCUddxNFuTSoGh5/NW6JoCNvzf823bd
w03TdZhZEDT3VCT+DhzxTrLKBVjTv+x78bAyhGpBFCqN0T5sw4MVFR2kA6WEv7TZ
CBGCpsjioSyn/t/MlK8sxHt488mpR54zedT39Fn7tkj0QGxDeVftif1+C2Pwi1/L
Au7mlb/l889UgbaTepR6Vncp/C/E4wydLyxWY0ZXs1TAmlFKTuKxGpS9JCoe/Ygn
kLEkiEWIQzFwtZJ9Ge07BWsBUpE6yYJLneooiwzUasgzlgOwcAKZVkylZQBZpWjn
sPqIzuROBRXOKajuZbL6iVyKc0OehcRI1YfXOhECHyo0ssZQvuQIAM3liUcz26ma
EqU3fhDRouNegb9uE1VjPqeVFa6lP9sAK2TcYZokpO/HvzCGP+leUafjd5vnAaWL
22ERNrckoqzvTqSNIvU53nJLpoukJm/mIV4ptV9g2aIh3BDBV09GiLoJ0Wmaqx64
gXwgn1FM5dihCAGcufQnlEOi0ZrlOdGATOg5HyiPiEJQKVtbad/Xf5Hj6DKhitbL
GC3RyI5vh1hFvYoQyYW1MXKjoaNrvRxJm9E7A2yd+C5A33iI9SxxukG1CFysnhSR
QFDu12RerFO15LZoHx8HcuxULKVWsi2dsQhp2VN1ndFRN7okbGtEdtWIIGsEfyOa
eFZ/BZWK0hfHfo98yxhg/MgGGg1G1zgiMQwUIJocKCx9ho07md1eBaXwiaRgUiZM
mnk9O0sot26jScB9uIUBbv+lp5MVSqveez9Ede36oFpr63jJWdiswGqmQ6g8JLJ+
ymgWT3ibGic6LJdQ7kqHBOrZIPLdsFGvww/vtzBPMI7wp6C/5zdHw10edN5tLHxh
MM4i8ZEuALiwl/F33BHF2O+88yY/Gm8ItbgrrSlD2qSbfo0MWS8geIu6mdR4fNVi
N723CV2sghWcEPhO3+JK+Vi3X6v96G8uFveUwUZ8hDXL2tQUvyT9M/3DHY0FiW4H
AuXW7T24otGNVAbP72OBRqxVzpqsxYNcmnCJVu2Kir5z8y7/YFKSgpWfIAwq3NUe
wIAKmfgjJj5iYiweNZZQa9WxO4OI/5zTBdeE/Ah8ZFOzpVE5dZ8BodY1mWPJVR0K
NGI5Qh+UDxV8SdypY+6sRvq2pr8J9Gch3rHaSmyzY11dHZIYHcYxHfOzVHQyG7qN
HlI9lIm1Cs+hoNY67TkXXajAtSdT8FXwi5dGBHocwra1JXYUf0sjPPdgofAtzBEa
OGp3JPWNopWOW5RqnRKFSthwVdbPotkpj0/Lg0j39RGE5sRAPynVn/uVe0cI2I9G
40m9PxMDtVk+qg7cfpM9TwlxJb1djT/xDq65IBELmifSqIi9R+tb2hVdr+mnfUtY
1JO/BDeZK65zJUCDcjUmbrXEdlzKqFIRpzQaVqDlpK1TRCKnk2jgap+BZrqGEGDH
caV1hiCJQmVeUgwjtrY7KkfzVRWcotr9LfV/jt1nRn9rwaeHiEPGLS58HfUlkkKa
hw69FFJXOn1XeI3cpcOPkRfTuJhzRyl+44wOnhPd+mXdq8D3qXKtSpvopebkqBqa
iS17dLk0rMD2qLl7t3ikc1/tpvDGd3XeSEK8UdCrPh6KlWZevnJZrNj9Qo5seS5U
QJBZ5nslKAvW9JP0zF3PtUBVQeYjM7nTu512GnQFNCurwCG+VqjhDcvqKUUrjZKu
g9kXIbnF2yPoJneqpOnEIPLLb+FHzolLqho0jGJik1ZCg9ZEqNZpKLKOTISm/DSd
JZd7/j+nOEMO8mx4v33qkp5XuGU4xcTrJX1NhY9Ocb4LNVd7Of04Pmm6EiX3cizh
nwddKb2Lm2QV/IUYzuU7EARTO9TiZ0RqGbyUFTUSMcT5jL8msYCRs+osQPN8sZZ/
tSvum8P3lrA01E5KWDZ4AyN0vOjenJwQTzSJQihj95g7ea1zArJL0OgGva/T39PK
bX1HeOKerNjIs2wR+ngmV7qhXiiktug77GXtxCITQiJ9j1AVhWrUP5cqlPtF3lje
wx0vnnI0QC4HRsPV/YmLLi3BJ7uxqCzY7pJGZxh8j3dwn7Bc4aHmskkNN8n3UIRY
sszRPTTtudY4MP9WuP12UdKxI3Z1iRkf4KXayzlTsgJH1BsZmCTcZvXnAJm47/S8
yaJfe7pkPK94vRMG3tP5t97PN3PpBcRbMjQLAlVIabLmcuwYGTyVILUUTB587Iwk
YSdhlSkRrrpF7bJ8iARk4Tk8eHF3Pu2aWdNDfGv2RjN1+qy1zN1uoDAWI1yegBhs
FlE0D2iXs/jXdaJMf0tapnfDf7yX4T7zsDsYj+z1goIXOmozIfRg51CrZuKTYFjk
EQa1eeSf3sHnzSriR/TyVZigKO/JH39xVdp+ZADGhS5IdABAThlMrufdDPPmiI3O
0tCpZWrG81/RFo68lXCCpyK80YkpoUDfT6Yu/Q5HCnNj8dyrCp4NFne2A9r3wevr
BLtb7Emr112ikZZYo1BmZQxAtoVzscpddm8JJCcIs0NbDqob9UiL1WPX8KSzSUHu
tiZqDjbHDa1B2t2T9xKtsla947bX7MrNEJXT7e7awBGt7OnX4fZQwi3ui5d1ngK/
BmDWXylCobrSFsScEUb5CHJUCTOYQmCXfJ9dhC0wb6n3ZXCSN99Si5xfdxw3caQV
ZNQ4adftCuWCCdl4ualikURp9FYIxDCeBIMuFF14U+cv6ViFJkrZp8kgZzna2qrF
JFIFgLpql9i+dB3eE8h6ksOHHjB0+qjbkmmk0IztI2s4e47aCxqkHJsWlt1lB/Ez
AeLU2Q6G24+cbAFugPyKRb6If7XD6+UIWuEFPor5jopm93nSZGpRaQraZU5ZzY7O
nfKQbeGaZOZG+1ZOX37eIF9I6ebEYUPWSlxC6z6d1rC+YQWw0wnFXjdpYGGi7HSS
s87/JsIGq59JEmCUYyVgrhOou65cHA9uzr719vi7JTMqDIOFhj0CmrndyreZKP8I
MsCD58M0Zb5zEBQITERTZ3qyLO0LUYBH8BazF3eVHybfCA2ohtGSM5lfbgULjt/C
kyjKThe3MiYnptCw+/af3IFe3+b4B7pRD8muEE67YTdk5HN37CLx2H0uYhobOZlv
hUOOYFBl3/QVq28BcjBZhl0/FGEhDxD7uplBfwmMVw55ji96gE4TtdGjGlaWmkaO
YFt1EdfeP8AZWIbI8g5PPbFNHbFTchgaVxVW/vnnIngaCg7qTM8pVVcoQhP1/RTD
mq8TMt4yl/NeLmA/u6uinen6y+YqQNkn1+7Jjm4M547kBQN+brJiT0PwrlWr5CNJ
pkLqEmwzmapar4wWUMH82O3SbISI/dyHf3W+ypJh094mmSG1pZqY52AiffDeROcH
hmlbh1MCF1C5K0g034jXDPiY7/SdrW48d7VXV78JtA1P4HUo5vS37oPnqnFKlc+A
Xd4GoE+6a0MoiBLQs6iEewxqwh3ivvD3q6m9Y5b3vSeZsLOjAko+4Ji+uBdvT+cr
peb+phN4VzffKeLBrhlt2+HoFRDQlQ542PwLTCF/CrEQNQA3UB7I94+p8zMUebPm
nKMwbBaUtfYWwg995R/7npRKtlqJ6pCdSqNvo8uBPHh0EDCfYlmYAzRulEWZinA5
uGKViJMf+V1W3wOC4kV98Kbq4frsvKsYm/9IYqP9UafnRFd9A+P3WDOC5yaLWAZP
hHs0qR5CvyLaA+fkISBco7al+00SzJCYo39SvKUdUJ8ta2Jt8ZlyxkD6mt5q6LpF
+FX2lAcK4/s/FryA0yfDKLrhaxBi+7ii9He46k24YbKjCRb49FLTLn7DCy4awC0U
/chnP7mMGu2HiFdbKL4beI4m6L7pYa01f55IL1Nui/blzOKVF25j93c3eKArV6rR
KTLkVSYKgkm6MlQ5ttU/ZHPEJiz7oDLMhnWnnHptnuufW/JEGaOHEgghK2WYQTan
ix4FGU6ULzkgzyzLCVEZAot2Pr1sOjWxm1VDFOwgYQH7UFG8f5mRUhmYEd5S02W5
hibkXuScI7kvlugd5jutAfjXzerB1rox+9awyrU40yPFUl4jt8szdK6bcE2+FBSM
2kfkoXFaeG63H1XNA8uaaoEKBaz958053k7wFV18o+DO5ACx2jx/mrUs6CXEzvIP
gNHkZDU0r2BzadjXJszhMj0znlGzxqRCgh51MEhJjhtDIkYjghdodKG7AqIuHaJ8
H5flAP9sw3AS0yXktmhUF3FQLVhwq4OJYVZsET7n01A2V0WMUimyJ1gi5FMapQvP
WX3W3NXqDMVuffAEvycL3INTCEOcDAG1hINkLBrfs/y5qmdeglLd4vtuzO64/YlV
MY+BmsAVS5sIm1pXUgUF97sYWiugkxDD9Zt3qvpNP+KBWWX0yRD6Z76bPcd/qMKQ
t5TEX5fqs4Ggo2uZfbzrZn2CaaDiROWRxSFyJjrlNH8Wv7jMOniDSR34uVB2UJ0u
/h6u8fMaCkt5cxdDMG6DFRYeWhgpTkJPouNpA7RHNmi3zaPsbhMPvQgMGWezxoUQ
vAsS6l+4t4+qr8XPQFCdR0JW2mAfLF3oz++6nhCJfxp/c700jZ9BAu42Cy2NxOHW
vf3uGm7PJKWBhH4rjO299NkwhkqjHPG7uJL9yM+poQiJvGgAa6+KYzUGDwIs2MMT
9Yp/3fw8qVUlKzj4WOTP/tY8vAB12Aq4beGfalphQZ5+0jshFvCjmD1w+qomVocA
ylWkGuLAMTSV+U2uR1hUoAPqxRo6ogKIbGWOqpNiAvZ0/1ll+TZPLc61JdSunDEz
qZwNXaJR79A/oNscHDKmS5Ltc00PSurkENnFcpiFqsoV2UJfdkA48B2Xoq6mO0+c
Gnj2jPu/5mTXgf6zNe5PGELJbP8DQBuNXvjcGcQ2EEBz9TV2+dO5O77hzWBWq6VY
EW1AhtPdQllvnLE3TGpexKVdP0VzUyi3INZq+88h1lUMmc1pwFF6+zUXJtPGtlwj
D+583AIzyfx1f8oWxxatEpgXcQjbgnzWVWMXqoI1A0DBnxJhYsVcqt4zXTfY4M58
fbEgdfmauxaKWvr/H0kcXLqVmklA/74DJf/qNSjcU3+CO7tJdwQW7aHmQ58F4F83
MSqZTXpiTyb+Yln658Hc/7MkTEDyTpoLmexcN05cGu7by9KaoglbyDwg6jTZTyng
CWiYPvGfSZp7gllm9sXHhxSEBQ75j4guNDi4/cYnW1uOtBnb2I/kJTpEPNJxE55d
VfCE/ultebiW+mUIHxoY1f8HogemdO7Eo74FKCQLInrSVGJQUM1zIwgt/mbRYDpJ
4SfYkmDULjjcsaUFoDCv1YwWiGEzozOp2wHzqgadLho2ec7toHhSZbHtfmOertlv
qURVkl4sfDGRqrZiz93fHfjOx3P3ndLQJF3rztCZBpNSt0gQk7zJlUWizUdIFMOy
6Xt87+hC8739tPc9RJIX6ZvnBJ0bpEVEgmDUforO3qOaZDjdHKpWgrcfMuIlZjKo
dU93K9n/Du7j0iUrzJL2ykISL+QWv7+Zrtta1csDaBO2t0BPJrkhxFKEzGrn/Goq
yQXo5NpS7blm0nqdjPX03hvemxxlJ9crLhD5jhb6aAJA99kWU1AVy8BJRGp2HhBZ
CoNl7QZLbNNjgVLovcvbhn/xxU3D6ACn7hoBVif6QAKz6TnwilelP9DjMG4Fiu1A
hSTQkwQLnbcjwB/3A9ZudccX/hnUmqMusUacQVI/ykm66UXdPqDTk1eAJ34t//ZZ
yl79pKMNolPsrkNSHpt1kea63WdMThkx+brMJthhHJRft76TRVyiZjKopS5ZrDhp
NF6U1bApiHNGHXXhFSL0xaxvMgmrQiB5YaGieRQAeARVRGvP5hMPq50D478MsAU2
QLtHLR6vmhxd/uAEdONrZ8AFiEydQQVnJ2adZ4KnYTKQx1URZmHr9Ge6m3MHW3eP
RMqc3Wo3WJeerxqpobzM2H3ta19L9nwfzTipcIiisB7R2JPk9H8Gtoeimvoijh7A
c5ip0BDJJgqGt2RnK8V7vjfY8V/Lm2+VT6cg4xxpdOc2w1y+bdNi9fLlEY8RCoLL
bOsSkIupn38B0QPWirWHA5vRDR5mw+plhllVT65KQW35Ypq/yh5gy7dOST+eA2aG
574UZYdGtBnkV2XZ8mN94mgbNGLpjCNGgmCMaPQqXTT/q83VUmystW0Sx7kjTzP0
9z0sLi0SF7RsCUr/am32RKh9CqIG59/8uskzdZAaBtEiKxXyWgPLmvDZcz5ef4eH
Z/bc5PpHgn4UwWBFgEQ8V7Pld7ha0mo1s5zoQwaO3bgZ3WBBfbvNx0zYX7kAP0qe
ZnFe8IpeD98F67hmXeit/s7o0Kggr7eFi6Z3xDEjZJEKDRrMmq8k4gvWZSBw6Afi
lopv0phyucDlV0a8c+kqw184vuLvS8qIZceoFNe1f0yMDUzzpyXg7ri6UHKdUchx
zTr34lfoY5G97DOvZj4jusljwgTkRPFeS/yS2EhMPGIacAMS0P9phFSNT5mICQoH
FXWtSB5VTT0D1BV92NAwjUYjtix0prY6jiOatUg+/88I8kB7i+xbMlX/KrFI0lI9
T4t9RIhRUMG62Vj5jk6SevsyUnB/ca+l/has0fDQGMt77GHjCEO/BNwZ8UMo+7MN
ZtCAfO0boh0+RejkV+h9dfYD1w+noST4z6CFOco4I8rNzao7027Bi0ruVC1aDPkt
Ws+233n1IllRXwAvrF0eeKKTtb7mMblSvX3fdKDWqBpt8I4J7VKd70MWLn/KvDoF
j1tKWuRrlOUVXsa6cxsQoa/sIZlv2cIDCh54E7NbMyrBwfaj4pqoKIsm3/6PbEHC
cJRrcxgRBG+f5wHn1gJVeZTb2lXDjoF2DCf3SmeiwGgtxSqrn0uRl65GoBrqAUtD
hX2RiJfsi01F5FUGuMqfNYMEL0ZEO3iR4nAcSFIFwRjjbqRU/Ct/EHfn8XylKkG+
hJV7D83FcgB+r2ztXOG6CPZ78joNhnNRjvcUtXybaeFplv/12LG7wslsawHmo97f
BgKkemGVrHkLdSuQfLXhsbyFpyT8qTXEEEaq0OpO1zbwrksu/nEVvAMVNW7Idveq
UjoRIr2vOkv+xjX2mcbNjKdDWew1usBbf4F1DTHyB+LMkmV6W7vMoSTuVCPU6uRJ
JPJCBLGk1/bOBJ6Oua9ejuoH0FTEurcCxYRkIkxHE0trHqPJ42S5nzV1CX4BrMUD
q1XUzn/BV9vnKl/zuGv1gRsyrwy4jZXmmkF8AJVqpD1B+UkJNewzQbR3ZKQYXUBY
7J+iNWPrc6FR5m+aH5flaTGIZ8Z7UgCfeKfTgbmM8WlbtO7Cp44xoe7kzIMtt9Gc
6ufCplyjBMTzzfpz1KfzQnEoZzn6MfJMlWfaCdcMhZFzitJOMuABI3uUyz8mNjDR
qG7XPNv0VCJGBZYMSG7w5R0oJm3dEwmYWJDbV9U4LZy8L+A0VPM60G7MpzJWAJIG
vo9o8qCDolXrehc7l4YBVQ78L8wMb55JzjNOIOhoY4W9iyIqpJKhq1i+HHHripzH
tmSTs5QkURp1z8MIQ17RmI3WPn3QpRkzPpS6MblDic4RO11KUSX0IeE+fwTfePv+
snIz88a6adiXEOOW7UA6VyHiek7+Qx2kEtbbojSMTwKtL9xToJgZUuC/CPFIp5WM
z+DkDrzD3W5LT+knos7FXAdDwpTrNYHXnDwIatR7E5PhV6vjp02CiFcKJvVu4Uxu
uqDB3APyVzusfr2H2TgXW+AZBKtyEYc4FkoMlHcsvlDM00LvLvCPfazj/dTv5P8u
cLiEKFPwlSzwPRPYkjTPHiFKRMkkBV/xiDhEw5LYoZkU5Pck7+pSvxMklBPi34y2
M1c0rk06lG6xtv6tIoMiYyk9PfwzWuNmfQUcK5+7sFRu+J1bUQuRw5OVfwQDss1R
VojajEe30F2zxBoK27SrJP0oXG4mUXxk6kzZRzGxcb6NGTPehJFr/47Na8XXbEDO
XLRXx+sVZttOJpu8JvIPpHFgjQGfiSlWpFVL2KCzf8iQR9b116oeJVKvPbaA89tc
zX5IxtgVjr4NllyMtXTD++0/79hXoHf/70hln7V7RUtDHbaOw9vmOmmOJHy3o+ST
G7kDJ/qTWIr60k78xLnhkd2LD4Glb/CBzelCmUFbhAvEzd0lKdpTXvnQGRGU4JOz
ejaChKFHRhK172SHHPfjyhVRqSxbhbBVzIFT+hjk8FDevegOFAF7GRp4JDkUvVMX
ixPw0rZIZ/s8Y9QeY6ZZfac+5AkzUJ3VXaDsSHf+3+/M5HQJAmshKOZ7cWnRQztD
yfKk3LxZdiw+MJonJCgBv6zyElJDh+AsExO1+g11zzt3Tl4pelPPkfuXHxSXZ1lo
4rqrdnFRz+i2pP6DhanzXpxSTIqnv5kRdQ9XS28Mf7zjPHrdB7b6ulYLeYstL0dt
ZflIlc94H4f5hLPqQ459k73BfbwkEv1vTQWJMoETMZJG3ZG9/TIfG0oIdrOBa5RI
SXe0v7hPAlWhkzqqUDtjRyCllFwXHiKEDaLQLikw9kXGjdM9qqfvNX0VuHm0met9
1UTc0lFXnFLkQUPwg+I3GJkXDAC1rhqQD+lVjXQw6JwLXJ07OPSTdUBAWBSXpzEW
ZWhiN64Wg/RXt9c6JR7DXYs7xByv/UAoMH+i7VdrYCV5xcU6C4wDVy5gC3sk8mSh
fAfi/6kh+qS4FPYz85KKfUpbzhck/Fku2j0ZRGNFM3mPUe3jCqtLNLPlcJqo/D0z
2hUSp/NDygObKilTQri4m7YK3uFxPj0oATyLMyImRIXwYzfCJeWcO8r1tAe8u1pJ
Ob0bhAWapxjdAb28Fqyya/2hcLDvG+VAr1JvXOMMPQ2ZMgMgriLBAGMbrNisyprn
Iuxkk/dJ0pOjD5UnK07rNrLTzSsPa30uW/AXKBRO/BqmtHDlqKMYmtJ5L8SPGwBY
Rikz9miVa5aJ0oRBbrEnynRIsC/ZNPXFRaFvNQbx0nO/UfbyoEeA4+YFii37+GdI
G9DBkJ9PMFkftUz1Wt+lmKfqWICMRsTUKolFumnNZixMttOgcqu2PfogzfBskPty
JRqjo/r8QNjZK7leRRVRFNBSUbBEvY8WSGzvCrtOpTosugJqt9W4UiFugPm7YZm2
Jr3JURMxGDczsN1jGJ42i5x67hex44u6stEj2xBX9HT2i4I+UMl8MxNKgJK+YQQU
a7ROz38NS6CJzJl8D3S7i1tyvrX84BXV7kaGRut23IPEalz7y2DftItZwYx6+tJk
nyMxjjjG2Xvfc+t09I8oXCZeJxBHovM6LF9nABbtln5pmaxv75J3YQvK9Z4nlAmF
E70zjEHcFrlp7lEX6cgkmnRfxfhEaZ3WM+QpH9U7XiwUElMVKlqaURTJiMHgviIN
6zo/19YQEq9oZLh0/tz0CJW739Xlnu0GoPJH0sVQPN1pNHabE4o7IVQKgN9HQTYr
2BLr0bJt/Z8DiOda7G451VSo2fkjHScf1v0nhWca3TD6cZn3qBy5YbODOOZQDOQK
10cpJ+BqfHylXGz9fo9JOY0XfUoehn2ub0t7+HLzhbkIFcrOcf339ibEudEJXMDS
meH8CdLwJsY92Cc2bbgW65RhB7HAZWY127bBRCK76tbZFNQ9BtOLcIphrP8+rZsc
W/bqGQ0dyKFgqP61uis4OBuwUDfdISXseKuIUuJ9OdlTmUvspQLo1EW10gYK6+MB
zAS9/PibDEPBiDZqQBTJHY1DAJn/Li2IBvaUA97kIrYoLSFu9EqRc5+DrVqa2Huw
f2eh3j40/78fYpeiMYV/La79SVO3ZBCepx32zPoHpD1SB3dtdDxrgdE6R1bZnZy1
QbeD2Uw1ZM8JhcCVNOgH33luQ64X03wk1HcsJrJPhin+hHQqYr98RdLywAG45aRF
vO4OwXAhGJtuV0YWT+iMORkcY/qkVCQNHW0QhIoT8pYoT0SkRJ2Fjr9UQgegtZUw
fW0PqRcdkNxxspzKhNgWw6lwTsbrPvQ6userXSvqt3LvYGjqiLS57e5RpZb1KyUS
ER0PZ0+GFXAFVOAdC+Fh6FHHCq/e5j0hcoQJOfAWXyoNdDcw59c6KlQyIdPyKitj
dDJTX0O21anBzIsZorxuqH2cEwBnGwTFhQ27WbBRfIeGhHY51Rzya+sDMGtaN5Si
E7IE8V0NwyFJnKKksiL1KoYSBDZH6/O4jYUse2ROVPuM+y8bLLvVbC4AGIhQeQt+
frB1quuBSfN4LHzHjFIJl9vVwNQKHOZpsqqPMLHhOi0bTvh6f/BuBh1NxelqlVS5
Ldfs3wcpl/qyx3kWRZaZOwuljpSdhptOkFxthI+iG8iWhQqpQRXMfnop2kqnclMn
moebjtCnlNM4bV9RIc8NWMy4U2z5iVQZfifg6pp8NtIUoLnFyXje2Z3xWMS1eWXp
olAPIlzSBccp8rD7NS7RjIWNGqKNaLHMeJCpxXmFv2HvzfIOrTkcbKT2az9MXKNO
J5WTHEWuifH9FRPZZFPITWCI/8N+uhK53uXnJPDgBEMfeiBJz3GKKYeQjSBudkwS
Xpbs0QMetXOHlMRRW25A/t39m4kW05JwCV9MrxaFDAfN3gD0yaZ+ZgAhZsF9PItp
LCnWNk7lAVuuuPjuYV5c/Ym4eqNovYR0G852Jy/T+8YkLTyr/lHwbx4hl6SAjamz
G5dkMdFTRfhOT//cC7/nCWXA5PYz8KVxz/NCtn1bhynyHL10TgANscBok/7QLHet
PHZsKf1HnltR+lP1H0Qt/XMAHDgJC+ypnN+rjA2iMDaBlU089fgh6ml8Iispt3HP
wZFnjNcApiZOEBohSmkzHc5IONVqHVZc9eUg0pea1G4junHoBKea+FImePUjIpS/
bVzS46Vw11q9MFLyOfzC+uvceqW/eOEI/ToY0K8xZZFpcRA4m2vO5h4B6vUeQRuR
9+xyOSLecHrDpcQHKtAKg8vhdzIR7Y7NbBW8AdzahjmcacCweY7ohsyvX3fOqSUE
0IHepxGN7N/k/wpCxUgBrUavXQks/zEuuqpqbL5uPFnEtJhgHHwI6TiOqLSm8S2t
MxmPpVyeNf8u5ja2XXTB5MSLLaE6iYC7KSxwUTS65+U4YkSYk+xxYpMxv3DvzM7c
41df3O/CNOshUjlQRvcLHEGBnAsg/VRAWtZmkGIKkXrVcCBGrawsBzCUBBFWueP6
Y9Ru2ABOSzvxIYUieN3FWmNYmtg08/WrZpRNlwVxaSQgF5JyDhVjtzgTz299kNVe
K0feLm+iN38fjfQqQYL6awYxL8D+snOE5EfSQylUtUmX0eCCitDu6jTO/4iujTJJ
QDuoJlFiscY8KLxDTutjmseh5LoipBi46F4/7qqbalLBMbi3N3Ib0dwbzTc0/abX
GLIOlNMwBdu6rBZtxhcdDqOMoZi4U8ovfF8siFAiQf3hFwnNF9UyoUwZXsFz4Gdh
T7st/3Q06Bw34xJlAmOrkMViiL2dC6kFoRnU00Wl8uygpx9xvJRPkdw6gnaCSRmJ
HCg6ge5lNIk8furB4N710beWda7/oe6Mqyre/ufem1QVE+DjB5JhA6qIJ0Y08NUp
6bt6mgyPldLi212c62xsjKJXAYTgPRx9KFuKjp9j7kp0EZUQ6WfwgGo+DsrVZHfC
1P76f0HXSamJB8RXjOwUrDAVh7lPuaCVkvF9ngzzQPX05VkqQZwyPd18c+eU0Xcd
9QVdrn7Ngp72fpaErB2Zm04j83viakkX7zVxzwbFnC1HY6OxRAGggKFe5bQlRdrk
gQZ6noBqYZAdzi5TJfbXvhURxsVYYVzgKfDDybjJ6v+bXBs6x2VjTsTuDFBE1P3G
z36IY4CnNx3rd/GWe6/7khwuzncJ9u5k3jnIJZQs5H6Pmdr0WmZiOXjkkuHlLaD5
jcwvckjnv95urjp2Bf5u0LJp66AGngOZe0EvHX1CbECUyFmcmcnNAPWt1YOJFdjy
pkF4qPCVDU4cN0CZc6x1sRMEjQ268Lys6owaIsaRGu0XwIYhy3dIDLlw1ZI3gjBv
/DfnKX30JCl1g1zuIfrNAl+W724XijkXxGLUtcwtlnqE2/uwtccuc82teoMd9+pX
uxZdIIoZwYfECpFvmCgX+wGppxne0rsb4m/HugNIh7JcGPoa8E1Il94mhDfpQLo/
1kSMhcV/M78uy0L67uU3rA5FRD2J0nVGaFa8EaQqSv2pLQW8N/XWU2ckkq9D5oBI
NWC60ffsxC4otISfOW+j7Y9r0+PcWlJOmeuNOGc4c7IgN/+XKz5tMpQXwlADT/H2
PAkiipt9rEjwsGRU60bntnyF35EojTBzJSanttdUERWFY2aNlCsh26iNnZc+faqf
pOZXKkouUaAjVy8fA2LHhixB1oEE345GpI6C/s/ddxXKaznayR2fp0UKMmRPVoJG
sKgXr78dzBnJlxUa7y6fY7CN19Ej8wDIsMxYEQUjk75ftm3vtRQ1RYx7LqQAtTIm
+1b/jiMszzxp+dOuCYzpVVlx3X80qRXn2TGGHqgR4oo8zsoWzbwXG/1uanjdtK/F
/A93YRFj4SKoJ4sUprNWzE6T3smfag5nu8b2oZqalSdmURI+tGQ13JIJWkb6AKRP
gmchzGIGmaRILl31YYbHf4l7BImGiM0I3H5w/9QMcY8VJFtkY/N2rBt5aW5GZ4tb
xxAiFR054S0PBrLAosgxOUJH2QvnwWNy6E8ftKMpzdLo50ut/+e7KT32OlxoP986
2nyazF4v15R/EjEhqmTFMzUE1PXBiR6B6EfKkb1UXSJHwbxyfWH98Qi6FESG0f4i
szF9Ie2DOD3X61po0WeK1e0IJhysfOQV8xZKcLG4R1Blu55PEusx69xvJgSbfgIM
Tr+7e6i41gKug4JPEIqYeqiLGgJglPss6QuXiwAHQyNV8KY63OA7vD8XGOB3dNoR
XLQwI1q+C53COoW+52aLPDyErbSMwcckznTpzHZSra1iX7D3sYQJV1kZjL+yB6Ja
yyxdrWgHIoOZKwjOqB1KiNTSGOAET7F9i+W1GNx7u4hlaEGNswAY1azO5ELhq2ei
nrpIDKqCaKKJEzAHqNsV8/+TEdHN40fsZ6rAjINbz3Rt9qgM/fXVBDxiLCfdyUpN
HsfHjLYAFFhgbWen+xyUN0HTHC2MWgea0FK1fgBMTBlfOXmpE6akkzqWjsjgZwWX
wIt0qRhrej0ahnhkgESMCCyroUTUTrqMUGHI0pUGB9ETeqPIFPFsdrRwMoPr8MVP
w7lhlfjj1zI8buJhLEVhtM8FxvVValeBremLu1yl3NBsGnD5b3RASoP/oRbgYkeq
ZKoxALhWsk0I4CXdceAKfWyGKUHXZfmG4FlC3sS0RmmvlxecWl42Klk6K2msGRPC
LMxoiP6e8Qe/BCnofuRjhuTfT1K04WuKb3T/BkU5Gxodiw//NQoN6JRAbEhGs5Tl
Lv6LIs8aoKmaReKfvKTkW55dWTzR/+RpIvsn9IpLKV7kxkXkHAoJh2KXe3UD/Ldy
ar7scb4FZOKYNMxAlUmn3Fdt/OQrqGuMZwC5EfC0js8TE+ENAfdPIyswqgTw1U94
c8GnnRdnHYHq5rXyAcPkwza3u+yjHS3/R24InMcmDhQcWqid+Wbvl7uFGYQAAnNa
MDtEFSeluBbTIxOLQ1cmCTUUoFR9lPobYsQNddyeV5gOHO0fdEISy1wTV3pmUDdK
God+n34pcsLjL+jF12Wz97c0ZyeL9T/yRWeU3cOjACfMn5mNXwsba74TMP1o5RgS
RTfS0gBN4J8pbLdD/fSmibskj21lR9hi7yW25CFBmkBP4HzZOLVMHiSm0l1lkHnQ
cBdZD9N6krG6a2SWjCKUlwxdlTZXI3ye4wJr2z7Kkx0niM4iBcTEt3F5M0NR1APX
j08V4PJ2SUQqEuRCOizMaPN3+rAzxEJ1+8WHKajl7QxSjuHnVTUaJTtskpRXNB/4
pkMuw9Gpg4DEGpiCQaEztJ8kRS1rMAvzsRYcU9oEmRJURYQCd303g4/IssEyeSKq
DPF97uHeIH1ZzBb38x4eJ01bVWulG0z0FaJalJ05Cly2njsSBPOWQuFsbfTIcZu/
9TXhzaUkfKStrUFctDXej5txhSVNghAmTcMpr61BNeNJmI5YHf9X/tJfC34CR95I
zd8XU+WXyhjfYxFjkIvxZC3MZA+Jb0VIpUAcmg693hsn2ziQD/v+9o4gY6oSVRb2
2obtaJOiftEmq4UF6jiiL5KQGluKaAhShNlOsG/yRqBXc0LBy7UZ6TT5xbuXs2fR
ZLGKjCk34nc0qRjHV9kRFxyMn+fgBE0uIhIzHj78MhH0hYAvTUcr6ctSacBoQKzr
PqmQGLgJVb2rMw53jOhc8+rEa8/gcdzQq9GNA3cgAGT/JQEj3T6/o4Faml8lA6bi
BadtjDAb0Iy3VqRsvWs1OG7RiLInSgJtLpOcHaiwb4eDiDx0XpkYrBYB1R201e9X
TqHObHfSB9+FD4lXVqXO0wFYO6nX4fem4cSaaA9PtGAqcrj2sKACej3wE0kPnMYn
Ums0GLR3FGnCCF3sWHmS9/hLcK5PvJ9dbx4aUF9qRRnVEfkf5o6pEOi6JbWOArPg
lbDZOYt3JP2FrCrQZr0LXEjshCPC6X8bq7RAwR3/JZfnEbfiVKZvauZc/wGJI1VJ
yYxRvXJDFemqhwZE8XtiEvy9N1nLoheJIhpHnqi3iWwyVdbgF931EFevwbJK9a0j
sBsMplmITWHMLd2CnhzxHxYDyF+2QmjGCidmBR+e7tywhkw1ThFSnMYrqD7sMXJN
o0Ncf5iKf3gF4vYGrCB0qCp1xfo0NWRuy1DfnYVBjiCeeCDzOdX8xR6J8DanmuRI
rV8T3/rUu8OcwMeiILUE1fBLyJF+IMrxJsQ/lYnZTmVokV6rZ/ywkWPuSVXkthGY
7yNs7cXuxEwcj3/p97suVYxGWupdmaRsXRaFIFlp9bPaseNb6FyIancag61D2/p6
TJxsDVHvdUNwPCrpjfuvLQtiyBB2I7U5gfc27iMCiONjp3Xc1qTy9j1YP3v9AVtn
k4UsziZvJHk5wuwB0op8zFJyxvyONYPXnX31CkTF9vqJ5ABmMg1uTibsn6a+U50x
ribCmKECls12RmAbF06Ud0a3nRPOCCRF5mAABysR24evGvOodD3lRgNp/wWrP7yC
RtCwFXAU01vikkjgb8FJMDwkJgHliHina5UZKuwHVuB3aDtFNQLcuEvaJHocrsrE
eQBpkOAacV3sQEWgCMGrcsF8BxHzNic3mE0VPbVvU7XDHFdlJ5FBq736ptKjSD15
jlXR9oiAbz8co3NIFv5s/Eg8iub+Cs7icB+Oxadqwg1z3grBx5XjQHNhWjfKCxul
dDZ0/Pvo+B4A3+M7RfkFHVN0zO+MiwQR9qyZjooCa8pMFFmfyQL+xns5JZkKj/YK
kYrPSVz0/ZDCyTIGepgDhHeuqyyi7ngKYd92OmHcvG7HrZkG/2FaEfzUiQg/P+EH
EBgdrSugC65yBHFyoMsGnDqM3ZAmPWiNgRGmhme0xVBXbgEvI14Ij4ROdJ1J6mdO
Gpfy+ezsl0Z88pc7Hv5vp7/jm7si35t85zQmfZVju/+AaPqnBeJYwtpiV5mtalj1
fe4BgUw/3aPsn54EseIdC5Dq+YVwf2uAmhGc5AS9bAF63655T+RR6HKa0P/IDUZ0
Nrz7Rsbqdi0waD0EIMJbdiP4SI+Ee7kDyogc5UJHPe6gw71T3nNgmL+ZLC8MqyvW
G/v/RIR3ZaQXkPSC4LDcb1lRcj4EkOIcNr53HKn+o8DwIrRf5pcYCw9K4dQThfnU
iI9wjWgltzEuvJaHkcBaDeyCj2/Ub0/Sr9rgeeLmzZKB1E9sO4DFXxzrFTfqFxnr
Sk9uASDX/cMfTB1U7m0EPHhsWI5Mo9Ky3UBP7uj6I1n0GQWpbTk5GYGamwTIVubA
4Jqe1M7mS0gG7+QsTGIHbBpo1jdNzkH42zs7p7YHE2EHEDIhEaqOGUICkqb/Ho/I
/EFv5QhwIuBonYIXWMvlDleMO6ihX5utRC9tT9AVEhCmvDDzkA8lwbQMr9bsRB9C
NTvsvu0rUU2yMQ3UMNUpEtYJILAaRv2mBjUmv/BVa3BUYty75U6N5XB/Qtb3MWql
wg+Uvvs4+TNcYItx9Hj/ceV75Yvfa9cAmjlMMqAGFKZJJZp4Xy2F3UniP5dfKS6v
PupnQtDUaBZW/KNSi5ixyP3Gd8QxXxIa0Z1O15UUxF0duQwEQZISsaaWDJhNx7O9
lutjZrpUqAbb1xcKt0ZyacvnlT6aadLL3LRzwlPdzM3T3Ue8UXsIuZB8VX71MTWB
VDMsUGVkDBnnVbxh6RSzK+KmkYi/XyjJWmdKW6B7gjUiPkSoTIk0VLneX2X2fraQ
m5NVGQTiK+qOW/86VHtRTUuSfkUAVX94/9zfT5NCcrrppdwPaY9QRQOpMfDX+/bi
y7QgfmnUyNAgsyYRkrzpgEbHRZ/dnqS6svoiMM0p5MOCtHt/djfcgZ2dkFO/tzad
IcGcicDAVY/cYg8SZF5llq5silXaitXpe56/OEHofnou0XZIjwWT+XotZhRy4Gja
UccWEIrviSeJCjAmL3MwcLFL0z/WswD0DxowBuRTUvSJivz8cs5PL/wW8aFDfu5v
NPwe4tafceuaR/pWuwOjU1s9WCaKWZQZJIQcorakYOZMqR49daUSKQJjXbpqCyru
CStLvIhyqnBDH3PHc4ECoW6IlO+Ec0H/8X/1o8CzPwJAzL8/EKm4fwxRowFRS7B2
EqJ8lKRQ20C5ushUeVjWStrjugHqTCQIiC9uOqT2hVtcfcMHJZRKasPCzWZTdRV8
mOAzLI+TMnIFp9x/t7mzCOvBo1dYl5tHvO5sWjX2NamsMRvUcrZLQghiahXt0gXI
PGaBpRmJcztVSrE5xP3axLQToeDEfAKhLgeY0K6lwzZ3WNykhizl84n/UMk/TMmn
jXUgi6pPiYTSenyTUtN9KXwNlF51S76gHEtxtVAaKxO8EJOzwvCmz1vdybn7rtUs
JSRcd1ANlQZfHnbDMAsg/JBh37IOK9R/p+R53kEGw5cBYvoiOIAKh8E+d5ilefZA
phrs6To9S6VhfdkaQKmT7gAM3PdjMS+ZlkYWMlGeBrtrKh6j4ZcG4OFfiwBngIpJ
Ld1/bGMsisM+G+dkCrwllqDP7M/L1jkXzsVl+nTnsFJ92J6gaqc18XhYWR9SlH0O
FIikqrc6d4mX6AIeEMxUhHb/zFKeO1W6QU379U7XvnQ7E07yb6wexmrRxbwgi4Qq
ALjPJKGrGPuT7bOFTEE/mH+DC1Y0jUHV7d4dughm9trs5SS4nUTOIE3uvsDK2BBq
WiqmYoiR62WjEj1QGcspgS7DAkJfD8eU2QeZyWZnTywCOZlSEeASGNcHEH23iT1D
y0iaV3WGkulKdLOW6XgD8QTHeHjeVbBf01C6b7USYjM33evktLXw+/vildqgmr5A
zMz+HejNOox6Gij8wI5oFHM7zBop6jnH8hSxtggwLW0Toe6d7UL5rWQPOx18w8J5
e4H77j/+3oIn8A+KxwQOnQaAQv9YERnl/vHjzKgPJ88iy4lnjd4hMS5o9m75oF8s
8YV+ysypILqWCmzXHnNChLrwT8kAfeDu5W7pkJvamuAngh9KaGwaruyfdl4940c1
OfmPc9ChDrOg/mXvqwAKB7dI/zOFwyF+qCIvHEQgTpfuhsvriBkI+izifeGSCAdZ
DcB6EuP0r8a/J/PDhuHpJlpfPSfP3HBIYC3lEoUnADBb9ixycvgK7jvuQXjW2OdM
MsNlCfuD0hbp05K+MQd9cmV0p0ZMg8dttH56M0EY4eSSY4nK1kImPlkfUDrojAL0
A4lV6JwS4zXpNUEl6Lwy4QQzEmKHrvzftqh/8Hr0OC76glRy5Zl8SSM0sfghh9mC
J8P8QI89mLosk0U3hW1Pf3kknxzH1i6aQBsUOhv/gs0hCnDtJvvofUN9z56f412L
2bT31tD4m0HaX2bBqJNBuxgGHKuFg66VTxbI3nm5Gt/BcdF09j2EP5kjhXIJzM6L
CVpkBh2ZacGWXapD0qcONZ5tIvRZPbK/PXWpK4jWK/vFWTespRPaKwweBUwJdwF6
ryMM123hlFyX7C6lcRbnpTrUXtf7K+hkBpnYn4HCB5uF1/IgRSW9kopKde2EIUab
kQMwTnGjSPhQw6hRiTEDDuaMtmNyssQ/VbXZIugzJoyUrhrBaQxjwVe4Rwke8h6S
t5ZsmWrBt5pOyibBZjv3s70kUhaEvxA4M106yQGzehDCV0GJvY4j0f7h/hb5HkWp
RIOWnqRH9R8GqMee/PfFKsn3Iy704w9FVT5uNoNfvWkaquShoOcVlFS5WK5xuH68
I+F8Qw/Yxu6EaWbtwVVfd/flCdWGJLpgHxMKT4wN0makeYwwHZIOi5W0ED02bBHQ
4AP6m4CHXl9AsQ8EIzn30FfRzqH/ePG2jazM8zEBzF5lLWMaTrZ/WkW1j74huxVh
WnnmV4AIS91jcQdHuyrovhvNWFvi1Ie1EtsJE8LjgdVy+dgxmC8kNsKz1eKXe/K4
1FxHezaO9PhaXTbqt6UKgdQlXobExCubIIcnDKUNoVM4HrJjxWJh1QNRgPlIe9bF
OeDZVY44RMMYcy2xQ8yt5bKPEj3uNCn3fJASWPlOpL+Wu7IroDmFyyc86yRQ8hAF
G23VzMyp04XiPvj1kXQYSDC0i4ttd7j0cGrRTRLc16ZxIvp6i5jdk/wmdshasHET
VMenYV+TyXuIEqOd8rrt/KhIImlKIRklK/N1SW9ZpME9dmnz3xUTnjq/1oiVSbA+
wQ2C3sqPmYWzQott2QONo/CsUIwbIMVbK/YPcNAhyVmCEA0q/JuUVhx4MraxD0gF
OM8nntcLWXZ6YrVtznlGZO5uMbJjRA7DamucmMHkU3ne+e+kUGwCSg9920AHulaQ
lv3rJ0+bZI0SPTRqLzNJgW70iAySp6R7hQqrMsDZ1lukeXsF2Sz2BkSDuqFMv0cl
H8ygqVn0ooXxRLIoG2U4l/vHZ4goOKnhk+f4zY/qRFI5aWgGoQCHqWvGy2c8QmYe
U0QXNspG5ShfIrsL3bmys4hyaYFNCx6zw5MIdr18+6h04OqF4nEAi6Lov+/scjeU
L7LUBdR/g0WU22r03AIqNBFKPspvXp2ztdCImByP9A+OpmJ1k6EeuSAmmhhwt3oL
itx7oGzWgKBT8VzwYpwCKij2e5Yo43rXN762fhsw1DoemFRVTibytHsRKxErplSi
LVn/19wX/OMjgg/eOpmdoyBqQNszvbsI0FR3Dhe0EwNUmCFvZu9CCk+H4SB9XIJe
QAm2A1J62kcLmQC8ov+tfM/Hqe72wulbhQkQXVItfu5YuJMtwfPvaVyNtj6THQqS
HRz2mweheGu8MGrYN04fHm0706MPRssa1PZcRk+nvB1gyWzYndzvJreCC4TwEzdF
jqM3oS/pKTZriojNTOhFhw2fUBUMhJirsrqzoWw7OfapASsDlFseHvR70qDKb6MG
EMe+YS9iz5fKO+11XMlIFb5aB+9C8TjcUieOBM/jXTu1vsvFvHl2ruZzRH5H8hQ3
fUqce7SWMdQY6WeUQg98GgPbX40Aoh6/dhhj+z+9MLktlZhZhFnZBRWne8Ksd7Xk
tG+kJnrKigsRFHFL9lTYSlb8mAb8NlBx/Sgq86lcYqew+3ZAdj5MOubZw5IxNge2
rrywMCzrS39o7p7LmmUszh0PxoTXT684gI3xfH8KX1rG54CglB9hNy1SM9CgmfaP
c0+pnOUZXWvn3MnfC0wmiqdVkukS/mORd9XAUyb2tFUUDKCo51DbJ0rtQMUegdNZ
kzh8JMi7jMsPmxQ2/EhXYPp8j6csBs8FyIQU1r15hRLMu1Fl+umsZjvlm7NKJsdw
Hk8lOX3bIHAzZ0TOCqFYiRVz9vIhq6CsM39TfgTvKiGM1VuAk4x8Xh/gr9D9WK+i
wIFKxApQHHHnOcXk6JYsPLKEoVtrjYhsLeTI7EcmnbYvJy4etjoqwsvxuVQ5HhuM
VnFfoFOOiG9sjJ4R9ZSThQnTfigC0yZgXyMGKgG06VgbyiOWAERaP0Qr/QXCvwnU
7ZY2ispQSvqftcwxNxq9LDbnxQbdhwIj56iTn6oVAb4CiUCT1jx4iwJO5j3QKJSm
RLN5sburggMx3gZSf3UAgZBSYpY8XMnshPlxUi/LfSFtn3dR6+HtRHW+rXOIIKxH
cQw4GU/R038swrejBHEnXu2oDsTzibsRmf265mI6YL3A6hfNcWFNJhuNn3Ihf7a4
Ea79WFin7+JhuOtaxl6PY5wDKJY0lCc3kVhwqcnUlQSuB0Nbdoivgw9TmII7wzaD
HYTJ97ZUHN8G8nidRlqKJ5nuGG3Pa15a4ABQl35Ld7yNMHlpM9LtblqYPKNXlMdV
Hygj3lnTVVr+kliyxsDeckmyIycWUlPwKmGnBtKJMFlZEuxsdZ48/oYKNZ3BD4v3
/nmQtoa4Oc9R/A9Sv1XsLv/LnechxsMjeScTi74E9GYX+r6ZlN0iEbAlJ6LqAUyB
A4l769BX8sZN7iLVGmUJKue5cK2YsFlrZKgMTBV046b1FVrursz2LLjJEP8scBbZ
tr8B9GeObzrHKkZ+B5PrKeBiVq6Qtczwiu2Aec2XXkqMpjpSjtwoQE4SxWCwqSs3
4Dg/CRZiJxG9JaCbIaRsqtnGMoZjZIda9jQbMjSa6RLB2Erp2d0CbR8sCkEOGkTW
/hnwlHqyhHb/UvC+ocsp2jloDis99mWoXlnBMncEN7pSICQt0VotzRjLA8OzuO4V
yuO5nDzD443WJ/wOJEl14uIFTee9M38PUyGVl623jbo9SGx4vqIKS+ryYEeUgQrJ
53RQZ/f/rczmsOx+krW4458UR5MDX89/+EwG+XoNu0JETDwvMJl644iVQnILkp5k
ZwZGZx8m8F82iRMQLKpOHW6n7ehlx0pVcWTUMbGJ8Aks8XyHYEFBdbqbFBTvfpru
BeQ0onoZIyEaZMX6UuclcKnKkskglPaXLRzoreYWJvLsgOMr+pfgTcWzN969ePJG
X2awcyPznZmftrdQCZB7e8PQXW4EMT0fISzD7MiQN44pVGQU6EBK2R06tZSwvJtn
+F6b6jfKo1syDbE1/n6m3NfSeVvCJCAmOJHAy9uY7e/ZoEdI85yRtd5tVp5KNvKR
GSpXUTe9Yi7f95mik74Be94nOlPX1UJHeYQwg6NJPrAPsl5MNd2OmUCelNdVTf5c
jpY/AT4Ec56aR6qCzuj27zYfE57CLjviSdWTRZTdtSKWdcgDgWxr/kD17IgFXLAV
9m2awYrGfDn6TWuWqyAwgdKcfGzQgGOAxWGVtcCmr13BcL8K5FGptNxRo8ewQ4i/
3b+RmDpQeuqb8c48Qo6WyQK5bnf8nV3zlnh6KwNJwRLzK3CRD3qTwmnBSratdOz7
eZ16KKCDxy+kaDAE3fyoyRTtguEjmW+N7sfSvL4XcbXcgRW8muysDYTY+rZStxxY
eebL1FvxB9ycMo8zaXYedooBFsjrcRxcceJ9+A3t5dl9aIcZrRv6KPtWEuaCtMOP
QwwVWN+mGjfzUNw11Ca4eruqKn15qYlAMvGKc1kj4likoTmyZJYzL5wdndtezQSV
KaTT7RkR4UObs4nTI1zhbleVkuWrfqC2URtGNhNfim6tykSepSDG2KCMQZ7+hyJb
bjlKMaCg27gYmSpH6KlqrV6EaUSTWZKzZFIqqgmyIFUQn7yfo/JbQLX4+3XuZQxe
iQ6ok9tIRT+OkiNNI7SSR1OzRxrcQFulHTW4CkBYWd7tYSLe8o67lnCObXxlzlu3
n2uhVn0eufGTYmlApRAHINCjYoZWxAnYK+I8wq7M/NaPzMpyGpfp2G32bhj1xHUl
fEw+hGlqHcPhY46NbOOhdCn15n5JnWVlDOKqddPR+SbVcLemg8YZ0q+O2ep8z5YG
x7PJtH5wAw7WcboM39GFUJ+0m+5L7TtJz6mJFjpLhv1cUepK3iVsf27OTJXZFAin
SvhECmiDFZFr8UIgh6qyQC0/AnOpaLWgoGOyjB4VL4I/aUXnO5ZNDgzVlmK0irHE
oJzQWLxBGPB4WMvs0HknnrYjIgrFW0udYTj6kwDELHp8IT/kUMjmp2b7/7OXi+cI
CZpjER9qa0AN/VOhTrSuuc4m47nZiXn+Gk6OS5IpqQGQlPxkXBNB4fVuJPEPAzo9
HqdWuUdC4zCr042iijujGWb2GthRJ8nLBqqA8SHHmCg2RFZ+3f6cJBIIKrfOKcMP
cVjPWCN/Fc2gnOgFfTXJOW7VW7U0HTAH6CsGTRGhMwRtYaraqZkmydcT8JaRV9fZ
pOukX5Lf25QldEvRJc490ZW2/WLOP1EP9shqzuJPmEgq01oQ2Q8ic0g5hm3P7ppk
iapnKwg2jq/+vIunVaCa7VULruJml3VfEr3oddULbF/xQ7/kBL+/NGzc1ySKJKTH
+hybbcHvsmAKTWLAXEfU3vGuhlPMnu3XHcjCTgKkwTCb4AHEO/3pQDq9jqZdjHUi
indJXEVqH17WUm6lsZkO+dKFGaQvX72NJNSJAeglbk9BQj00gBH1GGU1nSvKHB2a
9TIkHa+KBYavKQF0yFXeh7RRKa0KNocflgOnsLmsDrpYtn4kW6BmViD0klNQcO7k
sZz6icPNnUsaA+oypySLAZ1W5xZAdiGPVcuH2kWMP1G/jI2bxhKDWzHwKMA/MS8o
snQNuUIF612heuBHWvg0B8rOTae3vqEe/Xa0TU7Ydy6kmk+SB+H5BGnPIV2m1Q3C
VZn4N9ggoG6WH+vwKf6EbbYy2avgVVGTyLcuCKKVY6ibgY8IjC1hi6qhkj4bvpSY
VgA0h2fC6syPBHbIG3tMvQr0ndzdUYH4JoKYhe/pxcQLTxFd3yZOBhfpyg1Xxj6l
xRpEfA4vrCu7Q6GWiU0J/Qt15mKvRO+KmSYxNDatNGoB4OWrI4KGijN8MjxBM/So
GYJMfibDJKh8hj6F5OIeEG2kbd+6eLQA2ZrXa0hW8mFx3zax4Bsw/+D0yp1PzRzC
K6CaKgcm6R8yQx+RS+6aXFvcwZDtpfKwTpzylTpekgXrX6H8Fd/eCwp6CVtvZ/dY
cArIRJI2belT6rWzDJlMuVBR6Q1syzRXGftsdgoiQ9Lpdp5GkPrspQ3ZPliZa1VI
KdNzSAVzhZI1931TlomxhKDJ4P5eo1V5eDimccEqPEnoHp0j4vJA87p2nRjoLC+y
9kqHfsPNPT8ZJofSjIyzE+bs+LI0hbLObj5KMCvN23eR/zL02Hwetuwvy9XTN5/6
H2PSsIXIXMPbumpDJl5Nz8GLy8PvO7ocxlHfUfFRWe+Lxv+iKKr2m9NBNW5yISt2
k1XBkr/8PSBY245TTIYyS9LFl63g3zKotD++8NxKdeQ7JxWIAql1wlcraJxM7sTm
P0EVyyuJpQrQeo7dQXst9yN5Wjp2U8O64R8oogJiYc5TY5kPTnOD6NkP5VLnYYDd
o0y1XhUVom9sYwHSWejfmRl4sOeO1k8LoAEojh2Vzc2ecpsozp4sIHuCMUbpgopo
5ZxW/d2tw+zHeipWziR1KPrdcYbLfFopYie7cfIvOoXl3Zti3F7rDxDEdSf5BnGg
vDXRVcjuN1n4FJBL5iqtc76tJvDG6Z0EWekdQAC6Us+Yh6IzRg4f7Yt4BEH1+kHh
deMBMQzWOek8SWFzJrM5qVPUtJxi9EiPZbX72D88hZBZgfN0T3iWfvSEr5GYowIe
RrYJ8apF+XjG+u8i46IsaQYfjJKng3AxH002BDfLKPVfEERCmIjEqzHrvTmLR7lb
Ez30EThLJdc2rsHqSDE4f2adIilBHMI6YgmwvpHLRx0FL9ZudCIg8U0GjiSy7bo+
bTKkeiJS9OOAkUCDcORvYbaZM/2v8RuoPrrBhjagEiZnLwNVg8uCAn2eGXBb4m/o
uayjUJOX196g4cjg17h0fkVDYTvNulktjO3CPvOG85OJZxb3SQkes7LD82Me/dYS
gh8i0bbJKzxIbaXhdDDbs9jxPDnezYfBWMmKkJbH2FMOy7xnoq5AIeC+Sta1Zzuu
WpswU8EXX+H5pRCkQyGkgUdWNkdgptS0qKUHQfmmkZX1Pennly+42BUWr1g3WVAt
5K9aRscJAr9Toa525YCNS1xEmGLKIjybNIubkx0pSak3NvtUwMVxu5qqivDoy2GD
xbI8OqiTixGyRGptEc1HiNP6Yc6YxZ+RoFkb2y+tivvUH1gkb/Sr+e9EyjJHVg51
vxmr8bGQvzl/HMWGDXvQIBZcOuXoSYSMZxmwCpG7F8O+/rOGffPBrWZzv8rASYdJ
mcRMmDiN5WboTfwN7KcZxQw1B5qWn0gSgHvDMVRhYHmg6hxCl63S24eV61b9Oq0y
ScIAhHJyizGHid/pkx1gzG5vgyS1av3aAT3C4Twed3hUaM286fR9I3d+TupANY3M
tOwfvrdU9Ae6JImKJ3D1xaya8dVVPsqr6WJ695pTSkCsrkFxpZP2/UQV08RgxtH3
AA5AzZeEmL1BesRRCFU9gZMcivU1GJ3lCuMi1QhnmAFFQk3k2RLtI/w9gZUiV9nG
+nYVdyAvPaKXEfOVBO7ymWG3S4C9UN0+dw1NCe4YQIJc2jlqw7Aw95JA6ZFjkRba
JsuUkAiCLyGn4NBWlUzLRZYB0Jg89rKGh875DmK5lFq0ZoDn2bO3DUT7KQvM57Fu
pDsOBJ+32gHURRxLObOPF+NDb+9KqU7Ck9iflyy0hsV7+QYeNAfifa1+5AXoG1zi
7Karcnjz+9wwMSRU1z84qSEVrMsTE25JlAGNjjou1dhYWV/J20yzhwgpjUthjsdP
6rRwXyreGBGZB2yen82+Vhvh4WL9tQUlZY8Bn9ByMkyDoLqXr7nXZdSNHHBaBUhj
G0MlKFxkeLZIS9OFrlpenN56rSkelnqXJ0/8MlLCgFos5sA0Io5WriUMZvO2rNW4
Sbe/6ywlg6A2LbiG6WUeGrgSvRBR8QIFWrs02xCQSjU1d/ZSwDdNq9KvJhp+3c7A
OBLhnLF7/QFGuADixRz7VewxZT2ln7etGNfW+03gFT7AXExpg/BhrDJgN5Mt8AMe
oN/AFP570vHUMxUOjjvZT/CYxB+GQAXx+AmJHcqnDkVyuIPIgbfjYqDz9Cw8qAbu
xcyP0GHLppLe3jhP+nXmG7t1PJOnZS7C53UTxvq8HAbhuP4Alip+0iKM2oGmEMtn
nmuMl+LYcstKN065Vnkce8SdxF+4Y/JcE+6cAP2wjuiAeCGyzQS/w+Wwir1ekhX0
ilfy+9k894wNLJ01BBZOhprCqkmOZxSTJjJFLXSzWT0zgymzI1tOcizpDoXtVzp+
HK/OrIgFN1+qHcw33iserAoKGgvTaFedysBDvB9FNUaHKmzyquYsRwqygRG5J89Z
yO/d7ayUIF/Gx9XvYjdMEK9cYasz6qSaWAZlNuORlAy/isI37rlQUevIC2Vws7g4
heVVlAKmDuC6hdeu0OU+An6ODVVEmppS/SrdcShADPzCduxZrFWZukNlhskKvn/p
qTmC5KBya9Gk40L5MeFa26l5PeRDf/AnMxrMWi341BWqT7489/LLNwAE5+xVt/33
86uFH0ltIQwLqo9hbSUFLvp0wcFzmraVVxe1kpIm9KDYXwhgNR/uvB+w3dzDKzjZ
k/HJgUHO+CQDukpxHQbbFJ93kLWMYLMfRyek7hD8baW7WVKkyUFDMJJT84CRPMtQ
xgZS+/5AGL5H++OIGYayOfx4KX/OSa2Sl/uN15maUk02WmMXLGFpfm5DuzqS0KkO
/HiQhdm1V/iwvch59M0bNpg6ztlvl/J1PEcBO2OEDUbOXRxQcl92uSO44PWPqoIR
GoI/ZTxeSmyUSUKec6a9hif91WHyPUF3DogHiuuLW5eOaLa9VJWv7WGb+5UvhxNS
HHUvc/LaPB0i1ofjXczy+3FJPIy9zDbhyDnomMgLRS1yNyE1FAQhjO+Dt2ltco2U
lYFizOAMeU7x4vN0pGLNYF4EUmzoH3JDUnjpMG8uKeO70OGlDNeTk7PbzjlMbCzV
byyEoWPqW5UpSBPBzadGtlXrNm1E4oaKGnSdktiJNJsp3qJmJpwXSievAa+Q/DJs
ZyGrYEa1v3IgWdvf+3ZVeCg/eUQJq9Z4YCyEe2RSsZq8qAqDhLJ9mB5ty7VaAqBI
oqVPaWNbpMeNcz/sU4NN++9YhFoW/JCqmfhb5E+5ioEJDCENOtzBfKpvrnrXTrsX
GVjRQ/62u1jIRZRva0dVlEiHFVVXsZTVix96Z+WDbBE/oiTszidjPn5q9izvow/u
iES3ccgpIACfx1ptVnOtRbqUnYFjXfJf8lFyQ6sdG4e9xUrIYV5hlVarhq93bkUL
DSJ5lMv4zJ5k2AbYCqsto+/e4pnfSsLwNFXU7OeHtElhpqXrzQ94fFRhXvzKeSxq
kx57vOBZHGQ3SeaYoNQTwB/k17YmL/Pw3HhYXPSZX5t0aHhb0MSofyBa+MIC/C4a
uIcVklzxZPlQZRsXIAJiTRczZr1Zbe5SDuWQMCXhDJ6kQ/w05AmVsTEY039sSWKF
NOXQc6x3GTgUj02/nXk9zyj1jKX0/9auk263rmD7DAz4kbibXEEbePM2sHvkrkd5
e09PQ/YRfcGKbBDYgwwHiI1TFrelOPB0rbByHjpzj+FkZ0dNxuuIs/Lm+efJ69tK
NS0w00e0LkvOqLF5oYNY5cq+f5Hc7vdPR962D+SVfoslStiUanlFOZkn2x2lBxuo
M4YcbZgOnrzRThiAIShD744/yMH7sXtxsp4JDA1A3NQvaQ9yZddruOb/vkn7eWw6
1LC1CrrFt2cNYWezlTuB8+6Lud7qc1Qc7N4vWAppjNbZ8KthlZfCbGbswXtcy1+p
vDZaOpZeOkYaxls4ojPOOxKVg2SG1IfEgF9/a7ZQFryU8KV7YXB0U60G0UFTHNen
lv3u+yeWZtA8OHaU1/YXo6mBSh4/5h4WvKkE5I65TkNZjnhVm/c9kWYZyRNDihnK
JFNRpKNiRbaC8Souyzlbn2hlOL7M4CSW7CyEkmVkRrpUjLYpKoJ6Z5QPZm20bEGy
eC5lC2q3vpnzB3Q09ZHhBMuSA6zzAvuFKU+cBgmtRh/lO10URlUBtQBKIkVTGGkp
+AdhxfikP2QH4eG7rD2NbzOVvpXorBfow/B2IDqscwQGoSPcwi/rUFYZonqc7kEO
yf7/OEISHkLT8CLEuVQSTe+eJ2M40kXMx/AUkdxXKGjdjAOAj1yeKkre4ua05oX2
INkMKOKxzykKbUG6GAaxH8z/fOZABtTJVJ8m23XdB4mlF6TYdbJFqYQBlj2+dO0e
5G78ZXSpHVUwAgwm2NtuO55m58zbrfXvm2qr9hZlIkMMtBx5P4nXCVtlTa/vaMdP
873F90m8ewAptrl0ODKVYFmnjIIVOsZ/YnYyFXCNxSrOCi3f8ilX8BzBNxTdPfl+
BH0Xh3upCippu6gYxi/5+T62IfUH7Xt7zdDfsGlrL3SnHAAbnHBp/16Ftc/9YjXQ
GCZRdmfcuFe4zymVuKtsta/0dMoLln9+wlPonBU7MCBw5HsqQzgauQYy14WNYXRp
YZzCaVETwPZHdn82qtjpZPHDd49cHBAcsTNHBfxl1iH9YwNCgoro7FQFMkx026+z
loKNGsJdT8bzcDgXC0KZE73V6G/tCvWnSc45J3JiwKCc+hKChD7iPkXo3PZqSxt0
mE9LBlI5JxIDQjj7y/XMCpR+sA3FQrGUPGH/f/MbalsFsXarYEeVtmhucIjbdnat
ZfHdA5tTnHy2djOwPHQGFSl0ocdg5P/Sq+BkYqV5Ub/P4ThFJuNT1gmyMqUa5f+w
S16Gc51ys/lXXAKUkmFpnU/xwruMfMMrhVtiY35tHBSiSTFD4bx4Hg6UuZFILWTO
ISX70cYehZPxs3eeWJnBDdABqfWN1xyXo6pFJz93olTSGTtle9ZLme9uGQelEE24
JB8kSaFYZ9jTMDlX2nLe9/cWkLuS/E3GkHn1lPWdG4TbhNzdAnjnnLsOY+l9KcT6
KUZFCq7BWtss09ypp6NGl1XCzvgI+9MlS5CzIyiVtoNmcYNDBUKF61vahW9wJdiU
V/dXRSPt4SitQEgoKomGpMj4k9EpxDzl6hbhNVdRzSUjoM40UQCv08DDTT2Gs2bN
W69ydlgdA2/UYLc1Xu4a1A5mTZebHy9bWb3rDCjOwdaqFW0Qs0nUsFe6dtAZA8ds
8FleX4VBsQfM8dFLz1vR5MKLUo1FOU8K+DmQ+5gHKKJlLryYci4Z3ABk5RHYIqeV
YVDHEb6JzDvP9gWT/nej5yq4rVjaIrD32SYdL8zihOhKOxaZ2jRGAuN1bdKQjw1T
MabpbRl6Ixm3GAtEbbpz8Iv7zrvNDlOE6/FwmtlqMrbCXS1S5sx9IlIKtVsd5IzI
y6GPeOOGtIE4xAiHG0KWgW0AFmdHPVIk9bUzVpPKbKELcRDSkBUg2HCy8XuA6AdM
T6fag/qXPxhJN7ea2Ma0YuwUePVIXMKGYkOJvZH2sOb7YZJPBnUjKA62bo5M1lGX
ND8tk+UdIRCXjlIKwpslGOvZ/mIz6S6HBRxcg+NAoyIc14RbhjFpJkZVrdo8Zhxx
oVuHrdC7pUkPA9dTDbTJDGe01hi/8viDeyBDnpHHxw1uwAx/kltiaRRl6ax+203s
1FU0tSxN39X76MqahfQeKo86kwbTsER3Gx8eMe56eSpQoSk0hAWBcvxxaJDp76jz
W7N6mE79l4YhPEb27ItCTUwMtehrFOCVGcrJDBNtqSSV6abbYHJ1Ydk60ZSHiY3N
qa7a5YnhKEsluTBkDeNI3qvps4QbyCb1Amwhc6evrwyX4zE2apO3SrHPMSGnf7+Z
aOypciLzJdoPzYUpVjBI9YawTFCp7K1ky3Etwjd6JpT4gQeCe/Hn19RpaL6t08Wu
h6tMVrUENa0fO3TGwk0dyUuqLCiyz6UWdYtsF+ufm8FzT3/kPz+ZpLERl44KMF4R
MHlgpGxShMFWZIQ0q8ZWmBzxY8HHMTM3PwNgJgfhjrnfZHdQ38f9DutHuf0YbB5u
k/FTufBxqZTJVkd3Ae1b+GbncQoRBc3Te92mMCSRrhutP58eiuati0q83gdxzaFp
yCuf8j6T8pvz/4wOFjnb5Nau+VCJ2E6wA7fIVO22BGmTDgN2eRM/fBnYiKvWjiRk
07BlWo05ZG70PYjfFlUrS2BnKnwQi9u0Md0CryQEVV12HX+MWfBjHTqaVb9JRLqD
AbnwrqCAXAH/FL7lVhAGXSCnLWKD7kRhCp8A/DFgjW4v+6iOj2XkEOkshhYjb96i
v6EZs5rrUB3vpWCp/Hoga7YV6YuQuRRl4gdSjsOHUtYziK8sE0UDL1FNQb5XzWdF
QheBWYXVK5wM+bWvFTdxwSO54zdDeaB1Tg++SPRkYM5uFxvaXMjwL99hCnqjSrZg
rHEtLqCLbwY7aWex6+CwjgrBdAk83PLxT7S1ZM9CkisXXLEehl1mQlbR/0KanFkU
GIo114c4895prgLJ4IdbUyd8DjyYqbkwytixggMcSZUEK/a/TWmnHDB8M9EZoBNS
16EK+HRaAZrUbWo+MbrhuQrdEBiY3R2/bTABVXWkGMImLgiHufNPhzl3YN410Ef3
UHwZnd9DuE9tVfj39l0/Y7m56dHmIzAHZStOZfbSrxmzcR+dU6hc2PIW851ixv+S
EBG12vtjreeMCxeUxP4+OIbhB0aogqhbeHragJx6dkykf/Mgu8+8TUQx4GGziLTh
zS1bRtA7XyBEvDdAalF1YalKrvSvWfSKLSACaHF3qfBpGhqtZTpJ0fwk1L4LneFZ
Vm7LLIUnhK43Qom6SQ4KtPpVpnXd/VfLX8xSmjhx5pjGwEycMbatMFoL76kRIIUZ
i29daRARJVP+4X6ZofnGW54DNEiqML3WrAUww3EoSGZQISVrlIsk+2GC/0F24TQu
JfJ502bWD7cSpMh9sdoCXRV4rluFnvO01wmD7CJW02ti35Nl2j3N7rezslS3+G9k
OnMKO9BOl3nYC2fbj/bU56FuOf+fsMs+5LT8/4tOZgezUcoTrZkas0FyFchXSKLu
erFAciw3ZlEApkYGWQte42oyNBu+T4UeTjm1f8Om4oWEm0ZZ5NK6N4zY3kmLvi41
aklVTYQ5NVHhsvuwY0ryGhKaT1krKKu+FD/I/1cjA3pMLGjCzdl+oPUwfU3/P5Xg
GmSQNn9qtpC9xAS+sqzyEkkgZQaFp3/JEZoAsMFN6jvKX8oCtcz22KkKLkhXcSt5
wJECT59aD0bjaLWAnMgJh3xFgrYnws6ShtW6URwX8YUFO2rb0tLrf3YZ9QHigsow
aFZEIEcVuKYDy0zhV/PKouvpg0QLK4yhElWEnaHTLSLU/+QFh+Bohn7ru9TBMPKq
WsalYWJw+KIc0Bo9FxEaGFvz/0r2/GBEgdsHxiPlZPLRHeaQZncjPBkE0nCnN1P+
8CB4S5nn5qJkwYvnAbSqxudB2Gm5VPqENWmUHCTbbt0cws2wpV8h6ifqYMnwfXMT
rcXShPNMDMNDp+42u0PP1luTmXNBt19b0aLxcqHMQD3cpdRb7thVrlVhFnkkqueH
42L+Z+MrMuNMSk1Qr20Y35zGXG4PSI4ORsWVlnQkJ90m4XUL0QZd3l9ltcxW57Rw
VrmBnADCipVyImQ3Mhv9UkUhA4Fk9e5AbkQ/R7BQeYhPPX27UQeRSf6u7g2halWM
Vhuc0GgEsf4jTtI6VU//AYeVwbn2wAjiB0ry4UeLvBBvU1J114PoC2TCUBnY2Ix7
QqlAEjdXMqUB8Sf8bko/txmYgvubABcBZPpHh4fB27cf37At2RkaIW7/y0cdXPNQ
pd5geYtVjFGK3mmdMMmfmLRCF4BU623ljdXFOIMQycLXJSAIq94BovrEfNYN2YYi
2lTVvVBDWq5wxdPkQEbwklJLWwxVfHlDyVp8JOCasixlJx9MabTEDQ9xWkskrYlY
Yc/cSl52gZZnxp7geeb3b+zqNg0tZr17d0j5GiYdprwkf9mpH6PCQLOFU2RP+ZeC
W/bkFMIJhJ9maxDgSpXQELvr9O/XarIoYb6FP5/+u+egj1S18D8n+SBDn5Kux25s
KSmrH52oQ5khdjyfU2jlUHzb92+uOMIkAmlWmUo8MtX2VEUdvL5Je0RdZb+2I6n9
TRSy6KgVJqJtPMU+j//sA3kIjDB53ildeM40XMzwZfuMQ4boP7er6JdvFChIInnK
5ddTUt67lJ4SPZ1VQlKqb4z+qg7vicDlisaJvgOdsCfNxcAkW3pGsbxAQrCbre3L
7pX9trfj2Go2XKOOsLS4eZG5OvnZCqqqdKl4zhxqtKApw9wBkhH1k3+4QoNksm8S
OnpgpQE38ZOP1ZiaTliLKi53JEAitYG9nRzx+rk8/Y5Fdtta80si5f8Fpu/lKqP1
rk1HYYok6nSkMqp01ySHKB3uaB/xUCTocb2k3Jr4gqVq4dohikk7RCR7vkkyGqzP
HAjzPDypnUqyO/5Mzvw8Dq1ni+dj3Zm+knKcj/K+j2nKnhJfXfaUodQilx1InqjT
ox+SqKD25oNYNDlKH7GPFgFqN96PEexaMGNskEu7jhidYoJKFrIZqjvC2wFhTrwF
a8SR82mR6GIrkDgTquaeHTwX2sxVz5AC0uoaQtNtgAL7+E4aXD7/BjTVWRluNBbU
iA6POZO4IbnxmPQ1ui066VBg4Q7KxMDrBXauzg0KM7w+dXhvd3daZU5s6zOwKSc8
3bfjNk/+WZ9PDSOKuPdYJsZTKf9Nx3EcKbiznLY2kqwgStcde1nqRlaRVNA/9AkE
OqwYumpgHBwVbcQi9TVAjzaRXJnPZd2QA93n2Olc4Y44lNKPZ8+ok85CVp4KcQXV
luz+3aXXUqgjYQSlEgqkd0/k+5X5ekgWevj8Vaf6swd5ANhKWXTTk8goYM7iHnJV
6pEkdprxOju66PDNaEyQ6CCRG3OqVNCMlWvzLAhdy/mDwsWudr+f92pEC2deAqlp
BhgH48BueCnyIfgRnAQnovJ1gdiUa3PhgCok2Mtk2SRi0l/GqNp2v8/bi3N2PM/P
fVjUzFXjpxhoSWq4U/3yjN1+IwuhBT2gy1SHYbB2qVhB9alMZ23Brn/y9GTk2H+Q
GpqQLhAbbopaI64L3COcAK7z/r8zhIWPYOVJ0pvoXT52vx3hni4VRpYjx+jrVCDV
oA9d/zRBcoFOnO8W8nd6CtMC2cvfEINAqsMNuT/EDwaa6vgltQkZa5cRlOuw9pK7
joo6Nk8bYS+g/K3OCawZGbryq56tpYGWfPHWzLqHozVbGJ2cs6jZXHPU2r/vlDgl
+j5k65KNdMrdOa8UjUlaorKtz1e2GGEF+kC6HElCcdD/oXWipzDTKWmBXKM87NvO
v9K2pGVsCAIfOwe9q5DjD7JOGlHM3g7xkpdv34YuTdVMNuersMAwPWdFTgC6q12x
68EoWk96hmcggTB5VrDDgeaiB57ZVYQMYtJuJBSypgWBrWcMfslzLMUvBPnJldFq
lmXzixKJINf42aUpUANYhM2L4LYJCDMnmyRPLqykx436d/dAfQD8D7fwGY6uyN0Q
osxzeae7uaM4ZGrQigpkBubX7FGXdXejQjLgRAeJ1wJ7GL3rodbdGxc1YWeQ2UIP
SW0fwE6nNQIJMxVB+3x9Ffn9z2FSHwX9CLHQbZJboYVp+301y6KWLxodBJsj3tTb
RKp9JbocaJQdVj1hxjo9LOjGaiACBJjojAmmPR6bYfG2B8d/8H9ZTdJcnWSSQuAv
JPau5Taqg8/UM15wMZ7REsDCdjIXZud8amYVjpgfnIOy9gtX4TGMpVj2qazEt+BM
BLU+9cA45Zno5ETS3itUrAPSCNjzJzDyHCCwNfNPNDqo/MJLJm+aqY2A2tzF5Nmw
EglhYveKkskMBxI4zx1hZjWvz89e6O7GtVrXpQa0JE1V5AnbS4aJb0BrdUVBgEs+
PBJgPh3tslfx/cfKT8vorVwOoCrUnFuEaMFp7x7cn9FSmX8iMb61Z0vUarB2YIUs
a/cj/Kz3IJ9pwcsPBpsOju0SWoEpWSUkukqw0jUgTh1NGF8aGRdB926TL9AszsNX
ajhNg1Gg0XaZm17ns3CkQMVb37tiO8bqclOapP1O3HuEy7fxMkg28RrIbEZaD2mT
1A0yME7vycDhMVCGJNFCbIiGySUOMEanF9+FBV3BiaxqYye+PdWh5vLIo9RVEPte
nHSy85Rqw09tTlx6j9n3jSnU5NJB8DHGiKp9CpMXsULqaNLIl6PejVwK5nex+4ji
dH5gXZ098qQPItRdS8PhEznZllK1LpsiKBoukZ/qApxarTeGmIXhbVWlh6mF2Duo
BpvNu7ARrb6IY0JlWYMzc28UnNVOmNOmT7YUByvnGWCN9NNe5WYriRQAnHwvzv43
45oj/iTFRkzpcXN2S5TbyN9Ph+h0VXNPCQ1vGyJGPdSOm3AnPvAtc3z9YPnVRnyi
UayGi5tQj7DoJetrU3qD3Nx6RxI/W2qjDII+fJYAksHGq+dUa7FagfDyEJ0a7MB6
5DQVGO5vQfrTWqBfO5AQFabOV4Vcgt2XjDAy9RV5xfkBMzVF+6wt7N+roY0AIEuK
57yembdmoYXm45tf5ghT5XMXDdn7P24JVOksQyA1VYX4qCCfLv4DrJ7lg+kz7goh
eWzhkZzWbaQKNbHnB4YwpbFAy82ojAKsgQlSJnZSew4Ow/8nxJLrxCacwPm460w1
IDVJw/tj4YywVx2wMEDnKBviRjkuhgLeWBOZ5kOU270z09Gm8Otzq5dVbYQJtkKd
h4ExUtAjQJmvLAB5NnNJ16rArNTdFL5dBv8w7qBwZhWDG8mUJVkHWhxAzmiRkA+D
Uw808uL60FpbLpOMb2aLDzxpFSwHxp/dly6rIWSzCPvC7kMPelIIuQ1layeAro1W
gUAXW1gIzE7Hl64N9UcMH3EwYTfMBzjiBdHXw+Qy9RKaJlbCdYt0FMkBZbwzQ5XY
w+r+Lgk4V8D0pukN1X3tbqAHSB8lxlGIjbL202FHKl90xWIMjuik8VC59mmDX+GM
fPnnWMBqIkAGTxvPCjy2IXnisxPTaNlISi+xWfzX7yNxej4I3SUHdmTGiGd4Cr/i
JhRPeSTUcu4NuAWOcv7DmHRdME/u34ytaFziPnPWChDeIo0QOtBl19xcHIJuRF/j
5M15XJIg9cuUfZri7ZKHGKkjW9U28JGFi5CNyeE3gBs/wZLFoLctfeC1HEirAxsP
Ou9fdkPbdAk76YYx6hrQgT7VMM26OR+S5wUL9vkE01/uI0dVIuJE9yLsEeizU18S
nE9CPPk1WQGPtHqywvLYKuYMoMSuVXGyLaL97CKdgOsRV0aFBfbOtSrfs3cOC0qi
FnROsfa8coksikd9HByHE7r4Pr0bD/OOwdSz06DrsfkWZmvyNWdMGHoHZuumnupo
/goAX45lYMu4KKaPyuidPAP0kylXzFXQx6gCROrpTc0eMJLzWyR0NseaewRcG/3W
uLNASwfh/SiAJ7vRAOdJ/5usZ3he0qJLQo722cUvuduR3tfIigiMKSjSyDtISoJv
z1WhUTd95+D0giUljNOnG1M3xTtS1CPv/s9WGmC9fp4S2MBl9CEs0knBOuasgLrs
NrVuRd/HMJySnz8Fa7XGdVLFtWLQSuhz0mktuGwhStV6GfK/i/QXH3QpZTlQOafc
xV1Gle3eYz22ZXtkTOygzTquru771WciH2eudrmIW3y7Hz+8brkuJVAdihwhKRgJ
u9qJaiHEMth7qk6cZ00gHmXHtPv71Dpi3aCINi1EWP2aCRFC6PO072bwNtuYXl7z
J0ZeECZ3NSQMiriolgSaWDDsfGwQ9UcnayRLoWUlO3uwgjuUALQDJWFFanCS7Kdj
V1frMNQl0BjfbAke0QG8/v6Pr2vIeZ1TbmvkQhdYRZ8GiFekL9sLTlGHdr2fEPu3
NrRiAyAgXJeT2eZcMhqmC1UivCoBJ9DH8QeQldjwYNwJlUy4qA8EVQfK//6cTCMV
r+rLbabRLbqkoqYch1CYpsR5MTVu+14eC5tOHpJidmp9eo+BOSp8VynbmB9WStrW
GpYUs2TeVwHHLFmw+qaUupgBM0sDHlZDiQVwgYKsyb70G1VQpeyt1/gLOzLU48BT
+7PTyXFAZi50U7sxso2BtQpQaiUgKOG7g5Cz/cke+OmGqWz+uht7AU3km8gNi+1X
qKFI3RJgC+MQlN1O1qiD4v0yHGD/x9yxLrhqDXHMh9id1lLWBis0hN8IfEmHjJD0
QiBaiNEv70soVawSTan4zX2Pw7uZI/5yUYVSB/ZTNAPViAdqFYP3m2jSKk9Sqgjo
tmt0TvDOGMnDo5Q3vwYS+hhe8VI1JxOwXVdDwyMOGFRBM2Aq/yadsHQYpRnbvsjo
2W614VwpYRhjA3X/vvulevsfkRMaxyD7XLdzBcW927ueFUBsEwzK8VDMH/51RkRq
XsdJaUUhrEFBE1K9okUINFnMioh6ep699NxRRWm+phoe1kvX234UbJr1WVFyPVi7
4gbLoIQd72sZfmge4apvLO0yuBrB2BR1/7NbzTDEcI0kpMe4tUmCnRnEmTtr9tqt
HCLZL4dQD+v+vIEoRmFK3Mq3g6qQpyK64d6SdcxdIHVl8UQE29v09MYwsgq82or6
gWQpyqbT9XSJZ5gaw6Hv3D9hxSdP/irPuvQ6Ja6Lz4/nXOMrrJgRgH5jAh1u4tId
dkDcLnBTviMarezNhrQt55qflcm2a+yjH9wiD7MogslE3QIVNZMuVtqxMSdSYJNT
umTp8UFkYlk94cen2oABXbDLsWtmCK9UOaL/ZMJeFs6+dO4UBH01HX70bPtE8X01
AqcayeDigEtgazwcHOuUNZh1UTuhw6zgBuglMSLsOMe5Gc5utFerlHgEkLoydRVL
3G1hxkjTKY8LcDceKaOV2PSUTnzyDWwQo69dNVgrdBWCZdAWFUpejNOcL4Z6gfFo
6HlnCyM0pC4uruIvs48USkmA/sV3VaO1b6nqXXt9SHq26keOskc6e7bPKlS1GVis
L88uAG0zEWEKdz/D3vGIbKngNWxGnqUinhxPY5gW1cwebNRiUkpZY98NujgZlR3R
/mYVU4toZcWRTLcZdNaozIOkboeusLvZcm/JaGYkiJeTuZpFepLSAsFw40KbVyvE
+Wf6yvzugSu6908Z0Yyp5SK4l6yBDZ9726SXPRAd85xj6Em6ToED/FYkCEkcXMQ6
he6R/ovOhwe+/ySxtltKCkCePuKyXETkUdPwoiE6f7XA0DS/GZXj08SnSkezWaiA
DeO4wUuwg55l94vcqoBWXnPUDZfV7Z1VMehlwGw1erMDGhNQdT08V2rvACHaaCOy
LkHm6sGwIDHJbQ71K/EHauNjrBU2M96edhHLl7Y8NvWico8G4WAzfx0Mrb9Uhll/
HZxMjZ3kmn/THW1eJ69r4bDk0f9N5OcrwT9F8+2QRnpQANkyb2xvwMpU6f3OxeKn
0WpdUGmpQoyXg6jA2MiVIttzpPsq6NOLxBhRY555WSVjU4tld4LLba6DZVF4gM5a
zchGmhqxIgYXeKSYlsXMX4s38kI471e9EWgFSWxFeeu3nLKFs8+JzpKYVDvcUfaI
N9PaR1303p+HiFD3kK1m22ZV6bN9AcqPx1sKICUn8klcDr8eE3RrJuvuTtTud07o
nxPwlveyWtM5WqUpUYVF6R6VDNQW3A4weiZ0tYS8H6N0tmYJ+gWUmvg1jqJzHP74
1OvYNKrDTb+bgGLu0JLaPvTxagCjr3w6Vy2X7xWCvGPZBrkuFp4yEZJxMzZnKHNm
rHkxadYh9HnXBtDqIsWzwuFQNCBMYSUw9wFVETcXZdbrote9Yj35ifQFHoDDDmGv
fN2CBLHnAmoBXRRTfDXZcfWta9Sc0YBpZ/JWJnej10Lm+vclzLkhjItsb93XyWJg
rt8YMfOYStJmWjkjz/OCp2OOG0ahUfUZSE2wq6Y8Fl6QJVQCyh75ZFm/i8ZEsPth
HnLk4PytiSrn2cjMnYg5gY2tl4tx4SAQkqAgUHtyKqbepvPdBlueOOSMoExbS0y9
dMqavlbEKZDxc1jKYE0UCLWA+CRFhD8hy3XQ33F0Ps0OMCEuCHHzEn5bn8iDsmsw
y2S6CNJ7EG0VIXGUUHCQwI/iT4uI2VscuZPERWsElvwyrexsTgF/U/VNcBOw/NyQ
Fkm7wuVtXdng2X4G+Pve4zn3QbI31pg09gZXRAmxAXX0KSwtTK1D0j/Dt7uHNw1g
OAu8d3GBCGlTiROEZ2yyZCkHP2w8rpkZKzUZXfh1Bl0uz1bjThrwFdVBXt3C76dv
TJiqQKu1UOILk+ac4sFm7eCTHoCJcMSCAsIn9DV9fOvTkiOS2WsIBxTXVl5GGSN9
OpIEZ3yDf8sFwmThSzKpD4PY15hBv29nOFhzu8ohsEKF7z+fjoCcl1l6agJuibTZ
c+yMixBwF4fYVJkh1mujzKcxnopunXnFAgRuh8Jxc6Whja/CNv+YHly4ftsXmfSE
YiT6ZjRjfeg/EkJFectlo0BuhAicjwWmKFGqfPb58RvJyzZnmVwDrs/CJgq7Fcj/
MA/Lu/pcwZwhD61B4KJA3E7uzXfqTMiRb4NBmEL5tOIsgc0qIuvroWW91Y749ugN
tXOQX5Q4poKQq6W7k7IyzfQtMWWOZXAZhtlGDqrhZ0HUIeAA15vyFD0RrXzsQ928
JBvDse4kYkuaiW3vdC/Lusxg86nJCJqChTXCtXvwdVL36fb9aygACce11ago/XPa
szS2qQp5m4yw6rWm6nrsh6flm7nFE1gKPk8LySODbVc8npMc7/CgXR1oWT2mt2eK
KazlegOvV1sH/DCBNog8mbEXzBK/3nS+zfRHOWn7/lLDaSkdAiVasDeoqnk/IS8D
vPlqUQRuimllDARuFizqwxOuUZlX0DkrT9OEMhre1wehwSIKZvj2gklf31kTtzAC
BlkuN4VUs0r+ovoCkzXa4EZC/ecreAxKk37c86Xn4nUIanfKVRWEd3faSraNoJi8
BHVDkJHz9+yb/z/f3/g5NxIK4Zr6ZrjwsleFQ67yrhWGZzgzx9ufYaiN30UpCJ2/
yfmG+G7oMOwlTIA9+nabKMbArHMTcxyxUEK59Jw/YILC6+pHRbproZsJ0MbKFEQx
7JrrCYXudUoWdwUNUf6oEFI9DEHmKZ2t/LRN+JuQoTcENmExensUS+U56JXjT0w4
aNNDIv3O+W/uEWUkQc4ZMMhadX7EUQj6J487rWwJDM8y3lCmFOCjUopEAgP26yjl
78NuloI6OWjIEXv8kLcZRRJcq3s9TzotOyUiIvbanzGJVoJc4eWIKmR0lSgs8/yU
Vo87bgvGvpXE8sqrViMhBS+QKt/XzPT6xeK4caEAr4OEAlUTwh6A7s8qAgiQC8tb
Bq3jNFFYZoNlH64vUvPTzV47u9kLhI1jKETdILY5bYpRIFwzOkcXp8QS4Oamx/Ti
02MqAwSmPC7O/aAY+A2QCyNLYLQHUuBQOWr4FGl+YZtWd249xyTZipdC2kBZ7Vwk
6XAvKW6aB/LXNEn+xM66Es+lRCvYUpy++ekaoxjaKoynSkp0tQepsnk8KF6S0Xfh
r8CIuCczXGLhAdSITQ66dz7Sa2iAPLyznlN+3TLP1TRVzuc4Eox5IFIWgNTfP/zh
3HfvCWnJfVx7QxcxCpaJpd/qnbLaJByf36wYceeu+4aWfZcbf88kWYOA22vmxhYJ
N8mdp1U2WrnEWqkmpOwTM10bVdMcbpF+AfdQwC7265h4fyQmlbgxYNBNwxAe2xn7
s1h8wLcMYvhzGi5feQ9iNqRtQcNkIL/3ZQ8EKwFB+WJthWSuUIKN1ktjBEq8iMLx
cnIkbU0QN3BgZIEMce1KJIADy4FGLG1wMv5RjA81D4Hgmo7KZ6JYqVUrO9SG3iw+
N8w5PIYQU6KPOd/hnpq3fryZbWduVPyA3SviCExBM62GKy9LnuhxE+xYqkkoXewa
EYM0jyGS5DZuwBNfui3yBj4bZZzahFiGMyQDU3qbWKk73hd0hka0r08Dm+/g+BP/
HO4UxZ4mP2p2o5IeFBhTJVOqNNTr/Vnzsj03dcwoeIcQ6eigsYRv/bdXhucRO3ml
gtHwEd9VsRV6uedEcr+gcPcfgXzs92WCwcK/AnllTnwESnttltZ6jEa3tLHn6rDn
apWYa7YD6dOeA9kfNq9UXNYJbiboUy9W8bbEK2gXwSZ6T/M2fazv7LD/l/XWhtSu
lWZQzIJf+V4606bXH8qTRMOZcHYu0i05Q5v2iUCfbhaFBlstIAteIAE04zv0Q/c7
N+XaLyNv0C0csY/0hoBcDug5/uKGydALA6ujJFvZPTchUD/d0DPKPXa5IecTPluI
hFlscsykPL7thHhM+DZEhSSZ1A/Ak68OO892w49Si3kJ+IAgj2IdK/SD8qhy+wKd
8OOV77RdbMRnxwdx+labRTM17V0/Nq6RQxLig7Er0YmJrFFyUiAmoatZU3Wt2i8U
CAw7UNkmIFV91h5oN8WberJl+3toTiN435jZzpDvkN7VPmZXSkC/J6FJ0KjVtO03
lDt/AvFXnasMi7J+410r0jabvh7JX4HBHPY22wx+Amr2ZJ7dIwadVrc0fZ0UQh2h
kaOMR8RtJociJyCRf2kAo8PGJCSYqNb/o3NnHcpCiC4OTi0Y/n0NCG1fUm5SWaQw
i2bvVGn1ffp3wz5aePK5YsIQOSRvDAMFb281IOpVDPHHoZibWF5xCBWqVFHSRebg
6n2MGvTG1rgS2h9iP9R6MdC8+JMA0DwK8oRFV/0Y92wjJi9nDC61fIuxMhpd3o2c
bfCHs7RhTJUSYY1qP8J6ypNiQ89eEU23k++YeH4DYZRtrUXxe6UNYpkX3cJlj6tK
ILFFRkiFjWEHvJKR6X/wQQuMXu8wiCiscIumYj71/L3Q9i00Dx96YgIJzlk7qaZZ
zsQ1u75Tbxu+Koh7jbmfDs+i2iwWUrKonUsY1jbZj6Zt1WG+dlQLdV6J+CgHeijp
KLS0MXQon3y9rC9FyWue5NjR9WB9XdvKaM1MBoBCbZ6ya8D1xjUBfxONa40tUhnF
GXhBlrsJQj9jx2HUbr1/iovqaMBhviGrTIIBkZrOs9xWbdjq6NHvK5gvZXZ8Kb8T
dB2ERxEqrzJCPPRj/2u2xwnvfTuCD7eh7DxLkgffvh5zli/Oq6ixcpY5jytL0NZA
0iF2fDt+vuArlIQaN5fXpcTiANbSOlBa8S3TY5DM4gWajDYBaGCKB7MR824DnW2F
cilKnhewr58dGtsZE9HMMGnQzHYd5Uab95V0P0S8gh4vNpHjDo6wCBqs7XA6qznj
ltHHoOskOwDW/DP0bOyIVp8k2EpNZWQtoFSvSdyD3JR+2rts2k302MDGdi/05nEI
If1GE/8SrWwuY1sN1MpyQ+/biXudceWtyu8gIUSvj3/L72+eRRol37dnAE7t+9gi
dL5+bSLoGCYsLiCw9HeB+4Ag2yD/hWKw4RNUNAu06TQ9oCj32hVzbvTpoTGff3PD
kCmq/oOR0xBk/UcP1TIpbXWk7EMpTq+X8Y4BMth7Z3HcKdKZtyriV9lPcv5UM4qp
nOnDLe8CY6kKXpXu1mBRegR7iXNk3l+lJTkmeqyZwwKDJwEHB9sSa5HMS/2Vl/nA
XuPxVN/rCmL9C2LT7RzctQbtbUANr8kgplojuJpVDSVzMn3kj4BZuVMWrCQ3yVPl
j8pMPUhuAsDxlUwqrKzij37eQ50Axt2SohpaVvEsiS+PqWD3BcunkD9OFB0/rweD
FV8poaDGr4bdiCLyKaQN0SOKl3oMiu5i3HnHHBGVrir9RJlg68MmSblNYvJyESmH
poI8hHbhBkCvpY22Zh1QwgBneWEpjP/v6vANbb2F2cXz6fz3ZjPaPyRjdP8zEDwK
jLYQqeZkqaNGy8lN8DW+jC7uhiWiRSppt7RB/r02PxCviboC7QDChdopqsIAlO4q
8pws0sGin95CSmU0cEy/pPC3Olz3rm6i2pclFH0BD43p28Wu/jwaeJnqs3haKcpq
Uu9tLJZ4W1MVhK8WPoR2nwNgRB+0P2skDEXSG1e5VysX8VgMHjWOUstAWhJj78UW
p0KvZg+HpsyHQABVGuphiODzE7PCnNT6eA/qipgI0RUvIhQn5oglJhtpblOt0e1x
jD9IkhqGRzuyS+Uomkx5JPJORTymB8YnXUoQRgOz+OodMe0xat4tzAQEqrCmkood
iybYTj2dy48X3pZvCcfp0GmZfWsaDknINbEOaaIU/DW6cQ59/Du98QZeuLZvBcwV
g5aMcH2kChFhXwVa4fpSeD34KE3yreu0w9JAIcmJCTFlav3/Y2LFDDcSTLG6lyvX
XXIvbtUICJCA2a+cdn2o/fl0zYTKfeLLHvA2HGfVZd47+u7WtLuNMfZ6rKAZzlaE
`protect END_PROTECTED
