`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAWNWDRetKCPK/yWvJH3wC3MMq6kJ2KxyXZMl1JqhVqFR
a71U/Ho7OjFEqDci+0Ci10SiqSXePsB95t5aBGEdKNq+ba7/5ncWhV/GvttgHImc
n0ayu28EsVpu0pzDYXxeK5sKUIig+8v94AoHPkRsv7FNaX/pzvn+qdJ1kc8QH9Fn
qFGryG0OyKR8Gjxh36D2JpoQWsgzWd/aTmth3g/uTUv2rChF+jXKij99tFEuewbs
mDq7utGTGC4AYF04omE6NAMgQr5i4g2v3DsGV7aJDwZfO0+Ha1IcWfrSC89wD1TE
rnU+VqIiVcCrLqOka0o+mB7s+64u4QV+fFw1qsY7AIS8jN9IElgLdLvr01CBLEjF
G0bFPnZ7Vix3FAoQSQXXzLlYVTjQMWFiAS6nkRuqpHKe2ZjOCTZIWQaLnQ5+ktEt
QHac0NesgDOprv0Xjd4xJQ36PtwHC3aAQsn3ZNcEvmY4g3KzvzspCpstgOcU5CaS
VvDxGmXeRFELcLszn0w97fhz/nhVH98A4IH8EkrlctnJbmsvWIaBH3FbX1S6YxUx
HUGPwT5xqAlAr6I285eKPsuiuzCaIeNXVH+LOxOfGfKXPIzlY2xBmdmS4yfEvJAs
B7eAPLNnWrbv1T4+fgKgNDsktZA+F5/6Dk9j/U8G6wEdUbNeBj4Y+waIW2dD9Qlm
PJGsiV2It+B0tG622KVrBAKsAKaj00VI++HHorpoUBha4fk6vtDrTSC2Snp96Hrk
cVkyViFAQwtHzOb5V1VWcAX5OxFbvbx9+rMLXDUCqFLLgPFIxllv5mWCyWpJTH6d
IMjvYbl7Xt9vhy4AOT9N9N1EWScymHtveFyFRenSWzA=
`protect END_PROTECTED
