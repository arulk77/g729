`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePgJzuYEBvAvomkXTYxSDzWKo/7W9eD5fO4OVel59S/a
FD54vbGBTAefyftVhWCN6aoUzCe6dEKI2R59q/df9vis6XABgKKtIe53R9tgOUOi
TTyevSW3e+7uzREXil9qlKftiQWTj3z8wjwxyzKv6qbzH58xPewGrVQR6GQmeQT6
rEDFHvgEuaTu+0vHHCFw616WwfKsOU0V2SWxO1UeBjm4bXr0Nedf8iFsE1ZTegPf
`protect END_PROTECTED
