`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SccGu0kLPpsRA4gi6Ykifql+dgyRCVTKrXpSazNGZ6NO
pWAw2TcmvePCFwN2eD5Qw5xCN106aKMuE5k9n84WcUfk8J8KqwgqWcovV3GKceMB
C2r1ufaFX7SolVrOXPMfqn408E7iM35iZJltEj5MpSkCHTVJyx/6f69pP5pFX1wO
T8qFiPrA4P3e311xgLEDFEur6rBQLy8mGaLHKUNg6V3Zhyif0WFPefdgGo5JYBeR
2WdJEvasY1WCKO8lrys4OfJMvd3GvLrzxGDrytGd8eeJZnx184ewrDVUYnSa8aKJ
kaIMAxKXG3+y5n0vtarA5dxUXhY0WADGuGLZnq/BwRWG4I3XwxSNkdngK1M34sYR
VStV3NHcOMsc+W4iYrtTpPFX7jgtHB2qoyWcXZYvWcSIG/lZ3VJimZn9mIELhXfX
hf4KpO9U2cI3+ruTi68Lxjk6zj+5FnNk6tR3qfnRBZBjJPRTfVnQ0g9g2DeNEwor
Ps+SG40RY6OJMd7cbnGzDsK/Es8oaNWobwgFJdVFGKjYbKUprpOJUc2/k1vIv8eR
gY7Ey1BtkrDJqHCLaNFUQDkeDDLFXaaR7Pjuu+Ij2GL+Yq0Z0JczHCdzBN0mTOGS
xaLeMB9IdtiZGUnZwu19hfiZ//hXR/5otbIwxP80jekwqv1HBk6QvuYYcztYo+wP
Bgio8fVAqkDDDKoK4kJICwLVCxV7yc1K5lQU+4Klpbl0YkhUzoLNgwgOM5EJR1mi
Xj/7vks21AeRBUbLmqUUZwyb1hCXMA1XD3C3FhLoqJgwytOQLS+o5KtvacHEDxWd
J5LxgDdVseSO0BF+Hu3Lru4KVou2RAuE+4k6+q7Q1HVAna/vElvOiNspx/ct6+WX
HLpjaUbe4+y9YTIiroZKMRdYtNwdP1MiBt45F3DAqal98+fTeA2x8sGTbTLB8w2s
`protect END_PROTECTED
