`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
AM8qsSfgAyX7SuTM4ifTf6uZoGtw7U8QQUwjxMLEYn6xgqZaAjwQqhsgLE3Og0iY
Z/oZ+3TjNiSv1DmpOxG02kSvzdavu1SE3bx7Ww83kduznYVBRp/80ooZB1BZ1Sl9
dj2qMaKpo4pzKjYTQmhbJmWyygDl6un29qjhV3tz0RjCRKhIUsqRNVqgXztYaHp3
Zi2KaBjLO8+26PMgoo9Up4YbJCn+Vd9am6RryAW+XFFCni7lLCDPyoEwGF2FBnJn
1DsOCPrKnU/caJQA7LkFDhVGlEkR8bSsY2jTYM4c+3rS4UwkjLB+nUZXG6ChUNx2
Q7i1jIlYqJKJ3hqCuXSu/uIjn7NqXxrNGH8ZzxktnnJbH7ACcoT8kcdBnJGA3B1o
DAtheZT/We30HeKJaruqejvAvzlkS2lCXhbT1MzeZnjuxHg/tEJBpTilTzO/tzTe
TuYvEZZxn5jXbD2zEMB77eATN7qIUrQJP69AJpsCceg=
`protect END_PROTECTED
