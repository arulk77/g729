`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
gWXuTUT8KcG+z7H4J4P/vGcfzddNUJfpj4z2tydYz9weCSVzCyRRqs5rYy/AH6Zq
m57fF+WdorBgBFbDIsxyQ8crBpXXy2HwUxAgJKiWRyZZWFaZF60PRbdTpZBBWdQj
kIYmYUvvoQg6RKSXw+sXvlPI6t6X0FcN6YFBLVc5VALmDN64M068IriO2W4AGFeJ
rPR9LZZjAkDmd/mS2GZ1a5aBVkspbrwZqlxEsTp6C8ohaKNBwJW4dIPTpbEzGj3y
`protect END_PROTECTED
