`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGSA5N7l5T4Jn5lEIm7bTKMwiv7s5HVio4m/ezFFnOdM
TS2m5q/DbXBWpsN4Rh1do9ORfKHcPht4JKjgkWc7ub2qIXEBalPRS03oHyO5FzXN
f0RSvYRvXyzbh/0gMxMQubF4F/ZIIoMOHIzjHZQ9H4rM+SSw7bkh15nzfENJrZXi
`protect END_PROTECTED
