`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP1K5vCsupgq5MDLbv/HLOAvcL9yzOPX6D2JjW83Ul/J
V0POuEjp80ILXteWoBVcM2mg24sAN/GQtvt7JW6wcziDllFm0bQIBlcjptb6gofF
3tNZ8HvbLjbJetNqdAb4afMlsfO4BGi/KcJ7S6DfZC6QqTj+wV18JZUQJwLGAbgj
EtzJ+rJ7+xSk7bfAqXLteMVTh5tnZSNFzg2cVEPGa8+4PByutm+weOs9sFVvv+Yf
AoWHoYOjdxfEZEDFsqhbI1yJDAvJ8t8BvavXGdZzXc7lSPAckIc+Uiq/lLW7c5/C
eKf12SLRgi9VsiCbGmJPchNgt5hs5RQ8s7g5uW/SGN49ieoGXDi36o6xfDuZDkDn
Xi67ZNEx4aGDT3uFawUVokmaMj/Gten/vTtv8kKuxWM5nOdeL8URcSIjWg57m4Wl
I1inMhBCTJW18gPI1zGr08emZ6bejHiT3zcKSFb9M6tc2f4CmOUT4P82B7QjZZU4
`protect END_PROTECTED
