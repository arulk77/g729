`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP79Va6zzs5B0Kw9cjQERcLmvXqCW0ZPtnv9gyOiTHIB
T5csSeZtClyY5UcQs34DRz0MiIHVRefOwfT6vvwkOQAU7EFPHMWch3JGcDc5WjN/
u9f6wKvbiVRxS076Mhsbs73xEuqBGH/LZTcJnxHM0gPChlKTHEE76x74tyup41cQ
PaPdcjnxFH87dQWiEixg5f0O5WdltsTcMbI4oKhpNFhN8XsaD2URfSEl007krJNn
lzx/2S4ril8E17t0KqjveJk3JiE3LPtTRx1HVeraA7WBB1iDpIuweY+kVC4xLrC5
nmleH1UgiGFCd9lP9JWKhPbYJ7O5JoyxG4AzfAaaDMR3Ew3zsXJvqrQw5K5gcE9S
bqXazuEEyew3ZVntaaKUuNbPZHIL18irgencb8raCPQTYVtEuMdzs1nVntlClmhU
GAchixOCSVNT9Xism1SA0pC+lW8V4Q7+rbAc1NcRh+MhCM69XCNh3oMNqXvAcU4d
5+thwq7KHqgX3ZcstdeUPw/qqbDe8PRrBwZcyuJJRTMdsdHH67wu+t+k08suwn0t
JGhBrPAchs+bXX29d5KCVLYnZmHbqyJquqn2tCY299N0d728+4VZl70JsVmxxJxS
GBVzuQIvGf5A+6izvLRLs20xejlEzt1zccsAReWm97Tj6tP2C8+O84w3qkhnNbJW
bkhhh2Lzmb14fn9ooKspWvPitT+149f121IJiiichi+AYYjFVGxB5O77pXIfIO+f
fh6s/WivOVQ10R9QkiUdu/0CjG0wfH7YFkMKPRy2P3Jo1wMC8B3FqMFsoZGvFEg3
PuUzSDruNhPBZEdHhnn3tg==
`protect END_PROTECTED
