`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu454kp4t7af6Jo0ei75uKKEcM3eq6cmsCfR/MCNsUCore
6J9sXeuMEEVJfo0WO7b7TMhW6S2QgpPb6oUi1Jg2xR9NCxi6r0BS1zYA3ksK06IE
wd3HQPun0CSpWtjYRr3IqkNuo9rbS5RxmWyKZIpuXJujdpwg+Ld4TrI4LbVORXIm
shUik7rKcptVd3gwCo37vQs2ggUFWnX9qxEDeF+ol+qiuCuF00/MSlubeAXc9ZE7
1NFxI/Oz+O7m1018G/Z8Bq/iCldPMsjz1oYHFuIUQbs=
`protect END_PROTECTED
