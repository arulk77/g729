`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN8i/kZMcbMsS8Wuo/bRYRBynk3yW6biGYVwP2WCE5P3X
So45+ONxtkwQ7FDR8aqsjoDJDAqfc22Kc5RijmxXzIvdh2MxXG5JCNfuBEx1t2Y0
fUoacDDpbHrgnoAfvC0v9FWqWQW8qSMCKCX31+Zm49Hdbso7VVzwlyDqEGJAPFwv
qNp9bG0AhFOOCsrJzbD9bVRWysZvzMnjmMhTKPPrkM0BgfzoB9PYwYj+TMsURkzJ
sBIIWdGnMFkt4xoZT1zofT58re9nlERtW9Xb189q55nGAzpBuTcNpUXRWpUswHUX
SwB0DgCmmNC7KEDxqIr17yQ9/e78U5v1b7AeOfT7Oa9EqczHSESp+kRa4df/D/rb
vNcoGVHp0ZmvxJ7EIN6AwxQDCFkj9wCegSn7R7ZUhVcX3CVl2NLtWgs4hOZHJUoe
R9iTd/9BU+7udGmkli4jjXfj2DkUgZcn6IOqLdJEnkadapcT6cxZeOZBO80LbD/r
IiCIa5mOBptK9HYSx8dF7mlCfPo4Bg50NNZ/k6SCIeRX7hPCZbyLUAvprM++vyPB
mjUHwtDX/5wq3NvGnvEzI/NJ+0aooxSebnr3K5bN5+8Epm/ED2N891K1pF0lBG4Q
gT9b1sxER9eI0SLox5e+MHw7vPpqeTGg9EkEMuekPKULzPFe5Q1OSkcWRiaqDS1R
XegvPrEg7YD3R4KU5XdwXBCkeTdSljsXWwiQwHBVDHlA2SbBNBP2j4LIxCGBpLtt
HtME3QUZMmpuvG4au7/fHXB/2Y7qQZyUOlf3mZjgmZrwcSQG4hW5KrlaF819ZHB9
ZiOz+TdkRJyWRkE/oh0iqyFSvDnXJbBpz/5sPF3zPzDQ+1XOVREpdi3oe1fy0NxQ
3aWuTkGvpxIXOLNyQp0Xpgxgx+rZj263MejLisJVK1ZaoszvtC8roGB+QWvNu3gz
sZtsJUFdZPXdMt9zecSWOsekxiQTm4D+dc2cmkExS3rMaMC07HlLm9WhLYtW+uEn
WS77kqHFgYCTzCSkfLgk7qhFa0MI6X0sejb0cSE/95h5cG6QfQ46N3+nI8N09i4n
oZ9rDqvWCrJ2ItJwKWfbcYlAtecwKE19qkCePemBUh5MX+9bRHckJbby54VEgI6m
mqVtsUxNE25xjkFLOZKxNvKw4PFOgooyDUSSe5meK0lWmQVH4/ME+ta7Gcav9qxi
28R1RzgcZZFUMJjNdipJFr/cFJXOIZtCh/5GB/tGdXcS8v1deIubtwB7NYY9yjIM
OP1IzKLFxCvA7QyeXnj/dBK1WdfyRICmhmA4oBB/6PsNAX9KAw+3hn8KpEgGescA
RYdnE1LZJofwnvuhxgLaM1Q+VQieeFcAAmhlnpjEn/r+i5ZUxB3DXM0nguteuKNp
L/IpbaDQ+jv6LN6A8k24pzdlP9/Pwrh3Z7A/g0DYXJPTFVUk1+8mwYBwDKIkRiVY
U6hO/QNnPTk2vHk2a//wpoy9Wo0BkqsHw3RsKqekW2i2wgUFWKbCT3P2z4/oqgs4
WxWbhbB7/KdKbPYIDRRMYEaPvU3s5FCzfkFk/sjYsHePM5/fRctJ+4wO6B4VGbWI
F9vPXptAIxC+s7SmAPbD0pxS8sngiIw4Lu6hurUPdeP0FH22ZWKWLey17nThvOwJ
/aXi8bnLQNUrXgs6pLdAY4TV3pmo98Emvdw314GeUbxTJV1XWl+UAnAemj7Gr+iY
+N27Hwt0ho1ZPxQ9RbJX2JO4JjbRS/nrARvJ9AhrhWlUphtnSyAt98sHfa5Z5Lq5
/ntZnCh+z1wt+xn57f2F31Y5PxAwtxc3+CgZcEblgsT8ql1XL9e61Tpeq0PTXHHZ
cz3YxZwFrLjTI/A8Fj9vIp/HWEjd9Q7v8dLZo/pMFOlYdKv27Sn985RHFg/8FV25
`protect END_PROTECTED
