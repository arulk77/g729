`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4/djxYQctx9WbGBXNaPzJMfJ/V0i3Skw2yTBNdKcP0uGCb4a5QiuhT9L8VM6DDmr
H8fzNT59oQt3A702z4wbX2LmYCudCajLO55q7Ki0La4HWW7l4oNxkkheTjQqmXmN
wQCy6jA9AVi3JQyh44qubqRptSa75DrcimovWUzt3hjF7kjxa5Ot4pA6RHqJhogg
egT8+QRcVIHWNEKYOsyuZft/7eJQt/w2nCW+gFYpb60=
`protect END_PROTECTED
