`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
vQasLabjfLexWU9vu3VEYArmPfXeHmwzRU8DxuRpLpOCRwj+hdn2QD9dlZfgYteA
GziL7JuDzATU+m0ryZ5fiJgi5GbWpEDbpOoWe262QTKAjtDK4RJoNF22bkmaSgIk
VzPmOKjupYi4ckaPofcV5DgRZsz8zC02ZBNMCehZQTaH7VYdWDM8dy9SJvWJi7J8
+J4hy5aQRc9WBkhEU+16kmWzDgA5/D7ocjWv0E7+DTTd5w775ce0KO+KKYq71pOw
X1BPDMA4cRC2E74AGgCESO+Vx/njisIcSYjd3KKkLWq6Zy0pwYO3CjfBIgZk4Eke
joCghZsbMHX/bOmX6mw/RhmU5GWahvo5yr0GWy8azuQNwu/92pJgNeSKZIrSrGAQ
0+y1wXz3A59gFvGmZDsVhErJe/RR85nqdyRN14UXynF9DT+FfnPpjbpL2tuEchyE
DWwcrDZaqmblE3tlbGtnzLwOCLDCBNVUUMyXr3cH6WejNNo8KIfvLHGZGuB2BDYd
0DdEuk9RLD1ESnLPHwzqPXFWNLy8CanySC1ZOc/fw64fWdonHxUG2FYDdkShjbc8
sq/6tkdVOVdEZukcZr2D8Gs1X8xeP8/XWxNfL6Rd3VA3AsmHKVKDmjyUY6rXL0iz
3/Da0NM4wq6LNOPPvHjN+9JMd/ssqIAMg6/D4KlXJcJSIaUY973menZxKGqbk/mZ
x6ZS7pPcqX4rwq8jGRcqbLtBXSHcXJWm1g90aSbpIyhAOIs9eM568zfEpV4TOdds
MQsF4voxcapEcbMKAbaZOhlziDGfiQH+Hh4ZL2+xGeRXB64I4gxvWSmIhTdYHgZl
kpxqgmNelJEMcMEYW5U/MwYnIP9Hbx83FfomTtjSp2lvv7i+TlWxBlP7XEGiCNRQ
JXvGdauhGAsMY1xJLcTVNSnJs/HJvSNNctGGKSt5NHlFuwcp5rQX+wcYDNKpOUAE
uRKMcqBtm6kEVJI8ybLfLY8Sp4s8B/0TpxgYzVx/RhHv2FoBUo30aozvrtR4PsFY
dEZIGt/PigY5EBp1KfI8EBVdlYBtEbb831Vqo0YPyn66h1aelVgXiEs1t95wyfXz
`protect END_PROTECTED
