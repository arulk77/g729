`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGQeMgyQlqUqAJ1JQSpYxgDKUthPZXcnRpqcsml21kij
WxcuhAKi05Jj94lvgwrRbcqWkDudO7aKbI/lyIJ8vlAhl1XIzYUBaIZpBmtLDsCz
3X5GFYzcSrutd+H+JvUGZiO4S9KZc4nmoIZvoy6LI0tjM/DfNbRjy0BXT/Q48ahR
2UGSs66qRtEmKWZKk/Mq6jKcDfBibflK2Y9THvYhp6rZWEkYnrPCuC+sUSTXLmpE
cQLAkMUNTlifMzQSjKZCAyvVjtmlOkiBCZ2EDoN23UPHGi6fhwbqDXeWmWVUL1Bs
NepVYNHc2IWlgyv7EtFyj5dZFnT6fJcv2NFzcusuUQ83hN3epS4RL2518+WapWGO
ztiZAw9APxIVHz3dWsuFwVqZxl0yW8bLURxA+mZ7Y8c/B6kj5sWPrh6cLgzX3xHJ
JqD6WHYVncknfmJezNlqcJaCw7Tbv5qvNz34Wi6QwS9SEYnp+GXoN2HRQ5S6e1n6
/OhzA3A5yWBJscsFf+2ow182Yf1zPFMXVhLkJN3SzkYaiSYQg6x7ciQGM1IofUOM
`protect END_PROTECTED
