`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDApZUoUyilQNpT9ijOINndt3CblQ012sgCIPke7z3Fb
mR6WVwp4eDPGUtNaH6Ms9Y5l3C7d5JR8rL9N7/F9vYRNNQ09LoPCM2NdQqrzhZXa
DBbmpitthywSfZuV12Ppgki60gvZ8QX5T6+VIph4xGmi7M9SM/vir7lEBTVpKZz6
q990WPPsdGgIhiGtW+gJXa6cfRlo36qkY+s44amPgEpXeuqhquT0YS0C11HscncA
7x481k3kN3Ddh4QiNgNx7PjnMCLV0FdDcVS1YdKdpzWmzb8EhDJ/xZiO1bNLTvT2
jxT7ZjDe4C38ME4jiSkNMtp3F9RF9OVpV5v35oDz9bg7BzYY+zs//yS5YdBiK8dw
u3nrG6H+3sfS2p2uxrN4d6VnsgooiiL2/eqaUu4BTV6zz7Yn9eDzaqXnC55/0ZJU
Nr3t0OouTxaEThs1D3IIiYBfQiw11gCI/3Y6C7b+K+FwitndhrsKr0ru2YYISuQt
`protect END_PROTECTED
