`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43LN/t1EVw4dVDsJ1jlg7qxxjfg9qO1obFiw1tsLVrjh
8vkJ/ODQYKDx7XgtQuh1oDaXXZ03RY36YqsN6KD/swZa7/xGgaYbyCL+dVyAyQyp
Q6jP8OL53wehuDF/4IL9nNsqJ6oS+5p1w/l0v3czuHtWEqnsykSiZvunUiK4gjkn
6+Mo3Kqxqaw0LqqPfSiYFo5Ch1Xrej5Jh7E+SrySDQ7IYfFcwuwM0pRGK8Hgh3gy
qQX3V/2/b8ef8KtQbPPCfdV5H92jS1IIPRgKdpvUtRQ=
`protect END_PROTECTED
