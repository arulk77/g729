`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45/zU6hvBNtS9jwbWro+ZHjwm95Frg3w2rGPPu2CiRb4
XId3ijK/uPreqJEeyXM3OFQmoYFp5NHqjW93TYN2BncG+RQWIT8LXETw04aR79th
16p6Zj0txJt3aPUA6A0XLqrrpgNl0EAhHPn+JGod3mDiCPdczlT+sEvb1knwEWw9
sYjjSFsTu2ATwwh+MGu3Nn7eeod0f/7miZFDcdcg4KbMmdq95OIMP1uRLTrM4m0O
yMJonN0lqfDYUmO4W2Lo/uFQmINgg4os4J7iL5PN+o2rYw0AwMqwwCGfoKNB6s55
y3XN5f67bkkTQetNLaFpWJjXi/+hMlVJTfuM2gDGUkvoi/8o5X4oSxB5WV5bEYvf
9RtvON3dEBAPoYpNgk1BVQ==
`protect END_PROTECTED
