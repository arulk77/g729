`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkauwNnCqO6dnwtypLDQ/6lATVc3IxX/uDXf4t2uWIMsr
pdGM8H7lKFuVWS3+pRASDWeApVfJ2yWj/2By82cYK5UqQIaZyTMiGtT7XURf6imC
3FwPEVnBjxVWIn5tarRmDpT0aH2IBkN+uqUzWc4Dtg3ERpIED/gQK1rdxK3bqtmj
/SzOVB0SNgvSc+/2H+gbfpvAy/WVBeZdeqNPoxLWajO/rRRMUuIuuHtMC0SFrrQF
ceODVG2cB4ukv0OxlTBmuGebzbR/HAYpJXwnwGJu+GvmpaJlIX1kCn0dDXzgx8IH
3gFpYKQvAtqRtmGdJ1GrNznG2wHyC4ikJfaVMAPnCgSjwwlcgHDN8pYfx2bPvo21
MdDcexS4r1n3HTi2eS1LNi7uY/poWVQaJi9Sj9sgbD0gDu+CIw8AhNbtEwErY/gg
V5CXxFvWB/WpBr1uVLnsPAgqfVtyB7ri3it2UBUmAJZVLS//tmjwgY/60nbO6zDx
pXjPCp9l1uOWOS6SZRsx315bmjERD9Bld5bAJLtRSd1XugoIXq8QY80e5uchd3qU
`protect END_PROTECTED
