`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8ScdsPDhqoeGWJvHqQriZWIZrZUxrrinkuLQR29fbTuVi
DlX7j9Eu278UA3mDMqApBtMuWgJnb4s5L2vgNLC2Qlc5WSZ1HW/V91xGQYzQMZ/R
l2twmSqeUOct1MYg7iBO/8yWr3ngXrig2RKcbAiKIu9B4VhttbxNO9BHmS5FzT/s
DhlqJNcSCG/0rxmgm5kXVJQMG8jzgjeIid0JTz5JjtYphRF82/R6aQu45FT1gx12
Jlc+sJZZiR49xtfvVcSMEsGenGbWzAa3Gq67G2KSFlE5zdHTYP9GIT7UiTHNOEW7
e15vEAvos7SQcGYFrXl4XZoYkYy/RUoQxFqv/QgS8OGO1DbHidvdjK5pXopu/uue
t+/VYgIeTgl9r75RpPrRWhnJ5YCUoR/pNt/LjA3HvZkpG0en5rIzZFkI2srUX4n8
Lt59p4VzuVPEM2a4aAcGWkA1WZpqdE7L62b6YBcOWN/vBbPpeffCPcKCqBqea+P9
/1JbTWO9NMccgJhscIvelIbK0jwDPmSrKVuAE8eBGlI1ynv94sSP6957M5I5dpnY
FgK1ozxu8vA5sqt5w866QTtY0tQUt/gg6U/ZxRvdYpQxb4+gAEui2v0zrevEnWHD
wfpZ7PrDE68HMzAy20TD8zOkq+6hT/10B9/Nrl4d3K5vHaNOEkHjMk3U0cqafrbs
gbvUj3NTC+aWPzHWlkXYAJonRCilnXxdyL7OdG5n3zpA1kAAR1U6EfP2V4ETOSP2
2wc7iSnBQ2Uu4JKJCYHYAMppcqjHBTgrNwoqQoX2gg4I2BR2LLPAU5qSm0ojU/AC
pIdhY0bo3Kot9z9WKSK01+OiYUdPgbyDD7hZA+SWZlazJFCDLTWLN6tytockZUac
bKwTN+gHLXCls5uYnIZoFfOhnBoWxXIaM+G7Ez2hurjoeoXDhOAl3jX33ZbKNL39
dGB9vIRHlxQ+QzJxuZgQEWNIWodhJ7UjYIRutfSBKsnjHcF4+uEP8tqeqyKuP+cB
MGix+VznHYNTyVbFZKx3xG33n9zE/wcGQKCIRBx+o7RMJVYUx1X/HiustFvgTNrL
zQE6gJlC/PyypYMJ8n+NpeUvDjWtBugr4g2R1Ysm56mUEHnLJTCwJeEw23nhGK9S
JHAqbUDgw6GGrFaq8JsgYktCKfFbwPnDhmdhJxWmxr7+W3kJs+zevaQ5rF9BW6Vr
vP01UKQWxNm9eD8XxaL8mrsbvBICHaasekTZW2hriEcfIboEWrgdVxCygVC2ebX8
psliGi8wgRRuURk5TY02sh+yLBLBux0QPPi02NGudFj/8I1uvo8zcAftn8+N2CHi
POlb1e0o//QrpTcAMnQwYeBfqFtx7mS9Ua8r21zNdA1OwBHlCcLHYcPEJtO7XjfI
6gSeaal8URTBT/dV8QBhfS6GnQGeztz/XdSAnRmGgRvB9j8+psBr5piuxZIMaYRK
gpOKsrtXfKlzv5gSBTN+jlwxCHjDnxOT4izIEbSWoNKq1y+9QL/uAaTDtYBNOarK
zPt4XGdW6fNVOoCK0iLzo5SQW8/yTkmp2toroyGpJUs=
`protect END_PROTECTED
