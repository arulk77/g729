`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGiAtF8cTaMnwtaxzlZ3S8z4kYn3incj5MF6DXYyww1x
0PAx+aSb7Sx21jb4bhhBBo9s0d9G94XWGs0OSLo0AXILtnmQSquKLe7yNtb53Jkp
jq1rOV+HDPwWUOBsqEFM/tltrA9o9cIr7jkiylNL8qb6593QqyIPH4btCBwxYWmn
jcXhhkQk7Be1h2/k6j8blRAV4GBDf6zhakusUTyCeRTHoqMBz+MEQX/02amu/6xk
`protect END_PROTECTED
