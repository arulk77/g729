`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCC7UTY9AsonmA0sN47bYFM/AhSq6Izi30iwBNsOR/gh
9YFsFNtlch9CL6Hr8BS0hRcmJmf7nRbwInVnpgbjrVXO+VAilB45zV98Hc/ppPW8
Oi/tO2pwiBjL9RYYAYNGvoEx/ttgoRKUjC2qj7aT718zaOEl4Wi86QjVlAPP90O5
pNgL73OnBNnAIMEN9AcQShkN5VdSpW6ZGX37FRYiOFsrQgqrOGpVFs+JOMcyIGZy
ae5hLV0y+1HXXhgns7atBJc9kcvS6tefDwmLU6pTO0+JAP6NOzJ7rsW02l57kLHV
aHYE/szrDJ4pIB/G16/sgA==
`protect END_PROTECTED
