`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJT0PgjiCLNaTMfgAbtVvt5cqdoz6kPFnQ63LFdtQ1pu
TWJ99LMgU2s5XFV6kSLE9F6apGTOC2FNLmu05+LX7dbOgpH8CQqL7am6W+w7/K2u
vjw6osqsziaGupMm2BtCmmTDVs1v0vSXP5pH4p4lNn7PhFSBsz993AeUIna08tUv
dM+PBu6EiCjcxsBwAgtIWZyjpA3TLepS+eB++t/1O79yxVFFaJ/dSF1MBDIaXnBR
`protect END_PROTECTED
