`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
nOgNpicRhjMj9TCEj9siVdcLBvKxITWJHZWuRlBEZ2vL7lWQBO9JegaKRCqhydn5
CaFjq1ltdMscHZFE4jmbOdvhH8oFlBOT5FhKWdxPmMoqADzDfDJfJEhOK4fCqK6e
2UNKqpbEyBEBdtGMmQIFQ+MMjBwZzdiYcybav5baOZM=
`protect END_PROTECTED
