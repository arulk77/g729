`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkS99db2caarFX3uDW36cbq0zv30cpaY3IhngpVboX2sV
0Wy0D7eqzcR3G7sJmnBHPtFsGw0i8NwoBSHnl8l6CT1SkCrIG3BGvRpMXpED/hzZ
vNhYRNixHxRpEfc0esf6/vr4j8XQJWQia4/XFxBzEcQaHecHu/8YjRloJZGs6h0H
Lw61/dUJEv/NFbXiSyUPi0229vG8mh8PlqjttVZj1JbV+VVxkqFpDxR0dRbLg7LX
/7xO5e/kZkOi9Pjb1Au7jDnYrI9fr11/du18EkjFMez89nTM58cP5zvp7MpjtWbp
7TMchgxC8aPZfPDDnI/Lw8lhjUb6DjcbgLYBFOJQKPK3858RPq+QZY4O7VRVmpqq
kS2qRKSlxrNgjMe5oCG6px4hlnBhLmOqQ3fg+T0UQWAjfjt4tSbQ3rPN5FX4vWQp
9mxW4dU5uJqFeZKkYHv5/d56LU0OdImKZcPDT4IkRAcAhU8pCVnkSET9jc6GkojT
0FOSUkbz2RbaoUeC7HnocUce94tITXrpEXgbsA2nf+jPZ+9UGiCN1B4zpGlZOH0p
hRRtlSEfIqldmTs/YIMC+YNxjWrwXSG8cCywT4x+1H4mmyaHVCePWjnuSJuuFhWL
kr9ipFK+WJwx6NA0KegNFHEmhooCxoDJUrSNPC8nhPe+Ce9tsazX7xmWnHczRALA
9wwzyiJV/wpG8F9oMfQtEALUEqLCOSchUd5Rn+icDEbc2++QofejWlrPaxnbrfDD
dYgX0vvX4d7jrxE8LrQlxXUg3zE4URSOe/ToP+ttNxvEbjm3dwI8Cc9VEVBrgfme
TYjRnSPYMXGTioSdByTl19j7vzNoL4r1hQZ4BRz0lvpBxZ+mOHIVMZybcpccPfrJ
R6ti+m1eROwlCQrrDHg8rhQ8umxN2erikRXsagof8L8=
`protect END_PROTECTED
