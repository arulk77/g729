`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP+LJVEUDmHH3qZxvuVrRFAp6f+FnWbNhyIkSvkFyx/o
mXQVSY28krGW8ir99ZW/dwCxphJIs0cV7gQ5SDeDDZtRGiUV2JN7o5+w6ve5GC6U
56xbs91A2mu3ZvWwjJVNOEGHFBGBX/eq10/b9DiBgc8lDkulUs2qyR+rrncNv/AV
Hkfv8H83WV9ze6DEyzolkwrrUZb6goOYng/sQ8deE6O5bZOXYROMkd1AkYBtnNvW
HYCGHO10+GHf5YxP8KSbLo//mfsTdtFl9W1EthQwuDzIpIeTJJ1QfDmOX9soIoE9
18kwbBbIQqNX2+aA1Tr8QnKgFCymZnDvt4L0KWTKpuPKVevw/7t7Z4BRhVY5xm7C
ScDa64RHj0jXkaIhatQqraVC34ARMYebilWYeXhKbNxrvU9Ua7pyb5ZVvacA4oyK
dSZYRzUpP1ib8JhjUimMD6oy8gtb9WP/G4pp60ThMHHreTtN89CNw6+OGrRpyQYZ
aiqSQQraMwEiiQBjFBIf9z4uhHmiW0X4BLn/MvctDCVn5/oVDzuHN/B467d7zglc
`protect END_PROTECTED
