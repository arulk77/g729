`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
YnHJjWeYHzFEpSOFDJULgzanm2dAoi+64MP83zDC0eWuWhAQrPeM0qPt61Ynv3HQ
REQy26Z+pRW3V0oiITZJ3TJfsdctY1LYsHkAN5cu04z/x5yRjUos6nybLacdVqde
5Sg2HAo/OEKQT87k0OUsOvCsRsH5O5Kfn9jHvGv3WQeLLk3sP3TkPgZMeWTZxnx/
OwaEgH5svwWG5ptY8CzHliNfVvk40kmXPmwbnGOHnN+Z5SOZ0wQP6K0P/p2onsum
j5ofrCQy3V7BCVcx/nO93HKs29iXaJFbwJwBCFLRAtQShS2YpmKtjMQwaFGNISIb
b9V0gK7VSOLnLYWCIBI7VClDjjebFcz5N9Xs0XtL8TIGJwmIQnxUy9Z9i7LP/lj3
+cliSNqTvePfQCER3BHj03DlqhzVNFncfodF3DpN3rsph7CRgDz3hdqfNPzRI+CJ
bLmGwAiFLptXYpO464PrwOz7ngEx5sXNwdASpg2W9nkAn5Y6zTGt6OHGFdgPcOj0
EXf5hCsX3Aq2fj2AvZu+1PGjAA/LRIagj+azlP8TmgrBTfngb4fGJAJHCu5Zkn3m
v+Y+SP1XjF7l7a2i4gbSuxYhkIRT6pkkxF7eE8Gx9AVp6kljRK2Da+525QoTaQ7A
9AU3j60aZiCu+9TaZIkMwRgVxAX7ZfVIEbuK+tC88aCIbjixi1biVxQmleE3o+i/
CEO7n/6KAW+EIWd3jVblzY3xBYpohqv4nvbKh2uZu2Z860B2nhE5DJWb/B+9krsE
B2WdmZyT3A+nf6b6EsK1Mlfifylv2qDMLfB8PGUSREYjShf2ONENeio6nqpOcJCa
WjeX+JHKOrb3WqjDMf7qqK0whlPaPfhyiC/c4jqfElnleQRwiL1BG9XRaR4+ETGq
q1Cx4Y/zDX7CuGAqhPCLxAMIwuNgZk9dgyU+18l8uKUqINxn8jb9lW7gFwm/RmRi
Ada804PqbqcvoptUDzV/xivEV56Z5ppjgFF5j7TQlLkIVmiGnY0372+SfuP5ns+Z
s1dAK6qIZoRgri0Wdl2U7g==
`protect END_PROTECTED
