`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+4TMvXgxXk6u1ZLhV2ttQclpR0FUdEeE5WRiaSlTtSn
MstV4LYYvZvarfAByz/aTkN63q3Wuf2ltmnVFeQIAZldhjkPP5a0txY+EdCRHmTG
6n8o/pK7CE9H6mmjzYPDw4UEcoqVch80l9W4jpBa8gspTcYwIen5K+IBjiZUHQM5
qH7RPfbuLSzYtKwDJt5cmg7fs4C5o0HF1KdgBavXBj9rf/dvUa1UOyYWI+7E+/wF
UdJHLtCKmlNsLg27AoeAVNxvhjvW8K7ravLVf7UvLj1/C+kU4UwPdjAGktcB1off
TR6C4YtRbwvs3LfuD2h6gWnvTuudvsuyYXr2GCt01OUxG6r88LdC47xRHl7i4ZpV
Jm/Px1KbUz9Vc2s3ZGg0u9yoKsbSpKOzCV3md3ddyF6ftwh8bOiGzPs/Xzos22fG
mOGxSl3COQodBurwjSMFEK9DmZ64M01pdmKz8ElbHrEAjJ4tG2IZ054dMDAl6omf
`protect END_PROTECTED
