`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xel5UJKmwCsv1bJmQVQhdomMitdFU285aqohiTb3s4F
jhanXVqKDSAaGZx9/mNEIBPu3oQYBxZZj2wMR9MDCjWwqwwmfV4Fn/zCYazHQkF6
ASJX5ST9LbIPVno3E0Ew3nJCJeznpguAjfvEamXaNnEcPh4vH9UaGuNkYyfi2dPe
+qXmUP/VfU971/IAMYUIdH3cBkwYpw43p72CSBGd1fNVfQacaofH4yyCM1fM9tRW
syn1ceUTKJZFnMVaEm5c2T9Utb0CaiIdyz7hrF0BPNEPJSmm0h34pJ6e8ZDkSbym
S6QhGmZYfS78K+U3A4FTTg==
`protect END_PROTECTED
