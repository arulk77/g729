`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45Q0++8YJTfma+RO+gJy4TNMHcG7eXJVSIN85eGVwH4W
DC/8x4bA06kSPDSwrRvLDOOvxPdJ4Q+b47o7X6e4V5b52vWkG6seW0O7Pt1zdF/J
kCNPehmgPeVlgGuXCZ3k9TzVrOziKx2/7sdF3bo2HtuUMb8xjIxOt2uIHRBaY59f
6xj57DN5QDO01wmWrfbBLbbOvSjSUxuu2yKyECu/RzI=
`protect END_PROTECTED
