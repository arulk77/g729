`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
igLndomFzjGSwOgD0bmd1F1WFfJComUjay4Pw/HSOeXK2bKjpyPd0KOMGqAQaDol
/9ARKjVdQQFaAiE9oH3JJhQVxil+4RIlUaBoLaKU0PIm/fWILF13SIZvNgs40RUN
BRlW1Z+W1Z2GCNskTlp1EIpKbnQ4v3GtiYNTliYCvD6ggVvcAfzyB+mDc05fDWWI
zrYzq3kFGe8N3uuj8B85BvELzkflVK79rTYOEat1jbddEI75eKhAvQWURHDcf6h5
IXcsuaP7NSskUcwkewzBp3F4+Y4VYDAgX5C3nIqwQNZ/PI9T3TpiiXhFlzqecWUu
FGEBaTZLXVbM2rzP+SQhKYtCN7cLtr5B9z6yLFpd+pto1ReJTWDVzN/39tA+d9uJ
GzHv4TSSfpIuRyM4L4dmhWZjMpNOaNXYkYC15AuXy73TYrxWyivf+Gs7MdbCZh7B
xLwbgPAH7UpLxgIU5tCLMvd0auYuqbYdyVUSOoZdX4xtU5azJocnlF0Xtn/scMpK
0BcHEj7k8GRfabsdzfnX7DOSdsZppB9YreMfvhoFnIX1JMCjrYwBQjzmOzqtGRPt
/sB/z5wCB1D9WSA/DF1bNpOHcSpw3dkJvIoLDJ29zuiBStV6Z0heOD3pnhitQAHT
+gWw9XjAHQlvQwZpaKWv3d80iQlYG14P5Bdtmv+Ho9T4EOkq+kmIEz+PonhixG7x
52qCdxNswbOop9WpK4K38ZQzOFn26Mz806KUOA2HkYK4k48EfMegzJDY/+kEkft9
`protect END_PROTECTED
