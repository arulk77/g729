`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCMK/bE5pGCKnlOfsRxNCf/yb28T1oc1si1Fb1R1CdUR
OrpNA7cWPWVzhgngSAoBYxc/au7OAIkLgKT4H5tPPaBVSD7i6BNU/OHQCGMGGdyD
zpyf4ql0fTR4w07LlK4BpCfctbg/XhKnFNmn7GnzdYUx8Dz5joRzrSw6Pb+T3BH6
zCrylFFuMDH1S3YkySInjcvP1Nituak+C1M9P5uoweenrajCzdUmTwmXUg7azewr
SQOm62J06iGf08dyj+djCzQpvaDk/8DbAt3kntgiriV6yBHCGNtWsiFS0shXdIP5
NzuUmRcPvByAxJf62Xl3Rj0fx3F32NuRSuC6jNwfy+FLYRiVvnw0uzwC4Oi5mI1L
rkPHEbtGYFiygyilHxOZJORIotJn4KuF555mIOmVpDzxal+CoAvjaOqeY3JGcC2y
CdBEfR0GpE3EHsUreCnRQnCfXmI0D5r+pqU3gaSlMio8HJd4WiPXpCc2dWYu9T9p
i/OSzB7gR1ycNdSsXBcqDh28LpDlKR5ek+GhwXoD1RDEMtUGqJUJg/xluIr1ZMLv
XlCg0+huG7KJL3cagyanTdUYw4FwDqXyxX5u6vb+UCQZfmIAYH8WwzRFvnTBYV2U
b02nTV30TmYLmT+UR5hDVc8ySXejk1/afiXofmri4wtKIsDYkENLXpUjZkTY6Qzz
l8A3ryl9T/YsajiXVGnLT7HxU1XpALHOp+euLpfDh3mGE8uG97r+rgwuuQEwsllm
t5YogpZyHmAJcRd0eSis2Q6BYMRrFVGtmjLlMqAeJJPJ+g336u79JKsaEENlX/pV
Pi6pCFC4xa44uhF280MSviEtU00sRZv2W6waAVKK3ollj5d/E+K7av8JRx5rr804
0uX7PbQeQePV1PZCVd7+4vTlvYmDMEcvu9p6RzkWaEVHg85yrx6rNHUTnSqMB0rk
HVED7G7qqlBVW675MjE2updoetAc67gNQIWOfTdNKjjHsD8kjHWbYoKVLb00mVB7
Uc2wEnsnzvm1KK0VFbWtCIe8r2Wr1unIekj/k3suo7ogJEzVmsB9ZnurfU20iRov
2xC9XSHe22daGT/b5K5Fr9buW7upZbYNL4AcBIQJAVMHEuSC3Z0j4b+qeyrRacZy
YQJOaNndHlt5Ss3j5izr1t4+cO3e9rS9XyKiSpZcikj6iubxoSjm/FdDwkDsqAZB
n5gkMWSlrYqjJAAe1NyE6bLjaeus3xkaP2niY57LLqQlh/rz2OukyqyLjbxC8pLG
n6nfymNRRRcJUTxrniCPyoRVyqln75hF4aSFjy43i7RLCCTFDnfmW7MUnrsPWPBN
8jaqA+VsVUu9AlSFT5poKg==
`protect END_PROTECTED
