`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOlnm+V0OU86cu3lWv5j6Xn0eDVHYMMYdvfgN9h85nf1
Z3nulqMA27kkgE6BxjAqt/DTW2zeBhn4rQbfP7u3dOI7hmI/Xlo5i8I/+KmoDp05
Fux2MtRUIrhpbzAK+01PwMIsGGjWC30oIhIzLxUsievLFGtbgaJzhLR3rUj7qqZU
VTHuNOgRJuifWFTcdqGKDyNSjSwqzEYT6nG2z6AgAaGDmRLgkhroOxS36p7A3K0a
1NkW8JsZNvmQy8ITvCirAp3tsyGdkmc2tjQbJcvOt6NG6bFnBy5tDYWfPdKrkJD7
/Ac6tbPoXBMAOK7o0T0Fmi2mAgBc5Vq7I8R6D3RmPwKh4XCJa8jzt29IzL6lJFjv
whd0wrP6xQE0Wdc4iMkiNg==
`protect END_PROTECTED
