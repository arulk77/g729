`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOorua57fTvi7Lg/gQwV6WwUpHz5m4NTUjliemFOn17g
VeZArkuap6IAd8YcwQahPBhDE2gTlhJYc1qcLhwbkM7TJxOKrW1bKQ71HXyDae5c
wgMqKr9Nd/55vp9Tdx1YmykJnVFWe34D6JK6FwFo4h0toQdRuGVusMVsqn/ne81j
VZKlw0ymuNLW0rdxbo3c/ioxVXZGYQ45kuKSoL3F35c6KLZ2la6JlSNBMaxCM6zQ
AJPv5IUYHckoxTU1bgWEuMDBldFEyWK3dsGJNgc1oBjXQlF0FhW+0ei+Sj9YbeBk
TpzU2m5aV0hvQl2CMhtQZc71icRCl1Hl8weJ3JTNeMug49Aj2zNjf0AkA+0tbixw
Ofnw66BgvR/d1ZKxsnAC1hi2rH1WITHEqvfBvCcwSrJHLDdwkdb5iSez32hlzV9G
uxO5bwVEc+IN8wfECe47EfIA7vYPnL8j36nNdVfuiDNrEExqNrSvmdzCdJO3C+rN
S6cwtV7e3Na0pU/VUjptY9sgoWJT8KR681uWsjCBtxSMGRa3oE5O8heVmoicL8gw
`protect END_PROTECTED
