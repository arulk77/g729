`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEuOtihT7etdQy+95R424P5U++nrQAH//BNV6fC2cRvl
MFK9d797N4D+Ywu40CEkET0+l+zxlolibSDy5Pj4BIhZV7Og4O0FWIgHMiFfYvul
vvYezFajoniC7tKtwgyaGnqx2Zo/kxJrk5kzscIGXwx9MsrSDYi9SIfzf005uPkB
NWy1Sf2Ip6pLektSabWmporJ0dlxfJFVZtx0plPZEmWR96MlLBSfeCayp/M5Csvc
`protect END_PROTECTED
