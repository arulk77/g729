`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aRarnL6IosqTLHRKMuBJPzCgsk3KDcAdNOhWtV+VVRJK
WWiNSSRL/ox9HGhbVgYaUiAEuk9gUeTShAE7ti7xQaPeaexbDvxK9QZcJbgpkvAp
m+/2HGC3fI5L8SnGM8CQbB0A1DKvo44SYx48DgsKGLnWhTaUqxBuG6O8A1TKy2Nr
OmGck1KTPIdS3kprrYBUaBNZQ+/8seT+1rZDV4rO9yms7SEbRVZMIjG6UgdSxqLd
8dKEE2sstROcI/mRb9Q+s0Nd8GAbFGG9XYl45UtjdWynuKgUTJBcFrsKwkWQeVpd
Id86LyeKPO50K/b25TDSM2Y7yA5AWuhalBLxuAu0oMJOlk5tCbCHyRJ5Ux/BVNQP
tEcBXgnYbhlJqnQQr4+KwdFhpkTPMYSn0FLA+MeaPLAxoVi5QCw1U5kqROgKd2GA
luMmVosPTqlYrs3tNQDKoouRq4nfSAe5ojuNJFteRCUgzqV+uD815xHKkCp1sYdL
RZkrMhDmQCT3uVVU8CPHuTElLc7rfX5SuLhMb1Sm9lz5jVJ1i/XAKrXx0JNRy9ZG
kFrpLBbqvoSYhtfcLIhshT35E7iSMKLiiv/x+iOB5vs4opW2I0S8LbY/UxwxEOTn
OY65/QpXiwXPR5kN3RTgDg==
`protect END_PROTECTED
