`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNo5eTsfz7AIgPc/kBsPA5x+Ofqj5sLAWIe2RyLxrBAv
4Uy6wsZxBDj8DORyT1QEnX0iXD07uxwdSbsyLRS+DDpyonZ4n2e4Y2GMLaPmgwMg
pPnggUtVnxqPsRAAbo5ij6CdaKIqstOSM1RjwVUBo24mrIxwYNU+W8bUvnM+SMMb
rELLnqhsuAdxAKCci8XGNX2KRCjPVt3ahQMJjyZ67QmQ5UcFK2ymQ7irIfqKJEb4
`protect END_PROTECTED
