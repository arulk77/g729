`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLmaYvJ8epK9Bj3ndifbVUQMGDAU4YiAFOTcq+/cSfXd
8VTfTCckRCeb5jDI1HBGSeTp4u4v7Gw4K/jv4aTcgg16J4g0nBjsnD8ND7rdV6bT
A0i8x6EeDi0vJtPSRBerJG1zZwTyEe2DploJozfCTA/AoR2FPpYx/5Pd/EAVrckm
E0Xti5pWCUD4PAIYq8+AptzOM2Z5GyaJZfRh0a0B40TQKU/HL1BbzLwU/HkDYWVY
Z/47FZov/aZUN97moh1cR3j9ukayIC5PCJV8680mUuLv37SPbYFfMJnFt+cj9Lbl
THnHoRrizelKDC57JIRI26noVOrNXLQpM2LuOdX5mxZqgb6nbvjSBXkDkc5IeMtd
nt1gKtE7e75S0/O3/e3Z4UoTXJDR3BxGTFXm4PS/lfBk4Yb76e8/cKtgQJGFn1pI
2JPPo7oq2sbvviR6N7yqwXThXePJLQx386L3nil8sVFWl5C9iDkc2ruP/1hmybAz
0k06/qygi5ffH1EJdY7HQylvBl+EKZwajY10L5BfCwNhqGm4uBTAs18dKWbJObPo
ySVBZf5NFHjqgL3W84Ior3kK6FzBarBdDfLYrvQDCzrrl+a91B1pJgHsyZsSspuZ
JpzH9BjoP0psS0TtgP4jfrEEF3clFEVbHXXaA6TgjrQTIQcEFAbldyzjxSpek2ty
d2V1CXqbyyMXbofsc6KgswNnpjJgg3FxXxgrgakhKGmV4axF2eb1V7IsyBG7N6M4
8TFzdrBoTm2eWw4nJm894dVS5CDd+hTslAmtHvMTKkRcTPolynR8CMg8ex8SoEOv
nilnbn9uxdQRwOkAaht6c9kPtOJpLjW2H1CDabuSS2EUmCQEckEYLL+Y8Vy6BrZo
Qsddx7YzLX6Z8CZeomoGf5CCPboyl9HtBzg+ahmwIU5juZXlrr0Pq/OZWEyt7QOu
KbUp/rcj6wFIob/n6DqIAqXv/9NioV8+yQLPr/7lb7A06RV3xsjHnwe3uZrpNlkh
rhW/zTAO8d3NZq5kRqs9cdzAE1NcjsxVurcsl9zPQYss7zwPemUfUCk416gbGxn3
yK/gjSYYNNK/V7Kx3ioDftT07QTZ1qZsAb5rshkw51CTo7WP2hTci+HsBMue2dv5
0N1lPDfJKUKREAjIGcnVUvDJyUoOudOo9FRFrK3gf8dKplznAIKPWB2Zw0x8EoGz
c6Mq+AxSiPHWVhEZppMe996981aWmLJTjyP0GPF4aGyBTKBiiIa4LdkphqZGFOgS
4T/ybyle7eaTaHixS1DcQpapB8G4TdLMxhsvoeFdnB2i/YakEaNlZUc5K3Fjb+Cl
rsJ5FNtMT0w2R2YjuSJmzQIUhERwMQpXC9VZFuCObaNpYiF4iHqw/HShLPYe0quP
MnVlgnJfIW4MbBXl70LS3d0rRzgrk+TjZUmeB9zv/ndSNfXowsx0dwhzPJwHGfSH
U0uMwIA33j0q1D6HlPuIEdPncbmkMKUz8pJyM/DH9b38uu/WfmIB21upI0fMcx5j
3zJXvZnFuz9FCKIZDCSKE/glximD4SlMOxfcrbz0YtJJl3YtISCsD6FM0c8xyNy2
9mXd1mjbZWLu/oWqfuG89DJyrSgirl/l7qWifP9XyBI65X++EO0AihqIT4utNxr7
CBJKlO4Vel3Ms3o2u5sUQFRCkTckkZcemlQqtXPU7vgayG0pK0pZR8zrsmFVCeex
EUjIVH82ib1K03K5xqZUj8rsvT3ortebjeHbnFLMX1NGwyVXcH74v8VipnDa2yYp
SV3V7/qlmnYjzEf5Vb/hPNINbsNCmX6khNjl2xYUGTKpX5ZtgtAPZkMXJPZglX3h
2XidTYlT4FqNcZ+x0Jf8tSetmUqg3/7I/CxJTXsmUtZaOj09mpJX/WFwjDu568se
ag6WKLe9MEyASTIDRKF2lBbl1YHraXOK/VybubpW3hYaMAvuIvHewkI8NAQvINkB
Mo8YTMlikqvzTAEx0WJqSjrrlAcOnoq9sADTBdNLIgbcq5WKX7h615FQrWKO2UsS
16BsnIR2G+5IZV8GbOMpwLQg+PuLSdxMFZ7IzeM5RF8c/oiw/lcJFFAgkxzDmNZa
3lhx2YwMaWSS3sewa8vvrBze6JBDbT5zo2FB+gGDmPHLZPY4CuJzsZRGZTy+f51F
MNJpG741gwgQeWGyMhkjKrsx/DG2UMz97Eq9q+PHMtbk7kddmDauImSAkgu/gAVD
r8nlqP5R+UM+NBNUdpb5fRGlW8Y6VZqzraaT22s2rj5Tr34UT27uQFA9Jvbd4pJF
NbTf4p8Gg75zJ3jgU5L7R4OmQK9lt18I0SE8ZjWs4YJRgpWsL9V5KlVLFSY2KHP1
IN64j8aFL0Loz9FiCG9KQEnhA/nu0RsgSYdTzBzpWmw8/tPzZMiSW2s7IVcaZB4j
iwHB1d/5/XfA0eUToJmo8f2G5sHXEuggiyBP8c1x1YzMZlYvwoSglXExlU2xIKj4
uX5O5TyrZiaRtpMb543Bb51S60qgE6KPsJQE0sXrJTyv6UFcTQ1By8Dxw2GyH+OM
wM0MTwgLZNHP7TmYmvICgnHPWW++4FVETNOUs/6kn/xwSQ92iPswWa99cT7VXnW+
RxYzqqZTJQPchL/QWX7slc98RlRFQ+ohafFsYd92IzacicbzzTzxWyX9lOO1qdY+
yvMBePAo+YhyGiIyzrgRcwiRVp/lgk9m1DKDekRo6ST4g9QRpcTesk6muQa+GuZb
+dfGtcCvA+YtVPNrqEeDr7/VfQ0n9ZA/BVEoVOlwLWaeU31Zy2THuvbaA8+QrDDU
VYJZQ1bNJYW6dX7p6HWEvh0D3wLRaF37xcmKPQNY4tVPUWchsRn8eIHaszoqweAU
8fvzKDakFckpw9yK7V+puF7LM6y+jh2YukheOOy7Q49/eCB9M5w9wwV1FfkzZLKr
nNCepm7Ilin5ZvYThvz1rn+RwWOvRaC0Ln0hPKH3mLK7mkD5K0nMB6cWP7g3mrkq
9Ty747MPgvFiylojYI9GdHTqNgFoD/qgquj1vXUOpkGQAze2gcAcv40ZSOVdSjc+
nAd3gInNjVbBOhG28cIjOuAPeo1GimQbXOmRP5MzUGVTY6xa9pKcNhchT64YGJ5F
ycPg8HJ6sjDURkV6tmZg33JFu7ESW0b+1siOGjjDcMxru8JDSycZ/qv6m6l3Q14O
fWNGqoqrOI0HoAKP3u+v667/x62NWG857kuUU4fnMRlZAnvFF0BiR7tvMYnPo67x
LYIa54rJh3/ZPiL5DawG6ial0OBI3x5/vlAE1IAobIzVusPQUju0bfmg3QDSBV+Q
OYNbIwsTgT8haDfh3SC7ZUOCWqEXMWjFZKRPhddQUlucI6fxj67D/tqoaya0az7H
8+Ms0ckQ+p/2Do2Nb9DHtXC/D+J0vauxg5PckYZMdwcI+5EadOolMrfPl7Skx5fc
IN8F60PulJ5V0bb3qXiwAet8MTiDvM5DGdHuOccuroGEJxyPlskGax34E3rIstZs
H3X0IU0Og1b0uvL3iQT+lMl88XfvELA8JNwgsVt4Nlf51FwSNgmUK4EhaES0ENy+
aB1P9ZHMwKy2kbjpIMVRXj9KpTLS5xuYWHgFibwf7XrrZKf5jUerbs6A3sPWBOem
/y/6w40ibFETWrsThV8uw6LhYVuvTpz47kS/0n8UBW3fkWoS3Kb96rbZVGRRRT93
LXBgQt3HdOTP4FaG4KVJW5ryt3KCa4eXn2FUVyeFnwYhgM2NDx7a3K9xQRus5Llf
aNKWWFzpxnXf5eTDNV1JrwIhfq6WzSVVaxOgJ8FlyKlEBc0OxjZOhDev9tvvVNP9
sSKNFyKpPURBz0y4xmz70GchKAw+pVzaw3dnFyHm1FVP0R9ysVYAW4dESMfILkAr
Ec3BaJW5cyyh8HyvSROxbmTvyeT/6eRAZveBmdRisKtI4Ub7PU7OPjy434jwTtr5
rhlRFLGHnGM07sTntQweB3RVCL3t5eVMqDFk/3NXJAzBCtA9SGmxtfLvLfOxjRHv
SSeq6i9r0U4lxLrzGHgCFJtJM8OBqKAQj2MVldTNPLEZ86qrBAcqKl1daTq3A/Mn
SeYdXOXYxUH1M0WED2UJ9/C4gSkkjcm0WE6xYQC/1rhifFkeZRq00+pqU1C9tFIO
C1D99X+q9jYAGrAL4jQvfusTBvQCkzDUkt7Vbw+0wPAKwCExv1RkILMBkg66FasG
1hpPtLJA3d3f+fd0miGIykpqgwrOZtkXi88lhyrJ3cYtFVggkmLCnRvDjshGo34W
Hz8q3MVYLueqONY/p1FvW2wRPNNdcR8IYqdkvwfjwcrCLy8tpc8jg2YUJhKXqaTu
cZAr2HourijD5dmqPyi5CHTwWrRKAyXeIbswnrPs1ILhPzwk36NbZm3/CuCM+PwJ
xtHPhCBx32G0N+DpCaIVb8BeGxKYJpn87pBqbOynQmWaYNNfo54X9iZJiWxyD1b7
ohCrm6QJDM2vUU7v6gIGfY6X5On/BfanhM6UCdLfpVQy+04HiilLp/ctauDIdFfQ
NMnDxiCHcqbWwm5JlEY0uzjtDDr/wrA5JsxdI3xES6222VlJLy4H55iMkjg2jreB
hznZAp4sziQhm2pPv+8/NB4xFGb0ZyJtBFImqoBZP5zLtb24EC1No0OxhSZ3tmab
bkcsBHumY4wgEwlvgv4ZQ6eaSYPXfMt59P92j21Vp7X7DXm2T5Nx+hYyv4kznlM8
w+DCGuB/0kQ+Hh+nSbl1HzoZhApsPu7od9++gHLKdTAAdon5GuciUhxsyS1UDA/j
qTV4ApIUv1/b0jdQU/Izc+xFqmqjA0QBP8XUPSVqUDCU/+pLYvqTEzXg3uvgYJxk
e9zIzXG2kgwKBhYzTXXFU+P/EzhFZxjhx8aWCq6ZEdXmEaWPYljO05CHPpBiydW6
Dn5sGtyPpPqgfThd1X8Z0QDwYy8S+MZOJD8zWPbptYf72f3IuN/mUIkM8DG6/D7M
jRGK1XekRFM+xEwJgAsiJhk9yF/WPq1N4Yg0O8LS8tJQ2n4TIDEsgNW1XpIeA5LI
nJtzHQGO/rZ9Bre9W8jmtSl6KHQoTXDCS3fG8sAg7YO+TdaY/BKdaxB2la8cf6kl
+9lVV/plj2XZZMJuRbjMhhYAa2O1ODiP678RR2HIRBmD+IRkteTPzrYkQYJiRZkc
Bmbu/sHw4NisZeIvQ+A4wxbmIzUB6ETtKmro1z/+xEjh0gvuPRkiR/u+7V9Bf04d
5KdMX+1CVATiaJiQ2oOCzwUoiDTFsxuAi0Boy5MvvafgzbYdHoeosi7i0EmUrvzn
VFFc4PljCOtnywlm2baH+YGPdhCQB+FsdQeCrjbbYvO8dvqR5BEqjXR5XWs0QEE+
VeGH++ftBaxWbSnEEAn+Dr9JXQ7Km1oToh/jb6ECG2AGJcqJC1CZkRF6Jz5/iPTs
t6SQur3UMVqMGUYxW9bqjX0xBjJ3+g4gofVNeBDwFgzWpIyn3cvG6w0cuWNVbMgy
FuJhyoxltoxbd0DyZe2s1a4o0b9/xKHRZdR9iz4XIoK72uQl0lGGOVuqF0dqfowa
qT7ccB50bmPFlKbHfFueL47uLvIPleI9uuBMkryLvJfLvnGEin3iaEa/YUXC+Zaa
JYzN+Sq5d8+r2BMx/0BTcBN5kFM4P4nhai6ECslsiCL5FHqwkenaMhLmErlIHXIc
EcLfrZVNFJ0egWD6rIX7AMceiDEVOq8oSFfKWlXGQ2JjXE8M5rTNhxr9MqZLvcez
0uRUvp1RQdrbT8Doergojejse+guA98VSwlD8QYFjq8nd8CT9GCTcdGXU67U/ZtO
5cfhtuL0IO7dQ0CrNjf3bP13RCjfnOi0zxGGu1o4TKVmOXPCzNVxGegfEOil8zI9
9+Y91mw04zvXenFb3OPpD7qU05LxWLG5VIQQqzrb6kQRi61kCSBqy83sVZxsoanr
lZsEDTvxow2iKZsFvnbCR5G0ZLF9dAd6HE7z16h+tNu/w/1qPURlQUivHSChWH3F
+o1A28tQ5pl3RiejruTIqSmE+tMWdYtLW0yO3i+9Pch964KLfiRxK6AmH/3YXwU2
5ckyxi86tVEUJhagrAtehPWYsUfB2jty1aKl8hMz/6DYIUePt7MZZGj13j0aA9V/
d91yJhZh7RGJuNiCTMpeA9bgLxwHwUdqAi1cTuLIU5qqu+eODMo4Xa4pj1jwtwyr
o9W/rxJg1erf5L+7Czfy3t1QWmE9DuxWJi7XJg8yWbC1WItNRGtrflwaarJQ9hUb
8EcOzR+eVIMYkMnGMKhC/50Bm3Y3ZFmy7W2b/ve+c2iNQPPP4AmKGA3ezQNNUdi3
m528QjBxIk67lYv52yEwPnSm1U8jwYbTjVLV17mllup0pOusk1o8Y+LTcnJpf8Ph
+/k7VoYEs17ChC0fGIqDDpoVsfRlJiq/KVinIywEcSWyYl70DXWRsObW1QPAsHtL
K3oURLwUyPsLYaJzljlW3E7SOi9ZR1Zh1HhPHGO7m5T0O9pqeFjiThnPpyc+8LHh
whuCU72pxLTfU1i3r5dq+UOaSaElOLZKhkaXb4RNfvNQmzFn5m9IwxSbeMmhmf53
vuWSYTE863zl6wTfwAvi/FLdX9fRfEQevmhiph7h6srFC9aOYDgAMqWo5oGI0t5z
tPEKZsNhA4orVwX7guaJyY7AFbh3Pg7VgUXepj5bQxmyShk3Dq521faZclNTK8QU
baYfx47xIqnHmEqI9ufafmuUhPananSMD5BOq+VcpnHV8V5P/AuVjeTsEUfpvnVy
OX+JjK513w1iZ2apR2MAL35zOET751fos8iJDodo94/WK+PZrLmckJ0zQNLOzAmL
OfZStk6HqIA/cTHDEgMT8DdzFGs+ONKLvaNd8f5UaQAnSkqW9TZrLbw762mOa1c7
p9OacdmTZFBb9u3gTRmhbj5dRX5TyNX3+mA7yojGV1R0ULCHcOxHilXu2X24WZbU
E5HKy1Qb1nIU7o7dgS1pSfzM8yD5KxqJyPO4XY/RFTYnCnJmqBRMeCKPQB0d07S4
K7qVS1k9LIxcnouNlKVAfsOgDe42YgXR4LVyZIHNu9g+rXfU5RySFUWWZf49nIc5
QO9hq1nrL4M8hHoZ9ZF0r5kWeHPAOGccSRV4uBAdk1W78EeceJjmcoKfgCMu7Ng/
z8zvO9g/RZ0++jVPoe0Takqw4mPvXFYF9OVZ7YV+zuOzit4lalN2P/Dd6vLJjQbN
YALUjga3klByQa3iWODD3arBnfsJBuW0S66uvPjlHtVx7ohCMhan1n9A9VKyAcdI
nNRogQ1omJIJ+gfDeUjCMg53eLGJjsfMR+ZDcYFbDmLzqBkDxMDKxGXRUoStotuo
nnHm8vFxIqBT4jisgsq5xoH6MJO+sewQDUe5Rr4vZ/0TwKboGMZeK7jljnmpjWxM
MbQkMd7EZdEiecVdQWdGtZ796l/6UN8ozmV6Zrb3RZvrLL/cOK38XPtukwSoj4on
pHM3ZUP4Kon44WzvHSsN1ipokrb1CAvRu/uADJXThjMS7uXX1Jto1ERN+++PgtBI
XFjjNcPf4zpJyvG0elXtC8bTCa+TmsCGcGrmw8VlNsx1dhaZRybljcJwSbpcALpf
XD8oieFVeJtIwDj4dF6KOwd0A8UVRQDgBJCtodzGD0oZMpTT1CHbCcZomDxT+PUV
s/miwrH4wIkFOYRkf/vmLm7pxtllYQztkWHDHRZiIl84Glqa1AqJeb2raUdGxwac
7CjcIqiDxvyh3eRA+WDOGJJ+sLXpXYesawD3lEWJRi6WKXoV2qN/3xLWY4vWHy0b
Qw+TCrL5R/7dX8cOYpxQAzajDZ8dOxpGLpF1VW23EvcKDsXXW+0sxYvQXsHxC+iV
DrNI+Wkw7cEtXk5BFHEFWWvl8aTVoQ9Xwu32FeNZ6mUnI77T0zSEDO4Nehvf2YaA
YYh3LhwoyBN8w5+GGsNLqdKK5WmsPsDR+quDIl6OXG89nhox3iGNO6ZvnNb8OBcE
6MclMZQhyVYAF2y+CVWmjzZtircQEsHyoLAVyoMkno0oIN8Z6bW0zNA9v4umGPoo
btbpVaHYlUtpyuY5Fa688koGuCW0J1p4wcZbtLAxWAZ9QSXaj3fmWMn4lamzU6lf
GKyAy13qyrIRpcubZRf6SEWbvlZyowX3K9CBP+z2z8k98oAlviKNZ7jKvArXOURf
BD4j7u8m2OdU6yrVX8IW0FHX7WicgXnv9uDmiQ9rMQxnVB8CIHnGvwjQKHTSj/K0
PKRJXImncbEcU9zuIgu7FgYIUHVr9w0qOyi1X2SVdt4XFRKsojVfy/omLWd0BfCz
vGH59ilTRXG00iScPuQVBGv19tL88rX55ISXQeWxM3weRcwYcZSP0o+24WoMMXH7
7c0wFhdJrcwRrw/gnRmqYJHZ43jm/0jtr7g5FvXxlq9p+Ui5Rwc20ZQLfur2Y70R
5mGsoA6zVHjA0HBrqqTfjCZHE734JxZq7cyaVq20SIsJffUAWOGvXjNmwQMF0SoY
86LXd9SAR/17gQuhNmALhi7il0X0x/fX584/X1U1Xk8gR5X6UJAkQ6RM91fekSOZ
xNS+mOse0I4U8dmDqg3A4bLsGNe+YTcTob1u1lE83+R8Tpgq1HNB0WRKabsLkKGA
LHu/q4f70ycarFJ9T8o3qxcPouwNSdgdFkOhb/W8GYVUyDBMz9CcYLiYKOyTus5J
qfcqQcr0Lb3S3w1IZO0FyxcMZ+SyqsZ5lLHrIjeVnQbbtbpHDPvcU8trK2ycYjP8
j/L2ynkkYNUt5du8NJlR8V7/YhZfBHafarYiHfXq59bHkeQroyN9F0qbSZQh9I40
WVY0eEPJv/U+iQzP2mJROlrFw0Rba1UIR/rKKTvOi4FuEsrAycpX64hGLWetS+De
mvJ/I4s6xwShCcdVkjKGCApgNn1KLVEtwa2kaevY806iY96BJ/rcvW+ER8z+98Uj
8kl173e7bU51q24PFw/3f/uabPbyEVuvynoblIfQ2yn7PDj7hX6o6EX2m2cLqcZa
tuYupUDf4IuoKs+eCMk+wPcuHbUFWv5BZYaadFXvlRHnzZ9nEOEIwuX0kGRkJp4Z
2rS6wlxOzj0eZQiYRm5/AN3phSvOFhF5R4EN0VKAW8TUlEJ+bpF/pjaLG+ozP/5d
nfseNesegCggIabLGWdXV+vEPQj8MWP3HDJg8jVj+U6I1pPD5eg71R5hTFsAQpqc
GJ40loZ62HKLJNCZHkqyH6pUiOH6FEmhupnGwWApIfPqppoka3Wc0BPGOBUSoRRG
SO/Xu7Ycmk17Rrd1Wz0X6yocMtxLNQv9+XuWflm30Dhx4EmMBWAUnWk3+BSBWRJt
EppkweoVVlIdzZqzucjGXyrRKnCVpy2x3+7gK2b/k7yKIQIcFS59RXgcz/3gFVCX
edIjmH3JDvBzEGOrtjNt8sjNCF8KdEzSi6Tq5RDq6Ylf8AkVaryQisOXybBPr7eG
O6uj2FWZBGoTOCt4vkmthTiVICnveK0R/eRspTq1DLWqV+R6Oo3YBn01Hllktccu
iZlFRrzA6AecXRPHnZNn6JeRgZLWS6pLIu98Hf02O5mt3I4OhC9q8JIGIyGsxz3l
KHjWpPXQ1iQb1LD+um9UyTctqm8sfSn/UWWH51F+H1JLEwM94v4KY5pHT9FW0ekb
zN9876r5IhXJBdXKb710+nisgemtKHktTB60sX7N7KolsRlYg9nxMMPIvKstkzJY
PRT4kFReWdsj4/xIjswkR9bY/kVrfHRGSZjVL739r5HHxxhB79iWxmoGPw2jBzkn
YaGzcO2AFKpD32MHghuAdyW9Q5eAgtlkjhvqjRGrwE7dmujpBtenqXnbDeCzrH89
nQar1IyUsMUqdF0thxZQ3CnJbabhyPyiPoSlTnVL5TPGfmeC/NioavD78oPUwM9d
KJEI/sAT2elCtlvQhoKw42KUOf4PHfug3q2ZS6ID/3dH7gRU2Fy++QhRuLfGH3lw
iQ4X74Ei/+QodAgN1A3YiJs/DpQE+Pwjr3Iyktw4zTGhL8WxOFCsJ/jMk/XvCGmz
SuMKMmOF+Q+2dnheoqYIhk0cCR4j4NGzoFNoadi+KUAHTUWaRCM4Xbj4G3eUlZCB
onzqgE/CUCWz62EmoRaMJK6ParFRGO9Fh5RrbcZxUMWzbl95kz63Bve273fnDAsF
GKohPoD2bN4+QLdqrT+BfPtWNKKB+u0D9zLgyut2Edr0TM/F/z8AMAJocaEo8d8S
POGvVhK3IbBGxgbhuZPWpw8huVc0RoOrIGJ89rZoRbZVb/M6oKjsF9HB7Pbbm4U3
xQtWq6MRKj/Z2IgZZhQnfymf/vJ0cUvLREvQ4mbXy00MKI14zDFHsU7ckmH/zGTr
P20huG1YhktVFgOSF0xiN6gzReqa4+Bzwe1REHhm8WzPfZKrDaddzU/oMxe2E8MH
NdNtevkBoHlZzNV00l8Q+kdCCMvkFhUZkD6SCxl+z1YGMNI4sv65zlBZvUjRzKj2
b1eS4UJALw9tjv5hfLbXeOzOWUhdkC0nUwW8e+EbacoOxPfKqKzFVJl+RTdE5CEW
VHbiUbNkmM8491SO7drqBW9/9hjZiUPFjnqK1RDQvUh7hXAmtxAvKtDjlDFW51/t
7dRb9do/OutH9N/PMrMkFDvk/aGauIuiq2VS1QbLSME5vD7YpFGIpdrkOQ8ZYMoZ
Uep1W8g6a/clhnkyX7Q2bdZwkmBUEiTsIHEP/KTYqgkeklmCuEKNSFmG6kKd5ZiY
wQQpl4veeMtcXwtAwVH1+JMqJnRly7Q6kn3g32sWUQ37iKPyR7lIsq7eY2fBLMP3
oDR4jHH/04u8Asi5AE2AdYmQT9cK3WNTj99Q/QopGx9ealUxhoG2JNiSWqn8Vk6/
6V3wjVe+OQ9adAFjdLkFWcjFoPLDU20x5WHVLi16bbpn95Fi2q+8SChLsJqsQiut
ttacXtNpttWqZNRe+gSuocai8GSZT0WVKHUjEaXjp5IIeuA6MBVIwBFLJkfdqrxn
pBSG1PNHR7z/Q1k95eR69s1r00rGr/Riy7ZACBbvSexMKT0g9LSTP6GYLeSEj7v+
rDQgZrZ1y7FuGmhNw3oOeH1Npuj8lDhdaJ+EVV506kH35d5hnjJfwOzyWGNzEnKK
YzaulBCrZi2cdT3OGNTlJdEIh+WmpGt7GPNMZEerpl1BRRT1iWa+uCBz+o1QZbHR
aHroo6oSnEi8G+CKkhj481NmppTrmyONBkx6sL8xFTIW6XHEnMBZ35rTwOWUlQm+
RX4CUQcRi4meu8PPYJ0+CS1QffsInNWmYWrx0W+b/cGGZxGwdShCWwk9PbSU8/XX
W1/lSgZNYu1FjD6BILsydTuGtIBnZ+Z7PnAWEDnyVO/cR3Pho1siBQfDPQyrcpTM
z81FypzwCpeXLbnpQjeMlBI5yfgoyUHeGSacJ2r1s12PAr25edEDEAgjzLgRlDZ3
SLnmC0As0mTfKTbSq7mPahKi902nJ9vP4CJy8z2BbCysVK64GhJ/hkS5H/ww4V1N
wHQQuwfhCCNRF+/N2RHtM/5jNfCZwCYWHNqr+YTGE5Cc+faaIt3mfoDVqPjrmTeL
acGtqSb1yg2Omd49qB+10L99+i4PmapntvXX16vsq05NgP0TZeJ6zrbzde0A961N
qZHCaH1gnfENjadqawcC7Avm93m63V1JjiP4ViKeEAicTm/PlO0R+V2DaFkPSrke
YI7nCULydXYD6+V0z4mEyBR229bCWM+z5FZGXhMazlpjFukXwrkej1kYt6AnU+y2
ISaHNzMsuqgHZBp/NEWmQhM+THWP/qw2ACqWRcJJDqV0DUPQ8o3qXQj8D4xJd2qd
393A/sIVdT0oGiMY5589S9eg4BZSXVA0KeHocwhnz+Z43dCsFEEML0mlsI2kAlim
OeNJMbTOFH4bqxpY2ifv6o7SBapFm28KdDDpE6A+fTzuGXe9pxBwjtABol+EFl3P
ScRkosfZZnMFK8zMCRTZ/RzdBrKQ6P+B3k7uWjUnMuZ3pHogoWn0F/R7KNowg3ZH
4N/smX35PSgTZMaW5AdgqRP4g/Q41k91qWY2IvBep3F070fU0AJg0uYvmeNaLiiO
//cQpdZx2NVQtjUz6xtFYgS8+gNUg1zjG6HQ5RGQz6uaoBOjYJAUzzjyrKv3LZMy
gkCklAM+fEqBPb8wtGltqO5dG1f1FqEI9nrHJHpnnPRy9Fs9CoGgetpkQ/6FzQ5s
k81gzzMetaDntwUoNl4PcfzWp7x2yrax2D4Gxj3kn3NyfwJCg2EhsaonOUoukaF9
3cAL/1mvC2ziY0BYtXPv2Zm6fXSDjq7zDq+SNNsalXguHX/caaO/s364dUN66dmt
xw5IgSqDdmkwPgTDHbGhYLDjge9ogr1VCrvtcWnxhd0/OaUpYqNHW07wqEWAQbcg
Im1JmAiK4gZApLAZ5KUjH4r9VafhZF0PDws7cK1sN9UNHud2ScHVTewmu/7Ek5bu
2srTeO6BbVg+62NTwho5UKDN3jPcFMlSZmlI2MdeGBEcpUmHi1FyFdVvF0Wrf5Lf
yIx6YvFpONRHdKBk8KYk04p9At76Ed0r7KsjgqICOCfhvG2x6oCne46tpgvGeKHK
+RA9BVHp4X7peuRrl1Jy9o9g6S6pOhQzUFK0Daa1v9RG5Gb+HtH7bZpgDbFAi2EZ
HMoTresk7ZWnUFPFp5U+ODT6P9Ay2GHA/kKjDMsob3HvNquL25CT4Rebe/abjcxy
2a2xlzfi9dG5ffuMueeNxucoseX7nrDpdSqHkrQAgExg3qkHIpk8dhCkHiqFUs3I
PdDkQ33lh84D4p/gWQz4q1Z6HoZ0KU9ORypIlbUXjvjczTRUHD/N0YvXb2kAwvjh
ep5/D4eJTQODBGMS8cqVggn3KCNG+R842sfTfYUaguP0rjRzUZysiEWuZJ2mI4xC
YV2AZAPdILB+8oLoAkhrOq+lquHpIlNh1gCJ6zLIz93FMiX6DdzXldLxqzx9k4Mk
i5WB8MrMZ6TitujkceJoQvbeS8XJhLyrT88GxmYY1jM4W0nH6VV92ofKf8Fb1959
6jU6ZWFTPKzKLI8wiHtrQdKflAL/uQtWT973x624NqS9SmHfIuE1yBizEo5svgpK
KzcdrIwpb5Cd64qt8XBZuZEtdF0pcGGpYQGDxrjTbvEUXX44xe8ixsEmr/0MLSs9
T02BE4lB+1Smqy2jWq0b6fs1u4JhWK8PG8iB9fP4r3vwMtpBe7oXXIfgEinek2iV
5n1JvQGahLjxjsF1lEDFtqVuYLGigNAK5W5G4b0vgOETGHbEhkDgrHwCsu3hpunR
cCmmLyHWAaXJXSyH4J1CZs/5P3qdxQfXe1QjKO/yfpOF3BptEVgqH69B0UiJ4tic
ZfMCZa6MpuDIU/QT3NH+hoggs5gioC9p1XPUCbOA3sqEQ4ixbZauDWE1WFe0fmf6
fkwZAfi5MUkf4CH7ViJPPXSdjTYeiTrfu3QdiWnGsbFnOK+2KV79SVZ+Bs1TeeYC
EgX4zqT3KG0g2/Y7RyxtMUbrfJ/Bb4XSosCizp7XuVqNG3bAZc3wnlbG9E5JD3mR
6M2fzilBMsNWQZpr68dTADA7AZryU5FYuYenpbVD7/nCIQQanqBXBU5jeU+Rt+32
Qxy0z1C4NSmvmAvDimY3Ok4GbkkcyI1wUP/1DTlc9CVOQopuTELWleCvoRbdhmfs
mPj5yzWzvri8OXfGtUmKOI7gnXV0uCDk+MbpLXXzJoCM9/JtBkBwvOgFLQoS4sRv
iuInVJPBkC1I7Uj7h+7V3oxt7DUw5vVomrG8XeyrYKFqoCaa8EmVic2XpZmx4LiF
1KLSO4jsDZTGbrD52SCciN4gMq2VGUMQK5rK4eQtVfwGoLaf1G3/DKO6qDK0AwJz
tddOPdxNzoX6lT9HzvFLXlEiRQVS64qL8ttkqsZBS543EY1M30r5r9727HxZGLXj
X1AYT+IKGxkZpEMV8u4+Clrj84VZBEcNqFSlM83pP0sn81jBkn3xepKj77m7RPis
f6Sc63z6EXB1/4dLriAOQ+ociVaWCOrO8pK210T9hl9Dqk4vytyZ5To3x9PGIiVE
m52OxGU88q0eTuL042yT0xeS23JcDWsBALAP/zNe1ZOHf26khzgUyHXhgsWCZzON
/rVTqyEqe2qFRYBctfRxO9xEAs/D7U5GhJtyxq2MkeWVOAzCVwv3CqdS+jkEGKmY
xzBIppvEtSZwY+PYhrRCVVetu/fxDZ6++S6Zyjns7tqe32kC0QRDUbaxRlzdI5fF
WcujOQ7uHj7lDnttSuqcjJheW2Va+Ru4b7tjXr/rKRqhpQAVh2eh4NlDU1lGTvL5
itlMUAMdfgPKvlYSxq7b+3PLn8beyRWRwCq8wPfUyWDT2d8De/34uHCCSI52hjs8
DjXlVc72U7LsvuXUxOsWWcV3V1USYn2WwE4hq8Po5zmUyHHcKdYRN0VosdWVwdWi
b6WOKvQyOe/eBVfjZWkGHoeA6H+C0oTQDFWttKcwJvzk/mOyd5cjRbKB0BtuVtu4
3eg31zeT8JSp2sXZKdmjLBsjQfmEVD1hZ2xKGVU0F6aMBQQTmyDw2s8N4IUb1LtS
Fw92T+EHqzlPORNCAtVGcZMITVH3b6+K7ySLxwpDZyEEzpc9Fd6icWV0i9SXaC+a
0SFcq4hwZIzvAx1P7m9fGQq0a93c5jeAXqDoZwRMz8HHwOhknGnXf4u/42YZNlXh
DFoCTDDjka2OGA9w+FdGoAehnHirknBj6NwdnXu+oZi/t2c7AFtdFW6/a7yn6YkZ
uS9LBew4AxWIs8hCNT2W13NZ0nOeneNNZZpFXITk9W6IRmc9OY1UmCfrKs0vV9/v
BjQmBFVBSJRL4fR3vO3KUw8ea9daxOJOpP9y2Mo/Y5Vcj5zILI+kyabf9Vh+nMXW
4Rbw3XPmENl97YLtYKmIx28gv52WFqn+ZlJELw/Vxn/TJGpLbvxGnx9gYD+ediri
mcS0kSgiV9grZjwCyGGLIU+regudxu7UeE0LAhlQQfWSklDkEfzOWIUwHab8DaIK
DS0Lw5abXjywN14Waj3F//oD8VouSmo9eHufOBAs+RGN9EKjzxqm+Ma+Jg0I9gzB
eS4sSqsNW/f8EivydZ4eaiNigKTpA/RSKiL1iazrkImJU9YNO7Fod2tAq/5qG/rK
JvtDF+TI/uzaamv7IjkcIKADpCDnS5EWBIs6nhmXsYQal+bxCyJYXLiW/s8aqHem
29JsckYyjw1Bhk2YBQUGck+B/w1qbXQAKnUpzk+Cs3ZSazGlJX81MZXqf7ynRFdc
PnjPCsAekbNToYTyBCgKSYWlssUVmXBJJh/Z2Eb2Xd8KA1OI+HFa7oI6DIHqlkUa
cbK8m/Bc2kbMByBBmHt3Lon7KPs2iwWzZ+a8VdqTvDhndFt5HPv5XTvyNOvLrZcM
JivrJUzhHcJbenwOyQN01cOHMQ7ciUVjhaUIsKJQyzuWtMHuigoMt7c66Q8Z5YG7
B/Bpr1txPQuYqj1Iiwi90vkDbqKwJxK5uuMtAAbVic5t7iUFC4aU7UK1Q6GehBuU
FT8hJRccP49gMfEQmCCy+8bo2pUDdAdst6moQfdIRGaUVtnnPUAgvFKR8wBppTE2
gqi3MDRZlKjcGVyD+xHyGbT0mySNfgNuq/6n4LGOdUXFwRhOSAK/ayKvMjIq3Wng
0ZLwl0Cd0nePBe748MHAi3FUAlJfLPJDWx4mZC32LqaVMamH66YKsriVt4690NCS
djdYph75yUOB6819zepHI6L336eafFaAdD9CBZjfXUsTZ8el6ftiESqbGlmeXydK
CYVfc9V5EkmZIilHVscZO2yTDBHnGv/5vcLPefF6ABrWifzh+LAxW68c054VPqHd
FACz3e6UzNj+NJU+8fesPukswlOBoAIRU7hPk7z5gigVn/dcn2pHw8Y0f8gQNfc0
e81luMmIaeEdi8Jt3/nw2kbJ19zqnpNPI6Mpa517ztCc3uRvlEKGZ14UqiLCPUbT
dOPoCudVtgojxmTYj7JCU+X5Nzi5uIVrRr/BemphJz1i48+fi4Hzj0I/BKTM9PZM
r0AxhPlEuZcOmgXMlirPeWtoX8/gz6pTB4CjXXZmvKr4rs8pQQFgclYWg9hwZ3Hw
A2/OStuikESumzzl9Fhpg7aDkgYGccnlR8Hm94ejw40Xz6vKMugw2Ad/BESgBtze
FDTBraEfe3kmlCzIgL5/yVqCaq0YsVU0hu0TxgC0Xku3clcuEZCKNvZA3ecr+j+7
SDBhmIwDnVV/2GMb6uPNpUjSeLdI93+bS/KEDzh0VKD6/ZrgtsGCd+2QG1LS0DSq
0ky+udd64cGd+OULX8enzzqWsZc+8zb1iWgThCIxhlV4R0b9IeWF/N1C4vXPalP9
8ucyVx7e0XO/sDn1Ud1if7n2uGdWAW16hDxO7YIDO13s6QgPJDorjHmHzKUAsuM2
LJw5Pp65cJJ/e65HH8i0LLNhfK1O3BLuY2yWxFGUrhBp9QdRtedGykRMbhCHyo+x
i8JtuaYIeid+CosS5faqL1yey+sGj/ogTWGKZIWKk75mbAoBGOWGqJ5pWV1kHTZp
r0P7NktXCYGUsB9W8fp3siOKLEN3cUCZD+vZUNV46xC82jJVPCVQIGZ9gOmgLgcw
tEKqXm8XEi8imOt01OYxMGyvyiK1bkp3r+Er63w46i0SaKGvzQVUIwsmZl6oINas
x1XLqUfhZDzqscvwxkMbu5SmeF4M0dGdmHPcvJMs7Tz9cUaYHGED//b664J8paIM
VmVX+2hgUnGaOqFg8Dtez1E7tymLiynqyt7kkQIAz0igzbL5tyWMtOgdt1t4Avwb
6Zrn3CukGmSbKpVpFDySix/uEmrk1DREUl4zfEnOJUDh5zpmrf6yHT1Bq9g924cK
FSXN2U09A7YSqdy7vY3AT64z44zTw3yjSgR0SZw/qcRCOFWXsys+E5bhTHtX9trL
zsxFtedQJkN6zJiz26GFoVxeIcwYUApwpQX/qrXvlX3S0Hq0Au7JN4qZbmNYgbpr
b658H1Xj6VK44VSejbTSZ61QO005kwcwksjt8X8eUyOnKQvQz1uJ/w1YDvlaUN/8
U+T7vAx99qHfAZrXTij6ppjGJqDAUu/HDP2FIXtvLU0Gvc/MpXEb+AUqEpx9aRIW
lR5ULt8KY+A1fSE2RQ0b9nrLml0ESQu987EPBfjLstrEsSMCdOqOza5iblj14Max
7Jka5Gl5+fClekY9D3SsceJIffPC04peDCcmm0EEyGvDOcGruN2FCgO+fqtwSvF4
9Fsp4jepNXCDMOTlDTUC8c+O6Mm6azi8Jy9FS3A886KcDASEgMItxTimz5Y9KLn9
OYHQiWA6DmcEJtwE+ACdSwUepVa/dh88pTw9xcsS0Z7Nzwg9TNYfSvKgQSZKzKa5
zpFbOFRd7jCvZ1CoZJrZui20jgUYJYZIuSJAkSoPzKnViUfy2pJ6I7ExB53DF0m0
PXrPFHm3qH06fP1Qk9n9HVr37EgBEnsLAH1OOYEnmMAw3ostFFj28214S5Yqurcj
CnHkBAHGU3o4qjIIa+/8YjDqEtqNhY/yAdvGpiqcOcVp6PFNGZYb+c/g/6Nty0uJ
JiMmG7FRTDpVzagvwbOV4iHOi6UqGq5adyYjfrsIddRrb3k5onMMzAtdUoLd1y+y
XxjEfRz9NutTBuwYkrOMSsDdB1bM2qe6Fg84aJGnRdmLBs7tk6Gu2EpeJ9y6eDfc
PR0wr2VrMWCu+GX/b/RC9oSyB3aKXpS8cUX8LFerQXHpI2BOXIY+ibrExDXPbUGL
Ea2lz4LBrYHVZJ7StIxeZUNTDS70D61JTMqfuNVRt7ez3JF5JndFGumd0btQhGhx
KqpkxV0wHqRYwPa8eAdJGlqRYx+E01OkW7SlbU120LAkMLy7VZGJCrPoTStvpqY8
K20eDgBM3A5BbCB5XPYthdH+MSkI8qY0CT6qV2ftkxevpBmvqvbjA+DrGreVqYwV
sKaKSuup3r+qaIyjNWPfXda6anvl03OuQE8+UB7RTnnG2G46ARrrUDoKvbwt6fSx
sHnDGolbwZFguQYXEwo4YLc66IIAcblBhGy5TO10STU4opSNeaEuc1V34Kcp0+jr
ja67lMljLLtB5sLZ28meT+lZyhDOg95DLCy0ZmjqX7k7FgtTT3zCblciqmLVeto3
E2oTVXarPtuKUoZGzmJGRnowsnoqTZ5WwQGj3RZ2564XMh4q11WX1xS98vcCIjnT
j19f8MYlyKQgyB2+FLCnVSzPcwcXDi5ecP4fkjdnWUdubQctfA0l3UKFVEVk09Q6
ti4AtdX0sfK0ed69i9WPl9v3IP7nNXCGO03UiRPm69dLoalgn45MVKGJdbRg/h0y
6q/nIm1RSIw9Yv4tKsKz9vDGxEiRMX8WaEE9aQuP8F5M3JG5h2gx2zS/4TvU93pB
PjavLp15WpD9gyJAF5XJGxvVv8jhgP5W5e+UKyJbcW81Ansj7iavkIOgfGHe7nBG
9Y8Bajp2ksI4r//IJSSP/mk//LpRJBP3wiKmAJh50Axrmj3c5a+dwP27rXRgvQk3
CVc/wWVkc5JhlewZG/LST8AUkp7BGQuYMdvM+z+SQPBGU0Y/qm4Yiq7PQzK0taT+
U13AcMfI9Jz/k3LLjNtRVHMrJ9iAU/1h1rRnO2ATc650od6tLMjc+tQEyDkfGiz9
fDRHuoQ/ngz39jK3+zlVIgNuF/Kh3m2q5Umei4kB912BeqBzCuGihsxSTZ+sGcnU
ACwrnrZwL0JBlYDGSbN16ifV/n7a4kE4x0iAeuZQ4bO76100r+D9sLGWd4WgU1qZ
MMGpuk7Q4sVr+U7z1DGoEDrSxAseM9oDlgXcgOtmmzOH/snyUj3fuxHi430vuzp0
eA58OiOX35Ua7/+XGlRmj++JkDx6nRCIVssK0aOoVXibmZwV7n3P0DaPOUWZD7MO
tStiYFtXi4XYjknDGsYdkeavIpVOtQykg8kKk1fFNWD4v8ZyID01CW1nisHKtzRg
1XbsABjeoUNjygJxKxXUtCR6EjVQ50qJD7ritEZoR1k9YAGYwFlhE+5qo+ALoNm7
dFDFqdQzaUmtPJduZlFOcNJOAGFlY++nXbevqQlsqdVSv4pOAd3niqiVHzDrcXv2
ASPp6xLTLnDCtaHfdQf8r049s1TE/6nDFXtBT5ntkhQ7YHobC1H8TJPEoEE20XLu
m18r1KUezxpKz57aX7ixsrGLZVUnQKcZUppp/fZm/wPsAP+zrrZ9U9DCNUTAEjwm
sXsa7cbJ/rgNU9mpzfCEjqAqp+2GoeNfhtpmZSP0msPDl52siE4wcu1a8TSGr0Gj
xCyISJN9WfGhQuqd2+ctmCowGyRctCoTNpxGQq37ZbucUDw5oCNLM951yCwpZNvC
lSBPG2ks8ndRHxIe9uZwSWJC69BlapGVzGgOj1EDlprzI/uS3TMIfdIBnbDsvR3d
VMhMUgxw0tzfbu27iwwNFvT6vqRBrps0b/QAsq/qolaCbCgRTuixzD3Vf92MFTML
OSKm1NIi77PQgynYeCMP2uVOJ5PBPVLWDn/Vo0RgN5BNuOEFF4DKt6WCzpg3cbS4
8OvPOEIjp7vyj1EeZjKLxB5btcQUvCa+tCWwavGtITAHqoSC0IIgu7II/h67wE8f
vkJfS45I49BuXEOm3WHQBkXEVUKWcSniF5Lz7kOS+k5WxmQqEE49vAaw4sVUulih
N+vfSlEVFojdjYXFm1ctMTvvtn1kZJVOW3+wgPY7op1hB5PiKrST1WnY0XnGR7ML
JdQ1oHXbBgCdXkY7IKUr4N3A08eQr/8AtaJgBL7frzdrPnB9CtvmjXbHIbTVk/Mk
SRIacbXy6LLgfHkobgUjnljvZIbqE2U7jf38uTNPFeuqre+KI5hJmO322nxkGVXV
9BYmfr4xvtMABGIy/Jixw4u9nSiEY/bIvMQSh5N/mYKzajM/qBOl9bVglPTj5/mC
8/Hm/VtH62MgQ1eJ7ZQg7jEPjT8U3bWuz24b/fbLgKtbliFvgv0cd3a0+f7CQ4/k
VhFArZDkM2H2cH/6tOAwDW+b+8bUKZ9fEFSngqE6CqQEGVsMcGHuusidzto+bzFt
wWJPAYBAACVWXFEOnlMflqTTrfC92dygacbbJ0vtUvSdK2vUJnu+9TQPtVSaN5EY
UaDe9IA9JTh85IAoJgVmGAGbmvdRb05sQQvGxKhxDCvZ/1Q94oMBMRx7lZcqVOqo
2ZKqr991gM8oBsvuoeRO2+/SX8klSkVR+MGGbmRUqeZElp+mZRXV5Q4ZR/vpzBbD
6JgHMf8F07g0X2nNd8pvow3RjahijxmnbgajQwOKWiwmyU7LE2Vtqsyn6IxC2QJ/
tXzRObRPNVuSxihDPC6FXI6PpxmWQ4QdtR/0N9o72jdWAauwXrvV8YuhfKAijGt2
2pKgTT7c/JknjBwC+ujSZ6g/miNmWkD+thI6mXVWSfp+gvq1Z1LjnM7luckNMyWd
iOlvQ24H8KPrusy1M2vnb6Hk6q+2WNoSAZohNnP70cQamQzHxoyVkTDLovAm1IJ2
CcW928L1uf3vbTdNANci3Ixs/J2Xn0hd0J+0deslELbjw8zAN8ctD0cwETFjr/Z/
bgzM9c0dopdZg6vErbzexqF/VVdfMIoMS291NQljtm6n3WG5uU6J3znxrF/OCy6z
F0khMyCjBIZT4tJYAZRn7Co0G/J+m/NN/1W9M0IDzZIyhZ7qKTm+XnHXoTcWoQvD
R0MvwyQwNtzsULc2QdlNesdnAayJzZ5pJtUpUSNqKNZVwD6OR6HRhcKcBRYgSJdt
G58kqntyogjHhiwADuNJ5R0/X6id4984x3Kzx3ScBF9syrLAF7Vdlhpr08dyvvei
M+XgcyZsEYqdw4Q9l5W8S4+sEicuAnOiJSMq766kdhOdi6uY/73VzykVMflazoMN
J4AgcgndSujjT4ZSkxfkc9Jj9fzxuJUmb9NH8Ngl3Vo/OD4R3jGDHXhmdeKKHLYF
v1b9V2eXdZkzw/1foExTgB64IKsdSrhdaOYzML+XvBdqUJDN2zEugrijNAMRJWOm
qgFCWMOLAxw/5zdD9KevXkf99GxIgswdfNXrfz3HqWAiE30wQ01TpjskzCOhSEri
K73ajp9qBQqRxp/Dmqw97mDhC0eCIQqbuWMyGRbUBDzNIyNhCJQijEDE0ny9n3YU
3O5aUBmyBb0QVz3gTntX67mbXbPo8gYWBDpJSNGxBrKW7u9a8/DEa0zDp0wsSzcA
mVZoydh2cWdP+KCLHt0bbxT1SSDjkj0rz7UQplb35+3rYJ5CjJ6Amhf1PYKSC7oi
vNiWtbFfdn/LiT2q0teTSe1AaUs6eZO8z0aiKXRGSz5dDxa0t/ElVq7vibJOvpdQ
sqVEhw10CpaBnok1LQJ825eoiFQL9FkiMzxb96ktQ6be6aYUljxZ2prPbn9PC4tj
Qk0BaxisKWy8sniT86oDnJE4FrKU5WseyAvzBn70fVK6vhMjUICpHbkRTOxwxZG1
1j65h6PWc2RqGBBHuftNwVoWH40lKca3c1cK1Pl8xnWu5ZZDdA3/FgA8VPjBwYRS
9zM08hVOC5fryBiP58foCEuhkGP4qZWbmilVAe1r4U+qQ81/hIsJ3uqj/R/WKyFE
GPgbgbaOhARMs37OfahSG0A3RO/dCScMl5Ku1Ty/rP3RQs3OhHnZoIy8n+K0njcC
tyqZAh4NkwX7zmerDknpEgPGyjkJLrq/Tx2jx5wMN5X4y1WOpGVS86rYPSA8Zd7V
hM9+LqtuzVacjT1vXAnyRjlYgcCCxYVWhqrJhp+ODQZKAqvqMBwE/6fuo517ZWGd
EG0+WOqVshOPnRowCC5mHyVd599dN/gBYlqXosuduu8tMymQPbN1jJDGfjy7KVCK
/vfT1rGEZ3KlkfgCvX/GJE41KiXbGhENCcaUsx0z329E61UffuHkmlGDhSQ1ouxI
3b20Pbj/EoK/e5Tc5ng1oMe4TP5Zl0sBu5pOBvp2NZqus+lS4d2CaA9ETl09wuJ1
nzXr17LYvpHpPvfJSwsbyZcsP83bLW+bpp73a12tkyvKg8jqRXeDa7xkiXkA2sVS
kgner1DSu0K5D0fw92gqAaKyeGMt2EfR241xmKi4jj1yFUjeGnN66DxGzl4Yo0Hx
3WFNEurh0bQmiOwmmxNAMLe7GHkSvBJ4H6QvlICjblBGz+jdgZLranMtrCU6S8q4
xL+TniZAgF1KKn7vL78M/R5WFk20LziFzu+zSuy27eSpFHebJP16P8exibeMr91n
PZrrRSCOVjhQ1wE4ao6wYHoJihwBzl2ykPeNE/J3Vde3XLYlJp7aG3eut2MdKFwY
4SQxmQuVW3XaRDZG/+6QDkbR4XoIL9Vi6xsdHcsdSmFaEp3qZs+yYG9eIotW2ttZ
P4ZTXPJKL8AJYuWOGh7yFR7LCIZAGmbCoSE32EWvxI8beEjxmUvs0XBq5xmsMPgo
cc9az70blGTBkvVI0KIEg85D32v9hJBo0xcPa6txNmzMlaePRQTUUAmGDelNtQlr
Nvo2Vh5juaWHhP7RMKkPLB7AI0heKK9Do9fNsiixy+U3JwYoLeukhsNWoYaAqPEo
zq6n29GDNl7HIAmYxknfMxsVGTtDHnFfbQm8ZYQ0XaGXA0uZuo9ymPf4RTjNUXnk
d2T53e7uKoU1naCa4xdLOrqDw+WevruCWL0tPqDaJdJuvTc6VCtWhuv8JRBoRtYF
AUaSfBqzxxuMz3dQUxl/dWQGlUdhITCVIIWLiqWvcRcIVWr2XpjZMK2v2DeEZHtD
PBJSJvYkPldcwGmHRUY5GzmfLcoDjnZq2Je5mcNhcIKUbRI/4EJl7Kk8lgkaHn+f
3RoNp3UoePNGtNS4ciequHcegzPUZ2PQBUshalux8XYOXF6H1w0JoldCs6J4c65h
oeIF2KdXaKVTip0HoIQJrJoY25tCrsabEDIv3K8r2S2xi/10Hd+XJGj9twv0ia8z
uTZeKuusttVVwC9UKhsNvx7D00G2ZuEIXaX/BnQDa31fEZPCjh6Fod0WgzsKp9Ah
Xz+HF7L5XwKPgk9Tln+bTZumq4SfcDiPFytexWfZJp3VJYnSnYFk2lCPgfEm4QPz
WC7nHbY+0iAThRToNrVXm6gYUue3WrHHq3cRphIR/h9zNsa5NCZTNd6ftYKy7X07
Q5AaF+x1ai/MNVYk5UCrAZ48q251KBkqPc+oe/7h0onu3GEazaJX1iYku6gWdNIe
ifkdmGZc5YvhWfiNTB+TybP8TSo2qB949ftnSvqE9N4rEg2KoJOk0fsAoycTW6LV
3eMd3SW9qK1e92KWwxOITb2vdeRuNuBmdbJFBvtdgFYJThnLgSzul5mJCI8ZagVT
u63RW4xBls55eq/aqpEkLwHeyOnxagXLZ8O3/DIro7ogAI55asE9wenC0OjiBQBQ
rXPr7McxvRcplb/HWuTypdJIA6Fuv28I0TN2TwB8XXmGrcahdoWE0Si96XLizlfl
TqzQ43rxn8sxMZY/H4WIxF6u8zNIgWtmvjSrMXzB4qzIB/ybnWMAPgZPpvoOQ/w3
zS6tkv8Yn80wEf6x0fOeDM+3lVQag6mgcbxWAepdmmr6LkphmTYMO/wy3QKe/iKI
naDpjvSlBPxt4acVqdEAyZwnOYcVyriIaI75C42H5xJheVVvDjl4/mno2HmiFv+s
O7Jd1yCGNyv+A/wE4cPLYePsHqiEwWCcLKaJCS5/peVIqM5A23QK3rrPxYkMB/sW
8iL1AquhLlUYr/oOVKffr6gkQrN8SMhNaXD1wDTVmTm+o9Ug9G+SF3wx/Z48S3h1
pkoI5nlc/Pln9VJzX+zQ+r2eVESR4k978HkdS735ctNKTXBYEICFqhxIZWB0ILZs
1U+cR/0Yr1DGGgqHUk9RRjzpVwGTA2k+mf3M0q7pMRsOvIiv6wlcFxMKrqIMJlY/
ulgQ+FgbdpDq0lX6uTvbZgY0hqu0vunrj0+NsoBZ2kNsCgM52fNyhjajYnYdhGs0
bnRfcOki60IGqsFS2uVpBtKFS/gBWbMBa9w95eOavqIn/UySpILlUW7I/7LX1ejl
3qezUp5UGz0snLV8NcxQyE/YlU3nRoU0i78vLH9luwbMOd24DDMHDjj/Z9podEPD
+koMlAND5Ct8yTSBnwPCvGGPHbs61U3NzNFxZa0fD7uJkuN2kJuf/jytWdpBfb0a
bnBUyeZ7vRKEa+xQbvYBc/VqqIm+75cjLqwxlt7WABiwTdEa56j3gbq/Xf097LIV
1/YS6Y7McZxO0eUV88miLFFzQYs3aK+TENEJJADDcIGHcmOZTZlb7qI54pdVeswu
hsUGliyjhtlSAhoudXL5K4yO54ztDxlNDE+zKnah0ghjgT6NF8DiV/hmp5MEvBY/
yaOCFEbwLNFdgdZfa2UxLQ8LyUPcK1mfWq6IeRKAUJIXBdhn7k9lQIsSIk0tqVyu
wxOW+OMXZHjLr55WoYTOWQtrGYJ1KEVim4o1gPUlPtT009doATX+pGWJLhJDsWPz
TUIDJRCv7DfWb3PcNHxIuUCIMOqXCFN3jcy3qGWDq4T6Hj5J/1xETJftsYHno6K6
G5+AzWJhvJroSbmEF23SlnPq0hjB8un5Yps3rGawAAwpkGtOHNY/whmLPG53dH7k
RVU1hl2YWaIJcc4t+wg2eioVtewaQRcp2iTRAMO/Tq2Ko7K8b7YXZk+ZKjuFlhzY
6K1L13M8sSSopN/F8SgIrpniMC6gJyJPHd9cAD9w5/39NLvDNPsiJW3j6KeRMEuW
eOrQU9rZD6zvIXyWlTzYqtNzoifWGq3sDecHcI0n/NzAnlN0f5wJmhR8D5uoLq6G
QJjCb8e2BfStg4GiGnzyql7v4t9mRNfelJEPsnsAgJYhDGuRgZlbWJw/13dpcNmR
jqWNHGiwHxAGDQ4JoXHl/JgzFggRhvFutbs0YstUcdoQsN3Dc4EsmtfHdBPUJ2mv
RBsa8G3n4H86xVxO7LbnGZ4DQvjjYCfsHt7Muf3LdDLWi+z8f5vVVqsGrWs6yIkQ
eKWhFtY9paaEV33c7PVTL38DS9Ouo8ea+Ow7joryV+MKtZb7/PSSutafKnajOiep
qtrZAAldZ8jxDxoE5YLfKkpmk3D2toFDYOuj6pfFz3VI7LVTNS7S0RADmEyXXG3c
wJwjtLj/URUr4ESIvt8QZLiYWA0LJ1idPdEJb+Pv2Ba6Jll6lbe+z1FO2ja7tLXz
vmLWUxTw6OcHHPP2SwC/d+ThaMc4cUXfePYU7DjojveyI+UyJoN/IHK+1ZEX3L7G
zQEhxuOQq2BP14P+kzRko/0cMp8I/jdZR+lLSGozGuBW8ZmRnD65v5vk67/4hcD6
VKzfefwGuOYwFg5m1BVgI5T4jBE7qoBYoW0EjxWkSXxgKLF7a+fOqy+ScFyYRJhB
CSpoyYyLSbksyVehVRSjbxCvBCD+Ee2yrQvuD+JOVkgFt1R5mk2pEwHMTvhR23Hl
tepFugLP8M9uiUy5rk7NJo8egAPCs6LK+iUa3KLLUseCGrvmuIw87scGWBisQzu9
QuEqNJeOWwfz88jUM/E8xW8STO2BAJvm12/bXXJSraTll2Ex3tCn88BeSEnvzymX
RNHGr8JpeG7tgQrvGid7L6NwEJuVTqvtesCTWtbcG1ZL+FcjlX/8r3KnOqihtcMq
ueiWfeZ/8BlOtFDttPiJJa8PJq2hyMBrE1wzxaElMJ8zak0K9xWYa+LHuUSkU+2c
LsCb1ybnpkzRHScDzD3ALu+vJMZcET0lWYhiVQE1kAM+Mg6v8b7hqHkxSg78XGus
KXk9A+WTD4unWMvGRvstN3J1ptARIubsvB3+yvg/Uk749MUWwy1J4xoHSOSyvWCI
1JnuJ81YjkA5vTuncvy6SOn1NFrjJqi4KdaA21pqelPC/5oQYQ7iFaCNPUb92pe8
XgQCpqz48RLMQoANulBmV/RtqltCTIgHVWQMFnPT4Lj+6iUfZ6xWsvH/AUjnmjpe
Yko3xCv4pbfkGhm+pqQo3t21Jaf4klH+eZg9aEY79uW711M8sUZzZopVnC9s471+
ftuW0D9PqcEwyK1siktSs9nRnw7fDWHCJiLtt3yLFReUTBNVKApP2ppVuhhcNLrb
tOe7yNyc3AzRh5N3Xea5V7QyjzSgTXAXbuaG2k4g7v99A2NYFWplbJj2I1tyccGw
7fkZB0U16emOyDRI7Zb+bc3qPzCtMN3DiFEeKvQ3UkbGcjb9NnaMXr674vPi9EDi
LuPmg0HlroxzS7byJB030Gpo2M3nhSjOFDZYsx7KjCRsBcDLiRiapNl70FYJUA78
wgdkQvyRDor4E92ou/gWDKyejE+miFrqgSu4yiJY+yIro9fKDsTEmUUCHGVGONLE
c27DHc862fJeHLprOE6CDviEqa875XwMi7EN2fKhMuw92r0O7x898XEEPyJPYjoM
9ILx7ZI/7FAvabtRx5XW7euDE2D3c8YJoganSSmyULWpGl6+gGJIm/x7vBACbJoW
OgDc7z6mvo0DvynfYfVofzJwGdYZRcPB7Ph5/4MkXMX/WhqO/Q70L0fC+Y/xach8
XVLlQdryJm8HOBP9wLXVFR+ViLsR/szeLGT50dNJx1+Gl+QggvHPKL4MhZ3qJ1TX
Un8GkLPTSQjhQN9AQyIrHCMYaqcl0mO3iz4e883Vb5SdsM04PfB7C2kEVKQUTZAC
hkAtWcKqViFXhDV3RoBTAykQTXiyyLmPIjPZdAVFM35ZhDvpcS0VQq57KfWoEa8u
f9mzok5DkTG6EyEXynZTpH07PogcHvuWlYpUJfAO5T7miQT/WGCOCCFui3NvNiRc
tUNPZo9Ju8aap1JTiw+i2dVs7qVICmh02csiYyYzS0DsOhkpEFVr+rKAbz8U1IMq
g1kQ2XtBymGE8SiAmk0dHByaZYWjqqo8t11p/4s8Xp8/atLDAQAV8tGp33HDzmzX
pmPZZbQzhvWDW+bdJFqGLeX2XRLJYyuiHRQGIf4nnNexFye9zmMfYJsas2d0zIQ7
4binI6+bFN/SmeogfOyw5/N7RVmw1rd0xiU91r9p4B4MoNbPSswNc7Rs8NZeTZAE
Ffvbil/+sn4Mo1E4Q980KCQBHStIFdOD9QLIiBP8aU6IZXOEWrcvPqbR+New2OD5
d/SqW1ClsXe0SbHfvtKUwTA7B8L66+BcNbSScN9gGAkz/5BDWRvaruzZ0Hn1rCu0
0wcWA0iBVaP9AeztnGDLLcg395Uks6idwmtqeWH3iY0OfckN8JGGV91/ulMLkoKj
gfrHyle9tQg9F5hK9g/0B2ub8VE65k3W7NOf6C18Q6LPuv8yAsYoeT8S5KTwVpl5
voS2nlcNhtui7B2/mhwwudTjlbhyRwsVqOeOw9ismTJIYtbpA0jHCzekrr1M89eI
hd2kyAU+4NB70otR4a5oU2g564CwR6gVjfzlbdQZpyxsQkbj0jHFzQhG6cxzA09w
8Uzl/Z2NicSRmXYIg1buxSVxj124QX26YX0diuooTitx0sYJgvDbJN/w9w2RjoJT
Y3Yngpi/KM6Gb1TpyeVuyNq+aWHwa0uiit3IwoJ2zgXPiH57DKiFz/7Woom0m02i
jfabFHoKHtXfkVdw1fedLeoYk9uYU6+4LLDTwVvB97LI4YS4m0P/IwO7qC1IrFhF
f4CkKdeX/qUv+wB1DMtxcPC+3irXiEb8Xy8cjytIpQs0hsN5OT7YouZ0Q7ryuYu2
YOj21Aycv/phD9kGFVwojirJ+hIMaeaSt5rKQf4c2rASTuKa2iexQPELwHOYzf60
b8NrV3FKLAPJHFWVjh+3epXVFc8GxoIrAkAu3GsqjdxhUddhiTLyQf+9rN+D1qEC
bBCO4gOZmhvSYSmBMLdEu9COcnB3jRD7cb4hMLcShygFBzlDTRc4ux48fNSlgRoY
X6sDfKKHEj1ILZa9Xj5Uf576+5rWQOSX/eMRKYCq51m8VY3hIFvxeERCmz1n2EvP
Qq8qyu3N77yDBmOGjNJnEB+sfo3yNP4rQ1d4RVb+MjwoUHceDCb/VOLan3qXGiTl
Jnea5Nno/T4DcgLnUtNHznher19dXJJO+rzPm9jeKNbVBHDgRTBRg5AwPlmX0hR8
oGoTP2HxaG8Qim25/8UOtK2gTkkIuYhZba19OuhlxRU=
`protect END_PROTECTED
