`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42Fz9kWBik7SS4JBjCDX8f8HpuZ/LhcBJz/Y0M2kcGz9
8ilrrbP9KpEU1wqQDNi9iP4zwFoYiGReKzi8cQ4Do0XhaupggD/95vM3oGC/yqQq
+EBuPyATvjDC27oQ9pGVaTLVFkbdkUHuG8M5l8ljJTbaHkTkyZN9rYHfjpbfgUVe
HegMbFw5GfcenFrATyFI5w3Ljlvhuu+8lKcDA/h4huMEdVWQ5a5X/PNznzjjq++7
hz3R4YJ8RrCK1DJQkWj3s9lZ2H8u+hmfcE/l/8614gVD5iD4ri17/JOk+TEozloM
ikVmv6ooiBWoUgwz3Wyo/plEPJYAWY9cMhfpJ0ugimapiK8OJpKUoz3hOMoHYsuR
hJzjPlMJ7JNKCiqlgWyeqQ==
`protect END_PROTECTED
