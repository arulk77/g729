`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Hs3lA4rqSHXgGV62msSfckVPk4+HH8BWgAlCtP4Xo5Fh11xWdvXswX3EhBZgpRSX
gJkNggKVgobClCbdpEReqx5FUmEE0QXdEcD2WWTQy3YKrbygbwzvS+428WApviTf
72sRBO6YkXBHLRnnpZ/5GOltqyBwpIzyNQvizEDv2yNrcA/o7gbtCoVjM64G34GJ
lu0nFFl7iBhVian1qIEeEw/MIYO+Rxs/g8SCo/tvQXte3vKmHAczhV0YASPkd9iB
B0NsM3lMz4oNl5qQCRlEXsoLAbTWtaNa8qGLdQtXkWxavw0LzF/NXSvE0VlGvgJ/
J/c92qadKZumr3WOMLI56bJ+s5LOx29B8HO5481c8zZEC+lTbuZyuub/SqvFAdS4
UIA+1ZbLR+/yIvYPp4hte+Ypww2qZcbT28Wchz6nCSZ5PGLeFsfVMkRvFj0I19cD
eoJSbqAi+w4iv3rn8KNq/zL4idDPU19PXQ6uiYhE8Kt4BpBuFlfZfYrqy5GaIWOT
f7z6IDi4pFScUxOwiG2jAr4MHELPuiPLHt8TDdJzYURx3uWMZoXBzzV6k0PBORZr
uVgtAcN2HuGuGasd03LUa5StlxdMyucTlm84gK+6m8kw0HRr3VEsh5dTUZCOdS9f
gV8bhG4WZc2RzpeE3p4Jnw==
`protect END_PROTECTED
