`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKOZGSDLJrRRnsFzOSGHpwBQ6+Im7V/aC8dt9eMIku2O
zjGROPYEGRtiXMy61u/0PAxrdLYiFVuumQyhmdvzpiSuC2e3bKL3BZ5dnxXWuQqU
gTUfGNlHqW5xU5liXAMphSG/hOELKn+7F79vmvfuJ/KNm/XSEOhzxQgGX9BRTSKJ
6YCS3UvVjxYw+l7sYaOE6Q==
`protect END_PROTECTED
