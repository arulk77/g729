`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePdSQtWp0hIZzXk1o4B+T3wVL2NyUkwBB1tG9huaHbSJ
ETdhO9kE49bntN5aLcZNvqVyEFq52Y2xPlpz172uIrsMC4WGHQ2WpVlfAKd5+ct0
ACGaIWACKUEedN/7P8RmF26hhp1X4mQYGu6Tuz9hV1iE0iMnvz1JNcVqUXPGPEb7
bRGCsHCB5d/p7gNstcKlabsz7sVOi4r+xz0W+DywJspMPzRIhwnieSb0XrUDFYR6
V6AeLSZygVbh/OLwZGe6Bm+uT3PsWCfbMrkkhxjYnvrDjFgs8BgdndpJ0FpYQw2p
lMZ7dIfL6hlSwJejuNE3tA8G0fgFX5Pfycqj4BBwfMZb4vA1GxsDP4VBHixpVVl1
KdaXkp0kKZz9SwbqXXz04U3ssuso97fKNQsqLmy5WemLfz5z5AH8pKyzzgUvSCJl
/uqJ4SE6yFEW9TAG6hIVAhNPmLF9su7sFLN/6CLCLovfoWxOYo24CnUTzib7Ri/J
FpVu/eS4M4W5QLRlYhNVYfAza+f5V7OCBRa+E8L6g2b0wnM3PnbjCGYtoZ9UwTFe
LaF7ha2CUp1SU6fUJksLUsEYVA2oVTezHMul9D70hZgP5lf6IzK11kcLNgvlD74x
Rrl8+xa/mDLUOjtIt22x8ElqNHxDR8bhkWUV30wdbOm+T1YFtZxre/Tj//KCIcs+
`protect END_PROTECTED
