`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCL22iMHk/fPGdhacvc+vUZJHy6cOQ+nX/Na4xDb4CqI
Z0OQLrb5Y55wglXsjQBk2FI8Vk2jCH02MqPjyYeq/vI1xispfpv2s6g0BEr/sMlW
GYC2VLOi+8s7/965vulZUig6mSfuXlpmfY4JvWMzH4Ww3Raz7Tm2M2sQWnL82tGL
6lueuwQu7Du4m4IWekNygYxhXsK1It/Dp9d/y5zK0CmbzxA2AM6oR8cn8TH7rjN5
NJgnu9H79dLUHSpBKCy13noHrJrqIx+S2hFTprTA4hilUoXgMVrPDpTUcsFPl/gA
Y0NubkzooL7gEqj7fbDa7AX7gBxh4fUKxqO8y6pkn9yF6w29zhDfYQ9v81DOGsGu
g306KIEFn1HuBMtyQpOUyf5sG29Z2IMkkUqNHY2V3vXpGY5Fxr53R/1bCtBuQjd0
+4oXBc4wpXa+JjzY/c7fuu7slAOXpJT6/rbqv34u//uqAIzjj4w4rLyJ1kitN5d7
lg01KhJ2FqVJ9i5xXPmznqZ1RsS6Sc+5ulWiNwj0Udh4su2gM+kshKQh65li8dF0
ZDDZXNi5f0L3+BFL55eYcnFYYn1csBt5kINa+FVjPDa9+9PL6nRWrBI1lQYTTeiu
`protect END_PROTECTED
