`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEwm18WzxfEwYP1fc/WWb4ABjKPacckDYeTLVLbAZA+/
B7i8Z+ISbK9qqbWCeQ1gxEhrA+aSw7VjN/rDhSBEqFkiES1Fnm1JBI5Rd16T1iG6
PVHB8yoVSqSV4eRcUfw+cVpJELxEG0MZFE8G6OmlmaWYsolwPd1/XOr9oFdHUiD2
J0pihHxrZdFTn/Oi/yhLq3A44myVqOy8rbO+/MhyOj6hy+2UFunU7EobpSxbB4iC
trLyc+vYh86KMU7w2O9Y+O4Cs7jRbfl9gvkyDiBmDieHYBPX5DnSrBTtxZMbDaLc
glWWHr0KQIDVl5Nn1WlaRfRQIV4UfhZuEy8/3I99Y3/8AacDboP64VhJZZz1ZgGn
jfiJtbeA5SkPxwigz9meiw==
`protect END_PROTECTED
