`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLN3t2WKZ8LTqqLiAKaXJ9ftotclov3iwjVTZxA40u/B
tlHZGuKY4+vUcU4UGUdlIFrOU8YTzZB1uaPX3vI7Z1EfCGK00YExZOedqzC2jGyp
7GJ1R1ukG/7zP8X61VVjHH2eZ39iiVonRgDEWSPMKQlaj1fZwdy7SfrT2o31lYC5
K4Uc4K76ZpVtZEyj6aHVgPd5GtDKuMqwndNPGu24Nt8i5Wvp7w0+UUHSFtmU3NhA
lStn82nwiAVehPsZ2Z3bmtHw0wo+cAeDIwAqzXxmpYEGu2j9a3ExQgP78l4tLKAa
jcpLcY1KZ3QeuHMoxg4bDgRdUOwUhjBsx1Nz5rfnAkbqPMW2ll7W8NyZQUbqliuA
MJI63RgJshdEnwMPLdDz2upyzpMKjbS47z3x79FK6ZJxcPf1mgLq56tH0AgIllj7
mE4zX6BFXE53bXk2MyDL9Q==
`protect END_PROTECTED
