`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBsBOxtHy1BwPRs3R/4UoIZBMtGukpdX241nGWEx4oKm
RgrZaqpO8vND4EHpAOsn5KD+E14imyKacRCxwsXhUy6XXlzG2DUQwWZ0Wkeu1VX6
zeN+IqNVXiQGzFs9Or7R97300k1/C1DeDi4jzkOJd93y/R5Jz03EHyaJdvIs7UqK
rluBOhKIIBB2cmEnjUIHVeNehTJ6HkDKY0U4c2J+KBoifmdXaJvlXft8Mup8lVDJ
DdK/0dMDV6Zf1E4YBZevEAS8SlLo8SuFRWXk4N9Ienv7CnfTxJYOQd2YMHBdHMcc
XXNVQ0F6+nTJ65UGOQzp5n8WF7V6+kpeLiy3FMpQqUQuZjkr3YbETdPeEp5Vv7Ry
Ev5QCehzTeKyxmynNOfhXOrOMbHdFQp9Up9x49ij0g4CWlnYcOCmrVKsmag6C5mQ
TflARBzeeE1jM1aloQMlElDar7B8Bl8Q3E03KqMrJIz9xe+Tyy9lzZ6uOoJ6PjvL
ZVpdRtkRyYwKD6AYjwKJzsWbBXbdg3fxxM/GsEHpuWpaKLG3lsTDt5B3055Ygha2
`protect END_PROTECTED
