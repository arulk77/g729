`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOk0zM7Mt5Fq2rRXI3RvVlRw4EiLtf41ytxgQ2VWXQj1
/R9fiqa1FoUg8iQ0vEc1TBtWRDnpWm07KZM29xwDS5Sh3OTALmfOpOyVvGx84Aim
vPQWe5ittap59M6vrvdVBmb+wASbhSUfFKEBSV9O8u0MnamUmxMSAp1nBUZVFO1e
kWRI8HdLkIuPp9ay1mppgbs+yPV0IGC0X55dVZQLtMtAeCtGIgIg1N1R/+2jnXFj
Cfdk/pKl+OS0D4VXepbWcA==
`protect END_PROTECTED
