`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBmHd0d9mlva2GMUAQTtUgsn8mBdrtFVOPCu0RVQtv10
viCVqq/+rzlyTVn8KWgWWNJhy++ci6MK7ATaclWTiDzRyVghaVyTKvbsovK9IsHW
lkV+6iGE828Iz00yXKE5S3mA895nHADEQTvxweMWctUkwNwGFNJH410nT0kSbFjt
WtrszIJrdeqvWNJM3PET7xrKOpe9btJOZ706IjT7i1tTURwT/27zSh26CjKDJu8s
i/KCjmJI986AisGDOTJlvYsxrLIHbvvkKeOke640bYcEDcHR3vvJaGoFVwtTLQ8J
PFOsH5Nr1SYZxliFPa1d7NTdbftDJC1SYga6DK4NniEPxxcHz0vC+Bkx2ihIIgyq
a6XEV13wOeIAAQJelBD81lg0QXgH88VcTuJybhrAuD4hjWaef4nr2x7aMlkwgRzg
P6T4Zqt1L5Q571bQlToZ92atTjJk+C8rnZkP76BUx8Plgc2k4oVK+Q1psRgu4210
`protect END_PROTECTED
