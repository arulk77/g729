`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4ycGR4SaM9a+TjPbDBcwzuXhVb3fXDB+u0zWfsa97S6O
lqwjVX78WoT3c99Bj8tkGLaZFFd41/SgpzLL4FO/A5JjPNAGdCRPmRy9lRfw6+i+
i7Fwj/19cIXxIbvLrTe4H4hH8ybv1oQBzeFu5VRwVz/Xh3NNubZC1k9NS0Vh3GIR
6kvDQXz6rbOX63f46uh/33oAd4TxcdOv6TwnuH76DLYM1/Mx4XHzNKuYxLK7UMae
f6UzV3nrTuAVJE1Asuz4W9ra2PTAe/JjshST6hU4PZUOAm7+XDPIa4oVWcIS6VP1
pDpjxEpu2l50CuIwSJrLpA==
`protect END_PROTECTED
