`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xrDM9jhnjuFbLxPQDcRlyQm0aDHblHhVO5IR3t4Ma7O
wkBsHd57ppBxz204l2QKYNd/mseWojtB0aQVxuSAD1G+DeNUN3I+VkBXskSao/YM
BWzCnzx1Bv5tYDCOX1LQK3AGo34orZPPKN4GL/WPUMaiQoSlnCiY/y2Rj1tMvFhR
PUvY5dSbrBhE7Sox9+/VDgTX7XK0UeRGEICOF/PtNW/of21/nmcKouqvBMZCMXJI
dCi/atSkpRFO/uow0+z24i0a+lgYuzJ2ogqDnI0YHcL6IzMtaqmYD1xL1lXAuWaG
XPvcpX2Lv4hLQ6DUjj76oA8IobCIXT+vlcLdHy6+7WS6ugTIb7JD02Ej2Z8F+mTH
1vVZIgeft16F6vo/oqW1ZA==
`protect END_PROTECTED
