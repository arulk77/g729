`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47iH5iZXxUvjqiv/AX5rxC9rm4wrAVOa/Mjhz/FGMPxI
jLIJ1uPDLTL2Ul3o2wVFLD4rEOOiSrW9wolX/tPqdPKELFNjp5BA6nOt5aj+yJIE
Uc+jpAuyCMed7oUcXXpAMO2iaiITJqAjgKbdkPU0chk107BnUeSLQ5nzYGEim4jK
FNVez5Kzg0JNgJshulEHdoV/um90zRwFVrG4BzNRI1w=
`protect END_PROTECTED
