`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKPcVo+cWvJjI8HFXZk/qz9mmYVeLeX6hR+f25GvZQGR
KODmfZ0rVnsvgRP+pG/RvldOR8IWPm/VsinzsPGoxrBEZLDFdR2FXE/ajpaVgLBw
oXnUl0Mgz6BcSfV43+qKeZvFONLMF5oqsF2QsQ0itpATcs7vM9wYr8v6kKIB6C7r
1PUwI8bj4nSWN/kdTJw4HNqOp8Dx65WEDd7FVR606cES2pIX8QDxgF0fDb0Fw/w+
TSjT0PVkoGQCYJPKJiDellbhtSPyb41uT6kYM6OCcs1M9JG+il6p0pmIR4K/iZj6
pbLWOZvm75bWbVEV8y0hAtwmy1uECsD87Gpso+kmyDRy2sFhIk4kMEabaX5w4mVd
Iu/emWHncZkEtj+DO3t3z63zY2IE+6Gvz3qruqb+n4u0mNgge4zsvBHqdxlnEIFI
pyqTbDGuPdlbWyTInQF4nhMmIcuoz9xreSQYEr3ZSN9doXaXHyVkSYzDGnDURrBw
wDeo8jxbsXVBw60kWvawWYb2cvAnL7Pi49T1C6/APTXqC9RUUozrMOdZa3h224LE
90+SleCLHieFaht/EsMvyMVhNz1iIuGybjQxGALiTQ8kuRR9ZClpenpNQi/uTnf6
FmWQpNZVbBBaddnVOBG/2tDH5B9e+3OLa0gTcSnA3YGVn9WPsi250odO+xPjV8eZ
`protect END_PROTECTED
