`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJyTvFn7O3jK7OPK7olXHbQ5w57zExFQUs5FKEvdOm+g
0BIMHig2SiN43V6QyCbKqBEbiHumw0nxs/EDirmvr66km5+rT6W+dvnKASuMBgH+
8nICZ0C6Avir3Ixl3PXI5NemUxvE9MK16jQ9Xu/0PqkaWLfKpbv8Yo+hYN8JMP1T
`protect END_PROTECTED
