`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNnDzqt7CwtK1smK0+wsfxb9rK75EiC06T8iP4BLsjG3
QX0NbJquGwviMfmW6dc2nI0l5Tcz7zHXr4hwmo0Esi8cDMxLy0RJEeyJzUMG0T1j
JskmMsR+2gwSOoqXxrruhAg+AzbzQvhIrEJsl3aQgE7jGXCCkgtIKRSclWIYxieV
uWN/xXu0T9vfLsIcl/Q9PHGPTktCUT8xCBxSiiHrPRVu/ybwmPQuBFvOU2fVbosq
imbG5Shjzc6U1WvEzgLpiTCLCo/ApRjgXv/gATFhmidnDN5yMtwq0MIrEArmPtkb
xqXZ7jK2s6f0rJ9QiuqlQGgYj02YIm9s6yKZvQs/cCK13OoN9NJKCSshKUHdNtNb
P09zn3ILmZaR5PwAXxDKFkJynnRTPJ8afaGGJaGVcDs2HIVK4cyjdIhvPdY/WmrT
wcSI/OnIzzE0sEXBC4dtcQ==
`protect END_PROTECTED
