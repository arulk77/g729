`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK0uGVahN5NU3CkakZ4/uNeiceYRErQ8XCPBAXAV8uAi
RZR2neqzJ4MHlhLYo5xAp4xsy42jM9XvqBhNuRblIiM10azuLJgNTw5ecjhTuC4f
rPwGPyGRifOCizBx6Vf/tD7UchR2AZ2gZ0ubVyVYmT7hrDd4n8SAX67oYKh3aE6u
kDTSXuUP7nhatVWxb+zIFc3UDqYQVZc1T/kJgtSGqvKJBHo+F6girphi3kIiHSLD
7T/hQiDMZoxCJsawvMjqncLmzn4f9DQHpOomEP6CUr7loZqhzxMOiaDYd0SCZ5er
9pWebQm1xUpthGuGOweV4DvevovtE82bjvpRVGjAu1y3FgKiIxVtoc6r3ww5LGWH
RIHsuI5gyA0BocpmPLQi17QEnUbBWBia30DJ6z053rUBrjxVRhDpdsUXv+mRZnd1
cN861dwc34TQaYNRrt0uOrxT8yvQmgJGXoiGW88mvdn3okY+FrON1kCor0FAxWMv
cCz2b19lvwb4urB7yQ7oVDA+W6iAL3KmEZG1bik5rffdJlNN9xIizMwEwH7qr6Mb
LhrQ5NfTPR2JeXs8F2HqrWuJORb4MOrfOX/2EjOmXTVkeu0EDJ4p53nbi74Q1oaK
jfdMgiood+/vEVxR6Qy2WzwBq29T9WlyKRul43AmH0U0n2K2vUv2pTOmpks8+lUG
`protect END_PROTECTED
