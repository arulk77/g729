`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JEtC00ldjwvHKYhm7tvefoyMPgM83G+9qjqRJCzr8BKDBjtTScMO27gLxhiPFmYY
8UkXP+3AJcgzue8YYxk/RMfhVk/qJqIoAF4NznjAcO700co2QWoxQ93OSC3n4vVu
ZniLJX5DszQOQqB7N9jt8SIpB0GGKupHwJ9igDZriS+N9i+5KeJUruYGFm33Tawx
s72SEl3lnyqHa2Wmv3YlB0wwZ8fm7bjDd5t5mZCfuQxECcC3aStR5CfHkwLuZjC8
AIQ56zTrHG4+P++7kD3waoIzDxWY5z4mbOaLbPzSiDM=
`protect END_PROTECTED
