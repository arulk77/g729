`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SelfvVXVSZyeCBcM18WSpX9z95X6C+mctd7OR3uD5eHe
qpFSJTA9ZuDK4YHidgcBVNApH/oj+lxvDT3pYnF6zjoAW8n+k64Q3bqbzICoTeB6
AqG9x9YvmCehDCo3xaoz0vx55Wb7m9hllmk7yCnULa8yt4i8Uc+kLwLqxvhzFrHw
Ot47QOduu6sdudIn4oA6j6Olfo+fCCSZ1F+6NASUDFYxKyE1n99NL0FtBZiVnhho
W7dxRCEbKpVTyY03D1Kbk5HsIW1qSQ5lFJWRW9l7wAko01OLdJgNn399UGQfua0T
+DYMPGlcgHjwdYm2KdGyblLIYa6L2LodWfMXiRTj5PMpLYUVtMvHwv3chE/2HjVi
oG3AdHQV5zZ4x3Z5BGtPNWNJQLaecBW5h663HaFzUcg1/48if6Zby9p/247HvvyZ
DYdNlonsTM28mEfmfKAuaj3kLZdoF0nwuIuX6NU7hEi8hg0ClgK9BFJDirrr13Os
BJ/6k5QrtvJ7+e7fc5AABbEal0xiv5pXoY5QYNiaRWZjC5flhE5aJ3IwXOhkV2b/
7cu7n7duTLfX47AKwEhjqUbBcORbZ6yLnnO6gsJwIBcXre7ouFTSMizwQ4dhyojv
ifa9ChTNBU8YtmzkDb3mpr9HSpGzS/pevgMoFsX3rG7HlJay/WoWDzGRG4nMGsn2
gdZ6z7HiJ34L5PQRR8oGlhr+u51SiqpC0H+2hrKxBN5ftHuuFuLI5ndHw45l2q+D
J8bprP5jLOGc4op9Z4t0cLkEuRL5Wxrh9vGN4id21YIH0FhUzQ0dET9y8Vh7vw/o
awjbENEWD1a9BX1VpP/jucVPHg49V4GuMuWP60KFbtpNH+l8SjXcx97kpt6AzUdk
VB96ofs1kWD6qzMygvkSfxmJE4MmC9LauD3wGUaS48+ZIYgYV/bH+rGJemSqTc66
YpjNQ6rRnVbz5yPHP2Kpdq/LNWHW2XeKQxYEsW4le2tmBlNImPn1g3znLFbe2gNI
4zKYEuWwq1Sdvjfdd4vR5NcluGgN63LX9mnewGw0cfQGW1QYlKEbU4aUPyDgYyR6
mgbzbKXeiBKvX8p9nt1rMnd7LWV5bdLcB4KPxejwQ+BW22BMbpu5DMgBhgLtGtTM
xHl5Pf06U0g4k0kXzeq1zDt8eFtc7L1Z5od1N+0wDItCUYb7z6NvlQrkmmvjRvEF
GF7X4Ltj604zEg9DQJJtjigZVbUtP7hfAIsfKpMY2YZ2npPQ18W2h+zkPUeEWRbC
b7aNvddzKbY0gw4os2tpeiSP+6jY+BTawOHuYHbPwKT8Tef28BruKPpw3ZuA+4IP
qb1AtclUFD4ex1uQWkka0oSUi3gqAA9WrObzZmbE3q78c65b10pTvKvAG4NVLhDj
n81Ja1dAlCaBF0yw7JXC2/IUbQ08iVnphOpWQcHgVtmedB/j2DYC5Wrq15sFzQla
aqse+8HEJnMoA2SN5UBr8gMU1+qzcLjv+kfe0qcG+ZZAB0Is4VedWMJ6up+2Eaew
jPZdqcQL26Il9njgQF0TBwmwJpvy7ePYcVKulV92FAWjB05nsn2Uj2YXpnZzWG6H
nKUE4xeLP3KHhlOip3OUjxh8MRUjxG3OaqmPESiWIpJPoNbLYYfyi1MJ3vpyW2a8
CCCz1lpI/0WKKDpBGYH39fRMVIIrbTTuWps9IBfezXxE7aQfVmu8USbs3bmNca1v
rAnrVPzC2ajVDMxXdgEYvCeDPZrc2UwyUDOS8+q/4J+Sh7cqJ3eueFNI4I0E7F52
ufQqCLEpwtLiLruqEO7adEQPs6BGmKRns0jvCyq5HSqopOw11AlOr6OqmSqkw3rh
McVqs/J1UwLxz7uinGay49e+7DFZY1KtoRNFtXzFE6eX9o14/o49nnCNL3QF9Zo0
Ip+LFZi8/b6g5/nfwkDdQHf/bohacL2wp3hoe2qleN5n3+ZDW0fYuZ3PreNkt2FL
0yRKNouHaCOFIfdLWBj60NKIyc6l6Gg1RaalnMtD/W1DsCdzv29y6/Mo9OcJuovJ
T/Pz77C4fDyyiC7Mdnq1/soUPjVQ+aFm6SmOjWtCxxAlNw1GKc2UiqouctfMoN0B
Tm8SEPxjdw5EI1j8keB7T0Adr3sz461AejbxYfj1qzW9qP500nqWf2UcbDT6u3UZ
kHFnkf1tRgERC8f1DkNjwZqSaPemSwEqWl6/Klt0gOHFM2e4OumBvwN2+rOpoHmZ
pU7ZbB8ML2UDUsAKModTSUd0dGV9horN/FAq/dmSO0jGU6FBOd8QZi9GCiKeKvEv
32h+HRDhIZ8BjHAoJ1B41HvLGqNU8QxTK0095c1NyYc1m/deUSOfTlG+QJiI9gvH
09RLfVQAvggeOWxHabLbkZbt1T++GXVVpARPc40t9Rc3Fx2ktqPhgXYrBi5ODhTw
hJH6Y5WUo07KnmqOZsvA0bC9kuFOe+Wtv87lV9934DrZ7lZGPGMtJ2GE4IU9R5bC
FMJ3y51KFj+vGYINuYD2xoOSove//1g6pACqZ1zhObp1pTQTKO7BxL4ZzaALKcDM
xsUNVqNLxtApVDbmaMkzWaPWEttKYxUhrhwjUcWebQNugUQQS60wEbg7HO/0WT4R
QVHtK5wLZAM3OdN+vn+8zLnKGyyaMEhJokfil1KYoRDa0ZpwiLN3GuhZlC6n3rdL
mTVrg/s1d423dqnK4P0wBv6SVNwT3mvTbi9YzT/B9gGZXANePWAhxekEgzY6MTf6
Es4fSGqdqDz/gGchOJy2I/ADY6CFKbRK+onKs8raXTAlNMnOtlg2G3jIY7cZiPpC
qj943wchygtLWgXbthLhC22B5ZXMztoBEuM/ha+m0b6+PeRzdDMCiqZlk7wrq3in
no5QiPGtE7QMa3qN8Ms75qill2O2yGbFAelf/5c7ij4veo5iIZ/xPzVitDFPS4tx
YJ+OJhxz8bkQ6IJOACn6P304Ov/6BPVxrChpxAVLRThY3eb2sV9Vt07UeOfy02g9
FD65YMCYzkoz6dsSuHDBVq6uKZuXxqOisWh14k3x9t+wzIc81ydfa2VS1BjqD7MY
QolriRvMhL4QrXNk+xWdrwzIepV5YtKwn0WNbkNa4lnikwXUideB56pOMBVd1xtZ
/EvagBxauKvdC4r7KgLSznOehbWMXGpEQ2y3Qid6cR07fhzzw8DV7JVsYuwsQBxX
GotrTAodelsKWHcfKzOu9DHfLDrkGBobe5lOQdEtvxlh3Ww0WHvp8S6/PMQBTnvh
NERHabCH4G6cRGVc7lbnn1VV8duoZVhjkCAidfNd2JZHgAGLOHlqGReYqlfhSav+
LBalPDoSX1s8qd7+KWXQftfZtcUQAWrPGfEG8HIFc/VUVg4Q/mKEZidArbOFK45b
E4NlnYkSzTCZzvdEg1HWLUN3JICAcaBDBNDb+bRjACAx1BobUp2ksMWIqyV6v6Xe
fedydNazigK65tavEagiEPgA5Y+ZMIRM3lHEIlt4xORGKOufY1Sl/bBOXgXmQry6
BSL11yMJ17gKMYnKIZ7oCX0nlQQfuGKeFU0TpGpr5Fo+UoYqHS6QUcxQRu4S7rV+
O7WwU9iSGOQMjxLcOrULuu1NUZwFVUtaRd7VmV1OfwTKjo4ErY7xxFiD86OixoUT
+5Bnx8tUs5Ep0hwkCc1V//DMYvebUDFfIRkChqHoC7XV7jHxOKVs+HFPY0dYOxcW
qmWzUTKdMjaOanCu809nafQ1JVo2IONDrHlCNFTKrBWvv2m57WruirLseLWAIDz5
nnSaC7ERKaz1uJK/aalMhq6af5n5nSIJ75vzGQb7uYVPnMpmk2qWRIk2d6qyXcUg
n5Fbfj35QQ0nXwAOifOAHkgnOHwHAfDRz2sAOhP0W9U=
`protect END_PROTECTED
