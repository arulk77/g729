`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+vI5Yxt0Vw3e+ltQHsWVWcOm7of6sCFeexJ8IhoxAFG
1+nZlWnq8P60XGR2wSpbYk0UWUvgVcHHcmjw5fMpZY/VRCwiEvuJFGgbp3ZPYYxh
3aO9x6RTV3heFGkxLYk+l5RtG+59VSQdLlqCIpeHWjnAb/SwDZGYp/J1ccze6jqO
FGE8p09XbUTPZJsqHN3Am+UW4+BRwjkpWw8bV0kzP7w=
`protect END_PROTECTED
