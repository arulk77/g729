`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFlM8c0OF8m2Wz1xUGCPFYpyTJGyl8yEAE7dYO2OFyPs
ZZt+PZ7/hAAAhS5YkhlTWLoi3t5CPptQkjT7Mp1Hw9XtK/D3pd3GVTaYR9zDrCOF
wnZRcCDanhfKxV1HDaxVckyBQej8NuylNsbEiBHeM4+XSc8/3nEEFHmS7i16QCUm
tM0AdyC4lAhooIirolwa8A==
`protect END_PROTECTED
