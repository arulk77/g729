`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mlFBzCyNIVABC0bhYTMiKxrxVCLY9gVPlXDf7/jAbRDQpWRix5rHFhvG8JH2QCWK
3naYw9b4adUC/vFgq4ShEfyK0MoMAoOl9oObBDc6kwuqQkq26YuxYDm/MzJ+/QiA
B3SDNiVKsfNp88AmqiR+J+wyXT2EbGDBzQW07CeCyKfJP1GzD4icLUCrJV20niyq
yvCzVwTwULjMhOndQLlovlnN1GKNVCSc13XbL4rbuD4eWZyuSUlg45o6bpiaPBzg
`protect END_PROTECTED
