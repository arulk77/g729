`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42we2m5AbqcUi+rRwcTcZCmf1xyv4zxEfaEKZmk7H60A
GiwKlwL0txCafLuKSf2Fsdun1bSyvbG9ZsktOjByfhSokh5yFFzTdmz5wBEbCzIP
PUL1q2nR8yB2zDnXWYxBjfsbOuZMbNYOLboNnKELrNOvbb3RJvfFABM0um4PMkfW
9XHNIXnkq7dPAR5noZSRJrRf/vLrB+hlG2zPXbj1WZnJXsEWwIJsBP9sgzcNtfIM
4lp7UtUyftgwTPXM6Q3htcI83Ywd3pn7Sx9VlyCRCUdXKrp+gIK40farlnRZue3E
V59UZU0I20qufcgxXoVnOpKB6hNT5UZrIoBAmA8iQCzneL5uchKp75lVLsYwKneT
JudUVYxIxZBfeA3Z1XWxJQ==
`protect END_PROTECTED
