`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP5+YyuifJPsRLmQqsWyS/wMsYuoZqtMB1XAkNhpxmXM
CY7AqAWkIIgQv4uUjKKUxSuUCmbxLIkJQC6wEkSg+vRWM46YICS+EYMgjq/J8LSk
acVzEuJVWXuNRQdj4WOVJeVYbCCgRqdraLb7fti6m4Fbo2GJVRRm7183RKbmbo01
CHkY09eZYeWHhoAY03MFAgM5ai0m29F/D8xXO6pvW6wfn0+fGZjUNedhT6U/C++k
8PCwjhxcBHfHe9mhWIaWj1vkTl8WyWI2vtwgKxFImsAiQCJyqesIsB5nceKLYOK3
xDz3XqH/Jz/IPE3UucIXMAs8GqckCNhcQorDQnroWpHU4/KmlBdzV1hRQRHh5nm0
p/LUQGfJJ5fCAHKupSBx1g==
`protect END_PROTECTED
