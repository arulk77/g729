`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xllvNh32353y6ujGD97Z9/LUH1MZ6LoH8e0ryTo9J5t
uMxlCW4Ii9xDFfNgWXL9Fwnw4uRhwfhC0zQ8k9sQ81K61LJD7wuuHK6r34D7+gGR
DDWbnGXzYUDMeaksraCdITNfosJemQAbjk6kjFU9heIK847V4+UEgjF0py+I8PkQ
mtrKSqioAIzFrxawazg8Eombb4ZzjgMa6mfHmCOwr7N+VySNBq3dELOM7DXSTP52
45wKNT8mzU2jkQoa6hFSdIO1GGLoNG1E5Lj+SRHKp/voCJsZI8D1Twi4ucFadhAe
2sT5ChQ2Fti7uTdAxQDs2A==
`protect END_PROTECTED
