`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNx/c/DzzTNJqZQ92yPxeG5Kl4uMOYEzVUsxyc06KIock
bwOZMG2EfMDyt7dDi6lQ/yrW+Dgq1epNv8IidXJX3QDjBh32BSroQvHBd6lqI72M
aV12dNQfngx1QqemfLk5Ay1z/oY4GP1NtjQyt8Od/gB9h4hjojlCTv0HaowAW+DP
BlGSKv0ChQGma1G8J8NcsA6Q25oR16qHp+RI2Wf3Hi0FFQluS9PPj2echeLvlqQb
KIOZPekUgG/8N9CKWNwAYCn7Oed3sOUPDyb8NhuQrx64dUEl0U2X2k9STxk8CeC9
9uSkS88K3RIJUYZbFd3yHg==
`protect END_PROTECTED
