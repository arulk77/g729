`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aWug6iI1EP3XzTeZl3cLnWm92ztgXUs+BtWCfFHNjDTk
9YE5c8zyMP7Mx94ArDi0l6EDcpWC7OxoEKoA9+OXk/mLMZK1pkMgSrtNLzEjdEZT
TJTr7giRm79rzAuBIiNnf5lkWT/65xKsicw3qOByi4uYRClS6OO8K1QSxjMQPmPi
FgXNfpBusqVuTNqygCJa/VPAVpIDWs7H8cXdsQmiDslA234i4w3xiumBi+OpfRXC
VQ5kyjhuKLjtCs+IfMQpO6uHmtqp/IiAq/90npzOOVceA9cl28e7aalKQcDCteCg
a3/ebUkdK8Kv1AjuvyuvGntd9vYSSiRgg/ypCx+uL7kTPil4EP92ogpdr1VPEiTg
PAWBZfWyhLMb8x9gTl+785sgKZwpkcgtWC2axhOvgOluF1pxYFFlVHjdLk2mPJqR
BQr6Pk6wVK0XYfxUQ37D5nvhNcfMW6/gH0DgJr0ayaruWUjOVZkmxGTZ/xEwBxQM
MMqTebPIVQmCafWxBjMRbe51Rj/r+OJMOox5iJqlOOzRSeYGyqM6ILp1lUcg0+QA
TNYFhhFAXogbUPipbfvpjLApnJ5W4h+D5XITYCk+Je7oBzYY5K+/F+WkFLIYCThG
byxRJjTFSICa94A3so2G+qQ36yWFbUcAWTAc5AEa4Dj35RkjczukIGXscEgjKWi9
q81aW/4S4TOi2jP+obuJdZKFZF/y190gx5kwYRUK8E1jj9/HIu9ryMKCSuO0Tcvz
Yl/0hDN1/d/w7fjGuxEfazOVISjf9ssJKSJC2/bLwQLfwVpx0iyny0UJzH+tQ6NG
RtiinQZiMf5LneCO4Vd4Ojroinexc2pbXdr7YQCOOXaVnf6NeC9FJrRQTzbBTQ1y
eMb55bu7MiOiNwMceab6OJ58UQux/W7mT7hpFG5CaM3+2S62pFUbP44bfsple202
ywy7cVg6YgwhjpTGlbcG19xvzaG/Zl+XP4xPuacoi7g5OM7xzgGyNj/qLcm1X2lG
Ub+AbcZL/UYYrcUKyxs7pbeWbuJFueB4hsGQgWPEvnRgBxjWHDQvigT6Q8g5CIAZ
HmTYtmeO3Qh7y9zBfZ60YJ5EUx3J48+A6iZeEGayhboc7wmoXjMHDoIChnCPYbrw
1OvGtONlyXxA0FC4zE3nPaG5Pw/ib7nX6d9w2XuiKBsVg1odmWdFtNWO/nU99Q1W
vpBxBAjzFgqsgl5uxCauu8AOOGEQzSUeDzuRqJiZAApDEEe/ug+vlvT2LQFArfbe
y1oNiUH+1tOkH/fdgW/rng2vm9GykGS17eZgITVPjELDrf5dZXSHXeJIJSCBCI9F
S0iZqckz5gLZLvdxe7SmnPVgw5Zu4LBiMfpRs53Z6rXMBSvcs0DPRtJK9nVNFbPG
oi+qdrI+l2BEFHs+QitGfVz/iNgjJImp4XY60CYrDgYbHDrlOZuCp7c9QVRhbLOE
WMAkLe1nRg/eGcq3gHp+Q/vjdWOcoMHj+2n5LzoX9eT1NSIWnrQKPJOyWOuKHPMl
bgz/4P/jhkAzpxIMv62sI6jBT0FSI2JZeEU36ETct2yHQ2hVzS4FC6IjU2+dF+qI
eObAKx+3a/oZNRhmNwwHIJ8AWuPufrZfIkgxkAp284Ksr8cY5CSlXH7q9rqpW7kU
tDUQ0v6A6x17947qBcLCC8z7Qg7DpzUy0BEin1h8NGgJvWoqrK8NAxcSiSv5tUgX
SZ87OueQGbWXYyspUKTZF3QoARTqL0VDKPvjNrjRvPZlde/k8K7mY0+6YyHxB+/a
+IwuKr8zQIwryv80CqKI6jtuMjXCzmBBiWXFAn+XLTdKCcbwNV6tmKY+NDXbNcNM
KXHWwmu+hcpcDPsKHHHGpwT5Bkr4a7AFKCTPvDexh4qggyxqhs5ptOIMyF+ln8zx
c3tuGS5N+VRPlCWgCPa6otMjxxAVtKCp052v8S/PwGcwvDwootl77xTcf0Rqr5GK
BIefb6s1N680NuJTnEPo8RylyrfqcNoZFEDJ+4peVu71fXPsvQwkpbhf496tCOXz
DtLirgYiu+CpgJ6uINocrmwvO/0aEbVhbkS82x3QG0a/w0+YpQJ0qbL5vDPiEWQ4
OZyN7UNOkw7S5jtHNE3lcjz2xWgEy/G8HETC2vPzRHmPzfeR6jM2iOD9AeFxYIts
KzesdSHF1FzwNgIHxBpvIWdDcWSdx7kOfhh3EPV/8IRv6MtfniTlDVTxTa3cQ8ft
ToL/SJtIVqbFnN/kTb+dB4YB4miAK04AHFe4LU5bI6itb/UZokOevSXosPsazmmq
5aBIpewH0I8FbmUVhG1Wlg9Ii6pktJ5nWrs3tR0bl3XKYn8WZh9gkZGr5kCGIbyQ
4iTWYm4RTioUPi6lYpPo2LlDMNap02uHZCIma5SBVVy0OYgW1wuss5Fmbf8TZOPj
ri2HyQ+lCaxpopyJHdP7ZvvhswSD7/b2jVIAPw0L+zAsa8DH9tkwn/rO7lLyDtu3
P+kdRr16nrG4JHz1iyg9Vvwy3ufbjzqVNkD17fCITvs0F2vQfyCfCWyPSMH64uNT
vhbfJ0fwqRDp7SXuNGnsCRMgkxTGZ4DPQphuY1el69p9Pdy4Y5sj9WhgrkzDIiNk
rI+b7GMOqTpcbxdtZIsFZ+7J9U0RuwmoPKheWKppvtH81NU5vBJ0rtgrp8DfYm20
ESfcIXnHCifLUwZbU93vIsvnVX6YSKillr9nxF3nv/eY6pfLUjJiXJfD0/2+BXY3
tXwDRYMhAKn33VmnsxDMPI87hhmBOZlRBTK1YQt4bLSVCdWK93X39HnZ4ayq0iKf
+qrl72Lgd/cN2MbdTNnp5XFOBc/hbwKmUeCxeeZvJUYk6Iub9UYaV/T2qgPR1cZ9
pXgf0gl6dnGEZ1QX/hecTc3N0HMTUZHCP8a6jqaDr6hlvcIzdFDSyFvsMZg9jWqd
9vtROVYT6D6pluuryNsoWNzWO9k7kQ8HJIn3We+hxYVBd+giJf5isxtyARpTK2Ip
9m70fDd5iRB9y+DVeQIAOCB0McMvdA9zUC7r8NaEUvwkKsRfojQtNR1mj/Y7oQX3
Ros/GrOVPnMUFwEcR2f1GlfjDY0Usz7QOl5gdku/R8oqEoWf5gAKmwzkX0PN7Y5Z
lYUaBlog3wWtOW3lzlqcGjdAFfaX1prWOhSz6wdvnLLOakktlWphxlpKhlSLQ1Od
ZTmA+JSruz8hZHwmop0j1boDmEfy2IOTJySTTp5oNzwmc8z7yPwvijuIL4ZnKvCG
vqK9TUNLVXAIOx81O9PIaghV+1vgootGu7Kp2lDIGkmnxD/9Q0xVM1zq6k06Sr0R
AzIXeCjVGRic87oEWOZzA5APhEIjl5pksCPGfhaZr4HDWjnkslB4/4kEOsx16khl
SPSb+P32shGOKSJVH6BbAi9sX7EWODvlccMlzkoS0E78DJrIEj0C8MHIoqhN0nwE
+zeSIuWs8QZNwYV+ET2SZGocT9L4/r7i1UMdFddprTX0IId6O/u02k79B3PlMA+4
eLj0+Fi6lfexsJsmOyGAr57a8sRzPOB+AOA1H/Si+VeDfX1FzLDPFYC6mEAosBcL
PC6AmVxvslCe4t+Fn5+BgcIOUNz1EYo5wbA88xToe8Bj5ewWVHsyJh2XiTd9Tw8Y
7M9DwzSBMUU8GLKrwGYjPXRiHBLWTPb9sWcs6Ualx0nNgYpEKnUDdpyrlOpqjrgj
CYpB3Sf3qqOd+IIWv15AAU5FOHVjJoenNWCc7vcwLkFLho9Ok9EsbCYYvRZTMQoe
2ww7GG2f6foW4mANx/UGmo5dbfoeLTvM/6ni3WfQotqnPSgxhoGGOjl034ksuL10
zYDzFnOHTIf4a4bqrnBvIoq28tenGYSA4aSIIXd0wkrWqGKZOt5B0bT3Yy5GeLU/
TpqzhMSlUvCI3j7FLvt3KsQ1FALBmWZaFr/+7+mM7G9g3U8D4DyF1mFHcAa3MrNc
0CK7/XEVU9SP8EPuLC0FyPvJ8/h0ncWIQf0fUMnSv/9whx5U/bcHL/+VtxHuDnHW
+CoIOqKsPipaPxkpkgm+L2MD4ZimxC0443OLXoHR2auUJpZlzwV0lOUi08SouUh+
xKc2neiHEAqJ1TATiIsxGeWEl1XslPLisdPwlC/kIi4QL8oL/YFGBZpkGwX3ISDE
p7eQlbG4o35eZbBZutahIf5XcCu8bxiZDxiVuL1+m9LsaB/I5ZP8CaXPJ8L4k3cR
YbWGzBZQ3bkSlo/YoPEo2i7AMzv6QhMXk2u/BduEC2FRrwe7hJmNwiUG6W0SK6as
IWPRY1M0UIdwHmTCr4/xRg==
`protect END_PROTECTED
