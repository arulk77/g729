`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
TfWOfgUmUq6lQBqvo67589uk82Z6OF2JIjlSoyHH/Du7UeyJqnmi3k4RrYa1Siml
A382CQ9iUR98U0laoF9FvmQASuL6zvNnZSvqqyHsZyEeXe4rrrVbttaxT/2fA42U
rA0UmDF6c8yr8k+elVzkjy7KYg3ARfpTvp4foD2heausv0BLvNdCDSQxUsAhO6a/
MGz7N/AU9DQ3ZUvRWgh/jBVSokIa2bQXFfr7GgFV6tD5JlZAG0lvwfhlkOxcBNT9
vggJzkwsw4T+SoQMkvi5bn9eE9xls12bMfufcXHiQgOpGbWGiOCvKX48QK2MLXBZ
DLJHrgv3EKvEUz3UAfsJViFu2NHb/OsgRk9Qk9DNNfwhqUQD8LDeGSeIh2FIBZGA
fOb0V9/nvvxgI2U/7TATVAli/cfKBiYpf86VerJQ06tFeRr6LDDUggUFLxzSYx6q
np/xALgZRWZi52uHYqW/5YEp1Wx4YIOWojXlE1Pzv/6//i0rHtG8Bs0V6ich2wCv
sWNfgxqJGwxREYj+RX6QF4tzosB4Z0bL7WMyArs1u4ALBJLpmiH9DX9IW8zhBypu
PMObc/oTnANPl+lDQnzbC1htEDSaVkqB23tQdv98rTNP6T/4Qgx8iFwgKFUYvFR7
h+YiXj7fnkhh2PxPIXMXaUK8gOxbVcPpiw96QvZ24H/7Z5rBnqjaF/b6CZAKycCg
gZO2CxzyVrmcAseNhlpzDil2RQ396ncmQ5vGB60ja5rN/WMCUxgykZ8iMuU+hPPF
ZGsUSs2jSjuZhFrjyj0wraIRfzck9Pzr+GQtV5G9KZif3GMkO/6eECdMSHWj4DmY
5xRYR450v1ToGJ4wfvC0DcvRIza5sFSqR8LolbRwKAvBbRVggABO6iAyOQgitXUE
iuKT/X5YNr7aGqoB1oaZx75rtcVFqS1uXlI5Q3HKxlZPy9XCxC9dZnf3mDjdy3Ud
jTCoJZ530JLylEsFaOy9fOV5Oj95RUB1/uwnFHijDGIa+RKZKUEroeP/91KE7tz/
2TCN4D+r6WrIQMOYRr+CJ9M/rX8F3uWZ06X16VeSGsSDbrqDR+JtNr6c5TKb2dna
4URshixJM5Ioyg0ExMW44yVRp8DR1YlYTbiuDGXlJCOKbh5l2NAkFPYL/8u56eLw
QGjHg3cpYIKguRqhv4u9bodDhcw4QN/+Vg0YNT4BDYFlW9bifSeceMhrtAo+oAWz
U0xqg9IZNn57wU9dnXIfwnihqpqxmyPeOoezOJmBrz4=
`protect END_PROTECTED
