`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAZH7AJtQK0h8T6siYpK2l0GUNp/S98hqmBXHgiWqogc
D+M0VdD3FAjEMSmIohSewoPL03PAOAfGI/SNPxHzG+AMYVKit+/CYeuG+zCR+4G4
bCmavuLyKH2GBgyOa5wTEULalhOrQWFSMVSuhwDNaCKfWv+bAPiMzSAaOxYfoIoa
GQTMllW+MhjCBfPZO+kCIpLxLQJ1E7ubefMLeiF/rYbdezd2tLcfLTxyGzFhXVmp
lJrUcI5gzohnnulFbiqVUkByAXB7JJiikCmspcP7i1tWvygDb0gYyEETTugRxUpl
s+5ZchGtJjzQV45Yi7vwyplI1LpJ9xOCaOeYvHiNgdbLc/UrutKfB0OVkkN+Smhc
tugyPLoGi7B3YKKyIGnvI/tOs9OZhJWIWKrh9qN98GmYfLIlSK9RKTak9NCJHakh
39zovAQGAbil3fFLqDvQ7Qpj1U8tbr3aUNHa+r9TkIv86QByX2NeOSDT7lyUyfsN
0evxvRTaiQA9ZrY5Nz/uaDLXc9nci+9/bDi8HxIOxtzdZOKsJP5dxL1ETb4v/MQJ
`protect END_PROTECTED
