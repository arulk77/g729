`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePdJjZS3LLNplnriTyojJp3Whw6JF6OOID56ekcg4kWi
YTgHxLrj54dKfY5ODcG67Te0VbCY6OURXymeltzhyuBlx20UwMUC9ahzyF0FVmd7
Hy+vLeioE0c+VCGUyj6HvgnIUepu102kPDgow4IC3+ASSucGPI14cQtLLZC0Y74C
GfpRWX4fwVZ37COaMqqtTJ2D3UjfW+FBsQWg0XNv4t3a19xaU97Tpwfv+j2Kr6T+
xlzWAe6XaV3UBylJR9oMG/13bl/ZYrD9uNRQS0k5cXcVpeY5jrO5ROua9yDzyYu0
b3HB11TXW19tPS/67wMuhAU9kyaMCw09U6mFHxmo+KTuO8xlCFnno/VWIZeS+MFI
kuytdtkYthMedwZ9zXTngAE/6bjSLxBPtNtbvlMiaSYrJtr3pZKU0KRubqN3jtst
`protect END_PROTECTED
