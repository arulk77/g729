`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN22Fmi/Z/KTONfghawplAPflmgJg2M8hWgp6u3U3L/u1
bepmZPRqtVErkpMZ6lxbBbzhSg1DY4QMmjL6Z32zDOiD+WdS60kn662pWHsXvwt7
WMwdJWgM39q+dymjZEsJiktZasLN+t0nP+MPWkQS/iE02Z487TjNZE7GHqzpZNiN
SG+6SVMkZHaistpsfVf1zD7KmChsMmErU4/6GAESlCtLURyV7r+vpf9El5HAHWRL
Y6wE9wD109Q4Z1DRmB3xmIQdYATaBRrQyePKU1yKtg7szB5QgYGGcAkfRSg21K04
GNsbzol5jpRPPj0M2NsiM/g84M64L7m8CqZ5TyyXqHk2JMNqbAHCefXkPEfAx3jw
i4Aorlpeq+p16tp1wvhJLWEgsgYemtpDlcW525fyRBnyDINiTGpTWE2grihzoXO8
vEVj53Bfugwn5mR+xUoLzYNDrSAXOywlWW2YZW+vIhhvgCYZglEKfkUMcO5URJF/
HvdcbZfGRoWE5k3yEs0S4CrnRDsLL1m+U7LHMRsjaaA8Wdb1nvPBF3EczW64Bvzj
hxijnidvbouVOa5fR1E64L7wYl/1S8TFnSNTzvSywvMS/TTKERcYpoXhMzISd+Us
WZrIhKtJr2G2Zf9QRrnrxzkdQ9Hj19Z1Uia5dRlmHysRdmOJOLJ1kMtxRawtPo6C
AXq9ObvPicGXt1IqIkcg8jCpgBt8wtQgu5ZoBtSx0Vi/mpMdgJX6GAuX7+/fm+J/
TVX3zl3EfU9QBHFn4K5bv9tXRh1XHCX9dZ9x4YjtCAhhITKUmQzo7XdLAmEUgHiM
e9w4bEY4SALHI5GMXqGDHfTdSvgu4qOiLwl9YK+eIff39X22c2rVFL5mczG2clZn
tqmMxUlC+aJpbIbIJSrxNp/I33W+NiEkuBnlfOmZ0Nn3k+A/7i7C51HNTntNjaKY
yvvmexU72J76sSndg0jST3TkdnUmMJbEW9p+Om/zY7yVyTf3oIZMsaqbCmtQRl93
swBLjtOyKylJuirtR71Cx7EeR1HbmfI6lruNbMmgDOfk5Lo+9kjXaOjIC4T1mHNS
fdDUYOfe7jlPOp7/JBQr24tsUdw2ZSlHnZRXlsZJnlUgjaBPQ0msOe0ykxXNdVaC
x6g04l6ZjIw66n/+XaybOCIBrNVG2vcr7pX5Wn7+i+38Huc1y4stlgxIMjJoMF5O
k2ErUYhbyaVgJ2itzKERvtjhm151EPQDZr75q4FEhGJV4smYYwFH5uYyDDIVZn1u
CZGVzubNnBVdBA/XCt86yBWaMieXQlFjT5NrmHXz4akr6jePKx8dH24XYRmP9CY7
NqoRaga18L0mNzPA6vQRMOGX7k+MrNkmxTVKRCb0Q+CWhnMqiJWGuOnCdWKZ8xuT
YJlVXfVNqUYgvvLrJJZqi2npCpTWxT2IA2yYm1pGBVTdOb/Cet8GyrspBX7Tx1i0
YSmLz5di5uuZvREOEK6ixxN5/yBn+mGYxSvVogK1mFxJMXjNjSyaxjjXvdM+8UIY
t6yZjTdWDdW0BmegViDCgMquC7KViOoXWzBMIdQNjGu6IsHkprawnrtEuimeTxTr
lzLucl8lrC6BklIZ9dgfH1Z2ch4QKWDysiXozJSZcaP05qOJ5o0xtXtiESEcRhzT
`protect END_PROTECTED
