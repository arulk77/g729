`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bFIQbJQHTJr6UL3+OMm7ol8WVgZIIMdhkn086Dk/u284585ksOnkz3SbFpm+wdcf
r5VFH3lCrULbXkWrkTZ2nmHfuMcNJLhISzESwFSEiS+E2xxt+D6PHrOez3TziLsA
mCkoTjxYlHBjiqC4/U6ww8e/XAD03Lh3tkzzQJWBRGUC9tCpKBt/nfes9SnoLMj+
AvHDAF0jqWcPrEt+nKz1bwNDEIRHXBlER+7Cf4Mbo/0=
`protect END_PROTECTED
