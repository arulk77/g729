`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
iC/ZEDsOAt5W/x/VrHQOdd7o1ujlJqTxb/RSv/moRUwAwtunDCjsUOYJbBO9pCS5
XETwhrl+Cfes2sNoh8Xck5di6wnlVpzPSh49xDgUezchtEzzgiELz8xtVDBFrZL6
SAmWiEszpw606Lhb2oDELKXfS5aucTCe5YDbjOCjTlgXggXQ2AQ0wtvH7Wpo7sl7
60o11fFl49Qr3ir3mokX25nt0im5HshihJCCQWrWxdfeaQvdk908UUyyqc+mnL29
4H+V1sv/m35Pig0XETjzDOF/gKBSEhHN1t3eSRHhl6cXlwkXaoiAl4wIsxaB7vgg
liAn9UqsMBVLAs2OckJFFH6psa8aOktyn3F1wNx4SJDthdU0vSbG2CeDeZOG3u1U
WmvSJFqTM5VkYEB1V8btdPmnRWNtqN0ZOv1VE1WOlAxH3qMKArkSlbs0JTRLM1Ht
TZ7Cp3Fc8Ue0ncWjuqu2XvnEYHLduCcEEHYjCqc8Cf0H86FtDoPvA5/eNE99rjAW
YdaDZl9MQbQ782t0VX6VEdPBgqgWvks3RZkdhQD45gUuq+9arRx9EUiJOGQF6Fzf
TghtTZJOYSy852+OeA7rhDZF2Zk+oXz7oiFj+gtpngd3eenwYdPGNngqC7dWRNHQ
iFK79nNheoK+NeiS1ebx+ONJRBeheN7ztRDtnBw7VaQjtvm4rKYvvTjIxszO/kYb
txDilZDVRkkEErAAuQehcGyY1MXOJYKmvenU2mlA0HQ2zMtK79Pwn8U/KkXwKqcU
5HbPbC2hD8xTVsJQQZZhFfQx7ORYh0YzeLQf8q+jGSolnXOkW7uAx83jTc4GOJcv
XLHHpl1mzl2Y+gdNq4bGhsU2/3l83STgz3j0tCbzDtX7svU5D8yekmj741Ajcx+3
zZpQoH9oVA2SrbZmgR1iB0XP+Bhx6vTuYsvnvKdlf9FOfXUCHpgTHKKw1b0r6h1t
0kA9xweXUe5ZcKox98xZWa9gLipj1uzHU5OweINGnw0EWzkPwXC5nGW0IW5tivFn
EdNf8bEkVClma5a/bm9gV+3zzaotMAmAc0g0kxz2NlMBZkfLrAxLm1aLkEytnbN+
fHw9gf1S9UM5We5fpSP0h65Y9TtyypE3BsV8mGBSC/WWOoJBxvFJdKjeu8tmS4YR
BpLwbc2+ixix9LkENPsIJ4Z3seUgDTYc6ZmLbCI6jJI=
`protect END_PROTECTED
