`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxka4pR2Y9H69rDt8VwBKC/ZnBrKFpwcukA+u3ixWwVp2t
bS2/dvw1ORJVWQe8zSk+3q0C2w0hiLynVfsXbCyM0qP8wc2UslJChexsEyXjI9ra
luBOYll1RYzwReDMi8/Da7PuSJf4zW3K0fwgv0gxNXfTy8qNIsH0R4XerV4SBzTP
S575bWJVrkkXpwjAHzGG9aF8JJM9lPXOrWzno+gH37lPZL/+hhkdOxDukUCBgdWx
A/ke7Vhv47iUQuJWCSWpf0cWRQjhLk5OKkeaNBQL2/giZf2huezvUxU8BcqBeKm6
v1rDu8+jqNExCt61KPuKCR7hqUHG9QBh6ojUsQbrzodCA9R4YV0KkcZ83YlPA4y/
5t5B0BWC+GXilMc/2xn736QDmF5EjfjqJek5a94bI58MpeG7YL7/Rw9tRejRwhCJ
qKYGMVyO29fLV1slJJsBydNKfxgZO2C+Lki9ZfuCaHtQnUtJmPPlWOPbXMA+e4Bu
iEK1HuKQPEMax8UBvYMIotMP7/0oeAFrGiFni97zX4SKfHPz4X9HHuYahEpax5Uh
KMI+dRHKFtuoy4bKmk8yZeB1xpP10jsqSe7Mefs6Zw+jxQG2EQSLZ3rlCAJrTHej
tDvp1Fe52lQFgTyEmACiZykfNpuIEMF94kzvzdAer/JDd12UYk702j9FAGxdzKse
QcYIY7zlHo//lTSjBjYS6ECvnPoDkXbCh14H5m8yLKWZNmVDesAQ16mSi0FJ8pfF
wayxtQjN9ourgkI3F4rOQKveVFlCGUSHsDJi/9mugjsWMTwBPeqC0su6MkTW2+mG
hPZeUmUKIvh66ihqknAJIspqowsOGk1b2zHcmtdciHw=
`protect END_PROTECTED
