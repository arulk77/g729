`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JS6Ee/OUguv3S0KjECptSJn620YlyMi5Y7mU+v9yIGVvKRHZbXqKtHKVZttjIoKH
eHt+J3cEr7EBhPsyTPIYVx4aPaHL80KlqQTMSUh5anGYj2hH0+Sku3b/KMdriuJW
8k4Artuzv+t5xbOBaDZWFexC692iRBfY/DHJQuYD3aKxnNcBS0TUjLfcZcvmxWVA
Z24BFkO1aK9GURLbe9NeFMUkFsNBolnawHnus6IWbFbFqqdZcJ2T7ItHnI03nU0u
HaCfOpD8YWlcb0QHcaSof83T7Vqt9HDDPnCOo//1S2tvMX/QwagAVVZ0fg4E4Kd6
1hJJsv/yvwHRWsdEA0HPzVswESn7/esXg9Plix3x8F1CXKWk2jfsDMgEZoWLLPWT
FVO3sPWB6gAo0UbNblevAOLWnlEvp/PYEH1RP7OuSbk=
`protect END_PROTECTED
