`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+A8VTXuiauOxLqgjSxWbsUTT56YQ/iA3RGiVklWiobn
xHWRF9kaaVPgjz75YAYC0IG9uK/u5O/hO/vttitbA0xiRUkJL1j6tvNirHH0NYc8
7xdXla8gOd0hq04b8hzGPWfVrg+bfbD+IK9SxkgRCcL1RQaFSXMN4h281yy3e8Ma
R5WSYhOAeNJlZhP0cqKg+1jX/LtzBUHmq1MUmoq+2y9PdTkZi31MyyxNgkdgVQLE
uJUeXN1LzgKKm4LWB6WIa1/qe6k1OH6BS+3eGiGNrAE=
`protect END_PROTECTED
