`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wLQfvnzBkr/eG0VlK1FYBy+ZnVPGDGSSADstD4CT3uW
JBh+EyTxtCBtU2dlOv3Jnu8Ty07buliwSI3xnIZ0ZJjttbTFJrTVDTcqa75Vbsp8
rNC4VBjQWMNykPwlQAcpu0KGFkIrndiOFXgCd7q3Vwo4OXmm1XBi2FA3heIpOHOg
A4tbgDqrfsiEYsqQFxWBr+/9Vq1tGBELXI+vGoU94as=
`protect END_PROTECTED
