`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4z29cENYRZLgU6JMlNZsunkjPJP+40XKE8784IHXbT5s
B1kQ/e1VrrSmaljvEa1kVjpw3kdy7VtfyyU3syi7v2Ve2EArdYFIaDQpgnueCnTJ
q0shKzPfASwwf2YxxSD2byjwvn2eH74pY1/Vr0vZbUIsYutrdfCojStnKQAWiCZ9
70gbWe5WkaWcCytBh5T0qXSJMrd6XPc0dPBOpOjpCLA1aVR60xqYmHidnn+frL/v
WTb88fkbOgcWKnl3P+VZzEMN3hcGORZ8sM0E/thdqERb63rlSWUVqPB861pwFOD3
st0InVfJ/2ILaoXclP5giw==
`protect END_PROTECTED
