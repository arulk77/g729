`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
OEANfVc+r/Wi/slF7DX7FKltw+uXLHcmTqCgCakVy1pqWqxN+ReSVk4/wZjf3xnF
MxH706jqvwsV77HRYUtQaHQCxsJmrmyk4UxwQVOJlU3SUAmGPfQjrY/zNL9vCAEO
yl7slQYZqT1fjaV5pV9jG5GtIWYSuRQpffjLLHv9mfwIi7agf+aD3plyLb97cPFi
lygeSVgZ5I0ACD/pWm9aDHbuuxkHjxHaYLOKDufO9fUc7DQ2VstFS6d+FUV7hpQz
h7NJT3guuOu7lGk3p/ObfvAAv+M/9V+7gah2ZEC0/xa8Y/fA76eK5MIuHwV4dydI
bSmasN64/CdYq5KexcYXmahx3+9dF85R5ZbiRtLUyDghcjHVLHmwbxavbO9dLGVw
QLa6Ih7c9XYug2jkFzn4e3BJucamERebmE4Pr/qL0G5C2LDPtIVwSlp6mJaoAFGo
HGr+bm2oS7GFFiKDMXwRZvfHIvZJF96DB+e7FvwoYsWPMDxu9RytX7QuwlJMQUKn
mW/X5mIxfXtANOmRwpdzSfie0P4HYfKXzUVnuRAFXL130jV1AAJGmVHfewHNF29C
8B51UQ0m9ILZTyB4J6TA7PcP4/DHVun9NKgslQMHxt5YxAK9x3xXQf8ieBqz98xt
xcsddOzA1yKovYdouLrJPDsGG5vsWG63FWYm/pmitk8LUt98VGolR6JFHh3I2dXN
I/waFv1YxccyZq/K/y4j9A6ouXfjowIMkBMzEkheu29QiO1y1asa8wcBjJCa62p1
BbH/p4WFEhBNJGioh82WzDrnGq/n3MsBqFgO1JiIB162FyX4KcRkQkpT8ZYIyVWN
hAzxEYhyBnSMiOM8jPlQ5UHhf84ke/pkuQYTtF5N5SRFEULRea7Q+XNMKdyNDaP6
34zzYyLAXQY/pN7/BXpFWaJdiayHB3J4bU5CNJ1yuikuOXD4Q72fKoPJgXnFvhth
W0/pDsZyCWVpSsS0cZRkuThVEzTfzhFm/sCfN3A+UCrOvfDW5eKoZgZqdcyux7Zr
JpERUQ/BhCL25rsYQNt/zXqX4ABPiwJW6e2b7CmFRPNJZtHfYOVXZzk6BwL8/pjK
4qpIw7ojmaAszZ1+iiPuC5wRPm8O/USSnYrW3WhyOU7zFJP6GAU0TlCJ0kRMTC+F
VjQmwasDHcvf79HCtTzbWDy29c6Q0R+abFVEEcJt4N090eJBnEg3wSdT/o+lMSJ4
lLN5XNJEx7Ibcjh4r1ci6wDjZPAjsg4YDObQCDko2Yzep+V6nhvHUHgih6Dy6wm/
1gV2CWam4PTnP86KGEVz7mXRjruU2hjI58ZwxnOg0CP1Qs6rjnmIgGkJsxyRqze2
JaVCjWmVwTg2mAqzVSTIk7aOZ6fHakpxKiXM0Q185iK291++yCw/aDt/akn9CBf8
0hfH8cL+8fba9lo+p0R5dhm5L1ISdPGVLCG4BjieExXi8k08mzg6iJyXf/x3K9TY
9+UB4lWb4PH3uCxJuFd6WugFr6Nigtjp2gwvfHVd2yk=
`protect END_PROTECTED
