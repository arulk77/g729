`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
sCN6e8c8VyI48RAejMrT9RddYJNZhtKDO/PP/MHJC5l4JmoBchwyYZHhOQpMt7GU
qqzkHqu830BoikimhnGRgOfqlO8/O+j3v8Exts4bUoeRJRDGznFVrSHVnEfRWxSH
3EgfQqNSm5z3AK1iMCmSTmbki6y6YIzZcCij4+p0ezF1Al7sa+lGKt8sOpaBYuqM
PL4ZsLHVvM6G9b3tLgX9+T97M0nWfzi+1MRga9+ONqsRsGhyAn6KIGsu/fUOZPYm
NbFBuQNh+BCuJtNBAw6pSa/4Bd+dTbglAkb7p6n/gLk=
`protect END_PROTECTED
