`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJj9+jJS7HkJTLd+iNn+4opokcmkqOzgQdAk7aLRZ75E
n8RQ6lFBZd7uctVJ/IqXHjjtZZGHSa7U2cf0xdacW8I37MN8W17W0HhXszwIpM74
YU5AQwcFtYIibiKocArr5VjvOdPkQn/Ehvvst2xuipE58Vn0CD1BgMjXqcatlZsh
xMBTEXGkF6DgFLfbNPG3oIvIELYqRUubLed+y+nDJMeCcNP3LtwQIAAmRPmlUN3V
`protect END_PROTECTED
