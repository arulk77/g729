`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDDeaVNPCwwQYN8usb6f4js9UHVL6VKdaaJIcq4MW+Pw
OP7WJ5Tmm/isRIRZ0Ms+C8LmnhouyylzLc2mxzZ0a9U/B4MfVsi+mjb11e6ihS+X
8Ri8AR/1EX60Kr3azRUNp2My8t3Qq/mk3kO4FWN21fU7MjDJSZQxd8tkJJyL2k78
D8g0djMwPYLzTL7MBTmjag==
`protect END_PROTECTED
