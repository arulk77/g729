`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJnxw5NT6Fv7zcqS8YmWg2Kh4JS+ZVAAezAmHkekTGR7
AgACm8x9N0frJvFzcD+rFkKKikOjx/Td+u+T/S9ylB3sFPvvjvrkMv1ON59EM/pB
HezBoECD+hwWMszFmIMmcbShXuaAfEf3S1f6l3d57cz2aUBN0csVbLY/B9CefbcX
jodgSoLUF62upLrXNsKQ7h3nQQ5eaVrfPlbf5JHZZ+Y=
`protect END_PROTECTED
