`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zFx8Ns/IiHSIUvWpiLRWHOLOgwrP+he8n3USaW1kdzW
Zuw5Chu/O1lB48t9MQF5DKHbl7veLKlsY1++LaSQ0sIj6Q1/KnT3k+PzX/EFILuK
HxESC83tFRSpM4qfwtPKl8Gh3lxSViYSJuW7f+QWUUcQj/Dg+CWehUF3kGWelv+M
S6gA/TkfBU2O3C08Xi/bB9Tcw92SLkS0dxmMZdStJvQbiKsmRRZabk6tAfXMgz2F
TUNeYqf7Y1axsVrdL4sHQOekwgu5uscRfXzJyY6tyA4KAEWInnO3HOY2+L2V08L5
FX1tOL4VBAp6mpTb3lLidQ==
`protect END_PROTECTED
