`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD3WwL6pJwiSxCrR8/xgnGmml3xa/7mpwXaW18iA+N3W
ZaogJNwsR1TCp7U4ZNkJdfa7v8NbmzuB5BR2QIo+7jK5bK1bY2twxLVx5vapgWB8
TKE9VQ8GkTcPtgtJ13D9RUS1EbCMxBE2rfE28Hs/iQPCI3csEvkaR7vDIpQirZ5I
5ZScsujQ/2nlZ+JqVkz1lw==
`protect END_PROTECTED
