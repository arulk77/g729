`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Oc+KV2tPx2QJ4Fp/h3/bhKgo9YqqY9vPpWJldIeuuXAbFXw9h3d76Tl9Lo3B4tu2
YgWqbw8ikMkrM7rEhqynvUESkm9h8Dji0Fac67891+GCHf4/mMqAnbjeAxgDS+lP
LY602j1PYyzfK61JWYs5zlvyoOi8DAHf9S3h+qoGRvXCvsiML/9hsaddR1sUT4Ff
KpmRJ9w8r4aS6lcy6pKXV80v4xd7zzU3Zrt60R9sUOj6+k8IQjliAlf2KOYQ9SkJ
`protect END_PROTECTED
