`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMzzlFSN6QUGA9kD0EKyzfLY/p+5LcfAhAF/QtrJBicJ
zGAzxMmEsvOIPJFA2voPAdIAZqZ217w/ge1uILjFWHNBDOSf+jLG56OhmO9I52kv
6XGrK0HKu9uttbrrPCXJvJEQRO31fhaQ53wwekAzbxk+d4P6gGBoHF4VoPmg5aA9
Ja69lDZDucaMq1zuBXzQR/Kk1W4YpfGDr4H+WvWAxbImFpMdw7yblUFO4OhgRhF+
0JEKT/NcyP2Tlz8HSCVJTkySqSJpBLS9vc6UMyBjaLL0KTvr4kOtkaFkUpE33MND
gu6mPVEdlhwd51AIWUTNehMST5cZBe0KUjVtcmLRaC0h2HJ4fq03t+k0WYlA+0wY
Lzvx7AOE6DnkN2bJMAscc+waWfv7++4EVurd9PRcB3MswNW+ltKk2ZQn+Cd05BBJ
o5rsExCcPE6U75n1W29zyukXS9VOm6iqtJ9zBNGY+7okUg3BGcxGuX3i5jJyv6pT
pgkQAGyNx+4IT6YYg8Jxdjg80hs7/aV/48O0mMFu4G9g2peZIVaKcLawTPQuFoTx
`protect END_PROTECTED
