`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zI9pD/BoCq0ZWHlMkmKcZ2j8Z++QawfcO09fWWdsKFo
k/5cDaXjN5U3FdgwzsVfB+5JxBtWfh/RoyKpUBmXbd3OdH2xWMICs/PEa/MZ2/mg
3StbQIpkBdRJRM22fM8nRJ3AyjEf0W6QfozWT8AXm7A5MkgEJMVuLD9+xb/KyxFL
Z1sd2qYjeCBb66aenYLg/1qKvGBWy8SGwhtkfmxxhJ5jNMuGIyulUBc2VnW0KfD9
ZtyiFKUHv9oIDgMjhPJJo9v8ekrM5NOEy9BJi2ENelQmiR7OnvB3v+hHoh3nqy+4
Sr18QoHEt1xpZXENUbnfcJrMW4TcUPX30Cqdj7HcBQ+6jWbKmkW2TRgeuY0YExO7
OY656wHZ6e5dn3HGq+Td87ExL+joifNoa/YfuMBv+xytiPwj6W+f1R0dofMfAcRR
qDbIPUMmmgrf0u7kAAr1yg==
`protect END_PROTECTED
