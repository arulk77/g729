`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBds+11OAwD4il0Dki6nLga+xWjOSKt+ht7yBSzSoACX
+QLhu8+301WUnwD335n3OaEs3ASMZy8jgCYqNdZNlfoLTPzPMw+vrpljaXAPSklT
wWgGsaVGMGQphR/dNWU5qdffRdUPrUgQ0Bdw0ajN5AgJoIYpJt8Sr6PcCeIKRbao
RYVxnw5KUx6Fs6wrj1yTF1QJr0SNckd0/n9bCUDJXHWyqfLU7KSa3yAKrmtbspPG
DaNB2s8D86G+W3RT8pelIvkiLsC7L2Xx0EHugNs7dLyvbIwpIEZgmhHISNcw8A9F
ltTQ6/JSaw5GD9E1E4K4n+FJi24KyFPbtmJwgPVDbWOa8df+laBl1XXY9d0cv8h2
C8FKZUCVTdVLQAjaWh2l49sY2IsGwtDoSxBpkN+7dbfZcdplhiYsID8keB/8vwNQ
9P71VT1RhTAVChhxI/0C7Buxa9igJONHu7NDxeSOOrjqgKB46xPxcKlO5qmZEiHy
0bfmHUruWTuxwq3RKUhFicI73QoQuUi1RxbW8KSBp2eYcsIjyrvuB9W/BGQjvIyn
`protect END_PROTECTED
