`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKedzQw+WLIODasq440PhZ937f1CTfb1oNuO878LkTdI
KALto16knuOHxm0wiJR7jaE0jnAlAfUEXYKAyM91HPf6+lC7/oCMFfzpsX3bln/e
O4h93Ba7q1w+BiQxkroqJenuuS7tMPcN8lqPGV9uSt0xcXXP1X164w1TD1/KRAwq
0u5WjiwibCmNtiLGBsiOAviE+2SZ+B43kJQz2P636OF3sanCr7GkU7GsiUi6rFjf
x1VBaqWX7VUNM8qQLnqBwKTGgOtIWUT+6e+lKii7r5woNdhy7/5Wf6rVae/N7VY4
0zikhE7f8NRxWw8S3BEBIIM3SuKeUwfNRzd6RXXnIDptJRqkdyakE2oygcxjBv3B
U0KEzhf/XuRec+FXBUVH3A==
`protect END_PROTECTED
