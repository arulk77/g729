`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFPtpblNstlCzC2MhiCM8prbyYOjvKhZteADqBlj7AoS
3wLmmSL7rgvj9W2u2Q3u0L6SQjhbGXn2jjBj1jfTT7E88qLtqV0O0R/JUK5mGmlp
niiBJ1b/np7XSpB7l4F9LqQfblwwI4rjrp4uDLlxVkp8w17WdRPbGFxyger/6AH2
7iIclfyCqAfCyHVdYM4odWKE70AvcE0e6FYJDilfjxOYu2kP+Fqxdn/xojT/pS18
uz+sQDgrLd+fh0EGpr6+PZrQqxJ/OwCB1d11r2crh2Q3n46HemKQULM1A3SVYt1t
OzB10TEa7i8Uw8V2gsQtCYF3gTYyQ2BOWr+1s8r0XmBk7sWUZ/5BFB+1JPsJDr5F
ip6FxO2cAmc3vvUI7kq09pCrjSaZJD5F5PcnBT9RF21oebfgaSFyR59518kDirQY
yLjk0FYFLohyNErIIyj3gAlB/KM21LrVuvzOZ2wACHb46beMx1Mb/t1/PrisOOK8
FGO60LRgjmv+3DCeP2CfkgW8UWXYM1ytFAE5NGNBRukcboE7qtTH2dXHx57qugHa
7m1FcdpHIGpm5FRqUlJC4tQnUE+r5LRN6+q4fsKbfPTBAgGyjyz2YJQr4LdAJdbw
ihDxoIrBcSLwt7MPRUvt4Y+7RuYHF6f9wGeF/E5WT5SqBoKrMMBd+9819c8/t69k
dad1YGT0V1/N+9sxzk/OPjMlm72syRPIN8Z++eqcN0DikHFB0+wW+A4vk8BT1/hE
8hba2CN3ZVg3GVheic6E1oIC/9V27Agxb8l8wUJK+jm5g4ErRO5Sp5NVZCCL1EBs
0+VwBX+3SFLIDfpF1tVdiKveRywHAVC8kQKJql5om4Y=
`protect END_PROTECTED
