`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Acz3EXNnfgrlrBmqQuR8UR2ZuFiqXJsO+5Yfusg0qL5icTSSWbuLIYgQ4XQWi36q
k2H8GlSNI0YIS1dxKqUQANuxBmqSt/+z0XX4CyQ+7stHAFPtUdi0z3TDbAIbeypx
+w0Pk2X5gm8XLEuRcMsba/48xY2LFK0EkAA2tAeDF4S+bRlgVmpM+NpffHDB7rdG
e4b3Fa4AhHaT23f7HX4ga9zaaOiUwAbrOsu4qImrVPxuZqXmGBUoD9xy7WQ6Udhl
DW3mkCXMMM1jE9+1/GmnlifpUU7k+WEtNWuhxmDlSmrGsMuKDSp6afasLgiA8UvE
p3sAkvVfSt7Jm46VmPDpkhFU/HKKgUByBzFNga8STfs=
`protect END_PROTECTED
