`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDytfJxUegZ7ywRBV72PhaXgZIIas1400Cmgh1ZZXk5a
pediHwMdfXDwZysIV0IDSiKlTO8z6iEL2IZTXXQJakd64YyynfcmSyXuOYYo851h
/Ub7Rcenb7a4GL1V2tqbnaZTnlNEUqk9bf8A3wMVpzQsFk5KiESDUFckNIqeeh1o
1i3wgPVdheVgJaNIrBPptt2WTqcs518CyxYWzZcnNEWUrsazUodSfJYwjxUIR9GG
Plqc5XRx2teKqzzXCGoA7VMZ783wtDizDZVP0USOSeDcxJIDNSlTtyXJfiVb1+vk
In0ZZSA5vKrRyntqgLSAWmL0K1uIuKdyS9LPnmHUCq6XcDAm1PRO1VruB2pBsn30
`protect END_PROTECTED
