`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+wR5rXzOuYxViSQxmewkdlZqYo3mW6d03udtlrD4+K9
o6T4xbDCA4vcxHs5bZFuw82OHg2pINPJyPjhQCJh1JxRRIO0gsE4if1HoWZj1J4f
0QFJkxA8ooZaoU7EMyJPJdjkaVdIaHKb/YmT1hvlARDQED1qvPmIas0qMBPgyhm8
g7dP7W3FRl5vJ5L6JKvnxOQ/4kGsC9mQLPqRlmhvzPTPVXo3Q9iPewkOLignhPSv
Ur6mAy1DIGuse3d2iDtXa6HOzldM1fc3SSxSh8V538SgmxnL/bM6RN2opK//AtX1
JJlJ0PKciMrgywZdG95ybg==
`protect END_PROTECTED
