`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGav7fpspAH/bMKtUidtCBOs62Xe7Cwpf0dStqLG/GBP
iYM29YuVf7kczCWP+KAW+JNXcI3h8ory7+Nk9e+6CDiZpPSXHKFVS+DSZYs53PpU
g86qdpUIYSwAqtzg9PTQKEeRlS40Nkp/+Uv26w4/XJi02UAQ00dsCFNd4mh7SZb8
iOSHYH92atkyk8/OZ7UsNNyI4t7lkY+HBG3rao1ReILF4yMqiJbketZOfTvPZNEL
`protect END_PROTECTED
