`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
jNB3A/SDPdw1qqBZEKwWo3xBX+WrwjAOPddLvLXkLfosjdActN1dgBwKUMvTU5sO
raJzHFYS+DObWl8jHSpVIW7Lo4EAaZlB1DEOfM3tPmRqtSkodbj1nZK1hSrKyrSu
itvPKJDV6++LLWUW5+Eic/LQqyS8PCvQntK36Mo8dKgAPkaVl/02r4UWIyBM6hkd
Ne4BJAx6NWjpg6u973GbevAq4XnfcJ5re4Rpf7Sdvvpo8mJrDfHYxrO7/bAsgTzI
uy87lC4k9+2dxeKaVKPxTrQ+0nYxLD2GXJhfcboXUiIIoy0vhauQ2NOTqpxGDJuQ
NnlpDmx7vhzy4yz6CbPV4iYZSBFufdknA8VTuW0Ih99EDw0OEIdpXAHrLt+DiWQz
8EsIwe2iSDG5DoDg/PCr9MaVhLV82ODsjTS9p/RRWxuF9zjv2QGYzTa6TGXOqu27
ow8MAFQ6VZR+o5TLwVwr3g==
`protect END_PROTECTED
