`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47s5rdBGsTibUgxXL9rO/2KWaO+YeLiREkX57JAdjUsv
qjcjWKMuiHr3HI6bbZ1Hz1PLJVKcRljIeM6LHQ4W2OQVbK/58HmmTIkqxF5JQak6
FJzoFPrk9cX1jAbYdy+pA7JyiYmk92OD0BJVPFPZF+jrdm1eZS6qX6MUTziqR3cX
YHudMbse83l/XcbvGg9uvBGZYqj7olQD65Kg1fZUnek=
`protect END_PROTECTED
