`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFE6WCzUw9E6In+Zjxnue2QEmSKcEUCcg9Zs/4O1iDP3
JppW5W13/hWyrg1EZdTWOVDT+D4iLfsDQMx1R3c6MkzLh6dS6nVqTPQT3ImmpAW3
+AlnZ/cCt9dK9geSyJrg9ZOtgyNwPK5X0A5QqHjxyVAGKeVw6D6cxLMSPygL5gNW
fBOW3dtjBc8g662/Y3zyCFIL2aNsYNet5AH6lEzDrEZNg2I221/o9N88XWCSug7Z
JEl8nP9xxxD1OCelHOZNGxnl5Jl7Q8fvY4VRKImcQj+7jf86RP3zuw1fVHIBJGCl
MdszSS2d3lqsSdt7Bjucs1QDWorizeZgrTqSSXn1ewLvNCRJUfgSlTRr9tW5w96q
xicQB0Fv3vdO6P112s12u7c9XcGpzcLXnpOmlTvgEWmA1ydldkY/nOKsCFrM1u5X
WVtwLlDhrkmXoyjx52ZIJc1xMBVpFbmKUEsRvj0UpObzWSS0R94yQGCyEUQVkP/w
PqZNZP7/pGLn42zXaGkr38GwIk7e0TKUx2F+fjXkpvkWOExPYMFsM1qVO8WBrqfJ
`protect END_PROTECTED
