`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBrLFXgOkX4UFW7bUj0Kw5Wq5b0XF5zPWYuRD9De2q0J
hRHkAGxtwPU6bZtS4gPHp4ke11bBWI8IbrkhACnrqp1GiMaxUVBQtYPWU3F6Ky95
wlvSIgC931sx5PRPZeVlQk2/t2cS4mccDdXvzPrn8ivmEkxc958HPnl3UAG9AdZF
2Kk/pjXbpSbj4LKV4h+hAePmIBhpb+1vHfu/NmnfCOhgjW9cxAPFBKl5HFrpzZVQ
c7XkIn5bUx7iKqwKOD5qjefxeHjT225A/5gwKMqWpZfQWCoqcvpnlM4zGsgs+ChU
LqWjBciOQEeJ1s7iweE8BI9ZC2qaHvp/PX/bcjZg/Il748YXc4Bk4lclvipovp1F
anns/BgzKRiDlVNt8NnLah/ZOT2f9CP06JUkq3p/l/uaq5BsHTkl2/1Fpsdr7Sji
m4DfkYf0lI7zg4PFs8uglyJtWPSzXQrcpqYNfYMuqWXmVeN+TZJ40K1eM2yb2JOb
ZylEoFHnxQ3znt+utFtgXOZuYpEiwB2LCBcmaUalJJ6Yp9rCjd7Zi+db+NOezXWo
FKageQ5c1lX/o2Nv3aQf7BMyRktZPFXMD+tcczvtMBo2RY9Bag88l9mklZ+T1ROu
MEyVSE4VxCm6hAV6cc7MVTVaGpVBACuyBC5AAczSlK3A+MR3H7vA/Gus1AjxVkqV
QaRXAfZOCOagag9UXAcyjhTSHv1/fQyhmX+69rBzCtL7XiGoavzuGK3LyV1qF7NR
cxrKwcuIE4vbydJGifpIRErjLXL9n/mBh5mEr3ZI3v/mkxZjqg1wkb4A9kZG7huA
qANus4pOj/4w0gbKzAKVQWBUP76k8th3e5+bPrdfGUall9z3Pk16aVgzaEc/AvpS
/vZ6/glX4tjQJA424wp5ith4yXjgI32NCtSpfcQfeMg3y2cVjbzmVryXUbDFy8ip
XCLiIgB3YdWitjbFmN39B+SjTLO5fVYKptnxe8vorCqcrbVWnHnXDP2uB5t1ffnW
7u0WkOGZeKxW1TJCZBZt+6FuaH4BUivMUkkPML/AiC30J8g9+ChXJBwD3gD3ghGz
Sl/KUae7IPmo6+46sfbM+BSPfMpJCy0LwNgaD2Cjifs=
`protect END_PROTECTED
