`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePv9vpAkazHbhMgQ/HoCnInKHZaIfqw7nh5vhernT59n
ji9foF/xs0S6/wxIF+gFBy67gGXx6+HAmhYttx8n1ol6rutTqHyRlu5ITAXZv1v+
GpZRwywmhKNdiPO/W+fFeNX6Ltpq0KkMxsvevYjOeRfHJ3FQidzeKpnJD3PVLj7g
EtxAMUc0FxdrrE61HuqXcZTW/j0hzxZeyrYWsgSSap9BrXFR+GZS5RGPJAszkuSj
lY2k+rWvGvBj1MO6/9wfj2k8CyRsP/34CjaDw2zTCeRnMJ+rbqhlGOZmesWRZtx3
nFld2ZhCN8KTEoPrP8o04KjF3ky/gXkSxN/9kbY2rnFHmrl4UwS92m+k4AXp3kCd
4CZeuJXxB5GiRAo2B/aIj3x/WKkcpjrzN46VDFgUBR+Kc6R5aQ51lqdYsYAUeCQM
`protect END_PROTECTED
