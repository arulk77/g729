`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNz6ku0cgBt2hhivtGerXP2ogJ/UaTH9PVA40NVpt0Yn
hwtGF7begiE/R15kbtmCfo2bKY94SMNcGN+o78R8vP5bYNvHmIKMTUxaP7Oolzea
5AhrGSOsoDonZS+SiScWDYBncvmA4D+/CScKYmnhnY0Br9tm+wcqMizr1s9Ept/s
OV3K6pGnfMZnZehNLGmDsAKkYnOz6UlNMvXykjZGi4ZyECLsHI+oAoVTcZtKBkRC
YRQQIw9AqBIjTRixZpFdNOVRYxQT+VqxQL/10O2kBWI+N5ZIyHoSAJV/K03282wO
G4ogtf+HujqfZzpod4IccA==
`protect END_PROTECTED
