`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Ii/UvEg8W9+Gr3uKAWBLspPrbjVa3jp9vIvPZMKne0ZDXpkugOeqJAilJVw6GN8s
XEb4vdj9/3w37he1bEg0dw1QDzaKKSAnl/aVV0NvMG484Y9CJGsYkkd8r0Yedow5
ntttmdxshLGt2Cn2DCrho+x0xZbKzJJjzp5XDkZcT9yRSJ49ssffLQtqxYBOrcGP
scsSEJhZNq42zcMvUuiEYHbsJAXsHR+OaxvPoOd5kMw=
`protect END_PROTECTED
