`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJiB1jic7dCLvRmH6vfsAwMwhmjHW85r0iIiN6lP9aL3
HRGEDfiZcgw7nfJwa1p9PH+S2Js3G6NuELbZJkgZ/jidYF3uAqGT7cR7kz0Lapu5
rH+6xp3Cxubh+SLwGOF0aVzmRFgH6VOJKIy3Ag78tSGekmZdP5dOB9ut7VzFJYbF
HHmJUsxYtpiypepGephbL+j2otagIr/vfOLXJZg1/I5tu3d234wqnnGAWrDsbaSK
kJ1bmweWcpsqm4NOFZ/amfxhYOX0ouJOUlqc8y66cAIAovYQQHX4jFU5ZmcwOZyB
SuoKoEsYArSqT5sKb1ZHXZSsQNm881HKtjWseqRsUcMmPbAljkHedlBT4Zv7exTA
IXm2LdS9hq3qSGsZZpgdD9FJYba6X/yfvm7SybB91x+2bL0UwSPF4Cr9OD7IeOZN
5zZKODtuH1alw8Kek39Yds6Dp4DG5nIbnZEzh2a+JSiH4xwHPPct+bBddZp4tuDK
sgMnG8hCxricIaCpyGRZCqjRX6zekg/u5eHMskH8K4LbPltkJ6Iq++91zS8sg7on
P2BaaMQeZkl8iY/EXAC2tLFkah7MOqv45vQT/MPtuFM=
`protect END_PROTECTED
