`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
EcnZZ02XIZVXOn7vElj2Xl7LcGlOHTCfbuXBIashFPhp0Zmt05Y/ncCDWNrLobBS
Hjj5oKoSxOEs0+3QjSsiofYNx7fGYjGSYmaIKd8rGEAO5HQeAWX3Nsx3P8FfVoq9
HmYivHFy6HjKrX0bB4cITsJNgfqYFM6G7YkIxV50I4AOZtNWOF499AD4KhS60XiJ
iQvlZLAY8Dt6VPWIALKBt56Zd5qrxYAFO9D8Q0GjQkAhpVB5z59wHUbx14n0agO6
dQNd0EvQkDdVHTxileIGVty0xYGj633jrp6UlkX3Fm4MKjeOYzx3gV+3vU1Gk1lP
IK7iS/YEUA5JucWHF9vo3/jFAqGZjkT/beaAUXHrY8grrvBIaphJSEMl4eCNXEwT
8Ztwm87H7M0ira+YbBfhJCedI3skhdsH3yFLvRMAh5v6dzpcfdzyfup3eL0bLtQE
S5ywNQxSK6hBB2zXndRwOmy0F/zY63BiBzexFwPkC52NwRMDsGClhioxgHtsTWxy
uu+KXYjiHpaV0mq2zNMkf+BeHMCSRgh0HoKVHZYNpk5V4t9OxapOVhmX+eWQ6IT7
oenJrgrl4Y471pLZIK8fdA==
`protect END_PROTECTED
