`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu486Y41qgPdHVWYnelMZzZUpyK30hrWaAdtSrdYn1ji6Z
eFAvFFbmCeO0LHphcryWECcpZUUrDmJ5RPqJw9SnsjZwyL9PMU1m2ns+KA7wXyLi
HaI9Px34eOe7EXLRdtjlh52JP/51VCZgSLkqmDLxJCy+ZxnwY9D56CURJdtvLtAG
+Z9doviX/3/8433AV2NpLa+1Yf7fLhjz90GGqswheap4TxTLJGALDmtAP+WVW6J4
I300pRLkv5/UTJNUw04k56A0S2uVY+rrNg+MgPbZekeUZOp+KFbBVchU9wBkr7U/
q4o09kOjAycPqOekolC1bg==
`protect END_PROTECTED
