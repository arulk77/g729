`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41UoIQwmQLX4bIm+fsv4UT5n+tlFnVgwoC8ypxsGvfxq
fYzI8MIIRl6hX0jzB5SWQugvVmM1W9B1n6C/66D1Uq9hgyL0GwWUOB1cRqLA8LFp
R0XCiyVemqsOJs04p45Ols0FKqlSfQOUJXia4tHshTFcYPJqeKJvY1aAwHVwUeSg
SaAHTmNk5c3yjpc5gMSzf7760rEHb7vF/862pvQySo3kfl4lFJAa4WlcaawaMml0
dmwvG/S9zoya5wwZYRmHW5ZKtmiIylp/XM89cF5+kjAKnWIH2mRlVTRc/gXuF9hG
2OJZEG8Kdp2Eln43XtQiEk3ln1SkieR17zn70YBRhEPAYjLH4pP5Bb+pEo07jl8r
Tx3xUebxRMdvRWC159pP+Pjdvqhfoud/6heoSPi+R/ibxj+eKPXcxtW0lrfncFqg
RqGEcjTAKWZyNVWbQmFD4jWb7DVBlYUjZhsrq7K1PnPcYDsG02PKZX4Mr2bOSxW6
W8LsK/eK0aPQUpe5eRsw65XzK85hlrO5O/n3s+T3IXtJhMUdPGN9EQwoBMMqr2/E
/YKbX9whV9f3BlVH0So7wQWg27H9XmUiVVcbfKFAAmCa1fPq41apK7Apbs8puO/i
fCHd67HcWS3P7HwE0k3YPB0W1UyShsJ6B4SQrKuvtY9Teodkdr2p22Sj4xDu2OEt
pawXBqyGHIE135EsX7KPhPR9azHJkZam4vuUMNKRuRJl8bP7/kx64Y3MUDyT7OLX
ghuz5ATARyaLqFH9O9ugTdxV+tYOuRlA+9H8gDcRkoRoI440n0qsfNqtg3XlHIPK
MjEFbMTJTqEpDWIWoAeos+QhOBZzkG4OxR/xKLA2qFsWGwXyCkI2+Cg//SJbAsu1
waGUZpuMFLtZc5j/zC0W4PCIYVQqeWEJ5iXXToPof1iLyTNUypsjlJYCBIXnuP3g
wpBX56zfmujcH4PphyvfcCN9mWTAO7vnDaa3p+QnU8NpfA4Kw0TIBEy13McpFwN1
SgwKVeclsBI6X2VQ2mpIjrXAhaRdLl2hqwvVpTe7WS5HpyR25zFMF09qo3wkqgqm
KZbWJkCJDYzsg+EyxS+5c0Ih8pD6AncV5dnQ2zL6j8ZL6g6eEKP57tLZyTTOw/w3
7JrSzYs/5hvqZyaoQ2eIy8MVzBgT+WwGmxOdy1DTzLJQxzFKuW+JNlgQcJQGL4Cq
B3N+KNvV/At10F56/VjbdRgEkjkNNdip8tY3zjlyWz6GIziiXR7omIA/jvfFuKiU
uLurmhuQ5e4O5baNrijGVd2ygAkA6vW9Pwl4A+WsDgqNqY3I7X+jqNeM5kvI3Wzy
DyZF3IG64SYuGQqlAyFnET+Zj1uy+8SK88bWIySjWn+2r1b4ACCHLoIheIP9OBLQ
DqW9XQ0RUa0/FKSTH2mYsiquIf9OqWWwwH2lvkqCV6YSOHvgrWWKWsO/IyEOeRF7
uJIqr32CzzDDQ3BnZ2GZefrrnCKL54Y4oSQOO6TOvnTjdQZ+mPHDIrupEP9wupYm
ErPBn3jJohO0tGa1YNGO6CBviq8ZCAurQ3N4Z61109mcCdfNgib/Q778U5OLbrV/
6RS1zYGlb7t4dsDgppbv6evL2nDnzfbBcE0qWg2ZS+i2SZZqAk60bXx4F4RZtuLC
FMnVkm7CZIqxYnC0AA6kuT0QEpSvcUxNm7ajr7CidrmqgmVOFnFWLFMVrUacpD+3
tuRvzSAGKxhcNFzVI3IQUkP//QpNdgOqt9GLyi0GwU1FLvW/Vzda/GBNxHIQVxa6
MGnuKAbsVh197JUYg+u0iUhtg0e97e5Luxx/5kqTgJ66imQx+enZmWqu553JJMh4
YBEiR43khgOvtc5QDDh2Sf1NtvHyoWtyXGDqmPqTMeSBJ14N6xLrSR20/pt5377f
mErluRJnB4pO6HYzZ7Fu5CpndDz4PBkUrHdvYYE4l0PxQxC1d2J28zRXWxljXvAY
i+7qexCcMXQ80pBWpdJVUuORnJ6/7AUDLw9B9QHJxf7F2svLaF8f8EI5BImJThTg
/pA3mlx8B7zYJlNiv4LoyQp91NZQhOgQSG7wOwKyY+OB4kah7fpTsT/US3hhuNEd
USvdfu8HrFAaOxHOum8x3IHpG2FnIiYS2dthQFE8euhMXk+rbeHJwQL7pmVXE2bv
IKejuUiIV+/vNeghV52SykA3r3T6GcZV4XhfMGj3YM/8R0n3kNonicQCAbS8esn8
njl0xj51dPVEuHBs/M4yzxPVO3gIE+0OOlId6n/WkgdM4reVEPmrm6qAKTq6LmFj
HRk/bbgN3/4EBOQJ3vkw0weu2QaTL50tErh6jarXICjO1WyZcvoJ2iJvN+jpK501
Ccjg2xsGSQlKNKm6y4fhVYugiQPMEixoYrieB04yMp0iJzOJTppVKEgtRRgK3/TK
opluwsPzRt9tm/qssGkjcHleiZTliD034ilwNRrEElcdsyeAjrd7ey0YYKE7eDDd
wLrNLGXlftn5jnBsHAGFH2zJEiZrMamDo9+qlIhhlijanr9ffDeXExy1GdSlTJY/
ANR0OP3fP2Q97ql9BF3wrxY2ayW/sCZCvQUMkbyz2bfLkuybCRVVEcsBH/iFwtmi
ui/Xc2O4o1Fv3WIR4Bllzfb//XU/rx/LwXK8vntgcIeU1AEeQEX4ogXzxAOcvGp3
lzv21z3FkZNnR7iQAttrfZuEOX/6RhnG9kqTxjG35bFZjrzqK9Bb5CWOQIEKkHjn
irEe+4LLDI0u9C8AofWbwPKwimkmJhmnGz4F38DwgXpQOTldMPcv/cBUr8UUVD17
dOYtwBq4hHK4HqGguT//cvFEwae8YD+HZ1Mx5SfN/lo6SB5HnTVVHiWK2aHEhLrX
vQL9hmSZkZ1g11XjYv5BMzm9X2noMKju++l65WexFpqliaoW2o5QhPMI/jY8J4ZA
fuHlqX47YKZvHpsk1zkC2A==
`protect END_PROTECTED
