`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aR07FFMhkD/J6FC14cs8HpaVYvfvwTp9gTlBkLQQS18D
UtiNsEEPUYBaN5ZTPDVpAM9lmdh3vON/+kBqN5woDm7/6XCq5IOvxQllUEXR9ba5
fkF9HlGaLH0IyTiif2YZ/SbDiDX9FdTRuQZ284trfvHNBOGiBakjyPlJWvuMRI6O
tMcsneklnCe+WZzR/c0al17KL1fS2e2GyYY83BpSn+9U8M6j3lceY7cZzqHQp+8p
oeuv4m6XNkRAYHjnhkBt0EyzOn7mdg3mYqETrGIBQfAvIaet21NMf9SLSuSUo77N
m6gCN1wlcJzDlaagsjlW1tbZbrn09ehvHbFJ1/ysSpJ2he1gOfIgB9u7FmiFNTBV
p+4elsYAs9qz6orutgERTl7CUsu7E+SleYJ7uIMqGowotGoLJGsaM+arIw334bpY
7VvPpMJXw0RllAKYA0R/CHL3TMdu7hP/p0+Rx0dUF6ivToSw6x/5dubPF2LQOvJ+
d3H8xtGbFMoHsLPamXBw23Mqd3GmdHDuTrZDbK2XY2zCSpYBZEz9QCr+g5kdX8Z1
Sm9n6fF6Nc8EFWywlKWtj0YcQSOwQfQc1kFHkF/iEwxPqR0yBwOXdp93lfRPJ/ne
+FWNE2HtxlDiVrQF5aplEcEVVbdc23rwKNWY7NqMnuSQuTzXcwkaj3WCnFuiNc3Q
4uCYEQst0POlRi6pQGPN621dUBFtkw9B8ZiGA7FjJSD40+eHexpOfvcDzykdnIfO
KvRldRu4rv40N9MZhevykwS6acfbvEwxwI+lavaaSlZkFF/Q/EwBO3FpQFfRDEVc
/rrK3KAAzt4zIklrWkktOA==
`protect END_PROTECTED
