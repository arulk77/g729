`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAYVPZkHbV2Wj/Ke6PD6QiJdvxZDkAtWqb/ImVP37Ak+i
BNPktLGwDrI5ITVJHRMafODy7ConwbkqYaPjA+3uO9km+pU0Cr6DRIvXb3v/Z2gD
31/hNL0mYxAKD9+pMc/YldKCew40MrrihIIQjz6vS4Y1W89aWcoD2+K1tFakdKQM
Nn+PXELsM/+b819ZqHhrNovj7hhnvhmEWt55mOc7gmSlbOZ4Gj1De/ANQM+sZ0Zh
Ci0WUyURI5LMSRcQGmPEybd+3paGJ9hE5dlVZqbkY9GHATnTpfIvN77O+vv9ibrJ
vmLmcmil+kel+vHNLfUWAl5mID/++WMR090GzuVxyjvrfSoifY412CKacTwHk6C/
c7aOxSOTSCskVV7hsYpn/Ox6aTfeNeM3kUBHBn/HzUsb8KvqXBUBmgkKa4hil+yd
meFvBawXxT98Iznl3jcvc210icu6sZe+Pv6y0cGZwUY+JwcDG5UvIUbvJy7K88zj
1TZ34IGWQRs8A2BrHgJhJCtI8O37Kf7z/vuhh8KUUme6WuIxqJeu6quH7wVsqntD
ZHqB46PN9qa9R2fmgu+rck7C4dBxahipuROi6UPQjl0vkUhixJVSnWmOiuj8SnSe
qje81J4sO5nTm5rv/7BUymAQ65vznlkZ2ZsSNiivF5NVQC+X9NiKycltvWR0SoTC
sJgxK+A57h17BgF5ggy945zUIUZDI1BYSygr7wdpacZ2xBAU8IIuIG/28WEUTRHp
QqpfOqsw0xY5GGqW4u6DhH19w7I4Bc774xDwM0KHp2V5G7tyiNqlt3oJEfbXiMSH
ySI6k7rWb5WmeJ8nYeQ6bO+w3OSlYc3FINqrthMCwpVJ76KVq08qYDd6NOMVhqvW
LrU2AAmHKXhViDeBF/S3bIs5ab0vE2g8A6eQFoyHqqykOlsYVkmzz9SAyiYfNvVI
yli7cI79GieAm+rX8b3hbBjqdLx9E3PFC49rYVBNEl5yhOoUFDJIDzvKFTbMEV4x
eniJOfg8Pg8Udrf9cF0MDAdOHoekQOMZA+9EC9DjgFQTKfykFxQCQ/xwL6GrzbA/
/xURW3qCCI1O1HgV9BNDvM9svYECNwl6mHE5l5IfnuevhaGXAGU3lBREBYC/uchM
8veaqpCnM/ffF0ZCfb6fsGXjg4KaUN8n6g1pU1URxCnDVVh0tpZA3SmDyaWRgoni
hcTaCuG4uvrOaCgRENvbTnhB/WCvWY0VL4yH5EK0P+dSOaz96mC/NV7B6lcjxGb8
KX8Alk/zCxsSGOb+1d9bOh+S8oZzgFlZvaubnKl9OxuJlEFx3GEADm5zg5sSblXG
R5ZXLKnshFYP7YAtuIppA22G9g0J0qMA9EiOJBLmebdksQxuP5/XX7N+oxe9YrSe
xqHzrcc3tdnIWBny0CEjiMDsFlEBze718N+pMVnbbRt+D6GtnwSKJFHDJVBkNSt1
wbBL8kZ0qUVYSeeJ19iV0TY1j2tnpkYBxcQ0x5LRQzlVpcfBkv8rjFE9sFl5e4Ga
FiiP5YDHIXoJ/8uOUmoRQkUBqbAnQA4d8C4mbfIM59qVugAy9oIbNTT0L6BV27Q0
+/W9LFeF4KoE1f46ygJMAitwyePbUQMlcUWKp2Uce8QLSg20NFd7Qq53vadcN8+4
rzEjqTcT9/RBsQ92coOzF8UR7b2aXg+SLecXCe2o15KVt/OFCk3DW1zvIDozczuK
VxYGa3xHBGeDqL5m8ymgMbGEYauzjkBIqRdnwOrKZ//5+vkI+WxICUjLBsWJ7bQf
RGhanr+GMks5+PXJNYAQ4UJszXuQY/tE/8CAvRLhenL5Uwv7XpYlqmYimW7sJb9D
nizVInwOSWJlNohI56tvxiZzZJX+KEIE7l+qM7NLCaY80LjngSkyfCgCPG65YFVg
fx56C8ouZBBHfU2oPoQ9O0qOUBVg7sOujwjjLWIqN9gIBqxKMZAFVHtq/VkVzJVn
ukbBn4zYP+8RRuQo5ETNtgeBadQBlFHYWd4CzmCmLVfrOaYUDLF3cZiazXN9zbYu
+C6hq7KQPpg+4o38gL2Al87wZNWG1mYo++Zljk0ixD49u6/IMVt7z88KFd1LnQQF
a0CifCQIT7ui7RjN8gqa2CwTGozF23+pnx8FXXOBlsxld3g7WPYhVde9AKm2fJ1V
ePcvgAjOE6V/OQJOOh6LbsdBF8G+vljQZvnxCL2h5ErJOVh8w7b/s/aGDw5SXmSY
MQ6HJYLSlgrtC66d6YhkMDJ7F9ss4mehI51EOrATmEyvct8xie5OrS927KN7hgws
yPW8fUuklvJ/gKOWF6/vecg0IvX8EUk96/YtBmbZvYi38OQ/iKegaj3SrEz9G3v0
Ct7bCdpLuTiRY9rvPcwz0K4uH5SqoElmXEIevn88xyQ6Cxg0T0ZlDboRwiWwwVV+
GudpRzStpVNvYxMwx66c6k4Ulk0xIDmbahti/Uuy/om6r/B5m5LPDgyqfcXPo4eO
a9TcErrMT8RzY61Gsk24phFGYOnUDmupsI7AirN9eMZaN1GEaphCqQLYm5us6luY
Izfv0bwlEFYFWdLMAHV/H7upxrdZfZI7YIaRJkqoojwMw0DDvq8jGgsH6LLuE9dn
iuiqnrr70z77IQ/TsjSTQaWzp1HYpf3CrXnnQ9rv6hRNwSmfNEJVlmT5mGr8FTeM
a/2t6T9GVJeX37u3Gt3OEgvUV2bm7/UrY6dyLvYiEVeoEIGU4KPKCLq7dbOPyQxJ
hIRLQNvY04DLbTR6fGbrXw/D7T3r0/VSinFWK2vkHje/ZWYd6ht7TkSH/dDrdgoo
84p0OqlNfAAP7RhkvRcwMmXTy7f/TcDqpXkueEViZD9DsLgVFzzzcfAgKzn7x117
sAUGV0mcs0e7+4ITbbQdsu7Vw6O1w9vu9AN6i2VI3duqGeCW0kznZkIks7qpJ8jL
KnOYGIgUAoJzdmHwUspN9R+V+5i5+HiHCnE5ibVH//XGcoT2M9aHZnZKpK44AEfo
U4vUzoIdRLX++ao1i8U+K6B+5AHDyJjXCBrUf4h7zXA+KKcZGwm1AnA9fToDy5HF
a1T82vGbSd33qmh117bvt4oxKO3IKsBiWgNXrldE01865GfcRcnXok6DNuxsn/hk
IGSegsLOoMhJYFppHIS2yBg0cSB7RTPH9i4pBJBeguO/m+XCkR89xan/tvUMunuE
1jRWxKKSs9/sOMabNkhKWqokcMct5vgf5M2GjLgzavt1lWNUw7pQj31XNLJLY7VW
ONIc3OCp57EJ9TFYJSVGiOD5N4U0neeqvUSaPndLTR37SEfbrY6+1pbUN50JHIn1
9G5w+zNVX+WyvHE2E7WWGQKNUaOhBa482AllcksZCgRzDCi8G9kBZK6qPJAjXUzl
E7LLFFgY2edizX8ZMb7/qTQQHiu/Ipu7NwULpdbgggY7wyh49miAkgd2gty/7ixw
GJ42AL2jzAcw81jurkiFP+LdFC3oNdRp1Xrww1Z3k/WyM9Q1Uawz8bNTjOBTlq/U
czUD1wvc3QTKnK8L6r3HVVGFTdjUSolYUhqAAdLXp5CLi+uycBK66SzJfUuMLcLR
7LbsaY2JLQQyzG2SwxF4zA==
`protect END_PROTECTED
