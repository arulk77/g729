`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFQBAo08sp6mCTElmCUjMWDVyT9jY6vSGhU1FKiS8I52
5/P4DBbphAHHJvBpGX6ckjH3MmmIVqDDdxCx1Sw3AqO2UI0iitQWUyMh+IvTnrMD
RtaC8zQKLEbE+v/Hhcqxh1cutqlnn4XUSP/7LdL+/ZMYoxWj+igXVz6tjjySJZlM
Y2eeZKVc3Zx+PZLbv3P3o+ORDch/EJRmmn344MtLNx61hF1VavIlIoVgp34N5oMO
UIseFRKd/LDzPG8LcZW0IjnqZceHopuM9eJZMQ0CKICn0xRPw+DemJ+AQxsGp84R
TAz90oJYGa+k/Rc74giNFTnHitzfj3OhSYx3m03BKMtdzI3lkoSxoFYOATYLaxkm
MO3R7Ty9NiT9AHW3S2Cho/b0QioTNfMG5xBVaUqNSXVwrDZPVWw9TookhPeHJ+YE
zikzNyw9vnU/TWo8byr7g/lH9/kuUt6URgebbvQzZco1iyXXoWleYCdtq2zRvEgl
jTVpX2pLuJ7sV3cnEO2avLt+digESacVn45pV08eysxDdnbkSGdNsON2hoNL39l0
gD+mP0d7p33stsKhFo7Hzzar017H5/dWS7XjoWwfNupgvZ8Xjr540Uy2ueSD+yD8
8lb8OwIF2kOfU1PLfZH9JARW+e2iTRVpVRJculuhgfRCTjNaMmcxokCrL8b77Nnm
OZXklvsb/fqyzXH5DsscndVaYmqpW20y/L2ZesMISl5GKZEWOc73smeZC8FmkzPm
RdbdneQC/v6MLhgtkncuPvBy824gPyHumC9hcsTu6gIznKivzhQxk1XDJTXQZTKE
`protect END_PROTECTED
