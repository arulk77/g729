`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45KLHu9QI3+UnafMmOlBxw+T+60vDIvZSgAn15NAjlua
1pSfaVhTk6zGr1NSQXgYjOwVatAgzYWn0F8OUQjEJryGlcQXnkO6fmKZhDZgce4S
KNGTnRsSfWjnJTKsBjA2Gcs56DUTVFG8YeO0AhOQssDDzAUml9yXMbsuZqSU3WF7
daprT/JBaNhuAPC+DO06ImX7Rx1jKIrk4DLWign1Fte4agyQ6KtNl4uAHuFLAIl4
CNExuOxLOWq0nY8nnQgceUl8dfEgjZFgbOKzz75egl0S0rTa64EE7J075iXg7TPx
RKGcDSlaOgLr4BiOi+2vWQ==
`protect END_PROTECTED
