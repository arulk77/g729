`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN6ePoYNsfg+rN2nnIxssztHhue+WkKSsul9ruypldt5o
JZnw5mpHTGBVZUdN8vhq+Y5hCDOFBGUR5h5I/EnCqD5WAN3i1tcXq0hJ1E2aDcP+
KGm1FZE4C9Cr/5dEKJKjtrCHMeeVzH1g8Ho4EdO07jK0xkZ3l8kzKK/GusnPFOcE
Q+Df1GPZU3LG0IRpZjnQ95ChfJlwc55jerhIsbqBUE6PAkT67C2ujoMetkCDPsDt
e8m7bwz66/ru32As3M7Za6I83HCnXSNIyjiepSu99/kuN90Md41H2GHdCFR3EQQl
g5Aahz1mTxqw7fBTaFbfYH7aRJZgnriqpTAunpbQWmKCRt1cWVjPzFiB0JcDIDKC
vjF2PhcMzmD64z8K/G+Oag27gHJFh5zuLFQrblaC74mTZDOsXSBRFgfAM2bwlS8G
2bTzcKTeysocVwAWTZBrzi28oIaJ8RVXUigPYPaumYIQl0UGDA7i5J7g2QtWKzYw
n1+UJxxeVLNBnP1X3oO10wTIdEMjTR6CYBWjJsOLp45QUb5TVfzY067EqxhUe6YD
XA4OZa9UR3cg4St6ZJ4bDumUM4JZs6TgXfepa4Esgg9/B6vNtF9jb4a+uBDIAyAQ
OTOhQFVAa663JPwH2I5c32oLpWSUDac1Lg2t0SdYt11I8aX9w6cOnGxmRYsmVvqX
iWMUAbmceM4f0Kj3Aq/PZJ1KEVMzuvmMquKMoO+bIaQ8FWg86XHpFiZig2Q35QtU
qUvySz66liFlWtOc/ABkuUxggqz8FU0bwICHhMJiIqInCC8PRwQtden8bsYiXzxL
8/lISuN/dq8q0MNoSCZEPwuA/HqTGl7gsMj2R4/ualfLCaXNARiiF07hT4ss9+AC
w88Jy8x969G4Gfrr5O+qYzlLeSHaqYyEcE2OTFjn9VdajUy0qwi8DIcP5JOjqc8l
YixTq38jN/EgrnOYd8WEQaNvAu8xLt0MpEUeLRDRE73cbMz+5HbLeTnm07CBwqfi
nbmN3ob7u+8i4FaOHoqFo+l0aJhPZSQ9Fsnv3pW5umj/hgnV6LP65pTRQE1K86vS
YDX0GZe441T7VhVjcDRc+YtwpYMYx5xj3MveDzkaoIgtdLSPmldpnBbGpGRaXDzk
4G2uK/l9DiBJ47S+lZtKDrM0FqVqDJ9dCyqdgM+ngAC5UVBBxMnHCBMkQJUdwPE/
Uwm9I8feQ17CEfQXNVAPNpxP09A3PwsOFyLonmnU1bY/xzs56VKzsRAEpoOrome7
fxRY3ciAzsMq16rnHOtFrl90j+CdF8lva3hdjEqEMl8XZd7jJ/RBw4VXlAm1kxHS
Cek36Uwyxe72CKpxgv4J7/1Tt+7H8RF6OKbQdkOdk9B4lGUQpz/h7u1aKnQg6JLk
OVB3HUjpYnl9eUK2ERDZ3DLiVUKqDeZcOy919EoZ89mhysVvaQzoGLHxOd9Yf1+N
GIY3Gku4BUFHb1BC+NWJXHx0QOUqj6vcwBuVKaijuOeAlZAokxuz5R+YCAMdgvqS
aKp6c8Ka88VawGx3UhzCMl9jn7Xyhm1nkyM7FPtUboKHTN3Yakp2+1Yf6Vd2pR4n
duXhktH7Dajbo0zJs7fVxnyezydK+kWJLImbw8kHgU3iG6lf/8a9CNnrW6RWputO
sTKC3slWnddKRlt6AKmrznWCL1CiK7VWeNVC/zO/Emev15ZWw5hMMifUgpeEM5x8
cFCjrxqwCZ40XGyiVsfEROX9i0gKpRd5W0MuCt1Vorf9e7ghjYB8OpReqjGHo+wq
YoQq1Ii7I+Z7kFTc3tSRqcO7jBvk27eRHUFGJVCX/GT3rR/yf83WC3AvVnzmt+z4
rNnMiEUsenszKCwClGdvCWKnnH7Wl/ANFZTsgE29EPzpnTgqvz9YDUOCZxJeoMIo
g9U9ISMFZx6RQHj0mL9RFsW9c0hLZtjgJ9hA3zIVEUqhMqC52JnYKDiCSs2Zmt0S
prF0wPyErkzVXQpYx1Z5dh9t/qHb9HdhZmo1Nts7pCOIsGZgLxxoaU48R/V7IZyc
nJTztnWduitUEEtvAF/HJEdqqdYRg9VexyTI3H8Y21Cg4ba9iTS5ows3nfZ7SLZy
NDJrNyb4OI5VvhPCGAqXZLwEJLpTP+u28P5g2i1ZKiAPlNYUMctnpqljyotmuNp6
VvInUPQr/xii/ecvaqp7uV1bvgaFaAz2cltc518Abyzmqxe4GwACV5Qbm+qE70f+
+eU3xbY4r51fh1NL77cx4uV0rLpsG6E/ER/SserpJWhCWWe9AOcyhmu/h1oJwF0K
wjhNHCFc0q+BxNEY5845JTHEILycmkakoW1M6syIy1CHliiG733d6ArvQO+bSP3G
jLALMNyGlEqToniunjsOoagU7pNSQQy6o5qu9yPsO7lVjffxdgKimPrV+yZAfzyD
WtfnteTmStyvHxuvCi5+6TjqDoUmrUKLW4QBjoZDRCoxPoYkrhGqWbdeaLeyMzw+
pOWBonQ2Wvu1o9icatfDuknhyR0dBk8VDUpNfOsU7SIOzWhBiHj8zYlDl7BL/d0V
MslRLbbP0/KDwGZ3VORH1MLpAEDd3uIyiT5kp7bEqrhLbg7eV3OALKKk39SvkjOu
vTiPEYXo3Qj5TOoj3CX8yUNnwYm7TTJDA2bkAD07E2zWxswqfNKkmTL5Wy61VMdb
ncol5in0k/TOEeKQmX594era7YbNHtIYVdi196tvDL8UUQyVBDTnJM2duMNxpZIf
6T+rH/nB668ZM3Hxo2N4aDeNG8iJi1jXs1ehVXeDIdItm033KMcwfJw0q/L27oZ1
FDWG8n0VgeXtPPP5RHpPX9GPXUu+RbPhTAgPuR7ZsDzWn5quRiESl3u7rWgW5ttQ
Oik3rDsCcsDx0fJ3qb62VaWpUUOuY4QlJEMp9d4vWbpvzexzu5LmfvD5WRYQH0sJ
iirNaFQz2vS05IAvOUuEOxo2a/uNkm+U4cMIii4G/6kExL285Y5cwf9QRWkADltg
bdNEE3SREDEmolL9YUR6qdpafkTYKoyCURTSOqPOs+FGvk5KISEOWrjKywN194ph
WbVaVYByWacZLc+Hk03J5DZ2F2/HuztFieWzFSbvZTyICeVu9p+zXCMTqyBmmC7k
344md60P8w0RPA/KV2RrbPUDMfMuKx+tnj+Uerre+KCgwRMV4p4tPOzBJHze++MK
k/AOLpvxdO9llKCncId9/SjwIqdhLJKaLpQ0nhFE7SSm1tzQTJm0s8tcesWTmmNf
xnAQzmj8B1Ya7BvCseWh1bxszLW7EaPkbnrumbYRMnPVNwsA6wPtRQsIv+k78fpi
QZkru83+SibBnp439/i3cePJpI4peDleTN3EsREcu4ML5zm2iMXGGrLuhW+VQxoA
2sqlwZAajV5OMoakCxsicfwrZUXa8l+IfrXwBCk8U0S55ta3MoUcV/eclzAnJcRg
QA+/D0bhUHvrNyy3uOMvsHFuTjm+/O3HVN//8knSa18HWnOU6UqLWLwy5A8ic//m
FXcuGJsNiPMp0ukwiu7MPrO9j9U0dbI7AwIG521C4G0g/QT06vizAw8p1SMY8AHt
Ejj01rY+LwtOiba5R8oF4pDvp0i7k6vvj+90cpCCK06X3ymkoTnJtlo5OXi9o1Uh
0XAcSizxhUhZuGTeHOSZZq0t0a0Z3qSByc8G4gVBsKSZFfVNCA69gJCDLeNkqy3w
0FnEyszR0Fe7n6IcBenG7ElHwLge4JS0hiOtN3LyLgE5CUshopc25GGufbutGYDt
4ZDMT6WsS9kKKHl0/RcHcIXipN4GwMeVGLgNYgJCL9oFRfJO/M4aPDS29CHzxNdU
SMNL8cQs3e8vkhtkm82aVZCoYcdrT88NlkLtxqC9QrwG3rKrJOHaH0Z1vHuMFpnD
zrGnQoaWDZLVg/ogAdzvnznFLO6o+Y+yDEZZhoDpJFvC3gdszxfRpJaqCl+Kd5Mx
CkuYafUc06MMs1KG3vc6n80lT53gkhaw1iclGC9PiKWjNgWhN7vqdjUEqoyvYH1o
YqBd7HSFZnr/CkCDk9wGpDa4pY0T5Ni/pBX1Hv7Vidzhx/NiWAmZ/sBXFMGx2dxG
94u0z6Gsf7kEm7f1gEGaWPi2Vhf/ZaOShJn7e4KUJ2f6FZKmNVOejNNjlhIYuboB
fpsF54UJU20Z41Fa50UsURu8IS5fKWHXh2Yz+MQ/cytFXSlDGaKSufu5Dham2lZi
bm8ixU8QBbH5E/4KWOwpcW0L2iZwnmC4P7DLF4eb0b1HM+HIAhVje6KETbOQR2B/
OI9LjJb7HemTXgldMRpmYtBUaYM+oxJihBYnXDawEJt3MQZ+yJERiMPWr+WbU5dm
1ZVAicnOHg5iWmp50rG/3L4ZX/VsqTnh+ZTyugaLaFtuU3XVErhIX9FgrdIq+TMY
h70AedrIkftHEFxhmbBJ3kaHmM+4UiCccI8RkCfFNt/q+TD66B9aWlemUV2yCdTL
kM2oaSCfxd2OxCyBJWbapLSpvUypuK9errWlHCzJm6nA8QSNqb8d0H7w56oaDH1v
Rr9FzIEuF3mMH7VL7vTNk/fx7Qoal7eMxoFpebZ5AooCJoKcCyubmN+MEsoNlXC5
jItJHY4Qkbhgdze0gYMfwjmIF82+P71IsRJvC33eh9mYuV9oQPCuXErKWoFP0PlD
pcUoPOIh18nyw8aIxEmGXQvVZoLGvF0dtYMUxC1OacECfdp6Sk3Enjky+5OcSLkj
1lxRUTlCxuyZy44qaSc54zkD4xrdTR8KbG0qAOqBx4/5hzDcGA83IZOQNn3IzQ4b
xbffrlY0FUTvGfaAZgLfAkQf1/UqES3s4N7SQSEe/g3HXUbqgj4WL0e2okxfdVXY
B2yhHHZrUQPi6p3bUFO6ogpqrpxvFrizlYCZ60ng+BFi7NLoBQ8PPhYsMtRwHQxI
Ry2ZShRxWTfyDE6/O7xRAs95G8sJtVrE8yCKug6W/VA3JWMzRcEScCPEcOoF4rGf
Mc3tkGhf3VGwxqW1mOz/U6YEys+DSrS6NWiBe7j+7Rl4XA9nZiGmI8JTiStecft0
kwmI/FeqPVrSgoSuPtISM+3I0ti9YtVpW7THe0TTfzmeaHUsTBnadJWYX6I7UDj7
I8n4YFeeHdB4GKq1N43m8xZRz7ToAF3g56OFFc3xessFXQL9S+X3tPe6Y95JzJX1
QM5LhSfZDAyf7iRkrPN0LDwEg2dNN3pW3idWyLUjvgv0XHDIGuOD3LQbtwkqI5ar
hS5LYIVQxS8nYQ16wZsa9EOdcjno8V3tStLa8G2JRzXaf0dANW3Mltg/Jg747ogf
kSzj+uJVWsCpREjEGwHqJYWTHCqicwBQuoRmLbYHIAlyIpijshDaUG7Ld0lRAztp
pNiYyqHmA5op8VJstsriCuObkamH/Hc4hXujp10aBFcCFl+5HA83+nn5BcMVo1JS
WnkPX3KJzthz8py4EmBWVb/EhWTKoU8rkfjGQasLpTxbqrHmE9CC38Yl//9Dl2/H
u0PdqpOHIOj2WcSPdXoJzxr9WwoyxYg/Gbp4lpX7t7p4AaF15BjmE8XJ3GFVlrcL
5NVnvb27vMViMtM+tTVtGLQUoHdJKGGlO9eOXzlLAygSPArVp188ocY54QpqWmkb
g2BDi0pVzbjMoHd7xJqm6YQvD1wIIksUIinCuwn215d4DxMqJ8blGYBth67ChoIm
VlCFojbUvTlkhnrg+a+3VbT9pTducX/ccMeqRDaa1ACfEZJxdo5BwHNmEBuBSlo8
jGJ4wiWzi7BsScVCymesWrs73QuxOY7h6vkW1/Y7SZ6+7j5uQYsawmdxJ1gSv0G1
/b6goVZizVpzztswPuUjiSkWLXgw2SAL/ziZUOtXrOI70UiecGEdPrRNJaj7Bm4s
5NXWr2oRy1xdqKf15W72i4DZsjMY1tVLZdi3Tfq0FD2klm/KCkkynnPO7URr4sjZ
1W44mZdBrLR2zaLVKqBSeDStszjYXlZmV6aQdFCFfEflefdIhrTbbqBHI/J9RiPU
b7g31tTDNLPktVMJmPv06uSHt7qCBsmkbJoXZLNW9KxTK7QOShjC+cdt8t5n0WxF
ProGEMu6NylYDcobyrvVI4j1uho3PlbKdtypoXn4RODIR1KeYTr2yDBKiMl1r//s
+11Z8NYzBqncDQTX79LRT41cPH0ud9cdndlz978UMvkcZrj/D8EIk19j1sC8YDna
DQV2PbqF7fmU8eTaQR8UPm4nZd13/S+P7Xb1YVz5yKU9A6FX2ZcXHk4dLRxlUNqU
zcn+Go90hehx9hie0Z8PASQhxVjIKhMVsCjfu3wyvyJ1x30V0lf0QdcHyo48j5/l
SZOkS9OmNGMkqX3xtt6je+QQ2y4OH/kozEGGSwOH6VQ5sq+dwinLVIjVWvlZveg2
E39+FktX3aTY1d0vW02YxW4re68DFfQu1dL9+ylVJqu7d8ySdZiBGCdlXmFnsnaR
npbwMf71Mm1uxSOs938jbsorlyaNG73cM37FXyrMMHn3H4OyHHJSgLuDafDfE43f
3MhEaohF97o1I0YeqChP1/tkdrZebAAB6IGkv2CEeYAsbontr0qO4oVvuh8AjZEb
ZIGfn3nixEqb6YFPIbnhMBCotpb28NGR5gJIoo/R2hdpwbDygQTnTDPNuuQHBmSF
5FVk2TddZaty7g81ENLQQG5cNbFtCXx4z0rCFIrTyTGVIk0GQMU+sJv4W7PvVZJd
4LFdi+21JOcsJHKx52nNCDB5nv4ccCj+91dP1g97YCwsGXRvktKNSLnBnvt1vuTh
SYiUviH4BQ/kZ+jLcd1rtqecRgOvTnqTSkfMZpKeykBrAAYwDVF4euFGerWpJRqY
7zPIk9dWKhl28YvFMHBmMJadMcYIqIisznnNRllr3vKC8ETuauUiHtuf+epoIyu5
oGpUgsBzaBL1B1BgdVcnilTilo+GbQfI8Kvd+wgDOnlfh5mLEslNkGBYwFoaGWZv
Pg/tKdB5q3h272llj50DOk66UHhfJHb/gpkE3vvqHD+Zz99HE7P3AATnuR4n7a8E
csJKl5TcO1g3BVsW6wS1RCpEpICxseng7obHCjRs4OeJn31kuSjLJzCBjvCdeO4y
/g5aKB1EUlp8UIAU1fmuFTtnL4yQbX3LItwP0MgLQE6OeUXGq+r6C3T9vdfEVkmY
op84iJbrBEH2O7t2uiHNu2INhkqLKlrX1UFJnORjOWBl3yUG6o3cEArU9g4+eoGT
gd64A02x0756/PgLPMEGEvgIDBycplUwmoToxCRQdlPcXGsmqmlSem0PafDvAmyo
4cHbtgXGqw84TRDgEVYGs/1mnfHtCz7rNGkmJ5mil3DgJH4L85x6pzYDD2vmD0Zq
EOVETbk4D3z7InhQJKnD+lYBvFiNLGb0dH94+ZwxA4Is9pWsAVmLzAYXoLzQMDbt
0C65KlvQdrLynEAICQOZFbywMKjMbRI/vzqTI5qhqKG2OHt6iFlkuNfT7OHUC71n
p7p2RD33OJYG4Lb4EpS1GAYLn8BFyeeesk/LuX0TV+o+QQb7AZ6w3FCd6FOWuFbG
frfTl1zz6n8gc6snQOZ7CisIYARUml5IhDHlCdxQnDmQjaYw7Bv5EqxpA4w7pLSF
4l9awg1fPhszqHoMJOcm0dVE38exEQ2zd8F2aqNoemIcvzRP/ocT68JgkVgOAaCI
WSPLyqztJDjkil5Z8lvmw5GW4+cRnY4kduqkJqw5hLertGJ88PjimQEnJGiaVW2a
el6wNvX7ciErperRaYf7z7livTwAnPARb0AvCjwSa3wPvPW42v/7nom/ZIZRteo0
5rpSIH8de+CwjJEnXf1dPO3dmErD00vRuitRV/NMIvJBh/TWyUtL/vHiwUPGHFCF
3n8TqhM5uetkld4ZTqAzPgVLxqircCUcjEfe+XtTf/GWcXAtCFzXa7wNkjhhYdT0
cr2DSnTINJW4DTDDICUSQ8S1qQNnGfjlo9XuHMK9ydY62OtuvIYgMI7Ffol2j6tl
qaF53S+mm+WFktYSh92E/tAHntNtjyp70CWgmjR7wr2uSosnGUadGwNhEoCTu/Vq
cwSLqjfhG3LMexfmYeIMr2WbUnCjw73IBAQzbpvIe7ZC5Gc2D9+RymjunFLmArjZ
tVeORw5I0Ht8w/wEB5LFtBlo2Q43s373G/Y6H8Z90PJLVqfJ+Rop3QwM2s9ufZCR
zxYzOB5hOPjQH1HeAa8nGSqJ+zSfVXUx3G8OM5mpxEGaOVxbkXYBO6B5F5ZGq6XG
/ldQhuVYwwm1GDtGMI11C6O7mMR9voWqbr4AkMR4cAlp/CTGndnb9c2Ah/abYUsD
nM9a1RuwuccEbqjDZx7+NF7Cr0GLV14/iuUtrRg7RdeQfSa67FH8IvQepPiHqZn+
jiavL4NJt1wHO3RxOH0UbLCVje52t5VT6XEwzK0kBoDmg8KrWCyzwliJQ8dt6J9r
gOS9CsEVSkeoMDLCtfNAF/mKd8eBzIvqgvUTBIkno2bxALTjNIGA+81rG0Ybqu+j
j9PzupxClNPKW5Lkan5z1Gk97Ey9VMXeuy9jTgbkEsyq1JQLUfxbYKqWgz10pyFs
uFMCKpxaFMncQG6c7uMdzoJuzRw7k8VX1Z4OJNiSzZNwn7cquwjAd9ZazYryRlwQ
EhH776CcpOJEE9KSBawUq9oZ3hUgGKRN2EcDcFJvKpV/kV89Ua4p3NINW+KZbmi7
+Bwo/IaOm8g5ooNEe49HSS+ZY5AIpyKTURbalGlV50muE/wYFnztg8fzlcdpQ1Gi
fuhqCWVrzPWn/MsMbuLVXYyt7r2zjefwIDjLJi4LtTEcX6XB+Oc9JlpcxJai2QTA
XN116m3thabEGyv6IGURi8Ov9QeGR7mHn0sfl59rEF8ISAUzetq26KxMYP1G/qWk
7IkMGP00KVYQn+IPIuZNVSR8/OBbpjUlajaK/Rw0olqQTEUclJ1MAGOJVrbSWmCu
/8v609V4T5ZWvw3ZnXCca57E+9jsRFsHXMaIjSBpDfT1XoiYjcLiCc9VpFq2uJH2
wGaIZb/UsQ+8nN5M7owkxqow5yjssYVarvV3SzXGhhe11WV9ab995ip+GAPEFhz8
1kkE9augz2edW/M1L8uL5RiUjBbl++d7f1Ublumi5iBzTMJcua8aK221OBtq374Z
zoj3DhNGqOtwYrCLb3mDpalXf9wYYp7mwPajWl8fCFX3mxL6yt3o1s54xRnUCc9q
43OHmxRARuqIx1c5+T6uG86/QT6xCh8+qR6+awLfmQArBxndTnKGoT2i1tdrPUnN
DPfd6dS8H5Rh/tmUh9B9xxE8sBu+Jvhsx6CoPFFoX3Ejdg7dhpc/p7XuoWiMMnfT
Uah5CzllpYJr/FwLlFyXB7MS5MpaHA8wpm0KpO1UVD4wni/0xdJ1iPWBADDMw2mZ
xVJFYGW7m9ksJledi7eS5q/Ore7pbo+JNmndTB7JgHJ3sY+g3i5ZCtBYMqTX8NdV
10dyBru4Yq/Gl5ZweaNoVC/PryAWLX+qavOrZabE48mUiUhF5DwOKGDWNcNmHaPC
mej4Xbu46OQ0Aswhk6Vm3sUlCD8houE8lyjNcsOb2GUcRpeiJ0T7Vzt0Qm4fP2iH
fh7UEg4icXFEeLjzHzeWtRCqWXB8puZRwMdynUU4XMIvcTd4PtZFacUj/WraVSSs
CyX8IAlML4Sr8Y1ppjSO4b2aGrqCRiHTPCzg2k/pZbj3Q4+OjsBMAN9yTHPut8Bb
eGpaVM9NH1x3Au7BIMDQKUTEd25IDgeRTqrbx3QYqijTNzUwcHmBfyI4Fdm8BfT1
bV8ng/lJ9XLE+5dpaBzoTY/pKfzMFFQYX13cyoSfbLLVWHI/Ym3yzqLpO6OLHje6
ensZ5WyBouFgV1ZmyuXFz9GpuL2xXDILjgCfCvO5XQNFoVFHlalgWYZpnL1khxfa
UeNBNTJ2IP6uaXhINXWUKiYc+gZSn8Pu3/Drh9KFeglpFkh9dIblv4cAISHql9Yu
Tv6xvBgZR0JARsa9FsdlCE+t1fqtZlX4ECEYG0bRYWE0RDrqoDK/HTJriI1uVNGj
RjVjazd8MRAn4v1JJTdhO8Bp6Aw1gvmfMPWBl2txUdu7o0o6j5C3xmHlv+xzWmO4
Pg40KTT7JUU6hrWf8ZVrjLVlD0KwqfQ2rRhnZPDWAN38WYUOWhQ09zivMdEEs6Ki
A+X0Qc0o4XLaEJE6iSKdHsjUWuGzwmxdpTrF7a6ShIzMGuhfn4G+KvQoslEWq1fI
t8AfG+coo3lRtdTeGBDyUh9I9f8Fo4oDcG0/ZocMFu9Ldoibtz2AV/klVfYF6Dhr
AmzNdP0JRBMW8ZlxNe6aW0oPGvZc+2C2WmLyCUyarrmJyuMV8+Uwg7fMm6zQcaee
j8paRwHJIBsuc2NDCXK4xAWmy41R4G+eKJvb/A5dFaTstcxp6tC1wu8nJupLxxGs
65CmLchqliRJ4cahNl/zupt09tcAuYWoD63VYC+0fYhyo2+emmCDliLoqudbnUfY
HHqjLLnjmEOO6tAQ3E7TWCFqqT2xJD/FdDamkfZYYsJV606+YrtA6pouDkQq/oG0
0+GaNF3BQuCbn6lSKepvIloS/eg2ZEG31wjh0Fx+1ASWrFnTHBZIXCgzkmQxOHpM
R3mPmGCvNBK4sGt/5dYlIWy7A3FA46oWKBx2Dr0XufGO1GNJpoHw1MVobbc3dKtC
JwQ322mv7inZlrAcp4hIfiplDNOhscnMv8IeEtxYZI6YItUtyqVQWA0pTTUuLTSo
Y1/DP1NVi0EFyAS8qwrEk3sz05HcDxLmmeT56wmi3LcXvwhxZEz2P8UhQPDL7y5X
GSZn7uiWrME55gP3dfZQaDZR+Ttpm7rV2HAhwTSnDssKmbyMjSCCyF2PU4TY0x7t
Ahpv9WWtZ/4QcOFMotrKxOUV4SZlB61I6sx+rM8QfrvMfYmaK6nGVpt+X9jRhC9+
acXz6FljfU8gCW5syCYwLDYFBDPDUUzu7v5BSMZByrqF9jCd0U6/X7SZRzqUBWoC
EjG5DIqAA+QL3IjB9cpWC0tBQlmJ/BVFxCaBqvQQpN6esjpiVDQoJjXNYPICDBub
vkuGF/2jK+h5FOwGYMkrUnOWaT0o7rIREauSbaBufkHQp9SfQwwTNTCXTbN85ViJ
kNczLl5uEa3q9fGi5W1Lk0JeiUc650q64OBYcWq//mrabwCyHELv0aJPBSHUqXXq
a4KQpiYzWWYT2S/ZDdX8UKeSgym9vS9k/r1zRj+KV7yMrqU3OGXOXJY61SG0meoU
DJLL0hSsx0dArAJncEQ7/bLQ+xUSwRmZsa+hxyoMPzDU6L5PV05GrDTH05egm1PB
WSADJ5f4hE7QJm6e10GJJZaZ8QLBpjpznbAdsaWCWKik1XvKJMflq3kSvJxFhI4W
h9qzPHBBRcZfvqA8qq2aIeDbOYbxFq2ZqsJ7Lz0O2EStyGNecKVXCL5iYclLxrrY
E0xb6LZ761n+hZTIHIrVOx8f6qiqMeGw29sJjfiebMh7uS7GDcK9UliMhrtwb00i
/YjUSBRMvJ4Mh7Cj71Q/H1/nyYrMfqcjpZKV/4x3DoozpQYs55s6cPomD0Vfa2gG
zLB+HxR/ssR11rFO7ydCZUCchmKQv5MdNfZd4oFLaHbhqHyksKNg83+j+7JUpM+d
nAYdzhgBWrfp2dUyfEx9f6ZYldvEj/zRX3okq97O9FxCVh4Wk43EnFzulZUKg8+g
/VxoF88YA0KTQ4LlvjGon1/9OeL7/F5cFUUkKOIDNtH6G1kmjBNPR5htRGaJYiG2
hbLq1S3rRkX1X90JnAZ5X6Zax9lv+2L7kTFSHOzfHcIzMsAnxByCWQwg2MzJDRTv
VvrrA/v12WWsBA+FLLU4C6wE704BI9A8lQD4CuCTdQzppcRXsgVKmV6wZKCE2Evm
F72Bi5F6rWNN6C12yHCc8nXm8KIuNNxwQlraVk/cLzf9sJf0DsrKPiCwPvqGKFuj
DNjMURlhLnRxpdTYg74dMwkNeaH9e/7U474sai9BcGFbmI7CizNdPM+eK/p/t/yW
Xa+zWaKjbpywN5waMbuoabA2ZgUCIq/Zi24LmQZ7il4vK+2kB2OVHX0V/UC6eElx
h4YeU1cns66+GAQ2cHn3qBTvl0F6HhHDd4RDGUudzZDzlL+Dem4IG6XEMgplQaET
lEufGYtooRGetfT4yIjwgqkn5YqzTErM0BgwAs4RVkAlyjdkHHwh5MrJnqx+0LPz
WpMBlNGpr5rtnNWvJlWaq2Nh/mG8cHlj4epLaBFkpLcLB1G29vlW9iNg2zPgttg3
u0OdCCGz+pwu0oT+dK8nfPjSZjKbpFYioVRH42hS98Uvl+H9EiuKT/ZivomvFwZu
GEitzu286HRlC+DPHN+mar6+bkEXZ2XzIjlfL20RsOA9fh/oUbOVhlpOtobhaLDs
aFp1PFUw/hHfwUmdYmaeqi8Yx3CQBXW9/k3PXOH2hXuwy0BGsFADxTj3iim9UXDj
kjxX/4XcPMCXivzPIQUP4+1AB4TSlsFCKuJ89NH4Cty7K8uOlaTVeDnetsIf9oPh
f+1/P2xODmpagER73IApa7owoLhBdXiiF0yXDqR8tuy+CSxhlI+WKzA9t9dyGS2F
VUh0MqYOXPbyc7jLW62KHhOpZKa/tHTsNCoyeTDUpYxXyXuaF6EpG8kFCAEMiPH1
B4FCCEVPbQdgbfFri485hLEFmfIb2Y8N8vdte40d7w7dIAzfHKSnLuW1RInZ3sg9
w7BnxpqpVcxjY7FgCY9k1BcPkP8gZXGZ94GU88JaaurSB3TbLvSXrwCxwAqK9mVJ
AST5NHjQxkID90oL00GsUkLtlaeIhJuwX+2yVQvXn1lGvP5UgcUpGgEp4uZHD8PM
mJGWUWIC0FLwQkrU/IV30blBinuko7YT+qFVDeMRTBlfRCzzxaa5VJA3C94UHans
I/P4mw++InkmgLJlkMsKSchcQjsCZRVU+2OHvuY7y1C4Mpk7Xj9rX4PLk9gBD8P9
RY1MgodverZvlX90ESoc9p9BqCi/Cpj/wUy34dgMCXjZ3j1KjcCe+4I6o1yNdrYT
s0JDxawIXoeRHRYrnMgqvCks117MzQrrZ+5lbu1NF/cMuTi1icqPA5v+xnBXk9es
HGHG2K8kpTJXrGXj8JK5LUO70GghUV45u1iZXS8AiXrcL42cUAGIHHDK7GPPzOM2
9oCbE+56se633Ka4RU4wXxQ0oxGRUq085s9e9jHZsk+WfVZOFgqS1r7Ldv401zfS
kqD6bmZua+J4UdpGTYhVBmKg60RscmTTC51a1Q7d9L69ye87PjkcpYYIbnYXovfR
Rz5rZl0iBaSL6X0oek+bntO/K16hbXKIRkliDwyomNPv8l/h5wDmAucfakhIbSCK
31QzaPcQ4euoqLu77K83G3t2vr6US12C+TQZ0rLnUfaV1t8+P6VH5tsyBsgG/dv0
GPGrHkgxvWMnQl2/a3w3fxwV05xwvaKCGhbEmQHAulmoHHtU+OlAg8cBpA4OsOfN
0tbp9EfSLin6vJVbKQb86UUGRdmoNa0pkNVDaSHt2Bf10KaBvDdZuupzTt1IGnYI
e5kfVAdCqdcIz4/VENwIV+VLBNC2n3ndZ8sCxfwHf60xV1dYnXQyMPEyw+GTCPTJ
ymHO1Lij4/qQrMjkFkae9uXrGwRSpERK/yXCSq0o6IQx/kelrx8Vx96D+5uavO3w
RUes0YvhjTKIkYRLgEwi0iofLRION7+n3kzTkWfsx3LkWyxptbUTo8fQqXaFMrn+
fhq73a6GqPGEEeomKTrmhAvKBCXfbkx0D17ZWLug5QWAP737xmmAK1tloitPlcbA
+uUTc/XlBRgNPnVZqSobJmlbdu3nsqCmgxC3hobH0hm7J47zIDLSEdM1EX38UOgS
+0N5jDi3yzGP6PmtCeRleQTGtR97VR9joE+sfZVkger2gcCuzSEVGxzj+8la7jlD
K6+tbNC1jzNRQTjwn2PuKXQsIapgYEJzNkCjXstf4i8sfhT2W3BpbFYjdDHA64+v
hpULIW1GQ1d8xpDuKDuAqpg+2R2rjwUrGdw992dwZ4MAULzcDuYivhE8Wq4UiaLb
K4Hnr9GzXUmG9wZvQJvlk9p+9AtnOSKwfAqigp1pRFozCu6zfupeWQLDcd0NmuEb
9SHE0fAh3ZJZHFbMrVvrrSoi/uHzsErL6yZjG28kFLhQWbRdT/IOMqVCkSdAuwtu
iNkgtVad3GiHGYb2SARw2S73g9kvwZdQW5DlFOyc6WxyMVPekIEcXJlTtC63Uj/m
CaJLV8iBMJyl8vS31VyRxiy1LmrlUGzNfMoyfgQCRNmSwdBqSdmmm1i3BB1ixzEJ
r+fAZYh5WPk27SCGEDFF1riAYjG+iE5GLIqOcXKU0D8lus2CDCyyKYt+OGHHwe+/
RyzdIfPJy3phFk0Oc44PPBxEY9ETs5Oik7mr839cKk75knkD9CXn+8X9W53tajrC
m1GCJ+vPFGqqMldEWpGIjADsBJlsjGLv7CG/FAsqN7AQjusGG+zzpVF/8QEde26R
dVigNXInlBI8x0DKyVRbL7uvO1ndlPIqYySdlftWSJ0a1SwHdsAL99qnDQO4xoVt
oz9MDC1gkzrxRvwbYZES9rJpOIkctT4C2210+I6d84f0VojMQLepqi6/miO/X9J4
Q9DLR2GF/i7vhMrrl4/tnicoDWRnPWbFvVYQbuIxBM2F9EAzzb9m0PQrSYPdgpwo
8GUX4/Aj9U5Tqqe+xbZLQhqMXcFTOxXLJuLYJToEvZ+lUyDphanYOZYufDrRxMjv
5bDBoTtjLQl5wmoJ0WSw/DfEA+j2q7WoFEvGAn2Xi6PCaHBXNrhYvDa/cYKMnFLC
SnuosLfQwwE+SaChILWJ1EGvhqP9aGx0ng1/8FSMuiPZYSjNzIsBjGL/uIpCPU2a
LKBap+A+b8YrGK2w08UvV/v73J3tmHdgQWbDeUapZqAwvQo0fO3q1PTNU3nypjrB
8wvelwlfMcDEYeyY74SsKxiMsqdxqs8tz1VBofiVXRxJUUnpVdCMZeEaRYJtwkOa
6DrkkIMmDfrd2TNeW/8Iwe4Qy65fh2k0CLAWpJC4ski6w6yCIyIWFQZzR6GzxhzM
X/rxPO9EkIPz9f/mDHB3Md83iz97TZURzFKX25V78wveF/aZalsC2Rs46TwlNQFt
EkTXVuCJhVYfpFuo/eqGgVNA4NF+UZqJqbAPcLHwXr16CRFb4sAVLi2pmLONOFUN
3l2X8Gi4VnuzeqQf7t2lYH3KiPZGjgqD3mHAIAse9dZX+O6CgRIhULxWBLWAdwPE
mva1pWGEF5XguApXSndFIMI+b2h2cq9IkMp7uERxq74K+3LHjjuHziZ4J5HHo3iC
0XgJJ5BjCvGJxcIAhdG3VeG189yczLGQNa4TLIOtmhtHXQu211Aby8ELwRiNd/lT
uf3/UonKJJM0RQIWfwcFB+TXbKLbUzVGV5uGcGtTtxetFVp87JONINwvPSJV1mxJ
YCa2rAepak6NtPZ3yl0ESWBUKBwDtaTXQA+DRiYl0uID4qVZjpuP1aloOLgXzBZE
LXb/ycss7YZCU/Ma8lAfZnWCFmUACjWLsYGZi8Slt582ko4Jk7YaIvV7vZF7ROz5
FCv1eEJhSL+qeqIJK6aRiP/Si493E4rsbiYCyBlm0PyZjn0/+9t0E2Lx23tiMQtg
AmnnBmPoYXs60YX1rFMt4Q==
`protect END_PROTECTED
