`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
LzJAxTc7ckdCft4sNAmjXQ9lkmBgaNf+rQITOkPPqQrWmUqTc5aTcmD/EL4Vsody
wEYVhSxvKakh+935jtg1H/LsQ07y2N7q2LN2cvnt/aLlWbhG9EY6UmiBqGVzMHfb
7IbUIRqbHAjXZGIOrjEsME5KbCf/ImzMguclFI8IUV0iNqxBdTnjwbOXvu91Tn37
KRjzHtcFBRCfMaFJynr4EqUr/YAv2bwRcVX2D54cYAtcGpl4+lgpBjl3fRtOQMwx
OCf9c5uhjVar61VM+USixcX3oOGUMK2FAriG4lfCMLM=
`protect END_PROTECTED
