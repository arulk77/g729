`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAcFvnuTR6RpcpC22JG0760zHuwRRlEW1WBEIsfOSEcq7
aCAE3J9pJ+tJ+gk71VQAZ9GugNlwDrMRJh9FtmIXW5nKTMD4ymERm0ayu30Wkg70
k7aridQAZXsLbvuWH7UmPLs5VTsg4HuynE/293X4iY8n6MENXHO1AZBmksAIA0Ml
m7BFEtNO4F6tXQGsMyawpPuBMLcX+5eHlvbBleuTm3hUtV312GMYWxN03HUg0K/4
gy1HnJaicemmA2se8Nbli+SnjdaxnCL+mYd+TZ3VDW9NS7JEhINwtlUSgrim7SBu
Rvc/2AfOoPLso3fPM6nVNoKUSwQA3ieFeD0PM+CFmSGb0xel6RcGyKSHsfIe/zXS
FMskbwG1h73R0NiPMx63BhekwPACKk/Gw+c5OStFn0WZluzeXMIc6wN+IABRGy7k
tfs6dHJAyzbKytnehkuRW4xgO0CkXvl80vQZ5ZmLkde3UPXNktk/us5Y0FKCnMUO
FHFePIJ5WnRDWKjdTGvoq7TS3ZDgatY/ZlnzeRd7g111ncZXb5dc55rsQuhV+Iul
J4o9gT0MT6WVb0rMzjhjYmg/2OTpvTnlXYIZJXIT8n0pwoHNYyuEi6O3S/RbdBYK
7UaP9ldZsmlD2znPwBaXIY8m05uJ55K5mOEoTJILZEIb8RsJycZLWQ87zv5TfKKX
GtTyw3NWBph2SpHDn12kVIHDigp9OFG2dNswGwjkq/9GmTlDmTDedK1+BOqnd+Rj
URFktxdg9a8WJd09asc5YdZWWQb5H4kDeVJ8QSQqNeh+D5Wz8LX3PLQBmg+fk1/h
XQuV5Xi4Zhr82LgxhsujSgtCtnBKstCxDkoLqSCLd0JfLeLs+alO/FWgHPL3p22H
M7KqvMbL/BrsyinX0Ef/r55aMPsI6PJ42hiZLt5FR1dU8p0e6Uf4v5uEITaSaDzT
PCLQy9VyPrHvGGUWr/egm77BzIftbXRqPHXNf3d6HBEagxqptdvAjgg98j0NFlT0
w6fTSm1uZU2IvyMoM1EOldyKaddG9ykkNuHj1KF56/8cTn9tCxb3VMgp5apNwdac
K3j7roLRYFjcO6VwDf5jTxjdGsPp8fQn9C+yfQo6MDKiavGzNRKvnor7ZsbAhomE
9o/uXQMknGYWp47rkaMJ9nGY6Kas/+5pZylvTCRrZUmNBS9T2F/xI8Kl3USaOC5C
/0VfjTtQwUKn5/qFKM5smZell7DUR+nmnvvUT4g5n9HDuKGxm5hhOrhK+GXm/jv2
6JcfkLrbmJbhbAJ2w4wImSSX9UzUaHS9vMb8/z9+E4vbmLv0n+uAPMCCGXpXK2rw
qjYD0DoGH8kq9vVl0pJHXxkpc9r5f/Ld2wJ0e52kRMS5C6fMpxvOwAYl/KHbdeVE
OfrrScFsogC0AYDZOQr4oxNPQUr5fRRrbNZsWrVrMW940GFwabr00fxLbqtjsd/2
0xubbklIlvzleFn1B1JJC1EjWWW3WIcdwG9zgE7+O9QWozyFxK+uObUDo8wfLqEG
B/cdtqP3iTTIr8mGeZO/z6BbfVMHB2+FL3bRAAYvgu4XDpK5Tiy5T6xomEcL6MVd
ulAA9NSB7LNS4xXXTGMDJqtjODAlFRvg2+GExRfQRKv0OV2f+A5RtBxhD9Bq7L6u
3vf1yK+Y7XscQ+BCuIsHLZjcSVeFPhHZrBL2ynJxzHgF6uwSMeeacL+psj58TK/K
uLH5MEIXZ2Q+QL3y2WRPQ15CVk28E2vahcz8Uy6xDI/t2AqDNXcTUM7sJr0+0Z1y
rw2sOdO+W+MAML8l7kWTN5W0lbMfvxfBXCSy91w4heGaQ5rX0IP4PadWxuKHMp0Z
g4kQr/hCw8KsGzCATZF9DUetmVxLhmAeaqN5hm+khVK05K5x2g21qW6UFA/2r5Br
3T2FrbFsnR9Z5WPk0VgZn4IG0VEnRIdfLUNAMDXqBiM45bQPJ7cQV3fvpt6US64V
4GoiMdYBePz7hJSzFw7gAtq9p7j8YVuvkMvJ3A8p/IcTMWm6Bpoe9719ns2iLNJ9
RqReLIH7BD7mJtWx4/ilozo2012CtvJ14xIQ8xC6HoCIbBKtgvZQ4nT8REZv3gFF
IaQOjFI6pwQKAEM6ivbdfthGEX53Pu6cODI7ckhVAdRiOoaO6Z6S4Xo972Q6gqaR
hKhS9/hv+Y349AEaBeY2d7F/6acNe2J3Izaq6Lsw8+xu34Ml2vW7NEttxiJa2lBf
bjSvMbD0ouwLhn0j7efKJ61FlHq7ykUhJ+XcYlZKfAQZeoFDNaZZubE1Xl3otEa/
ClaUyMRnTGjljDFahgmKGAjD4d+XMUzz39agTvAxvDBN9LL/gZFhTKzlmWHrqVA8
8IpPNSvVebU2XLLScOwQozKpd8aINBb9A9vYlrFVFaZpLWMZd1tymR5XkJ+W5Cqa
wazZj/Um8olttI47SSu8z8+MjFMDXLzzEiG8ZSIDvBAmChOMuPqBoWtZWT4bNmxE
GZYfp4RhM3rKu30yqWkkiPORlU53cveMc7yjVArGTErTBeitaNPOBREB4qDqj2jI
Rf9hmbZ1UYiDjAvx5bcmNw3K48/CJluI7ivDuS70OwWRPIv8sxN2nQ1BGTrqSJf0
sczp2O+TzjlIRfKk5kgB0OQ82H3b853qOn0zEt7DdgJWTR84xDBQaxSXQ/3b98TU
1tWhDsGY3O0VL6LYnf8zPgFbv6JOp6q4Y4vPHi8E3jInhiYcaG8Qudx3xeGx4RP5
m2kdetIlav5Q+ILzsuTOMUWwqbaJtFT52D9X54q6n8HrHrl2Lqb2BYC+l8DxXoZQ
g4t4fnljzsurFjQNh8gcCb/stYdPNd3YC1esEYj5rsfuNB3Gg8+/WNq2fawcniSG
i//vZEwRqzHFsM6dtcm9Q4PwzRAalKbby++ZBO0npDBs5sD9jsKNvSvEfKKM6LM1
wd3Mnvq86gPYNtYtvlCtw3cBc3b3PYJV94PJZIQMl7on/KbZqwnRfpGrLiDWPYTe
D1+ClJUGTc9UrpVvzYv8ufSYO5PH2kIe9otHeTf3XVJffspO8N+z3wago0rUPhKA
i6hxAU7WLtY5tCHjye0u9EAUFwwbRmJGd8g5rHPuZg8nyc7acc7AIhV1hypQDfJT
fBm1wfWPnHPK444q+MSSy42ieqmJPsoMlMjDJacS06Gpv8OyTWdEmMAuiMjQSX5n
8YAizYJRx3tr6Z5M+PUd5mjTp7u89Roz1aYKk0xGlDHxfT0Z80Su6O6pWwZqVmPu
htQ6UKBb8K83tjq4kV4QoPtcKpzCTW4qygks1q42J26nd/wEnVRoTyHopOpCUS2J
1WB+krz4yL9ekqPJMpzzOTY9HJZJNeclaTcVpeWRnSbNNYxmwxrxjPC5P0pJHw3m
iXR6GDUSqaJLHac37Dz/gYUvc1+7F85bvhKNuTTIgWvBobEiG0lEQFa52GWH3Geu
TNoeKnri0O51koHTmGz65yTSEJQOjovOUsG3Iw57s2nyk6jjdbFz4tLlZrVNJ19G
f4XGDT7TM0/J5XqunRaaEgYVZKxjE8O+s+Sw7jsgzTmEE/vkvsQcrLHaGxgVi25C
sMmHn8sjC7/6ex9JcEsuOvL7k68wLnRB1iWdlE8u3BRV5bGaeS+BkFre9w9NxngF
4znr+MDBNGMZ8riPmrYOaxLwR1mEZsFtdI9lRhJrvg9OvuNbFAMVrpdx80CpCvHt
RmI6Eb2patwyuSjB2ijff5+8pnkEM0PW6TGV9jFDF0y99Hdwyk0V27fnZQRAVuAt
SU4nJ8AE57GLnoAHGaH63OUoMES00oJ9vDchErsv+eGvYM69yspZRqD2Ol2CuZ4l
tN713HWctJvqcIvY1zgAN9+n+bKymx7r3hC9MlEfOx0mFJ/xbTyVwWWjXk9lFXEs
NLsoWxmBvxNQ4kkc4pN9dBLGkW/NfnVvg9+nT1nZVPW3JNuP03fZAL/PPL3MzXIP
EF23xMQQGFqJMc9hW5y8ZLTn9Q2XxoLuosua5mOzNUB8aV4jW8R0NmQaEuZ3xEw8
2WqhLepi/3HJGbAUjAmxdvfhHDeGEPpbyKJ8JinM57aN8gmGbHjr2bGKJyLvXKl0
WPHSTSm6EBFTGmbrpY7otfizMDHFFcYgNuv8v3LLckTzmxgpgH1NdfEGrySFDkbZ
cDaknG+TThs6hnKjUw13LReERbX+yTw3FwQrZJvV+8Km/avyvTUeehorJeQvwuPi
JeLFc8+NUX9qc06xpURV/eilFSDVZkcLQpAWlv5lTq3WU3NV+alLyNdkkr9JbwiP
/ACHmnAODVDe+oej/g/SX+si2IixO67EzxSyjYoMwwRptn7Hz34XedHldoMPhB4P
uybTzXRiiUKGXAADUOIsBEeHoDWPrkmxTqhw76oGj7AytY+6BUzTTOJz6qwvmbmS
Sa4q6DHhbqUljWBB1Y3XtunnjJwuApDIHiGFEamBHRdUJoB4vG/rThTmDTrfTrUY
kLxKH7ZE36EMOYmzvgjpL6+7BdX8IpZ4xbknvwhf4Rf3jLj6lZcKrgHMqKJW6dFE
VogosRsVB7ZlsUfeDxHus5OLFrg2QE51fM4d93ZLudfKlcC5dGjXT9CwU7EWRdA7
fu+FxLw/gL3LnlbVW9MhhNHKJFOY6k1rtGieL/bShKRkCD4OrhTExvgfQzV4Sz2/
EFv3cOwuBprKJDqVqE6+c34pNKIPlY/xOaH+VE7P+BipJN0JlHeZixC4XNTGfAjW
aaPBkQVkOB/b8AXG45N9kH9xbW8vYhKogA9i2OzS5dqV3AaiO2H8c2D5a5TDaO4x
+Kj4p9s71LZtcwFFcP05IyCfCBvLFPDho4HbBr1xnvkUXm4zDEdn5RjfDuhBnil/
Zk1llg70mEbj8RosFawnczOCcHUZN9A12Mn1aRVwb2e3KYcoYKSxTbRVQDA6TRqC
1sc600NN4j7f98TubRjCc9KkJ1XZyniBGHtP37KwBj3gXntYPdCmLa3QjGngPt/+
gqQuuWGmOVYMrIPwuqy2MjGBj3yUMKvjGekcMeHtAEUVPvvYXiX0CC+GuXd5qL1L
LARbGDZsjYdbLIKBkqhFuJ3Q976H3iNttn1QV+sB4mrLR/LiAjjb9lRaGOut6Qi4
QchEjIseO2r43NOFKidOXP15Z2eMhqgfYoTVhiV2rJoFWANpY0p4UKvTHUuavvtP
QfTnbsUrAxT5tL50UOPR2VZNioQKnLaWA9iUUxMm2c9+tx73bFzWSvZ2cv1+Cdhc
lpnO0C6jIt9r4Pb1mY08M56ot2S2NRaUXSORfPFtoAWB/ri1OP507bGOq/wDV0eY
8181IoLufjrwzRAGLe85d828coU2kgVPmm5Lobktk+PTYCYDSRhI3e/9Idz4TDrH
ldAugxiojqcqWFvgEPqn0532nL5Ns1HAtExBGeDtwT1IzV/RHykrCB38Bnj0rThS
YQ4qCGHVUmvRf0Di+k96Y0vaW8Av/YkyyYsWsDJFU0n2r9W+Vprlm3RnzKhIpeTO
tBB5WB+X+/cFYKYc4Vn0eKBoqn+Mf/kPm4PV4dQxy2TvBK+kK9n12RaWj+3k7wtL
8RlRXDfSdcoeLtWdcn+F+s//AxajnhRDzUluK3iWiEFnX3Yj7xFwJixMUzIBCZF7
NwV0Flya35k1todzwWd7pwm9WqzIBdZOHFEdqDeNZLuZMgL6T7SVPHDAP82rrV1v
mOjbbi0XXwMRGfz2nVkKacR0pwPxkTBXkffxBN+ktV1+h7CNcGVd9BvF2t7GrFD6
UWEliraVAwZd1nA+XpRQXf6Lv1hcxnti4nuIG2az6wok9sGj3b2ERyulHspmlapN
u896IXX9xef5yHavOpO2PkzV+d1vTd8J8VWaIpALl8IBzlwp/uzQs8lvokUaxewy
m9wy1L6jkWydcQBuTZXHGTqYtZczGqGbJTkm3Kz+DXEzHmxynjT27kaBczqyRV/d
8qJlRLb/Ag/PgByNiBp97AToIgRO53gZmF70uXb91WKODGUlx/jxoMRLQ4vOlIgC
DgXHTPWBuuT3f+9KuTsJ968K1TwxD9vWjn4D8LJnAHeRHkrp/r1VuAZjPl3H+JLr
JredA9dwny54osnlqoAmyo+0TIRiqdvXxSO9sB2M0Jir6skV/oOP7mV+Uy/4zK61
59Ky85EDCZaxkwp8+70rlm8N593wp091J3GFpYF6kBgctHrfOTm1mDh4Dq9hTpRM
8AnhrK0d7kPZX4jySRW6E0qaOwWqe3K5hUXc2bGFIHP2PFC0lHp0n/btNI7DVk3y
n3BbTw+IUSAMioKsueSzCjcRCrDUNc2dSlcfejeJ4cg6dFK50gbyoVcfk2W82kF0
6Wmr84BcvMJbAGkG8lFXOTXIpQRYNeWRL1vNW0CA9agifayh/JBxuEidykHZNeXm
ZT1W02nO0N91ai0kGJOQv5uePsvCFwaKa3C5N3NXgEpLCvmarNd9SASM5nRmCgGK
2lcaz4GpEDnQsDhSWvI5Z5ceRT7lfMZD9ljfbkkN/ciCRLTWuKmjK1cLlNkiUr33
Ob1qBjlu+lCohjsHvQ7mZxxNP+SUKq1HoxgyKoGw+cqmH+uN7jwmwbrsUt+DD/1c
nOrhmtKCuCckUrkdtfKbTBOFi7+LkNLP0EaavnjxPS17/o6SRo15cokaBOh9eLBd
RbTrJEBhcMNAUhw+T7619hqX2P4cpZ7pO4soG+DMyIcw5ezW7IIe2ux8gDQjpsc6
5Gfj5Uj34DIZ3fvQN055yoLy/3AAg3KqFW1Wiu315QkKCFrwYTkhdIPgO/YxxJOu
iJL8b4V9NdyyPj+0JPtZImIAfMrZYKY9JQAPWqAosctvyMJxyDO+06p2exJYzRBy
zk3gH9FvSJM3ysX4FaPkpS/03YkrV/tbBi0lD1QEFgStrt+qazwJ20hg6CK5XMQu
h8fqZvQvVvR5WQTHe89GYui2lRL8Zvb5dW+mQGHoi3dB5oRCEHGmfzS/ZVCFwN8Q
8zYtCP9eZZMsnq/ayoHV9QGx1oN48i0byEQamHeyZ/mRRupx4hx//UPZ40ebTShB
iYn03Xj5QlPW5+WYn85D2vWCGb4NttJ3h0nRGD0a1qidWwUr+BWdMKodslZ7Roi0
wlYZX26eMpoZqUJVWIrKW31XbAi5Smn0kgapZ5fWA4DK4VuAm2x6xfR+96fjt/82
LDGgsLHpOm8ZNH4k2v+YQbzhW7rzQiaFCSSNDCpLLxPQHKrpP2pnHWYh5nO1R3+x
gPdsoYVS0N2xO9FoZ8ZBnXh0MrRQG8aN4a+wkIvKoJ7E42OwwgIZac86fGh7Yq9o
zL7ZrAUpcHh0PE2xzwHuteik83IoAn6j7+5MGLQHM27GqapHnvVbGv5nEmmq5Xit
GhUsEeq+PcoAzq+AkDSwC2h+WX3rJMvgTSYwuoo2ZIMCfNN4MA8WAZyHax5AMOtC
tcUAMA9Nbfvl7drp3ymBUWZfHzo2POj6pcb8iCNw+N7g4NjJu2/k6YUwXZtkkl7w
SWsn7bKmwEV0c5rV3Ol6Ods2kIiqjyNWcYe9xPDGM41R7ctasPz1Bq8tGyOfDmVB
Xpo8hYj5jsUJCXMaR+ozrBTW3jIQNqtJQljLI+lBK2XH98fKyN+IKOcVmaP73NjV
LZVKTRS0nfohgrfQMOl0tbA37fRmOShu0wmEfu/pLiBmd+PsjsttfFXo9iiZVeTb
I8NhFnryt+sq0L+uAJ6v8IoolKjq4bS/DS93IZtgqRsqyJpwcdzt1rT5iwKggPgG
8Q+tCMsbc71o6SuDz8FAOaFrTy7MLivgFiHbdIckOdhImhgji/AQnj/sX6v5Z+cv
NifdW9C2NwvAGDzljoksMqa1PKRk9QPZk2LnB2AihqzTVs+Uxvh2OghxGnOp4wOu
ZAYu7OVWXQzd4dumO+8f7C2kQ3IkIODj/gLvWjsaZ/WAIAFz7gNTLN0CkXy6wyJ1
BXIz2uKQbg74pjPgyE6oAUca/z3j3RjpSuRt3OGchkkJ6qx7ZRdLFxZkl2MqePXj
/0X1p2DLKyMEEebC9LmTnxOb5DZOgW+EmNOlzabWYPlC09MEgWDH9loGdR4L2uhr
egzliNeP9X0F2NBI8O++b2Wh9PXrlpmrPsLhcY4KFaDHqBE9q/yENh7hcqm89yBu
L6ZJf2ASsrPn4y6EsoM5SIluqaGKzpv5LDOyrVWuju2khCpKvIppo5nnGZlodcLM
lDkyx4nMJU2czPhrAoeS28Xcb12F8STPviQO1wkuK5WmwFgWUz0A7LXQpKu3dHZH
/CGnZ9RYXuIdTFdDtkgo6i4YBi7nbluHirTp6+ZmaWB/RpKYMnu/JcBJDSD+0IYw
bPIvG/5MMedpJMJAva/HBNd+Yn0/9khLU9BTkD3xkEx8QuVe0YwkGGMgl6pIuFmC
2kbzSU5OZlas0EJgiUpe/vqLcV45AFnXUX0jIdHpK6N0wKwt2TN+UdjeiYXCH9i5
cCqLd8rDcQw7Jz4HoEjNqr5oTkBwmsTtOyt6q6GRobh/ze+8LMjJi0ElV4yQqCxk
LgAD/F5NT8xE6RvdaRVLlPgcOcj6JBVrv4/M0qDZ4TXZd9aFSXFcwWW6xAm2+k4T
r5Re93PcIth3T2GM8W8w9dcErVmHG9m2GP8h2XQmIYSoFtZSr8a1M8m9iKVZF2nC
NlLLwOq4fJ/V91+DWXRY8y6G7kYG3ZDnJHoipaByTDWxdoqveM/84mD4Ya4kw26Y
sYf2BlIEfPoxt+2glRucZItQ0Gdo39Mhm7asGGG3rLfCaXB1WHmm2F2lkdkqCuIc
DISIcibKSW+e2YHO3jUddAkSjCUa1jD/ehd/OechUL06rgd4f277gJTx0AfZhehD
UUU7EIxKJz4JK2leseJVLnYE8kIJxlrHIG2d8pqQ6ux7gVQeSFOid5nfncpUFkgt
j7hQcQC3MJ36PfKGCzLrLMTwDw+qGrODCoKRCCXj3/6jn0hY0+nANKk8fXOWr3f/
4y7eisQc9GzQANb+blAikHZ6JM3s4iHsNJhiW2cw5uaALslAwtpSENzEXSCpG73L
Cxtz9nFyoybPMgWEv75kEFRMYsNsHe1Glk6XoUgulkoKeytuJVPan+Tlg83pWIgL
D5WYVxWKVj2Hf3ZoYQyXD+/dSSI2O50GEZ5W4RpOq5wnbnERqcQN9HHLx7qWvHXw
Qu7pzf2S0pm2oyZtW1iBdR8TELLiGVzylEvufyd3qoaMSKtIIeN59VLGpuzMgzrn
iSK1xfU4GTmPm/SDl8iKprTVLHVSbbWyVqfi0cWXQaTZj6iqUtUJrKoRoPLTa4mG
KHjm/vga+qB4J0qr+M3+6304pmCnTR7HIJLesQKEp4N8MtxPbT7py1nuXh0cx35Y
gYKWrtMJi5+oGwyyLXP+KTk5GOGwhBhcSLoXNIfXerI7LA5YBnRnyMlnjeFkh9vE
K0OKr0wBHY/VvIM3WdqxO/x10ahzb3S3kkXemJ5deRPee5qvYFjpvrifG58eI/5u
R5eW+iiGF3WI9eIarlxkM/VQ3MbLOaAy3WaW7HDRHoPCvWhxv9rONcFAk60XRsaY
qp1j8Lpldbt9w3Yc986Jpm4x70m67YexhEmFMvfyuRO27h6h7TViJSCgYDPrmRcN
hbCl/OVIbi/c3FjO9EKX3DgVzIisFwOFKJwpyEVIBKM+MHMJBHi5Bvh3WcCmJm76
4IMXjA1yH9plo4zbRHigqPtiy8SJoZZ8cHrxeQ1AidckENQ8mLX09YMhAnbeyx01
2alexKnkuPZrzmfD5MV6fbZLdStrq9Ubep1vu+yCuFGDsF9SNBDfDXm1hI4bLSIn
3Hl5ASEY84SeCxyWjkBcwZHpZItdyM1JGEJ8eXIrJ2nZ3bNBsbnDbvEKDILQPV6D
Y52d4qWeHOV28rCJHW2+AhtCRF+ogNIjqfO8Q2I/bpHESAxPLwcPbZOr4itp+9z3
BOa2zHhqIt+7sCwgazbY8POKgo/24v+QmPhJDZ1TM1j2fXdWydaTLvG2EvuKvMMW
2+kLhD7bPAvsEiQjKVVENVTUmLYiTlxnQrr1b3oaJWqvrMO5zDIZ6ZVMs5ZTz29x
D19C/D18CP3P/KIH1ZM9H0gRpzC8HxD+xM4M8+02GVo5+E+08Phg8Z/+AinDJUvF
srvO7W/P1pRVK9ahLP4QHTj8auMkgkumIXngM/IREFzXJ8zriF9CjyV4dWAsfyVK
dOykvm1gbbouL7nWsXHm/X1jqBMt2IUROi2WI6bqfVyK7mqwMhfLa8E1XQs3FGGg
rwwAgL49PBXZ77IeFsynpRJNLb56BHcuxHiEs0WDx+EBZqqxr7xmL/eCLTZ0sJ8G
G5KeCEvdpgnHyt8mM4+bT7i2kNAMSkzFk2jrExmMZta+k5xrXdqAWLBx1DOrhPDD
K8OD8MjedDxGtcJkIJMvMcvMPMga9GgAK6BmDfnsF8etP8UFA2QH1qaFlfCigUQX
+CtTr6cFX+U8qyYmH+26crisQHSsazd/IcRArUZC/q5cShenQl9LKo3rcP/roNn9
s+xnU/7QyiMkXDNI7Rpu4j91HIUEPkOG8pVpySe3yKamdzX3TxSiExk44j05SMKB
0sfRzFx8jFb+2AZsDO8i95a5KFni5kFzAhXYKoXu8GxgbKsTGbHlc612vKMed4Vq
Oa7FMxGtORC2O4fs3UlBcad9KKCvwLiiiVP+5RTOdNvgYsU2Jx3vj5vyKo1kktJ7
JP0kK+eqSSn2f2v/If9eTVwIhso4ZpZXTVlBrExI6cn+s5lUI6Q/o1ty3cFTXclR
Mbm6fDe+sdlV7nGNih7OCZffYcr8AkHCp22nBgUtX658CWdx2kSkJY3A2Ge+WAqX
IgZxZGrbgQfgt2+I6mb3jqScDzpsaMpO7fc3BuMmygD4ZUyuaH+Um5L4NqWLE/6a
hyzK6I/nM11UOvZf7gj2G41G/x7R2GinH1B4RWemqIvO03eNWqVKL1hRj2fqrJV3
eAcIo9qf86EdB8+QNGHRoWAcaF6VIEAkSCibng/fqie11bdNwpUNWEkMgxOGtIRB
zqkwRF9LcjMZUe/HOsj+VCDfUJ+LjAwz3YZKQ63E55gSv0zURdtFlOKgSbFHilf1
NF4oNdfjAOtBfU/o7ylrA+rBl49mwu47JLJbm34adK2ll/T4F1nngMvnrAsCI5GM
nGgV6HeQrdHaKWs3C8KxhhN482GsGL79kfWcXNaE82/axqgjTFU+v9FyUxGVIZiO
WQxlGvC9K/sf42mk8Ag0aBHNHkIF0O4eZCLw0j/DdmXy7oEr6U345p6cJjjvMbCb
xozBK1JU7x0HZQXY1Dy/ewciTVXOMz4UAxy63mdyRo8SJB0KUWxtPHfv7fHTQ+FP
ba9sygq/mtyAEv6MeURl741zgHw8FO1JCYaJeUV1aqdxReqHSPzVarEBa2uGXZ5n
mJzIE0TAvaHINvuzFAscjG8CePxiyteb4Kh4nk3+xb4JEF2OQge6TDoDzEZEC/dF
FaVHLoY2Y9MRoGEDPmYUUt9wmDIdOg3ozggictLZMloXPhmnfp7RYCOYg2uQHUSx
prtqx7eJPrJOBDFiaAyY2vAMEVtI9k+SBZcx6CByZ4EwgeA+O7rarCags6+mqK0a
2Uyl04kvr+JUArYol1PD5nrhoe5dUH9CzeW3lUTtLrv3CHOPeUc6uqKYUz2r/GN1
XBtCkanEQOjJU6GI9AUsxez+leHmesw1pGX5TelTNDBGcCtXAK2JeHR8VDc7JFYV
VKe4/H1nTh0Ad9TzTsAh9Mj5CdeR8NvDV47yfe5IuXfokaFxnH+FVt0l0FM0nnR3
nOl/vuc1M/uSQCu4PA4vM7TKdU/GojdCDcAcFktkGu6q0mCglaxATg//HwNZEbvB
kipyrICljbhijtckcgMTL/VF/E2tCmT/hFpOPmaeUbHNCVZOgTOIpRd0ZhNbsNR5
yM9s7R1AwO7jvSWnqkP4qYqwr6qzJtX42+OZJ1p6RZyEAcnHWBNm5+M84DKt9PvF
wLT1H7uOovzrU3qcEVgJmU+zPMYMALBbIS42TCj+JflkG3i+9qUr2RHNYzg3Kt7l
hPVMbTowPwdWnd8eMKXHVLR/uc+ETxhEnLKvZzZ586qDd1bCAyIpBxqIw+gKTUgt
Kv7ap9w/kNqlGDY4JcNzZnSrp6vIS5C07beo7YtlTr+qzkOV8Gg3hXh1RDaIyPFf
WweObsaa1Cm63f47zToVurwUoY7K9FS1VFDI8LvSVs/3r3OyEcvFtv41YPchNqQZ
gDzbBxk8GqN8Qc4LsZUArrPlZoPwzjaS7NAN53vQygZN2YehWx0QeFqeYj3otKxA
lu7s/oM19yOi6iEoSnZLUCVrVmItO+KnTd3ZSnMzJ7HPD+V4Zl1wIm7ApjInW9LP
8wChfpRrITLFF4R0WVKJrGV1RUWAvqYHZ1lQ71E19vOq4pKfn0axpeEo4Kh2LOKw
s0KmoZMCNDZ2x3cUAz5Zv5cLZtsSLTvsuek3JW8IFq8dnCRAieCGJPy3Hi2Ga7Dj
RHi2YXiEAqKHFPjSv+hCGoMlmhonqbw9WQyMbgo/j9Wg+5Pf6NviqjnTdDLYqUe1
8MsVXerDbf0UMxevL2TGRoGq+XF4H2FhlkGz3v1bpyMV6yhh4fuwldcmv2QooHUe
xQ/7jFn2HyIGuL9wN0PrpFZ3OdcpG5QwVEf7FXtM2c9dId70AUU09Pw1z5kG/3jZ
XS+MHLEhd5V+FsASBlwgkDBJzuFE9wZ+r5YwqjeLFBIxGqzWT/CXRaVdFPvQQEu5
VQOVnqfgHxjZRD6pijDCF1y80uS+hr6F/SYT87BVhHIf52FYdyOyHyFviz2CcTga
G3B/NPyHfpSgDwNhfxIShQuml3k3lVKM282YW/GxwvTlWX18s2exApRRaYcYoALy
7aDnKYVyAUrgQfc/SEmiTANzAWNcGPU4yb6xEsw1p+vyTAYHGdpa2lZhjUB8xxG4
RfzrzTi/uqLhyJtqqAL4LS34qJiONOA7NrBVR3Xjx2Wsa5cO1/6v1Tkid6JRSMK6
C4XNJjI7swf89AZfQEWIukhiyupwMv17U6LWtToBOjL7ERfNOplG05I6yrMnMEc+
u1Qivchw4JTLMt1c0Yk0K+1Qs/OFctZCTr3FsGgcdtWqXP2RuQyPlNpaGHgwx2Hx
9A0Y18bMmr3sf7Cx4Wt6oUyvTg0m3hXSpgP7vxrRsh2W9apzfY8Jv3sx71SQ1FOo
suBm5MdqJopW5EMZlUxY4Mlt3/vXjjn5ahi8V7Q/1AuPbSRQHy1n62g5yo0LKkl5
27g+cfvDLbANNErylYT9OCkyeSz6LR+kYfBw7vSVjsdFgTdJubSgk3yAABx05gqW
I9wxKOlV1Lo39IIX8s2qN4PQVoi1ArRLXcqvXDamuSWdwNGRRusOPOzUf+FkOvC9
RylR7VaOtybqGlQSqiJtzYeH8UdidBCObknEztgbyXS2qsZdlr4/ouiF8YpMGRc8
BGOn8w6TOBc2u+w6KJ4r1+Kni1k8uvVPgu0HlbRviSnldAYs01YlXv79qKuyUWYx
oRUr8VexIEqEGiXYZDCjyKrS8+XIH+nVPgCrGkjh86WHptC92Scvu+ZIp3iVSOZ2
T16r25wu1ZGmRonLEVWK+d/baPXt4mL2EbLNeBHnkupd4CBqFijqj++yHehlfS/+
HTCmabHF/S0nvI8mywtfOzU7OFyo8HJAnz2KIpX4PXlpvqel6ZbmNrtlUbP6oZwA
V8Vm6GmFyDu4U6CXeM9F57CHQETDq2LiYLOwXy8wHVf9wki7jmrRNlzwUOEjTitD
ZNfZdNqLqDr0quIdMz+AOW8vRIMSVA8/iZT26zb+WjCWT5uLwCE0f3P+0XcfLcW8
Fuq/9xpapFt6CFh9WxME0lVLi0lodRmhegnZ2JJc2ySCPOzQTAxE64pwGNtxlYzA
LkWzXzta7nBvh4ptSLuOAiS1tFS4NIhg3FeeE1CvvC7liLuPkGtLygVKyOsgssF8
4xpz8rC044NbbevnEopBIlEhfSEFYGLf6/Chd9QiqictstPrJDCbDavjybp+lKwK
W1lFcuAAxGuscUITizUOGXYeiu0yWrcO/s/mMuUKsJHMcD1FwqGYY653dOH/Rqjl
5fFmRtc0Gx4J3+yp8OQ109l51EbgtIIWPUsER5VTDWQv2mAhboxJcnOWrYEwDteJ
sAZc+uUBUY4l7X3XuA0xURT0ASih3PZ1uv+KmP8DY4YXiBXz26QMJJ+TB6/PWcw3
2xg31gSw3RQXwmZvwwRIyjXGUBjViAKG/EDDUR0HfrgcypJCcZy6VvdQDWVgY8ss
sD/4J7CujxpbAud+Fjt8+I+AGfPAFDoKnP5b6YbnnQeIL6juZJtRHjHNzG2uIL1C
/vvHJdYRIlJ2XLbJHc/vkIFJKFM0BDOczqdZwpJbdqQY6nuk3pAQJS/0ot1kPbtN
iHl++4k5lBBr7ERK1AeuP+doMj6Tzi/hNr1d/8v12opT0NG5kXMf7kHaVBYeo33O
7WKTLzlvDrxhrFBLe9YCMHh1R9debJzFdhz1/8G+XW9lfb9cP2nRMJOyYTH6Qdyp
+WkPcxrl0ZqgP6RwvJDIC0rieGNrR3HU5TvIoiWX3AyAyISnOVfVN2nwjRyLS5M5
VasuGqU8QbWLxxCdw3jU8/uuxcn7xSD95i+8CI9q7fMX07CW0mOrZeHEMCtKFrmt
UlfRLHt3VU3+Ofm6zB58gmWFSrlXyp9j1SvNEETzEGwsmsjErqlm90oapnKgusp0
vQo2V/pDFFFgf0tnhyCQ1wLo94W9BWed0Yoc1ij3HhIo0mqmY5W3qI5UXnyXtzWD
wTV109UNe5giaC+CRb2Yr1mE2XCae9+U9FLWx4ntejeckY9uM8acs70AZVpk70WS
6rtTeo/kGWmwyksCBy4Zu4mTgjf2NtOwffnvMr+Pj3kv2ayxn0RnFUrtzyVc5xlY
Gin/TnJzM7Ol/G8dxb9kL65UaimJY6Rd8B6E+DF7EEm3WALNGwaOqNF5YIWh/HW8
y5Sy1qkN9JkLLzVd9zq1NzIIpiyKIT9mlQ+PkPhNDcEL49x3Tl340/FXSqCJy+Hl
J0qmXdErd4erH8k6o+3RomK8pK5KGWb48f3jDDuYYgwtGvh3/luhmYPA71UBbviV
0AJbeWJzgjHReUklbRzEhFbUR3QlGcbJNWAJLrAm+YEP3UodT7sUTfwQENzqV4+o
CzinxaoB+2rt6A0qka4n2T903zQnWHsHpdmRywk23dloH3ABTbJufl8tuccwJ+me
E1nvui7enPQ7BIHtBZPZ95jhk6Usl6A3z/ApSpifv9zBUieIzJcF+6FafIOMGo0b
FYAwIBHCGnPWVPQTjn0ZWRHTJWS/bzgCh5ZeDBbyaFCvc+jCTvLHse6joa+BuBa9
RbJM3W+4i4qvPaavVz1bBsUIixjT+iQmGErzPLwTVXUB/Rqnp4UgQrWYKgUysEsO
Yo7P1tNbgmPG2rqgIdEOERylmx54urcvpPE+RGc/8+tgastgWpQHtHeGU/kKjaCw
RBw3X1QIOs1GKvAvu0eRCmKQh7ZrvAi3VfvYEG+3U13gxCs4e18zf+fCouQIDCbs
JKcRYGvcZk3azWGgqLifiCEbuI7ZScMSJrJ1U0jyqvrzuQBztdo1ySMbsN47m2I4
vWVV8xpskXjIYpBW/UFG8wdGqYIy7Wt1mpnno8PsgLjm+FmVKUwKWf9aoW42VIPX
PBXNcSNeFIxdwe47aQ7vJDaMb0Hm/freSKE6ChbvcboAocUIfhNrpHvKue/QI6Lg
sqSY/Iw8Jo7lTwsPo7Ie/C5f9hd8wMFlqmMl1PTcXqea4rZBXQKLuu8v3eJZVPAV
VJMw86jypidX+4FrnWUbwxOix8fYTmYrLDL3QGhTU0XFHcr+rQCDjaOLpJYG0Jj0
sJpsX+2QbyAoJ7wpXd2Nr8pnV1e5QXH/isFX+M3kP+MZrgXBOkaAGU8nRjhdT3zL
bB2Vp2X3EI4HjWYuZFAnvn9Odwg9N+p5OOZzwc8nxj8C4qfE/S39/WLfzkXU7RX7
Spj3VID7582gCcg02+M9N5RsaHpk3I7GpuOj6yRLbb7UwagFpBolxwzO3JWPE7mT
NuVpD7u0OFq+pulZvEVRrglBpvLoEJ/uJN9QFDekmnU0/RbzuJioBks82g4SnLRi
gqsoEx40nQ6oILg4M5Y8H3A8jjw04OYwB7GVp3hsgl49vM2c3Zro2fyc7kFQrveS
XoCJ26kIMFCiacbbxNjX5Iy4jWnaLLlyqWeEh78VfbgDpSm7Dr5UwjDoERRn6gz+
gRgGVwc8nZi3RG/vPlCrb/d1HEbbuTWHGgt1Csqa/42+DQ85xn+E76jbBPRqmIOg
Re5QwgswC0wSR04E3YP6ATE7pIkjvosldx5Z+9O0iB20/NRtmqoUBucOft2IrTtu
P3XFAS2w1uWxa+PA17azGNDBU4f4FDzF0GXq2VJvIruGqoRP6u5hvlIG3e4W7VKT
LqBBEA7BNcMrgF05A0Y8ZvX8WmEIFJXgUKaC8IPBVEj7URGYSclGTHAHLqGWumRD
aCaDIHqrNGwqzcvxDT6FHMqb6OnkJ700j+pv3s28W/iKY9h2NXYd+IvE9SOhQDcU
yhN/fFS07hce8PHKs/9kOiS2KT66qgzAKqqgtRkvrXD49XsjS9UAx8cJ2Eq8AcO4
60friKC5j4YXqK/0VTYc2as7QbIAsKFld8/BMRNHxkQ0llviajxfoIzAJ+wmjadN
95zDhNB9RIkFmAUZqyBz8D2Ys4zhqIHyv9p/ZFyjoEj+epTPsku6i3DxBZyuADB0
23eHG73bqrd2nxp8avWbmTgsXqonczDf+UvwWK9t5XCyAVEKQpMx6PirTD/2vTaC
vxgs/OoR/4MZtGTGbF2hod8xfOKG7EaduLY7MnbA52U8zyhx9hXwb2hT7VYgBm5N
Cg5fXPoQKee6cd9PwqEzLzTBH4jyl2vky/XEeNY/s1rDiS0oQOuSLuJ83qrKNGMa
pYum3Kmgzv8OZqZvm9ujUhnWJtwWvqx5aykt8ksZWg9owhDIcQzRocTtild1yxjf
Acxvx44oavI2CxOhSZyx6qZxjkPwwCabt4bTmVsVWyV4jDqONxNB+x2A9JZb1W5O
Gx6J5xh+kAEYhsrTgbWe/se83IsG5JcoeXVGfUBPZtcqk5GMhPqo3WCRshEeS/P2
1cduA+GRQHjDNKcjqdiET2y4tKODva+RFdlZdrOvBrDeqZ2+pjoIvt0zflTeRbAj
sJuEr4ZFBMouFXwBp915W3N34C4X5XpLwXbotMYh1J2HAAn7dbvC8Txzlad3LcGB
tPAJTCFrpx1sfMvUV+xl2ArBk3JqZnP7ctfWB+FEZlHdRs9sheBTUPxhqA6emhT2
okbZUwdBvPFaW3vVgXcRxrox6QQpH1JJiIk9Ek7xu3jBg1HLLa+BFqMaCyikC7px
q+j1se3OAxL53foxpdZuxh6r2goZ/kXVHEOq7lBAx3hgvwA4tc9eU9oWoF0s8p2d
oLPvcZnE0NcfTF2ef2Ioz4lYYooHIi9wLLw5CKr8Ff2XqNytEfOULxKecCByiJ5m
MZIP8UVtWy54Qa6GbtI0cMrjl+Qr62Wvzw8CEC/yQ12DP6rckZmS9WcIkGW0eWwc
qFoP9qmc51nYNIPQC5TwxVfjivEiByVno5u2gCab1qWM6KD6NpLLzicE7nogghsz
3jYiz5FD5E6VFzEOmwAUw14c+JmtmXMXjYGiqxR2yOz1AW7rL7sxIGEBZBrO46Kk
Fbeqvs/OFm79OSx0ohE6DZefHx8TcdAZLR4aB+1wVvmTkhCXG4zfIZ0wWIY6Ahqh
omat6qEGDvileybUO3SD8iPiP6+H5ONLLO9BgidaeiF907ER0SZnCXdT5I3NOdgO
AQUuUOKx3hKWr3WaBiFKPXNm3nvvlMmr2btRxwRII4qaQKvbJ7DaH00H8mK6hgO3
Zr8XmooTRgRsvepeCikBdEmDuPrM6mKX8zsB4HrTISBhQ1L1wX0YEDCrYD2zRpcT
E/P5jHdat8OLNxCz581XD9qbqdM/LNguodqHEITj37tOsN3ljz5rJCJeFIYxEaFH
65dHnwvBxXzKOMOoIOIWLk61N7UVrFPGX5dSXq6rdOMgfkgZnlHZ9ekAu99ubnC2
CCNqQEPvUgneQHB+1LHjC2N4HultxEGH0lmkO9Ul1qEhLZpDjWc72LJ6Axc3b0ea
/Sf+z0YRG+0GJJguBGyQydUtQgU2We+UolLNhPEGn9GXxuVum8H1mjgi71reFStz
kDk4jYSocvbWFrBX8SLnztoFihCxmJcoSAOCy947mDrS14VArWU8j8bRC+F9gWBC
yHLsKPn9HulqfKvCew9qmWmgW4jxul8imsqWyTsbPlpbXkymxHRfwmpQfIv2T5By
iNp2MRz6IsG4QRczdQM9PiN9e3LejjCDSxmK98hrXoldRAbqVtftM5hS/WpcO3K/
Md9U0fRrmKD7M4R0OAA2sepnzHabiKd9PFDU7h/gR0pM6FPYIcVvCsJjjelkgN7E
swsTWuc35OImAptb5Khra5QkbuQQgypi2WodtJax+GrLNxAIY3Qc7D5aFV7y2z+3
K6q2LHC/J11AKHALxK0ePEZjKGvNJ8/3Fd1+zfP7bQSXWRDD4WwUb524c8ntruoz
FGgAVkwP7exZ8bJosmjPpmJsyldkI2Tn4pv0Vlfbpb/Nv1j7WZ6sLFbdYyDHA0fI
WojMgTjfbSp5puNwFeLyFVd0nHhdSjlaP/o2K7UwAiNgjf9cYqyrfp7WARZwMsBo
VQkRj0eyrx8BJA2MT3mQEu1kYORFEy3LP8oIJs7BBIWDNMeTLqOxyvyX78xTIO+m
feO9rF7qgGiDSQtFSL2Smrys87zvsjjEUNt3qdUfuBP0QjMoQZwr/jFMcVYQQmAh
I476/g3esjJ8V2LbjzO/pKolp7hQ9w75BOPsBHZnm4Z6byaiMEaxeivlDA1xsd13
wDB3smkaihryKDPFapjKI7BbQjz7mJHsndyzwiTI9mml07KbAFhHAAZNgFN5M9Pp
fza7CMOmm1IMWYtARv/ioYHkwBMHcdjZRHSe58eMJ6dB0URJAFuGBvFNs3j8lwtw
ZZrC/uu3IshxlRANpCWclNh+s3qJKC4u2vtILvsG8LJndsrL0grSaWw0vzM5/qwu
cuP530E3pezCLm5sLNJrEOEXxlr6Ru7vHP13R2YqLNtUwr3OLG2Z4uCoWUVomXeS
BFQisd9Ldr3A5kydpPVTCrMdek93YWGOM31aRf1x75CVwPgtD7LePRsWBHi6PtoU
V5SOOPbhQjrr4znpiPlAzaIW90vlLz+ZoRE37fF25sI14m8iTEWhT91GjuM2xA0E
rcZaaYWhIspDgPE8XGwGZYLaN49EtgkM6tzJKzv6wddps8Io3SUZIoHC8g+rTeVN
3ljz/m37JWkPW/UyazQ0KypmxWR/TH7gqVBdqcgW/2WhZd6vuzCddL05Kcyd9EAe
t2dvuxV8L2lIN1ewOKYYeLT/egAaWVgWJ0akcSAZRcjSV9ILw+0C/eK61w3O6B7r
eTjgb4rtJy32EqkE9Fo11NxxkX70J/nCgeJHY1lVa6CzhepWmp24dz7S2SZs4Uj3
sAxEMm2UHZ0OHYvc24a9/R4kx17xkSjs7Q7uMO6d1mTajU78WVHvfRH5jZt5GwIA
AEEWnkZlvdYu4bdZRzRmBYr2CinUBALgIfUEAs0umdafnELA16Vf+fhu35laJpBG
HttIh8hwilaDKIkwt5O19pe89mENgugtRz6Wa4M3b4UCAz+EngDEcz3sykmtHCj0
gyr0Jsrc1fnrn+qaeC/fOilWbNezVjkGt12TI56riLuopB9N+z3jvA/rd6zh8vb1
ziO/Lj9DKKInBx51v1t5R2K0lAPKS9NjaVurd57MuSo0gdfxPbRPj/spw+fv9pvT
nMhRdGLqLAAeWe+6X8drWyR6XquVRmQ/DTEg6VT2tmatBuj+tTaWCN+uIuRHqzZ/
9D5bF3OMshKiA87j9YGvjFCTD9MgzKixnyjM0lSdWGUn82yJ6Ml9siUgZ7m/aTk5
nAdBc/DVl6a3oPGxy0vSZ7FosRV4IuNkjcTdXy1dZaF8Xkc7DwaKCz21T07bfgIs
HCeiZJZ07yfOT1DY4PNltg5HWjYfDAhGbGGmC1xDwHno730IRIseskMWC9YhiROS
Mx5HhBk0TajV2PyItSphaYjPTopYDU9vhexwGQkdonLQaOcxSzhV2ZIa4GRIgxjg
UxkbY/6r8YQIEZyOqcGgKvClS9dTyu4q6h7k/aUiSJ5RzOWbxugsm7S8jEZfo8r/
OWE+Bkf4ULMzSGssXne40ijBsgUNwgFwsxerPJvn5J/TSmTcir/o/TgyYAXbTU3v
EIfYuQSVi/vHgrQVZ58hHPX5+kWOx0XZqYNtbTOuuDvMxTVHuIJLqU5I2AvJjFWg
Ff1u3wrFEgYysm4KEGS3ZmpuiCJa0CtzTlLAeHxl4k92CQ4hcLzRtrmVgvAH0bY0
9CBMjPB4IEMNPKdtNFPFV4IHdCvDu7OSpJ/IcnZcQPo8zN/CbcB8WO4GnqlokaVk
aRZjrKK/+DpCMWU6x/cMmN/G8xAJjWHCkvmduWeI5BGJ90VDdEY2Pp9WbcO+zXJ+
ogYtSTwlQuFOBqx4eBL39CmaR47LZmTXVxNfDJEnEaQPujMvw1wPKtnUZ4UQhTKR
Qqykeh3QVWM/Ya3aeZwc30HAUjK768nhQY9QyMFUpVtGgvNQUWcRHKCkPixpttmq
qv0nYI0gYL2CgFShnswRvXnomtFChSJKC7KDIJtJsvh73pIGWUe512DVQIRa0eI3
PuJvo2otc1Qxc13Y57Q1RdSHWr9xAu3M4CxLseioBLf90Ym5vGQNLkDW+LC2rfxw
/3KNV0ViY9q3fqGoZG7HQ/WVT/QNWeKEcTsrURRF4HGbW1CzGJeZqfGr6Qg9mzhk
z81YOt8M8hazfdD7lHYFRUYUqN9M+DyFqy9e71NzPHBwV7KO+TJieElB8D88CDwl
yYXfGFYYn2dxrfslVGq7yQmXR+CnGLDDRFHGs2kPlLZcfctrpgUDlVRnWS+rqK1M
zeG6w0Ymf4gOpXKXRjJI9eycvhjv6WqHr4r+DX54nneRrWnxLMawr7nbVbiRjmqQ
98MIRuLa1ZFdgpSSoHdeBWfUGA+dXH3rK0Y+T7pKC770KtP992xU+FEztpnUeU0E
TBI2sWsUeDZ4DU2wCDQZBW0tFfrbSYz+2KUSLZLMd4QZ6C6vTPbEiRqrpbb/93/Y
5jgPXx4IHoefFo3Ob7xBWzMYb73qjjt4Nc7zf5cVvT6J1gSDzvyXjxwPIUI+M2/u
rqhBdrWDYTQ6CvFaavXaQ5l4BvJ0xHoKOTAzpWZ0NRNJPek/uprmmvish4IcsloM
bYeveUk6eFLLyXsnnqocr+SkrjusuGirskSLw8vE7Us7CppBrH1e8x90EtsAlEfx
srjAKpgXEGyMVxl+UzIA8KvEDbtOr3vVqodnAIBxRgcbJZz4TdTAHXj1wt45n5rI
ObK6QfD3QtiUmnk5EjuwN6V83TKWYy9+DtwjkE+TxV+1PYPU91MUs1VGCvUO7i0i
suGdHtVCJbL8gcR32iUAccqRZ9bD66eZVStRDxLAq4MjZg2figOVv85PDIiBOhpK
IDAdRUmFzJCTtgG8R3ohWWV4mGQV5pHYWuY600n3UpJbJ8Ub6hoe2aaKXTSo4Ad6
mnTxgrn4h4QD6Niw5bo2GwKJAaB+jO5Z+sDVZwvs/Y9Kftehm6gqznDuhB7oQcYD
n9/HffXENVxI1kK4b+/2oP0zp0NWtdJc+vdjjaclrofZ2rzCGRJa4enrsWu3l3gp
je0Q9bcVoJA6CHlD1F4Y/006YSGk0u2DszymXOrD++BPD1iR43wUXrCxseNtfX8E
cysp4NCWcDT6lPtJdYA6x494tTHfOiEDtWdYocoRtosYUZ2GWpP4B7vnSFUlmt0b
8JUReR/MEDakTBPlN/dejenk7d8VfaaoW7ms4+t4YmLeHcgYGWDbBV2F15EJP2+/
mnptxwYVTLTBmH4B+RuyZqOQ+LkwqRlrIkIL3VLPRcw+1hq++w96Fu0WupaHMuPS
gKKB73VkPZe7Q2b8wPOQgm75kbUE/9sGn7yZAJkCVXNyi0oMYPiyqLSpfpuRZGau
jj09uoLpV2C+Svkuhg8c9gdR1/oFw2gg8ZWNDLizZg8ESQ8rtZSLGx0ngWcDFg3G
mqYTEF+ZrBrKc31a4hJp9deDW5eFfStHSrowdKloPrlCk7Gy8LjploavgSusgmIp
iEf86RRMxbf5kTQ6kzeA6Q5QtKGB2Rwpoqkhu/aRlxLWqK6exFSJlEuQX0VbaMAJ
iAFkd5GCeXvYc9ieEz7nSUm8xi6Dbvf669t47z7QuAvdz4ECLoEq4mR0zN5s7ijo
OXFkBZuEVHRrIQenbwGHgKCiOFTWYp1Rbm1pqL/o/jZhTSzRXqlWn7wlKQeNIYjQ
AZqTBJRspZcInTfw/wfvRJYQv2Xc34NUFZRIroNRSO5gJLAVgCG92bAHF1kMRjX6
InFxps5Pc/90WFqwXXupR5PPLrXXnEUW53C4Ycl2N7Hzum3HPLbanAZhIQt/AoZY
MDSLNUIpCHQxb9P4Ml1F3h3aaA9cAdj1tnheWchXFxzYJc/Su80PnH18/AeZxoZZ
6PFViZldrlg/ZBQ80qOt+ZEvziYWIJoyidbUbnG7fxW3KJGLirBpNyHzSJrgJPFk
lxMYDVsBK+GUybPgX5e5RNMg0pQWjDVEta+ZMvBLjsy0Q4A2wSP6mpEsXtazD5Au
asV/G3uwPO++sQpBBtSRbAhhoXJmXAKIqq44daatw7mNxYBVWiHCYgMiJTiS3Cdw
qK3UzqDBJxuAnlkGLeH7+QY6S/BghFwhCbYyJ0lXaeYgHStu+Ei267O0xnb3w90E
dZMb1LpLigAM/NvOkn5mfTK3PQg9Hno/QfFU9ngZDO6gf0+Mzd/hUR/V0b6/SpWa
BZKso5/pgftUtFQdOkO58tucbvXF4L0zxsf2sVSfOSXzR9pSLbWJ9eBp1eqeuN/q
HFJVfM/8uJfQRuzS54YZVbVlI8xwqEAG0fEQ9Y0SIieotlC9+0IrEqFo+UczLlH3
1TqmBCSY4krbzF4uA5gppsy2Iw6SOIg+dlAtC2sBZhZUtB2GzqSq18bwr+w4/S0n
TEkH2PDWiqol87Nx0xI8PSY3dhRJR8Us+6mb3uqjaf5ADhmSmJrCq4gLdySn1Uf1
3kH6qz0SL0Dcvh6xpzxMcfNg/1PrWPc/1cSrWMx7mwiNPa4XRnISJwRzuVIUAQoA
+0ppWlyktD9ehAEefGsBHA04nugcAKl2ATzxzbBOLRiImh6UHMNXMiCi6fy6IgUh
IwHjhW6nWPSHyzTOmZNNj4YwMR/xdEleT9PiHRSrIZT8/21Lcnghc1vF1AohvpzY
u8WX4WfYAB8DFCNcLpsxoiQDTRnIOKH+qrTJec7AYcZ7t4NWHVJpAzzpL/DYuOoh
+5ckTFW/5Drwhq5K73yAFD7xUWcyX+CAAMGpTu9HymDZqlLGrfVULRyFgMGOMzmn
L2Sn2h6gK2riejk6lozluZFuEG0KGpy4GHN/9hJKb+ujJaZkxLWYroLp8NiPanyK
CJfMRpkPeUxpS3kdKiCquFV7LtyOAcB5p46YGeipSsq1WDTeV1mljUwlRC4RISJU
+zNpEK7fHjkGGNaeygeRmbodK8wvy2AAEUtDJtHB/ePfvqOaxUfX6a/QYL8dIaVJ
6OWavHlJ+W5WOCMQjjTxcqlXIq0joPjXbiUtoOC2tRp9plMKEoUrXPjmLy00leX7
JgVQVzCsB/eo0xX9p8G7pWviWXdD3mxRJffDmparQgE/xo1O7H6/67NUS/0V1ciN
OdsFc8+8bn4qhGR+iGUI/BQ2SQLtTbVh/rbKnxEwpTG/hcrprw/U7lYebEGDS5f2
LRCnOTDsBJsjVPJ1JnE2jzx4s75ze5bcLIN+IX8ZfGIF53wrI7b401x3zXVgZYbX
JhEICyq75R8LUl7jGUh+Lx6itKjGDxgeWKfDdC1DC2yiUvWKyD7Q8rbuMcI3oyG5
1sTU22GNts6YB/c5o6iWibs8ol83ZBZXjKo5d2JzaNrGh9TYs57OQdCBDswisj9X
Y3cHitm2DX0W1SvAyFuWrB9MI3msDyWhJ2x4xHz9O8/eSQ6Ifj53hTJaPfEqVkKu
dPoBwsNGbjiYR0+Z/163Tw2plSwi0WiAkWE5o3CKtfyaAyUZoGaJx+0mjFdiuffi
cmZCP73VEvp10bwXcCAGJXDWmIqIhoyYX5AOIhNQRdjp8iA6Wl+vdvnSVc41adLM
1/zjSa5I2WkCNWqCu4mvHN8rnyDLz7NnOYqU8nK2J+xNl5khy5J6xtsUYHKOzAuH
dwCV9Cm4oOvqzCCFgUKup3VHDLEMP+lMRMTclXRX5AXTU5hdWtRmJdmT0uAIiKvM
yqjFDqVLjkIM50IDIuKgCi5PPBFMi8ognWryorKQy82t2JKBFiQ43egoBNd6o0U1
hRzaRUnJam+pTzSJjA1viSucdwcieY1lB7UYLyhFuASH+BsK2JguhA/UEI9vr4xS
1RiI2jkmRpeAPG93mJSg+jCCxaL4lIhXxOxKXXHzzP23OjRpLk1VzffSbQ/V1eOL
8AHnkDa7yg/NkDHcIqREYqHetavXpRVvj6/JEqkrf7oYBlj2BtRJy/vT6LUYwNzB
DHcnb0HfzeKVOkZqsH0gKsjUFh5HIuaL4R+VRUFs/mr/unWaVNk0DEjO4UbBzUIs
ixjndMOuLdAxyBVMEscavtYzPNtMNy4L9iEwb+F3QxMTF6hEmfEHSvh9nl8KfxPM
i8kNnhlFD4s4EjC77RjIAG51srVm+YPsBiXH0YPXenBJi4gjb62XuVoZQ6IN1xF3
7O45xcIF4IexgpM8eQCxNlX98tKcNUG7M4CvLTRBkV379/eacuEHY4A/AC6KiJgG
d8ZqWMNJsml8yOKTgelVLrLggmr5lLeOarmcHRpgjRLPK+BRQJ+H6JACRr4an+ck
yFOUzXSQ9pL/8XM+Qi91GA2H7LnstX4fk8tuUVGqH9PeYGcvukM8NrlBzNQxkp8a
mYHrUr4/KHuvkkvu/lQ8ym381PrMRwvM5hmEH2w666NTYH6MoR7RMFQCmZgqrVHZ
vWRmRdPj8EXIEKj77xRNdrLLGTSJv/IeshPrQNQLChraPBz3Rg8wADmQiZL1jCnd
fCecDBVVbKCDceG65UKQg0Q79U/AHV9LfrC+2j2SHuBtn+1HFgupKVk//KTPaO5s
wjS5l+mQrykSsftPaTjPO+kSt546Ws4NS5mXG0isvSLf+0QkFy6/gF0bpQWbDh09
Dj/J7OAn5hYsswvNf5MKseA/UK7JCKgq1lBZdqSzKz8QB6Yaj13/o5j0qiZMzt9H
/W+7iuhMlGrB+KFfBZCgiWe7gjpN5qJyDiubLOo76HaFdUGvzxMCrxX8sIRKjThD
/S+XXx2TNXHfMkY9JVKID/XJ6CvHRzN0tAjy6TZHzxxr49tWN4dfLkYuhlYiCOBF
twg6QKMWT9IW15CrIxpiJkmVji4F8jBH02Islj3rOY3SPN4FBC1WzRWhSgYP4wQS
wtBVI97dWHWHOJVtScCfEK0ODVyrg4v7J9UB00mf+DNXk6ydiXsmPxso/XK3clxk
hojzDpTwr/T9AJQ18AhGEVb8vBSw54l1fL7Sf3+hQ9N/MKCitZzCur3TjSdypg3L
p/PBdGVkGCcp78hmk/JG/FK7Fn1UcN+iV7+r6a+MOeauYdsyHA0mkRnq1tt5Cnx0
thVlf0cyVcE9EBEKJMJI0E+9LYVj/9om5883097i3EP8Q74VEphwehef6v+d9aOE
6zXGmFHeMN2/Y99NxMwZYV7laazzgC2fNMrRxqcVJAa3mkJuxuWpXVB0XvSbP+46
Rhceg/LWrjbvz5A8X15dsDZK2CWMo/n6fRf7BWC0tj80lAT5ngm8IOcwIsqcVh0U
qcB/aBehvnovIQPD0Us7GCgHuRT1GHxKBkAzLCSsVoQVQp+tgMpwVOO/XzYI3Evv
7ng8VPF1Tgc8RfV7aMdbKCDTuaVffL8HBgutFU8mxGN++plWeUVVO6KtwWzXitPf
9Rx5xJ3UgmY9jNJPl09hFerlcoHxtWpsbN+ct5mSj4tn45qbhCCBC3aaIPz2ptUN
0q+eWYvaaqQZUThctvtPuZvrIc6OkCRxfpDAYM4m69HSYUx6PSl1Q/wf8QzxImoU
Bb7jOidR9DpOMDILAyP1ZgqihnBg68sHkq5w+bvgJH2EowwTastgJHWHzkSXaqbU
knZZyIW93x0tgoNa4Zf5EK5I6oNB29dzL4/W1z7B62jnxjBZ3Xa8qFHCZosoNL8v
QYhUB61CF3JyNlpm9lYvoNe2tt145cjU9t9Bi5oKogE4qzaKUv+u0c65L8LkgPqq
mrsnsi4/zKBpnaZ200l6Ngg7lgAo6Txwkvlg/CCnF4Vi+Y0T+3oEhyTkxTdlhoo3
vppdF6cssGxRJkNsvuep39SU0Z2ozOrEHnXByMD8jDN5I+86awn+ajKWckEkuqlP
H6ZVmD5TZxZ8zcfkoBeFNcRNUnkE6N9Ist+txJL+gkpfbr5pVY5C8K4XUz0WAHqE
SzCoxSDba5cDqcfQMnYMwITX5jbG50KrNZuugbyC/H+mseg5GNGvPLtuRJOdF2e3
MduO/x3ItHClPu8/TIChzOgmIKtdXn4ZlWsU0DQeky5tMCQU2tARHPhRqmcaaLAW
iTuB9LrL/+3JhJy/wJ1LptP6ZzANQC0myITjF8Q6AtbzEpHFMatrXQS0XRMs2vLr
5GZQzpkcPmhMhicVSpEQWa1u79sc1UbA922G7tlplKyQJYMsyspyfTfn63XBcGUG
90ui5SdYgpszA5ymLqT99z5xLTa+2V3tQFpEHXMJFgenFxucVFhGSIqiMBMjc894
Sk00dF2+rzwtoQBm4VGCSXOW6rwG+4DTRV/wk2pbXp1MJMafq2u+cK0vdd77Pe06
g+Dt7l9R/O0mvGslHFwCPvMLyvKw+ucMkc3kdYggwBEVH01PPaEBmcuzKKcmjqm7
OuQmgG4Tw7eRINIsVy0gmdY4qM+HlJyCQWlp8Nma7ufMfgPaoYwUuoYohbsOucL/
nDRF+/zSvP+X+tQ13VAymjKLIWaAKfos5bVL/wNo7X6b/rQSq7da1sSVFat0uSLo
yJ+DkHKzUxlSTP/sG0LnbOrRvSZuvVXOtpvuxwujxHv7kIfOl6OBGg5piRXiUh+J
qiMtxnIgSugqKT0ApPBB5A6FX5tzVChjee2MDj7F7++OvmR3KWTOWZrb2JwjgXil
mK+1mvdXLq5OwVmU6l3iVnbKx+JzuIY+i97j3Ndf5kj22ivuchqD82BIPpsRnkp+
tu/eCTg4/GP0w/Ca0a2nOgwUsqOnGJoTC+VKjdJlwUJgMGyTYciqaz7XboZuqDLI
vUBwRkTfRS49Rd6lv0MOOMb8CddXKFXznV2zs9lRpiPE3SP6e5/dseQB3MCZaZn3
5G7Dm1nJLHCusTj2lSjlgEQUYeqKfdmmmz168UfjKHSdyFVVWE9LtPXvT4QEFg/Q
8Wwf1yZJeN2p2a9rsluXrVhGqTaW/tjlH9Vi3Bw1+7hVRdXAR3n958YuuL5Pw5Zd
pUd7HYyDy4KE6oIOYjt11K1chl+HkrrnSOtgOp4ZMcqP9ESDDMzkLbub0q56tmDa
lM/JrnT/oKQaybSGsEehLvQcjMN05uVD85TgPrnhgslZT5eLbPLwtqG2WqFbaO+x
niIJrWMCZCswDQNDjDTAl0Tr0CLUTo4oj8dFKBvfoUoptG+h36TbFG7bOZCtjXQ0
irgWf3kStKEiWRWg5PKSCxZr8D2wVQhE6pWWBLVIybEyxyw4pMRe7jkkqqDZsrCM
Fc8rDvRopMCm7KDSrrWfPL2V/AZMQ3ktGyZwf4UPlpDu92rcLkWMbdLbMNwcT91X
jSJtRipUzoUc8WEX0LrAi9c4w4VsAI+7sx+mOD0l6M1RhhnJw5cq3UI3GkQJvdxR
2esUrZt0+25LvS8wmbEx3eBUhBfMwWG7i7RIRxOdVF1B23KV49VgDd4ZPU62DRNN
QQ+ACx5leoVU8b6ipVsAwHBTV7lUOM9WL7xhSDMGcnm29T4K/cDJIgatoolp3se7
jkyBK078oABvfUjvOlijqhnS0AdXirIsX73KUKbSUyOV3prct+kikuddidRM8AlG
cPQkRGPMn0h5Co5XZf8lunwW3Dx8HBkJC7/kjqJIa4R79McM+gTUnl+cBS2pL2pt
lLJBwvm/ufViJ3LJRbwkNg3MTTgWumr2/ptrppkpJP3ajMFjqbrtzKx5hyGjT6nm
A+0GIWnr5qOV0yKmruPowSt+Jes3yPOurzStIKMBWS3LS9yIn3STjHqX0VovkZzM
nplKAt1ZwLPtNK9ohfcP+e2XcZOqP6tj7AOBwDjRlgyPcgMzl+rMwJPVh7zaQ4Qe
5bW9J1vrJuY4Vcb0SrJTSkWNfcdvdB0UBTRk0BvYSE38DAFKIEcenHQA4N2/ZJVh
I28wJuLZf+KCWTpCxGDadpmCbcpwZMibz3lu2FI5gGw5ib7xP49TidAmMnZcO3ZC
jFnq/iQOfSMML+EDxfyb+7SNozclrlwvKgznRHNPyDWsd0KN0CksU3FZBy87sLhE
tx3Y9oaqodWdF1YfQ4hTcuUKl48iQQYOUhqzfJcfnxkPvbohd1AyDeXh8dBMVMvF
tsWTsn09ReC7xW+i3+nY2Hy/7NcdJw0dGVgzgg48vTELA5pRnStajDHaTehW3Aw+
GGUKKH3OYrYyE+PjBTrGn521hoXwEQ+KDGcY8V3fqjs0zHl2qZ1wVRgktecgMa8q
Aubxxfvv7KLk7f56LxwGxJcwdu+KSTAQSYvBV0kw4tWAyz1TqmCEf0pkzz6WPWrS
HINHXkDTP6y1DsqrzGkw5rx4PEiBHmbUtc9hlZdabt9rJ0hm2mHgCL4Pgeiqx9Rr
LXAWYANRu5ExVsuhFkucKS+t0UNSHv/zdFQHKb/VahynjXdK6TE3FvW+rQ+khN2e
jZOvs8DfjsZTsD9dzlZXRM7fUAOYw2sxYK8Dddk2FbOp1cX6amwFwRt9+maejHAu
JBXickK5R3oQp/eoTvBRymgXIAyJmk36c2sdC0H0SvNWfmaB4VHwwqYRTCl9g2f1
HJNQvZ1Obavpb1SIoEwG51u4y/aXfpUAMsDRSthzZhXyvrYRDe7L7NUqImomclHO
nU7K0TyrF+7sBYKiYhq2opQtldDb2HXFMsDyb5mUoaKuxR9FRL+BH15VsNGyKZ5m
+7dGSLd4F76rHsHLVnkojEAJVmgDRNnvuHHl4DJz0NsndopKrZNQZmb6xkAN2KdH
XvY/BLa/GPa9Oc0kitny/fHj6IJUixBZmH3+Sp7oCHTjMVtpmxHPT2d2KUTlhcym
xFBzTW4Hjki+KBjBivK7mM7IleZmx+7x84dUDgQXvTlrmaWVoq2gjHNydXBmNFx1
nKUIsXf3XtFR5JZnhVzCQ3wtHAFtiLvNgnmzYQHsxyq0m7D9D7mScYMHgCBO5huk
ILyCdx7HwlPJjNH8k/Mx/srIcURdZX7tBHLKHYI9kcgo2zAYhVlxr88ltjSL7T4S
ThWsqLkl6Q2yS8KKyDhdbCTctxjk00PxBFADj9Gi6LgPTKa47hOnSQRndDmflWI5
YkzdnRuNW0uiKWl3WaktY9PcCj5CMX9dbBU8tY+No43boQC9Zh5IxdpTt+n8hCyR
jG4k03CFQKpaJLAhjlpG2ecF+9crsa0ErLcrfRhRT77bwwtZlD7K0GMfCZU2NWQe
mdijSl0rnF1rbmtxMmAmnbvky3Qpei3cNFRCFdZZj5e+I3XRaHUdk5Z/lLRuzOlx
WkjlUtLUcmGJaJ0Wp/RGZl+UcA4W7c7LTaqyROGojgJR+AZFSOXXTEutjl2i6Yv2
KqRApG+uCnjTLFQxtKRU6/UI/K6Q/c/9gClBBdWPMgd/srP8NnEybCpqIek99VgS
g7IgMGlPOloKxD8ITSZasYZ0S2a9zyqVCZnxGnIRBsB+CH5XpwTTk7HrHSXgqYT5
ghRaKeTIYxqqiyX8FLmqPCY55p4xQqKfETOXWf26Jorp/BcVVr7OIM83SQBr1P9U
RDFcTWpm8mxqXRzjpabjOq7rtDuAEsoYsq08qAHY/FXPQaHRcq4R6/oB0BGe9Wsf
nh63BQiBFCW4fT+RWY5oj1o9d5UZ/C6JJ7cdnByxW4g1VOKzPUNGn5lu1PT8BuCM
8NXaZE87d7kIWUuinGVJL5xgL/aeSGKOQv7KF99fnYDk42w1k7kxY5bWhdB9p63C
x1PLWJBIykiAKfdQXF0KRqFx5JybBg0WOW/Yp6SdEyE0+pbJlIzPdZoWQGy2JesB
gqR/wXKPtUAdqtkmOYQ2+awCBn55cCAox3gJdLN3KLmHiUFOUo7Xq9djv4Cf8Mmj
rv1KypQoH717Ks7X1RQ9r7kykXX1egS/IYzM40yVGCtqewrX2A/mB2fBC9Wy7OUD
4i3SbqDS/gMwVEohHnTx1ZUerVpTi9w2C/kI+jnSPtyJntiLA3WIaKamJ3lE4txD
o0oOwYuH7K2AUh+/AWo66jTvJiUXysrsajxnTloiSmdVKTVjc7un+JzLavQOG4qq
YqDfuJCxSfQyVcSpbGrQBnUod5vDCU2TgPayUgVxzU7Qa2W9KuaryR8hX101a3OZ
DcdyGWW2viTU0BilVgWoFv6n++tQnS/nnsJIOXWzEQZ3ZeSiSpsSS3D8QcwGY8U7
p7R+YUCNw+24iowiVLl80/pfzCOLhWzSruokLQqObe8YHT+nS6sssj5kTMmrV9b2
KxTBFSwM/vbkn921a0UJDa4GstG4HhPKmQOW3ioYHnrYTXU0O8tso80RrTzqVrc/
NWy/OnlAG/3IFcMQuuKQA8dw10xfvIqAF+9HE9O1Hk2YGEo5DPJoW0ucHQWE/ATF
7fXxpLu0aNBCAPI3Ru0txQI/2DH3gFzi63ADyv5JEhj+gAc52ritEnEu39R53iPM
7+IiO17q3fe7zZzS7C5KLpq8V47yqAPDa8Wvye7T0d0Voe4UIE+tyky6Jt65PRmv
pvsIVOeojtszXYJaLaDx2YA2nuyw25TiIj+ebWkgMbZS0Bi29Ac20pSp1fj2kwiy
qcmspEbNX1s3IlE9N743W4kVqOU47y7/30HdRprDEtPDqF9272xsZw75DH7/MueC
Xu+sXnf5xds0EpoZOmknHqKCj1gePDzUwSLBT6mL2OYK+0poBeBlv4dJZbyOZZkB
1jxXNVUNJ7kPArJ/CwzO0ImTpM8sJEnFoxPIvSfEQnTNEsm8IhcAWvBTfJXtXDvh
Urmu/TlWfaqGijsAT234sK7KcGhPj3LA8sNKgrKPR4GgzoAWHPAN1Uyg/0ub/Ay5
dvMvR2RBbeu0d76xZPzrsTUhNnyS3OCs01ZakmgbeLtS4AF5h+Rfi/tGUGjAPXIN
1XicAx+aDALKKxGkhWlZjXpuBsnT31KuD4TEk45Hmw35BP1LF+GEzuX2o5cb4Y6H
aajiCSPpzZuDPE60NBWnMv+Ryt8OFnjbFjgGYVuFxmUKhs1Lgnqm8BbUqytfUW+h
Zn8ZYGk0Le2Y4wz2FI2M/kEkaMRo0IoeFJKWWSnA6FIgaKsMtgDxE2VIg9dS8QON
DUC5+kGc6n/I4U3wVUbFIcpj5n13b2YWSCHkORmA3XIxt7h7c2S9DuLtA0CO2rFs
zUUZld/kz1I1tpmnHtDXITSoPEI8oMVSJhbQxtl+c7XK5ODFSphIn32xn3e38kDQ
rlXo1p00ONZ5EhqLqm7qwhm1lq2kBKBjM8D5w9fUM2ucrPGBCuGzdnLqAZwcGkEu
DRHldnGmYM0Uuj70zIImX5FKLfS62imxWisr2J/0yUvsg/oOkXZ+rNdgkT2SKCj4
CP8sV/rtK2US7ji1g7GEWZc7o1LsZ2OmhXGnIFr+CZC9on18MaZm1Ws+VpwfydnP
dNtsSZwg8/tqD49ct+aEU+BWu3ueob1jRlvWHtYUgMyfAT/2KP+BDIRpcSsV2TQB
2u15GyeYAM5ITee9Nq6ybGZpSf42Ngj2QEod/CJdSnWjjRv9ITX2M4P3KNADDBdw
iaUQFRERMIct/2MMYFTQ+1YFCuLhgo+hbW1UOWTDJfYXNxl5d+UpOh1sjA5UCQwD
Me844JXLnNTuyKFATWJOZnOwW/KklWY09sBvYc4Jdlyh6ePMVoWRDIpxE2tR4kFY
1N+aeZVp2cYbX9Wb5bxevYC8YDvKB/fjLUoYFl9qgVuDeKl8bDhjT0qE34AweKxe
E+7Bf1P5SoZPzUS6b08jBc3s6ELFRbGH1P315Fa6mshEUs7licDYmHI/iqqMNcvN
2TganRAbTAPQM2tp3uHICjVF6NtXCEvYlyyc3ZSadRyz8PM2RuG9XpbDvEptfNs/
KsHoFoGCkYFBYTL4nd7rByEsvVjZ34IXVDPcOsfgpaVDH6KUJvmAuNeQ/4ts5t5i
gPJ1uUyez+OXiXSYE3pYlADIOMRbmerXX5p04Y9uVSKKL3bE5Zlaoid/vGC3ub3W
fo1SD18OQJY6WtPKn5nFdtjXqA1cSZiwJ+F2E0mTGLnZcxCYbbkfByv7ZR/MYf5z
Cgow4MCyJ/Ucve0FGspzMbexVUZ7kkEMR2Nd/aLPtuPjAOrw97L0AOfeA34yUjXa
hbAdPms6fq2+27syMF5OtdTRwLrl3OcGZYB5nPKxyRpAMDdhODn2JVLkm2mxtUpp
I6o2YHuH/tBXZMYfRQJoj5iyNyCcEU2NyUxygY3J31mQnLj1L7A7snYTWTcS3w3t
EKpPMCrLbZ6wNQLTI1PIHO0rEaP1s23O1wPu3AEydETf5qi5xCuZIHagURsaA6N9
m9DFA9PeF/4WJ3uNd9XOWkdl50aiYqn/0aRoYFjh+ltQediGcewwQHch8FgZxyKM
jLTHQ64a1WxeSDshP1R/tG9y+mM6Bx9XzOKUjYxIxzw3rPB4QXza+B/uSJ1FK0QR
vps9MkKoldiZhG/dIcf+x7iQ+BHCoSm6LOS8elcIWtb3U5yOHU5N/TjdGTdcFYem
R9rgX9dUioX0KgfMvVBxgMtOakdK4aFj8K/M9AypNNJiG+bI3LFux6OYkB/CIwfx
DUQvLnvuPglhu0VYvl0n9OtpsI7ToDN3Tx1dqOtRxuIYcmZhWPvq+W3KoD8EaK/X
eIn4s+/a53wzNmbsn59bB03fV7qSHUFLHpdlN5uFm1JkB8lhvRf+8TfuanpUru36
BMZRt7VCiQgSZAeqaw/u0zXsk1sC+ytIMqDtYm41tNq2TV7wDWO+2Vv6QDvtKn+9
RAVyC1ltbyiRjAf8G4CTSqPdXEyEziRZoTTXUAjaUk49IMMa5NQHP5nY9mnQf9p4
yTepL5DiZZuyTtz/aaZfncPUJdpFsuZaEfNUbYEYVFHdsyrbH+9uNIp0OKKj2omo
F5te9I3IwNivoWmrzSoELRBuG6EsnoEpLG9mSq3IAAtBIL2pS0a6ioS7LbYxXlOx
PhR0cT2SPFg1gHCg8TQHi0DmNaGd3K28QzLlc8HVzyCMWXXPtfzpkb6okBd1XMvs
gDMM5wdw6yntIxkjCxUmQaOI/66VP1Ve3HShBMctTSMGQ63uyea6RTec4/zDShbo
OhCIv5yBmmnVUrVKOGdloVKwh8fUKQjycSi9LMyDZRbXRooR+4lc+XS7wdxPJuK7
TxT+G28roKxuPfEL0RXy50jvESt5kanxOwZmtAMg1PCNua7LupU8zUfjEjmgCDjj
gRGS9ac3EnwFwB3O69M349jEE+4w5phR1wIpT2ZxRDgJ1BNSt523f73CkbEjNPav
BuzjDpoQGlH7KPxVEHv0/A45ubrGOMl5ReD0VEa4ScLz/00NXkaMoZnm5jTZq1TE
mPC8bm9UcdiXiSIEcOg+ok4B/Od4tH0mrmk3xIsQla8SHHyKYMcF4vTKTfXNBz56
PLwN5Gm1bnvO614EWt/5tUbtEw30tPTuj0JmrLQ0jhex0s4atsgwYv4fzfLmtQvu
ipOpK6Cgn3KJOyPfxDMLztDY/KWOrx3gSjtMwa7UdXWFewB37JgmeRoGIG7N4gAD
AjxUez3oCvrSSQkw01sKe9oyNa9crzNXO9c6dcJ5zQKwCW+9ySw1Jmg986K/lObJ
W6WcH2V01XL1rzufmsfubSy3Aaif29H1xMGpPCN1rYGf1PC2OSvRrGGTJSjbUeSw
zXpqu5d02bppaVnoSv6cgDZjShjKMIqt/PWruNUtGJDZmHrfmmHQRucXFWT57EMh
+1ZzroQPGd+wuzZ+dx+N36031Hfes7qwF/DAGQBP2o2VJRBmrtQlfABfJfsGdxW3
E4E/Ny9yEaK6mD7e/jPwG349L9WUQfTbjyBWavZzGfP7MH/ROG1r+c4/UhHoJ7+D
Gas49QpXzRYOXf0HHNeN+AjKp2JwxBUmfcX+u2RkAb9AU5x/TewCcZA9afthYg1+
6KjxPmKoy8VIN1/8kntnkFSurCXCnVaukc/e2rIq5UW9kdByRrWdzz+qZio++cSo
2T27FgaoowmLooLWebrZ32VaG3OjOgUN5H9YXXvH2bZ/KdYcFQ5NKIspGN4bRa/z
xEZFs7VWaAyhXF+2P5oPBOFXmTnG/JojSnf3omS0feov+dV9CMHmA2QcAR+KJzxu
ShKNxDGz+H+D5uCChm+U5WzrTUT9bQ3sLI6sWdhOYLIX44H9Zlzd02dMPoAm4xwg
+bDu298qgMjCHrKcGeg3eov+8S8BIQfA4XX1o0Xcn2bXNaEkVrVwPRuireojUYBe
j6nwA0xtI1iR/n9yiawXRrJRME6n6wbrYSL52MLe+JdN6pASDIqCvPmcOOVr4xbf
QM6QcJjg9fsDTTn7FfeXJep29CNvpK1MKYMTFeSvRjttzv+tHqRoCbAfrwdGAezl
bjFpR3fnaaJuMkOm07gZCrUrSVN9lupASJXzttHGIkFeDoDJxkiexVZO7y1O2+AJ
2rbbsU4abfznNhfFCfmSkBFmRbqlt0pkNxiX4VE/VzWLCn/aHXm0PhVBUr4GjgaF
qxhx6INGoScYYd8TVVVXgH4xcU6RuPeq2zc2DPhkpqPYTuGUJO5RtLmVRE2oB+AU
9q08GolItOez8aKi5g/83PDvC/XOzaKrEp+bRhL/H/x8rIsgOTaBfVR2oJFSxaxm
l4CXZ5lVjnmpq3CLsybLJDIsdZJNna7LuEdIZnFWNg23huhZoTseQIAWJng21+pi
hQoS5t764wEInzbK0ptMa+to2afreyvWR5bhlmjog9S/PKmvTGuYtcpZlqPscZoc
sH7pzhJemZvajxAeKbLexv7RXASMML1FV+lld2Vr9MfZKkaU8hAfanhyBzSvp/uH
QD6h6RYAengKVDPpcNhHIVt5nFwttVV54jN7BO9+ev+lmW0ABe6NnHl1HwDScwox
avgNY10qe8X89Tea4ih3tcIBVUn94q0qEpZVqPHtYR2usbKK1DzcdmAF/yWPbb47
pM/mGybmynsLvQszxlNu1YzZSJ1TCvNR0Dmbi0Jt24iKtJBXKh4EfcJflbOuFTsp
XvOHIyLjzolmiajMdlejI8J0DAai6Hp2gHziruVSqSj8QY8S8LsRt7470CKzJvMg
2HEJrNDgpVJMf/pPHcEiCujKXskVD8jziz15L+AcnCdKHrxJAMfVxm2rCfyB5SHQ
APlB83HyjeQnF5ct+i3aknTFIPOw93j835BLxWfLTzxysWx5U8UZvtmEFOPeq2qH
9aEBi3v9oMWzmzAJPtSTcnndtsHzS9KfNo7c0rX02I/E9eyuEOAltQZPK8IAdUsx
hNC9cZ08/Q6DDZEY0IDA0fCqyRRSH/5AlIdBEDjv6tpcbKMKhzmtvy86sd5a2EiC
aefhBA8USREi2jfnqov/kuSC/ETItb0DUfYX/jSJHxJs3K512T4cUyZp1xE9pJJG
sx21/nqiZod8yJVEPyGfJmJcBsspvBJFnfTkmPT9m0r50OlQ91xhz1kJTds3YAi1
bldlAYbWcXYRLNpAV2UoyIM5527146+LZaL8u/WinMdcWgRTp70REjR2kkd+voHO
0rfqcMvAHglLgoi//CsvzBvCj4fQQpTQFzsJ0BjdnS30zWlfBo76fVaChDYP9IDb
EHpJUbhLDwQvLD2MxOcZ8mDScxh2J5bx+g43LHtegS5ovUN4qrl/XIAL23lgCf1P
5Dy2Cdw35RE8RN6AJLnK0f8QF1OK0C7JwMwubYhtZUQ2+CyLDbTAxshU9VbZZWQG
7XhOcdyIrAqG5352pV1J8qlxxQbl/Mo2z06ib8gG+DdJdynn++mtbV8eQvi5MsdA
3bbsfZyZYN2/3D2f2JZNWOvxh57cSvdp2Saa3hSiufLv9qQ3v6Y0APFTHWUHQbr/
dLOmjx76Ofh+QL5hkzJISYT9wuopzNkc8wDp1QyOuMxGTY4dRNlQmSq5G7bDJX+p
1XTk2Pk18XSJHEuarpdZMz/khzGRCqR3bJRyohOYlyPQkXA0whvXZFFb+Yedn57W
okPwxm6IuIgHUz3jmRk3YoFvPZs2Y4A2zVzlhsc9j5fWOzzgb3i1Lfluu8neAI5s
y67VjlcY313SmDjKREJ/hqnqRZNZ1oJxYwfk6s2Tob/U4KVsNZE6naovVJWsDvgK
lAq64pU/FmxwboBUL1aR9B1xjtuoABxxAtHtF8dhl5B17LfokNA9uHQ33MXwNevY
VYl3qvRyUleTBNOUvn/kGWrGSQmzpELPfmwQwzzqCLriRB/sImAnq8OETjH+wT3U
9AXSoZh+l1vJy6ydnBP7o5dhKs1w/icWKSsYyvKxEAN73PViYx4vyBVIMmogQcQ4
P9OR6Ucdcd9rHY7/aS3QyThiNNJL77GN0M2/0V429B4KgtsnQ5/+cAaMKHBRonNm
CZxQGogakdCoM68giu8nT0CAvf0xrUkxq9W/NnL5J82awuGUzGPT3hJNzKqOBUl5
4i+7NjvSQyPw63TqObtCcfSQJ+wemlqRZ8n3iz3Im9xW20VozvyFIO0TKWsxjgSX
Q3FKc8ZqPXVLzXjrEWVU9pDuoRH0nahdsK4U6sU4KSopkjPKZzZZiJgXiT1lDcYB
W7ylvd44uBfyQu9ZDMygOWRZrO2sLc7M9+JDM0YBmnpuP5vRE3pkAEbuDYFwsC6V
86f2itMrnPKgAU9/tigST55GZx46IbOQcALXQIYhgwFMLhWtgc3rDEZWK2l0w5yY
spsNoEX4irTUt0f1xItLhJcrkPkNoH7peAihrc9KxXwGsdleLP20L5+o6dtkM+o0
HWLHIFkM/tXbWVhT3vTxKJln610MAGU3FLQpBd1pj2Knwqo7mKv79V8qmjjQMUVU
BVD7C67dFlMqtemU4V4xjn94SYWtF2eGXk09JJO3mhmbptcDRi1kIKjAgmXFYS8q
MtUaTF4eQhJMH64zK9oYqxyiSf/4EsYFcewcrybR9DNRo+BIylirmR6dVBxSuJTE
a04hKc6mkbVMEPZbb36Z/JPxXXNzk1e7f53HzQdj/TurfDXtgElxIWrJIipCF/jL
mAlgBO58CP6euZFzYykYAOGGSZVdKYzjFGnd+etNf74o4J8bKRMixPqgVG4uEXN5
txMx1bjuJz5r0dkc2wN0EPCnBsbDW0BxGFq5EP7yLkl6HEEzvZUDLfytVKOwx9OF
szIN/GfPpW4TcRBjo2MeJq8wPMKg24wL4ZUv8jAQOB3PDgHM5j6gQk/KFTfzIvcj
H38s4fSshSHEK85ZH3wzgOrUqWRGxlqRAsAAbDwZ+m6QbB0LS8IB8vpETPIkG2EH
rVITsrBhkL0yZD+SbIEDwZ1EcLLvoUK+4Rql+ef18yxJ2o5wWaVLSZB55+7NDe0U
FrU6jiy87AdmuS4owUqwbBwI5MZermgT5vGG/ulvi+7BsBLOBPJqKIqL4FN1vaDB
wPzXB5DILiw7mJc+KxqPwuVLcIWxlm1rYHJCvesOFk6HrcUHJhv8slk40nYQIz0K
pMD10EMzVYFtwvamDINA6BJj+HZYB7GwAyP6QJCeVS0bIrFAA+N7h2Ti2iTcxklK
h9a+52nYkB+3ffUkqcl8lI83iY7hvJ9lx+gFsacVw7i7DQPzQqU2mkTuKm7fT9mE
c6RbYsVPUUUUKZYbPR8fhW/6+0SN5HKG39sDIc28G8Pi9b0tPFtez6UgPm9FQ0mD
RiQCZkxrG3qanwIftsgCc1UWJV+AZqyL1uHPIaqvu3j0UpO/IK3GZl1nAuWHlsqd
0+YP3kQSHtGNTd1sl5tJB3tNLQBHx2Lf3cRH2WVDMf2zgwhrAAmCuBebXZT+Yx/Y
6YYDZaepb4OOs+yjiYn2MKT5FErHt4RGBd6RJmcqrPFBQtX07wOiO5VVJPhnd9Ll
sR1tayrY2JgpP/KM8fEonvh/6bVoxC6fXQVIpOL+/6fGE08j8iXf4jbJIwPLE0uT
3icFV7dM1/H1UApGeYfmuAVte8q5JBamogM4Kvg1aHbGI/X4ABVLMH4RJjzcqgLX
NRrldRb2N2GR2uiSW2m0pUQ4rTTAuTNca6Y9vM8IWhCU0YBVyJSqXASivipfKEyX
igdaaOh7CU4Cha0TAZe2+E6nZa6ScM7JIvt2RF7vMrL3CEyG4fdlcYLWydSeivMn
ZW9QWwS9IwQwbTCskx57cerdVAJRDWDjy5C2PKn6bv0NsQzObo17yLlTxGMzn5Lz
HVEOiDooZF7PT2a4gbcgACbu/KmghP+Y98fn2b2MnxQirbOk0ow4Qz7XO+DrbIF2
GvhmRwCV2sf4p+Dhsm+o14xwbL7Xo9pEQ0LXJfClwT2v3PbtcqRo1n9EUXKj9C95
/I9Ly7LBhHfVsBkkdASjCTgAEawdjmzx9iQkxZdCYI6HndBHGdt0oO5CHPQV5mxV
nVP2lbV9C3j1+5JDvbJ2b6K2RDo21HKd1ZXSNbMtG2LJ+iSg0tlh9gU0rvnujbKc
XSq3+c6sEJZ7iSfIqxzm/JjVG1BtYaT8kzu7a+zReWg7I8za/OGCCL0TyQdnNXYd
Avy0LXnekvvaDAwEJn6HIj7dfs3KLYC1q3lavtYAR6hg/1B6hi0KTOTrc7DgWnBP
SO4A2F64HULAOsKm8/9YKTZPTGFcz6oeP+x6pblFyJeBGOeuJeL+7uA46cDs0DXL
Fafg4xrAcQY/JZBsJhon0aQ/UxHggzl/dk9jOgZL2coMYrqfQuGuu9e5JfXl4f9I
PuMW4VZrYTjm3xnozJ9AxNxhpVgvsIPrQ29lvg3K6lJmn7rzPLJwXtb0G5q/pG4T
yH89jN0w8EFpRCWpJs/5kOeZ6d+BfDNp88EpxMaAsSdHBYX7/P+5KPHjyfPFjiuB
rdzuCWdfxXevxxTgDazPfzXw0aqcpsvZl04dXtm9JkQygt0lDdzW/+qMAxrdBFkg
HgYFitV4wA12Aq3ErTMhNbqSbdBkOb1R/LhmId1XQzbWazLQKMW3OhDMsZXsmG4P
BkPho1ZB7XkxsbQ77fTBuTiqlAHsmHtNVatGRUCgHepV9U68bJDKIokEcNPbSFhp
FZz+RfeflvGeUmd7arpF9DqgEJ0puQCqe6pqMkjUuwQzSNsKgjF/CNAwq3SCk4FA
4jkDllIvhzoqXbXeIauKkvO8LlD/NFmhAHbLP0RhXHu+ZIdOuykt8s9kR/YRwfYi
oz3uplA/D65l0GZZj1658YesttnraBr9b4b3KE7G58RxLfvXRMfzA2l36hFpZarK
X/ARJFErx+6VUs/kkSVi22UeTQXURR1QE4V9yuel6nQJBgKNP2B+1nNUBd80KbV0
/NkchFweuRf2uo7a30bNhdoqtcoYM3TXetmLS7Ge/k4eGiKx9O9Q/GHeIH2BokeZ
Nv3lcwoWbo7lTxzEpUceRoxVlIP1aIhBHvic0IG1A+qgFt/g/MUk8FMVWXKCNuwk
Y/xmAk8NIYa0BCC2m5qSC4WoJSfVmRzW78We5mtQp4buIRYdHRprOIa8w9KnYopm
Xm6LfJ8uuIQmGoqYAwvv/gcSmlDBj7XRZ5YfbJaAJK/vmcxsZ+ATAMIiPSGsgJ6n
0DYGImQtkq+N01mbeWmEUYaY5U+Xa3KOUB3i/0OpVlrLygP4b6X+JTKhNhlKbKs1
d8vBvfNyN1n2YDCe+tVr5bMKr3NDEFDp07g+WBTKEWFMutwlvSwzLYdXRQ2PSpLr
e7OwV+vMZgb+BfuK7n9H/+/wYsq6vHmrsNCrx1ZuL8d7lLcoXQKkK3O4JKi1acsp
1fIose++iY5vVTfzuUoU2sBkqHtWVndqGdnlhM8Qi0lChWw1R/64YZXx/WFMsL7V
T5iP2v1Vwtw2NOhQwGcVmlsVqL5+90tEmENB3ipV7b0jTs8a611nbRvS2VfGvnrZ
yVMWc97IDt9qncPjKpqaaWcBJlu0DJqSsJO9lCjSLmtgfrBPlxhGdS8+9xBsxSzg
N3kM8wTAo02gNGLkLdjF1YVFG/cGFvVrMeWG0pLm1IF0lZqp83gbglucIq1/iuw6
825R5T27xmdMoOqtWVSMSrPSR9s7znlMmJBR/osm/NM+8brcw3xOqs8V9uVgrmDP
pvirvJGlI+VeLiJf32It1g27bUP5hXfZEJB1sZQK3V8vpKfhhWsCqsNlK0LPpW0P
Kv1gvV4C4l0g1N+f5YNBMJx7MA77XHD4Y9l2lJJBpR9uaa681b8Esfx8VFQt03t8
yo5KgsFnZZUfZHziwMX/Wo32VmPbIfDft+/bgBbzDifh5CL7Z/I03UI4gVG9dJRd
hPXSWNYPcGAlHcEaZfEXi31MmvowCHjm2cL374PzcUnh3V/7+bGxPLwyginm1Wy8
H56cDaBH0R9HZYkxFmXElNjMdcVzXXWlK5ucvA36Th2FH2mejhy2jgcpeZS3bcH7
Bj7Z0Zn/Q8MZUKn8r3grIaI86IsUcrEYXXBH5nemvavAPd9gzdFZQvhwuX0IYQCc
RKfM6tjJndRXCKaZGi99VsbWtY7w/DTbENUKJRxj8FrI988gOYg8D9MjUjHvMyEo
FM1RBN+N2w8rtpERMse5X5wOQ+DRIvwROUBF6YodxZ2AWb4KUiUJZK+nTKMJmv2r
DRkA+9SR6+hM3HErGedftLbyyyQfMGMx9AJX7ToJ6xss33aYck2pfxavGekPP0GY
4e15sQAn8Mn4gqXkBDgcu1mCCZnlCrSYkRJSwflWeohwGO3IPG0/0Yv2AjuZiVM9
Lagf2h078t4/qh+CdWZ6zjceSxZUJyxoWRQKNS84/Yci+FVCQhrOAHCpm3bPbGgB
Sm3Rs5r3ICGyPhqN8artAnr8BHFUyWRSypXFZWgA56dPCYEmHSPe5W3ipzSQdelC
bHNhyWy3ouh5/5k8K/B6zsPZUziNTodmC03M11yUKbxf4uliPzHESUio1tH3/sBV
32KMQ9xuKznA7RmJIBwgxr3VlB6zkVDn8hWqZHIICgawHwsL9dhAQYaPXtdtY3fP
4jt2BFMYIG6TAXdfKKkLCgiv7rUOV1z2YL0lowOCIuDZ0u/WUszNzdX6GSZK2i5n
pIQZ6rUTY8QxOJcaWswOEWV7C2pUGqhJZXJZOdzLdrXmIheDZoisOd0k8cTvSLYX
TzTIPYVP2tPSxNyGJ387PkfNxusebcrHCGBLgczuGGEqhKyTaHdS8nBb2h7kOI/Z
cjvBTydCC7lw5T/piKQJEKKtpVQ3/sKlRM8RCO2HWs55lGmVbbIzcxLTRS5NeLy0
5/OUVQankgrHeHOyLIIbdjALm9Lz75ustFHwUCzWFs6hDoCcF4AhRiML/8snKbOv
7NXw/2eQ35yIQIfWWLvOLc3lvs2wClZGl3wRwp0S2YOZ4ZQZxkIWuYr9p1HML7X9
fkRCl2v39JizyNy1N65xqJPBL4gweBCirIRI14UF1MrOdwKmvi0yU3dkaPhOa6zd
6lbTflIH/CLQ71RMs5HMyCwiZpS4sKUZ3Ky1S3ObnOgEvL8gGKN78EZxN6wzRGCL
3qry+R3mg/GwhHLfHIj+W0YBImfPCICKRcK0HtkibV6RkpWFeIFMxn4PMyLHAou1
eyB3lMsLuovGVcwU3YwEzmeL4ApItcBoTgsErJJBMQoxhnZSPrVnAhSROfSG+A95
5BAAXSfvhal+vjcFpuLCdiKv0xFQndtxOUusprRZL6J6AwY4J4J2mp5m5/Q0V4zx
t7Ufk0H2Up0tzuMsczseMzucrZ1if24OGVPQRY5mPeBqrx3Q1P/CuDCUeYHgDCTQ
vy0KwJaOqEfDiT6scG0hM78Bfeu0VIS8rTIlIoB+r30eXdbisnzRlbYQjbkRd5+G
Y641kAkzNlPpVlPzONwaBi9QM+Y+baSARYFJl4eHq7jEDxYe1r8FATia4mKQs1S6
m5v3T88oW3KMasV6bbnJsdsZCG+2/IDUdO8JVWKG+gpCMUi1JEwIj55/NodNvwQL
rQDVidSU0TV5yhPMNwVX1YkywcVSVx1m4qCAV35o2jrXy16juefoAmBYsQ6skPGv
AAhC39wdKcPEd68yvoMBm12O/IXoDNwczm92lnRvyIOdUdnkpEW0ELknPfFqyExy
qI7vJMWhsLLVNfnBJMCvjO4kTCs/P0rnPLqE1b6t9QS8Djfuop0q4f3wtaYO1fb0
4mEbPezbXblQkW8yl557rP/BByee2G6jYLdqzOFkbHQiVLeHmqj0T+WRng7bD4S3
gkIkoj+izOGfu6vBT+VzZab1f4YUDLd4NT5qghc+VHrvkCPItFeNfdRpPelAjJfY
nasuR9wVlkyyYEthxmtM9NcgNrNjXbiaC48sfJEfUEcZyRtW1c4W69KogDn1gLKl
ZwIkk78XlkuOUBAdmn9Xsfvoko1VHi2+PQomaLvkrTGiOlyv0Nditd+lOLK0t1pV
nxLBfBr87Nlvrz/QRWysCJGGucKqtVDjiB++MYiEGtrNtwbdMT5oVpo5plYiYMdF
nYtioyo5CWmaQqW/9pabs2AvXdIjTO7ykaVetebDJasrJhyWD51HyEKkT/b7kMc9
XgJ4Fn0IVF5MMW0X39qf1rKBTUO3lU90G8EEcCH0pp1px30JAuBhkTpsFVjEYBK1
QxWnBayWrXb4hnvTqcFn3MTR6mmkKL/jGBiGlOOL41sc8nlTxjQeTprlv4kp+k4c
n3y8aKV5LXcnyZlx2uewcfJogpQ5Q2+3kl3MFpi/G2PK4MWdlR2d8Zgmz4MFWycm
zbDxUyS3vuxvZnO9wd9HxqZzTsp62bxMoiaYmN6fuPOzHK28qhqBGUx/N1t0YtJ+
pZZpbPBl4ToUGJGinLqFp4jpEN+1sKt1y2o5uc/VPjb10SeXJDrrJtvyPtLQwsNo
ZzO75jpZ2yIoWCAKuLUz3BDBX0JzBwG4HCqjxBSAGbX2m4JbHvFlvMHU7Uha6evO
QVop0+qEeITu6RlIGADEclCwA6c82tiW0x+Io8SUY9b/ralgCK7CdYd+5gizYlvb
2zKsrASFXUD0xRT1VV6ShMQNi7UOMTpJ9t+3lGknAqyVyHVMZgUFzjjlpqkCrR0e
44JFroAtgIWr98k/CozL/ylHRWWWXi/rY7IkfkrhBVzxque3NAvc7EERVd0tCYjw
5zoBs5SJkPazQYF+E3mBzWGzc27fJk+4Y3D1HveebxCkERpOm6jhnsalVLvDY7UW
l+G6Icx784THpxGtk/Kz/weCm23j2ZFqBCwPSW3nHABW3AG5SeJ4sIFRpTZ1JbFW
XqjZB1YtBVv6ogIFMw9SLqECu1pUm91WYuobsORvxhFFgMymPUG+Vjzh/Xq2C+Ai
dk03uKJKqc1Yx0sRTfSyUb7Ma5YvcbKM9Pc8v1V63DX9xEB45DyiTLEr0wfn9sxW
5HeN0xSkiCKy/QjtwE7RteZKY7hBuxAhBlRru17KGV3yfQ3IgJQDX6nexboV1iEO
WdCSGvOkY61yqZO9auOKcPUv4ScDcAFTDalJ62/i3/0ieqpTRd4QFlJPEQcsrAy3
dO9w6gwaAg/Q07a+u8SBZW75cGYK01ut4pHDJZBvQ/BPsuUWcdPU0FLvK83Pze10
GDvhspeZ3mUeZcSIYeClAtez/ufvrOzzWHm1ABigMQXw48R0emyTt2NFCBmFOxVI
kzzB422tzpX+o6Uhb3pLeg9hfoR4aYFd+rFuoAemcRbUfxNWlFwbdf2zp1w6Asgx
gbjyLdDc+BUiO+kg33dwa5voKYQuPhcpayZ18M4+pE9sq4gAYsP9GXVfc+3R2cXR
i4IMIc6eMfEox2URAtCEdJKRrKVUDHRB411M9Wki0OxcLoe5MblKyYlwI6eD5dKl
LxCQTwgjO07fdFKq6JVH8LMcwQtseNa6TDFpjaYrpF4WIlhZ+VQgXVc/cmOsJQvD
MJ85yFjBqYaUIQPC3Xyja0806RPHct1H1zKS3Mtmi/Vf4dQ7AX/bDH9dD55cievr
gtt1qr+nsD7ntsZ4tOYWrOdoqFgH46S5URbZK2AlSlpCrGKnykULv/iix+VZRcx/
amv05Rs/kWyq7m5pEDZ3DjRFm7fFeaUvBFRQ8r3AQdvh4HlwlsEVNQu0b3cT2nWw
aPYxtgqWOBST/ejB4fQ1dz3AwLQ7FVo5KoCD3WIIr2MOovuW16M4ei5i8v7/4hCi
TEUxmqyjIZBzaniYiixAcjQV0LVS/Ts8r25mh+jXrDuTsxSlLP0f3i0ih63vGIxH
Kofg8nvYJRgPLfOEroBktljGlQ3RFhwy1+tnWkmJ2gdJWGDgVwJMTXnaGiSQYSso
5cEP06rxWKTpT+BlepaHzo1VKncrr72t/ZlMqV6LCYKrKJm/JnhRTRuBAtNmhoIp
fC09v81ROccmOPjhExDRZoybSHq1Bk0vVIpO6NHZBs0oY0yhX/ASlqn5DSMLaN5k
LnwfHkvxLjbYcUI9D9Z2nZNRCPgA01LMs7+CcbogCQnyEZH2LNGenZ84yXFMAI0R
JrNgTpAynLD7IK/hy8naFoA6BsAblSXW0vdy9uxcpnCvuNPiRTYkJHx5W3PAJXY4
qFP0ggG9imRbFk79Ka4StHfHvY+u1WngmOx/Q6gZrKJJT6vrOkFsPV9Xbq5cwmfk
ihou6bv6tqwJ1GWAzOevQ1MsHAoLutxGydtjhtzvkLoq4eoQ3UZDLikivfx5nrIO
wW/4IzrSVmgb1j7uk2048T0lJOd42fa1SmDvjBgpKy/DFi6X0qe1FEaSCcngqsLB
upt4l+XUNaj/5N52+LRYXjuFRMPIkt7DCdV2KEjw4sOgh4ikDbZLNh1+XXb2MvjX
88NpuPwPqixz8nfvUZu2EYTHTtKVUx04vovK9pKMNxmwu5jL9kvmQP7E/D2eod8x
kYgg+Q3LHkW0SJap7E1UI8qgQZXWWN+402hvB7UoUah1VwNJ1yUQ8xv6TerXJ6Ro
U+cYDR48UIl6I37DXakoSFOkksLnCvSbBeAw26jyc2euCe7DF+SVh4LaAnl0yrDK
yvvgc8YeSNCO9ADQZTBJxYzJp355OVFppbucTuweSuVepJsnn8ExccUtAACJY8ys
rQ50LFLxR6aAG4h61nhAW7FupttUEj9ZUDPmLF6IrwbrPIvixOQz0YvVCqACoS2D
HzRmclMfSQEP5G80Lkx71NwUVmTWzimBEjF/o1tKtpnhrdLGBDCBtY95cx/48naA
VcFGw4DZKIFW9ysFEgFhI/05T4XkRHjBnNH5i6+eAXpxuOSrFYI26CvI/6QByb0A
UJe4oF7jhTPypwzQu9pMEMc1pnbhwwJicuehcB7mU3EZM/1Vrorub9m73Bu3nx7K
hfHh5kGHGAekmxS9MO+0BU0nON8syRsne5SuMYJW6QyT+g+eDLn58pyGkaqWnw2w
Wv7/fiMLOFMzEO7cFLK4GbOMW54WjcjdCQnPe6SPHfVCb448HRFzBLOzvSJlRptk
8aqQZzgHwJ5V8n8K8DY/qVPWvWW/erSnYfD+1M3D16aiWCsqyMUXOle5rZfHDcnb
ujVdBL426Ko2C0tAHS95qz98a9OY9dtJgL/eSFHuEHKYz6lqrJK8kgoxcxjO+swq
5xSEle3lO5W+oEz3wAle6t1Rvu3helEO5/e6Gk42/wXQVS60RtYFRFvrdYq9dlt0
VOG0qdukJSZRagoB8e0yTmn612Uv3Jmsi2PORca2D4hbzTE4XMqUmYvwkyxIKl/q
feFPbPXzOSv5gK1ki06SFYR68A5R/kcS2zw3lU5oh4xZfCX7ziAeFgtxNYUQlOeu
CNMwNJCL4LeOLFyC0r5ZJ4DgjXIwNw+SiwJHPEkHjGoCmg9LC2BSRoV95aIWUwkF
DilLQBxlnEBESEru8hMa882MjkgUKlVwgIAGZWWWwJl9t2lWHAMcJYFHSWB/1Atz
f2qgGcuE6uUypske/OgLuq01NXC1GMhP2dEYZDLsOoI/PDuV2MV6fZj/p8g7Uben
J0tnojkpYIXmnsI2qMRjFEed/HomUKjl90dArgJxGhAPlnN3IaryKNojDy9hPTSX
rjjnf+mCoyWtCmoFHhRdW6GwgcvsnAHvBa/axClccUAFUt4a5P49cplGywWPAXe8
2zhEug9yYmF6BCLQiwC/TlHemTgjDzEqLupjd1dgu5G051OQXAaMK4P/T+yMHt5A
5s+RURmlXpwxX+4v0IwwY1GB9ACwfWptSZv1vBFuKJpTvBWq77bzumnbFJARG+Yt
JJBlGe/Ed87lRH6DsN+NiDLwyQFfhmjBEM32erx+TQSBjUMtaccVRVJMEpanXgfu
c9c444LvMJ2Q8Xt9rPGM4DxAwcLRGXqP/N9pGdTOkNZU7FuBNiLl75G7f/0gvnRU
+c/g07UPg+kAWkTYZ6C/k+3h2jszuBHG60+FT+xvrTfEyL+NeWFnRoPCvisp3lXx
zq0/E5ovFx3q4kLDX7lTPo7u+F74Lpn8GuDFwszc9IOd3Swxer79iJCPbisnrRj8
j7vH23CWlC0L+NQUMhrNMgkDf05Z2f+rZurnkJEpyvkLNW3OfwS+1R0Psl5SzWFq
BJbrak0XPxFJMc9e6T8H4J6KYD7xDx6WhRaRvoeXHXq9tnXHkhyA7AWLwcjZN7HY
PfaeLIMlm8xp4ut6n9gK5hsBgx9DL3ZTR5jFP8itygrf0pUA6J0sPKu+YO5iCFZI
rWzqUEYRrhbQWnl3U3o7nv25K4CaCItFGft2RTT3sSk0qRlYwnZ6wDtuvhmbj/MG
hmvJ9wicpsaRZG9LKyqdy6O1du/2Eyir5HSNrpwEpgtRxKxIMEHmAZSGcBDaH+hH
bbfXuL3XlTzjwzkN0WmD5coOXYnLFaQ+MsQK8PMGjwfgiEKIa+UedfdKTWG+D32I
tAUV7NLxjLZ4q1L1VRNyqfgxxG6yEpxEwULZXOtUGysExTOlSpVWqCgi1TNfTG1A
OdmckFoeqQCHp6TGDosX9LgeVwyqtg3C68EU7Guey+Fvn4Hz70lgNMmM21jbTaCu
5yGvq0wVKlPNd0lQRo+jfXZmVMJcrFCYlw2LZ2RVE5GtJK47ORVKsxEggqk3+Sr2
JTL1jdxwOe7LcGCJCrQdgSiR4QC0IF7f0rTGNRLZfJCU7jmwJcF9CGJD+nYvbBRt
sbxKx0uV4azrxGROHn8k/Epf2155Px0xoFWerln35cd2g3vzo8JsK1ikRVzN0jf5
szk+3fOOTfBEFcC4mRd3ScNztkU0Q5kVUS2U8nNOD9xuqIbLRwxOtfYOxwDTGI6S
6LyatTZS631VIaeqY2PT72o1o5nq4zYwKF1R8Qn7iIWnngB+GoqZIr11H9AXh+9C
qBWoc+qDMqjgZMxWcU8V3v3NkHw6GNSuR55SfnMI0nHrsAtVY6x7uKWhzzDuajWk
1EOaRksV4x+ankBevVq/VdG96xR/Twgh9xpkNwpAzywwryuNKjnwsQ42LZ3QvptO
7gCuSzlDRI+080KXGfIIuakU+m4tMx0EL6fT1dZPxRxvQmoTdTE+QiIpW6wX+TmY
bfoQcVPnuthGdCDCI29gVO2+iaRU1cfwW8I8rLFfQ/WnGOCPSjzxWePPaMFbfBYW
T0TKAFbQSw9l/l9d7m8nz/bmqljBX7iaOxXBtPPWh3z2E4GuF7NweZnc3kZ207RR
OrH1Of9ikuWrYvYY9Wc0I2tlrgEQo5j8uFuxPlRIWIGkaaL5PpemiKZcpopVl1hW
o0DWR8t8AyEFtfyEXs4H8B2s2hVZFshyPpCP0t7WTXRbLHnPlOaX++j7KNQ201ic
MpGSreRuzAugWxu9MUx1k6AWX2PdaCxOS5ZZsF+E0j8p8g20hjC1oraUpRmrkEdB
nDerlaoaOCfSH6LLcS6h4NHE3uY+0aPylFQk3utKatsIY3H7WRb6VZ/akR+HlS8o
aPBZXYcRlFCULgA2mUHEOO97+ypB+W6E7xdx1gygpgHMNZ+LtuTyOqXYPwSPnzlR
WWYJsImNOl6NgBWLPEzS5UJTMZRYZEWA5tipt6dBlRhEVN/rt++51DgNSFrfEWnV
bEe2VJz9nTwCnKz/aHd1MuVrQJ0ZKkoenKNvIfLpDCxCMh1K3QPX03BtXvJrbTwo
P65cWE9wHekEQNs3SOScjuFMUMPwX2G1nSyvJu6m97rSlr9+Fau3faJpjPA2QFNv
7H7+ldxCQGcH1FLy9Y5yRuvQoont/XzicYLE8zOsb2DRorQPRZutXKNeAF4Tns6d
mb62gXibpBMdYHOcWdRVagLvsAGS5xIMCBFIkhy62CEIohVeLyxO8RuMj/56Ke2U
dh5p9neRXZteh0jUJoT+F0P2ntjWMSaDAuDP40dha21o5I6/yfkMOg53U/xCGAal
I8/nM5TgGA4TPiT3dKVafCwt2gGtA5d7I+JPKjE3BrWQ5zrrjZncbYLskVNm6gRz
aYUA0G/nb0nybuIaVDFrjebQSEnt2F9hPAGDfR4N/4WTfr1nvg77jfS3V0w1G9s5
+F2AMT41VJnT+7ZTvk3TUzs980jM41qTU208sICGG4iYtgxZSEAK9p3c7SmV8pBV
ccocQcQAs5hvQG+5deRNlLJQxPQ8Qwtnk2EkmMpyAv0MCv4LYZNZDjy+MyzzZNRN
uGbt4U66N5fDQEqxdS+wKoqau10d4XsDPY8IZg6AfqkO+GpeWY5mk5D7qtjGg5mG
XmKfJXZAve62HGRU0/53ithqIkcwXEwPRRQOXFg/Y3Mr8QJtymvLjlm4Iax4mwiy
Nor4iTL34Ecni2TIkREgJYHnhcuEm7W8uZ/fILDLrVhFPkoriPtVIqx+uLwkWDlW
RGG16uocE8D6AT4zWtbwi8wv8Y4xSCIc9ApANlNIIrXKM2hItl/cvBrfu7CRRP1P
r8O3SYnXOrey98e/pBJRb7F5k8DNT6PPVE0Av6G9tP/UKlVDoXSwZIAbgRKLY3KB
W17rpOtRJAa9lAaaiaugbSmffn3LluyZe53iicVB9GsN8HHSSGRK+W57Dp0Lpsmk
PXHuUM4F6MfQoysnnENwaxA8qGQW9gN3CURoBAWRs4q5phpFPkYuVpb8ueVJMPIS
1OUB4w8HHojZFbYNmuegg6ROLG+FzPWlOnA7+usRX7UMKoxCRsQbuw92hikfEhUn
x2R4ekCzfB9Rwu0e2VUPvqmfXy2mObq3bQcTZGAjSSrUwLyXBtui0dVeI2Iz7Ll0
qGXAFquNvlqtAuWTNi1SVzs3TBOkO3d37bLy5UMixraGhNzHNAKQu8zFht8dbUEg
3hfRlGUomJHkZSwC0GCw7A5Hvg9aqfHT0OSKWTiuPSqrYXAQ5KKoy9e3fS9vRvpR
dD8jrDex2chlwWQGetX2QC1hGbYcC5jo9RdqjR9rqUsjJ2QFCCpGnrwFkEAqTkfc
Qa0a2EtCEnk7tOKzJd3XYa58JjCIFTeQZZe8xntpDApmnG8+JzjTLAVYI69Zw2vL
3gaVnx+Q2ODqj6aPW2/b3t3wdWKX7v/973TTqbc89q1mmYh3u1Ux6Bir++PICLbZ
6iIH2IzTnmeAM40j3ikeqDesFdl8T4ZgqtFOe3JuJg9aaYSWvuYg8foUTeK7sCoL
ylTeUbg2Ykn+uXMlDpCPB4lenxPABUjyD1c/l28TqBbfKv3MibaN6l6LQQo3mtmc
fyLnInSF6keeo00Mqa4znJV5/0hUJytas5vFlIgfk220aHoeLC5pSdV48tadU+Y2
lITohAsv5WP1MkiW5xCgyAfPWHVC0OO3zh2bVnWenWpXuW+L55R0Z27FE22dvESq
l+sE9HTkwLxXggwbYSrqbbNu1OqQ/FruspJut/753mTZadrp9luJR3+3B88YLJZv
6NcwhzLA+mhDSG6Wx+HZQgn5Js3tjRAgRQY5/nXnQpb9pz3cGtfCp74gUja466iX
mtLFHdqUMHuki5icibDSSnaxRWjWkUE7thcSoVN1Pxbm+xYByUWshTOLHuElEfcO
l3ptw1XSiHyQQbIh5MIcLj7JdHSk7MrusSnEfUBlJnVdQBtIcfY95olV67pbcltP
ysDKuBEzpTD9LVgU2pwA9ljqwHc+M/4H8bHoRYRbQwT4bxXQsJ+OGS63Ml3R8MuI
ydNAUfjDn8455Obqx9waXXTXA+m4kKmtsfcGjSQWEQfYoF/yaGbrnkiev5C0JyZp
0qNJSL2wy0nlNmxfdxSkFHMvZDiEbTfHb9Huw9oVzQMOSFCSVWNvSvfLBA/LFz+V
TQC1dBFT6Zajs+d+EPGsPp1bwww/c3suQ7gRU12/4yNDWKUNQKr/a5+L2lcHXW/M
h4mh7lLZZTEoTBvaOwsBNb/kRGLOEy2f9duix9wHrTG6DduZGfj2fBEEuHSesITL
if2KXT7Zxp1QxgkOhPnPrbg2J5AP5Ab9Izf9vnxoezXOBmU2zaUXqNkInjiVLBrj
nbdczshvaQFaiEuM26/TsLPi4lyrLL2W1tRgRuXdP2cncIdtu11kTRZWkbt57fTD
WG4VRTh2NvVNevK2OBhAxIkY1lUrUcia58qhCfk+eE69uCm54Z7F6HZankRjK7nO
Pyi+TMy5ipTMZXJfauaYJhyQRodNOmiKSrhNgg5nrj1rBzQdTLmbhASA1Kot+xGP
oylA+8n9faN4RfpTl2UooIAN6MXFMSUWXW4usRYlqPEkn52BA1oA82KiX+WTF/rg
YIyBNWIbXiirwlEDXE7LEsSnHBWFYxYiJZyrF48TBqSpwHP5ZsBvNklz3TVF3Eqr
7MuWmcNH7oQsL/Tg+8WwvR+Mo9LyI1gGeDxZLoWEoBHf8i49ekTWiQKtEz3qRUTd
88QXnNY2ou4RbPGKrp6nBuXPlS5L3ZKkTnb5AHiGuapBEJXsybW3XQgQcEph2eHC
jFcqvqRQF3gdQy/RVuGBq1JuVX3Soo2h4qDHbz8pMXBmyJPczyKt/oqAExFC15Nz
kXZRLK0rZ6LAGeOLopt08Cbru2FI/779t0JW4/VWvexJ5SePABmlyeCjIus+KffK
fBjapgHRmRuxAm+aMHm3nShE9hR1Z6pCbpbvrWIZTTsAlNOF1ndAhDtwBBluD5xE
k5GzRtw8oQqfFakP+tSIsVzQyZvaOdH4/fTJPUcXJOLeHbuV2+zGGF8PYUik7OnO
wDNn8jmqDbiULFWQMYqXKXBwdpOVHjn8+q6BBG9yU+JcWl+o7FLxuRBqy7waB+3Q
huQHZFm+QzuBStEx94m6DUBssCclE9DoVQH2fyyzRJOPEpsdBCQsNW954evx9C9j
X00v6g6BvGCFrXuW2LWdRzbwzRofwVdtYeaViMMiYfthXQpUQn7lEG4gNb4MBd4V
Tr254S3cg46w+FnNZRrQ+ZyddOpOB/ioTj9a3J4vaGH9nhMkfz194j2/pnt9Xi36
nlXi6/UFW88VBb3K765Wy1DXpwY1ul9AWqY5KmHDvZUyiiWd1xWbfjjlYByyvf83
6ogUXefpCJshoEnTpEiCLMl0Ri0DIXKvqnZmPb3jqW78CuG0jkuGWjaRTg5g261F
KDjflI08tSbb2pi48NUV0m0yiirmoIj2luQLSmRXlFiEwORWAWyu3MWRcSI3Xl5b
+SPj6hNqaFnPYlBWAxUEB8qNoUj7WUNCo2RExz6PlvC8LYy4+qyRg1YTrQ9GKWG4
XAPwF/ARQS1Bkqt75HVj7MP28ZnNSHBSl+m6WbsEMfEeGx41KcKq94PH3bwlLJJG
K31GUZUttuVpzAL5A3d6fOEOCFmG7bEcSldMJE4Fqm/aizeQrpPGuA/xPZKPKJq+
4TyjokbOgEgk4wq59Y/vWYf0pt7bxhuqsL2dPjDWY4p9d7qwY+LFKsa1/UkdJHGE
UlofNxEmOOjnjEpMaUC2EfO4flHC5u8XmSrObO2CaKHMRqSoex39DDCTJpkm4owS
6SuVsYph3U5nsYNkbWsAK+6FHH2cOLoMmKhvzQ6SFFWLvJxApeJcB6ZxK6M9G9kC
PZyyPYv4g5tFQFh1HhQvfLleCenEiVeSHwTUZnY42ciDASOqr7JHr/OTDfLfiV8f
zgbHobgpGr09HTtxoriiV4La41tZIJpVEYAhVyJnQtnhOjUrs/EfNXYdQ9eHPF6Z
yTxO6LyEi6mtG0W2Syx4DB0EdWhxUZLIfQ0sFzdzA9IAvmjdahzG9m9rwi5heH+e
v8sOgMIcy10+5y98lJfUA/6SOrJCaIrxTdWT+teakMVh+oLZ/7vSTrMZd9KXdjXD
k63BGWhdtuei1KxcxacCFBwWFQbFapunwjAA0Tt1OOyi5a+q22XtjuDYdxLVUO6m
LMyiLt4WLm7zV6ghKRhfAHgseFmCMMg1eZk/dITDyPiuEmQmrESJxorH6NhODFNU
qfzJAjUhgjDfrinBbQDLoo22GdP07zmdSjEdpa7jmlulHyGrftpih9pIip7wpRQy
aH5UuXwHyktYpw4r+0rdNK2H/ELgqOwf9Ay1SeSWxDJC11yKIhpu0xg3qC2qcq+7
UJudonvtvoKRdWdnZzZKrAzbsgD/I65G2h2AGOS0bZwgoRGl7/Fqy1nqnllmvS7e
z6MZ5luu9mygZxsFXntfnYWsh7pYeGxIl427usctBpyphu4e2DrZ1gaGAxO1T7HX
rrGBq66pRUnKsNPNChFwF3KVX4k0h4LDJ0/7KDsgta9UCn4k/AXWfdf/ESP1MMVd
GE4Q+AmAW9sjRhrMA8gkY9eoPC9LshCgVwjdnQ/nC61H590jJQXSbPTO2sh855/U
m+TxLn1UHlOtlHriIbXac2H5QQZN6ZgAxZZ/ycUFxIyTJfAy6d3n/AwtQUXRVvBC
I22YIr8ZdbLfcM7yoOWZeAPrHi3GC4OwJCrlYaDbivT1m+0sivkxvJjzBH0YPzrX
vKPmeQmutDfS+T8k9u6JjPccb/gBg/Wrb5K3MLeDf5GYV6NCFv5XESYEUzPpyGOi
C/Z8CbCRuzD2cBhKCY0nhPmRy43sMrn8PJv+QfcoBS1n7ZkgCeoMS72C2c8We6TV
40t3Z9Cio0iLkbx1ghL40vGJk9MNj4aDR2EUAliC4My4u4snYP9XWOk8aCAgWLbp
bIYnicmltmBQy3ZU47FtIJrjs6y8KGI27nj7CrQmWLrnUmZ4eEY64f5Ung9oA8MH
wBJhXUSXN3Z/FVU36CACUF/1ClynwbuqygHHwbD1Zs9dKSjYsIwUS/0xJscG0c7i
eXfgXoVHb8c6mlGdnZ547Vs7LTcV+hzi4tLMZidLS4bBNoE/YKZ+wwyaXQoz9uUB
QnSR0zu1ZaBQ730OBNnuQb+Gpv04cAiswJ8Gj5p2sB0IhelwMWb49IywTCHgFttm
zSnjiOBj9UDlUJRkx7f/Iuhsbz0bkN9dijun9w9Ucl01qK6OWtSmKj1xPT8AJ8gi
dOCPzBe6DFrhqSBePUscn2SEgL5BpY8hAiVZkRr6HG+9mnTgYRNVSQqaKAFnD3zh
XcjtBqGtOcrcRpqA+fYILgRbSdMb1kBPmVIr8ft2q157mtLioW0wKWm36UiebjQA
B6pV4l+y2YFJjtJvWu4ZKmo70d5XiB7sUlGELzt+2WSZ4fKkhaPAI6GKW8S01EuO
UTL+2oUfWbgpel2ioeHLt3XeRsk0DciVvR7dCre39mMGaBcuwxTS4t7t6Kvipqo1
ug48XHwAdjCGLs2RiCo0zEa5WTl4hH3OmC8lWIjr3x8F8SRrFeVBZvJbfHlHVCni
z0Dx33dk0hOUGPID7sxlQLQPcLH7LQdikA7dd6zEnFXMSJT/fBlODmR3BD1JLO7R
Eni/AkrNc2icBr1l+SMlqgY/HhPrwu3gkn1/shUqbyU5QwJHp/pVqSNJWsu2IqUQ
xe3Qk9jQN5EpspDeeF0jSvB8aQdWQTDcix/Slx8Q+X1vdRHp8hJKBiXgj17G0dpv
z2dwh247ZHqXzhppVoC0T7bbc2hAg9wLJrqgmIq4wGrkTsyAOM0ie17A3ZAAmj+z
5hpRu5a//iLPpzNx1PnY7hTQ5q7xUVDOtRo1DMl8w/SP+2feVI0qMSD1psmWK4r5
/n5kJENOqFeX7H4iX+/WYsc8ifyLD//TuBZZe+i8bPgGa12R1DTWBEcP6EbVyTTx
KNj6lfeuKl3Pd5uwHDQiFAWhQqPTTw+XEk2e+LGq9NccRh0+UXLuJwrCwXsSUCOS
cTwh0XPrBDp5OMBnwRmDVmtomX24eDZatr8pmew4eecNgq6LnRAE6CB6kc3q9+S6
J2PPYU81gywnmF2HiZ1+r2YpIUF6SU315N8Ox7OXpwNeIqNhmeA8CWOMhOVlQvHC
RIijk/Kh2nd7CV9w4UxGZTYfFD4yEj/llGx0nVl32FaH+hYlU3HEJ1zR5K0yePcA
SQfJZuEU8J7DNokg+M3VhgWhrBb70EVa7WlVEF5Ous1ipx8bKNv1xwy+ymrrFbRF
sbvoVYn0+LQvUa5HIz9V0uwUuHGRw9dw/q+0QReIpixJ+HmLMA61T9rdOcfJpuw3
B4Ep5ZsgCd1Naxvx5LjrRwbMM1zj6JHOS3lYn9kP8hKaIu4BQsfN0KGVA3bO+t3v
yN1R89UCJlyfkn6/RkIHi4sxpzCFOfp3NocuvKbyPnxhWq4wLE6cwtppbw7AYAEh
PpybweVzuZAmj8kpaSL/2EiO1NVIT1IZ19AnMi1Le1lWAOXkH8UkEsPWLKZvaVoL
nDh54Igsp8ybrCcEKzjfxe+Yi4UG7Lm+etp1HDKnIoUu47iIETNF6ztvUQ1E+LC4
74NvxxjLugqjQg7gfU2e8FjwH7Z8TBdu66HQMvx4caDGXThglYeL0qp7sLw0ZkOu
Pk+FCwm2bW3iPssZvx0UPDik9FiofBLQ+Tw2venu/yVhrdlnKV7xnmnjJz+q6Yk+
waat2UCXKtTOeuNi5Cl0pEaeBlIj+5nsHMmWQ+UL/0+HzsRSJDr67+7JSZO8Hl+m
i0IoWIR4hmMTONORT8TjjiSNOu7slp26TpQPh4q9m0uEWnZrs4bvZoPZe5xTow+f
MNMT88GwuB0JH2rDr9RK3/d9G2RcftoluGbxDgQ+YANXyBHLa4aaPoqeIX1jepoF
+dWmAXTMixCCX7WTcTFDq6BVyHM4I5Hxkc/ETVBzcFlw92iv+EuzsP6wJuZOcJkM
C/5LBtLa8DFKrxVN4gIIqEB39IoI17gUWrzip7/PDc25Ieg4vD10au8JSVcaLvDT
GF8b5IykquBCLMFYr6GM4fgZ87iQMdBLFVZAwtsSlWDVB+YKXfmzicnd7AwqtS1e
b+HzroCci5jUDnUOgcYat17W+OQ99hArQpZG1k1sNgrhGFfbfTY9FpPi+UEBEpeg
3Zov1J3krbDlhFf2aPK6FCtm8l/yMvklze9HRu03qRodpuBrzOQVq92inoj8LQQH
cr2z/i/YT4wVOIsGmLpBH3nODl8XkbVQz2tQw8oKT+utqKx5uJMK9DARxoIA6hI6
7hOrhK4bYR17ZYGZ0YIBHCsD3cxk93Z8UWF1xF0xnBRSJQ9pDnQ2NjFAoU0KTjSn
x5wrcBnQRyZ3kbRPvbZCVOwzOWwFxmCYbOtkjcoFH5xeS013o+czA795kXmffQNn
PYypRpVaWtTe00U4VGg5yswjYZJ/N+1tnhlYTeTBgsLdepQziIip1EDFRm9qN4yP
rWq7fEmPkTpFveP78S0bJhLuxfw51GQsqIyi+Fpv6btea0VePiVGCz7kgr5YNcok
L5owGdLoLiN8uyZImevUHsyAiCdPnKYM2vwsYi9Ij+qoY0HcLUj5KQujr6UKAjKQ
y+qU8s8UlayH23s0DaDi5XN5ATjgF62cO1Pq8vv3WRjtDOw5zWwtqz//UiBGRnIT
mCThMJbtZy/iUkgyaFK+GdVtpc3mDf3UT5uPHdnHM2wb4l/0DoZuXQR4OlpJjk6P
jvdwMC0uFrTuJZbhZBUW/GxdVRM9EQ/03nqWWGINWGTdcZA8Anvp3NjspamKyWP8
v5+xrsmWlRqvJSo1SnBwHngxP3YNFVYu4+LkGvdxBFNsy1901pJZGbgYWbVtMKXI
7lDHvoTRiMKK4XDjED3toe90enovTZxe1sRAaHBzyXkq6VgyeeOVYNCXa+EY1QsL
eAGETTD0T7tL4M5/c7nsTLSgT8ucooC/waLi+0+J3pxLCuoed5Kx41btXPa+EYNK
c+KJFcluniU/QIu0sZnsXpUdUmw9xgcJVZJFq3BbjtJ8WGZO2Cdwh94DF7O9D73f
z27aZeiSXQU8/mmcmAOXhLTWbO9QIxo21gFrjEwbLhtKYznqAg5GMq+DyQnUuN0m
bcj9i25aMunPhcaag5p+t5D0RvI8p6vyL8tzsvzKR36V95O2XsR/eCfbqCvSx8Hd
dQWaJHtoiWV3C/xRUTLkYfbRj6nLZe4gQm3l9DeIstt+ZYUMF+n9Mqru1Syh2OBP
gxMtM9Ie/iCPm1TkhaGtE+rOsgLQr4ONlWF+/pxO1yc8gFWU7CqhbPHf3OuFwRni
Yj0oyxNK3vAt5EB7qWCQdi77Yp4VZ6DRumVahPAOuJnPTaHwczzVU/XVuqJ1JfVY
78O/jgZEEs+guO7iJiZw+pwLoyBhTIuv0WX7sLmGlxVBHtZ7MYZ/W80685r/N0hR
tNaO55wPdWuhRTJVjNv+PjFabQ+l3XIIo0vMI16wiQHBrqxZ+Pub/iCplF3CP+pc
W+T/tOVqFGqxasm1dJ3HqCUAcGgEBCrSpBTC07Kpak9ppMv8oHr9VSQKYTN1q/3d
WBMWaV39/o0YNl0ewXVOPFz+ssFkr7leHtYtBIeP7mP+UrnEmwN5gWKkmL3WPf6l
RAjCtvV/jYgb/ZGppqwiqRz6x/th4vN+5wYOXuBPw0EdDgjrrpttZqXVYiRJocls
sakDukDfltt6djPI76t0vQO1nwXWm+cNMwjZ3Bkk15aNDjo2fRTiZWr0Tq68h2Is
aASlaci9V/U3i4kHH54B9Q/rnYXRonXpxGDfhwkE866/mLZ4h0zOtwJ0nvNmKvpq
WSNnhoGnEwEwpQqgz30ldWKEcERBx0dDu2tORMmnIDeu4+Nsgl2OwOoffMAs11TK
h2ieUFMhEiHVxFvqF8DSDRTFtqGpjwQzxWh5TV4jR2Xpxy/WzUEBTOfKfFCAwWN0
hUVUhhJVUNW6CevAn3EPGMILym5a73oD7R3vbOBTbTJkVjqBcij4cKFe3StdC0Tn
bPM3zGSLozKqJ1fh6g+8EjQIqz6ucI+JbJn9G5cq3Pg2u5W+WvJqmW4BAkgcUxaH
hEAuX//W5jXY63N0pCJUrS7R0dRCkN8yZXrc4GsTe/qD82x1pEK+MN8l0NILmYzL
NfLIeV/2UjSfj8ZTFgRGG4cV/qBpbwA4oOMvx7CuQY9rgHMghAVnC9cWx2munwQ0
Nh1+MsC3hNL99yTd1z+/b4aHOIzy3G9UHCDfVWndKDjsUa0I1RWCxUTCCQ08/6uP
r6KEbn5LaFeT+MKfDewbpB8wJYnOm/xs11kMgJMoMJn0mhMbE7j/UGDOXdzCBT7U
wU29rN7HhS7dSNH3w5eYRFb36l9CGqzc6E9SS4K7qtvl2sR/Xdv1mSv/SCbnF64N
9V5lxBsALnlSLPV8bjFe3Q6cBM0L25NbZGKR4qnIe/aousrI47wir0t77Jw2S5Vf
AgQs4bPh9P9jYv07mjj8LRZjDtfC0FkqkJMvXux8f9bZRk7TBZSnpzQ1XQZW096I
13F3/gbIzkHw9eZ6h8/rmFlh6JitOUbkFIeniqXEzjPYfZcrrhEPJaRfDpFdVNBv
wL31n40xrvj5rA1tN+VyFqrPY0N/O0quOrYZ2fClJdXmIlbP6Phm6AtPkeoUAox9
f/5s9XfidNC+E5t9fnvG8//fJqyGhbYf62MYjX3PzoBtgwsh8V9wE/9YUpWiFN4y
ejK6DYJAl1QO7Ors5L65L/tnUFqwecFRCeVYQoudLAU65P36173g6QZB/21QMC9k
p6xS1t/8MEt5AJp/JRnEwe4FOr/SRlePa130RLC+Gqdo4c58UpK/nuGXB/SL5d92
/ue8nQzCFMaaQ7d0zjWlxhrCFVRW3aLiB7hYbDx2neF3xaNpeO/DhoVcVeZ0XJ6L
6TRukphjItNnrxbRxuqsDZmRklHDhOE4+esu5Df7D7J2K0pZ3GCJe+85yd4g5gom
Bm8QuRrvSuCO+2XHhK7AWKk/2KfFxMxB3oOMaI9MVOUybcLq9z8/OSEJK1LNRnu2
TiN0MOgZ6tYQ1nHOCntR/Kee694c326Y8W8kY58007Y48JbWAL4Bdzqq0J0Vi6Z/
IXKQEENbFo9kimj+6QIYSkO5DMO2NhZv+TJLlvoP1M5E86gH/HqBbWCXUEfUGW8B
8sB0Blrxy901zmdBnHuHTNl1ylB5zNjXXdmgIa6zYJIk+i1LkunghkEjQXj/m/13
exVlj70q10Tao42+Dnkq9Agn3FNAIDhzJC57szXdBsn/DjaShzJTJ7XJL5At7ywa
t9XVFJZIiZfP29DznbbkzCEIppWqn1X/zLo+mHvZwZ81+H1pvGh+ODS7ESizWOCs
Zg3kEe6SlafKXASfspcI2pbQrTF21N1d6eamNRm4e3HLJbpNAmOEzL8TqWYs0Bkw
mE6Ua1R/Srwc5Eru36nZfOVHfAO2qnhNYI2Ya9eDxLQKxj+ePZbG4E8O824R2RIb
V47lXxNEvh0oeLfxCfZMdymvVBD++LnIPIhUsMwxZenpSkuPr97x2MWRCWnZkqsX
9gklAKSYjdrManU41m6gPIL1hyFoohjpz7jh4+UPHp+MJ97NWiMGOVzDCGiN0rSJ
5Gpsq6KRiO571xY7dU0wMfT8k4QqXj2qPpCeELsP6N39q92jzktm1UpcInYalhX3
TJ2gW0R7Fhn170nr7t8MhZsr5smDKlHZcvtnyf6nCFQktUnwUyHl3SY8smWPgrA3
cwNuzLIF/F1qE24+43dzmkc3uj7PQna3tEb+FmZx7/H3dQDxT2X0aPcj11gowXFL
rhJ0b8e07EggxZRWzv6oXiEi9rTLgKuLRoaZO35VfQjMKcIL8doAx//0403cwJEE
OVEQ4vai01Lx1kPrlixDw/EFkRcSAHQ48XkvlKjB8eTm8cpNqiYru8UZrSo94cwH
yQjNaJexA7EvYwfEOD7EWZEfX9Y3Gi8C27xcYX8B2tpSOLT6l1R0ZMtM4jUKC5gc
DxQgRuObFz42an1p4l/zxY7HOQHbuE08fx77sofUCmq99q/VeXiBzkA+AfnzCuhX
n3Rik6AKry3YseHXT8s4oVrRsNw+Yug+3LEnDBXMNmnyif6vQ8xDJD9egc0lPL4v
pTUhQb7tyfUNo3kzgueA1Fwfxc7xQdYdTbF1wtGTRlIlD0GLnzojdEkR6hhOQzTk
Pi2UNPVIzqXIdpbl/5D0fWCMG5ydzLb4L/KO3aRF167MOFEvXcIzs3so0Jj1Ug31
jJwfvJRe+8aCzQKCIFt2XwmxOZ010X3GL6EqGFAv/gZZkc/y0Jw2dYCtIj0Pb3PA
2pUkmlMM7zRYUllF7vAJkT5g/NipzCqUabJIK+VkrsLwTYEL0EFVDIm9jvbPJxlF
taMqCi+ZTw5JrU48Dkf3vWgnj+UwKwCa5wFE3WbnzbBB3X//tvwVq80B3/mDI++/
TgwgHl2FRqE6Ta0juDfgye832PRcTX75FyXTPUAVa9wIbREUX0UrvDvEhs0xqBh7
XVLkSXDU1kF6lKxg/oU2eLDhchDe1ejVQjKulBcz+6nW8RP1sX2g+lD5NAezwt0S
5SNlj10p2mm+SoF25Kr5/KUu/+NdjoTIZrB2cwNLqNEQ02/m+q5kc27YRQPrCVaL
Ty2FomJiq9cl7169kY6HCZYcHokNfxt911QqJ+Haqt19rL+fPPwRHhXg3WeUtZOI
NfX0wqmsko1QUJk+qurxD2oFsXA0a2JDzIJITwLPzumJ5CKIWzeC09Vm4QW6JZsZ
O3iFpXvQgJ5+EtdpW/bC0es0PK4juSGn5D3P/pnqmfsr5gRqTL8o+sbu+/zeTFA2
YM0v62E/idnawlzpR07sE4ICr+hg+bn3Q6lmPLGqNHOmxtx7xYYJ7xEZTyGGH9sW
fn17CoTfzNnkaExgEVAXrkBlwPvUF7mrwgvgKrs3bdToli7/wcUwdbACzUE6V3CY
OsVEoMjNAIhX05N+egRObJWMF81ms1xf11Chmap/3ETg0QgWu07VOnmDLKR59BIe
4BRkqs3TCb4Q4KCXxzCGhOOmOq1LAI99e+xm6UzrLdXW3MfsDFS3txU1zdOqlv5y
qAoQ92PihOYI7RWbXa/mK0qBmFL8ilyDV2W7uWE+sEnTx9ta9Gf8E1vE6HUGz2QC
lIKJ1T1EUlckAMz7PPKGZTnyghHZj1U0nlSM9ZOXyB2yCsOR19r4GZBLhk6AE7kr
hEHjMFxaRMzZ8H6vlACLaVjhtavVoVWYIHxIIhQg3t4kxS6bciD2b/iQzFrhapYx
mjQrTBlmbt8O3yfFBQYMinlvpNQuh4EAIJcyMJlMFAXmLc1Eiz0Xt31SN47NZZu1
nDZN6j1J9MAln6SqaU3kBRV/RNdAscJXWZx1Gs8F+3ozZr2PiI4r2NVzc2keG6iY
rlg7ZiX8ugEFaPwYcvK16H5EWgdd0YUitjgsnKtCiEtiXdi7JWZs9kiL21Zr/jI6
hoTw6PNwhehkM+02HXRSNy6phydiBvWavCKD6nioFSRxliIstyCHsfLHR+o69fSu
p0ypPLPKoCyOD4FAvur/dl457Hr6V8X2nkeY3THv+OahEJY21rgg3o6stl6jlAj+
XV+D1rpEPfDzoIYCtUJU7WZYmzcIMEKHTPrVWEdLyKLJAx5UtbalkimcBEjl3mWC
vuDYuv9ZVDoVq/ABJKNESwjkIRia/pD3pZnIH7H4ytNo/eZc0CU84cH2ngnfIk3Q
72F2jgzFvKYJUzthfK7AGgzIDIzLHk0VIynU4v5gUEyvCQlalqup6bUwsLA/+I4X
AiH2yH3qtYvC+tbZT0PNTtzT0WBG71Uf6Vx5UTFAx0uQCIcjxMcUSf5etj51t+XG
ZNjDXJQseQVGrJhB383QGqoPrzqEDYTAw/q1qZRKOMNnewV2mvlLesh2gvnEVZm8
6vgwqf3MkuBZzh6f1ZlcpnbP8eUIQJ9T8LqYNghcK5FyWvJMh9qVqdv7Xgc6q5AT
WrFp2j7/lU8/TsYbuDFGZGXzTaod8UbskUrjmcCITFVYtept34gRYiBeYlSeIRch
HGQLEXfejVO2blJo5w1YdKjH0GxSbTq0ELUP3hAlHaYm2+Oo1XBwSfGtEeTy3O4+
nlIeZPPXOQPk5rXShvfIZK4ssuC+zugzXq4y8Z8Q1wgXg36gWzlfFXlhi53a8Zu0
IZkizuZ/F4oJ4QBFUwZVBZnQKQK1UnBBfwhbBGLjc9VdsuTZHOFYkDsrvkA1keqU
43X5vpSZ/gv4W/P6Ro8p6HxL+wFJgh8tSwPTJjdICia6gOO8HS8AaSgH7JHkUgrf
xBJ5GlyFary+AFJ+hG4rsp13tPSEav+ja3fIZ2bkLMoKZggTDR/9vRgStdA+qV8k
4mPaZflZunnc40T6fD+JhxrUq7zFcjtV4YC7DUkpCBDWu48qaeQ4wQJUjr4qVHQ2
4cJOSlyWyuPzQ/1MpF6I3MY5ZKzQcwh7UDuX+lkNkJTyMVmyhAukNuqzhFMLsxX+
7cYJmcRQVPku7x08PRADRyIfSPmhGLYjzoB318kkd2KGKkRvBgYb8PlaNy0utz70
45iauXhQ4dkZHnO+a1FOYksX3DbToX4vX/rOPfmM7Q7dkXZ9pbAo1A+i+1rjzFxK
cn2RP6L5w4PFuHeiFuFHCrXnA3SlLY4arj4obbcLqdH7UbLs4jKMc9owmozlX0SI
i2/CBbHSCkmkifXrmR5+hWDTkWAdhkZuaUaYblwQhV9niYi50Fl2KQcqBrwiRvIz
WbIP66+1JzvW0R5pLxG/5KXpttZAMVmSvkqV6KKnyFQpN0aU/Z4K4R1ZKGxfFLYx
3C0uEVrMN8YBP7oPrWz4ZlAmr3wWbRvsC2RQ0Lnf4KnNgiR0TkralwdQUAWJSAYA
LvMGrcOvWUH1+PBK0V8bLooHShv+kduki1EKF+hXFV9gZDCdXE1rSAxWcku08yUe
BtNSqmctEb037axmPQrEA4ZIaTHyDWEb3VaN73YravBxUZG12oNAOduKyqmZuxdk
hUoKGytCU0PJYkU0jcI6UsutqgvydEIdUvzlQlwa0osqD1Gjel//95sO7hUGufB5
NiPLWdzaW/Yih8yUkCVuntAdvgyi3OqZqGIyiSV0QNR4Tnsqv23j6zbRCtQi1iGb
1LjPNb3oFv71GxVZ99Wo7VUrhNTPuttvUyEUoRbQo5KVXADjOnBImDd/aVCZ0xfI
A7DjxY6U69+Xr4WxKMMkgp3ghY2StwzOdEFG9ykrFHqlYbgxidK22qAHGK2tlWjV
E3AA6AfrPg8NLB3EBa1j0n7dZLMYVFD50TTSQoDxg+RTztoQa3d+SpEsA0AHG/xh
aZOFCZPzPrUkDid9Y0Wlkin+lsH3R8lYvYf7CenGA/EOIu0ADxn692GZ0iKY4kh6
cUkpvtzaSLOe6TqBXzHqem5ASC7EUZpRTz+YfDgPaNJS4d+UxB3rVS8LAH0v71Tn
qFRA6ijsOh0hQx/qxEgUNlG7O1b6pCK0i/7XG7hEPCWNq5QL4pjxLm7cOSb5ip5c
8XGdq8weffZoSc7gXzxXZO3/afEX9gua0WqT9KH+AD/zm0fGuGEZllqmgYP0nGZR
C1uGsX9VlfltLcTagqWtFLNmQUqS7Oy8EV0rYdT/pkWe/vn2a4Ao2p1jSKzzyazb
RfnLtpaCFeNI35BA/wfnlLpOeV+7Q5IQtfsaM78B1R0kh7XpiqYD5t+mRMugCIJO
SewTQ2N9nYTYiInP1fKg0XPJM6SATL3/8GWDvxiS30sX2rdSrAm4wYybTmjjASWv
s1tV41Avza5XfAZMgiUTFrLBzs0m3FTTc6Z/orpcVAtdPTppIc4HA91f6LvFBKKm
U8/yo/50OlhNIMPRkk5KY8kPn8pkc8qaS1F50OFwpRcZMSvo2D37gSQfL3bI1Wud
IsAB2a5YToegyK38e8ebiVXzDWrP/kf2uEIPxoNRlM1q3nLtb9NSLtUwL6GOW08y
OR92CfR8lmmB2X9pHZs7AxJjC1FtxUgi6YHLkYi3Dh4yrSSyikendspq42U3bJMf
o3w/ErHQKIGYglf5p0klS2VihDZV94Ed+vi9XlTVtcLuxoTK/mkuJgf7Csy3/t81
34t5bckJABIXkLKTAGuiGUVHOKvI+WCIRVvEqGoz1ZxBXoZMoJlW5hsOgyQXvGdL
LSiUvGZUrQ7kT1HkSNcftbYSn/49ov6zxAV/1P+LXelfqUbReyJ6VzLYdoFhN/3i
joT6+PkkkvHM/sCJsHV65lYiruG9q7EAGf1I+ojZhP7clKHHbn0xfRJzbkNrVW/4
j8VBBbB6VS4WNxFnePBRNTnitJeQYXa0e29cCr+5eF1sf5hIGLWk270+EA5Tp5XT
NRBiXCkqttqBxflyxRa2ZzsSRwI4lHuAw1xyhAy3puGTiRXA55UMZDRIcitZe8El
YpCQXtlbqYaOM4DjnfNaqT6LWiYy4NAaOVarCsdyLgkn6J+XiLb5f6HCda0klHeE
7BoT/RXCev8ZF4ONDU670WhyESQIgBOTH749OFMR2hEx4jLqcBAIdKe2Bt8si8ME
08HudWL82S/Ax4C0fiz+66emnEQHoq5v4gqxFYo6+rRY8Lyi/fpE8bcbAfbfSzPa
hikYaxLFPB7uLvjZSp4ksyUWholCcDMA24l0XIp7prZolxJj9yWnllUOdJjutdmX
qx5MvvuAU4qXz2YpjRiKibmlEMJFhA4t2PwNYVuvZqypIJXLdQ57BYpma2dU/oZ+
WX5Lka9iTfs7KY/zhtXMz3K49gSr9xLtz3ss1KVSDBxmoMAWO220TwfG8ppU9177
PzyNacJJp0FuF/XUCYgkY6LGRIgzgA7uucJYZ1Pv9G2X0VAW+yoFcgmGAMTk+viM
+StI6hJRpXL2UOEDN4L0GGEhMVIc0baxDv7zrC7KekfCyuLGUUkn3cIM4ZiHbaAL
v/iD/CUttgg4EPWHf6xgR6FYpNwEToR1WTy8c1tLQidoTqTXoQOMgkXKFJKouRAO
gfCjPXkaOHR0Vriq4RWdj1UFlruGUadSN08FS9ZtO9DHTalVGpj2HVYwREQ3EepV
MFFVQO3+pBBxq1nNacYbEsPRu+oi69OB1gV98uN5+Nra/vxNhJ7S8/7ptDXEQJ7c
Hn5DgMQgVouhz0dDhH4a+DiYmkD7l8/IQQJBBYyT9I6GNqrmjPlFFN/iS01fHuwW
8G/1g4WILDXZcDfOyQeOMnbrcfDs3BDeECptpstyLO4yh+Ryz/QBbGxISeATLsq6
b0Ae8rhOpOs/JE1QngwpUaaArQr3quEHEVtx3S5x9vyLilLKCiIKGiDuKUttGqw4
aPxV0mTT/rj4vOb+4l42NfDqY7ATifVvq9NjqGemHoRHA7+QbedYBw9ZCv6s69q0
cGLqHvwZtsmMYgJfOLGb1nqScRVopFOifjVS5kkrYcezhQ/qA+oLqVQx69S2d1HI
pmlY94wobwBDcfMKoSIUyGVVDQAIcz/MaoC6az8Z20gNlkH5xnaXkty9ZWvEIt3d
BReeRD5+toJAFDcPVdJfJNFLDy4b4ukmA4U7TY4L05Ejpbds7mQuOqfDqV1N5r2s
Bab3wDYnmpojKfHX1xZcTL5hLrIHt8wxvv/WQEYksopDxopgVwJ8j9x1xMrdUczv
GP7q25R5DwAVRNBrKYr20ErQ5HcEG/BA+0Zr1neHEBqsjrZaqQ4XRA4eU+ARlIMx
a2/InEi8nUEXYcpRmSk5iB5HFI1r4xQhzH9T0h5tM80I1kKtPXDytK8y2gmRkx3Q
2yeVkfAXBc8/vTCyOjqP7uzqEhJf7nAFYPQMTF7LlpJHGCn27YmmvguhYrU4LNP/
0w0TOkMF8pcJpxCh/BfWsXvQfmEa5vx+gjoNxCF3rnGU2v/igKDxmaqsqsnBd4Hx
v14fWwNd2eSRWxyts7jKrGdX9okPDlWrQCNv7lnMVPOULGSSFjqjr0BIPaAFcSS+
bBtZhWhjAIkhGY5T6tnH5j0V2/nGdhPqu9/TmQ0RxgS1tHWEoJYOP+Dy/uXiD3RW
0NRAnVboYTGwUwvZjF1Epb4dzMoNKdvIUmAgfFNSMYsoGnFwpTq2eDi28tDYqR2P
Zdso4EiO3gpkER+OZjJFozfPFg+mXqN/CaVgRaHiS7eE7zcvgSYpGpGTZVrP1FCq
9LiRdMDxhPZ37DyQGjL5nVpcXQ40OyIhLCL5yRUXNkvBlSkJqc+IMGeLdIjmPZKr
NkZCk748OdePrbqv5sggqlOmhOfBb6DAtbz3xTdyeGUxYXx265iECzYKGR75qVZM
EoxBCJD1XS9WFk8BRz3D8Z1Qd9IVpuKSBKfYYGRRLs8OYyI7r0dmrki0DB1/xuqC
/PISzqrBeP+DWZfWoPofcEysjwnZFCob6277NgVkcZc73vLAhmj8FKmyDfsfU05k
sFYMrs+kn3VQePbMGTHmy/S9taCmOwLw6xTOTa1oH/IcJEyM1LyNko6tf+pBi6lH
ByW6u5J0mczHrssIA1kHyZwQWscJqpZ6PJJdzIfNmYfreatuM2Jxz9Vcu3ZT2ESJ
k6qz1nFGgBP8OMoJsZN1mtL/4pWr27XWN6HxYCUVUBdJP2I0YRdvwWSQKNnFtWSL
Heotu5zO7nvZzrlPiUQKur/1j7yhh1ohplOS2M9zZEnuVn2vdpv/iQKEKKpY4WRL
N/c+aHMydMHvhRiJwOG+TGkigHaBLku9bYqASTEDeL5pQge3yZ6VkSH5ze+RJ6J3
zO6MUXA9trwMraf1V7oBUdh7zSyAlyjI477pYzKlwqqXiF6g+Ty7zXUIKd2u1R6d
l1Ey+l9Bmvw4VeOPcZpRXebZ+9buevB7+CWMfjpI70dW+0QSqa2GjN6U7AH/i1PL
Yo2vd0gDXJHCnhAzMtNpRjg9NAvWF9VAgv2s1WUjVBTeW+DBDvfwl0F5S/ZJ/7Hd
BWEMZW2UdDMaEivIlNYTObh+X36lz2s9uZpu6xCXNG1zeUT4GLNIi1CX4gseyRYO
hGRTutG13bLN5JtlBsDxRt4qqhbw0b5zAYg0VcHopY20Id5k4rBtMNsRkpOEBR0l
AETS4XFX63NbveGrXJk95J3scb6dlbcFw52MravjFI1C92xq485ZUNdlFWXDE5Bh
npXT4tgB5hl5wpjTy9Oph+FfhM7wGMtpiLUrEEKBhnXt5E8vVUk89D1FRrKGpEwV
LxYdvMJpYpP5/g/owhSUs46l8GCiqFJTEEzLFjdFWGWWJ8/ltdeyLI6YmZUPvVAi
v49PttZJ7SEP751kkv2pDLs3ZlwYBPVYdup4O1S7mEsb2rz6eh88yX3ykw78Mjt5
/fqPOehgCuuQrTM+lbdZIrAMbhyDjg6tff3nFZrZ8tAuSIeDUvO4SyngUeca+hHv
LzP6SMj+QXxYHxZgnB2DEz6ORoq9y8eMNnABROOMRE+RYdH6PzofDPZLELz5VXeb
gdGcbd3MdkZObVAAYG3Iy+/t7osmVwyzkD8fEkPERw31WLAwmHeO6ZKlr8dY9opK
3Al/0VBanJhS7vaurcILqwf4gNr62WP3KrzbdNw+8pwJLQinTKH9+amcuDzrJ8QU
JVRFYDa04RBAzlT64SaCBg7V30YsmrvVqIfd9vdBMs/QsoknucFajHs9oMKFYbHP
BIMp20FgqAUqzP2F4mLrW4hGGxx7iFLev8lP0N6cPss/nZSaaFEHeMEEd2penrR4
bWRsR4SWiZ0CCkCTIgZkCuneLhuIXSkLbOsUFRXFMhOQbyT7nct5xtyUsYYDetTh
URqepuswSrNu7EY6PtpUTIq4Kz4R0vny9nBxTjdVkbLjEJWoyxcI8GPI4MSi4Zro
eQDs4dA4QURT/D8TzMmnT/HLJaialbhqUWZg2kBZNgXpppMVZX9xyuCnI5zvTdZo
060ipnQMKlRcQlGk/i7ZoZNy1Vfvf981jzAeC6c0L0YZJg3cOaYx/KEt3AVw60UM
no3f0l+gMNtvnYdr4hJsuYf28EXX3p2d+Z+O+aq8VUDbBOLRHLOn7emynYA5w+am
2e49PcIGCBKPeLy3F4PAhNUbQi10SZGRTDjR7VRMQkNvJZIBcft/2eS/DdwZjEkl
rnj73tqzznBUFm7kvS+v7iS2E+V9dpxhcKff4hU1nIL4w2g3uSJsHYWc75DPHw9L
vVobgepg+wrgnJ7U6gcJ971+q9ebMG6ZTqF5Hv+tYxAmMsenp1trOOf6v4J+CQ4s
LSL3WkZ3wuj17bgKVoRNtWquWpfXLXwY5tp6OidcYPoJlCnJBxVIPcZeXKLK+nXZ
GZHCCnbUo+0czld8fgMaXTqWtBLf/bGms9EKJ+qt/5PUXvvBumjIi4lZoO8oQ7+Y
0uBQab9bHIVDUhIY3Mi9C2P3OHjK1kGKSj5RGCbyLiXf3fGlEOtvU7PFdV002x7x
2Vtt7Y5Y0yrZ5ExIaocGUaALPNplCf65+WjtyaQWkGDbpGOZs5lbzuO5FqjI5EEI
sjuxGUjps5Qzln35pIBJJZFpxsmmI3P+bsTmql5RB6fX7LYHFYjsUL/NXP6IrsdY
NwRk4fzcnUTubi5iq05f1U/Z7Ak877j2CMnLLoN0hNCl91WS2+Bymz4ur25p4J6x
Uhsg+o1k2OCafQthC8mlZpTKlVvNxK+5wHpihNNe0NXtmOYVy1qXNLD3q59laB8Q
OXpdA90uydSBrJ36dffqkjQ5We36ncMPEKKIS7yPnX6J/nBngDM43u9oZ4wOFhp9
OT7P31OtHD1gSbuwvT6ub3mpfpux1mTd6Xy4a5hkZY1b0H4kyZCa352lvTOSuJF3
Ng/mGX6+9M9OBXFYIl2rGt/PHkLTNCLj/qG/PgaRA4924B77gyvBDkhKFBPppX5R
Pb01fM1ofzokfBxmtFgvBJacISXj5r2b03L5QrdAVmN7fjnnq2T3apSZvLsGlhJ4
Kw0euRnzAPRhDEjB6GdFbH/76AG6QzgZPKPR4ELaPG85cjaoyqjU4B4ZBmhfRx0H
aTaUSelZIGb+3+XVxbBvatWaEA2NoPe2xRS5XlGTBuqDeF+x/5/RziHBFFwFC0qA
GPk8VsNvoyKmw2KqG22ihUj/6OP9ZJD9HRSjOuj6YvYTWk2IUXpE71dplVrJvWmF
eceCISSTjCBybbRv0J4kd9YF7CEUWBJr9xtim58JHirPVeoiwIcSFX2RgRqNeF5k
s82dayk2/sc2Pl9uaXmyNaUpRMyia5iq2MMUcLOfGYx8os6ckOSu5lTqnYveWGmh
78ecy39S0zbQJGjsGtXa3E7iFxLPsSvFGvnq5/aQN4W6qOTpboPpIg3BfgfEio3G
tESJcSGTjY5BOjK/7W3TpZ7S2D+iqAZcYsY7mJVckeP47Lx+JlqKu4dMgW1xp3o0
RGE/F3YGi+Oo43ViCuDX3MSCu67hd962/CRdRTxI9fWqFEx9gbWavZRybXVsyrUY
RYmEMQXq2Y6hqzXNLS2caHSD+NEsJB6Psxe5szzw/dmNdH1ZD07fS/xyvlRdV3IQ
o7u5D2TEBdbGa+3wAVmeezvtDjhAidQqYzmUXyhLRVdXH41GQ2T/jBm4YqZ0ANgO
gP8ffSHCa6uP9khuC4TldifGwQHYAI0oHfMufNBsBhP06struJXP2Fo8yt9MQig3
+TXLDn2hpEYnDBNHjcDv7GY3oLW/I5Lz2GOTTzs8hEvX8k6pkRXUGUYyFL61qw+D
wgtNJkqUv/WFX8seIRuxlbn0GtUxvdKKTp7vVMnM8xIbPq25VBN0BSNVkN3HKgGZ
vUgWmefH4Kb4LJN8bb4X5YaAjBSmIAMLrp+W1oyGClYTN8hglOsEWR7SVHjr0Tts
K5Y4+QnoacYc2Kmx5VdTUu7cL1+LfuJayLk3m7CM5e3oPeyNm3LSKGqsEJxdCHLv
pDsrNYrs1cZkG6wdI8tMOptU+AYeMdOmmOwrUPEhqgYwDb9wqIg0SnC8v15Swu6Y
qN6bxN0m3CasmNSxIXwexbn9CseE94+/zaeR6XksxAq9rtamFKY0W/GvjzhtW9/b
kAza+dKKAgfDM3Voqts/21T/7TgkZeXtwjYAk94igUfYlAvEAzJLUK9Er6V/yZMN
b/eAp2FRs7gCaF0WMBAbI58BtRzvNd2uWpBZ5X83HVsEiotXJtO/PgTBeiMCQBJj
x4rYV42EHu3ZoDMY4D0shIBl91OlqiX/JJKP8+KeML5upNqf7BxPoypLxp8im6FC
GLgPSvM0H8yh9jA90848nKb6XsmLvzGPiIR7GMbIASgHgRsD9Jjz/iWX5uN/q2kX
ceuatTYHH13WGZO27AZA+XJGx0DmZO1dxodykQTFNiPflyjrdcUXSwlWcqRLUFhe
5FcD5NuFzUfqNAHAB6eS8PUq60IpcGO1ctVXvOrjL+LuyK2Xrx9jE/FoxhZTNLae
Hc32J1vzeaTX2goVjoPlHgQvReyS5mgVvEo/kbm68GJazNhGx4FuW96Ryhd+7q7d
DtRJ28cnp8LhjDqZk7F37YtGiJaHAUfmXBKFHcNBo/l4tMmVAeRZFf99/kTGuSlo
XcYwWbM6T0uIUq6Y0K221QgSWiex38FrzCZP5QH7rsbvjR20gvWxklYKBuDNUH+/
ZnDn3eM1i7G2TQ9e30oOESN4LrQARh6blzAfWB6vlaA1iSZ0mNqAjkGdwp6g4QoL
+8jfb62EWCX5KZ+v7ppXqU4+bOs/ciwILDwtY1nHYT9BoL9XpW+KLejySGo/VuGF
Nn595oGRZ6MTk/zFQqnpXLY2Y2Lrmt5OFbgDGIZmji1EfsrSsY4sFxB7I3f4boEe
/rjb54566T/ejLZUzo2bA7hK+948Sbrnms0iBw5F3N5FtW0KC6QYaIPmUY7izjtQ
Nmj0assC2+iM6263CcAvVIeNxYDR0qqeoySdpcc0d/LhiXWzmFwJDFXOjekGZWxt
oRj4z/oVTOpsY2eKniXpyujQZG1vWewEx45z4El6KLbFXcvyvUyEsc6u66Pb7NFQ
VydOSO6Rhypf9oeTVaZmK2uerjZOXqhGgpW/uX4o7ZwzpwsPhGQITLjwzselDNCN
J+taGzKivcbUB/BL8sGV+y/MJPOiyC5tWuW/6/n2dunTzZbbWEC9DKWzBD+uVxCk
C1cBqtW5zfS/Ug/RmNO+l+zpzpEndBJBESwYWT0rgUaZlQU2qyVefBupAIb+ARGe
vZNFqppWMpPcIqfe1D2PUo+h8GjH2FKyttUiuIc6ozKjHqP1fWaD9rZTiHTzh2Al
JlAZ7i+6Mj5R3YCxQZm58bh/XCTBbkagomZGS0l6geTILjT+5FVUr/qhXqg6tn+2
qECI3Jzw3rS4TSf6SbSejNn4VAA3lZVisXOUwNuBh7wAhlKsdADBG+q1rMV4fFhA
+N0inwav8k7gCMZZphFl2GzvI0CM92YQ2/JgjJu2KhTxP/uwco4X34yKivNz8Uau
69C41QWvm2F0p9zs4j5RZD+IxZwViiBsl5CIxaKlxkyPRE6DLZ3+4HaHmBvjugex
F0jLYbY7ZI9ymtZOPtQFk0jl3/EIZP7TBKolCOx/6/KEuGBKHPScafZH8RtV3sNQ
bBnUbPqmUXIPVI2n6+aSKbrDF931LpylPVqq65knhxrHl/qPsCAlmWMsFMCwJFXv
GvPN1DkmmdeiDg0JPlDw2jjAFwmlxrDwbmLybX+p4AAQA3s7WoKBSl37Zw248Eaf
MePxt9jU7AV9LU+vLDd+o/Oh08MZl2ABUEvqw3WtFTBEHilLlubxxInxkW/QrjHU
3OT+oX+RszgzvMB+7QIEPF3aNpraSxkqL8vu9i/7DMrB3XcP2ZbZ3fqFlL6U0WeQ
FgBBQSYZxD0O8wv0iI5PCQNjyCTQBFpcyIo6DnUuRJWkSV/E0utZfG9rdn/Ing5+
UUmVJ8d5mrgEeYzqZ5tbdpn5ZZkte0HwrO4/nzT41i5uU0oixu6mZrT+JgcqO0gI
BA2MUXkpFWPJbSgCUPZiyooyhYWiMP6RmXZBcF71so3hB+wSI55RVCIdXThjrULM
Z4fiInnjCmn7c+xtRlOKKfrFaOOLYgCvblTOaLqO4AG1ZGzEmIHB5wNkSmoHo3wz
cFUm3P8syqhEbwq6wGBcooJ1TQivePEIiNTncfAWR/uRxiDrUlE5up1HOSssZybC
Suq1x0W3oNlqto7Cnu8w3DJNlOyx1bNafS8kv1C00bs/ZeCH+OkqH/Po5htOYOr9
jiRV9B+59dJGL1uOuKpwT97la7iwcQd+vaQjRw60A0rKeSU3TYiZX4DwcZ7ZeEdd
Q6f/LFBG2maUE7ie/uELXYyYFOBYkpR+4wI2sjsxmfW2b0lA/hv6+XFytLf58548
XTEY6hwyW0rvsJhU59eEk+DknoRWsUM3bTJz55NGO13KltEcNHYN0U8PKJakgUUV
uKDyKx383hvWzfOxJfa/R6YvgYnJj18XqX7a6nk7iBsDpSyW1SQWTjuvJo7v9xa7
5dqaXkCkS0o0WZaFoV+CXCBG+ECEDs8qRyXotT5fAK99xJVxI9tbCcBXH5EG2Fmo
sk5Eu3wa4JB3gQNjZMwdMDzQOrLLQZ8Dx3Zh8nJRIn13k0zhS1HwzQsFqyP7L5v6
Dof5peBQHaOL3yhJwWp4ZMlZBOYhTUW/a7YTiMHlT7KugKlWSBr3LoWM4YHvKTdd
2K5iX51LU1J3N8q719V1mpbsqE4DoqL2SnDV/BOtIdxnBI66X2VtX9BkFQiMxIIK
gI3E2j/UV/TKRdq6C0NcULaqivt6cYcm++eOlNcYVBzopByZCyC+qa8K4OzLBiCR
OQr4JLG82fG+7B4hkKPYXIf9qa9RXS2wt2ay4afsbvS/SkReQUS1MhSGtFYwxg/F
4FRO+D3LMrYPUCS3vBpAwiefIfGq8Pvzg+U7B3N4uXmuLNW10JfXk+neEHHx+CE0
s/WEyBXEcdKah9pgOHNl2MbW15cnLuHIgJzazXeJ1yHwO4G4nZ0BDYjp3HwAb76D
5u9p4444p8WKEx71ezgdIrg7iEiZF+KqFKz+zOYF98o9b5IaGPsri+hNnnGAyrpw
tY+zyYEM9B6DQC6EZYJ2CJLWNhIoe7GWDto+bn4At1Puuqeo6ckNHK50ZdcFvrpR
B5z7cPfW++UgkWCDEBrVCjt42ZdOiYqGWHUDET1Xzf+mEzIPdIAj206UN7Abhotk
K9BL82hX35qhv/m/QfxIXuFYyFNVVbkrOLQm27jzS76H+SzBGtLkNQOI4tS5CQuu
/c12ujFWSWImMXy0tyQIxn7FkwgpKAZC5ssJJhJRrPsnl21woL5xlhdRszKQ7KYN
IH+OLUhmt/c5Lqkt/n9heiE3w4T77G++CEJiJY9oyEh8YF4Syu+wyOXKoU0JrLYw
h4ukPZ72GW2xb2ciXvoiyEIgdITMr4bb29u1zxWH5YAlGcpDSukiVbfqHWvQ2TAl
xnc1kdF1nE9qLfto99ZiZzf7DlRXT1oefVfe1gEFYi9Yb3tyZxNQP1QhxhGz37PB
2pTt+6FIf7pn3l/4v7e80TpJpxakh6/Ne8TmimzFK4sJLo6XI5OGCMdE7x1lL+cG
IFmFNbh1E8vTXZy/pLV3E0bQxOy1oXPrj30p0Nl8DVJPkOg5KxLybgekv8F4MGur
M+7ZMBUUzFpx7FqcDlDGJWn1IJ4J7y/EJ6kZrtcmVmHyJa8/XsRPFKXGi2UZFp3y
Rej9RbDYcQdgGkMMwbaU7I3J0+1ZzthKrMCPsddhAdgy6n1wLW9pT8r/lW3fx2QP
WDHgEZnpqN/avEM3iG+nPQa/cfoi+27qshqzvptyixRpXO+5ad2zELe+G7ZhIqFF
FDSXzpXjf/eYKA1GHAf+QUlU/Kq/8h6VsW41APzd7f7nB9xRb8T405bRJORpuaNV
3wuyPL7TLhVUKgtGQGSfEHs0v1zIwbD5bjPS8lkyrxr0f1ZIOE3jf7X8p/4/ErNB
iRrkgZFFPUt9mr6cX4jQ/W1JiVlHk0Rb7WYun5jS3QWMw0YphewcG7JMxq5XLSGe
/G4sIgwz9hRxG/IgRqGG8FZ3VMdY8czvZ0UeOopZWwYQmYd+6SrVX0r5MQiXnDZW
jIlUwB7LZExQy7BK2KjF7IUKh0cv/tbUywHoQlN9DFDlzKN96Kbvou/SvYaVoUMz
zq4zYbESxYpBI7EPHmyId3XusHyRs4EC47RQmtkA4jZpIVdwiqHQ+Egj+onrbPqH
cY9e8PvwvJZtxtMWUAFlKxYDPuZ0cAGgGWosirpvhBCcq9mbQHHeulRUti0GW8Pj
OSRiKylAxoOqgpKQLgu7JorcBLiXXnwCN3i16x4vAYVJKnzE5b120Lbkl0HC20E8
MG84NIwLteGjgYLm/EoqjjOMHoDl8b1vIONdf+kDZ/NNXQQa9Sc4Zrt2NEe6ERC/
c3SxbV3wZc1NWKpoH8QAnLHD7OuDCxw+1/YaJnLL2jKpP3nzEJve+ncK/gOgKnqX
y8FX33bh+JDTEm+erRaTRQ1B7dUbbs849h34zcmI7kHbdCGio/mNAfExb5Zr7rw3
mQ4rkvzk71wZ403vFu79iE/OTQro1ie2dWJAPD/BlPFM+hztCY/fikZrFluBqk0l
+2fxyJ9zQsr2hu8Yuad+GlDsBeEuI5IJBGMd7G0j3okByAvGg+tvX8vP4dkbcIV+
AT4bH5wodb/75tQosOy2B8LB86K3uNxeiOaMztpPMjJJLIgn/XWl1woScIiO52vz
xE93ZEebcF4LBOBnVJR8NQn7Kh3d4LruFV0dlegpQIakAGXexfu1D0m0zykwHynd
WlGa7tFq1gWF5qopv+Co2bPnOIr972XN4WTr2p4vOE1DsKzrsQrWxnOpbNct/OT/
tVeIPB3at5cHHf/A6yEtlkk6kiHQzPu3mQrt2u7L4+1YnsTNd0WZv928vaReO6TI
IDXvJdzmTZnUWxdUOwy7CWyDDJ4xOmle8eJUujUpV4NngKzxiodIHyhc+cLOHnre
qP4lIPPJx504o4TzaJ2tpeU0YRLLyeDfmIxr9v6+a3SniQUckOhjRXcFJr+zBQhe
WSHOJE4CqeGT4dWX8S1+tt+zBv1sh2J40OsqNQx48BeuyNzZtlr9ll3gFTQZArSH
OjFYPYwOoMu1ycYh1ypey8W1r4ZWOaeYnJA2ru+5bEnYDpIq8/0Zhudqz4ZqyTsV
itLsOAuhdYHiAuJfRCrNRdR7468dqEWhLIl5Va6HGEM9fp7atsb4xYxqyqYsK5A7
i9grx0w0vDMY1qh5E2sCH3l1eTgEbzjprAQogIWCphWQNW9C2WXol+bfG/odbBnb
g+YdgdSyslJKjfacngE3h1ZzaUxGf2Max7SysyxC19GsJt6d6K9egIU6IwbF2gvD
bD9hzUu1XU64vuqV7I4JX7BdjX8XxpOEE79g+L0UhJM6NqBOtG2X5SlT75wY+TXR
+i4wBlMjfFiHf8tjEEQQF8Af47LSf0Dst/JBaW9Qqy+CEa8HgzMw5njDjUGj9Xg0
Ajt2b9iFaw9rFGYI4v6G38wHVUb5VAsgY65fpRJUGLwmiumfspGBy9gpAzJgY19p
LNR38RThJ4N0NwCtaA+fFkXEvVW7aXrS1TaZJt6HQyi3HV/X41GgiqZo2/9tMWzU
3x7JDxooutt+x5TfVUS3x4Wa/q0criqi0ABOXEJfGR6MeWxHoQcvMPUlVm4LqbKV
Fcza6BTNcfGFrZbQiW6jkd3yU8IOuRxE9lUnKd1ACtsnbKaRR4I5xmRXiu0rlGC+
Rcp3vbpVL2rX+qtL6z1rubMIXBhRkIjpVPpZfA7nySmyKBZIv/b8unl6gbIFKJ79
HOumFPHp3AHw/Cgejs7byPEWlkIHyWDDKmxILLbBDxShAOb8Rv+fPAKPcW4x97vx
zzVEYOGXhU982CBNaATgS0zJ1WmxcNbOaqGa7pavYIzkaA+/sG7bkGUxscPspFih
2Z4AWD7IWHFO/UimvPvMGaQ6IY2kuACOsN/rfpYG1khO/A0XyVq6WV3aWglh0CJQ
mO8ZGqgc4+/DdzMo9mszRq85i/zMSSrCtpabmiujN2xxNFpqG0mNjlsBkpC0UXX1
owdzJI29m1Gj31qSSohpDFCxNBgIyKwklmxodFdAxheVNVgSSnv/BSSvG35gW6KR
BgTPo5EHszueVT9Us6bL0PgN6Jv/Me2EuKUKzJiTgIWFBHrveQCmRh8CWtbr/LTN
iVG2UT/OtAhKzepNQbM98SQYuFHAbRboO5Yrst6L0WaTUnKJn523t2KiXnhvdaZq
MWVc2ML/+rH33zNUB6ys3B+cQrlUeJEkvMKXjgYUvEQlsOJb8Jj647O9WiSIO7Wg
/VN8VPyH5C3ub0loSIOHHYBfoU0XoeFqvaFd+AmYcdxKcfdyZ0TD/nw25LZGZG2f
FxXaN8QNmdxCM7cDsFIAxeaQUWj9H7JReHb1tKM7sRynRxUSeKEEiIDHOadfgtdk
EL0CQ+BD9IJ1aRYVq2lmrMIXAAceMVPuB9KmTEyUzzh49UuzWN2Xs85SW1r7HLUv
nRycLcaCoHnlNDXtPbhff+t8xtGFAOiwSxkCR0FqMOtw00DtPH990G9IgN6HFT7X
NJ2AxETYR4uL8CVPCKxA/oz1ZIySfhcChUxZhw6ZgXC/7tFdKQBlrh3u0OfOYuuW
hsWiip1libNo3pzt/S/HdOYeRipTEkFv1JOksNbMRdJ9Z8si3HLktLsR/Bwf8ilh
24ewKYCpLOAJlVy6iZBj3v51kJj21IpUn77njho9IarLplK2mn5UUYhjbsipTh/O
0+3+4htG1rP9+2Pt3cIqJVhBlhwzrgex5miI86oq3X/gxt9dMTpQrNuPWoS6DvQ4
OaAf2Bhh1jxaPHmsIfjYCtoWj2XpZp3onDmQ6+T29JTtAi8QPjSvX3J3++X58lM3
H8B5bjlFdSWjZ8Fk0TZJF1v/N0BsIwBgiNzD06+6KILp9tqohnm7uMzAjhjV8dPk
9r788U+IMLBSzIFaXdCUuiyorRXNkDIeclKamIhJ98gp31jT9+/Q5mIChsm0ceWO
7jIUT6Iz6b0E2by8faIQgrqd+MsAVh+noVYYD9nfwPC1nRKC7xOXkZWq/9XxDA3q
uufnwpvNGzTMrYMO1b2bgH2ItOIu1+frXkRh/yHcDs/l9MIj5AAN4lNDhxX1BKrx
vq1W8B8v5dzOBkS+7jOu4HWigW0XJG9PP1wORrAb1p9MkwGdXk8lWFWO3vDz0//W
D47ulbOeifxIrko3eLcXDM6C/4XBkLEEBxhkIQvPfIcYEm/siAZBNnvTzKbDaD18
WWyMYwq/+UCW/aSNKum2M/dyH3pLhyPdPdhB9UZPSEje26vdgy5o+UsW92+n7SWr
CmSf7Xaevt7M6JCQAyRHl7oHx2PGctGt8u6V5/rEm06HGhaoYjYC5yAgYda6t24z
7rCwbTXjW7wF0n93x1t9zkBAunFDIgYXXRPhjrRsB6BpxrmQoLLzcrGOtAFIfLf6
qmLVRc+88HfKoeBaLlvV2oE861qY2uLnywur9+9Cf3HQ3YfB4NrRVYSkisbZf6z9
7ixvMXidkN/Zf/ADKzJVFHbcrERATEmDEIPzQEV1A4VRjDFvR/fYpBmqrtMzNVSL
KUHylEbvzgR372nHoJ02gjT8EvOXnwIUxn81nrCAlJ72LZeX0kkBe0WYutMscB5P
QnjIv+uVZV28OQYD1dg63xlTmIMjKaCIeHwiROqiEqKn68NdMTGKYLDEqK1aYuRR
u5mWEOTP+FSZgCTwLvBGW2aCvBpFsycNLjJae2y7g2vy4zW7iPlJgLj0RsrXrF/M
V7POAJO3t3MiyITv3QCGyZSG8fJvRz/QtZFEpev1IJmY1Bqm8EOo5S1taYBN35Co
niZX+OuSjjjqYiNO3Twvy853DMBm7YakCG/Xl8Vd8VpIrM5hlSTNmNGt3dPvoTwW
rWzV5o37/NmWqPR7JwrUBMNxrZLs76Li5NeThmDVqKlsUbrMLBmS/0tFw2Z8kYg0
/RTlLn1Gnsq5QegwqH2XplhPcUe7wajAvYagPVGeIAw9MxVm7VdUS4c9o3TUtzbs
9a4UD5gytrTTkawNj/PQTkq+GQ1Kvexp8cKIwVoSM30dc2UVV1a7HBc2LU/pkDGY
dZX3shdpfO5JijGJFLmm49VYHbdY7lKu36bBvj7+q+4roG29TCxUxz/evsGDmtib
Za3tyX2uHv5xIbN0aVgS8csSwfl8HuwC1a9RBnZ8A3a9x895i0hQBVYMIQx3Prs2
c+6PlEcFQdW2F6KV0RSWKy6LhVi5+JFOhyUdvrqkCjrWD7PnCChJQOBoDJzAce3+
7qPPMZFERclkoL1YsWHC/Hhpy+CURjO+UpMPm0h//aGIX5XomzfIVnHSG3T+2S2c
PGXIimwZioAElE6QjKKVahFV3yRWAPoDDE7nBrP7cWAQsUHBcmj3Uw4bzktPhEhU
Jk6US6v9PsR4xkbLSvMeX8nMVIMaFzRTbQBk4jcq1+8AG2Ko1zaKQwaFi8msDBKV
gw+HNlZfwSZkrDxaBBEXvl6ArbtZXpN1gWor5T2kZHAsG1JLvf+kV6b/T6TdzoDi
ytnCOPxSQip9QORftNBstTzPr/xYzLNRImB1O0oTvSZBqucLtvn6iQlSIZLjpQcF
9ezqVnto73FFcFpMsaihosp+oUKEbqmJLisXQDFKusSIwDFvDc9D2VzoBtqzYY4M
s0mMbe7dHebHHVSR1o1aSfCDkihfXx50WsEG24WTXbIUJU0Z7WzWcnPhNQMvsr/S
UPgMJeZSmHViNzlth7WqtX4A+Gwp7dJfl8mY4ndQnB3Jx14VTQfS4QuEFIyPSjX3
lFUnIGXwN91FKq63eo2XwM4L1MnjWKgLfx0mbtQYgnhe9eKi7lfnKy4ExTle6QXD
lJ2RGfP5gwftmHfJ6txBOSX0o8wWbHUja7PKaUP9daAqJA1/K+y8kzxaQ16UMtfs
GjSc7QqbjexNUHmqFwd1Vnnzg4sMzWwcTfM9/MfaSjrHSp2iV5yda0kJF5XUWCLZ
yRiImVmd8F/qvUOaYI4mYH9zlUhe2sguYAgtuNWoOjg2taZIPW431wUQnAteH+cj
pGRYKBQlrx4WyPnRoQlWbjAUf1I35q0b+fkajfEawQ6XPQ2rIq3Hx46zMCLDOpgi
PM2Mm4y75Yuuow22zqLofe/QEYxIiHPxIAcnfTuLC0N7UwzZ+7+75bEWjiKCIdgM
Z4IyUia5xgdbxpROHbpDg2SYNZIpmzbQeX8lRArPs4cXUWloFB+KiHSsis33jWPO
o53mY6wh5IOtAogwvbLbX9rZAh0DHOs0yVRLwf8z6w7XBDjLieRrfdKfcOd04gzF
qFQSRMLggULZLi2ADHhVAyuC9/PlbesVH2JLay5m5GEpQ/VIZRgbepciN1SbgAQt
I2A1s/AfeHG1Aojdw49CnmfWQt+vLQ9AaPQ361KK+IJvBGTDBjQq4gXLravCU/wN
XSLGpRs9EL1399u3Pl1N1lD4OyNJyQ1jojoBGf5/bYYapDqnSh4Zeftft2PowdVL
Hn6BnMoWP3P3JQnmDAjimtatSrlWNzPtaX8RqqCi94SsMW1LGUPIrXBSgW2bW9uc
TkisD3yn/xMT/T0Xi6CWxmuKAPAKL5plHfoZ2DqqFtoKRcOhMvY7UiBAkg5Xn2X9
VpOOs7GMLhqmDUAImto2gEV4xb3aY2Smc02A/GfPkQTjS/bII/d1/O4USO9I/tFr
qnEXdDNQDUzV3kW9Ul7AQ8NBFB0XRtsahkhU62Mwj9RquEs+CGejSB0XyZa4awUy
cABDWGyd8TN53VOcG0oQ97AT7S4T/g59zAAs0H0x4DaCZFImS8j8iVgR2rcK6PyT
hghV2RgbpQb9rpsNikduKV58DSrxVIlmnm9+/MeldbOHptQWgpUtp0Qxx4t7wxw1
MTTjyI5quNVLzmTEwPuHYkSwQqNf/xODL8Y017geLcANhasNwJ3dhi0X7ogXqn8S
CtWxHd8NcYjklDZdOPCwI3WtUBnL5QYvOEoBRxm+Pdcl/ntUvvlRSGLiiaSyYvTB
GuX+TvmhVDscQ4Zw/ses7zHIUbdKDaxmayQbWUCixhRXG9Aus2GpONPT6KyiY+Wv
8CEkSBdptwwhYsmeUKTNuHbt9zA9ZGnipTjj3R3ysYsYZDVLPvpj8mtIzi3y24LB
tsk/mShZSaMr9GyoMNGJJ6Ym2Jq7USNWhNBvf4hM2JjbIcBsp+Pq7DL7BNkLM78Q
7tOlzQ4VzIvgnKw2OeLk4C+afkOzqkgkzPs957ayoQDqyngQc5NI8Y6vn8ody2RQ
WNbEX+D9ne4qq1FUDAbn1kyzWqP6fbAK7JAc9T7h+InDUI078L8VAYtwxF3yaBrc
TexZVv8OGgioB9ltLgC4svbV2sfdEwxt2rlKTfYzvDytgWqqDDS0aQiE5bosSMKQ
aWm/iFIshus2j/pbFLe9Ryr+CGZfQ3bU/7SqmvxGFg8AajMyF1C+jJ7p/PB/LNU4
pubfzwgFL8zgpya0DtIXu2GutFMDOlqF2VmBom5YaVSvKt9g74L2h7XtwZyXGE5s
jXq5WGE0YYQ5840+JDoHUXGM+nYK/dKHBnb7qeiKiSv9U77p+DmTtK6ekrNhhHCt
06fX3d56G19j9tfBiawrGDOhYie4el7e7NW700Dg9ztTRGIIfutSSTcXdH49dFxl
lD28gGVZefLWKU4F9SeJRyNi12bE5iM5WlyoQFSFT4d7oLQ2CSfmTEvYRitvEhfw
oQBS1Q0tsiSfQh9yLB1xpZbzkwtkDpa6P36pqDZ4iZ1T8ijpuQqby4uJOOSzjloJ
SSsYOmrcDXKU8Hrapr7l/SDpKiqLSJ9urCrdxHHocG2nMZsIc0LR5U8djB/nhueO
ZmapHs59+dWsyjUC6rp8YZMP2U+caChKBW4hwrZoyRogFBf61RTL/6DJdXSguGA6
/hIvPz7tM+zchrizUmJpnc67BqLKBn0L1lhvDa/h6pnb7gltbsxvSZfdDvDzkgzE
bQFwghiBAyfCPqB8KEKzbDb4l7S+VuMLVZFyCmAx+YYh/9ues4WkKqctT9h0MAUx
5G3tHK0oT+UOHcOUTkgSKLGI0hbe/5dKTdK20PK36utDET0cUW93CIx5ZimlQCXH
Gw7m7azpk7It9nc/4bbI/ignF/z8RJ7m/bns0bWag/7igEVsZ7ldwugzMs1I+H9A
AWWbqAh+xZlYdTYyXwqUesfHjNCJ9fl+fLpNzQ0npCHW0AerkYDTzTAb2bdpBtOl
Tmqu8YM0BrLkRjYSHWpdDY7DGVqkLWASJ3fM+yFbXCIscIbVRCqRXFR+51Pnhzxr
m8G12GEftzy6RrrjLiQ5Jaep1vyq60bBEb5HC8g2xYZ2WUsZ6d53LTok2SE0lwa+
3K62NmRcvBJDRCepNW5zBs2l7FXRIsdKPphjC8JgmpYG1fUzuqflBXCDWCEL0n1B
5cbVjf6SjTSCwegn6kKjkC0HLJ4MT9bYV0gfR3gVssLElS0XyKs6/aNtpV9Pnwfm
oH1v+ba7+FKHPA4EehI134IXRfFvb+6bSH8jk6x7SUrnzPGbVjQvB2KZzly4idXA
i+GoYG3bGADRV5E2lAcyOoY3P1JM3yl6tzZaFIqEUH06KI2KfeHcbqfoEPnhzI4f
p+HpmWquLeD53YblEE8lyhhpD6iBrucdLP0uTuuE9XhOV4/w5EnEZXhm2foucesm
xopJF1Pc6NfFxifYwSTcg8leSZYTWZdiUmRKC35k3a3iVyqGgz4NnVY1+JJbRmGK
7XN9H5or8O08A3xW91n1PkIuYpRsvbz1KCU0VcdfiS92ogUagUfOPz2R6eYodVNN
LzJUmYx6syvBNyMrvPXU0/8Sr3BX5mVG3g8F12Q3Roqbh9okoKqIVCzA1Fh5kuUs
mREwuS/U3a80wtoyxwMlIhdAwVlOCf+wjn8hArWX0PVIBhLh3ybATZbz4tmCQNiD
adn+DnARU7IxMIgINtGyyxeuDlLXwERf3iwFGXG9rdFnZOxWFkW6f8H/pXmyt9la
Bq/SCWbeHpKgRgupDd6hB0rAVRoIVxquf9q4qdiQE+HbiPJXsGyeyJ4AHuvMuhgM
AdDGGW8y0La9ULiG4pWa+1IYzhw/k2dGtqCQ9U3wpILh509sT/8J0SNL20TZV6b6
JSFQpFLYadbHaqx808bQkv8RhBZXBrvST/0aCOI/JxAGdb+QOGHVrmkD1t6tB6Fr
vbyxuglWwa+kDrm9jrqsfe4HdrSEkvbBgBqKCid5uM3bVGjdVfa2oQqwwn4+oUCD
6iTWUkGRcHeDynGztFCdDlfexwiWkV9FKnYI49n8IawCGbILQgE1QqBjg240+f0M
hdfKtVoUaFFXku21KCvMlWvZoEH/5P9CiMQblugmKQaWn2tNtExTQqjAa3/EuOim
RjG0tLYuPHaKNwW7SuQIC0J5JnZUpI3BUAqPO5NKUWdgDDu5vUoLcWdFXwuCQ2AI
miiOO4qqKiKaE/cDYYbZffMBaNJtaHUic0GOo+LMY7CPjS0BbGbfAzMZLVrdEwQa
L9XUbihTi3pr8ph3hCw517nr2qdTRuLJNXPPrfdobAyf9GK+Ubd8wk2sxRcutRw1
QdkcQTqcz4EI44u42/d510bYQIXSn3AsrDcmEo0R4DL6WpB80T9dYhNLdoSmWU3V
AiQLnbHBx8DZG+fylh6UWwbjbSOWEwxYZikZKPK8rPFKLa5MeZ6HSgozDWABDTVb
xOE0nFHjrMeV02TS34YG97C5DrRqaG0hRURRjyAAPYW06EvpSGMtIzSz8fhodYNj
XvLGNXS2yI9OyuE8rSoDzE9H4lk8JNUmjjOhEej0wrbQGKNSB9VGs37BHqT4WFh0
kBraJa786CGhWukqJEFVAUVco61oAzHD5UqM+7IhUt8EvuizcSwgtRtXf+GuY7U3
M3iKRMAqDEv70OEEXucrtnew3Bi0APHXhq4UePgX/T8i6HXP7EUdNkIRNwD7i6s7
0YnrL7JDHS4AQlxF8rIMG+ijDrrw/HqzQoaFu8/JjFeLPIxibBCq2OQyBkduyrkO
to48brgZ3fSb4P6mWV6uEkuJ3eiD1VmMebM6RQXBIdPMrTLQR1Gh0GvCyAOzLh5E
SFLTA4xqwPXlFH4KAt4CBO2E3jAzhmIiTGqzRVQBazk4woNcDxNIkT27hLS7c34B
PWVYaLX0NVeHmO8gsAyNQFu2Mek4QJwwgrjh7thkEKjRN55OPodbUrV94QYvp34E
VzKOgOI8Za/mwQWBJy7f2qFbxvmvATSuccGFcwGQ3C2h3RXygfE4rXhEAGOwyRf7
bOkG+lDIRf+hyrhjYrTTfIew0i3pfl6wejhTnC8t5/EXWqv60frVSoPhmTqu6eFH
jVaMPgSbGd1wBmmao11tvBte00VMbAc3Vtb8lL3zBDJx03gftcFRsO8hS410Bgu/
Wdk5xPJuDaGw7CXbA1xplvCTazORJ+B701fuWroY+UXsKpiMBI6CQ79WZhCrzqRe
htVIoTg885AsQPV2IvhILWtDyMYhXHtqrplEulS0BDFPC8DrPTAIoabPWDnzvmwS
5eKdQbBVdg7SN17F2QiVL5JZ/2sH9aIfllRdzbPDZ20RONfL5VbyDugJabXdU7p4
fHP8rcdw+4fV9P17TItb2hVnnS1bCI+3YU8rM3qcBZXrWme/Uc+po0lPw68Psdhi
HVgzGVyypdbM9xiSTp3AlARUqtHUjbadpPz+hrmUT44yT3n+smsx4MI7ptEHuRX9
TNzk0EMscrjiAF4yyU75ogUYXSMJ047hgZRkuJT8bBB24WxPimfWllvE1JbZfT48
FDz77oe2iBEPzmZDSH7W5lghZoi9646D7Ysca5uJD6N5N8Y9P3/psoW2HG5h2qiM
fT5mT4YC9z3IwfQilPlQvNJO5BfXXDz4KnoBTycV7S4xFHKUuvK0EYl8a/W/P8Kv
vXg8F3G7Rgva3SXln/A7MYjaNgT9WDVfUFcOAO0xvRQDLoXPUeFNoybn+vg5A8aP
KGX4SeasWlvXCGpHy9CPGlMb+TmcsJe13w89py0JHMg89VF1+3DG2ynDVQeXN2R5
i/+kt4anXBuHuyBxgJn49atEAILs1oj/bJUwvl/uLpKNg/nDsq8pGpbuaw1vnxcx
58GjQV11fDPFzz7engclWprBdtbtjolP15mwT7xJA+MqP/Uf53uLCvjJOLcrLfmB
LzX5EQlEkyImp70D3zZRzF/Rd1qg2OksJVDD6DKh8m7AoASZjzOR2gN5R/Eo15oP
ymCd3DXCcBVTRrpLaI/ZwTtYzuaTnpwmYSwt8qV7B6AbV9aCxKeq39jQ7G1VLVcr
PiDAQX2As7VyeaUh/DibyTPbDUR/3inbOBndPfVNbY7R+jNM6Ct4JY8LJqyZI81z
1GGKFsj8CuzF1XTcTOJkVM3/ScUMwfQOrh6o43LGN8P0VtSdwAHpQHShlyRYwHin
MKefKnGOLb+hBRLoXOgFDMz0qEcbbXEla61v4EIDXk8389fmZEDj/DsYVSRafT3b
Vjt8LfHiLzXEAuDjkS3S1sZj5Twku0WajRKOZqXSseylxtguAQP319GlJP3PJmwT
qoAfT3+UYSWkazuIOsFRkQmSHShXoaiIjRHzkoe9iGvUoBw5LAjs6ddwxANo4krB
1x99XMEIeqQR3GxdJl1EL5olU5+5KfTeIUg56n/mSNsQwByUyw050iLN5w5JNb71
37dCtqQk8jwly9EBdycO0yHzidiM30CU4EchGSRFnXdEM+nj7kUoTyZXOjKOFWsd
iiajfXcwUadDTdGWbRlnSzYwNP+LF8Yx6OpRTgazqUhCv/UdxXJVmL9mm5E3M/mm
3KEV6pyh0iHQOTKr0XVQgMRggGECCVdj1AOnaPc6DqRiTk5FRiEKDM8eH0fj/3kx
3qJqka/hf8WqO3LFcEZgJofexxrcWGg6LXIslcyaB6uKkfABJX+dtmSwtrJ0yBFH
+ggjLmKTBxtV+7ReFsrT04NJJa6xynATsEz7qSRFUbGgtanUtoGAMptkjvrv+wCi
XXnglLR2JVbccNBMpA79/buBAwwC2H0FzMopKPJNUfan/Qml7y9ZGkw7vs0/R94q
Uq2qEgOrknNFAwF9SkCr9qfFP/2tGkeXTyGrQMUl+mB9IIGGsqOFulZ+hMZp+3X6
L+RQ6pG5T5unIgfnNVL7DAD3zEdyVl5uXQaOvy2avn0hNtesxYq/w5LkEYhvf+NT
PnjDWl/w7IS3GqRPZGcgUYcZgJY3QFDvNFhBa1X4zLPgHbDiUd3VarPy3S+VUPvD
znR+IXoNpRXiJGjlNaVl1EnNYni6Frcgq2r52VjeB0TnX1RfiKPH/tblzVNS0j8e
xHHl6vtWtkJxMnYoSw2rSPpAwLYEZ886rvZL71+iWLikQ2hQCiDK+CDAYcNfTtK4
sKfpDD3yokv5RfUWC2UXTZ/LBE+SMT0edMtq/59GKfOBiw3z3ofY9wc+US2GvkgK
6GWzJ5d17NnrwbTKmjP2RIxSOA2fH30gDfcXLGBz/sZIbElY1HIJQznkWYkcQnsa
nesDzPiCZQPKnPZYgs/ZIYtt4NaBSnK6aE+/j+QVkDTaRaMxTpmxC1n5Ojeb0zjr
Ax5tNUBBrtaw7xYDZOZVDCSM7I2PodjoNO/6bwyP/5m9MINc/zOJeN4LV8mZ1zfF
1GrbT2Ec2qy37Od7wojcBd+Ozi1w+w5jeEfDexGEUdHei3VI9idHXHkzsClLPJHU
hcQ7w91zYpqW+a08Lvdtz1GwSJp+eUckGyjiM+izkRWTlyK4j/N3egZWJkAfro/0
0a0dUACTKMqjfBuSboNA0QFtrjPfR9fFqlFBj2HRrMPoizL4rR+sSkaCplJL86i4
RWaNzdIXn+ZaZIoJfbBk0SfQG8xD2pjIGnc4hIOpHBPh4I7fUWwELNYkDij03YPz
q+yF35dVWCJLLXwd3akr/VMRgHnOhuxm9x89Y5vXW7h+3sK5biCmbtnFhp47WZWo
8qC9oIZ6dgECur23N477NuunCmcy66VwIlaSJvGzW6VH5c4zzQ8JNoZ5xcYUQUYw
aU9QehSyXp2DttRkiyUcZ3Qrr+29YkVmM4IyQveesrvtGQVu6Ey/y5j+khijTavo
ZoFfWxQ/HZNNR9IM7D6RLkqa/6fgZ7ENZ5V6nD3JBW/3LaE5LkoEU4kHR5k5Lket
jzFmDR0nS+QyeogYku/svbCHk4gancjgyhUjsVVSpzBVCqZokhyBHOofK/LfnAZf
VtojVNrQ9a5UPvxAcjnEEzZW++ohIUoNZq+wZfoXcYDErJRGijncNVhRIG5Q7LOd
5Oj7TNzgN1QSpFn0ZCdnFtcx8g5a9qJSFGxI8/h6SDoZSm0WpJBCOYRHAU6cRE28
ElX1Hessa7ux374VOqmtIlfd5JStb1PoEjiXCn1KfQ1tBXdTNaXYE6pLoU5FlVR2
mA9KNlh73ZZ+4g61M+JMONPQ5bz3p/WPLc8ARSkUIJyJAN+40XevaBQzhPOzOybI
HYJKAun1uYqOQdmg5a2stDEhX108STy29WJ3O77ZqmZAwzdekN3/JuUoiTMzNjS5
SJ6QI1OLV7nWTeCIhVtJzvHiZo8AZ0ZCnLCBUKTi2d6LfQs78sFrkxLRDZTdSTSn
mhKcDet14tldYuvMG+xOiHkGTbKDPf9588q1rQ8bLZMz/ztPiRrcDVz4c12g+v23
++oS6IsZWDBhFK5BN0i+7W44OYh6RFwZOCHzjv0OSQBvgLoNi1GqTlCzn/jya78q
r0Bw9mU0ciuvaXq0obqiK1X76xIW2tQxdH175F8Eg00gY5BvIWYTRrEx+m47kZN3
16mzxUmdlWJCjn+92Kz83sEdDKQFYM5vVSZq06/0uvErvA6hcbXlY434nT5dyHOg
8Sz3PKokvqjhAEBCo1RnZKKealyLuGHx5jOvBDWHUU2dshA6kc4U9AhkZ6zWMpDo
41WQvOiY0kk+pnshya3dOi77zHfzyI0UbJn7fyEbDpDeg48zRcx2B6fb9MQjYLB3
GxrvYZRfLTl5z44XuQ5FCWQQB1/S1R/czOg7DeNbACaIykdUDVmT2MWyb5p/b2it
36mOfYMW12gAnSICuJB6ZFdYmVB4yOSYQJeLzUszpJRAJSBfkVcZACOWmVgHQZOS
DjcLuvkCeT0NSJJVHAUfESc8lnad18WgfSooNWfUIwY/7ocxREXEWWywUruHXwB8
r38fQJAkZTXOT6+9Zr8jBJsCdGA0gCB0sWc3lf00U0iohWlH1kfPE0LtsXJdAMnj
Jzbkfgm0tiovProFr9pYp+9ZV3kiqelWFfPXCkr08BBe4PJujzfGtDNFNZ/1u62g
4336KkiiKJBe0oUQTZtloE+aBd4y3EH7GZd4z51F+WGB1CTkotBbJp4UsEwuRfXa
pUYZKyP78/ovWcAOBBPYlw/krODtY0RwtC6VYcsCMszJeKRQ/LrwIL/kjj+nzEFG
e8p9kIf07ndgawK9txOmgib6vu5AFVPdZ/8W73PKTRi8FRwjRCfPmREsMJzuqChb
Uj40jhLWddV0gx5IciqhQfdK8psI89LHnGd72gzpxYjhZ3MZ43XNubx1Yf0J1elq
oVLYTXAzphtjNT5vfzN6tf6Ddv0uVWGa8iAAhXCAAmqnrAUZGh1oT33GmYThdLDS
aWWlx/knXbxpNqa8V+T7h5ndC5JCgDoCdgs0h7KJbUJsgIfHf9fehpUsh4eAPXMB
J6PAkkC9klgVS56PMCYHLLjVEny0zVhg2mYMTY7lk02sxjzlaxGpczmNVdgle83l
Yel7GallQLuFtpT18SUZ7bKDbEUo4z0uH9NiocXHJXgUc9dlZSfGcjvBCj/yUbXB
A5HM1rnPUY8931q8JCG0mum0v1ZisLOf5J2BfnjISPwCMDSnPGZSfzCYJZlqn5W4
7HtAVeVHZAXXeLiQWaBp9ZkHgi+MUN01KsykMLoHkyCubqmXBB8TfoIi1/iBAy+d
Mpawyf0pY7h8sMvYhcyEvikkdukOP6c/QNstBax3R57eLhn8a+BL7Wzz+QJD7niU
KIbe56qnSNidctYzM8peMsNPexra8TOmJDFDORcjpbo/QKLMrAmeMHbOgiPgEBa3
V7r3jcaTcLZ+C9actOMIYFPLsrRGahXSdQOuJamuJauYVxl2y4DslxjnrOvoPbpL
zPTWH8snCnjqvtj0Nm8igt898OZkro3Q9VzfW38Stzelg9FSJOTgn5MEIn1QVQFO
3sgtXU399TCjWYf30WSrJRRsbrToTZSMO8vAK3DFcQiFgzF4i5IXKt2J8++UUS6/
QhykaD3mskmv8T+Dne8FVHmeDIPySXJGz8EWW8de+qeeFMWjB99dQBfC7YO7hSoZ
ItXlXeJuNgvJ0rdYxwn3N7tKmlLi3A+T8kFTRj7WR/Ngcolc4qJH1yCj+fR/bGKp
ROgGIexv5wfuA7DJ96qPTSZMGRZe0ft2HYqrm2iRPdniCueDjPg3kJhNdZHV1cgp
hSzqpZq0UDW0vZdPEbwIScYydd0Mx9QAKmeiEO9bjRPXW8FErG15EPb19dA0VcTb
xJRmYv0+G3rYi/RDf17NLeyy5dsNoXIad5K+haqAmqCnHzXwsRaU3Uol27/1tffK
AJQ3+gvT5MJof5ezQyCSsLs6ZNME/eGMWR6wYdwhoz19pJvvQfYWvVGHnCzHYouP
/N2AodBvhvZzjnyqj0OtRVsIETYAzymZxOg/4/E4mg25mic2ygPd+Sct9RZckLVN
/+LKy5rWTPHjK6UXXKsoj6s2pPQk1+tyHfOf6EuxWqN5p0akZdF52rB0PYJ1w4aQ
R8YFTRF/CRRX2iI7bRK9kDfamp0lv8NK9qrJ8UQk7K41qkx6YbchuCmf7A2+7ISq
BamUeCaXg7clSiZwJ/bkcWEN3sPNnqG+5kVMJpd1+2h2vxr1uDM8ys4XDHpovmBH
8ZRmIoKGp+8ym0q4m69TAgcRlnQVrUPT9nJIwIEBFWWnNPI08PDe1Lk2WQ+9ridu
48eR2YKfKrVzVgqsw2K9FrIwBnVsNtXeAUoLxk7cmEyh+A4DKljJ6R6V3+8Y6qzV
v1k1GhzBpF7Sq57Q8vGW4slNhqZtIpEqKJEYU1I/wzpywNOd8/QDAniTWx3yfa0f
IwHQlW+dz8WET/r5iKRfRtvrhoHyBBBhr7ywrgdy++MqsJS9q6jNlTABBxUzpWIU
8ge1nUq/hVBcEQ8cOwiuB8dtvwcq1adutbRrSjcAfa7XAnnTzgKb2plKp6s89z86
Tbopwxx4vzJNZubW3RGPbIJFwMFZK3KUzMNhEE9h7uIoDztOnF2ESUDAYYacVs2i
JDAUNGRKFHrw5hbzf99o0tVcIj+OutKBhhSnrLTBFA2SUkywz1euH+f7Z1R+n1oB
cnUxJkiWDgORV8nDMVw/VLf/tnNpVAmc0n/KBMrU+mbmHLUV3TFXXIXXQ/cw5i4L
nBdmgzUHzoCoxprhBYfssWPcIYvpLvYwQw6pHCbfw0idQhmMJNqQ5gGuDUfAbMay
k/sLpSrrxfVXpuraFzxvpBpIqHGDyRenFOy5b7O84XrGXGtn6OS7tafDHn2r26mf
gm4roNvJF6lyvYV+Izpo98sTRKRIJfpVjizaLm7TA4nAt08cjSQEN9vy6ZEW60Le
ytiJEyvm7g1SPgju1ihoIWM5uCJlwY/FikyziNdhzo+9S/5ZhZOzwMYrwIU0/Heg
dJcwM9aadaEkmYlHLj203n+s6v0SWmtgxRYHvTzEpJQ7Djd+fxPMxQJh11W6a1JR
sBWF4dP2Ci3OMIFaWEMdHvBiwU5LBsMG6YHOVSDjEqpRm0ioGFyJGldLDwfeUlz1
ue9+SiOFcV+PzGXVxAzx6K8c3eBSOxyLzGo+YH74JnTp0zKgKZn0eL3p4NtcSCKl
Qw+3eviFRH0DP/MNCtnhWFP0vVFKcuasrmO2NlauF0u9Zvigdi0UUQKmvTBhz5hm
4UOgCpnHb81U4QlNLy3obttJwgW78uXqe6Re20hJh3twpPoVhyiKj1A5E4Hl2KX5
MuIq45t0ExSPqeiRXq6ZjNCGDuJqbUgQDRB2mj6EA/NtCI62zd8THONsCkRRH7mK
Joqj4e6lObGJtmEFML+H1xQbh5e7dMdrtRuShy59xYMneHUpVtfgeLH0RxlBC/Ty
Q0U5pc5qN30suk5lW4GlZdI68qTcbEdujH265MJqHGqTwKxUED/nA6hUSH6nxMJm
VKGiYDL/v1M55iOxB+MekGDCVwxQxUJdRAz6mYpO6Ww/OKeeSI+UvtUe0sAECVQg
kDfwbcEm1zAzDmmuH1stW3ZBQWeUM/OvJyLwNT5C0L1sFmedUIJOBS5NYQC5L7CB
+acklea46lol8cYh59G70duQcHRsZKL+CyEk+da4Rk8GoEHeV/qOdLE3pv7fXL6T
T4LEFAZ3APvw68xclivznRNGMMnp+vZwsp1/mDlbGkVFWMJmd+CHhYzV7D8YU7T7
Zv3qXgEdflbIVkEiADFWHycPOLooBl+ILv+wIVjrfS+Vmf/r6Ljyvyx7J93m80zK
GjyQhioLeRhGkzgjG4nALJx0NC00tXlpedu4CdDQcUbZkDIJLt+LBU7DXbWOi8qr
P93KszSiAWpICE6baJWtPt2IVeUMz+4SQXiWFjjnP/qLx8NGiAFHMcR1ZwMpTl4n
Qekf7TuxY10U2re9hPIsp+/xl7xW2usoHwYgibSLP+0vs4oqOilWe9Y2mixZhrfC
cVIAEIbBYjjeNv/lzQi0lHoGfSZIVc+tCwdaqjTihodFCg6Bj5QXQ9o+IZS3kVZN
jCf6lcxoMLH8GgtX0FhpxSWEbs4dTomLDfOnDY/r2B4rsh9C6q3mmrvHYmNF99VS
ev+dcsVaK5A7Bx6RbhJ4/9Mp7Vp/0ki7lC5pOCG2n0vUY8VimefL5Z6ui4z9KPmh
9vCVU9Lc1H4C7+UNtbWTzfaMeu2IjSVJfZFIWUX+kTroKTr6XpOpjBx9L4hNFNg0
lNVHCAjE1EFY2BgJFkerKjzedEvKtM0Z6hLT+Xg3YOTVkzlujYbv/GeXSLmN7Ud5
5iSBjC4bGOO0GKhVdcwP0zUIgpbyw9mzV9XJXTEE4FGq4Cs+AJpF0LmRUDN6cBaj
WXX22MVzF9UJcejOR5JHeJfclR0lGDEm0eRgaxfJ0BsmQqUg0WPLZAvp8DPHvUuE
QBAjyPOwyac+C4ee66NLk+2T+nOEnyqWzuuCtDSqHcVn+LTxRHu+ZMzzTOK08J3L
MgkVV7hhUccggbiVL9OG4uwzrHeuPNNVWOBh2cJepTsj0nNLEDr3k4KAmrU26Iop
AS4mTOUXoZprre97iIxGSemlGwgzIcT7z8ZLI11PRAMS7XwvZNUWhNL7TC53ic/H
1LVbvIjTiGu/oWca2aBdqHYUhCm1VoEn8djqHr8TUlG/wZAAUgutx2tYY+RMnXqc
WqAggGqghL4S+GeIPCxYv4gi78tnJ90RRSsgRu7QwPwbpalVfNW4PZIy+csH0PgO
PVlT3hsWFRZ+nSMcc7XIT5hAkFUbSP6yshAMItvfUHvwf3wYmhOXENsY9AoES0Xh
RuIsYoEP/FQ8/ldSVlpGBxQCFrnNvo3/l3MuiomqDqUWngwy4TQf5lb8tgNgOCC2
7q8K0HVy/wpjyqBf3Mf5+OnK6EyRaaUYtcddJDnd94LVCufqhQvyoruXWCCfbfr3
5iyrWuAFZL/qHXQu8+swuyyAj1y9Lmj+3nBLOUtqMMUiJZkgCmZ0DV3KymALQ0Tm
8xkkjcQWqi+W1/zWOdLbTw9BQMHn2awn8mF5KKK9PJhcGS/1VKSuIcYOjh9DF9u4
6xagaptyR2CQqtTMNLnWJ+eotPPl5MvWuIghZZVGm/KHHvQaSfEyH4tvHeDkVEFy
T1/QzgcvRgbR+Gxe7/ENn/T8CGGM4+L4k5iBLU66HA48AnX1dWFOatd6JEoxtsR+
n5IfJyQoVcapevsG2lY3ou0ZhMWfCa7RdZmO5IbZxcNZhVZyK0Q6C+2VAkm4JCMQ
s03uY9j90TLItEuyO15s7Wxg/0NYO7id/m4DdMhtsXnYgu6VGDctrAOy+liBo4ve
s/zHTsaPXS8rwBBEOMIHmSsZB/X3NKy4eP6KbHznbwtEtw/x+MkP7afr9fytlc1/
68IsQkvWh2IFI+h5gFPOtVWS3gImG3DIpvXP3jKyUrazV/ciQqSoIl7P8uq6G9iW
eQNztjcSqO3Erl+YB51hRzAXnonzhN3f/ZCAG+o8dOgYRalYdAYy3u2EbnpVYMYg
c1FAkuLqNiZ8ltvnuu5Zp5yUWRLwdQiTchmFgviwwuV6L1cRaswM6+SVAQRQhNfm
HZsVDGlsoVaqIb2+lQB0Wd6V/IKpn8Yxrexb3M4wLcKlZco3SE4f0ZDQ0981htV5
Ndpc1B2R/7U+aqoZyfLMb32SQEmaask1ZcuIw55VgijoDDCZPIoceP22rmKDjXkt
jqNmAhm/tnu6dFSFnXomLZ1hsmMim+R6Z2jJ2vGWqKL34plRAPcNqOSliGxVxmKO
k0C51xvWSaRZ855+yjSKwEaD1eGbNCppktVZvrUcVMe8bRD3Q1ZBXPu83H7SW9vY
/mi7KU78fmOacGA8sixC+J4HEyvuOh5d4sR64+ClN8fGVw4stBq6/5OTmjF8r03D
wprDI1yUTIlQpkpESaFFz5Aj8TYVR4g5uu+P61ERDnCjvccwRoqxoYB44SUXyEKG
vs3QSnKgGdSelYO9vd3qOC7szPvMyG4/lWV1OzXwSQitPbRPNHD5hpYjLIjh/+dh
ZJq5NXt/7Vs/7pzb8PpRw7X8sty6aai0WoVDZJrZ6usnU2rxaDL8vN6mD3m3yCHI
jO2DlMRphVTQ/k2xwpAqiQu6OrL9G+cTSJuU/49jXs34FEPXt9FzisHVfIUigcT5
frGt4ENPRXToQ7njFwHoWloZ8q2a5GhZqPdHTFaQV7xYIwRDviCq8dMtVgGKeOzx
D7M6pcdcOkSZ/R+5+HNz4ZIPx2sBdd5s85hFS/F66AhEoNgAlQSgZggMdJyyrtcx
NbViPft5YBR5bNvrPKkbts1z1Gm63LEeU6lPL1Kwh9M89MCo3X7atfnGWz0jOaM1
7tz3lIiR6espp9q0b1+8Q91sIsnMDafFyU9kiB3OUB2mxXvCEHStmJmVGzlo/vWR
NEaHZipH57AgGw02dECfc7WwZlML6cm4J70aieM2BcMg6b5+pfRkz3Pz+HvVqfvV
bs/UQyszJTgqXbGPodIaI57aVHD3cFp401+QlxlgD64CGBgSN8hEggME+cIsew5d
cNsw99UITE31EjacE1epFtDswLq0o9YBGc1BS0Bfa5HDntsxEbwCgp/xWJMx7y2r
N1ohl3meqcHFobhV7PzPRD9tmUzhsX2+dGl8Vt0FHDV+MbgmT4lla+bfAY5RtLjT
XLwEbzcH920Y4YG/eKrrqpmtKibJamic7bk5Yeyc1hMb2nY3Svx5O4uz31AR/Gd4
HDyXm0OAaZauHIdLgU2FRzOhduLhf6ang6caZNdXI/g5goyj4pADIBq3VBlC1M/h
n9aOI4SI2kDOreZcK+JsoUgqFZ4RDm1M3uPWYXHO9AFJwBuvOPRkVI1/Roe3QiZ0
B/kapUfpqg7od0z/Qpzrr+jv7sOFCiqmaeu7NR4FRn+cwHMvmPFn53X6CVSRkAai
vHZq6sQKrtlG6nvfHbhIYqeZk4l3iex09zfQ9tf6yS82pq8w0EEMKMv20WPPn1rK
PojjqRueBBkjlAXKBO8Dw5xPbdO0jGboMVa630HxOr/vxPu1vkGQhU5FWM3Rs+KC
cKqL2q5SJsd/jtzXlViKrcbB/IpzVnGJkdPoJM61i23X6h5Lr+Ny043HSy5lxFB3
vGCvZhUsKvzd1x8bOrMhPSjScs0BxeENaepVxnL8wnr0gxoVvB5A/NLAuEIx+oVz
ORfPg1g5s5oJ9bNBuJlI/u8AJZV/o24ww55ascUSN0oZmLnvHJKsvbHdQOYhRAm/
KXCq8KTH5p+3XkfkdcgPDm/oIeVMZHOXvGNtoHyxxhLKLr+DgC0W8T33a6kFSsaB
M5Cut7apeb078uCf68t4anBcKXwwppIDxz2l6BateaxweeOOtRVcWd9XiXaIeter
Z2Y0EqTlgtCPEaLRoC7mqmcpIwm4eRcCsbzdmG5Nuc/ZhlcR3OnN01lnVvju/gLg
buXkn57bO0tSCXv/5emzkdHQnkXIaMxgUFe7uWOO+Ja+RvIxitHuRsDvg30i3+P7
N/0p8VfwJWWSMx0zmLKwiQuIl9YtdYCrPfFAy+e3aW3BlTNcq+yxW/qqynRfSU7t
W6m7/mgz4Yr0tsJnaeBc7OA4BKM4YggMMnHdAybKS3qK0xFs2cyDa4di0kuxROo3
SXx7zGrSx1f7LIMNJVvGaQsQ1gP6DaYFXeNHb7vMHpyP/gQfXjUu0m+oox2UdSPy
85UYbu41fFDNvH3SxFXsrv30I05DUzN9t2iOE01bIgCToj4DRIlD0wQTVjkDFt/z
JBqw4pZufcfv7gwttgOwqCG43ngQmY0iKn4yRy5DbfXTikGJasf75rSWDHmvwRrt
ZDvCpRXnJVi1Iql6hnQONL34QoqX+H5cDXWjlPNGWrGff6+s3Ly1OU6kn/tDomZ8
JdbXMdwiTF09GFERbAe3Vk9ulWnkzoPbiAmcca8d7fHTERtzjEcnECEhDTDvweDK
VWhAoghgnfrFnm/sQ5VK0uYnvHTuazmHpavHRkqPZsA5ppJD7YjfkMcN/bWAp2A/
yaf/l6pZ3JnKHKBIJN6Hd3XYgpSZN8iUi5fwnt35WUvyIvW+X3Z2ozrZBeXgiXKb
lt0p6DzY0Rh0rmHmjA/gAf99KWUJm6/mcyFDqchyKpgQMXvxEhRnjPyo1KdraxQA
H8l7Mn3hh4/bfino9k+fKg5H6vyau4Is6RScMOWPGWvrKHskzx1Q8VsMTZe6mxEj
C7VzpfXcIZbH9QJUVKeYAAsSNDAUgdRzXHi9jN/b/Xloq3I6LlYZUdEmnUcgF4az
MZpDP97QUCxoY9GZQpvZIPWNm2NA4p5qfBhpTKJMbW9OtRPCl8+yilZKJljGfjWt
TqQmrgOYPTye22dpLfEM+Vod/SNKtB0jBF7v3HcYcsQbJHxhh2861AQUBDfV4j5a
XODGL9x71XuRaSknCnBHMjq5+LikypxmdT+SYI/J+C9RaEJANwGtEFzdIn+/EV7r
Rhwy1gdys857zCnFZMOB2iGEiwu+Ka1dwnSUu5HjE3OgtUndkkXoz/Tfc4uIrhg/
EiloxovEDx4gWl8jvZqCUtEcm8UWNtKg9KljchhGvFZ6wsH7InJvgkUEJX/2ZZeV
A5u48oTcptVcs8YMVD32U3y/SodT8M1fveD2JMDaJMJmnrSsk2o2ue1h1d3NyvWf
gonCtJPDl1CXKj2lo0EQuARNNfzLY834sjo18apsvZv0C1ltdq+6Kt8hv68Gw+TC
ftfFVnHMFLa5jZP+dFa8QCacrWtT/OzKhR/spVU4rtvAlpcDxKYXHa1ODygQOiWf
mG63Ls6nHvG6kR/5IotnIsAixlqis37oWGmXy5AkMTzoFtvPXdP9MxyiL8IBwZNv
heQFl/9Qhd9V+Q7xecf5+mo7mgIBOcvwKGf0eoLifwIuPT1d5VH92yuGHDMhPSSm
BMkiYL6VzZWwOKWNllAR1OoqIOop6oLheZ/ZN8aeyBJ2oqPKEZF8W7RNGFhSgwDe
+goIcqXaMRLDbgRhw0hLYwzWEEGP4uI1tpeq17kRkphxN9iKc+K/uDjLP1KjQOOA
VJbh7Zp6GcAG8ApcDVSx0Xt33nHMGjcllFGADF12GyhK5aykgAo+pwTrsq+qZ3za
Jbe939tWF+3SvwF4ZkUKhiHiL8LyXpsu0RtNIc6YGIaDRXLpOVQKHFLaaXbnKWMp
uJJ0k5vHDGALP39C9GO9+k8mcT+XoYW+MxyVA7dDaNWM7/sWoI6FtLrdQ6tPyS62
KMx5iViWJBfqX2x9cS6R7IYpynvl97qsHU1xOJPnoRDOuTTLK5rNGN1GJQp/p3Xe
l351cljnYlp8YPAedrgih8w9pGQnNshH4qswOY38xmwPWxwsAJygmUITPnIMotjm
ATNpWDfx6CAyJ2MGBWCjPC9r++k+jI1+Z2f1SRJ3+C8McxZqne99QDucQA+hvxGl
KtSyaIHPSQM9MCKBElq8YzLMY2S1bqduifm1q0APToU5YqgP3fy1i55ZKt6yPtW8
XRlGNMTtJro1REZbCNV9nTejS97WCztUFfJEAr6FexwRBSN0TFX41EA8VwD85Bao
voR4PMfW6an16OWolbDlLqxwBj9+/IVuMF6SZ3qwYM6M0CltFiiXfcbGfUhIYnSU
nK6yYDT5h2YmLUB1wVTZ6HO/81MJy+r87NpsY3ZHSY/f/ObkPMqIXy53aBP14TzE
hujTttNzi9UoLDg8WJbkc4dJjiC/BQaXed6A+/yPHU+k9P7jMdAr0Bat9OMq+rIQ
AVf+tf3VSkFafabXhntWQoLd8E96ViR0d2WyWuh4K75loQ704fUnt/mc0cNlyuHb
8zZc4N+a2CXNCg2H98MfkytVoo+vQteiic6Q0VsmSX08wVUYY/XwqWnxODdDeYc+
BDqqQ7b0uopgtmyI+o3sNft+OJlUSa7N145OUh9EK7+DTA3BiPk2bk7NiQ/+rSua
wRKXicJry1abZUJg2c6CsPiSfmAnGwBqqeU9mytwMJOdRfFgGjneIifM7f0jXH/j
Bz0CLmxOFrDBuEMHr9VWRXdtVDY5ZR2EA12jNbPE91Z7nZc7bq2ftmTnaNru2V0t
H2az8wFiogP/Hr2sk4lyoBHSKlLyOm56JnZWpR/E68j9cEOx9/XByWn8XypfLaQc
pLxa7KUtbXnP2UC1I3BnnpQowBPWLcZN0aQN552BP3OPuQUAaopR7uDfRUCXpra0
+f9HrnH3ZDDl0QMpM26pJOkdhqJ5GBQy5HHi7ovYAEzk1N0k8bmHT5gRoqjw1zfK
xde2XnvJbmhUOCnklxfO0OBG91xsBgCTfsx3FPt8kFz7Ip1K7pbZYbDowhqqgjhy
cZD+J6L2Z5LPXSORv7z5pYwm8MINXv8Zm+DU08qw3JLLnRzEnozbRyb5kMWxm7SV
iitm5BxE0NLLOFsiXVHWZq/DXFtAJK6kJM7ZIfiXly7GBgUsNwwjq5Ugr9QDjIsn
pMR299WTqpZqZx6JFqZD5tT1/MH5QbOaHQqRj5ds+54AzNjxdWpfAX38WFUXnWpe
exzkkCohZtTCEYgUv6pHRRHw+cby0WxLU3UJ+VajY/aE/fAV51VS8ge1I2sfxsN1
2+1lWUP7o/nlyXTNcHsDJyDgceRUQ/vyBt4CepTwD6qhoe7RQC6sbjWdjLi7YDZR
IVdOX9XdRtvNfxK7JbZj8IhqigYOsxu7THpMu4eto88/7bHip9+XRGOwMAJYEdvC
cqPF3juG1pPbezYWiGmDpce6u7+4ReVhaWtHfYp6690scAS4chkC/L9RiPI6VGgp
dQ4eAUIU7Z+PW7hErK69WaLmWMz+oXUUcfK3mNRlmsdqLx3RrGO3lYkJNF/CiVBp
a4k7/aU93Hizxa6FYdSfmSJXE+c/u+PIItTLX0JucYSzaATay95kZ5W86fAr4uuT
zyf4Ia8qSZ/t29+qYh/3iWxF7Rnp7kYbFN+RCthTykrXor7K2MnPxxQJZRoHDyXt
K0PnvJO589YKxI9yMedW+XnnXrUCUcnAzxdy8+XtJVyBZ6KXTxV+67AjiOebBrTR
U/kwpBWpz/zOJ87cAIx/xDu+4lxlttSIJgIWVAynhoty/rzPRxcugn4CGr66goyj
YEOYHOyLtdH9ACce+UK7ONzVOwpNuRre2/ZOOFHE1J7kLQ2f71UL/9YobQkv46t6
6eWIz1bj+/+1lCh+EdoI6RwQae79aTf9lRpFMiNKmILJOcLu64XS94+u3YGic6aU
CwRz+OyrJEAN3Mi8w7c/lSdnjlC1wN3lN3Zp9ysBed7wVS3dWdFxhvARxf5hcjXG
+KgJPXs+VIBd2V5auQEEnBlvjRBwOV0LG6TjFDOF6OY0DsuZ8BXNxyNHv0MGNVHO
nWswJFZGxR3e2EcdZ/SJOFPfa1fPXCFzgRyW9rYbuK6TtQiAGKLI5/4h3vNR+UDw
Qd8Mm20ZTAzbLsDDYGkgET2iIDPhLGnHJa8fC3lKFGYvPMIAIP0I/N9O2THXzqwc
QmandUfMuY6CJjReNzAZXQAj2iz0PWBrDc+h1Q5baQnXkCs4vkQ+Ycef3VC+oMjc
nJFvGEGd4RicX6Wof9LgNvUiT7GvuIHue1LsHbzRJ95CXkmlSTMLZNk/GJs94ifs
KT/33xcliP2HUbyIzvEGvTardyGGE2DE/cLn/bsflRX5B/t+DO6RTfAUlD3Xonl8
a0h1/Om+R/5kWJB5kxDrPYRwlo1VMcrnfxGW0UPHtdK8vE6QjLnJYOH+kHbc3UPG
690EV23AQuYm9vfjUoPs+M27bZ8KaG1ogtGzglXay+o4AEFHORSaQjradYzOfqq6
stlyZmJSH460y62JC7bD23fXwiFhDCYx13hYMgqiTjp4difRzIO4OgVneotL2Imw
snTbV5vk3ojn4MBceWsVVXUI3huCfT7w2rWGra5xstTtkDHId+cGW3zoaGYePFoe
NWHi/nCyYzsN4Wvy0SC3lDgMMb3SBDwvqG88pTIy7ALjy1YHvmO3ZPQ9QnkDxle6
bo7ln7ktXnllQ7+VCRXwHsrrIYe9G+Sbqsk5mgCkS3IX995kyiyNJmaExxKgvvps
DYA/j7oJksDLn3EpgNBnARWSJCU3pxfmtZdqjGECeVOVCj+h4iH1Z+Qs7UNjaRKg
HnxwdPBoUjjO8QUSpiZF8keqpb0CIWZB/HmhGqmTUs9lxtlaXxPf5WBbE7oZ9lIG
XDPNBRMZWorkryjlZ7dCZNwOZ62ltFBpQDW0JXQc/7EDk/tf8K/sOazkc8oCgHdO
Ofs1g2zi2ihTgCfwHSKOmK4rb9IUoO8d/lbAQXDXaPG0IbHenOL/qhR4boMcC4dr
iE9FY7WfSLaPvlFVx9YvPXtTmQzNvHip5hc4598gyJGH6GQf513rd1PL9XUkASmN
miv420wxWyVjrefsFXwZfl54fj35SAHdkBsAZIAmzrIF6TO1dytF0KrpeJl6Mnhv
mCM2zay/XvCUtjKZkY44+iyb+Gw2c6Q08j3Ej1oavwqq5VGTexaZxDacVZJj6f5P
Kmf5PeUHkIxrxBUALvq/Q5EluvJLw3lhCdnL4xdpK4WMOL9oVhCPJ7JwEkhkdXRL
x1rGzylpUJQ2PEh4J4QZkIFN86MsbkpYAcxPv3me6CEc8oTFtmlspQBnmWDXi/af
KOa9obbC3/HY4z+9+sun90WkN+0SQbk8PdkX4OiaxnlHJn9pwF2GsryYuwkMcvXK
ZyjZEf3Wgb6Wkng1BQvD90sERo7rBEj+oDMFsDVjXmBt2UHmgw19bqBJWLzhry2p
jw6r4akTITJ4RKk0uGz7e/tmC0hYamL8kIkUV1YevROb/9zzWRskWc+1Z62nM8Rn
w5X6I6mUfxcgR0zw4P8K0yzyILzk1I+w+X99jysFXla5YkCxorb2L5MDlPKtnPbg
yYUrtPCHpFj22b2+vAH9ft2k41HTrn2IsRoUYe5M4t6TYheKQD1iL9gfAYrXCFcJ
PK2NiOIP6Offqv3xcKR6JwfFt2SUrnCssHJeLVYtRUDkTsYvwlqw1wJUGH+Zafg3
Ri+Ftw8HBJovod3K9RH8nNRtdkTvJEj/lM6fz7r2N8x0rHjHrKSaKxk3z9sJ0Z1K
WaKXcoF0Kfbd6j4+Q7at9jI0Ll/8li4wVcBNJQW/8aDaPF2lpw7m6Nftegj4Vlnc
tnSk2rEIMOnYID4P85vhKF+lDuCRoK6OnhT2EvyMwTxDRSK8TlcDJRdoPMy9Quxt
HsGT8/S9IvvLa0IY4gM0+IojEDozKKIjXbkbFxQQ05QfCZz1J2Ki39b9k/mukFZ2
R5JPdS133GcL1HDeEZ/tc7Dinj9/bqfdwy7VMelp7tllk4Z7DaRNnN2oXTxErgBx
RD6/OejWXfhaxj/5x+IWb8KhaTnldOVFR28DJQcGg2DuouC/ATbuLX3YJvuUI4GB
lukvetwtWdrVRKaTx23IA+qr/aSPlTXUA9Wt0N122X/PjGhkS1s3bNUxJ1Fh61nw
DS+MgY5GQT9M05ZnPY9u4nlLXYHhF1x+ipPuI9gmcidtyU+i0xVjSQqQjAhN6Sph
4VJNaiXTVi6t+1yoZsnwMk92h8XJqDpa1Hu134L1GjydKrv8n6ZXg/xfAN0B+hoq
rusIVirXH9uCH6peNIzPyuBf77VJny/xpyYzLHvD8beCO8pU33FXwpxMI4jb8rAe
MHq0Cm4MpTTq8px7yZvlJ+rGVjwiNSbu3k27PdgSEUWHWqyC+3rk0wYH9A/MKIaH
1j1LZ0dD0Vgi+wjs0fVwlop+ACvEt7KGBv5LfQazWppr997JrLSoCrDb9K8IWF20
73tm6k6Tk1v9nyxdfwpgi0XhbQEpzQCGZRuY67YYm/fYbtmBOZoUlIpuw/dqqf5H
EH/9ZzTry9FYhTcjBv9xFpi2uSXLW+mzANtVSBrwenLEo3gubuUFaI2FHQFiA7+9
AqF10u/6NgfiM5CPqbJefxoAn/KyH2SqukWc6KUTTHUoltxoBJWSw2cRBppViMjM
t6ZhmgWT7XA3hDSO/ljxaffY/MUd1E3VW6IfSKJs+LK/EsZH696DHTgkz3T5gt2v
iFIEyyWmckVCHb1exG2FnD3ouaZA6LSltm577wh5kTVPpT4xP3s6OGJ3sL2nNx+K
VNvtu6r59UO65gCvrBbVFJ0jykwbbTpkBxp52dCOmEpOqHqqGD9veQGAOL9pe36r
8ILjzCwEYjv8YwsC3EC5tr58Al7LrYMPM/GZbuCLA68B2OE9IkuUl63KYYpipVHA
pgUVTivK8c/WXUMZHWsDie9sRSbtF1x7jVLRUWNGKc2w4mbOV7DBu5TCScm18Coi
ekCmTOSO5XmRlCqO0OgyYXWyCM9qGDkhe36soCAdMpHI4ipOOLMWiMeePrETVDQ2
H8K6EOx9+/fAdEfJtQBtChjG3bdDs+Obv7H7YKsIm2u7fW+A6TVSdjPj0BCxs2md
Jb5LxDuSg2kkF+191ubk8XIHNLl82MJrTAA1xcoNiR9Regoc0sGFVCpreq6G1me1
8VJfJVPs1Kf+THvodSLSxbvuzbqSQxOiCdDjttDEhg7p8gtLQTYQRVPZCXa20CfJ
Zp5NyW/ufY+l6I5aQsq+G2El5/5MYOX7XimGjfQx5t1k0epp04yE5SPTlAC/wEZZ
JYANVZfm58SQN1+Gp2Sm0UMyPuZlqqMDfFz/Qhy4Hz30MC0iuF7R24W+IHmhoP7O
4vcKuv0xk84WLniUlBEGorNI1oo74smM4RRFSkmgT2ZSz7rEAvcWffIemfXsTRza
kh9QUlZsvJtBjNQE+r19g+LkLaXfkrJ1c9jNPL38+gMCzfOtTBCy0Wb4tXVg1+3S
vF1tqrY0M+3aBUY2gUpAiJ2h5I/Uhw6kqwxLy+BxkykN4ffFd4Kr0a0tpc9kl76J
5gkU+ylOfKpA8MlxCLhrOzks2Su2rj9c8rXRR5Be9JWm+C+Ne+JB/N2WB9I1oTik
gvNX4+T/BnXzDyuV/OhKqjsc9EKUHd+PKaGbtxwv24vWkpdj1mKBxAdzEyab0Er1
868uBqD0TiHwFZEzqeVWCdy3rsNzbiGE8Ajj/2qp3PTHfBR2ebfoDAn2w5NETskH
vp4mUrzDhTT+Ac6RPHaZNmLsK3qUdj0kL9lqCrmw+knGwvtn1SBs4IzEL310WOXM
qUDnG6MZNnwC+putApFAx0dMJbtEmUPihlAMLb6JDqmD5BgXC1jC6px1GIC03+rc
TpNoUQlxw4jf0MxUkpelID1D/AYVe1gkUz2LAU/90PEAPBCxmcZ6Q8ArbrJyfkhM
8n4PwlV4IdBaohJSFLwDO+nFbJaB4l/d17EhZCPnshUp/5S7SpMuobkAi4U4aIkV
//WUEyJdPSaQ5+kHUj3Ikd4YKmi02jLDU6rngPoRjGp1ut/56RuErdFGjKK4ivJX
9KykzUGFG6LxnQK88asmWbznLv11pezwu9bx09E6G9zXSkfVX/2T7uQn07Es//+o
5eVlKt5xSrKR+vJDyZRoP8OGIIC2ow3Xj9u5KhuycbtGu8/quI8MRmR9KPoAEP7M
fIOwrRy9ZLz+CiVfw+jxy8DMArES7C5gaJ0bgPL+iQEsikF0URSoPqGF8u+RNKS1
hG0SFwvRCGcbOIG7k0ARB9ZMW65gh2xrQOZ0iwRf1qDexkbvRnAWLafdm+iIjPDl
kPU1f/Q3JA0MyovJnUJBVSVhJVWk0RBWkp366p811CmhJZwFVzEsoStMOxPjYl89
626Bs20SAArL+PFoaU7bXhufN88XOp9/Nh3K8nJ/4TpueGrTP3/0jRUHZm8yCVfn
1Jd08bmuxPK/q95qEBGOT18ndvTjqiiKbQqn6NC/or5/14o8NRnhMir7NmEG+dZy
2eHdgzYZ1TpIl73DRw81UhZl1vemarsGZJD9wpn6xHI7rv3IDk22Lh+ZsbnsrS4N
nSknqDev9Q1tiy9Xi2ZBwg361hhxdT7uQDFIr6Wz2ozBtiuRn/n2ddY6ILDLi5QQ
zf7o87wJuV077v2f3m4ZCCWLwucwXKfIODrbET7/N7iSH89T0MPtVyUZ6PoX9dXD
ulHAjWEVMev0eCgkGruiWxBfi8P7Xhlov6TORU3zRmzHbQXr2e2UUXxMw1G4FBms
SiWmeXU+qaBSDrMNauCRJOAhoyAhsxowC/4q+32D60cuWvjDphFQAmlkTW4ZyhTj
AMIi66c7+iFfJkMiB3KRd8ixgMPkH2IhTSOdxQZ5svHh/VhCpqW0lJUFP1qRPDX9
Q3LAthq3tW9kqes+viY0C9Lp2jF4weIpS2FUWtFtm2qBKlNXzzdwUyKAp/4tzeCU
77Pj8eYqs2cRWKXX35MtJwny/8HIzcjC5wzXADWGsJXKY5RuXQiEo/Qns6ls5+iA
3Da8uLJo3A8iyR5iVSKUHIt4SzfJAKsnlZ9h10kWj0UbXDUmbJ76sLUfS3sRX9Ig
BJAOoSy64+ISOQsmXun84h+ekrjwJ8jSyjjVeImzLmKWCoyVSxq/GORnOBXn6GBO
dlN4s53EW2SlqPiyO4axbw4RmZgb48YqJ2E/a5cR9PMqthH4dQMcTpG7gM4DhxRQ
P8Bl253+gEEgUCRzn1q7FqB6P1hZ8a7+YhDN5vziTnq8yOvlA1l8PJhxWCrsiUdq
Eq2pzBQAbhMQmJcRAMOXe6EdnyaQTDDa+2BonjQoBtSb3pDuTni8Jgf6XDAFXKLo
yAAFy3V0WF83GLeCWOjvuUDUymv23k0/QHJ6fG/Ni7r5B6vdi7gtJXUcdlluJz/4
5IJfGs6fcIDI2swUiK8yy0bHh+z14R0X+rs8y/bP+oKiWaEmyd/tkapXyFxQNdrT
Vdw/QyMVxx8Cz2WIUVIvKrGXGhF0nqaD7krKt6v8kGhNPGdL12w0mtLXND/I9j3j
SHDgMtQrRBnCBxBBDAY6ty/Ty1IlMdIAceZasXMXUauLt27L8AAIe0fWYJ+5bstF
nFpGzLk8OAYr8JRQRUcZq/wqc+R9Qq0IZ8KPI4JnVsHi5/WtUbjlRRRNCy34mtNB
mWXC4fp+j5YzYkhCoHzaNfQHKiTBxpY61uKZ+7/2H6v98Qr49qNbzJfRw/AmWntU
vjaD0uL8bhdbopdrGd7hBMMdYlhx72gFe/AV3g7Imlaz5HRubBVtYhzVEegvdZFW
RoWUl8/7+AdEhBHvwPgvqFB3me1TTgGGpNVgMcbs3TW12st74k+xhCI6wvPaA9i5
BLAdwnpk6O7jPMjwuIrDmqF6azIs5y2dq2sI+xD1MjWFYalxEdaxjys/pvSrGUjp
ZsoDxJBJqu/qSX6h1qOvs5Vc8s6gBVPjrzqY2h0CQ7bXIsVat5L3xLoYXt52I6R+
CZv9op0tXHemXWghA7R1kda6h1MwYwa5zu8BIHEOgWL4R5W2MkqjcQKrimAiF9dR
55W+uhawb+m0BPQWx3/iMX6CCgfcbUsaWybkQKK3xcgM+zxV7sKR68n7d328GtKw
RjiRSMXgYvM34eLs/JJtQ6EAw6SauDgJ8ZMRGj6+mx+MQuE7DxTJ7yLsTHfZ6B3E
BqB4mp+VJX5cUsopK8e2/aiiTpwU2HGd/G/HSfzTVNhzjlVUX+GPX13nsAifBNjr
eH5VIu5yOyDJ2/iUp5w7WiQ8se+PO5Ki4CxZgAsZOfAL6HsojH5hgiEHfkShFup3
h7ek/IHLYF55z0xZELaJcxutekyKdlcjYAGP4+ptMKmEPI88P1CjPq2uKt5s2ju9
sm4i2KBsk1gogo4DYUlMT9/SRvLExbhT1zEE6O/IqI+ylGmmksBavqaOf7kE5DMi
Bbw9gAyNbEP8pLGnRrhj3BKgSIUzsrwrbQ4Qh5sJT423iGf36vDQ1M+HrIPoVq5i
Yu6ic5YcLplTm/ztrAw60Jarv6bWKBoCAD7FHDzdgBzT6HfUYUDweOwcDSYCrsoY
ESvfkuIVTW6qxFVWEHwQpfAYzbHdS7K+hfKpJAW/297caUFcfS31kwxiH2QVoSy7
KuyreXzGxEBgugmclbYM7L+TV3NZk/fULYq6JAOc/5eSdVX/QKdjRldAQRk2iKm+
h3J/RsXNIMSz0dY7vOaxVDyyZRdSwqRw1HdpRa3m91EZ6b14aTTGRqvKbWsgbG9w
JOrTBnz3L4qluR4BO7GSmiRdRmrptb+5dsGIP/9ldq4q7K0DRF3bxvPAG9dmep6h
CCA16sJTa/gOHFPwZdbWAEejFtmHByFK42mpyhohHeNnE8H2G79w0vhBoy5/R4Cv
vcHpxYTxkvHWOpmblXJc3gXmsaAjmFa2CTq2zwg1vdmuxIKwB7T5oeR/52gsYLbT
yOME8xHaBePOmJ64h0QwyIfIghw5GxLDHvOohOzxyYzyzVNUaPoqqH5f6GYcVmZe
Gpo3JrbxO0S+gIszFPWCicunmQFu26PD2K1PGdlu7OBHgRkelOwxF8S4aivbaTW3
Al+NCcpHy/Bj/VhhDore9JQOQce3zvVUyM1mAz0oamlZsy8HiyOLKL59qjbWo7Li
ottCTUQqGrudv51+d+oybmXdfmRYmj7O/aRuBkfa2nSvX4BwhPx4pwok1963O2V8
ABQqtcsRNruNbOOvHAAluU4M0KrTppTjKSpW/MaJwhMw10TWDjEOUw4gzMXZ75qD
vZJWAMyibDeuhL3uLLme91EnZ0U81x4YDOP0aLKq9NnkAGZ5tYDGwRiyNLhsOPNH
YxC0qUrjg0SX9c+8cDV1ynj1jyxUP0r2kIxf56S95dZ7sr2M/9Goz3ht2F40x4pb
vRATiAtaaw2c4+8vBzN7PMpaA1GdU52MDCvyOGe2wCIwotc714T66X5bIxs2BDP1
vtl94chBSIB/sDrKL+X7MaehddepJ2cSunTnDguLmw95f6YVzLMi+vm/ZLR9NwMD
t8HAncuSY3QIpk31OnDuIVQx3bsDTQcg0h1yjpREF/DcfgxhkCWKtTf88kZ2zJQM
FZi8ieovZDHvHBnzITRu5jM1fWfhkI4Jkp6sPpGolcXqd80vdS3iwzKVhl544DEq
H+g7wcSWVW/uu8af8E5pWp+sEsJ1Bk79owjM+QQl5WcSqK96XcRbH8EDTcSL3j0n
XVxVC5NA1eooAS+YOBHwNLb2IYV3o7w7VIMiH/y+TtBu3tvoaG3EDBr/JO7hzIoA
bfxWTwKgNf6K7KlGPBqRmpe+GtLPIsStBuCEY3nt5L9a3ozac0vuRzTkBYu255Xz
7+LwMjwJsuIhXUUt9lfIL0GAUSoJ5TQdkMfuwtHxfRBn52mk5KZW3zSWQLfVI0V3
Jd3uOrGEzHPoIqIKXViMr8rECw7en/df4DzzdLjGDxq9fpNH5DGOt6KoWcWIzIhV
C+37Podt6yjodxDDpLqXbKPIcdsbrKT0Rvnk1CqY2rZh7uy+XZeIX/qw9Amsj+NX
eD0ydhb0ICJQatOIGF+xUp8Sl+oW4OYXwDyzGC/EFlwIrKCBXM40aSJgi0hAKhXC
rluPbcPfGS+tVzssQ3QsLzKsAkIyKtlVszdLIlFV6KBZtYhc3rU8n1cg9gvnfcgI
n9ODZJ75KLPusg8nzE0B1jhYKcx9tPKTi2POaztpemqjfwOnZFRiHObit+Km8oHc
HQhxHkEj9ivKI7MAK21O6kDyr03a6R7ZiJHfDOushinfTU9kpqzIPXfGnNNUQSRN
28h7Hh9Jw7ffbW7PBgGkqv5gDya+NMmKS4N3Y+wkqCoLc65T/ggbEFwwwGn8CqQX
RAiWjVCMavIT8BsiKn84XTUR8uLB1Ln4SrtP//Y6RSMGsNFSvv86tGYU/3D9xaM9
RRi4rJ19gQd7nmNYDHGBQascNoGacLuGdu//ggOjkXqnNIIl6nFFDtiWkU0/BjRc
Jsh3Jho96NZZknM2T+TXJ+0Aol3BBsAQuTuJZxDZ1TDi451EMgeE7KVg9qEp84BM
AbFgkkKU9157BjYDjA8hIvC2oG/cFdtmzu0tW+dZG52NCpCfoVmAaMPqmkbwt/E4
Lqa1hn4T1kceRX3Nt2pw6pqlqO460HtgxdhnGoiwt3UGIEXZjefMt+ZjrnwY4YSo
yih/Ab3Momlee4wdSwf9pruXs4A6iYJ+UxtgN+KWUv4vbtG1YIy6p/ZcgZeFWBDG
nF+OPRf7m85nMu+kmpKO3O3Hod1MqUkgtENTyqcpVkdO0Z92kNzRREGYKOPsNsFB
PdsCCQclS1KAMf03//G80Ke1tP80lRI3uP99iwI5xZbdqQtVP8HWOFDBkxWON7bj
GHp8yVYxdu4huw7+qlWlHDOjJQ8OpxiQUq4nD3l4zd07ZZIDXv+QkCdxk2wK4E2i
G6R4fMSauXFpmlniPFw56VBGD+DjABf9dSGLGQg27iJtk3sMkXGtCStwyH4ZokYb
xcD057A4Juo1kNP2XFAZU1H9rJBNCxu/UgOG9OkE3oSca5UqxJ2xXH0ThHydzIoA
Va0RGyWqgZuqrAOLEZ2zg3O+KbsD8U7LJ+uJCH+gY1/2rzlBD65Qm470oMtPah34
G8lUfS4xODpcjyPLKsd/1Jzm9unwoYf0kHNEKnxWhK9ULV8L9nbxcxpg/1Lyn36P
HJeB9GnzT/tG+R7XvEubMNho4MtlEdaPZBdwCrOQEhPzQghaSP8eh6owNDawMP3q
CdTS6YriYtj1gksLjGcJVPyN9AqOB6ZjYWWGT9RqXunQOEnByJPCJQbYPHszhGdA
wh0wWVJgbsIXRcn/UsMEWlU/z8/nzmERa3/njvvW3aYNj9jDcTgJg0CF7UceDo5A
BZfBqgc/dre6clcBVGZkR4pNG/9yTc2OzGVKiIpLk4YCz0uwwaIe7npI91S/BHdc
MwFJqbzkgIhNLSI6hE8kyYN6kIoo5D93O2h4C9wwnj6kvmuLXmuoGfCpCd1pBMz2
fiCRYj/gPWKK//hD4eNpWR02C+QBqY8AM/yiegBsYKhoKHAOcy3DlP6LP/oO9h+3
kJnSo7s7DarO5KBnpNdK9uaUhUELswVi4Hc19iVpCE8jM73Qg1Mcg3ocgzlMMguA
az3/UsWMwMw8shD4qlL9Hlc9OXOnjUFWln5/8Sw5sK6nnxswHmf/NdwMruRJOfNb
JPc6JzkpRlVEg7ZvADcIVdzYU44qwiBnqyRSyUDGztgaZ8qY8NpEpffwovF4IUxd
fhmk/WoJRU5mpiFWExBd4DkLK/ahdjywZ9/UcOJgpbh8Zh6r6RW+82vwDGoBBT3Z
zo95Fis6mhTM5xi1abhJtivqwjjVw2RCE2Oy21x2JCjHH0qIQ1WXtxcGyG2Ei+1W
z01kUBhJwH/CGe+zbBGGkwdEyFxeS5/tRTKD7+WepFlm8d3KFXmOkCjLuIn8yDTn
GmLKILB+aXSMV/skU89T5kIR751bHMgVj8LRZNIwRcKHAzQRJAHeDcLzTk1EYh7c
jFQHjOYaz8JqKo6zHkWvhimsaXCDY2Tl5oAUIWGuRcCoEeE8Elncg4fnm2ZMpt3T
uQmlxjEQMK/j6T8OUih27Z6xRfx3UCvegZ0b3d7Vaw4kmt8dt+n0XHNac28Bzb50
KpZ01tS1FlezCCrjGZh6C9Otz/24JdBEoIDQVr0ULzH86ykOdFM85S1aaxPybjKW
tnWMjulZum9unu7ON5P+w4NRwm++vlZvzi27N7ifpFq5gZRWDRZiQhH+4h03l/UY
QL/+csqTPGRU/N0wcOaTw0C+IDzBCXLNQTyTjWtMMzNpftaf1VmjNNebeVjGZfAw
XQAiiVN/2XLUMUq80cRGxPXL4UWTb2mTecsanSNIb8MIjklfkJe+WT1Z3pVtRyqX
lm0I+iq+5glR23/jan99ZpY5DWne9NnHFBK8hAQOd3/AnbqFaIxC78/+viu5n5y0
zr7LdQcy5Una3tdE+rGjYsrQ1Vb/BZWWD/DGfFUYilPFYcOCSsof0YV8EsADGw2q
AYiv3VN9QBP8hyjoH3Mv/3VfDCBKOYkUmzO9csHh2TNj6szBX19VmbMia5sYzlaX
/4M19rKG13cxSar6rEoyVUTo6pU8mPUIdWd5Uqqg5KX7whj6NWeuliST00MFmYd1
1R9cRJWwoXFGMkG/Roe640/JnVa1yemhgCcLTvNC8rSoit29vGKT4Wqvle8wr8Ct
zNDvob3R6lhPMtoKkqjZjWUlndWby4ZET0PX5xaYjMlxw9cUaSzP+eaut81buWNp
Mr7xGzLKYGZIOs7pLXjkssPKvY2yNiyK/P67CcHYuOVNrjcxxH4wkvJpjgM9ncSm
1+HpGrwMuoY1zRs/IUwbffoYDqWqcqQboeduHEsLOHYM+V8lNzrM/OND0IN6C7gM
aMOs6kVkwdaJhS2rB7ggIYaS0A6JWNd+cFxC41f29ApKPPZSUe9ufExM5KXF48R5
w34sLfOr9rN06YxLfgk/DT8x2kyZjcFk0d3I3DfWyQUT5cGHnPMAvVpVUiIQVSmT
n3WC0ZVq+hz7Z3XLEq0pZ2JLX4fkgXcmGEkxsnq3gSJzaIS/f74xIVtwLqGz3VRY
FPL+ndrof8VHGW+gzmbyvgNEnsucUp5kQsjhFSqZDO9eZTDUtUWxfxTmkzIxr821
FHciepxStZgTj0RQ7MDlgONCw+K/wFpt9Fk3s2UGn6N9t88UaAVQq5JxKM0cLUtx
x4QKvij5LhYEUceaKvhttCgjqijS/FAL0AgkmHT0qvD3tbc9lk8dnpA1Gatn+i1w
CiSVh0Y4/EtE3s9yqzztyPVTn2b+MoQ7bPI+L5GgwA5oRZ14wHjVKRokvWbeilVk
9HFFz6u4tMmDd/vv+xptibNQnIofgtNOPVhxqkhbEV3WFu0Ku9j5TdUzvHDuxJ9b
oO3mPRjBcvl/xFZcq8/dr+y7UXjp/tMDEdTt2pAd9dcL2phrwruUGo257QcjUxrX
1PfoLPvIKPSzINL2fCSiYngt+7vZV/zjkzT6QqJtI/n3dyDbPNwqiRtU/GD3ARa2
rjz/62ECFqib6NmP+33lYmX3M8OXATVqNuw9Lwp03mCWd95cvQS+z/O4LcKKM2bH
T09NqKTkIsrdBmUhuifMbg2gEHXM7c3r4TFrOOMpGHfwUDyiOVacxU/mSbMtcUhN
moUQc3qkHc0FPpVSA5NdUv2BNgQ43yvevZmzdlIXEbyGaF91Feec4+VJvB/P6fsJ
hF0O4UeyDDPtR5mmQWmEHYCSlqt0TJzkuFlJXChEx2B16Np+yIx61L9LzLK4ng6r
iP4xkGEhGxUkHNJiQbWridYNxwosz24RQgCl/g/quY+k/v7RgqhLCQD2e/Mb/2ip
6Pr4m16s3tdbxlJaG01gJh4Z+qwNem1e5gVLtvxj3q798991wIdeeO2wQIuxPaqS
bO2Ccd9CwY1mElR0Vy8aapnzfJ51d5EL614I5mPndomXudTEIdh7B5lhMF4EY2y2
IEqnyIlJXrTpn8vMh4oScXKLKj9kPTaV+XnktW4E9ELNOAffHFdrwRuY5q74MBq1
PxZ8qsLV8gYoHFPX6qm4UZ2f2xDAXTooIqwdZ7wpFXiXkaRinOHZrN5MgX3ivJY4
58HxtEFQNjyUGr9B4xU6ps6T2ScXB3IMCq0xlbAOBcEyybKwXfeAL1p4p7eZGye6
kFiOFgTctDbUnemi3V37u896kyfwk4g1UXGdB5UydjdQSe7HbXpxiVkyjz3W148e
z6wa0+y8oaP1jsXpCQ6SqqSJRMG9pNpKVFzWpp3h5bwex4fTg8J+Hi0bko2nSRFw
3+n7w7rt7P3ScIcNlhXn0zpGGjJogyMgyrIlGcC/gx8lFagV5SgYymRUWAQA/lkl
DEXz5cZ9DwJDm/v9v4UEw8MUPoKqtadWt0m1Q/xLrG2tOG1BNLB6kRFxzi5WsHRA
dc10aTGx+x20qcm7CCMdDZnLSnG4PqMFIYT7sLnXhWybUIHzRJtg7ycWqRVoLsni
qDMoFIjOfRh5z2g7sR+U8anUUCGMWocNv9go0Bu6Kg58gHREdQh6B3KRokpl+zrk
r+Oqu3CCM816LKQP2OQJ19y/8sij03G0wB8ABQtL71/ECv8tWaxI68g1I+U5CAF3
7rnOUZiajUQ+q1AbGyv5r90G//dzQDQz2/fnQDHw2TrIWe8jYRJVao0oDkiU95Pw
5Xhk4By32rIGip2n2U7E0MlF0WJsJ+NL4Wboy7zRkQUTmzJV6MYJRSoBtlqFnhag
LGSDAXrF+IRfRzgqY8V0h8YUx92gL8Qvs3lU6Lq63W9iNueWdg4KbaKIKErd6V7T
OxlHP7qS7IilkHnnl7U5HQgQoNm486gUdV7/ei12xBFOvS6M/hCXKYKNPAFSd0H2
Tb3syriI8loYdlmLSRcNx2nYafnPvUEEjDq3WET7gmBleJQl8Ql0sWN0YGytX/NQ
4NyXlb/wxlUU/PFDZ4e+UgVcUXDNWddnN5z4tH3F2cmVvR3y3cqXsFwHl2zfNQ0v
lilwr6qprNfhAEmJB/QNXhvCf/lv1WArRhDASAFyRgS6X6BmuQCOSm5oc/vED5GX
ftiQu6jhsM2z3SIjxqw4VV5OW5SbK3pdcx/27tBZorxCySDU8ApQ7bwA9UlS+Wvz
SuiBLDFMda10zadM0DO1AloTnB7Wls0nEPiOQzdp2h5nFm13xgDr+QnD8tY2xrM+
OaAxtBQI3XeGHNTEb1ZvRqbx6tqcfszVPTVC00FYrgfXPuOBaCLdp18l3QbmsFaP
xQGYKfCEEpF3Vvi6s2CV45YvvsBDXKD9NF+E4Zq7rt+0hbyXydgwZcTPU3j5XjcU
+Y7oqFXf0lTYboRXLMHFCi0TZWFBhbeRUmO1wqZC66eIaxtINimeAV005WXS94li
utmzLVLYXnY8R/96SGQwhEaZDz6bXQ9lS1Bc4mE0d6TbIf5FY+bZFpXIjmqMKhUn
NU77nhb60JlZW0PXPke2OTIyNYs8oMZkK37v9hXNSUAeA5kkwcrkHJ7cjeAgY0aw
tPsVsi3OdFp3OiOh/wvsAkX3T2naHg9WJwiwY2QSmMoqb20QNqysmIm3j9I0kYPD
7x0FFHErUZf3h6GTrhRlBqtdLZlF25GAjLVLk28XsY2O3nVUielXlWvJhN7y/HNz
wZbOe/f21XnI52MNCIUPzUVdvlLlRFmjfkDZWIQY7gIjbPt9HjOhRCDsYpodLveB
kIFdDTP++iBqKFlcAF2VVKrj7cNX7hyECe5J1st2FG79WpKk5kkTgGxDGzlggsLc
5sNyzSnxVkdLNOrCqDsqI52Elx1cV3CL1GqObyhjwnGUnZLb4o3QOLaHmtd4RpL8
tIzrHcNr1/aJ3jMD6rzzEBfJwnoX4U3azlv42otK2ucA70/u676EoZ6POkFpjEOc
bpWtQyDQDfTPR6BKKM34pZDSZNp3PTCqxYvHoQw6EfiO5uKNy0sOL7ztnQ+3adoZ
7L5BsBnOxElRzF/w//2s7y4gP9KyVEmvwAsRiVQNIlfsADt2B/U1ZqJ4umUbz5SN
Bcd3BUI/GsleUMHdGWaw16ogaZ4FIJOJ8ch3TSks3NslITsYV2NosvPAh7Djtc13
mCI9Rsu8+IaNW87R7YPmplxT39Who8agQ/OomdDvLWfxrQ9X117S+bbjYMlKS2bc
gnbseraftxaEHpHzhaEJ7c4wr2HwXvck2/rPW8TXGAXAzb5UpflW3VaGu9FJuqeh
GNY50ib3YHdC5fgr7H8WJS91BIxQBAsNvnKR0R9LhuricPq53DOZ8tDV8Efw/5VU
gqG/4QWbYGaLnhNHbwetyzpikp8NEGhuJa48GNbK5xFL9AnlhGoQTpR7t0pJCGJY
09qH4nnQFqis/bTWt/FNPl+01YPFvkJJolJFtuwpCte8UEW0qRrba9IOIzPTbhSI
XvChgvXVaxf4uiUItW+lkfzCrJiUQDJqnx29gdHX9cfyQGq2ernvDaFdMvtyOMpN
T3MKVK/mZGGXaEscn2GM4RsKto462vHS8qvbknP6NW3afUTXBsAYCH7R00XPRFnO
LskGQk/CcBd8bFRRSmusrLaWpM+x3mfMY4DafGHmnM0bVniyuCHn1VAa6PW3hb3j
WrUSKy3Al2nQRrzJuENL1mZsIWPc5cE+quv+2tNAkhhxze2KkKXp/Dg1jxY5ord2
vMUScARR8wjJX9sZcSeFLRmF6pFt7gODs0r07Jph2mme/8mZQEYIUf+UKoSoKr0x
lU4yAH2qhmjazbWKvkM9v1j329AzdVmplYlTlwt1JQt5ONox3wQwP8bV1jTIrBfw
J/r6Elk3iXXX5+ahuPMGE6V5PCF4aNYxESDYDMdsqqlrS6QFsRd9KntEgZVxhRPF
NWknxooRSVu/QtIolCdYeF9zsBpT7T86q4lHwEpOgTArH3pk3QxN1MO3LiBU4UJJ
Tg0TyQ15x5t5VME0uQD8ilVnRRP1rumE+ORK65uAJezigBNNnuUL1xwrAJw6b/E3
o/haXaJXafnXg2xu5sXFIDqGTOCcUFP9SZxjrjRa+pHu+F7jbZZZQhlN9j+Kw3g8
AfjyqPLuJkBh2wcJrq1nKIViSFSK6mKPLD3jwvdKYY15jSjTh3bbm/Z0eRx6uTJG
W6OhqVM4zMo4s0fYVa4uCy9AUNl/9R39tTIv2/qZcqxRwapMVDGckCbg1YB6LUfT
M/pRoCEG7EqNpKdTgEvXigqwjZe3fA5bYi0q9KjTyOqfNasqJhNWf/qC0E4Hnqk7
Mz7n/YJ+NS9eANWdaDCX9jDfIUm80RcNOMkRuJfBZWaUVPIl9u5tNj/+qKdvuIjk
L5f/wGzcKyrkQW8oJDoBO1xHYzAv5PTOaup+dYsWUVJt3jaTjrOsSoxDKdSEmoGN
PjtP8RPskRX1POWHbyqN4xhdLGl/NScpDkJ97GH1f5HbRK3IESeAKjYCQRlWjE7l
K1vL/8s8wv9sBy+3s0iPhv/SMXXMRWde9s5eZhCojDKifS2AQRplTLCsey1Qt751
JbqzBeAOJ4yLIz6G5sb6JUBx9GXEmzbeJ0OBh6WY/13VzmsBoqX1BLrlRLF/TGl/
rLjWNFOAymRbHCLZtVaIO5TBFW82a81TLrofpSe74n2xhSKiH/iaxVxSjQcFEluB
4x97pXeo4uyGHHhfGoynSrbkDB8k6no6JFAFOvLEofPfyi288cHbac9LaIT8DL1r
rJ0l8TFfWvYJKWsDz9RHURBvHh+25pltLd7lRpaoYvLuQ1LePYcFSI2UKypmMv3d
mfqQ9ttZy96aQnketVT6ypTdEQibRLdb/Qsx8SkvUp4I92mHl750Tt8pvHyqFrrm
vtkYQy4zfYRjQnQcRwCcVDZq3flmpXO4leP5/2rLOTnj4yUyJ3IzoomxJhgwOS1h
Pys9pDbvKWf2wyb2U7MxFEnrPlbpH8R7v67PU/9+vrAb8jNLSH9Gxp5KN3h5MF7j
kUxgx730g8jRRTHmUXfpaM3f8HLdQxnOlS7F18I8KCCYD5Yt6jO01fw35CwGBvaE
jygk6tc9+BXzJMXw/ff8dE+71sAzzJmTiVbJjOKYctsas66zKPbQECyXkcUMq9Mx
/a+LUI9KEixSxK7whOmJAZsbhq/6g6bRivpv4HODTpaA7AQebrXi4fKK8NDqhvg9
2qLi0hYWqBpdxC71woRbGWsTpN/RkJMxc0OeqcoX9EGg3Qk6mn8F8exv2RNepAiX
SBJSwx0QbXa+TpqiNLlECx2t8wwBE76PoWnyG6zlj1AisBdfmaeinvyWtUEhBLyd
dH1z/42y/PTPo5O54J1mlb+XxtOll/zeMA9s7IPFxVYx3Rc3oMBHSrGWrirGLzIX
DyoxICBzGxU0+daJFLKR1X35bCS6R8T6LV5tHKnrfe9hbMllzGbE1N2YLQrBhgO5
NuHeXFNqiIX84bvteksmP+dntkS/U3sKXT8rHtkw7T7wqKcBpOIBfXfYff6ix+rn
prhkg3O4OFFe3VNj0rtrgEO1fR2K9IXaoqSa+LJl8PUm9zFrn4gDXG2Om2j4W2D+
lF2povBuV4eAAXhJVcKrJCB2O3FLFQc4BD+GJcTfYMo4UXIKhDQVAri/PhDDqGlU
G18Wq1MV8+1plupBKrMdCTGVIWdaD4mqb/rk6XeHcNjBonjWjYIXffSh+PIcYOJT
Bbf3/Z7aKl1wSGv0NDbGCbjGEhkcCwDKWVifb0p1Gdh84PcNMVjp6h7tpkQfo7YY
v6SKoYfzPbldDRKUTHveJFCLYPIfle5rkktWsZzf0h2ndDB4rCs3pZmg7HwTNYFN
BmibjMvqlg1+BabwOJW0r/X3O8J4LBQ/Kb6CBgWgOKF2XquAHSmSaxikZIS1HwNH
D3RtmuXpS9y0zaJlIsNqk8O3GEz27BjAARa7WmYyxq0GaCBizB8yrbRsx9y0S8o9
Ne9VH2/7zdMGnvhEaEFl1a0SF1rGA9RNAQvGmRJDOFbu24/iF3qFGjplmsE02fru
4jHRrBnwZHoQyw7Pg/3lI5JRssRevFcttGxui6HaB8vjBNkBKlASj9veqWomMd3L
/VKiyD4yT3TCe/0VUopPXQCFHgmk3UXOjvQ4GvLrDtcuFk5eaBlCXDsvZRKDDmZ6
wFDf4H0wdVQl2oJn3FXWqeiKvWDF2y0ThH6E1jxI9mxN7/uSdQ9rRcTFGZuC9N1P
jLLrN484VjymMaBDqzzwSzKOSPkEsEgOJMPvBteJur9Aupzo3SyuIsrIbC06zn9l
TtOIMJb2Tz2qZ4SRKAbC5y68mm+btWarNzbP11AFRJmwyv+Spxeitz4Fkju9wJg0
Z4O+EEX4ynrXBO5omPzPhKJ0QHeTBnKFlbCYABDBuG0EH9iGHEoIe+VG+q6XLS/n
BMBOC8dnhc46yLUt5aZ8jqau/lYmzIvXysWceDfIj958wtPfrjYzMr9Xeyzp6/oy
hgAuNsh92WxYUbdTjkMGs3qfV3ftEItEkYqaFHZmWVLdCju4Q4rqnMTdC0aWisF4
FbIrkrN7djn0zrWrJvDuPRDmWf/2xMbZjl7wNilppICx5yICRj3nB0vpSJJD9fj7
+G3bn9zN4anPlJtdyws3XqXhTIm68ohlCekm44iaVd6f7ZvG6Z/2QgPk51hXuYj8
GTws+5TYUwpGqCIuwysVNTftTf3tr1njnRHY9n3A3aaZiFPHrbtLC4elggxocGEH
AK7+a0QkE5ZgwD6+zp0lKuGZHtxiYx0639W/G63bRy/bX93uN7U3myT7+YbCI3fN
j/+tve547z5wGQvfdoph0mPWGQFubpnm81FF1KE73T8bzcF/GyKfD9ptTGh1Aqk7
r2a6xcvXNBfIllCozgdFxuCp1q7i5RA5L0zbrVDPmiVuPLN+gvbbCaxCNsh+dvhc
me8qHSGCDmtNumDgCx2d8mE10CDvhcQ38Vaw3EssXlNpQ2dOf2f4LsF1pJR7sqr+
t1yuKNBs23xh6EDvYUMmM2Lwu8sDDHDrZYJXyLSNoczUos7hcRMoaduqPEBOs/zl
PEaSBEKsuhZjshzYTCc/L7FWsojGvYINlXpgs+PG5ecBgB0eyjmWOQxVWDZg/7bJ
6A0LC80eVTcElwt59W2KHodaJvRXRwqfE+BgBCH8aRwByAp93GZ4aAbiYLYqfQrS
pHigeYBJNV4ujRUg4IXqvbi8a8YQwYERN0YTZBPbmX716oBpjzT0Fhn5mSWTl5Ao
MJU+AGTYZY4zUX97KjEYTt7Z1bUGyrMJBhSYTB5eVTSqstTgMt6AVJKooTosnaxJ
lawRNL2mdsRin5tjXLEMZs2HwKmjPBCUiNDmxrULSoQTLghjC66Ut9jRQRipmafV
kdvgsQqwkcGeunyaQtYRtVhVYXDyDjDYUkWslvTtPyMO4XAkGqRqtSb3UlLnpD4S
n2vsxL8F6/ktZ92JMWgQxBnTvG8FIvVlEwkN/VbGP5AO0KorW2IOkKhXpDTDhOze
eoJ6umrdT7iIRr1AMke3HHPLOexuuUE88JyrBv3nJw2LaQD2ztw3mnBFpvGsV3id
pJQE6M3hq9pyKRA2/W7E/77FUb+mb33zKb8Wo/VJ4b7YygETIDxr04fF6IIvWnVm
T0uAY3JalaCJtzV3yZirX7a9wi4MHMrdHOQKE+r61StxrU7iiGm29ey7kRsM2xz2
2Lqx/DisRj5bWfDVKPPzQdM7oUYP6Fgf8G/2vuIiYJ1eS8VeARi7OXs8pqHUr4gS
sC3Y2eOiv1TU68Nh82GsfOA3D3PSjrn585PUWlJMEKMwzg0Uu0667NuN0tPhDSCc
3ihSxDV8MCfDzYZ66LLR8mihRn2534Cg9IL2dJaoX0t4inkUMxAJYN4t76y3ANLz
Dv1oNdwe4hJpEGeaPxOurUEb2/nm3uZ3qlxT9larjCpi2ymdM7xGzjkWCx2lwFmV
AsCSQMEKOapzWobkido6fZV1CPhcTBI4QfzD1Bk65fc11EFHW2gIL/Zc1LVRFQ6V
TGXUrzCzgIXt9vhEZ23ykesZcDfckDdnTn5iQV/IagNmMjKMm3nvL+Wu9Xj6WBJn
m4cLj0ebPbaLcxuoazSxfb+VHjzdToyIY7nGeKU/l1Ex+WOoR0MpIRsM4u9XcZ/F
OMPdZC31g5YT9TO9rz8NASr8vV/ns6XIhWedFjrwhOU8697zv6jpo8xoHeCJTx+I
0Z7/poFaBNVtkicL+zYLrS4CtDhZ/I69IeBKouEnlaz+6dzN5QtGpyN/pxVL+l8B
pKKnNzwyco6/eIubMo4gTdW9AWMpIJicMpTedxSO8ffnVsHrwrKzLK8lMagxIn3a
nlL0NDp0XwxKT+x6tEGyC0nd0BeU1tiqlhbv2CJy/MQ7LM8XGBOxpns3unqfM48V
yhpCKWHy3+ahb4vECkPvwU+s+dWkec5RO9T2XySEJre/8eGa4exyEdPPF0i4ACQy
KiRkwdV/0iQnCyTiNn/MBjPzEbPLEszLNdhP51dMKKCmpGntg/A1dq1kc7af7zAk
0L9Dn/1uKjYRqB44I3yCMIi9BPDd9MpJ1XmfrjmXQodbhuVrp8rajAuEDKwGcjex
ZBDWe92d76GmSoPWNuaHBrqM9CccW3WCN1rdfu8q4aRCycnPzzhhZ+8wVHi/qQ3K
001T5QHQTzEkXHZu3wfrNIA8bBc7EqU9sWTPF7gF9LLLHARHgDIeJ+jPm2dFJfoY
n1eL9Gzvn7H8zynk+XyH0hJPt8VhsOEM6RQ9H6aProDuz6+11BPUWLAJ+zDHoYtW
vY8HjOfJYUkdU36cDrXNtLmoTLI2b0W1QwZ4lVC31yu0V37iDGyDeE6YwEE693eD
wvEF659goc08bwgGks4riDTALHaJAbtPW/e8lr624Ip9R9QLuogkW7YMbjte8IL+
pmbKNUKMWoYEmxM/KasdM4spa/XCFgxtCHowq1oAzc6l7akTnmKXDMZDVzuX+Le/
t5jpYpt6JRNynUgPfznOJhdhVFCNrFJZihQxvA62hHpK3shnrZLpO1dCcZ1udP3h
7IXgqua1TFo0UoqeBMsCy/PI8Nay4foKUGeU4b3CNIzswWndjTG+xRk+EWSjrYGR
a3nfJCAZzNfh6sVH/Yd1yI19MR9V65qJ/5iAE24QO2JrLZsfupXD5DbPgCo3lP0M
rizrJebs+qFUx3Wc5LWZWOnU4HZgcRezT3jZPoIjWGXzq9wxGaCKADTEwIgw+ydO
QsWWfauMpE0kIv6CxZfuucumkZxO2yzW7ocEP7G9l9iv7W+cc0Bkkc3X9yclsB4z
r8LVlFCwOtP5PVpKjcCy0RiudllhPuz42wDzeCzO1SPehqqN3kKeqxREzCP9eP7Z
mJ10A3j+qgPIY4fMsSqjmMcK97V3AMBuWtEAqUw4Tb8ays98TPC31Aw9I2cRDdJb
goRtu+rKFj+37WHq6GdgpF2Ng7t0vG2xdc8Ef9vt5WVIwG3H0WC6HNwdxo/6oWbY
SLjuP1LH7K7nn6V5AWbzZnY9tMsvWTRRpHS7YWUHTh3lw3As6a7DyV0krmhXUykp
O1zyO0GeXokf91A5NgPqT3Q+2VpXQm0hl8pCd2IexQTRXHJu7WRNfM79lZM2YlFQ
JnBNpl1gIHmRiOikt6xAYrpTpSMfY0zpS431+KDDI4UNkyErFE+egpSV4Tvfmrhn
YBkLV+kwwB4o5sC1aGQXqqPq7b20QNd7aeg7kF/DZZTLUp5Vha2UTxhLFbMcAo5A
qIhVrQjajYfUgK/hemT1lyjYlIARCOEyQWEgVEcPpp0OBaemz4nzMkQmBsVQftKp
312HXA+7cuIMR5fVCkeROzsNohvUFtES/yDZKuWfTanwhL7YPQj3A12A8JzfwJ8h
ojh8cH6CLf3Y1qEVjsOBiULAo1Sppd61wQ7sSvFciM8npuMZGpsdYLnrSed6W6ov
AaywjfewOWVb1XXQWyBr3x6WDyk1vOSHhagpYbw9Dnn4YVHkrDFo0DY0oBzM4Rom
PtZbmM+lF9ec2rJQGpmJdb9MkQvBogCrc75h6Zccr4J2tu+8CvUTicjv7BOz7k0K
vFCi+s238uzg0bG7wBaAcsbq2i3UsnK/vXrTV3XR/yMYXVvTAX/d6HXiaRoTdR4l
DjP4pdoKsr5dNHj/Bwt/E1RPb6IVOXA8oIJhv1xs9MMD3kAH3aGCFO9c/CLwk7te
I0oEqe1nZ+F31Ni5ExrRhH6ZBcKxeWAfPXG7OrSmB7bmpRbykA3J5DaXtl7Jyz06
Rn6ZtQCaXCdrOwQiw8AkbKY/oDI44m5/3nW6sP/bbSurwjg7KEv/H8EllXXfjc4m
7fzKO3xQk8t649KkfNO257JQ9QTcjqFk7bum9GeJu6nqLseUIeIOBykDdWx7Xl8V
2k6hij0p7YwATqBt9TSf+JKAMcvujlgAH8bylS/NWGx3AnOLk1JbPTlGYROuLg20
IoxQ/Sp+gRcW9q/shnDRDW+AceZEpiJAO02jqPamhTjzSzgTnfR+6AZGjVxc2num
DaslMM6GbgF0yxyrnf8OZYfM1GNr52hfwFTu+xXXJ0WZA5kH0JtW7npulFNpOCDa
oaDhwh1/TRwIGggFMwQDCKZkLMOmJXSonzN2KD/MIW6EXiLWF3LSo0jG+enrl/Er
i3nghV1HpxgFAS9uMTCIjwB+/olpWDxG2HSVm36xj67T8KRs6JTa4mMbUAGrkrpO
FkIvpgb2IYhcl3EAYw15LkscGL3VWzrLPrbMNksakczJs2kWkKlHaXm3oT+xKFXg
pb40DGYwQRia9YBPpcyZUxV4AA5TtPj951DiGSDV9vyCNPNfIT/CCxTED4XcFJal
hQW1pb5Ldw/MLEs3eUa2FDT5ACe3OlM9pv/qm3vnZxls6OH2mZHqewN9SjBZ3B4v
8L1/CKPm/HEnw14ltp7YypmQX4tLIMgwFaoguZmxhI8IeXcpRtEoDiirjadmXotC
fVYOpYw9BmldXcWAJIKCzTCRDlsQEiT31G1o1B8OL3ay8u8NSqW7a8PnAxZXmw+Y
L0+BcUqmUE5KgixxoINuUGamwfHPg50xsxTmpkvQMmHUplBHcy+/8Xuq2iFWu06O
QW0bqR+YPoWF131ndo4YVe0GrTa3fY9eJsYcJ1bVAh+DfKU58CA3fwJ50gdXBICk
kyYR5E+m4hlrpIcTeKT26+Xn6ddcgwL8KenQfqamlPT4eaGiHfVGxVv+OE75TWIh
yt97MbWrITZT/MplrnYxmdDpAKdXIFAmK/LUv9qXZNmuJanmvnEv5uVIvdwLrYe1
OhCkd0up2Yn1RAGvvG6NT6vyu6eQ2GmuDgC7U+K0LvadF+LtG5F9QOcG41vn0zYK
YQpqdrrvshohZGjLzkp5dOgx+00SYDag/m6zPpWNOPN/qQupzlzrx6rKVxJrzg8C
CsZZn0zNNUTS/pM60rUyUKu/1GpDDtCfvaIA1nkac/9EvkomqUTaX9s+/Z0Wb455
/FtGS4LdNXaNLaIrtqSvjCZvbGO5nPS6s1PA3a62s/Kj6mOiTA8/nr0KxzahrZMn
I8HApFwsSesqBc28p8WMF4bSBIymGr4wRAOsfU5cffw+PBLKNOFu+gzYXUAP6D0I
/LGXxkD5mG3JP74AKuBD3BvvIwkywbVNpgwf0BESTf21xfaGrNVok36rvv/4IFVY
BkMxBTxw0wjaIkICtmv0Qm5V1FUxjPT35CVTuNIuNs8t5sWoKS320RSU8Hw9219V
EVDDnnxQSO57LArILHsFjaV8cEGChw44J1jLzYYjs7jV0wAuTCE7BSi1KyRVALwV
QZKm7WsrxsWkyrjx74xxO4Za2fQLrU3HxchGfR91dVdG3g0wE+VMTranpeuaF+SE
03iQmKccHF0+qxENbHwfK+2380TxdZ2eo4UDb5HKs/AMbDPqevXyfdcUbxF/eDz3
RaVo5eYGy43T5si9zu+ngad93u9lWl+5IDGLaFJgOVPHFAT0a/hCpdDnEPZFGxl8
7f3dldSDWpH2uzAYI09WScPbPxbckAhqOX9WdAtNMTt6uLDVhSRLltC3iL6Ueq8v
rr0peZlSQ4acZILCBJMyx1Hl7C19WfyY8bocOk4l5MkkJ16JCT/76XD5GImD9U+r
zhKIjbE8V3Yk3q2VaNgnyna7CgelNb+m9MAvWMXesGtkuKNP6kph510lIKiueL5U
uxTPpOIXTGXWHjhLxg2kwutDL/0klJajtBTvmMP24VoWDpI3OzXAgwYO9xuCreqy
sB1Vd7tWnOJhZ8ssGG+IOG7b+kpcZytziziVTHTIfWF8BPtNBn6L7wKt0emyCfF+
vsaVIXuCqNhMh0Vfu+7atrw79ba6mCnT1fVIiikaXlg1yLMZsCsgbSGsYMxCMuMN
CcEueAl0xqMUfSVWCXDRxETQ0+lhfFsqkmklNJpxWohmbXJW6TC9AogP/YSMAmmB
mpsAzCxhSC0+Mj0IeH2JW5ueNEXy+k+LA2ooBUdKS06mOJkBJ49tMn8EeanjzKsh
Q3Gn2Y0fnh5Xq1Vmy/OS4gnBW8FCW+z3yY41aManplC/KZziqd7W87FjuI0v7HUV
eBGsNysLE7erMCfVcpFRAgLNiQs93cPeJDuYesKs+ou04ivAEvcXOdEqFB9Hk6sl
Wxr/BHi0BH7bbimZxXw/hebXT1J7wXqzzE0mI6wM8mQk/oVLCoKHPRJ/bOsBJPlM
WTrLY71Qb9hFN7sXgTg1dfiOVmb6lDp1HW7BztL6Mo65iXe3Au5zAIWjqlQ1y6Tw
PNvxsJMtK825g6zB9xXT0VYnI6oKv/vn0/IuXwJ9DNKSNKNIYyapeshH6cqskQsT
VUtgzay9j3KW2hynPtOEozXqub2E5j5wgkE/D9gzICCi1KAGtVLKRJPa9GhDB4cJ
o46zJWDFSaXF7AFN8ixj2VNX4qcKLnUNm9Xqi7cfTWJjngwwk9tkaUog7niCuxU3
CojjhpSknd3SHvgpmH1Jrwo4hbFF7JalMpEfb3DbKIh8loZGGn+gcZvONKEvzstb
Mgh2i/upouaP/eQVjgoCGaOpAjXUfsbQJn8+0396q8F/pBuBe3zcK/mY0QBIlRcB
TUr9eT+UZBCHxHpa6DKDAnufoVZkIT/UCLIXJzNNvxRtPzlKWKZIXB4GFipnyuUs
BWZSHatciNgG2BfyrpZ93pc5h9+geQYeeI/G1ZdATF9+BHetlxLA/oZE4C7sHcg7
f120SICfZpcJPLAd/3Qd8kPRKUox3FecevF4Z7p+/KerMgT9ctCl21PC52+tdXXc
tCgID+wP2I3g3ECMW9TTzLwrQteDeGx7pbH2h4z+HX43FViOlK8C1/oZUVeR/4Yc
guvbsMHrBc5n/MlU3zx0yOa3zdYrIT+fGOK3R3+p0jKjQ1hZMcQWZFzBMQ6of+0A
ytP921tdxwWqRQc6qi+2Fsl0fvIGGM/e7BK6BDfXq5fA5KsKWfM4vK/YvB7LRMkS
Vlncy+YMZqHK3j9lkmfWefWu6nvGeWFSYRqZuriWq2pMeQxMrC6QNdCx+mTIec8P
WKEbxlznCAGBOJLJQ/Th6befxDFCOdtjwX6CD3w+TIa4S/os1uZpNOpTBp+d6Eve
W7iHnPW+sjQ9D+JUQnxVwcRvicQCl5NfaceHbkyQYXmBnLvY2SSalzC13XCCU5Zz
6Q66tM9DOQeSMo14kJldNSoCZUMPnu9eUZmgieOpmiFZ/AhwiVkyfjrnftGMdLB3
jypYx+d/P6wXeWc2HZLZANDMJhguR2NOL20kFJHCR0gj7R49PUO65EJbwBzkicUq
ABcfCozC7oJ0wvCR07Ktc6u3bjieUKoYHAd50STcaVjt/yC4ueEUFwkcVdJehXD3
jNnU6SSK4ncXPFjqdTb7yvbA82jtLY3lh0xCA1dL1AZqKkg/2Yyq7q8FkaUn6j60
2dW80Tf9PZrW00fTQbra99vhO6Fy0HoFoZ9gfip0WKrr7xdbh/9Hpcc0c77+cL6e
peKAD0hcdi7N5iJkTNrHH8Y3dwsGfeNiG+t/6JVkkqZLtsevWZ50s4lhhTes8twW
HxfR2WipSI0dVWSNZBTEyQYu8SeTXqp6ETl3hLtfrw4M2vg5PCo86tkFj4zPS9uo
+aZFJCQMjvTtui0B9T59G2Ex9vLOqgncJdnaYjU+xksneobd5fpbLJZyD+rTPDMn
2twAqhDnbYQtZvjG3LazxZKkQYeHAbJS4ephJpBdhTR6CqAk7Acx7iSA04fbeZdE
cmxcv9YYL2KLjjo/Htjhg605eMV62XdnYvXiZoBqSsuMXvnCI1MKyQc5bIwZg+m2
aICI6+IrPFgCKf3A4GuHIaEcweCPVyY8XeIwp88Bf3GQTUJ6gqGSyvpM7nnfjRb/
zATqpsQHrvECLBGl9UAjabbqRS28XJX5/AYBv320NkGkwVEhOa7B17Onyepfcb+W
cpx5aSBy91t3RgyTsYBE/s32Y/jle7ZLjk8YE4+SBi9CAD6juWqbG4mbAbd0RiJM
2HmSxUtD5hhpflo9+1bEmdxhQ73L/axiHpFVagIcNoSz2DihbslkdTiGX19BsF++
geT4mxNsjtKgvrG0Nes3mMNY+99aPRuR+EiGLKXAHjmN8gInVlJ3qg8blGf/or+U
vE24s209JRVyrwSTaaAT+DAmGAQNWEjPakurZxInJOz+zZWbKoj4IYkbJ9eLVCRl
H22zt73Zwiqpi+qRXDL/A7J4+1LGO5v7pQdX65vTMMOl5IWTu/clHK3Gx6HCwv2C
rQq3tdXFV+lef5FHEiCrUtgAJdT4gnWCXKz62Dulbo1s/KEjuG2zccmijE5YziO7
WYziWxzGkRQID123+0DVOe1JMcuHoToX339EqXB5aVeXYWY5lPk5/DWFEKkflNiS
sGdo7fgyUEc+LpVdQXdfderD4HsEBiHYohA/QS6lTT+L0s6G0OjjdTMAYhb1xFRo
dqQ0ZDYi9IXNn93Otg+KXMT5YCkVJ+L4TmIGte3G84r0MUgV1JzUqBv8+/Q2x7yw
aSBbZjpRpqNkOsldxLai5yThroDXtBlO0UCaRAQ1ezujW60ngEqd6t0HwaT5SeDS
T+yX34iu23kJSnuGMxqapV2pavLbsQEpdCL4sTJhT1/hkpcnpO+PFc9Wkepz5T6v
gjM1ldwGeJ5hJxrHedi0JZTiCFkVcZ9noaSj92PFIqcyA7J2m3qMScJ6Lm+BwGxd
qt1qOy+Fjg44ZQTnILzvpSswqMwZQHzLNT34xcQo5LFJ9hAV4pdy83JjxKxXsEJY
xR4lHmJW0MZJzf1UJAvUsLw9rs35Knadfvt4YnBPfhO9Q7knMq7dqwXe7asNJZt/
xPR66UhcIc0DPfBp89U1szYi0x9yTf8pO7Jp+8zIwCmj131pEo+3ER8Uh9isDin6
RP50oe+VnSNyw8iaBu/PRTcic5zqTjQSbD1P8qYYojx1HIJm0fyleTmnN+eA0dbF
dH9tbStd22gakEl2zGgqwFFKjYRjfVo2UEooVf2Hz7Rbff21hrAZdofnYdkjNszK
Mp34KLvl9JoSXACfNAPdnQdfWJy+EP6TFqq5r5eCTkBFD8qCXNIVyucf+yPz9ryg
pWP5ncY0xubvKUy7pTh1fwzv2Bdc5oz7wQpj01GhT854o679URqQG49axdQRWZ3l
6tqwAE7m1mHevz2MRQFhXeelwkCH8FnKOhvcjVtGYjE6PoAq4uXQ9sCuNRkpZvXw
LBqDDcwu9UX9z6o3uGJNarle1iD92R7ndyXKzLjH7Q1uvBDNYro1UFInOFssRgqP
p8KK/2FEKjy+ZAZa+tBPvvZKUni0EB+JAOMNj1IC6h8cUu8Zp5Her3fasvW2Y1QO
SYOtXGy6PT6CzH46ffEb5aYU2i6bntQqiXpeminVDsuvBQkJvCbUrt0Qj4GyIaXF
JI1GtE6chFm0nVcxaUNr4bOSOkzoykP+eQE25jCg3jmhjHAVOpKCPLfYvCl2NXtV
yrvlUrMLe60CZc592DpN/MhZAeNfuINbd4/+PRWxsTbxyX4kUq52715BDplP/KSr
JOoRlWREdXpy2Klkh8+LUWAxWaqfMmpjAecPXzYYr+ebzW2W35ZcX42sKIhx1eOe
NQV9NsYQoSK8aux0Q8L5j1n6uOsrJOpGsEHCzKFz1YFji/hjsolop6oe3e/D0NbG
y4YhEyO94wjQ7sKbuuH9mSKnae3W+YNgSSCWeOCm7NTiHqChsYNYZn9WmBr/eQsT
tSs4kWV8hxvziU36fT4dWbi1zvOOHXsJzs+beKECDqueh5mtPxlRZ+EiIxHCzsbF
frehAssZUj0k0zKAIji1W4fDNM5dVH+5ORn34IpqeeexyAMDUYIF4HQOSeuayRdi
k1KZQ3RXEVx87/TJawvX31hx9XR8WhpkQ+pfPzpVlQe7ixGGtZoyenISD6QSJS0W
v88oI2Gj3gjLoQAbl23cWRPPlrGV4HrCC3xC2mbjx6M9HH8X6P21ioCE51ImQZjl
lWt9SWaWIYYk1wQRDKzlnZ1Znkf9lA6LUS/XvRq4wQxXGe2Wud2H5JhlvOyjbevM
cd7Xlui/eIqtywDGSBwD8pfCOwUHh51us44ipihGYnUPMnvy2mNNGoguoyMSlmP3
RkToiCklMlFJ6euLRrXlgYuJRKQc9vZ+FE61AxLGeJKAu+rFl6+Lzzu3Ruvpjv2Z
dshOd7lVZl8afgEgB/oOS6TpjLTrygJJUWv7SuQdfTaP4FEICVwfDRDDBqa4YRGw
NJLwEXAC0yzw7SlfHBhbnum1SWo9M7iJX0bo8aqMtqduSRpovR5KT/AdpQoAEVq+
7gGlYNWWKgqu2/TqXO65bWUUwcA2JgcYpXpQNC5+ZvWzj4Kp9CfmEIIZEIS8s2/P
rfLfavxGTdXg1iIne05HZxWttaPPkGfUuXEpYFXZmwUsMWg4542oYxmZRjKmI+Mn
zWBFqSMmux1vuYZOs7YTwxjWhwA0Ds+NFQahU6un8OkHGBcGjSRSvbcD6PoVqkyk
p6UBUydzV2xpC3vnmOVjqwSQmRs4sy8Z/7fW9y2jXF3xbnHpL36Gewg2nUBPH3FI
P2reAyjIccKcjg+nO2aFCufEl1UmWkziKVtTiEEiX+BSfemmxgUjRm7kx4ifi4Yd
JOyFwRJGKsytVZQFsIGC+5gsueevQ6+YeOn8u0w7QvzxQryaDmje8uyABpC6IrnF
Tp5XJaTdyZlsSi5F0vOab7CLN0ILu9eVaJeA6s6o8Wp8+jAlRQoWFif9hBgR3VHj
m4z8sDx7QvBCzZqR4z6KO3UMir4FfedcyXiVCvHGtEDGBCTu3mn9daHzMnyl8kLy
eYF6iOLVdDOYF4jQcsvygKrV1XbQsSi5niQUjZbeGH1QBodgx/w9slBNMfDQIV1R
ltOs47cnVxH49mo1utCcaaeUmhil2bK3yu6NJ1/n5vNZYVeo10yX0c38t2V4QxCB
QYoTwuYOtEf0lYigNsKwa6ws01a8KSWrTkkqh2+QjSIt0FqYLpgA81+nK1y8xhtw
v+zJLibKuPPEIX2re3AFocQfRX3x2Ix/bgLfWM14+CgQ8tUJ4f5bm23wrBux32L6
jSsAtUpiVv2FSgL64yS2hQYu96892K3GxvZJNy9Agqj/CMmt5d8jGTFxWYceVGIq
+UVbqe6n8lnCtWj6ZZHOqJovRegZXb1ExkjaI6vml0Lsuba15lZMVHV5NYb5ZCUF
Qr7hZEu7bl7XmHIu58KgsTzkF1HOZ/+qJcVt3MnenJYjDfCI/Rt8Y2Ousm9qSyrO
JUZSwu5Rzqr4Pm3Z1u1+gi2xAXD0mYlFrPs1hogzXKs3GMB054t16ZXSpMJpOtOn
pRKfUoSqBC/E//OwJRVBtTGM1rJ6Qv+kQS+rlNUGXvHgAcRI4EOa1lLwLB9/6iTQ
egs4kEGXF77jvZWQhaFfj9QVwvIk8aj00nEXyapYztKP2GiinCnFUd/utGOceHCv
1ODPZMpCMT1qN8ampx+6HdOAgcLHb6C10FEXvXxP+35lbxBE106UTVoX6WHLZbtD
9jOqciz2r71Rb8tEPyN3NFSwVVeCL1T4V4Yqf5CpX5IHYY/LtKVnwS7H1lYcj4SA
K2TgghGtv/OxixnHyXCWRRZiFSadrHzyH+TN2qFCacd6ZIGCPOZnTpzSMQo9jNE2
LaqkhLVc/UXFqJosFNtUg+qeQu9qTv86sejWmhtlLvtEEVMNXK68eCM850jNKNrK
L+KysZD2y7NyV6s++tmsMYtrN9T901iOzoEsNMEMnR/ZuYjiFVxa3NYRJffxXTZo
0lV+rZx09Nq9ErmLO40pi8pi6KjAMY7Zkc6vShJhRhapHLyLzr47SfFnUZjGZ5Zc
CB1DQ64e7nEj588K+UvzCfFeSdTKlrGTzJvlu8WRp++792R9zZpdwRD/fEAJXnH/
vP9ORARKW/7WAaaWPHlpONd0sX3+LQBgeBiWks4RRuUeWLGE5nqZGJbnsE6atLEY
htuKj0rtXZLu/F4iiui8DUJ6JBRtiEt5U4mMK/1qn/1iYNzZVBMVfeivSZ19reoH
wuCIdsl42YXpOIHKofZBjvV8534O7LX/BFI7ZVkiLGl5Q+gMvhDgfWvaIuikmaZ4
VufONxBH2Kevu2tBxd2O/ApHGJw+1ocT6HRkShSBLy+mbC3syaw/SrB/jDGBUvSe
WtdhyHp4j6mlEJ0Q3VI++fRQ6cz8p3foAKklKwCU8/k5kSPiQdRtgXIwEkllyZ6N
4WlO6tfIjgmhUJJ6CqCVEXoogTKjeve6f/MaPKjM9PyBgdcQDItlObxEjr9KH9T3
Z8kIKLD0PMK4wxJ2uXI0QHhgRWwrfKTu7VpnQNPm/kYWzFu7BrpKPhLkmiqPwTty
TOc8X9VHy0eCulU1A+IwDWtsE7NtOhkTme6AfPd1il2FKnxj6aJjWI5B8McLNA61
3JpriqU6ZIEJWhWH/qZEyoM8zxhF67RmYJCZvcpPpFZo68fJkd/OUAQvit+pyzHF
KdIcxJFD+9BdHqh11pLCyXUw+PCFtrRTR+ATG5Vlc9MwMODVzxOhmI/fhelQ9ISb
em7/+tjzsXCXVdxhH9/EWC61KsfEQMjtRofi1zMdVJK7k4CI0YJFN5GF52S97xuY
TFG+vyNhGfLvuupOOY0DSkmYjxNMWnTr672mwuECm6BV1ZgHYNpa9kv4x9LJvhMa
LK1ofZCbOBa1bTMy91tZICp/at6VIT764gu4LQUqde6OzCL6RioxmV75R2s5Gm3b
y1n9PH3WQQev4ojmTOiZQALoXMsPuxG9FuNDIQp2dJGKF1Jg+1QWqM7SgFUxz+pi
6sBZ25b9KpXR6ho99qrFt51HMsxDNwHmoE0Lpi/CQUQLjhGlEXbubkhcumVgoYYo
E+pzLGxi1+crw0KYZjYZlFn7yS/2KtS0YFJzSKym4z9Mo1fYe1SMGsD+gYAgnJww
Vv3bxU0/n8qM7FYrHvjd1Yzun+4xBY203M/r9WaUQSscWKRAPsZKmP2YdUa8XTjS
REacpyay+pEuLJtpOZga/IEGATNB+llWQ0/QFx3NX8OQ1W6p1yBhvG2Z46u2dYKH
g9fa5LrTkIBnT2YsRNWuPYr0LOFoYcb7NXNytCHmR1AbbPq0Df7EJm3JIoXulg7y
94QmsNi8wHa5sOeNvyYihqvj9Qa3KlsRVGTAj1a+GudjJnXDhpXKOqdl9VF0SjUg
khryUPnP0hPwTku47mqTa4gCwm08zuQvghgycM24SO1RHN9ExxGA+HyIwxJ4UFd/
+mwvPZDxmXmfMTx+O2EV97s4u15HsvbBx3Tx5aXkumeHZYNb7/Z1aV2djsgxXsnu
uhQ4WKIZ2AbJut/M/zHvEWuliHOcTjIpIdh3nkgyioVPKseeBgpdiVrJYqRdJFdf
LQQHo08WU01ks+HDJOxGsH4PD5n72PpklMK0V1oANbvRStPkGKFHjydTBMv1Y2GU
qz+lRgPFGWy+muNbgcjgkzLumrsjt6dTPfktR30IWhlu5hOdScgU3iqZO9pxCX3V
2YmSBG8Q0AdQ+JH0kJOTVpkrK/M9mxcdglhrZzWb9/Zm0jHnIsYry22w4YC6BT8x
r2X1eN65ZNrOraiQeCd69oAUjWdnLPlHQ6GOxeuPxrqQa1GAG6fRSSFmCjUDiSvW
5O1eBlQ3DRA1ISVfShC4DYtVSVjOP2H7wzxPs0ccfZRXAp7vDdq3uXROwnWA7Qld
y1E5HfjzJQpTuwTtRiBBfBs4+z9Z+xDErq0+CPkbChZynSBHBnqS9zrCirCIEXCS
/8FvTpJQMCtygPA76sQnUJK9ft+s1d8isaPILxqOSyIgedvVPj0WVUIYBTkRh/0q
I5kVjYgCNkyOwM6+Xv4BRg3FRyUOiHRuUE8GIln5lHSfj69I1kAqnByRLfgx8fLM
wAFRrkZQzVn9Ms5CTsRfdV4EigzL0U0nxkA7rDJGWFD15WSYThB8YyfmzzlFfxrS
X6bGjorGnPb1SGC5Fz1sThLrMV5n2kfFstLYj1oIwdZgAPCUf2EGK0Sr3INQSYay
UwtB276vs+eDf3PoyA7oYx4NwSD1VezzR2S8RIUfqpfVTKj5u9zfy0ps5frI7da1
yvhHPDLUU8WWT8TMWLo3LC/GGIsfj69jP+5oOXCjlJoOgV4dLSUpFGSs4QxtG7Y1
XrxQbO8R3JPv/X3wBESnVbXf21BekFM7F7wwha52GX1nnyZDlMnGgcUdy/CbuuId
56JnoojH+vuxYEoY3PC++iqendWaWsubdtN0aJz2R8sJ9NMbZzjqJK4GHmWHDO/V
uL04e3/EwhI/46Yubrwy2NC7ROfnX0I0gGxNmGjGtrgRxuXgqfoP2NoM3Hm9nw/h
FOGpkRtTuDzFQNfJ2A3cZiHIc+GLUcavumhkbCo6obK/bmiRGVkiCPzx/WrWskwk
1p6kpzLFnEiD3NKrJa7qqFSAPDBu2n1YCJBMtwHHvvT+uNU0ByKNM6TI8l+byy/7
s3CMwOGRjrQVIzETId/PVKZBsbOlUxo1mASwihTO8u4ZlKi+onfwsXDFruH/LRIs
Q0s3Zeeuiw9pnBN44yvlQwm/RzA4gGjJ5vNbsr+Mhe6A8MYKoQjguEt+6W0JRMDi
XU5aj0oswCGHrA+GQzNEK1JVkbLa1gFY6/bIcUpmsnLCHesSgKa7Jp0VtspW90Jd
mOcEMfv0B/tI+GQIpGpLgVrniBYlxTzOPjAHJq63uQXuciLXl6qTJyrxP9cWlnLX
LMxmEktzI3AHefSeZ3kpXyKR5Qd+oge5dNzrBy4wTLwa6OjVoBdGor/s3WYyfNf1
K5YqVHfMbS8b3PsFVJ8fspCd0Hg2IpD3Y8+9PK042rpKKTgj54g8G4jevPdCaqzZ
x5aHFZmO6bTES3kbgkEz4vsVRW9I51V7R/xRmtsWv3NmLlpg45b+mLVo8zaDwToq
wofpXybgyZUDFmfkIWif5bXh9BoEwCHHBo8EcnsvW5GHEv62tnBO0UaVBkyjAHqY
n0T/NFfNmxmm/uwQnrVPLXRbPddXQXL2QwXCmB9QUCmblfreXY0cZQ22I9FLz8P/
s/UDkUl0c9IXcmmNR8HGgvD6Nvvqg95dzmclcnOar1BEYoBaxzyRvd/5W/+8hrUx
S7eC1W7DeQVlAlaZrLRJ1NieXm659vga6Sy17vtRG8N/xSzD+0AzwsRU9f4HAOTe
EkH3+5Ru9gewPPfp3ZXWTr70ZHoPy2b7wuSICysnTp3NwxBMVfdVIddpB3aUX9Nq
h9PgKhbSViju9gxOhjRpwaS5CrJckxffG2RnnG1d8Xb1opl1a7kQLbfZ1nw528Tf
J7srWcSaxTWOGj6mNbSOe/hNAKldD+VpIYA0ClfGebjtCxUFZ+Wry53J00ADdnO2
bGMHoPS25kR9j9gDHZ84/uteXc6TakgpWDTl+okY/La16FC3hYMATVt5BeyLEDz7
ryTYOd+96HLKfadLZdbWK/mnSiBbOcy1jUVBFRjLdqoZVQSQsEj2usGySMP5sxnv
2NeykOQInRTKPYEcRYM+Bn0t93JdDNUlc33skUu05M77rPAHshrCfAbi33Vo7nm6
posOcfdoHgf9hBOGa+Aps0O+B2+JVSK8zSRC7ljpQzDAZXFR5W59ELm7XkwE3esg
btoaY+W9UdPM8sHZo8JwBpGctbuGYKQggXFMXN7LWu7GRB89psjH4aFsm0O65OwG
iG3bFQv2FhcdYIHXpOctWvFJH3pjLDAzqlM8xy2pAuAJsT4pEcWKpJ64RBDTzJnH
YioUiiOymGoOp/Me0XTvdzrGLc4EDZ098LgwJtFdA9uTGlW8q/6S4EWlVxv0ySe5
CR8upSoL1LttEhWuGnojGLRI0tHH0fFBLVs7J5cqqGzUtqMrjB1UXZ/J2rF4UAxX
pv9uJi8VrJq8NLeuAB0nJe7pP+mRrvJqJrh+yFUozCHytXAVd4DDwUK3Vz+WmqgS
TRMlgRkbtwnF4yZijBUQua9NHyb9af6K/sAlegmRXvSHfcE36n2eFo4bKmPL13/L
g6GjdPavHEwWdXFiT1COpleyvAyGIkDrCaTQSKuBp7Iu8SmNY1lVifz2D52KnMSc
YYSUsMS7ogDOTAccum101ELlLhyn/kPZFH+nZlc90hW3sIDApnaHCC74LWl3AkL4
T6jk17WafsEGahF19LdA2ldUQIuRC9TiVBwKD/p171QaIaPZxpnlzmc+ow27vBLZ
dQJxd7KewfmHmMkej3ODJtd9nEE9nThE09Jji1db91Uh2F+ALjnoDwLsrX4XaGQd
OTnwtVG+r/Pz2rTGUQefRfm8iuPIk4GTSJpaHOVwSyJDGdtIL7pxRZbZbBc/GwX4
q+UP0GUrCA0/ujY9zy9a+atItR8bZJcap6jUVOldpbb/Qe8gJXMTcf/AJL9NRPtn
ZRBlef3Td10UC4zohbnloKMgpwTARra2rp/kMEvynlIyeavHwOc/2+UkYou2/8lm
DR9p/Balf7cW+GiaK0M7E1VOX+Q6bNdwePYyQV9hjm72woFZeEm/c3gYY3ZuP+t+
DMHsNgpF9SmoH40RxGJSVSIAblaHAjbbBHWskdDqmZVJY1I2yTWsKUmATaIYSkvD
y/JF0dSivZW309Gb8z5Ebnwk/WhQukxYXLm0w1tXmbjGgwBqKWMIb4ESY5ICNS3g
BD6jCOSpDFCCuia/oZ0t97nUCX8amo4OplU6LydTOg+T5bkj3C0oCSDioa4ygUDs
hsdv/ur+cJ8Fw411Z8fSWKdSDhN6H5UjA8lZ02MLGGvVWUIDfBKDLWOBI8oonWdG
vZj33TLPt1kGsdnR2cQnnB6XJ1UUo7N4CRfFxP5YMUUWF1Vumb3FKR+STPd4DkaU
rWD4lJxZcMjL4HtD10WsPDe8+c0uKTQ81ZFx0PqGil28lGDoPs1tPYQeWWOF4/xL
60uY8Y7GBV81jJKb79QvUJWlwQaqWIP0+wsBfGr07zjXmr5CyDGezdbrU3mQXCWC
/quElUR+A0qdYGPS9BddhRRM7tF2l3uN8NbATJnIShV5Ra4QI4iH/xcKgohZAiD9
A9V4OSNEDyHdOKDKlRQEY+dhl3bNkyMaZgLk72MqZlGDzWAW9WAMC0o8J/sHAK3U
ayCynGRfGrvysHzT6UorCy1sLPG/7PPN2B8LnwJGvW1346KnopHYyL6mNuCCVN4d
LTtLVn4ZwFUgNryyagPzuLXYcJx/KLRxtC/nWxOwDt78V12dUcX7w+wn2VvJbi8f
+JGxEYI9fp79TS/9w6cdON4+qcp+JTkiRMxGOCCbBjU3CcYhyMOLV4MO88jB3wp4
c8qzeBOLrWxGlrCK2M+Nm6Qmqpn9pZBAs4SnQQ8hJu8txOA4XeOhNt0/7H+FX9Kr
mUoFbLAhzLz+0Fh6LSHmnSA2ObaCJH+xHuyabfbx24vwT4P1QS8+A6NgziwUjDeA
PvBzcVlovxXEkyyaULmCqodApk+xctyYJiHBh92kuomQjNRh/9pfM3thEdDh8oqc
fuBA5fpUfDLCPgd/6YunTb5JUeYrSzgeghLqqLWGia3DJWqFsV41eZ9WPx88OP5s
bGC0KdBgUZAv7J+W2Ik87N6+XBGcNvdMQp6aQg3u6QH0i2SdWQR13sm3ZLzC8R7E
hZ8JnFQUU+sm1b63jVtAPfMOHCLy2PpGRZ2MVbstihDSNYsmB+nkxvr0jgBye2wm
mRDIo8zsdh2yMO0kr29dJNaqSHtmxXyrWGIt16IiUffHyxTuDdaF2+Y9+VhN2rHf
b3EVuUP/DlEfEfoB8S3M8KKQ9Yyo84Gjz4qQig52fwLj9fo0HZ4ppTEQbzxaercS
vysj6yN5X/VEvHxroYV9mPOVgaB6/ck15DWqH8osHsgDX5vLvI2PLlKTZoATvyqp
Ay8b8AWY2NnJTdpcMgVM2iggwCykW488mOZ4uwYXg8wDSFsL6gM38NxTpkUJtQMg
EVC9C4Qcvzi3cJKV6zg2xeId6C6pEF49GMzHdu//diLEzXCmCjRodCW+F4D09KEo
wLL1l8q1xMzRV5zcjS/V2d3iZcRgwnL3Lk/M4tfFenHovGYj3ki2gMCWjS3lagwu
OU9N4SL0Q+vg1VvSuS+yS/PpucpC1UPG46YmMCrbI3ND/ACa8A0vegMC9krjylXU
x7UFA+JWWUqHEJxsUVdtZdA7gniLI9WITBrQn30gcgvrXKJfzgt9BFyzVkzfsvYW
7gHFocyHy6GNP7fHIoliUVSbtp6ny+ZF129qXAuWUP+GXFY5/vcFR+/b669j5llP
Hs/wvYESd1BvCGaVgx7y3h+Ebi9ojSioG4M0zENQC9OnIR1lPEGlc2s9T4Gcnr7z
IYLEbOf2UT7DpzTAW4KCde9Z3T1YUUkaxFM0y+Ld2K3rqZAP3QfoOZ8b7xJR1Vo4
Xyiw8TUCAK2T2MMGrRzRHcxkrLCTWNmpJty/EeINySE5zfdDGex1U5ZEz2JKEZQT
vCj57tRYj42VYzl/wvpvEtOrq3xP0ogApWm20h/FK133IBarCpCZyjIPv6QRHlwS
P96Eb4FkdS1+heH7nY0vFaEjk2S3Z34mj3ADqMwaxBDJ7rpvmmut1/vS7CNSEojg
meHOLtPIUyTYCAYpp1Yxafp6hBtfYgOO08ZF+V0WmSNuFKIpIdbOkPodc1SRk8Rp
nTfWi1iG8rFe6vTlZu0witvo00PHSKyRz0Zm1WmUOmbmWb0mbca9RUh1U3/Btoji
441zzvRSm7jWKkss/opxOiFqsjqFLaXNo2ANEtJj3Z6wcXNIXfYaac6y+i1LoF0u
iU+9by6W35uWfOWfaBF0p728jarnNGVZ5/TVX/++gps19IZo/K31FIT0N2NntDUh
u5I3wAQB+2cncr1ZAkBOCbqJxS/sE5y0JOl6DaHODJiqT0J2H7lTk9VPj4TJvS3+
38ZQzf41kyJAQcFbdIi7UKVu+YtIQtWALhXYXGL4Q4O5TgwhSMIV+2DgHh3RRu2J
p+pX3l9BBtnty4M6KGnzCcZ8/8EHFn195ttA/WuSQfUKagN1BFPFn5GyQQSZVUdd
k+FXs1OzVtI9V7eP0aLRA0FnNKLlE8eQHmY+0ek17EREy7wByLTyVzCY6M+gWysP
lCNp3HS+3zITQ7QqbiVxk2jlFxyeoIjsM+wGTvwG3U8EAQMnKu5EIzFaZIWVyEKr
E+/UfCJVZ9Ini3+XHfuzZbwfVtyyjkOlwyCJFXAR2C4kca0/9/lRHmJPLM7tg0WO
jFGFZfrk8oNQEGlnaKmhg7tgSQZlR9P0GF66HIrxKbxYEBd8s3ssrvVdwUJHleq7
hZQdfBkgWzD2nWkVhEjwd4NRDgPeopC3F6zbXbAl5g5rLHJYLDH8tmluQbKgsJOV
R7DWlhE0TSbTWSBfabLKB5Q6SlAI2HIM8K1JTFR45ChPNEGlupaFV68mEPiuzk4o
3nkO7uUloleCw5JU8xsyJqflP69V6uJd2i9AaJFKsWMTytAbrV/hIbwmOS7YTbDy
zsNy1nSiV84CgD7MmovV5dbX1tdsUPPOwFMI/onmpFEuv8bzAtQvC6luApD8gYmb
Z77jzYmCZPwnrMvpxjKVcT8j3OJaNU7bDeuObEvppieP4xmgvMjVGme8hJ2fTJE1
poMjt+/HU84A9Gfwf9BuLnfMjxeBgLIdZ/+s3ymed/ZgrzInYBQ3fkDpq1smif1s
pXCBo3Mh/gycpw2kWtTysAvcjth493R7E7sGm0UiUq4Y4n0dja+hWZV73D15VDJr
SmkuytA81xq5OvnZJEF638ymHZZYYOARQYgGOKLIkHULDFeBg6SnvPcpUNJLIC7O
os67sPOHfoKB/HyEyAZ48iT+itIxtCyPTKMSYYu6RizZSaydbMFQ4Q0Mnz4qBlUl
Cd89zys4wwGBX7F6i1wBv0CvS3wR8xNtVyE2XVjNXkkghtYm+5vTIAUPPCfTcDUP
Tq9OKwfB2+u8Ze2qEZIXbn72ziGcyvlrVVAvYRvP/aN80hQU9v9CSB789XhYY2QR
RXxP9K0NOyfdxmHugXG7bRp2XKm4xD3Fv0cwB6s5vDNqy+UuXZS/CUX2S/3ku4ln
+aLY7koTa0dm0UUFKMRf3bNglWzjuIZqq/GqXeeUVoT17n1SZumNAA1jDkmqbws7
KNeYTVGq9yrSTsAykN4BXrH06fXEv6QeLdN0wKy2UWZ3twK/krbgT9CUuu+Jh16Y
Gt1ypOohCcxPiyMoMslLK/wgtFfEqtUeHfCEUjW9OdTRayv+iGNUVYGPeDtciCeF
JLnKygMrcFOTvTRMrvj+u/s/t1IaPHLJhujw4P1kDlaM88q17GGU05YE4ERKCiw6
9Sq4VIIBUZaM3mmx0S6aN3/7c+5QHm5jy10UoAoXISVLKWJcDiiIDVIOcXqrIJt3
t6bAjPQxKyAYYClaNMukcIYLJDv633jC1O3E4lqOrThWtAEUbvb2PVW8MFSFgyGo
J9YsqyiYe6IGWtCun3ZsSMmaFLwc0VTDI9tmvYKYVaGm+5DSmZgXOkzZcsQpdGUI
r278dKH1fvTRMtAp9GwbXBjZBR3TEauISQT0wxXWIQ/UWegfkAeXOEsTtxNZueDD
QPABY6BnaT8cBFggn86O78ZRMD2I03pASg2DZo7SMmv2U2HyuCG4IraAa9Bx/YGC
14jBsrKaCECMO8JVx1VGLet+DAcIWY8JWg/O5MKvllG/v8M1Z1es2zt7Tx19p4Sy
4DERfcbV4jSQLPeYlgQ/PapT9R+KAbl3B89JsKhp9ADPDqRnMxGEhO5CdZqqy1zF
aO/WTrRXtcVr9HP5xgRR4G/HZtULpge9MG1eKYfxCotWbDUtGDDDtllo+iycVMkn
FDNSOsa72heQUkNpGhSi9RMN9G4BMKXUcFLYeNBXS1re/SQ/6T0aqy5kNh06Bq7n
kEQljBf134+OiNjjxWQxKjiPrTodYxwDkFhGwSYeLtLs+7IpXks8YCXIlvmSNw3V
2A8d4MlgaQbZDtZ+dUA9wueGHyPjmFjvITt0y/LhBnMI/iSPvffLwOTfgQBUUpb5
hD5vz3gdPXnrlWIerB83ahQfRy3e/uKgTX3bqrCoss+gm2mzodSxr/ovYpi8i2jZ
LwxR4I0xIQnAakGxtmaEKJCRdgn/OW4Cq74kC1rSA36i7lOLG3s3Ka6tqLtly7lQ
ByqLNgEDDzrckmGeKAg5fA3CFqCf8pJ9pFS3iUSaUfl/i10xEaExZkC9NyFbDfow
9ZzefUiIqpYcI+UjdO9k/5WWmGdm8PK2eYUjvD3kum/sxYEqxnLqNQKJcfa5sjPc
Lgz1PKqdkd7Vri14rr/wuKA2xaqFenOlXXyNLE44lzib7wivBkPAXwzD8p8LYjPu
zAyd6OEi+do4hkhI6QonKXJ8/TCbM6p833N3/+q3Q4EkI38iuXyruSliuHATevay
j48J5B6FcjlJqD9LcWhU5x/jzgu9+yW+0kZKWOgbSIrVWedjOMP2OL7ZvOzgwGyb
IqEGS5wAwSO6BFKNphkd/Sdp89xv/o5Upd5vq6TSrBsuZxphLRjLCA+B+Kw6JUcI
7eyWRnl/kFHusk96+ythbBiFEjH5++ymaRvcKgICxjWuwQ8qbBJjwXLc5xcEvCu8
q9RAC2d2HCmrVrddCGefhwGd5/f05y6rSSmK8CSEdWU/bz8ze8Tflin+dDduoSKq
NdYaKf9D4BCKY1847M6M7qef0jm53LOAQ1SvZi5wVlBbcInTIX5QQyUnrFkDgfOC
EkRywhmUfblH+lQMJUh0zKctQCyiaCCmKgS/mWDPzCSIp8L8aPY0+QeK2NRII6mQ
ssXwhnb3bWJW6eE9aORMXBgRiXPs2zOjhMsogqpGhNzmkA3rml12QfZaSBrp/8UY
4wv0z1EcBwxSYD4LJzpgqFGL/VnQnDlxIXt9b9+laE9Z6vw78jigR/t1waaFbEVH
3Ai6+pHcayTWDJgyZ+cododQ7N3Ry16IHc9yjbF8JIb0M8nHExjF7WvvENFvUNNe
TMH8KbnOhkXff1dbEud76NM0APav9JfzPVOMJpxA4VUZNPVsJviRXlkidUUSfH36
ig6rc/+nGJSS+ugP++OpFSGdr1YhDduzfvsTdGJvdARNNu2GvPdNG1/nQ58wI4gX
0hk2RqdGve9hV1GEg626LNMCPVNCAtCCKMpMcihsv6NG7Y8K1BbVptLFgVSfsj8w
iCbNf8YlkKZb+SczblVOxsw1cpRhajw2jPcMsdxImSzkvuxCsGyH2fB2KMwPvnHU
SZYJKPi/4vTvQHvcN3VEHvwqc7o6TTalmJU8LgxXCYfEDLhqjj+24uEqXXoBfCil
oU4qKskFmbGHOcr2FNpWLQ6DDzN/n/fB5XbikrmxHYj7yKGWr6cbhOiNn15O1KEv
4a7bS7etvGDn1C2A/V80Pfig9q3Vqa7siXjluDv2s/TP3mYwQFNxvwtzTgzrcG3R
nZVTvAsVMbU2UcTjnEX5bMe1BUlfgQTNtZZd9eHbDROEBcUn57AOukKpBB34ZCMS
eyanBMvBBldBEg7QCS4tsAincknAYJZb0denyslCnXjBW+dhEHE42W4SLAQrIamK
HHImSx4HfmLADhB5JFUr6sgIPSr04nLGrOTYqezrF3Ck4UCNCHap3yezv2dEvOIq
RTlODqUS8fr++TsE/zyg1wmOI0ddK5aTyi7XftFNkYjtpD3fhiaewt0Rf5jY4dQe
uPd7Tzk58dr0NO8h1w6OfHjZmRDZlHJwqj+PA2nLqVu0oQ2P9wDqO8jFP52NJ4By
jsNEBt4ZMml2xFstwhqH2C93YV65hOc0eBypPJ05fYYOuENM8mWoOIHlc01LDE/D
3+ZCW/1oXvC4pO/geMxljCEDwPVlYbY3HPQ/nPau7MuVLKOGHXn8Lstd0zMZ1n8Q
azTNDT4ugrXQVfwfshJv8/xRYDDndJ9DDamQU6yaIEIAUMUFqRJdMmOsgaefDjsE
FYjTLJzRoARMtWWwkn7JJCJ2w2jh5VwVTYWAXxmrjJ5leLQl3GRuhe6PCw6RiZxQ
SGg/NDjbLrgS42vnEhLE4iz5IwJg5QwOmcls6iEvbRp9VJouFRonETvr1lptj6r4
zpQ2UkoTrCvsy5O7mdXAZJmsOMJDp/ztHsyGJvSWzYwgBkAPUcr87vlb5a+AgnzK
KYfQvx64QcCeaf2MyD6o41/HD+m8HMipdMbuAfBja6fBLZn862YlK9NmOrt6VnD+
xMCt0T8dRQDn1DeD9hXoEYfSSBv72uJDiL9s7cNYJKRfL2gMwdU3TIn0ZYcfdxaB
8+HdLQUz0msrXKm+t35yrg/iZEZMXLWw68bssGtJflcify+TGpfMJWD5bwP5tqCo
w7GxLSB4WAGGh3eyldPMLhhh/Kc76PEM4WWMoJ0VCBOYZjE9m63Z08ZpPM1AEN2d
fVSqYC3rfqulTQQnZx/HPFhaQ00gAf1m2AA6D2LCuCeRgm2aM4olcffxovqa514C
9qJ5Luvy9K95YNTYWss2g42IuURNzzyS0HoNnFnLSVczfghD4252Ewbu+UFKj/cG
WRvRSX38SpB4qCoCWyMY1Xb65HkjWALyjz6HMYsG8EPlI5ZFRFZPzOOlZeQ265Gi
mMFhUiIKfsdj9eJOv17ca3N2NdEtkdNA17zGB3OeIqiCU2m3lgqwhY6cMEBw2lFr
Ig3p9KufDRwdOZ/1euTJTvdcAk0Vvpx92GOi8wRUuJRHpdcjlyT5oyDbWUpKkQNn
X+ar+5ya53gyHgphnPcifA5T3ajq/ZzpbD4GCofoEFiT8kCx8NdTrRNMxkeYLbxX
ZX8fJK7yr+EHg+SbF08LH+98g6PsukkhG7srZAmS5rxUuorlXZIR/m/DvjymWkN6
kIYeS+JmftcirZ5Aqs30JogssJaSsl1hfxI2fKJcj0TJVem9bIlRmXsWhjnxOs7o
facN+9uzb/7uvHIDdKwCeIt0DOTRaJSUDL2v+pvu3FFf838vGXCMx2lERIVyUigd
6qYrKKt1fKSkhHiGmjPqQDVUSrRc14PQ+1jKKfkIvfnNwXG6ssv4dcAch0OIGNo1
yPGO9bb55LjNG0YNSEPCq4fcfu8N9ky6Ja1VKVyGn7qJqyTzOAC0Aj1fxhqr0L1k
2gvT3v3KK6xwoxfArfu/FPeKl6vVKIZYpy/ykO2mLOsanf19hQFr0Vvr0P6gmPYU
oVzFTwLN6Jr3CBRF9l6YyP6DB+iB/oFpPo8KCgHJIUj0o+Vh/5jbccRlrUku7sly
ohvlI86GGLYBA3e6IoOi4+w8e7/rWvapBl6vXhb1ClwFukBkNZ02LU9WxRkrQ6j5
wfIvu4aKdy4BQxcdkmUGwVyx+slmPAIBliAjfqW68Z/ksqBDH56ksv6Ue+PQy6ST
czOjuAbf7KGAn2EWbcm0RcB4STgt+Gxz/1hLrrQD2Hj9+Nq0HnTLfnnHXuS19Y2Y
apmqVt6Bm6MpwAx5IS19zsVQfP762YvoTKEwuTOU16wsb3tc2/B6dDi2Dvooph3b
+H+0mG4L9p//hsf9S9yeCk6q4vGIdZdlQaa0NrEy5YBryEpZVB/edQBCqUP0q1Ki
7lbmZMVq0h7deFvkVJDi7sZvR9NLOCi/fA2ADS0HXoAqqp8bIvDJK8npWrCh2DMp
Z4NrmaJkaDw2N8xJz+8gAdPdVt6HLn4qeh5YAjDLR4LB89+wKflUQ93M56pkUk7V
nRniNRXPfPNuFQe2a7YlHTubWGnSmtGjYqjthkZdkWvyBeV4DrZ4MaovIPnZzEUD
DujKrLnUXYPL2OC+tJC/GM+j6H+ABGspxanb/KmVYkbWmFUngBvCSFQHOEeDYV6H
8bEOdS0lmdUK+zpGAyoq9Eoh0GlDtJegpMIRljVu+owuYF3Ezanew3t8fks+SEW8
fXPZMStODBhoTMRtluKsTSE4w2C/FLrLCxfzR7WW/Kk+jHukY98xAcS3J/uwddct
jWrT3k3QF2KDEC6GhA48E6uPjFuoDclPmZBeY5pkaQ52QpFOe6tqB7xWjEvoV3/4
Nk/4Tu59Nf0VrMDZmnX9w2mPWrKyipoCaz/0fejvF32vaCppf/n2in+eyMC7BsAv
sDxylOJEp1VNR9lHjCTSnJtrkua72HOQSLeinvlsIPCVJNtNtpbcvD66zs1GXzgg
kMG2QhmjipV0tJp+BeKO/BHgMbRyCUkLuwt9u9LJrBO7DAZS2RDcuN/czcWWxHfP
NA7IqUNGdCDbvM93cDiHXMU4xO4beP+evU+1jdr3GnwNZg4IruGZN9WkHNP1lNeq
isUBymqqN3FjXV9qPNQyLg7ASStj6vQlBdPsMOvpWd8lftjeSepqfLv1cSyp51Nq
/c3tzou+cDMnXThQXeWR+u/QAudSxIenQkb56kZ3CGov+FGQrJDwXXJf+dTnsK2H
QNUkhUJALHpsStr1f5nZl7q71h5hwRbKvHbzqQ+S9SyGSe9oQl02h8LMS0tT3BoZ
nBtSnJ4NJdwjrkHxTtL8KNxCSx1rmfkLCG9eu1iB4q4ZhFk0n8+zalPeGGDZc5Cw
YhDfSz30xnIEWS4alsTUAyqnd2nxceHaGc0ggp23luJP8n5Cr50klncgeUrdJapv
7TBiGCUOh7GGOpJc17/ZlMO9J/ZwgaSMF441CBLl+0rCuiZ+ySMhVy16QbvmFZD8
oN6TxskokBi7eP7Vo1RJEGa/7xmwtPPATNc/dOtP39WaDa9IDA7qS3MY+PwjIzvm
KUy1u37MmD68lkbGyhBeZP6su6KFFD9A4Ci8q/6nuTZR/yQ3cPPyo/KiW2xhA5+w
+414g7ZVlX92eBJ8fD+ioTJbyWr4011EH4Kt3tB1DtzpomK7rLlNEltRc/fNEeVc
jQS8Fbclr1n/AfhP8yCN2v589+ae3aDhQlHGrlXeFn8U5CHOS2cWFWCx3BTdwaTj
wRIeHxynQXa0PklJANAMYgdqdCYxDMMT4rg2ZSW1A2zI908pSc30cWH9SqAL2Nlq
yPekOyoK5mtrWzWbhW9/cXgRhZq/MNN/wKpwjTQA60D2RvJL6nGfSbFM7Xp9xKNZ
QQfrfkqi447nK8nlzN4v+wQkibmCi6BUkDg7NjFBHnccrmQzUoMzP64m6C+dK5V1
1HYSeXHGhuRypQysAswNEL9bE8MnJElnuQ65jpimE9d2YUu9XFmxhfzpTpm8umPj
5dOpLvhDO07/Jq+4Z7yL5vINA3TEO2K4sQjD/JVzm+PlnV48AABtUgSozclQUBKt
Db6Os4K/22w+IPaEFgG0pI2p87mn6yBoV+wgfpLkceHpFhvJR+ayxQSZphXqKqiG
K2lVq1TXmCN8kEcVkCOBWBGJIoC4qwWBVwDwY5TFn7l72MZAcA7sZwrfzt6UtiZL
XXVV4qss2NO1tBLGuxL373KmWBJScvm5LAwYqliUHvC4BKOm5/iQ8Hqd7dnlVY7B
eYg03rn6auArsXZ8jELxNrT4Kd2w8wVH/qGw/w5RejbdD14cIUvt3IP12yod1i4X
0JjBK03mrx6SKy8nTrDV3xkrRzNI/hUsoZ/Sv6upCRRbdSaecfy8IT9ebJzIF71v
oEAjdcs3gjKARmIVtKMA8xUNdrt54FI3fR63fAgFdqPsv2tq7YVRZRUgg/hJVY3S
T51cavJngO6uqBH2juNk+ugTuNHZwZcqSHWsEnhN7SONWLz4EKhaFJokNunugLi4
rDwV4ykkvLW8xPA9DG5QUTO6CoqIFXki9Jrmy24lJVvr8M1cc3bdaz/LKndihw5u
oUXYYSzg2Q3n/YlWvYxaj09f+aVvyaA450QbPqfOAl2nLqRQ0AUMVJ8Y6HKk7+tQ
znF4T7Slx7fWi4/lhYVuTAs+zp6lEzjCPTgbYVuZ9703afvUZlh7goa4ZBXHxKRM
aPSen5OHKkv36tkEtmvWRbKfbOVZnhW7DQv8xHpXVGF33o8rVGfhz2EMWWmsKI9l
DDLPyX9/Y2dD1o8BwlpZJzh+p+T6zdDdMDz0ZsMQgD2WGCvbc1FbSWfHGnBUO9xq
s4ROJNgJ+NxJjluvOPU2QBWsojaS5kxLrBKquXdSxjTXmmh7E6IT9xI7sGRgca/6
6QPdJtG8wVH7nFk7T6xxs3KGG04eOfYYKhozk2j5gzKGq/NJboCQHXW/MYKlj3U1
mrnxFoDCIDlQneDk3Msh7zYe/eq9tHs84iPWrOHZLWQoCPOYgbxQ9B6zIkjFiJpH
ZovEmdGDxL8Kgy2zmpRmHrgvw6lbXM7ctKattUsjoNYi58n/0R14BDhtoj+0icYe
1kseDp13vxSiu8go7N8aIrx93PzK7JcISyZwW+/IejCOzNEazzGTdN+YXm//o0Iz
8LaHx9ylzD6WxyBBpACdekts7b4MxNb7jrYDeFqdiE2hnA3UqmLm2KLt+0CeD1ju
Gb0DG7IqKHkDpTNrx13PXyqrt8RbsHk305447BO6CdVR+06u6KL+4zvvQoHFOCKc
uq6FANjwJ/Axro8E8ki2bOCx7ajnIjv7/E2i6oq458/PIvqUzzSNlDKzXh9oWce6
nAH3u0xZdVjb0eEDunzOrnUY+R4gDierPtlJkW9bDLxcUZavpyzdKpLCvJwGXouP
Fa5ybTF8FnZ7K2ymHfkdx67bOS1ASuUAUCT+Zq3XfucSy7HJmZVmo/eoaW1BvKkL
XwJ0fZtU4N6zasw8CUasZcCwtFMxyNI842Ach3cC9AZVrWGNdYi6CAh0o+Q/Gfdi
CH/lUPBuQt18kHSayYXYKAbxIOMNtexTMDcpa7ZQW5qVGUu4vdz7qO6n/6z3vRsU
zw06/uG/N4OI7AvXgQZ5YG6eYi1/HCwk+N2FMMKF3F2PgS534/zLmcNl8zXg6D3/
OrzuhjZUO9ahCYoPM1YcMVG9XReTXyL66fVmypuhD9wTq117bUj3a/AdqgnJYlXh
Er1ur/O4+abz9e/ueayRCxxxDvrRG+zsJOvwkNCsGDEbse+0uUz7+xyUyZmJHEXl
+qii+NYwg/0/Y/bV/7QeLKGTKC/b27NlhsKTAjLkmVYplCf2BnOTlb3G3o3yn0wc
CrDaxvTz1qsc7ssWlvXfx2Km0lLEMNcDSs92auXsuX1yVwBJCwe++zEWRuBXLYrO
wGhpVbSxv8dGc5UKME/lOnhNrEdTefwz5ZSTVTOuIe30kmpKEt62Aiq3V+Eg3vPU
TvwEC4OgoXmc2ElvMuT2m1rYu7Jn4rvmJ3olT5DYsdZN5r12rlhmHFsVLPTy8/wD
9/rkIHITIcg315VtEwcO1JIOlIDNiSP1WaixzOIkmX0SUzUcgFq2FoDP6dGWdYer
XiFc2f8ewi07/MRWPCFDtZqMRd59IwcDKRNUv+9y9YzH/N8Ysj+c+VW/rcM+waLS
VnFVxuUNqd4I/l7yWinX0Bb/3anjOi1D1gdroH3CAq7RHGxXYL5vqrVfYhr5pUQN
bsjg9a56hKe0R31sQ3UAp/bbDzRFGZVHOXlNRDyIcX/0+KuKhNlK3pnl/ywFDqYB
sDGAlTglKBgnWWXrLDxqEChgF6IT9fbowntcILMZuegPgEP1Pzjun2/0JiKLp3g1
Uvp553JT6zi1g0UlujJotwCLOw9pyku5AkEEQA7ApemAT/aRnWl29tdZGMZYhykv
QFWRoKe6tszoOQcQwNuUebKNu2KjdfSqzih44c2Dw7MxABAMG5pIOB8IwBJXJWNj
WhPdygbXCpSITiKw4w0zw6VCecZlW3aHKY1b2EDCmY4lXwb6dT7pq4ByJ4lyto2H
N8WjkXUfWrpEirUHuz5HzjxZwOG6Cj533FPeEx9nVjWNg03SBfiOCTokRzfD/ryU
yrOhvp1sw/IYkXMqAOzRpw58f7nBqImqnHErKpm5Nr3Yj4/MlXipPdmU7tEVaf38
4YH64rNg2P57utvRoUmQtoOYmE4faZ5j6v9CnlL7TMEm94VYKQqxyVVEW/ZET4B4
EN/XxPZtIjow36jdJmu38SkMw7Hi9kURMBFaUeabuQs9apMN8MWCVFw6FikOJ7cT
ltOk30lEanm1NawmBT9hIdG4RqmAn38wYkMSmrSQRGUehKVc8IQD9AqFB7d3RwNS
Od/Q0kurdP/wHI2i4m1fHuY6dX+ZtB6WNQWe1ad1hVixLS5NGpdkSawRX77zqHt/
sPEzN9r9L4HkjIgD4rlZekd3CsacPu/qQ+BZ8dmEmafogc5kM5ahebYusauNccF1
vcWOTH22ewgRDbjoY23AoVaOrJ8D81qz/XD7r4zuA8klrSgsTHQ85aM4rWi7NEna
Tbqn42J/GGUtQO9iMVpZNbHVdXm0bH+hQImr+0Db5y6rpl3lSTHWeVId0piUdPv0
6RjEI/kn7fQqr/0Cc+g0tj0K5Fo/QkmoWMM8/lpTR/70mkW3FHA3aT+DMvdmmEnO
O2dXAOzFl0vnIaeh4G921xdDMA5zfIFyGh8mXvs5Rsy1sg3O2r7JZP8q4MRB95xN
UYeYhKQQcdkZz5NwNAV4eTb6ok2RB8Saapr/momxFgN7kU5L1MSOuts0wRt6zRkw
1inNi7O7wovLvFx9PUC4nheRUi6WBZw59ITUxfuLa7IVf73tZUpRlR3NgTCDKxWD
wP/oJc7r4sRGB+2j1F9eu02R+OfHgRKeWOLc1WneXvZBD2/hw69pPEsQ0f4PmYZT
cFzZUl98juBHqXW5feoukHIBKD+2vjQ27uZUBiowiCryerHWR/L+HVSv1ENWzIGE
FEYYFq1MOT/cLjC+QitUGLdWJlte2GP/6XEyW0XeXqI6MdnZfglGD47E3qyGRdf1
MhToe+HMheg+P3eKkaAskhq2VzIDzAmblC/uz809XqqgpdTj7wq+iFDg29U3wuhF
X5KoN+QxywZKMNdqgsBrwW2TrL+w37wm05l9kZwl+te7CkX7vMhKJexUUd2SLN0Q
FdfTdXReDSG5jugsBbnqvdQ4Wv2cTzdtWjwCv9gdBilcSm9IM3WziQF2vQ6sURap
N+XJ21dNShh2O8xxs374g6kjzjvCVqAMasz0rJ1MN5EUcHMpL/ZWCuw1KB7GDpsj
zyTQv+UqCUbcgL/IsoJD2GVln5oNPHvofyHudjmAic7TLHkm5H9XKhSQgIwYCatU
6/lH1vyvcI2AtEcqS7en8Yt+bP5JWD/rjNx1/WozhmhbTXYygU/Glf7J8nl/ZVaJ
KiRQ6h7cJCyAHZRAG6+bi6e4kVPBfka5jP5LBa+29i/hsD0TOZJhzRM1+0WDplhP
tepb7bCqOytYYOh076hYzF9ufLtw2FkOPo654Y7pLa3fr3D5xvjFBxbdSN2Gltc5
2yc3I9JrNRqgTiOOW/5qvWSep/8FEZVG2gEOyrswAOR0eN6as9SqV2aVhp1w2o5u
Al79RuBgWod3yjiBxGs7n5i8Mm0MUcOFcRs81AvvROAsQgqIkiscsiLzwGOFqq8J
4I8rtKOyXL3M5LeO7xgUPJdfptwHC1Up07HwLE95PVotE3x/TCFOpDEG4OQ8k6b3
4nU6X3dq373pUaz5urUnMVwVRfvxbXe0myXo79VbwkteMGrgtQlWeydXnKM8B6h9
x24HMlfBBCErGVF0xS53pak84ksavLp9LDLqM9PJBXwNzAA257Qo61S6G0ci4EeO
3kgJMLVm4l3Fj8KE2xGwpXJXlkJt+xeP7QB0TZwi00HG9sLkBkAmO9TkzJI+cutS
hoxVAHIXKf7UtTJRekoPlJMetBkyDVEAuRayhP/fgNbkf94RCDE0nh9vrNycf71M
Uk8SL54VoGqVLzynuSwSJJiTr8juC+R+L2i/fQqmTa47cEj2yGbd6o1fkkwpqfnD
yPE7BYLs0PyQRdjcrj+asFQppRWSmhkAb5/2DdP2fMzZE1Cl8AltSRy38O47sJJc
OXqhXeqLsWUgIzYonduy1BlVGHcq6geaCIJa9U8mwvVrivepofrLO2CF90FmghqR
O+ftFf4IY3V/8lN/QzkeJuUUasVyU7elqNCaXICx7jdmNnLWgpvsqa2C95TyBm9T
Ag7XbzwrNjra0++Wk/CE0NtWH1SwNd/TM9879UIZXaf/M9F9kUj0wcScjJrZGHQC
PkAUlhJmS6CHIgs9yAHGIdcjyC/0VynD+8+buKx9g8Yxf/elwjIAHjiuXUkGB56k
aXtRAoRfG0eKKv/nsP1LPwZZOx+r99F/D+ucEoYmRtnMJxpfCr89ilAcK/V6mx3d
kXqFW5qk/Y3/eTNSkMtHuRbw1fmbTNNA7k79aVuC/YiKARniEAXB+q7WgWvy03YM
f/tssSFpOGwbE37O6C3dSOmsrNvyotCsuSQHo/YwEuv2kss75mwz4//3IMji6g/b
WTRp4gN2IwDTAQdOZ/2lGRL7Iqyo1omFquqb4heM9BxRwF9PMiRd9XFN7ZAYPg6t
3r2XmmTPcYciCAW+SCzgwLlM2j+5mTy1Pjq+zrIvip5TdL46GgTOLexmuItdeAVC
sKlhoz6SFHsVmVC03/WDk8TLrOmIEzuEzaNmdc069xhfD6VKP+mbp4FWk0+af/Vt
mKwPv0hkUadI3IT8ZTswiCwmMX6RA71IWLBB05V+D3T8MqEAlsXCXsNtzHJ3Zd/c
rm95MaXiwD0tClSFgu3BFB4ZmN5rCLs3F7dWtqEf/q0Cu7Pnskpd04Ivw4Aut00C
RELDymUA4qf5Z7epMBoZ0nu1Z5URoDRnV7H4Zrny8n+v6SXh9kydVGOKAVMNu1nb
qMq5wVlQHSn+5x3foHj0yQgR8rTsErrdA7UrbCbd5tjRyiKHRMr3R6m3S3vk09vL
z8RXYSO8nJo5eI/HPY2vA+F4TJkgztebXR/rSp8mN8vroEZKI3GG+QVWFNh/WTIQ
kHn6nIerzou4HLwOkZ8XX99rBx27hBwy6l5TNjHHCWZcNtHk63Jy0HQIttmW5mPv
UjnwDFrL5TAc5+AjQyx82VUowqgF0bCxjTnq7y1HW9oBc3aw6jQpVc17OgOQ2b2z
6huPlsCdsAALpF5XvgfvDaZXeFB1Q5bOPC6I0ezLpey3MyXVF2+X4Xfkm2+SmeIv
SKUTwVi/JDc1T8y6y0wbPBL6oVORXtZwnwFER4lSFu7eiWxwnxBzikPe/D+jXtfy
H3yJih1k0R9kQ1YJLMG/TmZcsMJw4kUYmvEGZw+GoXivZWr8SJQCVoK8pax3cMui
a25JTXd0zDZVl7vtKDuFFyjF0g/8JLWacDQl5/nCLilYZDLkMoLRFmduXzJy0Uga
AFm8eaLiFT05Ju4F6CkfLJNonScn1yhTXafM/d4RmSP8FbTbBdwzYI7ySXxji17k
skW1b+dHgPpxTIgaDWsy5xG3l/OsmfuGQMKeQ9pWdqLGmnh8IRbalLP4UgkznHCd
x8ppm/8md2N15F0AiuJXf6jt8pG0EKqehFs7DBKa37fy1ZvPAt5N8/bs+lvlWo5A
2KASomcCFhv8lBtbNmAYkbwlZjrOs0XyxdVyvdUK+kGTNbYXbumECe/XXQO4pjNS
EvFCGOZG+1EtahL/arWhUchuH91jcGmfShAUa4Cx3t2OUXtPpuEbkaWz4ePkVvF0
EgcNU9nwZuJyq+H263hY536aZBkkO5bgfghl+zNk+FMi448h0JZV4CgyqXxRq9h8
fdPNhx4oM9Ko/yhkfre+nmf7ziy07UnlSQZmg4XrSPpts3BeBC/YOcC3uAd5rHt4
yNoMZ4IbilZ9kj2pui5EcF8VfhYDvQyHvidev+UJ/4xcdrLvgagQAam6kM1tHUTE
ULcOOq8dwrvMxc+we7FNnTdHxeVDFY0anykLqopO31kBBnZ9j5tGxsLGiCj4crff
oTMamET/3jnOSdd34xmnu/UhIlQmJe65yI53+oqNpkCGGo9WLNVRT9UZ07kGaMQT
zqpvuzVV1z7n7bBukK9B52315nfJNRJm63mjs/bJQcobBPfCSSokXldteTj99lPO
SvaO1r4kTUDtEgyWewZ4TeHSyQpvQJugvsv2Qc08jUFR5Vl/xV9gvd7Nj+SmuGcC
qYSDzM/HJnuDR1g0cRyzYxA4OHoMpcSybKHcqoPFVBkzjTgFXAV1HcE326geCCpA
JEkmSHy/Ago6TeZFdJNqyfRK15Mhtxg3rYMw7fydff9iXjM9Re5+qkHuNg/ZjKEt
9akOBiy20h0Lktg9x2WFaCP97P088Ofg+CSLfJqAwExLYayK/fW4hz3q7IIFIgQf
gQ8vSUN5HK2nrLcTRI5j80Qf/ZhAtAxzS/rXaogKZX4REI83rt2KYGq1MAETM8nS
66bGnrjEYS4gUxiAwcpBHOYv4RonpivjtI0KlnUS3IVLLC8Y+c3M+C+4xvwNWvEj
k38al4wVc9vdrQpKt3qX8iMHEoItIeN03+Cle2YGLpEcTAZqg2A0jsHeVpeFhDiP
LN25RzyCUocWIRJGlyXA8ZQryPctFXpXhGe24bXBWoi3hPaqmesKe4L4B9NJqwsc
gCoE0G9D2jytMPtQ1PGzSo5bxVrXjY86lOWfUiuZCZKK29gBsMp+KvPKnMzq9tLn
AXVVR3bytN76Q0jamaDsfyxGl+q8D2MQXqI80j73tEXKhwdaJW9T1OXTw72yC9qu
Zr33IIfbCpibdlUNT/dj81oquLnUnPErSjvjibqpt1QK8Qza+9qOrpb9qE4YPBPs
NSCp7n5ChbDlVRWJLNFxJdk+fpzvh/nWqjIzd408Kjsdoi5qWOYVhu89ixqwbNes
Je51pfMIYErXqnj3iFwQJzoVnP9NDh0OKqqE9V8OE1I3Aqy5eT7p2tcAMf8tF47Q
zEf5acpxvVPwX/Rr99y70kwhnYj8YgxTrMUw0gQ8nyXrW1DlnWg1WaY77oZ4qFIB
FtFcnjj0vFHWT4VnFDNSs5tbpAtTfei98IynfBPQFZY1kKs/0SCgIx+EGvuAdZ7h
+nlkSNOLGPR2mjtMn5Lo4T/KogYk96DfktuH38pLZTv6kwSqVwYcS1TNP8BJLM3o
IGgCwNOLdDKAyKJAxxue97Qr9is4Mq9ryJ3WOASxhPpsx5iaTwEpFt8IyR6mc1IV
tqA5U4O8nb89drpqnkCYPanHs+YgyMeZWXqZhAE6axcye8MSKOjsAyawYgbN1G+d
EMTb/8spBb/COWRmkv3wO7d+oA8iNZ0a6hTcd6MJK6E88Zv0m5SidK+p6BmR0aVX
JHvBqHhNaPwGWaCJdTkkhKqnXaONBq3PXTDXOYGYhjT5h6vV2e/E+isW345unvAj
jxaNE6jFe62t7KGMnMpYG5a+AQo1SqtAUChayAr2bSeCWjukhxIvkGnWyZl/VEp1
+E1SKpyvcc1Ezp1O8guzInj4DMg+UimkDu3Bf7Km+iLOytyb4afXP3UHwuHZWCDE
MVRmjjdiURddecBpurNRHZvz9rz+OKuPE8bd7AACzKsfVlt5zCCUl4NdHLpBYfWK
kzX88MyxIoOntoS28Ijj7S0T+YIOWSBUyxhUzhyMKHBCRCERBIZqpQMGW6GDnuML
x7t8Wza5GAx7XvBboQYHH1TWRE9jmXUPF+FD2NAlNu4OVHkE2m8B9iX8b5kH1IHY
SLU7o1w9++YIGuEe8g4NpyjmncwEl+X9+CuWwkTOKu8fSsxuIMMkIucUEUpsCcDT
bcmRWgoKdfMN0tDtx7jP3sB13REc4lEGoqgtxZPQ+jN2k4WySYJntzx2mwPobeVP
1YN+CtrVc09RFrZ8rAHHP9KV/qXUQyPFwdUgCa6cUXlG4EsOrRTdfbArROfGU5PR
Bhj/MayzkLbWTpnis28eUP0dU2xGOFZD6sCJ7oqLtjUJ22tTn1xsU3cIhRgrdarg
I9Zvvm4Q/WHbxVlenDqJncx02rq95sL+FiLSkDYCX2konLcGYScsIrPxNxvKQRqG
ftyPvB/Y/GUkvVT8FoV9H4mQt+Go70mc5XK5qzq9eU8bxtJhBqdl+WKU5cMt7baz
Ldvi5QfkeGnfuCEPkeFRoTUm2dZObm3LlRmp3PN8qOVIBCE4eP0zVcJ7lcJudJJt
OpsYemixCudPY2JKjIAaHIV8hoydMldr9KEo4Ptr9SnKrWYP2VAW8NwIAJP25xjO
9UkPK2X+uch2Esu40DMBqFSxeyPMr7/ACEOF4MG5ovD6VYM7irbwPTVWhHKqmRYD
2+XwT7hHh1wtokoWL+ePglaZ5ku1QNx4oOGhMEb0+MdiFp1hhFI7gdU11a58sRij
IOwtak4SfP//h4qHTfPWPfuoUnQUFGhM0zTNxoC+KwSkevcrt0YCd+iM31lI3S+u
bl7YRORb77OYElaIkhtVTvkj/iw0yWx5X4X5SXH7QuhxOyOGa+mwI7117RQsCvuv
5aDjzFNlu1vLE+6VTZ++V6POHlgefnknHjF+RjtLRRb+paT9s+wSEvQBFvv1PONw
7pXUzg3EbkZCL4Uc60NxD41+xNrQcgfFkBSLQfDBQ/SB66cUpRjhMgL7AHfMG+xO
xqvb1/Q4b/CYZM/y+oYlfsCBDuSZ/XbLfm3/ad62mozTgVkSRdZPJK93ktv53CjX
pogiYTUn2Cu9VYC4/79b/5LvGyk74mMkDdfEeEH8Ah1FjPb/pasSP+n/w7hSrcwq
n325wFuM0RJF9zbQ0IYJdPkNM+4BYqJvnv8HTO6GWmwLOsLwFhDQbnZYrjcKRhb6
5NvBB2yRJzWkvmlwzBtDf7hMmBXtjNqm8nqii9X9zq8XeAWaWMaLino0p9dsqtxM
VOId3spG1gd/jVe+6LXuQga1Nk9geiOUh3RxqgjvaYbSbL+goo5HF42J6fQPqiux
1OQIUzS0OrUcLJX60jBZCxv17H7T73m/yPADi9ELpg/XjMFeSVdDLl+/uXi2efTk
2cS7oNIA0G16/DAqws3yFkPkI5cBADP15bL/RjpaV3cqPP4e8iZEF/Y83PW9bHDU
npaZ46w/c6/P9EDz6p9qUPNK8VVqBDzBFU/bPa0oru+FPekMXwKXvB087UIpRQm6
k8izF1QaDV+gl+rBNz9dzvJhR8xPrmflO1m3JMCHdU9uiVwG8bzMJeJW8Oi4yBBu
oV0buDx97oCJLGKUaE9JykUwNI5qoflaPS6YVt8lGCa2yUPm269UQr7n9u6l8uC+
Kt/+NpTdOY2/DjXaE1o2fQq795gbY94RQk8JsXlahtPlij9NzALKEMsoR1QFBFFl
bLEgVX6RTVj2UkcFD241ZmGSLORC0RU9wnQO95FNoyCF2GGargoDm7vZe52S5SjN
QIRxR6NR2l3/1XekXoCNY4WywaaZC7W+KIuOHZP6t2IHa/cfcmtBZzr5ZSU8xS1h
rcYbXRdTLtfOsGdZat03LzK4sS8Rfns+ma9oV6w0M+VxFmLXnPlut92jBbluiBPs
qP04M0VPqPur67PRhuZ8xQy/jgKIsxRmTiILM9HsdAevyyTUdw1h5VzDr2yyXPbV
i2knXg1qtSgXxk+c/tFVS7LU7eGb7rxUair7R4n5A3gBE/XNQIVV1txp2mGrMs8I
uToxPd/0dq2Q6q7xCuB8WKelLYPiZ3dHYxWPk49zO8SX687O5mwLE+qRGukypKUA
oY9zy4/plvbCam3pO75GSpgqGSM/onLYnekGKgf0+3XYSQG0g3rX/XqurpwLpdVS
rRMQ7565ICiwjMW3yVNgFqZem2F/7I3dEpN/rQCIA48IjRDKwgVl+CHP4NykL6wV
YaVl1TAI6d4K4Szh2ST0qKtbaqCThpJje0c/RnWQgCG+2HQEMaQG4b8WXf5aCILc
WTZhA5FwI4UwkNoIzdCKV4v/GcSPLY0dHWJLTwH82kSlJUTjg6Q9CZmdb86IkvDM
l71pK5uzZQDdhNDeA3mwL0qZmdq5IyUBE7go6R/v+gQIyNIoV7+TB/qABBBQJocu
A5XexEhHt03cyvLSGaGZT2ZX8d89ClAOkFq9ndqbKlIID3TynduKRdfrXt/NVgUt
vyDbHFB8aQGhQp0VWK45td2/MwIs0HzqLoiPCLr2nDFOeJXJ9PpcR/9zbZUclTYP
/+6GoltLuPFtVP42GHVkA1yN+O8ll+2B9n5L0t4MJ2vU+6aqyf8boGb3U+Fd6ot1
4eTs2nrUtD4uYCyhtflxMx1HLXqulGRGkgc+pNKtOwKNOoPnkogAmBOKfEkuTTWW
ye735GKg6tYmLUXVWXdjDZj6g4iS7Nmiu4GIJF45jKNXdK9E8ZMzo1HGbrzKb+4e
yd7WDCTphFm4/jt92ZvQXXDlKRNWhjdxoYtNeRtkeI5Mhi52avmSaLsd8n3e1dCN
CUAH92Rmrn5y4FeVwW/zZmbODWg9gKy02c6hNJbLRQndk8EhNb/lgETe3SgqRtXN
2wnwXDN9xFweGMn5ecnkB76W7LD6DzrtStUEbnBrMA/wgvSeCJjqOA2C5f85hokm
m1Ni2iAqraAFRXOprfDjVer50+f2K0H4qZDoDED6H/3ippPnMJxrtWsjBRvU54TG
WnomtTG+XDSI03IcvooUYztNhm7rhUoTXeMBNrV6DRU4RuVRTFHi7Xwl+sHC0a0L
/NgeR6oFqIHWXxyNMho8Qw6q5zKTKAbO6ed7tJVesIe6wo9ofOacDl2lD2jF0JVU
XrI0vKE9S5BG3WoJ8N84klfzmA0++lpWlRC4o/3nZbRLJ4DwOldIrKcOrMW4sxCK
2JMa5FoappR0aaE3a+F/FcRnHbl7bDnHAflubEDMX5cfNruLfE9pTI/JUvQ1sMDN
4moxxEj0mE5x1+tWhR3YY/1qAGJe6088ZICP+NFgpMPjCsbPIa3RQIVebKFcHDOu
0wsXHRTILzO3nx4XG3/HQUv5BcJy7oa0FKf6gVyfc+F3BoohlSih43iire9oMqw3
DtFyDhiuM4OM1w7vXvQdUkTBvScvwZk4FRzXAA3EOeiu7WcDnuhtZW7+YQNri7VX
4z2YoVfjdqV4JXDqcNN74blFCBnsPIw1JyAXyzbOmUqIanPvc+KeFvEIiZ5UW5ZM
MbvSwTPZgii+IqFMPMV6e1BYL+siScmRD/nW0LGEDrTjEQ7hocXOqP36B3gsjrOo
6khJTm3sszM6VcVd7tW4eLs8CT4aebVMpk+930s4KAsUK86ZRAghA7aNyH0yKgRP
dzEDLbNbcLk0RBlii0HfEoBprtE01ve8ifDxoFJIUIFHgcAlA1JDv5b5elOBbMLQ
FWoONREfLftISdCAlQ9NP/kbaGB7VII+3g48X3v7EpZw+zLMWiCh8fxY9mT4/rc5
MPJ2Bu8LH7dBos0J7rUcqU38FOzaynlFufEeoi80Lt6vQKSx68rMOCXMgwsa/6+g
Y4IoKVjieHwyb921vc1SP/PtDnaIwLXt0+1I8HAnccOre6Yj7TKE8LT+MbAc31sk
6G9jsZcn3RVsbP8avd4HGzBQjm7RtbPvNMxDuC80nT/JpQbfNIqhEOT7NDLKb76g
exrmxJx+ADtgK1q04DmLPjMg4q4im/Nkwqx1tb1j7WXZAJ7d6WWiiw5hrLqjGq6n
ww3rD1xfy4Xt5JkIUvcPuFx6yoDdoivYu9yF9TgKGPH/b2e1goN8SZFXsky1yDO8
FHQihoaJ2nJAhA6fDPfYTSlK4Z4QKV1Cq5e7Tva6msONHC1SKxnngTgdqpaKhyGH
9r9hVxKIUaY/BipkjImWcGRS4uWa2xues/9LP9OmktVuLEHBD4FMaJbDe4ZKZoPM
sqDB2qPurl5gseim92oLGj0BkX/1ux2q2mk0RKLvBM8Y7c4yazdPigADdgpHhJHF
dA9IxCL9kEnSMyN/RUaHEbLWuHMZTijjJxJb3xYdUNCkNr7hdwpGfQrIiXEY9zrI
W6RoqEP4OaVcZMaqMypkBWCYFgxznmSh+9QCYjbhiGFjm+FlkwylEeZQirF+utJZ
0TDpytRymC89dPHRJcKGIku8Fx6LEs17s+k05vz3dpYYV18fVAXDwnGNF9OMItGR
Nz4O2WBktKAKoVtaOW8tfKYJjD8B8CVpI4fzdTY8XqoWxO46Tdk+YmVe23DgpPSA
NnIs6djzSMDAT/3zOGi6lF22SdBtaxR+b5C8S9/6BJvNGJWASMyUVcSlwLOmC+24
o9OGNtqGWShI8buIklwV5wThRbR5+XEOv1ta5diQThUUpq56WPir6nx6vciDJSb3
Sd+IglpAzvxVch8POyNOnWshU9vVyeH/Pnz2fGVbTVS5LG+1kk5Dj1pzei0QhDXl
rkG8/FGgUbzW8G3X6V6Jd7yRq7XByBA0I4jP5+DkUgsRlnzYQrb2GuwS4bmfrjfj
jeqHwO7zZV3XW1729kfwtRYQ43P8HOMVZ/33J7MikT6ahEgoKkqGR5I1CDzkPfTm
9etmMCUXmmKmhRRBYZZdtB/7Z6GMhCE4cYXjclPMm8PFF5wMT3Q9zwNWfOUj5zyX
thA5n4Wx0b/LzQ/yRuL+T3LMiVo7tKFZ69eGc7nW/YfkIpAp7Pjd/TeVXMZqRWPE
7mzz+hLB85/1joOfrPnJ/IdB87Sw6c236Q+Nt/WM0lO9q7tHErYelqIatNFszFJ9
TlALUcahSGGdYWFMbRFWOvR8ayUPalOeQ9dIR9QvstPRn2vTjNYBpTrq+r1eOv4G
8Scwb4YI6uDPCQu9mU8nWYSgckTEIivAHTD6oD+VvNC/v/o12MXOE4IBKywbbf3c
Z2Nvyp5O3EJvI8kMJm0Igky1qQ+/ygKyy8g+mud/GhHUiv/SEOUePcDXkXo2IuD2
cXqZK/gAO6plyItcu//7DMB2CyqiP1+9awfWfNx/zPc5op4Qgl+DJg54T4ebqKlA
/KaMcv/6TvoZ1pDx5nr3QACGIwd3S3Hpj8Iick2Od1+FlCQF9SWXQeL855AF5iwk
omk2GwTf+O5octi5KuYMkuwJRZFYC7uXEo0KrAtdrz4lJ34BBEYe9di1m6EgH/pr
RHfB7AQnb/2FrLoaCsSLJlZ6BJufkmZ3a1FnBOwqdKLgQOdGZFOzn18tylPBI0ff
rM+2DXts4Jvr1hDSklIAg9SISLkra4CCDJlOnJrVc8dS5R3OTgC16kQ5X2kUc24P
Ee986okHmIadgvWpypA3VaZBNQSEJJUssL36Fj3D0m1C27SvhyFlAzLKq2a/jvH6
Ba68nI9/llwhdPU453Cfb9pFJa6aFfTJ3JFhzWTguqSREYx2Y2fRq6FY9gXLUJPa
FOaW9bjlV6fKs7gUPy7ABHPnusmqM2HatXLctd6R6DC5izzEC8DwlXod6TxT5L0Z
k75nUdgeE41vtti4HoKAq3G0KwSHNLDyJlNIJxKy4m53tQXJhSKiUwtxcNrKyenG
wUJm7nz+t8WDKjxRLroCtuTxhmK4GsnUXx1KRZvP4PJUV3uZGmBBkexGj7BbSXZe
LPb1L22raU7gMciz7zWk6D52+E/aq+pVAwUYXndzijU6sE2wP4QlcDWKVFguRkBk
EsoDU6+3uJ/ZZfH1aFq7mTit9gp/8MvEmNu50BcqT+2umq3h5BzivjJ54Od3J+1Q
0RnHV3Em4YHx8Y+tw5Ivxog9xhCiMdP128OGyNDXvBJkJCqmAkJ0gYmMQHu2blEK
+f3Q6p5rQcmqKnld/q13XX85euVUFGXgESa5JkkrIuWY+cC/QaYz//aVUSRwSEOe
Hnaa1NLV3Ne1QtKKev8D5+SqLEsQmcaEUOt8fflmUua2xdJkPdd/DrKT8tPGiGqX
eNZyM+95GkdYWzJuW/9f/DQVbCEc0ArJ+q+VrOLS1E2caMepcmyOPzroBjuK5YT8
O5HvdJj8G4ftSDQg6lC+vprwc4Gj8BpxLIHqczlzMl4J6aHughXVuZLaFK1KfF43
dsUwh4THuo7OYwBfHM3KZyJ5qQCv1/3x7CXcPbzyZRkBakF7YL++bvS+237ub5OM
VptIEoF/X9fQdkAgrirHdtmj+h8uq5UOfJtFBO1JIeBNprmb2HNa464bXwPPXVmE
iv4Y7XiMNLy0CG8ElG7ep9inObJ0r4+2cdGBZXdSGeciY/OIGYFdLuCG+AT3Y18F
uxp+yAQ/lHdpgVd9gVbifkDsKIMsziFzDYsUaPxl54zku4BWoFPT1/FuCa78YOSm
jpUm51Nzr1c1BF4abArU5PL+fRdbc+syvBfzYSeDdM5cYCyXjzfQ7JqASReeLkYe
2uWs7t00X+nEm2wn0I/DIjRI2GWfqA5MgdElwclBh5JA7pKQQGAEXW36FXQPT/ck
mjvupdl4iHtP0M8drNrL1s46ZBYYVX38t5CYtk8sCejZ9Wpf00MOaHLuv3qgCsfJ
iSzkzSHBT8qwpmMI2SLyxiWq+hT682jpDRza1n28QdyY2FjHPIlZa+0/tyhmY037
adLx0exnKDybtM0B0c/QDOEx5lvUK7ca0NbepWboCe3gDqXtwlW3ZZLlf7+uZxpE
YFMGrVXYFIP43+Lt3yc7y9E8bQza922CCAVaAziE6JMCgX/+GRkL64LVYugNaRjL
RJgD9b58kor2dtzq7pQJbR9/+TUayYNwyJs2P3XpCkOCo9dlu5tj4ofl/AIczVhp
B+4sl0H8UlNtp0JxarkfF8TXCQKmId7dkKt97FNf8FsDmXuCbZEn8gQ61Fux/6f4
6lH3TIuXIuwaxquxJmxdN/ygEckyCW26BDv9R4UTdkoDfq4q6s1NiRPCJUs06UH+
WOsCHMosL/OrD9oNIIOhTycVompeSscBHfDZwAW1egxUTA0JoWK1y8gHHvzaPIAn
GGSpXdB3eoja7XVSUjEwe2O363qhmix0WSYGmMP5OUXo9lna9OaWjH8RnWTcLdVe
y/0YJ9tcGTOUXZf6Kogck9YWfIqAKJXVzZjiVQaTpQfsQk5oPw1dI20RDVwGUx4X
a+ibQg2y35XvN21HVXS/XTo8B3I3ykjjltcPHJjFvbuQ88gxMo484tiiFtPn2WnB
N+Vibqpw/QHRaLXmC6ZP3dtICqGpPFUI8b1E0o2SZTasRDWTlMqOsrigOnzwB1kw
Gl0OdbwgK0BJWK5BkFvMsvk2CeyqTB4x7XImaxl5ZToWIUiJ9fzom+01mEFiuoms
WyrMoy+e9W8T+vxyZTsNm7CfRutKT8tzUJc8P0sEzHfjiShxHXWRyGiP2MN16stP
oDGbGEqwOkof3nqUpLoQQKH9ASZXLGhuMKjAsOiZPl6i4Y175C4TQE+SXJy4KLFO
Nt3Qmyo2PjFYrvnrijB2CR04ILY/B1u4vv6S3mHVm05zf44QQwkhi6Ex2YQ4HqYK
ml8957M9e3IRqttZ1V8SqWhF3/FoXV99ef1knEIHZGz790hHMuqS/eXL53IoKKyW
vY//lOPhd+/oMzczaBnMIclBoBFeqGurrPcRGQ/df+2gixTwmU0goooMc8r5ciUN
UyacuMbLB8DAl5Sa3H8xhbqnd2uQktVQhLwoTYe7FcmeRmmKlgW/I/u3jN+30I6L
r/PGlUdLFMJEXSrBgZ8Vo5KCiefK+OJt5fG8NVFoqJrfZivYboivuv09eBQv/Zp4
kpXEwoN8Wa+EVsaMA3b5NwJcdjjquaYJJNwyiHnpd9aBUNy7PSkNLbhiL+E+hFVd
iBQlZogX4dehBx8lAkYZl+6xvkkdSy4KJWK2NIuJIaK4oqLDwKscBJor+qgfeBO/
MhrIUXneVKAQL0zgQlP5ncbrQx8S/6LZijSOhJkMiU0qGg0Yag/sUsNDT+ttIrpD
PVfbpqH6MGM+xbFDwXYE6Lk9JVmS8zKPZ07GHPAO5WmJK3hDKM/mTX3nE6JFSeMS
nsre5/RNb5284C94eyLHwxOGD1Zn3FvfeXDX6mol66n5gTk1dX2JdDtURIdASieO
csg2/3o3Mu4k3yDzxjwmKBAT9qtta8lDxLipj2wHx6obbTQ7x4ho9cUDKXQg3dEv
2D0BbTwK95fe1tYpJMsY9e7G8BndTLD8lTTvGK6pLUoiutfiXkWm/NdMIn4MpriF
kXGxncpYIrky3cfN0ggmrbIU22eLq5PNZHWbZm+YAM/UkTDutB9JjxRAEhNsv4pK
i1SxCgXb57ZondVy9R3uZAISt5qS+xSTbIOfwfDr0Whp7H44BITaEjZ9H0X4lryD
WzGWLm+5UHC4qL0t27usQ9qMw1BKB8SlUL11zschuWkXxQu5iM6C2A/CBIJO48Ea
ZrGPQNUdf3FsmJL9CGg2Rg814xHYo0hCDtrrUC3n+7Y0n2EszYOOWeB53JJDbWM+
+xntWdYyeecgSrKgkTHrUnFOtl0DmgzgOtwcWObG2paw0tZslbe+L9TwSMjBJb9K
CDDQHmYybqT067Vpw4ZYIPTAJTSYYM1RLFUqb54VDZNA3miBMNLGTJAGwf5ERfdy
SEjwKKLLnWbkXDMwPpU6tUglYJLrs+Fh9EUgjohHZf/IGVZPqc2OGcDuzmkQ0WIk
D49EmuytWUp9L1JRD5qbWj0REUpKpfhTb1hM6DWULjWcQd/U27xYHjgQsGXSZ57o
LAs2Ddvlb0h6dRouXUwzUIsbunjgDzZ9VKKNFRPrH87OhsiF08Hy2Q4JJHIxiEW9
nTMCtRr2t3r8Pvmv8MvOO35d/bLWgIX1eUhPCTxvvS98Sz6fNeUhd3UEQTYDWNDE
DmurK4wMPOmDL02zF0L4KV2XLCKq9zCgNS+wKFcXiIXbQTtXY6N7bPiBd2ELx09F
8ZCo94MgglmR6GBVo3Wth9OiLXGKXtpSAyhtlA4lD459/Mhao1Gn3WBrgaX5i+Ug
tqLuMK0Ls6qh9IxKQtC3f3psE/NbgCzTAueCRwLpUA1XrIekXXFGxcbiYgstRDs6
oXhPuwIpGjmPeLx0BzS5oGHLyqOof/B5dYWiALMH+pB8pvBPQBIL6Aax8vD0DZAS
Ku8FItuo/sONMzY0aCd19ZCmm9zo76PS5HZMonB01/adSblrSx6VB2Neu+WgGu2s
c7XWq2WFrsUgnHY+GJp8WcGQJh68cFXv0vzL4Vzv392eWPtyio8ILnYL/tzZqnOb
pbrbF871oTF0IqhM3ouBPqzw3zU8i5SeU9iud0livJGZmmyp3wZ70E54OQBZv+KP
zJ1jy1p/vuXHNNJsg6mWooyBFyj0d1S9tZ/queb894CXWh6gv8uIZWDaJnlAMZUr
WT75uGkJ/C45TKvPJ/53bv3wpuNLM+Ap9jjmEEvIOynrJePGMMcvqFh/29mr4bQ/
aqa1DNikeYTg9yeGRx9JVXI281deJWei3GKjpdVIHsIVwZQU3uF+hATwF49xLsVj
AR69Cs07/MLBKsfhYNAuKozZUceSE2wOIDqNCLa12ZfWnhBNZCoAGMIk7QpMDaPe
LFpHoRzvHcht3deFZLzBdZ+31XJsNoIPzPpjdhtTWksIN8JOUTQr0T9Lk6kA9du4
81U1+ITiXrFmjCsUVwgJlfg+GSMIoKE1vFjEyYsgxja47LW2VQl1axGY8V07iSw3
vWBPgxs5dy/Xk+ggSHmfG/lTvSmpUqGl//Y3wwserxyxHCv54NBTynXv+yyZJnsh
ZzJTeNXX9dkKDl73ocF0U9fD6YEdd1YTOiiV8TFgGRMecn2+hEKc6qbmxLGEIAWT
ghwtPnXC1i4hSbew0PhJTSRNEY537sBfSeVikfkzdDrN6GtpLQjohoukeK1annww
d6rJheTqgr7iff4J0qj6ie/77ITOE83/J12m29rluUZyBIreJyiDYh9sxtWSKvj1
5cYA62SAPB0g80F+ivUilnq+PQkS5YEfvtPPWCHcP8g5w1jrnDSoNdPFiH/uKIvZ
PIygjDgTFG2PbrUYOYXN1WOlnWxwIcn/wQ9D42k31O0HPGdB/pkQV82JXNb+xaCJ
xO04KfqJdA9grsuTNs3bpi2aB4BOgBOkH8Sx4DfpN+NQTeWt4+3A3z5f8yaOJIEY
Tfg1gmMC0EuWGSq86OE3dBkFO3jS7BulNCjDFHkc4PwLLYPqJIHaTJbi6/IRPKu8
5UOXTQr+fvv8JWrarllFqB+JvYdiX/zg/X+cMPzS7k9xshfRTC5fNHvM25eUN4SK
gPhyjH3K+vr5zhx/uFxdh60//YeUBmzDxy32ZyCLZVWfatyI2YusRQHdtc019jE7
bgcufc/bBmOZ41Ybodm8nUmf7Zn4/HjRMKU89LxwL+4lH8MtWMaPFQYoQ8ua73YM
vtNARhW3ItJ8zcwCfrImv/RNi8hp9uinICZCZSMIdWtno2SLgz55pMXyov917BgL
Pzro4aB/VlbPIM2yXfxvB7gmXaudTaN8UWOJeTvNd8RKfYZQx03Uiy1ZsBSWS7RY
s0zTrJgYDMTfUIkvnUubckgi3Z89yp8w1k3B1t2wWa3/zmAmobjbAPUHud0D4juh
8MtrfOTUR4GNfUtpZIdbCa86Rq59Owg6LN49H9237BpkyjOkf8ET4TX439GysQix
UW0BaclgLYRDxlW5eBfV9YF8TvxD3J2e4WUBPJ8WzJ700Muaqw1BhdriypiIhCxK
1Xur+zwq5PhrgZKrUuiEL5gQCoVrHg2gal8+gYhwpYMvoRlk/NZoTe0lSAk5U/OB
HNArxF0sdifE9OUE4carvU/EAKHTvnlpE9eck1wfjQpVtsnDSNsvFCekG88On9t1
Bo+hibR9pVg2GqGuWkniY6NN1enk6d0MM8fLjrcp3soKqAu4sYrSdv8bGrUR9W4N
AOooez48uzHxc+7zeer9Qu1SOFtC2q3wJdsWx00EdWJlG2qEWHBuvZbjmUsfITnm
aGFXphrEa2M0CQlLmEZxtlUIeWZbAD3ZHL6UJLFgL2QPZ6ZUDFA/Jo2kjijY/28f
5GOx91yEHTlTbIaoAf6upAvhfmnYsjDKRQ4AYCd1sbHHZROJkZ8pyFUFqPbKdLm+
ieu9b/Tw1XUJSyI96oC8VTW7a5zeElBMNKcAULVRaPRh8rFfW7Rkmft5bKcOugzH
YspmrsBwU2gxSufMlMwPKxST0I5br8wAvh2ad3Q48QVdJ/Sq8FDaKsCn+izBufel
eDqGVFWcds5ds6C6U0UcaE5+0SkSZxGTgfYsOFKtTr89jPR5be7GfEtLjBgh7ZJD
Jj1MrAN6LWMLKlZqoPvovviKSBGWnwRgmRNyBN3jki3/nVAeiAysNz0FIV97BY3S
YyDehUkcPc2/I+DxOK6Cu6Lz5qhFZFc0KbeddWvor+LIHyGe7xlvuPO8CKRrMyWE
mwjfZmdVHQ+iBE/25b1ObW9NSzYN1o6oOdzCy2U7F5sXM8+G/wGKcSnQXB1HINFj
BE94wIbRdWpESk8Mb9fUN5d5ChPKeQ+8OlAL3BpcVVmVhV85R5O+pGUhomGGXYgf
hYXqnS4oogl5hSnPuTyq7hveVlNCqCp+fM+AL0VdGeDwbUmLcHCfUMnjQcZp2Q7I
KzRAWE7FeX1QVDrraV1sSSUFheNedz58etDyM/0O0LC/uC4pOhQ3HH7IS9hoL42A
e7p2QcoH/vHh4ppDWH4KQQr4ijfUC1a0qNoKgihD9NjyD93naGX2T+a/t+N5DmWs
jVdOio+mm1iEdoiTLOpVv/rrAk1rQSyFY8pdW7NB13PbmDtxMjtWxzgMtY84IhS2
dzAKGKkTqPtJlIAxOfC1DfnY1S8TQyPRL1dNv+k1GH9u5xEcAhUbmNxwhseLRQyQ
6N0gMu6go0vQ8T3MFJNeQpW4PsrIIfxxGMxOTRcPyDS0zCa+9pF7zJpb4GJ/rXhv
WPqxZADgWc0fmWTvU6/paaYEosI9PwWAOer+KS3XuOCMpMAGrCMgyK7PeEcizncc
X63i0NA6Fv9lE7AzfgWvz1l4ZJsUwDBxcWZZd3/OU5ymQFahPRcevHkOFsCBsaz8
DSJBwVnDQ+8d+KAEeJp7N6xtAYE6rFzryUi6VtV/xMHwDC5djNRDbtRMeJi6GSeH
1J5lEYxYkw/KbqLJVajC2aKh8+LvBQxbAK3Xqujelc6b2N+mJLCdT9I/AJ8DJqab
RdliLlH/VDHQFzsReqNC15yCRyWehTUKIFVgzaeRmJCPqdHrjjp35lcx1T//H5UH
9wHQGZm/kWA0xEfts3DUdwrPdQein8vAr+KIL8Be4KDmKKXtt7jBd81uAPHmJKfV
UoY6yRDuk30ey3/bVYAlRfu6VvfxJxgf/YJ7exoo4MVL/kcxZfcUXcbI/BXsvzYJ
R3zj6nnMR3WytUX0OmokyVr3YK4ZzDwf9J6b4g/qui4XcsynvP8jl+gs/l1KTHEP
LZPy/h7QT8nsLR7ch52uCKYC2ZN7MnC+OUkccRSUcJeCEPc8Xm8A5XiGdcjJxuUe
Ds38kUwrpg3B3bxd4kikWqO1dkJM4x9cYx2bhSkIRL3Od82Bzzy6si/pFkNgagip
KiL5gR9K+xLsTjsUbdggh8o8RV0yygPwdKc2gOL5/q0vVoBgsRosrPGYmgqbkaub
IpDG75PFv+3o09gSSkgpKZCP74w2MUcMY66H9IZqBAuLq1U3E96c1wwJDWW4iN0s
21ZCMdjlRSFZ4a4ycEd02LHenDWQ22FVYwISy06Va3mbjTH/Q5WTv57upInKxKF2
iZ1UB0bJPKcruZ50PA0A72NRQeTqrBkvihuc+agGWPkueVfwCzYcl0ZpNDPmK4BU
vRueCIgOSYbrBvOXS/cg8SY9/4Ya+HgmNm1BnP7Y4RVYDEbyXhIAM8ZbGlFbqfCj
9gjtPBUpIYElcogijrH0H85vkCqDXxIEbmCQJsOdgFm56u0ur+C5plGgsvVe3T1i
wWQZCGjPfV3Y37WsncY5rKzi+ETFXCO7cLkOwL5YMtM59ucVaflexc0lYUF9LlAC
FNagtuvftZlSzNcMJ+ghYZvvNjAUy8f6wL2nIotGrAA18lXgCaFSuDvvUkU/7sz1
gyJ4X+N2TrxgwKRaIAqFnZwxR5J0TLbGzmZBOlq2fII5FLF11NG89f+p2fZT8c+O
8yM/OCuwm6yzX3uwgtfGTDmUKRLszVo9MSrHaLDFG+jJKw0Bp4gyPb4MXJF3vu6F
4s0OfvxtlNQy4l7eJCQOdLCFFOv6mJ7ZRWJlWjFxVviYJ3sr3uEuegq7iuUX/o+4
WVIhBpfjdM/hnGv8RFI5iPbJ0Y1XxnSpS21vYliX5a7SQVNSH4xKRsl3wQLKD23E
YuAe8LmxhUdieQxTcHE2OMGTbjtwP31VG9YcNOyTW/lVEacAK6FwaWld7QxMvKTo
tEQ0K5XS13zMPw6lvd7vFladDm30rm4yrYCP7Iq65hi3CBWNHAzorFUWQhrqY2Xi
+ZECReS4ER56GlU+cH2TWUo7+OpTqgCblVzR7fUZ009fm8vacmChposvPd4On/vn
efiVFFcazv0ww6onEe3wg5ygyDXaYyZnsMETk9FD+WYOMvSxodFNxTY06ISP52op
N2qGSLPPm9ylzi/oDhqe6CUij7QR79j+nCBNOVjwR/GlBNy5lldam+2cY27qV5mV
ldeOpdqoznyiQupqTYf/k+eAXhf+CZoFDwSobCAT8NSthUgnjLS5QYHjyTlfU8yr
WcrOoj+fkSEvS93Kj4VlZlpcKGHwc9bewtb/LVtUIkHRAoD4M94eLGTpfvxplA6L
7j164crfHga7Gw7eAI1tiLcS2M4xdZCH8SRVRB/CQ7i0g0LqHeNpc1yQkNLNqO49
vFhcoapNLFXTe/uXkUCb+iCH6eSh8CnIhnSUJEaZ5njIwK1lUwybqKxPQ9rtjNCo
rZasRCqeqS16EA4wBTzIXkIkDHiMmy3hPdUCUCPIM0o1KUhOnue9Fzku5JUHgrSM
mXj7IV3giJoisan9n2dDYMzbl7YyQiZr6B01CpB/mJTdh9guY5AqXCsTYuowetUr
/XK/NTWGHsvXtKjquj3/jKtf2FpHPytV4Wn6RvsSxZs8Kniqbyr2G2IRiU7HjDN9
MOp2cgni8wEshCzMVFPXJ4e5ejC0ZfWwhMwfi/ahUdG9WxVzmOCcvv9NXZqDnLEQ
1+Jx7r+nCc6BrsC42/jtqcHgIDsJt/T0LjmZvRhvoO2P6TQbTDtncahZSYppTPp+
z0K5BfxqdAyyb5bBsImnwpk4FJrPJSq6+1IOsY+fG+huVHCJ1e+FS4HJdm1PAnlE
V3NbaDokVjW2X6W5qm7l4xAqBtUzzO9ZYl4jUqNT3V/Vq+EMZKuGevuuQ8VLU3tr
0DyfLn8dQcusnG2fiIUywHwDLTBDDpFkOtUpS4n8iUOLaUtw3enZxDXqHwe04wzs
7tsGyxo0fsJxXW1jDpL+8Bmd65/37rYewtMeNEGHI1Tl6fv8a1kmMxpflghnM/6g
G47A9sASXcgCICzmyMThgE7DGbTPcyfg85pSDQoHxbQNYD3lbVYJx3b2FnK1i7xo
+PZxrcs4QKmVE1LcK/udfOs08Zcs+NIRfKn/LlqgIAkm0geWOxFLMTCNGVr+iR1Q
EXZbwvObq+oY8w3MYDqrLaslzpSICj4B1NLAn1QAVgGYVuvUcatXwpLTFzC24Uuz
uN87PzK722YmF1bBTLUzRyR8Qid5B6eWhj6nQhhns3Oz20JyHpA6F/boCsFUGFQ6
3baI9iTnrp4NUS2zgTRs5V1UhcG6xiax0R69LwZ9uv96UbM0VaXkDA5j740IXZZT
A5FkGN9zjo8nhtjLxVpuKvKMclloqw8BBnVzkOugU/wJppVZ7IH/YkTDK2u3wrB2
2K4FxfnTXPrdOXa7RA9zKOuACZyq5izepiW8W4ymBRbGRUD/lIXLMN/Umr19Nf0p
KaFvXbAk0AD1uoGJNd838tVgBQk1nHQqLGqCOVJxsh36fV1KazygwQaFeRpF400Y
VhkPXtboECw87vT+IIyqfKoKZC5NABRE6QyQZoIiDCboZCFkVCKPPtb176bFCvbv
IKGN9e3NMY7+P4YUcEsbci2ZVwy/Bp6X73AB8IX/o5d/WZ4kAWw+3clgwEYeL93X
R7yhYt5OrmlkADTGa3Lz+Sq2XaBmFK6HN9xsg8dw5T6br8BOcFsVkPwuObM6+IEj
edMbHsiS/lZAkxD+TIeBSX1QgeeNoA4xptZMAvYhG6rDHu75XVQtJ66mX3JO2nXI
9WV46A3hAdG/y635TlOme3cuul6uNcviBIf4myAwnrXxjTXjZuBmyTJF+Yjqr68R
K/iNZ3jvgSDA849QIdGB7S9zx/FU5FHfXNOhD4zXhGubrlerpZhh4I9TltkWudVV
LHObR/8n9BLhZzDMW93XuJzqC8Faxv1duhiK61G+gnCz1Nvgy+XaZjX63NHexUz/
W7Rpz+6S/oWszRzcx4aCPqsQOmOZSnWuy6A3r6rCkVW4FfqoP4wP+uTC42IQncLM
oXnzHELKNlPtLbpcpqbGvaoGisPukqIEzlOlKAHihb/NlgKM9mEIiKGAiR1n+LTd
dPK3PA/QeA1QW3dAoGNntrwr1hUS8AfLvE0O9i89i3nV0vj6hNDiGk2pNpAWyCQJ
BznrakSjCKr+8jhDAh3PwYsUy7vs1MJUqTNQ6BsEzg/U1pL3UkCM0nNTXqMu6dGP
hw1mwCSvRs2IljTquIxlsy/7lMlbZP3dsv+NW4mxZVcJrihMUXK+96qePyo77nv3
ByDE1Cx3lnb/JM8cCDrXODhY39Z/yD9Du3QHqf0dE+HwRusalIf97z8WsYDpeBhI
g+STW8uSx7Re06jpedzUaY7A2BseHIdq11vDNrop9iKUAXrs6Ryg34QQtsokYKlf
3oQehj0gszce26xjNeeIXhMMP6xOYQf9XzgYjCO0/xaaCaG95M7gvXS1BkoSihsQ
eD7AAnpCLytQv46xQniqj6kdvFeC4a7M64zs3iFqTdvqOSS/Y/7MdkLm9cDHECXz
iRMIPo89//IwF+MJCq37Xd64hkB/1A3GGMHDwrGKCqRKOMz+IK9hO+JvFPRGFR0d
oTz9oattnZbeDJjOKx35JObupXkw+JG2K7U0yf195vx7aVLX5Q+3IN5RcwkTjUR4
WRwUc+k3jhBw8jUpy5FvbnuLZhkzBuwHEhaboQAG1f2qhjEJndwax4dLkrCt8kt4
40wMxIOEb7RSSdrzzTRwVHCsGQLEuDE8qUSlzV8xRlxn8j5GcUaOrhjM1yPEkzfs
ja28rA0FwLyUak5vUTJ6NJO+svZ7A4dhyIRbsMK7tt334U6jsJe+rKk8hLfUrdg5
nh5TEcnMHBZIJeaaV/0zO/9z3jRZgy6g21xY1zdAPT0KF+PfY+hGbPLQAVthDx/k
mbd+VSw5iaSgQip81KcRcqqw2HIpI97OOl2VAizRDnUqP0DhmhOLXz30ynekyBth
KKGvZQ2JnhoptfT8gImjKPviNU0QsBnn/lBa/AbVvKRend4R7R26SnxYoLVWX2hg
3WtF9xdno1GSiXRMoV6kQAiMTeyFKgjhgW8AvUFRKfZyJgHv7yUe9LKl+Y+Xb0+L
PmiXTu27CLml5lRYVHzg9FMEsAtUILWr1uZUi0LnTdDsjXBhDI4E8zmQT7SyLFZp
zHNiYjTGn47SZAvTL/e262UpqpqsHEhIOa/CQz4VkmAGyaHTAEe6AhgAFOiakrTe
Woub7genlXiAJwR2SGbaiE6tXB30e+FyrppW9YH9jHfSWEGJJn9PVL4aMLFLRnH7
X4G7IkGWGUM1u7tj74h5GoOdiO/qRUx74vtmtPgzd6DL7W04/OJo7HO8xHLjjtCB
1zMqZ/IdISpuYMvfuTm+K89dqHId/hBvWdk34vQNHOBPzkZEUdeshHTMOGPCrAUO
ps727mjzTdOWnCfpRa3AeMkvVBnqCauGe6/yQa9NI9GAsQBywvYazZBEJXt0vI9/
bVqRPXTvvu1DD3Tm9z+x2uHHUEEwz2cdu7wKu2oRXQbHiV1XqLN0Oj2PpXd1mkpf
NRjUL8vJkiVzTxwMUWbG9rP79hOndOyDjOXq5LSXBgO7//UgVzfJsIsjCBf7h/ql
jAQFkBtA3+QHWx1N7ihTQlcbEGDNRAFav2rOH7DIeSGn7CR1TctJvZOeejQiWARK
pKhIHNepzxWsQqCLTi/+UItbchB4R8NrpZURkeZie0TrWSpSW/Zd9TobjGNAXleF
FHxnoVwUu2iyitemglGm94CRLPng9oaUYEuzqT7uBkGL+cqbM5Twfa6XKTVWWYpa
6BLluc4xIkvu39jRNP+nn1dCweJusfhOb+TxdTJkxMBDckdsiKLS5E5nZgHLnmg4
Zre6MGaCmcJxddU9Nzn1OwzgCd2IXz4SFPQDKVjd80W+XbZf5lo3CkgyMGA3pVOT
msAwWRIVoLI/gmva4t99Kcb/AgzYkLyFLTVQJYA76beHnBcGrmtnPkmvmp4fldX/
R/uwry50CmyWmVxZa8tMIK8V9L0RXTjnVsfckJpVGZeZQ48eU/7+J/5EFbHWCWvM
4H5LQV+aeqa18t5jr7jfdN1JLIbLca+iw+hAHFulMxQfmuqCCv8ujb0WyAvNhynj
4I7jg0HAd6Hav95UIKzB1zeJvXTBElxgVz6x1lKKRM8PUrFz8TLZHlZu2KuK3Vdq
8ryE8YfSbk2FCaP3jthtj2OBh32OXkbc48esc7imnFzFhnXlpwknoAET2I8t0fJ8
iafjFooENt6qu3tUDTttRzCKIquFG1JLhY7Dr4kQUI0IjCXzrDNKgIA2O72FyEhl
4JvmojtUrghRBvytl5+SM9nXo9CANxd+wkx4nQNt0tq6I+AVAbAQBM9JsvabH3Td
i8qF19IYlZ1TrLrLsaJ0+AjGXm+CoxMPmxBGnu7V/ln9RUHpiVJYNgfZoPCEz+v2
sNqU0wcPdoxIbFIz8Fb5YONwI49bOl+bJXi7p1IefsLB7xd4Ek5W5AwjLIna8EaS
7+WmVF7CU6RcRoaZEKJrnJ8Mr8MeD49Oe1YoqpsW+JXCI1vKVcjD966WiqI8dkfp
rvhU97JXEhY9dI6ari91dthdsORsluNHBKwpTDtyKuI2eM8R3YG7xMJmtKhEx17z
/CeaoW+Qm8t56Hdugk6oByXDDkyVvkK+QEAt89NgEuYSzY8TaQFRzTdzObJWzlAR
X30qXi/JcEhgEsJ3TDg3XWTlxtlgKDt7HHIZ5WDoTQ3fJzZLJkc1gDGsjxbE2sXW
myN8KQDj1tikjOwZ9EEBwZQ76DLbG7FgAjXzKSiHQMIdA1oLHZ0xEOOzZulAG9ZE
vfA/wBllZNSGBkrlLZ3CyHwVv26e6KZMZBO1zq2nzlJRJrrN6LjkeIDJMEQLTjOH
BGz36/bnbjSGU3a1JQNrMUGvsjkqmVMjeZ7LPR0cNg7Bbkus8/nYcreddfJw0D4n
LXOokH0QEDStrW7vGIpwCgagYQ7w/EgLc4jB2Eq6m1AWkWZID0rm9VPARfx0ZBu/
7cjTtnW5vtaRTnCPRyJ88OTOoslpPs1YS6XJlhnW7gjOy4JayEnJpcqsS//w7dNM
J4q/FbCWf1l4VAgRuIw5tauyDEHn7MDKtUouL0dbkRx19CO0yvn4YpvF/R84Fhon
wgDHibfUv2v+pw3kddXxjQgPfHDm6hb5FDPEtCL2w0Q9cmzNfbCp/XW7AQPKaXEE
zAHPcL8p1V4WJrUioYTaS3uMllyVja3JwnPPfUG0fpMPC8iBAtlumVmDc9RsDBj4
wJweQR2EuqakKP881XvZoP/ztxqKNI9eWkCuDoXmaeLIaPDgWA+xUvzho0sTJj2N
UREfDg9/zgpGf/krAugWUXsoM9/4mRCF+mRTJpdUo6E8Xr3YOQFKiwtgFV2YpBns
m+bMF+nXdKK/T74OV9F8NIWNR7oTYTqSZdsih748e4obDL9gX/kqKU8EkdRaTx2A
x40MPMSfRDs16s56SuSrLwMRzTfY5plaS/BeUcE868xlrFPqPqdivvvFJfZtvE4b
ZyRwjD4EleRkFSkbCR+pbsrydBPzf5YEnFx5dMhodoy6v1HipPumeL5Hr8Inzu/F
f1I7O2m+oXB6KiASpeuVtq+zyaQm/vrKnILn88xRsWiBLLooAzBaRal1B1sSg9uw
3YpBuO7MhIt3RN1MB08NqqiRRI7yaFyDid69dISFjxYqoSBnQWNERHLrEfHG4Lpq
ZSQD0Oqfg54Sbcl/bKJnqxOqbCdSZIKHLOLaRTjMRLhLjgtf8xudCjnOM5VF6VKd
Vmv8D3RCXi01SRPH8G23BczQTkZnwuR121boE4SUGSR6oTPidyLfaJRsiSS06ru+
tfjpPL9+/6ngODoruPMDQO5hsaQtLPXHAv0u6y+XV3xnxUkSkECn2iE71fYTrPYw
hMcDVRHpUqKuDnnM8O9iMVhwFgAH+obSzKsPyY4zNO/JPuF4U6IiAgWytTi2Fo00
W3pt7DjoYtZdcERQLm/MLvTeb+IzhZj827w54fKU855Fj0xJQqaGsQNzY4gM6qWJ
/7ZjjbT+WwvO2kzFdMxmvSWzVVhF8gNrZsnfimskT2bzmVkwrpZ9qn40EW1a1OGo
2aeR8JuNkQ3udrezegm6l0Ih1Yi0j/TGWcKRa1A0bn5dwmPkGjgSGhALuyNBU2l4
tjvsWr8lLijVsvjVySluIMjh1YwrSdb0N/J1aY2o8baE7kYTZUGM4PwLweQhM/aG
vFhtognxgGTT0sHDFD5OJ6X9+ZON8eQtrh9RP3s67kR/Pvj1U5d7BqhNAkeDLEnt
FRnehssPKdBBSoHIh97vvKD7pNap+4kbzm5vXqlRU/shm4qhbWBjarZWzFsLsTiZ
JnfIDQ6sPEW9x1OXlvMM+KA7mut3Y+rNS0jk+//Fc+MyJwArEEMhY4jJIbYirGxv
SGqc01Q+Cf78YioJE3cIeILmhSnkKgCiGRrlINiORCntgGIwoOUQaoYnPW/zTvgF
3vqeyXm2fayYWo8WYkcnaY6hMLeX69E8EN4wBEX7r2W4c1pbIOuIu21L39zUby84
mkwRQj6sAZWgYvQOgks1sSCjuMSHLaz2OrK5PlfXy/FLGC94XfI0fLUB7xMU4zq6
cvHkGrXgy40Ese8GoOjpY2Lr4OMh9/jhiaDU47k0EPM7MdqZ174D1syKIRirDjvY
oNb3aH7TaivrQkgp6lZdDTX/37/Vpch8BrxlFG6Dyyrg34NasfD1nqg39ZTStrdG
zyb87QmxRHSDeWVS3Dik1g/EyoojqqlGlT141+sk3ZiRPILSoNIYr9+nLK8MGI5T
JYsL9ekIbsATZOofBybNMl/9puJN54NNPNIp/AFHjo9jwU64etiwLveBRzHSyJLX
pmdk0XSEBfQ12OK80aV2yVHtfcNc63KE016kv0TlPu6Rc/QVjbydDOnHh8uDvCTs
S35EPTRLueDzAdciruqaDHvYsRidWOHHZKBu9ofzacGPju5jX+9QWvKsaiAGaFOe
CaAgpjrVgS6KP/6WjfVy9ybLCl51877fERM3B2QA+Rvkv6V6+BbW5h0ZzDER2RPf
2IRwj/RSTr/15EqGvH8WkbG2dfRJcUD+cZr/L524oT3OdzbtSb5BzzSSHTnZaNRi
XYxYK3Ot2Udz3hLTla16vwpGgrA/ESXkuMW8EcFbecONZ124eXp3eTR2DLaI99Jp
pV6nFrY5RQQ0t7tFlp8Kl5VKqPiZ3ROnEM6tUcDUVCo6wXgnQk23DEaiVSizYAsR
iZNq4IBk8gzOnM/DiI3lMgoOnPMSHKCNxouV6D+YbCLYeom0NcE5/jmkeMP7z1M4
p1f3UuIv05uA1R47v9fritq7x/VCeyK6cw04r+m/mWoo+5vG0L7ROvsLJ4ZuyNnH
VgtHqfI5Zv0kSVy0oWmN54G4htlGGidsqcZ14fAeDw5hw3tebw+3WiK7960+B/q1
eW74xP69hPuh4/s6nOmIbkhrqz25L7zuJJluhDlFsTrJSQIQ/34CCjcq9aZoh6nR
ko+SiSBKJoWgZrFxJK/kFl0503rg6JG+bnaNNtANTgZmOkhbwvdV9QmUx87raUxi
VTDX7LNRknq3KNu/dPiJUruDJVNqB2p4UckrR9l+1WVpDHDw4FBRwaEq/HIge0Xs
6icfHgl2yNBI4qGkk9VUOAuvQrWtVW/MHFkQjFgz9GN8DRSAIkNCI9/BbUlftolm
FbeaxMI/OsjP6oN1bcGdI1Wjc6CVgpcRKEM2RHcAEbNcubwQ7KHFIsp5u6kFEwqw
JCwPyQcUw79zPVbfsReMmcU9w8Ch6Fd2NpixTXaKexlF1UKQz/y64H8L5WsO7sia
IMaj8EpBlZlS/TjUsEocGCLC/SSlx/VdkG5tsUYlDPP87lp/qLFPCcWwosHhJGqL
PeMVUtFFeqSvmD0E3uE+T5VgP6ffrNIBs1UoYPujiQ3x3U21E0G0DMGASGzMfGdc
x92GopwS5gc/bHMwrxsPMWi0ZSLncmd3G+tIrVMm89tEjPjSZLd1QODge+kY82kG
0KK1xXEs47IkhAMnj9rTYp80rDHENb1b/+zr2jO3UokPjG1rAwFVoMbOiGiRbql3
inKqIvcMJ0mZd8mJwyBwB7Bc03kr2Kn4dk4Kyk3KPC17lsydi90gVaAo48PAJEIr
JLht8ACqpppUvt9AjO2rFH6UeVjYCWQFTYMZ1Mb2qC04Lv8pKXExhOsE0vMVY/l4
WhCWk0YvLkpseAShlEizMNvOTySeWmXl8PcNRUAyTVkob33t90f+2Yt1Ig9CKfEG
rEe0USc+saDvq6vvlXfZsNK1Gz5ZAbKePTMJoX/WyOBdY0kegEX+SCZGJAY5A9Fa
jsGD42ZFzVRZMr9QUCPlvEOdbonPfsgtUv/5f+RXcso2BVzvUjtRkWNSW262wCf8
zm3tZI43Be/Er8iUQPfmL3Y4oEcdU8hKkGp5WLl8ZFvpV8weufSVj+34Z4KMSm4B
glce9/SfkH6Pk8CqNk+wk4Fe/I66f9ghh4YZbNTrgOdmt904CWPYhbk7UO2dymwj
j64I06ou4HnbtwQ91C03Tt/A79wd5QzctNLQwCFa5em6f5qAbV2lEUMOPMvrhYDk
mQQ341qpD+dyD4nPk6hBEpXvGCFzhBAX01+tFELULYZ51zfOTthYwMgQFmfIlmkz
Z1+/wWZzCYAtm7pD8oYlaPm4JYUm1FDDs0r4qp5Fub+vYPel95HLLUAs8m8QgIPh
E6fTaQwp3xS7Nsjsa4gtifymCGTEeOp2Us9fwBWvuhLaeqaV/c+RNSpNyZuk9Bz6
dztnTRPWtHWhH3ZnqNkehwOVGzBPbjBXL7gjaucSyhXVIj/fpQSdU2ArntcAh+3N
d/PFfHVc/GTWBGSW9OAK3Q731T2r0mPJD0oM8KVW7GJTWFruwSHchGgtOKMhoy+O
vvwAe+APFwL0EHnuYpBWTct4FeZqTAnRlfs5sDml7t16leTvZLbrwhNXPywGsqQi
aCAieP9UczPOUhh3MVU7cDZgLfQamhCPrtuoSshDD40+W4l2C+vB1JjSkZl75tP4
Ha6nubkorZr1QQKhcRVRaQwynpAUTlMT4B3ic16UpJ0/+rJFBAWQiYCtnKCu2LiH
K57cWdZ+V3gJkWFT33q5uSZ8oFHE8JiihcKn9rVkKWTqDpye8HLmmSSI2D/BpM0D
pmBW/RoW75xIqzk3TPdejtjcD/eNSkhcTyr6X8EsRYkc70eB8urkIWoTQMAe8KDa
F6TDiCeD7QUnE9sceJxWH21prmSExMRfo16iRFhK5+GtVC4jDlIc9fJALnmDUvx4
VzdiXGB/U+/n7FelvuKUwLgGT8x5i1vsEloO+WkI3eBbchCibNJ0+92OUtcm/eHd
fIEq65QxmwPG8GrrqKv8F0VeXh829/aNcAul8HNuZawnC7ghBk95Su2bG89L9qfn
A3wy/S8Xk/ctoCX4HpRoJQ3gIxGwqgcrkUDhZKyfOT7JGtlSiwu+iWi2b4A8ds1e
b6Y28RZgorg4KGUao1IwRchJeA7cVBZ4H4s3Hy/7VX0xKxVIdYmhJIvCeMHwZVCq
W2T2sqAGL2l5qIuUdzSByQxtQ2t+0xLmQdGeJ+h57u6RdqREosCCjinMLda4AcNy
X6M9DepfSfiYMXWLLi7q/hw4C4oE+iMJU4C+f43zaukCH/mCXZDOW0PHFKCZ5/Ca
T6zJ7lvTmlQW4RFMeO8OoPja925BkqCSzugW4jWGZSnM6h1UDSjJaurHP/LR47dX
L4QCjZqrbsnlQj7Y/v/4LNHS9rDdeN+axNzsE4DtB6tEnJd0g5Hk9PmFs8KO77bO
9w3EcuwzDtkvZTkZGbWYWRnPH4eNEyw4sdq1xhm0DAqjbGa9NiL6LtF6fIPOrwNo
jlSOvJJVWU7p59DIfVFLt3hhcp1yWe8dy5TYgQokzdqIy7z9+phKagupBW8V75Cu
90gnPc/CKCJJjtI9VM6NfUaiUZepqBU6Lt6M0VHCdxoh/0nf+rHoK59/Tvxx4MEA
ZGFoEV1LhtGVLp0jsh0v3fwtq44bj7PNsW0d7ZEzUc9g0D1WszWizAg/sd/1kAHg
jT6gQ1sNxa9f4iMhOOXboP2jYipHGnq0+G8ypHyHhQnIgzW0GJ8+5vEOFfWSp+jX
mvejQPgsAYYWUrfT5rhjiBfv+oVNepY4YTtCMDWQy5cw8r9suNCCS8YnDp57KBqW
SyE+rHjGjtobQ2QFWzjpOtmQQLkxNrYkdmS0blhMJIbM7J+QF5gPvuZZUuZQeMTU
YVKVKbZJjGqn34+DDB3zrbdA/UcKVxpMfeaZ1DAoIRWP2O70VwcRzvLFMjz6cxc3
BpzCxwRMH5ejwuGLG3jEIZSdM+4KBKzEWFdJ6vWlkEtf0y8uRyl0WSgAtNhr5C+b
PedgNz7hQpMYzYWfThbpJXPQS2Fre1jBpO8SfWbXflDtC6PB8BQeY4B75F5uup2H
tl/Tr92fpjpvzmW+EdwNUX0N08ZyO/AVx5bVg7b0a8aofy6CltyRohajHrqhoaWn
jnTtYM384+A2knu9aZA3ZfApZECjok+l6/eGdq/GFNmPuSUBji3ytlBA8UWy8DpX
fra1VGmBWlgzXi2lo0wyLsRjjnDOjWn+V/KNFNN9uFBXouKSGLH6k9/6yi2g+WLQ
5lsHrMsi3aUgA3CVWNSki86V9QvfrglREfgkJvUMGycvI2TuvGE7fHTcl7RVg7Fv
3zgxWA18MSCxXmNdkWrdO4hGkTDGEmj05jGX0Ut4A5Kq0PHHphF9ls8HLRAmzxFn
28JGVJJj6k6tIzkkcbAU/UuvFF8lJkMohoJxtqeSkN3rfeSaEQylCPQ2yO8+eMDh
cMJJG3NaNNH5kfWXH1L5gjSVQxsBMB2xdXUrwrAKOYWeKUI+GYio78LVWDxsM0rO
edBqIe3uiYre3IhjcANcYilnlI9CHyX6Zr8XiGFzqSn96dmd//DUf9yEq9lH1id3
VmehYExAdi48OPowxr3plctYc5TREKy/bkAoc2rvVdEbeRaSqLOwBZqUrrl7UE2Z
/0ry+fEwgwQ9oeFk608K2lPsCBBm4qt8twOcqeqdB5KAmBTF9fSm6xpHKwc6UWQV
8P0cCH6i+ioxKMFTLjCjA6lxKc8MyEoUsBI6sYVj3Jl2EmbKQJ4Z6ASNavBfAzNA
pQAQQGwfAwHWqnTCOJ50xZBRBvGYerZq+UDuJMMKqNue/YfSosruPNoIGFoFkwGp
lLZ8HYIth5GCWUm5fPDzWTouvzoMK+m050xbwo6jNGaPzeN6KfS3C4i91OIU1ZuR
opcPx7hHR7BsJKASfwM+2/yjWYSnhMBqAyWb+UPSHSigvAGRZOUpZCAd/o2hetv4
MZWJ85wA/pkQmFYIqLvhT7Lcb3jm38X831vRL8BxL6sw4jMozQ/MCWHmokGnfPaZ
Li9WJ9NfrTDt4cydFmzzOGiWE9e/cmpAJP/toBjmjQ0LtjQRi83bxIYqknLzr2K9
Xbku/ViLLkrBGHCCqSigmhBCg4o41AtIv1WnaZBnRgnDE3CTva9uYvrSKBc5l5YR
0Ll+6QKZt0LUH+bLYyQ6FH4LFM3WBCAn4Gs+me+K4ir1Czbu+CiWJva3+JBvjXIV
DMrQcluyh4sxQh2vms4kWQHk0UBkZ4079D9Gtq3N1OZqoQ/X3ZzKBx9utjry4SYU
/JhfDSoFgmmpz+9GmxUbM4DDxZGXbcZpeH6KVHszxCCUwO81AYSkoP1Zmj1Cnrve
i2/3pr2oyYonSynoyfGOcOP4leXbdDHjWJYqlkTG38RrnSMixRR74DpRqyCYl9Mk
vUndIltF5QM40W5lGTV+sZP1oOL4IG1FNf1OpO6sq2nZaWHGIaeeiUrZE+D7PIvs
8wjj2L3wnvhivZn+A+maGx3HJsvq85yihmVi92HudnTicDJRaHn44lwfESOd9/lF
1L52BCFYuH+iQcOYWDOssSnTV5QJNFOziIuYfoC/w6nnhGZiNUJgwZzHCn/L0WY1
DRDG/NFyvxtkqeJ4eV4Q81QjPB+5MA4aE2ijbKue5UW0u+Bs/OE6RicvFaILa0qr
faiEJ+G2ZvTCJLy4fTgdSAdVVebhNHPTkvFfTm1fxnQC5SveRq4zypX5eVMkjtGy
DL1lSnboJrKk9+nA5urDsqFmomHCWCgJ+2INkAXzYLqVqU3Hc6ZUm0Isd+8nCK8b
bc/2zbEUFqZXdnXEp7jHn13O8M/D3sLoQZpgPTGnN3A5+0tv4ZxtMpOxNnRfwx3N
XGI6sZzcr/jxPiCViiQvaEwWCGtcqspTHfWJYlksTYWEoHPlfMLynxs2iU0NZcBR
KmRUFeCnuww3zvpWPoCnoH/hhlDeHliEWREuKv0FvAwP64ojpq+w2X/yhe4hJs/j
48OsXXRI9+3dpuPfItuZYeKroWZ7O6couxZU3e2kLFesQL1RxxVdWrpic2w0onGi
79JgioQV4E4Mi3GoFDv1BQn0gWHTedqLqKxm1ftgW5NcgVXE29v+CVP4cCIy/NgX
XWHyBSCQ8KUZYTVhAyDFRdq7zvRgkVFUNeOHfgXk+XqP29wyn1sA71J6aRpNFbP4
nxzBeDA8RDFnKGgj/MAlwM1Wcl34RtqxBiaophA55QnwPpuwU0SDvQ05VgUzot/B
WdGMoyKxDlqbRmU0PZQkLOSXZEricS3juFtjm5bs++t7aV33kCara/Q+I4FNba2R
wQBAJk3iWKw+ve30Oe6rsnUoAINQ6l6ZSkL+Wo575dAi/ODSo8B+ZYEzCOLc14Oy
BXlX+i4yCGfsD0frZ6yXlKCLt+n7/9LwnxFFlWdxnAA7jfFPdzMeRClstdIIuXlV
+NofpqSjdwD4vOmT/DfPZP4akp09svI2EAjsSwZDmZeWzk+EkZg267BQhafUe0Md
sMEVbzrl12gzRv8zfQpY9KT4PWWTw3BlFIM76LQ4fcPvomQFZwLNAg73bv+ZTAzv
q9N2DInALBb2QF1EP7iGwOOx7kbKPp9txuIGQfcd7FRVeqNpAJGcBRzFtcUGi3Dl
u1Q+13GE2U8jEqOuFHhn1Knd3qZFmlLepKJRIoMe3DUgo3VAJqsGYov3zMd5F+Sr
lV6z4f8sRdNO0cmrVxtAXPOEpb2Acejix3gIGQwFAun3hf4juEvnX6vb/abzS+Vr
5s8DYO+KykQyJ5LdgK/XKiOT4aJ4nREY5kYuI3eNccSwgBtmUOVMWkYpWzlotjuj
Rz6VxyBgQgHMJziQ5bMPjPfJikMn/QioQedx6QgyzRe6rhOs9/+knE5oc7vv44IC
CTJeiF7/FMeqA1rMoenYMM0zMbZ8ApjPpgRnWeg+ZkeXDEc6u0Ofq5DekUMzf0he
gmHk3EpISrzBTmTuLhDMK/2gtNHL54t0lRiKr/YkHvYPttsY3GbL0V1Y5OHurnaX
9QgcOcW4Hj+9gXl39Tpi0ckh//wpOd0xxLz+EHwbtEXQfnwslYxXDprJo18Z7O53
RV/iJNzSXqhvCz6nhUDqEkWuGCOXu1y4c9M1xJYtnZBpvG99zYpFUdjVjoWKIciq
ZBlG98VgFhDUiO/m3dWQ8gVYXt/R99afbSv5qyVLO2mqWQw26ho6YbnPuOHYdcq3
RFiIzmy/oZlD9QxGcr20IOKimkylE+eFgCn7r2urdIolAR8lrhe1ArlIlAeer4BN
TtiXWFR+fKbI7qwz+U2k08y+8xACQid46SnTwrZ5mw/tXBzOM/zMBIl8SVqZ4/yh
2oTwEKAG9tLldhj0jID0PlVZdQ4EjcKkXrBXCsnLJliBBUoreIyad+Ng/KddpPOd
saGsVQv50uJILFXgaoXQbBngQec7Zu4FO51YkXV/u/zq8Vwn2RBwPkNqVfWJWXQA
Tc+fH5twiISvRkYLQoX0mSuhdkwqWaMzYNZC0VryU2SOeKLBrBZYXaYtojhqXzNw
OLkR9YkUbeXHhZCzJZyaas7KsYhnk79rk08t84lzdIhylPaeNdkYI5gvDgU4egfP
6b31wN5b5kaL0ZBIxcmwv7sRA4RxW2E7MKn7YN6+goK1pN7g5GGC8XLGJK0bQ3ZI
/FJw8ZGz8ut03T43GEZrC5vLR72CEB7wdeBiACMOUN8EIpBM5fmAbuPo9Z/E1rYc
VEi2kAzlG3ikiCunWoG2hNRh2/eaMWpi0Il431CzsXu1PGUDCXYaiKX1JHCfikkC
J+Vu8Veqv+3wDbme7pqVROP8AXeTf6SNWmLRqBdWxtt29XnBsZbi0eYzpJ8SbRxm
yME++GdSxtEeHbHZ5t50iZJDWC3zCQha9FcANAKT4U1bPGyk4oJ66p4CG334Di0G
f85U2S/92KNSZyM1TnjiHSxkpwsWiBYD8a6HU81uRQriAz3lZ7eImVArPu8MpPzC
2VxpV1h7T0V80Lsxq9HLCQggTYE0rL8sEmnKlQn4k1AgWkdKlyDvmKT7ZZON9sTJ
UvPmB/E1erMcntsZUaFCCZ5J43O9U4Nmyny4etg8xtVKWNvM0/wR8eTA4jSMIKg1
fVhrQ8DYk+B7Gqir1zR5QtD9+UDLVPmtNlROb1ANwY8UeVMaZugC2RBzNMzRwViJ
qdXCUdyrRBRmOejlb6qqu4pIIn6Jv3E3rUvBfgG5eo9mj96LjzLp9oV0ynRdIGJN
blfBJ94qIwrmM55c1CbDCKDvgp47kuz3wSdlkFUWEAHXl5g2KE1VnMa8jZOAypXV
Jy4Q87IgsvllJVZgeAkwlrw54v278941386pZ43VJ3v1DQvNZnveTs7Ix59TFru0
gl7PRHKmQSiNCVN2YDpLeZHqwOrTMtK3deiwqZpe19psnNRhk3DI01OZVzPnVACw
xfjBn0r3/uVHiIprLdQguAFc/a74xQcGx+xsriHRqoRjSIy+SKa4lBVIG0zeln+d
WOs+mZTNJY6VMRi7lsE3eiJakLbBEEcXCUJcSk/p4Xa8NOlQxR59GRAr0ypdg9bh
jCjsYY8Vm6kVXBbnmqCK+yI5lLZ/McbciLJXt3SknVZKTK8bt1bMlG8FyPENpOeN
++aOKlvf8kW9wrfJrG8B1SH+kdQ6b7+03off0q7VZ3jlNKnkAanUYv183ms7U/Kq
0+EnosnTBUgEWzjIWattt/peUpyjQx/yMIk51kAeHAYNx1EXa0Q5bujCz4v+Rg9c
AFXw863kGBPY+E3p2hpra2znkpdfttAXhEG/Y/00wVYlWPXQ16jk5iLLghK/Uuqn
j8VPEWHzefFNH6TZg44753CBJkX3rfIv6LZJOLCOuBw4jQoBxF7oS0YZ179KJPbJ
tHHeMqU4HFhy+ikWhr8hX/X3AcJtb8UbjMy7/pd1m7XiON8DvajTJK/35XOewxsX
Xz1PDr4WhSEOUxcEHa9m8c2r18vAFlru8jMQxLRCJZ+4CfJj4R1mi3uqNoj6Dybc
HV8eBajdIqSgu+UWvHrDiN9McSQZ8lVRj+rw4hRnSy6NpgvtI5SF5KRpTk7fJA0q
miCyz+ibUq/O6NkWXvjKPPl4YQNujlQp6v4LI+co1aIvkWipPE0txRhJWZM4/Cnw
GAL4bD4dTy6C4wpFzpSkM6V7F+PJ24BJCHyE4+z5H9ohXQpAuQjcVElTVsupjBRF
x/55HaenjJ4Uh1QA504vU88U+TGQQwuJoLPO0EcvtAJrRlrUjYwTr3/QArHKIJLd
RH3C97Pr2sbTxooS23UOfnoz51z6oce4bO+sj9hGUxmlGvCHxEeApl3YVgjkQh3A
vmHtfGDo2xfGkO3NRXJs3Vz614Krm1UutpkhyztqvcUPkocMo6I3i8eCmrkv/clz
rnHkAVF24R75Rlh+5yKVpAiAOAadyP71r7eCvvYF1IZ9Js7Fh9g8Tb4Q7SScj4VD
pskcjUTtBwVgx+zo6Ydnn6CbiLifiKIZ/aVo4TiTlg7S4mQ1Vr+rNkiIqpBf96g/
rJokcqRjtkkKNlx00nGATuZU7D0Y4SlueMqYi7zIQuOzuwsWbDG/JJclQsd45ZlR
nZQNaOMJPgr01V98Mep8rX5kkycwwCtjSXWKmSxoThTwo9d3wR3o1Sa46wBOJfx5
ukUq3I0mxstPdREyqaN9iENvYTQbONUmaD+tUODaICaGUfXSi6A5kvyfAVGI2GCT
LpgfiOJHi4RHczwRhFBU/R2AYNuA7gDuRK6ZcCcjYLQlNyW28d+fc5Wl7/Y0cfqV
7o0jk8jafitctk57lu72lGEqhTZLsRHnOaXqn7W44Uanjr9dOg1bUOYaNAnYGM2E
bQA9A4Slq/1KrKCzjarcJMGlEllUpQw47ihTVM+SaUerFX1o5kuaApJBvp1AwV/j
vV3YKF8cwN3RL9RSo96IOBkHhwuqqtsV642GFlisvdefTG0EOvCYA3lXZs9lzYfw
83q91auJEdTd6XOkHzn82FSwGJundYsiDpfDDPl/JsPWgClQ9Pu40zXwnSSoWYaY
mhgLKpS0m8Az2HhNlk4fHtW7w+/kHkqOxj7NbnjYZN9U4sB8B6MTefFrJsSoUNtM
yqJp3RsxQaqab90+lfgbiN+76xMbdrJ+uJYFicq4lK65dyFu1ZE/ph3KSfTtlhik
+0kXOdXk6kvzCW+doQCj1QvmDie8T0NM4pCVuS6S//P2z1nrcEOYCSe0EPIijI8t
fZKQVOknFqmQYPscjHW7sNfJvQzEHd11VKYKXN6JZFwOx0K2O2vz5j+eC7nwPsUv
OvIQVgBxxW/EOsYq6Ba2U9xbp/c75vkyOdO9Y0yOkLgwiGE6Pi2nSi6Ue60nMWFW
p+C00Uid90VQBsn6qv4ztk68VsU5X9Lq8gc5nWbJgE2d4YFh0OdViQ1NiZ76mQEC
K3A41sSfWP5l91tpHTB51SgQQM295ecv/dbrbdKR0LQJOgqIEEVig0VpOZkSovqP
daqnNvuO11N5J1MQr28MZ6EYt6IpV8pXVSbFKL9JhbuWnHMUQB9rUiQdwgb19ln8
haPCvSMTGhmGsy6K3jyxV5QU2OCIJe0ZEDpjJHXGqTb4RO1zJ1mmRCOzmmLcM40H
0ojfv9OPd2Bu3X6IRHGyRWkMix0QTJ407PHEohGBS+g2vko6Nm9Yk08ysM0ld06t
SrcV2TmmJmuP5NHQjF0kh69y7Q8drym69zHAwxc6946rQ6W4f6/Wt8kUBoqzS+3c
22zL2tMehzCJVDeHM4GVxzDkuUn8RDTODskqjTOLpiUO5IlNEjMTktkdhTZfChth
57jKDgwx0C6xbSKC5KOX47xu5KLl2Xb5OXGg3+CjuoMMU/j9YPHjnSlqh9ltPV1X
xX2lnxDgt89d2gviK0bUUeCZcyS2YhjRqKkEwkvG03w44HVZcWaKiKUcu8drUJyq
Q59OGKjMZdMnszU8uHDY4Ufjjt7VUqZLkzsD3G9toE5n31MuCKRe1JWdUy0VVsDG
qmDwiUG0nx387q0msQLNkbJkQiSSMNu1qCJWa4S9uXUuRsGqze69M45U266d7SO2
5sv75JTDCt0QOS9n5xQepVR7zJp2BmJ6LEPyU6QY+mVew75Zylod+jJpMyv3dsM5
9bGAaKYkEDzDwHZ0Z0wXNb4fq6Qq6uMxZzIm1GSxtK8c8eCsVo6O2pQMQI0W8tAw
1trfCnid4C5NLwyeuJSs0a97JwV+AbyyvsFMdPRolXidTd+J+XkpL2vNlUQkMK8c
/Rn3iJz7XaxVm3qMf4Yj0OSybZU2teTkbgDayOlliG5B+t0ebXmuu02lSQUUz+l5
VQil/bpC3ekVmvSGSql57Kk2C87XSle0CbsE0fNHKgpkChpE/Y5S8MrrRBAkkgbK
sur2T7aFiTHHKYGtHuA3ZW7wBdGQXtEYyXKz8Dp+0XsMk8WjGuz/P4KiA//x2b5d
8PB8AR0SbcqBQa9aBJDhimT4T35PvY7RfmHY100TKazSL6sinF0njw+MvOnY2r7q
+G7EjQwXsuJi0BOEgk7CQZS6T5ydV2fCqnSjnGxq9K9GyMpmfeWTCUIaiSpheFoH
CBlsjUcl6MEq7RnP2zi+sB7GeOj99YftGB4muFDFqfQKs1kLrOjwEWOU1PhZWeEi
FanG7hv3jMi9Mo5fA7jeAB7o+tZ6BAM2b2yGaWgGT1XtJx9qKmd5IVD/jM6Ty96h
X1jA2Kdz+v6OMiuqnio7pIhvHbMmpwycUSGVnU13nFjHC84FiJJfIWNwXbPWyHLc
KKqlM1gGWxe6hyCgKZNpNJq1I7sYTZIYxFrPu+xG/Y+G8txg1r+3rhqKMc1xnWAp
Aq3rlyITM+5VNNmbXIdI+ZHs8/sTp73bo1b1Q86+VSbrSbbTsEpMQmXhd4OXQNSO
f+Md+Uhl0l0O6vEEn2OE5Cb6qeY/SXZo9pHZgWS8ZMwUtBBIQoM2ERa91AOYjt0G
kQLdEw0XaD2+wsvCgw5Mv68KdT0F0zfhCysDNeMND/uqpT9O5DZuXWRylZuCo4Bc
GRIWpY8Aiyoo7ynL/reHPnDUkGmIqb//HZFOJdO0DhRpI/IutAxSDpSWkJtf49oy
3BMpikf3jTHghk3QsnpV8nMsFt543rlrl3XUY2avFX7MDorEZ2jswEzJaWKKEGGp
ezzPVY/TmTxo7/3lOBTpPDtluESCxPzRgIQdXYvvIYFGEApfKL+LRPSEluMGFc2J
zaViWqxuRfRjsoyvtkWXNVnKEpCkFwx1kFVWW5S5x4uhj7P3daaiG6WHHRY3IPRY
q1qs1zNKyMVUVK429dj2d7iiPuqM0xujf6eOp9tBagzLiCwVEaBIcXijNwWPz1Xv
uHVFkC49lIqc8MlqFg4Lm6JVr/XM6qwzuweOUP7c7ffeub6xnFlQAHzdtRSCFXye
DsBFCB4TLhskcTxqcVOL+iDICfXQQseE4zWQrYyFwxjEDBAgw/N4MGtQss8MDURt
eH8r/tbs03Gvb0liZjgzcG0jWzd/9miHCUK/rLuixhh8Y7/JdFa42hrDhybPo90C
pv1EI4755CUUrMdVU/u0I/y+JAwjGKVZP9kQLI3cp2XzELyeKnpNkkkjw5WEfYLE
QhKpBTEEtC5UV1yx69OAqV80DYRL2b+tgSzPBf3ck/7vrUedhyJ8AT0lPYD8DLft
EoKzICwaTmcXWwcrjGqEhNV3l7J145FiEP9hND/BF5hrIgcNIV2EL0yE1mK3xuC3
EZWbPVKbxK/hnd/zWaeJfxXKzwiJ/DWa/QZyJOowIJHWcAqUtHBpNWEmMj/RpIec
uEcABtzcDvF/jYiulVOvKDcB5C/jScy8x3K9W1Ev8NUQfDpT7fd5Pj6JR8nDnalw
quqxW6k+84K52NkmW0pImsLgVj327LVL0/svyhmgVP+AIb7G9OK7+16NhzFHaa7h
0RLxo3k3LD6Es2FBYPOMQ3i09U9ppfT51zLOlmxuT1irEnryVAtjcNJwKJe4+ydb
/6JHnb5epNJmO4LTxmWMnHnV0KmVkvhjhxABKp9tz+U/2VLqNAw2Y+xtCbi50Hxw
V1e11BajEeszhAcvxId7k+6f2qcuBz6qlpiWD2xzVA2IuGf3kQRFt/PLAHxJQ2/q
XpVc7ZSDEAksOaZPF0TnxOvvlipBZ266714ZIwW/nyIdHjqMH45lICSwOVbfX6cV
SS4bkUOqGy4UqoJEcMXqckly488iDzd/mLUpPRJ7dRYSuMPhafnyyeprEBKgGwU4
amDLs2jzGVJPEtOq0EouJCOHcZfNrO7SrYYM3UohiEVDjdxaUbqt77PrPKZm8BgI
XIUVPo+jPf2fpwMoqeMhv9EF41z7TUwtMGhN3D7qxIgfFufAt74Iq31ckdJTTsRK
oX0tVxQVEBKcmFia5bFJyBcQ/T1Ps83/lyOLAiEr5YWgfOgs+88+TBGm2sholjYl
8ito8QZsaefWbbnbKxVMQ5wPypcwqZy60RUJBT7yTcFMScV3zG+wTkNxe5m/89t7
rhAG5M8Uh9WHr9qA0INOoA1QgAE/IErEAH11OYXYvNRTx9NOWygQ6Guy7p6mzLZx
UGI6Zxy9OWHnN15ETcA1acq3R4acOQ5S3/C5dReW8/rDQLW7xThxYPCs9fzvHp8M
U07Y8g0BbfstorfWqJLiErikGfxpBtOJy+T9/ncspF+/BonuiWQmThxyQnfBkPLD
rlEc6CcClr33tAaJgxsEWT4NNVzsXCJa66UjaSYQwfUgfeA1kudhrvmS/N8OonR2
lg8ZGogJFIiyBZ8uhjpbmjXdOy24P8d4d5FNXK2uT+ZVrR7+PiKl9B/T2MLcfAj6
F/F9Jtkkve/1yz6eWepikD5WLl3bPYHn9pP7z5zml2udmEBvtuJJ1qQIp4KEtus1
y2R4xrr14gvOJMkq9k5r9MvSkPeXGMpid5HzoWZ+aQEKQV2NwMLM5+c3hQASuLe/
9A/FJVwSfdx03opc5UcZcoPHrr3fiwHaPvU+r/pTMZ10NjlgfJmUO9wxX+z6huln
dI+zQ4oKfiG1YsQ6BnPxJBYPU8Gcjo6ME5IJOzzN/aj3UPy47XjzRcevMdy9Hows
Mgr2BYfUkkXgyfn9rdEyvzr9z+0T/oQDhROHm8R9XkjI3yP4J5ynyORf4qlepIWH
uRWt4Emzs26pDh1+OPw0qpF/O2lVd/Ii3zmiiNFpCm5zhMF+wzt/J47zfVuHKLnq
16qgzOzfojRbVduc+2F5Xmt1IBca/YVByRnmEdg/zSye1+Kjpzxlc0nDIxyUc3Pm
/kPyZik+Kv6kdK0bsY+idVvn2/nQnnROKFTp/3AljX6dKhW+vbXbQBGlhe16rMxM
oKk4ym+uLQyLsDtvK0dp03cD+d2pnisGxjy2W2iXK0HayngIB9XL9w8NbWrn3Eg4
IpMqs1kNiQr9dnckCEcAwgLAZjuqvKB57OV/SXiu7OIZyuSgY4uvc0BjSei6DVeI
AmAywa9GcD9WmwJJvn1vJP3zGd7ZfPUsqomVVlWBgN9sgcrrsuFLZk6J/wVLDkZc
gtl/wKkAfi1Or6PZTAnONFxE+RMtOMoaVHln9ntcUnU/Dm1OvSxl47UbUQGqHTaJ
yxXG4x8rdc+D2UxBJDcpDRBdGI8fgSsXxe+IPRhILIspSKzwo2vNYPuyPDuy3lyE
/7e4eKdnF3Vnq04hRvq9K7LnwmDfk+U8DA71GfiFuJnyn4PkjDlZzxtaoMmuJ+Ci
xvnEf0bJFdxlZ3KuztFlVS7kHsHGHHGrMO19lXOraR2rbvRwn4V2VERVWmmvFrmF
a5Wf5joia5SNRS+L7VyZvbrFsdkGr60GdY0yWUu5r/evAEPWjzUCxA7eXg+SSjWU
aGUyyFlyrxOBAUwuJqcjuYgjrOMB5QQTXuNlF6AujSYeSxSO8aiVkQ4LRmEtVmfQ
8i+b9jqXKYKjkt6KxQU7ERGhkAqBKK7Y6Rdjd/vMo+D4PgNaLWd4lgDeL4edJKYZ
BlP2yGU4nptptjRuGWsbcTbbocN7rFEcJoFD0RpvahUdoEBV9Bl1iId4H8UWM3SQ
9mBWZCHMmaJ/n0p+tHACQ5kGxAm4cIIHK7rSToOjmvxFeIj7nL5/0b336Zmd3e1E
cmUQbrmf9elhBal1ivALMmr/mjfOtQT06AgPBkHff5TqfLWIoNaU0BuNb2CBSuGD
ZzcH8loafPhdyb0T6dmteyw3uL7+N6tDdHQBOSc6MJCL2I3JTsHSVYq7T9+88qSx
pDVgNG3zppMcYM1V2I4E4Sz8EWWh42L0PlVMJGwe5sP/7bp30gcM7Dt2UESg2qM+
yW+MtFifChy/xSFO4VGeh8/3w3ioM8IHfV4XIviU5KvbXV1mi8Fu2EMbZq4wVGHn
sQbkyvDyH3DT3yAGVRaQOoAyhPtOH8BrCH++mPwvBjxLrc31XAMsXhydhAglVwAU
X1NgNt9lkM8/5sjHVOETH9cYqzvN3pFNyEZj7phAaxZnsTDqIxZgBvX1GBdxP5eV
2C4Dyw2zVhxinrEyFj7htkHMBiH0gPOwzkjllWl1DnoFvs8X7mkyKwmCH1iGS7hd
7kgD9DMvopqYxn2tger204IKpuoxQMAic07+PWFI30+fYyS1VX0JpxTrJZ82ls+D
12SBDcyWs1z6iOOx8UFXTdTycA0Hz+pQK435G0PMyMrZb8DoSgh8g1vFd49Zf87v
YVg3VlgAhPC45DVsKuP8qm0T1E6HCSldLOxWUk/kRERtGrfmd6ugjtMWMq3LfMEl
Xg8pF7yV68SHvb7tQmUwdQQbHdTubhp95Q+url1R5gFVQsvdQeFQ5vz2qcpZBmi2
WC93lAH8FdAxOXHzNtIZuGPm/gM8r8DCE61VKzphG9lTfopa0GjM+7q7fCOVPQig
N6xs8b3NozrpVNFr8iE90VAWVI9b7UB8jSBFSF3PsE5EPvbpJSmvMTCQ4ghfp2YK
pJeMveEtD8JB/Q8SStrdfzgTPvGl76+avkxkA2AmatMh6+cSKmEFUVjAKS1qU7ny
Bww2uf/SjUw7vyVabmVBaVkum1lreC3TW8B5v1AEiHr53FsfnbHUNgB1oy+PI1G/
jpKbr7k3Tyz8gER+Mrp0ckp20ISoAsCczVRYVFPUG5mXVLMuLh+db28uHqLKS/7B
h5p9rBRVUB3vg4lTAa+004AtnUTg9YC2XTwcAetaWFApbUasxwn8N/1UUQOZHjNB
AMaqFTlzI1GRF/CkWdDYTlPMdo4gxdt4SuTWkgCYOpSUGLyX45oKQDKXkq7+1VDz
j3p/rYz5IMCpbh6fc6zBc1T+2GFBx9adtz0jLXLsGp/qXsR88EksGQOndAJssXET
Add1Pz3io8/UBHpNbdmTe/mDPMykNyoiSUP/YZZLg41uOUUs4h32ETj2jbAAalfR
an9giawdN6sSew69NncHfJaFIzpyGNh2WiU/kWdCmwRqysQHLJOKyRoeMJ3lP0TZ
POEx3f16fnu+rnOXwve4ivUatUjPOft1gxpXA6Jlm0NP14QnIkhPYeRiqrAOD85o
079/aeVq7btc/Xc+JwwR3raKxTJsT/4hy4ubvY7zUkbnANDmtlC31Fz3hwFdBe/c
yTNgJ7pVB4M0OI7/C74RV+MV1y/buO38mwYr+sEKLpCzs9ul/heGNhOskyE6IZPB
exu3MXSjdCxnamasngzmR2ARTXGvuSuPPxw5Fiy0SncCD3PuF1xo+9q+e+6JsxIH
ypo42N/dpeSuUbzM34JZ+mTKf1Jbij8NEbDDqjzwayIKEpEfDaFK1sC7MxQCazkS
KJOf6+aDSvxWCQQMpk+T7uB4j5gmYq6OsLTVFSklzHPpX72UXsK82r7VLcz1Lqx2
Po4RPlEOI1xNd/lzlLZ0vUnSrrxAc0IDK5LkYUcEnY/uXjalfERd7yaHdGTVxoxr
MPhL61SuXSL8W1OQ0Zmc2/6kSg54mM+bNzKzkdfmm3g0VWXLSoI87iucyggsT5pS
9NAdCS3unz5nRlOzlhJbAShWEDeplxu6wZOMzvwoIN7XIUV7bbNLUW2t4Xe5x7jR
hziWPQzb2+l6bgKm89wuzsy2IxBD8SViJaB9NTCX6N4bvd2zh5z/Kcz2njqUrLNS
OSFKbCKFl3ptKidYrEA4Tknn8WprIL4qwifpYNzAcdiVhYaAKYPj9FMzXi1CVEII
1K2WlZTY0chgAO+BWqn7UYaD4/dsgyEZgXpw/rVHzabc7LIPHfCGTvf/BNAdIMBn
2iLXyP+GQ5nOEBYaDT/3TPPQhuArx9/tfWOvYHvXFZD2lasS3nr3zbYt9fvzNW1V
SeO+RAbiZVLHm1M6gOU2shc/IE7sWsDx8RkCNwcrHbwj926bZRIq8w/0GaoRIzeh
RtRSdPrhDAeKbRZF5h6UT+83hb5gYruzqAEQuUQDsFBm6LbOK7ObMyYxSilfkqc/
oPD+wD8pBH1Rc0XOA3cyBsKM437SyufNzimDJAqDx8zXLCgD/r3bICSgRWX64xFn
w0g8E4C/m4t3b+JD4UHTpcyWlBZA7ugWmR0epTcu6YvC6nPnS+qVjzk5yvkug13h
60JsdmKDfhMD+TAFsWNkLIEcW9wRR3K6UDanPA2FeCbzajCpsVBMFSYy0BoCc4Pe
IqZnA+X1xMCjnF91kq6i7xFI26+Yn8XCQbnVTZH8Jxo8dtyF/lpKGB3vD3zfIYry
Qn8/bEGcbdHccF23yC1P4ew0IKurWJrC7K2pdNJMzXNt/K1+LlWAh2Dqdckrcvpx
yO5T3aLegR/0oTFp9RnmkCcmcjaMKY3Bo1dtVZVpzQjV9n1p+QPoOgIP53o7zQtQ
Kk+DrhL0phw4UN1Vi77mO8KtHSG6qB+vnxQdpliriJBjitISdjoIQn9X29osZ16M
fjhiR4jrlWRRbOxiQTersKekQ9QDgCbh0vRNpSc29i7Z6C35sjtgCnLVsm8eUhVb
dLHQLicFv1JKkrddjmxORWB1MiAfHoBtiqMHDgaTEeSfiEnDBQTmNBYkrLwa0Ohs
QsOxnAu5E5JhJ+okI/njKycVRT6/XrsE5qU+dCkrxGocBe2t/llSL5H7wwNXBtEZ
5NA7qJYWBLLIK5MhspFFUb7yAYIKOhGTTKH0/D74vqolAy00aLO7E5tOfQAYbBgb
4KZ+A44mgnh6cgJZdl3+xR9AuKVbpvkPvBkFjirb1421qn/WWXLqxqe4td/diTYv
zOGs/Z8z6XiyuH4Pq1AIWtpUuSmZJ/H6u+lyDImMDDo2wfEEQTUVD7eFFxYoq0sU
bcaBT+Dd+sF1jCp8/zDPaGfXQPCmOtkcni3ay5WH0GPvYdp7uKMrTPI+G6gWw/sg
i++xDzikalFO4Lv8YlzD3K+mauMjRath1mRCzxqaqRnE1IlEH4RIT6Svg4CqnPVx
NR1Yh+CQNSB3MP1XcHk7zlb+ttoHYvLLF8VYD9yZdI7kqIwfiL5K9BkAWUzXuCoI
ZdalSq+ClPQ3GmmcSQb8WPMUe1Aqnh8OkQ1h3qUq5GxWqxGc2NuP979Q4nic2jGV
SHeleScXBJDPs0PLUZN05XXKh2FNlGLuCj0q8ZesPORwznPKiUumHt7SMuVMLbII
GtODFR5mg4nrnPYGvMiVMQwiqRRpEItdNb0fxqrptHmx+z509V5+84oFV3Ou+xg+
9exO44g1lMxV0mj2ayaj7ZBtyXqK1CVArYUmRp6LBejmTUjG5RJkciY9YKxcKopJ
2WgN1AtoHm8U6gKcWQylMOjuMyu3LPz2eCGQ9rhxsFzLh/hgx0+x3FK80tA2M6Od
eo2FeNKcBjA3G6IMNylZgj8fGRhxvHWMW5CHjDfAkcekcYohsfXPQR+vZG+Y4k9y
2xB1S66WYqseKAGX69OevrPtys2WESVYUkS4tWRu6smdJNXdcVWOt65/PtHlZJTs
whmnsG+y8qVt4sfybSSPOiPHjRvzKxMvrKrQuvn6VWyYgs3yjKQaJ8SxzDxuesOS
igkCuZYn9i66Us54NBzlVzrsJ+wo6qO/x9IRYBe1IyU+/1a3yngFm6M4AdYiQUwU
ZKQOnge/MIKy+D4E/jwhjZABlnlCH+e1/jyf0Hf1rbx1URDVeRT7ioA9+KtuBliB
sSMVdQq48kltywpUpb/VJYXHRTlVVF5sjN6KdAwowxHa4EqwbIMYYxYm8X0yMhdv
3gZ1ybHl9JoQxZ2arPtSDxR2/BGPI03UaKw55hkiaFzApXhgCbldNVKap+hdqozb
Soic4BJkKT5J9IQfiLD0RiDZhI37wwuRqC2WU+j95LO4fnu0ajUpb0QQ3+fmMC5t
PnSYJNw90t0IwZb+FXjmgN2hxyHnAM2RBowmsuMJVIMpDIStWKYnI4rgWZDTcTF9
OaEn6RXhlYYtNbxmslPLarZzl0qH6xpAWwuyxq4v2cCiq3+JSjNdcVGYu/RxDgvF
vm8m0ufWjY3aD+I8lCFI4bv/0w//3g3YnrneWkvPGhRMi2bYVCn2gUYlJFOLHRT7
ydxkQaCsO0uXr9DBKX0mwUPwg4Cugh1MyXqUA4rBhgJjTluaPwFgb/Ws5+N5OLlg
vGTUVVawTa60NN01lh//ERd9cKjpihCPp5ZujOxYjqOb1ldDin0vkT7NyPeyC6MM
cv8OvrjWGtmxsP9qcDrmpBXStWEArCAe8sRjrnTO/vcU0QMbkJwGjQIcP3A1OzrK
SXSoHZskgL0aYJuqi3ZgHDodwKbQkxdqPmwJwlpjNBa/KnWszEmA97W0yCskl33n
pDGPgkVRH/KJAYHt87ZF3jEXBTzZy/sdMfGMYFX1Cz7xPv1t3MDxLa/GCV7yg2EX
iRTdTKouJTTC+TnwJmopPE9ccLhx6lkluxCgv2Gj+bnGMvil6OsofTWAdj0+7t5s
JOEIl4HTIHRPP4YotZjVQJ7Ai3UasJNlo14RrIprutgWWQusRFcYedPXQwB4wQJP
SCPJMC4IFauV6ki4oBjnmFZXiPE29Nfhyzh5Ya4wS5rvM7+ycNPtxhhDpV2A3ztE
Ij7+lJ/ss2BIdqNv1OyxwvBYLFBI7LU51dd58iCHEH8c9W3X4w8J3NhtsJadqtc9
fwJzw5ID4+UAqXGJ/xd86MI0Zt6As6LgpmfBFRcfO3+twIRX8MLFNApNKTO9BgJR
gDr6baX1NjcegJrKRinxd/7uOoD1iUL64Q3wSk7SOgbx/38aL8Fkl8QL8VRCGzmq
ZF5VxWhbKERVVrEzLeb0QEm0gZS9ajS12bk6J4Dj03yuoXpx0+JyVoB/HtHMtMRW
oSKd/Hod6pvDCJjxFUcdwD76hsoaqaqwgNDPc97frLy56QzIUt6tF7Qa1loaWxAh
7H9C/TjcS0OD5EpcoyyzeBoEaVSgbm8wMI/8O7+KsVOpDXdMdCWdFLVIePNeOEiN
OKWdjaj/tCPpGh2dkLzwkCkZne+ZpO1yueZsGb5jDkGEZH62DJlAQeeoG4dHZyN6
1qzkv0dwZlnryMyZiUG6ly4Aq5pPvofNkTjiSzjuf6wV1wgpCr5SAYldHIZCEH2B
PwZi7i6Let94aDLIYa+Ul0tNaU+v/oIHqpNc1QUp7DDnBhnXzeuPBTQJSnMHi9sC
MZaDsa7UhifOtj8/H5jqQm89Vt6rRmjeV0cqXc1Dj37IcxxZnuSpY3Pi5bdWi+YZ
HRtjOC9VU0mxXJIZ2Mgl37WnlZivPbjZy6h6tunTwwp/9oycHBkG09bZyfFASwYB
Ta9K1xAPjJRn42kMbjoTN5Nd7GfUXwAiUijl/7sWaCNF27YG382OpvAe1in6hjjc
RRSW0PXaJorKTM4JkznsoQqvezrkMMLamstpw70YrSISafp9/rVW7rPvqfh0QM4g
Av8k9Vczy96dLVU3FMlbZ2JRp7Ho7RwdF1VkyJyj+klL6vLp5fhs8CZzMDDgB+Gd
l2f6CDiEWKiQCL8tSbJH6HJlIUy55059fi3QYTLUnVFsMG27g5AdzCk6oWREuyw5
0wu27Z1E1890G5qBLPH0eZnYne3JeS8gv77mxe0Y7ctoWPSD8gzGi74UivYALw1t
00rRQcCV+8TlbS7WOXb6syjpWgRDofspXXg3erW/ILBnnR0EWeFBF8QNc8bls5yT
ScTGYax1/RZGyhWvi6Bpqw91fqFI13xGifwK1mDnAiOgyBzen92jr88n9sIGYkP/
yLUX7lp0H2tT4WtbknGYQX2GiNxs+de51B2sfQiiEB0i3goqBiCcfPas1F7Z9SMu
3dqahTss71NYm1Uj6e7dc6Ld8P0p3i4drNiGxbuX+FUyszaEMj2cBW6p18vi0kBA
cDJlQECeHUi53V9OFrat9jl8Jrq13J/9f/E0xofO3LzkhO3jn3z8JxAbDCZWDJLr
E6328m1qGDMSG7cD3Cv9KOFLDxhtgwwKcmRsHdw2L5/GBk+aD6YrbrQhsOMLMeOj
u5DNovJ8XGbYq7wqHqxkA2r8He1CeAOWGquLgIgMBAFnPnVLjhaWyCI8iZhz5wLI
/jJsiXoIpzWotwSLYcecPNbx+h8mPFZLexXzyPnR9oCTC9UqDQ3u/0Io4XJhClcC
8rPqaLeGBCSMgS9EIaNmPiy06cH8xsbPWZ2eca9LR1SnMTemAp73M3/bi9SMl3B5
lx+VL+DCAgK9sybrMG3vu4mLmPtRpwelZQe2XB/MUOCwABt48gNktJG0a52JaBtX
Yut9Hkk5v/23RdxY37U0nx9Biuz75R8OW42RqJ6uGIBeOecR5xtgiJTS3pJbzFN7
AP16wzqCLCzcElmtYy3W5aKVH+bs8IyTOI2Zd5aUBT1c17y+DxJke2eY/ma50T3d
jxTaHKIw7iagt4elzdwlJSFBiBv3fe3pZseZLmaIdHJOn/3SpgWxtHw2A8Hf5hH6
Q8BhMOuhKMG5nO/50dyIzeHp6vQw2A2YBIDvimsZnlVkaj0Wzg3QWXelMhQdb7Wu
D3GxTeX9wqGszB6TOKnwNR+Ar9YuWbEEbbi6ZV+UvU7tcdhk0aN4KJ8kKbOr7jP3
a/C7X4Vu56iwr7gKJ1ub5B3xaJCvtsDt7JWUq66kbK84hDywjw4EvNca6gZCsYxK
KOxillIzFmTOWpFXwjrAxg7wx0Am4DhYSi2dozvdKkfFDpX1Q98UxPXH1wa/bqzo
xiATYQSreIVBOVDwy6IR3S9KzP7Xgk2+WoE9RJXlwRnTthAMxby1YKuU15o6tLcQ
j2xHXO88HTToOVT79mtvC7ASPe0hwd8MJnINNPafpKvmupUCtxiRjMpvfYJ6cfaq
5is/nTvc+SiNhdBMVMjgtYq37j+4oox8rjwEvqeJPLVcI0wak480f4wZBSKJT1p8
5gI+SceKcow1aidDdj20SuGjU3PPgqiywlZqApzrhNaiWb+dS9HEdO5Ob3PIFjEQ
kT6aEFuh35SxUlWH0rHvOAFy9zOjqBvv32HHivZcYnCsuSYDQTu9+RWmTchwotUq
ltmfB0F8EzkZTwEF+feWNNgT5ig6anYNDJLrQh2/0HzSXjrWVvkqRDcwR3sISAU1
yK7oi28muXtseUhTJXAeNlmG+NvOrje2Q6O6GtJEu1Awyq+BTPrMrHWU7t3RrlCW
7ijyTy1P6JXWS4SkQcWRPxFKAjAM0iJ+CWqjDi9CYps/S6lIIlVH3uHR36s9WrqL
jWanfNaXy4Q6gUGdoG9nr2/DKMtgi31GzEzXuimfngTmWOh9NX2+sJS2Wxq5DkL2
EzTych0BLAs8lM23AARseEXya7aYt++8yDApjZLCvWN9mHjN3+zqqxc0YBTUDoH1
sYZ3YWX0tnpCJlvQMze+dxoS6CiQLyvN/gw/6XPCfITEpCOKmyOsqVXR0yXpN/b1
wsFG7ML4N2U6dP7KEuU4+oT06ag5uV2dpEF5uIFL3uhRg247U+8kiFEi+UHYeeu0
yv5oD6HUTLVvozVib/4TVrWMYloLVsnIkLBFPqQbUlFmXJdBuR18BNJNcw5/n0Fy
h+cyqLtjBEdK2Zgw1+aO+wiNiDWqiCGb9ll+tL/L3AgzttFA//mbDpW0Z6ETNr92
8tnCmlSGUPfSexvQDyzfQfF8F97k0ebJMzj2njGrl7wBbDsdmHSe35UbEynnc9Oy
0w2R0RkpiSIW47TjJl/mXyg/Se3SRhsy6bLqLKPF8c3sDu5bZQNBWBfE66CCpX7O
yonQoZFY9ZEPhPfZtwAak8EyIrVSI/nBKHbB7D2+q9vvYR/mlUNoUvBiLYoe2Gok
TPQLWH42kBcqhhnN9VqImEcH3kiDGtpYbS6lmaMgWrrGJMZaOF4hgsrLJqbAfuBg
bA+Fm75rtQYGQ0neKGXiRKVQOay9JP4o1gjMK52VgMpMPcnFaavWuZbRa91IR/2q
e54dAMWcTTCtYalSXzd+bjBUzwh7T6KwuYQVDPQtwBP67ZQgR8BBmz/qG/iQsMUu
dgKC+FBF9WIQ702bCDTIemsE1gIU8+HMg7yQa6j2rl/pIt33InCkCDXUGEEeSOEX
N2WSwQqBp+q09QgHx7AQFcKMJyEE6XV18/V8R+VeemiU2145isorGY34e5Jj0pc0
N5JHnQJ7CH0AIJJ0r7bQYK3KDJG6WtFqkRCffa/aqyKgk5W3dfIMAOJDkgkf7YwE
3BYbwMCinW6nNAH+kHaFffOU1heGVJmjA9YaRw4R9qZxAfKu4T25BgTpmVam/vR+
zEDYy76n/vrKXWHVeKQZEb2L5tAPtRI9pmYnxy1vNm55XXKoyyWIwzLFHeYzjVaE
DTCKgJB/QF2onhhPtqChFVm0vtyXIniD9aJNurVWWOcX1CnH5A2x9YX/OY5eC2TD
gxFrW5xE+bHHCZcN2VEm1Vh84RPhyKrm8jkiyrpLZjbp/1w9h7HF0xjXnNMv5py4
xlCgO34e9Hjc5ce/fWC61Pyc9aEj0RHMmgyr/Z0tx93Sc5j95t+wM2aMetytdrx8
JCWdxQ8s7GP2IN5qRc4BWLewpSWYV0CN68qq4pK3Zy6FeAaQPKoAmrrtknaUHXDy
avFwMaNhpK70NOkx6gKr0Cu2P3gBRdesvCgLc5thRxm4zyj4e+lwqrWY8nLyDe2k
7XKjZwA7S99mHwHWY0fk+nBHQB9RojhjjrSqc7AClk6mSUU4KwO+u3aHPMfXyUtk
izIAs4c15PcoO3jwWX4/n/hx1pfpiBBPzWsQEnrYjKce8rr1Fg0W2YeBFlQWAhqk
+yfD7nNiqkjCneOCsxBACnJBWBqtoQgJE60PKKQ4+2Sztn5wEnu7//5R5+zAyFYh
Za1dKq3yR/xCC2zj688O6trzqHjf/Z9JGuNX3g7OqktTbmGLBA7sLnO+Dd6HjG3h
sBz0GQSj6d6YL0O2BjSA5NtZV1KBBm3wNZIqVAyvMpkRLbsRTbGZJD0Z/G8fDwzd
NuzZCHvx55TIBiMirNfaD4bqxRhY+Ynhe7NPrl4WuZElxiCsG+V1vuoYhTM33Eoq
8ZPAqFW4c30awxcCTkOUlaePK3gDG2c5xEmE7V11g86R8YiTrv73FTMhVIyymfQm
7Trz7dfNUsmbPmxci2ba/k1TZRZ7/DnH8Pqjc9/vlzk6URwnaO0Ybmlxjz4qbUZa
SiJNt2ZKvECT13rZYGD03skKmgMPc3cgzPmRo9deDlj2+TXSCNbV9biysdFetqpC
MML72WNdS0Gsvp0/cSoBnFhyoEGdcRYfvMg/pFRIttTUE/3ZWyB8hK+DwlwsccpS
dQusP/5B9cEUL70T3nWiC04NCloCnNGoMD0KjRNXGlbtJJvmr/CnbMzGl8QXDhS5
c8PnTPKYaFZgGkqocLhl9xpFO6MuYMwaJY+YqI9Vnlv5q29XHOrVFkC849KOChIp
F1DhGFYSxUAEZi0SmDPJwJKSDjy51Bs0BhvT8xMhLkiA5wDR57iZ69kXOFhBa386
+xZ9b4C2T9oOo4L1jcRsJu2W0l7MbuLhTT8ZMcZ2U8kMrL6ItLEXNB4S5eKtXc0G
js9zc2TQZdtbExM6GU26wrvKJ9wGWcYn70/qN5gP5DMZHIj5ToPB2sBAKR4M1agm
6dXjEc6xuRvgPGbogT2Evp0X4Ov1faWz4rhXy+Bog6Q1/M+QXzzMxrWlTgibeYfw
ZTXCeiWBwUH6jZWUJ7C7voi4/V1zONS6EQwDNUwU97YA0+oh3yqMwiSKGk2VY223
vz0lvIQdK4WM9Xud1U75yU87m9lvbtygavepMSe73q0+xfP/iB3aIejLDECbz0Si
Z8sJYeIPI7FqhmUyJEdvbOwxgHF0N6boMhuCEmgdGbnB/Hvj7/0Ex1KxhMn21NGZ
d4GJI6VfTOSD/gdNQfEu3yxBfcWEZGLMX3w1USM9RGcvx3T6itT63d2VscMPtAjf
K0yNYqGs2m56vadoEH+dcmSAhIRhPEFHh7h6tTzB8RZP0mRbePrdPk6aaPvRzLSL
GL0Nj0DWfty8CrXG8MA7uxE4gAKDTO6V7CI+UTMBgDCpSeN02lL0xUFAKx3ERp85
mgu2J7YNScVQe60LvTBLT4huPv9VuzvOGETkVOj85jfDJYvMkBlnemyq/C7Gk7fN
FujbjbVrY43GeoZjKs6KAEOB6DbqXckMYTskqsbac4OCwA7llOBtLOAf+CDTxtEB
q26RwKN1lvDdswR9X+nLJrfs0Rac4tVR1hSPgwCngtNKMBOG0Ghfxa76bHwOSJ39
dITs0U4zIdXpwUHk3FTrcRnglEIUfaf3Lvq4XCte7+dR+e7CG1Eik6ltw2+WerJL
pfUaGjNPkVrqZfjEGH0dSLSb344Zv5CsZ7sigKFy2KbGxxgaHRqU60864fDXjYA4
Ef4R7TRPkJXoWJKjao8hsfdTSzumzz8z885aog0qvex90cFKvjDFEBIt8U2oKoAW
0OFwnn2fxjiGy/7NqX4rm0Ez3ufUCG6QtSFYyK8I7dYfgkKO3zPii3cgJ1xOuiWX
D1Wky08GjoocVNK5wUfYpTTg90Bob8x/GHnOEwaO+uD+gPgD0yIyEqyDZjIWrYPg
rc7YvtzTnlcfpwePY2/qeA7zU2tKRKJpmjsiAWdX/L2YXprYe80l9khfjbMY+1Dq
fadbMJIOCudM7T0ZSFQz1Iga2j26abrX9gJX9dL7yH6gDGSBJE6igdAJaf6tj3cH
uKPoXsKlz2eVLvkTRV71JPDa0kmiEsdsHG9MqqfpeVU71bK7ZBjUq3gCUbM7ZhfF
DLeAQSU0wLS1FEaekuwlNViQXVj5xV3jYRO1NxrvFi1i6T93VN3vg/JWo9anzCuH
W12qj32TCJC8lnYtb/NkUQGn7s/FF1CBe10uoyuLL1MXt2y+rxOxBKf0V9wTvH1m
5GMAg15ANIdJUR7uGRuDAWHrzNKp7ZYmNo3hQfMuPImLVIAxFKCibRTigi2fiATx
kw4K1sPJwhiRobi/boZxoc/CL2acoo8p0U5n+P8pAYYhr0rvI+2pokx5DtC2dk+F
qLmPFFZnhqGG+jk8+gE6zZwnpMxxOUM+ExiJPUCRciUPBzYpyiy4aaWBfaX2I2O7
p2tiFfkguae8PMGEV8+k/Lld9kaTAn1uwvJzrT6IrRFm5ET1hBCqGueN7JEIGLWh
4qq4nShl3t4cknPdCzs8Ap2kivZJK+8C9N/vi2JJhxgBVzWLdgb2s3lExYoLdoEJ
OCBO65Sf3I8smoXpTDWJmX6ouFNi8BIhS084JSqm0tgETvYWi3I8a2aTl7MFhENb
uTQ+1AIv+VI1I0dRpAtVZFEUbnppqAv6bANTU4L+A+hMALyz4x1+HuPuvbEoj+cq
vYe6aUuv5l5G9NJqgKOkz7hfcxxY72Uxp0rKeeq6XkLMELUi7iN7eFqYLQHKikkr
8qcvrfL7SwL9GMrHNiLaczUcv4zrhr8qoijs/6+9C8pushpYkOBkvMKRK6nVhUX5
vbI+2SenUz31t+dhsUz4TUzjGLFMv4Xzz0eXBi/1oYeorzgGWd5tKYAUNHDNk2U7
AV2Y7Z7rKp4v9KF7T/WXwXmEaKjhk7ogjTABzsJZBWh+XRmkpjXOWRWuEDfZp93f
WLUcQo4uMM2oRsBYZcZacoReHxc8UZiwpEUAbWqgoFOy7BUePtzU8K8fgUagZyDf
k8S7y0Vj+w0PoItO+srmYbKii//SGIbdniY3uQpxDB7uMNajGNwK4bH5qQsdcr1K
UTVM5AmLHV3GNeBkm6qpqHmgmUD0vaXIPcj1W9XqIU9ToQE0Bd1g2NqBv/wUnAQS
929e42HvRQS6IDwJ8US5V7Zk+gj6AXyiaDsShL6OTAkIAOs8Z85YTgVoocd5syAm
ebyOF4A5IVBr04dzsnj2OehkVg3AQoPzfeYfVeOUIySrnYT4eDDO3TZKZzgCbIpi
iTfWZ0n0KQPuMLY6NFsbLVXNfOyQXF0VxGEeSWrY8I1NxF0DUf71PgSVD7U+m54o
XmuRjG8m+/KXUj24xcRAqGtU8AOOS/Av0J806AAlz9CszPiGQC00Rm+0ngBuyIJ3
Zy1K+6hkAL+NZ1hWv6kX1YosI8tmCFAlK6jfHIMnR+carNYl/agXJvQPA0YPifd5
PQ/hDALeCyd/ttLY40c/d61VYZQbz/zTrUb8q+bCcgqPysX182gQqTRujv1DVkbH
UYY1q3Kp4LO4f0UfxVWqV5w89CUmABRXNArRvWnhODS2ptcWmiTLrmaT0m1mkYP7
sz7X38OXrmA0dyetcNTUil79pDNcCyh+iC9LGZuwmag+0S6YlR2SJviGBI2GekY3
G0cOQRteS+Y8rlPdelnPg7YbcCy5xn0XzKXv4GDEA1bzKyUvuhnw1+GEu24BwHVs
bi3BkcPus6qdLyoRF/7AHwXCOlOKYOrLVwmVzRc5zOR8LK0z7oqg1uc9+U61KG5D
SlrZgASf10u1D+/jeiOr6w7HIbCmmQk2vQHUYLYnRFf2TsH/s+qgN/ixdAYahNIs
HhpbIw8tRUXuiAKNQCQc7Ai5SXmsYjGLoAFa+9kcFyWly6wEkAhgUcBwngkCxDyL
EVmdBqRSi3F+yJp41PDyhSU9MYdtskCKbfHvfAd7UgS7thFKBr/W00RlptancOTV
QhrJN80D+kdtFJAXbCbmMxnqOdrc/CDRPIs11ZmgduB0nPp5wtuOFsA4iSLj2dri
h3uywfVE6Ae697WUHgHqxK5PzG1I9dffZEWUl06L3LJvkPIB+YhQqYd2D1BafejW
rWfcwbaGOMlL56+YybPmzFAb8vwaeOtQj5bMDe97erXU1wYkBoCCfeUkxSvugrgg
mWPPO2OKL0x0N4Bjzenqz9/qlgAYEsC4Kie1zFlJlczwDFD6PDb1+xF9wt41t2EE
ziAEtqD1oE6Ezr09G+sydCUUZPXxjFr8SzFTYGcHv4TJgFCDPFJAQYndu8MD8cg7
Hm0MVc1hPFfVuXujzXUD+kklbC0I7TOItu9UavnznkIp4+SxYFi+loi0mig+yGxt
aF/sX3I08AYPIj090ThkzprF9u38WSWxZI1ic7hBstH8qBInNhgKsnl5XjSmvTg9
QIKUWCoSdHflwMHzeCH6EtphPISN+CBrzWwqtKTsVW/8ZcOpcgfJhD+YoTnC3udF
z29ettRxqKA7UBwQz0ofFYNCJk05zZWIZeoOEToHPUsPiUmYghVxpJ1v802p/Bxu
XCQC7fv+xpN64qR1V0YO6nC0rBESRKxU0foEc/EB6eB/QXiSwK+oCnWckaLtKtuF
lL4vovVhPSBKo37P4y3spt2ti8xYYYJ4pZIXFIxfgVGk+isVi2YyRx4lTKK4Dw6d
9mF8lBC8OYybjH0ixKr4VnIwFXsr7ksjEFsGc5Ntnyn/Twk8fv8wzIA7e/FtGYG0
EeFcfOhf7Nad2JECOleQ2JwSeo6B3d75UedsrZQL/XGRSHVphdI9EGxpyrbJ/7a+
JW/kVPHhj/95/HecyTmkKBacT5pHwajKqFYBH9kKiTfoaKsSoVnuAOdew588ok/l
VQ1k4tApq/ytkleFYQl7G3CdY4igwGa7r7UnYx8993hf5qcVQqiTM106xDyZcM7O
PciwJTAAFuyrdjAxgeUTxhuGsfdiaCFbVCJBMTXEzBYfWZVaLfVA3yoXQHMvg7Su
sreuv4FGpSZ1e3Ga+Qx+ThEuAZpcA1FFTULgQ98tDR9e6/cdxJSSvovzPT2QhlvV
dfWbim0NJMqWUoFeMkURTLNMT6W66XHrBDwlhM/rYeYofP6GYoXJx8u0RG5y5ALn
1zQjCqQrJdSxFg8cP04VFbUP38uI7sakgD1pRFmj01FdUH6GrbZ1ribb25/cRwmC
q9+7dzSObffSjsegLKXuFG2xxxpFCRiVrI1O4EjE/Y4/nD3zRBW+slKdLvEeZIGJ
9Jiqx2kSdEYGnR/HkOKkk9TDbd14a4z3l+ExCP9pTrgi8Od042eSYxqyDU6OWs+j
28NheYryT0N9iVmbCXWf5Ra8cieW++NfTGXKjybLhKrjDKwa9cBJUEXVC0ZNnLPc
rwCVfIqu3v0xeo1fobQQo7fp2AslESQgIKHVjXKdBDogYRW6o6yi6hJUdCLj/wNQ
tMGZypch2NvUZcKHX8hJ+MKknMjrryoebPgOh0lVeSN73fb1MNUUfAPUOou6sS42
T9yLBYqAr3fpMfD7voHKz72RTv3WRE67NFTsak1Id4Q7CimQjCY0D/byUtA7tVqz
J+sQpfuLTO7k/DU9n0wvIBhQgI3BsnpdEgXUagXyCzRFZKhi+9cFoTnYdqq5qOam
/YXZ2TNdmGkrx/8x2BSnWWRmyWk7JZGMT5leuDAh9kP0pvABNolY3oLQnkWW7phR
nqvMU2Zihkl4RUM+8ApyAbZNDokArsACjzGLgA560zT7T/sFmozbRuI/wSHG0CJq
3Pa6Tpi498X+hbNsmh9NnRun21dcmRvYclyo9ur16/VeJylznnt5JsaGMnymMmSi
JkLoSKjGOJvdvRnWhzNtLFkj1pora29258SDJUBOQzIiJ2IMmZsoUiWCT3w/Q7eG
aCwEPoZlpp6JHGip0oI8wqGrtHMPUzHqh5LYV+ZexR4yZdX0G6a/K1d+cKzfkFwR
nwX/TUXRQ4swDZZ+dZ4jlQy4JZdwP1IRmQo6HwAsepQ7ezZvWuEATurVNhf6mitY
oBJZM4HkK1cmJKLEyt3vVZDDObCfgfY8riHXCJqtB0CiOvel0oDUrvgLdvTemAC6
02j2w07qPAKVw/tCsIbuqOb05cAtGcpk6IMF2dkexk76CEpslb19ia4Aahk7ebB6
EsJAP9GL743OlUZZYmO5EFE+/wGTdHWU+8CnqBQweDaFL0clJviv4R2ZvUyXJyMC
IVPyRQXRy5PxiA01eyWhhdFSrcYNpZQt/P+9N0mRN/NikfXUat2crgauDd+2xd7V
6M+AzJuYTo+YPqjGcP16eH5E4mHTrSdwQrGVe4LUGsWGZWW7nUU4Jty6AU39CqRo
4mv+WqTC77wObk73wz5T3oKbIxh7bziGF87AXt5sGaDTzVOcCoxP8zkM/mnrVjUG
tiEdaZaHmk3WAGWhaqDH3Vri8/Qt3Htb8yqe2aAlU9G4W2Bts4E6stCclPeMIz1z
CLJlqaB2a0Ah6M1HGEOgcbPz7LXZm5msMl0L2dHKgsDzcFgRUsjGKJJzCCRQLvln
T71U3vpDsWTC7KxVWy369TX+rQd2g34Ulksq02PgrRTEyz8zA5TT7RTQYZOaXuDG
qM34HgtGEo66eiqN0RxCQvwedESEwx8DhXb+3uUGu16oU2cKQbSFFXuXOSFkCQVL
DDyF0lH+zOWZSwYWbkmAX91IPyT+K1Ogksyuj9h+xZz3cVLnrFpAygFQVhu00FA9
LF72oOQ3CJVo84PYnu2ZTGTFoayCuX+vAhGhJhCXJUZbRb6L1fTbhco4FDqf2h6e
bn2vuXYVs0tfPHLen7s//msJGsZXPEfx7NayiAPoeAZYTye7e/A7wzEsvbj0kRtG
pJ/TMXiqiCGDiBUUf8bILeQf7C25yoFXTRwNyFvMcK7USUoWXLbGIKnHbgZl2jPy
m2OBD6wMjy1OEC6zPtjSG+1opQg0uAXTxwqUxPRWwKPzF4Q/egCLxoOK4yxm63hC
CMfzdlKgt088I1zoqfurXgk37EIRAJwMGqYKjv+rOXbcgoKfgitOF8aCzPBXMPuq
C/k3Nweg0aBwvnqt62NkqZAbuxMzMcrTqISMJlQh5TrcAeetaA7t6dQNQ/dVytLY
/C6xOm9vBmTLGyz3Z6O/QR8iR3eFgqX+XycD7F9MQODOEZk5kHk4w4XX2/vUvKtl
F/J+fFZGNhClpg+mjfXlAtegl9QGORKQhkmY3YBexxzs7QNk2JO4dA6rfpJkphwA
Mdsajx4ejPtC6GReyP0X5c9EdeedNlJdigziuXEx4J1o5zrt3k9R/+4bxZCg1bJB
eQ3fgh/21+sQPwp58OkSVjUfuOS8yl118QPCyrP7tYn6Cghu09/nTVqZ6YD3CXBu
G/NPQC/W2R03t39DC/c5fdx+0P+s4y5WB26eGKUUM5qBKPuGqIiLBfL84TmIMy2K
mvpS+rGiCvqM+HoVadafIiFZdi3i2mkcdxM3sy4keD42HRquw+X4BwNGbf7wBcMn
2e8Qsa2wmk4U2BXBkUhHdULXtjJ5tVd8vJg4sMu5wfxSK9QurqvvuoPFq90yERCo
LDZDz97PP73TblLPnSaaE6Q7RcSHjI7cpBvakmTWEGJRf5gRKQFQeFSrOnp8pgsT
PQSOnzVKZYQPLYXZ+9YYMNXOslEr+2Z4TNKbLCKNuGgEmoTgtYHIyrzQW75c3Lnj
i9OyVdVj+Pjeij578opLnPt6EWcKM6f/Qs2+G2WXtNpIr0Hyn6LWnLWZmFC0rZG7
BYYO+GUTooBiVGkhMMqeVSu4X2hF7hEutb1DOg3TENf/5Lr9HE07W/NzN4TxSj3N
yGwo+AzOaWXTGwNa81UXyGqkwyMFti6RGQVLWMfJSAWn/m1d8moHSjRUoUQZnbkB
KkNmCVRGGXRlmnGigN5W/CMHxGDqYLJOqlyF+jTar8QUs0SoC2qP9aOzx+TYwgGQ
a1yqk2fjXNG1WJS2Tu/TpRnGu/J8UB5ZwBLbnoHIK8Vv7Xn8WMhNn9ClwYIhmjTp
XExoS7bRSpaA0kk8zA3atCW27Gbl5XDX7aPeFmmwbcvu6J9GMvxr9BX7pT8XTJph
agCpSF9pRyxZfF+4RtnXp/l+sjXmGfbSVes8ubv6Es24Q67UoNHANHV6zj2pL9gv
NOY9rPHo2FeRS8+q1+kNjb7YMD896XOwLmhoj2yOlgNzWl+6e1MQTxDYkGmIE3Df
kbtvGs4p3qjI2s8DFeuUqo0DDPueC6hMaHhqwJmlEPZyAHl8w+5owUW1k9aYrpGk
iENtE9WTxrZ5KihPKsdKY0fYXyFOPAch/c7KNa54MrN302EfFB5I34kjclRBhGHq
sPvdsQtTi6CqnIWHNNbUJ+8P+7rgsP79BGKUmxkC6v+wk6gcDmhhSxC4bSxfTd87
pUTxP2QknAhC9bqCQ6M2/0IKxtyrU73UZvMUnp3rZXuy/NCbKkn45U7E0yznZwyS
M7SyziZt6W9Jay9T+Cr4jCeKiIsQSvVSmiwl0Cms4dWPtzWPHu9xLeM3EPzVEXKV
T0B5wpR9EvWYASi4v9Wli69hX7J7SkfYQ/gL3Q/xpdFhhk0g5Na4SVI9e1v1vNx5
pGKAbaQi8Klu9ij41VJI8Dg+P4gzfyPLt/EzJxLSzylHnQs28MbrWxSvXlOkGxhS
N2jkKEwmUIqWbjIHtAyFy4865qZ8p9cpEXS+GMq9Jn4OGfXoaOHuVcBmkTyTtO2P
kdRrx+sE6tbScNOHn/BSw0WUPnW/zY3LNruKrD1dXRmHraCNIA/b9UVKZc0g1gOS
ib/CL5bMhdGC+3SK7AnQ/CZEpeCSrDCSgMG+7uIjzHqjZ0PyWPuiXIUl1SF0I6gW
0VqWo5zokADUv3cxvLqPnzeHXvbbm9snGQ9Ixxm6G97Ml+tw69TTFVUQDwWAJcaZ
KbQ8DidcJkizS7GnjM7KYLh8Ungvem8PErGdOC1qo0Wwj6x482CrqmQ3PZvtagp2
fNxGEqKjpIgAqoBdodAySGHSNKcJcu0CUh92EHLRbvfPwlxuK04J6UPLqw7AH9Uc
GKguNZn8CSlEdDg658TYngr5Vv0bxkG7YmcdEg8OC5fF0eRTJUfWe/KFC4OhVPmU
ijHVU9NLliULDkjRlBvzdRHl0mlvqRtU3WROKt2XOFgQKUWAUAT13D4deseyR3Yf
wn82kcYiXJbHRLh0WRI7wGTjqkkKo0h54XlKe4STJspOGzmxQNEb6XK+gs4FJff+
BCceKLDX0Ih0U4PwlZaGQhpdv2bTpKxFaN3PofOkxb39otvCVeoYNol1E/bMbazF
oxuF+VoWb4LRZ8gZJ1mbj8FT551U+SvDWhqHEZpiWePdWxFhRhKHKanyFcHnA/PE
9btc9T0mO76o3FDhr+TBUNs7jRCiHVoPL4SfnX5+FJ4JIc/e8aaSEVNEvQD8KwM7
v126g+iNaHjeL+DupIfNBRv3P9u50RNY6BgawxumURwt5RdgDv/f3AsNB1nbRQMK
gBaGzV4y5KsEu2jaE4vGh4Y7KkcsS3PyKC7iMsN8aom7R2/zqqbTkKv5w88pXR+1
eTPTkHm0yQNNtGEuPh2rj7QUAIEtF9zYxAQjUv5De6wz/HooTQXumpBeimVxilzr
IcVGjsKxGRy67dTP61IK/JsMQFTAY5Jm48rl2fIEQPfqm+Tteid0JeF1akU/PSMh
q1H3QQe784ldAC/P16glSm52zFGNifw7j63eADbZxzebuNli1OI4speuXbkaehXM
tdX8x7dktGEuRe+TRqi+2RdsfVlkbV0syxBznHU5MB926Cdh/Ir/+8TdLBjryefb
5AWYpqg8RM6MaxKbHLAMYUW4V0hK5pAWSsSewy9htOduYrcql3/3gR1ID2TMfifC
M9U8JO6RjYcjCTBUWvBUZ3TwRbj95jGNVOTO4JcZmFBO6+ccrv96j2e4ZMUzyV2g
xSKWkESrvtrecE3LqlPzdMKU/WcpSZif0rqo/BzA6CtTfllomR/LwmI+Pd5lbYHf
rxrV/9KftvjIEixjBwml4WXAxaqgQ01jsTSE8S/qNk5hap5bjmWZdqo3MWwk+/tN
2NBpLjJj9BLyQknbpLPy8+Vbe7N+SVbX5TCkwmy2deTQTIVB+fCSKU7kBs2KfxIT
lVcgRJjK6bC1vyNLRN2e+1XWFcSr0ubd3oLDNVzRQ3EdRiJAE0BW2h2I0GorrUoo
p4ihOuWmsJ9GAl/93E1NK8LLwhcRFsd/VWCRva3boeDDNKoKfF89dlzWoaWXr3dq
DAlrP0X7JAD3ofwO50nexVOC/tSeQNIn8aAUPpFZvj5/jNJyGzet+XxCNTdZrMFr
wDd614V9fCzEAsZZu1+oMPS5jzFvdIpiPByBfSA4IZr7BPx7vd4yZzmVMq62VwC0
Nn1O6DJUdyPvf0gTIgGT0MlcKDeH9EuWIWJzTcTg6zqM1uJRQvbvsAq3KlS4yjDa
DpCVNe/SDk0gUQxAKixKX/jFD9qYhvN+AdIF8z6AASnoeNfiH3hHFusDvrp/3NYB
xEhDVXMCYH4Pw097MxbOJzmlpcyOFvwxoZhOCXyY6oTS/7i6S9odOZnn0+zgw0DN
uwqLlyLXkJLRtHPu7jeSoB1c/alD4dJKU5ol28egbhHe3BxjyX+jubaXewoLwvCU
TtN9B02zw+njAArFNccNgnVWj++A7tr42U3pzrRCy0rHyhCdXidNeeb4sQHB7554
DSFiLprzqoTEdSef8kp+5ULvjLwQbEqMVH3IPPa9wBHbKKVQYHujZH1F8TW2PB2u
1KqkmXbT68rf8WlrOrA0rMq2d02MxL2PYpL+k2OXNrgHbuiGHUUfzto4KT8aru2r
jLrjZZMrDpDL0ASrpUHLnhp6W4igvN2llXHJo3hj6BrSkOwSKGlnlzzDhDREeT9M
TSAmj1Ccr5v53KFFi4KmtEddQ21c2UzOzBFyxKgrfrx0kk263cRLsc9WW+vG+WRP
zt0BwfLvXG27e+zHMiRCIHFmMbCaVclhAlTxgB1EYV2rNeS7G7EvdkB4UhJKfFuY
YjtfrugF4GKcmQkH4IvdZaQ410/ZZCFzlh1tJex88zkUW5WOjXzUiERrGbkCyIQs
THYyDoVII6E9lrgMR1Y5mO6iUQZn8qH5uBo0kz7paiH3vxQGI+hnVuu8599NTHfQ
gG+wYOdK1tkZQ5Ds2QpWpWLJjZM2k5xQove/nh1uBuXpa5ybsoEIJQe/w5e1zIuK
XzyPGo+odXxt3dYkvt7cs9woZlVlZoqljah0rl2Q9Wv0CdAK97KE6tlBBwygvNvj
bXL0uHulDUd6wFdDfc9Mg2hZROp3xVVt9qyJOdQ5huXscCKb7j0+2NyIHngNypjH
KwbM4Qs91pmK639Zgpzk3Vleo4uQ3Z/PfcneRuvdruK1p0AEX+OpbEa40MTuAzMo
yPxDdWeMIm9ewsLnB/d4Oc1XuMxycxmhOcAoDJMHgvX9KWb4t1e3z2Q4FctM5luV
00pHUkMw5oLa1LjDLv0BZ9O/TxiVpdfsdm/vBm/qzXI6X6cNG3KhA0pZ9CPEZcDz
FP8lRqKgU4ZxLx7bV/q8b7xYleWormY7157szllbMQsdqMKlUX6XQXBuFKDII6Jd
vJikCzpbj4+wSTHbhUOu9tiV2Lc9zdW5zB2doVKadu7HB0SmBNvXaaX9EyfkKnkc
yhn+61/u7vLHG+DC3f1g/1g7rj+kEcWsIEOOj+JRQBd1I3sB2FUypDgBrQ0rQnKJ
wc/EeJiJRkZWeXJHDMQhgUlYPCiH5JGZkFWzLyBLMC4Bwhf3jQc4rvlBsYvqZvT4
pBibUiqEQhiI2+p7rqDkA2gV0M33saaEh8aZA/P2BgF4gnCRmIIzNjiQYT8IkNYb
R+w0UXZMeUP/sU1SEGVqjgADlhtnoiDCFMyBEeeDHDrwHZ2L9kFnhTD+AWw2px23
iErauNahA2Az3F4LxxpSSIP/zhy3Xsc8ZO7CToBNDen98u/75FU74rJo6Vc493PN
YZeSKNf7GVVo0/oJevB4o98NPHBeiQlyUOWdoawoTyyfcyrVHvn1dPF/QzeTmJme
FG87hm/+Ka0ioJc+tCaWHMwcjKqZdUa5aQinCFaHIR+dvtcKDUA9pe8bzMDNknXv
1e0JpHZjRMyOrH3TZ8IXmQEbepZoX5g51F3Fws3jwL0BDymVcXqWrVu91KcOAluc
bKS8RfxOih6JlokgIvCLyS+CDwa5+YmarvuQvTF+JoSDszNmYw0ofoQhAMda+ILW
L92Zxs5s9i+f3TRlnJCOWTRDZm1Uhobkz420CRTNk+aQuLxm5/WXJSui1GglVHey
6E3o9vTHFT02X0BYMTnuT6md3zqp5PiS5WzmIxHnom3Wm3c5C//eVGgei3oisThp
9Gci4wyqbuueWhGOJiI+4z5J1/PIJjx2Z0rtVinKWg7OrM1pBTQODoyYjTtDlF3Y
Qy2w8ds208Nybs9TEbgWTJXfPQ58l9h1SWAGa2GOhkh6KXgL0oJE8wxk3Xipy+Zb
miJTMzQ1jdpFRWe1NUoFISuaEBGza0YTZki+DRkReAAWHdH9ejzI8mnRBSEI+n73
aaD076QnyOaWkpHu8Hmw4/zszolfC7KQXCAGS5YcklzLN+v9RGmOLA0qq5ZY2PHq
J17zxN/ptZcDtDc6dEDt34RJqKUE37OXMWh1uw3mNezEtdO+CG7YtvO+i8l3OUiy
XmZOPYOS6YJ/fOZTm12aCkGjqV/JJLBCbX/DXrMAl/RNAFm24HYZE827FVpy6j7w
vZs8vgzmt7WoRXUfqpk1Bj20JxZgM1PkcyrXRsMstQgDQ7SM/yN6rz7WM1SCIiOB
g7lFzT10xg4Gun3Z9XW2/xQcGsNBZuajDOuHgTADXgevuIPwOWW/ursdKTuHjBnV
nCT30ndprLd/CvM7uWbbcmYYsb5XsMrxDtRn/ZJfJnqFtXgBzfdyi0g5OXwA8hpi
VMAZAgu/LxNpFZMdFRdNa4knC5Aoyl/xWTmEwa9HNy90Ca/hh0ooIONBGFAJXQS7
kYwqIdLX8jamI7TDOL2aSacTC1WKErUAa+Qfdf3OTI2CPU7RnDM65taCO+zS4Si2
Ko69x9PJU41HU3hf1gQ2aErYgZALCMFk+a98R8GluZEHO6y3mHweq/GXcbRbY3Q8
DLtgKBAvKk7+UCGLOm9/XMWRbYNfapVRL/j9MaCkKwT7abLzwqLqfweBsbqgljdy
+fqxK7tQAuXGDsysPjzBWNFC7DZk/d9u7kwpci0FvAjBmSj+vWlyRrbb4gRfRqhd
JLhjeGTtiiwnAH+H/43JKUTq5vLAGQTHe0qjS7RoeHHhCtvzz9Oxt/TvTbmWF/SR
KIQqFCucnccn/7U/SmCHJoXTvhFkies3RuzlRfIqPcCyu93G7CTAahYNpgUAAcmu
AMvk3zgR3qQaqvnutDblgtMOrexM0Fz9oJpyenaHuKbKbCrU+igeCcTqZeyYjw35
JcobPDL5jlpSAh8fEnanYYvGEYzS5YOKEZ2kC+3clTqjUTgnds6dDlDIcoc4sq4o
AAr2vCw8zxN+GLyEVHMxGaltMtYw2vsMvFCW4o6G988VGWUtHz+cLAUyLhCPfPKr
9NoFa88GFciMeymsbpdew/3NAby3Wjvp7bVXnWehyvH3mmrdaFkhTAk94fxPZ57m
3CrZTrsfncgfzVEQHqmqykkpaN1LtVUmFWwiCB9deJHpfiHOYEzesoqRkwFGYBGZ
ejk8dK0HQzP6i+fhgKVpn+iglxUfLZHAL6XN1Upm2TyEGlYkqaOvBZmW7c78+tcT
lKn33d0bnmF9+8jPtmYGzj/zOdhPQkqD46Q/DyDroF0P76RnoGqf84W3Xz88BqdM
qoEn6eURj8y4vlk3cr/nfjyPFDkl1IOzLvNCfTg0s79aF2q+e/tjpdyWk79lxssF
EAtLkYq9rz4IbG6mgGvTjSV1gOfepkh7sb8HYvcOiweYIRswOlBN5aVUZ1pZViur
PoTvM8yFAjSOhB/wwkFDf/nW4PxSG3sJLAfzb8PI5OPFlHmfbsQ1Wz6ys7R8YHcB
ShTDAsCfB7pSqn8bFRSwJqyhbvGnC6GUP0QblBj8T7tZ3c4rcBET1m5FLDwoN5cC
NnDWBc87yA59X/sq7aBsDgXMzbeUN3Z8fTj8kxRC3QADjQyFpDyM/SKlF9EdivkN
lSzcrEj7bt1XfPoPXFne6EDYhQFHA/aIyMrn/T7zXCQhmB5/45Q0FS6zZoLIZRAe
61yw7dA6OG147zzZMBt0YrUHDy/oyYT2qp4dmkqlkDH137oqPursnVnXSLXU7iAf
GKSRbNt1gR1m3rdCWK1K/AXLpGofg31DxIM3hz07wxGKIF1ca9fBdYVXN9LMbDfK
1KvLONrxP8zGIyK2GOgOjVd7fwHvZXrgNgQEDZP38/aB3VXUimFH6MyXR++dRYT5
+3CfIYPDbhJVqo11FT7TiPrtnInG6lRV+DKWahC3OlkpZKT5ohxnnnJTD5rLhy0c
uYtZXT+q5wFOMhe8uaSsSXOthupd81uGpBewnz/N0X9SbpHgvRx78F6vprKAa8VV
/LawvvY7v71dJt32f+/FjtX6oXe0aQABMbdon4FSCembsS2Q5F13QGtGz9Az1o4u
QCq+ClPDewjv5PvH7SMLsG0Rhwt6nwNs2Cs2ppi5jLtiM7bBIPWZU3MPNpeSA3Xr
TkXpPKtAoYWDbmncTcg4CxFgB7PXQ1609suVBJR15Wz4qboJNfiWc5MaJv2y7hfW
PNduAi5CjhsiAMzJzTtB66x/wI8I8RUeBhxEq0Wb2Cf8+UZoGkpFSm6Uq2YQOpDq
ghp6u5Y/hoQGbEycggx00jhwPzwSJgQfE3L1WPKY/QLaHNycuFJvMu0DE72IV8Lb
XuyqWvNmJGB710o9VX19FRrKQRuu1hy9fU2jaNptVVeqxWVo4IbRE2l8JpXulV6i
4ro/RKmFek6PFCpcmqHYyiIY9o+JsmtYKIJb1SVzlpf7nlL82ZRkJgzgtk1Jbh4b
9dVMTOT3g7yO4iLXYXgO9/ZfmUHbtcvzqVaWWbKZ7F+m8aWykQZ9c3T1E/ljxijy
7Ym/HHbOmVuPfWlGdWNG0HVBf6LMBQQeecLNAqFOjxs3c39dNAmdiES9tBhkqNuY
qblzJojez4S1ZmaVajm3h6NbvVNpAmsMHwD1YaOmi2XDqIXKqR79HFpeeHv1IpNe
+JuvEKHKHCJyVrMY+h+lLRnpzQLycJuoQZqNyYT538bW5O2Mx6Bal0gfT1dN/z/+
PO9s5mTU1rjk5rwKPLi2rrf3D69bgVaxqteTHGNksmmPjrtxMHl6djiZK8tMsso0
UGlK+QwjlVhBr3LAJd0RzQdk6gjyxhGORcVNRGmwQZ029N1kgmGBieQTu88YT369
szOC+W9b6Ahz1Uebl8YRClAPN5uaELfXmTGt//k1YlRFQ+afH2Blvb/k0JztXEMQ
s5K1eZ6vptb5BFyBEiNts/yO4rjxEIq2p6YySwt7CxspsSbeIawxKBwBbwQTEMzJ
W1KMziG/izn/2zikdEQQuFZr26Mwcrh8et5GcuJxwqJQBlQSxqMrHzI9UNNzX9m9
sraf5ZjLY4qKWfFeDONk53gogI8FyHV7EOJuSyzcc3jCIk6tltTvD1O3MkJ1/xsk
GRTIX7S7Z9JJ+WzCx2Cz5e9kAFQ54biTWUJFxL6CM0oV+M7FlX8zatHlfi1HQEJb
w/LO+XepR6butgM90HmsTNAMk8EohIJIBdI+VqftT3jjJnOyO62uw5Zm0UQF+bDI
nKNW5hSBqFed03b29vS2QZwmvCJufT8jRqS3Q38nPWbvQFdaH/ot8SwHOYMMA5YP
enuXkrgW8zAGQti0d/A5ShmHIeHorg6ENhtjppvJq3Di3sDCzT1qq4zbx2mC77cN
4CRjUCXeNbAVMPUmO7aLwEpcDRWbBvIaIyfm2HIuM/di0490bvUNRHDg8tNWB692
t9E+DYURTZ/FItWVju7+hgLx68/iKtsTYVGzBj4bEIowJZQPJ83yKLmml13gWQfY
skfyWyT0PY6PK59RkzcTh55xSQsTvYfaa/ASFtPWf/wxYbk5LB1xZ8cJewIg9G9u
CLlguknSz3h8b2noA78mH8OI+y7YwKRu78T4wqBBfjMelEIV2Po1GIryx8JlmW4X
S9NsmW3I6j2EsTb1krUvyOc6LA8dWhhx0IM2rq6qoDDaBS05Qil2+GGCT6vfnoT+
dvtzuWjCINCzgEYGukba1RX1nMQJrKbYuVQYfhtKXEarp8Rs8eX/QyfD2P5gjfBH
btvnFfg/N4pPiz6ksCXN63KDiJnNHN8mQejssPH0ebtq+h1m3RD1tVsP9cJgWGJd
t+f3tA7UcKCxpL0rPVyKDSd9ed8BRlQ7MvQFIubSuoBkDEQvPqi4RZsieaUto5ZM
+XKefOZtUzd17z0q//nq+jAlcywJbxDZ0wJHlUUiLtRJTPHmqlgq9KGOOvRupZ60
71NEc8nATbttk5jNtF+aWg0xX2QOsPzKliGyEtDfeoTXfRceDrlw03juK5D46VgO
tvl6x9rA0XXriqTS2AOyNzqwQvuxzwnTH0rrc5QdgFmsIZViPlJYhqKEIt9vlPEN
RYWB8yqx7mKgT6jDEXud4iR72bYzFKSb9zeMHBB5KZ9KXT8gXSwZ2ZA6PHIguo5l
K2Os5BJtz6667pmT6Of+1pJFPn/uy7nfxdVC2HU47aHsmKm1ZL37kzarWnKKkBnB
GhSWCGJ6brfiUtuws/AHnhsBg+X7GXLME0MSswjAG4iHfxrspfcQ9KxPTBxM4ZVy
ns7xYU6U04GvrsgJD7KnK3wI55Jfc/PRWFL7n5PHuuFVf6tbIeLrwVsn5C3FfsLU
WS+eBA69iRCs04/N3dmr/rTMX+h1bUoflG+wuLaynQFQ3ApaNKO+rgPNURYS8I8n
zDVSrwAn3znk8MQrS4x748RP9ROsdQG8t75FqR7pgTGyzFZmekMJpm6k7JqCTIix
EYfwNm4Lv8shDv7/tX5Pheniq4TNPSTYnfMHj4MdGTb/RGkXvTuLdgG1G0xbTsuV
+B4ZTAk38844CJG0tSBszpZRcDOZDg4BKyfES6/3J27NRw8Y17rT9r3PtMuJisMs
BZpUnVQzIyU5omUlQiwk2V403yXSxFiHpNUVby1wQxnnrFQDb13B/gG+hOyK1EML
c0OQTKVXVXZhn8cAEzpXQvgkYyVxTMSQRchKT/jl91ugRNQgOVWzBfQICYKTf56C
MFdl+m+GZJr5dtfNCjUbdJfLfdfsH8FaUE3QMmtejB9uMkqVOew8Zvc0kKNByaqn
8f9CYBGCQByy0zOLYkt7HHQL2hbYnyr0jYToEOrbpipLStvwQMSwQ2qFqVJQLktE
vzetmTeFIwv+LFGG4dAIW5Thh68fokiOSrJVTpigvh9V51XF9EMTVVOMasTjK4kE
ZkwnBntIbhquDuq6LyZ4iqWgvwLur6QwEmMNxGs2f+tVNvOx/RXekr2yr2YYBoM8
uzAQRO43uwNotuOzuBpvz8clLSlDKHu95Plapqj1tSSKvtT1nGcLBC7rdAJWuOJx
5PFzNPhho5Xy0uu9/kranvj78Eyvt+UCUFXV951F8GD5Q7lCtlm+SEIIyHlL7cjf
dxA4nnyY8p8Q+7XKIf73IaFW8Q8jiZYQ8lDU6uzUoN60qLJhHSlKVzos83KbD4t6
0BuVD5BlItmKe24kyYVYrX+2nab2fjkFmiJcd+GKc4FQpKXmddoCMBcJgujvJTqz
+bwiiYIMnXXpl2nt0JwqVaxXyE933fDyDneUg3E4pOl5E1L4GxLc0zTJAZd8+Ay4
/7YtU/AdB5CpNEpBzbVSxw+Ajyrjws85ESydTK8EjdJ/o9C03/XL5di3hheclvZL
2WfXKgE6Zd5+5rnMrz7sDcFEpZ68CKLPY+sp/NG37CPcslI+k6xGFv7dX2aOPnEp
1Nsllh8+MCskau1yBk+kf+h5SH03bOmg8ZU7cV923ZmyXKOUk5niEoFJCVbt5NaJ
Uy369Cd9/eUBN6lGkmYI/z888cd7TuWgGK5Uu6rArjW1+dqe7RLjb4uwVQLFOeiQ
xxTSi8B9WazStpCauDEHDS/4QJ/c7IIW0xMEan/HKTI5HDTtpTNZsz6ThiOGEg40
LmzA2CGDvvLkwruqGGkHJ1Mo8IcCL2/YqHazRpWwGgAl17R0a+T1dbmbHE7dp4jC
xHSUvTqbc720GbTDX/sIe20DbRHDMymtMZ/b4+wkWgAQVFosXOBm4TbdknBVdzmv
iIKLEZC4liw9JR9noSlOF36to8ygAEMrEmIF4q+OxlIP5D5zozi6MQIEFuk0Loky
Fi2ySm76xUB3qsQ2zdPPTtCeOug2lfZOOuJsG1uerdu7NvcldOP5hd3wcMq0TiE4
R5T+Tt4J1i8QU5+WR3pxsBTlHn7gf9fv9eU9/rwvUr7UPkojRW0ATLMfRDar07xu
8/vUassDSCvq34OOa/EaJ4sQKkOScMLL+n329v+WXvHBT5UvozcawTypqKSfCqbo
AlVWV+irakR4mVMRwPV6TEi0af0uz1lRshu135HsQ7p3VJGxPQ2s7cfO0Ca7wh4T
LW+8+K+1adahkesI1I2IcBZLbAO6O3yUriYRunSed54NpK+QfTlm8+XAMHnpUT+G
Xu6dBpcLG6hvyIM0/aYgHc74diF42O8oIqT7a3eylKSSCUmyB42++8s1s1q2uwld
8HW9nCozn0h3x5BNlxBcGNgHnN3MT5iyUuUOvFYTS4IkwtUVUvS77q4ed2CXH1PR
j8MuUVXCjx4hwu65ZazPAMshAlE3G7TjFpmi4LIBJT29tGAApn+/71hmVhV94OOs
uXyBKODRWvYiz1Li59caa3NpplmaVtu3QdxX/gzIqVKdiBrf/0ZXZU2G6Ub5POzC
K+WQDgIBqyagcewMjpXY0mebum4BuzI3GPC8mgayTU/9skvWr2kNjLr54Ppyctb9
j1IrHFwocNK8yZ3o9T44r138eI2zex3S/pWc6MrvrKNxp+3LUrDR+C/sJTnaaPt1
s4+5VkPWORRQVCXfLQFcpbmb0hdjKwp0MgZ1YjWrnVRWrLdSjpb1jiCB7BetQuir
X482U3e5uVtVi2Rro7FcuYNwr2Cr8MGPRu8+fKEP44Pdk382aDSkZLuqkqGuDLAk
Z2yN7IQ1vaB2UxY0z+bRTKbJzdLWsRUB6WY9kcE5nbdvMO04eVnWGSNce1ju/y1O
vIxOC8XVUwSCZhyXl4D85kTjzBp4voe96/pdLHK6lDSH0bk0+ki5TorHZywPekjR
jkCt7mCYhxJz41UtNmHD3vv0Ve/Pwo82y5y9RzRyI/RXn7Y3BZAOimXhFowm8G1V
/9OQ3DMQICowbjhBq/GzVakJ7WGearGZx4AHMCSmCrzCNlBR/QwbGvjknX4khu7m
nGOZfiT1xVRTtwhUd9xvKxqzD6JdvDLtZJ9svbZ7AgTAuN2hCdWNmcoVKFNIceJX
NKveJMCYOtnmRMPCyut9INqrH4QiAD+sTeb7gGseah4BRTxKdDkiTI9M9Ffa6IaF
AP0kQloUnXwm+6xifOwof3uSaanXvzU5U7ljvlZNhe+eBi6uZ3m1cjysrN2HImqI
HmvLnSVzI++EKTSRcTA+SAxlWN57ZRZjaFss/U8lwNyM0ql20Y0VgC9xhFjkYYyt
/qEyiOk+cFdaIBaSS6j7hivO6AfPmSriGrlNsUl3Utr0mvM26NVTifcOLl2nFYEc
aHSTf/ywbKlnRmb5bwQKuHbIC3FboivYV1Et8AJeH/+2p6OuXacenu1+mjNP6zRS
IWHzLAtOoB6jEPPvNchcjQvLaAKbihE0TT3P79fyjMcLmuhQvVAVflfgbDYQFMvN
P3VF7n3W+dw4MlDGinx3CYPcAwRViEVneITETpW5vbhiqZtpuGJ995REiRsCAsP1
Gq5Nqi3nGi6qoBUC6dW49Ydt2JEOq03JjCcIR/JYn9djmkrsxl+lJljlbxxt+1KL
FTV68krl2VPWd71WilhGyuHHPt/cOoT6/FfThNsaEW/FENC+IoWi5DiR6rlUTRGZ
PJcPmmUjifzh4up6EfKxapPUIy0K/22bJDryabE6Mx7D357wj6NeTAHmNJvQfXiX
R9YY7MmQVLH3V3I2cjeeeKDDrS5UIpLU0DGbTOb20Xgxxg10XU6XkIDj0uJUy3ZU
yfqpbwkr8PdSrEnMr6DAYTG4NldojgCLQSrfb6k3LvkWkUINhbK+x4l1NqE8MmCy
MzXimR5+0khQi8Yl1UKw4GhpbOdSoePO+NjtW7x6i9poKCCRcskQEbhphZUyMMqz
X651zi7n0++KbWNXnSnS1CbdsrXOuMGccPFEkpUCcxnsym5C54oWfkKuOAy9uKd5
NoLYs8NW52WqohVNxvPEkyEve8A7yOnm6+pbkXs3B97jZjmT2Lp8aIBu6ZGKL7IB
JoK8JUJ86Qe0JgzzmaigTzTgk+3KRhE64KGxxPjq0LLCxwa9RXJ4BV5VhwSPEgAH
Xbz2BWRa/92MM6GUmqrXVH5Of1zGuGEFeFTav28PTw8+7HFn8QrXSUjwV0mxtBzf
ttMMSshrBmISWjMFxLj7BdyxGF5iNT6RkUUrpCEavN+0ZorYLaX8n20WIzQN1n1c
+cv12xq1znSXy6NnHaveqD6iVHyCNyx0XQ9QMc+DenHqUvuT+RJ8KZ4r4E9YRpIt
jqeMZdx6oB9JhINQ2P31V3vs9qc382WF6jK3zoIPshqRQbNMpWKq/hL8fXbWFG1F
dVgq1TGkda+iMc8YycZcOAVagmOnN4mPArDIwJsVXT2LBDRueNlVyCPjcaiLXGcW
etCEKrpgUOPHZP+32Ju7dg3Hn4T6OwNn7Iw96SGsYP0efXrl+oGzp7/yQCCpnfgy
yK/TNQy/pTU+a7SY2mEePoSRFzcJ6yANpX+Ya1SEfP7sbNWFnWyTV5NugORAfiov
4b2b65tDR76KFBAtvEoZ+4sK21W7coKnfmvcS0hab7mOO82QwoRDFPPRFlxmgNxR
/jQlSBDHf4HgjRAK3Kf3feiA9J7POVHzoxdL+Kdfu7jSCXutSORix+xLusIldNWE
8hpkTqoMCOMItaHsSvZdvL4T4cbF0T1YHYTNFFnrLTEzEjzuNCCzUX0kyAdRofKj
RiINqY3iGrpsTQZyZNQegoYPc2qPAgS2WO8GonzjdJzP1SZ2MLAZ5hYmJfc7XDLN
GyIRpsjGQ8Axtb5hsoxd5t2ao87wPrte95yeHcXJiaEdivP9VyS0yIuSpYjO5xlm
XBOOCuOczw+PfjAEFCN/CTSpdDe45Pc+R0DGjDnc3HHd0aqdc8TWek7l3Pa5r9rs
U8pBVY2VZo76DCM8CXobgY7YvmWDnomGtyF0IhUukXLXfXaD8VbQ1pvyoZ8KMgFx
quvGR0nwzVagIHBQOWMcO79GdouEMus2NOKMND4ikS+aniT9UBRASyyP58mnJI69
7jqyFpAWXRsgfxYOWsv/6GQLLEvYJdoFz+llTrA7HBplcqUyKqLHCCIBRe/xPp//
2nGJCbuA1N32zlOFYxDA+G7IkuIVvI5H7Bbj47ierCdBUFksBmVyRGKu9U2MrhSP
pexaf9LmO2WmXCEJOSJ4rq2w/Dei8Wulj/osuDv6UuKgWkXN1U5h4vq/NFXjiK+n
+YezTqk9ZzQiER6h3jNeaoWhzga/fTzFzUOY+jse6oj+Isgwz+tdB1K9DxeRqxm3
SV6bVdXqZ2MtuM/5Sa0lZiezYiNVoWRCm8m73VZ9tHwUYnAKjLgNrm4e/Fzo3BJe
cMtlz0GlqiF/Hzxyhjtvj0mNapin2CvLxG/a3agpKb1FVGEMcuLsGRct63PfpuB1
o7G5VfAnE9s/8eMfTSHvKgYPwI+f6ievthbLtwv27v4z/qGPmji3nJAtGExDvGu5
b4DAjtrHxtyomferOjYk2sXR22AlSLnKuQleF/bFgwltXNcqdU+rEEwvc+OnTt+N
6Xi0i35wLA4hinRWx/R60TtuWuIJ23s3fCLnHHjDIQMTULAj9pDnCMe0o0DQrSVC
BG68VAtMmbxBy2x50fwAWvM4IzCA1McxSCFZA2DJ+0iWJJdabQG12v50iWiJwweG
6sORcLk1BASla2vJaRaDLfzASoy5xHLg6BNdcBFKtEPg++FsVsyKW+5GHlURasot
BMnXO28/tN2rCjY5UyGMJHDfeEVmuzvonKC4bs77a76WxHtSGx5RbKICPuRAm8mP
HauIsw2ji+293xGLtcVAw3RrGBgl0r/qTM5gicgHYBS28XRsKyUvtNjPsWkdrB5b
YGzytcLqGD2dMCEgOVkTotlFqv1RnYqEdp6SbMY47QLd65TcQFEyXQSnMJQCMNyw
+1R42FYQRyOCoTqi7JO6RSJxpViDSXmh8t17HbZmfMcQQbed8igKmsBVgG76F3X4
0E8uHFCQXAW7l9AQwBdXKDZNdkYs2JVYwk8h1eYtYYSTsrpnPCVWqwT1QwHJWLGS
v8ifPT6ilTsi8CC7yIhxZbo13ChaH3cMbOibUzSRQqZlwPG7GnMcbRV8Ewm9Zkj9
H45pO4cLBMAjqytuTlpzS1YKmFoOWsxC7NkFwAbEx40qbMe1sk8pjfPQj9D8ycr+
q0hTuzRLqq/Mq/TRmiDntIZiiRCXzOgXSMEcJwLR2cKAArkEZvoo7K7eAueX84qb
I3AsVPGtOE4kBznCl8nqHXaASsbkkfqczu8Bkfh9LA4++x6chlDYHFlFwIg20puF
r3/VZ009V3CisFEYyQlL3Iazs0NNkTGqlvfB3mw0MD/m/V1QR6a3ejKxnO6p3iq1
3FpfnpoAqTw+7D1sU9+9k3tCGCR7jqSAP1ho+PJaP9c+7dLYH/d4aK3JT/u853wD
wMuUMwDqwLoO4IF8+NWYyf/lZMn2aISjhj07eKqjiPCUrgPoTcgxZwXamTJmA3T2
/kjh3XXN9ospLVSeLF0x9TR2e/o6YmJcm9YI8AQA8kz4m+u9gPQaQrJTOrjhE9Y5
iYyAPrst4HFnBQsXTKu9g8KEimEyeVCuK6+F6B7v+dKzSQMtwTiNZUqLecM0c4gf
GlRzxpyrMnzc9C6mjR7GDJPELw3KaLnZFqFP3v6qdOlktWj6GOPkT3znU6lRd3lQ
A9HrQCtOh4JIGt1LtBygaCLjHN6Z8Ja5t/uY/lD6/ys7tMFxutbYFPmf2hBj3U7S
3eaDRkU8j1j7b00GNT4oU81UBcpEZtqd15NgOiinNKWDuUuQcZQ5SZlLsX5V9VU4
kXMV3cJmp5Bb76TW2x3yKi5VieC7hgxW4rtDxZNLnE71uFh6qbtsTq+x6lEyau3m
yGnrFfawfS3k8r5vRdTmnQZdfLqI0/E2uizFtVqUrMQEB8lAMwWA8yPV8jPHPQDO
kvmwZHOgBW5/82G3DXJmYkFJeX+LYU1QdGgpJxCJrPrNTbv/BxRltZ+N77P7+ky5
dWiDOcHvJVET174gLU6WyOzJ1iLDJ3chNDBhu14ZuLesg/HA/MV+giTjrNpg3A/l
D18PCIBme8Pxot8L7CSyTyO1TKseVK+W+0ZlKkimDwtCpC/K3auCROrm37V2tZd+
cXIqvNXq5la/QkfbKCFzYONkShWd4b+xOPUK8tFD7P/RUUXl3sKTsoLpDvkzudoa
n9PtylHkhBMGR2JjhbsLQIvu8jZUnaHWWNzsIgSRWgEhPqEa9m6/86bKbShgbWFU
wH0pAatb3psv3a2H0iepo2zbOcU3Fl7TG9KNThyItNCggXTLrDwxSMqtnSqNBbU+
aXG75pu1sJLg+8OjArm9Uw3xJukq13v8s4a3xdtoligWHbntSNL5W1mpuxNBNU/E
ufaxA51BkWi5uEYK9ZONZV51Z9EsuES/vVhMQX1Rm2t5hqVghi3sg4lRdmgmt5qE
ZZQbUaA0kyjOSyoGllyIgmAtZtpVQr0hJt9lF6xyj/6M5X3II1Ytm6aMzqK1Wp4N
AqjP3gy8wEpuk9YEFUXZoiBBzn/eeIf6fXRn4uq2SSVwTU85R+ypbE7SgTrWULBx
bdl4mKmt0AUe/x5tM8uuVi0NzAZ9011Gn4M2T/C4CTjpUF+xCftufSNirO3+HrPb
dHzcjNTQxXDSVXkjaqTUTGs51+mNu8dNdSxH1LBGQJ/1MjiBk0wMDc2q1+VbiE0X
DWDdgkhitSMtCWk6vZGIZMzUG0SV8BYZdJ+4LRW4vBnA8f/P8BwDS4tnw16LZKzv
0PSU+zMmh6bjTX0K2WrlMMCvlfQM1f1YfA55Bv+o/gM/KkfLbmnRbQ521bJrusDN
iJdWMw6zp23QsHnaHTupm0PSvDUiIESKvvvV+kXThpD3GaEfQGAxhhC4QRfVDLTb
NjaOJLfwLcrvBCtVAf+oG4sx9WAqTkOo342WuABG0v8aDh/xYFfQViKzqXEaHRNv
wy+aCRkdVn32jKLSO6gY6o/WzZSjle88ru2ra/uYNgCCv4g3aylkAzfThQUtg2dM
YWjQV7TN1RMsRVSnLY62me7hAJK+Yih39qS7GjUHTmYF6se9XvzfVoZalQZvezzC
nUvCJtFtwEAi1K0gzlAhz3Y7CVjIpPNSR1ZASjxUrt3npMOlAyUJ/ocRfJI/RB0U
bf9pCDd/ETZMB25CJLeeau5uUVIrRZG7YLcXtDeHeMrYSaO7opyUWBC2kO4IMLgY
ibihBm+28w1VJfu22EvRs5UJ1PqAzRsnMszgu746bkcsljiKEXV7PZFs5EvQky+y
RuyOGgUZNP+LeGztJg6fSlYi8um62rd8miabQrs7hwgW0yFuJ5uYL5cm+zPGqCHr
wX4SxN1XGsgX8f6XuRdDJmEGBCO2RgnlsOVDGBx69rmVCidZQlQDKcjX410lkeXi
7Y7oC3a1RfO2IRd6HJCxy5H4nA1cKdu+K/ytwrmQta5lk9rz9JggAClF2XWp/dZW
qbNmnUPEDnXw1aB/DTLgIdZ9fa4GvF9G3TX2kXey9GntxFCUDbCC8SIsQ6uAvVhT
5ECEnMvcroWjH63nggiPAoe4jBwoO/4hen57nv68xLSw5z4tPUwz00lVKULPb3QA
p3R4jJlE0oOoTdQiBIL+xn+lmIiunycufntqg82t718kGeJCSmTUM1jCcxgOT1cI
8UmlX5mAidp1DLPec/+uw0D+78BKIQYgoySkDi5UzHo4EMHOYBj4Lg//L0dXFNrX
vrZbjletbazBqxI2Tx+fwJHFRvra88ebiaWOgWSgWhWBMAVxL6lNmXD4vqoBL0tk
GpSDgZyUaLMImPvIcVQAzem89DsRa0VjhfXR0oal1xT7plyOorNXp1JObE0rjeLn
aK17Jhx2843UiNF3++MmrYrSLbwJqkEJdx9mig7mMPphDKBdT8iKAuRCfZwFlcYF
0A+sUhKKMNWU3LkT9jOdt1vmV7B0Vn596oHjXW1072JSR0ozL5n1BNVwWAGuTTOn
h4yPsIuHpY5NBoFDGUhFIl3R6+rLv+60OvvfIScYG6nHf3Ey2O5W1hDkDNIdzFBg
IIZ+VmAyOWElfx6PKCmPOlyGwCfSook2kUyVkPvEge4Gtxxlhi2lGUi09h2EB5hq
smjAn3YQACpL9rZmMzl9QBFX+uvs99YrvUnVX/WuuEju1SnEnhOtKcTBQdvDCK+x
hKqSPf+4XZ0lmXXslXCk1zwtCKq89SX/AU0PZ8k7tcu8Yje5pbVfXAldBuWA0S2W
3ONPQRBzRNT9PBVxRlnR/sFHWcUelv6TihOzh9Q+QfpZaJlKCTDGRkjydOw+fpgm
bbILu2kqifm57/6/98w19vnNOsiCGjymTuNsI4vpsluLJZgHRGWC57JRgCbNW8Pl
E9Y57+VEuNs1dlpQ+DDACVSeILqvIdJqi9Ie/iqhgxUSGRJb58jzmeBc9/XD+vCi
CMDNfs3a//wVi+t8fW0nqAFpcaVJPfjrC09JXK11P+oUppIG3Bxf+vD9+YSmIUAd
QT2Aa+jfpJKfrrpmrWnrDBTaJ5027lT6uSr1JH/1tH7DNbGfFj33jJG1LqU1Lsut
1cHlbvNaRzC6+xUUvMVbERuIeygkhWVZOgAlhyarc1fStGuDYqlz1eYOcNgU3eg6
NPcyFG/2wLnp36DOid6mQRn7oAnb9UGFrNnfAJFp6sEd0EoY+foC5hErWoq64X3Z
S6IZhdvGyqw5Pyg9XlrjKLP/gIkqWjbQaCyV0pC8DQK0NhpMbeBNErDKd44wTiP4
nzn4gJf27zRiEdKTxcHej9B9UTy/Qv3LGN2jZxg0Z3lHmH6OlotvyAk4pdVHEUFq
q+uPRNOskjCHPpD8NxP1A57KBgG2G4pZbI9UFq7by7XM0UzO/FpBE+5x7fjLwRAg
Vw27jadSOJkcfKEv0/9MSxJMZQjXaeuycRVBvWxsv6QppiTictVQWSFk7cmYDgaW
yL6Ig8yxh5/TGEIxTT16xVJjeC9YIu5JbL3PDbrpH/Mxk9uWwqHtutOnMGc4jQUH
pnc5K/kRSF1yojjD9fcSdnxr9GlXBQAGzJNOTUeJFZmTsXvLYXWMyRhXffYjKleO
FzpPGBPUCNluhPKHvkz5Ukos07Zi5aZlkntlfp1RQDdyWqHyH4cQSguCtNF5S/L2
mR0EMp3Ne9/bN2Pvzm8CLy/+dMHZ+T9sL96cdA1r9Xhel9ziv6xE3ab6ByRAzRA/
UrR5CTrWV2ilow+VoptZoBoasSOdfUxYq1lioZpCTJeSfp1y4npp418pt4AtTcj8
Fx6PY+93Kv///UwVGRfP0Cq5/c7gO1UjvjAU9ChuOnplJrjxpdoqUnVcE9GXNwum
qxyCCYnglNRwP9iI3ffiJRPWYrAo8aqa2IPMLzBqnFjq0DEiPRWa+BtB5ZxtcOzj
41SqjlREBIK9kNyZzhP+Ea+szJu6h3F2gwIdB1pbhO3S2a+nWbNqZnmagc3OvmEk
3TgTaWkD7wdC3vsjArXNXw5FUouVcOdpANgEIpdLZKGCHg4PR9stqjnrmzrTDgu7
3UqfYT2hN5f3Bmj07av9q/atF2A96Os6uED8mEfU7LOp2htotWeuQ/hCSDGlDRFW
xDkST4Z1+lI2FJ/H7WMnskCPbodBGupAnX6oQRkZpheFTKqNPjUo/ecVrwLI3+xx
44Jx70J1I84llfj01iu3fycxGVBxIuaLven+0/KjQTviF2SwmF24FCRc2aOZ0OSK
Rh5pKQs6ZynoZfUttnF3RCk4ftlHNCodlx3Q85GvpWJfV46RPHVgv2NBcvvIPZfW
HDot0NeEQUyVsOwMmwrzW0B+ivVbVApfw/Tc7iowmfoia6uMSVYeKBbSR4jfSaU0
1zKhh4nAu4w3oyY3uhZzi7exTp8TCB/ogOT2BmtCgEH2xpDLofO2EaAzrH1PLsvZ
/gwuHgIqiWn4Tw6JD5EdnTs5SrJGv4l+q0rYsavPQB5uXB4GfYoI6DAN0yiy2fsb
vnfpsRyLKoGDH+VsgNqETtzIBqu4RT/HLkxLB1gDbY8ybj3UIA4VxiJKz/C0sC3m
AwaEgwepcKoO0D+6DB3K1OYXNfcUZ1yn91rHtmnoL7V3uK4DJe99USyd0Y6Kun0b
BGYrB+EQD//2vTdMppraTBki35wC6YvDr8+tEQlkjh7FdiJZIUh3/MT/79cUCWzp
luVAPqjXPb0njdvx0/gy0rQXK7yvFcTyTOMdPHNn6jGEwVAeh2kv26v8MRokJz6J
7HLuJDnfINzmn4+hQ0C+eUmcC2tR7LecMUlgMTnOvyFGaAYdnjhgs8TTR3B2lr2w
xYC2anA+/mJ3siDcCX7tYW+cBLcBi12XQo+lRa8a90K90tgxcg3hLm+kRw05El0w
Whu1TI6Y8YJN9S0CbNypQ/aySk/A0vhhZzqNuCCrEIITx7z+NMBMfHpFKN5F5DAN
xoIkAYoMvCAT1ugB0qB2dKOzj/AeTr0Bd28AhG36T/vEzQNq7XjONVPoCLUtcSdo
NQ45bIxsI/o6VigbAaNLS8YN7XAMMtQ3tgTqaphcFO6H2KAfX+eXxB4i13Pixffs
UqjCYDM+b9JRhQ5OlPrMz2akXr4Tj/kn81kJVBluz1zvIDgyZEytMMH3tjQyC6Rv
IYQx+hZNCfOTp+Nyh2lK9S7QmfX1eNhV8/o4i2e3/y+DPSifL0UOi0mNgo63t/02
CKGxe5oxPZiWACYzAVZfLz2BVprNg5FmtCtWKDLkHCjvSVs4sPUY4Zututsz1zR8
U53OT5gdDJYyPfnv/xswkYoZvbsMy6MQwF62t43cpYBwHp9Rm0Ntw46PihAFSxvc
He0FcN6jhqNHvcDDpKRINR6AhGPNw29QC0Fp2MwPYJJHG+Vp9eeOB7g8KWLUeFjs
a1Ov2k4QGnc+bQwkEhmxflob3D2UGen7COU0TsMlw48RsXgObCmUkd9HA9bCZj3A
a+UBWhsqBixyl145uY9nxgF+CcDAbC7doUOPUWmtJ79KJ/R56pB/rnmikmcOiRnY
5VUMfsndDQvAwR12HBcuLbHkXdpAgvluy+Yzrk5Wp/k0TO3kdw1C5IvqHltFvew9
aJh+YY+ebwmH9hpqCbZn57J9VI11lUK4pAdXZhYa51xRPnZYcKjrFBzNkQQGHyPS
R9EjQA7UcoTc/4vdq15RBy66decyCguPNxX21ngwJNKP8AOWCWg26FWqz/obB6RQ
SwyFWq6ebNyFi7UQ/GXxjNwY3qDOgGXpEUPpWAEIDgqELEkNv5D3Ztm1EN0vS/bR
A2SVpgFnluoT54ICfNU5+YfRkND0nmtSHJtWu8SgWIylI8MA+ErBwwx5ioljOot7
f7d3v9CSgsvHOq8VUyz8yg1tT+d+29B3x0nEIxhI/xzAjlS81khf0ayZK92fdIdA
iEVxqnj5fB3xVWTk85FCODt9eAfa6MZGpBLfDbP4K6Rhx+GWs0HIdRdqJqE2ZiBo
MGdyn3NpFAXkzOSEZQkCSMh1hPFZu2w2F81TRa2Lmg9AfpjaIIrkQwwOiAVIh1O5
9iQlswH8fN7b1vYl83QaEWq955z/yemyvnTA/ulp4tPawhywyqJ2SsFaafaN1268
MJ8muef+mJ6e6F5h7N5agbKt8riT6foH7oPY+ad3xHbjsxajZIcbkAQzxlaQtq3Y
Dj/S6uGnxO8/5psmFl3ocVCrliALoUDSUn9j0Edg0XxMfnH39ZqZqNHos+4Mt20d
vIqFAhpzQ5MlZIbq+jdkVP8aex632bG0qX4t55sPRv2Zb5KKJSvGcfOEX5f6sgST
A/jF2o/ldwu86Er7FX3ooEIOa2Zs+Kz/GII2WFSsGH3Ajpi3UNL6txKOFBzA1/2V
sbBCK53qokRJ6YvucQQ3/RJkvBYNnKftNcFYF5QUsYCxYjgtMZKs2L1fea6gi0Tm
ToRhBepAki1zzCsiKTsIMIec6QJ6ouJ5Rys01rfRjiD+2FM4ZK/4/6p5uG9Q+56T
NWCDQQCgi1ZBbS5Rl3ok9OmwXMQKzjEcVwxctyEfWCDOfyd+vejeOqN/epT2+FfU
91ITeBovlGfwcPZbQ/cdKgXODTLDtu7BjNYPMwCMlz2GpIrAo7mvFMGMhxDo5ePj
dVQVQk/9gT9hyWtZhDcI64p5VjZfSlPCPDq/ZEJQ6cb7srEsEhN2TkwnWlBCk9/W
U77BM5kUA0zuuJSEfVXJT8VZHcwmMY3zBYyWb4HGIeeBOGrI+KQ6FYcD00dwKK3O
1cXv+qFt7wwi6Y1+KOqUel7QrgA9j4VQNQtpZIXE0t7hxAKi44QOlGjJiwtWgWZE
2x1iPHo1N62ANa2qt6HC5T+Pk3iHKj9JoRhdrpeMLzBpXy8M3/GByUE70gwRBtWX
mIT7asZUO6lSUQq7zt5AbBgZuwHWkZ9qrEcGiqOEYaiOrjwcqdTQqB1CHp4uLBgJ
higxD37b8GentY1S9A370fsIcuJf5DSFMA6Ed3FOw//Ngo6kMz8e85HPQZHtpShe
YsXq5jsHvRrfKh+/P2ZwVdtOjtSjhOM9hKd8o47n4t30/g+v9Bi9LgtyTnnyMCus
j4WbeCoLNbyQ7Frv9wa6/8D8KinSGKrLp7GoP/sRHSy2S2PGyp5dsqhoHkBDG/qn
XaR/bPeImUF0FWafsalK6Kqz8N5RD13jj4j74EB/nZnODiyGblTKLxpsTyxeQkZK
eUMFP3w4ZYI7bccS7OHPLm3L8PZCPptUPMt8Ck1J/EY8bbzThR1cN4/hzdY9f/YT
dT0Gct0o1/n1lQc9SrfnhS951gG+L1QVBHTany2PBFeNn3gNLCvkL916NXHGvlHn
yGn2KfnxSilp119kPLzR2gTGPFd+vOQLbf/mE3FtbFyMhAYxvZX+TuuChNxQY7L5
60aCr0UMt04F/szAx85MQot6IRw/R6KTOkk8LCx5cHg9uXtLYq3SNyeWrIGZ55rH
9jJqGHZmNL31nNGu/7xAc8MdljL9YSd/9jJ8+A4qmhDPEdzKME/sPOS0cf0tawmL
kAuzPG7uQ+ilipipI8bRlmNJZqAsQnCk3KL7nWUtmTOf6cyyxR9Yjbt9l2ZN3Ip2
FjBbXF8LnzxAJqR5zqVw5gq7Yz46sUgWagQ+gZiKRwgRoU0pk3OO9wJXiP5hOCxr
Cyd7SqgyL2xVJu8k7+LQWVgEm+iv2BYLOU8O4aKTVKzMoMnwc1pXFyhat83qmbBA
2x2ypTMNoV4eSKcmL9VCiq8HdGMjpBn22naQ4B5tKkuMIdP6A+gXW43L1wa9190s
zGeL9yr0DVJmqxo76d2tULe18SRV8VGSxYv/iTDUkw650jK9H72lsvMxGmPqBhSu
7M+rRsvmZwGkUBxnYs2S0GNuH7FbFwcWU4bPKyYl6keOqntpz4tpxhM2VqI6pSZu
Rxv8f1VYV+fFdzoEwgdl8F6fyaGzTUjgOgM4Uss2WjmkgD1fwn9DV46sKotkKg3C
m+p5hAKXkyHYN59qVSpsw1eYz0j7s/EwUsbEehaX6BiR+WKl97vKbi/SKArx37aB
buUZFSPIKlnoHiX8CEWyMJI3JRVaxcdbcgwGHHTcn13MnL6zo4SNMGnL3LIMKr/K
t8rmNiQpsPhY8l1mErJJ1KKg7/8CTLeA4KGl1clGDM9rH1XZi8KWbEdtY06v5k4l
GRWR1ercJRXQIkhLpcs9QliHBXVTkX0O0ZOPLwkUhM847WDcPvTBJygCNY0z8S+p
hYkELj6Jv9Qpb3NcXGmnqrbNFHik8ZzzkdnE4u/DN+JnFE1rhFE/vEe9wM8NkP5+
OmWkSowJPveNUQfcDxn8DSBB+llQzB9JkQCdI7SlLzTD5rQfwxnpicrOC3t5PgMI
qopXS4/JK9IWorEVLu+l33UYCPiDB9LOWTLuHg42Yigg2dED7uCaztcXPmiwLlRE
7PwBjrdYo/7NM7GrFiYSSksv2YtqC5C6nUWTEFrxnY3rufGtbZ3+KH7Kcak+9NLT
o8yOFmVwRdReM8lgEpR1nAE68/olsFbLbkDG9twRK/D5Dj8p5GPUnDe1i5ry0CNu
JnOGb+rMdMF5S0jc17PCx64YTfkgmPwRz28iG6KLgkn0F/DvgmhLyYhoMi7CZyta
ZQcYydl08RH68quf1s+np3BaB18Z+ql2LNEFK+dot5mwzXYZwQ/ugApF92gVJwBW
KKjk6WickkCeRsTnHzpNIHoONLeuqQhJ3gGpkfXZcme/qKDQ1kjnakYhRGoU3+z+
D3wt3+uROIwNlWBbdikHKmngbO9M1zW8eHUAdB/YyI+3J0pkgrtzVSIAR5Lf5bqZ
jmjx3mZ37zzbHPMKoYz+yU12BLKt9DFjoz8jwQQTkKP6pQK0qFghQ//WToB46ixS
aevdU5xeMQh92HcpdPqltNT8Flp+E7GacS4TZL4Q+sRL26vk5AA7T6G2VcGSSC/F
gPQIrTBsEEDWbSH0zJPwUCWmuoUhGevB7RGaDgNpRxOhd2weiQ7AqtMltlmcolRv
BA90O06iII5a8LCbCI7M+0t5kMzpHd8kOEvaA1LzGKN0mQN/xRxgwBv59XsrmIZ9
8juM+tkQRIhxbsB1lPbsLdDdFzY8RL1TG1swZxvbY98G15zgbMHe6m3oVpLNWlNY
z4RKq18n3+gmkW3+YL8N5u5wW77DF/C7/KbwDouS2V3S8U94DIiXYe7rm2J9bxwX
Z9OPDHNKXHPtIIQwAGtpjm6JLpDhmHHr91Wr/MaUwgNytXuJwNIp4XXVgUutGH1I
FIB/3TflNd/gaaILLB9biLu6HvJZym2D84DTk8Gk7aEEJyCTMkFXhD+BEOA94iuK
AK6KTrzSwXXQEiCQbepm8IOoszY6T+TQdgdLS7pyGgE1OFJzl+YZ7P9NABJylmwe
+gs/toYjJUBLPRgMwzbu876mQ00KboYw++wIvXdSVVOq9uBRg35V0EkArdnkKIEf
tmsNp0YFfDZWGb2+krp0Wy/yeiOVBgMz5sJY1+EcAiF9QAbeb0PvIxDCcU8YsXFL
zVYJ07aLZ3pw385IxzsSpOlxd4uxPtjdw+tOdbZD87kMCTVvTwBfOAsX5DTPGvRD
JvRnT8+K/M+EbLzCfpPcsUZ/XBBCgWQ7ZqKYbooad7Yegss4tV6R2b90kz4TZjo5
ini4g/EUjXTqeBqqm4M5j1/+2q2g5hz/VZH3ZOhTjwb79/C6Pk8F3s7oKhVqgrKI
4/WF0NY2CsA2b7rYDrfKRcDkvQqYiRYach7eheLo97FJyOL4ISO/UwiBrr2vhawB
IwZ0ouxqV6pw9tfuthXr5fTc+o5p5XmLmX98n479vFFK2iuftg9AwwILbDkhYaI6
zNu6kC3ec5Zi4xu9E4Y5P8pRHfkCYe0i5uI+b1yuLPI3LU9MQG4m3LMXV57ow/VJ
EDKe1inT8H3NIaJT9TzLExsPrQ3h5HAIkXFJsei6J/Gp1yPaFXxeNjRQbyGaHayd
b36PCNfa4BFzSaaoLJiTcNf62Yj89jagRa4WeXcaWiiZoxLKrPo+evktFJiZLpjF
iistI+vvUAshGSwWSgtqw/tUEXKFXzr6C6zurMosyRRJD0LFpGokVUs6vjIXV85k
ddO8UVJIosmcyogkOnXKo3aUW2yQoi6o6gKZq2FYDiRpgRw4Cix5SlhS+W+ED9Fg
9cX48Srnck/BrTYvRZmE4n5fdigrqdIrKKRAxlnD2tZ6VzcPBJmbGiMTsP9zQnpw
B1gXVNgmEMkjoS0cVrtMwemlc6YuL/SbdIBDoYS+1CfrCv6pbtypfbpQ/O+Ol332
s8bQzUimDRfSnSLR00OIEjyL2oMGTzXJToTnQE123AtYBdOeXQGKBMBfC0mpVg3r
nC4cn33r0bn//8AjyTOEJq8IflxQJ6diTkZaMUgTkXizjhCiF2FyUVMpqM+F3Jx4
xxNRGGaSVIUYyPbTTjtTtKlFAMFqkiQHbi8TdJlHxaKKydpm3EZf2i5EkYH3iqEm
vsNfeCZnej9xvh4jQT/1fA72GlA1uNK27/udOkXzIvjseiAzNiIasxoZGlXDWolf
R87JGG1ke2KagtQ9+9xCQrhXdyIBMpFGzvSUgMUmtXWGe8BRfbszHopzwj8hpA6K
hD1p1YjxfXmP56/TfiY1hR9On+HOFoi+TwYCE5pZz/y7/aKp5iUzL3KZAIrR3gz4
+2ZSFPP80x3ALUd33oaXK10pRs9fpZ+G46yhq7qpm13UrxtN6IQKJaVoRf/grfr+
8FF/osl3iDCBUb6jiZe3DZXO+RIrYC0cVErfpie5G1FCAhopuKZbvKkvCxpJYt6f
LEMAR+v6WZpqncTfvP2nKOapMstBkOwzbKyFtJooPBRMN1Nu0qAkxituD2xI/zlf
y9coxq9rwAKSwzUlnmWnywDAjGMvtzqE70Xvun3shzHNMkq3hzur3NmiR5P6YbYU
LKgsZZ20p02sHwMbe0mf1Ms5+j4yokA3IfRmvNbtpWsnEXkKQgCqhkep7TVitMoo
TUtdhiIyTdiSdEqOuDXKHgUPi8G03v+SPQ/TDYFW/JlUYWSq9/awY2DNhZ5muGSP
uygAvofBiIAOGlticQMNW4cWXNXLpxsSfypg9DisUiLnNwUbKciZE0cLJnIzMbrQ
rQgPshUK+C62Mj1MsvKEw/XBZta6VhHHwRTQaeTOTL4KoKEmFjVkPcBMH86yywqr
Hnwy2pgVfyk0sFmZ36ktNiDCEa8SX5V4CZR+WwKfnWOjIkVXvdihbNdTunfOY8HP
ntAyVfAW5Xuho70DAKo0tByGLpLBRqNposKjZQ5SXyFHcWcqA0rdhNHVP49SOlET
PbkNP3MSHNLPbr8fuQqz0JZgO91AcBqIoChsHFeHoON7/JbkXS/82JTydTfjpFV0
crnxw8Ij++4c2RjOleCXoWWQypehvD/Q8uWvutHhagPeDu/ZmhOeeCPm+BB6zx2L
ovWukoem0hkfu85F9+BCk3IqybUQ+FONY7XVyUHQkY/RaFzL8pTW78H00oYGx+u8
/Em9PVU9d4occXnR1llBg7naJ3h9LdEyxCgFbqT1lVT2Gxn4tKLQhRMzvU1s3tUT
Xfq0qi37ozoPbj0E0CEdF63s+4I1JE2MwtuKq15J59HySxjmuARwMT2SyIo+ggUF
jR1HDNdESD22Zrh/GB3nFBqe7X+Ir24DPvYndUCc0fnPYY8IOBHp3g34Aslp5WDV
oS24VQ/Rn9/H+1qhLkNc86kxEMn3DeduxpAOff2PmA7yeGEmcZw7bvu74e/AolBS
wnRIdfLFPg1hOUfWIy73qu5rqAkdhORKhJR7VfgCnr7e8OOdEHsX+3d1/j0JjyA0
jW+VWaVeOL9t0fZAOSv3HqWELI1A+4yjzzC6HfD2vD3HjJhiW21FeXhWf2Fhwry/
7SQY1SOSaXou045CP1+zlcHoLguZd0u1Vzhmv73FA2/O+qOBA1Hlj8OGKlUdh1Al
iXcReIK6YFtZjA91doXpmp79MMQHf222xmsHNqnoQCuzorq9wt5MP98h/zU6z/zJ
aO5b2OMBF308IyNujUyF6uR1qFxu6/2rB9Bm8Z4Wv/UlQx3f+ut6iY6QkSFOPDRS
lCcuMoakKkrb9ElLVirVEq0FUwFLvLb6G1MPDlDmO92pdHfwLx+KbtXzAHkNPv11
/rIkMRXHD5fA3s3vCsNBWLgZPhmq8oC7v4pUirk+3TieZ6vLObCJq69pvT1CKg+d
Irm94h+sNzUEu95+qIls67Xkks7nlzYpVsjNXZCtUnmsyuYVDc6+F4rBiYmxm1Ya
bRw62il9MB6pEdzxYnRLm5EkTqO6a2xf1LPKVPdF+udXhhLf+tE75USTRl1rdP3N
l5WMarsoljuBjKkHyjB/V6Nu8sVTBqsjdS7ufxMVjsJEmOsjBFXhxfZe8Jporemh
A7Em6vYQ+VJ2OVmUkA4E0r5CvDpxZQfdWRxnYVZ0PL4uffa5CkRqtGJzqfj/dBnq
6TYRqwiLN/InRMPAzpVZZvB8Jg2pe/LFMsuDavni0kt+VPyxljers9qzhElJ4+FH
qmIl8bG5FLPFOQia9t8y6vVcVsQ5It0J9FUdTggwN+Ea8nQFIckwOzKrys6oYOHm
fIGm9M+uOYKhmeqZiA+TT/YvTBS67viRmiVbSBAYnQgAYbdYKm1uocdQBybAZCZS
HFBNe6yYgPj+tsya0m/2DmFnr0nqmqwpVkPrGJRFXqBrz18nsFO3BDy6AEB6YXYX
hws+O2RUJ0N7dES3rHYXsS9kWrj7o2qDuvNUWbRn/RKgPCgPQ026YX9BSHFwvS3/
agCl9Vprdsqcid5gnnZD+au5lrgCVvv3uILkCrvlR89yfzFOE1eanjl2pjr5CrUx
GnI44aUTGb5kHleyDkaiL1wZD5qhSnW0uJA25x3/5ltafM0ckflS+4kLBGoUImzb
8we88ThopIa6UgVjHJmvRSzI6JIcZprdDd5ashtlHyqGQokxrrnEOlh/iewA7abD
Q1slbR/2NWuHeuyzTnJyRZHrGd/07vbmkh50r+irv2KLX2THWVPvt8WZ+84rLfun
GjlZW1UgG6X9QbQiMbC2MAvPykVMbbdrZdmSF8NuiXAoXjmGDkDU1GN+AfE2/Y9+
pV4naeiFSWlv5NiszkKAy2sY+BePJAJrKlsstjcJ/Gc7HgdqXelh66W0MyHH8Rt/
5d7tJDhtlxC8t7oqS71MKU3wnZ21k9eCbDRvZNQ7Kn3acpJyy4pBBzjtSjXkkpWa
sTkjgcF0gT2D5vBi9KC6Q5yx5I3Zy+Iw9MfKMPSymbWaRPx29FTYMEqTs+zdjq+X
QO1gbBlyMwPqTH3m8FHghSnPSZwzkpG7o1SoRJPc+6vjC8UErHSydltOmaShTqEh
/ZlN0DS/S7r19b64Ui88iSOrxO0s2Je1qqG74+n7JHP7HkcrvjfIxH9o/wEglLn0
sCdoSUo6Ma7QS8UjwHfXlW32vfefuAsNq+P9BvAKsYYXg25WC6y0KFkldanBdXUV
/MH7CDusMoipWp8gmWHjDat3UBQnAiLm8r/555C24w+dPRTqAVZbB7c6dDqtqONu
eAzWKuDIjKn3jogU8xidAbE4A98mJKLa+SMoSxntQ0uGx3JuSCAVk7bUkebwquY/
bzvRhasz2f5Hc9sXzxMPAejtCJRKE13oOpmrPnqPO40Gs4DNycenyXppaa6VHNJg
WRXov3134navRgU1g2VZK/CvIYdHr0Ov13oM0MdFcmbKRqd6E50vcAYjBOLzrERN
B4Y9U3PgFuQie4JTRLoC/UFkJrnHUz6NvWMuhiHAFZuA/cbZ3OH1wwvKvkTQPMMJ
MbJ1tgRKDVoRAcuISsbVkoIsAKTCSLCLLKYupgzizWxF8WdQsrbKdlE/QeUZ8BVv
0xSpYPUAedkm8ZF/VYKlQenurmRTWBcOeMTwhuJ1s9TLl30Hvvx9gOQIEtmPAYY0
4LHqIFDHtA4HWdbNySEkn1o2HRBhO4q1nRQfVovuynDpPmn7MZ9mzy4yrwXqjUE6
fryn8FmbFhnw6CNnQGVQyFjgIHVYFXK8XD58aiCLuttrzLkhb2SEO4Nsu0Z5DHv+
09/w/mWHrmhLOWz1+hJ+1+mMzy3ur49i4ukW2+U64flKp2M7WgF+crBSvb4WsQXO
T5KKlB9cwv0IiHgRnIweLdWElZYnbas1z4d1YJQaNgo2Jcda6cx4T41KV7aDSRKN
wg8eIGBus/0z2rDlAA3U1vICE+uk+VS4aEzNyxupSv8aFyRwcbqog0FwRt93ImuA
IKNJtcZEjz0riVV/0TtnQUlpk12ouuMoW4e+09P5MVhpDG1d+0dY1o9g77klJVzS
/IpBUp6eMvhqVuw9vkwmG2gW3Mlgd+65vAyRP2Bn0P2gwgBDD/LXMZTKlW7wiop5
E2l6PDjuKkGJF4WTW1gN+26JHKW0HOhTyAul9YOSnf9JGZYy0+48bgdehSn7oEaQ
zetk7WfgVndVJqqsD+/1ZPcow9nBof5cD8IE4qXjBqdCHpgCj7ZpZ9wI6WUsGpMi
o/yYqlDSkPNIpUujEMuEDgDGZfxIU9NdmEmRiMqHR/AtyCPJT7TiZmLI391TIrdV
q5bcwRXKwSaW3CVonMKVzn0pE+GHLRpYYHLEXNHhpqqYWBV0VnUhC8lLpYRW9kU9
ul90mDC2/5105F5a1pvDPqO4t51noKwQoPHnjuaN5sRfJgHFJ5lydJpWtOJHEMSX
h4fu37lWDKfAu+AbD9vQjw3X+xeP7LNyAMB9LthZjVs69lFfnab1gqTwpEC6DzwT
9xgZhMxRdV588meOw3xmgeIA85KhMK/2caNX4zpPWtpsMcPOE2zqHE36flW4IROS
LXtbk+TVS5Lm3utd4KOmnPiI40Cq9TuLBQe6DXSj27+uI7YvQ8auCYSpckcvH466
rntnZi9+6Ta4OKWJhQLuiuk5VAgkpx1hgVZg3z9+SrmhZcy/Yw6QK2BD3xn+9RmC
uiYdZfDEpxgUnXOwI/ydBNbfon2CVPMfNQ+H+msqDGcR7+pvR1X2BCf7qrOrosLG
uGXpV40L/sjsul9XcOb2UmZE8zuJLQj/7T2jMOmjeyhcVKEoc22pGw4z2jqzL0kC
dj9V+gCM0BjqrZWtpCUGkgIgaep0j8i/5knN/BRhUnvC753sTq1zagg1ynD9KwS5
sxOzSVSHcIkh7WN+EIUzZVRJXZoUL08gdQcRb9XDyJ9RN8QwlR9glTqrY4B8BE/Q
A/bdgdn1lxxtyZWfPERTfJnv3WBFc+JIVw2XTObSU33Em9ipqe+LNJlo6zQ3j/nk
Wzw9l9SP+kLE6xK0FeP3hUAio4pXqhKyc9KrYuKMAGHn+6Bnj72gl6DMC4QOq3FA
eQlNgZzDKKDculH2SJVern3UKy03/yQvxvCyXszucRNAN2HQWnWPr4NwaFjHUP75
JKHj10JZqFbWqF6TNMBtpHcd27iyzLkN+DWQwiHnEN9OcPKps8Ep5mqZ+MpTV7m5
5ZvhA2J5pL2ob+6zpWaXcGJWI9zRlkzgJFxH9Y+Ye8g0Igke1LIZ6qvPtRi/4Yr6
/MQNLGGT5nAIIQgTRkWWQWZWJNtluYmMH3XQzanWvC2LUUG/UNHixfhS26vU/ICi
0ef71Z0+BkpUp5Eb4Izo8Tzhc4wURkh0SUK1ZyZxe6cYUzc2E3+0BZlkmwuWlrny
NV1K233505wwH/rotsuDAjOxxPIOIxLK3NWQAbheser9mQ+ABFpl+BpNXvIzoaPo
6Cfys49KJD/OLaFFovkNrgMGHrARoLRg2T3QQwQy8Wt50g84ZATBB1xna3mZPCv7
Lz7EMhqyEnZso48gkDIJbfprAqnWyx/jKrs0G9/ztFw64UCJDDObKT7X5I5wyxrH
VY7eH1VxMBPp6aZ7raUOC/xOmwewkXx8JJQFc32CqC6cnImCac/236z9uDfiH0op
A8R2r1DEhuyC+ynSG9AHf3gLYYgDbel1IMmKWHfQsXUyWrmX23QDDVhF+2rkavSL
8YMgC27Q6G5Yr+H2GcVb7ITTmso51+AfQAoL3kyNTcy7bqhfimkyYF6hxDENS4lW
BK07K+mRbkIJVz2SNbR6GJSJtLUJqhcLFsvhqPM+1dLJ/8r/d8gCoUzS6mpMv7tE
J2XFLwa57+faMjkZebmvHbY2MzJsqOj1T4IOdYMPYJ5q6ILGK8udtbkpIJmg4hfa
L6V80YiR77wkLA24GuerBbf9ljQjzCqjIcnbXcId3Il/Zqc6iqrbGlpoKorm3NLW
J2w+Fj8Mu8piihCeBY7OcUHlBn93hFKFP/MuJrp+P7xlUj7+bW9AB+uZ/8srjS6k
2LQnmyVOfybzOFZEzH8VWc4C8Pf/DrsgMszT6EXLWF2hIbvqlDJcNdCTwpT5KrLZ
EHeaaM35kLetr+6+R/MTZE/hH5EahHfWya3gv8zuPjnEZIYg5TmUAvzRe1/U7pRD
ZfXI8YFq2ob6fmzjLvZVxsQKaJnSY136mzTCwU5TqNabDwASfeinR6qDb7tgHAv+
nOyYQXG3KhJ5ex7kSNjtK0g5lySd4UUGkE2auyiNqKjaFqc44E16hqE9ZBPphOQ6
j93ccOrEoXcE6Emws6iWWQHjKkIPDcXzziK7exyc2BIZ8YttYqrV3I97oEP3vfrR
KIzVUnYkWADvK7oXgEprqihz/X26gTxqA1m0lZ6PTQp9spWuHtfdNHzILRbE5dcs
eazQdsZa/FT0NiVCl8aK/dZt7F3NZHbqz2s7DIbAw8xJ047LzBJV3E6UzP6PuA27
/N6Jk1qSVQSZ4S0NsG0Hz9SzlKuw/uTmzl4WUSBIcdWbB5m42cKIe5YI0KSgZ+1H
pPKKtTWFlQ/h4QJ+dL8CH/gmG34KbEek3drC5ijOjV6ar9icR+MEq+IJSt2JIVJQ
GkUx2Emc15xlXLR4lN+GZiuNRlpqDW17JWoBhUL1GpCpEgXWAJ+XSyKWhLlmmwEz
TvTSkeZCiRhIArAiNwumTjfBFYTzRNhSVSP0locuz4VdKbOu100PQmVWFhsVE38x
fAVIx6/SYQxuw0LOuzctflfVTiA8BIM2ZaieNkc6QftlodgDwVJvPXA3Asav4Uul
qyVbxB2hcc8L50Dc8uOprlONBW9KlobBspYI15YJr9GUzpMOj4TndX7VnxhysE+4
i3/bffjtSajAZbCeC+8d8v+/YxQ0wsPy9mZYRRWeNj3xuAGK7ID9ea83UVWhVbT7
gyWoRyYmYDyEdELwrov6+3ner8dt8UI8IuiF1RQiLIos0zbw24MrUFUAWqKo/rHu
KD0FSEMqOgRkmRoxVo90bAYjBcxCp2AKD9ufypyiOUJI3wd+QRNqMC1OaD37Ngwh
hvN4zwdEibqsp+OCOs8h7HrwdjbGhAak4iHcaq0LfWgIvjH+I6xAIA3ndSDnRbh8
LD9D+frpz7NkVXUkRWFPg04LBIseWBCjImSRN1uwlbZ9t3V0TVt9ZrrpHHSO1EM9
6mVOJmdcW3oDKZcXnLw4KINnNAsXfLu9r3CfbLX3f58/f7vh5ot/P8vz5c4GMUu7
XUEICXg61iXZvvbu5pJSi6obiQ+b1cYtE39rDTzcu7w3YhCBkI1gMp0buGaYVrCz
E9Ntt/s5teFLO1ztUht5OW4GTUQJTMqfc3/HdaKHDtIOP2utZ18FDnbomXS3867F
RVUYsfbr4TISleug+0CZfY+OOWYaRdrlt6iEJJSzYmMlshZD7+5uRm9sOv5b0JKw
HG80rI9CSUqKR5dPz24GZhBHZBLdYQED0jWRdsmuOXJOjlAs5X7ba7ErPGzxYXXq
nGW7S/0qzj5KSZ3/QF8m862/B59VjYQuKocymPr8eVXQtxCC5h8vIj8woB56Ny/b
ZcMGtAQlzTujXaKVmS4r0Sl2FMyhuHUO+rw+UvVvOJcZRAqCki79tKZPz2XDKG+l
oapddj0Ldf6T3c8w6J429lG82lgcPNSHgJYPWKmG05qQNcue8HHBHSTE0twF3AmV
FSOIXzXLIphaHGD12hi6W81WP7zetLIHIo/S7APjMWYUvaFq5O3qpa45HbPGapgx
sTJDV+LaUJEdqH1jMw54pEAv71Ae1+DVCruLCDqU3UCVihx4G/YdPu3mYC3YukEZ
uAPi6kGQ9fj4ztv3cuz+G62ds/8ee7d/A5xdKHzjCpKmNbVvjq006k5JaGyelfca
E/kVJdRPYo6EVBxjodXOnndzhad+Q8QDTeP+FNDwMlm5HHsPZHfBJ0Py8qV4BPNo
O8yiivWT7AAN++gSWByD6mhgEY6igrB1vE+FaI9XmXrC6doCSHUIl0MdJ23XIKIK
q7ES+oKn50M/wR8cyAAr3ixDBj5CN0jm2Pe8sEISbPXMX9wzp/wMtIVzQK4DJc3a
FJf/HOVLeUeYOxepOuxAr9AWbxzCBp0m2zAsaxvGnx6dB4zBNfccdMyCgqDTeDoE
SmB9VEsAd7upMqxGQgN2i9Kl62MRehcreQ9LI+gkE/kjFjoLPBMN2TDI92pPdBO4
7DuH5wttuwzf9phwkGHDCDI5fWOO7ul0QOL6geGnj3brtFqPaxqKgPWUjQ+c+PP3
zVCpVHk0WAxJFfjvjJrqkhu1+KLkutuHQVS8p+6dTZYq5U0SK4s7cAvCvaeFsbyx
zUSoO9G5saXqrO3ydWKFiqXF6kl35B7/vwFV6bG5jUHmWCNPH2w2otd+VBkl0htB
XV8o4mx8GHEU9rz1nY6xBiYaIliubBBAM044xequPCvMZ7wm1NUQlBPVK6A96kxe
7/J4FQeyfuNAqu9nFRP3Ycwio/j4TlX29jRc+pjz5NAus9OqGjenqNlb8G3B6EXn
kc7HKG8PwJCL7nFWdaypU7m6f7APumco6YowoK961H6AfyFSocMVBkNr1uy8zhdv
Uyzy91xEyb9mdPQAfk1uKp2G/Bg0arQTPJjxENoBgBBMAsdS/ax+djAH2TRlfCLV
VeCZoi6RBzH9UPQHLY8Z+8ZSzoDJk1t9JIzfBuDVpmqzHzqnxZ7J59pTOnW8uBYt
DkOlC3PPtQa2JoJkwSeKTi0Lb9kMQ+e5QjU81e0X5vJBQtqGvzWF3qfq7fwk1miX
T1/EiVtP37AXCHSqzkxBXWoRFYF6FSFVli1gPXq4jdsbjJ2k3MGWgwop7dRj9R0y
rXiF1bjOLXXbiu0UnyhJ5MssRvFWffAXG/k6ThHv50kB4sL5KWXVfgc+njJKej//
k9yyipAd0ZpdscF5/HKPDuT3/FxxdLYYuRtzxVyd/CdWPsZwOj4gnC0b459yr6JM
xUX4JtkUSWGh9lqUD4ayR4ZIDNbqMVn6MdnXu2w1Dlkp87Ugl96sWrUYEgpy8qZm
oKfoWey25OxgLGKyRofD1Um9s3GvePslBHxsUPd7Om4gcZuJgrMVOwdek4Aje93C
ulbUwlOX3ZG6NBwqo6Jkz1WWYTxIOFkj5+Xqand61RqtrsvRdTqsWeT1XcM2FzcN
wlICE+RIL+hL2DoCsk8OF10vgyPzQSqew6Y5vnPOy5mTxbo2ymZjymFuCbhyDvSh
TVzBm1algCGouDreyI6d2AlsU+pEAvMXPVfN5hBbiarBjmyWm2396UnLpgzqe6Im
h/sxUlXX+PQCIaNkFX6y1sHzlSU4yzDmJGHZ8kEi4Ml1psuZO141rcgr8wZp7fZn
LTQ+yx6nOYax882bwRQ3RiJ98FaPVw4JzF6tsDR1Q1LergroVMuGLR4rZuDBPZGm
ZxK2ADP+lyHCPqYJdzGbTk85f/b0k58RIf0jf+ChEWArEor1jIuWDul1dgltNbZq
GM3QXFWtbGmKcOEgqhUwIVCCAHx5tEYJlq8ySvPOUAJN7qYPI7IVhxu9T+MEGnXp
PYyutoreHz08AdxM9yCIv4J9CWhXPCqasJMb65baawZDnMvw+NlRz5VGANTmNAHC
EKtll3goHtORmanptGTTJv/P7w+4VuZH9/CDz9Vecb2dYiRJ8c/kvleYHSJz8QSP
1Aa2HN+JXhL/DgCCs0HPLNUBqou4H4zHqIaWf6zHGbbWr1vYyZ99EEzwbaCvLPtR
7/iKmEwn9CvKOvjvzyx+gdHcpC3qKnINPdXYiAiO6vm4nFJim4tf1RMpZK48Jdz+
+eOznzMvrmN3dv7Yreggh6ck9z/Q1E3fe9yCztq124sx88DxQP0ZPJ9DtgA9oI/N
gu3oc+DZrlmjWahM4Izlo4x+VxrJIJvkp+Qqp+YmtlxnmeipDlQNRTVUWzP/NhXv
6qvIJ90DS9dg6IdXJaQbF8w0uJnNHpseYH92bfKLYgfrxHBhGG4f6oRFhfuXtGmN
tEzN8A/dDRcZKKqvsJYE+n78f34eAqyVUtgUXegvhdKXXVUO0s41yR6jyZAGWx2q
udu2akbX1APgLzAznFxn98/46Ny1u0G7HWwTMccGqAsqGj8kilkRCpcD08GS8ocs
Pz2bLX2bppJxCOwYt1XrdP6WqNqwS9yj3hbN21ZHdrYYyGVx9sH/VywW/gHLCks5
KSM2ux8nuzlsjRQw9j6D7STKCKi/vf5bKRecV5HLpPKF6FJKUwsQRR3N7bofRFod
jDdD7Tn/OOhhPcVnoe/asmYa0BaLbdMSEoG5G/jQFQZBTvL+ktGAv4pJ6lvqXNv2
1yzo0emZCArbi8A9v0C+1t1+OvrCo9dJV7P07enj1zGxTCL/kaXzxgu7LH5eJ6FI
AVU0fTsYjfHwhhrkQwZhVSfH0PRHCnBtBqeSb8XGpd/11BaqjVS99JMdxqj5AeBi
E7WZalYUJAXvMT121SgEyK+oGqohxXN3rO4w+ex0cz5xOK9Now4ChhhxQzJzdEty
QaRPOwDn9XefeD5xuOUT0XejeKI3l+N+fHzuyen43wtkXhHrMb9bIxku213xt3dC
Df2kKY2cOJ7TTXVOB01u0fHiba7IFHYVgjS1TN+FKr5nKylaxs5TM2YObn9/RsAU
JAFz2And8XQ3ZyhUkIBJc7YlwIrK8rtreRZhSwhnZohlua9tdA06f06Z9SHsFHtG
DL37ufdYGgTDknIybLVy1m26ey5ErkuEmsD7TnganVDbOxL7ZMnMw3zCNHTXXgoB
UV2Er9/wPdLEpvc1/lDhU3+r36ztsfrbkEbXu72mgYDTpzaPfGwJqaUyaQ5diRAa
ENrBqYUSQ0CMxeOgeti8MblcCv/IzwtBIhaw5GAUHAZ4qh6+eILpubPyzAL2ZEfm
1j7m2HtjFaxLDPwcZA59sL0qYjdpPabjsFoIu4YYoCstonBpQiv+oZVadI3g6f28
C6FUpzA176FlavfBeaC0o7If25E6pFToE40raPEn1iSqGiTxRpkBN87FWTlElILS
Nhy2AE9SArTGXomUd+x6DiRL4PgARaLKKqoHOlAyI1UAjLm0SCDxp96FO45pTs3O
4gWdxGpoYCpKfQxTaeGRo9m6M42XxI0gpBA9soHiJC6NzQptYynrqVPPAjI4Sj1l
/NqDl2Iw74BtrXR3r+9QXxjNANt9Qmdvf9Uj4p80axdLfuxlQwPb3uuN7xtGmY/+
HJTqYbyg8dgsYdJUXFlp81kw9lxgVrwb/zEypSHnbqoZMtBVGvU+cccjZ1GSlUbW
/rpppitoyzlR1NptZCe3d2XXfl4RiJoGuSYK9LLIxwe3z57yPoKJoFd7QhroMH3d
ng1ZXGGmcMT2mfrpyJp70Uaz0iKfS4ZLMO3/ywKZr+JFF6pfvom8GstV7n+8otkt
H7BBsWCK/GedBDLBKthCKec4HgSkDhy9bn5Hy2AK867iCCMFdVE9Y8MkK8CZhi2p
x5FKb+PQr6oaK6CXbJdOi/Z5Y1pCwqU3+bvUNBthXaTmgydwzyVg9iZkP7oTadCj
ObK1DKDy2tA3tz8hwcmbD/dWGDcGmJ8pu4AMa4XXwTY63pBbU5+5ZTMQNxDxbSKP
W/+sswtn3dVTnezyxqraN7Zqj9SJiOa7/LY+o8A5vpcxvR/p/XVuhPdqnR1M9PRQ
Cf2Anu3hRaNDpWUjJtCEMpiO0/mkzXYxVAQj4rXbwQL1mwGTzrCYi1qajECMTST4
yVXFSCIFjMK3ZorpUmww1twnDPoYmwVTyMkJLdKwyramylLdebmkB/Jej1UwQRjN
B6aKL3bu4SX3kSTd+pcFVk2pKyMdzAJL9+qk1lOp7fj3InN0o0W94jhki/WnWACe
gOTLxHHciYVXSLuaIjl5LbqyLQSRBHiZxI/QU8B/vat38pnl3mjuv+xJuz25SR7n
N5RO1TGxSs/IxR1RwHCbSuckCKR7BL00yA7cUGni98MiG5TlgOiiWN8+irKEwHAb
dSoB/kdYAaPk9HRkMQgn7Cq2gBQM7lCpiSYvS0jjC6dn4pjGG4+fNzLf7Kyi6TG2
WUNpuM58uKR5xXHhIcCGkpSEXQJxVSn2K4Xxc5ktUFRc8TKDq95T2cdAxWL75uLE
zIwWEmQ/aNI9dWe9KblhYRXg/iPv723zUON7sH5NdKTwcltQo1Q0KBZPWeYYIoUz
7X/Ds/4Sig4Q919AJqOu/6NXKEshPnJ/MsW0WB7fEdPfFhgM5i+uFWcuLF10VLaP
WPosd6u3URI0pT5iN8aeVMgwNZp32ReGjL7HaE5NPxQU4xV1lO4nPtXwELeoX/44
P3TTQfMD5HHhFQkhTbi1O4HqANsrvFiFl+2eiyS2jQseAmrnMI8Owr9LTCF6iJnG
BPp+liJeB8P3GvjGIaS5JJpgOldow/qdluk5RvoEqXug26N3kz8me9vSDpG4cMQh
/iuph1mtH4njw3ByE5AXPQWEyeLE+UzS6dtYHCA6+ZFUVYFkV174IkyPPe4s6GWh
V2Bre7AXGqcxEyBaDltqbf14OB45tap5t01YPWa2HqIt+uf1rR33DMdYwn79zBjK
QfAEikBaWJAD+9tI6CDOcsYcI87EXd3evrGqH8LbmkxuXLpAFgottxEgvuac78nN
Aac1iWtgiwCKubQS+//QCbTuZ5rIgIFUl3o4bH3aIcl3LQ8fkNc31GsHSUkcVci4
76zouyi2CvJOnx5A3i7cogROTEFxoPkbaLZfBj5BXPLvwSNXNkaUbjTq5h7OXcV+
/F6FNOJoW2JUrz5CQKJ6S2G5KKVT19iGVO3uPHtyUpjXdrhvlbNeH6nZ7wRSmeei
G2tJ3BnWxIfFKOt6qPZLuIxrv4NNdUzo/s0R1vxG11nWuLbdl8mAb7RTBB7fVCzL
noV+3K4SGEgjBWDkHmzPAF41GcI07w59rGde259lQKOjVidU+3ENDQHVMjtueCRz
1we9gM7iZH1p+6bScvZ1x1IySdCyaUosjEG5MQku5gMXXK29cZm+INAqrj/CKJ/o
oFgXQ1C1zRfsLzpfmO555uyMfisXDucir5IKWVH+bJuUSK99gHDem3Iz++Sk+mT5
q3IivVvMplGWw7yyg2P7l0C85CrbdMGpjl3ljRz8eD5ZMlZWRD0S/B23Dzv9KR1d
3YDe2g7+5UkKSIqxqAgUX8mnbaN6b57nKBCM4Rg185itqE33fAeGepER9V0lCm5g
EbhKWiaTqIlWaRqM40RWdoEfVHWnPFU2/bavZZOT2u0OVZlaCrrCu8oav1bWYolT
iYP8BTzv+tmwi4oqLzRjtPFX0PepmvDlDR8lhKSYY9NxlZWeluyMOm65gNHEdiA5
HYLQw5MHrcyIQSu845qvoOVM7h9Swz6SZ0HPHTJsQkz5VEjyuFydUv85uM6kHZSl
PH4PpNKU8jmYqHcRBorLXZijNCXPMddfq5qI5p8c0+Y0QL1q+3AuowkHugV9toPL
Pxv1bNQNYFy/Wd0qUIfP0VWvtVsJMTcwcYe/LR39+ZgATS521kHVyFGMNDC5fpp9
qccn47aZ8OvuDX0moxBj/NJ1NJR1B5Reip9Tan6kRqYFK3Z9twWSN4GJlUV8LY+Q
Pss0J3k54FaRu1YJ0FsYbiJsv5RzLy+c1v3VsX/5I61WKFNAaljPm4uQSn6GFeDK
cAQI/8OrU1QtyWvxH8GpskR5ogClHFMf5xCqtTQgOAQF5gth2560Mw6UM6OBTgEa
o413+pWHdBEp74KQzXy/d/vuuKsupDWCHVd0mep/ftlDpUBr9TJkF/xFMBcCJWSF
oYJOYx7Q9ktILPZaHFEA3tMObbJASo/hmCd6A5zxQ9WP+PyAYL0nuk9ZmwCIZwQa
tMAbMF8XX229NxaOK8VP17eJN8rvD+mMjoL7UEWNxO0uTJcGltS2xT9weebQb2G9
XzjlPhKzd2BQl/zSpxQJzxQHNKsMSG5pKQjbDWH71cF2g5YCKkogK0hat5k1feoK
9rOP8ip/TKHYueB2ijriMgTjG4IQti9ipJH+vvUApbzmZEzcyjGA/EcW0sQELpkU
hYorGKR4Om5rH/NT1jazs7/yPkoPCo0IsfNUkKqV8xBaLB/RB47O/73WqwihytkV
FR7Gbs+ayt2j5VR9CuK8kS/hRQs1HsG6x8wloQd4e+qe8E/BrAASN77qWMPKo14m
bjI+wRF3Eq0YhXNJ7y1NhKZ6B6RMnOrA/k39F1ZVc0DPfnTj72BIHTBfMiv+3ZEK
PEHaIhopJhlWab8Dek1LXU6EXzALJMPLSGDqmWwJ1uc4S/4xBbd5qqOQJsVi0c4c
7BNOT4oDawWaGB7JkHLfxoGFA3Psl0m/Xu/6dGuxXehjkeu/b1fZ5JcFD/Dhn0bM
lGDu9K4l3WTG76612nuqf5otQuknbYtEUeYpDPtr8y/QGVumOJokmFYJWfPba2CM
+Omqz6bTZeN4PGD9C2DjJ8CvCQGDl24vY0cCzwz32zt8MzK5F12Ugv+W7OuGwAMv
YcnMcSXYuMx1Un3W4mgSp/vunP3wwbUGJY5bTLQqoUR7Yt1GCHS8iQXgRPtnVVSk
kbQcyk5r/nEtJY5kPLlWAXplqTvxeEvuKMi4vumZ9wKnpNY14qYCEf170srOUkv6
VDtnW7ihD7w6KPg0yse4iVX4N5tiJOvLgaN3T9bp/pO/Bl5bDtRhIT/Tov1RJtDb
YiSJgJPhndOn+GungBumX2H7131DnR766eYxdygFV7IwKiU0edSUgxZkS7XyTl32
mngJ8fEvPz+OY5a1qBlNC9HhHBTW/tO+uHGm1pfrld9T3iXIfXlWHKXBG2BScmzx
IRouRgp9AsFa3AK2aXjhQ4tBl5DJ95tw90DbykK4D3caWXeD4xBy6C9hfwUA9doC
6KjazMIzwi8wRoE7UJ0dYSDgSqeIVFm8RyFmqqX/14cp52NQ+Wop2A7JoCJoDt+L
HXIDw+XFw2MK3Nsfqyb4wAoLE1Y1HpqI0BQ3d3wYhxBLxgXNKoPUjyqx3ps50/NT
A06fLqVhRmvk9IxMqp9M9F5S6FYI2C8eA7RcrnajKtFRjw+OfFAR76yrt6CfCoC2
rRW6N4SSAhlKa/X7ByZVX6Bdz9LUStirnkp9qfTymyPqPnr1LtLzba+GSAEC3054
GliMbJ/Acm1RRcHGn7x1W3E9eMeL+QaNGTkzjAH+Fot7euGgJb7KHajZZu3jZYFf
3jRy7gXFkKYqK1KJxxtBQdvN3QmLT4i78PFVbEApy1OYUG0X1AdoZFHnJnLgm+TU
2KAOZEy/q/v7v04EWPJwQLVGfCXBsXn7pkG4SpdakoaFUajOCkxa2dmVjj0Y9I8H
o5uQdgs4+num+85CPmtyAPnPlZis9YTRW64BEkLPw9I/IfHFI0bGwDgFQBdowZ0y
XHU+b2jaKUFwo6mD9fvPP2V43Fr3/GP89S4wh0PnY8WVZtfzLpvSAt5z2NwA4dQm
Cd9t4XUhd58C6KqDqa6yJkg1bh2UXW2KV9NrgK+WN70ugy6XcSmLUevcCHa5oBYv
VTNStQlGRjjgUrn1hvGI4Xci1nzeteBgz3fT/uBlpt06bHdFwxPPldsKf5vhk0H3
zfYjCytjRxxQ8zixuKFe8rzEhfUdFImvGrqkhaxHKFDVTKElWgLNMUceIBb5xniB
v9NPACNikASqaAiox+XAnnDP9I3BW6uk54pGSG6gGxlONISfrdrdMW/dQiSuDpbS
pYJI1VsyFpl9+qHCZe7jFVjRnLGyeEbPx9QOGxGTBKXvbFP5bTQOZxSveymtADgw
yB6khye8EeeOTfYM9po5R6Wd+F3gFExhinh7nrlUKCSY6FcCe3WCxCmmzEizIvkI
Z9QhfRtAzR1aNWrfJGP7HIU1LR+Q7X/8yxkLOU3VMy6fWu+Roivswn/jALdheIUK
J5o3RKF7Jv1Usmw3UAaIXoD8UPOfxJ3TMu/aje5/d68quWIDmYJBIdarVx+Bp/o4
XK3M6OquHa1pfoMGDYq2N6BOSx6yWUHTgTE7x5VXDjqNMzrOEKbZz4HMGZqHg4ki
0EJdyZjOvKYyTz85B4XouO3FCRmoAn6qFSsGVhWm0VNgcecmqyiVgGZlhwFXtuOH
V6T9dBf59kvdFd4A6CcFW81Fy4pS/fhBIU/j5xujcf/sY0ScqtR02OLldTJsckXC
iCpaly5B8LkZI4SPen0xCgkI+eqmdfpCQGOmMMt6drTFtuuzl3U+IM8ilBXWSh9I
viqsnkdi+wMv1MfPt++pQRMr3rlIDQgdtMbBMJ9luE7BSfT3LO/qEMUP4aTPbTXW
Dq/JEVepBD6P91q15bonNwnCLPH/e0ukcRYji5/uKiWAU2z29ufNCpZ9+8a2WsPG
ONHUo/LZWQK6wkaSKo2BvCRIiGlpKX6BziqDc4qzifHjSqUsSyFKZbnHXUsauh+b
TU8leaKgj9uGZZ9QWjmjnjCrj6MlTb5QwYyF9T1qZ0weSwr7uaA2lzJUSrvx7OE1
FXio+oOpfS2aWrh8YBxTCuxffp6S5NssGqiG8QAxFusvCATZobREUkj4VkaEWRYo
EBW2IzIMR+IfcmhuRZwbuAPj+Nhvn0pKJxyuA808iXhx3uw22ZOgWcdf7wBwPwrV
PdkKzXoPjIJvsXKv0a1vL7fgZuafjtvuxIpHc839zB5oIhnAxoCNOuG8zVvzzR9S
fpg+ses7ux8uetxhZ5SyQ4Ls1LIB+/hP0YwTF/9lMU/uL19OmSlQlvl6L5LUEEQF
ohbfTXykEp4aL7vm+QJKPhfUzWmTmr+GK7oVUyDjssCztKat+zYZ62hjdRWp0OdI
z15z+dmH1YfO0+97N5EoN+YugsYO/zu5CpFpQZZFKE4t0IkV4z1NFDTVrGN0/NOL
KEQOHGt+G0MFvx8gU6gfV4foIiu75Rz1Y2oJRKrh9ykX37q/eB5RmXq4Ct3xibfd
EUVC82V5/3qeJCBsMBM8K55AvF1TPssgkfbwfZvQwIqtpeOZgOiI3I1fmW/f+6tl
yxdSgwzKVWmZSPX/tNB9sz9bexM8RiYGQBmX4vdu++9ImLV7i7b2omEoGq+qCe0B
IBDwnSE5jAG9bHkdab7n0EZpRElUKAGNaBaRc0hDH4daq9ugY78zoxi4qx65zYH6
wSh0wgBo0xydOe0hiereGzKcQLDAiA0O0nxFLMmMJjXmzIV8p2bA1x5DJ9SsVmFW
JFdUR8z5eQBhnioD9CJ3IIOV1S+nu9alkvZG56HOIYOgJ4w6gLf6zbNWXoqoPS4H
MFR/4N5GQGzwjK6kC8fE5AsznwaGDeFQ07gGOulqs4QMiTiijONL2ftu55xjRWsS
okLV/8eEFrVE2gSz76LxeOFh4pNIvBVdOpXuEOPJrqy2tmx8GhouVDvwDFtmw0+T
ihTRi7JRYemS/zJrOeDIVPZysxRXVhved8JaTJiIL2A0cg8AbIfNV34cdpE3wk17
cvexgi80GvvUbtHv2bBzsXBcUXsnZrkuAKokk4C/p/fDkQSNIwVSZVrvqcLOxqe+
oEyzMK9v+kd2HAQgfWXp/BHwVeCLDzf7P1Zjr4bY2AlZX0keCaWiLaSZZG/vFodj
Zn+7u6kcx5olwTRdIWp/QSlW5ZZePB6YyXfzcC5KKE8prDkj7mX8mPLf8r4HtLlr
DMsISiFy1r4RAOMvSWM2vipODSrbXyOv2g58bjxQrTavkKIfA4dwXOPfkYyUcTP2
tH0Z7iHctGtyX1nf8kWeFNLUAlcSkeYuj2Z8dbfbIf+wRbNJT/2cEuzBk48/Pvuu
LdOdvT4QT4F5eQf/xMDcwhK9OhrTjlWfKhUxgtfTG3naRRyELBxomZUzvb0bwtgd
dBxbq/hlNonB5ew20mcdOFOdJE2l8qqiYw9jDx35kteDxEkwy5VtPtZZsyrrsbDT
gMqnxLuZoWnsfFd/J7JRpQ/xwMEItO9CrElZjUnibPU6fKJNvdB/wf5UPlooeGaN
vrJyI8VtdHFJn5Ka/1n1aZmE+qS9q5+CeDtAtm7ODgf+dreLTKxpJbc0JnzbJEqD
hOOXP03akvSP4YCWBEoxwgyrz3Qg0p6JJ9KVA6Dl9iMyIyJHoJWsgKYPR+shyyFJ
5z9R+oHXo/Whs2lXVgkZFlMJreUVeWe7hA6E+bbZqes2U4ZgVVeTBdLAli0ENX1Z
1b0jpBQ9VIP2YIau2bWCxa69TsRjeJIsbIObnhSRP+dJ08FbbXsst+XV2M+3/XH8
J+c5e4vzWw+LG+DSRA9ATW+UknhkmzZbnHSV74giNX9qqG/Xq+f27/wV0aemCGnb
RiSL8hBMsR6hwBhLwIvXkukwXzdrYkWE2bXDxy30GbdFTTYTLWXwx/8GWxzvQyct
LI9eP/ORKcDjO1G5+A4PE0KJjIye9MMLKXd1Ki8QmSlhcog4DjCBziXjv1Pscs1K
KN4UrtrXG8YlEQwFULCoN2l4Du4wMtPp3i5MtjiHUwoRSIjFYOXlRxK2MaEnNLvk
Bq2aD4GrHy64D+F6Wu2W18Sd+6K6r7D8tGkK6tlVBojXtKcRj2BoFEl01B5iXE6N
j8XzRk7e5u2kELQUfmY2IFBKWbpJkZ8XYzun/aUzYL3nzI9YVEkta6Pu1KF4x5jE
dIJF6rgoABTHqZrE6uDBJw38KqWGRbhUKcBpX9i6u1WGROgDyv+zoO8J3w4CDxnq
xvgsYoIKKiU4U7YypurcgVam6YBBj7vWHBfMI6qxotxOR7ZCsZ/36xKU7THizBGL
ZSsFsywi0Bu7DoFX1A9gd0iZLdFiuiHO7OLIOPuCPyOEXcm9YAuLBx6tVTUoK1jx
xDga4HcBA94RcQzoSNvPymLRteCkmgKZHxfiPPbvtRu7O529AhRoCXQmZxzh0KBV
MgEu9wNLf/+3vSVH6YgUFe8jIie4yW4sQQh4PWQtex0/qbVmHY8uZXKdmZxZ1E5i
pjWK05/FSBmTwK7KEJXeTxke5uP/CY2PsdGDjoMk9R2DzRZPruwn4X6yhdYxCHZu
hqkh0r8EwcYxgP0x7J709gWMCBou7R+oyHMowaXb7PoE0qKBPsV7TCjrZZCHA5sx
G6mMIYaDz+FouCfE7LZrtNrWN/Gnp8Jj1OxdlnU2QqdaT5kstYBBscJxIyHC5Doa
+BIk3HByhdU8CY12BZTTv44lUxKRfaGlABVz1nRKCAnD3QArcPy9kx/f248mzTme
FY//vgQVo3A1kroIQGiRwHIKZHt5srle0jxnCAJjWG4S+xvYH2SIcjsteFlTooU9
CYHa/ApOJN5qpe+eXPP8tA2JYM3/9izUklMsf7ERuLv0vcUr1aTCsKT/DaaczC9L
ZA+CfvIltQUBcxT+QN6GwSOQTRSuR13VrE2CFdbanHT2/km9r1zzz3YOTkwDYnwX
tdNbO4ISCX1xI9lbgMV8XHn+f/dhugSX2avsUp6Lo9WQClzG/WMV+a/8PdQLUEu+
0x0gli/btvoHlCN7Ep8xjysmFJzSQ7lDMZ2RE9jF5721CrLUHC9ufwNblhi5FRjQ
fx8ftJYuqLC95uKckv1VPspplGZmwZlxQoMgFhayWy6oxIfDbjSB0hFuXCU2MN5g
bkRqEpk3Q24sTA9/hro1WXG9K9Nak9S/brlRHpKX5yeHh58NX2cCaNFn2PzVLR22
gkK7GmgwXSpmd5lBocx349q8hbL8y3FeSfD576XKpwruro9fu+U46xHOBHwwdEYU
r984g2M5v0Q84+SMS3yoGkuE8xf7SpLhVd2psga9KHv0wNH7h498AKfeZqhiI5GZ
mLoSBPOXwIsvhUATNbuTxDMjTCG/rbdMP0hhhdgayT86kEmsP/Vzj/PJymN+nO+2
L1KfYvFDWxgfTRzLAnMUhjR6cixas600sr7wDOQ1uNwN5xaqwJe44NKkrWFkOGqN
Y3gC3FAO/XTMGZlJzn7OmwV05RwugI4IWRFtB7HtJy1jPy1Pc57NGn7D9pmrnPe0
0koacfOp4RW0LeAR3IQr0u25Pcg1+IFar2U51aSVbzb3j0yvVzYXlIooulPhigp0
98W0SgB+Yc5O0vRCg3V38km/RNpWNjnwaAs5RqxzaaHWo05o6zeLgf4C2baLIsJX
36/P+5o6vXc3+f73rHhDNLQnUQNwqKSl1wMpAE6MDKiDdLXBJeO6z2zpuOU6JUsT
oMuUtxqv7aDTPDTciiUswoKtvLc9fHmOFp6+Cm3A5A91Yd+M0HWliifBdQ+svymY
9UCN1lBcfmeMm7GqV1hg5VCrjqMMOT7IH2ltx6VWU2hPulqrIh1WF0UJ63PfevWu
YdSStJ3+uHbClPCYAMTmjwe9u4szf3LSMAbXzAcHGbm1RLfeqBWW0uhSUqskq3YC
6fLpPW9bsETL1P+gW8sGyc8hkPOm0O6t+MSLYbYfF12ELGUYXgaU0NLrqjGjdgPc
KE2/nqoro2VNHGhf0xqV2gGn2TJkuzR3sWFWuOXUL8jMptKHW3xXHE31xdYLJ3zZ
ZoDt2ZrRJUHLRMzD1UB2WH0C0Dn+wPN4rzw/h72hnXaWK+wutC58SKndaed9ZtJb
t8srUpK34XksKdH/LPpe23QiX7AwLT6xvErliQmXdoACxFpO8463EoYWsgAIbZv/
Fuy/lC9Dw7EVlmNozj4zlPQYSuQdMqvf3rQmb+QbAIgtXWgXBA5Y8Ik5rACGEwH2
mGVAktoYDBMiAX+dbD/Su0WKDRT59fZcwg+YhJ+zQewFv3vqT8WVXQ7evKNX35KM
pOk4wu3BtLdL/11Li2LA4OJEyNmVuox32QgeSCO7GSFERO5SujGYAx8dS14DfE7n
bxYbpRGRF2VbH9Y+2G75s18VhwxtRdbxZBMI4P5Rl0j9EeRyRfZ2ATP7QfF2v75B
XWm5zzAeb7fWfpSt3Zp9YKHnxnJNUWCveJAvC0ugKNCoznbuUsWiVoioHUgb3wKV
dj0+237b5jPEQyNeJiJdRI5ZJVbJrdociprxTs1XN5CnIURCkimTGQoVWggGd4P7
DFgzBXSWJwktsYAG6o20DVnNaeGEpulKV73MRPdvd/S4EUMbinT2Tlwk1LakIT0p
xdYIlNb2uQhxzjcCj5RALuRv8dZ8/8K4ysjPLetbJU3HQ6iE0MQysiHDOhUQ8ESd
g/QqS1OhpGAxDcaK5aZN86zYP63jVL+JeOsmQhCHXqbrJ9cD8h8vlScbUpIZoyl9
8+lTJIw/AwE9ll/dIn5bZrC7UqfK/kXP1x28y3K8L1ZUaEfn+4Dw6ajgtQeG583N
fwdmssIRLFI7rpZxpcP4DMHsEyGSsuTBjCqgIuSVrmIgiGCvBBR7u0C5vzlhbKbw
vikKD6Q0HqqXhdGU55On/rpDfHKtfwZTou0CI+MRpAL5ZoZ0IWVivGfDma5zUAZu
+Cvqc/oMzqSSWPCa8RMt7gzUfkMWHqSOu1VSDHrFs81v8ZK9lZXFEvsPG5ovcHkt
0fWgHv089780v/A2u+R6Ed0Yv8htO2EdS/LyEplc9QIHkpJzHOOyR2UPN01MJdeQ
C5VsOec9cVMUZ8LRGDm9lV01bjxZDXGlM51gAuKwi26xh8wI+3eFsLNNRj+hguRI
XCTUBF9vqatjPA1rZBsZ95Mze04uZjDFeTwvy4fYv0LaucVYNCJNu7mNhfjDsPZs
OaUOlSurHJZfl5qR1+HTE6rVqQrgtLB3t/MqSNmZq8QojL8mn5YfKEHJSRxBfZ99
pyBqjSZlzSJZC3NEiZ30mdvVJqRyfHMmys8iQ5qeLwTj9El8lK9CCLPwZyZEvg7s
6z9Lxy5AOAvT+Zsi8uaU7K0d69n8gvU0yAHarQ/VQntiG0ERLYXzBxpIi+wawXiO
qCq33vqRLZ7m6meBpm9KJ0oP439dGl7Eg45EBmZPOjp6RU+RW99I2Uvj82GLZe1K
oOaNY83SkZh4gFJinJWNIhoWK10jIudVqv1pmFiub6CEbXxuAIxpYHPguuLApIFC
zMg7e3m4jnekn64rjI7mt96VlX1M6MiVC4o3I9wlDZYNR2AFTegApJHlwZX1Sx11
eIPxyD9EEB0Esw0wUDdH9GwZPYTD82C900CJk2DKCjRXTUS9K6HkiBeLH7Q6yxkw
4B/Ao6ZcmoVPnJZBmp6ydItMInyUpO/VX8YTHMpvZ5875cLHbA0C1AS1Qz2P1uaK
bVIcVelt19kOFJ9KBB1G/lSSQ4oqd9Tk/I+gyBcxx+v80gjEqJ2eF0Xq3shfv7ff
YAr5rv28Ne2nKBiD49oEWUt2oWmGp2qmjuNsGvdQyU7E4iDt02/7uND2kZ9qj/A+
mRfH1SRsygpcOZjruKxViEWJESKDDLn4LN/nyyf9kM24drx8xDIebmuesBSeBf/Z
AGsBISSXj3cTX7QFoujdJQrtku407yCQvh7s7N1UqBe2LwU+1i8Zz3U/Q+ErtD4u
8YTGjA4Oa7PqDuQP8qRgiIxMA36gI9UBUTPULQ3VqICribXaFBQ+2+HtUgKIdNSx
ZLarlxe+T9ecc0vwX1C+w9GSxnJ3FI4R1ElZaO59c3BdJywbK10yzvsMjrKzTS3C
jHCHv0e0Ysk5jdn38uRD8YEdrpHd5dUsBPBnYiN3RbUFapsr3b7JrPKPWxlWiKpe
GeX50TWfF+ROmrp1h1bAgKLUBovnJXwPzFG77R8CeysS9II55YrlHJk/TG0EPNdG
ludJ7RogNbkzWAzNqguVwknGtMLIixFDakEFax93G8xR8m3PAMU65b3EDps7rEQC
0zZzdxiw/LKKrUV0X56cbRL91b51khdVthq0TniUth4Gn7NNmYW5XBaTwacSbZ+7
PdWbn59gGWcZBaaEfTGqlPLHBj0Lj4+8tmyPeLNO2+kWALfv93l1PSp3nPZRMEah
ESK7bpwUzTe/5JE/GB71O4FQves+/kcKPcuc5/Xt+fCI8yrWlyWxzkSkSWZKCT4x
Fi6G0TreBGT31mPM3fKmV+1rMOWDOgnXXcC9W4fy7nXPCRM43d3BYmMjCbtLh3jA
xk94LQVzZrpvalithSOmCJXF08dk8ov+7LvoaSh/mjmPcFv2MVsfAvYzBaON/qHo
UeiMNdmYEY489lw1df92sHSL3WELyy3qSB36k7tyF5wfTdiYCYpWt7TkMxQh91TP
2VY8unBeGovDEq4WZKPfpe1USjfM0BXnBOWIb8MWqjztPVErTC+SqlR+yHF3Ngip
13etVvOxHEyu7955jhEUpzquxrbhEop/S/z64FZQgfwctV5C8g2X8qQVRfvXlSrs
LhHo8VH/i+eG47Mv24yhcrj9O4O30fGIYTwQSRXxQ8+cpWvS/XjMiTjV4ICy6LgF
eb9b+MdyrcrsjVaRrSSzl0d7CEPYR/Z8tFBk94NfYv5Wa1NMRguGWQTgsXb9srEU
fW299bZSgVWINaiNGsE55LT2wJl/0InhchFflKPpIW9joKH2yZMSNlhi3KRrxyK+
5uNoiSlduZaFQv2T0I3Gv7rXkDWNRJr1jENJ4MHt6N7S6grCzLQ+WQ8Cak85kVTm
Ysw5XjRi3Nn3NM17fMyywJ4NeXfa7Pjz4kCaxDMx2nlprBGAeNnplnW6s36LpW24
w+Yo4pL3GYElx92j1FyLIi+XaK/l2XRe522SRJlEjytikv9NAEERvKn3lUjmgKq/
8aBFa7fW/sZM+eRuOTGjvK5mRgsJS3mpIIq+BL2+Du92fcIf0Xp9ouduv3YrhTqf
5NxZvz19XbnvNnZZmwHLn3hW1gHz4n/4EQkBkG1dizvlrCc+yf3IwAs6kdwoCscS
EPyW+U3QnflDBvnoYFy0DhmSt+mW7gXrkxLDiXQYd0GJW2WGX+fIKvDBJCDYiP7O
l1H8n4FFrKc5lc73w3k77Un/NfjRt13QDRxf16qqGKT4opCYoHI0sRG3UhDzidvy
NnGeBRLr3yEgzGmA/Tc8cEU4xEzuiNblEt1o62SsReb15FFYXSkmRZ9s2m+WEfg9
AvFq9OuY/J3CfZ50UE2vcYtGU1e/byHPbSiOROcT//0WqGu8VMGiRvRgBY5rT3K9
GDrJ3xj1uKsVJEC7DVgwMGzS19ytsE45YtOC7nMAm9F+MNXhY9VtXjse4VDnWpdv
IuAf+9rn1hxEz7OwxZFy2KZXXlBltlO93s62LaV4lOs1C9iexGFxjtk3hQDR7XPk
PVtZCgAZS9gdiNZEv47MTwYQYyYPn5PeCd47bukt3F+uUDs48ftYQGTRhpRftsI7
+H3BHwJZB5LxNfc/n5meRULJ5TDkJPdtT96hY5kx+LAljSJA0xDj6H3rYXpOBYIy
+y9roju1Rcg7/Kp1sMMLrSG36K2zdvK1EnjKpYEVsic4XnJTnYciQslCs8DSwo9g
APMyU+soRAnvqN6oaYAx/5rfWxzG6Lh9La2HdzzkyEfBxTMLniAJ2ENVvQVO4pr8
mSZnil6eSgpAEZoxixk/dPYwrvH4zX7lVPGxUwTH3gJLja3Nvt4SNa+UAYCZ6cpm
lu3VACC1BeGve/zZMDtdJmPIK4/rVklkCo795MaNkLb+BNHMx89U+bF17dy1igeR
mILauku5HalbIs3EnCE8gIRPOYEum22c3mAI9r2fLH6Eg3lQYXk+dSMhKypLfeTK
r9F4PuLb4gQyEXKZbm8qXpWQ7jZKFuqjl/R7AihAQ2KZnAevC7T+PNDeSqpdVYqS
vgI+K2A+YcWotLRTf3+RLstEyZmgh3FqTyLNcxg7gX5joq6iiKhZKmHRDxxK8R+S
z7zHNdPzaWNbXCJ3BAoTcU5TqqOvKvUh2WHVdvqVFv+GmNVkZvyH0LnLh7GZj6T3
pHEP+FLmAqE3i87NB0K/Md48aymKiIGoOA+n/1x6HehMEGdjk2AtvIJ8r3IOb6ls
UPY4HhONMAZp1s/EsyMt9qEDdimc+J0Tk3pGSRsR3LHVVQSwsfFRJTGvLYcEb+BT
ZJDhwEwYZIHgNnoQXUcbNu0CsEeeidsshy+PpyXrH5I2jNgZemXJKlC7D7A+abEi
nz3Gtuc5S0GkcMYNkSSBquI45+ehxVdGC47+bKDUlS1AHXjOyXnt3e+YPHVghSRi
9FMwQN2JO/i6+dfNTlXZGLFdugXUjoX8jy0Wcspwg6ch/mH0Xy++BUDFgOjK8IfY
fbglo5zJU4rf/DbudXJB5puzX8I9uXwlPsMyhoWKDIIeI1cJidjI6bdVkiqa2FgF
q9/SnYQ2n6dMdlffFEJgQhcoeKTkei4wspb5rrkeaUfDE5CD0yJ6iqi9YVqvwOVo
NEQIGKBpV2n3mvmjb1d/pE+DkQClUbWJvLBUjcaQXpJtPE4KGyuOdB+Ay8VRNqKG
ZomEtv4zQ7lh7L0FLygnfy7uR/pH5AKgOMOHOM5iJ8oVrsC8Yq+noG7P8CusZJ23
J/LiJew01W52e7WN/q/qyn5/ZIh26wBppcsBgF7ESTBiyKQqo0F7LL4eLeonwQzN
FD34+Nz5IGBZyLGaxn0QiCUUbETHtNdneInX6cvNlxsS5cvfetBSTIxBA4uPjfIL
Js2851fNY13T0/vPiYooRip3/lCTf6Mh0btmVjZPECBFu+dOcJTnU7xDfNn7kUut
M4lCG6GhWXuFRsnnorCQbVUYR54qqVD9oy4SRffly7CCpDR5GMcRCCU5aNqZuiI3
UmQVK5O6lgAkhpbYelRGadgMn2YgdkuLM6LFK/VgXrq6x7ByJSBiliERt19LprAZ
VfkQq/0ZPRlFHvpZdcG5zhO2l+cWdVRAuWS5Zp2uWDLPuIUfSncKjbBFUbD50hQW
8E5ZF44OYo45+VS0TlCIGh06j6t2C0dVhMJV7DfQtN3GrqnbJTVrCRzyLTvGJjfl
Szfv7bgkjTO17mLHJB1o8IIX0g8OZQyBqNlU5D3GTa2z/Goni8zIwnq62uvkbQPO
aL7w8AkPF1USAjICdfUwvkQlfUA/+b24o1OO1SsQT5L1uY4siS/aYZ/yvHhLtgp0
581t51P9IySTnSJuhLAyY6CJgBG4AkirTrwAgBvpNtbKPtuH9ebB10SlqhsiS00U
9sDzUg+bW2uxJ0MFDDblvVNIgvHkaRrQDuv1gJW1GK6gKKcreZuJwGo9+QfoOfDG
TUItE4LglzeYu4ix6aiZ67vQEhgU/K/kPVCaW9OI9j3gn6RxvQKOfo6ivy6lhCPv
dLep+o43vZLmAvUrjFZEQrgXvFhn7nOQyseHdPdlQxZ+nuSAOd2EeI94Edzg8K24
n0oHrHxEWzYuCrpwVRCjA+VynuZdHMtgolzqEuayx3eCM/lxMeJHWOyLYvUcN8lg
NhtBks/3rQ6CxdVUyJBjIJ8y/bM9m6soGG0So32/swNCEu6E4mPvuSvjLB5VFVVK
pHBYw8d+hwUvoqkHZalRlGpyk9Y+Xbgt3hUFbxfKNA0q3BrbeMp0ly5dF1Fweg8g
RsltYLTUNMjttwtKAAAEl3taSKGIhebpl02QWld1VL+NGnfIATWDG1x7xYqhLE+W
2tI9b6OQmEvyNT1Qmi5dobvXH4Z8Vdgi2ot/EhXPpW1AusCUF4ZGNn8acoWFR+1L
7IDamfjxWgEjsWsZyQTthBoFVwM13MCZm07aGEjHQTODdrkG5HlQirqDvV55dS7D
PRBKRikmJcTKR3bsglv0GWf+8sqjukzU31cSzrhSOb6E7rDYTi1MSuFcnE5H2fU7
iD+LCq9daLEBHyESsDj5I991WQzK0XFu0HfSkWjoBPQxwk0OY3ypxSdhAR1negy/
XLtRTDzna/KJuncaM6J5ZQxHG07jBbjuT0UArA4jKj+O1O1P+xkeTecBeN0rhzsR
WJGawIkycC1GQ7olslhheE2oXuRczlIB/8yYyuXcYKBCUMaX6qjHq3/id7QCJN3V
eglLvExB7qk5Xqmfn7lR8qAp/drAczq+t6xlV0lDzBlB5oXSr5+xQCrsMlfJ/aXo
GJKR8fdtpHe4HCh3+axAe8gPQmsZLyTarrgP4ZK8KBG1R2jmaOLF4j0CsyaNKkB0
QZw/rrX9REK3y9YK/7pr7fEuL4hA/FiGjQTVxxH76Yo62jcU6k69c18AB8WrzPc6
LD0uax9p7wkrxy5cpZlKfcl5PigkckIMNjEvPkOb9UxkE/OSr0by12cXX+8l7ZFp
JZCpbJw/kmgYX3TcXSxTqUVEMVVfYQpCOTtiAQjvn7lOxN1itjXq9OP755dWmpid
n7t9/MK4ZKE7XG1j2m/O0wy4tK/JFiSTIMYu7DTa9FBhD+cF+45HIC4dAEcZxddR
+cQkCsrOwzzjwj53Tsd+yRDt936mrrKFX72IG0443lwMzYt9zWErpJC44JqW9h5p
Jecs+/ow+fahlu8+pq0zQS7xRXW2K3KM+wr8KB8V5gq11F0k/zoDnpfFUqPcIi4u
j/rzspMVvdqUiehi9SvLZ/ukLVVh8eXx+kOfTsz5os85LNviXIgFHFA0aAU5qBHW
XzlBzJIeXK9T+ic4lK+ax+JUPkkWKib3AgcCegYO8UOV41f/TDJM2vb6SDGAmRLo
NcHcKRzZhTkRBfDBINfQYPmxzq1rADnim94oV3DEMLK+EglEo/3RyEK0h3f2ATyE
IIyf9R2mbCeuWZvgqcSi3IsXzruzfEaWHd7tVa7bRPU9zq3rT2sVgBH+tHBIyp/5
1/2HDiB12LIICnzNHuuj4ZJU1ZXpf0+hO9F4M/uByDrw7rWRJrKZXCEmsxmkUU2p
zg6XPbgzYIJxQk0w6XUYox7eM1wvnC5HRfLUOHM82H5zeRtInoNbsbfQkqVKb7N5
OTv/u+L3zgXNuFU+dsVRSSGmpZMTlIFlztkPwYEmKTBMt0pyY6wEQdj//GsO+DTM
L3VOMqcNmlApDcG1egEIOjYJtj+Ko10DPVbrgKrbqcyrqrU3bmhgDHXHCRWR3Ldc
Tt2RKNprLx2E1JIE0exvvnCRQf5BtC1ghwSJCQODk0YatOlnA/PBuG4T8r73h+h0
hMDfH80YLDRiSh39R+zQLpLpBYdMUV6z9TzVhskp9rA2Q7Z3qKv7vjOFHDZ0lgFs
sXBPdyc9EYcQCcZ7+DSBRQV/OgiHjyX1HrnDLnbvbSRNj0sAi2+B0i7KQYSfGC/R
4AxASkdVk0yG0GGbX40ekF267eSzOs7V86SXo9JIFiYb7wrTp+ZSzrVgxu2I2vzg
akUjMVycaUWDYhEk25m3vr6hDgAqeEevMhRdE5/CQdl/Ce4hSEzV3o9Fm2+etiVH
kpnyd48i1dSM8RNeGEhhiMih7tAafBarCASOsTodEQd/QUy3uWibp5bxYFbFS31b
arpp2Xnk+QqPTmae0zLpFsz8bPq00vXAB9+dwMKh37WHORlRndZ8cBdgZq0nDy58
12U2c4waTBjHlZJWq88k2LF8R19hPzlk0WKQxqf/M8JZVl5SKtZ6jRTepeeWGKrJ
b+Ns/R5vUND3LrRVE95Sw7QKS7G/cQA4gSKB/gJ7cNNtAKqJmMPIXVFw977GPUsF
eDyE2LK2hBKFyCOTJN8it2Hel9P1sX2ozqesLPo+2KJ2+6LlzJ6xrIG+c1de7sWc
68YOqTqxKAQADKPEbcO+9xf+0Y5rDJozc4KpDdVSYp+bf6wWG8+XFEizqfn+2sh7
bgP1CJhzjutu8j8yZnekxJRHzKp58dm8RkAxVu/lHlRI9hxFPMopecznnS0Ba161
TFlCn2omT7Fw/eu6eqphrhLl/7tNwDZve3XQiNdxzLieevn/5i+pP9HueC2TF2WD
PoS5hJIqOvzmHZxYykgPAhm1rcVcyhWYWAPri3ApATN3phsPHVYQjf+Gnfpw0/y0
RYn6V90kJ9LurOmDgm+WouOPGPgAQxEWUgnVPlpsG0AYyTRBghULOg1iGLamZ9MG
PU7eS8v1nCZIGLmSQ6ssqcl7qpso6r+2QKnf7YjuT4l6QFGXzglUQVXCnUnvEopV
toFLvbug69iEGSbrNkul2UyToxfct8zJ3w2poSOrYNu0slWTF4Z/1YFcC1hhoxqg
Lzvwf97JWJyUf1lUAGzKz9bGTALBHysLEx/cc6vhlZDFaht2ge5PYOxRhGBk9zI+
3L57j9qBXQLJhS9NNiByC1YAKtq9pmSLTNPcF1z8Rwy6rEj8dp52Tw8Zd6O9c7w+
4RxX0Q9H+Zpk59ez4qBIN5wfvRB+hXfXJeBr14jjS6hEjGKKIsCyYIPY+ZGhyS/U
DWdEwd7VRW2/rffXRKJTJlf/ZwjOJKFBWdRx1CkGgKqdmu+npGwpisStcZ9tLgGq
W7+MFaDMne6/k2C91ihClWIUT/s6rGr9JYwVWUQz8hOGHEFG5c2+zJAzdVCdLULR
iXe2Gj7gGTJgC4YzDdxM1Sc09uWLrw/SjmujFpnx55WtJDTJg9l/yZOG70gHO386
goRboOlYEtns8WdtIPDyNs0zbCmblnNCrGksWDxW4iSKOYQRLgUQ3urdHCV1U7Rc
8v7cq6tmDWOgFqsTv6DhfDxhWzGPKuKadH42lZ+FqnhasLcnRgs8vByf6FFtFl3P
pOc8ibtqExYlzXCJE3mu2gk28qdHGLZqrX9yOmf4tjhPqgx1d6eWFsexZTXA9gp/
lTxt6T74LgEkbK4Ptm2IAK699lWE7csd3jgEYMlSHES7iIaTaMdGWvRgOc8g7nIf
3Vn72Y+TpZC4w7d+eepE+nfI23xYdzbSjrQ3tTJVAzpXPi7AIfPG2glYb4HnOh+V
efO0Ek2z3Oe5uab0z4JHrlkwJl+9DvYRu35QrGZg0tLYT9vF+Ir+DFXpL1N91d6C
qqizHJrCbQW8CUEdRpZygEy7QRXM6ozrIBCRh3bTIQ53vhePmYy7n4uGVmsteL4A
eYROfUtJUt/wY9IN97xSisNpS0dxKC93TeIDCRoMTdgmzC7+41/iJCYfg1fDHIko
JzcCX4hKAluzNG4qgVhXoHsIwiDj47vO7uo7qy4ADgP5z8TK2ArqAB4Uy/iqnRwf
ulI8C5xIQDabvLLye2Fdoaf6pmWkt406LlypXUnnMWnvZplCoIkK9fYyIuWsxNdS
4aKjI5FUemGFWA/XSJE57WS6bQ9IUCXzOpbFLSrFKzPYfZlKGxndejVeW/W/fNEz
S/0VEP0G64pXNLehvlXy5SmcfMQ7YnRS0THIfBM/ndd8It7HCjEfm2r0JxUIO0pj
zdhPCrO+0uyaSbU8vB8YQu72U2ihUJQK7XAe2tQ1QBmGgoC8psYfkoQhBZdV40Z6
1o5JSMjmX04Yg3KGqJiDKqUGENw8ZiGMFVkqtkQjQLtakNCgY2Nl7FTuADZbX75R
mKQxhJWbrGN+hBgFws46ikWEBMBeLasNTE96r7QvLyucgCHWTkG2G2+CLI/tWmC3
dwa4UANVcm7SrCITN7Es+acZrbXtTXqj1ht/9JKPkvKLOFiP0nEHQ0jj+wt8rbWF
7ZueRevelFmJYQ7O0URShur3EyGfxn39j7IH78QP9BjcSw6MgWpQppCPupp92jvG
wq2ok2PP/0FNscQXrjExCnP13djiY44I+IIX/KK6Ss+YG98FQZWBz8g1J9r4pew3
F05wF+g31nqRhy82jqrKHqGTuGpyYw4LyMw8ADEpTE+DBA1txz/dut74agC8EWF/
zcef6tosiYcaMxxKv5byb3DVTjw87FVyfCfUJCrs0aKk+LK25+LlpqDX7xVb/YWc
l47wQJDvEe1ZacZEcZdgkRsG1EtoZwdz4u0964/A5NRydT9RqHRePh1q5MRGMGEf
H31wlT3SSJS4css+3ibVIN7zHq2qPpVXSIClJyL7vyBSiCn3irt+zagyUttj1faC
K5Ci0UzBw3MirezxLUxswGczOk4wmFw5dUMSa7fJZupCNnit9UQJ11bVUKMKDrUV
fxZfsuQih0cnWYK7LddfMyohDHmBrZLso6BoLx2gXiSxUOP7ZnxA7Oq9XxTrOchO
wV4VZDhrSYvYY+iGx5h6JZaM4Zpn/43ywz3pGjC13ZztesEgA5T+ylfehfi2mQo+
yg3gDIuT+bSYDuCSM5SE3mcOp6O0XdxU651Ocy4MM6J6AYpnW9GgwDRwlWyfc+fa
Zhb8S3PEkrg4GDUDLfzSwRYLKOT3XcGbqq2umJxvHhpaH8pG1y5nbGjUBMPpc4bH
DWBrM6ajobdQYX620Q3lfiqmUaqYFk7hGgV0Vp/UO82ni4+hNnPiXnd//bMEjcpT
2BLacf26agWL9N1thP3JXuOdg6CFcZAOEZ5pfFLDhfCcpvFl8woF5L163oQmb7dS
i8SVcsjpleqf1+WDEL+7Q8sIv8/gC7xsNqi11HUcqzU5g5n91+msyBc2KbvdiZ9A
OKN1joqdCN30Tg2RFaDj6gqGdS7shdtHjpRunJSVgANPNKxA+S7bjNSv0S80p11h
ECiPOhkWuAPfitWvX8u10fJPijAu4FecyVdTMQ9C9tAQk3i08ug9q0h8INdpEQN+
EBGzjFcBF04SBiZwSwjzJ3k6ZECwE3UhBJFWQ2bW6j9p/h935uDCqPnTOAbEMnQy
P5ja/OlyC5VRF1J7hGlKMeF938Efn5CVEas9qR+xk7znj1ZgvwBwwbkj41ljb20R
VcLApdohZcdDMrtJQ1widZ2o0NDYgxUoKFDTmfqPXZtVLfdNPIa1ZuHo/V/9VzHN
cEqNMDKvOJ1LHAK7ONjCSu2OaVig2YZS9yfi/7a6fOqorFvMuJU3bWTDROqPAduf
pNQiofbEOeLBlTh8YGdD+qQCH4DJ4bprufmxy2HoKzyxn8/pP2Duk3GfbRazI1u/
zN7PP3qqeZD2IYUJ4nic9JJWQc1+Z5YTgyDFBhXLSC+u5ww3s+bm6+w9Bf0c9gzD
ROKz7seybpXz2GHaIdnwi1vUzot6o2tqVG2DAkeP1kIiEFqb2Vpr7q1XlX3ic7db
wu3nBklbcozVUuiVAfYrDRjuoTxeBKUq+xPRYWE6zN2wsse/mkq1fgHhwQSmn/Ns
YpFx6gy7ihk+tIIEf3k0RoLG/3BUXzX1Ml+I1A3WxVhc4fFMAu8uYqhh0FqTTCh4
5bw7wAPzwK/Q8Q6FbnARAtsE3GlvXpT1dQpcNX31NWPmWHm5h8snRmmN5EDlQcsn
rnKkvqlSsqfSAyrDgCXW+bcw1H+tF9J60ufHUyCKcwU/BqV8sUuFA19rsnjb0J72
/OLcgz/1DzMMNAgzPzvRlpgwZmqjn5W+mr+lz7Ct2RSRpxrZ9QmFnCqdQX0K3n65
xYhV5v9UPcoNv2O8oxbOyjpsPIjX9mvRqi8IZTwEKWkUuYM0a/wvUzPROgEZs2l5
eAQgfb7RtphzluEYxXouJUqt2xzP5kzDMPEipZqRvhTMD8YQa19xRg7NKLBzoROO
TVbr8V6BPRaw6KJVdfGtvihnVoW1t9zqcxNp+dvne6WaDWgpykaDH6m12pte4zxw
WxpV92I8VPwKK3TJAQLrNmbyztA59QUQ4j8MGf9hQ/8mCRuVPtWHLE3VIKw98cJ0
IRn8Fn44nEauar/sJxU/iNgBOWfzYSzA7/pId3ZNcSzTWvrXw2ZNNUL/Xm2iGhZE
Zh2h0yJfP0etpLV0NbmjEDzJSsGSU8l8k1mFPokKF4SaxPk/Oi4j6mAkM99N1qFI
TU+jvhggj7sUJXJH8/nsqyEtlwLGdKOJGyrcnbt+cqu+XFNtLXT8sb8RPcxF/PXy
SZrYIf3xnTmayNjcuuSHXY5NOSgew6NobR2OkpLawpsbmHxtwWrY57RAvygWjKrZ
2o7yJxkg7wTT9qTuL1/+rT+O8n8yOxOSknHEm9DHjnokcq9YPGPrBLhIa8MNjVDl
PpHrODagJ+tx5jPPY363LpcExWkKMPpZIoRtT5WZe2OfHbNwM2VXZgsm7YkrtMhN
jbxqYkQLmMZls2LjWL/1/ag4cwU86hBCHtpneQC62sHSFDhF7M52qUfSC+hybDCj
+TwPzJONwwmjt3+Z416VpXajumhtK9I7XskjBHgQSZpWEpwph78ukak+RZUkm00Q
iN9Xcd2onTmNSkXW71Qu4LGFs+IeiUkV20HPUpIGeR4wW+wT53YsSSeEvePGPbzM
qll8M/CYDVtabZkyEQ5mALXpauRGJy7jads7TVTJW6q+2mqnkG0giGNn9P+2/4nt
dE5V6lqgi4Pmt2W4r+Lu9zhCsKMYWZBrvteaO3nO5cGq3ZZGxQkGxTRHQxzwgMCD
4qXIM1lK+/yPcXeyHqii9SIlEQMsE+wnIe6YcSmMCESX7jM7hb+h9cESLB+OVx9N
ZD0NQH44KQ17d+W6Bijnu875yOvgiNsYXbLigrJMDc32ts03SMARuJRc1JipeeSB
m13zRQ7njM38nkghj9jR57ROuH6Xsvat9tbkEg5Ud7zMo56wij+8KYMchlwar08B
mSIGjUf3l1GTAE/N9qYlXUXaYOOW6wsUKQilOk1MNEzmN225x11GYEpmLKgUEFg3
Kb/TlDUYfxynBl5n+d54gvYqnN4oPzfsg8SB42J1jm0VtdOci+sMB0vpsiwuJAFj
/piDxstA6zLQoXGjqtpGgnakZkGVzg7ThNQD99/Wm335uiZW0DXfiwUlHDXVOq8v
owwK/iRZkMeU9nDsxg6SaN/veZAlbKOdEOwIXXeze8j+pxkrcN8tjIM2CE9lc/r6
TJdU84A6zEcKS6FLW+uk9b3Ju0AMK4mKq6nrIq4lBkPFoSTeyzJ270ITuaXJwWfe
sTd7dDL7bh/R0xp24B6XD8fex8EWX/jEuKDQGEad/Zrmd4xbpn5Dy6OsM0Qb4pir
iCqpIEDUl2prqN+1oFZJGXN//ynxVXfZNJ16hu4v3L/ZzIeXbtQXxF/NAoGVHu+L
3Xyyo5rNcW1aVYIF+ThQp+9clMy/C5SKw1LXWClwlYDYCeZAdvZ1f3W1wmI9yNPM
yKO9epRB0OZ+mCzjWSMNfRirOIInsr/zdAhGyWcx6CjSa8vldYU6f5+6sbtly8/q
vtMm9A52Q5o6Zoi8HaKMzsKEPhJiJBoqHgLeN9cPnx/VolT4DJ5jr9voFYlmy25z
KOT3grDEACD2oCOPrw6P7m5tvYk8YJTl6CvEfXZYwtYe7bLCyjy4c0kdCcmOebBJ
nWqy4Z+Gzv9guRM5b7augOZrJx0DBZlneUeTBhIe7Z/0ArcJ0E8qI09ejwJCesOc
e711KAc7+HIqM1aXRsMrdIB6DRK3DmaoJvhZpOHFMyNTpJpE2XLjEoaWvNMYaPOE
X6zjS8fRPbtjsl4kzFMBLx8ovoCq0E+teOj+CoU2raZdm0vu2DQtMv+7gDZ63bjN
sy3QtHFpK6Begc4M0I1xWm87PctmssDsQGRInJxjVOMKoO+oUlgD+mUjIUJqQV7X
Nlgkk41YIUZUPIXjDpyWbi1InswJDSnCAujpVmCWyMiWY0I3bwfuAhGL7Sze7DfM
x4vhnnTM3NjKujZWDM8basrr9MMxuDq5oMc3nViBoQBbVfADtA0almp20tq1xHxo
ptui7lYGHA57pGpkziXCTScO+aLiF6SgWHY7sPYUcmkbTNqWXADbJsQdjXL1G7q5
PjaxO0Sx9WYm5as97gMaI2ZMQwWkq74nudT7eTGhY9HJizs6lvgEBbfMPJx8eJY2
5VJ2Aj9nR93FtckM1Sl/se/s117aMOaALf4bHkEx9BftbXibQjp3pTjSLryBbOML
z+rXpjMzlinq6ihXcP8SZuxpUa5VrY3IYtpYCgBWKduNcpfOEf1SG5YUcPe1qK5H
1IWoX2Cci6tKnt8/YrBjjNavU0bawcmfym/RFvpUQjRbz/y9NqW6D3wOPtROUqAg
70pQ29BVE8/mRooRI4xrr7OxcHSiYVZWP1TaJupILoT6wAeujWUCeWRtF2lPaLUa
gbNtWokDf9dAIKLg4aWiza4kj8IvGfgOqTSHaJmhJDaI5v32DT/9dcupu01WKNey
1zUzlDD22YmPXR1ettVYkHcJAO5ATHZiXQBr3BmwWLzQ9IFixGGXj/iY7vQRCJbl
tjlLdczDN/oWJD6et83SETb+M2zmIF/vqnBGqNTS1ocgSNYybN5oKQtcY3ZE4kvR
VpGOXmCCd7KUsQNkEFtKIPdtdvhv9xWKyePrA+hbOEqEyS7j+98K7mkGPjGTt2VV
2JzznRJGceHyc6EjEhCYBftp+QxPsHMaXyKKhCfx2Ec+00VEC/qqcGogMsOH7KSF
8ZBw0g/twEp8OQO5hUXgTSogWBkguP2zOhd0IVXQa5c36q7zZzxyeh3RhPgvcbS6
XaBJ7/VCgPRTdorKE72z459M56DZHjtImYa6MP/zpS0Fg+S0N8l5HWUj2t/9ZerA
IVFvZRvFn0xXWjrQ+emKpnlask3ALu6tmDv5y7NrMmPRANxF77JH0VipR2xkf/82
tsucE5qbXonjJUMGaKKqk/xdCEhw8DrkY5H0sAbQVenOJgnoEvd7uHJEvz7tGVNS
lkVDUaQVl1/kbS2oiuywqYz5yL+ZnavKKxfRv/G6Q6b11ddlFdKrwpau/MCMCx6Y
9GBdakeggU5DesmNP8fSIFpCux1iovJ6jIEZtYfDflVYDCpPVIaqNGTKl0cYp3Hh
SKBCGueWCj3YiSGgfMlXaTbS1VHQS1G6AeSwPf7UTwkVdtAK8jS4TF7pQUIsFamo
dlN9XpD1758K/H4ll66p546dfF9DH8pRE5zvWkHhc2j5qZe1dgUxkYVu2ymf5G86
FoOMToQIBAgwFglzWLSlaLiemcxkoRUOgZulTQfruFxMrQ7Emxl3KRBkfV0zyGYK
33h4tR0/cLs648aZNesASaA9gqtLqsdrpj8tJSaeLHxWZli/ERoeANHfnKNB3tBG
YwX4PuNJIGFx4OasL/gLJBnmx+esk2wiwWfWgu8hzReaXcki3jIaDqIi4dkH3/eA
WSAiKOdkthpnA8KE47feKKDFBvjFogZowpddmx3lWMC48VMYMDatcl2POijJOCKg
Tg2P6j5pgz9wyvjGtOnL1AjbzDFmGbPCLeU/sCNwqggf3jYS3av1hOW4aB6KbmH9
2OTEJpxE7L3SmmPPshs1e2OydDSbpIsgG5o2PRZ1LP2K93Xw0iNb50NmCCLrkPsO
7q6TLooHcz8mo5Md6PFDVCpB3eAJ88i0x0BWsroBJbs5jD+o7TGquG3Wu/TaHhiW
MYYDR3q1aihMqEv4l1SHohuEN1QFGLIvicyg89nhJYIOi0nbv49/O4YE/oqTce8F
C0f4zE7tnHRwYCByvp8itMb3F3M7bOVAkUP+jeRGi5ARt1PaMdW90xHCSMTv/lfh
ROtoHVhfnPK18aLCMJOtHmMSgXDMAACOJyVvx7INWgv/AYvxZim1qP35B/l2ctt3
vpBSt+aYqBIeVQK7j8Ee3aIloR6h8vhEEjEqbvvm2JaRADSTjIKhHC340L+7Fym6
YtmksehLDbK5zfAvPRj5wuyAJoHFwNmoqXipKjmgCtk+NaTsphnWBd2uWJz5a7Z4
syddlKeMliW25s8VFt2yZE+u1AreefCaixJTe8RsPaPMx9W/AlSHMf/v3vgUGzmp
feYNuMb43YP/aDrN1D+wnjE4IYH3rZ/tNf95Lm2PO+UXfLWOtLfOAbMtBeAYhZv0
QdInUTUh58HgoKHGJyQkBT8KpWK896vmgHQanYmV032NmAMEgxm3Sh/rBWNhcC6F
MT19XgROiFKlxlECqHHJM7uRCtYQ+ygpMXFWntbYQREJ+BzEW/QfNTP5D+9WofP6
+IZa+sVfyuPtyMIZWHi9E+OX+cue6JPeYy/yuuveUzHfZwuqqZWy5CG/wtrCax0F
tlgnp/lMp+sUuAEH+vQdEDoAc/BCuqJNfGQ3Y/5JpV7xQxbuehBtgETZ+O/GG94t
+6hpv3dZKwIOzdkieVTjmaa26Slig7HXeYlVRprWRFFHVZoqU1nbn0KmFeGNZCKb
4A9hqGvFmmSkjKtW8OfyzjTY0czc9tjkdT6PfgVDAJLveASbFhvlagpib1057MB+
/DfgG8lVF/YeeyFCvHm8a1ljZzkPu7v33KVtEiEmC/nCeQbljajPbwuoXegyb7Ua
S00VXihBSRfbFQe7hykYwb79b6IZJ7snhqxt4SD+4u89/IxxEbkn2wEhaFn3nP4k
m23PGGYIYKOJeenR9sJbrn8ZZPWl6CnSR383qLJctv2kr+rl+wV9yGkkQzCcofWW
+nuMI9q3NZOwUr0psMfbjNV1yde2occJNaE1oHmVlctNzx8uo3Rzct7JvH/+rdRV
+u0CoIz6Nrh0EA+Q4tY0LRKOhVAjmwkh9I+CnFF8z1esoHLD+s54S++CzOvV0Wt2
dZvenAgCezTz860XV80/f5ES8DRVBpJBtYwp3G5w3WYzQMl/85xLhrbQ/+MlePXX
3yNGNeWT35CmZ4aIeJgKqmOvuKChni64MxjWFpKFb1yf55fyoy2HfuEBoeTgWUh7
78vXgIPI13tAHsB706P7yNFvgO6l5NeFJ+rzrr0PQRM9hbHs3KMErDpHko970hvs
1FzQuF0m5ZTKOT6Z1WYn7Kd9JbYAZHymReLQXS7LSORlTZeliaMscqJPkdnLnFEN
J7O7WCQzLETjusmqQ3xlOGS9r3rmmUCK0owZU6B20cMjwWvYDSJWDrGMJ/w8ek+a
4IEWijrct5Ee84stnr4ID4PaLEgrFu7i1+EtAntbTqENSlJCCBfIoEcO9lg/0yhl
V0aMTf6T1qmGYIUF5Gw7bKQVRePLsyM7c3C4p7bHGxt2O1QanGgcenH2NU/cBKxU
UPu8o+xmFtIgIUKdJlL0zrHhC++blSYE/vgMEFVH6O7CNkFFeGpS7Zl/ZCtwmRQf
8+daRTARaqh7Kf1uTwmf7P9xX2TeRoTJsaSr8Ffb/foyBHtz6J5YVWMQAYkTREOZ
n/92E5EB9sONl809iLfOsBVE5GTvzmkNGtFvON+OnTakb5xYgNROPQdFUWwxXySe
Bv0aalHfBemFRwrTMs5rutAztRbv+4kxRAG054ksklGwZY161cD/+IDgXbix0yIW
MKHIH02aCspNqh7rTXpWpTZZBqWTM75a27VDdbRefF1xE2vUlL6dG07u44Sp7e7i
ACiAnUckO/DzCdOjqXpSjyIK+ClTGXqEVv7RPqB508297REDNvcv+OZpdihw/ae+
S0hm/3g6WeLuRq/z+d+wB12dwDElgM8ysBdSTuNBLAWsvkCD8oOPfETcBcFDS4l7
9s76ohOBsAnikwjBXckJLkQ/xPS1EubmFxa6BT8KlrJ6oxGM7+n85aMIQld6YdPR
o6hfBI/584Ja8D2j9hCv7rf33w9f3Zbp1lZMrsOEMIJH25acj4ufjyvRfpczJZY5
T9KLjvOeM5TBxqwF7LX9SWVWsw7OD52FZbndV95V2+u3w/O2cDzoysjSd286OXpb
VEXvuqAUNdKoiqoTE6ksUQoOh5mMxYxZip6e1801bwrOQhfIf31RroDOJxrefxRk
BHPL2FqWWM89amJwW5T7cuC633hTTqXS/YLc+24LSDathD87+zOleud5GJaZzmI2
AP1vWWmmeqasYj/i2n1I6ctkzm61w24SYykzzfrfPwaZoKfwTAYRaDKedEch6sVd
//mjNaqQCNMDNpB/1418XPn2L40ExHZHwqti4lUwRMDZ1TQHjwl5gZ7PgGo/YUyA
6JlXlZtwVEe9kSHimi2S9cWq2Cw6PtRTYqZiRLgHv1z0Bqv6eTHsAnSOu8vvGS2h
BZs2TEhF9iQe1SingCwOm9CIp7a758rZ3Tpu8w4DcBXWSpFKeCyrqNHLZEIuJm4q
u8dIgUUFMTwLqHTkWPD6FQEmhaOIyI0r3ddQrWB17Pzv/OhLj/CCap5arKLeRYxY
l4/EHpVGVN7Lh27fUfT2krZT8WWtI4BXSNIhh4QLxnwoB2cD/9GjDWQcRDhTiONx
N3QxinyCZNmbZrZgrmcClXv3k/dlhRZqnwYyJjn6m8p91U07a2rVyjt482soSo12
ww3uYRqhTbht8ttD0h4mpk0XuzLxaua57iKhzFK3usP8yHDGbIg8JfwkBcRLbgBw
DGdb3tJTJQnGX9k1lDoI3apTdlVkMASt8CL2UvI/O+B+AuMezKkyCPCkcwNTHEOE
g6RGsN3Kg7963iLImkmCc4xpZgo5K61/mVYqdgpe4wd3wHp0RAgJYczrCoTVpY7U
6pwi0olmOjg7ALTsmFliIv8K836nUROES7DyOM9KYy7XYmaxg9MgEcX91bKrz81l
TB8fAx/667NCMUx49ICzky8vBWzs8Mty81sR2wycytk/UIoBQoC6GW03s1bDBoCd
FNa6eHMF4FirpxG6+8TKtmIKuqlAQ8IkomkCYTcdpLGEecJzHAW7he8FvkqY+OE3
JRhWTh+m3mpAe2qPRBubfDpMizBcX72H9tS695RFk15mBMXOpRnc+t8UDcjiJ/KW
5MiB1AYaOiTz2jcVYlOuQEl8hscxBBarmvlw6TcQs/twna/xFu7LrPK8c2osJil0
Mu6MNcHfs4YetyiKwx6oeuB2w+5PhmYPASCuon+ynErqS7FMosiLz6Xuk8wKYPdD
Xm3zBlxcoVwTo1xU2umezKwSqFi4PEptHuMLd8V/uQamnqQYSjzuACJzYJ6cTJ8d
YnlLvPx3NtEQzxLmLYHxP/1Ie1ZEUqkOsMZBsEOQIRTp8oIR82YgJw5PIjcEqdsu
+QYayNSWNutBqbP4Pws27WAuF7K1QKn6Pgr+ibYmQPNlzFO47An4DWfVMTt5KXo3
fKj2/qA/lGsGEPqLZMqXSNLiEw0lD6UU47o5duhJ96msX2dCpzAsbXwtuQHe1yQd
i4iPsS+esjnOLMse11P72pklBOXFZ/Qz5D2hlQlCbnKcEprwENg9X5pN9rFtt5Fa
wTZZxTAUVxSEuBkw42/AxL6aU77O+6GclpwZsEXkpYr5sFBJ59FDVG85CAi/O+AA
3HupmhAFx4A2aTrBG+rXKBDalU40F4dDfNrsFaOf+C+pr3lsrrEiugWOaQZiP5Nk
EVvFZRmsma8ACeGslh0hefDZ/lDl8UzhqmXk6ByNz174dQGXO6L+G9pPT2vHTSU6
eiPmUK4csuDS9EJmiEIhd0cjGh8TW7gAvkQHraQjn8cBYvCsZzBEtf703pzfcjyd
nIMyUMnclPM9viEnInlQL40aqsXBkvtqFtgo6TdBYz1oviDJO8A2e8lDrroFv6Xp
znllqmGk4hkT8OR2Ab4rNxz/5itTXQuAUzVyxgOvrJSUeNRdeDguO+E/2VSRJUaq
/+do+UX4hZgvY/TQwpXjmKufTQLX6VQFtxwrGTngyCS0tCHgrf5deCetQYPORK/p
8hbQpuyhK13hee0D14S4y1wJroxlakyyfuY32wZy/VTabixOOZu1b22Xeezi0Pjq
sD3mpWRT2GX/cpFuY6tyeSdIzFH3FikMXzC5OhycUrIq4la/a920BviiuJ48Dqvz
VmfKnWhlxj96gBd0OrVBfZmUyEt+QobjQLK6ybLUUUD+HSVSIiMzKsPp2N/LWBib
+gFtgYvsn2mLsn8sLXFzrAylE/CubFdjRsY/3/zstqJb2i9tj6vgANDpDeLBFp+J
pYvyccWb759hMNzO80tpL5rFmaPVsup80iwbwiYhPP+9a1Mz7czsr/2lCCkMe2oU
S7cJhOeiAZzhTfSQl8BPs6pjHKYnP/JynEDWIEnKOtE0OVgRr1egJZWVQf6Anb+X
jTilz/UvzqamVb5VMcooT/XEhEp/kI1zKg6Cy6rRzvhLtFueuAuqb09+Et50wKMw
2SVTA5tfVAzOUXJLUIEPiPpe7lvIKV/IkuStJHYkJsfS0Aj3p2jONAFL+XgG1OdA
0GNg8kYEvfuAxf6epJIxlLDSboyr64u8pwiYZel/k1t2qNfUvH5xcmcM8yNTjobl
uokMXNRm2ioc2tP5g84y5vxH6EeW5BTSzv7w3yUnC3CtkIaeuNF9iMqlfz7gmYIS
yl1JrjFPtD8EY5mMuBtex8Fjyc3mojvXDR+KanpWAz1zy2bNG7bedlgWlqkAmvcF
sBRRf+OUFpdb8zjuwYuv0vbtDnaqRKyJTYIdJoT3t7h0wOoOYOphoOkYxOV0T5z/
WpdmH8jS44jXQZrcvpe4ewBb6IRDSPSRxm4cSXgBGWcguZXIu/kNzUaUVuTb4tD8
cvK0wK2F/GhWgPPLKL23UNhCtpMNJd19L8vpR0DT7dsXPyJsmTNhuv60Mn6ZpnmG
lIaMZuwq3+vTBakrADUTzUtBQyfHb6EXE9tfbT87MR5fFKP+dnRi/F7KODiSP0eP
4U/xoTBRplEHZ/3wI9h4pCUZl1VmbX2rEk37nbQJm5Wp6ndL/YOgwAS0OuPU0wcH
1uyof/7PcZGJBHf2AGOmcWQMBhfvBjJgNlpqmW3NdbnqA4kQ2woZTm2UtR8dCmeQ
hUKVRlswpXMNs8/+RVD60wpXS/XbN5TF2vsSVCVN97BfqjGmC3Q2r+iBCvt8Yfzt
zdkwbkFP96dEZRedE44quSneGYOGXQS8BtHO7ENMWCBwnNQEPnJviZ7l+dk3I34Z
S9KTkCi6V1JOZ6nyZEue8G+IBPdfavWC7NHgkBTXmX10go/XVU6kvWT1JvCqjZDm
+GLUZIN7pntC7CdLILiQu9ocwJ9gre87k3AeXv1EPuOXYs9QIVY1t+7lhXUoT8B8
D+MBOQ+nk+mDHK3lZxdQggh9BBD/+DobgOAtN22sO9YpYhm77CMLL+IxxxTW+hWw
Jd1lmN4ZZSq+BxsrrkUW3bjBJNyi2bVMoTo6sx4ITriO6S1FO3As16pjCdLzSPO3
82oJ/22kdKfrgC14hMuA3AGVIG0pF8HZDTOod8bcTx6i76656ZxAKEM2ZZW+JZSa
5sn2mdGWoewIwAABl7/4jAKmKH9GI373ucu335PpqcSCS3/CIUG/xqsfT6dhRjRR
PVc6krjKkv7HXpTmm1E5uzvOV1SRgfuS2hky8TEmLCJo3htHtG4mbi07vS/mwydb
ntj3rQxAXzYYnK5CPXXx5TWj3IPQmzVwspJm4T//pGuIMxALontbrqLJ3hVV+xD7
bgBFdjS3c9HYchpkl6BTKT18XDly62gG6w2qt5WHt+JdqsOZyZhX7rTtrADbgcj0
tCDC5+0VIeant16EZtcw9VN89nMeveGgvvpzEdFV9LQp3PCADUcWJTIOLKm+8X7f
GZnYaA1yXCU5vOO6Vl91WsNpbdL6VkNq2+Es7XHrPzxT8AbDOMQuY9u60Q79/gdV
F10H/bwEyM4vqFJ5NNxkB5RFKxTameJcq+gzbnNkTVOLVP2jzNShMJmiUYTOjJtJ
KMBJdr2bi1NJsWQt8TY16MaNi1U6CmnTW/tTACbejbpltmGWHJHMqkI7ORw3fhXC
9MYrDRCM7QNMHQkfngT+KvtvcWrEMiAks5pkoEMWok2oJW1Xc9zrvAQGiSGNnUzy
mU37EDodoWIgtaXSColJiUxJgUEKUvhuXfEAiJzVdhm3VzN1xPdTsgGf1oajaMwS
wlnGIMxCiSD1Nr21v4BlYr6c+s6dAPATUilcS9Q2kjR39nsLhBMRse38sw30JZWT
QvVf/w8yafeP05A3cntD6tjv0MhpmQZGK2YISWzH1NTXPkDSi1AcjK/9orkN2TrC
sR0Wk3XM0Z/udUmG97Sd3XK8NfT1EIOQBxM1UxgH3VkeU0Lgvnam3PmTABM2fp4M
k9asR3aLh2AAY4lNMIN2FkiUtI2d1wmnZGoU1R3b4tS74ojzcTYuAam+zOZw+ucB
GerXYFQu2zPwPOJmzLePWKYbxX7eLw1nZUtdwupBeS0+GwDwQHmuczwOSrJna3fy
oLYRCZts6VBIiOTsV1W7H6sH+znevykoFg5dhZYVJA4nl5c4ay2WMu78NRlyXOtE
U/uBTrmNuIlwaB43W+tpJkdLw3riHKqcWu7hbfIp87GW3DFt6dmDYiT6807fTfCA
FUyMHoylHwwNSUOr4geHgAnoFVc94D+eES5A3yL4f1075wB9dwjMNq5DbFDbHowh
rZj58nwPwR4NMpeOuvxGC+CpVKG2TyA2+tnOxdotypc8d+sN+B9XRR7XRwmrFBZr
XvkRJHtnR0qw58CBeTQSbjozYrNzJEJWdK2O3B0trFxGdNumf7pO8qLfrfoz/KGL
njiLTEjOU0CZMhYumloJEaC0yooFWQZv636yTk12je+36OfdR7rho1cfE7zLeFS4
gkNaznATef7R2VXGE4ltjyL+MlrmJkz7ynRn0oOxMIB0frbjZv5MLFfPvp3x6+LY
+hlEQwCAAwuhlcmHRHHgnsIFMSKq4uSAZhFQVKxw03ng+bNm1PiQVtHyClfBXeTN
/gAGM8sES3ICWBUrr5qpeznZh114VYeyCKqggewCzSbNJOqkKfDWNnNjqhhM7i4E
TjNgcPXVCPOn+M0lcnwy8ORxPIwb2gj6X2OxzyjGxAG94HWe727PY1qZ5W1ZcYzs
l//OniD+WV9xN5TxZS2zFxpuKRc0kQKai5yx7ISAUuCt6KR+UIndrommNJVk3rKc
Uf9Z9wTEpzti+nW0ll14IfMOEB+IFbyCCbQRmgPhondJrNb5iw0ZxZQGO3EilGh8
pF1qgP8xBJDzfHOuVfHLLY53Gfx71hkP+5tnMbqB6YpMR6AK/3DnpCYtlkNRRKdU
Z7YedyWOLSKDD8K0bi3CDKvZCVnqnYTuyv9E/CJ3uyGOQc44sVYTWhwsqAJmVZ32
d46pO2mONaHwwOEH28IFwuJBaDl8QrLyTjV1xz3OkEc/fkws05vjujrOtaz7Py2z
4EwF8Dvg4TWZhokE9KuLgkF6BbxlWffJST83arnkBqS/7JPWZFhaKNfiL8Odx6QR
e55Qb3+1zZKkd1pS1LwI0J1ImWmlpKS5NiUio/tenJrvYiORkSzjZepuwQEDD/F1
4lNaCYkL8LFOqy8UzKFg+I3Q46BHxVWBTELmUaOwPxNVIUrQDHleiTzSLlf5uMl4
nMgGb939XqSHFgFAOO/SDSHFs1vzZ6+BieGLKQL85gM7wvAWrJdQEIEv6w1yBWrO
w9oh+MR+5ZVo+g8gSyqJZYlibKnx9QILs2cPYJ22LBDC7dsEloLCuWVPf2wLLLny
n8vGQBqgNlozXUibinrnwu1oDZyTf1BHflEAMzbFQuiK8S57l4VyZNhb3WUaeX4u
klG8rXH+y3mO2r4wasBBJK/Uenf8s4/M6q6oI3wKAdygVzl64tKrQ897pHMz8ALK
PN490xm1WNdqQ3p1oyt9bvLwLTGwEDpMee+y1wZSG/bLKddz6O1DTe8kiFMPjgVP
qpH0FyRNvjZ9T9+7eZ4cNQzus1AGiJsZBWYT9umAuRLEtquDOiBNWx19NDI9t8uS
8mv37hWiVOBvRM5VSGEtuqZrPjL/bK8MlhLLONgz0quub/PvaE/JQbYm2pMHdIta
BT8JP5t4mmxqT7Pcq39/qjicQCiJyp/3Jt+1O+YPPzM7gyaeiO/8+kUolIxM3Pc2
avbhug1R76ApE2BNM8qMYH5TLRS97FZluujSJt51WzuQYU5RRMGbooZAIywX5PWq
Ey9iqBqkx2SM+a7w7lEDgxvAE+l//3uL4O+INJryjdkLvxPv3sIusm5F8C/MfzP5
CvoN01xQu5M8o8V31uBI4oslgWqgZahc5VGXU2gmhc7nXGxaxPQbbjedmCpv2EeY
Q8x8dKdAedSQkQsCVU4dojGmWgzbZ23taRXhA/bkYeF91YSs8+pQBNdxXOnPHy6j
YZvMlxQUTUZuh4J65bdANTog+Ph6Jv1G1ZT1vnRVOAyo3/mEswQhu0F5pSonkJbU
RdpOJ8WhDSZwYwvKqAFkwWpQqyj3a7dGpFUARZ1m6nnensa2w4MdusW0P2ZGiaES
bh8mqpXBkevEfUcjiQClbobq50Z500n8/12emkZBmmCxjYSjVycQaDox0THR/n3H
SwY7VBxY8tPnTSh/T2kdJZdHU1GZKXf01tJQUl9eZPMAf3UV0MI5M29LgGjbY8Qf
wgB/k5StujfdhITqhVHu+MXqeGdiUykJNo4bNzAEzPmapvSoQXXqWKjfPo//jhs0
IfzURiocHt2FLJY8VXKfMj45S2gSbyANjrivNbCyrI4P0et0gE3LGyirhmlSdkoB
zIwi3/ILNKtZH1WJVhw52Q2sfA8J9RajhlEFQZWG3cwgvnd/BPO3QrbpW4nbz3Xx
tJaIqvwYHB4X5ARo8GEu1mDi/Uev4D8WOY7peJKWscNqfb1V3Ib3AYqpeVHwvkyB
FfJY7k2QTGVlg9Tt7o7t11Ujmj7a7kqTBsBh7V6wYQzRfkm9P1xTsae5xC9LuSCx
+Fadj9NdePKddTtdrLYdg1wkagX5Ul+GFEtY2soUaPXJpE1Ufo8+MVI7Rgnq05xD
CSQ6pMEkdj0q8ghhbf1+m6W9clz7HWXf/l9s29V7MWvBICiUU0JLZr6+6gpaXoC3
Vude0BUhY9vxyr8ZrNwvvUHZ6gVi9ZIKb5/TzCJrhkiJcfWDpXma0uwQ4XRxq15a
4QlNa4FFfKsqhTz+bnwAFZ3azjBOSK34r94xhxiwedHFu4zMVk6F9hy47c+Lbl4N
x9KQULirHX4EuItaAi90sMnhIo0MSuBi8+XEvJ0URq5azrCgFEkn98PaUzNPYjRe
l7jbt2bwzwR4PWruNl81itxya582wmYnq7SGWTRtpSxAxc2dtM+1opkdlIhJlede
xkfZOH5WNCLIvOIeCfXKVifRkgzBfepnctRMVR3onIUsmMtgiiwYBKrzS6DNXVqN
i4K0ogijr/MhmQoqb8Hr75DewWuuYzE4SKwgYB4Ckx6NhsdQTEjvN47GWuhvWUXi
WIUR9roDFzwzDyRQ/l7S7JDoM1Y0UI6I9xrYCxa7MEGnEnau0u1djz7qyyuG8oA1
48NsPqw3hb3YIDVrQx+3c1YMdFiSogiI9tGEGUZk4cM6B+YFYe8/v6Doj1cOb7Jp
eYjN/IkCLLp0QBZod4wInWZjVQRPIemduNpoO6ArfqqTfCXBxzXnxUTgYzZOxNc5
63aBlnmzKLeSN/nASEI5kgceuW6HU9oB+wp0btfEkModOPNCLUfhclulpitB7gSW
S30U/j6nesua6upeFLsRcdlkIlXpmF3eGqwDssqNwTW9cDSKLFp27DudLH2Mth+a
C143v+bKcE8Lo3wxHSiQGW+ujJDW3RcWfPjmeAybMf8T/n0GYB9YGSEiyIrJwL11
sKJFbQxnxtH+d7ObQ5s4Lcxb3qmJPuEjfPcUez6RRvQ9L2z5YlWvX6CXzHr9bqg9
L+Gs/ZFArEv7SC+nne5B3DnBxaBfdhozJ4kKl1jIzsN0muqwACmryyAztlMJiE71
LnGRfDmFTG2budDdj+Apg4RCrMGiedoZd84MO7Fs5rv8hl2XVpczKTU5uAqUZ/Vs
X/SlkzQsV6KvrVR0yjmW8aSf3/oF/nGBi2LnRgDSKibQYWL+7a5KWZ/b+2t7Rc65
MgVmMXZHPetDhFhuU5pFzycyudjQhBjW7RtQO1SbTLYbiSR9da4w8pjke7P0/ucc
bX10DjQSmrB/T5lfyI9Y9/yOuA9enRbzJkhwdExoVg3w4TBK3ibVzYp0tEo57eHf
7Vk+4rbLb7funYFEdEKc37FuLDD4TjyWbPqU/QYKFQR3giSj6UXwV6VYhL09VnFo
OdGIcpn2/Lu77Y2/T5rSbGZq3W8SGnxCzsxk+a/aVET+yr4NN7kWiQikA3mRwFgN
fWge6y0402N9XwM0vPSkmD9FuQ+UbYNNeiZv4Hcjw/gEeyTVeZAwYFAojQiBSbhr
u24W6omSkwvBo7yxVnV6FpCUinRAuQ1hyJ0YzVoCZ+bbTpWiFW+NLMjwsBjTPx1/
sCEAnQIsJU2ESV8s6hIoGCUyVowXqfj7L5+hPUuccu/u4ceQCrN/Wh1giusJJrHs
7mrzaJTz3njpzSFoZp0uudToqarsbs/pWiGkTI+Zg2+JdSIDeetdeUjb0vAsQYyA
TiMQL0854Aa3MiajiIw4cMa4jr//KKHDXz83Mbb61da0twKrzTnrw4B65hTHqM3V
dskbV0VKyAkRFxAyovPGiGyz6Nyoc5GIhGT+tsGisys2fuQqp0JBX03sQrauou6u
xndkCEDmirJkNV7cN3s8mcSaI2R/b3bgJhI9jDjIbyGXHjPAPplxjuvWZ9R3AwUb
PwjaSiFyfmvuFSqqZ7spZSPdWtENPht3osJHZaGwFc+bcNU8gXP4MUb57IsOCd6x
CZJWKGOz7fbCDE87nx+0gM73poqI91lYKJYKI8QlS8aSPuce5lvJ7ouMCHzy6yuL
OVL4478pcgZVEGz/rleLLcHCjuVtJiDrkObVYqTdJVXj87CJtJG2QfUfIcVKo6r6
t8ek8Hf3sZr7sYK0c4BhkILAXxslL3++NL4XrvPMK0uwSgGlS3PPUKtQkrPcbXkd
vpGQdC+x+XNKYx9rz3W9JOOfWa6mwMAxk88X+IMN6zdCeGk0Ya7XkMByQMPZrL7i
VBOAGLScYq/79f9AD6mzWdf95Daxn5BivWt67rB/k015OQ3v9cxWjb3L6qWulhEK
QlCK7YNddEddkZKkBg3cKPV88ajlBpbuY+TBKR8qrvxGdqqqKd0WD2Ev7bblrOKF
EvLsFSk70t+g0gslNkLyrzFyUH65HZiKp/DtNVwEdEAdZ1iVQ5LZvNGYMDgja1k0
iBO4mV1GopK2EU+kE2jkr+UkG9kmigUYnyxDM16j+rpmS3S7mBi76DzVLWLmlcdf
57rwXOcCm9ZDgcAVH6pHb34oHI5yqC0N461xLmGGyxUamnMkF8xRsKCKvFewg3yu
0zQ5G9/1tBr78syHC3LpKoSKGc2xTVsHrOCcBFdLpmeebrTtmzWfJZRxXpW8+g/Y
EJP74Qde/WMGs1Dzs26GmWLwdzsPEkdckuzm5EcJwAKzWrQpAqezMa/S7T9fOAcm
kz49c47u6dq063vKAqiE6qcOKgdwBpGtwY6HWZT01TYwkZn77bafQ6c7T1zDN4Qk
cynl8lgR4jpreVv4uUoktz9Xqpk4LAWPnxeefAQspEtZUEWaI4q3V8DOzFTT6qIF
ebHItTFE+/oNo/MGRaJvkKk5S3L+Avgq55cUe2oyBInNvjxkrxvMDVPTCyhQcHUb
UJDsLOyaBC49lknV9wE8i6wsy0bjT69I4jfIMzrUs9+5FZK4lC8+9qjQRR6Y/3/6
SkeYF+ZBdoBWvRc7hhTvXC6tjkgCV0f/mMvJZ4eFjjxuvdqI6P889xA4kN1QCES2
WbrAjTmyeMUl3l/hPTfZfQ+QvXTGXzHibL/c+XLsq/fD2NTlHFhlb8GCqYQinnr5
9bmj39rOuf5AuUWuBDL8oTDZh/Ot/rWvK2Slv/Giliwo21cU97TdgLHpaxyPwwQt
InZf2exhXliyqH7vQtdoxDNe3E3tKWVXLe6nvQe0OIb5dV0hcrclGz/PsWZaBT16
uVizD42xprfns3uHUfc6S85wt8I9tBy9ZshM///NaxmsrR86YvuLjDF8JEKmoD9V
LQQmQWl4g4ttNj9uKq/VTYfqo9BlXAxAsFeP3NekKUJtR1VLbt2QHPuZ3YDc38+L
QrDnwOkBiz/r+O2oq8naBY+N1vTJDdJ+gHkZvwiY0wGBc+FdfYIpjvAZLftprV+y
qnnDUzpmau8v7ggKIqKVuWKQ4bp30U5HIKoHmkISITEQ2wDEQ3vfPfw7trpGc5Z2
aLXV2gFlnmWHm/F5xACmbqJkby6VUMwd6KK0ZRaGd3Bk2ywyqnAgX7Mv/NNYvb23
iiX+9thXhoXn+dX0llAM34EmCVweRtFOEGpREKVn62ZcELXuJysaOqDbw4NsrYL2
/sU2xDye6amhMHvSJxhS1gFtBriG8LdEaRX+oDIYxo31zt12kEVw1TPxPEz6quFu
TbvL4K9j5Fp4OfRWN8SYvCRpefVf3y63/JfNT+/wZkQElY+dyVMFrusg1Ddo0Fgc
ekjkY3HSMsdPjZxa5MDw/vn+mVqh8mbSKU5GSYgYnhEi055WN/pdVevMnJ8Ywn+C
HhyBYYwfONFsCjDq71PbiS7XRIhJZUdoBKgE091YMTK4pl8lDyuvvhFkGXhRrZSn
/iqsI1RDQzO8POXFJ8vcWlB/iFc5G4HjtXBCqQQdl43URoshKb8qNT76nfZBCZJF
z9FaXjE1fTvjLm5Nv2/VQu6lXf+udWqQQSsrHbuxyVr+8UqnK0sgrkweLzmorwwc
WqfvmenJ4Wd7KV0w3QE9ieiqrj2sJOskAQzNGgguYKOUQr6vqNWB0K2K+0j+WkbR
1yv0OE5LWuK9NBHDddcrG2MNaIOK6oHv6NDMhLeCoe0A5fQOX0CXgo0WNKZa/acm
/Emj9fJLUn0IPJVgjErLPX4YcS3LzmNtK3Se09Rlsa6AuRpVLtR2Mp1RxQm8Eq8D
5ehUvu8KG2xX0z2KfCzZWXOQn8HOuum3goli3k1P8gfYsO6OScZw3CLwygPomgxP
ciecDZtsnQiEuhaabKC6nL55NcWfphX5AqaXRlMZhs1jIoSIaIIDCJtgPCJr4zpk
nZCmrBpLs784zkXi8CegTOb1aveFj4OaMqs0hpiHVQDNJABXpkAxkaDK0tDbZoqV
YQ4eOVbd6Qz41dZ7EVXwRfDR3HkUqrV4wv0z8msL+srYnDZ7S59XZgjgygNiNB+3
fLMYp5LcHPhFOgMdNcM4l36fAAKCooHDovGLEUy4Slt4Yyg8SZYhSrPpG9+7CQIW
L7ApH3nJidbLqpDsEp7AXA9AgqqQvovYZ1QzjP9oe0RZ58U/vQr6xLgcKjHRZrfQ
PY5ElM055WxvXxLh/ajs5VtV3zjqJBZUEMmktBQ1RA50lqK1ATtK6CMeE8EsI40E
zZiFqMtetjO2VWKM60ptQxeLKjBCJXrKlItuyc981ivxZTcuA4Y+o49OVB3+E8yi
q70i7MqYDM6I9OZQT+hZAUdVdNX/U/gmKGflvqioc/zMtrHkusTtJmrN4MEBjflA
hMBrzFDUC/mf0pIAOZwJb1Hv7l1vB4BnaGNuO4LrD2ybA42LqFaRRTCYsEPyh44I
zuzMIAhVDRCj39cRHOlLiDNt2uacdikIDni1tGj6bT97EY6XXwJD6SYprYdrIrdK
C9mH7QqPBAnTLw1MeUZBCDT5gXeMgvyPk203zUma401aFAP4VqQ24tkfzI0i7RRh
3lQwrYedl7ssjl9sKQQcD5yrAtJfQEtZvZVdkBgSjIzWbziqQZKeRrB37mh6afjl
deusZSRJPini8J0PPIblXt0szE8IF1CiqscxxYkAWiTRo/iNqMeMOR4MrMz70oYP
b1LMMP7pKc7x0WGFw2He8ch69kg5CIai6R9zA2uIC4TGAo5feyTE+RVZFp6Egn8R
nqn2RlvKGH+FEgAfXpxPmxRb85lMKOmvSzsmcPfs44sOolA6/S4nv3tVqbmlRQQy
q2iJSliWTalKD0AQKciH86HXPVtq6ug2R6hCivTCReAfoo4Uo6ptQ1fCWTGj1eIU
4KLgg8d+aRf/bkzZePPiPik9URDd9ue2aIPVj70skp87rzqOVaqQL+0kIuQQN0aw
qasdx8n2q+XOmGGD/KhyNpxe+Q3lwEkKhzOYoccmZQs+s7bZcLzujv26k6374aOF
f42NrLV+lWVFoMCTaX16lFiwLq0lHDFDcRCe/t6u61juxKBkqkh2aZQNFqpvlfcp
sqKgu6YGfx7L1NH1zUSu/E8OV11H9WsPK1RSYW60NWrDfK5dKqDeLwuRxb+4jirh
v/EGH3OP9+L57BZGxXFUEI4CVroZ4WaKERSPioXMQ5OugkYQSTYiSVLVyF54/eCt
CTxNqjofXuvXbVNWMYgcRHsNgsJEHQLUDPvLSs3kqzbjdRABd/9Ogvdj3FU4eGJk
MaT7kKggkqDB4o47RGfiaVe/SBYGKN2EHzO5C0RErGJ3p6TCLELESqfx75p77xVf
xiQkl6DHuqg3dAyhFXQPVymyXmKPqZggYFWIbf26k2lMP1lyVyyLrl/LeVC8Pu7r
JAeBEtJo/tg9jaegKoeuM2PMDG5r3jYhBAju8pheQ0LbmUhF0B5fQZ6OUf1VKb4G
fyZVkNbDPVWQC6FSUtwYGnRDbiIuTRZbrpN11cEiE89IJw88pUqpTluR+iycwyba
enal4zxIRe3BTBvhaFFYmBMmCA/3Zeh+Zb1RFcVEOVhI5NUsLe6boWx1cAhf+U37
TsCf0ZjE2ZZ0GNULFfdVXcTlLgnzFE0DHbb3DjoM0DhNiL2aTmaxmEaQiPwHcSZa
RNLscUH6Xy4469zSrvEsUjyYw1DrFMBzn1ELtgyUgicHI1vxiOUhjmMzApxdnPRd
eW6fbHa9udDJjaDMFnG+DojbL9fK0uV30z5SzmbeSeB9cowviTK+M5L6TEcqr1Fa
0NSppUQGYkn+jvu5hJ2BQMU/z2l/7u6xTsrmaQeqvPqjg1YkFCDivC0nCxIzShs6
wkUkMnCYURxNqqSDeByW37PojNaftqivThrYQ4nRZtCl3nEOrRrO2fAhKLLoxEVv
MVMQq0AUVt+P6M797oTHSMxwlECVWr+hvMUBr0N2bEWQcBhw7sL8MwjWipLzEolr
X0fN+fN6t3N/y7v7dhHOyCDx6FrTV9CkJj0b8bdM5J9q8s1g8Igu2I/qj7x8/fPD
GBamYR8IyvUoibu/DjJpPqUKMfOd+s1ipQMFjPTW0lpYZw++Cp4k2I1EYaR1AMGz
AmpewNxw8tUuS2x3K3YaKJ3uNb93trCoSIwHWMNZGlCj/JNbpSavIB95MmlZRcxT
M8NWQYTAyZFIyqVFZaTqxkbLNyef8LTyunp2naxobQ2oSES29VOhKnl+mlCrLRBf
BBcCc4wmJmNnVcJxxVbRtaqCbXr7i3rVnmMLG0kABiV9glyDT/N8+zYqJS2UFhB6
4QU6uzMdfVLQW4GbSdJ039lj/Kq2w/vmAGfo/gKMPbo3edFyZEXNf+CCKkx4iP5n
tsZOf1YuWM+YRvC33AbIw465enDa9W1t/H7yNMmxaibzJe0wS7y4956KsG4Xo9UA
FfIPEKUKpGyPAca7xTG7f/OEiWx1+S1k5hJ61L62uUqBFI9v1d96bNCobjLlc/gy
u1nDKD17eq1P1iVc1M0tBAw7DILQPGwC0WK0B9isazMFkB0DO3UOHusOorljGVgS
HWYpx1zskIWN77TzRX4otWjlKIt0XWkrTH5R5TQtKMhXI3+c4m0xjCOGiB/+2w8a
SjJTdllezcUZgdZBEThzIi2b1QUjMr8eqwt+TADqnaCce5iRWMdQHgmh3CVAWaOO
aFFcyMzlT79ZHRifXlQC3T0H6Iyy9LYCY0PExselsWJZ7+Hnx4tnWNP9tDyluuP1
OyOfraGIVgI4PkXVNr5BakmkUX3wfsZSzImWgOQM2Z99IzeaEnt/omE81YU9ExJd
GZpvewHKb2omw628H1+tIdzLpBeGzTizthJgWDofrtG6e4x0glod2FRkeVTT8+HL
vtffRT2L85UeGhjYaCYxq8y7zb+9JleXxxhoO17qms/mV7x7bopUuQ/5iipOS6+a
NuCgZV3e9CPH+zF9e3Haztc2yY5lRm0b4Bu4iopDWRwJ7l6FI/5Ngn8VNt6AopxS
SYGpu3x6+fQ/r+qpSAXrMdfEUUNxpFZ3agXSvaU3wjAyfZl4N7lHC/kTjBMuiEXg
/JnthtyA3eNx9p8+vlPkFnDiYdMWDBdp9PDILd1my/QAm/Uy2LwOrWA4lavD3a9v
Wb6l0smGEHSN4vuym0qFivxeRvjSa7ZhaUsL69nDfOCp3NsodgbzywQxI1o1eEhm
O3Bkk0Hd4n6WVMRQsx7QMJK1cylAu69WoIbbViSzjgqF9StBc33tcdMTXNzwlK5n
IcMhbFLolLXujmMhf8v1JyfC0eA94OLGgsFvpz5m4vO3xaEROtZvKpRBFhqKwj3v
ju4bnX6Xr1vE56QOEu8XKes+ThAv1emCBbc/fMIxItcZUJr1FDyA1651l99a1eJ+
eBlthI0Oa1U5R05bK9FW+XADYJ8Tzn/vKmfoPlSvmwxooyYe5BqUz0PliArtBZ4t
8iqp1ITgtEayBehG00oGSFh76AiZUAekTcPUHhXXMLoDsKlyRzRauihlnw1UlzJx
QfChBofFIYS//3FUrfbTYS0R4ouIWZxh9hSCx5JVgTlUORCJnrwwSw6aCEvQRdF+
lj6weq5iuR5JgWc6hig34n4nXmi/f6eXDXZvN0Qy8e6TBllvjExa+oouTfHajfBv
5lm0dlhs1OTlYXwb7jmuOPD3xIeFYwfXfoBFhEdTmznNUP9Fu3zEIwymQMRiwPqO
p4qUp4dXqqpzWSM+Vo/aZSwMecRup1Ts0OGBTTctCFefGLH/4afPLdMOtCnMFx7Y
7Viu3odySlng6Ki/xTGcmNtm+EWZQzy224f7zznAxp4Kq3yLImbo1AuonUHmZkxH
9mx0/lgaqZVH7TSOOkqsKOc8uayUe/bPbRcXVwTGVrwuqppfxiqZkAd8ESdBP63S
ca8qpXj7y8Q3olo21rbTYbW5BdRl/XPusriuQwBzj9MS0Dm+yynVVQQkRwf8WHCv
dLj6tGgt4wpSQY0KM071qBajftlKsleLQUnb1qG59fG59fWW9veO//6QxG7mZ0eR
uaDQAgVfhoKm3xDjlVYJO6jKQfsFE2IlNBSdJrtO0GhtL1qPCW1KxXTcXDXvuaHL
zIfL8pxZooiB8UyUq/K9F1+4yV1eB4/2ONJjU8dB3J8XsjqWVQP1cwsnaXRBXWeh
Twn0b133SgswuNmbo1f9A70B9BKKlmo/yN5UTa2zSpLZqyEptAs6QQdspJ+bfwPa
C9N2ilL4MS1gqdb6MbUGWrcaSVPzBUvEHZYAtrrMD4Xk1S6qXaNomRIDpsXEjeGD
o2ZZiMoTUuFH7a5cfKQV1OMGNV38u5TesJuPwT/tiyKD/cUjHlKqpQZow85bkCu+
6YUs+SzBZAno2xZ8D81BCu7/6SfpOEvXZ6tjCBVXicsFh/FsjGUnqzmP3rqoWoaW
9K1mZxfhQRuCZq6cLlLenkpF/0CN6TAu0pLYWpdR42t6l9jjzxyBsY72lu6P5qEp
bwvBO83yQWDOo3sHQZ1atW6SbPWF5ULMmjGDaDETTsE2pHJIRAi9ihaw2DPTu5Hx
jjeG7G9E+pI6W7pL+VI6tNgutmxycnQwTwLAKqKFDW4TIjLhZv9nUJkydqileXjF
GsvWRPD7jhpNNRdsvI3h6CF7HA4yoiSArubeihGKKvPpAED7KMNKWCZXj0/BvlH+
3L8/nd3QgHxXcys2rZaXdRXds9HI0bxePKkjOXYEYmf05NJx/1yIpc+HaQBvBfk6
Ch9jxu4e3zPLTsB0sFtEI/I6IHNT5wOX4Q6lA83hdw7QoTZqAzFE11omMJvo2Jr3
K+Frbq3Hfhx1HFemlGIguCZP1xw5NVyxZtxqjN82c2cgH53IUa7wYdYPF3/s+DJs
5PUeeQqdJfmRoWVcwaj08j36lhxQV+twLFqQlxS5oa9JQ7lS7XguaesCTKF/pJLA
8V8sWUebJKS0msoXlgLwXKbiGZZMM7Ub7LKckvy48PZl+7LczFLZki4MY2u5Ac3T
qGA1QV20+fCT0ptekZlcTIDJhnTtiHHAIBXf0lAodt3B8+M+b1WG+ug3l9OdcD/Q
sjTTRotXBMjg7MNEwqbQj38+Gi+ZfbLcKyUNEaiOB146JMs57CLbae8Kog7LdNbE
Ja04+uUUW7xHteWhXBZ9NhNAiwZy42rzpEnexgDtnf0MFx1+C4aJTQtB+mpIgz9T
8XIGWXsSX/MilUbgA5PBC9QIFMpUFJzOzn3FaMfqS/w44cxrT2JcwMT9R/PYDbfx
XTWkHLiA79er0uiKmqfFRxl8vMgDEasasT8ArrAQzhxuUw4Rx5eGkavUUXh5RsUO
CsgQSmPZqPHK4oLKlhHC0PFQUUdxwlF7p6ovjj5XPxUUJf+568gDOLslXHeWwmGI
f+0lAXihYtuK23GGOW0dXLXfZydLLxSNZocCzE2Pe6sRDdZtnPB8+K1H2tYt4HmH
jYGxNY6wRt/W0i77S5hesLohfDICOIuLAa08WDnEMQTwfq9Nxi+Z/lau0nzBTM0y
MUXt+bwvlnavl9VLzfr7x00CYsA7V/wA1mjRi0sOkRL14+dhYrHbz9STbHBW0Zih
qLHwJ6HeTXZdxypoz1ooMy5j/pJrQeMbTY61FDZB/M1xjeWwurHTQQf7nzOatP3m
gLbw0wxOD4CcZOTHqTaN7Ophshv0Un7pvhZbDZxzDF4a6hDCNzmDHse6otSWX3O0
+P3F8YcBbl83Ix0sq5UyW0cOUuPthDwSGdIeGQfDw1v6LcLQjbqmdD7aLcCqQ1jA
xaFTHyJDutlJkKU+u5jN0KMc+rukgEvBTVm3pG5briluTdl6+qRhQIZ8asw+bSDR
yLtWAOS23yv0598plo76fgbbCwhBaEsCuYtB8fM/YVMy0ephxoaPVcp2zKt8THUS
i37Bl34jpRRT0YUEpNa5K9IC10q0tmur6ptb5ZKK2/FqkOJ3MrIM2CXsz63predh
29G8rYkkFZaDABOkfIKc8lZcLEG/3u75cZo5/gt3AFF/ewB/7J+rp0Nr9h5WhHQN
1njjJl2pJHz4/AJJ6pNUF3UzYs1y07mxSHygPbO1OLCc+7HYNI/1eY3j1OGhIb/7
nkZj8Wtlo1z+Yon0L5+gw6DObzFBL7+56oQP1FIw/wD+LMmQkhjJa8PoVq3QI5PI
wJ8mrBfaXo0gCPxT6UInTq4Frw3nkiUdC1S7X6Qq16OqkvezjiZiwq2eWMPbm/J9
3p9fycY+jFMO2fKI9QwksWEdu1Etm78dktax2n8rOXpCKeUPD4S7amxyoMPm2vye
zs72xeGUzNMmUdehGsZ8qwR7OKKXs+EBy6b9hPDCeYcs0mj5RK7Yz09DaxhaZpQC
7ETsECNQd+mxGJjoUxw8HKo8uzoaqDox48VMjnAWBGlkvxZlMaLbjehgAwuRZaS0
cjywK3FFwVZXqZrAFtQGQusovcf5w6rukLMnghZYNFwkCbr5oKXGluAdNgssHygE
GcADmyJjj00b5C2KyTujA9DOe8HBQTrVz7pR/3LB2pmwhJdA5rK8hVCiUV46VFSI
apkxTf2KN1+6myOtywfj6p1k+OQbMYVrdNC+MRKuCZFNiudFHWSGTHfBXjdbXdrJ
3N/++TFgL1RCup51xKdtno9/Cm4IINb+S5HhiJ6JSxtBP/8TdIeltaP6u6O3EVJV
3fSnWcyZ2q4UYl76/oYrDI8UQPVZ08MjrTKxCp27E8id3F+7usLaLMDB3sI7y0GN
SbgwZ7gDf3SWCYdu6wnxDQhVcJfAT4JY9/D34znAZfLP1yT0ml62T9/fdi2K9jQk
8e8pGe7aTwyqtFxkqjSeqjV+OKUzDYUTGMTbyJM0Wvz/eGYdM78lP/9YuOJGpNB9
xtn0DrWaG/gXu2tlEVGyyMCQ6Zxmedp4L5weghWOSRusIgSzfmI8f/7Fpq/zs90K
vdxqdabjhdohpO7eHTQb3+Qvvj+wRSE2EIXtS8pO/2wkb8rj0wWrhXC1XTEA3KfL
K/sqC2dl1L50rqM4NpSzgeOydW2EFpgt+3WShlh4FicEB1aqsytCrHFYxUnw6wD5
dMm5PC1bJwIJqXs17ujfDrC9+XiFX7BWXTVTQOCeSBlbp+5dwSx7c8Yh9jeMDTnF
2ydivmLyRPYr9uYYcyvJVDsL3pLf0UViT1RAO3Jdqustx6OuDCHfjuCcuTCE3LA9
rDJ8WzyjqLbSJ2QoamY6ufKCHtvsg1uR22QN5kItRJMqTpd6mUlgIRqe8P9Smn/0
hvoiYOZMl5gY72vt4FldiVS9vk9Guf4JMO311xf5vCf6rI+P8WRXTjqTDJnm8k66
MDtml0s8BzsVmfFogwYHC6Aw14M4IC4RhfW9hyvTOzC+8XGVgTN0L/1wUPu5nJRU
Y9Wi+LEZeY3Vodc5bMA05jsYPOOFFO0aywcfN/3c8ZSdVkmHupG/h+mgwW8guIqe
u5uqsFzc4NLyKGQqYmqVl3wSp0s4+xwfh8O5eWIVK4Hw8ASW1vr3ulRfw28kfAXm
3Y3yBNlrtDMWJAZ25etwTSdUYkEh6Y9X2hPqkgaKK1OWBygEQdXkMqmvF78UN+uu
qgKm3G5GJMgtzwFNtAE6Dl9ZILbZ6eYAUxpWDN/gswsPZqv8TPPPlQlr41ofqbHl
XyJ6q2wEKkpC4x4qOyEFnhR5Zan2dbGjeoL+glcbGO526uh1DTYEColU7eNHxwE3
drWxxwq3nS+wrRFgZWwHkD/m7lwh+JNl1S7jYIIrVW134An3XK8dGhYcKeGirWbz
0+FP9mP9GEwa8vR7Yk2yys7wkNaMVGBOMgD4jdH5DzemX2m0hQ3kU5aBiJaydTgH
nT4Gui2UzdNlU+u1o5TgyS+NriJRLidX4pz7LmnwCGVzYu3w7YO5IPfF9pq9FUue
6JBGgamJRPYFL9FtWkoqxKTm9I7WG48Io4pKg2ACpAQcCB3+FsGqAXUizVblsC8e
PVUrMiDGJF3tr7+y0M1HvHuigB6pfqFG+D5RY2bH+/43vgUp/8zjS8YmOGGVzZg9
FI8czzVmB1SzohM6vP5fnZOLZb4FOT825jBKScMPE7g7EVn7nGHaAjQqSEDW+tGe
tWc8Tj8mLgY5OqHzoElgY9D5V4pcCFJNPPtfq3rkR2tGOctzzQi6O0wWndDxr/Ph
j5RaaLPjnKi9E3KNZGKJl3exJ31qhffsQiriaNl9D/KCUGFhSvJTow53QcagK2jc
B8fDRIvNMCZFJPoppvaHKZO0y2gqOCL9VW3pr6qIgBoWIcw+iN8TUTGsOdny7VcL
8DUgpBElgpbsxXT8cLpQo/hNRF5jkL+E8L0xFSsNxZsEaX0B9A9QjVbL6o2KdtS4
9nGXihkTyRbfmkmBR164Mtwtcs0RkiRZnSU4hYpuXuoBIeD9znOtT7WiS2tG6Qr+
pUE/CXyXqtodrKpPfzS6I1qM5W55NueMHXtJuKeOA5ig00O9P5xMUKaoDH0W9otq
aTMX0VRxAGMTpk+z8GU3YaCJMaVOIR4VxiHJ9/6cZ09V76WdESMSFH95tTqtiPyg
RrhIC+R/mySxGARenpYSped3ipwlucKiDBzkZr0CKkHVD8B2h6oF3uNXV3M6ikOn
YcXBUfx4EUDRSyT5i2U8OKzB14SP1ShnFi3+XySXjlXmyJo0fgffUHhesEg2piJE
yCYUGQ0dniJRo1Nclm4gt+/sUWSa4TPylLkKPPzX8i97LAFGtdDnvGOH+zcm110G
l3rSD5K+qJDZmRSwU7iR1UwOS9lTu9L2cYIFTvnir/qgbK6diUcRlYyPL3FHOi+b
xgg2o8jCCoQk7PTpnnLFzdGis3OThs4WWtK+xMHMwauQVWRf63srmHZL7CN0Zl/N
AujWHF0zoUhnU1uFMOt5YUqtyMvO/Dsl8M/V9vzpBy8bp01xNsBnetAbEqL9D0xD
UinOKouPsflKhnIemJB82o8dG70b4faeYjf8ojqk/i0rsVa0/9L3RNCOGVPMb7hh
5BskiD7pCyCwmWOdTkuCEBpTDdNdtrbZyABxQTNY6BVQOpoeN4VyUvXJI0g4QS1k
BwNfEUvjfCY+Dv3KieCIdBIwgepN2FysFmGNVVZ0nNKiSBcq/U25O5Qd+zAT+ZZk
Jnlc2xWI376I0GLRBYj9cTtZ3m85Gzq9WgUpGiJgJSgDrRn1M3vnx+gYF5RUO6Hk
0y95x0GYoFFgT5vjQSaL9DsMWA09FsgsmPmcf2ZjSjZmb0o5j09sR1l+TcGA5W2n
UIgGTTGeugZtt795NKO5lhQQ3cdCXBNr9JvHT5HhEU6y5w6CD0/iXYPMjRRGUNU+
nN/UuPNsbUb9VEETmf19IjL/zlCL5aFGd9Yc2ivkQnqvLWT+L0vtIpw7Got8nejD
zkyLnd0CfZU/YJj2WEPBZ6URVZkOQAlXCJryCMNRdtzyBH/DDy2qHrVwdoOBLuJw
Ymd+repPV5suz4oeExj5u4wDowEJUhmyVEMW4BQ5cST5HCGANmPOZ7MPUcgbtK2r
KEPKxyYS3qxSmYdgEz5gPyAJ/Z2Yy601B9MUe3eRU725HgwFB3ZO0oyPYNOgCkYn
axjmNg/zljTrc7Uo+COVUGw7O9DvqTpeU+QI+CN7W8xbSSZssBuallZUaK6Gkb3L
wEdLm1rONVbfDVs3f64uS2M/8ZT4t0YbOyZ8W1JsBycHeOmz7DJztKpnfXOsDlmF
92eh1kHLB2FR6bvi+4yyrWnfvkzedxzc6SyVJ2HZ1QN8mGloRLdpKCX5OUiUpoiR
f1aE87tc50Oi4rxXG7FQxthRYXqxsGoJGdBkkGmc2v2fmcUQltTM5axph/+C0CYg
ZDbcP5lpI1gjgCd8HDZLhXhZnBvEptyR2BE/Vw2sdx0p5co4Ri0iKq9Qhg1TPQKH
JzMF7esTY6ESawXldHZkTGlXs+BFMonk7SuMPmMMf3qK6zF4+Xyo4fdjFpZo3bFB
lr6UJWbiUOnCaUdLSNIjzVMRc8GnJCwb2TPYfHDe8J2S587dJW2gbMX72Ojm1wPp
8kQ+F+YZZCvf2kz2fNFRTUag01dhT173MdsZLUIxtGIWseNbS5sYj+pf2gsGvEVA
CXc6pYa6pUuO8yv7tekxL31ZXzCHMqUO25kGI+PTWFMCDTEmHPeKp53ClktI31B+
MBZa8euNQwsKnbKauMvKvj3HYiHFojgvHob2ZNO6XUvgCILqSVxRAUHIHDi8qXUP
vxLoIov+/YpWSsjdGsLaK+8cck2Cd9VN+Sz4/Sj9mdyxJpuFqIHlQaZXV+uC1pbo
fZtWgKr7YFeaPFeIW9oeHZRmQER+rWtp9bXNKlbAZys7c4JK6MbWVzUmhRW9IpbB
CxAfSAkrmzNKTxpjyUFOmwO7JmLpOmW4m6vtPV6Ukcwhnl94GBUBLgsLXPGTvBij
sQMErQyhNLvG0Mp2Pxqb8R8B789wLyPM56+1xmefXl4eaIeZlo7JvIxytwcYuR4r
S4ckp7l00rUe+EiSp19zOx/zvsXhAiPNow9NTceNxhaofvm+eUyJya2XD2N3CEFG
2YfGIzvSNW9E0qC6+O+O2m1mH/oqZRrt6iBxSZkB9O6egDvCSf7ENVJ2/x6YvQfM
EIUq8mslGsDVPA4SGMcFpDbnIUE7V50YuqvMSlXnC7Y5+zEPppCVFTHm8L+wH0Xh
Z9fTDrF5WrcLlOT1nH84gryC8yxJ1vN94RyBC4Zn8AXLrJGMx3AJkcsVw2mrx2bP
EFseU/CZ6v1sPvnmJNjJFWi5x2KoasSyALo4kmd1LQuryGShvlEJzIwqNfsBJxev
cN4oxPmPNNAV4o4iT8C5HLaIqxNi/zP3XzFV+qeqRZePJctlMM6mE0SSFiPZ9OkR
JnpJT2e6dOor95UOqrAgXWnE2H+t5QH1Onr48X3AAco0f/bOsgmH8O7yrDAlytfd
9XgrcKwzUl7UQxgiwC0ay3SW88tpOsaiCMEHIrNq2uA74+OGopJzrRZiI51o5ElX
wCAPMAHbVTGtpoPx9W84cBVt3qABwyY0n1q3zWmcJR7FA0zm7ruUy7UEBRWWthnd
joBtpcAhwMvI0kTZTvJpE/tObIqb9Mz0TSy/DrE/Fb/HcSY/Oj1Da7fYmca0CsBG
rNtBdrOm3KaoJI21y5+A7xRZW7Nskz9ikcJh+GF5096OoFiiFnV0VQGKfiDEKxYX
2R9eWvtFOak8bud2VT0t3jIF/K6GPdNrwApywibWYUMs/L7sH710QeHXdD7i6aPI
RtOpS/tTHCWlaNxfYi4wyEc+mWYDSI52wVAETp1MX507LqzAzncaxw+7Td/XiIvt
gWWN3z5YNjwmpi3o/TKqBxqGkTXF6r9CG8I12mDeBjHjLRTReRPF4ZEYNAfhWPdB
T31MgxXT7N70rd9Rx0aurAdxotpjRJpvJ18ZywwuJswy4de/Z+o4Easc87gIO6MS
zN1uFBc5Z4os1sG3XIgI3CMD1Eg+QNw8dFumsrQfDTROETN+Z/wISTinquwirFRc
vt+W0FFM+/fviZTPwT09bp6WAXDeNKEzHQkDqt3NVfZAzT6V3Wc2/NxYzaWXDOEy
mH0bP+b27h8MF13glMZ87h23lsARwXBzuL/SyPPNrJH+1/IGRwpwJBfqJhTK1Ghh
K/GAGYos998Jn2gmrwl2Teaqi3i5gUGIY867+DDgx8ALNnm0MKw/T0DC9DOgcpBl
9ERNLJo5yQs/FMT6UK9UohpJdShqBXmr54v7zpIN5ftXgaaQw29FbWIEq6xQGkAG
16Yrqb18pqe/DbXdduwL+9Ywkb+dp8CHanEwjmDWWqqXSCN3eNvAw1WqhAjVR+7Z
nqf0BIeIRpDzgnNbTRbbgDtL7OYg0PnFTDPKG6hCIo2ifm7wqo+wygFBxmCQyl96
TC1GsZ7xPkeR0WV4999GBDKy0yRR+6s4X/PpGHO4CDvMv4NVp0fSz08K6T3wLcdi
Uj7Ty0N6bCgmitvHma4TjXDEl5cRkTNkISHu58B49LiVp5Nrd3NSf+7RfGSnoWXg
flUM/1HgCobzxUedVSS27AvXhw3+BiiqzcHvAOrbCjuXH8I5HzUYNlr6rWf6O/R3
TI4/zSLG6GEjDg1eNKcaJAQCESQlpNYMUw9W+4/Ul+8leCjubbTpMW5eu4z+CpvE
62blrr0C7mzLvG726OhfRVE1xz3ZESVz4oZnqOMWlzjZg6ZGm2aYZ2wsGVwCto01
1+jBVbOjlZhC3nmJ2nr65D506FesxAlEDnq3hm76cmCi+0bNeM5s5i7bdGmhgpkX
hOjm78fo7dflVUZvJ0/xxcp1qRJrtqzNtQc9o/oJk9NAVmOn5yCGsVBj9i1+rOAT
23XlVw+E3n3zp1x5MZmrT2olJIl8lKxBv0mfNtex+72KeX6M9b1lUCkuj2d0Gth/
sBstWoVrP7VW5Jna4JwNcHkJc02vmlb54uu5A8LVFwwin654R/1vd/fdHqLhK3uL
m8dRKG0/TscKB0LImEd69n8hhFhymy553F0yy0zjeaSnyce2dgFFaVJ2GR0d4xB6
oiCHm45mki1Mg8rzg1yHtAKGZcoyAE1wrmS2XisMZ6qqb8+YI1m4I0MAEmI8/IVp
JCOW3BT29xKFpil8UfO4TAbNFHTVVbWQGjghxX/oHPxXmvs76sHFpRbUgtA+amaC
NfLiz5Y/8vh09OgMkhHzBKUx9tdU54S/afzdc5fKKRodHEI4UDpt8oo/4aOwmbf9
aIuIeC4+ZYq6BniLu+XG7HXcfRkXw0jFWLcaI3jDVPZNFZDKKxtiQxGoNcomX6jk
uMTvSwXtOU2W0ah/ZoxNMA+0w57v7VmvJhCoRh89BO43m4LM2MuF719pqV+mUSre
ke+8qterDXGhL0T7zwFcTlZfnDSaeL0se3fHnSBR1mHYaodMxmRyoA+kc7qMzoSF
Iu9Z8fQC5S09VzJ0JCHrO8kYizNEGHwagCfzw9V5OrE2KcRWTmOA9HPj6jyZGrgH
6XSFQk89UM4hl2AAdyvSkgpmVgzq2aBLYrUBlEQWjMQ7AmTAVHkl927pxyJ08eGB
Idy4cjhr5UHX7hBvzysPSt/6vgA1bsVSq3lUpoUDuMchFMUS7xjrbNvOJ12h6d1t
IvhHwQl4jT1Y+jgMHEP30t7620Fmqu20I1MmCdv0yBNdxfI8BhWL0ueUf+taEn/w
ygTFsg2QxwjdLlOAbQZytQ87tEaKk+mHRJJIuhwQnS2wbJoucqPhMitLMk/15Ocf
RbCVB9NqeP5HxujfEPx68Rk1dnJDnmEoONU6GqHSNyDdR7k9HvSE1ipCAJhxNhys
xPL5ETcs2yf/N5cnP6WRGCyv5foOoHCQo3nSkOhEFyhg1iUyx9lI++DwqkumM7Yi
UAvFnb7QyWtV7PnjkCkEzqhUQeH/mnZJX55ehtg+JCkRRNGN5/K7ArAC0TxsDzXV
+Lp3/pFstCKnJ/hdDsOwDPp768waLuIAcwXEXjr2TOzzxSxQduP9qXsbyQf7NbDP
wmJl828xtEI+LY+BMW7ZIv0mwqVIVTRf3J9V5OEMky9SS3GARfnhu1obLluckvcE
qI/1pEQG233nOSToKEXoVANcVh77aC4z0IoJO2RwR6S/1Iq9hPwpqa8JCsC1J0ex
c1rAABkKnb+XJtI6uVZhNDpMTvVV8yBzVMS63sQ6J3I/S6yf5mR22Ads218LSKLi
fc7WZbUyoJC0nTOLxvbFMcyvDDG5W9IwMW/zDt1aUD+GWWQZM3vQg4FvuH/t69MP
FVwphOZisJbXx3BmjdVhbWB07N5mXbQ0bjVZXGPjEDgVlTaI78Y5vnWNk6I4ZC1m
7tju1YOKYurPhvBUG0BEacD/T8UhZfLZBvyp7W9NF7F0jV9p/90gCHyL1JdeOlzj
X1wp1GgrtHw8hyhNRUVMPszVqrw5P1R2sR0cG9cFmCBr47wKdzfGUsFH+C3KO+zl
wA9kGnseZqFYK6CfoXBfve93Rq562RlDGo7nWcZJQ5bbV6aF7b5/PZfW84WQMBn1
dcgnKVqHGdpPQMXat8xhPLKBGs4HCG455+/MFyltjQ+ivyfcWMN6gyiQxoGfQlE1
+aqk9YxSLBRz+KD3GqNau9altyoKJl+uIAX11Ce6iRicG9tXuCupEnHJw0zY26AU
7BKczzzw+dM7THiQXYl8L1LRIPHtcFPVXndvJ2rcNPRmh/pjQDWBZnAdDK3ZUn5A
tVqEP8uqyy8NB2s3Gq9K1qJEafzec5fdAHpqbQBVoeCSlcaPF+PudwBS1fHIjQsq
eoo/UfJ0dLvvCFC6Yi1/5sh9hyWYMOSfsNWfVB9MKftYgX3uiElIHtwO5JoMdLzR
PlVPr8m2UaCoMtbtdbJMvPu0YDaJ4Jx2fnCQkDGyI791cbCMh7uDF+Y7dsA7HsfE
ghqX6kSgdCRuKutZ3D42r+2hFziN+gV9IA7XTFq1stj3RYC5ejS3ozo7OVOw5qC/
XNRdFdzDQ2V2WkEVxbd2bbO04d1+mL2stERmn/FbjXkEvRmRRHpufZBjO6ubEswx
E30FhBrOm63iftS06Gx2xrJKj3EoLwUEMx0j/P28dx00tjvu2/jiDiCmS7QfWXKq
fYwDPz9VjJpZW9b2w3/Ql9uMyMqL0WWbKboXZwKmUbQm0GW8zqCYKL8KAJW7jRvn
xpKf7ey3yx/HJWVQRhE+N8Ji6b3HukKxJjJjBHwsHJ2EXtYymKF/79c4ZpQMOOxU
4G3MjZfIMS7t4rAOsgm19WSoEPMyfw0h3hxh4W/50sAudGqW9qmlWk1DJSHlOSgr
3HaaVeiFqX6DRH+PFQkVl7lkwqXvLpQhpbZ2U3MRSrOG4rl3fbneQl62R5/fGi4I
c3FKS/u5MAxXg0FLXBJ/sleX45Tmmo5QIHVRk9PFBOPnVEE4Lo5EOkSDZXynW6EX
Q9bAsbPg6p+g9mf/7RTSvysh9N5VxuQWRveJlONklw7QsEY245SSqVh4AWU8xqt3
nA0x2/hCE3kj+R1BiYkH1WovsaPDE+J1X5+gC1Dk7QqOGflEjrIFabT1Cbb0gOTN
i60I4V7ExbuJo/FsUeX94VO93llNIT03FAWQbhltjsaC/sEKymWJOOtWGUNbOyYp
+mFg/PAxMOUUw1MjB1T/w+Y1cxAwcPlNJNAvW6B/psv/h9Sxh5FG3wtUfcadcsEd
CEAk7/MEc5V/yq0SQ2N5wVe3TbwZaer/9+wgcNK3iEdsWNzcs912xkJakwPD6IdA
33uYLVQywJ2BTknlMtfeS0BiDrshTJcAwBLyisB0JVsBGJyJSidDS10Kl1swPdaX
1dw8RcekvfNbbYJ7i3eYbNHQQKWpG4as3pN43bRc/UqeCesruwjQw/TxsnC8QgS/
WsfylT4tCaI/kbsJJ1k5DVpgOcATnGcPH0oN5xXrtj6N8Ab6jKaGbmIB0DHqlrwW
WVE9bgByx1+FT3XJlYYaDXYaU+roNqcKgMNNpZ8sy+vLCOooDPcemjyxoRq1QozU
jL6htwXmLTZEeWFfPomzDgy7OvM5+yjuNOJx2P5U8tDTl447bClNjK2OvPBicWWH
EUt5gXOmBS7XLtg/zCDpIvJaX/1XrQL/TDYS+2j4qod8fKqFnb0GpS5e/lTI1viP
J6m+TIvfIm3Poz6q73fY7IZk4IDe6ZooZsT4K5jfXtZDAvU8Ja/rwCaSy5CKqXVb
BHW5rmE48RRxBAeHA5s6X+/DM7bFHIoN6473Nyw8N3kekIi1V4uNW9D8WlH3Ni4d
GgSIk/Op2OJvoQw3ycz4hwchgMJ6zkIbowA1vTYfvjRGhdGM6CDk53NRygg1zbgV
cBpxWotEodLCtAXc0UoSu5STju+qd0UZwndRajZPi5++g5jGtcWc1QcvlFf5FFGZ
HJXpL7uE6ZpPLxaaUmbgkxM9NxalmxWQXnd7GSPjYDozcX6misVKCAjyMX6AQCe9
/sTU6CWZruDUUMmt7jBePqOSbBlqaS32UG+TbT57stBbnn2fPsJL4AirQD62Kb3l
wO5fUH7y235YyghrhjhYStS0WqqGNoaURaNQFQEGFi7xXSNYVoKpPdW6S1qTfxv7
ANujNxwkyqVQ4eY1MECdB/GzmSweZ6rbDAF8HHLXL0JNIkX5N2IMg1xpEt6fkSrs
2IOkoFECE0O8C9aeHaQRG2SccWDEyBbOXlYK523k1fNEGf+Ka/VqVfHSF3ANhu3L
MOMBYb1Ixn/kqQugIz62G21Lg1eX+Gum1CfIhmOb/xOformRSY2qCLYj+Aue7AT1
6gaQiCD3lsPqbJvQlFrkEpdP4meM0ZEjhhaY4NZkU5zqMqL8f/AkdUhOvWaRFaQ9
8kzzQcR7ueJmjMane4UgJ21VUc/WqEUlXxj6iR2TDzwg/7JltBc5cYBxxNbioHzY
5gprGSirCB9N7MffFPx0FO5TEfsXtNIlR/dZcwaXySJkqTDH9lX4MUJf12LoWLg7
vtNkGQf/IWAdrlg1zJ6T83xJ1SJA6TrYGIcSK8S5M+yHupfuYiAAKbwnbIQoqHoC
601fTUKVAK4ZPS2nBugZwHvlisgfhGr7Ju/pnDEhuilMA25fY9GWKWYTHLIG3sTU
hHsAdLZNY8j+tkKZS7lEP2OOnXd4rhiATR/8Y86z+1k00fulQPnkqcU7D9IOrr5m
CVjYlletxv2w+VTvli+YILe/Jxinzx95u1MVxdXmNZoO23CWKb7OvwC8YnYzR0hH
lDOhEJPUQRSNkkKWPMiBPVunCty1zf6EMMugw38/mUjBHtm+PH3pwRtEr8y2JRgU
UrRU2PVWreJZ5eLHUKlEC7Mvd3DiSU0qEV2ZIdkNb0aBZ/o/DuuXiiisDkVIfHNJ
i9tpNOnFzTLuPhJMKogYjmpfHFegSkN4bcdbd72C2UpH9CFPEEnLQ6uj3hRpumVA
p9tO+BenwjoztW/KtraErAM3xPo5NULXAqN+rXspx3zaUSVDQ2oQ1dSRmSVaizxr
yvNYnS73xbn3QTsH1VgxfeQNHIyR03WwR2B9HV13HpRnvMeBH1tEelO62Y7Gb1aw
GtqyfXnLfGQHSC6frBiExcr5rVpq0tBbOSQIDmP2l6r5ydzsO23Kvc4cDaJp5d9O
zi1X9n8Y3wzINzRE4jdOUBCOWnRnieV2xK2mAOBmPLGV6fv+z+z2i0sve08edwD1
8YCBDrnH1Yn2cS5hvhNzuT/cECRsHpm+wGgh4j8iqU0nfJe9bD9jX2GLotlp/Gyn
YH3o3x3CKJE9jsoqUFoT5GqnM/3QRs6p7AqpqkxOrx9dzIFMDYkgNk6P9ub24pZG
KCT1CHAM+k8qFQ3L3ALx+Ms0bLaWHaBwWJJovL2yrPTbKsOSAad7KAwG+d8IlFBX
eWf8wqckAl2l8hjV/TUYIBsBf9swHRI5JlyHFDLexxsyzcjeD+ubwzaXn435x2IT
mBwHc6Czw8iuXC3s8xxAzkz8R5KOh69euLdB1V4icoz+/emPgQgUTrXyZjCLQU/e
04tBpz+YxbHmiKKWLf7z+bF5eKTQdFy7l4/vZMuUTHnMxGVJ2GbpqH9dgr0QTdVe
tgm83jCP+HlLlqkB+4bdnvs+FqRD+W1xkWC1ng+PBUwTW9OqwGe42BC121DrHbkL
j7K1wHHn6VMPmU6l8IL5tWOduy90uNxu6JwZNPB9zSYEcsrFb2xLPulwqM3SyxD4
cZFSAJX5FJ5WtqRXR4JQITFv/1WjlaKvDP1fAiL7fjwQ2W5IIHdt4quStTE7uTB/
MK68wnh4xTuxQMq+DCIHU9n9lmXaWRcq+1NvAbqlH3Xvm22i/wQBtpJwNg3wlRQI
GJ0uOvIXceciPDZ0sKJ5raXcxKd30kB9KOl/grY5pSqYfuJtwZhJ6t7PY1kVMRDM
vZTk7TXgugdhabzKRsnphQEzR7y9/y3XYTG2MGmaCGApq2XoUda9GFrboQNO5Nqt
ImLnHnntGQutexTkUeTKYo9NFRRERq6u8G0T8DXmNwaqTdPd5xjhIZPpA0gfTxKI
J++DHs8alH0GUCmhAQiiw8UXltd1tHPfqSIG1fES670j/kZ+MlCQwAx6VXpcYgou
thkV277YP6igMQ2AsfJr0etau2t+PLG/NrmVUIjCur/rx9T91A0b65/Iblx5ykuA
j8A4mOJm5LPVdbOmy4KqBBOOqb6tAIEKcbKIntKDJ6FP868VAGt5HVN1gL33bmNX
W1I9sb5+XlPINITF9fufuqmCYzLYsqTkrHfLKnAkPm77uG1yrSzxzDrF9Yl748fB
Mpe+OT59RoJMWaeKkSjW3tJ4cIVU6CAhs9uxQeKgrHdb8SiP6ovCQbMRZA/7iTAH
NVk8eadmY+CY64Ef+y1bKqQaBEE7DI1LZQev61bpfReScLaJ7UshsXfabxBfAdDx
k3C06WohyEi/go1yS3uq4IIKthF6e+7Gp/dpzo22oSSxZVY1LVS+TjE8VnhYOKxG
8rg2WiWwYHNQu983FQuaTHr0tpK01Yq4Rd3i1QKsbyJnZ1qtnpSInc/diOmNVceH
E4YY9IbOXH8l3XwAogX+CpNxwcaNJrYPQltGcaqQawxQwcwy8ZDNkeWYJbWp6M1O
Vpq1YTY1rB21oC4B0kYsn9wQK0SPG07GH+KcCAHthVlgp1u1XjWumr+GDvFGpJDV
UDeXFC03tfpDzfd+C7VY0q5TFGWUL3JWUO389jb9Ewtghq2c+Vlfxv6evBgfVVA8
f4SSs6T90kbLbLYU9xlFpsQ5ETZWOZnF7RwFnEtqbvOJUKCNRHcY/uf4dCA8kVvz
pSuZQDn8hDRubBnZPAUgohN2Z8y4Rx/VVmXZbjveJKICFcIljPLaPD6cXsX81JdZ
gDSlpoCwikY0UDha3j2mOIDTpLUhytSQNfqVHNkytA/7Tf9AD5z08CbHl7FxjyHn
cb/4Dxc/bh27N6sLPXcyaiWRvNy+9TuCwBznEwiPyDkseL35f6cIal4AJzzZwA5z
JPugSZ0CUTStFM3caWbU9lgOf0AXwoY7jmuwGNJ2Szrm9J7irUDpHlOq8bngbnbb
7Sxo767hzd4fquvDUZ55iTGlXhkZNjKWpytKJjmb3L5/Sgm6PrPuhdAzxmrInqLD
rItNjUGDxXnLF2KLjQmqq5lVKWTqLK8vqHbK3nGNulTv2iiUKYXfs4QRTgpJX5O0
IbgRyVKzgKnoiOy6a9qgjGSaaaSnesk5Ed/S03w7+R5uRoAaajiBrNkO1r+pcb5H
3cILKCVjI3UZMANjqSwmgliavMZNpOp0el7/krHGDxtrLetgaoEXYJpqyBg23UUj
cwW0UcFKfmIc+73/I7JjST/PcCIL+kebocQBWd9NQ7ZFbmU1nzQHtDsKfAVvI5US
8NJwC4WXTKzhdcpNA3/x4wpw4INelLd/mtZny7jMyiMx37kQ8I1jjqf00CVz+xEb
Ly0C6X8+JeAdANFzvJ3nSypDp9nCxM7W281Sutdkglt2x0Ulf+E2k6xJuh2XSApk
mKRfVYbsD6Z+jH5hgvtnhuuFgRmTCmXQxtKkZOqO9e+kG/Vnf1j6qVFqaHViaccl
YexOSHY69NHuNNyrN2NYGG0nChbHhbDmmAN5minaeRqwPAb+zuw88KKAvxLV0WWp
SWB06j0NB/2MUJdfBe+4QSvAatNxg+eHm1NBUW+TySmjgBNlY9vwh1mMpdUO4zFI
9ZYQvba/0i5p5FSFpRpggQXYKeVVurIYLkF4xrYMwVFcXv/XR1QQcqMIm4cH0N9Y
B7AFwTsUweiKaqV4oPIVTwG4qkNBs4qsBhRWRJeLzHkDOe4Rqx61vJXMDzbgMmp5
q5Ojs96XNY5BXN5YFyaYTj3TC3z9y1pOqFzoEE93L/Jr8oVk+/Hd1AzrHxlm+rjD
f+GUPes9OMihjA/4CQoEuQ==
`protect END_PROTECTED
