`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40RRlykKSi7DlI/IdCiDLEtX9I7s6Z4uu8F7l2zuz6ZQ
dMUkbvSc6c9xhbI/0qQ9j9HcDaJbIPrBu0fm5ZHQGQCylssDElicLQhchltPjZ0a
CYbBLI+gcI363RBOp7qNh+BKc2iDc5BRJrqiYsMikr4HuV6QboviGt0TnCerNxEW
GxJzH8iRBvkOo/NKmeh9u6ENzhI9sHPdxdFoLW4B/qofWxNKmWVKJGKZ4zyQ+BG7
wPfWIZXvO1Bx21bMQhidYaHmyZLXBvEbVHRrMf3GRUrXtx7bvrbE6V1EtnyEAJA7
uMCDll6UP3SREmLYtWJdDw==
`protect END_PROTECTED
