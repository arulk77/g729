`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46oH39pqrF42ueXJI9YO5Mdei4HXdQciR1OaYFK//11G
kSshAMaK9KdDijeAgpZorbQh10BPFyWUNHwzKHdFn3MP8gcOm1ABdeSC1uW+hsXq
QDAqe66p4soyJU+leUx9t1iLOTIsq04Z5OFXWPfFAAWG9yJcyc3zFgagz3tjXni9
cJSKIdsHPHJSRyT2Mwix5VU2uA9Lar7YQ1QPsxAo0/rFLc/pUEDdSEhnxL7o+xz2
9C5CmrO+5Nd9Hk5+cJKxuC0uf3/z1X6dtRGQWRkI/gc=
`protect END_PROTECTED
