`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN3HDoNCD8TvgdBGwaCeAwJPnqTfA+Bc+Uh1Y+91SGIBj
oa0UcbkLs3NbE2etC0KxATPKqgHk7kxrAP6fbjRbWwU3OZZlG88cyP+dCoZMMhH6
ErMAGppZSLwHG6X0rPPbwm4vEHPPkF1VGk3gNAe6PM/pEhfql0Uc38HCn7D8M8Md
oBoPzf2YC/LTt7w4nWmPCsP7MnJD58Z9CTJowUxaoEs5Pi+iw1ubYIHcukkiuQjS
erf6gSTR9udSfcMlZuGzW+NJ+qE2jodOvgIx9Syf6gPeFuS3EKWJEG38SQJh4Bfa
a382Jx6B681CefW0qVOUJYSFEJ3PTi0QObESGfOIOgcRQqfshyJUyVlTbVlNFyJ3
DlBVQJveCO5dY1WoQ3AGiXrFcLk3XOfwuvP8cyTouiMjazK3kn5/eNn55RSdnlMu
dRsqcTg9Ab5YVI1jBKmsGLXdsdOKKQ3tjEitPyI9DPo1t+Ak4GKE+tfaDgWXIghM
H6aWYr6TPIiZvvLeEM9CepOgSKCCqrM3YNveWHgXxgnU0szTuGpOQanTs5UuSk8D
Bhhi/QejQlx/uUJXKlEKv0Hud2EMBONjTkoWrezMk9NV/Q4m9oqxdCnDhWA+aKNa
cLSi6wNNv1F9PCaKTM5D0wcAvI7FaDO4hrtv3PLNJYq5IjGs2B9eUadnQa/sxbiW
dTfApCrJXLAQWm68HAa+5JEqbBgxs8jMses+KvTMdR7uBtL9cbc2lA+uFcJPIiHy
qywO5nxFeMGjcFRmj4mHMr737p2WUuW5zeSfFcZNWASmEW1tPs6hi27X7rE015Wz
eEmo8DlYlzAKlITVvA2hqMkxjyiau4PeNnE769SJ1CLGIN/IMP9pm4iM+/OP7OFh
iuC4CS/YcyjPMPq4lTShcOgOr7siezzwqtewWqaxu1DwQxXJRcFdTvt7TsZ8VBto
eJwAL0Hd3N91Sx7z3vfiLpKUxm2VAnA9QA/tlFDf5lSNo3BJTVo2bWjHuV3KXcDc
TjBcpGUQM8qO7Z3k+nBInnnErkKacFAkp8RcJ74laDCYEoHlEcvVf9WF/0gvd85f
cBfjRxAsJC9QOTEOL3FOeUq27jqJbLhDxQE45UTw6g5G5qQMlTBjAHcXLOjYWPLR
iVeS8P+n/vkWIIMHhF6ZMXdJtSUrvE+KCYR1kFDY2nxppFmU6S0ZAlOm7UUZrLcQ
yh+sgOrdPe2RGiHtzkfEmHZLzQ28yFZZQZx8X1O5sdnF/bJ+E/w8dbQztSXSZwnt
9jBbAU3bIm7W+HMg+THTzsNEEQnUkTvHYANh0rbqwLUD2C5aV6u4mU5hTVmKppK5
I3psb/RCQWGPecCEtj7vet5ntUS13ds/obsOwAwuOox/zWP7Fpxnd6mExpKnK2XZ
xQLkmsIeXzYR9OOrenQGBWSNfGZ+9IiFkl78l0RRRu3N9tkElu25f2A/ZoxgvIRk
2eaGfox/J3Jl8LG6JyE81Z8z4a+D1XmTwwI6EGA7jo5+NiijKt4Rb89v6mw8fip2
GBpwy3cVt2L7MDKQouNkze+EVKIv8bZixG8POCrdrkIoSgcTuw22eF6FoIi8T6qu
RcNScHM2rIZVVV1shOf2rL4TG/0V4sB0EVcVkmN6XgAcblyi1M6rk2f6QdvXId4C
3qOHECJYY9jI33AL/jB9pNbEyv0LiN5A245hWw/H6IJbhNXUYN7JR+3mNHkuGNa8
SrdPWvnSmMCvPBuSBImqpy6R1nbQ6R5ZLdafVpRZKwT4yxV2lH2aOqqXfvhqIh0Z
aiCbDA5n4bQ4myZThiT3jGI9VsctnVO9SNqLJgAcF+qcoKVjJXom77ElBirzFml9
ALK+euOhze1Uo8cCMRc4gDNOme7O4837/tAeRxtUOnvdkhDf/XJqC0f6dDiJa7Ye
hhV2LNnckBGUOmKVpgOD19k+UuTx16NAxBp24bVZqynVhDt96XYOFA4dOlRBhPQu
9dRIxiPYGW7s8c3TGkF2k7aJFBEsDuqJWc6FRIW+0MBIDZNsWVYQVkXiBjVEcSXU
2HlSxtXEbQ8yoBWGVJDYTvofRFtMdVd7eyrSXvBCHvPYNzh5rJtjZaN2LFeVzDDH
ETrZuEQFg/L9rbO3135u/0UGkXeEkibp63qPpggiKEIUFao/BAizMycGlzuXEiyK
ouij8jqNDt5S8fzxAs6wM+cF0W8js6ZPjXrPS0PN8gcuQTzqU9uO7JxYqOAAAziy
Rtctty3sgQFs7zXCLk389lqMN8WkKW8GKyPIYTE0AeQ5/J7mCGqOGc66cPZh23st
nNF/CDBq7pFordlMwsww3AvHsLAhkT/08bIJTGT0J0OcQAOrLYeAOmASDXCIIyRc
Xk7zVVDyaxKr+ifr5eg1m1bGht/MvVR8aaxSnvfihnXqHNPuR4VPzOyAdDWhWICm
WJBxJQkY2RHHTA4BS4I8ezEdB2XAMD7Vm5VsVkDaxMuxszZ0bSRpMdTjSPJhclqX
mvVUTQbZJodc5c11a6j2E5virzoPu5PstVW1DN7c3ff/WOfNZd6NoTfH+d/bw7BF
/PRhKRCAk5OZsSCIDbGsUObrNfPOtIym+9qVrIH0EuMXC+BPiN3xPUT/0bIaYR/J
IkHIBtEBHI8J9A1SgEHzh0oOSycqvsyg0m4PMZKE+heZcf2UBPLM8EhBDwk8beAn
MTuZWhds5yG6a0RxjkFHx1HzujrgWAMg++rHFCHhqpzAPr5Q5GwBCn0uB6yDhwz9
kH+BeOVqlpceGzLUv/WivlQ3btMV112TSctBp1+l+TeeVZhMtRkz8UcyQ5j7kveT
iDyzeE1AGc4YFGNsFAR++885+Xs8nZZ3KT/na9oj0MmWb91pyWdf2VibB46p0rGR
M9xgtvHmECEUK7JvTqHvY1XLsTKjK5r5VpfSALjXc/cTLoxaqYNRPQMI4ilUoqNj
6bm9N4xL1o1kgA2rMqpBY6WWcylJZGMHSG/A0WHn39Rny0IrMqI3DWgDEvLxDGtB
WV0Y9oKTo5SaQiJH1em2++3Nguxu3sMAf0vHoDI4Z+UVpNfvqDmJqwaerKeHsCbQ
m4nTbHIfFbEi/0iiSUsMN3pSWPLR+e2OD4Zmjj9mvSJgSaz6cGLXFEIbNnGI2ebO
qzw/5fqPhDgQHXt9QApCZBx9OZ35ku1BSRvsmoMkGSUvgfmZQ6Xz5fMMSoglW4O+
0gykyAqUMTwy/KxCgTy5EoGFl85vMsjxQxkH/GQLkaa6tRdOJ2BrqmoS6P2/XQE0
6JjFBLYXu+TbLvG3JElxhlac1ut+jZiHsI3HsAeFhmH5SKe3qlOF9wUP306L/Hh6
PFZutwI9K9jNgiRyeSBjkpdOXOufVTu3UHLN7k9A3IIMRyuHGIqPRtYqqjBtfogP
IHowYiXlo70B+HGngqFkE+WoyB77gxQQoWQlOtcLSXfHytAK/L4QyrJloietwEzF
nSCQuqZSV5eBEcVWRlrb9/MYP706cErLmRiqS2x7gbAVtd/YgerxzsrDrnc0FzjB
aSG6vfETMT+9rhjmEKE0h/tSCUu3fGaUK+hgsZZ+4cz+002gjeqXfQi3gNJRdZmh
mcVPN3CVJQU4HCeRkTvewh7Yw+M4W1sW1YDDZWc06IwIJ8xBAvyitQuDTas2+C8+
s2JfP0bNV4jn0eqmAgn74AnU2Iux+h3XcWyori1G4/I5vg0TEoveWs0tCx6VfifJ
pMTD7XX+ogjTCiavFOuEp613bUBIS6v7/Drr3qCeNjkCxTeE/8eEoN0bM+2EkZED
ymV8VBRdiDMS0b6/RN1vtJzLoyUl+VOnwt0gVJRt7kRGTiO/ZM8hvdjnF3TWLEwR
+dgLl9Ne2RX0KiBHSSCB+yncT9nxvCNesiVEVg8tSvZ9578ie9dFkSJAJkjarP7i
KirvqCk7m4lTZlSgW4iwmIixQJmt7ic022j4V3+WBmipyM+RFPJNvoekpL2/WvS9
Exb3raWRAVQVQgAsvqm+NGhBxwVhZ8WTs6g7ICwq46zz0CuWVSKZWSMZF9q/p2Hj
2YknT/4V1FJ2Uq4Mgg3YteEQ+bhXhMKegXXVM04FjeFopuA5ktvTGakYcwBOIp8M
Dm6BIDadg/88CJF6Nepau9Ddhv2oJm7+DXJCjcrF0yQ4dv3qRUwNh4DEZx3prQ03
Ph+xmYGn9U3LrXH3nDD9EyExZXxJeuaWXISPhggSyrcs2C2kYAtDh5RuONafDU0K
d6qP/Whs3KnFn6MSHN6f8P9jP7EHBSTd5LYNnq6rMzD+AWHNnPIuuwx74gvEvsgh
C78y/2bL7DDB6GzqlYWJ9EU512t0UzGsuwbkEGZzvRLW5bzFRLjU5nPWdJJVHzaY
A8HA2sQkV98UfxWe64zBhM0m4itUXpeVBj9tZqXayfVfVt+77BaT4dM3gYPBIzRV
QBI+u/W9MIjWO20KK02f7cM/nyazY7jZgNYPzXg18Xm85SJV4UGxj2k7vuoIDWE3
ScExOFIKXT1lGBwCF5eCs4uQvGmLShXnhsJ7UeUGdGCphbyeP7BnBz7UkBGXYCdg
Ly+h/ANo1qm9j8Uza3ZNy/sgfaiV7Kzd8O6cbNlXJWntZOuaCYBM/up6rgJRaQ9P
bcb+E5Do0FQZyYrH9v2qHFZdm1NiDBATyIwxZYmNxzy9olRaZO1oxt3/ng4R3zWM
uPL0isrsKr92wsjtbAEdFG08x+LsYPvQq94BskrYm4MYYQ23rEad88za0oAhX349
5/tN+RxTauzqNf0i+deSkGmXCkOl4m5CNgTWpGKCu0V2Iea1WuJ9ZbfxFAjnAgkF
FZ0kWFPpIaxjV5E7UEjlckZ0UdKG/FR1FYvXAtJqCRGYeKFzj0PqwxbWGXRElpHr
QfMFLDQJmBwVLlcX/zd2tpskN8b1FuMIvz3ZKNFOLVB6OaolwhzFrJrQq42fbqLP
5Np4i5bXK3FkboidqCB9Cj+Tch0oru0RIKAP41YJZZ4Qs2dsW4HNjy7ZGb3iemRa
m9aMXa/t7tLef8s1ePQV30PqClaLKRS+joMuX0VrPTjx1cMYRcn8MRgmbXx1eS7r
MKHN4ZTczJby5z0gt/llIlZkziz9TPvfWsItkdvhUm1YLdKY9vvhleoJkc62dYI/
tjEuqXks4WzQs4wrib2yfAkcyawnFxI1DXhzDhhZM0EEvNMu04/gR45JAYG+Iw4O
oCwN6Wv+wK69wlMtWV6MSVd9lmcs/2cL0drwevvIDFxb+DtSGZyBeSzFMMluCl9G
JUskTtE/uzJTHEGBom/DYLMFA1MlU5kwgdxANhs8z6Ik41cXSrbFC4goaNSH5ELf
1SOBtRr+gvSG/TGVoTyCUZMaeQXnylONf/kTChjzKfVV2kGw2teoil5uNxlgmt0+
Mq6V1Lwy653u81ET+NwJ210pXZLunhT93Y8iVVoUoPjGt8Hh4cQ2DjYTlxW8w7pJ
77sro6l/IcPi2ePqWrN2hhS4gUrvkHD948wFtFIvIdTJUe9o03da0fc6m9hP5Kj9
xu4LmW6DE+S7Ug4gbLt8zElVHOJw/NYwYbUfRTk+MIjKy7XLBqKsHUbgL2w7Ug6K
xq3OZQZLfP8CXtwASk9GeyU7CvrgjvwUj8kl3PLsP7OvsMvQsixqDnpyoMZK51nU
pXD5wVhv1uSy5HusFO31HE4mJclbVM8Mky+ZG+9Q2sB/6iMFIiBhfVENzL1PtnNT
+FPUPLIHUAX7h0DWP8nvIBROKWS2I68cqdrs7lVsQrFQX48ijll6rnEkSCPLFncL
vkcEobuH9/J8MSPM6PGztl7+0OkkqBVp4pro91u0CoV96ksqUnRNNFLaJe8EHcrz
t6tjQZ4j2ShStH4ytK8AURiFBgD688XLXUv30YZ+b5+/H8vZA3Z4mQgViUIDQI9G
QUlmXelv68EfcggFhgF/8h+TMyARjm1iEuRW697CabqGLa2KnS/qMgoDUVJTBS+a
0ah/yjSMLcOPYx4EDYMyiWGtZDIv3kPTCYoWipRRM/IKhubgtmFejxGk9ktIk0sm
CcfZelvtSiNuiM6gyQo1WI6x7rlTXyummsYbb9AAwSya5z3mrDyppAbmrwmcCSFx
GD7q1eihBaMYTyOyCiQ4478+xWNlnOAKg4qy1/10XPk/iSfrZLRAyVVOsQ5smmx+
deNTi8IQqSJ5a3cANRx0Qx1s/C/YOeC/ZSw3RBmbhcvojRbbF26fUdr0YUi5CYNs
iF5PF7HpKERwzxI9feSubHwWc5x5vZ2gASdLfUHT5InN7pu9/Nb/qYmz9xu4/hw8
W0S0CgLslunXDuxpa2M1WWEZ8swJLNynAXO1jWJpWxl+0OYWaKTvKa7YNLU+H8jJ
XCdBcANgvnQqvC1Q5vIe4wMUYiLYmBGvEf7jBvjhISx+v/KN0yy0L+IRN3T8JskY
IOieCjBn1Yl6P34kkhz+D/nX9XkwO92fAVcg36pJkJBwSbpuWnlHsdGq1jLd7w8m
a+kaRC+j0FO+z0wtIwltUOQ+os8zVAt2ZvquG7uTxV9z2o3OosVbAZMglXEhSPYb
UU2CHNQOGqNiRjJm/GVKQeXBjx/vbbvljI6QRu2qW1/2//Xuiu0ycKzO7lskfwFx
y2ZHPV5UihCBMZpPytcFVe4H63wZN86K6KYPtaYVoOLGGAGedkzt5HYTvgSXvI3c
rvDI6wyZc5EsSoT9jttXBjKTtGXZYnkNkZAoWh7Nlt7zUcxSvFezo6U1qlbyzYdu
cE3survRCJEh1t4M3veYQzoDQ/jKsx3dfrPUFe7zC1O2n693MKhmdTaJR7IzXQjv
PgDmZVQ4/qyM5eUC1eEusV1SdYGa22Ch6y3LadYrbGx4pjQGTDz2TvSM3CPh3Yf2
rV3LVM0h5mC0eS7mAbhSfnPlfFd9fjHtGpFjXsIAjy7Hw3oYrLQlmkNgGCIXJvil
Yn582RHYAoVl1h0JgNOw1397jjkYu0PfEBlFCYVgbHSe1gcRxcNaA0ypNKsnUbxn
t35CXcq8XC3ovy7l3Jyuk0rAioY9bdg7X2JZi/DnUyDEapmKji+veA+Vib3bfbcd
y7JIc0fRJDPLk2lgU9KdQjZ74kJCteStqRQrH3ZPynT7NC/VI5/fOYU8sGU2wx52
TUrV6UDpPDmhgjbImI1H2sr6u1hsTpa27Q+RX6/8AxZaShFjsCyOMbOwvireMrMM
GFffuHadq+6IFi4ZIKAuyJaFdfnbgpJWy/lKX7XvMD4rM10vQKaTpmF3mrMadKlm
Sx4a10L9ztqGfM23E/wVWuB4OPWqF12ZzbuhQ/4bTEynUnpR19QMF+/d6JVlRRnA
/2eXgc8UTuGvzcI877ISMeJPifwXSb3dreAB1hn32a1D2MoVP72rMDLPOKZvi2YE
g1Ndk+ZxpcJVI87uOa57wcIEROjICD1DE6PD4wWdtrrY6s66JBF+PxmrGPFELa8g
yQgaKmVCC31kzF/zRKplzz68gXMi2MWXkmuyO2OdQdtbAgtiNIFWGBX8RwU4ieKS
KfatUVX0/htafxB/k+1YgHfBejt4QrTBWM4/fMIIAXLmBkM+u1xIU7AYkgsOJHTF
nPlNbaKRAMj965PSgIAFZru0ViyJKwfN9u4sCQ+O/y9KxAIcdS1noO8QsIz7xC3l
hggcZb9rWCvUq9GIVNQAPz8cBYVreAV5EWhFJVUAil3ik4t4Ez0ZwWdV26/uPYxq
x0jq56ii3wCqQ8AhkQ0mNtclPe6+qo3eqXCIoyYJAaSy3AonVcSczIn/5xna0m49
rIytk4+zxaqect1oBd8uB048KP6GGHdmqS4uz4uDmvNFWgkIWTkJJC69ltmage3Y
yOdpQKRo8GW1+UycnEToFERaQJ9z0PdpUdT4ORz+tCtrAFY+kJkycAAa5mURRYJ0
TnQ08udGVHncU1IlOSBsuC5zGsx89yjY9zSicGMXD5iSmrUqBMbaebxcOmhsBOOw
CwO3ncrG7PBWpYauZ4V9zhs38kisv7188Nkl49Mid9QxOOWUD/RPRFUy9HI4OS/c
4dNB5CoDTZB4cfLjsuzgsZDRqsmksIMhjjOzm2AwtyKJw+URMapk2w5NAIVaPF9t
uiFnPVAUIA+fdeKx5y4N9cnHAuOOU9vJ7zh3+rpCCPDjtpLd6g7pSfUDyFjmTUkf
Etb+NiFpnSxH9ufHMi/bUvTNPw5LpcqfAAfFc//TIRos3qt5z+n4W8mqrdLlzkcc
VtwwKmjr0RrQGxaD14w6NLEkrcoNY0Q/1r/zGqK8KtAczVP/QPrnvB7OVdVV9m0t
hv2a1Rw/jTpP3fvO6JPxZVk2QCHVgrJS1Zy5mUO1K/TpFvnhI/WDSQj88IT+WGXp
G/le8YVZjj/7b2ETWY5UHBlwL0YlPkZJ8elanCkos2NyD1O2QprNmkorlLD0m7Ox
/cOZyXJfgXVgzZsDXSuyMw==
`protect END_PROTECTED
