`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C99foBPJv91+sdTxu189R3a4GxbX1ysmww+TP0yl84cw
Jep5Z7qFVcxjNV+DN1RhySsBgk/+oAUrAwN8V9f90pG1cZBzAsilSjdg3WRfHP0u
9q0Np/Nsw8kBJzOV08GWqHTL3owg7DGpZmLQ4VEjJ08OkRbKLv4inp/E3aSxI5hS
oAiQSckt2W5kstp9rbMcO+vIYYzXHKgtyzuIGot5NiIrGUdhOVszMPqcKcloFImO
Jv8YRRKhMLvTLO5r2FhvSoS0T5nrNArhbZrHAeJS0ssl1JWi+19Y9t3h9BD5S3IE
ad2oUqChP7b3IT1dxEa2ZegcWIHz3fDT7BSL8UGYB/awnf5x1Ys9yeu93va9KOOx
kL8IYHFv7ohSh/2k/KHyaJ+nmBA7Zt8NlkabMOWZHgeJFKq38zgbb+eEdaux5GKb
JJOtfSQV2+14mDLf2JUKNJWLzAWSdqEXXbxwuSTkcHhQz9EOkIkl2kjqX4yBx0Zs
jwykmzYm52kia89UK2ELJ8g45OhzjPVsihU8DuTaBqurJDc0+ZPwpavpMfde0pnS
aC72M1V5Z6JFD7A2cRQBqEkcnrzH7Uzu5V69EIW3iD+eyAqCKWibby57kolFrpWf
v2PjGQyFRZEERuqZt+qRo5RUellVY1rlpFuaJXMSxP/sVFyLA1oKyT/DHcVq5nyT
uf4m04p8LSkYwVMYMVabVwJRERWts+wUKAPJBZKQFtSOz0I1HkVEbyTCMXf6XSUr
s2cu+EG9/vYUKaVknawzu4q3Q2e/LNQgUlRnmbV8s8k2h14muI5TSe6tWYiGwlB5
qpjHY6fzGmwTvlrM+IK5oowx9Ql7Qnva7bFyewySJiajBJ+QJtEmmV8IEiSREPu7
9OxEGpm3GyJN65dQbG5HEBdWT7W/bUXfyf47FGwLy7SLUoSIdc45zNaoDYMFMWiD
Fc921a/HnxSRK18OB9UZp2KrHSWcJA54MjKoZ8erL+adKiHRabp5rk189P1Ojht7
ZFxCB+CcCjrTqeK0uCQD9tPgCpl9aJNM2XXT0Td0Qag06cVRdIqIwblULB0Yob53
V1GktlVC8Rh7l/jem9rE+sAWt+UccBXSvzjzWZB4o4dxJI78lOcGVpBD1fpJ1nkD
m7qykmKk/eOqjUFUgyHkRapOW3HtpkMLF9k+/vbxMhMkDCVwg+4dp4uMmMFGWnUg
POkxqoxYgDxsgRYqTN4asWmtJUOcBAsoiad0qMjEhlg8+OIhCVg83NZUQVpTTa9L
ldkVSf881z35QUkecRGjVjDNe8G3MTq4ddK2a9L48AjVmoVLp7Azc7Oeyod/YEJa
mw2AW61s4J50TGS0sZgXkIzeWhJIlRmxKAomQWr056v/dtmteVL7h02BjShU53Nm
8OSeWz4AUg2sgaLvKaknOqtf5G8YIM7N+e3jJofDLtolFinnu2b7QdcJDC9B2yvf
kriqHAVEnKv3psG506FRyqy4yHGs6nm+ZEY7gwHllIA/eRSDYocE/j905F7lerFr
YVBfq1rm2iq6oNA1l86SnuzEAE3t2VfQa/FDnfPA/ewpjrUjVvTs1sLKtPxUdSsP
jtJ1kc63OlnJOG815l8Uf5qHMUggdaEseURSjxwAqFHpdFBBmJ02BHw/7Ilwq9u3
Ha1ImSqG0L7juN6qBM3an0vBj7CZyHaVGmEWTCQMrtEhR1jEpleqKrxAIHrQwwbd
agvNJt+e0Dit6RTEsDv1PI0byjUapkt145mztZXTExdNLlHbabT3Y3sVpwIEImP/
8A5yLqYdZuhUOxgAOXQhQQbQYMhqsydx9Kw3fh76YTlKRpUWCJDMHcEU0HieiSFq
XDGETpX/VNH/ahlNvos18f3LnxxrwXutv70XehHouB7G4oD8UyrTZpsXNPSLnPnw
+5JdZ9hZ3NWA36pZZDf/9xxGyC9xZLqxK8NDrVRuErdodt6Ib9NexN3gF18P7HWl
8k+kYF2fBsrl7shPi9FSznvK4AbkyaTSgw80M8OILQCzmlUmmqvf+IPT5Lu23kHk
zB9Si527Y6u6tzUO8uDQF1mBEg60jHZEtlBvnyO+woR/Vfa4w2wPlegv8meOd8Dg
XqtktzpykQugZxZRaR6nkB0AauIQCnhhq9IEu6gvzgnesYfuhSFzQW27avcBRHxK
EH+UAuQxxos3N76Xa/6hnJtLf4+HSbuk/iXmiX5FlwQJNrc5dRySyiMHk9fos/XU
GtwKo4f3VAJ/0Vxro57aQX+xAO5A4w7eKaxuDppkNNLkUTt5keVjOnC6mcaFPv7O
90jwlDjHC8kv3I3AlRi2ssH3ezr8cRGFYtnLO9WcOXR59bU59RXt+ma/LUbf5Kx0
dTwdJe+70c1cZ8M5QCJHFxvfG1YRo2a0/SAb6RXv8I8VlNm8qDK05ihZDfwNso7X
kyK4NTt7tLaubi++AY1lWfP4jJAsrcR5qO5xHdvo0IPOxFOJG6gR2InyzqGWf5oB
YSAoV4i+s4LoxhxULbwVX9U+t9sL/3p8dr3R/9XANTnx5Tc0UAd60Swe0ikJ98qi
W5h3GoPMzmu3wq2ZOJc2sDrQKTjDTIfF7HLANZvmv6DcCpcCWasbY/CPjGielm38
qurWShquLHwwPPrxK+jnA1hb6HFhTXJ6wpNteEZ2XwSRhsgvJtiLliUsgKXiDiFK
T3yjio2yFSMispifqx0BHmKF8fekEi3A+T994MDvITbxS5AN2pmE8hTkQQwCMrFp
2iYcUt+95EF7/lBCXNtQc/tea5eLf901Ajy7Nh2sUY4SnWSzHOCK/c++6Kyz8NQx
auUM9oAUm0D53Bz844nP+ZvwmlrwH1T5/dE2LYEqcjUntv7cSnvGvsZj+0NlLGRQ
XH0GB7pl5IkcOUYts2N4Q64ExGulhuNnya4wvf9mYSAkOxrjLLqqjlxRqeT78RLZ
J2zroyq6Zc4KtmZyL8CWBMD3mz7sFDBluoYi4i9FbeY3vJPacnP2CvPGtk34UDyO
yqB10EJDtszZ6vBENUNUtp7DzLrIm1BDlUiH3boG6iIFzLBWfoXvghtwAW+u5Vzv
H62RocqNsegbmzCmJnGb+k28BPWIcasIKPEl61XiwYnaiiODAqBOPaJz10sVkCHB
txuAIkBbIwFuqEBdBeMeKh2TSUG0MEI0f+4DBMeXClKhDi9aw9XgHkkU44mc1Hgv
sjuqAh0lKdrUUrIgmlUHFKGy8sUG9QC294At4ckc+Zu974dYnYKw0ynkJVazNCTt
NOzUldBqDDL29UlHVwJFwhNAG3mTINkLF8+hhKmRMxy29vAVgVMPoLtL0rq89Fr4
a36AgNAs8+O1Ltvj4lDodsWYB425Ei1K/cBw2lKwN46tD2qF4GE8HkO46FvUX8CC
bOSX2hd74ZYKkvkj+yhFQb31GIaHpRfEYarUqMl/sj299Ie37Iay1a6w43OsaAju
/E7Ed5ygz11t2B/6tB06B61ZJV8zMerwS1Lqs4PLu1EPN/kNKCo0/obDHF8ij88/
0o6Ghhwhiqxpqmj9s8DjWic7OL3EfnewWz0NoYBfKxV56Q+zjCGo+VOikFCDXdgT
zRf/V0seJspb48+GAYG45OnuolPcNVCgSwBzyhYrt7Wqzvt6VBfUqp7hrTKh7HHh
n837lzitiruFlkezzZcfCVT4oKA/BE321HWkH5sw4CNScXdEyM0n0FLNmOXMf4Tt
MFzeSrNkYgiM246+5477DoMrRfNJZj2sgS7NN22dK3Qr9pA0KP1tjSjouWrkSh5T
xVb4jVEOtnZ7NApqO+U+a8GXErdd2sAgnwFn/vfpDJzD9kq82ld2j5O/Y/P3CG27
R/Mgw80yCv9jOA+8+2mpFKRWvqrp5CbEY05VUMhpsh5dGUCYWlIseFno3ULm3wCV
5I7n38Cl4AUVsp+uUYqkrzi4KmELhzF2WAo5aYbEqpKML1n+pKA8pCPbo0uDWJO5
f0dt8CDRDv8g4JlmKRuIdHKL1XcggVaNfs8T+d9LhXZxjeD0X28G7ac2jYnT4mtx
x9qyVR2nQs2msm1qN79ct+6CWIoIosVdmeyWKYoDDNspr1JDzzcWzO8K7gH3eG0t
w2I/Yp1e91x+7NPFcQUc8S1u8hGpt7TeePSCgkeTlyhT9xmFBkUP5YzlsOreEduU
vMDMHgV5n+N9EGR1Q8lYvLDUO8qNHNbIgBb9D5uQ1gV8fBd2foXfWriVbdbGsLpw
uilGfJ/RB+CxEVVYcKFF30Qas2Ol7fJVaZjjGEEjjR/gqw79EmWzGvpySoHxtWXl
rMq4I/pFkclmUs5+xn6sQC52O/MwEtwR3ZXFjMHZmK0V5BuD+cXpJnWfZuBpUbrR
KSJL7R9mtDz1H3hqRd6JoGoyTt350G3mkKeEzraAgtRPSoPTYWeYCnsqG9CUaySy
kLB2WXGgSCUxWrhF6RdLrXpl/BnlJ7dmGntiJI4U08+SKZvlomgy5EFcOom4KN+j
leYs6OKhWdWok24J9ikTplIjAfpkBDqNM+3f653BTPvyhDHB4FBRVT5wBnQhlS2i
V3LeUt/12GgjW9sBHHtTSm505R1ThsafOUw78iKqG6gm7W8JTQ8qVhkDoyqqv9ko
mqKC/vSZT2+QvPC4dblUGpoT1oyanWjl/fs5LEF5vNqtOdnGKfvg+sBoyaRSFFpZ
iGWJdS2BtO162oq73aB/5aoR+4ar3z+FvNOu8l4SMfQcaXWztIlVhYc2EUTrG0MI
C7zQfEPF3tZcu/XtK4zxtdU1weA1Rgx1ls1dMtFGfTzFnPAdzcV+eF4u6OhXYsDC
elwmeGzN9q9i74qtpaJZJ9hO9bry+fVaIa+yD+1cPaARHeSHGX8SR0nY37jAFyOW
V3weRPXNiv/QWIirnoCBlZkjoMRi+JGvE5ikGZVvx1lz2HmhuxYe3Bcj+XjsILMk
Ay6KERw30LOMWKwVruDYbYMYA82zCiEIA5mr1LC7pPF8njpFaaQoIcI9JOMTqbi2
Ys6sZrwOPyG2cjbTGMxu1GTSmV/Bu3tXZ8C3MpXPeeITcaghhw8R0Kz96+AeTL6X
Q5MWqTKijmIjYJadiWIjs9Ho4Qvt9wrLThqI53BCFOIb8FrF7TVQ8BiEtd19Tte9
+AkUWy6H2xDe3pCSxP53OWAh78kfeRefdQ4DvQnW5/vLFnKI4dYxZrhJ6Y+Q25PX
d7VIlAlA5XPKnK4zrY2G04N/5jx25G38G2TWTsO/GAdo3Y5pqqMOpU6UBSHDHYIe
hEiw2zehcrW+A1Q66iIn5+SFoB0K5p7CKQpO5gaD2Jj1M6s6C5O9Q9Ahq+Lhpk8b
PRkZm3MNWiFQlHqUKZUsQU9poD9eyfzODFUshYiaW9UMkYOaElt6CuMdROFgLoQ9
fvbhx2AmGI8pK7hVy53UjOiyA8c+hTFFnuay8qXAGTHrZG4BuF6VzCV/7+VRihgd
XSmsV4khTQHcEX0Tc/9ivVx40z0GFeu9YE0lDiQJWCc1TNULyQgLyNOi91VQS6sO
PDXmrnEBos8v9HRqPXUUxoQq6fTESbr6aUqLEj26DigP74vfprmMXJyV0B5kLqCj
2Gk1bULIpAdKBT/DgUwvWdnolHkMBUG2qtMQ111d5VaycoPWpZ1vXe2UKV0Mmnub
5fuMU+tkZSY7fDihoOI5Frl0VbrnIs8PVo+dE7pI2SzIqj4siElb3f/6sgezeycF
3z1Cq8NRiB+Ko22XYRbLsJJoNmdGdqYlY0tHn6/BPoVBitLt4j5Sdixf8wvA3vL+
LGpcuAnNBU76r6qGrL4KXBIyiHKB2tXWfMgCL200kOH6yJu82t8k0miDIdjPo+c7
sR5WJ478ABJ+1nxXQhrFP5bBTzD8ONHjA20lkkgA/VSyrjD0TQ7jk6e9znSCnnRq
zUSd7DPTOKAFcq9m4MC1XWsc7i9kUfGqSxWjywmUxrrDR7CvvkYyZTveYSkJnugK
s8sC19RQdBE45DzR9eZXyG/giiMYXmEjtvp2dS8B64BU0UhraIpS5VQEFmCJFN+X
rkq/O3lY97/NJ8JQcisMPZ7uG/dUuyfA8+QOMIuXfZgpkJYM87gDhgmrbRCylqJM
5JUB1ITv0gE3yNkwwVV9szY7M36SIu0gQ+5+rxeEJRk2vNZpEWysjbQG2R5SHcaF
XQ65sGOwZNUCmO3ukuvynVNB1L4NCtyhXZlRnXzqzlNfc5AHc1YgvnMlagBAvphF
XGNaZ/tqvazlYMkhimX3pJu8zFMSZLfdUDnOLCRiy4HoDEuh+7RxG3LIPQXd95PU
5mXXAxKKxGzNSrQKj4BrHzOEqd8c/mECxqdjbufFYqaIcaZv8EV3neb0lzMqRZv8
cQ+nEQnBoQuZu7dQ48/36yCpii9JpoBcqb64RZtMaAK/Wp/jfZAStXsPPs7uqDhQ
J6nexfZ6ZazbANWHkwI6RoERotAfI8kGFEuqlcTOE7sU6/Qkct5xAICv2TaNIsfK
WI1vZZqEgQGNNuIxsYAX7uaJ28Ub73nztzIwe/rJidv1swC7joQrLkSKSAw2lJzC
CuwGxSNLPvHqgwLW9TXsuJ4PycN2FDNwfgP2ftCBwtq4ST+cWvWdmmYs5fid3cyK
BXlF56f76SsC7V1l4BUGsoekNG20ADV7s1LRxkAe4BMPy3uGQz5RS9AdjszPbLz+
Kr7pFTUlg+L2dBYYAGbq+O/fyZ1QVVYWSG0lVhYaO+Qv5cazFNDQ/nCWu5wL4ztz
Vk0QptYTRwUthwTLRIfXetFn6DNpzxZDqFY4/YtbAZt0vN4Ud/eWeI5ki2XeIkAB
O6ODmE9v3ZJ7C9OgwKAR42PwC6OTvHkQxOY9ILy8rqNFn3xCFtS6MobS8PE5GTtZ
HP0C9szLzbQbhY7qCUrk0QA06BjtAIr1DuC4rRae9tj/nqHL/74xd7UzXOYx9ik/
pXdbMn0sLunuMPZ7iikDIVMuMUkraB6eBeN9HrmLMaFCWiBJyS260kkZzlNJ0/8L
I9HncLTowuHihRXYlHN/Vm06e9bqpEOpmPgC56eiFnz/bJXKcYHbJh1v/zTKJNbE
zKgIMJsPV/LSU1QUfx881+4PngH/E5mslXaH6x6RUn5F6qJlrLTDp/7hr2EMFvQI
7SfvgmBlNto8u09y0+ve5xVlBFLPXWio3k3wt6GJyGMvuw6pYz3MxF8B/30p541e
+ZvuJUAZSwp2hM8CfXueGkyisvb1md1AqHVNBCT4jaL4fNrIVYvpsq+nT9F8Ed49
YcmKfea1G9iC2mw9jcb0voNvpgJ/uiV7K3xX5HFfviLJ7mSO8HLSrbibtKFQ7RYl
C4bfUKzVLJaxstGq4/qOIPKMfF5uac727nHlLG8myxbNd96chH3hChdH9srGc0YS
Df4kG4Y92ayOs7hiAu8KSwwZ/vcUbQa11srbMwnIdVz1FGjEXN7gpqBWdVKM6Alv
1RpfFg0sa5LnUV1jqtjL01fXydczozMwx2g4UxTlUkYnHCj90UGZdNQy1OoTe2Ja
Cg7wHZ1hwfv6UeRI8bKE5giVIndXZ4judFrdYGXqSAylRzmV52s7SLB2KGyLeoH7
Xf3/XPXh1ZXbTqEmxyJnftSWJN8WtvigckcDIGBudIFGbriWMxgwqsItACkq0yCp
Y4dJigi8uwIyT9h2LFO9is0PXoOw0BuZSkjt2n31lpL+GL4qo5LSP7T2fGgYPEoa
PBafLi7H6GnjRFpHDdmMLR6SoKr0KXEUW+w2uBtsH1/yus8zfmHJ47Vw0tEMLDCj
8oX2sqGMphrYR49F9eNYTEj1Ell9mA78QlrSs4A/Rk0c3Mj8PR1gi+ll7rL2dwJF
l672FwOffCTAdabMWYmHYo48wbDwRt7fEGHepd8zL0S5Y/7/3GmhP880k8G81h25
GWai/K4ODf6T2M8CexmwvlmjeamnSoCydtfIQYoGoqgqs+PB0ox2Y829S2e3lKHJ
v/2Ld1fgzkO4hRVN/Qi6F20duuAnAGpgBPlNt/NIjHSmWN2qOXOnAPg6//HNm/MM
ZxdEHKhSzin73SvM0LcLZ7D7TqUquXVLz5skmmz3OocKlBuwnAojjg8NsoFDMsIH
lxFcRP735hovNDCpm+ujHcjGO1zlw0m7TaJfnJ1JFXXoiho0Ap8RayEs5HjYd3JF
4ea5m7rQR3LrnMONCEhrb9lDvF6NY+8HfxxLUEoSpY78ajQ4BrjMQ4OPI1Xq/ARs
TAYb0+BsT21WZs/lZyB2T1HEdristIll9oM+G7OjrMnucrrNwd5JYrSuvRbvl/87
CPzLhFaV4vvLWtkYZ3SGLCWLnESrawU4A3oXR/Obf/x9Pwd3d+k3TXHh5jjKpFYS
pAWWkKe0aEufFRMo9YoyH9cUU6WKDAVR5XMbyV91sp0wds9X3i4rsyBy3j5KDH6u
J+8eu/Gk2howvxJl/JdqS5+DtOx4LBpRJszXjR9Rf74hWTXcW5QiMnw8agrGf4S0
/HBmUHEDaO7Ebl6fKBh7dxcteYv4H3v+wDS+rb1ne5KctUzvUB3dn2aMQ3BwnZ+r
as7a0HKq72yWrxMaKF6+bP9i0NF/FoszPt/7NkN9OSt/ekT1NIeNbkjqVcQ2vkYp
pOrFoOGOLkRrR88N4HDHeRKrdzR69c48YaMMq1UwaSRz83oZZHK9e7AB7Lnz/Y6E
Cl34rc8U0l57OQ1bYvaCSDngbHdFiOGz+o9XFT0irPypvjYj3Wtaca5Zws/JKqyR
FpsIRNlVOPGhEXgpmCgduSHWwtsJ7Y7eT2jTXvBZ/KTpRMQFya111E5DJSl//fWw
7b3hKfYv2HGAQWUadEFLmnHiTQhEBv06SzFQIYfuTD4wHP1g1Er5+fWQIqDmHjMV
/TsiPq7Iw92w9r+PPuhIoB/+XtJkOabxCcVbv5SXJ2iPuZsC6C35RqwuCbu5DN6W
X00BswTE8tJhAL2RiY0gk4AkSTtXjpa1JbgxaJ/xBW6xaAlMvxGT3aBRVYdT4cFW
gJtOpDFFTkLvjs7xDyLTD30xPMiUg61zwIpjDW3GOt554v0FJO5r4y25PEcCk1Ru
QBEPzEn5GowTWF9C4ptZmR/Bj0hATf52/zRktDjuIvNB7FlHVKLVJbjkWPvhQaFh
zBkExA++hzJNDiEuhny6qis0ye1P6QVzpHwAnUU6tP7lAPpP3gMKzyDZvICGcyhT
sJ5+o1VmSXW1A0rWyHjo+P5ukN92azhAMvDiTUTABaMzagHq0o3HgG1gNa7399za
uO1bc5VKc/k7O70ztEdbZevqckLjA5pLTDw1nwd9vXq4KFgCTLJCI/HL8xuAhip2
uMRx53CXAOYsbGjWDK+vQjXwq1SvxP8Y1eiEeWyPcFLlMDOYgMU7DbGv8RGJacm3
jBWKENJBVK/u5U2UTxTgnMLsZFW392f75rHmVXlNOuF9jyUg/bXDKV9aB4NhmVe7
H+G9l8KsW4GDRI6jaR9FEydLOfhW5MsNSiU/1v8PlYRlDNpc5QiHRRXQAPUHe8MO
5qQesNRkXf25v3JbgymMpJoYB5eWTYAafNK61AxpC21iRovrh1AOMaXOLBRZ7TLO
Wzcd2PAYdbVLHY2FRAxDpLBFkBzM/KdyDzSTBszydz+0A2qesZ6DLJXY/sA/eL9B
N0gXCrwPwq1UpEnSYQbimQqX1jdoN+NHusqirG7VztZryA0gLtLTQJz8+fn7XWAq
4aq4CLBHfvClobh0m11u+srn1bgw8OJr9qvrumz0/2mtRYcci8anc3YPwXEcS2n4
QolNlmZvfcSNAfvgsacrQNFoN2eFNukvEFFtLEL+tswiPICv3RcbH6wHb2hnD8mg
6NPPYJOM+0balZHzhXlANJVdVQrRVgvt9StwOOfO6CbF1jVmS2ZH7eDM2e9HawGC
WuWlhJ7VVZ7w+CiDTgDhnnhtZl/4vzR+w1VOlgbqWQ7v3SJQJIcoaWQAjj5obSwc
6hgzWX0rwcYiCKrpTUnwhXn1C6eHZfNGMUfc1M1qj72J0PVQKm+wDeQ9TuyJLhfZ
71zP5WhTdMhnIybeYzSUCUd987koSF0rmF7BL/mzXLN5ELIPy3U4p7X0CxXSlIdI
bLxqRA2Ui5XFjN1ZkHyPQniJ/rzT1GuaBdRENsytYinSRi7oHgw3WLdKH6peFOor
UBOZYZuqjj97vNKpM/mU6gVOhfvgOsNNVj+Asdke/fx73xaBPT4RG+kuk63RnvZn
YZVyIudjThGld6PxQpgWueAtgOuZ9f6A9ddJSGp0vv3YsQa3welNKO2K9VXuGFj6
b7KpozSHYmO/5XFBjqtUIdtzdnW8vHpk9NO8+kN8PVQeTX/gIxEPDkbj+n9rx89T
qCFvnWeQOH5zJI7iNRV9qmxdfzmn4s1RZveMbQsnQrxUR3wDJub50AEccCOYqTpD
ad7bA+F8rJ0OSbgAIIvXy4BYonAd+x4riyrcHN4JuIK27/qQ6f204B/fo0eFUuVr
2YVRrgLggEvxE/WP4gCCtRskWB3edCkU5Pmjrg1wxrb2bc0/acxfZUj/p93d+/CZ
VmQs46bwcY1htAWXKjwTLajITxyDaGfoV1kl4LtkuD+xDUNcW6Ilt6ueXYYUirbO
CDXJEVMKLGvOK5usGMr30dR1nEWdIDulGFYYdRlkNQ28OZIbSU/OH7AzeYMhP5yK
vbBq37xmGzvv0ybUgSEobuC/zaaIZzFbeYLeIAwF0Yw9xUoPSRFpck8DPcfm3A4p
G0GYI+z/X5qXZzntS2+iHtw3ufbBCaN9H3ZouvgTzZL8dB/X0rJl/aDvMZWDfLjP
hq74EB7+xHmrYtwGqN6CSiY1Bzjl5wJlUdCnO2OdLaD0O6NoLtDvjw/7YKYnlm+a
GkCwyWrfZl09jKYCpKFzBfcms45xrwrpa36DmjVpLJVNlB9hoUMyn/AdeDu3Un1W
NWjgZ68GARTeRGLE3NNj9fD8BE5VAtbFGo+fNwB79ju5LomEOIuhIlPIebKt/rOK
zT0mhpDn6fdu+eY/zWxkP9kBbgiaqJlcUwSegI2pUI8ngXJOWgguaQXZbNadMCBm
cLnqY+m7MzMYJYudHPac/U+rN42kJmN51U004KhvvZcGIvGGCKvw3CToGBBWpRBZ
YjNCK+w0I4KgBvqidsPIxIuHv0cVSqCEjETwSaGtqDkEoup+Xr68/q9mUk58fDPT
uQA/Du03xhn3dfX/Bn+DhxKrnxhi3ofmAeCZbR6RzYzwwPMnudBlYI3uwhNXI9pu
GeXle5t11txyMJTNtR5PGfQE7QZs9N5oJG+KQXdIA9UyOWDyOizRRndEj1JqNA85
6uoqFLpSwL6Lji7B/0BAbxNrqw5G/13S5iadBH0Vov/S8afCRLGrGT8JLp710Ijx
lmMlkaB9xNmfc00beotaf3nMpzbBGOIoSYxu9RnA8Y0SHAo2L5WXTlQWGGQY+hOa
XnpFkc8ULqVnmhF0vz1G7iXes+kag8kn77X+tFYdEl9IeyMl8kOU1Co+bzXyrGI9
q/jNuf6pfkY37k+qOEoog6DijWPDvexFrwrr/nIoSGtCnbkp34uq7VNMpJQ6AVKf
P3fOOaTFTqvD1SrEvih/iSE9+q6XfWCcjH9uWdtFMkOAj6XLdBPhisrTMY/DD5nR
K0k41W2+ULfyZ2GyIW4QKXBLd12mJNh1X2wbihDfWeVvXMg4lWrcBVFi1YJWMUMh
MrrIoVbBxZj3Th8Rz3UXzmwI89to4NSHzeIqeps+2eqP0L0Gx+Ga0mz9Xfp03jSS
ZQqn2Ko2kvH4ejMFplO/B1D08ieMiQ+LNO92yqHIk+4HBKdVaJ58j69xfyLCPuzq
7l0FXGPpu7u09X6QTiAPMFQhxDDGycvF/dLLyyWqiDWWUZM3PwUNT4X9SJBtUd4P
u/yFiBDENUzIxwq+PbTjW1QIrAtpJtOVcclGeY3oTQ8bCP5026mNv+Ir7trCa2xR
kEFnEv7yeOWWFyQ240tBCoev/wvarqKj7gs1xaomF6vIdoemJt4XXN5aMYPqNdNX
RUgczVExc0WEusmGt+W+rDrRd/LxMX0UW/cLIoIPzDhTa7+imFQiOZcaxBcfT/iO
HImdRucB8aKFhU5UCNHsaNKbQMsabHGb+Bh032oX4lL5FjB/TQOaLsd1mXlJH8lJ
7gQkSrEotY6WaqmKuwXpEagNX33xaoB+PtjKwbVec+uEzB7e+hlvI1tZ/lsHCKBZ
Qxf9KYXLSRu4rspq1i9VrWKU298Z7riAU/cnCI/OyeJR2dXQnjUDkN+FZPHvolV9
dT1Qt4DGKE0f/vGpbti6GrUlbLPSX39e6Wv+M/wNNCuCMyxEa579G3hgM3IfwLFL
inRCEeZMAnHnBQOjoq1zhP92NCjcMDPNJViwkraJ/Rs14W4BFGQLPIzGEtvlZiiK
+1GyKSzlpz/rdkzAz1mk1Hi4B4vtOmJ0JJJwOXJGNXC13QQxehBO8tkuwuikabDk
Dm3LOR1JmMEJNaJ2BPbBZ0p91wsatO+IiNCpf3K+SI49YIEL1lECZq8H/NsPzRVJ
e/KZe/zjJWVaEwy3D0FFe0p+LwxAmwOrma/OWjnQh386O74PwFuVo73sxbRR1Z0G
u7O9d2YLUOkOMAupwO2cte/DLWUUI+XO4qVnDIepRM1vjRO2FibKS70NC8bvGt0M
nr6gb186uBRfscBvMejhStYP7T6KJpP/4hejKBfvFUM0YSnHiJdfLrygssyo6gtm
mSaU8tDDy9WXZBH8qB1NjbpCAbzEVhNo8G5Du75dlbiAjKtQymduCXP5bhtZqod2
JXCJTXEBJAf/PKDmc4ioGr7bnWTR/xs9/WRYAVIrdhRBm3xfqwQYCxDPmom29reS
hZ5Q+qa5wElH7IqBZk9k/hZTL44rC9m9haL2P3XcaujauwMcg8z0KYTK2C3dV2gj
zq16ZhHM4FiXnILMMrz/diCWwpklXoPsE6rudNdH5vODuYS4M6THxEBL0g3hIR1H
R7j2qs32w6Y0V9x8djWEXF1eROrjl4OIzFYHxOCu4NVCBwdNzL87ekz0v6hPAXXE
z8p6chfPfiiX9G3OnFTUmiW9VufkFYQMLLnry61HzL32ahXW48WM6zM3GQgTH9iI
id8iPZLSWpEjXEn9hc7e4Bl2BTm+GTL2Vd9G1FBKUs8eYk/KiB9CqlTYrXyKQKfT
vLPYoDwPn/jxSnICPs1GVPfSFMu/u9kwbL5E5EhpanVBGgsHirGIcU3hl1UFxWXH
KW26tk80FP5UIS+eAGV+sFpwPNUrf+j8Ze9nvXRT9Iiny+ygxYhBCDrwTYaHpfDm
DV00KP1ZYNOfdSXKVejI4GNMWKViHTggOLsxxUyQR46S6FPSH9hkvVsaloKw4ozk
SFkJRdZPTMOQflZIFwPL01bTQ1bEqQHFMfa5xYizOxBj9KKKsXtMNzVMisMUOytw
UvFxlCohVSZtqGlIkK9rR5trsSUzRO7SVAYMMUsC++Uq8Z+0Jrqq8eKXhvaky0u5
Ehs+PBMZ2rXt2h33yE3frOez3z63UtUhS6bsq+T2ykoTiYP5HaednjMgvkCOix9D
ksOTQPUZu7Frp9nVZmFoFru1htvN1rgtdWkDFVVGOGrR9O0m+5yGyDQw7k0nGaDw
Twc69mXGw0QhFh1V09oAZ6nAwjOYHg944N3X5PytKC5FUle1A8nL/0bTn8f7JIMW
/PoJAfVIr9fKf6uxd45D4WhBIuiIKpRShp7n8msP9eZeS0pPZAMjAlCiFB4TRaXX
spXwjZOPR2BOoWVn/6R+JZQ7fSCjABNuF0cAEQMNLC5gTYBM1JwhtQZgK6JlH928
0dKYbWHfE/WkgNfSFPA7iOhuBDfYV4bKeU8Q1rONmvOqDpVHJDGtaNnYuVgPiOdW
F+L+hHBZkU3mc/tTfVcajYXIYA435I4GBRvEGtPqIP6p/NvHA0t/s9g97W3Y356W
3HXUM9lW+5ot0HSeYgynlJWfX6e8ZNgtBUwDjX7VILI6tFGo5yrrn5ibKsLXj5RJ
O2gSimEt4pdeR2AWETN9Srw7tHiA7YKM+Qyf8JWLnAvKtamd1ej0iLDL56fj61xK
fqhLQ7116WMaWGi0oD1Pck95yl2lX1KmXCOHzxvMqmF2qgZAXolUMedFP+EXnKba
F7cjwcJg8ZA9qRsKPCZeu7p+qG6vyrX4XLOGQw1ZA1myTA9iHYHrZ6mOoBQ09qIX
8AnfSQJTZiZLsJVE3eYYTQdTPn6cyA48FSL/EJnlLVfg1p/LmPyxcuPYtLgWmx36
zQIO8gzvp6EHEcCzi0OMaZjKu5QHnpMOxnP/RRHr79CsMdzXf2t7mBg7doK31WSZ
edfoBoxt8Uxf3gbeBiIrAxKwP0Uwjn9lkikiyFQ88vX4kwWJ35kxn4zoH8yJR0Ff
ZkgnQpmCOeZboa2cfgKcAblAZW2KjDvV91OhGLblMDsRLqGpJkm3lIH3oNISFx51
zLZqFF/z3WfiqtuBcjFcqNog0a7+FOC3jAXDPPZm/ZcccjE5Yc3SkObrBzKmC0k3
WJn0IPNd5MqojzQUSOzlUVBqswAvowniuGY1Ja4yHx9xoQePMWysTVrWsJFrPbCV
`protect END_PROTECTED
