`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMyaToeyhSTGqyLsx5c4nPdfwpyL80gsfX7/0x0q3SsU
7Meeugq9FOFt475pWmR1cwzkCRgKQV3+AyJGckCEa4z/vBDOs3wyheeUGbaYZl19
pRqEwbQTViVxGqrVPqBkKun/9RCIydOpltZe8rao8mj2NuFSdA5q2QT2FDF9/C/q
DTnv6Zoy2BBuVgw/fT/jLe2Rty63qoLSJ4f1LpxMka9RiLC3RjieSOa4cTocQZYd
OocoVA7x/IjA/ale7tWpouQcfWaTPrUaS42cEmAIImoiLrKUldEvFL1vmTCx1Pwi
KWFynHLz5Frqthh5TcvnxzDpU8pasiRZFu7FG+HxNzgC0faAAUXh0CPD594knqCO
b7APvZhhG9j+AT9ooC/QtVJokthEbVNHqsqXEwfEbAoYXvvsu5u3S7VtnhuG57TK
Fxb2NZw1Bnv3sJTsU692nd7w40jtN37upLMqEjfl0M9NBltGxykZJuEaUeJznXxd
DIheCpHui65ybqC6C/HNJPNIgQzyAzSi67IksZR+1y1h1Tzbf2f1khGwQawzm6F7
GqE2n4DEoBr/du6tIw+I/w==
`protect END_PROTECTED
