`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yZFlit3YC1XA4DVB9sD8RssT1Zn/yJJfIdasqRLQF8e
7ZHt44X5iOxqOvGnFH7HkCd0UcpR1VbZ6rxQQn2JsQwptiuAse/kjSynts3v2iTz
iFa5je34cOYHxrsUC3y4LIf6lk7oPmygVGtPYUaSMr2RrtmB3p5u00YPUyT/UxLF
icvULuzhQX1IULDIQYOeFl3A9MEAHrpfeC8zZVYwssw=
`protect END_PROTECTED
