`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAYBwY0QpM1Xw45sIuMWRoS08vZgIaqo7OOqJTmE9FiA2
c3z+1+rYgDyCtrELsLHD5boSZvUm5rsqUqzZgM1HG/jgZPzQZgDxu+86l2jyCzqW
ePCroEtmOKJtpbU+uh9cP85VUMCze4a9nF+orjgX1fYnYDZIfxp+wNYdFuvilZfZ
hoD6YOx3BOGz0FPGm+6iyAAf58F04GoxSo/6Ejpv6eEULh3QQVL21XTEZggCmGZf
iRSNrPDIRwB7WbZvOtwVUmKsYcsOR+VkLvF15zw2JHVRE3/OLQG4llzheSi5DTIE
097lJh+Z4r7Gxa1E6z2BWe3MLnpe+PdXbwU021WLIJcvVJQjJsDP6SITNib5jKC4
gFBJtWEYTnsWf5W580O8Zm6W+n9x1T6EcLEoPsYeZdhqJNpCuhBTbUS7piNl4ABT
bWQUf5COQz0PrmGqEynpANiVAbBm5/6VZsgsmLlpqZ4HFVQzGqwu3VMIEK+TrvUn
+hmfdTjPDDq5uz/JFiK0k1n6ibZq0Yc2zagTn2trbUPJRgtNTWEO+m0f89WDeOdF
TjXlTegFOZG9Qy2jpwmnhJ1YB5IzrbY3+o8W9o16y0Q/fSN2oiywQ2pt/ccq2gq9
uqFJxyqRKSO4Mh+KA921P3k9GxRQny7c4JXMK4FEFQBU1OOILUpUMzc4tEHNz4jJ
jqrk6TsWbngIQFW8vOovvbipFSTkPcUyEnnNUADrVVKxD9IPPqPUc3OABBNjjhJh
455QW6D6j9tODdW+Rmy2y/douL+NTvuOOegUJDPkDP+ZG7G2yx0d9KyFlD/3Tg/Z
w5xH6L4urtQB5Eez6zcRb3Q/WIO2r9yI7UxYC0DJbC2viYcIA+X0iZ+NYHJaLtfp
+amQOdbksFQ1pCstQpDud6Q+leZMsP7vpiDsd1tkXJETNuYyjzfhXNJdBxu0W5fC
1zHaHV4g19rb3V7w9yIk68RZfE45Y2H7bkHAGMUuxrpXp0Ir/gJ4200uJEMtO1Nv
By9LBFIc/Sw7TN3o7jJnt0MwwJ7J+uWyNsbmHv+wsYnklNpVAwRxtFdiM+elykdT
kKWU7pRREbrN7MWe4M3GecWlAjZKUkh00ACxCoo6NyP32Xde6zHjqB+0QTl46KWO
b2JAjJOGJEh5M+u7h//othis4un2HkE+b7iE0IIT/KESLsDTeMTbHfHd++nenMyc
dnO9N4LJKMrVn3MKMWRSi4T6Q6dxXSwkK91p53Km39uX+tE01BBZCiFafo4NAhFR
umQWwbl2PYgN1X2iBbNl99qVdGaghtcPdkAo/84VOGWzQscD3OQB46y3MCf6Nl3A
FLq2y4PR0aY/UWmn6A+dOw==
`protect END_PROTECTED
