`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xESMuMn9/oAwXQ0Tnrg8t5mKnHQ22ElN4QIUnLqTX3v
3UVKnJCDFnRuF164SibL5OiQtrJfIl/Uy8pn/uPmrNSfSNSRjY/9J9SI0w2t59lt
w+godLr8z3DMdK78OAJtmWcWNEooNL/FiIa57cE33oy2eMUST7Q32KyCNasMevXh
luoIGBYJkgWdLYA4ZAUJhdRb2+RjPyFO4+D08ziBdL5U8dFvZTXPtYmQ0InGKJUn
q1SXu5R0Q1u9FyGe/eZnTI5PAZOVs80rfi3+o6CWAzRS9r0SA6NwAyKjgcrM3Ki+
85pneNVxkdPBCAkCnSvbkEsFHYUCi3fUgHm4nJieLiC1cVKgCgUdUP+Fe45MMctL
o5ZRzlaT4zg+DGwWD/6dPw==
`protect END_PROTECTED
