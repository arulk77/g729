`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
7y6s1nKGvzpxUeISfGMlvfkVbuG7K4gx3HBYphwFHn4KNJlvAZsxjab5KD1BxeE/
aZl7l8ZXvP7sBmRUt0WzPfBOJi46vydjW9y1wCbKDR3QPdc7igDcQDKS42Z+cyeg
h0fOq4myLLBRUwY2cOwSc/T52NW0h/DsDrW9Gd+CO+F8fA9xWxNj9plyIlr5Ok3t
`protect END_PROTECTED
