`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
fWmST6OfICxXWwAtzIUZGZIqy7GuYqcwLBJcqQf/e+3C+u1ztOQ1SM5RBrqaXBFu
tSqEOZvbLAfK6Hx3Rb6uUVXhGTHBGKgBOtEu3RjsLc+qS6cKtisD16ylE5Y4TzlS
xS6GEFvB/RoeF5dGprDHgkzhWoxoEmX/OvH3MED9vTTd95GjlKHKGZrMOOSSrbEp
MRRSvuLJcpFAAjlMHReYWorg9Hh13iyX6Sv5ShKs2+maqMJiMcynbuEQ87yGxzZQ
ajwNvC2/BDAfO9nMcW7j7kBA0uibuj4YFRuLjdacVVFikED/P+lrHBqk6eDPXllQ
qAdC471rPpmuRPDtyWXUC2itR3qhKQzVzV5zToJf5FvhRY9IfDQ6ZT3DjO6BDQnu
M0jla+38zkvjFdes+Ric4cAyKBwseIyvhNDaYtbbFCf3vax52lJHhXHlzbIMfcD/
4n1N3PG9bN87bmMDwz12mxo7QAqG3uO8+LxDRRdVbs8=
`protect END_PROTECTED
