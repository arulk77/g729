`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOpgQHvynx0RXqzqlqxw0m5Sr+WxUAw68dnSRWI3QAYr
1NY+tPEuyKuK4ELlydIwPc+tQz5dKqcFoUKbnUjnytV37xP2yPI+Eb6LY1qBIGg6
v5RUAyQ026sqSQWoxi5pVFn8/VI5hwVrWkXDy1q27b9/rzG01oM2Xv2KlaPB0RUg
/QoWc9Y2pGrQTqBGPfra/mhyAinbralcljtFK89qbc9PGP3WdiM6VXR10vcMo3Dh
wYR/f26ppGHf+Kbjgrt6GaZmGjKjSF5k8jmkxh+92QWtdlDy3SH3Sxv6cgjUXC4Y
`protect END_PROTECTED
