library verilog;
use verilog.vl_types.all;
entity GTHE1_QUAD is
    generic(
        BER_CONST_PTRN0 : integer := 0;
        BER_CONST_PTRN1 : integer := 0;
        BUFFER_CONFIG_LANE0: integer := 16388;
        BUFFER_CONFIG_LANE1: integer := 16388;
        BUFFER_CONFIG_LANE2: integer := 16388;
        BUFFER_CONFIG_LANE3: integer := 16388;
        DFE_TRAIN_CTRL_LANE0: integer := 0;
        DFE_TRAIN_CTRL_LANE1: integer := 0;
        DFE_TRAIN_CTRL_LANE2: integer := 0;
        DFE_TRAIN_CTRL_LANE3: integer := 0;
        DLL_CFG0        : integer := 33282;
        DLL_CFG1        : integer := 0;
        E10GBASEKR_LD_COEFF_UPD_LANE0: integer := 0;
        E10GBASEKR_LD_COEFF_UPD_LANE1: integer := 0;
        E10GBASEKR_LD_COEFF_UPD_LANE2: integer := 0;
        E10GBASEKR_LD_COEFF_UPD_LANE3: integer := 0;
        E10GBASEKR_LP_COEFF_UPD_LANE0: integer := 0;
        E10GBASEKR_LP_COEFF_UPD_LANE1: integer := 0;
        E10GBASEKR_LP_COEFF_UPD_LANE2: integer := 0;
        E10GBASEKR_LP_COEFF_UPD_LANE3: integer := 0;
        E10GBASEKR_PMA_CTRL_LANE0: integer := 2;
        E10GBASEKR_PMA_CTRL_LANE1: integer := 2;
        E10GBASEKR_PMA_CTRL_LANE2: integer := 2;
        E10GBASEKR_PMA_CTRL_LANE3: integer := 2;
        E10GBASEKX_CTRL_LANE0: integer := 0;
        E10GBASEKX_CTRL_LANE1: integer := 0;
        E10GBASEKX_CTRL_LANE2: integer := 0;
        E10GBASEKX_CTRL_LANE3: integer := 0;
        E10GBASER_PCS_CFG_LANE0: integer := 1804;
        E10GBASER_PCS_CFG_LANE1: integer := 1804;
        E10GBASER_PCS_CFG_LANE2: integer := 1804;
        E10GBASER_PCS_CFG_LANE3: integer := 1804;
        E10GBASER_PCS_SEEDA0_LANE0: integer := 1;
        E10GBASER_PCS_SEEDA0_LANE1: integer := 1;
        E10GBASER_PCS_SEEDA0_LANE2: integer := 1;
        E10GBASER_PCS_SEEDA0_LANE3: integer := 1;
        E10GBASER_PCS_SEEDA1_LANE0: integer := 0;
        E10GBASER_PCS_SEEDA1_LANE1: integer := 0;
        E10GBASER_PCS_SEEDA1_LANE2: integer := 0;
        E10GBASER_PCS_SEEDA1_LANE3: integer := 0;
        E10GBASER_PCS_SEEDA2_LANE0: integer := 0;
        E10GBASER_PCS_SEEDA2_LANE1: integer := 0;
        E10GBASER_PCS_SEEDA2_LANE2: integer := 0;
        E10GBASER_PCS_SEEDA2_LANE3: integer := 0;
        E10GBASER_PCS_SEEDA3_LANE0: integer := 0;
        E10GBASER_PCS_SEEDA3_LANE1: integer := 0;
        E10GBASER_PCS_SEEDA3_LANE2: integer := 0;
        E10GBASER_PCS_SEEDA3_LANE3: integer := 0;
        E10GBASER_PCS_SEEDB0_LANE0: integer := 1;
        E10GBASER_PCS_SEEDB0_LANE1: integer := 1;
        E10GBASER_PCS_SEEDB0_LANE2: integer := 1;
        E10GBASER_PCS_SEEDB0_LANE3: integer := 1;
        E10GBASER_PCS_SEEDB1_LANE0: integer := 0;
        E10GBASER_PCS_SEEDB1_LANE1: integer := 0;
        E10GBASER_PCS_SEEDB1_LANE2: integer := 0;
        E10GBASER_PCS_SEEDB1_LANE3: integer := 0;
        E10GBASER_PCS_SEEDB2_LANE0: integer := 0;
        E10GBASER_PCS_SEEDB2_LANE1: integer := 0;
        E10GBASER_PCS_SEEDB2_LANE2: integer := 0;
        E10GBASER_PCS_SEEDB2_LANE3: integer := 0;
        E10GBASER_PCS_SEEDB3_LANE0: integer := 0;
        E10GBASER_PCS_SEEDB3_LANE1: integer := 0;
        E10GBASER_PCS_SEEDB3_LANE2: integer := 0;
        E10GBASER_PCS_SEEDB3_LANE3: integer := 0;
        E10GBASER_PCS_TEST_CTRL_LANE0: integer := 0;
        E10GBASER_PCS_TEST_CTRL_LANE1: integer := 0;
        E10GBASER_PCS_TEST_CTRL_LANE2: integer := 0;
        E10GBASER_PCS_TEST_CTRL_LANE3: integer := 0;
        E10GBASEX_PCS_TSTCTRL_LANE0: integer := 0;
        E10GBASEX_PCS_TSTCTRL_LANE1: integer := 0;
        E10GBASEX_PCS_TSTCTRL_LANE2: integer := 0;
        E10GBASEX_PCS_TSTCTRL_LANE3: integer := 0;
        GLBL0_NOISE_CTRL: integer := 61624;
        GLBL_AMON_SEL   : integer := 0;
        GLBL_DMON_SEL   : integer := 512;
        GLBL_PWR_CTRL   : integer := 0;
        GTH_CFG_PWRUP_LANE0: integer := 1;
        GTH_CFG_PWRUP_LANE1: integer := 1;
        GTH_CFG_PWRUP_LANE2: integer := 1;
        GTH_CFG_PWRUP_LANE3: integer := 1;
        LANE_AMON_SEL   : integer := 240;
        LANE_DMON_SEL   : integer := 0;
        LANE_LNK_CFGOVRD: integer := 0;
        LANE_PWR_CTRL_LANE0: integer := 1024;
        LANE_PWR_CTRL_LANE1: integer := 1024;
        LANE_PWR_CTRL_LANE2: integer := 1024;
        LANE_PWR_CTRL_LANE3: integer := 1024;
        LNK_TRN_CFG_LANE0: integer := 0;
        LNK_TRN_CFG_LANE1: integer := 0;
        LNK_TRN_CFG_LANE2: integer := 0;
        LNK_TRN_CFG_LANE3: integer := 0;
        LNK_TRN_COEFF_REQ_LANE0: integer := 0;
        LNK_TRN_COEFF_REQ_LANE1: integer := 0;
        LNK_TRN_COEFF_REQ_LANE2: integer := 0;
        LNK_TRN_COEFF_REQ_LANE3: integer := 0;
        MISC_CFG        : integer := 8;
        MODE_CFG1       : integer := 0;
        MODE_CFG2       : integer := 0;
        MODE_CFG3       : integer := 0;
        MODE_CFG4       : integer := 0;
        MODE_CFG5       : integer := 0;
        MODE_CFG6       : integer := 0;
        MODE_CFG7       : integer := 0;
        PCS_ABILITY_LANE0: integer := 16;
        PCS_ABILITY_LANE1: integer := 16;
        PCS_ABILITY_LANE2: integer := 16;
        PCS_ABILITY_LANE3: integer := 16;
        PCS_CTRL1_LANE0 : integer := 8256;
        PCS_CTRL1_LANE1 : integer := 8256;
        PCS_CTRL1_LANE2 : integer := 8256;
        PCS_CTRL1_LANE3 : integer := 8256;
        PCS_CTRL2_LANE0 : integer := 0;
        PCS_CTRL2_LANE1 : integer := 0;
        PCS_CTRL2_LANE2 : integer := 0;
        PCS_CTRL2_LANE3 : integer := 0;
        PCS_MISC_CFG_0_LANE0: integer := 4374;
        PCS_MISC_CFG_0_LANE1: integer := 4374;
        PCS_MISC_CFG_0_LANE2: integer := 4374;
        PCS_MISC_CFG_0_LANE3: integer := 4374;
        PCS_MISC_CFG_1_LANE0: integer := 0;
        PCS_MISC_CFG_1_LANE1: integer := 0;
        PCS_MISC_CFG_1_LANE2: integer := 0;
        PCS_MISC_CFG_1_LANE3: integer := 0;
        PCS_MODE_LANE0  : integer := 0;
        PCS_MODE_LANE1  : integer := 0;
        PCS_MODE_LANE2  : integer := 0;
        PCS_MODE_LANE3  : integer := 0;
        PCS_RESET_1_LANE0: integer := 2;
        PCS_RESET_1_LANE1: integer := 2;
        PCS_RESET_1_LANE2: integer := 2;
        PCS_RESET_1_LANE3: integer := 2;
        PCS_RESET_LANE0 : integer := 0;
        PCS_RESET_LANE1 : integer := 0;
        PCS_RESET_LANE2 : integer := 0;
        PCS_RESET_LANE3 : integer := 0;
        PCS_TYPE_LANE0  : integer := 44;
        PCS_TYPE_LANE1  : integer := 44;
        PCS_TYPE_LANE2  : integer := 44;
        PCS_TYPE_LANE3  : integer := 44;
        PLL_CFG0        : integer := 38367;
        PLL_CFG1        : integer := 33216;
        PLL_CFG2        : integer := 1060;
        PMA_CTRL1_LANE0 : integer := 0;
        PMA_CTRL1_LANE1 : integer := 0;
        PMA_CTRL1_LANE2 : integer := 0;
        PMA_CTRL1_LANE3 : integer := 0;
        PMA_CTRL2_LANE0 : integer := 11;
        PMA_CTRL2_LANE1 : integer := 11;
        PMA_CTRL2_LANE2 : integer := 11;
        PMA_CTRL2_LANE3 : integer := 11;
        PMA_LPBK_CTRL_LANE0: integer := 4;
        PMA_LPBK_CTRL_LANE1: integer := 4;
        PMA_LPBK_CTRL_LANE2: integer := 4;
        PMA_LPBK_CTRL_LANE3: integer := 4;
        PRBS_BER_CFG0_LANE0: integer := 0;
        PRBS_BER_CFG0_LANE1: integer := 0;
        PRBS_BER_CFG0_LANE2: integer := 0;
        PRBS_BER_CFG0_LANE3: integer := 0;
        PRBS_BER_CFG1_LANE0: integer := 0;
        PRBS_BER_CFG1_LANE1: integer := 0;
        PRBS_BER_CFG1_LANE2: integer := 0;
        PRBS_BER_CFG1_LANE3: integer := 0;
        PRBS_CFG_LANE0  : integer := 10;
        PRBS_CFG_LANE1  : integer := 10;
        PRBS_CFG_LANE2  : integer := 10;
        PRBS_CFG_LANE3  : integer := 10;
        PTRN_CFG0_LSB   : integer := 21845;
        PTRN_CFG0_MSB   : integer := 21845;
        PTRN_LEN_CFG    : integer := 31;
        PWRUP_DLY       : integer := 0;
        RX_AEQ_VAL0_LANE0: integer := 960;
        RX_AEQ_VAL0_LANE1: integer := 960;
        RX_AEQ_VAL0_LANE2: integer := 960;
        RX_AEQ_VAL0_LANE3: integer := 960;
        RX_AEQ_VAL1_LANE0: integer := 0;
        RX_AEQ_VAL1_LANE1: integer := 0;
        RX_AEQ_VAL1_LANE2: integer := 0;
        RX_AEQ_VAL1_LANE3: integer := 0;
        RX_AGC_CTRL_LANE0: integer := 0;
        RX_AGC_CTRL_LANE1: integer := 0;
        RX_AGC_CTRL_LANE2: integer := 0;
        RX_AGC_CTRL_LANE3: integer := 0;
        RX_CDR_CTRL0_LANE0: integer := 5;
        RX_CDR_CTRL0_LANE1: integer := 5;
        RX_CDR_CTRL0_LANE2: integer := 5;
        RX_CDR_CTRL0_LANE3: integer := 5;
        RX_CDR_CTRL1_LANE0: integer := 16896;
        RX_CDR_CTRL1_LANE1: integer := 16896;
        RX_CDR_CTRL1_LANE2: integer := 16896;
        RX_CDR_CTRL1_LANE3: integer := 16896;
        RX_CDR_CTRL2_LANE0: integer := 8192;
        RX_CDR_CTRL2_LANE1: integer := 8192;
        RX_CDR_CTRL2_LANE2: integer := 8192;
        RX_CDR_CTRL2_LANE3: integer := 8192;
        RX_CFG0_LANE0   : integer := 1280;
        RX_CFG0_LANE1   : integer := 1280;
        RX_CFG0_LANE2   : integer := 1280;
        RX_CFG0_LANE3   : integer := 1280;
        RX_CFG1_LANE0   : integer := 33311;
        RX_CFG1_LANE1   : integer := 33311;
        RX_CFG1_LANE2   : integer := 33311;
        RX_CFG1_LANE3   : integer := 33311;
        RX_CFG2_LANE0   : integer := 4097;
        RX_CFG2_LANE1   : integer := 4097;
        RX_CFG2_LANE2   : integer := 4097;
        RX_CFG2_LANE3   : integer := 4097;
        RX_CTLE_CTRL_LANE0: integer := 143;
        RX_CTLE_CTRL_LANE1: integer := 143;
        RX_CTLE_CTRL_LANE2: integer := 143;
        RX_CTLE_CTRL_LANE3: integer := 143;
        RX_CTRL_OVRD_LANE0: integer := 12;
        RX_CTRL_OVRD_LANE1: integer := 12;
        RX_CTRL_OVRD_LANE2: integer := 12;
        RX_CTRL_OVRD_LANE3: integer := 12;
        RX_FABRIC_WIDTH0: integer := 6466;
        RX_FABRIC_WIDTH1: integer := 6466;
        RX_FABRIC_WIDTH2: integer := 6466;
        RX_FABRIC_WIDTH3: integer := 6466;
        RX_LOOP_CTRL_LANE0: integer := 127;
        RX_LOOP_CTRL_LANE1: integer := 127;
        RX_LOOP_CTRL_LANE2: integer := 127;
        RX_LOOP_CTRL_LANE3: integer := 127;
        RX_MVAL0_LANE0  : integer := 0;
        RX_MVAL0_LANE1  : integer := 0;
        RX_MVAL0_LANE2  : integer := 0;
        RX_MVAL0_LANE3  : integer := 0;
        RX_MVAL1_LANE0  : integer := 0;
        RX_MVAL1_LANE1  : integer := 0;
        RX_MVAL1_LANE2  : integer := 0;
        RX_MVAL1_LANE3  : integer := 0;
        RX_P0S_CTRL     : integer := 4614;
        RX_P0_CTRL      : integer := 4592;
        RX_P1_CTRL      : integer := 4623;
        RX_P2_CTRL      : integer := 3599;
        RX_PI_CTRL0     : integer := 54000;
        RX_PI_CTRL1     : integer := 128;
        SIM_GTHRESET_SPEEDUP: integer := 1;
        SIM_VERSION     : string  := "1.0";
        SLICE_CFG       : integer := 0;
        SLICE_NOISE_CTRL_0_LANE01: integer := 0;
        SLICE_NOISE_CTRL_0_LANE23: integer := 0;
        SLICE_NOISE_CTRL_1_LANE01: integer := 0;
        SLICE_NOISE_CTRL_1_LANE23: integer := 0;
        SLICE_NOISE_CTRL_2_LANE01: integer := 32767;
        SLICE_NOISE_CTRL_2_LANE23: integer := 32767;
        SLICE_TX_RESET_LANE01: integer := 0;
        SLICE_TX_RESET_LANE23: integer := 0;
        TERM_CTRL_LANE0 : integer := 20487;
        TERM_CTRL_LANE1 : integer := 20487;
        TERM_CTRL_LANE2 : integer := 20487;
        TERM_CTRL_LANE3 : integer := 20487;
        TX_CFG0_LANE0   : integer := 8253;
        TX_CFG0_LANE1   : integer := 8253;
        TX_CFG0_LANE2   : integer := 8253;
        TX_CFG0_LANE3   : integer := 8253;
        TX_CFG1_LANE0   : integer := 3840;
        TX_CFG1_LANE1   : integer := 3840;
        TX_CFG1_LANE2   : integer := 3840;
        TX_CFG1_LANE3   : integer := 3840;
        TX_CFG2_LANE0   : integer := 129;
        TX_CFG2_LANE1   : integer := 129;
        TX_CFG2_LANE2   : integer := 129;
        TX_CFG2_LANE3   : integer := 129;
        TX_CLK_SEL0_LANE0: integer := 8481;
        TX_CLK_SEL0_LANE1: integer := 8481;
        TX_CLK_SEL0_LANE2: integer := 8481;
        TX_CLK_SEL0_LANE3: integer := 8481;
        TX_CLK_SEL1_LANE0: integer := 8481;
        TX_CLK_SEL1_LANE1: integer := 8481;
        TX_CLK_SEL1_LANE2: integer := 8481;
        TX_CLK_SEL1_LANE3: integer := 8481;
        TX_DISABLE_LANE0: integer := 0;
        TX_DISABLE_LANE1: integer := 0;
        TX_DISABLE_LANE2: integer := 0;
        TX_DISABLE_LANE3: integer := 0;
        TX_FABRIC_WIDTH0: integer := 6466;
        TX_FABRIC_WIDTH1: integer := 6466;
        TX_FABRIC_WIDTH2: integer := 6466;
        TX_FABRIC_WIDTH3: integer := 6466;
        TX_P0P0S_CTRL   : integer := 1548;
        TX_P1P2_CTRL    : integer := 3129;
        TX_PREEMPH_LANE0: integer := 161;
        TX_PREEMPH_LANE1: integer := 161;
        TX_PREEMPH_LANE2: integer := 161;
        TX_PREEMPH_LANE3: integer := 161;
        TX_PWR_RATE_OVRD_LANE0: integer := 96;
        TX_PWR_RATE_OVRD_LANE1: integer := 96;
        TX_PWR_RATE_OVRD_LANE2: integer := 96;
        TX_PWR_RATE_OVRD_LANE3: integer := 96
    );
    port(
        DRDY            : out    vl_logic;
        DRPDO           : out    vl_logic_vector(15 downto 0);
        GTHINITDONE     : out    vl_logic;
        MGMTPCSRDACK    : out    vl_logic;
        MGMTPCSRDDATA   : out    vl_logic_vector(15 downto 0);
        RXCODEERR0      : out    vl_logic_vector(7 downto 0);
        RXCODEERR1      : out    vl_logic_vector(7 downto 0);
        RXCODEERR2      : out    vl_logic_vector(7 downto 0);
        RXCODEERR3      : out    vl_logic_vector(7 downto 0);
        RXCTRL0         : out    vl_logic_vector(7 downto 0);
        RXCTRL1         : out    vl_logic_vector(7 downto 0);
        RXCTRL2         : out    vl_logic_vector(7 downto 0);
        RXCTRL3         : out    vl_logic_vector(7 downto 0);
        RXCTRLACK0      : out    vl_logic;
        RXCTRLACK1      : out    vl_logic;
        RXCTRLACK2      : out    vl_logic;
        RXCTRLACK3      : out    vl_logic;
        RXDATA0         : out    vl_logic_vector(63 downto 0);
        RXDATA1         : out    vl_logic_vector(63 downto 0);
        RXDATA2         : out    vl_logic_vector(63 downto 0);
        RXDATA3         : out    vl_logic_vector(63 downto 0);
        RXDATATAP0      : out    vl_logic;
        RXDATATAP1      : out    vl_logic;
        RXDATATAP2      : out    vl_logic;
        RXDATATAP3      : out    vl_logic;
        RXDISPERR0      : out    vl_logic_vector(7 downto 0);
        RXDISPERR1      : out    vl_logic_vector(7 downto 0);
        RXDISPERR2      : out    vl_logic_vector(7 downto 0);
        RXDISPERR3      : out    vl_logic_vector(7 downto 0);
        RXPCSCLKSMPL0   : out    vl_logic;
        RXPCSCLKSMPL1   : out    vl_logic;
        RXPCSCLKSMPL2   : out    vl_logic;
        RXPCSCLKSMPL3   : out    vl_logic;
        RXUSERCLKOUT0   : out    vl_logic;
        RXUSERCLKOUT1   : out    vl_logic;
        RXUSERCLKOUT2   : out    vl_logic;
        RXUSERCLKOUT3   : out    vl_logic;
        RXVALID0        : out    vl_logic_vector(7 downto 0);
        RXVALID1        : out    vl_logic_vector(7 downto 0);
        RXVALID2        : out    vl_logic_vector(7 downto 0);
        RXVALID3        : out    vl_logic_vector(7 downto 0);
        TSTPATH         : out    vl_logic;
        TSTREFCLKFAB    : out    vl_logic;
        TSTREFCLKOUT    : out    vl_logic;
        TXCTRLACK0      : out    vl_logic;
        TXCTRLACK1      : out    vl_logic;
        TXCTRLACK2      : out    vl_logic;
        TXCTRLACK3      : out    vl_logic;
        TXDATATAP10     : out    vl_logic;
        TXDATATAP11     : out    vl_logic;
        TXDATATAP12     : out    vl_logic;
        TXDATATAP13     : out    vl_logic;
        TXDATATAP20     : out    vl_logic;
        TXDATATAP21     : out    vl_logic;
        TXDATATAP22     : out    vl_logic;
        TXDATATAP23     : out    vl_logic;
        TXN0            : out    vl_logic;
        TXN1            : out    vl_logic;
        TXN2            : out    vl_logic;
        TXN3            : out    vl_logic;
        TXP0            : out    vl_logic;
        TXP1            : out    vl_logic;
        TXP2            : out    vl_logic;
        TXP3            : out    vl_logic;
        TXPCSCLKSMPL0   : out    vl_logic;
        TXPCSCLKSMPL1   : out    vl_logic;
        TXPCSCLKSMPL2   : out    vl_logic;
        TXPCSCLKSMPL3   : out    vl_logic;
        TXUSERCLKOUT0   : out    vl_logic;
        TXUSERCLKOUT1   : out    vl_logic;
        TXUSERCLKOUT2   : out    vl_logic;
        TXUSERCLKOUT3   : out    vl_logic;
        DADDR           : in     vl_logic_vector(15 downto 0);
        DCLK            : in     vl_logic;
        DEN             : in     vl_logic;
        DFETRAINCTRL0   : in     vl_logic;
        DFETRAINCTRL1   : in     vl_logic;
        DFETRAINCTRL2   : in     vl_logic;
        DFETRAINCTRL3   : in     vl_logic;
        DI              : in     vl_logic_vector(15 downto 0);
        DISABLEDRP      : in     vl_logic;
        DWE             : in     vl_logic;
        GTHINIT         : in     vl_logic;
        GTHRESET        : in     vl_logic;
        GTHX2LANE01     : in     vl_logic;
        GTHX2LANE23     : in     vl_logic;
        GTHX4LANE       : in     vl_logic;
        MGMTPCSLANESEL  : in     vl_logic_vector(3 downto 0);
        MGMTPCSMMDADDR  : in     vl_logic_vector(4 downto 0);
        MGMTPCSREGADDR  : in     vl_logic_vector(15 downto 0);
        MGMTPCSREGRD    : in     vl_logic;
        MGMTPCSREGWR    : in     vl_logic;
        MGMTPCSWRDATA   : in     vl_logic_vector(15 downto 0);
        PLLPCSCLKDIV    : in     vl_logic_vector(5 downto 0);
        PLLREFCLKSEL    : in     vl_logic_vector(2 downto 0);
        POWERDOWN0      : in     vl_logic;
        POWERDOWN1      : in     vl_logic;
        POWERDOWN2      : in     vl_logic;
        POWERDOWN3      : in     vl_logic;
        REFCLK          : in     vl_logic;
        RXBUFRESET0     : in     vl_logic;
        RXBUFRESET1     : in     vl_logic;
        RXBUFRESET2     : in     vl_logic;
        RXBUFRESET3     : in     vl_logic;
        RXENCOMMADET0   : in     vl_logic;
        RXENCOMMADET1   : in     vl_logic;
        RXENCOMMADET2   : in     vl_logic;
        RXENCOMMADET3   : in     vl_logic;
        RXN0            : in     vl_logic;
        RXN1            : in     vl_logic;
        RXN2            : in     vl_logic;
        RXN3            : in     vl_logic;
        RXP0            : in     vl_logic;
        RXP1            : in     vl_logic;
        RXP2            : in     vl_logic;
        RXP3            : in     vl_logic;
        RXPOLARITY0     : in     vl_logic;
        RXPOLARITY1     : in     vl_logic;
        RXPOLARITY2     : in     vl_logic;
        RXPOLARITY3     : in     vl_logic;
        RXPOWERDOWN0    : in     vl_logic_vector(1 downto 0);
        RXPOWERDOWN1    : in     vl_logic_vector(1 downto 0);
        RXPOWERDOWN2    : in     vl_logic_vector(1 downto 0);
        RXPOWERDOWN3    : in     vl_logic_vector(1 downto 0);
        RXRATE0         : in     vl_logic_vector(1 downto 0);
        RXRATE1         : in     vl_logic_vector(1 downto 0);
        RXRATE2         : in     vl_logic_vector(1 downto 0);
        RXRATE3         : in     vl_logic_vector(1 downto 0);
        RXSLIP0         : in     vl_logic;
        RXSLIP1         : in     vl_logic;
        RXSLIP2         : in     vl_logic;
        RXSLIP3         : in     vl_logic;
        RXUSERCLKIN0    : in     vl_logic;
        RXUSERCLKIN1    : in     vl_logic;
        RXUSERCLKIN2    : in     vl_logic;
        RXUSERCLKIN3    : in     vl_logic;
        SAMPLERATE0     : in     vl_logic_vector(2 downto 0);
        SAMPLERATE1     : in     vl_logic_vector(2 downto 0);
        SAMPLERATE2     : in     vl_logic_vector(2 downto 0);
        SAMPLERATE3     : in     vl_logic_vector(2 downto 0);
        TXBUFRESET0     : in     vl_logic;
        TXBUFRESET1     : in     vl_logic;
        TXBUFRESET2     : in     vl_logic;
        TXBUFRESET3     : in     vl_logic;
        TXCTRL0         : in     vl_logic_vector(7 downto 0);
        TXCTRL1         : in     vl_logic_vector(7 downto 0);
        TXCTRL2         : in     vl_logic_vector(7 downto 0);
        TXCTRL3         : in     vl_logic_vector(7 downto 0);
        TXDATA0         : in     vl_logic_vector(63 downto 0);
        TXDATA1         : in     vl_logic_vector(63 downto 0);
        TXDATA2         : in     vl_logic_vector(63 downto 0);
        TXDATA3         : in     vl_logic_vector(63 downto 0);
        TXDATAMSB0      : in     vl_logic_vector(7 downto 0);
        TXDATAMSB1      : in     vl_logic_vector(7 downto 0);
        TXDATAMSB2      : in     vl_logic_vector(7 downto 0);
        TXDATAMSB3      : in     vl_logic_vector(7 downto 0);
        TXDEEMPH0       : in     vl_logic;
        TXDEEMPH1       : in     vl_logic;
        TXDEEMPH2       : in     vl_logic;
        TXDEEMPH3       : in     vl_logic;
        TXMARGIN0       : in     vl_logic_vector(2 downto 0);
        TXMARGIN1       : in     vl_logic_vector(2 downto 0);
        TXMARGIN2       : in     vl_logic_vector(2 downto 0);
        TXMARGIN3       : in     vl_logic_vector(2 downto 0);
        TXPOWERDOWN0    : in     vl_logic_vector(1 downto 0);
        TXPOWERDOWN1    : in     vl_logic_vector(1 downto 0);
        TXPOWERDOWN2    : in     vl_logic_vector(1 downto 0);
        TXPOWERDOWN3    : in     vl_logic_vector(1 downto 0);
        TXRATE0         : in     vl_logic_vector(1 downto 0);
        TXRATE1         : in     vl_logic_vector(1 downto 0);
        TXRATE2         : in     vl_logic_vector(1 downto 0);
        TXRATE3         : in     vl_logic_vector(1 downto 0);
        TXUSERCLKIN0    : in     vl_logic;
        TXUSERCLKIN1    : in     vl_logic;
        TXUSERCLKIN2    : in     vl_logic;
        TXUSERCLKIN3    : in     vl_logic
    );
end GTHE1_QUAD;
