`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Kl/9fI6f6n2YUx3zvYiVQ7BbiwnfkQuFj5D0OByRjfB/EH5WBaD6+AM6MwViOr6x
mciiLjaLtUXp4h0VKWZzcqftgkVlB/ePKPUoWHCyFD5RtqTzcA/A0H2pSJYX+VDA
XqkYYDTRXhrriqeJhwVbQlwbRm5OeFCQRZhquyt+exTTlauELt1bMJcOadBut/wQ
`protect END_PROTECTED
