`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43QEIQES4pfOOb9/jLYwYZx/ULqjcfGBsCRDSSztG3ie
BmWgTydVrsrj+mDh6QT/CFwbO//bTYrAlGFyy8KVgpy1/WwvvAGGR5Pi7d7+8BdK
tQjh+BLhpModSqSh2EEXZ9+9OEIJA1UxaNmt/6jeUp+/MsSeyzCBaeepYajo8FU+
WI5RRMZSgJeMwNF+1s7hAU1RZ6FN09B46wG0aYkVJOZrq+4/1PMvVMKk/7Vr/T15
Mt9OHgzIe/3zllu3etJPlRYGYuf/QbTRgK5db8odce9+O/XXr7cw7TdT3gvGYCYd
gjB2p+Kc0Y9Ilj0ANLVPCg==
`protect END_PROTECTED
