`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMtihXKWKwnLQ5Ag/vprdyOwgjgqEIzp1usoiIB4neqO
WsPtOuru+mCMZdlzO/XK6qs1xWSl32yzIjwcIrFlgSTO+1JvvF8DeorO+IpOLNdu
VBlJ9mG60qfXlFjH+0UMI1S3V+eoYS8Vcaw23Qa73f1mvmzKIwJeiEWuq9E0d3Lf
zXhjZDCWQkPWn7kHcj0bUakAXJJO8GT5VleO980ofJapnteMT+qY9vjftPdxUtQ0
BVQJncjkcWtwLzaSKQZvZ5LTHt9678OM6vbt/eh2nbvhiY6HO5ifNIjTZUaWcs32
OkHdPohSY/4m8HRtRIwyhFTWP1J8yUYXxMF9y3EZ0gW6iElzEoezgvgt0DPthZCj
b9IA75r7OiqVNET+aGCjfA==
`protect END_PROTECTED
