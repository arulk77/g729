`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNnYKhWnLYYS7v97APPojcUSZXEHU/coMJp0XLCM03Ow
VmTjG36KE7oyuM/9GTzLl386c+AZkXVBq+dx8z9Z6LxjExu1Udq0BoaF6wOoOTLB
Frqme0ExidqftIGm7RISR0lcp+s+LgyOrsRAxw4DzQbUdS/WGdK5LlUzskCawrxx
LAsRPN0d4/Og672C7O4dgDNPcdKl6IsLf5/v1GuU66LyPp8ccwXkzcfRO8JSq0qQ
MJ1EHd7QkM5eQA2cOuGb52Ktq2si9YJAeBuWZj6mNlr/+4k4qHAW1fbrlRrB9el3
k5HOAProF/Opu2D+OWLMY2Yr/dnpXLpu72hN76TkRAT2CkhtegAqJ0ymCk2V112F
RebNOFzkeT3va/ki78XNHEOHXFEEfhwSvUr29/7cg85G9vF9akO2HJmDxVW2m48Z
ghDRymTx98mJjSkFGpycsYVr76u7Scit4uaSOUsxizTeJcJ1ttm0SgxfZeZ3VrrE
`protect END_PROTECTED
