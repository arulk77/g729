`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43JGp9uez+CKK3sKJInRDCqVt/XF+35MPppFA0zUNXKV
XqBMDa01b3N2qLpAscnqSEhhkabNuhD50Ge47xoTwPsrAcu5Ngt0l2A4qj+dQN7W
WOusF5nwWos900eK7tzIwj4r1SF9fYG/TyaGSS8NpCVHMNSzV/NE5z2IJrNpKCbx
3yVPmhKuNy6/hdJb/P0xz/tdC0pU7PJQwWrVd5mV9vpj++EKKgRrndp62ozE1g/m
RRlsRCiaIWy11C7GeYgkbPvomFnuk6W8DNvp83FhMVU=
`protect END_PROTECTED
