`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOhAIuzvpPoxc2faCq5pWP2Mm4cedC6J5QQw9DKsnBDN
4Kc3cReEHZF4xRfWmwdRw9tFfIhNov1CkDqZ3+hc0drStsxsBymm7c8AOcuaCjkj
LLdN7e2KI5msefrnXJxM4j4CZkOgJoJJrC6Iu+3R9z+BybJgQ6xKTvIG3/4ZiLZr
Z6EIB2bS18DqXewletC97GeRDSlS7yWb0NBx2yxRN7tmuNTI19TD1WNIVj+e2kNC
nzggYUzYfqWvakadDeYYlVO/lRd9klsFAUJwwSzp0hHaBh57Ptjw+s/s6ej7w6op
uOxcHH9C97r3gs/a8irWLVe39NTkqy7ijThkUt7/tiuNeVZuWAEAUPwA7wxB0wUV
4K6i8T5rCbvl32S9jmwFceouAIxha02lvxSwpBunk15RpveVcLFhLaOZh1uRFrad
FkSdTZyZJzl89eMyf5dg/pAlwrkOS7TYGlkarK6t+pz4qWCvimAzTKd1HFXJKsw9
QcheOxL4R+gtFSzU8MENd66NEmzXM+Xj/4PFOoac3alP6OLic83vbFrfatAvL7sa
wU51c9DkZQvV+dT5hc1Ke10EZqKdGtuufjlZL9UdT6mq/tF4IqYm14ZKeTYsMCOO
z51GhcjXn48qpHUX+3uPrA2gPD14qbp10GJlX2euMLLiyo63HlOzdr3GGYZeH1vT
WI3/kxcwHXejW2aoMKlnutN4ztm/r6FjvRVKsFsT8xejLl7tqjV1bd+4IHD7zL2t
CAE+RF1iU0um0X2pTq2gFbcMcJbCGTHibbpfg2DreLATt0dty7LmGDK1emaBKquC
`protect END_PROTECTED
