`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46iRK7/FJaP0tO9eckyrlUM+ZPFaIALPjDNmNWFmIW8G
io9bJW/Z8PNY+jBz8oU28ymNbHJWTBde0VbF8UZZqfBur6lJmNXwyqimrKnSBIrG
H+gxgv9Ab6xsf/OPzqAJf0iqQVeMVoPSd+29d6+Hmvgxp6V0rsoZsp7YUwqOJBX5
MJwLeL0NTOAi9jYKcswElWYbpk9Zb2sy82fzKAOI+NvaVAbE1iFDM7kLW5OoD6H/
fzCYuc/6ZdaeOm/E5hrYAnxla/j2/1s7fpcLMGEVObHfqI/DH5LhCEFkTDQYTzFt
j+FGweHFMbcKn+a91XM18Q==
`protect END_PROTECTED
