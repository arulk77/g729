`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ErQCnae2O7a46wRXcp4+6tTIr+cwHQdQI/UwUTKn93yChRUb2eoO7x+H3u2+sZws
QiZcqOMstHG5NrMUu6DrqBbAyZV3puSw1FrdVZEE/1JCA3N/MoeVkqGEfcuXjWMS
qyBX/i/2HJ7U0nOz+dOPQq+8i0rmlSsEbRrsefZBtP/Lc5JTnbVNb/MYaZZORdlJ
qN54Nzf7OQzpuNbPpYJomAxN0ocDAY3IKLgxBImS6Cj+IU5JKVPZvefFGVJUKVvw
Fwfs0t+i52JSVrUM+EqyLVhr0EpIH49EX8UYJbQ/n7220YN4cGITsJeqv0/9CE/0
hygNoisPZo7RVXAF7rvlQ8zj7n9dTuHvmJujfQs80aaON2ROacoEpRu/IaBPi+rx
d46vNsD83Xz1I424Hgua3ghLNI1GcL80xtZc40ZDIlFVYzYOGL/a3FQQT/mG6uOA
GSmOpuLcbtgUmwlH6JQeOQRNpmL+A9JXt/OqivBNugjsO7uKHoRr0dmp/yMskkpH
qDTE7NoXRWW/7uXQEKF2CPJVkBrgzIFlVCkz/1QJKW7gjzxUpN9eNSQVCfNyXsFf
jdTip1Ia8g5pYg+ie/N4FfmQ+6vU5DB7vLt87cpTs/A7Yijp4fSTd2QWKE8438wV
MwqW2KjLH1SfvOOUo5zV43SxSHqYn8B2mbive+lSWd/Ha0BCaE17dcp/s9jZAZ84
A+/eKdV41i7QN89Lf25Ox1DSQxIEXPJGZrCbFLmkIjgFuHuvS/2AXo4UnT8XPbnF
`protect END_PROTECTED
