`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73Cw6WqXieDdQVTeJxG8oAAxVg81bgph5Lljv/tCSLYWSO
F99QHwc+CNOFmOq4pgIrh6OIGIEZ/veDDtJWudioGfpzLwuQYv+txMyhAVPLv3ow
Cc9CqcOkaZUiwJyths0urzzHxCjry2wa0kLTZoWvjwuHVA6XzBq8C4SkDGvCjQap
7VwwGjEAbixzwOhdDa+GgUh+rTmCSeZbwIrawYPJCTx63qDaRCasd4+YtyEc6jgt
27z6Ww298OQraXpfCv6P/dHhOD1iwdgQZvYHL5mQG3+u3gKVZZLC3bUXe1UIUif8
TSvlhf262xMDMWpZaXN6+w==
`protect END_PROTECTED
