`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFoK+5GlwfXvYLZsIRliPulMLFTTxlcbypp0hFIzY3Hl
bnZ7B9cYjkZc1VSStd9osQVsfGMZoV8/5D6tkmJC199kybFTkPXt1AQlEVIgBekh
QEqLSkCJklUIYzfUn8T1Mw7pVW/QrM7h06m54TZzPfMy/1KJFe9u6IzvTwisYiEo
YmiUBGrJHQfXfvf2F3bccbchaE31V0CrYN6yvX+JAXFYpRtYhGoA87IciCzZac8u
`protect END_PROTECTED
