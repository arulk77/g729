`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
tcUfD2UpXhOd0wpAp1t1MQnank9whNe+MjFHS/fn7WP9oWyeZZ0FwpVBj6vWi0ei
u/4/Pn4/rN0GHVE85M0C2TurhtVp0tKQHTvIqI4/DdRbmTwk7KaFdM8+cAh5Dj2d
`protect END_PROTECTED
