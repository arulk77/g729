`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
kEcT7Y4BO0j8pWo4Nc/720rSdldVGE6mpdJ+9HVWtSPs1KceOvN7ErxDR1nBGGgS
I2yVmyFVam3XgCnxefpnmrkrs8D9dTG7T/1QH5YQ2JXveYIJAjh6h5qrAftQwwDl
VeZgoQH+uZbQENZkFIevhuzFR84vy5bchEij6hTowAuapeVq1EyHaJciOyPTfCtB
AUnVz3ftrmg0hsM0rBctSfxAg+DrnmAYZUnDO6GgZvAeq15X+m+n/XV4pfEGAX7H
yq8pVpaI3Fmh/NkIoBTizr2ODia9bKAJydlACimY22L5UH/B76nAnyyeB4giJ9XC
Q+uF9KX5oidV+bnN8OSbZw==
`protect END_PROTECTED
