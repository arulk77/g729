`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGU6yA1my5dVC4V8qz9pr83W52dRZWHy6141lur5/DOh
WKriqHSYjx4Z5/xiL6oV2EUKR9/54he27+XoYa8OmLzKHNViWL+B7gAIGv5nHUWZ
n7gk0JvNsYrxjWQWCX1WYF40kYouc66Q0QdK0flzkRHlrO8Q+8HIKjiPNx86+jJJ
w/NG1ADSMXPrhbsK9DAgfA==
`protect END_PROTECTED
