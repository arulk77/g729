`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40XM6r28g9drhb0kBIB98PKITZhMGvLwuwkFs+0iegmS
KOao5/Rnx2bJ08NDFqyVGfI+vtPu7jyc9XArWsmDM1hqTmUEzCbAc6LhyCGovPs2
kkCGdQ6j6mj0WH3UqUy+vjdtS1xQzacgWcxOWOQ1fXvwP5HkKHMFCmuZmWTMVNHY
J9wiDXlKYFJo8/hEJSuUN4TxtOht71J0obzByU7qUbbrGqigetK0KquDaeILgtq8
gyxPMfLQMSrCgJkbc531Nn2WvNohvcFjoNyFI1Yw/ImGZEtr8I3GgfB0Ly2VvQSq
QQePPlM5v7BJgzlsawbko2ukMUZ7yf938/87du5rsJsQctGuGQIFFJsAMJOjm95m
bzr6XqOBpTPwbKBFvNARrAY4yGUq+5CauOuc9ogv7qbcAIVaZaI7ZLa/lCsykeL2
sLBOmrGKCgUjQ2OPZM3KHN6+hMd2tvFwcskDtwnqyDlaus4pSJvfa3ZKxhUfsnQF
`protect END_PROTECTED
