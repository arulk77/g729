`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLFdedLsd+8+aMRbeWVfCEQ6NLVmaPP7KrKq+mXGTbrO
yKxLMvlfobu7VAOlzoETHaAl/yblnIDH3YIRSHE88/6N29EcR+0yRms0TFULSJbt
PWm8od7UOF1ae+owkoahUvjq1VjMr6M66j0xLurlPzV0J+7xfhgLcErEdjzbrBNZ
ykEjJ6+FEgX+gzKrTeUw264gcF8bJfTvo8piNc5tTzUfP+8Erkl5SuGBUdm8mXSF
gc2aBP0P8PY5v1mRo0NJnxPu2kWcxqYMMcGkAT9XxUlBabO1S1WkcVmh1NeoEaea
VKQAR/Nx6n87KBa3CXuoLq1O5jdK38zA+9Pc32AFKtnxJaFwDwFg5fVVU3c7lu4j
pAduogu5vyNotA4rZmbTIQshBBRT2PP9H9/R0LhPZ8m/Sgu5l6jBgXZzcPpymtKj
zIbv/RlK9GOqpWJU7J0Dapul7+NcBxhLH7RgYcVeKTO6Pw3NKRqNVAkVdTdi18kA
f7fY2bSLyICzJxWf3YWjlHrJhua8B/IwS0JKPToZQHeVsdFw3zDc9yHvWqE59gXF
`protect END_PROTECTED
