`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJM6UDGOqdDEyN0xsC0Y3Qw8ARYvNFsN5kFc5199nbD6
/B5LrUvoOe/UDZbjl4QA4Am+bbRuGmFYYpNh9rYz6GPAPLSXqhXQ8w0eSEj8ytPX
D9TIO2pL3rfsDCWzUmzrlPN6xRtFk8brZwQfs/scVpxzFYfF+YgFrdt3HGVYFV+W
1M2Eog6Xnt0nzpVarWyPOvgEbQB6v1ITO4/R79tFZNWOA6mKjo+SN/3FGMD9Z9TG
BvnorwB7//Iq4CZDvstftvm7Gx+pGKX/GAepZk4Fp7KZ1yM5R8QJZ4Bdt/zIL9FG
o3Zcrub8xIdlMn/su7lziqdbCzt8dRvPxI83ZJ+nA2024mskRN1mAqLpKGZIJEqM
r9+//oM1bwdL+14PiocG19IvdoIxluV+cxwMdwwHcISVKoM3we0GYlNazffnSDrs
8YgTAstyGFr17/JHY+ms5kjxmI/JLj+aXgp/l0p1NkNfLibXB5+fv7i1qD3SD3Ud
+GUkWcJvtPoOHtvmxt/q+ph744rzvdaO1QOUJeBirj0rPL71w67xyCHmU1aH1I0H
0htuIAsi0hkxvqx739RlC2MpEUxMC1auJiiCvglZZP5PREDUnmfSlkde/02uOVcC
jhyk9EkZfD+9Uwr5PsxGqt11Yk3Zhth9Oaf476Dgg/nJ/9UwIVON74oHT+4R90HL
`protect END_PROTECTED
