`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
SUQtNQTFx8a6VbXbKmpbHrkVFF/L5o3NnZX9X3y8bHCSYeE7GiSytcWrAPwTDNO0
uUaCTyyCXvCDlSoHMy95PzZHpoE0yAPihpGhmYRe/Nk1YDn9x73lsJ4CWiFyx5Cp
b5JisagpcMx0px5EOlXgDl5d+rhrMQUX3OkmmYwMFDlYhh8eXKOADWb/ToBeOPrM
Fa92grFvJXh4teXoZAvat2/Sci7w63Lkq0YBblg0fdZcb1dVW0QMPRQ2/ohaevI7
f8gLTIT81tnhHNyQ6+VVNzAOEgwmOkEqSbAxxvBNcshDbctc00Aq800WxkmqY8FN
5eCs6FC5CMI+IY5rwwe52EH5jKuLwyVjoHJYm2NH+jwKxOAv5IaQDefrnpOXMhVu
s4BDBawxlEM0HIxzvckmOtwtWyqImC1z+HS+KEEnXJ8=
`protect END_PROTECTED
