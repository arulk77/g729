`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePtHMxjDyITrjluUFtnkUbiTcs0aWUABhr70huNsouqK
b8voHsGlCEPVe4O5NwmxO7P5dWEES+lnvvXVS+nsyLF1zRwd7ACMm7SwfPgGDdLG
7H3cPW9J8pMldVmONSQMWUbV0tTiQ1vP9RmZaKrKtobCGpmsYY7ixBLX0gJDc4D4
LfcZTuKfbe7gDQu5TTDY2UxdXDrQ8FI+zTyuAZu1i8D1pkJp0tYHZ9L+J/sVAe1h
xM4bTrExwN6Ugnm+BvI8P9MZ2pIEPSarrwRe2v1uamLEl4nD9nMrEaBnwS5+fx9j
7slfeQVj/qEqz95KdqQTAWo7voxmVCP3gN4NRl5UQ5vZEm6M4z6Omnf73f6ElpKC
cvDKfL00UbBeVvsXIIO/jKHCAmQMYmw0nZMBq875aAud9Y0tatHornxHbqa7v1Q6
j2F+ZRLWRvwnkzVvAyNlFaGJdWaKX3nl79EcHskNK5djV/ze3+VDf7M9S3JSjfLL
w0bEq9+nKEC7uwOoqpmMPJy8n2MP5j8tOUAL14PbvElu4OTDTodlbxKhBJHVV+LZ
kS7H175BaqHCLa7LLPN6y8oCOq06biqlwLRnM2RaT9sk4yZXfKFU0wDDJi7rwrOG
z8jJBLeQHavARIeRsa5ST6sDWYM6L9/eotCndi0eqlDlR2wk9RVD0TyZbkSvjRD9
c8vjxZrWCUH2UYQpLWF/h9PiqjTt+Es8PkTDyrylYtANJhHrV3VELbEmR7PXzAAn
8xaSdefeEb9iAhqX4Nn2uuQ0j3xf78Yv5iysFG1gCICBgSzu9/xkMxS8Zzza6Ren
4ENIh1oBFBhFLL72HJ1mIh1p165k/xyZ3OwjDI2WVuo=
`protect END_PROTECTED
