`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEzA81dEu6pdxIl3S2eDIF4Ni/UEpLGIz0mTGT1omHE4
CtPhtCiLJ9xq9LSg6K8R8J2q702RUZbcd/+QK4tM0O1Fbwp8YZtFQsJ9HkVdp5nP
b0XpBkMEt93LEESbXBbkAgFSAci3xwmD0aYLU+jtyAkAlH37TkHM1zHvFYEs48m7
O5ow+19Ypeei9aze3U27Y9fCUCXQrsktNgoxKy8F43BpOLbsUxVXIdvlmNJbAxzD
sbCOE2YBBLTiE0hEqvOfqw==
`protect END_PROTECTED
