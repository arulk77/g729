`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL8w8VaB9yi9UYkjRD89uy8KMpHyD5EgHqD3AQCTSjtfuC
HpMh5TAahpeDdWgxBFkoff72ATwH272jFdc2a/KyymJkxHZ6Zjnvd8CIc6SM+m0/
qtLY7Tq78058s6YeuusMQyboATZXipWMz1xfcGc7aCRM9IscIt/91ubKlZoEQgAm
PdKgv5ep7snI0nSvWQxuDa11s71MDJCPfrEoMPoSyHC072lilkT725t5HJ7Nmj/w
nNrSTzqcOFW9lBeLv1nzj41chiGoMAji3oWTDFipEchfX4fE99JZMRtkbO/j4yZL
HcyY2nckBH8LUlLyn44XBxzne6YYUgYcM3wORkcpP4Frw3w6COheZd5E6Fi+dpCq
oBhbrQA2xZJzJI/Hwu1nT2H8HBLS9uFnEFQNISrWyZ6RuquFZ2Y5CedYTenL2aga
6iSH6xGzDiyTBpmXyld/+yDRZrZ8IalZKbssSkH+zyVu6R/FC0EUMSpGBws+SSoj
0Kqm5VtqNAwdPZndYKwBbEkSgiPr8O1gLPZhHSPBBaNITpCbIC7WS1hTMW+rCZuz
6BfkA2d8tylckvCaI6SJZ24CuueUb2vFQPD2bKgYUoZdnEIeSXgkZeyFUALFqklQ
MIpqi4/tb+nXNzdYJ4YuuUvBmR25MaamzsgK/Nf3av1Qm+dMNDQ/gr7wplYfWY9P
nF7eBMKNPUcDYr1jLnC3ze88qi5n6fdcNEHWX1CikGjeUqTsSvr3LD0c6DeRQfIs
uxirBm0kuqmQ2yvuvt2eeWMmODOri1nBGvx1QsCMx6vWWONTnk1QanrAhHK4y2TX
NKNlVwPe4yY593KvUIBWwQZ0tG24tWc8tmcWrvV3ZoVZ9t1ShmWARfYo2fTDpyu5
VBqhy3+Z8jar4xC0ctm6mvARpegrKkxkpNBvYm9rjHjHNhN4HQgMo2OhaaBikQrG
ZrrMxOOBUFCwglF51xr78p23MUV/vIImeb4UAnca7oO0RegcDicCP2kSeqLGGhEv
2rg5YFG/G/y2sT1qJ8gjDls6tLE4o4r/3JgwRM62qq3n4LeCAT9ShkO10oi0u+TF
45/JaIGsGlRy5GNiUCtmMlwMs3l/dJWRjER/rBPnf6Jg05NkZSdLDhYpTXoPN4cB
Q54BzP4W/2QYe4ypcrKLa8uYWgvaJu0az8yRc5ZPGUT5PYxxPt4Ofesc87lUSCZn
1tClXuRkJDb81DEp7bomhNBjp2v6a+lK8Rq8ltU64dcRPoxzhnxgFAMis88ZzwV5
gEWUwxT2oa/pYh+AyaAtnlci+cNqx00XBSg8pnLr5amFR1A7Nkc1yD8/tp/I3lmT
dRgz1AYA+n+exmSj9gzF9zo2r5DB9mGtKBKqdcmcLBa/xD/4Fn9rfhMl2qaS2gY9
MoX9UrMMUHaMl8bywX3gMe528cwGCMQNZGB6RCpmAz6kZDRsR4vtQ685Wk7w0cu7
xucH0e3UdNJB6fPavKctgkNeWz18/RNA5LBLa/JJmxChRqbAj/KVbtJ45oRNmfZo
CQmRYZ8wImHr3IlfK9lU7VjE3mTzh+gjIghXCwOKd2WFwwoYtTlICYdJX6GQI0Ib
Gema8yMBDJpJ5OpehxJBDjf34XdLDa+zch3nIDsyEOPTc721/pJ0RmTOO0Z+NPj9
gezTJMM0HNbR9UR4qzNj1R37EiEXZiEIVMuC9O4brdf1q3p7J1TOIyvtzCtJ0Amx
j8l9PUp4f4FSHXr9VagjMXhA9wet5U5YTKK5uVtBMDclRssMDQjKjVbUarGEM2T2
tM3yw0O36wxBRcWrzUol14BCQEv9uPhLiBy3Ue+JLlET1tBij14yOQ06lVFu7V1f
89baWq0Hmxf3AhldV2C42aa2QbBiO7fV/bM483G4UdQJFsiNMpBx+HehlI0/eGjB
S9QHaNxNtXsN3T+XaZ80Y7uQwCObcT3ZX+d+HW+J2Z/qGVBS3dmRZRCQH62FUcVO
zN5+nMJlL5IXomn9LsRwCy8vtXt5EXfmvyOXzbdiZ9vGxRNi50WsZh6n+d//wtRJ
eSY4JntkyOhwAPTzSYoVeeoUxVjviTrIeD/gl112hwB93BWoBfQ9WYZg4oLow1Gu
InjBnooEcmVG8pTHenbQurhoYVZ8FpOSJmKgloZb4Uo+sywxReKZgkwm9kNebvxp
Zx0OtV0NgSMDqLPD7adEx3ZQEeqph+mFMCY05C2RtKE8YSHc7PN+WX3QKjyeySk4
iuvvQqbx1/OS8YTCdbXX8TXZTFh6umMtNxqvKEDvcex5jHbQ67eqAknr6A41UnvB
AodUSqx6BuSWMv53OLVSZg==
`protect END_PROTECTED
