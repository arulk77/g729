`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGPlJjud6Q5WOp4hSuGWyoMBaGRH2wUWQjF7m5Ln+JEQ
r5fuviOMKjdahV3t1TEvHTqWrc6F7oBUls7O+b9AjVe9UYwhgkyE5Xc5+NMO8j/V
B30/LO3aV2NcOVneoYKAUPcf8MQGs/apE2mZ0b4oa1/OMT+5YlaURK4Rp4PkDKWG
LocAzwmoSx5mIrvIif+nrN6cp/t5tZWZNiaoT6kXNMYvKJP2CTX5xDUy6PsvCc2p
PNZh66X035CVqNEOkQcyqC5oheoMiwsjWi5JY53sAvyHYS1own0kxHQ1GzDkS5pr
8yKd192BhuPD/olOpAybkMe0s99XcHrCpxfOPd5ex5sB2qmadGzuRf5ZTQtX4sGe
D4FiMOYDfK8aQV4Kgx+9nDP96foQASVUZGspjLtkPo+scedZTeftaZxoxcXiFR+O
tkC62eWCPxynte/W3glWtVsIOWSKqL4T5s0q2P1mdWIWh0Jdxk6nwr/tvp6X6w+x
dJmfIZIxg2LHF8vwoV8gyGoku9/H9T2SCGxrLHSNrGOx5i6NEIz5vI8zkSVGXPbB
AC49rzipAZ1dJL5+b6XyMe+nWmyyxjUcCNCiF050sqdBP51U840eP63lb2uq58CJ
TW08Hju1TwUvri+yPSqSkj2bhy1XWuLVPdWAtn/+T8QQNrV28m/k9KVxGyPL7T9K
`protect END_PROTECTED
