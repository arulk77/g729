`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48ND3jP46D7/JjCFRdyATgSpy15JdnEmIDLlJyt8BLj0
S27udH/kQkmwbmeTgsxEg11CNu8MW7Kenj2/ahyQTG9sF+3NVDe5P0cVq9Im2Pzi
Br4DS4ghjztrlYud48zPjiYFIxOfh2BRvRGmKiIs7z0hmXJWO7mCIevcOi2HLxGh
OrC2RnUs0grII3Gqgge+Udk462LN/RKVowAr9yrFu1s=
`protect END_PROTECTED
