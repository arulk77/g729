`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN20pqOgovu7UatXM2/ToaH4GfjEFMhV+hLnA03xh/+0
Bhidwd89KqDyKEqL/AGVF6+mm3byQDHCCz88gFU4/Iok9BPAh1dLE6NgMk9C/P3D
4BbDc+FrOZ+cse9WvuVhIdkF7tW9xVDN8wkjDhfhE2apgifzy0vpx3IsXmhBk2x8
0IGRCAts8Pexc6ZJBpW3n2oSPq2NmOz/zoOWvEk3M+uLsZortK3iryh0uL85H1TL
Xr757IjhYE78uwNt/0PBYKpB64INtykUYbHqvMpLw9ZIVV52oAKJB0X7wS3b0fjg
Ds82kPN69ZuFpVR0FgCkyneDRhKoiTVx0KrWXVW+ZHP/iaWVfsMkHQGy4b03dagC
0fuGFH1VUFpm+296b8/MwE0Hlcee0v5jcBbZg05IGQaHfnPXpaXamg9OdGq4r5o/
ARh4BfeSDx9odADt7OQuNdN2FQz2TV92iOhEu0XnINMNhr5XUo/yu80bXqS4xOKh
`protect END_PROTECTED
