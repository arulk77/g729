`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLGVpYuwzRHy6h4UE7zL/INdL09r0oI43TjBUwUs//Fa
oCCNKXRLhfbILm6001wVcWIcufi4I7ga/0gGYh4rqSTc5KpkQDuizAmv/XrB8xQK
MIdWZDWL/OUIHCreslqQS9eOAI6Wlt2k/vi88jZD65C73zCfs7RcVFRuiki/Uobs
rVm8lZ2KD4u38cR2DX3DQnIhbNMXyMZoVUnEkEg4vQrth+Y9eVx3mooSaK8b4Wtj
`protect END_PROTECTED
