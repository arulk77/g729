`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN8UMODUrUoIApZzmQaw5Z7a+HDzQbscZslJuVcaTswCA
UwIVY6cVhzlrtP5lp1YWnf3NrNNSJwM3MrIneYNv3TiBRmkIpHDiIM4n7AhfNRxT
1kwHnU0TKY8+JVz9lpDayzkWe6fQDOFRIbvS8eyuzkpQMT7h/29zxIH6Xm2m0umR
ThX0zpiFU5AxEpMpGWxWS1DUGQ+o3TZVamPYtAlVKn+vQkQ2k/hKLTNSj8lBS6ye
fr/R3kcjs9ucdGciYIkY0xNwo82O2i5cjBFfUK59XPTEJoRDFcNsEGVu2kAThtPo
1j46RYvryFS94abE3/8OcA==
`protect END_PROTECTED
