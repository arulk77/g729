`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wA2BXKyAwziPe3HqzdboA0n/ZJXHnYFc+SYCKWciN0m
jsjiBp5MvhYiS2QfzIOlHFimuSTgqqHYzo1rHh2QC7OCBBaiBJdjj/N+PnfLLCIw
YzLpWAd8zItpAq6wiqhun4gQ6+NGdkH+zEcIsxuv7lQDrznvFUofBdcD+6cie/5G
74YayMKtnB+HCzT/b9fgnrz06u0rogqftVHJy0SVzYYH9yVug2rP63pF0vIgIlMm
4xPS7VEcZi9H4yPG9tACqDbk41hxUDy3yces9i5ssKzi5+tJBl2l2CEDx67lwitW
tdhFYNScRKicPo3Oz6ZYFw==
`protect END_PROTECTED
