`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCUiMdIGP89oDTz+cSmgEHOvWdiMdKG/71D7Li5rRtf4
BcbBCkpFkfVWmQ5yZzX5j2eJ11SErnqE9tWqCPChNR5SHCnZk/Iysy5//Pavbc9M
lau5d+3MCLZz/clR+9llaoawzA8pXm26EpRY4J4f8uyBW5jU0iVaA732V0ywfNup
eL3fvCN01AWf6a1+UiBOUDwpgKihV35hiFqMGzNq7/SSDYR0Obcyvo+FK/hlOF5a
au8PtmUuyl8uoKQf0tDqnTwkP1HC+XcxHAiikSMX7D5+vlVobDui1BROlYN3H45N
3svzA7UGBiyUfiSy7D3Qjon5vFQs87BU6Hjby5HUeEm3kO/0tyqRHP4SVSvZE5vW
`protect END_PROTECTED
