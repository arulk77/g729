`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu471BhlFL/idKVn/7B8B3kur6Lq+N330a78OR3r8x70ut
Sudz0U2/nRMvkHay9RJlXSj+ZIS06d+y6+C/V3YYeEFcBHXer/pdK+Si5tdL3sdn
Znvj/PxkKu12Hxzs4W2RS+NRrw7f6sHt3Mf5P/iiBokbsBjEHtn+1zl+PxXQcJP7
B1P/2IXkgpqqU740G+eP82l8/Bv2G5zgdtDhBbuJaeD1O5tPzLIpQ6e9ZQF0XQ98
m6IFCzhKynGpv2T7w6WBipQz/gzoNB6yJL7Q2EGrccLNm2cyRbIQ7Xm9SzAR3Hpy
Ek6j/CTU0jG6HWVW9/31L/bOCXR6Z2nzsCS6QFM0Pbfi9VUkWtYgSftKoNurmdBJ
YCLEccX+hVxEe07JFXbL4w==
`protect END_PROTECTED
