`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveChAB48ql2othbwjOLoWigBuaEuY1nW/2GvuJCF2lm40
1WXM07huIhVoaE/VQ0ho7PBdICkgipDzOyIvhRX3JsLjykklO35/O/jd5EygoDI6
29pag7b7JvA4DfiV3gvOohaZXc/AZZ52ryzHil7RIGYbpqKWQdmrdXXsX8WLlLI9
FbC9H2L7pPM9LW9o3kj0nK010MeHrCz78iBSQAtBM3WBaRnHKZ/EJyh0C3tmXnJh
8WyVsNGeMy/hpHdOtXekPA==
`protect END_PROTECTED
