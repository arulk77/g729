`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
1FzKTBPmLy7UbepIrsWj9f6Ci/YsLtPZnrsyt2lDTF0eTe+Fk4JOqbjZ2xHR+Pol
vkyar9WePw5zJDGkxy572kraI9bLxAxbRVc6eBn0g0jleuVgAVYZi/a2TVSZgIQR
YaPJ1chez9nRTqsR5ZFXS6XeE24Wl5Lm6RjB/KCV34Lqey8WhOlaNqqCWzN90SgP
uw7mx1EQ/bAxI3zGEHb4Exgx2q0Se1dGyQ5CJ1AWx/tJSjyeqnqrXPS4u5Hr04Ln
IE8CNgtLuttATXaVvqjHJp7JTxfIKGQI1H1wRyU9ZF1qH2AtjVIpvxVHzDt11fLX
9fYop87+4W94hMotUoWgspuMVebCMN/JoYM4Ldme8Jk=
`protect END_PROTECTED
