`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43vPAWdzdggQMqjuUGPf1oUmo2GHUfhZZTEgCWlBjNQr
aHpaPR/L82g8p0Ak3MxXbJvOUox6VlWPVRod8KXXMhREbfncgwfW8I0UJVzKEnIV
T1H7TkPzd/M6Qr2DEkXl+E7K7ac9v8lqpi5dyjDz8RdYb1wClY59LFhjcr5QWpxJ
138xWv1hHpFm83gvU1MazKGfZVvw5bBLKHXCEYisbfxDKCoZiwBQNXEsGDrS31eT
OdH12rSHf4xxLp/w27XTFqiaGpbSCHTHnKuzM4YsSC8Uq3N2dtVU6ehBadTVQFqx
5wBjzxvBRf1QAc7hXifK+umRaUcpwqgG9vQd+U3+FNe24zSc9eKtVx7t3QEI0qHM
bU43/Xd7Y8bEzeAgZdB0Pi1ACOaASnuBIf2r/GUHfgYy3XSBQt0WwscTgOBWnslK
2GJtzXWGPkh9hEiMMDZWBb1mg1HEyr0pFDREkbY2B1yWckAOdTYywmTLl8wS94no
XRtpI+rC5uWndLr6nGyI64B5DjPUaK3uKvlzwirfFL1DHGVD097offJHE9xu/OWA
toNhY8uTRbvCAVuPX2fXvs83eT5BG+rMzkFxCbKIWvnw6RkoTmQFhOVjhYJz9N7m
f86TmGCMD3LCo6VQ6GW9gaeEq3KkzM/bC+TscRHzO6knu6Dve+tVnOyas9Kw+mcM
eVQo27O1flNPZP9x9NJnWu4z+b200g7IF0XSoJafZDU=
`protect END_PROTECTED
