`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4589LT5K85Rg7x1Fi02F7H5IkmxamwAhV1JAYcf3Jaik
9lLHI7x1COJSC2gwfhSmjgp2yHcBa2BsRUN4cE2Qq+r/O/y45+ECTYz/x8GYkLwN
YImybAcpQMEaHBtYtTU+LxxwYtKbovzWmNQbfz7ngOcWvUX/yUA2irAgNsF99htY
69swZ1n6/Lgwm9kgMhfEiqBqdDCItHxRxgqmT+xcFEYZu/eDrGZ74JIjBVuCAz+E
v0PQD7ggewvJISP0KSM0xg==
`protect END_PROTECTED
