`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JYHNhZdpfp5yNRQ7buW+SIzFeFe+wB3GRm/igoy+/ye8vxik2f2inpBHuLi+pZxn
NRYkgvH0U4x+Q7FfUUah9+56Wen08RYhEgBs0d8K6A2ojx6XGWxBi6Po8MCPMep7
ah3EG9wIOkzCS7bx++sbHH6T2g4exG5LGjS7EWNcDVANZp7JFpStNLQm0WUJl7HS
4x8Q3HEEx5ZC0M6sf5qJqqO0FoT1PtV2fvdbJIAlPt1h8jLk78pHglqNSxGGfo09
Pz1ePmNek5sB+VMSz3mbxj8UHHHRv4mqgicNBkh86mQBJAWUgc4O1OJqnDVV1MGo
YPPwPM57UU4eBshQwHo9rYw5YSz+bp6rDxSI5bqpjsQ=
`protect END_PROTECTED
