`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4390Tnwt87jTaudIr7fADeGk9hcC9i8iztPD1BojKYLG
MhfVu4LZ1/Y/3rJ0HCfLmMuZ5r34gYZf1tLRXBIheuayizeQY8lvuJ9NQvuFezHO
70UhZ/ePfrbzO3eOhhGyUoYzmNDiEGMrGtAME8sOdCbq2ALQi5h7cnqzKJRIG8l8
U0ZZqnf6mzcFt56rub4n23h6yca+cP4tk6ktpQ3bnF2DOHlhC/DorvS/2Dad7sDd
uY4w6ZEypWniRrr9u7xkOP2QkvqBZYudXoZBjMHbm3FthutQEI/iyz8cvoGM0o6s
GWizEJkB7LQ2JY8yPxTKbw==
`protect END_PROTECTED
