`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDn9vcMsh7FhMhqXxETDofnIkUDjfhwFj9t5Cmev/f6Y
UnBXNbbXxJfnS0BsteFIoiQgQblfgy28sAoEd9/4oCOiO6NqWiyUFK9+lh/TF8xr
j1hgGOtDonLZyJE6ZOM109fRA5k06VNRAagO2BD17snwFk2SAgep8xPGPJJzick8
w+NR7bpMbAU0sXHPvrZbmzW6CF2f/ciVV9hFtRwLIbU2wwdPxlhM19plSFPMyNV7
rmOrpvf/20h5YjUESUURzljZm31hu1p00EYH/Zqhl5TKuxR4rdDCFZo6YpWHidRS
LdOKqbU+uzaNR2ggTVtUult9fql8oFaBqL0pnH+mzry8RSr59A0O5i4ebzmQ7vnS
wL78SfE8twsoMxFuhB+J1rdRcP1sdqWuVE4du1glqzsUwK65H6HTAIJY5Y8EaxOc
jJzDzkiRkg8rlrIsy2m30NcncibUvbwal/3mQTk/7y8xX1igdpujrslOTw2pnorK
qwesF4oBRuWo8xmi3znNfqjb7OHuyr3WSfi77KDGVGzu5H+UYmU3TOyZCCDAcHD3
hrA5CtD+L3cdIiVEybzKJ5QgLvVOAy5OOoob7QMUBdofHCOvC0J3tQGwrGu2vd3B
G7h5zLeV/P13ym1Km51fk5p7+pr5NK0ptIWQZi7+fdEEM7nvipDREzcZiodmzLpd
pLjyzLIvM1JbDgq8DTUY4YOqL+nZpkfLaSsyXueBeI9SCRFVxGLqbi7ZLtpCgkJW
p54Te6S2aekJy1Pso8MRxROPQy1ak83iyAZco4OkKZLaTLiDcImFLuQMynPrCHvX
0ueODXfRxH8t3KsbtIqWz+wwweXhz0dvAsDR7INp1BPQnXFlqImwZGSDkCdaVsol
twE/aluQuO1VA265PsMJy1Qg8hyv8aMTeNUJjs7jmnMh5h2h4uDLr3dR+yqtgtOc
I7w0/mTF7KJ0mIJrxbxOREe6WtNqqrJ6bvyD21DAFUeT/aOpZWOZSgMbhyBIRYuG
nW3kKFnORfJGFJc9Xp7LpncUfO9eQHuRJTzvzMdY/BLY9MGFB+24B+l7T+HS4oT5
itL5e56K10QZq2zsLPv6c7WfRLJSeJnSdzuv+56m10UM+TwTmGI+zFXkmELDsr/E
507PZd13DC3YeymZQlzOCBhlt6nPmcCTQSNCiXtdsnThcZ9JU57U1978vqYoiSPh
dqqutv6Yq/AjnMVvys5nq4UcL/xWgJrSYkspYN9eg03bENok32eeysK1bJTQ+8BG
CuKOMzNX9ajd/PRf6jORSRrzB8OiA1/Z/hHk2uKtbUXZYDDgxy99llPfjG+4PVun
mUiz5usfQDnOrVfjJhtJFylp5BJfkrtZUQb8oglp/1MY9u2VfeQ3D9CkjpFfHjzT
TuHj4DKjMUqi6eBfIAXsnbVN70cA5PRzZ2hmz3UGS+7UhIU2E/hbUyHAuu7v09Fh
wbkakmMa7WWO6zO0vHGhIFXunqMOvlSfOvpQp/zMg7BxZnCmVlhwCma7pgYZjYBE
pUm9SalPf1wQTjBd7pRL4A0eUddLBB+Y17Ps2p11rbOPaULPbXfYbPbf5taVzrJG
77dQ/xI+I08yPdU6Keidsxuct6nIvO3h9zSlNE1AWW1ePSQvDM9o47F5f6naE/8o
HrZYiOL5kg9EOTSqadnmCymH8uHCODN2rBYOZMTwsnlDIfp28qXYGqAXWtK8Sdqw
sNLtX3W2EzM7/Jl+A5jZPDb5iVnSHyrjgGvQ1gbMrfMac9Geui0OMM4opPqVP8NU
QeF5DkrhdX+wtDBuP/cKXkQb7ldwLFvRThM9Em51vevzSO3epWnM47AMH0I++HmT
SQAI2bTRrIrHOjbBgLxuzPr6JKYusd5uIDLwjYJLd7waCbS8+WN99nFIO+UF9G2o
orFdZxt8ClBMC2f/DxaDqs5MGM9FbU2HgS20pKRLqFaEDzzQO7VLRAGUwYZ3of3J
zwP8dZHLGF6Lwm+9YbjuetwYPR1yGcpPiy/BpFf5f8MVvXTf/rGxVjJ+qRhFmCIk
z8UyMVIPamZelvft72mHNzRO74i85Pd/d1VM4sFpsq2ckSbtFWp5TFGYxrGNh8dW
yiEXYrLMOu+AT/aPcMEUKvL3YWzf61Rd6gh8j25AWoSNTT/8sJojuY76ppcWCmlG
XGwnIky1VLt86FcQUCHzvbDufqxbum1XSbcOKH/Cu0ZMHNHvf7yFnH18A9VgRcMV
9t4lgiMVRPlQyypgj8JzCuDBwDOkXcW5XGXb8EDcYH8Rr4VQMvnXgIJc120s0lU6
Q16vF04HdUJ74Xyy3KMBVMOIRHj+uLsKvG2y5DKEhLvoox0Rx2znRR7HMAmIPzOr
pElQpwTeohZ4U1CZ9fvedK7GWfeWkzIIyFaZR0pTzPp4b43eVFdls0PeirSdsY8U
3ariTV2VW3o+NsACTx2BhjTSee1zlY3j7y84eLb3+yszABbNP7GWwkOXPtYPBJDG
xVdJ29hcQTnZuZ0h7ohI513NMutXUBUSs8hYKHiZeXpBcZa7BNmqqc7dlYzAOE9t
6XyapBA5LKdH0PhuCdbSLTLxKR5FfF8v1qisUORtkCLjvqQ47C2qnJLKka3RUBDp
DxUYQyhyJfPlrIxHJtyWmDyOxZA+rRobexfX20H1Rb2EwcoNxphRVBugP/JjKBKS
i72IwDrb3KO7ckpUuzUT+XlkhZZmVdneAJCPm7B0G6dksSBgHSN/8ix+kDlbAM32
bAM6XGQKdbc/kmtm/yVdnPNeLWQv3iKrU7CkRJydTsDRLfMQNOHafXqPPicYDZZt
QBZ5kAH3GBWg/zjd1mptesZBE6T+S1Ybx+vYN0Jkew/D/mUrUt81wnVl5+FY9Ivm
jOPyaMzaw+7JEaNj0jFR/6he+NwgitEcIUnK5yt+7K3Pm1vE7yAavoVVTK6zrlVw
S/52a5CoSB8Esik3bbXi5x8fCUwlIXSsp4PtumOUSUJWxi+ND9r46eGWRira/oXx
2JynkppYOVy4HymnDB8olAzUu2Uxs8yLaRDyRY9Mq9hRFwA4HN+1GPVE4DoU6KYv
UrK30x6pObmzR3oXnI8EDWy78x4Xp7hQmJ4e+R0yTyMZ8LCH9mj1amE1TSveJVtS
XdCnhrMpHCE+3ulaLglctIVMp3IQK5Z0KwE0Ffc0b4lZpqnq7cXjRBbYsYoH1zTn
bptdMcnDxMOT9nK5iP5rzQQi5ZZP9uXxZpsd6JyNtZycOg5VhkASsBQgSynbvHbo
C2oqx7339lJ4wBxRbImBb0/LPI4x1n8xfFmzStiVcWtdI81+5EQyponA5lIVxX0R
Ymv3y5uWBl0oezAHlFcDFucIDBxh01tfP/j4OlIGwWUEWff5qEJRe3Q/bH/3X9QA
RsFcqHlV2/T2BZDu020m9ngYRDznR9sk47vB98j6VH7zf/yhCgF0+47E7PXYes+H
yQhwg+vmPE9YpszcKrKloZzQoE0Eq1aKjQC3hZcTcKZWL81zcr9zRQ6uXhaW8YmL
lwtEyYhEJ8K4NMjlrrewTCtB8gcONJvgff6eMrJb3xEBkn6sF1deoUTq6O1rNTBg
GcL2wsFJr7BiKtxDG/JibLr+Of86Lpv3BX06Ebe+SE+oH0OVipwrlgjGjX+Jw1ne
m4J0mGfQxH1ENAWO3CRb4UM6jSbM7+/KUNddtiVicDc+jchyqvGtNGupV9bxNygl
`protect END_PROTECTED
