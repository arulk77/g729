`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLmk5FGdAfKVursyAi/bQ9FNdJORP83DpnTxzKTdBjlj
sn8CXQdZhnZAMj5aNPNlE4xGHlu3Wzq8S5l9N8ixQzNiw3O529Y1nzX9fr5upM6J
W1g1Bh7VPYhCbWBKiU/6HrNuCMgoHXWDRcdI7OjhlPfIsm4Rvy5YWdNvVJSBGbXb
yUVybJ8L70EEycz7+cQKEZrv5jkBsmnWRtiftKdZGkPGqWt7ni6lY9+ULjPqr70T
`protect END_PROTECTED
