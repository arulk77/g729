`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL8zIr9rSOWiRbvI/Iu+e3ttRofe3CUHVcafEQXUBQFOww
ycgq4Lh7Z3hRoLC4RUaiPCfXNwdlvCh0rdQeY0ofpn0hv8Z9EcOWYtQn1o9YQt+k
5Dl2RJ3fDBe5uWvQ8DOmMg068+2SHvaOLTLaYUX+wkNWOSdn9KHluxbG4nGudJZU
8CLjKjloshiBcmxTPxw2aVtP3nM3hXHqMe6exr5U5uFLoKGE6h7l2lSCFHFIN6Yy
DaTekwCNGYER90ato6xBJT23fFtqmhUkfX/7HYIttJE=
`protect END_PROTECTED
