`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+SUKroDzkuNB75du13ZAAYizfmgoD+4grciKiLHWkdC
mTmsntNS16iIIzmIPh/HHU5P+1hPv77hB2CV3/Co2voJ01pw+sg4fulh3PUXVkdc
/3DRxRaQ+aaUItc/M8Wv7Nx0GswCAFPtCPQqwTFLyQZsuqbQHL4Awd86jnmX2RT8
/VWSNlt9mtwk4Xy49D31g3ZHHJMOlnyJbcndiXmSCBeZhsU5i2kldvph1scQgkFN
8ddjOv8pljNmap2VNh+xoYYUHwiougOAfdtLV2YYF3ITSz4WwVY3pStV46ufQ9XS
d+F1sjG2FldP6ufFkc1bVysDUYCIgSXqSNk3z1bRmJIRTYfvme1iVCbH026cls+k
a4Xz5z8Kc6XVVXuvSL8kHUtnh3WkXz8sCuIKEara5yrnqs7/lCJSnueKdETVpQ2B
SDWB+lHumKHsyuPHQbUisQ==
`protect END_PROTECTED
