`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
EpivravZpLujpzuwqovyFPHCy5jnn+wCN8yBQb5VwvufiEf8XSKhvF8E6jKLliKp
TEclfBc+rbDzEe3tDJuvvQsQ7vXbbUnUKJTO+Kq9zXB4pvzH0ddZ0ehfTBZGR+ti
5TN7N9KpRPSyqj5hREREuy6fJLVbWsC0AulrC7FnPLQImokWWuh64TGh/uOdRAVM
`protect END_PROTECTED
