`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
a9YB5EKFIlopW+P7fdAw1SWOgwx5lXCW4YXTMHoha1+viMU4vxnZRKRsM3hTco+X
XSbP+OLNR3lKh8/9CjI1r45aGhxsdS8Nq1n7RM8qLndqvdEqVruLASPs7WwOIRrx
vV4QPTQr7z2ruLo6exeRJDXTPLrPbwM45q+amZpos1+Eq5595rpEiuuT9TLnnbvI
i7uWjkHNGps0gBaKrFfERT+TQpsjY68z/mGCcz67bW/sJIVNMD+AXZr2XPN6KrP9
aAZH/dQMfPRmnzIh6W8JX9VUCKY3TsjDeZ68ZTZdVYL2ikB0YGAlV78yHrGiKEUM
48qJ5hsrasO0kG8JIE8e56BTkPXlwsHfZAPoJi4JzQsPo/swLeq1mgENrAQZgE4d
4AFSRJW7cg/aUb5fIBomv1mBmnpNspRQlLByAo5kb6GfYe7G0nN4WaH3I3hgb3Tg
xnvsLoYjbLmf3DLEJqdefq2YeBYo4ToMxpPsc0ALwcFTdEOmGO0qbtuQYJpMlMO5
p/SLUgp8+fmof8IH8amYB73QRP3sM6BnZXEE/GL58Z/yhqkIC4M1MAbiEVT0c6uv
aK6goh9UuHanrtKvtOtXwL3YJtd+US5P71BEh9MXyBSRRxXfXjvm56rNYKhM+bLC
999QiJGY/C4zmUgogj5vkoQ9cVBHgGCd6W04M5eXkA64bF8Mo29DL9wz/JOQ7eJp
hXSkZFBbz0t3LB8O65Ff1LBMUKvB178EKzaqmN8aiZ0n1v/AGCLz5+Njn33GsAN3
rrCb1daDQ9wS4XjNoKzN/CsILLZ/iyTz54H8DB3SdRyVRj27K7/9uh6Fr/KUhvq9
MSWy83U1qeQbHJO1uB7HSd8dwlLoxv5Uk0Vx2rhMpw0Sp0mJEBUIEI3Ky9XQaX6J
WFlXDCPh5p0ijcT2WNcLjie7lIQiip+e1ow7DjRTzPl3lCgyZ4Zp4yG+WxJM9Tba
fATYRzaBlOKvEq3oTTkQoqKaENbQT2Ac7wZRRGSR08k7J9kxYdDla+qVEzyEo+i3
+yg+wCrJGHzw6PE9YGkTV/ar95M7/buGbJ8At/FtZyArIoQhl60SeZsnJEPYobuN
pFKlZVCbRDsVafnhKkMNt+WaaoQ9m2rZDMFS3FRbsOXt0vK2njbAvggoXJYNSItw
YlvTWzruKGwkTa3ItiE4R1EftdTj1BlrIFIBU+bHtQYkKT8Q9iSiBSvmgZgXdOwt
iy3elvaINTg3ztFSCeufPrVE3fy6uv+JmG2f7pDmpFpa8xFl7ZtaVxI3lFNn6SkH
EGRwR4hn5ZCWrhzQ9ZYKgr/zt+ab/4tknGw9Q24HKFKeLmrR0S0bF9yLhf25afAC
pFKE2QKwquUzfwAAR9vcUGi3I9r7xCKNkRCU37LJKK3rKAg6yBStzdclqwPo65BO
GoE/qpY9f7+xRkCaBHjo5ou9U6Fjfo6GvbyqGnAe6kQyWe5pXZV1xCiMXIQX0ixW
QYIR3PLGyneLIeWCnOVAYG4vynTTWWGNNS1gs8BWl81qlDlR7h8NFVBMbZIFIvcW
qT6Nop1KArXwzMLY5SpzVgAs6OmI9IgQdLMQdsZXXXnbYrG+VeYmjq3kNWr5rS+u
ZCywAoJz0bwd6mJ2ZbpGOM4wl9DLZmdowx9CYmQ9H7rR51sVirjnhjtmLzeiS/xB
E5nHIIvx/lTM6bdFN+1cqYYoDeEsjQryRM+9Df9wzkO+UeqXSer2wmUmhImcstLz
eZCsBmDO4eUX26/7+wM9mre8DbXR9NrJ18QkVJ8w7/V0UKyeY1R67Ivrkr7BLbMo
cAmiIESgAun91AZ41pasEkUkiFJWQhIfCyqwTEVCQSs+Wzo6nooxnkcyfhVHUnrY
tvA5W0uQKW0xN31AbdaO/PWjwmnkxPxdHxaS+98KxoL92Wr9yn6Icj2LhVXwqo1+
IGZEWpvjD0PWcisk2++su3ZnpKAmUJ07zddkddZhbBZXaXaiK4MctgBiJ7h7fkag
qJdSn74ai7XSD2ckT2LMTZzHwp4+eciCnhlqR1w1mka5gEBZJTi5KAap8ZVxkHAC
pIG2tlYqN5LnzjsJOFyVMAXXbgRbdeM/43nlP6IdgdlC/YAfRM7Z+VZNiO6DjFnM
uXRQ7/SWBDF7OcATNMSv28ayDe4MZ5ruZHeNOmh8E2FMVstCNMDwwJui5A6G1jxc
vIA4DBHsxHJdfmEYyj3TM2uPXo5JGRyv6uyXQ+POvlEoc+8ooVfxncY1LvqZjpL8
7KKUxI9aUETO9wJEjvRh0duAWDymz8kEFx1X3iUyLge+dAoPzrxk4hGBPoYkG5oF
KzuLm0VUXqDOgha0t0Bs+44dJWdNjciY3N07mpqbUHq33X9gGrcZXpylXg91qY0O
navnvSDGKUOjG64UJrIygHnEHbek7ks0SScOnChiXVjsUMK1drRNUn5vq9BjMFRV
m2IfObFbmSJDMdci7lq3dSMOmY8frBi8na18Hs727U1m8aWXf5VZDO1HmmVmCwPu
Ti5Mv3O03NQuWKWKLnLhlTt/sRPHh6CRuvbUWI3+fog30QeQBKGRjW/x2ZIYtNQl
3lBNLP9zcse+q5fCdOqSTeO/9P144Qs7rDzMOdk5z9IuIS/NZuLzkP++thRqKBqD
Vbu7WflLdssU2xEDVNs0TpmLAudpzQFJvO3Tw3bxHy910LySEESQBQ94/OqtzcCw
PC0qII7L1rc9nWBhHHV6LQjErD/MHbTm2WDJ/z/F8fyf7yyXDfZ7ZJqrUEeHZVt/
k9+N7qjMixGm5F8zKF6saevGGzxz4eUwdHdKVruw4jWV2gBy5DRPy+Zh3fqiUOUC
8C1FwXCrRoPmzq9tVBMsBjyh7SZdLQkEspAL5/WXoMoosXx2s+smYEojg3HGM+wd
GfrNWW/sVgK/UdRvj5yQqc+HJ84kCiORTxfvGUDOy2Q/ICNpBYv4j7xosssdwMNe
NIwJwu5/gw8h0Phaz/IjKttzbzSDbHtPAmkrhGraeU525FS59IbnM8tRs/PCFTw6
9kI+9M3Wf5k5mJxV6rpnjLJc6wO4b94/lBc+yf/t3jE1+WYhQpm9nxXkScK4mGSM
wBbCgaXHfDe7JQN2nzuyggllkD25FwOHH7nHC2f+PDQP6gQ1X9p9mebNNmh/aB8j
AgGftIEYfgN5Oj33Njb7okCzuQR+HFysrR13OR+Vsdo4fydbPLsvts1rF4JcCN8z
`protect END_PROTECTED
