`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEn0f59DS3tVCvBQpB8mlsYXXdc6URk2k5wQOTP8h/cC
dk5wM8t/22tjWa6RFUC6djWogsn2UUdVW5qPwkDY4TBcBy8FP1TphJ3QZzKaScg8
CW3wZ+F0gzsW06A32ypJY6X4dTNV08yuewY9QsM3Y7txdVJpT/k+RmjIsRDpFbNS
48DJ0OgZAwzxGk63uNGSVIvi2putISKJTCrv3JmsK8yge/iCBjTlmbOFbGkgf4oH
rupZw5i09X0/R/CtW2D0JRRTuzZGSPkehuSkIcHOe7MdyW195ebXQQ50OLYWoWCw
4t2p7T5NTIDV93Ev0ZD+yx7xPsXpWTqWbg/RZr1mpAQSsQSaIzLP3en4heW3V9Mk
E1nxyD2T3VIg2kLeV94ODioAc8hIMPW4BSnaszJnQplfQLhcrvhMsWxym8alpZ+i
Mlos9mqzXBsjetK1ZgqiHoUjkli3UjB4KqHEJi87zADB7eAEjn6WezztCUr07eWQ
KIV+tuxAHGnZimBkQJ5KvcfvnoRK3vevrE4QnNvzRaWjzKqoKybpKvDthQ7GLBFy
dTHDieXzz2Txk3IGy9YScegyCOJuvUGHJX9tozpR4OFTTTXElfOMZMcNmeFVLQZz
kyZAYLTWB5+/T2Fh6y9/kus/p/HfJvQutFNawGXierWl0z+zeHnUuglgN3AfFEe9
aSNkQNGa7bKvC68lgtrW3YUgga8fUrA5g51hkvrOF4pUt++Ax6DERJ326w/pWU05
2lO4lWEjhcHRWJIq/Vxhv3e+JXPOR6pBF10fYoyth4akIuzx4N/l4wTTkqm2qV1w
`protect END_PROTECTED
