`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveClR2YP6q0lw9XfxXKqgu7Tvo2N6WjikRIR1ZxxBbTIW
x0eLBezhThYrSfY6BMgd4XJ5MBnUZM/iHOK4ZtQBNt9joUcb7yIPL0FGb4/RzoCk
YJ5ndpwFirFJOd0/aYi5p9R9k3m1D2SrM4rqVHGbneyDBF7DClRzWcQTK1aI9t9v
TD1rod5/XVzBu39cmHSHonyHfigwgGjPAPKzoHFuIEuhMHN8foDq9Qb2A4E76rK8
PLImm1iBYR/gCxun8Mhq5pSk1BVVnU21syeIRcJf2uG3HIhf2AyS3MS1vuB2b8OL
irOGXpePqRwTohdiiNUzuIznqZd+dhTHNHSToMVG/6AJ+/KNtgHhePDOuvlKtHZV
15Dh4+6lBV0De2hj9FvA3ujKw0CK6/hivJql7VdGBZqf3kAZva7MRTnEVLLsWUA9
eVz/xq3vyhqQf+hz/ea/hUhnQZc9ldcqJAv8Mk7PoxDOkAl2ahWaDxeS9MjZkwsH
`protect END_PROTECTED
