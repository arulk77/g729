`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveA1o09Mxr8dmJ4uaF1za/QfEsJ+7pmdSZ6xFJPYVvOev
fTs1OvzLFnU2y8+MmE01TFumBC/Na8qkpJC7ssbccf/kl6NqpYmy1mkJFEPFvEbQ
mEMVu4MiuhFZVUTJQqr+CijaIu7gbwy6T4Bw2CeNB4wGUwwI+21qi6aDK9WfZqYz
VMnuvHd7RW0XsbCZTUpGM+CPn01PwP66ykoYJ3+kI5UlDIGII91wnqcP/Dxl6WMh
KG2PfMPZFkYi/TnujTnvfTVI2ZVK+0a1NpqkGE0AzS0seUmRWWhqQqfp6Y+PnPb3
Zb8j8GSH45/klABeUEBRP0QfynGqEA71CVb0Dh346z3bQmiBgNKkjg4ExprNFdD9
2phWTzowlWKiLf7GaY/psA==
`protect END_PROTECTED
