`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C1YbSFt4XpACehjPMonGB1XMOu+iHwNn4oaLLrEW/jMS
cfAucNE9tX3wnK/JFPZSTKbGt0+fAcfBg24N1k9YimoMGwCIFQ1XWFRLZJ07yzLX
qVU5oYCe/Th83mOz016GebaIqnjnp3FR+ppHryQbmvm2sjlUqq5hee7u3MIbgv/d
V+FNS7UoIbuNgfjohO30P5xm4VC3TZyJandUSqZBykTjWKDyhZrOvUfFLKGRCQxI
ODZrrPpgyxxr0nQ0FolcqluXsizEzbx+6dhDjRGADh6yepC0NZRvDQHHo2hMqcE6
nHpxUC+l3kgatboe/R+X9Q==
`protect END_PROTECTED
