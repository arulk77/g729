`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
5skro/b+6GHEtwSrpmq3ujVNLuu61VyvOwOrvdUT1wiKRWjCAWo7nIrjEQKM+apS
WrJ9KTfzANHeQd4aBP+Rl6vKDKjeHPHU9AHnTHzeJTaC/ZSXWiUFwAfHONyvx+Xy
3eTaq1UqHpWJ3CyKCKRQd00aC9TgKCjyIdO4DjzP70nUwG0nUEGv3caJfEnpL5hr
fN8gOkf/DXefk8XPp8yUDD/cfEzd0owZduuHU0UQZ+VfCmcG/0KpKkxRCDSRxbfV
yoOMgvP8KYL0zCEaU/08nkIe7L+z13H4ucrba5wLGNI=
`protect END_PROTECTED
