`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJwdpJbfRAJL1MmCJbPJz/ZlwreeuzaQ9YsTft/g2TXv
zzDbpSlE4ZtEAMUG6Qq6UFcEWMYwVyKjzc7T9YxwhIyhBz3w6/p808sTj4DPsFsR
GINllSYCo5GMiiXXXo7KmyQKYvTnJmTwZAEnWDD+HFfxwkze9SRlXJdYPz18tM0f
mWI2t8LDFEuoFommgec13QamTa9nPIWIAXHIkjt1FNuNTYpik53/YPeUEcXNdmCi
/6KbPb/71EAbjZ4aq5yvOQRIjEcE7M+GBj7IPAoAGfL2LMjzKyL+OqgWy6Zy4DxL
YuH+oiVqGEZq2/kq8Rk8G9K3fdZYkpsR07WfnEIRyOGDm1CBJIkh/oAe3FKkSd8U
VC+72jC7dPF/1guQ+proibY6EZTMYs0uaJl+N5BlxOtNEDsCLWqhxSMA+NZjvMXT
d4pJp7JqggtUXWC7TbcX39dEE74fW8t9tFPrFwya37Tobyk+U+eVzI2gpINLauUr
ONxJzbjZyB4RiKBpF/Nl49yLVz/UQC+wfVVqwtNNNDPfAuczrTw58B4j7A80RuJv
`protect END_PROTECTED
