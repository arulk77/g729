`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1acxWC0j0Sr/NMdeERtumIfSw7aQYr9j2xOUwwLVF8nyw
l+Za8hTA0EU8ybfXBbRKVkr4FRkZEYTOEh0txvVjnO0dPJo0gHCGhY29UxzHRQS7
xaoAJA8xKGtGCGUacoV5QNeB404DpNQk20fUDulvyYrW5xFp5TI2seaSVXbEomWy
+se8gGWuPoyHj+D+fNoPYExjZasulgbscwd5l3NDLGkbPKJ1zWcdoKoFmWKw8DI7
`protect END_PROTECTED
