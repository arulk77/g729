`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI9c/twzUI4n08vJ6yXxYYGV8rMKu4vT8RZ0yWIWupCT
8H3b7X1cxq3zi7ZVTZCOe4ZlzdeouZ015UF0p5duNUUmIWnI8I+/5+5FmvqNOIAN
QRy7ESUGKTg4VoOon9OSDLA8JF8aukIEFgk3oEUyFLPlpJKYMr32aTmcl8H+SLfd
XjR8tWphR3Moo7JSiLfclhZX5uYFtVHA2a0Rx0WhAh/Mm5DPe8bYg3/mDGYNj5Ik
nC5RORt4nJKRTYUKAs35xQ==
`protect END_PROTECTED
