`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SdOaEAR+MAr6t2MlNI7dTRi4Y6Z9VS3EYTV2Q2bjz5qc
o3zzazn3tcqhUcRJN5hPPTXFF03IVUUjsFa5fX/k/m4nZlETcAyTSpQ8SiC6MyQ2
0mxSTZUDZ8Tep850gbG1JvBeAPScKa3avu/3/CYXIE3rnYHYB97uh1dXlqMnJXAr
Cn32aeEX5uamDMWlLe72NEywZWEds6TFyKClFa8IPlTn0ifvAmWIG5ofkWO2mLKk
cCZif4zkF5E/0O6N8tXDJlIn/s2GH8LdGlbg/pVsTSSDEyl7Xh2RSQswTqJeyXlf
F7JTMSM1DYM2+oUFSjG4snTBoARDG0lxJ+ufYtMBAYnVz2Q3inUQl+HKqNnf3+6x
NypVM5OkmnJmrp0W4eU7M4HOCIspCobD6IpUQszA9p7edJviAh9TKanyo2U458qS
cNdnBrN0AiEZ5vvnEaxrst1Bt4BPngBO0XgzvXben87inVOE+aa1b2HBPXytz2P+
rvD8XFIDOVXdpiXWS+jU9z7UJ1KINfW/+WJ/m/g8zr0SIyiv93ms6zqFhV5kAO0K
sdOxvCCwqZU5VQupEjd9KGKGrlFDzKwV5+SIITYa7uJmaQvnnS0MOKw3Rn6xeEie
jKk963N5sJoFKX/hFImKAHPjDD+iLVyBEAKviFlz7+MSvydA3tSjIHFCBQJo56lr
lz98CptT3RJFkG04y3ARWdxSCbjOMDxEdgXG1p6NdPG7ewIYumh3wT54FralM6GU
/pyDPrOpzFI/AWpzT9cPk6m26XZujjRBftAPyfecYgTDpsmrWkGrHSVRLXzmdC2q
LLJKrJPQnI955T0KfL4Ax1frONgJ09afSJ8THS7Wd04w9SuZlDk598UG1wMnqVAS
PylQhTI1UiDfR8gI+C6actZ5ALMmLnfOdxhQoTHpSV3cljlmTEujgwEakfNq9JHk
7T7UoCTIOLhaTEzcGjs+2sooD3mGzVdtxJ9reN1+v3DnYxg2ps3Mwat66JQvzgn2
pHUc2JPS/P9nhD8NvRHLxLMOLwoDOZQkHzXE6N5UMb8ISjGkMKH5PF8lTxUcfuOb
U/YZtz8pR6RIh+yqtyhP2FvHjOH4h1UYWdAo7fCCVhYBCUQoG9AD79OY8BLeRE3H
dc8bADj3LFirMPbykJCMp6NPlb25FisSxpXa8HOOMiWSCHoDWUgTR1ZmEUxxO9wu
vl8wp0MyTCYL0+rPS9RVlb4BH2BRCAf5c74ywlDn+1oN0vQZy3DF58GEQLu4etaC
lYceVbN5quZ/moscqGO0mvjhSP700PmAE8KrV2f10Bcw8qGLvCViR6qjRDDmbr2k
BQLc6s7/gKIfSJLZc6WQaBdxtHIa4XDyoh/lBy1nMEi4Gpo1JoJpXlU0BUQwNT0X
I3bZbLWEwwjPH1KU33wY2bMwgFyKS5g/wrifRgXWaDXz7P6uH997HHdokEgdg3pn
aXz6Pa12upoHIJxeYAUkzPrNvxaR6wWwHw0vN5IvUufss643FhaWS7XBnKCi5Wdx
oat5CCnffmJa8Bg5l2xadDsoqhELNm0a0AqwZbluvU42UQHyLmUHXnH74kGATDX1
DOTRT6MQZ713abgr2wbrF0qSDHmy7ZqwJSTxkig9rq+2AvYRXNMCLuihiptXHADU
39GtxxZSv2FGdyt6ocnBkW6JiJOvNEf0jeRLhCkd5xWRpIZ7UOYJL15sRV+9D2Tv
gN6mf0frNpTIzIe2ubOm3WHc2s/10IHzjnKHh/j4J3RLB/8MDpxfQIxHfBY8oPzP
0+AUEif8AHkkNObe+WPb7sJiafpvyR7afky606CQyxakfMKOMOrzQhKiLNVGrcTd
43pzU+SKMUtN+7DdtnSgkUq4CIu1QgDK5XXbCxT1Tsvs2KPRgadIdRC7RM83uiWt
m8d2FOapcuWabyVIRBFvjVOnOdOI73jML90JbduwNLDzN3ly/9tQkFWer5RkpQqd
kxkQl/Ks5s+tMr/pRqrtuz1LbRJXymSdTMR0hC8/ibjaGSo/2kLh+HaQOdifP3aO
HAIQSUthw+lM7/e4j6RU5HGdqzKXONRgEHcqfRsuWQ2Ps6R9d6vMHyA7GxgM8FFk
MjOr5lrgZSPk419gIplkUhRXJlOqpSflhfSjSzycIum7BWmvhuken0XYjFtdEcty
jwQGvQT1m3YEYxMGeDcNPo0onmtcPKttx1eRhH00/E7kjzpyOuPYTkaSEaIYHHg0
/YbWbId2a3DgiWh+gwt9gTFVptswfoUw7qvjitGSKk/Dds5Y7wD7AokuW2BIA2f6
ZMH5MYGN3j3r6oABankVLj7yAmxFt93ubVPIS/W6zxKz/LAQP8CdtprSNrynLWLP
gnLO3dssZ41VW2CHGmwUNtkmhNMvPBQn3peVe9QI86qhGJfh9gz6c/vukx4mABuC
oDNRIcs0XDwXkCnCFn7t7SD8at86Ude//KV7K2zQrNlzEuswEu4A6Q3zl0hdgdtD
TT6jmwZBM9A1oHjL9koaq19uorXmsH0OMdz/VgJEfe23KjrE6cHZrCmpZNmGILP+
De4eaxLG9YDiu3ao9lNV5yhHpnqUzZhsLjd+aIAdEFU7GYoaL2wG/zZfIh01e7oJ
9+c3y8w7v0pPWX4QOJROLRVtv9EZoF4JhbuukUwdXRGJibQp2l0/9k2+297qkPY9
YC15W2GRwTYPdw0HRN4wAPn1NJNaKAgleNVVsMfdTlGS+oI9vpY68NKHQAA502et
1K05cGl/EG/srRVV83ixZmI9XjEvuqmJhLtylkUaW9MSW2Ey8pjxGbxes6/V6so+
rkUbZE3RY13M+iBxKvnrZze1kV6hEMelUzNWlXnFYN+Tm+ibKI3H4b5zSQXMKylY
+DUovJIW5jfrZ9DHR0q7zY635uWZmtPZzOmYZ+TjBo11cQFVnJGe0aKnaQFUvfwj
Zw2u7uPx0QBotw55hXcdjyD6OXsZ9tZSXX+8aJ+zQWY2TChuz3eDQXnakD3X2cyT
wqr+Rv8Anfx5T5I49ZOENJOHu1qZ01GLIBuXkr/4AU/GW+DFSU8FqURdfkn6ZUfg
BBX3wHYKg40NRM4CbHApSsY9iXMfgDE2ASzFPxpLg1Qez/AkUsPiEr9k3vZ8HKhc
bf/DuILtNO0apeYsFwZtm9Gy0gqfdOoe1D0YiphVwJSYReTsFkZuRTIiyC0/MqLd
F2vSvO4mLRhB+l8M8PLuDJOVnvToULn7kACwjwJw47DzH223OyatQRN4s9l8ch3j
6f1/3H2Ut/BrHV0HXzo3twYnCoggWjrXnPafStVZRLnr+pqzG/o8qKtAr4K72vgw
s4zpBvoFDwFRSYZjkjR1R8MycgQ91FrcDPiJnba9EdK3XO1OA7LV0nN65KGyVsH1
MiL80E0Uqy2AKb5iHCoy0ZFfnsGWVHDR1QZTGUDzTXISe858nbfJPacDWZpLVOcj
HmwtCr+tucQDhIgdsNHSOoD/Ln/qhd2G85dyIiOGG6pBI7oDNYy3LVgSb5HsIe9N
+pZpF+J5c0NHRjWNxPslkKpgleDU2jYftxHimt4TE11k5+VMzYU+FejVYSWCfOHg
P0s6fQmqz36PPqaHykXLhwXyD4zy1v+QFwvcw0EhDB6t05P5W119K7J/LKxJfT/T
eEP04tIyNMfav1GWaST2gj2HpFMR7p5WqZjFsulh/PjFN6I5bWMWnGrrO5uKCR6E
3gSxH7m6OHR2Bx149N8FOM2ZFbjBBT+McrcZtsAcvTlUbSy/InqkeQt71Wyi9hTH
3LzRREiNWVfZqMxfk3BqbMqZpUUv7x4dLYy2t/5dkLT5w0nu9i2pHoyg87DXnNPf
2WRcvSDYTImYYAAAr0jcoLzH2LixUj4OhQtDws5XhyG4Ghrn1IL/CksfieyoLEpL
dayp9vjq+KJoc8Pg2O0Yiu27GZSs/77ed8D56+qa8g7RrgzmW8hVpzU8GZZXd+y5
g+RoFUuBgyJCyPiWZHv0NBybJx34f9MeSG/FvfKOXOcj9dXpalSOx+jgU+Y/ln+x
HBGukQFQ7hdnKjqR+ClpwHVDwZ6iJ8eOHScXLzu5rbKdLGC+1ARK0uh7fzqVtGc6
h60mNdpe6doD2lE8Y3la0Fsq+vN2dOyVYC0OA6xIezGvFBc+h8hsYOZzYZbnBapw
8wbNdEiGVGpY0PmSHw83MzKCSTR6O5gooABKy6gbcYR9iEnkUy4VN4mY84GCmbRl
kJ4DmBvu6rylfQpQeDdTT3kXO/TG/I3gCwVMG4f/FlrtjPgekH+9Qg0wBjCEaBDh
G0Wafhkie5tSmkvNhcX7vO2oZ8h+0dTSzSOOQA68rOuWEUENHzvm8f/2YvClOc+J
z+7Z2PqO6NCYEQjNVdC8RNOC1fs52GmepP/XKNeuwQuFG8Kfq5b32IxF/9DHVyvo
NZQsw6jEcM4nV2JzhZj1tXA79ugiROr03KuaXaeps93YFamK7J3r0VByA66B3+rv
MXECXh+8D8YofY58goc8WS9FAMsPW3srOsSdb8POQnXm9e0sO5pEf+czjiQqpUSM
wxUkevKNkeOZx1FX+dEVdNcoaHicF5rV9zxSYV5e9SvYFadPSIrzQPxmoQH+edmz
kLkIozmSJvym9AyIAfEtCZ5M5KcjR1K7Ovx4XSejUdahKNrfDY+AYDC7eXk/8bTJ
0M8G0nEG88Irh1Q3QCFdVBCQ6vkj9hqEFl7J10qqKjp04mR1MUJbW9ltqLlHJ86Y
lfeGeYTOJKEVqM9xU+UGBMdNKa6bpKofpYa/wBWIZsccd2XRfX1HKcVxBz2OKIJE
WOxKFXpJcJpdD80mGX85WOP1Xw/xrcHWTcWVARnZTcFooY7WU2s7lfPROdkxA6C/
bZTVaIXgzmGdEBLbHKUwTtlPgBHxfglM8gdJ7UZEj2IeP97EJ5ZTwNWbyZP4oB0A
c2HrbvR8MQv7JXnV2ne6x9Ew5x+yfUtX5Zkmza/ZT2m/GvHZOUtblLSU5sZ+RghA
j9zkasFIgpXsju78H0Sckdzw8KphbJsl/ffEQVNlZnlQtEr+LHgaI8T9pEKS+ATz
rXKssnUCr9ufx8PPOPd9/b9jzuPiIMh5OMaXlteXr7ni1H3i5UPSvZiDBHqxbfLy
Xs/dnU6zzlAHg1wnY/fRkk5m6/Jqpl2xtd9FOZnk2KN3yvrryWtKkZzYDS12Kggq
IaVQS5Gi+R+u8au314jvdeLxZRidqVTpMurkeb0LO2U064HB3j0zIiPa2AIA1d9w
rMKuybWQ8ZPWWwBUPsHEvHPSY3d2S/8bXosKgF08IN9pmp0J9lRjkmMfIrDp16dq
ZsOUHy0Bic74dVtvdwsDwv48nnOPtusvmF44YpQEGK1LN88NbJo7ns4QQVx2wLPK
GJTd+/CVa81xE7B5Dih44kPwKF5U4/SrM7r1qgpTz2M+PwBPELt/BqN9Qha1AqLU
kyelpbaOqOENxEI5+vReLgUNcLrjo6A9kjE7+6mB1Z4e8KvE6zeeSGTMOZlE++Tu
X678gBjDTvVhtqTwNcTzGDuwmfdFof0q9c4nsjt0RxUJM56gk+Xvdr2s0+btaNrO
1YxQsDPFInpEWskwNDb9VB/++dfKKs5ROyGQne3EDJAKDVOZPXeq6aJkUbuwd2SW
FLbCKXDZxg3YSIR4OL+BvD7b3w7gH0xMlYCWFMT/LN8O3cSZKbZkA6DZSEHMwph8
b6TUdPDSvI4guRukRNJZtePclOFhdYHmYfe6jQaVVbtt0BBWZDyco2VZc41l7sZS
rcVy0ZBavphn/BoFOEnaVctx2La5Kka83g3W4fxsOY6v8GKfIF04Oi8T323zgSKY
AFBgA5bnuViREf+vYEUciDr3jakohqOy47bDXEQ6vY5oyYDatk6pkoYumBaxEM7t
pMfVG5KOyWaK8Jvget0M9n5GmuXWIBNjJ4yH8S+3qhwphsD6Ss0F0MRR94TRWbyG
oGBWmX01x8RxWKnSg9KVNpdsvriwVw11a7fNxi6R1uvsE7E7ApoJRbqEYQ+ujZ1W
BZN+lKXPSd+p7lbotcqeEf8hFBLLEWmpJ/Z7p2ts/yvpI4wGG9TwpWQMmma8h5sx
XwW4nfLtrnkaBzfV9zTvctP8Caa7IvlPOqGjc9I0rNIs1IgoaNYZ6g8dNHkyr6rl
ZIZWwjv7Jv17fhTWiGelnbeE1IfjYwI1Mqa9JIFI1UDWbbIqg8bzHuFS/nsulX8u
Oks0NY4oWCCo2HXts4b3EROw4WGblvtCKOKvkjHGo10ddb32mYxDrYWdUkvUNG+i
m2eSON69Ys09k82A5xf/nFJ2aH302nlS865ef3rAg+G92kjScKYox6gxWAIx2TRC
SQ3Q8mqDkFC4lPB2gufdCjjz5A9JiCCXJrIgl9xH5rVubLluiC3xZJON1b+c0Q/C
lZlO824kDwILlUzj9BHKc2sZad3Hi7qlDk2dEX4Htvq78Fs5n7h6BIneZw4nQFK3
Nt+AyLOzSj0BVObyC6OKt4cb6K2WVndheCtwdxtbpY4jGVfDuxhTJmMLJ3s+bNwR
yOp3KqcQvZYwUzC0sM6Oc7ZIw2T+667GcSaFh0Hx+GzXZ486nl4iDqGkJCkmcR/6
PApRJnTLVPyoJftbyOsMp4xoNqqXEZsdE0X5RnVWSnbe6RGajCTsXn+BMmR7Xs5b
yOywybSRHj6m0UBsMSzLkA==
`protect END_PROTECTED
