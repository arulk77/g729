`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEwx5hjjahZENeNKZKK4KkTk7Z4dyL4PTL+OMA57oGs4
4b51208NV0jlX8Y7/HIe1aSkD5ipy1g8sM3BxL/dSKxKJgod36gL3M18l065UnIs
UYhwQl5nRh5iA9fJsT+lEG7MX24KS0Y/IAwbIXAM/kxaEFZojzR+DNX4jMhAgcDg
TsbsVCXLxzO4oATK0e02O4NTu6g7o8KGckHfKmJu9lIwpl8IcZJeM+z2U/kphuLu
`protect END_PROTECTED
