`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42NCQeU213pPIQmcyxrhd5t3q5i0guD+50ChsQbeHRAg
PguT948wfC71kxYmkAFSVsgKs9oPOe/32NmnOHOT5105KDRXrpH60vf2Dd2Sh8iW
p5xOtS68ky7AUFiqphFc5nuocxQniZuT2yF3RE4dIyKedI74Ukj4tXSS4LERVk7I
6e3lRvxjpU6u/seh/P8zBeo+aH+v4TA9hdRq420fOFmFGb3OLE142rZ1ANeMGMra
TOohZObps64kpBC35Bx13k9ysKutvxXezTMz+VIfeNi6NKEc6dAkgO+YtdLIzORH
k9ywWE7ph8URdmiM3FYsig==
`protect END_PROTECTED
