`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2RtTiaLwZbJSuPbraFO4doeXa5xb42B/DEgyviW+vflujQscJZ+WmhdikBpI2F6q
JDPXWSyaHbO2JbJJrvGunLRRAn8as1qv88fpIEDbGat5BJWYhl3FLuEKw1BGewgm
3NnuMuWfpMr6fmM+zVeW445JJ1Pt8hT80N7FYZLgg1CyYuXd4QbQCrntq3ReaIFm
`protect END_PROTECTED
