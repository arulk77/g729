`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG7LHjMpSlm8DSt/EluNXCaM5qQZFdT0+QvkzXLiwYT6
3ThXinbfaXNInVEtZ7ZouGYbvJ7da4+L4cW71bWvQRQT+YneDF1Ur/8SBruXWqyv
VP193SPp12E2U3Z7Oep/HhcRujVz2JUhEBceLrPrzuGkmPXhcpIIM97UU8NsKzH+
PwFqDiKTPiKfQdecZ84IrtubTXFYVN1pX5tSeMzUEaQA+FntBuj/pbU4NV9Z5Etg
/46j9ZXIwCyEObStEktmZJR9YBXtoUvinEsXP6y4A+/Ny3GkobhO0CExg9YKOddT
2knpCOrPZ/epoK0HY2Bgvw==
`protect END_PROTECTED
