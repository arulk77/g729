`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNNn++ohdZtyQ7ti79EOgd3qzVYXivdnRnssBIVXmbY0
3DT6qcA6KJifG+EzwA7WxvR+FZcq3uqhYgmsCBifOv/jCvl/v015TYzf4CJyPvnV
s0Euy68jNE3r19sYcI6f+2VYkTdueNn+wyakbhMD3RWeq+lRq9Oyuoj9366HlJ4V
nwV9Iqa6LvIYxDjWR3k4B2SpJbiSrqh2+aLXbsDRVZ7xsW8YMchWbSJBxAb0uLNO
UjBwkyRbIubGDewwmBXa89jzoEmbXGJdLhW2+jRDaNuWZIJkiO67QFH+Bqncf2XK
q0VmCc/GrlV4OXa+w+k8JlmK46ORBMECYlvbYXhTZboPIZQHSrEhFcvdvUWnb+5M
`protect END_PROTECTED
