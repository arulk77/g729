`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
fH7XSDmiMqLDqISl9EFhEiFu2MBQLf4eu5TiJG8I5qNc6RC08K9dFj22me4wDnyH
l6CYstkMVme4s5x+9dQRoGks887B/EOM1TgzTFgHfoUiFJbIuu+yZ/foo8EmfpG9
45mvUxoj80xLQ3nOLYeVXgjIo4fnXDAs4SbyMFS8jm5dFyxWhzeOllyMwwOCjZjK
2QF2vp/SoQDsbrWdKP6EzJwnCEHQ1FCsZFAPlMUaY7/E3zzST1GGWpSdYd5EeCxK
Zcs7p1qe1vnFHh8tP6jkSAA+rRmwfKAqKS7ksNJRYMo=
`protect END_PROTECTED
