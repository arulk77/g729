`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEJud/7xf4Bjy4YXEse/NWDk3gsbjl53b9ygYb5D/tK+
74h7inDOunOfFXkdZOsuLnrXXYpS64zsopdL1ThWSC7qjyaoqJ3oZGqD8PPcuq75
uW6CRusizlvTjDCZL2lKFsGXvyF3x5MtGqdF0rFCUw46I//GEVnsYJP9V2hMIl9/
pGjMqO5Wgy9h2bLDRnuSJSCBDiShdBGkH2Yr4iniglYTF8eeBqZGLo1By6VhAcTa
WS1WYWTq7hz4s+B1l2VOvdR8ySYHm5ZPn3jn2eKjT1p3g+VDSUsTpebjzZMTeLcR
FPHR7YJvjbNndzyZTX8nst9xnI1l05DRGjjYfTVqAZFtTQQOXv8gjIAmfFD3D69k
i+kLk8IW+uME90GKlprAntV26g4jnE5sm+Xp0P1qwI5g8wzvPsPf3s/Mr0g5Z50i
TzLq9hhsA58e2VL6soifQIF49Dlk5ro3qbw0ELJmoRT+YOjVtmbsF3H2PrfPCg1h
IrLkLcHxgV4cH9Eha+GIyA/U4SQDMMsFFkTaatvxpFzmmzAG9NLRNmDTuwBs1obY
Dv4Vt3N0SZWXdzr7Z4vRa+jOjjEpYJLFquPHeflA749OMnXs7a2iMUm1Ch33XoZv
AjP5W8oBiRsFfhLpONlFOnihMVCKqAnFc9iiID5QxfDRtlXXukUiQNtlKGZ7obUr
`protect END_PROTECTED
