`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBUsZpKAJbs3fwuH2p2ohYL6gco65OrRdcQiyR5mJ5u4
7mPiatDA8tGqB+tZHKEJeJVBIg43RWnhSJjeq3nvkt4ISImOD4Ju4jLRPzshL51F
K9A3DV5RIox0hQo/btMw+tHjDuGTlgSlbMxy0DlqU1s0esVkKRqzfsoD+/bq8022
AWMar/8tGiiqwpFhZbu8vA==
`protect END_PROTECTED
