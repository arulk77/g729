`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
f11uP3tAS38J+2XEq2c6cCF5ACVSaSW3s7Z+xGIF7dKgH94c2RC8kiRfZHDsY0Z5
sSqexiuTFuFAHSB61GQYa9bkfffc+voeDxOOsiY1OdO9iCxJ4Ko0soyxiOBTmQNw
LCZs1NGvB5TbYldQUj7Ygy8AtKoU8w6cpXLNBGYjzt8nkiGBKr1jj0BTQRdjXhRk
`protect END_PROTECTED
