`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAZ+q/W9GLlZJPDQ5TkCDlAonUMfIDxlniIKPeNuHVW9c
UYYV+mm5Z4D9KeI/ZHd8ziqxlCH08/oFUF6Grv3kM5OrXsNkmTdr4DFwWgREOzSV
QLKBeLPR1dcsoLq1H2Ys4IuU+59QKMG6cxWqjtDHJj2+Ju7XZn4GnLuMGubqwIxS
K4VupT+pSucHK9vbsn8s5KYZynwS18aJSi0whR7FzEdRW2FzE7ids9uPTUz/xMeP
4ocZlMGvEHaKvAib5bgAai12nPhhUzvzyqbxTzEdHuEHqYQXTUifXde9YNJIDPpI
DIb5a5JRSlKwyKm6LfEpMGiQJ6kE60Xi59p22y0tjMu3yzLBtLd6E1vcGQtJIaQW
UGudCQjxBhlkPYlPhjimdVO9Xz8je4zAt4EOWDEylwh4yN1YSTh8Zk6eIo76LFAD
oC5y3KMQzxLu4H9CjA6hg11Xr69LkJK1FfOoy/5i8ft5Zfvubfe3gJWVe4MiUk5R
jqW9yjL+lin9y3Qo/h3bVlekE9DB0TAbmF8egEVPVA+IjNhtfZejan0z/5tbSnAa
ExRn1PN6BfqZ76t09Vlg1q9nX4W6JLyN5EqcHfBPgebRnHhfwbtfT5Q3a9rts1IP
Nb3RSwKKxBUlgoLD2E9e4mOEGZOail/VIhBapoCYnXakUpvmxaVe9BZe86+Qe2Bj
1rGueZU083eZvBmvJfToqyORGbUy08CxBKSc8xmf6D42NL0QagpRaIBnTdfNAAJQ
dpcQCzmxAE4OpECsarHzcBnvsPoPR8j9IJgVO6lZ3kirxjCkXH+UnRJw1fzw7CXY
0bqbV/G2cNOX5BldAuS5AUZey6QzR1DiZt6RWa8P783scjsbanFmNj8Pzxc91uM2
C/wrR+Be0pd1st3UWIz2Bcv0i5E5MtpVImVJiozkEYNS4WGhz3esDprOmOD/Wjec
P9CboWeRvBIRe/g9lWjSIc+6olkw9VWfTEUqDZGsoFhzs0Pl2xh1UnQiGSAwnmnB
BDqzoQoThU3TmjpRh0gNN7EmXlxjcjhqtxpjw/JvgtRKInsERN3H9zx4cHzy4wvP
J4KFa6amghlHz/1JdIbU0WzUgC9j9hcuEX2Z/eD9GydmpnqUh7dhmJDCXOa9tLms
axnJ5MOraCdyU7kt3qmADQpuGjs4utl7SHjuiH3ERia1iJgxagVqlASbTysz4SGU
MnMjSfLxjQkk4/isMzvkNS5c9hjbmsEo9MjbXLCu8KUyVbYUU0GQgHtu+xo596ln
2aZahbYyTvzKbtFsDwTtC3Tz2yIp4MFDeH8tsItyj9bLPUu6/8EZLiCbEgJum+D8
mQM/ftUCJxdbbJNPInQZ69KYtTjPOdq+fz8jLMaatzuC6e0+HC5wO02waU0114x3
c5gMF5EO/H1qgfUYOfY9syOrhGXdWzrp5tgLEXeW0kJrTPVTpSMCNbTL6HH308Ge
fiSr04zNGt8cjNpFMmfpdLB7ENleFHID1l+1DJwaJXtFLmr5X4k+oiXOa2oaTgv2
qSM7euAS++FQOc/KYvBoe/dDOQsy5nSpRzmuLfZQqW8dHsR3hR+dJ+GLdP1ENwqv
PNPTiOGzJ2kXEMAyhwjc4nxb81lOixgdyOT7gcHAoXAvUHNR/4X7meWnCcPsucdp
GAyb2PCzere8EJOaedGf9HZs7mfNKN7eipI8MYO9YXnFyxw1Xxk/2c+okaj/R16S
7tZeheOtKjGN/vH1RM/IkkZtQY1ePShUYINNwfTr4IiXAGOzsIWge2fRmJDut+Lc
+d9MbLsJJVUrNW9fTi8L7cS5O8aqX3pSMBmoeHCGMEXexHuQo8Ujqu0eTROxMrNK
BSYpQ+hXrc5O4obuiZEtKpX4C50/kxMu6J9fXsFWm36zVgpUS6apKjttdVQXFhgx
euKHzcQZYcLFRB35GvnZzC1YiKifjTT/NjDJfqXNkblkkiTcIj9woOSP/IsfZ4kp
rZjlJbjq02KW+0DF0z1NdSSAg8WUwxy+iapzan8uiGju/QJlymfbdDhu8rLG7Bsl
+vUVS6mOlQUIcX7LNdaVcAhyHZbgELyTGhVl0+WfAsTFVjud2FIVukUUROKUyKH2
bBXXyCxaB5usHfMxpCmv5GE9MKv/z2KX7jVtFxbo0UXzQM1xj2ni1QUSmJ4j1JX/
w62YQgq08zyZ5CkZ7i3I/VQrbuMH1GPd5687GqFArp/dlQH3KR8gFTElGfxAtdwI
UMrjxuDjb8dsBsv521zYWdDeLIO5ZZCtGHBOYaIANrv4OPJrrnoSkFmK2CC9My3p
2sy5+4UkmLbP1Sj/AYol5G9AXl8ApMRV5A+whOoX7+MxZw7ZFYPrVvJb94OWGY4M
3pVyv67f6kLgP80QGv6cfCI3AFWHiuat+1037OghfZEwVXDfsUSW9UTKGjv/6d/O
zrA/mO30Y+MJC8YmIOM9qDC4zrrFmgJtveDgbnVE/eemFZYTtBiyvVvb87rHLr4B
GXTGbuErngvylf5mPwSPCLQA+yfStn3bQIlUjKDpHXttC22L8H6Lv/f+XWb6Wdyf
5utUNl/JqIa862fej670E4D52bydi9YW8W8TWuLTP7dbIoNgEGDZgMEQQA6gxv1d
IQtTQYntdcTdw2DkJjRKfVADIKxPfzMJZInT1nn1ZT4GMBbH3UnFKyK9bAvmEZGL
bG+syfzKxID0KU+3HWRJ3IG39tRO7lfW0QpOpPEBQmhzYWD8d+DEkOIhuggoGIu3
zl6Z17CxjYWvonx02evkvjtH98JXHH6JDJF2B6Gd93+82NYzln5Qan+cSu9tCbrt
ktQci8to/J8gu4YwHfJ40jAyEJ8SoD8X3PQb4KR2a5bEtQwfV7f4D83BGBX+ZvKm
FL+447ettPYubSBM/yBMlTZypCcDKZ6AjNbI6+DVd4NLv84nsSD247PPMXoBR8Sa
sszQAGDZ47gUjNVR1Yy/53N8MJ2kqMh0OqK6tsLSY1hXgUNx+SDmWfibh+Ov3BIr
8w6OGDywqVC0Zy+kOfiheffe5vdJSrRzJ5T2yAPXMA4VBSG/+UrOG/6nKB3QneKo
ByQl5H0sKSS6lQLUHW+un0ynRFwJaXPUDYGu7G5HfqfoBmR4DdnCPtKGoRaDuA9j
5gFlzOwW8i0UvU1EERhTR0tK97IS9KH4YIoI5OxbVj2GugcHijucfw/CFWj85Y/O
KCi8t2rP25PSo/HkbIxS/DF9nZyZBlrnfbNwYJquXgtkqhhpJleCMMja5hOWtyXT
LlRtE22oRK3HABWXzx7gc7Ua5AmVXb8QMCuhY/GhkM4jlRFJN42G0Z9+9Sk/BomH
IvRv2RaKqxZs2t7PEDD61Ldw+1y392Ec2Q2uULlaToCzHxzmcLHxjyTcbJ+uI2yZ
oWNOuRo8KFzUJ9OPPCwfGw7+/yIbhu8YHVhqgzIC2fiMM3n1q5sROVYnLMnQM8Wx
equ980xdRYWsefv27Jg08Agbh6YmfkGhbD7mtoo7b2jwpWfthZpqDzOdg9Tkicv6
`protect END_PROTECTED
