`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJi+VQrgWuEmeEWciFv4LjfY2LXydxUxqnLlTFypx7GK
+wtgt55g9NWg8cdDXGw4LpcPcoEdbKpc84xIqSNp0nFQ2RlYMcHCymhXQ70jJ3E9
Yh5otWgCYKsVU2cSpxdXfNT3g6LcHnHJOsyNfpv8l52tlXFJGhNBfRZ37BdTIgn5
bGEUAwAUD/kPDnXjZpZvBVLjDcOZWgFHtO7trCS8LZjQMlKSqoF4o/PefimCtBri
ru7e5396KAokKqGRkATQ6ManykGMemwNKPNwQQrt3QKJ7a6glLm5K5dn3Ca4zo7v
osZVpn7a8wWI5Tw59cVymOCwKbtihXeYp3oAoW3BspRgzC+Be4QaoW1LytpzfLur
m3Xbwr+U/teom5x3sQPR1Hw+TxaoysI5det3gEhrDt8254KtWyKO8ciAGfNO6ntM
J2siRfqvokmuisWmSwovApW8OB16Kjsc2wLFliBv0UW6hXqTbfrmsEPHWGWefEPM
mcxQBNGphAZm+Zu3vcPqvYmK/gQl7G8pJVwsRAhQVxTqNUQL/nvZJnb7B4f1zqdW
rpTzJAS5cQ64t2Qw7vlg4rlItMlvXvHLCvsGcJYggyPX4KEA/+kRjUc8nZqWi+AN
NsYgeIuWTXh7ZMUnfXqbN1BNb8J6u+QdRCpU/+ONQUT++Xz1nwXvhR0OEM51T8/r
k1ONkcorhK4akUioIn9WIyHPP2LkZUwYzeDQKtjLWgGuFsAO4uhp1yrCMlQfRC9J
MwMy0EtlLQ5kSwNJa8arLtb1B5TdwE15RoUmWrLjAc8GiJz1TGXmWA8kiuRW1jyv
hgWSQ78SC3e9WOyDH6dPaS3M4sNzd9f7W6CTbfvuNLUfj1JmPR3PYgx+CeCsCxIz
lSQ2/eHPVmwiP9X4N5lbYiZh3D7O41lajrsgaSeNz2t7WZP2lo+WOnVHBuzlJtbo
kBk2mXG5KWMM5uLVZW3YwtNuAdNuQceNmXrRgQsKqQvldPFspI9w4ztPKLxTfMvT
y21QZ4aBQvp45w0batkbPh/Jn1ne8NQx3x+4oWkMb9sHMPa6YP2eHt2EZXsjedmK
irQxQWIRmh29nj3aVh1vKHsVNCqIgGDOsNpMZVuVxZdEgUx8zBBFY8pCmm40Fdte
sPBmVicQxktRgz4o5MNe5t1i+h8NNisRygi6pLEaftwFRC6JOQNsu8vW+5zjl7cq
MnLi0T5/4qkD6uVKni25xsN+nH2qBEoBbuAHYwUwRFgDtRwk71IenSOV27xtyH0f
JK/NnqcSjFAglrnRzV7L2r0dsOOdBUldSdwRro2TqTaVktFqw1vq20cEPoZVwCr1
iVeBOWf6lZGT8LElTDfSpo45jTUI8leE667oyuZkPFJrXCZKKpmAVpokWKB27NdE
pXTEMJNYcPUkXHdd7Bt2ZnnrAasLvb8SRwjcHP9oNuzG9Ma+iKEuz9iD/l0a98JQ
0wZhJIwn38fr6oH5E9OICUgCN78I6HkcLPmjHglP3azq2YrZ2W5pTsn+dm4+KaEA
5GbYD9+ItcJVqyZ94zSFgGsVnRHf0MK4QMlcplGIlw3W8iMsb6leD8Cv71qukk8K
kYhNnijt31qGG9hj/TTiF6oYxHOabfErJhClvqiyNqUkBtgU8EHPqAlJrAkvmPT2
nvFv7kqUuWRFxbqxcwCcKH29c92jYG+GdtkBKWa0B11v4AvgjxGruAlAcaTZaK/1
lgBti7JgYQaiEx61MiF72DDX66bRCG22NlE1XnyegH5JQvGOMIvareEG7dKBUlXd
D4mBC8tRmklc/Tu5TpkZJuINKHtVdpMSN5WZ3I1L6viDX0btOadVC8wHAmbfFkBk
xmKrOABV5hXs7HDKcoEKSktd4D9r/OkLT4z1SCfJO94LlNLMeevdel6BpSmWQBVr
7YycB9pBbaoMK6CltdE6ONxwcNCQE55Ky8hSxDOAF1bxc6ugeJSRYj+vsz6vfXu8
dkJ67g7/ZnQGbKrhF+mr5MNii/PFpovhBz7bXO2dm1/alA/FIrEZWybmkbG+PIo8
lFRbNA9uFbWhdK6fmm/mlUo0JNPGBmuzGt5UxDw+cj1C7K/27sG32rlzJL70Zw6m
TxdTkytv7FvYjmno4qIzOxLf0rgd0fJ4d3C7sM7xozqRS0NnxIxUrExE+Mf0w7YN
HYfwae9cRbMlfJ5bxx/97YIGAJwUGrJiHDD8yjLqo9y+nG79JdF9wjyzIb/C9Gid
NP0gCmjyKlrLfdrbOIfGkVIxgK8QbFX+oeTf02D3WInE5Hz33weV0mKSorLFJS3h
TNqk4u3LYkjcAKO85a7z1cqKIvyJMms0OLhGKc0DKde6am8XnMM4H8Z1doxM1baI
RliWqvuOx9JQlmQ9bQnKqIbtk4TRDnDqslCzlPp4mtuk2/pkt+d+ZBVAxoXD/OiK
nVjz34ME2qoSZr2SQThAjOZJMW0stxlWAmoBXhtEJkur0xjEOMn7y/7dsP9NqiBx
WKZa+TP3w3zTk0gmGXM4fRis//xHuBBQ82ZXL2eDd/BmTPLmsuMEfF3hPi7JW13C
l6pbirsky9xgNueG1aeYfTyzQfxAibvwtqtCciJbXMq9VvYd5GVrrGRIqCrShSLI
aDrK1kXI0rJWCW0kGI59FsYT2CU19BQfuCulXo9P6ARHVplbp8CGs9BM/P7C2sDg
vaUp7WVqehN1lTytbEUpGf1qOhZyJHr5lCv4ftBzrWgCgghdRUFkZWgWdTXLpL+s
KbgK+E4BBAPZSSgywb4yFV+r20Yz+Ad57yeTbI4Sd3MLZ65jUwc4sOWMfeWxN4Qx
CVCVlu5vMyYOG9mDo1wl56DLsT5mwyLVxuRWTWxRyEawoaEEQeLzJZaHdoMxICUU
N2mjBTLQSQrXWKQ1OABGmojUATEdP/JaNR08fyuRKChEXeH9iWSAUZlapY6Ytw69
vPw/BNJtNoEXIKR+d0b8foQwLN3z24G4OfYJ7/UscVLrX0z8i/tIYOGikwduZpP0
JpfaDITtqANlSGnaif06+GoxexwX7YHO4SsprUe7wvfpL2B2UFuFjj5zNR78WRVW
Se0n7onSxkwUQIwHOwVHyOPiEXLO7of0EqqW62F6W9Z9B+aamCQBaZ6LqA4nzY3G
ys6SCO1T1i2bZtA+5Ed0fN3A4wl5Ie4yBkLXGBJAl/StDAwsniQWmkoyU2Czcj3p
NE1ZIxfiLVAo+fnHXpikxGymVLMYS7k2SNKZkMEa4GHHIwcVclI1cFSHaCkg1SdT
AWGkWxkTLJ2i9Azgtq2KDHISepBdlTg3FqYCkIF5vPGT7NgryoEECeXurr4QAaHy
pIxCuOM0CE0C5uc5hx/Xa6xXDj/UpmojaWnV1ZxwVCpy7lvW1voFk6moAv3jUIvk
ZEqu/Vm8Mt71KIgp3bbr8raae4bd0y+zP12d+5AuXV0P8cGa/EaegLH0rnrYVF2+
Wm1URi0AQkUKtjb89NZqxU8798s9A8TRz4q+xKc8/UTC2sEPzPXlSZkdY/LLBSo3
n7DM0EwWbzAXSkMNNd08+3yScrUibingohfo+0wN/SBRMy+7tRoN5AJEANT3x4u+
XKZ6SE1Lebx5ODqV9Flhk46bYYsBg+bz69yzKxKkxy77juc8TS/zFYLqKpFGOWhc
EruNRC8mERfeoA4ltjlyhwosGnTiYfR+u2GgOSaKtvZyU8BrDWfBUEcrZ+/OImNm
btPIwfa03VVrhDxudpyFkLingQpfgjVpyiIu59c1LLFaavK8KJ6AsKnpt2CZWABd
l2W1FELrOwiRRi+xFOeyWTmgmwrBMLjbeTgdFRqEmCLoVrgmvkylakmvEd5Hm2QW
9jk2tsrnl2CSNo4iYw5y1owOtjDLllNB82x1XKINqxYn8kB4opl1mRwjurJoKByQ
Nh4xsA6T/+wV/2cxJU5FhMOIQPqzXzz+7RoWzoTONJhbdEcaREw9tPwgbRK6XdZw
1aE4H1Rd78Cbe4yQRTUoUvv2qI6KfqC20cuUmTS307Hqga9UB4sEjtvlxyeA5trN
I4AUjb2RqNTpuL9WvwM91TW0BgTdP0PUglSt8votUdA5n+VtgFM2sbOlk0h4C9hC
Tk2A4RWCyBv+iF/psD2lh9hU5UZdpssITfuIul9aZ45Be3Xw7ufbP5Z1C7Fpt/fh
tMuyn75ivZc5cIqsM9fc785HEG687KrPOC6/77XimhmDW1pxc9AJdh3cWtw4LfuD
Nrcu/pxqhOeZh1op1Eu3e01U7b0KAGUoEGuNeTkGh9qiOKOEsS6s5mqnOuBYFDrx
JOpFtZoNrXfz37BHIGeD1cN6EdVJrwcNRBToX6Sd4FVfonOp7R6NglcfXmyDqQDr
9+WCQ3TMC5BgLiYRQs4O3Z+NmRnhYpQOPMFGfdv6V2KbcVdr2PanSpL83hoqK7u1
wWWwPfzEJFlOELkHaDaaJGuwHGxr86e8+fWkbyRCxtNDw9ImGneiYzEIHmV30HsX
Tq7mCyQ/qmrLNaz0o4PKehmsTDXG9fI1G51tkUGijoYfmm64V3NKyXqkGBM0H9mk
yg5qygXzXw2sNCImDBO/I+pc6OEotBQclt9jaGZ3o9sPsMDnLykAp/zNbiaDJLdm
3u9OUd4XAmphMoHNkHb1aatdTaJ5N8MFkYLhKQnsWWO7+mmSIOB9GPkblU9Qqknz
QMfZm2bDBZwO1mThTc21GcT0UCVPx+y8hOttQaM7FotcMTjf0n3FzCMK14a42MqG
64RWvEJhyA9G38ISR4kpoc18NjSaUXeAMDinUpVambe4qDS6ce9GEh84n6forsyJ
dLR+1vgFm3z9Wy5vMvrMiBRQqy8YuVkEOty6fI+qlczadjJHR3bElutNYOi0iY7h
Y0ldAo3sdy4CPnmro3v3I43/qHTMMpBZ+x2vCiuzZWpaZ0uzcYwXJCM69aqnx0yw
UITBuoKt1ROsWmZ0vcTnNqisxKdUJtSZohMZwoL3lcP7wmSXEof70uCulVFsYpue
s5yAO/m9mSY5YADtPKf49iM64fKbbN/xNnF9yOt3Q/JFeU5+AsAiZ7g3UVtGTRru
QcJBgcBuzo03THNG72FrNKvaPy+aP9gDAxsnTGD0xEOU6WLFzU2JHGNx3mOvPwpi
n0sGesXE881mMM408Q36kKfbkbogef4Se90bML1+fy91ufEB/x7v7T0bHVWmHWd5
q9kofVOBm+45hA7uEd86j/OUS2jrbbkW+J/+nQL83obDmo7NjlpYaJNr+/Ei/c25
c2ZK45Iht1guYFZXLqeKZQJcmU9oPDJtbBlfOVJrkOPNCJc8nEKjQ7Xak/fYmx6r
xodQ0tun85EMRjUg818lkKYEUDLJozRMbYktBmV7DZTGdXoiKzp2hisIYU2broYn
E0UBGqJ7uythPJqWObT50NK5qJAdrhwrhlUbbkTu2WfLWV/+2rNz6AOAuc1qsyPb
xeY3a4NvugNOkq1NQmP/JkVRKVpBUnn1IuiPMnIH7UwJUPgq96PP6+AEWWM3NVaS
smr+eRATkU8sodYXHT8nssqItg/kf+EMRUxTUs7q26xYbtyLEpGhrtruFnFCSTG3
3wqVCSVh53SR04uow7LK1WrHbhEkR9pZLa41YgWNg/v3jeFmVBV1Cl4USw/3y2oe
+C8SzIOWIc+3/fSo3lgFvNLUxb3I2ORyxYCID2fLCKdxRIvrI+pYlLx9kuKbKRA1
1JLhE00S9nO1BeC80vewEYqPUKPl6axa1Gd0YOI+oWwW29kWs1VRgsG0HAtIjXmz
TsvnUT8Vce9Ukl1ILdiuPYXIUqTpbVgx5EXuhPMwHVvPVtu1DJoTtq9ajmjrAFNw
Dfgp8tD4oaUIIdLN5dna2+ur57SbVac3UI1bbfkDz3lQzNd9FV+Zc8icU3h9f06l
P5NXy1oNFbBIEtLa4ulkNKL5obWfcMmkcmYvqJsow7PCWjf+bKveUB4t7OK5+Knz
VPUsYv4SRT8lpZoCigCqUbYrFSYGSrl7xdkNh1djhcYTUVtfbOAwskEeq3CTN7ff
pLFjn2u2Vn8Y4QL2Y/xBrZoENPFB/jlEE1rxXohjC7EIAwg8HXEO7zNr9SudWnou
8TynA4h1GYgZejYmwWABUUtvVVPDlmq5qse9ogBksbRpiU0L4Fd03E3BO38rEWG7
bIHojaAvetyRkojdQ/VhI9W2NNBcFALJ+06VegjJMMXkvS95i1cSXYDchFaHxbt7
XH2Abexdow0szB81MA+r7YFVYNXyQIhtJiARF+ZN2hKd43e+DB3xLicJuxMxZE2Z
rxNlrRfuc29zeTI4zbkBKq8eFi/+42XKYDV6rFRZ+WkAb0BXqRwa5Bo4JURci/pR
GoOeEUSawJcTsK03dXeNMdGVGkyaXVpr4j6N8j8CPthIdk7Ooi8RkjHf64iY206R
bPowGgkNhl86ohBMI1J2H2VzQqX/n3gmTVkPQxTEwg4kmEmM0HJXOLmqHF4VPM0j
vWT9GmUVoclaZgpkJbm42uXC3h62uSxtEnbZ9qluM9h09bu5R0fkImiCEAsoxq8h
+knjhTacuF1+oqZJtkNj8ow2b3H+mDFDFLuiRVVcGO29E27kjxTpupELWU1O2ayM
+3KkTjCBY/Hi5To42zMwFqr0B2AX1HlHoKGg7rImzzc1ZBYpC9v1ZP2ZaJwH85gd
gaOpijjtGl7M1o9gcWBuBaIxp9j7cCSp2H8zsMSBxLIyHnBzZEuAXuFsTUnrdXnD
lzGIlwqqNWQSp3bLwBiZyvySRsyR1KHw6I5F4My8PSg7A716p805tthAgN3Zpyg8
Mo/Z24BWDw1TLEzZeeITtihkwZ2avTUjExLTeoi5IzzMO5PlJqygRyk2pI/1nHKz
+elOMwboy+FxmyxNQG+5jXOHQ53JsdZkVkww7HIAzRcDbZ8CnzVPtTL79aHMFjBA
5kM492u9c4a9pjgYYs8lRO6/b8cyaypZ7QSgCClzp69+Cap4K+DK2IT5r1IT2Wbs
vRDL5rDKiTjsz7fQ8wZXo07V+uBkD9QmCkIibXamJ4Vb2EyvjhdmHZgMt2CqKAXL
+lBzkV3vMzi/wEVncS/Vrda66SwxAxqBpxy3NzV/3QDtGoHgfuo2YDHpcB7uejWL
EO7apQYn8HUOskd5uk0IyouFlPlhZq3hTZXmXYrXgwtTF3Z8eOZEDSuTUfENo4g1
zl1CSa4ha1vXfxUxdVfurXCHURmYgxE1nrIojSsjDCXwM1qZ4tcBvba0VAn2ZT7W
mtEzH8f5+HAeGHm7m5hwKTrZzI3GvefyWfoMzlv/2Za2Pdi3SiumfXnlwGzQHsFI
eiJmiBjcDfEAEV9mCsj8VPavu2naqfZMuidPhz64oVrbuXCsbivVAEC870AypgJn
ZB/WE++r3hHwL6WvfT5WTYUEZDY0PISSHuEVWC3YvtM5SoqaY6lslQbKoA7CUnlX
YtMAIRrhsVV5MDcUBeS72wn+FXIIZBpHJsSqHdrYhlmN7DVY+JKY5//2A/s3ZVNS
xMIzQX2DTqL7dfh9zS+S6rTXNsF9B6ykBoU+DyZTr03jjWM4Pcri+7U8QxC3cX5n
oF6uQ/fL/rAKewKRXHnVpUKBMsE/P/seXButcaCzcjM+cq7OYt7gsUTUinRGi7DG
DahcS33n3NlpsT4ahV3y8YhXdVej4jHr2fyTeXAsKpqZCb3KgcD/HoTYmifrCycr
dz+34LTYzwYnSTVTkQLTZf4E/KZroPuO4LuRyPbjVcH56ICDs8sIiUDWTRfxD9B/
+0aaHjyMoMDU5ngvgrb6KUHz8pBVPfNR26X2OsOtvbUkcJrZenPgORUSILOMqWuq
ngX2+WWMfH/9uzFJkVqoMq5NCYl+5wZTIFTvqFNkxu8TksHYn2CyVIwbH9aAAI4/
oGtCFaAmkdOzL3lgLj9/UAWWpaP+bW2EIWrMPRl3jbbhp1ucBFjHmDLqxgAq6Mgb
dOdrEAevr/EwJPNRLkd+h1sqa0SOqHz6SCn6k85t8PcuHa+MQMWT3GiGTAPCFixW
II1V3e1v1JksYkOxGh1ooSw9kwJjSKf9ptq3CmB3zkRH4HCiP5jXMxRpwek0iD9S
RmdhL07gI/b7in+Ao+MOs4Zu5YNrYJSWT3NmeCS80+rTgzeSyuKkkuVk4tJOKGUe
9LsA1Qz/LvL7lQSPhpr9a9dDSVobGHg1iS3OYJHKNDCAcqXGLHpwb0ZDEiSXG2+W
SYUPcmaMGDgueUW+4SjRtXDsOOjgPPGRnEiAl7UDYHHcUxZj+f40+9nS/AMZhCII
zK0Ls1wh9RiSp5J75q4dcqrVXpr7ifWPlrh7sn4MI77oDRVRTAiQYnPaBCvuO3SI
XXW8+iSys+snQiXO17YINPEIrn3gSxPRXlFmFy1p10AIgfSsiPVQrVgt0lkbitDN
M0Svm1AhxniWAT0Qw8qeoE+qikbpSD6xkk3SVbdqjNnbtiGUUYNboN8EnHs+WWqw
ShCc29bJXM0NX9CKhZTr/cPE8f5CsLY2Ao4B2jgTEiDGyC8dDekPgTkvuCvgwrRs
zSTSdEJir0SSSydDhCgE7b1FDOOEXcjIon7fTwDWAU1XbO3NfDCUEBfV19+LKUTY
fa72aeaWKE7B/DwvN3SrbleXVEiJBgfThluEL1NJs4xyjAMFGIC0FqKmzFzmANhR
nqBx1PqBDLzdusWJBSSKtt87RAsU7pYghZm4lTYhH4TsNNHO8NbHTI9yid1hKdy2
q4XTP6PzSbL54mlU0r29+qEkJ+YDmN+xJN2vQmdkwe9syCOByy/vS8u225u/GaEM
p7qwyRrLhePmkyAEBSxy07KHgOPj8b4ZlIFnPssoKvM174vn33kcCACKwuf7Kpuq
JwRe36TnETPgCxfUAqJUXUawv6l+mMN4iV2nB5RxQPBIPKiTkfDqi52VwSm7fxpt
oXfsmmX6kV9gjRIciGBXTeivko1zMpOGpyUXUaQPUSC0BrjI/GbRro98uRL2RYSN
qRnP4tL6rA2OG7Sj0clW35hpz/uMwBdR/QN9DIgIC51lPWcj3OtbNPNnCEkIC17S
zc2AuKVpeXKeKSxapdYKiXO7oJeQbaTyIofL4CUUlofYSSqq4yHm2fDlH/OPnfvS
kW+41AlxmBfA9/LkjHEIJgt41hdhFJ/TyW5wSUyWuB0x5N/krvmN1gfDkTQnJK49
Y0+Os+qYEt+K2QXw7J/f7k8s0I3IWZ1TPjP0LUY1CLJw7pKed/hsWAxaKjvGLWQj
/BfavrB2BLrR1zbVuMyYTIWGFzFUMbJkVDTn16xYotjA4BExHlf81CeQ3bhys1gv
eMw1MGIg1phYiD4zvZ6dMLu9FGCFCZfm6BUVH/5KMlPyYQRV7GeQ1lbEMm8T+2kA
7ZOCvoufM0BeeWkU9UePsE6FJDFa6ZaFq3hd8w55OVDiBZuyjy7dQbGfys6NeEhg
I4B6A4SHj3Xwh1ozieafF3Fgj6QgaZnqNBng1XNdJjDJUQDfhrjJnO0TfP4IcKxm
ulH+ySiaXl7CyjAGBGN9tEoMsdJOywNIssfRHnaXGzs44gzCNU9ISgwr92kmvegt
WH4jZUYFfFRtBGFjqf4+EdafW5ot/fxixzWPFPeSmAXKTDsXwYGhQe3gYTCQbX1O
qvSbi9jpKQcR5OpOcWEXXd2jq+jhcURAIqogMX80MWaengfhm38DISddI3j2xJ3M
U/0qedyJwspdobXWxsIm9m9GVDAm1c/B35pIojBFgIN3wdM4Y85mBPvx8aqCuc/l
zgmdiM9av8TgTO2piY8ttVURFctyzclVfVfX3xdBehV0g1RaCU3SWwowRTdFerbA
iMRaQO+M1TjHX6xeL4ZmoHZtGKnSMkBMvQqM/QEUVIjy1KR2q/UYQAHDmPHblGtn
tkAFC7eOTo6J5UkTCgztGuc+cBkisKF8GumVwGP4SrtH6VNvJ7654r+Kh0s9uEGV
Au826Aabcc16+Ttzrncs1QAj2keU4lweIAs0n1ZBQV2F2ZDTng061OxoesBW3O3Z
AwaqwKe6dSZalsoIy3tq5JgDc/sD/DGyNCZZHg99QSka7kN6RAC8yrKJNhjHkQn2
pC/XYlNJu4cDb5CfVZtxxwzWuzWVYt9wgjziytOGV4ZJM2SRcRnPQEiJTr5ztVjG
8G0XPne3SwyCHFGY7JELCoXxV1Wp6s8rXSvgPtti1WqygYWzbcaGdRmxrcBpSM2w
mKcTTJDatEyWqxwWEs4HwJHhfeM9uY+SeuTVCba+PKpbf/xZbOSW80unpXE0SK9p
DwDtX1ftvUf7HtQhDDiZS22iaiTwUq65iBWguMgVktXOZu+cCIb3qDttAldv9RoU
49C1KQ3sacDzROJPGMoLkPTMPF6egSRvPSEP3utCui6N1J1iiHxk15QNkAq1o87Z
bYdedCv8B5tOxXPUvYEX++OIUpArZsExL0jZcRkMkLN0ENuD2L/2Oi4gSxT5y517
viSjXn5+XTjKYtQuPDUmMJw5XLP67Fv0a/tSA4too9+yuiZ50MxBmvfQam5M0eyW
IYfi0Rd0U5G6RCH+yu3EfJucpEqp+s0j+2yEaaj7UTTYTQrrk64qCFuG3alfsk2l
iw2oHXflSjqdM28jC1/XnmmpnzJ9Es+khPVe5tVphMcBWMHiXb9YYbuoqJlc5Env
MU+tRAoAQ4V0P/9X9UecpREZbpKZuAbnJwehmBSa1X6Km3zRyhMP7Q3OCq833s4Z
w5jWTvi7nspln0hC5YmyuCe3gPfNKcJ+bDZL3tVoZd8Xi1adG9AhVs0wVuE8VX3m
PPT3EoBSwAb/XsmxyYRLvciP5ZJppaOxe8jK7f05JJqezgOBNg12f8+TJhxBNgfy
f9ykXZZDNwcYawXsaWa9wYMGYj4XtjkMoJlsoEUjol/RRn+Xsg2zPwu3GZSUBNCH
L2SCTzXPpZ6kUlVa0vcBHvzYxNXFoKjizt/YSbQrvmjygYUkQBNgB1Fkuk0gjMSG
skP11eu1ZvNragvGX8tw91S3o8RZZtBxxlYRK2pST5ipmDj5sEc+yvzpR8S4N/P7
wNls0mI/oXWRwMxN6REKVjEVNhgnGRB0PTnWR/2VEI152gXYSaSczOTqURb7Yp3T
NzrJ343BXeK/UFIwxIsoFkTrn90v8rCtj7FzJcBVv9uYD2Ues+qxSWwSlCaMwkhZ
qp1/zxzWKcO7W4lbIcWhFjst3DVz015B/SNM9IPS1MEKetqdejmm37kjI7bYMMFf
rhfceh+k/u2Ag7m2jgbbbj5gMPfJ+ZpqW/QUVwtgowNNQlF3UmlIGs3IY7b2ZR3d
P7/OssdUV04KPg80SpBNlAEpuxpHByVmu9z46cunmzKr7ECXGPAhXRqYWE9J2uow
dBIwue7BZ+E/bEzsJIHrvNX0Ip6B4+Q442mIkNO4nS3vFP8uPe/xI8yUMI8geHeU
t7cNASX34A+fTuVBQjgd+aS2VI1xRWGuifCr6GkzQ3bd8n7hOajQuHdcDjjm5CC9
vICuQP6i/yeSmNIMkOJg3h+pqn0m35XM/tS/LUh+M6XFBDF/hihg3i2o9isF5fLw
U3HN6ArOV8QTNfYAx2PlwKYff4D04gZuqjVRVFzsA/DcABkhEOJh7kw/PA7pkMFa
A0v8dQiy7nGsS4Dj6yQYGZt8G521cA22xy9ZdHS0kOLz3H2cL4/hPXFbEOatiIId
DVMVXviNWUT8MdSgVSMN5ynXgkIOK+3K/gb/3yR+w0Pz9f1g+29OUOecDADPUHlw
RlfSSdHiamSlgxzlKm6REmdqAhzpUi5bnRto9PDOStSB0E1Z3CQmkHZlXPQrXoty
ClLdsmdkTN7TSt7pRnpmsT9Raoua0NpMeA/my18ZEe0XJELYtaLlsFTMxsyxWG/x
UOYjXz7O1QZtkmKd4WWxq2dzThsaLUwwAAmzEM5mQ99aYWL5zxKENwHdHeIb76yG
wAT3//kaujV/kJvWgYiHBwdChNOwB2UpNKt4acoSoFdddT+xsCaxys5xjx+z0ZqD
I/dBcYevA3/5+4N61i1oJtFFblrmhB5BDqq5jEIF/6GhGLjcyl9MmDlg8ktrgvEd
COJrYb5SkYGycZWqmqx3A0VU3WsCBZoTHvhSn2tJNFPuvSVY0DBLwzirN8NZiXca
CjZ+1kk2lGr5cSVGeMJvXYxVXeDf7yrMHgPO26ymmLPwgDfKbT0ftVUEX56OYMa6
17f4QALdOp1jA8LGqjATxUWMrEJdaM5uT8gowoIxMrKVC/WAU4f1pcf9fPIVYvlT
u/lGbIunywbh0vCuuFa4zbXuCP4onoRcy1FS/Kvy3PMAuhZbXwbQwXc/Mf3RdARv
99T9ZR95RfqmoBoNGrXtx6TGNp8NAWwfW1E9EqZNE3rGj+qcNelgumw2rkSzH8jG
fOWDtduZqGotVLTU1pxEd6k0kEkWnaXMwRzCZppj+lEwkEPXaEq10ejwSTDoLSTN
uwd6SR0Q2MCOdnVadtE22+u83QyVIbLuq1BI0era6Tqosv4sp4Fj96t+dtilsfT7
0XsLtKt6+lbEmUqKRIV8EjYKmnRMskXO3LAuPf/2207QTtOhvSq4LeojsN09OYLo
d02FcrHfSaXaitXOCo+FlOtc3Z3WDggsWOvd0PsE2zGXaNF+BS3DrqBUoVUIqUjW
Zbiw+CEKAC1uWL/yS0CFKEwVSs3F5aeC43/5tgOxOfnRDOxf54opt35yA6ibl/oX
wlL48nyxV3XOO3NNazXpX2Z7Ab8HvqiXNx5wgkKDoF3klMJdXtWs48AXkVwp/YJI
50Eijtgm8Asot2AuUiFUHc82OZCfn7NKDN0eXGPsn/YVPlftd61jpXDQ9hU2U41B
p4Ko3PYbcyNbwmqCHWgBIQrkyvQdDSar7cmdPSYmh8JZjvofKgbbuaQD8U5LR6Bu
0eOCPa88U+muBNMJMyRRTJTaF0IjYwAeQFXd0QQ1WC9jbpeFpFz67nEiJSDwSUBg
tGwZzlGf0nBK8J431sK3Refjp2LV8bnQcXJ8Ka23xfrG7Th2HU4cK2RF1a9Ez++O
0eXC/cH45Sduy0sXWmRbS43IG4wIkrgVOm8EllSsDOnXLl+gUKYPkMiQYcLOs2j8
W58o9Oqf1pNCpJ/5P1Yhs4ttRorkiS7zcaWz/3Aje/BAE1W2959QQRkiuBipSItU
YqpuvkhM20NAw3hy4kBdl5dUqGBBM6Sk9YtxwFCgVKfChXBI/805aBcHA5iP3UVr
cFFkpE4sGpvzk++8/eKbPFmKPLXZL8rTlw4YxZLuNa29Ku9mEE0moDNXjvQwJuiL
3uH/wUC0bxGFL6vQKQ5LxIltXuTDdnE8mYKGxdU8dCBLVxEkwU9dKR9n9MjDaeLn
NqlYqeCO9FlOpOucp0sRLSfZTBu1i73wp+4sAoTjWo+FFrjH7EgO35cv/FYt138Q
f5l9QiH349H8FfNN5+3J3YYMkSd0HY6Oknoi9BRAPhAKiHjTBl0KQz6h2lWXJTsl
Z6SrjaG7gF9ClyTQHhHYv3413IljeIjCFetel3FAwdIJC1eFJJrGrYAgFgIArxq1
/OsrrYvUWCkR8z83phpxRZ+sJ7kw+FZ7w2zjWi+1QhXMPjwEKcLKxn3AX7ZdQHMo
UssSZ+f4CqTa9D/WuaI+QlN8xuVIYaHoMuSVEoKw+2/YqY4BTlfaFEP6KINLVeUJ
BRn137zga5lIFDbHzhnz/D51HQIE8i/9xpT9HBAm3ufEhWMNqITC2HxsJ5K5xZ7R
/4PTmpgAZuDBOGPax4CY970Ibw5TsOhzVIpg2aI0WmtNFbXz3ZxqzaquGlsP5n+C
d0fwKIliInRsuQ/5lyler8wdFIK2bBs398//LH/Nlc6y7I+hKHqaKkQ+2bLWDRDy
gEkVY3jjnjB1se0a+d12LMjVx0o9BKYhavh/NmTuZy/MrPlR90QMREIlyG7nSghw
h7vBk2QK0fQL/+PRAxKE5Yh3V6a9Ob7TbjnnL+AXaVUJke5o0pdt7XduBiNT1Cqw
tmwlIvux8VdilVI67X763ZpfGHWH5hd1H5Yypx0M1gtTnLwERKim3OipbGxJ4IPQ
FGazHSFsMVHUj5Azy02IHip9xIl7O8wlyNbDm7SWyBw47j7wkAd3ORl+QKIfMt6B
jx0AFmqBlwvKzRRD6FkiSy8RMvhMPtWk2vb9702L45H7Hovac2Axn1bOq3QYenQh
PjSutHctLvywko36Qwcocl7z/m1K74tg/XJwDuuoTF0IaQ9jVqR0OvrBd8AUJozH
0mh6ULnmZx32wxVGQmMCvyNif8DJsiHZOLIJi7B54q4j0hd7M+qExbeeSN+0oT2s
x+k95R8H4Fi7kJ8Qxkt9C5p6GMeaBAE/vMs9LOwozPqaqzc1/yTDRwXO90dDDeWL
5U68WWQfDdpmdS8MtjMCrtYuHdO+B8ED8eGQd1CG36AUe2ZI8fiP2a9hyhhXKH5W
/pa+qLbkAgpRSmYzwWiIl+CIeDQV8Myo4Cfimv4kRibVBKne39clXU76IMqAn8fV
0kdymM+GikkrW/QeMQ5WvzsruWMeBj1fLhKkew6u4au2OfmDtCDgJH9Qyb1zDkMo
ZnNyZ4SOCUxXL94UQju84owsUCknwI4fEKGVVHkOE4dB5Le/TZmOX6uwf2cfbJib
a22rlmnkoFeY6Yr9yM1fnGpgoykfsNUOV6fsRJBqidIEvan+Rkuyt7rRJ6NX2w8f
eRspv8yLHFq5URJ9I5Gl+CWHNdOkA2exdF5Ww8ZNR/jxVziR9MiLUA77Hg99HLRb
m1n5n9ubfBj7X8t+VUFTgEtXzAvt4DlDpqPc1kMEUQO31cWcrhStYq4Xy6mqACtC
JJ4+v4AVtKyq/HO6HtkRcbfLSTi6TDdRgWAoYBZyKsfuxlNwlUDGjHV3wQdv9gXB
CfQ1ippz6if+CvmTNVRHlq9zjhL95gZU2BQiPucCoz/LBAF/PvSlZ4E1kO9412pV
wB3gYmY6iZyC1zF07uF07Yp6QljwFDtG6baVDOBsAyjLEKje2L+2v9aMiKMpIkFL
fw/nwj3Raof9/Ut1rJS5GVeSc/avbnIwGDawsKGTIOmmazkBbn+184idGOjsN7op
uy5HrU0tZFsMXWb4nSQRbuadMmEMsqxrRNJizAPszn3u23Ex8BNyb8Vi54HAvi1f
FQFxzrb+6JJsfyhgHafuJQbVL4aHOP1haFnnVuVTMGNz2+0wOFXDRmaIncSGC9rN
pj7cnttfieeAP4R018pTjByxRfVjT7Khjg13f9AcJc4Rm7jjd9SeGUCLzaf5bWqa
Nz6SI9SqX4NTS6DU21EM6cLLamTbYRoTgyKHNTzhgB42m02B15Chcec+3787QPki
XmB91MV6MhzjTglviOBIVy5DnP44mRABYGKW5MG3hOa6u51P+w3BiKx3oz5USDdp
pvCp+u/Opu/nbvV2CC1Hj7lwF8YnHF7qUY33DU7Xxikdqt4kukpg2IrSyK6nbAnD
UEfJuHn2jRFGn+r3IK3Z9eqKyu4RSY2a2NfrBkjHh4dX7ctdrlMIdlMIS+uWZw60
JvhZPHT5Qu8tnpn+oNIDH1DjAHSlpPVTp/7vi2j+lYK97VZ/ZwBWx9ziOsjUL6V/
UHDWSMs4Rn1vib6k3bznamd/dsYTDH24s8/ySRLD3LyoE7cETHJBc7cn1paDzYJ2
a3DQWJ7su02o0Kzc0EUYO8ZvZ9JRcm/l6NU8ZBP7d5er1V+BCg3mzoOX+JOlP27S
jPeuVuWglU9o4qBPMkqsxrs8vh9YT1W6oDLmw+gOwvqudj5unEMkO1Tbt56dVmB0
kyaTRXTER1Ul82ZDvyunigSQjG54wtRV7jg2fviiczeJYM64y1CCKtVRdwPq+yiU
kfHt7U2b2fm/TSETuL3+NQ8qrrIaCxN86dKnGvuUPJmIjhXYMKG/sVcMO1eFKkQ0
6HqgQ0WxH+Q7qwyB8MExTp94isd7DM43sKXnHvGLPoj+I/O+Owlz9P4i5Ui9Vd5b
BipZ3IJ84jSyQNEaAI3ORJCXXh/o04dSbe2s+vEneCq3zZMQWvoYQ6xeM+qrF62V
2TJNdjtUN260axnMaCqdAbFw3wt9oLpMea3z1W1sLsydF1c4r1eZ8hX4WpVdytul
bvUvuCNK14F9x1YE/LhFC5DgnPZrhvU2mCCI/Ht/HZenCfvKfdHyz4byDVd5wz2K
lssuz4uuTZ3+Iw8Mwrrq/HZ5FhLQO6q/oY5AttOQGMK17P+GeMIQh4GV7c2ZVCgX
oZSIT/fj8L0KMQjgqVGaFCMN6cTJYfiPyCfODJRN+rVxiO0ZfaK0xRQwQrQgdf6H
SuCOZhupT91OMolkaz/yYCBYZXKoFJA9voS7oDpn0/wSCWtb6Xt/Ne+1quJXPPrh
01o+g6WLF8evHWiN4y7Fon7AuJwc+V52M6D9xa5EXyVEQ3x3jLL2QPKeTCgZ1rHt
2kfIvAq80bbOrDqXV4XaSagDbNM9QPPwOkPoW1wjO/z2KZHpYzx3HVxULysX1064
TMoUh0pjkPryf3oGqXOgVyWg1FI6VIdMa3LzAJouIj29EgohmrU7yrI9wlloYr8Y
kWZZQyC6+Kc9E6reVsL6YtUdFLenrWGS12vCtj7fagomnR4fDr0rnusymggQjmRH
yMV33pGnJpRDQTo25I1y5V5DU4ZExjoY3jBcz6aEdJHx3RyjpVyZC+PGqzgpW4a/
UMBYdsbukbskF+JEdBth3MaAV/QwffiEuLFREBi9R5Yj2+5JirS3oMTuddqSV5Zs
WNHc95En7Wr1IHc6kCs641oSODzGo9mLF7msARH/0NGSucXipba4B1UcKmFG8u47
gsGDU6/77BEjuY/2VRunYI3Dgux+UT+BsiZYn7ekPK6GFezXnoBQ9cVBYE0HEiIr
XLJhFaPPzbx8ml7BgLja8gYkH3/rxlkIXaHSWJ0K/JH3FdLrss1AEgPRYPT/y5Me
Ds/0hBwYFGGcjXRbyhLy6Dl+Qq5RbRMyhF0/glX23t7q3/o4L/dGlVeGUCHGUIzR
Otd5BRt72fcX+OMLrxOdSCB83F/nd8GjQmTAF4Ct9P6KQ18Lc8przUxwaO3ou38P
v7ln1k5tj1MPY4Iz1ypsWoFyzk3CKDWug5fZo8osoAHMiwfvx8c38PhWGvfhaXAH
gI/m98/Hru8c2kpOCE1+ro9C4FDgZf1jMOOUJrW89xXjdraQiDpAKM3OaMaxEUBi
YtDpQZWDNnaXgAgddKEfXN1cDbM5wvwNmq52mX+6beHuOrvOOKaPl/yxU4zprOXk
/6Nc6GWkXzpVTCBELAr3EPZIRQVcqcKoTXWUT5NvoFpposupAZtB3Y6xuZJ0B2EK
TorMocXfQSsrvTsksiAf8goGx45GLc/Ft74xO6hr8A/SC+QZo9z3BKtmSDL0/Wk4
4UmQ74mmxb8YvSnAT8LrrUIyA2BoANaqWl/Otu1C5dMa3N+SK3tqjPfWLDSH6r5U
93N03NiY+UIDkWJOBbEHH0q8CiGc4KufzoDue/TDNaDGHmkznVRseS66u+fS5KB8
YuN6BUAwgdfWHv7w2JoaNwypLsKkIt3t53ftKzrOTIRgdBYt9kF9sGpGZ2C4X3o3
+Jxc0O9tTEbmtIIwQj/MxLTtxCqZ/bFNN4OSW6qyvobKIIVVp/NlCqynTe5Bveq7
WbeOGP2yTydRmqMJHc98AHr9ZLOgshDNRxOU2UOCipbKrciMQzfhqmxsxyyy7IvS
uUTpEPKp3JCeAtEH/PxAZrY0IxYiI+biYroyxYek6upnajPo9T/fL0Eb67/a/kfB
7PoG8crwBo7SdVVeVNFiphmwah34D1n5wO2Rh1ZN2EZiIw0LIStG5ZMfHj/EKyI+
fa9BdjMHH0f7Tk7kKHBcNRR6j9JvhBwZv5hWl2+pybDl1xckQNCrylFgrcGEFvAL
rp0kog+pxGYyvQ80Kg0hV70xIyDFeroeui9/8+mmsHbINIvP7o4Gm2qkGGJWfGf2
`protect END_PROTECTED
