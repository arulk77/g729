`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
PzH01JG7X0gwDIdYA9hjmYzCo8tJpAxgUv7CQNEAXdq/UFHVB1sJ0MR+tuYYa9xM
glVwWknsu5zl51/wCeT4/QcJvVeL7RVBA9B9jOSFV5k4kb12jjicFmRaYra90USp
8LHG6pxEeHyvvLgzrUQ5KILsjyrlqqJCusrxik1y/mZG8p+pOQO5JOqElXW/LY0e
lNhkieHf6TcZJUqi3UON4muwxJ41rjXRwr444ueMnL/eiIrjCza5y2Fh/lP91N/T
u+zLZR/NqTepNBvsWhKk5shXUs06WJcDKZ6aqzkRsxPfLmE+iUbwG/pghOOOrtQN
yu3E2apgDeHC91ZOMA2V2JIu1z9oGjVWMy6FNY2JLiI=
`protect END_PROTECTED
