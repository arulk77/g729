`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45PK7MUJYPfxOhwJ5LyUsJuO5GGDBYo7IxfwIBgazZW2
4BkUdDAoDllzIJ7HVb8L4MQzhNCb4LfJ8WSAc3Lc/o9P4BFsRtAGX0dBjl0mwm0i
4GIvGBQXm85jtWz2YM5C51CZk1sPEc9B7U4Z484gNkAOrmyaj3EDlAthlyk6kjW3
LbwMdMuOVYNCdQLqnbujcRaGpIDwAsnMfUzkHpOFKUPll5gLfkqsynmZbX6awj1i
SY8kwdnqV+JA+6piEOIUCg5EctfCrKtCAtjcpvyuRI8=
`protect END_PROTECTED
