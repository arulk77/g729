`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
dzkbPpKoSD1jfb8vG4yMRsKXWrxvJBDzB0/PX9QWZ0opSdP/05egqCiMESzwNplD
8YYk5xgh26W1tXUzdqoTcyfic6dLQ/ezKr6ujcZLVkHzYkhxdAQ8zeFChQVUXLl2
7GA4CN0hsnrxdavppLjQqEsaZO19u2m9HH3qktaTW/YHlt2E2LKlGrYSFaDPn4bb
25Y3PqlWAVxNJcLgkoGR3BPECJfjcSLzBbgB9y9L76rbmD22HSjx/ReW6MNPy/EQ
hrED2id/jymd2Ac0rDwnj6orQyuo2PNFbH6JRNh2/PU=
`protect END_PROTECTED
