`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
1GruGSu9PglXC1oa+d2P6KMpoj2iewbPDQoTJc9cvjC9vj26DyhVWAb68cD1sHDn
tBVrYwVuzMjFfQR7jiih72mqrlEpRhlOkEiihpHveznSl213Sxuj8sOU5+HiqGZN
7+8Sq10EtVUZ9U4GrTc46crO6C8a3ASCKCkXKYWRJhx6ZV5VXNZzXWZTIflptF50
Z2eTI2dZ3cqa6W4WvhlEl4OyQX95K9WCPSKPi/862fVuyPNoQHHUjAVMGnFOfGk5
cc03gDIAJdJiVL6qNiSkh2G95waGOVsRHyZLHWY22aN1LhHDNDf7zcdfrBKWBgdA
eklQiM7rKwjl8A0x39XQb0PNNIpyihayc5yFFeHY1BdyCsWmEQEhIIu8Y6INRwwo
Vju/Ygy43R2iSEPove+Ays8kZD6Emw4sP17UXfqpCV9phfGQK2sSlUZxiCS8LwqD
WMU84wH4I8VHm3JNZBj7hcrfolhyf6L0LLT73YtEFt6uzdnzU7zIjEkkLr09aZIt
n8gyoVxwtm4MWzUpmAklgEhy+KdrsS+WCX7tlxIquA6SQX1UzFWRRTpxyQzK2rLl
ZAV8bI2LXKUvxYz7ZC0H7d3zAcAbsFknc8UVz41jG6tXffHaJdYrYo6ALAStcLEn
rtiznG6yNF1lX0oc/URX+m9UQ2r9Yig0jyg67aKTnt/hNffitytWdgjYZsodfokv
94lQlT0ANlq0EzO2mzbSTTrWw4iAh8anZeR10bB7ld1dZ7nO73rDBJz35/BNt9BL
Bl2SETzmp3KT4l9btRtYUccs0TmMXHGx8pPvRk5VdEk/O5xZd7z12ccXMHgHkc53
MDCkzZJo6RyK+b43cFGy4IPdPxCayn22YzGQOUrI+Wx8O3kIYGNKJ9vOmqmPJ9RX
lv63k97IS1Nza9LH5mQCJdYeChpEbE+oJMIXt1DiB4ydUcnmsCu/YlOHn3aV7ntM
Uj7jCz43C8IZk6Y9Gu8Y2kAgPBW3raZAADl/6Vdh2BFtZt4CzUDiTUPHrUIs/0oD
/ndDN2q9BGvDrZ0kgcdVFYWqE0wUjwg4mIzdqKtnJVzM5mUP5Nl9lMqCRbzDn6mi
ki0RLi9TYG6PWd88UMAnR218dQogD0uTtG4Xuz3ME3Wbtdh52PkU28jhrdRbMy3K
UVdoixvShIRJCNeHyFzGgyXV5KpSNoCiHeOaL0tqduTQQaf3RZlDdc6jhguTLu8X
0Jgf6BX2zxqVXkdcSTQ1uDGUc1Ko9/+a9LPlcegzrSkT2geykrzOYpYAWMrtskDY
7apkMM3DpW/ZL9tviA5mgDmeW40ovKk6IROzN/bSwiphBTBBuhIB4MmzeKCxZvOs
rCTTxTOrXxRwJUhBiRLlPxVh4tCTAK4nGC2kRXbAaJfnIiTbB8yIcXBkoyB1Uix0
zRxf47wQnDQIQaqpbzB/+ksF8h7o3tvJiYarxThlHmVqyAod7+vTgXWTfsAbbdBv
0y0YKVWrzQ8u7ij0DovVu3dG4fVKVBcxbg5jsuJai64pce6UirWCThUKSEOajOev
OIQPd7iJHxSzKTzcfKb+KY4J+QTLLoAKJcXawQGeuBIp0O52YiLuDpNiLkc/EjRg
iwJYsdisOGl1ceO9sgVgeuSa0+1Ef0+Ob0Vk1NN/6Xel83H1QRw+q2p6VVjvFAZF
xhUxgavNDwU7Xng6qI+iF7VJ00MzmRiVQh0IauzWubqP3qr4zSViFbKFgULZNSli
nyumioLlPtB8eSCx64Q7u70xWFYwdeh6YDHiL7koDG8=
`protect END_PROTECTED
