`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43MpyMQfeUDPxDQuBiqP3hQdvGv1ZV7jNWXvvPV/v7wh
1es7jum/fili0FmjDaQ6AuexGf0+U6sVjUoTtFdC3fm0HscPjBbP/VM9tMzFW4/f
CSDin57UQWE73y3uOYkfcR/SVLC9X7m4JUGEiPpEQh8o4CIeENeMuQURs1ElSlpw
f0DdnH14kRL+/cgD0CFyN8K0L1hVmDGR5J83EqUhjSfIC9R+Pp5H6Gf7CSKlU9/9
OgZQzdVWDaKAUpOA0tMjgEBuMOV0AQT37M4l8tAO8l0=
`protect END_PROTECTED
