`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBjjP7r4jU6REdIpIOzHDbCGkkQqiGqAo/LcfAL+Zrar
jNE3j28cgRjamXmWS8RI8EuekyVYc0CDzpH+aargBqwUmXBYDtEgCe1fBEut0GwC
9KRahInVn4NhFpn8gF6TP11W47bGpSdVwH5Jt/L9KW1TCjO0pw+lOWqs+p+UwjwO
l6V7XXfRYEDNsEFAHRwl5wKUojkckcKA/deGtv+KY6wvnpFHEbDv45/ODB3dn1wz
Rt9EszaYocbo28WxphjED8Pmlq8bGxSz2KIHHhAo6zBpAx5EepYiwkY0P91v4u7p
/j3B38FRuRnCLOLk49EjU/AcxYIOj4SVhi9U/CwNNFoYyTral7WBqD4V2fV5rk6I
7qJoYUJp1luj70/CtnAWcwwyrLHEUltmNMQll7dyqEEaTNeSeRCLFqq9XvuZIau3
kUEiGouvE5AuQiCWUt6CQRws+B0Y7vWM00VfNvFVSBEKLVPKAezgxQoZw1b7WiNZ
k7eu4KgqBlsoG/xZu6rw0e0REDOnagaZPpiEdx5akAn0LAlQrsuAaga54T0yhc8G
iOTRmjAxhg6UcfAdSFl0k3ukbzXcvrbL1xfyh9Y3eOw9O83Miochm5yCTqgMpnGI
KjwiegHtrCpsJKcxgU/4f0vLA1U/EQHU4SGRGAP5k6W8/5zTiW8MYLwRSrfm4ByV
gYp0fpDm8OZTQkWcLeB2tb8ASjZR/IlUAoqhfjj5Y6LlxQ+bTXHDPA6wKxY0fGoX
KU7Qb35efM0gE3g0ECvfLPOFBJIB9KLt3PpotrANvrvaqhD49q4aCD7xzBvbx0Py
vUnvSXQCsh04rSJvyF5G4HXVBmP9/xoyob+Nn3OzsIFG47FIu8fz0B5LvowgE03G
4RDoxPA9Ge3heDsdEKD7hUggsBX/NRTrNVOL/nzNFkRgTj3jHLyGBGExmDXaEGoZ
mFC9G4q1XheZdZqD59X/Gmv37BIgrCyei+vKdITu+d8KEddYFMFhguchZA3QhrWk
A8h3lMcL8CGjznD0lCHEMX2oN05Cw4eNF5x7HPdQGJu+Q4wKfYZ0SBVYFlVT5XEm
SrrgnlNh56kJZXjfhdmWuxm2nlQOpWzCgfOWZjshUcNr7MQNRq9yDJaDyLWMVtOm
KIT8QDi0BFpvWj6qDAZhMRSgXGfdyO0srIHBqswVk4gjfUoSn++vV7SnZ+ykbGsI
Cop0BO3sACdqlpXWvRDlyXh1UYllY8VIeP0Tq3SuF6Q9WPfIZYovMl+SOIgzrChQ
8Q3PHHtdPPevq8ZBJBzz1O6oKbc9fsWKtmEvvIGkTZ/dqI1rtvRGmHMI79DfEP1c
l1eBMklQBi1DDBtS86pzFjZ2tVTGDWo8gw0DSMkNysh7JMq9xfJGOTg+xsImiRwI
ubNPSQZ7nyQdLAlC9s9m/S9XdcTnjFbpTOEYy5eY8jWsgRw4p08G56D8lkVSjuCy
qP+yfwsEZKbv5S+C+PtBAxQWTl9ANgHbgrESeDV0VJn+lG06Ckd0YB2IJB3IYrW7
eKyHRbbBkqa/n6mvAq00USasrFJPNTgX4BhNrQ3+VrlXwQRiVT3XASedkTc8G4y4
NnU6P0rOoxv56dX/HIxZPJBrMQVeNDwqVQ1ZX00IGykrzPdUQnfjLOsnGAnnsQP1
MwdZVmyUsnmcipHNGySXlxchgkivv0OmqJ+DzPdNnXkiW650TLhZcddu5h0g6J+g
vZXVQruBFmApxowuD5jV8HIO7iFXni4vYqvd5H3GEmKugtLcoaS61S8ZAiyFRQek
8to48k3MjrfTm2huE/B0wjcYcRDRqQYbVhMwEuU+4+ntI074w1+D4Qnxvm/3l0On
`protect END_PROTECTED
