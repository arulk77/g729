`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAp28LORrBJ5ylRLvrsLAUD7LnwAEFDVRS/oLM3mK8Q5
zSCymndYV32QpyDKIFy/3fvaMvOGuUBZACapKB1YqxrQf3DZ+N1K14ot2dOpUb5Q
y35mHyiYuC6hOlAxH8083c7h4vGlbBwdloWAw+eIlzj9glccCe9x0ApWuXM0KQmz
jI3jBz4DBjvbcdl6suIgcMc9HpjCM9476x4XUsxyAoGBFtgZ+04FPpnJjSEcBluu
bo0hAypWp15pzCfF/iHp994O2cyG/wEPXl/K/oFQeEd3ohHkb8VUwM2kVMo731Rz
s23S/YJZdfOeet8Ej7FYN1NEd7LJdNQw9934hk8sWJp+Lcj+iugv4ywR75MgVoQ4
ZdktbgJfAO6W/1mJhdV1YOIpaySFX2e0sQEMIoiCQM6AfoUfnE/g/SVGd6SL0tJm
Zzxr4uue5iiISrxnLcU5eMi6Q+/3GFvH8z1r5DIYmYV9PI0haFw0s6ZlV/GZbBnS
`protect END_PROTECTED
