`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Zi4MJInhKvZrflDDs5uBU53eCkZCK/Z6FTvh9tSnqAVuKptKC/hb5WH15IyEKpsC
cbYZrm0mktjqtzwv9ZoqD2VM4/kB3BIgHnCKFkSUiY3r5AhOkPTwIAQFOK7SJGiA
7kbZqOpAjtmvL+DIk5WrBDgYmTtpBaf1FxiNjSRIgS0=
`protect END_PROTECTED
