`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
rLIi9h6UQw8JnHeay55uKDoz8TjO6yohTRWgK/QZ+8AdXvwk1y7KB5Qj8S3oFPaJ
iMA0qrevlX1bZOZmuX6HngPmnPvW6sIng0zc8aQu8WilPMf4UNjSzg25YI+eubqa
zhENsNFdnZWAOE/tDU4Gbf5gV3HprVGwSTDgJ5NO0lA8q2kW/osG+tdvwJBRQRj0
2iehZbZ98H4akfPHy8yrUR8ltHpwhVwx0BNPb2kd9X+tyDNGWpd2sMlpOd+Ft2cH
CZfoXl2NZbMdkCFxIkY1HdB91lIP9tBLBSYq2+1sLY1xUmTON3kjBx+gqL72xXTy
FmlzUVqKeUxznPJYuUBWOn+QSiZk765iitBgTTU3/EGbTo9OmDjIBhpcPKy1InL6
Z+y2kFFplQKKVVDcX/eV8nven62Q67iY/LaiKIznhY92U/uehuCi3N6tGBxORTv2
M3kJdYGt1zObBzfkassqZQ==
`protect END_PROTECTED
