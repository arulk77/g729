`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47PSM/gs7ZrKPOCw6VJc+zA6QUM3f6okVT7l50WaopWF
qGvnY+Ux9NP98fC06axi7aDtdBkx6HWHmNIcMXTAK7C+tGYBFBNNa7CYLIGgfyE+
aTSvr4xvm5vHyDUgpDZMXt+Ojm1GRaEeRWS5EQKpDZ+SX8G1jJRCb9WpdbdLKTxW
cbiANKV/a3W9llWU2CGtm8ntzTMEcjznlJHtgJdXutM+WxrzWgewfVnBfDK182zg
LECAsMayoxHep/Dgrwmw66DrQvvr+7DsfgDa6g7Ox1uB4OjNP+YntSMZS5wPvZcF
awZU5q9mpUY6TKJzh0oiUg==
`protect END_PROTECTED
