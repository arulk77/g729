`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePxRjlgTev6CeZ1bRrxtw3dFcVCTrMpcRkHHbs3scftt
yX3ejnIJstr/EwFxpp7f0eFsypdAdDQi1XXzlFNReYsN/KjUI46M/O4nmmFOc+0F
FLK9IktbKA1Pk2yqAwD5tO4Ym0j+K0PdFtvkYYu0rb1ixISFpFgP5pCYkzfmRUO0
codIQ1XzFzoL0Zfi94ARI7d8yJj6j+5yIsgeV3c+GcEn+TAegmObGEyMJHfh+1bL
RGlc06dEUqwMUweI9vVRYHFDNZT1Ad9UGoYTDJBbOnn/3bLSrw6+EVsT5/rFk5Ga
H04eCMLDb0NWBAlmDvrdR3Ubd4zRcgBFOY/7SZcRPN8KG06ndRGhVEdRRk6OHwFD
aalEJTcLZEhm31aXDkkqSw==
`protect END_PROTECTED
