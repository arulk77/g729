`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB4EeKvnwTl80f3aanwyjmFR5v6fVbFuRshckXUKfm1B
huAwBG9Uuee462IM+Co41TImJ+/ZrrHjM2gAcX5a6ZFbvjSg5pSZ3kep/lAqk6Ac
L3WBEDSIF53h97PETNrB7cM67ScCDibDIqpn3/qWDdpTxVfQF0gWCHwWwxa3BuEp
RHulOZ42omqWudPqz9UQqT1DseeQhJTAoeSSV2Bxfo7M2beDHiQ1THiHAkxd1oww
WxSmD0bqeSwUQS1nUhXSSg==
`protect END_PROTECTED
