`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJioGSlNuyse20VDOQFBPJKlaHhb1Fu274lEROY7ksU8
Lfofh6MS/Cq3bLIEkcVeK/Ce4VHyR46fN7LhKfngT7JFs+LgyzT53Y3/2JVojDAD
vW3Ljh4T3/Ti1SWT+nfaY+NaYJ6OIJwwhuvtdSxI9XJBzWA1cNUjRWObJjfNB4OE
IQKSEvQpRKn8i3q8PlEnOd+8eWrR1XAeyVBu4Cx4V4cKQ6xIoEw+L0faMGxQDYVW
`protect END_PROTECTED
