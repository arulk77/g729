`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
nl8wPDViuYhFIDHPy+fhxtSfHB1tO4HIL/zYdPVMIMoA0MD4swIax49uYP5rG9Kf
75bm0hRfSQXb45vPBps2Cg7iXIwevv04XGENyOGFiLeoWBa7kY4d64Y7CmAIZHnF
/FKSVRZYSBtAS+gekhWPm/EOubAtZRLXOn3s6LXOIpfE03B58IsQ+fYj3Nw9fy1/
ZDcXOPDkZyV+TnbkR+SHU0ywyIIzBBJ7x0spWrToMFy2/7VaFWlUNZN2ssx+/C6V
xEnl86nei/GXd6DyWch3KPdnUB9Hf8bYGpXdwSWnNts=
`protect END_PROTECTED
