`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
cJLJDlxDbjbGXTCmkf/yr8sBGkUCIsUyx1pVhaeltA0VlkLZav2609JqNHWUV/OX
paaAG0vbZTYktU2XRvqDWRCCHTm3RgFjKaEMbAw6LbskArbPZRwNEka5nOOxnOe0
a6ghDtakEr7F2zrl1LC/g2/cMSsfZ5Cb28p/2wh4c8L+a59zNQxAZ47xvh2geva1
kqBCP3LaxqCfVqdharf/CbA4O1tav9RbX7jCSHPTtyH+r5cwLdk0weayYUHWedFb
UgwIzcVVrFpAwrt8vgTnkhAc1b9iD7y39kvGeejDkxwKxXikgqKjjYVTXwge+ABM
AlyOD0zEtQqSInWkgBk1Lv/ZWq16XI0gChdgKJDJSc94xv9McO8gBZ4F2aS71PpP
Thmr9Nnp/Y3qimBIc1F1/n8CfE2UqhCCvbZlFztkCP0FwQvsGE0LKIhX5MMCdmwp
Vf964UHBCNCcFo4lih0d99ZGmjQgfutW42IlrKeL3qe5IiKJAI51VVIgyvVeJdxg
vQYP4ZHZtUQXyg0VwkUu4vmfVc1o/+gybgBhztd2UgdPixTZ0ytSYAqgZHICoS2K
rtJW4LSkID579r2RWPu238VRsnbZJ3kuB7OfTr5bYZDHCZj/L/dlgOOWwT5+JGuY
dCVAoZOo020NTZJOBCnqR1oIDgycBK3OAKrl73hr+bsmbFgABuZ6NM7gkhz0OEGh
yJWbvlOWDUMvTz3EQq7jywnPdh+b7fOb7uj7ARWf3smV5SlmXDlZcL/fj8KoZqDS
eJhvKsOCGEDVAXV3jTuiVELiLuPW4IArJ2VZBiW55x+uqTyZfEdwqQNvatjF3NnU
nFPuZllD4j4nOi4PSSZQR9UmTDHebdUqInxWT1AR4Q4=
`protect END_PROTECTED
