`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNG7Al7dqDSvy57tprc8jJ7LbVBLO4K9syqtROiCc+ok
Ap1Tf1zg6sTLgxXrOpwOK/35c3N+wyj93MHIu9yRCtXLmD9zubEyN5FtyOIJdrzj
RLPcoPN9XCeO1QuwI0vAtPfTXjE60vkznp/5sOSMUSjUPMVLLgJl6pRoVkQVtTpR
ZpZajS9a+nWqPt3U/DPu9VV/Eu+nLP4ECncgLtmXPx/qfXF/7HTX5lxRwYQQpD5z
`protect END_PROTECTED
