`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOOHrb+0TuG86Np9/Wr9VKtNdCvjBiE3F6/RBHngSOm9
CkiP1+hIGgMZz0jdnYBGny7+l74JkWdsKMGD+LSxU10FX+hNS17h1JrHiUpH8S8c
7P1VhKExaNOIy+lSjzB9exmULL0NsfHfULACRZXzV57EOowmbX9wjb0dd3m/kLEM
uqxi29JfA7Rxbmus1Yvx0UrVojz9msCuXoJy48LrHpLXcCqKzJ4KeZGeg9n+qW/C
7mhsotgSambct0KfEyHqCbRZNCooqr5ov/2eVlz9htMuPE5Vh/qjOrr2snSKUzDJ
Zegx+zNbIi73fM8fePpYSRxSbnBEPOSvNi+bpslGuLd6GVkLeHjndiAQHNby6x4w
yebi2LQzADt07KTlkfCRri7sSodqS9XSdYj2HHFb1nvsmzKQpgrqvaZd2vQ03TTY
yCrhk6PZSoy/IbQNW6OUDZDTT9p30G2fx8sB42S3DD61qq3pwL4cu02OqYbUeVRu
2RTujxj4ENl+wrx0pgb1ZWPpuYHjXYkbPpxbkYgsruWcsOGPI1VAJsk2Nw4Sy7uV
jYO3eSWv4grJl+bo16x1GVJwp0/yKIT+sds5CBHjT/M=
`protect END_PROTECTED
