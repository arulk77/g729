`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
LYriZfFBBcfird61amq6g59fFA8kuEXUAsgM3dl3Y1OxE2RxzXlbf3hbPHWRuSCh
Cyafa/4HnL0oSSNUsFj1g2SdwZtFgI8YWEfzHP++5AU3c9NGkmBCI9Xtt84QCyZ5
aNUZrCli77UnWiM/onT1y8DDgh2RemoE8Otrl4mp7SLFsNoHujq7xx7F5OTpz+V3
`protect END_PROTECTED
