`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1afbwa6NTQ9iKUA87ZC3Oi2e8VpJ1wLtZWgFpteJ3d8zL
tMJPcPRwnzRQNcoF994sJNNT5u5twmr2ZJS+D6ap13wxjLv+gmqlEgOyZCtfdnu+
Q9CvABqmLoGYl03AucyR7iKXOZ3kXMYxJxeEFUkTiY2RfV9fkiBQRMnj00TFbAHE
cjqMGqOkvSIByo1eAdMeu+c8pcD4tCZWth4WZvb5vX2UlfRcAqlccLkD6OJywNSy
e6XR2xjYFc+7O78/p7D9/dNyzmN7gkqNQtHLYl3uikhzonbeUp6CTkFLPUtc0Vr8
jRtVt0026coufs6neJpap0475julYulZJzrvBROjR2neacwGhQcZGeuSqXgIf9U/
nj2553MuHcvaSyqzQh735rWLCTxsKdeBuZkzUm6Slxqnqdkfmlf62OSSq1fssFKi
9PAkM5u9nSWTnGZOBk3P7KNWY0uTIJkSZn2PoHafUPttzu27uGe2qsW4O/rmNJ2s
msd1NvFONWAFk09DHDDvlqFoGUoWprFzb407OEYRy9M=
`protect END_PROTECTED
