`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePYUnQLgWiEhfXBNas9rvuCI9La9IA2oHsvSB6c48DSS
3NdaZrI5DdcfqSFHGjl4q5mZNTlpncuWONcScUcZaBMJsB/nUOAiTHc/BrzpqrEi
EbnDzlFQ7KneNiZmKAWEz+h77uxiC8mIqgYLui7JnsqBZbm6H3SBY2ejjiEgyyx0
VjRN5leqKKAB1bg2zMi03g==
`protect END_PROTECTED
