`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJp3aK0FUnYdO7P61gBs+VJdjrxpjGMxS/IxsnJ6qDmp
n0JCp7bvKYwAvttTaiHfG+zfDdbxHqJXAswnCMm81tCuCyT2LipvK9kNtnicwPN1
ALpYp/RrDrRJv6KcE0yNp3NzD7m/ELU0C6Hoq/08eICVackj5+bLzZgaSmAHwSVB
CCwRZYBs2NezyB46wkQ14Gu6mI1fX3KuZIdftRB9MeBDAiqhOMTB/PbV9FEh1i//
1kpbHOi4u69rHZRSp/ZCwb4uq+V0weH181dDgctnthOJGvXgPNT/1cCANilIvA6t
H1NeCtVJo7dtopXIbnZ+pCQZwelcm81sA87bRbvZsgCTvoSyZk0FIfd8qTihI61S
Pa4AhrHP56nVqJWdHyIN0zCJvoZ5j9KxZIYQRyWt5UVAKoG0q9LRQc9XFnbGI5Cd
`protect END_PROTECTED
