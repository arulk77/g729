`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBbJX+/S9de2edxOw18pMJZnAwRvfmi5XD050Lv13ZjP
lkcbqCYoYp/4PXS7+zpRl3+y/3KpQ38u9nPuTnY282MFEjhAfZjV+6C1IJbuBAsz
JTGoQGz30s2jk+i47Dk/6sXR4otgQK/7QrNy/on5mQbbGEu29dGjEM1N7dVq2jY1
7HA8L4QgYaqy5+kNchh3nAlTrENc/N3os8PCzCgEc9O9S8rDUKwVQIGG3v3RnJuX
RsBR0RbHY4ntk1fi5L5ptQ==
`protect END_PROTECTED
