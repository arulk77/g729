`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zYs3n99/Bk4xMjukODEXEolvIdy7SqofuNmGN41GRmQ
LmkhF1sFl5XKMKjLJcw9LKUG21cMXwqjQhWidg5Sh86zJB5iuY1B83NLwpU28Tqx
xwc6F/RDzsAj2IB7ZlSNhJDr+LJtkF34A+3sz0zfjH0qdBJ1HG9OEYgAA/tK2z32
qtAppmP5bStVjcBlQEbBwCLZtxmGSjSbh2TJ8DKgfWZ99mBtY9o7SZV6T2Nt/ZpE
d1QYXXil8T3tlIAJgasBv7bhFYUtKQ/MNRx1eqYkHszyWPROtSxC6PCbAacZU302
WUc2Tg2KKRKeTNyOp4U7MFl90+IcvhoZaSOjrqfKVW9e8h/nuNHSk9Ie1l1EPKvj
DQ6cI3FGWYOUEvbZ7xn58A==
`protect END_PROTECTED
