`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73CzmzCSDW6o2H6FmDrNe0FvyA7137KhvQWzvSiUZw9sBy
BzwJnmM735gg6Lt4lxh4OrxLpIKyWwR2ZaKxq9MT5z15sudr5uBJ2SDgpcjz96/R
OmY7q4CSZXDrfp4gBI188+Z0VDHNNtfguo5vJhCrm04Ikw/Ed0NV4pDQruVAWgkr
9ITBnhpDKcOKdT7mqODu2bIrVCUYU3RQxdo6phVoOUMYDaUe7wgOv7uU7II787Vc
3MD+pRePfVIBY7LeZ9WecbHO7W8DjpTwa/rHNtAz+Xi25YFO0EnQzGNcZc55VDAN
wEeNiWXZC9Ho5VsEUCQcZ9GhDJ2EptHe0ONm6bDmUg5F27PKJLqwMjO5HZKRbnQJ
I0asE4UBnsy+L/k/AgU6q3H31tWh4CGzq+0tguOoyImSDLsPcRoP246tYLABXxOK
2P7LNuowjQPgpf1dqsPpSM9e7AVo/22wRjYHDiWhxdJ6FSmDvHsQ9XSbcWIwCeDl
6F1F3I/GPvEXJVTX/cwisnN6VEwcJdK/cO+w+2ipCACoUaFsfK1jR/G74Ac7dS5y
RxR+WvYDu67R/XVy9nqJMfcsVJAu8OxwgbKbpcEqC2hJvFEn+XHNQQ6fea4KJaio
tUCEG1ARNiC4ax/BXQblukjhrGs5OWgwWd+83WefjuMjgjAhLBRqCfH51GYi4hXa
t4N4i+whp+PxMorP7LE7lVb8Wz5kefvGp66E1Oezt0EzylFNUhczLNfxHN0/mBrV
c76M/UUuDz46TQugnDwoJb0wcU7dwdDxkYuBMIzN5bvpmPim7TVEWKn+YoR4p3ox
mw7Mulh+mQoeFuRbxriAkFdccqWZWUelm7WKBAJzqO7bPhwcERTSt8kHApynKdKj
tZIWKNcwMTNaygymqtQRlDga28nNoMZQs3KEIS7fArHo4HJf95O5shLxE6KEuIW0
QWd9pjF4UvLziQdpROLhqN6fHoJRQhFXYEk9MM+YnwisWOrOCGnVBfHmEzPuCGD+
ReB0eElRx5eVg7HsqdPkYTA8QjYJJ3Ao3o2RyqQBy50YKZsy7qc1odevQZlZ1Zm6
UBLBmRkmL316cVYwsmu8MEaTxrWG2oYPIC+otc1BlxwDwRygFSn5TuO4pXSGZsM1
cNRUvzvPhD7mNAEKFG/iSnXGzk+pDNgT8wF+256NmtV34sZ84tNcZxjEJQE2b3mU
p+xCKyzcIv5eHy5UrZeRtxip5rkMLaqsveNMPekGogXJ/RSnW/OOvVqEyQsCISay
v1IfxoyuncnTpH4SW/aXLlT7xOH3XCt7XE273g4MqCC4d/G6IvhbBLwFdktnn3Ir
dR/WHNhPujY2ZOtCMacKGtUNO+ERN8R/dy7uYREHaKjwEwKreJ8SPwVRjbI7dtU4
IA757V4QWZllUuk7aDbbQAibmsGTteDuBNZvhHDUFiMbSFJaKKxr6szDXbYh1aZz
y/dDgHDpBPS2bY19hxSmAAW6i/hx6236waWAx/rPtG5DB1dE2ul8y7YaoKA+jjp1
v7Pgo/SDn/0SGbBwwNTPXag0C4Q1rOTywiz8f0PAWuw4pkBfCXHJ/f9XVrMotpWn
Ax+hA0yOmkt0QlJ8DaQxK58kXodAtmKTFDnRTh5GbYQphhlZ3D5Rha0C0eSg44bT
gzL/kMx4/Y34Tl+ZutShU89QK4ZXfHnr5+3LF/5MChzQhf3h+V3jWjr1t235CdRc
2rH3fvc0/64wwSmzVHFhggyk5VcHeRyT5422H2WnU0cagyNzN1YsehidIlweRpxm
UVHH/LVPjmkI0FpnTjxgMXlnPHlls+BJ+zgi7VhV5XjBqSZbLj5r/1i1frw0qgNL
bp52bIe2FK8yYmaJHUjScaqy4ZIASxDGvNc6BXVyu38+XomwzO9nw23n6TVRH73P
1XKkRNxxlU1YrB8Pce/30+DkOG9IinuOHDYHxA9ISgsxHMjqQ0M1L/4oEd/Jluqs
U2xjenHWbRSiLJsd75l0PbqA5vivmqeU2EY5B7Jl43Pl+CI5j8/yTQY94eeOVk1t
UvuOiQkM47VqOatuLr3QH8Y/k+VYxz/mF/aIv0A9mCxRFwtKjto+EOBycq/WnBe5
j6+aUpjLQGqhNGiK+tfl0d5itCJyIpx2WLO4t11xHU5QT1xe1K7Vq7XRpZ0u2IGo
iPYvIfzjHsOvINQPhs1uECIaTulF2LNxuW2cLwB0VsfLPt0m/1GoINh800lM0701
Z/Lc3xyhusWSm9ZoFxrxwA1H8vdALrfpsq+oU7+RYMV99El98PyhkUBb9LjIyRhA
997dTEzXcNxPxCSei754TjKqzFFiV+mWv+UCOcv0Un1wQ332jL0RoeBonuBcO4KL
1Y/BxdWd7poMI8rcvslFWi4zN6uS6QV+nYqyR1dZrJenONCTo30w8QUzLrxLxMRq
uNCYVIoVZmHx+rUXkTqwulFRpzamPcQmzLL8Y/q8f3g=
`protect END_PROTECTED
