`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG4WohdzTIx87oggjfA6gcpdJOPfIml8sqbQyMHkEwhZ
xn1RkYumtZFnbfdfk7kbKIRXko8K2BRg35Xf8Emi0ovxFkn4AmUU6rT5oWkcx/TZ
Xw9RM4wR0XJFH8E/iN1Nb6dBKI8EMjkzK9mM7JxOKlAxV+R33otxhGckcB2bVKFP
6CsR26UHPTzTqACDJGkAM8YYF9+5kOB/hjk+44yUya4iozs6B1hHvGZifzCUZ/r6
LlTRrugvEseCZ2GRc7equj+lFfJ8tR47s+XM7pox8kr2h9AEhOlEr/yAzeNZxYgG
SQmwJbYWGHsqqzP32qQtzCwmv0qyLLgOkYdzB8fUhNuPS7dYMXwgUkwY6EuvLDbp
Nezm93XzuOtz+8oEq3zzxrh5LND5mtlyIJxYboT2rRREENi7hsjImFOBtQq89kvj
5QEc6d9inRVn8LoOOx68v5BQWKKHC1rfN/gSE+fsKpP3jWR7mCAVVA3UOXgysUfm
`protect END_PROTECTED
