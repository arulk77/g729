`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePM2QwkLnUBhBkFCQqhZkq2Gh0ZeW20w5Slt6w3SVhtr
Lc6BxIk2KvPLvYbhbwZKoVxIIX4KNI+5ZYfnX6WfA+vBFbOOwyBXNxo29KTVQcQB
OfE9sGeHH3+G7XzwzSfaMb+nFWhLRh1xz3R04rZJrunFhd7f0vo/zPssbnnm9q/B
XZDDoj9ECmAtj2k4G8wboKqhd0P1x361TNZnDyVpiHV0o6lnE/cD5K1iw05FRdfc
FRU6oE4zrLQrNsm0sucQfHQgXy7iwIXsnzY7jEAzjbVOcmhlT7Mafz7mJwDqi8WC
bEfLJtEMqjtjh0raJkh8GjtiJKpyC7h152fe7AYNf4oOs7d/jEdYHoAHz7BAkN3Q
CbcS65RjFFE49LOICPf+hrYj+Mj75uBSkBMkjLKq3G7xKeD27W5Seo4xRDcittkA
tMkyP03Xrgf9qpgA33dW85sdQ6DgL5diaN5flbsjGgLzL082WYhXpHioiP/pGQOs
vEk5g/pPrSO7tTsscUdyP/IDqyWP0WJTt5Gmw5xk6GU6gVCxrpR8CjDZt3c3kiUQ
`protect END_PROTECTED
