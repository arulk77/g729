`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHvaujb60HAtCQbmeS7L/JpmuNi3bivaZJpgD9lO9IsM
R+V6te/YQg3sZExtFdfO/FffDrWNxEceGEo2wXyHfeOfbz/uxhVBnO+uPA2w0kZD
0x4xZX4Qs2Q0M9Fqnp6uI2mbCZXzRUkB4JMiHAn39v7stoZBROjVJmCTpb5zRRwo
jzFS+ifiE1txbH9W7Z3lc32LxpDYS9wQlh066VsQLMCfGVd0SBb6wFspEA5N7DLA
PUsN4vhu+6lq99ysWCWyaQ==
`protect END_PROTECTED
