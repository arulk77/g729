`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
fHY+RByhTXSSaHXeCfbRt7SgOlEigYTQtaHITPtm8kwhmmbAUfkyByeehd2rj52L
67GP9qyQ5IpkxJr9dSHSwPXIbkp1/mftsP65y/EWla2ImiDYkV3GKaaqvPM+v0h8
Mxf6r9h5VhDY182IE9gesBaNNBogNXTySY234VJ0NQAE4WHGWBeUA4+tCo0E2rec
`protect END_PROTECTED
