`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCE3bpl4Tid9JAydf30K7UKTKVi9FCJeTogMVrkbrwuR
bQ6L4uc9gIFlGJOHbbNFtil68JZvUzcpbAMni55qLreTNZBMlV07ph4qib/8j/lv
DVzfLBL7gKOIE8Bjapxs0MBzNzmMKxrEtwWwCxHcHpOU8NV+uhBxvLd8zxLSpmDx
1EHr2mcXX4NZR1jEbmS85gQbWf9/S5FboaNlARFsPG/TwjFyGfzGyo8k6s1ehTGR
C5nvgwqrCpLCxyPhEjhWqw==
`protect END_PROTECTED
