`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCZQ4YQ+zqP5hph16C73FPJYFjGHYMnTpSBJYfWFE9xk
mRdri4iMCjCuyo3qwP75BrPyBdovCiTgjDzUyvYMqU+zsLZmPbYhVwyAzJnm/I1s
QTuZ2zT/Dtmk8XdfNIRpLQ/pBwtymUkK85vPl2kiw7ZSedid+/zoomjjKsJxdrNk
s+fHHa2wiAx2Rz7zSuNJm7Z231ECLKcSmR08E5a3RjTun+4W0HRtQU7PEm8ObrRQ
Vg2tbWfhvTF6cVFXDx5eHxW1774yR5q5LZuNzERrDWA1/sWt1o29DJjou3bp5ooQ
2/VKXGdOHFo6LetGt4qQPrCHfT2Ebkjfc20u7uGBwa6Z2t44qLIjBzCAI6CYCssC
`protect END_PROTECTED
