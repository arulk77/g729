`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDSV3h97Gfu5CoozaN8qiqlnf1iTHB/Wzt91roFmdtA2
DigojTnhoPKedvBYmyCobPGX6Grk5W0elfkE/UyjDZes5mvzbRhwWPcsbrvkd+ZN
iEeqGngKglfe4MMIFD1dvTZaonjRV574tUQIqwnPJqZC99QSLWPf8H4ePKdM2liS
XHokTK9B6JZGvq66ptpETNuqUOpNVC5GVdVec9v7W4B9jrO1uVAI1cvmSVY6EEdq
tc9Z0beiiyV+BHv7lJaFlQ==
`protect END_PROTECTED
