`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePlvCP96HpV8UtXeaBCI0S3r/5tBNjTymtEUJyL0tx/L
9ezXO7sqsQuJnnx45Voa0jTkcAHcSi1z4VOGvYiGbyQC4hwMZHmBNtjVD7W6hCtQ
yyB5bn8kmv9k0IlG6AGAFoPFMqBZXO+/EOFAWbClYN7aq0NrrtmzSkLcrSxNKxKT
ZFk16tP2Cl38BSGD1i/j6lr7SKq+m/2KVrXZ4CHurXl2WzBcS8BZaEL2QI/R0D/x
AxwufNOm6+LuM/4XGzLrjdWAErR6w0nbSAkrkcG2C5OpkeZs3fC5sS9L3cfWu8Rx
pDXBu0yqCyk8DD4HAreDedAI0wBXcaECIjZVtw3uBCn6Ekx8PCekrmMqIg+YlzCX
`protect END_PROTECTED
