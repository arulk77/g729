`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
p8qgxFrlwbf1VbToxwhSA9lPa5Bi+38FCOZhZeMGAY/gdOuyqsrGICRpHtJAN/qj
vLJrFD1lPwdo7ehXfk0kVG15iJfDSYEp6+ldPWWVMLCXaQsLB52M9QpxgubL1BCK
x+h+Btj5n3aG5BW3dAp7J+S+HU+ZvnJnyAP4a4vkq6QbUnsd3FOTMyfDnig3rj5t
3MIW0eD6WavUg/G9BeqRZAxVT1dnqTcFhFSVs2Ba9OKXc1WRBWf8Q/NDMDUAYkNB
NRseqpR0nu5jrtYQpqby3eiXlmdDQtQF82CyZDKdam8=
`protect END_PROTECTED
