`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Dgo1BIlaWY56ziELruyh+nIfzPbrxMLLH/kWlSSJ2hhyz+RHTV0drMs80v4qzf7Z
mkC/SCI+Loc/eCnbt9ZWPm3QXegc8Rrdt1YxTcf/K7yvGEfRIjH98uLciBFMhA3B
XrtPjAeSIQurqw4i/GV133yuZE/erno9B4viDnB+smrkrb9s6U8hzSUMkV+Mzvhg
HAfulexPkERDqWnTRwtw4VXAzqEf5uduKV9gQVBw0P98k7VMHeZeruBWQtpnqBdb
fG55NIROuYcC7J3+fXVo6pG1LHM07VG7mJAzDlbrb1xuEEpYvnvSyU/OhmSs++W3
E6Yh7rbQhOaJ8ccPODRl5hoefOy9IVVxcCxlGa6gNV+pL4uwRAWxxSF4/Criqdg3
tbVzozKAud0mtCz2fn85Wutw2egzUD4JDC6uO0IVe/0ou30LDiYfeXeiOhU7DHkC
63cdzX/OhnfOUwjzywYpMjGLe4m24ddocX4AiDdtyusrpkVlhVJxfwwK/i0dvV5x
4IPWqynEoshjTUcMTEgqUxxScLmRxRrlM+5riC2iNM7QM+3SdfAPciYuRR2xcg06
R5soq3neIkscVYWf+fC9zpSuQ0cSRBgLEpAHNnGsoUBTg3tuT/Dsmli8S95gvsJ2
E4uifpKZ00lvO7eKfNM7tfMsc3F1Fy7F8Xuw7QsiIxQ7b2p7NaWceIEWJGKslJBz
+IBZrrnK0zglFn2C1l6U+9wadmJcILNwkd7mCCutqBnBTJmzOZWid98ft66B6esS
auatE5bb5Oup+UHrzkJJ/SyrMjriiT9SlzOnAbTJb9CdBSKgrXRNEQ6hPVOltji+
BmWXfXmQEC91ncdyC3+QgptRMN19NWEwz09VEu0KWwSyFJVJd5msFCBure4SD9C1
`protect END_PROTECTED
