`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF24THtC9DOcFNu4eb8PSQ4Txf8IW1Wb2iJGYu1V2yuW
VZYXPKu+gzP2TAkIG7ycwvMn8eAZ/e7XS62Bh01HoOiXjxuxXfJT699QOgt40B4y
lm2W/8BXAxAMQXCKXjULRl5JRWUj7CyNi1zcil7depxeU5cfYRHG6gXLjP21J2YL
c+CN2DCPYIbDeCOhODClvKYF4+YuxgKv3JPyIG0+eqU5yLxuiDZ12nq7SqlCqhxe
tckgxhQUwOiuUev49cvRjz8/lPMAsk5xRfWgLa3a7B4f0FX9HQUWOQTWcH9EXJko
+xRWv5gNTK767AVNFWkUMx5o0lpvi40DH4IrLAhQR2KmvyOefc487hbdOGYYn505
V8Z2izNKwdkeiIdnpaQ3oQ==
`protect END_PROTECTED
