`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDARbAC4dNiZ7sv2sdDxMf0zayG2dEVwQo6HL5oGHxWcTl
KotXKQzTIcRGpf011XM/yvYY+JWYWzp2IgGIS+tTl7ppiZE8HQPN6obDr/DEKTXv
txkYrYtp1AT6tcwiuTHuny2F8wCqdWlJo98coKCijaIGRAK6fa6ai61Ao5AMQC/S
1669Ij6IMqXd8M0pw5vX86o8zJ09zc67LbxcW7yVNx8dEc67BjGVNoiPmVZ3PqvR
zDwrBlowiKrz9AB+TBO68ssn4lelwEAzscZb2tXmxM50tt4OGDfp4gT784nNzibC
mXwFInQUkV9dSMekphp37y6JMmyQCymXnJI3gB/5ml3AOwuPDDoFZzJk0oACQ8hZ
V/irv6rin7OmirKr+cOI1NuP7WXWBLeNcgulKwmQgc6/T8fUlgkmp6FghM0RVEv7
eG5L6I+u/333uX7OuHj9dKoWA/6g3YtuQ2yenWyM6MkEUWlDKcRCC5W4CF6ngb1K
tsugrbTv6FJtith9IejuLlUFQFZy/anwdcmuQHJumdQzohsnBca2lvp4q/M8EmnI
jkf2GwPUtJ1mewopCxJMA6/uZX7jr4eK9Q8md2u9+3+IGjYbbQvIqiK8XBxI6AMJ
f/1chpLyyDOjxkrKHf1+lmpWYQHtKkgvKARFUJ3kkN1uUYD2eym9zPuzuUWX9rCL
RgZtOWDovfRLSqY5nlcsNUsmkGlQevdvoJ/LNqonnUB3oEiG2h/VEdCRsYbGHQw5
1DhN0nmcM6L1Y8YvzWtxsKawL/bahOG/UPflT4fjf4XsJN/p4+BT5HOoI89KN3Rs
C8b1Hcj6HFq/uQ/LKqEVZOf0CUSr1llt6MHVtuObpDohgINCDDStO1hOBCzYWJiY
16qsidrWU/MpuIyC+uQz5F19HiKPhLH4jFjCwz1FRZSy0RRwGK8NkCDctOgMpwJ3
GhVZrDrdZ3qZ2LP/dIDlSE76DWb4oucij2Vs2y9hBmgUgPRHnZMpJ8dq43lYWwEp
9NwYIwxzatFSNBKwOrMvQQcp4Vg2890s6n2tawbsu8V+WwUGympDWHYnfUcbWemK
+FuiTEXpyqowzpqzoPsFtd7r/Qf41j1uRRnhBaUe/oOXLSTRmgNUeFfB8Vt1lirv
BRKSN4KD5slx0/wNnD7I92HD2233cM0TQwUYX42B70t4ghs2mF/Oc+jldCyw8Odh
mhmbrXCebDlgYTE8uNE9x7i5qrchoAEbSAwuKBJMb772AD18coCPLmGcHliQ4wus
hTO1gulNvY3Stx8pZMO7z5H0s+VWUsqGQ0mnhZwpyIPqFTMS8vsC0Dk1bmI7o18V
yQf0fQ8yuT5wSgRuIt2iCPnmVRynz2caI0g90QHetriDRY7DeFmNHPF1vDd/ozhN
nx58Er2o4ZXNIbhKGV9GgoYacZwOoRwxHklhfLdWePj01F6m39mg7XNJWtYyz+di
FQtZqppxnWnvJ2szGCR5vJbb6LYEXQoDkRuHGBgbPPuW0K3lhi3xF7HAUGBdxSYu
wlOT37pnEZDDdajyg7FXyzCPzin+VXQU4TBVnVnJHKJxSlStxD2kimZXYi8qe93V
zPrGs8zHEUeJAdAN8l7k97UrkHRp7JMDu4nmEm+VvhOdlfHRqPPj/iiEnfAGUmuH
H+nJ52WPOaca8tUqBLi2zCLyDcSpZ6Lz9KrcoIhyLpbsrRbWTruN30hI0/twoAmn
ayuBUB4qdQMxas8KU3Zu6t5eZxW3/u8kggMGqZW+WkMLoErB7IRKgPIq0pWlB0HA
x9z8nVwF8JDEEr6VaJoCr/Mc72Hnj5fFQuuo5ZUX9XqB/48r2bx49P1fYRJIpoWG
TAId6CEMIkgxollVn24txXz3bwRo83C05hoXcfZnnqXC6CHHQ1LceafoxILylw2B
y6GCnPcVEroB7o+OvIr+/vyUGJD1Xz78XrOeRg3DgU4YEGxQMLMAPO29W03U425g
GuPTpR7E2U8rm1jNgesMra1mfHtwDv5J8gXS3QI7Q1xkiH1vHElYf4nSI8ZCGxOd
nb6iUOH6L50IaPgXOT7sspjPPTyBRkgKhdjK6wvgSP9x/GO7T7tebFqxKeQjVbDg
+tHpQmIIjDKR5ftnGysyngbeenBlg8DzWVjdxF9m+jNVOYVPst3K1Y4EUQh2ZuQF
Q6dtv6EHB5dBz3eHLQfKhbshpFG3TKN2k8vkO/KZRSWSKr0Wf9kztibkRRcas2Pu
aRT1UpCAwjIX10tgiDxnup+afwsbOYDJXn34gqFwVOgrcS4y996d3DsGiBLMPi+Q
GaeF5mi7WBMBQgEhfICRCTv2wiCqS7Z5tx2FpDTu3+aOyHbapNvRXb1PPK6WZC63
u2zwtSohvD+Q7gvoK2GWouqziiJ+V9/fCnreCgmvw5gK41/AN8SZZHFyzCKgkPNY
mMX32MYjTS+LsWJzy3WIzhLYbOHdBXHj+y9ZelDUJhFAB1rK0yxWdW0gUdeTmASl
FX9wXoTarBzepeP16PbwkAnVeSGbEsnAjRX/auRQOdNNKpSveErmx5yLsS0ZMtZG
Br+1rier4Jc5NUiJLc7yVMH3DnsB4fpL6yGCATnGm7eRcx7yNO8ZdwjZVqNTCRr3
S0rj+xWp82ckdIe+mhGkFjFPDJr7uKs3vF/CC7JOlTAYcVwSpFxT+hjOxo4DX6r4
3+1ejDhD1JF68M6/FPLl2QBe2cWlC9hi3OLFZnD97Rhbf3tNp+IDQeapewd470Ef
8iH9YfhJzJCwHx8dm/g0dubYbodlJ+Ub6fWh1pH5wHw+f1FvGXyMn9iciLiMh11t
GO0u8bGjYvdwshnMSxJCgL24dcYhxMT08vRoKHCfRzmXIugKqyHxGTmv+8wbYxV8
H1JAW3xUPdPnqhNTAvNkVxmu+CibSQ+wwq+JRtM6NJLoUzWwNEDsQHbgY6BLGpv+
+A85Sd2qOO3zZ806GUl0bnbwBzZ2acuxpyFJhME7koJwKqCttH9denU61/SsjvJ+
d8Ggu3i8vy6rtL5OKyOiAFfds71PZXBuE8S2ya7ulku4V7LgNuy6L0ZKmknSSh4m
aEeHz/Hc8XIO4hWMkQo8yd8QuDOvVDj0ZhDdrrvNtKCa32FH2Ki6ayfA2dIr9gxV
a1Lh+oGBk3sNxPmRV+YYm1bcsWTzuGAcMO6imGXsGH0nUvy0MBPfKbzbt66I859E
o3DCrsiXAC5IJUMiKc/XfAFL5qTtcI7m6gUx6jt9z1xQRV1+vGuA/EeL4joNwM8q
d9b0bGDi8CrmECC2xm4ivRF3sRA4OdL2X6TMcaYaU1+FA9LYt0P8PAd8G8NWpbUL
F0HdrKyyXmIGYMGNHh+Qnq9H60mH6vNnNzBulAVatJWbbNDRV7OHt+J7hBze48bv
vt2zFAvQm0ng1dkETit4tWEajl/gIHXoPwLzGNceicDPoUdi/BGCOdFH4Sb6+bu0
SG9kvWuNBq30qlVxCR65+fBVrPx4+H1lL6YYgg3Pb3VxrfIdV/exWgRfRTSSFDrR
BLxXa/BdjXoI0qPq6maQgNoyVN9oAnuByxM9PsT13kGwgV+0qWXHCgSE8m/rz/1W
KgnaNSGDYqrPljV19tggj8LrCoCIEM+5Lowo0VCda0hUpz/U6NaDmedCTJZ6l3P+
X2RH+W/J5DIjwa7u/Zcwm1P6i3T2CDk8v/UJKzWIXn/XCElM8HTUsW2R/rRCK+yf
HqnLtKw8M18wZtRZFXEw03Al9uCzN6/PzJ25i4BA9HYKvBNzPXQ+AENoN/vOXUTe
7pw3zFCVRLVmkYJQDlB1eoK/IJoUhYDDtPo4p9XMx8YC1s0JAlIf2BvTpkpPQM9A
5wUC++o2BeCG73d3nIAAhdMyF2MWtyBfgjhf1rIAQl2CrqFJrXlWwxIL/f+pyS3U
eEyHAvcohx9EqJlLWjqfTSnwdPqqTpQf2rb1PY1EK8KlFDFnmcOEmv6TJQNGWxTJ
QuQ+uod/bMeTjQ6DlH9aAHJo9ohABqczo3pTcWVDruzW2Xp45KYp9VGvkrCcxNdt
dUeX7BfuAZjXBOWXqA6t8XsUtHPhStWH96+unsm9fWfjPjYecHSc/PWtq3NUnGwP
a51CJkKNXAcgT3Bqp7f6IOdv7OiRoQTg2eztOQdDL7HNRsUhyn9cSGFuI1Av/WVa
s/C96TnBTfmDa+gnc80eeu+XOs9p5g69Lz/HD13e5VLaXjGfNCMpfWCb/fAZIN4c
jQZh3geA/49RxMRcy9h9PsdP4dNwPjukfU+PJ52bJhOGgNiUloFIrlnXq/1A2vA6
XPGJBvZtVJG8xC05GDXRP54rDjmjTMF7tAD8kf/HGHL/w3tlvar26v/zFxV7M/f7
tl/ziZtgnHD5qOWvjSvCN5DHzv5o6cE0PJSDKtKvWQE3Zhim7uoREZWCIAsKAYv4
TJVQeduH2tWDtl3JZpRlG0DgXZBOrQDsCn4McaBcP932g4TA3ol/NrmFwEvL0YXs
BQ8UshBx6eDraWNP/KPSO8m/SVrzAlSEqoQ7S24QkceXfOwPJJEDw3uoUzu46ayn
yOO9eFln267CxVQJxNR/deczhLaTeT0H5VETqj/2sdzMDzZYtHYWba8XbaGiekqQ
b5Y6DF1OroPfovNKB/rl2WYhNDZk5xyggHzzpCojKi506H5QBVqZp+LqoKytHPKO
C+fTTSQRxKmKWn41ICyDS9gSzXS7IgFE/aSD1Vg7K5M9bWLVK9Y/1HSkELNhh8Cg
mKSnVcRF2h+rGIKVt5vpBCNvjkWMPF5tkzVqij6EzsrUZL0dUhx6hogFwOdhMrrY
CxTeS3AQh1G3ETITrfFJRgsAmuzw6QV2HOfSKslyKZj3fekeOc2hX8LYdv1qK0rz
OeBkNREm1f7D8abZtw3M19Cfh9dfWR+lYPYUysUaTVM8clLhFmJfgWVYra7vu+4H
Ye0cxZZ/xMZ/hhVVoXycrF6sqZiuaJAmmKWWm74dLFObRML7mTrIUqTARXHhlTdI
/nP5L6J+goFZjkzfslxiwlhAbd8Bh74szUMbeAT76hDIoFROI/2kiRNUu18FrfD9
3zqQWBN6dvwHKC4Ad8rAhWcPGKvszo0lvZtxaI54ZFoJojUp3Q2Pc3YpmvajF8w5
0uGqy6swbjgnacx96wWiIO0k4Mj3q3HIy2vaef8akbCkmPiY8MTEDZYnQyDP50bk
U3oOyDkOF1ub7U4hUvLJu7H4OUmEIQ/vRltic0HzGSjmX6Dy6IL84biqEYPtluaS
5efqceM0aBHr/dCOi9DWF/ttXnz1S/soUAJHakqHbzuq2yvnhOYH/w6vxO9lMp12
92o94q/ianCmAvnNjb3YY9ecC19hd6+uwCHEDtaFIF7vIGT7smwE5SU2kSnAdTK8
3HqrRfjU/uHleIMeCEYTXAPbZW3d22qwd9CGSNn5ipCfu7kHTDUPCz+1gjsUyqpN
wpYbv9BBBEiom1vGh/yjz85vExAcbcJ2cQQJgoNm6LwDr5XWS35+nVjiuJTpRWoP
S4W2Pzfk2ueysq5vi69L5rXIkGolfhsKjBrj2sVkRboomzVOrg0qroKFRXEyMlxy
yx7YynPDt/ULAS/qY8azu7YCZaCjTeZus3/To0nM6at380e5MVc2l3SwVA8sY5Bi
TmAs2eOFpSJl0VognZ3C21K1lBBaD7R1rygP1rIY1UeWORaNdun8taaIpvC4ZZOM
VW91v8/tJZ36nY3fxo+vLUrDPrNbQ2LEW/vy9LHimNSo0YrJrkTgIWjd9rz10QCL
080ykyhtwg1VXtRy/DQo6TPi0ZHg7Gtr10hr8pwLzpSmhiflUaPEBiiTWyLkXzkP
BAi71UPNin0/16+PcXxA8g3mlx9Mu/8yai6Y8ol14gn42gxHkgcQWCF7UHjfCV2F
+aBql08HNH/NRYPahqpxoW9hsDQG/pwUC0qbxSmrWVGLp0SDIL+mz62G+XyZKgJn
s+W35xEhCcS9TVk1GYxgoLsh4klIIp2wvs5UpKXnMyS2+aJ3eplMOeAIwIZp+YGp
rODoU5/yfObGqw+V55LDPnGBYP36PLxHp43Zs3xAgroy4o7ECVn4TO5UM7QOdZI9
6GEw40x1pCRF0oaVil3e5/iLUtMoGj7lTmPFQIlXxICWdiaFe3NS+MmtJj9/MB43
uv9+mOau5qG8Vl3/ilaosCuutmg9CzbfcuI2ydLbS01O9VBGiUVyyO7Kdjb7mpQt
CWeIM+zyCs9lNUVVgTUF+GGLzqW+qzbophAr8Vwdzz3e/oYjPoo6Hr//hiKyzF7L
2m3A1AMn+b5cPZLVY7rkhq5b6g3xJAHRo/ycczOr/rPdv1ZO1dJJryQM3svLHyBq
md4n69X5Pyq07NVJ8NIREg60PTNyen9d+QjbJxs2Bj46x/XAHXk6skqJi5qbB5kJ
YMWL/DfBpAKHgPw1b728yDjs+67r9SvrNLXokkq7FPxvVRvh053KBWZpaWRlqSkW
ce4UxVwjuax3tVosRXOEuHvpMglVMeoQVtaFzV0glOYxD6fnEstiB5BLGIC/RA1d
CnrJ1mtPWvQREvXe/M9H7bC9cb5ah16ERfsD0+jRtQFj8bkSRYWoD/7bOOvkleke
LBNRGnI6kR8MhfvX/Fj31X6n9a9pnzcOqcRFok9vScAwSfo0fUcNjxxtd0Gl4g8+
GrKP3hBldgFg+T5sk6+11F8YUgEENhSHHt38iDbrALrefE5GLYTPOFY4Phuq+MDC
4adOK9UV+DwMTm7DfEyAL1UUNDl8NogvViOlpfpjN9YlXebbMhkRuMFgh5AJt/EY
SO/5uA9uc72lBUOGdDw6BwSJUmVS0xWQtetdO5llxGoGBAbdUOvt/5tKpq1OPF8C
vRfd/OCVzVIiX2HcEYhC7aPMOgpqWhxU/xGwGjAtAxJdhTx090O7byvnj8rA6UXY
jzv7YX7tc0AnFO8YGrHixxe2hoznqkiSc4jxXpfrRAW8250HGhFOYsjsnKOoEUC5
Wwd/ExJzs/QBw1MrCQqWq/wHm41EjRYxgcvfBi5eS2bHo7lBVg1V1r43vQBrcNMU
n2azELVj91hEQEN67zMd0f+LkPisX45QFTO/O6SmlBxHIT2/BA/2SjH5vmKsf785
ysnDTl5lrAK2wXJsKMi4O/UoHMF7ec6Gm6yoghmV+AY7zGp5kc1BGGNSx0RKD0iR
OCHDL64c+umRGZXnuKeY2v8DF+aPSqLWkjF3Q4280LX2lndj9to/bIDW0ltuORTG
yE1pDqRH0okSg5ahmdxcTpIgrafy6B9w5HKMr4JHB9ZjpEDHqwNCLB9usxGODpvs
aEVZ4dsaYAwAjWOHcYOjUs9eiVht3A6lYH5UrkT52IInR6tDOIPdeDYWqdlK4viy
V+ri2vTX9N4lAns9KjufnEETyDb+Iukmg4CZ1k4FB6++WLgbQYGN1x2LQ5GjULTZ
+5V8f7pXmky/rof3z7Wt0HN9VJVOc8+aJ5nLs6LBAgxyqWgeRfk5YKKRGhulGPNf
7T/xnI1OTc8gpTKehWv6NqINe8oRF7/tM+XN4WrUrKu8KnZmRRrxu++bMYolUVWP
ee2hq3aMauFSbpq0SirhsSJaAhq+sPsB7uMJDByAYIfhu/Wu9m8GT32sNWsWLmZL
478ouriSr6ROtW6ZQUgvhxYauQ7Pwfd0ug2KdNLKLvZgSqhiaVy/6Ib2lQxDG0dE
pVIomVjVTC51v+XJAdwaLGv0/HgmtyrMYjLf6EV1/XmbHL3q/j/lW9mOKaIqt7nn
EGNJDphJYv5nyxKDxA49Kpv2tpPlswGmnN/0OVH6JNAT7zBukK4/E2cFGTfwxi9s
pHG+H8mw5Sbflgh1wNWBeFj3OGzv49z20+ui2TWlyl9qUFv2MZuKLKO7DLc4xYLO
eHdfQZ9SVcTM0Tfn9aXkqtz0WtZErspYr743+HazgpHDkCYJRDpXUmA6bGFDT5dq
s9vxAcUspZdAtOkgzvB0W2fBVuTZPo2tw1rSCazB4Z6bF7LQJRQFUCEHkrs94hUk
5OXcEByBm0fkdKScp8QimVXow7Xc8hz2XWzQ6oXXRhtHEdDaod5qe7m2l81BXo+U
Tbqbxr4i6/Ai4PBSiPilpNLcOhmkyNRv5lUItqGnD1qlyoxsrhDiwK42dAzqfbx/
qzM/oVrIAUu4gDRdYSVYu7oR1L8iysfezkETLt5OnJ/sUsNYkoA4cBIO2cx/a//2
OWzK+VYVX851OmNn16YzwSi0MpqxVEcIQ5DDcK7kJOw6gFi/7WgiDKFggFYXePh2
NSvczSJ2BC9OO2hqcsy3omZiNQ4rVvUDoswgunYI0hZjTxv98YYjst+LF5x7gvSV
sbjkCHlmVzDub6ApHPCUYataMLLKfbcmjWgo1kEVMVynxATNtR6PsbfvuRca6+Rz
2iV6lOPkAHiwEEUBOxdz20Q3nFzmpx342pEOgYY+XAbX2O0NJgnw8MQEo8qKWnnZ
eyZBFLoU09yK8btB8zB0qXeXsWkwu7S+aCMSPAjdTh2PCyus6EfdEvfaVfK9kAne
V8idLnN0Yl5tn+48Pnl/iNNFQXFlT8M6vRXgRne7/Kyv5IU6L2C5sdAE3JpeIhHz
t4FwY6bnzLXy9YnHfB+8WU/JWwE0JQ0UDmQXaCq2qJwsM4T6uK/BdrFoJ3Ju2pEP
l/Q5i0UGX9EXhiTRLgxgNT2hxdqAsSn6fw95rCnZRP/J2XWuZqh3CrAtUPXT9j46
ewKScQlfRzgtnexEPhzAyt92rgGLlGEIV6ZSXeH6hoZjO1EjHjm9H5KiVLjBCCpe
QKknqjToDThjfytlMS8QByvslNgbAm22krCBzfmNgRBI+84EC066lT7fFuyuiyMx
ccH31/FG3m3sWEkZMNqvx8YE455Qt1BJDCM+6HimZwA13u7FIrGeNqtZvHVdNn0q
yE3f5yUKuP7qWnXEE5JND5l1xoJHdiX08a1EbGdt1Uhp4d2MgsGJBTv/62VzdN8Z
mMIjtLUDo5HePvSaFAQqzg4apJEV7iZXuXjIkBdVuZvbkKUI17Egjt53eJOnUvjl
rIaDkbkOdi/K7seYYGLJ4mmvgu4Sf6hzv6mbOzWKzBF6wv8tQTAEBkGVa0sLyy9x
Y1lohD4ijfxzvw6M7q88vFb9TDQ24UP8wXWv/IDOl5Swp2fZv8hiUK3B5iWvf9mU
/btB7aSCZAlrBOizIZC4TsXmfTGtcUfNhYT74EqXuGl/rRoQjjN7aKOhiro9qibO
aVfSkHaIm0KFdx1hy1zl/LfOITzglAXkNDFvrrs4Z2fiZAaTb4qDGPknHDtXyuyw
rlyqABoEFxeml9mmpfy96f1rvxXE78gKi9WF8GrQ1RRnk0kBUmaxLMYRtH5/qv2P
1D/ZuXO4GWaqySZQba7GRYsQLrucDiFXQh3MoKhWJv7xf41qqvQI3MjSvcv00d0s
R3f4P98tyRqgOnKvqdyeuwQFKEjT7Kca5w9ZYoo6Lgsk/9es1Wb4C5yQW6UF2iv4
b47A7ll3dDAWH7uQOLUesq5XvCpz876zhY7qXkcZC2nLdu5uKk0AsiMvBrm6yXwg
bv1UBw8b76Vz/BsHNHtzDWVob/VYt7jNXKZzCBkHZEdK1xYg2MtQ5Y//D0S4I9MT
Ch1mLhAG0A4bYA4NQu2qiOAD19nHiBlAv649BroViaPMp6o937z12uwFSOzzGiiZ
AS2i+2ikTHQfgwmRKIHYdwljwP8fDzbmBen/XoD7nnaFxZ521BzqF5C05BBRnPJ1
EyUPDdfd7fZFBmW09bFflBwA7LS6gxG3gDS3DUbGqghOkpCkXY+8sTZ7LqVk69Og
T2KT+vCvxjdNb17TdB2HvazQ01tyCsEQnr0JAm1oOv6AU6U1ZZBMukq9K4vJOJje
+SgrS0CGWp1oJTuVhnlJkQ4QJqNQ+McxD5uGFtXplcfE4/SnBlbHcoZOc+3RkBao
f/bJquGbOxt08e4TcGAKQfYJlZWjGYKWqIxOw0eqH/Z7cEdsq2KdRHDHta2b14lL
8XiPWztb0Y/2/AyQ4Oemp+VbIAqNw5bi0aRFo+sLUfjtEuy787JWAJyUsakhGXZC
JQYZXv3eQHdviy7IwuX2f36W/kAqbYOKJO/8DeOKSV5bhgMDWjM+aHAhPnGwAbs4
VuKRRDDrI9eaHw7JtWI/o6oXhtMIaju5jzy/yqyU/9DI3utAOM/HiFM/fhRexXfN
JMabfMwtH0aXSLz0GVN26gIOC/4HCPK8D5VnmpZZxe+A4uKtgJ8Sq8u7OPYEzJ8r
WYq2gL5oiCkGwERk5r3QurDCOk6CkHd3W45P77EEsWaGIx5ZUEDjo/8VH52ATQfI
dU4QpdZMPOl39iG6EnDHx1iuQBAUsovaahfQGNWeyw9R5QOsf1hdYPJuPfUGJ9va
s6sgEhp3hkgmx0n/FkBnyJw51NscC8iFiSDD75iaBNh5oJaT5DcRqTSykrX0vBsh
ZtkqigC3aqGi/zpWEHIsweKWbgpKZWbZT+Mu1hjg9PqabzyH1cpZ/99f0z+Usda6
H3+lJEc9eKoN9n066O8P1xpIhg2XXlFJ8pLfR4s34n7/vawDnSEY4fQP6mA15lCl
IWSRRnIO3dENfiKFsIJeRP1e0PdUT9Qa447KL8dck9SiwyovHJ4vwAKG/nXe73qZ
erYohklHSEeBDikLokaBouLeYfzY5yvS8FthnfG/nxH0WAyEiMD9OdHxaQiGSxbp
9l8HBU0YAGcYE50lTjW+irXibu/t/Vo2DHHTETpqbwYn2IC6kTMY/zHXXYcAv3g/
8r16TCRMDUrHNxSOrww7o5a9OwXWIdIIwOw2JK5XFHA8wSvocCQrvckldP6iHJB0
ZmYOpUmrquyy4L/iNjuETtsv1oVXwIkP59aq/bv6Yodp1GeD45thC38YCvTQM0C/
q7BA3FHM1++HJf2XbRInFI/NXl6PpTOlcDCy5J62uW8FTmT9GMVonoFeuIg1cq+Q
4q2bfIKdWXMVb+YAljeOUJVOtVJ72sLk5Csyzx3wVQ8nyYPZbogO6aTegNmLYwff
BS/BwYqEBAVMxhepuWw9o1N3K8Z/O/NDYIw3pdAgBpQJvathIsNomZNi6/WCCRlY
QQbLtlzCKVkddK4sCagJtLynjeYgOIxqrybyArbS90JKvA5OMGbZpQNL9xiOIwGf
VvRvyiuTsXK+1bKkMVyClfjepcs7OFSoubBh2oQXOuiSRgIKvYcbd9uu55P78OpX
GUTmxb5PWhyghbKBueT2mCmkf2615HkCYfXGm4kv2B8dFsdPXsP0za+/ey/Be0qm
p3z0VwBmRt7BbbuaepAcNpEO/V8LPWGEmrr22ld6tGNm/kTJEQ2SbD2qLyfMJtOA
OhfPb2qOfmKQIm8ekobAdKkrVpoAILn9mX3ry3yaUdDvccoMIlDiNX80oUGyFG2x
vk2IqWjItln6jiG5WUBpTrkfSzniZJZqq7ej2HHdFOKHCeHqXJewAib89r/m0Aml
jqnl7s/U3T07NmEi7MpKDEbPZRJrzhRgvojcdzcmXLdPqbBxwDka9atbK7pQDUcB
1FfQds5UlKsso6sePs7DyE64AKyUN71sUbhCOw+aYqsdUUOAozWHiOq4YvCvIgu7
d9SSdRAM3SsdQkEy4pDTWrZxNu1TKYfqbJQBZjQwp3sGABEgVC61iUwyg8GqI9ZV
gcQDR55TYtNRXl30Pf732lDCDDOkSb/MTMLZRJBoEmSAzUakPfMRk0MLv8VoPJFy
jvEcw93unTbwJelv8+CIX/KFWraGjZYnZ8uGFTfkgTZJb4Uxe6W1GH9Sh5mY78ET
Z5v3vTNG/I+CAhQwSbwGiECAPIexwz2dKZPaBKpJchkAOTWe37Fm7CkGznWpJvn6
yaNP2W3fy09bHtl0Qrrnny2BOfvrAFVMCUMqUH1GqgW5OMeJ5IVrOWzvhpfKacq9
AR+YLtKgsRb1fFUkO1PUJSvr7WVv7j2ht3GOvfyFmo6D9m1PmJimU2kstkNvl+xJ
cFVDWVUDu8AQY4LQoWZHgwgBj2t/K4EAlkWZsXztBsv7nPVoylYrxSg1ioU8w8IB
pAy2z9OzfCnYirBQBJIaxweSHtcu7lFjLewudT3bDjZA7qWzw65HJWqHxrmXnLWW
oJqNsFHxW8ubxzazeQ0JCo8Da/9hTMsmY0USP6loLvHuhiSaKTzdo6OGFWmAGekY
ESHQ2jKgLtATFZB2uEclFACGdRPKuWeNQ5CldLkokAITdUOo+siXk1/DUjg8Bps0
8NlYUqXeUDruK5eNVvsEj0fJX66cPJo7O/MxUOXe27U7/NZSnivWeR0LFosYZRAk
/mpyTdzibpRSwAAhrMTPyoAmO8FIRgRIZqJajWhRY5fC94zNFJIgW3eTzvsYRYFE
Gzz/SU3DepyI5leqvX9QSb/6WqK5IHtXX3gOjFGwd608VL7Hhn8M/Bxics7a9KPd
oHko2EmCp+lLEh3SHADUvjtKeUFO3v2fZ2q3mnvXyVWK1LEuBQerUzsFAS6WUEw+
XitWiamj62BehY5W2ciB68P6f3f9NlQ7f18zx6z5YO3AIO0WpdRIMJzkKujV0jd1
Z1OhfMXSeFZSj1CFsgOMq8EQmXfXt7tx0D+xgITx+qIP/XxIfG0c4hZy184ix7VL
V8Fhz5A2WriXq91H0OdFNmiclehdDYlLcvywvj/S9U5CRTgpKCtEfyzj88V95qD1
00nGtvBhbXswEoCR/uBL8dA2pjGDJFbkqjn560RTdhLjmWcD/HvkKOsqj5YqGyTF
JI72QYvtoo5wOPn+4yK66SIWAaL117Ex7ld7BzCuEsMWsT/6KK//bC9VvdmK2lLy
gn6szBECuN/5EqdFe4wUVm/s6HgqUfm9Xw4lwYimSD8ADE6zM1wIFqmCVSm/REAw
xv9LBu9ud/4WNJZj+fxkUPrJCc+/5bHZojfn7KZuJO4cKBrYZv+Mf1+RiswUz37z
9EVhH+EICsNwndHy9BSlXe/ogV2QLtIit9sDHpWnRdlfBQCA2FaZ/V1/AiFx555A
J+Fuu9g2R3KCwCFwnaOW5U8AltAL/1TBFgtaQopovmctm1WZeDsQceYd2PkN0/2u
nUzfQw4DGX9qy+0nFLtDOp0KZHS/g2xaZNH11gYfIl2qsq7SDzPVEVDq4/TjsGTv
DfcyTH1JyEU38hITPQJtmLq23CYR53MWyhJ/AlKKbXgRbeQFwkF1R4ujyIpZFxlj
naMS84iL5kr79JL8Xem7RhCdJgE8WSXOh+rKNOb25pPBhvCe28VIQkTjFO9bFgS4
pvsJE6+iZgnojk6u27dh2Y3eOxpFrtyIh11+E0AKmf0yYLSkHQevjOJ0saD8941T
F+Li/kL840OT6BdrmAYzAPfKwXqw7rgyJ1XLu/tCHpRhXzEosqIz4Rnn80ZJ28oR
bxL+PMOa/04mx8Lo7Dumrl1plKCizI6ecFVjpiTt8KXrKrrGHgHr7s+i+fgmJ2+2
mJhlYJwNrb5LK1zF+baekzdw76zxS5EWUYtz4+sf9vi7Obh/mCPbOMa258v5bqCV
mevTSkqXkelGhDapmWJFEG9AiYIDNNE/LrxDc7D30jtuJrW6ctljCUOyESmv8xFd
Ghq7pqx+XOkCzXs+9CorLVRJsWMd+gkaio57Ez9t+5r/f+MJbnIQbB41nfEL1OZS
gu3CaC3jakl4mQO79iDA8CrzfgMip9ySHk/SifN1kXmE75EgLb3HBHQW9TEjrPBd
46lRkOkr0v2tdoCqWeGkbBBtD+7DqHSfpN7h8idoxNaY3dRCGRfKOg9BGQPCcVl8
nUlTKgJyGZyukXQuQwrI45DiyeP69skyRVmLhwjLlbBDvB6jJNgrve3zFimG245C
+zM8oL0K+6dmWoh4fmtsv6PA+if5UspVSpKQDvzYud1n11AzEWqcKuuMzB925/Qh
+VmL/Shu+yLie2JZ007Nh8T18P2Dx27YerOat9M5ZaNEMfFiyEoLLM25GMLshclu
bRF8p53jqRTbVyTO+ohXrpXxDidkly7oH/2ceGL96XtzM4py5PReVj/XTD0AjZbX
gl74lN1Z3wcaLCh3tBNUxXS/e4z+owebZckm44Qk3GUE+1z6rCsPaH4g2dfd3zH7
mfsjHOrnwPdVXcBXwGVN/kHVvVI/wbVpHQtKKErjmv12flWOcS+BFXhVxU9yidRM
8MEbkhHUrRDmrZYalyvpeOKdEZBOFW7PdVEklfwyFh6MOS6viWA+7xWt7mTlYnmY
F7AKGe3m6FvsMsw+JIdYhBJUPSfjvE49vXRyKg9cmYRR9Xe5gYCmI00C6HAsvQRU
HfD2Prx9/nSBy59RKBzs9Uu1uiLZ+hx8r3W7RnhwQDmOEoEw2doDQhafQPg7Bf9Z
2BsQJkuHz4EqdFb8kdm8B3Xv6lLNXrHlRS6jin/RMOv9PxG2pMhow0TP+SKH1gN0
EzomKW5eT+7D7NcdO/3l+PF3/XOyz9E1wjrdqfOPv+PryArRpZTjXyF+2kLwNFxp
AY9EL8p5u85n9FoUqDeXQMlsvQTuKbvHweH39Z7LzzlRAc8WKJMYBAxhKFTFIhk/
RCsCaq4vas6Bi3QiYCJofX+zkI8iTvtf1M/ar9WZuHpx/if/fuqvwe4lRW7cejpB
Nx1rokL05DaOeJ5c4y18BkK55ACwu7cjFJeP4WP0sgS2NBAxaUFCmDF1cNgf++RY
KTsuf/gleat5qaY8e0gY9LcN+OMb8rmanwj4BKQXhcdrCUXyeBHNtkn4XRnL1WsW
kVqxQni3sHFYfimwH68OLb+Is/aam0N9yukf2wKzc84pSiPqsMsSfmhp/wDqr+g2
b/xPoJjWMsO161FwnCJ+v4/T5/NZLQ12yHZErDEltSFm2lhn2cYzhZKvJBT+b4Vr
Z0qE14XSKoYzIBIbSeSrjQ8crIHyEaEP5fu/3EDxp+JTGCcUAKQak8GYFaaQw4jT
5e0YDenwklUWh7fL84LQSY+9b6TOlgxkQL8472R0fuDUoYhCg2yh98rd9+izMxpt
KmdR1ghwIjfkKJoY/TJZmNH5M5Ea/WdnSMtXfJF4is/ON8WTiuFXDh9bG+BWBWNF
PnIxrZeH9w3eOnfQB9sRAg3IiGS4SbxNsJwi10SJQQQ9W2zuDzHs5Z65QKBgGOC5
fSQI+/I1sxnkW5fek1domr5SWHFujcDJVldynPgFnHWC8NkTL4Ar8Lj/41KNVG+N
Mwv+eRaWK7CN1Q5WB7P2Nx3Ay9HROCHrR3kSmySPLwWhn33Yo3XCENulwbOvcpE4
W+aX1gUBW+i7vPj6s4fSDiMwVtTJ55lup7K+ougKtSdZGwN3S01syLCV292+M9l2
JyKh4Zr2HPNY7WMoxaRF+hm+/zrnPAOzx+LhNzPN5tLdGlKLkn/Anuf6cg6Av3Fi
ZkTzNVQq8MkIhZwFI965hlszkOwEyw9K+AUYL2s4q0RgS+Ry/bNMz/0aaPdn69CF
2H8IXZBAlpFBvmAcxpF9pE4HXpV79gA6dB7lw71PMHh2fvWtZs67nW1Ke+pj1uX6
vIYr+s030Koy+Cj8bPCBn3stERSa+QKz7RuL/fP4ByncIXp8AGGYmSlV9MOCk7eU
mPFQ/yyQfsRVZl8FAyW8GQbdboELVgC8r4CPvrEl/V90Yowvj3mh9XX8qo3fk2BI
CXYopGasWPLeIV7J47Zf4sys1q6LSLUah9bM8CptT7dO8Qvwvz0WffXd9XJa6bsV
0omEJt8R02/EuTFwn+j7IqJGbJk1XXfFIqTtJHMhIH/x0f9krc2yMBNVy5GvdGk6
vgWHIhcyhpMNVJVJpjRIMtawxUO2kpHIjJzCZ4JKxJKuxfuTNFvpl8ASKow1cMAM
Ui/l5FPDgbWU5bYvwahovjkXA8KvFObOSie+MCg7QH0ewsg3kzmOzBkzpqIojbPC
pxrjb1gkun6BLf1oBaSCpyGtRaS+HJJU6YnctP4/yzdBXhWIO/ifpp9In9eLmRl8
VrA1hMIWVqvlEahNyUMGgvfeu/NZnlDMPMeNpJ7HA2dPyJidz6gm/e6PBXwv2V6u
wI74Hd0i3dCLfJZ/zIGcDpsSJYeTWg5xy55kiKARiwDLXQFt4QP/DIpSm+KfBQm+
rpkqta/xgOEbiEh1cAaXswqjJBSUlxN9uBeKWq3yFKr9GAynzVkggowTw0gIGQ7D
jgmjjJzJ7m+XGA6CxZWq2XgjKdzyYs/U3zNazDBgD+/FsS/kpqmQ3khWyc01EGGj
PTd3ayNe4vZLtLrRNKw9G4m67yzzh5knvj8CTpn2zfAI0NPjAASFUJSWyFg1n52o
if9B8iEaJDZ4wLyq7cZ472yFtCnqIm1lhiyf9nsM6zRYTGp7i1oy9jD+fYHcOGc1
SrC1XhgfQupVmHdf407Cv97wwWWMiqo3VO9s3aDGl+JVRNyiMfS7zoJOg864cH2m
43uOA3PlT+t345KlNI3CGKgTPmhCZsA42ELczXjJ/fiLEQQBq4fAqgE/LWBPBYmF
3bduX9FFOaqgzVtYvvY8hpIrTLpK9mMxBWvdRJRKsLZeCUTGbPJttY/Gi2PqSaPK
xnNu3iSMQ7pGz7CmOIqw2C+i5xFec38FltnUQa/mHQmJvwsz5WjAHLehF4v+EfO7
T3KR/3/eJf84xhhP46kRmo3Vaeuu+4/DPFM0SUHcOs1NoD34zKWlLtHyfEU682Y8
nmRz/wRAuykKoSoEC1BLiOLE5Oqem+rJJtBqR1UQU6rMYHAioSZZLhpfb63CUUHT
UnpWwPhsjpNFw4QgNxH2h3CcMHhrkhnmaXlXFQvWP3Q9k6G2vZ9n3B18DXDpyv6+
r6mlOk7SlgSPXKHhNKfnKfdHpPM/OcCLNn8aO+1BVoHvaQCXH2aR2XuEOC+cicJE
VtaYu1NzpVJIRH70lhfbrz8AgEUG5aT9v+mSynZ+RakheG84PskFF32BdeDDSTKA
Dnb1Zk8LR8ICvuPx4ngDSKTgqpH8u4t0tI0jrzJUzexXMDZuqi5mkVNI4DNCyPl6
galrcW7UHInlTdIF/+i6yvL2YvzjGO9XnHGg0IqnfThywYzx8FnYk42f8leC1HDZ
IEiSWq512ClCXwCyrDTDOIM95Kq6cHpymYv3We7uRpYPSodPgYXIftcZ11qsLJqa
C1u1KILG6D06dFm6emqpq82NVINItLeLcjuVXwpeIrNOgW/L4b7zyEoGnsMbtQDD
jX9Hpo0QM9MffSIyO/sxpw41LPTejAcP1kFKRm3RaT7h7vkiSRibWFwNMeVznL0A
xmvfRP5318FbCP0dtlyU7GHVSfJVEh2Bdhzk7f7L817rEzMKYh3kyn4z+raxplER
dN4ISb304hlXmV2/xbuIvbP/duV1dA4LB/M6Va8+gXWUsWBT9su7kDtNW0h9dBP3
TkAeQdbku7iYWj7HD3/9i4dqDYA9gmNzlK6Jg9Q1arWVIJ15M0+VE93NwNnMA0EY
7IuehtZBj+sHy0XZyEpLF9I5ez8cjHK0Riej6m6ChdGUqT+6ZWxQtCBG3XbBWTv7
cjeJ3AoHZHU06NO59/b4BrnX3cGkORvCN7dxNtkHaxbNeUsANhFbmNa9GOwZa/5c
jgQQHvwKm0nbRwaTyzZlRpFq0lD6rakTB0TmHndaOMm4dCHqk7Wfp5DmTiiSgnLP
8TdIwrcUA1VDZWcrQVyjl0RcW9qCGWIdXFc7qPXUhtKJ5x19voo1N0tLdzWN442h
84E0fMnjwird1w+CuIzKeTBrCJ0ZfWw/+k8eqRrElLDqMIIN1Bs3P4fjvjCuPT7a
uMdN2Amqn2fn9bLEURJn5erlzR64R5csCkUbBTPYIS11DcTO91qZLMBEnZrlHZqW
lOz5lfym8lqoN/1EiYU8mcD1eeYEZdz5KmYLTkXBbvlhnQ115O9uBZFlUtkWVR7q
zHifgtVs4ucqfIusgDowWyAzeXEWAP0AkH1z/CNVb1d+K4JS/59G9qBZnwTShy3L
5IYxSg7NftOaTSGC9sHp08LVDk6YX+oRJBj720q54tONBbaXLvAYqU/neZZb933p
zJb4Px5pBOHCqg3vPAYf8eUsUfgBnSPUUQz4/mP+jYfMw4hM+ZBy409qmldLeE+q
Vvt/rqwIP+zM9rSPX23CuxZsWppB2LxT4Noc5dLwI7/KO32MLmH7WJpQz2FeJFeg
sFtCE1Nw5H7Ipy8rKTJTUXvrrhsP208apyeL0peoJ/Ygs2STEPx9l5bSGosfPae2
LBeT1PwKyNwAfRMpGq2PKSo4zfRaEzJ3DYp2BJo+oy7R6TEUkJykbWvLlwqd13ch
jEPUOx2jpMSbZRXDjJlogB62XjYT+G/4h90A8FLO9bXKPQOt6LVnbPeghXagC0c2
XX+G5raDNNvmrq2OiUpGMvfXvVoJ+HeRNFrY0jF6S1S48FgyvOjeM7S/I3A+937H
DtCQ/yL0obkVoHUGj7VRMhVi6xHP/n177rEY1P/tIRyR2skijHdEe8cZ2W9CmUU1
de7/X5g82xOxlzeccHoYjhn2TGR+RUb8SGSuhiqDzHlpRiexf+XTBTAa8r5bxsCm
M2DfYjWKdey+8l9ammsP491v1iIwJyEulnb4A1zcd60Mrl+hHis70hNf17MSRQHn
uGwSaeWHCOXgia1JgwoWDHXcBehgGCsgV/x6uYBFIFu3tUxNP4fPBCtgczHScCfp
X9fEKPMQMuzbnAU2zNX+ezb0MIrSHWY70JRk0ctoSTF1qZ3JrCiJJMRZyml1Vop6
mZi/3DkDUibIjcoxrHMvz7aHh4AjjvZJEwWPSg31FuW0X3IguOgXkUtjZ5s3G1bz
LbPAq7N7t/EL/i6A4rQr2gVdtTlmOV3nuSQtlClTf2Oy4qXbMMhMVotLZFtoGfdO
LuhOzqvRCsfEvLWBfFH7lFY1wCQzsxAcqyC2Tkozf5iRyQ0gPlcp7ZlUBwb8lUGf
q7n8K/6469Sj8wL12UH/ymWl0asqpEa3iNqWJL2pPg6KhVIqqHhJlAxj9AWW2imi
1VcY2Y1+WRJcrKUANvkWwZgK5QEtU7budcUDXFecDVGDjSZykoVIisymkbXqFPw9
zxG31AIxjpZ36QAGpvEtFr/q9hIHalWRBIdgwV9Kl802oUuyGADVH+YuB4JYJWK+
dGWAxpw8IcoUSE7BbbvM1RYgW1wrDMJ7aDZ/wkMsCFe8YC5VdIY7BB2upew4+1Ns
zeWu/38k5kDWWjT9bNtXDHbi1NK+kXztGoa4Zata8OXB0o02gm86GdzhBqmyj+NC
WEnaoe7ZXKfBu33wI4FI8nD5PDMo6aWm0cN0jsozRrVtz5Kh9YrMyaE++oZe9rEH
gTzCyKDcF2czRwoJgPyJsjXnsl5Bm2B53JM6qqurZ0WhHyJdEZM7q7T/+5GdkqqZ
YSLUZixJJ+CIQ/KHPsuq0j1VvqSOgauWNPnJ0nrp2RppZEPKmIsZiXu+nn2xS8dn
VMhOy8lh8wpEWX+z3jG5CBz4+nL02qzyEJovX1xK44X8Khd25I4u1FM12Py3GpWf
PvcR7Et3V+oe6afUlnqRsLBgKhBQWJ1QjxKKzZjqzyKguxy+nW299g8VkRrBG2kh
U9R6c88ahhRyy/t6XGodtiTTFq1G6HLsoaylv7yZ0W7PP9bjYBBRyhV5cXWxrLzU
YGjN9k9F8UqScc/rcs1f6KZ1OQMHewIVxmarTX6Hq2LIGhzM8VwZfPbkA+FDUbva
MB4eqYxcCh7kukYSlw2USndouW7Zjd6rNt+J303rbKYf5RIShZcq/6OYproq+Gnz
YDlYhjMtJwwfRibMNrEUqrvj6J0B+Omin+RfledDMgZWrhicirLVSBCD3kQDVpvs
M06pRrFV0d3/t8KIoE4xCNI0Wgl0ZHYE/egodC92JbVrfoAZMlJ2K7d6zAxyLfYw
RGdttAbO+RUXuTHI5DYZD81Em2XdqkpSKsmj1FovI88UHUoCkV2bHMLxUZ7ChGAd
GGQ+QU23iXFtbn6Stw1PtgPU3BUoP3YFQeuh7aEAdIj7fyeNQyyIt2D4JH2htU8Y
rOoVKbPgCePIy3EXMEGBwnaC+7gHL1n/cLWwWz2JBqtLAnpokclZWf+GET1TiWh/
qYhSWxmUm1U2yw9Lzqx1py3Cy1V6JE3RE+6Imvpb0el6CIprB6jpDvmjWtRo3Azb
3cZ33tFXGr5TAfYjgpErV6nd+SSdom7aqWX6CaD9gUW65EjIxOvsDLJr8Zy6nEve
0Gy67Clv0BahdICxKMwyW5Ot03+roP6CURoDn6ll+GUvJQBN5JB4GO/LASfU1rOo
4Ctc2e1XRrODIdHPqBbvLOqJ7hof87Kdvm3GosWMtntaiWdysqEoZYs+HXSb8uF3
s33o6zU+Q1F/byt1gZr0Fww5pIxXFjC9dijc9f9Aoif7jKe3IfWSFdHBKpa5Wll/
VmtaTbm+sd1djPMZjObnyil++cyvZURrVxzuYSXieZgciNQO13GCX9BfsU+zWfTK
7QkLI2mltGKCoMWB+PeYcIjaagNeVRjKtc5r5/GZsdAiJlqsaw487hbzLowkd3dX
K44pWN7ZRN1NtDyYMUPV4m+GkfcZWZCEL+53dbTv8PHKRV+CJ/zAWm5gQa23fpnN
x8J8ZkNY+5ll1naeRH/aC2cl9mV062IrZgImxALMPbkIqkHeSTtR3sGLQzfWdREX
uR3sFYjHGrV4MYKeIwdZtZ7rUX826QSeMSHzm0K9fRqbj8U2tsjvvgmXt/uc6Q2+
k/B8F0/T4KkkvR2iGFLWQHqRm1UDkWZw/hILeMDH8Wpt9ChEZsM88Sk1LKrL8uIa
l6M1pi51us3Jkxi8x8q9FPP7sXTPyqBB73ltzPDfg9H26mik7pbC+q8PPy5BnRXM
//VYnaZbjrU+phuEUIz/B3C0GmVPFSmqvDAY7av5fAJUBuOqKRBS00E+7Uf1AyJM
plt2Z+E4ybnYcFkIFWwxpA49rfIwr9rMitF4PxfP3H9ZzofO7cjhsaBdWxGbT/oY
oEfyEMLlFgjicdXz6Xe2aukMGU7IUxfyEhCjkglLxoanDNIffm8uFtn3UfwZtJ8u
MPBYA28t6+HbjGQshXWmjqspQomLIBspvEgD8BydxBFxuyE0fYOYTPZFUTUhrH1s
oANv+rvc6gM4ce1kVVgq5eN9XFotvpnHC3okRfFOcncOrbX0jjTwvEC0rmPc8K7Y
Zmc/Rx0dhlmu8lN8qJwZZRvUumG4gJtx+wRu/b/Ga2AMnQUSG7tNBkMecxrkItVE
dovB2hoeg9GOTOCClJRRHfurGZlRkAfrJ2DeARc8/pl5zzZBrfo6fCEhD93AyiAc
p/e1e/kD4jx3u8VI9mMXh1yLE1tOB1grdmnuptnFmMHq+X0WR+dxXe+btMOs3y4S
ZZ/EbLtAUBij+5OXV+WqL8JaRDGRx9wf43/8aM83uE/GDwS8Job1+s9O2+Bh9N7H
02+WTGznVY/Ejq0pwMFDWYfzUeS4MWHEfUXnxIBB8+ELwHLg5xymys98p8O2AQuR
FBn1R4osqzuAt1ouZllO9zh4RPpKBoGmUd3BK0tbCqRLeq7g2VD40c92nZecmti1
hsSYaF43sji2dvzk/j5/gFut270Rku/n8wo6TuLX246859bTOo1vgkumdxk0EpXz
OD8PM+I8AOYpOwJDRPDiyTq5rF1ZrmG6HOD5zgBJIyipqvXimTALU4wPEln1nkXy
2DVZpoTbYA2hJMn6cXxqZNnyvsYpuwS8IhRaFPBkLncIIoaKAE9ReouxdJZgIGmd
evEG5pkZ61eiqzWrKBvRlqKH/Txf//CCCkqANRm6YesjZSaYt57W3F+GD1i3lnuK
cJgyNBIybRqNJ/y3V9eEk9wp+VV3i/+ohTmaVhtqS3bma1/K2W/xHkvxv3uokY1t
doIp8EpSgtS+Ylwhmk+FAhl8F30PJ88UBtphGucaq+fafjkJb6LPB8Hl58nYxej1
77cyxqYE66MOKVmx738q0EAYKu++2IK2t0NkGAJAGlGQKPOeC8Ui1oR3w58DOjxe
Uiw4//U7VoXFlbL8s2leiMu98B2lCe+0IG8by4U7gShLQLQfhKxxY0pIfFJC48t+
NROte43yJKdnbjs8eZbONiJDPo/lAw53/hjaqrS1khYGJWBWPTpIRub/fwkC7OTu
ek1wil3CjFfhenqG4OfJNYCaYN69rfHDpFHbCvV+pb7Jy0AkgBc67CECLrF6DsWv
BGLfxyD6JL/ZuLz8yPSmn9TyzGAnlN8izI4ZiDZU7KchMbTlIu/T3Y9f/oFgF9Uf
DQf7yI+Q8qGzZuIz+ckmzxeae7eMOjDGatsyayE05617/jf1GkKJBFwSGDzoaBNy
bTRH/2pQ8vYB16pwcKpBGHtUuUJQ9C09eoi4wytc5NToHZJiRjfG7DVgswV9U8kD
+Fq+kVxhTQngVqtEAOpi6/qkCFj6d2iRLQ7fVBNa9/IgadSgt4sW1lZ79PH7QkhV
baadkUdx9DLIIcFsbs/2Py46SNPPfwPoOLTg52LMKuAu5YdxHUyfrT2i9pjWNtQQ
0DYTUfIyc9n1POX+ebF3FyeRi45+Qtk7UpwnN4gWBotDfU5FjOoK7Xx1WmSMHqxA
ePzasrDJaaZoEpjvYmUHEM9RDuABzean4lCKV5AZYXAzKhI02tqPZhj1KB9mDWWO
DNcHS0rg42tDdN8bwA7vW9SG5zur3Hh5f167Oa/CtmsVzXgzhNE9B1uOim1PlbiG
vxKWWDMvGkRRnHgUnbPwrqLEYh63n9bOECK9jaGcBy6a+2MPSisejP+tszcCXtcb
bOwPooQxx1VMXP8+lmQd5YMV42KSy5g+STXPwf05IBMy9qH+XC/k30ayh0bm7yAq
Q7zDgZv+KatqqJa1pRMn7gBoFp2/sVN01Y3AFo5w3yvmtiN7eokp8DFQFQ1MUk/A
hKEaH3V03TlTLDH+Jf2pxdqk999RhDr2pw6rT6Dde7rEqw+O6S4Hq+2pCC/Hre3w
N7ckka5A0NNwL/cIYtM0O2gKh2+nmyLyGmaFSLyGu6DHCfDBnpobLkKLuQczl1DY
Uffxzof9JoxeBnehk70b3KGtP6gCA606Eqe5fpu6yTNLuvGwJbW6vMY/y/KgU/tV
RM24ICtPF8RzLo7SNeOOWYBcNlpWalArD6I4QKLyy5JjA/oA9hIHStMvbtopWvzm
BepQdiOPPTKY+//bU+id4vI3Al5OtKQbkFuaVFknmKtUj6a7O3K+cWrVXj0dijNH
LfHuxjvhaKb28FZXCk3PtDayLOMd2OC+NJ8sZTN9FWW2zGErjbfkJ7ElAD7tjBmh
Oj5JwZlB8FsQ7jG61yxB+jpCRzlNPYytDaMIeUwY44rb1ZlzORqmHnvGa+g0tb3w
bHkEAlef080T+pVK0+DT148+J3bHhQ/9dwfQZcLmgg9MyiJnkVj9rc22/H2U0aDX
M6jPeFzDkBWbRH9SNUkQKBU7SSX1i6GucX8TZXE7QJk9mpvarLSthIQ1FqMD37rE
mYymTtecMK0ZoEBoQX5MKsNv2Oc9xRc/t6ZzSfhsEEgahw7bGTUdI9LbZ7Ccf6J9
QSDFy71BiSiFkB23oNPibs4iLbATLS9PT2NC2pX+Pue3DYEqqdTGF4sRqJxjypWQ
0n9dMs95BMc1dsNgcwybZFnGDtWu65m+GRjwIGzbVydlyKm+8PYycTlTiQNtofwZ
ISMKrXI5K0sulwQI+6c6AmPJL2sKuYe3+oraXPwWfsWc47/5tpcIeQG7SZmQBSgh
b9GQ/a2XVond0JjlpnDJ9h2VUYGDIdX2HRCAE82a2a/Mmr8iasCdPReBu2p7vDRO
L7rajAZo11ekUHk/244B7Lz7OeCJDOfenDLbpwP723oNk5AdsW+Lg3RYtMGcmiBh
X526yH+d+LAHUEX5lPHdlRqTEWlBhj1ilzpgSUnVvBdQpXAeb8GkOJFvxq8lvyyO
pjkh+RQufxCn49oCASeC5kExZZTfx7fCsSnRZ2nA0CtSBPkskLkeSO2KP5h+kpzL
INP/UtkBSoZxYoMZepw7Be5Qoy+a26S/92sWR48CkV1zY/gyygtL+RFe13j9TOAG
uGY7EuZEa12y21GStBLLeSXIMfX2ss9CwvyFsXfeJAuhNBhjKqb35NnmH1QOfCvY
Ps3a8eBWsmuvfMjn7KUAfoNM5RGyjNNB6mhqhPE7JSvGnvZkfAt9n32BIYUJKbeq
QbTefWd+Ogbr40o85nTttwoHsy2WayZ/zMYDjcGMFE7pLD7lygC8iNQffYPOKuJg
LNkTpctJ8QAmUwFAa5/2lri/d6ZSwbceKfjlpi3oDcO+MqJZ2XG24kbrk0BNRPrL
MeqB5FE98ii72AskSZodgyv8S4TqRE5iedEG25VOGSb9UAM9Pgps11SaE9XHb+8N
8RGyQYBchq432iJ7f/bnw27WnEPi6TNvxnsefuT5t96SzKZ3TCxg76lExN1An5qr
HYpCCegzGCtIjROgYWkuoWYKUIOJoVwe4MrkRfXPcIjdFcWv5hzwZ1CQzQhU6oW6
JZI+tYXgjAnqa9XlR/f1W3nk4SBWvMBiO+qEVhRmh9LMur8e7wYn/shFRkY8sk+M
Jz3MOCNAJb87luMS7CY2BlxwR0rO3/s0HZcvCjNlo90zxVTmrC4TiqUVyo647U+u
A5AOaSYWF2W7LDgyuPxdLWJ8xjVTh19xe8LqI4o64iOGqdsLJASSkUbtSjr2084w
UEanaGkaSZvRLjZ1iR/tbp/rKvKHDkAbcecZUHFdgnYTWMOsuag1RVQKpEG6PDVO
Dv8fvGRJ+DnIFYgWHgNfTzAB3ynAO1Zngj0hpXw/GajpRGUK0q0h4Dyck8v8I/XU
vJ6ySZxQWN9qJ7oFjW2qiXdKWHSbkbDn7KVNUshr4zfOy6NZWn488SVuqcz02K11
P9auvZOLf695QZbcQLnbFjymaQdfr3ax9owx6vkqYEzVh+oDJT+j93FRWZwjiyTI
r1ePaRyBptY0he3NQkvVaQuhU+OhVGXcZfE3kjjXsgQzi5x1IIS+C9zuLozkaqxC
AHZK5IgQ3FIiKOT5vCeLLT3IDmfOcKKQmF+fS96RdItU2x617gU8WkcsVazGRa3B
9TcFKDU1qJk54iwhO3a5i8RMO0N6imQtl9gt5A9HxbqoMKLphrwYXNB5muckbkBK
t7L+B7LoF26CVLaM/eKoIeEIseUfanA/9aYyKqYkR9P7h2PzbG9d6bhRSPXHx8wV
A8WT8z225DqWWAplJZeEiTQwXjWybRbCsdmLrnTA8NzWgxm9bqKcnv5O/xy5Rvkk
2oefK0NWIj7fKMstZkaCuAfzv2hMUlcTbgRtMkwEInBuIGhzlhFs8+AiM1Iml0rZ
wTCgvAk6zPnufSdeaRcDh6YspcehcS/i/kyQDn1PB1GAEMPxlaTr84685HdXGrUa
yRH+5vk4Z3Zq97TkFfsWq/wimGca3cB/APvjEulNIN3k+KwUSWUKEg2lDA8lvQ5k
Us0ij3BOWMb47NYzCM7HvNwFB9JlQj5xMypxor6ZZTGcXytwz88t/Sf/Ql34iLVU
9pPCDithYRUwayXl+jiqRsZe+hLnXIQmRTRLRDnXPvncfnrnI5qcdACdWxZVE/rC
ADAwNl5WtvlJpqVBO+A22Pk4zjQeOaYlq7IqSP3VjDKlAmq9VZ7KUCdGBb1zk4Uh
OZgMr91eaXfwWu/w9emjRkgeRNi+BMXHDxBVaw5Mvd2o2jks0UYDoQmDEDLD41iX
yRIDaPsto2qmb1MbZrRPNc1yw159zrSpMCevOtBx8/vamUR63EMCIlD2ugCh0Eeu
5G6pHsDVL7WvZzz6WdaCpcpCCfwrfvPpiiCvD1CG06MTGzOJVSEMhLcrsn7xZaPo
pkj4D6UaUx9GBSgsotKMhzvVZBx0hbBBFEOHMO1w+XtbZA/vvGxERxX8s5ImlmA3
tW0hBBP5xggU6P2Ak/jrIH729ALt+Y3NAnQ7Xtys+xac4mIPdp9IS9dnHWc1ZcDj
efLxqovzdYA8rhnDqGMRav1lSdwzRysP9wY+R1gOfvNs4eGwJDuJPb1ksf9Sq7WC
NomKhrx1T8rCufPj2UTek6kPZSuTBpTWLsFq7FLjtrpVQDF7KSxw/BTlcnUu1Tgy
7Xo+GUSD2RaO7mH5pULufn7wlfA6i73Zt9AYpuX0yau4rZMU7Ldyld3edXzP76/U
MLdLSchUngEVv32xdqrgm2EyySRqbL4MPaXPmlP57YeXwZkhmc25ntbkqd7zkMoQ
qQlzE9h49FfCepAi6mKASc09cFTNv9Fhi3ielWuXll3OftE5fic784hrp7RF3rAW
tqK4cMPAX2VRHE7H9RnaTbYCZ3bM6kK1aFFAoAa7pYTQJOWAGj4sJQP7qyMbJHEX
APcQoUHGHk8DVtE0OoVY7VCO2/rIFiv+Ls8DHG2tbNUTYI2jhS2Yt3RLAtv77C7Q
vJV6KgcvHhOZiCXnJxj3f+JJurYq1rpTGTOPP+MPoxnCATR3Kk6Sos5O6dqaF/ZY
B8M5t4rmRPX22neIDULLf3eBs8gSmtCkc58u17cjJM778flvkumQZ6Uj6v3qEDvn
1YK7RZnomVMksgJXpq+i6grcpvsMXxL9CmhE2ElQV5KNlk4ihgR6SDtGU/vzcRhS
lQ8utTA3vMacFf/cw8BQUpsxeiu7D9W47zm820GPpYNMmolxl1vE9bMV25X1I6Jc
buHPW/rabh6a0TwY1/VHwRgaYYPwyPQ7sGoqypdnnVXB7oFdK3EauMpPNw+H2cxL
AX2U82HKcZY9MydgIY14xrI5a6FHdzeuLGaLQJktfMiy/AKTExD24v55z7CblnqS
7CUUwTEfJxLxO0pMZr4Ap69YyhT0xXvARIOO7nQS47C/KhHDaGUBiPArq9GYNV9e
Gp4QxRqbFO1znFFVdaOE+iCLQyOpjeUjU7wlEjhiIlxg4dQVe34GsDROrAokXI3Q
uBx6j3Sidh8iEzAs6KY9HIJwc6hJ8MVIZFZz0Yw16naJvs0QIGslwreFxwhdMUE+
JA4XSjEo3zmKU9VyLVjItdhiR4Goe0qaoLiNKhH3T7fqX6aLQIgRv3y2BnsOAiq3
hfqTlatp73dui/F1981JX9/aWWpMM0CUiCdHsDRbIgLBadJxK4s9wLSDHgTJdzUq
+44pXX4ays79MmPx11Odcel3lZc5bjHzUv8Zb5j0Ctx8VgdEv1B3JMgIgiZi+NcP
RnVmozg9dL7l8UCztq/a6q517pjxhoIkUQCHzKMJ1TxB5EGUJVcd1SIujz+ff1P6
xB47Xq6g1/qE22sGYYQA0q/o4xhMNMGi5mga9Qw9IwxVoLzVS+YxhUQpb0OZOw7h
EAPqAcesWCyobUFapCdG+P5QyyzbnMHIdESRBF1Fq2cxQDi2zkmVcGi68epGzNww
b9a1GBLncLgs6IAAlwkX3yFxMrP6cGdXMTLbbW+GczemAd5R2jIT7NVse14hjweN
F7ofOA12GF1az09fIlGYfSVkD0T+Gcbqq2LnWOSjS4Jjp5GKRKn7IbmWcflrU062
wLLpuA+7DykVUVCPKpiqlN+bkynVEhmSxVngLwsbOx6mApp4aFMdo/vKzy1UwfGc
Vgl/18hjxNYD84uHrYYK6kO6TknacgLBKyrmCWFWL/JWg5ta9KRw7rA6O8t3NTUn
5olIFKCrLyZRUs0wyk95cJIzL6des6EvBzvMPRQN3V/e6DcOeSCIGfQpotU6KmJD
ZLHdsplQzrUO80RA+wIOYVwuPC/watN630gRRh9F5MkOjuLFNdMMWHE06yiJcFL/
9RBcgNuj5+2UsWoBWHbkDbmIBcp3QMfSWSBg6YrnwIij1Q8BYAC42CKnhAjQKZDz
PtyyJXhiveYATnhdsREDIXUvU99eoT+4+U7RhUVAPTV8WvgYLILqGdKPJDV4Godh
IsXZh6aR6SdM7jdgKGrGhD48uWIBt9zFHo9rY4BQKEj3aAC+Om1PFyfylJOjn8kR
U0+06sqyOQeqQqwIchTN+soCNCeOD0yZMK4bBG5RIcn4xwLjfX9IbULJvWQ/Wf9q
gfTOKOsMOx3sfpaN/S7HhexMITDFEf8g+WHLB7MlU3lyopHCqsNdiZCRy+NiF7Av
FwTYF7rKFTTTrILysVwP1w3Vxj+6saroF3xpu7GOUiaRLMjqbepU035k3lZ4rd6n
nZD0JqkGaXWQbK01LL53EYD9ouDxcB4IroqrzqoogncoQYhLJi+xTKqCAyxmMv2N
nKW4TNCwh3mqApwR7hta+BJ1VfqhsWleCrj8MIljI5PGdjWtMo8TKc9GPxChw3MY
+nZCJbfYZoZYTvlJYKUH54k7fllBGKRkz7nRXSftUd+cn0nyMtXsHmoex4wrR3ks
IgtS2NZkWEA8brZBM1pKFE/WLafaFf49WLrRbAqPUTQJW8CE7oSsFJSKttiGs+Nv
hTrGu/koeDG5R2QwiR+3hXH4UqcupvCjXzK3zvOpb0DHy3VKZO0raVPtmbC8W7K0
xrG7y2QQ9juUi6ve95Ii8K6eVCACr5TrF30uWiDso8/5qXwQ2ojUktmKbAiSh+/C
ENrIclRVJLbjgcjMgZgCVov9InxkNHjG80gNWZJNNcpZYtDa0iEWpW7Il/WIBguv
+RgJX8J0Fxx6tR6jOgirC5H8UXL08q8NlpLzMvJPuex6NG4AaZ0uVNmdd1wtmXk3
rzv3BfVt9mUZiHddEAwKn4FMkUttpvyZQmxj3D6hv7klaTsuJDalvzUhMe1qS5e3
4JTG+ujajX27gkfvNRxE13uB14UhskQ3wErGXJB8jXLic7SA30fNM+yBptB8Ji+P
uZNS7x52Y8ex7yAT+4852c9dBHGwMKk+cqBNzINGsUckNaksJUhNtYTuGtIA/Ait
mnWtU8pRsc4t8una/vrLL4XFvpH5jddnbd3JJbUv9GYIBRGO2U0VbROIOtpPPQEA
y6Wbw30jqm5OClQJLkQQMl6Eu2XKjhJoWsEMIj5Jur7zZ/71g1NS5Dil/gPDCics
2pHjd+dJSnM/sQr9lLusnlbap/oiA81hP1HSd9axXpujsoABXhv6clu1UBynIfp7
3ci9GLxaZkG88DH5fG76yIjE3dW1rxdP5jcxLRnCcO6gp8lXr2tKGMoPRH+caB6c
uhwmpAEa10Rbm+cHd0QQAJLcy4F9RLSCrxhXJFenlRqoSTAj4LI+l26YYfY8T5o2
kw5C5DbMjYlWJCdQJI1gx4pueIyDhfn6cMjd5XRAdSp49kOiEUsXAqCinUlC+gie
BG0SmdPzxVujkBf5cmc7SoYUvD2J9hWSFkQ4vNaiL9AMyD5UE+2k4D8GQkEjUxiU
QIUt/LA66ENjlDXORfcICx9oNv3vizNF6YeEEaHC+o7dxD8ehSsxTVjiflTKanM5
3L6l08roe3l9s9OhqJ6LVLsX/XegMYvwq5MxYU4pdrzN9mr14lBcjii2yU0sT4Sx
LgX/Pi1d7QCEjPov56FYGmlKkpA53lBixBn0nvE0eXKAspuPF9orX5D8InVzrEo4
pgiOc2z0EWZpl6FNUqkFVZp9yLfTCLB5OkCsVOI6pmXpx6pIAzOP55KXgFGxxlcN
WqVPIetQNpDxR+hHiJqC3xXWri77sPRe237EvSArgfMG5jTZetqtR6hv1yWTotqy
xh++uSl9vK6IjLeDcD38nnawXWC1Dr42+DRusSqvetmb5bFPqP63evCXtmRM4lVx
1ieXGO7Y3FFjoGNfLhFwAv24dbfTCPCGZjXJbJ+zO+kt3LZMnM72CxnJNBI5Pvwo
VdKNMQfX5TeWlKkBvch7z5rgnqq0/scwb8IFsLtun8qLB8aZYOfCFdP6FGJrO5xT
vT0/HR2mrKkZHt9gxLk23rHxfIHBaJaYYQtGm1t1RO7QCfNUFlqBNzRfpO0ALQKh
JYA7Dq/e9YruaOhO1eb88+kLmAM8vLBVFxq0/JdpkWrAvAGHTxe4NsOVOGaLD+2O
QvPXYuT+NTfBdz7WH74WE5e2wrgOLGYXkLV2sQKDy/MW3+gfcM7/m5WctEmDMeqh
Cmg+xOOlJ4TCyFMIP396s5RJobTop2BrvjTu3o7+bCB2r4KEVE3sT5MyzQfFal+O
9aFKaIk4kb/X23RqAP7YSf/PP/mwR342ItLMVNu/uRVN4Aac/OYb6VWMeHEWi4MX
QEHufpE9etZhN2jrZ+KuNPYgvn0NH4a6ZYl7xEZuJl37Px/XM8fjkiFvTHp8b1Hi
08xSRfsPSpOXuPR1b5q0TTq2/M4OwkTvFDmRrFi0iUBiHrK/YhFC96ps609eLP6V
zFrdhAJ/FKVKRcgTv4Rcb/IiK2DdQebLXcb43/wQBqa3NCCLxtXYiTm+tg2faxH2
gV2KgjYfpiX2DBsQar3ti44XfZ7SdhFzaOyvBKtyXfP/tuZOjA4BZ8w86aj5o3S6
0YkckQX/lvng616IiiXAe88IyN+m1NLovuyQTxeZpuuOGvU/Agd7Hco/kVEyNmbC
P26+RTdnOZeoOrf4vYRqcqSg5YKz0vwwBDMZkI8PfHiYBXfAMOCXH1Qb1I96RgMz
UZbRPY1JNjWA4rhLnWdN5zaYjd9H0dKGBOMAOWjrDQ0ER7N5bT3qMN9dZveIB/xO
feC8sJ00MnYuK8reOAPTvlzDzeRvoDL7eSeAmgYfUSVnymRNSmiAKkMrPD1eSOMp
1IR0zS210RaednyDnnhS0r7GNvLKw64GGe7O135cw1b0wSDaHU929OUmUmHvuFfW
9olC0L97PkMTo86F65rzx/U90LF51ZWVenc+eUVghCL+1pNLR38xSsfrS+CqKcnS
9d77NM6kzbC5HHNDknS63BAOFgHx3P7OLFzTAQZALmXM4/7RCZvO0Wq2MUDWQ0kb
bP2WjJURWzRweskcaaWAS8aQw5M3cJzq4wn6q44sBTAzoZpWYzUzzCnbv2Iwxc6g
aF8GK8nQa+7i9Reh6gY2Rl0VXvu5atf28T0z+5ITXkZd7WBs5RSPwBCPUNUaftPl
kbrwQ1d/MXvjVNo5WHaBgTD0L+otTJuTZZYMlioVsG5aN7rVhrgSdt97W6chkeqz
Lx/HXn5kQaXE/3w807YYi2MeNmbJdSNOZZaCXHvvsR/5hX+nkzdaqy2io//nYojn
peJFYHdPecJtvuMPjCinmlMccXQYyW7LOtYYInkSt4adBnERnerYnoOZpvnwTmRF
U2ZkPxKXQmMXld7mBhMJNL3YUfc0/WoRA/ZdT6FXtjFVlyUJHse4xYmGw1Op5Dup
ekdnmG/QpfkoDMJdHcfMnbI5WaK54IX/HpjEGoSvv1xrdEeuKNQiagXQk93H8yxZ
59gLNtGIx0JXG2E26QH6VH1mHFQtWKEkgkyYDfG5rsPw5Zm8TcfpO2XOLvQ6ZlOD
BjhoKoN4mYCKOqascsIYV6k/m99IMw5s1Un5ScCoRcPPD0Yr8N06HDtIw+1AwZxa
o7K8FNGKkdUq50xkK65NLka+HrTxTj1XBukYWks/5+M/6xjED1p4I6Pfvr+HKIUj
N/NIZ39AqpNXa47iqPQtY9vrR7u0e5VSKlVu2wHWORCPG5OhNRkt4ZGHz8QK0/0n
Dtj5+wdo2WvNaJSivNwljW5iYpWqcDkLT96EAMFqdQhPnWuH6RKlUZGeUOFCFzDn
VYlfI8sTLEcVS9LWV9VnTVGBGnfuDjSppWQ2tdZ1bAIhaj7L2OzazhYZUCIt07H3
vGaZOj4ZgVllmKE6WTWYX+jguxUxO/XDJ6RPef9ofed61rNHMTdoSwfm+3MJVj+N
nkHT0jyKNlqxMKJfCVgsBYGOo+zAFTamPh2eBiB03ZpFzD2Q26k5kzRf1zSa+7a8
ljhO8uGDIkaol1vlESm+EK7Xl/TDqU6dMua9jGFZuE8IbhXwFFLOPjhEoD5Fz9sB
qILViOdE8NNCSYK5IqmHME9Xu8NewP2RRdwO8AXdycZZqJzGGBcH+eofHdyHQy6V
pLB6u/dnskhR6w+j46OUa8eVDlmoP/O/m2aB9aUgxCC71iW+HD6mPxL8nCUl3+Fy
C/Z0luUfoNCh/N27zbDHfzZJNLdawYOib5wHUIYd5eSSlmWDdiSRSPjFmCCFiATg
eXWxmpEtftLqqOROGGNKBrcthVqYbZlbO+6mCTN1DM3tTxWYphwMWtQ2Eph4Vi58
jrfb7CTGfIYYUBTFuY87nTRAey1LjesdACNl8kKefckLdDIBS2Cf9b6dZwmz7T1m
4/xNOWsUedsdF88Da0i0LNoSZdBM0Ta3WfHJSJ+SSTgmXShBAS2ik8YQKzwMw0EI
tcNwqbk0vFEWzVDiX0LoVxivnf6PpNI6ExQ+A9EUdBgIA30XsQmudHWltP5J09Vr
2byEwpDTteojA7JexVeoDWvs01GVhUZzO/Q6P62djuasFz2Zh6hzs+E7Ys8SucLN
b/mh6YlB1BGdqVdO0GOO47fGM4FH96WyipfkrZdfEJgwV/A39UjRLtMa5Y1PhG5y
ZSaQy5l7B6Y9vHJOP9a8e6xGYBrwcmlg59PTCblQecs//2pFn2zJ2gVEyd91AaRO
So+FDLMxTlkifYWaDoB5497njEoUgEd5VeJzFjM2E9I75PIrnfVaU6xA/KE6ba5g
IAoc/N3Rzdr3aVC26pQbMbGVRFrenq0MbMMdPn+dImjXVlvTRGQbQrbJ6UQPocGk
HzX3LLysEd0fXvchombrVxESddfmBEQvCWlc4onbAGHHItAeEq7HXGNIfSi72eGh
rk1rh6kBZsGcps4B6U4F3QRdU+Bub3+2Q+6YXLpYVAlRZOH0FjSriwT/l6+9Cfcy
LMCKGBQzTrhNvdZnHTCi2I2sa77eEmAIXj5rI/ernpnuMFqO6oVVDZ4KZamF2yUJ
DD+zHxmCR+rPPhkJdIKjdCiwYtdrmgm1i9YRASGQanA+a3F9EPtrXQVWMFi5xbJH
DM0btUzbdjWuJtMk6cV2mnZdMKM+sraxVXlUYwJZj9/9KER1gbaalY+GIB9ETOSt
KY0sfEHJky24vzsQRUrf4pqU81gK5uOtcwlRVbtWm+PdRBI0bK1CnSeHYVlnDob9
P0rGXkBiJxkuHaN1hyOMIBXQ3fw70oOGJ9+8MaPpicxZM2kliyMr4PSggtL6Mefy
YIpnFG+bbFDvXA2j/K1B4OEDFngzW55/SYmA0I/0XnHZkqQGeyz7As9XdA80Vfhu
8TOqQ99SS+2MJVt+24N5UoOmwHlhHh/bwdNm26ehGDsAiyWkihcWbq6nf4DlSFEP
IdA3UnRtnWDyYZuUpaaoHgZ0P3gKS4t0LLqTjSqFrJeDcMA+Y/jQKRlQutQW1rVN
GSivnkh9WMZYNbRIxxSpfowt56mhKdJk9Or1UerqOQGID7hvVPH8b3A1VzCN3869
F44vOhSotQN6NC+G/Yi6WbwPP9taaexJ6XxNZRbUXviG5lDH6giDdNH/lFWyd2EL
Nit7zhax42aiy5WVjPJhzDiH4jaZnktyjeRg5g+H9EalMQRrHen/+5mu3obGh39/
UEL7twJfRP2KTg7shNKQ3kqfXNWgYZb7uc1VTAC0j2fcAcLwCD3DXABmdQK3XmIv
q4rmF0mCIXmB+ThCee5n2fAc6bA3LL5+N/j+4J2zycxBK4xVPLvT0GfyCsUjLg5z
rxVfaA4FQ04qReoVw9by6V1BR1EDod4OLm/SwwxFzt+N4yppU3dGPB4qw5hmAj9Y
bywmwa6xzauFzzJScXcRC6GvkDsPRGbsbCOOh/LCgNV+K020oUlwqd/k4ja6tmD7
TIKiAyYScklW4SOSii0+Zdkylqeaq8470p1Hv1O1x6/WExa5tFXQLt9UTPnnUmpo
xEQyT72tTXIsFeuBK7a/D0+wFZuqCRXXxDL6FgG+SMCAjBJeVizQTsq76QRnAScC
LOd7qziTXuif96SXyrAw82swbrkGszIKcH6m2wUsmCfIU1HwmcWl0YqqecG20Eme
QWO1l6RRh+2N/VY1lVEGORaXe6ElSNAWFHzeVhA8jEBFP02FlxAnci4CpFaRqUXQ
t9wC5Aqch2W+zA5/dqRooVFiSlVMuygmVoEAdpLdBwbNm+aJAH6skzAI57X5SGke
pmGikQEKtzEInCS7+v9WAmYIhE8AQVjjfE3fghgXyvkIZifp9aXvA+nqRWWALmRB
rfj1Hq9eN0RrD4Ot8DhejraEvczEUWEghO/rjweuG4hnD+CS3+orkpqGlvHvAXhl
9BH03t9lnjRAa62mdsSMN1YtKcUmxsTWg5Kd4/DO6hPnFGPsOAq9PnirpN5y8xjc
9Wn0Y5USr1rmIbCP/9N21hQcCkLDQquRVcdU2IarqpZ7diG8vV/n6LemqMz7bRbk
SBdGv4n08+/zv9+h468miqE/194dxiLT9bVGFVLLjSZuOoy67yWEWYkYLhkz5w9t
t2gVynUA7aeN1ck7UO2bwfSjVAH5ayialKelLJSepLSa/8zTFOkr6PZAhbsvtpK+
Aa3ugbpxJGD1qn2nzKrYHWmmEc8IuDqhckRlKSjlMhbIer0dC8Lr5RQivOJTnwPx
h3zNnCrYFOLHqhHaI1bUVLESsLcoW7t+LtrAi6+P+hWImXOKkDvT/K1jNSW83Beh
QoeJH3fzUsX3E66my0nRMEAP8vGGj8ZL5htAw+0L/JfdNvkd6AxWC+T/kUDUL27G
2edn6SmSgvkCZii1IWb3B4YeNoJiIPa2jyTQbYarjHzpF6la+Tb1b9sWuwN0hKe4
GvoIArwHOb86AzV77P03tw/oMDJCa+yDYsiCVxb8+jIrH2Wag3dZiBRCdit9mlbh
C9TIi7ZGX0lOc+pJhZjO3t3Rg7tpOSXozIc7FO0wBD07rcOOzP1omEJRt0cKiJVm
dMXhLws4IdIUpwc7kUZRVzy82cT6521nVFqLAh7WWZaRZAjDTSJrbQplijo+jZ9W
cu7A7BGxjWwcyOxB08yOdsN01OWpDLp6rbOSSQwiMQdEGhwd/UqgNiADqCKD+U9J
I2Fwc4FRXq/0P4HG/ITyNnmEagI9FhRWKVDfR2rSfWmED9mxjBPs96kyitTIMJkn
Dzyi0snzq/bHzgyWZ3Qka2gsOIusKC4UvDV3yrK1gWvJpyWr84dwm2GeNc1K/tgz
Gnv5pJY3OD/NCyblYjBS27X8mkJqKxFx7Xn1747MHEZ5/AB9ky2L7W78V9thl0so
mrjGTgr14Z/uvIHB48eizeG3jC2FvavykxmDG2KY6i8UTPi96ZPHGK20LqMHOYN8
7SheXWr5d010tkA+f5BkyokCBgW2w8SmGtdHIg7/jEr08mHRZTKcOd/R5cCsUutg
rLez8aQzlJ3JhK6dMNX8AmZcAAULpP5eVmEN1qGsq/UT/mlql0zYiQWTiIoJ/3KP
HRf8qSSMBqRtYhtCSLNem6OxhhOjheiH7WeATDJkiYDnrrj6NA/dp1BuBzeVSndw
LHN0HX0Cnn66ZlT8VNmtuyolLNotYaWSyH7iMWL7KgUaAaDPK6j8OvWVljqptjSF
BKj/xXZJhBJUUXKue6YiMQ8kZx1NUL9EDZ/S/VnmYKPHLhgdkllfQqeyefxgOx6o
4/l9n3Z7ojb14npfdDIf5J/YYkyF0kaNidOTKcwGKTEbUDQZ7EZFwn9X4rwUrwG+
/PvBfoCEhxdt16biPfAN97bE9jVNm2imvP1smQdR5NxRs1++Z/IGMH2BxQiwcPkB
NXR+hDbVabeHOFVcPMUkVo+xDSXSZnGWCn19o4BSIFJZ7+WPvEEAf0Jb/I3ftGtI
vNA/lZjB/2pUTymT+28OQrz3JJZPuxoc8RDj6mRO9Zz5f4ydlHXV8NlxnoX8DgaB
a58oKMxt3C3jnX4RyJiYoG0otAp38LioWFERckOtSxbSttIH2IF44WK02OqBhdYT
ht89heG/ZVu4NVl5KvPRXHPsj27APIMExgIUxgCNWTmDm7uj9TK2CZXRBDanIbSa
d2GfBj0TgZGqwqJ79hHznxaoyRGa+k+q7Qdw4yu7lXNL7yC1vOuEPKudLVqPUK5L
auF9tL1A8WVjgqLBZbeZAtrGV1CLwHCYiIu9t2f1YlFNdYuTX3Dcqpf40yH8qf2m
A4gf5u+wVuscmtJL9WZi68ESjJImylDPqgeBgWfUO6OeJfvFmDgt3+MeD8kpvU7g
Hf7za6d97PJIiDouy+1qCDRsRwBJMv5E2+DyqZoLV8K4e5asXNxvTT4ce/j/Igto
Q49fy5HSupwnLH6/7/KbmQW3P/6pMAijoHqm4Plnit720rkohCaquAuQbBk9d2VF
NiuAXZr6CZMCMdoY09VeABehBGDy5NHJdw5eC100HU4Rq06qtKHwp/EcFSjlN/8/
A3/+Ud4upmwWXV7BBKb0niG/8XMwO0RO0pPqTw+FMBSs/kUZ4deRKbS0NuIv7Xzq
KHyExLg67Ui852DiVu76Rv8Jd1Ijkj0Z0/y9nza6oq+P2/77S/N4Vuux8FmJgwfP
bM0KBfJvAZkAfDhzd27PY+xtaVvNhFawwHN1Y8znaYNMcj4KqJpBdqU6ODZKUj4W
3Cmccpa1XJmt7dUwCGHJQUP6y6U8JxNBT3NW1GUO6JPSp+Rkt8fJSa5OEgb+zgrR
6+079xWrvna7Ec5Ev5NUB+ihcIsn8S9Kp6/fR710SEMvibqmkiH41iTW1uZsYcqR
MzF75UUK0ogVVR9oI42OJjUTrO23YIjsGqf1/lDMaksJreqFynWUBYMvR4ckthAm
8TYaxgWFL3WLpJeQ9hzi3qzmTiivniU0yTg8pJq4JEFP+yspR/W6/2A/acQmW2gO
SObj7b5ZhlzkTaiUmBogClAR85bZxgAxu9nw4diwd5BxBFVqN+rOUiRqtzgWSm6w
/pKKxhBPVeCvW6a079sDy+OFGrn5GrMeo4ZtEVRL6ODrbDQJGb8UFgVr1NL1M4xv
bVxoc1xu/u2IiqncgHJ+jZQfdjIYAud4tL2Mvl+V6Vg5sg4EV5XGPBb9iQys20bo
d5Ebw8urGSxZI8hmSPwddEDzW2XH1Ndyae+q6Ua8ewAlEmgZXDtjaSIp9R6HCOg8
2pkGea1dDqJYTPHinmO0FqkZMaa7d3xV5z2AhH/4ETlF5u81pQFSICaoo4FFSiLq
+h9IP3Mlec0lpUbAnQ6sSNw4UxKwbMswaQFgL4lsftJ2qB/WPJjh3xzpLbbI3Ewo
9pDVP6BuKF+ALzOzMr/oY/EQIe3K7qA7neXnOBbVOL1peR/L1VHE2/YGovlcVLIa
1TcJPqyRO6+jge/RsxPFSUYku9pN+3FlV36cm+ncDC4w1iuI+QwBgHlRhPIOr58x
S4GdY+qDdiVxPWs79lWIRDdkwLjG7vKrk86w03y/eXhl4pFBXG60+YZx4TBAUXj6
EqGEPxKBm/EoVwHVi6sx0Un6NDITy6MSF/+PtkWk0idohkADLB0tNjJmy9+dxSaf
RvJ/1PaRdmnwmoHFr3KR/1B1IxtPyOwbRj4B0yIPtyrYObx6/L5iOZSoxyEoAFo3
4UfSg2ThBobwmdlHYwiy2ow38dS485U+7Wwqjrco71J13g7s0nKwZWxBwbO0b4pb
bARyA160euV1yF5UTq08QWSfi65k4+rqdmjH+KtQVq6Nzdn7hrir1pWXP5PnNN1A
IppGDjidVnCNQDz7gDhyWgyXvrdAFsedYU45qzk6YyXWsYuXT2oE/Ml173Afm2d+
C56vPM+orJlegGaQPhl5bArHrp9i9jldr7FUFN0pAgUz37Va+2UerggNEQlxMKgw
0qbJjcEE0wxa2Jv+3pWAOQsqFLgUSnr94GmiqVwuNxQrK++0wGiPIiKSb4OmWcgb
S6Z2UVnYYScgb6b8u37UQKJCF/IOHp2Io7X4wN7x0YaomHH2xhT2+KBeCx0jXaPE
sazoJ6yNAhHJdUzjE4U1Q7+djrCwDvlDlQLcaLElOz1Ox1WqNbwmMJ281DfCGACm
OTBi+jarkXFuvrPF0bQ808bTOpjapSW9fyh0lDafJHXdDEqf2pcVFam9uVxGUZoN
To/ZqnMfhaH9JnvYcIiVug7tQ5DjXJ8SdKbeDyCCuvraxWwJSfW65dmDLGgA3I4i
O0UC/L+Us02ikrCZKPAhn+PKeKjT3DmyZtsJ14QKQP5Zs1TrNt1OoGT1JnJNmV2+
UNecrJys/om0QkxKXU8aXgYAVRp8PccKG+hHNQYFRsp01PrUvIEZ7zLfcLAJKX/Q
CUpIfnA/YT4YKT45FgrdrkeSmiIS0mq4ps3ji9ZlEhrloeZ8sqPmChNGc/8At78i
OdqKbk/ZxGWliXn3cLEuvStrJ/11SBLIg0LR8YmVyRLC1QUHM2IuaQk/s44VXjWt
K8YwL+W4wInns9F4EDNuTOW24P0si4oTKLO8C+Vl87SujYLYERClTCUZ/MLLGYPP
SFh4tRFc9e9i9lDK4CE3V/0E+SYOk7L+naLs0CtDrxkvETZulwMwkkrRj7RasuOx
IXWRBTqdkMJBHKbPBZ4HQCwSC5TDuGVs4UMiHltnmBoHDZtY7kac0rNJJ0GkVert
iOvElzhWGyrdSRFoR21+kjjjDKWwYREFmebCjLAN/0zFMlpZE0S/D/+OOegkTX1D
gyLyu2pvyLIpMQv1YJN5Um2VkHwV0kXWdP+oWWbQBaGJt9qvXVE0HM2ZuupQU8N/
h3u3+IhIzbAOe4hlgb5DJdlDwW3AQX3V/PwXoXtxsI8evmqw5FMADSm9XV9BOKcX
xJi7o6wsYeEzCfOpdQPMe/TvAuU3NUAEbQbBWcKirXBlOVx/cMuk7VvPnZKvKR5f
rXA795S9Bw3lDHHxsIZIZJa5DX6Foi16jejvhAt/VR0KVR0wfsbP6ZMxEFInD6JD
DyTUdDIi1FvnMjqEEwvW0OFOiluvPopaYfxVFjD69Mdr0fBsr4Y+Ycr4M1KENJ7n
6qMQdOc/+WdqaTE08Llr2aLKzGAK0sz9qxettZK0sZvZNCsyeVqHw/sBld/oJLkY
zYuZWYZThBUfgFc51fxpH6WDkQJRtTQg8hrIyse8jsmEAMLv7hRUHqG7XjDrLL/b
7yjdfJf3YulXXn3pyYbH4OJlD5j5mflFIO/KFAGTJn3SRw9z1Deof7vHlQAmjHv7
NNhjETx0vS0cESsX/tqp3uB3KXio/rgzuGaoAuufMFZRtt+SR6Uu41Wh4zFF3hOU
JfHYVVRtc45xtDC1tP/ezQHPlfrQUFgvCIBvcyR9ulxaQRz7ILtFMHnkce/0fHQv
mxLG1vsk9gser5y0YxdLZTmaMaq3WHRvpySiR6hgqqyJuiZnnAeZrdmT5B6pwgQt
7PEk1Qo4YIwVlEbUVbaQdkrRtH2OVltu45qfeXSwlI4sZr82vQ0ob1ux8VKqUbbW
IvE1o4LGntv2I+IoyMh4YRqN2ufmKgStmqF/VbjVnmusf90IehjCEpzi1Mjj7Hzd
JUpFOfiOzsC/5Csy0y8Bda96zzM8uFXGjGlSlbP6PwcgfSIpGrFb3NXarEGEQ4IY
ozMP//yBoA4/YFxpTjP/iUTdmXqsBDyccIVPAHZD/U5A1yKaXOJiEDru/esoVDvX
+ya4Zqe7ezV2cwlf2YSckgRZLvvR7RDkrY86wv/WZ23PqCvtGd9SZkaAn2xBp0CY
wZbcEQERxxV4QL26rCglkGGIIK7hlYIjk4T44mBj1POttw1EJu+smCQEDuuTHTay
0qhEF50VtZgtTUiRZ7IdVBkWLwH2PjJrgL47YbzXSn82xxhK8Opm9MtwokQB5IZ6
L30GsGPkrOKKt9cU2csK+K6FV6ZoA8K7FIrKRhev1cmYKxBcEH5F8Fc5HAolO0wy
4uv+5dgeqH+g9WlnpatYevhSuEcNgxdJwyVoVOGW9BWVQH6+VNGoL5ZXV05Pazbb
DrUX77DIc2G0jMJ7wb0uhcXxlMMFUyqaD30YTY2rpvsnfGDaq0L4YmIo338WiLWL
StGdvy20RcwSb+BehoyaMBqFnm29WXnFH26iKr7oAve3v03KjaBYGgng1s9IaB5k
PsN3ifB0mHbVcYX9yB9PDNDznuY7Cuj4zPeNXgz+CBgvOESP0ZDKnPbGr9Eufftc
TrAJYVlaArie85ktk5VDOjw4Du0NeWwMuJjXleIIfCsEBlP3hUDZqKhlNUNG97UB
oAUAgqXQtGG+0sq/UTcnyVQ0QZO/l20ozayAWOIT1Vp/gpLspnmEu436og8SyqG9
XADbeqoCCYZQIFR2lOZdQhYu8YpdJgPq+o7rjHStOBA92/sTaQvGZb6cMKFdoM26
DO/2a+WsKQadLq8zYQw4sTMUb7J+PSB3tAJKICsO7Krn0WoANzR9Lowe3K3cJGx8
9LRtv4TPY78EDMGQ2ZTivVxx0D4cPYRp3EDC/u6Syi1D2GvHq/5/k4llNyI+jb2Y
m6ZmmUNy1+4WFWVZetK02XIYNBY6icylr8yfbDpP0U0qlCmI1OG+Px2dLUWceOep
oLg4K7swyQPuxemWArb1EPRKZBSAHe27MrwZPadrwJD38YF99fWBfWk5bPZDEimy
sXVlKORQIBKFfL403N5Knjwgi9S79fRw2mYyWAX6Taz5ruE4zyIYg6YRSCBKBEUn
N7oYuid2OfDcZBiGByHwiBM9D4l0sq5nVYmFH1GbTYnz638ijRgSZ7DaRsZsBgio
Y4mvUD7bs/u1hrNiJpy4DArjJkyAOW2uzrWXsNDXoTfwQYaeuIhDg3+4Q+gqa6gi
6Zp0G6iN0ayjRijiW39y3KEqoOn7MU3uEY8tFaLbF5s2uITnUpjatU0up61Y8VKk
+EQH7iGZEuM/TkRbN+P25/Woq2jxCs2z0NFOy1uPQ6yxWvDF8dXvmLApFZsrY6Qc
vTjE27PbM9+eJauUhA7E+mXAkM2tjL64VTCJ1Au3BU8F8fLmYxdHCXJYRV8tvv3C
YfpVX4tL+PVD1A4JrZGQgL3hSstU/8Drn3FD5UeAYHAIfGQ9SjXskMyOaS53hGYg
QN143qzqXERr3zT1Uc5f94dZ4AfBNvsqDIH7PonZgg6UYeRZSkKb/PBigHgvP2OF
KY8rIIUfGYcNrzVO6BjWXblklyQfYUuXEZHViZE1YJW5Hh1j5Qd/Mpge0FFhSSCe
MEmBTV7n0cuM0ULNanCtg8YGpUBjr22udqgu8VhpEwK83Bkf7iW2WZOfczF6bd8d
3nO3SajiSTUwsc7PsEu85LCHslmqt3H7KnJW1JuKReJecfaxGBvZ8cwAhNGKr0SA
it7y06qlYmnaojCwIRn/UIuBctOKowVz2YYdkRmA9BlMGStcy7lOgb/nLFLEzqdS
2BCR+vmc1QGEpLUuwQwEiw7hdoJkSAkMWDyjU6XQeRvMohzcPZm77axPUigbKcIN
/J9vwRrBKaLV7qV8mjrr1Ad2iDrYp3SKRvCA8akmEV3b7WstAnTe/g2U8dH2T4iR
9+OV3vltdKNsFsZkv9AjJ7/C7tmoc6fyQy3o0VRnHIfAgdEzGa+A9Lv6tOjGW1O3
MhKCyZU4ZONXuPRSGa+jtfo9fOPEFpxQVaHNNB1TZ7HIoKVaU2cBnFnH9u07cTN2
BhqicdlXGWOT2tSQZMXaIt2E6LoMlpiBynQLITUccBw1SFunANOpQjAGTKgTYEo3
xnBcrRBV2DCu+LT8XgZ//p8m2UhdIuPY1eNASf1OQdexE/c797mUpMVVZr/8E8IQ
jp7P8GFsEGpgzDMB0XkHh/H8rdMYB+w+nJioaZxMfDQpwqPnyjZsGImCV54JLlH5
fVrVdjHLO5bSbd7aAQKXhrRda+Uw+IUcXo546qD7FbTsuXdX/N59cD7wk4vCgltw
F/0ecsrRqqtje7DDzF53Jg25v9DD/mVsaZczWeBxqUeZpZqk6QrKrnpLyKH/CCr5
ZmlG3QkG9CfaZdhABMNggezMdoHz/sjm1Rfock+C+n22pglvNUIulHAPDWS/Egnv
aEHVJiFhMAlghyAd5bV5T/XNQYnYzYzAHpx/iN+XZEQY6UPFPd5BhrKSEYoAYx67
op1ynKTu4i4Nb5eKpgTgILW3sUEVwf2enqZ/hx+I+c+fd++E4OfVpZN4wwwAVioQ
RB1VpcRO/sYwzAMzyxYDQWC04kKt0IJ31xDWZOIZZuHU4yGiSN659VcXd4Ioi2Qf
bksWd726eBhMV+55V/Jf9zhAKHmGTLEbWb0ZAz2ERHi46VopxwaCR0u2CsNY866k
t1HYvaa2wNfQgGmGYlr3trLJAuARVaolh5yYLO4prtTFTg19Tsq+xACVLRVuuhXt
6s8hPw8ciadIrxy9kSDhlRF//ElYPZJyDooJKrIHtI8IfqQH2HGE0Gf5GJQH2d0O
N77A05MwoSbac3eqAapnJ2OE9zY+NXRuch4wTKIcg8wt0b+AFBi0ID7JRh+0jbr7
BRKBaWeaVl6QWALsdspmjtQ7xuj8UNcZR+9Cw1MaXs69c8fIR0YYHvSgsYiVDS2t
wuNeSs3I7GKXH0sB/05rfVE7fBUzGBEdagoeNessukfGwc7+u3+x88PR+7n1L4JH
QUhttbGnOIDJ0+ay5IjX0cotNHhQOwjsVzxbMul3lrGVF7aJ7ldZcNOouHg4zqws
VqcZ13TcHjSWD7OLrv4GTr7aJeycGYcgtvtIqwSpH6+MgImU3tg2cM+pHYSJitbj
IQSx5BCI5DuYfZ0PfsArNgTVmVImkHv8jnGmyaHEJl1TH4ULsUaGypz5eigO6C4r
YBngNzHEEg412SYUTGgeEvP+sX8Z8vQgGLuN1O96ntvwAYTiKGx/6tgOVuVP1WRx
Qtvb8iJc/b5UH8cBFz3eUU98Uz0Ue0CQBMPqIDV7bRy/dWOibymGkRu91MX9IoGc
pwdZDL+cl0lHxYqjAQQijfnOGimgNUR5p/rQDyQkXj+vb2ZfMHiFGpnam4E0ltG+
twc68dFPGoDqQmcrS5whppq0HaeM4TEqeFGodKK/SRyruX9jzt9Ir4BJhHfdQ5KW
7MwACxrEyMi5zpR5D5rzbStG8EV/hlgRTINHKrrXhk3v80k68IkTleszJFJORYPQ
BbAcKoamvmEyLMhMzWlvV2wJS6rYLIxsfYQo6M3ZDFiXzY5396a9/WJKorsq+en7
o2A9O8oQdNGZ4vrnlyFgfpxYe9eijlQnD3ZXl14CBJQ2wHR96hr3DN9ehr9THENV
hoFhKqm4nVWHznLsYOcRoYGYXyAFRdOPNNES6B+aZ11ucy8e/KT+CDl0Nl83tj56
VTHr7f1GMRnkls4VbtIxtcWdcyvFantDUa6YHMGVTvkb0gr0vF+ZjgbXBpX6CFI7
A6ah11mKQjO3uKtv6PXhDGXxcuDBjnuJzhN7hgLo2I/cQa0SgNxP5noFAufEAXCS
7joLEtaROq//umId/pMWHb6bDl0Lq7AplEu55ZFnoihTygny0pySHQhiiW/r+ujI
fm2tdKn0wOwe56cRxSwzhiRKHXdgzgAAfIeJXGVju2VGW38re6IPJ/jQ4Qn1AVDO
FliJi3xqdjKCshwIV1kuUrYVq+r2G0mLUjkl3/YdUojFcSDqCfe02f03rv6PIwm8
18I+EoAX2RVRlSVj5bE+2mAC1IYE3b8GrvJJ/L9nkSOwf8oUEGVft0FxsQsG/wtf
OxZ+f1Dc9JcUvJRp4c2t/9y9C0ay8yvb4idcL18jnsRCTRUqE3cLXNlUU4GGy/Wo
Ly66JOjTaPbl/yTwsCmR25MDm4I0kbAdAyqjopEBleLKqtbwSEOq0P9ySa1m+gFL
waE524gMsLXaBz+6LcmNK6MFasIdYzH58PZOtqe7IKAOwzcEgssHH5KBpqv+2Xs6
AFOOTzNhkr6jy34DFA+p2kEB8kRC8KxMeqXSI479o2ZoFayryOk5UtvLnfxa3Lem
5UJnercDpVzU4mFhuASwj+2eA4MrzcyWePUiD+4TmKMCwO4aJu3y6SzuVpYEzaNM
oy18DvakUYTzTMkGl/QnfHzSoztReZjaoaLozV/jyFA1ELCkKjXKBRMVF620ZaMF
w/ze/mutxd6wEMj/9SMCvrf+B0kcTF9Z5uHPKzB4M8kLKKcKvY0hpJ5QXzI+XD0B
ovJfJQsy5s4Dg7laNJkB0cix0Ke4auN+PFJyGBm7jf9vfbVMs9Eh1xTBCktCLokm
Xs4eZqJdQjhkaAG+vRCk25wGU9zF4LUq6VDuxQDWHWM+Y9Fn4n7K1ImIqs9kOh2S
EY2tdgke9HUO7mo8weiiC5Fa5rs+bocAKnZwjhLLJFAOuQr2M3UMRhku7wWRNMGb
t+F6v7bJJArCUK4hAjM/Y+jQBW4zjlGeaCv0QHCIRnIHKIFBP7oiPhhQJvnaNxQG
x5OZ34veIJ3xIG8/jh3vRJB2Soc8wdDb0EnO57UA4CnYiOuINal0bAeX4sGr4Eeo
u6hKbNQg5RqgfYh+8fOwz6L20aiF1ckBccvK3Cu5XKsCC+Y7th23kBwfoQ7Dw68t
95F1FtbnAMUgBTcM2+lxPOmoS6pJH/FravaR7wP4VigFA1extGozvpgqnA+Y7EMe
nz1BqhCe4ZgDL2vW0sk5MrwAmVcQUifWCjkeaCgKCzvPOIdVZD4ZnlJGrPvO3O/N
U8/XJ9EjfZcq70YcR1ajjeDpjrq7EtUML2fzY+kByhIevexfX9B+ge2QksEkNa7m
cbnghXKMZ0PRn8Z6rV120/KBY/MwgqWSlEKwK52UXXuvQxrlJkmdSiFWZk5auif1
z/GxkbQcW0/su5n+wX8F5cRuheEYwuhi7kxPsvay/NfC0axLulpxOfavmlqs2HiJ
XhPuznLzHDFAVJE8iK9Q+0Yx5DBtADrB9+O+dwp4Bj803TiC3x9xIblUOI+NcNGN
1oHc7Fo/jC57+PcPq3nSmqyM1Xof2OCoewtlbEhKVGx3Y/lqmVsHbAdg5TtJV1v/
Kn53dCBKYOv8m2kJvwWyg56hvHfAPWvFUur3vBktxyxBSfH0oVVv89VKHpldUN5w
2+0XtF+Vwk18+9A8ATO9D0dq3sGl46fKUskmWuYRePQ7tOoLJv81js0rD5IxwEFx
PzdNcDTDPCOzU84Ab22iER0361JfNhg3T5tIw1RLNpRcr8+uU0DBRn/HRmW+VGQa
7gSbT3ZNkCJobYWHxeYm0DTs5JRlLF/0o6JqFMhqoJEkrr+J1nd26GzaZ6xHQShK
Qpdh+KDKphZOF9V+Wd2abqrd1EF1TbwlbrQZDRaeL081SsYG79iMyD2xIiW1adBR
LEPnR9nTeMacmzBnFKNqtjpiiSTx2pZOlwMzItUqWdXMGTYrMyaintCrAxnvKnDA
DB5PGb+T46+OS4xpE35cx/EepPVV2fJUraS7JhYvl1wUcumsfmXg8/tufXbdRIa3
jayvdieIk4YOuYVQNFXCTS6uoJGmbWvDrtwr+o1Rj6mT/r2kkHLfyjTV7x0jJElx
aGNLcA2YIBT3n9+0dRTMOWbTMb/YTlr4KIUZ9oAtHKNOnYdzZ5MaUDGltgW2Z6fp
8RrbKoXRvcovUF/fe2gDzayE6AylcvGkOiE/UXoHzBxgJj2RL39WAli2Uc4wTriA
uo7pfpTNBNrn6W3Y1VAW0SCBdh926W/CAFVM9+j3VIR84sk8HGD0uyxKzAE71SXb
lIv6X6C1RRLGWciLaXjvTQn3hPJGnH8CqTuKWZxzLY499fW2HeVNj6fKUqjSUG6V
rZXlELaEqjmm8K765VSXKJ/kmdNPooFBIVtGXN4qpScyKPcaOOoqf7nQScGMeYo5
rqI8LR4BMPqZ19kHgobdyJe5jJngsb5fF16PK4Pe8lByyXYPuDEzuwLZuOK6OU1A
JQygEsvbIij5b9vRwTxk5ozrl/pcw//+LwaUHMtnqzNc6goLh6OhbPpwwjx+MNF6
5RR1Y/K0ZNxi6wYWsFPG/o9PUoYWV0RCYGcthuf17Zfzl44KEyIB294eCPiYPOyz
1Ux0Vo1pHmQGEE8gioAwb1BWeFM3XcT/WBJc4gbL9s5OdLWjRZzwmYZE1hDLvgeR
NT7PMzF8vd4vW+bVBF76dvB4xCg2TKihhWL8FsM2Eik+vWrjft8iKDIcg/eZK8R9
AZ66RAdenYm/lt1o9aeqdminRZzdW8/k6j3WHh5ciNHBExPVMJA6cBP0uxnb+eLV
PI1qWjWrSrcZ3ciJRNPb/jR+s10vFvopgZOKJSVbw6GKa1KDZ6J6K5Xl0FouLaG5
NZqBu06CURA4Q4nC1Gg2/Ok9P7ura8KFp30nTZiifcLITpjYhxvhsnetADEdo7qU
zUrLcX9QS6O8K3f+BuASUrU+wXdc6+oG8rhkVBVSfQgDjBhphH0TQnDk9wiCmkIg
3L9JOeG+UU6v4KBN5iA51GFDkbSrvxn+QqJzdZ0uyo4sL+WVF+GIZnCbbu1bwIwo
kIPZhihzk/2Kk9Ar5/tDDeHJMGo9+zRyni1L8xWwNwhxY/+ltTFz24DKUBWCNj+J
Uf1+lW9Iv0r7+NPOYTz81v9XL2JhMYc/K9YdTaWMFAAR9Af2XLVdilnrWam+sC/C
0tGAgDMtNeT/rltSIN6NZ1qTm0TyJhcv/6Kmd1STyTnfXXsU8v1z2qxIVYvhbUx4
rkMFZbyuWJXt/bR3I8Siwcg1kD2RJV6553bQE+f46W6GAhXkTp0XmOyWyNrWI/Xk
AyG2ZUQs0T3yd1XP/LxQlifGS2dy3RxriOIDpZnIGuW9dOwydEuh+USDGmaw3oG4
18TleItGMCHBUjMJoC8WbU8u2Sg2lgSORHNosIcj/2UtkuKTQtB36cw5+qaSN7Rz
Ce/eZ3x6hClOEplsjxVzDn4QAa9lflyL7NT6NIG4kjcltSTHZ3HZDIWHNy0Pmt04
HC+eznBGUFNSOjz8mzpyT0a95EAfPVCLLWWbaicUH719y2b+YTi1L5zeDROg16sT
NEzDeF8Cp+QgUyI+UG8BbMYecq2x5dMzkcTOjKm0CIJxVJwmFMK18rQTT8VlDNrf
ZPeqiREEEH8FveBZHc/kCbaJBX39Fy1gpBEJTCJXNlpdeJyRYaNkPOZoSsmKV1yv
e9//fAsqtqZ0YWvxFjgow+SK/awCxOKprHtnIInB4v3ixfzTnWbVTQeYTSlgnILH
JCTRdpmOjjPlUv1DTd3zmDQKARs0pNsvakSWnU4m+KtM4pJ7J0D75hGbmur8EX6v
kNI+E3P5QTArWGEosDQufr2mIdYVF2NECkIjrZ00Q6dt9S9agx6cXJwDSvfBK3Qh
6MCpZt6rCEZvlmbNCD9XzJERoR3X9SrospMEawE3wu7D3jiB2EjJeDnxoh9TBFK/
sTe8gMc6TKidjGG5qyA7UWh7H5da5x0sbvls0olXBKeE+xNYcddTC473bP5p9hHC
M6jloygNs2aK81WUj42jR6is41a4TKu8JfW1ueAZqzSFw3q1qcbZjYA/gQLwJo2y
z6EETVqPRa8HaEfQuTisHGd1JXS4ka2CSxAnusp2dS0vkDt/MSK5N3bAuVt2mfvM
gMyYcvh0DhIuREJTVnlhQ5Z00NaujmvM2YHtdaL9+MxqzTMM8hwfzIJ7NC+VERW7
JLNjENWGHa+q9Zu80xDr5YuYwa+w0TLhNOSuQpsZAQhWS4T5msw+iAorvLCYvcAa
T9tx0NQcApvqoKeRohDE4rEkTlD3YIDbs2/Urh58qdQTKLXKvUHBRQXdRA0wRTBF
T+aEw8ocr4CDuwz+8vJkw5j7lCbxoPCWzNSgVvniavrjBovpKtMK3wpE2AD7eC6l
I5jQpCqCG1vXZB3HYnm6CypWtq2DPbjFMWZbgDaxQ9eMPNllfsc5hodrxM9CH/5O
WwOLCduFvSnYKrrvDRP2MDI96xLe5FfyVBA3y0QepKorexH+6LBwQXzhwUFUdnkr
HjNZ7WukbuiD7bsSuiqwTMoIO7yP4W/zSj4HejwSFCQvGFMoI1ZBjQw1PCrpKsw8
OE9pDA/7v0KCn8xUD/0PcLFpYIrQ99ufkBczlVIrkiqK4O5JsrI/i16Qu/XnHQ1S
HeYYCaBH/eOFL2u7MefxKUtFOtKaN7/9DxdRKDXuoLXWdSXkSSY6pAniq6xthhlK
UTzEXvPxKtL2cOO1XZZ2zy+U11zFaWa90SDyHuJjVcoCb9OHWwHUYe5Suzb6VKx6
+tYK9gQqDNE/c51XS+R0aQ+oJgRWOvJvj0gEydh3VKo77ACtBKBARIvE7wuXVkhZ
VFspkUjmsgFgiPAb7CfcSNKGLgIaxwzK/BYGixt5sOGMOo8P5jw++2qkR8gSBxNZ
Y2v1/NsLGz1NYteGj24uoqq9hSLF7Y8aArqofR/bXHtgzjBJRPo7r3Yot8YWMpf5
3bJAmt1ksNGWumJy2DA20wB9aRBX9sCHRfXpsDqSCQhtrulwoUfu7X9qNSbuPB8T
7iijX0tRlug/QMIqIotl+a6ipd4/MjRQKhEbzxKppTFEcSCW8NQHfrf2o4pQQP/F
A2Ru5Bb9Pm/TP/eALfIaiTj+cJMVMNRm7O7LtBTlWKm8GTgjzFW0DwqublfXosmZ
jYMp3xh3+DSTdQalgIo3uoFmyCKFte05AAPYs5BwMrhyd6ciHKdqtS7CItGnY+ik
jljLC29yj8rPRcmmYesX39cTIXZDfoirDPHV6rh4UE/uyOL2HWFHPSWbe08oqA3a
c20LTyXuOsX9ywudfxwEVawEQym88viF3JTyd95+jdjjnRYMcaoaXa4ULSY4CS/o
+D/Vtb9CfKxgh1oKh4fl8hF32ak8RF0Uu76i3s2wz7spsIfkzuJid9hbT5HZ9r0/
aWwY8B9MWoOHnceg0H4mE+FEGbcQFGo445HkeioBLbBmLvsLy4y85NaTREILUqg7
Ftnq5PaORhYp7+MXQXsQ+30A2CSQ0nI+aw0MB9mMkKlsdvPnFwLkeZ61GAt+37rN
d2oa6sr7g3y6JDsLfWVXpr2uQ5S59rBSbJ4rPLLMWevWcDVlCr4DaWtkV8li+4WJ
NTLWPY6nwAD0TYZEmdNQft79DbQK6wKhgWvG3ncXWEbbp2t/BLq7pm8QChOj2agj
tOR7p966rPSICJ/SOkxwKIs9PAYbke4rp0cDHhl9xZLoHrupnqA35EQ3cemIn6Ln
HV3+zdxNYFKEGoiCBbGJn7AXRYz+GTPAoQ8NqtdtaHX9SC/mO7OG9NYrlf80jik7
KW7+bC1k2udAqt4XopOL9rmrBTiiYdtP+ccJzep8QuxG9OJTbt+fOorjV6EtamBX
oFuBqX3OFiU5/gPKYzHbPrKV9qv0atLf3q/KKc55fumvqNv/yhO/DVGwbvVdryKz
2NqVK2a3/AhPWvJ88twScTOmdPQxt5lh47cdWKeVU1Q+B3WJb+KhqrTiHixFqh4C
6y9kOSLirU2H+jWd4/NMzV3TCUZArDFK0IE0kjSQgNef3IawWNV84Ayj2hXTaFtP
Tce1VtogGsLb8BlOCRBppx5+POZbYIbkkSlx0D86k0XqLpLiCXfQT24mrlRA8MHD
A7qGRIcVi4eM/K8mBlhUxRK20axies4EouNGTxP2/cw6hoWGl68cEXttqfSi3VI6
mXxkP4TbOKTDem4IUxNwZv9j75015cNBs5VrkqQXax6wBnC8QN1dbDY8VNw4yUdP
HOo7f7xS982C/vVLmk8jhfT1XOvuQ4HiXf21SoPN8Xv/wZ+MFHhhQ1eROML7autY
wadAFKV2de8srAu5aVPxCwWwJxQ3TdNLvQU/5G6VBeuIMS56Av2KPcgRgl/zhG0o
Z8pDPtIwTD/7BLABGhxgXEtN2Z0HDoRpmwmyYHKqJKjzu2oBlvE86IDGcgWRqmem
5x2vEppBApfqol8exwfxbAHpQ+obJIuamAWBLzWFSujNBTGYqjfd2HNIjY7Uczt4
+vOFjMu0n+hX3Qb1nrgKF0Fc4h0HgCxOVTnmsjiXU2tvl51liVQ1xa0Eu4ywXtrU
rjYPrmJewvzvHCscrK4pEGFUzJUJ9KR9g/yrioidDjQ/5oksdhkcmMT7LBjEniiB
somKJq0eGfy2wb9I1ZPvWeaKXRW7VWWimZYeyqgyDcO3Vl+5vd++/QupRSgEriwv
pGfG9qY8vYdeEW3uxrVQvw/GAXrwEZ95sljVmpCT3HQAdlC6E7UuiwuTpqfJU0BI
R1VWvIp/sXYwaTUXEU/NYwMvFsFcBJkW4PgFKkTvwNsLglnTECQJhU5q8gAf9eOk
fdbacQ8seO5rqaP1s2eSbRrqzh8eSt67mq5+FJjgUNMXDipZ+4XQ46Gt7ZVMp4eD
Gp2EgO3U5i/iOleEtyjHHeym9BSR7s7qbRYh1MNMM+WBT0ctfZIg8OKvGLk7Ac+S
0NGC9XtF/SZoWMZKvTcMkXe0t6x0m6KcG9hhvf2hY6q6ksjfj8PqBNvolNUEf/Wh
wSutxtoEIjFCrpLgG8EjmzpS3akrKUgnoI/RhgehaCMryP3RL1ODE4Uz3TGwzft8
wSbTFNsdsomp77os10bRnYYrH1xlqWddZdmIxaH3o6nhjRzXvOHPNlzph9nO3Zv0
KZnoxkpALlHSiCN5NJlA/wmhYS096kP8AQaHqXpWgtQvldlOgEfzXwsagkm+TnXe
f5WECbLJSjtBY7F1gyucJfVWwBozkro8UJGHpEhD9Gj/FFQLTJw4fuEIYESutbVC
WpX43f5eXbbrgHNNvjKJ9YfIe4wENE4gPdowiBPjnKN4fPKhvgw6hPD9J6jwX64w
LuZ3uql6TqanMlxqX/3IquOZ4fhYkvapkGheC7aEbIDyTn2pkJQ/gtReSJ7jqdnU
DeW5WLi2unb05JkwezyODRpnHifgpYbz6r7T+ZOA3ILdfMUFsm08PuacGj8dFD7f
e22NYpj3t3ERs8RwSZk5YXhV2q59iE6DaXERoKqSKeUmUz8N36Fblyi0eRCSYpOK
QAnzq23F484BksLlCOu65hx4E5tea88+ga9Rj0Z53SmGPH5BVz+a5Rm3Ujv08xW7
FRw8Twvy9+2RWoCd5aQkn5u1fGLOkPr06+mFN3RokBoVU6rJLjYovJwP0S+HV3sy
MdKJnOMfnX9zomrNdEGVnadH/JPRfso2pJzxQeR/dT6Teg1XEARWrc2wXe31bX2Y
dF9OMm9I7s+1b+g2cAZqEz1PRKtcr5PRdpgT8oywk8tPUarLoGsjojHVkL+6XDh5
GvxaLUGeXiYv2nsaTrM8g/x/qPTwIF/B/r62OyBv6hnVzVIvx2clpDkAhUtV5zfH
o7MKOejtHpNAAIjKhLOGhxXduvd/143+oiVFD0RaXwyjW/dsnAbADVjH6NNG/mg5
IbfXSKjfn85cGwqPXkb0Z8583srb2xWIxRntLHTMxkxEep7mLu5MBtBDGSKfdGYV
OF3wU3By2wN+68B24oezUYtGnD2JyLmtLgf90efQbdUP2cWLqi275s5uLRsaGXN0
SJcobY1izVqC8yYG1xImjz3bN19O2iD7sVclDHHhoF8bpIjlOC1yP7nLYHudskEG
94TLY1h6jtXeC1ji5IMLUxceIhuurr1vFiXAToZqS+0VU95+VBlr3Xa6UeCWTR72
Dq3JQzX9PQ+GtSBmGeoRRU/4L3PMgdfVmm6tm/YgtrHIjxkdkQMjuD3UV4kUye3R
dS8RAXHQhRayQPWoWQp94EpNKnPzNm1KnooL17zqTNoF3XR9MXINqJr20XL5jo1W
MHvd7MV62L0g0A6h0/fQ5YG8tQYZ6/WGz5NOtduCt8WWi/uCirXlIUO4gDQKHUVZ
d5B1iH/bROLGf4dQsv/ek+ctaQ0A9ZbUNXhECyu9+popw6CvfwbFn2zzLgn8kLsT
fWwaS/cgya7SeeZhO/jPHOP1CzCPv7CjOEnx03J+er4vxwJsLoB+m/+AGhckUjLv
9ys/Ioi+84cpwOTFdlu0ZiJ9Wiqv6NUyas4AZrevnv0cPCb+2BHFnj9VvKkJkChi
7LvQSHP2mB5qzSuMCUwifmEw17NPNVvSlgwx/xig0vU0+zu+Bij2bsLjDBbUlFBq
Gqohf8jTav5FaqM6w49rk3s539f9ADcx39v+BjTmuDc/W0mr7eWL4pxHoMQPByyV
UUmwnPd1o7hc8aIqRI6PTlcNo4VlJsQu+eQp5u+tB5IBttkajkbvJDT9sZPw8/HG
eURJlODIJM5/+0qZYdgJTT+aVizrL+sdwJgjjeeJ4qZYmmHwoaKVc5IgCuHrEXIi
XHJjiERKqpwnGR8Y0qK1N2ABlYJwlQBnEJ/9XlTS42WRWBeojLIqBiUSP3oeKYJv
da4i9VlYOki4AmGWge/4trwoGt0Fb7rEWnwZ0st9kvmgfQwE8bsmwloE9osPbwaR
pdzppzn6MgedMvgnDJ4jwLKhn/2etIR9+3ipq28PFyvhtQLZ2Jjt9W/05JzOHT56
Wbik7fq7G1ESqqzcplT1JGw3DDI+oxjsUZkIYY4m2GE86uzYdP/HgxCrbDAvC7dA
w1YmPA4Dg7SWOzfjU9/0SFiQXyp5AadwybllfAaKPvTMNVZKAxT2nZZXGYMHQlay
cXPvg5v1awuN03J/5N4PSzVbxbvaxt/hidsr96PKtvDExJjbJ1AvKmey+Y7wUYMj
JiXRS4O5wy1KHg1CIQRK+H6TO9dJjZ4ahS4XJBCFjlS5GffyuaCebpodBgS/HFGP
vhbWwt5dq5Un9svQLlRhjdfg7rcqfjnlS7G5dfJnjrZx7Ha5ilc2Pf8kSm8cqt6B
GdoJDPhVo3+ZOs95cg6r17IyO24l1rPptiGXOqRojNGFhbf6WGtsu41VsAF91dA3
+s62ghcTVSLD4R6xUrrCskrgzqYPP1HbEjEG4XPcqbCWXHyWXZrNkQoG63H9X8i+
tKK7pd2h0IfHXLOB4keR+YHDBeIjp+dcthBKRaeSCVoeER8oRMPquGm4YPlX6Dt6
Bdr/4TnmfKLkvxCkAw4Qe+XHJcU8m3tp18jwn6xwstdY/OiFIbGVomqsAMIOqTkR
ZGo+HlHUguaO1vUr6lLvO3pBZqB8Clsn2nuRSnsSRoi/8ZUTnqL8/GVcMpXg3MJ1
wuIn7onEqFSSWmZQIhMXa+FnogEU+Nk60xRjaJBNWVo65Y8pkrMWq/6FOSbY+7x1
JITFgEf/WE3gQWFffZWhzIwHk8tNnIaKQ2dj7E3Rx5875WCymvKK4AvtwWgPF1SO
P9m8/cKykj/ySKFMRTj2cFZj9o990SJHhuU4C8eVX1t3Ou60jRt9loCnaMEscCNR
FwrwveZmBYS8fsxPDp1+T1eyZiOxxlp0+DOF+ZvNv2f2xlc8JcZbthJ5B7BKaOvu
k8Y0F913geHQ7C4phN9izFXkLgRGlDvIQQVMU//fJlGC/DT4libHm+nU6/a2Px04
gkPSRjCSmu7cTn4/2Ij5iKttt9ikXE4apd0D1kpInkQB5bF8h6Y5LdamWL19POmA
PMFSdNRrSHYSXt8BhTNiV3ePyysDMswBuQfAxFWcuRP6B/fSRVfU2hhoDb1KDSfw
jowwKwhYWcd0wU1HqS6WBk045eRodQq1CIEfkIQEcBg9ExotuGoikVH7/Cuev1EO
8NwYZieL5V7jUHV/afT8LqXjHLh7toX9ZuWQ9YDxGyPSxa6Ick6SV6ReuddUxm+W
WPG9LQYutW/24jh5psXpSx/bRbt1hKqMQ8Ow3tIc10lydUcz9t5lMsMhHHBQFLKd
PdVfhANSNpq7vKJNwFHcFR5epkd3GhPabkZGpriagTsUVFYKUO9gbDRBamj8aHS+
BSrvt8tGCHFkFxNA7j5MzERdC31m4+BSOalA/HpOiFw7TNkNKc2TLSpb01PA5UMU
LbRa9WQB53/8GPhFwvYJqvBaMAu08VN7L9DKJXS6WkZD49OQD2VT/5btnF2Pr3ZI
7UnoXSbpNLskL3j6txiuTthZkp3hfH48pBBlh5fvcCNpXpEPOAHORIn2Z7WqDgmA
HrGSItTxhODik9Lm48ao1WGBvjxfvzMOITxEIKl0z6LxqZoTbLpxqaKNuVUzWMd0
nEVBSz3nQPUV+FLE5BaGmPP9n7OTmmoahbbyBuoN343AMsOaQp7mweNMXYlW+lSV
AGBMy24z9W8KUqm9TMZrCiEmZAhlNBMAj5mAjWoaFoltH9iloeTgvghWUhjq+/Gn
xEsH4HXoeIXmFPixBFqfxDalYwBl91xeX4Fq5o10ihOqYQL5MehsOe7m6WzLuut3
s6jSZoSwkLAvIDSyPSMiUUvZzcHEl0d6PZ/woyyjj9yPWNOXnQK6XhU8zGKjySDJ
/VFjUfryAbKEk/CVHIW2f9O/Z4EPJHzCF6KnZfV4vbZ//ZOosbwLWDoFdS6xpl1j
xmfoK7lMaOnsY3Fcpii6k8Yfm705LedNNcPnRoJNiVPUiYJRvUBua5CJ+Zlbj6Ly
rdUDddVvLQZn/gnXD1lR2z7k/+4t/eoctr9p1s/fD7Uzc/ox+b4AIVkQT4fsrPMl
k2gO1RoMqut7kmhUxDwdWx0lvLMX5gkfupSehwWT9mesyRFjiacuyEMnQblCNjuM
eTi+zO8e7YuvIUXijnoANMv+rqcE1AoRKHJpT8gi7iTMSviF9nImuWbfrH2lAz6G
uwYFtcszlHFAfTQbLVOtUArcBYJwvkeLBcHaf/G0/u0XDUFQlpSepnl/DODYCUIv
Rfus7dTcHpJNIN/KrPmL81+/vEJkZf/UtcMBX8L9EF58VcG4KNG5xHDyC0/TYBbD
SCGpNj4Ur7WbNBkZ3uWTKXLBrcv/UWJGby1Fbe1tJa074mhjBtdGLitZIeDqSXxC
GOXmtmBG0rF/al0qt0da8ja6gMrr6ws30uRqVrIb1CRqXfc2fgj4hvFoQJgd1N1R
gdw3I8ltnqFZQhtAFjhDgfJyJu8PDBQlWmIFLV5ndbKoQHzkdXuMeZUVxotvkCyB
HNLW5MSgEx5zaqNmuM+OWuw6c6+G+pan9c7quSeL42WtBI2frGZ6M60+EPzvHl+B
BSf5EafIA1hFOVUqxrXMLPu7OJtncDrskc9E1tT3CVY+58viQozlR8nYGZTKRgi3
anzczpuui9oBQlJovq624v4i1h9xi7Spje4UliWiABO3L0ZTmZJAqHHvtAP8rKwy
M3CX68g9aRLpflx7251+r5/uu90iG+hdCrvR4JLsvDUVOxkJZoxst5M9qUZ0AYZR
0QeDQZ50BKhttcduDR8yhMZn46Ym3g+47EnMo96hqrqgxgiu/V8b4FiIq/EUOWFr
HbdSEbpyne8l83mTvqbjXFFJvvbWACxT0uba52MfG876lBVh42i7Tx6xkMO9+Iov
Pf8bP0rbr8FIBalLAyLxlO3Lv0A7r0gnOJoliSHYlc0ZEmd4n7CTp8JWOY2Rc40j
24iTBbxlahyKL/nCU2xLQQVBPBxKiJq9AhC8feinvI06ZhbKU0djlbDgZmxrGohw
2zack7zMxvZS2G7ax3AoSE58X8nrf4FtndulLqlWC8fRHX3giFqikcE9EUrzrMc0
X8XNNW+fmA7Ptzh7X9lIZyCh1yzbNoypB7h1UIVsLZSxn5+QZFtwuEL0dHp7qItE
3/nna8sjWF0UA3snsTqhhD4fSs9tSaxFnkWDDCIEydaaoEa8qDgl5SH5dVGY7OYp
y6OrdKQjnuT82Z5DfKOf3nPzJP6iMYOMLk3u5gYE/KIL8VbO7f5/JWJRixfpYqsQ
35neWAKNuTIJfap/F8uckyYCF15IWjx7a++WkTp8n13WB5FRU/7A8mggVVWkDJ6A
xcudIcpFNo3W01s+2t5ugk0o0AQR1+o+P65evV0eMQOQsLWjRTTgsuLYhxCqiGwv
QS/3xQaPRjtw/G7lDqvH916ZkRHMhXrHvWxgiMzfbME2n3U5/IPRfvsR/cTKF08p
9Vq0myWZveI8FaNUuvyJDdyxxUS4ZfBc6o+R0jXtMAuDJTj8s4WKXCKT6g4Oc3g/
5h5UlSvUfRMQn4GC9ANKiuyjBNSm+XPoetC3ZmLn6WlKiUz0leTVRXUs5LfZSmtm
le714/Rq1vG6DHpwMin+UI1y7fqzcWgH36Mr0RmH1qfvSHho3BYrAdcQL/vEXZt1
6vpMK4IimxudgpAPCoPsBEQzHYUx5qh0Po6tZhqZ25LkGD14RxwqNfTRV06qAo3C
5evzvUfK8qFI60T9XT/ie3E//35+/EnAFypDYGpCOfdi+HTcB1Z1v8mj8ljwrPxs
znIM1jGnbqnXDo7v0uW2TPDmWVoyCTd4HH5M7ip3ZTsdE2VyD9lwu9v/g7ZgTVbM
qlQIQphQZTWr3mPlFRMJ+qGd4MvW+iF3l4Yl+I28b6iCh/oEC9M4V7NZLEbP1uZG
HDIMq7VlSJt0c5UzigiCXBHkas4NL2CKHi7kYRqxwa+d5SaOAeCacEY7Je+KhFa9
Gb/ygixlfaRtkOT5rgv9zboQglC2mO1ZkZ9wVFbDHHlMb+C6l895lzy498dBiZrY
qt5ZgS8UotXLa9CuuXdyWFPLgup73NmFtEIUrCvb38F7vpVtpgx/e15b6Jlsgm6c
Pgk9ob91GyCZ3FnFtnCYWCa54ZzX8hcozvb+HiT/7jNuUOVzO58ymjxerdvEzdHo
0qiGAhi/+t1Sew4WwqKvD6jqU05EEo0mTdpL5lmDGewv2e/L80RvfWoaO5OA+5Ob
aCDrpoWwPdSs9T4t28XXoilCfN8BiSVDkygKrc7vbgfhYHNWl+cqfDMm1S7lQTz7
xeoUJETkWk8y0xN7TcbTzl0VeOEmoF+pHZkvS09axqtzobF6NPTPVUykMEgTU+SR
IBzyP8xuf5TRBCAumi1mJh4XZSry2Ba8zBOT2Z1bnjA8a9PBLsTGBUCA0w+jqEsA
BL4xtYOAR7PrRNCnrs92IQbtvx9oWvfpmR7bnmHKV+IoQaweFwqRCzOda6eghZgU
LwKpQ5HayGfCNokKIoqFz4f787/lKA98jOwTlV6nlPEse7wigvnRQtGHgPi1AXJ/
TxXU1d9oh7e4JHItSZtqaaLxRSWiHP/oTYjUi4mRyhWSCLu+WS4aCa8HMu4W7fje
HVzjwcm4pMePF4IRHMqx65qYsF7/MKpz+wf/ch2cXE41g/1neMuT5qWDqsClI+IB
+MxNwv/d1vYZN0FzTykbDbn8kmkko6+iEUxgHUbwKQl1fJ8ApA1OZSQxpDYfyJi2
3038wEQhsxbq7PZuf6tnQvjRIq/cUVBovHjRa4gR7MaBCl71PZ+coFgmFdS81AGn
wneyQLptZpuXrhAd1io5/hGJnFN1dEGjJ5vouFibeHUaFqZYNubl3SF/gwN5EkoR
6EseNch2yhLhtIUl/6fAQ7osrB3NTSErFCo17UjvU0F/t6+brIxoaW8v0qg6SsdJ
5SZMfCjaCGkHVaSAR6eSy4C8Gfojp/9gcjymI+SjNMVnJ+qrJaNG+HZJbkVYAYAV
j+mERvxpM+ERMFK7V2xp/uYbEjczwsSW5cHyFW1Gn/13bwLzuw7uGolQUS4wEzOL
N4aocDVXVVT+ps/FoYT3b5Y7rZwo558HgtPlQ2O5SV8pHOhF/rjjin93qH0Xgqea
DvGLKTZiaabvkX1Ep4vNfU9biG32/cQlyga6/2pSiVZXMuTHINbAL/NsvQ+6GnX5
k/k5u65O5ziTVU+Nwmv5oiZ9xbwUQ7MfjJ446+6t5WXV3WSpQGNBwrro9qatyEs6
bLI2GRsbLDJLxw/nrfEVg+vZfdFoAu/h7WFWTtw7AtKfNTRbVUksU3jSqQ8TOLDF
8ixWQISMdcQWa4tPbUOOBBnyLsdmLXVlfKgrc35pyJ2gZLAZKiPcwsNVDgdyTO0R
H1a6dtXbqplxlBuy965beVcNPYIJIejU3PJmS778QdPFQ5zKxhZMXeGOmTtrfHxT
WW1QXeZixdk7SoVgfivUGrqROrS5rkmT2wvIUN6dxlYaiECrU0UStFFeMb72BRDz
PTOzFtuBS3b4zCSkjg5V96t3j2ACNFQkYB6GNslsDmtp5XhCJtMGMRTtEHgUL7Dp
ROtKeKG79ZzNUEY4RhwTYPpvzQK0rulCh+jn7/Fp+7slZLfHz8+GFvTfveDeTKFc
VzBoBf/ueEazHeJapalV+lLZvb0e8KTOZdOLGreqn07XcB1idRPclXwU+LeW07Rk
tWKHWCr66tq4gztjdPQr11oG1aU7dKplcg9OYOKk7JqsZsclfC3QWVssAcLzJ6l9
vNCvhlvPT5D6WrfyvUPolbym5SW5yW31G0ytWVXS6ARTmVhtacGDBkdCwag7y53a
oJqP9gIE/UKAWpMo1H6ivzO2GpP3ZyVrXEl4v0Aer+W1wgM99dLNCnC0w+h23Lb8
4ri3qnUTKL9ZHIUn7o+rZ2j16eh5Ygw6183KCDRoLhd+aiQQJl/pcRZIbzyDmYmN
JFuGILS4OzpsFTbYQKjtk3G2IYQ9Jpm82iOqZ5pzPfVmTPL0BheLrU2GdFnZiZw7
sAjnYscy+vWZDbRSf5Hg8sxqoHz4JlwniKA7ekXvoe/xF3xY1GtMwfpZtueIXx/k
e9gWc1bCrC04ys8QB/+JfEhI7fvJ3irCrBBmjgfKdPr8MOBV3aO5eo9jbvQjy+dc
CMjo7l8+mkjTN8PalG+wvs2uL3ebyxzSmWKqEj1i8oAkBSqXezekHZkwGbUNfUMg
BhJAtkikN+hjjmYZaZZFsT0u5TvQovRtEuq0iVuNwr2PC+DIp6Urp7ZJf7Vb/dB7
Zq9rnkJv7/G65yuPzdY7l6cF4YO+5K1M1jHB2dXHJY6QYdOyYn3O4DzoQqw6WcwG
ragx1pGADZIHVIkhcSbaFuKbSVkz21vxN5o0T/2ppXJEDcyLAnVZiGiutqb5++qq
CEpK3lL0pHqfJ42X0f6h1chs4oqWI2t0fqNUVa4ZaqFgsUw4t8VKaKPh2htRP2Dy
+UhRaSl/HEiqslQGsFdx5bjjnISzizqBcy5qb6Z+RCgMF6kiAsLP5eeFiHLE02JR
kyQ+SkcJst/7xl8S9YGrOn5wEb8wJhp2Dq9lQ+hPxvCwhOmQdC9vdrwPpCeJt9I2
rn31tQXZZ+3Ts55WljgLAx5UtLD8JMO8eW/KvRHjd6UmFntFwcEeGPkLKX9STjZm
H0mGHXMSN+We6tv5gKBQYmCPFpZiAPM3n3eB7TOpjVWhQtbJrgxG22ysTVuDKbNn
NOmHs5IB13a9da4Qd9v05iH2NCOTMQW9fNFNYOslm6AvnsaY+O3Nfj9+Bv4fwdCm
sgxSAYJ6cWfQ16lV5IXrg7KB/zVzqbDJVXz6bn+oCUoie5HpMwQEAMH7RasvZklF
W5pDk18lesbkPq+i4/iC1N5/hCPOsWw3Hs7kGwX3B7XqGIpQWWIkY6ThSifD6jJV
0z5u/Bgo8Lbi1Vm8qqlSoIUGR1QyZLEnUCeuT5kfZZYsr+mn3GS4xKp8dnd6k8CA
XIx/2dDk6Xc+cKCRHvqwZcX81O8uq5b4y3g5/zQXBeaVxiUjc5jRD/sZmrpsOw4o
YGEGFmBhApwYABFWPaSHP8FK5E9uB0DXHng8RttO6NunswRslZA+5SWnJlOtq8Uv
VsZMPiwn1JI65SOQ8JHCldE8JFCaAu8f//vMTqLnENOo17RSssWZABZmE3DG8aT4
bOL10HLDh2C0WzApIL8H53Xt5Dotu+Gie7uxWsWCJGg0wErdYETDZ9utdbNlMbEp
uC8T6SzbT94bhc8sA5WsdMBz8ypfWjdhqNUqg86SvbZiofxxiLMqLXdV9fLNIXYh
lDi0/txFXUnXQIhFiLD2muIY0nMJbGBRnAxfculf1niZ+pcaYx65p+i3L/TwdykO
PnLLDduJ7m8/9ENVjdwKOSgCZSe277616nsvY0Mq8WSTUfwu/DCqVZxwzGXAKh/R
TVH0urCN9qBlipXEMbKVJDwIS6LgdcdYAIuxo47MS8wmkgASVVlV8aWPHlWmAGvT
l7lEq+m65doWtaf58lESE5enVbisYPdOdh41YPdYEqD0wv8oh9IFb7OUR05VxoPw
4CLhUx14l/iardxsuxw6lYJqFAvysry4/9jSOZ0awQPus53l6whUPEqE9fo1i/MB
Gg/zAf1IeQi0/3AXgUCPEbUt1K31fuNBTeYHL2c5z/L4UXSfqmK8eICbTeJb0cuh
G1+5NwGYByVipgFCtMEltQyZ2JMjtgUGKOhTgG6yUP8VRsoukwtMBycPw4QWxmke
CaKexK8yo3s4eJLshXIPX39QFJXPekaE5QCu9nZUQuu2tj4HdKaEZ94/kHWNwBy1
gQnYltb89loqWg8V9N8k7TQIUUJ5uIh64jFRtpJsMWtLqbdL3DoNOe4k10+METf2
Efw+nIaJLvnxC4iXzU5Poe/r7fksZz6qMWU/+pUGcffiC1A45oD4Hd+KUWt2V72W
okHfNQKwOEV9O5eeSSOuGrLMyqB4WzzTO7FM6v5c7gvS+KFxDb4QX5G2etfr6gUm
o7rWDXG1EWCXKAb8945MbHa2zqGFAx6nbZxW/+ChXSzS+fi3mybOTnCcQ59BSrhW
ee89NZ8qVp6ivmiG9Tk3THiLiFZVJ+o4/D5QSCq5eJFSzihHKERq4Rk/WyUsKIQv
8s8cevoFY2CGdCaIRNIYVE6OjyF1K4cySsDJ3R9c0PJs31SkLAzMq19h41kYUkKN
2O3zYweYlSVV+VNmDgIlWnqII/dZH4yWvF/QB1Ol7DCE1TuKdBTFmYOdc/yYPtIh
phohI65jdjFn6au9JHUg4DUAuBirIPcHGWorZci9vYo4gziZnphNpl9buaBOG81D
rpbWRUSb8A8bGxaGBXemJifOQ/tDDV0gG7MQ9iGfhedav5gG6yVaAGCcPSmIVei5
uToBJLCTJsyv5K83PSHT5fkquHlc8xMh/g0wi40bGFkVhPzXaBBufHus0rrapGEk
60sEBCZf/agKpVVnOtDRRKR3HJzgreGJ4IfIUGQsRwcMHxUpZgIpSU99IfvUV1a8
+boR9QVPKeC9HlYvfOGtcb7CViVbIjkFINCqu5f0bL5h/ycL9oGOQ1tWWCVMT5Oe
NGihvLB1c2nqm/6j7ALQUV3SvcaR+n+QNfwxrD1a1U7t9txXDiGSCjMIuDpJzrOT
Dly8QvF+K1ty/O2ngT7GplvPWDQVc+btLMIWf94k1Yriieun5RkGGv+OOJFdhLMr
ndp7tx6YkL0bLDWRxv+jaqe1k4TRyvdIi8/LbUa0Q4NMhTNPWBkJtWiBobZFzC93
8FtYMejEYCwb5UDJHw7/PeTxOhdD4qDvxYoqbvwrPYTn4/MHlRVb3y1RHdcPcvFS
HxNes6+hTSoxY+/xRJqXHxWMXDFoUEobr3dPPS2hdHVvwt1GOyLCyPeS7xJnoDBi
rbw0VkuDUZ24gAt9CgjeEuVtSIVY7FObo5LeKKRmUPexU2Y9U4GhFKZAMfJN9VYX
GzsP+1RvwcBJlhdhAwsV4jZAY6/uKVteMvkpCkELE+FV4gzvJoF8n1x3fac1ivhj
ElmQHTMPu0C/LKr5bZMm2L5w+byE7IHQaGUjxACPiDvP1hemE/y/YwrhDnqNqekg
JkzwobgIAADWsgMcEDmy97Erep6+8526mNDpvHKbetVl6Mgo0zExHASyyPwriyPv
l5QxaH9n7gdzE29366PuU84GAY1/3AXBLL+1/Q9UO+ib0F4HVdmOLjvMT1TgEjMv
wvY/+NzhJFndsjty6rCmhb85b07ADvYmfdcgn/k5eyMTkKFDd5DSazs+zdbOZA5S
UbDNefKogIK3gLUVFj6uK4+qsYn5VKqYM+Na9QCxTuGFGCOqmffek6m7C1/3upB2
vyQhNHaUO2V6OcY6eo4ZX0Wvhfa7DcHKHZDD44THsQusUvoVBGSk0n9IT+SjILBR
mYHGOMl1xIPHDpdubG2nk/haOhDMLATX9wrkS/6b3xXyQCNEH0bNMcSX9cEruBop
y06ptNrTooSEm296WiI1P0wAJvJep/KXL7Y2KbZd8k5+UM81ZJ9F4ybbtYyuIsoj
AvAL4J1xCStHR3NvvpktE4gJgQ85AoGxCSYLmluWqhoz3x67ByvTi+4M1qFp8VlS
NM3Ztv/NPIrkq2ChO0dIT+BuZ/sVBhREn/MOBFd/2y6Ard1S05bkBWYf6TzzoXF6
FdouSxB1u6Ab3r0of+tMTO4VLYF2Bk00/un4ge86k7FeH4jUWBvdtIVvYWWw3Jhm
z2ZVzMxacWL7EGuc8IHeWYOci+HiG8b7szArD/BWaDXCjjAvfj/vCuVl4CE9qeTn
sbDGGn9XiqsRXZGy6pGbVB9AlvLYh3YsgKvxesw9AX1edNwZwmdbfuWT4twNKqoa
+UirAONRgDy5NHg0WlNzW2z8cT1oZvNnWc9AXj5UYaXwDbkkTUgvNFHA+r0wduT7
rnORZ2S3habkh7lGoetqUXjgrjkZb0/loqDAiZvRZtImvE+sW2ez9vtE2GHmxq7n
d/Up8FsBfIRHM/DWVjTznSIWqyN+qXkZFaYYna+gGgHzLy79ley4E2+ovamiezl6
SSDiRzmvVgIiqjwNAv+6yAWvNrANMLMZNjosyJLxREwrEAr9FXqlQIcow36uXoKZ
+vynIM168mo59qCmKJgcltuRQREa3YiB7G+HVxsEPVlEwnSgryhuT2r3zlQ7Ww7T
4T8gjAOPNl1kWAbjDue4WCi8v6J8OyF/8oC/VRzVrHwZKPM9q4/7gu/HHEI/dNSH
8GIcahRNu4pFjylOkZYZRWwjrGTiP1XKiqXsSWYmHd4xa35Gm51QTHy8fGCr4Bnk
iT0l1Sn51EjRFQIGur1tuV8+PkmGshE6E2Puj+iORQ9ysLShIWrOytmtcxc8UkWs
VK5zYr58M1pj+Cagyvaf6C1OGANnh/X7NK2N/20zEBqLTncAkErD74hCjR0ZtIRn
VEHEwMsBXT0C/h68U8eTukNiXD/irwA9odu+3udU6ArZhFW3ZP5nArlPOQm49RC/
A63Dd+pGUenv6W48e/fXBlAqBrSb09lTQlU0VZXEqsJ7MHct1/QJGt9MbN5P+9gr
i7K5pYU7sXFpka91/+NQXE0ykLCvgk14nqw/QEHo38Xu64zuenYgaJnqgvbEl6gF
8KUBgewywdE5y4nrfY2zePRGUY++V5a/QPMOH1+4C+r305Co7lp5yhUZLnQgDnO2
5kyti8ie5RSRvHEkcR8BAFks4XGCnoSjuJmNcZ6ri0iCYYpqqJvsqROM3dJD4qcp
FCyhhtOFUZuO0BJLDjNMCXMSbkdwgStA6G3/mHPwsZfWQJ5/a+FJCgCzcVFVRyoN
SbiLW+GblppJpzHKRWGT1uBsjR/WeMcJEt3vFvAmq++HDmOtruJkjFq0dx8rVWDk
3iOl63oImFTEhrk05K/L8oSaAiTrhh+uq76tcsUr0lUlM2m9AWXqwbs7yiP9pgTw
nR0FX9OMxZgk417BcQV1JgNy8Ugz0EqOp1oX8kOE2PdDvHSJRDIaSZnHMzOcSDvP
m4M0m9Nlq4d/D2+QUd5ux/jxhsGmtjgw1PZmFREE88eCEWMfsjdka7Y7VYVhYES9
so/bvwpC4woF2+eP3byXWroRjR7E9kZ/gBdJm5xxygw7NIaHhloeOaV2kyze1f6B
CPuQKaslOJnXCa6E6ciIVDPe/kU+7v1ZJ+awBbTYHaR5xrG5csfXhFkgUHWjStEs
1KhO45o1SFJwc/T6hT+64f5AAWth9Ey7sNy7wrfgHm+ru1cc5Ws+Zv/YCEr+l4T4
+DTz8IPm5jzLOxP6Vb61efqFRceZKlvPbvK6/E+1t3xvr8qZjg/NvvLdqrFTLUSA
PnKpEldwC8Habv8zlZCa+kgQEMSz1XCxlo5l6tCZwzLHDbzAqc4U8fUCSn7l2auY
wFzG8yKzH0lKdcf652MKxGk/6xlyNbUHsItpU6CMaLBMXqdo3MVidDHYPksGInw3
4+SNfC0W2GjEtaaINKnrlM+dhFctfSmsEBktDk7nlMPSx65CYvg4zGpmDCMVW3/v
rwDEtvvBunPo0DUyfg+lJAFg8bHZ3EP6Tc8/mE1hgc3ie6JKqheTh0YyenjqIXle
dYzX3KJbTT4Vjt5YxkPcOeozKjXs8CDbSR58QH0dTi66LUsoAALDtrdte36lGU3k
vT75hPdl7FymPJZHlLqNiz68TRV+NYeGzlSpfHoB6IcEEO46ZE5pvhW/pFnfHcwa
7clyO69GK9wvtMaS3W50wPu4jGqobR82ui1jA5ytaL6ZRZwA3RIqUQS/6Cf5OW2a
9aSo4Q5P/U1MxCboKRzpZrkUZfrigs//n3bdyPAt2tH2iRgBLuE7I4MkcVqL8tgh
j365Pu8sCLCjbKUO0MlJIeMsG5DFmD5ShjuH5/EYiYZeMy9R/CkEi+YOoxGbg2t1
ZBPMrxuoS5hLC9UF4TNgnGWClzkThCrwOBGh/InQKDWw8g0M20TTe5Qvc/rnoKql
7dfQ1IcuIj3lMVa0VzlreGzBqABagGNsoeF6FcnefMWrbfZUkay1omWXt1DRL8Ct
FubIgN6TMdq1PsWU8ovbytEBhuZB1Jhb9DHv5nhL9MykowBhDMdaErrgbOKLBxeX
NcPQ9A72U2jUYAcFxJ6t20B4BduHVGeupMcr7v6gizse8vnkugTYWuGQnJHzj7Mh
QAbcT1zugRKnOJKo7vJ90rZHhTRics9cx6sunjImgcxQIXYlrma1cwISc8lf47xD
3r+dEkZPEYObFRkpcxvD1KgmLjUG6DG7chWgihPZmIUpH5MV/WtWqrBYEQ0/3X2K
BSWtwyelv0jHJOKU2rjtd8J0GGZHdKoh7sLC0xYMTY+D0JioXn50rnRfZsNbSYuY
+eMUajbdPvOuJXwkwymq29jQ+CjoOEmMC8Tg+m3Cq8UtywgybBfPsolIVR2PNXEG
tUO2IJ7ZD4jUFQRkpoHwBSY5oH3MfyE7I9qeCAKjVRQEefLRgnleYgTpMee7S4rl
MzXzFvzsPp6kibO63StPv5I0smjqp+TeaB7onKydcXjdse8yUSKJhrLkf3V+jIqC
ykLtbPqpC1yBlBy0wt4jCq00IHc6HVssv+VAo00XkxU2MjsOEEm3qwnUpEeOSqqn
Qz8l2A7fOVMgjythiu0/KSOdvf0+nR51TaBNImHEmwTTtfQ9q30WZpXuuOhN52HA
ewRiG+0x+EVgFBN580sL/7533s3MwDuOBebxiNa/TS06EqJLCP7QAlciUlud4Uw8
CY0SO+6RffQFrgfe3J+U43Ay2owVqPkiQEexd9jGxeOcOuRpdfl+RYd9gsdz4aPA
+kz6fYwMLIA48T4xxevzVDqiCiel/NSiS/HvUetcZiIZQVBDQMtWpApAPi/qAcvw
HJfBgDm2Z85qxXfiM+VTug5Q7thokiEsR7V41n3GAZbZMWpdxCpaQr1swUpNQD75
U6bDZ3my3gUcJaahn8XtjVupSS4m9jmjMdPfA/NVs3s5yisIfc4SCiwVzQZEg0FU
Y5Rrhfpzs0IFdahsN4Pyh+TTnsHMmurGdFB8AavGHT+1hOThffElGaXl40Ak2TMG
wKGBUyrrYWOauf7n0+RHGLr5gXn3uOFn833n39ZI6aqBT5sC8zgwW/9ZMNsbHy8z
XhePNMHNdy7ssizzRxGUqJD383h9MGurU7CchyY4PyxInHeyisxin9Cqb0NnlxTg
hbmIaKE3kcU0sqQoGFEoe3W0v0WH4RuqP/p0z7IZ75K3XTG6I2xVKLWwJfCEyMPQ
ZmwNf5cwPiT5V6kiGJrw/8E7ctNZErAYuV64+viP6VDjod7JB4noUc4SjFkl0xcH
0A9uwc6g7ufT5FqWBJaZ0BmLw9rrgrMV9EFOjyt2AU24QulGU8AXHE2j7OuEl5MY
09JMCyHL8H/8dGQa3lsB9wlgls/tivgJvl+8T94+7UsfxHMLsBFL5r/IEinm6XnR
aA6ONQe7epByvrsaqXefrBJGW1LrsGJvKewuMEn8Ile/lJjETfdfpWiHZMzgkuCK
BkPQkGyKUTns3R/jpbJqt9H38m57LgWKwYnfvLD/Aw2MGHeg1UDYSeBnaA1z8Gsr
1iiNNghpet4IWNb8e2T3jhxGtHaXahqxIfVMXYGU6h0ApzmZrJyiHEIc6zSsvs8J
viurtpKp28TY1Vlubv5fuoJ7hgb0SKIyGzAOH8kbIW0HdsyA/7qsK+ST1+p7Y4ON
q5WCdV+2xuhzZHGM7UvjgKdAESbA4DVi3m2SaVvrzsvKzax+zXO0eFYq9EG6Gl+4
afKFn9LwXhrFDK5OgzHQsQnZkpR473T+kwb5r6i3nIhazVwfaFZ4GCkaMx3GlobR
mdAfdY7msTZ6Mo/gYHsEPm+Si5Sw0g4RKjDd/KC/3HuKwYbbpLfLvXrG63XN1SeQ
2gJwytmDcZXiHmNt+4DjPZfFNG/jizeFcJxzZUt8lM5YVgwLR58Hg6Z/Ch9d6BAx
Qqb3boaxLzObDkfT9PoLqcxhb76EJiqYVwQpxNlz8NZnHLw6WTI8oXlL7x59E8a6
2xoWpXfzE5cCPjUqHCWgbCcFJ1VLLD+tAFLhgfmruGjPVsPIHTk+xcweJ/AejaEG
0u9AKj0gYeP7fWEbfktivoz0Kp8gW9377IZlmXw2gJqOR8oJPhmcr2+JT5Sv1KaX
BQFMQTYPUTzaRDX1eDAr2SKVUvkI7yv8eON4tPexHfnCnjBbmZLAredimnKwl9JG
yO3qnfDywR6p22PlHM67/o6G0feAx30JZd8ibEodzUSDHkCn8reRZEHKIfXr/Km/
brDgKABSV5T2N8TrIo4cDFchj8U1ABaMYk2s9SVAo+DBIQJVEW5g5UEMq9XQyIpU
GX6N7m/+FGUKV8EO35iLUoDUHaOg1Pill7FzuHW/mlxZbwCN1OlMMW/RkuGAD6MT
uF92WmwxLhI40n4yyH0hXCS9VaXvqNRU5aeXYjkn+ihXK9fu8DRAm4SXmiP1ZgDe
H9Bbb28ZjAAifTSmtmKQA9eAeXnChRA3g231g5QeHgLSZMo94eKQu6z8KSh/8mfc
fc60hTuyZmJqDMbGiTPTSy07MhsNiCfGP6MEpWV1swYPO0cJHq0TGstwNUcA7DBu
euTweYVeNuQEyT2fuyKtuCGcEAmlLaVIWK9SeITZfdawJbysOjfwSsE1UIAaiis1
q5FVLbbm1ql3ci6JLFdrORTokxIDQSzAaSnTOQ9DO7N0qphh6fiavDMXjjjmt7AU
lDuxGHkqnpapyl+Z16ygenHrmABf3bsUNG7jx/RpKMH5Gs9wMwIyyD7f0wfwxawl
E42bY2QfViR04af6RXwR3FqcoLRdCktfs7fbPSVyfiFuqcKX5LYd87aVoYlwHBO/
DQU28DOtSVCEksukUAJE/nrUqPkYUCIkoZSDYiHgV9ge/O6h75s7CXehOxIaGTuu
b14Sjv3IX8r9Gnalkv3xLe9m8Gt7i0iyuj+JkZ/leixMdgIY/tOTC1FkoOg/egWx
vHdpdhZ1Z3Fzjd7d/wQMaYgf5V2EkHkH2ua6naDjjLqNs3m8cHBJDpCN9WR1hlx8
QBZ8F4crmX5tSroax+FSz6c+M/tZiK4fvh4aWj14NZ6V/LyTeZHdLzsrV/yj+3ou
qsIWVIndVCYhRVhp8MtvsZf0a4LstgyJcRyWBiZYXnxom9OwtrpssbTsZla80AhQ
/G0k4zrlVn5iSKDTtbhGaDwouQxIQCkSA9htV2lPwXkFAmCrYLVdnpRbd7LELVKY
FouVmGNKZrOYXl4nbVTpg6R4d1ZV86NRommcnY7xdeMV8TGqXefC6+FJCwl+wU8q
SkB8F2ePjR7G1tTykv1KUPTmD6RzB7is1O8/18Q9SuZZ3qEUCiqNrIHro+ymgfJB
IWi/fjYhAn+HLw49PogvFHJhybp9fmvTfddRJHFCo57+AuDO4n9sDBAv9K94aQad
9cRK4WK1g7zKkGg/XI+5aPzyUk8kl2eDYZ3TCZZYx7CtHDnZSkXavpFPNWaqTGlE
DaHAHJtkGzd/SxBtyxLunp9iyb0Jp6Sy/zW1+WeZPyogRiOwhA8C6GaofBn2bp7D
2EWYDElfoqitVodDYOZU/sVBU/EgM+85GIemSj8wx5GRpxjgFdueMrCF+KrT5vdw
I0S3i8mhURumFqbzT2WyjEGtD7C9cpjCGJmOmYvIFmaTRRKyc+J9phIT9AU5Oic/
eYj8K2rk/YTLuFdRxjnLHc9AIgkXlgukHDhlO5Q5aXna+GBpkfdt2I2E2LP6T8fG
HUFLcA/GrK+rHJJh6FG9evFp6gI7O2g+Fio5p9lLZZ5nkmyEp8ZnkM6o6YZzJtq4
ObwYfC+B90t1egPNyCphcSrv9YLJXq2jm/oowQt7+GotdRW/rKmMiV/Kmf3NptAd
01gc2QkuOA7QjaqbJxYoa6OyQpqWlWG0DYtGHu6ur5+Ynn0yuq3j0ep7cAId4nqC
c4wXG0uQgX77xXKzTGjlSw31+K20qC5pRdBrwN1gxElGX9XMEZEUjSC7PZ+UDnIq
q+WFhM6mfaSRP9gpqAZk+KskwN9tHHrmjsj5TMPON9jeRwiKg1LHIEC2uaWC+81G
3geITRAgYsf9fVNXPe4tfSThMefHnlFFTnbAUqiBZz2AG2BUngN0wwd5sJVaA87L
+WMtRibUl0UxxeMYlEoepw2sNtHlSaqL21ZU1lMb2WlsilBIn3elfLsAez7cqOOB
dyDoNZ8NAuHk5nHYJuvjUkyF9NVS68o0sk2Knia0oXrb5mAGDategKZSteXaKscu
kVT8Rwx4nYBBddpdTz63LGqzQQ9h9YEMdxDp1h3Nb1KqYTypi7WobxFzecrXdtO3
IM1iexmxtrIAy2Ux6tVHz0S5lm2tTw0ZZbilGaJFpr/dQPR+oQWJ3qkxk3gXvVPI
YHHT1aMAL40jDBGRHFW+giXVdcqYT7p+HOvX8+65CeVt3fhrz1vIHze/AnBhCA3E
eX3lSSyHV1DDVEwZkIKwclZN2rQ5sSdFR6w800+QdVnrXuA9C5/pTeiiDaSIEJYu
HHJtGdo6CW4cP6g0+0tAbmcI2ZgaQq++NosKC70IoxwAhf5cMKrhJAtgeunoSJEt
BIoP0sbn2kygQMZjSLVXxZVe0B3eOIArYQQE4mFFb6mFL71VT9P+wUC4Zte0QiHI
n/XrUy30hqWnyKXkgnSU2ZOBcrruDj0Jw6hGcg6s4dtzq1jturiBGSZPXOTMgQ9A
ARFeLsw8CuWlcLOMgHR4E0aGv/hUsZj9pdREOCXC0GqLKclYHP90Rrr+iYrZmU2G
+wZL2gwPc9UNZeBWoIW0LmjhjCLvm6D5qI8QoDaOaUsPaO2PhR6th5s0VJFuRiWN
UmVnK6XTTD/pOI5ufWQQ6HY1xWWCrSpfgRmqT5gc8bW3NT8uiA1ULYMafZJMKPGK
qG/vQlf9P8ovl7AIMu4aM2AXRCGDgI9mKLRyjvbLSdGG3u+/Pt9NguJYvgDRP0Wk
pYuO9KmqDoqsUQ+KZhDFVBZ+FCzV5cXtvw2JyteZNzpQXtEdbRi+cbJQs+6Hguv4
6RTn8nGTNAXb9AxOzNZNzrqEkCg59wXhUOV+F2qtreAoPKXU0SElpzdwhxTdy1Yo
ViBzDKjTjMcg+4Vc7NnYAnVwmFx7B2W61h5LYnZOtkISVhIMTTDy3GeNRap+gvJy
kQQrg/LGinXloRBGGFjxz/ShkRLewfIb4iwtuDV1AeLxlCJfmV1UsKox50WJ+cWl
8VnjCi/XjZtCCvt1wn7DOt9Flyg0Saf+1nGoE/ToqqPxyeNQ5AKAKlYPTlIW2Qny
dn02/iuAScTyik8tRDRK5h1s2soXsbMA6E6NdPYUOReEqxpU/GH42ogADcRhQjRz
Fisopz/ZW4iEI/pNVEVZoEvxOucnqSGdGR9qV2CIJg2Das1sfQ6SlLuJaKyiob5k
q6e5eA+6vIX6PPoPgODJAz7MEl5X+wM6OSCnEPLna1AoKU0ycqK1+y37jJeR0EM8
4XkLG0uAIrpQLaidUG9s/UspHrEpwWfA/6+vWtvk2lgAbkBULn0HKXCVsQvBOCbd
/kfd1zH3LhEqZvKAENFZpvPO5r7kDkosvHCuJIZnYHRA/lCYA7nqSFS3+2sbxBQq
B2KGtZTlcx0Df0XQPpao98tIYZ1XXyFjou0a6pbDvvD8oorSTqea83mG4K17wvjP
nS2ipDAWBn/ekuTw2Yk6ZjaYzNycI+WMa3+L9Wbjn+CohOUHpYfTtpUPqZR7TlrX
LfYfxkEeZDWF3hQxNYds39yS6ErSiceSPTO8pPDHOSA2EKZdk4ZGL+3QHIsbcSst
TSWwn93xvblIk7BzPHtW2MCxYI7C3CKasYTJOrqVsGrk2me2/psymhMvI2bMTgxx
o/b2pLxioyRYNcJVhjYPYbsgLEvSK1AeWGtpEGmIl2mafVSN8xJ3vINGPwF1Tump
GyQaWCGKk79VtaW+fTGIdToBLm/QJK0p0ajg5d+IBUVPAHDi6rPVQjqXIivhd8vm
Z1G3h8uaUiCnrMk7QZdRwONJ/nr7LdtrHcVlazmPyj953Ikv6WmwTgmpstR/W7Qw
4shNw3LpZ76t3yZU3/bK89ep20VLQ6RSC2Z0TUQGN/zTp5i0M867PrHUDyoKuW0f
Ma9FhkP/cVYGVRgstv5jdhL3LYHk9QO7B7H0WjkaL34BPWSKvBtQjbZOPBJn47wY
qL5txbHtqD3I5eeU25M43JhN2jTvOAazDZ9r5T/VqvIx0aq0HayLZhaP/JJVffxD
PWpaOVrLVqppz8xHP1qIT830vb2o0xe/ib3CgiDyjaOyQo1H1/QPDae1OYoGEGT0
BLrdMlYvhbxk4r0tBRCRN9SCGtBKnqvdxxNUFjZhwz4V6ai17l7oDg/UOUZ4Xkgr
dL71qyJ5NjQouB4Fe8VAtJM9kds7J+TxEevIh5lrX2VmXVeKGlXrLVCJBw2uVFOS
RFnGQni+Pe9LUILwUsPi4jATmbhb+PFyRMM98klPvSXziCdLWva6nfh0L90uZsoB
YlHm2zfQvsJv3mcOnIypWhDCBXcqOr8awIvAZl68NK4dDSrh/DsDVS5wW6guQ1gn
6+ycfGJDK7emcJHU4SiV2anPPa7/AKNwI+KCrYpkbhhnmVdPz7Rs+lkiLSIiuanC
1RBlqC/OcGyp9G0NHPicdjYZKyIZx1balw/D5Jjzdj3AZUS5MMEBkQZU1L8FIQ/H
A/HJEtWa3p5xINR17II8rr6kAHxue1g4XdKEkNa8XDrlZX+2GUu3Mb/FIcYZNSig
2LH4ovGoiV1D9yUTLpOVJVPNGCouRO888S/qOha1m+jwF3C7K+S2PeE5bRDeYG3R
LWvP8urS1eAUXxCc444Wi2b7V+rgo5L+X/ZBP3QqTakXM8mvGL1CByxYfSUYzHqq
i3SFVXLS+RyC01P3eWV2Q6hLxCKMOpMn7T50zYnW58KKbJBPGtpRmW1sCYnhKZpn
02MEj0TZFKi6flLHIThTrIy5i9V9blHSUYCe0AKccpgBFT2jTnonlln9rfl6YB47
68RpepbDWJiySgLrrkbEE95SqJ0c+2DZ+pohXL2wraqkSQG2HF+s668ZZwZeQefM
lkwfu6KRQufJZHiy1ariT/4s3JFoOGNbZ9itNn+iI8fnFNTdoJQyyxLR70YdKJqO
5zWjoCswJP1+9t1F268beFTbLh+mjyYHI39l//Te+v4eoMc9Q/kuL8aW1Fso3XI+
m56vfCxBXFg/pjG978QscST7VHflKSqrSDLLarOSHjGzCYkaHT48OUFv6ii/+Kbt
OcVijKPrQb8/12iSFCYwQmmhf8l1C5uDeIDRY9YQUlXpnqdL79c1A3Vxs1sUoXT3
zKxG7ETVy+8RwTDvzHJnRBT2s8Sn7FRdBKN8/XUF1x0MSf8MvcADGTn1VaOfjSJA
ItvapROUW4hUpAGPCB4Fa2Aax8smibcQeLyNCER+whRcZjxN5omecSERTzRBRc1M
c5I0tkIJh+3TSxqIsr14DiaYtpNJUfYggtiSltQe3kCwhFDqm5FAPiKe8PorNwXI
1S/21UE0KAUerX1L6EaEZT1S7Pi8VZfht7Wm6tEp1aa3Z/aJIeMJPJke5S+yKOrW
4kdrrCdXvLv4WFGrn+xKvBTdfVelG5Jt9qivQQC9Pum9OLEKzujVMfJM6HztISw+
lx8B05qZRk3tkzg8vpIlY0QcvEvlAVI2ddpQFLQv0YHwla0ZGon6VilD2jPX1t/y
IRqQi8Dhv/XGE+TrX1nAHR/t24YVKQhJLjw3M05kh5PavKWscKRW7Ko2G6sGGpPn
Q5BeNIpizj3Sy1n2vffIu8BlFpsAWyyq1TRK5EJnvW9wxcl14K/CwggKlnlVdDwj
/jx+TJjwBDLhORBBklCTZLH86kRduG7wtCN4BUcQIXf/3ddBDvHobI4j71lg38kc
ghGM38BsnsgD+5X5+sN4PrIDhoLiTY2UagzJ/YlWqpbVw6+br7zPBMbRnXiASzTC
0/kQHSdiM5ab5H3RejKtuMklNIGLZu8fSV25e33SKjfN8jcDgZQFoxjzfp+d+wmA
I9jW+ir9enni1Lk2hG6/n130E8NXLHUtQCtVBPTes0cIgbhs2s7ePRp3ByFTDQLQ
Qr3wJsUd3eZHpj73jXkb3g0v715JCZHcbrdJaM9pZnbLU7GIXftXpPF2RLx14ZDY
NrsrYLIoRTKeqfJfD949i8BWIxH8NcaJlcCjkhdiHmUe4B2Rm2m2jNLCOxJU2EX6
kCmwXfYD79lzVU95gqESJ50ncIll4bq4dcEKLPT2302L3zZC7gH9QCZQeV6Q1jw5
0nuYdsOb0zxx+cukqRBcnT2o+OIIXl0hCWE2QYuy7Ir9AXpl4YUo6SHaATnc668B
Vdr1Zj1eSDI31i4T4T2rPof4jD+d02f5AXrnlTjw4psyyPk9gXifyOFLKH3Lad1H
11+YaCsxxqocLCD06r65hM2rtOu9VWF43gY+Hl2lDj16aIJYypeN+OpnSkmVTkpN
fHavy6nv4DVhCefBVRfTFiPVnrz5TfwwB0cjg70yrwu3QV9VxuTqb4O+sNSlHfw2
QWA9dcN7Hj3q25jYoagEU4mYWInqZhug0VFMTf+rK6Ra6xwYll2vxJjaTY45kF2l
P4ovlW49yGhzlPT1z7Qb+6U5p5hbj5UTt31IMIEDLnY+nCzFFbv9VB8LqI3TecIb
8BR5EY9NXbC47o4N2axEI0Wr4TlhS0RtjCiG99aAlf9ue3gLpDsSATfc2Hgf+znV
K3wcFb3E4guWcYRufsbcsxHnnDCSBTDiDrOBqSxYxmMVPnQ49DOxBesuwqdeROXh
HtsSGkkauHqbEYEgvh8yiCgg5c9sDaAMU58V5mhYC+fP3h910BMis75H0TwXu4Co
eJjyPsIjd1E/nAFKs4a8jffheSb1128JrdN/LxIj1DHaqC65nUVYvpkZCS0Zbc0H
Qqlmc9/EsXoOqXljUkn7Zh4ll8taYEVUWxMdICdpxWoE0cnKOOjqawJ6c361dUdd
f+WeJ4ggqVXMWuxabr24UH5O266aQbRo/E+cI0rNBUfLbdstOgMTTOybekxHDZ4W
F2SgkZhzYzH/831TGRstgSjR5lMZtWPKG3I+/0VP4ZhUb5wNcjWCdsez1Ucb1oqu
M1nT/LtRxBlO+6mWtueAxiJWDELQgWR73/2+qRBhzB5Pj8ATMWa/rlmhG0Tk9ZsJ
xkbOIsAMikbWCw1+1COs+aGQzljvG87z+DMH180HejlYKrg+6SmQBiIZUEgiZeAA
lPweMX4x3ntQYdcwM/+Tqpzwz51u74AZFWudLJ3r91L07bKoJJYjIhEeTmcFNN8q
gq1RJdan2miIqm3HgrYSmFYzR5F7vgA7LNwQBpI9jWBkCPr6xFXykhD4Cvc57DON
VReURpmykJ7dEEbTapOCXHMOo+XtBsXo9MzV/Kb5yKjdD8sXheUgGOrjfQ9HsUkw
0XVr84m7Pbhj0qS7v71jD67It6ASrTIY/xhvlhHo1HtZGljn37gjnZw2DuNYPgPU
IYbRj/Oqd/zEj2v2rDxghUTDe46bz8OOqQ5SZlzsgr64+Pc6SgreW75/TRQqpxT2
0voJsdz961LVe82UeRBIwTuJ3vTGEMKaqLnBbL4nnnhgAvBRmAnVSECka47IbioU
+gBv1x2d55hs5UuflGpcNNC3f6KAVhRicCyEJWrijfUMx5YXYFc023WYXbuZx3j6
2FBwRudxmtWfDbyqfbRL2f/R9yn+81PRFPVYIPemHvyHrF81mmi/TfNtNRo4nEvW
+i56QTZyj0Zbiu8YyULdhxccE/qiG3GYhfe2/okVCGSZi/5sb0+ntM7ABVP0YfNO
AvmytNbBwqDZd3iMm0Zvk0Emg/lmiVojyWvAw5Nq4n9rKhFOEpvyRDfE1hmS4Mdk
tnHAHTRAoNo2/vk4bg1qzHWNTLjHXNYY/bvIok7NAUoN/N3Cy3uxm2bsmKcl9uuB
E9JXc048W8AyK2gx2S0XUCdbm5mZdyLjIz7pPBWxQPVrWKEeeoqo/mxQSYqaK8UF
NxoJDgCa1e0QFp2ovn3pkklLmbdAt2/1SR5Y+rcpzi6IepkFK7yN7BVn3GqF1At2
iiAxlBeqSzllO21EUeKtJpWI8TVG4NanW6eeRt8cZPW8rsQj61Aw+rLNzSdiYTKT
eKB0xNbqGJWhULx/Oi6iRQKHqNbTkYaggO458bC7xtVZmJEy8nAJqGqmSO1c66VL
zOxbPyIIuupL6IQt1fmxo65t1i4PUwh/QhdZrbGDhAQf/gHz96yVzfGUrZGBZeNh
Esqwm0YD86YuTA7JHi6wJGlZ+rfQXHr2RI4Wwut7NG3Epz+T4F44LWHFgVUBiWXh
wtVPClasCoJXcZ/YQo5zXgHNoJzuSyWIAuUQlAMGaPeUHwv/y4bPshSHayK+LmCy
aqQb760epO4Yh59r79z+3GqdC7Zd8rHv5qna+JtHI95Qhw56TSntTwdtqW3art4N
MPbKHs0we43ji+L1wcWiYaSIMp/l/0qpkXgAHrRgWXR9sCPfX432n3wfsslCLVwM
Dgi0xILeNCeEfIgvLlLtRDb5hEhKBjWhatzi5jBve/EMwmPXUtc9DGvMAMfiE6yu
lkWyaR//3fFKkDutic5+UrF9oe2t5j6EjNBNYs0XkJajPAnZz1s1h47LKpbtb73i
8GRYJyisrMZ/II9ta9dD1s+L/LPZa8zLJnIWjtiYqAuuTAAjJM+Y2pge5gp0Q/QN
kpw9yewvtU1WvTQHdqMxrjIfeM1pzgBC7CK86J7E2UaqcDyLF5woQ3UmJnqE7cgc
gvR3wEFD8FxBnehp2HqrYSTrveb3Uj/gl2G5l26m/6yXqyh9RtC2wYc+3hTbX+uI
Qd+KAMpho0MMcbxq6ZLsJjE4fMn6/icGlCggnVGJBp7L+BUSrZE5077Iq8jwPb0k
2uZ5kyThVRP3mZltRCJFUWHRdyHfjccJ3PQw517z6bsoTC8GAbBWrynspfneyuNp
TlZz6hUJjSOLAZuv3M1dZgtl9GjkQzfOrwBP5IZGeWdqLU5Y688PDE8umHiqUbaE
xjijTeofbixCEruB6tD1dCDTfdpF095nYpiK795egZ+1UH7UG/jqQQZVxThNANcU
PeJDuJYZAlciVzMJVOvLd4xt2U9x9eQnvrZ1fXP6rMU4rmlV73B2xh545oIYABRq
AOSq3jxx9KvI2Uqf5EGAA1ycajmmrUCL+V1KFHYk8d+KzCMV/bkbZA51jAw8PXN6
uIqvpQg16NKrkN+D6LsgHqqiDSQMvt9nnWY+qKhOz1HKlk2jth16TOV3161Kip8p
xDRXpZdLR65CE6wfJXxq9Mm8wyEeGryEIDYbN86oOIOr1hJ0eV4h66Pbzt4VXWok
99AreHNVbMstKyK9unEJgX2d1xI1sXHt2ZsHfUhqHYsKw5DHxhsoKE0Feu5pEsWK
ZtXi2V4AcmIOrB7PW0sJtAboaY1kKPbYt1ZHpikQaOiS9x90/5CspPYxvZD+j/0K
5a4VrIVUztDH9Nnz36cx1ZC9HhwK/Itc7/GVnDJ4Cu00S2S45wAU6c+ysjF0wyjN
i3LNYoVmfUfTvbaOmU2sHxWBpppnCWr/PgW4OQUz4YCV30o491LRrHciIgknvQCg
pStlykvWrcK/dBHAH/DmPvvdktPQ1J/7PnJnqrGAPUXhog3dfnrKBOVrkoz1IpU9
wKaui8Q7ThfVsZMkxn0SxrWgGNni8TCw8ROtkbOEeQkXSsIvEuMBUGFV30EEObZD
h/82HykpZYxvYffMJO40LvqVBNoShCsa9CXMwOxmgt+UeoH+dUcKYxM8zkH/W1xV
izaYPGdJKikT0uZBw3/WRgfn4dmwpZ/Xu23UzsbVSvdP7CDwgMUIyyqVrATHxk5Z
TPk8zZHCNLMyQ3UfRjrBljzYro2FHp9HUU82XWHzrZoWvrhynHLyLm33w8c2lBwv
3uTwcZ5ihXZnpKBSr9j5jc7QmmFOatgJqIpS383Wng6/L+IPPLPmA32lMNsVeuPg
BY1Uym64sGSmloy/N6j8pCIc4/xztOI3pIoyHZUQ21AY+TYOqXY7FcwToknKMESh
uw7n9CdOovsujqavx7m/7m/SH26XfrGaer6igkTMdpo4JCdiSJ6cK6VDbUErLRxi
IzBW+w3WcQs0srW334y3H2rHn0omElJdTJn4ecpjfm8S/kA4SQLMmCIhmVQSxeG1
dV00xX7Bj49Cu40umxaEneiFI/82FNdWMFEH9+J7CbpV2MxX3+5CUw1hap5ND/gx
S2y5wUS9ecawm5uXZ8jOi+XFMueiZsS8m/bi321enVKlgDaEnGvdIh0cB626gQSh
p5vzlC4CTbn/5LQ3RdbcI1CouYQv3eCPWz+X0s24QtL7VUfvWTJwXbUmGlPSBof3
RTJXhsbKr69hHIGpTxSv6h7pgzm9n3NehkuQqAR5cs3kDuzMNgw9A7iQG+jFkGKd
geXb18ANBEkiRy6J+Qp93xAdG8IZrKbDczhO227Xqu1ierwzGzB9UdsAsb0gKrg2
w4FQfb53Qhc0gDXR8Gg3dC0x5xCwmPl7K9VZpniHtURcDLIrTj4DGpaCH5+KG+MF
2GlM7q/h0/b0ddpTmkZkOUEa6OjGWKLBTWJuPQaoikuAnFuZm3+ubSQOUuB46I5P
LCin3DxZdSHOE9XhPoEE4t5xNTGMub/aAvfxDQe/37lIQtatyVkzaJcvu3UdrGEV
6kpCA+RYPzj9d4F9f2jSJLvk8lNBwjNkMP6BuifuMlKOHQAt6gxL32In+pEOXlSj
amnf/U1wPtbpJxracU9QQcIkKVdogbUfquUGfloVFh+HLcr43moe4Tq0X6fb1Pgi
5dsb25qRBAdgxYCsP6P8BdwKvwr2CHWKy7gzNSpE2oVNZr2AtCSgq2HtW/+HyLJR
5zmvr6l7TBTbjHlYZiYgkKBBifxwB/mC9DOq/nf+u0q8esen14whDxmwqYUaY1uP
kDRzI3UChwN3Z8N9hI58X5mk11qQ903gGdE3LJ+2Ylk2L0ZBd+jMXIxxA5Bz9sne
iBQkd5h/L5jupvV+MEl5t5aVd83ACIejQwiSI53cfPfCVXWIYyz5ABUuaoAvzZ6M
80UnInrZlpLSa4DXIqYM8/qVQY/RbR/LPtOfz5w6HIDytOhhQlsOX3dmj473neUo
wxipFW/aTYT7Cms4baFHAajlHIfh5ZScFjQ2ymMuwBuJ1MH6/1EAd/V4+SCXTvh5
1bX44LpmQCKeblzQ3mMaRh8pYaeT+a7fynuoWIJzCtZKKKCNmcf5YvLwNgi6Jeyf
8otemHT4Krd6QG6wGlPHTlY/LFoalOVX/yPC9ggaNaHm3LJ2K2bhFh5fcuavFZTN
KNNmOuQ+ZlUz/NT0kpqvbY3B6AG2C+G4kV5RfiU2FvnnBLzrGbyA5krNrHPAY+4i
4mkgcXHI5yM9jXnmW5aQXjQIDsJJOwIQaURqqSFFFKan4/sgD5iC1C1zEVJnRFFd
bTicBQyFUKMQxDNC7KYkpQNXBOdsm+3NJGoGvfbldRi4pROCGyGBWgF7P9obgFPk
T7R1VN5mrKID700jwXCsHxsDCjDi6XblvrBXNTONa5KbZjKZUtq4ZZYLU/IKAdbI
xcwjgPYHpF6PVC3MpK39/J19sKzgifjNktjj6zGXeGBn3PbiJnjlCdkIOAfWcWAu
Nrz8VNrdj5GF8AUDwea6aO5NE83A5jWgMuy39TQUr7e26yEb8+8eJn+gIVq67Te7
X3hTiFF/0ClT844FYSEmZ6aGsT/fFlJKtR4u9W+5uc42xAkGhDu/5sL7bgYWra8R
9tVMNrDgSZI3aQHHUqs6Z8cpn19epl30HuYzrV+4lKppDGbq30DUUX0lHmAQvGV6
Gdtuq5lnV6jibw7TJXzrqJb24Hp0c91tB+D9Aiw3hs8jh7mEKKlfGAIxAg6zHZI7
ONPJDjjRmgo2ihrIkjVHTngtSrXjxnuxvbrEvgJxgLvGq+5NIPaCKlOUHGoIpgGA
yoAblw1rflRvUl90d5d0A6XL9AFb5JRnH+NtQDsTlreDFGnOS9WEeXVJYJ643zJ2
1ajmr23lp/uDIaExWZBtc8rBIeIBmzRFoTmTuECXXnv2FY3RqikH5agH6lqeFEe5
zrm3pjwM11E9E0hrfWr4+xIqkY6zQoX6P4qCVYIBwHwsEiiGbrlNBThAid3Y9RMG
qMGYyQYdLCjObjfwTX+s+6mFnoOVRaNQupWRNPvoQXNJCJNtyQsuwkNBbFMoHusx
sV8Q9MfeL1mswJcL4BYuhyqLiWJlCzkJbFUop9/6MmcI8YgwbeXTMA9/ugSLKeGG
jR4GuHFYDUY77oOszg74O3wklAFk2Lu4CGSSVkX+gKk+0cEN5ljaYo6kv/LDmqjn
IbaGOhQVwjxhKtoqmNubcQwX0SMfUHrmmqjB8Ia8KinKedAKAyt9YRqQ8Us7T6IE
5w+PUhqbwWy5dLXnqXdX69CDen2S+W4cDltUqfG43lafHL8iByB3d0s2662RVxzK
uLYPF3EC3I4RCsNov+UvAiF6wwhvzWDX6F3fueIZIEQD36KXsHzdeH5tGGIENIxm
qG/eLMgR9KCsz0M/DCDJDpuBq843DIUNacYp39T6Vc9mUdKavuhQloPWVqPjFu12
FjKSayfOLo8b4QnP47giqVWJE0hBDwF1Fm2RQkl9VqElDxALKlhlXRukgM2hCLr8
sppcjrmDq0slDP7Qmk/ONK5Uhkzm3/+OudhRUaJnX2yYL3Ow3q7Q7Ov5yEGUpC0g
btwBW+XIriKU+HJlvdXYDAAYG5ejWItLHkqrPiE9NUGKGmPsdHGSIk9mAapOiwgA
W6GlkbIw0HOOZSj799U/Hduxve2+hQ0Iis8dRu61F0kNsOi+zsAQAr+9rPh4AAo0
iI/7SyM8x1CDpEyDoAnQ6lFNxCLgrADaJ+z6baydlKXtMwL6j41j7fiM+ekoBTLh
O4vq7Qqo/Byl363Axs7GK7AHyUdF9oT+jwgvRvp9KhBnFf/6lzAGq//oXc7MOIfS
x7DLZR2DqpC/ws1+D9zbmcasDpjbYF1C8qrw8ygCD+WVR8njNLN2B5KYuxniXYYY
RPt13rtqCesDzbZx7FyQa6NpIIM5KgPChgCLs9QkANQg5TZMabEpZOfIFPV7Kv7G
hUACiQtc8MkvG0H97iuhaqBgH0vA2059LcaPeLq8u7OxiPG3Gb01Et9VQpiNn0sM
pdBQa+f4oCkYX9kCJSS1Bn8WtGwNpy5JWfUKhPB7ULhDg8GWvjNr86SQW8+A1/gU
3Azqewej+uGlm2KkeFgmxxIA33v9o4KWzO4GRJ/WNySjN7Q+2lPNksB6MlqIo0zJ
jn8sehrJwo7NEjwu4L1txsN2vayrX/mNfCcx6ByCdmUX/WqKpL9eyH2KizFD3TXy
D4/wvHouV1qOge02WZCIi6lAewP/Tn8VxXVZne4e/OzootIYQX8tMu9N7Jbpm1aJ
KaY4GbcvUvQ4Yff5ilKXIscTnyAacyWw1QXVVNGRGcsVwOtXZBA83dph+oXB/ukE
b+eEEMc9CZ4TdKcdKi0hg7+JXvCKOeW8gNA1qOqTM16PjPQlDVsPOWSb8hsC7SLw
GXCzIAC5aYH/aKBw2KBt88mwKAXGu7bfecyn5Dx8JMNPDj1QaJ0eVqDoC0GmHLtZ
cA15A7baSIKSso0HGKfvEq/8z+DcKQBTHqpI6PoV/NVkW+MjNWoUj9dS7YGaY7Be
ZYPu3uFSx1rQIrOkvF5g5nA+g4Va3apRpRBiyNSYBdXSOTOgJhuPUELDezD4vOvf
NbeO6qR5vXW3UaXnjJ4798oEMOVKb9KydyCOxI+xt2Amjkr1A0PnzAJ4O4GtnVyM
kH4NdbhIYYywI94g73nQG1YouQ3Dtos8SaSPx9rNvyoEH6svVL1BoMYe0Bm11yTR
N03Qc5q+SUVB8nAzuW5JLXmSFf1gl8vLef/l8Kg18PbRUN6sL4iwx3gCwXUfHn70
NOTt8tlXIcJlNKWotQ4AsF8ClDbBYOynxlWaNAC34CMKQkwUcNyubuDXL9yvNAk7
/YNufLywOHn6e8lcRqySo6GzoFnHZFiAxxGyfUNM8iV5cv9ACWHbgm2bCw/DgjzO
1IGeTbBnUdW9ZFuBn16/3xJMIyJwhXoNP2ZIUCJT4R454sA+pbX7HJ7LGLmJuXAl
2lRszYODsB8VagBIdHnXHDUcwFgsa27wzCbr2hD363d7cN2enAfql4gg9I+8AUhz
EWZl6G1/jPyT/USBb38gjRq71wXMRXwFKTzyFuBZ6Or9Qm+C9fRHdRdtMwhrb4xm
hB6VdSwG0cpZTS9Tu7TsqdsVgYs+0RokoDDaxG0ggXMVulaZ1E109gN01KdRxQw1
L8+8rZOt7Y9S2c7wjDul3BAlbl6PoZs8+IxiERhfRboCZNI5cfj8KMqwqllrqoSI
38tc3XPXyLYUTMMvuyfchiKN/DO6k8t1YYJE0zUdaBiYznnVTXmNxwoErgjeoswH
xwjRVjBL1O2IJsLhkcac/Px6e8BUcSXU3PYK44l4NgufPb1Vs2iXkzaU4ocV6Oj8
VusY8rXfCKeK4OZs/C8j9olOZSXqYmmwkvunYiM1iLS5hIP/DGOTbd5JS5N6ga1U
DUqaUAYxCUHQB6E3Wl0pmfYPiOClBrZuYfxgOYHTDlOfCq+exclvFKqPpYYBb6kh
EZ1hmNsYicDVYsQYelFr6/AMf2nxNR74Yg4gzZ0L0FvyjvCHrLtsJ2s/NOiS8bqh
moRBCvVSmJ2l7YGHuS8x/rzAI9kzMP1IwMLh7dg4LNAD5FPBLOYZ1wPSaxj7oQtg
uJ/nuK6OxxyllokxRTsfN4N2A74hTDPXtkzA3CA4N8dqftLO4jvq3U8mkpot6NJN
tAopx8CMSI/Ys4FW6lIpYD1l8CXubPToWjy93Q3MxzIiRfrV4JO3gRihHpOzkm44
JkTKWoVYhwureC9nbv3NXsCAerYczKz7xFL0uk8jw+Bz/FULs61DuNRj1zQpaVu1
EMKLDpxLT8L47VoUtu7njwybldrTFAuRMvhqAxsFDdbUXwLKPo3NSAADs2fqtUnm
stqQc2piwSN8k5IuYRcE94fhuQzU1VBrRBNoK5URRnA0f2Gywmlis/Wbu/LZFZi4
jCjqysR6Lc8E1wCOUQKuIStGbNgPYKzbeEhkHv6oZAO+E5H4yjNgEx0kCoM7bx0C
aRFdvvUGvLB24X94OdKNkCWDyHHJ6dtZNsZ+KDD/IorbxcdQuhsBIdlCh98syGOr
F5eFSz0mfKCtukfn2OGYW7c1vnX1xCs34I7eNXhOua7cah+PC05u3sGHnLR1OHPB
mULwZlkuS9jH2SknrK82DOXmySerTBfjs/68HSu1km+ODxqJATvcQGrp07x6xrKg
yyRsMk6PgEPyampmTP/wxetaznLve2fHTneLF6DV2AWew8hBK2RP1uLj4dRTSjXz
0aFWEqtWIsdjM2fT/azjzpI2LnqmEFUssApRcKIJTIQ7VLBGHs+vRJ0fPR2+lgBq
pubzndZIoMEdWRWhRGkqZJfqqDDVhWEC0sbwEil5hw7D45//c3w+fscPEXOGgbdU
nYcWeh2qGtALdwjGeU/hUDZSGC5TAdpWpzui/fHA05CtKmotQxbSFJuzjFj5A6sK
NEDd3LMvNNF8f3feIH7dmyIQ7Y+zCz1VmCix9uvHzsdkukNmiHVE5UpWDT1gX6Tt
biKYicrYAT1PyqZIRgYasfzZSCoM0LeQzv1UvHafbDMwKuhfKSRkiW4B5oXQy3Pt
rn+BiNnUKErRcYiDWL2aDT7K2QYDIUExxtKSxxMtIENz+EnUoWb+tD4MkGzSQXUJ
vdoS4UV0qbDR5V3ReQy/q8KgtefWoVHX+vT8MhfO/IxKkEvqmECCysj7LnaS0t75
gjO/V1MMQng0SCHFMS+pnW2t/NSz2FhqZeB7r9b/x+3ETwwrLN3qMAn0rJB0Wnox
blzVh8dZQ2R795e6zXu3iO7RkM+1vYaCMNoTetLc2ZVd98MZQ7Ad6JpAzbzhEm+8
zlf0IOSnZfk1j4tbZIkpIavo/xaPpoR1mbpq6u8YkgeNHT8PRaO1XNkHbeSDSD3y
wwYEPgsgzPfv3QdnVgLJ52Xt1Zj0aTPczFTGnxrpeNps1gE219uRkjSMKMQkjB0J
g1Z+NmhOZHLdFzFyOD9w87DGx6A4BwQAqPFHdA/6c4XXtaWMCmkd9nmJkmWdxU1a
dea2Z3ELj2fH189XnXF6NFdozISFwtNM9swNjGiBUEvIwCGuXqBvO6x27+Vkemu8
TStifIRLHOJ172QUu9MUdefWacYtrgbKiTO9lEQwdRkXXqJJNqFhJZ9nHHkHAMKb
9hefOMZR/xHnHXJbOww8ytMYZWojxbQ/7UkpqwvVm8moTrcUcPhJcBM1Q/3dg3bh
AWH+gPmY7/e9krZiCFbQ6dWvqF9NY06wkCF1cNdQCTu1pyK6XgIhSaJ7sn82zcun
RRySaXarNu2kJgMBt758T47bvCe9KfT2bS3yIhEfcSKdhSsLtDnO/1oJrlVlWRuJ
UhYZPr9EkBjBxTDyJ/9rRnMHJhXYNJYwazm5XqiMejQBiqsE92X+mAEBb0fBQ3je
mpwLyaQgGa5NRryPj9bSShv6hAq2x/ILYioB/sFHPPkLdKy3P88nbY16s4jpq3oc
GxEgKUVu/WZQi1wxJso+AG3hq2P7vzQXn8qwtGrO/HRlCUPqSl5bFehgg4IgBsfU
dkd8245kWhlKXT8UlEchYt9kzFOvrlRqD24ZyygrxldDOzhrV/aPA1D2v+q1DmdS
A4wFnbaoEd+lMukUqLxIFMH4OpvJ0MBpBfuspJCafjw1kaPxDDt05iIAG7sftY5v
W4RWi+93jHDAsoNYER4rKSxj4hwrWxOGaIpld2NBhUK1SRgXg25J2NVVUzLrCalJ
az5vbPGw8NA0cisBWdAYq7jLXTheAQz3A2TyojDsCe1BJfg7LXoKNc8+F1rk+W4m
NAwGty9MFP+DxTLl5MISlrglk2YbDFxjZqiOIWmmsvkYWiMQRtr96EILwriEV98b
iWnbRrlmNbLIrkPU4s9RP0AT25RtadNb4djMmHdG3pxRQNziUddKBSQW9BRMCMUm
FC8N3FvLe97aS6HLgoAPyvutF92SAM2iqm47PX9u3H34O9RyzsIwTTCWAT1RCgeV
3bUqP4D68aJsedKc52qdiXRH0bhGgn98nH947ElPlzy7PLPvglgI9QJMaxIA8Aop
bJdHUYqUJKkDSHluGGBWRjlWkaFWpWMvoXdf+fA0hHDiZhe1PJ9ci82MB3S4ewhE
6OETiF8Z0pEUdkpYjD9zGHqHHNe7oQRHKxmczhC9AqU39LeVv/nRweFfrUUr8j0z
D32SzmsM+29iQ4nye6QWVdCevLnv0WZm1rPFrr51WBRkgCKk/AgYjjZGOsyw/jtD
hRVTIj143DGiU5QSip9pCw8Qz8LYk8pLTwU4OcaCB3lviPUsmqrLl4oV9Qy6kYan
P0NrygDGwajG42VJJtDxNr6vMIeBuQJfEz/H7Ut7lVFTCUjvhsLyK6fcfsBgVAc9
d4AK0VMeUyOXcRjsQ3j+EUpm/Z/Uzntsw8VP1HQI5YCqfaQdaHV6IjIrN2b+tArk
6++43c4SY3gUvzGU8wV9vXPYRswqJLD8TlOV5DbmqxBUNExg6F2ssK7+1UR2v8sv
HC20GbqBfgE/0162RolXpM+AV6b/ATqMC0qxCKfQNmCsaSXVyR+lFZjarhn+8p79
SVqIPs9rlciZz8gVAG5wq/y/m2W2Wz6O0B6DpAzelUSPjOW6AbldEe9V6iyZ/Q94
E9WHIg6w0SzF4ZY7miMnu9ehAGkIFjUAo7hxlNLu5BXG6YWSDLFYxkz196PUNnCc
UX0DqV1WCrDN0uHgNtWiWE7eaGnJQ2wUI9vwyD+4wivfAzC9hYoqAEe/RkFm6Bvj
vBxfw65iMqL57Ez8YNVQeZOocicyy2ccJ8q8H2NeUpDErrz657VZPYlsHF3PwQPo
FSmmyyzh6aOQhzF+tg9Db+CV2xPopsNwfzsnltzTz4182Yo1e+6irB+CdKwhxn95
ZJ4kIJnXeydFndSqoxCr84SDFB5tFMpoSme2TStz/m025qHWCYTf6AcV7QQTSHtP
Q+j73X8waqJedw+bn3t/A0oZrd7ymJDhwnHdxTeWFo9sBmufmASL8vE2dAXUn65i
4lJ2+mZ/FD8fkNu5XBkyC1EqTuXfK4kKaRjEohz/5wsDBVUn24QVPGpoexxl3Q18
yNho4o4z+9UskYUTdcp861iUjX/TOw054UtyrLgmzNEp6NqaIHlx46y75rgMnVmb
7zLhSTFvXlYpBpctC6sKPuNh5iot+AiIEYTw4YcIU68Z4OvYlH4B5c38ht3vScOM
RTmwejm890hG5RyXuk4wDKcE0lOHyTg4o1iRq8LX5Xda51hDrBK+dwXX6ciZp3+H
papqy4og0BXLQCGKzKZlyQEV/dmp1JDreqwWGjKWL6SUhg4ajauJfVvwjo8J3zs7
GbE5GKVl5nG575NZuYAhqRilR3HDScNuvTeWVaG82KXorvwbqunky4Z0UaI3qBqx
OAs81oUJPR+SQWgrTMN9HqzcrcmN2GFtoJh8UQtCRLV9dUeWvF2/OfzY95olkC1m
zFGT6tMViOMPKO7Q5kIREa8Y8TMjOZ9OwHvQCd2y4svB3KTL5xN3gA5MsqYZxAHh
pfGVA+6wOrxEGFEyXLjzx930VrMB7WoJbvZJinnZWjhrwISSWH6saE/O+sLLzJvw
cWpNXBHgYf3Gj9iBnfpZsfiEpUDQK63WkVXQeqJX0JTaUG6/E/SFXBVCnCU7maKW
duD+kTXRStQFUNYffCow/JxSYpM1Cq0UYyNyUAzBAYK3ITQQ5wuZgph/j3z/z7vS
ThTLB0d2z7G6s/GJd+YWE8PpWaQgQtiqlYxXnSZZI2U3LAQXu5balPMCWp/6QTbe
SAlPv/r0AE8HvQ3Mn4i33RWJzz3t+hcnyXcYIgyRgF7wPWHd5Xx/HcggpZE0kV2U
obECkUdONSU/XaoJ+HC2XW0W1bC4EIsKAiJIl/L8YuM95ivZL/bmg+FI5zju9P0o
GbGvX/VFyl3ho2OKAqu28w0MXOi5627zj4iN4uJxNqFzmgPZ43o0MVsbuzkOlrta
KHJ9soc+zEB8vkBtQgK6SbJz/yqgT7DOMmomefja5RlY6IO2I0ULBXqtQah8XDgJ
UIPL2GFvhedv8Ae5Fg0PqMkZ17vgtEz/5Njy/veVUB2NASj1Q9L1RwsUeTeLxuhj
RTF1tpPFAIFzkW8D31kzV2hoZDy95yey7X0WjLB+TNGq929AQQfM25+/CTgGzVIF
ZKhqzCmGH0NsWjaY2/KWHEGucl9PYbYwwHBXGk8cJw7/lJNuJdFsZSPey84a1r2i
sQgIU0NoEsz6KQwjkbKTuTFu5p82EMGX1yOrLOJDdmAGM8BmO9D4lSxEhMDg0SVP
dN6BbLJmL09vBOSrAN9m/snynPN1nyvFP/mpoPn38uC/MN9/zeRobtELxtiyTBOz
DzB6P7BakaKp8G6nxlJ4qXqI6/VjCTZ3AjYSWrGijOnn+os3wXib4UkfF4DxCvO7
CWWEBep7oi1FYEiKv27wzrign2KSRy2mEHCHVnsWq+HwHR4iqAMRnyUoJRIdCGTs
+R9pBUWOUZ57/zKxiI8WIOEac8FeY0IxC+5EfW12UrY5Ce31D2/cxdjpYTgBxxct
V+CimonVkiyLvf8AzgEs/XEpmRYtMwBAjyJyBZraQMFnOSmoTJ8Dkq6IRFzRn74W
AT+GbxhJOBcPnLSF0mJO7vn5zjZPvBkfq5Tc7CR4dZnktO8z3a2zjRCewuQOvvvT
238hKqziHPb3uCFU/dlBYwDbKDPBYglQ7bbU1g9Ayl9LZ5oKmW1oZNB1lbzd7hvR
uD8ZIkkYnFm2FqYYZ1adMO/N1sIXHU5mRC+0kgYD2VeqvlLKZDjfDy1GDPtOuaPe
87coLoNAbKVBTitccSBkml7x+wDLv8cAI35Q3YuQBxHSKGD+zFLomzx8OMvRwb56
kn0PbmfsQUf2xGrA0xgTQ7NhmZ51lZQLoMVo4qHCR7+gFWHTJF9fMz7t2hBkBHGp
bwwTANiVWONUxWym5VbFrM9QpcTMnCfeUusY3cM825vauyZZ+RVqUmLinF4ALK/j
eRIIwklNp/YA1ogmHMEiYyiDjdkT3J4idVm1QsUF1F2+N091e3trzSNmun8NEPBC
vzot6GrBTULB45s1XiFsmC6fWfwpuXHhdoIUE7ax13Aj9LdqV159WUHGOP+5ginS
kfsdx/EVYT+X3XpD/F8TFY7N/EKmu4HmboHlKxC3V7sYJ23FRGQPqukVejSQJA20
zBn2LPXWF1yUo1Y1sllYR49VrE1VtfmoxAVh3onBSyTMm6sL5LxQmVof28AWZYOU
Awr5gQiLCrzsBvcI81CIs06hlkGzS1LaJjcIqOll/rfd7BiETBE3BDwGuOpRWYrl
tVxTUJmJlwI8bErIEpRmU78k0+oRmKQouXrd8Ogi+wypyRT9kuAWqZfoP9oXEpV7
ftryi2DU3lXfqVCRzP3BsqN9TquOuQcegqo3F0gGRtCOrYxjPHD+ocLmqF6UvtWl
uSYW21VG+JH3eZuIBKraPffwwL1bxxPrLOZtN/4zt4dyC96jWU1cymu7DxHPvSWX
Cdjoi3Ucp5vUcy41iOw+mMFq+LjWRWZEsPcJ9tvW4FWl0MOmtpb1a58aQEyAsnMI
lteNrqt7zZEu4+g+nJMn7MxAkzDJu40CWXj7X3MIix/0NI7PvguJPIRlKSWbwwWU
pVc+m4RH8FXvLQIPDnGuq3RL8mHQxJCW1mcEXrw9gtvMgG4je3gO7RoioayuXx9M
bQhPacBK9pCkD+xElR8EM77FVVUYE3v8IzTqqTjpnWQeRelqOhn2rx1MQxrZTjlb
/nnolCWG+9dkhzdr5sRicIkkJTK1r8MP04inlaz5VWwMEm8Fo/LwE99VJ8gJJ7nV
xfqUPTpqDMmn93KG9sXjF54l8mJ9KSmkqVSOH7COKCP/++D6SM11QXOxHajK0G5N
NWG3NHy+a0qzUV6KGKoTStK8hS9nmIVvDUrs8AZ5gHvQ1lqiYGM0DBgFeG78IB4v
qKN9mkq7LM1L+okWwI+dUAwkFcJnmf3jyqPuXv1RWxM8ptwtlYEAx8IH/cwEYAb4
OkjSmh5f9CBm5Pi8EJhMH2bgwVtSX7H5k37IqRUelHq2NSD7zNz1YPDPou5G9rt0
ddo0/WoTdnIeMubMrIIOnXfZyprWKhZvrevjCL0aZl2yb2ndo274x3KleA+c/tud
SwLahObTIqGeR+O0B3QFQKluUYKmeeVbFr1lLWh1K4yUNn4So5HiM17H23qIKSGl
mokYff1PbRQDE8vhRU+d019VoVJbS6b/dg1+O1zda8kNcQ4x8ishIimiaspGBqak
D5aG+lP2G5Iv4p3RlEum4lW+cJ3aUwW6RhNuR9JZ0nNOgZ/2EVRCL5XlN5I6aKha
jHDNgbrC2U9JnBdyEzE+RzUKwZtv+KMDbRVXNM0oTk7HJjeJZp+vi/w1RhawUKNh
cq0IZYWsGhclgbB3M9YerqZRsMJfYrRkTdIcSX9EU0Fk8vy4Tg9DiARDfwwnKEDj
DvOCM3Zkl/+1dtr/wuQpZFsdEBEMkEODMi11gSI83UfQoQBzKM6lfpDeZKw/KL1j
NxLcxcCQamX8RNPbfZneuEPiWs4oSnprO0aT0pv21i8wy3r5WWj1IvXqjh4dvIyW
MQ5TdAh95JMIa8bUk9ObZWNRiB1g6rynsnUNEMlmKsS9Bv1rNvxHZ5rqgLtG7Y4c
AC8vxnvh2uymoCMnGbg4O8mAxYO1hjfSi1JTB5rKF8a6WAG8RIeU25GG91+RqzpB
+e26DuCTcAjPMqeZPfnvA1rypm0TXmDMETUGsvD39+Uv4oguO1h1ooE9DPsuYcKF
V5ehYIb5sZvV+RS/JiB/1djgI1FdiyQix03v0E9jHN2ReFHcIl8wHx8C8jEN5iAa
Zz0lihsnFuYdi0dx95dvURTymK/ryBSLTzghtSyl9OnqG7PYbt9AhliXgJrKdQoi
8sXpoY/Kw4chqvGvdzMWO0Wik6/kRurYRMyaa5FsM8rgyfmow2HaZk2TorpdMyuJ
75/C7JBeprtS35ffyBehYel6zJMwYyw7IdGvlkv5ngN+9DGbIMS7zB9ibP8RH4HO
+w4q1ty1itHqStd9kRrChEAr+Z//whrVet3E6iWiNTh3xPLzRvdQQgl7GDrzKDMv
aSLJSUkoFQAo4qIHXwP/EuURZxJ3TSpFWnL7VPqVBsNEkCK6q+hCysYWVLzUoVeF
3dy9oNNbIWH2wJW3H0gQEVPVH8dV4Nwsi9RsbFKRxevNP9Im2oacOAsrHGjTRxd9
hnIhUw5XGwj2nrCmifv3KAMUlCftnhX1EgyeIW2BcN2w5i7s88ts81losAR7JTRL
/whShLtxWV8nh4bQ2nI0G08hxzADYDEyPHCky5R5Medj8ts7DKwaPCwwTO1MyCDc
EgiDYZcgJwYfDrKIck45mOc8jdWSXvtdNqEaApW++jLXEMb0gy9n5MIhDoBnItcy
BC/ZyXP25fKuFwfOtbLB/BSZRW9iWZjKP1pPeLNCKYaInEmmahiD53mp6qJ2O6eQ
fmurtebdysrQS/ZTNSQEfSvcKTdK7VM/NHcwI4nCKdiATk0KP/veDgG0tl3A2LzY
nxUWwmHEtBzp7eUw8HFaa5OAJiwypj6mfL4WJSkhBfyQzFtHT39/sI3DvCfE3ur6
Duna0gyupjDy4uN2PmXlgS0dXfbhrpOLHCL1oGCNnwJZBygT0GJapG13ho5ptqoA
qpBYeVlgAgROaXANkMMgGCXTo2JZNs5g9eYyXVifP2B1ncsg4COCdqJPkWoJPRO8
Buc1qqJN5GP4IBNW5xQ8aJ8gF8j2x58NE22gItdp+nHdE3eqRS8qZXURz0nR/MzA
3oRkd88ilAYzTEypvByGH6ze5IE2gs38eMb1t7bBrQjSy/6+sSR6tQ+N5QRiO5Hf
5VD8POP8avOUuhDB/byBai3eRoLoNp1Cn6xNoWJQHqnsc7Kdqeh1T3APcPYf/o2G
AiUkwRLowjmy7OYufUzhhLF0CYIp5er+toAjioSRSxr4+6Hd2a0fxdJdcZdElz4m
+l5d6YZFAOhRiP7mcBGQwTfaJRE1cglxNq5eoy8DnD+11l1pibnorN1PUm1bZwQs
R6/LeOfkSQbOMXX82LnykMXUlY1V+TTqAX7jbyeqsfIZznfDtMwL9YduaC3VdjBV
kRHeeDv2aHF3Ni4o+8giKG8nx9ZELo++wKF3Yfy8Ga2gm8J1yaQwXXnHE4jx50OY
SojyBEE4a6WG/w8Mln6gi+yI6iRaquou+MWnvgZUarrzuEajh5o+ERZ1UzpIWpPa
Hn2gR/sgir27KsC3NENFbbg7PoPIpXBb7zODYReq0amhJMjAQvPuS9vFilPNHWIu
C5ICzMGuEKD7Q0gpCxv87J6F9J5dBr2JL9mc/6jSdEuhpu+SHNcda9SRO5eWIQo2
tdxaEY6nlrQ/5USe+NLTZmhFMk5MQF7bSktFDHqafPVJP4fxsqskWHzK0J50AK0p
7eT1Ke3OGMabZfjwN+Z4bE2BWHg9YcPQx3WRyzO+2HrUogE86vj9r5rUk5dDy/Ed
HVeomE/ffQmL25SupwTNiYUh19vP3o8wtT7lfgH12EXIeko4lrp0zF9zEyYVGPAr
L2gDGrVOaA7Ujs6yBusPn5jbF3qjwnqJPAN+yL0CfO+bwUqUPumezxioeFgkeMLj
4gQobvon3IGgZr7WTtkp2Qcwh3djKklrxdmr9nNuW2eFhiZcv0m4T7C4YJemFaQB
MLdbt77s25uFRd8t9wsxT7Qi0sGwSciOvsw17sFfksQAOM+vQ4G9/AxFtk0k+n5h
NuTal7hzYRLS+J9g06pD+NwVisXHx47WVWMcNtspIusWwr/LfrTwSM55votUdQoO
1SRNAlc4yty07BNrUWtugUdaDeu9JnppaU7rW3+sReVAU3NK5P44AVv6jkBBh6Ab
hQb2mCmoQgEQKe7gZQ2wIYkS0tNH9nbUwT3gSpSSXRCzSwikrR1zqsTQgMqjgiNf
1qLwT9NE2bhcM26BsntfSg0v9h7WVRgSMSE8fBQPRuMbdCGQn1SBXVnh/RwzTI/n
7dRyV7RhBu9vNO5pbirLfw6wikdz53/JnsQLHPXJAgBJu7q7vr9Ci5F2u1I8iCSk
o1QGkofixDmVrzhJ7I1YWcBiurCqVWChy9eHxIcvNcoTEqE2ufixaas+5mz333w4
cy6gDMm0Z3dSPbkfQxFlVPCQPfCo/WfGkmpQBBlfyfJxOflgKeG8ZNVr9tlF/yUZ
jAAfElDxxpnT83KHZcg9fPweltIqZtIFD3KZ8PsySasHhn3tlFmVftmPxkF0Ze0b
zJNk3bsFiMw4gvYl1zdBryEdyzEVRGbtTKIuQn/VeFgxcAucmyaMWqWpdU4mexxY
WHrt2R6Ck7LcFEXie9zhKOkBLlfMAHfC+B7TjU6Ykjotue3Ae0jVXTU6/zqFTRiJ
V2IlyzNq7smDMSjFmRbi2nbKN6U0VNZV6C2+SDFphTXTnESvT9OhlOR/Jj5eX/8w
TYagGzqkDDVMwriWreB0VGmooJoR9Cyx2cUzmoo/C1GLoqz62V25b5QpfTxQ3Bq+
BGd4WwGo0wDiUFcG2ZElI03Hw201QadZw/1tQNMRAGw87lAKn5aaLolFgbDgC2jQ
w9eBsnn3ozQ90bvz/eJtMU+vAEU3WtE0fhljlYMA0VL+akuLKIldJ80iM1GQ0vcg
0zYHeRvWl7Th143SAGMJCYgD2yyRLGJKO3eHA1YzAf//zY2Z6VHqBmC3rr3jI3ph
u3YJJItt6oHTChF9/QnHAxcnd31K4XYCU0eOJJOCC32vT1nkGic9GlR1W1Vm7dKi
fMslQYtvFwNpHq3ejKh9Mfn7zAJ+bY+AGg83bhLOWHC7/+pOif6kNrVNlXcw50/f
iTzjvO2DwNiy4nvRSEtlDdi4Ky9CdDEnjltoqHp7+VOn781Gom6P82b8tDIbWGZz
eVmWsAj1wZZpGEEqcAy5jHdTXclWlFKNnU7B6GhgJVc7IlmcFae3WQ883l1M+HfZ
zgOXA3h1dsJq63I6LzWE+vGoco2/2PbvXwEDNBS98Sehm8gjUFoGRSH4VAPOvufw
n5gBjQyPcY+FGysnbnkdGkHy6OHzL/9n1y6AJ7dwLl7VKxx0N649zfjzQyqk5caJ
iSmIyd1p+kSpkBgg9JMKk5ucY0AuCt7jHrzFYuK0WJ9R4AA0VFozW/6Gz3yDEu4q
vf2D8d/N+aiDP08/0W6GDhvdNyjBS1B5OzJodoDtn32Ocyv00g9rPDrdM9DZxpIV
JKhpWo3xhDmNwgrZDltYVD+E7BiCns5pHecQLcHuVa1xsRnx+dJUyTbkM89e8kab
PEWXs/nq6Mn0wpKeXs5X5WhP94EWo221ILMIzZINJjv4xLFID7Jd6vW4o+oqd0Y1
Q8GXGAaJBgQxLCmmnlCYERMZEYQuYexLsR78eQab2fjrkOoV1oAfzMGxuQvYW/JT
aiXVJUfNsPDtHDa0ZnI3VX+nWWKAPAh2zXqFc00Yf6/5ZH0djZhCTTMENcLAXV6o
YI9YIeR3C7AzlIlK7Nwqn1GvUQmEN3jqyRZ9wNc8FKFRiIkg9KEqK74VgAphOWQC
bTfrT74Ekxjf0h8gM2qo9p+jcTBfmWcG3Hsmb++M0l8RRmfYPniirRow3rJiw9T6
/kBlq6Kp/VG0Rue7NEZySbrkcXiU712nzQdmLrxFN13EtbGya+iHVFidkzdY//nG
UXCXapduYPYlpQV3XHBKfaQz8Yg1q9fWc4vu+WouDMfzY6KhsLsxKR31JaT2Vrtm
s5MC3iFe7IK3JwP5SfkPl6exe9i06gTKw0kEDB1aBbtP6E/GVvLbbGs32r+lBJdJ
36Q2SUUB0SkBvG+WXkB4vc5X/H66zXW/f31ui/j81RM1Q9SsI41M+zNMY8CuFQt6
WOQW6shxhR4FumDIUesR6/OSfF63T3WmFDFuRCAl/DTN2e47z0qoyd1DHFubCmMt
3cODTTNftl5Sy8sRmhRZJOBgyUUQtUMcxL+A3nNmkSHvuXgKjaOtMKewVTl3mOX4
KwaEdSAboJ/Z84JJCjB6AyinmXtbpRzRi257qIKucTwsH3fQbSLcFJ8mHR6QXqgG
Xed/ZY+iU/6Ix8vciC8pvgxj/RBSRykRllZq30yVQkc6F7HeecVnBgN6u35yW6i0
M1ncP3gJudovfNYFQ/9mzJzIq/1BRaeypUS3iTbN3EA915APVUX2eNYOmDX0c5yd
rtvm3cBWCK9IxqkwlpQjsPC8ic5pISTOGJ/+kLXgJmWH1zbn8J/49RgkclwaiKUq
vVjs/ba9vltao2pYZazjK9emn6L6ffrjWsD4EaIyUTE+zVNLF/B6mqHymPdRDZ1k
Dj+SAu4n7PJZLVmpKC3+lOmj+1OlNJfPIyMy3Vmb1JN8wEOyU9DeLx3pwAbXG1O6
6MEdOQ2/yikmDLf3dCBcFnT5GjIEPBf8YOtbS/x8/1aqictrZ6DbdiwYZA3QQLXT
FBOymQNOv8LK0q9WZ82sYCud1drPRisvTnK3WEhg48nAI/ubW4XqVyATlgcuzfQR
GMG9N/tcVb+l0aRGuwfdhu1+hTx3TmaUpupL0+q1NN8N3+e5+2h23hQ70fU19TLD
x/D+udySwCsLlLlf1RFkScmD5hg8RFNNQfwsuHOxv5vqk3jpfmpzlC5ugTDxxP6o
W/gaU8DZR3udcbNaF1Rx5ja1ni2aB/tCoWwBJ7+HfNC09VypDehX0kQ27kJ6lr0l
SSs8D2pdu4X1N41MGuMY91aljWZUQEtnuxHxhTlr8XTvxsiYrhorOfJj7DoDSf+Y
t4+pWPWGzYhHSIapzX/Wr7xvcMjwoJEplEYrtOSSBfIh0Ld+OdDj3Y78yqRD3SfI
UpSb4/0uca+KR7S0assynz+7p5zXoreczKfjIG4KlvujhMEFNS8SXE9hBBoo/qtk
nCNDCk9eBouPl37xjsIWZpvFOm/zxLfU5LKluqUiJOdS4IkNLxfRsK3hsrxbdGZt
ZGXnmEmPHSg9DuGHJ40eWz/heJ4QUmgMvRwKFi33C1Y7FZxQ3vreoK8q3L+AES2j
9vXE2PXYR0fdYjGA0G6feebKwi/nLP3MZW2Ceriu+RDoUEjkfhjgdCPnBKMUpa+J
Wp4ofgOAnFeyxmgpNmN9lPqJBqiFV3yry/xinRaY2vClDQII7tp4bPDYiwVDYmHh
n9Ft6f97hBEmE2Wm3hcQN2BItqs7gFRLwY8OEbR2GSCFabfIfQgl0KDcOvhZUnTI
7r28zfQjNRIjttz9wdSF5rYjaoBduHj0aovdRoSngGKozd9iCuRRrBezl1pQ5W2H
iaBIQceht29EIUUy8/5lx5VKkQ2Sum34Qul2lulAUzIdf0HX1SWuIiVGw9/pVe6D
UeO+QzGRRS5WcX5ewLl2GSNPRJLqJMNKJDvx7hMNhPp7DYfZ0CJOu2oZLD8MG1Uh
2zFBDjtyynJLaix3GE7dvpIaHaiibGhrFipN7V4kaV6Voc9dPIQ8AY7V0Qid+h7u
faHwJYueHh/jIO1fn+tx3EXPKQwjeeORlaNPVeBi2sx7Yrf7bXA36/bcJUW7Vdyg
z/gqfEw9CO1CKodp3ymKOr9NtXl3Tkxg96nw+zyWK/+0/wx/IqRFx/HePW+ia9Gw
Ysjtu/HWLI2SE7I18B73H6/JBFJd3KqvjNMLWUnsFEQ0M/B5dHgLQq0LK0XznFTN
FTS8jQFFoS2EI3TdQ9gflxdJsyT7oScHbDahOUBcwSVGefMSplrxi1Wpk4sp0a43
hxqYxD/NO+ye3cPxW2SHLOu3ohiH3TA9f9tOtK4W6nJH+yF44gCD6B1Uhaox/CuO
6/8kAuiq++boqA/ieyylaOCYeCd0ynajKfDPyvZENcd743WZI7ISofPNFR+cCQE5
ebmu8nOhyzMd75aMPyaZh5e3ZL4Sq0AKZoLKM6c0rTMVob66WTDG5LVEx/KAflun
AfHN954OIDOzB3iU6gOSgAJvYNcpdNqNgoDKgwhqpm6MgSkivj1FRKyYsJld1rk4
v7DUjLRrptGTU0pcSPgFYFT2om9muDXHkBoQ3l32YeyA6N0mA/3TdLpEtC0RAvNg
xGO4sclIFV5VrZXbCksWyqEQMu+ve/Y4/wCHOsC0EUmWncRV+wBj6T48YwF4SlTH
Iwlly5YLetWP9FF4ADIy+m968hczg7DhQ5dMV5DKKnYM5aW751ALDVMq3/4tQydY
iHiQ5oZAETXaIP1Nt+cHATiQBF/KyOl2zOcIqoxuUXCxoTPfJMnb8ljg746Hr//L
kaPg0uSwn2iYkxVfCC/WkOBlHcdM8j3SoXkHkq6iCuxwVWzVp9hbeGq1PjlnCfvB
homAxhK3bvGEr9B8Jyb8oFJdsNGgpw6ajiNaNntH5YMGM6GRbf8R/nFToV9zO4G/
hkit2v1iCvrfP3WByA7qSzrKv8Tj9xbfpmF/XyojQYY7rUNCL33jhNKjauoI17pW
EQQxQAX66yqp3YyFE8tVj1Y8q+/reQYLMO/mNdI2wpFQcdhXrAJvVnA4UvMiEl5p
8zUXI2JSMzFHDhxm0zSStt7fVplwlPjFdsaLSSrFnaegCVfWJkheyU5JEHOKiAO8
ZP2qLQ+OGejrDyMPvXKf3E1UJYOf69u5MiDKzot5brZ8Kx6QUJ4t7QEENqgNhR+6
Q+tm9W1mhgb6RHHDsOCm6K6sk4Zqykrgy16PHE9Z/EBfMEikueK1O6a7K04nBRtn
7IloPtfuHcPgGwWyUB45oKp00WHzNLAPixP3QdQuG+/v+RWuzlCaJGYzXpmgYQYe
9w6R3O6RLKtM+vbz1ZmsxglUStn5LCZTVcz7lPSBBXnjWzLp4ZwjdwLfCDEPtBOd
AfNsOuNozQU8Hp7YLC4Tj44+peqr1mpdZWXeqdN1kyzIcieVOPWfsiY1I7psaG02
sPq7lnn27W93CPd1RefsHeynv+55FvTkd5CSQcuSfopxoj2nQabBmMIF4YxZYVwQ
eIjveg6594ujKTZBcTDesgffiEjbKhL7iW8W1I17NJTbvSjsIBXzGYR0V3wfkaf9
Ytt0a1ytSlovWsgL0G+AHkQ19QyVLtOoPqwhfvZbrjoKyB8MSvOQdIzQZgKfzQnP
l7m2hL4/qtR/EhWHpp0zIUxRBPf5f0GDNf6GB25KH0UrGf1CEMY29JrEd6+RQl92
+eCPALdTUebZYnWHlGtxDnccqo4Uivp9ZB5bS/Q5qT+Uyiy11gxfLwKIKR9Fh8BD
944pNWaQgdxWG+1+KbLpRsM6Bbh7NFWpOHM4vCEV8vR14S985NTkjStxACN5OEiA
Xf2msZB72smHduEuKDIENvO7FD7NrgK0qn7S5dfEUOwqygQPtaYqORbKJSobjHzd
pvnTlxni1t3XzDfR2k2jhqZkNd/ZUBCz15TD5dnYmbg76LbFofz/c5h9y0/M+hHt
3rKkw9rfqry/WTW2b4pfrTnn3e1/2xOLT3+VQJMn9dj4T8jHW6fl0Cm/2lNnSza1
T1pdzUthwFNMw/9Xjtgz792j2bDg1jehBwG7OQ5Rs47ctcTbHRDDasxxJQcUgE9m
BK9oMp549qKyiSkkAV8Pxg/RwsIsaxsuDZ8n80G/YRq2C0qlTfMDLH33x8WuR4Ne
894jF25ZWXr+sKCCwi6g09t2+HsyOIQcvxtNk0FcrlZqxkM7UwaXwizZUNisDlF9
55CDBz/IelzZ3NgnRLoIWO9M6DBRYAcWGqtGlsDglhEQXmvwYeO/1zvUXbyRWH2q
HJ2jNyUHmIXc1dgZpjzERvEc8b+VXai/Ey7VWYymuuNGtlfO3MFX+a0Sn1Z0aWXW
AFm0qH1L0bOdOwmAMdjsWy9020Prcd6szEgdpZsHGuZasww/lmayUK+ZR51X3FUx
DTJXgexcs2tZFjHbgRmVEen9CsX9gEFiR29t/5J/exNtRpIJ++RaEK0Kb7RrUgts
jFxGgdPjAx4PiPR1R85cLa3pZVsv7sncwzMtfkcC4j32vtPPuKwJSblfnPktMGU2
kcDZ4gIxzEXLz0u4mj63swWEwWyPqRThfVVvRtoMRgAi9HLSAsKg8LOfUF86wVm5
j2ytnoO325CxCv4QQlekuy9e6V4QK9f3XzHtCBmqd4nzvaOmht77xOMhM/Iqoa4X
5AVcyidzpSU/kqI+XvqNXruftXkad/50Svfc3455X0r+Pd46SlZLFK2NXHyyhVv3
mh6B/xp8oJ5THPoKSzgxvltGu/46fl9kwQdjn3FsWxKNEjvn1KWmfBJjE8IFBNG5
UPZU1Wwm2TgR2XoeLrEMcNW4mhNtpggl3WBybKUFPxfkLUdAcHNGeiw0mu/vOaQ9
m2uig9V3mRiYaXB9w4oJLJy7MAQfarcvrdXWYKCRAxAxRl/3XmWxtZNlkXgZPJZL
IDZOEUmhFTANwONSe2wKjlp2MRVgDxQK6gUqLiiWFH75d6mH7qO8KVibbx7VKlYo
Dga6dUVTLxkcP9z1KrkDOPiiCz2TchCXCg91JBxg4KkUW8zgG0TPL9QGCCzUepmF
tbNf2Ap0k0v/YgtGe7ZtDWi7NOe3xPJ7E9Y+5hbOA0mmtF4fo+Mru6Ip57xMR5k9
ASJ54swesKLVKGAA60rpC0My4H4GstmqA2Kw7o6ynsx2BURtTZyJpgByQFldqYaF
xKL8VdAifWsXx046HWBKQv7YxJ+o84wem7ndh9Do9VAq2QxUAwjuGT1TmnW8KyWm
NtqC+M5fj1+mvfpNzg0GOgceABHXKpT/xwnpCwnX4wLdAyUP0TtkKFj45H3N5/bl
8zpJa5hmEfSpceG/IPV7IAgDzC7e9SS5ZHmtRvC5wKWE8gPwa7P/Pg6SVxLDuIiN
nZD+KNQGxdCegVwYFdQwrgBkXJ6dor+PLknfGNT7EYh8bMzaW1EDVyK7i748JL4c
BIntQM8IpKUImYylNswYULv6BWmM+7PR9Fnt4wdFivTAP7KOOgDtPXx4fs77UlzZ
dDBAVDwsK28xMUdswXqcdn3HxBit3odEM/VzLiFkU2wMDOIkEolHSuxhHNDnJfMu
iDu54pEEtxFlPZ5mgNkpd1V33LZMm0JFrDSgOsEftGzksaBD9oGqe3sGPPZ8a8Td
LrMK4D7/j73cPtOYJ7GSYvJp/nAhG4WCMalBkhQfCmpOCK9tXF2/CyQckVBaXt33
AliMzeXyGl8r7g/NrJ3lcXeAPLdXcM8Hhg6uO053kzm8I9F+ljRxfBZBhzntGAh9
VB5pI7FxTJkHNjG5ms23/Kflk8NIIC2TSyB2WGfHdSfJqJetWp7mJZPvnGeObOVJ
rLQh55lG1OrlLHIo+fi91Adtr4ghzou+8Bfl5bbZ083BBhXsqOUcXcvo6nIF3LZ9
8jquW5HBhw5ZDAaiktlr70Mhudro3lkjy88IlaU9EpRfzCk9r7mbbe0rEZ4WaZ0Z
N2T1JwqGSEZcqtjNXt6x2MVdFsvG9mK12vCWm+P/Eo6aBsKGZs0NlVJuul1x2QEM
hvRSerjIRUpRHjvx/pQYcHcOx54waNcQPXhP5Uu+m7zLj9oN+qtQebVCOy/KjeQy
Lxi3Q2dnEt6o8GrKEOvCA+ZYw7qe5LMJdv6ipTm+pypU8lS0r3OfIhWyLltKS9YK
XbB0LYmHvSX8z9Onm6un6qn3kdIxXDuCIeWHoys58mS+RnKa34bIzcpM+sf2qCyB
+cIHDmHHt7nFwlXJQA5EP/SyJb7rl+rIR+IuFj5gOW8sju32aeZuwL+QsthnPEtg
GsKwh3ogILkJXrAzabnfoeP0dGjAaSz3tUTb1IjN69xnLHj4n+bRlToubJA94y1F
C+An0i4AvOw2c9LN6lC8on1bB9oBql80jz1DHvpwFQS+NX2izTJuqDZN9q2mj+7l
aaFL6u1ZJhjQb8gLLRh8/d7oyTvaaI2/5yBogwb/YO+yXutXZT/pDxyG4zkpR4MF
qf+qvpHQRjiomYHVzDJ/5UD2TKNK9fdd+rv6jNkicnt5dYFsjmHK9mdjxGWBpKbE
mvo3pR8yEum+h6ae3btneuG9k3W/m1r9SJUbyGEhB3mVsu4qPqOopriTd2/GlYwt
qGeLycxl3ne+y6gMjtDs4plIQldRzDoDHSitnoU1dJ7vb0flQNd5NXmWSdR5liiD
If8Jh5IxB6WhYIEK46+5nRKdYxjMm2ip+vMn+RZrh7dpeVDhFbAaWv5bIE+w3zod
tuM8NWA4Jwauhz6snvjHBzGNVFYABEmU6h4W7aA4daoTHY/vrxUuQ6yjqTX++VWE
y4aOxSafOskijWGXpncCbyQDJX6kwoTGFGztk/Y3NdSiFeM1/6w1DP16+9a/mFSC
rA2bnIhAPDV0k5DchiIEZ+OKzWBjFN6I0QeKLwxvv6tYl2a0JFhhNPOdgcaRKD5l
62P2c2VomWNdWorWrCudyg6eZrKhFDBWxJZmlec3JJnc+H75F0oLbAog0pw2y1E4
NwM0u5kgIExY3EYKo/khbqe8V1erSxJIAawqNiULjagu2OP4wnANy/tYmsHyvA7w
6qcMELf5Y/IJkvqDH89Iz8UTT/2FHPse99EnZ+xFMjEmq18zqpU/52xFIGntdJiJ
h+Y1/kvq/TA4FE9m51u1CKY4pzabeOYqwyw0Ge3+ors2DRBpGElBmXd0KF4sojhm
+MTHefwawX2kDE3Z3dr57zmgqVStv5VcOLuaOZuxxiPc8rW1VIrGOLQQtI6PDkCY
ZGMvA1YZmqtAWt25r6OTrCAz/rSgEugByuAEz4n5/ThZU3tIAdhE2LZItWn7lNb5
273/yDqy0NjvbnQIczgtg45Lc7Ix6or+zSt4FsDySj2cOONQTjDSGIk7TK5Z/Vco
nNaciVln3DDTmXv/WN9PQkPhU7vJltYuwWZmFzySR+V2DXjb5nxX9wExfg16ZLCD
ptxbwMlyXT3VJ4i98tXbmfnFtzwSe0k9YAIlV6RxEDshaWHY26x2yvD0f1pkA9qx
liABYmb2pdjF/HpbFU/1C6RfSKtf9IHGU3x/7n0OZmF0Tbmc7qkzOqux9vxOQAeb
8QUHX9Zd3PDh38ZKwVQp9snXFnpAOOcYmZFooeGfohJGiZ9ZospY4gnMqGUIVnby
5xWnTVeBchbrRko19r14sciDed2dff7utMXWt7uftjl8KsDcKtwFT7VtwoRnbY0P
qcsr22ttvbcIvdF/1gszWszfKEcpC+MIKx5cnzqtwvrmZZAfUFQPU7fIvnNXZBrS
5KNq1fWoVt9DWtwjzWApmU5+VH550LD57lQ2T9A6HTmCdQNEzZJUrFV73qiN4NZs
f5xcrRaDLHjWRqEg93kl2DdBqYBmbhrPoUsoXpEu4zwmW1AbxEvXvGka2nK3ULos
UMgGcpwx4mNutBlhu6u/FzMyT+T8Jj8u6P+5/tHQtxbe63C/H3XYC04QzKuWinOC
SOVDa11KZF6bNqKkf0025k7QwKzcBzATAMMleHOI9Y2PbnByGJyoIYrMQAHZ8PGV
7gmrrjXysesm3hE5Ns07PPpe44pklNU13P/FQJAtxDZtacwGl27m5zNm6sNxahBl
wbPDKnWECPJ5uxCQieCv1yU2bZYRRFxaBoCP4DX/p8yaOEYahd7VP8O6dBWhKwiP
jFLewXttc8xr9AkbiLfr5Elesnisyu9qYZ+h0lBpS8x1L7SbaMggzSg/8SrAH4JV
LvgnDP4qMam81F2HWmddCUj+pY05VkH4wOGJkT1zzPSmktvaCvfO84IVFm9Jl/g8
HGjsc1TphVNtJbmV2AcItRRuIkvrqR587xId+Kxr8pFHY83GP2l6N0HIAxwiJUwv
INRAsxk755J6PXRn+nIhoCluLFEFJ7e2CIrzOGz2COIkIRhU5vM4CeN+j7FTUjP4
7NaEk70aUBLxQ6voNS9dqNPAtU4dqwoYR+HdWkrmTg30pslcXnVeTOog727y/2x3
Fa3wa9vdlZS8E7EYiP8NL+h9fmQGEqQSUseB4/lfGoSnY34Jt5ARnkVoHkKeIDIX
dphQYaN1UNVw5hpfQsQzl8dRqCbQzCi1jsdoQQBR8+cHZq2MkTD5lzPy4m+DP2/l
f0FscP1C7cbggjlWCBVywC17mW3MJFu24SAqWc9bH56uaXscEWQ2szItOH/LwRjI
Da0q1rUW2sd8zSqmzKdkVu1t4pg5HxLWtgimBfrJqAuP1O0HZCsCfT+iYaAWcKHM
59nxcQhkSp+m+rWRpuVVFzVEWVDea7TS5/k77jvSWlUUTR6iZjsLgY+zcIK73EAw
6j0ZkPEsrstR9ScXaAmUc6ZxfdDWRpJCubRssD7+hWseY4lkGIzKiMqbUYgk0I5H
9x2BZ6GAGcLmVeP/gB3N+9x6UYJyB33+s38D9tRtAd84BoYBgGtO/3zfGt9lG8fp
y6GDx5uiYPTKVciPGUm+liYPtB2hZAU0L4VHB6q/SV3OHAKhlcP9yDoQL4G7qHpt
GPL0oDTP/KZ8eIL8x4yyE0t8jUnFr4P0vYVaSeLA4HUGSmp2Il9BCVRv76IQEQ8p
fOuB4VjZaj2PEqUnwXa4WxMg1Uw22FYXaZHc05qqxqcuLAKplXkdDJcBXjFwwfaA
mCAHeRQgrhoRN8IjQ7vminMcvWMWwudnCOekhqVMwaHd0DiQlt3rQMNDqXZEmxDq
KlIgJzXWDNtjuq9CXn4JOM4LIfDb4zI4pO7QVNfKXqXepg2bPXqecaum8jwmt9iz
LfCGhH6uf1aLnbwcp3RjUbxReeDq9ai+bovvU8hJLbiNWcuxtU2uz2zG8r2MfC+8
Xk4GYuKv3VcEJt5340bE0wu/qUZJ0Fw8N95xstFf3uMsOi+HoBRgo7k1LLO0GUfD
YyAHYUiO1XTI69n8CF0tw/zRaSi3c9z3u0MT6SuTEPmhd28+l1rtylJXCnNKj+nS
lUJsgQxC0OAaFaaSTv3bkh6G4wvedTxNWZmQFs6m2LLmo5obpvNVeNd/2Jzl5Mzl
pKkLie5TFkuM9ZlfvsGDyxgPy++FK7iI0b7pPWfSZajoKr1kNssQB56/n3qeyM5s
A6z+qQHJWctCzB23/kMqNh1UFnxwYk5y0DCKIIN/En+Vv5OstsX+zWviYKHazqId
hLJ4SwMWybQCcistUFJgS5hrqmL5EXocwlZtTb+NZ7x4ynvXSVdjwhn9/cbFO0sU
fPqlU+yL1zgLGcb7/RwSabTs5J78gKEMMNcWcbexYpc/B3cMKBKNl5UX2ofmiNc3
1Ju1dJ5r553A1Nf/0a267B+c7mN5VwYTKzaOBtFVvRGMCNZZvzCleq1ToOTISUc2
aNKKZ4BSS6fMfxfF4pqqgIKVgdlPCRMNbds1foOMGPz4+f7D+JC+k8OeTOP/tOIi
AyGzMkjlqRlSVCqMiRAegZs4ebAO5FWgBsa+zdeLCw8yXPwOsXBf9CjZyqW6MmT3
9UEHCXHtdKdALC5Wtd6KLqcyPxVf0+7weYck7vFyaWmWuEmM2gzLZtFyhOo1RTS3
LE7Dwg6iElb3LJJ6vvHDqkfk9g3WPKtWsoEMA1f0F1aUuEUCzT1WB/az6v6nYooo
LtJkoDmYYYoKw5QrkYdmccKOTwsMDUV8LVBV0JbugvAB4sLgOqUgE9TmgEdGPvKm
fMvjl8AlzKsETtRf9W0N0iAWiOD2jxtMRPuKtrxoKqN+t5BaF5zTkN/uUA2vxCJ+
jrqHMy7BEWDc3YIesSZm21aQSXIhdzDlm2p3e66AP3stscyu2PVFqVvLnIGDTJ4L
/ganZllGJO+0cRCJ/V5Vshh570xNDLi626j+5YgvCq+dHR9W8PKoRaSVBw/qqnzY
8Nlg/mqygMFddUvdji98bh63TVt/ejla+swIJWyFWgexofqY0kxSvxs5SNPu1Sg+
6N+dayG4Ret4vdvYI8HPIJ18CDQ6LS6GmGq6sM1oK9W0uDewF3rPP6hLoTsk2z9+
SuCQRCw4QK4TORAwwoy10+FyAytf5lpR1/THSX28PIB2AEFfz22/QWergF9xCbo+
R/YpXpZgrk6OhauesL0jXXKSYfSyXeIKyJAwZXI8YFaSBv0Pb/GLSPrW61r0ADcA
iKZ0iqPW70ImH4ugXxHaaMKYRDgYVkoRAkU7gNt5vTuBym21cNyEOOw+mL2atHv0
ekmUeSkXUz1NV8Ql44IdR2J1hRmRsQRLgTagiSBwHPNlKOGr+v/Q2aEu5Db37EuA
hmTVS7tTa+0khic0ueUI3vW/ypRy90aw8g0mmfbT8yOJz1Gj2/MiVBkYHxas4Wah
cgBNt6ffrNEAX46e8ZCXaTr4C7BvpPnsePDoJN1sPsGXMCvcrT6MSnP2pf1bAv54
LamgqYrTm9l+D7TLLIfNGdUhIWeGrWa2gKU1iboIRCTwo9pc6sg8TMhxCl4ji5Rv
nmZD03wQBQ+owuoPNPcHUXXN4PoUl8mCTrkzaGjW/rSZ+mDTnTRH7pIefJdZxNsZ
DLJ5e3RU00mzwgL8HhKMVTBeyaZHwzuDKtZobJ/BofuNHKz2xCavwBTpz1FuRGhP
1lOx0GRmUQateVsVNvIzn8XW974oz6AItKj1d8u4ex0FZ/x5wLKp9x4KpQbNSzIM
Q/kCs8MhuMJBpnU4eStOvc9GNPQlcJKAn2wCl6IgaDKIlm5j36kfL9yBQtsenWC/
spKtSDsd/jFRu24AsEM3yi3NxRWqCRBSTrA8h+mJ4PRYPEPhRy0F+KV5okOLvpwV
2Meyt11jXhyIV/t8BmHU4IKtzUPUMzUBKdN4CDW/Twm/LJiV4cHLsR4k8uvVq2I0
GsSRj4V06y7VkXiKvSDUgg/2KzuZOCKGXa9FqQjV0Luem81OgZ0Jq0vrPEDA1pOp
/zTUxWTe1ICOGjD4P3WT+f/K6VhX+bQz13yDodwma+VQcUfTQWd/twv6OljsSqCs
2pA4UJXD0CljZnZyQBW2fKLhQqsVd4Pa6hNP7RuCfrYKKTP9zMnHGUW73sTM6LdZ
15dQ/96kM3wJBkxkqFG0yrpvEqZLQ22IH9kUnzL0e+TfS4MCl+cPCAA7xOO/IHYr
eAHSRJ89ANReRf/tFTGU5gts0Gr244TW6U303UsFOClvIMvl6CVLlylKBPlvHLrw
zN5VvL+wqAISQHGD4uWPLeZ4X4a9dfEy1/C2BYMgn4m0uawXndlu0Bj6C+xdbNuE
SmKaqU/ct1k3aY0Rr7DdZYBEXMtKecyqfphW2GaBHwdxxaiYLGnCWWTeB/2Y4+Nr
yoplaaMKSuNmJrm3Ud5p4+CVvISqgTlVEsboKATuczGzwAg1uafxgEzyZpXlnGfQ
LqxfI/n9NNWhGnPYK2PU+4jU3Dxb2i35lPoSsTWhqL8PGYjBGM2kMEsukzwJHP0t
swGzbMNKpdt0UfC4Fk609N4glq9xtG1gXgkbBCb4GShnRciiO44ScL64cpQNpM49
bsodMiAsH2H21mZos9uz4RCzhVflgkiV8tejM2UoxAwkcdrld07BCctGBM5/3eCh
dNGjhJMuM21STv+QV1GMTknGMLr+3YmBI5kJgQVWPcFXy5A43jtj1c/HHIrY9r69
HzFkzDimYT1icCxSWhaxSsR5iKw30fuK+++rsQ7eU/LgmafbAqSQ7ZTnGPwUZsxV
GdA8c4HwUXJEakATMKS3Zz5+cHn9I6jSashW2RLp5OT/Zts5EtGUI3qxIvVTXp+y
rjeoHvHSKq5mcRf8n/x+0eduB6/+nR+3CHcj5xzrEcVIEk3OC5gjUSmYbgTJHlzd
IutxlbwYRHJ2U32hLE3AS2HXHAbaOuNYWk8q7KN5TBM15Wbx2w3S8lrMkQ5SOvQO
uWiwusRmxOy0sgogqSIQNCgtxIrSn75FtDs/09iOz1+p4/OkHMKH796DFf1fvZjT
xkvLgdTfIGVLCcjwaJWGv5KcKpI452I7fv06hG2OUoUPyIee1U72yhGEdQubo8qP
5otZncxd1rr/yj5Vh9Wa/BCK530nlJG40zSH4/r/EXnapBtRLW0Mn5n5YyOZABWA
k+nWQtj7J18gKg5EYZ+Qz6B7PXjOL1p5tw5ATjUEvbbq8xYmOr/rtFGA/8ygYBoL
IymnI4eCyKKxcqqx4pPmG3ozA+D97PYCaqqFST0nwREi6S2WMmUVFCeiAEwnNrDH
I+Fcu0n8joyX8uBrfbiw12Fx/FA8s87JB9qlpo34F4/AWhkv4n2n8WChp7G8AJox
x3cOKJB0jYRisR59jdlhSm/D/x6R0qB+l0eIy9S882cL1B4Dy+qZAKAuCfo+WCrM
4tt5oEaH7CLckK0tFq1nd6D2h6Hz5Td0g70JOnzSHV+AI9sA0y4yy11Bgc65IGXg
pX0PDmcsndS6JE+oJQI9cHQRiiwF7Z1Ak3An8By7/qTpqOH+nOqCwb3uT0cib/ZD
QcvoBahTSzrvOpI27mHenjAt+yl+iBX5fJqABj7+z5PFEJjsNR95WSSngQqEwi37
yjMJSbmuNTsqBnMWteqp7jeqSTqZsY0CeMBWMo4DcnlC548ecM3VUnQLKdFiEpXA
7hMAc4vbqQSgKlXnLK21Uvopz/Oom45ZjJgVGTkAqUcN6Ir2+PAffOwXSAAtVpP8
avnoWRqKb9UhQ+EKhAOu/nJssIepf0hVwgoeJU2Rc77ucslNYnbMYS6MqFsy60lZ
yoxOfbNfQSxfM/7fDN5W+6XVhX4W+hX2x6yWEoquWNylFMEuuezXRollxorbLJtY
N/jb8D8e6G59eLThKRW3yD00JG+85lyjvreWBeb23HngjoDdQ564flfYS6SKuBB6
usIAOZA66mMzV+2jIpr05F85ylBrDlVbkPS/AtZuSyEKUI03gsGCpMUC5lPIhdA+
TF3nN2f+FlNfAzc0ZvU4orJ6P4kfZuBJZa6nE6B3XMqujtwGWi4cdGsHhIbdf+k7
4uKEq9lVg7GVrDJRKGpp3i8oRGmW95uArouo8r7LgjyX/ylu+6WKd/C9M7P4Epcx
3kUDfPVDKyrlvTWxgbiAkdi5FuRq2WkOXGUOOm8Df2QqI036Ra1jTkTdejjzpGuL
lBXI5d+LB9J1FeAsZjwcxArzPbto920gxnR+iRj9C8firhaogfEkqXJfXjwllE3s
LmYUDIDrwoxhnhh2inX61OTest3dpHy1/anwKcvKjfCYFqSuJs6Xq1IbHS4Xw8e2
C/bSF5Hk2COpQ1BVi/0YM9RVOjOR8ppoo+IDBbHMQtCI/+T5qljuxnemqKh3zSQ0
OT9g88uIp4sXEoIHeZ787huSZaNbsTvVz7XVnSyVPwUd/SHUjVJ7YO7+sNpnhbsk
M9s39Xz4NBK+fGO7MprEzQqICCl+fLuEd+8JZnDEU3BcfIr2lv/TjD6Pb8/NgUzx
7wX4UsH32oOBBdZiR+1ScTCX34Yz2ULKJKRjuysvtu58NksxoGNb8HW4yhEUcSDG
qUR9Jmg/YO5lidqMEMVWZFrfGnEFXUW0Djj4IqksmNGV7zcGA/EUwlTO1vnOPtlK
RBCEcIAmxFAMNFRHbzsrF4g0mt+AAffgBOqoJ1CE/RFde54YEaPlWAe3MVRAs+WS
Dt/nrawUP1T9mMl2upxB/6nG0ZtOxdcmfFuS51IqlNlQpMJYM+DP8A1FxKdT6Hb9
tnsfl5PuApmpH8S9X+w9WYASzmnRmhjft4N0JQtIf+sXHSZnOXS3Xb/14asKTHxl
m+5g6MYS4l+AGT+FMW75vm7yYGVqU2vJQ7+0zQXOopymIAYRDOfoZlXrZaIYyyg8
Pv5w6a2QTKLMfqlejD+nrifpxM0VVqYXUfcjwdLGzWcHxW+YSFNQCfhSmoxNY332
tb1jBtfPg2BmP5lpEn7TcW0nCFXuII65sposSH5Y2OMfaFrezMRREW2EiuSHOTst
78IPl9ZEvIT7QV0CMPj1rSYZXaEs27kYdhHKxt2X1h1xxNyTx4DzRAWfh3/HQ9/Q
HdM719eCDRE3PYs/vW7yr6yyMWOYLHIhMELDdPkcYohy8CaCe56uzPz9U6TAg1ys
X6mVOqRvpc4ydXEvUeCWiTLWo3yRRCvAofAG8XO+17bgbot8tXic4MdhQL9Z26bk
6XXKbjfT/cWGO873ErtXaekvNVtOzbcXx1aCAYn0ZARn/zPbcZYm04FNbp8bWYE1
UDGqV7zpnHEAgwXVtiLLFjFmEvSCwKllR0HCMWSEFkS6G/kF3dgBh6XKyacjhcPx
kHNOFT4mlchUTmdFapNrhuQOK+z1Jx8w5CxU1SOPr2JGT4tLlwfbsLqe5WCRm4t0
Svj1vA2SuGFAvMKraU6HPl0meJQ9LRvEssICavg5kyqLbZJKkVUOBGCLFbipZH3h
FtPdVxN4fuUr34yLXUHIuW1y7NL2jd0od3pFxa42zjbSYzmfngyE0yPzrPQ9s5qy
zP6vo4k78GUG5uClCc8+STw7l2yHxc6ph70W0QkCeyExgpc7YoOQgw2T1hMJsdkD
Kio1oRlODNQFr9+m1MtxzioReBFGMR7+MUB0rHCnRgR/QYH59KHzn+fL+2FZiVF/
PBZSuyFYsQ87UtZDQXkTMZgEaey2g9bXgPE40OYZ2krLTuNByuBGMVucugbxs3Df
z3yr4rNOx9ad75dvRTr9XJqBLxcyNQb1CP3E4W1VJCRb45MwHT+sJhi1dwIa5ygg
7+0utMS1TNTWan5u7ftlzTkC7kL0o6H/OB7agYRixkc/5YmjPCXITL/Edsw1AL1q
2sH+KErb+vjSNmdCGV34R1NOk6k+Fx8QqYeQXwN3dckXWfLYg/JWFnTCbaQ01rfx
HBGevnwD8N+j89kFyIVTaujK89g3Wwjl2Ljdz9cNcFWyHultJFSyAxZ+Xxa6gFQw
rQW7817JYT3gjUWyscVdjAxthc7FKEetykOgp6GLPt6nDqKkzFCnR1W1QnHvdEQ4
mqosMpU11ITWjGovj0cxgTtal01TprZk+0Qsd2YQcIDJC6EXLvJWo8uwe+u8N6V3
1B6hFnFeOBE+4Ef0P3LCtCWL9/nGVn6op6MiP41WGOHCtNDZZCaZw+zdi1b1SOsZ
XM23DxyarW8EwQ86FoiR3WiEI69EUMWIUWem06pLTEzrS1OPATRvN7tjQrZjJgFN
D6kqKnXaZ9ryixMwibU1gcURfXt3ZzwaBmrz4N16y56eFwwY/h+0lRWRKPQCMapN
mw8M5/SDDodCC2Bzhp5ZynqfjUdcrQO407LAMpdCosMJKaTzBuUvO0fLdAzVEAzp
E/YkfAomanyOvEiTJFR9JP1LQA8bNSKLd53A2tgGTuCSN6AIyL/wHHJ4jk0FG5Rf
gQyiBRA2/Bjd4QTrVPIjzDGpvzWufRlYJNPajMmEpcN5hodlKUNCwsI2HrqGTsMk
y1IytYYHIlN72aTVjNAMMg+jEvC7AW8MKudWBbCvJzL58mAOCyfZRhXlKJ5/c3GI
aQbvKh6H/KwaoSz0/du7mlSSWxPzBflT7hgSKztk8odr1CLM1DIMGsZ2mB55M62J
KjbiOAFzi6PpQew7r18MgWsPi78unk3K5V8ZmVuzq++nOWts/DeEo5yxvYrBXYoz
DCvhxNfDe05Jgs23rJ1oSf6E2vQs68E2lIiQwCuX0X5eFNtiCsyJV794xH3iHxyS
xAKH3dlVrdbI/KhCY1m0zFmPukdSxT9yoi++MxTB/Ps/Tt75h16HU7nUlNNBs6PE
M50GHVTEwYfRPj3hsdhB4ngG7g28r0d0pgb+jWh5Ifkz3KfVQxaD/mi6PEozmR7c
NkzWaRnso662P55IFnfaV17kI1DVLbpdTC8/WKERuCJfvSLzoIwZFHU1Hd0PAFVL
/lKhMwomH3Zw8ZGYV1YMEnTpd1U3rtUBhQKLqDtrfw8ZvPweI4HbXDBoK9SgNckk
KJuq34cY5dOhhGjyfHzAMq4sqSPx44RQR4k+Kheu5MMKaXc+gzOJ8CCMMXKaQ7Yr
ykgp7Ew1tb0S/yCWL1omzS0GJiXZOA21HOZPBpn/K0o3tchdnd8pCG6zR8jZ3glu
SpOcIRRnPfNq8jb8LWZ1qjl7qos0mikssnoAREPMM42R7sg4fPy/sCzNjQHobHiZ
EobIYpuwuw4HRtpGk7UwNdDymq9X8aIFNAUuVwZX9wqY1iJoH24MBAhv+G9yTZ+0
zy0Unc6C36Q20PHmlDrbyuZhmyo+Q2+j8NgvKlWwKgwuBvAoyQ49ziVKxhDm3s2x
+TQUrKScmGnCtOp0LnFBrlTjASZne+I2ARn8ZrCgU2r9yIA3i2kzWXpspMId8MdC
TInxX9gHG+O3Je4RHZ/WnZVc04e0r812wLmDmBcYWSB+8LdWdW+dqw74k4vevmVM
FWGxuMR7T3pR1h8W7n2vErIludIGpwx7JG+QBiytAqgCjCr1uMJoxOhCXReXOWrk
+uOz3bzxHQmvromvIHlFUQ/lUUeS9ByDWHM0FNTOZaT5Wfb4d0lb9m2C/aWNFj8j
VMe4GH5pGDWHF/UhK3DaZiXPwRDZWRMAcKqjB5AUNvnVoj4+n2IBvjhgQJhpmq+2
GLz+fOOq9p1G9PK8Q7CBQxuWmWxfdWjwvvZZMn5yg2/GclkQ9eOmf82uo4Np9x3M
hon1Ra1bYgzdcVwU6F6aqpu9i+V8Q2nq6XHIu2YOCqXfJA4Ikm9H70X1pOlU1fqb
wjXG2m/tkcAcNM35nF8InkyuWpiyXSN3yOar99Vw0Qo1tQXiOaIVrP2aQKplrbMr
lb827D2ScD6zA631LjWaoVnDORUvO89erqTnTDRqwF7a1uySBOGib6WQ7BMLvvOE
ngcchbqHneAPebhZGlFf1Z+tWuH8TfG0JQoTmdAjOgPGw69b5Vp3V1SASmVu/DHm
H5BwFEdeYlapmX9FzuIjuRBdVnBHtLDYrDBkdIHbSeWX/RueXE32Ix5Qhy0y9znZ
JY9jUS5BW5yA5/sUSpmHw34je+CjBgMq4L6p0GLPET0fo90FWpc064W0vY3Y2ihW
UuLFUjSP9hLl1TSUsd3m1LBjc1irEpaOrrHAtiZdm2u4O4x3CHXBVij159uNg6nP
3I0tsXhCv4eeuW7PI5aYGPGGOZujazkGkF9XZ1LDu2iuUhelNlDrkKo6QD2Z2GbZ
4tkjAOrvulapu8OOT55FaYcnWok7mIo5cSeSG3NX6PHLvei7fIw/hzZ1eBtOL9tw
RX1pqNfict9srGpoPTK3PS4/g2GRp2CJ98lNHCEHbcaiDz9BBd9/yT6BFrr5GZAM
MKrUWH8KU39IPdM3g0sDykRbFS9CVrxreQm25OxYalhAdme+uw+JEEDKDFot/9iK
d6sk5Onteo4eGovLfDC7oZyHCn1ebHAuU2q2QJ+bwTIvnv1qSkX/DHmQ7WPCDm7Q
j+CM5KqX5bphHOiXphM8v25F67H4D8BNgviUwk3Yj9shg11n/WW1N202bkKR8GHs
jaItm3+rlPPd5mh4ItpM42cOGyhNOUQMuIsf8uSz/0WpIoDkEz4VbCTkSgamvsMW
5gyoq6cAAGtvJgmD7ljwzN2txEFeMdG2w6+Q/PMGsziHw6OabLmTD987kG1lEapu
v3HMO/VyDEMTfxR/htZkaOKwynZ3pKKi+mPgGXB9ha6rMLKo1emF/OldvvnmrA2X
i/m8NyRmYAU4ydvQ0jB5viVxsHzX+17o2V8E20OGHJkpFVe9laS1HlyJVtrkYOJg
j2VMukXOU2gQwPZvOcdxUhYRbHF0ilpGH93V6jt70hPVF5cbdWXFkRlwS/Umahko
1PjhRMYCbneVcyNWi61uAAfQ9ZIO8WQbIsiXA7yvlk97yOqp2ilPVQmfzY5njoSh
CnZkp6KNhZrzNzcz0mIYMOTz1uYCFDEaJZjDqwN35lr+xHjK2lHlgvJBugdoH5F+
dWOukW7VV8ebwsnlapiUdjrFoXwGS11gu0miu1Vlwe/TUM0HQnsYVHu9BSgAzBK2
zHFIEYMXNPpY1j/TlfKJora/0CrFAz0QNLHgB3kVL7czpnfcoEt9w3Wuq57ic4QI
+s/uika+dBNKNPD4KJ/z/iU8U23mIPb4Chp/kCVizIOuVzyQ38KeIorQvn0X1yY8
L4WgtN1etEzAWpLo5gL2MzgkQmUU/bg3b861i/pIhdV8xHWSZLNHS2uD+jBVTCZ7
AiwLnVOjOTBqSci3ZaDG/u33URH278rQX7fYvEPsB80f2XyUFneSTR2cLa+BprAB
OpFyezxR2PSgxuCVqXNF/ekZYnIKkEOQ5P7IB5VDxWQIx8z1Eolll2+GPdsADAsW
DZoX+v6VmaTgeDQ/grT68lUp+3t5om76pB1JRsFc2xYpaew2KE86+P4wZ0syLVbw
+5hDePG30+0EbBcXhNCDOOstaBt1aP+HZHpsKYMM0g3g/OSNxJsY6n1OT2+hyXGQ
BMZp6KAZMBIwNINmtNXliBCXSMjZ3tMWla1XHqtcnbti0w1APzXxrxa19gLZaPw1
sSKQCMC4Jf1nTnexLRnqQA4TE8I7KZQ8oLzrM0ZMkMwKEU6bIaWdZ1iMnUaKx+in
HO8EkT47FvB+diMOSoyJWMv3hH1qQgE6znyUrTf+0+ZxAjw0AB+Ko5aRaN5ddBeZ
il2yAkx3+iOnN7B0ZbXxtWTdwmBkQlWJ9EpkUNKcpVg+Ag/U2q4vNxeDfylZVQtK
jecaqiIFCTDJeuzTc7raa0tuKTzz+7ADtrK6DBUkLaQwPQvUKPgO+kFHGSwsPIz7
bSTi6/L2z5pLPI10Ac5zI5oDdp+pj0Jr/LbRkqC5cxrrHgZptzhKt0U4GE+QI/j6
LoN2oWKPJnUCUWaBgwB3GTD/exCoJkDbyPOmW23Js7/yDpFQ48XF+zgCvVLvrj9Z
gZ1HPXi+oypdhXlXUzwhtnQM9ZlUsQUz41LcXg87Kyc1N3wn1P3Z/498j0v+ih4X
9gCezFCp49SKmHiyJDaNDq8VowzfU7s+YSLyFIRNgEomu0VaDg8CHiauX2eoxwdh
CCzXgZuotp2i9PKbVeXeYnS49A4gWeAsiOJAZ3jQ1tbWe9PbjIF7VTtlYmqrz6f9
4mYKJdXplIMJEusEa6wVT3dEU4U3foFZ3MNSPRw41zcE9TewYUidFPNABKYeXcOD
yH037th2CYPc3GmD5wudFemBfvCIrOZIHyec+rKxuk229yVqMlYqjoR3SYG3tOyP
d9fMJe8UOG9cQ1R2Mce/Y1j31x9w/rNUyTJODbuGCbt9HK6KMXA5wvbMPJ1Q5SSR
nn2hWBxc5wGPazRVEUWX3ZE2t7ZrmWPMiJ8eZHqSRfGJ3UD5qeAsiKLmRFzhZlLe
c6bib4cLxEFYJ4JcYDGskc7G9gDDD5umEQsLzt1QolvGFzNM+f0M8uLaphVpedB5
l6JLjO//Lc8pVY7CvuWzEzqBZ0vmVGQwkvYgx6BxxwDnqZIN0kqCEwmCtIbAXnUR
9GEgFlXmGt+rUylHGRXAEhWQmERqHgGb2xfiKVI5XQZdDEv8Ue0xY6gkhN7WLTxn
YRjeEU8baJ/yLdK/1wIUeCWNW4RGU4PLPUUib6lZFh1u6eVtZqByMmCDVm53jjql
G0pcFfOZRrqjmboEq5ICGsb+2ZOXWwDgc+HiARtSngfzd3ZKE5fgRR1ijet0TcoU
CxGJI31bj7qkMxx8iWWK0DawzEvc5kW6N45Z7rKdtl2QMxzeR2YDxDdiiPeBgXzY
wgpGFDRFduqB0+fQqVglE1uAsEorGMB8Hu7pEs2RN6ouKs6+bv6wjDhONEpMZbT5
xvMwVRkZgcf/h08FG5zWIrskPRm9zuEhJ45cuujUkuok62D/sDgdZ49WH02NHz+y
WpSzSRaCIxICJO8+uvArKovrrqwEpaU+7vsND9oSYeE2U65DlMuOugcyVEt4QUU1
5qOYYA6dQAqjI58DYAdqpNeZJNOoPl/682HWnvTJsQ7+sgG6ClgGSsLxjNBGOe3P
osYd2iRNpzcZOjHX8/Hn623HRM6geKLX5fI84o8xGHiG3GfJHvlSIXtcP3x1Fxip
j6IcU6u1ODeloJiP7fofcsihSK+hBMq3jbP4xWFJwwSeY+2uuEB0RHUj6L6+4Y9u
KxhgnA0UmLPnr4YzJV2tcBLGM+h0oakgB1tregEkf+H/1/LbU8paPUTanLWUR3Eb
bxp1hv88eaxiBurOEZvTyViMuAHGESRJexdD2vXOj8yaFe98F7GZr/0svXVoPOdX
zF0UvmGHRY3OUliw6qO//cILipvqCwgvXFKoMKWok+nMaTJEVxeaFOPr3mMYlQJK
eCLJZXq+c1N9j7c6LhT3M2p1jk3yKaGxCfqtSKnL+5YwbgWW6jD5TXT9L5aWkjVC
Iwy3uq7Jj57mTo4In6lFyuOlDSs/YWWBtKPBtd/J/ITFAqAhsN/1QAtusW4Y2zjw
o+GQ5bzVMse3SB3yR3l+CFjrcoDZEEsINf7v8bOAVz9EiNa1OjoocFTjbnMLmMlo
uN37dLZ5zohPfpSHozLgSu2Zs9x2djRiXdJYuV3egpeRWrw47cVNJ9HogTHXUdty
wjMRahPZCzaI0mbtycLHIX3OiT5a4w1uLAeli6SIQleo47S0dLNSbD9m0fqO8RD+
Thh/3K4/aovVdvtqBLlWtoswDhg2NIv6+X4NAmtBVEyO9RVXfFqc3/F7ee7mvS0Q
NVipkCc4ppCVTXTrzaKfWB9qh/lC4aAemVFGKFi0oMB8SUcae45MmtpOCZDAotMe
8lN+ZRBeZRP+bn3qFuWS3Pczx7RK9pBx118keRO/jgDSlDmYUnud/bF80WKM12hp
XpNl8b1t60McC24GA6dy6sK16FzDkdjjeg3efrGgvNpk+Ojxq1KfFenQSZh/0tL3
vARsPONgamb1yq03Gf59hL3U11aXBG34SlmycMbuCvh4ANCbOx0K+OqLhH4bqJQo
KFzSrraSvxKk4Z0mMiwO51usHdyt2dybWLUgduLC03G6elHujtOePyOHPOTd+jY/
XVv1NdjUsGRF88jKHIBk34rlkUadzcea7UgHphbVDdIIb3ePXDF2khgv9QaYka9O
AkhnFOHy+gPXKZtq++PHUE1MZRk9XMm0hSppDtZoTgL9fqzMYE+03YgDPG0cUcAz
Q/cS4ym9mDegU5nmymLNghsIvxmZNTBv3FKWqf7tysh4TBoi12WfjgfHeAJrBYEh
pNcr78GtU22k3gPHOZp0MlbmtAx0I0jcL/3VCJEeudWcWxjVD7kdF7A9lXPIKvl8
dt2mJzOIKpxO1OjiSUhkzNvHT+0VM9ie2b6/fXuWPuqrl3YQ9Gb68RiAQ8oW/s10
7sRlLsnxZd83mS/3O4tNbmcQ/vM4AJ/CMt7JWfQPadpvO7IbWytR6RcZPEAo4qQC
MpDRrJh7hut0t1pnukVlMAljBU42sIiurWU321Lrg99uKNOeS4SJlce+/H+N5Nyc
yFz2XJqnRU1yMN7b3MNcoMur47Oz5EcIqsjleFlRgZSkq/niaVpu3TP5Hk9V1Kom
noo/0JSXRI4yL7d9VRJHoSIXhP1GprbTDAhpXcFussQqXfPNKQWjs6Wx7Q56MxIs
gbcSwfvJxy9gnMlFcq9Of+JEb0YD12Ti5tZVpibBS6nqQA+KNcpESpHCLNh71nBp
nS3yhA7bXWf/SBalO5iGN2bSa3/VUA2cGOFuI40IPimFiUkN81ksuCdNZONyVu/o
hfTXkgEODkhq10DeLtu65ATNrpT5CHl/4I88quUfGcm03DUMjrYIz683WV255S9i
lxLgnBXcSd15Gd2WHuvfECi3Eot985zsgiTUYU0hE2/zns3emIA/62t97bWjus+k
JHSPZTvIvx2PFvj4JRXaVOJfJCvznC8mXbJR/24btr9VAk5tAaSOZ3lxLKBUGzrv
DwHEP5myEqfSiEIkZZzhqGFKKcUAOvWxLX60woXJrcsjubIpVTmBR24jjvCIvL2s
c5G1OGXaGV6bxb+t4VRyuvbPDSan6okc8JoiPRYx9FqpKAfXVXgrX1TipwdMTJXe
sxRCAdzfKHnnOmWkc6knTKeVstOD1i6sZ9V3gyeONvpqNc4/58N4Dwm4dxDbNUQj
8Tr59AuMfcScNiQXyyWOe4cr9ibGgZkD5bTGbMGOJ/AA2R4KKKfJbZIgH+97Zj9V
yVFnR1nA/cryuDscXDe+kj7JudEHtKjw7jxj8awnAmVLGOlcYJAtA56eMa+BRWbi
TFopDwkuvbWJLP/GFbFLP+Rpa59bKaXC57jzgcaf3yqVFRQDGTas65VR57EMk8jE
4mjg0z8lIlpbuG0nl/CbG738qq3aLWkk1gPhdm4ceEaryBJZ0+7WrFn1YtmfRNQA
Mh9+COsZ931kc/JXMOncrKUIH40sxRO1XDDn8HwMo76rQM6OsVcS5EbbodcnJQnD
XR8EoTvMWKD4jaHSR56MhIbduDd14IKQHEry/wcR8OEHnTt94BFXUOOa6oweYeP+
CW9SPUvJOIdhTfuWstUcDU2gMBTLdiAgzF5IpK8ss6x8CHPkBq3/R8ctPYPezIc3
Fr4DxH+YUbghhnlFEH7w4b1Nx7wRYDuaRwxX01tjWzh5EUzM2ElMGCNW2tF7V6ML
MeoeRYanDKCaP3eJdBj7iXNgmA8jox0Hx6rr8k3eVjavdhYIetZv8vF+VRWIUVzz
uDVPx6cg1n6sJNxL1jwp9PEPzNkhfSRvTJLcmUT+XMX/X8D5kxLQceOZ0ZRhNSo7
Wq3E3h6yXlkAZiD5vrqDR/Z4pPdtmEe++Y+DenqItstjEPl69q0Ed2jlmasOOT9m
X2UrohOZm9vR+tndTBceyisKaM/Mvqr/Q0WRM6Qnj19xeOMPOXk3Xj1oBZr8ZtBv
hbu/QWwfF7BGw9Mx0fwCLBnxr2gE8SXrA78yEWvBRxuSpMgtASEtT9WB2kX+/U/z
0i4vDaHk8iBXvg9aEe9kEP5X7lIWl/lR1RmTtSn7sQGq4imzM+VtQl5yCmZH6s5R
PpRptR/H67Ixw/XtQBB3ko3aENg02ZlQlkBdpgGa9D3e+wdbK+OlWToqbhPLunwH
qBvqCk3FCeIvEFO/x5YCEi96hxPGYcJg0tjg2xltoRaYYsvQ3iNvFKJH/x71iWd0
eX1B2UdbbQotrjhitl5OIF+G8/SWTBpxXN3PmX5pJz0ygNo1a/VhQgfa11OtjhMQ
rJLMYfMxd2JVr4PndzROtmcJz5AuxPlimvrynH8qdbqrCwnT7XZb8aMoaX+k3pWY
Mj0wSPcQM7n2+nrTr1hXm4rkAnqhWb1pLbiHRSHSGKcEWiO+usQ+qjwt2cwd0NWp
Co4Y+7xxxPBqZSt70qi5MedEsacyv6Xqqccsfta5qvQSMyvmtpY74YrY8EecwqvN
YPd1ZN68DWINi5s/Lb4qCX4nOCup6LdWJUWyM6EmoXGrFYSEAXmmialGZCrWYUTp
CLywOQCyUfcEunmv4vfmDhRNW0eiLOAd6twwbdlutG4nL2xm1kY/+eCIh+GiUueI
76XBLZsjDlx2tJ4peLR/phVxd6VHleBSdKD1EA6sgDQZC1mnaryigIaeO49LQFHV
Ln8y+PXDEptFG7iKZe3ywDKErxj9NZqJJWTka1S2U2CNmhVBS1uqILOt2NXVQbmz
rRx5MvnlrNM5xw76yRXUjdGti2QYzqa/h9RkpgOzXTo/OWVMuwLdLuNi1BW4YVEa
VrWqWL9fZ4suGvHe+3aMKDGg8QIuuHoQLdzRr7rcQWkWjdPqnHOqVdaOq+C4bLGD
n8g5CchJlS+h/XMeoIOs99QrCf+gzhKBSIhzaNBY9cgbS2HYU6UH6MsZSW0s2yCZ
huza7CxFwTNE8zsjKIY5+kXslXPEyRiHdJhzDnOZNIxmKjrHxC4Y7UQON7YysAGb
U+TKAwJ5qqxMhCR1NcbdEh/4z02/DKP6DYUAo0/OtFuMeDBAnrcvcV32rFts2IHf
4B83ykYf2xoCUCWMVtGD0qreMgfJxbGwZnv3shZoGPq+NfGHv4XCbyxfRfdr2188
gjLKk3qyOqp29OPTGUZOGkgN2vHe7ce/ko5YbyzsX5k4Oq/3iPP0xWeYTbrQBxiZ
QEhMQFdOXViFT9K3wit4K2N+J6zLY2K7Qh5T8rolv6XBV/S01ai6J1kwjOKuMDP9
hvHfTvJz/mgv6NhC34mhIGhABDeFMmjVq1eJ9FK17DOwkU461g8RMdIXegllXBej
YJT1tMiM20m/5vzFwD2svNO0cTn3OK8dfB3xGy0pYaG01SnRCque7Y5G1eNmswIH
RqY2V7hOR1Hs4iYi08XKq6rJFzkA7eMLBmWD8CiPJK8w1+GXmYxL7zauksD+C6BS
1mzEWgTm+brJ8oTwuF6zEDlxAOqY9BRpyRzAJdJg4yksKmX2F85BI+Q4EQtNArS0
aqm7AYjMXf5zy8LNufjLjn58+nXJpo2v9x27WtFFiN6TQoZSk3ijPjjWLXBmzePo
1hcsoUVG436/h6DOOlUYZCzcHctw9ZiVvSvbEaeIpCRHQZRCno26wDRQ+Ypnp7FS
sGj916inrr+YcxYoeA8zViFY+HpvsqQzd6QWClaVuGqf2HYdoFyTQpLbofhLGtPw
SX0qAnwVF0uO+fpCKsbo1cBJ4obbjzgoUaPJImwG4/itqAvoTzqRjTlPx5osV7wC
j+yFhSAUzqqte9q+zx5vVG6093qBsyXrfrDtPDoCRFU+XcIp2AXy947jBSF09Qzh
1684nJcy1i3ubLjRLoeMLyM3GASh7LJbMEYEwpe7yFLO5R9IG0W3sVfMQJhrWWjC
o1EJb5VWrHnEfMOIuKR7+WAlRWmDgZ9ZG8jgBFP8IzapNVBW+DvVt3Baj20btu+4
jCqB2dfd5iWuKPaug0PscMmMyybuyh49/Bd7VtpFwkrfna3iVKNPj065ehgB26E6
IG8tLIv6hTTuF0h8EgDgM7aKQd55MrQrW1pVfC1ZrYY0PKl58/0cUlYdAc5JBxh+
calI3kp13qvWwMie5UE7LCWHS/njEiL5RIVpZJeJmV7GnpRsAPgynRUMgukllA3w
FowG22OWeKRKlvv1S9zDWN/NDw7vE8C31/3EEqH+FUq+hMbhCgjYEUZO6kzH4JYR
UehyVs1XsXVpHdRIXWSVTIVrOaGF91IKRXZN6YEzXcj24pMnzp7rqW6YKC46zySJ
H/fHmUsMlhQupp3vhOh+6CgAFnu9hEo3hCdV1HhRHYwZXEdmymvJV6feWeVET4jn
PKX20wONEhJ+529Vaue2npsX8LSuHhn1Wn6m88WNEdFXDlbWcddG9nXM1DwMzprD
pDwI5VXhlF9xgIT+4zwgAJ8FhIrttdAjI5mpxkS8HpZVw6Hn8vxTo/bdRGHiflYl
dIcmiBqrBzZvpHMgGwYsIRaCJhRflDYpc5bCyNMRb0xF1oeWsQOHqBWoMz5//cYO
lXPCWQ0HP4/gNb64+FXCku6wJU4N91/H6Zyjhw9k2Q+a86dBcEQ30yX3N/qZ2Nm1
Qsu+/PQS36R+FApXf+9r41wOnHenh3dLQ2q8Mz+ueNN+qs6pI9mPhzJNkANfrImt
9uOYSSelBSIgm7mWFQFgSEiarLFRELh3x+Ld7TJgjKZKMntVo6EI/CEwga/WLCsV
1t5odVwuVYsFBGoAGc+/YKLWrJqs47fjdVLmvEMjW7HDhbsx1MaR6enbtDa8/5p6
D0o8/HH1rsGYZKYpxtzvRzBybpr/9O/DBz2cT7qfuCG2zmLTFJT0yocyOWUVZufp
C4FTps/xjcb7qc6i4u7mtW+E0iEHEytzaubW1Vem149cs/7d0HS/x5NxWagJ8NNY
dQ0ja7IlOTsbhrVBOXT8LfSMWD4hKRrWBMbFXXlAxpKCibjZzOY9PiuS36XinuVA
LnpPL9UNRRxgaxetOy0J8CFndQ2Pol8Ze/h7IxMlH2+xKKdbvLAZTcKGcK+yfOgt
G++ylPQMk/jCsZ5ZtDcooNMkC8ySXN3yBBnU+gozFgv6rS14Q/cTMU5E6h56L7B4
kNT/ojvlxAn0opqdN4cYEoayxR1UWu80rvRHIO+bGkF2Qo91Ua+Jup9a/cnEjBsG
0+JFnmUMH4QsMCXUZQnjpIuSds/qkArtk9g17cx9KMvrRdePiXZzzZudDJjfU7qk
8GGTvsd2nVdDZUT2vAR53lhg0CvkUir4f/86HQ+am4EW9OxQYCIir750k+avHFnA
O2t9zV9uQxTeZgNI0bZvYyZKGUtu5jEVcUOIJmQfPAX7NBwwedkzUWmnfNk0odyb
uezMC0T9iB0NXKzl39PMd30QtUob6lhkNa3ynQhzmFtivHvc4RhMBcBx+9nSE2BN
PJbnyFIQMsIB6nW7MH/S1U+PZ8EsA0uoyz55UJHA//6J+fb6vKWHSbMkHWE4BEIt
4OdcwazN9x5hZPwkl/yA64KYrhbnMdY/YO43rb4uSN3Ex+lX7zhKGiyXsPGznekp
w7imQ+EEheiR5JfjF4qP8c+vRp6zGrrqs2yUk5ZoZkaqu7eokkRHJ78K3i4gakVO
AbrhU44OaeSgyaG84EHLuJU7IvxPIIosKfrG0R2jBP9qwyN4VfIswKLJX/kx3ysL
3232mWzHpN63H4D/I6ZjVejhC79Cw5fIy8kukKvxnaBb/trGYZ6WfheELkHJFzYF
4VNzofNZfh4SF9OCuvrKaSNMahzI1mI2hH574lQqOswb5lfmC+ZpfUTA5N0YZNYy
Z6KJIz/kyZUsMqpcJYl52H6ju/XA4R6qp0qO+nw4Hz8397f2jOQQjrzZqFvIu8YS
zvzG9Sg+/6OsWZTaAHrNTWBtmhVgeWJc0xhLy1G96Xq/57pxO7yk93XNuOxhmy2f
YliqABWbjsO6i9rD+esZbysTS2nQ1n4X2jesyxB1L/ddo+mt8IZ/tNfGqnHwr8q2
VMqzKUIC9B3aacWRnV77X27uKA5kGUKe8XxYcO2XqvB+H4i+jvVaQeoq6L8+c8gP
UJk0yvEkjDEiKwuw8ApmfWcMjoCQfZwLZFgw2GsMTiC75KLXqvmREJgryhZCJNCp
HBhFn5gKHTOScBLHJWaGV5T0aaROGdm4tRWewlB33/shx4ucIaCnV1fg9cILjQxM
kx3OjOJnPeVYK3uJA27gRQs7fQhhlOD/E1FrC92UnFlZGPBPu6d6G4f57jwRrsGh
9dWYJZJyqx4OR0cIcH8lqj0R+1l3ROAFl17Zan8YiJnkxqFOT1pgBslZchxCtRIB
kchvss/YBpdE58l//s62QqYzO3WUyXOSN8jzjSCx7luiBw7lKolzQ8tuxjCaB1f6
7AgaYHCF7RhSjvP4Zc0Gka8wyttM5qcSsiMFMRe+sVj/mz/9eYjxZBWDNiHoKHKh
nYNM5w0834xPwPzZXnsA1l5HqgK/T9DeqXCcxllsYCb/eZAST2Ve5MIFiZc0zC39
MRAl8kzsMyCzLvw64uzB92Uco36n7bouotIeYjYETzEvN5X++d5IG5aN1dwzEbQf
wc7scSPvPGeJl6rYVdIOD/Afj2Ht/PnRey3SvgmP3ocElf0PkFyxsSH1iY8Q0y+0
sZqPbIjJgiI6qzvxK/sXMOUwoymvfwB7h/c8L9vqGNJhm75nIsW2aLP0jnBe9X0w
bc0V6aJZ0hdmTuk2iKQInmhxcbnEPkav084UpwNAQJK9Edne5hSY2iT6iSUtvbA4
tJN9HZyx4+BZzfH8wY6yCdCj3AMYj1zBynO9i7doPNF2/Um9qnXjhO+aIgTFaeFm
knhAdQ2xlBqXb5KO8NPE178loMv9q/tSwotoS1IpRLk8jLOoJ99THdIwbX9Vq1WT
gd6iB3cRdvSvJUDsnv1CLR07m+9QC9hYjfyG8/qtjVj93CQjaq++uBy9sOdo92Y9
3yvpGGEVikKZXgNFSWy8pvy4FPgjgg89ESdhQ4p6nC9ukkAO/TMPi+tCll0AjPI4
xQkWHi3rS36EyaJciruK9ZtCDLLSWkBw0M5yPlZKczYHI7OeD7pSGpetRz/hDtms
69JTBS+R5L/VJ2hNjgRPKnpKW4u2Ft4ikRMF5OOEpGGNcisJybqulamWI3715teY
3aUV1WaRRGzD3+hyVhZsCGNgGcytuX5tb2LoaRzJbNtpJ4wK6OTJ12IKFplIcixj
1vGPWmPQlQwFxBKFlYQYZoKuCZofn4eqlX9raURLxb/QJxz/oGqhkZRMpFP+Yuxe
NBMQ4cqQ2sF3IQFrRfDhP/+39Zey19pZwdbV00L6yWy4GcfC1m1WPycmjzqv9NOS
WuiJ5RLOGOxUhPBgoH1BPprpxP1/7gkeSODl3zjbfnfGXbZQU/thQ9LwdOYIdygv
g/D5crRItvvL2W1+RTZnGlDsq7R+cdJ+kDEKfPbkeJ2+ZMHjR32itV1/F3o43bfZ
SGGH84Dy42jJkOhlJ+TnQD0uniDr85iqJwst3BD8fswrfSNawrBkXGTw+hNKKmQo
6j7q+gnb3h0R44m40z/CXFR5uX2el+KKt0Cxyu2VaTrjkTTEzk1omJF61IHL6SEF
2EUIJf5pWKUhIzzrPWXWd7gxT4IM5Ul4PVJ99jH0j0x8VCatCvp6DPv+xwYJHkkL
J0HwPsuazhMFTyyurZieCNpiGEGk80NyNm0pWhMcdec/vx6oxoWm074aQsAR3W5F
gXyDE6tUw/r0Ili47qbQPweqV9KkCmKMnneATO2SO2S0W/V4qqooPQlF6KourxGI
XEm0ORkxpIZM22nnrYW9dBQvWFg4/ex9SEXxNgyHrN6x9Y3Zn6p3llGboXwlDSPk
1eVg/VGaEiwJ08kwW2YBDro4pjxB7WbnuP4sE4IS7c4j3xMj/nylSGsvw8t3EU81
yxfJmPtu/2qMaJxD1rgP/CMqyYO29pvrEPhyocnyjSzn80g6XbMhIFd11AO8U7OF
EtlPMZ7YKP/a5CjFMLmRz/Wou3juw2tAqWwRA3LVqHifZfRiu54nYRXlo8R3n1+M
lCqr3n1PRWnSMlWZ/SeL43vqEhvAyyZ4fqwRm6zaB7ZxLdJXsfck8NzAyn/hhvIz
fscb6CP7Yr0nGhDaYG0C99DN9/A0Aq0peMdshoQm3d3lL/sR3TzDcOzQRcBGynSa
MLI5wx56PxYMZu364pw5C5C6IoZdhMdiXo9lX0+veagMJI0RCmAlizcibTEp0teA
sf/8sw7mniAj9PYzR7q8rrC7qLMYAXJ14Ex0crYGiLcOmFOX3J7yVF+bW8JC5TLD
N7p8/20Mgc4jbd9xqdCHlRUqq75Hnj98sXcrVZpOaIKtirKzDfGY19q4fzZLMPZT
cVaJ47w5JBCbnVkxF5Oh4hsYZ+VNX7U/G+BPLL61lt6ekm+fTf5QzCJxImrdwr09
pRsVaMAZeQxUvwWfhpGxKfM0Igp1x2wa7QaY3ccry05ePVWLnNS4hBhfRGEf+eaf
e7Jj0CfSkHUjpGBQq2qvffRGjX0xhyh1Wgcvf4gL/I8quW5HKpChLNbt9ylbM4EJ
AVc3M0+inbPqzhOXCqZ/UV+LDlxYC8e5gVUlIabTDJ4XX9jYOp+Tvm4Y3T6Dvsyd
l0HjKANnrh8zRaPlEw5++HHSiP9FdyOj1MPDpQU0EMHQSYwDIr2Ghl2xj2I3wk1W
uVw+5Yg272zQyua1lasMWS4SThQgvlyst9eMwIZ30YGEH1Y/vNn1wdAJFoQlLHgB
qKXinpjOAfG9mLMrgY6K0C3sTkYzsIDPklf6rfQsLDWOWc9FBJ0kQwe76dYy9u/B
8vA2a7/t8/IkkuCtpJhSbumJ/lGQy6UBEVKdYmEQh8JXb0Zi35bKTjpTvHhck+Yt
oIk4958vy/3GOrqbBRjg32nr8SgClBXJuQLi7V1tDXBFRTq2r0QP73gkvg8zBQpg
9w9UOt0es9QFJGpcilDNpm5NQDzUJ2D8SijguIvzzt8NSHBEFgz7+R4ae2bHw/dh
K8lGyCNXlwdNc63KJIbHkf9KSzZAJaPGGF5QgClhJVUPz08SFLP9mz3HNnGHH+Jd
RRvKpAJhlXqYsiwtAmIHfnDBROYZk1yBlHh3BUmNaSslSYN+XjwU92O9x9wnvqzt
UUVdFewGUgxI0R1cJaNyF72YKBTnGC02GBsmfmInc6V+5fR6PNBXkr1OY/b8NyCB
SjZDl3YKpYM5BmTyXTmvK6+Bo4nRGojrKpdmVKmM1AaRfz2UolawUfORZk7z/92r
Nekwxq9YNRE3z5HVaHFQX13RrwA5HerblufQvVi7Pk0CDWW9j3NO9AmKffA+r1at
jRp4DqHpZVFOsgJn1gOcsCsNYzd2/uBgap4ajPMeTfeZR04qDvbloMjJjvge0GsK
Ri2X9u9VaacESAp6ggpIuerpsI4h7wzqeTJwugZMXU/QcoK9gzOshl8QtV8IHMEH
63PDRxmDnwJVccnpF8Ez1zIu9M0SjwKVDM2b7LkAUC3ZLAhuK9Hh6Vtb+fRdqHcj
Tck8ib5MhIAAEuTbvVBlOvGVQZQWAdoIzwVaAn6cBCvWqGYwqosm8/IMsseppUhX
rOe5OfTxnTQfZ6meWJUNF0JHAozaKOtWfpH3EtPJMqmtf+kLruM232R2YckjRCTT
9URSMtfn/a/OKus+8BqBdNKGSZEHSzUGrVTTEPaToJmxaT529XEpJPM0IlafbeXk
7sT9tGG4qTBUS/3PXyr/IA5e7yv5y9+nVBxVlbOl5vqtk8BESpfJW+ossHGdgU2B
vwE7obfKQlT37LBUZhnjQHBnEbDpF549g+rmbUqkFz2rTHbZgkZLr5qZMPOSPPNe
edBTyW1hIWQulwh1D8I3VF+03UWHAU97eh765KGBAdzsqlL/SaQPG094Xu7djHYd
ZbwkKURnwnitbjgAycx3unjCz2/j0ktgpsQCzu8JBLyC/h7XeNWk0ehciKNLZlwC
xF1sxXnE1fENi0HCw4CxoAxp4HR+YL6xzv/BO3yRt1y7E/jxVIWl2bVz6jlzvYtY
MrkWs6cWxzGLKRw5FyMjB8WPcz4dQD/EKRL1dh0ItywmV8L6Xn291rGKwuCRpC7g
JET+uMA0dbWJI1wyjAZ8UjAvteavG4Gj0Plu4vATh5K03SSHFUboiT1EdeQRFLp+
Q6HVDRFZws1NV7Vxu8kf/OxFX0s2Atk/cpKM9U3DbnqcjS58SPzkg7L770TWGqis
I3HLsEKEK+T2ZRNp5zStM1f4RLQIHTIjH8W+ywBM/SduvHTP66ZiBCIJD+DF84Cf
LC7SlBJu1GMXVCl85+lmy3sSwcacXOaQQX8altETa0bxrGt/Pw1r2yjFL069eD1O
JjT5xsP6Qgae9IaK4v3WN+HOdPYEhLYJkD4sHb282prrxwVqr9LJF3hkHXcJED+i
500hIrxKaCaDvnW01PFN/wptUqhoboLSWall7zI7f9lRonJvTEr3RF7tiFNn6asZ
bCd4k247WOBMQ0M/Njd+FjaRJI8ilucekFS7mmpQtYOuIx9tpYHcHll1ZGHCUR0B
E1gkpLjuQRsLDOIsfg7qXPCWS7wrZRTOqovYCwDO6AnIwqDbdLK5x4w19iohCQuy
khDwUUAAGfLlDgqu4o2gspak363NhhM5GgsyZ/1m+E89xJRnosDNMP+xc4tkDiTs
FTNQxk9d1QacXQql0n9eQH5Wgh7b0NHHQT+NQ3mpdscO3zbILeDksnRCPgv4An9n
QIEZrrvQgl/MrMD4GeLqdl3Ot5CsdNWPCRPnbvuZgC1EiYJbD0Y+c5WWBtjGq5/g
11aY6+ZBvlxcrlYILeoU0nzJzx+CDf0l0QTCKRngjLzZ3MIBhd4GgZihbpuKdRx+
EG85ZWrqkZtVYl07rQTTuNGb7pzr46muU1G5EIR71MgJcU7S1yzHTcIBt48XmeMR
y+Qk+qFz7lVIlxyxv8aO9Dsl5Jt2iTaoo+2NXqbNU/nDefHiTuag0qp+NqlePx/8
pYaGOUBJk9tN+orcUJ5bCgMYWjey5JcRYnkMOTckI0AabVsY77NUN8RRAq6w81/4
2AyVGMNn9BzcGbO7PfBo+6Vd2sa8l6cpSxxrjIVym67+BtATPlCUsl5NPak46AMT
8hGUyD7YSxW5Xc5MryKHgHCpN/53iWHrGSoHAx+E7e6XV0/zzm9mGjRXZaMrIvf3
r78lBlWrc5kyKNvtrNlWmWE6zkA1iEwr2g4rVq4rIUsHEa4wGLCbZixrB2MEd3Kh
EKwTHvYXezMiGVAmqi5/rXrSVbtohAJ/ZJ7yAH8ITQdhM/c+UJbRsA2JZxdLEkLz
yQsFHTDNPeGkagetRU9+LmNBzHRBvMZRFlbjtO0juSRVmpST1K/POSdrGXF96aGP
CLpzLZa/0aNRktjeeRhWLwu5PFUm9v8z3PgWGab4lTt/3C+sfRWDLtZe8W+zqfbL
BUERbqHhcfD3meFfSlynsHsgVtiwixDxXUc0+o2rq1cd2v9nOXKxPaIl4MhTfZR7
03d8224iyqY5qxFO9siBJUxGtmodIrUxLvRyzhyhmcDDz7l8D7uH3mfLH3Nr3ZhO
Ajnv31QiLunDH1PYtAispre6K4eUR+Lx4eeuNYVrtYj8Zkl3g3bM8PEKvfW3KQh7
Aw0WWiMr9HxdKPZu4eEl2jhyiHDN5MgDJTW/nA3seD3dC8sV5jurucg5Lciovipm
149fwsXIPAv4fIh39nQlCDV2eXK58Hyi9PlI39zKBbz1GSA4olJR5q5iulXSUBAY
U442ixw9G21TvNMDHTcY/UT3r6NFUKW2IV2kLHniJort5BZ6fY2xtv1jbJ5FYNbI
QZpqpSnoPzgHp3lgyBHQSln9DATSucry2zSEMHjn4kV01KojOinpUW/5j9655a3g
wQ9S07LYAZfkIsEa+nfSRxL2yU/8Bx/cUnKnNPbTU6jpfBlaJebfm7avVyAeS410
L/1/rr3JbPE3j7R0WeGyM5OOTYWCNcKgiPVQg+Tx9ju+973Zz7NcvtfyCKUJjHrE
hqC7xMZPq0ATMOL/6DlH70RwB0FZvkgM2EZ6eJRgIWbMjHAMDrj1Nl6GOuNhNkh2
/2tCmGx4hxRzFVMM+Xs553oHOv6gLpmiqq40WRa4DA8uKaX/r50L9mdFkVDCSMnr
hcQtIrivyaxJtmQaoWpkBp8+iXzABMSi1JN2RGYiiUk4q3W/kjuG0FVy6C6uGBlI
KL/AzvpIPD63txtuvkbe/Hv3LRmu9+Edz1usoHWHk1KPVot1QlirKlgrwsNFUlzP
zmmcPkIbE54UniwbfWdWo6X/sjVGR/L3lBJE8cfBuSG44utAWuCQRUjZnzliEeVV
q8fgwFKzBRESFblNGHa82CUhc95mFXfHj9pb5cAj0aWyCz1EJPWfIofTxUcthDUS
SLBklDb5u3oD5gyeQGzJc7jipc5IFzCSJOa5osYrxCBby18A8mL38/4nHVbd+6OY
P1g6gn5Dkb6J8pOD7l7fcmyVJtwNDXU8KKV+xRUMut8EUW3/Xx0S3gR9FRKbA2I5
hYwRFmhx5ytAG2MwBrsk539Asu9nxcfaJMrK0K3VckzX9o5iUra4nzQqLBtfef5k
Nbn95xBo8FFu12Bukh8Wexj2gQX69hjaryUYxeTAWlN0qC57uvY8p0TGeDe/EiiF
XAM1XENJQdrnTPoW1PUplSNjV6m3yvcEtRDy3+IEcc89+yXCYEJeHICfMEs5a0Ao
TePGgOXbF7hmKbCaFMNFc1EUquQCkd6bJWb0VBNimRqRMSJ1cgQJTBMEsgaKLwFG
XqhmHNl++v2gPnz2s7ZaLoBE4k5K+cXO67i7PmBRhtviITU9k/xqxN6fKCVLaFa4
v0s5FG8gbWn08srrCLV3v3glQ7DgkElNvzZNHg84djut/oLtrM8ZS9kdCl1pihVe
IsQBoZ0N8Ovsqfu5EAn/nt2HDcJSwiTGWTlIUYdJPElfAyJq4/j2f+w95z4ps6Rn
VorfP/kL4erxSTBC3dfkT6+G3Q5VqtEXFjArEyzQEXlQaucQvVwRSJy0efwO9o6T
EU1eTOY88cax/j4cn/Isrvke6mopvJmAZxZblMZTqxuJ3Vm3Q1Y7GKEkkk2a/Nvb
9rwxQviP4lcFLM3CgjDs7fUGStxUk+wuG05dXJdQdkhti+F7lsVEb+qbThn5YasB
INDcdDUtNCOh+6EO0rV9EkPRnT0z2nfOFGHO0om2NW8fBu7kIG57BTinu35owI3L
mYAJJfhE+64HdsMITXVtIJzUijlY8wF1RxlbjNd0bDEf/rdN93UH8dlHbE3BAxDE
YLUMlkkoLd8uXRnN14LPtNt9JabY4ae+sC7zuSppyvgqsvw0uXIV+kXaedy9xoW+
VdXw3uIHtztc5s50RsBNBa1+3JJIeyh1WrFDD5WfHPwn1B6284UXpUC0MQyJ39gA
4QJrJhFpEhSKj4OZbsws7KXM+AH7nh7UATX3H1p0lX6yKCyMEOegRPV6/oO25lUF
eSdJYpWYF489YbyCnNNu8scDXXNtBc6UQXtjwjAOG1RyTnra+ehiHbs/XXUr0qDg
wBqZkXhSDjq4P5iYGzE60eDQPGymsKpdeFYQPkQXK5MrhHy+Px/SLSq5aCTvt4pg
dSvITUlP+BSwacPLhW255/iqvLH8BW1ZwPzn9SsRqdtS/vgm40KDPJxGq+XgwVxn
mGHLRS7ziu6Fe+iXYML3Et3CMHzx6dK1sKedmgm/RL54lS8ssZgk/eole71amCf7
jGECN0Cl5EfPYrdJHnGUA1MQDT01ErKTl/Z4ujr7hUiGHzODBVdNHasIQI3gxVN6
xDg7RfVzful50O828+O0bn7p0u++YYLk7kvmvfvLaN3wF5/xBfD9CZ4cMT1C09f1
SgLNaOqSNABlKbmROOuNAISdjbsgrgEA9M5yHIJ5u5JUHQJq17TbXqpawNbvZWbn
pBLqtltANCSHkn5rbnxyXGrcAQdhUA3kvxYrHYmjCRGJhOgFv+Wp0wJnBem6iL/Y
2yxljPTIDiXSgr2dNtBkhwXVPircHTMZDIAjS2Bq+DdYFHeOo2MO26cqmI5jMMuK
2PmQRz2fHxVgLAsKZRfflbu9RfotK/WOkyiMINMAyX2lzhDOvNy1uppIy+8EMr+z
e3lKJEUa8dNW1n2EMMDmLeoakiqkyS2edZyuQ8blKHTyXT9BQxadeyohginAHeVi
vvFwsWpF1QKPvq4F4fl9Ei/xVn+RKPB6yWD/e8/Yva+kOCFUKC/3igy37cO/8bjU
mEBit8tgPi5SBfLbDZ/dZoTi8fKojCWzzg5CMIPdlqXdbNIhPcJxvXHCKCqI+UmY
eGdZPCuJUzKcZZJ6W4nVErNbw8RHhTyLTAB1ykNMRoN9csiB4eCTtDLLWxT82WiK
MeKKrOXY1zQJUoWdRrNUimvPgd7Bp+Li+gEbBLDfK82ceGH6gauxi7HY/PEEC63A
/iKHQo9bQjqtLeftvypxc/xm39OfeW3Fz7+KkNUdsSEZl7Zn9Nzi/qjXG4oB+zne
wUigdguIkxlQAYcTAji8i3C0Okb00g6Ld9EiiVqQHomN7FRMlnPLOHNWDK5fGXdB
zI7aosiBEWnkKkpR+lPCNduLXtpjHsoWzUSFf28vgvf5bLI+jkplIAZyIPfvQFWW
ZQxvOlySm0PtKTCOYgPaFrfcaPrcCVNPiQBmwzoXdoxg1DcHTK55g2wg5X+OdHze
aWQ8diNvQgs3yKBBOKfMpvNNRTycsEvAaCrGvdccsjSsYJYrXoz0K+PZ2YeSwi2S
OXFsJBIQ9TBJNvb39eurrdPjvnO/AY+4MiVaR1jWcI1zy4nEyfuK5arCsVdGiBrs
6TM8USGDZsiflkOSluWACn1eLRsJhyji5AV5xAr4EmMu/lJEfQvYlxs2Fj8rhDcs
TBEpfYORt50yRGFV4EsHb3nGR8Gobqx2BesKBAFdWH1jO4BhePaZi8MEdlgp8501
VpsM0E8TNQIQM9q5d/mB/ORY6Jfn8D5G4O0odNHODD7MiQAbnunifUce3kpHb1pK
5E6IYyFtkaS1UlSTjl8v6vaISH/M8UAR9EX9i3jqxuNeV2k856fZawhiC4JxNLGV
6veLARL/51sRTPFkb9LkmMYHfI+XPXYd8ce7QpUIowRo1U88HMxcV4bjjHErdr5P
L2F6Sf4zvAVGCC3v9N/Sx358XyDfJ1LHWrWAPkM8TiSDLCjJbGDzSVcPQUr0xsbq
OrwtIigad2tJsMCB6NCjlPMAy+JaDnvigE+6uqYk5xTmxGKmiqGtnUnphYF8r9+W
KKinbL5GK2FS6IoZRvXfIGXktoyvZCGfecc9zpkL790rjxNlXVJye5R1HNRulcsU
O3UIpneBHyEPf17D1of7trKMPb/MXyCKnU9m7FWsjLbok2cOmAz4VOiDq6XSXUzm
4OOjkWc+Xo3jJ1FhDkD3zts/1acn9zGgkziDcAJehHjvAJrbXVNWFxXEHv0q/ftb
N72jhyHpiBAluc1mWZnXUtxVWsg8irsO12G1XB8KCAeR8jjUkAs73r4JimH95RcG
gN+YL9fJCJ1vEKF5ONoAhfyjkTresc19pcuBbxpU90U9DOfMep09PIfybUefJoyD
Pxdwa7kC3r+n1uKt1ycB64VZahYBLhZ1+pVFb+7UCt/cpJOz560ISar5Y3V6Rnm8
L4uTB0nAMH5qplNACAY8KRYrNJ34dIVT76ZuDbcVfnFUk+ne2kxmoUFCKxpClput
jfcCKx1FesmYmXEUqmjXjS39xnT/RziHjJCkjTkGSYBnmpdZX85NnDivydNC1xNO
6KUbx/efmCKw4AVcm0tFZECAY0AMG+u3JzoUOckeXM5ay6UGUNV2Rl1U1GxJGffe
k7lE4sa3H06V9s9CmZwF8AB6hZmhrmSYRedknpfR3fmapouLsEQyI0B5EP+eiQnw
Nzqht44BoIR2p2gAlIPC2WhHUB6ZyuQTPJC2MX1bXVjCebjA0JK3mPYfiYO9o21Q
Qf/0a1iCcYcCaeeQYaUihO0JjaJjnw3dlhCvdqNut0S0bk312knDRmSgAS+onjNh
FDINSGdjocQ3i/c5jZQPZjoQq1hxLE8agyphTxhRlDxzufm2LkenqbJAq1Ypw3Jq
+SrhRif1noZOY23tm2LEH4xYmhI1OLw+Lws/c/umLUwCefBJIpYMWjA3HNCQE6QE
c0LKIjSulQTvo1oMhVU4OUCZ/84Gf9IX/GuCPcWU8I70EKWdIHLpdE8RWPh6YsFa
CLQ9dHoMheDxP2pEDdMZUkjpRL1ExWcXcFcI84oZeWdwAnvcGKiOg9pikYg2Jgxu
btUP+x5axP1ZQ0XPKWh9U0PKep33G+mHFw7lvqyywpD7Hh1hMgl57Z+I/3uNfjpP
KYoPdMJefU75GqtuFtQ7D8qgOHsmxiOaFVKs7A+JeqEAMbT2VGG+Juppk3hG3ntW
FidrkOqBgIhb0c4nycYw8RHAUGK+kHyceT3f6Z0+yC19qm88WF8EtlQ7ITuCPk0/
nkegZS92elz62WkBC+6+owBWVswRUxmFjghk7thPpxEcnNdB1UlbLkL0R5qGJjB/
t3f1uXH20Tlm7MtxEsZSsyKg0wG6SS/GF2zOs3Ep5iuqabyfunloOjr3FIkpZ6Kz
Rz+R4JhQNpfJ+pJ1UZBrpoRAT4S0hihJ1/SwBU69FWKKJNaQCBMH6tWgSKPqNjqn
K1yOgOKAn7vxC/o1stDmT7DPX06XZbANpYUDZG7LP13WecM6BmIFdD5fqI54blrJ
kNRkGaKWN547+tEbVWiS05jPb3RJ6rPxKb3FK0Fj+pktXdvLVHtAb42FsV1QIWoP
0lt/ATpxoNR1e5oQjUu8mhzYz9azzQ3w6FiJjUFfCHpA9/DRcljrg4wM5xYq1anw
IeKxNbv5JmOVmR8gbYn5eH2Sh6cPp86U7Gq8cTy9ko8K000q3a2Idg5PVZoB9qGk
XDXUtv+YyFb0j1E38XsuaulnkSO5bxoUoPTCPiEbRAU6Dyc56dSONtz5Ya/7Iz4+
dX7kDDu1geL9bd5yOgCU8kzx4k8cZfg6o0JB7tia245C778KzYdwtIOgcmHUh3MQ
Cj6XU0jNJ1k12cQV7QrdhfmQlnsVmQTWy7+y7TOI+iDGUIeQ9B5RKiWSFl4PmDN5
NajJfr2YTw9/h9cYg0a88iV9hx+s0EYfD+dC86xete2iq0yoQFM7lTrGer4Q9fqA
6hXSe7kBQlyfZf4EAXQB2vNZRJ/1VtzZ89/K2jvU5pyCdAxlWfYaHt+IBmHgpLmD
S7rHMMOtogUr1MJeQC7fScPwF5U7xjyvrcwKPaximYD5JXsxvXJnkIwxVenp1l/X
O2WQ5YOs9+SfG+8uLqMiZPlP+su95DjEAgLPovdvH/sE3P1vtPaq6+gep529H9BC
A0nKP77y/OWl2YATf1ea0xFbcHHo36u3A0DqATZeDm7txRbV4br6fSljZ/RcP8zB
xdlHL7WzG98+sykiCp6nRxTqMNMEvxlBSzAJV8HiFV8ndQNFIZzPeE4g50b6I4Gd
hpkFVaxorK1VBtjSVTpCXs/61OjFODoaWfYIwOhsuZAEEFJpz9pBA9ppIYIxCy9i
skBMhHYTQYafHQtKk+czLcawuD27sMpkjL9p4xgQQHt5U6xbxV6fKWRp38hhamEJ
IXFz56T/wtCms+RdRSGUdm8sVfJ0tbOQ7Emg0nT40ve4UmEO98Y06M62L3/MXaiA
cSE9kT87RIGNk9QNg0iKviKjM5Dy06GIO1AoeHUQqNwBaVJ+g2qSZQ6xSTLliYjq
1tujz+16gIIF9PIi7LRpqAX4MMNYEIFXpS1Tb2hCP6LhRFTEIuY4ZOxb4cBGr1n8
YLUrZu7Au6LpZU0ZY4z1QVqBK2JGqBoQQi++bYkcJVvUfDRxASP/Qn0BQ38UtuUe
hwjA4VMNPCJsH1uEURwD8dzZOLkqcNf1ZuNU1LLCT2/+CS/hTOLrQBeMNSzmb0Qd
W1Xjg0yubXxwnA4gLZPBISMJ2WJuNp6T5M80CD0DYLBw+0R7EFd0PcQJqeR8dCHr
69FzQTrvQbvA8x8zLJIwZvj0diDP9buk1YaEqTH365NPaN9tvMbSulkvL//zC6UU
AmZilmQN7zYbqHlIPJ3fT3oPNtdEzRIhTcS8hY65JSuYTF/+/mBBVl6R5D5/CjMj
TB8heX9qEsxiawPHK8juZkca4dzgANKYWbrgE+co0Y8z5GAB/5EG2NVhWu/RSk9g
0peHG3fyZaD58T4Nrw0yqm3Uqub6YNweYDwmLT2htl+eXSehU5XpLQGU7pJaWUPE
S0e/vacnt6sH95mHbJTqDPheUjPcqCGySrq8Hw8WZeOTOOKr+fVF1FaAPhkLW0B5
zOXbOPsTp+pgPS+mbgbNfGTrfNiHHLWx+uMA/TPnQLArnCAByjIusCPAOYRQ/wqA
8UI8lKtTg/PmAaeHtqjPcGmS+oVSf183BYsz9DsKEo00LLdjX4K32sfS+FDNrcc+
AtFrLdE4c94XMHAXmLR8dOeoQnZ8Ydbhh97UDJsdeufI7X42KfLzgxFR3zLMx3tP
wfXOGS7S76WGXZ8HVqjS94aAYp2c9hV49qvONnfHMilw8xQ0jC0vNM7LeaNbQj5Y
Nd1e4iWJKs5FIB+Rz7mo3K2zJkgMtoJNg1Az2/UpfZ3/w59M0kUScij9CkVn333c
zSBJwl1RmUAoS8OF4q2CF+0ERQhIkjkG7CzCzk5A10VBug9I3aNZE9TzVHW6WcVe
LDy7QY11JDwz2QTkNAlz+DTR6u82T4xJMDtM4EPLQoV1CQqFGdKAVXqxC2yqHxvQ
eh4x1rMcBiTVxxLlyfWtkBLKwnUkyQrM1xzMBnNBK2k/FOA3w9UhVCQXFzlkj4jO
mhkk0Pk+2gm9dQ57jUsIamZQb7RwpvTHNuG0r1+QcK/52WJWboyMgpOgLgA5SfNH
M2KqMRx3bX1X4AhOBZjmubaEGEnBbtsk3cy5cQ+TBM6PFFvaE1R/0T5I4wlBc0nc
U2ol1YZbavc/Nq/C1c5EPLRMl4CFg6j0nCcFsryrhaxFPL9Rluxgsnw745TpCqGq
/xaS/fYwm1rf0SRY6UXUYraxt7Uytfopcj6Oufh1S58BaaPfH8Aa/LgxyGLLVdDN
WKgVoE7tJBYed7MwopQWAunVuw39ggzHo6QnvEZTnAVbiEmLG0TMK/POq076NCgl
w3+NQcgDIUNa1CA33bSWvZM8KDRimaJBV6HhgLJqZY9mnRvfDILyvcHLaqo2PMpk
u/jk9kCYzxTe1KyujMYNnh0BvDH2UwH52g309otyBHJXuxn0j7z+Bn68K3maXpmY
ftk0n6g9/5jzCvMX1esotKr0aSHWIliv+hT/3WXsPgPao9yoE9itVgYZ80v1nK8b
/dEWl07LoimYohoxJ1wktXdn6Z5RHUwzopXWSzQp2W8e1w8ybpFzPj+rrtuBzRHE
aG07V1LgckSta+zDN0JZNobSAruyPpqogwFo9NeDbvintAZ/eIPvYzF9QPbmBijW
vPcWvNTIPZUeJvo+HGnJ/TvSJ92ZxucyjrW3c/5Md5Y3CUi4+w24Wk819dkoZN+0
g6ZAq9DoJ1FR/68ZFpJDx300p1yS6hBpUtPqBNWNeGd8h/aCkZxHkhXL8IiTN6W0
+zKJNUEjehEmL3MlAultd4I++1PDV4Rt7/FHU9yRM+lp3hShU8bhg361TzWnpC1q
zcEDGvDz+WqKr3vEVnxqbMbxf6ezZ1urjNIoEdq+Z+hVOaWDaH1X7IQn+cQVUtsi
LCrzsR30xjHRf3h22YAzxjGCLiUGhdXWirjw5d98jWTv9FtgSUFobfKkanvXJZ0b
KYdFMqgvbB4v1VfguZC41KGcIz/QgNaiD8lR/6TCNenq0DWMv/dtip+jngYtzR/g
rOdvfUAFRu+kmzxD5uVWci9yjFWLZDJXhSHStUu1gA3++WkLF106G7PQg3DQshPD
LG51xNCfFXyuWEK+Ck7EQWpVaQ5elooXlA8fPLbcswE763mpRBncLhvbRFAzrvIV
EaFFCSG+DYMZHIQS0DiwWd+p97uhLZqm6VIvR/btHXc/4+IC2hPAltXWTOsb27JD
W0pGcbI4MWdIeTEtezdJM8XixMfZ0nFxNhSC0VaAOGlAb/67mOwriID8/Y/Cet9m
OlBCwNpWd/XRIEeD12t/Jqz7+wMoZ0hEiTlTC6znFZS6Jr3RoxxubcD+yDd2H4Mj
wzpiuGvLSzpgljy1qQ8V8iQ1u2rDL/SY4OEvaLxjgwqn0GMP5TpqfCBsW6x038Kv
PczVpfrhNM3Q0xRCTZo8dHpH9xWra05T7e6Lpz3bxeHD0ILMNxYDV85hgwxqFgV9
Xg5WutsETNo7dhZP0f6b/sE9sVl2VzTnG6drgr6/T5zAUA6AuoO/iuAadRiSF43q
mYeABfBFHZIOMGJBz0l3b5VAZYgkuikpFYA171EB/P2f+nN7HxZ0dQjIlIgQH869
f8Kkwstt06i2FXL1gLY+YqfhbaRPh9oqgrW0StZeNeiMfdC0vPsv756Q3xfwdLm7
ApAuNjip7TmlTF98qfeiVucnqXCUgo1YnHyuE9BgC1wCe4zWwvXlYm7NoFE4GRcV
DavAxSq+Xcl/vJnfrr3I4T1RpCuFiKoi4ZfbnaS+SkB/lO2/nJeSqwpyKANHkc0R
TNIOUm+zRfeRUjnLG3Tmb3uhxPuOZ9K6WgivQ68nOlirnH3omvmZLPakprqC2Min
y6b4HvbmYZebIbcve7d/mc8R2gVU5cDfPBjCpp4ptai7QV/XoMnZF4ZtCOaK54Uq
OQh6Eo/OQ4a3RstHAD5zd7V19PJQxLZuIOrbszLBDpU3PX43A2m6MC+1ZK1sgb0u
SG2ZmbKPBbsjgAN9+SVOZcTh/KgRGZgp4NAuHSOqEKKcXLbiByKO3+mQxSYcf1m5
mJokH6uUOGNaoAnNEU+WRY85nQwo10Zyi9zxggpjCtzp9BhBg+/NvMu4t5oPdXeC
OzTr9CI7E53Pc1JkAKCTOucEP2jGXlAzn+cbF5ykq5e8/TmGP2TZjrzMAB9dlxiW
Q3l3FpGHJhfgmHlW5tK0bg3mdKlYkWMvoSN9y6N3sgDNtt4j6FrdT25EpfJktURJ
Iw5HmnarysJx4hXfAzM8keEveauFwsFf6GYAOaWFPiB5dzXp6Vzti1Wv1PPRftkH
/xF59kHFEJcW1g7zKSpqp+auI0u2AghTKV48bPeA5JZpxZx4QgGdfxRuMitVm9Zb
sLFIbGtQdIAZF2pu4J87pLCWJU5KNuXsPak3XW71YT8+nCsJhmxV38cX8UR/7eZa
b0JOgot7PB3DfBm/fKvoiLBI7XM4MdvRL/bYGKeivkz68KP7S273+II9NNKB+nm9
UqEaV8vsw1mwwdj6vv4TzWjl8NTrasxaghAGRrPehoC4zF0o63bwJ0TVNil+kVQv
UCnHZjApdW2tu2UmfoANf0zcGv1/AMTepBGyoJFC7ronxjHpn1rqFYko+K/EVCdL
6Shr0LJMTFBas68BdCCtFaND1B9gjiTQhBSUAo7KHV4fXI4dZSI5fVZwRypxDk6y
LjVBYXARERzKvAZqcciC4A+HNI3aOv7a0N7hBkVyjJFAUrPFiou5UWZ/siSlZLQy
8joDFPES4CFfzeYQpj9QpgsqabUsKdNmt48zgHdCxSSGDT4zlkTbhs8QgjYtXhxD
Io3qwcwi0iDY+0W5R9EEYE6Ikf4N8EF2XzxPjAE8KEispfrtEF2tfavRQqcJQM3V
nzCRBFrTnw1nOWoj34BsEFAWSmTL03RwVfTHgrqez5j/rPqjw0maZTAcWLGds0Hy
6wH+riV2nmxMBnKPm1Obt7Iv+BwQ23wuMln6Tne+PdMwbPMDfvTdjQDEnUAKvYvy
hAQCmcWujQ/dGwmg4ijN7i+VWc9hpGxb9xvfLJw8Xg5Dlest+rKi4fKbhoCwlsF3
nDuEdvW0XMBnsRni4d9qIJ5cs+sjPjTps33L4QV6pIPuy4FwjOEVmMKjEK1XdJZ4
GijimoyAJ06KLz2DFu2iEubFSp7SgCoeocqvHY7dzTf/ZAfgDDn+U/ddrXwrkKJS
bBVhTQonRyGqGcJRL7h5tLzuo4xE7+AbND4tD89VvOxZzlIqU1khWWMFMFdHheAf
/SWGjBzpsg/2H+Atxp7gn/SRyf18ECWP99rxdKtwdpm8+BnU3RSHn8jDWKxNR46/
umJ8VRYtzOdegT+HFg1CcY+cUP0SDeCBU3iHq3JzwZcapwhroJZ18IxCFhzflXpT
hBPMU2M2tmep0cDYMoI3rdRf0nLs0oSIBg7XyZzhA1AQh2u/wC6WaykfMSxwJOYT
YPd5AKTvCxloAG9wegqOk++LF5Viu6GMU25v7qYC5qNm+QvhIBnfPWlNI9gnt2kZ
XBSOz+HEifDI1SYrq+cJGRyf4FK91Xcra5ElI9bU1MrG3ksEkAi510ytnlMfqWqz
YgPF8xBSEhV4/UX0uFqval0pQZMtz99/ooMV8LGxLI13YSDggozGCXNfdHWjds1F
SjxHWF2jDwNufWf5KyMBZHvE8646/v7mBulVxH4FQYja4bceWNbwQGXCpwRfAiy5
xBBZS9UhI+PKCD2bgG+KE6DpFt0zzoVKW5WAyEcqGMPqidzruVfEDxniquUdgyin
JIMSqpxJsxMxb9S/EbckISQjufhWC5D0jSc1WZHmljD3snBkfncgSIlz96d8wyqC
2eeV9yCncLgohlqHRH7oeS4aoVGGR4oP51wwLKE0TJ+GG7AHb+xxLP7q7itzRIZv
l0bS/cwsCxn+3UbGidFtG0olDfDx/OAeUfPLuPYdM6F2US3fFWM56+dKeoFfFxPK
iUJBcWR6zr9+HFVjANBPTsQJqOrmtiH6fE8v+d+gsKYCFyn+fJEzI+CFbvGBuUn3
HQrBPVLL9DkG8TW8LZkDhhs7pUgCHG661PLa7tjJAAodTpx1NRZIRRaiCVZbtnyH
XJU9UFxnbrmfZmgTpBIkUnEBQ266vhYVD48Q+FawdgbaIkwm6x4Lv0SI66XtYcEv
NIOevpRJpmhoLiw1elNkBp+pFYhqCHNF4JORtxmaaUE0KErfjMbh6iGXlZdpLsAi
kyjAA2Y06Kh4vu7mm0RhRVkhd5T6zqGuIb+WUiREZR2B42JEDyjPFo6NJqSRwNEC
2pnqLzjDTzIteLZ8mphkzbAWpCR6AGA+aR4Rd8sYXKdDT8dEGj51v6DToUOy9wp1
/h1xMSPoqG9xtOrzLnbrZqTl1h0K0xCyQW9D2VdY1+Z4rSYkr6WX4kdZqKgK/vtg
TtFPaRk17D7hNIJSHENnISOJ6rWJedfBdbY2facqW7ZOvSKZmTI5SI7je3jIRuO/
MVDuL8FmdedOgwpM5JNUBvyuQFvSO24RWskfJe5DuECZ8nSGjjdg8vBxffQpgO+b
d8XKuS8pKrStnHZcMu1GIhdcZrrXDoEUk2ASPB++w5xAOCVWf5zX8Y8erorGiDJL
G5Oqr3tlYyG2yc3sXntm2HR/tlzJdoqr3O9NYxygW/keizHEX0vl7IQkW4sSTdOy
oU79TCNm1OEh9ZlZKnguINAZ6XLflj3RJ/mGLZ8eW1o27RDq7J16veJdtsidScb2
ITZbf0T3MFuLLSuvnLlSmf55VUdTy/wWo9EA4yGjHv27baAM0j5QHnk0AFPffbXf
CC6X12/f+x9+AZdc8qlwg5taHZrJm6lKA2htyGZMeDmm1UDdsE+NRChz1/kMGH95
0c5Q8r9eHFdja98NDuRhVg7Xmeo6jBKLVOiQVXli4HwAdgT+L3Ein8+qAI/M3VZ6
E5aunhUx9W9yW8zEwXcfvDE0t9ZT9eN5rRvld897IVs1ReoVnE/xy77MeOmrufR2
NXgi4RB+pvOVCOkTzPdbnqqaIYAFWCCOvk3S/IrSQuT9fQqAwqtEKGIu2wlb7F/f
0BcDDCyS5LjICSOoDACxPvfJnHSI/Sod2gHAZa8NDtYF0J9Yl5KsHKNO/xktBT2P
/3599Si9bsNy3UlBiLJdkjoWuXQFzOfH/DsNKCWBgTgEt16wQ4Vw1xB0yzlYmlXl
+yxYeYgovKYKALVD2CGn9gL3j79Ai4ZpxF80Ar64VDFD4+pig59+4WQzcymiS3dN
Of6F7RzZHAWGwqS8AWWFO9CO1FXZ4ttlgbcbsE/aOv2pCi0gQs5Wauvz8nokki5u
uxtdRn5aBAezoIQPAwUdxZgQWKqDKsSU5qEKgRwwhlpHg48JjDuky1rwAplNPO2h
oE9Lw+5tmYpWklBa4Gqb6CcSgWmmpF7+WWDN3j31zpfg5I4Gky0hmp3U4JMG/EQG
1KB3lGLtsUAOx2xt/Kyh6MVmRxbbMjIH3KHqoTuYCwIRrBiQQq0VcuPK/b3LilGi
rO46e/Ed0Ie2FD4Lu6gOSY7ikV6yRqEYyvHb94HgzWflbdpHVHq0kgwu4QgwaJ0b
/upJ21Djb1x271Kk2b01j3dy8sGz0oGg9D7uRUshRmJiMPbmbYrviKHgltVTgvoS
mdgj8xXLfUU+N7psP4q83cQ0qIRFZl0FyWSogW7CWiSCNlD7yDwtz5Xf0VI5OvFA
N+s/1fB/JU2/BBTQa2neIEg05bulW46F+ClvFqZoemRhnzng0AHLCUqpkIgG7EHK
GRnQjejbrtxM0/xEC9n7NI8WGF2BUdRq4Cs+FLLw7HzVp7gQmvdI1uQsG5icq3JO
UaTjTBzOG4wmRA90kGQ+sq5c/WNF3hbvQhMWJTly21ugV9kjUPftwkTkfjOw4xLN
lqAkMxQdTaLoWcm/hobnB3NFXllClxDOOVv6oO8CjJBvP9v0yBDuAen8a7+psFlq
/BojzXrX+Qxdqe9IAlik9lHv5zOAqwg8cDxWYGD0VR7FCLEJLyYgjY6KEcQxiHXM
7AQuNjt/CeQDQTvQE/CDeV/l6uYTgvI4q3Nwy5fOZ2ANRGKNtCgDwUDw8BMBodgm
epXOjDEYHN69qIwdStpbsgEE/huSSu5/klfDz2f0fvRLujx2F3xKgG2skia5szR9
F+Vn3wmMpc9kiYugO7OizmvmZXT5L8AN9NCMert8i3x4SYuhQPp21T1kGiD4h+Bh
CldaS8Gl6KFAH4WsOAsrxOhUQaaOycELIfgn+Mf0+rU1iq0+5gv4Jghu1Y2E/L2O
v9UpAcFsCxu7KWww+HCmk0YNkI86t4ta2I5ngEjAVVHYPWb4nXYj8+Siy7xAvZB2
bVLNi/YwWva0XcqJLHGQd6IeGv7azXId0uaktb7ujtwN31IsY+sE2ev3kUqa3M7J
QbucKphsR/2Ghy731M0WFvKcFUV+pLU9Vq60xsvG4aftldzjxwJLKlJVRFQbFOnt
dLdD4OgYPNWhotIRgFM5BWLdAxnNhYcj5VQgpfIBsE+YOdzILWx4n3t3EZEkw8oL
2jS91X974NlBzVbyr9IBnJCqA8mdMaXLmhJJVqKduubpayY/9LNdbUZbGxt8/0qD
A2YZp3VMN1DcAbhkGQCVwaF4y6r7q8DgaEdxg8YmXVajZ5jd7mHYbm4/Nb4EgeQQ
sZTaxhDslRGl3Zh5IoiDuhTT2jgaGX7uCT8xHn05XzwaUPIXgcUADBPFpqgsOYNT
mjD0jqJn+WC5w38ovXDYfvmZ+P/pTi4bmJYlkFW1+Pq+jiXYe9NAlrkeYnRvrFCY
IAIHj22i5Kv1UPg2lPSoFov3kGJI4rbuesBen6mbYBuaji7sDQi3uzyCIkGjx/d+
ZKVsD23EgCpDIBVUWJ1tDFGvEUFX/QY9jC2DRNbnalBytpjwozh14uehATuuCXKZ
X/K27G4OjeqACZettf1LQ6hJJqGrb1rhzC4X8nZljvlXl38SNNH5wo5Ef8fhg66w
lLLWkbvYas9ifKcw6uGn0SUVaev1rxfi3Q99tnBqAGZba7Zd4/fBQA1ayO2vtOtv
jbf0LkaUhZSZozMqsWhXZ6oJYXzDbwl6krgiI2Jw2LIrdZ3t2w0vjqmSoFhWtmh2
hHPmSe/EfhxXiVXBJsqM7E30TYJmOcSjeK773qYFFgdYt6mxqTo47OBSaeHumjc9
rkzlGj3KcQSEfhPFtzXn/dr5eZNAK2+pz8Wx59hDPt/vi6B+SY7AEzQEyv/RoOGi
uYhbEztH8mBei6CqDkOPbMu9eb5T3KgQDhUUuZWdUDsIeeTOAizPeRXO/jVCi1Bt
RZbAljaOXAlVVxLiHwmwjNBpAx8a/YUQIfcxdZu44qCfylke1VSCQa6bd6V5WaEP
03AGGnA7ilnPSzswCa+j1K52bXQpfa2fvFYU306pIXgiPdk0BP8zIaWKGJa8sNRV
1cHb1S0SlD+aYrgSpNTNv06KvGJkND/ZrP0ZUBqT50ccO9Plz9DaNzb1cpNa3zQw
U2J7St1ehgt/SQVf61NMR0/Ps0MV0cmH46z3uqbltx9DQhgGv9279XimbbvTlorI
3uJUzaSOAMkbizbBfjojzOFSB3UoLiNFl9AsOuNMPxoMdRIHWL/X3q/V41TzaVkG
hAhXLWWRlNOQo7xc7v/+dBq74DlD3hG90A5ZBp7ges+LtRoKLaX/TUSXYRsM03JS
EglZ/6YcWYi66kv3Uj8PpYbPSQGINY5eU+0NGM03Dv99/mTqNFrS5v6XjCEvSpZk
Pz1FyCsD9p0Y6c59Kr/xVppGwd1F4haYvQ86bxI7Zbbo+F5XnQ8VjkrflGFb4xsp
GDeAVnNyoptrd3KTm1/d8ue9EDt8vCnQT6dNncSh8ChFxaY+Y3ksOq7iGlH/risU
nA2NOAG+C9WKer/MWfzDJNallwgka9t2AIcyuSUtFDoJRKcjw6dZYa12QmVcORO+
2Pqq6ksyT265qntjcI+4PuykPQiWxdHs4vwdUFsRXh3R2T6+zVPmPlRjr7UdJQmO
FxFq70pyp1j1Erky08xsE809QpHYuWTRQPF6HNQRvcZxLgTxOTJgjrVufnQ0QDC1
GHDnnrMjm6mkbhoyKivQqrN671JYBdW8HFYl3+wT61paJ3BacAb+AsNPR+vUaBTz
PidKJd65HZQF+QbMsC1A5TEwE7U5IwdxJ49TFAedaPE41oFUbZMLIZQdVP4o/FUh
jmXmkf7YTqsApmhuqs/ghbEOngmYe2Q8yGem9PZDLuoxIWoCjZ2Tz96S+X4tzfDB
3g93E/BlZ62fCQsfDbkLm79fLA4Q6NYiySYMwEqC9BwQz5h9byyTt96ZZrgQRDPA
mwgxRjjKtHrSlbiLn78APTcBBiW8l8QD9JdFROXdaukcQFZ8VNAqeYDbn6FK6USg
i7sJsJ7vqc465kThif4fBw5UTnHrVEIQ1Gh34Z+LBsL14lN0X4QjML/rMZS4rgPU
YhE+4qG9mCc+nvt9JYrpz3Za3RLmtgVMDh2Bo+/dpZR8rwhwX0gqyfxs4rt/6U8U
kfqHgpJFa95AMWCjWIb1+mCAAJ1klfqEIDiGS+MYhNpkQgi7HD/eUXpWVoJiGB4u
Unfh/SpPjAFkCZpb0NmrZKaKhLwYZ2sKXvziPMJgtHyl9T3DyDx1sk3AEUqspn0g
xs3h6XpMHtCNRvs/z8q6AdpWo7J6Hk9U7FxcIP7M9lhXDdu8UUahfEHtNpScmtGp
TNzskyA3t2B1Q/QKBWEMcNOikbaNjofipagFBB8EvheM4I0PHKXVLoc45OKyPSSM
d7i34ip53EIU/KjDcI9rekNWMhAVhZUUGS004UX4V3zZ+o7TbvTp3BITYD79qgmn
m+Tuu3Mu6shx4uizJhqI3uFu1VV8Q9JfAA5M+d7NX3rVTQPbFdQevf6vOOHcMgNW
mdvPeJyJtXAr8x+MTm5IEzSVV4o8lJi8IQpfUUuoTahntgLsaBqRFE6AIOwWzVVF
CrIaEZhHlmd+arFHfn2/LAmfGBtbho3nW4HcmivMmzcqRCbCL1xClPDKR3yEGTvz
Zv+Ay6ehXw+6MvIdRff0qp6B6wkM6fFhqzHE6E4XQ217+rCH0b0ktKXiNayzwylp
JAp+BC7Z066StBoNV4M6usfmec7H2KaehsW1XVUj9F57SQ7+SjFNj77CRIHbGII9
23t2JKe/wz4hRe1+hydtQActTWO+Gf8am+Sy0ohmV2GMiLenPPY3VeYo/3UBgFQk
nOBp+RVWFl5na0MBDGW6jrOF4fymbIBkujaww7dZKzea9frjRFkyoFFMy9FIYtwt
bRCa66hA3flulsfmV9GABtacVZfA5QXZ4sSZxtm7eRxbblk3TsDENlSElxDa+Hx9
ZcK3tuk+78odM0EgH9X6NOWW+8SQ/0/LrmpfcrnD2rAS/kUF0yarq4GE+ANolNgQ
/ynFFOSEzA3WaEay+9U/f1qJoj5c2NenIaCjgSz4djJaIoMndrfdcEOKYnvxGaCh
nR8llMI93n8u2xOkhFBIJ8dhyd4eW2tYd/NN/d6W36gfQyJ9bSotsLXMQt/0gztk
oK9xY1+hpgbz0h8SCgnsHEi4PsX/Oh3mVNoPO5xCOhpEXd3whzfKTlj7f3a1/HdP
3udhO+1HzRsI6RRc/ylp1TGdn6Tb+CHK05rxW7OZOOJkVQ88APonipnZ9JhYeMSs
lYT/nbsfH7m3Kv7Xka8avKEYZyGyNGitmBAGKV3aKJ9IOMmcAptGnhOvD9wEUzW/
2u7Hn3En9dC4dwSDBmxn5lS3hpXEvf3Y63JE6JbdGvxOu9MBLgjlIeTFMoxwTp3x
RyEjy0OB6JkGScjzf9K+yq76zRFRpRvxfthgozUwcXNXTkYfovuDF0c64qswdu7O
rdq4BYy1QKuJEVmVmXswj8qb0WwKoTvdfCpUEmaNUxFrfaUTKwEM6kAU6wPgfsUF
bByAwPIJHXgRoc++wQk4kYSDw7lQkp3n3D/iHG1/tpoCYzjAbg5sjc+byTsnwW2c
QkDuwM2hlKKSjQSXmm/na8xYHbOWw/z1JBqDmS0+iG2eEwdbtBQ1s2f+j+IoXce6
i7yNanaI3pjq6dALuLaE7Ghlas+CVCssJMxRqc/eiZAOxYwBsPwYYyL4wFW6AtVR
7f9RS+Kxngr9oHtEkbU8jBRB0hEnPuDuoB+gTnPiGDcda4MkGbKnKJLME/vI0xTv
pSXjEPRWbmrdOvy2g5BmrEHE12Y1EkXVCGdLkjMgBC6IyYT4KXBvqstDE+fMKD94
pMgXb/0lYZagAKQ4mPBVmpPcNMX++BcjSkxevY9d2UDkzJe6KF6lfXItvXFEPXQy
Ra398ueEic+LHBk+fLh9O6mJ1EoRflqmklj4wS+HKekyaK1TcN6xponpj/n/hHN0
ILuUP2cp0S0VsPqOJKcY3e6UQ3E5IshoeuDioD9ZWQ5AcgJhAakCOTuJeDWFz/0B
Oa+/3SSBmFsBxVTBJXLUxgOoW9o8hYlIGYeSTVGzOIyCgt0HhKwnQ0w0KQq+HvyT
94TQo1ni5Z4PqPG/7sF1iltSvJ/oqaXLe3CReUBW1Ve1/ecMRepuHFG5cb/Qg7m9
EDJlEbwr800/grzyT522Puzn9xdRw7XhlT8xYQW7EPZnjNrfudYkyew3HKu1BNCO
OtoESqlsJLBSNnUwRF6WZO+qaMuwXWBMHUA9QH1pH/BBizmVcTesU77qxyfQkFgr
khvdvKFptSulDBxGOPWKzBzoP/f69y9+Iif2HURaCX0pVrz4uPrpDQxtGd1QFQyk
EBmYUfU52RdBbcqfWgocOpY0rA/uxj/BVChb6ASWq3kUHrljxK1FLRzKclOGFgVX
TWT27ji2JszhgPzpkBZtROC/wMf3KA/mHnaBXJkqF1daI2waVoIQjAzAYzqG0wE/
ubRYu+nvaC3qyl3Jv11W7MYiGBdjAJk7sLedk6+mHqKjRZWCaHa6tCIkcEHRabgs
RQyIgnm0JdCLevYJhj8IhubxD7QAzzvvP4fRw4YI6e/JxuwcirDG2pIzknlKvtLL
mcQeuTPTmYs+N9Tms6t4BONLsEX4MG2tKK+JPo51Zi2RdmvGuTQBBU59AK+PcYTa
jj/riLMzJBJYBnBcw0ityDLoz68txB3pScHmaaV4vFXn1ENTOS5V5c9x0w6Uw/Rr
tFBG4E5uX4uhsnsSHFLcrfNCfsGub7vN1F3aJeWGy3FKBuaGgEkbK1JXAXgKlnH1
rneS6U+K6OxoI5jII247FR7QXdy/TFY+9OaV593+O63kDy/2rajIplciWTDfkOkY
crpmUcIf4Mutg/E4W6qWLqlA6yAyCMCvOvQ29LTWXXE+Aayoye5RJPIgzBWDVqYa
C4kmz3Wod+mWrAhiP2z8oGQ7/pOY+C72Od8AipEU+6HzGVh+CzlxjibtDhtLco0M
u3tyKy5Oq3GImJ8okzUwJ7ca58cL0/nZa4VtoQvKZuU+3p9Dm2UnZVjgHpV45uY7
oSvjrSuf7WQbXsDE5B8IaNcqfgbgdoFibsxL6iKIdHRD1Favz0s6y0dj/SJTlxBf
HRXSK1iP1lNsWVWTNGauOI1QC+6bUSI510c1rcHO93rr+7LMKAFuAIgWJ8QzfTN1
fmxqeQhzqyJvlD3dOrW9R7TnZhnUYucAXp375CCIzvEVVZWCVkcNLFLqJ6O7YEox
+PJzblwJ3sfnhyVUCoNRDrGgwlCppXbfCXPSCTZrCDS0qmDSDp2gnVq2Te1CSphl
Si11aikWiFH+Yq7TJyzaQLfBIsRLH42r5p/A0iHTdYdPPRP+GJgAbDrH9Y49Psqv
OsGBD9zeb9IBNDgGZ/RneF87bIg+EGPbqyLjnnGy2f1HkpzZiQP53lJVBrLUSYT2
MjO9Xug+acsJrHcX1HabhHjutoy56sBp2XkUvdXjKOdgz0wuzsaZtKfcqncP/eUK
20fxm6HSlFz5KsHRSKPzYZqExS0J16dxbXHsGEoDWsk0t5d5aojkgd+94SpeOkb4
Mtfnca5YTR2kLsnzyEan/+3OCRG1uGv3LvThdW4ji7Lp95ct651nCmddj6y70CeB
UWAmuc4HN1u/HakY+aSJXMN2MSsPU7B6tFHPnCQ/+Cyj32/6Ss7oecqWjJb/gzjB
qBcG8QpYEf/OBU20VX4lDM6/hpnbzn2f2LPDVmnkWUZGsnmEftNu5EUQTQhNyP0c
w3bHkQ5NvlrR8MPsmoWZLJq/uvnleB2Y7vIDJO6KkJRO1aLEF9+XoErhkUWpKFjP
o7CsW15xTwRiQb7ynm0A9oGUk4oeDqhw+oxqaPNzMreHLanJv90f21RvHR5vOFA4
BkaWYVBGxTY3y2NRafARLo1RYoA/M0rZ9d+1O12i2ATjluRmixQuzqU15KWhsrTZ
SuVj239aD1Z+85hSozvvWU2DVcfIl6gyqX5Xoys5BSi1sgmKjnDSTpwsmrHS/KLp
YVfbOZp+bGhR5j4wTt71oFlIblBikmppL2k6RuEtRh6f81Daapq+gCdbX+MpAo+6
t2VtgR5TJaHzNd+pnIGKZaALKL95+cUUmvXqXAOk7QcQUqFhuWLQirqtsMAmchKi
NyJ5eKX6bxflaRlkfA5nKxwdZLBhwPTmha9dONE6q/95kQfgegRWeH0Vd0yADGVA
4TaSIxm2FuD8n4T+zPBDYAll7vDLBWlT1D8xQx1t9zgQ2zSmSUc/AmJ4aPeQDLRz
cYxTO7epWbpoEypv4HHS2Az6sLsM0IEQ2Rmglzt7PaWOKy7nWhLpwfcBWJehHCKw
lg7ejZPZUg83bKOLr4Yu8Vvp46jqs5m5IKcjpuTJh09Y+61ML66+sxP/pBqhroc7
9WK9rhH8xIciVVq1FjSk7JjKqycPJLc7Qxx9wb4lyvSWEbmExp3pcyGy3F5VrMYh
gWanIJdipXfO0cFEXn9kUx0xUCYS/ojdOKf2xMgzbI8FNSWo75Qb24qMyylguPjV
SXLfr/06dhJ2rHN3m/VVufEsM43GYZ7P4ubcYlvSOAz2/up8x0A8xB/NpsgLXOis
DmIwUiqkNfVEbbrqXVYsfuq5pkY44ULY8EEfWTHnyblPmlzo1B8X6bcniREbwrsF
LbNgetVguKgiebWnHcfQKDbTqKDvU8LauIuktU1IF9N/mFHdyR21Vvzf2HeoqDkD
Ti20C2rVJTA0k2zn16r8KcPAB2yVmTqzKbt8KzQYR+jTgNmxnojT7zYuxtG4ph/v
bua+Pgulb1kK8qYxtCuJr8hmOJXDORw+Eh5jB7vQCGMTMTGVOb4Rb+vPPp8QeqFw
JXkv1cgQ+1p7+ZSI0jgOi67NnOiA/o3elc0uwvky9AHTDGas4ty83EzJzgVUrMqp
HDK24GXJYD63yII5UQ3G8eoNbnecxY9FZJg1RTVm51zgUMS2YCBfNBXl118UEwWI
vKS8gJyTCxJqaN6Ch3Z+2QIrkrB9uwfeB3B9gtUtHBs2mm0zHaxKeTPL7b8rkKl+
D8I5xQbBVMl86yS5xQ4gGGtPg3CrpNEs+TNoIUPqCx0GlTGSb0GecnwfGzLmOV0C
fUFhm5vmyT+ae00FJ535XkweWHlU5MDg5bORYKoJSHA3HxbdBOWKLn7PRPf6RzK3
PkQSVzFf9HnkAb97wJs//BVCBhbkzapDpTwhU6XhI/wn8yiGwgQHaKyWR+eKAtjc
lbonpkn1cMUg/dziZ6qh2y+6dW44X3LEr8U3voS1uLmbiQQcSZ42inWhnf0ybSi3
AxbHvBkZv+mGR09riNC4X1JR9lqZh0Qfsk/bfpgRbLZcFPXEESn0ucViU2dYfmK2
rEZiDIxiFZIPD4msJhBXPf2MuykldSIvCZcQd26VuhdCejlKn8G/7Y4befV+MLD6
dF5qp2fceIWx1H1zTryXVACJXuOXbqf/ciWvxN8pkBfOHGjohXbB8nmRg2h+NP1z
RJ07LEcL5GKS4BThRhZKUj5k0S07WmtMTs/dQqZO0nBSKXMK57IaKtsWEVXC7aCl
D6Ua1TrIGQn0dQsLGNU2AaDytoR2H5lcfURLgSddNOjjNV+Tn9azX1TfGkE9V8gg
oH6qSJYHwpwDxKtaoLLt5kKjtFzNblsAHmPDH/4Mn58GKRY3asdMrjlEtno19e+/
Ehqno6PO8LcKpIgjQzgQiptuS1mrZeNCgpx6aJ/2A8y2u2rJHeawxeCDyxnJcEh1
WWhNTsWO8YNezxHzCvKTBwqEdlVg6vSDY+sw1cp0Ad0g5bedSLZOlS1DXHbWw2qR
vTJ8/K9Q7lMC5PLhTn7Nyyq9Hs7bQLbA6rL9qyU5XZkVPYaAB/tl9y3jUvN5owFy
C7jCw/mI+Nf+ZyTMleL+tQsfD1vX3huSfJn9lJL9WAEGxnuW3shPJPaB35EwTlPa
VoV2OlgpnnDcLK2xfaJPd7bSlik2PBRx9y0XqvBFZQFp1oQ+aMTmRFQP+ZPfx6ku
a58Pj29QQcFICv3Pq2jt/6uTz/KrA3cXT764Y9r4NXuvChPPLMVUOBJXzvZA3d3v
yGdSKlIkyTXsoLfvwFYROCEfaEvv1PaTnBp19KfgUp+VOa+KQbWoZXVXAJzclU9a
oeKjuJqppgdhZDlm55jlgEFfhhGp5/ZP4aOwwUNM9ujrhkY0NwSnZwF7KFrMxa8p
xC7fgVDhDXJEe1LZiDdPSd49rNzeVGEZ10IgH4N+2UxB1UJlTeKfzbDjxU43xnN/
suOFpQBjS2nGDODQPChQvuWaPxUEUwbcTPoOsLKBMcsEpyBGNlPP1qI6m5u4FWv+
zhY1DRaP41Xujc5+QkbV3TFh7i9RrLvSB3+vlcVo/Ce/G8u+sixlW7HzfHqbvflo
1b5/sy5RXcbVO8xbevvCcMeuXkdtrjLOlYkBeWisDH4KNcqlywUHBS/paIodC2m0
54+ZmAOQrBPlkTZKgw2uYHIlF/twDi2rfKnkx3M8wAk6YJjnu2wzhuBP8N68m3UP
4VFQ6EQYuiMV3SkJX4vPxmrNOXtWZynSl715jEh+hdopXIQHWyAPi+p/0wgRV2EI
J9KuefZUY4vUtRKSvMe02E7Hwr/ITkgle7evOEylkbkSHo8bVMFi3/5eKe8ydgfa
RwwobwpMaImlQ4CiSYhwlAaf1ZVyp4xA5DP5z4vJG2y8zqDha337vrlqqxgz4MSf
R8npaTPfB5nbHdH93aZzbcB/1Ob50ut473xuRI2Wf3RMYu38e6mr0eTeOQJlCm+Q
VaRaDMyzsT3zRPyWZKOPCTgOi8bVV+rkE5crlZvzw94N6PoOO7lQEJSYmc084nSc
oVp2CUDliQcChmmB5EOxDkyUjqUUnhEHhjjgUNc7rd9f0Krk+sWjmD1HWGCM7GY+
1cnwvSk+XIVR+pPKIqFtFFWuYnM0OccnNaBkYzqskfDL58FjfqQGK7Nt+GV72W79
ww2j6jWHk0Yyqal4I4q6RbaVjAZTujOJzYe4v2Us6+73fw7AlyZJVOXyHK8pU1Ao
5EAJZM4+uDShZNQAT9zm2aJ1WcR34o0sqqR69q31t7bbLn6UQtfICRaNl33L79Da
y1mKZ3gkVI+JKgxaAiuPd+P1dj9+3BLfAszgQQlzkJZtSGr+euK2TyXvINsPdmHM
I+hXsXcOjdgmBoLh2OHtEmAXimHSYGkQfey6/LhbE2o9Gkwgqoq4ILuPsBnTRpIx
7N/B4dyuH4WnW5ZnRFf/5oqO+mpJHKTZ1VLXwViygV+623lUI2XrKuXo9JccvBKa
6ea2NAAnNALETs9nXaHxBwXLj+4kCDJezHiLr7VeBaU1xlDl/yzKRtTPHDy0+Nai
8vbzzqIJpQlOMNuDxsTBWOr3t8SJ23q0cd7m9qhfoeJnCt8leKoIIo7Nvi3AE6PG
VTRvnl3W+uqIHID+TVaqelJiw9CvZBFGi9dPd5rajfar0klIbfdk+Q55txS8lxif
OImOp74fexaD7rjKrMHsFIxrhbC+9GZrGFb6Mx5VrDheSug7X+M2E3Ksb946dXEO
S0f00OUz5h/RG4sE9mCDmvRYV36rXVgmoX2reVGJ+P/OxMGR8/Ywjk2gvP0fdt6k
KTA+63rKvXKbEDHmikNKd20L4kCsnOs2repb7y9BEprJd9Q2hfHzfd0crbMn0F6w
07h37u3sVpeb7PzrS6hbGeJbSsQp5Pv4CWVZWPRunUriNmeNTKtBtGWkp3EZKNwQ
V97mqN7bkfbariYFfry3yvePZAezbM3yw784tK7lxJjdjMm2MKMlUsGTtiYqYUtk
HZJU+IcwJd31AtHeyiQM8uEV/bDStVMhr5a/RAyGZhrm1vExAbp77uYb3stA3k5v
PQT289MAMPOkk5r0l1HwzpjthvBwkQLTK4mf3jqdZqQ1HcoiPW5CLiW40WTakd0t
yWdm+YhEx6sXunrG60VTqkgGfvTvv4EIw+u2p6lBEiFkJedhKLk4NjePl4fsXK/K
LC/SGgSG0xbfd/FQ2C6YYupFW5IzUltjSZ4JHKIX0ZDNgagQ7z6dxBjy0lRGlzIy
NPpv3OHkpxEhzJvg9SJsJnausT7as21uDv7GRcrG9XcLhzNGRB2dZ0TNn1dNsQFP
vJcwFmEf+LUt2jW9R2s1wBBDzPT6fgUjrjQ5plicLckBaMO7RSb+4uMp9zaqiSRQ
PjliRyy9rxF/AU0NDnfo1laCEFtEdqI6bQcrlo++e/oUIvfIHpGYquUITN4KolDO
k0Q4AuEWmXjpr1lZ6pB17MaKtWuDN1aHAIelHG9Dbn9VdcJImhJt/YRtpyGSZmof
OYgPEkK2RFULTQvC+v2yJMoVrcaNLHEPAy7hCv5vzffG8D1l8FV8v7s+Nk1sfkJZ
CxHf3x/X0Ce9JKbkrJQlYFNfaNEufGBT1Qazl5HPbKhKKgXwS9T4D1PLg7S0/b1/
UMkfuH146ig12ewo3mlryeVRSNstb5rRXfTUusSkhX6qI3kBx8I4aLuwraNBxIew
VF4NxZVLr2duS0ViQRs7fPPyl4mHNSflKCp2rMY/lLto1XacnHsjHYVM22Yayu5q
IJMkw02uiVbsPwExs/ZxYE1sk7V+I6r5SgSMPbEIoFsIj7KM2mTGn+LdzZEboJ47
Qtu6H3UwB4kDN4kW3iYN1gJz2lAlMgM034SxFMcDkY1Yhr/Ol447x0L376oX8PeE
6E8haJkrhOsxmWQikbNBvCvnyFNPeID06oKnrG53XjLP0/gKS/Gvt/k/2UCbQMLP
rO8aiL0mQtFn7U2vIupU5qENg8mU/VWpeS6ehzyoL5RTCnoyjCWzxRO01lBfNb1q
L8fvRU8/1V+yKifOgJKQW5RO6VbHKY0zTC50dxRn2lc145M8g082MvjJ+ANe1a/2
ZTYbsMJJT8dqE/YPApl6+Z+LCIat5b+qabC5R5Mbmnru8kaKI8M+ZODkSy/mJdZX
waY1rVkvIQ0LgQSertUFMeeRBwhVTa14TB2rauMQvweCDSK2696nM/OEdzU58Rai
+w3qXAKpIDLAQSoyemV0E3uXVhtodm5s83F5oWaFabs/RZDHLkqdVf2yZiG/QEk/
8BM+rgx3Ya8/qs5PJdUAw6sHVV/VZiM7KBWxq/xoCGQLfIlbltVm1Vqk3yW4hLAq
dWfNbQqRu9DXIeazht9pBtfwKlY6pLSIzfxhO1VXQtYJylfBC5vCK68Gucjmi0Gb
pvSLy7vlCy24VrnSG/KehfVKrujzko5QrDuv+6Q91NxpQuIrcUx5Y2ZfaZy9w02u
DtHBjwbLbCCy1l7lT5C5hEbPO31nf/7NFL9d07wuhe6ZbaIFXzixwrcNPgtv+yVn
zGS3gmol7Y/wx8pbHvL3faycQrf7e8PPilMGGmW+5Fb/LS7ibOSIG24yC+iZB+Xe
z/xFU1s2MUpVGYvTxqZR3UlCYJpb3fZ71x9SRrR63P0H3TvsJvZvQTuFnAgTaMQo
BUgKtxXST/E/ExOtiop58tLVHGfkCnxmE5kETe4wqknNeo6WhWF4LujUVTcKhS6m
Myr9ZbGtD1o2ZEkorVfFXt6XwpOROnRBDUdEwNJ1cvcrhoWoYvSSh4JKGUnsFd6t
1aOQJYZo/dZFvP4nlNU8FSeDBeU3otT/DNUhazdM5Nt8GjwZ70m4aaOqbj2glGaD
cVJXV4pdkSh3GedEqelbSXEf6MFYZRBMMxgzeXY3eVSZsBCE6wEaTizxadb9MdJ9
Jz6WFA3SLQcxkfZk9XqCYlrjDN8XlUU50Ifc/MEOHiaI7TjzHawgxCUkbbb2z6Bm
rCq24nSA5AnhHg66e5snKW9NFqzisQFmAlHa2xoao1XpJAJsP9bHZUmaMydc/bUz
s2X3f7xiNmGJIJFmyQagSnDddpF87rDtCaxGYW+QP3uXivaTIqmvPgO9gGfVj3mm
xT1X+No1a9w8ifhLK+0SpXqfFwTXErCRMcYh7h0EyvICZ9N6b8XQ+BpIkquc3SS6
RUb3bqrHDXpyG7dFRbIEUx8PPRPpcxWkUgTl8Nn42RaqWGSFMLQWdsJ2KzAksI/e
HW9hy7NIiJ86nRuOkLWai4H/pVu+9s1J8dxiSSHBL9GswuYQ7Z5WLEX59Jxdf4UG
gTvrLm3fcYogFdXbmVH1teJwXtLlWobTlIEObfHNFJTpPc3NOJ9G0oAW55zYTbQr
1Q2x55j09SFoo7QDGIAxr+oYrwWbot0lfMnksFVGYNNbmKa/BIZE8NgLXQS2DOOK
ncf91tRC/w8Wx+JTr6zIEGi1b5B3G0W9ObwBbx8a+V72LFDicA/05zsQ+dcK/NDT
WlqI/IKldvydQ7jQSz3Qy7mjdGnifteRgqGXdJZHCKtKc12hv2bIONoghAnvA94y
SSPJvJciFREjjiW+b3seqU8SDFRsQj0uLWU9NkLR54DoJ7diaz4TBbbDvR6b9KB3
JFqO7/75X4BDPRFwFxonej0JoUPqEFMKRZnQ/tKqvQub3cIfMc6BvI6ozbiI5nNI
a4UYk6XRXMCC70GTnUH20bYxrK12MkhTou4EcQp31qzI/WTo1hrRQdqNShsjNk2I
p/OguM7+ZzDSiQS2LSaQBTjYEl28GTY8T1RqBWrlkvgaT8P8XLYyZ5npQcS2z/Cl
Ud+f/W9wYh4PYOOPh4FE/4ue+JlgkeAtLCPpQDiWg5FWpIiSaKxH28ZrRPyD0Wji
Vy2sZQMWR/KiP5J/PLz6vPJlqeDe8Z6pKNEf2Q+IF+4Pw+fRxZF1N4B0ctQo3KhH
DVealJAsM3yjvnJY+6dbppbXM4pkH2G6CZg4bD1brIA40espT+iztqa47UrrVPqh
ZZVmVvZHSkqYKsxX1yOdJ8BQogChHnQB5qbGecmrfJv7h13PlhjzN0xttNveamFa
pFQ/lFI3+FR66ppN9AqhbFG7bI1HfKKpWdaNLwBRWDHDyq8W0zTAIfhbA9IHQunn
Bd78okG3FUZGssElTYuULGrq2mSk0jsmJglixrtjrM7LC6Qcu3/0DlJjtBt/649A
pXz5qflpIGnOI2mYB53KM87rxBhF6CeoK0LLeOLl+QmzmVaE9Magle4txJdJvycE
vdmLdBsnRdc3J8+aHhEJPQt5cQhCeX1xt4yYd1d/m2/mDZQYhF8hTNnLO1cKXIPf
cpiqfrIqwrmURLLH2sRZTWbIALYZLBTA8dknS6Emgi2BuR8X049+ZSE6Xyn/+lz8
vOYIEBguXAmbmMsXC4NmsuEo3YfFFTaNsheX4DfXSvaDibM7E+mRpNsyxnQDvYQT
bjfzSspWVnRYO41/lPeZ+3+WwKXbwvnhU8axOU/M3Om7AC8k/c+8cThjxVWTnISF
gd+zgUC5gNfJYBwL2+jRapTmOIY/9nIlUIv1V/bwb3pippafbY95nOD68/VfjGFc
JMsD/aZUIn2J77rbFDspel5N5FcjZ4yTnLW4bW/IG0Fac48BChWRupLqga0+1QTh
XJ4BD4pat2SWGXSCBuhB00bYl0xFDow7vRSu7b+znBMKLQdQiPv1IENG8RKFD3bR
ruzczLwr7h1r8vrr27tsnIBxtO8pbZ2CHkyBmtk+Dxv86zzjA3kuXXRK/luKs7K2
5HErYHySWk8zC7/pa11X+oARaG8mszm/5p9PRU7UBDmHcEZqk8EKykXYGIeERmkq
FTzvnNsgsES7MBLgQO7ZLJaHu6Q/wWSijVUZ2d3/uoeu86qx4+Sr4z/jLWEJjuO1
mfKD8LZQ3RAZh9rOm4zFZHOWAZe+voOyh6+e7xymP6S8EF2H7yRwMomt7bD0lBSA
avjFQkNOeN19dCbBbZr9UvSB6uWRQPSHR7LDOQvZKkceEFMUV7NKmkmRX/9LCfbB
k6hVzpSIDbss9cdamelBcq1LdyqJhB+iI49xKzmHSpiLq/09Kp29IA4DNx/caHl7
LdiuoE3ZvKTP7vp9K7XHU9hRdZH3bi1NAd98MT6uCPH60I2B8XdXpFD794SFROeq
pXWP30va1o6Ccfrj/g8aaphPAwA9kE0F+tt6GEXxrcXe/4OdFeyNHJke14pV4rFl
OJoqAyZVg8kYLmtXYfKLn1lwHVM1sOqJamy+cScU+vfFMev+4GmTdYOMR1KwkM9n
u3dzIQZFUgPA7h2o2WaVsJIVxZQx1MzHppBj+Oh8202vWUxbwWJ4jvmAFfslUPSE
Mr3vq2ZWI4gpSXetr4UtuGB6RDP7K+j8jEucj/HFby3vStEWiCHc7bPZ5fGIV9Rc
ZId8CCyAzW9eDieaA7TuDeS0bPIeQNRjjmseRmEem6JL1pMUg9fknO8Yi7ZT0kmb
JWqDK+krwLbXDT4Mc6SX44wpk7BE/tHjp/esJ2XLFzoXkkV5v+sCcEnxQ84zROti
t8qcSVm8ytSq6Ud+xcxWDCISTTWShNAbMuvzhMMA5za/I0MJgWrHdPPHQCziWTD8
sOPFcnCviDliqwSLjavUc2LnvwYOIGeNWiwtlXguB91gATIeT6VKt8JBk48LnHbf
bAuv59eayFqHfzdP5/paOeibbsnmZblUS9pS+9F2uT2tYxYbMU5Kqmxya6Igc0zY
uLrtwKI0JDUl8g6TwWitBt13Nr9fNTOLsofZ8p61YetA0jU/yenWTPzxIK+wALvo
q0ftFA1NXdobfHy5CFcmISvv78b4GNBT2KUoKweJL7krPOPheVUixf6SZQMz38pk
8Ljp0ElelnyN6jq+CDxlxYL5AqXDGxTJMQoouL8sEBaW3rxRDuqlC753eofTnUOf
GtmALoZPM9QqPTQhEM6fEjmYGcrxj5ZRLH1f7q8COM8puNH30KnkB7q14DWJKzmW
7KpkxB37rsld3z+q/IIURA+Srd9vSALx0b7InWFXox6pxAKjUTk5MQAFPSDrbWq0
BXbfMe86MTJ/is7+k5XvkpLZqXo0dfdsBMSzUq8ZuwF4o6DgUpj8QsmFNlMLvEdt
Djvyz7KM4Mzx2P1SaVfjK+S8CEM87yfmJwRSOkk83Hm99/Cs2HsYy7trSfQLXRIg
w0ONSfUOn1VPlDQErjzfghr4OgjYKI/+2un/t2xtrCARde5BOc7Wud0dviUh+ua8
Kev/Ar7412cOK+LuWAoBWG3J+iRCYXJH2poZ3X+6ETWywwtvX6mJWTaKI0Y1y7is
O7jwbRzWCzfV4RJDMyVQqAC3Ajtf5T6DPbBY9Ml1Vcy6GBjG83S94mAAbYQ26hIN
5yI2UAe8kcoqTIH5TScGKf3/vqF3//8x7/vG7kD4NqclWwOrreVYdDQA70Dz9QWL
x8E3NNDk68KKoq9soJf5ztOEkuIIWlJkFJmnwGLBdgHyWgQXE1tM9nPYm4NC0kLR
OvKATCGk2bEnLmq2IkanfpLdykhMmN5HeXE5IOOAJ2PSBvjA84uEFDaacHX3lsT8
xEFP+Agaz04jRKF/9VfnxW64E5a+vlV9xg4+runz3v8x/+45B7hbuUxkbSEpnvrs
y9La9WcoIEYK2gPN3TQ/qB67BqodiH7s7HhuXTOGPSUnQMs+8SxYNCrYDGD0WIvp
hh2OLf6yqhWySXXHGeVZ9KebPdaYhJAr1ARA9t+jWk8hvVRnHrK2jQ178qwJysF6
hi1TbgiAwkiTdOgBAkssmC+P2act4jx3ZF21pqA3YJ6WXShL7SPNWNrAWjij1/qa
ayO8dA6yx922liz/kVfLdnidNkNhc0ogqmZ2FsBtekyrHA0iDj5/x3vVeSP4WR2+
z8ulmHz4d6DH3KGvs4m4FQ9gM0WihVi0V5L8tiFhe2CBPT6Et45ZaubskyLdWKwp
/Ymp49P+6VcKxOaJdQey+5hgPTs9R8cA7GQvCVpMtlm2mCcQvOwpin9IR2XkP8Ls
53iRKkHKMWJGc24yp1znRKTbRmYNvAt7cbYmWbk4+Qzk7Dw2Rb96RERD1F+hT4M5
ltlPW/9cAvjE0MvJaEDCG3gHN84iCxzVYt539fe1ijpXvT9nGDU2obyhA+TLaKIf
zEF1g/jMt0Sj3C1ly84t3yTOm8vWAVFJQqPJA86fB/7AZkXfHa5qlHuH9JFF6Z6f
Dz59Cl7bEEmDgLJthsezK2YuWYTsm6gtcfCGWRnUGwpTtA9pugc9+7qJ1drTAggv
iREjAMWbng8bc1YGSQpY3Tw+ICRHxAHr4yFjzbqzMBoM1KAyYY4HgtR/MfUxHWBz
q4Y85/xdvMhmaHeMno9R5XA/S0+FeVOw6Sl7fsftzcDyoER1RpBIQGvGzwxZ5olx
LJojuXlwHRGJlUv44CM1tmvLnR/CDk+eohraM0OQxFL8/T/lDMKiH64ZtQCTU8Ra
sXQ8uPLTRuMIUMFwKWubTuHq4QBhuOtUTDd0Y/qwio2JB6BOTTEuwhB7/1E+N0Sh
hywW93D43/umowPWgTogIOm7rtPg/lOZfq+tLIFPZm6lsUsjGxF9agsb9f0ZjDwO
UzR9Cz2wy+G6EuGLVJDO+o6ygPl7ii20wR+11oHmF1nYmUO9M3rSHw0pAmuhA0CW
WfBtKTM4J64Vr+ko8q7EPR9ONdx6Bu/6qZcpkzEcLOwOx9ji4plQytL8WvJihtsb
I9KOmj8ItB6mSOQiDjyUiQQihXdCZduYViE3/8X7QxU9k1HDe5vn4WfrH0MCe0l4
PMCvw4x5ae+WjZgWCyyGVPTwuX4gcNvbQUin1dGwaKYLV4jo/4A/jyMS7TmhyjTt
iQf4btappmbf2uuc/E9aqBkwBwT00vwFDv+LR+jixbtp4uotCwwCWVdXULOQfrEo
Tor0TiBw49dk9KZRRksRIrjBgIprzQQn1J8qMP12vFv4jMgCTwR9uR15m6EIJNnT
8jIeRHykKGwgv82bvsyvgHUOcqeRVrkLGrs3PC7363/ZmLXlYzAcu/p+gQ9PPI3L
jnYBnoj+QdPtfN81ig+OixitWsIzEsaBt2bSoVihhDE0hA85jD4g8F93DpQbVygm
lfg+Q31XXllKeIFJBSc0uccBvOcXSQ2kYDnL76A0Bh4isR6U90KHwr1s0dTpcFja
a4s2HkwdSdqpMb4W5L8175Vuu2vtR4K5XzoEGLVZYNadf55aDnGgbMUoq33sMYJc
oSWuPihKDORc1ppNIeRe3owpbqO8BWhjc0P9kCMTD+m2Z4K4OSSXq3OGlLZ+Rc4P
R1ji2i2VzOTYnTObrnvKZ/CyrksirkqS2h4BsnKi/mSGv0aHY2X9iSW1zxiNem+0
fgP4iJkyE20Dl9yEdaSYwVUsuFzze4MSvz/LmNGerGA0QC3zw9RjoixnN5z9BpZF
ITNq2awoPK0TBALFL/HAiCChtELQZlTC66Q4k2MOl/SLDaem8Z/K85sjPiHBXMUg
RkhpGY83VPjmhli87wPMi8HZ2wUs+xUhHrFgsjt34A3Z5kEm8SN8MUuLO80Tmtik
QAe7+I51cXEUkCpY9gn++UnEagYq21v/u3+020EDNLo+iTqt/p2adIO3RoUAd736
kureFXeRgy2Rcqt5yOaVngDm/wH84d1aTcqFyP/fk71jrleEBTDOS6QeHTNW2jeo
rvgl8KhNx04rR1L7w2Mq6cBFigY+bgYY0pQ8StAYgiKje+HIWaZ5Wwx8MmSqK11i
hNRDLZJWc8pPLtiDEQIlBIZl/K9u9e8m05rM8tr4uvXBcfbwwowr74RR/Y29QUMq
Pfvg7ybqyu6kb8US/yMQY13vCwsP2U0ax/uszFmWZIEouDYTfx5r4WrPGs1WIeb0
M2yIddaeFJbuyP/6BAlZpG6LNt2tA7cR7BLEeqjY4wb1aMzdCfgBHmhE2BoOsMG4
dIYeVpBSocigLYIPTtCzVhJIMcHowl4GBk5+R1t/iPZPKT5xhyfXP8fFw0dTr0g/
pxKJlADf2CwFVVomIDvIIGsHdyEb/KBGmkkggxvNpK3xbNx0msrMuzuSOZxma0Xu
5fwSWSmZZFVMoc17DNbD9/LSUB1IDX53Que1pBGcKdD3cgXSQYF0RJHXChFRF9m9
t8+KvUsrWZeYU9BWhShb05O8APAYSq7qsjtN87ccEaE2BCF6h5G1KUBvNRkdCory
CNgxCyqzTRqT/9n19j/2CdnggmV3AilUK9pAJWX+YwWX9Kqty1mcZVya+mKfeNuU
4eRQ8lSvg/KZX92wl/dVcyEMFSPAWg5rtkI5PcVkLLFJ1MKS+3TnwtuP9S8gU1sD
HDYq1kWCrX4kSGuhyytWFOoQByHhar/7i5oHs9XHj/zrI8yXWwvaTLyON0oPInfU
U9I9NoAnndp+vsfS5AGrMQlpuhit1MTeYjIHowxdMhgO5ob5/QGb9R82XBhRABaA
SkpZot2GfQ7QSDf5Zq1JBwhu1MmsUIgMpClz1gR7dotMgRFs4jEWiZLPEgW4NWU4
DQ/CtTAqaMdn/oAhxN2VGDc9TyYfFqn/OuCyqjJoCdKkpInPi2WyzhN0oNgsN/d8
1/80ykQ7cX8HEr2uARlVA73UL45EXfZoNiUAGWtZmbORPcC1bIk36D7tMwSr5sOC
pkE55mKO0w3qhdXjz3HhwytRIu3vB2VbqvhAwxLC/yrXYpzspx3R5LSKvYxOXcPL
qg7PWzEXzYh8FAG1HJh9XRu63Y75Qkf5ClKSjAUjoSJC0nejvxGxde2LXttbdrUm
ADnHcHnBSs6XKUbiYMFh1sz8Z+LJg4mKCxoJ+w4cHjTZQPTbaj4ox5HfnZ78KcOP
UDT6i3mN2GVtofrqLizLBRk0dEdoab4u708Tm21y6hdTn2qKfPj1SnjSYWqFbkhl
1DOtYBcyc4pQnFevD21wvQFy01C0aKPv09O/A8zJ7tmriwXpXVZXcX8+YbADcbh/
H2S6N+2UdwFyItNmp3XJvIS+z67NC54072bqB2+yhiaYAVDd6pMNoCW16QN3orsA
H3WW+tedyop3K/s9uu1hfXzfd+bWnxBP6yw5wkxRKa/j8LhanOojv3LUjoRrJdst
riFqWJyeF/ICMExNcVG4gQKMg4iYKJN4a/0Ng/1poVCMBvGUe9hOldXopkpkAINC
IfL0NEnaZ1Cxll4oN6VohFzSA1Fnh/SQMepGRw/IrgV4Kg30muV4a6pB+f5dzzkl
80p2jzd0KCC4JH1Fx2oIPAeNIstqn6USKmxR9qzYasALx7OiWnJUQctYqkRmxZN0
7qJ3fn7b9ajm4HDWZgXIFuqNCoECuNgDD25a14VJWNGlQ6LR2m0eX+aRK4oey84p
6St111keUuMGUSIJ40+WAOjJPO/dR0x63YGpOX9FyRdhVCdCp3/OMR7RJ4H3We0m
gf0etud4LCnYkyXjXO8NgpnaoVo9FLY7wOefM5SkKc7x+DW9ybj5UgPyPCjSEjc4
akeyBIA6gdPRnG0xwvdkV36CtTQMbTojqKIP3Pz69Rv3BwP1ks5Mo1kh4DJY/w4o
+7BbbxPyaoN6pavcCJIqC1ZgKzSYiDVJgEJVD1PvG+7eKWcwNouvQF5G2mIA5lxX
4S4D3dWJJRtmCepSDu5xZahvBR2LI5XvHtMEWsiaRjzk4mUILFwHNewlIfbcGMib
QykiyXhp7CyXaSyeLlTol9ZDLKwo8gt4K5Ky6Gqpj1OYfXZZz7T/nVYgg2XoDNiR
HOXjbBDWdo37XQUFcBhVeePfbRTMgg44bGgx1RBBNkY2OYsKqtuMZ9GA5Gm9eSZ7
Kh05pv+SB4W3X9BtoqnJiiW41+Px+exAXkQGrQR1rVQxT4OZCFcWMkvYbCCIUe7c
PNaL+9hZ3av3mifZd+Hed3yzTSU0ZrDrjSbh2kCRy1BIKSqrxCHQVIWuYAV/WAyA
yKsxmcA8SRS0C8dneLa9BBMAxtXUvUKKdigaze/diiOP421CnkHTzV60FhI9yc6m
j3wtn9V1HE81auOVTd0xZfk0YaqTeJ2onMLW+jp6riSaHvQQTgRJysN8tOp9eQQv
nvqv01V708x9d1CqLAgwIM+wgF+GeYHrA1xGs9qmV3DAVbCiDNaH++vSOHXcZmGT
my4el9ugdXOeRxD469QJLIXv9S0OF58Ng6v2n9sLX9fT1+iQW4tHJF9ej6J/0VMh
8DkeT7yzx8ZzBmu77p0nmjvH+YITW3Ye6EN7CjpeF6+2LUZJMBBDD61YiGKIetbV
6cnXvlRaqDAIp+Ipstf+C5ZE/UUz97alMqicDRTlzlUOfol+MEJ1Zex70J47yV8H
raPLrSmFRWXLhVyuEmfrUkFG0s2zRMCHT7psU5ZRnCpvxAnv6N5igS+tlq2xwSq9
hRYlldqzlISNtfHEqMlFKiwnVY00TqDvuDsLa7KfKe6KNDB2q1uVNrubjMeoesIf
o2Qj9n9frxvG/tKVH/VXJtRE29pTmSgErUIObfEwOii3IHOUvBgE+F9IBrSalwLW
UqrtrBZ5n0O1zkE/BSN5c23YGVJO87LbTnXgfGsbm/+GPvDFXHnEGq6ORL7muZtM
nWISLhk51VBT/MaENLuLqndC4MilmhsNbPukFtei48BOqb4ZrfNdnVQUvdTJGjf/
Cit33QiCPyLq2gzUc9IRw6toR45vNtajQvQNZjOfNz4LhrX+n1cRy3AcVcuS7M4c
Va3DDOhDZsQnvtLxUKML9vw51ZweqKFVwt2rVgnX1JZTsC2tfRErZr+QSmGWJzSC
pgjhwz/ufLQyCPA951P0kPLQSFDqns6shPmTmHOzr8nR4XkzEXWcMlEBpHSRtbe0
JWfjCK1P3LKuMlrZkNN2I1fTHRUCs3gxXzftfyey+4d8t8Wd9esXogS3nOQfv6yw
KwtSwj2pNpExD8a1Q3IxSV+/+9IwAlSRjFPIURj2YYEeeREeNxTKcHmwnpUch24j
CamrRRbe95LpoZMP2jiD7Id8+DGB8Er/b54jQe6mVSqobi6WyHLS0RhsAIDnKlSm
aN7B8muQOGnngPp+yJZuoPQ0JXh2l3aqMvvG7O9fyYhixzbRvINh+8UkP7ECyw/F
embhE4q9bPo+6ek7hcJjE38biBRw+dqtnMVI/tOWGLFu9Q/Y6UddE/wXGx11nLiB
rtjTA0L4e7OlcH4+4yy61u/oo+1eFj4FqieY+c7gYJ2i5c0q+HpUfn6jxGLkASVs
mr3eibkuKHMICuis82Dpi/t8pkTKP1YA0cKyqkSfbhvavmQ+Q7P9ZWi5UGww9RLc
feECcFCkjVpqm6NJSqOXIgMfazrg72tlb056aYlIH2/NIQU0msL1I9JAN428I1DE
IddeGbkVCuwuRNe0cuPrWfQ8h1nvEE+HVgeuD4mH22u1EEjfjpG4uv/NRXNSWCfz
txX7k33RTRKUpi8P9dd5tms47lV/KPQt/PTNphJk+D82x4OBZSy1CgQ1/YS+4LmV
/hg7rpT0CQQy9TtU0vUovcMZwYhp/gUMFK0/mJXCpJGVQ6oNpjDZHEsRAIyrd/q4
oRd7XB6cLFgECfSFLpxmDXa7hPo7D67v+DHB97T/lynAeZ1QZApodXkXsVbF9SAo
TLZErhII+DF/7sCp0KbZz0iqyKwSl1GiyvOFr5GN3NMWkffZ7WHmtB2R4CgfJTx9
2WdRDAudd8X6CMEfSvyHwxJC16dwytjmoNFRbWynYUfbhxhLKgXTpcETqO2tAgPJ
k5u8NbiV1UUrkJSuFC9bwdmMGUBWhwFrh3iPsDx01Hgdtiuzk95bBUUlq+opcPhr
STg1mXYD0trL/zGAf39SKspTfek8JOEvFfasCVqty2kmYQKc9M551SMGy9IZ8hqy
z/kjKmLnu48Qno6syqsEAHTFj2odN6MZsitxmzHVDNOTxgvCFYAvAIDZYA7Zm3+H
P5WxT7SL6DrCV26FsmpdK8+/BzyDrWtdS5cZR0LqUUXRTIiDjv9UvOC6Ir30GuqK
fGsy+ky4G63yiiq0fPNiB3AxKLiru8X6qqJc5Pjid16jjIkS6yOeJo0865LgtB05
0MvODNHb7vFARu0lsnsuDQH8ctgXmtapzJVXlMiR0pihRR20C7uPJ/LEI+zCm/mV
4fiKplbM/aNbNXWhZxVB1IU+kkxoFlkE/3bD9fMUe0Pag5dr9FUog0F1CL46xSK1
sJcBopyMlnN3RwTVYriJ/TH4PHFLOMQZef1D5R5jjUJlXnfkGTjiRiVvTl932Wzb
NU40ZCqTEyww1iZA5eKb9eKNJsuzlgL4JnKJEUaHfO2P8RzXvVy8Lerg80U5i7ZA
Q52QPEYI3sLdwgKtBtyNlzGLfawWrhI5wGyZm4JhNjcaXH3Qi/iW6bwK5WKHrsSH
QjLZWDJKdppFOtKoEYV0jlvIciC38EdZHSo+oS9RkSKypc3LZKyXCxjFeAsEqJXh
StMqzfkiVqFpuNoh6XFiJcfic8mdqv5j4vJ/ZJTXu4jLxTpDHCg8BoFH4TiH4NxE
BF00BQ1XShrKBdzmvlKTW6/bxurJ6DBKsV0kJj9BLxhGTABu1FNS5RBiAUod5H/C
FnUl/1Rwn5cebf99E6uUrlIQy6NeCCI2HeNiIoREDnCPfagWJD3Z6IyQ7ixGkzG3
V377TdAtTS0z7I1v+JAGkWoqBjX1ZixiytWCTBZcptvJdNka1iYjDiKBSy5vLzG5
NwtgX7dZbEn361qrfBLh2/o5SnrA89BDT3hrfadu9Jv3lLgzqxxL9eU1t0Mo8iew
OPDOjLHTm+rnZWmPlXtj7oZmC5cu4w3dajgf8oz2i+P+/NXmHRw4psj/XBeSCnVj
6Ug818Cb6J6A7f/6iCfhJ+CAToYp9qxvw4mjFPy4HP6PRC9GhUdQMR9P//xDV+LS
vTjZet1hcnH6/f+gE0cq1PHxtIWCMiFbdeKEFSe+09556XJaqD4p9xEl8lyZe0I6
EbHGJCo56veo8ZHNcKmlMqU6j7YGRWxCe1mScQEelANmtfxRK4n98B95DT1W5LP7
Fy1Ih+CyvXNVkYT0tdWK/yHb59gx89LO7j4Yv9xLjK2P1437fwsHO6udLI8Sd1DK
KbLAio677wpc+kvYkMFqI7g2am+FIaAChKnFv4/p41GsaeReqJmrdZzDA2dLbBlp
YPvrYTNFXEEs52JDi/Gx6Apm5GAi6pi7L0XZVp1i8kj9mjOaP0K1z78FOW5eMAk4
Sr5bH3CsI5PkOu8+DSoSHqv6aneHXXM7ZHyfDpEZvdN5KN4qgY2n1km5ZuFsZpWn
sWZo13w3mC+8hlDLjkFKqcSIqr2XMYJB9Y6kw5PS83EhQWAAi9zDHNWwVNphHzvo
Yy43pqZCc2YXRstnrr8/qaUpunBDOF7N4Bcsqqm6pZBr74YgP2IXvEDfgXXVBPVF
syHLh7czXHukzfcE/nLr4lTM8n/LfABxX+W8fa0h4amzPjsfsH421VeKMz13E/jw
ujOj30I/kKSmpwnsfF1MMIuxbMG5usAVHX60Ui9Wf3kqbniGP1MI85pXD3JQdLPV
18IRSenB0jd0Gvg0ZQYJrxrI2B5adaMq9y/rZSbO6O1alNKQxHqJjQDfZc6Bjoym
9RgbiMePhasrVQI8T4JoJ+T5/ZU7leTNfqvaetj7OdaCJJrIFV7K51bIoCknm2yZ
OzE9y2WrQW9RrEH+8wNTewwZuyCbPQzXfFzpwCF1z6DYdT3UVfrvcqxWiEGocQpH
Fw/rXxUXIQCS9JBTN6PT9JAvXvTiakyuIbfOCpGagVVQv6r8+F3BXNeFP3gRPg65
2W6DrEi9ye2257dKSH5qQECybpAe5Bj9K77ms565sedfQX++4hAF3nv+1iVNMK9A
FGpZ4TpLORRsIKGqbfjDRTohQFUjXYOHHTzlZB8r150VjuXgsoIyy06Bf7InjAH6
1dHTlAhYU/o3Pd6R3YqovkWYPDMc+yo0tg6ZrmVNKSm/IslWMP3Iq+VNWP0l8zJD
zLM5U6ouARy29BYjmgGdwMbmAuvKYCogoAo9/dn8V3amPcJmTPg0HwNAAMRgoLUH
6H8Q6O7I+miSWPusfmcBJRtgv29R70zDKh4gsfPzusYozO7gWNQcFvT1MSG8pIv5
JUfgUof45gOIaFfvVbVIFGxz3wyK0k4iwGUsQ+k07WWvvRTy1mM7l/IIQnpr1Mjw
CP5OGeM9EXYm9Iea9+GVOBgsHLfWF/6mfLGtcLaTDEkQOnGcN5gvTw+yEz1NTdFF
RzHlaUtNotyMNKwVAdJLby/xYUJFw7dJFkO0KKeJSWdQ7OlvrJoWQX6ua6zmF6jL
/5lfaZdVVKVjW0ccEB4mP/+a3p+jqiP5+PAfVTlmGAQY404NTDjDR+gMLu7GASjr
IsN5UnmkeGQUGGX2wjLnlicoga2XLtA9dwLr+QiJ+c74kgBm8LjRYp4PGTm2iHti
6ZmlWaEJRcqHa355q7u8mRLcGdVm233KYvCOQcOABwJ3LPu+Af3LWi/C0mjg8q/W
LjkWSiCNPWomZxR6YQO/RNL4faninjdLKP48dFpR3GEBApoTR8879vaWITe0kAiq
S6VpQBXuDd/bSTTba4hH75RfNhTIND5G65gthnsmq5moh8/pqwpDHUCHJBojTIav
5CIkODHzvNDs6q73Wrnr/xi1b8S3LKoWZ0SdfYqiMhSzt8btNXe+KNQ8VQ+P/TXJ
1ROcEgu7DZmqN+ikikkuxxQgYyW8A67JTDbRud5KuZhd4wEItK3tUNH5S3CYzgdv
uK3xQkyy9iwhNTPwO7LQR6I79aLe1dinF4rDSjsYWek2QwG4BpG4C6Zetp03QS7a
LZl7IFWekT+OIUPFTXXlRYjurElEUrkv9UMUuz1/w4oLPdyD/IgevoiR7XhlhY/2
yFZMULq3L15WRiKy3G7WqLr7o+dhxrmP3w8WZfRclfgr2QbNMt3oa0FM0U2fH0C3
GKYk2Nbek0bvG0zN/7JJnY4+EM4gBwgGmmQQWEh8Ks0g10okSh22w3cSRKRVmHYC
Y/t3ji9XUYG7vdyMbRMxVRVvyOViNF7yVqEZfX9nzKvi4laH49NTjpefycgVgM77
x2DTcmprBjQzmmF6qNi3h24+jrmZK+Kb1tST/swX1a8ebArcMAPccoOJLehqdrl4
g8PTDZRwypfxR8UqdU3A6NE93TaxX3osCTvKpvL73bJDeQkbNv5opUzK+iVTJSqY
pTF7e1zN7+g0G1TKz2CQafPvWo4QI3O8J+ES1wulZ67EPyYAN4b8XNzvoIScLCYF
5hprIHWlkE7WyicUk7G9gpoZSf6jKN859M9Ysed2+0RFNo7SS8Mnp5ZdGkjRavDU
GEmVDMzahXPTjhWSS66rsspJAMtdblmUQt3tJmuIsArZ2G/WUBjwihmOijFKBRcw
ozikPOuWOxkVjtbHegnUhKgoQFkGH0F75bJIgBiEyKSiAPGdHUgbnPrAIqN7WGFw
ellzivDcds2AhQqESu2hVw5T16wDpU4SOfODBuQBOvPaTjdVjXvUGVsC3U+Bi9o9
3QTjMWebl14ISU3/e/2MUDzbY10+CU82mf0A/SRJo3nfnHp8V6eW+bt8E77j65TR
2O2rKwKxsUZohOBw4PD8pJqAHfBRHfLy6RmatXJup3CbErZ8q+PJXjrx9EsXnpB1
ykHnDN7zoriT1Y/h8D3q+ILWOV7e9kts0kr70ERsUtp6b6eQDS//1mtsxrnx2RXK
Z9Qsuf4Ka+cQqnMob04xP1m/+AjVqMnSESoo59emhqfffAlrIHdRCfTn47/GjWNS
zP+wEyB6lq7SqZu917qx204oTMJMdbmvv9xKrr24hggN1RtwfC+0mDCXzSSOMfmQ
hWW129M2vaq1AhHF1CETZweGGlLKJi0E1lMpVOEZQ+Dg2W8InNwJRZNcWVX2zJYn
LHdcLFpJhmXYNWl+2BEsBzGDdwNUcPk97tfmPKlf0J3I+ubhaPe7t74N8wB/mb7P
BtVuBCEz4AzXVsUFdVhLd29NIw/XBjmo+5Fm9zJKhhz72/JOSQ56lZRiEvou931p
AJPlnSj7Gi4FR2g2jgjLxpeCZaZ6YSX1wYz8s/2MAjHxoNr3BiSi/Q39kfgfyuA9
0YvhTU5991yuNs9PLrfY1ALisgGNVII4vCQvwERYwd0Q+0kog8iQ0hxUx4A0etlD
+sLAtjOXvRkCp9N6/JeJh4fjemt2wvh11h2tA3UcSVQ5ZtNtlcq/r1BLfcbtmEzi
Uq930rE6PFEPfMfkpZEEXuBKEQS1sXvQtBYl0Y0Jabkkgyk+4ZKzg3QlXd7/dydu
WcjJGamnQv/DMnzKXtcrKci4fGwwMvLO5oMJPk6R0Ggz5MsYH0n1EKvLkXfGTP+3
LUn+zV8ly33yAOWAReZlEatpYdsgpqS2rutxpWp82RUj2Bz4u/CCasS7l4SQWye+
sBPwSo5azKrdqF1DOcgY3YPuVVC0nBdqT0WwWebugtsM0H6Rf04I3svaaBP45KGV
lAfq0K3eEUeAW/+w/YFG1Og5RavpGH0WyXf4h1BTkeoDpXFsAQpO/C0ddGsUyhrB
VuDdmtVfGc5XWCgUAaE0sRlHPGHr0yTq0e2TTUbydtnilFgub/Cj7qDGJwTr8Oo4
cORMTAOnYuuJHiR0fbdr5zfsqnZsBOX6vWrVbDspONoC/f1B8gqLztl1gvKzAdyb
s27yqwEFY7Zv5a+EqjkroaQsSPYlUESpacVX/k1hcOXl3LX9E9SQW+UEGvJypPsa
hCaOVaqvup873nPKlgTsf1tcP2/DUu4+psRyvZ5VIUAvWpq9BtH9LvftBya1pPAv
Rj4sHiOTYusnRtt4778QoE+V1yiWM8fjl907MI6yKqQufk61K9uyqT2KvR/rhe3V
5etCm5DugC3KDDWJmnVunlFWctKzoo8alXW0B5STGaT3tZKpbMflquamevWzql4x
GfulOE+iHwSzHKRPkRxVAxxkA/vFAe0XkGJDSPoD+magkoR3quFyspaRFQCNsFfP
92oGTAoeniZqnRh6CDO85vUw5Ic8t41wHrYE30Q5hgoymHq7guL3CXUmMKHW+NUg
JPVeK80hHDtjOwKGrMqT6RMJRrfabApkkQAbNqJqmHAlNpK1lRB1gSsklvLpZG/Z
eaDbGml4BclLaRcZKEwHc0almrc7IlClOSrOFEtNw9wbkYVUYJDUaHlpWi+5LBUR
YIQl600uj8y7VVXapBh2BBF0ufx6T2kNBF1vRU/hkCzegaAfMIHCS4NWWZjAYUk7
QuxX3+vYM9/DFnZx6FAPGfKHIg0u7Qp8xsADjvOfLuSrJJSJAl1067tJAfPtjNgh
qYj/bzeS/i4q2ACIwk/Daw/kzcdFPKZKOhbjA2rGQCrjSClC66Gg11pzvPNh5Fmw
YFnLWOronJj2YgsNX1fhs7/LSNv7UGniRZrfkj9iYls1+2Nsx0KN9S1Q6W8CHPRv
RRao9zdHJwYK2PMw+EP9w3SmbgNr5dduHLvbTRLfMhrM14wz41qjRwJOwXgQoTSH
qOB+uP1fBqxNSS3IiCTIEPlA0bsHdknvx+MQPp/Cm0bHp0tWhSjS38ntGkMuTgqL
dmn9km/Z9/sPO46W3JXG5V37zo8L0RFSeUGUhjEVn8exCe0OEleXo7Kag3DMiRix
mBcAe61zXXqEKBK2Mslj2tuRHPinWaIv7zlzbyUNa4xiV06uSS4khEvUdBPYqXJY
DT3nOQBIBUvKJYqKN/cb+SMvTjUlnhtZS6bhW/STq2z6tGDYshwlkoNpkTN4RZmE
eFJ3zohHPxBob/TZXCx+flhaYMEuJo8boGy5ipR0EuXpVYVCU6MEsSzQ5aXppA6l
XAKfSPyKKH+/kdL8jW0CYCcuv/nCi3YAVaXszxPVf4jIXjwT9afURwDb3B7r8LoV
mEj5Q6vYZKbGT+4EZTCrSCxfCdzgDe+HxXCZPiYtgjSWZxmdC4WacgasHuqfdh0d
o/X71/ifiXCsDVC1gLqJ+4Fa1j4NWX3W1FmoAZssCPFFWWwdjHJu6wW3rw6WTIAa
QXTDWO8XTF8Eaq6mjctTq8VvTUHeXK/dZN7VQfueZ/AJ3d+EVsnbVtawuG7dTnrP
cPZPISNP9MizqMhqn8/EPCjUgpA9kMMz23gjA9uZlTxlYG1LXrmPpIReqw/RaCJy
TVxwRp/WCHLu7/pLidHFgVhaOUbt5pTQXpa1/DqCCdS2cjTg5yySz0pLJO4oLYpF
RJFtaXd3OV2mxp0dC6qZ2KKkDD1P9rxjYUZj78PhNrNwSfrsi4Oxh9JWQF0JTZDA
QBLBeKijKqIsi+WRsvlHTa77ztfc8nCGbj7GfNj0R4nHhq6dLu0lHN/BnMCg7/jM
n6k+JRmH+1o7o5kn3qcCMBK34FTgOl6PDz9jCg8wVT/5BS4WqyJIuuakg+e9N56i
HfPpuTpMn6/EERfnu/k/AxD1vQGrjdcKyIhPOXwxgnftZGOC18IXdy5PT8Za28WJ
Pn1UPqfW1YegO0Vt9ZmQ5odiXlJQSK0HeECZVxgnlzOC1w4DEQiTNPTK+uJPrenU
W6A2EZErEYAZpsWKdGp8nCIXGsIWMk6TKoAlmLEtKhYSqia3ClNC2JnRs0cf1a9e
L1Tlf/fc9IBYQ1kc3zBf8GuGzomleQQWZk6ofPJ0ak9yCs/eYox5eun5KjzYaaxe
c+Y1TkNXrGSpmAY8ZWgULXm8SbwP3TOkM8UyDTBhnmgkZP+lKRJF6aiN84JXLYOA
ZX2QtiPTNNNaLoP5c1xQPg8k7tV4Tt8pxBSQHF8UBv8NE7Yrs9ZO01/MIBrZRJAx
pUPsvCWvY7a22MGn9Mlwopwqn5eoztucS9OwIRm7vh9aLtJjxVTxcnDzyA1QSPNy
dx6s5aSvguRYmDFCJwp9UxYgQhl6Y3hFruUAcyYZVy+ZPd3a4dXtDf9IIOfVFtvd
dTyrl/n0vwlDPe2yLjrNpQgtEx2zcSdyuRGPCN5Z41z3BqGqXH0zPFPB6HfLCpFE
EZSIhkPPCFr9pONVLoijTG/9EcwA08MxchNH7edtcWD+1v46GbDeseQVAfuJqv2T
HmkYU8bC0DocoUCHFjq3t05N3Yy+mXw01DmPmAol9dsgPlBmIp+AkIOISX9g53Pk
BJviMPXmiR2bU7iiE48Vbeqn6LkuyLXQzK+UfvPZdWLzhaA7PQxATgV/U8hwBEHm
jmzzddgYqOWepMPQ3EweN5OgalNAooFyLRaYQyyxakYQDiX95wH6vWRbc/6c/Cy5
VOxOumGYOi+Jhjx7gOVrVY+bm/HZYLXFVKHU7R3IJPVWt7Pm1Wo0Qg5v0RQz+In3
t12mvqT6whhvfbhC+AB5giTvJrbr4c89zpMJQQYh6lZ90VnVDHQbcnW10pene/Ke
ZBfTXmZxoegXxeDXho/Uc/nq4UCjdJ7LZpgcabCcSV/tOffhpmLfzd11TpCXdxPt
NYdM1kYZZZ/nnX/c0qtdnThdP5kzTY8lKqv/aJ99V7sedW4ICXOYDcm7eEXIvifx
ZHUbHrPC6jYyYxr1e3dvjN+ENsvJfKeBnZenbMn7uhouoFbxhc6KCGYfhmBuO0JV
ZAnYzE0VzFulBgo+NrnYIencVVsPqhVJrrW6UVMyjCC8Hv+xiMlZylyiBCYLIa/f
YIgXXutDxamWYpTkHUTHvDbb00YG3p1U0y6d7ZGgrv6XNPjFfW2Vfvw/5HgWCBB3
fT1Kn4XBh8O2uAA7Y46Begefv4zxS80tBTZhrQ3Y62/FLVM6IP14Xe1Uj0EwGVDN
29Y7wP8eOq71zI8DUgK/rrpgboUkEIhzQRFMPYMcxQq1qxh3PrsbiKeNYrUr6OAc
fH0a4ju70xJ9KsZIXrDQtUULRW3ELRyJ6SSWYeBJF6j/gpfCTBdFjh4ZbxW/4ve6
nlOBvD5YYRcNR2pHCSBdPq/8+dERcqgg1yf4mue2utXW/h5QeyLwPF6XWJuAQ6DK
TOIGetThg6n7xtUWAsaqd9J9EEARzxm2H/avz8Gql67vAbjNZ1cVw4AJM0m7dAsg
HLdVysmcLI+4LCm9qTysA4JovKqkHEjncExTflZsBrRFOtMDF1PNkwJgq0sL2j2S
mJM8HQ9t4SoV8JO1CgatUbii+XTDxoxLIuRA9lnPjpG3zmUzM9bMQMa6vIUGtP0V
3MCfDW7LWNA7Td6afqnyCXm2prMMPEBxgrbQ6K4JpJRHQn19vHL9mbeK7ohC9J2K
9c3yfWZzvKj1JcWi3+Elrpc3X9kvQQ04MOEJkYTqBiLJ2RjicENE95JkswEwNh0/
iQKgHdT5D3phAnzBv2xQFickBULikuFsGNQ3GUinv3EsPkYGtJQSeDvpEz9Cu9Mo
8260QwNhoCJb/LzNeZRGThIaf4qbpKshV6ArSbRMrDPKDJzd3tRjWYX+7G0HH1Uw
+/+olxXgJr42HHjoWHi9OgHOa+7X8VnGEucvAryXd8J4JjW8Hr98hLGtUKQWmCrx
doMsxxmXX2D9hM1HcrBnO01lT9rFtHMliuHz2vhAbX8w1xD9RtGnc1frpxHG6CpK
JVpJOV2WiLAjb7VVlj/rUB8sv6FXTsDaw59XF4pWEJyiWoqo/gZwLPtPgBasvXzy
dOyt1UmtPlURKjKkoY+mcyNdS5h4YADArCAJtulAHKWq436vMtBIDQ02sjYvssge
FKEVADbgYIjxiJ0HAYky9hbBh87T7XAyOszxOrh9CFT9TSXEN5MoK5kpnUF8AUoX
/KsqeOlzy+73+MeVRAWipW+64Q1O/GElsdSWlD4eUpVeattnorsM0kxA3WuAsbGQ
4pBrkiTOUwKAYTPk7bdj9X3H4TD9myKC59sqrPd+vCQUvFZk13lM44cTJEuBSgR/
UXvP9X+7TIRHJCUz6cjRzzrDlhIzInEZMl5h/nvpmuXpP6HiW2kR+XnRUvAHPWDD
9GYo/oaoflEu2tXKZtMCHw5jJlawHRbBXaPA7CTezdHLCh8Un54QJlMfKLRSJzZk
FgoknJHLr361gDnHdDbTARvP/HpfUOmJ6cqfJQr85vM3x+zA1SqAQlrA2MARO9sh
nj8EaHqw2FFDirCQDFiGNYJSkXgfSf8K9tAayQFS7bvoA27XmpWyg+fIObYDiY+w
5EjRxVQyAhdvFMYnuU+jNRAoWXcIBG35dZwr4YFElpAuFNdLSB4BUJO59SOmsAD/
5Cz69EBZQXE24CDt7dhgCYu2U7EjN86qN4N50aHrcQVC2hL0TXSUgiHhJgx01EKj
wiHlgF0WkZbgVjZCRjpm9Gqr+OGt31f1VMeOwmRpCh9vh3TsZX6JQD4y70lVIIyy
ypqFc5uQIuTehsK2/kkxXDH/2k/UWEOAdhzBibr/+Vx7d5/j8tf41K/y4ZCZz3Zc
zuY3YP6xtjBEIfYL0x6DWANTqFZsc0YAsppVY253r2hQ6JkjlBmG6n3BzhdvZTXj
pLZZuKIjX8jNVlBIGwXQYmH33DiltmWND+bswqSIbbA/Os0kaQu39fZDbWHeku2s
2He5xGaw1DHNkKm+URYyar+Lh3PqjcHYmJoh2JW5UVz0NCGNTc1U4kbL4QPQ2SaM
EW3cnWoh/x8Ap7s4FkHeMWYOlAd3FNjOko1s+2L4Q5zdOLIlK4dHnex6JYd3zC29
58Et/esLKdqMEvS72O1iUtJhX8Y0dxQWazslXuYIdDVje1UbN6X89sS+87jcVXCa
Yxe88K6n2Y/DxpiDJQrTOMiOA59o0FZxEL/bgjGmPXGniUSy2bIxeiGA3zKBNFB/
M6tQs3wZJIfo4Qi2SVwdORO2VA5nSsWUNwl7oUm4brosDaXebhvBc5oSm4cRh1Es
h8YH0d9dIc5zQaw9yqMEhsiA+H1noXi/Px4WuSm49+UZTc+QPMkNGpkBiqUDvagV
FmqE2audhnyxlv6j6mwPwoDIfTp+4gZ3P6MaBvg/n3i/kBJECZgPxaTRgwVj06Ky
LyRxMvlDFu8xbNr0vtXjOsjhVVXTrs4nT6Xkbpc7H3FiKFZEvZlP6xbjnT3aiE0E
lsdK0vQBXd0f2O22j39l015WtV7PfII3WQ3Ypf71sWpLD/gCaBoRlfcGw/y3dGcO
hgbSfMVFl7jnzVnYWZftQG4F1SlofCPM5PoHwsh+k+wFIpuhrV438waWigkK6A82
r3hIflHqpk1Cs9IrXTuNhvy1KK/pcQkdKingb2gNgUS8LFZKlc80B6LO4FllLCvK
IbL1jvS81UVG5q19lLJgH9Da28PllYIdhr9Tg6FomYtK0+vFtYI/aQz/LrC9lOua
S2i83SorfQAX/FeQHO790+ODAp68CkrThcxyMu5RYO9Ci6uxnSCBPZPMrzc0xcCU
MLA6dzUKt+pJfiwT2xTVQW4hP8NFrr3d5ZQCb3NaFJTI5Y70adX6JRxhhAtEzI8X
zpIx/QBv/zFvrkBtznaHv+0u5HQvcExaf6AxPOupUVgj8YlMKRaOl+KtfCIVgzCB
HDrlLPrZaQEEKaeDJ+vDdNJwkg2CwdexhS3Nya9QpWFPCxNx3ysg9nW4bWLw+ma2
AvmqalgxZwyD+ZX7lPPdcOnImjUT2JekW1baOMAfdxUd/XqE/8x0LQR+UTwI0AFH
ZLc9wqfL814UIMx8oXFxREltmvyACOjMlG7qHEKi9w5k/PDmwH+CVuOME1TtaZUo
1zPmWHeQ5ImviVB9qrjZHc08uAd4+wh/f2CfLOghnLeEqrlLFcNQhwHnd8IiyBB4
f1QE2nvTQWrCYGquEIxNpd9itv5RQcvhG85Hh7O4O/jAvLUE4ye4jNv+MOtuGZI/
/zomP0A6+2zGOv2D5q42pbHySnk2XnLAyagTwb1/2Q1ydlAmm3Bn1NNcWupe/hCE
zKQTpdURq2vwbT6WxfBVub1Mhq1BwGpGRmNhxHORMIC1x+9I3kTpHCfRIBW5rnWJ
XDjy6oEMRiq96ZbCVzwfMbFfcDGrnAeHhdUJKukVzTKhsw1j7MfiVtaJsFyp6F4d
oVxkffXlyyMihuPEy3l9LZHdl67COFDRl0w76m2w1PUHNWZ1AAJivp13Wy1XBNZA
m/zQe0sIsTQjFJ1mzT8GoKBKHZ23KlSzfv+m3ii9+SI+PaZeuTsep+Y13SUj8Dz4
4HXGjT8HlNxrV6a1fXkqjneWRffq2bA9B02AcPV4kw+bSzEZBRbNmpTgIXIrIQ3c
dr71CGalGSV20CYSOlnON1oQN+xeHgCHPhwi2v/iF0Z20tq/qHOZtQaqput83pHZ
NwtK9HLJm9TOyM0aLbFqpbg0TK1imt8rthHtswYQR+QAYxUel3ZFUNjwWsOTMQk3
wCAhlHYFIxypBppVdQ8h3QKW6eljmBYuCbsTcEAtFSsedSUsrWfEsxnUTlvo+MEd
NUyUUSsy3hulkBIc3nPfcVFnlzXIU/CVrA1FV/cNB4c43cuVwzEIuKRyDLfvPNEz
1EDpppWTYglYVhF/JIDPJgpCwiH7WK1i90Dnk6H+9iYLHJEwLEGFuWxZJaH8IWND
klLu3/3/PQYmatHZ/m4FLpNezvur0EcpIb2jv3dP/ckQ0LNN0i+h+Gdsf8DlBcqO
sDJl4408g5tmndoAdyHyINVnbwiHMAmcIZGtCSy9WaIh6nxtR3DMvB1HlPilWoxz
+f7zibesxeO7ve3pxPc03sxTRbGfsmU6QxxDR1dO9Gn6FFn6s+yrC2Y91Q+o6wKq
emPHI+wIXcoxy15gvH3EtRl4XLBB+uT+ZkImF2sCxwOj5DTcdLd5Ag2GUV5qIMAv
cY6+Y/pUL/Dv6Zs/b5aTIzuwpv9tGbiYC3aKbBYGu+NF+SgTOpuppa4IIPSh6ooE
i3scITDkSKjm6nNN5fKjzMeqCYonnn4Mekm58vEClR+gbQf47S1zQAbW/3T+deo7
iJGbZ8+eMk4aftrbEG4SCk+ASxEGjQKElDthyvCaeXM4mf7bgdexFZ4ESQ0oM/hQ
3Q57Xd2o9V5KSrh4DMIxUIQcv+6Y//ePmYkn/2KNIaN501hPDjQ3+Yxqr0IXrlpY
HZS/6lR0chKABOr6qjBMY0MPf4rsgql2ZTNZ2RdBu2WL+mRev6rOXEmtPn+OqtfU
b2ym3LC+YpgdORTtYKJ4lSocK5d510bqsleuQrZ876QRfOUj0WM8rd71OcgKcsKw
hPrusFCa7/CaohWdjtZ7anCRufjil7LjKYL/YJ8za9vLWL0qXUx3z64ux7YQcrBw
ayBqSWzgR/fm8S/V/RmVBMepGLEr/5JwCfJeM9yFZ1CaVjjRK3RQZFa2XNqC++30
MyRBPJHiKUm6nHoyFt+lT7Mwj9UlQt84BKRCUIZhET3cNBAW10eE++D/SrNNBzxv
cU/3GYyvWaVf9WggZ9NWEnfhb1LHHkRHxLRuwu5It5Tdmk+79u7h86weWqzqdZHU
CWOwnwPLMpO6A8tPI3CE/ElVjzqcLjSoT86jLFN0udGZOdCAh9nX6SxQ4xtw+fnj
6jRy81jW4sCi6QO9D5agGN08IzWaFETDiCNkAuv2a08iZcc18LD8dMsP5K2iqd3V
aERNtsfljs8VIfOk1VUjzbc4QnhVnW5Sgv7bGLVNDhinO4UAEBDClSpTBMSu5Tfw
yfRuHBIKTaUhE2KUSaGqBE1kB3Jp7U1bbFFa8kOhUAInzfvE2N8W+S/3x4tSlRfy
ad64ave1/Lq4KKXx8Qz4zPOMoKSDbMgahbSqz1BVMztdd2mw8PSYokz1QnNlWiNg
QNXD1MzM9CBSOlamdCKsp5ThH8GAXKgcumSyZvf5UITSnDxGfkhCnqc3P4B9+Jhp
N/Q7i8jXzso/8p642WO/DiMJs5uelOQm4c6wmqWBj124cX1wNQQbzaH3ujmtau8E
2p/TL3gZda3et3Um6t8EpkwhIoQ9e5c0josevpxODFLtL6ICf2Ex9N43mkHhaBLO
U0bw16XFA7dbSOnurWFDLeO1jfhHlLbs6pXV4NoYSo5cT+gqyqg5zGdJKRUygTKh
rJP00M6TbzAMASDWDHd5bcsJsYjd3oKpme9fP03dkWdQ3DO7NNowWkZ94uN6B7EK
G10CNxVFeu/p7WZ7+s+CRIaIfvcK2doFaytHxc5OSApb86Naz0+Z8lyITqmbzwP3
Ey7lA6Ufa5qsPMLtlCjH1t4/OT5gVEjGNmIjODkWSMXDJfsjxDUzw678uoTVZ4OW
QFnNCuIg572258aVcE+RQ7npJxVQpt9iKEmAZPPrCPIBMbfaHCc80kyeIqX7GFZU
/ud581+qcuec8NGTISIzaFva8vXGSMgHfQ6T0G+iuQx6YNMcm9TbcQeUaGQUS1Hr
mjD8r6k0kKumLq7qdXGqmWcltJ2PE7V5YwwylRiNsJ/S6xE/QISrjeXHIsmI9Zys
WPoOJCQmEQLc/VSaC5knqFOf/kD6RLato+caMH7Xhz3Qozqs7WY6jIpfbRbxPExr
DUfj7RCeQpMh1vtfHXUq33ZfqzPubPPqulvc9U51M3xeGjbyfeabL7kpnLgylJI1
cImVb0JyAPvZ59/fz8mbsUvXsbBTVMqEb3Nwc+HyyYU1Qz+BhOgfdF8yHbEx4DrN
4nVhiG+g0jnzqEPXlnqDaOtEmNYMuGLPBc/F9IHq/hwvrVVDaNmWjY5xesdlXvbC
7TOcdZLwk8/QWFh2h+Q/taLKfdBEvMaBQGUmU3RzLYDvsK8BY6bc4sLnjUtbj9ZF
p8QI5ZYwWxonSuV6aINmO/uRSVNL6hfZp/O9ou+uobzK9vIAALMMdOA4f3hniLlj
PdjUq9AMUwluzW3nlEjfXJNRd8oP3ICSOtYT49Aak7VOJIk6DSYWK6x00aCyTCJt
ni3fwZ7mhuASHv59R17JyBMnqYl75PL7kU9Fbnqr69jqQ2oFfrrL6evpx0eqO768
XgUasUX37oEptPeC8YiYTIpjNkRGJ9nau3k7NMlS/M5BZ+0OnRjV4FMcDney97YG
kEXb7oNdAoAEHBh6GkwcnhkArTBY9ZtfA24C9jCTec0t6J4WA7z1WS02nSmEbWCS
7mZNI+/pDX8UH2Vw37bXvnP+LVjoKvhgaPUeiU85Eu+9NBsDb6YTofqtynVeRlBQ
RpHlz/F5G9K+np83hg02YQI3ZHWNlTDh6ZAehMo7l0nXl7EhBzri1k9SiyBdNsg9
4aqmtTYbOskDE/Fqfx0njfZ7T4GC+B7GvWNo2a8wC/T1jIlowOJ3wREr2S4mLNcJ
JTP7dRjYkTeFRPpQpWl2whGa96UtE549xjBf6mUz6859ShhkEpPyyfX8oyN8bqDW
xjgExYk+uLeqT2SHuArx1LPzAvS0F5SOU7rPGFG8m+pGKBJwGqVJPtycMpmEiMuN
NY4szzeYenD9imyH1V+BcBZ+VC7XbpULNxEJZpVWP3dXMCy8x0xKpS92VlB8Eg5i
PWgxJXYRYx4us4EZpMSnylj3JRBxNOe514eUMFHPENREj+rwjLuoFf0qxvs3QUQ9
k88JAN/e0J50CP9iHSbeOR84WulDrOkM6LWsVxtIkP47rkD6auSLgiTqDHY8ituh
z3w9iQeyMGIaaT7e8FDoU2UI/S8MYu76oFy1toc4hDi/q9vPhoEQUW48qvVcUtPt
7/FFE0PuXW7dkPbEJxspqQAqykdkviNT2tvjqyO+L2U2NSIWN6d0px1jfvBEyV1n
j9TNAKglLpUVPpbew907G+EeZ8XmnUFvB1ouCwVUDow/r09F6LxzBZNfF5NLxEaE
QIq93T/4z4peXYYXDtDx/96jAT25xL64HUpQHBHv2GfkV5rR7aYS2stPQ2cMXwVu
DXhdnSAPHW8yHnp5EUDqzXyYz1pXMUSHdkoVO+e/U6lK062OEJX7pRj4A/ML28UN
lmylp7bPK0l22fG2THjCdel7/rTeLPM+6vViLgG0Tr91aoN6lpxopmvn+0lCeyej
JZgUBHypQh7Qb0Kp5T2ul7qw9U+gr74iDi2lsxJAUB7780fFCbtcU7PsXaaLm7wq
vi5TlmYzrqk3gfIACP1jpA6rn+lhEoefDTShrFttyMAPyuYXY+r1LiUy2iefEpnv
oTVbENU88GoSXWsTwek91tBC5eJTA/V8Ehl2lb1DxYDSHaFth0WXUFte54HhuZiP
QV9x7MS8RcmlUcdlmtnXobIH3VfdJ9wWBCPpd3f7x4adl2wmhM7VSblCKfDEgtR9
UZI+CJjJj1VaUNnuLcftL9o2LlCigyeRPLy+ukq4kXk8KBZdeMp704s6/B6QPYE0
OEE283BA9q7nnguChyq0rRhfS6/rDeY+0rMmEZgUdhr9V+teNyrjIy4+1xr2dkW/
qTWLZCbN9SBRaGSGdLZZyqGlaELypdp3vE02LIEQg7YdTBgwNatNROTlrW81yggJ
dj7iAkX1q/6R5AaZNDP7xdNuiIHlXl7s96e+nKV7Jg/boI1Scs+3X9n9qrbupDgB
SDmp4GHRzQZmExpFKVlLZ+xhR17+lf414fXyJrnwinq/TtpxiCrKGGS7tHabKP7z
EQxqlUn2b+swJu+PO6cQ/lvTBNGRsX+DSZozzGbvZaSo2ZKTbtXpH7W1OUvidhDv
CjeT85PQokUiNtKAGsLqn+/BpwyykDz8ytrtOt46MTP9eB7Krieqs2b+cWBh8Wth
2yN7CMxhbvx2AZ97f8Pb+RniYvdyWRpNDjs0eykY/Z7c4P/qUrSXs6Ju1tl4FPq2
2BuJg9ySaXLOkBDncS/BI7bH8PdFB0438m+FW09vvpRt7MrKBkdznWoXzZomDJDq
BRuYjCd+Y7kbUpTu+mSvleMtyuYyEjhD76UiB6EzXKCPyKAgQUdkU8+JKZjUNEDH
CqOCY3HOXad4Q/H+EfYWZNl+svvN9zEd5CdC8XbuL291yWh+YnxCV7dtlbYOX5QL
Ipjp0jCXOYGBbDnwasoaGP1SpIJRExJQ00yyOorvc+WjvcnKbtT5nGNkYc0RE3La
WdO33+vpjc1sHOl/wBqF8uT4cd53Ylo2PaZ4RUryWBXIy/M6CmTsGzlipxf5DECA
HIZaZ5WGwNNcngQ+AtkDvUowlfFZ1fbeab0IQIdfFd/rppmf33+sFLiZfK91i0Bo
nW8M3Cttcx6B6xnQ4bkzoLoSsolQ1oMuEQyrm6v5TAJAhzqfST5MT1pqOyww71bu
tg5yELh5CI0N+4Dlic2VQsQ++Cr/phOC+MUOqJR2UD1UpwfJISDuGmuQIJzCcpRo
sIuxg5euNyhh9LiSX0AWEDxp6Zoz5xHh8eEp6hzRvRlrd17MSeI4Iik+kh8n7+yf
Nup4Y43Zs88kYVC0N885eCNr3S4AsFfINdcJTgcKZqJJe8qUlqmiF+GPA/TJQlme
pZsyWcNY4mKC8p4mmhIQCu6z2ILGnIYadJWdNumzh0YV5SVDHwZgBvlhfLdqfyys
6XwM+y6o1ArH5TjZ0ZIFXQxonUNC6iXPGdKYGl9yA7oN1Fe+37NA1bwZxvtm7ACm
l/jvQmAsJfX2axVhZNYAFqVyZ1RnijFMgs7ZpUTg7yAkJeufBDeVhwo4y+w8KvjR
NRLeiIVZs1dv2svdqYIRv5kxk56KwI3E3ppXemt5e8l6dToblahiCUT2hZcsoDvH
6qjsGnxR1l72DSuLajI7AFvvt8SzOCLBXxW8zPrjMaBZli0KDXh/u98V93/9QhcA
OpsnxJs7hHPzxa8GGJjnBDkCAD6SYJ4aR8JUU0tyk8qWVQSJyGpiLVKIIz+JRT9f
M8vip+Ej9NssKW33haE+u1z8YZQ5klBuU+EcJgu4J9zOEOxncNEz2lLQHb8j9gij
zs2e8MYdTRQpGAEMwiSLZ+P/mwwgWCu56TN7BZwZkYdSaly6ynZ1pXg4m2sI+q5i
9Y8VfUGTg08Xe+XAm/pCjXRCqHRDYYs05a3HAppFGAjeUURO+iDoChIb1TpwNQqK
DunSSNz+hXy4Bu5ibct1+ArkCztBez+0OfXXFpXqM+M7X/7gpSXdS++1SaM9UiOz
v6LgUiwqvUQmWbaSc9OTOrwfQ6+2cdWH/npcEDAO+h1LsWQ3MaxL0w4D9ayWQFeT
0B2TgvLJNdP5/CrUNq4LsaHhEeOHLFSsRfhaiqne0i2NftpHO8BpmsU8VcpBrlfH
zAZRorICgNelmx0TzcdlinD4dNvHqHYeb+6d/KH9JFs8NzuGDMyELLeVbgpx1C63
QpU0xARXitptBQRSEWR7PV7X1qq1nkrPU+24k4mArccQzznYYnpm6yw6iU6gYSJ7
4330Xop9fjecs60H8naaMFq6DRxF+3ADn16to2CpXnVOcLox6kDLqsl4nQFCPlTk
fQNP/Uf4hsirDrc03r5kZxe5X5UY7472ALClQGTWspzRV05DQViQot/Zh7h15vey
oJLARHR0ynw45Jk+SL/mcmP/SWWtsbu8M13SkS8lCEXTFogF1pai/0Ki1AOp4+ak
zsVpQV1fyeRXj21OqHfJQUf8Um01gnz/46NNdcEiELvMsWhHn4l0xPoVw2uguf3x
NQbuYJ9UvTvzvxgnX5BRk21lpWVMVtTgkeCIaxE5dfzp7bN3HS7b6+2MioKCPszg
rqrgLlWm4iAHvqWME8X8VoE1ePsFacTmOawQKEt7B+hUd7q0Ilw9Deg0LdhhVyA2
nVkHxIe/HignKoiRZpcRTv0F3+gii00vjcGGZ9iV89bZdjDlDEkFLMX7IYDY+2xq
s+UFohIMCWNVjkPYvpmPuQ/J4Skw9Jm2w7e0sQI3twrDAWTMK3hZpcB6dSrjJZM8
C2FCrAbTNJBEuZswcScwvO2kNDpdPZnqH7JaUrwazF4CbPnkFt6CA3mVy01BLR9E
d+Cs1Mc8Uw9ODLrervk8wtBQzdKuMVlc5Hz80ZidtOTzsh/uUJKex1scR2IH356T
mJEaXHHwm7WKjlhe7sYfC/Z3XRNdUuD3XT8l6dM5JgZNMp9cB1lS40qArFAEhE8Z
s91w4vmGZ2YFntvtkSQXkVDNy51eP3J65gDx0HS/KD5Rcm8LtbYJyeEWeCduLhgS
w3L/5cNaLYYagjzkwsnYgd35t3zWQSFARAZxcHviK6rXncNAO8xnpewCAC2+igx2
XdxEzoYzEYuw2x9DtAV5D5ZvgHdr7UcDfd2sYRShMixEdpyYkhDKWF6XfgeM7yqO
MA0pzKthvCH3Brg4fQEaoFhF5I62dzas3sIkwolwZRFzOWwRlhX3K2NrFMv5eu0L
T5zyX7fV1kkeUyCL/5xWGfKYNqTRR0UnbciFlqRkBYgFyBxxFQbvlVbqyF/tHvCt
kfdxmCNetWrQSqvD81quEQ2NTOMbF/BvHcoHMeJfYQ0t2SmVPkCwyN61YiJywDfF
3oP98BHXh288Er8GduDo/DUrHubAGpLY19DdfE3gSoyUhe1fNP6xV+7wz/gQ9AFb
HGlxYr8flBtubt+mZEzudW9q3Zo3WYMVal54T8WAPxxawsMqE1zIMkHPWTk7a98d
dJYxeWHS4kAQlLRHuNPC49tev3jyruAzTn1ULoAjrW2U5AHir7iq4o4FBaldUEYA
pshZNfxECSgES0LwPgXUsuCyaIQcdp7Zt6gjHHIxpOU5HtGbOABUTareRy4e5V4Q
1VpvKdXZ9qosfQW4SHR7PXke1FtzfW0ELn5Zro4FtPlu0k7fPCe8rFsLm55Bvpza
AE07o/MxoWms1rwix8dFCdpgmVQ9NAgD6jiEM2cBwaK1xVVDCREk5uttNp5YAmmJ
SjrsTaLzWk2u9V8zwEKDZbeDJUfHksbtSsZHyoUUZTJOMg86O9Hx80nGnhO5bBrZ
+NPCnY/RXhDz8wl3Y9RwFna7GpcEHUi/VqdxwDjbB0AhB+JfTPb6tIU8ifKKJzTb
ebogNibQO0i5jJMAe9l3F5d/uvMKuy2NHlUkjs8RwBIolAJgwl7QRKeQgzovvD1b
Yw9RuJXwRlTvu0QNrjG0PcEUK/AYE319SLjj+S598su4quYJPZYFH9PoSYoYtHfw
k01ldKK9F97jWk9zBKQtyGwB5pXPia/GOcfZ0CarEe+NmsjMaxKR53uDhq4UUlfW
8jvFkyHkzDcXRWWJU8QyrdoN+U8mT19+mIN2DTOE0aF+JcSLNaLRRM7KCEevFya3
6+EnMvoortERYdaL2JtWk0i8NkHa4F3ljb3x0rwPOywWzGyPATd2qyphENeRsDjz
pPg/4/buCfsoB7yFr9GN9HOrvGdbcSEaofcqQXZGPpUub/K/99T0++Ta5zXMr5AA
5ghmYZTaMpiILGvfW1XY0CRBwE8fY+4ecgNw+IG92c1AfkxrLYcR0EemkDjwBr/+
oDCFrzYvBwn5NL4UZsTgqIvTXPZqz40z82NFv6ryi0mqFvs4gqEWe1jUdzSEHD6h
RrTddAkxshN0jmjvzUzrWTytiokVOzucEYqnTcM3YoZ/q+rVcUUjCqB1jNX+evnL
2fw6euIJC9vkltN0/rdW+c2PzfaQ+buN9ClUJwoU6h89/MvkCedO+QoIixssJF6F
3dVT4qEZcZVRXrK4oBuX54XidDIxjTtLQ6bDbKTe896g5bT3eUvnFjqQ7mmYsr7X
F4OMth1x4GvrKK14VNXqzy8Eq5bvbk6Bzn4sql+5StoY56b3YZQ9ql0hMBLSQqjL
PQ5AwUL/HvOPyjx8lVurXRZsj+ZinryofXN1eXJERRvoS9IQCnX4yzjGBjXPs/iD
EyMLMxWAzfmaLuse56OmC1fid3ehfe3GRYS4aqGtsT2Q1BcPHtt7pP7xLLf0NQ8L
xOqf++W4RI+WnWtH41jaPlOJjTrIvp5PhROzwLtMLcH+1YKG9+MsFVwgjw9HCkQw
qou4q0TtbAPT8wCaQCw4GzYAuSFa1hTNao0YSDlhKuzw6JXS30U7ZsP6+5sGxAo2
27lWJHnDWGuVa1DLiH8SMylGtVGAjGPt8p0URf5DV6/EIXqEvPUPM7puZ9rgrT1q
MWrXHkQn/VH+r7BbN57pxHxQ6HGZ9nDWFUfrN4YSMwC0lqg4zhNUepLo2MuiJfGu
nMesD2tr1OKtXpq9h7ooMtCWqROBaREZ4arKCJYtSdpq/dMOjYg8kDQeXhyi1QIL
3kSPBuvn3qRT0/r8+NU2BjffnI0JLJdysxX2O1kLYh9r2Xv7m0mCtrfMcV44k4t5
28l/fmH2BUllRrHFrgykbPkYfC1rn3zASq1pGQGC/K/4t5eXdFTFHLm2Y8pS5K/l
G+kK6sSuNpVXqcqUheOzbXKHoGE43X5iMYu1yh1aOpDcCc/2F+90bLy3OsMfI80E
Rc3aRT+71a2EkZVBKaHnWqe/2usko22lJyPpza8MnN+kqnvkP/O6qrDCl3MA5UJi
XshJZL3WxTUygNovdLqtu10v4iW/aBDn0wOx+nnThtGenlipOeYyzvYkV16HQQds
QAp7nVGHHRhVrPMTgohAgQyhzrSLULCUayfvSCM1lDfO8nbmIvKIWK7R3fktqBnt
oodHQQHgs1QqGQO/1Il5bpIMqCErWX0JdLX0457qU91UsVpFwh2xEbUKtVFSLYfo
Rdb7CtTnX+KD4hBAen2XNJYrImxmgKK/J9RR2qWyUQzPtS+wCZ69arKocaPpXexL
CWLDxUCJC1SbYXPRIAPu3l2TrLsnP3ei9IhB9mq+Jgw6XKqeVm5ByXOePoOo5nEc
+01MLh+j05TsbU3Z4fVOlBzhYo0uIraZKQz6BFu6NuOwoRXPJLbUmJJpy8Gcux/C
NBtq+z2wRzjtVLkIoDYziCqrnXKCDKwaN8SjmRfG5y1wlOeyDCn8odAWXPcDto23
WypAX+lMow9yMzLqzfBTrqu59CI32AQbgXx7bCqmxA1o9deGTVCVpqYwvlUf9Bom
XLzMF/Mhbzenol+2VtD0lftGZD5fiaJYhTPzzpxXE6ZO/dLpmClQlEToGSo0s+pJ
gqRXdppseiMB4rdm8kLrZ9nE1y0GAglVlXCg8rQ8tMUYa/VjZoUlctlL3sbJEiTF
rUeXKaexEJYQaXxSx4B42vMyg+1rD4cN2NAWvclQXFaSAgFLhrzfSU5gcEXR1L4P
0nApEtDhDG9LntPP8GUyFDlQqxJDfzw4FTV63Pcvi9ZC8vT+rXOBgLn5WunEhz3R
CVlMk93xvRVwZoKAiOpSqHUN0R41Vo61o0cbMWzHitmjOrTfN/Brl7qbCX5+DFUa
GRwbY79SagnbXwASWGgayyWZVkz/mvdfMogIu2TZWia7R7vFzdiilrSAZq6k/FCZ
+emymeZQybdy+tfthAi/6PpbfvkR2/+sDV/PetKT6j8zG7/tk+u3cJrrG1Nl2chJ
HJmqUFNIFkNexwNClek26mbCbGJosLK6N/ZT1m0LKRTicTCxqEr7b2VWkHbSOSD0
McrPW1b+SRsiaOTuaa8K6CKqLAp4JYBn0QAO7YvrfJeXfIpP0MZ4Vc5mL4ehnb+9
NNf7s9ykGpLDUZZgmgCWt8nwTWW7hALNj4/XF7nEWSXJ5Z90gBSINegkZhlO2vhG
pOLir0Bm5EMRL17YxI+emCA/6zT/6avlAU+kcJVq2y1aDY9DU0EQUR7atYqWqmrx
u5J8e//Fx1+HuuIAwncXKayml4cgwEVsjf4TC/MgtmPQoBNckwXrneHt3K5L71mS
bmewy6TjR4WZhBxHzWlfBHIari05qb2VJLch3mO8xTt2EGcSDxE+VGd6wyYJfUcG
Uk8Tpf67q9IfaObskA9FhpRfpYz6SbX8P+cn9c58CVcckkRBX5Eg6tB7JXso1Xez
VTCrrXVy1ix3pzsCm7ff/fAAlNTGg3GTPMSfRtaPsayLDg3qHoCnP6LT7AJ7s67M
CCGK+dOdy2Etke+FMYiRQwolojCzWWWIYUNG/4HgdK/bvSd916uK85cL6Yb6gt0c
eg19IxGjzrYp3MC6IR6p78P+lGnJ5nBOayGwRvd/t9+Y6TGebZFSMysNiDTrbhoW
2CPEhoUSR5ilW0DLNz88qeoYP8QKTcrqCc+SrpWcpf8HP0DXfIEkFjYbD7XqzVUY
ka3F98v3yZtRZrp8iaS7xJPav5vwoO4f8rn7IdTtmW9ZIPmn7owqkhQsWKwlK8ZE
+Qj0UK3HbifY01EAzzSeQB7vKO0yrDvLf+tBKOTrjYOSSaoceD6HDm9rZGPw8epV
suU1fkLfpgDb1PFoUbouuWUfJK7HaM1g0oIgMkAAyrLCjLXtUSdtLRTAYIhvkz6O
79gy6e1NsfI2Yi/LMoEF83PiNkGttPaSQgF5mVMcOwWIm845wgPcG/HApW565OQr
y25yRUayzn4cFf8jZSI117mhI6NsQXsi+GkDCajE9T64jB1i/WR678RTkB5fiuBX
4KKW0q2Lsp1SFsmomNTbeTdPJwkplSS/jA2msTi7rlCN7lRkDBNubx9PupVfG3+M
nCJVPu+s+LCyNi+kJumtPOr/TCHdmt0il7BHwmBiBNckU7tSzYhwpuqKV5oxWoaO
2jfzv+nR7HaoblwxfTlWg0fNgWnkhsHVuvWrRNgVZynXv/i5yGOAGD8JEd3MnTa+
Jt4QjUBZdK5qnUgVSQ47Ncr9jgFbRDwMOOhhKzR5w3TuKj1ndoJwxXHUHExgrR8/
gNLVyTwv66m3EmNSD6+k3SppQupHg59iMgewQnDPZkPNQrYvelLKXSkyXN6OwLb/
gztDWZ6DkX214hBw7Xrd1SAolbdCy5kn+i6s9ndBk3pUFrcaOff1N63orPuAYi23
eGeoChroHrZeIBe84QzDXpu8+HAuaEy3K7i/gBp2ZASrBWKp1k+w+n78oIXUyRTO
X761DLZLiip7ZTEDLK8apa0CikI2hASZIVaOSA3PBUCCV+ZqgxwTN+S2R4AbGruF
9qB01LCHvcZbf6lcYpAVk4vNhBxf0l+QVL0DiyLyHX2cAL2AKUbE7BVH9sHdK9iu
aDzQSugPueCsThZKUG50t2S8VG92ntODvmXL9pIRalHhH+sfsw9o/k3MJO4tGtjE
nl0mZFfvRqUE0x/Cf/rpUNmGqYZv0/1AAjXQEaP5k5LJMbYu++D6HGW4Sv/gPz0R
mGkfgCK0qCiSwwUbyFQkAA/o4rlNa+avGvTXx4xYfsUJgZRvljxFI1D5zpmmHdgD
aF/Zq4xSQUFRMudaNV5m/+H9MlmqSs7ILJvJ0wtJwLOEEsLlhxNTnCzUWZTIOXGZ
9jGK+5mx1c5a/YFrwK9FCAp7S9tBcp6uYwcK9YF8OkYk16A+KPPW8kXAuFfJnv9N
M0Ux/MY9F/fUiyuqXC2uccxJIoLsbpIF5YDj2LQz03WZ+ogenn7PjrY2WMCctIFt
yNjmYDTKAfyfPm4wcDJMaNudQn9V9ufF5WW/v6XKFNRydoGNpWEt+J2rMIl9Ed11
CFSM47aXH/dNA+T8DNIZOmSx0ZBK+rhFbGbd7xxo3NEhhFt8yu6wC+A4TTv6QvPc
NbdIYZ42tfupqXy4aN/UwNT9kP4IhoSXZ7ac1DhaCtokhayYEfgG4N1WverNI+am
FnMPsXE/9sxXvhgq+CR6hqGhDwSFoFyZ3DpFvHFG/w9fZ72lxbezmLYwgDN7zvHL
DlQYw9cGDLqszpbGRsKSCo/M5G4TyIThz384zsGkpICRVV/U64ckEhtQe9zQs5Z0
NYZ4nupu/1H8dHONGg1kHBBEqFItXTvPqAgKVSfrisjtTQ7ZKG2ITL6UMH8ZhezM
KU9HFe8x1Q2+bSZTCfLl7t8xGb/Flp4SSJ7OgbR1+xetCR3zH0BvuxXhE0EhtjYc
5oMqMHDOkiNoF1nYq1tsuXm8o02eZ44H4R8e/wbT/G3UhTwgsb/KvvgmpNhWVUi5
8JCrlMs43K+GICunn6Px8O6HOGscCdMOMXyNV/KiOjeIqtTIHRKkgB9GAK1q4dWZ
UvtVIik8zyJ6MlmZQc1+StWlO7DnPOGzS0FNEV/OxpPMzsyrOYvkFkmQl4INXJfU
Uoz7/uy0j6lBd/SiqJe3FKV3C4JYcasnfnTUgfxfEbWlf1d0YDnirWWIWtMJe9Eh
6XyRaAVFx3FcTYsyGMQzwHG+kW+ADDdV5zkQwbw/TGWX20X3tmkO9h+zzfuvDELx
DYf4NL60pnqnC3Iu4MRZuNdUTq1eyryOI88ICU2wr2f8/aqcsne6aUi4y1v5ZHK1
2pSaRxosNLIxBA5tX0YgVB3K92ire0kHWHBwcpaIGBnf6rQFGOkt/KKg/Zd7qcAe
stm4X3Fa795CDMssSsrysq99uOir8NOlCEPxiQ7BqbsBfwwQJXB9+5ErL0239deo
/QWJPPlksTJ659FQEP+OAcZpWKCzgjb/Zrh/q9r9YX1rnpNtuxu3c/uBLH5Rdbe8
JzyUY4DFI0WXnCXlyhbQ4uombaXOw1Mv8m2/7Wz4FxJA+vakMPHcbV9SpcSgBMtr
KHnJlMZIY9khPRHOOV2QhzjCBJQkhfy1nfvtABsrKSaNrqGOa4uVC7D8gOKJAX+S
gpsxPyrfNWck/dXBi4xlJ0i1t0tIrrvvKlvsfd0N/7rtzk3sLHi8fOE8SpMnopeC
6LmJ9N0NmS4RBf7FfI5Vug8ivVyjAMSnUN8qUcPeMEuyK55ZKSjHpZXColN1CV6R
pWyaIp3LMQdswEpF73DL+j9bP9sumgN1fimuRcta8YFVcqtPg0qegRu2pTM75vMx
W2GLUsy53VtnO/YkslrQyO/+xzFTo3YoMq4/kQZD87u6R0I0APjRvxp8QyRDXHfm
JllgAguVpNcFXusyg8Ygu04ZF4YBYBxHJBb18roMo7u+qDpgzmD8uZhF8lC4/Her
ncMYTUK0WlkDtf84ErEWNc4ZJa7U0O586NHH6P9XhA25YkIMTqHbPshuoIeGfXOS
9GRYXPfvxfMOTT001yE6ifnLpMsrIn5KRo7cFONAF6X8qWaE3m9B5Ilg0H2nREGn
XtxyqL3qrsikuyWH0ezuTDFCxe04NpI3vHRHQwDeRn+0RXmMuH7b4PPjobP2F6Ps
4Lu+BUOlt0cDrMnTe1FNedqcgWbiMW2CUGU38YAKV0Mtcf3C1r6Nrom21kXi9sqK
Flszib4gpfflJVZrGAMhTANEzmFgeN6nIVzmMPcxS/WGTfQx2RNzkLs74/yWHbJN
Yoi0G+pXJ1smCam0tKTOxtwasLGUriae3NuQcQHCCLaJ+JpUNBh+2c/ddiv3FDib
kkq0yJibzhPNVY0y+8JPkjHuI8ajxMNZbbktXqgKNzNzPs6FKOJY4b9+OEBSh9WW
LRQxGZHtet1TeRR/Y5/N8jxSG+ymCl4d2OalyZcjzTgdCtRhyUiHQhpcRQGO4cOK
gMk6QLRMc3Ulqzx6T86TBkwSnvl3AhMBpgQVtI0PSrYJA0lDxR3kyxU6UkwDEJdD
iUZbbXrESfaRTSrii0XmcE+fAQMughqkDsPnOZgW+JhNhqQ7ttI39GqcO5kdA0Du
nQylFeKviZg45TwUJtaVywjmF7lDumpUoPNkWdgQx9bmenzIUqkEx41ISR/c7m0Z
xuIit9ZKh/00hCinKR3sO1n9apsSIcHnh0P3oy0fp/CQy25Z53TJcdfBVPS5wufn
g7ZnoqL1HQelhil5i6DpL3kpNfvLVwDgnxA2DnyJl/43L0bc/yMllHWw6JodniSL
QFtItWylS2bsYShLhgjoUj8W+xIMFRRsOEu3Kfu9rp9ajDdNxVxW51iscgC+fDx2
BrXuZY14KNSPAZYKzj6IhPZUGbHh42ikv+YkWMqv1wYcBORaHPXVoQdHsaypSGPU
7+C/HJkeCTLH07gytR0kjQ6G1UT9Ph44vRig3+Hg/lMIwa2QENwcxpuTajx6ClEl
VixsI7xcfimfaScEiow7tSoMh6OREcZ63yREGdmC4mzj9Cx/VOvuMvaBg76SXO/s
RrGCOv020OeFlpmpBN3+87AwqzyWZIsjiKXdF50lpwc99S+xb1z0Kh6D9gXkPDyK
82Bu/vxXyh23svi7PMmFepMMSdYYZLMlDv7TSck/6IFGyt72VkaGQLxUYzPq8grj
Xl+QpHSiav8t3OxXhlBzIXYt6s2n7ocATyr07xDv0QOCynO4lBXNCMu2SNCwv0LD
+cSjVEtKDvYb6WEh9PrdeA6S6swSevo++0hAw3lQPso3KFHfP78EolHQRX+u44y/
sf7ptX7EKfrPUwES/VxlqW+ZLuqVXPJUFIHiUdvJ1KIHCCF6XfzAxhZQERlwLOIM
UfYa7MsBl9L56d3U4Y26DxoyGpTq8gvk7T2gn0yF1yHWXEradmFg6oDP45Y250Ee
3nCFNoyNYqQX5WT8mZfu+kkapiPE0ChJtiyzlZDUGxOAxm3/8PYwQx7W0jMNI3Au
BNciGU1HvuJ3u18G8HN/0JHkAmy8jtnxgNCNYaipRTVdBNj17O1Ohi7GjxieJLRq
eshyTHdY71fci4xg+XRgHU0Vha4Lfyr55csJIkX98ngDI/wP2YUiOkCDfnAJSw+4
mT7lY/COUYP6Bs1ZpVZUd4k15nGtynUyVxvk4CVaSi1QOtAsOMDl5nVmMgNe/3Pr
9pVoFGjYkj3WE4ckko7JlnxlIqmpIIfb6hdfAQj/Z5QUQJmsJXfoOxOqPY2lfO2a
gvP2uoPTmPb0mpHYa/yjRZ7OXRy32BFUTQNTO/fkbNntkSJrbpAHLEEFhknKZq7j
GoK0uIovu9UE6cNGuN8kFtO0P9AWt6WeBgQ6qyWCc98a4vYg9UYPFfAtHCOmfwlF
i5CmMPXPrxchYjGO1RBaJeT6KSoUl2nlxJLgUqkP/LaxtGYz+94BD4Ydsg+8Jj6w
yHdtLfahnPwzKXO4dm3sEJa+d9VbqGwuvHmsLJmf57yPyUxt84HvlypWM1y9sUiM
8WOJ3AbFeGsZjc0yYeoyKOT02n1OOcweUi+ynsLFlIk2U2uq+hDPsPBiWRtR+6vn
4qPqidGQw9izHYn06UirWBZG29jEvjzFreTRa/lQgf78n0kC0mOGi3/hYecEpA52
LgeS6TCSV6xUbb7e6eCV41UMDOXDN13JlotTwOkwXQMNYj6VfoqdKV1H0WM/5ebS
xA0dDmvaDIISyReAHtzxA9lKO2NVYCKQWf3+DLRLBhvS4GSQn7D8irPOmUtNnoD8
eDH2jg9mRr9BqLthbx/9e37tMKUTXzVftTzOdSUwCtn5nGVr27XqfZtrkj/MrSYp
qW+9ZRNHAl3F/tOpKJdRtkl1hCn1kuYfwQswEJXTyosD2JI4OxG3bti2eH8xB+8Y
7isFkLoGVapouK+tr9ExIs9HVjyCzSM2rL2Do1KZkddRmMPWBLkbiuhfvRFvr960
29xcG/l7KhEMZT1mn1D2YVNrcB9Npb4X2gaNjP5CO9o0UXPCK0AIxm6LGp3KVOsR
EWGiKeyyj847X7LWwRIjKUtAhdcdVoqLpRMi1JGkasK3WoCI2FVocjd9rLeoeQSh
B7OUFuU9LoMgtaz+WHo/mbBWtRzYH9rkYsZz7MPUEHv8SrUFHMiS1ZU43u10SMUG
G8Bt3n+V736+tvXdES4XDMpw0MWVYbr4yW7i57CDwEj/p7b+okBz+2lADrqmZGsi
ztbUe3cxddV10rUX/R5dmuPiMKmShuuKdeWSAzpQfeR5Ou+19ulo/kcRx1Dkh+8z
9ZMjkPg/lwKys5QCGsaG3x6AwlJnx5JZH80JLVZ5j6wueI50w4w+44/mNu/bFK0Y
Hzr7q2qrADqR688KjmsM2w0ZpEu34j8z3BPdubOqrM2RF/ERH3G7sbtT5XRIm82b
aAVNDg5W5tcPf34+pIHLi3YTuBXDsj0bJO4PzKMTdbSGND5o4ppBJg3ZuweCYMf0
AZrXN7hz6DVe5024GLGvnmYBJrxvOM1CKlTRanyWf6hmQ1j0FG5qndCjVbf52xio
UR9WvWICtYjwZ10s/6zLbLAOBSyajkLSrw71qo7bEkKUpkRRWUQtvVRvhYseCUZR
7ynQYsvqwcQLskJnT4ckfSBqvGc7CuATHHiVMdNbFI+EONmKg2o9IEvco5XVc8KG
MF5owJ6/khcZBvpO9Zp1DV/af2fE/sBJbVMDDNQLPwA3cPQh9I9uSx9GnMxZLuZs
gJ/bhIM/cpOUzyMWDsKBTHIGLeFiQL92j04L+YYTr9wqfPsMTcgxtL9rD4giz7FN
/yPI4ML/tOW9cf/bIm0KmhKvJyU3hFyx+qw+Xzt6uG5Vs7C/GvKAWgtJkdm6YM65
0tDqX1PBub6MMiB323Gk9TvHf9aHXNNLfy2Z+EmBe0xhRUU7ZcigkDEBSzyy9KXl
0KPRIrTSnURNIAdp3yJsRpNuyZPjGb75HbJaeWsygICMOpiuXz3V2Ym49P53RIBB
iN/4JO3QNw8fHhy4idvzFV1pIMlaw+6XKh68YxtTHl4RevMhtR/nTnH7dBSa+rA1
KxQ/BCNfW/UH8q4wtsxCAa07W4WEEtNnxGuTr+L9sxNyJyqa85buOWmFeankIPtF
q6Vi4CJErI7e0EnGetyUxjlJ3gQRJvssIlUt6st9fXmjsnncJCuSO5fnQqwM3aLP
KwcI6JsgLxSv0GhofRA5EpGeRFfdblE9SJd2cvUt0g4j9fGrXfN48sI1qIS4TSnJ
FU2kudj7lK7K1yDycXI7c2SlaOqy19+BUW8iCq5MtONCe66/IabaNO8UOcIgy+7w
GD/wOadjM4bhnlBwTxdMCeHM6mJ6+mVxEo7MbuMbFbWigSklr1g96QxHoFvwCfpU
ciLxAZVB1K9/62gJxbXZE/hWDTc8GBl/1Yeei8s8lZ6Oe8eIvXA7H2HccwzaTJb2
RjQAgWIST02PNlNfAzUfHtwPbgptJxuYJ3gn6em/pu8WdgZoExmBzGyoKCVib9kK
U7TtZcKVORRbtzVfLT1bTF0e3vQZvCQAT6GLdaJTrMNN/GgCJI1YomBkCK/7u1o2
q9ywyoj4ogQddZMN7yv7i1Pxm0XQRSyMBXeLvXMuWpB4waohWI/QIhFTb8upAw2E
hYQEmVxw5LDqZDlfNWKzn8AZS9xldDOwns0vOEY49UnB6uHuP6en1lShDW2Yd8bn
1I9sKLGvlu2gMpJBGC+pizBcNwcz2Ru92nz/MLANkrzgVDWyF8u/otGbI0MWhT6e
Z53K2b1ZDGSynicS4bSaQ4Ha5mP77SKw8Pv9DD2LmrtWiD1g6UH3MySYr7E7tmba
wa4qEsR7kXo7BFBTSrJxHVdDgH+DPjPnAdHjYFYcJ+2oVlk+Hf9ldrM5T72ayBoj
QAz9JTDeZ/v1xIamJn12XUc1A01laMuYRlsH2I6nrjAOnVVUJyUQXpJZfe9FPFRS
9fYt/wv7mcYMZTopVzbSEECr17ng6eGREPxoV/JTYDVNnwRddBFiZvhTU3SKe8T2
FtwTHHEKtvB9LNBr1/De9SXurhMw69WWKJ5QcYAdUX4Q0ovsgWe3j/wyPD58ylMR
ySRBCFapmdzpJvfY0H4H1gjzaQqXVwZ6bWZv8HCv/H9X1oIIBCSHfTx/Jd3KD487
xVh3RPZryqKh1MBk9ooo84oPs1x7S6XIQreAeEckvq2nveU2QqWL0G2u7XCJIwlL
YdfWenP7boGsv6eb4bzxYSOgC0lJOhcbRvKhTnXm+pWjxp0T5Ft3wJR+UEKkIPVS
JqE1s4kDB3GaZvj1ZK1ySnCka3IH6ku1YtINI2oeMaWLGKx7WY/bH8zLTb8Y5/Dh
kuIp5hxUsLCkZSK/tpLaRelduRbmadp9tQOu5jhBCxxfWElvTibsgpZ9EYKWq/m4
8I6hvQ6yvK4ssqcvYWToif+UsaYvYtqJSteYkG4DM5Ge40JUnFjnnOaHn3zfkq01
QwiGHmrlz6O/ZewP7afSlSs24Ep2IC6pbGLUOWbbBBX/qOo0t/eimkD8EzAgfaH6
NUyFqu+SBncRHtkvOOKpYGvBieaPB966fFkPG+zG4AMuGFdFKENt+KgM4UmlhS1n
HpUpLc4yBEXOU79EOZ7PAfN4KH2fX81MFXgoN3tqifMhvUqxr3R6n17AqevnmzLz
IqB5xIjDxJ3YxvYgwQNbIMFOjAxQZtXuhKMJz4Dp+tw4Zp0spA87DIP6K1xCzLK8
A4F5ObVI6xOd80ataTuKt9muFUcY84zax2MpEHKdT65zjCrnTNFP3wwP6Po8MxF9
1yVGdgI4OKdAxtEg6t60dn1O/AogaPmfc1dZkN9xyZYktC2i84r6+iUxmPOE1WAN
JfdjpToUCc43W4aJW0vUYGXuK64WW8skmhfE6lSQ2mFpNRBxxLtZVCjpFqO7mb3E
ujKx0ovAEse3UhQiSeETbvCDQvjnZeqOUCRjIXJyIFR1ORlePjshU+waaIPv+k04
GGSojmgEIAIbzYya6Nq3W5TNCL8ATxiOTdUoSd7VUQcsI7NUJiCA+WGNZeYonHwu
6XbddF/MMXn3r4SabctHTPVMmFxoEjS9sci0etpvsz0iZ7U4zrCRmaKqxQb2NGMU
GoaBbYHAEjaQErK0kVlwogtOm0XMldfB5M/W7cOgzm5poBus3+U6xx1GqBQCLWQU
UulnwgDXpgIIJEv1MjrL+UzqUEBKxwkimFrLj1UKd1bqGBRcNqbjyR/AggiUcbXU
qQ6QVJBIMFvV89WiBdhs6HJOOTOKYowD/1HKKCxVEon1/vvbb5wKoEExF1yJZtgZ
4VmhG2wu0RAjg3u2Xp5kght0wSYC4BCpyj9uO7RU23GuM7BhfFGD/R71+jiRQAsB
ELA5vBSsXR8x2DgdwBKWjJo/P2fp7hbT3vp5L2o6b0PAkpGeaVLfkf1Ho0EkQRUk
Tc2fCUs15D/WE5ipmGHivCyGGOeg3d781IQLg2NHtrHSFxlxB2fEr0HFEm7F7aZa
U0RS8dQksDlSR+AEvIwpAH60xatS78AvW7S1YRLDA+K4qPgn9AG5f5WzR/Q/3YRV
COK3yVHJ1mzbuxennh+dcqSW848lW+GGIYr0BBqDWDzu0gdutze4hlpv4w/UDqaV
Pgtx9NZjVsyamOymWoOgLuTg0ltFJtSU33KaCCeBpLYf4eQjmNiLudoYbyjjp1tv
pLYltRfPIK/rBg3uE1aJ2q5C9OCIrS+FWDrHBWr8SbF+/f6z4t+QIKJPOwwjWPOy
b9NgZK/qnyblIJQvysQuUiOk0muof8BtwJQ4Hqr96ja0DVhtFri43ZHMI3gm6mrd
bi/rDX/FesALwb0Fc2mzs8U6MgnPXamy55NP0TbV8S2c59AxiXxY6Jy4N+99fAhF
dbU+Yr1dSS3LmGVpCmPEWHAhEGIf+E+4e7wgYk9SYC2cXzYDcNJDvJwI0wp5WTm2
P7CKL1/JCj+nT92PzcV8YUIqZFuCjUb/nYfJ3tmJZC2l8zv4iRHGHy3KzAJauwQy
KGmtxJyZeF67bTadqxII3CTL9fMNvXIt58xzR4C6qKxohAoJuObCCiZ7tgXCRLzO
O3CiwxqncU4UGuX2YG/mf29u+nc0pgJnaBxjnLxLmi8FpMwYYxTXJeMl/sDFeZ6q
b9bgbHf8oPl+Gx6UD6zkW9VwtvVGbnOkLBM+E9d68KfEjE5qXKpupxvZF7hpnJH5
0YSamZwqgwID0OxQW7OTpd0RSQaBxoUG+phcDhaY4K+/y0Hx1YEX9hmckBxziiVP
oUzrveWa80CEMkMwv7SH9TlKwMt0QrJ4Rz1wRYuEZDZSOKVdTwio7++8S/rpbf7i
y1c6b79DJheBwJoJek1l8d+jkjYkGKDfAqKCb1v0koB1vVyZoOqDNKVdZRHZBF1o
eDmChpoaVd/7bbckbhncHs9gkgAbKtl/A0jvxOO1h1X5i4Hw9XKdpAMi4ApIAF3f
dP51VNSBCkCPKgLHaRgV+53nWex0zBdFMmNcMSuGSJ1MOZXR6H6pN8h7MSn7jV+S
E1SU0up1TXJzzZ+Tx7JddPja6KqBIJHvi9A4RGApsaLqqzfVYd1cuU1UrpKfwCxz
IXpqe2o/cP9CpgGEqgMdybAUATI7ik0cfTZU6VmT0N2iC5Ang0H6+FF5EBfUwZkr
WhLLypmC9rwTJdL/x7mV469R5qWUgMGIxhxlZ3iM2vxQWHPCPbOlivBpReq5wU4d
Nj8ecBDwFTIjm/8syhqkV6NjL+EMu3s13sMWzgdkVSZCaUh30orTiv80I2LmsQbG
6j/e/mbjfemn2Bmz4wYgyX06WsUy+U1bg6ujqbl084/8nmUfe5QgovBBsPJP9ARF
CXV19IQZaz8DrXIPrWf9zvuHSJJbx3WzLvR8txQ+Rx3KCXFOxVIg8uPCMAL/UGBX
73A8gdOOrR/Uj9cjIAvcApThbRwyzkcfnYz0U/J5Q+iWbiqidhSpQnliOlxY9fb7
U1WTJulkTqpwlSjZCJciZ040gSxf6i18v4UzdAD/NaekcpPOuyof764U8z2PG0cP
GhtyVcHuOyTOFBiaxRMF0TDIutzQzVB7OYaqG+LmofW/RZdq5zvgYfF9kxZi0D8k
EuSwl6e+aBMggSkV5eiOxt5JnDX6MQSgdeC/z7hPyC+uTWAU6rBSDzeco9FMNOsf
eLBJRHF2x+1+PaoasDqF/kQfroxZn4gtofQnKwQO2QoRPAnwpNcqXcU+qBeLzdLK
BI6nfi2hdl+/ebuUC8f97NDO4wa9evJBQPyk0SC8ipzLByDNMz9Li5fuj7fD7i8r
23c+LIqLEqy1K2hrYRjKwOg+0qUBUuO7gYXBF7vvSSEJysyOrB3J6bRmUh+ukCOK
c0u7k08nvwPr43DeUjJ+sz0apGRJ0TUG98Jx2D6bLyulPcO2hSdPUj6mfGX1Qvpg
DaD246RHMYfZY9pvC18eTp/AXvUW4wj/LgTHwZj0dhMHp+qV7b0nsJg3j4gkaRlV
pWjH9VJCMya5MXKruCaCu//T6YRLe9ZcEMBuFvmoljxK8nbChYj/LfztA2PTrJtS
daGXykaQwd/rAROjK9StohKnWB2Ph3E0Sv85gLVgzafr1SkD1YbGPMWQTxdqC5Ss
+z2dYww4EwQqMI1l4hIiKctf73wQM4JQ5O/V67c0AiSMu6GVKRnv2iL5PSlIrx0N
b/4XUzEgGYOB/h6kQ8ORlKByZJ0d80lGgMzNOJFUcw4OesYn9BuVolWFvXmoHFHF
QOgKc3LNrR/wvRAW7PzIVcfMoe76DryTYcA+DhaTPybgoCB4smprtAj2nLo/sSXQ
nFiT4wv4DKUaud84QDJIhMpHC79+fAldPrDfQKDgqdcfKf0RqtWKUnImWEhVQVOL
XUrjHVsYcQXBfM+kIpjF8qUsu3k6m2ZiBW72JRwAgy0tW4qTpIN0g/DOtkHOsmSC
Fat+f3soMGxID1ExVOfm64oBQpTxwBT77GwuroiLLKTC2zTVJnPdHenBVnuytYOc
CFA4T9R6qFZktTMIUXneW0lkxpgpSpaYU/siqLInZJCytR2EcvVu4zcCIhd4Mlue
hIwxzW9nZDvLNcb8qGl981FfYM9K39kL+PU1Fu7tL370TlvAERAIdgywd89duN0p
C16dWkf2ZhjwxiWc1ZyRx7vlpMkfOT54SS82W1LkI3GVDYBiakd+LzLW9igVZ1HG
jP2/LhB6z+sL6cRet1I1UX8fFaApw7bK5r3mOl+m6eptbmZQpxBGx0YHmT1XPA1y
sM325e35EEm5fnCA6KgIDEuq67KD6cTbalouR9/epYGF0tOEeuuZ+YF72EWQphKV
TaswaCyfMF7KTwepC1ePXz1zfRTezX7oekHA52cXZMqTeX9gwh1N3Zsag1o5ZKoF
bOd4G5f1iVVjfjFu1Je+s7dTGkJi3tQtK/PiPqF6Q31jIkAoAnHAU6LBDSmOvxZs
0j0iXNizmXM1iQBgMslJoeurJqLnCculyzApWTxolgl5WRPkQrqSsIzxozOJH5sn
el+EsOgLWbpqjahssHAhHiUWNrirZYiM5gWIx8jZxCQcXMa9LzfLQSlh1h0C1keN
WLGKGU0OozH6AzHj2Bca3HO0s31SeTbpKIu/5WdTpoAT8Xv5thZdfUGujNdeD6V9
rfpSFQM8B6ufjTH/7c85TXvdmD9LZUkRltKLJ3YGj6YRPveaiWGTzKJ+CaUIK8lL
mjSdlYVmJOVkDx72qLZzNN+gaXdlTLXgBzEUG+IqHMnS86gCDdNyLbvMjxhU8YST
oObpiBJLxm9QdTmAGsaSiUYp8VkaXY22oX6IMKAxNHzK1Luu+4FWEs/YRwhulZvS
jBIcmT3lEuoOvlA6hP0SLW3wK7ozXmlpxxYxGb3D+S6hns0Gdb3+pSZ6rLJkYNFv
snC7kLepfmh6tnAot/fUb7kTT7oZOHvT9vxd7cyXeWNOO0qvscDso8VGyadXDRKz
i9WQBCXq8KBXXzbeq4SkyThRfi4IwX0ylQ0PVSD9XS7x0DFxHrPCEzEymH+eql6O
wbotD1iN3OxpST0dnzDxvFBV3CEC8Sad+xkpKj0ySBUEmZt18SQpLqwNmjZnM/bc
6IYwCXdBdf9l5cJxYv1YyrZDlbxS4QHm/3XPg3nVU4i5yzrL7kvq4VX8O7Uk2Y2K
4qChU86kHUzCpv9XINbbFTdwDtfDhyuxfQ99bhgoB+NDgO1dBGPEfyjdvMA/ytUK
HaHHchEQRuUrmz6VDBliS5/S74WVTwBugsKHOHpzEif4ubxE6NoIVK8NAsvus34K
SV2545mi2URxmYC5wgQNqK6lWdYBC1alKCcycvWNuk047U6tdhGv8/y/iXEAVbMM
m0YoMy/kdmBbfr4EZX945jZYReMTGadl+W3uR6/D4Vapugcd7IC79FY1pOP6Wqiq
ZiSzOoPVObW0ztAL2DrQ0fT9SV+p/IIhE4BBKC0qsRwLoRY5gV4ybMCYEgteKK4y
N4WFGZzAnA4FGL1+zuLKE0nr/9+Sq0bnAK66tJ+RnEWN87gVHtGl/7fwzDw3pXxL
+PbxrNysD1Kolq/KDHRphBCD9oL/DhcajZxr1ANFv4u7Av7oZvCd8iMfux800h3j
XzFkafkKk5c7bAPOAFFBqUFKCO/PdDc4IPgaaLCiXJGcJs/aXiUfxnplc8A+bpdH
NMDJAd6EBaH4t/Uge/AI/IGK1dTlmXeI9g7jtBd14DAhkQ6FVi5guUQbxoypVnHH
h8bRNhufrw97vs8gOHoVpugghEPlWrZpqjkoa5DAVjpCsLBYojfugbfPlXKbV1eF
buSRe9x6XsspsvxVR24vTFs94egWfdAFwDQ9C3/pp7eC1V+SVWYcROfKUcxXIWHG
7b0vH4nnNRWV4wxqRSdSVAwpvBxeJNIjKzzMe+Dj+J9caHQMJeG8QxP4nimO5wgc
jQbtwU3Sw6QyqiyO750H5IgOQGokPW5mavL76fUQezFfJ6D3CfGqua1u6dxQznMb
eCqqGhZNMi4ZQBCHyJrkXZH4V7qO/z/qNfKQNlxKvBLJ7skg6tdWvKGLw9vTJQ7t
0fDZuDIRmYpPJV8i6ylA5vtT56fcbO6cYMD/S9lFfZ7doEY5Zgd+VrNMeqdhYq89
72PLg0fWW756o2Nn3Yz6GLBmnBfqBUhfNCqj8I2LMlACyDhg/fFi9ERsRmPVeD8s
EuXu7rBLjkw1u5pZzQFkklmVwM+ddywkYsks23KEN2ptrfmjyEC8d/RkMtr21HLZ
palZg7pOK2OLnO+Jikn6A/uxNhe8Ab4vA1BDcSfcK43a9obSNWewSYfEnGigLvxH
as74hUjZcTI3+ZCul6AdakZHZH+K2oYeg52EeewxsHCxGuTBzGeqNUHAcD5UhFyB
VCWxPjgaKqWOkKDnm6ki5+s2U0mx1dOvZP7v0ujcu/hNsSaQvDCEgpHMNf6CRimC
20a5+x3eKjXhQWdj8R3LvoZycUWLVfo5Wyo6dr6DHRm+xsuFaO0Hkv0EOCvrsXqR
RMWZCcVgMBcHA5OSa1a+i5ewksoqpGM2Vsl9UB5VfmNK465ktrL0G83Gdzac7b+c
fgldseD4Il4L8CHZCFHN47wUxLIb0MDynD1YkPApuRmVfdSsyM6qjntK+8m8jdRj
SlMwDLl+ZgLuW364z9D8+ppq6+93x3R7//0+f+OcrlcjSznfphv49oUs7KpCx01A
D27rxO/vG9nsiyvGvtv1Yn0jlAIig7hret0+eZAfmAp9VX0hYID3rftxKwUWt1J9
1Vb0zmo6YLECLjY2iYZvtcAY1LQno2g5A85VksjxFlAkIlQfSofSwA73jF4BSytX
oGzNV6+fc+3cVihbA7PsUutrTWa/ED2BDVyqx4MvQLvaouDc87mCGxdNxlTyxgxm
/MqH1llfosUtL92+JOKZNWaIvCvQXKsadZ2x3WumqjhMA3FiPKR9B0EcmRz2Tyf1
QlrG+uZvQhMKA96gXqNDpc0j+NK48HFJzhv7esnNdNfALHRF4FWWrS2+M5lFbOM2
tzNrrweTbunv0y5ENhghnEfN+r0wTg01vV/9uwKMkahpgJglV+lIQdpLH0jmodMP
0v5m+pTIdUMCFWYqvg4DJgYuDdAfgEK64wmRkFkNmgu2Vu7QmsZqpBYa3vXFIChS
nmaRctfUaI/3EncPk5dlGY0evg4V+JlWuSOXfJkseyK/kTlpb+pAwHFGSLMeVNQN
z7dv4TdAL4MtYeCHozbQ3u6tgN+tW388ry0+Kv6SMEqygiARZFWHn5ga+sEThO67
ERje/LKX0L/oW3LuOgnvEardZIRZye2eIGDLoPzIi9AGfxf19xsQbU2fKwUsboju
Cqt9HFz/25vmmXVFowav3LPLf6nMnbPScORj9CSehB6gfAqOcjkaeH9Xsfwh7MuY
uooXW5psRTWAdm15SoXuA1rhHa7gdiJOVgiBE88p00aM/rUe4fF2V0z/W9X7mViU
ugyVumnQ21g+U8sCe8QNZP8enHjGV3J0vMqxO10N22IEovARvjaDrkCNr/UtqDjf
Jfh26kXyEro5bmi7GRDhlbppVF8myKkuUowuddtYTGd7+gQ2P10a+FbK/E+dmCwT
BLEvd9W7Q8ATDGK5RCHO59PjRclaTn+yHk8mLh1gQR18alz4Tx6az9AoJza/ocB9
atQeNQ0/zx2Wx34bGu8h/WBX8eQy+M988QeLBY6s8xiG74T/4Imw1YRez6j524OS
ZXjpW7H0yJWUanbrlv91AEBFIOGL7H1qyO1s65NhucbXghRkCBJ+32f156ov4r7J
LK5kX2YmVOujnNJMa45aiZY9L97n2w/Nz+YwcyMBqjJ0u8iyF/ylKVL3odBiibs6
8xC4njBT7rbTJ4IDRi1/dSsAMQ4i4Hg6kkbYPV7Ozq/Ivu05LHl62AxErh805NBl
ilQp/6s9l35SIfZ2IGMGx33tpyzp+Qj4yw8b5XQpsceEuVSUqALlxawLXcIHWozi
3TGNDD58M7cKeQRKNUlZJfQgqR61I/H3FprWNksRc2Tl7rm1+9T76HW0RuU5tY+8
aojzHNgYF3E4i0fK04Yc4z0olOcb/G6TUgWfMpRgle4CMoAB+q2w/m5xSKgGwa5G
DWoqCtYIMiu9OGCP3wFk0WTZAIet10d7RmdzdnjnzmRhk/kNh5S9ET/Ca3KKWoEi
40tSo6z/UBzblNgXFIQFQYVAx5DHI/fETkt9qXRQztgvzVlb1GGidYCncXcZiIyv
wKrVZoh3BSz5DvB72elUoy1jiJOcGMX+2sTMqIV1LOoMERe2t34EORVMU07qw02X
zH5Lho4iGchZCp7shDzRlrJ79rHU70TVeOMpA1OnB7A2uOlehdviKP5cxcOnlrcj
VLG3a6Zq2mF3M2RhgHjoDORrpRqAITIWmkUdKaWSjBe3txjtONZA2ki7PjDefj4i
ISvBdBqILbyK1L4dQyrnOvuSrCZv8vvIzQcYOD1iKP8DCYDpfYEPXV6NJMI7nqwV
ji7NMIRZOBhWur5S4/cyY2BVVY69odC0du4lSqB+ncHmeYhQmY7nl2BenRz5HMGI
15WVYAmL3aMUG0AnTZotmLlm2SvFPvC3nk9bHI+Rp/o/Y6X0wHPPA/5ZpW7osgZS
dLxi/9ZZoe6smYILZmN/Pe/s/1abi1zQnXLJfjsz6IIfcWq+tFbs7gmezjAsZcql
riY5RjJGvOGoudo67NHC+RiDMGhSGeaiMrnKvzk6LBxA8YJbxT3vqN8oUFxkawKN
AUs6PnZfmJGQwiwvFrowgbU/vByK0TkKIk6tvn8P8WxTEfzQHGGS+CuXdbqIeB02
YIsOqEcsgMWoUOd/nyBlFN4tbcQizCP/vhjVKcA/tmTSxReRe06K7A3bODrH7WBw
X+aptHAIIAZ9tMzALZziTSWH1KasczCvwwrw2I7UytMTXmZNFazcTz77wNaLWPwZ
ZxwUk18CAjEPXN+/r+MbPass8V7LdmlNGbju1uGvz87mtkWcl+sggTcHAj96+Q3M
DMDxkC+OC6JKf4q79n7i5Tj+K+jkwWFqOTOCJYXQlsMvvuVYCEOROhQC+BZZNi8s
i6jwVZn+HSE4UX3kw2iXJOM0k/zUzpvBsxgLkKF0mzA4HW+9/HaCE4fVjb/Xtfea
+zCkpZthpw0REl136PyoGkJdFrAgltnn98bhevmmnhkOChpJpyPKrSHp03rbWiTb
FijxAbtb+51UiaZXvQsgSFuxyFznL4n675z1dAOKdCGe1eHbwxN9bOIZrmJoqY23
n7YSxsXqH29kI92XmWINNbd1opDFkeFeTDzskp9XgiZJCgWrZbw8KGpPv9eWT4Xd
mQuL1vLqSqbR7VtLuN94cLLv56wG7/Hriha3/wjRRp/cLSno156svli10FXtwdya
hM1h+nrI1zr+NpF3jSVAYwsccIGyhMDd9vG+W2SiVN9mNL7GwVg9W/NvX2uFcras
4CgOl/Bhhlibbb7LdM5cvAzbm2rnecJ5D3R2SXg2JBRK1egfxgDiu0IuMsmG6uHe
KWmNbkpt+dKzo/N+dgjUDu+tRGnsY+gbszpkEDW4gT/vJ7Qe1vtBVh2GOxGwyTer
r39kZGxXJsztdNyjbG+99v7NT5iSxIpRxLb9LwYFS3vINN7KV/ttZltgwqGp/uFJ
YaBGgPOv7e2AyGfew38NrHI/AbMyhseB7CU6qc6toCGUbRk+CQ3OYAZLbLINk+Wp
a8KCgQcJ4VFfGtGPsehoSTFDEj8td3jnzQRb2bI08al4L4MqIMIpIvJw87VBoPGf
y7JU+dDqE3UJdVCO6uwzoMJrso2LA36aUOVk3on+xJdqOMvUasenxb7R1/StzJXJ
3sMAjgkekkhv0KLluxBGN7GopwUnGs1lLlERJSO6WXtLlRBmlWVaC9Y5tRWeYStV
tFsQ2y65guiIMr3096pmZV0NP0opkJd+WnFi1Tk+I+TRSYzx9yW5l5/2515SikpQ
ned0MANYEvPZyMSuRFHNwGUXsx7MBD72FxY1MLdwwg+IOSM8/1d2eUBAkrmZFLzY
j/8dJ39oft+v5dlKYbCu09S+oVV1u9WaSN7lRI1A4RPMnufmyOqMk0OdcxeNtyEW
+qiQkJ6iyYQjBwTH/eGyJ9OMPPZBbkX8g12rCilvekWi1+Sk0Oz2xD0QnxDwXShE
NixLbuh1S4qdzIZaAY+ZvBaPMLmxZ3cqWHhENVGyqPAzoPj003/hAaGb5hmZG/vz
YwxDvLx0D6ekf0OB2Iv2lmc1BTl9XufwbpneqrowMJmFdQOQ4Iv4o3O4BOUWX15S
YGk8OVFQSOKqpQL87TpQFXwqAo4djwK7gjtYVLCCkIdktWy6mdmalgzDcsrbooy3
Yd40a4B7H7RzNokgKo78UvD4nWxRbVNXQKNkzisVgAwL4HoMnDjeOE05ZDlMWKKS
C8l1chL2QbVCMNEcGrvJgpBp2O0M+dfSZScMCco9nfxCcvWfBflx59W7oddGEyao
uVLr2UMrQeVGaZ3+3VdSRBpcqFrBDK+wJt+XLPKYKNPyZ/87cvsPob65piaY7mST
J6QfT3rIrGqCVGTt8gAR8wkuWkc33NBgMRjSVcvodToXf2sOj8aZluM78P0s/+U2
6eLZy3fA+vwXaR8LLg1BGlJYKtPIY3iqVqrdRF3UbPaSWglGg8/cRey2OsOtcbCA
c4fcCWq7zplsUol/i6X/Y9Ssu+lTluwndnLZQZ+7RW4FHtUeKLnuSF5JC0rv5nkT
F5/qtqn5DXq8fXqXa8L84YqhDzixMOzad5Tk9anpSr/ATq4TgLstC4G1ms2o4szW
jYsMRih9DgdKG9bzhF0v56FnW4hgvPnC+t+a6c+HdsEioLgeDZJaXmpyYkd/4ifU
uN/RFxmxXD0+VGQ6cyQeIA/V9asYnSMVR6g4yPjiq8C1NfaK9M10ZBKnsOKTv37f
U+27sU4uDPOxgxM+4Ryhr3TdhRLe7fPTu9CjkoUe7x3nRVOySDhDJySs6TeGwZzh
UD7l4GnWsyemwpXBUpxBEBmPzkjHaFpZlqLIGJkmF+5DnrWpnQxDIO+Kqan9jo2K
nD/wIP52i2yqZGKtrxEPME5L0onK+MQfty37Bm7f0Y7U1C5EGFB6aGCo0+H+V5RW
Swh/lHv5EJCIB+2mlAJBkQidaX+g09eKFHn3oyx+LdeSJI6GtJgtBl3F9gvmM147
UFifRbuHwY94RzvmvplGHQSMQ41GDcMo3Sc1VzJOLTbGDLTwGjxnBZ2vW28woUcR
3CDsNervYEiC0exMAcyQUiql0QwTCFFBjfrlRYRosw2ClhOIqZtrlIKPu/Od/7UQ
1vdmXo2r+FrVX+HnIml8VKrprZWYymf1SIY7mvJD9j7coXXg3j5x9MNx1/j1f7yx
DdoBW8MUfFIO2qkSiMq6fVmvk3Ue781lJsuW15VpYccTPPA5q8Q2fkgBmSpAHhzw
MXWT70u8OtJQeHbKa6Ax1LR7uouh2iacNWu+qoZbeK0fTbaSYunz1e8yVceKe6dJ
AL++LuMrHO8tEklqLuPQoqd75HHJe84H5VaCiXE9RZ/KNwAxjTCSQOgpSQA+kK/G
vOQs7cqUJSIlwTXqIYUjZHsKsUjbC0y9C3Zbp4XKbdRCzf+LsU3suOSr1T6zyqJQ
dXahnDTSrI4Vd6LqN6eYqItV1V/t2Y6cYLp2lH3zi8qRrb3sT/+qYJpvqnFheVQH
cipnHgM9lDA3Qp/mSpXnhoaPtE5C+1K/FuaOMw4qui11C4+Dqy+CK0BTd5PC+Jk1
Wl+ScwWhFdv+ZUCjWOsomiLcwxDW9j4vCuhn/w/z6aFATadg4CL3WmuxbKVRlO2g
ZXl2zUEexiq40btnHkdmNHHwdShVir2qW2wCaiIUlN4/Yxoiz80exvncRR1ZGmL0
V4Bn1XCLg0VZKGri/nnE3X61yIxRTFjL7LNZRPmVS1kurF/hvFhwMsUDwpWzENVV
fZOSkbHul7SWHtIlFbh3SKxmV4aNb/VdrwozDH4yjKav99Hdx4ODhjfX5JdJh3VJ
X8PrgxOPlJXxV5gR0ECvN3pD7CtAhWI9DW7y0/zMPjmoDZ/fRHB8CH3ffKf5wMvC
uNF7hJlzAleHI49YqIv46Am4ZFONRSadMH5vYpOALYC6PV8mSQFj+vEtG1513OIT
YjrabUod5T5tp58tF14cfgrjp3/AVJZNABdRtIorLHTu3veDyRkErQdpnUvXCe2r
jX+mvOkTmdE6bPaQnvX64cz7020h7qSdJt1MfF4vAlhTyUi0HzejRmFSSM12qamJ
q3ePEdkbEJg+i7SG9TWHbs/KU1XqrLcPIHkGzSm6PiZG1E50p5MUy+lpaReAVhOr
bTVUVeiwnRKw2CCeohBOx+iVYB4d0V04xUhvqLBHJoD8HrM1bKHeVWZMlVYqQ2uI
J2dr0uVOQgoEMygb7M7w54cExWpDy9vcdc0jNoE+UbrOb33oNryoFZAxJsPoQBLQ
6wg6kszaMrRzXjaNpKKlstn+T6gGpu6MccdoBLIKYt0tQOM8zuFkEvYkduGCzmAl
85lA+KTEZ1BjBUfH5GLWRnOI7iSpXTtOlPhjpQLZpM6JvwR8rjmvqkl50wDt8sBX
/egA+nTb3PtqA3VD9inxE30yMRpkh9DBt3+p48ns9ebbogp/z07CJx65Dfbu/lpa
IsowozElfrZNmjWD3KgCJxNphw5dlNGm8qI8LAFyDrN5riAvX1el9c4qKhH/h+16
uIy6832mkKgLlQ67igHfUBnVY4qsQCMiJM9GtmVVQKhGVOQZh3Ejq6mor9gmu3q4
h3dq8PWTfQfuLsjQMVGOcaN47rTojt+tlLBLeE1cy/eYw48dVJOuTa+dYMx+NSmM
zQFonHmFmN7P6+H35muc4T7XLW3LXUzDIJVEz1iIdZfNkJ8d6Di8Ay7T1lbsbYsW
zi30i95j5WTnJFK1oOGbv3Aene2eOrmjepU49Wg6WY+NkuG/tciBYogX6MthLsBC
LXBx9VUO0gwvlo1Jsx81LVHj2NvzKHokGWCTBwQkEroiPAioY/n2v8uQ2N2srulC
6NJreNkbq7z4R0XYoKxeSYnxLTXdrhlHqKfycFazMZnDd+VdvKoF6PCR+NhM6wFH
pj3QXd32TBjSCPty9Vqxc9+whXiVGkK3apiqWsMdrrrOd4CExwaB3YUzCyIEEEpg
A1oebjV7E8tGjwAafZI7/hNcjOAIa9KlERVzL6z8/rftH3hr5I/9kLCTyMZ9EDW3
ANk7LUb5McBbwe0ocNIL7lun+wf4jnPEu/ZOsZC3LiVpjjcB/z47fSh2zENTDFgj
YXj7lWc7+jcBoACt8UuCzBnggAG47spmqeih6jTC4h0x/CH+hX59O4MQZ1A6bz9L
73Oi5Nl8DahH8cK3MxSrD/AkLRojL7wsY0iijRRB/4gFUIGMDD09HKGie9E6JTK9
44VMttxOOXjXMe/QfBTbOm1TE6k6yUC1sXPOqgDYme2mX0Tz7PEd8jrjEzDzZuaU
fON2LX8ho361tsCeCs718yvnDCvFa3yWEKgwd8UlMOZiCPGbtTs1HqsMKI2LVe/V
1NWKXz9R3n0m6vFw5Q2zbdF1b5XxK6i3OeyOkQCj8uSz5cszmWKoa68/2vAuHm6C
rzVo98eO/J1+GXzRE4SGeJo3r1gm3NlcHPTBZuRVi2GI2hyQW9mFgnmTnWNzbguU
iqYOY6EQ85KfFqG3RawRLiMNXNusvL0U2BaFbWEPR6t1XDiOwxLqM42dZdLiL3Sh
Ateqq5GjiKVFF9yiEV/nECUlFuIskf3yJ4F4K+NHUJ/+mQI8/piAQhCXj3KpUheV
Mf6rXwjfFfzcN00iOxg/NtKUxL9hyYm8GuOfc+Z+3IGb0rBJUW+pFiuQeZ46rCVt
aqUi2y9Lb3hHDKvxW/oE4k7M1S5TEa1CpAF7pA/sg5eUBcjrbmq/UlkT0SWOTtml
d4ayYoFLWP3RuXSlG/xJnEsguVFxJxpywLY5FzZ2oNuQ8uFUH3mijCVnTMvibuvl
z/cMoagaMP5AUplGg50hXSt6HSD9Na1hM25ehtFsMsy70WYGKMq5i1pfFfJpAr+b
mlMi0n2/BouAdMZUESKz4hffg9ekncgGgPecgnM90nUxo66Zvt6s7Ki9HB0yCFns
H1l4I/e9zz9dHZsMnInUHG4gnTHmtHCprlw1w8hemfJ7iEGE9Ybsa3YTvbEsJoqq
XgLyHvk+RybbkCsgGCoHo83PjLcFq/yGON22OD0s9JmQcNgRazzxDGgYWwiZnE3M
i5mix82Ppd66qHF/jeP0Jyc2rRbkg4/hZthbZlYQnz7lxHNKmlQh52PhlPJT0uz4
GNpIQkgtC6guhr+1+1uh4XyOvS97xLpYSY8ILuKARCNFKVB/MYw7XTgk2VYweTcR
R6T+odo/VT5wUQkw4HVNDHNfNYiQL2/WgX+UYLhmzOqFS1p9xQlnMj/x8Kdm1Xk1
XaVjf5MjHqg4P5wAFS1rt5phGaErIRaaVTuUyjIzcox8MWRa7noJyuruwpjm9yAF
J+42TjfYp2P44zY4Y6I5L1UvNZKwzqVeeUxILhb50ZvVGHDCBwCj0U4c+Pb+Dzr+
SHT4YhsFVneCVu33mMiljfEe8LlMMNxcdZ8tK69i8ijh78Ooli2oxR9Et13Jpv0N
ZNIuwL1Hy9sU1Bb5Oz7bk3gMokQKRJZ+FRPeQSDXffHH508FI7BXTHktLUaybotU
3Wi5gFCStr+pJVPue0OUgKk3LLhfcsG1LUUWiAn7lbdYAqxb/9DwObFreMtR3oH6
EsLhmPsO+9fTORBhmJFwrpeHsrK8dkRMI1t8KBsOhn4v1iVV3vss0nPxDacRvmCf
3amqTP7XPjZgSJ3sFyj4skBzKDzfiS7RPCSl3JcJTlAIMgKSHERbKkhotqgbdI4T
wiKA24ZKAuTrp1IeR7ujJbByaFL2Bykr8H/t08zkgTzTigQQHz/v9gS22BBYNi9v
T8s2rAzH8Gxg7bpEIp+FOWrHbcmukAnpwTj8P8Guai3RZo/JPDojAZYnJKHaRYwr
9x+ARJre76TGbogY9zUohW08e9u2duikeXZBDoMBwA9A56DSZvWKvYe07aM9hCsm
oXlme+bnrpBa+MMsR97O3L0G+JTbLiT7RWWM+f0XtzckC9GmEiRWxAltXhrTwdpV
XSIndvPzGZL0kqItYYUAUbJxvyondJBvzI/W2PNTw2e2XBIr1uCPMdTcWkjG0q2U
TapaIri2GG26t+jW6Z4k+NVmWLTuePLzIf6sJzDsKSv+EHXY3G43gbgJtsBGZlnl
FvjDK5p4QDrGidVjxICA3PtDgQtQ+GD34aWymlXh1Pc8LLatWnwRSBA7ltELR5VE
reasB8H3zxCUHTGUQXd7K1lgV2vPFAsnETzjzB1jdf2tkFLNKATCHff7tsaopCVA
BE6EzWkoM89yWoOLk7tlpZKZmyu+7zrTXCgvb+0VTUl5aRZ2GwG+GTjphy0XZ2Sg
bL8eLCIFNMQmogHeQq5DIITipvKYJnzqBYYqInmBEV1FyioG0K5H9t3kEAb1BBPe
e7O3uTsy6TJAlcrYCexP72A4JQEHwjMoBHblB5Xuh/n5tTyFFV7YIrPiDyjzKN01
DcgDRz5J2yrR7e8kjpzh7EGV379wOfFUOLqI5Qq8S6jzR272zk+L+kqMD72Vye81
8FSyUfyD4bprIpKaRNIzbxYaTEPo7SF9I70reWG40ovUIW8+QkzcauMWkh0fywyL
udwFqO8SY1Kv6qT9afoeOU0tclhZcE7oUx9ng3ZYL/S23DiVS/GvZVHKlzEaDZIM
l8ikT9JxxFkGNw0kf83Wj6lp2ceLk0430TMz4CDvFjmVp4YTC8Q7tdOmV4c+d7oV
qTRWhjDEk8VPvTvHVJXrM4+4d+hDYQaL3i+FYvPaveTZyVIaFnP2/jZHFQ/E1Zhg
ujmyvKhxkyjww6feigTm+HFYaNsyZDNgnzbGTrr89x1irhOmrHJpam44jjV/GgEl
FNcHKTMhuZQWcdKKbR3RLo9Q2/zge1wXFSrN3G7GssSUMM9qdTG9Me1q/OgvcjOz
t4d6G2BPBPeQcGTFJEvqtYl+8vbhbdZt8qrQXDDZYZstby3JPAbHDtdMZUmrJyvo
qWWyp40+STKJEGe+CGVOG6UfW8o9x9laAZhR2kAJ+4av0C0+OD7jKQ4t45AAzdkH
EtpQ55C/bwYlsYySY09Dpw9GdBsDahHHKIxCqKl3RVbKj9hByynEmKXDpt0zTMRb
3zyLEGYn7J2K454H7dkY+gxcV24ANhCNb5kDfVoxxOGv7QsMZto0pbWDjUezVyDz
sUj8ro13M2Ur1pTL6gxmxAfd2wHZIivgRO6wogwiBpAtSkBvvX0Lo5A2vdZso3t6
TbohJSM39PtWibLrXOf91etLgzIbA4FlqZE1K1Ff7gh2Bu3ofXTQLNtTcGS1xiHV
MJX4ZSLsR89isygLD2kwXHotQbuWfViqPPoXQPgcxlYOxIq2dtVVwSXK9AoLkrL5
N9mKlZj9B0Ag20xb3CEPEJ+TvQ5acbkf4biLh+n2H9K7QO/k1i8D1eq0EcEhQmdu
wlSeLC01btEETo+igDZZtoMnGRXJuWmmML2fnM9D1ie7w1Q5gtrIFb2E1BfU7xWD
2C9mC1HbapIGZKoxzMDlT4vpkmgJ1uBqKsKuANh/Irq2EEoVvNvD73U/2d2Okav5
Fr2rN7Qoj3ca4Cm4DMPWJrCjrZhM/eOh4Z7TSlubY9nVasQKRgzmJisEopLfWgeG
43HmXsRAizvNv+6HH6LMmHJimG7qBuFxPRptSVN67f6M6MhCY6eCMbJ4Ym/mHCyy
QziIQFO1uVQmEHIRCv+CU3zgcDJfnWF6RauhNBxNIiDd6g8oySHaaNDCh5RRAisG
0Yfm1Tz992HgGZO+AKNWiT/4CIoDZz1+VsKnBv0EXvQaUTHiFwvSW1S+ztkr+l8s
hkLqmrVKBVw7vUtDpONktIj6WqJd9iR4CCMmmJfLwPzaomSVTOYTYjBV40KdICa6
yVmWPm2lBSBT46B9EgkflEnLY4JAFQFU5zkEALIABpRzxYV0NSicbrtwFJ/xjCct
8pKyZt0c0L85Sq1qgUa8FGsgtwQZ+63Ej66QCwXGuZ3Mh5vaA8APKrZHfXOre7Vp
bgzpymRSGOXo9HKf9Vei8UuvEOLMCHSgxiixnrKt4CX+Yc7YgnKyR84JLrfWqwI3
va26O6RqrHl2SiwcME4Pjmmu35bVCtiX18dcLWGQTutnH2DIH1Kges/BqocSyHHO
vxDVq94HSRdLsef6JEm9ADD576bzCGyZDLbSJn//PkDEhhoesd33+dt1zcKBJtuE
ufrq+PUYmSyZX2h+PhHZVQ48aTIm8AvTRO8bSe9h9N92DshSdfkaufdTnAqU4iVl
aMBWkajM2lLdzNsLDF1pBwuocGdtEAlS+OA0MZRkZsexEHzI/7NsVdpLgz+G4Yvp
jvuf29j/dMK1OMz+5QHU1d4tjSylqV5Wj/Qhm+EC0gRSA6RhXfR+tUECc+3l9EFS
APGqHp21zT8pcc1/Ra6pLRrFX20leRC6HCW26JCnoq56j1kxrYtFtD3G/9dkFYcY
Gn7pFsDY04DvqqF4NWWZ9raXRpCWlw0BmEetg1MAOlg4oH8+VJfFfdgjkvyi3E9n
oSNtlNNpDJ8ezCxqSzNvCDlinKsSMjjXT5qh9SQo77DACvOiRilv0OwFDjySaQKe
9TuqzkivFkPEzEeL7ZOxSGYcvKbcWvpnCk/9XIMDT/dl78iOtUTkslW1Cn1J3cFL
/Topl1omBPVjseI3Jt24woH7iAzyGz1UVvx3FU96g0wYozo//BSL4/yvfjd5UD8u
g/7yd9l0ILQg+b/6m8oSng7xNTPUqyqF9r5AQ+Y4MLurlllM1mtCVf1QvB9SLAYu
/ndfiYzDKy4nN2bP5/l8u73KzfTE9tI/e4DDyO1Vuc6LfZeLmt5A/a7HQXy3sLm7
sTq4V/clhrG2OAVH2MKLnZh5E5O3+jyKd4QqzpprnjrBO//KABIjY1S/HrHpvENX
8A7jfA7fOqmBUpLSR4kLYT8v8Y5x+xrxzV8z6c18mVn4bO433UZ9mhU9AoGb5KGK
rt85CyukOiFs9R/Ok8ycyeK+Y5B9sZ6zjhKEO/XwIECDfis8Nnx9eKnbTvxovFnK
cEJjyr0d+tbTsHrc/WOQEzEX9BqB1yuEH+Gzy6PobNAcgtz/x6EsKM616Ijz/Ibc
9rmVu3naO+2fdvWAhMw0Qb3hdOvxRPGps/S3DA/seTl05bhf3cOmb/ZAIeX2D9Ub
ZsDDAj+NWtER2wnn6wGmCJc8Fd2O8SlTCGBDGK2DpQPfxYafhCDcA8EcG/mN6Qpu
nWtjUJ+u/4BPBDQ/HT0dv8HVvjRIXPGmoU5DKkM9uto+WoEyk8RBzrvtX1BG9M6G
9PRjN63BAZ9+47OTt849QlqJgqIargYCqZmDkSxsK1xrqKkIK418pBFK0DkJAt51
38536wLxQJG6MxaAcHuEqdEPPOceV5IcCRYyxkWlgExfwU3i3I3aqiFK1ivKd/Rf
Zy+aJp91UtoFb3G20Q5uVM+87EaUFhOTenHgipTt4n2pTvwkFUt/awvebHUM4Vhq
rJUd7d3gz0RN5t6/boJfd2DMmWCcLMwrxxvB/EJ7GBAR4nE88WuOn7jesyx3Azzm
bY6Ew4NCCT8+jzsdXpuWfDVeXh0rgMqRPJbU7tO4QLGuR3gikseGwFOH+h9qVzg0
AXWackw958ocKZU1FmuUn5V2Dh+KDW1/UlFjuRnnq708CXONIPcjOlKZXMOaWklj
7vLl04GAbal5k5NGX9ziLDa+/Ud4bE7ZVRRXfB8KpP8gXpHRQWGON+tGG8qZnK+N
Bzp/+Zuos1dclE/08aFD8sZaN23a0N3Dj8Ap29fNhYVgmdBEF4JKIti2LINoigPq
fIRyk0RG5D8xZWoSmbm+2rs7Kmt0L6sL6JKcfo5HHnNrDpY92ItX6zMKBqCXJ9Ph
6aKGJpt9CIWORYm1LaiBLFLPnuA725X7C2SXntb0D0gq885orIbS9bqXdiDgoOlz
TW5HeSKUy6x5DeUyy+R4DnOwQqG0v6BIGytMqsp2EnB1y41obIXAafIhxSH7vzos
Rweh5XRU0Jm6+T0ccTf4nVJMHcgDM64ctjnWtoRhYSQoDOGlfr0HkeUUtvYCi8Xn
8dq50z9hAbFs+HnxAX3yLWSAw8pSbhW7hIFmBbPrS4YgELbHorVQGGkZfW0RdQRP
d6ajc2RmMpn8uKsp7+XqQgbaHR9jyOfU/8tpw6za7gySsfrxxmQxexYwg5DWR16A
0Wio8xzXqS2SoPxiMbXtnW4Xz3e6ytzofhMvRO7snw5aYFFMvTFOs6E66rQ+9w/b
GXHXAjGMZbFXvBtN/FRtYpBK6B3HdBkcQj0n5JXLDwTi1LBIAjcdrs5TC3QsPCE6
KFo4S2huCu7HC33xq9EZemOa4nMx8PgN/PoxuWH37M1zK4/WZZnQhUcIV9X0SxY+
3/xYPaHDjJCq5+A3lVb25GefLBcnkgUp2LBkCQE/gR1xXKxdZiG319aJ/QzEcjK7
5ExC2S9MfEyvRY3bYx7FrP2HzvqdF1GNdIhAphKECc90dmpLFOLdlw/8RhE3S9IR
nkGTq/aBNjAVu1smKxiNsxNaMcmPeSmU045V1j4vLuXnfUHcPzu59r3xhIL72uoh
4OroCrGBn7tWpkd6WYpOFLUdtt7woFyl9jpRZTSmmKbV0e0FKKApc/0yDNofsS/y
S/dRDvDCze9C/8Bb1BcItbczxKuKowF5agjs+mxzqSICi+d50nITn7LGisnPrqX8
zyS1/zmAuHhCESZOA3qqz6azjkQAE1smc48e8ATtaHMfjApNyY+sx6fkqUc49XdB
B7mOAR5j+PUsGF9Ow3cBURfWDbDpkelwoYE6FlsyR2SqDSOdofI+LKb6+eSNwjfk
MERA4YFdze6PaKIcKzuqeopeg9vtjplWq7mLIJEI3+4JtUtrzCn0kcE/9b3LQE0T
m531HaFWIhozJYpSJQLGKBN2azc2BFJCJX27MibEhtaXjDe1tdaefXJxL5yROnTn
lGOAZhQ72Br/2hQStm58p/3EaftsX2sft3Qd5RmG5LY2RwfF8BH4zzK1BE9EsN19
iNKVp2SGilXkWQwZqOHVwywTzCZEt/BNACnGOwfgEmJUaIduY6YgIdVbVI0N06D/
6oPRYxia5Iq6nRq6nUyh0g0OgCohO4HIYOPV3iBzdol4ys94FTGKy95XSGKnEKO7
pokF4BGeruS8bPzpnqv9H/IrR8JGF781ozxEbKRD6S47mq6GzimPTUwFh3NyhD1V
Is5iYD0/y8JHRswwPoY1Cu7mRO+gIPwkRF2/tRU+wPVqIaIk6r44PWcbpqKTkEfP
O96FiI4h7I8tSoal/cua/DLunsXhEMT77vcLzSvNrETCGlhg0EO0RyWOmcD5GVvj
IPQat00xn6FiGlBiNtSacBbnH7hD5oE4EoTuBqKCWK7WV+ve2dcwc0u45o34Ndaa
zYZxLY/zGYnvHBzPpJCHHOJuem1HS7DDhkXMwlWLPK9K5yumviofsPbFIAX8T1qO
S9VWn01sW2qGAUxGixIHS1e/oup9nLxoMXA9CUx2hiZFwefjYAJ5Z6dpxZHu1YDf
cF63D5ICosICyM+GBu1KabNNWbB8AoDj0nUiSvDVbMbcG+0qYz8MmTX3DwcewVe0
cz3nkfHXNkOkzzX6+z5/sazYUhmQB84U8F9TUctT3zRfeJtncK7WKcEOXRChLxLx
Erma26Dufbp8xRr/pPIHJIKOByXhrBiCZpjsP603Jv3d1PUVfgas80w0h1nNUWNC
3OzYjeaOkzqfaiyXPIZftkHhUlZ32m+egnpVEov6Ej0zk2mDkayYRjqoxbTjYOic
UQqYy/hAVDej7Chv3LO9b4HU+zcTgHYA6OUTn991z5ImDDywUmArRCaeI/uW0M2X
EwiY7ye2ePoEhH8Ah5Mr0HIfnyLWW9cKUdHDzsAmiarcM4H0aLKTiJsWUG2FEeEs
mnjXCT/U99GLEaxsq1SNBEXYsoBNcqz/Szso8cxfSN159XrODlfcpqT2RyYug7PM
Hxft7H7l9otM0PeN56ww+0d5ykaaf0VwtSh0m3EBdWaF0f90Hrpi4SZY6rzKJVuX
mlYM0SMt/5UX15sejb+/dXSslrGZBB3zhG1Z2sICumlEsIfHtzZxESevx6CjQhlq
rNK0UBgC0pjCPmfswF7yABISeF0GYKulfAEK6qj/6QgM0uOzl47215ExnAvZksG0
5pY0nzpP30+nh0tBxPRfoq6PIISDT0R63dvn7PYBY7HyqcIuTKF7wG73XP0SrS/o
1nmGn2/lIwgvBO76Dmda1Vk5L3OYoPfFf8qeAs8ISkZqMvZIoilySy7ArNS4mu7b
zNHoWjEjPrdk3hMlG7ha1r6RRr91n82dt1rl1lPtJ9yHGc/nBsqOiDeKQw9ToYxi
j/M9UcOc0shOMThz3hpFgjKsyp9g5Ea/0WTNqfrb0AQl9ATbioQv41ng6yb3qRWZ
nmSrsEXBduL8/mHAG2DVGMXJelIBgac/ugvHl1V+k8QBt0wNHO+zZIXKMUY9NBGh
5Fy+2ZrLaz50lP73QDmoxWBLruwhqPfDfEuWrF05glXLliaNjeJmmP2pPgfE+tpn
5gHHZaW0oG68hk46T1xea+a0dmeJjzjJDaUEYOM0ajebRAWZ8LKiHA8MNhWKvne7
qHnk6v4iPacHSYyclxdOM4F+nupPP/0HLrwrQS2F+tOFxSFOBlXl+pfi5QJr4tnq
W7C0EFT2tmN9+lncswOvhk3mzhrmABpswupIP54bSTs6DkDtQIxE6+rtMXXs1qTJ
Ff977kzy40V2W7/D2vH30tLeFJDBIMN8uSLERuS7GbLJPrbx4FXTny+TvrbEBjWD
u18B62l1MfGRiemUCTEwP0OThaUmJvAJD4yf0F2Ky+FTlL2VYeTETmRWikAyEfNx
18erMN9izWk5RMhjQvujYgva7DwgIg3hpTOFaBgvO48gHO2wlO7XfOQneQIMaskO
/bJBq+yRwbdTz7lwgoHNGQGmN12PPOoN1ClXyIIYHo7vOxnoQBgjSM9035pYjhyW
kA9l5td5+/OICX1HlsxUQJ7PNhufdv5krAE3iaqJvd9I4XHgY780qtoT/PIdwG3M
ZQzFlc9FyJFMy4c7l36S8Uq7IBj1TXp7cujyJ1xRB53dbgbxJWatBhxlA6km94cI
gbHrObutYH167l01z0qFJSuKghsYLTKx7R+YjHxZ8YtpYM/jtWcFiWw8CwIPsO+l
S3tEIR2G03wFc17rLPYWIsPDQuZoXfS9VnP0WemNjpYy/A4VrLuPltpHcuTYCdw1
oF0PW/4pXykIZEVUJ8ldlnjRi+iR/oUHh2fB7TW/SLyKATkc5D5yUgOhnaQKq406
avDGmwv/cDm+K0UiAa7/nk1BF9KG8F2nhzLujjUz7MI0qJ7/4vCBBZeMaq7HhXXF
RchH4P0klM2XiJYwpVu4RjgzTKLuvkZKXR+zXXkaWwnBNQ6cORtKyIK/l+N3uLhH
hYxAiuy6omtWDJ2UHy6EWbCHfuVvV+KvEO+8MBahrlUPs0LW/JKGvWMBGkH3beaC
3hGByZb6ov5Nz++oPWbg4RdxiK9JgYkgzjY2YUtSOU5LxM/Ywp7Z14/8b5gga7VR
kIjhUJ+UyJbC8+xRzBQwl8ooeyHbCMbkmvNLF4RzSZpsJpEbZq1CZsp/sVP3BDKm
kXOOzojMQgwh3CCEdO9t+xf+Bil7rpLQ/aAMOSL+hdtoudKvHmyPYLjz0hz+//6W
ZdrM9eFO2z7XBxye1AX26waTgUp5WX7JncgHcwKwcmudIfXtoi3M9kvKPAadATlT
oX4zS/LQMBMvms+BrzAm6Sp8KbUrLOB04B2nAmwObIq8247pM5tsKxLd/GlkYuNe
qHw0WTLksS3YMH6bTzKQSQEG1zP0ulRivZpdB348P4UbwKMIgAvbu9px/E43Km98
rpl99+gUmSl3x2fEJAWDXhLonijU0cJk3+yKnxIQDSXm7kamrqIF+7x6bHhMTRhS
a0G+DXTB1BWDSYYGkTvjaFb350ZtJw4dTdLUWZbKBwfQd4+4JsXDBqiRbvYzvOjn
K8LeGVnXO9o9Vr9er8fgFEph5oalj460QY4QCN7ivv0bB9A4l2HFW19Kp/fZlNuZ
IpZgytuG0jyMi4PRlSPopbIauFVwVOjm/7SPFosLWEeYCW8XscveOOqUvmeJkniY
2svEqR0/8TVEQK8UBLQaREAVLjRVUBm5j6OMkT5+spOrxFLdOsaLTppAjtcLrtY7
Kc6qe3MxL7bvP6QK0i2nAajVHDR8EEbCvQ5/pLtVlK+Fmu6PZMES48HG7JCCgM8N
1atZWMHKRR+Yml/DM3Ih3m+vvyjZTj3+aKur8uIdjtl/eNuMmh/PYzHoo2ttE3wT
wLlbhh4I53rKE3/7Y+3HspPabzS5ED2gfU3c77EznZ1NG5F+hwIJte62AsrL2jfB
PeJdnTrYV6+OJGJ6HKMA02beJ1Pg9O17i/2RWw0G3jQaAwtkgM/+h81Gyl94mqqn
dwHhBsDT6VK1q5yj0HS/CU9uyM2nJwOGrbwcU6W6WgI/l/QSfZyZkLLmrz4SaOf9
dUgcSggTiq9rnrx3eobLSZO6XR2NxsHbFN1O0B7q4DjNbHdw9PVcCEEPAuviDJML
AH+QGelKtKLpTGl5L/80mW4LklTnedXpss8XI220S2adGoOK3r7qtiIJPzVlyiop
jpEo3xWv914C85DXtxVODTv1Et6/2kOzprX4VwdIu45/xbPVfZe0Tq0jTUdPAVFV
jK4L2fu2VpkZ3ssobpMB0oF1G3OLrCFFm6THLEPjHNcU01VR/+W8LPTGvuEBr6pF
hY9yG/3biXbV4cu6RJFY6nhPZkIo3sPWgxKGDvhJGGTQFqJWcgPTiWuWPUIfgCAE
hG5JDH0xP2gMS+1PrclAkkEQ2tLVFIEmFHJZsqv+gWHdz/R992VZOo9/qCxMHfbr
PB8UIziwzELPVP0Wl7YWsTlTWxWRTTVhBpUInOKQULwEH1j0KnGCiuUs0goLj6Kz
2Bv1wMVBAXAvFtMEOLc1nlwH0+CLVIGVBmCbNSl9zU4U8YMdbGJqLLGcRD77BGza
kgVZf3EfLR3hE2zzxOrtkvn1slG5qeOTMORXxfTPvPIyiUGYSVeQbo29wBmJYo/C
l7ARqeU9QnBiLODgaCKffB+Qwpm6hpoQ/qbo1nuzol0XKmZ2IHr2vzg6xDtYllfe
4q77FdlXIbQyw8c3MizNpnCu6wxHwV0bLMNdchjdS/NYUL470ladl4N3M0hwUAGg
ZiqFjNaFdupGIEEJ7U9HAKhUBI/APCQMJ7nsUioS+9PsUEtR+XKmmqYv9ADCkQk9
g2mVc+Oo7Bw6y8OFgYSh2mKZRlZWBqKDZQyCY34N27K7shzIzLPIVSZotN1Lji64
09EQ2h8/IYddAhpH6NgbZhlXCQH0gwPFdLWNZSF5PNB9RIPVk49VbR6pAV+lxk2a
ZaTFHmBur0m3tyuiQ/lbeiUcPTACxmSkzzhzVAhV2B0FmZWEj3rj9aU8XbPdg/+i
lcmU+PeGSJrAlTbwrDp4ErU3f487E7RSCNtgsLhZIe0KCZS0a91LUiATW5Oz6Zc7
55gMMg/WTyhBUS/z8No0Znh6+bV3Nb9Ntki2pw/duxqWbTooKWNFDq+W87jmBkfh
3ix0NWhQq8iPKK6RoukPlrJvPjC1p79ebSNum5e1DNVjeT4peE0Ll6Y9eGJYgVq7
oQdZkQB0RMreiBIgiwesKO63O6sJNzsVmlFO6gvufljpss6FiNMR++CprK/pJalj
qjrlar3xP66Hz9dE/O6bso8Lh4QxXue3RvdOjYvJazNEm/mGhALp85jMoZMInLkW
8c7a0n7tRf4e8d4e2RoFJmT1Q1nFkvv13ttYbL3J8+ff7oL5aE55jdI3UKZiq6CE
yQ4PWSttDhxlL/Wd1EAvqMEWMPB/mNbbSKtSFGtb9An/MDF59C1XQfV4XAP+ajkI
VHNJ2NXIIfS23XImJtojz0KomNfY8X99U8LOQTQbNEmXLia03DwZ3/hKEdfWEo+3
sRI4Jj0dpvoGShVVcdz9O/o9sYXbTzq86Zt1ULnzdtJ/p+7JBGrBKJ0SjFqydWsM
YK3s/4hDYHXfzqDx/DOBb7BfV3Oe43L6W6eYR8nP7eB+sQCH/lrHnDqqAn0U+xkd
0bXeim5V3oGgBJ85nKWZOK5z8ZzNmz2sSLwTRsx81uqlO5GJUbkX4Sb83dbTq4Wd
26AnxWMBYsvBv4RiAlpMgwmFTRYHzgsUf+cqQWRe/JcO+vEWJBc2cmrzQjRMT0sp
Xb9aX96lBRAXnW1D8e0fA9zkheUlh6U4zIffja81ysVcUi5ygCb4NaYc3/w59LQj
nQ6DKITPNbU34WiNh8CwxEQ+lfw9vepOHD4Asg8Z2P1rJsvqfAJ8Kf+7gbrwcbau
YxAO4b9DMhcfhKNkGt8pHSipVdzgH1sRoqSUKhCENBodHuA57Uljv7wi83zOVPcZ
NYg/4RZccuvC/sNnwnD98+mg08qVg7yYk38lgn0RsCdrGsab5Nz9wt22W6vVjVEk
HJwK8RxoAQ2K5FNjDzHiWUYG30QHiJyaLj/3Hb8ze8iQ8F1nNIOUE0365wkV6r4p
pcpFtXGSQhTp5Kmk1qtkYeXJcEgUDBaAhxj6qHtSPjZ+XXvn2eiS5kxvuCg+fCC2
fQZKyfpwDopEMgB8Oh4t1BupwfR6vw1whOd8L6X7HmbUWJd0tcHGNwd4PQ5CLeWT
MNUbFEePJ/gtZ7Fnl28cBPNPNeiILX5/Ifhf4dfpOASVMClTNBbFwmjfwxwudjc9
YgxX0Vkxm8kvgvfYfpKYqKVmZuVRYr3P2BHZnJQRYYtgvzIwMcbES9TxkrfwYP+5
MiFioSU4t7rx+LgduPtrlUDbfguyZ4vd/ZaTj+jGzP1r5wIwiN88ftDQP+aW04F5
rVAEcUVsJYEeJCZ4ZDn57ABsJ0tAG8xBFP27gJBSXubb0tmWYkrylksuIITtIKSl
R2L5puLZ1ftNT8RKGwVL604U7EpDRrzCu8Lwpuyig2/XgRLh0GlXimucfuEVjQRO
WZwleA8uquNkNcJQw4jjMu455QyJnybnJwpz44CIIM7YNAJ4B6uDklXfLa7w/ThO
wKdNIemDaaqou25ro4C5K2HdG+GkasVZK96yVcCesO8Pht4fSRNY/SxT02RnKxkP
bps2HS7rFQ2K7TknXOIMNK0GpKnPtRFLX2iJ/NYZ2v+h2Z409InJCKYAJejuPAHU
/oQZQHaYe6R6f57ATmaOcDKFkJzMwhcv5l5BUK/A/iJlbtcDgQVZ7qt3lsk4oJPs
ocjNI5u046fpTIPvHuDE/G+/DRfgqz9G1vMlHkMQtR6cgJj78tdeSDzVW4BejHaa
TLNgPw53lvnZWNaZxYzzEplNa07/LI8dcVFfLAzcGPwVYCFZuMEqvZyEI8y1yqjL
yTdJJlDJp6TMku8MjQCu43Y3hombf0Ia/GGbzwozZMUIv6Yb/eDFc2t9oRe+Chuw
u8jZ62NrODbayIvZa9FD+0qhOxs7Yi5/ZJq/zgNApmooBLHHhrHlLcHWTtoaED1E
6Pvd+z78NxA3XnKfeKmCxhS0v7E50qepo3MLnQcSSL/Iv5zBHNz8Fjykq3R7MoBg
bbZ3vPbWLM5pZWaWLQF4PEwLLisB9vZ7R+czYts4UyLvhmg8qvrKZPpdZYJqjdlz
HzuYvB4udIGXeMTA1EqB/XJ3UzNqd3uEZvf9caiNZibaiSKz2iNRYVAUI8NEXCTz
Q71OBiGKX/qBeSBIjO8/51OD2AOld/8Ndo9Kw1eAvQImez+wAquJHEinV+f2EsoA
6ujE+NUDoUA61CVZ8jcflu1SVYzzf8dMJI6f5M7U/8stza5Ckkt1CWE6lOMX0sNT
eZMvlDRAkmadVznEBgHszh+LQUddJuPC9OkKb0VIbB0q4Hmu45kVsdfBjp5kSP9o
eAfLp9FcQijYPlCss2grB6q4KGKMDxgMs5VKXqlKtSSX7skLPaW8cR8cRuONSWAp
mM312IhbARgCA75wUbbGFmru3ZAeGYvognL/pSbsVUAjaVb2IT/Bg+bzPLMCJ/x9
9HzWGHBzjsXBoHrrIShD4TtzrRBlhWxVgUWc7xDRRJVzJ64ALBVRfHVlCo0RiEwD
aw5JLLDRNXOGNQ2tT9f3mOfWKLrNPVGECJ4PkVUVyKEaLw2y/7N8h2BWHjhCcvr2
wnHggYn6qtpI0jsvHlMPdDgZDHnkBoFUnSXt3+rMtRudDshFQaEOZcWwZLx7b7rj
O7NLX2lBE7c/qQ68TGqzolP97XjQ89CkM94UEDBTattwEZvJs4ZVYdkNVuUU5Rei
IkEHpMygCBlNWS37Tb4h82NwRVL6zdgAeJOFtU41dSxKyEXOuworb6Rmpma8ER8z
dTsNTYsDjSE/TxVSfqFC4wGvR4b4LS4EOQ2huvlYvRLDXdmuigNGgrrVLfDJRmWA
jNUKUeWs82xyxiqD4CP6Verqc208WYNUE6q2LPbEOrOSI1ZAF3QcG481eN6Gs9OZ
F/Jfsk8Si6covJtP41r3/nv2K5kpY0OLhI3lgUHsScVlOR5qtodwwtVr7C4q5rAz
G8qhTp5ngfaGA4PLrbN/ZCb+Zk71dsm2/JNdKOS4Hr6U5PS698+t/ggxk54Ip5PC
etopVMg7TWYMHQL6OVl485sLt2i5y4ZfT2PA6/L9IvQEZ4e5H4ntJveSJjzukcug
DYt5KbFbgZvnlRwKYk2DItuDIRBby/sfExhy8rArMaxk92GDG+/j5/61ZPDDOesh
97UiQmJFfgEYwuXE3LVRgV16nMn2p82jU6Be3Mg/X6uZoU475hWmW/Xrl4IlTlWS
JWjaCr2Zwn8uxJskElvyd4t7JFShIQxXRDm4ya8xTawWaJC4uBDFjT0OdJWhzWyI
6bvvX5nqEAxqAGsmuhUjTJOzRGj7dHnNCUU/vKhEfa70G+lPeL1itZMsKt05QpiP
TcuWZ/enPOoLpTB2McRIS63hma9IFUfT6hDXF5esDfbqOAdBotzllSGCcuEPoufh
OWg/ee+JaIHmK3j68p+AoqyQbunp1t60vUN+uDFLty6JWCXyCv2SYAH5tGSqK2E2
5C3iYS+51sAz5GRUn++e8HGmTZUEstMknvxVwbMZUtGeR/HdbPY6aCKgqwTdRpNn
/Sctj9vaZJKBMaVVViFmY50EKIrAUpeLB8/arvSIQu+IbmPDuMcWVxjdoRlhbBNN
BwUd9qHkHZwwjEDf5+r1JXhrC203V/Yea7n17xkUY17DlB+cRi/ULrxjWo0LjEON
dNLQDR5LV+kN8tum7knjjx1aI5KUjpbvMhcivxpIhxorN7fNx/a5OwSqZ1zEmWHe
pBymzCidv95qvSiutk+MaBSdN3pFadO/ut+qTikEkt06/yTY3d1r3oOoArTJqaSk
FmSsDiLi/NwmihwSOmZw9WkF4Okh6EwhmXx2KaWaMeT+A7Q3LP9Y4vv8lcAmY6aZ
eaDd199LBXAW7m2b7DpPv/On4NrOEMyy9MrlRuj1YxijC/W62LtXdwxwMZVPfuLU
gPRWjCgxv3/Fzm9J2yPcOS9Qc4txhyXuZ8U1QXTr9pifZxkO/yh1hhozhFzEutHE
X6mRXs4KgJSPYDERTyOuv3Gli8Q2SfizXxSoHq+utCMlgipKKDGEmCuKryvCv0dS
FJ26oSmC0pedo8/s/74GJYHsoDlZ836x2LCnuh0bhzmacy1hh2v48SACFnu1LZws
OUo5w6qlBTEUwwaIcXn3zzKKH+KvyH3Zj9SQga0LHuqiDSNAZH/fFGVJwBMbWUEd
mW0CVoYgkVboJrzcLHjZguEtCABtodE6GXyPjq5dTKuv8QGiMLF+1/vxjdjE9ZSu
y83rM+nizIcIVKq34oFuKZ9s/aFpkNvSKZ87tae5CB7/wIgfNOT8Re0F+lemOBDm
N0IMZolhR51pfyoygt4R78y0p8B5N5bFWT9X9lZUfbPREAEW0NT44HPmjBXagqEG
f8PWI04K3vZJEofTxruJUXLWIM2QyxCwBkXStvRihp2n7FTFlXZvqj+11JHnHrUn
bDIydfugqTyf2tZZ6rB0ZyLP02Wl6OdboPmpYyIjkSrlgJx0xwk0HYYkdIRZnvpx
aD6xEsEhLOwEFd8IkBmsGfHS2cIgeM9n/Q4ePY5C1hQGjM4OzVT1I+zk7B8t8PIv
316c/xwR/vRKH454uO6Z9j09l8V0IHof+5heqnfuNdJZ+U2lAnhtXwRYVN5fLt0i
xrbTNlCJrhifCc7Ms+STsM765HaAUP6JBHZjQWuIXFnRRtvGvujRAzwpfTsVBISL
AzifZGPLQVTEAQWp5Nrz266oUo2H1YnveT+kDqv9iqTC9x/Z6Vcm/cgHjZb4O00L
3b//5PcxFWmf/f/5b597Qsp/4DdtQTyeJNjVyjrI464oo8tVOewwxUdjLEvtjA4v
DKtTMQAq8U5VFoaIsl0u+N4jrHvi82ktOZEELs4FHJjhayxQDu2MiKGu5PXFKEe2
0js1uRlweTBz8skWL7XsvS9m85yFEzFQ1o9Y1AL0sX9Ra0FegRPhkh2wb10Ws0Ga
6FTI/wI53pPhKpvnnMWyHf53v2HFNE49SDdfgP2BIH7dyBKhXBRD2jGZVMEhU7X7
vXMli/htAt499I/LmjLvIBS040jkooJDJd7YiQwAYv3tIA6CK/PtBpW8YtNldjpP
J7ppKVZFm9jhO3fJKpHylFo3vzNQWfAtszsrNBo4VaanEkUgMAmMC+01/94zHIFo
veuXw76ZxSttuAHB3cj3bm/tc9+WP/ji9Wpmeo+ssSL8yI0XMmb5X24+kjwOSya6
NSFTITfl2WY8S+k7lA5KPRVeG/OYTOEpDFd2TmeE3tfjkuuauCXezC863fzcI9WT
an3bumuPl/0uqBelOup/8dd80wj/y7i8FA80SyqUO5ze07kF44ROTKbtW73i1aUA
G8tahQnYg2Oo26gKpczMQ6ydELn0lk67cMbUuBuGhLfzH+jrFHOeYCbMBUZF0Hqw
ZWEbDAMgswxcSlEBXLLkg8z9pIxowhUcc5BW0tF5GYolGQdfEZY/ip6wfUsC1hsx
f2XiFMaVj1J6L3AxE3DMY1FQH6yTW8dHziYHq3FNIc6tbiI00iYg4wyDNhJiimxs
gExHm11jKnkuM378zIDa2cNGXiGk6dozeEpJYHbCAf61e3kNXiigXRd5a/Yh1Mcg
n/7oSyoD18hPyq9l3zlSyKfCDZ9OEcibk4OB7IS4lOh48/m/X4jhYRUgSRQ1e4SN
yH9acz4zOVM1LBRnMWhuaQ3GOUOLYfm24MbEYZ+eqCrlt/o4mx3yd7cusJIaha0A
wocXPrx+zYfmzFEfCYbYW7zwVbg8W0R9qDx77xmEFYnu+OgUWWbQmFwol7RmlRc0
3H7sAwdd1nOrFYCpLpBx9l7/lXzH83KT1LKmuevB3nU6sphSXvEPejS7UmNod8WD
FVKqJ6oIGa0o+zfuJ2OdnLkrZu3QpFurfOKp84wIkpk0fjmOvlZCH8OzaeUaaHQl
skiKaZ9L6URdccGP3Xe4/43/Cd2tsYYOmdRMCTG9prr2EydTn/42ms7EzYvsUPfp
gJ+3tsY5upwKBgjflQggnOYamaNc89C5lGzzthJXr329VKsNBF9UoaxOhAAoQJ8J
3XxwRxatCc/oKXftIkUh/gS6aCSIi8MCQQ0B4jWINPC0wZrBEX+suL8k7W4md4Qx
SMxvJ4KZDopoDX26O3+X+hbAEWh2LSOljdFq5TzNdWQ1xZlMrIP98pHMKQToVpKo
FwRwi37QpOZ2oF/n887uJ/RQNtyK0xi9PJ98UonfqzkKOIHjDIqct+BLKUf95mhc
gempJz0OjBBLGOdK+CNal+urWk73v6PHSLTGyk0EHH5zNv1ReWbmmi+ReLcURVYZ
fDuaJR7eRvcZu/jixB3Stk7RlI8YdBYAO21/r3895MM/SzlQZyWEOKs9Xku95BNr
Mv7Bo44UkrVVHesducw8Ee8uKMAdT+9rKWxyMxw+iXky8Jp2kwRLOaUVVO37gbLD
nG68KcEwhfxjs6E7x2ZbpQ8CwGCk9bLman8pjKXlyKwQXOACcxNBPFgbW8QWumEc
7u9HkcpiTCazaf/J39jow4+hDyfsJSr4IProIopSo7Kh7AaIoEzlChdO3Qmm7qVo
5hOcU4NryXoegS8i6kojT4OdommliikbWkxtDmaga78JjDyxRyrii88OFuRRaCAw
+/DNpmxyhoOswE6q8f+UYOd7h3+CtkRnGEKLp3q1dZYl+gv6dSFM6mkVuPKLiGHG
R+zkSD0tjFK7zHuJeNcsqdRyfsQxrbC/jkLEOar+U1/hLPQoK6vjoOn8jdI0iZGA
DylSWBFQ9G9xsCvm70NyErxnbLa1NXMdd24bdSULIrXjiNv1g93h5xxxEJxqLuGk
Nobv0NVre8yYsL8qJXJ6Ow14T5wdbT9NsTvFtfswEWXZJFC/bUkDb+M4MC1pkXr7
ROoo2pc9Da9NxFUIpvjoPbXuuKys4u6NjC3Pl20oVM/VyAOceSXl/hmS3pM82he8
sg4fjbKMC9kpTLEqdWAM9cHT0qDeEJpsELl8juvCbwKrEgfaCT0HFAmK7hX2SA06
A8iN+bqp8EfpIqvJQgRgj9KIzWZ5GuEysojPEB0ji9H6OGWBZrOk+fls3ddD6BCr
J9BRYUJPNUNMzTX9b75BhoxOPNlrZ8cUBBUyGATRRksmS1xxdLA0EMbr7+JrZnI5
TFW7rwAjfFSzORuB6W4dyDv6C10lt+/os5haCmB2BkrAYP5IJdvQc0jliMrY23sB
zmX7QT//dCmhJxDRLA4hSNw4TBaOCLjTB6yzttML0Fl04O5cIe7N8my//OBHrVto
jrNwO6bKvgRHqgZe/FgINbY/uJxRo8ws7JARhEBTo/V9fHShjxAQRnE3eh/krHRu
aF08uIzOYbUapu9kGKJIRfwtF4TcVAuukqMdds/2+TpaohhQSgOrnl9yZm9Wfk5K
5vPUXm1BaaHe/AJidWzYLKAavFn6sTFlpwW8ufwdBXpJgEwGF8sbTWGBKaJBnzhH
uz4DE8hPnqwEkte8FEYn06gR78J1KHetDNdaTqoDyA2g/dNY2UUPFONXXajMNAP6
IVKC48uO3s45Je9LxeDnCAhVIx1nBOeFIUk/8bnhsskIPB1oCsYcD/3p67/FM9yn
uZbfqe4mHTlXGBd3kB1YdJNHy3uUpJCTTol3VBoM/0w6fCERNhUy2itkwf+67D3b
5IzS/3QNuhVm80gK/SrNq9k0IqBupuUocryJTYtf/BkUAB6TXvA6/wvUPyAIOqhR
UHkILL/0m0jzT2ltUJ0HdIkZ9ZwbztoZ3HzJC4ZBfa5uvtiYFgknFGYoGs0ZHnBZ
5H7qeZufzVkyIeUENGa/iI6Tj6urBcWlKenUV2hhAO9Ue+zz9ZGKcgvVrCDu0JMP
c4liTi3xsjh1xQeDjEdMdj1cZ00vfujBn6/jIYgKm0cko1mt4XcUpJTFmycrc1aZ
BIVAFhAeAqk2UwPSe5+qlEPsNZp+8bOvtkqk4JHA9jabjX+tBKk86Zt7A2RxWp+i
rzDvaPWbsZdAFcsdb88IOisbbhtXDFICB3XrDTRrk/Gnq/kauh01lsnl72pipdUA
gv6blGKw/+kRwspVzV36E8J6bwttM6gX+ceOj/atyblXONKV3EeEYXryCCBZ5GDa
1zJS9WejnkAM+AkOvXL7tlVGL6X0MjyXouNX4fv0xrkKvX/3ZfegZ/TVNqPxPBDq
1WNt41xedVy+6zgJKDd8CZ80EIFo8tVKjE/o/a97ZglkXjrcN8S/1ks9pYVk8zUQ
s8dXys2OZ8f3dxiWPGEF0P6iBs/jmsX871XJTxRyDBqJ+YIFr7n2nhDRMEehYGbj
Fi+2tlkj+om+Up58ch15n1hCgextHIvBxaU3aYriTYrcPZGhitiUuphd9qpkcSJY
TAmMFu6L7ZOEITrjrZkvSwovmebM79OSWdVzLCJ8kD82jtNua3nalbMJyLWEiArK
Qqd+HWWquqwTNDZKIC7/I/7K+iSENY60mXIb84P9wRxzB/SVxBOTnjza1fRJdkqv
r3LqZugtJZPwgRCgRB9NSq+pl/MOU8PPBGfEBSc/cINWZ7UWpc5dWS2XmYZmYeBJ
W+huacLH0hjS2ws0Nuy28ajhA/eEwZB283dMdvNM7lXqkqWqb6/hJmd2+tB46oq9
aZK6UxFCMgUKv0rcQ8+eSGJvyUx3c+fb3hZG9OoClobFvij2zPkB96Uz2yF6lznZ
2WG0qaTZp22urVq+EtBCIkQqF/81tQerZzbULZM3ABu4O1HlM6cuNcJIAINqNojg
CPBdbJodCzd21Q2lTUyy10QNYXwo0HPdqIeyCSxtbMVzNKghim/oGLcs0P4DEEOs
MaIVr1GFm4sLklBqqu2ItSmtchkJQI8dSMxZEyPYCblW4yOz7SKSpgQP6QR07oLf
d7QU///PhW9MhX4hE6X+2X0zn4TosGkdMQMgqtwsFFc9mYYGo3niBsq2TTKhAwX3
8ZLae2ZuwmWNiLz9ufvxo7jZVXjVqVb1UVNk8ZNkOdwjqPErBhL0QxF1xPbCRAAU
GScmQQd1AXs31hxDq6nCU02l6nldhe3eaWeA3S1MvnQ0fFFFAg8SmKP6rFpPVd+C
6H8lHjUSCJujUDF5E4RzmOs3VAR33hknHLjrlJ29QeFKxzl8C4b0NxCYLHmKUhbO
Rf5vtE2v+GY7CVPtgtNja1ZJ5SoRV89ANGpgY4dk6eKb/pi4+JXMLel0XDNGOftm
CA7bfVUy/99eNL0ACiWrGHy4/6ZLLGj3DtpPL91MCQoB3Yb2DW2BbooeprEjgzaa
vV7In2HIViByCoXOUkRi2V8U12Ce49Jg/vFLaKHeZ17vnEPYvgXAI/TSEcHF22nw
baxEaCnCTGf6QXbWzcR8jxw1dP9kGCX0acUqS1VPlI7v3HWTgcJ/J/ldTdH5PAQu
E2TjZefl244UbEmhSctKlMmSshY765jcZphvUAKyVI44SiSmDG9cuOL2qLDhBlO1
zAbZnNvySGvaRpZ75pctVpoij3yN+KTtDsFbzLzXrFaldhQKyWBScHhK5ldoqWSL
mIg7WNvfAIOH2gTzc5GBEB9/SjwIOLHLV1pfovCztOBn4OjtOT06lQhXOGfuaOFy
QWiDa/4cm+GWj+bUOQcEqqDzX4fE7NewXtDZoYat50htrr8biXbSb3qa/XQJGqUW
4viBu9R0qQ0haTTRTPd5ZGhIe1vj/mJOgqP6vfm3HC7Fm6VVt6PBW0j/3v4UdTnK
atVmRj4F3FjRoKiTQVg7mEyK5FJ2hw7fatHb4ntOIni5BPom6PEb+W8Gv1zX5dlR
W3bjJ9ptupDbqj0uL0SkQNV8eSYwcMOZQvgdBRW9ZRBjx7H9TDnM9KDg2w6JJc1f
WUe2Y2WYP21dGjSF7WSn42UvaN0VNOUxJYZtvglk+lh/Ip8P5DLbiVxxTKVrIKnv
mg/oTb1kGFiU/nn+LUdXxl9pjw44O8N/Y6j53wvL/8a+uoigrdaAy1D2fFjBYma9
cPP5kKzZX3vR+9wHd5eLBSpUK06e0SieMFoTTXTHlIOqUh6Sh0Xq5eQSkBFly5CJ
QDf99EMSPKeIWGHJ+J9qWSOe1iZ7gmVGYoYyZ5tqll9XD83y2sFdXElL7CFdT7bg
/anL4+yHc1h4RGlcCS657xyXkllRRRFu1vZQKYNbagxr4WhuOKEAK+zUUwW+IXkm
MhsMoCk6R225bIa1AreZ+AVQl304FDWj0yFQZhQGyXbsTcb6xqxVpaZ8AvB70cyn
qBc8NhhajWN70YwxePHGUFgePm5vxCQZpQ3JdxMChQ8yKSxwponLBBxA71BmGPqb
qorx9PpBBAhN1o+TEO0qimc6rei9/yBYmo09Eun4TU2u3YYfwVycmLmOJooDs/KB
yHidfvwPfDwh0mqHnQ3aFNfPEUPXDXBqhduyJTOZFA066UYqt7RFMtWO4MyIvAsX
8R8qQLp9J37b2bxEsvgBwXNzbpZ3kEoilnrkzorpW4XzUySTyF6re1cC9UgABIsi
BgTAZPYhPvKmR19gBfMLJtSEuwNfX9QnTyAQJ64fJHgsGh/i79Bb7AFx8l3vZro5
nMEqlGxNAW9y6UVbazNztIPZP7BS8JX9LWdvkQm1oPp9OmJ8nyLeUaTse/oYbFWE
sF3pBQlPBDjgJc8KSTA+V797M8CQ/AQRskXlC46zeQRgNMm2ZtsQbBh5Z2XCswqW
rojpdyhRXNLplStq24MS34RnYw1WUs+PswgG4XSczOStgfm/+n/TmrXlw/mKykjh
0FHqUbSTJmRmdojkLpNHhHLDFksI7RCI+9qYmHH2GA69t8739JuquezrEBkj1jeg
eVfZS4l89InLLA9Od2tGuv0R/nn1xdnoGz2PVOkNEGEWPvgxan7aZRdnrJTXcY96
y140FWazt0IeyguzpxlaUWkD7y6XjG6oWb1S+5x/tjjI9Pb6PXE0NQFqOuOiAlg9
oTrjCSoc4NTEV51rkzDrHSS/GB83ARN+QoiYHbUNmlYfEvQObCiTKrnSXUoTx8rd
i+1L/TMEw9r7Np7/saskM1EFYO/UlmcjPzd5yQTnDvGFC95P0Mv2oHIjfkY1oXb+
jRN86cCO+tzPOcn7Fe0X9E9zavtuQID1/ew6PoDwLWn8lp3WRwqvZZvibscMHlOQ
eyrymXYd+fOxKbxOIciMfsf++yWxobX5NBLw80tj7GTS9jIVaUqg5Ey5DbkymyKU
4Zr49tGcCezxflobZd6yP2qjjrZ2dk0XRMo3/5R05QZqjV2eCRvzYtrHCX6iWSwQ
xKz+0B1S5+ytS/PgEv/bL/YoHDmK0A1qh9sdHBaYRgjW3h70fQB7zaWP3WNIWqCz
VKZVlR2LkuDDE0vqj0zzEXN+taALsw+TWnHdWSiz9eDYfjVuqFe58ZHes+nPRP5n
AhOrCEqKgytjf0a3uoJf3tFkLxFvwBJwTJOA0IF3ga6kCmtz7PY0RQ2EOUA1Skl5
ykgeC0s+AfApIy3gC45Iym8w6mpdbHgBHdMMk9j0ftdj/ejm7MmEub36jFUr3x/g
prjK+giKAvW7vrYs8AgVPi96vmj9iOIyQFGOz5IqGaIq2IYMcytzX6ig+TjgoUch
9vS3uX42CRCiFPraKwtM9WJvc3PoFsVFOP/1NlN2/yin+fUlj+t/6YdxK6nI3PGm
6uPc7P9+Q1HfJfOduqIligkK9vLG+CliCfuyoRNiEWCTZ4MzMVrALAh/Y7e4U/gr
ma6kMRZtv7fmkQWAmPR6L+1eX4EcsNV9yQoz0Azp+PpdlMvD178GywrgGtU/Oe1x
UBOaCP9oJP353S9O25sctA6xh2MIyMc+KUn9B8W5ZJMIWMUl4ikiUKw5cFkGIx+U
JJI4OUjM8a8OQ38WKq7L5kToaQh6lTeHbnLMfMyTbFQzrOj2NSntljNI23HRXudD
w6x3bxn3kas548mbMJr8NCbJ/RoVuL/sQySV2oFuKDmZZzEFh/rpvtkICHRyfso0
Wt6ZZy4Hy0vYqJrLmB1CY3PSwkgsNv6XMJrvcn7PCpYTC9jKDzVYC1FVrUyn5iFV
BHjQXavc9jKIrMhQb6vh22qlJ9sswPFaLOHRoP3UWe3l8U3SaXVVXmMqG6s8pEka
rGKdgdAzQL/FFPCmiq5NFMd8pn5f4BnMI4xtcVuc8tROoKrYDLL4r7qVqUu7aYhp
SJhm16PeR6NVIc0wX7vu9AKyV6vn0El9I29XinRF9/o4fbAHHeSnLMktGfy6bBu4
XRmPCJRIkttYjZ5SHFg2pscbuT9NPo1rjWNIuXSWnv2bD3YcGJjJ/oPQzWBHczve
7MEVX5U1utCYgO8kmMiNlPG+lvYUjiXTmVtfsf5NcZsNoXfJIWa/bMeUb+f0rrJu
bK9J3MlkOwZ7FK0bJNAco9khF6rHyHsZq/DmZuz3nhy1J4+nNe6CuMAIXW8bnc4l
90T0P9Eh/FQ25A0wF/N5ZSAbMcEDCfqp0uUMje3CVeT2ZqZ710TaCbLkRm5PBfQt
CfyKc8zR0vImhxMOF2cN4fL3Attq4OJSqf/DHOjedKgDnqN3O/a07Gjj26K/QUSN
IpcCeFoMQQjwoeajWtPsThRBHNFbeC2+4TO3RrNoVVD3VSlY552Nmxw7MAp1SnrY
2q9sKERBuVN/WvBdYD3IS3SGbv+DioKNs+xfR01Kk/ZrKX2Y9Hzr1XOBZtIKXojO
vcTWtLpLvA6RBl6M7hUljAmRiXPlfNVP7ZFjm4zsDmR8XDyImDcyrFkraWqIySZd
tX85Y/WK04Hc7rtoZM5d5Vxeuor7fm/8jJGBh0mqomOVui4zoh02xK4cZ81cClRG
0f2mOAS9ncYorZO5XCBhEDEjWfkK8SRAg+AiG8UeLw5VdO6Z981+IwEq9vLURnoJ
/GZMZej0ULureKAQI9hHD7iJ49RyMbUsCACxupgXjMGbAgzxaDfMyoYRmfuFv0IC
Q4AytgGjQBJamvPPoMjBzDyRenYHbFaofP67gDavIUu1Q4LEDgaNC5vhMEIZNtR5
IovpVJeLZzBI9+d6ap9IGmF46qDzpyb6RBTiow5bEeJUs8nE3fClWugdrfih8raG
jcVAf9bqmq3qD+1QSF+B3TJKA7jxSz4GdY6l6IfrJF9V7Lj8y8kX1VSiQx1Bby3v
+icH6ZKR0aEnswBEGCowg+bxb8CoYGnaDDjqwvAv4Kk3174rA+pCrUOGgkzd83Jc
NS0cZG2tdKmhYaEgS9Q0KxWzFjjsYLpNYZg3K+qbAlqR/z2V+7xqLusSBbh1C8kN
L9ARa4wvd/TBuFGA8jxj/onvKk21x3/wb4pudhOEUer2DOF6GopIxAWwxqg7GFJH
blWdH4R6pB2MdAVQYwAT1v3F0C0XihED33sTOHA9Eh9nNFztik6DFFUisp4jwsFq
ZXvu+MRpc8tyzKVzpVvsLqstijIIACDHUfVDgTL6SX0MHg2u5r3UcmgltNtuwqhQ
1mhSKN5FR33zR96levfJuC29/9LMI21grq2qFxiSOtF6rw6LA/ejff1zVE7ygb7R
EXkFyoWqE/A9OEbbZpg+TvpfItx7G2FzlNRI7YxLy3L67duJ7qbQhoQZd+PO7+2W
E1SN5ycUxjX5777jY97mPrS3QaKTKm6jmKJl4XC6EQI0NozVnnRxmK2e4XnFeBfO
apMWCFHPKW4uE5azaXnKkglbPjgrXv7gQ/EnLxUNU/5ySHIYwJhkE+3Za70bm2wf
S1KJtZ1hNOhBE60gBgp4xQrrACPUVU6HZ3vApIYi11thySdDOePqTMWsFdrJoF8I
u0gCEtY27XTp88ox1/56hPtXGowcxpd9ARAujldCKiCUlQkHgDVOQxQqRWS4vDKW
vQTc9po9HjMdtwVv8KLNC84J3j4nIaIGFy4uBKag8XNia0urTMjw8mfmFiHX6354
yMqZQ9GmHyNiOCOwp/ESBVUzvfX59k91sD6I8dn9e+W0NFA6UFs1ccxDY+Cc9vaM
qyOxAC6mmKdCtvvQc05qKVH8G8fWSOEFUIcaXOdw6xzrHsmwXpuXhD4EQ4hubrWh
vByfzOyheLFAR2g7yx2m+B8Irm9w9UsxySsrcggUre1khma86pOXpUJA144BHrRN
v26gznnYiYjtArO+2RdKqs2FuaUVr2vpor+yqeWvZ0rJy360rle4KswTKSff1yvv
oV41n0s/514nHHJ++l8pcYXd28PZMT8GUWTgMqbTUMyCsCruX990PUvfDXCm1cdA
Az7mjq8kYKpHKF3vb9s8Ir7e/a6aJPvJRwputDrwPD1HAm8TXap8gJL0KHjw5xp8
Ezp/7b1xG6vmyMv2VZCEbAy4eFWtvwqhYCjpl5lMCZDuosfouoWSH42Gw4h2pi6s
5gSyW6GPOVeTgITgtyGNvEED9VJ+AXzZYp7uXQFrCusLSjFH41X5dRt0EMmfoQKm
/PlM0BbM+6Cl4SuQvH/CshNge5TKlfZ2BZHzhxj9+TCnnjVOypu6NJvHN1CGdCfF
gYuXLmuQTU4mpAMK+A6hdOQCFnPrGOvj6GqF/321sUMKerqUMbVJ9SJNKUDST2tv
kfliO1X8xJg0t07EJz0VGPyPPjnJ9jxpuidbtfsxDONyqo6T8whqvMK/GFqEfqvv
hTm4qtqxvg7ZbvezvO+2ivC1MiT3OTPKE2LxXIptTPGNxE8/pTYeOm4DlAlvNVk5
Yd/uR3/NjkyAqHT827nXzdlA0hWAg/z4EcDXOaI6Yw9ZkN5B+1M3tbAQn8DMkjo4
B3Q1xV+OH5GVJ6IYd6nluQfupj3h0VJVHqT3tsCj4ooxmtIbLOuZ2srb0VzgAOqF
uVv+2L53jOCfYw20KctTCINdEDDSfgAo9iOvtzgeWnP6uasjklYyU8h+ETi7r0mR
gZU5Rhg7L9m8arjryRqdmawzOqNWEKp9Svi1c8BDBMEn+jykzpZ6HLxrHpjV7XpR
owl5IK3L7MPizlLKcUZGZ/9Zla6Vn1KoLyfUcLc7WXW8MEgUFVKrDJrdKJPaO8kd
jhPTQflna5JibIpGMDiJu8+aME9KTOpLd+H4klJmfLoMgOeqL62dzTCO+bPor/ug
6SfQqzsWlsUdx8xgKeWhQwakVWT0XXToq1/dc+CfsMZx9z6PTox7moB4WS9s/nj5
4YKq0VEtufddPX1T6Ol5FZO4e/5Ekaayf0FWSH+qopgkI4Wg+2IDR9YLrqQXeTin
CyvY4EsslpMPKMtPJ4rZnSlDFyBP0jSzKxoJNj6L/9y/yeOnhf3BQeWvET0KT0l0
HpZAbXyxA7yw51GvCg0hWOGRTPJyQeDrhQ7sEuyEpbEW5O8a72etfbboqqKCxiva
elgfmnrW4Qih4KJ+oQOztC81+pAJvS6ajKCxGf5ErRgF7tDFuU+c3FNopT9humLP
FzsyhgTmEVMjEMLdIrOh/rAd82BcWs+I/UwS1WfZTxaUc8+feWqRJ/uSVOEIIRNS
L3bbmPy7tg61+KYWlssmxuhrgx5jeyQxHeWxU1OhWAqFsnIqfc+6ytw72HNKXD3M
5ru0ep+v0CUd3uQRqOmT0kn1Fmt3PgTzE8WGLN9EuZpAW4v0utPI1L4147iTWMni
IT7HnQ5KI+sdvk3to64wJ4zA4w9GNf7oSpUePOdLTiPoMmLYp0G6ap7siBZCFZwU
a1mUR8ucLmBWtMxIUZ2oLGjmC9kYsu5weJRpM8POkp+QR/x3NmEOttE7zh26+uUE
RIeCGS2RJpLZ7pjS4qZfOl8S3u3TqQSTjnXVhBLDtw4U5UJuQhFtt3w4OmqFSsBd
fvQUd7wFG5aMGyUEwFrWXJ2bZ7AXV5FhFcX9p+WYobvPIdLX6rpC7dH5MTAJnFUU
n9U7XPZHXO0VaL2ODP6ut5AxGGpcKUWEwDpAx0r5Q9XfuYb6KumWCguS/ZmRKMe5
AqJtpV0Q1qo8x4AePqjUmJwvCWjWgj3u4MCFvEbb6K0iad7nS0UJk3fpeSkxhacE
EmTV9YwZBTwQx5dZaTF449FGaw0OBhUnGzNLg4hS7fZgID5UQFveGW/YyIzdrAOs
C+yrFo/JuXxX5oYNrcpHITxHU50fWdSVIbiM3uJfuuqtMfT21NBsqB96+G9NPZgK
sP/Ax2G1BfNgZj62dSKvAzXNNBle4h0A5EiK4JMWK0yEahXu8VacFpt2H5JwMQs2
KsoU8tc0N6FIF5GHPbgG9URwF75zTn+N1AsQr5MJ2rSQq1N6A/w009q1bdTV0KR1
+zBMGqSIpWC3wLpI2R0pubEJqioCb3v1xujyHelyvIz6EH/kCHbmH68Y2YNF5tUh
6/TUeTFKQvM4Za0AKYx9z2ZZpHIE4LfmFyA5ANWePd78i/zS0umIGK/YPsYSv/Xe
8OjvcQH1vM/2rqf3IDrBBEHcdQSINpZIgxCjBjjywNWLBscmlMhmyv4E/qZrN8j6
GuIsOYaWhalRDeT/fSjVk9JybGpGKABn8DHTbtF2yFG48GjUmQ08v6tABKmspIiM
8tD0j8RpDmDD2N0fuj+LzCQ83NP6jKqQvjNB1DFwima9JCwAZNnZV++dU5DMLDnI
DLXJVtuA/jKbLdII2jGIePOkTkEXb7+mLKF42w0x1xQtWpJnX8GJ94t3BEvkaeOg
KLENXl7ZSboO8nhDbG9akU5ayKw0NInrUclQ2IglI3YwGptTJTuqZ9OrpN91IRiK
SnI/boqpXNgV1ykiwlZJgRkQ5R5Q7qcYLSzTTEaJs6feRWSMMf4i784sqxUvtAGZ
TUpRx/aIDiaLISgir5S5ldxX0OWxlhHEx7ABJXS+sLiq1oByEYi+tUpDnapeBBSY
aPxNLr3Eegn5CJXiawdVjKdDNxnvxDV4jwZqOM+Za8A9eDc673TK8lrQkP04yJcF
ICaqlyRgF5h/XqMp6+CKgevUydirpgRNljXLtS8MMaboUvrEuW31XbNYH6/MeFs4
9lRQ3FNUA9R6xvja7GGXj7fWEjxDk+FQ8WzKkqHLyH68mTTm8gqpMOxmlHpjEcUu
eU0b/DecX8JtohYj7txxa586ayvjFMHaqK6mZ0R10K35AAA3G5JNsp1z+9KRsBk5
+PG54/IkzUv2OF9Kq/Zylw3YfosisNFUR3ec6L5l+Cl10OAVYV/5/BWl5nAY1W5C
VcxKViGNihDDEVbNb9KBfq7NOwLHkYocBOMu3YuY7N5XN7lSx+vaHOXQ0t6UPtqQ
wBwHlE44ds4+GfIM0HPHZKZgFjqdwgzz9jHAjKDn1fG95UChyuWAUKg3dYDOyaiz
8XE1kchsgSaX+RNckv9Fj3N4QAFCl0a8B96PspKCFpUrn5H0zRmEomEuoBG4ky3P
4vvGuG5YhCAD5i+gc2zRze8hnoiSLcoCbXfmPlLDxKu9t47KeukTzD7DenDHDGBG
hjRRkdBhsTYVKE03vUd9w3OpyoxTqCZSNRB9N+wgOjKjmv5WUqNxx78PgZBprqM1
cWJIL8pMf1V4qFjPfEyHNwF++fitM2H86eSL8daYN8aJoJl9IMcnZ+Wz9zhGwpii
lofJdKYSiodBH841TaXzVh2g0DapzG7l7Zos78cSB40T9aW97rX4+M0+7GJzoiNx
F+56t/Da7PzuaoK/pVs8xIRD2BZNNi//4gKBiwwwPZ3bGOu7dIfNJxKejQg5Oi+M
iUFGtWehBERoeU95b5yCMfLUgWjqklYM23TavLvBE7xyDnRNYepeL2HNVdxwzBdd
Rv/t++/aBdX7uHrtxpLDYcTmrxNncJ2CoWOulY1MeFqBHccKVc98O0ZmbYUOcF0k
ijKJ1XXce71ygToutWw7rnw34cM19US7DvvDmdlG1EPxT1olO5c9ZejMpaICdxsP
pUEL3mJbWwMkt5K3zd+H4B9KWhXspwjRjnXxgUushgDhpQ87W1PEDnDv2bHT1evv
SviM+AQn2WJyCcX+sYAI438VyXjPccjpmuA8lKsPrY5xJXxRBXYAjrlY0pDrNKS9
cTSd9tFlux9LdUZ8+AzBDLMZtENQwsu/7oo+Piw/2ARN+P+55GcwECbWPO37qpUm
hUHFAspXwBXdA51vwN8RaHKBqzIkClEXAor60022AMra/aPDFI9wwIC3yZ2Uf+/C
fsYVPk4Uvz2GSOVw+3QCnWUPezKtrVr6KNFIUjCaQqWOWip4t0B8TDeIBbPOPsZ8
SgYEwhVZJ6Ez+9cGEt4JHW3GfQ6RfmXhOueDAw6bviIGMdAX1OBiclvfDrQoZZl4
7l7wDv4RoGh2WYTGs/+vK00AgwoJKUyffLccb40LDTsyMwRtBoOLAb/DYWlZbX5I
CVdYqeQh/YlxVLTbiT4sR7bWJ3URPUpnpkQZF/Qp9LiB2T/QMMVGyXZtXo1RWbFl
K1ocqO3GN6l3WDRO3tsiXOeWJ0ufPg1JOrRmSzMPEL5JcdZq9IR88K+Aew80Qpti
q6XitxmnGektz6HJl3bkyJadNKvGDkFXNp6zxMlXYkTApmP/AeTbvgHeUIVY/yCN
1c3PtmHNw8lHA5YWL9lHeHmo8amruazt8b0HrQg1cGRXhJveH2JOHVt0oCmVVio0
upf9b/8IJJ2Q1+Qhmj0IFCR8S+m1eX8hlSNF96X4TZU3d9lBnFXF7eCYNUNVHAF1
vcM7OqVy+D/ynTl4BiM4+xXsmqvgIllQwg10d5K1Tq0FnfKhQCkeALNzSdCeWguS
sHbQac1YFoaYbnNs6COor2J0a9bTw1wMutNXKTTA3vdatoP7r8kBnUUJ8i6V2Dze
NbJveBqAQN5Z2qMJ3pGEswLuLSI8L2RzmhbRAZu2GzYHdB5nozxS4hKpTlouhnBi
zsJ3jGZPAouXmVkmmq76zNQdfNPSMSk737RMSyhbCVwtgq26xqjpfCQoiNw/Z7yv
CID55vUO3dcEcxIua4UZDl9Dgg5d3qA8oLdp+qno/5W5PRgDbaeNZuBIbouEW/eU
kof92qFHFcWXGpKiv8TocJAGgBLPPPE8elcRSnE3YP91A14i+576F0by0WHukpzl
jIqjFMmrJZQew9vBm8jyqW+MEcYzA+znqYEboXpOuMU0XtUF+CTQdWRVOaDdELE+
4CvCK/FLNNL3nUvNmwFquiqja9ULulMUrpABAcA8aU6jG2eCrhpnfPd4oEcUPuO6
9Ko9W1Fp8fNskD2tHCF1hobe+UnThxeWKm0xqN/ilDgh9gX3Q57K3fmeMAgQwiNA
K07lp5+guqiUl+NUFaUiHG5upiOCIS94zEichye3SGQkkvkoKg3OGQyqZtBrG2OU
6/dupUIdy6nZh76qwXO+bvKzx8wILFAkqZPe+qwlyTP07O6n9X4468lpF18TDCWj
glErCXn5/CWHRhx+Wfl/DrKTDlu/ZW+HxuQYh7H+sWyH1bpq2FDJKaUgqryfapQq
bRoh+lfkeBCTKNlEGcSXw4b53dJ0XHjj1m3eEDfz6cExefLule9nqHWiujE/+JMP
p+H4AJCN13+4lMOqH/Sk1Wuaoo0SoMO5bfqprwnXfDTwjtsRx8uyaUvbmhHpBv+i
rOxGHiCv3iQErvLqS9Pnb0Fhu+lt9HkrVj4ZBy1TVsi9S31kpOCNpzA79rxHTr+L
eZWa6k1TP/cPeagPtupsIrn+iHJwJ473PUM67wocpRIXsRUqXchtSHqXSa+mu/rw
eCxEhEOnWxDH9e0qcGfct1+TdlJNwFeMXEEdFJcR9JAvDbDiusDlEzMUts0QzJqb
ayPfxqzwsI9WP7d+LGbIrONooqJtzAxDSfEonkliD2YPBC+7ZmeB90uW6M//Li/9
G59bvB+m5uNgbIzjuukGs4YaNLtroYexkYDOd+F7Z8DUgD9KvYu7zx8vBmxpJA3V
5yqZlj3F0EFmzM5uQPIQ0jSCAbisHyP2qgVwVz3px+lNyhwfQHpi3f/knQSwJf0J
450sUHB4sH4kgmsTJ+yCPxHjSwoycpAItUSht9iMT9eKaDIuf/CO7liT0Z532TyT
nWNUPA1+0227D2+FE5bfL84RSE1CwXybc0+jcxsoz5JRKYwlIy5gYPnwyOteskfp
YCbKx6b2Hv4HrFQkSZnfPCRKdHMlP+3aPJNnj1SRNWOSTk9nZiRImE76MQISsTkg
Gwv7Zy3PXM+AMnKA0cPddfvHyG0K2Hgqk+VSHWZe9kL+cmarBmuKygtxlGx2ondN
uyewtgl05rTOfqcsCrUw+cNAyNCUHICo5iKVcCATp9Vicnrem8Y6N+Yqcw/uFeTa
1JCmi74Clf5hmc8DTfCy/vYbs6VYT/A+c6ba9g1VKQ3+o9XQ3+UIl6RBRat6E27k
ZfJmmlAMVu6kwSKSS8e2zf4ioCs26lVa+x9JIm5EdMSCbQSyyS+RJhFJu9v+N+XC
FeooaMVgzHIkFHzE399F0XSSk4yE+/jDTSHsi4GfmBjBfYFTfSH4u8hDZPqDei1h
dYztpXn+07p01cSqjVMcnCP8q23IZiZCJVWA5KwvBuka5owfwnLnbeK5tMjbDEi4
NxRQtXlacOYikh6cA6Abs/h/5haWts4GM1GU9PnO2PyVb76EFQ4L178PtQuHUVLt
wiR1LKMZxMQtyaDgZ0gIntrBwbpVFelOVRclDtDblbK+tIok8mrgYdobzKtijXQi
atJTr7YtWwyF0/fbPSRelNnaXvaeR+ggK/STWNA7JSM2qLFcHEuelQPSx91+PLPz
usdR1CYUNV4blUH9yCuXefWA0M79q9XB38Vxfm0bvSasFjXaGPd00qbD90TCedDM
mYNUQTPHLx62qf36sqt206eMdxwyidTWry8QGfv/cZAw3ZeR8tKnrc1+ZSxw1YyE
4Y3T77g0EoCVj9gGxdg1dHSMQArBENHMLk8E/9L9n8dv5t98jD/zM5TSb5XSRCZu
xg7DeonJFoftTE0HMMMZ9V5nxMnXOHT7Pg6yP417n71Yj0QOm9agi5YBkCK270bl
T4dwlUmf0VqS6hUYElUvdu6+48LzWEIVoy2/exealUUSpE/wUJ/dzc72MymGSaeL
z4J73+j9elcsJnMS9Zs6aNSmyuWo50EQ8n2GteqN6tuuuZYlKyXlbkEGlCLre3oV
nsl4bWhPaiaeCWL6K/9nGboBt3MOoOewP2d0D7VzEP7e1cvjRQLZweTzLM+D4Iwl
NwGFIQ50fJJh9sE5hcvXSTX3l+ejp/10FK9QXMhyyRuD/9zSnhkfRTezPvVZtnEC
/fA1CZnplBZZfQG4nWVKghA/YzS3CdyLJ2+6aRjqC1qLt6zIo00qpdka/jtPnQ+B
AW1JLhyvjlLCG+0lX1xH/gIVQjC28CCC4yu+vQkBKFl1AO9NZjDaDXyUdvi+iwkb
T6DxlPd1hWunEy1lmKwT4bcfJ/G4SYAq82YJqkPYzutPx2zum1XNUznJ2XaKtmN2
4bZzbQKdNfIIfYU6tufgM+ZudaSka+IlcsWqP26P/0zpozqbEYeUzCywnjQhd/9Q
aBqus8c0ipH0RIdmVU1wnfGG1d/ii/S7PpnO95mY07lfNBJEvHduYor6YXw29HRr
AOu3sPO29/oEnFWpofW4dlgJgqyycbGaJrBhaOEGv5aNY0KMCh1jwsC6KfoObmg1
YuWZXMKiQuerWQrp+cW4dn5OMJK9t+QLBcEMw6AZ4Mzj0cnUh7GXVxDkNGW2vKaK
YlDBhMMIfLGH4IAn20ioBZe9xplX5FBXAN4+9nrVSqStKfYPyF4ajwxp4m/CLypR
mZ+N3vuRA+bTK3NzQHNUGouj7RMOgL8VhJQAg0NRKHAK49twU2xI8qwGBqG0Yd8N
68guT7FXxPWVuGqnfdOeTSJyQoJFPrj9Xm6nN3MeyQY8FDpfQDOkXwuP2Rn3xFMu
eFbrqQnDMd6Xz3iIkPj8vrvFkDxZBCMIMCsmC6rSf8FMuUk2aV0FmuVUiud//iY5
cR4quYNPtuJawqYB1xUqJ9OlFIxnACUE0yM5LDH6Yw9MFxE39g9urOtNoVQHTnDc
RMM3gzmsNZhj9M7r9YQhFOzZavMAhDpDE8e3EmM8BRTH9kOch8Vx5vS0sp5+Mx6t
R+zpZ6WDmoJs8BIZO1Kn4znrL77bJJMq6f0NdmsijkFX066bSWhkCDCE+oNDl7GC
SNUGL9D7ZD1n8DX3HGpXObw8bOSvdinlPZI7mgc8ROfrOHuUvcFUMjxEN1Xwtak1
CrPlWhtIo869KgFos3NrXlLPzOno8ZjaKbyKm6GVOUOO3ChQNtRzHntctR/6yZuw
mvMr0uzFTCMdzocmN8ztRPFt/0s20ThqCAiWxkaq2GKdO3FoLiCjfIXqmljffwEJ
vtVUQzZvVAIF/q+7ivdWW20QphcWNtkdzP6FoIq913Oo31RT/egyEjIQNu9ubReP
BaJCI74CRBVP36her0umN9HR7tDjBNELBzXk/ohx4exraxMSBl/RV60cLe/qOoKp
20JBpCMiPKwD/GBRplJAXnroAD/t8TqL+QuNByPnnlHG1no7KNfOL+x05jSNgMcR
yvtiFwNKUmWIqoKlyG6GSmJQExKQ4DGw9fSxTySt/GrTs3Eb3aR2KVKkMciM9T0g
lh8ACM1yEIACVA/EFrWFJKIacmAMqjt3qCKcYBilUFSfHHFdWmDaZyZ6+boANVUw
xrUCR4f/Rbs9mSXMkhyyuTcx25a18G562dtRveTfqzuBjSheR9GeY/hDd5irafCB
p1oa6vYDLUiGAB0uNerdpotmHLbWIKC/SkN0PIBDHia28rq+XXD53U/T4iKaJDSf
4lHaThFSXMe86IS734UHiJ5jRucgY9HJhzhrX32qZwa9aT1HcDgQ0S+iFxVrAlHA
KFQJHeregTZyjTOIRY3fn1PGD0/3UbriNwu3jZlNiLmW3HQ2PhucgAo0zIeYSUDW
x3gT1AlS9phsTjzEXEa4JGd8ZOG8NwsU1lQbv4qgQVgFHAh5qwI3h3P3zBu7oKIj
F87LJ3IjyrLSENOBZczDlTRw2N67tt6ykSALVHBCA1paay9ueLgq58DOoJz7787p
yCvlIR7On3kzSLuBPRwKCx7HgWsR9Xp0+uejROiOsYk21/6HD23C89Mm3jYDH36w
zB5Pw6DyZZEJ7FrCCxApvLfrlSkUNThRkKvdsKiBqfj7dXJyM+e6hzZYhAwYgRAY
Dtc4Wr6KWwpX3prEVkOli7Ni6kdTtysDMr9HQAGT2w6FLDcCotQjrBOiLRhfeZlO
xdIM2BvlhAvpf2E7iuTlncGLeEIanWwtF6Lp1uoLlrZs+Q1Yz8cGMe/gnAP8hrsY
ztcK4yQV1k0TKxxpsg4yFIHe/a+uFS0Bq9H7fzgOCJJgQ5mZ9fvZka7Os87j6gnx
lenfz/NhHOKZY1Ic2ZJUq/HeIM4uKnssyrHKVdupjtNB96vdhA5VPf9zVLwDO9Am
00YbndZKkQX5piGMju9BsiOMtGc59AGdZHumzQJ3D3oI/JSc26k402Ideuaalriq
RAfWrjRnWibgDvA6ZkFzhun4nEpCPS3fNPSFnxkD48h4QGNGyWX3FxV1FxWytFkv
3bcNncjyXt01XNAn3RddyreUc1q4HzhR3IiYv0BXWCPQDCQqqyxfV/YdzUaEUbJD
CLVcfxE8rxp4TObkxnOhfc4OhTHd3jm6udoXkY0eXH3+5iPaGmLWDaHBOHEcf8MV
Q2JilQyLYhPwqtq+hlkeSIv8ezperjKqUF89eUZnxnj1GcoS0xLFIL4TJ/08/bUW
r1rfOMd2W4mk98FIKkMScmWSUDjJuEyd6YeVOVknGN46uYX8YLbaX8XicTNcJbmK
a+y4ntel4ka+UEz71Qy+uH/CRahZx1QD3sJDRXejA1tTefbuBTeWosMcLtZqllit
czFwy3gABUtQsTRzqunBxAEi9nUl0ELVmJuR5IIqjsp/KFmATY3EqHk9Zv0yhtoG
KAm9knFyvWAnynfRV3ukAhbjMOKRjY7gN8Wl4ItyPNPyb7ktq5bmqOj5JcjR6A3o
PDwgpOEKQepybmULJ6oJu46/S123wCGAFpwnxnph3Bzif3qctwBZtxQvcz9+RsHs
DauKJ0BCqWecUt0BE8NC2Vl7xqdwNTtxnIo59gi52Voh5mWxGA/be4BYfurmae/h
wazXaEW5A8dapXwqhAeNMSuK1g3R9A+DAt4yLQ9R8cbs+AxpjS0S5Zir/TY/kD0u
hlmmEwVaxC1C/DGOcGlGYWaL87Zi4WmjaFC887cOBDnEJIif2lfjFH0RYCLJgXib
T2VnVqxwED47NQNt/LGAKgT6BbnCzeJqqhtLGE7SosC5QwMFmekB51iZuxbtHnlI
aT6yKjKBvSKDnngLnCCYlT3+TwGyJX6SG3YLVifUma0FBlwa49QHjOpn2XIGinqI
5NTEnQk48PiTwLOzltxMDxZmnffeSGfKfG1Mx0EmwL61jJcLojfRGm2nlTs9zO8c
+hA41gdTX9Z+KYUtAYtFlZukgt+zk1T0tepASxWG11ibqNs49sjhUzT98LFjrIyd
OcQLFLRrhqYmDVGn02FApLtGO7OiWfNt3ANNlBbeGpfb79DW8Zcer7epJaXgH68f
UpXhY04HEtsaNPKpsix1APw/n1LixXbmGW3yNkPcPjyXHeYI5BDpIZ9ecOFW7OAf
8VPH8dfY9fJJ+0oY1Xc/bLa9sbHyCCFDRVUpDSGp45DssNpOItqV5DBsAqDaIAxX
9HeXOz1KMz0eKGbvWKGMpNMVVBuXMAU2kxy/PnCqH1lHkCsGkx2VF4UdCb5H/00u
7qyfFobyKfsMZLJefNzIPDovNNb/ORz0fG7EOf6scVCR9Q6VQ2x+jUvS5QJjdZ1+
9sLGfW0bglG8BQNYqgAjI1nXXY+92FMoi5F6tZ4UPu3OZQaBnVXlVZF2RNE2C6Ah
rHEjJypDAZs4WQ1z/JXxrVEc+EpWqnRkXJP3kBW4mcMIdTPBFp22lhnTk8y0KaKP
r1PjXvoRN9QNqftRtKz+TPbS6fotnIZUfJUcPqQ0zXq+Qh8G7r3cXhjw5G0So+f9
AKkKe/GnZUK+NSfiW6prjU9ymf6F1jjtymHGY5TsBJzs5cI7K/zLa8valcPIY9Fn
3A4jI94fjMCzlrI7j0SIp11wVzuWtjdePECXW9aqI0rTfvbVbosQouDyz5ZIvOOT
uqtJRjuAB1KmXfHqws/UT9QeK52wDuOCDNg24nY1h+I7maOpZsDgVw1n2Puz+4Nd
zd3XB8Gm6/0FggoHwPFJkSdiiZ5wC+xNT8YzjPiQZPH9r9KetlhuYqaCg2y1PDbu
8D+aw8j7b0TwSRbd3fO3o/cXUkTQ2HqhipeVsvVTwjbsz5t8Cpkyu4Tv16DGTb1k
EmR0utwGmBB+vG1GCj1fri3+xBoWdHc/xBJDIATac/quE25KkgNEyo7pe3Iqc/RA
+bRwellk7r57yi/1YD/ZdWqRXg+eHMTlHu9EHUVjr2sUzGsg9gLxGU9zGPD+S3u5
/ZMjeHCSvVK5FVQ1TaAXglT6gSN7JXaYey7yoJGVWHt/7fj8Bwbw4H0DXqK6Ucd2
ub2OLpyyZwWuwSOVxEHtBqCBCaZ5UIKv9jyJ2Rbgjd6cJLVLbPcF8hFtHDKFb9jW
mL3h/8hOJLujqSbJ4SgVkaktPzgrmYhn4KjtYUL7+KdxRhhbpUC5anXmm54or2t8
+u7kh4w1bP4P0UkJZnycT0Mutws1q/iztESsc1DnYcSErHV/VognAjse0+36DmJN
fqSjr6vI9E983wMcblhmX3wqjuxxEnN9TK82b19abWQ1R89y0iu5Un+IVUDseyJe
iDRba8wCowpYsw4TdS9huG5YfJD4xIl4BDXJcOe1W5gR5SDpkfy6s76fCRT/0p1z
vYkkiRFqkXmi5i0Hk+1sxkW+h3fdu/HNwHZWmtvZ8x8SsMnCNPSq1DNqm3pJoDY1
F57eE2tfNaqIo98KcDdhYJQTs1hlLoIznuwi7tf3h6CTkizFBoLId4OZ8ohsGWtJ
DQftn355wULPL8GoF7NnqPfQAHUgDmkcqRmbUsqxu2zLz1vcBjXe7gOBVOTlKPgX
mnVyMcYLekQBCuh6xncSCIc4VDllMP4pwoxCihfADyYKRFwhn0EGHD816f3LlwdI
8PF5qbjjetN2ywXAuKAPy0XZjRfQOFra8xcXvKI3Htt0TzKpTmp1Daupo04OeFO5
CUW/xGcHBjTpogZtFcgUDKid6aBLuFxsAyAFnFJbSkieXcGpj/tCzCkaseP8ySSq
vr7iDTTSuDl6KnmUVUCOwjVk9WdPzPTymvI9QByhGIqoswBtjhSO+7SMSrxFkQZY
qvZK/vkDv/ut6VlW370t9WbluJmWM3senYXs5f8VUDeW7eXQnHSXeJ7h3h7QU/jX
++AF+PQteO2Tp8vM6KUCzs7ZNoKfEVG2VgUfaL5/1HsAon43toBrLljGISy7wRnn
1y0RnmPmz8k4ZKbUc1LNA/MmJv+85ozCyvvS9xjGIk+R24LEeRvHmQBgkkSZpzFN
qs8yQgE9vJpKbdEe64YpeLDjQYuSB7tY9jYtuUKIaXP/0JttYbXjUKqAtORMpkf3
5imHcPhVLWoeURc78o+oOODymTqGqus21pWWPaX+f7K0iuwoV30bs7GnoG38q5px
CozVqePuLQVlMy3UYr54WpCE+inTDEru1Jz8bVBSaeqwY7kmbuIPeP4j8uHvizOX
UOMCdaeqHQZ/TRePylPUddSFoR264fNqfvIx8QawKqyPC7AlJsYUbJgUGIhZVw9A
ThsL6Q1XfS8jMzWkEOd+KO0qK7JSH//iWpuUgg9+AKXIhyG113lOilRsANdPk46v
i3pXN7w+eXCuJGgW48Mrt/BWezLXrRQEDInKz3pxOpDOP3T+Hj4XL6tiVA3cDljB
hmcgRZ24ZmjhGRU9DZI9qbcZ+D+SnCrzt5maP0Z934YkIJWnz6Dy1DWI08yFhroc
2GMYZX/1RIDIFcsX+tf7V/22a7eAOME4IUUR1WrjsnfpXxGYwvetkl3A2ePQTbUc
c5EMNuNTTssdj4Sqom80a/QluCER+zhWUUNdoAfDE3Gjfr8NNBo06gULlaRzq9+r
UqN1N4lpTaDx2XLhPCOeNW3wnpBTEJK1SbCf4keKGQO56/1ggQBv0n4EmJBd0mLj
mOGu491kJdglGwqzBr6N3frLgDbksrvZ+0H3ji88Q/eOb4moSbhuClngNxQ+zPtU
rQCEIMWzXS3Xcs/5ATwZ0Wx/dw537TcwmvLbIJr0M8HnsenRMu2KhCosmig3Wdt+
cxuaPDpoq4fu/Am9MbTlVk9O0e7zB3aHGUaXiwF2qnQBON/ZzTla3GXuqXsqDhd7
L7t4dNp8ccUaPAyD0UEj0lGbehiO2KdrjkZZhzeLOdgwgiLEvtfOH+KCvnADd22D
VvbdmOxwzn2rSuimX4azm2cqlMKMX4nuPXHzPQ0BEgAwij21I5n6VTSphuu8mM+o
5I5DwNcUeY65ZJJxGmqL49LOIPW7dmAcSo+NikRk030V1cq9ba8D73XNetpcf7zl
NFUd49J0E2Mj7BdH9Tp1WeoDh9I9oZvHMZBiAzcrgWgQIzKRJZ18db7QsV6SBzxE
U7reLZwA3SB8AnMlJdrwGafRD1pmWly/7OzYl5ngjtI1WDeNahC3BZmXRCR787rO
aHdpmj+JqH5G4hkYmxDVw6DQlz/QgjI9/AwGVqp+DCmjFlQ0bBYTF29neQ/pydtJ
W+C64I2ii0Uxw6fFGHwG+hcO9ZaTCqcHdrQdW2WoyINZ84oUjkXc5fdvJNO/t00e
8+hEDo4u8ezsVFw7rIq1rdHr+MPpjGH/WInirF2/v1VJ/Fan0zuzXXemvOO8moV5
e7wffvZFAsVXYGw44gMN5QLA7ps/JG6wwWN67ub9VzWA5D4+OhtCZeV9wiNGjXHn
MR4OYFA0fpDrqsNLKKwPPd/rRWarqMg3bVNZgpsKR2b0vSj0YTbpGFYAy0PEch/d
ia0X4SPK7TyMtlXbx609XKmHhQD2Up+voXVb02rVh7NgV8a918LQgSrTnrRESYgk
vySsd2Rx9GKhbMpRo+5ayd+0Qee1C9e0FxY9TYYxtotWP9IdW8QZuHSxhhGFSv2a
HepjqH09PaMdT8wqKg1S2QGw8dAbFe97lTJHiMOjsC+ZIB/TqoOys7NKvb9GC5YH
tz4J61JAMDhszpuVJuGuBVDN16JdBBNDc96NKF0dhBYYu+fcODInHvfAXlIi6EaV
KkEyO8fvgUsNCwPb/l6IBtQqL6uSOBnZDjgQs5S2NPQTiBQ+1AYhIf788r0Tw5BG
tW5tgRCf/paUjhEoxrvjqtF4vMZRDPif9B2xLGWcqqj6cdF9i82uaNVdhvEFs5UH
fZdy7SRoeh67U6MyM34wFJq4CUG1+cypMRiXwsnCF3yVPkMwatgWgSKusYxQKYmK
M/wqPo0DFyZrusCw5bzXJH/3Gzz8GEODgE7wvxYa9+5USXkmo5Qlj5cz8SCNv2sx
4KY7tlm41dUqSz7Rzh6hAZ75ewUSHCVbRoxPUlaQ93xWwc8KCo8sY5dEiNzg8Fej
ny/i/TkbkpDwww3a3Jc5XIsxQFJMWuaSX16ZiSJGjvtolrnerF2qyAhcaK0lx1nG
LX3kjrtaYfT8NQ7h7auXoacYEXKA/lqhBiI9SuXMg7xOL09lv7NHKhz+y1ukxRoI
ScgGCDrr+INPSttr6ALcrydOWMnrD5Y9xUcbVIT4jBdY7BULWVfz56uU0d3WqXBy
UbgwI95CiS4jn8ktp5Xfg0qVKf/M7k4osdW2l1HN/1KdFfPoUL8p9VgMaqAKeIMS
+Dd9/KL1tTA9aPNEdyt9nY1zizhjur1Y8+pZTL4X4PxPYhcZreJzM1s60ojE+v2w
l8ew1PS68T4rggrxZrPxoe9iynHdR3o/fu06CBdhl9B1fZgtTi7jllr3giiMUKcs
Ek/5QbpTECL08kB4tfYLbJvbGgkO9dLedwyHA412lOrMe/OgFo6NESokrPaqhBrq
jXdwp+9J61rMI5Y28Py55Gm20YXUvDbYjPwIJuEauqVbqPRPjbTY+AFVv1+g4x0x
yzIcYYky822W2/kt71WTCbllR2/ncsIYKGmfxFt1qUiAYihH7PklmtFC7hqChoSe
qryu1SQLSL2Zl7A6mcEBqFZLVDEHpzJKF6xFS/JRYEoSJojuxCsk54RQpahkRU1W
Lv4PuyfARHIz5V7Cg7iu49oU+q6Miwe7qoTaOBSc8b/ETrK26eiac+hNoWVQZKCU
4vSGezkCV5E9w4fjz00e2RgnAx1/TCU/HIFDUfTv1bESFqgafsEBozhc658R0EkA
ILPI+uRyBEcbf0V6600lY+hD0bQvq2zZsy1GUPLtPFZlb9KH0R/3H2q9hVmNu5Ro
6C4AEI0VM89cu8baaXvaSKMtbj9L3rstc2IU1/QWjmoQyB5ZsgktiQTR/eFCOrAG
bX/9ihlBRR+gkMRJg19xeLaqKqq5pCAY9Dk6n8uYExFESIbvwl+M3kHppwG2ME23
d7QN+oroNe2AUPpWhBpc7EMHdegsZvQYK1JLTFtSVr4Qxybk05JhchGrnETNU5lV
q7+KK9veBx9/+i9K1cY/yGHpFB1IKFErMV2DebR4L00iLhIX+VutdOTOJiHWMPxc
6MStU1EMemnBwzs7S/AVrNdLhKvBReLTd0fxK4S0v+g9o5qPqYGptJqzztYPSAjg
AOfD4U+rtuJo3iNIKhjcJBcTcCoMftot/1XfIMAV+Rz4TukbGajXL7zu3SSFHP1K
jdmjO1+LVxANl3S9I58CAzXjhg2gu1Vtg1tLRRA1A236Lz3Kh2nd55ZFgZrT1ugM
PETm8b7GhCUoF/SMq84wXRNtexu1RTejlgTjzZOXXkULngUehIqPY8UpINjMIiNY
SFzSrPZ7Eiz8o9dVkpM7TgnbvuuA7GNRI6PQYHQh3/pdIe2BsqxIpAnL/Cfp4iRc
il5moTqJtdgdCi1yK11DzVoZ4Wr8eCEx3HBCU1vioNROWPTn1uZacE64TsAsdRnU
zSNCjdO82fQnLo5+eG+9sOmNjKFJOmp7C2ICl2itnh66JCJ5m8phJM4VViY/hw1M
XyWj1jGLL9DyWM4/9WWcQlqcOlAxJ3NMms96GSxsqC1DMgLftWNxuKRC+Gr94Eq0
t9dL2dQuGvOlN12Df+h5DH3UDnUTlLK6ujQmzCcMX2E1rpSJgFVTwsgvBrcRMCID
lg7yc1WKPO5zHUYEcbhG9U9E29FXG6RoiTSDaLgZf1MUeOgCfLgVDIFBH/PvWGeH
yS8BJKvTL3qTwII8X96o7WJ89E2wplsp0L7ECLv/pIeW2Kl2KccTqNA7fBr+opUf
+H6A24OmOWXnRxR7tngMX8s7tNNbYN2H9ewu925MA2WE8zDTn959hX0w7M1MHQUz
li5tE5glCNeuuW57Vxhy/FDVAlTpE5lw5lY++Zf7U0S8745bPiS9WQv1GDA2EWPo
1+PNlclF2EaWFG9aWVb85Hp6SbnQotbjACGrLnLuvU7Sw3bdeiadAbtwQXj2MY8y
vW6mcwFngwAoPMMnEdvaWkHKEbzy+KnjIvE59cJz8ZIBh7RR1FsxcpMSo8pn3gxW
j48/y8QoyrgbKxYckbKaXoWPEah7Qv74CgUowKzAVO6qxhsqopU0rgkLsvZv+O/n
ruLKv30ehC6GYWEk61CBgFlAp/WWDKFjMIKDe/0C2U3jutGHFjxJPLIIbI/L/RsO
OctURjuAlYP5Rmhbt09yiPqmKqNRcncjOivOOIyFkZh6IOIM4FjZzHhrtZvh1Nz9
QXp6K4PT920QP6c71EmRwTbCUQtM6S1MNXKogzHK0b6MEGeONEWHeUeUF7AjRNrx
EG3XTa0FFhkwGi2s+v+UZTvP4DKizx4p3C8L6xVrvDuhpEDelr0VYMqxIjg5wdjC
I+FtlI/DPO6fboDLO9X/A0v2EXHgJpKdt6tPRK0BajhNP81JvuzSQANflqKEMZRj
NF1AVpyvtFG7Bivm/tlsMitDzNJfAZDrO4LW8KNWSUtrk6L9j6TRITCGgLQyO25U
KYrghbLbuXl6MFWyn3BwMaD2Mz5ZfI0GhBu/xb5TPlj21EVU1amwDs3GIPUo+d7B
SeqUnd3wbhjUgJtPm/DWDbsptppW38A4zSK7Dk5pNOrvw85WJmaQjXuj8/t8XxKT
bhx4cDUdsRp4N22dzpChQzEZiTV1ZAS2jAds2Xs9b0h3f0AIbnTdLvROzocpd5CS
StRtTbI0Y51KUUFzgoMueer/3gGiCfL9eadHt8L9mExnY50RQcgz4J2MkUol8bJ7
pDu2v/RpO/MRLF4ZBeDQtuNKckTv1q10ktdf+9KkEZi5CdGxNvBeSluHSR9GWz5F
HaJ0i9Bw6Ncw/bDDYIr/UMu8s1o/kmPUtmNw1/hHXrSDz1ui1AbZy0iVZpXQgEf0
AAsHtbys6Rpu/dpOpD36iwUAIQ44OHn4UPXGnh90br4Qyl90+TFuuQwssM+0Hp04
OKQbKXv9jujFgt53tRzRgy9MTHS+5vzfNpc9+oAy8OR5DvElBpWfB2+QdT6gddPI
h2bbIRb4EjwUr7nO8ntlxNmEufuh7HQ2J/VC7LxoP6QRraC4nJjbWaCH4fPVPSfS
rY3uAJhD2+G2GTYvOkPSIwXdTvMx70p8m7+J0hZH9jpe7cp6UwAyBuAbDeT/ZGkT
01U0122ry7Ljyj/LDMGLZMqOk9l6vCOrWMAEQphhTTSaD2gATSpvk6TxgU5qgCbR
aJK7V3KKe6qNuUuEfBytRCglewbdh4WTAdJFTrjMC3DmdzwsmYgU94cB9GJatVCi
KYKlQHaAxpyB/JSUFlRYmuiiUJcVaBHYlt8gNuOYCcxhCL0Pa/23Icalyn1KsxAD
x676zI/S+yoABIyQQSzYOsmAlsIODhgWrlXEamLxPhbzhCAuMxofJ++tnOD7QMgg
UwPf6kvLJpyYUF1t9UWiXyBK5CtCTI/9IHraQxYKeWx1WzRV3bTEug30GFHZdKv4
B0Jv0qKlTWt7dbusYtCnbfU9kNTqYBVXRc7CHOQJ/hYHXmsIKEuPaF9dyi9AxIZA
MZ9/a217XhfvK43uuK6wiSzIgApifXj712An7Xp7jtj5enoUk40lBLu7ZGw6GdKv
sHRPKIBkitgMgu5Gm8Kk3MTazro9J+d3Sj3LPf4VL5V7FBRNUcEltvceOwL4Ayoi
sYIEq7lrTZok0bVWXYffyjESXah+FMQ6c5a+qa65nYpnemigiehPSIxzn/VHr1zb
2hcyIRi3O6GhjrXYjYpFuepSX5GQLdKVK71TgAwkS7M+cOJaBdVPJ9i0WxX3JzkD
lBWAp9/++4orCIZ8xNcIm9+56aV4X6GY4jPfvvsjHcbx6fzGQF+3Vv09I/VC9CvL
RXTbyBMHmroudPHupYlpOsB07P5q+j/KRFadFyVCmTEm8dYpTC5s4K3INeG1HBPE
qL4GYJvJLm5EPfODteLm+WT3/M2ep3rL1us4P/7hE5ed1+8f4RVBVaTJt/i68a/o
oDEPkdHbD80l8bYb0CCR8r1jWGPYJqT8LdXqViZimOrvwPOULC9Rr2/e1GFVW+Fs
NmFDMHqB49qA+MEvpZEM+mghGYiFUsJn81p9Ii7NZYAjDXWnuJ3D8SuwSiZyY7XT
XzV6oeROVbtlhN+ov03EYSvoT3pbLYpqi/hWqA/9FX36bjiMP2Q6+M6wEvvuuiTJ
vJMbkvjME42/ElyRLXuuwtnHyeV9iG9ki0GTzLNegpMKfdxGe4LqyAR/rgRIz5r0
VrnTCoxKuWfIH3wek5l54mQZkZmsHfscx3k9n/EV3v0WrMpTZE8eLs4F7Gj/O1U5
PWCrlI0RqkErJSiF19IsYYtyZhMy5w1VpXXdQEpX0imgKZMLPdJpf9aKF2es8oZR
Lsr+Cz0R0EhQzdxz9sSAnO7IdZlVebL5L207lRnbK1XDpfnsWC+npGImogg4TEud
4vsU4wpzcKb+5YdF2sDRsDiachFshvg6tnGHSRSVn4wwihvhLtiuSULZ0Kfb3uG6
hZBFwW37K9tjU/3tq43jUSmc/j0fDc98dArl1sabPJRETCYbaUUl9qlKCGJjPZmP
AunUPa8XTe1HHsJeYbBoSlejcalJAFdJtj2qKywsQuTfWpqqGdls2iFa8DsOqXQr
bJ0UvF01bXyIgrz4buQ1eAJ0vkrGD+Z4JhxKxtu6ghvgmAXsUoBZ02hG0+FhraRU
UsJZuz4lhpp/doF03HCUuT4hEcxO2J2XbmQNOuUW79dzeMQhHanr06aiCidVMczW
CcaikhgNJCQhI4oc+y8bGfPzJ5yNw8Siso66UDiw7u/TO4lP3F7AgZ6a0jOp5a04
BchNzo1iMmWuprUDkYeu+94vr2SZTssDSe5wUTlUjccU91WaZ4xM4MZp3+KCq8ES
IEKgFeC+A0d2iYpioZ7njtzkFAyYySKjKNuf7F1sZKMoifDYLdyxvQhLKfiby1G1
Xz/aScJyueursAzuJKnWkiMigqALwKckiVvNNQEYErbz0cgla7Gr/69vmQXrIK2p
9adJWjVmTpiyZmlNH8tcBj4a+ii/cL1LUMX3pSZURSQQ9llsyA6G0qFUyibalTvq
ZO8Ptt41ThBLefll23BLi+rfUZqFZgW1DLy3AcrJgxSGH6aO6rZTvKb8L1LIPavy
x98h7M9Hl6usS5bqOXKFmo8/EmRk6bp01uO4CWML+sum8d0fndy5qyNEiAoiIZFt
m8vlqCLmktCurORYrciM8DYJmNrgbwVGXFWXrha52B5UNrBaPdJZB2xpr8P8KluW
Itv5ZpiJf/ZdmfrKiKGWZ8aOg8pMsirKqTX+U1rsfcKYDIgoWHJvsMll+oyG39lx
KD1hNYIhEfZYqHeDGUZyUTGB4qqS/LNZ7jhO6df/SAMScnNELZbEU5SU83r9AdyO
zrjdiSJcuk0N0XOZ9/4vpRS2AeGQo4Vmw8A1iDHyzLt4qGYbfvNuJnqie70tCX8m
JDQl651L/KSh8pSJeYFB6lXqwS8fzoGPR7A3ySRsWvr1xupbOjsK0tV2o2WEyDlp
aMDP/0jPiHbK/iVQNglOWL90RMN7eOWGbPO3xdejt5nGvU1plYVOthi/ok2rg7iT
bu/2dsNX0okWeg46QjwDWuMwhMOmWN6AEFdAsgXjDBZ26m3W3WKWdj9DKvGXuy2Z
4nRSPgVCmJcMP+qHqCUuZfvHNKCDQ28nd3LFwZWArpterVljSbvfglxx5HXifT2+
9oT2yZ8WUQppVHXt3MYsao5FDTwh50nHv83Sin+nyFfvk+h2ezPzM8nSN+nAyjPE
SFi/8plNXIh7A/cJBogjPndAl6BRGFrQWd775SDkm6VcFb6xGS86mGr8r57p+Ww6
gifVJYV7jBJFcu4hsaU8f5Iqc5tcJx4gn39I403nfridrgAOANHv3tc7j2TcXYvw
uTs/IOXZPZft99/vDm923C2qCPUPp19suvsXyJy3hpWBhIHChMQuxpsB6l8nnt0k
zH/lry0LcREqSJUpOprJD3PcWMDM4d0H3tCSUffccH0s9e+bB8kUdsvWDuIPm/BG
/EoJbEZ+Fch7Gdp3uEt8mAjp9zrDoUB3QLO/BpzHAWUbe3Ms+Cgr0juSLBNsb8G6
bu+aGgzVyYYRCn/uwnymwauVTADF8s/89KCOyhyfX6x2wuz/BMYrjg+WyHJRVZb2
01yOf96nQPa4RB1jXIE9IATPAoWM2xPb18n755G9ujNWSGGf6se+5QOcBFM88xgT
Pj5vr6/Ksr9z9gFk5qDLJJOCGvqd7QyenDyGcGSLo48OeDBnt02NZqVajj555zav
EMCfFMrzCdx4hIVIKoJqC5356Qa7cvGQvMv9GPqckPHihRzPFvDmce+EIsZIy4lt
lhaRBroGiGvT4+R1CZTuPc9k0wRy1RgGWoTdh/Q3USSH2TzHFL2/bseyNOs+x+b0
QobihlEOzw/xEw7FbUDGDRK2vehPVhWNLxxIBDvN7damKO0kyhlWIaEEGvgijMUo
wVQbOK+EZPWJGgl40QSUA+aihzCZEU/oDYHPHnnULkNyEDZ+DY6AKEyTw+NOJKY5
pW1vqqi1ZyQkIBr0S88F5+Ku+QDuefva1okfA5Fi2GbqTiEkW1O+Rr4TH2WoP8Vc
mGyLkoQo3KzH65OA/5fQqTsyahkJGbF+KHyxwwlyKBnI/6RiEcdjqDEgY7sqXYEA
c4ZL+muNVugWiP13/buZLDLrhCnQ9iqe4tB0IkQ2Y0JxqJAdyuVfmVqEwTmlSKMH
YTXQUFU1CC0c5OBAitgQY3DCzhuzmx7360Sj2U477cBTkOYOWYE6FXqQhLeXEuNd
pZBVg9Q5h+CGAhYhjaqHStKeJo3UZBOKli2Z8iwU30b4Dj2rlIpaOf6qW1nhMRrp
dEmzN3s+3lXHRkSg6tyoy7eaqQkfZPepdzd8xQou/PE+Kj70KmjjjhPvFNLJApe0
fUDUhhOL3NX9qjUwqFITwMKBYh8YafCWLA26MNEAeYRTIFC2JthSopRKDcQlyRio
MOCRHclPmWeNu6EamnntEjUtcfkcrRHcZDnrJ1hARtTsQBnMLqt270JPCFbjTENv
zt5qjI5ZThlew/sZCJlOtunrzv+rUBiiE5ch1x0pTP5tmZQm6/ToNoWoh3XweJqR
PYhxB336i6J+mda8adeFJPs/YBzMIWYT+C+EAKwHmIs/wMsUKdrD+lvf98aystnJ
IOK1xOewMX7cc39+3DUnPSmmlfhJycE8zhL4bVBmCSSHW4y1YG2/2NC4oAIog7vf
kIvEhyZMH9Wz7uyrdslsv7e9PPeuXCqwnG5NPQP1/IBH001H7qtQkr6Y+lglFeP5
cEnB4nZoVwF++jqYM67LtavQKe+53q4Ty0ebrBmitO0NihHvNeoP98PJeQE8nlLs
T+BTF1by46WLBe7uHuAT1WNAS+BwWO/fs0m399A1NhPI3w2RPXm2+WP08OsM84zl
j/MDORQEFzDPmfe3J2Xfjgi7NRb8ZkktzpCmSpf5n8f6d0t3XaxvjVM3yPtEKHiJ
5hyeRu/Qeyvf5BttDxnNyKo1C/so24Sa+YNiyig9dagxG5VLYv4we7ekD1dKQqZf
TJ80dBSL6Ngqmh6CT8PkttslKQxihvhPmPecJnH3v3hfyuDkgaKyC/yO/wh7TX2Q
7Pw1vqtA7cxWGoYsgltWr9G6joTNcQ/kaLbTglWJ0X15W1yOzct1yqW8MeNQIkur
YlTHfS+Ry6jqPgTmo9eRFsDw86BlPl2oiLJa2q8n1p2BR3WB9PaG3ir/KmGmrOi6
m6hiIiQSFVmYRIXh/OLiQP1t3XibF+/juteHWVRytkaNn49W0MhFGzlpbvBaVrr1
3YJ5+/DZ9rEbcTA+dongLQqIckHQZ9q7XnjNmIb0yE+kHJXsX16XiZY7lRg3H7mL
7Y2mgqrt7URDMiEvSu1yfTWniiqs4TR0LUw1zZdHCYSCg5ER4V79u6hlCBba99Qq
DPKwztPlYgjvqA8+EeyY57cy9xhT/TUb5bao5LFvPvm/HXuxRUlo4ekubcydMgeO
gA6H1RiVVKhFKTL+nb+F8DTw2oej5F8HFcHYwAXqbhK6LT/KdItPD/v30yVaQuna
G/o2pbfAc4GrMCOLphWiakUL9dKH3B8rUQ34UKiSFsHcy6HKlS9mH77zsy4JiZbU
eIvICwxBbcD78jjzzoKKHbQTLid8lRpWKjCt46Baitv0fuks4ZAaPNKPVou+/Rm7
8sW2b2npCW7sagXT/xp3A3WFiuJT3KaWzYb8/drrFZyDJ7il4CPcGTnaqvkWRjrm
G0S3VjZutbG1vk/chF/qw1VvA9ii5q7w5kCntA1Jw09OgCGVLgNHgv8lRJ0oIEd8
tAAPT8JdLhnDDBodAa/q9KU4JOGjd4AxSUf8MtPkPNSlcUvZsHmaZCN1uwEcVrI7
RzegyOgCN4nLtWj9hO1sIHooyh+ove3wuo2Ug2SEwx2q/074hnYf6/jJ6XMTz1Uz
yOORbOfQHVd77w0gFfJwfsrzZQ1cxmJ9oWJ2uEfzEeFLMAYwTkf+iroQiSpgpbw8
8ezND89jnE6umGycqKt8nZgzE/BJugqZ5CHtkooZOyxtUiXvev6doGcmOtZDdsaX
E4INwW4SidcucI57hR7b8vxEuYxORe1Hc15b3vDIq7dRFp8y1hHs9ZEXfJx9M3uw
xz+WdfqWNAZpYFXk9cScefySTt5BcNdZRU8rK2eX5mqvd2Nu7wzolg8BS558kdI0
TsWcOSU3XrVKlyFszU1Bog+DusidJOU/7w+tR1cK7i0Ntf9KpA5OdEM2itIOhacl
uj7CkNWeLFbYLNy7NVEQz45eVRNVbE1i8NsSuEJCKcaIYrdWsVB63uC1dkewAiEb
c5WRWEAJb2mB4ilZMwzB4TgowHrq96Ickp+fz2/u9KNkUowk6MUJVs9iqY+dNBWL
C+3xzttM+Xv/Q59ihUWQ/ZxnfoZt4+EKI2gxuVmFg7EFBaI4oveRepuZy0hnUzaz
eIzIgLn5DCuNIpwbV4MPfm2gKMuaZ9JFq4EejjUNwaLliG9jKG3WOI3hmy+n4kRS
Xdmv4uYPcu/RM1+ZQla0IyIMp0Ah2edow/C0kmCv1y/VVrV9rlQ7QBDLw1X6bxry
UbJqIzlRllfpUq/pIRH5HU42pCwl7krtckTkGAbWrHtCLQaJpgZ9kF7SYl81vZ8i
J0DIdhKvdu7HCRnxquLZQC5Qux0TYWurkXljUuHRx8hfaeJDt3xGQLpN1pj61Jmv
wlTGIbGI8g0gjMEqWvzrWqYFR1Fu5LN0Fy9RVPkCDYckEuqjp0Fw/TyU4WCHTowA
kK2Tx12pnEUR6J1H+GImgOdY03i5gwIl9UA2Jf29s6PJ3TVpJW0vldkdjB17U0g5
Xu5QND+p9gK/HfGjLi34GZVajQbfA5GV7fD5eicRQ67ijqB8gqnCiqBQWgE7WC5K
vMJOXaTYO4sh2vwETYjUu/xVpEwYYQwbaCE9X1r1M6Vf0J+Wwp2qjxn4E3hysbfG
xt1FQpm4aQkbRyIvIHonsQTOUXTb80BpnPzsavj62eUHnlFmidxIUTCxgIOZjTJN
Rw08wNRjFPkIo1g7cS6iHemcPnmVBQsyXytQSHV3/S2kmvoqx+ZvzedwW8GqBK8t
nnC7ezqo2D5yUkYnAvIBBPUeLv2OH1qPuhsbljU+tsxXZ22fXN5R3WNuzK6pWz5h
9RVuN0a/SXoPVWvR+OyrrGoriS4eDS+ew9YUBIhVNMdv81G0+X2KXvxugdwBzZl5
g2ykC/oLuUv+s1xEt1W84WOMAqVqwkCyYLeNEhMFGJO32z7UsJgXWdCsOoDkGIMK
WLDppaP3FzMsBYp+8Bv9nU1mkRfb05OUU8FRw8tcw1RlHVEN/e0LHDqy3E0s6O08
Ix1gaUbFmF/fSDitm8Cj8l9YIRJeNphf0BaxV2SJ4JGNKOjV3ch0fAZhUZjJgl8B
jGjrnA2NwtHWlIv3d9HIbQNEP+1UqNR7L1iyGptPbGfrB42u60+Nv06koRXQXsu0
2HqGrpSDe6lqN5N4YCBqXzlMCMYk65b6hJRIUqA7rTBqNNL0DmdGnU4pTOn5kV2z
mM1RQEJKGpeDWNSwGjilPtlyP41sOFo5ggBQskJQDolLsvPo6QPPo39h+0E3DH42
91jynOcpQVeqlxZOJntB0hDaE0Ukzkx6ibXs5sRsjSxy69v+5FigvlImXg9Oi1sX
nFZfj/jtA6TJE0FObfe3VHPSCMj70gY7BA5k+OjV89kvBaC2AVbp9KfDdwq7MSiP
uYOSS2lw33nSceeIy8oIFMeKa5pTvVFxFiuk3exoYecMO0ZPP5iNl7mnlxRKCeWd
fBr1EjB2PWkEq4ZYBFENNt1YQ1G0cDEUaXt6choKpmrbKBwO2dWnvuJfkXFPg1d4
jq7qxhHYQTcS6Zl0nir6mxzEWQvWTvdXqTk8He/CpH1PHmygJJj0urU/9A/esYfM
ACCtg4xt+eNF0Wb6VKRanBIbJ14ynSvOAkRv1qq2zczU54DD3nd1dmTM+T46k1Cy
m9j9o0E/OlMfjjwkQekeICpMQpwxpypqIhLbTECcq3v+vy0XAdiFtbrUmSmCWvkC
Lj0Z+Uy7dilCkOTYg8pWe0vYegSQk8vvhi2w61n7m9C7AUxLWUtsoTkYVjsfeO4P
8QIFCj42/SGJ36yhQ1pgFdDTrEtJtf+1/Y+7FvjbCrEwgUQPO/lZgX/N807NV++x
OqSljki369V0KLZBgAAEVt/RPOB4d4p4T+xMwu0LHgcSWaMH5r1bI5PZVCvHFnfQ
ncRDSt9OE+ilF6VXQrQP62lH9L6pV6A1uvuVN+h5sW26NuSQVtDTJYRFjfiQKANT
lUK7MvZKusrsPqru62kG1rhlN5gHDu8LN8wiywq+i0oZ4hz30NmIUbN22PWAwGsr
J0iqTfS3eq+HAWkF7mvQeY8iaErCbWvQ1RsNN0uXxmkhPm0PKo8UK4Fiz8pWN0xf
Nm4ei7qBiZOeVff9scvQcc4YqxfA/2k8d5931Y7r+C4U/QJwHX4Pl7VQMb8Z17T+
lidpi1nWEYi3g1dGKEEbaGFSTM+LvcPiqv8ZiSxi1M/P6Ms6Z2SlFbqWlXoE2Tg4
rQRM82J4Wrb7VbOTmQg5RDXkoqRtu5pL3DrtSYbdnHykZz4MCpWUw8i5hbTV8Wa3
7pNr3gXLBQ8TxzYkhQYiekA41JmJGqONZJZyMkkptrCqIIsCp6DDBpPRw5fxbxsD
U+tO//13cD10HMtXTDPmScBSPPu1a8R80CAPha7XvqMy7w3ZJ8Zb/L6F4wV4P7uA
/sma4s6flvjX+brHqhYWC/5xuIRzchT9vUKaxeNnBQDO0XGQOBvytBOEw85GGCtI
nZNLSfBvRng1PbMyOHXhOR6DeBq0hKi6ewqLQdHTkb1/bA1SVStaSc2qWppaeo3m
G6fUselX4BnoYIo9siGjacEaco+tnexDHxtz/Z2E3OEVG3ey0d9L+hIK5+SaqSlQ
eMPF07YMfgP8RICJlZo2nXSW7uZ3DA3mvzKPaMEH8oiaQeWaw56/CFpOwt2tOmGG
x0tG8Urbd5CzvtGKpzVHlY3QluRVO1CZ7puQPrHA8eDXxfy/ejjWa+b1TQ3ZHAXr
NN2H1CcREaMoiUvGPGzEHAbLfC+TsLp9WcPAdJjtfXmUxPjGEZcLc8q+47GfNE41
FnXv3ot2mQVcwE3LNpoZfG28g+Cp6GaF8lzlYvOC/ORIBwPkb2uMkbrsK+kX6Dm8
zKd3pEVklTuGPvrFzL1/2MD6yNoAvxeI4B8IIMfCAWlBTP/pLqxaZTEflc/Rx03t
i0qLKBCFtus8yBf/6urLITb1bwpNvjWhTidqyPBwUkjxWx5fvIi1TdfHlXs2TPUo
H4LNoDQBLCjeTG6U8UjzVG8q1T9gXlDWra9MJsYt0zg/5D6oc1istpVssZjUXbdZ
JzAGZvuMuJwKqp4Hih20TGnl7Ki/41BzQZhav52rIADHojyq1vugDchpWSiwzfKG
yFqdok0y1nMTSdhLDXI7cB8bQeitY78HAY+Ux3Zo/Z4c3KQb/LjMe2saWVoh0s8f
XajfcL2SKGP5L2ZaXTmhwPDQTHL/ci0ToRyvhAUXXQPJmeO5x8Wc1ylVEy7jPfSQ
XXHAaHKyS9R+SEM68NGLHKSi6A8e9R3oNDY74o0Z0S+zcNUOKfz+JgdA86oxGTfG
g78+BZK6ppm1/G7OilU0ilB2VNfWLtXHUjRpwRC/eilPH6Jf08JNhj/78MxVTujg
8TnVScLS+l8GDr7AeVvVUdMTpu/wyaTJZ2TLovVPLhVgJPIPk70hR6VvGM5Q5ZU8
aGn/KdJcsoH4fSVnq6RdjhKZGrOGuNDCYikN9K37bJ7HDAR+nteaKKsEMgAoO5vC
BVSzwBSAz0DxB+uDbgZn4JVGieoay4I1fuCvlItGetOpHH9+KQmPN7Ce6xwIU1yH
E3b/mYYqHSiKXLIxNgk65JP9ONyN/9fpGT5DX3z4o3WipqWtrM0cfdllnyYpIu2b
xgDMujL4cVjA6hCeHk+Y3NdTygac/Jf3HlJyuqCJui9Xk1IMHluBFjGEPLmQU81n
7hEBAF7fUbdMUoygRf01ldGQ1bPi1iFe7Dm1prVcz4Eu5CMeEzNZJMHiMt7eO+8B
7ENsFHFMTq+oLeyVV5yZvHSLY2fuLCFKY+mKfwb6p7jCji44U77RoXMvBgjK8OjI
RVo8rwoSr/rc7HfU8RQsup/tL6WXYhz1pBRHVjse8Tv87DXqWXe+ykSzrfD9+cZw
EB1YiwQcovzlx9urrSMndCP7Q8GKP+YaC2dXvGHzQUY9dCSiT25RLCw0UUaCaW/T
TfnRS3AGtsQDSgQmp1rCBRAI1HryYi9fJ9q7x9sOB8mOBixGSO+VfAXBmdnARm+z
wtR0YIQFVYWIl9/sAx2gLIiANB60bM0q5oWc/NeUO8ySKShG3ul8b3DOkkBvXvRO
e9HxsgaXt5Oy/n10F+py/fNweFXEylCNFcI3MHbNFa/+ZE7iR0riBlWJJ9fjsVIz
f9IeUz2nLKYA7C/dT9X0SlLyWgaZopmrJxci1ab9TsVzr4aqfUN0rbi0n0n84taP
AxWKndaxHpqF/J7RFWNLu2nVtLbk8iVZ60XNq+FSr5JH0KAwE+jomLOlGkrJn/U9
BRCOv4NC8/tsVsU/KmohvbeIN7U0Ea0LURAXErD/VyhyX8XVfNjAJX4tXddTR16j
5+wpSTj2I5rq7K0A7llEy+oTZgKb1rfe3FUTyS0bElKw32o8deLjR5tM9+wqGz+V
dE/gZC0/lGozttGH++FpwcDIXco4RskGRlPCmaRmGZp5r8MFKtTfWaTOps4o553n
c56rFrSksY4hpB9NGO/uLNWupL54JM0Z75VnlbNmgmMXTalxiSlMWj/4PBC7Uju/
iXl9Bb3KIfDg/phHFYcUkCYtXD3M/o8pLztmegwV/uoClyBMiqAjPXYv80ysUYFP
Q9Zec7X9SZedEHoQO9APmBlS0bLIUqOd2k4aVsAwzODfEom6chdpG1s9Me1oGa3b
iMrKtsISJ0Z5tZE1EN7USOqSSA544dcZZbAOVsQq1oEsZ2m1HUrwx3PjP7S2orY0
67rIefU4DWLXSLIM9E4N4rZd3eSit9stRFEseUF3vfO/CyAaaRrdSV8JP5DSI6R8
UyzQJ8NCGLLBm4VnAjDF9uQ4jYInsLD3r7JmEVfPhTN5iQN0lLhOZ1idUKK+b/gg
+gE6YkE8G8dvSAPidJrfNbopl/OELckVuqzuKk8JhsEUl5eh2hzOu4EjIcQbiZeo
dgSxl3rHAnGPGrZmjcL2/hAeBdV8eXCoJ+K1lbFT+B/twYv+dM7vfD8/zVTuuS8l
qXxGTIwQu/D5EKSothI9JSMYuSreITPEIRmECwCukwZl6RjCWPh5Wlb65XCKESME
a8jn/lKkd3BmFEnNjaeW3kyZ16yKZTDSrEHIPMnp2IDFrLKAmel67TKdrKmtf6SD
2edb5oH0CCBYwn9qVgH1ANRJXMtdeG2a+EOFH1ci0WVBGax9Q6IBgAQz3VbuLG7D
egDLWutFR8VFq7bOcCqRMFNah0gp8/5PGr41PJm1LGnqDXYQ3SAZjgsowsduPdZp
s8Kit7jSy34u6wITz9xKLz7541W077JP439fGtdxTOfT6NJbWwb44jbz/xjRmpau
MA6vGkpJ7rf/GxDhXMmuT4y/0hiqYly0i1INHno0ohjuiNJKZO00PB4cCUXylzeS
hy+qJ2z+6QqS4ZoTJDFYkAvLLtw3YsDzotDJxDa8EXxRZ1KqQoLrVGOOukudUrA+
hZfXziD81Ck327hLq6hqxD9sFGiCZfDe9X3K3gw+78OOVbGLhI6DfrXpV3j0+Z0W
MMD1xcCS7suB+pBZg/w4GgbxwCg+7wCZ0eSI7c+Aw/qIty8o3QSsCvSk+sGZgh1l
GWv+efu+wGU9/wrLU0PMBMNixXSDT8OxUHsvSHSYVtPErrSRtyvbRbZH/osvFfsB
DzkPSzGwXnz8Cf4laJzrYa28k/DJpAGpWWWq4OFBzzx8Dx8Eu4SnZ2URxOhbJEtw
Q7oGLxm16odzvuhCLJm1exzHhxKU25YNMCPzgIbqhN3PcIPD7u9uTBk3WSNkrO6u
HXr9ysfnSytbu9FFjQrJVI0DDguw5OuSclztumQMPUzLxt0szHgPNWzES8W0pf+q
rPLy/NMm/g4M4CN/lNlbnjsWNa9oKMjMjQomkd3UWIVhQ0ALM2kjt1nO7GFPEzWu
4g893kw9Y+vZexVZzY6QQxW7MI08YGlRwV/x9cQVWKAlW/7zjsgNclqLob7D5lko
AwzVnnyjvQwNGDKASGZW6FkeV0ih6g/0Za9Jpxb5w4o7npmdvOeDuj3xs4jTeNHQ
OcEP/241R8YOG3zbaQ4NGfrEHsX5I7JaR4YoIEQD4e/fsjo2bC6oSBRjxjogdqXC
Gp0z3ljSPDvgnMSpuOMyEaYmLSNngDT3gNcyYbSQ2ccepmjPQ1D9Xx5Jr8u/PxhG
cd1awgfvaEw6HmoTzwspMud3qkx7tCSjpN8DkFgMZT8JgUlA89Z/Jgbcq4Em9HPe
2hlys1ClDLotxo2vKmWTjryRe/G37HxHXmoOUR6hXGB4hPgM2rJ+8q5M3hfUev6C
mqnVo7l0FbQBsxhyEXif9JAnY4yfS+LH/ZcVQ+uIza5pszekGDJfhBpzO9x6dsyV
c9lePgsxGjl9sqOsE89UrCoFrAQaVRqH1hB7GcfT3ak/pZ1j/tQKlM2uAs2rt3eN
Q89p0L18rnxXqBPXjuXe7Jac4tyXLHvL1eC/4tcJ1nxVs28WjWW9+RWXIkUpqVnB
dsk/13fVqboDiLKstFoo2ZTGq5XHxQ3SGzJtL0RmMkwj7wR656bqg+Pf+Iq9etQ3
LQaKCG66uXyyl7YI05mxdsk1mi5rtRwqnTn7D6977sCMkPzk/5lYD8QpT4xqmW86
CLQnXTBO3+LxCg4+ceDtEyen4S0ejITMi6wH07t7Apkb2hfsfGYMBwIY4gOcVIO7
22ttMOCMiz3vKSlISakO+IsWffxNolv1f6J0kEUgtUxQ1VRp2aCqhy27z+p52wtM
8oF51Osbkc5fUIU8jGNCi8C4o41NdDZB1AA0rYbJdMMoJzYrAq0boQkZYmKxFkc6
EWLAkW6N2jYVsFkRAiCizmU2k43/GgFFSMvoaEg2/NZqGPcsCwkmAeitii7Gqfoj
B5AHTc3u6tH9dMBJ6jFRNkxTNOJeWvWIOl7Wx4nOAKrfANXE2TvvZ2e+VKgsJEim
YyKb7Cs8aPXgv0nxn0odoqcTyaBX/2axl1EtOcqVdBMNU1z6wB7vuOx+W7m/zEuL
uXfxQr9QSSjaExH2m3ILRzxf+FQrPqgEDWFucnf1uhrYcB2uqlsOGHgfS4Aa7tGL
TsQNkft84uMuGOXWbqEyb9Syw8coPQdVRUviYISCJvWh/mnZ7YrhlC59I/cVn5UX
6jb9Sa0yT6w6FHetKjFADgoI6lVpzQmHWuJlf1v6rPjePnJFvosMK8mIlLsxF+tr
4Kugyzuf/b9VybQv+nVoDD6bDgaZb/pkWtI/r8auXX132THrcJrQEzIh2jLi6bNv
xTXK8KAeNNen/7QFkla8LhMKAYLHquxfBaqMxTo0vpd6Sxgz7m/7mPguBKSQKVPV
eWfLQsYlJpjT9+sqcvAKaBi6vODxJ1KvF7JNNC4ncWWbDoU8RfBzr1FV56lH4P3D
YH+zilf2XbDjcxWHfT496BdP8dKOpPu2T4BIzQ/Ts7hg4xd+cNjZsCJmoO6Qf2RZ
nzjekEZNElxRGO0qeB23Ea0FfctUbXTd9jaIrQcELxGQA7LDsGB73nE+fIzA5Dzd
rFHvJrYbUBEuxDz//91woMyxHf+l6WrZtuezEZ+RXLaZIFAdZW/57bqt9C/GF9cd
gg6wJRwHH3r3oK9uI6PcNuITSL37RD90MmpM4sLi7QO0a/OIT1ZykZYZbb8QW2zK
fr8208mcjHFpwAXdTGd9bPBVtQqsIxfcxmTLuULgqpKH5Md1T/qEGRyHfZk1kX1O
+Fz60V9xeOlfwGn1bgCItQ9vlAoLmrHoVG/FBl32oUm0ZHezxq+UftmxrikQyp2h
oXNo+p7N5d8gKYIToEqz2GBeS7pz9UTe0zhcYpKAA8n8x9RORrP7rc1v4SVwSxuf
Lsr1zOucdRbyfqBz/6dmbDimi2MzJ1SE/pjbXNzHASeGgDug3Xyet8/6ujNJRxv6
noD4zYkZCpYMfIrzv9D1HNfnS2Wo4WHC3MmRIleaTGVs94b7uQFQy3TuKk8koxGt
PHTF2FcSs/Ecr9hoMbgf/JEYw2zDJleTCqCVd1Vb+4J1KLl0449E2YdR12ksZlzX
W23u7J4xDPcok0vmavwYoENjVLer64aUnSm6iQCxpDgyxkW7jub4hA9BMiCrMdZT
uREc1acC7oH6XOaUj8K8VyzWD8xmClLhKGMRxFxdHAMfJ43jXg7p8TRbXttV2rBg
uIHjgJU6s8s34ISfN1UJXsWzzK7KYp/WoaWTxchVpcbZYHsk/FuMN6tRkz5FYCi7
l1esCRL6N/YOOZb4xLfg3fgVBjjNLeG6Eql1pJYh/J08QrcWFBv0pwa8F69bUNJT
a3TMEMpBUTdOrZ9oWW9H64fnuoLkaBcV27uIKVgUJNpgoQqANiS7J5lgUEPCpSVl
/4WaprnBAqGcgLJuQC1RsFTYeSwxcXCnevMCoAv+xzVHAZlz155K/ajhXvAJdsfT
Ry0RF4b+VvbEnU652SzJhbtz7p0t0ACVsPj/fBXquQEwXsG+bOHuhGlkjTx7h1uV
B0hOUoxnBrHxNc7KVgw4t4xPEvpiy17BSEg+Jh5jswliMPhlldRbYrmf4GvPdqk5
zK0t83rhB10ukwa7uDxTDJL4irdgppzLooei/M4Qg/wq6Vn2lY8cckP0uc4tJJ8n
JlkI4hbhR2JcY+ENuLLwTgJJYjOvkfugFadIAL4zWNTST9WVDzOuRQa6/MoJL+1F
8CxXpWMP6B0WH6vjiQw5EGxNc41ZYmYVawcL5wSdP11H3A1JU6dBCt6oa8psd22j
9c6Nw41yWS8zXnK8CBrBjEmPi/LJlfL7Q13KEeRMQcMJWS0GGUMexoCfBy+K/9m8
8U6hesRdTxdmKe01lULP8Zzy3Bkk0bpCIvkYI7JAjOepKVYhEl9N/uhffpyUc8Py
lgBDwJnu9lC5UJ/2da1VMDmd5YQaRIYk5T8+xm2/F46j/XP9Gyxq8udGxYgAuvYd
Jnkt7FfMm9vxHb+Fo4p9ceBeLPu6YgWs3EBRIKMk/9cjXvkrMaXgrTdMwVWqyRMR
w1+SMEOqu2ORdlIOERFnaRClFDMeX2blmO6kx1dfhYZgOVX8QsK6QtxsHFtFTOA4
fWhL/0tW4Co1yJi691vnRL6pcDzkEh+E016plTzYXeHLtwHgaPsQ2sEind1s2l7+
WvZahn9nw4eo6XgriyVwEfb2cBfir5Du3OTjAGnLBGCNNB0mtQ2+kg64NPDIakPg
WdWzoh3xgtgCT+6eRfDlkOGP7+W7Agrrcr6BX6AEXIb2ean1DCNVlb9M/MRaCMsr
ysFxcrdlycEgskceA6NYlQWw63dPwbEpWHx9wj0NBjZvufhh1N/puDB82nvydyt9
FB1POChl6iLPD3VMW6IH1sKfIaI2PIymzFKJwhIx53wSdi3pWkQW13iK3fbwWWsl
6LKT4sXUhTNtuer55sTO4Nobvkepo0/BHcehpFImaBQG3yZbkLgb00FLg8MDgtUU
DkgVLjr+nVN3wZkJI/BKsKlaANEk9vVPgoMBO1ZXPtb0mq/756lkQyIJSuXuZRDF
X9T9GPoQ0IFXVgI9N+NzpuLSCaqT49yy1xXl3EHboQBepg2K45iVGvNXkdvEb1UN
FpA7K2KVVkBVpQmrKo5D/6E50ieq992egmsGazEyJZFic3z+njXYgr11p6kLPlLz
dCGW20uR+dBFpfm+rTe9nyU5MlKgDBugfE1zFplb9IPQoUgVrhZVpBc9uxMR++48
rxFxG6TTqkyehNA1PX3PnFZcZYRTboewPmUtcIxaC3PiS8CX++P1yTfPDxbqbbbb
dawKlfDHyDO8uHWaTP831aO+wrysPh2VvG+xjluxaYVUwTyp0t//byCkkSrB2Meh
2kosJusCvC2/9i/bKHMtWWRgF97LdZdJyAnw6j/4ebXqXLjwYIUnfzTIld6Q9p0k
QhopbzXSdcSGFlisXelwpL9OAtDLQcXX6IMfv7K4AX8gS4T0W/LSF9fFLmDVgbgv
8IRDK9GDrEIU+qDbPhK2G1X6ppyWrZgPS4yMFXIYlR7lOFh6vn8uOAFjJpTsLXL3
7vn+zyYzR65h1NDlpsHN40TNn7C70TAJ0+HHmFPGhYjJOPtRH1eleE7Xt83rm+1D
6wpFHNlQKquMPuWnCiE95DQLP+tRB+JX/SMPNr7nYov9q7xTY6xhbnJZtRF9x0Lr
4s/fvorBZw98VHb/7fp9pA3Aud9SdN3dnT0H0jOKGM7G0bWYux0mDu54+IEDaGUT
dKyDXK38GWYLaJJvUifG8mWd6JR2FAhpZXdUq+VqG5ZyMsT/yKDC5ON3RR2A3Oej
fkDbmGgtgSPBlalM86Qic9rac7aEEiPBLWXQC+eXdkMknlIxx7nOCuqFYyDx89wJ
ZjVfCMK/JV59GwmIgenEAAGSh4OtOAQzGdVy6ihLM1C9OyHze8ZRlRO5X1rjtzWk
8a+RG1mIUPbl/jHSoGWilNXWAGIAjDgrt53ySdv4bZC/5025qdNQ3On6Inn/f7bI
nJfKNlKuWxzuC2ygCMQv/+W5Dvni2DHHFrKYvhH0yqIgAZ2BOx2ZkTpOTCnaNrvd
wzI/FknaGWErTXwxAQ/WWU8jl3aLNtlzF9SD+hz8pJCgisy7G1XJhbNAyHRj/+Jq
rLX0Cn5TRtH7nqcvHIRd+lhhobYw01Qfy6gJEbqi4pt8Kd2769GyALwTNNdSKC8n
LuqJXeaCEZr8Q0wLcHTqT+Elsokd+lp3nd6QeypCJNfb6VgEWlAdtjZ2mhU37dfA
5mCWuf9JY43lj1u4qyIglWEeE0lMVbHkRhycM665MIKP3T+NltQJuwIYEhcLMYlC
Jo/T4neNKVtoZIsV9i1csSZR0YPQ2YLUVoB8+tRfQ9v+QFRtbFwDI6haZVPSNk+M
9vClbjw1wrx8qx9cDF0DndWcJRKaBa3c0U1i1QjBxE5JaiwIkaFPzN+KfsIsssfu
auCN18OXMfk5+iSB87mOO68jKEpLd1Iw4s3q7NpZZ15d348BYEDNgNO4621urOwW
dwmTFlcN9/0jSqxT6Ra4qIN6fWAiwR9TRLz0kFZACwJresdCfHAlJNeRPONnfIHK
bZrB3AjmKj0avBrsOiFuStimqRF+wBw2RvVFEH5Pd4XBPuNTcuIlEgI2rleYYUJt
dWvAmWbOVa4uwgTuZshsnezSdSFE+wMz4gYyOx3c3qumvm86mrDB3SAc6YgvXpwK
nrG3Uj/H9p9m7fVG0wxndfbFruAfwPK3Nkg/Pit5UXZEMis2iz4Q/5Wga78RBhxM
ai1NKwV84bApqwECIm5GZuyi/HpGNI3v9DTj9zXrpuYi3KaUrZ9kL+2E3FjSnyVo
f6J7++hagEmkb92Xk8in6psdwfLXmVtT4j/7XHaNa6jgXYWNHrwZsQ7XXkE/+Avf
Sd0lc4+bZHm49KS8oTvSqXeuNYCvm3tVQm7GyeKHciFG3nZAuef5olqpTVJQ6Ahv
JmX9iZG1CyE58ZvqupbOsoHVYzE2Jfgomgqzt7nK0tBNf+L09oarPj08LPjGNlRS
hQhX9U3+ErccGJ1/xEzOOmf6Kp5W/YGLmcJfmyX1YnDT18mo2TpYd9K2QJz0TvEU
+QAba9qiJ542z+Im/NKh0Szyj3G9e+7uyormgT/SBfpgJz7fRxB4SktDyLFKZBTk
5OtVoKf2BkQuJe3kkOiVZAiVklCPXpflyIQwF3eX/iMoXz4sbqP2PSH2/c6BRxK/
8K2CkVQZK0BPTWPulWjX58gNuHEqm8nWCJp7GacmeniZrA3qZZBuigJDOYKuEBTj
Z+bg5ZvvRiCuD7t+oLgbZ9jxHwhduUWjt/6kg72Q6FT1d3pTz9Vdy/Qly6+yORaI
L6+FQ8Zd3On1w4/g+QIpGs3cC8lsstvXR7Hwey8rkEnLCmVZ11H7aHwdvp/37Fee
VSlA3MTUMndaUA5ym1PTQAAQniTaLjX2rGlN+PTHQbulwnKwQWtyRWJ3VeB2JzN+
fLcqihhZSC40+kef7/0IVGDXpCcnC5H2umzmuzlJnYwsOGjmJOh7xXB43iFiZQiT
8Q0V9G5YzCkWlsUDdeynHiZnsvIvGZxLhTqrbg05k2m52GoxJbC4GogA47HgKTjI
GDsOKuTMzY2JoVijqSYtV5jOzXuLs/Y6dmpcuJn5vfIFDV6iNmcXI4fKUA3jWLKE
/RUu3efTzcxVfG9+PCuFA8YRZObJP7GGxaflPSqAOjxJToYDbZkj96Zf9C/nOjx9
h/mboP+zukR30nI1BUz8ZnXN/JwWP4A4ZMrY9HJOP4LWprjDtmPwb7fU/T1VKA04
bVkacCoVjc3Lcj2vQ7M9rsH66cX/uIP8S5fj5qGtLAn71nDm3WnahKX2HCdMUCqh
bbfW3RFwF13ZPAxzhn+X/g1W83kSzuCurX7z8u6j+uf/Uru5WXtpx44rsBWDB8RB
ygWmD/aX9PCJapKBrZIMNtxChanNzP8uBXleiDCYsJ1YbqflU0TQS+D1EWVqSbIx
LzjaAf8bvpiDcizfW55czA45biIxR4MLCloF4c7CQe8T9mrTskJCmDn5rAdEukco
M8EANXFJgnLbsoEn5KWdK19dt55PdmyEURJ3fP1GKNS4z/cMn/ojcRStPkcUo/t5
vI/9RnmhqMZDFyLjN/82zHBhMwY5xjMOs4UT3tRZcodbmWC7qyN3wfQZ4QCjGw8S
nPy7rrCrn6kYTUfKaekIrXfO6DmoBviZQWDsfpIOYcYmIrYS1na5h1idzUo2barv
i4r78vmJul1fR0JcAsxI8Evjx1IYaZ9mU+5/W68p1kivJIMBmtLinXdCAcW5updq
KxPlQo2SEvN/B0Revj5VIifgxX5G0momzwb9TsiC7Illei1cA+yPX74SRQpTm7L2
w5ddiMUy+ecygDZ3c0Nl7KvU6WB+7n3uDNsWkpfI4tJsH+px151VSX2lGuLcrsx9
WFFjK67LEk7NmFW2yXqhA0BMS1FJRDXODBeN9GS2vmQhlepE4jU0QNWmRvLkaCSk
FS2KIOdekiE+EjyIcRvCq1HxBOWtS9gLn0UYJRWg5agDnZnmBreOeNRQU0FSEifV
j+c3GJe2zivTyjUGf0XEghgtsFC5/D/mYZCQCt9cEcdnDmUtTXO1lLGSJ3qiniOq
w4M2yteS/EDWQl8+QScyUk/kVa4IZ9NrL/ZCQqh7eMnOn9A0KdKWCjnuIH2/d+G/
7b093CGgY17YyQogx/2/328tEN6NQ7YbTkWRv8lRoFli2xUqDFW+fUNg45FBnvqN
46jtfYVY3bY8mh647FCGy8tDvU/4UdOWmpjmNO4hSeqFw58PCdzFTkeoUs3k6lYh
VC3ddUVruvil6eWosyVnNMLSj3d6x3BfxY1wf6ShFFDpf9wglO4PwL4ieSajwU6Y
XnlaCHDxC8tblXzbtRpZI/aNvZ4VvOsKOPYEPlBHRVxCHmCRNYxAwvBNgZTRhjRP
r8Q8vStA+PzGAh38trPERSjCbZ3KmfhO75qSbOUgO4ZTJkzexK/KbVV2OSk/cB8G
OEnTIAAmx2ExS9HG9evDlEUbCH1M1uTTsmgE96IdfDCD0OBHu/k4LeEybr43UtMm
yKZ0qTJ8oNe+dLHxW+9gX4KaYZ8VyI0ajkboWlW4vSR86hGBQaPaxNnkB/Hg7sMt
xkb/m11N+I+DzUx902Wy4K35shvHXFzniPWz0QHncRTp61+FJRQL7oZ12Yu6ACpF
i5QP1eOTPJbAV7Tvz6FWN0NYj5HA/qjB3FqY1Qw59NSajy7aQCrd5yvGd+wmsPhq
xgArFwScVSCHFr1GV/jl7QEbEjF3raWsD9DOmntg4LUMSOTN0TA++oe86SSxpAZO
vfl3F0ijwAHcD9FshFRd3TeNXkOHx28YWnFnHs5s4ClzPpHxKXQltm+/6ZnsoqU8
KQUgOPg/4jnQ2TMPwZtDfVU50PeP7esP00FKEim7wA88Sh1DMADX3Jc1KNsvVxJD
QCgjC711L78qAlTywBIe9gxpZJKUzv14/zS4exJTkt4zj/Hb00oqJ+ec7zo5/oln
tKcXJegsVetUkEg5UhcARcW6+9HL/kIPXaJ7fUEm4M3EJ+PYf9BdlpmvmHGLL82K
vMyLMmjv+EGqba/iYC0e2VLQQrHzkqE87cd7/MmASTjK7kQwKgcWyas7PbC6covT
ZvNJmDtDiyw3d9hkV+uYAIFBn64C7jymjuxabBzWEsrPQIGG23uM5WR+NJ6wB7ZW
nfurpYF5kA+kWYduEoZfiz/fJgtym/rtbcXh1NIc9iEFfdXh0yYkkw3SBznE1ayq
Zi/PbLhlZsV7p6nzug4LsC5yTw456ROcE6VCghXMENegYDZll4JX8aJXZFsrtUa6
f80eujdyqvJZHspj3rFS7mA7cBKmgWH6Z6bkM1pdAS1zCIWSQKM8kfMdt0jnkKqs
K5spf6KlUiKm5VOpt6YI5AkCieFOiszkPNcjex9v77+y35Ny6uMgRKAviHUgMGIF
y969rWCO8gE+o9QTUp8SrUwhKvqh/XszIePJFdSkJlwfr2DTH2pT6FRUaqBiPjh7
Tn3JyQYCQkBb/64dZikQNwr2v1MQuVb+5wvl4xPg/Mhbxcj+CS0O3jyDYBEGCU+8
lbeIy2bfACXoZbrqnZTcNK8texS9Jyw56mJUZ++pdrT9u6/INaMuQ7JfZrLz7wgu
3Z0mBPi97xZQ5E1NqwqS0ZVrfH4F8mhclydX72VQCFHNtZnWEVV+zBUXYUqsq366
bTc4BR6kAhDHJ0wB6ZskTgzgGharUBIXJS7Mok/pq/kmcUR/Jn/4BHvGE0YwvgUD
xVIFppuPJn/CLZNHuA5BXNUNN6/UwtQM3tezY7uUjSx+iJR7qR9AzZia3Yf8VXO8
lp/5cMHGAiTyaBV0exdaBLWUpgez9H2bmGjQt4w3GAH9c5f1Xm+Gw6ZC4fdUXE6M
/C81XB+QRTXQoGf3He3b6MuwhjUkpDbSsZRtZqqbCNHrgr2ryaCz3WMTF8fc09Eu
LmxK9vVPiMKFMp+kXg9y/HqTG51m+v5dU6UosJ77U+UHSBgH5Cu/LHz4rsveIurl
p+objasYatCJvgZXchd1hdtpLEKCDsV7ChgX6QJxFc3CeI5iWJGcVrYHpjhBzLbQ
SdlExXL/Q9bd/lD5AMCndD9wK0TNplNjbI/CqmFGI5XBoAyeCXmhXuwGU/TZfned
9KXp0vkwFJShzCqMIffrbHsAEsAW0rKdEfgIBOEXDahBan8dW5LFGYSqFMET2GV2
ih0ndB3JNZBdjs6JsVxnDI5+SepjD0hKNMsTJ4bfrHfaUJxW24DSHMYCf7v/g5F6
lssb+qU6gDYDtpUZ+iU0O3TQ5G9Y7sV7bRhcb/drfb5cEYLyhoWUX2fOL1iFEtW9
iXZY9O1rk9E1acaI5Y9Dst4Q1EOMYHjK6MvTgg3xCwOyRMXOcIyguOPUigcBNrZZ
bHZjALovxI3c3+eyIYLhWEVxtkmjdreZqeSpc8EG2NdhNg+sxmShjJhR0KGlS7CA
x2HvhAJdPhpxs4ucLrpYUV5m7+trSMp91H+8E7sjrURcFlGi2KzIzGy686dkHiEA
oxGCzGC7/As6+K0wUvhgoC1urVXPQbYyuLcfea2vrEjqTeKNkuQuGhEeEnFcSrss
OFhG/XswHfzRn/9a/1bhOumMR31B5PKbpBZKL3+9VBp5NFdompHHVlP/7CDWfPVE
aKEBjcaVJhmE6vFaQaTScM9v14lQsMtatK6ON9K7+anBCVm1bV9cHjFQnQABXLu3
wIz/oZihO2Fr6tzuAO/dZsmZjKV8yCWo1kNfrPjWIVfbtWl+5m02Of7752wr1RIV
b4LioWke6ri4CJU/YachZTZykc8Pxh91EYkbQ+hZgim2UGxrHvaOYHhxRtwjousH
0ZalxCBfvj6LrxYAoBreSOpbKUULxthKrG0Akw/iydgx/boh967Px/7zcM8o6Gcg
SoRhzM7xD5zbX2rYAAMo1iwLlb5AabqcQFwJF3ii9O9Mat0vqjSRkjuqAVQlWdap
VsEXmFxrdax4FA4ZdjWlssf+BIeynZ2XLHwx5iLrsGW59bBb5j0/8sXoBFzuUu9d
AqOQZukO1hVVkENtQFnr4ZEglO615FIq8teiuwanxHsTGdI+RUK3L7IhRUIypmJ3
vbfQVIvPX6Ep65KKYGpcgfyfl+Yo7auI+x7rS0VNSDf9mM/FIBkfD1uU+iS2BUDm
bjlIJZbmlz38wPTvGnPTNqCrc31SK6EU9iPrtGYf2mVvqd21EBjYmqS3s0ZVqSY4
WyCOQBm6QFuWfQtrd8L7l2TTBOYRxc9N+GLi6iJunowkJRhb1E9gHvqE+tyxu/vd
k/oP5Qkwj6YYR3/Z0ijiqdL/Bwk9QsDCPTGHrSAMsnm+9VhT8773GYaio7zfO4pG
+Y7WrRC+/rU6neFtms9+euk77h+MPSwR7/iXOntZjAHppBr6ItJLOzTGlaE6Yl+A
1tTa+bgLiu4EHzg37LhH7g4Rv1bW/PVv0X09eR2RlKxkkwfeIu5nuD9UO7eACgxx
cVPn2xXRoZoc8ni43m3nhWblUfPi3SAo1HfBiYBnj0XdCRCVeGnb5a8yr7LkUSze
KuaIaYlac9PpUtoGdLMzDkglRZ33m8l+dY7V1Vfpo4th7TcR4bBmOa0JJfVom5Hk
AdjXhdkHJFPeGDsGS4on8zV82QrGQthmTQthWuavRew+iHgI7MQMev8J2w6jmFwg
RlwD3wRXmGwHCCsa+m+5RnaQw5dQoa0dM7w8dVyhx2PJbTpF8flg7of95b0J4eSL
TSCna8B2Du+KOnby8rVq1w6gOeyUeaMi0ZoQnWeaLqEbD4vnIZo1wnmaKIgwEKSa
z7w+wBPjUUfk0CieMYi8mqVCuHKuOVQmU4ZBCqSkWRhY7Abu65DPuYj53J36QLZP
9AveGWwC41E1dOyDYdTYpsIejwWu0mQEQpJPXnzhSE9jQUe9x4mUEtpisb5C477v
Dx18ubYwfB86euvJ+LxAO8PETUwItc4uQHJgDa66HLuwcpGij6PnCPM7wff8QAv6
uGFHuBr/T2Cd6jRSnlKXnyGEwrnOuA/9IxfGtwGWZqapBw1L8PDUZtakK5QBMUX9
ueFjf/7s4pGQ72+a+2z9/zD3Hr3vjXFw3q/AF44IKESlhfGkEaytdb3E/NW2+c93
5tvnJOV51d1dYl+8p6evUOum9EndStcZVzk5pLxcXncI32ZXVz33k0IcE11hhBI0
BdhBiwtmlvlm+FQYsUjHowb+eFf3pQ2C8GLqo/3VprT+iX5mS5ir3PtjsICkNJHK
slJYv3eXpkjC4HNDvK4JgqEXKJQ1mdSEazfDy6ggOYp3ZClUFkEu/zO+5w0txa5e
W41DkgviLuJYHF69kkZKee3NtgdZ3SC5nzBdfM57GfCy0z+763qwoZdYIOMC4gge
tE3lYtnvF0BiiwQrUa4C+zEJVOWnawFZ1CUjTWYUzT9bjNGGc2PW8R8lVTJ8wy2m
VK2gXtwOifJ8VuorvURSI7jiZoG7/y4DYhwNmCWgFgukXFU1Wafu767gDDTK+J1q
m5d8V/8pbIIXk+9NfTocO5dTxIArORQRkkV33m+tw74Na8arGBhHBl79+iZwa/SQ
7gf70r1nxfq8nfSDFVos5B5Og1et5WEPvUbsHQHk1auQe5Y+uMze+sh/K/xKF+Wy
2O/L2zHWjbudDhrAkret2nAhQTUBPm3civ0GNjWPIH8PIaJv3B9dgmwhkGGEp2lQ
pH0sqUm7P9s1krMPvBCHXuqkoW0Rj1TtbHkoxMRmxAUnmAyHvZLUXz9QbDKOFeVW
WrFZKs8TgIFMNeIiM4npwrNcsBnaIJ6c+duaKAEHfy1Uf24RkCmGt/sqUgtEKXEj
gZ7NYHsNOLkKPB01WBDaL7aWvYO47U9UUcIGVDaC8/yX0OK7f65M/2uOC+PUemUx
lepcohqm0b+soQeyvNKjjJNYaCWIaE3fBD+L3a3Pd6e2j8oFHJ9RidHLeRee4m2R
gSvOTSrFlpeW9Ey4pSZclGQIKKaLQgSBqV5jot7AI8l9WKcI8/OTUo4D60tsWbT8
AgO7ma8KnbHexOvAbyzKsOKRT3g/HNG3ZIeOVzaktBIm9GJS52n0mXJJts7fQ7yX
SgoxwO0UCCVaObwrChOKJwNIH+VsYkjs1uGsS8UDCLY3X2c5joL/XOAk9ZtKL4CD
ftSopJCpgOmYMfiRwMbtmnVWeDHnTXlvotmc0HluayR62soQixu8iy/HJ19AI885
sdt/syGXgAtroKD19CyLWZTh8Gt0dpVp3IY+QFc7WCJ1zV/lLZ4jC9RnVYAIDgej
NdA2N4OqpJye7kxYVX3cRIqSE6nDVhEz5zo/wILogurRVRfVqTyo3+Rl4Y4g2WKH
N0PpGUZrRacPzz1qV/k4ExaJLewE+nWtHUjtGURQv/WjLOzOIS3sOjn2KId5361E
aOvKMj5GC4gYEBi7dZulBE6miph9JeEYxHyLGGuEC7n2XntGpqnXvbdqindAfJW1
9ON5ox2C+v49myoF6mBI1n4lhB+okK7PKSCogbll4AapD9iDPtwl3klog6ktCb6W
uOQM5ndcwMsHivFs55BL0+bwAfaQyPeVK5POL7jEmOdOdr7ndxY1sXrEnbBt4F5H
idDbE+twqkEVKBFtj9X8PvKQMBcGyCSQ9c2XAEI182wtg17uVWLElqCeNMXlxseL
PtzmTlQtlCrAUgzlln0i08aXhsOhabCQxcYs6Fa2nKZa82h5tOxwp8Mzabf3qhjr
UnYEQn/tf9v5f6otnA32E9zMyp+SxqY/QlIaYaMkX3PJqvi9Dck1lMdMJb2YmsXk
+UUdpa/b9zFPg1ImI0qNcfcVu8gPzAjEt4j9dOCt5XgL2lOiJ7+sC2QrlZuv4Lhf
4yFyyhBE+TppMtpuF12Vxiu7ejxNC6k5CAnvLa+I3Su8MxUzevQ1nHb3t9j4cWOW
qoyRO67wcsJDz/qks1fRFdu9hIa9cq5bua3EW6sDCZ3/sRWX37haboxPW5vjpFXf
wiJZ6Uz7bnrJEud0r7X/aNzZT5DLovevNFWPbeHpqSLU9u2/4lAO12k6c8ObDkzE
kAGwmItXJ3GGR30X2NYx3rQPRzeYMILGLB+w6OtUtz9q7BeKVPi4rlLuJtHekSU3
2ss77yS0I4/JmT/apkkANDWpueXPzlUwcOg5x9GFMADrm+JQDWw5EkSlHCyc3jvM
fco/cRtdE4pJ7ptcutoxj7gqKexzIny41MkVb/hEgBzVgXRG+EgEjivTVkPLaPpZ
zIJX1BTUrHbA7ozTJ3hA8lHzLbqFBkC6AbpjGFITGcCsnu6vIGo4Adnf0vjRmGLD
CQHMBHIZBmkZDDWDYXh35IF9+nhl6Axfsj1ZSgRXLAbali76HwE4cKjecSrtdngm
tbJ+m8yVXMtqAsjo2TDOiLukVW61WOYBpPgI2UPWxOXIfStHEJacHk5TkGR0yhbY
YmliGq5I81c6b61KhcCEmD5FMZQjCkvpUFKAZtp8g24s2QiQyuV6nOGRSwlS3Hph
DnABbIFdXvub7VZx6+BC1M0ME/2+tnVSI+3KtyVrOQwxgwlKZjy7eL9tSwKKnEYH
uFjPuMSH8058f6L5bBEzJAq42s+ast8iYbO+B1DCVSUdKh3yD/0j+lR87v+p4d/2
FfN2cZNRvDBli6+4Rme/2ohhCWsRw4ZM1hQDCBSpvUkKytJxjorMPBrhLjHYESLX
4cs1K1HtfecdcWPmP8Ht3eo4n/hrLOZYcrbF5JOK31TROpWSrq4dneWyg54Jtbn5
Q0TG48vYoITHu7gwdCH1jNUY4VSJdbx5kDJE+/PL5TzzMHRRlyodPnxyHm7nF95o
ldUNtOM5oZpvLyFLrJoMFx+yIBYlRFfL10twZBOEHfxmGc0D7MiHX/kX5kY4yhe6
6+lMYl30YzMWDiFMWdpjqMJYmv2pFBdxHXvkYjoMZCvkUxtWhoiPCnfbqOoXwL9o
IWmnkfnVi4BGZXwSBz+CHv7EK28SooSsi2selzl1MhHaYMADUlaOiZJsw7BKO4I8
/5AGs32h9N98YxAxnws7haoyBUeC//UtdGo5krQbi6qx371a4EsUvmUBUb+4hhdd
6oBYVgMQga21rudkxx+6EHLMIanf4Nrl8NMe5VFidQ6i/AZQ5hwFMH6puacFzavl
1K87wPq71BwnTkGrBOzzb+vdbh53LXG5J8colYoq6nFdI7e2PdWsWZKjQ5tXsJ9G
YFOCR+w7aGMF82NcpDNxF7nCXq1LzedoIklR/Cp+UjD6jYmspN/QQAjPJxWFDQsA
vS/kEVO4UQoacnNPm+8xyjzmYJiBl69rA4Vyc2CEYwMK0M02UBuRu6DvHcBL5oo/
WjSNC4hyY2x2ok1Xwf2G4Mko8J/vHCRkbVkYPkvtnXDhAJhlKnA9qapByRKvz0dS
iPpXHI2RS+RlD+8Ym6LAUPbKlMEeec4Xkclcz2uG3FMI/sjnR7gWD2o5P9dcbm66
F7E3CW4lsEMWjyza/5roBiiolDnkacPFwBo2USoZVKPHzvc6p+/gGBdgK0QhhGdT
Rp6oUvXfVJRC2VgJt+atO6c6cn0ZWzcJb/zrOU/nX+TnIzV6n2oq1hesgc1BjFA6
lUaZVYxZx/yXu2wji0PiwiFMnGtlL+P0DsIVw09ebuKcRd3RtHK3G04WdOYgNhFN
B1Y92J8lj2oPsrLZ578B6y17dkAo4FzR3XFcmcvP/aO1ogs/JWOrajLpxrHo3Lv7
yD5vuCq8B1Pnu9tUFFxVkvexMii6pdmX8dtMcW3Yp1Y50fWT3YpPezQD92R6nEa8
BDahCodHKPu+Rw2vROs7dXSMYLQs/BIYo1j/tX3ahlYDLoxG/teWYIDmzXFRFvUS
YsieCJk9xthjbTWaL9PBxIBJnP20VRVAU9Xx14uzpmfXePzoNnKS2kR/e6ijHgO5
E+xVI/L33IYf9T55Gb8pbhr0cG5sYHJcsnlVkTf3qeBUmMOaXUJTDmfhtSBSajx9
Wt+L1o/OhvfZ722287o+pv5rZSoY1iwkJs077sAFoLXgxyFCSEyirx0sJ00uVExG
gxiOK0p9KgA2rqlBlFRcWXaAWB4gjMYu8T4JOEfCrSrOsAyqqCzI6Lj6BSeYsKX1
OmPV4LPArQciqWhPjUPYV21NX+YFjdsIwZC4mv39SZLvjCznGInqMD1tBligqQux
CVs3HDq9NfUiEvn4Q7DgenIIJsMWJuP2dmFXvGS4ZePnfeB0w3nS7ZDA34A/Au4b
rtwyi6FdPxECT0jM3qdcdD6dyf8MAadc64USTRK9OhrSsNjl9VNnI0mCtdNz99FK
eDwBvZN7+nbfOR0dJj4nbZAwLwXqNnFC3mmFw/uA6giAmCL9bJJm11iaZGkE+Icu
CoQCImJM5EwwNeJEpPrHKSuVgBN2DzvhPutXWMuaz/qyo4qIHLRyeBYtIqAgXXxa
DytdzB8AgvKiZabowBz4wj6lSr/JTBo/ctYjSmEv7AXWVGDPLoYoaHkNnyhQart3
m3KDepq/nHq7YC8VPIwwQsWUmmLAFMJv78n5rNt4ijY5kEAXiIMPXtM7MQk9N/Zu
15Rx0GhyjxVpGmFOih7R66VBU6+4CpgW9UAHVcPP8ZiR6SxfVv8pnFwyEeitNZPT
Jw2sP9fWOTU+DDGuNKRbKdZqqJ+FgUAN6FkVcmzlmRST/xZ1F5xQ86UUx1YGCwXt
Qt6l1JIW9bzyHQ5LshNfPavDn631VX5fkZNNCrzTkdg2knVwH9uxKFmlGT1D/k1d
l9XxlMVYO+1tDAselrsnfuqqKENEI0tAbg6JFAVv0JMRyULer6csD8Y/Nhwex0Q2
PO2FZJYPPTJHsagdOrQpP0bc0mIdHCvbuaC4Nm+OwhNDFHtVAFMtkIIC3vfM064s
Kg22oGo79BDy9bDMCd0MVOHhAIMp5A1M0NDnrDXNg0BqwDXXEdyQKKuQJgp4IHHH
FUCIV1qeYODHmiRguRBuuSFeUFIkWtVZA9QnQ91hQrUbkT2F8ithTVDUQjalWgWR
yyjeJM8D0SItMd786o3NWgOXE93a4bX76egi7c7fKwHRTv7D/hu1Td9NVI/KhF7b
pVNAgGN7pa+Wi1o6jhCGkvGkwz9miRvYaWM3iujcE4zipes6nmrhB/MZiFkbRh/B
K7mkXphiAqUdbDXR9decjqzrBEJNxmA3q+CPEgqUbMmMrsNu0ZN+8+FhAyCXB/qQ
Kig6aE/QRNz4tPi3vP2+w5d7A0GAPQedRuvUugVnZBytRc0jaSQoUy0YMXHuVWyc
4zwbFsBEFOGWzbX+QOgATgdA0hhki4nTkcsLkLj8f7OCWxIRcSoL6EFW5dFjiP/M
re8A1dGZ9TCcjty5xBNM7F+jUbFTFSwqkQAZRYSCA7snuupgx5/NXQRzw6AUyx83
PJgtVbA0v755aQiVTpwqCJ7laxNlqHuqaABl129A9Ca0s+Z5aG+MV2L+GvQs6sEW
p/Jz1CZkehNnzcu9T+H6YeEKYEnRx6UrJ4Sx3Ru8kAqfoWJItOgo9QqLVlMKBw+Q
XBgb40L0sLgFdfpgijvZ8jPH+VK6gxsNg28nn8aWZvIA+XmcUOqYuvvZuxnUeLll
rBWGaWF7KFZNbQ/XpWik2TTKH9i9SogEc7tDfUrZ1y97iKPPbTVVoJbNKxb0bUuc
TXOB41xFUkFHADHpafIEv5mtUk1Xjf64+iWyUNYJ3ENBZfypSN9lJgwkMwfCMvN4
xfLowvpQH46FtIvOE9QbX+N+NZ7nKRByeASWWb/LIfHzAOsGfANBv/OlOC7kUrPt
8CU35gxpRjOGXmkKR00UbgweU6RvRtbvcbNRsl2y5YcgYqfn+b+KkR7e2lXrBJsg
AoYq543sCAlt1wzgwwzLO3m506S4ywdm+370Luu7jfeeW3Wak8bBGvybFY9L93ip
Me65ioRUbpjfakgi1/2ey0ek4BX+AeliiotfdbtTNiJS2xlgkWMs0QwfAiKwAFAV
GCgnQVnGwfGMQsqEN0LKmLCG24LSPCTLjZjzkzCH071ViXHaV+aBKT+a0sTSNcAB
RjZubjeel5qufF40T31cJKHhDEJWtBvSXkJYftQDT/ttpHd1GlZsSxyVd8GEcm5E
fHHC4gqXOX9LKcnB5R2yMKgbHm/ii8Cu4tgU2oBHSl/gkZeRc/3/jKuz1BQvXrl5
eUUCi9g6k7WYGv9fhaVA5iFACzUyQITnNttCmxlxixwbi4cXGK4kuHbY/91OtypU
d07Bo2SBy1ksM58ssUlC4Oy5qtFJCwI6ag/VvV/xi4UzhArDdykfmX10lgsnA832
GDefPqC9OPoZEDEuW6DHk7QEjOso0Qb8ncFA107v++v2RkmBSjOhbxyFwUcwQP5j
MYlpTw8kdSmyB4fBYEUgPqtLCLDnZ+MnVtMQjivFpg/Ce3kr/yzv+FqotaL8W5IV
Zi5fvWVU2eUb0eh/Zb7lQ0xvzd7gpv70jnVYmfxdQKMMTJ/GMkDcItfvtQOx9adf
1Y1w+QBi4vR5oTjUC3Bk9DmIikD38ULqqppsaW9CXtfEE4A9fOkiUSOjiSSjcB7j
qSLOFNQt8OdVRE/lJwUJ+9VTmvuDdZD0pGAn3eWImUBwsyiTIqql+Yj+q9z2zPxO
qM8KvjxotpOSUsJomkWFKNoGGk8JyybrNweBKyNRyv875VcwEc5YXDsvK/0htJ5t
hSCzZNpPSlkUJLXCP9S/ZSC9hb0vKntVlVPEicEPBUr4rxcINVN/+OJxXyUUJtsA
TPAAaMC5qtyIfGUOe5Tgdg0qM4JhnG1IGhqGMAK9Ano3Sq+I8PXbmwGu2UEL9h3g
Cu48LwVwyO46xrpx6YhfM2PdD0RgCrkC71IIg1jeO/A+nbg4SVXMdcd1VQ8kFF5u
knZEMfh8mGceOEoC0mySn3/vqONyXdVF+HZZAdpk/IIBSIx8Y60d5vn1nFD2ZaVx
uSLP/2csBZwvoT+A8d1fx6VLbNT5iru2b74bZxZmpKRtjJhZyC8hvt4wtZSlQNrZ
BWy95XJmBjq1gQRRT3jGnA7vZojqu6abLbPW93MrNUcpnn3/2opTIa/D9y2ACD1Y
rJSZhg9i8Wc4yOCmN3kyK91VZr1ekMyf4Ey4hGIa/YtwiP1doZ+x9MqX4XCxhtGa
i4Ugcu3KKT5bJbYJuiu1Y0ZQAkCIe3sxm+AWPIQs4qorigC4zBq9bphBBrdqLTpK
G6Dmsx/CKYH89lB7rQzrLSGWSdOHHummiJC5iAB4DJ8uG2O2yfE5Me/Cg/uuC5KJ
3ZXd0p3sYdC8OxlTAL3Y43LgFCDWTrT/cPCi6cdeT0ltWc/72qlNCX6TLkbETWbR
qT0JsFejP8PPrhS5MFSoO/nQzJIbMvr4rHgl/u8OBLcOM55ngoUFmicakNHDJSHR
CLHaqLez8X5koJ8h1viYUr2pl4cja2rMiQnBir1492+pPZkciEdKTFnFHyQMqydv
BYSoOiBrzE3oxsY9XhYQ3zY2HFQIq/I/brRaT0ySyGtjtxmxS+Gmrv3OC3ZUHFMo
jBXUJt40cYFfZaGtFaswr4Qip3JILXqAVMKFQl+HLgfvlDZhA/oG94tlhyhtpF31
uQYT5q6SoSOeU2RjnsCAHRvYI/iPgem5lTfKQmS70gAfRk/ZPQ7BHd7LBEVz/1NQ
EdiRegPsKDhpL6H6IdjNzpcq7iP9oBGqAc23BOyT3Godl6YxHFBWbjHfDii72dKG
+8Wxs0J7yVX3Go58lzj3EKnRZXFb616PviZyjPaOxspablnnxNeGifQAKMcthq1x
fABRQr8YHeMG1JVPNSh2RWK5xLVl99YSYFug4lzCZ5aSptXJhisG2lwK8zegpAe2
UK7loeZbMLKapxDmeXFa5SqMYpFHaCTrIOdzZKX8T/PdGkErg59TmPx4HVyeKDRr
Kz2A6YrxcjfDWoUL3v9V3LvTgjlkxR0xicwdgT7P7QlFPSR0GvfmHsKpRlifIEpB
v8ClEP6Qne7OC9F0zOn2goHLJhyrBfL76AA+BvMJvS7TnDST39bHk6tBYl+5sE6y
MH/M+4rLWN1ZPvn1pYMJ4C/+MA2t1xlJXsbD5knAs9g5QXIarnpPuo1WtluS8Kr1
jDq/Zk1QvFN6a2BorP9LSmlq/dWIe+UvmVHKA/xwqvWOLjA50Gcl+ZNfYx2JdYq9
POnkaG2TtPxKW1TJL26Wi5UTQcfdCpnkXqXhCCq6uGUaELeP9AMc3+ThlHMzyus+
0MZNiaLDdrYZ/4axwUgCp4OeouZNZKI+8bz76Y+HfB5vjTrJDhuTr31NOWUyEtSs
vW+8voNvYkCZIax/weL8i31UtA8xLJo/fzC46OrLHDcqgKqZCaXf7WQYUkWIqg2O
24PaP3nl6jHrksKuSaTy8Ys6A2KTjuh3/PEoGBvXD0UGXyKHroHq5tC5xse5nIog
vdDYpclh7uBMNcU8H0ahp7vgkfdAFwDjjzXQgcO0fDZFjKaRh/H4+UrPh7pyqlS7
6Y4wcs9wiSrOkdNnFr2eyDHidBZQQvVJaTfchCrRJM31ugOhhmLo28wzjujlDMec
I81smkQc3LSn1MDdghle3MGmXN+UJrm3C7LR6ogbC2bnDoGWT+xLYQimvihyUjpU
Jei54WCsvIoNr8mjxPq5NdMgBy4OvKEp67nTBGB4yBwJP5olrcTjs2hNSePI4jHw
68WXCGuMfrA9wSpHGduufSifCw8EB1k7PesCtH8KQI6KaxGNP1IpK1+tjpcP8z1T
fWgv9Q5HEbQjG8Hxll+YhbzXyaochh+FLE+Aecpt+gulez+J1Hl8bM6q8lkpAAWO
jmfYiKmpRMMj+XpIEwlDungETOxxbGA7i0GS3j91rlmm69A14kwyy82YJ5XC0UDz
g5N7K7pvAi2LsOL6pePpCSkarGbL1SBXbRelPp0qkgRvs6kUC047Eo1zwGfGGtha
xAypbDBI2Mqou2rcyVv3u3G2oHdxGHjO8HVzCIwWg6hi61G2IcNjK6LvQXkY8Muy
HWk8GnH1ZJQUOGzC2KlBuul7IlYt5bzuLMNyzJ38if4LOjjYQM757QrgjjNj7noF
QoWqhksRub9+YuQpPPIPflHz5aS3HgobF+6j7Gv+GeRSOz9a2M4zZQdSnGeXj6MZ
5bhLl/KD59lIE2k49wTbx7anyY4j64q23AOMm1R6oYYTVd4HSwIXEBgyFc4IYbk5
+SvRZpMPwvfLsw9UgA1mO3j/LzsaHkJ771/zV8Ao+qjW3axLWdmw6fObG7Al8Kq8
82yCLGB5JwIF/fAmogcfQOJq4Q2CySiA8/PkTDXIAstISlkbvBvS70gsE0JINC96
HhrXPmJDIwoP1Tyi5uIJBYy26H8sj+lIB9TlGlEFfP6A2VxBPs67ajVu590wRqKo
rxkhIU2cUXW9wH2x2l8fay4DLD/NlG5gcE2pOeUc6ri5lh04F5OhpifMyJgLsaFP
J5+rbdiYD8ZAwXr0lQX88QaoMHbqSvHY8F67FcAilSNvEugJpR5/FPF8u+w9bd1C
RbZl9lblMxEu80P/AFoxFrqyC34LOMGxqIlGJB8NP7NoZK/GPRnWFmGCJG6MiDOv
Cjrmt3Asz2/TMMEsPR32TpvJFIBrMi6mA/mtdrbQstYNVaXwufiLTZeFpjOGI7QQ
aEx9qvOsKWw5mTyCPtU53dcU6rDy5QHGyerdpXECiuIfvl1V3XWZ8sWmgB00h6/2
paZL1s9gTWi2NSearEZknkhjlEIPOl2yI82E/hCukbg8LeelE0ozT0MfGxhUG1WL
S6q/G9LLDo2HJUVwJDisKF0AShnYfmlK6yLz9pxAAwT7Wj0wvWb7B2NHja+R0oww
SVk65W10bAGaR+hXkP4wigmE00Luaz8WZhHZZWzGDGbjNqJKvhV2x+pSHWZJtLk7
B4RciwZgPUfyB7188jU/fVepLU8jb+52zr4Fzc8esLT+SUowxsqRkut8L7PxOCq3
gz1cmV54aJqUxKwaLlAeAmCZDwNhXQVMi5Jc9ohWWtpCU1QkUaTGNP5/yatTGz1Q
YKazZZO8x5ELXl/YHwPAKnOsCBvLBt4rKMloYVYuE8B0x/8sRHVJreL9mt8sQiDS
pY35w3fLKMrfk8mi4ns0W/2Bzj/kXZT0cVwb97spkslNTIOt1ZlqMrrplMIcU4Va
lTfQrPkzfrVzYFdzs1s1SI2wp/JBVgnVwIei64NEi47zO2gQDwxl/LEXktCs1v+y
pAXKXdj+tB9dBO6vwKYFwTn0mnqqyaHugf1DK9vnzkk9sTo7nNfe94nVW4M0Sw5S
ZRSheO6VBtr9n659ESD4Ylb0CK4CX4oXcbvWOuz0KqmK/Xa+1fVn+4NkMWzQjecM
iaxhpCN+jCoA41Piw28oTxLqzLV3OUiwKHv/SosoT01qyPP9If9+etq9sFPcp2W5
1jGOHASkzfuXFfN7PwINWgZRxWtq3RTd1GtHFjd10FTQJecGYGCY7gQ16pw/UgXW
CW6ixmjWlV6LAEgNSW7hz5hppCFOxKYOQxq5gxjXSSk5TicZ6yRzsoGUaKps0QmA
kIDVaEvsugl3SULMBS1pNt1G9Rt3PSKXeofpz5d/dohd8HsPEjMUFNY8K6EE4A6W
naJ+vIwbER2nep2cBOuWwJlKCozEtbIyccNVzacWfuzuR60HcDtX3RZWszbR1b2q
Cd8ZDCO7E3zmg5+0b+t9+Nz++drcGdZrnFneI8/ZQYgWcQq3pN27jsnBSSZZkox+
BN0DNPnJVWDIUHtoUjt1ZPL4ZWSNsZV7TFoFQpMmm64hcNwPrDA2kgKel+55nBA2
3KQY1ipGSCofVP27l5rj2WjsfeXub15KXB5Mjd4eSS9ssLPpmoGsvpVCOom3KyhY
MgUQjVTp2y6craWMeUNB9xT6m8FkZLsNbl1SpbLxvNVAN3TbZfsYCe34Y8eydI2X
0tlza8JHFFOYRyOeVLyMHmT6iCHM7ypuGuz06ebxCS7+G4rsdr2eaDp/O4xRgbou
TAQyWeM3c61+DTFc3kLW595qAL77sMSAnrVczV3tWhCYNiene04GuMsGbaxpuyA/
VHmkVw2YDr+6fLOm9VNpmqStgKfkm+HAXZ0L1+aSJdvEUyipqxhKbqLCzplDgCzB
PkFMlydq+YyK4bbW/RsobLLyRYBwQ46RLfpTU0LwK7hARB6Z+q/ls+ZlQJAByH5m
a5veV6JgqLOglDWOUsshI212UKptm86lK4BKblDYBXYctDbBvJakxaW7TFkfbBW1
AQW27mg5bgYi4yFXzt8OSMsIVwqyLDJft+TCwDTzP8FhewdTzP0cIeXaTMbegyz/
xxeKDUaa3Jz6oQ4Vtb0n8QkbM78c9ySfjQlDnrEi6ajWWLgXKQACayMa1ljfRUd9
Juzr/M/nicc2YfFgLznBO0i2VLYxzDoQLYfz5KtUEqSU7BLyaMsRlvr6inuIE3f0
sInYPQjdH6bMVVYyOSxgw+sBB9Y7gHfdVs6BA4LpAAhMSoxmVIkO+eByK4Fy4/S/
H6spRhEcdKI5+CGys9Q/D2SI5SlEn2qNe9YkI9Nn+4fVHT4blGc7gJrAZYSq4hM3
R8DtukL2JEhF4KNLVuDaof2kG6IBCwKkSb0K3cfrePw31EVudoYyzFHyOQkb5kNa
I8SyqIUcaLjMoEMy7fHv7DKYCIJSASr7ABiiO49X+UM9EMrVLu3Uwik7V1GDX3dA
aiyisWIXCzP6ePlwUJWbYWAjPwChUz95qCC0Xacd3q4Z5sZJJAUgkKMPm21PMJw2
MXSfeEBaWmnJ9IVW0QXvS3zUwnUKj5aR42eGskE8G4c0VSgw05fRrvXwUIpSaNOv
iRpy9M2wJYQtDdawh3mifs1W1toyn+O3sX8NhxMgTMPaj+MSSpEGdCC8xeF6iSlq
9nkXszrkHjqMm++QCrbrRZ74x8YA27daePO2xm2FbnHDogfHXqCMX95TXyZI4qdR
3U+B1CvDIaGJNvfzTPpnZ2T8BJ5zvUTmCC4X8Xccq1ebSlR0ENLJ1q8+8F77W1Lh
qaWhojDI9PHJMjsZ4i94Kcxvuxzu8YTp072GbC1ig/zDB3VVVUqi87c3qn9ivNwk
CDUd4Cs0rBm8/P3vdyP1XXq65nfBZHKBIROSpRs67UJBaO2ZDcdaZM2qIK84Zyc+
7FiYlNM60GOUWSrB5smhFwUrTR9mxaKZKJB4Z6XsRX7jPBmddiB8yZN6IW8zZYW8
79CzFNN49ixNxZrAjrh/ohV/z225GZuMg2KrY0uTNfOkAJC/zK5mVGhgdjUKBKg3
mNoZJfrI1W9aSuzUJmqs6iq+xL3uTHKfPAB4wI+7KhhcC1DT4QKB0taRua14/AIx
jMLyocXL+KvrrGYi7xNmIQRLHq4miuFnOSlK7JOn1EsyPSJ7mK31wCrKC2FfMQTv
3Qvzho8YUSkAypzKRznYmVYAuR94m8YHocumMsUxpGE7FHQDEnbGV6g+AhKJb23U
IuA1XyoMvTnq6S7kbe+oSnBuGLlfY6IWT0kZXtdvxuSLAwZzQi6YqP5383A/43WH
d4YOB1i3stFvzDB1a6Khd7X2rMplKXvGaolJrXcL4uj4tZVUs5wn5rrTspkGybYN
iHBz7qoDiRpE1gRDucOKbBknbnolmiXigOgN0MbCn4MPy4MVAcdIswRnKSajkXe8
Xsfg+Mp4MoW/tINwxiBfGFaIzQc0rbbp6CGSQkadFIaKS+0wNwwpxfv/OElBDYDf
yWiwWjz0txC+5qCdQ0UNBvIhuphh1eowG9EZjMahPxJXJFnmiX+yOw0oQ35hBt2L
Cw1rkgz1ywTLGUFKZkqLXe3vH7x+X1xZ3ykFVi1ZV1PagNk8x6c9XHGMdm/2wEyE
wTIPTYGd1rdUp3zNYzwveqPI+bAQeYI0otoUk63/M6X9EBs40y29Xg9eOGPZrpy9
/LHzW7TGvxeduz4ZWTpTTLiYAAMebW7A+lIXrI2SodW51GVB1VhvGQv8UfLNrFof
PgfmQWyGuhFjm3B4M5u9j5uW3PYaF+r0dKuBQGuQTH04gAZMmogrwhKCjiski0Zm
flfjU4ZxXBkpqTEBz3ijxGhBYZP2AVqSS8EkTHdUT1GmmERHCyS2Nfgo8aScLeay
qGtwN4UVo/ChTbeXvOkDqMWDZKBuVfdCUvgU/htpcmzYpV47ClqiNxU6Yr3iEaa/
A07eOuXmOvFfLSdj3d0yeG2qVTQvmkc67iRZztUxkbdbeAPBFUtFSqmDjYYC9REM
hVTDeUzLV55jItbBmovbEG9ITGSXOYQ76eDmGmPY5DM2+vWIhjwxCmGRukMd4fim
Rw8QY8Y4wUJtayD672qVJMFaiWbOCiifGP7mEPY3Zm6SbcUHmrT/wlSwWI8c35aA
eH1UoamuOtZJbeqDTghftrH/1eYzg6FINi4k2ADSqCktrbQk0tLhXCESktdQFq4z
jbpbbNmBnj0+OjMGSzF33MsxTyMJSWwJJfki4Y6krcE5RP+p9PGeeYsjRAhlWkuX
6O8ZcVHTkxQOAtjEBLSiTDBANWao0XocQnuL6rrm1HhgxsRKVWLcAG8IcpKQTcKn
kv6Lpgihlmp97uhEYJuG00YPc+cOb/K0P2684SZDqZgn/sh5dqMPg2rqmZX4Q+zP
QUmMisFItnjl8TEF5E6WIjB1gm0p7ybdUibtQQRa50ic9/0sj2d+Co7ersoHmZw7
Pn3U/POCy5gHQ/FH6LC74m4ZvqYsfAyGhCl6AUVeAo4e603tT4HMLZqdNtD6MqLc
l4l95g2Ii0d8mJhzYGQlPeIO3VICeb5XJbLoLkxgAEchpa6jmDLiicD18RPlQn2R
eB8Y7dwPFGUxOtPtwP2qIT3m7L73wrax5O96qpCt8BzS/JMFZ5It6G5F3OeajR1W
XrGWqTaZcKyaCLg44I8vq3B68aYJKmpPbaXUeMh6MA7yDwKGcukyAvFMcr4i6GM1
45O/Vb1TbIuvCbvzGBmh19oXqge7ReuPZYHXjaKOYAT+mWH2QKCKj2VAAx/OZb3p
QX4BdA1MdElOh4LM7i2S4ryuLOaucKhzKJE2/JUP3w6oRv5sLbma3G63xlKecb2R
9VvR5lcvKlyhVd9+XHTSozrfMc3hjkgg48aGEFQF7uovnxmYB32TWDnpYzHuXH/x
GC/lGG1WYH+2SUwoMDeNZWMzZPhUGOtZ6F2cxRuiRXe9cDQr5oEGkqpuBxwVfcWf
wEmw56TT14RiydTrDJ39r7tLz7vmKwNWY+hNAZEgeFlwoDKhGLNEe8QYEmFKu+TD
N37kkOR+c58sgBjuCEevYjegWFexASXul+Dgq+rcw+bw9v9qmPjJKJSK49RtISsm
JgB2SsR6OQxHQ42P9d8gJMeL9/pay4MNgL/+7+/bdUyx6JE5c8JTs4BHJjq4rL85
WkgqKK+re0dtuJKg+IR/Ky/6LuZv0+oWUNHglCbCELZEcwek/pId1+/XuL/tUm4I
aLYF2U+BkUkRdNmzqY9x1BzjCdMKhlxH3gwuD2iAuqUWItWACt+DCEFtO2vE7at4
VRhJEEFEatfX6HMFYu3X4hYNJq7ICBUUb/9br33EIPH7tkjIFqKvshnpbpDjgN1B
YSdDTT4++I1ePXv7N3WjVik2vdLZTF3DUbI/ptGlOZQ4SbmZGgo3brO8L3c4FZVH
tL9dbaTIYo+ChsI8zXm3rX0UPuxmtnRdX44mtIgd7UVsrx5mzchDlaHZ0HNYvpd1
SkY6LJbL2KdfGl6UGzRP3dZ+sdfXce/uTrSLZ4d7ccLYHn4aCtCzsfkS8ARnOsiN
DX7QVm4w/QsIGOrjejn7CEGwGYIys3Sw3YdDf6jCMDDOpEVov82MeH4dnZO2Qv3O
hFwyKHlLmS0Q/nH/bx8j09nrLYyoGmXYgCMC6KkqvB1IC/pYEt8++UW99GKu3EfK
/3k2S1baii+C0AxhUlBc0qMEsvWdVFcoXiXv+2Zs0E8cFuZ7MkdDJPQl3ERY2P3Y
Rx1jUcb2EhtI9E7jrogE2j6o1kdxoM2fy41I5XhB2KVWhjajj1bJ6fBJcG+Qc5p6
VyIYCoGZKAQitFMWhebpzamQyD7AdT1iwp9aiRcSLnYuCKccxDPJdbnNjyPHJfvq
yib11L7voWRY347/FNgL6RS2cR7qq8iTNmpJZjtKlERbyxNzW9BmqhTObhp5O3C3
v0pERiHGStf8Wu22vRB/SLNf6EExkposrAAi0iIRCVwEt9Sx3Rz+exT1aaj0tw5C
KyRY6M3WP3L2MugbFuG3VhcKkVFDEqtZmVfW2iPGVtSm5N4UG5qc+kqeyy36gxt5
CickC2JUM26rr22KE0O13JD6FE67OnPU1wnbnFEBq5A+lqPHjubVIJ4c6tqDQNwc
WwLCZZgzEYwvw+Xdy4V2h5cB7Usttqk7eMFyo9g3rRwljcMPHZCsBI/LpQEJHZBt
s9ZY/uo2ME/Fs0bJYLjJalQDGdXxowwxvlct02je7RENQL7Tl3JRT2uTC7erp9Zh
Sf4AfsGBZphlpW4qCRB8zhg5eVY91UxgId0Hf/LOCeBmSeLDjfEKb+UtVfbrnocf
wFkYc961MnB07Abv6mHubyuS76JeQ5kypMKIssNeoNg6wWFRK9TtnN+4GQGfb5de
unlRsu/AuVbvq3YgwJz1aiHzAsBf5HBdYOY5HzytbA3dlG1nMgLpwFmBV2L+/x2v
902uWKl0wYvSuehrQUhBZ8czpzX/iRntxypO4sp4y32TzsPH1keFpLx1qOSnT1RU
2Uoi3eat4zdQMfwOW88TjETjxBkGKBPr0r4RAmASBrXyDhpvPqRJgQWQ2jrCHAsU
k7e9x4ShahR9J30LrW3wQ7T0R+EH2FVOMQUHI9p27H453tYcZrzszO8roPvd6JQy
Bs6uHI/3CHwxDdaxIcy2Fng+UenxZr/u/PutZV17kajEzUtG/i4hkgCokZtMMrIz
vZw3IOt5usPrTfHnnRs4GOK+deujsNH/34cg+/puchEdLRhN8gzquqmWZYP15bQo
RA3SBob8ZI1Bryw7hCEEqbzFEiLVyG5i4h8U+f8T60ccMHGGtHnnxeyB5yc8NFiS
vGZ+zZUf1OjNvT/XAxsYHdxOlcqnplK/RRlObbkNlDTa/h4ct9TAje/TtD9OWZFR
Q92oWmBPJ2jc24Bwzw7FDSZouXrZ35OzX/gQbEKcL3BTIo8kEiebm8qHr+SyP81J
jkGzON+CpqDAGFvkopuDS+p40ghzMBt7Dkx44kjrONw6kguzWsFt7E3aYgn+GVpP
1lw3ljwN2J+8ax4lUb3flDSNC+YGJa+ogfh7jJblyCgZPj/erTt1NBUsSflFqA6q
jB50JlMB7HzObRzRa3zE2Bj0DFH5FeddrXp2PNJnR8WTfzb8opdUPosbnq3IZVeA
c8Aao4Q5PPQ9Kj6L6MNXhGDat3rMr0dDIvLY4Yf/Weq+/egXLRl1sAJ3Mcu+LeVF
oNXKwJMkd90f5L2iJbaXTZRrf1t3/0wXRY90yuY+RZltsvBQ921j0jc1PMOTf+43
Ev4vGPmkufyqT02ZeWEmIWr3AGNIalpS/NSZ2U1sdyaN7BGuPXSRRf5vn4DfErfu
Y78HlJz371rBoSLPhr5Se5ESU5WDcxQdY0+BBbLapo9nkeRbIlRnEu4Cd++VF4cS
MuguJG4BYmsNybA49QbXvZU34o7RHyojTHW6XsB3jOQB+7R19b753kqXaCXgXv0y
0b10Dl8t36mMaN0AbV4hheavdOAPdnaSyljVInfgPc5xgUbBNLcu0xz8UQm9spnZ
wuIgFaNIxbnMB3gjd7eEdlXcXVg/nvNPDKN71KnudCoYApvu7nHzTaqjqJRiz4KY
kT6xLFVcIQMhkGNF3cYe3whMPvXOtPKTwP9q+eotHgw2GKYtKHjwJKaTFuaIrgEU
zqk/CfCG8tosUzCyeQSOXxUNWKoN5tJV8VEy/5tSHgKliiH3SV8PBq+hnLVnUDMk
WB1yRhPiI0zRwwoTrMqhruKTuofRqVhLfQ/9ehIOfsChm+yr4Jv/bPR68RW8yfRG
/a1x/oTvXVl8QtoDk8Hcl+TVlU8tNotDr3BqwpX0uYdLJZbkF0T9p+Xa7MLE1r2W
0ikLLkRAIsUWOVR+9bNCab57C6loIi0zAhW45uHXY6xjzF4fOaE6vzC7UOX2OYtC
wkbDpwmXnzTcQ24w8dD3P7gWomLVaTTZgheAtnJMGPeyJP2J2dF4PUyuqDITQQ6y
w18WNlfqRzz0Ic/ZCren9jC8OPc5sa8yTPUrPBfNXVExpqui7ZM5+aZC+50HjL2W
8172lamDUW6UHQUjMEVUr5A9B40KRzC7yRsjXVh28WNJp0TkfHhrtLk3+GFSW6zz
qPtoFNLxXUU6RjZIn635aplWgUg401O5VXp2apOPTw0vpc/mN3XoBXc8+OhjBAOv
9mS7DfKmOudv19ZZetlX//UAtoelLcKon/zufQFSotbgc4ukRo32j416ayKsuCaO
1UT4FAR+0p8JA/IfeVO0A+xZ6iCeIjxvfcQUr6+ufGs7MUf99qLluGVaeKAnexqT
l/iq+xS5jsVcUAXmrJfipeejmVZtEEwyI2JkZy5p5PZBt5lQ5E/8dT1CrTYRFjlV
neQaeQIMtK0hnxdlyRFTE7sHNZut2iatjFzag/wt04DPLkBs4ouZMA8CDs6R59rx
1qxiVOXqFikygBGOJrDAh3M6Mkv9mHTR674DUq6rH/8c3ScRWYSNWdUTIqlUYb4T
ayACOGtYuiY7vz511HmPDbHh0jQqQDUXg3YPr5RBTS2ViUyiCvBjTZ7OeBbEW7rJ
zJ/EiLu9L3m29Knzp5gLsoxLiKvtAwaHABxUsit2SihMrbfXsHvErc1ZI+Zdu6bE
djX1adqNlPWSUDjbTylCKtsjR0gjNulVKATXmo4rDS8ccU399xqpy6/fyWNVAOu+
WktcelsfG+tCceuelDg3IMJaF/X5/iepQDiAAu56XrpcSD+015NbY/3gYydjPWnN
+kVEYi4mCOT2Lb10JDfsehcy690YGmwVttO69ddtYSeR1iH47KHWtMSwW/ICzSsJ
os+Toph2w/nQDw0lTmdU3bMYEm5QCbmqpvA1My9suQTZ6HPpOYDWwLNKd5IL8FSD
Mu8bJARkEJ6UC+PhPA0xpy1XDo0SSDtPmFg5R88Aawgl2YBILxqQIM0IKEledigm
3Jg8i11cl8PB+ri/NoOe01Z27iJp+jbXX+49pSs9EjFciHiZplMws3Vl41wxPz4b
kBwnJAet+Y1AFiIojKJc8x/60lqQrk/CcKCcxpCEBXcisR84dppE5vWhs2XzqyG5
o+1G+aoGeFAWlbhYNS7Hl4SrTsktzTANXDOeqwka2b1WIw8jbAwN/Qq52Q8Q+xAV
MfmGW3l0cnXH6Nhyke508k+R6UlK0hLbdiSb5cwULfkIrSlSxOHfmWrbBO8HS+G7
ob1KVq20B7bYGbXqThEXjdgH5Bd1JoiISlFBFjkGoPHtGFplUd7o6d36WrHNj4Hy
pPTvKCljx2Mej7OwNlyHNfQcg0Cyq5+1z1CObjmB0svonjbZaTLIhu2TYul3alsR
kBn68or5wKB/RMpzgndMHulliP/nI5IW2NzL3DaP2YevaHn5UQ+5QB9lhd8JB3kM
S0FCC0iR+l+msY+B43Buxt4bEri85oZUJX6JLnYtqBszcsA/YF0j6mlp66RPTg0t
qKm/MuyZXDZRqjkunjAOK6aVC22uKyptUK3AYhb89AyTLfkaobHbE4/a5usX9eTi
8ewv3rJwiMPyxyLunoHX9/LaE6A/EwpSgZneOb2fyO0xclQKKwVHzYCg2ZpnKZcL
zPDbAH11LqKJaeCNoQ9BtmxkFDJCNXLEgxXLOM6e+IPf1ToY5dAitM1YLQhCOjp2
StZWgp8W66iZ5iSkF1/jotMerTWRsy9OdMbWM3+PsfchJ1lqK0sN3+QVhh9ES+M0
cbWxwmT+9GnrO3BdTfES/yrKVYKt1+Sr9npd2dQifGGfCwoaS9MrCTip52+LQIPz
oFMzNR7yZnBWjrIhLZnvY8ly+164fxYN2aHgftLDZQqmhSgPtJRXRHe/32+NQsHn
dNF12OTjr8G2ChoSAbM0Er63jwbogw68DI3Hb1a/wpGEgvS/JKU0KKWumw/bQ99M
gvHBJkM2phykTLNEYj1zGVWNF/Yp++Zs/6qHm1yOLP8i7gP/lVWj5kSjcE2G2b+7
6ns0l/GIxf23MReD0rdV3gHX/SscBgjk3T01Q/Ha0NherTXKngKrgHHDlL2a0VsV
sX2aqrYpuKzTCc7A+KNmGfOAVM7Cc7+rCZjOqP5dpvS6D9g4084+oGlpgovNMBl2
QP/Dqi54yPPdfoUnNLMF1XJ6t8o3isEpIf7V6vVRnWiNSdUrM0msqLBzIBVZKNNw
MVIGalrYNeJAHuTsK6Frbk5cL4Oj+REdvqd0XHLvz0TWlEsBwlR2hrXdbNhi8jHY
D1mSrutDsDNTJ0EuFkQuJmlMizagEDtP9TXUFq9vd6+hccsreM/V/HH2Kpoy5nwY
T2oCijHAqEiIN+QTLGrZoKOM5RsfGitzU+QhsCdHb4oFbZwrsxX00/pUP3Pqdzd/
fg3fQ1Xy2+xrc0tuTHdE+lJnpedJsgJmO69z+CFUpi8pRs0muhgB9B2bQeSl1bgs
IlPbre1x9jkAe2+C2N6QL8kL1Cpcgiqehr68slVvEWfafyGZ5ihqWm+fv/LvqZwq
1xQW1FeuxcsDifbLmUQ9ELUalpCB5EIEnlsbIgb0JEQ5CW878SBJyZ7ACYCfZdvw
Ewq/61bSRdIvzvykGIyLgis63v5bwPuRWX/045DO04yM4P1jrwxg91wbOxmX12Az
2mtFN/hd06jeWVQJ6k5Q+4GDTJEZqnMRbLFjPc6kkuTTqaVUUOc9bw6MqIsAaaV/
Q2oL+W/PgYmURUvye4LaAG68jHHMqfvTn28OZjp4tolmiVc8uTyfwihlbjLGWEKY
iwvjYh4yfoyU2mwwgM2w/gkFiAuP0zeLlKjlHOd85H0qRt648beSyqwpz8eLQlcn
PS2zPY+oRX0K4NITBL1r8qGa2y8BytvHQ+GWIz3FfCDIzd0KmIM1wXaSWUAq8hpE
s6yQuIVkD1/JmaEKp53b/IdyiKDgNmEshxxDNd6VwCDODtcnoWS8IAw/hzg2Jjdi
ortkFoa4P3wzrL53B3CS1Jm8ZgkVs0OIWXKis1UxVWzYJuObcV0HrozTVIotziM6
WKGEZK1aKdczXpFFg38zqCDuDRc81PWsneJ4hJ73un4rl3Nee/4UlTg7rbjCuSLS
jujHi6LL3G3BzORGJpgnzYteh9Z9YNd4hu+PcKC3/0i/B2Lt5xNJ/VERwWDkr0RI
1wmcDwIyBvS4vCGfQM0zLhAXloBDLnL+WLz7pg92YVypAE4/plW8qdEsa9aynJPK
RFjMPChNfQgKElU4TNqOqyCL1a5QoCaze+OlVaer4Nr6y6XSJ1aM8U9icCZwHS9J
I/Rt2EwOnhDt+M1DkG6vReUsaSvl7s9+hAmwRbHJjipUENILGrZhFlqbBek4Wjyn
JGdBeD2lV1S0MLN4HLS0xV37PxGGxPGXrLJ/MaUB549VejOt82ftpnfRf5aqBzDE
HqfJubVWg7AYlXYd/9mA5VLtJI1zwxqOD6rQov0RV9++85AoR+YLG/gVOO4Ln9p2
RgT4zwjIn32xnubTm+Q2ZWq8kt1IohrKGBQcHXtOUAnZ+on5K2dx114YFbmJRvhE
SAEiQ1uzNweTE+iXONPgoV7XcXqoCq0Bu+yk9Ij9aRCdIvDOgVj0Y01x44mRiIrT
A/mPfmO916dWmm6eubQJLAGSbEW06EiVeO2BR2XihJ2rMCMY56dh8p4g4Mm/BhiM
s1AkMr73qnsA9+WzMgdqQSacEPW7f97yH6GtOrrc8WdT1Vfm1fIy9YbZ58DqvG7f
uD5X7yIs2fVSwittz3GY29W58RbG3AsOOIofCn4LhRumE/HDhGV8Sz649KkKHzkU
nxrmUEH3uhYSpHjmZlixVoSRKsXCTIbH01iPBqe/2EFcDbsJXho6U+68oc9mA6XR
7arfFR0nN4NqBwfdKsiQcAdO9Po4oQTRANTqKZrc2gB8sj6cHkGeQF2G2927MPbQ
NZ/v8DBH0uTqovKa77/fpVizqiCHYuPXNc4WzaIN19SF2MQN+gL45yNcQDDP9s/E
fTHPWYTXmbuLjHVENfqzwm/GGmw1PkAEBsHKMFmVvkMf94GWldq9or05MPo/9tkd
0Q/xGaM+GcLwEUGmi1VXQf3GAAjWCYZgPmLZcat0AgJUAtIZeU7NzCr1fyThoAwf
qeUoBnIn1YK6V1sf/eOgyf2vR1NZTaolASkkgAJ4ZpLf+0f+bKrDU83Z48w7xGf1
Dey0RlqCR1vSvWMg/GdcpZZPS+e6BIl//MC1CVa6ts0aJYhkAMs/KNk24dvP94/i
Pz45nVAOOhw8j3DKeqPeAPyyMuZ5Ab9kpWpIllRoJ0qDHsSodBttHNeaEh6bVfJy
VIB5epKZKkKjGNpsO1F6yskhVAvJ13928L0yvy3bqjZbkYBwL3OL1L5OaqlDp71Z
X8xUxNJoghn2uXNpH6Z+fRgXjn29Be1giv+5EaP4ZI6r3JfLcZsjQSkN4txkZpyd
hdwyBUdY/Pas+vUgr2q76dOZ8FqENpNj/aQqkqz5mi3L8zh4MvXyMGcij7Nj+Dy6
YRcTNw6xT7EWDAL6IY4niGBDoaGKpyr7KEwFChATAgO7kartX1i16651Jkr4uQ86
jt4PFrgFewYl8ezbaRsZjIsrM37wBttrzQqjfII00EpxWgWvc+hUBaNuv03Nj0yV
0ISYfimZAlTgg4CwWMl18g19PcVswRe6HbBfwHcc+g1X5ljHrr0hGChJUR1po023
S3yseJ9pQN2iF6yb1auT7v1ynUithavwzME1LciPSJNJSBbep27A5c5+d3AN6HyF
H2ik2SjGLaK72Y6KV1dRKDZVje3ffGUorm8eQWXvh0wrwy9+cdfyYAVqrLvIbRV5
TmzfJ7dwP13lRtHd2SIlVpRdBdaEOd2a8t3B1gsqApyWrc2gTnTn7mrsn6U/DWUK
puHpGA+vw7Wkm8R65LnoFBPxVGak4ofVatK/ATsDDtCJbD+7A1mzW8SadLq9dDxf
q8wb5o3JJsSS6ZJN1KnNX2gcxHGf/DrMO/4O1awa575oO/4fNGg0uA2QBJ5OHDTR
MUO6PK4IkymkYGi1xhg6UkYkOg8u1RLx7g62qoTV8WvsUelX6qxZKqbS3BMe6NE5
/YgM7Tu+oQuOg5ph+a9x71ptlhWvmdLTqqFf/ABeKZXsKVY7fsLTG6PMn/v09Ya9
ls0JNrKmIkRONUeULH2D0iOjMBLqctTjvHJcT71G7S7+AU2GloQcckUVxfbCvQZR
IJ5OPyog/LR/W/7zlKnPr8FloVzBAQ8nmUiFA8joon3JlrOlMGRG1Uf7SRUv0T+H
uUAP83wyrKDi1heKdm2Hm7zJvjS+mL03SbUf04d1FhR8a6Q3ARBixTUp72VUlUd5
owdOUgRU9n5p1NvR43XQnF2AqqN4JmTrFSPf47ll46gBo5K/MWLAy0rGsIiBgcJS
ndvK1jMXhFbr3GUt//2yBxdHQ6IcgcI4XcQBJdOOSow66loGB0zfV+pIsbNL7Lz5
9Dv5xkT2u0gTxamQOriScatP1ya3qR4Cwb93w/6to3A7PiJS73mEHhz4qb1hdgvL
rnW6XEmxOUED9t1eQFLP5aCoEFX10bAuX0PSvLX6JUzlKPIF+iCV2fXhY90NKFmi
HMTN4/YIx0kC3Hn3gSBIgROXv6bHLbRFBkaeOdt6LJJgO9CL3liY9EZ9IAlwdgYv
KU90QlVBRLrkygpSpsP+yITEMiY2bQVER9x8bg8fGZaniFx09cgz/C5+J3EZzQ5S
+2r8v0BhU9iv3adSe2RJ2b1eLeyyuYp7yTDR3MgahOAJD5fGh7XzkcI2syzcNcx6
GyDeNqWD5U/XjyBlxlIoOOTrUZ+99HLY7JbW0xBQ/1ZyVx8sXOeH+rP2UWXY90gR
P8wx+ycsyYw/bdRpbYJ9001VInKniEX/Mkin0l96yqgqJL8Nr4MIPkm8ttsyJx17
r9W1PFW9kaYqP8VFqvIgVzv0V7B9m3MOt76DSL3zobNQT9J4BtccEALLWnfIwzL7
BWzVAIecHAyxqdn+roaZwRIX27KGJmxaedO/28rgfV7rEHBHEPmhJM4nBsd3PmZ9
CrCY/d9KjiQ5jlClqcE9Q8iconCKVemAPm3R5yk9w1jhXZwmOapEqmijz/B2X5Cv
hId2mKuhJL7IL1mCbhWIqwSan7rhwC1ccachrBmSWMO5/nOqWKJFNije8GexSv9X
SHoDkHjSq9MuspwrWHGe+sKikSQNKCRP6WeOC6S0sAmypAYceyBYN026R9h7XSym
sT0cOcUbRW3p7UKkcgMBxLBH460tLNJra/IZiHlSRPZsbx3kaix8J4en2F6hAjQE
OtwRVb7MTVxAovfXCuFeyxK9Es9JpSPbfZGz4SdPrQO1Kwz/GudQR+bJ0XjlQEs/
+TVrcsSmHeuHXyE+X/2ccTa4fOONVac3ogtyIXodbml6hmLxygPDUjadPhtJFYMB
7LouqOC2culW/Q1twf4ojmkJeOckR6ILxBkKWAMYnJNSqc73FkacRDnq/AZd6OM1
0FSJs9rm/ZW4u8CT07ux8ji4309thJiuwAduiPQd628zh2KhosArOu1wkpM6R56Z
d31KwacmRoq94Jka/lEHjybzrNuJ4p06TvWzU1aVFLhnt8q6/hZjmKvh6L+450fU
8t7IRghizxNXMZwazHN4qWmDb1St38AP7XCCA8bKb/IiJjRMd/C56DEm+sihVEQN
xPXDoY3BwKk5za7ISknvtO4Qxn9YYJsOn/hehGe6JDvuI61vP+n57pRpumi9xMGW
GclARYUIj37Q5Z/9rxIrCMx2aVXzadoqda0CD7ceg8WFEow8pz2KzKtRDSxLNqPO
CiR/S5/lCOxvFvXkoQPwKsxnCCQORHiEgM9yKoZwId1aB/33Jfb2mgPswXfboMMh
JQu8lIxEgCZ7YEBPO78rYF7x4qr5o8t18wWghEVrQOGCIV9qRCQakBgI0nRnu3W6
8WDTqeC9Obe+Fubjjr8QNI9FEpBUlK1TDoyRGSeTn8/Qr+HvcHahP2c71/q0x1lM
5MiThjm4KlYK7DSbtsRGFkLrAtPCN2J/oCez5D+jZzrGIL0d9nGrbi/A6o0woRrs
3XOqEYp2LQtgmJfuE6ynBA9pe2B+sTucpZBPAKpkjNKJsjS5QyCrnIaL41+QtqBX
uUs87T2gRrdtSu1yqHk6KdPozQqAev3PKZ5vvYrQcfcrDi/G7qYJgsVt7ka/yyvi
VpES1k+f5ZOGF79CKJQ5+X1qdNcuGA9bz/T4S/eRTJi9l3m07dCanNPlHwGsjFSp
UoLwzLwurs/iW/Pn4QAeMjADHRwnnPTOM00pAmWnYLsHWjZZ8UUg5WiOOE/E4Rgy
RbOjpkXC8chJsTG6MmAFsRHlae7ge4SmIQ8iVEfjsD8Pd5EOL59prGuxRDEWAWDO
C62en3Xo7Hn9vY6pwBCZClkynEufC7EaR+9Fjizzvt8LrB4iXhPmGH1rnu19Q1z+
nPw87HabN5uYOeQwEV7mXc8sNYIhGNTkCql2btJNsy5Cm81pI/yVCoiafOy8RcSj
BXHqFvRhGfkCsIigXKjIbF+hGOFpwp2hwKLPeEHwV0EtvSlgXZ6svaNqEocAz+0t
rLbIwawkSmFJzGVp9Y+Lqfw5/kMxdkzeG4wAZZNObYBqzq86+FUnQuK0Zh/AkUn0
3NqMoZu7nBaDlA7tFQC31RIZPnCU8L+sKkr42vyJdQv2IrD6o/GaSJvigaQX3txy
5dlqisE7E2O86y5t+c+g2HJJJrngLI8k+v7jBe0H7Pd71zq0iw13ti5NmAW4rG5w
lqJDJtRaGuxXY2EzCZNQoycOkh7iNETOVxY0AtCvUPBAiEhdtBmeUn8fReiwkOP0
x5Q6HLwvy9vvXaFMkT92Br9Vs36SDjBXt84fvbvC0g3TYBAnItrc1pu2b4XduOBO
haa2emiIm4P2Lbe+iyl+KpLbMV+F5yJT+cT5Cyc/PoNQZm3W7teVuOfa48RfNCso
GNjJzi6xphEbGoPHcclWikZ9utm8dnWfaExuUA5P6SK6tDiyEK1Veb7PtOSPp+Zd
mHaBuh2SkKGinmDJcARqxdvdF/YOvVZf4+lVtpbqnkha7rJ3QksbO2zk3yqUra3l
cOEqggFmaGughlT06FA/BqmS96J9X0vCzxA8eXFOV9wEf931NLbztM1ikakXwDpw
UHG5jjmX66K5aiYnQOZ8/aWLIfffcJIQhP5H9UU0j52tREVoPDxYVLzKe/6qodKD
YFgX5pfA//lCTNNTu6c+QriDWQzF8LM1+vDl5Eu0Fmm87b/padEtjQZK8jfZQ60K
desuM86PVe0hYEt7jz34uX8Z+dG737tcSMEh8doArRqAcyiiGYy25diogyN4vhUC
UaJaSxqxNvrFBy2csmirkwXIz+eaOtpI/zlLcfhPLlsXnPXtEudCobrP9oy5q/YV
atXu5VlHaV6ac/8vUdcyyqEMEAmuntAcg7OZiP1AI/iplECP7jSBjjSLgdkUjQL8
BbcaRppaguHDskkk+vAachIghRDDgx9rcq+3Z4D06W3pd8Ml4Ih4H5bQWodL/pKl
yXk6FuKaqJodjQAOMrsEFumThV9v0CJOyjsgzz+EB7KCUDjTjHFvCW9vhjlwLdYe
IvYpzih6Y3rP3nQzisx3DJ7hbst4jf2IeUFx45QMMmTm1ybFu3pLa6wahlBZykEC
jec2pfuItFL95J/ysX9KEtZ858f415928uylpY7u9fiiIJOzcL/E5syJ+4UvqAdQ
07zfu71VHGfNZfRSvXE/dHQQdzQYB5GH4DxGGfqDJqnaL5miZbrhHWE8JYgRJRuu
xRZP85QmX4e00KcL540ATaA+h4Qk9WV71P1bxqAgzbgWNBM+8bB4fN5Oa5IW8rdz
QKAJkLRxCBIXLF3leSQXh/lYLCvTX147+saXqHHrib+cugGAoDnR7mNhKt3V3stu
UAXVnNo9s3kvuXUYr0yWmaTUJ/wTyBOyw74AgTv0Pt7l0holf0lOwHbgpoqDCVKb
+Ml1SyXZ1x1hFuyySlZas340GTb/ok595pJQL7xcqXGqVrB5lfVq465Fh849fNaC
dIbxX7NZNsdzI4gB7pqJ1xap3NwrZ2TIEfcFUmRhlIrtW88ZKQqPgSeu262TkIYW
gNR+KIp6XP7sehfxJhSPhRzyyFsp4lOstGqe5iQlT9wJWs5ovSrVSpPztr0krLHA
ZSN5PStuSml3G0GmQpQB3aqw23mJepIuShNZ11cHLKYyDReSNzNK6+oZEGj6qI/2
KbUPq13eTm93zrcTIbKR7dGjCy0uCKp37QfJApLoxwfAFj6prB6ZjqDdeObQyNVE
QiFGeP28V8N8VSgfEqGMKHQE4+L2Z1Km/tL+I0AB3VDHnIDFynoMvky6n4AMNjf9
F/TKAHZrr0psQKy+2cE9CLD3keskDxU8EuknlDd6ofYq7slfFHpipT0+dGabKo84
GgC2fXKxJZ0KKAdoSGYdgys1Galt0ljWkty+QGNHDzZpJOVZIdssDdvat59dqEsA
6NmmRiBU7+FoHB03RWRI5Y4VyZwyCvjL3ykcw04Fkt0w7KnUArAaF06ek1hg+jlQ
clpW1qBdwysxFAxPxjucaD0LfAlgbYAzHPzoVElMujHcEzgAQgmD0DF0DSVPHQm/
CD9bCju8vHJMRFe5j3QDsgP1mPVwYTDz9AC8bjihA5+QCTpBUA/zqQXgZMvc0k1b
4+r/5zFt4eDkXXsIoPEJ/AuyuxRWrYfdgLfUz1IZx64NNmDGr1WtdDcrWMcymUAZ
tTDofftetRG2Kc1EctmcephJEAkxQSWiG+stkeiIO6s7vLg1Mhj8Ya35GjNpT5q5
YTo1aJ859O+qFhukwCmBr8CNQ1o2UAix+DY3ZR+gUCsho4he/rhHDBWRAjoaiX25
fnxYwgV+F5J+J1T4TRUlklD1hJ/H0BvKMYwJYkYHmm+3s+Z08ZauXl819Anl2WHp
yoGsjsFp4CYXlqExQfTBi7/0rp4+fM9WIRm97Z2EA21wiv8F70ghAo1Q0EcAKexA
DRU8nObe8c23ofgk3RY4/oJQF0sRLJ7wy+STuQ7NXWjuZcwgbHIiDrcuBdqYKzzm
OBa3yxBmEMnM9ZmIg+V83V0p4MPxYaVZTqevO9SMMjYZt1pQdejpcwrtdE2ZNbcZ
PKlQDJaYgX51cUGxE9vzkPwylS9u/0iRYh57tsq4wRTopeosm6ys9L4bjCnP1Cf3
zJyJYY9GwiAuALcC2NysL7xWJvf8Sjnt+4q1RpszOwSEG3aNwFjBWRLoGozBJ6BB
MkFkVRdQodB6wAZmPwTUj+m00GczeVvGn0aRAPUgr+bzjCRD4hZ5dj77IqgJhWRx
LoBN24nb4Q5TqGIbL4yE7yqnHru8ErdhVzrgOo1dLpUFCWEBlvcSXErnbPNJNOnx
c9kDka2zoKgfcR7wV7Q+CdcRl4Ln6wX4KyvG41uqm5ups5ehEis1Kf3VpAjJaPBV
V+BvbVXgfZGWJ9iMf48ERHviX48JsvilPeQGumzrIr/h6+gzVTVXF8K4L6vYdh2j
K7buvFt+1FACkalBNFLKJLbAoUnEouW74+SGTcdBEHtgecBKhP38ihTFB+J4UnEs
w6aTjoHVoOqtI9lTBz3V/6dXknOft/oxuqd2V6bZQsVj8H2CflaxueP4fkrUWj3P
pWgP1mvQbHy5ygTZ4iZg561k5yTaXU2wUj5opeITt/DaG+2aW/3it3bN+inptc+X
0xC83dxTxawB2+qCvt0ZqEXvI9Q0JTrAdWMf0pcG+D/YaNzHb3gY7lAv0c0We8SQ
xVUW94Ff5Y1RF0yQPu7ipN8GMJRTUxBkcLrGwMc4TiMUCfx8tNjdIaair6HQPxSd
IYINFJnkZuFGw+MszgKyhC94A9XrQ8iDoHKcSepppk1U98PvdkXHnq181Ro0s3zM
ChtzGZTsb421G22S9H2vYq/69uWvd0L2xA5/+PtVeUVV0EkAK8esh5RxtW0Zr56N
D3kra4e5A0UDXODnTKEBlUxvqTN1dLaxo2Bx+GJUduxlQdmdPSjkDzdar4OuykWI
3/P4yMkPcYgvK9TASW/QzQL/Yc/mgtKktwf6AhVdZ4NVQTsd+5mY4CsDijze6OuJ
nsJQCF3Xy2QHAjxSE+VpCV6TNVzoiwgNM79caV8kpJYYokJQA7oTzXIg8GafUiFW
XZx+f7cVJEBfD1F0ltKCshVbZqX58DeOT2i6e0uWWzyNFgBQloIn6R3VwmxrFHoK
wiKPMfNIgCgMCE0SzN3MkktJi7VbdOI22datsKje0WjpsCn9E1xVoSu1e8ncM3hu
12QlS5LKsyaz2tUKk12pfYrzOKNBcOUcWjZyjgSzebaRHsNS982ZQw3DnFfDUB9Z
JxRSA9fhHCrDC82Wql30nb609ezywKYwwP/FEFJqF9K5wCpkS46Uprv+1Jbb40MC
uSKVsNJ2kKK2tfQj2Ds222dgO7aVeMpvTIoTA2oxh/eKmMjmRxy5UF5Cyro/K5Vf
cJ0Zw67CUv1ZWoNoZXKf47HpDY3/wakrKgZ0sGgvu8dSNZvGPy+dF4e0SvWlsmZ7
zDA3knLx3Z67YH53Y26zFyIRxod0W672CF7L5jXguhAtwAqf/IVM4pzFD+wT0qvU
+5cKX0QkwLO8dfSS5EqDGdigxFIkTsK1+i016Sn7Yf2xsGGdvLKgqmBJ8l4xsquA
96EFG7zsN0iIFXKJ6qTqIpRQjNkpDb/S4anCHtLTiTPuKHut6tPDUrCa40k5ss2S
uNDZ1z20yibDYBrqTyhaix2nnqSvaseCAf5nA03UcBkDwFMhIvmZ105PEMSW6ddm
bPi/KKE7v4F5TIwK5wQ8LxidkLIqAzao+EDTTgS2tSXWpvM+swVBnrNyn6FodP8X
JhZDs7jGFCuUiTgT+N2TjX5sMB1PyyYi7pNbp363EMqVlxBbRe2glXqzpkEFzcpk
eWhqQ72Nj8g/ziLhEsfhyknTzP4f42XriRAvj3ozdSJMKRDgHfQ3ZOF1thvwdb4e
QhBiKm424hhwUJ4lCdeETYDTz5P83+93/RCimgF4+NpELZFaVCbfT5LZmBuJJ6Tr
+UVZQ9rRTEFY9oFau8DNLdnccFtQlQlV+kbYgLaI30ooXWOf+WCkUPGBTu1wmSuN
oPbet0/HLqhkKWUXSh0NDtDczan6mWhTsLnW5Mn8z0+aT/3lWMgWEL9htJhMQl19
f/sXsQRQYlD/cZbyYwJJmiNV67bh0akypw+J8Ku6v4iKc4h48dLTvobubBdELaJp
PWZh7KijtWYZeiOwrtRJdA1q3qruaHoJdBIPU3GtKK24tJXqsy6a6LmuvXUWv5N8
XuAhjvxJ0ab8KXAZMX0Z0f67pmr0TDFxb5ch9wd1WEJHyMMcK8NH6I7IR2+XDrrO
i5iOp+P7mMrWkeLABTSSbRcyC6y3aJUkQwJp+mcen2rKGh448/ZWfVNA7MLSdr9c
RKbSIJiMAbRKC5Em1Bum682j/Vup2VbccJFCyuGQuXNJWA1fTaj2kNviWymFO8zh
QQx2btDDXS0P46fKOhpb1DJcSWEnkPo6wT5RpxYkhlhSJVHo/HvNnCNIRXBY+3PD
JemvTrYxUlLDnP1iyxEA0Rhb4q6YfTwDjiHz31zP2jabTcYkza/gWTW/UkjEYWP+
o9Z3cZm6wGWcJ976pAoXYhD9WK66HvruiTf3Kq7V2q3jTmhtMz7TLZaBxI6jc35o
psmm/Rm6QyJF0A5DEj9x4yMw0MYsLEJSSLublHEML1qmQgMFS69z2IjjS09rEAdJ
ySN1+Q33x+ibkfxbktw1XzJjLin3RQJj9i2A4/DJgJ4rbap7mtL23esAhUgu1Fz9
dJJ9ZHvMGJhfFjxT2KslSWzOvFQc99/OgMavCQZzPlqDsDF2rOdj8gLBKuSVRjFX
pVBGWIZ8xe0esp4ylkVnUvo/7B9HctM2X9GglCaRxmnl5yXtr7Og5dkTL1dF5JQ0
ADyeLXl6Lq2zZv0BxAiRpcZgOo6VK79H9AUZceIH9+lZIpBFFyU3kO9K+UX9156F
FamlJcW4XrgPySzUnCAQunAPLkzaltj2NuBHUvuCZvv6cS9m8lGkDC9UKkCU/tgR
ft3+xF8fIpSIPqXo5uWeCC1n/fpa8DDiGbvHavKf/jnP/BRaG1suf78KarbQcsht
S0Jx/FZ8KPb4z6zqTrJCpaAgo6f2doIreJIDYHyI+EuuDMFTgZ1iYjRXi4GVYt4n
SK/W5SBSS+oVdPAjvgEm4xaou0C3+h9yxiMtFT+sG8fOYRa50QoACSj5LsAill/L
0ymZx6Ihml04Ql8ltJMTGuTCd6gVhfkkTaW8zxNOl/MBAEQJ6kyEFo2/NvOIZpaf
Aygw/Ac+ibQOL5Jr+NYX2mS73kN0YwKY2JMSqDafO4+rqgI4c/zN6x24T1uz/W1l
pfS74ftZ5jIDJRe3j6XkdD6VJjK7grM5PFkm7h4UhDU4VddFGM3LB37mm+vIp+4c
hzjWxODVCZZHdmiwczx9dCI/Gu0CbMjdVvo0gsEkZKc90v1k/h36N9qfGZYKW0M/
IlV04zt0Y2jwniulhqV5CkbHB1gcqY7V8T5wxewkOu2NElCbRrNRH48tS4EEaXuM
aTVFnh+EQEnPm9MlAhtrXbFO9Wbe4suVj+U09qrcZ0ZWzncURycjqxikKon6i97c
gCJjMFIv6DIn7JvuCYa/VKIU8PSwbAcaRcIqjdb39z+Ca+1KVoVJJZZ7nJIZ11nH
bhAww688egkvrZqTC9VpUjvJgY1+iDlTYUigf9EVKbF9oL7iWqgSv1Hv874r863P
3dWi8Vxnh8D2nkxxpeXverhJPcYF0f7lIVDGEJoLW98hcqkh7WKxg41Pb+0q3tEZ
ru5KNm10MMEa6PYQ4uU3+VQViV3k2AL6jq+WvBREugURXuiRZQ0Lx9Pvg/Pg0FxV
eqgXg59yU7vLIH9tQnBzjk16sswWtthtHBe71GH2QzFiH91+pIRngujOXC8FG8uS
SIocwQ49M8J+6so8TfSIDXo6+Y45gL3RYiHylWrQyLL/Dbt1dYlQBFEAzI5G0aEu
8kcmZp8Fu3R+Ccan6wlb2lOcNvWIsqUxqU3qTOgvz98L6zZz/HnCw4S8QyWoQGyy
kpFukoYZuSs7jvUtP/5NmUIBvEhFrCqzVHUMbFNpTGxnfjPIhNwtQkmfm/Buq4gN
v+FsFTpQCGk5esxLUAjOZnmneJIBCyGzxxD6gvyuXWkqoKHRFNsy7hw9uxV32jaF
GCAq4FCML/IFxH4JZZbblv5eJ4r+qSjkYKKbHqv2orbQ6XNG9zEW0OCsM+uBUWLs
o8Nx7MDujVn60E/BBdvxgkpJ68zD10gGa0dGSNANNPG8q3lVfroyxCg8d78FrtkC
txhoMo+9W8BAiIXCqLFthIQi/ODx9+PKvmmt53otZyM2rj1q4SSsnGmSOYR6vcua
tbDXcq/P59a4NWII6vpaAiwDwtQXz6sQ6iZSnJNES688prBdSBDnPDaxo7ZSUYKN
LwP055kIjGoCz7bDg1niXSZLxzSMFSKS4BVKni+Dpk6JE01kcSZOE8d6wrX/SVdu
A5ai1Hsb66W9CXS8a4a3Pp5fevhcEBRrtSejVNHfGdFTjXjQ6FnOwW3NJ91A/gHk
xBLloVeHYsF6t4XyabzPMufGYGRBlbDlpYNIxJ7QR7DGENpBgivxWbYGk0V+y1r4
7T0Vw2LmzRkm/GOfS2LqbqVcWa7NjFsXSPhUqlKfLwsAvT/FHvjsBErYbsNs17Rh
fAmOlHFyM4KI+98tGjsGzC029EFj99imRd3TQhjOl2gmb3/dM3AVJTePZNjdD9f+
HaPkf8OySLvFQMHCKuHDTAkHYANmzQl3fLy9RcHlPBINFdsHNOpBtlr2rNNWc3Ab
h0W//IxIyi3zjJgudMlAjp80qOdWkDSEU0ZKq9pghuwTIZZvGKNZOJCFMtKoA0pz
x4H7XeKVlkha+dnPFXA8OBffqBAcWDJ8+YCyls5VTK1BodtmxANX7MTXZFploG11
auLslG7K2UOx9TS/I7DIfwOy0QmnTLdYSzlqrS1uJUMQ/lBoZamKivWPfkuuZUEi
mViS8ChaUHWlkxSAg4aQPN68akNdCZHVRL9DLcGBoSnXH2sIRIivzHjiznAlzJty
zG1vlQjQD6kjBfJnZccFTeJzOvpjJJpAAhxkBSX0jxqNMlvKa4bYV6J0obOXKQb+
csaZYW5xESth+uB+fVKZrHaWHfDaNI9DZwIByVtgQuCBp0kxnfZVaSyvZPYEpbTN
OibFpPZ4ka3g4prQFqEIYr6KUzJk2zqLnS9acHNG7oWe1C4zLxlIW8xGeM7Q/m1p
zt+abJmU35AXyQGQCR+Mvm0kc67nzfXkOKR+Be3qqUsyUQawNMTj3ld6aPeyXlFR
jKW0MvOZ5FGYfs4zJAyzAA2LVtldkrbvdRvjbjF1VkeKgwLSW2coPKIAWIGM+aPJ
uYpxdeGQ7UR2N+uikTm+yUHFFWqA/oxz77JjrGBdEVvpLaWJGXaWWkr2R6KpGie2
3U7UJB4xUvhYucln5kgz2bHCCYVfJeRYOiUgaMUyx3c1zdI2mj9SD4t5DtOvhgEq
sN8aoVFGCxHOaPAjsY0LAnOGH6fuQCd8wxYCp9Y7jd+0lSrjyhiMgwnsixFqNzuV
vig9V3gAQp3yeZK60lmvm5jNUGHZ92Rt+oFG3/4639Iqqi8nFNOwzt4UNrLS8rIp
kIM6O2nEoU28oHQ7hAQR3s2U+HbNeICxfDfIh0k4AI9sblnjeQvwb4CbbVLPcpu7
tM2iTEOACPRBSFCppeQFnN1CH0b8ttlsCVwIBQf7hpk1tSsQz8G42Ay4zLNt6G6M
HCdpwg6YzacwAkZ+r04KMepeIpJ1qhuchl1IYiplGZ6RnDOFCLSbgU/zvgT8AT2p
A9Knc0PdPDbIqS0vXO+gTCbgFS8CeBNdSO/besHz7NZhFSq5F6NIwZlnpPqpeiub
Qe8Qh1uzwGez5kIElN2dEwBQWjcbfpYS5zIt/WG8t6Bhu03mB50dHDIBbGhe1yUW
wTdbgUl4PqmxIX5psXpIVA3SUW9GvNMX2AkViZXaz7V+/6UalEBAjxl9IpML5xR4
sjs7yOi6CX2i+3CgPPaCFlle0isie1a9ORoRrW69zPY2w9ZZFlxdqM8qG+7SkYJ0
wvdpA+Cc2396wnpDsg4eAuAJbnskK8HJzsuWAN9P+23Gybqo57dAZoFLhnafi6wH
zX/nbJALiWIFNXg5C/XfemXyMCbQ2EzzAdvScYJ+f/ebKV7oLWuS4CKJRoZKcA3d
CLRLCXXs6oDw/edUmcP5codlW8YvjYVRVmjSFtc9YJuP4Y5qQNClUnCmx4uouXK1
PwxGYfsB93/tNrdky7tJ6TWrHKZQQUya6nwYUWpfYW0g4v4HJ2OyKUKT2z9ouQ31
KSPjxvrufENI4HDvJcxrU+PqJOVXsDL+OBogR8e3KucBBTTsrd4lNx4TiJeVa0Ll
j/AzlabpgeUYM9heJNCQVs21vK3uzLFcff8Uyihj3Oc77gafRIZdj2Obth+6wYoT
mat/IXZQk4xezyWjxYXIZQRBpjuWFwzNpKjVaMKo3tuQPIjfoaOl/bdru1oPMdpS
gTbryYhLXKnzx4F++sdr7dWJOULtgBDJckH0bGLNOtaJ7W78n/t0p1r9INlRm+mk
LhRN9w7DS3hFRSe2Dleh5o+wWjXUmVQDbZjQ+B85064CflcoSOOAIcISdYuUUBOh
H26kXEAH62AW/J5KkZRjYQWqSWTUw3O7Ol/bfwcvw7SjpfvaXk9S+dFhMpNNJKRJ
7pqb3LO8mKcJXeb2QqTiz1EEC1t2KTye+Fp2mM7UBjv862euEmdOuPQE6YaP3jFm
iS9kBkqtX0zp3sGrgxoCeS2nP/lXrBR1J5JlDF20PM/cogLHrqKiWihvXfpzF14f
RE4WvxjzbGOlqGGAXHVxRTYuPVkhdz3k22Oz03veIyF03dq9Nqf8BDCwr/azKUwc
p2GutYll6lmBPVg++x3xnEoQnbqyFg/hiQmQzncu4eKcvl0qKyz7ukwmu48jCNrU
uZR5refzTJ412DR6kF2Az7mQZYMZLbL4FYwxwrdMik94G6hU+0+uJfz6DABxCIKc
w/6/XRsMx34mDsN/gAbQ9IziwmcxKWhGl8D85bqai31DVJLT7Zuc/VVgnFglITRK
7XGVPAP3CAcrlgB5RhfuvHQ4I3AgSmxjd+Ao6kQxRtzHNLb1qyRMWHizJRmNI0lc
dXRq9TLRhC8r6GSSztMMe23sH4NHKKYr+ZaQWzouDR1rIA1JM4aayLwkue9NJTyd
xOkVxXDqVH/FOD9yCJlWk1vIodrxW9QSVK8xPiZ+62GmZAj6XQLsK3/EGqgFztRt
GIUsLritORtuqv2sMoUlI5YLlH24l46fQzLg23rZZPYvV4OXdUWq4rl7VAHnbyKS
MAxA8CG1TW2EbIFinhJmihYbt5Fk3JG6cqKds+nwRBrMgaAnYEz68LBSnJdKdosc
7AOYmHdQFVhezdaD+fnkj0yPbrOcGxlYevCsK7kPURim3YKh235Kp0xWO3/yIYFZ
hQlMHqQI2B2rzC5lVPJWFUCHeYwwsmoHIaKNUK0AJyHyAgiIYQxUAypyV2wmJ9tK
Vo1rSIvchGRfwDSjxhUiCf8+S/S3G66m4JQRv9kpRpHeR7RFWAtgFyZViMg1fDBg
9wv6SOJm3H5F9DU+dz6w7SmWe9o+sAJqdox6czmFrT2tTUyc9EBcxUquEp3Hn86n
KfEzXr0FKsaGwcsGaCIq0E7TSbuMroXqBYngtio7qQAIWbBh+PKQZyrJJpTSu6+S
bSMk/sk6otT26XSVlq1zwj7Udkg+1p/DDdR3KDM7jYjhw8NJRlaRc8dqFALJmGqE
xr88xi9Tphkr3k4RLH+H6visj8TJnWY2trET79+8BEBp5gONrAJZFkUEFI2MxF3Z
Rm8n5AJkdZLz10dnx7dam5mJ0mKjlH977gLYBy33/w63AcQsJz+haOD5yUlpqoIS
y6i2b39glQFpoL5Egaf7wKV1E6pdN5gvtAqca+Q7jUy++gbyNWtVxUL/VzzGIbWT
YzjxC6dm3577MXIkwwOwc+Ns8ZCjZ6z+gxodVKeuSt6+MW776FxbqhrmmxnKJHrE
GFhKJ5SxHf6Z7ufsxSUztGlzz6TwOjflRC2PJlhpybSwnUTld20IUtRE7G7COlcw
Q/UYLxu8MLYEBBHPCNiHzJjxIFs0A4bHNGRP7MEOEnB4/BI8I3eDidTjq5BzmdxK
ULUkIuIcOm8o4qJdPxF3z2qTxfaUsmtYNTxzDtyv9YhvOGHmYuJ391RTC3laqRp0
80UmVsfDbhwDsVLkyf5tksnxNx/HeDB/UzdklSqAcm4Z+m85cRyVt8qmPnlTOKCh
jjHPGVMvoqZQcyzpZ565+U3zOVuPtka7yu0SM/Af38gStz966q8AOW7T6aaCDZrG
8m/MABXeC7YvBXemrpzoRgDzJtWcNefKF6qt8NCe+IfE5q85JvWdUqWKgGPTJBua
1QLZ6XLQ8IN8WR2ZFgTB+0oMW3SoupdfoChb3Qy02kdNh7P4HSrUfv96PTGzqTeH
HVUa98X2bZ0/wogs4GIkjJlCYRJcPY76gOm0hwwP/3up7MvVLr4NMbzgzG3Vyn7N
pYK6H57ADfzu/OCvrDwDztQEBtZphkZJYn20CBc+xznmR6zQmmZE65teRWcWBnBI
TopSrTv/CCKHk3esl7zk9U0Du/4+Mf+n01Wh0PjNsjJN4Q9MdaoaK6qrjS4SXgSD
T9I4QihqE+dSRb1DZpeHVEC1jSjYeXCs/ghd9ZES/j4h1tHNhI4v2PYRQln2OHgx
mnRzmomfgmwefamw+OL4gnVSnp9ca0XFfufL8n6aLtqcIqqbjbwOh35IfelycESQ
QaHnEA1XTKzgqfl1NvFUZZZRdpyPi2DyV925m0sMonEQV6Rgdl9vpM+Sdb9EQhMA
J0L87cgBrFSnepzEkfOhXwF4shktG9ulCgMBH0B2lO69q64uKCJR1Z3l40rwU//E
6rUrv+LQNKl+ZamtTUA7pxueZtZT6DKOZn73UlUl2bppofXxwrBL9gRgSKIw6I0J
fJdVeiU400M0tFAUGMSd4pp/TNBFHa74liSYaS21Nf4LLKFZh61YpcT8ehRwdpNX
BncEUyWA1fGcO24XS4f08sCf+FWZSQHOmP8p1uQf5rl1xd8Zf1TbfBZeeogen+GD
/eC+cQuq4ystwes9/0maa367N530dPK29D9gkmbqAkzvBLZjzoqk7yvIE6Ac76i9
jmxr9lDmJDlO6/lDYVaY7iSQrlaja+myMj8nn142u2Zbgophwqqih1tDUORNcNwo
Pd+6H5Wj4DAAf0gqXzpwFbVf07ofKYP7V6G6KmKsr9mzNcGbkWxcF3E1XGJQc8pN
Tivo2TnDUFHZoX8zJxD4welk6xSUpsgyzOgQ1+Y5EcHN2Ex913LPya5in2zJ1Ptg
WBPPohcWG73VmFce5HCyttsobxIovIALOeWWy+5JO8E+mSmWrIfEkwkh4/bbpEFB
Y1e2sRAUVpIV2LVYS0lMDCcHgU7ruIb6P99yvA2yTe9SzNShpgVMN8058SS+XBDK
M9l63FbnQzo8/9NP4KRvlUObSUDXmqSAukneEGq0Hd2ez3g+c5QMeKhVG4kLya1S
86nV1GHa8iR98w44PH5oTHhZvSuj4jqLfHBo2zMYli4sid0MPjLPYURBez7ej4wo
ASXQnBO5duPSGbNwEQ4I0NykcXQehUiTPA2sSkJD1MbcLYVABZXakpLKBgJuEQIa
GtBPCpezAz6Ke85T04YVnyIhvfLq5IHyp5oOtGgPPP488jJDF50nPnuefm6fbrsv
V6qT5tDZhVvt4yhhqDR3oDLXLBeGcVVZHROJUJ+Pbt2GOAdIkM2XmzhGEPNFCtYI
gfDgYBBzyg+4mp1WAWhGTm1FqYbnrbPAa9ha6bjnW45ylEve/3PfBu6PKloKv8QJ
bJOKgsGJdELi1JAgF0ZA3JKS2lSbiOyuDqj1QR76Yrk4Vq4Z53rAGlxkaTYROS2h
S6O4U2Svhc8DsgungtRdLcBSjxLsByhjt8Q2SLfNOzOWLBhLFheQ+6jnRbeml0sV
8tqQXKE732jGArez/2lrKrceluLqsRxdUsmb4vpcadjN8rH2+u6kP+cK44UvpOJy
pTz0/2zlFc0bfeXUI83n24J42jXau1GjmZFFxZirv6P/voSwictHNYAaqTG2eyrG
e6Dkpjv9AlKltS2PyBT7Qfo7GIIa+oyiAffeZnu66Sc3LO9rlc/qrTFKabhl4LNy
jGBQFiSbX9iiDuSxoy2J1h+DMQ4eFH8qLw23PFquf+0ab/xoYxr0/IyCIB6Hct5o
ghr+f+P3CWVI+87/wMNOYWFK1vsb4vHMQk4yWAzLQukJZvp6mROp5J888Sww6eO8
6rn5lWGSn7jaK+on474v5HiRIzl3Fl+RWJns7umbsGSVUKG9q+yGD0KLrizKuBIZ
mUkHOMamvoWsYME4uHoaE/10Aj07385wq23f/pzXOWUBT1OvVtHetNHOU2HfK9we
PyYBCJP8p2QYvRSyp2h+kX9BRNC2CG+ragOtfCiY7egFuiPf/3h25OkpLISPRqQj
6mFgAVXB+Ma3G6maE4iesTDHuO9mFHCSbcnAvTw4Id2Zn7o12W6wowryS8XopLM4
ovFJWJznflbdYaWCzBGtg2/zGZZLnRNUBIl9xORX9B0+Mm86PZEasQfm+fXVYnIU
HnQ/zjU900VRLMtktnjZ7E9t4Zs55MdHCvZc4fW3LvnP5MBbq8CJw20D/8OiMSFn
ExHRyrjurM3CDDptHKTJLMyRBB+1sRHFx5YEEZkGKPUyCb9H3EXcE8SfZKVFcvgy
/sB6GK3KpuQXRPpzhDG8obcrNkxTo+wOJ+qLc0CaZUqGS2BCrcGKGD9hnG/ZeeIJ
JkTRgz6XOneH6y3uLxNheuPac5UCKiTjNP5+2wIh1Ne/HkxPmnh8ontvfHC32Lvj
uMwnfjdhBUFOIg3rGIboRC/Uow9so1ptYZ4HVF+jKtPT36dbOrKJPliJpWVRGME9
5TpRJ29Rq3D/dHAfcphLJdTKlbRTC3nQi9QRO4RyVyLVAQOdmzsOlzC0LoIF0DmA
d5DIt8iWSucPziud1JaaPEZZOObB1oi74WxjF93G59SS/am22sxPEfitMDXst6lO
sMatxDC23sYLrn3AANCLA265/nHlZAOHw4eTeHfizInPNBJ6CaLNP12gy86rpuAf
1xq6BqRAtLg7qI+Nxcv0XoWCBuL3IQD144eLVbnnep1PSCA4PSS1ZezJKjxAS3i2
A3eoGL1PGlO5REJBkJ7C8VTH2EO62UBRQUWYiJl3qpoABWcI+ff16xftP/Li8nBJ
c8rgBgs7zsUOdBcaN2ye2vy6qX2/kkRaJxDlPj+6DNiq7OkLqWSCJDDoGXcwjfhR
vBDgMe7nZcPi9IXj6hZSzl5gmcDBfrSmjC4dJHHYD2nw8ko4ZbcW1p8GAqLY3lsa
/p/RLYXS1+2E7xEm98msvFAUiqP9HE2VK5i2VpVzWbHLR4JXBWdSdQRFfk67bR8t
S+rTk8+qQWBu1nubKCIDFHa41T48kxrLbJykfSxQpGxlGlvPrbW1t9MFMAmSM9u/
PhiFfoiqAAfVnXjWOvbe7CKxJVku83T2w7IwfDvkREn0x4Yh5T2vxZLjjzMH7PIe
kIQR15k/+MzsLzrrozU0fDIHM6Vp8CX0ydZT7xIuJgE0/BCTCnElilJHNq+/RLV6
3T+duIblb8wzpbgEr1VwbRPxIiDnrAsQRuw9OMokWXYv1LdVl6ddifWkH/K0nn10
tqGbm9Au+XNAI8gBo8togiec4y0T7QROgJosrMFyEvvd9+jR5X9PmmISydy+5+bV
f6ypM36rBF5+OOV4J07rJ5n8DRQYPyXYrffku0Jd+5AvyN7f8ATwVRVuzAtRmfQm
QcTvZZ1aTHTQXVNK61d290G0r5FnDZjrLO+WlCE7KtE5r3K0686VgJRo00lLuoeI
RRBm+w3V5SIWd5lMcHwEN31fKuq2/3Xyb6JbJgy6xMM+zxSb+hkNhVZWaNbtoW11
yIAMQ+FG/P0KTPafM5YA2j6KdhA428ZnAG2OsOtGNXs/wTgVy6B9S8UVQH9Bv+vj
c29CBwXWX1Oh9sasXWj4+m7nS9bwoOz5ur++YM10X7hBCWImkllyuCbbz/tALjdN
LLSP9yzLoamOg56oNrmHKyGpK6sPNinf6mRZd45UltCrFVbC6WYX91RpyJH6EHfU
BwPILHpsAXiQr7YzzT9X6I4GFb+fPZEvyfKNWJi8Ya98yw4gYJgcUaOLEkr7WyBO
EfntUO6yAgaZzjwnPtwEjB7TcfF5PkdIjmnQo7SrDfIkIcDGHBU5NNg6n71Cd0J/
s/dVOkJbrTOqRyEOV1hb9fNzNzsmuhNWNHjflJZVCbmaMs3k9i5rpXarphwfgfmm
T9QtQPpu9E95DdirC4PRpbqXOd3hvIIBVCr0DL9QjvKxblLRlWqWLUHgX6qDpEmQ
pdudmN6KDd61+tEUJG6I3+BzYXXC5NzLymrUQUIky0INQFFCAw8VmE2tSHSOX2yc
9C0pMz1XbhjXLlyCHAiepHcBzXEpl021lqV3rUQvE55xg65tx/3JHVNbZxoj+/35
WL0L14AcNOvCa13ugfrkZm3ErKvkH0Ep+JoeuytRs/89M0zTV84j5JRsso0RkC9b
Tv3fSGoYSoIGgHMXXAG2E6XpIJKswyN6F6ogMNqQ4YWZ6vAazLOVYdmp2yo7/1ZQ
6XPcKsHilT/OQzz58Utc8oKYBp+73FToOcKeSBZX3zk32DPhV9BAUMowhjn5Zbfp
QeRoH7M+iS30BzWGA6KEIp2j9rgVtnqc8v4F066LfYNel/4PXaZ7lgtoWN993iVa
C+lmjGp2LwFZcHESOf4FKdcOVbmw1SC+S+5PZHysMnrdAqZZ26CZBxkgqL36XfXR
IXxi/3V8RAFzPyjuZ6pmHacUDRZKCz/K5VBI5psTBr/iAqLJTq9P/2WDcpSypG+0
PbnDdqvwQS7pWl9zSa8Tg5oP9sF7eOMsMzfKoN2oIx7a6xrplkAk+68bTblOlVrr
AzzbAv0FE4S83YGBg+/PReOzZwcc97qwWtmMitYCI7f9yR2+mEcoqO8C9l9BiHTj
9e6x7dfsu2RuVUqzu46dbz4jyQQMdvKdZ5waK29zUTuqnp6OR72qHySe/nHSM850
fZaoFaMuV3Jt0pfPBBE0sniaiqV2aw78p/v4PzndKoIwcIsWISwX4t+0NP8R+Ps3
+qhTOtVFK8+a6LCFrr08hMqMCxdblLlW4vNzW2qx1uUm6/FjQjQrCNDEB62F05uJ
SN/zXi1TwJLhWsymFk8co0jRR7qOzNrVwtZ91WkoMYC4eSKhJ/2Btryb6e47zaDb
u0VL5Gme1C0nbTJyyKrEEu1FNlYqaoTJUbATXDLXRXUMuKz5/RhGZyqUbpTHDdQv
VN7q54mAD9scYdtJ2XAbf4p9H9W33quxDeLd3OvOZPIOrqHvxuNZPedP7j8YvGNi
xHboROybQAaISNDuXezXGDjCbNrpFESx40sQ1hWrZgMubR6FgsCHRskvYKntLikI
J3IwvusnB8nkOPsIIeJg4rhdBpKfs+UTTIMmmBmEA6yovQMQ4BQ16VoX+1tvoQpK
FalLi7AqzYCsZocQnnhqUbovMxFU63Q9zp38HxMAvXLom91S831qYOgRbVcfpkL9
/plY0NOwcJ7seKt1+uHVcPYpS+f/W7gXsewx9emTj2jIxAtZBzkApHINk0V3/KwF
zkJs48/yCg7JB8q7SiQ9mkTql42+c7kQtjX1pL5qF9i93KRVEWkLs04dGppCCb9a
OlAAm/DKFwkThmB3EkcuSx2RkiR1lEagE99e05H7l33FhcWMape4U0TTH9znT3N/
w9Ikye3kxMB00EOJGXE+7epUd88z+sBHspVIdcDLry49c26csmrYO0nFk9QVMElg
wJgoyqdR0x6NfrEVN5fFhHHRNYHHVajf2tCTRaBrLvTo9OLGtWR5gJqBmHGRC873
l6DyTtpaTLVwXa93balHvewu3lTwa38Y/snwfwebhBcHIbhhobpSDnZKKgWqxx0Z
fgUDV2zZO+4MdtN8FPzz0wFqeUemq3UUkd4ntpWvEWKwut5DXQMmG8+7doibu6FF
rS0VMhcwcIpWgRJHBWhZ8BlFwjA1kuTgxMzyFnweqpqpPK2vtFkqaUl+gJuZrNKu
1/Zejni1S9kZVtba0DJhe2EoCDZ5rrl4OTx+ND9XvQPOxk968Z5JpP1Afb5fMQUO
0Nt48QV+TBSNlqb3uhzlzF/R4KJDiEVWUjgS2anh4JIVAWVLS2cfFpWGilS86EJp
hmvXDcs+5/oWxPXawPRuQ4wa+vLgc00dSUBoC7LkKgc52U0EeRmKTV8RLwuEwi4C
n4pWMqrIgEN8buMw0U+kEhhdCnJfDv2U5PGOkMw5qL/jBBAau1U0iiTQht70DxgE
7qyjw2Gz5ZNeZUQx6pNFJpHpJZ/B4CB8vUvPFr5wrrHUGrBC1tO7voFBcCUedX5z
H2i8s/DQUE5qB3icfQHTqDfeXHJ+XC04jNpi9hd2Pp5VoqU9uJiqhGpsWZJytN+T
hdTR+qM24m8DDDcKO+JQ9wiGI/6s0+B0HGdUTWbYmKo7vbamMCwrqpdayOBFX3In
xkuJ/dacHH4RfCD7L3CKw3zie35QfT9gZv6Ld6vKiMbt4LBnTbIGuthO/q+1zjSz
dz6W31uh+miKj560KiLfjFqK9D1HHJyMPiMn+9MByISobTN9GvL7oSf7reYzWcfs
TrqQE/M0+s2sMpObb02TuZtaNZ2U/uq2pPh7ogx6LPG5Y/EOyP2929J3P4MUc2i6
zi5yTRRO9r4TBxwtEFlLyY/4u4a5aKsfW/xlruki3YDxw+zElVp/vBk9LsCmUrGR
mFfG9YQoIvNM5uFbOZ8415VL5ZMs83sKSKCWp3ppMYBwyx/v7LvjQvPbbtLnRg6s
GO1NySygKZl1LrOJv2Vi8uYnH92pcs9aE0l4+nTYFLypiNyzpBxNSQgLZNSSQ4Wh
ZsPC4jFEa0Oaaauvq8ytYLCJDljIJMSjOaOZXdCdgA2FXKQAOQhm+VE6tm0UdBOD
vE6zRhjU9eiWhl+O2/Ic61Ln/RxA40OVZrk9xG04JBHdNyP3XB4e6KLOJI0xLnL3
/mI+5g+wz9E2AgNnx96I+P19U87LY6EXVA8No93JC7vbNPzn5aKwXNYcCEAcpFq6
8bFISEX0OHBY36nXqu+VJEu3vjddSjwYDPdgbVNMq7jOHzb+paziLa3oJ22bDfr9
tSIGOnQzd0LQLbrUt+RTXBwOZYIILcPo0ZgNqMcNCzhzsBI8n5iSVJ1JUd8zSeyp
YDABOYMSGaFLOpC74RUxxDmNijqaIOQyLKnuwbHBRL41IZo4axqTTyPgpFUKAuFE
kQWn3toFAtW76TOXruFceAUxUwTb5POhCu4NJ91Ofh6Ec8p5ncpmgzqGJkVO6X8j
+hEFR2q/4qH0AVoZrorcc+2O8UqwY+UBvjwNKXjrk34tjPGniR13zrdseOJVsJWW
I5RTGf3ri06Q0JmXfwIiFTVg+/6rkGQ4BMEac0O4fIOmjV1vqCzrClyy9bZGJ7/m
3BAwm6NbE8T4uQSWoMqu2FHE5f1/XRjMnOSTTR3MHAUFK4zUCSCykbTi5Te7Pljk
+zdCSLTeWQr3eDC1KYN8YtVcgId/7SB6tNA7aRCfNMBLP6Yrmthegr7EpRwztIqJ
aSpsARaZB8WWT81cSZgk18HDlOXw0S5h6MPtceBHCiiKUUeRFmffnwPrld/xIoZi
k0FrmIXpYdhyFv7hoFecZRnwIOx3PziWcTBTQoz5dCeNmrdv5s9tv8z4aWoYBjup
c23Lv0/qWwha5E7EIj9VJH5LfXZ5Pd50DG1ivMtSYXaTbjGfa/ArdzxzEb77TIXy
qfUAF2E4cYSL53ud4q+ty/JIvYjDPQ4K3yO5yqlOjV8FZBq/Tt69t88yFa3GFFMc
yPlAyNW59SzcjLWPNNRjgvNSeACBZJJIvrE7Kww8bFtZUIxckOBjo+/e/1+W/EHX
5IkvW2dprKup35I2lbiTT6d90y+pav2jsMCRt7Ht/fsgd9mVYwTqJDrKy05hXp0+
Nwyz5eUb2vmhdBbr9H1nQG/pWp3v6+H8ehy7XcGuOiLyCWlgF5PYYrfgydIgT348
5mhiZRt54dGzP53P2VrCTR27RvETxsEhlOqTF62zgbMMqJZTbQkt+iWiDefQi17L
5jiqh7aJ+rq9aIh9z3XUzq5KnNCvQ/+ko7K3L+HZZ2Z1lDHq4x/oh5kVMcXIN489
mg/d4YEWNqwqE/JH4jur+ire7nV6eruQVAnMhknGJ9JUz6ZLu90JF+sJBLQgNoeE
LehFqHZk3Z2FdZ4cit9qEfww+Mb+d+BMhcnrJ2OyhpuLcNV94ILK7pl3trGfinZG
rOjZk5/GM+8fA5GQbMfUqJuq/ganEizb4saAemlmW/8YJ4AN+HytaccKnKFk20cq
PaF89v0bz+bBrW8qpYvCrhTIVXRB/MAe1NCDSocIZuBT/KiAEvzVJWzvRllQKD9o
U776sfHQvqzCG0q+zA5BGlcZ57w6n5fo9aoYfw/UDIweC1RO7FszP9UuYlh2mFnK
9D8SDq79BKgz/dC6Otwt31HAl/65QacTvLp/txHTwRrDJBlwkG+149OIymJtoI3i
711q38JsN5nbYjXJKfU/qD9SILpj67Vh4LfzxkvKitY69/m2Fk+wtQ6Z6g4C0X0l
APVcAq+mwY7sYRoErdP5DmxcMFvmx2fLMPxF6+gSXD9db1WIGw1diTTGYiOEKzDZ
/xhzrsfvMYOAjhZtUlS+aDIyNYVViOzVsIV/lcxpkiEaiNbm10jun9jGix7Kb2Lg
VVl9dUTYVd8BWlfsvsnLjVb4RvhOsV/jp0COplFvCZJofE1egKuA/7BdkvGxIiKl
AoxnG1ZFqRDQHaY1jWsjzaq0vWNmreJtAOCBGYhfYraoOJ7dgUMPBSOXYdeLIRey
inRpS6jp7VTGjGhS2snTWO5SD3oz95eL7pHBAz7vGxDN5CxXxFH70cOMV6cMyg6l
8TK/gCbLjBPxbt4fg0J22zctQS04PFpk/j4M96xi7xVhqxfxzGvgYANWg0Sd7UM7
E+M7CMvwg0B/8o2/VOz0552xQdnZQ2kq5qebAA0SGU0DpOmMiLj1FA9VkB0k/nmP
g87tSojcevq6ciB9XV2htxrX+dVoXnYxIq+8ZlV/P6k+5nb4tpV9uSKsbIDRGSzS
10+Dp3qACOE3H4xnWNSs09uvgzXW20sqEub9NI7OofYKXL0SmrgWTWmrUXm8LwCI
yC1HxumyiAk1urAXLq8iwAqa4REmu1PvgWMlIeWOcews5qUutSPAxd4LbY/VaZNe
pHhwJCIS+d/eqxEMw/uqhtdEJ/ViQI4oMV2/e3IsAKvcbv8g4asyynB/fhXnsgK1
o0hNG/cpzmdel649um33gnZ0XQS0ss6QHA3yvn6nK1LEzL8LbO9gYzzj7ilVtVEg
ZZU+QmoV043W5+mOMaV2kbevcL1AQ5OEsGy9acEVqeIU87yB1d97/EPttWhEJNu7
vJEYB0jlSO5ZPex095eVVMEasDEcSKlgqqzRFPiuyC2n6mZyLRyDTBqb/jHV2cZq
4id4hAQKDxCxSgtNU/2OE47lcUK1THoLN+4BOWpa/Luohq68iM4bVoUIRVlql4v7
d02Mae7fBrD5Nf9BIBhRucrWnSdJnRNte50988HhNdhe5W0B+UtZQ5pmHu/HyPI/
OOA/qy7D4JlTYqV97NA3l4lhuOtdZbCTaFATBNlJHmWJYJ9nlStrr+JaQaX/eM2x
w5l1kIowu7ku//0rQkxSqDavQCDdRdHKjo32oEdGg+wyILWwGmnWLODoTUNjZ9Cr
kwawBzyCgJg7PBjCxUdcJZqyzRK30Ye64//7RYtBnPVI2EbCSHVH1jIaUEtqOFwd
c6/ibelGqqIF4vDD1+ePWDc/OWOhqY6N9C9KQg+5WmwmnK6H5uP8xs09yUZ99D5F
qsNSjJ8iKNMSEACwoxn4ZUlfwNqWPVL1SnOUAv4Gq/0QGLLl/d1MVZkDlO/xPXio
qxQch4u3xaFPDxqMzM1ZBl94DCbqoY0tqw2zsnJ4CB/eifFW8D6o6VGBzD8mj301
qSolZ3FZnh/hWxEHK1bbcJl2aARddEJsu5To5KTYG4+uLHji/A7ND2nTpSmTVhUK
NYYeAkofgpYIocEJN6+JtGSV8qMYsxMowOPwDZx5skj/sN8Tg9EagzE4vZ6N6wk0
/cOXV8ySGbvI0Re4k7xBrf8dRqXYZQONrVPZaCxqb8rrSaMYh/hYlyfeUiFGaCDL
v9TV6IDHdAJ84ersEbGtzALIotnJjB29oe4JSUn+NfAaTbbf5wM0baTxfOMcDw5d
BrByrGQUQPaqxcL2vrtra1X2ynHYeIUoRPXJyV4bArwPz9TCaAklOdZACBprCYsG
9jJg+sn4hZ3XSv46yZyf61ogG4b4jQR17alVyAkoEqyB5nT42z3fNB66fh7id8q1
RhQOc3TUeF7f5AczAC1jPQTXFlIRN7Tmr/QwhB1LGHi15oLkmSf5NXmVrm7CuN5V
1PIOYwOlAachsYjHWI/M5HiQHz7RF7Tfy8ezPmwjp3wsc8vJOu8KURCeHrXRi0cf
ZyvcMNSDCevHune/J6kZsADWNRfkk/J06ar6uk/GaqOYXk9DGkaKze31kgDMvuiS
JyiqepdBXPCVMF+RGPg0IvXMA5TijNUKDiSuiQErgJnnUUwRaP+sUlvZWlG3vDtw
xFY7skx/IKQpnI1bpsjbZ9UTXc2S/kg9xwQlCF20EEDu02dBJEVoICNGR45i/9Je
nGRlGrEb6KCE2Kffq2/CGJNVG9ozS/I8PGFBn39193yGyaaNHSDRkMsHOvZVEOm9
JwV2P6FFbBu6UcdiURvN0DgailttWj74ddWIDxbytnJZmnZwgACXMjpX+XRyUCZ5
a2vQTz7PUfaQsh7mKi2v+aFDudhbfRJOGbuh2mlHnip1CTMHQYSHKGESKkIesgcB
ONtxW2gd7sRFe7qEaiHxbmhAEHj0YDuTToYfZ2kApCxMYBNV07xHEkpiqDF/TiGu
CY/AAQILHYvRS3eciHWCnH9SEDQDjBwXarMfxeBxNdPPI4kXyvhKdJ6sHIlJqhCS
CST1fh2MbvkwUwu2pkhI+uJTGTVJRw1VG7ZUjaKqpJkD+uaLVLyVeFnMq5UstuC3
q0HPgexLJwFCu1t061PlMbNOXC1KmsaDp7nqcwiC49MBK2wvm9emsO4yCW0cRWxm
orwmDV5S+HbtG11ImN8ohfgmsiLB0vnQBNwX1tZEUNi2DpZYr/ExI4y9oWB0uR/C
4/ZY6neiC12Nc2LYEPLZncGhvQH8WGI8sH67yZdhgvCxVZhnH7A4x+pcLjCGsdmK
p7CYZfDd+j3gKJRPVe1ac3J6yz2OrJIRUadnuVQUXqPPBvEOAiA0rxI6rNmYtQCh
75a+eZtBQ8VBfH6Nh6oOjvcVcKTM1uqkyk8veaL1raEoHOl7MC4sp42g7ziCH9gL
JeZHAsrnO1wd5otuIeZQ8MLEU8gEarmakAL2y8P/Kfomko6HCXq5r7VfAbDKZo2G
FVN2kggfWgpFRlWG+OvjR78FVT5Z5RbmCvFpQyVXxIEfB6jvgpqTRLCDG6eB5fkk
/txKaQAdgRqS67bUhQ3z8TWrhfzNh6AMH8opMJgxcRgbDFTS5YaZ1xMTxI3jirzM
gTM5wEnFx/XmDsyo7baHYWzgDkUHwPWwO3Ogu2UPlXHzO4y6NwM21evzODB7zlHG
oWKv49Ox5sHz1NX6bH3eAuRrZ5QhtV5H5nkzAZ64A3CMzLT5kjoG+1vUvfNvUtjQ
22YgHEZkhhgeQoUAl0jPDb9V/VVwpH1lfPfBBxlUNpxa/zFQRJISbOUYuc7DXEyl
Ygyc1DHHeXJUh+l4CxfW47PGrOEORlxtvGHgkpb2gIHqMb5StLzga7w58XxB7/vz
Jyi6EyrAli3XtIlP8onZnCvkkL46ZQL5fpNch66iSwVH0Hu7De6YPcGXovEXe9j+
QT1P85TshtgFjre+jteqRbp32X+P3BUemeXQxnXfwLzdkazLr6BCc70NJPBz7YGh
0cpzGJRstxX1G8ZQoR9+3O+m36O9LIZ9SO6CV6Ool8qTeeRGrwM+PavuV5JN4s9M
4LgzLTuCUlLKpnQnWPUO46ZXaIkf30l00W0587bh8ZEUcZunepvFOpdHdihnzidF
/Hawbm1KcTsQjtOUcIjDMdcc1MZrDfxpEHu4m6lXx9k/cMZFWdmXdaAi8hc7wa6x
PIHi3UxsrHTfLGfnA+K755is5/FcOy57AzCqaRaiDeu/PNJRIToxrnQ/Hyrlt4M1
Fz/GaMFdqY20w8UezbdHnL2CBOVvIOMAnAehft2Ujp2k6jGn2/aT6eLLDxW24Nhs
At3Gi2d7rYI3iVuvqxn/KuD31Cp999XXPtUp1fcrGl/jy3hsp+V3wG+9SbbX9oBp
ZhhSO1t1/FJKEUU71Cc/WjMcS8o/ng6wd0ONGMy6yiqHVAHFp/+nAEgvPIAEu62l
EbBCxs7G1MUBA9CT0ry5aP+3810gibcS4OsmWT/IUA+E+pYoyw2djRIJkfuadENc
GdsdbcXiBl0OCN4JO16PgDXePzPEcojJzYahbAmOwrnCpHPtOe4l5HNjzQs01pXA
3n4fA/89fXFLvcDySMo7q9RWPbzic08CDG5rYR+jwpbOhahUMKwXni0erdJ5ilY+
ezkiPQDsexLG38bNp5ckU0dzu8C9MQKfz6tt9UmXhnIpp+Kh8Z20YO/0nyQE9nFH
lrazNVsecXA58a5JwJOPgB7rovx9hIXIYiC+N6Hb3eWbk9di31oiq8EK/2SyAk5A
fj4zeCS8q/JMBg8S21cXCRxwfAw8zS97jeL4e1vOg6tBkJUpk1lFda/dLRgSf0PG
USeR+tuZeMrlQGEnIAX3tf4wA3C+2xRbLksa9aCyXRECoj2gSnAUzVrpNAvg/7xo
QlO/sLUJpjlN+TearAPOOV5PB5l0QotRJLGGGkg9iqDuxOByXftOZVIw/stPrgiz
3Wow0BPEmzdkt+0kDfyFy76EI+p6QlVG/Bx2mEnCCBq7N7ClgapGPCFoaVtZ3Tts
t8sBVw8nCtJTxCC7OlvgUd4RFKehXeVWyD/PWySAQLzFknNkJPcyRcwbPuZFUl4L
bfTRr8EIDZHDIFrH3oOQ8yd8Cs2skHoZNdyTR3zj5Ba1xVbU7dGAM2x7cTp1wg3G
k0/hg4pnn8K9lNK2V5o+RypZdzeAgB1QTyHLDye361oj6JBEV5wXFxwssQtkL1a8
uHUXlSBvcdgpqWLGrVlJaklyC7Vq4E9H/KxE7B+vxaEEVxIqHXdVtsgDQnJommym
NJ5rlck5VJUYLUg+/FKAxrF/iW0Vrxk0lK8NzV838HaVD5prxmeDDVhwZwiFfI7I
Jg6Dc1seBiP1h5BGktI+ATqnGonpVHFnrNcy4n8IqMP3PiirwSkDcJCLJiasGHCp
b+Wnn42fKmxtCDsZbw9S1CV6rrue5l8eCJXzO3KGRBzYTBGR3Gv+5ISMots5VRqN
4y3FI6fNNSiWjh6XiOep2xATH1cKbMF5GPseu53JjUkWgHWsHBqmld22oMBAlExV
bTNV0rdtHDagezEGw0gXOxpvBRE06Lc8n4999goqbc6kugurMchPEcVFWPjbw4hg
kzs3x0U3PII5iREXy7R+zW1EqP4Vs6s3sHOisKxkYKA3rhyEaQPwR4a2ZRLr5klg
28iWkNTTH82dyEEpW53aw+hPxGJNKurPrFtuMOzMPEX29SAc1Eg61SOWUfnWGHL1
3Pqg9EDF4bO08YQgxEu2uFL0cYgxhZuVyssYOC0NfDOtL1kQA3r1pQH1mCDDoHJa
54NWgUkPApkjOy2Gp8gj00ZAmS1RYVw9cr8wIfzeJ9kI7y1WLAMEYGxj06M6nu/W
+vxYD7O2t7lFxoZpttRquxsDLtLc/thUpuNQ7NZFfygBe38eTTfzMsP1BRJVK2rZ
lxpbaznJtE002tQdrRrHZzeAmpTZT0IphbSL4IpiOxGo7LKrVSusHX42EiW2rO3f
/G2xpJN3/3gGTKFuTzStrjFkB46e8R0u1dZ+DNPilHhQhD1mS17ZBqlY7TtL+HuA
FfF2M2vruvhFpIjEY36TO8aWFsh4QzyyioXkcB7hBALNTde6bm8Fy0Tw/vI1f2ss
Q1bIiYZZ6PucGvzAl6JDLhAipRRWzW8u8fais3G7z8sOLDRxrItQktYfSEhrSIrq
TSlT+bLceCVpEucbsfYkxQpeoeRGZLMDdcwfoQ+NDwKHgHh6G/YaAyR5RpXwhdTM
qCUBj09dluXMsNQcZ+ztC+e2FtVz6InpatjvomSyqOHeAIKCmBTzNN/A0OBEW2MT
eKGmHrvX+muc6LOldyv/bM+QuvwTGC3Ya4czsqRphpnwfV1ZER62Fi617nv5Rj/U
qZDlegfHFoWMrYhseGwSyXt7YVCQ3rb2pXB9MAavOswXZBtM0iofqzySsFwMdDZZ
shbZQ9zdDXRntmN2O70blyYnEanEkgx6ghj7xmMZJZPS8Dd/nFYN7Sk0OaNGLXHg
o8pVxSFNWi28QuKVbfVB5yj/7AjvHc1Uzk7kuHPyqzj6xUn4G9AYcXvOhRAN3Sp5
2gtz+hgwmq8sUEHoKWXJGlFBeNynoTErIsCQtZicXWZ/zBV850gmMjBTP9A7Lv+m
pTql603CtODcD39bORf5qZ1kGRSSLhBTfz3cffs1hHfNN2r+yJPwL2cD0b8b9d2y
51IxAWeaeyEgcm80seqDC9xiZNQtH6W01m3mx3kWwhr+Av1yWvzWwsUoEs4xxZYU
VQq3grYqiMe6ESaHPhVlobSwLaCcSHKlgszRrJmq1QdqLU9+cLmC919z7miPCi5V
Yg1TO/TPIpZIEJFSsQxYqPUsUNMj2KDSQCxlC57k1g2eR/0icurTitojclyHYfjd
24AJEa1Tf5Yp5AIrJ30WkgERy6LHp/IUNkUE7BZEkxb5qTWiZWY0+8Lg+PlYIBZh
+RT+WiGEGfAp60OsyMPOA+KoRE+acgpGk9uh5IgJOYipGUiUxB/Mg75cGwG4lh/O
qDk2DdfTUUzenNe6CZDYhWgOWP0CP/OHh6olaraXWKqc2NYsn4dI+ud+apTrPE2s
kb/O2u0Vv6scjhBycsXZQsNJpuk9wI9pm2PdEnE43yOAdHUgBqNa9ilnj4Rxv1mD
umxBkMrf7J7x4z8EvkC/zEGqa6NnalX0v4PN8Rl8l7uA03TABpNNWz+lC1Eqn16l
SzM/NfNH0gWM6nksDcDKGbDp6+rzw3qovThAxjO84x2bszDl109mbF+pZ7mR4kAe
1PQNGYw6dWRvo57oJ6hB4y6FT9B2aqxtfHW4Mftq+pcZtGobpfAJrtPc5ykq4LnM
lqbwsykcir5oKIFylk27pRh22vfbNtp5yWFq7DGWHhq546CXTyX2Fi7V6eJ9yc9J
Oi4AyKOPiAT+fYCkX658WMiVMlfL87x0dh05UH4yYBwODh463RWbfmDRaHtNF0cv
lkNz6rkg2rEUy7vbdn0hCLnGFVjthq2Ry0F3z+/v5KwylfqcqunEf9eeMVcn3qdX
WJgs/tXkfhrd8rFl1Uvw0590hPRnpooHiQpqL5UG1qzpB01xRhgErcOsaK5spY06
jLHUeIcW7PHu7mUuJ0Qq1TBXWfP8EYeQP0h3AZDCZrb9U/vZ9wAPlpAO62HcTEN2
uaxzdz3Vc2l7g41sahpa7uaqd+kpq3edXYoZFn4FU571DCWN6i3wwposBE8DmUaP
LuhaDf6PBui97Xde0yj/KxYKs/vw3EIJdafHzkGbBLKdt8bf7nrVKTiL9aIgzQVe
xi5NwOwWpWrR3nXn7ShpggzBLWwEpRhG3QhbgTmlBVtAscGkhXkUJT0Lao/JR5tL
MoHIVEVLyPcoFfHxBB6rcgjNLCybvP9TkvQssdzsyp0gH6Gr6YpYED7aymDEatD1
3zE+oZBadtwHZ7ScvvsBM9ivN9uQ9VId4nBjm0z+J59nr4+tob8iwuCQXC9z9NGE
Yf5N09A7AqlnxIxUDCb6sUtMbmr7Kzr7+8KMFyPVyAvLH5mwQN4nW6Naedatt+qP
hqlFaE1TIpZWgbr4XKxsmEZQHNtFy0/eUyclx7PQ04/ueIZHnDkCnhggkij8Y+RN
l/nkkjG0KVMuAYMRtow/D+s7rKGC9CkDFoAkz/4ycV91OS8QUtjp05PnFW0hH8l9
nclFVaDWYta2baflKwdXToE8ebJOYMVVWatKOePB1ap2CelOyZVzDRjeO6LZxOkE
3RKQ+r7Tn4oumbLnFajtFI/JBhPi902rZNdSA8nFGHEHsPgV1bBuxv+rEVf8EDn+
1lmHhGECH3MisUp7p6IJWJX/ZhFfKo9bMV8V6nnjGcEl4TGh4DMUVUySri2XR1iA
F2DKlhOWt+dQol9qP7Da91GIh64VfRR5+b9xyYjDbvPIlaBCVFw2NO4tqH4TL+hp
dR/Jea4cbXzpohBrz+W/cmIUhFl93ePXshmNNudvsSneYbmiNRrVnfuWEUoLUME7
nPf2Tykus1VFaulcb0IFE4yV0YNjd6nQRkZ1iq1FhrLwejrGBIqXy1ZRXxcJivi7
5gs2Mu4/9Nz1AymZL+YNMKG/uAEY7AFnpCSU+0o+38W8tHNsXHMwFoinjgHK+XiX
APQBDUS3nBkEagA+L9DWN7TZnekE+7k/HVF6KK8edhpWwoDacPAK6PjMrHVwKRBr
KhyXIkxEyA8dS9CL1Ura7Cigmd93brygJe2/UzFKTnyLkKaaKsO4f+g5hMGee3vR
AvRz7I/n9Mq98LlYbtmqfoHPOw9WhVxEcTQGnMgrbu3cdn7HCvsRJtqvJTT9NgAY
djFnda9O9tvruuspn+12eOV4OL+Ck5hCKPDPhxKQ78xHUIiVCiRxAZHqrjiefjiR
7yn441ODT/xBEat1yZOvKHa5dx04i8o6SwFT9wOGAlNJ5KqDq/hxDzBIJ2DbhyFV
mOJgY6EvoHJSe/2w1Z36DBEuWnu298i8iJUYaWoviBv5wKJGXoWuR7orSI8cexpK
mgwkHbCK9R6RSI9pU6ajG8s7tSohJQiq97gKLEwuGIObasc7+A9LNh9VgHw4veja
7dsS+01ZrYXz4bOa6G1l3eG92p8W1vPiAX32zYa7R1Q7scwlYij9mbjGDR5xLNz7
hcJGjWu13UDrOW+lOhsS1tcRDo0KGwMuxOdBP0nXrZLv8uGVWmlQvGhmSOpxoUdT
BO1VfaHNauSNfZXUj+sZXmGvqNWEqhdf+DccqW09KQDTyewg58P+SVqQk7TgjEBj
4OtbRoslE88AVaLuMRDkGmZ98OnkkwMKdJIRnk1OXbZqETbv4L/+dwpWJOQ1qgYo
qsfmf7ckDYBzhBBIOBa/uGspqpXI6hzccNP3Z7gK/8fqShJm3zYPUAfYk42blkCJ
efoj8nknskYivH9HR3NY8Y48QPCWZm8MW80F/FPp6XNpw4VxWN+HujAo9yyScyJa
uJW+IB7bZgcZEocuFUrq/yqLkF9uIN0s/Tam0rzR/aKyRMAbVIiuaAI9AWHb1UOZ
ISF7HfwvTiPzE2iAYKVXq+CPKf2/llFbecLqNDWWcCpu4T10iI0c5ZVdUaP1lY/v
R2JNw/h1zzDFV0YFIEnQVg7q1WGOO7MVPxJWmS/dfJqpeCR2fa8qHEdr0agGEWET
QENBBx5wfQU2o6aEnPG9vt7xYbo2Re/3GExjdsNn+rSOdyaBU/r7RSFtL8simF/m
GA+uiotDikc0rumCFO/NMGzx6iYWMD6czFbvlwxdhpbTLxQK1TpFPbEZ5r1EIv4r
+wthWjqj1dCvucr7NUa+/KHhY4bq87VPISEbAScOdasXDcePSOCTSzBRcPQtYCZw
9exwm6Cc8jZtNDDuV6EPTIR9siTDSDozQTiPAZhjh8tWKe0U2SudE5nWNuiJcsdb
UlPv5QF3Pb/f2fiNsHxU8NS+MWgG/Gdr33wR7DABx6Zf29hHrHCU/dY4cnXWuFaU
5+eeGd1x/zLrF6rCov14kmrVIZeDwDtnQvpUadtrlsN2jUZSjOusy4R+VxMcC9Oq
hCOKE1tiPGy/UuoBc3JbJtvQ+OH5gKqO+AQBw0VMjnf0/bJdr72u8V/i5z08mtQR
0oOBCL5gNBie++B12e+9dQIBUPJ2lwpsffY0+eyHSF/Ym0d9qebuvcx/YpiL7GeN
XlIk46xNInJ13HNslAL0bO/JywKU0M3RCQlKlHnKuE7b8JPm5TDXqBOFZPDavq7z
ph+dD4HTG4e8WZ6BEpfxad7HBt9ZhLdVC8UWz3Zh67HUMJft9VRH+GRu1dSJcgCU
4pVJTiW4xLrAiuEBXIcnlQmWX+vdXuaRi3ukU/zCmgjDiFoVnFJP9enNW9veyXWJ
GnOl0pPNOrdGZ4sm+2mdFBOsmyDgwnp/MEPhpyNyui2Cxdel0Q+Cg0Kum6dhk+9y
wI/cv4S4t8nnU75FN1W2vhSnfxi2E0mOfg3Rl/rdKtnsxPGbZIocppQCYiGD61NR
kskUAq1x6uTXntKrR8V2d5XIPid05tKNz6+5lcAF8fx2cVHDhcVJlVuRmWdEBeiw
nMUTZrwhAckQq1SF6ANSGLJM0WWKJ4aLSdfkRuO1qnTI/QhpBHkgs5TAVhcCjjQP
qxw6tqYNXkfmTW4VFuRaMTnqAx4zsfnY10LV+DGJ8cvMvbhNfst1sTE3qLLrJLp4
PIOUQuk5+MCJwVzgu/21qZ8quves5PK0QIjq5lrd/dB/ZJsj3CsTUqkB57uN2reJ
P26dNswXAdL8/M2TRg6tZeI+E8T8w4/bHYu4KAVzOwgzfhywmO3Offh+XWWFBcYB
8FMcl06otCl2x9c07QSxzVCPnrIkfB1WiLYKOGBwEKAIJBP5OBHIl2Z/f3TyaVMn
6nYqGFE78rgvAeBT2/Bn1AaKvtTwpJTvoxHzx+JZgd2/Ii6n7l/uThz0koTul8qT
duEf1P/3eax75QKWuMrS2iyEHmW4vIEBPuTBt7KfcFbgCBsNAFpPY+jaVS9C6PtT
TMzUV1NGN97kU/8nE5GYiuxiZ1HzidpQSld+iRFGmriMe73ZdC/ze0BJTYmHj2/S
JwwMQ3ctTJx9pDUzct7Ee25d+pddgxA5FNqHcjRjktB901MNoT/NcTYapr9UIfej
EpzZqXxX5JGmvk3BgPE8Qam9U2e19OBXPHyBRPXzkRBUGcHns9XJdvCNzQUAO56r
rCdo7Ba+rEW4x1ZabypvHj/GS7mDEN5hvCTigmpKz/QevjqEooTrucvi0el80JPS
XBB4sO4i8YQqIfcy0HElpX91kXEUKaMDlCpSFuo+yrXRJ7XZM6hSdcVmjhb/W+NP
OqjuJAa1Ty5qae21/HXahriiJROgZdpBtyLwz/dq+rH7ocR80fM174dMPrUDlbhq
kr1E5rs5rRtMU0GfABPv3pCNAzQSFFmjpHx4fPC+jVyzjT1M5kP1X30PW4+/vL93
PEH8ijod4IkyJzV0dr/v8fQyI5DIvp8mxh5diMu+bMUwZmgiuMGvi0ZwxGA3jtnx
c5SftVbgcukfk0dl6JKlows95EWY2eNrFXf7AXb9uynRunViHjcudW7PygGHCKlO
yVbhUd6lqB7+9iSW1KbPnFNjNTWdaITLFh27IfOYW7xtAS93S9HVupLx9v8kykgF
sganZYrhfwmX6bppByDIKjTDRBMyd+e3AysjUYEzj/QxzGK2CyBfmHQ+oz8d/QxU
h7exQJrn/am3Hmir+GWZgFn5GpH0X2q07LfuoctaorEktgPgSQxUPZEJ6LSeZMMB
Vx9saJQOXk+h16RtvCvUqbVO3Kw84bhzZONF59EN/sB0Arlt3k6GYXSoRWbMIK68
yPuPhQZ/x2zAWD+4tfZ+vg6YkowFcKYtLb881tg45yiTyNWGxlA6zWE5fQ2mhRtH
RCRI9iUCeRVywFDSHOzjuc6XNjlaCRFSSicEJPaj1U3s25lrj2/qL2k5MkCca5OF
SnXBA/KQxcXt5g/aELyOpQhjS7BsN5yi6hqtgVUXKrP/SSVnvW+5E7PZQ9hlb8+b
L5tbAlNBdF5NcC1D+S4DuIsXPTjsVhI7lCS8aBlpm6HRZXFvZ4ityeQLKnmngV2o
P4kPW80RcB5roOetlxQzokRusVJT4Pt+Ohy82yQDygFYnYjFVceBUtpm2E3RbnDG
ko59jubROYZJn7m/0kmBErnjZRZHAD8KpS6HZY+PXX1coPkXo4AtD0/4spmtqQW0
0aNJlL/0RkAm+RmNoMa2FTFwBg4qp3NR6VKcJl5QbGjauUckpx/mxl9QbkEi3RNo
OlUt9+RhZLz+t7xqC8YgEbR68duyfDdrjzM1offZ9s23WE/cy3M9tsvV6kLfvQe9
XYwpoKw1hOnSYsV0W0y/UTUIU516QpFEMIfc/Yln7o8+tjpKIsRMsiPPvWVXM2YR
2z5wuU71gI/VimKlWwgMdlpWw4LIguohxnQhVhkgFDnQqHIXoWtGq9PxiG19hIP3
1+TgfGbP2rFm250DhA5OsXalpSTXu3q/byk1fhwpor7KVG6uGwqpFSzioog8Ty44
V2ibLiQUbuNLrHZ5JwqgKJOsyb3O+tTIAsR/aHsQWwN/+qwDmhUVAOb6aLPAiNmQ
PJR3AOxJoTlboxuUC5T9h78CiWl+TL15ddTHcFxbrYdALTD5oEBvDlrj8cx/2j0B
T1SrD2FlLkBtoVYrjFl0KVys3Dl9m3HVAzq5QucYu0guj9MbhnFGu8hI3o49NMZ/
mUmZeim0IJrNBT3DYbvxHG/s/vRvlCruGKH60txJNnL7lx9eQmk1J5/rhKJeKdQC
I5Vs89XdiahpGnB1ciYjxeWH+uRFC7JHlSpjckti5V75/t3WcOBpHsYBOBAJQRjS
edR5O13oHstkG9RQ0MFPe7c7RpDlmoBvRAc2fzwL9Xj0M2eKVtkU1Ozm7i5g98bG
urb1vVyrmpUtO9ZGB/OC3oUdFD8qfMrnY9EZ9BkHJ798gQhInxS1dlXh7/zRt9Fp
RRhRj8sgX/ixkayAlXByzQkZZ0SWHnaKtE3lYb67sQf908Lb/K9WTnK0C86gk+bB
QpVOk9NKUE7uLoPs78VdiengyKoALOggItVl2/JHEu0WcM0VfucWaROx/mUX4bC6
vrzmGmvqw6yUor0sGPIWINSo1yMqJ0g2mfjWccnMl9PS9Qs+QSCP3dXsDKIfyHmt
+XrahFeMY+LusM+d4WPqi32K/GUwBkNHiGpAovg99C689CHN25frq09BxFnWqkwF
Tsr/1NinvOBmrFJzTUi5jpHcwHTxlwpDZgo/QSQMn7gZrpVbc6byFqFO4dTTW0Ja
vtTjFlQAUzL42tiOLWxWhHP1VpSVNd3AE+jxeotDxwvLKtWHiK9MjG/7uD5o4g4x
fUKLoX2DNVV+is6Nm6NspHl9oYpCT3qOvIG7qYWB0pziB22OHnefqIR1I3YdQLaI
R57cI3hv3FCdRZiKDebt6H8+ZWW/fMnLcnnxtQIActOYO3qdqFYiDy+LZ2wuGfoH
p9AQ7WSs/REGrDHbY/4vd/LnPDVP/eYtEb+k8j1WxPHNU3uQH0VWVBWGh3yOmbHl
yq7HH9EJOV2ZHhp4uyl0QdAJND3mcQ/vQgbWGf9VjvDbhd3FwvwBVg0vmq2/8LaL
9i6eNLTwq+7a7BH2/3QPOUw7e3hxMwehQly4ufy4YWvoVMhyfDRjGXXu6OsSBtM2
GtB7/lA9RAvZGrB6m4/O92PeG7NFphf8QwE4bQtyItf+MOiNavfWjDQaWrqunIR4
RFi5PBqRvjxoIviJ5CpCJYLz4yAas9RApu9pzRmVzsrWgxsdYddFFvfV6XSaBS2u
C3ZWrgXELtDVIe+UQlbH6n13p3HXJKZPwcIoZ0ozyYwWQMudm4Zr8BJcykR4opSh
uAOJFNlZZe8awLEa1qKmHrU5L0oBXEinXVg/RkTV+ksTCDjfnGdPLWfdEKABqMQQ
ekbesBV6z4QPk68ajQ3sOC/2ywaZvymdNfPMW4kNMh980dtjCVD+QckVKeW0cj5d
0x4cRltHIHPRNnE01DB24brm5HptOoPQJO7Tszu1VjkvKBjp+0+VEMCOC34RIEpw
eOVt4w8ZDfK+aUBanezlTJjannwavM/FKu26UrIe0tKZkCcOZrV8JuA+xEhr2sg4
X0U3rPHV4L5jgGZQWiRzNdMvTO93bEVrl1lCU4QJhn1bmvvo3yqXx/adEN1V97XF
LglTyhSupaQ5HKZ+22S1e4SIHHy1L0bVByGyx44cRiTF+luIziQWW3QJ3M7eNp5B
3dPyXio9GeVORDqt4J3g3Fkvh1ejtpiYoZxvWQ0csWzii/gu0NB3aV3f8+XAjBog
IEZ/4mec04BDt4WLi48vRmBJ/TIJiUEliH/1/ldWbalffQgmddbzbGfNJ9xyfUe9
eFRLKk53frxuhjwzO9SJFQrdRzWFUBHdFWeuGeqqscT9XN3z5/mlJ3vGIuR7ERyp
THoN9Ib7O11N4uBaTQ1e6asKuCnypd5izcvGINRpCIF2AJ9w87UK1N0cUyiw+P1n
MPDWCDp4A9OYEfbT/FhtSrjEpUdjDb5UT5TsGUtpTq5MN7tlCavMW/cNsYznt9lK
+UGM1X7BvmknaziLeh1HFo9p3JhcDtvFkY4/rvScTsW3yqPp4IczXn5kmwn7PBMF
v0MK5l6z87F82F9pQpAWhQtulEpmSIpXLDl9U1g5+hoEQQuNjxyn3I6JeTd2JUkS
pAJtxmHMKNGXa6yQvnDD+DLyJ0DdrQPLD/EHqzULXPVNFW4i3yemXdM6DM+6sPKU
YIFrR1hWxT2i+XUEa4arIdopT9vFOkNhVxAoVNrAcXd27GaPOke8dJ65A3ldQuI3
3GYDZRUoJerbJ7UB279SJs3EktYUGI8AooEo3yBOTbpts9keizI91lLK5KYdyViw
/9pwCQqQvwycaa0xipCibxaqp0CewgONwbEGuz2oC5B+fKuveu2yyfteLLrjU9Xg
XDyQhyPQNbYQx16UNY7RIL8AniK0ILXy0M23LsYJrPdrrbVjoEhtuZr58nrFfrSR
uspBKZF0CarJcHFObzmVPBbZmBxhs8i/0vVU01Zgb0p3BBDORo9bLoNujyc9JmFn
n7kQbh9lHLycvCJ3LGBHKTjNo0BgkUmJlTMZC6TIOSK1XtMv4Ey5wbswU71z2kXr
uPAXVJzsM0SFgZB93n9Zk3Mu76M6D6jwpufrpzIuuamkJfEt7O51kJJXXganX4lp
yKq6KXpNPNRNFisEISSNr7p7o/97XTdvRzDKNu+0y17nLMOkqffnCFkOAo3aORWW
ZxOu0AC6sdFFILKL+qvSG5WgFRE5G+LtBWOmarmZDJ2sWon0c6PO4j/nX2UIPgzV
/n3EHuF+1c/yQSc0KankdMiCr+9N5EYMaF/Q3bbGZA0N/IkVkQHxOnldvxO7whP1
Vttk3gAyZ8EAoxUX50o2GY2AsVGlLh/Jy+nZZE8uKoEJQZvEJOLXNNQfmyCt+QVM
uVlvuzVdDbl4fncUsf+Yf3NXHCug7emGJ3tDdE1Mg4wwJc3zE8VsrCLtpEwBX8Av
W8LrEFfGL1p1myKhI1B1GIkr6MKUi/VnyWTqYhjbGuQpurynfgAA3QIKXqkp5NWX
4iK26Dx3vP2EGMJvNrmqGhxTUncd2S/s5uSKzhP28hkxDEHIKDtGLlj35DVM347U
rTekWkKoOteXig2Z8cUfLfMhna+I2hBD/lXsOKejHZL2LxKg92f05pnupbGvmTLG
d5R8eLT7HXkXAy5FUKPgibXuPb38ruC1D++6h3idyMFr7p0iSu6blx6k0aFm12Ma
k3H11rxGUOvypbXixuot0M+g1gh7BT//BxWX4Thg7xHZrq3i5GO7GqIqHC7GZ+64
8zb9yw6ftwZCiZgI1nx8h1gPsc0oHID0joRwBeGa4syLfsKwzS0oJeq2iRTtiHG3
1kCGKlfEi7rvIkdlwI5lB4D8dJJfDQ+1Sa98PO6GO7+z0lPu6EtAzgmAxUd3QKsy
jOfy3hBz98W5EgHrLPFc/8V6xN64k8qekMzNO0Dm1ZGpoS4PUZi7chAvHmrsTpJ6
CNjg44xvnzfSyj6j/dgUTngBO0AN8tjvnU4DZ/8uqhbm8D5lzo50FM4lAMH0D687
cxN2T92BY1yaAmmFH1cDu+P4lBPmNetUUCyDL8N5wrWGCYtgyzGZx2dwZb2dmJiF
loZm9ClvEbLbQDLoT5qgRsNfD6Ke/Zb/ig63lS+kzXuKjWQ4Lx7HtglVf2O5jjJ9
gfY//9DFjZJB+aDC1ONBlxnVqkMKs7lIJ7He2D7hFJ0YYvBoV/sYrURmGbLptcMk
8JXGS8BS5HnxPt/VJ8X1+POotsjhC9FbuiS+2uA6r1KI/vqPgUg97Ds++bMdCGRP
F8Wab5H5kocZLQCZmU829mTjDlnzenIC8l6SNIBQpQe/sVMlesK1oH5vpG2rXJbs
jH6J7/NP+TXO7/1GuMJbuYV1p5ec/98H0muSHrqADfQNeqj68MM/TXcB/opZZNxq
h5BdHzT4KID3yVNSZehjOm2n6w9kIOODFawWg3kjf4GO2qdDEvlnmKQCra2voDhR
pdbxBBpqm7UZXOw55E3ZCnF0Lg4epp8vaPnishWA/s00FH4UJz/z+wDynFxgRP4j
g9fkehZ2KK4cUtAoApuhUbB/+o/lNZEApyoGLjQrnF6P0ItfxXRmN/X1BPHNGWYQ
SSVWpLYhlMyokgfCTyZ43h5MlCY8+Xw6KRDVEq1cGkSD0mwufmFD8cdw/gqEzc59
pD9+E598xk66bmV1Jzoygq3ojPmLxa4+318RosgT3HO0WtMyXrM2jnx1tcoiboDg
MtcUF82KIU3LXejJj4O4fjyGXgI0IKUN3lV+2j+wPozn9v9CfYmNn4dOZFqZ72FM
6DvSAaOxrg1dppJzj2PW8E2L8vKas/Eh7CIjFutJRC7dZlDsQvTJR3402KQjLY3m
NsfzOi5wd38rVK/ibWgMf+EauVgP9PcbK2bMjB1I0LzwUzONe8EIThig4zsmXwy9
t2HT05kFEpr+q7fNAAUnvBm55h0M9VKt3PTknDGS/trPfmo6Q3Ryh9RpQ7rrxQfM
jQzyV1t534md1VIfBXuWO2phFfbwmrap3KyugenOv/5kDLeFACh1xGn859ddr5Ym
RtM/JpDG/ahaNqv5LJjt7df5emwrtPj7l02cAW1GKeCzuhfZY3M5kNYN5eBSaV5Y
+UZ5M8FkI0qGW8RvYJgsqsTu20a7gBWEmxR+6VNOukx/c55DyNqhQIFccvCxrdVj
13MEzgWy05ZszTY/sEgjm9BLNqi4Hq+qM+b406Ss0Kpx4qU29ie8+a32g5hS64jW
0jTAZyrd0D8GgG8eCNHTAakH+aQdVTdSMMAEEI5B+Fw9LDaHMBGwMpFZHDIRqbr1
KfC9Q6JN/RnMK3+F31snzcw2YmyRgGO5AvPVWq343tr/GK1xLa97pllcrgnUHCHL
z7jAXdRGv5oiRViFxQcg5UQs397rpe8UEUb0Dr6nfSAWvpt8kfyGql+RFAoxJ2N/
Kttb0FDykExGTDyjunWEg4u8/AWS9pv+OLgXw0NVbHvQZ47xeqVlaC/793CkslbP
qQyS6VyP7pBCB4KisbIdE+SEE00zb8IbqMqOO2IQv+BqX8Ts65pbU/H3MABzhWKb
kJAqGjyxep19wedvqG9brmFNtju9FFEJHj/tUhjwKJALAcMaAIYFQ+570fmo0Ehb
TGnNqa1a2QzhhnaX7ZA202DNeHxSj9sNiidlAZxfwIAMni+i81hxRvMtuXDhx9s5
rvJFZJDr7yPDyGIDpvB+HMWUCTJ4jjVL6x45vQemTSwooNCzdmxbqlUnJK9rAL2s
6CJ7izCUntWLhko7R9Zaz6X0u4Z+NpdJPz0ODrdMscT0ZpCjVOYe7KfuMw6kSkrw
eCvc2rQ1Utc5bOswN1B+TF4J3Xbv0obbDZ7ATBesdakiA1OA3VM+Mm0Zl7tOSeBD
sjGS3NejnVdb3L0MSlf72pq9YtPO8WUlktP0QQS7+Lruf3LPXV2yTFSJqei748rS
FvY6A0SU+QoOrfkqTX2+afIfqVE2wyCOqaem924mrHhu53wMfFKrsrY1HZw+/0u9
uNugZY/viypaBc3HIV+yteoPpUeRVHvOvsympPTelh+TQqIjkxZqGBoExL7iGIkk
U4m5IxPlXV507UnO1Wu8yuilKcqtNXj+KnUgdkqfLZSF3GhJ+GkAXd73C7t5nHiJ
RT7zxIedWJBWqItCHNAU2ofy4EahcUzlacg9atsxsbNk+70azOMNawWtLtqIIeYZ
RGIghdOmDe2OJX+kY8BSTD543WH4mwKkQu1FRDMANUWTUwP2/l8u0AwHlY4tRYDE
xv9OY79bBFxO7Agx5C5PW94u93pUGmUrqN+syYSfwg34JqbaadgxsijdbF+geVlE
9JFb7CKUIaOJyaum9gNPx7b/bX6Q9mz4ai1FUdtHucYnBAc28SnyNFRO/dMBJsWX
1694UqgEMxmgWiYAmqK1cNorgYRyCXjGlTfrw8JGAaD+YEQ2PTNZKBvZ9n/SEL2R
H5j1fWyORYRwEv3IxRwZExq11pZy/0KZLUDJHLO01VHRLY+4aDnHVYJZr+eVItPj
CyvW32168ks+3slceU/JiiG7CLKH8iq2yOxffQsNItiKMTeE5HTIpQD4NEecR/uo
T5wYZYfXLQ2jfXLUHtA2KkN9o/DzqKH8Q4esStittIHMlTEqB8FG1KWpcbD/zQgz
nZG3QYRGv7FpIlYP28iqOassZUZJNatkAtBMCa3gSkpMmFNNXg3OVSCpWRugKk7p
bMCzSU6SkSO/WX0DRRAQ6kWzNF+uE8N2ZYWStLzNBEpn8uNqKOLCHaRogU59Unq2
xkj5XYeVjTwhwhkVESnn/uvzHHBLLV4Z+ZLbAui6a8xplnRp/oVFHreI2aHTvCTD
mS8BGtVMS1vNfW3LDc3J0pv59bWMLGyfFodDArZJd/V+3a703zSa78FwzaVYtwi4
05mqSJjcfADa/VRGMvsrCwOdJpW/Bb1J2cUyBu0aipBmgIZM2t5X//VFyFvm9U1E
VjpNdFIiwrD6YiyrvBf9lcV6R1dLgb79NzkPN6PnU1ek1ofYsAahlY3DLdFddTNR
p64Q2sZfvOAhdgKk1qYnuM+OG96PQnrMo64ezq9KsV/gcuCvTx9nkgMu2srBiIRk
BzRb5UZaDxh3fFVTVgOAY99nZxbLAAmV4e2IbPhChuSA5f8KOrAxY9fCEtHS+Fxq
o76kKBfkzXDf38p1thJkn8tuM27BgrLb82LLwYX9b2vuw2/AsW+3hYqMmbTB7aPv
G+/zjRuMULlogitqB2hRBUGuxfuntyFszrbEP4SSYq3h//mJaQQ5UqIHQBSzCSHw
WDaX8LBhLv9mHgEEc5hqJJ/9g6vciFcK9m8ZWVjNawWZy6H5+c8d4YQ3305xt6i+
mr5+HaFzviwa6ArqrLfT3t4nYLCxDVtyTnrbsrUcFrvWdrf95yYm0EPTSmPDm5Ft
/UmVGVKEozE89zZ0wDIXaXlRZ1RXFAP5FpaCg7M0RpSUGnj38hAGK76PdeuwMU5C
YnZxGjcMV8g/Pf5Qg4XT/8mrWxnShvifgAxC2uiEc8g8UQZNSSXy6Ejw8INziU0o
Z/Ik+PwYeI0oElJ4G5UL64MCa8vJlcOIUVld5CwXT02pxMK7THx69t6PiQlPG8B4
ceHnD8FxwoGGagzqtA8TXTIwXwEyEUtSAhZFsngRYoz8hIx0FU7I70bRD4C4o5J1
9bTujx3ZWOQ36Fsd7BwYXe36YRLCCZsJD/v+d7ncFEMTBfSEAYG0GORD+Qlne4jZ
E/6ZPo+TFkdylMe3N0Pr93R5yueErxaDjNOp71zRC6ZFPNiDzw+qsTe9xL5rZRmd
v20VG/9C6mWkM7rxVmDbpxbNlCiZkwlLbSJMqJfXSNt3tIP+ji9jQgi/S3cQbj9y
9j64lsRhfZuRlPZv1IzTY1iKei5+6LqXK9D4HyyI3lEHjqTLf2Uhq/JFXIGwM/RN
VateJ+Q88T6+LKSlFGQLDjL7J0XoMw7+rsrVObWcCpVoA2feqqg8MJXZKjsLQRDm
zaC/2cVIX6XbfhhfT8CwZMPVzHLbqnCb8nyZBTPTavxpy/TovpgaB6R4P8BKD700
Eher4HZrnxAjEYJ/BOWG9t5fcNqp5nL6SyYbpKtLvj8RPJ332QMPBThbBJSm8Zl4
0THth0xKFyXp5QAapWghlFoymPmc9E55mBo9ph2NgYJJ/XV17qBTo1HMdZnwySVl
WmAnpvy6A1Ss0ZpkDg43W2/F8RtVosC58sN183mQUYA6/HtoXJRlunvkYPHjxl/X
gsWxQiFJsEhTNEMgS72/eroNhBNsilDhEhrqJFkrpR5VI5gDeU3OQCSoeqM9P8fn
E99fG1CBNMLcaHNKfMC7pFttY/TyaJfJG4Czax8zDeTKKX7soNZ67zqZGn0lBm/V
Bar4cYZ6qFktTF3ZRFXoCJE10rkmbuBHoKiZldsnz0dyzQwCQLoQ3zZerKh+PHRr
ZVHxuG2XvnPLpYRv75Vun501/BwPdm36YJBqgRZNuC2MTdRroy3VvfR7izn6jFzV
I430orV9Hja1mppubmIG8yfZiisE0yagHmT7k+DlldLZqw1AHSNG915NSy+ikxJw
xlgtlvf5TQ5cwQm0SPNaH6OelAAlimUs7a+kvfCE1/Du+PygeSc41qQ8jsTvdvDL
SepjjX0Aj25JQWlA0aIRBlwXUKYim7YJi49DVkjOlr3hCxro7DYx8kpOjGY5Y7Xy
4BnMdXgFssOA21JgXp4A3Qy+ywxGYdFPXjeCVG56oITDArKkKLa+bAIc7xbcMiSC
LdlpL20rBFN5OuvrraZT7Tx1SJHqQZ0n00HbxzfvufHDcC7wR2rXPV1u8s/wal74
uPoMEUu+PMCSYVnuh1Q22qFEMa7wMkVYe9zm+H7ryeR944mI4Wq5tjP6hUKMEuPQ
DxCldk0iJJo7lJZozTcxFY88tBB5mhmZXBqV8XssPO5ikAekhhth+1Pkjy/hx9mA
vBysNKAAplqhWjlGCQfWRFYd6BUruoq941SvaYyrouQC0Vy7v6roQ78WlQqbLf04
Cs6WTkBCtfMzAuJ4yf3kUXJk5OfE1yWn9Dig7HeW0ojuDhFmRC0SmlXo2WhJs0Wt
8mNo1xdOCFaFrmI/MB9Etr+qn1pEct9aZ505EntMNH0+j39O60yxr28ZmAk+8ulI
5k0r+rMF9SQ5DnIvSRs+IRbhKv7rQr8D2lSo+lCQP8sVJccL+GW067kCrsC3cnx/
GM8tBaRZHcCVNvYWBhHinPEsES7lgqp9rby8jeUH4Vw+VxJ8L9un6jHTKJjW0kqY
uVwmej0TwpRkPDP10l0Aau4zvBtErUEJJvobhW3ONDJuDoUyGfGk2Qy/jdUanmuu
yYZ540ZEg4QwhhPmUKeii1uEGlgLeCDUb8ymf9Jz3hl4gTAfn5cBpheBpEjgvyqU
fUrhoKKjuOGJWWMRIgCgbfxHHAX0l9P6vvC/r1cvuDLyXCkTCarMEsAE4xMuzWNr
rOCbO1QTNo9vsnMqfX0ziacdpfCcBSO1ia/tk9BSu/VsmKASEKE+vFzqOpV33/RA
2zuWgqldTZPZbtup6r3PhGxdvev2VMa/lumzQg/L/n3NQg5u7fCifBg/wiUR+OyB
o3dRCO1CUsRMAfzv4naZxcGkd9quBbmcuxhB4CJVCmVJD0Pre0e0cczC//51O1/S
mLvFld2l/DiNm71dsFogspoWR3qP0ndzboR8yAoKtSEMJMHD4cFDsT1WT5UyjP0t
KXYCCUcxIluJl8CFTWQREnhsGGb5BY522iHPI4gdoK5iiufPie4SScnsc+HvtwH7
7rxVTRcZzvt8J3AbZb4Skj9OUsdyaolyn2wI8bgsqiU45gaq3akIuxOjm4YRyPDb
3TywPPzBJ+Q7w95QZVD0wKAtiF0eD7TnuMl8li/k2XbNk7Mb7ukEwzsNzUPLIiQy
+ai4uxSN3CmtDwwkUUoag5nysEx+yqSHGlvvi23a2PAcJtm15+rpkJR+2zIWajPo
xt3mMt9+ZTGZ9sp34A7YxXvu/JafkOTNLkizDnu4nfIqCjG6mOlnTj2KLzUV1rtL
+1Sjbli2z6psJh0+qZaSrbFxwqGqq5Z9FWKmKJFP8kIXo60+P/4Mgxoq8iLSfuhN
0UyUI1uYahlLXlpftb/+JpD1zR1Fjd2dH7+N+jKcCUPxW7vRnYmRCHDUYjyeaoPJ
MhpDdHOUz5mtxDb3XT8UCSooquk9x4pfmPeECZr8yKOkukq4atFSkEAQFvlaQM4t
SBDfZ1sV55q+q3B9dnzSEMmQwduQ5kk8dXfTerQoh91qCrtAg1lPL7lu6Dy2jDB2
eIQ+6eF+A+ONvYIm/wdRvPYuFrxVAsM1IIKW9r0nGorXOkqrMnaXpCLzrsMCl9P6
CUEgj2yDQmQnw+bNFuAklJLllXUCcgF3j8UoTAVfTIkHENEnDRFEzcHTUo6BbCMx
P2ScJM9BecOfWLLGuN5y2hliq47ShqrD/sVOCVBvbYpWH0FlQN7UBHgS2eFSN89O
WWidGhW2a7XJ6qnJjBWQERFyMvS8Wr27cyJVDuWjpbUzbFRboiik/U2v0lTeug9S
xnODd5j/F2NuikMT9DS3UQaTDKglFH6sUg+1xRHPgINPK7KYMHitzb5cKzFlfUdk
wDGEtT4z+K7kKQ25aFRd3wbOScaIgQA8P5teRiGG4KpwT5STc+FnHV5GzJc4sjxD
OSnyAAG/N6G5dBiCFmKXziM/hneDEe9iLntYPpVHlNZQuhF/7WEAVovXtmwSbhdI
UZNjYQWWgUgqpiDBN5LkHneqXpxuSTZ/UMwomI5mfjBwX0ipH4rTl0X661X9j2cr
T78Y4NNc3Enut+A3HQmL2jb0ymMIvSBprL63vVcgeUttezBW8gTH+vZQqQVod+Xk
4PMhfX1kcGWg2c5jb2uiUYj2mJ2iU265HJ8cZM6uEpS1zKyzNuEgsD60VAVTW5Ax
Pa3veH2J9h6fmtnA0ZdYkFcj1LcC9ed7Y+i35giz/bIL6EtUYBO1otul792dCrv/
58NbYYFKbZLwmVR7O17mh184Vdyip67aYXb677pHw5PadT/vhqQMG9/Lqj3g+ylf
BcJOJdWgQE2Kcgap/4kMJwui87gECNg8OI1BxuBXIMo3qknileH01a4klTCGWASy
aXKMprreEHK6VyorErArVD7IRcTNBik5O/yJu+Fyf5Z6QU3tJo2E5cst56NCabXr
jc3y9cAhxiS2oTmrihDhaQHi2zlloXYgM6Xs8jP91J0hl7MIxoZdaUPuJz3HTIAQ
6J+dLFeCsRhew6dQPhxm3PdlAOXkCyP75aXFjx0RNBxZxjK509apneWrLSzh5q4P
6lZt7v+Wa3DGLs9rLorNoV4znJXc7YUrWc7YVwbkdh1qLQfUPsaTN6h/qGtrgV5n
90UbqiJm16HUQD0kmyh9GmAO6KvCWH08c4+KDuHjDnK8/FAZcbdQ/CyVi/CmO0YR
dU8PwP2W2r6AX8vHiWZuknbUMHylrDt4T96FQzGCvbS9IeroFE9HBS2h4nBNKTRR
Fj2wJlpIQj9/F8P/DkjnncZAzvK7P18guuk2DbNtvxDu+FEcjwPVOpU0j/YBloLL
Acy2Xe6uP28iULV7oL7jBksS1X93K86SjoCmcOp+RjQVD/BN22u+0a8eY6/YH5NZ
oIIyHbsjfLJzya00GUMglEcxm1rXHWidlfPVOdHAwmwgFhonubzN2ku4LECeqDNq
O3883q/lRws7ZQwjEWd5hxEk3oy3gNBfBk5+xGRtwBew+3g6CWO0qXRfe4TZjeq6
iU+Ao3Pgh9I8rrIV/0uyXKElEtR/XsYqCsOsBEBfKyAh0R458ZFNR6wxG6pnMNxC
JRAoSxxlpXliHtjka2BbVQICvfPuGPYsatmQSrmajexFofAjxljiQ42KbTqd31k9
t+b3V6xjm3Rtnih14g2Hf3q4PQkcqiP7YChq7iAKl4dlLyq9VnXy7gaT0CZq9Z6G
J1g3QEhue4yeUH0P8H5fH3x4YZzjCxu2+693gGDegBsk0biplxbMIDhdNAs7q8Rn
RgbR1JeDpJjlV0SeHbYbUQjvYatDrxHorJXlZSGfQrhUfBP26kNKW708a3fXflmY
QKF4zlsSkpb0PObYo8mSVmkH9aklZ1nYuHfjaHmZEcJ9faEdnNtCu1ZxsyKHuF7p
E1hYBSJZptO9ys6TW4wcXDYD2cLFH1LobGWxT4ZkSx0GPYYxzZcLLDyJreD/bSEw
HSohzdYyd7ISU1cPRFNEgKdGRzqtsNXuqfdNWSayTID71lJFvqVeEEx96YPtImJP
k3vLxCrEOC8fvGKKg6ilLUHNcFaYHi6+Dy3JPvP7RWC1nK+Jl/FouvQve274eqVX
uDQmNJPDGWYMtX30pu6bsnlivSf2PcJIrvf8s3BjTSZCgU7yKCSFkY2IQHdM3ziY
mCy8kF/TL+iA9yf0opzXFagO+ip96k6fzwM36y0uuXo8KviBrgWaepZgNBM5Ri7E
qb+nwyHGhsyPevHzFNgNHkSsu0yQD9zA6qpEB2DLTFyLgyrYGW1CJg5PKPdmnlWJ
rGqZqo18JC0ElUFktyLA6rYBn4tuekTGLiXW9FAzNkr/RaTITyWTtsaFn0gQxDVV
OKnGMgI398ciNES2j7ZWsJsSYVNuW64oB1OsTjfLeV4xzoXuwPltFc+BReKLaAfL
yRAAJZmGI0QAI+7jObTASD7rDlDUobfWDlYzp7Wc5pQeVPI4zwaUqMGanxDEyqPW
2TUQ97vG1fbmt/0AQ43X1vSC9OyThP9SrjV+Iy49dbbG4eRHirj9PHee0hYb0v6U
3raZ7oA0hm+XNFoCdrWC0YX17L/xOIx71FzyfDEkCBtfiy9b2v1SaPu9WLAEOPv+
eJiexl/Gy2htqs1UcDDgrZTZ5n/klpsZJUm439xA/Ofj85Hfqh5WIdxFDGIYkmXw
Lg2Omo+B+VtYaNi6fYWo2PFXcEs5av9lyT8B9RwNMMNvjgn16xs41+8optFJ3SBX
jQ06l8aEB82PpTLzjM4OwMNcTYHyyO4t19AnTLd5BJg+zQCT3XRCOucHUhVy4yKk
O4Baae2tYTBWRWNIycKd7uJahAQGfzz54ohxvEMhnRu/AF6t6GIFM2UiuriC1NpR
tiyNvGTqLbAzEC4eEA08gvsbKGg9Ou1aDxe8g0/d+pIIo/FwBLULLMk5CzvvITfF
GF0tadnfgmantp7xfAfs3/wxm2iFOU9CfolBLzXhYp9STmuHNO5CQYwaWOWdQJ+N
Yyxxuh6+Jzn8sPXp2IpeChAa8+bk+aA8RYP6gWT3AE9zUls9dzPG80DfY9sK7B8c
Zz8AzxnKtfliDBpJxOK1az2Y3VfbQMexjaJehYpqtxqmpkhVtqEkKB8cAoLbWQLh
LQ7FzZv1iX0DzJ+U+Y0j0LofAwrwQcUOmD0Z6H07a++V4C9c81qWcnzCOU65RjXo
LiUaqjW7L52ZkNHRLenKaXGd6PXVtLMufvNddqoWJ5Sw5p9xfNHyJB64XnS1y3+m
1jJrvHF2iVU9vyjNTSx1V1bJfpNJGOrCkio0GoUKsp0UgwlQs3Jwz0uaG3/MbWi4
vTYO0jFAh9o7g9LFkXgj1NXD3iNd/uApfRslyuFMf+7gnMfV/2tmc53IzOlsipb4
czava0ciQsXhxaKWmdbvPT8e6Au2MAGgb4bA6x7Qtbw76phUNbdwu53H8GwnFg6+
wDN0FmJ4JSXfqNvMOu1LWGjWLas+Vww2Feyfy883XBHObGZWwXX3f1CyyfBc8z8z
kHJW+h1yrpitMZqD6w96y1CJekgnilB6xmkr5cAtK27sAYvK2cZ5i6xSGjfro7jb
RAYddDRrBICcS9y/lrlwEzvQ4hCw5TsS3r3INyn5CZ4W4j0/7v74yTNhU4kyiSsO
jhlnj3ZsMsONI1CRNOwzi8ABfYzIYpLZDIW3Lv393bwenb8Nq7F6f2tzM9Kgrdv7
oX//JVyRUsfzQ9wz6bc9Yxq6jZy+o/1sBTCaIi4IDPOM9GgJuyKXBG2CCldoU6If
BJEC2PJVY5/9ZyivJqkNvJ/cwB0TCSXcXzANKG9beZpKI30IbISv/SZefdrR1jmO
iNFxqbqQuq65/4BhX+hewh9QvCW5zwaIk1zEQ8Lh+389AvHO3o09tWzbQ6tgGEIp
Nqdnuq4hRJI/L5Jkqif6+vmH9r2xdvU/t8IooARNo8FkEnwEBlQ77NON8cM55gyl
+/YKNpTRSlBTiYug3UiPx/YY8pZBIHpmyrDnq/Ae0stoKiW1ms9o4OSit1p5f6s4
mL32SDBuKV8DDjR7YyQ87eYj4cNb1I1cg9ZnIknhdsCDDD3VW4mKDBHwo0QrJrKB
6f6PBEK61pqmd/AnnMsmBbyutRUPPb/8IHUkFzjDntxDfbhg1d5upTdFwIWcep2Y
jnygWusNPGmZu0zEg2g8C2Y51RqKfadhlm8q2Das3YwO0nJlPZUF8dp04a/HpTHF
u175WCo1xZiuxIP+lpQAkgO0MiwxlyFQwWJSilRAsj369kCX1cUSb1E1AOgXmgQa
o/d1/ivpH1kARUZ/wSf4d6yneKIcSjSeJWrjpWI9wYXsGk0lL/itplCgAVfQw4fT
ch62Qlt4NeIPbdnqMfFctZLVibAAN0IVYNQfwxdOa3cFSdKk9NdGC66rw7aQkWcN
nxttqjClBZnKAb84nM8L+4EzGOz74ABzS8f+/u7/rm+ppwGDWBYhmTG6mevW2q8g
hd+hA0WzbpE8VUbCJLZsL9cSJy0a0jI3+1BnWwrA13hRNtgzaIaa/DWMkknU3/jf
g4YdMH9G87JnUh2O6vlB26shl4R9vJfjWm/XYzTHN08IKe4kFZa9w72LCN246HHY
cpMA31vtJueWms75QdnRUItw2UTdh9ZWpNFipnn4d0wLpp8UwOqUn1Q4gWjr7OqQ
0uA+hLwFBEN4NOCQLdC8unXEbITUuZ9PqaZBy1stW7b4lYJkKXhhQDvDR6cikcGu
8lQxd8rhvWptMgQdsU4VMs93o5B8ubaHDhV61v+LVx1PlSCC5IdVNf5k3wRZRblZ
sl9wzx1ZF0kfRd9ziW0NfE6jZiEsdQf2WWSYHsAjqElJOcvXc+cwSRkal85GJbgn
Bpes9gqbctka2TWQYHkcr66w7971P3YmpRme0RYH5hYHIgTl8PgcSLvvJNpse9eE
WBhDgFBt7XW8bheXG9i9Ajtzoc8X3Z4fVBU+Pp06XQVwwTm4mJjDiZimBZb+wRyL
pCZWw4atWGSp3aIOrwIgkrYFKx7igBMjqxGjecJPlch3lJGDm18RSM3fml9kUX4l
VfnBWhbk3KUqQLF27YpGJCLfs00Ux7LPcYmccUaE18izjAp0xwIp2XdkXW+GfX5y
6PqnWQvijbgb7zYGIK29N4IwyPbF45fncgNKi1g5bJSxqvaIyVVO0tdFk2zb3Qys
OOC99ACAG0Or8iHJDiX9K/J9DVRXc1+AG6xgYatv5Zuiqj1p09w9IY43LZ84s2xp
l7ujahab2UKaLf3K8d8Ru/L4JQWY8bsbr/tVl+3A1rJcGtWnxT0Zwm96t4f3NHAN
MyTf8SEjuHdhJcdK5moLY0QyS1ZDGA3eTEIpzGzSILU0glqAT761VZXoFvbG2Abd
0Jf1c1gcrxh42kxOxViZ1e+UYTLm6NtWZOVesv3dX0J7wEhuGdaGEXuqxxK/Ztso
LoX1jOZvjKuQxTQYUNqiIlQ76lltBp/lldljoETHBgyaF7nDNUXyibI9RPUNUYPR
vGv/gpMUaK5WHdCXTbQKeYQgS+Of3JkRkaQs4QYGIkuVeCxbtA1CTarEaQLN7FZT
UgH7UI0fBU9vr7NsO77gpwYvnv6ekCHlxusBYh/c7rwa7c+DL9SsrhoJgr8Gkb9w
LzlhtOme67+UyI7wA48r4jn4i0T9DTrSMFLnLOku+AOaasAyjk1NbPKSGmd1hbKJ
q73s0nlzRv6jdCePtk88B1qR5Mier9LEqs742TuQNf86Vk0GNwZDzIhv/Ob6okUC
CUi015pSiz6c8Hjug0/uG441IfovPSbpZ5ZdrpAjQxtwkFmxJhmpxTKAvtGKptyj
Li1WhtOmVCGcqYGkjvUlpmQxQmxIgaV7UARgkyv/e9+XoGBXS1qTTNcBIQXuBNFj
AFVMaJhckzRgxbjSg3B8XvCQ0O1LryfZFv+UrldntmFkwd8PdxtozGmIFeZjpBE6
qKxFgdyRNo1h4l9smySpwdFZ8+ewdKgY4uEnVjmHe0ZSR7aeV7GJqunGSXnPqCtV
MGJKM7tLi76ZGt1GKRVkq6rThfc7RecB6NAYNzQp9Ni3xTPC42X+UthSSnn2v7Mm
0FtYXsI0xi5P+XPSDzOfHOLV9t6TPaJC8/oDZTMvxXENVDg4CokG5RQWs75t7tKt
fE2FwMJPR469ngbfE1Su2mKT2RyygePD3WIXx9XKSHtp7Ipr2d6UqiIf1FJqbL6M
jvAfLOD8CC/JAhbesRgClwDBJB35hP4uQkHRjsBZHEN8MubsiKVAMuHKyePDP9re
acVX44DUw2rmJUpa0WJE8ybQKajQlltxccRxZFe5gMFmibWY4zGNLvo6DrFBxvmc
XOA5B1pjQPEpiAW3Mldl0do6hCl17zuLZBqoj9wrY7wfNaZFZ+TrnSztDn6AYdSX
haM3QwTr9WuVxV1aTvx5IEG6tFAGcRD9NQX+6d6nTWHh1nmWzGGwRwz8zvc2/i9t
iZyVUULT6BAzSyefNkRn11o0ij1OHWIF2R0l8MnW4joGIPyfg+D3p0WQA2DloBYo
GSnaIG9Z9II90hyQedf0TdCWsQ5SXHjGRPjJcDHQbvCYpWfrTYvAVekjqImW5awb
RKOjp4QcR/L/6edITB+zfgXtDNHceyq3lk3k9JSv10AK/M00CLpdz5TVRiPUjMiY
sJmbgUxLWhOjqTsQhSz2nZQ/mHvG3Z/sTY1LedGjLw7av5te+0tKfxnr1bPXberq
iCe4E+9T85EVWtnYr1bCROjz3qAbHAmFLHrWGgZ9F2wEiHiWTnRq4M2I3qIuq/ri
+KNU5dxTMJycD7HIodUC7Dpo/SEx4pVmgyKd43x8Qg+FLB8CY6i7Uk2Zo+BhGTGJ
Bz2/IExt7AuVhg2UkifvCZc0JA3gz7LYZ0t7kePFRwcdF3OzZsdQU7Bl7AxMvvo1
PaAjCZX2T/PZ73vc2a7ER/ljegK3RBhKd1bK9w0dHZ3E861Takq6qnnRlOhf/uon
k29tmoqYpw9L1NX+RiWomntGrZb5CHfJDMgfbgx5W8dhEEM7XVCafNDIOvX3jD5N
INs49+Y9DgoZ4Xl4F9+0Xu9D/JGB8v7rK3QFcQyr0DljDWv/ttlILbQaZJds9nyC
E4SKAWAptjOPZQuiLs9pNsen7atfP2RpTKrdkq722/RSkyKxQE2lccYI9zI2bAvK
/i9Tc1yWW40RSBvATrhYu9TTS4gV3fkyL8VdoxCbK6/L90c9AR+rj8tewXfy3S9M
piK6ueaXRFT9WFB1Bp7rAlpU+m2JAT9XTc94hcr6/SNYJGMd1zMCTzzqRM21MgHD
WJY+0Wo7IpWxxNp5NPzAKBnqlDf7GPC9WUi7C0yTZwdvXpA1ysqA3NKBD+4yvAiw
hl08sILfCes1GnAwoP2q3BV2wFEkOKwv1ccYrjpfblkXr8VsIqP5kkaieDFWntTV
V7RJPeRDmq8bdM86xux/d1mXoICYQ2UlQKXKV4h6NzhlQK/a2ROUIN+eJjEb3xJD
tOeuBq4psKlUdlHWQsbHfZkoNZesMqj2+Yq5YQyK6H7qBdLwuk56suWBO5A1pwgg
0iLJTbH8mwn9nvBNMCA3+NDsW7fn0IA3DVJU9W5xNhUcAwOq7zlvWXr8OrcAfpGP
T5daDIfozzYOXfgrV3Ujn3VCA/PrNtC2DhMmCwAkBPHI/S1Ya0LNji2cqo/zfdLW
y0pznmMloVX5Yel4AJfoGwqQKnCvwDh5TTWL+8K0v3ZSBxUkltw4N3txEvnmXRza
VFsHaHVeIGCDrvvtbp9IVe+KapVpZuiE3GwsLNOSURxhNFR2Bznw00M0UHgC9Mk6
v1LYLOB45ySOOggbh6bEhdsj97iHsxCSQM2leTq+HEnaqZpWoDTzDE0NnepVyCJX
NkuD7SG/FrVfkvwZyHijDT2Lh8fPjrRNsWdfav+EEcOb5s7o7cQNFLyjBOj/zv2Z
qwT5vDDcdQHRuB4V9rx8Ks3YmjBBjGuZ2WdAUBNmhwQ/++xI6fwbqW32F/EWMGGd
hs0rdiGwJec6knhGjQCmTWPC5vXX+gnvgfg+0IJzAIG6PRgeUY8o3Ro+KcWEmQYM
t/snOxDwwLYpWYdNKvIM9VweVHVNNVpxs+etwrGYrx1vHc4C+DTPtwMwDqzn5N0a
9jkyW4XAQWuSJtjlfU3IQ7IUp0N662zSzesKpVeMYuJ4AsMaRG9R4ru1IXGoAq/r
jj1L7THIxWx2go59esX6Sc8n65GH6ZOm1hTVH9svbu1ayNhcZRGoQM/bPW7Xz5L2
gcZ+DYxnJQx4tXP673cX0yR8e0kt6MnNZD1sCOdFCpAkl5/zM6z0yJRUqqzORw8F
95APNzWPEIuO1G/JeiKQTrKUz5vLXO+4SkGKZUr4pPf0Hu6PsdHdz+fMCZg7H2f8
sUn4QKYKO7PQMJkWQybmVRe7nAxWj5orRSKp+wTr7XxpfNL91w1497x/ps5lv2ap
HHPpdNhAmvAYCG5a9Ss4rWX7M7MLOFzh/l7gBnOWwkYm+FohoitXX8BGpmBYV5Pd
ythdMJhgZNH4NhwNUeTOEvRxwjtjwemQ09ARaTVaZC8rNCE4KiXFXioemYOXyH27
gKsyR+uDW3PH521h9RXU6OkiDiHEVbIEs21CsUtHoX/bJ+IKvdTlXiWIJJ22ST03
UTARDGbTsUM/Pr5XyQIAB4lcUhjj9wzRC1srqF979lYfEGnmBLz0cvUq3giCxzCo
5WlSZ9HTmHu+n+ja24W712fdPZyc7X6l3aI8z98vaq1iPz8CDHBWHwJaSeVybg9N
KblzXjs7M2FcjfkiL6cuQ30cgv8AnLgVqt2E3B6IaWon0c0SqrgFvy7IA4FTEGsj
O7GCH80zF/Qn0i0vd9gnVVZRDJF2G/KUWBkKMQtjzi1a9w7x/aDEVlCGG+UL2ggH
sMeeqw85zULt6RVlXA3/LsEoJfA+k0BFKVEKeUIGM8txH8Aj7as7uLF+qlCfoVXx
EC79M2AKJAft9EhSLhhXc+JhZAxNT0E977hjZELVQ+rPOA8gNpkC5BGmRDW65+ql
1EYKkp78M16OQjVajMt+UaitXyIchpY+mZGm3UsNnqflNi/orGBeKyxXIZVz+saJ
AIKptQmuz9d00hHex1aztiOkMJVEHQBGKGtnJzLQtXxvIADEd+Hm1Aqg1IbJTg5I
NYbpUbXCkOZfuWbyQ8RIxtXM39re5C6Cp56f6+ocXwG9mrR7IAvL2akagttB5Pox
hDWR/gKNKNCZnh/Nxlv/+c+R2vJXwg+Igmg2voU9TT7Ts1cpbc8NevEcwOB+RXC9
rE4x9MCJ26XpyyzrRSZtqQJnhE0eSx7F0ppOupQJUVs8C9Rm8JVMt+bXjmW2X0vu
Xqzfiw5XTCCxFIW1IPwY0kWA6b5RQ1Q5T9NrmcvJm8WlILnAjbaj97k39KAuuvWK
QgB+Cd8WdksVbrWk8DjQ92b6TaT1ituk+TImU9CraBEOiR6hpp4G2dKcxjCLD6qJ
onwBLCPx+73z0Rzo7zxPbq0KWzfis8NwPz7m6qnm5aTQBNB4rJODjJOiPmMxgJ1O
8qS3C/UUOkD0m3NpPkK+WY3RVpHRK13ucky/GMKk5fuKgYesczOkeAtkNiOWcrxX
F+scf8N+r8L/y95+KifXkB3pGwJHfNWCFVclJMqvk7DGumMtTGcZ1mxyXCCpbMjm
PWvIlDQPW9YdDFO4B6ptLlu+7ypVw7clhP4eR7YFswr8ZtaNGw54vPQqxl2kwIT7
RtRI62OzUhbbZhmY07OC0wjVTAZ/0GXKNWfSAwxMz+SBOk7z8RxVyVu/CoFO2sGN
xYuEgrZ8Hp3wSwSN3Gaq/dwYeg0absh8ToByWye4JVxGalFMB0jY1vwX4tnJTcQC
Xlrttfo+tOShGOz2M9E3a4QJkvhL3K2wl8Nsa9EzDFcuND1/oqUw6n5ubxjBfW1E
pOCcm4AT8gsi3KZgubyacMZEpsl5GQ18tLQdcS83+RUcmaaLuXPMeLBIqZ6ePRvD
JZUT2gggS63soKuRUEVNe9q/ASRDxvCdUR2nzOKF7g8tCNmtcQVhClIYincFlNQc
bAbCGNVE+wZHPzuhyrhag4MJOCOYkh6FVx8XrhF2rmbLtNfo+GJ5g6BT7cdRK+WB
HWzwg/N5IxQgi+zMsYtQQATp8o0FT5rFcg+ukrYSNlI3OdHzkp3Y8x761hZT36f2
ueh5+ZaJLjl+mDNu2+kNi/D6oh0ylNISEz8+ME0QPAz1RsTNEmd0p5W9bihq56B4
C0KriNRqex8fGk13Hysr3VeChjukGtn+EsOl9QM1K/as0K1UU/mJIqkwpfn4rKWM
hfz9R8+gx/lXwFdSOdCxEI4TlHooo1/FdcsRgqU2ARVGiG9yfHNQpM5qLmiwDbVM
Hh4wJX/+6dll/ZQnBbyZLpQ5l8PufFtyVcJ0Ls8UOFl4fWHyLQgZVVtETOKSZPi2
fsjY2YYtd6uND9H5uZPvESt8G8WtoOXd2ckCaSDga6ZMWsHBisHZYOCJd/FJlnK+
MbKRkW4u0rR3QI/eKm9QXcetmITovR15Fhs0VmU9JJk1mUwkl2Wz2oE/hRpTVbJD
gFy1PhN3nVwHi5KjZjchicKtbUu9Bhom/ZyKHO1SUUWkdJ4VnkKE0APQnatp2jGp
Gh6/o/Q+dtzhj8GhwMoctu5gYSRIWeKh/5gK08Ub3wt3OXSsgFU4yj66f/D8n7LQ
N7EoY9ot66orqn6awrvs8H77pwXDiRON2VQM1r7QA9oz3RnW+0kFOoVdn7h5uTed
vekG8liVv+nQ80z/ubdhJJrouIi+dmyUL46b4BR4k5Ln6RzQuvh82TzmtV2pRvfH
5LnnWL9fBrIlAK2uueNa6+frz1dA5qE03Pgzs01dtWuTUrQf/9yYb8RUpmYRBUoM
IlMIceIRq10GOpt04Wn4kwtA/7AINIrcyPzsZpdfInOtlf2uHC/hxDZ3PqEDbW2P
qZfEKGQfy8Aeo2fnoHGO6g0jnyf+TIjO7jnQyFizLL1VSXR3caqQNZXdT73/w4GM
clw/wFZaQIMrBM4ukdG59WucubpSJ9MohNv5FPT+I3YsW5KfnYcAK/x4558rNIwN
SHvbEG46vSe0Y/V3f3l5p4sl+RbsmwpxmASdmyZhUU5jTd3WeIvd5Za09ITKGNAf
rbU7AeswlvK4OYoYU5WslLuQ9xhok6hpztFVZgQAZDGV/DE5Nhtb6pEt+pfxhOfx
66W0Rt+Yi2rlBLgxV7b0bkBte5sBkg8/yBS4BRBppd2uCuVJ5po/uIXEWpldokBH
Lp32VGF3b0cd5XECnr0b+pUYUKkyeo5tm8TKDlkmU8XEtvoE6SL2hKAJvJ+7qfp0
lZPlfTXzMAc918+16R71vOfkFlS7TmyX55Oh5uNC2Y4sNEoo2yuJr/cBzz8eUuS6
dO+OKr9lhlfel0Nd8Hk538Y4PEzN5lNb0oLl7YrTfNGHp8/xnVBhLwTGAKyzoQjv
Y5x6Emwg+7Hs5IbaEvykScVuPTSJS+93u4BtNlkb8ZQcFLcEb0mfcQdaT+a/4dxf
DIZCjIJf71/pWoBpB/QvJMXaD4QB3NxU3aXrPwYSZ2jFPn4LJ3QOsIDSzwPyQ1Dx
ewSM7DPfcpgUz8H8w1/ZkIVCEc0S9gg35hdMIjQpYKFzu0UWlLa5BrNsDDVcF2/s
WH1KunplyexHZmWFz+Oh9YeMHKMwy9qWARrBxAKCzJBtsguv7e94CxEDiJxg8s73
MhXWG4dnNBqHcsHJ8D6uiBaqBJ2FjXjaMJ1FrIpIOuJG687XAUOP7ud3OJz9i8Ee
x1Ra+X+3xNM1cSIa+F8g2G8geNaqcyJZhcNe6ZVbKMLrozofV2Qn0qDkgqXPIITP
2LvobytMZ2JDzPR4E3/p2JB7tbm9SVCVyBofBE8uwesVBNqqfj9I/e7FnL3JHsUc
AuzK4wUf4zy2bhsBs/xI+jnaSex2jYIzpqWSrbq28ZS/gUhDvEQRH1JncxWIWKu3
AiOYzbbfmH/PxuaJ9XStUZK+ICKFb01ho4XPF//M/m0dUXy2HrzIDabmeYJlbBry
hv3bQnh8DuQz1pC9ROdsQTP2vNVSRuRftCOrxLXTOx9OvLK4tKGbQhDoGKsk665r
lrpJV0pnvYT5x5jBp531LxbbZEuJjpgh4Oj0mTVE9VU1K8EOInUAqx+YOzqCTvKN
2U0X++CZPp2ZhwW6WWA0GNOYbOWyNO54zN2tGJtZaGaBzswGDUMOgJqCCeKz095/
s+3lRtlQRRUuXpAt//3rtJSiG041uu2UjJGlI5YONpA5bIoWiRMBD12mhLACM7fW
+vWq/5I+vlZOIkhW/ojkaaHC++HV1J7Pa8yYcLNA7R/Hxo9/aOT8y5pP+6qPMjaW
pzwawyaz4mY4MbW2uKYT+Htbpo3JkKa76r8vhpgnJpYjBjhch22cvKWpQocNqhWc
/C6skEetYB40FWCxRo0fuyvaZS4fwITnAN+xoNGAtVIyxe+UF38sEKqeDkv+yoFv
7AO5hWI+nYxithGOm85jy5aXfIClh5GwlaoknvX1AqAX91ZqkK7wHBsHegstuD+Z
8JIbO59rH1Ckh22kL7FRouWHJxlhV/vPe5yiDI/9JU1DOftYe7lmy11/fo0K8/V0
2EIdwO8K6+HZO3BE3RHKE2SdpyHIAQ7fmoVne8hn/Sfj0fgwhcwHH+Q1daV2+7jj
C2iLm2n3iGPv+/Yb8Li1HBIrhQJ9+v2C+HW5iC6frAN4EwBQtHK2z1kGaXJBKJ23
We/CJF6/gAQAmy2oMB9UuhVzAVQRRYfl0h8x65s2Potps+oP1nPIHShYLldO35pt
+1petN2ewuBJFvYSd+QCC+zyYS2cwNkqY4JzF3KMvI3H4TrbmP+poJgPDD6rfLW5
V0maTV+6cDRCOrorO/guivnuiOoJQniOHLNU8Q/rNTejQGYEN7J5t74z32Q29yYJ
EpjU7KoKCZX6icGfqQ8u5Qi9L7CxtvG130ewsX0VG5J7itLvwk66kdbPq1UgMbMX
yAsHbFhIz/WSeYghLcK+Jms4JomLsJQtShxFMC+58M92cL5t18Ky3h2ePdRorUUQ
9rLiUz5DIDxoMkQBEh6oBtvs+7Km+yXJa4Q5V35sGQS7QhabDoIGNhPgtF7Eh5+v
BhwXeYqZdbqcDEkV5wTxFAXXWhteaxiTzux3eMRMpTYBwNNWyKDTUuGKLEiU/fTJ
3mzPMGWHzQ3xaE7p/Ic65jgqnf5715esdcl0lXSJJPJWFnSAqyFvaWntrbpodbUX
WbsQKCC2z6hRdjWSMXcGdPffmE+Ccu4OMx1fYip4cOp1Om0E/Ldr959hoZMu5pH7
wbTw/3rnh/bBNQSKX4in6Aw4iYRtgIZ/sjkThj1RsDVrQOkc84yEUiTZ9QfwylA7
inOOrER5yWDhPjMJG7T+lAUGnRA6XJ8BeCbJA+Q2+9xaip4sJ5qNks0vHv2IJ1dK
MGojikzO/46abTFMFw5vkK65eI7s7BgrldhDFPVp+BB7BCoxYl+4ZvXq6y2y4ta4
q/5ZhdcQSoIC84mdrLCfpQIFvWRjY4GKfeFy95SOVG/XX6IkCFbp8iApPldP61k4
C0JQi9IX4AoGF/SAt39/0NP0NP3w1Z/K0lJZkqijOb1p+oBYPazQ0Or54ta5Z5PA
0GUFZNyiXxCdTkbh0ePz2aULev+HX2lzC33mYs8jXuwvqpvQejshYz5UrYm6Z9Uy
8BUtGYaRk+/FN+VWV0X4h2ljK7gZCExICmOyjsYJsoFvJNPVR7iB8B5Nqp8e4R0s
6zwVWVDuW0lE9ev5jOsGVEVUdadwB3VeOHB0xVzNLH+MBfQqwsomjwf5WveR+58w
NcODWwhvSI0AfWWm5hlYncFJSTyhPxKG0UVV8O6S1RDzMSYKSIXZgVWusF6HeJW+
QuaSwID0o+aKy4RSBpRQtoUMhUYOHDWIWplp9Kwpxnrqq2w9JUSeava8upgZOJwV
lA6wZtasullW3v8WMbi7GudFcBXHi6gI6/sIpqa/B2OHJK8smk2BR9U9nZ9r1h+t
JNE0k3IfuPEWbzIhQNa5zXXHvlZGipA5ArIOhXRGQsZPHYAKk5rZXDTGd6LNETkf
Yuj0rEpifikTFrrmNS/pt8hbwMAD51Tv2GtQV1ggnUzQTi2ux3gprUyH9qSxh3Kn
fIm4N8B+rinmVNeCb5IxaDMdWdpwzaa8lsA/lSb5Jzudes6PRHoFyCh9duefYQnf
mDO60vtb2AmrcAbhMEp7m3HDcwNEve/OxjAxG3A9Nv5+2N87ZvVi2YjNXnflkGhN
ZYkBjdTWHtfYhJ86i538XTuYCMmMGfrEJ+wMx7QMcW8yNWBw2cOARL3GGSylsciS
scy/ZT/DO6M3JKlLz6avdl2EHKnjBekLwCmAh20P58ca2O/pqNQ4N5+mi/rWQQFC
vn0JyT3Vofy8mGsEf05AvXlRPbCB67y1w9Ksp0yThfWTMcyWV1ik/CA6GBzcJ/NJ
Lt/C7iiyetr42bZy9stEGDe5zQdDYIeL6jx+5InELNnIa2M9wzGkCtEORmeAeTo/
kwbWevWy+rhBg0azbmNPSIAUZ/Ngu/BsLbGBfJHVCyVwNR69zr7S4AKGIzM+3V/p
8AH4zFD4NaGzJ5EsgnwA5CGO+WXjwI6CQh1/CgjuN2weYylnEdSuv5LsCFdeMQeW
otYI5uoCwHb7/MEG5Jkb3pnS1UmTW9FXYQWy3t6PDLq9muqRwQCbAQkkTE2TpZmr
a1eBN/vElP71SztJcvViVxASYCZlYL3PmCEdNtYC1ElWsMH50Ef/F0Q9za4vkw2W
pDORDhxt9Sy57yGIu5o/lxWPCn6gyZ/QYWm6xVQGUcmpY6KmgRwMS9jb2oS2SAqn
PqJS+aVSubqTSm/gFX7FJ14hXLLkq3OS8m6WXpcMx6AuGqv/ZSQgF9FiEgN3ntzo
NV6zEWQUZDIUWK9XcUechrACdMK9F+Bxy9Jz6AUDrPIxKPRcTQjfyE0BYm89Zx0y
vvAyI+3McpMAW3gNJFJ+8BdkGMeevIYsRPtbPHM5Mr+B6V1muvDiJeymzbg7sCP/
khI7JjiFyAMy93tFQQQZeAZSQlPF0U6M1w22x4yC20fGO8S1RH9lUMIxXFRGAg9f
CiEiS/y0b+OKUrlr1t1292f4iJwWHVLhLS69uiIHBRpuO1gBkB2U7SpK+T2Hzcxx
9+fvLLGChxp4IvsubvgMtGIJ7SvHcWcmT6mAsXrsy8G8BG6iLHO4cBwvhpLRgp6j
MCZl81UnJ9mVP2iSbGCoxaIjL/rwGCUAtk3JriMyGU6ZB0RFGSDNSaV9Myswrca6
IpCjSvq6X5bjiOFNRTmH1mRPQ4g/0Q0VjJKeoF0vqAlSUk5G44h4yKqWCCM79BuK
mN5y6Q/mXNV2oWooQvHFnlytKiyatER7HAHJUfeLDxXchnEHj5xHiGxMMPzvkCSP
gcq5Jcu5fWylDWhZd90kU0HT7szbWyIM1GeiQ8tngPBF5/51Bm1ekcUKQHjDAfTE
xpvnZbNtkdYhvyydychrXZM+D5qnmi1CB2+r24xAtlHdA+/6/6IJ2f9Y03NXyZ66
IIQBHdMa7MFejYA4u+YQHfngoceMqf/HcvVqajw3WC3bkX6sul2yMjCyOzeyi2WU
5WRpCCZO8x5Gd3JsN1pkqydC0h5KMv1uxyB0+N9nGdqKoUirM/A/E9WyQ32lfxPi
vvb4zGFrFMNYzntmsnan69tYhaYzSTw7UQgfNDursNOdlS2jAdJbWq1HxiUvphod
QTB0c0YeKtIIup8mPrCvCd3qnG6wIUolnMvCSRFUdU0yx4jv/0ykTYLHpUudPGdW
i4sESLLezdvtu5DCSzRO2jxBeXD32lN7HBdodNlpkvDjdHdU2ZgFO/HQJ/cQzGXo
KAoPYro6cOge+Mj3kPiYXPW8m+F0uupMrjCZVFMdClL5jXw04in/p/CHjn+7zPUN
CopYk47j/0ixDhSqnC58Z6DpduTlY448OvnKeQRmkFJ5IVjxT3HWXZEdu+nlraG5
iisaO5Q/QojXmnSHL7vaqiLXKZ4xx3op8EzzgV8iZIZSuWgzx97bABU+6/qBbvUf
grMtJ9G3JiKqVGnFi+Kp4U5eKakiPIWjqQXW28JATYurHXS2EdjLdcruEVZbW2k2
VvJ2SUbJMKfiIkqPXiVpy1QKvNGOhgei2ZM3M9I1WyxdMxHoA3zFJ0YxUesnHuW9
3dwUKduVODaMVftj8dna7yBKtzpvTfDj7P2NlJAfsjVLRlukj2nHuG0u64X6+x+d
NYj3vSBhSm7NkHBzxzlQX8d5R4bVG6o0t4IX/FOdzFDpNe6M8PVr2KUT6w6GwHyG
oqMRNcsqYU+bSXNrUySTm3HjVbGa+PbGzejeqxzUNpht4O+ZxCeLkVPnuEYtxaj1
9c3f+/zNR78WCKvhmrelBbQvqHQOHvO4p4IkY7CEWTzhOANb8FDAUdUvnk3fCfvl
VVXfGzxQltLdM/OnOGckucS6ark8wbLPwu++kzsfvM4C/AD8JtWHM/gKB1oSGSbh
PrOBw81r9BjJbVDXw7dARCESLSjqZ+YQEH8fcS3BAo/zTZ3cSiOD6xvj21G7f7JO
RrOA3x5UUr32YGAGMsw3mA4lHoj3kiX/+BOVJoQdJlhOdRshoYK8AZ36zqOyCGyC
vPv2L/fT5Va7DcU9eK5AGlCVrx5kO4KUNXjCmRbg5Epme1A/cAts7cHC2hnTnMFO
KgbPzIV3E4/3zVBcqIdU8kOUxlLt6Ul3FhMWpzINszAKHuP45k0p9vBuqwOSTSsH
1YEQbIqTtMN6oGjMfMTVyevGCyE673xB0kL6A6la4gga1UC1tcCqulxxuDrPwpgr
uI6ow00X8R517XwNjZrh2g70PZfT1bNeWG4Lb1CkNxhC/eTZSwq3+tbPjXIMIbhr
Tm/JIAZlvGQ9uZAD7/x+Jm8BT9DRAN7FcjP/u23ZhtJ9y0cLAAs9i0rtfc9fuURM
gPuzWRaMAdb1+ViQibLBTIFJ5wmazB2YykKoHTgwSz28mKMXQKZ30gCal7ypedLb
rDujhQeJ4iHwm8N9St3nIw==
`protect END_PROTECTED
