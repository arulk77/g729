`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zW7TSUNThoyoDrAd7YV6lW3mXmuSye1Eh1L2YfiRPHu
6UZxMtcXRc55iH1PiphNrV/n8L9M84FumkG4jvXOZGCa7L9BAAip9CjhOfmFc7Vo
dngRz/JBpxivDWZUaCJiwj6np40/9hhWUPTvUmUXw5K/yT37OL8y/hBNCc0rtOUV
8aBQQ1eMfT4IwGlX1SaCQJC65HpneB+9CIEJTdTzI2PpFh8CVhmZjw8MWk3iB6tC
HAYkFPv3HRwc+rBTEf6Hd7IQEv2wPdrrCmN0t2sXk/LG/soGjEUmhGynjy3jqnqX
eOYBjQImYEH7YUmHda9ZNg==
`protect END_PROTECTED
