`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGDHliBeirrmfBnHjTxzCJssL/MQGPFqLk9r0HKTjH1j
IKuEFhBO1ET4AycHOwTnrgYrNQCEK9/ZhiFjHUONRiIQ945eUfLuDt3h/Sm9VdzO
SribZ20XHhn7uGvKtfeaIT4o6rPPGQZ1/OtvipNVjTSWmehK714ibgjEwmq5YsEM
F2knE8IULBDfWyniemnW4Jy4QjxKiZg1M9UF1mKpGcoBhjOWj60mr8UIGnIT65H/
88VGfsPbhF2RMI6fMXckNnytyVQ5amgv28zOpbgzw7bBJC2nv2/256Nr8npQF6Va
wyBsLYqDspYOF3Fi1SuhZgd+LglTX5vnHZLr6afP3UuQIE2NoxlnIgSA0Jy/eVce
`protect END_PROTECTED
