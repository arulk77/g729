`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
jWt4zdhWj/rkxXtYBwtdkPVukRgTaIWEOQ4eUpvMvR36YLTKTdMDTkQ8MOHyUSzr
G+jxhRnpnt4CTqVXb37Im9APaAmtkFFwH3+8p611qeQsX5VWo33T8rPJwezFkNWF
2weQ/jjnSZChd+91XjvSSeuvHy0isb91ODtxz1Lf9yU7Lwz2gpCOq16rU2Biyc/T
`protect END_PROTECTED
