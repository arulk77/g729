`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yyj8OugE8QSwxd21LagEhd+BolUn6JGWoHLJ2aBNghc
ryjJgm8EpOjAiC0wKHDaQQNGoqyyD5109UXVSQU6pfR/zeGegvKDuarCHhH2JeuN
57XJDzPcz4AZ39GZzv621nQHYfFEswht7HN2UyoeHQ9/mUqcG/GDnnjVhGZbDhKR
beIDFrXL8NrbGcwy5zdFli0F6d2ls6i7zWPgkw2OjOKcGgyn1Q+KU+fpKiwGvfsY
6lrKdgkqV9CNtDvaJpBqAEePIYJCyVD8fDkOlj1wZ7LvpApuiswbxCMMQZuL/ku6
EPx+JfPfiPRC9pjYTUaMOoBUtTulWrXk6VbwfzB8qkA+Ft3ZZ+mFf99LCeesPMdm
B/u7ypOaKbuyAS19ty1FLuC56Ftyg3O/SwretqbGecQ9+kcx3/A8bwMi/t90SG0n
KO4cEpI0YF+1Pv7r+MQSdJ4DFePdFhqbXNTdoi0eeRc/cwaE9UVVpISB++MT35zU
`protect END_PROTECTED
