`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xRRmt6AQx4Xpp2VAgfv4aVoqxiD/62JuKJGZXlPvY1r
Mj7OiLSAnAbbRDuw0fvcFAm80adeRAV19x2X16ESga8JdpLCyKVmxnkkYAfM4Em5
mI7I8bM/T4nLT2FGLUlTQsmDa0eIGMtzhxJQ5Xm5hvxBDTI2RGFhbZa2fkiq2bZ7
Hsk3Lps4J7bwGEt8m4EXjHBxGawDJPVJAoJsphWO/SIbX5nbUgWLLxn9RwNDUjpK
63faiejuNlJKYBtb4ouFlproshXhqRAebLbRLN4T7ECzG65Q7I2AxUXSRUymwFbq
3zLy7/qpQrEvj/IG8ME/erjnoh9ESxzTfrrrr/MQAb22A+SQGL9BuOX1BFrQd+oX
ryedVEOn5dmAJw6sdavp0Q==
`protect END_PROTECTED
