`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
e2XlA5ytclJpIcud5/GbjECFHFOjyzcnNL1DsPGffMErwQcUrrE3ORrSZU6FhdAD
9I20ldb+8cyQtkbAymIW5gt3/REM0qO3oM/NNxv1bW2YqxloCByItyKUmx1aLcPu
hH0li5MrqJI+ORNANO61Hlfsb9kMDOfLfsBSAH1hQFxEJAcwUnmJqmblgxY/tBBF
BrrMX5iwLytK9Xiqug4TuAK1hnS4gGo9PzpWrxeG1wFP/kkrd8sM2+Kf7jzZjFUs
qL/xh2fCe9dxMiRCx1HBwRdQAcG391LHcudcVbWzbBNs9LqGoBsXW+HB7ZMRvrau
`protect END_PROTECTED
