`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44/dHlSDV4cT/SeflUoGDrimQ8r4H/ItdZ6jjrfQUlbD
a+hcRhVdpe1g0Thn1RflAW4nJxIhXMxYa6EAB/3ZcX2aC6W827uU9mwR2wIMXHPN
hColN0ytwKFdLBY2emn7S9oXui0YIdI295squOJx7dzIK340ImwseamYo5Uct/vk
+JRSScZM80+Hr+XJ7NiYFiWVwYMo/u4pu0DiCoKOHOgSuMGY6YBbWIo1Y5hyv/XC
5FPIo9ZnXNoQGwUdsYBIQXyUnYTUlE3G75CB882VCnucpNZLmi18PWfKg7/MlFfn
oWRNxzvOviy5NqUnJbGfjSOCZ31gx9BcmFRh3FFWfS/TLeddDav9cW1UN3zmc6YK
nEAbMfsth/mX2d8HQe6f1w==
`protect END_PROTECTED
