`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIfBjiqNzLbpQfvwDq3oBMN0Wnu4vBrhKAUCq/GNkF89
n/TUmur6FLZEKsnBl5aHGAaCN9WdrkUcdLb2bRlzp99dOTuap2jwHIj2OI/eVb0z
73Tm8YPt58TrzUKhsyc1sPYcGclZ10H7p9nOmFf+X3UPczNmDb6dtylvBm6ASq6L
fcf17XATDGZvOiejP0stclVLXreXBzrBIcQUSw3qBA+ok66ZudITt4M5xqhjv4ni
N73cZQ0GKDKblDbSNQLG04XBe5JR8ugHsHY9FXLR4bY3GYKe5fJt9LvEFL43fDZT
NsneMAWv0TAvqrC+rJlDmWWvSnuKspLoeVwIHAorWtb6r3vuIRfnO5V+1iF+41kt
GdtSHpvE9u20L8Ck985BFkAYUTrJ1p1CYx7T7umfSdiebvty1xf6jgWlSTXT8lh6
Ax5nm+LmN7W+cUPq6uCBHYB4WSoCrFfQrV4//cB7eU0Nonetj1rZG7soweAmmIQk
Gebkl4rrra96nlwLtFUzQj0unesbX6EzQZcXGWXFvcroPxYiWknSBiR1iBQb/9kh
`protect END_PROTECTED
