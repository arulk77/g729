`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
5gJ4bk6PZR9HZvmOF4+vh0ZaQtaEzSFYJ6b0220Piy5kqo7st7RoN+VGCX0Ljv8R
uIrzvDl/eJqiixcabQFAK6iyK2bcmHKfuTFJNVAlxc34ZznkWi6JkDdFVxB79OTe
A08t53n3+tKxeendXFHQqOX0Z0DvgwWKU+jwqjhobs5GNH+cPgKy+tMgK2bHGeh+
`protect END_PROTECTED
