`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL6QQY9ihBURZeFDACKjSezcbInFPzVA71jG0FhfFO2P
LYoDakFqgg/ojTNhfgUYQw8omD4A0LPROAuZbFuSB2AvDDlvKlk643GvWoNn35iu
6X3rDvuE/lf9Lqe4cXhpYLNVGITM99Be0kf19vf4skOu2w4e5qE/QAALhUZPSGff
zodOS3pg1+1HhxQ59Yl1DPRCCZvANEmFrpCQ0oq4O9mcAYBERnhpbYqiRkCyfHd2
OpbJENhpuFoWO16x6MeozfqbR2yo3NoUbG9cjlyDSyLbKmOQpgxmnfmaC16PmkzI
kCxyqZkMWKysY6fd/ybWHDaGnE7oSlpktXLEy66LaPcmXsUsLCKshHoDyHJpLnDM
R6dyx1B1JJH/zp0V4esOag==
`protect END_PROTECTED
