`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
y3fNMism2KAz/57xN06w4sBY8dXMm61bUIMF6dDizY7S0S0n7GafymYz5ryu2+hN
rYiTevexNf1CEjwr7ABmKppzbD8ait6q9byR9PViCkfjj6GNJXT0tnjZMdLKRSSe
GqXoJc7hXhq8JS2Z5Oe7lVGBiASBgMJNM42nH9wOIi8vVe9hmWSNqbIQzxjY9Xgg
`protect END_PROTECTED
