`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zihopCZu3HIIR4/hG0O09Nu4hqePgJX96q4owEVjsx5
loC2K9XuAD+lPjaZ1OY9Sf2oQYL4hXfyRaO2gFXJmoUx3Zm5i01O04xEjnGRerhm
I2hdxhHcDvqO4/CoFScwFnUhJ0iQVUwoLXCIjnEHMrYCJEqtCaQcoQ6yHxRQJNCx
4PagIv6raFfOpPJ3JSYr0v/jtGqNiYbmCvK897I/bJ+XPknJv3jo7f13TaHjWGX6
ucMZoAVXLNFHSn2YjxfApQ+y5xqIRfpdMY780rOaef0x4/j2OurMkjyqGnRWDG5m
NU8551ZkI6rS0RuZ1r087A==
`protect END_PROTECTED
