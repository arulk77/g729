`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
1QDqNzACiL9Cg/+dRWiPn9aIxQKxEYmhm9K8Pxjg7mcpiu/JUWs9+X/LtWpV/mkr
fbS3nITN4Z0fg2NaKJCUCW21ZM91zpz47kG3MNJM4WlWekA1J8EbZ8GpYFCbgH/k
cbupmWg5v8FGg++f3jxiQCCc8UEw7tGyP+/bWzpjgB9xRvUVD77Vz62BxiIJGT6M
sVSVs8bYmJPUg5zSL4OK83yiUdxX4wHoaP8xXvDQ8LyaH3FsHXBiQK7BZD5aGNHw
sdJWyslTRbwVQevhOwipPydY5ERvC9TaXXxSJoA7BHvTf5lYvrWkINakxI4zr5rk
xoHXg12gutvVA06VMkYIWlYt7yDw53tdei3kTD02aM29k7qot8SSuxjnpUAWs6Xi
JcglyoQw1aFck1j688ecKCqgJphBnieaGo6xpw/cKKhfBiMf5/YzFRbEHY8kYfIA
`protect END_PROTECTED
