`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42NxU9WYMzLDYctWg8DUFOzY06SI8Bu7RAgfJ+Umhkj1
xP8pChM78zDA5VTxxtV2u93oCi0/G7ZEAyD9SvDjiLSYA635w6sotC4l81e1ztV0
ancQlWxORNwLt4BiEnCFnp2W5wZvBia8M3LsgIE1gpc=
`protect END_PROTECTED
