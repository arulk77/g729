`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveH+0c3+cPUhhJGZt3NKdQlRERR1/17+xGnNfIxFt7GHN
PnDQbkeWLkPHl7/6z+xSNDqPEh0xFq/6mdnckIkm7tTtjusUhVsk9e40p2p1yQrk
/cGk11wKjNYjefTpTyBdfN2YpKqU04lK8S+uKsw+m1Znm7+8Z65jKOQoCFM8TrII
1qnojaNws0uu59fgZL5gpaOD9SKEl9BGY8XMMiypJ1fo1LcSaAGZm2n6smAATm90
`protect END_PROTECTED
