`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2OmpkLaDYZ6ZLbe8rKj4d23E+TANpYaYbCnwZhrnQjjzAd38ijAVF+BDQ5PU2/MS
Ie3wC/rlMY+6GZGV2/hMowiAht5OFgw5lPFzxGWku/P9Ba75mYUYqQCoxKtUWV87
YruZmS/SvSobyCNUjh44y9Y6BOqD2o8bAeC6zhFk1ynwlyapWhzS0C7G+m2ndPzp
HBJnXt4kq8xSbAeTwfcsdAbYzVuRqg6tzNTQsn9z9E9dykzB1qTMZ4yKRQY/3gGo
jcQqUPD70xTRjFPy2LUnzPizZaDbjtkN3YirHs8W2Rg=
`protect END_PROTECTED
