`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDATz/elSRivQmgj3PLrSzv5NhV/DTwWOwP49/MLEfFS+L
ULHWSJm+PfvjLJzTm4OYW1b81iuPpLTrxcAOU3gu29PVgqTLA4QV8W1w8BGCDniJ
e30JxiWo8wm/Nkpkyti8mOrgcp1eBDSAenTz/2j2SxkwuJw8SnUq+jMrCM712yQp
r7LYLJ30w59DKrTHMPeEa8H6kRZQ4p8uu+WuhAPvGzZ6Wa2cHXaC2+b0z/Ig2Qxw
Epu542wIJ44YxwnzxGtQLg9dyz3uR9lnQcovEzhwrh7A6WNv3vITeDzP/gyuH0Aw
x9iWbqTEaW7MP2h5tZ8DMWedjXvpJigxU5gyWys3k3W19VihuEs/UwWFU3lj+F3K
Y5SXceHA7/cVkBRyhAsazyh9xvEsZx3t7W4/OkOEJNzqKJzAV0foP/22WDtO8pgc
jNGqz7rE33rcdl3V6mUOhx0dneaVWenIO0ifMfycMGD/VznrjxZJEw3pyvO76tco
BslQF/Si1mMfHZAQxpBCjm6uSfQZKMAZ+4Ex5VPMNNqyNhaxe8iwQ5wJO/61HtrK
vwCZt14TkCvaONkZ/YvRKaSTpUiGBKW0Ja/0Rn8LCwb797tx61pFsahgO1bslJm1
vXFEZwpqFxNi8DIoD+/iF6uV4A8rc9JgiMYrdlao/JRqMkfhNIMHnxqynpA53uzq
ix7qzdBOzmjVS1gputnXhqpMEKfNvrqPSjrcogOb0HRSpOV8FOThsQU7hPJEO/8T
aE/A+qGD8lAPJlh7lk87M/d4vuZ3FEMEOySv4b/nCNEUOTDbihaXtz5Payl72N75
e7YrKha0Z5z3MxUmvsNj8z/nX4cOn8qVn/2VnLVNTuGfc9sxJ8f2cieezmsRyEg1
pkeUd+ZlydmX5MpBZO9PezwAFAO4Qrg8z3NDndt9K1xYSCgxto8KoAaq3b6HIo/E
8yhcoIhDGjKPJxQxLRwgCT6GLp3C7/RVHb/AXr63h7r9tArB7gihyYobisIPufmP
ZvEDKoX3nu0eX28cvwXrmTkVsr4o4l66/83t1gowL7KmpynYeQVEWTpy4HK/pFQd
oPfIUsk+wgQ5OYlxF6IrIy/0ZTf4WefGrQZN07GoeDazL/p/2kzZRJMxXlQ718Jp
hJAHonS33sS43p/7TgI82VC4NpDVN2zm0dHeQWKgUr5BemRqVl6aTCStsvgUXj4v
v7vJGbZjPQ6M7ya5oEFUi+m1ZA0oPloU0DiK/+iSQOowxkrNd2F1QZEa/kVtk8VE
ZMOmkcwAUBjYdzy+k9cDGaWoenYM/thhq5PXCmEkWpBJUo8GIjdBNfkXfz84dwj2
z/LbnvZWNOc4OPpVEAyYkWJA+72NOmswi94JQB0x3iiAE+Yxi4zdGYKhahBQyMeE
AdzYzL8NjbUBSocNTk99xNPsp0qCzGOnZqwN+bkOeUGZipszxCeYW6r08ljSSbQ6
UTjIbFpDS6zOfWducRZ6e8/tnTh32LU9JCp+dBeyQhTJDTSCgVxwsLSGoW3nkQv6
NpOYGmzuqOeGu1KcqjvLtUtYH0rP5HD72yivXZeLaiko1CH7prgrBZc8LaGPahBL
oJRmeDPLqSyBevaRNXqSl/Wxmb3kRSgMVaAdidC5gA3cPx6Au3jkxcJG5OcyZAM1
+PwO9McW1i016poStRD2w+HqZ29d4dA7CdS7I9SX8Gd1PfdqErX0UQrpbMFknnMh
h7npBldRO3oLHuAKo6TWwq8tj8h4qsKxO9OYlJRFFaHyNuHnp3CHzQmsrAd8K6d/
fBsvDG8IwHFIltIqTRrKYP9ACOiNo8T/1qDxe+TUnt1iAqBJ37OEwtP4fNeGoXIq
3j1ZmRLjYT0ZVWbMeukf2q71eb69UvkWZQ3+BGr8TtONsF/gbQhjPYC9naeXeXva
PTVHSeYbEBx03v+xQsL2WSyDC2PlNyPwkgFi6IT//I9JGKre3j8+CYz4cc4U7m1v
skwyk0hvmRlInlG2kO8A+lB9HT3ATOqlAZPCSeoJ5Kmlwfi99u09/d4Cg6kAv7B8
2c+rXWO/+ZbjwaRReqU/zUm8DNHE8E5HWOTJOMK7cqGEsUSU78wvUswC4ABKnGue
aSsUAD2NdrzpbpPbHAr+CcXXuFfIZQHKOBtI+VZ4J8D/FnXaqkAp+N2XTSohx6tq
8/NjQMU4Qc7yQ1/sLDEIqxvSwHAcaiaiZHgmUO74MtaxFAQFJxpNB2Yr751KCiy7
89o48adRw/PPE3HeVQH8r4LS/lskQLRboZrS/KKMT9/JR6MCdU18tbitJKxCt2jQ
Ngs84CSkDKChMXOmPlKrr17YIeWgaPChPQF7i2iHWlXO4TeYLPOHKtsOtrWXzBPP
8U8Pfs1Rtyinbz7RaiqAN4tSeUjmyUKQ+lXKltVhVk7YMI6AOzZ6H12ERDomhBBI
Lv0mm3B0QTyjP7rTHtyztfJVR67Cmd5dmFSogYhOZ2XrIwzEmNLVQtCftx5YdH1q
S1BckIzMLiy5ftByHYTs7xIJbT3FEWUV5TIAlZCVVb213rzOT0BDZ8cSdV7cJapX
bMFdrQiAfitDOafupTFhz1gbygi8Q0IfHzE4DX0r0BK0pDXDfr8VjcKeTyHC9rIt
/7QpqZkfVlzZ26mR2kmyGNHZb90zoUdH+hkXVWH4Ur1AXt9ogG/QUhQ5//nmjiND
m1Kqg06/9QL5c5pqlX5aYcW/UjK2mN3QIEIqw6zvgU7c9TCtRLGOhh/XsjHHYGVL
XS4J6vuPFPAfjTnRLDbw1PS8PXoOnOPvZ+z1whLmWXBGgvlW4kYuN5dBdFpwcKP7
SyfL9b/KqrEt1IfbQbioO3J+3MIfhU8/3rYExWBINMZGZDoQPJaxOAg/lqdacyzN
MEhM+bRJIQYdGGglVPh+TD51onISAquBY9JHMz3sb3V+8kfGfGC1T1aayqMWRnCH
rGSF35oi+7Jnh2zcHBAUqr4pAJeEkoOaORwiQo9h481Fq+l3F6BYgykrs0Rfa1zE
+Ruzrcx55k0jd2LrwIfQTYQffJ0zctETXKJtM/R0/J8B4u00T5lGuNz3bK5woT21
6slUYJ8yd2EJBy6Pi2jhn7uIVUrBVDdOJJfZlJL8dANuiEkQb3tLBlA+E4xKIf51
rCVSIOuIo02xIDq+oYDfqyi3EhVFpfQPM5p09TEEEojXEuMzD1sQDCKioiC1P1tb
obOPoRF+gOtHIwRzJh/clhgCVm2H1ywa93QFgvO98eziY8bH4V2NmF2UcQe5QikX
kqcIMy+KsrhooG8bc/lRbxlfYYJpivqWsJTtSIfTAhQNuQTy7q53p+RXKEk8YP0f
u+Dd71AfjKX5AGLAlsx5az8vvxAH4Hc9XZo46t7uq9KmayICsCTu8T8y+ruQUqan
J9VkeCIqp4HyLEX9M5ftZ3vd016yZhtUySDPM9j2eWgWqkl4pTVbRyVMBCIgcVXg
ETBGgwme96cV/qpRf5g8TTNN2a127kcLpEzNGo0JVp8NNXIKnE8eTDHijtH3mKwP
WnH6FiykQqWWE/Yd75PNdYnwEIfduKUmr3NB3nP/j/BekUbG9LtrZ/pOfiVnzW09
65VJcFTCC0ZNc0jFVZW6/0z2nhHjEq+qnbwsbl2rE6bAdOq+2IrbdMgJesqMD7Ha
nbswmHdmSkKV52Mv3DDHIqkTPdOJAFFwjrjvq+Cz5QAalMuU3kQJTWFkLQb9qv2A
3v5tXNCO3M2YibSCfjfDmfCiF60YTVSegmZu+hE0w/bsBrvbfmvBCsS7i2a4V5Sh
gSn3haIBPaatgKrjDUnoTBWhHYhk12ggsICliKTXepGiFHVld+tNzQoZvp535DkY
VrN4aSmfXHr4eJ2c292DRwGWnusoJra6r3BG/+rL8czsswaDISDiKzG9BszwPvk8
xpoh3OfbgpgFnm+9UFmQSH7Sz6NdEF5Khp8cM9zBOUx+ZakGUxgFyuCpgMSR9M7F
4boXyjf7Bw4GcQn7Jnd49zPlJuJyQznsJYcxCfDDY/KzfScNQeUv4X4gjYM066v+
kVIQkb722kcgiFBFwd5TzgaiwqQ0RUeCLOlBHH2SbGSAvLeECZ2VQGuAVLNoHpdD
QoEMjdWnpPVNO6DWWNnKY+rOoh/4cKNdEWmLxYqrZ4hgEb0vHQ+nD1nml6tsGr6b
UzvQyC0UHRRg3ACHodHXD5hh+EeV/OO5zUdC1AOPXA8vkc+jtPB6VJtyYrdnLjeP
PdP2MOrj7gWrV0+8s6i3RM/RZFCYxyqd5PdULwU3ZZKdfrcIz31+Hz8b+d69kqqd
0l3KXP6nVVLzwRejwCkSIbmW6szt4GsggJwVWI7tqblNpqdUN//OaaeQh9mppq/x
RDDfrSLRsLD5LAQPnYYXc2rHAQAr/GR0ZiuIOGaMwlcEp9EnDKbxymVUYaVNd3zS
cRf2DdZpIsC+5REIvdp0Sys9DjTVyVkeYjvQE2QM7+5nUfS8D0SObsKBjjDk96wx
W8Qhwg1D8GEyZdfyRxZYnW8rJIJ5Ye0PhuZf4DDTdsAZcQg18M7Rltd3zH11IzCK
IqYcmRSDfRuFX/d8a05GB3GeM4ctDtAuceTBITDdvLlpHzvInlUJFfZ4P1HFseo+
HBaOPuvK96Rduv0M4b1ircKfXScD8jM1vc3qAwVuBU9kPttYV9N6pwPmiqHV4Z9Y
f/n0K1woMTxz2Q6+cdYW5rnQQZAbxcimQOhGvGP+KolZ4+l0b9Z9EVWgZEGihs/H
jB/GLLjrgKbhp/ghpc071QLvQCzg865Mu9BdLTtnWThklVx43m7yKaN8rNvzWfR4
bS4eNIBIqRkJTinAv6GZMmSGSuxJcV+fqaXE4pGvEiKs2lgPlpxkbl0E2CRiWY3u
7oK8Ma+WCQMvR6s8PSvrNQf2gty0TwVpvxZiwof8UvFpDFxVxPEquac/Y6pqoLKF
tyUAVFKYwyxdE6yy5SQmExJol9/GiKMJBIjr8T+zvQQ61sQNBeoKDowDKOjPnYS8
YZiORttPjeMK/N9PXRIow2AW3MGdNPWhIESCtcrB7ecWcAzm00zaoOt04XLrzj2A
2PXS6vNHDDTdo6+dqcpnvdaSgpvtw/keuCPT6NWq5VmfhgfGL7Tu1OCC4WG44Y4o
tWWQ4jQAWvXss3msMFA8T6OIP8NfSur5ZcnsF1JO+bclawRg/D8SQFSZQB3FIeEL
ptthNMNAZOnuJ6oG9OQMp/xfJisBL78ckhQCo17/xQ3J4vR0EzLN5Okl71iGL36Z
QtSMJSDLW2j6fytr7aQATslUcLIVuwZ8fQ6NMRBl4k25ehmLXe0VR/STWGfRUF1n
3hrefnd7Dw55XSE619RG6ewOtscn3T9fWZtxxYLcM3fAUBoRyio8UP+leYVOcnoO
qur8FY43FssdCYM24QHNQ0VpZqwSdYvEbYIrDALCi3Jwi/qqZjOmBGzIEHGiZZjK
fxEwd2VUD2Q8gZsSWEl1trWB45Aq7BExvayn1R89dFpYgxkqZ82j2lI0Scbx1OY9
tjK5IVZOBw5LZqN7TqnZmXEOmP43KkRzwP2TX/l6/sGH3EIYG3MhLa9KVvvx0H20
vXAJuDHlok7w5HPLox+7pDup0ZglCn8/P9WDKIpQ4HNAdmCywz9yz7TYcIM50dZK
wiODSiG8Ur9ExaUkQi8ZLkmDsWtaK00K6kBv4pwhKYWeVLqD3YuSt073HwyJLStf
DTe273NG9WnAo383nAkdpVEJKp2TsWiM+6aOdvDnuW8yDC3vfHqeJ9xvPaHQgId6
LOfodLr7Uc0tJ/h88poDicAkG1+QoJdzGgAeo4Y/2uJkbfsVbPflrid5lEVvOayM
XEhl0KpE0lk5PzoPAC/H04+cB3MzAxGHrtmkPTwKmLBtm/HnsXZXh5jXobaJCsg5
Nd3mMG99qrjSSpyI9X0/vpPATpqI6PIK7E4Jpv9octfnZ4v8CaCW0s47rbpWDoLd
1uoqUtoFjE0KYVGhd+L7De3yDbT38Rgjyy722h0PZVPXuaInV2KR1K/4dyK/4WJs
b39O7/YBbt5qraSjPPEjVzvEJO4jNQtr3zB7K5NKuyoZJoDBWYR3Jpm/cwymFACF
EbveabE9TXLD5na0BQYU4CUChRi1YjZjWwBbkEVzZpt9atxNRC57MY3fiQ6mYaRS
AwnonQmKtcFPUFRQG6T2jCcfE/2MsMUePP1P3IGnwRBt9EcsHvNQMKJPrnbY17+G
xBqf3PGWNgh+tkUqJa2DO8gWQKoZAbN4g35LqF5dp5hL1SbdJ7EQXaRMCn0LIE6u
CKpXK5jqv+RncMD6/PtCaXB8S3YBuyfZ5I2ZbPoUb1kK+WHtcmMuhJO8oCF8r5ig
yhvpL0fAkI4Q6e7mbbeQL8RJY5BkhDHGoBXbxlIkjh2VlXikWOK/xfO04eJgzqlo
Z82qnAkQ5Zrk3Cc/ZrEYkPV8eDTg3pk9+M6z89rargccnWcpZYjbm0UsUTaQHhQg
AO1qTdu5bZw6YQNRAMqT04kWB4Ax9x6dFbLNpIU5u+xOlXvnaBfsuQfqpPCb7j5U
IdQ+35qAwm2C0n5g7TukAlJxrJkxbQvY0RlyebNJQWO72meL944a8Qcw99g6VLr6
bkxmCAbRGNvvMlbCAABuXR5K6K0UpX94gSk7G8POdCdsLbU1F3SMH5PaTMXN7SSf
Sw0nACp6hhxxX79fFWx6rTJwkgoi7Rrqv9Qr4mZWkV2KLV7R50I6dlHvMScRGrtQ
KSZ290h/K5VO0VdDbkBLty8UZqy84PfruOeb8tta/KB/6dwLXxGA9E+iELPmO1Bq
7qiP9lIoToNjaXtJnIK8qTIbuwqlP1Q6D9M1WXypwR6yunUsf1F0/kDqjm1jTQsL
IYPhQ9we9M0QB4v2mcM80hkNpGkAgVLtCTzkP2wMKqOvzMR4TLIcxCecESA9Akwq
GpCSgSKQ6SBkFY/GV/j+iCl7CASB2QGagidcGWxuLbFBqnwh91ez+K/EZEaHdJiQ
gREBO7EFZm/DFlVyu8FfOk1UeigLtd/La9PXSvGeRpig1gvHicILkhCfHvKb6Iv8
rd47KRyOXQvC3AEdVcyYLt3B4W8bCO5CBNuirrNp+dStrBRcz31nCPVnmW+hB4nu
W+pn+a6TFABwzOELRlarQw+xGWxz4vuWg0aAWRpLoVBnWEH5g8UBq15bfJAe9NIX
oUSyff3nNVnvxrSjytxLu8aTCF+DLeu+dc0sm3LLfmNTaBXDK8yReVAWFLvNXsLY
d3k4bMz1kUtphIvi/yQu16U/h9PZbOW8wDLMLsbrwuKEfskXA7x0RZL79gT3L4Ja
S6J2F0AQZhW2HvdY6w/ZQjtYsy6lbEW9/qLrfiGbQZGhr+5NKpKWdMlVSZgMWPT/
7gsy2lNHsAqJdMJomc1QhXWUTg+5AbpHU9vRnykZO5Ahw8KuAsS7vxitinh++ALp
0NGbyj1iizlR6S9lcFdvYZxHTSKMCNnaZuFHitMGfrjIIw2BxTtu3um4O0KuvuEj
+NHszCSAWulGd9W7yjVdjqdlAXRUvfvImUYzJylCE7M3r3sN4iU+UNlrpkUNs59d
ZK1bkIJYPx9LbNuevrbok7OxPWWfu+TwssQ9noguXk8nVDgSicLG9v1VB+FLvpKm
dMHdxvu12FMQJt5Up+SrmhyQBXeLVDmyxes2daB0IpFGYLgkqSuLsrHMyPl7yXdh
QICU9npXYnFJvKjiB4+BpRsW1HyQj1A9MXMKSmnvkpx2DqYq6/wKrMLDESNyKuSJ
NHt2CCVU0jDg43MG4EY5xeTuDp+qEvcCCt3DN6s58RkXXAkTSI3dRN4GX+cJZpDt
X+l0SqbZxxDF22E28aFM/poUlZeIfoqDvFAtZnsB3bp3o6/zmpgXvN/XJnY07QWz
RAkpH6qPg/eBUhjU5MXI8Rhy6++foxpNEWeno4KOYNCMjn0VhnF2HFKD/nTxnnB+
ROQyNx4u85nTQ//ioJGJJ/4D8QHlD3E0ER9+SPv4lzCNqiHisVtHsIhGBgizUZ9c
6C0uS27AyJvNC+oYcmKQAAxYlAH1T+izGcS2obdTA3T/I3XvCmwfXjheGMgsuOne
EiA4aPKQWDfWYV9VudjH2D51j1wPxvzXJTKUzzZfqeRtpkpjqm5IB62XwvFJtvWh
GazIl5C9ig+0+Ty0aOonMw==
`protect END_PROTECTED
