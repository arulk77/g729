`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBIHW8Kp4hRt+9D95MqIncAAK7X5KGW11AVswgzOpFPC
Gq8kIXjc7dWDDQ9/EIUWRZ2xkE8mtSNkyNOKFM1Swi+T1jXrzX7kh+B78kNZy97P
MWgA4G5AeJjcIn/0y8zskaNZ82tvSUB5WzaP8T+BvrU0VGh8oX4n/6YH9QPTmUaD
JoYWhiP3eHpkrJDnhWyPsCdCv4FysBYs+3+JwpKxnRltyi+1hUHMfFhT0XiL6gMM
M3yF3IKaPBsHzUUlziNkSoLo0pUqi8P60rk2prv56MryGA6ghG06XBoQLBD43VDQ
pAtT/WkNPwkhsMo0LrCfkp2CR937osvuWI9DBTGxRVEMSX1TSO7kJH1KcPUyb5NC
`protect END_PROTECTED
