`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCAkWKILh7xKOskIDB6+c5RI/XgZI0eZSJBNIi4gMNBU
QJxxu+Mfr/gaTNJ71yRkRXB4g54tFAQj40108lqW6ZKeldbeY+ya5q1jPst6Dq0G
iPaBHfo+nwOcoLDqNu4wRTuvsdwPanG76g+kGKmBYzfr4eEOcOkLyRTP21JigY0g
wqFdmAGRSPBQCICLs4GkV5sQyokO1Yi1zluEskqlmDuBLNXxgnU2n2B6/raPAbon
eCNkn6uAHnYdaQZtiDd74ApKsDWl5qJadNJa9l+iMFpIQGUsMeF/EzJwxAUbBXlf
wCKEzQ9uUqlmH+NyslBfCg50FjLjQiGP8a2WCkrJGc6DbsNtEv3lzXJLijdn9iAj
yvA+6WHlB4DQe1RI34jzfCgAihOfv+tnMnPHo5XCuwA4eHLPGvpp/XiQvznlYoOa
cAwgxyQHR0vVw4xJZ5bKPcM4uG4XR9D0qUF2GVXjkbR3f/6vsjscL8QMz+KodBoi
c2OSvznqW0EwO4QaXrMcbts0dqLuCVxdTNTOL1Hg0J7VQMkTfTtoDXakYWXNcpfJ
6e8AUofEd+4PiR/A61K3ek8nAftF496NDWKt9sEAGq18lTesbojkKv9eeknPbxZd
gS/2FAQsZpxTB01G6+R9yKKFnh7X03Eoem+BDx/Tk6erk/fOhvJebIY3vQBzlQmE
A3US7dqNGJckQ2vUkeUwe+iSRyqV/H2Lm0UknYbheczeDqbBoXdhddlU3meXFiHW
DlsnC7dOfLhM6Lqsji6L+pINgulBpG8BrXx/23FtpydgTlh6nyZTgjhlPxRQoHVu
QYth7KFcwI0bAJjZFzapkbdcIc22fRHV4w3WWw57NwmLZsHetaUHdVam11GVkhGS
7YhadT26UYAd5Y8qZittPNlVHpb89h6i1w0GbrlOqux/PeNQEVtnRCajhDOM3Qms
tcx4uF/GHiKpFjoEprmqEJcgOCwQ/hUGWZQDQnYWRZcyozNK0LV74bb7N6p8AIKX
dApJmn7Lug+f0w2bCAMF6nWFKQYYcC5dTEjzhR8KQzc=
`protect END_PROTECTED
