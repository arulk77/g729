`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBVDCWvGOE/rt1TUiFFQxugnxYP2hC3GNdiq6CJXHKJv
Ta/1PDUTU0NT76Q6kB2RV8FMTiQhIEmbGTfhmnFBqFBsXazsD8hf8rqf6IYpnrUb
lWsgohyEtFVB6RkIhMA6PW3Ttxmk5vYs1CDN9/XPTRXqnvlIOmrRIDsq9WKsTC6H
AwygwJfY9JNTtnK5Qnp75/tlPdaPZ5HUoIk6b0WfXbPYcF3ibRR81NmEemWZulad
`protect END_PROTECTED
