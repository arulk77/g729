`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCxDYJce8e6eolDZB01zsDduKt9C9DTi4p4DS4pIKgru
zIca76iUdiDxIGjLwO4NpM4EaiaaU1PkebRI9QYUZtBsYRYACkMjx36Fg+/zAmoF
cNsYkrhwoOtOuT4dhQ27iyL859G4FajbzBgFfz+R5lLkfK+xS56/DUJFGGOCcsOf
UFHH0Gg1pwW1f521um+Y1RWS7FAHjP2vNq58VISSu7Z66HRDoriLu3ZugqqW8DUW
hDhUpfgcGJWMsUjKiml4rRTZ5txTec+bd72WtvVWvUxp65++f6rC+eH8oKJ3Uv9s
OPVYGqYtt24g0RIWCeSLiAcPbEAdw8k+/1ko3ntWOsxhTcGKNpp1wcwtrlObW7bN
rCVB5lif5bl36Exu4ZrL0pyFswms5ez97azvVre+VAdXhQpJuCMdl9HAXuoYfVvY
Y7lrTP/irKnH+6/nwEbTvLjj0E3Ee9Cu6G0WJ+j8JuJdu24ZxzKgwB+sHZVRTjAt
AT6mna3JkRGMIhX7a44y0K5lZ9NtBa4hEsRg7HvhWpx5CX+GhJPg9HiVv1Fe70YJ
j1GhmGnKXbHSzpfgqDE31G3QlClrez4coER7qAZg/d+EszGyHqelxu617xm/tD5H
PVwqZ2fx/raZ7FaoZQQwLzwE/9yYfjp4ODTLQVmUL0pMY/IuTl9NVHu19y8XyFQB
MPmyd7KXQOl2RoDQw2nawNm+DBxlSHKjc7QF5AZOnBdOC8WKPJxzOAZ3MuVQgizz
p/9pfwXVLF2vYwdgkkjB2t0mFgNRM55fWlhvhOOv/HqX444XFpDaoYDBHksSMLzw
L0EfbUxN0Ghu+SstStkrDgM3Mi0dU63f93WQAifEKd5rXA+NoNLCLkwwk/MX+tQ+
lMjEi5siooFYo1TPPI5LZwdDFZlkZXKMirg0Aqc3TSbzOa/P/GpwPzQZDhPjSSK+
5miM0PnxF9Ug9+ugewaaSDGrFf/7RlWUTmwhuzJp58qUY2LQAdx+l+j1Yumbtzun
VvyrAyfXtsC7U70j4CO3sw7Qza1aqffM9Cs6mJDvG4+9XyxuNupHFOSv1fSPRT56
RZG2JWSDcj5VnCvcE/CO2Fmir43HDOLGofNUnq14COd51QbVDCIPbo9DGSxDOZ6o
HFXzV2DTuFDurIM7zfG0Vk7snYYwGZrBn4rqzwQzXJ9QyhMzU9+85haar8knoXVS
dNMtlhT0VGy4iy4QFlEOXdmQMPw4Jkj3Su/DW39t+DIrwxi1P3jMvTqBzF7s+rGV
5M9iAsekkmdoAzJbYBKHTmewcEuvTfm1QvkTHqXVyDqpZBO1spKcRz9ycgqitjN2
Eg1uKiV4tDLZY+qHDGfzmNBH5ChMUhJFModj3Q6e30NJAJaArXPMUVSJVmCcokMJ
8x/H+JlkgxSzPnLZEbilT7lQzhKzSy7zx/y5P2XsO2ALS98IoPYcKk0qWeRqRUDf
McHzZsUPO9kCc+mT5SrQ3E1SWFJOry1ow+v7HhFDy3WoxIelmEqhR0lEZetCittj
sHaKT/nFJgLoBWVWn530YIjk0uK43ivcP6bYMXge4Pr6SNPA9txM+To0FMl7NMLp
1Ll/m9lIrpns2SPe+OfyHkrPPXMz81OsXPhyQbwwmUJECn63l5XbGlD0FVxEPbxa
xGiXPXpILopNpv1VlCJGn29rgVyiE2worCGd/iwV5YtATpqgkaVkWqNbqJuoPFqv
pRx4iOdLIojcdE4DSkyfzC72QN4stoUzSDPrU9xESielgjjVxFxUa+QZ1obVjejE
7xwEtRIkpKxW/gTDm7/fMVh8J0grF6lqCASK/GUUHx0BiuuzsaBSVeQbPbOHo4H0
tDifZAetk0scRao9nnz0DjnTLA5WoIOISZCxbw9hhKIPmHPG5vqj64G+pYI9Lwag
W2hethJcy5X6TQ26wRvA//GYJokDCQjgJ7GGpBVdy8NxjMNJm6vURum5yd5kAS8j
W0Hq5ftT0C8IbondpSyfyy+PRTMVnAIrGMugiAFhuEcAwEhd1vDwgX9+di95iXSn
irYpUBxxIb3esYUMB2pLogDS2Oh5jEdYjM5OvSU2eq3usdF6T5YU/w7yGF+DUMR2
NQjXN4wfWOs3j7fTopS0dixryyrSaRihnxOXBboFj87IBIFH8EaP42rAzwWyc20x
jSLm7ll5p3RgIHzOKsGntKPLqa6F6JLKI0D7cxCUTO9Xx8mtVaWAWj0jDGeXm3Uk
cAN/txEjQPulBIJx1pTPFy3zkykC0Eixft27YaKIJXhEFSOmiAq1LMvkwrNqDyJE
vNIiVbkIU2QDLE7qv6yqPZkT02NLYkoY/zsjrDj1Y4s/YvJovBXo2Fr9tpG8RZJ0
pDl3uMDFwhHPvA6svU5ZbpWqDBrryxkCBGGUaj50URhRfToFUrjBwCcx0G7rVEEA
CnQVb5MVSkV3AEsw1sgs8tKAEa/x21p19fAS80ksFZWGxZrmkDdGz37GilON+c+Q
TlmQevGGfXBnlSOnnmHRBnxD88xkkzwB9Jz0nmEqWmuEtOVFlbfw9hevVR4Pe5Ph
UJxN3gdjlMbNmmhtTeo2ADhToprBPGpr9P7AzcPe8F0jB3G8wNeNa4WUfEuwod2i
CSF/cm5wjimJ+cHA5/Zq5/c4RhhO5tDARIAbRABEUARKl+vMCZlxGI9mXppsMvi4
k9iQf+KE9OorAvbKyaBeC7YSik/vSCgpI18m/KAeKXJYX01QqOhfJ3mIYbj1xCQ3
Mp1rDH0+K8vcqAC0rGCfgf7HNCe7PBVn6QHJ/rP/cX4jDjhBm3X8kZKUqhCm66bt
US1OxMe17VnjW6tln06U24Xf66E+/c0axqj8ASWpCU4DGM9xw09jyMhgB3w/YC7c
4YZuVNte94HqEIWhYr+Mbo5UB3NuyRUN4F27UCjZM6a7JZfY/82auoon+mCgnXNg
oR56hS2y7IbyGkfJdcjs5ck6U1CFtpcylWNja5QWUNjjrU+jKl3i5ZrQ5bpJJvMe
FJ7kJEne2rHtf3XTajQsFPJ4dksokGJq7sdgSTU2Y2LICkFrGGZaPciDm4yqSZQQ
hLnn0+FrBtgw8/UVyuW/cV+sILVtRc8bbuL2hz8bWh06n9EiQhcLSgsh3SsgXTjM
EmVXc3OJA1dN6RPEABJP/oYUjmyFfVJJrv2KblMlhCkwP9KDyBdsQjtBQHKAokmw
gGNf5SxYGWl6xX7YxQ5gWAZQ/xJrCmZhRlDRRRNUXOCJiAFgyYKeI6ql3Upo/6ID
WiXBMJRM3ebYgFadtzVMqpCrfBx5yfkRhJ4dOXczRPMORfOR0ONOQi6SSzDlkQZv
UK6/NnL9YrZp++76OzVPJxu0Zl3UKCoCQL5KnuOeos/kXfnKDbCvPpBQEzr4+Iby
8gj53eyvbO3hkJ8BlH6y5yJMGCm2h0SEtIebVltHHIaUyCIdd9nDP/9NXJbjKKNw
tWPEu2Y4KYYV/ekBDgZj3k3WkDFOljklwyMcQBUVMufzk2Pkm+vTFCdufgQL5JZ3
ZRC5wkGQ48Y3OFeufxMNwvxC/pttuon/Dv2zsdunHdkuMzzWt5lFUXiPiaYBr1hX
lE3zI0hajHRk8uFta3Ne+wzcWyHMNd5HSq3nJ7jh1lg6CS6UL6j2q5Ao7+ezN1AB
f/blp3zWupVI8BGdhH4foDweahhCs76UDjBFLqWTSim8uAoily8uynWARt4RwQzN
PTRi0IbWxuaa79iGju3vJU60BjAFSA/RPjfWw/Ig4K24MsQhWUAu8Y9gJPY+3ajS
dS0U6EAYzNyfFIECvc5OgxJaaEv5BoGVxgC5cCVlLOyMzV2uLAU2YlPy5YDD+Ip+
DcewiTXZppL4ePsZgkTcCtVCJ7SJmup4lya0LVQAep45tVTqSI2HXorEJBqXLz5o
SyDsLHkEFrJGOO/JOnxGhhwhK1El9Tqw7PQ46Ly3iihdarpfhbYPNMcoYJMJybGg
4S6sAgZWUn8NR73rtnUlh6gwSZjpk7CiFhZUKUKXkfe9mqfwk51WInCvYN5rdP/K
IDCaUlwhkESAavuwPESn10QiMmIgtiVN/rPy+S3b6ufprghvX0j0Jx9Gtmqnl68m
imDhQBAd2hhG3qOuJ1rQ9OWUIew81zBG1xsnCFKT4r9wZ/ost4esQtkGBLFuGclu
oxIjLE8JgGa8AW9aUhOnLP8lCmNn41cc8M2FwIG4R4P4XMAeEumbWRBzqaUv/xPv
GlTzx1xN6g0GG8k4KkgNSc9jOjmOLPDNh57mgdUg20PWAeeOq1oA1tsXWp+0A9tM
JV042OLNLFM9ak0ofqvPiVCsqDNlGKfGiOThU+MXUYNJs8NOYRW78NiiyngK95XP
M7E4TnA2D28mRZh4yLc+eZCgWta3OksGchRie0yaRD+WeHBIRts2MIGwJBceSdck
AFN1IYlxllBf/mOFdnO3RZPGFrxKPQBUXB7+7sAGjdwz3ofXY5EzTCe70zGdio5y
asqCmvYAe/ksUx05cXXYCADdphgmUOpRd9UHC0I/SDeUvPGU7ovhiwAwnk+S7SD1
/slzUV6OiLNXbkQTTHQe2qfDMz0ITihGOfVsKZ/dVa3yV2Y5ug7NkMD3otofbXc9
qJ77Dv2cl31M84moQY3Cd2wizZJxXlYRlPXqZjOnxjUxsBuQMgdvgyScTSj6V7sI
Qmb8CVzdhyQwAn+rHQwZewLJSsmoifJCrPqibfEOjJS39k/3ykOjky5zDSl/g9ch
MJoY1Q3/3bf0OPfLyeEJcxzLTVFn24DrbHgjmH0VIsZdm/8KidRoYjO8Q027UAqF
8O4riNokmmoz1MXEGFjclH4Vmh9yvx4vcoSHAjDgyxYes20vaO/sO3lCduo34kgg
xFF7MyC5M0j5hy2ukfePdTex8ILxvsXtYekXR5GMXQZUnN+KQ4h4UMAMjqDNKp4r
pppZx0v/XUFWtoNiS3b9yvE6Cvfl3FRIWeFyPu5KRbVXT0cEQS+aq7jF/eit/E/v
BouvD2mn1ARbplUrE3pSlMs4NtmjQq3xJhHW7CG9jTVYiOfxWE/K/thOQGRQQX/g
8y+nm6cjigtCO9pdL5d8ByvE9B3TqQaabJoGbL15ecoJAS6zON8bGQx5kslNdlGL
6M42cQOSDikq3doZJl38woUcPvz8MuW4gA6m8ry303+bFCqBkqzchrz97zXelKnE
nGDcbP8Rdr/acE8ffWGvCGTMQGjexnsT8o4O336n03BBgTZF7ghyEziVLjSNwmUb
PjMXbVL8hyUrqYEgLOU+sLtilWc3HdH71Iu1cXlisoAebVz2gWKFKWWfMKKfk0fG
uHsZ7st6Q56+oX/des13ljZLNCgNHaubKJZcFxFbcQyEUk54CHi8cPcngZIyO1Ke
/6TohVnnE98SRktnWjm2G0u8uBEfnX8XMbjmVEkfkXklCczZiYtFzLzIfkkDKfyf
/qV5A3u7TDfcHv4reIAnJG55ZI+i3SqlMZE0vEk1iZgl1/DguHhAHqJFc96qVKhb
D7NMhIv/Oyox48Pecbi5WZN8erwUNOYb2pMe3ebVaB/j+zr72L9fZqlHyQjjkMuF
9/Cb/w9i7eZly3a2Kkguofc2VKPAnFeqoZOGstrZCv2lGioiVawG9S3BKBet4Qsw
sBJ8EoCYigNZpi2m4yP50YY4kSvfwmZg36dMKyK5CUuSBFlrdTzdqy2KVH/rgc2N
mj41t/xGKP/l03RUUU2Eada0w73jXksmUkdxzRj+6mjPvnyzrFPZ+IOH22l5sB04
woYnFcuYqklwm5wKZb0xbVy3xFvMaxSZv8RiNJK//8qcXUB44XqWQy583b8Dl4sV
c5w/AtYdEI5A90zHz+QoLc4aH903gvFQBMw1Ja946KymRcryMdi3bWGKMHP+lxcq
NLpBedoQjj11ixJO1OR+UDjC8kJ2NQAEy1Yzvn5VTXBtmUP91PLUSwiwngYmul9Q
tSgs9aSLBjg4zjb8cbc/PqyyUEmm1A/3/IuirMajgMz589UcHK2L3lpNFeWdD4zO
qY9Qqi+PfYrVUx0opOH6xSXnf2Dox1mO9fP/xJuq2woRU5jzafBUjPiP3rz2uJuW
nH0KkzNYMZ4SXzRS0KKDlqM88LxxL2ya802rbmdj9cmBZXALV3RZC2E/SeGUR9RA
gk6yh+VnxTZfZL6ebujJdnUGXOJqGb3PbCrrbBTLURNrj9NuDeMJygDMYBOGvJqz
HWuUhpqaDnk5HwabrVuN/Ao4bpKi82sf54vWU/Gvpfyqbr9Xw2BqMOb5CS3Cea2E
PRBdpjHVd9Ei8oDKPOB9v4oDSvFa/HOgrjKan1Lt6QPqJ+s+rAeqF5YDm9hVl2ZS
I3uZulnlLMVtYk1V83h/cLVMGNN+/ywJMQxLEJWfefUrk36JegRBDTIIJEMzkC6X
8z5SifrtdD0l6/m6RH2HfHsNCDFvuRZqBIbHvSC9YQynRAwyLVVRylPeElNZc6Iz
2Nd5Qnbk9zsI8Noq/Snw6FlHPDK2P+XJjz6OAwSzL7ciiKLof4ooLiw8r0WednRC
5DmIabcfGMTpIyER7jbrWAIqZ50w6Lrw8GY7qEdX0Mmhg6kgdAtetL4zbfyuem8Z
wHpb1lBvsjB9/ZHvVvOXenC86Hg/6Y2SRiH5vzBRrvyx7vboJ1ov/MEe+bkMCim7
wOtzua0bKUOpZosruoKL/PsHZ8zVayGHVo/XsZHcBp3L/YG8nFFKBMnTXz9UfAxF
K3fZi/t9ySU/afupdH17vSfRed0WnSH91Wb6xlJ4qucHbUx5GUJonVGBsSwFal/Y
hrykT/8/CrgNObb2qvMPRG2K4ex+w1yVQSyJ+kQ8ytmbMeYu9EFGxPhGdv+c55CR
xttNV2NlCt8KwyinSSawtRwRTEdT7jSjETBv1QTE9guJ6J1wNwn5Yw5L0Yqfx/3c
ANJN2LF8V+F7vYilbRY9Czg3U4l2Y59DbexCToQeP8YtIdoA+dXAFNcG0moi+Lew
Ds9tQICUCzmVoUvBJpNeNwD248URbO2qeGCO0nVA6tyOhz6L/bVTomUDCxvgG8Lf
6UbEkxCjE2fJjnwY1R/bi+Fpwnm1ZzP7X6DaoLBrRkjpava1vFgDmAxWPLzfjWL1
AMU5hGwu2lcny05lfP+HIa2qrHWIQbwIiq+UIgC7+iUHk/KFAcEiG8lGSI45EV08
0ixTN1aHDc6Im28FSlptpQJvnyJBqtxdWaaqdEQ70t6PUsiMGosdbAUE3AB/XmKP
GLwWtb5sM0W6wlIDZTVB6ek5Mt8ewNnpVGmJkyqXTP8j3Ec8Lc7oCjEZcx7bEJmn
hy6i3n53gHZLqczJxwkzjJ4pjIlQDLPhuVWFmibj5lEfpAXlscTE74exi5c94JUT
wR/XjIRpQzPN9y01fl31pbnFPyKUneQzl+8CIohLUqFnBaX8A1cgDJWUD0nCDWiZ
Mrl1ymGxV38oPeSvx0l3TTCgXb4oHYqlJUwbquQ1lv1pYjwxM1TnoX2q4c3RHb0e
BYec+usMS/t5FZRpcoqoKcQYtTSbZAoTPa946UagesRiBETv6mi/6hV1pCQxXM4J
vg8fR/lhWorg478mSqZLuDEagj08VEFLnXQe9YcQog/2xJEVeAAApH2OIS4/5lzG
Jl/29bLU94xZGdtZK/FuTIOL1CguVnd20r2sfBJAnp/SsJuQ1CKoCwUKOT10h8g3
CGWKvZaSREnoPuWtQqYOYXtUYaYYiPnrw7grVlzYt8jHTAZjaylLLbJE/hbYbHTR
ngC5D9hzXQI3bOB/vmX1Ss4Q5ghJNkiOB3cBvMPTBmRKWo7KY6RLpBEaJSMqduFg
fnH1WFT1KKIgpPUqhvB5cJkjat1K0utHGaH6clirScQFCf/sZWtptkbc5JgCA6VI
ua/Vxrg8JTX3u12qfHMNtGictD5Xy+ZLBUj946TxkLGmOCEkjPtuFtmKCCNkGoXN
hHmKB2VWDF7lRGMh0XCnHu4IjmL6bgkdaKPvRfvNYVRw+dNSg5NYohqSUnIBkLGa
l8+N3ALlt5uDqqNcqzx+rR/fyqXCZK6YDRflKWIGseTVgIy8yPkZ4plq0br4zaVC
ty1D6OTnniromWSvAzNwvkaPR9TmXX2knoXHM2PPi4Aiw19yhVll/N1jyfE/lRJw
wBQP4a2m9o8HmH3SYGRO9LkOI6/ZT2D7nakAJ9JFlJ+fNJ9vlSFpYkHTxPlrP2cm
xr24/SmeLqwZse4TXnb9t6qq+1HwbmaBJrrOuHnGqEbAcevRof8SUPzBUgCdryTV
63MHVyuVXUQXIiFmr5/8NTGqErM0XFYQK644A6Lyb/mB8z+9CfJTLs87T70DUBfs
C8LVbwxeeWCZ+VAeiQTS6oL5YVnpD6x5dRJwyeJGdXQI2KtwqjQtndzqu1wAgAXq
a5wgvDoK4+oMvmfoo+Sz7XTBwdgv++EMepnb2aDyFIjZgqJDwHU0DtLZCVBzIMzc
gAsFthw5gaQZ6vjFbM/B2YuIifyqIRWgKi3RxrQuh1GXgG44AH4nZhgI3rCUaUwf
pc1aqPZztOFCjzDHDu169FQiBhTQxj3EkJSYwxqHI8qAiXoclgi4Kw4UOq3/bPfd
PTciLwx9EakK9uM+R4SjnSmrYH//b0KwRRAdIw3FiAsq3Y+Zy9bzNM+PlSMORt2C
fQbE6ETDYLj23SGDKvJSS6kT6iqatjrEcH4csA9aiZ6Ru6jJorlci5rGoPSuubca
YLVURcg7hh5UQh9JPUVi2xTR72AQwJ7MlvzDjL2y8JS/rb/r5kulM30sAWnEmyAK
bAwdJOB3xgWS397daSTxTCHIeU0v/x9NWKFIauDZjqZYXMrRoGPG+oSLq9rmcx7N
jE49eo1IeggE/jC/Yr4ftPA2WTMClhcBph247J1N9G0=
`protect END_PROTECTED
