`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK2b2Tck39Gi4Q96WGe/+9lEwzc/zU86FdN+3Y+p+IKE
rVUI+DoK5I49OUZ4qCCtitmNyK/S1IHBBCANpIi6A7ITcVa8jzueT22Q/xRc1sZr
IGVStm3Pl2BkJ4BXzhnJY26xn3toaRv9MjsWwgqTR0alyPXRmjEU8gbyJW5qdhfr
Q6IS3G8ys2dx76wdrvZt03NFjoDXrPBz1FT66nuBCI86T84P8JIIteTp+XUWpmnd
JV2aoU/9yS/9wSmdrfjstXkK4PauYYujynqzeQUhq85u23eJMVpt0HUhmrmbEfTl
VamqKrDwZg2JdPDel4oXE6KRk6E0/RaUgELIKz5WZI3K+z2NiQVYoGhmclcq6c5I
5OIc0HuEf44AR1xkxw90xwg8RI91CpI1pkIz5i6h2T3G5t+J/62OuxTt12ZLsxhP
jgR5Vu7+Plh2GADJ9roEi62O1U34RIth2O4s40AVGN+lcH9D7NPxuIAYKlBdhv6Q
QpqmJBukp0ETpy1Y5xwF1TGc9Rio1VoCeeDJCpuDRuHW07DazYr2zs1UijGP3NXW
`protect END_PROTECTED
