`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveByg3E9zrUhBB6IY9paBL2ihDGPcvDWecOXw54MMiMZw
39Wm93DswDbhXC7hEYrr74PbGeyerbLnl1RVjD4DpU3t9OSuEJHM+/VMl78h0jhM
ySFv5WFsG4xJcElkiIcw5WcRVZ+c31St3hd4AsvO/iplLm3iXXjx+sMuF0hYrqCD
/3FCsLKj4FfG1EmKf53itWEz4qrlfWa4cd7KZIjCFMz8+Rl51OMqbbTY0KA7bgNE
gusO2LiuZtLC6SFYP9L3XPARQMxwYd3tBbN8IDo5/RZ/+JUyG2E4jUl0Nu51Y715
BwE3w8do+nNBNI4UbFhngSJ6Rr+0p5D7eEeeZcDO7/QyZiR+Nt6kwW2abLABlFat
`protect END_PROTECTED
