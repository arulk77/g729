`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4z8fPEvRcAmGj6imGTBRSy/uegTYMsHEG00nTvqU21Gq
3QKr7c68KNIPduwEv6S9iB+gkx2QKD4QuE56UK1+wvUnq2bGA4zXS46Ul534Paz2
sz4sRIddlilm/+iKhCZWH+N1Wft/gjQjPSCQZ5e8jlfZH24kbUzIe6XSuz0dC0tW
mkBfERcsqjUUR58qS6wBLPJj4w52KUEGqc2n/JbRpi8=
`protect END_PROTECTED
