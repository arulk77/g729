`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveECnVZFWiBCxPIaCTSYSQ2pt9nF9OT+9l0w8dwW3F8yl
/VWthHtBgZPTnFo48WuPRY9WTbJf16t2a/Y0e6Mb0ygMxXm0P1jAdZOkYhDiMc83
qTXDNtK7u+pdJeFgOB7HdQw5bqcZgaYVXjuN+AXD4/KMG9vxBUObH0qSl9Zt+w8h
k5qvWnmEWTLjhNU0kkSC06qYRHGXhl1jUbT/qvg7eiN1sgUpSYAe3bQFP5tDU8SW
k5pxrroPRdiWnxK2dszsmYgxuDONk85s4TPilPhQNUvVQk9bNSHREBvSpSTgffQm
N67p8IA3MbIlyb0kylODItKiXb2G3Gu9Q+uonuIn8S+DI41nIwTp/SfjkANpFI1Y
`protect END_PROTECTED
