`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN6IWIRzW0MWtkScZ8A6fg8kVbOMCIwIXCadylFHMQ2QH
veAj3SC0YnqrOzoic1u6yHDovNhOvNOblfgrc2GoaPYPHvRlnEq5M8/zJKadbzEO
hqK2ilRRZo39rc343x5oHuRYISL/DRUz/HUY099M7R0Pl+9e7TsQC9Xv52y/5RDV
Bwydx6RX7iC6twUn1ubhO9z0etaFUwQqxKvLJDCckKTaJg42KvegvaP8vbp86Zps
2XvdyV/5QWYy33vE0k6T7gFCnf/w0qqaJiCJPqSCoeq6zh14AoPAqMn8wXEZVgPu
ZVIRau6qS1YyeR4FNTWlVRyvtkTay7xTavdshpUdiB0UORwGWmBoJx1adTafACEm
6RzckyvIv8P9U41+I5CQ740LTezx8ax9xAjvAGLC+WenAnXQF4h+6sOr1qcbxjQJ
hx+OtCLUmEmJs3dyAM2CBdiAd3aqVYIBws3S139UXd4KxyEFtQk7nBHq2vmVkVeU
tsahjZkPhmWgWMt2fNNQihUHDjehlmzdE/HwMuJMEFKbhBv/Npl2OQ8ETgZIKzma
/xNcKS8PEUugkewt+Nd1H/N2vVNqbxf4D5X+l+QfNl6tzFOY0msX0xTdgwTd2ryf
sj7pbAHNaRB2U6cdR5vbXVN6kiCNuZz+gm+NXSQBz1hyyMcCu7VZkoRFCMI4enBA
r+veyHOyLXSes+z5BRfN1EKXwxtE6nl1r8ZrhH1u+hgjHNmJ/cWDKNN3XnQ7T4WP
5uoSjAze5iyrYLOJqgqE/12Y+TQdD9Ij65MpCZ3EP0XN9gIfIafgB9/Qc+CWHkt5
hO7n0SInpq8f9CThEdTMuwbXXTSjEjxppSJB9AOtfC5pgEgCMRMXjdFRMvn+ALVp
HCTgC24i375AK6mtZkQe1J/1N+fUz6hCHiWF543SkzAcJGt4urdCf7KV+LdWkShh
nt+TC2FxC5yRFK3XuzJKYq3p2YsdIJoOLRp2h/iBWpFw74vghxcLr9dXD4W1o1pB
DmDwN+9ihCBZd5KWNjuQMKjSmUJSFjl8+2m/R0MSG3XOPAKEG4CK4Qyf27Z5Emdu
7OwgqxN4WpJ4YdjmBF/MUlIlLk7eGjIVa6RQvvPY3DDkBMg0+UazaAyljj+X7wAU
xDFUd4cFi7jIQB1ujLTGjeC0Dy0GeIVRtC09kIFYCsgoznqysnPVJW9JSajuGXWY
OFZ6Jre0rAlsaOMicoYUZij+nll2RO3kXpEhIplBnoIv+UCM8SRZAUaWCmIrlFTq
VDR1VaZdytq0cag4/4Z3B349gvumHwr4jkC53t+86trhOz6OA90EuM69Yy16UsgZ
utXknf6lHI604QtbBG0AOQNWjnDBsDyPaK1tYO8T0vuywb1v3kf1e8lbF2yTgb3H
izUm/+jeDu9jXtsxnLLuqQ==
`protect END_PROTECTED
