`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNzSF5srE7ghsyPp1MjvazCGDIRMnC+rNi5zIoNT2xxUi
Iohl532BBVkPXv7M0UV7Em5jk5JR5XQF/3ZcFvAMN1X/+a5MKi1RcFld8XIBON8+
CnCK7qXW/H7g1PHShQ2uQgjfLQ5Y+Epwd/xfWsTY3S2oBhZeXK0ErWBznd83fkFI
vPTWEbl6NvRPnFg5wLApqhZ7BUsaNyCmf7iQ8A5MEFDzoVpN6UVPljeN8r4IUmi4
`protect END_PROTECTED
