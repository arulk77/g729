`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aSU7gCO6gmEeQlfO+sg6bqCHXtUujflOaRr5Cp4+FQGV
IkyFwIfoIe9MRu1oEPyCupgdeLg8OFk68urbwkl1LEFxKsm8c/GcVYzPgWfeXEek
fGqTHMCirxxi41ucPxVS+34GxsfA65cC/ekBMIjQAF4cMMgV+HlI7b8DmBLwr2hJ
Won8QsBhcwzEa9Xp/IcvSxtdW2bL7itXShpfk6r3wglR2BbUoQDtHxIF+M15rNzX
qXKFJxNeyNr/e2zvpmiIYd1yKvM6t6EoKMky+ss8+ogmtcyAS0mOetwCMv9DO9EK
VqnLGHthlsqxci4tJNaGPD6Oqn2uSA+pfYiPvnnuna0JAqqfsEjYF2dAv/AYiSeX
+Wf7klCe1HlVrhtbPugOfWtcFpltgq6FbgSYnaUoPHTW4b2OzZS6/K9NZdmyzNBY
V1nHpBeq0TAtxGjlmPZNqKYzOEYMjJQWIoCCGUqGN2ZwiqBETo94kcuZCmma2FE3
C+PkqzQpMQIDmVIBYJQQNK0KCsu6E4mANkMYmYcGViU8kXYFm3EBbWsT7dcwgXV2
/JH29AwwqAiZYqwpond51QKiKmaBZgyAyb8+rryzT4bnh0quDHQl41ciH41ozqpT
hi2rdp6cD3wITlzQFGwoD/Uge3w+150lBhAZ70HFZcPiduo6IGUJ6VMQ9R6kw4zZ
UTJ5oFLZFww9tO0S1uYkRXVPbahqjhbgeurhZxkOTxO5/ubS5warGMT+Zc1c4795
U1QE70uBhXNnu0/uphfDrgvqHXklH12QrzJiyqYJG7mJ/5CKfoGm7wFhILHk1t3I
9/uaRRX/IxcoVh+m9ymqoDYObVhVRJrgvk96G/ewOPBlytz2tJ5Za5M1moN0JLGk
L0J9Lc2rWbGMyMz70EIpWZzRE2Rz3GgOfDpcbDN8VxKs6xMS9hngD6RFkswANgWB
s8LI1o4PQ95OmOPloNpi0Qv1pznrR6UCQrE4cO/IASUA7pAYITzr/7ROMK3NYXfa
mUWV/7EYmDygzg7/i/5mIS5qeFq6z/XtsDE4K44PmregupWGcaOJ6+xkacRIqZlg
g+8CXzaY7WYyhr2g17J6orUH4YmqQI85tHBKq4d9djvfyFoBAi2bubAQh1zIcaBl
0JUqiWpHXEUunDMEcxnFaw2k5MZs+vM9pm3Z2rb+g2wwXjbhwKlld6QhKryWoW3d
iXJL9EhDYFKk+nQ0/EuUdDkYmnS0HxblbHQI0yro5e/8yZ2a7nxK6VU7xuGGr5hF
Uq02cEnuchAbegTYLBR/9uCSEfcBdax1+DNiyhlB4gWY14KfhA1hTQRF/+YOFw8o
MIQEioV9vHbnWebYCgY0bPoRofaSh9nqMzPA2YvrPu5UBpyVrNEwXihIIFKCgNlZ
D8rii7ZlXJmdka19jyXG8KcDGDT7BaRYYoFP46dGdJ5iMlw4Uc+r3oGRkhJWmmZR
bn3+cD4b1o2mkXM+6jKvd9dQSYvip3VFthMS7yVE6G4=
`protect END_PROTECTED
