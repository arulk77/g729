`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOTrXj7Fr9KcNDYgLB7MKO5AMEeAOXx2fYwGrtthkCgi
WQpGHpe9qUAFVSsGTfVwBqG4EPfaYg6g/cECyVVpW3XEcrxUua273scKNA9ZTkCs
fkyZhMjC2rHUmW810mrcDmvikxTNelhnSV1fvjw7cG/b0Grkj8qLH80BhO3sAbLi
7Sj/480Fos4LL4YXEiKJDxgwDdEbrBWSSwoN7b/H/82FY0OxA1MltywrjrVHgNRq
rByJK4stQQ1jloiUuE9eOepRnBL8uoJrf2YHzgIdyj0E0FHazXfsA08Gh73ST/xl
6uKKxuTwfr2MjUWRp7CQ3gtT+fOxZpqe/G2XSB2y5xIhMeJH9Se/KBbT7ZLBmTxg
TZOr1qkX0EViqscq0UbNohuTrihQ5Y7kixw9Gu2uDEqHTDHkEK9AFKyR0B/DHS5r
bBNxTl9lN3nRxCyheOwgyuM6nc3ZizX7+JhFOSE1VjNidk7qIgQaNJ9p5jbxisAK
ely667yAvj8Qms+XcPlOUgBkE3OZdGO/9xe2XClIx8ciGIxONRiFRUcbeBt8fcac
oQOaIepJcTt+ifXVEcxwSqNijUVx3oMhqE0IE4xN2/AGeUWxVaSaxPFy0G5+bnBA
`protect END_PROTECTED
