`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+DqtKcBnPOMlcv86EOfKmSESiZaWhbNqX/jqtaAu5+H
7KTeLiQ1TRKKVhcUKSiLNcbdQkj22ctvlr3mbgR1mcp6vf0m1ggHe/pI355oedz3
E5Fl1KD5vvkFvgkIFVOTrPnL3IjEeLAR5YCVzaBfVfCzLbMKk9u9LLiPVLP4twqe
t1FgbxGdxo1cp1e+9Xb2sJyCIohFf1EyFATeM+iSsOvuoOcMwodEx7g+st20UmcJ
2xvnk0yCJqTkpW91jx2NZSmiz7g61rfSI+sHzq9ejA0=
`protect END_PROTECTED
