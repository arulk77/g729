`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMGaQOcL97iO9JCpvwefCynkaMmBllABoRBKTDRD77fa
e4g6fkMcH1LRvOorJ9LFiyyz+YU7+1Bhm+od8zZDNkiU0zi5RVB6MSOiF0gydKh7
U9mJ/ygWcIWKSAFyWeHUrnnj6OoDCN5126dvgUBj4kpxxdGXQ1s1StmHnHmwsyMs
pxOx8LkSgasajdphHm6X9cePiNKjv0ZgXTVw+BibwdE6xHRy23129/U7XDuy8qz6
WiOzHCEhHoaGMdDT9nMkIvrVxAUML5bul/99SV4iANRINNiSJk0exeuNpi6lAeN5
LXh0GHMrjwc15zrxjaN1Z2R8bA9vXuUWf17xt/6qstDMBvCBcs89aU3cxy0Va0E6
3+xAIY4jOpgZuj1YGnEBw6AYV9grd4l2wM8Cz1QDPAd5AiifDIS+iBnTDqI30p1z
VCpLbvfHt6DZvFJf7px2F296qecBSNK9oD3x7xaKGh2R7M5DR+Q4IH8qC7cD+z7C
YEryBbeqHwroB3kN1TNunZxOkMxGv3/OUl0gXNiwonjvUziqlhNSAxcrqAXXpH8p
n9uYATF8M3Lu/TnzNOPUl95F/Ru60GpfnXoHrE3gYGJqEwjmKnslU8G2tC8hwH9A
appB3RWglCnu1tB+RMG+Rcn3tPfIp0AM/UYK1plPtDSYrhsW0FgtEOs8bNC4sXoG
`protect END_PROTECTED
