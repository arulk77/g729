`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44xHfxNOM6ZYL+fGCzpA90oY6fxj3f8txYrsKsWA63Dv
1ZwX0DAIVIg3d48UYxX/JXbmv8CX5WjQSbXEA5zVQfNvB5oCUw4rngg3iuw618tM
UxJMXvKd7WkWmRS87ogxv8EO9xyHHTqSFuAX+nVlB4ycq4vJO4x+2+wY4Y4PRjCt
KPrBYyDTPd6rD8lNlzY55o3jlXjeFIPymBhTybhA6GEyLyClRQWUp6a1zD7N70JR
HPKmpOD98vxGQUxjC/L8Z37RU8QiiKoGyuEX90uAnvju6qZvuFndEZZP/TWql29h
buIOiV8zdSM0xI8M7YUmu04JiF7QXOS+J8oiqyay3fc97rsxPApWPedPtNrJvzCn
Lv7394Mgoqgkr9m6a/NscXtesM+mHcChTZ1IgPnXpPNtSdOD1y9vyi4+sOWWNqWD
80B/JhviJbcc1q09PjYA8abBr/YetpIDmtd2TWBpZa+XiNcdbgDFAwwYj+0IQoao
hUtZM7aiI5UxpJc74+zXo4CUbfKCoSAxBrm9TFhi+/Kl1DnDUu1eS5N/eLqLqFZe
5gt86ltmhpjR7ES2x7y9cS+N359uJH8VYR6sMuQ5HHLGPChBQvzkPD7oUpvboEOI
`protect END_PROTECTED
