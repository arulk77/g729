`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
radqBApGPVupM/hLSvtAMhaO5c6mKcEf6tg/LLZe/yb0tENjsQE3Lvco0vsYVLnF
m3eF/R05Bb0kVgZSvJo4RCwOMn2Adu4TN9zHdLf+vFdevDpFJWu6K2RhYGydYW90
P0VCbHy5EWlL9vtt7WcVENvJJrFZW8DqCTzSgg77Pkhd0i89W5cFLVA2Vb+xIxwF
a4VPuzPxjj0JqJoBR0gsSf8tn8V36o8DRS2Jc0yGfkk6FDWskVtcQ5FvWVVyouZO
3Umr/EnFO6R2HcNgQhwM6nRYga/yofuifZr6kTTr+ajjxpWHQpvMMLW5vBbjUkRQ
pSC/sfxMUUiWbLCdeSa7RwcrHPpSfwYjILnG1EF/xuIblSM2LZkk0BRLNDwGz3ph
b+HddRWusOSks+ceej7TnGWU57k7ueeT41zsz3fZqx3ctZ7U+P4wMFaSrfwOaiPz
jEudVepfwfYwZJRoydv1E2KFjI8iftzxX9RLacqSltXjDFDyxZ1xiSP1ZhPpxQRe
loF5PVNc1Gd4FegIC3nc0fzMSPk49MgAP1e6wRCn3uUAv8fA57kmF+aUTVH6XVIB
Vm7Lm6vNYCPjoDbN2gl+Uyvx9SJWspMmKHhjYBjVGikYtnnn5NjWPnR2Zht4vcey
`protect END_PROTECTED
