`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42DLa8Lx12ua0uFA8BtH/DKMGUUwqVKKrhjRms49Nmdp
XKnw+BrB02UlItolaI4r48uVUcOv4Shyz7mAWq3D86gSC4wGPIJ7nliSLly5PO01
LV0uFb+x8FHNLsvabisRToLYj0ZxvXmvsSnI8oxJtQaQOaLHv9NfPVEG+gKPdLYr
3uL81mw6xW/XdrlnjQtNb2AxGHthdnEBV4aquPxwcTVQnLTkco3sESweghHcbw06
Y4hFay+Y57gT6Fv6rHaoTWvOeRE/1T/vYXutr8y7Q3H5OQ4B0LR0OMa77CWiDan3
Li0MP3jDqJAkIGYBnZ2DZP2tNHBsrZDhblkg7Y96C+/G99XGAEs2YvKzy4bspMXx
laekukUMKmd3NDPP9LVvHA==
`protect END_PROTECTED
