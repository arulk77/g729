`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN+ol2YQPQNRQK5Cfa5VPVtMegwZZI/L65ORMaGSYraR
AnxXVx6OCcXy9ix8jeHDhsry4RDYySytm+1YE3gcWTrC/UtfC+/83Drvvkip7TgK
HBdCONB+5w+IZY6beBpwAw9nx1ZFAxVCv8MrMbkhC94IO9tL+uXjow65DEpWG3Ln
d32AVcqOhRt4OX63jeWyG/ZViDQA6dyKeKHCdtw9UhRpAwGL8R0yvd3W4v/cBCmd
7f21ga8zTXGgmGHhj0qd4nzJ3c0hnB+AkQrQGQQNa1EjP9dyI5x/vMOtZWbI44o6
1JPnNoJPRV+CYULzQjDTR0XDGeTSui8OFhqeyNpedPDW6R4OFeoQOScGmcZyBYho
oF7s+YyKU1aipa+QOlrZ7Lzp0NtReR60ICJRjW14kZZoV5M48ngBvp4tyqrzJv4r
F5cQ2zC+XTJ6R+wy7toS6RDQlen+I3CkeObATFmCCegva6ulX6DaPQRp+SM9xJVL
g8FCxoR/4uU2CgJa5EGZtZRvdbc/LHkqrjcbXuaNfAx2lmX9fcnWSejry/RbA3To
HbI2afxMS2iVzhjambVMhOsMBnVYO6sOWrZqgF+yJNCO7FjxlekbwSLPeHtDsOsd
BDE4xdlMyFXdsOmgOD48z7fgrnTUFPB4E8g70NfzSeFhpD4QrJcxVSE0z2w/eEMC
`protect END_PROTECTED
