`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAfOAG25IYPX1gHATGSGGl/FZWssa0PAaX5vMvNVyYWfE
en4BsM4Traq59FiZDrSAHsNrEldPI2un4cpToz7mYLLTB92SDiiXA6qqZhMwP5de
i0Vcrr+KyzRO+ewW4xH7KYpnoThj2HDbZFkNWkzEiFGLJvzILC+CfQf8ePuGor+N
HU2gohivSZlIMegdBkHtnHW6kdyIQHbtayp40tmh66ov9TjVESWNog59/iDJqrsk
QjWqV1W+qmxHWxMmNhCoHaf7CFr4Tx+kODSfHpkCOo+yvOzTadJlOFDtCVMOnwNx
DrLAppEVyKT6JJGN24qca6HIO46DL40sJx8aJaZVu2AaVH3JxSeMjHR49bFR4FSd
r0aIl1tMzvaUX3Q7K78cxqWUHQWrO8ULUzKmvmql3OERXjne3VbUrVMbQe1hTTpp
KhF0GqFRD7DIUbkYDxh5BJ3btvZiDRQ9i+MuRO38hLs=
`protect END_PROTECTED
