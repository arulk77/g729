`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
xr++t7uBkrZm26Q7QH1dmgb0Um6Vfn/8AsYyoaqcFjyKLXAN80VUMHoJGvwr7/BS
qfu0sJd5aa3Ykx5gsUcBnHIv37gRMIkQOcCCoFGGaRoPeC8CkO5CALSf63cLsSOu
Mhe2Ab9d0KljL3AgJHkjUw1QQvdtanfT4j2GmhKr1H3CaMoIaemDjrY50WSGBTW6
`protect END_PROTECTED
