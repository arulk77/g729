`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aSdSbgj1ItHsVlr0i7Fq0HfPxFpEU9jXgt66kiADojku
cYzhUUHadtszAa/fmkeMmEYBz4XvO0/pOKQT0h0234bgi4PgebkoXAw5ev9Io7yo
zQT44Fs47NMnO87owdqFABMX9Tu1188CR1naEpzc9LI0eToOqS5u+QYyGy6/mepc
qsdnErPxhXV+W0TvRiwctj1dsrFRWYQWU0LndbyKXk5wXxbPyYSYunGeDcOeYZFb
3pdVQtnRjXKvjWqpz74Y2ey++ED9spbQPpZ+6eO7kcrCL9L/YVUoTkUVXFErjLlR
wqNxsPqAxuxEeYDLaoM7hm2fMEhfNYJdUJ3kIj+MCGoTuCgLHOBTRR8V/NT60Lu1
QXw3HwW4s8Oqq0XK4253j5yuYblSQjbR0SuFORFITCNMMQLbFyqU/CB4GbagrF3I
sts8ygcI94lnHHfBzEFLC0ir4lyVZlx/GaeGpwYBi1CCxJuBFVByNHYkEOGveE6C
3geaizF/k5vL8gp5OOBnWaJEJHIRSyAFtdM/MFDkPAdeo0H4MxNnAePKC3YTqYPq
iBZwVP/OM/Sf8xBNHsi7KlqqHPtU+h4g0wrMkuq9l7QTOlnPajynAiaGt3+DyZkM
zBLDP9bZtdsTxiNO4uXqC4dD13e1jrtZ32dzp4A9bec=
`protect END_PROTECTED
