`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDzJQAIrkrIdBuqrgz4mGi70DDWOmr2ne9R5aTimygoS
zstIJoUi4bKIkPuhfzyqMEgmDENSDBj3IfL7oSd78yYYGzSsAFVpNWwy9vug7J4C
+tRFTWtU1C1vF8qEEUoErt1tR3MbHzJKa1aTYSoyWl3yEVz0xPJEctdwRMzdynPo
o3kF+fcmLjTa8k7yoFlPvLg5wAb/tdjxzd+DZE/jtiaf0D91xLWf0JJALVQfRc1Y
EFSvKjfp7N2gVKYsDS4uwDMjs0hnLT2B8untcEZLQ3UzyhZlKZKxGl7zHKEL2aC+
ji+8wfvA/SQ7GGH2Il6K2HgpWEMITz2HPLQZ/Jc7q2OLnc0+OzBK1DNjqTBd5UmP
gLPiHDKF71ItKl2bhKAiuS+poVFzT1wpTytp4ImXkzsvqKXPDSi6/s5SeSMcsoRb
xJdgbpHWVN7WOcuvqzzobHZ1vQuO2hEgUMhTlK/GqkMq1SUmlkH3EAjZpg5WEFG9
cJtrBOlPaB6+FQtsA9IwmFuUTylEN+gdKdmUNGi+XEfr0+4IZ83iMIbRqkew2KKe
TzIdrGEWINb6F7oFba8pPEEw1OL9vUbR80zJde2hucWtg9a7HCVImKOLbNHFtNR+
whk2lPfckYP4ZfRH3eQy05zBUXynp9gk4O5AowQj+12KXZzaprR9QLR+d2h22bTx
`protect END_PROTECTED
