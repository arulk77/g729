library verilog;
use verilog.vl_types.all;
entity GTXE2_CHANNEL is
    generic(
        ALIGN_COMMA_DOUBLE: string  := "FALSE";
        ALIGN_COMMA_ENABLE: integer := 127;
        ALIGN_COMMA_WORD: integer := 1;
        ALIGN_MCOMMA_DET: string  := "TRUE";
        ALIGN_MCOMMA_VALUE: integer := 643;
        ALIGN_PCOMMA_DET: string  := "TRUE";
        ALIGN_PCOMMA_VALUE: integer := 380;
        CBCC_DATA_SOURCE_SEL: string  := "DECODED";
        CHAN_BOND_KEEP_ALIGN: string  := "FALSE";
        CHAN_BOND_MAX_SKEW: integer := 7;
        CHAN_BOND_SEQ_1_1: integer := 380;
        CHAN_BOND_SEQ_1_2: integer := 0;
        CHAN_BOND_SEQ_1_3: integer := 0;
        CHAN_BOND_SEQ_1_4: integer := 0;
        CHAN_BOND_SEQ_1_ENABLE: integer := 15;
        CHAN_BOND_SEQ_2_1: integer := 256;
        CHAN_BOND_SEQ_2_2: integer := 256;
        CHAN_BOND_SEQ_2_3: integer := 256;
        CHAN_BOND_SEQ_2_4: integer := 256;
        CHAN_BOND_SEQ_2_ENABLE: integer := 15;
        CHAN_BOND_SEQ_2_USE: string  := "FALSE";
        CHAN_BOND_SEQ_LEN: integer := 1;
        CLK_CORRECT_USE : string  := "TRUE";
        CLK_COR_KEEP_IDLE: string  := "FALSE";
        CLK_COR_MAX_LAT : integer := 20;
        CLK_COR_MIN_LAT : integer := 18;
        CLK_COR_PRECEDENCE: string  := "TRUE";
        CLK_COR_REPEAT_WAIT: integer := 0;
        CLK_COR_SEQ_1_1 : integer := 284;
        CLK_COR_SEQ_1_2 : integer := 0;
        CLK_COR_SEQ_1_3 : integer := 0;
        CLK_COR_SEQ_1_4 : integer := 0;
        CLK_COR_SEQ_1_ENABLE: integer := 15;
        CLK_COR_SEQ_2_1 : integer := 256;
        CLK_COR_SEQ_2_2 : integer := 256;
        CLK_COR_SEQ_2_3 : integer := 256;
        CLK_COR_SEQ_2_4 : integer := 256;
        CLK_COR_SEQ_2_ENABLE: integer := 15;
        CLK_COR_SEQ_2_USE: string  := "FALSE";
        CLK_COR_SEQ_LEN : integer := 1;
        CPLL_CFG        : integer := 11536344;
        CPLL_FBDIV      : integer := 4;
        CPLL_FBDIV_45   : integer := 5;
        CPLL_INIT_CFG   : integer := 30;
        CPLL_LOCK_CFG   : integer := 488;
        CPLL_REFCLK_DIV : integer := 1;
        DEC_MCOMMA_DETECT: string  := "TRUE";
        DEC_PCOMMA_DETECT: string  := "TRUE";
        DEC_VALID_COMMA_ONLY: string  := "TRUE";
        DMONITOR_CFG    : integer := 2560;
        ES_CONTROL      : integer := 0;
        ES_ERRDET_EN    : string  := "FALSE";
        ES_EYE_SCAN_EN  : string  := "FALSE";
        ES_HORZ_OFFSET  : integer := 0;
        ES_PMA_CFG      : integer := 0;
        ES_PRESCALE     : integer := 0;
        ES_QUALIFIER    : integer := 0;
        ES_QUAL_MASK    : integer := 0;
        ES_SDATA_MASK   : integer := 0;
        ES_VERT_OFFSET  : integer := 0;
        FTS_DESKEW_SEQ_ENABLE: integer := 15;
        FTS_LANE_DESKEW_CFG: integer := 15;
        FTS_LANE_DESKEW_EN: string  := "FALSE";
        GEARBOX_MODE    : integer := 0;
        OUTREFCLK_SEL_INV: integer := 3;
        PCS_PCIE_EN     : string  := "FALSE";
        PCS_RSVD_ATTR   : integer := 0;
        PD_TRANS_TIME_FROM_P2: integer := 60;
        PD_TRANS_TIME_NONE_P2: integer := 25;
        PD_TRANS_TIME_TO_P2: integer := 100;
        PMA_RSV         : integer := 0;
        PMA_RSV2        : integer := 8272;
        PMA_RSV3        : integer := 0;
        PMA_RSV4        : integer := 0;
        RXBUFRESET_TIME : integer := 1;
        RXBUF_ADDR_MODE : string  := "FULL";
        RXBUF_EIDLE_HI_CNT: integer := 8;
        RXBUF_EIDLE_LO_CNT: integer := 0;
        RXBUF_EN        : string  := "TRUE";
        RXBUF_RESET_ON_CB_CHANGE: string  := "TRUE";
        RXBUF_RESET_ON_COMMAALIGN: string  := "FALSE";
        RXBUF_RESET_ON_EIDLE: string  := "FALSE";
        RXBUF_RESET_ON_RATE_CHANGE: string  := "TRUE";
        RXBUF_THRESH_OVFLW: integer := 61;
        RXBUF_THRESH_OVRD: string  := "FALSE";
        RXBUF_THRESH_UNDFLW: integer := 4;
        RXCDRFREQRESET_TIME: integer := 1;
        RXCDRPHRESET_TIME: integer := 1;
      --RXCDR_CFG       : integer type with unrepresentable value!
        RXCDR_FR_RESET_ON_EIDLE: integer := 0;
        RXCDR_HOLD_DURING_EIDLE: integer := 0;
        RXCDR_LOCK_CFG  : integer := 21;
        RXCDR_PH_RESET_ON_EIDLE: integer := 0;
        RXDFELPMRESET_TIME: integer := 15;
        RXDLY_CFG       : integer := 31;
        RXDLY_LCFG      : integer := 48;
        RXDLY_TAP_CFG   : integer := 0;
        RXGEARBOX_EN    : string  := "FALSE";
        RXISCANRESET_TIME: integer := 1;
        RXLPM_HF_CFG    : integer := 240;
        RXLPM_LF_CFG    : integer := 240;
        RXOOB_CFG       : integer := 6;
        RXOUT_DIV       : integer := 2;
        RXPCSRESET_TIME : integer := 1;
        RXPHDLY_CFG     : integer := 540704;
        RXPH_CFG        : integer := 0;
        RXPH_MONITOR_SEL: integer := 0;
        RXPMARESET_TIME : integer := 3;
        RXPRBS_ERR_LOOPBACK: integer := 0;
        RXSLIDE_AUTO_WAIT: integer := 7;
        RXSLIDE_MODE    : string  := "OFF";
        RX_BIAS_CFG     : integer := 0;
        RX_BUFFER_CFG   : integer := 0;
        RX_CLK25_DIV    : integer := 7;
        RX_CLKMUX_PD    : integer := 1;
        RX_CM_SEL       : integer := 3;
        RX_CM_TRIM      : integer := 4;
        RX_DATA_WIDTH   : integer := 20;
        RX_DDI_SEL      : integer := 0;
        RX_DEBUG_CFG    : integer := 0;
        RX_DEFER_RESET_BUF_EN: string  := "TRUE";
        RX_DFE_GAIN_CFG : integer := 1576463;
        RX_DFE_H2_CFG   : integer := 480;
        RX_DFE_H3_CFG   : integer := 480;
        RX_DFE_H4_CFG   : integer := 240;
        RX_DFE_H5_CFG   : integer := 240;
        RX_DFE_KL_CFG   : integer := 1008;
        RX_DFE_KL_CFG2  : integer := 805889386;
        RX_DFE_LPM_CFG  : integer := 2308;
        RX_DFE_LPM_HOLD_DURING_EIDLE: integer := 0;
        RX_DFE_UT_CFG   : integer := 32256;
        RX_DFE_VP_CFG   : integer := 16128;
        RX_DFE_XYD_CFG  : integer := 16;
        RX_DISPERR_SEQ_MATCH: string  := "TRUE";
        RX_INT_DATAWIDTH: integer := 0;
        RX_OS_CFG       : integer := 1008;
        RX_SIG_VALID_DLY: integer := 10;
        RX_XCLK_SEL     : string  := "RXREC";
        SAS_MAX_COM     : integer := 64;
        SAS_MIN_COM     : integer := 36;
        SATA_BURST_SEQ_LEN: integer := 15;
        SATA_BURST_VAL  : integer := 4;
        SATA_CPLL_CFG   : string  := "VCO_3000MHZ";
        SATA_EIDLE_VAL  : integer := 4;
        SATA_MAX_BURST  : integer := 8;
        SATA_MAX_INIT   : integer := 21;
        SATA_MAX_WAKE   : integer := 7;
        SATA_MIN_BURST  : integer := 4;
        SATA_MIN_INIT   : integer := 12;
        SATA_MIN_WAKE   : integer := 4;
        SHOW_REALIGN_COMMA: string  := "TRUE";
        SIM_CPLLREFCLK_SEL: integer := 1;
        SIM_RECEIVER_DETECT_PASS: string  := "TRUE";
        SIM_RESET_SPEEDUP: string  := "TRUE";
        SIM_TX_EIDLE_DRIVE_LEVEL: string  := "X";
        SIM_VERSION     : string  := "4.0";
        TERM_RCAL_CFG   : integer := 16;
        TERM_RCAL_OVRD  : integer := 0;
        TRANS_TIME_RATE : integer := 14;
        TST_RSV         : integer := 0;
        TXBUF_EN        : string  := "TRUE";
        TXBUF_RESET_ON_RATE_CHANGE: string  := "FALSE";
        TXDLY_CFG       : integer := 31;
        TXDLY_LCFG      : integer := 48;
        TXDLY_TAP_CFG   : integer := 0;
        TXGEARBOX_EN    : string  := "FALSE";
        TXOUT_DIV       : integer := 2;
        TXPCSRESET_TIME : integer := 1;
        TXPHDLY_CFG     : integer := 540704;
        TXPH_CFG        : integer := 1920;
        TXPH_MONITOR_SEL: integer := 0;
        TXPMARESET_TIME : integer := 1;
        TX_CLK25_DIV    : integer := 7;
        TX_CLKMUX_PD    : integer := 1;
        TX_DATA_WIDTH   : integer := 20;
        TX_DEEMPH0      : integer := 0;
        TX_DEEMPH1      : integer := 0;
        TX_DRIVE_MODE   : string  := "DIRECT";
        TX_EIDLE_ASSERT_DELAY: integer := 6;
        TX_EIDLE_DEASSERT_DELAY: integer := 4;
        TX_INT_DATAWIDTH: integer := 0;
        TX_LOOPBACK_DRIVE_HIZ: string  := "FALSE";
        TX_MAINCURSOR_SEL: integer := 0;
        TX_MARGIN_FULL_0: integer := 78;
        TX_MARGIN_FULL_1: integer := 73;
        TX_MARGIN_FULL_2: integer := 69;
        TX_MARGIN_FULL_3: integer := 66;
        TX_MARGIN_FULL_4: integer := 64;
        TX_MARGIN_LOW_0 : integer := 70;
        TX_MARGIN_LOW_1 : integer := 68;
        TX_MARGIN_LOW_2 : integer := 66;
        TX_MARGIN_LOW_3 : integer := 64;
        TX_MARGIN_LOW_4 : integer := 64;
        TX_PREDRIVER_MODE: integer := 0;
        TX_QPI_STATUS_EN: integer := 0;
        TX_RXDETECT_CFG : integer := 6194;
        TX_RXDETECT_REF : integer := 4;
        TX_XCLK_SEL     : string  := "TXUSR";
        UCODEER_CLR     : integer := 0
    );
    port(
        CPLLFBCLKLOST   : out    vl_logic;
        CPLLLOCK        : out    vl_logic;
        CPLLREFCLKLOST  : out    vl_logic;
        DMONITOROUT     : out    vl_logic_vector(7 downto 0);
        DRPDO           : out    vl_logic_vector(15 downto 0);
        DRPRDY          : out    vl_logic;
        EYESCANDATAERROR: out    vl_logic;
        GTREFCLKMONITOR : out    vl_logic;
        GTXTXN          : out    vl_logic;
        GTXTXP          : out    vl_logic;
        PCSRSVDOUT      : out    vl_logic_vector(15 downto 0);
        PHYSTATUS       : out    vl_logic;
        RXBUFSTATUS     : out    vl_logic_vector(2 downto 0);
        RXBYTEISALIGNED : out    vl_logic;
        RXBYTEREALIGN   : out    vl_logic;
        RXCDRLOCK       : out    vl_logic;
        RXCHANBONDSEQ   : out    vl_logic;
        RXCHANISALIGNED : out    vl_logic;
        RXCHANREALIGN   : out    vl_logic;
        RXCHARISCOMMA   : out    vl_logic_vector(7 downto 0);
        RXCHARISK       : out    vl_logic_vector(7 downto 0);
        RXCHBONDO       : out    vl_logic_vector(4 downto 0);
        RXCLKCORCNT     : out    vl_logic_vector(1 downto 0);
        RXCOMINITDET    : out    vl_logic;
        RXCOMMADET      : out    vl_logic;
        RXCOMSASDET     : out    vl_logic;
        RXCOMWAKEDET    : out    vl_logic;
        RXDATA          : out    vl_logic_vector(63 downto 0);
        RXDATAVALID     : out    vl_logic;
        RXDISPERR       : out    vl_logic_vector(7 downto 0);
        RXDLYSRESETDONE : out    vl_logic;
        RXELECIDLE      : out    vl_logic;
        RXHEADER        : out    vl_logic_vector(2 downto 0);
        RXHEADERVALID   : out    vl_logic;
        RXMONITOROUT    : out    vl_logic_vector(6 downto 0);
        RXNOTINTABLE    : out    vl_logic_vector(7 downto 0);
        RXOUTCLK        : out    vl_logic;
        RXOUTCLKFABRIC  : out    vl_logic;
        RXOUTCLKPCS     : out    vl_logic;
        RXPHALIGNDONE   : out    vl_logic;
        RXPHMONITOR     : out    vl_logic_vector(4 downto 0);
        RXPHSLIPMONITOR : out    vl_logic_vector(4 downto 0);
        RXPRBSERR       : out    vl_logic;
        RXQPISENN       : out    vl_logic;
        RXQPISENP       : out    vl_logic;
        RXRATEDONE      : out    vl_logic;
        RXRESETDONE     : out    vl_logic;
        RXSTARTOFSEQ    : out    vl_logic;
        RXSTATUS        : out    vl_logic_vector(2 downto 0);
        RXVALID         : out    vl_logic;
        TSTOUT          : out    vl_logic_vector(9 downto 0);
        TXBUFSTATUS     : out    vl_logic_vector(1 downto 0);
        TXCOMFINISH     : out    vl_logic;
        TXDLYSRESETDONE : out    vl_logic;
        TXGEARBOXREADY  : out    vl_logic;
        TXOUTCLK        : out    vl_logic;
        TXOUTCLKFABRIC  : out    vl_logic;
        TXOUTCLKPCS     : out    vl_logic;
        TXPHALIGNDONE   : out    vl_logic;
        TXPHINITDONE    : out    vl_logic;
        TXQPISENN       : out    vl_logic;
        TXQPISENP       : out    vl_logic;
        TXRATEDONE      : out    vl_logic;
        TXRESETDONE     : out    vl_logic;
        CFGRESET        : in     vl_logic;
        CLKRSVD         : in     vl_logic_vector(3 downto 0);
        CPLLLOCKDETCLK  : in     vl_logic;
        CPLLLOCKEN      : in     vl_logic;
        CPLLPD          : in     vl_logic;
        CPLLREFCLKSEL   : in     vl_logic_vector(2 downto 0);
        CPLLRESET       : in     vl_logic;
        DRPADDR         : in     vl_logic_vector(8 downto 0);
        DRPCLK          : in     vl_logic;
        DRPDI           : in     vl_logic_vector(15 downto 0);
        DRPEN           : in     vl_logic;
        DRPWE           : in     vl_logic;
        EYESCANMODE     : in     vl_logic;
        EYESCANRESET    : in     vl_logic;
        EYESCANTRIGGER  : in     vl_logic;
        GTGREFCLK       : in     vl_logic;
        GTNORTHREFCLK0  : in     vl_logic;
        GTNORTHREFCLK1  : in     vl_logic;
        GTREFCLK0       : in     vl_logic;
        GTREFCLK1       : in     vl_logic;
        GTRESETSEL      : in     vl_logic;
        GTRSVD          : in     vl_logic_vector(15 downto 0);
        GTRXRESET       : in     vl_logic;
        GTSOUTHREFCLK0  : in     vl_logic;
        GTSOUTHREFCLK1  : in     vl_logic;
        GTTXRESET       : in     vl_logic;
        GTXRXN          : in     vl_logic;
        GTXRXP          : in     vl_logic;
        LOOPBACK        : in     vl_logic_vector(2 downto 0);
        PCSRSVDIN       : in     vl_logic_vector(15 downto 0);
        PCSRSVDIN2      : in     vl_logic_vector(4 downto 0);
        PMARSVDIN       : in     vl_logic_vector(4 downto 0);
        PMARSVDIN2      : in     vl_logic_vector(4 downto 0);
        QPLLCLK         : in     vl_logic;
        QPLLREFCLK      : in     vl_logic;
        RESETOVRD       : in     vl_logic;
        RX8B10BEN       : in     vl_logic;
        RXBUFRESET      : in     vl_logic;
        RXCDRFREQRESET  : in     vl_logic;
        RXCDRHOLD       : in     vl_logic;
        RXCDROVRDEN     : in     vl_logic;
        RXCDRRESET      : in     vl_logic;
        RXCDRRESETRSV   : in     vl_logic;
        RXCHBONDEN      : in     vl_logic;
        RXCHBONDI       : in     vl_logic_vector(4 downto 0);
        RXCHBONDLEVEL   : in     vl_logic_vector(2 downto 0);
        RXCHBONDMASTER  : in     vl_logic;
        RXCHBONDSLAVE   : in     vl_logic;
        RXCOMMADETEN    : in     vl_logic;
        RXDDIEN         : in     vl_logic;
        RXDFEAGCHOLD    : in     vl_logic;
        RXDFEAGCOVRDEN  : in     vl_logic;
        RXDFECM1EN      : in     vl_logic;
        RXDFELFHOLD     : in     vl_logic;
        RXDFELFOVRDEN   : in     vl_logic;
        RXDFELPMRESET   : in     vl_logic;
        RXDFETAP2HOLD   : in     vl_logic;
        RXDFETAP2OVRDEN : in     vl_logic;
        RXDFETAP3HOLD   : in     vl_logic;
        RXDFETAP3OVRDEN : in     vl_logic;
        RXDFETAP4HOLD   : in     vl_logic;
        RXDFETAP4OVRDEN : in     vl_logic;
        RXDFETAP5HOLD   : in     vl_logic;
        RXDFETAP5OVRDEN : in     vl_logic;
        RXDFEUTHOLD     : in     vl_logic;
        RXDFEUTOVRDEN   : in     vl_logic;
        RXDFEVPHOLD     : in     vl_logic;
        RXDFEVPOVRDEN   : in     vl_logic;
        RXDFEVSEN       : in     vl_logic;
        RXDFEXYDEN      : in     vl_logic;
        RXDFEXYDHOLD    : in     vl_logic;
        RXDFEXYDOVRDEN  : in     vl_logic;
        RXDLYBYPASS     : in     vl_logic;
        RXDLYEN         : in     vl_logic;
        RXDLYOVRDEN     : in     vl_logic;
        RXDLYSRESET     : in     vl_logic;
        RXELECIDLEMODE  : in     vl_logic_vector(1 downto 0);
        RXGEARBOXSLIP   : in     vl_logic;
        RXLPMEN         : in     vl_logic;
        RXLPMHFHOLD     : in     vl_logic;
        RXLPMHFOVRDEN   : in     vl_logic;
        RXLPMLFHOLD     : in     vl_logic;
        RXLPMLFKLOVRDEN : in     vl_logic;
        RXMCOMMAALIGNEN : in     vl_logic;
        RXMONITORSEL    : in     vl_logic_vector(1 downto 0);
        RXOOBRESET      : in     vl_logic;
        RXOSHOLD        : in     vl_logic;
        RXOSOVRDEN      : in     vl_logic;
        RXOUTCLKSEL     : in     vl_logic_vector(2 downto 0);
        RXPCOMMAALIGNEN : in     vl_logic;
        RXPCSRESET      : in     vl_logic;
        RXPD            : in     vl_logic_vector(1 downto 0);
        RXPHALIGN       : in     vl_logic;
        RXPHALIGNEN     : in     vl_logic;
        RXPHDLYPD       : in     vl_logic;
        RXPHDLYRESET    : in     vl_logic;
        RXPHOVRDEN      : in     vl_logic;
        RXPMARESET      : in     vl_logic;
        RXPOLARITY      : in     vl_logic;
        RXPRBSCNTRESET  : in     vl_logic;
        RXPRBSSEL       : in     vl_logic_vector(2 downto 0);
        RXQPIEN         : in     vl_logic;
        RXRATE          : in     vl_logic_vector(2 downto 0);
        RXSLIDE         : in     vl_logic;
        RXSYSCLKSEL     : in     vl_logic_vector(1 downto 0);
        RXUSERRDY       : in     vl_logic;
        RXUSRCLK        : in     vl_logic;
        RXUSRCLK2       : in     vl_logic;
        SETERRSTATUS    : in     vl_logic;
        TSTIN           : in     vl_logic_vector(19 downto 0);
        TX8B10BBYPASS   : in     vl_logic_vector(7 downto 0);
        TX8B10BEN       : in     vl_logic;
        TXBUFDIFFCTRL   : in     vl_logic_vector(2 downto 0);
        TXCHARDISPMODE  : in     vl_logic_vector(7 downto 0);
        TXCHARDISPVAL   : in     vl_logic_vector(7 downto 0);
        TXCHARISK       : in     vl_logic_vector(7 downto 0);
        TXCOMINIT       : in     vl_logic;
        TXCOMSAS        : in     vl_logic;
        TXCOMWAKE       : in     vl_logic;
        TXDATA          : in     vl_logic_vector(63 downto 0);
        TXDEEMPH        : in     vl_logic;
        TXDETECTRX      : in     vl_logic;
        TXDIFFCTRL      : in     vl_logic_vector(3 downto 0);
        TXDIFFPD        : in     vl_logic;
        TXDLYBYPASS     : in     vl_logic;
        TXDLYEN         : in     vl_logic;
        TXDLYHOLD       : in     vl_logic;
        TXDLYOVRDEN     : in     vl_logic;
        TXDLYSRESET     : in     vl_logic;
        TXDLYUPDOWN     : in     vl_logic;
        TXELECIDLE      : in     vl_logic;
        TXHEADER        : in     vl_logic_vector(2 downto 0);
        TXINHIBIT       : in     vl_logic;
        TXMAINCURSOR    : in     vl_logic_vector(6 downto 0);
        TXMARGIN        : in     vl_logic_vector(2 downto 0);
        TXOUTCLKSEL     : in     vl_logic_vector(2 downto 0);
        TXPCSRESET      : in     vl_logic;
        TXPD            : in     vl_logic_vector(1 downto 0);
        TXPDELECIDLEMODE: in     vl_logic;
        TXPHALIGN       : in     vl_logic;
        TXPHALIGNEN     : in     vl_logic;
        TXPHDLYPD       : in     vl_logic;
        TXPHDLYRESET    : in     vl_logic;
        TXPHDLYTSTCLK   : in     vl_logic;
        TXPHINIT        : in     vl_logic;
        TXPHOVRDEN      : in     vl_logic;
        TXPISOPD        : in     vl_logic;
        TXPMARESET      : in     vl_logic;
        TXPOLARITY      : in     vl_logic;
        TXPOSTCURSOR    : in     vl_logic_vector(4 downto 0);
        TXPOSTCURSORINV : in     vl_logic;
        TXPRBSFORCEERR  : in     vl_logic;
        TXPRBSSEL       : in     vl_logic_vector(2 downto 0);
        TXPRECURSOR     : in     vl_logic_vector(4 downto 0);
        TXPRECURSORINV  : in     vl_logic;
        TXQPIBIASEN     : in     vl_logic;
        TXQPISTRONGPDOWN: in     vl_logic;
        TXQPIWEAKPUP    : in     vl_logic;
        TXRATE          : in     vl_logic_vector(2 downto 0);
        TXSEQUENCE      : in     vl_logic_vector(6 downto 0);
        TXSTARTSEQ      : in     vl_logic;
        TXSWING         : in     vl_logic;
        TXSYSCLKSEL     : in     vl_logic_vector(1 downto 0);
        TXUSERRDY       : in     vl_logic;
        TXUSRCLK        : in     vl_logic;
        TXUSRCLK2       : in     vl_logic
    );
end GTXE2_CHANNEL;
