`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Yj5aFJvvK+EkYaxuxgQa1myrU7t7TtmNF56EUP149TVbOaR/A5CodHQtqRtgHiYt
/30z/f5SC4S6vUnrxhaC42HtNAG2iEfyGlKEfUHblDjXGUd824VwmzBqgvgDWXfx
/VQAILhrY/j17zzexlVHWqiA+q6NBCsRjUcamzok8H2frlJysb7R57ojZv+s0Ng0
n6Pdb2689OWtoTrDfoyskavJRySZgHKdfU2jHfH9D4PklPfF6BZTHXQ4ik/90O38
gpf2xAupO6BfnKy790pZCZi1Q8JBCHJNaqpiKqED0cg=
`protect END_PROTECTED
