`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SZE+HvWaHDwBrbYo9zrK5KPlcy2yM0aJKkTnQ5hcIBPv
ynPg9V6iBkT9rDwAKXeETNhHdvBF/o+xT1PMKNh1kUi2g0SsfwEjSGwDWRJLyZJH
YTdTgspgNbFKZ/zqheYlzxmxpzRbxcGYDROe/1YfWE018IM4MmeYisQiUPDA8FNy
9tM41Le3FQH52dwdh6hltbl0cWgoqS8DIIUiD92hAG0UTrEyWPJnVfk8484njehR
+Ix0S7Kc11WSNW3tz2IWICzgdxSQX0cpSnPHPFSfnXDp3jy1qST3/MPCNkUVGDZz
`protect END_PROTECTED
