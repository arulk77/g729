`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aZ+uaZkk3vy6GPgx/crMPse2odnChRdQVnbLkNaDHDgE
f8DyMiPqckBPyOaDhGEH4Ji2mckEngAi07Hf2cH1SoW5DBd4739indZXy4bTWyCD
G4zgxj3pugxDtxaudnvnE52Utb2jitEje6E+ek6W0rbzrIqrDVo8QoKLkZ0Q1K45
tOr0NECxxtGQyuEHRvcp/D95j1qZUcTyBWDl7k8Lgb8aGH0OHU9EAP/n9ibjk1Du
xhvPPjHUwA63RqWvM+7TOc2dOZcg9j4/3gWGsT9sgGTPa5Ykg/ANn0w7T6b0XcEH
YbzHsUJpHRvkP6zU614wygOXqXBC7/r41mc4bsbei5krNrOuIJQ0/fV/f0Wq3ZEr
67dgAfqDZN5CYmjPgRYKg/9PKFi5ftNgzFSVdvo9LucSYez/W94nV/pgOtAGe7mN
zN4ulWD9N/4v5UQo2cC8gZnB6iLEo1YOgNAT4xjbmT0=
`protect END_PROTECTED
