`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47X6Ju9rmgHDiCcS43+1+eetXMTn0HqMlW3j2wtkDINE
XwpNwYf+N3DRKw67i4ebkq6t6uUaNAUYKxefQTX2JCxHkqmmrwfplD+SA9Nnf74M
eMnKLy9+5GgHywwNSzfO2gwfI8xNKyZop4Dc6Ii2TjjZ6184rAGxXs1GLWLXUxoF
a3hVR8LEqNyun3H280vphHP8rwF9ZkkKyo4lvm/5SGw+BcYUJrslQSMdjHaWHyad
WfPZnZS4GRNgxusnVJCECXWgw/dps2SaV2PKVs5Y/IFar/Rr5jBJ6I2+yceawt6x
5p2P7DhbRFtq7KE+UPu3QQ==
`protect END_PROTECTED
