`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN64MuT20qtqdqyGDOfvznemEXWsAEgHs19yZ9pVXZ0lE
pVuoCZUshALcmKlEq8NS+2xGRvhUG/iFTdprarysk8jk7MzOv1fx7AP57oSetbqy
XWgZbM3mav/s//dxFKsTLi8NRnRPbuqY1XNKjkHBx6IjXTfqAOx8ghMjQ9X7l0YB
va4B+y8K53Zce0qa9BlXmCJpjvWsKKWmEOvFJsj1KX0QSCpyvunJZXvisCyR7Y7O
Ye9iMIqDbvkqtychvjd2cIfU+maIUhE/MflxFSWHvnIC9gFrXFczN+/Cw9VHrjs+
YiqpARheXIMVkIt4Xv1DmAVS/uW6RzrQ5IIcRWpvbij0fo8790jVNgzroqG6kMCL
2tlBE95vF8JWGJVTJ9RLmdXADhTaoxY6V0eUNH67iq7DsnUXTuwiENbkM1fowU1f
ls59S8VkHZdqOl0K8qt0aVhgRCqUD3MRvqDxbqesqwM=
`protect END_PROTECTED
