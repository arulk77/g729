`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePLz/iVCJi8aH0EVYwL5gTYnyI1Pb2TMh/J6PGvoAoTY
wAvxkadzdKeWIUXJrU+r3f1aNhzg1snV3EzdFADFaaghdS6CCr6Ni7Y+/Bcsh/Yu
fcJuPlRnl2pUgJ0R97WQRZOpIOoxOOF4R1ZwUIs+Jr12Gtdx6gHSm0yanbN0Y/CO
d6eqeybsSP5V917rIjUjqDQYz634xn2bvJ6mue4xOZi+Ool0RnNvjKYyFOzON+tF
shHs9GzdOhPO/0AGNx4qQtMRGdGPSqY1jICEB3VSjmPIzOjjVXD94KnN7q8c1v+5
/IFeIlGVCqzl/H/OLfCqhQgCi3ZHI2MzhkW4Yi8bwEgrRlirKGT6bmlescQNxNFu
7/WyQ55Z/V+FUg5rpMINn9csTvph30BD2Nc9Ed1TGQ4RV1Eux6zipBe3u2VlLIXt
kNkNl+4l+7eZ2omTCZ0uc9xly54NoZsrM7h6Usr2w8DizZgMtSmZQelHv81ekHLG
`protect END_PROTECTED
