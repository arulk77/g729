`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKxg7ZM0r+yz1vni66SirGsLufYeA609r9Upg00yHWrG
BR3QBsyC00Q9mK/+vYcQaWyLVx3GGTJJo4Ggyf5SZiacibI3WVY7pP5rCmno6PP5
hkZsWFOp5A1jbHfF6gTdgGlypb59hPABDEc7cl3I9G5y3XCKNW84VV8Kfsl3Y9UV
SZmTmPzbpY889PaERNhqxXSZSBoF2k2NQF+SgsDSnvZy8aeeshzLkmGLPDWxpQJ2
`protect END_PROTECTED
