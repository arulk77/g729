`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFINtRXFcqudY1iDOypuysFw+DBVkTpeBwVY/oaDrJ39
l/EnrxfkGHklFL9eXk6hfXpImcNTRk2hWCTJvW6MAjWEHzFQuQN6besdPc341AvA
BafSMDc7w1PxZC7UIoyptFkbu98ZJcXNEeBnpaiQIDpVrz6k9fXj1vW7qGxXy6lE
8PkqyFeA4k6DYHOFesRRJZE+YjmWkMoxRl6tFh71tTLr4h3MEAXjNs4MmDbj5MG/
KXvqP7/UNEPp9R3mPUC52w==
`protect END_PROTECTED
