`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/ePrT57aLeFn/qVQdIi6OtgQMIJn4ysLB1ChkWdHZ8h
0ei+SOukVnVyceUZa1NoZz+aLHuUL9Y/DprxycgrTis0weeMNK0HDt9C36Bg7SY1
Ss888emwukHPDUZfxW5q9b//FrFIHcpjtFiqOPI1vVtXA/Y0nAVoONQjg8hhzkDK
ek8DJxpsLXUTrxcNsMwz9TvqxIo62f0sQILVkd7Eqek=
`protect END_PROTECTED
