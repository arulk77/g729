`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveO5+nmZbU8t5Vv5MExiiFh2gGozJPFxWjkwJOr0RWEio
hrLvSQpO55XFtTjusnk4WqEO9JHUv3A2EkbJ8NdGA3A6v/w02YwuqrxIUdfQZXxw
MBUdB4tU61s/QzAqqE+PZ2f32RApMzDsF9Zqbxo2ileibOdF1rBTxdqRwEOmyx5+
EeXc5ejUhBCZt0IbxBOIhD3c+zV62YnDolvB7d6KQ5DJtf/5Zd/jcS5W+4uq/R8r
SFCrNDlI3XwGK2UkiJmNFekeab+juIXq9w6C2VT0D6HGLTOLt1QFJ8w4OZsktdT5
tDcVih7vK2Oi3G/qMIWsb1iTVz6y/PMrFVFp6iwzTATJZE0U4OeKcxCqmo0L8Ur9
+lBaJz1TQprrb22zwwVRzQ0UUPFQ9B2YrKY/dMzyMJ93eKUWgYDn1wR1lz7Ozhx/
NFyqGkzBUQDxp/CkKFB6vKotvJnu4VNXpS+5FwSi0JvTSKHT/gJWbC28SlMnduxT
zeSvLWvyEYucBE91jtpy/hbUXAirXjKsu7Mgm7Q9yh25+4HGQh+tmtw07HA06B3m
aE+VI17s/6sPoWUnBaRigw==
`protect END_PROTECTED
