`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
/QuNq/E6h6cJFj9EIRvn9HFo4u6LjTIfZ0MLueMHlBec0SHrb2s+lIEOR44B4Rcx
WDPq0U1q0Hwc5srIo7hTU7DfN9bBY76wcbXmtvgKpeq+5HmuCVjxB1xs3sEfR81u
`protect END_PROTECTED
