`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePOpzXQj1Ht5ljHbXcXk7IX5I3fU3hPmE99QTYBbaSXF
24hEJy4aeKF3bvTW9jD2vkl2U1FlfBRTv72gkAj5YsLONR1d6smA+0qX9646Sp1E
c2fKXjtdmLcrjSUIuuGanoSMADxL/2Q8TjoHxBMMOeklqPOpp1t/+hn6RtXOw5vD
DJix71C43elZR5I8KqFhI3GmtKmdAzXkE7d5Iw5jQ6StdnEx47cOwSHWOWPC7B88
kzrmumq2zAdVRCDr/Jgn1H/dRAkrXhnXdofDtQrlBQlyVHsyzWFQCsAMdpPNI1Hv
OUV3nzseVFFhiIESRTyGy2+V7anSlvMiUcBEv7G2CVcy4W4f8qGP/FBCr5EEXtre
2f15UYjjJl5ksIM4hiepbVEPDZFjS1uBtmZBMngzP6hEfpsBGVDsO55vrrEMfLZ9
EGEoH3X0QgW0r2+j3Srbyb+WGBGwzquf/LdHcXsr0T/SLMAI16d/kRLV4jlUlP0O
s+a5561xqNIWZjf2Ovy2Jw==
`protect END_PROTECTED
