`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ab3t38y2wf5+qsH/48ktMGFFVEPPKJd2VkzBMqM4dXjttvCBW7l/5IP+Ry9HTBjg
xs+hUt2jkvMGzThE5LThE42ZxyVzQF0dcMblsh19QABhuk34RwvCVsiHcby61MYn
xvvRSedbB3+s3IBpa2yJZjI2ca8LNp6spyQeY3RGL9H+ySQz/SmCPoSNq3gfcySD
NpX1FKVt70SPkHlnkukX3nbIaCJLED9o5tGBudrgu489H55a11TbeZGPLioIvIsm
z2/QeiqUrUP3CzSEutwX+96X/9IS1YYIeT4lZCus2f21zVH20C423LPH8I915hH9
rLmFyM0hfwzA3I6KuMCr/H0O7DqrYhfYOClpdbnOsonn1SGMg6lmVtoPHaaH4Zcz
CC70Km8zjL7lu/Q0bIG3Ns1kI8cea6XYWQCt7HsrrIk=
`protect END_PROTECTED
