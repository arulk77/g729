`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
dtIYeFtD3wfdsXiHha27Y17SyIqwLMTzxYyGzzuEt45qK3j7WFB9bGWlgxj7/nvz
o2qKPav30L8B2x+Tu5gBExLawLQWBmSxj0YeteGABy3PdfOFmSjg11xekM7ImvsG
IDcHEdKAQ2BUZaxzrKYjLUvNqWwD3v8g2zh6GDqqpupB6JcQJqdOERWPgpk6g10M
2U23OcrnsyG0ETdlMuz9tHbw0aizQ6gj98VWGSp5b46ADXU8iqns5QI97mdtJ6SH
5zYCY//76KZ2CheHhfFkpcOVaGttAoI+YaiQVXG9NojVTCOA+QrJb95dGwRDDI0K
OmgwkvBfyeLRf+mJPULE1fcd/P/99zpfGeIVYe9V8TJHcguRfDr//h5uNGLePSLV
fVnCV0NwHmp6asgURaJPqpDtGttIjthmoOF2FHcSnNs=
`protect END_PROTECTED
