`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43Kyc1KMKvf6N1KzPO0h186I4kCyxuOccyAjS8Pdzb64
jyyqvscRQQ2T3wCKPrAQL4RABojQ5CVhzoxAbIHOc6D6cnSs8SrqJ93y4RM3qQS0
lkaVzjwHYJh+q+9Jv358yVb11SrX+el1VDY8VhS9oP4vV0yGh7oPhc8Ea7MLdS40
e1cBTSDT1/zAmRCyupvkO6WwBl62Vk/a7Pl07g99nNbEf0bZoOlE0kd/ntggY1Wq
31kb8DVrpg9BMz+DqRDxrCvSXo+Kw1CFWHO02HEub3yAIj+oYtaPxzARdPBXwLib
BjYYnlp9OrepdPL+iJ7Kesq+dYhJAvHRWll2hbsh+yH/VwnsDU9joTs5p6JPueVL
xwI/jzn4ALi44VtWKSY8qGbM7K05K1OSku8Q57tWogWr2EW2E0cEKzQO5SMc2ITR
1B0iCv5xjI41tdacXfNuFDCqZGyEVodD02GkJich1F+b4XIx5T1W57Gih0AQLIfa
pQ8OQ0nV2iaj3C3dXJuju483YTwj1qyOXS7Vpa2UXAULmvcB9P6umDZ3lm9A4AKt
I/9uRNtQ1xuTpM4t/qhIrTAMxrW4FCY1MQQkfVUwbi/FP6ha52mYVi6TIFzu+UY6
uFOvc6POTJQpu72+mTF8EmaLvThXusIXQ470nm9X7YEYQ3wC1AafZ+Nbu0x3pJyc
aw8WozSIkVUHdt3y9Jd1HFTPN03VRiibiWP8dSRpLmqze2j79wy7L0TczQotE1an
b8/U5ifofkRwH9wXJq3SNg==
`protect END_PROTECTED
