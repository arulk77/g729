`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aQ6hPD2pMA6cuNpv+tQbsgA7/wW/Sqp+I7SZqv/JAbvE
N4pxCQlYum5fVJiMWjsOYQMLQhOphp4/WThB28aQzfVEOQHgkC2ArVAW2NMO3b45
etlaumu5TAbz6RhgLq72k+MGJqxw1rZcLZnJWsx0kRq2s6bmyRGbY7VAc1VgC/nW
c0j++8HMGIiD+V5NclPiU4ocOkqLRC164CD/SjFAgXfgHptcu6n8DbOpO1jrF82N
NAy+HVBpe2+jP7UiJ/ciDvtsQIei01uSOoCSEFdfS9A0LlSPuUloJL9u+/uVZ3p9
ZnM81rJevlXqGqhQ2D1mIoxBROZUtiOVlnF/t1aycmIgPSnw298lKqllNvXdL54I
CBcZapFT414a3e/xBgZNCNTJ6oylRR6521Hf9ZCzXWOpk6jYjpQkz6sYcsJoL23G
2IeflAB+nJ9/83EyT+WU+oQvX0UY0ItPz/+AlsIZywAgEaoxrogxC1xexm9fYoSJ
T2JS7xGkFQrRagRlyzukPCL4lItx80FWPeXDLpK55wmteYPPbSLaIoTTuzdf9qlJ
8qORpcFhZJ1ztV0cxuztSRV97fMjskyJSKOPEx13IMbQo8VY0KdD7DuG1+kQq95T
a2KbSA5a5I97Sw8g5liC/zFMXrnlLBWy0GtxK9DSs1FjJDGmi7+AeUwjEswYCmd3
JHIxzQ6/QTdxd1xfwpH/3bkDbF5qHJU51TLsQDSI5QngU4nCsWhJOhkPTCgM1umq
pq2odKwq46cYHi53xjFJwewfUN0P/k5AcOgcr8uEILWGxBXXisj3MtS/RJXR1omF
DcuKbbdLrV7duVhgbihw0m/dzqRP1c37aMntXVflIBNLd6Gpf7LzqqsmJF2+Krnm
4K2n51uRcwQOldl/47pLFEUT92XkY2h2sMP9T4n6zsIkzkT5UYJJrkI5IgFMhfSN
/LbcYEH5iR1u6Sf7qVeAQjGQtVnacuw/yZVcFxgA+8Z1Cw9bGAs1RoHXJ4p/e5Id
GAwk56Aj02yRjFfa70TD9XY6dnlKd4+d2isYohT37JtctNMQylNeWG8KByuJPpli
sKv5gL7OaS+sSTWJ/Zr4fcGrxbwyY8yMjpRDLU52GdZXBIYOlBYOBOibP+exZDfk
MhevtKdK/l/MFnC3UH2npbJ/g7V2BZK24DBo88J+09l+POpYLbV21bRxHWQBHv+k
KpIbnd5zInO4NUELwO1+tWeBqGo2XwiWWbz+XekXcsj/T2zFuEbfUcZkrfQXRc1N
II3eMUFzafLA2feZ467RlTbALuUAsDdmefVbo98bn37vqHSyn23CX20Jo8WPDLYU
rOJP2tqX1Pjt+Or7VuIRlMujxfAOVZGfUNkXgec+1cx0kfFFJXEtzzH1HV51bHzJ
PFCvYxgr3wHwFy3mWMq+Gadzi/heBUBKiZrKu1rtUVju7Dx7VD49q4DG4n11C3JV
GbM+yx7xOq2Gg53zrLtSN+tBp0Hbj8l46DISxsktr2e4l+fEml4nhtM9hlmcggob
Ou0rUYQw39WhnhWFIgUcW1rCR8s6nSC5fnqBTGOHchU34iJmIBQuEUC8KY/Pk7cB
ew2pX2F4b1KvwyYiNqhV3uYC7Eu8hJ31POR8Sg52TPUhPW1W2ptCJgfPOdOpVwa+
X6Wp8KUyAaxEwJGe9sbN2Jr4Zxj33rS0e4pH+iV23gyCuZbsxDYSFlKsnjeXFG4A
t4fVwfmSRYsV5S281hUMZa9y3pxUrp0scBnj45ICRRiEJ/NCRWeAwVtHR6h1HNIM
5fVelRhe36IhUpze7yc1642b+G5alqpM4FgufIahp1kcrlVGwsV2GBKAIt4Vkjoc
KNnXE0JoooFLDegPR02oZuusLTrGjo7pAttGUQLiebzXz67pMm69cj0wK2YC52zd
UFViL7wjvgLbP0FwBt+hc49Fzbie11xnerPsy/qGl7GpZmL9hScsnIpM9LQ8U/Gr
vubjS9D99F2nrf8S5HdmhdW8mzuyMosXqapbNwttwqWmjH0TAyZIn09VxDGPYdji
mj0pNzjMoQoyNQbWXtIqfyokRUzD05h/u7mmC2oBG5K3u7koF67hmf3u1kce3xDb
Eme1AgXCj4JKTydnpObRcGXpACgB8gGFjbEy7pfy8E8WBXEMoM8cVWk35RKxJIbG
1ZG9f3Hg0O3OmgEcX0huciNjWip60kTnyQ8/l3YIPU4gJUFZS0Kzoca53uAOvr04
1jjQubYWbzmvSNPwsrZ4uFMOiz7AK6uXadjMGVFYhqAkNXFTO4j7hUOv66OC2HWQ
7RnX5mhjTp8DOPgUN2jRKS99ErCKBRWsT5nJEzlKWf4VKjKwa34v74NaRshBFqTa
3m5DeKY6AgPHDDTZnDVDUEiQwmHU2rZ0dIjvRdSeH/UXq2o0x4qoYO4M59vchwB5
IHMcVTJvqDGRfpck7gIFUXyReVYdxkk7umQDcb9OfE8IlgmSl8b9TOXpiAaLUjwe
TOeLzANETjdvEeAHPAJAS9kNgTY6hrhCQW23PokYoq28GQbfUQ96zDemX01A8RFI
PcZP8T2EknRp3iSBAZgO/4Um/+emq6Lkq+BBgyXJN4MokeRVm2d9YVrFSjMOki0U
yC5u2dMyGNdYXNVZAId2g9yAHuHhpZZMy7pG6YTfwCvJFFEW1YRGu4lzTNPkB3DY
b4pGXWaL8ol17zOJ8Kucn/uWT27VSYRxjCNBKfypp0/qMzfG5QabRy2CKDR00OUr
QxoiWabo9OYx01LwANvDDy4sGVFItboL+OVpSHEeC6TcPQ2b8+5G7x4PDYxfSG+U
c5OFLgXK3ZHaED3NmP7/W8nq5+RWu3EvMIBWtdy3db/Hc7jnfiC4cg5DidbasPUb
CGbqhh5OUYKTkLpcvgkgRI0XDCRL/MQVhM1WtlgBMB2ZvJ/RTV4EodT4fHmZjREH
Md7+Uqoh3UdmpxwLrwB49EuWXx4XaBil6u3FP0u9c7HVoWDzcb2hiz1MKFcufy0q
hNJ29nWnUE+jJnJbJzh4lsLc+9sgdfB+ssCX+zOtfFBDttnIyGvJTfUOK19cYxb/
UINDJi2i6+p4frhx1sEC/Y7dFE2tryp6afkBpk9dUxGAVS6bx0iPyXxQGdsbMKtv
aKNF0XcB84wW34rdUNNg4T90iGm0zQe/Q3GgyLkRUTNPuQuiQyntdyEaP+M0Ed6e
ErNOm5uFaYtIFMrTE8QQ/VGBfsGNb6ucXxYDlU0kv59NKxStAn9DKFmd3BJoPhN/
1vZLEg+0aGqY8sTIE1/stJM2rmkPXrPrVWg58l6cRkC0wIhM9k03BEncav+FYXM9
a/fZGtxucG8iaSs+lMxMMKTf9tlx73jifWbeH/EjzlT9YX0oV9qzDcxaRUIIVtKn
GO6i4pqfOPUCm/x+XejiqrO6vSEkBblxKm7FNac1NkdvSafYfWXdVEADT0MOcukF
fX9S68IlqvI6jWR3ivPnHOA21h0hqI0q6Ax3F5NW3LepiftsnQuwWufOLHM6X0Vj
ZOHc2QFaOHR4Xu2C9g3mu313Axn/vd4MrB+lh/yg4pu51aQ2h35TFD37W1UAKZt6
C736ZCDd9nkncK28nSHuE7GVYohRsTExPl94St2dXBTay8h2TG3fIvMbBgqfxB9z
AjbyewPWZnpApvHHSLNx5cRAWW9XHxv/y5OrBSkWyi2N0xWFejYYPlK7pzkKaMat
BXAppcV5trOwHTJXCl6QzLH6waVWcK5D6GjsCcCHRC46DdmgmK4Rci3qf8SXhrSd
DNIW7sdYiI6GjMZsnKs4+fS/dsBnwrplzDE02mczHFOhF2xMfToIfpoB4R1X3g7C
GcpY3w/hJXalQPPwCnrd9t0xPfVTmbgp/mgrsD8l0brpbFOH47/NycyT+ce2qxGK
E6NUPFc08SsRqk+f8AIdzWEFGgh+9izTXcNxh5l+Z8eFQMfNeEGUtW7RmWDBcdb+
nS9ArJonuWnTlIFiq0sHxpTJ4NH4iB1JDuEQB7LLPpimuid/9YVKv+LElZolGTZW
FOEynflkWkp5SLM+fBjaQBqLO+qi0AabqYn3RU1chwbp+MLDJzgZO5uDdHy0Weh3
McTJTPn8i5z+pFoyoVJ0ntIppA3YfWQdeoTvPS/Z4xk8TXit670reDdXmMZ9rACt
haHgS45vqhWB3+FY9kL4Ma+VUtq9xm07XSOr/+rOS/W0NWLZRUiYPrLD2mlRGVmL
nAu06vPtRBynVe/9U0gf5km/czDqPYPsFVcT96PwaoEAok26HzH4Q7E4vCbEW/7A
KsShSoS/8Y1jV8rsJB+VFgd1UjRJcqVzBF2EywNYf3di6AGUh8AAVtK65W0iXlqB
7711jJEEjS4oFQSOZw56Il1sb3quFm2IfE7/0vYFlyYt1poDMN1yPyIYuhvxiymU
U0XkkC2TjgsSz2EIrVi9OnSvyUxbfQQQ/z+2J6zIYUzPLDRRwjCD35Qs8WIFBXSy
FnhFt2GbCQ40tCcvNJKD65MJWGcJVFnmsOoeKJkC6KhjT54Hq/uz7kQFZniet68N
BuQB3M7KvofglG4IdErgrZMtr23yND0BLmf9JtOkWGchaJepP15dIjyWAbqBgCR1
Xon0gVYCkjWpcjNF7WUwwZjl+bemlQdu0qhD2V3CygXnGPNoRt2U+y51cw2QBs/w
wLI6bqqCB3CYTaef7qbw2AHNmD1G/XIH6rCW++tjrfRQeqd8zxPWyJ1fCp1tZr37
azCqoZHes1IGWuCyrSs4uO2FOlp7WyBxxTdNwwoMWxYTlrQIx2T2mt3n/JxuIRbe
5lc9TjVdLGSi/sNNEOx5fi4SJTb0dDmMxT2Vk3Wqhu6y07oX1ZRSIHhGOTfIztt3
P9dY+4VWtcq8UPLY9wX2Y+55kGlWBt46I/TC+qhu2/KzUiehGaIwF07cBrg1ZHSj
umerJ2UMs2lEXM9GYgTlWjGbX8iHAngjXMo+8dBLcZ24UB8zdbr9tLcJAoIKsYi9
Kl7D51ov70rY0a71LfqBUvlkvqQGXO+2YcxyndXHA0lsEsJF8EW5II2Rnyk1zM0l
l7md2qfABA1AgMtRbfdkmL6BVIQOIF1UokvOAq4zCbk4BIc8Gz2VnL86hv3JwbvY
zWbOMN92DmUL7ZV0L6OTueRiiECqzlCubk5Ws4WYAbUfkqykW4FAncmBAqjhNDSr
EJLL8Pdiu7mYG58fBrkpETsv39R/hvpq3nac0d3PkPMhMg3Ye9Q5HGIPa+DIwZe+
Zlw0O+LEGtaCLCZ2k2mkMZ8/qLJPcTP4TqOmgiaG29OeYWQRSO2e30VaHLWSzpE+
P7aII2ocIpx8vFAEKyRJKCzb0bU3QIISaFDk1NyePFFrnCKLI/td8Z0kGVZ//K+r
cKuItNtGjU7+0mqen8K6OmttxocAW7/t1naDtyIxQ5mk6xgr/b3A8MZF0h43OVHQ
dva7YPy7PWr7Si2l5RVhUM6qo1JIG9nTufmeHhoBKh4PVKO8vzNpVcZmBIzIDNWg
VTpwqGdq/aakOJ1Yh8lX+wOus6DKNlQ0b9l5b1oN3BW0CtJAVI4JTBaUERYvteVi
mrafm7LLDBDAKD0Kx8q72BqWbo4jb36ViXJaN9U3tCXjANLiAIhRLw6mNt/G+heh
6RwjLqATCm9FyoI+Eh2B5+3B/YE1SDIqMfNr1BzkdQ7HEFbhjqrfavpLJ6fw3EFd
eCZFFXGJ+yfqwqyOGXQeHeB+Ecb7oCL5B/k9Ysd10m60h5aNDPoij4Or+FqXUcxm
jVK5f8YjVq6zoL6a3+KNwmAT2h1MtWQIvOqr4epslA3SbPCDzJW4emFR+6VDMz0a
2ita/XmbCbTAqXGF1R0gAhOunNB4lXnHiyGkk5bfFF4fB1MXUcZr9jw9zg0KMm11
vDJjEnroyXw0G+ytmtqPDKILzfKNx6wOdhfEoMKjWvW9MTXt7XIBMJqJCcazSoWy
niHBmzquV35Y4W0S79nbmqXCy6L+gxDLIxxL5hLMmYTQmq8IN/xaDbMa4i4qnaTv
PLg002qvH6zGWrw2GJrhAjT7oQrj7y0c64Zc4tF7bC3KXaAQj3+XlvXZrWouNYza
mn7MU63Q0ioFRwMG7WfFJ/VdyfxB/RWeP68cOk6QDsL9t9u7uvVWocOKtwWgEwbY
un9v18sAV70yhEDVb2Vzg9UAoG6iRcXofu48egAOAVPN5+UbMhTuxEnbexNZxc4V
2hTr1OOt7qUeYhtcVoCyZj+foC5ghSngPl0kHEa3arQCMvFMmC/wtOYdg9Xm3efa
hk28IukXu6UHLPuUzhfCXf3PCTs+jxQYVT83/nm5h+RKWGag7S5g6hEwdybYq1Vv
e+qbVY6RtecZEo1dPZZQbQQMh0vKCY3tUAbaBT05cmdM9a+2tjO0TMu+rHocN6Dt
+BAHsh3MNeVjKCKZ/GKHsqfWGMMEh5je5c/X4eyVzEPTkB6ZgwY416UDhckwx2rC
L9VLmwRg8DfWcquikPEGRxFcc7ABpdyV8rVtwP0lVO9oX64Kd0xeo5LW1NWwQEzq
f6dH9oidchIho1a++uy+LUmiBsY8DhNejSweKeC1RBcP0u7EO/euzuHEqByK5bFF
XuBf9g+AwhZZrr1K/WkSXzKBmdPc3qwgmjkg9knf5LcrQ1I60/uSLhtXgbfGNngF
aLGDM9hX5cL8OhNmz9WoxltHQnoy6e0scVJmkBN4EDekjsa/n29Lu54dX7+aNEns
93nj5JxOCfx+S4UEMLiuJnYVD5ykF1f/31thRCEbVnywKpFEPmFyuOJzvXiPTYC1
JQUsnQ7Bd0q270YgCU5Oigjib6+4uNjZnnayGKUVh/4HlsDknoJZEwZtDLa5YI/q
NGI/Y68EPJ15BpJtplFptAkUwXTk9bnXZh/VkHq9v6CLHOGue41GobZlaHF/4iEu
UcTXG5DafvLtBPqeL991ZaNlm+3ox6iZcOMn+Zp16u/bsG//NS0ML3rfV1oqxgio
mYessdPbnvX8sqW3qe1kv26yPGL3eE9jBkAeJi0Vy5hQrFP6MDaaxKl7Jur/k7Lp
+LUnB93CmYQaBGx6R1PzLyWRBT23IXGZthxfssgd7MBJd1uI1k3RUykC18h48g00
+STUewuonpgWdSBd1i2hxxfaYwnTcZG6WgNbEYzlf2kEj3Pyqbjz8hdCPDe73DMk
8PKScxT7k4t3b09HYa8/tT7its1QLn0fjGIiSDALRBADq92QJfozu2ngMW7Cdtwu
pULvbPqn82mUTHfrv4PRc10JRuoKli8i4ya77RwsVjsqBWhl45BJiBE2si+dErLM
tVgJeQQeXG7721GN6413B7LY4BdwX+ub6oAhOPhyrot6tutfm5HPkCXta6KMCJ5/
IPb+bt60KXb8RtgBZBaB+hpptuy/gj4Y7jkYE8jO1ojhSyGvNO0SUrrLnodllYzE
ZpXgSnGqbHiGAgDsrUY01/5+9zrykxYPcra8DChGkboqTwrsYiC4K/RpZPAzrS/W
TVrX5fCcrzAKG4j2ceKNzWW/aM8kIcVx6aVNvORMpbUNkGZ3wC9OqViyynRw/eGc
U1oo3IWHKbSQlCTEtlqMQra8kq4SJC+QgAQhAVLoIUvFpfCRPhZFfvvTQup7tgE2
rryk8sHC/1l+Q7wHkPZBFel8TUHit7/HTz+gJJA1YwzJIs0NRUplGZWlvYchTBY3
Emh/vMEHTl6g0cJoilyRxmny3n2xTiLFlWjtB4jwV6zITkFmNHiUjVDxGER9MfM7
/i5XhzsYBD46sVizfk09lysPmJKt7xH65tue6rMvzCvAHrEaTWBVoNlGKl7YMDYX
/KFt+TMLZWPSl2WxvadGbREqD6L9ZR47m8IWQE8FWeS/Bzfum9A510njBIP1aKr/
t9pLZZbAbVX2G255jGSmaaVcC4L/e1Y3h73tBmyW9GbJZFVbXlTp1JbPPa3iUV4v
HKAr/J4mfrwYweEdVKb8lh+2Dq7lqu6+SOnEaC3j04Yg4nX0aJNuZZck4KuatoMZ
DQ83+pmr2iyzEyrquCQaMZ80gde0DEKAJDKscdWNoMr8xEvpR4/kvLhe5SWAL28C
BGCcoPajtfFhUxvltYZSdxk8ygY6SUBL72OlQiu0Z5+EK+bTF0l0fiE5BHUj4Lyk
w25KbBhR13B2VuV8XP854FSot6JdAz6OK4Fmu3tiUtyo3fIcVbeSOS38/6pHXYTw
3HCS3yA9aCsd3p/qiEmdMsNJxazxGOPFNo4pGHRaFB0pzWjeD+HiIbJEkjo/nGV3
XOE2FcfsmK7rQRJ7zu7u8gOZjTJ1i5CKZ/LSY49IMvsdIAtF8x6DO5Uq4kA2SmlT
+QsRqOysjoD7q+ZNOc0W59rA1dypWuMOkcVJ9buIBn2a9YXmQ180U1I1NFsp8F5y
p5xG6dh6shkrrnQGbCiShCWDFpMv2RYflTydoGqCGjivDeSzsu9/aztfpo0/85AT
Q1XvZnMw6/5oclqiz/uxKoSkyR4xM6ZQVkfGq4ntjypaF4O6+74Pkx1LzLvJx1y2
Hd7BH08RBddTEZvBNlQPgKltuJbVXiKXxzafKL93Vk8dA2Vqwwo5saY4iH0QVq3z
UGk74Yf1/kqL37EPwLKhOjW6dVAgIKKDdTv1IM3ixGe5OR48mHS82NNdxOvzh0AZ
nJl6Rq4hEMJz4MaYEj97QbsTxzSYbuUf7VwmMDX8aA1DWBVq/65bJw2k9T1q2yer
oPFPsaFRYGJrJ9RpvlWyoK71rWOLGTkcQSVtfr2Nq2HVE/06AtgqPqFwGsQy4b5U
+ByEtVxnMoJDov0stmsPOlRHz/h5ibEFAU4nrNTzZ29ABzaH51S9X3tFsYSgXjmz
IVKi36x5UXeBY7Ghud7aHPSNhGS3RAQsNe4Busgx0rLPkcejNmQF3AXuj92vYTyd
lCSvSfHZyOuPtN30cbA9t4x78B32j+31e0PP9WALG0fZjatd75GoO98mTBhvJ60D
OX/L1RkH+3r87Bjar9SdCcxh+8kpvD80upkdM4kDZCGeeCv+P8+FiQzqgXcteAlp
zaqJdshc85oCJLKuIJIlm0ipHONPRwYnrtRj9Hi/wQJY095bw0yE/uZ8TOtAOfLb
WyZdkiJgm45xfFKS4XK7VG88fC+31JxV/oLKtn6iNsSpz0/joDl8lIuAIM5h8Mj2
qqxxv6c0loRK4R+cqmaLcr/9CiLfQ4MEH453LLfuxX59P88ECMBNCkZTf2rL1nWM
WnsoJvqyCPS5yUdvS8ubD/qGVJ9HQ45SkqGkww/XMkiHq3Rhpn0K02sSf8dHuM4v
9c7JLT/gKaUWkJ2QNkAGHu6LnElCMH9oPfsvQ8/oNXQSD1P0IsRAJucSVg/Hh7tt
H5LazmfVHRVSWnDYNeUvUbbfNmnwkXlFIhkJZVEleOOWcAq+MEQEzaMEXfHj6nb8
wwZPD1ZXYKEfCbf+OHotz/uajk1WCUGAwA8xT6KJBwVBV9JG+Vvk9Kxylm8+GHfo
uF8FSFKXQH4ePANksP3UfWwInQiidr77H1a2oYQvEoIgC/cBG9em6rILvgsKqj9Z
R1M3bs/6+RLmH3T7yCTTGQ67lbPJ0g5lU/solZkrgJcU/KuB++RqFcpBU8mHDPNm
jBcdkBhxdwtArAUIgq4d1IXs3R3myprdckuUqoUYqYRFEcklyhG/Abrp49eyxv7v
WnhAT1rDrvLFm3mBoAwnxJ6horOjZn2c6otvSDWJ2X67Rc1magc3mAIbIDBUgEQ0
MgnFuYhWxJo9V5XOmzJh6YjYJGyTSE9yQwOM2sW6BfB2AS/gEAUDQLf3MiTgLf4z
9I1QnX1Cq7ewwLBWkc/3rf2ieovTYaCSAEtFoBYEm7w6bQb3R7Iv+9XSYo3QhDRu
pycDQiAQkgFNOJ5qP/frnvnlGiB3kVY1/4h7mwUMCEKUTQDwT8xvEUUj84ILABLo
IGP2MTPUWgEtoEvMlGS0CudyLF7drIpS4/+dYUyKZz51hPVcSxO1qaAK4MGMqOa4
MshI45F0SPbVbF1AUESU330ICT/BEqV4BKO8p0sbRdjlpgdk0SBk2GvokOsNqBd3
ZRIQcIggw6xkta1TjbxCdb39vYQmi50fFZDI8D0gAoQ1tfjPOt8t1NHNnCt977l5
pJcO2pBd1bwsT04N0f1DDjtFkwcS51/SV2HA9lOrpGPqbs9zrDbOiP+6fbo1QD+b
jLup6kJbaMjFpzdMzxEQzLtu9zgemoPkCv53DZJFLUBshWnaeOG98Rgmyxrjk2AP
MtshXLWS3w3F+Ct+mf10xq70pH/RSBa2QoAoGjvCjNKAchPMHsRUe3fZEpSiT+Mv
DdHn54YYC3IZsRJzYSk5WpXm+UnCbBzJ0n/BPS5jjtUkUJRVxVCRtX0pjOsCYyf+
hs68EtbE6JaUhWkEEoGrJvmzPUjVlB2fQ4eQ5AfFJjp7nz38AttCTAOYS1P9NyEu
GZ3oGunHAAc8pJ8/dP/MEEF2oIfh3ipJoUXkwHRZiCfTYyPcO1pWhokT+Ade0BxF
3VVHjc11O0XfyTMyuw6Ef9/M+fnysMB3C1do4xQY6JlGxjCI6inGH5FbccEvyzwi
ivOe5ZEGXqqJ44uYlSHyRURBJptzPHdaLjnVkviGEtqHUWrA3fre8sn1Mhuyc/dL
CZvelGD52utxGCRSD4b6q5nlYxZ/196QOH6xmx31XUeL1NkPLNvKi+AW60xxDv3a
poxUfVEWPdhwlV+g4SROEz1nxipmmwTb148K1f95omMGQvMloRg8PqU5qsLrZ6/M
+GHa6FBrv1jVS47C2KMNaSAa4gbGwVmLlt31TY90uachX1ds8g3SXxOXMD7xNmRb
5cQQkH709/uuJUFdGFHT7Wh1HMFTBT26PD1MwIoLR0p8koTIBwxHjhKWir9JaEQy
rIQAa1xLkzq9FHNgbkzHJVqleqzAj9m+1vRIE2EpKfXJKIVephCliLJG2vPfA7cG
8v0cFuS/k4BB/hl+Mgx00pXGFkZS5i5xxAnvrBoIe9IMFHic8GsO69WOvxLJz3jC
195/IVhwQ2CBljgrVarqmOQS8lAymxMsv5PYMEGFMUKDoLVlu8jXVzdI32ty+Tgv
hXKYXdkwY+Ij4kLTVogkpKNRrQwuh6Oon/zMLGFdheio+L29+cyZG3SzbG9wPqgQ
ylsgjUaBzGw2MXzwknn8Etz6nk3XxFrUeNeUSNuNdv9+ZHWkIXkk+0n0hL2xj8At
k0MMEnXSW9pGqRxfP8vV8LtLdMzcIKe2vnN0Tazpc6CXp6HsYreDPtNY9gHDfJdD
8DpNMcPFQvUMSfkKvZSRPC6xlUF3EGDvqcq2Rxx4kl/+ZXzYUGKei8wfrATlET7n
LYuGogurbbvxq9ESeUcmYlG934BVzZ/O77Ioo/i+0HGFZfEzvBVrJL8t2wIAPD3V
9sYcOnG5VXv+SzykuAz7iU+SpY+6NK6+PyvG7T6W6UN7iHAlV2rnOlUT7FfUZKmT
dY617zDfRsZgNOnWRqctw68iVbdQQYRYsFgKQMuh9AOLG0u4FbZhyrdQ3jQmdUUz
zRDGUi01XKoLBfhSod8d7EPJqaVjRbKcwpu2dBfFToGHzKmjQBtQa+ua4mpQO4Xc
b/7SPRoi1Odp03AL5FfgwSxQnOwAYjvGB2jVXKDxOCFctjb4awRHR1uIUMHsUoh5
XewyDkCI5+wJvulI7b37hhrCCMv6gXPqPTPYNNSapWogDbUqHeZMdxDvNosFFP9L
C/VCULEWSnPgGpTjImIsyZqRvhLIVa2hLM29VTx0d9LKRLtStbEST4LCjklyJu22
K13rczoJAvFjDAJHGfxcIW8HVsU8cyaxgI7YiC+F6WEqzZIuzvySjADJENO5/T0I
IG/2BXigvrqCoVFhxqjiBFGySLzgWPbKHRoOc6cHncnZ+2ZR5JkYNf8P9QGBGgg8
4n4KGG5IrcG0G2H58hV05Y1iFyTXIbs2JdHQ3X5+4c5Up3HPkTRMnzsGwk0LjfBo
yEDQduwTKgns+w+hTgQl1gZBH8/gMIHtgekF03Dht3yzodn5/+Wot2b08yryzegw
gJRr11XgNqYnFI0BBQHe/5IBPiEFkWaKGRWK6qXd6Mr7XQ5jvUeQq6MrJgPNWZ9A
npzenxjhTdanR10FUBvQ5uqzLZg4qSCKNzgWzXm585n01yYvtsBgHMnyVLSFgCq5
8SciWTHM9demtkhttuiRmHgjjhbJr1FH0VVBCdTmOLAao+RuWIkT3RLIQCxKUs6f
NISzpjXmVTG8vGg76uwgUZ1tOtz1YAWUsj0moRNNe8AklX10jfNdtUla1zxYZ4Ez
4FO/tGKKzZO5WPqEjAsdWOufQet1Ljvtc8LCuYb0fbJlvA2qlen+wLNwpYB+SgBz
XVEluBfAmy65mHot2e5/DQBdE3W/ne5ijex3t2sBbusInBhd3e9m13QrtvRCJOT2
Is/7JXf+wiVCXDRFgt8X9LtB9qVOlem7WnV9WN9lhEfo4TDOVqBwR1TlzWu7yiSZ
IxiIIXVGS8cOocbYi6D9ZCkCkAJ330lNr0JNwiXH7cOsDql4bHD6bra8YRZQEICI
e3q/2VDzpM/BdqXOn3GVhbX7uba+wieCQZWGZWGdryonocua8w185j+VjFHgSwMO
YYiUrtz8gnaGAWc8vlp55wVgWPXQ6E7jhxjtvRWoALVs01WFM+nT7+ZNgpicaL6k
3+i2evmJdr6lQQI8Wb5E9/I72AcbJpGzohA4rB6QkbAoyJMMStp4A570kzn/Q78Q
qeZ2OxR2t8T6sKQRf/INojMuEQR1NHxGBmCa8RmNQeSTTFQPZznE+50VYmoksygF
8sQwltkVt9o8YQc0nRoF5fGcyZf/Fszs3htVsXayFC+DJB7ox4VuqbKsljFGV2nN
NoQc87k7IyOWFJ0TLtb2yTXEd/JYjD6BX0Pf9zazZg3rny6Mp1AAa1CadIsUEzrg
HeJx/f65Ju7/HKAYn+1QYCSmj4yFTSjye5krjtSFUPCy9K5gU17rEZF0VjsryStn
OVdyA6nsHl6wRDdLaUm/VkNQialbXan46NRNSgspJCssj82eF2t0x8eiQif+cWUC
SWYp/auTpsbagGcULs6l7Ai8LzcPanomgdt9zjUzqwmUY90PIAsLJmt0H5VM/dlH
dVZ4D/qxq1uFniaoQa7Ve5SGyDtK43MTxEzVdNovclBG1/dGv2fXY60xRhmnq1QF
DUOo6duB4ipF/HNSGLccKNSes6ornJ4iPZfMKWrz9tSBGw0UzMaSMgiRwG3hUfoj
`protect END_PROTECTED
