`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEdOrv0yWUHZxaGAg4XcgTETTYvP01G2QBhWvrdGWwzI
0rrz+6uIJ6Scm/5jz/gKG31jqnp+P0RlHjOd0n09FCA1MWTCMs+wolH8E19/e12/
tJuQBga+CQxaFwL7BrDYr88jb9rU32HsuQIXKe26d6P5WcFjL5x7ZEA4Rd2lGSLc
SIE/zyhoTOxft2WfEOHKRtWLpuGwcCB/ihnxuMM5oMsE7NsCfDTFy+pfOUy/zsSV
XxtIBIhKKlpyHgZ1br6uzpMC18EEbHJGBi4CtWlZbkw3sZB+Gu7va98RZ8xMdbdK
E53gKAlqilDp5ToAo02rlxB6+kA6z2qzFe/GKG48xbv6vviwFQ3oaQ2v3AaGtCBG
gaSTSHaA5l8bnpRKyVn9ilY6y8NCGviiwTLERJfxT1jP3znmCfmCEGr4uB3Dn8Xm
0MRcS0wMOZU9W85eqcGtf0qcfgiSm8xEQKSE7iruO8T/3b5ygN2/e3T9BOttdSXi
uDKJuIArgmyeFxuCsFoa4PevmgQWtwduXCIS1rPGp2AzR5OruICEKiRfEANaMQDW
LPRwhaBm9oVjdVMLcsqp2qyJ1x/A0PC4lQWr5IlAeFff7ML4wdIRJ8/9dIqyDG86
NSzPO/7dAU77vkWkp7E6csKu/Mut/9GdqgeS7dEB/c8sTRoRVHtwaYk+rfdHNnWu
cj+19OnYtbIhv9xNJ+04lWjHJT6IkA7a/tTZy3IVJBL3BYOYXdCHQ4gndCYivmXr
A5sbeCXDj5mY2ofDukJ15oOUz27Fqauv+5vkVJMxsdiLeOJYVoBF4h75lHivyswI
tLAI6SRBsltvDVon2gZJBQdvtbnwV2C/peX9GAwdv3E=
`protect END_PROTECTED
