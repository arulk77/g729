`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
WwByT+ldZGlKIY2PikOP3JCYzxUFe9++acl/BGCkVGM4pFFx7dDEtCdPK1YB6Rt9
oCIrxcwzLAl4E4BK4d8pSquTJKVE+WOtMd9djQVoj+X/Xz7sa6ABQARIPRTXxxLq
Wfu12qIz2Y4t21aOtO8qA7z+AdrYDxnT/OGBR1SuBxx5yJZy7FU914y0d3kWLMI3
dlM+R5drUs73n2qSrJU8wnM1hm4rD1LopJi5yF6v5hAbs9+aAle39DhxGWEeSdv8
wD+hL9tvsIIqreY+Xu176/SAnrfBdTJG3GsVEOES+//K3q9cvCjbrOYLVg3FCgcY
5XxhAWBtTJKd1EKscGYxrPu8M2hQx72lbVwshKVDRhk=
`protect END_PROTECTED
