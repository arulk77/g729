`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
haMrRDHspd1e7e2RO53oiHEyF5nGV6oaFmGk5gvt/DGmqvuhTqjLDvhRVTTMmgry
ChjcIhC87FAa35M2xGLRrpeSKtSJbzuiosO3Zq55B2YZUvzQcZ0lejr+R8oASPZc
aAvfuydSibyI6Xj1GmNOrvl+bflG6MTnqrPz8WykMEfvWb35J7vnSPozX1MJ1WwR
FYcAAsuDWWbj6ugUOvA2JBoNVu14JTp4AH1rmzHprAvYS4DXOGxiOMZEhdORxMRT
PlrUwJBmpDd4WUEnb2VsU3FMN9/Lq6oUaPBNx5JKiEklaKGpp+UushoLgI+9faYL
3EWNxVF3uf1Mm3AX+1uJ3qP1KWicsehPRzFIkfFaGrnvIJZ8h2zoX6GdU9A8btQo
WSKFYULcGzQ9d7NVT19qLkZEwFneISPnQ6/2Dk6McBzS9t5W7l7EofF6BV5Js14a
QywjE8qhmQqWRCWuZ3wCFx4Zqsrx+GXW0XicOrmplbzF4n8cBINYg47jGvnatFid
r1eIUk4O5M61dUAkv3TmULnS7KD6o/nzynkUluYbajMtHEcxTu5XExbme/ju/LRK
hNuzlVY0yeOgcFBuSEfTHcpixo/KXR1fqX4P5gH0Mb5fc5DPJfu8eu/U95Ust+zE
y990PkCM3hVct0Ph8kDtuoMFUiLiHJKMxVSas7hRO6tDynGMKiqgoTvnjelIlAwU
pRD6XnaJsG/p9azMdZlHZ2CW+A66b8Yd6OzFOU2RFKXOBOjjHeeBQC1O6WAzjJWt
uqJgKM6IuX1nBPgXiU+dvw==
`protect END_PROTECTED
