`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAm0te0xdTeTHab4uNgXXCjJ3YR/gu7Y/0RWfGOD4rbM
WSx3d+HE5Tz/r/0JdXnrkth2GBbrsXz7j15gksSi2VdcC73sE6q85jBIuc4Q+g/F
XoiaID9LXXXrqfkusKDBKADKRO7hzmNgln6/NJ5YR+ixBQG5+fRUn5vVadJggU6y
rRk5qebOpN7k7M15NLlQ6aRreglJkyeUdazbasCvCbUpFInUJMTGKfNl09bKCTVO
Robbe04I2wTSLWiS1IwdKBl5YVHE6aILfW0WnjkUboH7qGF5RaK5l5dKf4IgjfLn
9+zdpZtXWzBpvHaMlv9RwREKeGt+k0ol4oIwKRtp92xd/hvaoUddZgInl4lSiyNj
IVpMd3Y45oydRqGocVKszIiHFd2LCj1lFBuL9NqXO4L3vWXFsNGDXaUnJFwzTLba
2FETXmmrEkNX8XON3a8AXvRUDxfC1cSfM41HrouRSSiDggdWAYC8csxoAj9EnR3S
HQboJ0gbT5IegkuPEhYcU6JBZjAVPpG+ItoUrskWcYaq/rWknl91kDK2G9kcR/nj
fOfcBXFVAdJwmt1XXB0yjqZJnWdKxsVcKrOVooAqotA=
`protect END_PROTECTED
