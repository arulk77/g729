`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKaEL8HOsVjLT8JVJaSs3DdrPfZQufEihDpiXF0GZBew
12I8r1hVDx87G8YiLFKvn2LM8bzrv9I2MrUjMdSUMu0T5pzRPGlo+kihNZjxikFx
pfElD2zZU5hzKQMCNiHar/6IxXV2uvC2sVZL8GCkPEXFhinZosUGaK6Iq1dq7V+9
2QyZGqnI/5C1yGULoo0WMyn9APXqcE1iJ5FsUkxD8Jlf4yPz564GMtzNF6x68q2S
`protect END_PROTECTED
