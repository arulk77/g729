library verilog;
use verilog.vl_types.all;
entity PCIE_EP is
    generic(
        BAR0EXIST       : string  := "TRUE";
        BAR0PREFETCHABLE: string  := "TRUE";
        BAR1EXIST       : string  := "FALSE";
        BAR1PREFETCHABLE: string  := "FALSE";
        BAR2EXIST       : string  := "FALSE";
        BAR2PREFETCHABLE: string  := "FALSE";
        BAR3EXIST       : string  := "FALSE";
        BAR3PREFETCHABLE: string  := "FALSE";
        BAR4EXIST       : string  := "FALSE";
        BAR4PREFETCHABLE: string  := "FALSE";
        BAR5EXIST       : string  := "FALSE";
        BAR5PREFETCHABLE: string  := "FALSE";
        CLKDIVIDED      : string  := "FALSE";
        INFINITECOMPLETIONS: string  := "TRUE";
        LINKSTATUSSLOTCLOCKCONFIG: string  := "FALSE";
        PBCAPABILITYSYSTEMALLOCATED: string  := "FALSE";
        PMCAPABILITYD1SUPPORT: string  := "FALSE";
        PMCAPABILITYD2SUPPORT: string  := "FALSE";
        PMCAPABILITYDSI : string  := "TRUE";
        RESETMODE       : string  := "FALSE";
        VC0TOTALCREDITSCD: integer := 0;
        VC0TOTALCREDITSPD: integer := 52;
        VC1TOTALCREDITSCD: integer := 0;
        VC1TOTALCREDITSPD: integer := 0;
        AERBASEPTR      : integer := 272;
        AERCAPABILITYNEXTPTR: integer := 312;
        DSNBASEPTR      : integer := 328;
        DSNCAPABILITYNEXTPTR: integer := 340;
        MSIBASEPTR      : integer := 72;
        PBBASEPTR       : integer := 312;
        PBCAPABILITYNEXTPTR: integer := 328;
        PMBASEPTR       : integer := 64;
        RETRYRAMSIZE    : integer := 9;
        VCBASEPTR       : integer := 340;
        VCCAPABILITYNEXTPTR: integer := 0;
        VC0RXFIFOBASEC  : integer := 152;
        VC0RXFIFOBASENP : integer := 128;
        VC0RXFIFOBASEP  : integer := 0;
        VC0RXFIFOLIMITC : integer := 279;
        VC0RXFIFOLIMITNP: integer := 151;
        VC0RXFIFOLIMITP : integer := 127;
        VC0TXFIFOBASEC  : integer := 152;
        VC0TXFIFOBASENP : integer := 128;
        VC0TXFIFOBASEP  : integer := 0;
        VC0TXFIFOLIMITC : integer := 279;
        VC0TXFIFOLIMITNP: integer := 151;
        VC0TXFIFOLIMITP : integer := 127;
        VC1RXFIFOBASEC  : integer := 280;
        VC1RXFIFOBASENP : integer := 280;
        VC1RXFIFOBASEP  : integer := 280;
        VC1RXFIFOLIMITC : integer := 280;
        VC1RXFIFOLIMITNP: integer := 280;
        VC1RXFIFOLIMITP : integer := 280;
        VC1TXFIFOBASEC  : integer := 280;
        VC1TXFIFOBASENP : integer := 280;
        VC1TXFIFOBASEP  : integer := 280;
        VC1TXFIFOLIMITC : integer := 280;
        VC1TXFIFOLIMITNP: integer := 280;
        VC1TXFIFOLIMITP : integer := 280;
        DEVICEID        : integer := 20560;
        SUBSYSTEMID     : integer := 20560;
        SUBSYSTEMVENDORID: integer := 4334;
        VENDORID        : integer := 4334;
        LINKCAPABILITYASPMSUPPORT: integer := 1;
        PBCAPABILITYDW0DATASCALE: integer := 0;
        PBCAPABILITYDW0PMSTATE: integer := 0;
        PBCAPABILITYDW1DATASCALE: integer := 0;
        PBCAPABILITYDW1PMSTATE: integer := 0;
        PBCAPABILITYDW2DATASCALE: integer := 0;
        PBCAPABILITYDW2PMSTATE: integer := 0;
        PBCAPABILITYDW3DATASCALE: integer := 0;
        PBCAPABILITYDW3PMSTATE: integer := 0;
        CLASSCODE       : integer := 360448;
        DEVICECAPABILITYENDPOINTL0SLATENCY: integer := 0;
        DEVICECAPABILITYENDPOINTL1LATENCY: integer := 0;
        MSICAPABILITYMULTIMSGCAP: integer := 0;
        PBCAPABILITYDW0PMSUBSTATE: integer := 0;
        PBCAPABILITYDW0POWERRAIL: integer := 0;
        PBCAPABILITYDW0TYPE: integer := 0;
        PBCAPABILITYDW1PMSUBSTATE: integer := 0;
        PBCAPABILITYDW1POWERRAIL: integer := 0;
        PBCAPABILITYDW1TYPE: integer := 0;
        PBCAPABILITYDW2PMSUBSTATE: integer := 0;
        PBCAPABILITYDW2POWERRAIL: integer := 0;
        PBCAPABILITYDW2TYPE: integer := 0;
        PBCAPABILITYDW3PMSUBSTATE: integer := 0;
        PBCAPABILITYDW3POWERRAIL: integer := 0;
        PBCAPABILITYDW3TYPE: integer := 0;
        PMCAPABILITYAUXCURRENT: integer := 0;
        PORTVCCAPABILITYEXTENDEDVCCOUNT: integer := 0;
        CARDBUSCISPOINTER: integer := 0;
        XPDEVICEPORTTYPE: integer := 0;
        PMCAPABILITYPMESUPPORT: integer := 0;
        BAR0MASKWIDTH   : integer := 20;
        BAR1MASKWIDTH   : integer := 0;
        BAR2MASKWIDTH   : integer := 0;
        BAR3MASKWIDTH   : integer := 0;
        BAR4MASKWIDTH   : integer := 0;
        BAR5MASKWIDTH   : integer := 0;
        LINKCAPABILITYMAXLINKWIDTH: integer := 1;
      --DEVICESERIALNUMBER: integer type with unrepresentable value!
        VC0TOTALCREDITSCH: integer := 0;
        VC0TOTALCREDITSNPH: integer := 8;
        VC0TOTALCREDITSPH: integer := 8;
        VC1TOTALCREDITSCH: integer := 0;
        VC1TOTALCREDITSNPH: integer := 0;
        VC1TOTALCREDITSPH: integer := 0;
        ACTIVELANESIN   : integer := 1;
        CAPABILITIESPOINTER: integer := 64;
        INTERRUPTPIN    : integer := 0;
        MSICAPABILITYNEXTPTR: integer := 96;
        PBCAPABILITYDW0BASEPOWER: integer := 0;
        PBCAPABILITYDW1BASEPOWER: integer := 0;
        PBCAPABILITYDW2BASEPOWER: integer := 0;
        PBCAPABILITYDW3BASEPOWER: integer := 0;
        PCIECAPABILITYNEXTPTR: integer := 0;
        PMCAPABILITYNEXTPTR: integer := 96;
        PMDATA0         : integer := 0;
        PMDATA1         : integer := 0;
        PMDATA2         : integer := 0;
        PMDATA3         : integer := 0;
        PMDATA4         : integer := 0;
        PMDATA5         : integer := 0;
        PMDATA6         : integer := 0;
        PMDATA7         : integer := 0;
        PORTVCCAPABILITYVCARBCAP: integer := 0;
        PORTVCCAPABILITYVCARBTABLEOFFSET: integer := 0;
        REVISIONID      : integer := 0;
        XPBASEPTR       : integer := 96;
        BAR0ADDRWIDTH   : integer := 0;
        BAR0IOMEMN      : integer := 0;
        BAR1ADDRWIDTH   : integer := 0;
        BAR1IOMEMN      : integer := 0;
        BAR2ADDRWIDTH   : integer := 0;
        BAR2IOMEMN      : integer := 0;
        BAR3ADDRWIDTH   : integer := 0;
        BAR3IOMEMN      : integer := 0;
        BAR4ADDRWIDTH   : integer := 0;
        BAR4IOMEMN      : integer := 0;
        BAR5IOMEMN      : integer := 0;
        L0SEXITLATENCY  : integer := 7;
        L0SEXITLATENCYCOMCLK: integer := 7;
        L1EXITLATENCY   : integer := 7;
        L1EXITLATENCYCOMCLK: integer := 7;
        LOWPRIORITYVCCOUNT: integer := 0;
        PMDATASCALE0    : integer := 0;
        PMDATASCALE1    : integer := 0;
        PMDATASCALE2    : integer := 0;
        PMDATASCALE3    : integer := 0;
        PMDATASCALE4    : integer := 0;
        PMDATASCALE5    : integer := 0;
        PMDATASCALE6    : integer := 0;
        PMDATASCALE7    : integer := 0;
        RETRYRAMREADLATENCY: integer := 3;
        RETRYRAMWRITELATENCY: integer := 1;
        TLRAMREADLATENCY: integer := 3;
        TLRAMWRITELATENCY: integer := 1;
        TXTSNFTS        : integer := 255;
        TXTSNFTSCOMCLK  : integer := 255;
        XPMAXPAYLOAD    : integer := 0
    );
    port(
        BUSMASTERENABLE : out    vl_logic;
        CRMDOHOTRESETN  : out    vl_logic;
        CRMPWRSOFTRESETN: out    vl_logic;
        DLLTXPMDLLPOUTSTANDING: out    vl_logic;
        INTERRUPTDISABLE: out    vl_logic;
        IOSPACEENABLE   : out    vl_logic;
        L0CFGLOOPBACKACK: out    vl_logic;
        L0COMPLETERID   : out    vl_logic_vector(12 downto 0);
        L0DLLERRORVECTOR: out    vl_logic_vector(6 downto 0);
        L0DLLRXACKOUTSTANDING: out    vl_logic;
        L0DLLTXNONFCOUTSTANDING: out    vl_logic;
        L0DLLTXOUTSTANDING: out    vl_logic;
        L0DLLVCSTATUS   : out    vl_logic_vector(7 downto 0);
        L0DLUPDOWN      : out    vl_logic_vector(7 downto 0);
        L0FIRSTCFGWRITEOCCURRED: out    vl_logic;
        L0LTSSMSTATE    : out    vl_logic_vector(3 downto 0);
        L0MACENTEREDL0  : out    vl_logic;
        L0MACLINKTRAINING: out    vl_logic;
        L0MACLINKUP     : out    vl_logic;
        L0MACNEGOTIATEDLINKWIDTH: out    vl_logic_vector(3 downto 0);
        L0MACNEWSTATEACK: out    vl_logic;
        L0MACRXL0SSTATE : out    vl_logic;
        L0MSIENABLE0    : out    vl_logic;
        L0MULTIMSGEN0   : out    vl_logic_vector(2 downto 0);
        L0PMEACK        : out    vl_logic;
        L0PMEEN         : out    vl_logic;
        L0PMEREQOUT     : out    vl_logic;
        L0PWRL1STATE    : out    vl_logic;
        L0PWRL23READYSTATE: out    vl_logic;
        L0PWRSTATE0     : out    vl_logic_vector(1 downto 0);
        L0PWRTURNOFFREQ : out    vl_logic;
        L0PWRTXL0SSTATE : out    vl_logic;
        L0RXDLLPM       : out    vl_logic;
        L0RXDLLPMTYPE   : out    vl_logic_vector(2 downto 0);
        L0RXMACLINKERROR: out    vl_logic_vector(1 downto 0);
        L0STATSCFGOTHERRECEIVED: out    vl_logic;
        L0STATSCFGOTHERTRANSMITTED: out    vl_logic;
        L0STATSCFGRECEIVED: out    vl_logic;
        L0STATSCFGTRANSMITTED: out    vl_logic;
        L0STATSDLLPRECEIVED: out    vl_logic;
        L0STATSDLLPTRANSMITTED: out    vl_logic;
        L0STATSOSRECEIVED: out    vl_logic;
        L0STATSOSTRANSMITTED: out    vl_logic;
        L0STATSTLPRECEIVED: out    vl_logic;
        L0STATSTLPTRANSMITTED: out    vl_logic;
        L0UNLOCKRECEIVED: out    vl_logic;
        LLKRXCHCOMPLETIONAVAILABLEN: out    vl_logic_vector(7 downto 0);
        LLKRXCHNONPOSTEDAVAILABLEN: out    vl_logic_vector(7 downto 0);
        LLKRXCHPOSTEDAVAILABLEN: out    vl_logic_vector(7 downto 0);
        LLKRXDATA       : out    vl_logic_vector(63 downto 0);
        LLKRXEOFN       : out    vl_logic;
        LLKRXEOPN       : out    vl_logic;
        LLKRXPREFERREDTYPE: out    vl_logic_vector(15 downto 0);
        LLKRXSOFN       : out    vl_logic;
        LLKRXSOPN       : out    vl_logic;
        LLKRXSRCLASTREQN: out    vl_logic;
        LLKRXSRCRDYN    : out    vl_logic;
        LLKRXVALIDN     : out    vl_logic_vector(1 downto 0);
        LLKTCSTATUS     : out    vl_logic_vector(7 downto 0);
        LLKTXCHANSPACE  : out    vl_logic_vector(9 downto 0);
        LLKTXCHCOMPLETIONREADYN: out    vl_logic_vector(7 downto 0);
        LLKTXCHNONPOSTEDREADYN: out    vl_logic_vector(7 downto 0);
        LLKTXCHPOSTEDREADYN: out    vl_logic_vector(7 downto 0);
        LLKTXCONFIGREADYN: out    vl_logic;
        LLKTXDSTRDYN    : out    vl_logic;
        MAXPAYLOADSIZE  : out    vl_logic_vector(2 downto 0);
        MAXREADREQUESTSIZE: out    vl_logic_vector(2 downto 0);
        MEMSPACEENABLE  : out    vl_logic;
        MGMTPSO         : out    vl_logic_vector(16 downto 0);
        MGMTRDATA       : out    vl_logic_vector(31 downto 0);
        MGMTSTATSCREDIT : out    vl_logic_vector(11 downto 0);
        MIMDLLBRADD     : out    vl_logic_vector(11 downto 0);
        MIMDLLBREN      : out    vl_logic;
        MIMDLLBWADD     : out    vl_logic_vector(11 downto 0);
        MIMDLLBWDATA    : out    vl_logic_vector(63 downto 0);
        MIMDLLBWEN      : out    vl_logic;
        MIMRXBRADD      : out    vl_logic_vector(12 downto 0);
        MIMRXBREN       : out    vl_logic;
        MIMRXBWADD      : out    vl_logic_vector(12 downto 0);
        MIMRXBWDATA     : out    vl_logic_vector(63 downto 0);
        MIMRXBWEN       : out    vl_logic;
        MIMTXBRADD      : out    vl_logic_vector(12 downto 0);
        MIMTXBREN       : out    vl_logic;
        MIMTXBWADD      : out    vl_logic_vector(12 downto 0);
        MIMTXBWDATA     : out    vl_logic_vector(63 downto 0);
        MIMTXBWEN       : out    vl_logic;
        PARITYERRORRESPONSE: out    vl_logic;
        PIPEDESKEWLANESL0: out    vl_logic;
        PIPEDESKEWLANESL1: out    vl_logic;
        PIPEDESKEWLANESL2: out    vl_logic;
        PIPEDESKEWLANESL3: out    vl_logic;
        PIPEDESKEWLANESL4: out    vl_logic;
        PIPEDESKEWLANESL5: out    vl_logic;
        PIPEDESKEWLANESL6: out    vl_logic;
        PIPEDESKEWLANESL7: out    vl_logic;
        PIPEPOWERDOWNL0 : out    vl_logic_vector(1 downto 0);
        PIPEPOWERDOWNL1 : out    vl_logic_vector(1 downto 0);
        PIPEPOWERDOWNL2 : out    vl_logic_vector(1 downto 0);
        PIPEPOWERDOWNL3 : out    vl_logic_vector(1 downto 0);
        PIPEPOWERDOWNL4 : out    vl_logic_vector(1 downto 0);
        PIPEPOWERDOWNL5 : out    vl_logic_vector(1 downto 0);
        PIPEPOWERDOWNL6 : out    vl_logic_vector(1 downto 0);
        PIPEPOWERDOWNL7 : out    vl_logic_vector(1 downto 0);
        PIPERESETL0     : out    vl_logic;
        PIPERESETL1     : out    vl_logic;
        PIPERESETL2     : out    vl_logic;
        PIPERESETL3     : out    vl_logic;
        PIPERESETL4     : out    vl_logic;
        PIPERESETL5     : out    vl_logic;
        PIPERESETL6     : out    vl_logic;
        PIPERESETL7     : out    vl_logic;
        PIPERXPOLARITYL0: out    vl_logic;
        PIPERXPOLARITYL1: out    vl_logic;
        PIPERXPOLARITYL2: out    vl_logic;
        PIPERXPOLARITYL3: out    vl_logic;
        PIPERXPOLARITYL4: out    vl_logic;
        PIPERXPOLARITYL5: out    vl_logic;
        PIPERXPOLARITYL6: out    vl_logic;
        PIPERXPOLARITYL7: out    vl_logic;
        PIPETXCOMPLIANCEL0: out    vl_logic;
        PIPETXCOMPLIANCEL1: out    vl_logic;
        PIPETXCOMPLIANCEL2: out    vl_logic;
        PIPETXCOMPLIANCEL3: out    vl_logic;
        PIPETXCOMPLIANCEL4: out    vl_logic;
        PIPETXCOMPLIANCEL5: out    vl_logic;
        PIPETXCOMPLIANCEL6: out    vl_logic;
        PIPETXCOMPLIANCEL7: out    vl_logic;
        PIPETXDATAKL0   : out    vl_logic;
        PIPETXDATAKL1   : out    vl_logic;
        PIPETXDATAKL2   : out    vl_logic;
        PIPETXDATAKL3   : out    vl_logic;
        PIPETXDATAKL4   : out    vl_logic;
        PIPETXDATAKL5   : out    vl_logic;
        PIPETXDATAKL6   : out    vl_logic;
        PIPETXDATAKL7   : out    vl_logic;
        PIPETXDATAL0    : out    vl_logic_vector(7 downto 0);
        PIPETXDATAL1    : out    vl_logic_vector(7 downto 0);
        PIPETXDATAL2    : out    vl_logic_vector(7 downto 0);
        PIPETXDATAL3    : out    vl_logic_vector(7 downto 0);
        PIPETXDATAL4    : out    vl_logic_vector(7 downto 0);
        PIPETXDATAL5    : out    vl_logic_vector(7 downto 0);
        PIPETXDATAL6    : out    vl_logic_vector(7 downto 0);
        PIPETXDATAL7    : out    vl_logic_vector(7 downto 0);
        PIPETXDETECTRXLOOPBACKL0: out    vl_logic;
        PIPETXDETECTRXLOOPBACKL1: out    vl_logic;
        PIPETXDETECTRXLOOPBACKL2: out    vl_logic;
        PIPETXDETECTRXLOOPBACKL3: out    vl_logic;
        PIPETXDETECTRXLOOPBACKL4: out    vl_logic;
        PIPETXDETECTRXLOOPBACKL5: out    vl_logic;
        PIPETXDETECTRXLOOPBACKL6: out    vl_logic;
        PIPETXDETECTRXLOOPBACKL7: out    vl_logic;
        PIPETXELECIDLEL0: out    vl_logic;
        PIPETXELECIDLEL1: out    vl_logic;
        PIPETXELECIDLEL2: out    vl_logic;
        PIPETXELECIDLEL3: out    vl_logic;
        PIPETXELECIDLEL4: out    vl_logic;
        PIPETXELECIDLEL5: out    vl_logic;
        PIPETXELECIDLEL6: out    vl_logic;
        PIPETXELECIDLEL7: out    vl_logic;
        SERRENABLE      : out    vl_logic;
        URREPORTINGENABLE: out    vl_logic;
        AUXPOWER        : in     vl_logic;
        COMPLIANCEAVOID : in     vl_logic;
        CRMCORECLK      : in     vl_logic;
        CRMCORECLKDLO   : in     vl_logic;
        CRMCORECLKRXO   : in     vl_logic;
        CRMCORECLKTXO   : in     vl_logic;
        CRMLINKRSTN     : in     vl_logic;
        CRMMACRSTN      : in     vl_logic;
        CRMMGMTRSTN     : in     vl_logic;
        CRMNVRSTN       : in     vl_logic;
        CRMURSTN        : in     vl_logic;
        CRMUSERCFGRSTN  : in     vl_logic;
        CRMUSERCLK      : in     vl_logic;
        CRMUSERCLKRXO   : in     vl_logic;
        CRMUSERCLKTXO   : in     vl_logic;
        L0CFGDISABLESCRAMBLE: in     vl_logic;
        L0CFGLOOPBACKMASTER: in     vl_logic;
        L0LEGACYINTFUNCT0: in     vl_logic;
        L0MSIREQUEST0   : in     vl_logic_vector(3 downto 0);
        L0PACKETHEADERFROMUSER: in     vl_logic_vector(127 downto 0);
        L0PMEREQIN      : in     vl_logic;
        L0SETCOMPLETERABORTERROR: in     vl_logic;
        L0SETCOMPLETIONTIMEOUTCORRERROR: in     vl_logic;
        L0SETCOMPLETIONTIMEOUTUNCORRERROR: in     vl_logic;
        L0SETDETECTEDCORRERROR: in     vl_logic;
        L0SETDETECTEDFATALERROR: in     vl_logic;
        L0SETDETECTEDNONFATALERROR: in     vl_logic;
        L0SETUNEXPECTEDCOMPLETIONCORRERROR: in     vl_logic;
        L0SETUNEXPECTEDCOMPLETIONUNCORRERROR: in     vl_logic;
        L0SETUNSUPPORTEDREQUESTNONPOSTEDERROR: in     vl_logic;
        L0SETUNSUPPORTEDREQUESTOTHERERROR: in     vl_logic;
        L0SETUSERDETECTEDPARITYERROR: in     vl_logic;
        L0SETUSERMASTERDATAPARITY: in     vl_logic;
        L0SETUSERRECEIVEDMASTERABORT: in     vl_logic;
        L0SETUSERRECEIVEDTARGETABORT: in     vl_logic;
        L0SETUSERSIGNALLEDTARGETABORT: in     vl_logic;
        L0SETUSERSYSTEMERROR: in     vl_logic;
        L0TRANSACTIONSPENDING: in     vl_logic;
        LLKRXCHFIFO     : in     vl_logic_vector(1 downto 0);
        LLKRXCHTC       : in     vl_logic_vector(2 downto 0);
        LLKRXDSTCONTREQN: in     vl_logic;
        LLKRXDSTREQN    : in     vl_logic;
        LLKTXCHFIFO     : in     vl_logic_vector(1 downto 0);
        LLKTXCHTC       : in     vl_logic_vector(2 downto 0);
        LLKTXDATA       : in     vl_logic_vector(63 downto 0);
        LLKTXENABLEN    : in     vl_logic_vector(1 downto 0);
        LLKTXEOFN       : in     vl_logic;
        LLKTXEOPN       : in     vl_logic;
        LLKTXSOFN       : in     vl_logic;
        LLKTXSOPN       : in     vl_logic;
        LLKTXSRCDSCN    : in     vl_logic;
        LLKTXSRCRDYN    : in     vl_logic;
        MGMTADDR        : in     vl_logic_vector(10 downto 0);
        MGMTBWREN       : in     vl_logic_vector(3 downto 0);
        MGMTRDEN        : in     vl_logic;
        MGMTSTATSCREDITSEL: in     vl_logic_vector(6 downto 0);
        MGMTWDATA       : in     vl_logic_vector(31 downto 0);
        MGMTWREN        : in     vl_logic;
        MIMDLLBRDATA    : in     vl_logic_vector(63 downto 0);
        MIMRXBRDATA     : in     vl_logic_vector(63 downto 0);
        MIMTXBRDATA     : in     vl_logic_vector(63 downto 0);
        PIPEPHYSTATUSL0 : in     vl_logic;
        PIPEPHYSTATUSL1 : in     vl_logic;
        PIPEPHYSTATUSL2 : in     vl_logic;
        PIPEPHYSTATUSL3 : in     vl_logic;
        PIPEPHYSTATUSL4 : in     vl_logic;
        PIPEPHYSTATUSL5 : in     vl_logic;
        PIPEPHYSTATUSL6 : in     vl_logic;
        PIPEPHYSTATUSL7 : in     vl_logic;
        PIPERXCHANISALIGNEDL0: in     vl_logic;
        PIPERXCHANISALIGNEDL1: in     vl_logic;
        PIPERXCHANISALIGNEDL2: in     vl_logic;
        PIPERXCHANISALIGNEDL3: in     vl_logic;
        PIPERXCHANISALIGNEDL4: in     vl_logic;
        PIPERXCHANISALIGNEDL5: in     vl_logic;
        PIPERXCHANISALIGNEDL6: in     vl_logic;
        PIPERXCHANISALIGNEDL7: in     vl_logic;
        PIPERXDATAKL0   : in     vl_logic;
        PIPERXDATAKL1   : in     vl_logic;
        PIPERXDATAKL2   : in     vl_logic;
        PIPERXDATAKL3   : in     vl_logic;
        PIPERXDATAKL4   : in     vl_logic;
        PIPERXDATAKL5   : in     vl_logic;
        PIPERXDATAKL6   : in     vl_logic;
        PIPERXDATAKL7   : in     vl_logic;
        PIPERXDATAL0    : in     vl_logic_vector(7 downto 0);
        PIPERXDATAL1    : in     vl_logic_vector(7 downto 0);
        PIPERXDATAL2    : in     vl_logic_vector(7 downto 0);
        PIPERXDATAL3    : in     vl_logic_vector(7 downto 0);
        PIPERXDATAL4    : in     vl_logic_vector(7 downto 0);
        PIPERXDATAL5    : in     vl_logic_vector(7 downto 0);
        PIPERXDATAL6    : in     vl_logic_vector(7 downto 0);
        PIPERXDATAL7    : in     vl_logic_vector(7 downto 0);
        PIPERXELECIDLEL0: in     vl_logic;
        PIPERXELECIDLEL1: in     vl_logic;
        PIPERXELECIDLEL2: in     vl_logic;
        PIPERXELECIDLEL3: in     vl_logic;
        PIPERXELECIDLEL4: in     vl_logic;
        PIPERXELECIDLEL5: in     vl_logic;
        PIPERXELECIDLEL6: in     vl_logic;
        PIPERXELECIDLEL7: in     vl_logic;
        PIPERXSTATUSL0  : in     vl_logic_vector(2 downto 0);
        PIPERXSTATUSL1  : in     vl_logic_vector(2 downto 0);
        PIPERXSTATUSL2  : in     vl_logic_vector(2 downto 0);
        PIPERXSTATUSL3  : in     vl_logic_vector(2 downto 0);
        PIPERXSTATUSL4  : in     vl_logic_vector(2 downto 0);
        PIPERXSTATUSL5  : in     vl_logic_vector(2 downto 0);
        PIPERXSTATUSL6  : in     vl_logic_vector(2 downto 0);
        PIPERXSTATUSL7  : in     vl_logic_vector(2 downto 0);
        PIPERXVALIDL0   : in     vl_logic;
        PIPERXVALIDL1   : in     vl_logic;
        PIPERXVALIDL2   : in     vl_logic;
        PIPERXVALIDL3   : in     vl_logic;
        PIPERXVALIDL4   : in     vl_logic;
        PIPERXVALIDL5   : in     vl_logic;
        PIPERXVALIDL6   : in     vl_logic;
        PIPERXVALIDL7   : in     vl_logic
    );
end PCIE_EP;
