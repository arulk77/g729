`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePx42lvvBMlfJm8zQLpWxeacm5JwId13xOmv8E0+IyYc
ZJ04ptocAtmJkAvkiMlVKtRDHGEKhsTyVcrIfIvcklTuuSPR/DUBFz8tjvFl/BUq
OM3NLjAMyeLttt4S7EswGiRgh4bOrlKxTLCZmda5MZN9THcR+1PY0gEOMSC0Eee0
SZFInH86w071Flnxy0s+IZLeO19N0Q4jWkaYQAYPfZQtUS/f1zCBn19dIDuVF0uK
`protect END_PROTECTED
