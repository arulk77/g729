`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48Jf7DVNdMSNSWIXI3gM7rUgX2zdLa0MBOptOAF/R8b0
d9I17Bqxa2P8dVsaeIH3v76Q7dgB6Za7YRji/RH+LraSYPLibgsy38JDd83oC/NB
EsC1chNFd8ieMGZfIo9DLX/pcFGLLRX+xG4CkP4ABsq+SftzFIs42CchgrpOcqFv
vlktae5iItMSpGkgBKu0BgChwevGxcZjdIdtgaQ8NdUTv2g9DfpwZXrPYQ4Wwsjh
g1zBEUu2/4bkcLc9QiJshMij7MtmFdyyHtqRonh07bMKLhQfBaywHWtlfo14aJDV
x4JnKbpoLu9tL19xxGgMKFCGnymYPmma49qdGUSOkmIC9sgsnzC0JuHDMIy/Y4c8
COSK19rNGON26jQMjP/fwbLc+bgGsZrDoVuIiH65XtMStROq21XPKJeyCmckOjoQ
6m1SV9/8lY+iRQOzXkNRUA==
`protect END_PROTECTED
