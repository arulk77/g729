`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePxdIL8twwZclGgeJbPkmHJHGEDhsK7QUFElyN8QTUN9
qalvPNwWf0V8HMhK7UIebiWw5zeTXyBXC8qi68/LaX/jdF1B/x+H+4xfl7zypeKR
hCkkylO3HFtl+j8pMGuuO7ycHZcnclG5keBV47Sj4g63Z7fYseqwv8/kblSDq0VQ
+M9d+65nXqtzFEDXpQ4biin1WhsxiptOlsQJQB1tOWJCKO++yeSU8Zy71ZUZw5jj
`protect END_PROTECTED
