`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
SD6Ok1s29F08/c3sI3L8AUEdgrrvB1S1QzE9tMCPUgBLwlhzSHmaOkRjDrWGoO0w
JwF11Z2CdpZYijaORY2oWVWisiLv3LSG9/HPYFiY8lVHoNYtsIUNTvT2vPDqOlRY
uVOnDmqoLW7MeVFxlwDzNozNnBhiJXy3fIwyDIcFadw=
`protect END_PROTECTED
