`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xcD9uB0U8YYlI7BDU2y9iSl8HFvfTY8pTDZsDQwx6C2
PJ25qkkkaBViUHusXsmNVUybf+D7gqi83e1y7/oz7yUR7Dey6voSOX4u9R+E9nYi
LWnJdu9zCiMsTTQ8jc+mm7tQpoNo10rUIRS4Yd3YFh8WI9g511ffc4TnC2sFCfrt
oOw31RsVLPzL1WIl1vQVbdlgvNq1BM3jbyUnG2+Avlo=
`protect END_PROTECTED
