`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QYjNd15unvLKpC4Ff8J9upZHGeRMPyHWy+yy9fiZrNvIwbLj8ewLRbhnWyNsQj86
vqsvG5j9OKrhEFzilz8lBsXpbjEPoSAsO5grTkXLK4M+VnI3hFHDJNp2ex3vfhVZ
U69ywWxyDRO+YlY+wV3WyuIJKXvDpLlHnyDbwLE1Mk1Qv9kR9T6UhUkhzt8M9Rh1
NRCJcXMh71N95TxZJbGNTHMuCMzjni0s8xOzz3t6p1nzvTTIXNmMSAkNBCAp2jHc
V38A/s4L/VTm2vatF1hMvBM5nyxqsP9nWQnSCIoR5ciMydVKPyXCOAHnRgL/6BkK
mzBxcaTNQVTuqpO25KzfZiMT0/kOUxtM4yHPLMDqUQKDp1jQ8kdOwOd2fAYcqSHK
gS1jr5eD3i04HzN8RylKXy3rfRubtWOUbmuP5vRYR7ch+dlmob060T51dIktKjl/
9xDwDACFHXcNDAN42pVLuQKVyUZ3TTm4YcCakB7EVjbvADkhWGNmSKzRTOk7jtmK
CE/UJIYf4m/HUBtjiRPad0U1P5S6rm8nx86/Qy1Qh8+68VUZstkwqihFIUrIFIWF
ObeHIHfAfyzWPGoeqMdfZdnkttDmV+OH/zcfRgFfPoJYtrjawgo+e5JX7CUmTin3
qc5TrJYJXWfXtZgAWKnjkdVkAqpMtphzSiF6fZTOfFNNlRInAjGoe3EwKVDWHL0s
3H4UWfpahZqXvWMipxk4eq3hLUcN+StOblPfCfhGqEm7vXXG1Jg3yZEjoyomVRGZ
i05oWh/NDR8p2tCTfk6IczpJyqh/QV1Zx/blhjxN0w8=
`protect END_PROTECTED
