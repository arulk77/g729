`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aG2h5kRBNfXQktcrsDOicMYe+jOh2Hv0cV2JyryGA+Oz3Or35vd7J3j6Nwy+gaOg
tg1X9lH8Lx3UMuhvooy0qqghS4Grv2+IDDU01mrsA7hDrz8KpKQMi60P/CGK2e7x
GlAdfAx/aGBx7tzy6UGWkREhX4byCGyBO7UWmhBVdfpD75x6OORKYczShwIYbYvC
`protect END_PROTECTED
