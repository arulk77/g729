`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveE9hi0prARF/ATBrjKSVqeR606/B/aepN7pLmm7jHBY/
z1T8BgoeSzHaw4PZuQtzxgpyjV31vK7ySmK5KG5g3DEA3H0LekpbRf5PXZUE/cv/
ygVVCDodTdH2VhJY6ZR+xv9mZUq7U/073QxPupdDKFBsLND+21QykgnHYkFZIjnk
ObXX0QpXJH76vVZal0hKDgF+zzSyYRXrCKNBN5k+4K48BqDq7r2zxUM+/mGqQOWW
L77XdqAD49u3/VSYkNwSfn3PxidQHG2mqjRjEc9xhhYuy/TXUuxaWLhKgpGxGYmw
h0G0v/8LCXXKYoswB+3Cd4YdG3p8SndaOWIifXCBCW5Sm7+WUnsoeg8SNkbmcoVZ
`protect END_PROTECTED
