`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF3mIWB8UVozAbqrOyfRjQn9zknatKEbM5+MHde15XJe
37arMjOLFOnamAxlm6xtvq8f24Ef9Mo3ozog1mFFs3qKr2c4z89F+hJ1xLCZuR3b
5CwbCTF9zUuSYi5MmW6s4BELdT+JisbmgRcvG0t020vlQPWuAfOeXuimwOvR4SiK
dqHcCH4LmqNjctpgpJyHk6G/GbVORGgAR0G+y5RijI9GxmwlALmQ5wSwnpEBuFt8
rh9kqn3YsST49eux1MgFFsBMjF/I5scMZAZ4AxV6wu+w/mXu7/PyTXi/8fv7XhWC
hdFsbFTOVHXOqQuGIAlXZ3jq/jNHJjySEJLKA/IvGFZIEJKNDeK54HOeaRiOX1Na
fpDMEYr8WWS2wuxLlkhZSgg5V5VLIiW77NT0lKgp0wQczTzp9kT0bPHAvqnB5qY7
HTViuLn5pMZ/bIvlWXUB77K5PXyaAOz0SWptXOOce7zQKnkn+f/IiMmu9+vTO/uc
U3+dz0pjQcHaJhoCh9i2EYorz+Ul/z3kWsZz3+9aFXHwVghgLFYiotUFdcOtgPhj
`protect END_PROTECTED
