`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLQBYvv1XaMsDhRxwaVPgYJIWtOa8RvrzYf9bcxRWd+v
dE3D2c7DQe1vAX4gi8XCSrhiyPdqlVp0SGdOJh1Z9P39eTZBpHkLsmO0Q1KsXchA
MS0Vv/jRz9VHYepZ7hS4CKKbzEFljxKRPpqCeEc//fGXnPjsXv9UiM+mCGWm+XYy
pM6xIC8wcukLlGdKo81wiw==
`protect END_PROTECTED
