`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
BWFrwiuvB5avdsjPc2N56WPtEbl4Z/d2AsQ4iuX7PdS/Jy0BH/Pz2QNM5JjZBuOW
wET4E1FK2xo4SuWdFnJlvmRepLQo1g3RxsOhtXiefpQiMq+zU7A9W6FMNqyFXA7P
Hwy0JIiLMgBvY+rSQNlU8hAtIsMHpEWfDZ0XjoH8L4MDOT9M+Fbh36SCKkChYP/v
Jiz6fSO0R5M9vkfloKWS/246KUTtr/mvRZYsA4olrGuck+OnV4x2BmxQnbTzuUrh
1vS31cviIoRkrT+QPKGWi9rQIX3f0XrY1lDt6sl2t1auanFEc94uo4FK5XzNWxd+
NIPOcqdAkDMArc2QilGRM/PW72kW2oJ9dT1G9dLttlmLdOgAvF7vGmOFVERuDNAB
3UuHCFtE3HL7D4WdDREB++sACdSS1SZIxjjZvZwRtw+g0BhuieJFMuxRqgFxte6Z
ZnmV40KHyTyynbj7x9aM09Cl4/Ra4pz0/PoaHaEWBSmy+AWKZAAHpWMt1fi/xcRn
cmSVxmoxvhsUVhNtWBZcnHbYKKdx9umQFlinP/pYDotknBwucRbAbp+f+O27VTUO
yMnhWdKOPLlyOPN7c+1r4jqBos4mYv/Ve9a5RwNNRlBc3yvfk6eAJHj34BwjDZ/M
BAT8S/iOQwVOC/eZqrCuy14iCEH2I2oxiQSbARRmZw1vzibGDPxtqQ29NLE+rOUy
K3Vj6McC3eTl7H92jWCcutrNuMtzGnMN2TOjlNDOyqDY2hHWciPgVnoMTyA1sn7q
OFAnuYkQiPspbsTy70LPqmxbMzeg00t8dvMAmdpDF0IHMfLWH/7ZrMe/nyEzbnSd
2C7zly8i6hmSLm6yMmBBHR7AGFjf83kfN4AbMveOMcLI6bY6gfUraIz/ajQHfkUI
YuJIZB8Ncyj9RtNWhMZ28mNE9yPt424JwFBTxxD3Pw0=
`protect END_PROTECTED
