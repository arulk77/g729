`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47M5TnOxwhiJP67Rmf9ilYfTQHI9pDmOFqf7vwGMTJ9T
e3xRRYdTiLzpdLsK/AcAHNN/6OoBeXyb9WXv7BC1fUWKINHZi7OayWScr2wTUFHu
D1aTzR51cn3J4TEDeXndoCCnpIjeRwwqYNwSRIu5gzgF1Zu6uqip1dMO0zfmmSl8
PEaRSnT2cebFChKxZjMwbUBrZqkKYUKTS5MKzlC2S8CNgbAB7QLadXYg6v2dyUuY
oQ0/v3viaCV/FCkUdAdVyp0/Ufp4EMPLkcHzgXq949dtZT7+8+zL6m6eLQ5iKLKm
j+kLZYNTS4KEIeLidz/GHHAMj5YiisuwWNPxUtTt54lfXB2/jl1H0N+xI5dVt7Xz
50080kihtWo9SFICsdmTfw==
`protect END_PROTECTED
