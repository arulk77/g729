`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
VeT3PwTsA6xLWGx9az5o9IVx99TL/B5562zhFL74gsetGuFmjJ0F/xq4Z1JexVe3
Ym40r5sLF8w85zqKDcQ1KAxlapeWYWcFWIPa5GZLomEYpTt7mQMdEig+0cU5XBwZ
x/oadPn9Sxp0PUYCb09zzw8PrHW0zSjut21zHchXVDLqD+grPYp/PsTAnR2HDXMF
IZqfq5uybMtWJ7NmyVJiW3AfaJ9O7InJC+UbB0hdryBVqbeN8JQV6m0gJn32U3R8
n1pmqXQLtLaMNpkaq3OJo0uKqPTsw06vqnyorElC1SMu6tVyOTKHGanl/NAWDvFV
KTivJRgAnqgeiuCDVHb2BoVtsQIy4GyF5A0sLkv6SiwJwR1GOun/UmWN8CX6GlQS
eGUz0suQ9SATWb+ucQi3jLk1jpg4ha49rkmTbjXPu69lKqoTPjatexy4x9AkocKT
CmrxFlprSKIUx2gSPLUuQqezAFEUagx8LhhhqSmjFi+b8YtuOdAJq5YLWHzYt1Tk
8kT934IF4Dbk6SgXxBDq0Rk5IFfvZKenhOqko8jfUxur9dPnw2GWm1jgqgrH1bLe
XBqL9jWZSNlmZCjGlBB7WOHutf1dBYIcX8ynBwiSMa7I63GGEHfLB0Jak5eOk40J
5w9SFFyov3Ri8b05d2JQIiLsFHOckngOCYKGpa+HgYPC/t86Fxi6VlDhgG0HfHZq
4wMSsJRsrj2IYbslkexlEtAIqhWb5XRJsgNaDrRdFkKgl2i5nM+Ijy93KPsHi1Ux
B3crWcQaF+feODg4XEqpjkE0D+Nz8g9YkMWoMb9UaiJznVG8XXtuuESe2QS4TdDD
`protect END_PROTECTED
