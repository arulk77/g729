`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
X3qmBIkXW/S1CJ1RaSZbIvKyLyADWMJaEHZGVN5A757dSPF+HevMOcvTK/Mw2n6y
AkOwEQ2eh1+tgr80z/Bd9n0vj2m4b+WmWTFdAENntc6i1Wpjh84Spd7CYpzEyEly
YCiCRkJVhOwyvTi9IXR5mJe2xStWhvTZHne0O/bAwAjXzkz2fEd9SLAiI4zQ94r5
YBCwyeTrafoMPW+7nx/a2xyTHGyxjxJGp+Fp8qGRxhL1fc18/mFXcJeBiYjD++39
3AOLWi4kIUUe8xOA9C7kACxboH6QH+nkY3dsUutq6f4fB+31ZYxaB02xHUAghIIU
DamOWha0+MKVf2Mb5iiqUvtcDRQlYBPwlPrSmFVQQcgKW1zxzxHm9XAqMxvyF/I9
AzEhgzhYLXlKl+ZpN127RtajCKzY/06M+eFArVvirdLInTHk18Q9EgMFmgQ+Zc3k
0/4GfZ7b/qlj1VByUDAsWjoN+tokSns6WV/NVkWiWrl+EHK64cP7kTjda+8c6h66
Gz6Yrx/DJ6Ys63cJ3MTYxmus/DOxQVIBEvV3g7qJ64o3BQdU3PyQtlovJyB/Gtfp
q+8pQ0W2RVvYR+TOTAql3TrEkBZc6rWW4dbul89XMVxzY32i8JgEVor651xqtZPW
1GwD3suZo3Srxzy264ExyHNQqPRN06JGvH+oGoc95jByPKMQLa0iu9/BJV9E2Ghz
GSh9RvItAgpRpK8ZAHATXj876bcADOBTiHfivUuscgK20h5gc4THRX0V2SOMj6aD
56QxSPRSV2U+KRo5Y8Ud1qFozj8h4DzZS+qLM5/uGLZM4USNHWcV2YEm8znu9bRB
0J+5ZAwMm8+vTX6mkUNY0yIBtyWZ5OoCLrIpF/kYUXxBHfjJIMJEeKEwS7UUzUsM
aKEFJkwEf4Eb4EpO9dhOjK47hUo5JhgPKhLcsViUPOYCJ838MbWe9/R+ibJrLc2u
t3R67wve7S7gcAxrrFtxObP92R1+G8xHNurEaMUEK/JXb+ZDzcNJqC7Rd/EmccdB
JrE4QNhE0Ha0b0+W+DHMileC5wwd5WXW2ERzaga1+WZLdXodyVGJBRqRzWQtTVCI
4rqcuPqLGFTyzT8/ex83B6m2+juBtiaLZddlWhk+4b8qJGnry0E71eQVSMnDFKBn
nOMKG7nCv2eRGoWGKL61gYdDrb3/Uu92PoBeW9j4zJG/oyp7Komgl4Q0bwVxphUS
3Z/623PvmKpTupjk6SGWqszp/UzAJO0fpv+z+z30pXBqjeTord9OBhgJq+EY4n8b
ftkYEvQa2c0R+7w198H7Fyw339jXdXHN1kxPKtqBAPSbYazVB1X9S0cIPnoTWCJ8
8Hcvm3xHQ38CJaxVNJxtfG30ThoQa5Ppi4inQVPBNPUkHQuytfiHPCYdQckoI3Cl
jDOu8sXKTTVRZmQqmvx7goQabnyZFF396QxTglMUYRckEwZF7zRjKMWSNn7TAHA/
q21RwUnuELrtPSr17jSwtv5X/Xzv/gyazUNXti/jJSfiC2gSHvXeerSDLh17y+4m
i+Yd0RJI/CT+YdKBmL3yJa1822yqj4Xx/KVrjrbvNruPeuYLrStTwFPzuLL678fV
mjTuLCXEkqPLw/64hK7vbKGZ4miamZhlMtv4mHUTWrMSZNvwYdHNb2jaWf3eIcGJ
5oSCKrfTGztibo+JAFYaDM4f6t2Ig9J4N2/myk39BZCI9vZIWe7nJA1Dk4nJw3z9
IrhyPJeipZ6adYeOFiWudpy1UMc6JIKX/z4Mep1Ybu/BkGe/1uj90PXwJJQdtm8q
PZUN9UvVqZ0mfza+Pcgnc7mNUwKku5HSJTQ9UPhQfIo6INeT0AxB92zovOtHDtuk
8l/EFqCUmVZLU6xOXQLF7Lmgb6bWPhPLJInA0/KDCXSW6rmZXfa1Oxe3+JTiKc6x
gC4bijoGEc1wVcOWQWnMC1/pwRcJ8gMbZs+AkCxBXE+raRDybBXOGx4gByUV/j1o
3Ud6JlFHGk1EyC/r+ZmH63WMYmEWP/3/zslW4WaNmyt5tirp56wE25gXIiy+oZx0
GA+G8dBpZAsluHx8RrubELXVSggQ0Ez856ZaYpM6R15yBVlnZ7yHzgfPxc43ME98
B5gnaFqJCdrTHtIfAKnEvavqVtqoLRZLOI0iinWVWPOieaJsxd3mW3Ru4eimBknw
XOT+XSBKOXAQQ5FGT/J+hTJm07RytK/Kn9QUQndPrls6tgIMmVzOcdqlKMevpRWG
8RJrN5e7KbyMjdd0g4LxHK2wwNrmvvvC4arC900B5mKzHDkK6iNPJxM9qLyxxg1B
n0sbrQGFI6JE8gWedzGeIbXM+lmkrhxEL3Lqe/dc+h6dDc4HFPToudRz4qi9sucY
Xenr8aELkwQ9vkYamHQrI6Sz5jZsqrT86eTzhU6zQRRJByjwnJssplKidhrgtRtd
AKaVK444+3xPM71uuU6Csam5k/TeuFk1i/87LHux/7HSmz+PupK9/7looKiZ5DpG
XmE+7SiqRi86vQJE/YFxW00szGhalBO9wQjiA791ol3seD9RnHFwHByi99M5SM0V
NsJaNkN0VVtnhuAz9xqE2eIz1A9DPD3uFVw3Zriqq615mgN5lhKh8Rdk9ffZ3dUn
EVkYRiTJKApidTi15KKFH1YcUbXqzrqcApcS5X+J1Yoh9WyrPUtY3WUz7f9Nmwky
e2KZ5jg+/4JOLvrIrHSgmZ/yQ7hUd2J7XMHFUaP2YBEvwi48TPOqhPsPEnd0M+8s
y3Nv1d6qpDv9cLLCNXxGf6edOcTxXWl8Ad/dFaKAOsPgqJD/iUeLVQzcc4SPS7pI
o74ZNYL14t7VQ6B57eobpUZTlFRk4H3OHvaGTNGGl2P0ODvPdMtfowgq+XabtJjB
RuudkdIYrsilIKbtwjafGxljXchy9welwJdbNX4iGo+uheXShCzEpCk/IuT4JSDT
HXQRrjSC2zJfpbGWp4+9eDdP7D1msixfTfDE0sbiCJXEtW7LQYCoWGZAmsxsYmJq
9V67wRsRcq/K821Pgi0qZsKI/xwAnPHXJxoW3b9l60ZGqW5P/0Y8ASiJ9DtJ31w8
UBUl3mahfUsXHR/uLQn3ddDwE0cUtVIULasn8P/8N229XWSJkQiFrm22LAyiFxCh
BgAdhMjU06EuzlBTmlnpozJfRBy/ax7L9u3a238Vw8byXtfHIGEoacmupIEwRSpW
SpzlJ10ah/rHv5z7Z9agoa2hcl86vQe71E78+bTdoDEuOCa6dpcPfyD2fymjOU0R
I7/ETA+yE+p+wDOi8v69RQ==
`protect END_PROTECTED
