`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mlFBzCyNIVABC0bhYTMiK2vsW3WPEY5A+mLZq7i8J4+z1uzvuHjlIFBw+EfOz7Hv
5MFbuyWvvuRUNsec0RWFSjyARiXhimD24a1GIWAmrj+NDGogopRjv93UailqzhfW
zedIwIvAEBYRqeYW8+nOR/7RvPv8RYbCTaKktJC99U2EgLWHimrxjMoOE5SZ9UaT
Rn+DWNBsA/LXpVh1+cej+g==
`protect END_PROTECTED
