`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aXlxJ20TBptpseTnyb2/VYPDnVo1sjQY0mbTf76orGs0
vkTEx1Q2o1gJxFLyH1rAJrPN9+TyZ10HSHAMkYQ++5Qtu6q7GQ54xt9gaIypj5p0
qd8IWxLQvloP45xb4D7tai971o5cjv1yEN7FTvfYObdtV9Lh23yyH2R82W0wcDQD
9dlTcK4gvGRZ8yp9WmEA1ggdxJ4MJmfU15MKL/sOQjmEXeph7aGZfwZS/qhWh1+V
rQvQN3ei3z9HK0UbVlN53iaukdshYaaibrAADeTAdFTWMT6wR6uidUcJEOyjxNEQ
3S+rrTb55YF+7+dLjl2mm54S9MCca/w+VzkfpTsnPT3Glu/0DPO/BY8QvszQ7eOp
nI6Zn39Bt5+2t1/PC05Ov5co1bP28S+P3jYr/gMuoxI/sDO6qB/uzfa3cCKXsQhW
TzJV9psCLmyrIXEluDBzgtBJEfcVTWJpjRseanDU+cn4006DZfiqmNJtGYdyeaRL
88LJZhjK05tDb1NFZ1E+tztIy1qDSqMOZo5mmwpRt5SXk0gYR5b1A4Au8K+aazGA
GyaIUsGIP+Z2gbB0z5uBQ41qsEFgtUP/avWCDIUTRRwrI194CXl1p7MEZ4rc5TRr
2smOdJTC22KBzT6hu9bK9bIovIPPiuSucTFgkfex9TI3a+h3sA+5zp9D6kmtZc1t
u2We0bQxcqYQc2rKp8L81207nA16K8T2vKJ+JUVlNHhNUYTneHsVD4VBfKWOOO1c
RGZUHX6fwXcJBBY65csYPKLGoYvXHYlsYFJ6W6wq4WzgdASw7SD8RsPdOl0juNY6
CF0GLFpUsOGk6ldthfmrHg//HfhApOVPbCqkuemnJ7NKcGhX1J6+BZHbAcs+O6PN
PNipviXviJlWdz+GyAV3B3ImZ8ye9pKtDlsn0qD7tTqjCq4TkfdCAdsebnc/XuZ2
bL8oBoaA2lFfzwDkOHcIpCYzeEURZEoT5RviI3u5CuVNp49Jw0+gtrFeeA09HlRx
jdSLOeZTxOKQ+E/Yd/vjPE1wjfPIg2zfZ4xowpZmhyFhWBtj2jwg5vehJ2r5JHWD
O0weJRBLrDWCeBHAo6g7uNjTFY8OcIcNVhUc+u7dEcFLwp/10jgO6iM9upEVNLq/
WDsRvnlNoJGjaXN6Y5rXFD5IReHZpuF+TOdFXeeXweDAbOYR1Y9ROPxqAV+M+R4m
b+9IZ625GxxLmQZKf7ptq+iD7Zbch6uvaRMzsucCSfG4dCjJjGYmRXxx5woU36/E
wlH6A1Fd48Gr++tK/xHzYWPzpYA47Ri84Q2i35p/xrG5rm+HQCUlUwO1P+hYGiPz
NvMCwbpB0+2jakg0k2aWR7XyISN3NWF87eVGXoObaC8BOBKXPHcsGYyvTSo5pt5A
F4q9hC9LJPwyUyODKX4vwepZgA/dRe3iY7UEXUW88ix+83lSfo85vRttRumzx/UP
MsunYxwR8IaFyqqtcX9JIWAXkMZsBhAMJlEM4U3aq1n0F9/3Q0hX9mg/P5ORiV76
mhXhXO5o9pQa71iXoO/aNP8DBz39V0yRNxO1jZnqIEVuWPTPU/hg1fNoEgNUEeFQ
zmbS9Y/7loUu5s6N8qikskxQXIdvQYFcuFxXVaVkU/d8Lpv48dr+6+5VS/XeTdp3
FxTV7PXrnJ67beuR5jTWtkbFRfio9uvWQdLBAxcqZ6VDIT4JCgmxlOxOMex+5IsK
yqAIh+6mJ4RQ3wKQ5v354AGDKVAkpy2x9lIkqXjOPREdbUJcrljSpLY6nVJ6R8xS
rY4qStP5/hLlwOANGrayaY2oNHR0v0VZhAlYPn+UIf7d5qvTsGdLC0qp6Ow9zROA
0fRRSLN6IeFaJPrl7BKtOBiSJiLGBscLFwE3dXAsLZzj72ZeoTGqlqZHnTs4J5qa
pTUEDivARf+ycH1vjJon2vPNYDHsHabD3Krq0wD2vFdvLaXnA7BArKYiDN/2ERld
Aw3Lg3X23GDxcjuJLtYW+SWuVPQrZfyrgvqcMbrVSoaJDljustWtoBZdLrvbuFKW
7ritWCEK0A0yKKjN3ysfsD9Peyfyz9WPk+JTSZ+VpEE=
`protect END_PROTECTED
