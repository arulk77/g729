`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL855lengHhL+9xgXZ8Pkhmcak85la+CWdt0I1zaw20ZTk
x8/WRNPTLsrXdz2ze25V7sOL0EWv/G+bZwBV0DcB4zLFgiBTMtCNcJZbH4r2ZlU7
k4Onj9fTmnpWA13idl64Y5QGv94jR3kvZTEXQx8k+w2Amkg8TGrsgysMaZxVwnlL
mqDGEhTHggiw7YuziZTSxRtcsPN73e/7mnnNsycwAbwZacVKOuEdXA+ZaTw2YzQs
/9hPDy+yt5TCIyqB45pzeYawMwhfctlhsq4gN3MSD7jayPshHW7kA2gi18KRplZK
HXTPit7F2v6EM57mSlD4Mg==
`protect END_PROTECTED
