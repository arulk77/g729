`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveClRvVnBMHdyranqCcFo/XLJWNCvYmw179QtucdQHMmc
RUBhFFHmpudVeFcGZEsAK7yJlKpyNFQxiD43zCOE1i0e9aiXrD9wg+jGahVgs29s
+k/+RUPEbRNVX+2+jTbNiohQJivVrmSpH+USW7NqwFXO+SxbJPQxXRvpBqDXvs26
g5GUSJse2rXzKbJCsnfQMIj6xyo8e1tXGZs9VengotXmpPocJpYkWyPJKvZ6ejrs
VpBdP8RUb2rueReDalAvBuxRP9JV0s04GYNJq5m3V/rfgHkd2J34GvP/uzYVaRpd
VLCW/S9nUGsnXTGgZ8XfSlqi63Y2g1H0XPKdZHQ9vYQw+l7pRpG9FITBiHT6Ra/S
e6GXq27A3KjTv76bBwFwu4ZHme9V/6sYfXAn9BK19y6uBH0O4X32tZwTFtHWOmht
GxZogB9uP9mnrtN2yV9GLA==
`protect END_PROTECTED
