`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
yy7YfcErnaHAV5XOHXVfo84Tt3ruW3Txh4cMxHJF14v8QL0JzJ0Db3zcKASnTh0C
o7c5zwx8F32FhE8238AYVGJGAqa583L8gulbIG6cDMilI7W8Ar0zZqwsiMfI+aqr
NwhdqTpKBIUXSuZe2yTxfQKqCyZv6NUcE5abmo6tpG39ZUhKTMBHNn0Nxxq9EbOX
TSuQbj6TadDneQSSOqDnug90JoC/OQ5EyjaCB53t/8I0kHOfCGTLiW1Uj1IwmUTC
g+qe94zV/n7YUnHkpeoGn1HMM06OsqH9XtDvjVu/KUY=
`protect END_PROTECTED
