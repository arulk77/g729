`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
SfmFpXuhToiLQYIoY5KO1CydeBbv5n/nLjNv6Nmxyd0jKDOsHgvaW6SY+UelrnxW
RCpdDx2jEv654XifaeOiUV4x9HIWMSGiICI+shMXvefntv5GWNdma07K+xQfexnY
5a+rVZ8738njFERXk/q8+SZRaDFpI8tOKhs2oQ6y3rgmW/ZIt6YDKnLd42bogYJq
91HmOumaUd/FWWaJbCt6IeKUT9ZNTDfH7AtZsCIPHHE=
`protect END_PROTECTED
