`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
6rvgfgIm1zzNVCOyFmzBgEdivosU58G7Q9n2+uWc23tmFP6KNQVbYjC6fzUrTyE2
47kWC+0RVdmtQcyfY82wjQ1BvIiuicTx6u6klJGLHVVzmtpT64AeLIaIbdnBAWs8
1h0s6L258IOJTLJ9xA3pDxaCGjDsVY/MWQEerHy1pEYOoKqBltU0uLUH5JM+c5g6
IsxWpCJjmRe6Y8vgB6zBTHEEWTsEuQDgOUvAHD5Pxz978ofqpXg4EOxKndR3nZuP
Lq+7IawjmidSIDrXewncHI9dpg+njeRxN2M4YHS1S8xH5Ag/odTxRfbWgb8SDWo1
YHegFtLpUTbY57r3mnPj2oJiwacIB7xIjxrytP+HnHc=
`protect END_PROTECTED
