`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48MmG6JWEreRnNfCUP7IJjDsBePROIoHl065L/il6WuG
7LFPl8nJWd5qLK6Bq/ErjweePWbPQzvQ8u+XSouC3rD7gjHgVoUA4x5QM8hgzm9A
Bwkw9dLGjzawu83xixo/4QMVIe/w1lL+ENswKT4LeqC3h9Ta36DYvkoecTY/DBTw
yTbmORJyqoK9ynaNp5h7XOEHTI3mXRwqH80WB3a44XrzPS8xjCMswZYPU0CLFW/r
P0uvYmpHQ0GHe4wsOdc8p3FnaF+doCU+RLz2P+LwDo3i0gsUxTzdgD70aMEFc3lX
dHM8IUhz/r7QbmybPXrDgw==
`protect END_PROTECTED
