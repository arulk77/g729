`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL5fTeMmAimJW3XtGsgPJ9k+jSeEKAa0egD7iLyEvniy
nll45tR9254oi8CSKIJhFKoeL3PmOzg2mdote1yDyDV4uRZWzkJRxd6A5hxPTlun
1HpyLEza9zD3vdHdIvghNuuQRCd/7z/+gl/BnC9S7czxQf7gkPlVrQEyHAKQkjxu
kp8v5blje4O2jS2VoY1zNT82RX4RXGNK/wP7/punnYb9OK0OF3JPUQH2ciDUXGS1
e2w3ksxcUxz7BNUQQmGtxGL3IUcAmASybmGDcm7yujDeAWw0RGZodbPBostLCjgb
dhE+10fjYyRFUhJQC/oxKgl8zq0vQJ3yP5xkG40mwByKZCOAI3wppYp0Brznp603
yZpzZ1jHobiZZY1joxSLCg==
`protect END_PROTECTED
