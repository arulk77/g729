`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pnyY3jxGyCgnwWklYcFi/ePv4eDyU6SyTU/Evcq8vTIC+xDBrY1TaHFAAuPe7fH6
DUKxxKF+h/p2B7+lSGzdHs/dooYcsqWyCcBw939Eb2xr5CZe8GOx6HVAwQrw4Uge
CHIKMSckNX4Lga/6jepkVXT73J6/5rv2IEF3xjLHDJ42OmxX1cQTBRmDVjmNvfzF
ZKhKl8sjFWJvHxwGw/2kbK69nIWms/k+L4ErigsdJTQvj8lgj+h+3r5LYph98KO3
s5tE7JsH5X1XmbCPSuC9oeJ5Z9BIAEjZC1l2z6xJQQTHu7FAQG4GbKBGoihLNjO6
E8WFaxepWOh9Sf2OJ4rtJFupHDCM9MoagfJKFC7JqgCQCB2oTgUy7ctmGP/7jqyD
`protect END_PROTECTED
