`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu438sq+njXyTdWBCpGUPNTxem9flPEz3vvtMr/X9Ni0+G
Nl12WowTYDJmmbFa5XgpeWDvX0ySfcxtnKX0rtEEoVD69LQZU3lk/kicPuco/Ziw
UHZkwoaRwqLaCGev2mVWqtlMvneUBdqKY2KvC7CcwEjUk8UHCPHhDQdG85NzQbPP
j6KFgg+zqKM7+0gd87h8H543ev83SiMRrzTaqoNYKjxOtjSWPqnHp48U00/NB6TM
kAMcsp8nNAvhocJHYl+nlz8FgiHBRTW3v2y6TJljsPgyooBeP1o9zW0C2/N1aYYW
a/JoRInqK9oFRsrIP0WjNjMgQQZeGcMci7cljl/iYK+I7FC/IP6wJUSHx+hw1sQU
Vb54CDJT0BImJtvLqY66tQ==
`protect END_PROTECTED
