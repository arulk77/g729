`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/wan6Sly2iePBCo4/mKr6mPeLiEPfGfS5j5ONV9RlV4
dGH1sGNTVYQnPmBH+3S9/MW+5s6d7bgBloQKDs/4mDXtpWbEaj16UvNsbIlD0WJK
6xOD9d+pFAkDtjAA6Didu4uuKdzBoZkPn+41ckCdtj8RMr8lXK/xxCisUm9Tv7ba
ARP01RDmAlYLYcU/AlRsibnMqhdzckszIb+T6sBXFIU=
`protect END_PROTECTED
