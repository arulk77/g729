`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAsKtCY7lxS9kMychPa3QRGae8RpC07VGTxAZM3bjjss
t24o+o3a1W/Gbkg/jivrwFwz8uy84obI4kH46EM+NXbsL+G+dwQSezycXJz2nt8V
R4aDElP4ujx4K/FM+TENSmcN8BVNrF1bz7+UrvcxZFD+qk2gq7YlM5oqVGv+vsOa
7+GXLPche/tCq6DS6RtCx/jXFIqSXhnoVRro3FtCN2uvO+kHfFGSeBKqCQMKZqMG
QvZBYD92a0Ke29wTGiZ5T2ne1XRZwY/dcqMLdQRQZZSR6HSTpLbKY6QpNup6wLW2
aQgyaknRt9Y41PPAT9duXQ==
`protect END_PROTECTED
