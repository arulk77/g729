`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
whfZdEhQhIVICrvn0VMg7lP/B64Y/8NSHoksUME8jgdPhjYmh9Ij5wFDxvkS5Mv+
Bp1FnkHnG4VTTr3d40G4jLVfqVA/dTMN3F0/4PQumqOTht2m4aYpFeed8bVHp8yL
IGjQOk4bmRMh9uFQEcHFWOqhMRBhsnVqhcCXxltKWr52gyjOXX/0oP14WkvARfgc
pnCXpXFncQGemupWjkQrWSvpjt7zOdNAbtgliQuJVicIrEsSnIwuR++0a5kpddsr
duX3n9dGqlYLxc93DAC8gtI9pPqUmTtlZ4tm9xB/ubdjBU+TMUxst2iDlnGMUXi7
`protect END_PROTECTED
