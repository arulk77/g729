`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C1HFaUpJH6+tYprmoy2JYPe6jJUbgOemgQ1Tyf+dtoJg
YcO6f16ndWX1oMHQiyf+B5hgt+QCInnUmbYsOZe7w6E6NmHEZoIaFFQ2hbNMe21Z
HN9Bcw95Rh3+HKPyaZIknodYnO/dwh9QbkCOVkRFFGHYY42+3VdfNN/Cp6xInkmr
c2HGbHbdWj0A+PE7dHFVoMCUVRl0T7UYFbAioTHylWIFsh/XXmAi/Ywieg43sqYj
vXrICVP5zVdRIxioEIg41o6WDCLsXFtXx1p1vMX6hnUhmyRVJzeMSXoqKymHGYN4
CoVX8THeATrj+70O+ZzAwuNiW2YHiOvdPqbdtWoRb77aFYSdamkLF1fuZVfUVEAh
hwd3Lzsh9+IVYPXdeI3rsmiD7wak7E7j0fNZoLkv3gyMTRH4RVGj7fnWRafWTC/h
jBZqWBC9mL1WvKVySOEZnZ2eFcYLZ5VRPn0mSxLUr8KNBTnLje09vx1xIaxQkM4a
ETo0ErHBtcsID3QdGbSPj+CGDXJzwiOExbojKyIHE6qjHU66wZsDnByGy1u65XUF
p4XGt0MangwdmrilKCHxGGP7kNaNU5m8PznBUnYZItgZXVT/oN7GPj2/iOb9y1hu
x3jrZc67tHt/4vxs6gic87lA51MkPrxAh7L15pLgGbds9OCTdcAHo1cYCBJMCiCw
YCFVTDaL5mBEwbMV5Em8flvi35aNwnlLwkhj3mZwq+qI6lBAuMIWUjTuwKtrlNLq
uz2n9dWnwtXE87ko22pBa7+Tx7JEvDs8bC1UiOIQIG2yuFFFRbFzxs0nAXrSn8A/
rfTFDSAvKOMEwf4sAb4Hcg==
`protect END_PROTECTED
