`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46S7nEtR4NUFwlzRHdGeUZNmNlh6cceL4Q3GziWLrsoQ
MaX1c+cpRNtf7NSXLjh8u2X3+ikrYnnplPwmZw5l51TnItREHVC8vzSOfa6RJplY
E20mEvBa5ghKhAFQvlq2ubYjeJxtb1/iYxNeJFNDmOI=
`protect END_PROTECTED
