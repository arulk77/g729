`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49+E40FvSrmkH4MYrXCcQB3zOtD8cQfCh0dSPD8AgKV0
QbQi2Dej/sEKXLRhwBwZ2UfgAYLE+CGt9Ca8qCF5KjfSh0IOjIVDodPV15f5Efl2
ycuN+fGR0XdZ6VLARCNt3FZ59TWZM950++HkorOis8FmTd3QmC11yrkb54TI5NeW
AOlB/KuxkNFotlqbtyNg8hBTIf8bFRwKZp8W3Vs9KNZAGD9EiKiRBIDnEuMZkpgL
E+l7vd+PxouIw9bfly9QOpjtsHI9qGlnG53FZZhdaJzJnZr/q1VDUXwNY/rUZS64
zraNNjWigQjRqSsRRWXCFpE37xDMPanM99O28/zBtt3WiXzwsPxLmzNQzrKD44Hc
6JgFu5McLNs6qHqaBBCd+A==
`protect END_PROTECTED
