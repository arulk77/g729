`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49wbK/wQDivNDU4EgBtr56ynWx+OowWVEsD47gA0ICEV
OzH12uhz9I9Rm0yb/YDyXKGxiKAbLtn4Hph7I/63EkhYVUsDKINy28G3x8r3SA03
iTRkkpn7z9Kt3wtnIPzsZk8pColBSamqD5VAMa1vgWzwcYeX9o/ZlNhB+Gz7fQTU
RSiiA+JP2y1+ArEXHuHf0ILTN/GHTddvheJq1XsL2Q5V1rmoOZ/2UPxpp50EoYyq
p2MmNu3TyH627nf0XNU7cSHaFYB6tR2Bu13yFjMYsnvUm/t/6fYWUZyHKkx3dIB0
rg08F/BJy7zKMtGzyQ02t0hjuvXBvNqIbF5l5SQicB0vdsN3YrvkssuS8ftj978F
rnu3Wmt+zdzCgcoCZonuUg==
`protect END_PROTECTED
