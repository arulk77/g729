`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47bpSjcuB10BFHecSSrwy2ENLj4doFdXSmyKO6wwaVZT
o8KWiHc5dj5P7/9eKm6eXx3EoB8kRMOroZSdZVWDZTAsGl5eRxp3SoHmha/e7YK1
XOpC2mQIlgUe6EtL4LriYqd3PxaD0P7Dted5VJD5rH8tOAGORtAG294xEf2PLUwJ
USk2OHa+QxaaS+Aj9QMw69XNoSxR0dU2smPZe73jeuLItWPxAuHZGE4e7/11TJax
o7bC2j82AI7RwJ82UDEc6y2SO5znUGHou9NlrKyvSVo/N/JUwISTqoDEVNLnP9G3
DHYq0BpFn+WEZWmiw/nOnA==
`protect END_PROTECTED
