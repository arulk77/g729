`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDdP1x8SiF1rBg3PR0B9KbrPpuKJq8PTqYRF1et3tzBv
6PGGpUGgjogaMsQPxD8RKLalkxwMW4JHYbiPum/SHjdSzzas2GXGyFcpyHK7AEiz
2dwXSqNxV0Hzmub46r+LM9v2KI4q35n8pWIPudta75k1h8yCyBRb/NS1El/uB7+w
x1T3zexOZfYApmJkFjOcuBrf0W/r+sCxctQ5yl8FCXLERNJwKF5hlENcCri5BWGM
DH7xJzQb9xLpnuy96ktl/jwryubYiRk4ASrd1o3WAdMYAQGxWUV/JBZ18nc4rBoj
H93FC3zYdMhtCfUoGPNcsXEVNBo+spNOgjsnt4CTitFTGKomYB89UtWLzrJDKpDg
hQIn5OkewaZOqFivTWfwnvj77RIqJXQEHagj9dHTPb9Dbek1xhqsK0iNfuaGFqO/
0zokHRzwSSCVbeogfyRFEELxA2eKmwpiaigAsCvkfVOwxL+CEDUsg2fZ+dSCClhn
fCZQGP8YW4Y729/CCUh6rr7DpPqDq8f0w4EmHAAFv+at0jS0EeyPv9yUcEqemsQb
`protect END_PROTECTED
