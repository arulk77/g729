`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLgOcrzb+6D/Q72PjG3OKQy2zJPYxyFog9cGUUMENVS7
two965nBke6K6fvbTictIVXGpTGWHJ8pXb46N7pRpgI7btrQxdFwbe9W5DfEgM7V
24sDl5chg2jJ1+qmJFELEhv2Q/NzV2c2IznEMphVSALL1t10rmxPjC236bO4dkiN
bHKTVzow8kAxdMXcHV6NGA==
`protect END_PROTECTED
