`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNThvkDGmPwuyz5lyshM+suOhH7vHwJZ5m/feWLX83OQ
Wpm+IuOYuZq8N+W7bn9NtNzjwSn564AQgQD5SzEnyyrPQ75NYQQXlSCMWxsT2lie
ONodfKMIxnDd4tLbe5QAmsIZEGKOTwHjORW9w3qAoP7+CQ8QNxRM0cfKPnI1Jqdb
RrVWlIsBjVFk76G4lthv14YGLmIMgoyCRL2ngDZBLeEmjt/cv+BSH3segM9aHQHb
`protect END_PROTECTED
