`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLSNqy6v+MGpWomy+UXIigrCDPplAd3WRxijJi4vnBXv
ubXbailTzzvaUj0Rjk2akf2ZFyg3bQv7Dgwl1dhHQTq7EzZwGc15i49ClUOIshFO
mYgPKmGlDxo2ZNo2mLWWi624V3uQGJikn5I/yCuO0DRuIPp3uHexwIsH3OGBQgeE
9pGZn5sK7M5KOf23CeTX4ZB2cE/zjqesX4+ld4WN+qhmn9cfnV87NA4KVjNPIm5Z
`protect END_PROTECTED
