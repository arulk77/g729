`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48NUiaiCHQ3gKT0xRP6mHJvv6c6CNO1/uXo8LfXCbli1
s7rc3eEHC3k7m/UVXaVUwH396ZAtyd3XTPiHqYyfulaAduz1oxMv32eLtpugk/NL
6ii5PZi6sWBb8CMP1y7lrrDrVWdKSud/d9+sxBI9Wd7jkDAi1GKCfRlu5ABAFcY7
MCD1vrZh05DNA0X+yR5/u+YC2nl0iPe6fat1YwmMN5D+tG5bPINjae1Dvv/rnC+o
b0kAba4vOLCuYRWGHuCFy0MuU++oST6Lduzjnf/Jst4JhT2PuO5X3EUgNUaHCEOI
11GLAGJM6McMIG5BQgdckg==
`protect END_PROTECTED
