`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43H2AS5YyoanmrUIe5//1BQmpiY7JM9wJQjbqAXd/PIJ
9btLmCn1+/s/qheIhmpirHS3lAcZYZTYQYYFvM2LR1Ux19xkYrsMqvV1wif8hraa
5eF1EFIRZvxcCbygPkb5Js3k6+9qRjdq23oMTcPDAcwJYvqf1UWb9/MfOyaP/7uk
JjL8a4ppmyrF8DGwaiNe2P91yNMgx1LewiuYUJa1z1mwuzAoP67BlD0Bd/100/Eg
ykFRWnNNIuJvpdauBMxSmoMD9KGQu4VWi4likBXz9g+xClQLuK4CRXV4OeUq+xN9
LRDrd1OJGpai/A6Cn2NobQ==
`protect END_PROTECTED
