`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
idpyHPIYi8+KZsU3r+08BD8pzeEC2e4BEGRKXDtbOoCH+5/k+05h4BcZ0+lSJ5u8
eP3OjsSkr5XUBMWN0/8t52+zqFF06CId51+YDibW/KIG8cqlljZB5srZAJMRz4vh
9iB9btf1ihN8XWHkJwEa79tnoU8GeprrLdr5T5/UlFfVx1V2gxvvpmzWc4LVynAK
i4KNL/o3me2W6buoPjkOGsJ6/BmiRGxWq7p0eHIwHSoA57EztEdklZSRKJ8j6DV/
9535TGFJYLCOsyCC/+27rP02f8L9xwASc0iFxkz3HBJv7Uo/UuxljaEJJVewkoCa
adeQdN8qWH7teRu19K6dTYpZSy4GqifZ3amo5HIgDcqib3vJt8cUJozsDn7QLH5K
972QtanGH8Rwyvcu5hW47o9gCvboOgGj/pkSVunyfVQRAONAKvSHHD6NmQLu+Wvl
eN/MuoiF2AKeZ2b2dgdVV6PqWfn82tNwIOI4RFUuRSy1QjxieL8uHOATBhiLhb0S
lcjnBW/RMblKnvjmI4aFXsmVDdETUwS2d22nHhegvpcWFBlirN0eWShMUlJD+i68
vpuy2iqIMOrW09kuG/Q2gmCnJUj+8JLm8p7/Zy+tRBkWX9byRC29wd4DGHgcM3nY
GGt7eabcLx1jW0tS+ze8H+3V5KwW8n51d9IMsS+2kWdf+rlX5gvGe9dgNb+38i8t
6WLdkaA64t858NYtKQRmUK5LfxvrZZ42+2kWtaF4Qq7pNzD1QG6Ux+KzxTkZpYua
yjUIeOzAad2WBzeSMiVFsZLS1X/06d6sj0bFM4XiKfAQQSbXUhZ5VJQzhwLyOvUY
PXm8VbaVgQj0GAoIQ5HPbkc8Opt6N3mlsK/7DuRWNdS6q5f9pARW8e/q7UpmlrDM
1Un5gzlmsR9AW2F6m0HtKIKXirwXN+r3AWlFVBHwEt8WKLdJyV5Gazc4dQzfB4Z0
NhEaW0bF0QqzJz2d6nLRryEfo+3PZ5EmtP0RCQXq8hOXHg3lcrkqYsT6euslrCVI
fri3RRXSIMI0Ub0ePzEc2TvCiRdYB0xucpgxNa5LYi7sYuqNErOQYCKTtuRA2owA
O6eNrs7xSwGkCayQ8XA7gEoj9+Fv9ZH5scVkMqJKeEcJ5MIpJGlGSKtXPEwzAWk7
E4pJ0bu73dodLiYy8ow2MEWbu9vd+Al8DlOrzZmgnQqxWL5D1oWmNLsYEky47du7
lBK6Y/fU2bQO8t0LSHIlbgkJ5koMswI0H+rDqZH0tX9P4jvzr5xFdpjkJ/Xg+wkF
8bzLamypQrMyUZgd1S680cD/h+TdMvfFMQEzge7FDz254lNRwnbrBi76dfzeGvJx
/lAJEE+ZJloYF6p54PVXyqx5xVuhsQ4cx3q8FjC/1LE2re5l28GHhjtKjtITgHqU
JYNNFu/7WbWyhMHz/i3IepyKWWVBwRJTdWoOOZxkRDDLjrDV/NC+6Z53+o/7dR1e
lcRYf1eshsXaQEgd5Kp0l3d9FrwtpsAoi6W4EGqcHJKgQsihpr1PJt8KTnsPAukl
u0WYvGnDIfv6/B8/YoDfK4SpswdwAjVsqjn07EnUIvXEiejcxyPyFf7e6bDTCZaT
7gN8rwaIXqM7aNkLY0IDbcIVIqh5mgywHtyOKawWVnm16TlQOWzifhh6Gq7Qu7TP
z3DHofRZXOOEuKLYsZWuZ9d4ajseD4bWvcgtbV2dnvVHv8+tokpDQ6EXg6Vy3eff
BpqdWLhNWeIYT41MAQAHgzPX1LV0jfXnbxmD9dxKlmrz0DWTNszG8MYTdrKvcfpl
zCftoMxbCt4wn2wkTLMEVDaKexQH1ye1ZTLZSxIyxXw=
`protect END_PROTECTED
