`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGYMXacCz+vfjeC3RTuYl7yn4KRJ0By65I8Od3WIP2Bx
Rspj7a+TTuGkMygcjx+d0vNvI9dUr4yFbAI5CKwYZSMcgcFEZR5x1x6IEv8s/scV
KpTmlH221Lc6vDyFehhzHVXaKcpU1MuxILHOjrXFWim9d50WEB3S/5mlGeuSrD66
shGsC+hRi6goMtlsOcQz/o6wShdwvR3dE1ubaRHbU/8oHktNcaBn3H6F2zdFTjpD
h5c5vhCkvS7gJC4I33Fqf1WfRkER2tXb1tY008hm+vDEveux5VaT+BY0y6bouiSy
4OFBe16RJtna/FOL43SWeob6ZhR3JmAEchk3X+aSUxKnWgvyZA/otoa91iKClhRX
/mumrqA0zAxhfN31Bb6GLbQHdM5NVNevd2LybSogO359jSMLcrDHAON24uM4WPRF
5RITzm8cITl52yp2CNLRIJZdMwhRjlvmpx8mtegbt1GIgkGQqbPeqNP2f3Zw5M2B
gvFxTjWuilBOFA0D67veps0wn1K6rvxkvL/DYct5zEw7e0G+ItamyxaYAtWoXLro
`protect END_PROTECTED
