`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ySuT3C5boxbK7UCqHwT5dm9dxXIuremDgZfuODH7dOYMCGeQQJoxjcUYxkN3A6Hm
6K2hGdTgbPaeHNSPZIemdg4kxjwbfnfQIbL0eMVkMxj135NziuOGJ38EsS4sNNP5
kdM05PUQe8VT5m+K58MvPItRyuW4U8xn0AoYbwMpd9CKiRYEy9VjSULVEz/2QVOn
DwrxnEdPDIvWlCRlr+8T9hBvZygUrk5sSgV5bIDfpF3LIh0EqE9hUhk6A7gs3n7L
`protect END_PROTECTED
