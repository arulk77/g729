`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNH71diV59tfZip3ILGeq0g4Gg6g3fzuofjBLwhrbeGX
aeJTXfuTkKBQzs/0heP0ZNCCMMG4cR90bQmrnaPLbsIBA759ksQ0Ul02W9BlBMVe
sci5TXuylTbFqlcxCBX+3zSil4j4u89VlPdqqwGslldm8VE5y4jxpDRzLChzqLcf
aRdXeFoM/hWHGah+TCyIbfKyZRr9W5oGkW7fbqHRY5lOWWIOB+kPudujiTM8NGHI
`protect END_PROTECTED
