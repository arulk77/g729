`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBVTxtClSinYuSnVaPWF/B9U8Ov2IbRYFtVwyCb7Y5Gm
ggXOVQL3d3PcMtE6W/TO61jPGwBmPKGzrXKEl1cj7knb5b3KOoNpjFKIaXqgZ4v5
IKNGrSL1ONHtfYxB+DXQGdQtKSjXmBPdEYN7XfORaGmcc/bmTWSz1hECDI6jfgcT
+hopxGNw7YogrzunE/QF6K6/Q/kZXbk+tjIw/QgzjJTtcWCTGtDpimq49mJQFV+a
`protect END_PROTECTED
