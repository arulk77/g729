`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
v2KxMY6WQiu13JS5GDnZwOpDfGdURK9APz+6yr1Ha0LRyhl/kIY6kparQKFpzgh6
h/tjnnrmmASAgWzRao2g8/Z1cJhPEpTuJYhIfOE8nnj18iFYHRjfGa1ARE8vggSP
Nk/jn6zucFNMq4fctWjLS3bLWojlTeDDzJJ+NSEkk7IQ952g92OfGzjg7pdoIPWi
EQn5KZSRXwP8gMYdbeffsosn0YHSkfJ8eZZ4979iuE8HcYEnzosqthAQNOH8egmT
ZBPRKooBFZme7ocpycPrDkhdOWLgxezlqz5aTJyMFZ7h+yu3w24gArLwbr0l5oTR
G5VBs/pbVPa5sdf2esPo7pu599qfx6vGabQelH1A/zU=
`protect END_PROTECTED
