`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePSMAteNl0mHs4wKYhajLiCu/TgWf2NkGxsMU6g+v3V/
2VsQMAyPNUENZl3Qn0VkdwXXb3c1OZjZpp7a7iqMWEhDmjV+rQq+r1Z0WZ/Ju7rM
14t1LyjhGqv0ze8RuEG5+y9IqAs+uRmnNV/73f1fgzfhYjiKarqtiqraC6iAf2eM
ykDBQ0oJHEN8z792SgF5SqUnEEER+ZbYQrxMHVkmwWRtM/3jTFeUiRkoifvqB6xU
`protect END_PROTECTED
