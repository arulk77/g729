`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOUfbviXREeclyz6qyfMcZXdwNecMxZgWbmLdAPJu7Sc
0uRohN/Sgi5dHEO/eBCvIWsLWmdjRw5AvZEOUGIoaRrmakUopPp5eSwH1hTe9q6Z
cR6tIGlElRmETgBRrl0wcvN6T4Cxd8wZC5G5XIJvHEdfyprpZEuP1BkQ8Dj0Ch0G
QGaJQAa9GOUlOjgk6QHQF0SQMHxvT28YVfW8rQHfuGAU6BusQ7aHDU23tOOCMo7f
q5FyWWogVRAwPuwpa6i7bA==
`protect END_PROTECTED
