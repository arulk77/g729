`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM5gt1sKFMJ/GXv+G1jYtp5TR6TNzjJznUJGBBJKDCIF
oqkp3F8rQorGPWSIvAdMeKxxCYF2Kb4WZpp8yNn73+ondvJOSFG88HyXzTNzQ5DQ
+mxfOuA4PfsgQPZor+P2mnjDR9/xZn9FSCIfz+3H1TXTj4VfW3nHVei6/Vklf+w9
Um9t1mN0lft5V4SEg+k8MSknWoJOhQ2stLaGsEWn36ahVtGgKwmTkebSBx+gJq4S
ugHA6YuXvYiuXlqK3DLjY1L2GnB6jru/tx+r2gz/ly6Aw05U2ebtYOuupHRutBbn
BMD2prAaLGgCWNfqUP1O1fZSPH+1miXnB+LVeXhJwQSy0/fL8qwFuWo2eqMEfJ8S
IyEZyyY3iLoAsP736Mooppc7Io24l16IjR5t2umgOhmHG7cIrxEZ2u7DYgO9VhPB
svLgdnKgxPvd03uUkzGuCmmtHuxdzd3uffQEpaEqAvD5tFtE+PVP4tYdNCN7uGXJ
0wQ91/rfAoTlV53sVFCfaW4L1d2QsMsPvEbxlE45NCSli/qlO3fkl8xyP283JRaZ
`protect END_PROTECTED
