`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBcgsURpL+Qvs6isaJSUrSPp3qwHr7LxrBIWInqsSjpj
2mM7q+i4zqqGnXWHXdVsiV82fwSvuzUdT0xfz59uAVcn6y/VfVV+3EBASm7IoCVu
RgFwbgJHpTHgsmFSc7UNZFj/DlsrydlCzxGXcbC+pFRepRVa+n56z+rO2ukPNfvM
JVROrW7bFOlggUlBQdnknZyVHAqdS5WN/nm8wY44Mf3scIUt5vzAnC54hjjMEmIG
`protect END_PROTECTED
