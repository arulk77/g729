`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73CwTYc43N1zY4+Upi9aqyn+wBWeLGNrMnzVxJlPx5R+q0
zmvVIUTX21db8K31hH1bySvRJCXXtfut4bZRX4FwMoZVGTjI4Zq0MWFUszmSx5EL
T8I0YJCSAoW7Ue+25iwhuCiQaFTjGJk9xSmGxxxzBJxsSE8PoYe3BXxgRfzQrRNh
rgCMNN+beBO3n/7XCWlrT8W1B9tbaDMg9x7Wkl7955QQ/w/Ay7Xn+GtrL/FJFiGb
BrJU9SGK85Tfd2qFzTVZy0n95p6ToV/E+UD5wc9LHhjjcKrcxxIEhBOU+dccol4r
eNp0txzJbfId5ZpTGyr25OzznHnynyP4u2VB4tLZG1eGj8xIq1q77/tWgalSmCpw
qvKXbcftFDBHbTKwyXHE5X9KsHzvxuw6viyJ78e03keRx8El/B/CCFHQLl+LeFwn
vk1LPN7zIFbr5BSirY/jO5GIst6jbA7pLEu+6J2ua+p2L3af5radCFmVUO/kRtiZ
0mTZ7UNYCnHSRYupMnxov2V0LpXX3CErwjfiTX6DO4Sj3+Igxz3YY8GWqViMJsXE
AFDEBWIZJQ7vRqExVZwLWlkvmNNOZrkvi07A/MyKyb3K+6KXOtLy69v61FAhGDKK
IfyPOUPCOGEuZ8lYfy9TscE0J2N0Xb2esQTG9WMrERBlUPmgOplg0jqrq1Z5rP6g
PCwXErtykAjgSxzcptQH7eP8FYmVoFkUCcmRcN6VMullamUkA57Sr1sY/hSzaOVx
SZ9rB+CurTo/DpePIgRr5hDVeeRnKSUUL1qWhZq6XcD3lZzIC89Py+ijDA87+2ZQ
vRWzx3EXoNnAHgOU3W2vF+Rf8dV0zD9C0HTCw4+YiRjgIoaDCV32hsJrJ2kgTdLS
vEzzd/MQwrYAbOZeF4jq9cfqL7egpXEiPErX75l4F/fYlBhTBpUvGB9m2o9hLEBD
kfvi/bJTrvPjVfZCNzeMdlYng5BmwDJiQS/BAJKHoYLWqc1q+a9SKhTpP0gsp32+
EVRNKWPzJ/Pp4cy7huPhyaH8O55IOFTfsKyNELf53GMw+SvgKCK8iIhmghGGKQ04
Gh/aUzXdixBMk23UpQyyzDt8y5qYAsuMZuxfZEWVk+q+Eg30YU9PS+ejUsmlDr8x
MJwyKKz++xonWAZ6LbDKuI8eY6K3eVFZwHARUEpWkXO41c1ZqB7wAd8WntvhhgQy
HnBkR0/t3Jk4+RZKbCx4fb3vJN7lxAXedqiJTL+bTi24TbBWj0jmKOowuXaz7HzF
cF/GHsDXAIK+bPdCwqyEn/yiTfi+YBADGe2dHYbZIqhOoNeXbgHMIx+jnRWfTxc0
jnQrdIKNwK7vYoQmeiHUbRxDmXeWdY9NKl3p6rcVFDGnieqTaRWZmWEjlrAG3lBE
lI5ZDQI5ZvZWEGVHlLkmZ0WD7/6mRjrmgaBr7hYKDhD0yHMGxPhTtpcTAb0ThYid
b3ch6AEV+6zryCnt4+KcG2I1tffiKOCGB8F2JesKxsQc4joj9xhhzPcr0K0RvXk1
JNDOeR7mMszqdLH1hmS2YNrOrVccS7c6tZpksBU3NCTlrgQjsqkvnwXkr+3aNVY+
5g0shJVNlkmiAxokYgFt71NS8qRtPdRnWqsRr2r9Z6eElBkI+jvPW0omuzUocGLt
q+2GFqPgyZA9JTO+Ue+HLcGon4FjJVrLDRMIcPuevYk3m8FpyYA9P9id5okUvj7i
lbDcQeS5PVCNemNLwtvFrYnn9Qk9phDi/ZiDV2f3VZMrzhD9OoyE4TJ6jxeV0wZv
dkmt7oJoTD4LdG8ayQ8Hqtlxbf885OFA4C4/WWY/FOxPUfacQY3sY0Hq+O39uvYI
k2NIBS55MPgry3LGTUiM10X5nux5o0QUTuBL5utKIu0lyczBWEaIIH22W3ReNAF2
2k+1ra+j5o1Wqr9unuimn67fKojO6hybvdU2+dLDRnZ75l9xhhaU8bfYvEql9C+z
iqVd+FEZsY2y2Urz+32A5BCZjIt9n8Mem9y/fIfWOc9zIzRV2UblqJnDQrwq8rON
1ZBlk5Ad2TK62N1jBu1N84BinNnTxx/ab9LUR3N/lkzjKqRgSZcNKJLo/rbgzXZP
55AOIcFUR8eXIrxRoxoTacXU9rR1glO/n74Kz7en7wOcsNk8mEjIjPVAD9Gie02w
PBQhv4U6oCPOEAKx8w+ZFczOadCM11lqmjx5MCYHOlckgNbFZWEUHLKEgVMCCDvf
EBiDf/Hi85jR2VgdEmGuPleu7iwHwLpwU+dRBf3PYf5PHipqSauZE3Emj2UwHec2
OpMQDMzYIkJ/ANGQXG7H3CS8zdXBlyiAwbyzRkjiAcCgn3aXN/jz704GPTtPDXn8
I7+PWT0g7stNokjlSbN5PMmHmGJR1BQ2Z6CZ0wUOrKgF/gRDXTN73ozUCgn3iH6W
uTkaRNjCP4/iLlUvh8/USRMhnb0EUzElgu8xQWEzgseXVuUsG7fKxX67vmMwVf/k
iF8FLusJvhCHFhSlGo5JK/1JMtpdwO0fiwkeseMo9SLZPnOm+uD1SN4u1XfBQ9vn
SGRt8RIRIkNZng/5z39n1oZ668Ey1Y8MMk/gkRTqyPNeGppcq1ECFgTwrqMzNT4l
qjyXDq3JWv1aHEkYT1Kw+8YnIff2NtJPYMGw068axbSmXDz/KH7LgWgumbPmLJPm
xbp+9mJa3MRW/d3muLQpR5Cr6LJlFx3NwLcQXe1YnC4x+ZaCc718GTJKyzx96w8f
rVup7W4BWhI7z7HedNDo4LlU+mMVub9fWRRYHpbgu6FiqAe93Obfm8RLaffJKfWF
M+7cdh3kkfRvFJKLqfbCC7y/W2rSFrPQMy4aC1cLPtsniL7kLA726G6fB1IIdENP
k/QaYoWeTQ0X9PZu/HFA+NdDn89kIDvyolaU1Gmp/q68GqmkidtuVfRveUR7Eou9
e/seyLA46CMa4YfYRn3dQ+ALwlZv6J2cM90BC9Lk5XOfLxv5pVje9Y7NVLwuZcqj
WhT0wK6jH1VIwcmcx6uV8U1NyM1HQinYkr4O/LjEHAFNJ4dzcmQ909KSOrCYgSBc
zQ74I8rQ1vB2LKGfJ14yhsi0TrXRc0HjtzM9VP1IK68s7RjgK3NfRndW+3Iu3CCM
VoRQqszw9Mlqwoz7qq8f8HF/h9tFvTQRjmRpOVMtSIMHtdnOSfKu64uNHwyVSYDk
FZUsKTrVpfdRTD+7QAaQoBHPwyuKOpcRF6ZJ3au/IXm0OkOZsuv95sd0Fux3bK6F
LTpV7YoWVmL92ETJW8cabo5mRK15FhEC0/xklbHaoFxZZNVbbamUE33QdsU42oCT
iEwLSJMN//e3z+m1Fhxx7ohbX/ZWsLQ3+xHzYK/p+zMuUOS1Wq3lLAN0N8mA03B+
7MacOosuvtKXIPoK0j62X9reMJCd0PEIXZUFrZOCZIpm3fpq5aXYgEQ+vlhxLSd8
ywfFO/yc840d8CF96X0zoiVX8qz0DZi/HcMBPVhoFUg/g+u75Y4uXAnTHSIRs/o3
CEguDBOpiN8OZ/W4EEEIl6BebPyvFWGOyJTuRqMVTAv0geEXfCUjCCjzLfFIvYj+
dMyfohRYtdGw1rK63peKGCVZThrer+CItP8cpNYsJDTu74V349OOjwvL52oG6fkW
QFj4QQqj3BxVW8ojyuTR/yzQnHzWVVCFL4mk9SfRWomyb2vQ71hOArYYK/+kcTBd
ng/Y4j5bgFxAJQOXYBnq1riupKjHEGl6YmznUw9BD/M3xz1U5rzwJhqTS7JVcW21
lLSpdtaiSOKx857Dg7H7ZBwXVdrUWPvv1NGAMTNypSNYEbkDRwMsgTXnnqq5s/zk
j8yTITWSEzXWYRdoKll4z+0HmQyDpt2CSHXHmNerLYGHHmW4g7J4FGfm3de2fHf3
KvqkP9HR9ySTtnWpl04w59xbczIF3SGrE/wyrhkfUE14Rvr+vCU9M0YQAiuG07PV
JY7scz/LjfReAakS1O53hmrR1th7V6JUgO+/IM/4db70FZFpAjq98F6b4h+5VZnd
3q32C3Kb2bsv1x+2fMAHR7NjQ125kkT6dkIUrgCQVs+FaTCtGWlpnhlrO4I65+ww
4XuF7pMLUNKbw9k8fDlTP68uRhKwalx0b7GkbH3hGalNI8DOV1QQztPdLJTgIawO
u4/8TQ+cA4YmN1rCXwotkcWQL6v6YREPDAjh1ENpLkQaBfCxTJao2i2SX26m59EF
w3YrBBRsAeZ1UqFVNYwsUhc/JoE/Uzf+66fBAVkKIsdFLudo8h+ZvMx80XQobExE
j9Vq0bT03rsEXNawFXKTfawR7u+spuXlGsb9XgJBprPn3gzarcGjChdzykZKLbYt
tq1stU30b5JFVAZnYh+LUKlj8Hd0yGiUaZ3/953yFfIManlgtiQeq13Hdgo8Fmfs
FL+0Rn1w/cLOAWrkuKSAmv4rsauGnv6xmDvYGvvV/NNKZFYwH4fL+AZFUkH+X7V6
ILjECNhlR4ZOYEZT97MzBa9SRntvZn/J/i6zpGXP9innnrLRj3VS45dSXDFffrf0
8F0BWpB/iIw61l3eM9ixKuattEoEUL1WrOyTcbIXm9A/b3Y9j3AYoqDzeMe7vw/s
/eWIyi37jUUqdXK9fJaOZF6gQumPnWTE8acmTIkQ0T5LvSHCsXlzorFFua/LWBo4
kMFcxYS4rDk8CE8qPpSQc4xPvrhMMtJZm7XgJERLRX8Gk9zq48znn32ADhzGAS62
rmC6ZFF8kUcYnhdPtSbusKKkagWTsNnHWtiwUViRkpiClY7DGZ+3Qoq8DEXVZM9e
9gvXXuHZSxnc2imqDJoqSZKvGRQsNV1ZGLY/Yv2TSvTQy1A0InOsUZEMTu6t3o4h
tYAUp0nmGBqyrmj+BmG26XFhdUCZHrDckG0GWblLLZ59jE4f58XPjF0gaMYwxpWT
MJX0fKWXP9s4CSS4LYhoJIe0pLYgpZtMkZZcpyWxV1DGEWc/54nyr1ZPwTESHJxP
`protect END_PROTECTED
