`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41yuj6Au0wFMbNiB1G9Dp58AXn/QIyClY+8XKWWFwyqS
e0ydxdOvXjnvWf2pd+DIYW/CUq3iZLT4CLvhKF1SCNQbgZlLYHHdumPS8cbZMQ+i
biQgky1ZHh28LfvSfztCNDoN9EY0aiwMySJTiG2R10ijkyaFIUCMZ1GMkJga430e
1dT+qtWyrcXCTwsR4ocw3hsDY7qmZo/Guac9HR8ncC9bsflUIt4KRgN/xMCO2klr
/6vhUbnW2U/zQXa24tGAsh7yKWwwFgicwCEittYj3fM=
`protect END_PROTECTED
