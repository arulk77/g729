`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xg8FL3nS+hX21DHGvbY/qTynsV7kKIirRNHZBak2fzq
WqdoO660kpNk0yZoJ85QOMe1rxCkkbh4QY8tbwx82VbqoB2nYXzwOHXcZ4RKHfZJ
fPlK3wnny6gur6E/lyCADBepfRDI/Ba9bkN4+g1z9BQDZA41wqS7uqxXG5yB83hD
amz0qw+ZVsCwlZ5FaOTB8JlX+JJKutAmMW0tqRpoT5LDPVnpChI6c78k5TjwlEkg
JmIQshEd/34fqXdMPg/Zej7vkpJpocm40bqzRl+qw+U=
`protect END_PROTECTED
