`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2EBoZu9tBf8wFLCnm6xiM63LHihYlMRJIG/TA+B0rjj6xvYbsI39y+BzfmJq8WB8
iCYPuwZoJLKL0ALFP7woTjJQxTGerf9zh/KjnTXwBLFYa8am/ZFZGbRLSvLvzs/A
+cHMN3fvEW7lvNl02D3Er3r7yzEXeutKVcNmrlU71ondfNinwoYWB9fY05XaqzFN
blrDwsCjsaL71D9UO1tBL/M3g+FYgtmqjBplU3b4rhUp5oTNwZx/oA1U9eLqhI8T
DGmX+3vsqB9b4BcAedhRzezepXRWWkMGHI+6DvavKD3ZMXbmFw4NWdnsEi4WvXF6
`protect END_PROTECTED
