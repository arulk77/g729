`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
DxPrAow6Rdk2HfSEn1uvxKQLpwFQoG2+dQBvSJAD4pjLR2ycWgPmpxWmKV/Jls7n
6apuuH2NKnNQPxjlH8PYhK+sC4kBOIVvUGtqJ/1NBlOhJas8Q8JlWuwvTcE0Nn5A
72XOcJaplLV1fPPpsDvaJRKflM1hYmDPkjZCfQSuco5QgR+p8KlLJMNIFWhVEDbL
rNQ3PmvpiNVN0OezrbqCL3mMCbdIWzCHdmivRj5xI4y8gLc2Mfug/xZjgp3Gv77M
RjHy/2+6rUzBUJPmo5aY0lLqoncYv3k1YGx1VpudwcRRirhbk78WXzdPoIZVMTUe
+wBAM3Z2i1c0JNpPl+1ePA==
`protect END_PROTECTED
