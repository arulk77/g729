`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xSxxTxydpkr3U5ZRtGNMEkkDLpT92rbRxD1cdU24TSc
55SCW/gnNAowKcRHHZDxGtY41yfikrBunIUfo/dftQXWa/9anjKoIZn8z1oHvbrJ
fJ9b6LvDmw184OnC08+NqJufD2kG0vZKvNqe84VjTaXqtvboAT9m86W4nFbfm12F
zB81p4g4xjuxcaByeSzHoAT8sZzgMLNEr+t5hQhKglE=
`protect END_PROTECTED
