`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aVXAUoR1T4GjJhG4vaTi9CfTUXBJKHgggLqikTMT0Dsu
daFx4odePsIp+lKSgvNi3Ooa6AOG4OXsxCXXIoxi8UB0rualDrMSnBAINocdpWB1
8EPJABrWZRNbq35eZujMB396xr5F6ky1l/Wj9sWs8PFbV7bmA7xHK63X1q1vafbL
QGj9V3vtjtRp1KoHsNSuWJZdhsJBRh9vMSOHTO9emZEsV/ViRBknVCR9jMg5TVU8
PCygSflDa11yTaFmiFEaYm93A9s+Kxp8yQU5Ae+64MV9SxOYrdn9bvC6aAphi0a+
n3ykYu3vbrk8XHLgSWY5Pp942O3nADt72IEyblK9uYe/LtzZLFj1i3dBSxjncbwR
blMtANQRP24nDZBGTxb5GJSzY2mNkRtoNVwEk5ME+tTjXXJpxsorhjdbFfJUikN/
CFM/NLgl82obSyMwjBYeB1v3zxs9Cieni+3J+0n7iXjkS2Sc1YkJzX5JCuIV7hyO
wqO2Lk8AlGB46nXiKuFxGKgR8qUc8BERCvCHZ6n8Z3uiB8vav65iliWF/xM8V9c9
A4WUpKCO9xwdM1W42+eOu0pN3aSo4ituralYWOO6L9svm2o7tL0akFGv95JAU9/h
WNdTEp+9UR49jTsJ0nhGYr0ZI+lorRM23nsZWmUUO9YmF19DX8o4cpM+wD4ndDiU
yfggq9ULtwPIYgwKkflkprBhWx7OglQKe0rjGfRBNL+GMX8AjVeLRzI9bKrvDi+/
014fnTLnpSVD0VGQWy1JAvQzfguqCODfQH9gCeQM9Bdzw42m2dwTYjJcERT3QVES
CDJ49PcwgKETdaDGpU4eW5TLFOapi88MVYZbGj3iw907FIYQ/6fqawg9b2MEk2kV
36G/FUTXxB19RhSha+Qw7DmwSqjSTog65y74PAU/uiWzuo+4+L1MKkTn0YuR7xZs
/lwjWkN/B98h5p6vv1n+2IQ39jTte+RF8KiX1lNY1p4eGQbzKh2MHDu2Qn7bRDmq
AQlcEKa6ztqr7iyKWJXmlMNMqk/jixrVN2Ad5PRYVqCsObLhCPgmxtWkOpBmsoEZ
IjKulaH01FP7CuYgioEUu9mqzOf9H/32qB58SoHB8LDJdz4APbsNd7mmvzrFbdhl
7PqFIIfA0hTR34dfCnFQUxuAhbq+aQi2UEYueRz8O2L4MhIcEdOIQz1QpHyvDIlU
Mhu42LR0VaTxOz1K+GfGZ7CKB63/AkJVYGyshbNMu8KZzjRUC3F0L471ntf/V/Hj
6OihdHo8mNFTQysoDtHWkXsPF881XWomOZ1TLb2UTfiM1seNWTaelZvTB9tDjmJh
btGQBzPsIHHmKHrU29AJqmGxH0ecpgCAImalLOj/TJM8cVtct4LRZWK7pONE4ru3
8LAFGmxbezqnnKYCVOazUzYrcl+c8i/o0q7YzDkarEn9C9FsSW50VcRsHrDyJqTi
AVExf52cL2qNsdZHrClotzIcwDLnL10m5u7F4B1RlQksiOXtsT0Qalr4Ey7PQbSD
oYvG97rj3WkvMiHv8XMghPucv+9rLqsiNGnzaK+ssC+F28ts0ytx6BtP2sHkgyRP
Y0Bli/PONeufcPYMzezAek3NvD0w++TFZHtYHLJK2e4mbSa2rE0n+B9DtQhmUGFV
xpt+5DqsJ/AUnMRV7hEDEO0tD+Xf+OAXVfUGNzdrxHO/5mXXhAE2mFofvbe2iptK
uy+tiARsJoQNlSYHQJccZkpPwZqTKDxJPh4ic225GK1qdroHAgauLRw80XKrpIt0
n5isFs5Z6AvBbE2+o5byvWnr7EhYTZVD9qSOuPg368oQ5uJjY7AQrT+4FJsv1Bo4
9YBmov1SGGcwVLCdQWMHxQv0y7gVLVV1B9aUHxPuVo9ZwK332SvW9oZ8hZ2/Zose
1rvYtex2Ww92sWjXGzO1SjAfvr6x0X8g0plPMw9UbDq1UuR2D81dKzNmG0CUkfbg
MDwc4GHtuDpgDoaaVcD+utS19Mt7dLUTFtABTqSH9RB0AZ0cOVAWXmBtRLkj6ooQ
QSXmvMr3F/ugGV/tslFriYB7opG3tFIIHf5MqQ8n/C5l8KMGbQ/iR/eCclcE0ydD
9wHb0lwEYxRv3WBsWoeY9asuypiIu7ny0NTpuSdhOz2nDPlfmoVFr+AvE4DkYAkJ
M89EiGgIbNZqyWzEkUAiCJ0itSLdVhInnzsHenGMDDVRsGaGNhfiIGjuNh4Pa5qj
DnBaXQxNnEZJcxChtTxq6I2mA/r96YmDFq180zwGkIUYl6iQotJ7DJkHcRbUFNfE
PvbJwjP4KvuifljdmwNyI2UTe52aqG5KdnZ526jUZU5ObAzBg8KeJT5Y9342DU2+
EoIEmHuetyEr9iYpEW8ZLXi1/XNlWSzQBNht7SoB2nj5mQ3GloXQPsGzTHK9dWJx
YRCM72Y6d0a11CEAs5zxBlff4Ah2PTVXFTNkEYt6rwcv1hKnKil/SO49IU6Ao4SP
TCLiHW/ijqZ9tWMBfW9gyEsK+cxw6JvZfQJ9qc55wtk=
`protect END_PROTECTED
