`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49r6UZrO59Au+OOYUlzzWafP+SdJv31cNrqPmh0xM8Nb
O/QW7C/30qD3hXjz9bbndBcCdlZc3WLb6XEpwllPxi51MFx6VG9AnxyOlWcq7spo
OYSOxuzw/VmkDunkaQWg4f5xkaGgT8KuMfF0VmYurrEQqGEfmqtUB48RhR9ZLQg5
S6Omi35Ed0RYOKkp2FIx4J9OTM+STkSk6+Yf0eIwz24=
`protect END_PROTECTED
