`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3fD41N1u/Hva32Z3/4jZXNqURJ2AnOMObwW3/M8u+21PmQ/5i669PSJwwDA544vo
n4njLcPXEfCduma3NQyfkmUdUWqDzq3CwX9+8nwiBXPd72j/E2Lz6HERQnK+VZ8p
xcJdJFM82dB7xa/EGiZdcEc5Cs+USVvinjCzvxHaul1NC560Id1SGHvt+n9HCeih
rHW8WaiPF1T0C/X9PcCbs6Vv3hZpkDLYVEmBUYn/g7Ok6tV6gnIpI+K7Gm01WXdK
`protect END_PROTECTED
