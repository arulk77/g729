`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCDaCK7RAPpgFLEqtaqGTrRXiMxBTE3kYPyYWu5wNJqs
xiQSPR3ffCRdnnh1qgGHLGMHSfbfBJUWuzuy01gU8R4/R/hnuACwN4Fg1dL9xzKV
kovuAytIaXkRMgRPfrhhx95y0DRxovDizryTC1tikMI+uOPO8pMX79aSoTh7U76b
o7ydzVCvBMGwkgb8c79nGXh50fVjUWNpLR6KlHmRXtkCiwjPceIG71Eoi4DVfHuc
B7IZ4H44hM8kENg0U3DFGj+CvGPBiJ7odVZ4Ae4OAuWurFelR/0jpz9MX3L902+w
YOClM/zuvRnRj8/5s3jvc6WnWNYbG20IB5WmeTDxjPRat4Ep5kb68k/F6WToguzO
`protect END_PROTECTED
