`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEevyIRYNoXKzSG4YLzmRTF+UblOpkzBS54Ib7fmbIPp
WVkRlGDypyqySFHDbgojgtJ3hid5vGQYFdIWQCcKV+lt/HIwaL2NpEM2B+FxRRyc
sJxL06jjfQayYv7gmr9hJJ1FIhk6ui2dohSsg2jmSvXGLbXX5Zmy54Mnd3nkM495
9TlAp1Kcg+uhHG6EjENgn8R5+kg2aPB+9j5rEPuIHEoOLnuN3idHIsGuWLkGJixP
0QVohyUJM2itGH6ZiythaVt3daDFF6r2hvCHX5IKSp5r3RsebbC5B2Ebw9s5BGwx
5r9x5VAgQE8+kpPq8kNylHT/VVH1tCrtaBj3dNEGAJ5JbBmOawWiNEvR6SAhCbz9
Av/Uup6BynwkfHCCUBoFSoOyLVE/VE2InZzMgc8uv2l4H+1v0XjBwkeRj3lgv6+o
nJawW0DSGJiL8ERyahN/EQ==
`protect END_PROTECTED
