`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNkY+kAi3esmZkiTuUzF4JY5+OzW/gBoapWTlN/yFejd
LO9gg2NneGxZHlYwsI/zr1paoqyg9dEuXtqzujukcHqgcFqOHFEvrotQo0U1G8Xu
AWGv6YjUqcFJkja/wCOZQ1MQYC9bTUdPMSBzvb5cyWjVOEDtRVT7F8NginIDgLkU
+OjPUGVTum9UHrx+eheaQg==
`protect END_PROTECTED
