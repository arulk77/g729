`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aQ2hGJlvb465HNJ4rQZNRY2V0hkSYx948aGBA3bNyrTZ
dKODFeUGtDzqbUGTCzT7pk/+hSZivn6tPOFHXzeugzxplEuwSTxzB/K/yHbWNRBD
BGbpJoCQmDDa96WnVK4IkpqugQg4nAkXOukinF3K3wu9IkkXGwiFMlXyFNgEXOi4
EtQDSBgg8mgRL9+WbO/BJp+T+birmgwBLa9RZAx7OZ2Uz98A3c3pCG2GC1ledHFO
ASj5MQc9T5zLmsRjJzI5C1TrJWSyX+EUexaj/f8EM7PfYwLZWVCSjmBnG9M4/WI6
+HSKXJMkHuR+HRXcRdzz7VODRXFcA771Lfm/T6b//lOemGXpf98R/GX0POOzCijP
GpX8PVqupL2g3UAWpUUz/E2t86k1c/r3zgfO+ocT44etZ9BUjcTiktz1voqLEiMM
Xw7uSVpe6nObY2PUMEeqK1tRNXdNi6kZZDKYzytcAIki/rBCykk8XRmxA4D2JMzE
Fbi4+nxEnsn+q8p9jrUDn2aYRQvZtyv/zoMGboL6YnTP3wKkI17VjCGXb9wGpZl1
G5CZdQTP5FFNTc2M6L9CfC7bisibOR3iOpuiMfNr/C9h5o4s9+zsSBh1FiRcLjG5
dZF9nDS98qfuaRWApm+x2QcsEIyMM54UMaZby+2weRxyAa0TlvxJ+AHeBufPINpg
dZIVxDic/Ja2tMiefKHnd79yxwcMVFhvxjiAAyNAhdW9YinTZBvc5/hK5QoSTWVQ
Mko5WqoMzaN2GYJhBdXdyDIeCcmZPWveEsk2r/an01UbQDfgzDMTx2u2iS++RCyI
49ioSbUd5qNG3QK2a6NWO4JAcMxy3YZWKDsF+JYOGp+3w8iFqFg1fM/cNJcRSgz3
9goe4HbRs7MZQusn3TbbsiIHvNA7PzUNF00AE8cGobQ7dsZagZGd9tcdHXMTKb68
3xSZkvBXWp8sTXWhEsVkTkfeIEIE0SVQ8M+nN4AYsapy5Bjuog5nfk2UcY0a3DZ/
IV6dA2JtWUC2BDjbWXz2TX5+X7WkneuxzgPtzPYAUB5q2gqwqO2YfgDECG6F8TtI
dYeo6oIDmeaeRf9IThAcUHlurBFY0CRsXvjvHVozgzJKquG8YjQ2RMneJj64OHkm
VHQ90EGbSMWxjkPx5bYnCEwlpDOCuu0fx3gTcVbyCqh+AoXBaSfO0KJj+fAZOdY4
FYucrUNOeWopatFi9kk2Am119XIUt9b7GuYpP9zvYrszrKfDZo/MdeOuqKgETqLg
+YpHJQpZrESQgLUp5m9yCQ==
`protect END_PROTECTED
