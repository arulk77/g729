`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEolABxzpqICD8t3zWuF0tCdLKf4aHU/AkRnwJ5bbzLM
DgZfiSYNWreLziEn9Cpo0TTQWpxCHM7p3nICbamjvkinnYaC6ATGyUTeV9vTpPLX
DtbvTuRRsnZgx4EScu5aXvJtmGwse/of3FB4rvhRkvBRtqTZrzs76Kn4JzDVZPba
ibxuYXjFruVn4AidFVxonMHfOMGUTKbMsJJIzRnutPzxfZJEn66lnIdu4T+rbjav
teNRbSG01wn+4/owiMKY0lP9yWbUETzLJaASIoPdd4TNXK0tsu5StLxjV3GxiZ0F
xos3I0EWiHHietE5fAF9as48nr+fXKHj3aMdqcr358rSX92eNbYBzlYJ8quv1Lik
xUfVz7Mf9JiUXmTMZEQSR0lgl9YJZHVpMgF9OU6oyYSbBkGXykimGr6TsTYwM2l+
c5wj2NGcSEQ7RH/rAnl28N0y6zSorQBxNhC58pdjyYPXXqFi5WADgLEgPk1c+DzG
74l1bH8x1m9K6r+1bCP2/AM3pcy24Thdq5/sAE1k71qKypgeGRwcDegAjKEDdZaF
S0dB+f7kkSAf6iAmMyW7JES9/aQi9yUdje2HS2z0bE+R9wLbvD7TDZ+dNDDmAU1+
`protect END_PROTECTED
