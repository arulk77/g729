`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNN2j4hywYbceGecnmlLQBhyDvcNPeF/CNbY41n3HsN4
NHzBPT60Bxq1LcraTBMQVewV4bppbAmad7/G/tQoSgg5/833BdJgBZQHuQJuVFZ4
HcW0qR7nvROYw4SgpmGrHjvTcAkjirTuB5n3elgtUOXRsb4/AIHwPLA5x/ajYAo9
dqevF9pibpJ/0zo/u3NJEQnzV1xvjRQCYNydDJx1kVYLzlpBZ0cIF3f7zdGBJtEp
Wv0zJx8e6dK1BpeZK6cDiamIP39FsT1Ke0KK2LLQ+thg874wKNOtK0hrz8EyWWAx
KnjmYGePZB1rVRbhpO21lGfy6NlpQ95J49VhCxpz/wm4ffnRBra1cHVtUqlNB3pK
pOXyxURxnp5OuF3aiOhfXD5GwX0nUHZFWEYSPIvvH76AjNaci1e2WWbrDJ5LqXNc
fdffC/yjuaTuXMf612Z1uDAB3N1+WCAm6TVImC2iEnFrZySGx0flYjckb/u7zO9Y
wE2l9547mgc5ryV61giaG5F3n6kM99N4tNalYrXFaTRxW4oj3r1oNFMj5Iv7JIjc
WpfTiwWLj7fJ/etyJr9ykLIbZQaFmuD8eTPNG5i7OyrI5JUUvm9rGSf1mA06t06r
gL/6vrNDk/J33qAyDfIBst/klhjM5YaWdC5xE4eavQkIA00z2thDvbxwHbJ+aMXv
rnNXFqU7IIUFX9bSsP0yiuDyBW5stD5lQTgSzgpwfizf9e3Zv7GoTcVQmICabIyI
qhIqZqJ9TmnnYWxpK48KeWA40UB6olIIa7T15vIze1rlUg9+tMElEJH80/tnqp+V
WriTjZG7DWvEFmIlY6H4AOdJLKtTpVDoNkuV0aM1EhU/f2me+6mv07uRkphECNTo
9FzoZAqJP03LENbwSy0BToG3p6OBJTrHjizaW2pwWiFClKWQFZKqqPGUM0Dksn87
8EwLYcTixBcrOETr3DwnxrXDqT/RHGVRP1Y1iR8R8KeKs/sRhCJCVkH6ZtbdzkF4
e5WBkSsqOUqKKQw4TKTgPCRstxdKZbsei27tvwtAcn5gB1nmKatb4tQAt7ymCsWQ
9bNmgOwO1jl3PfgFZK3QRfmSYkdWqFMDuWak9agev5c3QnP7/IMX1PuDsWLP63DV
xEwVgs814DR7qIHyurirgMWySqn3yLqN1lfnSgMxNrnd/hiybZsAEt6s3REkaQRp
utkZXR8MmNl+6W7Id0DnaykSuB1O8pntYl5Y18UWijxQeraqY6jm9ULXFS1tPAsr
PQHRl57xr5vj0bj/v1vXBn1q4i9iCQ7EQ5PywjRU0cjtE+xFke9R+ip7NyaqpSUR
tzhrZcuAwroeEnmC1TKupwyBjru5S1m5rV+XnKTsB7En7AmulGx9wZAcfXEmvmr8
4YJasptr0iTTvckg7zPpc6Y3NF/5zduG2Vvsu9SHuI/2th19FfP7xbd917ShFCWp
w9TMSSZwJMJdf5WrLoTtxT3yXcLNxbPLkugV9ZlmG1GrxH33C1xfaKr0Dp4nlVm9
49Sa19cgIXCReFn+jDjuFMISeFhpTKhQMxtQarxGnCdJMjZY0Urvf/pQ/ldhedf9
cCP7B6LVRgNfJ2oStnzKlLuADKFZshraLKh+6x1Nqu8=
`protect END_PROTECTED
