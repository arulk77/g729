`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAfEjr0boGN8oh2j1HVg75fJhtgqFGfWy0ObpHuOGsQPg
uEaeq2i3yPjxINa+71jtrKZ6jOofodWvLheFmKb3iHfGZUf2Pogm3sAbddEfXwpf
r+V3Oq/hnr/SFGPvP5wdOXPNojBQPUh4a9V7kYchbcKgg7PZpyMEnuP9u5SZ3UHj
06TfRj/BWAKjIFZ1e80m9qEV8OFeYyweZw9fv5G9V/uxvHnUIn93OJNeJLCnIG9V
jVd52m5YonNPG+tcpXazpKCU59lnRDnMaIrz3yYR1qi9xqYtiSs6C1/SXE8ZCRp4
gbG8a3GnC387tmdjypisrHeSV19tXVjQMbXyfDBZ+NLl2yVAqE4h6Ebv31vePwJ7
ByrU4WTyi5L4Q+9vO0BK7YhBnuMm9qSmkBaGvELlr9m5Qts4dv4cH0mcHLOrWKz9
VxhauJV+7qndPALIlSAqrhwGWexaQ7YPTt+HnLErPHgHVpmNL6cjQRYKufEnMlTY
5JD3lfHsyTlnKo/2PrAIieYZfdnrJatADOgZrfA3JuVSw6W3brtRYQXL50R1LJU+
TnFbnF9L2oynTceTWk37DwCv11VIw5w9B5oHzeeKaiXPYQf0PxA84DRbXULkL3XY
ZJ/y+YOoctQGoisStC7nooHR4/9hceszl6XB9G2pgHQmf+bkWT4PmI8hu7LsHxwK
6jGgr/NoYh6+voYawrXR8bqb9I6F4CTsSB450hyX4CzyRucGfaW3FPFPesXb8vWI
e8zIXbyxksZZ0NQPSn646kpyIBlwOVNO0QQuQdSQtZkWrX5L4b8WEb33R/Vgp73n
YcfrHqYEau0nKNBBWrPMFZKq5bd5CYJb75B4zcho5w+FPUwxzEhMtqfRir6eDr/E
Dthb7Q1pkrdT8hX7BuzjW9b3NsPTK6hFCjoNLUd0/OGMz0mxn7ruUFT56xSJTeHL
Eef30VXXCCz0tqJUX1LFV5ouxlWGugCSl9diciiK2iwmSSu9OkkshivEIt6WC58F
EGV46Imv/GlKMkal89aQ8nrAdWkDQVpSIT74z548CW/zuKeiwSGgEWC/13VMp4an
nGC/4yIfNAVdvqXO/MlcL2HEpDZyJP8AcRdXRRwCFGoWR1IEOgrZAJp4Y/KOofWC
TnwLZ3u7aw5UeeuUrMjRc5VplH0P82QxPLN6Yd9ze4xFM6eRgmj3K+elEH5rDj4m
YsQ3GFUyAtgbHrgci6wuh691VWSw8q8966g6XYROv+5CyAn/mqamd8QUgwXAq3Bv
ODD/+AlS/8BxG/TzYdk/sO628EdHv6M4bPLnOfrvanG/e3EdCfbXxwckSnQ6mm1Z
X3PE86XAlma7L0Xc5XbCS4Rb6isE2j4/+53fcUuI+1ItWBvkehXUrgW2lonGaHqY
iZVquq8YQ0lu94HG+HgaBB7DjyhByO9yB1XK6UUcjSh9J+fhqR2lHEFAIfS+UzeY
XqjCLCKcMajxG9Xcf1vHt3lpOy+tmDjGUypyAag81kay4Aukf/6YhtWbUrQ7hBuX
shQvjMIc1be60/Q/B2fQeXLqdXnzij/IfwOxANC97ZVVyuCNaVyqNg88pDeoIqfl
AqIJ2tsxJnneRRb6gBYZKeK2xtQXVtAxGP4KJoJOjGpjpIP9orQhxuAHgH5myqfA
jzlGgRTKpLC2ckdI7wo3jvIlYaVxXpgYsGEamtHk44uE438/0kXtMnkyv4tqz5nn
Dy099qsMQJKxwWmPkpAX4KtJplEvVEtqvPjBOMhgJbEEQ0WKtEgGLhiS4ESmKinW
o+pbuACyoHsGBGBEqF6bMof7+Ng5d16xu8hK4y1aH2AxL/z3ai6REwz4pRXQBETK
xZ0E2rPgQ7BZStQCcjaWw6AvIR5UBrELYqSbwPWnz4O8JsHJjaJoZeBYf/pP0tIA
pB4sZMFT2BOJQ6FMPdreSUxdChh9AGDKQ5XwDQH/vkb/NKf2pA2IwyVzEhdw9L8a
VdE9ig75iVQMHAFynC1BD4CH3MMaILbk1HS0645x9b2Zn1fKiG2q1xiYfpxd3zr9
uPBqcVaKS0yUCiwRdrk/LZargXfOsECkW7sZW/u+bd4ha/be7blA6t1T6RAJy6QI
jdA5vJG7i1WDbbRIVhGCdgbjQPOlx59vqCxN0lbYe9ODKrli3C6trs9dKzDtslV+
lhaReASlonEteRIcIBFkCHgA6KAX4AgvC+PjGdzWWibJC4JgJY+dfyiqrKI1No36
klUglc46waBwBl2RCfwb3rVXmZF161xnKJmv8ffMa19OwVilBZU/UZUvIY8QXmcV
eaoFXY/6gFDzIQf3vmRkG80mFOXHO4xVEim/saLS2HBHnPfJCKOFgUTDbASo7hgc
lqlcyrUAIvJZml6bqKw1ilitEhTFSdjyonoXkI0G7ty1crIBlEq/H1se7ARhDuPz
JJO44z3J3KDwjNTvwulAzR5IPXDEfyV3XtDHj95M3qRwMv3/9vNUMxj5IzjGOy0v
Zm7o3A3s+vV13hoReiF4yxDvTDmhQCFjlY9zEJQDLrCIL2WehSNoPjgcPxDLbYfE
NgA7S7HQ2F05c4YAbc9KFd1V2hgV+PiFNKuHglkK4aTousS+x6cLoGIcgOBAyvjh
TErxiTjfFPH2e+sersMsw/4VkWyxX9HBhbZGRE2qrStQKxH9AzhDVSUZPMWB6BRK
beuH3cS/hNKFlbFz+XqTTaR9Y/XTHSvB3ByMsbNLvQFsqTaFyH/n87+HcwZW1cOW
9YtR7uZUtezCnozgqR0AjbINDvZJQnVr2Ts7HAbnI8/eA9gvCbCFZCwvoL6I6uRb
pVvliYDK/+d1To00PkM+K0pAlmfaV2cSKRbRuWM/lFrdg2I0YU13NcD14A9LN4wC
tZ2k4J++xp2UPl+4OmlMXRxw8BRbjYirRmFb8vZPPtWwhlW6Akv+98lWSq3dwFR+
iaYDmyaj8iEEMyioA6NbK6OCsPraaE1x41mYpLpGP2tbupvcGi53YJ4NXKb7id2B
eQJCMYZsF68Cq4kq2lEw5AF1+aUTdh4JGlz+Knis96t/IqOfUl1qTEuIEvq8ydD0
2Hp8Q2C47OnVkarHAJ4QDStb9GgVoZsMZdP7/o9yroOhPhLMBIqGiE7Oi6jbdIrN
FPYDoovtbHwm8MLgXHv9JsZQ3D4SbsBauhQy/ka8LDzNOZrAB3272Hu++2MVosjB
V/5UBtBKYobo9svoolSU3xyxGpKT/9uKJ50o2ePXjrE0n+dtLeRJaLFSAKaj6NVQ
wpNowobAA81DRtl7l+ERi2+Z/r7uwZkS9qHgRU4NJNx0pVmTUKDNNHZyZfDNAaoy
WaH+n2Ti6rJjU5xHr4QjNDW2HP9aha+CFBdZ7fHQ5Iuq/RDxky9K0foVjCtOGyjK
WbyVAR3hcBAp1IJaEN0tkMm744oZTNSd0yxgcsUi2OYcnxRycOS6hhv/7ZXXR0rt
BSWCCNV5G/tllTa2TWTBJT2t4gByvFA/ifNlDzweWO0IkwKXs262oFPcg//o1nCy
asYae5Jr42CU2TC7GKpZ0CicHzmWifvx7qzfxG93aqC9BvMm8Ishun/12bFBAeva
sNAYO+7HZt+07tfditoucDDIStREG5uxiwLXdlO7GJ0OkoShbzTYlv52uHtzcyR3
NqIqdQ0JIO+x+ygewm4YPXvQZ6Rw5i8Rayyulj9IwbSXgEmYSgFYQ4QepUgiQxzr
dHnJW5WX1MDZ7dNyQ60uHzIlkJ2AA7/cun2q1RsArrkzFTLMdtZlretgFka59Li8
0r34BYUdkgs+nrWirNRTNrjGD4dy2ZIh6KO9z1VMVvEdpBbxcnXqFZ95LTbIl/rr
x6c6xBlwrS0pRoY8kS9097bFI7xCwpEeqAnsc8nAwgLyZSqs9mpU79PToE0b3rR/
aqeC7zJggXYrnmDdB5fF3SrBMiJysqUnHJXXpcah4ptXNdfpZRHFMxkDYfnlWDj8
9q38B5byy6s/oF2HX1mcs4yD9gqA4GfcTZxiYSzZ55XLw1pkxSAFAdTmYQ314pAZ
AoPbXXv23jmoZcG/wCtuuRCiAg8/OSdwdI8QA+lA+P+OjkS9UXIKwIGsesXCtjdG
JxPx3fRE/J6AFk19BFRDWHRxIaJkzIcBmdwVYR0UkzAl6AmP95Q1Zz6mIxIbqJdZ
C0Oi/TT93G/XIPV8YffnVdbEgF9l1s2fz+lrmw73tu2ApGTqDtiF1FWgLjwE7f2+
C263/CN3sQV2k4NPMdc8nS7T/bN/0jYtrooTEmUWX2OmlKic98kiwszsLvoG5v/c
4+aZ8jpLhqCdeSYY+VV2PfKG9Ulw5hCBEWQqXjWEZZQMDyNA0QbNSeSSjlZPGtcn
8y+VYgypsdwmcOYNI78DNr0KcDjPulg0ihLX11FiuttYoN/oowSSggG/VfmW1ijB
8HmO3luiPkACgI3T4EO9OFdZsUOqT8KBSO886VkpeVGFtVQ3/krVAsqK965sRYB1
IEW0lf3TviaVsiSHNiwTWBV1lPMFK1+V63LFvfMwfDpHG6auxRzOZyDHjJrK582Z
01YoH1O2ltHOqY62kFVtPR2DPQ5K+dgREc5aaCUix4QXaiY3fEJ5xkSbASEf1e8J
nC3ZgdvOcEa7q74FTgiAJZ3KqK4Zxik3YYEXEAW4aasDNrOGEUY25g3Ed0JLsMOr
9aRZFTa58+YrzwZw9giOi29lcLGg0zdMFgtDAswcnqBTul+yHQPmNgxS1C1BzFEC
NphzDuLDl8cLDWuNxaNcgxhHEb1Kl+eIcg9xLUO1rfTTLoN27TQESxSpEbR77zgN
eSDhqmssvmWKMOLmF/XmbZbh96JBFvpsn2u7G7Us7xOXQ5tYP+usdxzx3ELcM4hj
3To4V2cv+OrsupgECMpCzV53PNCojRxHXhT9xzzqagutTuDeyGk4ZL6gjTeTgAX8
7UYx6N2yR34eCGjsVODREtx3lg42SQ6AE8cLokV/+HN0mHZJJi11V6K/4XiJ2sxb
2YwJkBlUTabjvbopIj3Mu8/A1yTB7Ywc24Fr1gdUQrHoU7+s12cNZhbRW5pHSNJM
R4EOvsQnxITTUMz/POC14q1kwOGGrQleGhs21cAExOBcjsit6pnpgIFZdAxhlG4D
Hlnc++UfZsQaDL5/yoCCJIYKusSZyGzh3HQZOpGf2d8vK1YNGi3xhL+oQTLUIfaQ
Vqw7ocKgCP426bi8qxc0HVkEyKTVtOZs73gqeeDiYoJiEB1SsCNIOxF5LuYv0g2v
jFIq9jsH5LHFU5lp7YxOIznGjfTdzXcUVfQI3W+iUGPBemf7Jry4LQ4vpbDCMsBO
m0p99je4n4yJxdXcBta6VpDx6TS7xj+Thf8WWg9PJXj9ZtftO/NWlox/bg1i/Zzo
PTCAJvivihQF0HXLdOBVgA2uomTNCDn2jvlFY3wBMis+01KtvpQl0ESc0UscbnDA
DVBRT3foSV79fxZmwb1SPNNmDZYFjCXC6mwUZhnGpHNcoIr/cOhvuqkoqj+iTq1n
D6kGsAMOWt8gGVHTWGfEW/d1a7jm3znTkjrZT8+dpV1c6GTDlZ41JHJAJ+Vpv1+W
8yzWRRhsZOMHrLLnT/O3Rgp+Icv37MB6AUk//ZpFXDeIhg/I1ntuvJs9RVJ2coPv
GcMRQLE2ZmcjkiutHvl9ItB6wgSmoH0ePD+MzUMlZiYWEfNcpvFKcm7jtKq7zAP1
eHtiJbjro4FTQk5yE0xMVul7lH7Ku0OgOxf1K4986MRaQJJwU+RHyWqTVBmRUNGc
L3HfRwQNq6GL+PXfiThCcpxvJjoW/OArfnrm/fOFlaJ8ULGjE82LPbSWqBUqOMB6
wT+r4S3e2mP0UB4u6Vp39XYhmLgr0FYXrgXWCI6p2PirO7zW8gzmVRJ+OS53p7GQ
Gh00F2nt76muS3v/6p5OdTDAdclXXhafCwxn4ALSIv5OXc5QxHcafxGg3DaS0y8s
10S/+Gyl0VG0Im15muSzfN9p7Y3Bk/XjW9gu7fOiKoXuQ9pZ7/Ivy2fHUJ70Mey+
OkYy4Ekjb6O6L+vOrgNrFTnvvN1KW3cfqH6h2cGZq0I0S02KzhtIFd+GB4OX9KPG
TFhE/48WuEXWJXRtSIiY+MmP+dLSi+wYNOzdp4GqNahftZDnKEpv6VD/Kc6eGVbs
PXH4dR1Pg40dsAQuu9itnYuOTlYnwfC8czi8IqDZwiBa88s+iCLmV2+iZZOuThrK
Funmm608+0vdHOk8ruhflk1UaYOUFewRO0jAzuL4z0pJkF8Q5ddnRUDrb6At9M4f
DuE1SdKOcTs+8V//sNHPoUyO/qhJSMqjagAenbtY9kC2/G2hGst8OrCeR1mD61mw
AV/ZeRN1bv6bKQRdfEWd47v47I/2Ayy33rwUTH+dALGsn9abN1yAowjmRovF6Hcd
a86VoqPFziUSkMQ6pUa+p1rhtgc5dSSDZPw+nubvcsgIxuL4doMqElWjJSNximWk
kvJ9cYmHZL1srTiuRUi8UGcDDBfKTCrawBfcIKO9+7xsbG4FKcttgKoxyAvjK0tM
pDtxdEn5He65XH3XA1Yko9aIU0toRL40BwiTbowrknsnN2HcCzbMWYjcQSB7+f63
zCxfyAndgut18bF4zbY+MVabbqxWx/teIxM1iX+VAS8PPTc35s8olbVvkyCRL5RS
uwocwGki3jmHMh8Lx8p2SDZ5hePJ2/XICYJvZwBc5rY6rn/sTywp91vBGQbj5YRK
sVlmggtvb1eiXXcJUjJ2La0ul38sWEi7PqRYOm5m335mr3ZDcm9VTL2mrTrHSpAK
yhXBewAS1Ll6F9UyHUucFJSZjVF7JKCggEwiAVi0LT/Vzer6jXHvCrEw3AMVuqmY
4RMf2TsInA9VW45bevFK7ElVU1vFuN9y73Ryua5u/90=
`protect END_PROTECTED
