`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePK3WMEwgc2U3Lpqc+pI0RKrba3GI8Ox+nc0hV9doBBQ
kSL6y6YzBMrdh8A5eSCA8o3p2tHn7jpbFw2wKUNQCUYv5A33CiB0Gh2DIC+T66pv
i1OGUppeKQ9xW4WO8vhtR8Mq1Z+//F92Qy2iloLksTV6icSKpVYFyWKxntPvk6wy
BZrs2Aw4yE2DWtlDEwF1UZxda8cY9ej+r6aA3VfEbmY33wVyKMVwZSrz7JQrgOV/
kesEYbasupafKKt/KLLes1fa8TuZ+ejI61sZNmW2TG8PR6Dw08mf+yTNbDV6oGj7
0jSa1QeaqQKShdmxhOFUuFy2c6ll8JfNTNqI0W2cKq595Kz9Cx339tR0QN7oLpFK
9Bc7BggB18Dbv4Ke1zAvlqtmULwcM512l+FHuN5Ejt9sjZ46Go3klf+ZJ71q6Lfj
cc69brPKAvDYJ2M8yPv3ouwCNfZ0gKcvuzK7O0pkuV6i1zQ76X6Nk0Lgz8LjjClS
tZJyzV5WBEWSVdxcvIHtzjGwc0mi/scoe5q7U2F7ZvC7BPsIxBQ9iV5TauC66JrL
uMdeTsv4lu17PPck6SKRobrNU1kucXNPS5LcaUFLxvg=
`protect END_PROTECTED
