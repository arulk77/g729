`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SZsQE/WjOc04Iykc/tuY5fbIrysR2Sz1d7xXYfSXpBKz
tmFTt5yut2Qy7A4RbdXsXx1CjrZClTUmO+1WKr7g6OF1RZlbquVMO27NMQsSRlXn
GRrkHdrgEG6cjl56BQZ0QMkWl4AtDCJPb58Vbqhqc1LLLeMiKuNF48AhSlKDj7GC
RWZ9lMdlYRr75JnSK3P/XhjAIPThCet5DpSU4fHM1sfR6fuw2TK4hurxDqYEmUxW
Q+eD6eCb47KhB7jBtdLC0M0okAoX0WO+WHRqXekSX/gbbd3ugn+8rJ2QTSpNgJid
ZJncWg/FfpPYeWHhzrBcXj+b4FiQMdHPBQwvJULftYXoQnFIKpSHuceuYOp3Z6ut
M1EANzU0D6Qn0hHfOBhmpRvfD2774fjW+Vbkjj54DUnqwVl0orResf7D30whiK00
DX/Il3Fjrozb5GY/XKlffFl0z1fBNZdTvjYgJNS4+cjXYaUyTUzfw4N+m2OKkNke
scvj2Vab6dxHoCkmS6uF+dnEJ82XM/RLBHHfBJUQqnsklvAB20XkKzaQBMzVmK7R
vb/wmEcNlQF8gyfOk3Pl2OU4qDQ9O8pBoxErS4Ng949QpxcNd4agsKIoeyv1X1QY
fI5Rq8xDk4qBjJIKB5HLo6Qz4A6eIIE1OB3705TmK4tfD58hqh5/R1DNwp/q4aUo
LY1iAUr95YbJZQba5E/nrD8z44TyrPQIxt+POJdbhK0vAUluAKzT/tUQ2dRAie5f
Q+dq4TpVsrsZnBpHxqnTlhMNx31xDpZBX3O4r3HLzGcW+yvY/4DAnVWA6ID8hON+
bUh/61sQrngQ2p/kqrUH+ea4Zs/wdxk2tQLBHtHe7VWUGTXbWoummojSTtDKLzEn
OzJGzr7+ZDCUXRjXUSRVGfdcNv2d0xWISOf4ToNJHDTz3n/vAVZSDjogiURONezL
0ElpgKARGaxev8pLX128yUOZsqhavWYFOHQWK7cSK2z4NWfAx6Jz9oGHER5RdK9Y
1viihLDzND/MxbtaEfBLayp45Xcdkfup0Am+ahFmwaaBqh+FMBSCcY1jMKS+tqCD
ElHsP8dF13pwEM9/tgTy9JWBbOZ6qqcmmw9C9H8wJ7nWFZP1elEPXX3lgBQYapb8
oRlrJMxMlSN89P0M05F+np5JZQ0N1ZaCDmWxOv4i/NCtfA8JwmogfnKh0HJraYuB
XOX5ELVk7N7ImnytZN23KSZzXi+A8c0cpt3ZuMp++9MCblGkCnA4k0Vun9fZLWtM
NuFlv1TH+3I+gekpUKUK4yIwP+aqyCBwLKmRxFK8s4eueOz99PLhdhELZb8GAjeI
yDzEI1GhUHOJRwbhwIdQLu9b7SvUUJ1MtFc57lIJVSs=
`protect END_PROTECTED
