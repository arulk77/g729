`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44btVEDqGrqROQpuPcD+QUKXzqch9BuT6KXQOgS6eZ3G
8CEs4KmLwFO/+dAj/wIYai5i1K0tTzMtyJDNTsKxq7qJnWB2wtdQKTPr/wvhcPCx
vd/4ndgVvSOlr2z/UxAOUMRI0vDc2dT1jFDQwscmZhhS2eUowSaCu4TMlemk2j02
N3HVpewXa95Q4hQM/0TIiukc6YbF9U3k7aCcuvN1lNVKtkiWTrnYcd8x/lML4lLZ
3XokPFtCZEaMgCnqcrlNaONZdpybShH3gOGWhZDu8DCUpZJx+9eYXNSC1DyDsemJ
/4h4r2COFr5DXzMnUc7qyiS8ha+A7taUE8y8DTqgNXe57wgZ11zejd7iIrnTsihu
eRvWu1cjNaL2MjdUkyc7DHSmndCsfCnOw6Im5ZhSJv8Gp/gFH8OTPCF9SbR9Zm28
KgjzBfbA9WuIEU7A69iKqX29fdarHgdh57+3PizQjvUKyQL6mlmKFpQKk85A5Cmd
j5Jnnm2B17mfwP/5cc6e5apRfAiS1hBAtBo1o8iCpqw3qKW+/eaeaWujZS1njRQF
s4tlQ3qCjMGUcYXewWP6Zfv90GH75QW+acy++zHE582kWPAF9T8XJIFVAey4Seq0
ACY4n9FIWSztb69+N62hNmYdeDPRGzx5dol7x5iGYduIlbcVWNLvVewiVx9xfv33
9XOFqQCoUUwKocgWvHtOtGnYcGTDMDfzIbmuMfsCp6zyIbHYmAFziEvA+yEIfchV
AfrgavCSok8CzaDZFc+oQaMQ65Di72bwd3hBF9Q0wk4upNX7FQlBX9gfa7sTZ4/7
rIi7CK7BknW5Ww2yvPr91SL4pjjsgRrnfgJPPs/Y7OJIS4CFQu2JsaIYzycwwlxa
DAfgZOAaTEP7S8R22mzEskfJLLFn68m1zKLJJfM+6TrzAClTfei2LEEazq2NnbLg
3W7ETqDVouEfs0jh297gEcfr0awj2i7esLr+Uk4QopJVXovPYQW6wf9oVCC+Nifn
YcbO+YQ0IreeHOgoBHRJ37ymV/CCu0r5ZP+9qgN/9BVR65Ua/XJ7P7yGSyNBl6TM
tu69/WLFz6Uhb7tRQULdsD3bgYyf4wquDB+YYBxpPHxjAOkybAzrgxTYj6K0oCvF
H0DvBf1/dFYWPgSjNjpihN6vkh4a/Ep5gzkGJjtjcoFJaAT9mhaXXzHzGklaIdjd
oqU55F02caN5QYLKTZ4KBkDU7JWRtDWTEP87HicVXBeoPopff5zfYS51NNu32Ywd
F9O56eqJBG4W3dQq4YGrhJmqNA/GdyxxD1BalmKxTPjSOnWwEoCWrrgIad+Qc93M
4d1vP+hAPXmlYbo80ZuHoW2YxXLZtDQy6yhjWgtDCAT4OpODotC+qFPJiB/FkJXf
o54HH0JMCehUu0M9b1kIQ/xfsI0YxTC58Srhgc7DjRMutOrSCpWk7nkq5M4OMpTt
wsK06NjIOHE7VCg5GhwXPcHTdarFYSsyiLw6Hcm4YKmaFeYns0HfTYe+Ttx7FGSq
a86RyPjP1UWxQRAot82iN3gMQxd49j66qz/v9GZZvqLB9WfwdySR46Q6L+5HZdTZ
kwujla+3atBC82R7wt+YnGzJLqpII5Z147ApqmK75U6zMOIeb4DjzgPV0IzEfcuw
og3Dqm7/EheWk1Uhol6JrOXSKgX/LPmUMUrT6U869K0+Jgml3rJYXj/FeOQLa4M7
T/YzBy0BuTjxRO4WjDGBH6K+MGD8MWYM00ciuahQrQ8CG0INL1Gm2x7h56COb69S
q+RU2iyGX6hqrK+4gpYUDkVBeQda40OwHfDRP7Zyc/e8DG1spF0acv1LPa2kIUCK
0GL4BZBCXMoqZ6yiJcbdWDzB8fN9VDRmRkaYHrntxvpsztlPwNra5eoN1RPTmmgT
4klHwfUnBbdS+w5K/9gOQfmrgJct2uPt/00y53cN1JIQvFZz4tS58Rv7dFfRnv0n
Z/tayuegogXskb4SNCZOKIKAEdpz5nShmuaomzOC3hZWpbBg4AMaSikPuuNA1nAi
ngb/yTlLYul8uSY6Hny1nGZkd7yi6lq41RhHsbhLbGf1OW9W6uL/aOLB9OtjcZOI
Uqc1zNwIapZYR1YMycz0brIvyRYMub4JN5YaS6AHKx6LyeuARG7klMP2C5Xa1kEh
GDub3+zti39l6BxcdxwF6kcS/KmkYhwW8QgVNAyBhdrD0Tm07gAG6hXm5CqdKV3G
tAMBVschcHNxVcXn3RktJ4g4UMrJcAthkKdxNdZZW7H44/r0cpXKATTgEgxEHDnQ
yvQN0FhBzL1rBh7WwrOCY1XG052czuZvCXiavTW28wF8oIcVumi7/wsse1QZwxle
ah8ug69QKUZgzx15PgiHMF6EiyiGlUdt/9pjfX+IBl3legzI3a4X1nGjBa80y4cU
LdJAqKamW3zYNN92gBlpfEkAft8ejwxaF5ss/d/srX8P180WfZY1CwnKhs0AXzQ6
f2BVlHpKwmRcx2rcB1XBf6Zgbxe0Q4n4Xbd2MmDhIYRMnRkJbjWmraTiz8HpuwM0
T1H0Dg+WzDzrKIgFpz4WbjpunyN90zfLgqWkPaTn7zFAam+C6Jo5+zMO+ytgYAoE
vsWOKIIZ88jLmmMY6QtVvZWX+aUYEs0KMJFsB+FEH0/te+VgAjxwaMKgawfLCSya
YFHX1q0jmI4eG7vqz2QU82hv//6rr743Ga0kp01Esjky8ZPKY7POtxLX31EVDczp
P220sXPM2zN3wStk8WrFzhjKBNjw7AlrW4Qp3OX2Qx1VYQjIi8jtvsUaRqkXlfEY
dpvBYHXzWfJ/Q/5h12+zLqhYMsP+cS0R7wvk+yv8wUs/afam/hT0+7kEpbHJdgyY
SPV9SCv/DOLQT9Bhd/ubUfG3FgxWHk1AKNgpmzH4Z0Ndl9jzqoKYoAExqWgcqeDA
IGIUei6T1q6QdsOjRBnFSkwH15EzL6tN6bIRJ6TxLnjJ/BhuVZjp0gV0utzfYxMt
/fNj6u/5yWwbvp9K6zG8YKE1dDlw/hS39zPhWBnijiZwyu0rK8sdExq3X3AgfFX3
TN2TbuNLcG7tAVl62gxTCSKZy8YtZ1t5qehYmuG7GobDORgH/fJ9590tY8gxRjey
EWxNep86gLHtx+n7vVZaJQYp4Nj4EFxWQYVUfpGZFauDOM2RfSyoKOoZH7mpYe7q
Esm4kRM6wk6LEcO/4zDd1c3RnjwphblfkVHnzKuiPf4iLz3iJEJr4GWx6pdX7/vA
BQAwMlTDQRW4cRNFxCLqK9ZyQHF9WNfdPubwYgyALuXC2fsDwwYj9CrHeJG3s71g
bXvaBBNJfCQeynU3i/42GYLgoEou1EI3KlSHMD7DhpSeKqHLN8/stC5/zlXj6E7a
6tqmRmNrqTLyi/0xMKEJyU3055Afh1I7gCfUwV9tG4ZnL4gN/D4QmWxA5PHgahpa
t0zDurAhzEdhHT8asbwi4efPPTTyjVfI9zbJDShHI6vZTVXOoNul6eqM9tnmuM4U
kyyDTgKybeGVtTWP/ldnPymEZHnTlYadftfRa558HyMjZbCn7b0sNqjyu1zl+XV3
cqFAGlxL9K4CZSoy9lWxMB2+Co//HsdObZBZGXCLn06WziE4p/dfYLHE64HZw9Nv
ExYUsklxgQou75y6EJqsj2+p3fJ9tvvk2R25j+fesRaGuCTuFaM4MjRMmxbk/bGS
/1EYdqkoMZoXaypjk0QapED16eFTDCEGHLs0jiFe1ddTmFGgPBAoeVfRS3/PE+NS
PdDM3Fue0sqvYqscTEaTpjx7FL81CALfXSClPd5SHXAz1hoylCDiX+87j7H93PAD
XdASJfqVwZZx3DoRh9aHx17vKj1jzIUREmUHT+hEzVOfCFUDQv4HcukgSKNstnR+
Qg/yQ9WLn/sW/Xq0mF58QWKMzs3aA6ViGe04GTo70xj4LmTyolle7vR/7eGEv34P
FOoLzF9TbMt6lUAEtDst6FvjIKmdTLSpy7vNfXi2Ui9oL7oUNcaBaxY3EkvmJA/F
2gcQuKr1ll/ZDMimhIwV8WpYKsvmU0d6RnBiqOuxPjU=
`protect END_PROTECTED
