`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePiSpHTJCGZGfd6iOz/b9LismW0acMjwRY8K8Zq2d4Cx
BjOtxFdqxzZRqWrxtHquMdwnaLD/HO9zSGPDGsvmMPz6KNoZNmR0RR6KGokvlt2W
cLVW70S7Du9VE57wFt04HH4ockwuYcI2SNZVGJ1ZFd7bP0l1qp/jGQL/jjOLKmJN
XF9+XQfIgFe+9h9b0TL5oXpCisFt65RlTTNSd7mqsSvIdFfunjvSR4N9DK3JM30m
pTspVMZba1Zbagl7+WyTs9jK7TbvAnLr2/Bm2T6cDX7F9bsMGmmoJTZdmauVkMTx
YoOiDNJNpbqcHVWiY13irdF/awvG1hmOt06DLZxLOGsVzDPvcc2sQJzhSxvEx9wX
`protect END_PROTECTED
