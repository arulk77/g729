`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42pErQB0eMuFTruosyt4KgPkP5/8Did1NPquLEPhO0YO
PXDM4khBTgRSEy/mG0EdK35u79k4MKPJ50PW71YfP7Li8u0i+SHe5IHiyXiSp66m
oy3sRmgum4soO9JGDkPm0wzIx0HW8LIE7ogLYm27r7zNgZLiGvUGq8q0ZPVI85H+
yS5+LGVJyVHeWw7UmXi7Cdj4p29UBg6iTvmTyW8PQ2sFJ6lU6Sq9JVmyIDK8veVd
s0Zz5rNoHPr693zlHkiZmi+KEj2pXHLGrNiEt3wgZaRtKg0LY5emSdZfG57EfVEP
uDdDS2E5QMG4bQK5M53HN19+u48kEkqH07y+MDOFFKuBXBRPDlz4V0Ry6okeesbG
MhfIw04CShVm60SRRvxlVw==
`protect END_PROTECTED
