`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOfRXF3gMTSZNqzis6i/1jrf9e7Q4++wJjw7cmKVietG
kXB1dE/rWR2oZtaFrlXsBNTUb6u5r1Txe1bpmPOcoyCHYqokNuvWiHFEBNMdfeON
1AwYT8pyGCzxIZN377epRiZEuBVVM209hyIDCRndZNofp65EWF72iN/HU3d4G7kx
vugbPGlgUXuqG7cm4XWtvE9XFdbv7vuVnxstLaPToypUT9zO5zQt4wZ3uknjgffV
9SzZ3DO6y5kEdpodNx/FY1ug9OtFOGKN4JWl+obHfHI/SoYXTnH5W1TUL8nPkn3X
syet5D9gNyblIPouW+mG62HJolVh9+nKeHlToQ7DXOcaBZbCSLR4gFNKjsZlb5MI
odz4kimzCAXlyfCwqK8Cbn6HGopiIJ/QE8P72A8JqWC8KynyGT2Y+TKX881fq/CY
HTtp5PvkvAHulJiSvGk+6RlYU5nL4QFd2MbfJU9MPwGQ9nPg+USkJYSXmmuwMtCs
`protect END_PROTECTED
