`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveInvC45caTTxTUwFx47zoshZQSn5bMtSViQDQVY7r9fr
LhIjkDD8jfTV5YpoMy+Tcxsoc4a7nDmWUgCIVV6r4ROqhRqT4wOMHvwFkpPPrC5q
g51WJ/cJbg1kbcjt+4/Eum0yrDlfjDAl58Bt+IqKJZbreDWexMaERBLUS+mhH9e2
Bq8PT7FND8vSBmC0nC+Hhw==
`protect END_PROTECTED
