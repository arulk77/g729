`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCxTwgz6Iry2MKBq1Mo3obZDVJyHZdMuX+D/rxYTr9Sn
OYB24cEvKR4M+pOEMe0sg0up3cjRzQAyqmXF3bU4CAJW4jFjsTU5x+cDb7/gFfRu
tyHuZOzBZ4YZesxm86ssHwhnc+78zyNHtgaVwadsBQ0IW19YMVQVwPNv+1/i9l7E
6dN4rJY7z3x6rvR9fXQakqmLSf96fmPNiZMUENcuArCWYbd+l9v+G64HXHa7o5dE
JhuWD/9xzdH3f5W0jCct3H25aG48b1/9MnxYFrm0BpyUo+ZvmdlyC4xifsCakBv+
9sZRtAwo8LnDEQ+YulIPzgtYFk80BIl6xQ6tFcmfe1VefcnS8YL8gQ0G3axiwNd0
5zBp+fQf0vTlR0hu3isu3g==
`protect END_PROTECTED
