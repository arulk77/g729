`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4Hjqyl6wc6zZGR//pfxR/9JWTAikI8KW1qMg2bggZkER8IIFhfJmfs7v/fYZemrj
GjVuogTqLDc/jB5zZOAPMTwlHH/OsRwUHRqzUAzfCk5GL/PlVGh5OHqB5hSqNnVQ
q7IL1TPRg92aOo5cGM1LLV2xI8pTkLDKgXOJ6RE3QQO1m1IZKgzUyTQdJY4p/Fj+
BrFahcc0DKXuH9UjpgiJIB4tvE2sSu8MDkiu3aQ8GkuVjli8VcPVlG4p87bPhRxI
38aGFW770XATztLQmX8TGUOojh4tKYnUrUPzMMxuapitRQ1iWRgoUJCEcP0efHuC
TT8gaZ8x5XISGAqsfYcV+XuTgTflcmLdHPX+DNmnUazN7ckiJd9oR/cUK0Gsre/Q
zSrffcT93ewdkUsnVSJoAZOgZd2H+/PvPT/RL85FfCd5ShbbWpkz2+a63jAOZf2i
He6vjykb8LTnn0geKimkIWDgU4q3JvB/Es8zRXoacRGQR0BtxLv526crje19sOyy
hgfpHsu3bvmjcT94El/zs6E7LejZPhUxjtDM7cYNchtJ2EDJ33CICQaPDho6vpyM
MOF35AMkPdzeMVhEYUy74hxFyOawEp99kJTPH7O70aizZr3w4tJ1NGS7jc2GR4JA
mKtskBiSdL1YCKkgisnKDzHGzVQ+VyeS8HNZYrJOxEvvP00Kbr94n/vFB7vg6hi7
wtNApunRNzXq2iMnOXr3G03APunMU6E2aUR6LUBXQnBohvu2cxQSjcmOo2DCJ9Dv
`protect END_PROTECTED
