`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8Sel1g44Gdw2fNrQKP1Mve89CDkqccd2rGT0qj29CMkHm
iBU18A1Sl9K+SAndaIPeLaXF8HVItyBLRZH0uFqXINy06FkxGNbHEM/cMsvEen4b
+NlIAKzrsPKzpM/R1yZ8f/rAutd+IUj5wc98/hM46eH4i/KijUpDBEkSMjspDtOV
DOFx3k0BXC4ueL0/F2qXNJDJP1BIK3x+2Ir1MXtdNEPXJqRGBrvlRasTMhqYYOJ2
sEddFewdJpLDzd1gIiZSl5e5x1U/tpslpHD+0pHYfDrmrxlIy0xEEAz5WnG2ah7t
9z6gcjvFWNSxeZ1nro2qOO4dUxMlTrIanhpR1nWqCPQq4zQQIJd0POakdoEbI0rC
Rp7Vp2QX10VLPzpP4g2yA58De2fcFF4zcAcsOFyMRTJFMGjUzYs55yY86tt5wTwk
m3biEHu2a6JyDP62Ku6+HhRev4fIeFTFSIuOc1+xWXoOYPwCB67zZBG3Br8zoDxI
9P51k/wye9OuKGIgxrug7+WuifbhH1iGCSnPAkMC2r+B4ZvCc4oPfttCwfI1nWzA
SIkfM5FhweyPKe5gMsqmeWK8D6MfXmvX35U2O4+ZqG8CDO8ibme17lvmAY6bFy6V
QZxyYIsKsxkD7bsGCBLHQ5WvXvo1/T+WvIHhRVVoN+ZrLhhpJ8uA4N2CkrHUe6+o
2s7NwwtXyO2i5ZrI3DjNSLRNx2kSSFYoNKGQqKSYvMSFILwOSn4Aga8wv3/GZ2ct
Yx5Js4ZH+/GZFlqHqD67PmVx/QqphdlTeCfARKS6U3oglikkBCTcUQq5jBTNpVME
XcHPA0yHtFFedf9fD2i/IWZt5MYI8BT7sZ15+XxEfNqv2kektlsJA16loMZyAMAM
FvnBZF7AAjgOKH4n/Km03Wepzm0i/jI2qoEQDACBy2LfOD7FESfGpxT5AxnokOzW
A8ASdBIF67tpS7hK++Grm7ZBZYM42HB14r8wr9kbzF/IpVF6nZpLkMWhnNLjw0gH
cPSlprktLzUxe56G+d3UHHXSihWVXzcAlxwmPNEo7Pp6SswWrCQ3i5hihtHxw6+7
MfP3yuw6cL9ccP3cLPZ6YMdNbEp+XhPPXs69+pxY88qnna+yZWKHIa3n4onIEbji
nrf0NfEiUiywNJWO7b36de92WlqDS863WaSB4Gzex/H3HyNg+Jrxi0CYIerHJzTB
riH3tFpW0hSZXPHy+h194jfOF6sBOiQ6LmKZSLaW4J/HCySczl2q3q0sRnwk5tAR
clr8MIZWhimV1+TgL6amGLOL7Pz0ZEaotWa9I/x5/HZRwKsP1mv0JVkSwZwHN5/d
IFQwXHYYgHMfKxadV/3ZxjV8FIxLT45/fIsh/Lu+YKzgPfOR5jxJsXud4mmipMNF
Lo62sE/LMCtXlJet9JG8M7U74+CX2ig/JwNuxN58WeOJEDXh6NactKapcQx0XJXa
s05sp7uHv6ITpodEHsTM+wgFluhRyspDGtyvOigMPxyPo+4rrShjg0QaVlpJRQAD
1aToWCMEzNHHt0MZyo8Rmw==
`protect END_PROTECTED
