`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wwXcoVrRjZ6Sat+f662XKGquO3NaLCc4gjuD0/QNxk2
yxbmgvsmow5lSYnLqt1txB3dY/hkK4F2H4FYcfyyhaNjmDJ/qpdW70aOSJO4nTKq
6Y3upq43JEQczwksRcI2EU0oQC9xAqhawl4vEPqwM8jgr/ObKchfu9fcFIGCvqoH
Jm8GMMmqwLrJ2MjfydrPxmDfmUDrfBYAVaiSBf+fbeGCe5uFpzj4JVlBAak2qrOr
qPLoH6L6qAq8RzhayaWm+o7QCHAMmm1OmD5l7nT4dDk=
`protect END_PROTECTED
