`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
iMh+7y8FTLUC4g2n/ugwSSnt5okHMeebMnZEf9Yja0vSIl33YUOPfsFFV75GFKyH
ld+zCxJDX/ppKKku+MlmOk0T8Z299eOiFh2VF2X5h+bCxqOIxO6TtxyFoAsvUeGr
NH5UEIwqa0Z556V52WCsUd2pX9F14X12cTxVVTlJ3GSwD1O6t+fNsKaakf50Dy8L
D/v49j06d9EM8gXs/LECBeI+BIKNXjs+7Am0hfWozeaSnkjnaTcTEFyDdHLraH/f
+vd7G5pA8/nPcuU0XvY0sOiHvz8RWz9pB6wBj4YkyOCDWaIlLRPBLqMAWjut+L9g
1CXqyWMspYRoe5RcdtdJsaNb1FuaZt5Xat2eVXLYRTB+nevcFsj3+6jCT7gJ8QUf
28S5fFWoJPmj7gi8G6Fy3Z7fnhtA4rP6aGVN1VrTkR+fz/eMGj2dSv6yew2jLWGf
vxEyGpYDeStVm74eZBYqUjntVm5JamMLvR+yJWo36Hn4O9V5dL6HkJIkGJD0HEZo
5EbogfKxkbDjQ8gyNXkgJrcfvVgzQsTjOoZjLnPkTphJ66p61LLWpc56Fso/ft5O
EniSM0Vx/KvE1i2ZwDmzttDyWStIiy69/wNcCEHeNlnfIlwOyasAWAq8vzXthTYv
xmt+V+LOZDHnSjlI7rxQ2XsJMmlvf49dSC1/SXqeV+gwad3T11q5XJ3B+CpnLSnQ
MVqouPU3c4K27enI2Ak2mdoj1l0NYl//IwHSaHSywd6d4GPKt0n6YLKzfg1PbLVP
2nlxhgjXwm+UEAtM6keMnoOMtUh0HzJgntPiV4DF37Ftj7BGeXw3z9d8l74LbXpG
DoAuM1cLZkaet0OmbjVKNaGLYdI7Y5ekhLLoHMihbAY18MaRDdEyP9BEzWFo8m7b
gGmhLICV6rNVvlMxYoCVfww7idZ9FOBFon+8EoPvPGde9Kz8F0Oyh+NMg9r9R/78
wVkX/aCRxautAQkh8GWEK3LeZ/kI939nE0Rqdh2Z9ddcWyKS3gYAEu6lBHuKAbST
IzDvSsCjUw8Wi2AkvJeprgfBIDMACVbpDr/gmqf+m5U37oHz8YH0WzmWj6sSoV0J
D5FYT2hawsYIiBkUpNnZBBFoGfgZ3+s8w5JraR6MJnCaYOhLnsHaQZEKwuxRY1Wa
VksPryHvyq8ZCirQUaC+mG30UmyTbLlPRrfwyQ6LWNRvgSCGGLEjSwzb+OUm7wKd
nP24dqCPwXdMgbWJn4qsEupYTcchX5OtgzzsOmmblNL8L3yV8qfqJHG2Z3m68WgL
c4VV7OoijUIbtscwabwsiFmXZXA53wb5axfHea/ZGYnc/23gSEvTzUYbSsx0l4+x
H2UQ1p02yagWVo8eTPnrdOqwqo0tuu/Tac/fs08aWYDbTrRoqASz8lryL04eMY3L
J5PeB8NVqP2miiqu7AcMvvnd6VE/tKZxgE2gmG4c+w3Qea2NK9LlJGKQz7z34LfH
7pgS7jaylkpzfw7A5f/1xl3FYcE3KYcqRqdBcdvThh68PJG4s7P0NJR0ZfZEvBDt
6GA5pYjnZyjkMaGAvApoOVvatx1weWmwDXkdiyhxFbWzfPvjML/Gdf8YBUT9Td/d
DVuuIQnZuvT8eb2xby4AfHacosZY2yWwXycvwD4Wp/MI2hDv1t4YResC4b6vBqte
aZibmRkG/oxWE/H2pY8K5md4RbplyePpIokImY3+XYIKtVQmqFv5o/822wVTmIwY
NapJxLD9hcj0l3Dibhio6rrBVBEZBnD8I3sZpcY+UlkUlJdER9CFmYZONpBqdDGQ
1gZcOSZcWR62Y0c9RNOiiNJVpQwQpjuWhIJXE5cVaU5C5prId3Ks+DcwSqmKIAwH
gRbIHXiypOhZSJOBjZmZL9Tg8Vr8lXP6CpqBtMim65YF3/14r095lAIUxd98kaAA
MSng7aKtQbiC/grb0EQIbL/7UQaCGsBU0jjj2qZREGCZy8EqYAMn5gTnSocvTW8s
d/ssfbUK/EQIAeD8JRB1bw==
`protect END_PROTECTED
