`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDMMnSGpGZZ2/xH0OJDHsSJzOvjeuudxyZalv0UO7kgW
g+D+rQbgHMzI73x8ypW0FzpDjY+v7DkWivC2GwLqL18o2GEhQrks/GJJTPC3Kop/
o/iZPUZMDlt72V/GjeOoSRTDobDNJwQrXZFbmEKIBhLCi5ZklZ9ULZfB37y0PZM7
hf8ocZNsMSNIt4wppM7xaw==
`protect END_PROTECTED
