`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK2om1PLy52DftjMFaaW9QuUdruy9hSQWkBGkhXAB7Bj
X/AI301Vfeocs2J/mYza1tySl9GvzcQGLwvcZOm+Mo+EN/YL1EiQTZNcrCfOIw8f
EL1ot2BYKY+tvJXQgzsTrjj7APNxJvyUojXZCAE+Ei8J5MawbP2pIYXeqn+bUZDV
akjD9Fhghim+H8qjF5dDQw==
`protect END_PROTECTED
