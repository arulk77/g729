`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47NoBuOoYppqEnzegPPtacJi/CurbIfLmt5mvmKd3UnG
Gs3vwqEZUskLnMUSWdxJNvVNsMXngogIqlJ61DIV/hfyGG+5YVfx0zKkTO/86cqm
e3bbrB/V3e8YQLxiKCbm1W32e6wWUpe7kRvLfeAna40RAFEJD2rvxRyA3jj/+i2/
oUz0cb3GK0u+u9tfMV6w7hy9rvQo0jIieB0c8SddTeY=
`protect END_PROTECTED
