`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLyWpNm/MTEICefzcJDbpdzPxCK2fy4CX+4NOE+cMVs5
0hPNcCoLKW/XOP1G91DO1CZXTf7bKtIR/rwVt2+x44jwN3zD1DiYXK8PS3Fi8pAG
kPfIKUsWz9NkTar5/G07D+1t+3AqLkwe14h/7vj2Z4oEqnKH2SrIWAY3mYd8bnKT
KWiaY+X2WTbie2AK5ffUCo4tmy6hcUMeBVUdfm5R7sbluH0zT/tkEgAWxQT3IKJ6
cPBnR00Zr5R1uhq7HI5+sPvffpPnLxd7swfGhkHnix4p1m/X8h4pB7f9HpYQHjZi
QWufCAas4bKifr8tTNetIJrqWaaq0idHMPd1Lq+JnsBh/MJd7hbk25GbQhsP69C3
wcN0q3zEGciBytgYQIP2WI8Ta1QT5CFewU/JsZCkFL0DTFqMvCg9AdN+g/wKw0Wi
bKeA8Swkw2lgSW3tPrvNqFWI/hWLhgEw0Ew3KEoIgMWNIbPkikvlFkWyEa9/biJe
BE8ijEXsCFUpl+K4bd1M0D/jNKH4etMJNA5KnCHFiBaME/JfeLlokshglU4PZJAg
`protect END_PROTECTED
