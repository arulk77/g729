`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47FVyFEMewOhonNg4IKS+txnOKZHdtDiEYbboIcz5TNP
hvlrS1sFQeJY+I4LmIQjW1vxXMLLI6VPgVJ8M6q0+w8bFeo0+g6dAREEM6521+Ye
HHeq1H8Meb0GKyKmowrqt73wz4g4Nqs9d9eFeOKn+6O0YE285Gci1AJDl6nqWj0u
pyHejVbokkig/qDZ8lTfiHPFMsyeyrABvrFTmindOyMTF01/eKhS25+P6HDB0T5q
4kWFx2GZwKfC2eHOLw07MDl4UZAkC/rEnszNqXz8ffCmV6NYAJeHDEPb/5oXmbON
CnpFBELCVEOqogKgwUB9zA==
`protect END_PROTECTED
