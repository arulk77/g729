`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB9WFV5gaTlELAQN6+SLhZQhZw84etuH8SgTEIdipApi
6yqSCHvMJpXSK55/AR0mefStELbbbMzyofXpShnp8//UWQuKVJ26rBkWuhe+7D71
aCnJv7fEYQxF494tXMhuhBmYm+66jhIxOM/sjC70GDGKjHxGr87wOg2ki/hZGF6s
GA8dAdx+rc3Di4EUNiNB9Q==
`protect END_PROTECTED
