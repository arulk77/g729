`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
sc4IqbKZAd5Xbsc/plXQl5B3p6pGg29fhV2Axs3jXDJfGIbqnsSMco9mbXBHyYV/
Kel+Uw39qwhQxgJvKG2flkZicUge6Ue0MPI/DjeaR92dqNIvghxw+F30928VYktB
xqa2BTP2waHJFxlnFx9pRGejjD81mRVhAFFz/YLrFRPjsMr/tkDa+dLxn4nB2K+I
3SnuYnoManWY+zlowXde6ARKv5oQfTKHcb06YMuzz1IsCKDNHdrM9oJNnTk9LaNp
70XS4Vzb+kyEIE9l9fBvplxn4P1ZTbi/w8I+/ZJE0/s=
`protect END_PROTECTED
