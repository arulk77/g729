`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42YWMaYCg+9BD5CrQQNfHwJDaSAi5PJJ5b80wjNEVj3I
JV/cFmAqfOChLcbJYA57QKeXeF7TswST9XYjvb6drKBz61swuofinpPtCOSuoee8
+MH9JYxfC7AxiL6/MGTcQKIK3Aea2WwWHMS93dL8ELIHRJAo1s+neRD5pk1nPt5R
xZchevmbiG1T/P6ssN1Els6uG0tQNhxO8O7UQtld8vHaUNJIe8OjF3V0C1e0eqsb
K4e9x6MmTA8Dl56N6aSuabFtG7aAFSp/i8+xEPTPwqxf53Xz0rPkvaUMohxFdjXA
HFYtQTdv4D6J/WaLUsifiUiUsTKBlbtmBABube0MhBujZT0oeRjG7VTU2s6pGgL9
Ao4+l3i4Uzv43io1HsnJqA==
`protect END_PROTECTED
