`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGrHfou6lszZyR0YjjTrWksd21L3a26qM717Hj2eXb89
3hKSoQ19UaNpXK4vnKLN+G3lSioWEwQwGyipHTxwn61Qx+JfnlK0V1HylgLTIEc7
CEjI/ZRvCOqCsJCB9MGq6K7trzHABKrVl+OrE6fuQ7ZurxeUi/1jpAJSQtXijShs
fJ+xhiqqhsBsCUArYb2GE8BVzEIgpr2yvXZSG7FrgDoNXXgvOBdyX9NioMQykN1b
`protect END_PROTECTED
