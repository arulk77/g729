`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
elWc5eeGjAl0pKPj1kSh4T4aon917ao6dxudYE5hdGrhnbUZlZPdsbn/Pli495n8
bL1CQzHnvjS0KY1DCIfpr5oM67G1CSidoMkcmIJUQK0nqVdimiRxTkZ4kLpVVNI5
Glqk3aC1ZW/aDNDFmrx74s4qbTbIybhR5DbGVAE9I5Nd1KbuD50x7gn0PSK5OWse
`protect END_PROTECTED
