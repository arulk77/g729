`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCEzNzbAuVNtM/h6HslrH4+BDDbS5xFO4T56xW52Opya
jT5VgwQ4zepHvsNmXWSMA1HUbLczdmsXDst2ZKQ5StyQFjAESQhwnMOOH5eeaLUw
5epI92WIu9sMYkAmXeaPB0PIsLU5I02/7DENu34nZ0MOQPO689CCL1wsOrxrh4UU
NM5EjugcY4kEfrqcKPh664xW0mPGm3HAXnauBu1TDf4hSVmRv4Ua0fZTAeUK3fFL
5BEsMiKYyYtC9feDotmzuqUu8ukuPeISyID0Ji+y9xd1CG1OAQO7N9SCYals1h+I
J8eynHb3mQxtbcHwFfytAsWRwHf21G1gSvrVkeYR9z+0Rfvghi1jjwrwbDmUzmMq
WOCkRnTvZCxsVeY2rMSIZA+KX9cky1Ubn9ZiHWphPTCHzSqVLoGFC5+nIRVMfzNx
BP6K3++tSo+iYmTQpS0/zYjuN3v/POIyzQoudouazsZKxASk1HpwgV16TF7ea+FU
Za4ULr1TPCb+RMsU1z7DAab1S0e5VWeit88Mj0X6M157CwhXWNpY8OIOTVCKpOkx
`protect END_PROTECTED
