`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
SOy8zRQkPnGeDazAjJk3PPJWe0Zq81uh+tx+eDrwCIa60weTnWmy1o5RTzfgeR63
wkxW+thmL2UnbpJjGOL9IJCHdrof/BUs6utaqWy4TDN7UWvhFxO0HsBhWwnnQBB1
XRhexrvgBsgqEgxfjS0/5INZjhDY5FLaeFfwVNUxpRYYVejEmqn9YHmohu64a555
NBZVIfV6/hvCexMB4K2K5I1hHiTBdRfzQqg+0p4hjKgq7BV4CDtgvzKTJJJV9k5M
0reDEGAkhS+WXVkoUOye8+im2VnjrMTBhzEl5tMv3ZWwhizr9XlgLUAp1JUTBJtN
h2Cgb9vAYP/KXmm8VdF4/oxa0o/B+DAg4RGg4YcGsE3O91LExOiupigMKKwhiIgU
y7LVOmT82eDtkgxcarISx3+QAnfuuyYJt5SO62VdTilFpa4amsZXGhrP1hNKWczd
Fm7oWYOR6psuV6CtnkT5QS5xwb0fKNcLI+iSB7D/4d0M9UK9Ae+X+3svOTOUT6oJ
8WlAHiRDTnu8JXCDCz8AJS0tEIk3F42XOf8SzglAumZCmwail7PbgVrStNKdR6Ng
iOKXG8+F32i7pybO7TlvM4Q91Tg374GCD3mAZK7Cr8kP1hbRaxJn+mz73ba/MUhO
f6EFsVCwCQ39xyUQwz9h18FO+UWPZ11xGNHmhrg+4DAJqxe7cuuZtp4/fvFSfodQ
K6K5dCvRoVNFQqUs2r8eBgUM3JTVCPlkGCC544yveNUvWsIjg5ZCxBpLgwZCAYdJ
`protect END_PROTECTED
