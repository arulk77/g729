`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEW/C1RQLq8pnF1qUl/V97HdvYc04F2yVs3HiIaVQTlz
3Js7XVU25LMTxlC9OKXzpqWdSMxmh+wKNco3PBd5YOrPrji92/aW4adq76PWf+ik
SjeUb/0FuPd4qK1IDVEn9lYYo11fKuXHT75b2AsFw/7m4i2An4N7KRgiKgXA/DCG
+zX0lQqRjc27qa3UxFWBPx1CKqkLv4ZoVJB4vD46QyMzq6PLFq9iInHqPUytdaEt
`protect END_PROTECTED
