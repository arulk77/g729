`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKUKLa/1dSryMo6CwGxBDvDLSGp9ay5kDbCKjieGfIrl
Mk8qNXMi3tVTU59eyjP8qr8+7Ymi0XyISHybngt4hnddLjvA9Tc6NG3g3mjzbRuF
XbEfKFZzOmN7qZ21Ct/QSw+aju6hJ/iIFuCor4k3Xh+mJP84uVhSVPm2qpLwUO1Y
gqcdRFbncvsePWWotTFaCZj+tSxqkYvuOb+yLb3FKdLVMgjfdwU3PcuEy43SucFt
Ew7Mf9wHogxUjD7IqfVGHWVhZK7ayxUh6fra7DktAw3HnP/pFRfao2eDNcX8F3+y
mrFChx0yAY/+zKZwqtZTM0rIBSbQDh+pTAESZRJYCwrIEUBlRiUB4G63AbhPzCib
IPIW5NoE0YB+iEkH3s0M9A==
`protect END_PROTECTED
