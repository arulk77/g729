`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGqc1OOHlMue/L1SH3ovJc3VTMSEFpcoMUSIE5KLLOsG
Ovy5M32aKFs/lbnwMCqYXRmRx/+C/ok7RC0MsqrwPo3hkHMy4l1sQqlnOgPgVJr+
6hJsuvPzsLgRqCNjA+eDppZrwqlBD4GqO+fQ33Z8K6HTZpxukmK0eSxiS+LBSW6O
XhUjg3mgA0WUf4gwjzgs+oDVXNgAm7Op7d12Vi0ks9aAkBti/eRlffKKbppn7hzb
zl37m68SSc1OdC/QmBuhrUTtlSrMNpV1IrVJpBzFNEk0X51stdlLGmncG+kx2Ka3
ksD+Xf66MoKvpBt7QsfWjgqzwTQP1bXV9AlO4ax6OsFwR/SzWWlaYMoPR1EQ5+Yv
ni94f0lUOWHKYnyHZCuQ81j/AAlTO/+iDOQHrZPDGiihwNfAdVBPl85O1dhG4Sb1
+Dfwtj4YyypowCiIY4FrKGyMOUQCJQARLaZSvT+7JcRLwMQ0XMSgB5QEAGzBdJig
`protect END_PROTECTED
