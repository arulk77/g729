`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK0jMSY0ymeCopG/D0WABe8CzxuoZx3It3zAkX+43/I2
0KIFXpa941FnYL3nymYvZC6rahv4bfcaMiKwVDnOfMyfkvFocxgPVs2SstquFi/9
/+Q0SELy80IulB4gpRe/ns6+mqoe1M5ztbyBG3yO2x4yvXsUDQQt2xuXreNDCbsR
kj5Jaqqj2mR3MWgFwGEyzuMPYMJiuNbilM1vDTaO1YI/ZEH8i2XYpKfHU4Jklx1c
AglhfkVx1gaOECDDJVkJY5aEg0OR9V+6EuMr3iuYRBMqkzO6Ay/Gf4jaGsgVJtKI
FojFob1oTk2uLrQSyESdbFV2jOTYGHsh7RZ0EJ9xk67JEKSGRW6ADabK3I4U05PN
PjvGnKvwMW733h4rZKOvUCxFSnx7VugW8hSTlA9h/FgbSi/m8mE3sOh/p8UB93if
ApR8NAHWOmkH5tue9YwRYQoS97aMpB46U+GBW/477dA+hSXQReF0xCtxO948m0I9
`protect END_PROTECTED
