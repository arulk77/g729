`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aSE8n/nhjHsO/RRjAStb8Wsog1+ooPMiz8nTfmP1r3+6
ffD2E8hr8SBae0Feii/1UMl0oT+iSTdGRMNSVcoS9w4yzrhsNyvdrGEv0rpbZHyo
Qluql3/Q/l9eCN//dZZwpU4zk78HLU971K1zjovCk4ItWwlHizdtweWq/449iZnL
NkRnL6mU2ufiPPwNMSefS1N5qRdgGV+CxGrwiHCb/6itzF74oPWuTE0OaECJqy+c
CAIg1vVK0/OsE/GrQPsC4uAIII4dyfYs6SLoSPuGX+vzNHNEmkZ0NYSCWShbiCll
RwlQh33Ny6WZb26ZIDMi/XpjE5bGjBFubgG/DUfJFRM0oLhm8FSWsVjVETQaU/X0
r6wU8JFe4G0G99TR9M6MgvqE+w+GwnGNNff/pJRygJDLZk8wQpipppQUUbG1fuVv
E+bf4Tv/9GGXy8zm5mxmzX+WuBwNcFNviKzrU+FM8ah7ahl3Py/RDBzCgSPVz416
glRUW+bLSmSfImYrUhkv5zUlm3e79jzdK4377cmmRr0zuaw3frTK4tBVHmWBO3Pw
CpONN4Nm0XL4bX8YqjEnGcSRorUytiCAyu8sBfn8JBqQgPYzX0TbxWf7q59ZoLRR
ut8t17iQm09th65gL5tEVsJido+AzZKWU49csTC81BJ8c5cgINQZViDLhpwuzSSO
82JWv+wuIJCYFe9tW2VHIpAk2N7Erku7dBFSG8YwNTA7fAhX8emL/hKARXaHdUTY
Fq3UcgorMnJP7Ct27iWwSl2kMyF0wVkEba5ZjRspmXzrHm/aQesyFBq0m5Axxc8D
0HbqT3vHYGOaTtzuOq7JkiT6/NIwe5rSMNTxaWwyDb1Go0RK90zif77EPx6Wh1a6
PoBH/aghGeJ8u5pFqiO58zjbofTbxEd3ySI5EDKJcM/8cPWz1Qgt8AVtZMSPrMg5
23SoTsvQzmqnA8ZbHdCQHr2mkQ7kJd7WVznI7V/KaScMzwo0CyNGq9frJeJrxSlM
trH2GsFnSjpOVe7sKQ/dNPxNZOGezyL0TJam2odw0Yz9OZjPOV2WbrXiv642zD+f
n7sdR3HMscovOwLhG/8uofhEwEeJf5tdIw7iNm9aJU4lI2MY7zYIAsptsqud+Tku
RDaR2byf+0NOr1e5n+SRbdCQgfArPGvux2ji0CO2q6Y=
`protect END_PROTECTED
