`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
36A/U5tO69wVl401zVMLLSMkyyZz7UahWM5yi3hu9xGoyR5dNCo94yI17o1XJYPx
jqnI/xVefFjzyftqeg+szygGNbGOunl4owEgqrKSEdP0eCluyIWVFdWzQMcjGSTG
txSv5FY3AlwFcruhDbvTx/wmYsO/2kpyS6B9a57QuFidKbOoq3suAw/ZhUccuJ4H
tZpng8kkJyAUf//RuOlNNHDfyZZmhu2ZVQGDkgiJgkDkY9tlqsGwmCiEHudMkW9G
/keoZcIjAJY5rLixc3QX+Htem3HAUiBbuPeQS5xJBKxGdwCJkIlyjtFmqGELxF9W
tk4UG1IWnP0XOGDzO8ZWOZSxw2Ev9jfGXyI7rV5sF7WQ+KgW1IH4iUOauJoPnllO
`protect END_PROTECTED
