`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKaW9FjbK5UYHlhjqvSK3WiDV0j7az7rhRknyamKTKS9
+h0eRcD6PcIIUrseE5z507kZRqY46zKNJnzO6HuvGpQzGabZ55DVHr+hzMPPPLBq
xdxcbR1msa6FAHlirsmj2xPP16GoxzUwUmou9Rwq7OkNFWMnwLO74RmqqidZbJg1
AY/I4c+dn1g3eRiPQDkJRCvBnWdgfjirBSW8S0OrNLwV3whmfwXDQyI9CTBciuFf
Ye+43VwXYgGXNQdE6kOTtw==
`protect END_PROTECTED
