`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAfnOmsYp/a7QowZO3apCrrOWQjPNdX9HbfLyXRUUGGz7
3UBskjPByDa503GoSlIa2v71kbT1QUF7yuicGjSXh1oIkcQ1Ib7Y42EaVnWXMX9C
GZ2kCoFkEwD/ZW6HXeiNB5WBCqaOAJBkYwrK2kuW34204d50670d6L/bMvb5+9IY
CAXChTGeqe0wIVmAHXNAfGV+/eVIVG1Yu2MYs4D2FiDPK1iadzsTZ8z9R6I21VT6
l5OcjC5v0bmBtq0RpcZ2+CXvu/K5dJkp66FxNpbdw6w2lqwoEhODRckgSHTbRXbo
+54RIpqQKBOfFg2BP0PcFeAaoBc5j9HWd4CDetkbSgst8EAXzQIAX3edhtHoJiQH
S8QsWFxobP/xs0FgjHD+il2C3WKW5L2sxnFQrkhW33A9kVCiIk2AqnJe41JEFyUF
AJybcOqFU19QYM3IsPaG/VdU00viZ3GI3gGEFLj9VM8N6QR6hY7yi1xy6C/U7DcZ
nPXq3GHfZ+Xsqv9zeJO5mbTUXhs2zsoLYI6pOxIJj4IueDO9/H4XkPnXS4esyRwC
1FKk/pmUjAn28QkftAKNveXV/J3e1xR0GBiENGo1fdJ+as0cAVtCLMMU2nd1sWOk
dVC+u76JgWRrYUY/Egt3QCSt9T/qlTrEHgq/L2cPw1hX46+lTBwx27vOok1nSn1D
Aa0XswRI7GPDkqRdzkZ6BKxKHhlL2FTIsWH7M+RuOA6qqhBdNZorWqduhajW7Sd0
2/ZGfKajtQyDDeY8Zj3rWoEKb8gcAvAG6ZbnRgsjgeZYMVDN3FK7SAS2g2Glz/DP
tL4l4I+Mmo8Mne9iH7shocYIUh2bhEKW6mfCekwOYh8gV1giGhbNa6IKvuDLZXu+
leWncCRgvXs9iXLN7POFb0mxVKz3P5H5L5JQkOR0qsPGIMUc9r4WiZRZzrXmn0tQ
YLfodbBWjG1BE4+kVIgi6GonVvpSehrhfiNSKWwL0uXj1a7yyICEurxhRHoXIzu2
9y2AEDc+DzPOO/HpBN2HinA0bhXBX2txJq52W5noxMFMtMgonQcAsdu/TIfbP9LT
nTLIGb5J5LiSV9fNFCFi9vPFKcPSd73rrFB5Sr784mqn7of5sZGRjqi2eiyvZ70X
zOiriHIWvJFlDF3hblQIawYOnCi8JWmuCb6Gl9AVrxWBw0iaUFu2IVuXu4Gu4M5v
JX4zMiqGT0inuPmlaufcGfESMVJledOdmyt0N+i2cGfNO+/aPhqw4hnPuqP7mpAe
7FHE6bEVPcochMRTbSvbX12j9UrEdtEH74Ztr+Gm563q1FJad4qjxzOcJUT/+kO1
X5cgLUpIutKeatDAZB1A+cmI3StcQZvV9iCc1sjaEuV1tZOXkUUYA0LGTvAiAbzX
dksZ6GfqyuBtpfLIwR1RNh1Z85MqkgPkT+OZw3u+MhyXd8T4vMmbdWaHraotGo5s
bZlqnW3Mv0QH1/bpTdthpzFtlW4LY0OxO0bubWxSEtTy4nqJ9ZxhLW718EzzBq4X
GNareY3nLjEiE+naEUaFB1OsPT2ES5J1Mg9aLU+Zuyfxs4gGpQsQdATj9umq6EbI
ZeD8o9s1LgPIVkwlmZWB9N0kYILTBpQBceR+/LN38YButwHWL6XryB025ssGz7wq
2v/Ewm0mgIDF8KjcCAijwopjKxqG4makqAAb361O6694YToCNWbno4o5XlaEUttt
j7sLcYdZ0B2oq47jUpIcp19hlfApGPcqpTo/RFoKaVsTGm+ea22MvljCxZECe1B2
YaPiw4w/scpwuOgt43AfgDLnYIyWH5iThOjf6ds1DzWwG3Qhf+KdtUTgdOk3G276
vvHkjkBSONWIuGtlLh8vQjL2YTBc6BfO7xBhdAxxWCxvuZMxLoUvbUK63koyEzCe
9lnxCyBQQS9UAujqdQJ8L/TM5KV+TmIu7zMpieE6U+agCAHHtE4c5F/LsjnruUeV
P1I0VHBfYtqBGlcWD+8yckK362sf4y13jGW8ebP578HfMl4gZFEPGZRlnCicir7n
teq7Y/wx3MFbPXSfinwP0sb0Y6JJPFU5O5UqCyH24HmM3p9pNyiiL/EfFhJ0fvnO
BoycvRQNAyDBBJohCkDS+MDQd5b7FS8sHMvldAxLFyCv6MNt8FZDqGbmNRLQeNzt
gPMetPntraTN9ZaXMFZCTcHNL4GgJNY/5k9r1wsbAYqdY3LbgT5orW3hMiFli8xo
yeAfZeT0K1oFQw7AukPloCkXYjVGjFx5UmQ7ad8bjDl7uj9hOofYpQiCL3RGeTTa
vbqQp4Wbm3/1CHKqyz3ki+HSXCTUvguR/dhIHTZvgWEKXDRnoZpvBS9vyzeGfPQf
D70TWoqJhHvMed05cRX1wA0aE2RlXGWvlYIJbsVEJRR3qQ9GP+PXBbWmC+ugtrFp
/vAPJDv7ZmScPNUdnD1LCWn5eBlsIEsqwuyR2lBQseHzUOCrtz5pt9r3gnQJ6egJ
5RybWL1wiU5W26Beoqzam6q0J/DBQkrlvYOx0kW087THCYXBBvle0U3KYkRGMl/x
16icHLBpnXT5LuczreW3/uWGxZirv9NXqyRFOEZ9uK3uQmNTLnoAVOVqKzQT2koX
Tvd+Cd/GhPvCV4u+5mNE4fwMk+0tXg6o6v1gUI+GDWu74pJ1mwlCDRMeDEF9bgXy
ND8crYn0cUFt81nVK8RROT1UH/AEzX9t77ZlKPKmUYXAgRU9CAI+SJOXRxuYA28O
4gSYj6KiSZS1d8d/IE8geuUpnbJYTzLtdbt4r09o7EIE9ssHF/bYNxRhJof1MoyZ
2sgXiwqZ4erDIMaIVvPnluQeeCwPMvYn4AIVRMaH1UsOwPQ4lzfdBwg5ddbV0Vwe
cPqywWO/oKPFP2pAul2dd8hQ/S/NCpwMLUgRw8TI3SaxOpLZJTKitsT4f8pSFW3s
QspPI9P2FA49Kk+2B+zOiX8vQEh8QciDp9AxyQ084PYd1QyYfcO/9fikGgYrDEh2
NOgHk4EWRphU7EzXvN8PbCaNUnpsnFTxiq3pJ417dhfx02jBbmS95gp56jtzjQSK
tWhREqua+z74qmxYIoGb54IlVn1JgsogVlvcWP4jlCbg1LGm9x/+Rgvjj4Vg3JzM
z2FJi5kn+kDe82M7O4TQlXOG0OrXRd88bWeAaW9KntI3lz33WrImke29656uo/9u
fqEr2pHTd7bg7qihfBnT4PwE9K7UdXQfA2LMFIf8M9AMDuEfvINbpWm5hE4wI1E/
Z2IzfzGmKfrHp+sOK0Qk6BwQgks3QRq7QS/bJ3aSOFasEs/nLtav9jZqcuDxYY2N
mXpSNH/tn/vQwEvYFDkASyYN4M5n5qfb4YDotnZYgLXH+8XJOfOQbZcghZrDVCdA
nRLCYiJLdv9G94SQtfCLLlzZgQ4YLHWLIxMeBvi/pZ3o9sPN4d/R9TcJvXXRj2NG
RzQ5kMxdB8V4Px/aKoyZ7VISOfZNfxWw0B5fAWXBnLkZ79VToACm2heHA2cU/0SF
inrvSmIUaZtRX/pQjRHMM2mzuzN4mDQGn9p/JrZRoN1dpmXIsot+KqGlgrR1loh3
6ujF0DupjRKnX0aw8GgF/E3bfxJlkHUjZD8EJrxAy5qsigAvFFCEgou5wsmOiOsB
ic1C4flLrrknLVqH3d8hnn7OYTHEFJzV9l1io8P1jxa4SWU/EoG71Vea6xEAxm55
FCLcZkqB0Ycp8FRGFzZrePr1P2U3rwRgaZvC6byzXmO9IXDVtPzrAHwpomy2plFd
mIaGLHN7Sj0DTBOKPPy+7X3a41L5MPVZeI83odGAhMCu60FgR6ICQn37RWOfMePI
YsL4Tcw42pY//yDrzXZT9kUIAJwSftrjoPYCsk3IGn9jYhZcU4E8kCNDHDtBOz74
ImZ8fmxIr/tGUpY1GZKZEjlZUPKfJrfVLptt1Fon6333kHK0hvG+6JIhEye0zsPJ
5V7d29+W/rtpXVXf7U6eG0uAbpazlg++jKHCPihf9sl6E0u9To7cBPmve9l8UaKa
MYRoR7BE+UESgwz10xaQ0Cgi/7IVBnDGy43y8d9HJJen/W4aGs6VjFF7fMLlwYM1
EceaNUazsmCuZpPCkfdGVHuoY5rqbOV+EPhir63IrD4pEXgqpLjhVe6O5A8jxnhE
0XyYk6FHo9Lc7Z7sESBh5Na2HwhGs5Q3oclIqKISK3RW9MybEIOgLeXB298dEyET
vqhEFufJYlLxbFagPo+tM6sL6CYm8FOBLha6pKQE72xH/CFqQ8ZZxBLzFxOEtuEs
BNsHOcv9HP1jDP+6QExS/k7Qu4bcZXusn0j9UkS5pl2KIpMfWc/F/R/XYq6vbmtb
5N1Ellqb4Ft7rIhJFDDKcZ4DMYJ7R6+ckq760r7chgxYEEo6InGdV1WZ55QcuKeQ
wQT2TIY61fhq898YAnatLMlErXDwpcfU1J7DxfPbf8M+DZK5rmp1Q2XeaS5eH7Jx
YbuKZaKn7JQ6xbgih+fy4SBDqC3seA4rVw8J+/5H63iymIlY01CrQENkJlWJari3
EEcNTvUTNXSh9ZL4BmPWwtK7WcRiH+JKR5TgDhFfQYIJguQI1yOgEcf5XfaljIuy
5opMBxelA6vx8Q6ouxRYS8kIAPCe5uwiQxfiYIdcM7sfMPcXokrhEg2S9aZblEur
OkCWzn/YEP7eQRq0ibFxTwJN0EUXYLft/iGz+jv/10zIOUMWNf0rZDskDtZFb69s
4gTI7Gmap79598l+YshcPrdVQ8AZLEqlc06xHlDXal72CHZXef9qXAlQ8S6qbZOD
XU2t/1YXRAU9uhqZjKEYj7Y7ihUxWOVthaEOb36ELcsYY8dZdXhgcwJXwpERrH4h
e7HRWn8SZzZEMYUxXLtz1zLGjEnvLHUb/fCDCOpiZrzaa0I0RWV5qTDTI5joCtIU
5pqiEG5318Q7Q0ETOGuX6QtPEcGKkltKir4J5hx+BIPdWlCfFNI7c0B638Jdo9bW
CXu3GGQAETA8oUcvnTYYbw1MFgmv+to4Sd5392fO1xseTuVHybFPCes+9GfZ1Ev+
E9Q36WggWMOUuiDmcoSKiWz+vTwg5J3M7Z0QOvNmCiNfomdcjVPfjqZFQSntZxyX
T/WVnLevPKkuuqk3m3aQebxs2dPszVTk4HxlG/OJzVTTuaS1RJTnfftHeU39cU3b
tdcwvTUCI5mIqgmnWMrfivWtopAbmEZ77KoSFJ2v7Jn75Twp2Y07+m6ez0erYPjs
ai1WoXIpoX8vGrpKNvGXaTxz9rQ3ahWHzjlG9PxpCagkPh6q3fmFFraBcfq+ucEs
NbboTOvrEJ9oNdprNW/ZN3Z19ai5aTViFWIa0murIXukII/Ye9MR44wMgH9NVL0l
59ez5HBquDkHqnCT7HlowU5+g0CBvFeo/rkkrm4Iol2poMMPntJ5evIcnWAhUU6Q
hiiTNNUDXofxc0pPCllC/X7ohUpG4GewBQ/u4w/rZpKO/QvVc6vDyhmUbuqppAxC
Lx5LUFWXEsvnZEsFUHXukofJSftuuOsnOiXUMvSSfmk8XBBYGL9A+y+XdEa1Him/
narJ6gHsfKOElEmnGExeFUeiptRwCoPao3YM8eyetJGyM4WZ1tEwsOw2gW/uUnGd
`protect END_PROTECTED
