`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42Bg+PTB2MByQJZFSmE6UA+E2EYSz6gMjyj73VTL6WNa
7vzskXjcmE68ooqK5hDaaoiw6GLs/WYUxQzFcC8ZZ5p2jekVB/ECk/bG612TFIPF
6AGF/GNxgxepLmZ/hulaSOXyvspRT0f05je2LnEQxIq/nCSFaycNXKzhhRSAlV+b
9t10xW7SXSCR89590sTXTWiZBUS6AEDFo8C02XhR9wr1jPrZqAfS5j/lOM2WxfVT
EFVz25BL54tbAefUhnPu6KbQim5eZpXQ2HyPSfNCOStsepJfLGhhBYGnjRfPQjFt
w6iCRkBSHGKCnC93Hzq9BralBEYmDR4lxECQCvjxCQy0U5lnKMjji5p5l8RYFrnT
h40RMTOu1nN/xs6H9X7kKCohey3tJbMUbx9UeACvQEFz/oawXVwrwgQfD0Ahpy5W
aftXc7AUDk3U2vudWECvBYzEjzCMGnCEl2DCVhx3qZal+mCMLI0ekOvHojDVAf50
f61uyF+wl3J53FC2gTie5qoeVG1Phm+P4U6KPZOjp9FuvOvckctZ4E2BdsAIfDQN
ZZR5mOH3donYFfxQ9K/X3GQL7qC0wHgxdLZmCl/GG1h2D3ypoFIyA8ezQUnkIBjc
`protect END_PROTECTED
