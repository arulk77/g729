`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCJa1XhZh4VEfBNfNKB55ylZsdvd+8w8Zh+PKoNhc0Wu
+0XtrG+VjnfHbutUD+Rinjz1kvqHqGTk0u9+WIcXaHVqCRov2MeIFm8VXJ1YQsKr
0ld/wo7PtAI7qZjjerOUwHgGAIX/sZw0gf9B+6XVqf62ntglbyZJgwIY/GgYZ6Uf
GNbTsuCt9zq8cp67kB7Sk5GUl/D6+8jeqr6xU5loDgvp8+yfy5JPImz+eLVQOK6r
q/xDsWusHawiUYoT0fGvGcsF13Yd0t3AsCQOQkhNF5mThsJEyKSqCRNrfXbv8V4k
eLhatfVg8wYHVFRWfvoMYezE6bl1fkZhBzVa6EmE4ubSyt6pns0kZLYyILvxtbqT
xWeiBY/BOw04UnP5uTMil+LtTrSEgL03s8Eg2nuj9GdkIaEoNNbyVhtc9tzSgmlb
J4/RtK5uYTQBj1Ea6MNXOxqcpOMp6Rth5QNKNoOyKHngVCim3vwnKTzLSP0XoqFe
xrvUSFu3SRFb9fRoQ48oN6oymRymf/KHqofBkN2vVaepqxdMhsg3DhJsj5tRS2YW
ySO/1YYKPfyp/VoHkSlvjFvuMGgXR1lStBrrkp5srWdVnkBZ9S+jfUZvwDgK1He4
`protect END_PROTECTED
