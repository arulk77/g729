`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C8LuT2edql5ko9gbYDzBO07galYUlHpQZQfi9i3RxeGT
PTnqBBDzY0gpr36MR9G+rEIR+KJxQWwvImraWE+JIqRnSpiJGkgTrL/wNXwpy9z9
nBZpZ5NN4T/grHfa/Guwc9g6oGhAguRVISqhx4LHZcRANbMfZv8jRxuq5IDEQgcD
DIQ0LPlWNfJqEXFSeYYMKCS06P9uzq0s9FAyuhEnP9TZoNRs/HKbU9isb78h6Jzk
MuTNweaHLkyY8oBaB894477eTiYkmkPrElnbIwkogYMullmu+2HZTVw4Kfj9bLmf
787NdUlSho69Gsp8zXqMZuXa3hTnZj0OwLT4RYAoDV5Yqt07FSE9ARklG11DMFpl
OZWgla9zWKPc22IssCpgdRtP6yw5LKkac2xw+sh12JLk143SYOhzv5s8UnPFG4xq
k61Y75BMyTZhlx8iUIVcruYzJ591UnPt6qUWgudHIfkOs/FhUm49Gj04uASAfueq
RGM2XTymX9wApaLILyWZn7RZblEA5t7kupDol30d9AA8TOPljcZXPVZXSQYSbcuL
/qVL5P6y8Hi9dzSEHQuoPrTwOkY/U48YYSsB2O6ygC4J6Kvd3gWN5MAeW7Jl0Mgj
t3q/8YtepozJFqddwCzHuS7zjMQ60xXxJ9yGsDFIJjLSPtSPnc6CUi8phvHrGVXg
d78n0xW5VP00YhR3YKup9oKW7PThHk3nkNOoZl/LiCVKtlBwmp7ZPfeSvubmc26X
ua31iloo8XVixDJyd+aJWSxHM9eFG3VWl0o3/hEQ3fjvKiBcgknP0VN64uXKa9wZ
R1V+L4B9LH6d0gQS2wqNQpJF+Fyg/4L9npQTxjyaCWBR/PI7fCKVTXYetbIwH8Hh
oaYvFj1CfaY0VlyucJwlBRJkDXqzKJ8QiE+fKTCGAHGFv5TqK4nrKqy1T6gSXjhW
DqeGmVNiCEiQE5G91Fl69Nbpn/ruKDk7aOzHXB+dZkd6ojPH8JPitDW6VXN6skAM
imCbmJohbZ0G7h6sOMm8G8sNZsgPIrTfNIB3CQmtoaKn4VDr+fmdg/RfL2N2pW42
XLf2ypDgKrMcn8sR74MnPzVSGsHnRdnz2SlhRV3J63lVSPeVgHcbwymATUWXLZIb
kXUDOkKHUKK1sWLrFhnWIk3ICOPs6a8XCggvW6mEFhei00c/lfJb8o5MvCZp6FVH
DwP/lFUB39jbA26h7UbqjjJFcKRPeE1tEdsn+fSGdkfjIVDxBchjdOGm1Vp47FhB
t78yvz/ocL6RflMe3eyrLxxuLyCfbaPA7WW2OiIK0elfy4tBC9Vx3S80r0ggLd3r
7PmG1J7KghOivrxVKLZ6Ays6MaZfk2Qj/Obn4rpJipJPsdQxg28Khwyd7r0WvOwR
Y6cDzmyFsbOQI18PL9B864J2PsoKAErCvNhLe6VxbA17Wopq8859lIeyLx89mEIV
9+Xuiu/aNahaxnqfp0d++3XkGq6vpfVKVN95DokTS3axoG0dOVt8MmtWv9Lhle9n
xRhNCB9sJ3d7hK0XlD9EjevxblqHqUvJuGL52YUfKzpW3ffTSMjgyhDyW0qNl380
Ad3WKi2EzsXnULVo4bBuOehSHBOQoxWafLlsheSuL4X/svYTnZ+6pFzmsRC3cQqc
bsxKERgF5Jb9ck2+Vipa3ZWTOmstfKPFzTRiyyOhHmeuYvE9VQ3+L6VK6QfVXtCN
Pb7eTi4kh8VS0V/CCqabrrTS7tQiC9ebl4IUl//uuDEfMWlZM/VQ1t3UCZzPH7MZ
oMaIvlonhyL1bAFdM4AAi1aSfb5wOIZFVBlcQwPQ4dmHeZ8SV//0Xmn9NF1Fv2je
5qwfPvyAvYLEax6lFYFKgqAbff2uLKG+lt4OuqtoW8BHy1cyydDVA+eG08unoAwE
kxX0AaHHEearQYUD31NgJ0KZkjf5IvUcptrGZAENlgXMnkPnTosFvnjTnYC9drKH
X6zZvi7k2k7nklX1nk5Azy++ZVNV354wN6MiDpApxNwbGiwog1jI3UK0vV/EbT76
NlMNcd6O2vyRqICPnLFqGoEcH4fUbAPF2mrn4gBOzjD+DyPOIZxZIonAzgn5BWAt
lAAX0Ze8o5lX5MechIbktFX15PUXruNu18qrH1tRFJ2YVmJcNYLJ5w5pXg0dB3Cw
guIODxPVJQzhBwPg9fP+6OZuL0adhYlfYak69JEfs0qmFu/dZLx2D/EGnvrXNeir
GJPNS0KLlAh46CocXeCfP1y7lywYybAm+CeSWIwC8oRiPCLqdD/8eTozwgUfavet
+HUKn2pJa7SdEnegyHgB+PAYsa3ZmSw2NpmxCYDwsRls5FH4B0WCpPqOZ+nLq01Y
VpdonH1PA/3av7g/omXugwJTfDyfGWR6qRf1v5eN8HIs+svMULxpnFSamH5xErqH
XSe2JK71e/lJdj/MQSiJ1xB+XYhqlZRCfRRh4vSEIRSVMHCUduqO1IzScxBoVSBC
6at6cOLmp1oo+y4xQJIY8/kNjzoHqeDMP+dMDRg4o7vHYP6Vigk32/9Fl52YxwGh
GHPSm2SZHMAUSewBANM5Pbgil9q6R5NqvS9ys9FoWqt7Nh+dtGsASiTkq9fFP/zg
lqqtwyEz0oFfZR7WiNrQprirLv9URLC8wX0AxmDmpc2aadBvU5PMc3a21u9+Rn8S
iQWBtCOPCmAcZ9gldwrTVM2GLzPlnOIlxePncQqVgLwo9RzOjA5koYkDkAy046Bq
G6rcU8NfhCcQnVSDBRvbx+sXAlvqbpKP6IlQmdIN0GPhjaOfC0s2WvIAGvSql/Gu
6N/cKQcatXJWfUizsINAe5N7pKhE4qJIm6shsbTpZLVs/X0DW2m0SGpR9FpehNDU
lvry3SptoPRWKGxmnSiooxstw6aucX3veCA7sCiaEXQAETxGs7CKGOOdK2NcmDGM
h6kN1cpOuczr349B7m1xSlguaUCpozcfRyxP9BhNaCFpoMDKxZlTJV43z6diY5h/
LP+EhDyrhUeGlhksBqWFLLpRyjw6e5uxuFiNdHimbpv/WLsRvsTSoo33hcHuBzd8
Ozd0mCFP+CdkvwO4PSD9vwVsQPJrjcwyzY5FWks58Zp1Z9TA0Z73D/uwI5KYp8RR
aPvk0fL1nHPaZ6AI/ShujA==
`protect END_PROTECTED
