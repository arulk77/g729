`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
PQcLXZSRMBYbNX0SFFixwf7v+IoHjwGbvzbdkgMBxyzWduPE7REzZ3DevcqjMEt2
z6k3YYck9kePsD+7KDOWE2qmkj7560c80dqWbMxda3F4TkaQbmU4BEbZyRd/gash
I/dzi9XL/8jA+9XIEPQI362fRwaoVFmYXCyftlzFsO5VdmHHZ/ePx0qzzJHnBYd2
ni6NA++b9luTFzqM7P9PSxqhRN0GsYvAdlckySyzRaNdBiuV5wXEDz/+l0CvFOUa
a4FyuNzUQpe4qRZ4teZc+g+Ne54vZF7GgATBUrI4WCiUxIGkog47/D2kHbNaPcpg
Dz0RjeY2jViKf0gtUzWkyxFmjTj25RumQ72v2sNbHblF+V8zdYbYdAJB9HcRxskO
FzwONk6MOTeZ711UHfUtp1wYM3p48pfaocLJqwr6/QKVxRq68BsYKu44b7D1imk3
lARbgmPXn4jWkdx/MmA90VEW9KdTOkHNAI/3fusBHthuydEPzWW9kzTsVH/T/pqV
0+xzT3OfiXsbcd+3uZ6bpCwFWpGXV0CraWsyvlOwS6I4Eo3sa3KYuGpHhgrr0pka
6RJqjYXvc61V9mDpOGpRTS+g3bqgl5MmomSwJPd/+S3DQFi+G3WWxjTC326I+Qk2
g1dYtBmpeDQg9OJF0/2bqRn4YRom9AvNjgq93OPgWRxfc0HZUb7YBCONk4ENr1lE
BD/adrZzdtJZkOhsJhjLUr4qIBK6Fk05YlGVNgU1BJl70jUBLumL2PSXvDxwyxZo
PSl23WycYADAQFMCF4bgEm1KlfSG1TR4cWDW33nDAFQRW9YfoZasVasdKRqXPDA5
eEnrEt+pocu4uAs5XRnOWGaXRxbqU75i4QWUw9IQPT3BqCITtVrEYGj0C5aItTFn
Aa1DxoUicUmwIoj9PNHj3PhBVHMqLZ0cdDzQEgkGMCvcSfSNEBen1K8P+4rVf1Sr
Wf8rgN5sBC/frk/8oXuSvP7wzCDQVzCn+corsEIXiXHm9UR184jVpqYQs+CJY8Ss
FUUhhsnYQ7AZAAik+ae4VpfCu2U1oPb6k6q4g039N8E5i7Bj2Y6nu9c2rCp4QTuV
kjvPyVrBWJ9D6prhR3O2nHytMP4N36OUMzjfSph1/PZqrw3U9rJiFix70aqC6QCj
vuGWXOTAc8gOQ8epSaZbiU+123cSmPmG4/vjWe3x//7TOPRXkMs5GIBOCuDFlgFx
v6G8sfyjMTSirZUgFHP7aFM4mrl4wOKvbM1q1rmPYnz8LfjwdasEpf8/boSzsBod
7LFXJbQsl1bAbZtCLpi0zK8RLOCiBQlazZxqgg+CFdzWmHgiQ36kceDKI6dCcIoc
wmiLXv1ht0mV537xc96hJmLWL0BD8z7LSM4078h2nwfcRYlUb0j4ZH3YHgbkOBb1
WLIHhXb/Obe2EKW9FyToVHpMjIcG+CK9dGnmQbQC/T7Vfd6weIb3phtLw+Z6IuYc
bqecmtB28QBTXDOOR+EjAypdT61eDslGFsoWSMfHrnEV+EhxdJ+qZGw4UiryBnNw
HQhmOLxiBz38SY4ZKbY8fh39bYaUISArihGcRFiGaq9wV7Z7fwYLnR7niIGIElKI
1H+4v3ol4KUaH9hKQkQrdzVZjZTXwC3NCX5vli31W8kGqaY138RPQ20+Ssr/H+RP
`protect END_PROTECTED
