`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
FRAOjB+iLqIUa7UpkgWw00oXCj9/+/YRlMpRWydkCMApsT4RALFbvBUqcccSBSVd
Rc7g+rpkni2AVKffPgQCKrCk3nkd8pcbFSq+T0b9Ca2D4MrYGvHFFaqblQ5lPO3h
qhomgR3oEX44Bgc4FSBoMPBMTlpK2RelU16gG/OxC/bFV3eeEDjaP4zFQabQ29bM
GVFV0AKUtjc+WLHhuqiEI1xgERytD7FsEraV9myloUI7/mSDVCIKBoEj6TsJQcvk
OOoo6iITg9N4yzG3U0FXLvzvnlse4tWi0NUlREIs+LhgURE8/bFYu0Jr6ynVrQze
sa+QEO+9jh4LKxv4a0BHsvtQhYfbjn2StePtgZJJJFw3E7Qh7TQ9osoiUrlYy77o
+p139ivtn4mb7rVp04QKEZDNB9FUprnMhLQMujaFvFuuhTWsvVlxyyGdqxvI9gtL
WScTZWKnchtY3kekd8YcK4yzgy/xDobn3JVVX5siSOXJIub5rCEW2jszCv6z6iDk
mMGMbcCCG1ToKz6FyUdgJApEM7M3uFj4u6XZTEd6Ue7heucc5lNt5e/Rv4W/SvKa
GvN3Vw2RJoy7Qo2GTenb/zp8B9mvKZCV7pKNaB2BzQmYO4P0p8QRJjFEMWZV+XaY
NGbIDoT3P6jhSeF15vILTVLJTNiJe4GoQTJvfOenp6SQKd7WOagGXTdEFCXi50Z4
4pYBGcV6mRX/nZA8YUwG363++ww0+aDpq4cdEb1x+hO7skbgRpNpEWCrzqRQ33Hz
PPijJQ0QCEJWcg516vNA6c+xupnyybRvGpwwNyLCXHzYJ+a91Ke/avOwRIgita86
KuwFio+YpASfXfq/dQb8AXEEMIkViV907PJilDOLB3XqwSr7a9soD+wU/QQgTMMq
R6jN/SxcUU6pnzexR0pC+N8pdckUYr5mNzYHQcr71lZi/DCESFb7XGtxZPbF7SfF
9sBZ1cWmRhEZi+GLPZJgnJV0Nq3UG+Ck3/B6Lu87F6D1kmDyXbJ1BSEPtFcLfeBT
LVcObvUUkAl44R+0HJBGx62vZDJdsbMXGMWkdV1GKy42WZgAez/MgYx/9GuGIWr0
jRXyw0EjCb57v7Gf22thWo6Atp3tQ+zrTdVmnF/r6UQcY2pHGUM0JFQCCARc93e6
oJhLjiLYhtzH4vEa26pmSsN40Nh6sAG4Tuxsr0xO25Ik9FuOK7SDt76S8cDwFPEX
fE436du1kk4GbgUs2cFD3w==
`protect END_PROTECTED
