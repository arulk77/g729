`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mdujDsR/KvUeaBTnlJy5NoFENFYuCpfS+H7gG3ZcGLnh669mxsnkhqRKjdw+0KMD
4ZONz1Y/ryqzzFPV6lbgzF+JBu06pqEIQdLO/ftx6cl6h4OGjP+Qz0KFhQn8vRRh
xHwW9ivyPcLwE5sn0rIUyNdbul20Roi/iFscduF/Jys48dCB1l1m4jAVMH4jCbX7
UEF1pf9mazo3Kb+9Jk5Z7xwMYGSQPYXESmd42uJzpqEYQe2YyiTtnfeh9x1y8PyG
ffXnpurqSL8vUK94H2LoZ2C5FP4eFTb2E0PpI9id7C0Fqplvw+h7F3fkfdVpvPP1
u6HGxmRr3h2Z+yaEX9N5OGyLBUBjmuOuQjF4BC+pU8TN0uPEexgPR0GthE3wpusy
SHLg4Nu1l2d4s8UoONprz/iwv8mUUiLZ7aNmBjoYCIeF587EnfKCPqPRPl7vXdgi
4R6ARtmUoyq24HR2N9gljReY2MrdzsJHJ81JQdOWjKEw9STDGQYCdttj7dFXkPar
vYI5GQMfxsGhWu5r1Co6eg==
`protect END_PROTECTED
