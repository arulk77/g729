`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveO1Gb5uA22Nd+dBSlGZHLd4DjvC5GXU4v8bzvXoZm4cL
5Mrw/9Y7EhHw3ldUgMMFQhv3x0TrZG7Tu27ZcpPgdW6n9Eqoto/8Vtozj69hhOp6
lbYwO7d9bW2sdXL5++tjh/PtUS5XNR2Yucno53Ng5fKt2MTuHghtbd5cjzPpv34S
VtEpljg+iuap10u0AXwfPw==
`protect END_PROTECTED
