`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNdN5XNx+s1/fzO7LlTMo9kLrxiRHF/Fwnlbn0v6lSNT
TVMPC2mA0YCX19bKy22yKmELelD6xWR9Tual8wAEdCzI7dYlQGhchtLe4x+GNMX9
ekmQuIMj7oHBMxlF6ASH9E8MOrIEA0Tj5TU6vBH0Z4DXUyn5ndjigYaf4FKUM0KI
8AFx43hgZzGfaFhUXy+ea9nSG5NHNLvOn1tsCNohQzLMsD/HsdFNSpnFitAwaLvG
edq6GKxOgbpUUJU1zyVha8Y/HGbO4bDxLqyqsnXQrHUvbVC730S6BGfthsX9fQt6
vgmq+Ibsa/LyQXqPBEm8WFLUxK2yq/ueDhwq1evxw2CEjPkyb4LhXP4sCBF7e7D3
sFeMJddW5QSqo6XcCTthbA==
`protect END_PROTECTED
