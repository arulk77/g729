`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGZzkoUDCEQwBJc8mfwi9rfzgDp+keFAkrNxgXr9veFj
jFyZ4NnQc0PpPgh6qZACWzZD/EvxGXKo5Vd6c6SMGI8r4LQYtToDLJvT/H1ZrAFH
S8FNNJ4L+vjeZL9LVyN7AEj+89XhTdc4HYvq1zCnaOEnSgjHfZRWdZDGiZhv3yon
gtfW9gPQK+FoV/bzAMG1cijBG+vBUWFoMbv9r9ZqdCg902Er71ajbUe1ZIrh5ljX
eYBztsGeC7txOiNcGf+I4pIDJJEe/seExZEilaM3e1jrPw/kJSe10X2p55CKjP1A
m+H6HWXJFZuGzh/EnYZBvcb0j/GTy45Vk2el3YAu91HDMuSrJns0F0RhZyWiGmYw
PhPWo66YrixKLVpMWUk4rsllfp6xLu66lmYH/tmtfRKao8IJ3eDsGZHCCTtx5La2
td2IB8zVyLb6D/3wabbiY+ZbZ1pizddMvsLhofgzvG+dphBIGHohN6gsiyWtOHpH
vyXpp/pYJK2W/rAm3eJd0sxR/TPq8gNvH1UR8j474TSEIA8JOOeMgcfYYEEoeLSb
mAqi5KWZj4OpRGkn2acB+8e8SMMxbwsbyuefrP3huq6LMYgrEseKWkBkFAUdP5LU
5R/za73FiW2nO6LZqhJ+mqWa6KmVqNM7zCoGhwcs5MpveGHTpIPJw6dS99GDh5Zs
`protect END_PROTECTED
