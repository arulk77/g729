`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN7i32WVhyDgsl/bGo8TzymC6h2mGdMEFTTIqpZ7y4bFg
q+GWh0iDGypmLJW3BBIf+1wQ773HyTg6MPO71mU0SIC/tvH3KMlrT4oCPU+rT2TU
/eCj/wUGgjSzDDAH2dFYYKjbUXwOxMsFhdxipyum4PKsQfcCag8vj9MXTkEgoiJW
Nr6GrFSHvJ8/uN2L2Mz6Czm6qWGtTPwHLlFqOB6s92r/PVzbXPW8B0eMeLywgqbw
YGuRsM8RNSfdNB68ck8vgtWHwkY9pCzcJAYYlP1EcGuVuR2iQds5jSVTaXnCWUS4
9bMFh01fNKwAqFZFSILB/3nB1nQuxwBAVvBdKR+Pk0g1RejTKZskcN7+T4JEacs/
geXTOSpgpv9VYZAhKQGHkB3rblxsD/1XkmQF+vIrrLfkrsK/gQsNxHYyMKxTSSuM
du9IIsVK+8Ejc/zSto0/+uymiHO4rKX/5VJfmyWUjb/KgzA3027XedpyxTRi7qw0
2DewIsWfcy02keTP++8dNzZ1EGYn3t0z2BJsW6DhyyNhfs/zGJbqa6dITz529hwR
aS1mZHuuRGyBtNHnGfSzd17W3SdrSXG2lAhLLph9npM0O5UuJ6NFpONC/5SLOZVH
uPCBb8b9NYfRRi9T34C5DwY7BEDRJWO4Q98WWdfDnNJUNjZR8fEUme91A4r1VaUC
go5UZhxy8Q2Hze1MLVtmy3msFGNPr8BgQRQNiL2gKlFsVGx/GdGddnM2gIIaOHgE
I38Jr1XL0jBbOSNq8EhVoD9VwcX0GKVSvndvDw9V/6lK2MWTdVvHCdR7erigE05N
w9gnTCF6XQ8Nk1tmb68SWXDusHhQKkNNlmgffRjmtMSq/mgSViyqqsaWzDydJi3l
domCaHRW/W8u+yNq9TMedpXAnKCMbzZDaPhcXf3eF0cEDXQ7iwVAEANOiBqBDOU+
OKPUWwwYbPX3Gxx0koVtpVlxuKDbBi2/AFqim1xCUBibCDmncJxCEYDtSnFMhN+0
qrrfLg08WON64W441Ai4wWSpQMJ6SrITfCDaX71/FeAXY0m0CNofMf/UMlzZiteS
v5OJZmS9eRYc56ZQ9uVvfe9sfJYivdo6hEj4mALraO4ibwIHNnfXOwvT++HwSSIc
QjoSiZyx6Ipvy5e6AnHZjFPNtOaMxOnZeWGy7DujMkUFCDmSF7z1MK9bHC2wrEuB
NFTFbuHzg98A+kHWvylWRAgS4rwtYktFkkWcuJ1JX3cjzPfvm4ZZ8u/isUJ1kXwW
mj98u1gFfOqs4ExHwlIlQ251Kip7+0I2pFqlMYK6UlZgnQODHBzYcXzrYT8+UpLY
2F2m4pCnLVQZZGLSJ7zGYwEmKPny1sWqvzUZtYj/qsTDjaMy17W/QdO80hhtjhkz
mqk4v9bdzTmokiPcgchwJEqMa1E/sjU6Ns3Qd2Unia0YB9cOJh/qB7n3jm598xoP
h2CUIbqyTJseGhNsoH5fn6QZmtjLgcT20F0+VonTZVrHQHI0yBY72qijShLGjP5R
lZjxTZy7NXplmD7F8ZbKah+K1T8e2mgnYkDrO52W0SoNuHDj1KkB393IrdjDpaQ6
2yI3f6GQ5MvaMV7ufwTHs19c0M3stkVqHpRcqZOlOB8Xq4Mq2Hw9uHygt0B9SX1+
1c+WRtVCB9YNcPFDAfLRCvciARvcd3nAn9WbBhlczrghTurWrCXqUv4h3zDV3LWQ
uwgLKhQ2HnrS9l03abBw4YzlK3f0XoRzOahd+SkWEkzQC9+ngVzqNkpOshTu418G
b+FBOQ/imJ5PqFZPmSrai/7OoSLmMDJ945IXy+PMW/K+QVPLKAUlY4TcfuJY7SJq
0UcAkts86jeXL/iU1d+mCHHlUVLzUQUow3J3Quf6F5KjDH66WkCnAEEtEqrHaOYf
/YoeC7/hliQsDNA3msZhG0w5D8KiIQt6Nxp0/IwDiZBk24YHA41X3Bjql8/cmHyx
TwDVIratS5GXTDEGhVgT53trVP4U13dzD97cXoVJk2rk4S6tPpqn912eAkxrTF4G
kVg/P3VmWbNEolKzNNTLP8lJl4kWmL0xPRRZxcYGLgaHNW54NE6lxGNUmDmBzfg+
vyhAbOMI8Dn2NSokGH/uZnk/auurzEmWOdAAiCPaKycfqY2TY+OMCxfvZiXXNF3r
tfTwVcS6QDxR7cCEIvJN/ZaVWuY5WdXNJKwCi/Be6AlfNZvUfYjotM/61nYtQwwU
7c9TCTZ8TmzVa7x5YTf6LE1yGUhhc279wHWsXw2POkN8j/cd0oBw+pbGiQ2H/vj5
hBQR0xa9sVlmN89eEpngEsALCKyF2ezGvJEIYRqFyMlYgj6deawrjx7LwE4VcF6y
b5Ik+lXEt8HUov2w2q9WrQkxa3lHponxx+HWSq4TYHO/KeP2IJLb9VJ2j3SONehw
yIiurEAPoCH+ZK9XlsnicBqgvrc1eRLRXYir2JfdjIUSAnCei5vFTvOSEvISkGDa
jwznCSgRP0ZBXtZCVCLu0BmUJRcVUnPYoJJ7V2tb73SnfyEDi5DNLB0HXutTAM0s
rtFNR6qafLktADdJNM/vbuicj+S+hT3cePRxH2iJ/yXUCXsecN6EZ0FzK1X2Guwb
wMhJhQ4P7nHn02qqF8G2/XWD6s/q1r1SPwR0ewmnmpnmSJa9y6x83MEV2aHAP9Ph
sPQ2HF23UTL7NPOweJrUGUg5/LWaW6+KKswnjGlY6UDayINyAhwq6ZIdMhR8XThv
YMoYG/2b0pZWO59WPkTz9ORbEdvgw07baX4cj3hqGy+yGqu6T5IS9VRnm2yn3O3O
Rh4DuVEYaPzQeJWI68NJMXCxOZYtSW+8fqqc4uYBw8QwBtIUeydqD0OaOqxqfv4s
bUHeyFK8WQPetXH3vxd5XYAhNDBgSCeiPZGsRFHZq+E5U9ALCgw1giATG6kdpvK8
ftgwaUwguEPuY6M7OLqa2BvSnJTp9OwyR/HbWns2/XpM/KxbBSJx87YRtBT2Wmi0
cq3Z+6B3f1DoJA3XmMcnG38ErNMEJdMh6BQejkLzTsas26fc4XoXTmwB2mFXzjHx
fn8dCt6vFaeas5N7SpjLMIfQKFxfEEs/eEZ5rwDkLtoDFAaalTMYAu9tyfNyDSBS
5Wn8Pd8o14F8YonchPXt+vC+MBhraUCtNFJE8uwEhvrnYjOq8JCpeB9qTrPr0LG+
ab7vTkIl9jhickX4IL51UoQGVfOfhpnM2P4pPvoLIsY3aX0pOkZ66Jgb57vQ5LBX
4jcpd+Hbny3TVUY7xcJ+w2bYtTYGjwl4wuEPuhzmyOWfwtauPAJtYJ9nIaIABJd6
KG5UYSJE1N5affrX/JgVP82SRLl4k5kjlun/NalE/nxsjjiwQtVyHZIJMhxXQIn4
8CemQaIOLuRBrrEuI+KledVJ6c7rDe0CGKLLE3Pcopbx6LLdqYTbxslOSmFP6obE
ERzyN5nNyKOtjgQcFESuMdLgvjBOuPU4CKUfeIC5TklgR2gLGDMUnHGsbj4RKDrt
XazXFatZWf87XnIzqWFAKc3sx6aOSMuhaMjWBr0gPPkxLaw9puwi6PUDY5SoDuuT
EczLHhHX6BC6odH9JyELO6RTVq/2u2tsbHYiwr40YX909UsREWylV/zTarqoYmZo
Cst7ePgNyR6B7KqOIiy6m1VRQYiek+WbYc6QfbSu7A/ey0KoK0N+poq+DhZAuDBh
/1JKBjEf7y1V8xhvChdLmzuBADAMZ1i8OHByaRZvPMaKv74+mdUePWlGv0eTRZUc
V0M8p5fUU0KuMOqqL3PGsM8CFUAmUguN2Sl2wI+WZcBYZc/3RWi3mrXlp0PDGOC/
1lQTVWRocnMx37hS+WVUtIqijb1KQo/qY/KfAeFZqUXgoQtJT10vR7XD514xuPOE
AvNpvGm7OiKPJmOmVGHz+JB7/SWDyC5YKULci4w6QMcTweRjUQE4FGmCvCR3dJdm
AEhFICv/iO2wBC9gePf4cr9vDDF7aXPVcEixmkB7xl4XLQoouLGTzYJEU6dZgf2A
mOO1BuPiGFzF+IQ7CZHk4VhB2m1QG1cesjQkc67JmmwzuSkSGwN0XuRwR/8IMg3u
Mv2k0wS4es8btRNUBPBd3pGJ05BGECrGhLWXoiArawDnwCiF3B5Jt30izy5ZC7pn
BVi8Df/UxOKnrEBNjXvlxZBwCYfKFmlrhoflB4o2PgJ0X/8nCHKwbBrkoluGPl4g
qJTTYH+sT8veYPm4x29d8qvOh2Vhu7kCxXtwJJbiB+tyh7E3bbRJvtBEDisoVQOv
uA2ii551o9urzxKL7E0gQWsWsYBVgAK/WdniIrqyy1ajwVuOuORBANKB/79rrMCW
YPoZEqLlP+ZSvtHo4vOugLIczyuXtCFDrHMwS0y66d56lr6D6F4Kb2pI64qmwuk0
XGhe+d0BeyHNmyCpwR61y0do8W342GUwj6NLwg7x187m6Ti5Egi9O080FBez3G2Y
JBN21jKZK19/VlUKFV+b0QWU6v9l+p7AIPrFg9WSn3BScMox5U6qhbZQlNRpTtLZ
sOrefKx62UdhThNvhQZJRb7aFd6qg+fCAjBU/AYkbk8kdqESBo160R/akZPAsaQ3
jEk8KhhlAhu4PqXti4+ueZQ8JsJrNFHZKunmrzGbYZhL1YtwIDjo+BB0HOZnG4+A
3PtOQUzS/JVfXFwBb87qXnkgYqtsqpS8yKS8H/MegEfonbLDHouN5XaT3bI8kwVH
UiM1bK1jYP9o2G43kwjSIBq/eHBt1AY9ihGaIZXMiaqlSZJLHXo7CeUd9llv132Z
TkVC24eqhup8QDoMKxiPhIlSKQH9TM7twDGlPcoO2vLpz1bwN7cdjSBlZS54OySq
ylDG9v81cDLQcRSYpzljKtPsXRTxbdPodt0y1VHgd3vxYM/q67pB57oaqcabqnUX
/oNNFefDsZ6/GJJtF6NwxS/QnqWKBVk3567dvyekHCNN1b7As+V9Zw3MGA3IpMgt
BmoQgl5/c/uSW9v/ao+/HU/Ds1nPoYIhXFKJyCkrfaGT7oMgqE+2+E0/bEFg09Ok
96JpvvHp515fw9SGQCkZ5h3LiTnAaeOvYyT0M7Z/OBOiZvKRpC85tOoB1RdlH9+6
Gq4MB6Xfs+3ueFwlgm6ZYiZTpQ8y6PBeYVivlzrxF7vrtCqXJQnRupZ89l76+3mL
PVFvXqihBFxEln3yuJ+2xlc1clkl5rfr+CpoFCLNSF/HiPK0FsKNV43TpLxLQZTK
blHpeK3pN8d25KY6lSUA4P7zjy9MatvI6nISph+tsE9/F+gFT3vnswd9udWe1YPA
/a0uWmJaqcwNBqOw4SN79n+tDcq/Eal+npHtWH2sNr46am0ro0nDiWKKyMYO0JPU
HOniE9OanJTbKLw/Tg5n9Bq8hXqftJOBlKierVYxLSaOxSLG82UKgqHTOmbdqvAF
FxXnCCwSQttRXMPyRvWclUeWr7LqnootrJ65YxXh/YpXTlyF3XQy2LO3Vn+omGSM
KGaeTqgnol9SSQvJK6ljXfhYr/hxUvqnC8GOD+GVHUR3VyIQwBxFATnrUOOgkniO
JOrmzx93f8hJ2NggCuFaLZBl2KKE4ou64bS5juY2VpHODIkwVeRn2k/9s3sxnvkm
g1beMMlz+E35xncnYsMD65vIAAww7W5kk3ebN2MvHmWX3kiA9uLfzkvHKZ0D94sH
Zl7nFXccH9OLmpV9hJv/r+W0HnSgvOGt5ku48FgksGCP2h4gWeW165gXcnw/7AdQ
H3dPYuz87TztoFOYxSKyrx0xHuJskySXsfe4hqhI+Dvz0Q8BdxFsN6N+m8RK1O9l
hKsLJocSe+hWPT8/CIPs6QkH7M9cOug0woUZh2o6U7zyeW62Cy+0hhm/kEF3fq3u
I3lZZcKYezprERruj0EnEzaVN2JnYwpT6gH0ZmtcysVjrF2qG2qM+dxaEN4vCVIg
dles8GNOXSnQUTPt/lfuCZ9Xr6o6uQkNqeYR/T2TvHfVvPXh4sM7Kg6tfrGNBzmM
gEwWH1DAI3oB5sJ+dJRe+r6Eb/idTjadSy/Le38k8W/ELbBNxwZ8/HcofHpu2kWx
vkP4teZRT23nvqgf9T2sxw1OQh1txJnJ6paPueFV8Ryn7G6iUYoJgyuUajfi7AxU
1J5r71gVNmqkDMx2wcSlIZ82zAl6XEAIV8GuzKmbSP3YIZ0NYngZzMBO5wQ70AuX
LIgvlVk5CfgCwTEx3xcqrucFX1gxRk2TylFaK8wG+p7OxdfiSAQT/t+GSpWRv/mq
LosoB2oIbhE9H3rtRHTXI+Z6AIZ2LhZk1X5CtdF4kG11z0p4cMQugksWy/vOCmfc
9q2p9Ci3UHqP5yH1iaK8Ls0aEY2Gcsa9cfN58kiZJI5FAAPIKWBCQotkENBWBsuk
ucx5vjXKUcDawnbXcgjGGgX6qK0htEVzgbhdHQ1EEbwCrpAtMB/ESqGVWQBSrsQb
ZwoBIe4KOyUVqClEBbBgc4q6Om1fsnpZhX6LYSVi2dp4rElZ10jn9YMxrzer9KE0
7lxWZGo/dkugjZNGwYyNikoWWvzuzVJovCiGUGK1+OtKoFRF38kQg6tuudyfZNrm
STu6qd3e6I+3UaAlF9JB3/Nh7THabS6XWEPG2sPmjIQQXCHMeYCvcdD4uBClzYIK
L7Iu2Oz9+3Yo1VA/mHk99Fg+9pvEBdgzLCzkmhQyYgnSLulDNSPBizEmQmehixDO
1Z8CtDYyedJRAASnauhpIAIh3CmC5Kpnvd7ZCCj7p0coZHhE9f29A9gesgADVVPE
OtuPDadWXmBLhZbZAk5qzaIHwEwfHOhnOT3PaWzWJEzpL2PMG85oy+1Gqk5QNhkT
wpmP2wKvlytSv3X6+Ewp04SdsYPzzQFVtW2vNTozhP5kcoam1FEyRmfvf98soYxQ
qszz1ZfSU4/0LcsoRPVZxOmyYhmBFBRF5ZzmYmvDFpk9ZfzCzE3FwRQxojVjzwAK
VBo9sMp7gOYYBUX2zCBhuLEKATsKilLBeQFYcXMKvAg2Gwc3RPvnhc3IeWENF5Sh
2zdDO8ZU8zZ7yXKN9Xe+NoIEUyGKJPsMukpjKV4e4xLrbq7N4O7lFfoOIjMBW0cQ
wtId6L4xJz+NcaZ+4CQpjyyNiT/+ESeOb5OVEsWfpOH/c4Sfu3zJDpm9VIObGHdS
zcem2V/wLy378P94DAc0bQX88KpXHkG+KhElPuXYdH5cKir12BawbAuZSQm9TeQT
ncBMCnJbZSavSWRvSZGeK0eXL/M8WxFMll7JSYFgRA3GkkylulRX4m3Nv7cm4kgl
l2qLzkD6Z3ZhfgdZ+nJH/2lYzEkcq695LzS7QwQu901OdM5qCQEFzRYJY+SIEd4w
FMB19s3eFwUs9lFD9QgC7sn4CisvKquJfNVHaJ0y4gNazQWgKTs5qMUORxpSqYYB
40vYHIck6GJ/SOdjLng50JY9YjRS317LBH8ecC8RYS1tW64T0dsimawUG0kVKSMN
onk6KqM3wu6Qpt2w7QzStZ1SEa84JxzCNS9r9XBbCJTPnFG/n5NHqWOrghz16v5T
o86KNQMVnoUUfz1E38sGVP/cfloPoGhZ+o5CtY9eWffa+b6O0zZI9KtuTK07isRy
7R39akJ7apiUNg7Letb5sZ5XDLVl0a8/sTvBB+XxaAN9d6uN0aTMaMgSbQVkIEAk
QxUgwPw07t874CwtoX4khkFd4stiRtkFFVTXuojnbq++AXzJKiE85StINBPT3u2z
KahuC2a21FZd4qPncXAc04Ul5BIOWgfEluBr8wxv/IHUFQt9P1VreR6M4CvtHt6I
joA9TeGt5MIS5N7sqqjOcefSUhLvoWMNF7TuvRzRmcZdv5KkPPrI9FPLRRWStI3Z
6kH4EWb5hPiYVQDK1VKsb7l8omZ4XzvPhuR9BFwWDl3tp73rU8VxEWLpdCfkvv6X
gixhRAkQ5bQOf1/wGb9ifOiXxUUlJZqi/p8D9WBvH3UfnzX5HmyH7F1LqJbu0MLL
sLNzs8s3v5R/DWbBln29S5ZOOAPa0S+IkLcOibl/il2ii0L8ZM/W2iM40wq0Txdl
CE59SgybfoI8/L32vzjVbhezA7PFI5XPEzwGdqAm6AurfG46lt6XMp4ZHP5bcgi+
XRa0LvW7ikQX16b9XTG0JP1JOE0OA1mn3gcHruqBEt1KLpF5EAdY994Ln75u1pau
PCYFwi20CbyA6vF+rpz0B5d9psS8UzuqyBouah54WLFWQW0A4ti2fP+w/nC7vz4C
qUE6k8vKT5ipSSnSq7SzJ+aFjGuKyCASLbnSQVNIs1I0HS7Wrj/Dd4cRAJDj+frP
azOk80HYqW5b70jwzyLs4eoDY6PPqBPxfnDKGWO8lOnRTde4sH5kxyx6F8WN83bL
OD7BnlsK79JkfFqOiL6Hj7dkPxbcnw8Hx/OJQSjbtQ0GrrkgAtXZEjToUt6sGokf
HZhldmdLMrGu4rA0yyIDoVzSXDeA+Q0B/yGVkLXORmFH+nbcAcMaKvjShxqVT75y
g0zVo5u5XOFPh9XTFN/KsudvSnd9SyQy0pn+GCAgpxucez34pjBXYbCECErJ5qsd
CL7MxpVJrg4LvsoYn58sA/kCR2QjkklZkFlO7ZLk7N0B0AFi2pjG0Vqt7rQHiwan
1mfVKa3kWidUtIaLA+rWTMJDXVReUlIr0ChEhKeY6RPbw1DxozUnlam3JDAfkdfv
9mKeLQPWqJrOxK3yDg4nRE1Uja56xQaPpxO0fkF4QE410dJ9/ZOjpj0tnIHIq2nH
Uap8eYckEy+TTaOSBMssZO8vtiBuFIwzKX5Bv32gQCvtp8nbU4M+1m/Ne101smCo
tazHeYmBz53z/vZIvIDENmV58dm3w4n/ytq22qvEFQ6vNcsV4foOBRxEpZ47f2Z6
GRQ0trc7/yxoDO/DPQQjVbf6MFgqc2xnRMmu9fU8KvMRZzSTcM/zDeO+4kk+PtJj
ReOuceB8yir8L7K4v6WJiINUr98vdpExuVcbvGQdYSTKXL8a7hbwdUe1oi9nNscG
sdGUYwq8sn6GO8gp541FXLSK0l734bB/QPstkVJY06Vl5uxDQXBAydOKSDxhauqm
Ll06cGH/X1c07LCdtKziJQQDzaqXmCQn29mOiWpc9FLIvBWIH3X+Rk+s+rDDaK4m
bpVxYCyO6aaLSDHzAXS3AU3pFbxWRHdRTE9bBRa33tHAhlZUL6R0EToPZHcFD0bL
7JUrmawoSa6o/CyYRhTFeJi+KqAJnznBxYfL0Q6k2GE=
`protect END_PROTECTED
