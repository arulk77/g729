`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG47j1YD+lAc7EUQFJD/5C1Ac6bubbjWoEw6VBGM8ekw
yrKnVBk0sti3cUqZL68OJ8fKNpZdxW2pL1ThZia6k1HYZ2iSkFvrRH4hkEWa0bBv
lqeJxEX717E/t2b1SRj0IqYCd9/CZ35vtqImaoR0irfmVUyvfR6s/PLgeaWSxua5
`protect END_PROTECTED
