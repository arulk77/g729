`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDd2Mapl2GFssy2dOJ8lg0DuWw44nvsn17YE1hEotlzR
0uCeIkbJRnmP6CsxnJc7ONTnuALElHHSQaf0CteKXd4G9gREhBDMwguwKHi5HdWb
bcxtOdCqb3VcOXKXL4maUVFagiioQeGGM2y9sGJgwndh6falNnbRcjZcSOZCTEkL
RUUKvqTrOnN3aHHMV1D1ibvmoNtvPSJcRacxEbGHeN1MDhwRtcqlE54c7nEMOo6G
9rXltp2Srpe1wvqhSVp1wOD/V1lTJlOPl/Y2M01A2aIktH9/eBB9u6ZdlilED1e7
JTKZvA1TZWov1NYS/hJ+LuFZDc9/4pvIJUx/FDpgwidB6c5uePD0Ivgq38EuaMpi
b3/nUed57UG8r6wYc0svhw==
`protect END_PROTECTED
