`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wdrmli7LJTJLzjco3q96+CrOv78DkQWs7MjA4/jiz07
SBMLkXorbSzBJIRoe7k1WAIEQPVIRW+v717l+zghWyL9ZKhoN2HoegvqFnJRab0O
8B/lR9L0uqVCq6EG3fqBWIEUiCkq0WPReeLhYqEtoay28/T3u9/V/h1OXonHSgiF
TKeZAIHzkv1gUk7zIR45Ztt0oTBZtxYWg2zrEtLKMuz+7sgsqGZRC3pMd/KYtKfx
atxJJflF5cyRk1AABCes3U8chpaFKFbVpLM+DnFzCTqDJwT1vEFi2SJa+oaynz9q
D6y5l0zwmG+8MpUKrWKPlQfsk+3cr+l6N+6ruD9knAnNpUyGZn5Ay4hbzzvx5PtY
A/SC+eK7b4igLq1O7S5fTA==
`protect END_PROTECTED
