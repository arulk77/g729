`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKW+Fzhf+wdvJoqdIsDKdi165brf5PC2+mX9DjjQY0nT
1rJ8Tqw8nah3j6+LisFyYjisPZW5g7MjqT1/u8dRw/SLgxeasB6q6FD6S21Onqv1
sPNeXuUHto33V//WY9w0dKx/jaztTEmWcTUHzZxfdjiGutAvZ34QR8v2hnj4N1jX
ite+odGHWTbUsgkki7VjwHhpOTBIXmUiRXOzVcoE3Hw+iha/kD6g+iWG5g4gY2PB
2N5sqW/DYuJmWNvbdo2IfHwxbDv3KQR0KdCEP4EGHVQmZ33149RkmSiEX5CyHcka
E7PUq+KCaKJcnAr5o8ywi1gBKh7RiLwQxYTf+XuNFnphfj2j9BOSiK2ZROSHqHnN
xdmdDuEHtPVsgC/1oj3KgqkmimFCca0rkolufsVInUOVVkal3GBRYTaSKNBLsoOM
mY4HZ26BZJ4/VwMp2mCJuw==
`protect END_PROTECTED
