`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47RYx0Oz2hJyj7kiMIZY3YTxYFjsoushYzX7TX+kVCNl
zat3/me3mfeUB/5wOKUTBR0rc9JDDpyP6p8REhOkVQvrHwXBh1lAXmCLdw2i/Hh7
IdMrjqDOjjK+FCbh0YTtwRMwplKa/uZfaWuw8QFSxPE3DjMjC+noUiGTWC2BPkRg
cmwIezUBK7bydNNeoIV2CRKfzrAWuYmJcarb9YZZvI8UeRy20Y/l4F0j+6mEAp81
bi9oOiTNFwzDQHPKOQDZLg==
`protect END_PROTECTED
