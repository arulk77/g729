`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHVw8nfC0t9tB8GYuV3+qTy0ovTCG4KYT5X4aZKI+cBt
mQz7LsMUG5mvIlmnalrGSoP9+1drmzigjoBUJfWpm1B1fqod8s/Rqk9vKyANz5nd
7cHSRmAEK9ecGW6ipSLPrloGLrp9YJZyVqYWq6GpBBAj2o5/I7z/q5JhafN7PsEe
Jdm5XHI9mPCiQIa3M27tZVcY3hVMhiSR1NIvWUbeweOXFG/fWGg2l/gKI7Yfh63F
KLxMhnDUtP0P/y/5eCu23oZuF5Xf3ZPQ3SuoXRf2oC5ij30TnIBX/L7IehYr+cOl
vWJqXClv77qwDKnmK4gT094oGkrNEqs9cyM5cM7THC3Fpu497Yn0wV0jRnvcy8/N
SL0i+aJux0IViCqih6xw04vRRMzSHNUGdAGD422zENSGPpMJZ07F0uNCLknVEljf
FjnojoL838oBVpJaowiPM1G5wEy9638SK1kYDvHPkjw7uhrv5NcQHoMV5WNvJJXX
Bmv4NiM8J8e5waX1XBPFyTEDSmEPXhujvzYtn++/A/E=
`protect END_PROTECTED
