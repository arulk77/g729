`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu488JsT2HJQ/mC/IIUzQvFs1gYfakK4WJKmFMosdJUw/9
s439odA79mfFfc7j4L3dJ3pLtJmFySuom94Gq/9Cw7jZqMOY3WhO1BAib6yFCTef
e1MrA4R8ihATLsc01zBpEZ9d+6FN7et88qOSRLWsOId4jDyaI/w3tdOaAfMifJTe
RL8+AwKl0bgxCkZ4y1caHzXLEae3RXs+0MBMGpykzV4LB4HcfZ+7y+9mwfvGkPTN
CNNGO0vpLR4409kYwbl3OdLIzq5JNP6DYYL7oiuSnVbcJ/S9DAKEv0H92UNHZ2XE
0J/LPF75EOB0ZEAkVF+kVyyBtMia6OgRdWhNo6vJKD/Wee9+B7ZuMs/sqWQP+WRl
rBnyo0KP6ReYuVtD5gkk+w==
`protect END_PROTECTED
