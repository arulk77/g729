`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu471yk39ZOcCa7tlkc4vbu9691nfukAqxe3ha+5hEW/BM
BdMVekARzUhD+pjftf9+5bb22vNKV8xF+pzK7inqWLKeJxtT29dGAcfJldsFRIhq
NZ4jvyBM1UdVKu57tz0P4WNSFBwAq0OdpOBf4L3XkUMutjE8BY6jhR6Jp7562lAn
04OgENFvDiq2ByuRCJDH6R7l6dsuAVgdxZvCCas4PbtxjUBmU0qfryjvWRS2dll7
C/xr14PjauZamXAzshTPqp2G2yDuHLEm7dcUNQFZnrA=
`protect END_PROTECTED
