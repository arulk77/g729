`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4166DNNgal/mP8BKp2zzVlclJUA94UgHa4uiS5rkgFDM
nprdX6PHr+4xsKrzqkqzgoaxTV71oIpK6T16JQQUBwjPT59axeNYoEE9Sbz6PcpP
gMY0vf1XCFECM0QT6uZXaJKp8+EaQ6N2iiNloHshgm52pBURlIfG9hKL8j788d3t
tnUO/Qy5g2ZF46Rdd/+7wQbpqqDkttPUmMABuvVhRYg=
`protect END_PROTECTED
