`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNag6lIXiGjwVa5vcBv83dLFQRhcO/0OIQSGvpbxo6hK
5WLnu8NO+L3DUNQDoaBqNFo+dtvqPcfQNB1knCvsLbH8fJTB/P1kVjlGxpjdMOyE
ElgJFzH1hncV2r+55Usi9+EpTEK9aQPWKLJQY1WsDxAGscDt44W/ModvVVn0dX5i
DPv6a1bDlNR0H1L00lji5pd/bcSLG9ImxMYH28yxCMVitm/AthAEM/Hh5CAesK+O
LrRAszTjQ2dF87LCmUW5qCYyiFeisDkjxO3H+AsbO95n/UU7/AYm8S0NMsNOkPAh
asRwWisIo0t7MTnLG76E/Ql9uulrQidx5YrjooPr4bM1LU7zi+bdsTmbwf3jJ3G3
GWlZ6F9CirB5dRgF+Ax5eA==
`protect END_PROTECTED
