`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF2O+EOq4P5ujhFo+gj5YDACYtcI9+fOV5s4/79cLqYZ
W7f9cR/wC8Hh2s1wiJQU2nPJ1CpNqDcNup4+X7uH8ZPEVzt3h/8PXcNyL5jeA92w
w4CMbdF9AVUO3NIowwHwMXdMarfp3nB/uUXJfXEfIA80g5dOVUau8hrBJZjOFIzd
eMKW2Z82jX3QuQeJyV7v7UXKV4PUc27KYl/TIID4+/piTylybfd3HG/S0tkW9xoP
`protect END_PROTECTED
