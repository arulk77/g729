library verilog;
use verilog.vl_types.all;
entity PCIE_A1 is
    generic(
        BAR0            : integer := 0;
        BAR1            : integer := 0;
        BAR2            : integer := 0;
        BAR3            : integer := 0;
        BAR4            : integer := 0;
        BAR5            : integer := 0;
        CARDBUS_CIS_POINTER: integer := 0;
        CLASS_CODE      : integer := 0;
        DEV_CAP_ENDPOINT_L0S_LATENCY: integer := 7;
        DEV_CAP_ENDPOINT_L1_LATENCY: integer := 7;
        DEV_CAP_EXT_TAG_SUPPORTED: string  := "FALSE";
        DEV_CAP_MAX_PAYLOAD_SUPPORTED: integer := 2;
        DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT: integer := 0;
        DEV_CAP_ROLE_BASED_ERROR: string  := "TRUE";
        DISABLE_BAR_FILTERING: string  := "FALSE";
        DISABLE_ID_CHECK: string  := "FALSE";
        DISABLE_SCRAMBLING: string  := "FALSE";
        ENABLE_RX_TD_ECRC_TRIM: string  := "FALSE";
        EXPANSION_ROM   : integer := 0;
        FAST_TRAIN      : string  := "FALSE";
        GTP_SEL         : integer := 0;
        LINK_CAP_ASPM_SUPPORT: integer := 1;
        LINK_CAP_L0S_EXIT_LATENCY: integer := 7;
        LINK_CAP_L1_EXIT_LATENCY: integer := 7;
        LINK_STATUS_SLOT_CLOCK_CONFIG: string  := "FALSE";
        LL_ACK_TIMEOUT  : integer := 516;
        LL_ACK_TIMEOUT_EN: string  := "FALSE";
        LL_REPLAY_TIMEOUT: integer := 1549;
        LL_REPLAY_TIMEOUT_EN: string  := "FALSE";
        MSI_CAP_MULTIMSGCAP: integer := 0;
        MSI_CAP_MULTIMSG_EXTENSION: integer := 0;
        PCIE_CAP_CAPABILITY_VERSION: integer := 1;
        PCIE_CAP_DEVICE_PORT_TYPE: integer := 0;
        PCIE_CAP_INT_MSG_NUM: integer := 0;
        PCIE_CAP_SLOT_IMPLEMENTED: string  := "FALSE";
        PCIE_GENERIC    : integer := 0;
        PLM_AUTO_CONFIG : string  := "FALSE";
        PM_CAP_AUXCURRENT: integer := 0;
        PM_CAP_D1SUPPORT: string  := "TRUE";
        PM_CAP_D2SUPPORT: string  := "TRUE";
        PM_CAP_DSI      : string  := "FALSE";
        PM_CAP_PMESUPPORT: integer := 15;
        PM_CAP_PME_CLOCK: string  := "FALSE";
        PM_CAP_VERSION  : integer := 3;
        PM_DATA0        : integer := 30;
        PM_DATA1        : integer := 30;
        PM_DATA2        : integer := 30;
        PM_DATA3        : integer := 30;
        PM_DATA4        : integer := 30;
        PM_DATA5        : integer := 30;
        PM_DATA6        : integer := 30;
        PM_DATA7        : integer := 30;
        PM_DATA_SCALE0  : integer := 1;
        PM_DATA_SCALE1  : integer := 1;
        PM_DATA_SCALE2  : integer := 1;
        PM_DATA_SCALE3  : integer := 1;
        PM_DATA_SCALE4  : integer := 1;
        PM_DATA_SCALE5  : integer := 1;
        PM_DATA_SCALE6  : integer := 1;
        PM_DATA_SCALE7  : integer := 1;
        SIM_VERSION     : string  := "1.0";
        SLOT_CAP_ATT_BUTTON_PRESENT: string  := "FALSE";
        SLOT_CAP_ATT_INDICATOR_PRESENT: string  := "FALSE";
        SLOT_CAP_POWER_INDICATOR_PRESENT: string  := "FALSE";
        TL_RX_RAM_RADDR_LATENCY: integer := 1;
        TL_RX_RAM_RDATA_LATENCY: integer := 2;
        TL_RX_RAM_WRITE_LATENCY: integer := 0;
        TL_TFC_DISABLE  : string  := "FALSE";
        TL_TX_CHECKS_DISABLE: string  := "FALSE";
        TL_TX_RAM_RADDR_LATENCY: integer := 0;
        TL_TX_RAM_RDATA_LATENCY: integer := 2;
        USR_CFG         : string  := "FALSE";
        USR_EXT_CFG     : string  := "FALSE";
        VC0_CPL_INFINITE: string  := "TRUE";
        VC0_RX_RAM_LIMIT: integer := 30;
        VC0_TOTAL_CREDITS_CD: integer := 104;
        VC0_TOTAL_CREDITS_CH: integer := 36;
        VC0_TOTAL_CREDITS_NPH: integer := 8;
        VC0_TOTAL_CREDITS_PD: integer := 288;
        VC0_TOTAL_CREDITS_PH: integer := 32;
        VC0_TX_LASTPACKET: integer := 31
    );
    port(
        CFGBUSNUMBER    : out    vl_logic_vector(7 downto 0);
        CFGCOMMANDBUSMASTERENABLE: out    vl_logic;
        CFGCOMMANDINTERRUPTDISABLE: out    vl_logic;
        CFGCOMMANDIOENABLE: out    vl_logic;
        CFGCOMMANDMEMENABLE: out    vl_logic;
        CFGCOMMANDSERREN: out    vl_logic;
        CFGDEVCONTROLAUXPOWEREN: out    vl_logic;
        CFGDEVCONTROLCORRERRREPORTINGEN: out    vl_logic;
        CFGDEVCONTROLENABLERO: out    vl_logic;
        CFGDEVCONTROLEXTTAGEN: out    vl_logic;
        CFGDEVCONTROLFATALERRREPORTINGEN: out    vl_logic;
        CFGDEVCONTROLMAXPAYLOAD: out    vl_logic_vector(2 downto 0);
        CFGDEVCONTROLMAXREADREQ: out    vl_logic_vector(2 downto 0);
        CFGDEVCONTROLNONFATALREPORTINGEN: out    vl_logic;
        CFGDEVCONTROLNOSNOOPEN: out    vl_logic;
        CFGDEVCONTROLPHANTOMEN: out    vl_logic;
        CFGDEVCONTROLURERRREPORTINGEN: out    vl_logic;
        CFGDEVICENUMBER : out    vl_logic_vector(4 downto 0);
        CFGDEVSTATUSCORRERRDETECTED: out    vl_logic;
        CFGDEVSTATUSFATALERRDETECTED: out    vl_logic;
        CFGDEVSTATUSNONFATALERRDETECTED: out    vl_logic;
        CFGDEVSTATUSURDETECTED: out    vl_logic;
        CFGDO           : out    vl_logic_vector(31 downto 0);
        CFGERRCPLRDYN   : out    vl_logic;
        CFGFUNCTIONNUMBER: out    vl_logic_vector(2 downto 0);
        CFGINTERRUPTDO  : out    vl_logic_vector(7 downto 0);
        CFGINTERRUPTMMENABLE: out    vl_logic_vector(2 downto 0);
        CFGINTERRUPTMSIENABLE: out    vl_logic;
        CFGINTERRUPTRDYN: out    vl_logic;
        CFGLINKCONTOLRCB: out    vl_logic;
        CFGLINKCONTROLASPMCONTROL: out    vl_logic_vector(1 downto 0);
        CFGLINKCONTROLCOMMONCLOCK: out    vl_logic;
        CFGLINKCONTROLEXTENDEDSYNC: out    vl_logic;
        CFGLTSSMSTATE   : out    vl_logic_vector(4 downto 0);
        CFGPCIELINKSTATEN: out    vl_logic_vector(2 downto 0);
        CFGRDWRDONEN    : out    vl_logic;
        CFGTOTURNOFFN   : out    vl_logic;
        DBGBADDLLPSTATUS: out    vl_logic;
        DBGBADTLPLCRC   : out    vl_logic;
        DBGBADTLPSEQNUM : out    vl_logic;
        DBGBADTLPSTATUS : out    vl_logic;
        DBGDLPROTOCOLSTATUS: out    vl_logic;
        DBGFCPROTOCOLERRSTATUS: out    vl_logic;
        DBGMLFRMDLENGTH : out    vl_logic;
        DBGMLFRMDMPS    : out    vl_logic;
        DBGMLFRMDTCVC   : out    vl_logic;
        DBGMLFRMDTLPSTATUS: out    vl_logic;
        DBGMLFRMDUNRECTYPE: out    vl_logic;
        DBGPOISTLPSTATUS: out    vl_logic;
        DBGRCVROVERFLOWSTATUS: out    vl_logic;
        DBGREGDETECTEDCORRECTABLE: out    vl_logic;
        DBGREGDETECTEDFATAL: out    vl_logic;
        DBGREGDETECTEDNONFATAL: out    vl_logic;
        DBGREGDETECTEDUNSUPPORTED: out    vl_logic;
        DBGRPLYROLLOVERSTATUS: out    vl_logic;
        DBGRPLYTIMEOUTSTATUS: out    vl_logic;
        DBGURNOBARHIT   : out    vl_logic;
        DBGURPOISCFGWR  : out    vl_logic;
        DBGURSTATUS     : out    vl_logic;
        DBGURUNSUPMSG   : out    vl_logic;
        MIMRXRADDR      : out    vl_logic_vector(11 downto 0);
        MIMRXREN        : out    vl_logic;
        MIMRXWADDR      : out    vl_logic_vector(11 downto 0);
        MIMRXWDATA      : out    vl_logic_vector(34 downto 0);
        MIMRXWEN        : out    vl_logic;
        MIMTXRADDR      : out    vl_logic_vector(11 downto 0);
        MIMTXREN        : out    vl_logic;
        MIMTXWADDR      : out    vl_logic_vector(11 downto 0);
        MIMTXWDATA      : out    vl_logic_vector(35 downto 0);
        MIMTXWEN        : out    vl_logic;
        PIPEGTPOWERDOWNA: out    vl_logic_vector(1 downto 0);
        PIPEGTPOWERDOWNB: out    vl_logic_vector(1 downto 0);
        PIPEGTTXELECIDLEA: out    vl_logic;
        PIPEGTTXELECIDLEB: out    vl_logic;
        PIPERXPOLARITYA : out    vl_logic;
        PIPERXPOLARITYB : out    vl_logic;
        PIPERXRESETA    : out    vl_logic;
        PIPERXRESETB    : out    vl_logic;
        PIPETXCHARDISPMODEA: out    vl_logic_vector(1 downto 0);
        PIPETXCHARDISPMODEB: out    vl_logic_vector(1 downto 0);
        PIPETXCHARDISPVALA: out    vl_logic_vector(1 downto 0);
        PIPETXCHARDISPVALB: out    vl_logic_vector(1 downto 0);
        PIPETXCHARISKA  : out    vl_logic_vector(1 downto 0);
        PIPETXCHARISKB  : out    vl_logic_vector(1 downto 0);
        PIPETXDATAA     : out    vl_logic_vector(15 downto 0);
        PIPETXDATAB     : out    vl_logic_vector(15 downto 0);
        PIPETXRCVRDETA  : out    vl_logic;
        PIPETXRCVRDETB  : out    vl_logic;
        RECEIVEDHOTRESET: out    vl_logic;
        TRNFCCPLD       : out    vl_logic_vector(11 downto 0);
        TRNFCCPLH       : out    vl_logic_vector(7 downto 0);
        TRNFCNPD        : out    vl_logic_vector(11 downto 0);
        TRNFCNPH        : out    vl_logic_vector(7 downto 0);
        TRNFCPD         : out    vl_logic_vector(11 downto 0);
        TRNFCPH         : out    vl_logic_vector(7 downto 0);
        TRNLNKUPN       : out    vl_logic;
        TRNRBARHITN     : out    vl_logic_vector(6 downto 0);
        TRNRD           : out    vl_logic_vector(31 downto 0);
        TRNREOFN        : out    vl_logic;
        TRNRERRFWDN     : out    vl_logic;
        TRNRSOFN        : out    vl_logic;
        TRNRSRCDSCN     : out    vl_logic;
        TRNRSRCRDYN     : out    vl_logic;
        TRNTBUFAV       : out    vl_logic_vector(5 downto 0);
        TRNTCFGREQN     : out    vl_logic;
        TRNTDSTRDYN     : out    vl_logic;
        TRNTERRDROPN    : out    vl_logic;
        USERRSTN        : out    vl_logic;
        CFGDEVID        : in     vl_logic_vector(15 downto 0);
        CFGDSN          : in     vl_logic_vector(63 downto 0);
        CFGDWADDR       : in     vl_logic_vector(9 downto 0);
        CFGERRCORN      : in     vl_logic;
        CFGERRCPLABORTN : in     vl_logic;
        CFGERRCPLTIMEOUTN: in     vl_logic;
        CFGERRECRCN     : in     vl_logic;
        CFGERRLOCKEDN   : in     vl_logic;
        CFGERRPOSTEDN   : in     vl_logic;
        CFGERRTLPCPLHEADER: in     vl_logic_vector(47 downto 0);
        CFGERRURN       : in     vl_logic;
        CFGINTERRUPTASSERTN: in     vl_logic;
        CFGINTERRUPTDI  : in     vl_logic_vector(7 downto 0);
        CFGINTERRUPTN   : in     vl_logic;
        CFGPMWAKEN      : in     vl_logic;
        CFGRDENN        : in     vl_logic;
        CFGREVID        : in     vl_logic_vector(7 downto 0);
        CFGSUBSYSID     : in     vl_logic_vector(15 downto 0);
        CFGSUBSYSVENID  : in     vl_logic_vector(15 downto 0);
        CFGTRNPENDINGN  : in     vl_logic;
        CFGTURNOFFOKN   : in     vl_logic;
        CFGVENID        : in     vl_logic_vector(15 downto 0);
        CLOCKLOCKED     : in     vl_logic;
        MGTCLK          : in     vl_logic;
        MIMRXRDATA      : in     vl_logic_vector(34 downto 0);
        MIMTXRDATA      : in     vl_logic_vector(35 downto 0);
        PIPEGTRESETDONEA: in     vl_logic;
        PIPEGTRESETDONEB: in     vl_logic;
        PIPEPHYSTATUSA  : in     vl_logic;
        PIPEPHYSTATUSB  : in     vl_logic;
        PIPERXCHARISKA  : in     vl_logic_vector(1 downto 0);
        PIPERXCHARISKB  : in     vl_logic_vector(1 downto 0);
        PIPERXDATAA     : in     vl_logic_vector(15 downto 0);
        PIPERXDATAB     : in     vl_logic_vector(15 downto 0);
        PIPERXENTERELECIDLEA: in     vl_logic;
        PIPERXENTERELECIDLEB: in     vl_logic;
        PIPERXSTATUSA   : in     vl_logic_vector(2 downto 0);
        PIPERXSTATUSB   : in     vl_logic_vector(2 downto 0);
        SYSRESETN       : in     vl_logic;
        TRNFCSEL        : in     vl_logic_vector(2 downto 0);
        TRNRDSTRDYN     : in     vl_logic;
        TRNRNPOKN       : in     vl_logic;
        TRNTCFGGNTN     : in     vl_logic;
        TRNTD           : in     vl_logic_vector(31 downto 0);
        TRNTEOFN        : in     vl_logic;
        TRNTERRFWDN     : in     vl_logic;
        TRNTSOFN        : in     vl_logic;
        TRNTSRCDSCN     : in     vl_logic;
        TRNTSRCRDYN     : in     vl_logic;
        TRNTSTRN        : in     vl_logic;
        USERCLK         : in     vl_logic
    );
end PCIE_A1;
