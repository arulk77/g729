`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C/d5VNCd4Lhwm2ktOUajO6sAU5OLiG3iDXHUDqyHfL6s
UNQxRUyfwVcUEqqxr5zcH1HU6HBDQr5BPTec54I+o4NNB77saUIjzF3UDlTzmo0x
tf8DVBC+xYbip0tDmKVZQlCY7Gq5rjC6H95AxfV0JDrRVWc273jwGb5wz15CLtFL
MnIg+dlgfI6sEAY3r5LL5OQc0n58gRLc+X/OMbWpC1kMrKa3o4VdWZhsWNpPF3BQ
CFgJA+ttRLCeABzS0a/3AY6ZDl8ffQ8buBEs8AOqgcNhfz1hZdJ7FH4bFAPZ3EP9
W/u/RCE3YMK7MX4oAlWrVtUyHpYT6vIBENhjnwybYVLKltJdyUIeSat6B9pKl8xU
co1kLDRFx7VqSM1/Kc2uQk1yYYwWGEtfwO3QG5sfULn9VYcdvHTmxvrSgBb3D6ob
a2yvMlsJDSJyXWnyIvH+Ws3J18VsQ9Im0RVIa3FmRpfqEhrQiOaPi9RKmAZcyzV+
i4DYStVSEgtq9it9rL7dyIh2fuv4RhnNLk/WdQtubNvBAZI5X1+Bgsv60wk+ICty
+Vs5YlL+6Q8UjswGHPgbUzrhrpDLzjxNWxK1ilvgAj7/9f3wOug8vkhWEjALFdL3
vrIdcXHSHWYZDwydloJ6SO4arfJi6Tf3OGdm4bIDNtHj+VeEbum5pzuMBGhgiuXn
xFuVoh4W4R6qeBdP5kIp8A5L7aBjqWdWgVBJ2++t8g5zozZvV+1+362eyvB/aZ2E
yckkAveXQlMoPj+++3E/t/NQobSNhGHZ25vyS5K/wQ744l2ekcEgBr2EAFQ8HHAb
5NQOTJtzHO5KKUqxppn/Nl/LmM4yccYwo/1nmyQfGbQuekVUA/dmMjODuOgDWsvr
zM43dPUK2NGMqpbKaL+gn1DOtEL88F6BNAahZ2EXO4HNEky0fpTCcZmJdkaE9ItP
csOiR4ALk3y/4fObgj7GV1KZmG6xhTvlEdFDLiHYFYK8Xh+6npBK4QOquqO3Gc9K
2AtlRhWCj4ngDu5gBD+IJ+MkiGEjhQWGyCOH/FIG0LgFF3vu/1AYO3UDvi7ZucFi
JwS7TffppHQyAcZhgBmBIF5bMD3zJjzy1haA7ZRJylmmxivw+6NgzZZXrRxKRnyj
0k+9W67ER5GEkAY5KOt+OYT+2bS/SiWn8wE+CpePPuZcgjiFCQ+3Xw71E7XZ0dMH
qtBmcB9a1Qx1rEuQuH//VFWyvrsQ7Ve6dGn8Ri6+WufozC+tAkIuxZfQmmegPhUS
lxKBgRszM8o+WBKlQK6ER40a3GWuiKNZQI7HBQSVZeYlr0QcfZ8Y8bddanqVwFGg
Wfr3hVQRGTMDy7S7XlcCWZjqCK5M02gyPM0VwzJJpQbp4T90rxJSC9HDCWYqXRcI
e+AamSmyJtN+WB8sG8qEOTYbbdzmsnpJamm0cRa+FTnUDCC47+O/FUmK612zV+29
5lyzhSqRMh2FfuD+vpafYmOlU7Yb31MZPdEvRiKXPLC5iIoqmwfjcYJftV0T8PAj
D6q7Eb/que5HZz2wYw227zxNXKhN3bM4DZBXNlXk6yFMkpvCyEqyUsrZ/OaN6AIi
VekQGOfphn4qNC+nXZCVcCiRcDxIs2UFAYqYRCF+wN7daT0ZvuTiPhR1P9OfXGKr
NQAPvaZQA53xQMLxWxuo9X6sLTM9rC9YCqMYnMg1U39z6nYseYT5DxOwnmh+nX6I
VvKg6i2Ypqd8rQ11R6Sg/q050fbwi1FsZmACGukh2FmurzNLkLR4EUtaiaEYsL8O
dKv5EQUXY+G1PVfsTnGtLX5yA8z2FuQTKTPN4BXiD2peyr/zcLIjhZ4C07TGPd59
qfxc/v1FWi8YdqBGGgUbwfZZOD5UQSO3cm4ZsheaB8pt/5u5ZRn1rBxM3FxSo0RG
cEji8NG+a7np04zurVukOkoeRz15klqg6Lfzrlv4lrM=
`protect END_PROTECTED
