`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
rmkKrAQuSppLwL47Z4ST+8TusEG8kJ1S7SNjjWYZJjA3ugDai1wLoLamG2dONZXD
Ky0AonM0WDQLo3NvP3hfraBswcpMlWA07LwjiBKt9Dd+Kqw4Wj+Rx2j+tQmZ9FWE
OargeMZbeXqND39EQ+Esbh2mIjxs9Fx4kagEeU7xJoRiVxENF8HvenNtrmy9bKzP
mNAntZN+xTT3O0j2d3q96Y0XE4Y9WvYH5MgrJ1gFA595qvKezt5wyGqUa4hhmo1C
PlJs6u6mIgrWSrLLvDUhfcgbBzcif5ONwHGrHremHkY=
`protect END_PROTECTED
