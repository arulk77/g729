`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
OjxKa+7wxg82okWXvG0R4SrUwt7GMgX9Bxrdd/r7S4TIChlmRNDEBDY54WoxEp5a
g1u6bCcHRgB864JwpnFVBEokOfG9y0jP0XPAvwe4/dhxreVsD92FB4OC4BSSqDK4
dEdB3Ee6dvYFcLFWmGeobh0kn/wVHDe/zvu1CnUkAA8eMJ9sSfeC2klWdDsjhWp6
mAognEbmExedHZvL7PLC3yf6o34iYmfgFKTWnaM6tL9T/mLYHepbfXX+tNCwygY0
Tk5dvJcRDRP2YeTxkjl57/LFp6sMRY/6u5/U9PHEd1rOPzKL9ogkjYAw+pToIBiw
TZ/HHzW4M2fffiwzLAXmYOCu4C3rejZzv4sSKUlcvlnLWx5wPlJKnJuKEKwZdCbe
XjTxOWupns+Ry2jyy1vdiSYRRs1SBU13+Rqh/IKefnC6ellZfCIcgpb7foKQhYi2
Ef1kpDahJazBKI6HnRW0vyPLvB8DcDNGZyymJS7X9EOTvqmk4xJ6erjhj5P1nEus
+ijE6IBaGVfvlmq9LHZePsTSbVTlvep9aU1PJr5Bb1qGeQ1KUO+uhUkhWfY32M4Y
2l5slXKuyWCc+TWsxwMBcal4EQKPO/uLd06yWvByuUdwguHOatZgFsBinoUfu3d6
Xz3DFqlB9Cle6pbTXzhHxVmf4hmylZnCRuR78elg4CsM4+rXP3/NzZ9iWbnJz8BA
HMgPKHcXaxV8TAn/fADtMaayrWXVv687sBC5J23IHSX4tNLMA3gxhNVZnPlAlDf5
V1GyrkjG61ef/WYueUCtdT8uoD6/nOOMSd8aDM14i/ZO8GPKkHFM0KaeWP/u5VlH
GMHA5chsjWxz6gcEhQhLyAkEBvUBE3wOU31WtbsPoqbg8kC/ioqkXJZ6yQUWBb+j
fz4ObccOwmuNR6YsOv9Qstc0CbXRVfZVvi+vXTQ+AWTX88TAv858+XcL1Gsbsya4
eC1YRZiXE+MM3eFV39i25eT6fwjyeFkKzk6GUA5kBVdq5ddJCSck6jhcZbo/v/O9
`protect END_PROTECTED
