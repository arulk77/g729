`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xrrWEdemImoALHuUBnb0qTRH0oGrde8eUqJEfX8fxrD
hWfH9powtrO/qy2Hy1fiR5kJB8MUwgc664MUOVuUxg3UsQOze7r9eqGQvks5moIZ
tEwNiUGjkZg5jfGwPOqreFdQJKPVoetUxpGH4Kq9MGqYwtPQIT466kTYS/RP3HiL
bln/zUMf3xfo2FbR+MOc4WHjcLJ6CVfczMckr8G8nsQdgUWN8cWLfIa5Bluvijxc
6+a/bw0lvalSXmJmTDMC1N1+yQNVQ1k2bdFQ1C2N1kistJjQoWV8FPO7fMxDV4Dh
VEps/CBlJYkeIcBYWwZYro7NfufAUFt5LrfkPoTfvhkM8rYXjXmeWJyhu7OqkzP4
T54qyNY739j9RBllvOJX6BD/cGvKd+G+gXs58S0cpQAuqicjR0TRWnjclOj4PcQD
hC1dZQeu83R3ULX8s6Yq4w==
`protect END_PROTECTED
