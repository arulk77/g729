`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL6iyGrHlGTd4FRJDbHt8NkmAJ+L9iYdFkqipMl4Z0cF
ZZ2SFlCNINET4DF86q4ehXdE4IQrL5NmV3meHwBQg6Rk0Y9mNDlq8y/SvRPctq1O
VwusZ1UiHpkgnW6h0O5LSfVFHcMWfHHi2UGyghULqib6Q8eQeTG2a8Kr1Brk6lCM
v5WcPsi6QEZmxiVXdv1E1E7QZvwhWD81gDaIn3EgeCN08RsHSO4iq2G8b+9pbKo9
2n3GuTnkOHGUVxHIuHm8MBPb3vVxMvyMwP1wC2najy6g1MKAg3PTGKSUM2ABbb/X
Q8TY0zKZ2IejElidBEZ/IA==
`protect END_PROTECTED
