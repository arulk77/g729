`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C2M5Gxk2nBSq5HylROQYP0IyopF43rJQmMlOrN681K9W
0uPi0RElIYJGtORTOkUFs1q3xaSdpA1BzK613Q7itin/I2UqO1QXHuf96BBIBQsU
JQGVhuqbmoVqgcRtUOlR2SPsnaotSbvVwxGvyGOEyxjQ7Oa5jtmMIBUu3hn00zmO
QAvGRSl3mHcSksHW5NDQbe7spxqp2J+/99bGhp31DWB/j7tRDXjB9N/gymD+lj0j
Sh8uIWZfcPg1ETl2OafaDRRmhT7LXYsrjCHFd+TaFkm7g7AkYZlLKOh31hGmBFcN
ljhVinpN5wa9JN1Or1hKoUERxf5vvCWVk0QHY3jukXYPdIlBtEAP7nOV1oxLRtIZ
Le+zB60jL3k29OL9nf9iRtiDlrMeW2kthmiZcytzunkb4rZcfAH2LBzm1cM1ThdX
q1YvHg5wzlJ176h7F/CVqhqQfnO1YW8cyjDx0YNCNiGHfBnjLrWaZzgNSQg4kEjW
LF/ByxPBoVcRzDRZF5DIogYQagu0YoNOCy97nLGdO1E=
`protect END_PROTECTED
