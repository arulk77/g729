`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wz1EKHKbNNFx1MdJYi0U3ICLF7+5bEnj0SQ9UDOAgOo
ZWArcd6lJF9HL1Mbs1lNFsOpmawQsLwgHePNZkT4DZo3UYj10okSA9bE1VIhOHJl
T81phiBstSG7JJ0CZV61YxH3kZvS0n+b59+9Tb66tOx/agnKnweVOf66JyablujO
HtmeOc/ZwWhiRJdxxYWVGEXXfZiOHy1eAHKqs+AxNqdGdQXGOf7ughT/BFjqozJm
hN2gFFdSgt45GefssFA46vLiHY4tDcSo5Ezd+JP3L/TXkKqhAMQPD6qLRlGqg8RN
UGqrcR7wXQEOOob3KTEdoAUdpeM/Zi2w3fPfUQcbdbV7MNVekSk76qTStaJfY9pX
Zceur4JbheeBhAEpwRnAy7wgCHzDnMlVyeiIQylYRDUrJlTFxSCeEZYy5MQpKGKy
47eD2+NPgFPNkwhKW4Zhvt1VmG2p8LhzEAuPsIYEkwu20zlqHcGDNHJI1o/BbqzO
hMJmFJ4cssmTyW4mhh2AB5CJKqpSCBHnygSIseJ7V5U1kDVLbQvNbGL+dYqbLyuz
CGFzAoe9v/U7pyrL/gwvxjrp7Yrkcc5DYSrYo97vcaJpWtOu1ydv1RnnqwJW03L5
/TlJUOBUy5eRUwGFLYjAtMd0sxZmHBw2WWyN3UPD9hoMkEzf61C57n+rmAQQlcOa
ArZBWdv7PLW0k/d6NnL4otLgE9kOwtvLLRz/Rs/ZJBTu/3WYcF7FIp54yuCFlGWE
RMt2fpx/TXR1ffzEKru75MZVDbb0ZM0e6BN8CRxMk3MXAXeh/SLCb88EecRnMGya
ty/AncCVYIXpMQNwwfOtEBPD5k4mQTdoTFB3Bv3Q/4n5zdsXneogT/QaNzmqRQI9
EoD73zvCmWFT84u/U7CHE+x2Tss0I+SwYDFliTBOiRDIcHiN7ikmJpNbPbSYIRCc
VLgmIJurxpYoOxRqJzap1ZUYmNJPqrXwUwockOzvxI6oPq3zqoKCjR1hqnbUb3W4
8E45fEVbeItPyfo1J5FjSg2zboGsJ6Pkx8+gBMbukbTvHbAXB1lQsD26HX5cbU+j
4Ih9shVYCtMTXpSmDRZInbn7gxP9oh2uD/jfXOSiKbzVmwjqv3Ou6CppFm2gZrhS
KuSjLja2KkQHFZyH+R50Xc6mOakPFua255ACHREHG2LOvzXDMjcXv8GCaVKIh4ON
AC2fh8amyCfT6/M6wWckxXmGbf+PEsIPISyyN9nIhg9/isJ9AyKxss/5NiIfMPYx
tbOTg0GAio1HFQJk7XfjTHLtJZB3nmf1flD+yfjr8+QXuAActYKpaWHw5dGNTVGH
yYgo7reuGNo9tDvAEWD4lsxfienpbamMpdpFqiHdFpjUdS12xTtu2u5P2lye735B
tIgSDBs4E5IghFkAoaZfwUpZXCf3sWRO7bp+94nqxGBB9WARn9G0GRdFw6wnh2uV
FErZ8Ty+bPHAAT03yeb11QiBqs6ZRHj5HLiOS+26R0uFbvSjTOw1WrO6tK5CDPnV
iAxwjLmpdq/HmlHPyyng0y0gZrYeVqSUIAfFcFPFgI9i7wQp/71+0h19Zkvua1WQ
NG1x5RbgDKoviAAtlIqfZioIUlz5A69BXUnhRbOA9xox3B/g/PUjRFqKA0jm61Nw
UOsHB5rb1zsmPEyNvVgmqFbc0HboPOgeIZNBsAW13//L8Tx3CQ079JBPTLTO5ooF
4+V3FNOsIICn/xLb5vtmEK0fzMbagj9y/1gbu87MjPSreCYZTOoUPxgGe9jiKYvL
nOJ6ZkflOM0KVVbhDDMPxQROE/SUqdoHYfDv3QzNuTpz5fG4GNiq1NOeVvYxveUj
GvZUC0TieXv2ttkQHh7lqXIFc190Ut4XBOB27AgJgf/b1X6EeArC8+38pN+aYkBU
lj92VxjoVGDcxXyxEd+j3iArczVsTUOAkXSrhnNA9sNFj0bK82AtToQAnl8mIkA/
6ZE2Dpj7IDY1zrHjU9/YvdlzETVWERfGywd8tB0q/LXd6bRef7Fgr4qlThoAoXV4
UHrgOE8nQSbUTnuaIMXNhkAE2Oer6bdd+zwlaR926+pKITA/3csHWeeqCw2VJhPE
02YxmW/irxM2r3ZzghOVqaHijNP+OED00Pt+eTSr3PrnuWhWGzDzFa5YzWE4MWAc
/rMWTuk+UrJC+DUN+sw+Z+LxT6Nma9tYNahK1W21BhqjQjtHGmnmKIipHNuvYphY
htZ8DhHr7dmxMuv7CZAgDAiCDNYW4MyQgZYjPOq1LvjWGWhvk8cN8Rfyj1KFPeuq
zYFd/P/MfULnQRbj8z5eTqlC0xJ/1aiTCLjacVuqX+9govR6+85uEBzIp/1Xf1BW
8xsCBKyQadvWHyw1zcogo2p+FUmd9NX82kGMTVw7JOp3MX/EyyJPrgwZVhLRA+vH
okT4BLZwcfzjH3wXFQt9runyOKuqN9TG7JnFLblvRAq5fNKYLqbuPXAEz0naEFhP
W/24E01lREHXEGM2wyhKIm2HljDiA2NAq1LFv4EKPL6AngTepNI6MxeBjChN3vDe
jKrMBQVhf0L7iP3Pz9qWh5crObRqxkt6C9oczuG0Ma7D7Naj822jioxU1zE7hya1
CwZcbZpazDTSjtfqoepSkGBM0DMXhhIi9ghUsvIm5SDDHQeBNtZVqpplvkKe4/Ie
dwObxq6CQgVEKpRyLa5H/oydMetCk/9YUIHrDGcttY4RVjRgV8RUYdsZcC8CrAuw
I40qA4lPanXaIJqz0YZMhdkLEasRV9VWhv38fSFdp3lZO7kSRhzUEdwxiUVNNAMG
iHRtvfMt/f/QNTd3CaFAHanAMK/sqdkdiv+kOBNjVrNqeUHg/cEQFdK4/sgNb4ns
/NyNwoJTD9OZ1/J8A4migNqWL+E4l8/2H52AT6MbsZSgi0K6mO3ZvjSeIGLUBTQs
cylxdLncrQS035laJkRsVy0GAypUem+UMJiKDrpwuOWh9d0Nc7Fuz2q/SFMe7bRw
KqQdNf0yvhbTrH7jwEvTMA3kii3XPxRg57JS1GqIZg9JIA3CixL4aJiFCcM+WSft
fWxWquATgozgcFBmDz0BGm1rWSdGVNkJhLzTjeAMapRwTkxOA4Qr0pD6HeD+IGON
MrlII/Q75p00+n6Tu/Z7z6pLnEm8OvVyJbmpWSvtV6yk3KNK1I+LwK8CmBfuaTEs
R48jQ+mMlXnvyy2KT8DrEuTHrVdqO+lq04O5mRDPOOFqowtUS08JiD3TB0+fu/8r
qGiFqNVlrDLucHo3Lcb5mMS0KL6XDoIdj/aFQwjfw55kBiL+7WMNUkPXA+4AnHiI
B5ru3XQp5myyQuZ/bGgccxnUIwPjaCPpHbsZ/rfSGx13pOjpzVlE7914cJtd4GNt
461AaU/08QLGlSOhM9fJE+SClSxJdQgTPVJbKWmWsHcbEBlFU68VvABCQZ3NLIhw
E2+FeDeaNvPY2J06TpCF6FuTv/z/dufS/96sQwdSyVREmswI3kBCXqyOjFSPHh0F
UBTReojUSoGvRM6dXaK1sDw2WjbFIs/kQ4+/13D/Rtz4V/TH02R71KCfQcgS1s3P
8+zL+3+6g+SfaddHiRlb6JvFD3679rkz2qzl4rylTcF/+F41wklr547QMQMOpKf0
XdmAkeSQpqPqMzSxN6H0d7SJao9wAYebDSw4OaRFWwRFV5q/MVz1XZz1uziJkaKc
ldXy7leBuV9u/Hz5TL2vGacl0BXxj6vkgSBCRwPueztIcv9ACHl9Liwi3NSkqiyY
1Jm9KaqKxpB5xe9g5nFhHBN+RDTFyPocMHGFNa0SU+ftDn+yZmJ9RtsKJ338inwB
aPi2Ls3NGg4K08IuAEZVqBnt7WTKwIzk+hz2P+qpYsGc8NWs942h+jn7EKF2UYey
PDcsPlwfiqS8Wq8Anynj4kbXG0K2tXC/eUnEW6OxZkxZDH8bucMfgYQWRL0gQmVV
huf+DQw2SZnNWI6V0XHxcRLMHaZ/S+WCYBchG0V3aiH9qeENWneuzmVjxSiwrRyB
eLKlW5fwedY8BxH43MymRke9C7MBfGmq16CsOyd+Jp/1fjfu3f5f4VnqGcR/yzEw
2WGZseZ/z8RdfTq6fIlbNgwlokyFAeSJQnt7ZI+bCcLQgC42ycmbah2oNfDVRiLc
NBJwNOkznpaDdImRdg8z3qL03zqeZj/IEhpMszfnb42YpE78sOn7WH0MZF/2to4s
EkbFRZ+0ttGi/D7LKS8XhCnWT+t3mCzw6ehHC7U0FSjjukVrmVTAtD8gyZrRRNBk
UrgshdP5Xd2zRcgAoClyaNkhOST3osodVBMzArXLfikZHBllM9nwiJ/pMiFHTBAv
NTjX0XqMR+dW7DJEm7BENkBrESkhPvDusnGb6MSw7HQPV+gj9TxEz1n88iL57Jju
pJZv6DfEptbHD1cHnipjph7oVjYnRvzBLM+IpMg0DJprynnD09Sx9+KZqMQXHnaW
9g7eeGB5bgnNhbaAe4H8EebJxHu209DyDfrJKatiEkd/yhSmw5ceWx5Y1PUe0+bq
GW44rH4wmoRVtF8aRXHYJiCErTHh9rAFVReMmp1uTRUBc467mnbPgLfkC8bVyBeY
WwEHvDRpaV9tMYpX3z7Mq3fn5tlTf1Dl4N8W2BSdH9lKbZmjs4Bd2okXaCTee6R7
9FrWs0rcIgy9QnMOCi03BRooq6dqHL8Nkmb6LwEQh+uh/+P6rFYcxMx3fh3eqbN1
pTEIKmHpMt+pSXeRC+yrchQaINX1Jceu+Q7aTcvBRtRDNgPVbWRHaDYlat47Q+Rc
eqZV/6MIGxdg8h2J+6I6Y4gzrxlGdmNkaCMXzzxe9K4hQQ3AB+N7FcE/YpOkR/Tz
VKOO1avq4T4dFKVoT2v2tDo/Uqp9H8zpGHxroW+jDS1MOlufBTizDm8LS2+H2f0p
lNqlf2RMxG7PMpokoulErxyTQ89OyQvxNVPy7SUcYf6hSaosHG8kPls9IAGakDEZ
4s9L91TMh7MV91LK0QDgJEKFos++zAPqKDaaFkXBapM5Ox63icEqSF+xk8CRfjLa
nWXY52XejvhytBvEwO/n8xgHlAa+sWG5dpmc7yfuz2KAld1AZZWQTDeAHA5g9pTi
B0aqSvLYA/vQrF3XnxD5KLydEuR7CzZMfjsIadipmtSR15/Y9xuPEUGsHD15ep1A
Vss6fxj6xlesqjgc7tq9cHSoyJsSR+YZuLlfdZp6wyEDWi8Z65rvLAe8+IwgODm9
4vrbrYh090N3JK0LZAkBIWU9wOv+B/gDd7aq3McR4fJWsG7x1/HglTlrc6qXBF0W
M1zVKoBAC5O1KNSxK0sBK6cbUTJYA3K3orlqLUqVOd0wTezBOUpDSE2ePDS1mbYQ
DEXigdKom3snp2tdke72TFvV8XQKEjjB+z7fz02sVd0Z7KuxbORklPoNwQ7AS4FM
Hnuo1FzVtWovMwYrMBGW0SrYS/f863yGuNAx4CEkrNBUaymq4CI3K8LXJLATqSFj
KzEXbKbbrETWVQWd6dOxqdwbrwKhBh+fI5uqjxwj/QKKNhThNafyvmHDNFX1sdak
R29jWr0ZWuxBBfwKvDj0DqXFiHgp9XQcqgDEAJJg5bJrHfKZXbmYkUp7p1KyfYCG
hVwrvyyHfvFc2ECavehPWNPJhmOh6CpElT+F3o5lxLRf/tbIIlbcEgSxtIE12DL0
A3lcrmFm/Z9U9HwibTMaDWPSMGmcgubnvrTNFiKBC1ENHGD0OYrnlrnPg3PCawn+
TnNKauWK7Jkm2LqvPbknTgk6QaYSFhczJ0sDKlw4Nk1bRPtBRQBhjNaaZhVt3DHE
IRoBVHzngsPXQIxg3NVu2xGlJllx1/vSoNxaNgud2YoLtC/+A1iHtfAAIm16icHm
mHVpMsGCciw/4cppbReJ/799H2omBytlrzEUMbK0UkjB02LbudjwAlvFI+o4Th1m
j+UfF4sjpcpzla58AXVd5q7zq6gWtYNgMfaA5nUlLsAL9Nqxujx1NLG8X+zfcueB
kr8eald7TJHJyHAAhNL2CMZuVrQFb1jsXDawPWMfh4D6iDdwqwqjvM6fcJxbUhS3
VimprXdNsaWN3IA/M+GMtd6rZnK63TflaNuUHw98PdfbsYPaqFfRp6+GNk3nBm4u
gsn4ff53w9TWz5ni32Yil4b2Y0fq22GMRdYInCyB/wBFFs9sSZTD8LM2y6Y5n8bQ
ooJAdGaeJGo6d0Va1HGVEDbtHP7og+gYU43P0/fXQTli64djGASE07DXXfDsiSrx
XhInvN1/F5y1Vgi9dIjn+NjaxYa+OlQrThDXSU5tQaJ0hqSrR+wxjZn8TVB6F47W
LXs9OxGrYO4tuoNlTAH+3Wb9W561ZRhmXJYJXryWSt5lJdqBpQ6WyuP3xcrREX7M
2rYdmwYr44dY663gg13KrbU32q1IOTJtbBrF0y4s2RWDbnm31ZHsFtm5nBgpSDuN
GQHPRzb9yK+u8GtG8SIilNv/y1SMy0NcSS9KAcySHB9j882189zt+CfH4TMxcaOH
3rynoTDcFoOsMKjBBQ5VzZsy3JJ+GKTjq0cvrv40vjYN/b5TGFzhG4ueJkqtq73H
iLDYVYBG4FOwouAh9PPS1regwYsVdS4Q7LUVwrmpLKEjnHIcduhfRDDAJIwjBy/a
LPsnFGjqt36o9NQpsKtviv3BR0MXswYAvD/uR7Ju2T2kgXMY9BuP7cPSsWiPEs0F
8enr+sB6r1PvtCVoMUR4WS6dmU4iMVFY40XvmAfQPUnpsVxnbEiNNz7ab+zAd3HK
pH7wtyQIflK2hv02A6fNvzGfbgZXcnspv3SK2ASIP4XVmir3ZqihQS8rUNundbBC
bBqHJXIfBu+mMXZHWHQatwnIqX0k6CAhrG+DLlj4AbdjhGzj5+sdCA08IZdcyA2z
NLcZCsIrw7ApMkceEM1V4YWvy9fj+tMkUz0d+NILAlD/6ZLT1iYz4BDAOJ/KDxe4
Zr12qsf+LQeoZgGlpCqr58nByLCPjDyXz/2FAyH+KigsmF6HkfCT/pQyR1jhyQga
Z4Eiv3RerfuCi7lL32IbXZl91B80yOHO5T1wb3/S7u3gOnNmrI4slQXDtx5JDBy1
JHoqyjO8Fm6EnthRkzWDBBXPeCO5Em8Kjqp2GgJdarTUEUVNSdnC6ORHpSAEjdau
/ECZiSo2Mz59NaY0w4zP1YExfj0slPPGPXSlZZ49v5WzqBimwMGyME6rm/XJFLtC
zjUrBj2I9vyd9ZkDDxoV9c1nBSPesRcvStDlS57QbRgKaxplrw5CbBkcckOuLgrt
grU0f616IaE6wv+iopajEX3fJqhrDGxBH5vLPx4+Oz8XhfhUq5vrsH/J0y4rBfNo
Uar1TSZeo7yF3YxORQodEYXTnVH2OWyWDAMl5393uLPEMc0WEj/2Glowes9Zd1gC
cgAiqj+ElRUH+h74+iY7DoZKVmfenC9AkyMLRhkIQdpB8oPTCyX0ahczNjf3n/Wu
51VcCd1W9QsKQpgx6SMbBkfWYX5AXzh1y9xuFRQhGwWj82SYsDE2IuxZkBvXst5R
Iuh0JaBNSUr07ZlRMx6NlV/Qc08a5uT2F/+S9w5zJyth5mCZD24EMGOQUj2mc7sm
zVxK6i+y0WSeRnuTagSr/aV1mzgu1+r8r4SWYPS7ng5RqrgP4LyGXXUbSWWgxpxi
VxKDcyIL8vG8F07/U7G0XN5Om/FP5jOzEDJ6TUtRuOTstJpgP4RhjwSNlB/bAPGm
`protect END_PROTECTED
