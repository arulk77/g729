`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAo5S64hNPmRq7e3k3KET+2nhNFqWMN/mEV3oLXgEQqo
u3SX4uplNGWrDlxp7RUqLzt/tZfbn4w/uigBkRMcCUULzKUcr7K5ajTIdWGUDuif
8k+nqVB6V2ctGs1iKDsBTiAIrOGfgPRmI7XpgFeGzKwS5G8mHd0+yETAK9Z11vZy
X+wKy64s+/C0S7Odj+ViwWtyfxasn7PonO69dXiF6ACvU4ZfD7IotW5k/L2t2c1o
`protect END_PROTECTED
