`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
72DKe5MEZSH9IT4s+0rFcClbQG17GYTilvdo+wR+JYJFoPAy42c2KsceHkKELbs0
9Ykv27RcqthntPme7AF0TkfzcZGYX+MTI+rGJEp0ZYZDECbd8k5Lp2Q2Mtpi2/Jw
vfa0h3Vd12HxrSgjioVMXMaxcGfn3raePXYRRNGvs2uVyWh+ENfd+DtFziibmzAr
drFjEIyL7ojTuKxdiL6ly7Sm0Ks/GSKgPOnB9iCyXZRR9AJVNXzZ2zXVJroAL3FA
xvuVr206aeX2bqcwcGgytsSe8eTVbIOdaxc6dcwDT3zy0AIqc44Ewv7I2N72rogp
Y5yI0osIupnxr02Tbqk3dkLaWTaWwYzPK3mNMh0nRNQax5oyObb7BuBgMzYWmJJ4
`protect END_PROTECTED
