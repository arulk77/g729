`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aRXj8Gic8LMnPzzEkr02UB+H3iMIsjydANZIVaIEbOws
2jlh/AImLqX/OjA4JOUe/Rjg2HNdyB52wXcRbUk8TvTBRYXizQYufiD6pjm7Sxd8
mH1t0M+1yrnsKQBLetPYVFeigHoFrn0z37+B5t8/6xxiCu08sSBEIXG/ZBro95u7
iFGQ7+JIQM7F0JuWZpvRYoyIcKbsNRBpJWMA4YFxOyPbBmpGOSO3rE+ZSLP3EtbF
44rAIgVWCDSERVFVlj88/35radrLsU3cEPmZrs6nCHCMYbSfUbGyQ4L0mbB2hyJB
WKG0CJV3LGHLqUAU/YDr/7rsTaE4P+vg2i/OH5j1c+IcuV+XKGSEBfnwh8LHPVA6
G0hF/lC1M0AjvbNwwAWxoIrQ8dxAhPWvmz4Ul/kHRDEoIBTGjT7Y1Zt2shpmhLF3
vtfqz1baoZ1/gkcRfRW9tSJZuZ/6526EDC8jXrI4IgKZhbUsSlvxjM+O4kavm3yx
3BCDTvijIRukBE2hldSqPp3vCc39GX4a3qfa3UDmyTROkHlMNwBGpTuDi6COxEWA
b7bxgca4gYX4i+z9Lfi29V+uaBIV3gWWe2sKr1yCFK5YkqxAp4BN9nDuFl0dq/8/
TEugbev9LsF1eqvhb2Jz5KQaJuiF/J+nzH5Gp9frLrVUckE0wA6wabNMG6lXonkZ
nUBLftszn7ZMYaocxTYXbECGJgYyOIqCQ1vjC5dQiC8uTgZ5qFi0OuMA9IH5cUpq
WvrARCKAOxqKpkm5ayvzZn+qKoyS1XHV5qfdlE3JZifWL+nquVGNBPcjOFomeNvL
sIBty53e6pe+l5QGkvmj1regeHFC3lOYmHzR5Y/CtlQ8osPvAcZod+cyYGV9w9zc
/N7lr5gzriu6HB8PCx/omlmbQxKAiKZZzuX7178r5VtSfPqRMwdxtvqL3f4TXUVJ
04+IyiajU+ZkS5hhqbww1XqxGOOWG1iINV1L9xkx8Fg4NijnTh2FK+Evof8JzeB1
cdYoEMYu9S3Ve+gjIU9AbRum1QL3FGNlwtUByUExmphhZSuA9fYus+zv1LeNeJ97
Qulj/CyjkYTkSyMrCsuO0rgO9Ud39zqlAN5AyHna6YgB7pSIeJwoDJb00HPNyKTf
JodoDyd2GoylGL7LATloGOC8xHJiai5Q5096lnUoC9k8918uDkSPHQY0Zr2fputA
vzjUP9ZzxEYoWiojxrLpBq+z+fXqvJUwynne15rXHT4KFsU4P762H1dEpiiaku9y
onbViw03rcmvxTgqM//nTCIq4C+xGLvYfgn4stNH5xDdy0YHjeaLoORhOA95Bx6b
ww/fN2KTVV96VoLTRAZ0B5f+v6CCIuMB7vABAQ5A0W9EbiAOU+kz0uG0sY54B27d
buwBOiIB23tSsf57++5kSNGaV5clzJxpKmOUm4qzQzMkwRsA8wjWpoTmcrRiopNZ
v5NHWVfavXEh2bpO0KuQCR91fL//VgOTLnXOX6aAyACkZwheTETVFHJnfZwRFPxc
/CUdilkjriZxF5TUhiSQJAyTAlGoiY35gXjzhufbld546j5dC7xZU1wmTp/UuC3f
ADrqy1JKCoE4b9jVfq6tLwtcuwBxJF3q7JDQ2wk2dhROOf+/WqJp1tA3CiEX2hdb
ijw98OF/9Zha7ndg/BAH9PTob+PTEOUxob0874wLWlmwy+5CbaahHNbPk/I8rORH
Pvy1yKeLA0m5vZwC9SlpirGqURb7JIrNkim6O4i235Fn2/tfUYf/0S3jU2D+XDXJ
Fmgs+bWQtdRSWHmr1XsRg9sLEmN/hxqJzwkF/4McTRRVW3TYKBwinTyzhphkrbN8
lqHduqK+j/acA1Zr3ie11NDArrRlFudpzvFZpN92v8U3qwSXrLiLM35YHYcf3Lm7
79yffaOd6e+Xs2XLuYMWeJbTqdOyF9epKFnPsUStpAIyLehIAYSkT0baCINpVxHO
a0EGcO3TGIqyTXLOziqgjAnENZ5QVJ93I9+NxO34Mm2/WkZHF+YQE4p8PHnJs8mp
Yhev6oSpOvqD8CJq6a0VJzw579WRSqPHqigICvS29Xy9ciOqUTRNzdI6I4C8l4Ou
kpQ1atzLLiUQ9Acmz1mLVF4ow+vT/MvaLBurT1Mki7P9bdEPbBqpMdSmpRLEkKq+
nMWz0WriJ/eYpzfjmwWoIogsH3Bb5NYNrRFAeEFrnca7tpNhcU3AQaoEy20NhE/o
WzVRIPAK7Tvu4OoaV9VUbGUL1Pp6Y7x+PC2z5KIgzv3xqydtppnR3nCbFDtUKqdN
gJYUV6TAKgEkP7kAE4kflTz1A426HKIN//yVIHNfofaYcGc87NPXdW+OgUvTxE8H
OkQMuUSrgQ3v2k6js9tHM1yHHhUFHSDaCcmxKd1u2vNs4TvgLL4dbNLoNjkRqg+k
5dhP78143POp5W0OVVVsRdM4/gBjN34J01y5cYxA7TUt8Z+Y6WiGTS4ctDTUsmwy
GJz4pVFa4Y7uIQN6C9Vvr042H4v7/HtDwGyN98fsyKeDuQ0sphszoViaHNjBvbO+
s9lO9b0J6FFOTxFOr/1deee9soHoB1tUfhaVBFwfpoLWPNa6JZ7b8/tIYIIZ7/i4
vESgLQAgCHY8Bq7BbhUoWOX1kP0CIMVxK5dSb+w+zQiHXTeK23P8SmptjAMzSPZZ
HQMzajKCyid00HUIUDg7Ruofue0NbjDzTxYqnJY4PCL+QucnZPKt7aj4PaP2Tg+W
oBBGupHekljYFSzfohG+k72yEz8KTogNIol6QUMTuJf/ccg8+m3cycfTdPzcZ1ya
p17sMe2uR/YZxqhNy84GMBZTv0HIZM/El0koMYncHT69gt/S6Rkg3RFvR4dSSrFr
PKIh6OFbAYhP45UzsmaZ30GAwirAPgl2Fl8sHB8xCDc/rnxaApTf4wKtt5F8d4Za
Z7nNz3lBspWv3VQnih6hUtYHEXfI0AgXXlFbdPSWAi3CRDUDZtYCd7lVADNyf0P+
IU4xZRMXmoXOJSqLD9Nn86kp5N+0Tk0aOKoxZCpmVWw=
`protect END_PROTECTED
