`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMuSl1RAJVyv+3lO1Kj+SssjKoyNISZRlEsFHncf+gAQ
eDQRKQ9IPXtYnpA85rNVGU3d4vd8xidcGJcWdvPBTFkqIZJcwtEJzEFAgBtEsKQD
ZvRZu8CHwI2NzXdB/II+R7m6N5WzTxtqNVT0uIHt5YGsqTnsweLveLzX2eT7NHwb
CkaQE3miLhaUKKoK6obodBO9pyV1YbY24M+qmnMpfDT5Tgn9v1Gi0cfTQh1KhFaw
CBr68wfD7iDpL48Ghw+mt15sLmNfRKjq2qgbwzpJIuFlYnk0xjY6RgNHxvdMhtZy
y+oQ3yc3WLB3QhViONpNHiJobTwASnSpkPprZw2S3XGUW1vDt+IDEtKaHoINnCoc
kO6SvQgT7PzoSKd4Ckv5hqzk93xcrCRBkUdfCDt4HXcwS76jm5U0KOVmJrEhykhw
lbWvG8iWEG4NYXFUP5LHqAhP/PVvowEJce2YBzpG3BNfKOw/3BqufTZGF7lFCTNM
sNDTXxPiH39Q4lQrgm/bcFjy/fbvjcVTKMxqxUAmj+C1qkyTAR73PK5ovbtmYNlI
41f7rTE/DRNqQloq4NrlrmcB7LdQ0x7tRghm7rT4axLx7dF9E3ryvv0edZPwgSpy
VZPjY4HQ3bvCI3Iir3ahUC1C2Dy0BJpGkP9+7ArEYVSuhPA0yEBfq1/K2rD2yAq1
/lkCd+9a8YyzLOgH8N3mUe+BnbOkEt0wdvWWiBrYooJovEYqTpvStpxyWIIuwsW4
HQ4oRKyHj7ph2rPB7lDk5zmg3Ly+SEOQ0IAzyAgqSwcOvutJOZHfLjbA05KnkkDh
z5WVGv7sSY1xzrg2HPpS0ECUgdKUcLiGLKvn6b3cK4M=
`protect END_PROTECTED
