`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOrerDh4pPDiI35dGuPePXy63LOKi5BrTylmcNceetsL
YChgfT0FxwGL+cxZO9Dun9XrmHwAEmgutaE2Zz0ED0g0/NL3CvR1nKNctoAkIi+M
8D+yGl6LpBvLBcI9coQmwCBtWeYwufAvJJlL/dVdyuSZnXZK1KNh8Y9S9iwxXLxT
wM1IOWMzJbNYdXQuvkA1Wn4qV8d5/71jS2DqHldPdEximsM7tgqzk9l/B3iHnDO/
+bQ9BkN1ZljrM8FTEsciq5hDTXfLhYl9XhkknTip82jRXGbycBq0p3+yUIF1Fa2R
2UHSG8dGcrLbgMMjfZJ+lZmrnV1FVDIsrgTB1t9xjIzPVG8R7t9Z5v5UN8S9Jvlt
lOy2pVWCaE50ipSgHLqJuCHW230vvODQNPAdgBd8whodLTh/IkVYx1vtcyHNZWHG
DJpOLT/BUDeY9Q54Tl9kGRc35tUjLoabbLcb21Ga+0+48fOJV9XAQF0PXC9J3N8v
u9IfzGahiLMAMvKeXkNI7A==
`protect END_PROTECTED
