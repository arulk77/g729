`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
DO1J3NoB6qL/VwpjQ3Ddi14sKkbN9aifPkF+zXH1CqvplNmkyjc0X+L9X9pIFWea
dPKXuKzmbytdeRhQz2LbMujugZ3xUxHFpfKLWUTjruxIYBhfdGvNlEsO8YeyFbi/
nIgQSGgZQwaMPVUxaK2Wl9mnXezIjuyrIYccjDEA6RPNQjKoGIucNHSuM0Hocl+o
GcCeUNZTl8tUwTm4OeJZvBquVqJznKaD2QRp7g594IkvxglfcPQ0DkKgi4JmF7ck
zp8EKrdXcTdQy1wVOGOPFJvMj6Q81qSQwLDZnPTdrxk=
`protect END_PROTECTED
