`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bjVKth1cZgycmK57Rp56+XFzQzkGAjYbyF7zMKhdkLjVyVAzuB7WyTOvgoNdV3F5
yh07R5Y69G34ZAO38licuKfxlzK3IE6Scb+MzpgpgSBrX2nzH8L4hnR5ZNQfHsfd
rhyg21DqJcijZVXNGWKR8rm7XxCpZUuVXLhWkYehZYH3E7FBUu/U87SihJ4Q73qf
`protect END_PROTECTED
