`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3cIP9E1nepUubGBK9azHi/V3DMWvg6wj8753Cr5FGVxKHVLIXIh7gxHPY8NTbdp5
QKd/vYSm6oVDhjCp3UIiMo2WsX/ufI2zwpNWspG62mGfM3/d0/y1oKB4D/ErCErz
hzTOqBPx+cousD9AMOfC+LGaoM5KuP/tCLHyB7cRDO+eRtnEdcDN8LaecVAPpijE
95GHqX2DCRhjrBbKkBjiMBWxPqNAXP7zL8unVf2Pm3R/KxeVfRDu1uAaGKG+Ta91
rrGr3PziwPr01v4v3onMlLM2rXssOuBheekTE29yJIOBjvGZUHDKP4fcAwAu+zAf
sSDxgp8x2s+00CIyRNxiR+tPy4/8S34jqQ8njSvyHH/bhwJn/IMY145bPeGfeOiq
MY9OMog1MY21Mh20DA8OI2lL6SX1qAJJU/YQw8MfceqNd8gyp7/6Xxk4NVQDaZrh
hQOrp938yn+uKcvCUZ3WSUmaFyyjJlLkHZsPzTOAK3OMgaG9pe68A7wfTTCk88Ju
F+TZ1YsLDEwwb9+VuT5FYxBw9fs7WZbFV+vG7JSJgNonyB8g62sGwY6qmqdr3VTD
zbLclN/Rau9nLgcZkYtLl3exknw2DesGSvIiT3lPuyrlIpWICGl3JzlajXNjIs6m
xXf/2xFKIap1Xn5NRFYjeAkeVx1Pvt+kbXyxsSFfTSYQmnvzQzu0HpjcrY5zR4ZM
CDSjfQwEMTPotX61JIpKIp7Q0J+NN+VIBOujewdzDqgC04d17tUZPyKT9HReL5VP
gxdYsNBi73MiQ1o2iKP/lqqELsHQalRBrWy58rB0/I71GugXiTdkHejzkRLFno2s
+uyCrtEsMxFprndgeP/apRPlO36sXBVUniH5DUOkm/EI22AuHG7Dn9uEe5t2Hcg2
e5oFG2p/SUepMOK5ImcLaut4odou91f6/xu4cq+UhIAncViQXLD++r5S6bAvHBvS
GPVomYTbSzJUGosgeCA34IvOUerM08fy37qSrLJjYY3ofIIdXrfz1ej4h/5WVXPS
oDM+WFV+bQw90Sr03E73p9ZKOchfcIC8tiwBQxwZjX07gcwPyxwiyIfIMrlFkEFb
0Z0QwILbwSI+66bltJGE/FWcpPkwZbh/qiu2WTwyUW3Mjb44MADpFytMz4gndbMD
Ssvx/cUqCJRZTzmkUk3RFMhse2qHmFSVah2uUPRypa/2kNpbvKmkqO0bZ7GgBgBv
puPkQxSaRuBYDQobC48SY5EVZlGRbtyDyI8QUsS6kGTDqh8TV2iPvQCNHI9XM70e
ZxCC9J6Zs4666Qa2u8Qr7v3i1wXq652y+tQOLak6d59UNZrgdsK8DuJpCkqrcDn1
uB/1Kq88tlvjxs9bBGbBn9LuD9dlsIEHVH+PGXDUm3kRkjIOwWChokf8CN6E7Z86
e+IM9G2ZooTXnhOniyaEDEXcpcejAaV3DNwHg0fzXsw2UpYjXVAtV78s3Oy+ORY3
gFZ4PW1RumnQj8ADxGmuXI+KTVIHd4CgnpGf5iDIKrm+Am8E1KVQ1jLHggfTFDFN
xBPc9sO/FD3X0mDgB4stNxHWBWE7OgpSjIWQ1M5D5pWZEMmhmejy31FGu53ILGZV
5N/gThie+gE6UJo/WXZ5909ebpHT5+U4dushMPx/aBRkA1KAYD3z2hynVKBCksFs
8g5tSAnEQmFPzAHFZWXTZpYstCQshb3w3KGsPDHpM/Us1026LBMDs7qHtHdIO2L7
fNonOy3bwlLInTv5hr17WLMb64pZwZ15RaoSk1UGTu29rzNVkhqntf2uwL1U7OjL
TbCjL7zpZgLFxs/PW54BH5LG1yy2UnGTeB2NAo66S2lH1EvYLlBQl+Pnwz4DXScd
jTequPNJlSnwZZ3Ilzf8ghYdD/dc7Jsgfyy3EQ8eP1Aqh3iB8/MVsLvy14Uzyglu
gkJeMJI021V6du6d62zzYw/smv4iAZhmUDP7ZeKbdaSA6mkCHq1jvmhAxzvunFft
P19vuD3e7FKG5SnzwIooPSuWZF8kAAb/F86KUgJ2gpnWn4avDy5Lvk7kHk9Sg/Lg
cRvLMpnRWcUuKgtI96YkWXgN0+NewImA+c92Ov/7+1ApYVwvZCUmSYST7Rc20ixj
WVuHhDa6yBCb1BzgwtUuONtowAseujoaJji69hT/aTn+H4/Ga4MU6OPPi6iO/976
AEFhb5TBcT+i/vtVnT5LKKTL8rVjDIprvHG/S6Ng8arecUSQ2ocaKjE+OClar9Oq
N30JWXWPpnkDF3SY/x+rxKJVxVZfXXTVuuWcXQ03pXud7XM459i1imTrN1re6G9y
7JpElI6/CU4wXCpNiyfSCKoHEh4Nmr0KEPinwy0aDgJ/EFFD+KzxTJL63KrnhtOr
nriiCEQNEGPqICV52knjfQY8yAKe6pF6mdDckQSwlr0Qq2ynWZH4amR1ZS/Yk54m
IHmHPcWYG5hSyS39Zk4XeD6/0WNXM7w+rD7aeZZrQsG9SySw7Q2zn6cHhSeZPF9u
DRaNasRTBAgmj42WfZflFvd72jWmNrdRxCmGjL+2/zBZ4TNUfEdmOL9uU6NfmE6w
JesuSedmIP05Kwg4jkJjC61Csb3FQC5/zPTHIC2TtFXx0aekjrZU0Y2R9UUkDuR9
tDIAOaeVdYzclZ3xD3taYIjiJm3LCnbC2DYuCCZHw+4OZgtUHtxdeGT2ItBxub36
L+paUGjINYPd2Qmz7Ibi00BTwHbPsoYUtGAP5qxgAiOZWUKGjoUU+tQRd/HMaLtW
Oaeh9KVgq1TUDeeQRhwJV+gJLfUwSKQP/cSc+loh88uX1pZ6f+ldbkB0P5B4uy/+
eRwNBT3iFNNKE0QBzmDuzF4yqU10ipxmKJ0+g3wYLW5b1jUUqOAkUfgFzWLFGuWO
BkAA0+xqOG1tp8rki/lTV7HVYv0nUWmfrWPhQWxcFgZed1QFHLN5ca8R0Jb4eleR
TxrjdnqeYwyol4mm1DpzRv9GBwnubwyNSQx10a4V4dEI8dnaRwC4GOqI/enxGfVP
n0CN74/dtQhD0zyxbz/yV3Uv3YCWazqCRvbtKqWUIhaKxRm1MhN6x1vvm1aJy2dV
fukeB1PZQLjVMIjHBwoxi3Bbz3ShWFcSdTYpRla8UBB6FvRnaJTv5KCop7vaVCPE
GyjCk5mlrPUE+Pe9J5AbB1D2vDC1vgRuzMufm5/uZWWED2He1Q90g0nq31jVFZYA
VUqM3GXEeHWkgWK6wPXZtG/8uAB5pBn3n1uaL65PwJVtYAsmay2qbY4kjXoa1hbl
j0fNOUiJ3ObEQLblFsmiXLv2DkY4Yw3JKAd5+sMg6lLyGmnf2li2ES555M0Hm2Hx
OBOke2aqfEkoQwevr4eXWSYADcDnyfqkmjSmFLYVzIbDChVR8KXhLLnYVLbs6dHL
NqjcF8pqgA7ituEZWW16svP4qQliGH6YTNJ2jc1CVy+/M1UbCdRskmrGakk4Gxca
vlMF9Ug4VvlsKXN2/mjQsTamGNbGlSlkP9lemvn7FRe853eOpu20wp+8cpOHEIAc
zQsSoZpPkM2w+3FeNREUl5rd13YjZHk1E1tmdZQTT3kTViFWHfUtuPGVyIe9doL7
/MeygGV8ynwPJpu98p37DDHVD/ivJad4ZsbNcro4KY0lltMP6VPUcbGcuiDO2dsS
BKnaSV2UBaW6QgB2JJByKzb/emDnI25LcFsAxtZJRAee6SG4JsAQE++pHggDzKjA
NPnyKYNnEOOyRavpGdMm9DUG2RiqiCUjg/XDLw4oZTZ7CfRIA411asYluDmnd5wD
69InvvNaPqSNZ9V+XQuDzpgvWfxj8OnzngABzHkSuSZO7XSVciEiBV//BKkNASIJ
wf/oNqkiJwal0Gl73EmaEV8r1sQJkV5F2i2fJsuofKDDQuJXJKw7v8ChY9yCscIp
Pa8yVFeAPyGEwHdwQPFZJXREeatIQmx5J6HIeHzerAaMjHF7U7WJQf7JJp031jFo
e3eznl/BpsLfelR2tDQZ83nGICzjTP3xbiF11iDDEbM1byxD7Hul9n8R81akJwtd
9YSdVAWyCJi/IN52S9z/8ihOsoezYGSkwJxRd5ltG01Uh42W6jhA19JHi/1WstMM
nj2MwR0qG0AxL+CoUQ2jyfneBRCuHZrZS11muF7UMAThSpRag47ESQTUlig/Djsj
SP9Ap++s9t9CVCr2i2dTxOAQkoNVvxH9GKEhehdFSjM7Rmd/Aax6eX7eZYnjgQOy
Os+U+0cvIacSQKPKrAfbqpbS8KjLFGEonXxyWSFyUvQnotZMcVJei/1uNzOnibCH
OfZEz16vISlztA3BHu5IZRhsIDjwnnzpM+ZN1Z1RI/uzt+2Cxb0BCfKWy+XY8Dwk
b8VRxY4K3lJKFmvsmK9TY1ZuxEp/xt6R3S+CBF1qdo5GPTWDHsxeiDRjiwC403Dm
ZGTUzpqiYI6TSCXq3JaT2HH/XPPX/KL33NbocXaaEWKSCjCwXIQIwQBSuMDKqBud
jAAKaAHlGE7w4yaigfLB/Ja8QBZW5vXGQbkYXMLaqS1gIvLOkn7zHV/Vw46cVak7
sPSpO8L2bmT/xT07gyecd4cRTet5JU5SwZLnpaPiuduaY7LzQXXB82q+WVc9ZIdY
ojlQfX9yqyoxBk4funmFFsSKwEZcVxNMxDjj7jxHIfzKFSYa3VMNjZFVBiOOuse7
NIzgLinjScEP81qSkhbwv0meTgPTy42AoeNtg1FIzfJjhChswYgNQ+4rOPsKiVxm
1nGTj4fO2amtJWwxjwj8RU0SVUMsYL7UlXa5XMkKgjvcXkLbwp0YuvFRLjPSoENc
Z1nGZarnxm5v+BY2a+gkgO2TMwnWOvKpWA+AIXJgc9bsMUo8/iibo2k/SucfYGWX
zHRqwZC6HgOv03urU8BYG5wJzqDnJx+tklOPQo2SY5yiFY4KiqryNbESuzlwMQLH
9SuEaMplhVn+bkAMk6afoG0tZjtssIDU2B1jIStvjl7P4HXwaAjr6xWmxyU7BEPP
f1EHFAxgh2TNDkMXcvhgJlwXJL8cjw2SjrwAVYYEpbLjHA+W8Vz6ydooMkzDBxTT
iu9saKjg+WFTHdiRAno8KtpsKDnV0QcfrEos4zxRbb7hrRZOLhKoLaQV+cyDMdH9
+2Gf8ztLkuun3Ana7VlWH9wZsojMmBUpnfjLfb3jDGn83wWyPJmZneqGXkL6PzPY
yk5ySLQNcujaOCBrrzW3HIXAseBNckD9P3x27VSy7hUGm5DEPwFYBIMJZ+34dsl6
OfULoUcxcOR8eKmAT2UAcmchiByHFvPH2oQfgq037qFPZL2vO/cEfl3yO8CYoL11
J+eCeUr9Sg5JKD6mZNumFq3jQI7wMOqSbXEX1/EvwYZi2gZlU/PlB76/V39DgM/Z
BMhi7Op6fUxEY8QyTHlOD20OmqplBQQzw+Zg7I116njOyYRewrjBYDkGdc3rKivE
bqa6Eyggm1Aza9C3YKmKRiJRkWLs0+yNy967aihcXZ/kT7kpwsEdND9N6B2Wkz/0
IQJyTlyFEPKjjwtLV9flHAbeYa9OXud/+BaDNK7fRHyWTkOAYwRzNXJNAK/5Q8P1
AwQZ6c0fhQmYLGR2xEzEgW4niA8Or+Tdy0UEHlbIXRnzWjeHoQeDs1E3vgHGR6Kx
4ah5NFkhTHh5Q8x1sWMEJ2M9BJxURNfqHFQFXnz2NhrvVbcV2bX/+0cEGCSVIsSi
8Use2k3K80V8WAe00avwgezDcI2wMYm+1d9fUN6+6q3KGG/Qp1MtTssQrTf0SoaD
3Kyf+hGKevRNhkYh+AXAPSkg3tKzZK57vS+LmHjFKjOk6S3xhGYbh5Z4CItn+HCG
oPajA86CiQ3Q5ycZlSVf1whoe37xqj3a1QDtL4mqbboqczUSEm2wsDfgsKi2izqm
175A2wRLd4xkPUlvhaT5PgApplbvWACVpI938hAR1Mnc8yXZAObFwRJG2dw7fA+0
1Sw/JtVuGQOdF4T1zuesp2eviVOcb6d4Dlw/65BEc0Fxac8TlUoVbaJW2csB+p0H
pJaOypHDtMoKnAeAYHGfDhL8KIawezabeOa7IoUzCKP4MOqmKbiJBXtl4dyPIw7a
NcbDJqKt78Npon8acSIW4Qfg4OkAfU2Wp2wZ45cwfSPUzUR2lZr2OxDzluuXdfTP
ApcsNc/ZvJosUhM6PixdQJPSwvCJaDBW9tO3OugfUO1gsARSi4gkCVNlvzDr87l8
X7gAchGG1lAVnJAX2MJZpFApChAGv3NtVqOjfT4VHQ0tqlgeLKa59doZ3JXXT+5M
Mb3m2guxD6LjXbKLdA3A4h9RCqCjOc62VOKEBMuvSp6orK2gr29FEK4faymEgpz2
BQ8EftULafqpPtcEjC5C85GmhYT0jgacuO0mgmFLpJOp7zwBKfG3R6KW4+s3hY9t
MGUIdBX5DPiV1QeRQLCwvDXzqDaWaoAYrd/IGGB0nnu5kI0SPJChd8qpQTdERaQv
SzOIDqzmitXlDvYnZdXH1pbNi//UV2HlpaGB8BAgri0SXsvvTzXR4yOG6u+1OLm8
jkycSmk7O7dYEdLvOQUEhmsRl8sgqtXimLJRz5JcUbrMrfpVYd+4OMsiUZc2oJhD
pHqzoPYPJM7rBTR2zK0yq6N7ItbIm5S2voZUZtL51lStA62+AqvFBaPgB1Qe9mHJ
eeVaXIZo8HYaLRS3sh4sFTS3zIXkhOx12sX4gqVCslEDsiPVMUSAbyTM4lruW5Ao
VQUvSNHWR9rrEYGIfiSpDOQ/8vKGHusQOKlUCaMJ59ai5T+qDIPdW4IWPf+LAz43
0TbI9p+4QaBWFc0PYCGI2bAYEZmHYfF2A0FOhfKxNv5+313pFnEjnxBMI33uozGz
7qPpMLUHTy/cmGRVQvXuU+zHtxMx/4VtJxqVB+hxlcchLLk+U+HHi/iFClYI3V7V
8t600yRXkHLd0aHUJV+fF+k44e1CLfoDJUT46mjDX6eQJfKH1KhpLz9hsS4ElFvd
wXpEFZOZWYI9soZMtmvY84H0UgCvJhvI2DhvnFaQdPhoscL+OlLqy1gZEAtWQrP8
`protect END_PROTECTED
