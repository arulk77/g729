`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOe2cOT8/Y9zGx2SobqwKpuWZfxPGY+1zrxQZxOE8NOj
/7UOfc3MhK0IJbe6cOz2EZCWhaUNd0Ia/Ndg19hllIzdTrJkt/cdoEjgVLbGzWNc
JvE2YO0XaLyZLA0YmUBCn+VET6dZt6pfTxMkn27k/Fj98IkSxX81Q6BTY857OSsF
mDQqcMVg/C3iiUvww+z7dpmmuiuRtc5O4tQTpNu2uBFjvC5Wn2tVldGqD+udDNTq
bwVyntaTEAdXNZv2kPXi4Q/q5BAW1H+yJ0ovxyecDvGjd7gfohrsq7wNz9w9Bc3u
t1QOCXgHKEYxrhUPiommDYLoUHH9X9qo3EvacA7peVBCXk4hvdFNFqPk9G18CAii
`protect END_PROTECTED
