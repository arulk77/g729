`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI2Qz0daTzRB9Mv2xvDNd6ZEhuuuVhi58oM20INdniq6
90bz2wVONpp4KZGF+ToazvilxAsOxbKdhE7JOmhCQi8tZC5lrfElfNk1q1upwvOc
fP2a1kZkZ3gOGQ77buzPMoHiI4S9LvWtMgyWdZpAsEm7Jfv8xf7NtZFDyHzJwKuN
XIjywPCV1go0CYFehzhlM9s5ahELLTUtYWGyzpWWIUerls7kqxwKj7NKgJE/TGDB
KKw+xoBTl5Xg4B5Ju9XLWyz6v7GImRSbm9oMU95gQof4fnZYZc4kQ/imqe7AYz1g
OzQIh4Q9kezpRPe4stqJhbZXReUcz77JFhVYeClb8f9t7YCpI/TVedrlDqJQDx7G
fAokp0t4zyoSuWjq/qZIiK1awhTg2Uy0ZscKpLIPwutnDWbzHZt6Vh1Urqejcat3
JZHqvmuhQ3M4UbXiH6Oy5OtfPpUTgQ7z69AkAOvZgYbZqfI/iAZgpbU7BSL2jIPu
IyKNCx7XhcD5S6FBOeUnQ+77SgfEt60ny0ZDm5K59tGa2F1IpKdY0q+eHD7vuCok
`protect END_PROTECTED
