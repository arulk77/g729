`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN3Wuxkx6NjiOZAEknVP1izMOJCrY8XImVyd/nvI9UsV7
z6Owv44i0bPPi02HO4mMoUBXx4CRo+xTjfR64wThMwkHvQQSoB+2uXxEbEVLJ3o+
UN3uxfq8Opf0BdwxQBIvKtNZjgnLVlEg99UvIoyEUZwJe1fddw+rRoGyeqp+gtyc
5HP74M4xTR1wDJX5WChIXN+iWVlKLOsUT9vmTKqYwBPW4zRj81orgUzMjrnrMSDJ
xL6TdqZcfUIAPbaSwyuv+aDtOOH032X9kCuyR29hR9VnIhCLG8mR5odFGGYhXQWo
5Q86bi16WBnC6qHE23t78jhZm24kXp3caoJTRRGe0JdCOYyvpW/V/ykeJx9io1/v
yXzZaC1ejC3H7c2JjGH61PNFDQqBfEzldNPOgk+2YI51Si9RZ+PTbUFV+J69F2Vk
97bKXqwu/1V67/B790+na5wYcFCbeB2yNkdggZn9bEh3sLpEis0Kmt2C6WH5kjMe
wM9nIVj7YnP7wtOegmowab9diBSnCqcY3gKR/U9BmCm4aB63+61XJ5jZPSBNhCfJ
8ir28U3p5oi0irDCyJvhwjsO+R5i1JbGMPazMYpU1VNHIUkfqpQLTT5wt/10EmJ6
470luZ6niUYsVWnD5K5RoJMlMoghkRY+aKgCjBY2mxcOuobdIwpZW3Wi8tH8/ndC
wDG4/7S2hHn6YwGEJnaiJbkem9uPjUWo4/4XPwXDS3/ndtzyfk+KiEOWPdO3FRlA
GLPK8TvPLZsVA0/8r0kdaWEDrXZexyA2iyjN6S8kM6ehvSM33+zHzX5t8iCOh5iP
l/9hBaZUjweOJLo926AjjeCTI+/Hbwk061Ofv4wKE0w+b5k3zTP8Mq+YKi/UHo4P
X8ObIbiKvMvjwDR3zVY5GP0j6Iaa+i/fNGsVk2hTqw0wAI+hQmOBwUMb5mq2+9UI
oDYXYaHdf7Dkdk1IZZzsydK22CdbazXLrVyjMoa9bg/xrk1iWeWINebhgzF67h14
ec66SFQS8jrZ2Es+1+41xKvnm7Na7bYpi1t7WWZ3Tl2tFhyRAkHm6HUvDCWaRWzK
3WsFrQmVF7zvqHfdyUqv2rD58LoZhdxeviVLE5g+euPB2evZoy0TdDFII2um8UfU
dFeynr0OxtVqtt30C2PNToKfBKlrGAysaAMfq64XB4m3jvzu3e3bpBxmqkxubTox
UbzYy8qrLvOiDedSXZVpZ07gojKXy1KDr71dm4/cHqBDVf76o6S2kKT4l4V3ox7U
pbKpxnk1jVBglHnud1SQhCcAggubhWp5uYaTNgMztXkLjVdoufbHPyWlak/yzOVv
xKBVuEVoPAp/3Z/QeZnOIbu1slh2LzHMjE7+49fO/HftRjSsxOmfrVDpht6uQcIU
DhN+M2bVk029HBbM65MXq9/IDchoVpuvjsgS7sGLaHiV+cwHvnRfO16yKP3zZBQU
Dc6daCo/VNIqAMRHVNQPB6ndadKx49AQIrRSXdK4x+wUWPJLs/MhHzFaSbOTs+52
yv9nJJ37zhpSr3b3RcEwm4SOXD3ht3k9OMcvmJopIAy57yuZ//vKCi6ZYUqHucEy
z2GlqaoLeLCWC61VKXPpxZkmASMZNq9ey3c5yQo5w+bgmiIpxV3ihhTcls31QYkj
EwclUdy4xH7dJCvFItf1T9bjYep0jMsOg4vZ/mvAaN1qA45a3+Z/hgT33j0YbahZ
TrGxef6hWdj5Z2Zl89Q7dsjkvnepMIP/ZliJSc74WA6sEd58gLJt/xCkMPsCmocT
naHe59yaOwt9KqbCy5LYHx2ZjR0fmA15tYPJIbetX6kcSvYsZTFiVF3smSss71pL
an1phOstxDKCzEtwQIQWSjM1/9PTkvObxVTLnz5+oyw=
`protect END_PROTECTED
