`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOOEKX7OPVu1ZQzAtjiPUqrEE11/2pK2WE4ib4Yqsbyl
x9BXSmRKw740owkcvD512AthHOkcxK5+4ayA+GYZGxRRriRisCGAI9qfhbtO3Ug3
19MWFp3KLf4/bNzGvD+eIEYRt5vblfVA7/aXwtIM0887urc5Xdv77IoCDKLit6sY
xxjC4dNqMV7zk3Yvkq7N/w==
`protect END_PROTECTED
