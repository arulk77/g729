`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
oBrDAVsukBsesE8loqWyU8mXI1oSLEZ5YEGeqq7H25ZSwaNhR18YNo1lo4QtHx1z
cc7Gu8IzIiY+pVaW3QzSqiEXYfZv9O2qx39HPOFna2IZMkpf2D6LiCsf0VqdelWe
ll7JkIJGRTKxcg8Yd4EmYrqO08WPOBEowzZ54LxtHmDKpYpmcIwNz/1/6YFhmsXE
uOEKW3bMTTxqbhkYhXyRtf8FAMmWelgFEVev7JOTZhNheBpH1vVK199RNrNJbdl1
6b51kY5h7W6SY7C/OCmcuOoDGmrLaYbPnndgdnSYRR46iiOTdcsMB20cVNu4MN9/
IijYsHFU98phaFJGlf7OPfGgFYi5xf522iZMUInaIfkXjuakWQtAdI1U0jg5SwNa
k1Z/0ffVF9oSTFfGWSvOM1GhVuosrsv/Zl5Ugqfk66k=
`protect END_PROTECTED
