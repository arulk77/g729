`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/7jM8aO84GI4U9vKD87G0dfjiX6UD8z/cGwq/fnK1DJ
5vBGBZCbV1O+dc8jdI4fez1Ft56vVmwU9ENHYkdln8owhruT1fb9kRiA2+y1A8ri
KvgDJtD6bwasYaAnXb+ks0YTL70SCuwJ41Vnacu2FmdAWIvwCdHJpqmS9/UsiWB3
GDyXVvbCLfnEYze8f4JLiD1OedutOPaH1XbXxkY2Yok8W0sSf0TjGmMKT+2s3Avq
EHIaDthFbFm7TWb2p5gROcoTfcS4zhi+JkLto1cih0Ox39ZH8IEEdWVEx25L+EyX
iKIt9xq9X+4lgMKvQym1GcqcCmgCYN+g7mNBtz7RVa4opVEOw0aOxqcAjn6l0JE3
1b/3he/jAcUW438hfx17c8ZGfXLxffnjvIN4WzfTKBrxxsDODnopR/gX+qBbNfZI
ioXf6pN2rn2JEu8SDFhJSTOPpD/8JTqoo4i7haxnWR/WMRlm7rGhriz2FiQO+/ZF
`protect END_PROTECTED
