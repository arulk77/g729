`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHvXi1oeBQMCh2jLB0hvuCKwnMKr9h8l6JcPFP95PT6y
pPANrD8hfGxxKuWM4V5dv0pdj5G0Myfr1PBZWrPK4BOKjXit7/HhbS+wsfMo6WiV
fEqxxNiJnbs9itgCKH05TNFZM1XMcTxaoE/jfJt/JxC4IcJrkUeZETNah3GAikVi
G01bOgoO9NRirV1iQKFJNhGeNAshVSsjw7i5Zj3k08zQkxxMdWk9qBW00pIfo/vQ
ql0pIFhMpvscEzbUHZrA4FjILnRD8i9jd+UDdCiR205g0equ2JJ1csLKwW+PP2GY
DC9MR3nBfEzq4oNN0vUm29+XIKY76HaQquRZXn2g/FBkQ5K91ntj1vR+cUPCsKum
gQalQSk0qtz9TQ88KtpNxp+535P5bqH/d8dNOqVbW9vCqXMogExv2y3PGFvxi76h
KBgmZ/p4j9H/xpaM7DblyMWvf8DEpBGb1R+kIdW0l2BAxu2FXPx1GWqqW4vFyxqD
rtf8iodgsm/82TgACpRhg3UTtkkC1kRIWCBRVznUi9vwGkaIPiDv1G/Yit4eFnGq
`protect END_PROTECTED
