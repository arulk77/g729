`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKuSQY3/wX0/2i+QdKl2tM5I3OW0pjm8hPuW/4i9lpiX
wsrjVS/9yzt5WFWKVNrdnQXgCU5p7UYdGoxz4zJnNe+4Wn0Y9E6ClFZSr53ZcbfZ
KiymR9sq50kytlSlIKSqGBTjdzx6nuvkjAY2E6xJvXARIzvNFfvisptGi23pVcYM
t/CIfO8cHKrOxqUXIaQhvggRC+/zM58/wYC86jjKdivYOJJZfRc6dRFwTvm2tEyY
tZHOfdHtr/JYxbewxzFd+1jw4HZi4F0GsT3pn1MUmbCJnsOfmasBqi8CHjJISpfe
LOs/L23ksSZdcBfcSjzuc2D+cwUbHM4dkApKQUCPTlYyMgax9tibwxH314Bli9SR
uHYEtAH4HUyVN5UyRePkO23fVPILKNcbEm2K8tQt1bvf9007oPuOgLgoGgi+YU8P
FHgr/cLTJv1AEQdDbJvtWQOHYQnrwrjCFm28DAimsFKCcehwowY2OEV0+9qJuFdQ
kSmje3R9q3wz0gEXLMM+Zvozs2merZJSPTbnFGQif+bKK9O/5fCOMqBJlBfqslpV
b33Oaic7JWoPri5w82HGHl3+vf6SuxS9uges3webJgh6xGoxJnDcE1WC54wXndoU
`protect END_PROTECTED
