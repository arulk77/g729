`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG2ohsJfOujmmONG25MsSknAwVILEFbpnBjZVk4MAl6B
dOrdu492dZ/lvnICZ67flOmE1XfiOgXT1yu5io2jkU5vPVTBwHSF07C0x8jR/VJG
ByvPuJO7yGFt1qnGk4OQ+QABzaoqfXDxEqUj5iP3g29RFFKDk0A4hzLdZ8vbE7bJ
SffOyQWyoHJcMBlAfa0syAeoG5G7hPX44jpgKGux3lO/5+6F+XuD5NPKqB1shRPD
np5zPDaQb/CipAWV00/ZjhXO3C4qDpBhmria+79m8KERG3vugFwRTpngTHvmGfRn
P4ySXK5RHItvJJ+yBxEewjQB4m2MA+2QYjZwMCuWho1vwt7OwUtXW90PPuz2pOp/
5zBc8x8AAFfsVnVHpmUsI9n69iaJS0CqZDlgaiWa0VPZ3PXmWdRRfOVJkqGi7Fkm
PrVF0orl/LCH091BbTBioLvciXSp/B4Ls5CE/wqjko0GbkoJJkb1ZChcZDhceOCJ
KS2CoWlmp5iICw37wEEDuADUOm/tz/ng9zNhyj6R/lfWpZRBPpycjLWHXkJliEdG
c+yveUTpKbzeyVM2HHJfIgGfGk/CUyhKIOZVw/AqVLEpy/AoU6E6jLOLVgxE/2tq
0VpAu75vPjRNfEoYcCHxBNS1f4MYwkHOCY2yhqKMdbVLlbbNOj4KOJ6fY1ucOZSz
`protect END_PROTECTED
