`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBEY6zwzKLTNEWc2cs+xG5UD8IqLIFlip9SRYGOnVDt0
shYDXxzLlaPptrM/tgXWdesP+0UniFATAuREmamhEPIoE7zcOqJnpWcXdPm6OHg5
pStEmuU6+mwpB0h7Vq6ix/tQoN8x+nVNuaeew3GiEhxtxvvJeBARbcm3PzLytFA9
GuuM6LUle2aG8Iw7FnpjqVNULKKepWxaNodLiOHilXBd2f3CpGsyD+iMAFPnlXPw
bd3ZaLHRs/fRR8yPTbY/MTP97kU3CEhBM+myVCNpSs5hb0vaLTK1rXHyjbunw3On
8EMCCo5ZzCtn3tHEIXcBc55A2sIm0rogX/YmV7l+i3nQJiW+EThPF6RCVKJwc4wi
5Y8+bI/qofeFisfNGLv5E6GUUUXIkilf/C+rw6FJGle9xaRAWuYPN+9Z7TonK2hv
4FjW+f8uYXi6LW5IKShA2w==
`protect END_PROTECTED
