`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Hnxpr4IVWFyZd9nIQ33u90CW6ZpzB86PfVZXmRYPzV48/lji1sizM2U+2aggZeP1
44ThCYJIMxgwT0QFeJqj51iztUyxlmsm0axgnZRqXvgAm8IFwFfZdHj0ihgmaoyJ
gXAXuGzGvK9L0MZ0zI0mBBlz86GxfrHC5AluF4pnwW/CT8LPTMBEbCH0fCfXhB4B
oV0T0fvCj0gEO7pU+HdFaXY0xhNBo4fVHmUgGdkqkRy5T6DoQFLR+6sHTM9rTGPn
ihLhBGDfMYkcEaf+fKVeS7MZSjEcU4zg2bxGb6G0r2L6LKv7NwjHtyh/tyUC+dsB
`protect END_PROTECTED
