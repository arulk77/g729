`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
UgXdLbmEAKUu7Z0Fw8YVuUQ52uR3CyrBj9xdstIxCKdVl0Gj2O2EzvBcAu7MPVnx
GtquiA6vofti8qLnbhLpJUzXe2UzjmCCHNTaQBEVgiV/rI6oRpfi3pGvH5F22KBo
OnYjpoxhrKWHe3cyxxo8ewW6bxTpnlL9NImtIYIUYJnSAnfq0oYGLCQEgN/pDE5b
BH1LY3vi6SEpt2Rxv6v1iUvD0VqSylBkKaW8jjeq6y1kRubjFrxvU3Uqc6Lnro+U
WrnyAxasaV/FELHEy6K+8QJLpf6fxYh8rUj4Ps7JRJ0=
`protect END_PROTECTED
