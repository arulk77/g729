`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGdaIguYtH/fSrLeIs24Q5o2PI02f9ECAupW2BwhJ369
TNn5PadYwnjgp8GiWOHur3dUR3L1a5VvcJ2nJ6WX7c0rDLinz+pwOC0YQkC3dU/M
HqsgO4i2p85BN+/9d0aRoDGVoIO+c+mlb9+frnywNAAlZ3wCm2nby6teS7+hCfhL
nrUhPeiYPEVvbdFMuJaGj4qkPRfxZYFoYlSvAnu9q0PM1yqkUUyHZjYvzEWOuJwp
ZY1DjKvG5wmS+aG6G5JN7AVu29kFbe89LDjVSKJFWUzPnJLc1ozdoXcePmrJiqwm
M4ulTnHVsLbU2/Yi7solcg==
`protect END_PROTECTED
