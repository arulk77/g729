`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNr46i923wsqyDCVkzsrtqcDClrUgNMYfBOp9awP8/Ms
PazU9qoXSnGqJIsD2V/S1qDGnl13B8/YvlGlu1B4hET1ClMZVP/5AdaSV9Lx9qDL
hZDN/S2cF+YrfJbeVUCPm3uhA6p/R7Wmd+gu75z0zTVak5wWSFTrfO8LINQqkp1e
1xG8D6ufCwWSYTvj+6jA6T+RU8Rh5dnT9fnzuMmipwevO2liU1Xp4Z72DWlC/CyB
XLdvkta7RyJjtaRFQ8J+fsSftKcxeeHnmG35EYly3zCS70pwd2WSTY76y1/WvW2J
s6TFwGkAAd0TSni8zbaBjP9L6tAioaMQXNLRkbpFgSq9iY7LkZhe/HjcZOGeCscZ
OoGLqjQpbCe/sUT4oI+ovg==
`protect END_PROTECTED
