`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNn1hLtwIDas+es5Bzwd9CSUHMPx/5d/QGmG9ZbmISOe
ok9gy2tzU7Dwg09w2VVuOlXgu6TBHVLCeR9i3iHjEYD7UzRq8bXE8OmjHu/SJj/M
P5O+EfHpIyPRD0OR56WZj6BB0pCC7/6c9Qx0NFZVSL2TJTzHlh+ym0eGcXbAbAQK
AQ5B2kEjRO8EC0Gjy9LEHO3iwhTX/ihBh2r2epZospO2CeJ6bmfwdJ7suR0qUhq7
`protect END_PROTECTED
