`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Abm0qZdrzc6MTWUBvldBz4v9oFT1D7xxMPDLfKqsaPBS2UpqxLn3aoEFBXBG0e3q
QFxWiFQBwreuY8n98XiSui26QpcrihKBjUNc2Y40WBF4UkXo8pO891oN1FDVqDOF
TK3Jg3dXhyyy+NuBcDJ8fcY8Fw+Bj38hhR0Bqa/UZX6wRmDfnOkQDW00TnhUYeYx
MEPXNmLyS1h4BYHf4ZKryfyJRv+mZ5Ik6YYXnZGxbmbfkmblFQSdPuoRmDY5WEbU
spPN2RD2my9G6Cv5LRqOQmEBUBi4PUDft9wQflnGRWqF0PDo/KCXU893yGhnSsC7
NNNEUl4vQ3a734YeIb41Cye3/z07lMNwQcE/t+jJyxc=
`protect END_PROTECTED
