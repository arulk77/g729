`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
UdngEdlfHVuFz91hw69ZN7dlYtHlTtyAj6i4ObWPQDqcAGCeiF6IYKUUnkBZeeAS
wbyUSZHLUAotEASuwr3nrY+Fuj03s+2N5NM0qWxvpq3Q2Ktg9+O1zAtWxPS7Wfbq
6LuLRZTQ4xEcc4BQTqA8e5I2k7Wxs6nYczQSIP6OmeJNqtpv88gABdITSq5miW75
BnwRPG7Oae+q4hz3ZCsQ86NjTirmilv+Yuzr8TGfC77aRxqD50D9b7z4jlKBGveg
Dc2PO3Ig7Fhe7aKV+dsFBLw7aZMeRk6Q2jpr7ASEwLI=
`protect END_PROTECTED
