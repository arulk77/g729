`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG/eR9z93pPcw9MCpSzeua2Xdv/T4F4v0nvGfsRi6Uzh
v0Hz03vz5mS808Ejqk58Ny+zBIJuIHlpz2zq3f0i7jDjT4d80a+Y3G9qzxoO9kC/
xAPE7R70UyDeHlV44vWUKJ1N9Rk7d5GKWWiQgHgRRxrj5o8/KNSNya/v1WF+48fr
XNFO/oKCBoD7IJ44lUdayF6hvvj4ZYeXTGHGYzWUNnzNwshgsN9GwdEVnY68Ul46
k3xFH0Px03uMgoUtEnqlFw==
`protect END_PROTECTED
