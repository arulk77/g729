`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
6VQBftK4xOfU66SbsPaPIX1Rg7PWie3Y2h47ykji/rSkFx76lRjpTr3tW2q9VY/4
jxXb97SmJRaCnkBZ1h7egB5bX7QwcWZK8mV4d6VVQkcY4FDyOWUVQzpBqgK+SdFJ
tkzGWqfITF4fbmKP0TzunCGJKN/yhorV2KjxV4GQ9uFKX+6DGr4y8tSsRy6R1tn5
XogRODCK+Eqpb15uO2X3J1AledOjvUOvZ8Jp2rSManzKvZqwrCsfn/nrZEXQodtQ
6hnycNevdh2ihCljDah1EYIGecuy+efuQ85f70llBH0PSXQpkEcVA8WzTgzO2hqr
kmz5Oisa2VvkhVzS1RMelhVA9ESBhVxSp1z/uAI1JJa9ozhWbF3alVq19nkH+xDN
zrb/OvhltY+dIlTEQ8DYTHgL70nbSPDQ77vRjpHaPkQ=
`protect END_PROTECTED
