`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aQBjRZIoHZmyZLcpqkkLaa8Lc58zt7XOPpIIajU/HUXm
8RcBmzgpH+qQ4CEn2h/JsG5f8ZZPWdhlXHLXOqLOjN0Vbl6syyJ91LVj4X6V2IDU
5HOaM31T7TbTKJ/9EkrtljDit/Q3gpS7cEL+LM1LLlnIRIt7E29jy8D+wsQarUM8
rfPcoFk2NmoGtkD9ZmxfgsEmo0nCdMoeq1XvPvmbf+HzUgw1PdG4LbcM8EYUBBfO
ulbXSh1j0f94Hgteokp3Pkkmhxe+uJi+9LDn2qZs2jslP51SP249Fz5K3koPrpLA
AGVij2NbiYdNf6ATY3aBFAYXLPlejb99VnFW0r+iRbRwqnqNT37/rnggC3loBi/2
+fato0cY7Kzl5xc7YX8tlDIq7BcRC+F0DRVvWxASEzPDzt9zg1u6qrVcTmuRfZHD
u0pCoX2rdavCWL9Y/I8vsfdhjbhOh8xMAQ2GJMEQ59r0XVzMAzEGzgH47gb0SMXb
guGGcsR+FihREOZoPmZkjb8zkKX5mtegVRmLlNrG7H5+rpeuEXv9dENhGdMCukUL
hOl0UUy76lW9BJ3Ic95R2p9XCemc7TUAiZordDdCMocsjscBIrv9VRVJ7SF0wq/0
beX9kzvPZhshijgAhdmt5W5UmClELehigl4IU2dr3lGgjVp1kkN2G9EQiXUKsZax
RX5DjtmIHeD+DHAMeuFuwpUclOx2fRk+uBakhf5gN7TSs6guXuwJ6pmPLbFQ3Bqq
4HdCHXCMandVjdlG9dOTPLOxTCAvUc2aIyNWsMM8B3GL6EkBadkadY4S0tLIF1SM
rmIc5n0STc/zUhTpyehJvaEdvgxPn6bu+HLFRo3aKaL7EuMmQotT5dpaL1I6aawy
zE+pIpy715NYnLVmTE7Fb8xfq1EBYcPKttlE8t7b7hHyaMDLkz7oUjbLMv8IeJVp
tLPdEicFcErrKOTyfpEj/DoT5+askIyLyAB6kL6ogshTGlA9spvvEF3ReU0U8CaU
8LwdwpRSOX/O7FMu637XuODnvpz/mBjnSVjh8kqHjZhgHiJ58IRz8GKT23JrUnyD
nkNvB3mdUOZWU2UGC4cN2J3kwIVp5AzJMjlmIDnwPCEyZULB1kDd2Bj8C3AhlwRX
L8oH7K7wtACA61cNh6Sl5uldyGaY9uG2BGQhD6Nn8d1YyTzgBIsqrFT+CYCKbfu4
NaNgLWe9J5rPJuW+pTaks9mr9uCdRA81FkqeD7wNW5+lIbU9vuAxZZeu0IWeMInd
tHQl1l5K2qujds9MuysdJX203flAEemBHPMHkxosfiOfU3B+lTlkcs/Ei8awSJKH
oxZF6zl2bsyEHphVPOVkY8xTksyNBrxwV0c/YfUloi8+QUlp84IzL+yS7Xf/lEYx
UEIFmKnclPqXZPA11mLk5QU3wpN+oaiuZKX/ZqF3vy1YBdDd6dTzYz+xlyVJMer8
Q0FYnXguGQBjHqEBlEcTsHRihSEfh1xYIUj9g3RTpROmDhnOwnqwhAN6JWBmDWn+
8pM7k7OwWiEyS8aeFHUtmR1GJw3zfU2b9d/u61v/soo=
`protect END_PROTECTED
