`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SXUABaYrr9lRAZGsU1+KEfb+4sYPRVfVOJO51lw9V2Ia
vxvuCZTOVl3S/+iMrQRo1g64SFbM8TX7Uyzphm1aNEvipuIBa0JznKJemcPAE9xz
lJPwZO4q0RfAzM7VpaapBli/eSyNLbgcRW8INCBIwjdIERwBw/3S2EfcIn3bK9pj
G/7r8tkUZ0f7idDaLDt4v1zkw7jhBw+snbkbnnMVRiEDCDnp3VH+Mjabx5pM0qp8
fNYF/UnwO6ng9Io7alm8G3x3KVMVLA+gBb9yuGpx6PVvcnZA4ctQBXKsuyni2O6I
TG4mvh5FOVzo/xMdkzEtJ+QpHCPwfD/V/P6/HlsPIi0gCe/SaZRfRlf3OtgFvlkc
BlmLvVaZZdVnfcdRaRxvQoh3YsQ+LugXRorC1Dpww9Ux3SsP97q2baX7GLMvP/Cz
3YZSS6UQ1C9QY14ABiAn27YSP40b30DraKjx7yctlCzMO2Mp+LrP0jVsvy7VFZL2
tIgZHtUwl5gPFIQmbsDezC8y4h0aFRV+t4og3J0IE7ljUBQxj0iqAu8mRPTjSJQ/
0PX8zvHujVE3uhaJ8Rxfq6iJTBIo2fYi8tDdRbqgyI9dg3cXqavkEN4eeY0X+eJh
89jcz78+Zhn2Hjzq9PRyv02YR8+whhGwobvF5f3cLwNvsQdxUoEq+uKF9jPji1Hx
fgfY9y40KsPNhz0KhZgw5pZHnjBeoG3MhbHIiQu0CUyQhY3c3ds0BC2q3ySfg+JU
d5LuVRHC68AyLaH7tp1Z8qHrH2RO9ZGftphE2fkzwjvGYUhRhKPTrC5upf5ehE01
Ph5WNa5ftfg+2tWPhQoa7ZkCkLSu5YQlT6wE+4Dh72wBKyN9pvVvzwlhSgXgEDs9
hf3G0JrxXcBVxelMz+3qdBLy1U5Bmpr0n/73kxEm90a5t3ujexUwxAIClIiolMES
rMvPV01T7Wwjm5g5kx3ynFmC8WKsbKv2ZGOhqqhHlXsznbaMwEe2APMYyaITh9CQ
SjZPGZcDOYl0gs/gbpZV6fyIzqUmLo6wuUK0FqtC+6YLTYGCmjDcCgUYelGarGJd
iLXc7BTJRQh996bX486jFrjT6ukXyywhMbAs2u1xXY0EmB54+N5yenq1fdFh/W7T
c0igJP9CZevCcF4v/YJSim2O4pZ/0UgzozAuIOr9tXbUeQcHxAi01sLcIjxyP9Dp
wBjaaJ4y8qsbFDa5xtDMGtq0CcPMrjbb/fCvX/QONAeJshlX/kc0cCssqxB87Ik7
aBIgcBZkGOhHtFhrlggPs2ccw1EzHWxE93XaaLhTiNRBur3lU3M1rFvwqpQHWEbN
6CUMulnoaAdXYGv8p850Lgs9TiZx1dhVC1KQPxuHPCj1jdffkAC2WZ8fNN6oIoHZ
EtmUI+sjc6pGafg7Ff+yb3A8M8OZsazw7l0l8/v58oflmerDCMjScP4Mlpf1zN3w
Dl6GuexEsbV3VPN/H/zcXmBaEA2gc7akmEXXJMLRpuu4XIVhiFcgrbIxxFWFOzZQ
Gk1mgcn4HcCziqU03xl4e8nnNBuV+APFe2hrebsTS4WVXmeD4zYO6VXnYvz9fcut
iHg8mVLMd3Hp2IcRd3bGECs4pAbdlLk/cco0cTDaST8yfiekmTKAPahwkkuC7Lk5
iYg80qxtnFCuKVk4HCtpvd/gsidSoCcXV2M4Q+TCRppkRH9wmSPno5A/hGpocpYd
5kv0jsqtZ5+ANEi8FzOJyD1yeDtbt4MyxtfuegLLrPV38sl0LjwY4fxiBfWJGKOD
8r/CcfjT1MmbupI2YzD4kPyh2+MBJ/YUpac0xfCkEgEEJHOEAtV6Rsh1X0czzAtY
A0ouiNJi4hqUz8LuL1tUJpuFurlqfEvDgdJIO5IegFn0eEc4+ihOXu2+xOxXbnO8
5qEvFVDh+4vdjNbV05rPls/kzR9wNGX1zq5lncklbkCW5RaJ47MSwVnkXzzxC1iA
USr8Bn++RCmwykN94P1GAfm9E7xSm4gzdHjFlTMo7yCpQKnavYrqKS5Jrc65sXsR
JkbtLLrTDACxXuvSn/2NEfpVknFQvCY1MNAwYhYr2PXegkNg7/RzLXkPjiOhSowu
gGIh7+wXvSv2oosSazAh809LPySellfIvsQmM3erKhLtlr53LGVuMIztU/RB3Gxg
Nn1AbaWmSJoG2UvXXVjOgiMHdaj6at9qsXKq0roHkKDo9e5fPfHyaPzyz7OIVD4g
PY2qqYxSWemsAaGYg/QD3I4IXZx2YuFFMWkmAGrjANHQT6D2UbZRY7PUXxOceRdz
M1ILEO+xt4nZGsRSgYsn+Zk0Um9K3xCShOUuu/F1B0d4aXjjmxfOS2uW8+oarpNu
ayx0TUQyNts2ENaeslyrkTc6zR19tYhZCpNZEPSESsp7rQvuJYlGqrl/8cpY5uYc
Z7AS7IuC5ZcUrNUIGwLgSqBJrmwy2mTav0Vp3P09zc21AoRCqkPs8XlYCVM4cgnP
oUcHtvnr/sMmcWLNgsascfNdgUBMDVqR6G9NymjtlZjOJMph73VagTO5Bdca6s92
I4zEjuwa+BFzYuoWBX/Stu0VptpSuFvpwwyZgKaDICxXODuPCuV+IRpk4tedJ4km
Vc9wOttHq83y5SKqGNNsrBzd5J+Cfh7BlZKU5lN+2Q3uKBn1dojKGTucWybXGH5o
Eq1PjNYnihXeSruFN0c2pwBrE8p+SAl7GIcS1i6kJBjP7USLdqTg4heGxbIvd6L1
efqomJddbTNSWIBN+aQUplvbgtbD/D/yy5O9+Rky6unRC/P/443+d9TbPEriyEYK
GoFh6/Cu3h8AzbWPU+aJCqqEJdAI3QLeBHqRfZB4QAYBxoAil0QMHz4rN/7l6AGf
UI7dHlPIB446HRahw/dFk3j2OIN4HSyarEjwmtdUwWztY/W51THCs49lVR9wdeKe
UQJuA8QgD2FqEYtUHYsYq31ZCR80mSxVVQrtCJldWq1CSXjE0QEirUzDjmeC09u8
DkaLXsxV299j6sVjW+o9nV8a+yp8sUrPvAQ4HaP0tkviauK9OhyEb6BKQLXkhBAM
nASBMHrdCdr6ZZNnfdMzZBoCwAp8YScQdky+rRYzg4xD0HbPKBMH18Q3eoc2j811
Z8VIRGStgI2hjuMxcp8JHPjftOXtgpNXtywnC63QjUMoipqGTVSFeP+qcSdvUQPZ
We0MmD4WDQcoOXsbLrKLWx+cCR2gOt3zd7C5kn1AuTLKqhUt55icSVUdoajr7/aP
gDxAfVitrH+GZlZaZmT5OsRD1jdQIDJLLDz1dmGn05CZFE3Ia4vjMtKIJAMi8q4i
YFI4n67ZME9Ti609N7CQzWIAYB7Rwr/4tJqOXE6tJxCspIKJup/+A88AGa8I/eIj
41Lvdg8B0wNF8h3OblkMpZImGRvQdlOfobAfO1R7JxzUJCHckZS49on8VBL8e5S7
wXIRyf+qa+uESGOWc+YQLO9Qwdzi40y2EG97/WYyG88NtEv8p3wD7QnamDWf5wMq
CYJY3VU3o69CDg4vkhaVok9mxki9KWuQwKUgC2aqibm1k8cJygGReVwvl8ux2Mru
pkD8zHxM7+P5L6QmJx97PRoFNRSBWh2Yfa9gpy/DEtPFcp8UlD3yorS1J8tlL3B0
WTXh8mCT94Vt62i0hkqfq/bAzSIx+OydMrSmZpP0jEVHm2cnaRsFVTdr8yOMlmBl
7dM6ERC+yB/E4LvgdJrNnHWKP4lmXGXPHz9dQwXPlAMr58/rIjFpLcbOUMn225Q0
AHuSNdMtJN3khvyFyyouK8kmxmtjmBMEAAK6Ej1kZwyfn3UvjnYFe6bxOWetKg9C
`protect END_PROTECTED
