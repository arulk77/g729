`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGWmXEx1O2IUEFX5cE2Z51aKQLZjJJIgXiDkpEx3h6Cn
45Dsk0QophnscPi/fdQBMLK0lEpmbV+YlECIh7PxDxuF8ia8+jxZCOgvJQe/stKt
OuUSQYtE3PVH9FdLN9wVCoHqim3QWVVecvd4Mdez40X2dccr/Oe58RVZz3sUjoCM
4PpwIZGxl9QhCLajMsWTPQ==
`protect END_PROTECTED
