`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
XlUlDuss/1GsxicsdH3PmjRzykNqpwFAmnhAhrxqgC3ggOXfCNMFk+63Ru240Obq
eUDMUAE4pQ+nbyVvwQX8UIb8ROJ9fSN7FQ/2Up205LBLU2YAddsm1gz63XXjACZw
1lCHYlKRBuEv6PwOdGO4jWdjCCoKehXk+vVzL2NJ5pAQc/VUFkIRm0+Jc41c7+aO
`protect END_PROTECTED
