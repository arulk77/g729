`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
if7OW3neLerq5QTb0GME9y4EPbbW7yD/SnK8eTFcz3ZlxaVqlqB9lX9TUgn7i8VZ
NS+xwCe2B8K6X7LS7gK/imCymf+79WGC8PJAq7gSYvVI13aKF9CPpeJUFh+wzQ27
GmCQreKzXcmBb/sMSqkVvGRrdAcpl8FquNhmaeO2HoWb5LhLmNgErbRUdManGndB
PN2CZrD51IK79GeuPyw8h80yGZzCjVpKFhz+nbi57zcwO5PEtzI9mEJOzaGpxj2L
1VGasmjULJOMyP0drQ1lrrTRavinl2M+7A4MuG1INUV0hRqv4jC/OYAHfOGlBTzp
`protect END_PROTECTED
