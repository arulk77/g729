`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAU5iAEZydJ9c2UicxzDICuM5Il7EqDdbwNE0jrKNt0Cs
nnD+5t33r3pL2ieakCbdixu+eJr35hcqQPamwjrAXYrUGr66h+2wDgq2I+cPZUM1
qVl5Ej3uOdvAxU86yy0PWSQetNe4axZZeOlJM8v0ZW5EtfxClwKenLrsmHCwJY1Y
pEfMKsA2WhlZrvQMq1D/hnSVug2nol0nl8DYIJIcwlnzYme0dNipgmvIUcJAuH+y
KG7ylpXxc9Z+LHxokNdI1kDaiPMRWxOQr+kfKJpnjaNKy4fN1BBJwOjtnw3M1w9d
WXZPgmWdqISimP/ltB9SvKa0P+2Nec88TzCqAfXWFSlO8RivdfPixPaNJ9VhCCTH
+sz59p4ILpi9X9p7y7jYIZIvgCdfydIWbjWA5UPl5aRdZHjG9j3jkqAKm/2/mHka
zDflmtk1bbohiLO+r79YpY112GqENjZjl/TDVn/WBQmU2kMDlxULyeu48pFxfkg/
u0RtlDv0NDUtG5roCqosryFQWD5QgizcQUaS9HsgZaRR4XRpmKhdmmEADP6wmrvU
A+h8dhoPx37Z0ePDlxJsN0sfKAkX4mk6L6pGWGqHtS6e9WbZ+W2k59GfmoxTwPpK
bOQS/98CEFtWgvZAj/gcf9hf7XF1H8b4LYIs/W5L3QBpGS0+k3bQ8V++9Q1zG8Xs
8L90gps0GA+eN5S/+DxUPyE70P0kY96aR0cil+PliNN8/VddPYueQQN+wH+MSpTU
W663fhDexiHjIWV57gNA1DkTD7kBwdwBzahnNgTSlXvkgEOg0JMeIO5KKpHZOArl
7RK33vl8cwntZHbogr8ZPvOwiv78hlxlcoWc/N4DGc7Zi8u/7NeQlKIQfis6RkDq
LomMhWoz2VwBXJOAhjn5/s72gX4sYQWBzp6fKwzgFc0tfzHQhhr3OdUEmc1O/XHA
Af6E3FIBU2HvfmpPk1stIyMQL9oQClN385qLP0N4amU+phZjWXQNeWbP6C4B3LKS
gqoh+UNRUlqIkool+g2CbSulRbIWqNJP1QZJtscsybZWOd3CF12NUKiMpSW2hmqR
3A+JnriQ1dwNlI6z7S2/13lEoStIOYNp5K/akODBn7fYntYgIMSxnxnP5qDJl0Eg
kmc+QIZTJVncp0/HmGR4j0U9anyX6wuPgix5QufKQTKLyPlt5MGP3AdN42GFu0Io
vnnA3/FWUoOE2zfLsk1GaQ==
`protect END_PROTECTED
