`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHdh3M9JdoLCGNmXrEATaUyF5pYGGxWX8P2Vk/fl3ZPo
NoLMmv4JNzc4DNxB0WdpTsBhMd7DQF8y5O+QGQPZlmO8sKiQ4SxI4G1PD331opGb
ogVfU39gQqmL7gM3DlYuyXu6HQNj3WNknS1HP476/8Wg3qK0+EdBzwzTkfaDm/UW
SuYrReTazDDCLJkjx1bRKJE8Y2AyxqWu28cP2Xut8jdKRVJe7xAFfEhnxn51JXbF
QIOzB/KLkksV+OlpFiRFBbPSRgoUnQNHKPq7vduOLatdxn07h4YU0lsY2S/Fxmgi
Xx7m6EwJhm3xbW71rKFAAQ==
`protect END_PROTECTED
