`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41xoT9ClG4Z8bqoQCIXWQrNlI8Qqdtqs35COopSCQDWo
Nn6kMiI8LNEmfj86gDscdaulIbFLAnNXqbw6NNRkmZfrGZKGzGLGppAV3iq6zgHO
+m4O14PWpNIB57StGiqg7FfUZOdLjcG49OcWV6ChnCU5ccj/gH7RQHEs/3IZng/8
4alturZ0A++d/pYILghnnuWjP1z9oewhR9SsVEpAbeI5OrYDGgSSNEGiSIzcqe1A
pu82WvXvY10moqv8ltP1Hsye7rBpKToJTBg4dcgPzyc=
`protect END_PROTECTED
