`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
XsXGZBI/x+yr0zDcx06S27jET9ITd8eNJAjTiA9v//ugcR08f8Q77LlFXsUGsPEx
/2Ukd8CW4KBcCXT+2XzM52Oos4ihmz8klj/A7pvfIPk9nxz/W/gNJQ+ADb8NlhUF
VKfWReS7bbEEqapmNU5owN0bkMkTElXB0AeiFAZVtMbrHtSD49K4kfFyiqkKsbhy
`protect END_PROTECTED
