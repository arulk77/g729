`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHRLNVq65TuMHDchLpWLcn5b1lR8ylDkYTNMow9pUsE4
Gu+A8aCR899Tgarr3t+hnrvjb41IMI/r5l0MJvdKUdTBh014iTlslr87A7q3HXDI
7xSsqx3bVVz7bix3imvGS/sEDWHVX+7jNPWSGuK9Y1m7XjgoCUXwuhT+Ejg7rtcv
CFXHlD1Nrm0o+HCSxu2rhLgd0koOg/vCOYVqDsCB8ErD0iR4dXF7poH+G/VSU3pD
sP64OHykFn7wbkmSK/k6wZxMmTujgSMqq5AI/jlXVWgvT5ZtdNVNXJEXkkD9hxwn
B9k7WN3r5ZbC23bDplc8SQ==
`protect END_PROTECTED
