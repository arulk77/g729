`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C5Q9JLe1IAhy2tftAPYXq2lPgi/4fyFE2h8fMU/LqyOk
H8NaFxUs/+zHX+z8z9ymYiddnRVtprZDeYYBV50BDlaYfw8yNMj9UguI5SvAJVL/
pEEj5c/vE8ajP+qsxPzkQuKAvS+MOzaPdyzHFKxdCqbFM+rHQhCxKrrghig2TibU
dCgw2EImE03Qjw2ZH1EBIdYPLsoeI+Up7iyAo0Wc5KHIopvbuxIfuStvne4is79E
ltie1HtCcBvM+YDhXEgNft38uxg4yqM+ucDVHb9Z9SbOCdqvw+06tEKACRuNSwWb
HOuXya6JSMJGU+MeJeTxhrwDGds6jHcfsG5iQ9rSGGJWZwgjQc6hB1YRwKHQeG4m
KJQJwTmHzZERDoy6X15q6cMGTxgivb2MnT/ur93ONt9m/EvJqun+MKevVl1nyvyd
SQpfFtrykFWqkc7W1CrxW5cXzu3juIk3ywOOdYXvlV1M27I/cjlErt/JvL3otxt1
4ld0OhHHdOOFrmKYqvcZdasXj0LPvcKx3HVYXxS4wsFt0CwfjKI2ChZUURuVblhT
PrBqAh+Q4Xue+ILU1v4mW3hj6N7zifgfHUuX7CrIvrXj+ePmpQFmDk8b+GqhooVn
D6nrxiUou/UK6ssDEPMZ9JvJ0gSw9G9O8mS08pC2bHw=
`protect END_PROTECTED
