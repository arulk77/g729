`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMfueTHJUqRbdiX/4UEL4bj6KcApnY2ZSbMovj6qEKSE
/cvbgeM18BN/uILOrkxYdzQO2LLcyj/1eraUGkNrq+sXAfusjpX6waw4YpyOROqq
+MQCUak8igNt9yfi6n79EsOnsxeMtYzlCCKFrKLFKpNFm4k6PF4TwOBv7wEyDhMh
`protect END_PROTECTED
