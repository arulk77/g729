`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCN+zQxIUoZg1xAQG+IMR7TcbHXUkv2zpwJ2xsin2FUc
tIFxYXpc1/r39BfUh1JnVGOTI+BYo1d5bUKDkc1Ng3Fx92e11lM5dtqU4p/ED5U2
xq43fHRrz9/IoFGaMNIaej5XC74JhHOQOL1V9eDrdyb6VjKf8gUG/tq2WGrYvO0P
`protect END_PROTECTED
