`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCwYLQnhoCl+ExgnB61wsiqh6/LK1EnVmxVujIODNerN
1LUTEifwPevcWfT83LwaxmLTX33NLt4NR6QTQmROO2FXRh2SRZcipWSZXQpc0Zbx
3hUfXguMWFWCYCa4u+5lc4wiLoukBh7ytsog9+OdrycusosKuWt8fgqey2ZteX+g
jPReAuwth4UCtHmrfrEhdo9ZZYD6sYiWrcvlBsdwIZ82P8slNQvLzPpnepj9UTyD
R1Uruye4+ewe4GlbZNpHeN6AIsZqSzN3twRIxNUc7Phh6+AF3uAp0ALfcg/IXv4+
0g6Ewo/jso7KPSDrEmVMHOJnGU32PSvj9pI3jLmVz4CWBeyH3a9gYd+ccdDr/bhn
N4Ah4ac6TbbeM7RsjATmKw==
`protect END_PROTECTED
