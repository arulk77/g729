`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40t3kuGhvjfUPItqOStzM6Yl45QrJ8WPaJ52LCCM+0jV
mVnVIowzk3UbqpANJKE+88nmJ2FI0500MgKAPWXP90mqDKImKokpGUrRHFjzAk94
hw0GLr7jQiOZs/2bp78U5FtPsdxAaxWLv74jC5b2NeyGKZKs4bJ1Ng7QfUovTCpO
GqRgC+MlBXABGQ0MxGbVfznGilM4X9cTv23Gt09QDyuYOOSB1FS7eLWWp350P3+b
wJ+7gmwrqr+vxDSAY6oxHL+WDOlVNLFYCXOAyx9oMik=
`protect END_PROTECTED
