`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIJmQyXQCSDn1msYMJdhZAQ55Gz2WadsKZ0kscgix4+i
lGpq6cx8nm4aiqspo1eM2aqX3uvFcxjZJ2aa94MFBtyAuIbXSc0WSCczjZs0uyvd
GhxP1QYf7neKej1NuzYwemS1j8Dbkh4jgF5jwXyH8fHT5LZO3s7cETlNyrpEptX8
niymbnjD3ypwLTSvNznlhA==
`protect END_PROTECTED
