`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C8pJFH0GD4WhpWC0x901zwUaEWO4qC5Qbd1rMrq30Z+9
+LlS4LCe8vfJqDsYSHuouBwfhPWwVRMsyb2ho5ZqfAjtkF+WNtfRsVi/EEY+xPRV
okOVDyZTCJNGUZlVvb7lq6rYGbaExDsrE/gjOmEVTUCatMh9jsn6LbJ3FATKgvhJ
MwvJu5dqqYKBWB1JG7NQQIqCeS95n5PT9HdpFcOVEUw47QYHZkhBZc5p4QyPmi8E
HIJHf2Uxhx4nemVS344y9Z7DXy4e+tRPZBCI+aaa/na+Shd0kJLF6MfhO9qbl+WP
WqHOEUsBuWmGzU4ugjMWZxS9emfZ0prMZzVHEs3doaUW+/9q6sj0upE4DroOYT0D
V0T55YhAm0MZWjgM6ZGuDGjccPqtODrWgC4WaXTMxLXXFpWS5Siy7QeFowsRmsXA
JvhlwUtFWtMWnfRPDBG9t29McFtCukkRAa0N6wMFGCMqvtzwQtXrV0aN6TVG/36k
4LfSXTPl5PlaLABMsxthI3ixs9ckhnlWnYOtyYFJTpTZohXBS8GFFmjDWMIjsArf
6huodjhIqam8/Jw7GP79yBPJMVhTC5F6tXBGaCsh2q4vz+5IC7BiwfU5YH/T4KCT
BcKh5J18qAoETw/0BCNOH8fynQvEUeTnkM9qB70FsXe+Zaeo6Q6gxIxMSmNrdKfi
/lderYqy4pbxtTW5J62iTp1oPKUlRsuCEsd30VkKTIVKMN7FTAIa00EXlcAjHdrL
ffMdOmG2WWnuvyED+p7PbtjI0C5uZZMfh+yCKcgoHcj15RfXmXl5003ywGnksx4V
r1KbvDVliqbbNpjj7grLNnjzH+y4iWt3X9jEohlEgUToEBmRtMJd78QqHJI0He4I
pdO3PGIy7zd2P6Wap4/CwhjjfiAGmrHQmIFuGdXqMFu0g0EwBei8oIohBupKwrrO
LlJpR3OwvpZ1D9n0c0zdSsSwR+a/08rs7jrq5KbsfEckKN4cYQetSJZ/ND5a6SyH
EXdLl5dRmvcm5vtTh/eyrjzbu04ZjRAcMexYffa0fz2soG9tvOMSJTiswQNU7Thi
HO1Pw4HIu/LyaispsE6oM/m437zI0J/A9Pcbx3JlbFax6L6UhmnZFdyvM3k/ziAL
obpgIUhh3eUIjLK4fTpN7NxWtCsukW9x6Me2eiR0C/XVrq5VQBOHriCxwHcAUZ+7
jRk5zkeNBePPgOMrNoeIpdncOpaqp+Y+lFwYgliYgYPQPebBngYVlevDDe60Xuz0
CPJDRYNjUdnJwjtIqB1ggrO+orXlLemEIizUwtWXqpVpQGWYnZiXeIYcYfowF5JG
Uzbhyzlq9E3TUPj6i6R7PwZEHMjCkvcOjhReLoXpCDPT5cBGrXFteUhHDXuHsRK0
O65v6Ryp63byaVwaHIudmKGcBkqAFVf/gasEgiro2mX/wE/AkKWSSnmXNZlC+bQ0
8XczoMXfFDStz5cwayiqCkjI2Kc0A80WzM2bRuCmkGJVG/7rKbMKjo0WsVxZhIWs
XIXJl/LcjVusArPBY2FLdxhHK2kSJCYuOtcTs+TlLnb5y3hAUBnS5Synrf+uUi+v
dL+is9XUZY1KpbA11njk0PpKE8lJMXQYbv4fcQ+Jndt+zgWnQEIvulLi3kQCye0k
CLSQJGHw77HHcCGeTpcey2RG5pfxjwvtR3mQe4wJhCzVQ8fI6bENNJGTxpavozLX
iZpADPjBcQemFmlFVHvcvn7XcDGPZQT2UoVasqqm9p6Ye7a0yUqXDeiSYpMY/391
CIUSQvCTsjZYCNVny1xu+So/sLCUTr8gw14mpw/dJ4jSpZIvlncx6XVoNuh/zMNq
J5582PWrKoJkVov3snbDheaJJPF9dr5y6UNTTFzjSTC2R7YTW+PDy6ddPVR/9vEo
ExKXbSmJ6K92pqaVa7qqv7KMRrhhwNGyEiUTfu8j8WdCE+GKTASQbpLMC2RnDalf
XrzLPCgpdACuc1JsJla5b4sACruN1+TBNAUf7syhWOTuIkcViU9auT9+v7GJB2D2
MqxA+/7zysiaG+jZSnLN4TwBWQ5KL1XXGXydeVFIUOFJ94k+P2gy8icxRukTeifV
J+vz81Bnvhp9xs/MPItwMNgU2A7d/1wYg9UejWJe6nosYCvZPUjFFh+JiuqCe1Xg
E+wv24QEqD54cRUlKjlQdclKh1I1ZU5CPfsaONfJJae3w5N5Kll8NU+tvYBLWH3b
5hHiuJEbalGDxrhVvfXKbyk0NgGE7afZiITsH6GYpOaimuKYv1i4GAmEa5QtNekD
JYkeCeeZ/X6WTuR05g2NJQ9gb3Bk4TBlTtDdmT7MD753PmmKpcRk/3xj4kHdB57J
syXXQ4hhcslT3g2WVBP58LhmYVvisZ2VytXsI6L22k1U23XiTtQ+iw64FkhfzefE
JblU6rZLN/pj+QY53kL8x7Fbkqj/ZEzB9ouChtF4F1xaEL8pcPU6VgmU6/Hnl0cp
DJSI3AUSI62x0PWSDhqULpZ4L6w6wI18Hu5lYh00O/K/cb948FB9rApPqlcU13ib
swciv+ct95lNMUTNTVhLdtWsle8a+X093xl88gtbGDVke8Z0JTHppmCnmuIVMVyc
YLr6BsdtUG13ltZQuu2ZoOGtjCUWRwnC/o1U0s977pDrNVxgRPLz/+s4/2FqJT8T
yZQOtHqI0g4KPNf+iuGCUjjqr16c80rxlgGOP4wDGCT1QO2phX/Rj3mMcVYAFpdc
RveesL4QVjIka4ViyvDdyWKQLVYnOMHwSS251Bpva7zBcOdh+VjjMnvAb3Iw1c+q
F7H1X2/0mpNsnj0cLrX1sLiKGxDNzruqZUEZoG/1trVi86LIm/IF81XVTbfiOdS4
xXLPtH9PIILNh7nj5MMoL2UU9Rtp20SqwZQPUlB/ESPRcGx7glgxyzZKBDZOAeTu
vlIrYFZ29eltZ8a7KIxkR8Q2V+akd9k69Wt/uLUvhmSDMya4ZqpMozhXYeYtOo8a
ZBVusM4XMFvaMKcm20Av4JnoIXYLs8Cluk3vFhP9spXpibzj/sHK8YefVTKQJ1Ph
naxu5ot4EEDJrJxnxtsljhQtRPCc1aLjMkcyd6NMMofaqaLI0e1fZpSwgBI20Dls
QSFn5y3yfbJd94Klv5AjXI02XmJ6BQDg1z9xsUeFfEHyyS0cQI7tZaI8BdWFMDST
z8HL17emeX/FZLhKgsDFu27Y9tHluIaDVoB3Dm4hxGyIesesv+16RnLBAg58sn6e
T6RI54eANVFTftwSMHzxGM3NmH8f3w1ENYd7MYG54lUxkCa7+MA97Hk/7/1Bkvzd
ESUN4GyW9rMswNzOgFTxwjnofXP1BQd/+rr9cFQnarhwhTRcLMmb1IW3L+yIjCyp
/MTeEUapB4DzmiMrbKZb29sDHsjuy0FNcPSqebZm2KLkPM1qUvKEVhY7iQibwbU7
7gmH6l15zlEZ+q1qjlaapwH/XmJEFije54/5xxssgqlNJryBS5bibKfiWC33l1H1
g4crDoMjBwXOKhHzDBqkLKbd4VjNOn0+aLOX19GsjB+NC35X4gvC5PUBwJjaD11W
YXTN2UlsMyrV9I4oBnoHlH7uXg4hx+FbaEPU0CVnHqKCrfUP0gz7YGK7ZGu6v/AW
eUe5DGVZ+CNPr3guKK2fo85g3L3XXcFBjn0qKTSjddIcwqpCdjRcrchFSJp9gfUA
2Y/j3CWan1yFI0fKqki0Dy/OfvH+/+EdEddu2nHOoREg3Po9CALxm2nBidTh/xyV
+uFXrIec0E0Kedn6Bbt48gnM3AM52erjINUhMn/G75nH9Xu4JP24OzVDbRq01h+8
wdGtg1oFdDAieFm2h9YE6Zc+l6sQQe8KyGTfESCadQDCBppipi02/Lmnxif+Gn9H
C7DPYkQVos8mq1vZmksMV8bd7WF6aH6kUqrNk63nWUnD4OXjmMM+5jIMs5mw7k5L
IdfXnPsHQ9gR+XdajkFZBXFmbnm64aCSTJx2yIY6tMEeYzuyKJc1X1Nj851sykup
Ty0E59D0wfso4PsXqRfH/A==
`protect END_PROTECTED
