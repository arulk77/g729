`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2RtTiaLwZbJSuPbraFO4duGIj6u6kbrSctS3s7j6/1hdjThu4HB6EQfqTBDBBPzd
+AkgbhHU4joXyF9nW5YzkjNkA+8Fzm7OzBHocOUhgtAdejU8/59C+nylnYAdDI0w
V4B7mvT4hQ6xQeLpDLsHJCCR5C+idNXbA6O3GrDkYTtUwg9/6Isdp7ui7x+Ofnvs
`protect END_PROTECTED
