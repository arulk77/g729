`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNxyFtd+oGJVITH6fN+QI3TKfMnNQX0maum7iHwSaEOa
n6yYjesUewiAaowV8nWJdYoLhUCK0ZDzIdCB8hvmrZLLgT1IwaqsngGUOHp8gWS8
P+lv59A28WQZNyDqd77gkjUAVunLfG316OkYPLXlCfqLeztjxmu0zGmOkZh9LXz4
WFVbFKhlp9fldfXol4vQFoSzfWQSumULH6R9fNgf/jhA4PCz5Wu4BBPRNjIUaRE7
5dtDVdN2PxYSS2YgaCKfzGFALsSCh70CGUFG9AB4Njxhws7pPTt8XPAY5aRTU0vz
UHt9XOvwdu88FhcwDajGZwwq+dkhDWQ2us3UW/1NgKMEOTNvEuZNtvV9oQZwYx/Y
uSonZ423LK6ryOAIzxueeI1roGrPcifYjYYFLmJRuTViYEnts8BcPadYLhHG+WrT
aPwhPg0tPvYXGTmYEHaxuPJI9DUnB34yS0vXZOOUOTZVWDO7p6g3SUMoWQauhTbc
P8kd/pKBV8ZICYkjKrEJ553/HyjgT38KidUqKuHPqGpEdlQOJEFx0OzcHYEe3Mz+
`protect END_PROTECTED
