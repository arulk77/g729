`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aYGhvlOKw1kSJFv8yPXnbLjN6RbH2ms6aj8mi79nzrrY
47bMIGmIA2HV/512r13Iuz2azaBTH/14g9MBfj89bDPsujEjs2bRERATqltBuAG1
ovrLqLXuSkGKn0I15CLVDj6py6DDSIRKa3aCacIsW9ZNkJ9EFOp6D4uTz3zd4umy
8zb7IHRWpoOBJW23te/60ENQ2+NaklWib/EIp+yY38KPE5Epky2UX4PDKzVLAAYV
ZzMgnRbUT8uN7gUKrHPbOR7MArsxKwXfQcAHKbiwO5N4uYbEzK/5hhP0NSz9nCQr
rSFs8O0tzqI7tIf16YXdX+/Ei3WkPcFDvt30XjlmPOFAq6t4Nn85cK0hS49poDrO
3XV1fXQk5/GIqru8HmRZJuQ637NIzXNm39N7wzNfBTU2B1qgjAbWLYH2C47fvw9o
um1Rym1ekUDAthtOFzZpAOPXxRJGiAGJUG/mZJ2g5T4AoeVfwVEqiOgLWiHzZB0a
DzaxmkWoFnP4HpLoSuRb5JAAU0mJZFk3xULMyRdrSIkSMtQLI63AgSmhhYQTBbkj
n+WXLuchKFIWQO86Oumg8T7lgluLVccA149qUnbnUvALahW5WxwfpX1z1ujk28Cq
fuOitRxNYHs2vp4WOatgj87gbocFO5Rmbq1s4AHB+/Ja4/NOSfaUS6C3QUDZExwW
qPpeJ9vsIvWInkdtM3Rs9MXaQLTYo3Ae1486jf62lmuxzykQuYeZMdaonSLDl+B1
A6m93mdMl/Q4e62gJkz9959SPuqGiUIOI8mNnUkU+erU1RQqPZ3eyhrFxGLS5VWZ
CxEUQOtLfgVdOmvdok/dVXQ2T37+SNet6OxRb6tNd8O6+UIPNNKOBDzLnvdZfuIW
X3ljxh5PFt0/RrvsI7UL8cYbYbPIQIegJNVALlHTclHb4LF2r1pBCGmSvKAFy7XZ
X7g+1bPbten+BZjUGUA/umRq51GX5EL4sCFi103GG8OYXIbLDyZZ5RMT1niRvjrf
febOb/5/8fqPRIijx/T/EPt/36YdJfYSFSX1ETiLOBu4kWy793S3RaULmLlSFVGx
nphyYgtQv8yrkVT5h+T1CsUO5+H6bDpSIqWO8Z2EmHrsNFQF7v0dbnzEDG7CmqIk
QNpoR3wZ5U7F/L5zBRWiaTwW9eG3WLf62jXavA6fmzzAuPhng7VuFKz2VemO32YH
K1n9N+d7dTxq/YlcJexVmc3+a8NFH9ChKd4yNWeSSFtdom5GwoeOr8bEY8retFq2
j1W45/hzI4UXpap9e99T4eaMcVJ6i68zJAr/vnLZjanXLfUo/5kQxQYr+V91QwUU
ripmTOU8xrERef01gFFvUrwWtbWqABCGXQz8sgKX4O6YniO3kGjdfSqdx9B3+Vu0
tfxhzgjo0yZD5CyLAeRzlF/ghm1Hi8Dn586y+aI6zJMXwaNQuCgNx/uY5QjQNMSK
WxAb7LCuJVAtygLzJCiJHr+iNt+I/eSa44jSNMAcXdQSGI40XASjYE4AdvIW6Wog
EijDA/0OLDNj0jDAOeag8CbXTibQgdp7zzCNMZFmThuuLlUGGN8giD53qPK1J9DT
AP+I9u/kT//1HY73VqmD/05vlQo5M7k3otqynrVMy5M=
`protect END_PROTECTED
