`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+vQXnNdCG9UYAKBuim+cnruXVAhYQSIZEplKr/+1IOA
IvJyuBUH7RN1IBp2j5u6+1TMpZzckG1+n0g1hE0h43P8M5OKHumdkqVgbI23knrw
9DWE4+ix9/JiFZVLKP48bGyAbr404rGYniY5heCcqH9f7l68th3fdt/9i7XLHPs1
0pyH4VJidO9W8gcReAUNnF1QuEnADU4wY1a2NsGIpCw=
`protect END_PROTECTED
