`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Nka6BQRJ4bO5XeNO/cedEKFc4icWNYIj021yQ97Cujaw3+3pJVHrhosZE93DWElL
MxB1h8VsruYiXjfMRqNcXs8r6TDzfXnR9oxsj2OLHm7YdPz39iIPhf0mXcpQ+wlU
9F0HkPAxBas0i7JxhZVZyh0xdr7B68TinJgq4eld1r5SsixWk+7ZUzybXypu8X53
ttd1fIya8OJxAftQA1AzpRXF+tPsIBsEClK2VhIjTXc2uY492vTBjQrpzZwfvR+Z
H/kPe2nF8RyMJrVbFVb9jcOa9Mm0fziS52untW2XNpIMWsl8wHOPnz2mpxrY6juR
wqWt/ckDPiMA9nsLVovzYGNltuW97t5IEL6ruAmYLpJHgecOihkpxhWWf5x8Tb56
SrxsU+IsyIxm01bA5e4Alq3tPCXKGKLyqnfUnE3PdW0i55LVlmQVZ8JHX6ToTj1Y
vgf1Lv/bkgTfO2HvuVW28A==
`protect END_PROTECTED
