`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOZnjWTECZH4anqnVJ/kE3iyw7nYvMm8MOwZKlb9lE/2
pykIRfk7Ldr9jSRcnP6KnXfBQL4oobAWEIqp3SGL9DHEEJc+Q6GGWZyg9UcNYJKz
CsavqtdQkTeWFoglh6bVQUbYO3JWRmc+rt5yhxFT2nuOvUK2KNs8NSOB/nl4jelm
ON/IG3CawlxuDzn9K0NEGX3n15KAfmdZMXjf6ViytyGUmV0iLeu26C1e0GuIoJOZ
ALyKzdOwCy4kuHVoSTsu6clWqpERaJADZyNFw2ROOE1EKWuVYuIiUEOS8MGUc/jZ
fXkb/M7o0HZZ5ssQ/i8PLAYmS9m6g+CFnXxKOoN0Wk4nF6ysNfjTE76d51e9OFd8
xdL6bTo19V1dgnef2eVfhsIhPwsPjh9DwZFBa48L6BrT7+/hQWr/WaN80jvV8k43
HbkF50aBowvX10pY6hhsOgMn49AdDbOc+qFtIhXJjKPuDc+5E17adlwDZge5RqVv
kM9TU+rV0jGFy1dGgX4WC/ClaqX2VCpj5UnqOBxkhshOvHgi6JTwATpFBLz4FOMx
`protect END_PROTECTED
