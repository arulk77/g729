`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1af4QNah1ILfMXn15V2TxccI7+WQe9e3b0sAxpa5Fv47N
B+qGSkzFY3jV9cAbUzBENl7dIrX9cSDejQTL7kyMrmtj5QeKVTSGHfpt65aSKVwF
VBM+ExVklZzSLGn0XKTsBBKJUv/0NIsHZizCcv9LpGebLKuccxokTL9bUZkFPEjr
aEkmmELGGJiB52LPYeSgEM35B6ak+RoeIJnF+juT0N81tdANEx1frRVvD/Uw7kNV
ZTMlisiyFYv5zbG7w8s7G4v+BsApqppSRKEENBpDo75/1cxMAUxdOomE5MagRsJc
oMKKwFYonzqgxa4G35TgZxPtw5ctOmZpJF27X1Z5fPwlEzgb+0F+HrsIY85QRAPZ
t5lox2a75t32OwPVHlqIusVvmWovjttpHErochUZP61m+GY9S2Nk2DMl7U6Xp82/
8/UGZMbtge4bTcVOvBvG9BzYVPnX2hT0F0pzQ7hr42HOCvmtJkRhvyFxwPJPi6MA
LdZ30GvAEKsO083QtOSXmK59proT5QmyYAlGSXAVSYgfNPsYZP57Bsy4kIFNHp0Q
vzLd2auJT422Nysh2nvGg/1em7dRVcq8s1Q/aGC0/wlDqMKhTJjiHTa1HRpqKiC3
l+I17mGOxhcvGtD8JTWGwCDsFyARiLL3KfHk0NXueb5eriLIAgd8+nBokWPj0gnx
kjaeenPndomIEZB0lOS4J2C58V8G/GQkun53CMyuQHXIJ2RY8fB2TlNSKbAeB2Iz
NiGl8lsx9i2WKLyENQUyI9vzdf94E55yss850J4GlARps41HlBJeQr1zyoW0vHap
VWjLGyz2r9U2JmbKcnO3GLaAOTJGuuwqmXylyTr5FlGAzT3bRCBFTucDDVWYdpb/
wJ4hmTgz4tEg9VkM+6lgbrQUDitZiU6s9u5trWkte1J3KYL/LU9Pd0rdIEIOEbGs
KnMsRk2uWcBUM7iulnwowfvDQQ5Uky6wYujfHfnhHXYU6+BiOJvDILTElmwFQIKW
wQjf3fxI4tHF5YAp3xWAgcY+TYKFgRaDe1DyKxFHh7i13jKExU3HbhJtT2dkz8k4
MhM33LCbdFHz3uOdkTcq6j6Toljf6rOMU7iVgBgehMxirZEU42hKUs/Lp1uM5dua
3tSm2NM3VQ630dLD9bEqcTXolZE71ncha50e0YMIikDV45Vp3+ajnWur4M8RgxPI
R7uWKpBH3UA+sNYt3jEyCuTrgBNSwUkfYFeg3gLUxAnGM2h0BVZGNPxPENe/hpTg
53vjQVUcEeldk7ZYU3SNgk08UwT7Jda9cJbzn2AGwNmCWBLUVw3gPNUOCnAeIqyb
mTQW31bQW/rCO2RCwmY8iK/SQ2T0ixSGNGR0ZpRPeHKoTBJLkg1EinxfHEmQHQSp
RWj5oTemrC3tvrNqtMgqQaMjw0Ebuusp6blu/Y9WC3lk3rK79XReRsYoouLUneXZ
5r1CwSg8GyYgeFhZ42UUyOjMpCW/Yn4bUxUc4nX6dHkckva59TFGR03kZF/wQJ7b
rAmUEhU3jOoh2L7bQ1UU9ft6FHpfdSJzTr8zA1CXPs2rWVQMsr6Pod3QPJbOva5o
bsBDh22GANvUEobvj8aiXdgSTnNiUvOyN/blEymsJKtG3zbkAPw2M9Y41OEyggkh
UBqqwGxmatYCbjtlnZswxwBxwyrDRUcP6O9NXf4xcRnNZ/enRos31vliH4OX9NIz
KiPPnscz+4rT3qtf4AKnaSKuTeO2lKTjAO/9T7YVaKRxiYRZeS4RR/IJQ5mrShWQ
unBcPIGt2o4OjoS1v8ZyLwB1RmkXW3G9QPRg4tQ8fiY4wg3IrHAu6YzK7/T03XFk
QrkLspbnDYfu+kbuOwzr50cQHpCr2nLNKm6NHC/+YE68h8s27YICxA3GnunJMLnF
ugQMnnFt9ekBb8YFja4hKf4v6ROAC4gHfB1eV2aMd1rASeeO7uiJUixO7p9nkRlO
fjVKdd8ktiU5r43HK7kytCa51IV/RMK8/smBawx+Vx5v24IhT/Sdxy8grLY5d8c0
hmayhKNrssOAkF2stdVHl7lLQoRtnrSv+WmYwfyKLwizJBzVVJxCBJ9v+taNJ4FU
I22KbiLh+RTzx+L+bL1XSXhGhN8Bb+9udky2stFl/MxjGCA1NE5Povq9Tg9j0egt
9oFFfDR3xYlBFf7V0ileB1vvRHaqT9eVDI3Lq+rSohMpS/psgMhEqPqmbByXKMLM
4tzFt3Ryhs7nMSgjQKE3YZHoyDxk/t1nZereFnPYijEjLzdgqg3GR/sTlUjC9mcK
8oNSYPjy7ejPIB+mv2sQ3NX7BHWpwizIoR8/1FOHuY1XKXAeIuJxm/vkSH1nd06w
tiQUyFDWlaxMV94X+UhIgEl8G3+bUN2xtC3l14fByXUxEuxLQAe+3WS2xV5pio+3
sqPr+sAYDttuxPx8aA05ulkRe/FrLYhhuWPX/4G8+MhwMt/auxbls//lFs9J3aja
YO/g/eqfJOtzr1YWHBjWuwEp9p3QV45zdi/G5a7dPqm2HIeqqLWjHU4aI7GOWBjF
2SOcclvO52KmMcAdS96Lt1XbdMZccurCrA93swxtELf+OgNXJNZYuqAaKsMZhERw
K+f4T9IY0h3zrBnzP0pa5Q3494DLZsdtAU9A72hXQ3TUkjpIM494rjsWUKgUYN8X
/TIW5G+EyGHz2sK/W3UDz/wtnEHeMToGSsGJ0rWN69IT6rONpHPYaFywEGFmwOYD
M+o1ofYVVKlPCP979/g229o0da4ccbkjA5TLOLKCzSs0P2vuSlymJEjwVz3AFK6Q
DW7oKT9LZNFjhmjjGxfWfpo+dicdlbuR66s1aNzZnCth2TRxNfYDt3/zP35EGkdV
UbDVJkROiVXjpIZgfSXVM9rhDFU3Y8JJuHKPZITJ2dRHc89208opcqfajiSu2hAP
p0RWjh3TLCAGVCsbCfA/Zu96R41J4bzHzvXHXaEHuuxgkhEeEt9TvSAMDeyGPmKC
5uetsFSDXVV5/q7JCIyxCwR1uc/l4adF26WdFaMK1Nb38rdbF3T/NJ6B2neiTm2B
5ZEtNoZEnvDxdK8EQ1lB4yEazRimL4aSQq6QV0QCgP2x+WukM6J58wUtWXN8NMPZ
5YrGHk3RirMmmSBbtrzO3Pjj7iIwlhQZfxR8kPnXoM7BN2F1rfiGvHxCemBgp4Iy
TWs8tnCGjNwLmu1rfyUCojOmbvRKz6ukZW8rPiMyvORdv+LNrqcFtiQUSAVvp1Z6
X22qf3W71fVcm/mC8HQfurJH1hc0zxd/Qiy12TXY8PlQIf36t5MonDwg+uRWxxo3
8poIlWp6kQxb3Hs6qDMXdDgxFnQWv8P2c0MDeesjvw0GB5jCZp/b8RkkUo2lr9l1
fuQpWZcaef1BzsLYLJk1lbZWiBKd1Crmemp0x7MbgqBqPNuViF+hgOdwPsFn4r1V
oWZ1fHOKHeYiousXATLS6NeakJ1gtqkLqon6AqinF8LUdnFNiCFX6aEJigT1DWtD
/pg3lP/qdrmDfCKwfRJm9H/EagyJvNlzt0dusTFb4J/Ew/86F7eXdD/jMs46bhE2
kMSpKreKoCTrJLWWcI5/6vu9e8uJu586jJG6kI7qEiTgimfZgXyx3PRU8IzAaq0b
Ny/Vk2nDpO+1WreHL7V0w2xmYflyS492XH+l8gp6ifb7gm4BqcRpiDjDSAnWKUS2
rsdroJbU8ICPy3pzANH7NNwNH5SL9kfbbEUL9hqa2btj5O6O428mUAakav6QVTb/
psHr/qGKaVbF/7xn+F3lpyeuuFKVh6WWZf8wSSLyQvXbohSJ/UUH78Unn4np10X1
L8mHObCsnWH9UYIM5D9EOASUuLTQvzLKTVuXXF6A+v8oPqVx2WfwbKLxKAlD9Myq
j94jODQuxpvWBiHkFCxAO2+nLLhao4dyXbY6boKRlKBz02u6ht02Zxavd1Hh5eUB
p+jZ73PWU567acFBgf6XAnDotQqAE4AMRsuJiujqhqoL8NLjnFgtV8wtIwWwVsOc
OTOvIfNByjd0m2u9SASVKqkEWDhe+kwJOYav6B0zHgC5JMcDJ6bJF6l+h7Fh+Xl7
P2s8eCZu9xMe2jES3urcUT41TwzHRRqQLNLB2IqcmazbV12Qb5VGe7mKCmr6rwD6
E5GOVbuPg1jIGfKFd3pyFZCPSM8WsZcN4CbvEO/1eQYLxBVZ6nGRMTSS4vIbOy7h
5Yi+2y1r4W0end/T7KisIWZ0dgNEiTadg+E3SGoL1N3lTgqa0aNfbRzrFH3W4ESR
F3lEDc3ehfWNNwGos+m753jAVg4OwRyk/5HLiMWsI7yVZLHhMy4XTDx/0J4iuHTF
W0VwvdqH1m/5zBd9AtIrtK+H76Kw32c6qX8lctIXrjcFsOFK9EcZiftiKkqaGRRq
FVtlAdWC0Sjq7dX6+SVL5Xp5UpsA7BiFrCK7fGSmdJHUu6gdRiKiB1Ia3meup51C
/1pzwxtWeBo4wCesZwga6PuKaIVwWl1R4Mi0ET6EyzTFLZAd/KC3rzpOZYxjDg4L
lXEtod+nS0RO/2r+UbrNMWMbJsqQLCeeyO/uouYoPNmQe+JJ11D5kSa1ZFMdM7IH
gcyRrNn+vbEI7IpGM8lJ/sQCEKLatnhQeS+Ji+9Sf6HOHwRxd4EgRvU1VwrvxDWF
kKfjNGgabSTkRbhzV1n02txsQfpKmsC36XIw1mi4l6P5RWwugBBngn39TQm8ozy/
zC6A/tu8GswyBLepHX+nYF8p/mMvTa824OQY90qfp8l/4/2WiENOME4IJAHWP5re
GJT9pDswJP9ZmHDyd152YdbE/gkp6BD0TfaYkwD3w+zAFNJfkplWYmnR9Lq+7AX6
kKquufrLp7UJwaR950Vy/+4hqA4FbFOHDpn/8FN6O/mEI01hPHH1D26zEQQZcAmS
fk228GlWixH0NkRkyYiZvKZkT0M44AdvQLUrdjSfP5Yokao1jHjH63uYlA7Hv/da
ct1bJfy8jGh0U89oIe+YkjMSTZx1XA351AioRJ12+AftHL1Gc8XiGAqXNBNp+i27
lhm1QvWZOYz1pUGRArYQcG+tHq9iadqbe5uYREiBrjYdEw7uBUsQdtxZnkPMt1E+
rzdcRL4+GBMYEe8pO1TwRf9Bsk4aY7Xb+QjH5mfpr4iFeWO/c3mZe0hf4CSL02Pr
54ShDWl0sqQZ2omwFtzuUaFVbzBYGMHB/rlEO/WkiXN1F/5bW2TaqXSJ/RgCFhk/
J5LlJsZijfMzByA5lGEKvK+lIywPdCnA5QA7dgUiRctAwebFdBEyNYTApCnCDxT/
dnvrSA1G9Q2TEBVHx+uiJXq3V/SaR1QGFPNjlgGrGiBo6+4r+ATeg1aoSE8NMNJS
eEXqwWUHVmEddVKj7d4xRiynTWosJj0nm/kJ0LbJ89iYRmMzDEJuqijPIOsCy7Iq
s3vS4waTOMLHpG6bv1LgSDDij7Bp0Kp7aZiLxl4Xe6za8jJ1JLGFqnfnRvsZRkzs
L/+leGP2R/jwK7D9splxBu2r14J9vjriN7uK7j5D3bOmJxOLaBZAeseQdmlOoRD7
pAqbDUgVbZ/e8hFRT5KKrbIInNayhXOUzNWL2mLVZrU0qGhCXQZnOra3hAHo2Ssm
/RXYm2IczcqqmWcNsdC0OL5/62mH/7PlEKenjFHIQcOcDkwCre5OD9PBb0eG/hEP
YwBZrX6bBcn45SHRZxtl1IbSlHUy90VlVTDldnwhXbHuf2G0bC7N2JithQSwzot7
uHWQ7Sxm8vESwevPZy52NOvJSqMwMdUl6S/aTioOh73FIJVN7wzwzNSNpUy2qexp
CA+97kr7akvxgFHGiCYiESQNvj4tGg8A89BIiiixvyVDjQym6qf7Ve2DUP4EQj7K
nPr5//ua1OgGjd9Z5T+gEGHwYCsHlSH4DlvtOQdeMrTldZDuT2MtIS1vzjM4h4/k
QySoAw7AzGMGbZYmNbAKffnnBKwmXw8eRL7PakZfArLn86hz2jTAvHUKMqzDPMDY
TNHSCTEWm1QkM5ewIvnO2rM6SEZdLR7k4iJSt7hPtdzx4l+dnchEEZ2oO15mxHov
WM2sb+W2IjPebnUtaJJUOUrGltHLOO+8SO/3QO8hdGepsO81SU0tZZrDLxSPzw5x
YPT27MTW314deyUQ/M1it/LVFFwZgbusXEC71VKx1yoWiSGrOVfYSamqSgN4EgLk
RjH3p14iUEhMJtaAffXDEhsK92utg80xDGT/2K01lPkah4ZlyVhPGq82aGYmPIEm
U7+UYTIn55zeGAQl9Eh1hHHTTXODANAESz+ewwdFebPZN3BSFghvLu2sQ9CBEhmq
b5uHdur/aLmRAW7b99XqIVFoBpCIQitdxdf2zA/U5Ed6+Yl1hfr30rgMP2t6TCm/
iXlEd02CYA0FGvtwGwOUfLStGhw1Q+3vXe/W9cSOXSJNT0yEouI1BhhgNrm+nj3w
2hu/FOjkIE/SRfUDWwUhWURKBd3aPi3AB58E47D1TvpNJ7Tg1vJAS8gxIsRrJ5Ce
x2rq5akKXAcgt4ZRblfTLoPA4FJ13vGrzj3Sd+Ya53hz71qITD6fZ76nG3jbP3Tq
BPLj+2XtgiWmDZbIHOwlycnTIlgFXn8v2nRJ46aRYlR2m4HRr0KY7JLqBApBUON9
ubpvY9Ev/vWtNafqLfdw9qEeZnm+wVzFQUo2+xcCKIY9FC8jrzeYuMxO+c42n30n
jI6Y1uAnVcfPb3+IrbSZ4uiDM/uLS9Xyhy3ylbeOTD/ufVk6n6EDBQfB6K6blzmf
axPn7I0o/6Npe/hTVWLz0y09YdZmWak76z67RZOCTl5rS8elzQElJj8u3Fa5sGYP
VgBnkekYJSo8605lV/uEisJJbV62NLipxgbIKoIGD9teGIELwMI6BCXSfrdKFe0g
ZXB4dhdY1UNS/u4u2pLY6jiX8eOJ6H5AIZ0Qm2pChTxhhpnXx3mdmIiG/OXakxPA
gCu5vonnwOK1lM8ZfUvrN3F6sxgMxjqNSmDYN2tK9ZWwGAzldByJGqrV220XpGbi
wi7XIyzvf09Sfk26s4n6LKIbOFkwHNPC9TleIHrwfYOiltQQaab96CrcpxXxU2TW
65xLcVhpyuqeaPL8RfN5K4ZqqiQMC5yerHtFydNkqt30RTrzfCNE0/bwDDABmMwY
lZIG+k+1eMy/S+QeQCuVdOuZf8NbDliX2Sm4TocseFbtnFNE7Fp/ETgwqe/epDie
yl0huSh8GUX8G2a7a2maZUrQjUebWX5+UkN5fBKpnKRtiblq/lEO5Yl/tWD58m9O
dlVcOFwwppsDNGp4VqYjcIXa0RGLmHzIw3apOrj7zdb91KvI1rfRJ/6KuoVxOoWd
m2YPV5E2Mi9StnWpeHdIamwjvDeqqQ0Rh4EqpyNHzV0hHlT0KXV6VQv5Lx2vzgQp
0qRVFUpPCvczLtbcdlZ+PbquB820Bf4Se/xMqzdditPN4p/Tq7s7WfhgyN60rM3T
C29lAjvTrxE+AknOcI/Vv9IilJXwTkaw6tOctpcfxp1TyBAakM8HwNraqxH6HUSY
9X3lWpm/eDLR377ZTdoTCQdrAE2zcuAOO1J4K3mpQoGAzt6vSPP8uva5XDhDXnHG
B/UoLeS1MLJYdUh1xe8H9Ofa7wY2pn3Oue6jffnINrGIefyDvLMCPgyzqT//izd6
xp7qwk1ejSGSBZeKs3aVBa+ljTCPWLsfZEBcs/qy9GbEEuY+6iq1hp5tU904hSyE
o6Sa9CF28unHX6zuNnHawEKH5Pjf8AnRD8b7J3YNkMwD6PXuqjhe9ClGgkNKdVYt
BPigrZky3n6dqIP+VjOKQuchrFDw2US6FwHrq0dvF+LG/XXhD7UK8pKeFU23idpT
e0VEdNKIZqiA6AxJtlEvFBA3vVCGnU93WFixhmShGYhH+s6LP8HCWrZsaH2Vnkkk
8JN9S+4ZA0o6Su239FZ+n/cg7b8e99k2DKpMCf09eP4fDdkqRhJ374/BX3qEMK2X
HATKjfQFnY8bgGen1xgKhphiN9E4tXtAfR2LjYUQJ+G0L5qDIKlF0HPePAL/bIw5
2ArF2dqngQ4pEFHeqhmHMOszb24DkL7AyafVXDXvKkhQeFIWD9cebIks1Ub5HYDw
tG6jiuR01PiyK/W8QRhVEGq8sZPbRf7cpeF4IavP35YOzPSJe8x+Onj8l15qqeYR
TLrCYjQESJAm17Sr0lFcHrMVMO/UUxt/iwucejPQ9kAF2Nnfx0IPspGPHjHIg/WJ
PEJ80DjWw0LNMpIWgP1aM53PabqWJvBw0Ue4JnoUeVDgFmqtrf0/E4zVdE6OgQmX
HD6cyq8VORcGJOs/lzp+nxnGqPCjfBkbo8sNugcdlzbu0+z8aP3y7Z7Ni9O7ZVJv
NVh9W6Kyeblr2nNonNT4SxTGiankQskJtWdPu1AqCYROWWXt5s2v+weCSjbOPxhk
cIO8NDw4crAvom5UaHqrEbmPJb7K7FmLsC0AT0AwFcnJf3Ph8nifN5+qXyLLUBPS
ZILbBaDvdolkdKdhgaqIU2lxgxsE4uaE4Wnfq3BqG+xboTFWa/MaDCTRIIqBYlkM
TWr1UY+8+g9r88AwjEgXHE9v7CMijQEcrfUhvsVfbBBiMHxF0HRYwx2aRfDIspLp
vssOawD/2b+jznLILES5GWod3Pr24uUXfaY/0y7+mq8cD3lg5LTFktzgel1BsT0A
SXkNDQI/ShBX7C22dtk2WliB4gp+/3u3A3z+y3PfBDz6z/JsjPb2V1zw2r1vhAJ6
7BH7Qe731Xqblh5xNbBezbENzehrczbYwK7tTi+B8HFpkpGJM62PTF5DTfxQxsmB
atdDJCAPDgQI0bqdKbqGji1uAGWxBNeUdUQEuUwrxYLHMvJITaDYNozvghDSo3VI
o2my8aH+sapKDzE/K0w/MUkf9VHwaDdVZgOaPm6gfcAUuqWbAhgg9LINZVBt1RIc
ThwI6HZL9TAL9LOx2OxpXEMl4nfIN4Um0ed4tRdh3E7cR/vD3UsAq/CoV9KcUWFc
M+AhYEL1FQgq8t7jMnOPjLrNY8jz3uqZpcZY8Tbs9AoVpnPsfBVyZq2t4urCVpAG
YEXF9WsBzqO2OLfFWZEMJs/5Jftk5ltI0F5LWq6tEL+Sxq+TeZ1MArT5YFCyyiaV
KGQZQZ9w2KNCsa58vW1c7Re2yoaLMO+txSpN+mra0Usq1BsQyasqwEL0042rhWyx
+0vBkPuFSttXb/xvEwHytYuiazn3TMU/VTOVYmIb7L2qynKRWzNRxNkHYrl1DuGv
oaBIlIk1cTZgxZBUHbaPskvafzzsA5bZryljtJU8sjMHvvLfJBlZHv6Ec2ttzw7i
2n3uiyS7Ggifu9qgCs4W81AxXzqwPcnODsUjXbxh1BDxT2L1vFEBqac6hw2/WD0X
SJDmxYjk2xguyDcIEjHBilFgCPH29o4cKVLARWnq68ZWYlFgspnVNFy/t3ypflzJ
YUV+nafoMuGE3fF/i7q0lWm+9Wen4xQ6a4JvKXWwvOey+NDjiINv07pts0F+FNp8
obg03k+cTdfuIQ4TCbmnRKHSk5bj/gEKHdcstC75ogxxrdUP5hAMAVRCaiKYKtsk
KMWa+fYQZhS/ZltV1TgK/2sc6hMF6briZ8IUKYD1S/Y4Gslms3bHR0BLUJ6pJY5K
Lk+c38gnTQ6lf+EAAjarF8U0ogXjWo076ubK9y9tn6BN92AXB0A8TtmS4XXEYrTF
z5+gXJ2b4LJQfE8bsh0vKTcWyGwjet+rDphJGEVzMQf1Y4ykFiS/i5riJOOQUCle
Fcezqg0UR2+r9gFyrQKy68v4KvKUGW6Euz9UbLKFbl63MeCPJbNQe+1E7PZ09vvt
yTJHMlGBtrcJEveoFqiV+a9Uy2QOQtIPbyOttv2Z9HGvE9LAQ0sMldVaUWRpPINV
nMNlqvCVDj2OrFI9d5TuAJrJRSXMVBn8R9nomf1ry7vqgjEw1+DoZ5Bc5lRHZzKw
qH+LTlwMw5QYbfynmoU9ilogz/RF1w6dVPYNXFQE9vyZK520BUluEI4lNj0VJIi3
qsG1w/4g6CIDLRdbHS/AQi/qZ7lHXrTrgnaZG30lAc5uuyjWb/IBPtxLuOBt3jW/
Sdt/EY0Ul7fTLcu+bkoaLJ+M5A8twF7y9UUCtncjUFyW2UA6TKpxR3lSfAnoynSw
6skltqWhFjaJGUC8+xTR1I6erDLWD4jree7Fr8yXZ1t4EhAcKjbueEGPFP+PKhZY
CtduX2z+S+MkEQXK1FMHYE0B9EHwCTZm3IpPKpdStmp2M1urVzWdW/xQZTFf5ywA
LAooEOakJPL61jxYPgwzs0boglzENp2M8vMxv4Bj8Md/2Ey91xCj/s9UUloffcsC
pKXTd7J3EAhsZ9S3RTIWk4tJoXWB8ciai+W2WZHbRxatl33YtGMLrxGxSJshi1My
6ftpu1FQYH+pty8BJoawNXpZHC85gm1GZp+CXZVoHLjMB/BSuCAcU0qKlY27Hkcl
C97K82QLZ/s7hX7gYcZ9hAPhQOE/L8v15qH1eG7LcC6NrW2lb9HQb8wNamt8H6zs
z3tm5J41MgGXhOFPQcZ0icruSEnZs17I0KvKuzM17nyj0cIAMZAKu0LQTgV0ROUX
3tJVuN3zon8VAMMnmRVJM+N6qQlIDc5xt0O8B2Y/G1NGTdL31mENOoyz5ORN/3EV
gtcAtWc15669g1aZ23WHIzXm+l2o3YDoSSpOJuoXQOrMXLQusBJAAb+JtmVmlc/+
fA54GvKfK2QoVtduP2oUzjYv4kZ3MdsladrQ0n5pUEoSxPVzHQBOhbOURd3DPM05
w5IMneT+mnDxkCehEezOqMOvmrza9tyGB/doLesYZCT+e5+mGncUcZED2NvX34Q6
+x5HSFLn0PzWbW2+VLugGD0mcCCHTgn0vkcPB8xo1JOgHP4FRZeEWDCXAsLieazH
9SHVDj7BGvFG8curLu37de4XFc6MGoiz0RhNKw2WqEBkxpAixd7DMuFDDSpIU/lB
4i50i9S0tmaZ7rE2tcaRZCpbcBSZF5hVz0Sz7a1uL9Xh3iDAM/q8+W1OpgSy2/C3
0WrOy5S1kUNGC/dh9dmH61Qkqp1YFFoNrhUr73AlVkN4911+xbTqtG+6u+oISvvm
hQ3A3OZcWfNjQs+vDIgqGeDRm+S9iUwYZA+fH8lf219xAZYGbjWfS/6PB/JvOx54
y6NxMIxRI4xQHB9VXQ6Fi6h45wNdqgA4MZ5E5Mw4Q2JLIBCr8X+bmJdnJXJrZiee
F+GepbgBZQ3VBVfZ2wOo/xAl9WLNw0qo2F1tyC90GSDEdbubv3L2hxCJcfzXjLki
tXNHli7+K0zfmwX83RS8KYOxCIHhqeb42AxHh/VLCvBCpH1FbR5Eo2qeRPgUEKsS
hIgxGcIC4fGneh3NgVVYAkSlCy60/qSoA0gYDzfZJSy7i6/JhqxK4oIvqonDQpae
mqmN2dC36iqNixqnnFH/Ih3ttE52mVZ48OMcK4dKQ0sPEHmse0AOAPlpV9rnaSLF
oAChyil3Khuhl9+8a1mfb6fawNjtjcnEkeX97zbeWAEhuVbP0KWg0KdAxNbLTNFW
Tm8RD8qHYdECNHwhrujXojB7Nu1m/4pGTWFMizlfyWGCs4vGY8FHUtZ483TjprRR
EKSlBh6O5iTwkvOzgMc3Ex//OzFmWpcjim70d4vpmG/pHgGnzT5TSiEqzJn6XuY7
q6ZPxbWsKraGtFesVcPiZ2v3EwxzIBfzrfBhaAUvLQK2w4NOkhv5d3uonszrd3HW
npYM70nPusqs8W/J5EojKONuqnmldfQl6biGIq9b8mUqfrAANYA4YZk5u/QKbh6a
tXu8vzupCBxR0n8ItNT9rbVwO7SUrPsvC80Q5dAJQDy0joaGV+iykrVMb7PY7KuN
PIsCjaX/A5tt4Hn+dbDbFeWc8L2TFhkBPt2L8As/vek3SK3ziHh/2fgOTuK//GL+
KPTyulHOrJLZ5EdEdnl63uvg1NbbIA0Is8TFC2Ryi351p1poW1uLPxoo1rA/m8CY
G9RP/dGRlzRANLZrFZxzrUza9+3/ou1v44yOq4NOa8aigXiCfzyA0IqpCsODYUUQ
NKG96ZVUijuD4gdUA/fF2Z8wiaLgrW0GUMf+sV7Fr6lTFJuIZIxokhBtvi5jNhsK
U3NmXahT87/3lpUxEyBRbfNzHwMRgYsbXbQl7YFG7jBuC2z6zK+qJi5VV84LGEkj
ioZw0StBAqdEA4ryKYZUQJMKN1+YBWKdHvn8fGEHk5eTQXQ9pLMqzJxejp6aeAWP
rGwooDJ+B1k3X4LKJ6J24t/G2TXJ+yBvqHLGDgiODdHZyS24YsrDZpsYBs2R8kpL
EuIV27pC3kxdNbZL7vlF8TL2fTyhw94OHb4vapWcyh1RC3GjHlCIKQj2Hh+QEuqa
ITBRzaC9WxOzrIGhz03jD92SR0EBw0SGygCEqEXnPCnYITPZPAwuqdfoG+r47lxq
u9CLkZ67GgYD6hoVF8Cmsu1b6ylKwPTXCJGtzfRm8NsINO7V+iot3oV3n9COa3fc
pbALqf1UozbrTcv/Up6cI/2MqDtB3pfbrkUh6+ldKtb8KmsZhVc4JmNIXGqugN7w
qYliaBYQSH+Ok5mHgrfcfrWEhFPSYpKJ4nYauVBdlAiGR4Gjh4HTMOLqHpt1BX3F
v1ujqA1DnZnMekuDeo3jP0MF9Nuiz8jJxSTN2jvwTXj/jLfsO8SjRz05msEj9bbf
AFeuv4hJl77kCbm7txiuTDaFB2zEvtaK5NGc1Iqgl9HP8C54ctGSR27Y370DRtCO
kL4Aa8Bn0w7Yhf4JIe/7JK6Z6ThtfPhoiQg/Vn3qaaNZis4hZwi2SCsEopEHTk8s
t5ltSVigQv3fVAopncdf+KIQ5yeKj3V54g/HHOyhCGTAo3e5Ttlk2fadjAbXAIfl
GbRJhfdPAA0CBR+59UJhDXITaLWnE53H59Bbr51LDNsVQnXraF13GaKIa2UcTFN0
z7BfNjqBfyQywFlWLTOCLxmyGZ6St6Kvzol9uLp/wkb3zmh3nl0QQwHP+E68LJrm
zo6qfBdqi4/JQRg9AaOhL3vZlLmyRy0jqOz4gtZruaBI1X4jSrRsVNJF4iZtiVsv
CKuPCJ5baoD1ub0xOwMmmeFcRXe88cTDV7k20KayDeoUhQdSNL3UKgEDbkft71h2
/k7i/gegF9/YSpzbknDs8LZ2cvSdIpcNZFM/rlSoneLeyjx5iSnyFtbWsd0VXLpz
AXH6yn6XSCn+9p8ZRtymfkYbU7xTAlclLBJiT1Sk1QmXHHuD/l2J/poiwydVehf9
hwM4bu49NVPZCECDU0qyzlCVTOfXYqhMHP93et96j10Y5VlvwMhJ4vcrrTLLbztt
e3VyUl2QdyDGun2pTHGp957EgOGNlrS6XuEZe7lJUED5nW4YP0fw2v7/8zs1IYFo
cqS8/+g5Bx7HkxXkTuAmKJIc5JwRZLwSiK8K9h4DGD5zYbD0WO03jZXR7ztpPeCI
P2ftzW5UGQs+IVEM8sBlNgjrmtBMYdwQ9HN2E0SWfxdARY60cLODnNAaEMJi4uWd
TFytD30OmYE6IDNVUWR45yzrWM+1L+m1VCJ0nNSpz95BZz3P7MXjZk+M56+wgonT
YOpKW40Tfve/+3/DXsOh93XCqgy6tAiZ5SO7LsQMMvgIx+5poirfZ/ZdqQCg9BXN
WIhbUAQfeO2UBmwtfCFaGTqxudeGhfbaih543KAJiQt4SB9+I/UsvF2+XO72HJeX
k0SAZUzD9e90Hr3MIOHCvAmrnzk6xBfX/sthXFu/t5lYRhN5yM1yiKNOtjRjqXf0
QwxsXVqJwpqXiUQD1SqF64R5qUdIq4yzyneVb0vLgZqoQRzz1oVoCtNoN9uT1Mli
U/kHEg5piQXmSaI+Lvo9LIQ8Klz7aU6ftSw8DjZD5bg963vGpLnNQf071hGZsSpj
yFZFwXShMj968fN5OEwG4vgcz2MjPuoBzTPPKrr7XI92mowh1javH/prz+X8Xgxn
jeH4sbtGfcDffS4EJbx8hQA3K959WXL04PI5Jix3JV1iQpXbeR/ULH8xpjx3ciQD
A3nkQ4Rk9NnczYw7MdvuDT6cpxlntDuKOLYWdPWHoqKGREL6oNnTYmKeXhvq0bLv
l6Dd1ciZ13ScejUi60nw7uqZPtPjIsGaZJ+QUIw22h1OiTHnY9P67OeHEV3teRdC
ud/hdnMpQhxFlhJ7gTA0GoaYT5tuYusvCPSf45356aH7qnC3S8wNIvtPzj41EpVv
qDowIBGjnZfrNO1ifqcitB1DeWSSKZnF/S4DKC+ymEyjxQjLXtxbiWA1mLphT2rp
lLC/mXOnGMGJnBBjaDPziQs71GJaOaT7jmdIr435SDH8PJu4eQM+OZwY59KnFTV5
PqPkN5t0knsHUkVyK0a/cKSsoUmsJ7At4hDq80dt5hDXvijKtFtkIroVLgmIjopa
4pi89MCX7bGfHyFZcKC+XtrxExNcKdwu4Y7mmF3a3yFAEwaRdqFSLOFHHsTvBzev
DbYgqp7B7dIxsVQhTJTxpG5ppenK4mAXi0FnbAHrWM3z1zXMTLRQ2SSNKzwjpIhF
DofBRlxNzMOmGxV0+jyv+LW10W1Esn3UVVBckVBldA85ctqO+hpTDXIkkqsMXV90
hN10JRzinexlMTDL4izVlQyjvoQ05oCigX/HZMUfa1hPzO81MCFY8jd+0PxvC4Tm
pM/t996wlpr6lCXM4+h3eM1kDDo31EVVOwl19bi3iDEKGITN+5Jyk/lYE9aDGldt
Lohy4RfHvRsVDISWHJaofHH6bcOplr8LyI/FHSwOZMqmgIoryzm6SvoL3wKchfG4
7LkvmOk32r2O5fkaiHWKvdiwlFqPwPDFe3vcyk7LNtvaFkzqVoCVQ7AWcZFc6K4M
YD8WwH3JDG1Jl8l2Bd3RffrjxyDUICJGxLFEzftyIWRYLzw2ZIlQx854sO8RTn1m
OCwi3w4vHeRuhwjwSGRDx+uOjRcRC1QAfvHvCO/lUJa/0ITTYiCSDfPzTyvgihba
CntKzjKLq3CMhnxeuciVkSive6DIDMvOEr5l3WoIcnRok2nDJnnzVkLlrsCCfT9S
G9ONQ5HIqtF04/VhKGrtL1PNU4d7eBrMMas59RRUFGwgg815n2ZOMrR3FoxdoimY
LV3zGqnongLADcXk+x6ZRTOSo89GdajJkEB15j19ADZ/dgAgwjJsJJ+v23jjb/fK
478CAhspfdlGFf1AeJOm+IV75wsY8GFmtShF/jAobiUHeXgchxpNKtkW20/0JZHR
1ISMh2g8WOZILuH4l6Ir/wwZqGk+CL0OGHS5bL6DP988OOXyJ762yaU8SwNZ2BBp
7TFY32XnZBZSVPDsKmyO1/RQlmRlGA9EWomARqXlnx2DY0JbRtTeiWsU7O+TrswF
5xdGRwjo8L6uMxQ6d0olabF9/qrJFDbgaRn5/HAI2zcQTk+OigL5b7ue0+tgiWZa
ynMxA2RQj6rie7Gu6YvjqoQFgjEbgY3I8Vp+AqxQ0TIKf5S2JfcrFHDpsPnpU8Sx
g/JpoWgpCneIaHEymh7/BFQokZp62jykQqcEgRJcXUqVJJ4MC3ZmUu8jRWnwqO1u
/2kgWElxvFeewWKapl1I0DlrMT6ah68jIYH60rc3hL/SjYAe/kClpZefvWkf/PjI
AL6qFd16AACGO/rULSgwYuRjLVeBWhoBeXQPDx7B8+SkZMtc5fNjPu4fe/Cjx83D
cpRIk9gy8QF8DhQwmifFTte2+f11p2LMakH7K48gKT0XVNE1jUrWROmLl7qsN6CJ
M8anozok5xdDftzWT+wIQG9W2DGvBiiubW1IRRDN9o5iyVLM8hC1yB97++Km5a6D
IQ5qh5ydChQ59192PDrz1QIs3PNAMDP+8KdJh/3NZ0yUAZry9ADi60tum2PMnc8+
mQzVh9U5/5NBBnrizlPPQo3MrLHPQmbvkaakGR+V69prZM0ac6GCO6au0BGCTtHo
BLSHbdjOXaXfmIFk7pCZLA4dFzNjtddCAzJFVhV4qDoDtefe5hZ+qSycVLAyW7uq
0QNvkJ0NmrGiRroEutmccm0zjoxf+crzcfCIhPfksx6KPB5x832bvfp5Z9/AIzlC
KzYggIXRwh4VWpyTybvMg2ATYWGOr8EYqojnXrfMYbGDEfQLfhmc23mnJyZWQM3f
+r2xdu3ahZw1rR/KgVPmHyFBqJHiKIf6xDmR1YcwOxTicmMdMG3iySwSoQscaM9t
QHpJmASx/gY4AVFg/J9zHjPbNSzS11VwuHjrAoUnhntuvUjYt6/WEaqBK2rVcLNi
iTkDEC+vjxC0f+5MxqyrIht1UtfU6Z8iZgY9DGjq2Cj/onFH9mtL8rrja40zwt6o
gSg83jbiGlcoc3t9CMJxPAKmWrwCKWf7Ypl6DRxOp2jMBcvzQhUHNQv/vWnmSJ8D
hgjajTA7drC13Utiq6qNTLpNwmWItAoMWnBiFEIAsuJAsLfHro2GAfeRWsfbEZne
cw8kwNieCaj6lvGnFyFuo42T4swjbjv9LXwtJfr7GiCWEnkD+UO9phmTppmIOnOG
nZ01+4JAfXwi9jqZHjss84n5Nww80gYV4PGEe19l285DxgLC+Xisb44dnz2BAb/F
W1C8S5AT0+PjAfwm5O1T5/SI5ByBARky793ZjUcEO3uRWTj75cFexxf10+0Mvr1G
cws5b37j8B65bTzzJK58xo52LSYF0ksMBbdOp2dbttR/PUSb8a6vh7GTp6fJdfWs
Ese7MVJ9FwvwDZuvKGyL7cEI86f/Jk5y4WY2E2Y9Hr/gOPa+pFJMeMq7aYG2PMJ3
AW9/uLnfb6hqqkpJlh9nJWGQdg5HVzR6urJvEu2wokb5iZ/3lPpHwlcG5F0fchzb
FjXVoY12TXdocjSRy6zZ0539bS/IpiDIQjA/aSixOt40OQqAfgF8Zf0rqM02IO7g
dzFuHTLLikUyZrT8jgk+oPMnnsJKPRrxjy5tCRZUFJOu/je+7AB0I9N8Zc0COCBh
2qt6DQJ6q6kwpdRf7S+g9h4O/coaqv8UADHF+8WFdbxPdzbI4AtcemxbAdSFfylu
StA7tcBRfq73s3FR8ilGJhTU052huwORDabkMxZAtmDCLkL/k3f8rF22BuTqtH3Z
pEQYNPf2gqfmRNugDg+xJuDUTy+wp25oyoMfGUCDAoDYnOm/CtDV15CGfgK/daR0
BYJKdIKIazj621GQoajAq7kh63HtdmoX+OgLQ9tI49SmuNsYKbUznqqYgH0TdMXs
e3ZW9N3cqh5/DZQDo4eHWb7MMcSZMLOiDHUr8ePB2wtXKrng1cGE7K44vY5cHKxd
WJbTRTj48avGq4qjWFccaW401kpikEN3lkhoXsYIuE0UDNlksq1OR0YveTSOamiP
9p8LpbsAZ3kTAQ3iUx0ziQQR6zlxFp0pqE/FsIwM7nDKphbzGXz79CwcJiPUaM4X
0nbc6+cnnbEFvPvwUbnpg3t5cnwi1feWf9rUzYaD7gZPOLI85HZpPsd20145RSKA
4nWDxUDU2IoSYKVN7e2qNk8mI5fyWYr5t+Pm9GNh7ViWNBOVZBkqTOM3k/9CEt3V
Hn7850pRj5yc7jhlPw/odVwglVhDPZAPO9SNIoezX61+WH0efokwp+7priZJZ8+H
m4FWHYsJm9d7DWruML/y9GPouBFTayFR6z0maNHeVvUbzbIu3um0knvqv0rzS1ay
4ZIaRbrCgvgE49/V6qWvn4S3ggzEfPbXKiS4dRd9VpYOMHdXUa5YUfuZQZc5Wjv9
5vNBFbRaDFokuzuvuYqzFOFclzP4xIeIZVkTUnpAMdzVqXiX0EKU/dSbFFhDazou
0rmBBL5+N5U71kGlmeuf3Z4//fCjzJnqhXvkqW2dEfVjrhCoQnCPCGvCuNi2hH4A
sstuTIj9EvxdQET44IpOa1psIte6IsbWZrQPhcPcLSKBUNimKmNDl+ErEmmizKkO
7SXRttfSJ8K9nGKupDACvdq07T73P0tSpbheOpT4peIHSmhd3FuVpMhLmu2TKEGX
wg6D6HrLJuAjYlDfUDm+RJyR2aKf2gIs1084aW6D6Y2LpebN7yIFHBwaEdAUJwVz
JuH+Bwge/DC6rKad4QzFpXvPrR9t4w2zB0WRSqEXGsl707iCPWn27QsSYOXtwsKU
vFGph/TOwEfagfPEhZ3HAx+X2q9BHUMUUDAezAhNgmr9lDs935RDy7AVs45q3Se2
I9SulKNUNqtQ9mDdLsMEFPymT9yb9Qf01rwyKUycEZy1J+YFIBGnpsY/hG5BH95R
87YgCoeqjkOvlL+TasC8pJ84iTE0w2JPMJemaj4f8WXJ0Bm+ZS1c2Xug6NmZVmLM
QEQ08Y23n2jvI8ZwmyOiiNaZ75Wrk8UUWn12+gwga+Nq6MLRV3E/ApeyVw93yn3R
x9+r1rMuNKu8G+RGpuP2QXVXL01m9znbsW87QwbrD53BJqVqoNgJpoLFFhoFxTmw
okWiCstp/HhDhTNihDHDBvLDBMG0KmNx1dUjj2rXWIRc4XBDw3WwcwHEWl68ObwI
dngyp1ZMx24NRn/HVAQKt4oIMZsvW05+ch1/MXXbe1VPq8c2i/MKHcGXB9C5UPk8
K3z4IEULMs8yRBXQuJJ/G87sEdGg42PGiRZg5BXogjuNrlN0uN7t0f4HoT8FPnhA
Y3lDPMj3QPAx+4jg7+fCvns0QhjJpmeri/5wlpf479Ta2gDK5UtTUQZztMUMHKNg
gNS5+4zd9uRE/IQ2mr0VAGbG2WEb6N9to1nhPFxY9uuPi1JKJYQyvPBeT/IaDd8t
BWzjzit30r0b2GDnNUdwZ/hRdoRc57bThCSNTrzg/vl4nP8Whr2mmLLhlu2rRwSP
LJE8kmDzD7fJGKabAInR+9PFUf/P7v7FFzMykq52JW9G4O3qVerWLk/zSRbzKnGq
V5aYyaJZzVyRtwntixgSU7WHqoij7ye7pOZ3v91Yx7lpeKrOlhXmO8VEbLf67Zhs
0Wd6mfd3e8Y8jXyjeEv0exn4Fd7GPXMDiJ+NzpKYiAisMoNWKaf4ta+zY/rGI5pN
UsDO6PcGbtS/i/q9y8+4/F/Rq8Z+bPDwsK/ao//lWW2Tn6QqThPlnq9if0TGdaoa
tUq5qwLSzNW5Z3RpNBHKqJPFcBgCXlLEzfAhk+uxI2EOfzGcp6MXXcYXDNEVzsS/
0QEQvMttuX2mM12z9k6W33z/xr5oyAlbn6VehI0mamdMaVBHevhbC2kk1torTS+/
smijrwwVyQOnkJxA9ksBCwxxyMT0Woa7+3DwTjveiGNK1PRDtTmNPW53VeVM+kbI
lQLh48qkeI8CRKLXdWB1Mwiae7U8gi1PZXIhC3BtHD5DebjXEsIo+T//wFzRflYE
4M97g2NJpLlLa143axcP7iZO6aMCaUaPcwuhd5XRSuTW0KCYlY7kPDfGBTIVg6Dv
OnT/7mA89JuWaSWBiEK9zHjHCOma+g3YeGcMt86Y7FkKtp74fPkHslyhw89hlEr/
PCxN1Rah3gTiNn1wCO4rDthK6CR1YTz7V118GRa1gO2te7xRPjl9n2PdrnS2Cffj
RSCtHU+qvOuUSmJgFEa4uTKnOeSMbNmO09HtMjRjvw5nMMk1o30JVjIXCmojaqED
ULKCcXVGrM4OatehWNV1sytO0UcTXsek9PFuxXriu0LF/qRNzP0kK1GaJD72NyCB
3Ksn3PVniLCVPdLG8GmDWLHbutTlMVK0AZ+pbSum6L8B0OvXBCTRag54+0Jp0vX7
BlWStO0LQssUkl63YDz6PnQSocAkfhTTeoVBujjhhsUud4bw54gR7CbCwXoKtkAX
jVIZ97k1WBRYDQ2i5+LNCNUIscAoAvsF/l2ZAw2kQfA+Cq3pQSu+7G4/lCH4d4/d
Hrf+5hPBNCvyqW2cLPV6jPTYdOKcuTLYgyWiGyApcsrnWbyH0zzusG7DiEik5l9M
iLc012trmIQd1julCy/Gp/NGboQHhiZh9Cd7yfABosd0X9c8O+hRNGyaYdjB/NQZ
+myyxzIvovBMSuNkh1zGWVgJOrxdsY/9AJksDXopCuAzQ2EuZb8bq9GyQFr4ggTl
Dee637w99TI/9qRf178PDlPavo9KNO+ijGYUnHFnfczhbHnQ5tGtQgykPC6Ct8zl
97ZOdxaiwFBqw/3tWU7AgBN9giHKBSQnoMak99sWq5L8R7d+RinnypSpi5L0DcCp
Gu93G5dOrkh8x3mh/7z1G8UIs8KmPaTef+IuqQjunsYoUe3oW0/Qx/hWUlF6QgH8
fryhyVeAKJhCEDHpz38RmdL7HAY7RVN/D4z3FuahoNkQ8rTjeQS+ChdQeKiLPwji
xe/2iJTxRArPELC1LIVQ6ovFTCFBpq3HEycM1+Tv+DXGqS8IVw7fo2CsWgnlL6Wg
/zKweMRk0RAF9VHlTAy3mIw17g5FDhUlK24r6qxDrWYjPIY4IFoeduG7QGzqnrmf
4vVvQ63hDNA33+9AiwqwMYTF81aEpiBF4hmoYZfH+ntHXxtDgj26yQERhOjfmH1N
rwdQ7Sjp1OmaEv7i6kJcpyY2ztLNOK/lMSHjQm+1l0HYKAEq5mPIXXf9YK6+mW+a
j2otb+6os6/WimiXq7n4fxi5JnHLDInq/tXJ2v9Qt6BL1cw5Vn5pb/+vKFg52hKs
RHKoHNXtt4DGtQ/899PbDFRNyZZ27XK2DIMtR7twWe/8BIcNzUxSFpn5vqT6mE/D
TU8dJICieIq/5vs1RTU6G8nEQjfereMTEVNfwGF8AjUaF/2YNQVbbbxYtfxytuDn
CEBLZsUwWffCVYcg3pymUohGZGnU4JSIBDNxscssL2lkBRREqkbsg4Jh0vNGYl3k
0XjNoz68GBKg7RfzA1f0uMiTK4ukqD4CD0MMA79Z9Dxr0GAB3jRoSY+dldLwL3uN
449d7Di1MKk/XwDgeb5NFRszDjl4czWUDu7Hsl1XI8nRMl7VAF+P92jRKRPX7nWN
HkEi4Ux4fVC+enfGTKLBIjtBdzxb05NqcLfghbEM9mgSdfokRkoRcKwaArzbuNm5
KTix7eTegyJU/Y1pfxbtV8zxyCP/3kLQ/xLW8ef0/mfYtb6aPq3mvUnpHOAx4Wvm
1RezkVrCaREn5p4i/5Ba+InlKhSHPR0Qwgt3Wccgq5jY6gPzb764MHxEzqnPg6q2
0/EmFcmNTr4dxRugUEvIp7K5ZRGA/0YUbigZS8MwfHOgG2UDe0WZYXKJS/+yd9fl
oj7LuTbdr1IVopaUUjQRUul0uOQN4Z3tR8kJ2aD2KMlCFFRtzY2PRZR6IxJVdD5S
UB681DYcEx3Q73ZbqdoqoZhEJLEUwjVpXMLRwHNk5yYY4YQaGZ+i+/ZxPABq0vgU
6Nc+pAVyECY/wVVkC7DGfEqNIP4KEVpSQZz9TXcUQAO5HP8wlEy91m4fsDv9snXj
Mkmn+0Y/jkbFoUHVqLmRPmQVY+8kFIHb4LQ4g0adJ49nQ90v6SSvSC96r7PHMXM3
NQNHhLmWzcLSByN1ODPC22awJYd+Xgafqnj7hJ/HSHrVPqZ1kDCK4UfVu4ESMY+v
Gan/io44X+8S9TR4yg2ZLckhBlrh/cpssCjodw/tMfOuyKqSmH6AIh/TesPWcYuF
w2F3OvqHKpFv00JWG+u67rcq75436nYe/vP3Y8SlfWupBMVxTxD+2TK8WqvByoFG
Tk9Jl6mkMwRCl9jyRVehdwu+J3AfOapgTqKq8wx7kOBhGiR73Vawk4+AlCpI/aRq
bZsB7YREZ0vgYESZWiimyRVP7+9lhpCeOl8kOsggtYY0tqjfjuuYUFh7nxyceL8F
XsP2r+1y0YLLQTJf1kBbo/NKSY6Iru35hRyQDYPwGpI9+8oTho8DPZV5+P2P8LJx
clYdGd+AoI25bpJ/ts6xV+QKjbS65FGMCX4KU4wHMuIWZnxkAeHaj9obptSa0x72
fgHz0gOy8p1rU5sQz8KHSZZjmiJFfueht97HvRvPuIizLfpXycfeO560qX1+AuEi
gHfIQOOZGeSX56zvbZO0/m2zNGcHJVoOiML0VFKnxqjTqNT/jwYviDGoe0T3u9+Z
5V/xuUMSgVU6S6G1DUcXu+nD1AjWa96OyPQzv60P/Efy2LwVLU+ji/wAqPGwfWbH
BWQXkpvv5p+Q6bS5cwWt/eMDmeoggoSUdZMe3CkKHwXaiqwKihsLQ1MnlVQ3iY9D
FhKVoAiVgW2J+7uJSk3C6Fhc2V9oaAmYcTXkC/xSSOzYdGnPMb5cdASd0xbBRMzR
jkJy4sO0LV6aYEviV6yZmxR7didQ464a2OtZa3ISTwdCaEHHp1gGHnKhVi0ADBKk
/LAEGP50+7oPyDFN1blbEWeSaBjrOY/TccKI+POdGZwsJnHnlzO/gxPyFwuPldSk
tTRHtEYcTEh+vYioZcLdoqSDboDedX3+R9WCH9Hb/9DoJKgs6OhJYSznY/Kgazp7
kn9EJC9ymWCISSN54DxtfNzDN1XTJCreEfq4O/C4kzX+irjm1zDG/uJqJrlbQ9tE
urktpUmD/BiC0KakkTp76k7Nr8TiOmMGoVwEgMlyc2R2TiNbgQRcUZwQskfwDqSO
16dSINOa5hNPsrmET+a9WcAmCGIXrxQAY487feVUSU6xL7RNZcQIXtsxCyMM+ac+
Awu4fmynvXYiEchfsWbLVP/8CPS1MhP//PsAGitGncxZPLpFCEMa0jvQrJDg1gxH
G05YNc0kyZgh1lTLSNwaBsbzuxN3iJ4FIV+asiPUEKcLKyZGVjapUXltW9PfMvVi
mX0lfa43lbkgRcmaAGOeeWoDfPuGLFlp4m83b8mmtvmdyqQfMnlFN8xmOs6iti7W
QzOnRRo1xw15NBCQtsC7kgAkc47WwaKc4qifsq23z7j6Tegs+zme92FWA0d1GHAU
URrt2xUk4diKK0//kzVj6W9UR5O7FLiN5tFbjJL/AX/AYqDxOxBLREOW7rpzrReP
GrmYirAO9NJqvcGHjmIN/Cu9lz+ujtwSq1gFoUIHbFihcC88cVCHK38Cgo0XkEv6
3nA5t5jsdiLQHMUqGy8ApVdu59bcLJAFGrumax7jLFzDUw/h7Tq+BOEWAwth5MyK
ULntRZeu+o79o+8kg24GnHGaW4AgRGcFHYzMSM7kiaysLE2IJkYXseIc8BdvMic5
OEARZRa2RzLHiY6CApkfqdu8AvlVK5cXg7Rdet/kqoGsRBDATZU9IAzgeq/sdZbE
Ih0IlFp/2Ku01oeOweHSs1f89Ay4WfU/DVysm3sTuWEskWkRo2HMovtqiYPjRIcM
o6k5L836WTUWoWWeifJBGbMCNZ9oxzhY1z/Zbbsqp3vdi7UJ0W7NspuJ7CAaPBCd
IZTIENxtOaM/yYOAPs+g6wbJ8mQ5j+LPbkCHdEfWi5BK3ywiOycTSQfVeK3Qmpw2
//6qS8zOc6U4PuNrminO++34Hq5zfSfF5MXcCSsAa0Jepu4ASS+ewU0WEb0xjTi0
LmyMsm7trLxpLmLO37VQbFZdapDbTdidNFF74G8o67Wi8chu+0XgiBpD8anay0jT
BTjyttkfHi6we4ZHuts3jXFB8GrxPrf1QSS67rkciA2kw07fuHj1DnVok/Iwxoou
e5lyyJdNdkHysjKab/4ylfkz1OiXc0bxfY7E+p1zwlE3GO9uzzDXY8KHK2UKX6Qo
ks/J5Rzz2Fac8rWdkbk5zgHmU6aIKCV5de1Ozd21q6b3qx8W8NP1gbPJXzCgM4of
MqGOvzkkBm9fuNujdy9t7NAFqf5jV9BEosv9N9GFAcG/NlBgZ5+cXlkqzJ/u0a5z
toXHN+iwz5k8lqzLHpuxyk2VUqM0JrWhyKVsO3WGBJHh0aMmRIbbGnyvkxqkf2KO
CukcMXIBqwisyXc9JXTYaxyekPefbSpo1jcvWehVmtSduh9EeRisbIOgqfJ9prLS
UVXVW/4ftZLAiqJOwSGX+uEyIk4RbhvZVvv/Z9rHhnuVPiBpw7kxwG6B6P8NIDAB
FhcjQmV99z10vjFGBJwuJ2co49dQjLtZPtwWjq1Vc1BQIztHVr6xS+7svXuwY3sF
OIdyBd3b5K7f25wXW+llv8IH7NcUuzKKorVxLjnKsfkonw8G4Epgr/ApXnCjtlu+
z7m/BxBEcsp4stVOgVmQaBAHEr2gLneKjetVG9i7PxV+p69oGh2aI7oTxRUH1Mpj
vYsoD67f6YKdRGalKiNnVK0gm3gtnEmj+5E64NaHghya7Rc96FVI7MOhKYZuukbQ
1FubZB6MFoK6kuOkkGfJJGIfJjSD8o0cpJNRiZyaN8DQF7+5EN6XgzDbaZ3o4jsk
tfTIapDXt+jdCeokPrJ8jsECIQKuKoImbRdylM1ak9IREFdE/RHDcaXfrRiZejkB
0c09ulgw+LhNnzGg5kRCW8+0nLOse1tVGP5luHps210saZImpS0kxArp5HCCnq0r
oSvrdvIvVXWD7lTQ5PbFkF9EhuT/VPeFrScfEMyuSQaIhWN0cHN1cNfgoT+y0ftm
5z63rSxy2F4+hnbpBp88YiCVGhZhUrg5YaDkd+MoSOL4OWvE/QKaNx2CzX4TzjDX
8GW44GY/6/VD+8FfsbOsZ2wKAEnEGxru7Yckyw0nJaPQ9om9w42k/34awrSf5f8J
6YxoMxsjaYHLLUEfxknbiRcMQLFZZsDFpiLBaHT5b1DxTNkrmGbfdLJIw1/FwsCP
v6bqGh3jCw1M9cmlQLKRiPHIWT44MvQu/Y7pzXF/lH4sMalPAsXnXfESH/SZPKQ3
iD/BOU8riGrug2BmAUAqkiQj4jcUPuLUg7t81E+9CKzPiuBcJyswZiBnYifb7KvS
dtDOxJwNElIUKvlv1T7Ol+pOIoekpCGj9VhoiKQWViVT70epytHtetK9o2IrIqm+
qk0Qsu3emHu6XZKdTvcq3Gjt28zdHx+JzFdmqAqiNvf6fj+VwU+gO6+7a9Euz2/e
s0tAtbwZM8Ic3ZQxg6v58r3giJq+4prRHL0PBmqOJaoW8xAQGnuwlB0NREIiyfbh
4XTT/8XlcHHyWMcG9621LO0cj6IFB/Ap7vRX8F8A8hqjZ/NdsQaGh4YEIZasjuF2
ugjxlGA2pw7gLEJxv+8+E3dakXY5iC/2a5a8HGbbHZomj0OoxUswXvVASVZ0UcYF
gH80iqwcffebL7RVt3sCHXahjf/GdCyCyA45wi9tq7AW/VyIGvsw1G+BbKjGJRRT
Z5qJwE5BMzR5KAcLlkvbNEqQNO4VN7YHANV/jFI2hlreGcIAbqOceshlBFHoO/kA
+M9i0MGRZg7vfNba+0LWN66yNjKdI54RNEiz83DppbInB6esHyP/p3ld3bjtm91R
fgM3/kSgKEZMVw7wPlAg++vfxVV+412U6sVY9f7bO7oMsrf5KRi5G5YIntbrJMAN
uXpwcLIRmn1WZGez3TiPj4r4oTBgwGCy09ulIljPX3cFUFZ8qBHeMuVFOjDFk+OX
4/MerEMbFMcqd/2Xc+nikrH86t6fTtkTQffTsUudsLl19r81bzv4gOozDQcmte4v
7ULlnqZFNefQ7NQ6SisYpRAUAXV7r8pax+U7DpZyqWa2deLRzfq45+oHZx3k//8a
jO5RKgRI5uC4/lppXMwsxeHTEqdRyvtCsCyZVmT+FhoSDtY8OmdFG/tD7MIwJFFz
LbsP3heEPEJvCw7N/U3YkgdqCeiJcJc05RoFxCiWDqOnJRgQzZ7PbpT93sMCSyUg
Yj/8Cu9zTZkupc4WEYl78n8a7fZuqnQjkgaFhVXbxB4kAbyLsucoHdB3u9jmL4BK
7FfneRWh+wGHTQlfrsobDqqpfg5EFyu3A9gBn/9m2EtnNx3nQmGFqTR62x6xWaXH
8noRy6/J8/UO9Of3zsMhM1oZ4yDeX24Ji6rAXbhRScluavpzHDwoazsUVDKLZf8p
Tsm8F4cIOYAHB0/kY/6AkxrqmGNfVSPIcHVqC+qHkWtCgOGNJVAB91oCdDRCI9Wn
OY8xgDILVgrZwOhAfI/8SBNXD+3FZ5u5KGjb5KoWeskAMxG9myJaCDf+iHYWKwYv
sQNF6lpIRdJEI7gnkQtfoBnzLn9aqsiaa13BGnycK7Al5hs5BOaoLGxC+ULgLHYV
1Mh0Eete++joct2KbnMAdjj6snEedqTJmlCfdogcJnHBQb8de5SO9spaJalt4FXE
TTIIwS9vfdn0ny15SQLr9kwl1de9rbmsPvjwfVYBNZAMgOne9KNa2NNVbeTmv2GB
e/HyX0DWGd7QZMn2dgsVl1h6BuZcNpshL2HTgNtai4kLkD/lCZJ844IR7amZxruS
Yn9s8EVxxfX72OgXHp0xH9kAwaGZ7Ty5wnpWtQ5vqW+1daaeV3fmxGQRXMAuqgij
Bmz5NGQOP2fQNf26meixCUh8gdGC+5qCcBz1wyU7oWQsqVIYylfRsttJ7d+p8PZ3
5FWNUWZIFOsWridy+REvOJFMe0tR/UhSFQNGuytzNweY4htTxyHtJ4XDPtuOB8OB
wnfpcSVV6Zpx9ptuFTDXwnbtLh2s8k5rwK6/hM6LjthoqpSN0zYjBQaMElO6iLRo
2uPoxJusbjhd4rQBVrTIrQi56wFy25MfyvizTXaoyc4YTrTG5dELfw+O/OEfV/U1
znQ7/YcPL0CnS4TMNM/j9mFzNl5By9/nDNthy1onwHCsxT/VcVkhD4IkKhQyHD78
arwv79Gm7ufmFCo7RTCexfaL3zvcPTcMzJI6vs2c2cY1orMc1tsx9KXUbYlkJL5b
mN84chqXUB14qBnlI86ZOCPXNDSrPLsYJXGs/fhZvMizQvl0FVHWD/onoGB9pbmP
nFC3HtiPHZWJ2tDcz7wEXCd0cETxW2GGUNw54Wl/QqlUHr2nGOBPBRLnLbsPKfAQ
K5bFkIUSa2L4/bD7qhjgylLNwT4FP6M4YR34WBo9qjZ3JO5xSZ3r53UFvCXRWV1h
aM0nNAdjMNigIT41pgvo8bgaBoa4wdUSV2hEVTC745P95upG8Vo5jiTzoMqJ6JyW
KX4cK9dGpOWYK74+EPMvW1vA+HkifnhuAW7dVLicLBraO59eO2MwmoGDpSfOIWVz
W/Xj1+ibVi3n2u2LFi5aKEkWQm5CxIOPdqQQGKI15ZN3o6TxZ5QYSIx1d0kmCvC6
WNG1R3fevJxBdpNaq8YxItVGOj8SWUzeB/MlW021tZo2w0hfSsSzsh+WgxdWqZi9
VWRliOg7jU46y/4pqGhk2ybdZpwF3f2AFxFe+sW++ACu1uwKEiBuwPipBf1rlHQv
T3l5r0bh/u+yksTKcDAPB+hz81jAigVNmNxbeJf95ntgHM2sXVlGedNvS6tJW+NC
2jlHw21TkOhTYL8sWX2KAg7l4SnsrBmHp7kNh8ReL2LwsRxVeles0QsU2+VgmuxE
1Zh3+dt+o+DkHEIoV52rho63XUSBPiFInOTVqwZluKpKFO4Cac+PWSbyy7+kh0Th
H4EMsgUD6rQTPiVPLp7d1U9IIQ8ZdiwPUYPuITzc6byw+k3lFCWD9MFtGUlew5tZ
XNwk8RDC8GqewFKCpqcVNEJuIBKJzyVlAyfecz7rHZSo8dsiKzKHsEnVmLdNeYSD
9OypD0dYuX226VZz+Q5dGPTxjwtJ6gHP8lvsk49Yf7QLxludRqLEsK35M8d6L2Nd
wqXLS6bmCcup4BB1ZBfmRnE5eW5n7k8dQSOWKslL3UX4RESj7GdKfa+f9LHbetdx
lz54yMyPZs457OKL6TODcvZrx37knW/brioZ9avtWWSf4XMKozfSgekj95golBnE
vLrN6MV4Elwws0TqsdV0KA2x3BW8GuiIpeu5cKExzglRU0l/4dU5IbL8C4hYHfLJ
LOnyhIu627ZWV/0IgSA852e8XA21bIl29uFAmE+fTrkL3LMscHD9znzMVmZdzr/s
QgFEuEyQwtLhLwhDQ+b9CfaDsWQrPGjhCiojy8wZ4+Zwo1tSonMZjaQjdMKqZ5Ns
JN0s2vEeTb/qVVj3BcugrJqns6uUIU/KeOa3dCRvvnz+Y/R4NU8bE91qLZ9TEDIC
dlQdHsAFwdFIjG57GAMZGIkUKCk4ZkY6e+c3XpiFETbGPYsfkVJPSDBV4/jy0Px3
Na3nCc4uxGyt7VKncjFBMvVsdPN787I12S0GXjtTGTeXaGEzr9hfzgpwwYq2Y2jt
WQ9YKQLAi4RYW1rUmwV+SQkLM7vbth+GikXihPj5+KdbzHbrt29Xdgy9ZrUWlHZ1
TMem0BrWS0uerUbGAvVJaAeSdRU3oglW+/8DGevghVGdsM/HUHUaC5egkGcwCwEw
Ntmkhb26G10BVOm9H3JKCqe6RULzN8bcx4jAOpI+4V6iHr2dKfKK7qU4SUUMrlbi
60YTBaOe1Ml5smzzOMstGc3TxbAAy6nQ41aVwrApyi7d0MS7HttirFTjvoBw5Nwg
27DB2d33gf0HDz6pWLpfl/PV11h8zctL4CNJiLVqr8CCAp2dKmrS1px7p3jnypQg
Ev3TUyFxdNMk2l1X0TFbXqETvFsnn80vEHVpv7Nr13N5RquCxfdA/MkOM+FLCRvI
i4HOR7ppuMhzPGhbPwKDUK1QAtJk4pB4n2T99YHkusq97Oz0ksKY66HCaN/byjTj
QsflqbinI6NRUWJMqXhKEnbOYX7jiKDhkO2oG0HbPEhxfX4Vw9TktahuN2a0S1c2
VTwaxAJG1KPWPWThAkKVCUcv5Y46inxmFBHwxvNO1WAJHiSSpX0OG4nptBXJYbYW
Bt/AeDznIWI38WNQD9ZCt4dF1i145PgepCsMraeqLbIbql0CaYRQql3yTK8Zn/ie
2i/5fJeNWysE3Z+03R42FaBI5Si0DHtdNW3IHDv00ArDrD+9SNUY278coeYSQlfI
UU8pTQysiCt2F6SqYv2Jx8jirODAzII4HGp3D319GQebr3XPYodCphKt3mFwqJfy
01t+1CS2uEh+97De1v8OHj8B5qRAdPiveA9hZT9aYbw6dFpP1LjgeX3e6VzYBCH3
54P5cueY8visNeTwfXdqRLlD+bpvGecFnAW0gelivjz8pr/39ReXVAmT7ntiFtfD
mn8Mqs2zm5TjFkw1x8UcM3lPMBuhfaF879QeJTLf/R8zz2JC9CB+cR+4B1kxhyW5
DSc5GIIWSBylr9GlI1KhUqClE2XIebB8OUd4GGElFjVtbU0tiFOqCZ75oZHz2Fg/
1Td0enXnAFOpTINUwK/Mc3vYkXI3/naZFcirF5IzW/CrEvZs1B7daN2laupwWP9+
XzjakhtcL18DNTagKhRl/5mE75Trj9/2Ghhrxq8mG0hGjZsIMxk+5BN4SBgs+mrR
4oh3LK04fr7HHcfSwfJrmvhbtg5rYK1ezfpXwIUyJA/STxNvqDxCKdqpy0rF1v8L
/X0A6M30klWuE9G05rOV27Zhgj0tRAfhdgucgTnMVF7zylFug0+MfY3o513JmbZA
R4qA/qej1l+rhwm5jyddp1+7xrukzvZ7AGfhn7ym6Ru4KOgLuyWW3L+zt3t1N0Lw
mwYwtR8N3mBOvYkmaEF41SdpqqGSsGloETLfIlOlnK8yAYC0rf5gDQX8fp5OhWpH
pj28uCLaO40AQkF2N4PQnlv7UvamBXXEza3oZe3z/R4rGzSHVeMD5x4pyxHed2S3
bkMwwhKOKRzyUJd4RdnEJzHmquhA85zmD9M7RasdhEKk+979YqkIu1LtWBoxC9qW
8MFs+1ifk3xt19dsDF9FjBlMM+m19je4CowZHzK2hvyYcQwe31ZqF6ByO6Yj/sCT
vJl4h/6nee6NrqwGNjvU73gnjm45Rc6aPmlIK6EIse8mq0hLm0vQX1ttQd4ghEk1
WB/GsS+Sr0D+FkRD2cDeWoqPuZu0tv7Ue+9SnPFCbBIK/D10zn0lypG4Nm5b+hSM
I3uoeUfBYVgl5etpqohMMBgHX/5uYE7gixmkWFh5cIvuxO2XAO6Ipd5d4fbsZ3TY
B9X/jvVeqg8JZ+H+QID/QoHMsEJq+v/69xvsn+axnHAemIVCtGVclHfYKdp3vbFg
ab1sb8rt7JDdfvgKBjZQ4O0HuvML+em3SpD9JdIaHqkyQnxQBfLKad5tH9XaAE4t
A82A5sLOxazTH/Nc7GwSBg+EFsp0VLQM1wlGl9o6ykYboF9lad6+5NzEZaQgjQCg
dMlMnRQW0vPnYrMxFzav1ey363JyxEmcRGBW39xxbpWOBQiwemIkpt75FjyqJl/m
Qrgwf4I+LIIT1ofVBpZMkFSU4ZoZsCSdaoQZtUXSlSxyMG08kwomXq0a8kusIbNu
xm/LqNYkmIhT2sLOLoN3gQ5FHCnbYB9tAAEVI5yNdqSITYvaA1oEHqG0We+/gR5c
cyqq1Oy7kMggrqPXYd24p+48T+miGTljI79eFaXPg+DoTmeP5GN5C1mKuYSeSfcQ
82FuuFhmm/pq9WyvdeszAmJD92e2jysS2sYV91vPkNaEUUXD/Yd/R8UfwkrWCyz9
ISwpgeitw5oPqstTRTs+yLT4OMXNdPkOSwDIee6BxhZiUDJzl1KM3JIYo7HKZnWl
JFfOcFpXOTvD03zrGfK/Ez+b91Cw3iC7qlUOsH/HRpgoEWSIsvFFEt6EorYAX0Yg
jg4l0mPHD3ADJpfR3W9vRTn84QMRqPz8qN+MXuT5jWJt8i6ep+JkjXjTuhWm7YIw
o0L6BlwjxOXhkqd2Q7reMSSgnzhGBQN7N/OfQOvEM8he9VN13fe0N2ScWFwLiMmo
PtVerzPO2+UTBsSoinNOfypLhqhRat/AWhqOZflfkfadmh/iDjIvDeP2fMbpvTjH
57z4EjgrwaFaRCFuT6KR8NiEUvk+yt7QZas5d1kIqqjrxLoZWQW8WBmNdIDGkg6V
fWWapIsrCsoZctSkQwQn9U0RJ3jBLjV7Rqy2KCo6gKk3DLBel6vCkuhdY8sU5eX/
M0/lPjor6k/dg/jq6oTY2zia8oICRt0DnFGRO6wzGtSnKDkqnlfQUlMIEHDxHTSx
qb4do/+j9cQimgYc4hh29BE4V1QhCuovPfCGBpY0PhWu4Vg2dTuC+xtVXcK6lR1r
shGSHtDHJ/7n5TnxbIlGuVx7XNRf6RoycuSzsqxd/44AhNNvzYvsto0ZOJLu3Ulo
O3Eh/EC26+OWe9BP0mJZ2nkI3paxJ6JyTIlDsQh8RIsWXePFZ0VYA5cjvKfpI726
ti+oEnhLB1MMat81WfUWoIGR/TVpvoqUvUH8O4YggojoVjYs1djSjXKjO0x/Xjqu
9Z2vPWmexffjt4y3FBPN5bQ7T0qqF2P/mKJTYb7AMiHAISTEYf55dtAsTAd5jVH+
wAGlGunAYADqCwp+E47UR9HW+aYRRpOWuiXUdwE579ABfQz/f8FWM3STl9s+7Nim
rqM7QHbPgWicDAgakX2hiyXMpXDBsAyJPQRANcXYYCJBGDpnDGpqJjF0Fg9xfnfj
gJRwl/8+opvgvBckBkJ7WbJgt3f4rtLjPSSm4loJVts1O66QuzFLevG5mCKEuJ6s
jiOd5IUOhKZ6FQupt7h6fc7N23YqAfouTHBUD6Jvz0CJhGRvUcGpgYMxdyrszTjh
rAxiMimRdLpSblghIkGnKrkenioeJ8Jd8upQefgzfI8KKIAQUwe4rih//wyWh5ho
lYt7RBWsbh23H2p8gj9p57l4XX/4AoFIU9HZBNVlPUJb2YV0MrC2cyPt/7pWXzpP
aePbB0BIj1IENJyRhn8qRdufbWi5TPj0QVAsa7y6h/wZB40J30KwpxDk+na9X6bk
Aletda/DjYqj6kXXrVnes69q4j9SFwcF1A8+HedoKq/yqGTdDRcZOkgVUJ+M6m7m
aHN5GD8Af4VElvr4/wHNlKJajtkEY8U8kOwJh4gv+y9vHC++OGx+5rNEzbUdtuLw
QVY5HHtFngeO7RF7OQP+kf+O9HMl4/9XbbqVhrtxCcZxqEfo3zA7VHzRKV/IOFN4
WqsxBn5Tn9XIItKWku0B3LigNNES2t43d0VQcnuT/B1omHRKrsJuUxQWxadH88aj
1i0Ow10hH2J3gTQAPWdCkGBjxuaPVCEsK0f/09ekIIh8cx4/p235Q/OBEctibvjB
ZXsmIHZKBQXybMVGJZO88pI16VhCM3bO8WYfJLKj60ktkkuaxUJsbSI1KTHBGYjg
jHxoBkC3IbrKsJrIUqAJxkSnODnsi3pmD4bEGke3md5UJCeFaC8aj+6IBcDcZBYT
k5CXyi1JQQS0ndb3X/hrRhnCjk5G/Xg3urTjp7gTwq3lVIMFrqIhXY4jALEdyeqc
lnzoLqaXi8he2oLgSS8nQzgI71O3/+SsfMsUoYEXXRnE0OfZia+7Pnj73iEX54oz
3qr3o1OAfCsV86D9FI8bVt6/bF1wI6w5qmhajCun3q/3xG0tgroM4NHZ6sMFng5V
+RRA9JzHAs5tAt/6+IUClbHYrRRLAGSnspQUtWju7P0=
`protect END_PROTECTED
