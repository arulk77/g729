`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN57w0dcHfMIIYE+FZx0/i030KTAUsahPxk/gqn4vQZk
iUuqX0ywfvZnXLx+41J8NQvnZf8Hk4VHtEGQ9+SsXxZX0ORkovQGOWvHcBKtyI0p
YtxmvBv0mrU9omaJnLumvLbUmGFKOTeABl/97KpmuectXwjyh8sr4V+4eFS+7yUI
1wg72z4Ua0EaXUc7x2dJDied7f7U7RwrCpYFgh6KfRetaUvCHJq3EMJARfNrgZr6
`protect END_PROTECTED
