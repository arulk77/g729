`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
0/wt9XZV3slncST9E39Wg+1QYJjHk7q3Tax5L9w9JUvZNYmkGRfMqWO9/IS9x4fo
7/x50lHEzVq5gV45vSZdfCVUdfVRWWpM+DIJO/cQ0bvx91kB8TqCEssBzWC8G6UG
sFOohA2ehK85GjbUCcRo6zJ7sy6U/l5rGXFv1uAyhaxHTJGOR0DLwvCRzxftm5M9
lG90DX4Yoglgn9fFZHSM3MfErlAI9+PS+0vTTb0lSmkR8GUROA8Z5J+v51V1BJbP
Vx0o//qJB4dSeL6vC3fi9gLwOVIMzaQzHoi3xWW/NgMfLUhgAfbED8hJpCnxuIVC
E3koyu4r0KDBkv9dEErp8dzLeojNuD3fqHuGdYwDCj8=
`protect END_PROTECTED
