`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDf5BJeKGhwDUGOYvxw25o8MeNeY/tTCqoERgQLzbcRs
SDDPzp1O/7xpgbtogNkO221nehDHh/kD/U1z7WDQ1oEWtNrPqG6+IWVOE6mABv9r
k7/f7ML3iG50c3ZUGBFdyWTMOOZ2a+zsGl0PTGhQDAFjTv3NyZImrp/aXShX5HIx
1NC/VqLzBHsVIuaRmIsm9vNmdBRzD92gfWqNFJrtWQvVFMWNaPOJ03jFcFahKL40
f4iqHhodhgaQM4N1brOJFuamoN/ks5ZMh2bESyfF2S0Po3tyos0FBiwUsGASi1l8
MTVfGZbPaM0NySLlPqUhuo+Cu/nM799NugCMope5TND40KayiSYQ9R1VC8kD5LNt
Qwa3jJQ7Wfy9NgQ12NTISLNHWosDTW7E8ZJvDNgjkFykttPcpbUVgorY+dlxLMCC
Ql1c4+08ZP2FGjnO51woGgk5CgliSq0YrV55HHWIqIHTU/YLbvs+MRkwdmT5vmOx
no3Bbkyh/kQatPpOa2b7VNpKSSD8pBuzlcNzrPVoM9oGzRbCdCrJIaaN49cYkJqv
GEWIoN9sQg7TbF2Nkce01KLGwq+biV5YG0cRNrxtTY7Vsvbqi/8Ymd/z8JeI29yp
lGYnui16Gk/qZ7y2b5sTGaCMuRpGr6tI0NHk4PAl+OsTZT96Amdm1Yec11SbEsjB
7qFUSZ44ov1GQPBAdYKaxm0HLzL4gaGsrqH8HUKr1vIE8VglqZFuvzMyYvo4TjU3
XutC1Kic9jkEWatrVHsZZwwc8/6xhsZWR8AGB9QICLTvdfmoj0SB+WN4DGZTvcUW
7i85BCHwTwmGAdyw/xqG9eSfCX+YC50/bgBYl+KQgrfjmwoevrQHFhFdX3z8NEKa
dXOXIVK41t1ZHI6RxUDH5Mtu1uy6n/nbIc5FSy4oSAk8aXfOOXCxAjfHS5+g6yx0
OtktKK2un1uSIDCtacXRVFVQTsK6gObaUyCZ7474Z9o=
`protect END_PROTECTED
