`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
5pma+bz2bg49bGmqIUtTLQPh6lcMqW1xSNfwV0nK2N6n3C9/Ji0Gs838f5a3Rh8o
wbJqMZlLEynzXoCO4mzzDhv/MFmwzwWucXipNu3Is/lLwZeuBDxLgL0ilDntOpSa
ajbMHFwfmqmc72KiHIdp9apvKrHE/FXbbmrT6fQk83pZt0FRgpiXEkp9LoruvtQi
WeqtigQt/vxWOfOjK3M5PbJ/L2/4rrssHJRGGD3+miE3DA4/ICYEqCeuVGmhJtOP
teD8D6WWTWMMzqw+qWvX3huJzWE4gjMxUvzsMJNFkn/asuAPOjO/Z9VpstKTPzV1
TxUc9sN9i+XXdkC/iYs/2WmEQLFL0wAJlJ4kuR08vgQ=
`protect END_PROTECTED
