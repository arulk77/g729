`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMwaUXuuGuTkekr312o7GzsFQk8OG8iOkl9m1vbVrUR1
Cz5FXfjCWvN6FXzh10MjxH2BOB/QFVNCKMv7Cwtee4pGsm0Hr+u8XQSMTq+P5MKs
dI7XMTaLc2fiL6PDNvMvIKvdavNsVRiyJtZt3rbyIp6A5QwoG4IUIw3D2ecnImFW
YpStV8zHqG7StmJq/tZ2ZbRUC/VyDdAbtkO0RM2pTfC/Y1hKA3DJfU7CUPNVBNGp
IX6R+DBqMLMTDrE8JyRB+xw0S+zF0UpIxs/DKhF1wNg/FiH/HpsaOYzfEH/3Rd53
4xoGcNnODiZ5yKcLi91GbQKDQWlZ+Ns8MGosjxTkE8qvQAAo0VmvAopIWHJOgY8Z
`protect END_PROTECTED
