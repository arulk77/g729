`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aTk8gok+oiWQuw4QCf378lwn4+YMbOeaLj5pM1eB6xca
GxtnKImKqpQna73yh3PY3Eowl36VEo+OZ0g1BE4kcR1/j4/f4adMPe4rh1U+wPmQ
9sycbKff8JpqAFgwD1GEX1vyowYwqa515TvMg/QrMxgm7HZHVkEcOoBmYBbkx1eY
O8tqQbppSUY38DhV347zUfAj/vGqKUqdtR7l6JHEtG6BeVmFwoDMgXE8MeSEZ6es
eGxyu2T0vQvLRM+iKbtM6XVvqXx+vCcZZijF+kSl1AfCO1mwYBQyxx1HSFrHP5mP
`protect END_PROTECTED
