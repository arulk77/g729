`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMPuS4Hb5AUcWnaUbGqy/u/MT+ixcaTpXzX+dxsjENtz
egOcepIgyBQmrexI4WwQiQ/TCGz8ILZB4UlG7Dj05J5n8IsoRTBg1hOHO7Zbz/nJ
uixvAZEbPrfpQHEeDq7a8fiBjwjRGuo5yvZKFi1IkUQr25z3jZHyBKrMD7rAMhsk
VAHqDoSTbGU6NRQ29OPEnK9M7lg5AF5p06JzjbY4mONxmSbbQXJ1YmTrgIMsTOCS
iO6KhNDXKU0WwRgvxlqRb3s4n5AuIOXvzWKC+oVxUExB0SZHB16zA8DuK7Gd9FtU
l9KQbxrueKm17kCMtak7PC3kavy7B+Gix8sxdSsX31mR+aps9qfjBvi3DAIlqb/6
ze9AtAsC25V56m3Yvb9d6ra2f0A4km5djsZXMozltqTvJUxBiABNCEiVl+uoRcph
cw6HN7h+Pk8pyF8r716pkpCHU5LjRCrbCJE2jydsGSg=
`protect END_PROTECTED
