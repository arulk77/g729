`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCAuPMGsOY0setvMDCZvRUVIwqtyHlTKS4ddaOMegyVi
XniulSIBCIpibMRwqFWC1MkIsYsPpJ5br+XOwLOw7goodkk8ynX1zInA3kFt4OK7
5pjEzEQK2gRIaQdiuiROc0g+zGd07fdUwV3iIMq1a5x845Mg09jUz2O9zUOrqXdW
j5yvxp/D9YbvzZ1osgsj1MIGgzxvm8t8Q5RXmzE+WOKpZH2JR/OnVxmV/6OZs25r
q8bC+mth0NXR6Aq0Dv9rVP1Pdir3O9SRNvDWinJkbwEFDfQy/GCyRt/E8pQdpgQj
GiQ8RKU++4uTX5m6KtpoZUVl5n7saW0WZihLRHbDaFWeDYTE5/6Z+QtzHV5dxi4A
OmnK8IwEEA6YkBFkz8w662vBR3MZRmpWyL9RTsNwyehKl/AHQ+p8rwfD4cSuyrQC
4y/117e1y9ZDvKJ4QBxV+x5iPzHFkvJrewJOX3CcBC6cJjZ6oekyEBsFDpMes/cN
3E9jbpo7uFg6nyAl2vdSBdUPViSsh45pCUsL1sQtf/E1/3dtSOL/ML1SrCi7PT7S
`protect END_PROTECTED
