`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLQj9VfFYcCH8RQuAzPlH56ZPz7DSHT499TgZuIdvLSV
NmV/S2wIkAx0HZcLQXDzz5RxOGVEjWjmCdBx3IBn3o2OvsdR6fVpvLP77/MwFhMq
rnGbHDiiav6oAO0Ke4FKaljEm6oD/dUJR0c23BHK1aBlV3zDuiyV57n6d2aVIaNU
j1dPNoJ/D3z4nxDHO+TrM4Kryl3qzyZVYZ2GT/OxiGZigxA9W9bBeAHmqfzvKAMh
1+tFVGLQ2ayS7u4B4MPEoWc0sYS55xJQqmNkN7klbvudHprZES1pEURY7nKTqwEB
QFzT7GTAYTKgbvMTQsXrdi1FwEp7lhiu/nlqsN9StIgS2s0PYqQ1uM1JARREufv/
59mx4thijxIWI+Tx8CF2Gw==
`protect END_PROTECTED
