`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMXz8C1TEYjznI0NxlojsIMDbPQuMTng0ZOhI1kOHD5C
40on7UY3nK9Y3IUUlBO/7sh2uZ6C2VUvxCDv/lECtBcUcCXr3FgMQLLlpAknwAeH
U71D5fBPi0W/hswXDbrYzgr0TnkNAyBp4zSAVfXpsvfI+58tk8uB0Yxd+jw9XI0X
FPeHGH9w1EWLNxWSTDt5/F9jmEB/uJdn9SPiOgbBwiKBH7yMNzg/LdA/tYmaUkzQ
V9ILoqiF9e6i3DXjoCh8VL0+FS2A2h+rXJM09TInU2kDKT2YQi7WQMdy6FC6OvRs
`protect END_PROTECTED
