`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
YTi9sNlfgsGXHgp29xERje+QqEkJQmQsVygmDPAI1emReZC5ZQQAHVETj7SghgEH
87bAv3FCmH8skWTjfn4qOmuWzysxL94teK6qV9upLP9L+79V6lKXo6yXBHpLJdYV
`protect END_PROTECTED
