`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveECeYYH+fQg3utlRz25u2QQ3T8N/StqOPtkOSzupCEHR
09nY+ZSjcbBHBzalWRQK8NoCLe2p8ayw6SaPG6y8WiNjhNmSmUU9JDE+zjpQ9N1M
jHfbOF+/tn9sxqJaBTb8y4ch1AP8SdquQegZPasSntib1ln4khZBIgIB1q97P8/2
VpfIPiNHyOe+EeS93uPtd8vPnAN12CNumAJ8ed/OXEXjTzuNng9aek16t8/5m9CB
OXkfe5HSXEE9w7Fgelksihs1+Ui6W9KRayui+Xq24J/E6mV65U6gIssK3n1lmpis
QcLMJvuQmrIy4MRvFnFua5WbLwjgCJoa5m7vBUR8QD4s8SkD2ydQmnxX+eAwfcid
50bDrleCzAodsXZ9PiYy/sGRIS7x+hGYCJFDf6lbjs7cj2diKEjudjOtsDGp0JxU
jFdIb5uzwxgGu1cRBXDhQToHU5MD2ZdKHvT44cwGLmQUtAYd/76ot8DjtPcF//9g
/4aHEN31CXpP9QWRXXVF0KanG37MG3gVfOSVDsOW/UlyDuKAHkj7OdeQuf7Clu7g
/CixDCfRoGcp9/0Le9b0xnmHlm3kIY27ufNTHQIw5ktTsrfIBODPdMo4n3ww3v9S
sW09XghB1KA8VSZS66RyijZcqkWAR9xLhPmTJ2g2VXBq5eoKmAAFG5qbGwPGCuoQ
JN/WWFzercHTxd0gjDCXShnW8DNy5UdLmT92fjvvB3tMRX7DUIiUlaUCl+2qrvVN
/4lcynOJCGz5Ll1hTyYVfKLFcr72QLY0e+cp70HDbKHYW5YAIyBZ0JlXhUYtX7bu
8gu+83SFSQuBQMkZz+6gQcjywx9rN5gI/lkKVBdQyzeemlzJW+zXtStw2MgQm3K7
`protect END_PROTECTED
