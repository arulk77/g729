`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveA+rOntjU0vMJwWTXowxasJHS+E3fu3JRSFRBG5rHQ1r
sVjsfThTlOKMQAdola0Yn8tXMCdfJoVo8KB6SCKSJMgYuzlalhFVPOmHy3JepMrc
tw2KfGgqMHBDR+keSF6pzAYwYK52Zq/h4DWSxj7akiWTZsoiRYp8w8JRorZoLgOO
xjAN+yPXids4TnZD/HB7v4jk69XKOxvE0zsdQJEYZ6NpzG/weA4H6eFfeopcYV07
8LY9HdB6JoPVFIGn7m0JgTJcsN/5dNcthpzDJMv3WnT5IJY746id+LIdDwgXBsQ1
tyig01pSTJcuXANEgIPUiiQBWtO57KzJFN+iPgEdaKtA4KN3eaJorJkMP01HhVPD
`protect END_PROTECTED
