`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
6O9xi18RbEGdoLkYYK6xs/DBlTtUA/A0CPcUOX7BBowlahE26hGjVzf+YQ/0PSil
UjTKOMoW7M4032dhuli5aEB4orX4Pk9U9og3aGPQ/j6ps6tNsTVHVrl7zHx9P7vz
T9coCK5wAGpCHKA3LTogxRwjIVwBzAtlxKRSKJ+PnBaDcV5hzXvCCLXJRUfy+p7+
7YLDeuqUvnKvRp4j6CnjPz31tuaXteWr22JR7ur5S4o=
`protect END_PROTECTED
