`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yVYUhYPevGFTtCJvV+s1YnhA7sFLBHiUaK+otWK2Bwa
0scg1OhDhYPfNWumgT3cIiqVV8HY/6EvOVAtcFYAqhLKj6PUi4Jf+l1/hG5Vu+XZ
GYGtH2LwXQ4xMl8FA6NT1Hf9jevCITVS0L5TU647DlHUCC5GOAJnZmQCzO/Z/N+R
l1881SObvqiR+SY31ozU5GJfszTevt1CQDr9hT7CbIGG4EMKE0T6fUIuCHZVArzT
2ko/6zFMCQh+RKq3oLGX/67makiT7qJpkrLPB/GuzTzY8/djwsqJ4FlIRdW9GvK6
Vt2kFNg8cDRsfPAjSDdBMqCRzj9noJi7LMEKW3mYz4ya1zJWI6Dib4HDi0fdSQ3t
6bwhTPhIqsSqEv983iP/sQ==
`protect END_PROTECTED
