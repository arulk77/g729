`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveABvqdOE25xtwdZXwnd1y/eUg2Y7HtjJgC1LytfcwaMW
vQKPUtRR8DEAe8ezp9q5Q4qk006OVKE624hUCHP3KCH2qHjV/+NO5S5BYFGXV4FZ
4e4aqg3HjO6x5JXETMDFwIBbYEV2uvCgS/Vk0+Md3CyrFDom38dw50XR/vj7oM1k
Xcvyy3pN+NnwG1ebwlNoPFtvjgIjoMODwS1FAdYmRowNh1hNM4zIgSq0HeFld3P1
6pjTzuv87Nft2YnRoKG7uKhuv7xT6xk3n37/CGLkKW5cBw9gLO1wY+ysn+WIGEt3
3SWfLwy4Uc/mgLwtDfIIKvdvIY/RkgQ4x3YYgCh2k9hPT6WRgPpERxUHR3wiV15I
`protect END_PROTECTED
