`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKL+J0PSvi9d0mOHhUf183abpHuZ8uSFoVyGbmHhday+
UkWM6t7vNjdF6OynVmm8wd8bYqgQ/TIfuwFLVp9Fis3LvR6zMlCPb6aVr7ErkGpH
GwtM/4/lYiJxdC3g3Q7PB/DRuXqXt8ReI0XAd28TYmdeiKsjhpCrU8CH70E5fT6b
xi67Pnq2GChacKPfyO55o8YtJFvnwEbZniPY6LPPpkoY2mQZkc3OZ5AmQ1VhZOCg
NyzpIZZMQSOg9C16gD34Jw==
`protect END_PROTECTED
