`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1abndi9g79EzsLa6odcThvxNKlmD1oXVhTKsfWTTi5qkh
DpxHEJME2h0B8hKNElW61rtFShjuB0GqQB9+rMdOf/mT+Hhu2YtkkDiFBuSnwHCk
flAtxQ0qGwrLxd7o7WIIQONJ5+Lhk9CMDQgHwMce2pKpda3s45C3nVlsEvJPG/ij
CPi8A21S3h1keZXWLj6R02WuS4ipHY8zbfQPd95gkmnciYrbRKWasFH5ziBxYAaf
4GkAQTtiYNb9UyKjOau3OE035dkQlIaGpbfNAUrbQSiLQsgALgPKsBbrFQ6LaSpd
bpa+KUSgb2yvbRpQYvQgwZUnTU864KXCNM3vK0GvXDW36auITta6NvNK0AJ3QTRQ
Z31sFRvz8Ol29Xc2vEZmzvCnPigBRSjVUheUJnNFGAFabbowbcfUFMEPxd8a+/9/
ziJvixAwDPNzxAXJKce1crPuEJ846PTmTQs4la6Mzj9cl1b1c2shPW8WsHsgqtpp
9NvxXOkXz5w8uuvf4jdatdkHlqc2b/YpWP8WS+nEQGFyL19bSj1MbtAiiA2XLnUd
5UETh4TA5Nb1Zh1UNDo5/XN1B6+PrRMHqumDcVSk4kfxNXPTrwFu0HG5zCZAwJ8Y
II8yR7GebXPaXg17cnJ9ghfjwW3A0GK2kh1PTsjBSk70huhVAV4ITHuw/IW+nGrt
FgaKAnQU3OMhODUwA6uI1SmMTx6kJ8uQaI4dmVa5Uc+UHKmwtgmn6afr12zEZOwk
WiF0RWglEawihYA1zkFI53qDF9YwILyRKYUjekzyc9ls2JiXySRyeML6CIZILMDz
PhW76Cny900O18pfCNAQqwS3uu6us1aKHu4sQrbgt3Ss/9/zwNCrmtskr3ZeYhcf
X8JDmiXI91t0zzIq0B9iQUzu4cX3O/a9D77rzsyZDjmbcxeRkK6orjO77D/0aqJY
9Nm+XfL6U6LPl1ojC0E0vexkM50WPuXrQNmh851KVYXM8WEjc/l1SCWtvQhZ7DPE
z5qzTtJuM/KDlfexeze3FowC+dxpXVGW5XEWIVTRKHXD+0+6pk50h0DSIHSaWkA9
dhe8Rc5qDG1qio1RfnIgLtinsBEXLmmBRq+YGE3e5mAC6Jw6p2FzAMGlaUId2zgV
lwekczcCvuIJy7pbAA+jBg12JELMfi3VQXcP7ttJZjsu53ZWM7i7sMOn0Gxnhx3M
uqsF5eVB/p55PR4K6GEQE/FMa35oN9Ca47/2eQhHscVY298YebTq9TvtnunrQlbP
YzB1wa3ZJbz2iHUIl4QGQHaE/aAdl23d2/miBChv4A/6KM9monm6C+qTI/oJV+vX
F9fUTeT4gmNy+gMDSLfEnG0JNfyJ+b137wL2Q9InyIrp2EQrTEgnuyBw3Nytvd7K
FR2/4QKARpU9yDA/lAvEKx8o5yUVZVQQhr0QKNX57/87xKnBkiSg7lSmgmYH0D+T
q8VuvdEsBbnwVELucAe2iwxry1V3KP8+tH5MErMPsU2VVA5zKvdj1Hfi2ciMXAjM
1K6Sp8/022RzSV0sMr+s0pENCDFVh52lxuZ/KuuyLRJ5JT6Z5sYsHVnzOF46OPj2
6j5hEJEjalaxDVRDVxV4gVK0RD3hstMU3DHq8JLLE4ezCyR6RjEWkPVCZxDVbtjX
w+BEKVXUfNfnqKY8WWEx9IGpS+09aJWqRLaKQNXlkxfqsCVwJy9B089Iq7zJyR1n
k5MMLj2K08B2qYv62x+r4eIzZYH5V3+Cboe79/bIU8v6NSKLSh+vfn7P2ikixgPI
3JAKNvYjn7FKXosrQNFmGsVw4tEtfG4y6oy39xdE6ALJPDpj6GW0XfoJtkwNwGQf
Dve3BlzHUzSf4/akUykFa3W6IDilWdkSWvGUGJ0M/5W49RaDW1BqSdnhsLqItCS1
+xpdQW6KBYkZ8oNY+RONIvScucAZC/Hm3wWHk8Ko5kAodafrLo7jtPj1WAQsuYHx
xegulozpfMWSHusLFPW1QfYIDJzc+6e/McfMGKyjz8webakNXjCNi4JiY1uiQ6b9
TXntgBCP4D30mCprygajx1eVfzWIZoULMf+UOlHmTrpJjq3lbXF3VyALqIbBbWFt
j8nEUD0W5+O7pPd3Wq2LrECJwC87fyAjghMpw6zrkX4yBT9QnwsfV1CN7e8a3aSG
ZghzDIInRpr5ODcaQ6oEZUZuG8o6pbK5Ng4G6yD5/8wn8ti57sDLW9gSoGX56lgr
VelY2TdznTUTQtH8AGHI+QcLHIwncJl2uStgA25o0n5UOAVLYf3A5ghJapvak9HQ
/iVREw994ndr6DiKdxGL5KQPFZvU8I5ayzSPJrMI/oMX4QTToFwCWUdXgbEm6Ej+
DPvTyyC50chCovBVTvTLSfzBZitSJSiXeSZwS1/mdFYp1MxMezFRT/1gLo3VaWvF
EZYw5V1LUsflrBVh+8WO6QWmbJ/gzUnZgQkGbKn+3AZwV5ZiQNTsYmlmcwyGg70c
QxNTixe80jSt6fLaj5zCZdK1iD+8ZiX2+uJtJhbN4griKMQB1SWfxilWgtiYMuIG
nG3CWg/iia3h2u1A0hjOd0+xznNPDOJEupqxJy+HzLsNRl67M3yQ9S49GjR+npFH
un+8958CvCvXhzxyfIi08RCIPi1jdSF4rDW6+dc294JLJhCrwnsI/B54g8uPpUky
GLLiqgfR5juzLcYQP2Irzu4D5ey970IZAcm6TVLF0JPMCQjKcNk0cMGXUUPkBpDw
n5YVutPEHdXw1agTuormRwbIuDNgjJmVKato31uRvboOqCP7EwF+xEt19JgRaIwH
IHb0zCKhGBrRenUgvWcCgkG0mnGhwB9NzZzjW281u1unlWRGZSAuTDKO8o3xBKPC
acPM8BBP0JoyZoIkgY4HnV+JDAEZ742Zfa/7Hm5SYBCQFBV1IHeP6D+yUL3uoAc7
4jB0fOTB/J/xlEzIUahaJ72EXOBJdykiXOZlRaJ8B5aiSaPThgn/HKWqXHF5i6wl
MxkkOZpMHHxkR4+8fhcb7bACcA9oWemb3BxraHb8AxHlg1nBKsOQi0Ve+Uic5TZH
z5mqEMrUwgnOGUW4W/H92Re+BrPHRET4Hp+6ndZU3erVgskJ4IlkQBGt7rMSe8IL
iklOsWw+QutF2n751Hm83w8KAXCIDh48Qtj8Vw26fyBR3utiweOQeMjn41ULcVen
sjgp7VBnpgicNKX3AydXG/5nJs4enZqyR9YWLKY7YjCfwiqGLkXYqfZrMDI41ndQ
AvN9vq/irU0pVisgRaQYfyDJSnamk/Jxtu3RqLH0F4su68KX6WPtNQ4kxJTYeNgi
/Qm+daG6gOq5GnUq7rXhYR0Kr3d7mUDL8rJ5/2s1avLk9rUsG4SXpRByxBhbNBNP
epAo4iVI/0Hh5plaZez7fEoP8w/dlZqHy3jIlg0IKeG2WcmRRvxFxDyV4vTx4h9o
g1leFkUmxQDnvNCgZMSzewLv3/fJ3iSD152RaKgZMru+x0qlGpVg6a1eCKIVZJbZ
Bu904yD8tZ2prC+3NaM1wWczwZfwruWH3j97hJn8MjjpXTJ9CbRX/ATeZW4N77yW
qhsy3w3if4mYooA/v/4B2AtqhX1sqMISDEqlDbn7tdfrZyltivCcMU92jgUa8W9o
t/7XyxLcDt/k/xPJZPwRPVuhT9oysEXtj83/rhnfFSPSE8w/0XdsJ2JcMNjcqC6K
pCLL2k3Zk/j26ZDNpWRNSFHS0GAoaZOJ4JGnBU11vtW4VWl6drzpoTJqlt9LzFj5
QRe/zX8PCc/R5KqOkkuxVbhbTYjglhUbCrIJCWc5C2cYnwu34UNOpmPM2AWG8TuO
cne9lVUIEm9fEUXvMk1T4jHM2h71BSU9y21cY6+CVSJiShIWvbKgaGeAyBlhmpUP
h1vqXY+yoDCHFLj8KqETi+jpjO5ZKdNMc1EpenncE/5mNhj0okHAmSCGXhHAcu4Z
+ZmiOUY05oHZLKEnPR2MeB25K3345iNDUHVGtjGNa+PZ5YJWmBBGPz6Oz7d/2U2G
Npr7V/zTpeU65vAlyQCEqCb98ozI+SYfrDp0utmhpQAvhFeAqKTARzi9izUau7qw
ZNqUTLAWX/k4hhJaQknufzDDS3UqhB7Ja89fPruio6tBhzfXijuFGfiKPRDhExRR
VBkkpEzAyrgqjDIYv0LxQbMXxiylS3Ylw14739RF/Fp1HyQIAuz3+h5oeHQahKWu
THfWArC52Ppk8+U12hVmpACZfeGtipATrColuGCX6fabSOe4mQq4JM/BrlnDAG07
BHu5XuUY4MHavymR3p0iDO5s2S/TmZlZhYS7vfmViAF1hdiQREMyZByIgaPn37sP
IHdhFTbNsxjFVwjlD+HIW0qQbOLSka/ElwK7GCkNDhlqqClKKCj3oJ5IFhhDWr/Z
oNWwFnh0DgmHrRhTz3U35QFGhKSQbvNX6/HwoKMeo41uFGSrsrHaLgnO4i3qEQ90
T0+GYlVW+SFKF4k81/POeyOMxtxbTajd9L6SABEep9SuhmvMCMllPRiYXUccH6lH
EinnkVecMyEEOAXZFfFFdSXMWOQ0L+dSv2wHO5nyF6BgaSHvUV9hJ8UhvDhi3ieA
QwUcJJd7nWrvimfLU90ywwh40mKNFw1f2fDy4t9WM6okuxDpqUVUn7IEF0OuUyid
e6kjrqrl8ebDofh9ZZahL3oj93S9SUgx6y9rNnjpubcvdqBLKygky9Xqwl57gwUh
gnlVDMXaCarJrHHadzIOZTXFZq41JTX6fmbhtoV5NLIm3HgD9ND5BXU24AI7pjQW
NsxyOOo5RZUL6+TYGPK6hshjeBxlFQsSaTMzGGNUfypzg5oytl+SjbaXj31dbUq5
+yOrozpqh/iFgJkpMqtGof4Vn4qzovIwSvnhaI14kNkPcPVqI63ojSModn0U9qkK
i6COpuY5s1FvMdSBscUBEaR0dnFayNZOP3JqnudikxLdGwUsBBYOmC6+Gp9Ba3M6
57pZ+bAL93nzH1WjL1x8oJ2dyt+5IFlARULPCNhi00h6pUhPDOyAOnj2A3LpjHV+
U14lZzhnXR0oNl4wvb7rUP4MxCKlBSrVVnJamr4xNJXfm048DY63w1k9OGEy0dpb
wSLkZCD356pu7/fYcO3gCh8SCINQ45NR7e3dDwv7gZ3g6Q1DcK+BwCwOtnjmqI3/
X+UEk5ovwLMwfsoxDOhmgYxra+H5yoaKlzhlT9J0IH69hfIfZMwlUdX33/9WYp6h
6t3bsjw1/gQcuG82l0X3wMq5M7vVCI0cLSnacM5Jxrf/jNiCLFJ60E5nlJdIYUHa
41oMxAX/P+1Z5H7j3eVBXX1aHP/4e0NH2v5xXWvgUVYL6IkXUNufNFv5Dptplnpt
74FB2VbrSSidOw3hJ9oWQyfE1IDDcKhtnXIs2fTxrL+/SVCdkrBHv0myxM5nob0a
GhFuwCMVsL+0ZuBJ5Vwqqie3Sv/aP0Wb5K88zNcuRyCEPjwpRN5LM4hETZ/VryMM
pT0h8R9sk8hGlZ/P2IESKwIbqsIu2h+jK0SNHMi1ohWpENPkzxqfh06FXU4v5soH
BPQose1pi9Im7Z5ITcWSVjcpUrXjEApS/lmuzsjmy2H3Z/dHQ4Z6zCKT0RbfgEsT
TF+sYLtMEwL6DWFp8NlqbYMH+pqQCCjECJ3jVRtJoZjMyZKrCSPnyVoc6EL//MO4
6iim9vADut6eZ4HuzN5EcRcLhuubB2pRkWuBqqGFZsWBr+lhnhlAUpm8WHwp7rqO
BqNNN7Gmca8tmbAfs0Qjffvk/9ionGY2cq1CxM/qPlDCpNCpUQWKB72+xBR+TrKq
R8wCkl1qOm1AMNJd2Q4OyU3T0FdGsZRpBPMBCl6UI2iTZs5iRQl2p8NoS1S1sLBr
kLdwfDUaUk6H0MrunZCulEmci7jbt3L2vHuw2p8RskzPQEgOTUVwFG6Fq1hi2NwN
`protect END_PROTECTED
