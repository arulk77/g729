`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49BGfeS2OW0hCHDeg8TXZpuN+mxAzuZLKYxeIHlDdsST
eNMotuhVGHr19ro/wz2uuMSVE2/lcRuqtFsCBrAZ6vVRZgEfFlMZiEY/GX+TEFP2
BW+CrcMGw687bVEbxrUhtLLKuIBx6jO1Il4/hPC9bpKf8P6qg91Mfw31Gm8J4KTF
nB7zxMTTRFOQQJX6nn4NuLQPQxSx1gsd20YENcvW6fa2p3MR1SJ68IU+8rznKTo2
6w7g0it8X4Pkesy/7L3WRG3KljH971KCRx3YCCcICHY=
`protect END_PROTECTED
