`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
UYlbbMBAn51MCx6ui1jwulKaoVbLDpf+g3GnPQtQ/7NVTuFsXzVpDkJDjPOWUQWU
QBlB9LzLQGkSN/sxtnNbs+05TBxKxxSe6znz7ajkd649CL93rkKveC4fx3NTM6bw
jVcT4+xz0GQcVTQyTeYqvXGHWJ4fqt9Y05SOfcxO2EEyDnBlgGpulDmBr4+aas9J
TrRqN/NogCtcDAVzfUpJSnpnT/Egh0NescO5OFsFacpjoWLvA8KxiqXeid0uEHaF
HR6m473mFEnhSuj9k0jVYBwf8XP3O0GwfEpW3BcZeEw=
`protect END_PROTECTED
