`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMjb0SU9VYoQ3/h0xgk8apqyEK8eegQKksPgIW6MtdkU
L1MU/Sr0LH6IzwLsPf0f2pApm0m/VAIKM5wX74jfI/GBSzfg8P/FXezcmCQYMRDq
PcYgP9nFUYvbNdp0+qaB6Afl979rTY9hasbRj3iHxMaUr9Mz7OtkFl+mFMQEKGCp
KEBPpGXvLSUAByZ6QmZhuNbdLZKeSVgf1mqnlYtJtof3KwDU2+7MDucOTePeAaEV
zqJPlgBffPdXlq2+CUGYh1P6STiA4DHcEimPR3VS87spPjRE8gdH4D/XnTBNKKSA
IsHGYrMfBOcviYkM1ptU4SOhDeVIzedbsbPWcLP1Ytp/p/NhVV2FQLh6Uo9RiPp9
b+YpIYeWKvZPNshnvJKCOspV3JxWtcaLWZfE/WyVCpymPEI1HrpZwK0zW9aiaMJH
Yk61df7om7lD55wbMCABdA==
`protect END_PROTECTED
