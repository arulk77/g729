`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJgmOZE1M1AuMfJ4jI2BY+Gj7hPmY2dYke2QqH4Zj3Ot
d1gomWxBK8ooZOyV2rfC7Sla7DzEp6O+UpCV1D++xLPGLH857JO1mZKlDnV8yR1A
O9K9eumVM5BN+5VEFiLrL++HuOYhKKAyy+46BTgQhvBIzSuHngxwvWpSj5RT09Vo
obkDrReTvgAKgh89Mz/wGRnCVSYBiQPfhaD/dC+tgju6WV7f/Xib6PLo/WBXg2/U
Dy8JGMUEjQIL6/7mHiCfAtizDjwJ2cgeoUh1LP0/5w8MSWslZz2C/vDn4Yu2YSv9
Zhaw3b1qmn6nm7MYrOv/BeZCEN3WWdm3UB17IWnLIlFnJ+9fsMqk/R6kwB2nZpfC
jGpfK8hgBJnHlR7Vsj2Ozl/HabCAx9361FoR5JEsDSRTyhg5AUlaADIENK4jV85A
74AWQ22+uprAH/Wzv6/xY8s2mmoeipxmVtCPcTEr+MV4lGYrKHttQMk3ibCxsvxT
aW+4kZxDEH1Ol9MXe9YtE/K18xekamGNe2fG5DcU/WvlHc+jDiCAoxMzRkaF3hw9
e5iPqX1eS8QESvmmxVcvAT8IJHjt3NnWFkZosPMLibwu5o6ZO/nrJS88NJSwzgEl
`protect END_PROTECTED
