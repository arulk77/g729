`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
tJ6hSSxbUp9/jGPC2NIa9etXStHhRnaU+mxrbRzeRtCkaHKswFwJ4uzxOQtIVFj7
FBB+KnPCVNCpqAiahlQ1zd/E1P4v0yjcxQJ3qrwFNmeULI/p4z6RplXJ36pcQVJv
tr8E/t6DBfw2ya69RftNECTi+A9onnXQ6RUxJnNLzIWK4Bu4TxZd41h3an5BAj3N
3QrdvvziykwDYnFiZ1/kmfU0gP1ZR2N+xmqJGalI6ioPukjaDLemhQQzaovz9lXI
zYyua5EGM2ny5Oz0bhU5qSnzRlJ3AKEGLvH9J7/DxCM7dupU2DiXmFzV/Rr0TMyx
e3kmjYBJPkwtau91+pH+1/rQMLyQs6HLgk+bV7PKM5DpYvgjoQXhOPUemy7AtnI+
TWYIbFAZTMlNIvpVWVqI8ZAs7mImYrXHqxWcyyFWN4g=
`protect END_PROTECTED
