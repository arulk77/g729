`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Ia1MaS/SV3A/sKchKE/MkmA1DvzYxKBKatAkn3iUlHbPJBjToJi8e9clpClxmOAs
oDH6pbXeKdJgxj8u/He80iuVmeEyraWd+XmuqM3xzl7soMocnsixUHZ5BiQcB8yN
F3S5zBF6tG8wG/XqqPAcR+BoUtBkb+CHsG+J+cPstCGTr95A8CLTkPcDS0wcmyo3
MR2A9TobN5TeRgeuutkrJeN7E89Pt0nIAXTkzvQ93rgKsV7wdFZagJqh2udgAXYz
`protect END_PROTECTED
