`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFPtCmArM+2DQyNSJC2xmYENRQ3OYJcjTutMZSHzgOPs
CE1CSfmFlVMNMM9uqWGJ9aTub4sZNvHYWiUHH0w+gmHQFcPoTmvtc1QBfPBxDZdq
sFGGRsxNWUAGG3IElZhQPmTdWnoBC0HgJcKWgQfB+hGaaUY8TyKmr5ToejF+dqu/
miFuNe6+MFZ6nn/LBMIlxA==
`protect END_PROTECTED
