`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
wrYoszT6KGLxnW0sucCjC4Bv2j/Ogrs0QddwhB6ljY/BFVIdzXmsdtlULRKKX76n
U/T8W3n2+3C5gf3754pJ5lPO3GqJ/8QIPL6e1kLzS6zk8h+YZkpaVfPRKAO34TK+
rNe6z90HXovxpy3JWe3Mkn8aOD1nr26NsuMUY+w6F61f6U97AFwbN43DdMV0ZiiS
yxO533KNIllvsN767Pr/ylmBkElrXMYnJ3ac6W1fJGCA8OMMJhl2E/uvYYl8xawM
qq+FkuXkPFyKq1qF8A4n5MjzYnQeTeplX3snHYDFI6DMckUtnLrXTw+D1j82y9d3
TIWjNv5Ck0yc5gfZmJIIaYkIze76rVOjcTrrKo+cs7s=
`protect END_PROTECTED
