`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCXPunFMK7LLCJ4wpYlwKeESNMTE+6yPkZksvQVhKgKK
Ceea+yPbs1lqcx85VITjb89M2VNr0msxPfhQkSAzzBLRD+ZdBf6wGVk5SS5ED5fy
2iOL2cNIdR4M8m6UhDHFdDq2TviQMWJFsS5oGNoJ/+Aro6tJ4NkCsu13OXQieKZi
Ka7HLw7YUW2jdYx+BfID4+5hfb+lt/aVFqhqoMPrDcgix5uXqqBpYRrUjHGRhNx5
Sr0u5eU9q9DlO/M+U6B0IWzhfSTMOompX9i8aU2bkyfvJ6HCiYx4joT63RxMSXuu
SWWmJuU+exKAztZqsvOdM9snZsG7Sxah+pGYEaXPOcWF0ux0YKXkMBhDYe9ipa0J
QLlvmWNu8iocA85aYPuigObTSSIqCSq+og5sCa3Dlbebsop6UpnN3cGCK+glj/nq
MOMaMcQ9yciS6QqhTEl8yfzZ7UxUTW9SQ8dR1pcIK4kFv8zD32Y5LYtlAhxegTsZ
`protect END_PROTECTED
