`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOT1UUDZUycbpW6ta7zoGfh09QnTl8j3Q31MMgzvqcU/
CwoN4mcTNyQrGXX8yXRD9Dliwn3SVJmEtp1ONrtXFGp9eZ4FIr51ET1O+Xl1VzK6
77WqIp1VwLccb0OLXtQufsOIUUMYPFgvC/0u49rqx5kxwoBSlNSdi2I65g/W1lub
XPT9aLDfciVHCe8VypxpPxcaq09UUYQ2QdfEZ/aGXvfdI5CPwYzvymBdgr0tFFNV
gyQcVBVtIHCFSgLhhur4QV8YWS12cchna/7XD7XTltSDY/qhtg8nRzixfo67tbBH
BL4rSlgbN4A3K7HNze+66fXGmO/wxs9yGzXRNwDZgwWYGDv33NQDILwQw7GbG1ga
8cgEovpJTRYMFq0fSh1CNHbm63NpVU62qETPi9whX9rI+jww/4l2ADroiCMuBtgq
6ytIHcB6SCFRPkUI2pgWQ7HtprP6Lso30DS8YECTWIYH8ObKIsD0bXF/oaR2UPdj
`protect END_PROTECTED
