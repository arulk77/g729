`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI6X1WWW0cqh6/mdeI2qsS+VK8VgXB5VR0IWKG9ArRAi
OqKK3p7nxlcW5NIXctg224cDVaBux3+7hw4/SFeYjLl8fEYpD1wyYnWNzC68QX+V
4PBfoDiYLiQR7aGxYBa3GHlVOqOnTLmZ5erlTvxdE4pva/H1h7uGbCSmmIqgtiHG
QhoYbJyO+H3kgbnpr8LjoC/ItIaVj7MTa/rCiDsh4Is7btSpqdcFcVq/1/dWvO3p
C8JCPop/PmmLuzOzcQe2voNfkPd45ZS8g4vHYmSIb0l2uRm/HmcheDCfECpsGnb2
SgoanEK2542eYpyCaiwf2AYGTlSBDXo3gjj3wwia2sfA/d1vaOQrMkeousiNAv/3
UN2BK0jGHN2ooTXWT7bhh9AbfRLVb/aR3DVL4i4AMXMC8mAgB5WZPdtGqiXVVgwf
eGncG4IQtSJh9TCh4POID4fNg+MgQhoxarV/TDZXQpVfEFB+forh5SO0Ab5zNHV5
SoNMciwKouXsQLWWH4htYbQUDhm12735bm8hFw1kENQyflvN80EbMndtgpabVz2f
5lgpL3GnOK0OPGdeRPAZN7pTy8MOs306SX4oHeKHEl0Veq6BhzPRB67fHg3kpI4R
rG6XvDIRdIkuLSXKPF6wG2JUzsaB/7t2KYZxApZAwPDsk6q1G1cGz3dQGCfQyL8E
`protect END_PROTECTED
