`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ZXn8YuyL6A/gG7NM+8zVrDfKkDfBOTENRiH5Qm4E7KNrDxc3GlX54ZWuh6mb87cF
4rOigu8aUAhsu782IJrKs78ZxBv8vY6/zDozpX4P66Bm74QmVOVvvF4ol96SWB1i
qA7SlwM+qu8W6gOk2HBAak252rzACwFYpmiREvoAc3v1u3Qt3/uxRo44vFReiQf7
cm/vsEa+w+4WRz58ro5h9cT6u0FSBgocZK5b8E2xf8MCslaXV14ANvvlYYCSPBP4
N6fI2k2xVoKwIH2rQXsbVsyJxzWNeiHfmQcwb0wIQgEeVu7nEs01bOH79SiEoR2b
Rj1RtDqHV5exb+UhewYB/rkAtTUhyaO06X+WOoEvVM5d2oMnuW0gjFu5XT2GosKa
uc5iV7ASogA+dZml+ChxbajN+Ncwl4rt7EffzqVjAZ7T+rNQdsZEeIR2xVa7a20/
F7WXEmY4URZ5F7zvdg2Y1LzVEi/viKo9Hj8sWSImSeI6iGiGnT21o3GYTzADzAJ+
wCjLMv2GSJNcHaQBEHWxRq+hN3aE2L263G/v6IQM0zRlu7+lj48w+jIxkvsUjZ9O
4IfHWQ4G6tpo7qpEqiiDP/0YJ09vvp3bA8dWwWrsSR2qF/GX/72KWg4sFvaZUpH8
+7irRK92K5dNwo4Wt+/dg7LBKSxo5NMyNeHchHYlkXt4zqHDHqPV/3L2Syt1Sy+x
aUdRu9Gco+o3JCQnbWpYcszos8o0mzgtQPzXSkkkB1o31E83lYpu4/++HTcwIhga
XZCJhxXGz3ZYL///FVG/MKIm8lizHUx064yGNQeKRlVPPDQTWkb3Phf/yPotSKeF
8UE7YancdeGLerxVpnEdL/mSBiIxX32ViMkLQA1L/qCYC4m2ILIxv/JLtFF7lGbf
ZLOPYzQtdugMHfwsgvL9ylizzHU3IoIrtLw+skxoDhVyTQ2FQa6n3Vo+lLpCzRjK
nKxtpg2C71+iJt1Yu9IprcqAFafERKaRuwaLRNzVeUB4BJc16XwsXYTyEeyoeyqH
6/JO0rtYzfMUIpGYmJnr3tcL27hFnB+M0/+pV/fq4DxNVfwtryGgqKyDwfTynaL4
1pOKMQt7ZOOvSPOoeSlm98yYwslyXG89NIBGUe+AdTiB4zVhd62jIIzPbafNmEq6
RJHj4Vv1hoo6UgiDqVbiYQ7CYvYjiLj3kqYV/2kv5/wDtS+OpCRaAgb7WvU1HfXq
s7j7pJ5x7sXaRsjPVVHnbk1EeyUwFSwKtgsFrE4xC5mxlgyr7VfDjn3nj+p7YF4I
t0q4Ufq7HCdTghwJA6uyHlyx00G/60jGIlqMq99Rf9FfOtnAQ6eITCVRpJCp7QBe
V4QOx7XtKvi1/2j5ht2IayI2HB1mPG+bUnp6uhBlTT9ltbFp5XI04bxX8+Qu1EZ+
ztU8cboifq+m1xCAhQcQUqwD7p5fG8GOP36kGLkEwL7CB3qRUw19BrlP+69VZNxU
jT0a4nPhE7HVvQorAOkYLxOTR/REi+gtN7Ft0vuaNqzcZxeX6xTyF+DKvul/hMi6
0ZWwV3tq+vz4jZw07EVNfQwL1k/Kmw9gFX9mut1axJJxjlVstAAnUsmOViyfBd26
RgZm95BxHpeePOOOanI95+uJ/AuiqVCoj8XiwEbiyblkNEeIXfOg47kKXJEOZJz+
UACOXFDXoSg+ITpCqsqFAnMc8RXm/tyydGbGlS+6v1GlRf2z+L2xosCCrdMvhpoU
xnVAs9j1hGN1BcTJBN6Fi6PHkF7jQFrO/ohuZCahVfuPJMQshVk1nyycJhqBXRJM
LVVSLm1/XLfX8oicZZUeg8mx2P1lxMLCWhA/Vvn0fkQPws71Iv2KUJ+FF1YmLgrR
hpt4MDa2PTtbjyEWF494GfjMKlVkh1pgpBH09wfXBJ8+lklVmU0I0JlbuBAZiWmi
Dr+ooKAkkHc+lmJ6jRpjrsl31xIYfwQ23z72YSxJoUZjMquVcplMJtiUXEJI2PgZ
sUZKOtoN3d96TKZXoDAohXC3CJxvYtW/21alnfWJCHIqTnPO+KxXeryt1DFbJGsx
TOPIGIJipiD/9gonuB3s1/o69ydKlP7982mIP0K9p9NEf1kbXhXHPH99hDn7+oIJ
bTcN8WoYFUWCjPLCzHmiBiZRTaAAyHMJs788WoqHYtUWy4WCxFENoUKhRaEu5Tyu
uUywYiVGmUlVaPZ4bChR6dtVZCVmFGnElqF24km1BQQf9e3x10Q+DUncUYl5e6pW
B1ekNcJfITME8Ko7AJVvIk7F0gVOoycYHXEnmxzohYqkkwUfqOxs+JUhDPPTG5gu
aMdMZedf0k8Xg06Wk///Cfv1UARzvVcK4XxbKQ2cewrkg1m+4WcALMiWDGwwnX3w
l2NZFBDNuya9lLYu3SM0ifmAyv/K8l82Ax51X/tYn3LdGcPY5lLv+YZRca2IKlfg
MjRjdOAE29TBUc71bXyXhC6NDir81lG4rQuk1YzzTUXaGVjjPHyYbTUuWYvp92Ho
BELpn7hjIQ9wlogPvaRR+++77s+1FniFVTovvkSGLvanFaI/j9IfuKE1yu3HXVmu
XzietpHnsqF+kas5ppnNhw==
`protect END_PROTECTED
