`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
RRg911hbMbO/naB0XSMVl90B88B1UQpmaVNkkJ7Flj1WrM3KIFPl03wuXV5/y5mT
TjdIRAx0uyJOTy1I/3G4yxHesUSNKN+E+ExcKfI2QbdpPVgmMB9lrH1FNU4FY+N6
vJFYtjh6Rz4pR5NInfm31lYBhLneWEh0XrMcmIIJj6IJCHOG8gQ0AOjg87ksI3Un
HwRtv3A+X296IKym1zcCrSpVE56dp9Y3RpMTMhTVUcxjbB20s7UoMjk7tNnLqrmq
Byehj6RQyAVJ451R1Y9RHWx9QV7hjTjzpgJOz0ngYQDy/W2WwNWLCZksGHsKlhMN
8whvT3VaIeQbpQ3YGUr1EirMrmr5wdG1ErcLwZlagrSQVFFwZXniXPOnRq71lEDl
NmPKu+L/4/tInpb37irZTu6Kb0aWI8r2z8IyXKbb+jkugTbJkKSCqqTbcPQB0TZk
ssrRr87tVqaIgbdIhBqxke8uS6Ct17XNA89suqPHOZ7FkN3PFz4LS5xunObeD2LP
C8qQmj8RyWKq8hWMJVxiRg==
`protect END_PROTECTED
