`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHqWDvcdcmlk/RQBAiupp32v9sU/aLxiFVthVPLZHk5/
z1pTBq2YJqT4P7XL5WjKS2t7KQAi9l/7/k1Ei+RWIb/AAlaTVbrqM9Jx6ZBXkjhM
6Njc+KLTj2Y1bObAhTsiFMWiAC561VzyKXQItQLTtqVEuVmJ+y3s9Tqx9ZrrMTOo
tZK1sT53EjX1IDODJVo2BRT5v6Y2hn15gsZ5Q/kQgFIo+4NMQlCN1YPO2t5w5pni
kMGlvtsgmmRK417pNPA4IrhyzPJf1hDFGYrtcmLXeHlwVpsW/C2/+coYTAu2lyNX
KLYmncePr4vGP+ev415H0pEC1URf5X6UWVOq3XJoZnc898WYnSMA6hcSFivDAub8
mzl0pc/+V5VfbDsewEM/rb8PiwltLtBnBO/NFluZ8P4wVZU5XApg/F3EBWilyNsP
`protect END_PROTECTED
