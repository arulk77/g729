`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
iAkvybeHBFx5kDfJdg0J9qu7hI1eokGXTd9B5JqDA0jw5oT3U7K5yZGGxErhnYAg
xrjFnZysLKtjr2uf6u9QR7N7koVJjvqla1hBnJmDofssacANjX3hcIc50S4lSK7A
jr886bACGkoHV5GYrR4YZFZn5q96TnpmAP8Dd87lbS/sZ5fDJxN4qItnT8JZvacC
GfbDWB1Bl8ELFkfQTPBupeAmMq9ujnw8lhnlu/99A40bD298U5eAGBlncjugh/Ms
6RNc0KgairuPblBl9i1/MRxTwu2/vsDB7wARK7mQKPHkRIweb8H5F5tMyoSvPC3a
S5S2g+3u1GL3MWc6RbeLJv7F3k3vBipEE4pb1SoAWWtaOHo4tz1TjG6ZtnrofGeG
u+mJgks66P/bCpLIfKguXxC5hFVzOJ04oaIqqZXv8/8=
`protect END_PROTECTED
