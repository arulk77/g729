`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePKwqU+D8uV3lVruK0cFty3k+FCZ+py85KOU6O/X3WTP
aqdTNqU3TcE7avjslxVOiROijYAzAWC/e2M6g9TT0e8/qDFiMJ5l77UdgnDIpozZ
DN1OV6Z7I/BI1gtSXEggzyBueCTjmPXRfLhZnrZuoxn3aec5vjoGiqvyomniGedC
Cj++G9t/10dc6PLo51TT+Q==
`protect END_PROTECTED
