`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
x/Dyb9ubVC4uflIE4q/tkT+x/g73B6l7xQ2IA50e/0wjH4Q1oFrvGhpVmRvg4tGN
nNP6Rl0E40mephIZ3za1a/aei5rppxkas53I12nPoE1shf7qa/4Bbg6QAs8X3KJF
BDWynNf4tCnSqzBHIObSrNDGHjKim/uo3Bs2ZSYYx6uAHAdfYsVgWQfShpIuANyU
lnRVqFI6I9u4ANUi/9c7QZm9ihELTZ1bjKxcbsv8EA3b8M/1jcCH0t0faItoNdOs
x2TPFHJ7uTdM3cupHchrItYAqVgb9waBs6eQ3TjG9tulHLK+Yg13HLOH+5yRy0bz
i+GkQO66/vanwhu2vLqJNArzmQOc++c7uLYSqvPyWJM=
`protect END_PROTECTED
