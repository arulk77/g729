`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMOz7RI10KXkcfBhQkyXHewgSBBir3mxIsSMKsyGIO6Y
eHosIXhuDG4rZJueOlodTx0X7ypo3s7mhJf2evTo12yg3UxcVrwDNvoFEkrwfevp
TWe3NEitZim+fg85BetPjRF74KQuIa9QyxwAWw/917too/CBvLKZd+eVVUQavKhQ
FbaRnrLWp5D7G1EkMsMCLbTxVEbJdH0WUi1zd4OFXDqHvj9uFRlUk2pUO+8RcMud
BYXfZNdhxc6HuVpJOmBo3YQCZMQoP2mZ5Lgfz4ljAXyIb4X9xNkb7Uh6kHwNDq6L
ww6/nKqN2oxg1m1p9PoE+aAVF8pS31Eb4kRi+5WW2HMX9xfHqIx7GvNWZXvhoFBF
j1W5oU9GS4s53lYuoHyaTlxODZKCiQV6viQD9zVkIwzfzebCxP3rVcUYf77B3sGk
YKdasdwiDacsr5fTHI3d+z9h8xVBpVsxoq/AJmVB80M=
`protect END_PROTECTED
