`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEqziTKvds5yvZM1Sxj16ZIoAckfWnb+bEeO01EFB9RW
Ko++j1Q7Blr72WIAC9Ap8aBQwZPp//i1EYJRMYdoM90a6HmlWCKdkzX4Y8md4oQH
xmsDoka/Q9cHvkAMZbtW5r2l9YiLQqp+oekZB3sv1pv3s1EbuX25OR1GYFuqA7oK
VaoO4znrZ8LKeHD7V+l93acjNK4UvTDZ3fF1X3jN2uqc2acVuofjQdq2EQ31/SiE
An4S7XXopZ/Gd45xtZt0RZGxHYGLZRLpUgibPfiWV+SzjLLnTq5jbXHGin6aBCps
nKj+nmnW9ZN8/dK7BRxi4g==
`protect END_PROTECTED
