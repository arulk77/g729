`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMQ7gcRP8il+VzvGc0cS2EGGzIMZs03g5+vBy5KOgTu7
1BiJyJNg26lZ+GTdtFSHMFJQ4+cLzI7Rk/IQXFUAqIYC2dOTD72pXNE8ZS3uEU9N
O3FMG2/RqitRieCua4Yt2dWUaQBHffXInK2olK1+FQ9WvS0EwChocr0fFOTd+VZR
mu9LnlvLbeIlNuqaQA/u5gr72/PF3vfmBtLqY4qAXb3U2Kz3vIWw0agqAvwsBsFK
`protect END_PROTECTED
