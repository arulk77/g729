`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCaV14PaW/aFySnmN0/6BuLUJN0YfTyF9jjyAbF+tt2R
3B7e+2dn2DZXVHvKrIZPWBe22PRnQIsQJAPjL5c4DGi/VJ5ItV1uYXjFTw3TssHI
K+ne2QokPeh3wWyd8y4xyfw8wrfaZkdy7XFpCLyhtSFvyHrIddPYt7cs12jzGsO2
MOPCUSKCH0j48onn2v2+csHO7c4xtCXVBAIDTKyk/1WK6cyuau4Hush+ZGJ/FYvK
pwHSnTTwhviO0oCT0iD9ERW/ho7OOVKrRMu6SOf+cyuCPYd9x8wBdRscurXdkpi2
uOWAbPVk4vhWTPIru0O6jRJZsrNDY7ovX/UXZCVjraLf0q62b7RFaUh/cwFz9ugu
pK5e1+6lSQzMnW5LUluIo9a6Hr3v/shbxXJajDRIb+3wHSCmo9UJgb7jrq3B78go
IF3qHgV0PsVPX7Su91rjssrL9IQU8MN4xQgsiGamZU0ey/endCtxULg3txZigxVF
oNZJy0Qkl+aKOakuu6D5ABSPTifLZ2qQ3cL7o85HQw0giM9LWEbjYS8Jp/SJwkSA
gJ26fVmqC2sFNaWum68R4zDA/qI+2HjACrj01aEbizybQ28FdELEML764jJ2g9Vz
cH6HjMlEIT8g9Eq4ub/f5QOsUaWMHN6Ww/8PBLIQI1cmR3DJ/C5oHdu6xN7uKTAQ
b+I+MNIvC5HBsxua/88FXrd2PKHdnNbS9MlB/XHiZPdboaQ52TGU0QYfRreCfAp8
cT6mPAfVV6qL8JNcBgJbyPCuVwB8gTyXvxZPK9pqY7/uM4KzigK85zZz1iPUzbkX
`protect END_PROTECTED
