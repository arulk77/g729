`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveA0gNIDOEF65c03HUE2v8utKdmWsIOW8csm8VCW6T3BX
da+pseLsk3nimA5bF7mRHqyq+NpGfzJSaToc2H42eBfy/CWGeL5/J8rQkjDO6d17
kEmBBhLH4WMpgBsiqqE+iYlZg+/g00gDKbC+R/BYn0S5JMsHFO7fq9V1sJQCpOk+
cdBHaWdzlu0p/HD9h+mrtZvBlLlZMUldZbYxexlhxiItYNemL9lejytWNy+uSLK2
`protect END_PROTECTED
