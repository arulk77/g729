`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDh+94bf60dLWpLZI4T/FDvyOoizvlSdKcy0C6418Wf3
EQ1LX09WTRgq7k+1CLCfQNzSIhOJ+/676EFpgiYmsDPWSMRhb7hGEcOr+sKIjksN
DddC8UBiSic6E7H7PO2ymEjSiPDBhNvsTHQu7+RHiban17Ou5hC8D377wUE7zmVz
09spUyxOGol+Ux/RStNpw9eXTaRsVs4KHPc9y9oiForxOVk6UHKw/hCpdd1tnDkR
SfAVdtxdHgmmi8gy1vm0BSZQVEONqL7iS5jpkJPnbAI0G0Fn+mWGOnSvqXFDH51T
qBPKOb9+PbqQnKG1uCv51oc/r0CQYpuqiaEEK6Eib5N+XABgkBbBc8SkzE1vqrJ7
XQswQ/4x0YjuQi2Vyy78LvUPaxVFz6cztisw5FThHDG1kgp5xkDvW5VSO2nrOpL7
Gqtegm3bi/tmd0f9ZILRowBxZP7bAF1OyhnxwEyrDOMq9AbJnUCNvZs76t9XZkcS
9O1JKJFnUWLG5ioqw/w+H0VplQC4fO8NijyeVsVWO3lTDPQQ+c1UajqNj4+C/6d1
`protect END_PROTECTED
