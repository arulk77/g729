`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKkhajp5cl/4SII2qnZ71nyMOMtOEtigHFFPGWnszwQc
HSOxvv5oo8eESDGTnRui731KEOIZhAGZHn6qbmnuaRpKfMi165izf7GHIkem5EAO
bkdbUiLA3Cr/zij/WsESLg3cxrZT3mK2v9GXSPyzkC7edZ/hdQOSVbJRi/6OHzsR
ssX1R6cCuzfG7cIwxGwVpZIABU6SYCRXMTbqYCa66/U7COzdNlMqYO9+5z3NBEsw
2/Q40e2stxEaiR2EhoH99anwf2Tfb08ODzYF1CYLKPAI+0kH0nDky3jbjkwMpAhR
lsxTmmGsbPz5EOqU24+sVGNfRgvFWy7qs6JObZeBTOfmneOkJRSEGE3d2gcx/tja
`protect END_PROTECTED
