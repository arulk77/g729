`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45U9vV8cy4vOykKfDxxG1A6AzMltIgMqEyIrn31HrRSt
7eZ+xS6OMpE0wIL0eZlT3999DEJ1S5sNNyd3S5TE260Ayl9cIzTOaJ5WWdvugqk1
xNyEfROm3GRkTUwTXVDVS8nDV1riXZKkwbA8yDCL4thN0rRY+z25+aDO/ousRCZT
eQ4yRBhueb02OSgDsNeyAQGgcOIdzQU5oLt20jhD8dY=
`protect END_PROTECTED
