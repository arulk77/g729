`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePQG+51Kzh2haVtXvVFodiJtaveYbgODkAqmJ0Lcoywj
gcmjNiKvA/NToKCRO0qKF4whg9Mjrgvzf75bq724hbT3LrViNRRoQz2g73KwqjD5
dPyxjPGnzoEZ7JcoPSu+XdBPh3uw3Vdjy08yASWE5Hb8VkBoH12+oHrI2ofLxHDC
cW3gdUKDPHMDSj3kTirkME/S//6iOJ6LQtkYIcWlkgqZh/nPD8j8gPZz8X4bdUdI
kRWZ+OlpH3k37qQzGd5Dq8gRZEKUCI3s0CPgzSY48bXXLRuFFhgD2L1/295G9tiV
qoqN8Zs0eYOtlVG2sGRwiI8FR7nA8b8BsQOdNvuEBF3vUC0ubl7VwK52zV1yVG35
`protect END_PROTECTED
