`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCSKQjmiQoHVzGtgpNLluO0TlSMKs31PUCibr2Ci5C/u
ncIBIDbVgss/bRdNVlW3P4V54n+cb5Yz8xodFTam4sK90hDW+bScNG71A682HWQi
20xDP0ifAOzsQZj7Nd5GSIzXxA6m+zT17sbg0dARYL+SKaLEGSQKDPsKyCqVO62j
57VsqWAbAyjoX8iEg4/B6Eo044N3fY4EkQbbvqvSOX3ai0ZfBAbo79UHIbTLlRCR
oz3dmi8c2Mop6+ZpDrVZM2udqXvngDftYlOoJpa0R/A6NKCwFEtXF5lEwXyITL6M
QTnGTIp0sqRjIELZz+/DLw==
`protect END_PROTECTED
