`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48JwOH8gOFHerT9mpW7n2o5cUv+fZ8ILB5+hsk77LAGy
EIQlDwq6L7WjG4p2MQiQ7ThNcsiXBkCkC7Xpf5RvVFwfYiegePfPAIsXZgAzHoa4
a76t+tO0hiIWR71/lSlXnwNlgrQ5k9yEs6m4BT74CXrllkOTA7PlmZvzv0Uwo+YO
2IcFzfJfDK2JWALphs9+Q5hvxCwKrwFV3qFq1DSDxu0fBgvQe5WpO/Oh2exF4TbQ
Guxzf9w5C3TIuPtKWN7OuSBr/3muqlku2bwOA1R1/KOhxUtcR6MWElPEbo21AvE8
9FyCRN64T2CGms80Ogzmrg==
`protect END_PROTECTED
