`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
XQ5tZ1HmkJTvGjT2CbmaK9opmA6/60y8p71YUnR+tTkdovfn/bofSgK/Sx+M3Kav
0WdKubf/GELWtAyVoiVd+wPZLPoZ+DU0/PgRO6fKtP2hUg65PW6cN3saJETagMxj
2UT0lEZrYzgzcewJZwH4WXwzyPGaxvGZNQThJoz9sprgGtfhKsggfbNszqp0/LWO
ySZufyaAu23YqG3Xz6cR5CiD3WGUDtFJtp1sJuATdN1WXdY3C/ygUYpkvEo2pYcS
dVWb48apG4tnayn9fWvpCkf8rjHgS9cLYJ/N7SP2MgcRK+3Ogu/lMiFAshiAmEzR
SN5ENI9Pz1Oe9nxtim+5QgAMjvR2B2vKeIwrQEvaUO2SojKJe+6cDesvFxYuG/xQ
lWBcnYNCn/XCZ+v6/YPi6U/JyKf7RquDXLG3RjiYK/T78L6drUTOQ/WcoWYCEXSd
aMkSLRJrRi/eX0YQ+TwSVHltw26bkpG0MAeDANpBGPznOARzSIejz6Lz1BMP2SYO
8Q5Y82Ha09bsnsprJblyunNLhRWA93wQhBfvBhhBKXyo4WJNrkWPWMvyXu1kVNt5
j1i2mFyymF0fhp2eb/6KyR/j9c555qGVhjaMCoxDIwnrmh+heft+xqKsCIKP2gKh
GFJg1J2c/VZBPfido+0jXpJcjCgro3x68ofOJJFgYXkG+GPrIQO2r2swV54pOPE/
V21HhqiRG3azryBFEIILf4Xa/TEx2+YClDihcJnNcevt/r9MK+dMu8mQtxu9YEzA
OFPidbSE33RcZvMjzbO1/emOmEj3p/nJQNN1k/4Bn1pMMTAaVCEHjoeb/OgDlKoC
OgfZpeWR/Kz22BAzmHL/y56Nw7jzJOTsD9+CMBCqQ/MXoDvDQ9V/QAWf7rRjI3dc
oILZ79bN216JXqlvWlNtOyg7nZN3j17fjkdeVhZMwBnRqiMqyef9eHkCdma9W/FZ
2WIfz+w5bI6yUS+JZapo1g==
`protect END_PROTECTED
