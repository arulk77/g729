`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C++HUFsWLzeDmhRkU0DwrOwr+zrYgl22r/NF/I7um+tj
d6waittMkGul2tHqbILeNFqoOHQgzssjpm8Bb8tqQ+r20SYbeS9NP8aivpb+I7Tx
CMaC6Q855z+IQFW+U56xNfAtnxWCWvxaNf+TjllEQa/DyB85GuuHI/Xg44SePp9d
OcLs5XyEUg/RA11b8C4mdehzQAvOfJGu8cXx3Mmxg4P2CedIHaBt0OgHyPQjzhag
su2tb6O43b3Djsk4jSDEFXqUCe4cBFC+8J/C+nadP5vWLtK3d3ca4xv9jra6W1Vz
ULE0IbvtJsQZd4rtucsuIhTsNMMeGjEfa1Axmo9gyNGDKQWwpB3EwiUrW0oSDZTt
fmJgnEEo49OhA12SzzdxwuOnCRrFzH50fnbOzui8YZvlZUIzVt9N9Xa90BKMZtrg
DIpqZpuPvioRiFVctB5V2DG4qTEOd2Och+cjFUMGE+NiC3FOTwbQvrXk1GCpZdpk
twJxAU5ina7i3ibYqN4fLPnut5HdOL3n2TbG+xIUxrSvUXW3ZPICAjP8TwHr9Sl2
eEYjiU5YxE6b+UyLXpCGZF5IpQI2dU2H5rHzctNB+x53L3BDZC7WLDNZgdrVhu9J
emuLZIMAfY5vWEB2dB41lu5gHZJ9I4i3vMNxuFjkmGl0j7Xe/KBh2HxUN6ASqU6A
SYgpRkLLU6mICrJrLyN6BWz8S5aDrPJeD9iCJGutTuoXP6oiF/jbtOJyEuSqjXu9
D83cGPTDzycF+LeZT6sXmlOX+nBZeWghqwt7F6/TsLiVYHxG+vAp9jWQb0/4sPNd
Fzjf+bFcyPpTYAwlI8OOqBeE5n4b1/dCHdSDvpJUu1A=
`protect END_PROTECTED
