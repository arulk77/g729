`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMNr8A3XM4H5NLcPnpWZ0DLSP/JvNOnbc+9+6/WYRxlW
z6yDBxqFEWgN2BJay3PJCzstS0GIx3OHwVNmSdX320TaIQgiUbc2MygdkeDfJRFo
NYr6nWQmgv4n+dKRU2i8fv+8rzTmNziThYmJj/C4kTc4qPXCoCsAuLKxdwQBInil
kVlf60ej7gmxvOPHVmRHFkAZ+bJ7y1KRRhMosFUmXPedG3IRAS7QVDH79UJskMjX
`protect END_PROTECTED
