`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGsU06+TXeJYO/xi65NGV/Et+0DjJzAMiNbtkSlQo8Wn
SU6SSNV/jMNdc/2HAC70UUthB/dYQs7lrVuysS2TsiDG2qgN44ccs0PdJgs2d0nt
IYxyZTgXZH6dkYNc5o1esgNVUtyL+qaEkCnroy9rEC+Mt+9C1zOQm3hUBMMUnldI
/ZlBx1PYyD7xogY5owd4B9ku6eD3t7IzuHeinr7np8v5RHFTPEWYagdXwPdOlrj3
INhZsg/fCpgjeJQ1t7WX8QzxIEPIqphrpyHwUiwdYkQ9jONfc6/Sa46Sq2ly2rCC
AwPLck6X+SBrb9ZCDl/OhBb32IpBd+D5nLcTB399a/SDGKhlhKt+Aj99xe9+UDgs
HafSyRehzeiER9Ps87eQugGiN5shHmvPe+3PYTDAeX3/zrVqCJZYtgh2H1DHGUAp
tup8vhJA6ZX2w3T3vOrPJLkLMTMmhKKqfESdxUF7EZ8BPVqGkrugPhPZetjcmJp+
EK3Ijg6rEo2zTEYYpgdjvubqI+5vSUmiGDRS58tGovLqxr01t8S5fc6gTndpO7c+
IoWvWpl8mPXaPysw8aw2CfKe/Dntmd5kK2eUwqRoQuDMJpqpTiXTq6hVRcQfQPe8
ybXzS0zVh1PFd8H00/sUVJYHBCYn4Ct/D624ZYJ5nYq9gTTK/MUJwoqmLEU7KKhO
`protect END_PROTECTED
