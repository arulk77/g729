`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePOoX0WfHZmjLnJndGTFOCuH8A7+s6HJ64JxYcIZhMsX
TAmn9hAqjUIrXCEtSbUk9FqdxrQbWmzEbutg7Ijr5LOjyNc7EOVYmCclwovu3f2a
070rSJ4GkKWv5qjxj8ZaFkU9i6bgo9tZoM3tCjANRfmgb65j9Sv2dTqovXaw40Ou
Ll5foSOzQy4BD/qJxwi7o+oNVuKbgo3YIHm1G2ELSXZ0PBA0ApQU0SwUabH9Vdlr
vDCOtFTFfHR8+wUkHtAvmbuxlZCBRvmiZbh+bBJ/NbAPJkE+GYPvUweDj4jyrKdX
9xtYxtMFAtiLv7vSFAMrNDM5fC10n68ufDpbPqySfkSiUP6xE4wtrfX95BMHgnts
`protect END_PROTECTED
