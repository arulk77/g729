`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
b+2AGI9b6HT4k5oWC90G9kmv9+5s+quVxubXsTPPUcgIrXYpePm7cVdLqCNaYfi/
4lYucbSByGEaMgeVVk5n5gwAKJ3p8POa9rLZWe14J74jajSfrvzH+sXEMns0Bjfj
8kJZEVJxQXnaDdSDwhFwS8saKRwEP+9odzuPZHSrvMpelPLJobmjlxwf1cYu/6w4
0wipJR1bqgv5kxLnNyqjAyVt7WYv0zMnmiil9L8foexjbwR4fP2o+7AvlDoFr9CY
Hb2bu8QVsftvMm+sEVHr5azuovBaoRu1D+1XF/bM0Kx55a4oEQjIxufxMRuaSp+E
x/xLkr/KYQp6538cgSH0YdkGw8hZvZD1Z4ekVzjOVWYb0BDN9No9wFB9CRDCzkWW
sAm3fMCjLINtQuWtMEmJgTkpaHVuHlyzTW4QrKczFyIOiXBvspalRQewsV/gE3h/
r1IFPHJ6K/ekovuRm3w9QmvnQd/pvOyhn1ychtrTv2/WiRoz75iRp9sOaYeRwQ6A
kxEheuyDwm4kSJ5c+kGutFr+XqR3Eo4Z43J1wkHhIYAvW8g9zrHTScXYShoS8Bzy
0bhNTv7kn7CmiajEBtabh40KpAw8uWbiLbU2g37XVmwn9JCc7JlZHc6Dbh9X9ioc
aCORGmcJ6+NtA2z1Ozq+QZeab48IhcTsuX3hY5Si0Efh2wM0OVs93QGvhJ6rApMZ
3r6CMrOcJMep0lMruXqJzr9cWe3AmPIc2yq6EtUmEB7rdfLSrLaNcrwOIAk6K1HR
ZId/g2q4GfgG+ZUARix6uq/G/HJ5WOvKqvCdghWJc5QnHythMwKaHRHt4T8y3E0/
fQVMgmLvffsI3DGW+tSZJwj2vgaM6QVnIwsMUYGaI3xR/BZL+EpQBkzbb68PDG8/
O4FSYvPNn/38KTZlfmR1QKa0HfTBbP7yXmjOHLbbcRE3LF4KYTEaMvagD5TFYvqJ
lt4jm97OZ8rFeY/fuLJxUN2dng4Wkv2HOAZzDBjAY6AT61XUHvCVdbx1GBgIikp4
4aLUcj4MPnlbfXtBVOPCgEcwbZFe0489F74DCQaZRywxTYMu3YBBX//VEI6duiHo
0CexJx3g2S5TPkjM8Nq0YrQR6uaqxcL7G3s3oqxUSGn8tYH6dz8Ju31GgXt6eCWW
lTGsszVEk1QUg5FeKQsMUVEeNGf/yLoz4HE7x9D/KT7Xm9HdeYcFpKGmtyDlOGWs
rhmTngXmHwn2Ls0igw9cLcrdcQ254BNa1v7B+HR0jGsMv14zBC+ONpUHe9YsznBq
DmTpoIEA23YcQFYb7k3h92NEKeWKjXA1CZ/D7GqDKKD1idcBJ3jLUL0szCFaQq/s
MHJSsCNIDPwHsTAQUtqBG3GJVpir9p3K7fJS/ylDj3s/eRVBjd2cCuhJcitTz2R5
Fr5/nCX8QFlkyAMS0S/L10nTdYytVAPlWIzHlYu+BApeJGZ5laJ/zGZSqocyP8/X
RybNkMj79gRFQPOmUdZjxvpXZKlqoGc4LoBEqiXzkdA3/A+5U3QNHKZeIe54q3sh
kRxzwnkuwNfVYwr8Bcr4M0a0lseLZru4nqxgnehZNP3E0pnzUwCS7Mc5izQTIu+r
eBc0zqZmPVZTb7eXv70tFF0gL2mf2Wq50qlH3OtAuBypDSUKStaYD+3+0ZyMXyzx
GqYV75rvFWN0JrrUOF5i7BbVlqbyPZYjbQ40UrVTxFy/2FZ8GTTwicVQiIMq+sFA
sJuqGEYQ5YU8ky9HNPbDOtV/ZsuyeCt7GP9dCjCVYPSlQmhs+xjAV0m9qsbg7Tiv
R1Xn2Z5I4R74OEyllqhTm4n9bD5tjnz1lxCf4HY1TZO/xw5rMYV0kuOH+nF3jUe4
d0B2IYlx2b3Z6szsG9IYe700fs4w8zFDjoViJrnx1vEOOLKH3ONl2bj7wtEwa8wf
vOzChRaW0H7s+VYpbgQaDD5kYeAg+KpC5Tf4YxKvEbgSWCM9Nz50IthIKQuBLH1d
yv2Ml/Y6+nOIiNZyBtfYCXpBZbg2p20Mk6ifOtb8MMXWFvtQ+/78ZdKlffTRP4l4
jjbckvg4FNMjYHXcmQotTbMng9ISSDJlWe2x4albpA04nsQKJNpBW+70ladCP1/x
zp7XfT05aiYb5IhFCwKeTfq/PrFNkIS14O4svYYbYw7dxzHANMeqa86oFO/g52pI
r1ySZ2i8msfZS23R1AVsbZ1BqnTDI+XbhUQjTIfrYNlU0e0JzO0bCRbXcWBZuJni
b+69kx5BCvTnpQeY4rpMJ1P5/CaZPeX0cNviPNYBHKzDfUKWX//1A8/o8ko0o3dy
s+mNZdc1eJV1pgeGzeUe7FYwCc0xRvy9xo1Ui0MiYENEoE+wZvsvc9ZwB/QVGQ6a
LdKMyaIVtpTWtz2JvLJYXVlj6n525k2ovsKnExTKj1RAPNF91305RrHqL80Jcoan
+r5H8y7/KxKNlzYG+hNSErGTNfh9UeMrYsEmdry7F+BbxoT4HfjsOdOZY4iV7kiD
X1jjSC5wKU+H2YX5ETmN9kuI3yZ2cceZ1RvmIw5qiFWC4JbGFt6mPWSTDww4MYWD
74KJidtKUjSD9rJOfgOr5RYPrQ94OrqFBYI2/Fs/0UC2ADE66uAcnBCEWhR8WG+0
Lyj8UJ8lnuzH5Gwi3sJ9bb8XJEkkK4N43JUdxcLXxbImShQPtKOzXZ8yi+lD+yxi
E3iInGNAWN+pB2/WPF1tnzWnqKzTN0uVOkKEtf7tH7n+h50n9sK3HCIYrYVCWmFf
7stmy58XqUSD3vG3WpYAK4ouBJ84HPvX4Q8jWb0rKJfrYovl+Z7k1gyTYfzLgMNm
6S88mdmXtftdr6tGeLjRcUrMWaTuA1M+Ambl4pqShnSnhSFE2nw/XZgAQVloK84B
mUIquBOckc777aaQKTAdutuSs041xzzPhlWgtEoyCgTMi6RwJZ8rv19lpfI5m3le
IYI1VGjsa7uGR9dalVBwxDaViox73NiYlr7SzJnoFPJCvjaHBIpkN8OCSZs0m4l5
Gc0qr/qxHH+OL8ePmPaHe/ygalrKYfUWpmkah9StF6Ig63rGIgsC4hqNIRwsN0WB
6Z7uen02geH52mF2UVsJaiVisXZCGUR3EzsMcvQExv6H64UT+bXaBm0cMyVYpUCJ
La3uprv6nhoyeaHHpiePYqm4pq85vCFwukksgQEQ/6QZG8BWFoMrQxv74akERnEX
f3m9QuoV7Dignjq+f4qgpeNKkkiX69dKdHozQvxlV4ZSKugdFO3CRHxi3ZLH1JdC
2cpAfpodXmdGFsPFj/LzxcxkOfWGq2GL0Dh+2P83Khkn/CGK1Vp+YqIxicASiHH2
Bv1Ihx7S8Ssb/+TjCXWsu+1H+UWCjJ94QzMvJcF298M7BAeVhW4mZoclYImQhx5k
hinplg4O8zfjGBjzHPAML843+DX6tgdwvBP8hD9Z9DLX5yY5Vj3ZF2x88CO/0lC0
I3AhZzrFEXwcwW/PO0BKuobcsfjyiDALxhR+GeeX28zS8AMWVa4lGa8/RV/SVaBN
dKMPXS8xuo1WDhSTp2v57cnPMSvmW/66BP+Qwrx3ugf76nQ8/SkBGXyWcyC/+nyj
0j9E5bmIFqtEMI0B/rqrVcDOoaHHOuW2+hCIhO2nntdvDuwrCQ3Mkvd4yzzQHqA2
+nQ2SLYnENpwkR0qmnLtEFMtpKUuhx0wq1qENWlqXpXSb60QX7ZgMaXMc0ZkuD6T
XatD3RZ1tLiG0akPvNbmN89XlKOvt6C8EPCC1fGiX2aEW6AqS1SvvKW6rKdvnjR2
twdfWd6lOdduVEVJuWwIrYh3Gg/CgFzkzGb7Vl/HKSKq4CA38eFbDtuE1EpxdjTn
nUSzUi4Lj/T07xSJpicONRQ8avsu7XYNhkdk0S7gYGFINWXEN/5NUSTsCQmxVMYo
vKsIncXREsjg4aVBZvq3hwYnlSbqEoza0VzS2oHi2oWs9q13DjvzaKhU3xrU7w5g
mPYtMvj5qAiS+H+UpA4+wlnuc/zgwKSuR2854/7q4LrJBsACChhjU3wiF6GX1JoJ
CBUu+qqoWjMy6wh2pLq8f5zY8hYlx9qQd7OZWfRx47RSvdp1xDajUGF/p0M4mcmL
M2Yvm94GLNcwKdRs2j1MMvyz0Be16/3g/zxrUlG402Ep3w3k5oPgSdOggkSoH/6I
80pmtyxp7vewRrKLpaLD+Gpyj9OtO+paIR0D0ADdcuA4GzSgZUaoqYw3Xyw0YAd+
cuOo5rbUWIk6l+5okLhhZdwfYnAVGaxhNMgLqYlIMF5aDlGst2ei/ar0iFW7k820
2MAjgIHbrAztocsVTwqvCLE8dqGG7zYP2d/D5iKehCMTwRC/5v33KEZXH9ElyNwi
2UPIucp+9ntcEp5N551UTT7wgKrN/TPKsr7s5V/St8LjqET99apPqvgFcMSQ9ETu
s2J3oYk8idtk3hdY2hZgC6imc2GnyusWYc2e4tVf1Ydueg4TA9zZWCaMjXOhmNgY
3LSneHJeAEUP1dVOKNWnFA==
`protect END_PROTECTED
