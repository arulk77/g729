`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
7k/+ajGkrYguhGZTbKtvX6LU1vuG/pf2RiYAnqdXWKKMqQXOCIb7NeReeMRpwo/4
D7O5jNMCuZJ7x+fT3AmlKtMXLEV/7/u+F0kI1djxwqxqDCZq28Nrg79GR38d1dfl
O29MOPCcjnnkEothuMJaf6Xk+j2TikjNE1AJwJ3AVVahUX3QDOU0H3GthbsMSKZ3
h6jov4V7QvX5Ma2/JDGY2Le/59uwnU5nZVMdznRxtsnYSrmcr7258xEGp2G0EcRx
o0lJsdAxobkcKktiLaUd5qtYexz/3tLMdeD3oWbdwfNUrCcUee4vXUc3/SNLAfkm
Hc9ZLrlQyRzIpUIqJfUh5A3fTzfMVP6HJiFWdq4ne/AtJaWCmi+fjUZCyU4ehiop
XbI4pi4byxWedQ0gDA23EsohNVzWslUCAfePaPsVqo3xadDDv6u8GwsBak1t1P4a
U6Ec22MK8ue6/wIQudyUly9H5CuaAuWBMWCRsZcnLdlo0GI+k3Kah7DWuesiClyB
hkBtV6i4ha2lLnu5tNWpgoMMM4sQRhefkEFjxXwRZrQNCvCyHpFAvwiZzL2vNGnn
xycmCrkf0VZfq6xYycr9oVOIMkCrRqaA3L7VQ8n+bmO13AHaftTZinnjzNodrWol
BjFZjVaZgOVqFNuhYIFYC64zWmj/ZnvPfygrLNDh3eQVtc3qoBZMHtzbWfAKCXX/
nGGqV+oFyU7AqfIMwBFrY6qRsS5tlINAzooauFzmO6mjPSCj1aB7uB+ydBF+flV+
elq5cTpAGUVMje95r38i7Dus0bShy+jFzlWeW6kIzr5EzMCi0hxOFCjPFJNXPvn2
NFOXU9sa/eoQ68JQj1ckEKJZq8ZxvGVNb2aWQsapbxZvnqdStdLqUc3bid4DGV76
YEnYlWjgFaD/gRosmmdC2QoJcSZouKKokjAZaSuwEhqJmqCzEhV/3kP8qiT/Kjco
oVESAsAARO2FpMlG/1APhGae50qMmmryGDzeJhVwPQJE6WrgrxsT3j4dyeuBCxx3
YVimu6Qg34t/fINDoOWetdwQPZsfXo57AzmdLVUaiCW7AuU/YKm9BlW/YwKOqdL3
U3F8MUSeQnnVD/nCBH7Laoid3fivYXrqGN9RmYKsG0h5g0E04fs2Zo6p2UFRt2TT
CcHChCmP+uxK7cDQzvVoNuFPrR6MGnFs1CVBkHYJxMj2CTIzbXyH1D3p+y7CYGY2
agBTjBOcFAV4Pys3hScjDnpvFPlqdmIksU4flwwssVGxypblG+AFy+5n2ps4UUZG
dW4fRg1RymBLw8TkS1Ru84TMoajYzKV0vsWxTa69UESjTSstP9kmgfq2yJoFclAB
t7I9oyCuaZUhI6f7VKqbaINo8WVjLTvUvRqsBpp5STR2ETZhVgGI8vIcIj9ijB/9
PL5RP/ERfE/71agMW3V0Zvwp9/M2RTgriwgUGEXKkbSWJ+n6qVLQzkyIaDz6WdSq
JwJ32O1hqK3zu3w9nsehgHaNcCxXa0JYisRoYz/eOMHWF9fRbzPoQa/BK9ZkR33f
xwEiXXLgK5zQbD0wD0eiwGdki0j2FuZa+jNu3fRigGH5u1LD/PWKBy0/zi8PlBJL
ZRllkAEh8QWmQjFFaKa89yjVrqAtAx64qAOIpFRq96WCPHZyP45+YQl88f3e1W5d
hhTgMFCs+hkiATZEwwyptH4IkslQGFcwIhDHu0NmfFiY4KFJdWEcIMVjdh4e3vw+
IrJSnj4LLFFao2a3H6kbSlrWDc1ac+9omxePfZ9QgqcmdRI81uoD2BVQ/CP+WjQl
H2+9ECYIctwMd3AE9ofsuMS4UeFQu6UJNsvgzReYjK2zRGz8QONFOSSHAIWnqPcV
sja+0wr6PnzWrhpfNPd1GJ40xTNQ8y5brYM5c/M8JG9NXH6e9QBGV854D3KHUGLW
xLlOZ8WU1qHvqY0IQYllZg8Dtxf0YJ90vC3D/Imd8nSeJAkKwwAHp5Jkpq4Pg56H
k+jMvmPomuv4sHwR0gKWx0jNENiFoYjmJlDjZmiK7UlrbwWeDi6T9OiwnnPQMuyJ
i1nz2PodTQR7JYXtO/8fwCPCICjSI9demAEaFuA38ESdwV+/2WK7M4apex/mWD3V
pRWVbK79vC0+O6C6p+OPYoFuXxkK9SYaI57r5bfgV5mHHZW6qimTjzsbmLf8zII5
UFyCsxOupxK40y2DqkbvqLE1EwkbLseuSIimFjAoLFiSL055ERGac9iivlmox6H3
r+DEYPGzjiqRnVgE/2hWvkY6PYoYK4BRJJVPNCkBDdFpc/kjmGiZgYkuH8BSljvQ
KAw0VFJqMvBMRa30wDQSiDqpTJu8obXZCJMwv1FJih/W6niIEfhVJQAUE0vOFBNs
T068eqH186Roohu6ZvfN3z7ROlpdyKSRFG+inN1wZow0nXzpE/qc/iROqIDN5RrB
YlVQ+km4fyoVY1SMGLEOR2so/CEP3IpsNwaEn/XPDSordnd5P48OTPU3gENGN3Lm
mAhyrm2L4o5ljvXBhT/kNhwJ6csxmBZ4thmvP7eJZd9BQqMoeu9Xom06Hti+5SaO
mFaLkKObskMiAa+tyQYOb0CojLqPPPc9WSmxdJhicGIM29I0pcVAX4UXsZVy+WBP
xRpeZL1zjvqJuVALi2SNkwD7WRRS6BR1h9FXRqXqiK/UJrq53ywOnefUZ4FlUT2I
bdmM5sdjM94UPIB9Mp0Ac9okzTyVvclvb24iK6II6buvWIoA40Gnxq442pADL6KK
2l9r953jGGxa9gzqAIcNClGazaCnY9UgawvIbMQUZXIeQ8BSILbDPt50ANltpARu
krFtltpsoPuae8SBkISk7MzY2Yxe2pmX11ob8G7dxxuhNk5lG8yaCNU/38DVvYos
vbAQBzEVEMqSlSp949i6Ao4DG9fYf4nAa2SLn0kYDN0ngkJscDFJQ+cjsCU9vHkM
1K4WLKw3UyFn00sLIHH5hPrxgj0tjfzDKpM3n2eVq1jOg0BCN5iosoATyQSO21JB
ILlntAixXXY1QKWfoduv/5SlPiRwAsESKfIcDhGrSLrarpc3Rkm2h6wkJFC9INPV
YnexKF/kQ3G1HZg0okeHANqNKq5wOzr2RxIxwlV7lvVy9jMwVvUjqO8gBfaqFXip
9F085clgAYEC+jVk8ysuJe0gt7a8433OeMHDsFcV3b40cjhVh+sZu1OsidpGBtPl
+5P6bL4LpswCOfimIZCSkmEq2qsmw4liWrQWW+tpb9nJllcvgu1oW85XJv1t4ZVh
bRhcTb9PrmTzbM3MQQ3z+ERlxrAHXyWQeMB2+wJzkQoEiSf8AlbKdruVbA1ENtiW
tyQqAJwi1Ujq0KqjYgQk5q1oqqP4vWnJ/r7ayj8XapC/1JGbCuNoEDtSR+6Gl9Ge
5tlWFp7DW6t9D9KfvR5vSPNwTUwFeTzwFGnMm2xrkX7Nd0UNYc++aGfdnrGOx0L1
VRA9jerSNhZ8Dtspcpp6ovzuSLwxQ7Wxz6r/fgwlqeFts/XBj3wwmXHvkj1Yx+tZ
RWqG2Mws7xVNnaLO+tDX62LmN7sVrOjEjlLsXAiio5ZbSHcw7NJqkv+0cmmIdnqv
qPZUwlNtxBFxhFxhR5+Bp5E0+3SWi8K+ZORwgsWZJPWlfUICIQ9dEtWaWE1M1RlS
WHEF8HpEPQicbtbURW+lVwHb9OGymV7meZN4iISoRJfDhmeHR3AYrYIvarP0v0ox
LH7l5f3T31gXvgI8loRXPqpQRhv4oDLquakvdbumYZKNMLFPt4bwefMuXhzGGZpa
ZMqp9hZiy6vEB9xyPyI9LZ0rapbKYhBYEf4kie/fw1NQGi9glGKGWpFvUu5tdwMa
9yn1QSOmBHWq+0WRJaa0iQDc707FnTOnpoXlL7jJebUauxDrVdoTuWJI+xv6+oaT
A04vw3BsK4KQ4cZA+uGX06fqAGNWdZijeqb0dD6oZ3TT4UrbkC9Q8ILvEFyvc/wG
SmTKDRh8VlkXAfqYP9aQu5FlRZaATIqXS0UFU75rF4PEb5zkAv2544UTfLWckIo1
yS8i4Xj2U6Mc1NxuW2OTqPwjLot1oGgtb+MT/fwY2Xz5e2wzfoR4AkgSqGzOYj+g
0pQKptmxRsouRaDqvMENBfeCoSN6mhbWJW+FLKOo6vQ78qMrmTX2MUTmx5V3hxuF
xLc+WSXImej6nHuvLsnkiMtCqkYJbg1O5fnivlFSpmr562J9TELt+PbXnrp2pj8D
6R9eM3oAKTIKM+tnahFxQmGCjngz5p6SmLa+c2fai/XSlAjiTiocM4SkP9fljv2/
bgj2eKEf4I6hn5k4HZpufglj1m1UyC7as9RSdmtUPdTFSk8+Ujc/jqssiwmqyQGN
`protect END_PROTECTED
