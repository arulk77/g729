`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aTELs/W1bsG/Y2H7yWkiIt9aL9ixzH02vS6K9kKjgcy3
RemNafqV2q2E3kd4W2SvfSm4/RJKKgWeHNJQkQI8UNrSgB9eyzP1RUnm2pHiwP0C
LTbxEdPdUWUNOD0XQ2QwLfkPaLv29YFyGVQc54o1dkxiC9vWmNaHr0V2gC9YMT6R
AJ/RC72XlKJPPB6uJhmEHJj6XmvpRt/l0xDu9+lnWr3heQx33SfuO3J3WB8VpMwr
stHO82SvT66n1xauYlDqZcaG2N07WzQ8Ldu+ccS7nGs=
`protect END_PROTECTED
