`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
nNeRV5ZvPd66ACnaDGjp5GULMYb+UWclsMdeNCVW1n5GWp9dJJBlWAqAn54GzmBm
Y4M5ENmXYYBmpKWQebf/1Fa7d/2P+VoD3PiK0S0PZQY4HidP1HOKHv9k5BkQpTOB
mrZNh2pf3JWfvgen16ogD+hw+w1+kLuKdWkIAw/4eVsHGPvmKOD/9uEis0pWu9hN
kYKWZk4MU+PNfdpH+VbrOROF9HI9Vlda5jTazLRCFkSc/dVP05TBwM7coSPRkUHf
`protect END_PROTECTED
