`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4xPbG1ja45eCyQ4wkuwapdEg51f1HiHcGqw9MH+ZfOJ04llq+hflvKzxZtueAGpD
eHy8+n5cO9gILeUw6hH5BjH/BqtCDk+8BvFT/qQd8ElS9Rkzw90ITUzwAHTsrBqB
khVYSdHU6L5wHoHgDpye6GNLAmIi43tga9YN9fJXW/9HkVpzqS/+Nx3py9bBxNmw
frba5OZeioZ1Pjhp2J3lG9rDHOM9mLmHoFWmmg9aayM284sd3dtXwYVljAK2/ik4
AoPNtmMdk0XMtEplx9B8vB2v7D33MNbkuYkYzi0r4WmKhj5T+r42iNyh8/iRG2I9
RZgZ4QSGTWXQXgYE24gy6jQzs/F6zgMILe5VwqgwLEbj7oOwxNQeFmfGlTJv18a0
iQs5ItEJVav9TCiDb9cmhpSQSOgMJoHaZV4T7cm9RpotV9kEK4gCclpSVDZjXeKt
wGAthBhPi7YvNl7jao0SIlDuMfh1CdComtawrflChIa5fo9Q3FLhz945Zf/YTms1
5Gf5Zvobgas80apvN47OsRnTjd3OGOXuGnKx8O3OZhLalvjSuVQ//1QNw993HOzM
J0NmxMyr5KwKDvUJBaHXnQ0MJBBwRGYVYSD3ugSilnto8BYNfbAn8UZgjzoXcL57
7TQUTDJwj+lMhfcrIDnhQxig7BV/64fwxC4BDGiAvwdgk2iPPiiZDdLvuu9pGUoi
6UJn/klKl1ENTpgY/CqvFuqlhZA4y2sMgfD9mjv39TYepqblF0cN2i0GFGzEgf7y
/3qD13GGA+d6vdXloORqlldIf/raBqg8kWTILf+/P5h8WNL3YuINkNG5aeDAELEa
1n2JQMqHuYxnhI/gNs6JAWr1kG+i8+RSP/krgLIaB4Dd678wcvQ1CZuoKvSEA9aT
6wlxWbFjXysPKb3Kxwrjh19PDxfCgOJpFr8yAeosgEmQgYIF0Xtu5t03LTpJJLlc
I2SmnVY5vCvGb0a+1DIKeL19sJQohgUv2boUtBgnLCZqd0NvAkALl6lA3jJSL9UZ
y/v4/7dsgEj9PGiL1/I5XA1rY9WAF07/h5v/T12CcAuG1RGxfY/Bf1iM9422LJQf
2YRVSSS7VTHbtJraqXNlg3Qscl3qcYNRyWqMNJKR734LzxhWdUhVrEMV/0dKKuen
u3WOQ9MwVFLgb20LMifBoQ9bmaBvjhoNoWe3rajsgIARvRBrTpJ+2wqwLnWs7Flg
y9xXuC9MJLkP+10vETT6XeZtHUoaFRF0tzkzEbt5ko3UncF0BGvp+0tLLiOHRvze
3cNACh/jIf612+cpXKtwS8T+kVUyeTFsVfcL/DTcxP/WBR7cFXXhEhgDwtx84pcB
2w5L3350HaexDZPXiBxI4tO0RTsmc3bUaK5OLWyoeFHc/i4Y+LBY4deo/8VcjBbC
16Sk65cfVXNTQoQSWiySZDV1qrZ23BAFg/SJbGgwAQaxJP7eOc/Ns2suGqdFqDGn
tFeagVfXec9RMj0uTov6Eq38vzcmqMGX6SOjAE6Y34/+eipiPIq3KL3WS1M58lIx
SmBCY+gw8+gLbI0sVBIYdKo0Gldkfu7iLjX5QXliJkXr2RrMg6zSlUGBPozr/2cW
PEo7zeDoRaHn3YCz0/23qK5vDYT7yqhtq+ldbHUWxGonof3NKScyWcgHDMiwE2WZ
zCIP0BSEsEOwtZ0IR4DqHI5XqcuYwjDTywrx0e36wnmvVrB83bYi1RhshJemSm/C
JNwuIvv3pfLJ85t7Lk+79Qr8RqORB42XyjrbyVlLczbJBTaOftxg4WycjJxdEghW
u53+aYE8zlRGY0Gzb25emn2Rre/88HDQHHxSot+dE/iEYoOaEZZ6gBHIMw8hqH/B
KaplYA8lR2yuMmW2KFtMenaNQ5CBgaktupkKOS8RwXr1NxiPEXjl0XnG4dUXIM75
F80J7nAluxpVc11aFtZgiE5mu/RQV3EwjXLGpJ6ba82FLKv0s8IMCW434WK+qKxe
tbV/cJ3pFRU0Yy/SHqBtREkJMgAdkR/KB+ncGA+qkL2OMxNyANr7lfrjCQ/HssHv
MHm0QUm9b/W0Lbw17MWU91rk+czefST+PTARC+uSO77cpwMOgaGXzIksd5hafHjl
Zky4Pabk0c3ogbT414kHXhGkQIcicC8HM+tV8l3Rq72SzyLc/2CYQj9n7W2mFE2r
42/84+cejthOdBqsRtpvODTJeK84dN3r0+JiPscb5wY6dbzWCqkbo9ZYJi/V7685
a+DjHCM1BuJQH6AqEf3dodQGnj9kbZESnmlH0t8ePczhfizjp8v/UFNmI9DmZrLX
rjxPmFz/kkl6HwWVjL4Po0ymtdDqfzcRaM7BaQWbW+ZMS2j313zMwtIcgscXj8OQ
JnsjZ2vcPHfQId7RCYdBt7enOZZa1Fer/36SMogrWx+B8vG5yemNvsLMz1htzClM
+9rylCzJ2J3FUWYrWFBRaC+7F/HdER8+GcNvfC0UicCMuy9teS4yZiFvuDpJwT9A
ameyZmzGM6UhhsxqwjKS9Ljb1kZcURBKiuoQ167ECXzGCDp/YMwQ2u+TkOHlDNG2
9bjPMf/YfR/QBFgHL71+Nb0OvkuI11S8NJJN9c518Kuk88lRRAXh6A1gAywRZtD5
Nf2lnPOATLUkeVXFD8XIZYixbQ3c9LYiYBcB7X65IL5E6aN9dpreshpwQSsPbTI6
rqUQQWs4blYGPzdT7U3d4C8kor/lG2WOz/OfnD6o86QQ2Yt8MSV8v/YXNPD1U9dx
EQA8shqL4FBvR4ecAxqsQzlOggxopX822NWJ9bimq1wP+05DAOg93kh8uUFJt8UB
CpHIV5DsuEP/ov11eSmFtGM6xZYMz2ZcNnHKJN8LsLe30CF3ZXsEjSSb0hEW+Qcv
BdekjaqQZhT3otV6olXYJquEXbTJGh8Q3CloNTBSoPbGh1Ak4zZCQchzdaoKEp31
Dlzd46iZTA0YtpXUuuKMPPJOANgRdl2JK2qWXB0yITPEFoiGJL0FdvdidZxX/CaN
a4HWsBkGcoCCBowRT4yp62eKWwn2hmjXkrSPoK0Qn2yzWxbucNLpWtk2xEStHwXW
4o2NWJNHUSuja3Ki35NNyUxOezzzd8qif/UfeWKQRm7lw+vSOMFNMaWVGZZNtAc9
HTi8teB4p2KuvEJqgUKgCl3OL6wPFLJQSLPjwvg0YB0E6yTMkHLKx4HBHRc4+ib2
FP2jQ5VddDIVPjZyAfdwdPsAg/SFKcxDYP77mPa8J35AlwdQKFrsbHZm36x3zZp+
i4M1JSNdEILoD8+wdixtPvdf33t+B563eCo5gm/3Uu2CEPSFO49aySUjTu3G51/1
W09xd1uKzIWbgByhDBf8cw==
`protect END_PROTECTED
