`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ClBGNQkz0yNQnoGY/jaxNDo6IkUqdX5ZUh9SouFDo+pVF/wC3QJseKGLgZUlg1bi
LQJNafOhvOe638HpND9bjYPcvIISYO7EAgvWBdJ6vMb8UpKNmU7NThs03RAaMWWe
7/HbQQ509wUSJJCCqvyHV2q/kdZrrzTe9n0NxXge1aWkxhkrqJ0F55CrdS/fdG5y
27//ZGYBgimFN8KjNdbJ/sOrU5Kd7qmkNwufDRiIk5fG4U6CmxvmercMUtJsO9y6
NHP359GSH7YMSg5DS4jn7ZtDl/e1RD4fxDvNeA4TVTD5cWwsA+CsT38xtuvi78MZ
fifktVJJNhohI97SronA3W30KzXwN/jxhdmzh0gDobeJh9vXkZ0SvQCeXm2E5zLX
7vc6gMupk+2vUkW8NSFNGGq6K//ZRa3JsdvzuNUt9vvm6sbZ8LlChN9Pm4hzfFQq
XUOwpvfPe4+VOwVDygWsdg7N185AZ6nHNNM98OJPxYbIBk9mz9TB2SBXMX4NNIne
0Y8YnyjatZG9bDOXurPQgiNOSFmC0oSNQCoBOXlxMx3BRcUP7U7olnecRSVMieYn
MgLXdimVm4Y61osKXiG3V4+pIBPfM+KuSag5cvPG135y4Mely5CQQgIXkjUDhAdB
aoR6YkcbjoTfVW9mSDeUrc3l/BCcJtu/kogVOBUuPC4UZGNK4A3Zm/mLf5exvFcy
i+iuLnJ+yEb6hNA5GHQbKi4wkbRulGJpExDpZXbkQGEaIBl2pvkOy0BbRI7QxhA4
YVYANCGKy++b/yvdvOmMz7DgOu7kcZ1ahOdXJ8D2AEFRkrBYbhNzkdhhk1b49pek
eD84QHE0zT7alS7O6SgpYtC57GYynBpzY8HXLiTQvcLT7D94TLrEkEonBHsqNRTL
6Wnht/dlXAzF3hgt57uiRe8Q9rLAPfLhJKgabj84oAp+pVojhToV5E/yWVeSDol2
iKiwP23NeYulK7LMjXW66EWcVHVUxOrnYxhJjdRvfiGFXdQuYZ5HMNI9jx3e5f0X
ZeKYUyRTuRBHHA0Zw5aqboIoNciMNjFEwPHEkIhWCTKTNV/jPIg15msMWpucE4gO
J4gcfsazGSS3sVi1EgWmO5k0LfTRlpOr2v4kDWgrQI2E7hrjtBYynjY6zhxyVwUQ
1eAt+mBgCEf4hCc5l2k782dwD0vJbFqlKaBNbFqjnettA59h6sUqEhD31YwjtrzG
45l7BS/ART6z1gMY6rnsIhEjcdprNgFk/NaGVOyx5lzxwGkj97E4YkPAcXA6szXr
Szz/vzi3WlSV1pZnMc9ATt5ZAZLEcKAaRuvpAUDHc0kiK/n3nv59ywTCIZLfUptN
ITsTwyi5vdcjGZ5d3LlXZGQbkdKDs3+g7SbJjbZ9/zKLVVVsUbrOwCpnGWBhQGyQ
+bd0YXGlbk7FIQ4neOWEMH+7rG6Y34DHpxSZmUqy037i4sT0ZoFuNNCrxR+4LZoi
GhyMBJsZlGRAFxB9LHSEUfLhrve9cDNbM0O5JZokSg8w8tZyY8AP8443FGx9kXMP
PU8m7wv9quydSYZX9h9z6u8wrT0TXSVmdvieRsuN0Ur7+3gvAH2an5Au9GwYRJ87
E9YW1m2tJA9iAXBdt9P15YPMntDgwE+O10tQYPRXkTr7xVMjLwPn90m2HAKvtrwe
gHzVlp1l12dRBFXe+ZtIXIoZ7HIKiQvcJW7kS5qbd5y+Xs3oFklX0wF5C3MUsqQN
TY2qwVXccZqkNfUc0A3sVnBhHMxrAZKOKfbQ+BhrOFdrXehZabLt0HAyj1qU+qmW
HREGPPEUd5L0FKIwUo/2axzEfpUqmS6uYE1v9O7TUek/xohErNdRYLMixCJ2WtDI
VviNsPiWL8GOGRfAlpV+gw==
`protect END_PROTECTED
