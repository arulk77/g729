`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJI6k/Dn7cT95g13r4XGmlE+2NjR6QmCWbFWqIRv8FGn
oJ8Z2LBIWpqEgmQOQX5kk8jQTvnBtU0wyAgvXUq4hqQFs1P5oAGoUuw+QsPsxu6E
54M1hVIPciB67PtuxF+oTGcEFwQaXM9jC5MwxfcODR1TtDXN6OqmAsHYX1E5Tf06
ylbExY3H8pUM9hdmLY2f7t5VgpBkGSNuPUaVWOFhp4YZzcRwpVVxRZrtDG1cFaN6
dfUPVBRQi+D9BWzBpYJt6Q90Enkf3s3S7Nj0xQwCUsKCcUx5Ibv6T1xKzP3fpM8j
jWOaM+HqiK9WqbRDYp7OmX6tJ7dRMmnmZLH27kQzekvaD8rbgiL973fwGn5OaTeq
EWmeCtVlb8Crv/Uo/zyGFbLQk2WOG3yeo22MWly1GuTMemsjWiP0rACCzpPeWTjs
LL3JbNgad+hBVIRJJdE7AYMAi3vOZaiKh/ZcF90rBEGJprh0HF8yUJliy0gjlL+e
rcdjawIeSXNhnqQqtz21uxW5Ugq/aV8bu+kKV29Kp5el3Yf86Aaz2cL1bpBmPfyb
g5VIG0E30wRUAjXCtFLdOOTfSn9qkL0OzgseN6l190N1gBMaRkvbiTph1BEVEqEG
sAAeDPi0scaf5L9LOIA9IbNaLckxFVqZ1pbN/q4HkVFO61D1Hl3xDYRtCj2+1t0f
IHoVos5lcL10U2pQqAda1lsXBqhd0Yg8f9re/JCPhjq3/jHAKnUjU8/T9mgN1LMY
xVMk9UWueWh1hUBdZf8EyhkckCTTSEOGxT30Jd6czAJvawcNlvYciYP1fGLQqp/8
4kh412tKk2V/XSOu/zG7zA3MYaRyZVoRm9/UfkYKvS5iTbmMwyK+O8UalPhPC1bT
qO4/VjhrW75S7rzhOEkN8YA43TqXIcUudoLgWe/1gMLC6+gYOfDpkIp7wergoiN0
7SZjABfn8w0VkTxGWS/Ko+CaGGnLNsrDXgZ0PJ2c1s76BQvE0ItDEkjAhrcch9G3
Cjk1rUHQLaiFsbdug9m5qyKlqDiGkm1pjXIpHmYIa1YfMHTSdlObJge39+VKOUrW
9Covh5joGa+qvwecgHz6QKQJqZca9ajzCwlPdlDQuD4dhmiEjlV7YF7HnFTEDXFw
w5HUGdT/FY26Xqv/oWoHuDsAKtFFTP2cyvOKR9nbbRj/FcqjTPnECAFyFVY5l0Lo
9p6eZo1/1qSzijp0z+Uy+4AIoqM1mYbi1LSiIsW5uxBb7R+uLQ83+10t/MG7sn6y
3i9zTP6Op7go7RFZ93AlPHx2juvUPgocDDUmgY0h2qLvlPWbj4p9H4RrlEbO2MZg
xfzd0mVOTHv5VqH9BDCXHvxzGKA5JuK8G+l/1zHXB4VOUoNuog6RP6sLERGdCzaW
8k1M2urySHSlQazU9wHa0ZXZnSkJ7ZKRqZMeogkLgtSRbt1tffKapZ8PxtqKSQB+
1szEBtYXQOLO8QGjWnSNsUKS2ZTZb/imAdjXnn7uktEC1/IGqh3s4tpH2VUvsfuN
Gne9Kstk8PmiGF0Ae919IPZE2fRX+kx4Srm6B36N3HVzF/Nl6pwnV02WvtnxwUIM
YSpqh+lLCRyI24bAMM703loU+Q8vlN49kdUrGudQqYqQpE9mylGKhxbYoa3JVj6r
tUrTA3Ngk7b/zFZd6ezuiBLZeS62JGG2yE/G3MQffzWr6YP4kORN9F5K6dFIGAHG
z/JiCsXCaL2xEzknrC+SDOY1deh4noeolEKsg01Sl8L2e3edhXbwQ4O62ddb7z8k
b0DrIwVdMsggZY+75eaR3eBqMxMdlj6aKmzSrKAnhpHveZVXB5m5ehpIVfEgiutI
ps3rD+UT7bY95vDz88kqr5wh4LQxm7AKfhZm0dPzRzleXH6drgndHRHQlbcq5uE3
7AkOP26xaNczTGamjXmKUPv+tXsHLPs/scXA02uIqbtss2VcUgSI8IAPFwmuK9p6
3yjmxVIgwyCEx+YU+2zlVYigJ4KFJ3FgJk9UtqBlpHbpwr0YGWHCBLKewMpZhu4K
kA4yEAL9kSWKOhehDbk1YnW/zJOkhqBwVXLnwcd4AyD8M90S9ZpYS/Uf/vG6vqFS
FtGb9zH8kJ1NzX/2Y1nVqthpFWXGQV/uCc2VCrf8hZ/3xh0hor/S9DRh0XnARZrm
ggSnaG4CfdF9K90SRyNcem75Eufsih9WQdskHeIDHoCBmsi+hKjjAEdEjzgH5TQT
k5+8bP4rb6lahsG3+KZHdfZVkUWCVeofx9TQHhuZBQqWOM42qsqUdqIrCnShLM+R
BFtF+Kqx9l8/ntVZemtUsnK1YyJjTvrJu1V1cDc4UF+h7q8H0vsNtPiKjO2TjBoh
Ytdcl36VicCNoigDTJWm+r4pcVMCkhYYr4/iqS09Y2wErKQiSJS3TvZomLWdMzeU
yhcOCfS59CjuJRsJqFWghIeUDJ9wpCWWZs5zJsz23A7r7khcTHAa/OWEKQAycFqg
UIbENIX15W0rDeZ5wDfgo567e05bVKFjaVOoI6XvtlzvuuCt+9/CP/u8AXMjgxQd
/reOnQJfwZONWpe09T66w/MO7j4XTFZor1H7zDM9D/eeSjdr0Zx7GBoDjehXaSLZ
TD/CoB/YtYfH9ggzFvE703YfcFA+IEBYw1S/Qp22PsiNBAj3evJlP0x9jj15Hke7
j37vtiaSNxPQqv+BAf63gw==
`protect END_PROTECTED
