`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN9tpU+ZsNkJl5+mpNxCzC2lcJkMy13Xkg1cJbG+WqUm
5np2l2nax+FgnVmBu7vxYBI5ubQ/ZVXnZHtvg/7T5tYzCrUC22Ao2XfoTlh9wD3u
I2j0tGJ5VlIM8AP4rV81vQpq7wDo7ePopNfMngURa9xyp/Qa07Wj79jy4MnIa1gr
O50molFiqwysrl1tUZhc9U5mn0Ix9Jr53dZDShc6xGOwESHJMHanExJnDVtevMJ7
BOIE8jvDz6hPs9yRRrMhUBVp0Soxsc8xrX65Q8dZTTgQdgoRt1A2XGAbnETmujYu
6Qw6XIg3BhpblxrMj1aR3Zgv4QpUENjZs58Yw+RSgk4hjX2qXTXYCxClDki0T6lD
NjUQetjojPaEbxBQVuKX8WCwmtDvMQhy2tvpzSvuHK9m+a9UzUT/5OE+sIiMy7K7
vzGcVJLY4sCjodwBDoJJXO+3pmt3mFbNF44EGDMsiDm3yKVg3APDw5dZSXyDCS9f
2FNMas4oVwhNaBV84H66vd9tLiGrnClqb3rcAZkS9/HHtGKKb1xYRnlRWnrC2RWK
`protect END_PROTECTED
