`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42NratkL1bsTULEQVLMW5+ra0GuCj3TDpCE5pDmumBPC
kgd5pY20aoP56ZOZhtzlNrr3Gz10hRb6IhSELkkkvZr+NtAtHdj5XGd9qlsNIV0J
uquYj25NNY6+n26dpc4yjum5pUhTdRFPeBB2WF6jXtDL9Mh9j5mc6h/v6/dRwK2x
a+0C2Pxzdt7TZX4QXq6mKa+CMVTJhg269TUwxafO0UVZsc3XLi3Zln1Zkhc9C8fD
jxtFNSPFu4l8vN4T2CMu45/E8t24S5bZD5d/hljW90G93HiFT4IM+FRahdP3AepH
5isKuIn31h7uHcnK4OYeDMfe3kG3yUkqmjJjpdAprN0O8/X1sOlpLQLprPf4tO5Q
pClMsiyAwGEsSSmV6sQ+MaV2HkxzauHczyL6oWkxCHEtwGf3aayL3Vd8Bg5cGTrf
sS98YLAO7UhcIxmaYrPxPg==
`protect END_PROTECTED
