`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C1CK4qNG3+gct3kcvLKGUoVawqS1+JdtbNoejpcDXW9E
PkLZLRL5+wDLps1ksZg7bLBZ2tZF11MbFyOOKWZXB8rx5mcI25vNi+mzFVcn99i/
V2RQM5YN00axQj0ukeRIsaDBPq7Q+iXIw6b7Lm+4QtIWZMFM61yIeV/XATS/a+3n
LKpKgj56c/SfFkKImxEpjViW7Z4i9oPv+NsYfA5fulWxgBVU8dY9y2JJttPf1vB8
GsNZ3PyOBXS7I4gxheyCFPP6lG2eYB4IvvjDaNKF7/BI3dJ8HJqC2oYOfABHecyn
J/UZm1TdxdhHHwGpujOd2Z344V3X7UsSDEA0Kv2JFpKMc2rSmsGVdyxRylX87axo
b/TrNwQoV6hoJMJSn/p6ST9jx7732Vvw1CZMINsfll3HuffIG8FofNCFwzf9AXuj
NW2Z7Q6ni72ArboK4E7J4UfLEclqn+b42+vLEe+rNCrHNIHsBeKSuxNjHeCUanYY
AYilX0uPxqDVw9HKope6D1aBFfF/VMYqGE4Cy7H0/UzK/4HT4oU/kBR4NhmAKoJx
81rh6HC47jGaw3xfZn/GH39k6/mPC9A532OoZKEI4yHHl3uITXI18MdoTee6JzlO
HKSXMcKMhGs3+KI13KJGBhW+KjQsmwNteRkFpI/bKwNVkgnRxXs0uiHLUm1xfi0w
38O+gHE55rLfXuD6KgxO3FUeVr5YtC7R8zGs1rXfPU0jmDGqRY0Ef1rSdvWNQGxb
WMHQzMSHCIhzUXlz1i7xH6GQmxDYHfZt34Ar41dNRmon8jRK+BjJzub2yXaibaoo
o9U+Yef1/UXoNPzl4e1qC8crCKGMNj3A37SuwwGGAq9bX1MWK0Q1nRL0rrfWcNda
IfUF0hZySyNozdfe2FMtFp7v3WlJ0kQ8aBwQEM9JnPzO1PLg9yGnVQUYBBrzVfEb
suxeiRLxW9Zz3E74OYPX1Ec9OTuGiqozr1QaBhEfd+u2Oukh/zOrId7wbIZYaSJs
srKcfb9nEXgcR7x1rw6A9pP5YjB44zj3MeKIv0LtFQaLb9VXSe3RsCAINreMXpDi
4aOyn9B7dxm9zKMuhrm2Vl7eLDZleg1ULgjlMvL6f2lNW/SVCHNG9Q0P2mHBCy2o
ewZdZN0pgct5gO7+Z04EWnSnFfNeR+skbYjCKlP+Exau56StjMv6nD1h0T8l/WWd
q3IHVg+hST7gM8oUlNmMi+GueIwXZO9jj2py7WRtaIV/mt23G3+1cdUZBUZIYN72
RU4g4T0/8IE8pv2ShyFyDno2o+LJiaHcLpQJJY7lFY5bcp2B00mDlZkAYTfPAWy1
yTKQifnuDiabYzBb1x1NoLY5DaFQHNYG5uyPaQMS9Zz5ATArgttVi9V2ZuYHruCj
mYoPI9ZZiYRsB8DdqM68502TyNkp4joZWZ+EzoUqwOSs/lqmaJiIjti3iCZDn7pK
Zm530ZzaZ2HBE3DE/SeXUoKcBQuRcBoz+BzG3eOQlMseZIMh93YqTo4khXLV6TrG
stTsPySMAYS+WAlIgBWHrQMF/gH892S4rD5ygjKkw848SS3la1Wb6zGZKIwr5/YL
ysE/IMwSZZJec+9NVZ3d4C50fNfCgkqfl21EakwXXCqpBLOt9UOHELC4mQddbThP
VhpmKAjzOHtCWMLqwi4A/W+SsnVldml6nULCWtAwEs7rUvZrd/ZsA2BbaA8ROsTP
/KYH8UhCmDozvQyG1brB4RRfWn3Ztz927NHcV26Zc7KvZLl5J3SGNRJwLyx/E9CW
OZzQB1S33xlSMvI6rGyR2xTncWZl5we8hTGl4EB9RpLZp4BDA2HQMD7+vwoecO6a
xxq4yyXFr2IpA/VhP2FahHEIYTMWOzWjkBZoGyVEFX2q9yRnBAYERoojXorzrKmW
pwUJxyUprzuo4YPtvkhQxHNygt7+y76rMYtRi+gU911sf+UdTkvrUcI7oMvmM4PV
/WLBN+gjd1YlsITAkgJlrBca5XBUHV6Ghzhq4CTcoSPRRSVQ8wUKB9YxzOsfeW/3
n5iHCNg+4zYaNlS2OR5ga5rsX8Q4OMu18Fn7hER1lfGgK3IgxeTPlvtPmsFPw1UB
JWXjtPOOIg56qbpiUF5oOHfaHTBmGHo10PxxgzbdClnUnTK7OTkpbQptulb6DaV6
EBVSjArHDUEbySTBbN1H4PvDWOkqBvVS2Rz5CYtfkIndOaX7/454I4mYjGCMySqf
2iTPcPCjAgus3lIFvQiWBanONEmj3p8plj4qdkfTTUma+RrRUE2FKBZzZgIZHVuB
6NLW+ZztZXUP5vHbK3O17gFZQ9O9MVgJ1zOm6je9nMC29yY/VC8obKhY5OidWvX/
sJjMxe+w9o2RyzZClIxSksHCkXb2PoZnqePNXbrRc7q0cLUALe/wpArMKrTvTba+
TUJ/JWjscQBmx3EtzaojnseN6iTiu3ClstR3e1s3AoZEbaPnqPJ5ojdl0mNZZqFb
eQdS9TCtSbt0YDMVXqwFIa0g3Cq1JQiVbsmUrlcKO4nQlOCRhVTIRnFJX4EcUZAu
gSvOw+47zlBj/E1NHOfj+V09rtZ2WrDfw+mKRNo9w+xbXo1dB11Vnn7fEFjQPBeM
ozXHo0VtlvfDuhXprhXPz43RAsnath6UNnc5Cgl1ZWCXrblBA9av+fk43MOC7gIc
60UyZNdUaMqLENaXlPZjeCWuDAno8FHVONbN6ILUIOYpMziCtCHWPyJk3fFPffId
6ZeACBErzVeOsf96mG6AbsVtqZieGvZtPRlym2EQ2YQpKIFyrk6bmxWzvmEvfdc4
dmwgFmIz1uOkueucgKVDOJqmxT97D6ONJk8FVAkRSzLgjmoqDpLHrSR+ce7khDYD
Hyn41PQPBsKPSn2RGKdMkZvJOG1pRaY9bv2GnoPak6SxE06r/sLxpY7mK5YVvKct
MYhlpKOvRlfiXZ5ZZzL7cHQyHk0bFqnl7JCVAPGrZaZ92LUuJ/WPGMsNEqUJOFjV
DGFgoIyHy7DLuNHO+L4/By+aONsd74dqlB47NJtcT3dpFqBY6HpBufVlfIuIaKwS
yUsZBzCMixkzMAR50Qen14oWau4qsBz/gCNpS3MgZbs1xiM8xKI/iLg14hGYZ4j1
igPBwjqOeKpkVqbdFoLxmQqXZ2WX20fvLJXex6eODMDbvmzal62OmU3IcH1u+vNp
54rwyyHKCbkNN7eK0DIttNa6U76C4c7OPFNNjZ2tHy//rIWPRAK7A5qucmAq2u23
ADQp1H0GnxOaqbcNLww6mFasqVu9WYR56N8fFqEzUjX0VVaot7vhLL/VoUstb3c5
gtZa+CVOg1lqqyGLpO3s7IY8/gN5peAuGsFwEVITGnZbZUdM2mPasgNNiiA0XJ7Z
UXBt5gSezn1YUi4Bir2zTi7XIvePDB7SdsBeHpCpyWpS/tm8giwNjizFNxc/XSjZ
vQzdKSa0txPqZIHXkhv0TvNCbiBidvljgwTp7TtgaTkjJ06pUWhz20HtOfvgRU+2
iGMvuF4m0eXyIQfzNbz3A1LNq2j/6UzaQ7yB9tvjsg39m/da7Yi7kmXnioaC0acs
0ygRuHA6Mje6xqh6JHw+AP7Mhbv4FKu38JsfEa5TUMmyhMOnNe05GG8d2YKSa8Hh
04Rh6OXonBhYYt+asrCQeRVj2c9Ccm6HNEAMt0wv4a2uA5/Z8PrJG8yF5nSFxxjJ
gJM90KQ+MyKcEfgKu+6+pj5w14J07pHpI0RQ+EwTA+hg0n8Zj8uzzHE8xBMSyJ/l
xKPoIslCrtbuh5KZ94/ZF8sprNuSh9RFD7yLEmzfL93ftNsOLPFaOFspgdZ+Y23C
RNB5boAOHON57A2+YXnziJZYnT2wI7VxeJ25oyEaXpN03XCg+5zeLQcSyw7Swd6N
4QRxsdPDOPwO2cYoiQ30nGeH7sTVjzpPzsZ2I+UNT1Lm469/eounagdYBny2FzRJ
+XMCX3+bFbZq6XUf5427lzr6uWOmKzIedjTnwmS2w993Z05ekRnmVVhNK2opaL6A
9g7BQcmaPY8y3OUtKrSoo4tyZ056yqVni2ci2jl02hJHFHeC/6XQ2TDbB6vSpw36
2QTysfEBoL7riBbAwSy7TW11rgJRPuSdHszdVQAlVky2qh7D2sgKJikLVXGFynVU
vRCny9bplRv2bAqsULJhSRpd6Ea7EzOYFHVStYUg3OANR76XLSpiGeapQCBtAQsE
vK4WZORAYe57kESC/4zzsW7CtVHl0r99emlmfveWV4uWHvmFqg9JgEBKmQJBYxH3
Adex9uEeiE4GQpmkYGeWgswZAVqADDkJ5hFQxrj0Bnx/qctA/ugJ9BsqA5HQdtNt
GUpL5FowatM4FcxzI9A2oLagJOYoa3v2WTZg9K62QkG2qQXtFMApxv/2EpQULQQ1
/0iVccWS1AcshEfS7CuKHwB2QBP+t0tdoRUA1FgfoMbSWyTZhoJwBrwKCzhyN+qq
gKi+zHkzJfWJnsiqdSImwcx1rM611oDrIvhm9TY00WqQLcdAZq+FFFzFPhtTNxvZ
g9WM7f5111QiUrF0S58KGmrogdTWhF1moGvcoplNkhz+0LKHl3KLRmmbd9h8zZCR
wnf+TCgKRsR03Ds7Jxygqe28LsIWoR9gq9UGrClW+a3sooXSvq5I81JGKTeaqkzA
kAPs6kMq0MqpHvU/iv1SWZH3vCEq4PhUTU9c8cCxE2kobqpnqIgwMxOHGdpvluou
5+SPd8VQoertFe8bDUnjURElb0Wi9P2A42HndzTtTgNCj9fXql6Hdm5n2J0xdRdO
23aT0n26gQdzhlRVA6SQeQ4sqOQR/0WWtYWjtBDhNPfLq7cXsjKs3ImDTU2DCDBr
BgUOtosmljBbIkzqDAkENXCAPnPb6ZcPbwDyJU1NhcKBqtKqZ0b/7bUL+VWs09A/
BAEywPuJly5vQUgY5xZXBJVthn3+Wr7pLNxfrwo4KJvbJd2n17mWYUBU7MS31lng
6XIvy4OhlEjVERn7kCOQMxOLqvmzbgETbw2VktmY1IjNTfeqa8Eb99wmNYbMyN01
5nF1Any7sOcDrNVsN2UsAysomZkvHBKM73icKWOPJh2nCGb8Y69z6Fi0KHO03UPC
yTYx5fTa3XPkcoQzd8iXebbLJBZ7vwil7+9Z+vpUJ9oUpMnyHFGVb/W4ERveC2lM
14lBtd9g6ls5oKKhF7bvMa0EYwVlTVrFULe6PX9B+nGIdPqN8BSnznCwco7PmFjO
a8TJ16aiGWVAhCnCOkygdbvjRzUSzgrMEXw64cth3wsfGq4LVv4STLRfTev1mFNc
W7orTEml4qtz1l0B8M7i5MScr9gH5d4/C2v5X6SrYGhGAOXXJQX8ohrEiW3/hPLV
nNgjAJo0yrig30h6SzYGgveiOqBfiJSnRrWhkReNsmyN6WeC2QSTAmV1jDjdlUVr
`protect END_PROTECTED
