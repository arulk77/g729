`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
RbTCskhYw8kb6iz+PJ0VOMgump5mG9ZM1xkrOPbPvgeBeYVwMixqk4MVEE3owfLa
hvahuHmpvwZO8sywhy0r6z6YmkMip7//n68RgcKt8bYBZignX1xW2ayCim/fMCm1
7PJX7Z+i/FPKKvOqMJE/otTQQPuLO+5OB2o+sesT7eya/iew7lLlpGkds8q28H0W
ga3VdEDJgGJS9rRwZwtzf6FQFXIfPXaI1SiCH/jyxReB0tS1xCmczG72VYGA2pIE
ewNV5EqsMC5t6cpyIjeMNSbvgZ37tFDkaFpXkEHP7bDkC6AJonHjdgYik5vOQkna
u13ij6l2tnUw/A/xAlT+NsK66afpEnqzEH0x2YayX18Oz6DLxoBqiPJmIMdXHhzH
luELGG/dDRtDyslcef9yjtmJNUx88pELoz5OOrVKajI=
`protect END_PROTECTED
