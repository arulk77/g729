`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aOI2aYMu81xSDl2v7OLppablYO+JNZbIVXLhalM2UBpAm373xyNxfvPVe39gC8MN
68q7tTNlk4cXmcGdiQzYDKZuZQZuwgCJGSgg/CuGCprpL27/tvyJTDTgPw276kza
Eu2Ss4iqocEd7xFeUGOk09IJKNAKXLWiYcwBsfbv80py+NDN4sQKAg7dhNdu7yVa
TAf7r+nRAMI4IZOk7FrhaoxEsHtqRXC2OFLJlu8QWR+uHtdWsowGBxvHxNoLTfoy
kBIoDG242C3HW0u5GxgrBuwf/pK/sht1ICIkE7kdZuIKfWVmWzfHuO2hYwknXehW
saxWs2SYg9is352RexCelq3nr7RqMYQ4wzQ3rBBtzLkA1zxDTc+3x16lZE9lp8I2
41sMKKZMg2RQD36kLO67vJk0owNlMYwowCfyV45xZMdFCOg/efmIv5h5t2/HAb6M
t7ZBm2mfhWqiT59aHiF52bTi5AzevlxQCQTJN7tJpl0=
`protect END_PROTECTED
