`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
yr0iEjEQTJ7ZS2CiBX66B63t/ZOXFlbfKZoB9AQUui7+8HIvzSOlReln9ySxqgag
LsRBCUXQhF0uwNooa7on4k3OOEj6/eqRYbUCi2RcQe6LSUpOqDQzOmB0ChRQZZvH
L3Zi1Hof1SY4U+C7zLt/s3Hif9GvAS8MbLa+d+gRi2oQQDFQ3MnLgR0I0yWoWgp6
JYTKdN1HQ9PjfCZPrsVZhHZ6EfD9DCt8w++lX5N7sod8Hjr6/0Uql8z2Jq0U0dmt
YMLiE2Vne6d63EJk1RV+yELXI1rNqz9vQ3XUlaw7Io/to1WpAY7FfkgihtfYUhkU
SRwPd0b6ge/1/glfz9Aa46Xq0gYpxXibllIfaNpRW8n4HzKCqnGYf1VNBffd3gGL
u6/uS78m3kab0g0e1FjCthBTl43VT68vJBMZof8XLPQ=
`protect END_PROTECTED
