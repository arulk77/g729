`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48/PQ03R5XMWN//yd8L854OpIrOeSeEc63QSeTM8aUPj
gVG5R9Xalk8kV0SnmLRJR/oF5LPvoNdYNrK8eT9zXutIuMNLpVRxWpmUooxB3/l3
wJstV2Ttd/8/C1Sda7lRtt8sq3lZnNIsKVf//5O8FqpdXQF26VBzsMV0ZSgGnLDa
hSoIW2SUqFdK6EehNZRst3Tw/BLJISbMAn3XWp+kisCAfr+Ac2ln58MWjC7wpW/W
HogHOoET2WvursJRQNp6SJzB2PLyha34QrtMh3+wmOQGVi01SE39WqqVZf78WfA5
DmX5UodNxOD1C/zLiX5If03qXRcGghdUWMAHUPXzEr82SyqXGWm/bnDhUYeWZDt5
I9r36nUnj5wKOL0Fp6FEW30KUWTfkSy3UIDhqYcTM71cp86QmQvAnscNv2H5bxkE
pXV1PYbIT7zO8d7TUsOjYHYutE8DK6keotcYUA3XgjPGAnlBLk+wAeGFvE/iBaOv
eVWEIe3ZhKbrKc6GPswkPF155P6Sj5yloqspXyIAfPABWL0pt144s3B2/nF5lfS1
C/lUeCsPU0yl7vfC6sHNJO0oze82vDjq7qpoYOfE7Bc9Oe/Eqzt3MSwU+Fhbi2kp
UK0s91KRkqNTtc306IxpIsgyqGvauiCJzz2b5T8O+UywSJH0fZQSF64RGBlaENiY
cv8epy71HHe8DsqKfPxTGOwiJ2l1gm/URXkrKiiN4bYaQ5r/mogJLQFbidCuq7Ek
4vIod09FT3AazDKlH1AsTpHKq13yTNUGVJw0pDP7e5SSMr3AIWnKutDlTHzfbK7V
scEdbjj0dwYI2EJTGNjylxadQNNsSQkH65DEDimF41KIMFgUdXaaO+N/4u11nkwv
Fg6dGAcChI5zhVzVSS+SUpGmFS0Bhid4NTFDfN392whDwcjpd4VHPDhWnD5cKrcB
tT9xKnEx0NezmMNjtjiTesa46fyAtaWrIUL+Noy6K45BLs4uQSjFItPkEOvEbenB
HKvi2cXWDgbRAHvNuyCbOdfHzkphpMWcSBwqszcrjunR/d9rL/NFQLh/pdm2XozO
/FTGXdy0Sn+oTaqnON13FVfXaPeVK4F4wqthtqnZ2DTtBDoKgCvfMzg3C/gVYKKh
HNL9IZlXq/VRQqfHw4YG82/pdA6Oo3w9BIhCxNCN6V0M9BUtY9E83HyeyHs7QIny
D5+NvzZWnBu2Rk9vtZn/13DvIFRFAsOPVkOUhmnkPBUnX8OQYva4FNlLreArqBKk
IYOLVK6LzEEV4LxwNb2m8jOrwyb8+6UbLGe28GhHlMnbiixOy0SQQCZuS18dft29
wcaCknn4AfGwQJgciBkyraEN/4ex/LnO0LnzPQqkorQ2z9nbWRwy32qDWNwRSqry
p5+qZImt7r62UVUSvlgEr/FhC4lolTeMF301NJdRi+drTaX/3fY0ITh78BFBTYvU
r67BLztJ3SEbbq8C5APPSFJu49DAEcatBxVo+22zWEgYpdLBEqbKxaXSGx8NOovH
0tzn4KVbJqIVWOmaf7sFDEaNqHSkvrf64rHlOPjcnk7iYHOT3dKtIaT+vgqSe97k
/sjJePx70m2omuU5AoIYiXPa+WZNzA3ObaLSavlPv+UF7XAqddb+nb5BEAOCwnDl
MNZ9BWDfhPpNnUcvfe+ewAlhAdlF3YCpTCRwZtoN42c=
`protect END_PROTECTED
