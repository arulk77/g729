`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48OYHZF7aaOz7p3zAF1CH+hlFAfKMecTXUDcEVRtI3lp
+dLnBee3tSUyhjK9pmOCIKfLPBvdN86VVBJkNG/AWwA0ORG9COAFJhG/c5o1VpiF
fvz9YZEXlOcESeDznGRLQpYLz1GlnAg/eyFETtSRlstzk2pECr4iI1eFMdBV9rVP
875UYnVhu3SJIUqoAgIvPKvRkg9j7q7a6E40Kug9t6HUty/MUZlkeQrd/YRABNpV
cQBoycD2G9e6I19wNaKulJ05HSsAW7Txxa7+2QvYqbAMRArTa0qun0WMd08Z2hiy
DX58Z9G6UPWgRnEAuMc/Kg==
`protect END_PROTECTED
