`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QfoId/zzuDxLO/XrIPvQEw4MEnk+UzCzzzI9bDlhSbvRbL9TpT66Y2Mj+r9GPsMj
t6kXKDwp7DvHqFgY7J35vrk+7rkSVfz5KQSz1yy4QZ5XfHuuH8z5VedS9M89ZZxA
n/Sy9k39bjuX97rSwZb5sOYtGHbc5GPMeeWVCNYa8pBxBXGCNf9Uyb4V6VY3jZfy
E3EDUcPgwakBqBpK+F3UoPnK4kERWeJlvN4T367cY1CqlNU3700YioLEwP/4tvHY
BVzD91pO2vDifcruX4i0wI/ATpj8Ych28H0xbTLkd6K01LdSrS6je1aEAjqpAs8S
`protect END_PROTECTED
