`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C1c6mRI5Qm7DGMAI7dOGq56Dd7Q4kgM7ypRnsA6P/vs9
UqYeNUmwJNOz08fINqlOar5yKI58CPmAJB2S4VS6wUhInW5IzL5A+RPuZk5lYS+C
++4MYl7U1otoHo/1ywTvqrHGWNHWHEIrnW38OM+mwmVrPUrnquNGqa6hZ1H34ykP
Hpoujpxh0oX2QdU845Uz67vFeGyWPr48pJlLckebYtI6Dw6hRzBLdvVLbyXh2i31
uvAAMlO377Gs1QBdu4wnRc0Urri9+YcgH5EpD9fU5CulA6esVeRbVHsnZWeQ/CPL
7vsHljtF77a6la78fDHXy+5tlC+oITRtbRGI8OHSnE8OeRFw90p95rtT7Ud4sIvK
cjlwMpad5v4ZDFoyUBpLjzxRngUR3+vLfu7697H27divxZHJmwxaWlnRNqcQXlqs
bSYXcqiMN1xPtf1dmi95K4ofmSgUwT1mIbZ5wWorVO3WdieaJ4WXTo8BLchR+6oy
DMiqnujuFaGlYRYisftblmxfoqsd3LUTpaFSOujGY8w6aFP/mg+tbjoAkP0oRdGK
CsPl2QO+1cS1LyQtdv5heMPoOuQiwLkMbPpOSxignk141diM6EMtjAYDspcEZkhR
DC+VRGN6Fjuw1SzlLUNmqCEWyJ2jntb5tTGqj1PcxqbJ+uGWuus44h/bqBxUitVY
789mIvI4kULkO4T+AlgTf6q9sFiMaptZ5V5qbu90OoyH/bMoDJicPeHeE8yUMuXe
j47od/3cWgZ5O85RyXyMtByvkM49j7nhhr22cCfr/mmtYqL7WHFvkVQqT5tUmm7i
wtFd4yBCweD3QwUzSEzn0WjunEh5jER1aTOMR2YCBmIPMEyRhlVHREDOaw2PKJLd
5pgwN9bNe1TIreDJeQP42lh/aih3JXLQqR8QwtkQS24lkKxc8lCNxRQ1CbWcKtxu
w3qjeYTvXE78yGDPJemSWi7dSZStMY0k+rLgZiGGS46OW2ClE+3CsatCODSE+Mbf
rvO7BYEboYMmLGcQGUye45QPVwQv5d++ooQ9jDG35DIRCduzBnvMTGfTWuiwyvXJ
2yN0yaZgdM89YCeGobli9uEilBgUmli9Y+p3LPvIUtqJUJ7wZni3xKz3Pep+ENVR
jLP+qnTJJ9lP3C6yXqyRTE+mto5EPpyojNtOa43BgOLG8HSx3uaB8m7fVCV4q8H0
kRMqs6vUI0kItAJoZMYFF+Jw0+XO4qJh3/tyJ/nJ1bb3PXgQhSSNEQgIui1Cufuy
0ZQMpToeCYyg89r+1iNMOVLEZat60qwoLqdICDvVeA/Gw5XsBSKeGP2Yz4Uo2KlG
b1rAqosdViimgUo8A1wuQUS9fV2Mo9E7rJiRkDsLYHoteFxo1mqxyr3AMuaGKQ77
nJo50HH9ll1/l0Vl5iHwnr/mfBcBatCVI5nJXTnXT29dXjGLRddGyrGyDSYk1Xrd
4qE0LQuxdWmT8aRMmrdpRcFsbxrmhaNXGnpLmwID39vr566Hr0bVhn4Fulj7bYPF
Xkd33gf0GSHX3mpvRU0xqIPz12DivdUH2QXS+iZKGvVtArNO6j0ay8/K7+JG455b
kLNU+yylEiKAnts3cKAjg/K0AQAZsDCtH4HdkY5cr5WhMbK6X5jq5MLgE15jsox5
cw78F+Scrib2WPeUkBGvHdlWqtgbm/sD5etlg3bYW9VH6i6mw15kwNyms8kRL4H/
5S6DnH2z6dzz15OdZNIlQ5pJTJ9XyVC9wCAY/6uHqwkPWicou7IwqnBKEbdwIXs+
qbilt8Jadl2DDGt3EmXjJC7FMAZt3LOHebzuJhpshT4KapqB1T0qUs9DZ9ZW6NQZ
NPtqV4mj8o5bg4ObHktBPy329yiwH9NwaVO2BiERxsLwtJuRdS7zhu+jUezw7tvy
qI29c0+TowpOw4xat3Rikqhe3dE8xz6v7+AYcNymw1gURuf0BjahKtgle1j0oKXN
vvSgMpIHJbwR8KoXLuvdrw3MCEFoeTCYqlmVjRTw9/k67mKjXTRH8aPlJo+D18yA
ntTNsJPT+84xRxjE8szURWXX1EMwzEU19EH47CbrrgxUy6PHa9oB2WMte5227QeS
KvZ90d2AW+Rc6S135L1BGYB9woJUFihhZ4K0DCFWv6nuqOJMW/JC3S+JsRsq5+gH
6hJ5xl+WkTciVq1CHp4oqPaVbbNpLyriCeVB7Z46Ug8LFcYySF4zEMqHezx7I6V/
/B2/p9EcOy91Mcs5NpJjIHeei9w2LWFrR+wNUPISFM3LJDc9UTAZNa+Rcbf2cP5V
gPVdGErQgHAGlkWePUHGgzRgR3adTug5dm2p62cejyNG0/+BE5imjv7ucFyo5jYc
HZNE0KhXiq2RqEF5j4fqFvERhRNvrhDOhXIH176m4lLUtamv7ffZ49Tp+xQKLlhY
vg58JQc3asHCJgzirZZ2J8GUcGUbvxCrriFvkZgUFOx4BHpFD7NTQ2x6F5jruzeM
rP4GOZlTM8tftezAtmyBhrdQhAsofATpC+l+f9scW7+5MGXLY2Pa3EYx3J7VyH//
humTAMqTuwH0TkRYLCekIAlG1EC/BLKcVwgDiX2SIu4eYbkeUhd/9minG9M+QRmn
nRohXn1CE15arqKLFup44xMMMGGmTFdSrYSu7OOm0TNwscLtJo576S84sa3KRwHe
PmdGHaP8uZsIXvQtqRpWh/u6sxQ/rmD1jm0V3SBtjzzsZInwarUiAh5M5AX+nync
I2VUzyUvbkaz1A2K2i8XMymc2orVqDUxvzW9VISup2+Zm6c2SxtXiErPJ5xJ5giC
D8ggqfBHnrlCgJ4chzJYf3sJPjgqzAJxZcImwVg7Xq6lKgHDQwuN3v+jA0vxAbA9
WWHOKD3H8uIHzLFyXiAcV5iLqxi10hdixvX/Fgw/pHnnyYi9IX9c1hpSN4CzSc49
amxlOxBgWUNGRqVS6WOxWGuV7RHd3nlZfVUEVIKsjDhr+fSsj+vp1p5CfVavfTKu
u+BdfPqYmc0tiDR25iuiSNNYl5HGUyWkZlA0e20F/xlA7mJqIy+HIaseFS6W6zC1
aonVc01swrm4K26AvYb6A3Diy3A95dJvuVLP4FZzioI58Iv1+pzCzSeaD9sA1KP7
N5ZdeLdHLAEQeNImdVHld/c7eJkabQrcf5o5fmZ0Blt3Kdoiopvyoj08vcf1Abt3
b4NVBh9QuTfsv5eVmKboep7SLI/umvi9RZSXQdst8U48ToR4qGwlBFNMLXxYo7sN
qRZMthFhsHmR5SG07KBcxRvtB4Xrx+/UZXAdhCnj+3GDN3QZ1MR6NAjmIv5O3qGI
RnMtaFPC0X9IrtimpxT5rTC67vakasXTWdZ6u5AyW7hIVeLcculix+oglRrDtloe
+x+a4Lqat0DsSUhASFbr+RXuIRmACi5sxKw+un+49cLDOo82sB7n1EYaVRrcVKo5
ZjSDbS6CNR5nFXCJkk7JUyqIE3LtjIystkIy1ITrgu3ArR21GA984ZkaAj+luXzG
AowfGqusiCCjLyIN/KhqrKk7zdx9KaK8LjeLlTBFh8nCixE9KEprUlAsqS/qL1Em
EGGcSFR6BaFIL5KdoX87xaOXUYm51N9IeUaX1VmJrqCGiABGGHYq+FZcrvjG3+2U
7DSGlx6IFR/jam081GrMvVvPxWj8jpt6dDvuHFwa+Wjp3tdAU15f79UPvTDDdkhy
DpKS5SdmbbAYkDDFcdzu0PKZrctXWkOyyqLe29b2T8EuzW64JV0ZIqJ3sJol3UQc
sKWR6olCVcwvTTMUZKlqK56D2CBaccI+tvecqkWeFCvh/34OF3oitBIHoOWkKmK4
kuUPBaaxwegWMvxkorrwXhQtwGnj0LlvHtva1CYthbBlrByVV5RjNtG0cUyH4Z3t
rzoJmxNb6K6Zi6DefXhTsd/8/ReD4pQwbVqtPQkE4CpoPdn+9zT39zrCYAe7k1t4
/orR5M6YtI9Gq7El3Zr7KWHB2fgwCW+8A+rvoQtVT3dvxfdE15lBSY2akRScqbFk
R12r/n6Ken7RjBhEwU64KrEXOeRhJ3ISUXReDfAeEpAMJ/Nk2rfaPcCYkjkHN5MS
evSSy8tSj6A2fbVGF3TAQSV3nN4/T0rt+X7hL5y8K28t0MozAqSBdIjXtNyy0dAI
rAqPuMIiGNU1KtdUxBFy30Mma8jvYZKJJWvPDkmeUL2Xp1sL5u2Z00cGmhkTVI85
PRM7vBhNPpudnGBIsSaAEoiZjj4dKRnWFk74EgVe79t0C6GFV2XzC1uFCt0mn7p6
tJCdlYe0aX9iOMeYzHsHaMqpxq9BODjmf391pL+Wco9m6YsPqaHxRydPAOsihKLK
qAUDyK9HRy4H9jLNy4Mxk8wKGnwzZ+8YnwufzKmGulQMZB0ljO+JQ/1PiQwoi632
uWP3qrIrsMhWp9KedbNsuN8fnVVInNN6O+g4425ub72P2EOscF/fDqc1GKHy2/ce
XbppGBGmDSvNL3dzdMn+T4Bj4wzjFBxuGn6ySiPOegTVU8A+4MIMSx8GED2LeWWh
c0L1S4uY+G0LoVLnCv9Ji6/zcKZsMtkzbhV3c2GRDS2k3eGA30ujB8dIFGZUG34i
RIby1Y3ubgD3e/pqAyZ96Qj8YjeVi2G3TE2BhLVuviGrF54g2mu8szIx8z1yeEhd
DmZDrQq+p+qH3tfKQ9TBN2O+J4kQcX7uq/Pce8GI9KbbZqyYhwhzIBHepzrcdqZD
bmac5Z7iUDk4HPT6xIJFzMHmjJ9q6ct4roZdGP7tPkIYXn/OnkI1Q0NRsW5eAOny
pdVtPitaSb/YKOrQ44t2R1TlK0N8HB2c7r0jwdXAHQFp3iz2zfExoe7m55daFk+z
jTpzvltsjsPW4fMch9MC7TZN8Fw84pfkf8TlVGtyswRcmPoSNlUeL6JIZTOd7BAI
g3mH8LLvcOCMrQCRwS+odOgcQbQncI9IT07BWJruzoUd1O2DI4PBsLeU2YlI48YC
87iD0TbTRAQ9EHUYtXRzcP4tu+e4obBPAG74Xe+Hl1qDC1l7C0mBV4dqHBCOCb2H
iH6jAYLE2o9qNN6VZtS9XBtXQ/VvOPo3YPrm/2jg68okvQq/x+uOS7zCP8fO40R0
Wa8i41ufA/zcORqKLMioiZkcehXVURZdUj86mEOGeN7YvFBSRNl1z04PzMEM04S/
dpi62pFPtEIZ+L7lflFDBpYi8vx/eojPYSr9ZwPwksHEK3qH3iLwORK6k4QahNh5
hGyE1KJGD4eIas5WGIx+sfnTVFxsr9xYxVPq5jgNo1vRymqSArU5GL3X0EdttUWc
GY0XX0ZKXxZx4lTtON1AdJeu5H1AZg9Ha90eNDnWkMVbmA36k23Ng3TSMRn+pIbL
9CM8GxBwV8KPCAxE2Kpkqlu8VlfRt+Nof8TrrE5vGAzWz7btUXQOre7LO2vjbrUx
uX4H8258i4pURelYKo/DLmKNg0sHQWoxuYjnEpZ1cDjfLrWTBnZ27P/KUEg90bdl
046ZWGxt7R89NRjjNnqbPtMqxrb4ApCGOmjNLsTwPpetMPO4r7kOUSNuLG6QIVMJ
7sjuP58GD4lJIEH2W6Ieb+taskUCNax4WeL86ouP6tufudtJf5KzMqqMUQJGGYSJ
vR5+ZwuWCn/yA39LjTEPKPaMSDEFFRbTYQIE1tYxRq5ybsqrKkFfqUhZiW8P45BJ
r462e+dwIm1SSUGTsusgKs5aJCR4qUjJ2WXC1WPiVdH7RMmsaK0LO9wIKHia/d9w
jA0oWm1brMF6Q9vIQeDee4O5DSyHuBa5+VL177QAOm7hperQ05uj89lfAAKiWvoR
5BTSPpN2Rq3YxH3E6hnndq5TYSBSA8nAa/95Uw7ML+1Ja/ajscuLQ22Lx0LN/DK9
2+2t9KCBGOok4cApxyw/B/7KM0rVMft2+mDD7erbqnt9Lxf3lHS8EHIZukoCjPqb
MX5KNkdLhOSSZNaNEjyJKUv1SkzzGIP+p2ZEyAJpEIZl45gtQTOxilRh8M20YQXT
cLoh4fHrCJOv9gmiufyadqwGyoEWLNg6g+++L3YT6nIXXemygGTuccItVTnPwzGz
Q5Sc/KCNpVSH+bS6FRfSdVw6M+hUst3y/DrCwwzhd5NOn7BWc/6TKTk2OmRezQS8
I3wMi1+4/N5Pn5ZZXcaI7f8nKf2GyuMfJvgKWM58FkkGWPNuADHdkN32P3S93trK
d62lgAARWdK6hhHgc3twagUlaOcfD0LBPHmTofcsZC/gh3H8HBUPne9pz5cn86Pa
UkRxjkTa9IoJWbNZbntS3tcLwTbRvoGgjxKMDccxIniZ7IZ56rnJ1IxElfBhZIgC
KkeYYYzTEQ0ck3n3y0ULppBin2CbGj/H9NKbGfNQG+N6W6IENiIYDD8yQgZlTNmK
6Mw3EEws3zA6XeIy2u2OqrXV0CbT3su8SMSowFZa+SRY0mJR4BQlWco0vYjFmG5Z
ifZ+yEuLkHhuVjMkCC6um+gd6H7V8fg1jl4X1ZvWHIYpJ9yK3dlBgtGh+4Zt259y
oPjbkcqC1i14WzgvFo5UyvbWvrehvR8ep61alOBgv+XHp4PxFcOQOf9LhOCpH9EP
rdlcX1H4/J4Yf0eaIbLRTC2HClUMlhGfN0e92Fbh4NcXkIt3fZQl8K3r7nvARFLy
TcoC3QVQfF9FGDXAJb6r6til+WgmvRVUpsGZ66fFyDbRsSaBb22aHqHBrMiD8Y1U
C/IfWK9YTmYM05BgQDrV6/0QBshN4lUL/CuIb/mxI3uHFYdHXATGCuGWUhW325Ie
V8uHFRU2Duuk/fQBfJAzyNbZYYuH10yxW54mTC5m1nBlbnt9GDkZ+r61wtIfq8+f
X9K8Blbp8wr9TnPt921QpCeAtlhOjokiBCwrlNfep32wMrgraizx8KBeSlS03/vg
o3sqHroonX9XTJHXc9vemk2Njuq1PeAhSShDHdmupzp0tNtajtAsxy2soeKcIcmy
6ggQ5am4ZY53jTfu0aBDf0C3ZoC+9bR/1MKHefN5IUmsrN/Lxlcit7nv3WkbeXH4
qjyhlpCCZcvuEWueRqgDJMLRSUvl6vG1UbE7UEYVjUnv6OATP/F87pRsEARzxXh4
jGp2wEgFs7xL/hle+plFNyvbQrFLsArIclEHBNMj7Ajl8kgZpKjQdwCyLYzo/lV1
IgsNNJ3c5M8AoaqDITBAVO/bgfoX7uXvXjJv66XvrtSxlKtCNgTZUvFFWopLlSbb
ZJterTgR75s0frZdVR44TTl03Hquas5aR0aQA/bhrqKLcNvLn7T1jsXmo4SZ5F/E
idnnQWXPU5Vy0O+08pxPV3d7ev9oplL5Qdot8L08Fyc8D9/+ty/05SfjWIbB2Q/P
20LZpRPiSaNkyWwq27Tbtpl17H8V85/W9Rj3vVT+LhKTxYOPM0lcEpINV0GLdLDg
TBDjJLC6afNKSOneuwIPbhG8GLDUJcQzWMSY1wZ8Z6vFnLeRr88ryXROl2IP1NHz
0gQ5VVqWhFd6ePb5O+nFnbWfOmPEiHGOmiXivHg1EGjdICoTg6n/9VnmeVFa5+1U
zeGZuhyw2xiYpGbehInvynk/4BOJ7lATd0LA7+0EuTQ8OtS1wpVnTgN8Z5XW3K+M
tpewd8t46Xj8+FVy8iBfr9ELMrLpiJ4dVDbNBktRVA/ESRcgYhiDkoHwN25XdEyB
RJeAI/2V2Zs2yKYWEkqH/b8i+4lPGsazLczE1g7RkYfqtZ0mCySQLWis1SZg43Vf
rjG4QeUwvQh9haMfPs4hrq/zWnSk0H5V9hMXN22Wlek57bNP4160uc839w+z07P2
miLOR+9giHLlhnLYUCp414IElbEG5t1MSUCKn9DZ/3sLmJJHs9uml7sUle3FY3uE
o2j7YnmyBgmtvsmtq2qW6Gux+sWmMln09eIc2p+xLm2z5SUN5izAR8AQG2GAlMlH
2nsBQbcvsit+Z8yMOMzlBo60ORpu9RkXJCCZTSIHekmNSeNHn1GUMhgSVbS5RpdQ
LzTDmBwHL3aijyJG9Y/vTJCAvS3pWmzOXKdk/CnkfB0oMXeumqyp2IMYTCnC7hMj
iAjeZBPjSRFbJ0KQ1dkWqCD8kNXKJhAL0jJKhxidNJTEMYcf5Rt19DDGEE1V+riN
mDeTx6rZMLq7gAWARpAPDo29Ldlpagi+dBgv2UJZj4TCbOXx8g/krdIyTdD0lbrD
rXDeM6p1X158HnFRWKFoeh0srSz9iJu5uqcC3oVDnzqR1ESa9t5WOWdsbp7CLnmE
TgN+JXAJSdgfdyJtgkDXm1c7+dg1MJnMnciW/XT/GKahWVNLnbQaD6QRUvdHa3dV
eRWQa28i5Ht2MUxdCJW8++c84La3IqymXBKVKViuLnHyg8jK+703dZQrkO8f3ImH
sxnnKTHoSWNVhxWQCE2oHFYA3Csgncc/4aV984Lt+0WJGDJTv0kUU0s7yILruJ1g
xLrO9gB8GFYWiSYAd1MZu5ueNLubUWu/SqvSbKq8UnwkM7E1VlQqUQKssHuADskv
W7WgwMIQoIwqBXXTE4cOcBDZvNlRRZEmLMbvecncQS0Mf5k2oVW176yFYwf4L2vV
7EetT750uDlD0ohkkoe9/OYim+TBEww5hMxDqznnGkVgiT3bfwy/kVTtOYsWgRBy
dsgI9OLf6yRHgBEzxa/+PXHkhtrdNW8Fv7DJm0Z7UXRirzA5GmAspFMnOshElY38
IzRDwx5JUD7xibz5GovIfnfL0Aa2EZoVXEbBDr/D0nxPfS8NvQZKD6yQ6oAFTp4S
JHE4agk7OmLAoNcuWDu0O6HtDkNXlP19VfdytYXeYTx0GFQ6LEZD0iCL11MjZY/l
0dDsSd732VfbBwusvzY7J0kTc5FSriGE6utKlghQZvpUW+aDlsRqQSBDlHcaz7te
yH8asU5k95M6L/wlsdmdsOKOMRHW49tpco1x8ehbo5JbyjPnAL/MVTD5Zy9N0nTe
gxE4svGXqvHm8a6rztF3qr00ohPUrNEEMRepRCuW7AyoDNWl/opyqc36MyE04XZ4
/s9zhvDkMBtZkzptQxkA30t3XEZTPi0SJxkTpMUaL0Pd7n4AdkSSAuQsPwA2K6wF
e49nNqUyhzuhSSy4zlcY/L2nALs8w+nYhrrN7Z92DChhuEohlKoLukH8nfafusuS
rtssjqjJ5TqAaW2lBjbGY8WxPm/XV8KLdzXzXppEtOmnQGdihuLMQD5WTX4dk3Og
+pdtPUXs1D1Sy16sovFhbpXtN4952f28AKfJTVl1DeZ7Q5SINcQxu7IPA+nzHFLm
orE+1Co7/Ee//fUQJYi+CQ9RtBC74VItOouKTdH/oRrOmnNVEfQViY7NDvMiGIsy
NEOYDhgkN+OARr2oVSNNk37ZkMzh5L86xHHbo5dflc7RYO2tEkXrfKG9QgUKqWDz
6EtzoaKRyLj4c/0QIZaULFa1jfHmabBzdA0p+X1qnrFr11GiGuzUTlShJSG77Ehp
CuGFnl3cOAjyNez/bTuY4nbEIejANFcKrYx+p3AXn+mdInObbZYdGxQG1PualQhP
Y265FPeTN0LHF99/2D4vTCezoDttivdpQeEWem8HJvcIj4eeV2wq7Y/VeIWRe/ap
e5dXNo+hx2JgSznnVXFbB1BIlFAk4xiwIGdH6Dhmq4ABJYYm06y+3UeZVVTkbGY8
vJD25aDSQGrOlKymICc+A5IQFnjxnuXLiv3hPzqz1UObkjdqsNrMN6UEEzqTSWKI
Dks/0O+NImuTCixWHpEeWDma6cFyYvrLOUDyIufv7n5NH183bGCS/cdLlzJ5QCTd
O+D3lKvgobWrwtaR+HeUSG6W5Jtxhw1F+sCyrReqDGFLPjTxKPxELcOptp6FChk3
Ln/mkpIanjzm8yPfxoZSY+IRvSfiEw5bH1SGAwix7kftKFc4BUIv6huhtZ2LqQ9u
iXxuGndJ1U+qFejZXuBZFEapPc3DFM/XINQCGKgROMCkuG6YbfoMFGgbkw0KHntm
M4DSSU0hClVulvliV/0bBoat+P/ZAt/HjwG9KRLQCaRKVn4sMCcgSJxJGhYf2uG8
4HYFtBKlMKDBePttSvmhx1G455ngkQNZqIYWWF7lzURnU1w8sAxnRpErL2qudJbc
nsNpLRH2bo0k5pfT/M1SDkSy9V10KO7MR0NzXvoFa4F6B7Hg9tyxkKF95g2SrdYT
sYO1QagqFEpK0e/LSGhQtUFUiZ0eqh32YGiUhfeBXURPTTARKT/qMqnrbhEnGYLI
eYtG/HFQn5qnlkg8HsUBc740K1V7wQpboz4hmy/LkFRyRsz83sy/rng7skTOQJhI
zF5S4bvQv+g1LDNztXgTElzNe78nf05xn3H9QUgyOC1j5vhy3L9dzOkhPcN3pXZP
zuKzs5VWoAzBE2wQ/eKQJCyZx/Cg8lJbyuUPdy8/WvP7IO+BqbId2bQgYsq66WUo
xMKTXzrDDBjvSvBQMjle+yrrlHm6eiPD91d8IexOKCZVOmjuh6aUc5bqFVYop7CO
NPLsHo1wQ6ejdgtjn/CPHb+qxLkk1SB26daCD5JZXzmXA2oQGj/r7Q0D9ewUF5ms
rU5SAdmx8rHJsAOoCxX0MkWb4/XaBC++BBh3jbX/2L1tFtPAcFmaFUFIvH4yaTGK
Bay3xfmiOJODhKOE/yWtNO+/k5OV23tSBnMMrz6KVKuZJJORBX9XfveOmB9aZSbG
0cGt2AcQ8iRYizTQgYJTHn7Y5FFaLrzqb4SrXQ2BanMysQElodG6w5zMcQutdeo9
NvgOpU2neix5CHyj2OUipBi/UWCsnhaGYJJCQtq5CrUNop4ahGzBoqVTa2+NjWat
Jq4QIave/hcHGZZ9vXn0eGL1jhoL0QQ8oKIehFhxFede+txGPC/8eUJ4VPbubRSI
chscm5Uql6SHtCvNHdGSoPr2KVa4499SbqdofhSk9gX6uqjwBu/sDrfoDAU6kVO7
1y6q6WRxXH8FMBmQ52axh30xsYmv1MvtTX5TExm4RxxBX1w/MrEeM6mSmyGQswlj
ihc/DWpkEnMPXwZMmahw/w9ORLF9w+qlLDFmjBa0Nud1gAmjJMj1QiN/1QMwk0H9
3/386zVtP/qmq16c8hZX813tQhzS1lrMSu6FFssCE+GloPsSbZUdrR/BjtDpz/O5
r7WP3uVi0MLKeG0clpu2i7mtwnORlp8+6lT/I5SkPabpRaHdJBBMCbNbLniKMxYQ
YmbyMBs/9D69pS2jyYoV0M9U5VIW86leDRVM1gVlI84XIjrnIVxHzGh4c1TSHICX
MIYEqUoi/ri3WXGqCIKJG1GuKdQw6Z41FRmWqQzA9i/3DBs7McoAT9SoA6PSGl+r
jRTwluRje4y020z1fOgTI7IHcwcSvi4SGzJDbR/TquAvJbkfB7QcXhesynn+DxGT
3L6tdmX4m/kNreOto4riLEiEhzkVqD0VYAR/b96P8nGdNGAHOy+xurwjjsgbajgj
aNBmJK1MpXiu5XHlPq5VyMdNhhcdzKX2i/Q54YdxT9XYM1Sk4hou64dvGXHDt3BW
g+d0zJ6lk21JaVs7j+gUab9zowt8qLBwkhlU4Zkpuo+KBZjTXSU1yszSn+F2hBTr
9OCgwoZgPQi2Yk7PEGnPxq7wnKdAwXdQFrE43QTb7sTk1Awr7RwLsIh40V1viSvB
hnkKJz74e1CgKDpv1LnYDcAjAu3LS/xe33618phZuE+58RKSEARtDjUB37hSDSRl
u+ucw0xSgZnP7+ojPBi7kGsASQp8L1LuAcW9r370clSfL3PB88R3D6na/fDBxP3o
ML7YlbWCoJRu3iFT4tshrIzE3cATH5qTNSEbGY/DMjh2uTBg7KV+Emr5fizUUDZL
UYUMIJ1RuKbyV8ryNz+uBfaBCPv/t1+yhsfcIOAyW6j8sXcQzi2m/u1q/i91r9p2
JGX1tK7U2gZ5x0UJBAPs9YTEWntQs8bgm+Ba9TwqFe4U7e26G34pbghOKhjOUHW1
IPhhPpMUGDx9dIaNQ0dEJKS1L1wfDhKjUQ7c34rZPODFQXDhuvt4riEeMfLE/+UU
0ef4CUMgqafeDZAxZFqJCgZC0ZiaoF0OXKkqzGt6IfIO4ydzePTBPLY7+AfrHytv
LpZ04O/I318XheUaetO0N1HSrafDHjeodvr4c5IJ3PuXRLwqPsoh9OvONOm6XTS5
dYCF1fh7znV0FNd14cfvAiKlTHXEFHUcJ3mqbK2Mx3IcYHtZ/AHwPFO+NTBXYxPo
SDkdpBcD0/sqG+yPjcHIXt3NR7me8GCsRzDLrxoTnwoE8AakUa1uu6eW9FhTQPCq
qLfoUITSKhfrhSQrKZwMyq1WTGqUj6+IrGwooObSCY0cPBglwRyGMJhcIU29SIPi
E9X7M+RiAOVVjVPAieibz2TaCPzyLOia9P+Ux4+mS00K5U8ALphq+qP2RaxS3G8x
JksnCV1y4oJHsEq4eMxWALX+OixfET4NDNivhQBNjoD8xfjAN6bvmt3kMlPtf7QZ
4+EpPukqoBFxTCT5j0nkSTSSoIP6zelweqwxuxMwjSR8xpLqQQTbRK3DoaNXZfLa
2+VpSDZVL/6lgTo4PGkoe3IUouM/WGaSV+uEMJMab+2G/wIryRA6hnvLYBPVcyfu
Fx3tMH4ZZAUEbQPsRZ0l7zVwfcCj4rJigTJ2Uu5h5PoddrtlfHY0ALpVB52RvHEU
0Tp6k1Y805kP4Ldvsqj0LtN2aZ0bqE1lKPMVGZyQqbEOAIFAm11J85g2NPMnKgKq
mCaWhEu2Aw0BjBn5EJhDsken5eZrNQ8/TV8/RxgH5EhBVqfcT8QAtow9eINBp8Bz
gB94sOrRVNC6gn2ptSny1CQ9GMVPEHTSXzE8+Kmx9t5MKAhkzAIyczhBbVVQF5X6
Vph8B6MixbWyRt4jCBya8P9yLRdfuG8vcn3hzgQ1TjQAKOHurlL6qqgX/sN+V0nZ
phOZtgko1WlytBpMDf9jkDsCluIc63oBX+C3wxexTteWRFGYHfDvLW/KJdJ7qN5e
aavlZ42rB7oRBIEtzrWaXSFtekQL2wecv51MD6y2b3Qxbp83kV2QebqjMErY84Uh
Gj5pL/2o0HrQGapEcwBVxbnZQ1oMzHGgLufosGvteyyFcy6CYNN9bDdF0ZsblKRL
OufpSZPGouUCX1QSfxv2MUvnT1oYPbnWsMHXhbFb/gOBut8HMVFocB867JjYFMj2
G02Isrj4Fxh+YxeKTvb4jAuDyG9RHiowF5unmlFdKCjNjYKQY+2lVmwcsm7bEESV
wi4nAgygLrKaJ6W6gW4uoXlsdvkPLRBpqR2VIjcVScqaF20xmBdx4ZiM271k2gDW
EXD0oWNlBeH7gKaUslpKb1lMv0jRr+iGYTCxpuklVGdC9M7ApGlvG3CRE6S9eOT7
tCxy8YnBrt6YSNC8b7etw582mPbNRD+XvzVY2GJtx2oqfqf6U8SK9S8T/D4eXEwA
476GSDEiyEDyMqqVVYG/lgef0AuUqpxsKvI2z3gqdPoD1nbsq5JZQr/Kypu86msa
LQRCHuv5/Y0proTVBG8YmwCXNZIcJ+DCdNn5/XiT5lLL1S7QR/Vzs5pW2w5sT3wt
FIiCDoSsBPweKPBZ9ffRJCOwkl8dquCnDC9iGIKt8/wGGM+wV1+koP6hbOohy9kY
LB/lv1KZF64tZCxkLmErzKimIyR6duljmLEH5RWO08kUTg3pmpodJDqUGTAT7Vkp
gkBzJjIA0KE0wLtSilJFkEAEvXYpPAXulFIu+0AgkkgP8dRJw+K5S5mqlDjjBMgW
aOkR4lwIYEpGWX5JuP/f7pfMwhZsIWyAot/mPwafs8N9E/EzUvtV8pO442fL4muu
J3J5002kaQkYhRKYVTpDvVo1uWj8xoSh4zrpaDGgrFFh9QsO5v7unsU4eycZojR6
TxmoXzlROyn5Ymq61TeexGBthKw5TX+re55pmjV6/Jf4GlOvXJC058VKQ7Y/jjo7
4YESA02W38YQ8XDpnbyXpe0O4hmDxxMGbVpTj+6rq9N8SIMlfOTS7pRaXvtO/Jfy
SnIDgUJg2I704RcUvoaSuZEmXYNJ9DmlNe+n+NyVbzTdk6Qd+93IkxEhl6KdRSco
OxPtv8r9BC126LEcEyEKj/oAxo0/oS9UPKL+nXEqhMObKq8M5xhXjrKEbF9HRy+Y
Eb5Hnmge0IYYq65cUoPwGnkZEreJyROP2wfIN9LfVfXvGXgpFmgz/eDZSJsOMKuH
yA088ciaTvxnzz6v/+erizVM2TF42KbK8TkFkiqydoF6KJEb4Zy+DVs7rarSa0Ch
nMoVukgPtB6CvH8pb9FtIrCsHdmEOsiz8QASxO3LHZwzbSfaTyr+c1B195JTTmTc
o0OkY8pvYy6Lwoc3qD/F3hkiRdmnrtbJ6c+1MDcfSQZWwDanIHjd2c7sIc7x3kR1
djtp12ve1EVcVXVTiJrOtAbaAwXwOrtYMtzW/TP+umDjWFM8rNYcm2nRoeyYBOb8
EE4mTvHKzsMbXAegdL1agIPTB/i9+EDOo0/0TQcMl/wumJTgSTbzfXsTd1pXer+W
kbpdyYS7n0sJVO+oxD7ifsGGgaEyxfO2NCEXZv3Ttx9o5B125t+KlHbD0NkM2uLV
OFEbT10aPW70Vt1gJsKm/lss4xQmbjLjGq7JVJts4/9XzWG7RhdWwtJv+bhHHclZ
jiTqlyszEfZQFiSZ6YkiWF4kSuR+cTHGp9e+ike8BcEJtndK75P66L+Kyh1cjg+h
tRoDBFpha32afVk4rj05xu7kAwKi7yC0F40xvtRfkPIRUqUoRUlZpm2Ywmjp5811
xgJEG2auhIoIzbEkApK4ksPj/tmJPDmskX8V+NoOcF4wY40MhZZZDpKE08pOIWGj
c1KCAC7EuFM5lm1JfWmbVv+zCWDHOpgPSsHTI0QnTEc7mmD2F3Aeo8XpFecIpkjR
edH8Ep89bAFEIKuWnTfIYWWyesX++M2+e7Hntn+vlC2EeJnPJiBPV3xP9O/CK1FT
ht1Mes+Kj5yDDN9aXtX70l2F8FulcYpugAJ+pDy0gvtTDzFggFX8znab4kfJhQKM
5/dsa3IidAlx1Wehat3w30ADRjD/9jX54KfUf8kNcTKb01thiFQrEL8lTLg5qUHr
BQYQXwQ+QHKRTErs2vIc0St0O+3daP44QJPCMXjDOP0jMC7gn03ZOZnE/dJo4fsZ
9Nevqr2PvIWJ9WZdskuw5TO+Z+d/GExFxZMsAHUikkVuDl3HxYDyWdXj3Xyd3avQ
flixc+N0Ia4jYE/CJGVsk8JuWKYmPixKx5X2uUtT10DbiD6Y4iBHglSGq6Vc0N4j
yMZ6M8xMRDuo5fxmuEYIW/2S3kv3d8JAEd1InXX6NByn2x4rhl/h/FoeGmuqvv3G
QYDlEAIMlzzo1cTa3qPyepotjLe/2dUcPjJvwN93lrxc3rHVSddCKvXHYqrAj8K4
/RZWd36utH9Qh55oJtl0ldlLCbKyH3Yx10Ub0e9feB5OWVRTQ8CUu4H10y+C8xa5
yWjF4nGdZa6aTV/MXFRDBsyhc6VxZvpVkRISl/LVVcjGrEVc+Y+C9t7KHQzuZQzw
MpyvIVB+ZjWALZaBlAiECoQ9+UzVE00OEr/UBX/p+kpZlqDRYP1niMILf8p95d/X
bxJBzwBCgLYCEROnE5nLuTomiojrWm5XIrAwAC2+RgXW1Py41tKCzVxalG2VWMEG
nlUPR3kB8xkKzU3E0tBqlPaGgV47pMNgg7ayrCJ+XgvM2Znm5leQ7H5v0Vu2doRm
sSvkQcP4uB0vK/IYcJaxBDnM+UhJaKkYQ128nCOlotqB07hNV3+Gr479tKL8zX5x
7woxcbus2pdWxexB+HuJtEtOhasdCxaVI/EsQ6C55K9PzMK6KYtkS0REr9CB1W0f
DVT8hr1DpwDcYCW56CsmzWvYlMgwvteXi6U+JuCBwtSde+1go8Fyo0AYOd0wiEwi
Kmp/NO5EQJLcoHY7wRQ5dKpeeNXckTbQ6u4uAA/UhbPZoaB4jCPZ7uIWyxkMq504
N9tcCl93gRxEIZAjXpwujND0Pqqj+f+xQx0ZfpMS2Jb1In8mgd3vhh63OgffCbVC
0qqc6MC+XtRERvjwpf9W24oEQfd9IMtWKUAf2jrnv4Ov8Hzd7xcdtNhKjxrEADtl
L9zz++57qoV66Ux/filX/lQShO7h0NoUMZdv214cFPEirzXL/KEmedc+7CmXgWdv
WIh34lKue754bb/m3Ird2Wm90EVeAVH92k/MhmyVGKl05z2lpJKAW5TbwLI80XOI
tv9NZJuD1PCLt3OcweuPMtGuCCkef/ebHh/utAptFJW5kD6u9bmaGr0ZCN5bB1bv
Ij80jIPUi0rb03cNXcZQJzxGnuOF8UT4asVdgYWry6uzWZWsmqGepZUnsGS5RJHR
ZWV5X895TN6LrVJu+ScIWDMID1bW0HiwLoMbzzEW7oglC/nqp0ovr0Erl6VpAdIQ
CD7ps6Oj55BafOvsWfH8YQzseyMTps4zJaiRVqirFYiURb5J/3UK6s49HxeQAGr0
NhL5ziQeSwQVwjiNGK80YlZC6CiPDbc0BUiKl+0O281dlUj7h0nLhB3AnmIgKDWW
2YJ1oHoH95ia9CNsQ/+5kSjC2wfJHhG5TRJuy2J44P+Ry36z5lvKU8H5LXBzlocb
qUTfNcWRpM2mqtUKGXhfV6MHQAWweadpyf/2EBROUhvT+Va3neVzTZS52vnlDA3c
gAQjb79Kp5AmM7kFtf6RqRp9zncKCFfQqWGDp83btZJCSz8Ixq91NkCgAg1WUeEO
Yiky8P8w2kNkWy+B7M9nyZiusL2iW0q5xN8QptwmVmKTjAgHxxrEnRwsBwwfY9go
M5E61JwIjH2QsNdn3m/pRarkJ/CtX/lgX34XXT8s7d326B6MOEobtjEaqiKqwerA
AAkIpH87RiQssC+Ev6IwOuLLWIG9HamcyBl9obpLa6Q2JVJqRnmNDh6zUkrTm3pD
sJaqSWU6D0Li5dxlBU+Ot7P9nBFuHKwSis8nCYpXIcBszPNAkcG632C8MXNbVOy6
W+0dzQUOKRcUZgOm9GqYzKKVHRq+OwmTjWSpV4zLaSBmOoR7UE+D8QkF01SrXqNS
RRfVcUq4Z23hNvXRDWQevo8Jc45x/jaUZ4mzEs6IlcRdvqLkQoE6VVamhTosn83z
ix499xxfiCCOBWFFpnGdUk2ayyO5JUPUB0jC5lq1buY9wKHZFYL7voD3RAc+d+35
VustHgErLB6n1zRQMtJWy376YI/GtfTs3S+MxsYXUP27Kj+SHKBh1d4WgnQ2jteR
m9jM6AWEw+Fa1n2xNy38Smnh5cpLLIrpkwUNNUMqryavl3a3I7gvYhIw8ivCNI4O
/PeE2okrmaCuK0LxqhecI/qeQJ4Fzcds+5QSRLTwpR2z+EVQHBGk2hnoN+E1zIRk
FH9QGIjvvvErOcAQdF7QU9J4cDLqa+1lW8pSo5XOCRtubOktjMj7+zqIdCKaP3D1
TtftKv1k4WCyOjAIFdAW8Nr4AmMx6/G0NZIKFFw5u0mP9LGb6wGg6dlLsM/Q/I4H
xOMYH9c8bASxQHQI21DivU/P6rOlaBeFt+2J2RuTyAcEKqgrkBDLaEIZu33tVvfH
mD7rfWKnUIvfTFw2B8E5B1ZOxZZY2PIDX8YNP/+M6LbESiSWhMxVFiLuE5f19lbs
i8MeeMNuxBF+zCaU9dpXQeXR4Cps7yZEXCXYbkaA7ZpJDUIhrABlySl2dHrzmOeo
yXoENbPUciJx+hZLMb16fbjAnz3kvZjQ2Yos5W1alPpoZhnoRACV4DcEK2L+PGax
TUVPEzyIS9IVoJjcpRfhsIL2Byb3CNNQuEZDddco+380MIFQ+R2HFN1y9Awqe2NC
LkDQuFvS8debHQm/2AZgw+g/HLo7ZKmBfkSzObaaNkCyM1msX+7e+BqUauGZVhQQ
Ai2E0lhQTTrk4KRuPxzmFeO1gLf9M7tkcjdSB7iLqXW6ddHlhrEwq46HoZF+4Xkx
QzxaHv6mrF+KCtdl1AeP2PZTJSnE+wg+rBp5YYxfMaaRCyJh0hQUE5HjODLkIgJL
795Ud7xWzG7DQCo3rb0LEiZRNBomgm32ysOYduPw/lsa6bI3Wf0OTSRUmTKwuxda
p6w04PI/6fe4KnJI/78YgbZw8Q/2SKFpJAzmWftSlx8AZ/5RXx5/F5sWTY03Bcwi
05tOtHAl/qCS1h1d50W4TAujPDXwSc08OcGyCKbMx6exirakdEt8QCGeDu9yG960
lwrUHpia/qhCISaJaDd6u/DvIZlOH9rlRR5a93I3824wCHC3t7tI/qbILigU8AUp
YnX3UKkIEA0rRlWVLNqKW7055N2fIWD1Wf4XeAyRZWCajxOjNVd01LqWM28HeT5y
RmcCC79L6ovKIoj01q8+l+mUdQSac4YcWLW2x9zsNsafM2bPe2GLBEItm0SFaaiu
XJfPIr8yAKOTi3CjYfWGzy7l7GPffOfMeGmuO/XfxU0ZrPdm9IrDKej6vkPx7E27
quAbUEdzPh8mHjDggT7Gh8FAh4fYejdfZqy6T7G+s+n1BhCfFi8g+fX1W6xAkbqe
LM2BOGOrgvsFdm1e4MpnFmGXvQlGFfQffg9wHYuezXiYBwRAuZzY1oP02jZktfN8
7PxUHMBrhOanmxGn8kPCMO8HBybgc5heLVA2SLDRP8mo77clcddvQeaEltBEgJTd
dp/efecyuWSEFWsPwE+aRZCUZ/LS7dJ7bGKtVJlZz6FZR3dFeV7yFljWOvrPT9mP
AKm5lYYR2mP3TfcbBt5AB0pUFRq3uqXI083Pn/a870tylObbUfS+lBNI9Ydq6AAJ
+InIaOhgcO7aNzbvB4GBdo47AT3L08XfeC/lgSrxLBvNEzGeFf9xpyc8pxy9jbxZ
o/CrhAmEv3BNZMtsFTH++CdsmsfTxzHb3PWi04XjKEBDpjkSAj0Xpau8tpu9/piZ
bTRsGg1+pRGsTgHvNz1NWizho804UVclj/CzQwImHFMf57acw1Z4YrTMqYdT2/9c
TLTAm6AR/HjJIAcE0X1NpXs4wlWZLL2Nsuc6JEuEgfqTnJY8rTckLZJ67qHpfwbR
+DP0J4mqYb5kxiGyHtiW+FE7xGXlOdHnMJRzvKBVFSBp7aN5vUVZ7ktLxp0qXkCi
SOuDg/IoWCfLx4nHnv5/gdnrD0yQrmrqbU8AgxIYL5uyeU7qem/goG/Qm8p0gLdF
h8bvsaMaMDiLvsa1S28jqpHTNegv1MP1GSHaUx14gHKZMZzRGQiKTPfeakCiR2CB
QqF0EaVowYRZMd38O455BbtIsTwRqLZDPa+tEqaivCYzasEp7jSAd9gYTPaVjL+O
UwDm5xfIhpwe4gNacm0IOPAKVytVaPFaoCvl+qedvCG9yKsMXHpUKDcnAvGn200n
jUroUZA24jcNk/ZQ0NE0/G7I4f8EIt2L89U6MtfkFaVzum1SD32GBzhZYBhoX1Et
9Sy4vZ77C2trTVmhBhlPEd8MCS+/LlIKuZr67oliw5CxTxHPL6IJcvMAkZSlarJT
I1nk4kvGujEF0kY0dKFN2/NHcsa7jK/FbyNdiheZFdFpFEgBHHH3QX+A2vKNJ1mD
7PwHhKvuEA9iwkod1n/HT4viBNT4I6Sgc2mBlTimi68tBVxYndPybxDf6NhQvxCR
VrS525O5fAmPLGnCosnjgY+xOm6fif3jn1QzPeniLkbw66nnsUIMkIypLTs9HlKY
qLFvnBC46K5KixS2PTCGWSEnU+3CYvzka40oPe+rr91/lzcVPh0qy2v6IPnBk1m4
/WtWnb5mwmduScMzRKtGO9YZkWd/47Hy8ZzvxbAJBpZorW5p2H+6FDXEkbnvaqDP
zO5Ld5+plNC0SsGyAYHuoNJXptJgoiCU8uTZtUm2QoNQ83KOXcv4gAG1mYlvc7yG
vnwptJ58NR+sV7yxwVzwBBNi87TkuTvgfDcNgdgd4st+g5t23uGM3hrGKl+p54tj
tvDxepS7K6qh79NdZVr3YT0R1YMcrA+jScnUvWWnxz979AtE2IVSCeznE4oHaaKA
2S/acn4FDNA3hGxPW0PWYVbMNQN0WVLuVnjCzRZ8m7iYZq5M37DlqTlS/V48JT6F
iKWMfoI3bNZaPdf5a+lILUB6kYXBT2rLhs6PFvSyFr3FGJnbbWkW2DxjISVBPpeT
VXfzfIXvsgUHyw+4oBS20/6BpVR4L9oCBni5o2oZ5W3dq/eQOeMrPug8OctNSmSP
cXuBUMrBGBYCqyJ27zTPnpdppaHJqXyd8JB5JPBOYzLs+OvAixrb+ppVNZ3wxnhJ
S2nj+tiiH4YwDsUN1HApVf6wMPF5RXBYdOWCPt7O0iYsaRViR9bSfNL0UNq//lP6
C9RufoFccrsgRXRkJhZfB2KIDlPudLpiXP/zhY7e59Fuhei9eO3QwCKM+s+rAC22
EEtuug15uRG83Vm+ZoRxE/CTdlXcx7C1vGDrxFXDAdWXYO+igv+c6yMLItBcq4iY
koev5WZIWeh1421UQqIffvM4usxOyOvTAYMBdFaN/iid83TLi30pZNC/l/7h9+mP
mJsewwkxl+RtHUxzSJp3eiJmIQiMqsCl0tiStmZ4bnDlBHqeSgBzioy/EhriTSu/
w2ZmPz/GEIkwe66aYycVWOnL7DylugqyWkjGAdtb3M77hW/YCclffD3XbxzUf8S+
t6Abdurk6Iw0S5lroYhOfVPBOiiqzYjXmY3TkeBWZAmPdEc6zLtYxb+UIsltUXCG
xe+4Xot69CEVV4vIBNEclXgowqxtR4ySaa/zpoFiYNOa4CY4pdpeEmdvHmPdfGTb
sOzgQINaKR7uBDf6+3C5OL5kK+SUrW6670u7L5s3ebsseB3z18G4CNCrWUohU6k4
I4ct1NBnM8RpcWo4s0FS5sDbhy2yzWz4vxpZEYs1cqiKSJSXHSH9MO0h7cd0pVhW
N5Xw6cxKD4exp9Ki5/S6O1g+Ob++SVa77SIJ3Tpdv7Qb3iIN7vs4RIYrbBbzIRnr
d2wMxJm9a7EH0fqWKCydw4Tv/bVb2ZeF8/1GY54bYANaU75HwjBI6RLZKExpY3FL
1AIy6riq336+8O9Z6lJ/5TWNELaeuQvFdKa3v+h7KRam6n9ZEQxGBkvDjESVn5PS
9rXToZqbt5oXOpnyeobwZ8izzxqwPwNOzzXb+tE316EWkB6jWRhguiNZT+tH8vyr
eROHOKFP1PTvSNEH7R++9wlRr2re/9GYh2B+Jp8cLe9iC544GWraBPo4vB6hhpQD
kJGlnKwtnEMDIIke0Zb3FvcmRpTYog2m7TxswWsVGE81UebT738sdzozIS4mAVib
uWCq9UoNZIE7H3ahuHirUtijxDmTPKu5Iy0QV5YUNjtVQ0UuhHSL3WcRmOlepIzP
avv0TI4B4lQCu7FZa4O3efwQJ9GywNW0lpFurvsC2N1XHaUaqCq91nJ1rwMy0JvW
kghzHdmHRvdj7IqcqyKbGP5cX8iHnyRVRLXKMJ1VWQnnSVwW1B01O0eALKPvycNk
g9omM+zQdn6FWty7yvdxS/Bbut7TBK3lVXuoKqgDATAqTV9mW9XPNlPKqXe8+vNj
C1/16zEk0cIzjt2zyxEOjaRN4Z7G0WAeqMUoHFiAPCCQ10iMOwaiwYieSZHy0+JY
VUcTPyFt54Gzp/Ln9o5QrwvWoaHyhfJ/erCBw/NEmN/2FE/9r0Ge2epFExhAHypr
q+LuguV2EDjhEbfJGjeyBLXyXZZ0JtGiOMzPjto6CbYv2KTdtBciRF9nEiBdQGht
THP7m8m6R1PJr+phBLtsFnhAEL5qxB7jPhAuoX/fBWhQF0vwhoBCuTEOAtmLWWEX
iHM9grz79uB5fhEeM2avkDmXFyZBmZ78B9NFfIkS/TizpclJROjziDBdDhJfN1BU
fppss7hWqnTjXD1lH9K+FGc2NAv5QiuYdrRvPxvJA7CShrX71+HFNOnJTtwF1ZOn
6Rj9yXLBPvelTHileuXyX0lShHcSgUHljR2956Ug3S7Ifspx/HEa4k09zqFdf7ez
LcRymjsRTLhE4garMCA8UWShstsE2D6W8/LH/61IlQ7wmKRcEeKotnp5XIU+n5Gd
Zy2iO+jt5jfsLZcxau6DY6lRNA2+oY3IT533SYgk0HXWRpWHg0Em9e5lSXM4rjS3
IPhNOyGjhef0qE/cUYvnjkKr2x/nXCjnBzIfW5+dBCvMdfRQf2TDYoyJ8BHWipSx
3DbnIR9IVh9LPeImvcTF0SDVjvmuzrlTomHneTyqDZ+kMW/XyBEtTsH0/WlVu6eS
zu4VQUHHZUnT0bYt30uhkSuoCKY+yXrtUVDz/txCDI4Q+QbM/9pA/fbEjRKixXp2
6GyVvucFE9ax9lWiiGeQ1jSHOFVEirtR9IpIkc9V7wRogVnzu+twbZzKWLFtfHsn
KL1QlbxJfxxopnvZMb0aNvhvDFrBUTGAyFmUufHQuK66JAXrupdJrw8HpC6+VM7r
Dnh4W68FrdVwsQURTTO6fqkz8qNZNPl3PQQTOW5f7yF27I+3xxR1ZO452Ydo/Z1m
b9GB/77VlygrX+fEz21Cmqpuf5KQxFpTKcZAS5yNkN+NwKlYw3IrJVylDidx0Hng
6AUrmX7rR62/9ekGcH2nYB8YzJQNIMjkOAN4W7NOqzq6LXtEJsp4PnwkciPpxMyr
I9Wwkta/Q1BuEVVKyBB5G+2pWSbNj/zKi1pwTvHDhIqS5TFjZAlLi8KndqBy0zcA
wIxrYJ/gTdVDfFfblp9W3s1PjP2aCnbBtuE1icQ+mLL+76xuBDDgwne+779HQL0X
fGTIYwLNrihznwtzeHnpL4hvXjgeHW/o+DpXPm80H6px/xgcFgGWudZmxfjuCCFv
XdpXLdvd/u6Tz48Rf2/7sEeX6g0vxSmVw7TL35zOy8lWMZojC8POkSrna6gBhiFg
07zJ1FgIEoo6fYWEYfggZansYx1NHQZmEZ12ekb/0WoZA3sr6WLikN5HWrA6XSVF
1wyc+bidJ22r0T9qfV3k3gY8zViVfjFyPHMpEgGTDRtIGdyGV0uBDK8Ch1sj3AV6
+4yDoUHZq/lfk8udREj6z0nyRhPzqI47tvi2ilpfT2IgC98xj4Z9xhMsjm1lvWRT
1NoT2XoXuPKavXGSsD1UEHem4GZ897Z7AfvVCTCew+zJIppOgSOsG0FLxfVIlj6I
wcud3Mz9b2Q9ipvsyua68+zPlEbR2+5HXxT/AOd6OKUBtBX8bBMxArzsj48PNysx
sPIyIcrta1c5WnVUD6IWUQJFPsMzSMZGGRBLSN5D2eZAIf6iOyvsazlX/V5D+8gk
87vQhIhz04t8svo2MQ4Vnk7F5pOzG6FVdUT84ClY7y3/UJnptRVjgJR118OOOzg1
lrmhmDBK9I9WrZPHC84VqabwXS+JdPpWguBNacATbwXjkiERsAf/DV1xJ3cqWef3
20E9b4hgkY4XVRvk57QQsCtlszRLK3jAervIQ5LWq265IGlw2rCoSVBM4ZjmgZcD
JOGkZFdiujnzGvM912AsG4kdyiw2Dpa++2oW2p8PSGu3crBt5CLG/iDyKl+I6AG/
rscCUysR7jHBTUCqoMnXEVWTiKa2efrF1T88VQAqifdVIEGMRd0bKK2FcuzgA3oU
0tnw1rBBu4cgGFjJFqWsjxkK3d8Y4R0E/svsdI2PquX5dp1afFYkedTepRr4X4tm
7wx/FtxNcGH43p7pueLdDSxB6MNmOcE23x4hwEWb8T20+irNpcnzAIigYcCzcqJN
T9Z2jWNbNLHIuesKhao92Lf9ANqB6rWVVZR1GEMKKLiCscxwn192QQPz8LXm/eOO
eaUti/o1Hg0mlfI2Jx6vu1W0vXzzYhG584ayihalzQOM7Q35sHxGxDMnBBBccSG0
aTs3MAnFJeXHFRCIzA8QXSQTkKVMRzGQcpCKMjx+FUO28pleHzjKC4whvC6QIG4f
kBWSfbYlTtGYinHm/NamvY5dWZXU2B6ER7f7ldRspYLz30t0XGHxcRqEeIWVYBS0
LtE79oEB2BOXCQWqZhXr9XKzuD1LRlu8hzEvM59U2UL+Ku8xM4A7GW/tFhfuaLKH
rPm4DheY9YMYgCkLpsV3LBDRQXdzzTj0UvoTOqKA63GlYZaiTzMkItG9cqtmZXog
of4Z4KkJxY4mWfLliLMPas4VXj4pfIAJoEtH+XBreM+k303MvzE04kEzXM1+jtzX
323FoPYgr1hL6D5+gKnzYRReqHKUqjw/8TUrIRA3DfwJH/cA2WLPi3UGo9YZAfSc
W128MY2sROCKpbV0pIhoRekaGSr+vPIhYsZ0OufRpdmXoyZcgnIMZFkra+vZZfnH
KqljoZqCnZlgn5jTTTFP/vvPUq6RhxZR+JpVfZMMXUbPuVOViOzt4KATzPrpgUjb
hBIvTN7VS0c4ycr7kszoqO7QuT/IoGMXa0Y/nKpx8CC1kOVEqD4Sd5ZNpSQ+zWIX
i6wtA6xTI48WAyLCnemQ3glyavoVmIp8CEQqOSpkGxyvJCdNRkiNd2EbAVH78c1R
4cHAh3wsgVDS/E7ynsvf1AEvTjYTvnnwKlc4rMFQq330oet4GIS/3eK7lDtS2D0n
tlJvauY1JMwo58axZZpYCxxnkbiToDbrQiFYAeIVAam9jHtXg80bwOvhITfWI9Cm
TYu0y+ksGpe/pl9ZzdkVnMycrPgZimdzwKD7fJ3WVg9Q55Gcv4fGdXGgdb+XgvXv
rzLv2rOUxeDAf8qy63rZponh7YoiG+Pnv8dzGIJaaeFlc6Th1tG85we9dkYSVlaI
KagZ3oBUQ5ZgwX1bTcX8mgnp2ra7Xi1Py0WWEzviou3oe1jXB8hzVjUr9HTrNc/0
RE+HwPVACVDeQ1Xr9qyPKlRaoBhl6GwZDqY4pUhp5CcftfTjCZ383xkHk0ezgt7l
mn47q97MIl2Mmei+ZHBFm7x1ZPihQb1QGeELiu/WXe3hyEuWgLZUqmHzlAFaj7ty
dop1QR/jo0DuZPzcNuviOkiocQyI3JRnQTZLgV2jkaH83H0GLhqbVPL5gDwILFXr
kgpMVJuczuTT9eUDHEpS1SQRSFSZeQtywCwJjV61i0kfaRky5NWLVtpiIk/zROpT
n8gp1qIxN0vtTZfrGfAdaEaRVSbHWx8u9wMGjG4hGHra88P5Lk4mxXZMo2rfV5y8
5iXAI0KCVN+qskGHlnE5r0JUkNJJENyH1r8dcM2hnfhRWdjKfJYR1eW4FzuhuTER
SvruZf5WbS8Y+eOV83eopNVGjAVz4h8xdi5ZUWb00zsFhPR4Cg95CQGDOr20Oy0i
BtxiGx4581eM/xdb0NZ3KpoPhiU77Yc0mBvWPmak6aZquK82nTgS/Q5vrbzBwJ4e
U2uXUajC6WUP9OxI2wUV+olp34ylr2evvMnWR038lTw49T9PsDKFrpbu1LJW9qEy
QDr6qiziHGV0+hDizkGqEe+zksLc0F/yKvGGKlCq/Ge4Sp4nsosbT5nLY4G9tboN
ZLo/4289TOCzyJHyWT0QltVWijfKKgQ7x+aOz2VdiPrnnWdX1/3ztGwMM9+HpcCK
yHz9Q4yfpJFmf/NRH6hTAMmRj1EpdsrjPjTOt5bAMNBAmZn18IDQaN44B90U8A1p
mJv+ivlVikG4y/uWYc0Swegde/mXNCjI39liqvKp9ClzxVy/ypgpZoSAkntdThii
AlPHLCkWv4GIToW8CvGOdMFQad3LVH1V/P9Bhp/UjR6vT4L6/Nv87/D47HREHeuh
S7hLwCrKzssH0SdoqR75FN9Dz7YAShBTkY4x+joBdjrUsEVghvDP6PHClouBKktx
OptUmLoWMDaUpu0H1yNXMBKnppfzmHB63J4GODl5D92NewFr+zdl6yC7XB8zjAhM
1vuNpA39VK71QFj/poN7EE1unQ6VnjVSEGrbZu38xBckFo92kZvKokyp+eCP5+t1
79EsR2GQEx/ViuYc5eNPSwTnl3ruHJbacQM45UWW61HgNOM3/wM7X51oFhu5SXDX
C/B9rEnCi94w+h+FiX/4UsHWcy/HD2n0iFtt6k2Hrm3i95uiZGYzJjrU4jS0Mf3P
VnGHuS83uMcu1bd+EA9sezscasggUDyVvsajXRPi4z1+AjEDrysuZOecd7Q+xEV9
IT5xUPqvgWoLuhEwec1ZlVqyhUc8hp/gPmjsR5CbQIOK5e9GHAO5ksHbPq7YktjT
c4FZ5FQBsZ3r4wDdVLtOIB/uZsKYEu9/VT3EziqJLNjINd3vz2RknB2IzoTmitRl
ENZnfTHsyHBwAkuBD+qeleV6Si+XkbEY0uPbIt6gVnpuAWG21558Wqa420TzELa/
pOpTSKqD0GavGLjTQKI4TYu2O+5qsl2mG3JeI8ICYnkjVAHSUu0uVU/X1pC95gTz
adpVuCLWNHUFIXzvTuNv7w3phjIPfX+XPkmS+bQhXLE30WpxVtTQhw7cPNLznbuO
ODBj6cndnfEOCQPdsFHxVURA3JLQnombAJMxLFDxfenhiTopz/dIgrP1/iDg+u92
jJz92XXXec5NE3SqaoYip21q+H5Wy1x3MH1BYpgXU2YLOuEeOusVdSSA+0Hpq3dI
JcM+Avdiq71ESu98KNBAOLiTlAyVAmklf8yvIeHQWFeN8sPar3P9ssK/AWMRYxFr
MLfYcHG1SzdBizZfJQgpokJ/f3ou4ADScFIzTDI6+IQZnQnjOjM/bGBMIgSV47DH
pG2emquP8b3lVwFeU5veRNtc8xDoa70GXyhepuxbXQ/RY1bgVw8b8/3UZEkFigrU
kuFiV/M9MnRfLQ38oHVMx/8amyM+fxUe/Y7is/KhX8ynJ9ptYQyRTIWA/I0Bmm0f
kl7hLbQFfVit3qQOrdJ+qR5WiaXW16V65qDZjYS364EOlZnHaL0uJOxcE+3ofiqT
ygb23lebFbJDs9UYnAkBaRyo5QA7ju9fWDzEtSWZA4hhboux+r8Q68k9BXA91lvy
L0/fayTynVDD7+Cke5PGZSO9QB+73TjgO27us6t7db3Ru/lN3J+8uRPyChk3deCp
NjmpwPJwplAsbHJuQZLEHFzo8+enzZGVScL6hvmyTzGGYJLF4T49PsupS/uBFPxF
Av8LLXvYaRb1rImZkxAEFDL3qs+zuMZVTFcqTDfZunAofAluHtlKg3KlvqDRco9A
2Tu4Q7at/ITdmhe+nWKQ3wFc+GAsXS3DolahaTsw08XaXiL06I34NQH4Bca2TDKV
+1RSMEEjuOaoH6dyl+CCsSwpBJszlrNZwo1NjmuPtfFEwYgib253Ylh3RwBbkyZE
IB9YCN0aDn64OqqW4lQkHe4w2uuLW21IzpYDE6bip33J0zxab6xYd4eOtUMcc8F6
y9ndly2ZrrhQv6GnJgdY7odlFCrQ5AXUs/GabTB5l6XfrlyHPfBCTBoxT7JBdfY1
eGlIqU3YVybi1WnpiPFYKGwbePJKJxIuJcNnL6jyJJjOEMZOIQJsB9aiUTBpf26y
CQe0iRPiWJl5LnsapRsjdUBYMYkvvL4+lcCOLV5R9zHpBVyI/+So1+kFN610phJl
Sx2I2UqXYNTGXMoCqrqkgvxKKvmuZEkTXqzk7+uxQIn5HVLSJ6QTV80kRX5+Xyjc
PQCP7rbom5eHzCeqcMIruab5/w4G+tU7kSbceFCRx6aqcCWwRUtZE2aMBetl9asO
1+2TLiEmQU4d2I4ozy42EuUV2Y6jvegVw8uDcFoaNOb1zYPsn6c2qwGo2mim+rJs
r5qcH0RLzxAlqjvJPErcp9ePMCrrkHlPtLkfXovZUTkRn36t7NFzAGuT/1TYNyOV
EYwFRcmMQ9i4ArNr0RH79W62G+UrIY/ATHFKAI7YrBzQ4/m3MIs7B/QlOVS3IihF
kR4fDyr19pwUtVyjjWe0xzu5RaXjfG1QCNdLkxNMEUDwJTvmrbSJbCS3Gr6MwD7G
tGS0/SydSIy0FBVQW3U5jGB/hiUb/gNPVaZ0z+cOaivM0kkT/qPLbgG3rj5g6voo
xc2ZKK8zqx17PtMw0WH09eCY0k49TFHWJZeKZodV62NgV8KoKwkAWABizUHVzVGT
mzHcIs5/WiS9+F+YYR6bjmnXIzQz9eIksKEFCBNNHkXE5vWAzLCWEEP8NnjF+c/U
zI55Ocl9NI7MZ964VhAoKuQz87T5nZfLjoZDKm9EozB6h44QQEmXhAbZriDyDwqC
mUgurO685ylearNPDizu/emG12drHt8xdPwPzYNx3HEyhl8sbASeKQ3dacNNYu+U
eBfY6F8qZvSbqSHoG325973jM91/AiT8KCLn1rZUfwf9vho9n9VvEyXtvZ/kcr5Y
H/C6MblItbUIKM4W90f96we1LaWgri59cN8h0j7QpfmVwfdXPmzuJwOIRbbbcsp1
CLm4tBUCpYPg9UDQNRnbfXzOR5DGXMGIBxQvP4dTGM/lQQAYZVdAFWz8J6EJKj+W
N5r/tHo4v9g1JZQI+tomzOIaMQn/QTyFP1nuKqjAPJLPdV+d30RAbV7xrDxqXLPB
81LCaQHggjASf0fyUDuhbJP3EKKET/Uqz0SKkjRt8FzWwnfp4EQhSFUAtXiEjFxD
JrAYp3ZSl8q329LrRjgN2PUhYw3OfwudfwsLmM3kzJ9XHEk23+JD2D+iE06VWKSA
7fKOsgW1gk60z3xk+C5V/Kos6is9qXgvFDt5Coq4U+ovBtSwzYMsOI4v5aQxko4v
zFPxc1o6R6U08RuXDUKOD6Y5E9hyCg0Hvij8/IsRdgH8K1Ro05on4T3jzIbrepEv
tAxL4mzb6HtJVfr0dtwvRDGPmz70SE0f3R0pkP4jiuYe6c1s8XsIHLQkGKtKBFEE
mJ633cADFda96mNVBE0Qt56C2DCPQnU+YcAH7a2ssqpjnWX57kLf3iAv917TuULw
PIF5hByg1SCgflpr4yFVLuU0DBLfbO9Yc24xTsPOZKHFalSYsNtazFNLq3VIV9QB
2Y/sbyBfjRhWzBprSpMBRDXJgoxjBiVa6QyaCGDmiNFFW1LvF6Pv+P/onjaEllbh
CQBvFkCOCrBVoRhsHax5Bg/F4wV4iXpJq9mXWSlzguMsT5GDd/IgrBjrsZ4swGvm
KoDOq2pcfZ7Klvh9Boc0bmAxpcbyGAHhczMz5QXPXAHLCHmIj885h0z+AmZXxWVI
vHcQEaRywOf+0cFY+FL8wbPs91OGhS2P7xLE0Nhm9DvTr9B5AZqQ4xPR3ssaw9YI
8LpV+17L9B09Z2J6Hr+rBVp2EgUa6PEvG10nrf2uGyEDuGbZHatOD9G4NZCWH7XE
sjA3RFT5s0yIc0ZN0Hd3pJrXa9PlS3770EdqH0Cbco6uWuWgM2c22sjzPJVYzg9K
CugQhANp9motpQiX+mGA9T6BqB9vriFh2BGa/oowsDx74knuEWalRLHrFhRMJLzp
0RbDTKkXYSD2A+OQAStaRT7c2bZdK4Z83HQPQks7zNYZ52W92x+fbMAyIEJIw03s
F3dkGLLHkiqJRupOc+uFhwB7rBbOjFnt+AaET+TTUAjS5QlpxSorl0Ton8zSp5Hw
eEl8iFqcVYIMxunszF5PCdKEtOrweiM1HyIqLfTIu5J9MX7csZ5Dcyo3lE/s2sE7
siVcQNFbrCUBBc6PyfoO5Zuh4qIFZX+zScBqyqMGzpBYw4y+Ewf/NBgDeihymQJz
khsz0Ot5iiRg45SncsiYP7ni1HilLKMNPjFayhpg3e/FBsNJSYyEoN6tvt1Yr7HG
ufatV3/8RBliRq8UQ8Qgf5IOazhZZIABgDLGIIZwFeSgPXrXpfM9aSbRfhLBDJLv
aWoFTo8cuG07iG+UPTTr8d/FjZwi1yLOyIShwzC7UVLFjz5BKTFpLFCUVRbGDcql
5Pq6Xl24TJeKPjl+QD1Gj0B0aC1kBjSZEQASdwbgdlLzpn6RVYZyrllsio29tcYE
SY2LXBGbunvniQe0zM8IQP4+NJbdKyOhL3e9R+l0pC75uT0rBE2k6KoWOMP3Zj9+
gx5xWCYZ64edeZYJO8GYLnNsdf+2bEp99rn+Yh3OXQxejGjjje4p873lnZppHbX6
gWrrm47WhdYEz0TPnjCqw91/dRb5BLy9XFYJ5qG0r+JuKfUFAnlfXsf2duDvuieo
LWBGcVGLbLrK6D1bYkJoAH0o+wJ3vldaKpadoxz3w/OK3Vnf3ZHHAY5bKlV+8o4x
AtdRESVdSD8pCJZP1pND/iMR9OtmM11mdr/JxolqzOpaBQMknEwNa1gp3ep5kbSt
ClprWDUChr7Zhny6UbJeFxIKWhZPH7IIKWavr7bj1Lj70VpYd/uZX/W0e+1zuxj0
Zc5TdSNLbq+TH4/p26HpjFaTQhlZY0xf5z0/H/YtfQtc+hVT4Usz4dijLs9zYJD7
IDA1ENCybOmD/68KTYCuiKnCaoRbSA3F6nMMVT0aWV3+JqgujRfiAVO60OPYyh30
LWompUXjh6vkLr2ZP4emmS2ooKSmyoVHS5+Xgu5f+BRlweWl23BA4DIJpQVDyUAT
UNPpn268cRt5Inj+1n++cOZomy2VSo1SF6Ly5dRTWV7JTfJFdevkM2kRrHw7faY6
`protect END_PROTECTED
