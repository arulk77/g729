`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveE1JUmSwpndgqCwKRw4tlvogGyUgfMn/z/TbRsaqQTmE
C8ihLsDvNnTYMAnU78Lti7sMIitC6wyvYtejjOUBU7VmJar4Bx8QHnrvzdjS2qXb
E09Qqa863PzDksl67M2rqclOVv6uBPeb1zfiaiYPe+UeWsQVdTQVnDUP+441eBwp
fX1htUdE5i+zm9+g6wvpumfEP+Ok/2epnfLiXR4fZ+m5vEja5K29ZPuwfJ815GZC
MuR9TAKlgbBnuDXOO0KU/Y/HgR0wm2GWC8Xhi4hEIDeu26odvnZwTQ4P/sP5cUPI
kQbVHi3+Rjgdwt6+mfc47Q+oy+Ii7P2GSPZQCVDQ49rDnLNHY+CXy6sLHK4G3Y9T
t/3nQYCxKBXhu+gKwsZz5HsYjabpGOXLDXJCnD+4aWm0DT4KVgOSJelkrIfP1a8u
xOA6d/evcTLWxXeHIA3xNUJW35JG9UxBCMCMTChvbjPBBR9uwcWJK0wR0XleNR56
3hdajYgQ5xdOK+R/xtML6Em5TSzmpbT6RyxoO2VibSM=
`protect END_PROTECTED
