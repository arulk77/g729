`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
66OCmbiD1wo7n8KRAOex/zhLTfTL/gGhKmHoFoBDe1pjSfJdQ3BXzuDVpZYP8KPw
e734WmKTwfGuLLJTaD8ph2hLexsskC34l4QmMFQ4Loy2zKo4Nh3PLjcNHgEGIxij
Uo1IFXBIpxrc1MDFgXk+7FCR9SWHTPAm5nohDaRhrjKpXvjSRgT60w02KXZcULUU
`protect END_PROTECTED
