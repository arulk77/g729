`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFll4fBTw4sUqmkvXf/R3m5TKp6tfW9t5Tuo2B0scJFI
sYMCDc4Z2QoZwTegH9b3RxZFDk6RvGUq2mpFpzDUVrSVnMkiPjl8X4e8/Xm99TmH
2YMWsPWSp7LHxMWo7jtNlXUoFkyIWh6PKv0J26wRswtoer+JtlVuD3wzc/p3En+z
n/rzzyA23Hotmo5GuqIuKdOpXMRPROew83Wvocu/g9ItiqayDLAF/aEQxEf5f6JC
pi9vu/2xBYXM8E5emxe6T/Kc3dOodHTfkYG1UYCUSkqxeql8Iv2KWz77X0/azMbY
GI4kTqRXIyGUv45x3qn942zMI7IdXoHoibZAFkxpMBJmP+LMXTG47QjfDjYhrkoa
YXFcBzEgQXQPbAWRJiGqWHXw+TYvEdP8WgvC2/Pu/0fpKeDuwuYmktlYXGi8YsrU
Q/R5rkKLgyNcUXrBNYXtzR+sjJcP/d3RcfSPRTgPFS79cjqfI3rlkSusu8PQq6wA
wc3qlmayzs+zgFXdKD9pMtRP8nINTpMZpiFmuAtzy6QgRZynVYnNVSfOoHRwMhW8
`protect END_PROTECTED
