`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN0wOpOYG4AskTcvdtAgw9ScqOhIVTMr4J7kI7YwneWMj
cvE+8rD8elignup+rtRnAsgzCrV7w9coLcKrLuj7GXo5ARbjEb42k17Ta9n+Jutw
aWcRtRlYyVyH4xnIH/dG9GJXSEnA2wnj+ZU7U9skyqQ6jVF9s0UbKEoHSqRFciQ5
SNz5+AtDEuM5iSDENz997tWBueugOXd8iulGrDw5gbnmZ9yeCE927f4vO7xI61ks
B00Ct/CgBmEg6YNn+4wFydWutGHk4J7ll1siane568AU6A67G01gvlX55CO+a+3f
3odcJq1y9MOUslxqa9x+iHkbnKS82hSSP28YjbmivcRawl/KxA2OA7F0EM7Ukg8p
35UdkhKwWvxjETBU/xA9RjRsWx7bVdH0UamYO9/GkRwzN0xw3hegDMgOTsFp9Mnh
neVKohY8sTs/RbfmUYXIETMviOB0niA28vRHyZMKfxqV4Dt63+zJjr3MQERJvM3T
9YOkqRbiu62Wr6RYXxaGOhs+MkmHk/bOPXSp4ydVN3E+jl5bOglDhW9o05IMOyp9
vonlXrLmNB8ldTkrr+hWsy7JuZj6EWnFGY/eyG16itFn9WCL0qtY8gb2WAd4mEnE
mOGgk09aNkcZGKy9hRCUyR9IxsKy6wnXCDBHURjP3zV87GecYcnF5dWNDyGN0xz5
CtfiokvN7tOUmTMCRYpdVuR+2mFibPG4obq6qj8GB6ysNAepJWW52uoWRscR5D65
/nCLrzjEkVYUNEK/G6+6DuhTbVoNczQRlk2gV/Ma1VUCOKcOG5NsLIjAjU8kyLSJ
unkWslIvfgtb+CSgy8xsi8hCqw9FdJExrqKZt8YSLvxiFrGnveq7N82TXr6PFpfi
jWDZoCgxvodE0BR4LhMSS2qhK/2wyVN3RoyMtv7/CLqjTU7VL9ZRGIwvrefFtxDo
Qi4XhaD39EB0n33H/um6Du1MatpFvx1W0M50Tf2cMPpkgHWN4m5qbPbZKQkH1tTK
jdSHPh65LSf3RZUr4hLcZNUsp8kC/sbh9uRhyO8RXgxfzvcvWK/MEsQq/ommFsMR
kmw9UeSdvxGnmLCQcpSG3L5raWsO2WV2mBLQ/GCBjtY3ZLwnB16Ff7gTmPScQOS7
np8nXMIsy2IwMW22WuIlIn/6m+JMvsmluEDE/bLibwyBfd0Ka7WKSMCCZki0Fc6S
Q1wK+yJhkOfwN3/eAGyJAwd9tg7LLlOxWr4HQzHFfHI=
`protect END_PROTECTED
