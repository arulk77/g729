`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAiFtCnBa6IVLcxavPhJUu+yNFive1Qf2ZbHqeYuxfMp
IuqQopwOgk+990E9Y5xP9te6ezDZHkXXtDn0KwUyGNHaFVnsde4PbLlxQGiOYTLq
kEtQBOU1/fd4+0TqUYSibG6kYOo4D4C5vXb4ZXuNs0aBMKVQWvExrf6LyIIzNyZ4
+mvWxL0FVIr17mcgsHVz5KRH6cMdDmmaqZ0n+XW0IyTScguQMAEmzmD9/2S5+iFD
dKrazw6owzTiIdL/ZBD4sQ==
`protect END_PROTECTED
