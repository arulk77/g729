`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCY95y11b17403ypLrgr7arOg0kuK4jK1nP6seuu9Thf
6eKaFlZkT6ukTOgGTVNerQPRU0emgK6g4UsUb4TND5Qu1NH2sNptFiuiA9IdJi5c
Zs/+eBARU3u9Ra28OQfi+B36a0LQ8Ur0MVauDASqmriHLthmHpDNCa607Lejqh8b
c5+rbX0/hb0tSlYNlm6pdB35QbLjsepNeSCJgY01zWgwP95BslIbyoC7r5RKif+P
rVEq3EpVLt/WPrtJ6EvW8cqC7/udUYkDhbrZgIV0IrAazULH4g0aMLvczoZusbVt
F3L+ImhsJYvyuGylvE+qNZem6X4Ixmouz28SHbRFrCsglyqWR49EnQJerEITOCZb
pethi6//dWX6iugfZdrFrPKTvO2JkXv3oxUDjqoKVTAD0ka7GkaA7F2L7qJDfvzJ
UgtUhuxziFQ77Ai64u9EqlYIQgMJMJtLkSgmYW4ps8avfmyvs16yXlGGNKUBaBP/
0ZsXwy30eAsgbs5rBqMbnQE/3fe6zcNsdmtXQrHzZdlUur9fy2dpBnA8K5jOM3v7
rfj/3t49w9NidiYOCEWnLN60CdGJty0MHI9CfekwHxaPdBhHvuvH4IdndBMKjeDj
4JB3cU9ka8zDOyJt689L/4jKCO4eTzUOPp5FYtWlrvEVeDOsGRapWiLomyXW07Gw
`protect END_PROTECTED
