`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
tIhGgwIHiaJ20/hYB1Z+kTTW7pWCIC6b/U7FRZKLgJwpysmdbpOwplqb/fb+AnRf
F4chlptqaYQ2PmODi8q68TzdqTlHxB8uJrRa6n1D//lzdN1hg1pgudEuoDadjscY
hyOn9P6OtzxU6NVwZegNnVNp5UgIWZKtL+sea482jIbtX3gTxTzlK4QVcdQwBLtl
39RPvIr/RlwoSGxWBSSfAuLQ3Us1j5ucaDfJqxIZZFyrRzI06abyAOzepxh+30bO
+w+fRqj9iHnFsIT7ikrd5U3XmHKGenS7rin1STVPBbMwUpXbugQw5SnQpPjlb7l2
NgvkHKbnRm6O7iT/C+kCgMoCbYPyOKh8si9xVOBPOEBDY1vbszj6EpmWIuUPwULu
PxkiEj9W3KdS39GeuihUpemojmFjRMZRkRWUN2L+83btlbszHRfYTb0rJHbBleXO
I9xfU9i+2fTVQqxO8UXd8NiRQXy8j/L8Zy138ZnAGCXAg+Y7rnINq84bCZKyFdXc
BoxuU3nE+E9aUE41sMQSlplMO2WKVtvPCUdROziOAyMUsKFZz7tJKDUMvtnbqpk/
dZDl0wJQBaTiOW15k0r688L2CtCUR4U70moQ1J9Xy8tbDSkgyAb4khSM//iWYE5n
agunE6v/d6YB/3EsyenCHet2xmf+XQOmwA7Z7sya6cb/H3J1V+piwishqPsZ9wZw
/KXzerI1jCUU1b4hUDF8yMf6iXGIeFfUfsARvl4UZDk=
`protect END_PROTECTED
