`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDouqO1dvtJTo4YvXh34UR05gu2NBvxjxQGzFkwqhIU2
6nPHZF+MPnM/cJEFyB6XqHsc+hacBk/EqtuSh8IUwsTA1nCPALiNh0RxAbGLuKxN
V1dpbOWXXup3HLeNaKeu4rTZMl28Rng/H9uo1ZmP3u/hLKEiU04kAaFHC+sVZPB3
iL9sVSS1XI+i4eWDqwa02YdXhuCPjwNXLW5T6lAo54/WnTbfqkgi1Q4kjkW6Jxd0
`protect END_PROTECTED
