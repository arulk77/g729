`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNyizsxM1nTfVVaALctQbEkyscoqzU6FlEa7V3XHj6UVC
fAtM5cHE+mKGVQih9YFJPQemloFQ5zRlkWAdfeoX4NdU6pIRslknEXc1v3c4uxhi
IH0O/mgyLQpBcT+1xyzDq0QCMXZUaP94p8kjelZmfp1jnUri+GdOn9E+2v8+5US2
7dXayxii0MEc6JotwXWMVMazm+4DT83tSMmXNzhbz43FHgQE6LAv9awVRFx5G/ZB
oMWZKWB31m6v1NvFyMaTpJ2xRjU/B0hJ35eo+lQ93DZF/dWxl5bFFfljd7nV50Eu
P32kKC7rggbE2jgVSM7s46yMeqLHRBLZn2kp3m2PTCRug7/lE5633/P00U5I96au
gyutN0OYyXKgZ1RjLr113BFelglqYuHAZX8x57xOFBzI5LL4xjCYMCiN6xzfN9i8
/jNF/zuiTCpJs8J3KmP5IAGWUZFrMU7idmbVEz5SGSs+kMTVWYsLwQ1SqzS4EjAy
UMMUxGxW+PZ0Wm7Y3RQWs5UwGV6271AelmzuynK2noUVOlERl/58Ju8Gz2c4ZPHF
LHHH8RwKZPYwFECbPCOqP8zKcaGFTy9nf895rI814T7fgPc2tZ/ggXwM1bvXjWDY
C1FUd7CZyjwEEo/DJiNoDbWjDHW02jeljtWfCwKDqMybCwt/sBcmTn7H0KvCShEl
gY68GN0tBB2aPnCQL7M4AGL3GCWN+jqjhw93oGimYa9rcI/RMLyAp7lkIwlHlyPc
vLsztyGzv+VV7CQRNoM66zx+lPCiBg8s+iXLuS49fpaksx6A1QFNnZzb5KbMBkdD
0jWy0LiPRuqSQMF0B8Xb6k9WT/kwTxRI2MbSf3OfNhRiT5Ww8cr4ed0LzIxd70fE
iAMlTJNmVC753zSwJeZhDwQqLWWEorGa1Z6VJNjldrQLR87stc4sXmr3n3m7NjE6
bpiK8BEhhCck2TQ566TkUydeG0HzSTEzQ6ZA1B3OjDCK8HILxGuDiNdFLzvGKG2p
PQo+e9EeDnE6PnE2O22wuSZCUNbSPE49nhGChU0mYvpo1I1J63tQAtIYrlm0kpJs
KpTd0eOF85h/RYIMX0BmYTvRblzp2yHGeWU0NklBB6jSxndxz77PFHj0GRKAAY3z
/xLlh+O/n1KwTM9B645dipMaAZUreW0mgwBMDOygoJwGodcWyWhGZVlzeo4Z42iT
isQN7qk3ls3eHRuHkua9Zo/dL0uQ/duPqdZOtAI7WNk=
`protect END_PROTECTED
