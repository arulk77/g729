`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNXLt3tRQ+AUKo6cxh6xYSJKCChKRgNLdUjlRrQrCIVI
4X1HuyeO1A6rVTUd0teFA+TTxnTXAG+/pTQNjPPEr2zPf4eJLnm8dyTT2CpzO2Qh
GX/dD5xfp7fTl028LiTvFLHtj5a56lbnwMGUAwAZe2Ja6kYGuYZQx/yjwl/qxvH1
VYNPLQRteA4tTmuqKVfvf5zYVCYdig3nWM2UzehKr7v3LAyDuQsDE3CL5BdqI773
`protect END_PROTECTED
