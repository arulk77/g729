`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveE5ecnEXROhpXYiFRa+ku00ikErQcBfTFHhIgz5KJF7T
TiNnGWrqfv2+XaCIy7vjfwx4b4GO/bxxMKYLWIZUOeeMETelXE7s15bExs5taXXj
UK0FXlu15fonk/ugvnie5MhHliksJTyON4IWdia0QgkZj/pqCCsAdEptRvGKAD6b
xZg0uTXTcIdJe07P1FfjLoaPNxvO5PbdzTJbx9CZ91vPY+7+IE4OLtYlIICfpAv/
slqQdS61KYBsnEwdUnNArQ==
`protect END_PROTECTED
