`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBzoUTJYJRZU5lU7r2Pe8Tz0TOSHz1FysPJEO/Glv4v0
sq526iwBb//Ll43b4Z90j+75IWZ1Bv4KbRbEwEk5t8/Bvab6g1CHchMt9jOTrkVd
W0oy9lQNXACdILHCih0Y1h4eQzRcTYRC6puNgQX/QHSQiLfisHhpQqyIxd/m1euj
qEdt+ZdTItJvLxqYLeTlwBt8TnBogVyflZOH6LqOgE1prSqoWWeZVY31T7/AXsV4
gFo9yfKRY6TyISsStMJjO8GxLrk7er0o+79kxR3u3bMNeylCl5d2nP38vf29aqnY
ijLPkU7DydsQ5e0wmsHEaefuTpOkBNI+ONQ8DgCpWho3keJpQ1FoRAUNSyDwQB0E
`protect END_PROTECTED
