`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGcBhNxTRZrvJB5oxCVdlgBuFZTUfw/kx6jlGk9OT1rb
2C4dqsSEPvolPFEGx9IpCXjo5DtceICIxzT6y5teXqk7pMXH3NnSL38Bcjzop4kG
YjYm8vSS6D2+tj4M4pL/aNyx/D2IzS6zfT7ltrxEDNSzJpPGuAeTNC7PbbJ1c7SX
LU9ykZC4eYxbuNaCK8R0gw==
`protect END_PROTECTED
