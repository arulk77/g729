`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SULUMQRzCshCmIWNdKD36XQjCvKzJFjFJq7JgSJFNjAg
LTndQaCiyGthDfuFdZqOnYirnWdNMF3YsyPVz0JoBNHtT2eFPOyngwVfSgvCmOy8
LuH60ZndberCV9yeDCYelK8RKGlzVYrKmYvbKHFZq2HKWCC/p7EmFkn7zRLBLIXU
NUEkiZ3mJ9IRI8dfvvvuWDRsllyj57VIXinH/ZHrJOaJ/hnA5ss7seeYCh2rTz37
QUgoQbnxg6nCUvwUqiTU8LnIV+gpec6D+ne7nc2SV8spGXgWV0D5IZz9pdUZx3Ky
WeQUYgUvbwXNoiUhWpw4mnYAfuYg8/7V0c1a14TzfxD6TdV7iaBBXrP+p3DN3kCA
RtjS7WyUb38OUECrkgR7pt/luaDMRdcxyhn2JwyfNuKLEaqbeSe1TsEM6iaPV2GN
8sFUtXqxK3SCwUMkudMrYoLbeWWbBTUmHwBjprvMhOJ9bzDLOqbZkKBX2Wt4NpA3
qCcQmzWKhPyrlJFnKcp3N+EalQJ8/F1/1NfyuZCcz5xEaehGHHloNUI/hc03GwDk
p0n3uUVNWCyG/o7aXwwTljPRQg2DJ8IZfjqZYYEB9iuWBYi5FsQOVtgCJgfWQ0Rr
YBxJhIBBaTzWzegrz7owVy0r0hMEoJMso8safFJdkIkkme/aVV3Ce6W1X1HCR7B4
q46CEiVLh/IgZN8/V3Z1YzvxHo5++7GHJ0ohlU18/u7D/5AbFXq7JR5pi9B4RtSn
tM20eNJ4CV3fxCP86WMJ0Q==
`protect END_PROTECTED
