`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
p2KIp4ggWUXdQFKrbI1jfnE54IgtMA7zWJZ71VLKvuXXNiKnFUXQeEj5Pni7L64v
a2i/dj4eJJsTs0Z8BHhbm0eaG/P6dGvDbi5+GIhq1q9ceUWHDE18FERCrOOhdQb5
05fAF1r9OkVqCv8KuCuuQdUk3z3mIiQlFc5UaybRHRtKQO9CFI6fZZM6JRkOndcI
mL7s2Q4pMytwQ10EELUMbl99uiQjCyE5/PbpK5V3PHzGLbUjzbc9+U0Vc4ZA+pTs
dHO5tZ4/ehIogNWGCx1hnkuyEwREi9b7UD44hi+IleXIJTpUq5FVbggKhXBaPkbc
GBwsxj0iVb6gSl9HpytZR1mBahzwqjRVuC0Dluii2oI=
`protect END_PROTECTED
