`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
GzyfJiYe1IOwqJZzXOqptkWjVZ+U11F09c/yNerqb9NZgAgSRuSEzXuPDocPbu2+
+pgcGZtr+T/cFsR0PqChyDtIJzM3sfuCtquFlKK0eOUBvgZ9RlElyUstGZeasiuz
nMZVqf+B91F8LQZs5e4HpHN2EOzk+2woYZAWKGwo+sPuq+Njxdxt2Cikq7VVyoZ8
TEKCa2HP1an8Cp6S4GCB+ieqop1FMbMLwOgSYTZODgOX0l3zpYclefnthH9zhAtJ
SejvAMQqvMJ1wutYie99a40W+3RjGtNxPG94YIR+pY51WOCRj0UVnBsOVo1sr7qq
b7YZs72etvylAx/5JaBK+/9R46cNaszonXPQqsoc6I3vPK9RIVV0u6y86mbyGZyZ
93u72PBZJsEe3p4dhDeNhotsuc/i+a/gxweWCTIGUB6W11R11Nmtc9nfdnMzSZmT
xHWy9voqbik62cgp55BFrMw8jbrinWHioQaBppwXN5FXhMGe0SFhhQI3e0OBTNWU
I2Hkw33ZPEAhOfMXBHt0AViI8X+H3FaXLfpPPgT7Ut/qO0Hs84VD95w1yXtlvQlj
oa/jruyWAFFu+USy8MDPy7OqIehp6hx2rL73aKAEgsoiw3muv7vO30qbfjg7TAgF
MV0RDtCubRpxGHbnpEtxTVsOvELQaVh9hHbmNeQALUtIIjjGxlBEMk1gvLwFyjmr
HsRik8Um2MFjB2aKrkUVXCt+obCPPS51hU3LUvaIe2bK5j9zuFltGnbj9lZ+nrvf
QqW9GZlzpUqTw/Il3vq2R3Ak61NTfeM+2nCbTe3iGziItiAwQcLFTUbMKdsBRJxz
wSvzA31tOuMnsenBXWwtOAssD2/hUrNd4aTES/LvHaajDNbV87keLOW/1kh1OEl+
/r5wnwyuq2/Tm6hNuAXKmv2VfuuE/hgrYY2eGyKm2hXpnjx6Qo74gmZVJyNXJF5m
N8s+VUvRb5gMNWkfCRRvkUUzTVGxMq4ZehBy/tqXf6vvjZQ0AqsuLTMI5umUH6F9
OxCVMaCFt+Sqz7xT5JkA+9qPcBZ09F6Wv4mHMl6t6y+InvqOblCyhdiN+qK7Tje3
fm5FoDNCmsQG6MTjaNBDSZ3KjEnW5yER+jAMLbdI4v6hD63He2UsIuPenT1+FSkX
UQAxnBHbbGw3VXsh+q9jr78jlXw3cGT96cky0/TB77g=
`protect END_PROTECTED
