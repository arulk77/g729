`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
zUozn5XkqRgfLnaGYHgWfkuo5V51eFCaxFRFOrF3wiBO3Cok1x05fgXd7l2Rn4Ai
z0cV1TyiJy7prSjzvvyP8/6XjLaUsn4k4iJhNRNI+d9kswC5CzJktiQFLXO/mZ6k
oYcsOUyNqdio2TqRuOTThMlHLgSKMqANar7iwacD6PEty6n8EAZ2N64VRnamhT04
zbhrO+Uwyd6n2rw93I0shHiWUbt43BPdr+4DyOSMeW8=
`protect END_PROTECTED
