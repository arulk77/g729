`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM8xw2Hq+wMj0ytH58ZVpJXK6Ta/PdLJ7q8i/SLcKCXU
bto6rZYrlyVd8adn2Js7VZSUkxW4Zu1dzazSXftRnCmg16zt9131DLdbbPPR7NAU
VmT0CpDAxcKe6yxlVuv2ZhAhonXmsZSfvCguscJLqiHGXp/v8S2Lh7UXgnQltXuw
kq10Xxe2ltGyHnz8jAJofLFvMdZwdxNo1BAArTUfq9Q/3SViYCZSHsetbCxEK/Cy
DEKJTZD69IJOolGCkexVmBWYJsFHTXMOEN1Qe2DNLYD8NZf/lprmSINb+Gmjve3N
VMaxDvsciv3ZIQQ5kuUWEZBOz92yTjRhNMMwMbSBZwM+/aJA7ELG7lBvhgBR00r2
SHWkENdJN1+Qk35s4EqYdenIoYAQngiiDU6sQzRwq1+PcnAzjtLuYhlRG7xk/Eg8
Njbp/fT9an+OJDh2SQM2PCJebJjSF9iFOeG2/NZvMPVBXr/3ZOkJJTyL7to8kG7e
bOnEpzOuWkIJSj28VHwJDMKV5wGA4cKiBOBkZvBFmYA/64kCa1hE6c+VO+IabftZ
+rfmbmcRmVgnw4HvYUJmJts/jB44UN4UM810qCG/SNQ=
`protect END_PROTECTED
