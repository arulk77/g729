`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aek1BIxuG9q3Nccdbu/quNABxauNbNd3Jg4q0VbP5PuC
i1fgAVJiHKvSDG+NfTVL3cR3s2q2wsE3AzZxhzmkUBbG/velrVwNoWWYAqOr2Jza
e61kSTLmYHXKiXbiZdAAkfTBnE6NvA36S+BkYMKPKdogw/7loEHdPZkKmXoG2gFp
rbf+0xVv+Hw7BwnQJMDA3wL96A0mvkgtiYkYaptaU+ltABxdJWg5RCvIwyVgbcdS
TjTkOl6CrCsjM4VC6d14li2LMnuHPueN9ClkLU2NgfGGR8u9t2u6z6hKFvqmj+o5
7oGHYA8p7jfBV6iwCXoHhlQOGuvR0v6OKHNnFlbpNxWbNzWlIBveiz/SUDyG4fDX
NVVSylR4icAG/yUOQ4C7U7fqUiGu7Jyzt1hMuGrnOcz+HreAwlH+Lw03OZPLJ74o
LALm5sZXU1jrU5zJD2r66y/FrO+pD16cmPI+3MNRhXjAbeYwgxbx2fA+KDaqmaZ8
7ZVLWQwocgyWzoCzPnYRGJF6kFKnGO17sUeqp0JIohWYxUvvmQeslEJyuuIeggq/
0U1cOj+2ZVGrOAECUOq5ImUjo8Vj7ap614GVth3YWRo=
`protect END_PROTECTED
