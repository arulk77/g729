`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMWnW1IoTh5/8itB7hPVUyZwhkUtbnG5BNQlB+1B+pvG
bR9nv5T2e9mP6BiHdnT4UKEh4jmxoHNu9u8SlZV2HmjlLYs+mMvaRcVv8xZdXXze
f9M6lVltKEQX4rGWfP+Qui+PSSODRVK2jUvpW6Q2iE+yUUoURWfGaWr8tofTY/W5
aAfsHJ6K/JmMpegAf8J4iQVhXhjGo+IP9tOLWQQ7KgQPWI6vh8xJmamDKXM9x147
PYjrrMobkoo2CvuD85WvKd2iAdvyVbbqRdmPGE+oL3kCi5WneMfIwp+5uVUIjQSZ
i938DKv8iAIOK6a78q8RaG/ZhaBNfsTaSoZt0OeWOtI9tUfuN4bJEb5hZoU2njRm
ZsjysYXKZd4jV3VpJ9u7TG14H/H+2+y8dW90pVYR6jR20421443ri6QAr92iiUFI
Yy5P6Skb+tTM5OFwzIUXFLimDbuZKJBlpFVAGryRQoTYCrxBXTqEtMYsL5MQTylU
H8xhTGWFj9TMNq/3bfUq9JS1ehutA6WKgo/tyRuFcBMGldNJTPazq7XebeuhboYD
`protect END_PROTECTED
