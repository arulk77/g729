`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49Y5Im8vgPKl0553WGujTKJoNU+JKDrxoDrnExdCUXUg
WzGbz6q0MVuSMMe6fOL7AJvEk7SjRHxmOZbt4/FVac3hLjASRGsfbklB+mGYjXs3
qgX3Qrq4LYKQoDx4/Yy8pisJRzTLkhR9rnKXg0cFpjE=
`protect END_PROTECTED
