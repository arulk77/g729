`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIO9vEAsYYJw9t/FJB5tSz6bAHyNUbPVwqFVeNeyQNOy
JceOy6+zJwH7qElgiy1dw9WjZCeyBI8mtEmGzQl4Nagoj78VCmOe/0FhHNwk6SRD
+skTx+HMRa0BIkaspn8GhCVUdqCFOAbANf1c8sEFmFddbJfBlyuuEHP/JhT0BCSx
CxvBmZBA6aIpH+ljqxRJ+31RUiJXBVVp7VxhlfuzGLnHwsY/nyTlRV9p5fEApN4m
UF8qvudj91Cyx4ccjcOpBqa/NeKM3mBoEaIgGmGDT4kU7BgsDWYN2xeGFU0hAObG
A3ArA886VT64RitM4lqHWgwXDs9psexwe4YXxyf89hsQ+k/t/EaBQ6mYIftyM3XC
VTY0CNIHjQiJAM4KBaA0cGpH2KdJfHCscfnjl5eM9Xv1Plymkl/UN+2cYeNnaR2e
jEAB25qpxSqIzvnRy/pvgd/xSJoRWEnVLAFvXVF6GXOhFl2iI7yLgyMDWXvnlQW5
iluS0Hm7nHavg2YsVgO6nEHTVfCdrIbLkhVKOOiQxs/A/2Lk4ZVBlP+LHwGcGNzl
geBk/+HfinE9GW8DO6xeoN+XnVsT73CWYX7SxCc2BhZJsWmtE8Ey7cyGYtAztESE
audz/fky+GfuzBYuvvgtt9Sk0sgxeV36wgmVbUN078E9nB/3JqghSvY0MxvLQbK5
xVclFSGIuadET/+js+8G7kvYRIYi5PhH2Yh+FSlirIbon2P2irAn3Gg8p1WSZNEx
UwW7bJmSccTyA9RrzavrxtVG8fRToI5f+s4v+4K5prQVCRLleXoDlmaSWMyk12Jm
MLQNG5I2dQ/FyYswVUarw524czhCQLCCRbWtMm2TiA63YhNe+6M4XqGmpztYQ+pW
o9kPxvIlYSPrlZWIFfLmliJcCCkUNn4BoFU/AtuJMOpnQRiHJdDax7a/8ng7ZccI
wAZA3l81JYshczZyIRcomPTrVqfOLghEbCfjZeZ5f3FiunSczUsNvu9Kh5rD40TY
G9cEB1KWdc3FSuJV1iQdz4HN0yGGUCtskLeBIrdODqqPEgZzari4XYJHPrvCBZYE
dwkr7h4S9cGsCfwqvoVKWeneKu0jCYoJ8tnJvGKRNwx1W/5EclMfu2Giwnh/iycT
eepElIUdC/UsLCHVPyUfz6Witm6FuAsrEIDOLPExcJBwDN4vsTczRRZ1IvklQo8U
wYNrFTVWU7rCxSuUco6SO6EPgHgaLtg1U5ulMz6yTL/Rv9fHJTeXVKvlcSyi5ys8
`protect END_PROTECTED
