`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wJ1i2ElkWCeopk6nnlXL91scMmctLz8JfplEmj6th3z
vBKFiNSWH5oRglwqUN3j7YgBiCgA2zOgE0KGr2szgAlb6jbxAzrbsr63uSTVtobh
DjfU3i3lPE5sBCkpXXpTBOVkgdsaxgOwZfbJIfw56pvxytUZ4YB+F+fSOrg1bAQu
1RZ8lcoYj9kUaErutSY803ht8Dum+SFVfvnrpUJJyxe10WPY3FMVZJIcFACKbxPu
RH8Wrq43zkU77GOfmX0OVF+SwkcE8kgxIyYYPmunGW3CxwKAN4TgGcKmFzfpZzIY
cx9UhTmCICniRpOlE6tBlYlSWqUeC/5R3K6UKM6Ryng4H954hr8lvlpKgQPeA2sp
p1SXHaTcAkuDrds2PFGFNdg5hqOXrJMlN+hZyvukKr13FXCP6qMY16sZZNVsfSpl
b55D8QOHFbhBPRceAPo8UDa31WXJ3QWTlynIcKDVyKeDBt+y39ZB0+nRVozxkZYE
`protect END_PROTECTED
