`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yFETMOsnJrlgMpuGo/BarSkw3o+zGKGeGnGKz397P5a
fx+vTdmmCx/AhZnmh1btGuk+AajylwQLP2rOaXqd+Sh061LsFHz8SwJk9wAhM7dN
pUbw9WW0nOvs0Elsv6/jzGWNCbKAf5hH4T5bVzZ2RYAa/UwGRIvs9ZCu4ldDlAE2
sCR8A3futm0Ck7YAHCAnRijjOBxDmBq3J0Qq/iXFPikcqIjQVsGc0PSMMEparsV9
/Es8gGctEp3yUkPGSnLGE3ov86j5XHLDqEiwCWCgO+CyKYqLs4S1+8avnu6Cm7pu
FPo5yugGztUGz/q2Il1HVcKGAaKVIe9qKk8hugAZcvgaf91lmtoKCM9dgctUbvVf
Umkh8cX5SiL173AMpTXGOw==
`protect END_PROTECTED
