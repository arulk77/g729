`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKhqKdE8qNsQSw4XTRNCTxrIGpwVb13vV72KldQGuPgW
qGlMTFGVTB9MfOB4sFFwYgEYpJp+bwmM8eVO+GzUiH5uUfA7ZOh4cGiTZAdPgOzU
zU0DZXV5pEOoQ72/muof3NGyAc+H0ppY9/bXEPxv7pmqCHxQdgnvH1GowD8033r3
2yNptC1sz38OHtpX9UBGTwEJhqApOofTvIEuBe/sFN6ZFcK14x16faN2COiSa2Gj
6d3uHo1tUkJg3+/f8RLH9ZGVOwBNroqGC3HAOx7QjPGmQ9A8/MrtO9FgNmYB3/5k
AYS4jY9Ugr2Cevf8WmAKqcT9yrG+kGGIFVVj4iPOEZpKGCX17nlse1Q4uGLUQzu8
U8hbs/BnEiYRBa2Ybw4e7XthT4W5JMbeihM6ay96TFPuJWpayvLuLkg9eFoTkwuC
7PlFeb4Nmn0yUTyr5meZxDCU93bPG6jZD1EXVQsK+VAwTsOPIEumjvM7j60W1eJ+
h/npJVM5fH42JTNrqIr4TI8M5BHKnHpHLF/moFSYwq/5LxyL6HnfZPFfgVPLB2sb
eAJksnsZBdjNO9oGM8NdIg==
`protect END_PROTECTED
