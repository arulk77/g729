`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN1lcOEY/9VvdU7yiLT3Ez6fv7kRZAad4o37HbH59kKcf
kqt4mgsFDQcXRwTaSLjuY2x6BSuGZ7B0/jlmUvcXk4uGmKl4OsYmw9bsIgcnb8z8
X/s4aKDA66ldWSeefq4yulo3yt6C+I001Vi9irdQZ+ljHXpZm+gthevPViK3p7ZV
yFNAyF9rNsRAUSk9sZ+JuU26pBbixPNrb8upqlrdu/lbaNViSFYXUKm484Q372Ct
/Spqb8CeH6guWNxP34e64KPXuFzsXUjH9J1LkZ+Uu7Tbmwez8tlq+dxNODUEHGUc
YP4lvfXkhIYdhCqEknVBt5uVdOXcBT3UCrq5GzgbhdW18O18VNYuA60f31gG1eCg
LWhuXyy08/QTyItvWSP2LgR2f4JYZcgcyn0QQI8qr5/tvaYoGnv82W5+4ThwSlAz
OMWWeHjsRC1tK+nbIMmRin/W1tuPTPlltbkYgSNj4it9IL+CuMGi8i1c5uDXoc+X
uxPY4GhQalMJBSNe7raV8S+b9XB2KVw2mHRhIXMxOnrcvUiRYkF7ETmTOtBOVhOX
8AXhLZxJ2MSztmwiTvjIJ5nXVIvLYVMHP1Y4WastUwuQO8Ur/Q0xBvQANV+i2pH3
uN9kuWKK/e5k3Uj2wW/5cfIQfH0hraH5epMS9vtKrSfoB7dmS4kwQzRFzo5tQl+g
haJmeaqVgmsaNYchBsCcpRGCiPcv6/cn61hBeBawhvlWthWlsELE70sx25T9qciI
akVhx5p8IsCnaVypvGY7MXi+9CBcoRWKNLpVVjHCsuTjXlpIaCcSmVeBbEC+J+of
m140sE6jvzhZVILUAKLeuWWRbe7AFMV0g8tsTKdD/9X0BszeFw8ZqkETzujKIGmO
o+286wCZGpD09orYjJu9P61k3OLx6VhLY/DiVwEyodeoFoGQ9jr0xxHzZZFncrV/
KQ0dHWsER88cuEBrYr2RU15/6fi3XnQiuGprKp6UG+kIPifuQHl2rFy9ebeZlGmj
jSMGKh2mRYxhmG3g9gTJQO5hf07llDvfiPHLQVpJc449Aif2VZAcrDz4BdeCrq0O
9YUYe/iArpM+DzBnhy3BHSh1/Al7+l/8wmLbrmyScDXsHsxdQFRvGVY12zg8/nYZ
Pc9sIiLEKNZAYNWBJ99YxaiidoP0NLvwiX4m0BfCyNnieERjuo7W2B57YX3lzbar
EF8k752TFTTRCH5snB4RkeguS5kHBqF6P3z6ToS3sBubLgLa2tktvNl+SoDJfvYc
6Bzb4xzP9junuxy/KD16EFVUP2BLvySvMcCsky+hTGW6fXz4TnuJnb1IOieSS95o
1va1CSMbHpuG6k8Hc+dULsQfxm6KP6LONdI+TyU2RuWlzrK90qHqD47ic0WZMwUc
qkZdT1pzbPNoyds3B/sFNi1liECSs2UkuxJ0Pk1y0PcysBdBIKRpmORsy4rsGmo3
A6FtaWmJJFzOuRQhBZg9pIDHP7lY0619r7dM3cUe3Yu6B80V5eHEgwy3uCoiEZXd
pM6MMMUSlxufSuo3A6BRFSht1g5E6HPPdsbklc3wwso5nk43QBnRpXsLTa1Lp4xn
Ou6/qBu/0GDtjq9PEqU2gxQM8gHXovhh+27FJyU/weQQ1VduRSEAIN1umL+ytKd7
p1BHwDyCwTgZAXtRniu/RlXRTxL8/UbeVbGlS1aiOdb/+I1rNVJEj1aM0S3fFPuV
QLtKJ7EqikxgfXat41+PX80VETG8nVqK5JVCPldRqDzJ+qxdWFMmZrEflwcZcgCz
/JcGvFBZCZYOm7ZS8tKeVCFBnLPJF6/1IlZyZxSEKsaOs9Jz8yHjSxx7dWcaPgCz
QDZ+gDuRjL07VLnyltnwHx6qs0md5tAHnieFaycmUrHAK1g6ALRhgWV/xUMtrkxd
84nCJvdiZRxiQwRsfYqpuzAH5W9H3BFTZbVbX1UYkaQbwNlQE/MqhmbFY3m1UQVp
OtHd+oiWFNxzqwcx9TQeKWPiSAbkn4L8bYzgtXfxMW0i/jDHVlzv8N+ezCiv0apM
g8TArAPKxCfyVCjfdRcvl20XkGJMwl44ETjeM5wsmcEVRcqVk9Y+viQBupP5CXEy
+371pE5V1P46k/J5J+OwPxh1MCyM21VNmBhJnYadvVbgfgh+PicXf/tsJDNX7Ho0
hGr4zTUzIc1lEbG0yGKYt0yPdDCIMktkOCobFVinFCi1wNypuEAwr7zozxy2qSyr
5GNO2cqy/r1haKBCUXzU8x/4ioaZXbaX8/Z22Y/lPwniRcxL0gHo4EwmDQK4m+fs
yQZ8/p3t1+7sGGKzTAHY0BGO0V+dPiGwADu8Y0w0NxHGQ/9jG5ajk//d9MDDPhkW
VY1bO2pEP56+qfny27VThYk0FrVx0diTXmDUJ1VdODs=
`protect END_PROTECTED
