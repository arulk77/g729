`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF/fybG37Cr8/GXIekI5UxOEWKR18VIQaJpIBUAC/SQV
t++2XNOBL/rQ/yqbR229FyRNAvCb+8el/KdPCbWPKGibStFsztn801Mt/w+7DrrB
Bl9Mbrjr11PoD2W6YTHDaVuqg+XLvCRoP0w6V/torXo/hut1wtwWiW7SWK0yeWzk
JtKH4sIi2UtIQVNv7DIPy7CHFf1rkJCmy5slBKfd31gTMe+BVVTdiscnb07xwJte
5TQKOQ0n6vbX7+Q2w7ehjLeF53ecrDzaWFT8rH1VVyZEPmfkO20dU8hUvcUIcsJ1
zp1nK/ElzRWAODr9ZzPA0fEniH5E3CxHgmVORFV/uU/+UyVtAJygs3IitFVQ3DTx
eeh9Xr+v9SjV2f2spXwIqCKHc3yKiTbHkqmVnyqaAZU2IV9DBjSiZOa3CHi/LCrx
9e6Y0/B8nRrQp/K0HQv+KQ==
`protect END_PROTECTED
