`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePCp3LKuJ02yEAK2b6UMYYoVyIY7qdS/yabUB5/ipmvh
y7O0iwngfQKe06KePtplebXAe+Bi8pw2Z12HMPXnFOYrxMUj3RmVo7WGBeJzEkp5
hmghEQIrUVj0FpK7mgw++/MXS21gdvxHvs10aTs8mPEbtPnIdRYtA/o3CXxgP1xL
`protect END_PROTECTED
