`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJSgwuLEUO29aen1SSj8JrHHc33KN+eVUO0naY5QEN0J
ANtKxPc9BedM4UsKkzwhUgGj+Kxfx4EOPCN2hjFHu1NrBAxMHl+cjtTL2Vu3mite
nq5pYi5ReU2Eop+E2YKKE4Xz5gy5mZhSfsr6Vet55UgUPLjAH3QrSfG2awd7GZ4F
RpBSgLivycwir/AEostyY4o2bRfDyzyNZBpMp50a+UY5uL6O7fl56JAOouam4lIW
qwgVTySs++emOgvFdUXwyJ963Q6G4xx2Tp1TPFVjGs53rBxiiLr/VBjg/9YbECym
qPLZe5dsQE/AHv44a0qqTkxgY6gZleUz6iGGlxSIPK+IyA4W5BcVuoskTDHbAK4N
gWMssQaD3V/xZITQ7D/BiQ==
`protect END_PROTECTED
