`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEJ4GG3QPR7hVExH8vfa2WgtmCjPNv0SPPodHC1Ykv/g
4SQyF4msk84RBbMLwKv7+7vyx4FsvzS2/BILxVTqBbz+y45gsmlzGQNa78jEf23y
JbPg+Oriv7JE20ql5XdBLSOSF/YBZpBkCE7y0RTCnHIky1lQAkfegnXIZUnqreef
O0OTIWIAT3fJL8YKyvSl2nYmzTS6uK7xUD36HnCdu7PvPsqPEkVRg2VBPhlOZPg6
m0r7wVJ/uSQ6K7mbf7oAMVKJrt4TH+Xx27fthRwu9JXjfsg+LHRqCDsNzVawqhhV
+pJGtdEZMcBnZpb3WA8hkUzfvTKYveRPVSrstyslhNo=
`protect END_PROTECTED
