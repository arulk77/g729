`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOiDv9w3EjsV2JfiyXom8GCRGt3i5q+mUVEYRort63uE
PGhzGtp7pd9hVkN2bhcnVXLOa5b0v/tlGfSiscIgKrSYTDpVyjsFtnj5HW7dpVL1
PcTIh5spk754SlTDiTYc4ApoVUfbGz1IWkoBFLQF67y0Q4XcfiofOYxWRn8c7p3P
yIm2leHK5HgiDvbBecFCU7hz1vsbJmsxmfVtTQXJLKdyQSj/bwTEUoZkf0jpnY6X
`protect END_PROTECTED
