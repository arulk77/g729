`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ3Bgr6+JeGxm1rbNtCuQOHTBKmKpXjKR3HoclkjFl++
tdLjGuRMJNnpE0JRp4hCeOjip+FVI2d32+bVJzsLT7D1fztBbUquGC9N6UIurr/m
4VcKmYAYdwley7G+P+Cmv09ToJabD7dfUOwJAL21HWF8/DXcOv8FrgdE5NXx9IVz
6aUmROTtyJkYt6EDAzvR3she27wFAy3WwiNOPdFqs1FuZ23AHSnHNvSTMt4wcsvw
`protect END_PROTECTED
