`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43CRbzqAZKOaVVIztsJqIaWgZ7a+zIvYuwTgEGRWO4vQ
BmF3qRDTRZhfhaouJXiStaJAX/Lt4VkvDIPGRzcjvsuLHADNb79+SeVyfcHWC9GF
IWPq7oAzLyn05lIf0hpYmjr3I4hww0waqefXbNwm8ZQr3X29/1lmf2YU2KYuKkA1
5JuB+oiamWK3CWEg7cTFhoNKBg6gVfN9i5EVsaE5zTcamk6PUcMSGQzEHH1nGW6H
RLSC8UnJnKaJnYluucicpAnzKYynIe+mEtfdky5SDmQ=
`protect END_PROTECTED
