`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveML35EWwlJgakgs5WR3O5aGK/hAS31EjhJeSz20+3Ft4
IrFMenGkcT87deE0MPCk44+Jw2rEnkVfsQIlkFUg3eU4RL4x/39krp+EhIsGW+KN
kgbeAZUUEMJG0YlWpThunO1U/LpooFPMgY88BRPW4jBimLVXFkMHKX3rzoxu9SY/
eXW2BjYPMkN3K47GyU7XxUtnvk7lEzG150jwcRV63KzYmfgesmQh3n7X8ZGF581y
AjVBw2fbt8r+oDR9mhWy+GoOdiFJTj6kVJkt63yOG5kiKNi35r+BieabsVjTyaLN
zj9VrwvNa5K1tHYcXQj4/aHQGLXoLyscshumAN8SxGiNhLV/JXrC84hatnRbhKUj
6eG0Dk+iqSYH5NjrU6guRJNVjGrbDe0InDwHScxRjCBFZVXoMvp/MXlS9UNRYijf
FJrKafRA0L/Cq3jRFKWx1qtHd/ORhTf1G1pdCX21sCERONz0/R0EvaNbgRIG9fwF
GBddvq1OHDKPQhPYsatH90LNEusSAygFsHoXgSJQKu/hp1w9newokMnEYsv8Vrx7
YBW5RLR7fQ6e8r22TYT4yB5xWaVEpKrUYLUS+Fn/WZOcmS+3/QGhzn4B5RmqLRt5
`protect END_PROTECTED
