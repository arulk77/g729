`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Prgb+lMGK4ankHVaNnLDqw1kDvzpPFjtRlxCu5cd/0vF8T5adpdm9z734O8Y2ENt
aKiyK4NN3eLbKRQnL3mNZQFnCFf8OJ3qmIZ37R9r+W0gg2xqcl6bGsmiQgm6bJvO
Nq362byM19+/6/HvbXRkKUfV27hFhSgXwWulv4t92C1Czc0YDvbP6xf/XT4UuSR4
MH9D/oF8x+KWZPmt1074dpF9bX1TdjJF1f63h0y+7gpknQU/cr6Er0kNEcFQ12uq
`protect END_PROTECTED
