`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL8/HuFemwcyjrtSVR8ungczBCHt8LFb+5uAdBaagWvwWq
LKJxA8/OrWHDszOLlwzN+0JwKsCkMYPIaD9ywpLQ6VL758pr5cpv+7/wAzKuQiGu
pQv6oO+hZPgoigQ9Xj/Ho0qX5r3SUPReoYrrw3PWf03BNv25FxqmlCILcFNp4tjl
+/hQQkbbBAslCl+w2uM1Apchm47K/hQTDbz7bmYzDF8PqdYPssF5NG64Sho3CUv2
Yv724cuE107u1f2un4cUC1wUJq3/4Navwk/YBtC7t1zZr3NWceRYJysCroFXCnUo
CWt7X7zuuG2JN22/UMNkMViG2S8nqi5WDG7NtKqi4rB5aCqZl2aKcA8W6SKKcAbI
XoaMC/knJ+WPq1cdSr+z9FBfmGnjQJb3pPWsA2TALOTgbAZ9h1jaM0t/k/RABsoB
u4gji7hX7WVHviIHjWKh/lLzFk/0Pu3hwcyI6ySzbGQpAQN5bGvXj4fmx5whfe4J
wIdyqkbQktG1AvX72TFl94kb05pezF6rZNiokRb9o4xtL7AHDtHvePEkfmixGkXt
a3zrDfmxzmWi+qO+JR/Sy5qdSK8vO7xcJ28oZM2MmmrIzNBJVRLTCCnvomU9fQHA
Qq4GL8paLSS1gHn0DZGQhqyBeU2a0X4yUXWrbRXpPoc+3YvtSaQuwTtenoQye+YF
SyGTh0qR5JwXlWoXbn6lKr5wR9dmvdy6dOs1EEfO1xxgwGAdrfOE5c/qM2PeRig5
7Hm7hmgv5fl0Iwri5pukZ7YPeU36sPVhv1TYnJ7DtxSlq/mlElUeXR8wnY/Sn60i
T1ANlRLQQqNp0TBF1+UH07yTl+zreNNBSAVTRQbsTeHnotZHvX91jktV4JqIad4t
rLR5tfegJAgVmg9kvhVztVo/cWubb6g2JQiEIY1JRK2eU8No52O+CQNBeW4A/Cnk
t74maous0HzD8GRkOVXbdj7FRf/yM/5E+BMlQuUa9ptaa1X2Uj3HB5lNfldPYLWo
YoShH4oPT8djQAXY91TRLSoJLXSEFOnupD34DJZFZZmGEjD76yU3f8A3XNwW+3IF
lL6RV45ftirsOuslBYTf+RuEBd5seYgbdm8Cv/oWLPpfgkfMGxM3aWOKP8c5kZ7x
TtOlnkfD7SG+Z90I8NwYublriIOTbU6JWGMLp/Dq5zon/GOFkZ7jEiD5kMOJ5k5F
vK8o0HJ/UYIIUEHvIAMceSOfMKs3gZQZVY8ptWtSK/NePQX3vCL4jfoHAX4nTrJD
3n/PCgMH6+Oy8XaFsI9sJyViiAyVAu80ooCKax2PHzA22HJh5Gw1I/udiaXQwf0r
w/+i3nhZccV5q2vaqxGmeRBJxeknxz3xDWwQLx7GUj5mUfoNPuSfDFQgtmXz+4lV
I/G5MV+7lH47qXeW3zxe/fi0aeMuRCZLEx1YGBqSVy8CCrjyKsfrbCRKoWIAcQLM
4rTBL+zBo8kbAL6gQT1gUnvkgRHhboJr3SR9Qw3lOjyW8S/gZO4czacKPHC2gPcT
6Piu+NfLgdESgC/gt74KRS7pyupP/fduU37Y2l6dO/tF8Sb5wcfl76PqDwu81Vuf
Q3LVZmAaAL49IczCkhPU8bclDE9EF9lYJyLbE+2/MaiFl4yHsjRdwzkkPP7USR3H
EvsmBBB2BudvjgXTfp1tR2YTkNYKxiseYNAM3Y2fJ4R91l/Mdf737hpqIg4f9t3r
N45haRDyreFV4OvBxIwmRZiWDgk6nGx+BMBrlXuU4K1G9B77XTMlmMxc5UScOIPe
IFavbEaWZsmNrAoLgGLSK1LGI/sPkSuKwlBUonq882JJwAzl3vq/BSnCulst8OIE
sJ9eSuGk+Eq/eC783HA95VxcUPg5+spEMkF/xiqKO6bIin7r+Y3UIgjkZKRUpCsD
zpfQlBuezVWHASKGGxstXuP9LGHDW4Pdh2TVXA2HxWFhPOPXggTeFrPjk2jZE4la
riigvSGmmlxlady9Eay9CkC1bKk2Q5jBPgJzChzAcoXxWVxa7t4e27njP76tDQ21
kz2daynu8gDtQvtv0ANPB5w+KR/r/sm9CQHcxduSCukywki6L0czmgsCud/SItRQ
hsCcdzYrOqy4uBpozeKj+IPMED7rgPikREvYarWSUgB2E6qST6veKE8Qpf58ldf5
`protect END_PROTECTED
