`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAe6mDtwqSxylXqkDZ685g5+Zqsr+kWFCo5mWEzMsPkKb
qWGeLQXuxOH65pncZnOkoaSUahwwWn4TLOXbGHLgi0Q4qdQTOxSfS8Yc0MHxGeCi
IqkGDV1OtVndf85kMVjrTzM6zmKrJ83zLXdusP3a53UsXDd+7X9l/POGpUIDVz9n
HeeJC0UqmUJJCkxJBWBcBZ0tzqM2usMRHV+AatvjV86mQXbTwHxdmmHpLECQ35en
WS366y2SlMOMjULKCUXjw0aBUOnHNAEYOFb7FxqbElCcvcj7xpeFlnKxGE8Gn3Yr
ggMHQEyXIyttURgGTI+h+iKKB4FI18oF5l/t7b7ybnqOWZmc4TQGsWJpKiSn7Zs0
gm9mksPp/my9Q+i4qkuZp9d+5WdEKpo7zGQwYp5YoSIEQ19c6nKnQ4Am0FQ8owiN
zu34t8hq0N9vnUa5Dn9QrVGxeMeyVlnEcrJVbRM30eeHE4SWq7MJX6bOLELTBVbs
tC7DSXDMI7iMbmM29TQJZQk8RsP2ADU2IL37EuLa5ErYjEIyZAlvGUXmGFR/q0RA
yFAjrHtyCEb8kslw88XUDWzpnusIFXUytX3TgUEVAg2hMfDkYw1i4ABPRQ2pHqCv
l3ooqYDJFHK7ySmHthOQ6aGWArHternbKTJ8xI7TAdBtfsGW5j7kqF9rZx7+Ouuy
jZbJHGaKT+15y12YgzQlgqOjPY4kWr53AukiHCBFvbk/ffBqn+mCYNMm7sOahOTd
cPZh50jufChl67xYt+as0bszMonaihAZm/KJaB9lvaipmjxQGb6TgCIKOtkeeL87
hpKukw4GyJFKOfd7106iQZZGychyrRIRxts8EVVEvh306H2apOql5Bk5OZE6hdx3
nMHDg5VzJMY8KYc3kJ0Sy7o3ocI2hzSiK9q+l5XmGgnWxwxR3cQR8r8MJsIF3ZPp
JK3LJTRWRIyWpRSuHTcZFFnwGM+m7GmihBElGmWFwmlxCHal3407l1wd3cUpYlBV
aAw0azvH9udLvuxuMj6A1xknQ/ECqmdj3kFJflure6u19m8QORsysX5IA3+T/utQ
P1rJMvHkawCfeI3pxjWO99ftPPVMCLb9bSCbJKf0Rz//nWWTqDstIXydm21ZD2v/
2AVg8Hklmm0ZQs4DIUxbjM9hg4vEoFlTprX688dChZ3PV8Ov2SE5N8SuJVSDAVxG
sJWDCajSrXF1Phqf8qEGTztCDy3Uuped9aLzIm0lGCpaG4bQFqdj/aOqbEdXqins
tvQtQm4v8dZN4zI0I2rjjtX/Ob7/3NjGoNXzL/xQdIxZodAc2O8MfQhWyMm2KTtU
HqmQhCwgMDjUoLY3DNhvYQb+filS8TXU8F7TXkMCCTs3cUv+rhL4W7gUNN3FxghZ
wfMlF7M80Xq0evt3mDv2rCXyZueRM8tBfcjN8EksMAHNAMHRivZQ4QXqlt6O2BXg
Lwmb0feag7rJG+fPq+b4Wrzi8bi/5hOWwljad13NTRW3XFpNZUz1zrMLN1JFimlw
Ry8qOFXPzI1CaStOTD6UwG76bt0Vmoay/Rvi75lSKGkcT03wNCqLOx5NSfL0YFex
00LNVPVTGlx+A8aoXOhxFd7ofvzUe3zPpkogvlmuhyWXU8/OPxeLpuOrLJnQW3Q9
5g8dDhELzss+hmJ5zJnueiGePLXKj2MLAu4jYoIKwYhBDvQ1ayOCaGlwZkqBxwYM
TzwauvX5Ln84m6E3wxXuxSn9rfnx8evkjeAMiOv0jySn2cDTiR9OeVrQBz4JCY2c
vbSGIC5WziMS/KtIQePCPP/xWuuqlMRe2x1qi1rTUivv+e/ZXehKBj0kcww9Zmao
KUS29bjKy7X35mc847Kk+c5qlHeyo2SaloKkS0Sq/ExQvWQRdLeiIf7LJPzpJ2Er
7Qv8OUE1aH6lU0X5ivF2xqrEIR5mYgYo/oU3MfisSEefO7QzVGVtxF3ur5eFcuXU
x/rbh13s0wsr7Zpmd+nDEInqW0NUhPWrKlfqNsAm4eIbkQt3BAD5EGXFlRBwq2BS
Ulk4trYtYsYlSQ2MiKNP6ZjnZ3G/8ngAcAYWDpGtTo5I19nmwJ3cig33DURbK4p+
j8y4jJbDNKDbCHq5MmHi8Sm4D2yQ+QnBqDDn/+R8d7Xyc8K2y9I3JsyvU5O3YFwo
sDwLhwf0Kgdhy03QpYLLSlo3bCZWePbYjFg0Uc54qYyHEhMghAqu8FT+CGULIOlV
IRQ+SquxbKBEFmjvZu+fyh2DJsBQuAicJXk7c/8UKHBVxQlIVUtW8gY2/9ngsAIe
j4OJg42HxrzTMo7mmGJNAnMi1gjjMA0MWnVc1xJ9RODpf8VGsH40EJw0vIDftXnB
Oqse0PSXpI161DfxNf8ElX6ETuz3CFZJzFEHW9NJLyALM25hoyLMwe4GIpcZGUPI
8ozKbXnpGObeDfgl13Sdyson2UG2z3OfpO/CwQko68ClJFBKesyibSa3bMvvzzIs
DQquwPVowjWG5429LyZsUW1NcprM+aThQfYlC2pamossnLKSJDwjGM/7vlJML/J/
poBw9qvdL6vO41XjT92VGh+X8qF0VbFzjfU+ToYkR+CObDoUCRUpgg05OCxsgHz7
91S7g0tygGx664dZNFFULpzViObq/URriJ+xK2U3Rbw0M7iVc3BLhwZF3e8kHwKt
PV7WU/jVGRLBk9Bo3JKyDTKvR9iZQWw8wcSaY18v5cy3zdnaO/ptm0tXzfxcvlQT
CJzLNwsyFH++OtmzTxunmq9fgDtAa88SCrnfDiWCsMQuJtMmjZKMzwKlHRMAgyfi
kIWdWLtd1+rn6vK72/B26GOF05oA/2Odd84h0dy1Ljz6UIleU/9F75F+/8KI3QFf
LFrPo4gf4H+gVJr5ajmWKeVWA6b/+yxT3wB8V4Mx9apSr1WueKqAaJwuBdau+0Zj
3CaHi6rL9n7isG9U9KjV4HQZnxW/kG/E/THA0gmikGYqeLXM+cNF8pv5U2ylM3/r
Bj/vUFvGnglgwqcMXDWjQrDCl5VlUIfwRQyH2s6kTmyMdYD+DyHzZa9JESa0cLZB
t0LZVu7OV2aSinWDzvvXvWtm5PenTIJ4cOqTiJdfC9epd3DiUd1PxraZC8XOjpQb
hLgD4GRQo2o+OCymBdRAzpvxcYCBZ3zunIpF5+6C24H6ZqLqPUT68THBiXu35z2e
SK5g5eyBOI/z6CbjYrIWAsA+eFH5AfR5AEo8N5k8wHmsl5VIV/B5sXzP/RkXKLt2
BUVfRRloEkXkuCFwAo6ryUxlk+bdiEe+7NnG27baabaKz3EE7oyRoKQBYEJgHjbg
+bLBikj881MhFR3ZkGuik8VgxmaM6OTGIk532naKYMr7Zq0XqFwO67k6Jb9Z7ZHz
s9hPyDMzZrT8O0wmCesqiCqGcsZGyduathQ4tRf4o2ntAO0LVJYT+ESH4+GAeGtU
psm3YfWcR+IlqNnQcFDK2VJjlucLrjkuqAB1vDgI3Axu9BKsSChpHlB4cDKuRW0a
aNZXE/hRl2Fy4h4hM7kkbl4tS2RVe6aZ1Dfdsj1oRaLy0q+UmHHUINehe9wtl34D
QbAYc3KZiFWJMHyDZ5DGA/OLMqE5JCziADQBMjT7R0Ue3VzUciKFDj7RSOg6kiql
eZ5lnqCoae178Xjo/3P/YcFngszInKJ421Bd84KHEznSoL+IOdpql+ykPK8iNWq3
cq99BbTSEFtwExOzv9YK+ckfObgZtaO+c7FjNzMJJ9aTf16IXWkF0683UAV97Kf4
aPv+yp8cRohZIkokKpaB2GRgU77gauEEtpl3cuHZyWK++Gi5yfxKj8IyYc2WII9i
3+wsYKZ6DjUU2DVsEdQYdYsGT8oHohhSWbV8FVrw9+4jx7ji3Vqng0uJkdGemCjw
VPNOtJFP3ecdrlEkPBjFjsWOfJi9jq/0MjZY/g0obeNeN2lQsh3S304Buv4ub60h
K+y0hqnYbw0Z0COhp9UUr+RzOq5fcgt/rVZiFCVqMKk7U6OHQ6HOMfqUrlUx/MwK
yB8jlbIPWkuY63MM086Fl9tSHbkOmwZqXCAVaDsGGErcMMnI1KjA6zt4YRjzzyb+
RG6cL6dqeTP2hVq7Wn+KR493xrdGfw4s/deicWDTDrfX2RA+hqniw8gR4OvkhTyD
2zdhvugElbluv/JjG1qwUwJTt533wSlP1wGgSEZfRQ9IU3MbRCkyDbWlnB+RZwxH
W4boiZk3yXYr4Ni54Gtg6pVBAiRkL1Mgr5RwdbE8KP1O840emaBsbzwRGtzpICdH
mmS1J+W7rXdnmHT8Yqmz+9HkRneDDse7Fi6JbgwtyTjIdIg5npZMZ8/BlW1Bg/YJ
gj/1xi1hxt68OdlTCa8ClKsYXDa1LzkXivglvtMh4gmvJFeEM291HxsbYAVl6Lf7
9wU7OxZ6Ahe4RtixJu72SuT13NWV9sQ/opUDzDNTBU3fW2WOsohb7PvP0PfkSyoS
K8k4dCqyq0jmruPS2VDKgYK5Pr9QoLz9lshqG7ZufQMeZN2kbSyQpQ79nZgWIO1K
d02s6Ts1oHiHkodmKPX0LHb6XrtQats1z6dt0WNg3s7stusgf8B9SdP9TeyyDSSN
wzkOm+liltEuk2HRgB6+/KmshZ5FLeO4rEfqyUDnpL+YuhBJGiAyV4oyx11Il3AX
xSOfJyK5vuzMerqKkNnWMxigrBzyiarTQ3EMuxj7uoZmH5HRcpdqaxjswmwb1P4p
rZcjZqR2jwQ3RVPSb/+ztXVpcXNCQJlHyLGcjfz9eN/jtCRnlUDoAeZ7j4hHhz35
HtIdp9eNzDQ7pE7H0u2Xcu19NOyejHORgFoOK8WrjRWJAFfEut8iQsNqh4MaNL7b
NmVC7HlcXgEB9SFlneZMgC24wyldyRazN3PYl3/5n8343Xp4mECAMvLUTNZ3jDNC
S7Iju8AOGecPQP2+KFtadM7gn6FmfIyr2U6R/NRMJE51MIbGPyiaSrNknm2Htazn
X8vymMCwUMolvuEyqRXiXmhwwOBkg9AiiUDe4LIILhrb6Mq2YvknTaww9y16hnPj
MqRSMiLfhEmHzukRqq5j0NTHWYFdMyPKodKg5BMx6xHbeFkmNApSpz12+k0Mlwq5
UzDhd2ZqA36zVRThQ5qOeSiJjpnYYMSP7rhlako5TzCFbOdk+Cyf3wcRWgaihk62
ANeUoU3ZH+6pbRGg+XjF+7fP0Vkg9jeS2sl19/ZOSfgm5d6x3WF88wBjAakuMxVn
21q0V+1NG7cgE9jZcEwxs3U0r8XNCO0GNH928yPxsE/wi2rIDsYufQrJF05Iybjj
FN03J+f++qM3tkqNwMIAiLXwBOzPm7R6qOSlsBEx0wAzWm4C0YEomZRIBW1uBE3U
UMcGnWBcuEhwcamL8WxqTcHw60Tz6euRZvTQImDdVzXQIzgBsLjl6CU9p336ayb6
bUOOct7zDUbgwhTGjHwuJC40cSkSBElgoEX8YfuxaSH3eF49oGQFXrfvAyNL2RXP
ntFbT0KA49xn2W2j7yEP9qwkttRcmzzbIVU2IYF85WUnV/COCgn6/oSM0mqX9pC+
AYHoEHj9yIPLwfNvUeXChnX0928P9slYQFARHBMaq7awQAZCxc1sOQmN498jvFg4
I+A5ZCkCUxpMgN+289E9aYw3VNegP4FaJb4zYvCm1vCE3DDD5d3koDopBsDpCl7l
tf/WPz1QWbYJgJuULsvprWNPU32KrTqWpp/pFNOm9tkGpYHnLQv0ymnmfc6mEjpQ
Y2HvLJI0TR5QiMFoHY1Kb+6qen2eFQbC6EyehBgnSk4Q5APh6HgULQtvMBTK3q+s
asa48wDwTKKKvZL0aBArjMTZq+GK26NGV2yVT0gpXNzaP++SHHcGOWEyIVL8Run0
djQyOnIjkAR1aNkeMzu782ZXVMium/J8f7/hNgNsXO4bN6e81T/yFQMCASf17ixd
WNASEWb1P5Z3Hf6Z6ys9tFzVA7SJqDYDWmnwIjEDW4XnG/mfoxrS4YEvDI6dNk9o
dP+0BAqVOoRbdwda4WTqIDGqpfhxKn2f+KJD8W+bFv2/0v370/xVegAYQmMjhn+G
1XWwXIMIi0hjfnkLRaSa+EZyzoWnosS9Rw8yLUKv+8c24xbH1MLs34HeBp9jhRex
0aw9Ufcu+k87auSXZfP8FRb3VVVyqIBcnsl4bw5+ZdRqXaR9jGTWvmha7pJYU1gk
6n1JYmMu2iIdic9K0WREuyb0yITvfMEqtnHI+bo9OHIRqceRYsiaG1lumG0aMtfw
s24IrKjc2flVcVPisk3jynLR6LnVkYUVufs5ncmDVXFuXR8d+IS2QzXxZUTeKyL/
98YU//I7egK8HgpBASwdcqx8FwMKQ5XPENbv+EN9h7hc7gm0BTFMibxc+Xw9vnMg
uG9Vkj58W7/C3SezmZ9wBj65suLcDx4fye70Nv1ptBfbRMDhdArLxVGjDnH5+e3y
t/7prdH9kdfs+YBAPjsCwc6eiU5iiceGv2GoNGu875lKo6LAMvhY5ald8v7Ih5d3
PYp/h/BOSkMM7yKv2cI0u1lWU2j706OXwR7KwUkA7lUf118sqk7Rk3j3rcIILuLo
Ht/0ymIZ3n1/lVx24r5donHgP0hnVZVEGa4A1pV8i4sOT9bGLLjmlHZc3S039uLd
jFewhpQKe4pySKcXFC/mQSLycZirZI5WhSK7O5+2ClOuVdWTXWs6jXqg5lrqsQ3K
6NnjHXcnMPUimOkP8FmrBnYofxDlLDvgToBITBnCF6zuOGQwcmubQ3XFSC/E1OQ/
sCDB/METpTyAPE8Bp/BqLwsysY8+GrZ6tGuVMpXcaWGWn95pnL57Z8C1wbdoFCpw
xLf4uqhZ0SzD9yNmczt1+QxBhNn5zn+IxMzI6JYxuiVF1hX7NxA6ZWI54DwI/rjm
n7SKRKrmod1jtvjCU/1WRGPNLePzD3toXZkXwUGxEw27duZ1Won1pxWzPq5J515t
wOS+3dVIGUZj+JlXf90DFahmWvR64VLmEHv/MH6kJTnblgDUN7uOFuJ8eHvlIjQm
jZgljgjrlb2OMvFxuh+VDDVIPQbTNs1tHN8aqQK5oI+7d1eRyX+ubUFzvPBSTmnj
hzolwI2eLHAUwHNAKkpUU6bzzI7U9ELHYv0LQWrQOFk7dhC/OxsdCqqaFAG7Yxa9
MZSngvogSWRnvHpXhgtKzaQv2fryauVJyI9YkOlKbqDrdYG0Vzha8F6WdkwObI4L
44TWD/hpcyNy34POFTVXYq/ivPKWrlIhZfNQjQQbptZFNy4agWAiXbgxfpNu+sZD
ZI0G4fWxErbgpKGxSqNBL+9Yzqa8ZnuYZ5VEWz6N99cvv1Co3IQMX8hVpZ8DqoSk
InisX1S6cP7j1OCnwLyMhNRq4XhZ3/M72yWld4HDVeJxfYCiLNdFa7qMpQkwhOg3
ifkPQhcj6OlrrV7ZcAlPA7G5hJ6Rg78Lp0oHuzpsaNrSqXgIGCWh8QA0j83/cas4
WAWBMHZ3EkgKRIV10OoABHDBH1CWYmHVolsBgmMn70cBsfTRH8j3AlKgp89jCpWh
Yp14sNwuzFY1E0xQVUTHbgACcXat0I7DIU2oZVFSGjZSht7di9XCawYg2Tf9mRLy
WholciK92Y4IZzmmDoKLyMPpLbU4X84TTmil95YLlr5Mkr7wgYKhzJJ8rC11UO8Q
Chq6A9ClKOU1/i1fG3HJ2wV5zM3Zb73Trtq85b+4TBvL7uQMu2tPfiVqMiFNL14b
GJ5++/U3PxurdQk/KWRHThy00RqplfBlXiWwraDoK6cc1lWI3XdlHMHToonrL4wN
cjCzL3z48Lj+2HqGSE39yQiXthP4A+rzThpasz3a6jq/gGpB369RFokRuBwerZED
OCYHtp0IenGQLifDyaThckzHGDshNtED2iD9U0NjpLvr5uxqh5bgXc5eW77e1ust
ugS6EOy2ukoXZPjcBd65tFNsDCMHOxKFut69Vjsqmt6KakbJnU9QWx07LDRmLGjG
2ht8lY44PLQA/zEOXVoiih29DS165wTbr1CDUfgao7948vx9WoRU/WU7cJBmpRJU
jP4LY22vWUIzWdzpJcErCOskSF7w5F8scnKhBbga3ehDRhOHJ0mO1q9DUtYRnSO6
YdHmaWEigr7C05W1Nx4rqL/DaJJz9WoGIiYJ8nK368Nr6hxaN+4jMjzYXTVip255
`protect END_PROTECTED
