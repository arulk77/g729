`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMWu8ZwouXqH7Ch0X2gpjfTn2sDLbz2IidKzeBpnZOrN
3DGvd7X8/wjGwB8BkIuV8hrXzOcELkyq3TC5pSuxdQavun0ayVQza2mMR1cnNK+X
ELLSN8U70Lxq/0kZzmcyixz+WKF1wDDd/jJVozjkBsoNkEkJ7sWBR3rTUXA3u1x0
W/H6XbrG8RYHW4Se+685pJz+kokTBFIeGV6vIkBFmXM5BtBXGzLksCL2FpKhHLXV
`protect END_PROTECTED
