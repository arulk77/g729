`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN7E6jBwuJS5LZUxRFKyJMsZVtNycwKWszg++9g8cHIK
cGgS3xuOMW/M/imB6xOdY4vo+YIsmYE0i7VlrKyerayNs4/jOeRLBTp/jd5xMNrF
fvZmImPJy7JqVKj7iH/VOgreQobRcaNwY5U6GIvSBeYmwJOJyDw1378JtIDFCBMr
MXPO9yHyoFtmDb7S47ib5WwKIb7NnT2pTU7yd1GCh2EzVLvKpVh8Y6bCuDKSWk4m
Yg3Xy8V/aFAi3HEwc02+E2ghFi31E7q5RSzy6pnCDqSWB4DmEH3m7IwKD2YmF2SQ
aZhdgU/vwKl0OTM/AD5a8Q==
`protect END_PROTECTED
