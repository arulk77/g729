`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1abExSeQ2G9gBIvWHIfcoNpNLLBarT3ktS+rLR+a/dTvc
3JoEsq8r5g1VAiwC1C6cQYy9HAkqt/tjMEPljdEbG30ljFr2yrOJfZYbk04SQ3Xc
m88zNeCfdW/dkK9LNFZD9W3kXLLfc89sFPxbUnZjZXEAXErg3j1foYRND1kL+3fh
e5/64CGTbq4Ve5/JAWUz4PIR60mJs+lozoo9D3NIuKsxwWwVAakPz9LbrmusFlOu
ybYbrz9pVRZ6O0FPm9cduhJxmp4wqnlVJby6eWfRvRNE/AqaLo5FXozSRJtd+ydy
EamQcvPNpHGACDf9igjA75bx07BrNvaw6IclyPSKwBIr9Gu/92vyyAw7E0vCHmCu
tDCj0LhF+UcpaWBIghFYhaFiYDuQTXyxXw35yPyB3DFNJ0upGVopKcFHNfGLKKC+
wmaPs06Y94LUSfHLnucLV49V8t69wmrwcEg2kWj9Y49hnr9EV1PI8YUqnFFVxfmo
4Gz7RzxR6ZH3GhBoQIIVBPDO1ah+gstKxPTbjQKa0AK6JBZ49mbLZAYAMtBEvod2
AFXjV1QT2OUklSii2GO543V+SetysvKwVkXsz2ZqG9GsEoJ4uN4uIcom9b2Xvbge
lGXGxXKHIGaZmhXM1KlLrp2JDqzlleVcz7e8pdvgtT3dN2TqX6L30QcriWJB35bh
DnOodFMc8NmcRwvbhWZSWB74TszSNenp2ul1ED30NXeRBWddQg0saPGP8AIbgi4h
Wkokmjj9YCxhOU+AlZ0ITOARTvDvBxXZBJ0GOeq7t/IJd8ytd9pQLKYWvpAAx1H0
BBNs04jCg9dKGtCydKx4+xr3BTDJjVTDLKTzQyH2bxzWaoClyKV2JyRCB4dialCZ
sz+ZuFSaOwN5QBB7b+pVGMAUtRRpZpN4FdL6mMIQY+em2FSsmnTLGxV+0cbLVtjI
sqwVymaZCvt1tkzPvBFTP+LI7QDrdE36t45bXNsJaOI2MooAmts1G3yRVc0i2sj5
1r2LkrN16FFeCrOE3EKI8LjKVQy5C81IK5TYhMnmYJ/jArzoELIBbObYBlVYgDYl
klntr7ywDiT47U5JfvBurW0IimHCAl1I1N1EgVOA8mP2FKUyBXFBnxwtx7BNySoj
g/QsnklSLgHl8C8WM0/zVQd0cv7Z5PKnCBbCxOtdLC9S1HxbqPt9+W8WdObL423Z
q2QcZBXByfOFwT5lFKKoHOPhKGBYYx13jm3L9vDCY6RP1aiNzYwYUajlEYKHGJcJ
xo7lLuerOiAbojsAQi0KQX71FwlRmldl80OkTL3EbtD8984bLTNEuW2/ik7LfeWW
3orVWrHWqxsc5VF1MxNqerQ7NtxbMk6pQeWqO17DLn3nLr3rccFW63l5gTdwmROD
yJiUYoT0VDu2FiOJA62SkP1FYZwhNzC7lpVwZBDogWx9JMV6Q9QpJEBXypJlESeR
ioB/9X5uqoFGlGrMzxGqjuActHbZQdJdyqT+ZBr1GP0gfF7cMh6XrHYVwlgGfTg7
jCVrmqmKn7h7uLKnXDcimDP89ltNKNSDHEhdqNSJ0fw8eKDD9nA3k+Ax6orlAoyX
elYgo2o5D0qvz1NGwgXSQ2T1cmhXQKNzk2QUoHEjVvLnkTk1XzkyB6CXc5nkTLAL
uemnudBEV0J/1EqdwwVG7vKsEEvmbKaH9r7CX/CpSvBBEJDfN8TsgvI8AvS7e2Cw
0ByS7+cdouD/1B8tSv+uLCMXjQG74DnF+KeST25dT0BahyiBBs0iUHUW9tL/LRtk
lVjPCqKMv3RQpVSRkbyGbGC2o3qGVg4TphMT42Kn27GclA4vDS12kGSKhINdW2VU
RxsjaqIJSqpEYZnYrQf6Po4+2jNPRJrf6V4gvucRWDRoXhIVmct3Aw7NGrlVUWWM
M8oq8WEDmemiRereSHUmJcHi47UhWFAz6ZtUHBsDT5NwHDkx0N7x6xI1BT67qDqS
f11oarOzT26nF6Npe1iQWTyy/Ddk6WFj14hSF2xdII9fJjohY4j1b7yeeAhsIaZP
y3BB7EmVMlc5w8zELcmMhuQ8EUyKY9BZ/iYDMrRtVo2eBNdEyTfBYs4rQ4s+GGJx
4tSBAFP2hqRJUapxC+nAZfrL9oBUUMQXQUABD0t7aphFqxiJa4wbDdmUrzetSnyh
fQJrnB1NEFar83FU/MaOMz71Hnbx55tNx0YqD5xHCSXkSBFZMOBrO3ZrfJKwGvPx
wL59nXtRWvMP3EzzjK/2g83S7552aUdCUkuBcJwkE5K3ERfsp8Clh93cPKvBY9Gz
/c5aFKn0MPgGvrG5ffusCDptu6HwjVFnq6pwETUoIrKF7IJrClO/f70ZvxyUqDv1
Xv5quhxbZTpERpndxtNqysjdabctbYT0doRSpwj/iMk1ojxNRMiWdCLUc0jQ8pFc
NSknJMQQpj4y/+iXgK99T288b6TemTdiDaUf8u/HnDItQ9RDWYOo0heh/NHe1Y7a
4QuOVCwfs0vVUVxxVvcsTWs5e9QxNk7Yq06HOgW8fAT3uRDEYTNyD9A4zXxAWFsM
/N4w0rHbKXOSxnPva6WhhBmvdm3qiPbb81IwgUq1e3g+weGSrHI+3WuFmo2mixXs
s/nOtyvdlgw3+lHrWKA6Fk/g+OBMDUG3ktqA3KtoI7M0ZGYc0zjlwpP7nrKXEtrZ
yjkcY1GrqiyYOgLk9lGYPEbyHcyG7tVKSwxaLnWTPGIBNnUo36t/AiXxKC28mAlL
7z2QQcxO04i/TkozPyuyF8eUnVjcb9GR83ZczCvLetkVZpODgem1D3kTqbmO0/Hd
yxY6u5ER1N2sK5RYEG/vK1ani1xHT/opfM6bmwjMGK9Qv5bParzhypBVU0VXM/Bp
3qR3mb1fclwV3EQzXOIqGBy2SbqJNXDckOg+/O1bnxsLFDNI+5bF3+QAmg8abGmh
rG4+53dbxTM7FceWzLhuNcBxuG95BhyK2vuaM/64XIPgp7B53QbaBQWm3J56zUew
Y+SPJ3uYKIYu9DAb2Lwljd5CHRaUa4QhXyGxujWGudnkZpd4NM3UUGUsfaRiW13F
H13eI++tj5+kscaMzoNwScGrSLiZo/0VJT4qyXdt8ZB+/2pUqtUn1e4Fa3hkPQKn
zoNwXXdJFiM0/zIe/vfqR7zY2CTdYq7zonfEOgXCgZILaikzjCZkpWnNVjpv15mw
76oZ48vbCguf1mJgdtKzQPoDJbDooEjnrzRqZ1QV3WepNOcYwK7qAHarT/4y+3mH
rPfJHJFC52hgpz44i472TCJ7+aYUDOoXU5rbwRxTTrY/+iScTGrdDxgE3mCCS/3b
jI3iTmDWZyMoQjFZy/egikxVJ6Ak4quaTrR9j5UBDb+jrYfnCcmCOteJTTZFtPwD
9O3Cre3BgsGeCkeQOvsnjBQEzFScnRR3h3aUQbJ+OhVqQoK0yq48JFDvn4A/w6ay
aOPXB2gBsDvp8KpBri4bmmSpPQud6TEcmOvinjj7LGD9cZ2BsL7EA9SUk4bEa6+f
VwnP44RkzA6oo13zy9mvYgHX9J9kroJGyTBMyChGdLFNWuluHpF73E75Sm6Y8hzv
nq4J4ar59tVM0p8EkRSW2SCv0oRD+uccIyOhV8cgtooaGI0AOxjnqxuGLlKETse/
sZtrpca6KAwp1FGzAY+vlF0tC1v6K4Ml1blmLOU54rPO4A1tDhUaCeiZB4l5n/tN
B3bDX9jNctGXtEYImBORMmh7qrgVSWeYd2/Ma2Y0MWEPuKJ6GboRE5YeRK/AXIhZ
WazrKXmaJtVzQ96qnSzGB8XErfzICLOlGm3ykjf5wHxSlyGSbW5+lfAsxmZZR7Eg
6HsRg8vII/x00KS5izDqTxKjVnKDL23Y2UUGvEjL4IE=
`protect END_PROTECTED
