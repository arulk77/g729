`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveO+WdFM3EUv7s8zouHX1wF/ay97NcA+YwIW7yXimLUAu
sYlRAVBGRd01dQKE1uIzuy6z6yN+xD++lfiKMWWPue9ritJMxgLPDtXFqV93/68u
gTf3TR/mAcEkK+BVlHc0K5w4j81Kgv2cnpUVEvfEY1+8D6J0WYxhrlFTGOUXWCWf
UfroFqcKeDAmIFej2w1dpSyC8on7oeJo9MtQdlIyjSJ/wJcgTQ8aEmuZYDmg4n3H
Ul74oLtssdMHBSJhxZkMgvqimIPxFJqbVDsjw0PlZBGQXYUZJeBPEpi3RGYmvjzG
RgKec72OaXcph30X08FZa9hQPEXTXzzqEfJqbAlNER4pXv4EPk0jKXD/8oBexTHQ
PwYT2DcMy1p8t4NmdkJc1waOMLVntXJKdkm3mv4cTCOwBbOXRZHBLTsepKfhR9AG
LKTVaVxvzL4SDJ92QmHNSWv3eOPCq3W1kUtzTG4MvOsHnjUxHJCoqehGdZsK/lsM
dpwRxFw4Q6XbMbuzSU9/jrmo7MOx3DrCGewn+tynIR9Zcpto2NeJx5qgZ2K+h+kl
o+0E7YVtVej6blFKhSbv1snsI5lXhf7MPYoWNB1c9ntPRKpC07YpNV5x6bpUzzhK
QZhR2JHAWStQOUdHG1Tn9aXub7KrXtOjaQGVwLfRSLsy1wx597siI3bWardk0RUN
0M4fQtchK4+6xY2ghCxXSg5rCMn9qNSOHJJKOYp0ynquWwq3FQdSm7pUnHA+IRIz
yzztQUh+G9c49PrhXLPRLRYV9RfvS2/Mr8+7mWZWeqzayXrX6fOazAJO7kETo1fN
8nTULAS834Lk31Ji49jjz893vXsL8RRpOBk+zB1mqdI=
`protect END_PROTECTED
