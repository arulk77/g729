`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNznW2IdTUNeiJOW6feXJ8Y6SRL7Fl8G+BNX6KHb73T4W
rFEp+eT+nnRZqB7njLOZrLlTbPS+wyHPtfovfQTl4RS4dsVWuZLqvILEqqZsOlHn
sWiaFYpcvPKjwElmQn9c+ZoGSb7G54sGxjn7y4GUejrR0JFu3L2yQ9rUfRLRh4dK
C+wLL4DXyvj1AEqXdwynzweQzEn8rJdZA8s2YLClyv07PRQd2CSqlj/is+mKreob
0B9K+dLiBfFrGqjdfoF4SZaGu+8HEXkjdI5WmewZTFo59gwX1MeZWLwpgPyk8RS9
Me8R6pm1v2fJd5y31sVf6QBHJb3bBdW6WGYBU8USuEy8dDa5yluir3RYm317wONy
OotUgcilqF3TTT5VVG5SxPdFmhYemnbfSIO13WbX7l5T75NZBSbyvJLtpK8AWLMm
a83wwkLaQ9mbYW146NMJnnFlexuNc8iPpHpGmtM0TwB/N9tVRXr6jnNBZwpBwkak
d3IPe6B925RnRlRbqdCXx39c4D8xT1WrdgtCehfLJGDqg2U8tDv1Wybi7o6FXhVG
CIRVCCkNjwToj/K+ltUy3g8Ybb2CO6ZYu59TWBD5/sFQQuOwETclubmBDSLrmlFq
u+M2hgEQB/smy0YfMKNaycDUMY0c3FpQ+WQHC82j43Ei65N27pOcw+ASC2SqGPuA
ssJX1m8vWlV+nF6hC/QjX5oNhcH1xHUdnbHzgguGTA2ru8XucbYOGfCTyoAqh7p/
81/4dffBuX6cfRQahc/Du9xMMd++vzVzmEMA38jAXyOtqbFTCEmaVC+thYXd/gtm
iJynZIzsI2Vwf4Vh0dasdRMxZJMh3nTSb/a6wxWgVTINJOC9cRE3cEJMx9GlXVT0
eZKZkMgQDQxAN19j0as43I8AN8HyzF1B9v25FGMpd395gUy0zokcPKNWYr2y8f3H
b5T2g2iCD8olmDZUDqEOR6H5kPSO0XxW8P8yE3iGEg+03+kp+2cYVJ7bg9BDH1qf
ssby6eS5ASPfM45Y/GSfBg3XAyrKaIorZ8/qf2bwWgPBy/9cCYWfeda8IpQijUXU
TNu01/Y5FrxzMaN6yzUIg8EUbDb2UAAYe9RooKuHAPgSnvj6s8iJsaekxqtKe0ZY
4UEuegh98LtAUa8LSce+hcXx79MnhVov2GA6M8ZpZB6dDCFZxZuisPWxv5qDe1J/
QgGfDZ0YJwfjZcNHUCnyi7PMSoC3rlT6B8INuFxDGpNV5/VMTNJgNQlSaQLI9yMm
8a+KTwfsuUrlrhlt/rfQoV9tJxSrC1KM/Nc6RnKCqBXkc/yI63ApzPvRbeQHp4Dv
IH5SpKvL1IRSOZapA6c3Q+8GekJ+hvj4kGTNpiAIgogD0mfMQbvOKjzJcEHvrXRq
5IO6Gy2X8HqS+sELGgtB+kRr2mvEZhIckKvrNAhzkjD+Dc7hu1YR61gOHU73kc23
V9VH1oH3eXko3HRJGPQPmvrW6jRjKFb0rka0Xze39KCMs/pCGi2g6o3VDwqcxy76
59Ns+T0SbzhASLOxohpY7uo4uO/dZxgUqnOMNPDc6a0GcWUSn7qUPM4I39MZi5dg
ZCRXqaud8LOyDWhKUAgnFRQHdZq3byUYdVUQwW5JBABV2wmyM1A75TeY5KYqsala
/hRKhLUpD4yuGCJqWFPpB1lwHmmHhHD3cSWFv3snqfgWjd35myWi7NnUeXkkNa7U
Dab91VAxLdVdCZrX9lNZNG/gyi4At7k7jwos1JCMb1jdj/K3zxjOPXkDNbvgwo3/
y6oSAt1E7ZoanHRbS4dgemIMwrX2rf/lc9Dz9mbiryZlBAmSDKxWWLalyHPrKWdU
rxru/+/jbEAAEykgqdZa0OmbNjslj0C1V3qtHadsPLVc2kUeFske05DRRRruuy2L
VM87iNjVF1CB1CAsStaRshOdJQp60uIlsReYgmx2TO9LoKOOcRZ/vbGfjlgS3ocQ
842zRnt9SejYJqQDyS21NyQY/FAknLdbYuFj9cLwg+mw384EEd9sZQm701N1mMYO
OgVy4PQ35ALlbYtUYpfJRZ3DVw/54UArq9nz4Vpb1vk0YqJglFS5dTTAjGCi68BB
+dAI/XsrhWz3NuGwzjqh7Z7YySpIP8Fn2kQuvMXPL9drtyYtcvFhm+anu26CQr4j
idjshZ8rL5pjovoWDkfUQaw1jREdC+YxKdazh4S9zozYCUMdtqMDpwK2yFrQo6ZG
SlQJBfQFb+FxsWjlafuAZcUtDB4o1nN2g3BlWLGOURIjfwAVhtYV6xrtz1cc2ycv
BNji6eYB6Eo163nWZz3tjkTth0LLAKW/POGiLhuL848=
`protect END_PROTECTED
