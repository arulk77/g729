`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDD4nH5b7hwyq3prVo1x7CClcewfhHOcHp3bfh1qWwGW
Luot5WrzhUTGIpJFdhAo2d3aVcKt4+S/lsfdUuEuyTa//5JyioqvJAbJA30jh1le
YtAoK0Zn8aOpMxEJS7PlADlU619Zl6v90V+BEo/OFzetDKqtb2a+Un0kiHfRU3bt
CjxBx46BAeR1Or9ZbwL0Aazv6KCCVwSKZFXPTKBg3ljP7jvkqAnDq4qIWBSwlc4g
cyCBHcRKIzGtQl5osOwdsWA8t+pb1gnQNoRWj2SI9oKVq80PaukVuFDYIf4XhCcA
ciA/jFKI9fbRFPEPaH1iDQ==
`protect END_PROTECTED
