`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aymsKZ/R3EmObhbt8ihLwBJEcn9s9pYo0SNUgtId4r3ROSVCDKaxnmgJmebziQeV
0kI5CCbEtmDmIb/QychrFZkjzFGlzCSXGYODjJe+/HtRsOC1ddm3bDTlrOEOBu95
RBXo45NcgSC0bqkjFY/+bQ+3Q4JtJ0+iWTY0nLWnCIAJKSkzivtMTH+UiqGqyu7f
hFrptZmjzT+gHWtehIBa55PpDxypZpFoxH4hoqQZ+gSDUtyEgHAlcJxVQoQwW/Tz
euy2LrE/ww5hBGSN+xxsFtIHOjJotPjkeD5BIftepFwxrxwVeLDIvBAndNyOOfFH
Soo5vzhh22JHNaYadkanm9fUIKFMolPd6iMuTjtkWkek9/U+UeyD240m/rcySkOh
gwmHXe5aGsY8TAxdtqQJlZXI2QmHFONevCX0eoHxLo1/x3VEpDmpy3AaYJ10yN6F
thw54d1DYeq9GMeiMd5d/XfMb+m6/M0ziRW620JGHowygHtC66RUQzxH5C7E8kge
k3jLBUbKsVG8U3QyHbRSgw==
`protect END_PROTECTED
