`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SXCLWUrh/MW3ofSpa67PinJWiVrsNoDD9YurjMzef83r
YMU72hRv0UEUdQOn91T1bZHzxkBbSWAmhJi16734ei7CzlZBzy+ji1DuLxE9YsUM
rWIDkAQWMuu9L9GNnO+jk/5JERnRTcmd243J5yOHV8wHdIsm2x8OEO1BHBSpo6RS
5Q0QFzu5OzZQM2m6NpEnxNbeol2GQhC0TanPU/OVEJhWS63StEk3tEKrJ/cODHpq
rO86POmcw3ZAeKWKB0vlHq29B6ZeQXYyNDKH9c5LsYwwZ1V3/QwHzWgV25vy4pXc
Nwm40LDq/WRPSODIsrIAIy1Z9J9ozi+LE9vU/D646xKYfFZ/xnIMM2vME3H8NjPM
buHMdq1EOX0yXZFlZyRF/MbUHCr3PRElLEkIkiONa/nDPptaR8O4VV1aBcUeLmF/
qkuBfuOgW2B7xxptdrOYlwMSMlIYSirszZPMYJ+khCEn4q21M9r3z+hRho7j5cXJ
F3cZEuBaS3mor54nnkuENPBH2Rs/WijKq5oAmV+FaqgRd5AU/EYTFiaNyebs1isC
xW10OaTlkuu98lRs+p3FoDtIwvL9A7KVNFu7BGV4rv/sTBt/yy9LxFPgdc9hx8X/
w/Pw4+yQ6nj00/aB7AxAySiyv7TQ8kfbva+dlG1sn5MZH70SozRjI9mzPkPK9+jE
3pMwGIsk/UiQg2Yvhwc5wHOu1BIMvBwye0RlWXyobSCKXFKgtDkxl6iemDgSdIao
BBXnzG235r2AVLVMcDJe7U0ihMPOJCCECoZYHd+61IP6thcSIso0hdD1F5xENu+T
aQ+exUF9QPi1O+GR00olNEjoWQCyjyrhXxokIEdW6YpWIj45BlTVfQzLrK9vRO3J
JlOOufbsXevIkOFk35TnsQknkqKpcef3FVA60bSyyz53aoL8PYN/uYGwqhRdd7q7
eJJjvBhdCdB/mBcr3/PeeFuvmsHIhwSVHjnMnnM123mYwdgx0wXDkpRVgesU+nx1
gQ7SBHpP4Zt0y5aAV/4QEbCs5sw7rMHRDgSGa2j3Kq0Q5aWBZcKDPaGT0hYWXvrq
CYWSB3lOyZmErEGuJFIEq3BTLBQJAMPGU+JAZA/VwEbFmW3Fkgj6gLuJTwTKb5XK
l29CaiLOWZOwi8b5uUciRf7B1rwVXRYJHT/gTgAOPsv2pgwo3SMBRYnRNtp+L2rF
rSqNgTZx6E9nuzGa3xeOp1naAKpxyPRzt32mtcLqxRteKLJs8Q1ObjuaFZEcnCUP
wKrxw4t63uPvBUHaWCU4iALMwwvLR1QfTBQbY8T6ETL1CO4qquqKD7JvuxDURVDY
CPASUQPvYQ+Pej+vKK7iwp29nlGGyOcxFsaaozAScta9fWcoNwqaAq61XUR45eDL
eeH8ItYCCeH54JhjyOZ+DKPrDj4v1/cTT+UhClQJXG3oQW+td31K1lkCCnVHcmmt
LEfoXNUixcWtj9S8B8Zav1kW3DYOz2jN2bI7Wtc07F8YdErSEL22/mdtVZ8KedBw
THMhdakNKFTDIn01nfHbz6qT8o/Zm/mTxZyCAV8gCRWilUc7gg7wGtaBKrgAOshr
8pIjiv8Dv1gFxSL5Aw15xhtrD9w/GjmrDPZeazT4+dE4+GrqWBuTNRQ8fVg4crdf
Ygw2saWDObEdSQpLWwR1eT+XIagMaQBg2qq0t//96Sqt+F6U4xRfHwosSe04ll6H
/uxa+Dex5fiUAX8EUQnezNSBvvgglHiRNplu8i7kIHwAP8xIyKLS/VokVMA9clVI
qP00ePpKYSVc47CtgitIBbWL4fhd1VWmqg0npRESb3UhtZ2UVJcFK16SVYhe/xx4
h+p7wCr/FwLJVgXcRdUzqW8GtZwRhfIsvr4oNluYIxXF/AKN9B8Y5iADioNm39d0
2TI3I86vgWCQi1FxO2YipXAJnttgUn6/4p+5yiiUSGvBN9QBMeoft4mRNstzTthb
5me7k0MbS6tzV20xpr+uFSf9EVsA4yt27NHWzUWwCc8CPAqps15rKpMmAwd7HTEh
QHmOA6ujWMZ98eVef3OVCUnOuh4K2mLcaEYoUo8Wrz2KYZ8UjcVOE7r1zNTjeUcv
vtD4UwGD3AJQDuEeWBhnjVLEHM/gKpQ2VAArKVOu/++g4FbKvugml+6RQPk+ha8F
VO3slfGAVMUMUys+RzAcHWmKLPtm55rwxN8txrSyK3zErv16yvQfaWGDvnytjQ8+
jYxOHPykg+fnDHYPaJwCvNUyDrIDpwdxI7BuRh1GJXNzOkV3NhGEdnvKvTuJbRa1
+lbwLh3fN6ETlgqUu3B4fKYHl/pCxph77FAG1197uFQAjHDhXQpVCyu5vC+BgCe6
HIED8DIvmn+2LDAKbc6AEDzjiXxA3OD4qSAKtkqjXMJri3WK0ruBuyd9NUV9zdE6
qrZ1eS+/FYJuCN+3j60RT/y7Wxg6HKNtz7zyouzGieTb5Ex3DkKdO1rEYcw8R0qD
8K1kyafbFiEUP9ZFCKtbgZwv+TVy5dcOe6KDQA7o/SjjE6jHBTQz7AiL8tOrUtYc
NS3c/72iqkg5UJLKCh2ibIiiPl+Yl30NPm/jYuGBRwwHCEjK9RkmwbU7uRY+vdG9
+uWHExDhe4X3ElAE+aXlv+a6irb3Xmb7zmUOJL46+KABBxdS/MSmzdru4ytDVSfk
oREk4KhLfTjv5u3CEhc+9vQBl0Z3SzR3cGEXTJIKDTSoV5O9TKciOBlWr/7XDO7j
HX4wWcsyh9aaw6J49PtKxXvFgYZdlWB0AMXU3hfgEyeBWsLQ9V/jeXhIUGFhi3YM
2FoJRUzEIpXMabdHDixVKex3TViJWjXCwwuucO1J6lvNzeJbk/nPPjFbawnvGc1b
TctdESeV2MMZbRW9dmqbhKTz1q3htO9TLHO2x60n+rlHIQN4wFbE/zvwTQik9sAd
zI3Oet7RxHin0ccx6HpMxHsZriBcsxWUFyPDhAgChSPhXEGO1DrIfZcUu5uMtvvm
UHFR3oU3PPVQPU6B9nhLyx1N+rK8HsgJaoIA89Xb/ji0mieFwfKCv7WbZR9Maz4V
pq3l79dk1rvvtQYsX1NXg3jbvZYNDmPDm2x8pKM6dstD7ZPu//g7sdPYyjX0Qhl6
LdiDx+WjlQJmPjd6fLXCz1RYI06QN/3ZOU52IKiYCNNqkZU2QqYbIJxs783DQDsm
zTHevuqemv8RwybfwQqapgRvSIcmvyC+VPiImycDCbAgecwFyHt+VQsjAsoJlON+
WGqDqOZeoXRRxzbmXZ3TZMXLV9TQ/KSb2aiecko82YYunfP7eHjHeSQg8cyCVZGk
bLS9dfEEW+P52w0+aLjG+5eKhiI8ntRPlnH+UazNA4CKfqxecf3bo+WW68dQ8jCG
9Nx4phpantp+hI0gvF1D9QeWw3pI0x3Qqw79ajNbyRIg/YnEn+WHFsKaVE/cygJ+
YOiJpxZTMuLYf32+H23OSEn/7V14GWk/CBknw9//Wg3vTUkWGpRTKOowIK7RPZIx
vY74U7JqKnv9mhHTTDQvx6Bp04+P7hCH+sg8vdkXpQTNR17zP7jEgcE+dZypXY5t
zLfUj/LHeYF6Y2Z1oqtnZXgWCAYiH+334yamov9ccJ4MMUSGgXGlf8wAxt4FwaC6
tUwyZhtVKJwO3n9mXB4twwC9Rd7c93gaWcdFG0aVMHKdlpaKOcsAWxAdh8gHOqV/
V4GdliKCY1GHBbEHoG0ME5MjyzvEm8Iu+mKpTtJAWcHpxjS4Vn66msoqZT0eRQt/
pxR1p2FYXR8/LuqGfzr20evEGRYwUoSVU8D96EiIdiHZu1BNA07STkyvong5gP1+
7Jdy1pr+hPH2VgbmfTvPlCTq+pvm8NBnn+vNCkJIJE0dxqsol75au21cOTM9qmWT
XhIAJza7z6UxpZ0kJ58KM6Lp6urS5VJOU6o4LbdE+2dTlTI+pS1H0yjLrraxSRsB
Po/sy6CFHseMukoe0pXj7cwxbK4tapiCd9woY2reR0QkhGDF9iAm7GFLNB9hmwR+
Ua8VSX+h1nbOnqp605cPRxwDw8llV/1DSQ+WW6ZVfWjT+xRsyhtycFqC62JgRA95
I0yj5zLHcTlsJw5dqLisTm+fx+WMwP9j2kcQc4ogG4T7OBqXHr58maxl90aerikt
C/BwwOhOJgBXjN1fSueRnUYAA0WibxM6lfWh2KLEXLun0w5TZ/2M0/Ry0XSJ5dAZ
wp6mRcwqHDHKstqbOc9hkZqzpKNcHvRdfL3nADfXA5UQQmkz+UlSja+YMX/WGe2T
iiAKV1B4EI0lqEQ29JQH74UvTK/KkWj4lGVvFAmesPbWZK6yDsuUc5r8vtUQLpH3
Scj20P+kGzBYa/RJE4WA4iJGHqYcXnwF5kaX4c/YFbiiU/wENB+bq+4hg0keR/jV
JJJdzW5jnfgl4FBQkCL9tLVS2sJO0JouT/on0X1JOOQxdkXn7e8Fiko37i46sckk
MJwm2kte9KqMrOgVU58tatCl+fTu84pWvoQCg3Myre3JJrnTSGdhmCAHNMCLg1HV
tvAhkQeKdtBUIRVp/GbYS7VUME/6VtWNUSMHZeiU2bGZ9B1Dv32Cl8M01tNed18w
ECIhkSlW6o/7TYqYllaVrzUiQIU2LuoMcY4G9uVahU61EFTEe8QwCwRxDF1S0aBB
OFdQ5dqt5ZE3xGJy/gI8OHYTbSGTzlTMsG/zaWFdxmEtM5n2CnbAu0UFf7s88V1d
yFDGYnFxFtIVjvCuFW0oli0r+5z90OOSOh9hsCbDmilU6UtbkbqhWm1Ki5cvLCjW
xNw88qeShiog1ubSmAMQPYMD27De6qJEZN+Tciyqw3YDun7rKF2W1sI2pzgk+hu8
Le21diLK7g7DzWKTzwp7nYdpXSK1eZOrkMsABGJpd8CJyU5WVxXtuY7JA3jJy0Jf
naFPi1Xp+OEMr1dSS9hni6LXMWViqBP3aAp6fq22rzfrdKf4aE8lDdCKbvWC0Trw
LyrFRT/ZLYEW2jrlW0meuQYr2LTogNg1Yf7xogCogkSLVQBzfeLvwDDR93tKDB9w
e0GzuP/EfaWt7LLR9SypaTA4HpxCc9tyR3fFxXELocHnWzC1INdUNCP+QO54XvAN
kOCfexJUEQydBXMPU6BcfjLdLpgwCZ3vXzO5Zjy4bmwDEGCkhIMe0aj6SsIopAhm
6N5THWUp0n0JjDBSnrORPYzDQjDMME/YAe6ZmRfCIM8=
`protect END_PROTECTED
