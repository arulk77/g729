`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveO0pozzQiQAH8dabr9sAoQVQCGtWvxPkc7QZScLlu0Qk
wJEOPJapMI2iP4t4csMVk8obA+vhcbhVZYIz65/smWB3ihNwJb5QmQRLI6fgySSJ
Aw+dxalcQ+sXsyMeIadm/69EQYSNsT3ApTNr1el1VzNeQnkQGtGjydBl72C0GIme
PPyLN04D8XXWRETe6Usk4KYnF6mA9V3X95O57yW+a5j27jZBx7p5A+fx3b31baN8
Lm9INJicnMWMYeT+IR6nKBCIScJNKY14lA61kT8r7U3k/itnrKZQrQnWiQ94fWVg
NFUCwq0RMzbbmJ1BTNxSWhTa8/1t2vRP1eancOG1t4nqv/qLHJADHWV8U6WxXtAp
IzsQI6tYK2nWI62qHiMpr8iQ1YzvSah+xjOnAVFKnBPQTO3lK2ad7+DL7FAcH2pg
`protect END_PROTECTED
