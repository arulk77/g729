`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
OlssDlFlz19Cd9IgZ5CaF3NmQjO66yODin2jc+tr+YN2sbPJJrypLQRH3FdqGkic
Ywx+P2kH2BPLDFoG4jC4SFBOHwgJBUEBjPDLLLdOEGFE/KTb+dUQ9Ix3dPl+NpnH
AbPzP2lQ2gxeew25+J2kTH1NJeZnlD/W3cED1OqEts1Rzy9csav++xlGptaTbJyw
/qplv0YAJnowoiNDFw4vfLp3eWxy5h+57Q/NLEp0OSQ=
`protect END_PROTECTED
