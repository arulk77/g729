`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SSCfJc2mHwCmlv195dBzeRrMGnmzo7Y3N2hqnVbVPH6t
zc/yVkJCw64dl/C7GEpvjBJPA+v+Grrc0Lvkc+xUDcMpx1qrJ3Bps6Qu3EPLW80X
z9mB6UY2bYocfhYKot3RIOGp1Nv0IqnaPe6rducQcvp43jvoG+gxTx3b6oDpEljT
KGX58EjV2n0HdB115+iCIPfynGa+6RajxD54qa4JePPrOp6OSTExg+6zvRq0va6Y
SAfv1x1wRsT3po3uuiG51ICZTzsqQmus/38Qhk1HacymugI9XjEYFEbMd1NENmzW
aVQP8h8+pCictM7m5lreuHwFN/VZRsRKa0ngIyR6PZ7ckP+PasZsdpE8owr5DkkD
DmQ7J5K1RdhjQ9irYOsOjqHM1kFIZKoQvvup8W7hDZ2dw+FSeaaW50Vx9luimNCs
VhhUwDE5r46XdmRVZlNkBRUlTUDUxtB9xNMZSENkOxYSNM2Po8mi4JqSAUOoFeQC
mL+k2BsT7Ns/ki+aX7kTefpSFCKjZfTxbl1XFXxCS4JQi+XFdonuMsrhU05/FRB0
ROeKXk/8rMFK/+8f5YdmVhzE7ArWokjuPMxBIK334pqZh67ZnlokJAc5wm20+0j6
5QzN7y7jtFk8AWhZCzT4KufnxTa/a6m481z8YQDG37Lm7qXT98oenRX8CgDKlN6R
OCQ/P9jshpiehYF//zB0VKcieHCk5I9N7QKACQwzRxa03u0TTBlAmIhtrDDUiFTi
sb0E6JE4yuo6i20ihHndwPg9eUeo/plGvbTLVHLCC4KPzk/KN1aV0SF4tIgFttsy
OZurhPHnUXzoZbgBIjE6lnmdoPFnAvXQ+pqdsrYVc1LAXOZBoDbXUVuw87sePZC5
FIuxBgN6Fa1nIm9qzPbdaunVtewM5RcZp31e9TxEhRpckXO26p9Z7QBojhfyBiha
zFrtBxTZONs9iLLPZq0mi7IdayiMvd5D7lIlZMggqlpuUNzo0NzH7B1xF3T4BadA
bbXzE6so5xkX/pl9cAgs/zKrO5AK7Vd2us5+ELUC6A803W/idj7ZjtJqw6GvdKO0
YQhoVGZ3hequlU+fmCdcPwdVVd3J5G0eaQGOMqnSZga1WvWHkcK3+sfIo17IxaEV
Wbw3w92PvnaaV3j5oKnKGYcA2FUqy3Ijx1XUZarpF94CjTEFFIIWg07BYdMxkvGM
J9D5JPQSJmdRIPPzQ2vwGgglUc/9jooBpTqkWeW/KDibn4Cw3PMdZ1aZePdLTSqk
m+qniQeWLK6IUIkLaseRvK2EsuvHYqgtdd+XnTR1A4gyYQcrMUOLlpRwB6+AY2Ej
O9fmMInMHcKxhkgVHU3cIkLApHHIVuco8Z1b2tiSimM4/mZqTVglFmk96tI3R1hU
wrKUTBWb5RGmWRUJnYUiX4hyY1CJgPCS5M/QphX4yJRL3aOaYh8ikFsXpeZwpUxV
CHbsa1uv38qYhzmtUOOAXr61ohxpRYZ1tYsPLV6/swkh7k63TSktN2B3q4SdW/6y
Z/7Bia+jMc2sq2zIJJQnZfRIXcqvV0dDE4P2+Dq8+czJWY86eoEOyksVsXY9cCga
1VNRin9ujIrE9XSqRSLzXdqceTiSgATnXAutCd/97MqbuxUfoW54PcZ/1eKxpHS0
/CkKf2SncxrhFTwk71ROz0hMkSmA7fWRULr8uH+hh1pL1RfiTx2ZlG4iNUr4NtWb
RRsVwhwUjohPc5tz3FW9/rfTbZH757pqtB9xp+4bClWKI85UUWy6ZY+DPU9M93TJ
6bir5KJD15bgrL7HHX0wvLsVYybTcsUv/5jJtA8fD3eJ77W3qJTSjXf3LBrEoEHg
jbWzfog9q0H7fdmn3FUDdzrdggRxJENkUyMA3PjpauM57UIegxLdprnD3QWooKlP
Oy+9npU9uFYzAL0plXT5bR+aOLJHdKZGmpBvmlCAg3Ad/1fmcngLoSS8orGjZTEj
CQHaFKW4Vydpd3LCwyoGyBrs3TM36NKlCdE/Uxev8FHrNJOba4xKYrGH/kSHfYr1
dTwIpMfMhfhVrhks+/QGmqZQzg3guWcmD25FGtQqwIZSqxdgLi1kKHP2x21yeKv/
PLM+WWzAbXUNOQlQaxkRRxYNKi8aJHhTrpDv97Uz23IZXwcWFFTBgsiGG3zd8jep
mTm1j4ZXvqNUI4TOcy9U4BtDhcwBZ5Lr4rO7h3jThSXYXZn6SWvhpwRuW5IX48Fa
hJydPQ57hfhuUYVbAPvGe0hcNCSa1ajtSH+0bHO+daOX58bsJRqnOOpAoVHRTyX4
45aRQjBQSOI9/dKkBIZJ7B/B6WAjpFoOcagctNrWgIf1qxl0SewZj5xxA9l+HIHF
Oyf5AuAyNwQVw+l8pgy3FgToPYjCRnaLrUEmlsyqWYMelCY29LFXPsKULaX3ZaAA
ovcQmlTZAPsoxmrn2HbM1FzoyAy5FQFMf4e9REl2S5edl4WoO0ZJAyqkXjO8U0TA
vFZ3LPygATmjOeoePPXg5Ob0G0EKAfST2Imxif6xpTCWOUmGvbhCMLBMtc/b+vRN
PJVDKYh7yOWIwV0kjHBDWmNFNtU8sdT7YjzgQotaIDG13d1+JdwAted2wNzATF+1
bepdccTbf++D/w1AObMvoxR3vk1hocLQtjA31WpOhzZyAB9vJq2xZ9dho3fMPe8v
MQL2PQt0Uo6aNnERRg+Gl22Ti5VDrK2whTm1aQ/7JSprMv+Upp9hvzTMgHC0Cb2X
meb5svES1qNpMF4r1juwiprZBSrsJYFjmqpcTKiTrciY+ytYPY+xBTbWPURWsqAf
cxuqdCH+eb1TRkTDDmIFx+57BHHvZX15iKr/yHz3e0MaXaO++xTwWTMjVODDkRXn
yn9UU5yBAVheboC4JWqMG/j4DT1CeQMPNPOwBBp+W/blO6/mTjP0502Z2MN614ZO
iAYcR3BWb68RLXrwAD/dv00AFUy3u7ID5YfARbhPs2RNWx3PuJnQvPRC+7c4bPxV
wQMR62r6doSDqIJ0f5/h6bEfQtWGQKqTCbhl35+2DuLK1mdTGhqPbn6/u7iiScNh
dcQazMrfI7SfRSmRJxLx+juBrnAa3cvGtlH3wyijA+EBbxN057/Wyk7kvAvjwiXx
6nP3lZTqSNotrHqOtx6K9C+k9c/PBWw1h38ykA8PdT/DXB+1cg89+I/LytYpnl3P
2CwMnHXOL6fjKhCraGwcrRN9MPL5itZXFfyRKUCeEiE6WNUqFXSGu33Br60hTaWd
IZjrVfHzhxlV+qxmPoBHneFFhMV5RWn6rzThpytoS6WWOVWLr1/GlStRTutgQfOm
3AtJwm16yLVffkgj5KEaOHIZGkJbCuZwGdXb7uSSDPVYJVZ1fXOkJbZKu/0V4tQg
H9fy26Efx93iY2Ep+p3/lkmhVf2FuFXNSt2LSmErcpNukNHCs30hUCO68ssTMPVl
qxE4pcJwRUlxkUPpB7Yr80UBA7RVq9H4vmkSiLmzTPgMj9MK81AWAnVFuD7irm0r
VC1FUt3DJS3nvtJUJN8xVi2ekpD9ke4fZu07UTaHg8WPcghsgm6JYouqOEbJbTXO
3gJhSx62/FFTN9Blq1SxtteboXiJULqDLgOidPYrD3Dro3TqVnbcrSEroeKliLay
Re6k8c15CY7vtn4r4cNhZjrKlBlfbbE6Tc8jJN9T09/Lj+He5IqRNDwhrhNddMCJ
zM2eCDNwy5Hw7AWp9IFqMgLHMbW7VdKbJhu8EmTPpD/3nhKr6lkf8mdXJ5eLwdnU
6TP2lUph5HaaCwejthMMmhrUYF1vGKcU+XkDDuO59VuQXylFUmpt1kxdkRtnBpvj
6PrdLIHObsRpu7tPHjFcIVZkLpAWRTiw5tR3mYtd97WqKhBIeeJTYejcr40WIyBQ
s3FV9hSew9b7MHugU0yHQ7LSuLefDKypwj+4N90m+WFz2ljGYPD0/DGdWUUjvyVY
D4TBR+TxhyqPFGD/eWGApWpF7HEBPWjS6Zb7Y86l6Luh9md0xgK5qmDvkDyFWXBR
5uv5lPa6ATNtGUuVF/gEWLm6OgGdLmOurLSc45+Y00tZ8IT10mIm/gV8iotbGawF
6vIRMgAGQtmOfN6Jh0SBUgqX73L5kgMsxZbO8kMtZQCFJIWyd6StBCNv8aZ3EVun
bas+AYVzm9P2a//P63rSpmOYR5dgEAJiUJOoWZUPytRACzt85M8Fw2ZmMjyhnI7f
srxIHFbe0gfuF5fNaaoLkgvw35luJ/y2yaDpI5nGaQicZTWjE/V1E4ns1pv5pg7U
kIXNYVGcOnDYiFN6uXj3ec+LyAXRDlzONTRq4jBXWcDdWaadePXlh48eLxG62ndQ
jGLnYGPnX94V7mUZOvoclr0804OL0JeDB1ZCbQxlpJR2F9cywvTz1CzzEoSZMALG
h1/vLMXpDZvEzor2YPTMAkjLttnOSpBeYVOSdhRWSDr1hW4EIHdVSvhiy4lJsAjg
3AMIOPn9Lj9562P5gslarjAwEYPCfAPg5KMHCaAQ+I3vZKMlGfTxf9nVTrtt7Cgf
EuvVluf2hl9lX/hv1UrH6oQCFf0YSIOiQACyr/ttCewjN0+40YuLfBWpat93DnKk
dCgbfumEsoDRVWSpVJ3QDLZp8PBWNhR3+Q5zx7+oeQpQa3HYqEFHRfw6CLujkfKr
58IdXNwxbggmf1ADq6EtsUBXDqNDosJDbBKF6xA3LRtxz2jvqRh2JM95lVWZflbr
nW7aeUIvAxikxmU7DZW7eA13lMJdPsO/T/J011yf3TC/+2F2HqQL4KVVx6xiEzZW
3Rj2EuyFrr6+gOcHO0HNUFFyRzy8Myo6NNnEZJILXtEGexvIkV0/IRbUGsDHArBS
BJryqjUQrOaa80WTCoKCKU+AQ3YVEQ81yG17sdWJ+UwyaKkkiqmAPo/MEOVyveIC
DAkfkYW85y/3f6CaJXLzZSOJ/RY5mUaA67xsfK5AWEyb/DQvsolBYGdEupMO8ert
BRQj0zPHqLSZdzxCoZvF1K3N4C/euHtVmfexDR+3rpsMtp6jklDq6jPkJQL8YGsK
Njo1xEEty28UIibd+etvjapZEy0C+uCqKrumjxVGsMx7CQ35baTCPJFNyx+tbzNU
OtNRO8t6wBcFhD4ZHI7tGkGUoRd30MbiSEP6Ae1xkx3qUytzQJRU/p6S+mzEHy9v
ppJOQ2eXi2aFhdspokBPxTNIIO06VPhmvHgCFS8o37wm/15E2u2Y6m4rCG6wLKL5
6AmzbDilXcikaSJsCRh+kav2ddsKNPqV1eUbrgyYqJyPxCVzwkLM2fe4ZUMLZkE5
7cVlvoZGXTuhl21GwfrzsfPJ9y62JzY1RtqOln4K47zfm0O+wJLOhr3kW4jX6Df3
70hmyaG4j9y3NzRkoV9ZVDr3tZdh0eEndguNJuJyS3+EGbaW/hfcWHmWDB16puVv
nt56aQj5fzuM6kYDS1hnuueWFhzGRn/v3j1D2pgAFXWP+vRBvv5Oa8lxeF9TRJBf
4CmddkaV3Gf9Mj1nPl35HjNVXbLI/aXQ6LGIyC/mPmMnVhxtp9zDnIXaegjTwTnj
URDDhr0dxexmzS1LlvyoBkmq99mdQR73tJ5mK0cAetf1lf+z71psF2HJdNPSK58a
3SG+NuMSZ//rE0D+Tgtp985qTMG9yt+xxOM1tO0eOY3bler4EtxQmW0eyL4spTcH
C3yQ7cp1C9NyX1akdVro3RZobtz7yBnUc4HmMt1sLiAZtFa8hr9NStGRwjyQAzki
xxodOI3jm0Lgq3ndpSVhfBOUt++bueqP/CrCm9C+gkikyMx73DE/mvy3sXbYugXK
BUVsVJjGiMPUOF8E3iMlAHsub8J85o9zu352D7yAQsm5gbRkru/fd0mHzVM3wtUO
1YKhk7Xo1K8hoyCmC3JIPxo5I7pTUR3ORq0RstJHsdpkoed3/W+GU7+ppyXSlIZU
TcCpKf/IqBRZyiH1ilYVrKzeCJWbSvyXa+uDyvNpA6XIH56t2Unmciu3NRsRNjrc
Pq6zeD/ZJo+//q0QX5E3bPOFjgTSuDsKKkt0RBeNpXUwUzu9MGV2bkDAxc/FNfWm
sgNEpqQprBy9XJ5Bt7zKaOjx3tOsq+Y9xtbKLW4hQMNVESordD7tpc7ULWQ2y5wc
5jkV1FtxT0r7+DCc9A7RR5tXpMlXC2NeFW7XlClY2JrDolnjclzd2IVxHjz/dQYD
sgT8Fsy8LJYefLTiEkIZD3JhAHnDGZIeoPZf3WetsdDhq1cvZggTtuiT9Ruams8G
e7MsKw5/2P32NQNBTPKURN58I1s/yc8pE3A2l6hodnY56QGBBHZRUQvjKNA/KU3l
ZNxnUNY3x1wO5OXjBQeE5P60t/+EdAPXISBuR7du27K9DYUeuXGsv6unVQP6v50f
JlezFGSqcUF4VIB4BtX96TkBGzDLpNIen4AEZG0Y8U236iK2RVJ6xXy98xxzL9IJ
K9eGX7QRU+cF0rUSL76Sq7+mRkjiC8cuTblpV2YCg9cXChxwuKH/fwZTXzew+vHi
NjZsqEhmr5hK0nlbnmQjnVjoAH7v7BKJHWwGHWyY5qF1N8es0b/4+pN6/KvQ+pek
ofrs/75zmwLfRTywCx6lXkE4Vop2hfzg9GYmPBOSA2nMprxQoRG35tV3P3D0q+86
b5OYKnQCIVdG0CDZFBWlcPjOov0XiqdGc19eQ4vtb1oymwqQIb8Ugp706OQHiKM7
6h3dVcXICvK4z8VTAv/rk43u6sCwIoGpB2OBEdbURYFay4gz/g943XTcIoYpVXhQ
X8VB937AsnhnaTq7WSidJNVth7jEDTj0cevZjKIYfgZ1MtdjItCO+ZPVunfJURcU
hiFUn7oy5mUJ0zKrFf/S64jNtaSxvF4O4sbWgiPAY5Y6EmwLEhatnlG34Sb5cyND
HMYoOmlo7S0YdoOM7AKmYa/srwEAm8TOjrc1SS18CcledrQVug4kXi2NxgLrnJ/F
Ap0R27hSEaCX7zZfRpQPPQfzDhr4ZGvJYAA+P9lbmPd+bsmn2aS8Qs2PoClTLdsy
PJnCdd8oLT6ulvmjSMllOkwqDrMuZeZEcB3WJjxcDHbOsH1MnmYhyiXbqAab4yJV
X071M7p2hZMzzsHFrvAoZLUqrFM0RS+hi4M0UafYeTFvHZhR8puZzKAqj09JvH7z
I48LHSYpFzOUrwWT2IwmAjsH0UyC5TmvufGC/ryR8pKHNiRWR3luRBjMtBwOs6KU
R80Im3T+2NrJe9OamMPTTc9FFvAS6VcAtzz8H+JTC7v4z48CEaEYzq+V0h2NOhtN
rsBvC17Zq+tRUW/h6X8KZw3xKfucjkU25pVx5zYfS66o2UGAhRK1wzBxH6RieXU+
vmOf+as9PeoSKoKG6q4HrGxP/fU61bXZctXo8DIBnBSWVzhLWPLeKqInd3K2492T
Dj4U9luVWPwXv07f5APil4NXPuJ1jea5bfnMWqIH1y9xmREKe48EtUdsR9q5dajS
xnVAvTP8wMPDRcgats9pibtmr1HlS6Un7yW5tva3u7Nhcz0uov3HdMZof17XaKUC
2K84EafkgafCeg+IVashiokbhgvbxki1wldsJE/XxRYDIWs872bmQ0zfawB2n+U2
KlHjASr3xaqGqTe9DUfKrdSDfLDm7QavacMSlUdpPWksfYagcR3uPTwqxJ1w10rS
jEXvrhV0ExBLE42cc1t6dW9ijRHiEP20AtJ3IcppXgQX8+J5eoWl7SZNwMQ1wtLH
E6UE3odbLK7B82nauTXCle29ognUezd2e+T+RsgkiaWKs6UYHLXSUQgx8opp8Ldx
Bg1Sg1lJLFS9M91gAW7Klu3LI/XqBjptUS8MTjnBPyebiczaUB8igimKu06vw2Iy
MSkuNA67+ATdbrE65ylSuwz3PLZwc3rGVVubbgMqkjNMLuXbEvDQxJ9da2pDKQ2Y
/xSCh1vRH9OjkKYUh26LcSfIkG3QdXFt22OI/ZQxZkY0HCevtETEr1Gx6OCS2Ua2
4gBvt1DQqjmWVl5FY+eb8meDy802BQQRH5nqi6Ziz6+qr4it5yRJabhsCjAKyFtI
9zmIVWUUy6UVDPW0oK1gMyCy1V6/U+UdYfdMULtaccNGdaSQqJDmvGlb5gtPIwTO
D32WrZfyuu+7WeHJ1rnuGZwbRv4GX/NzfRLKJ7d01qmJrkDz2CPUgSAC/gvWlmjy
hzfLr/JAujvkUdU6NsXM5Gjs6qLwif+IPmVUrIiFDAiVA7nH1ih/Ig6bViwZlAMo
aHoxoPpnMJWLx+BJ9b7luF08kApBLsDOe/ZRN+eBPoZIB//Jd3arRJ9tyS4HF6LR
KbVek27vTbBJhIR8uq71ssoxmSso+vCaQx1JLiG0/Gg1iQcm4OO5kr3CtI6GLpvt
F2I9wPL3sFXGx6ylYF8NscJFH8ZWIodJi60ljF5NGFt9Vv+NHRHRCkiUJ8VBgrbc
T16gzkGX9I0CYYySKY9QBV0Cv55LSgMysaf7UYOpQT2mXXxgDaVaPQFkPk5Ud0hH
FDW+ANFwundJ3fG+uwSX1/5oIQi59KQo4ovWYi0CQ2h3HgnYaQCEm764RvmhhL1I
C6gy5LiMvDqCunVAN7kxYFcw5uIs0YxZp83NsPAsxf+n5kCmo8fiauFF0MWYk1Bx
T24JzuZ5UBtzW5ovp6FI8lM8yTay6ePrs/1fSqzPLnNWIdeU1v/7ugESJUrTTaHn
EkZEpzbCucdC7GdKeRjHbahyk83kQ3x4kIdq72/C1wBE2PGqTwrDjz9TYxKytIKd
hXwzASpK03M8h8STgI5xOI8RmLDwlcPte69VJO934qPGzZcaXULr1UEitF0ME0D6
Ba0DWWZHjS8tGtr8Cu0/IPDsozDc4R2N+xDV6W+nbNqk4oP8qZ6sz44EtV9e+An9
oL7+kRnYQ/RN+pt68HeOFh6uj+OTx8zXl3UFTZzTDGscMd6QDQLvWCazjeWj4qco
LolFepd1akETGDF8kEKRG9ZmY7UbnJPIYqyyckT2JC2P54J/jbk9ZoOQiay23ktS
+uqh9bIcVRekI8DCEZ1ZAmuyIH2knnalQiALbxZLjOlVr+fS3Lm4V1vEnu0BqH1k
C/T4EEuAnK73asYJ8pL3nl59GyBSzgdBb2bLOT243FJnnDuB/jOct1wad2nvfTlg
uWtVbd1OE6YF2cf+XmgrQCj+whJwjw8Fvys+crbcFyxn34gd580WdRouPmL7F028
G+qa7EP45+usoY9qRK5U3LtnFi7Gfk9Ch0zVESARjccUphC/T/NwfeA0U2UUBQML
kB8sMvZitLSWDo1Jj/RpQuHojnM8A/gV4a1VzDFwf8vyzfa3Ruasp+vfO3ORZYmN
8+WQdHQ/cPSqzNSaWbaMBH3CxQlv91kSZb8bJouagPI++Kw6aN2jD/zPz2XxbVjc
Ec143y2jfMFUQs7kSjhFJ8I9q7VrLsN1AvA74ns67lOze6D2rSretybkHGN8FVR0
WZXVmPU1h/VBSPoaiFndwhUl1WY9QDezLGm/prTuVaONNV+b1pTrfOmfc1krGwYV
9wN5D1H6ulfxdx77JegxXLDYpHWDtm//6s5AvkFb09VAmnYriSVIiRKWYd9f6MI2
ak6jDzK1N5mmeYK1ZriCW6uO7kiuK0YevY7r7FufK1zmRw3ARsErYDhBOaXDyvUB
TMvaPF018l+s+YoY/SY+KOlpf80WdUNrJ7QVeeEsyYD0zfOKZdPqu6VE5vXrH8ps
r3BPJVmMxku0XJgL9zZshXtEoZxXMFBUMTskgeY0zScsJThsFIz13AJn6B+yfupU
BHBR6X/vN5/g48pRYj7i1AWzXs8mEwFoFgh0sly+JmueK8kSaUnqO4c4W7CQMXM9
Atn9ozG4wO44MP/xHgV/uV48iP546zlBUvyFTri/sUt9PgGebrOkjy4gmlD5K1S3
5GAP2i8GB+S/PYT69CUEnw+LCaN8dwSfvhS80wbIXGG1GWFEXhbGPr2/0G2QnG93
54XZdr67pWzBu4RclkaoGTAru8BksKP1v6bh0sY7s3UeyBeBUrjlc0jYxL8t/8mg
QwQvW/NmJreZJYbPMyQy5DjMbaQYj42bNlgW9KdV7Fm4IW7wkydY5lK9hfnPNUi5
KIEGYBe3tzbVvBzTi34Wf9DHoJViOTwHV4TyuNiAIFiWzaCR7Ue8tciCV5l2SDp4
v0BZ5nQDzozDoeTlmPwAdu0z5Rd0jPOD32n/IhIT8UBSZuih8W9mQ0qJdkEfqqC7
h3ZzxuNRuwBWgkPguK6PddcuWHiy223YJxG3VqrgirAMlJxN2ZH9bxH3xTaFa9kK
Z5G8lQuRX6bXAA0BQTObuKgcPQ8o7lnM3rum2+uchHQKB5feHGF/sxUgfmw5LFv9
ifG+WMq5uyLwVGrJd/1l/yIbt+nEzmz76q2xhc2HD4A6otVUcoQ97dWAioieVclq
Fr6pitEF0PA+oYpG7PnPdplB7WZhIZxFLe4XUeGeaF/UizCst5asWs3JZQf9IkjG
t6hMYU6lfaTSF5AnfwJtXNzNo4lPYIXGNpPDtu/imCYl/nzGNMg/QN1GMdrSfyMk
dq5jE0lYQQ6i0QK9x55QcyyoSOrQwUKpUlC3+1H/pcX63XHZBxwRbzmd3gVpXYxe
fyMRyg2auWHjoVbYYDBXH1Z4PwzCy4zDtWeM5cHs8UGgwDph/Q++dnpaYWhZQIGM
qEtEqR3SVTxCMWYRNI6oUT7UPd7HqqYDUey0YAvns1+X9JRaWj/o1gNx5yB9T7QT
T5T7ODUhf4b+he/bqC7G6IJHs9TuoIfPugNF3VmdJK11tPsyIXKb6496RDgEH2AL
iBa/uKQKYoPKIZXj7qRhabc4deuIMaZ2oMNQkKCggWkikxJY/B0hmpjMJ7F9lmqV
dLUMkVSsrEpiweeFNqMQ53MT6c7eQ1vJC3vHmmG340afpopGnKmTJqHshN6lLfgy
KESI+WZaLIPu6GakK1TasfBTcwm63Hs//PoipZsyZm61Vk1jyzLIQJ/xDVWyAI2z
WPx113TC2uRRo1+5jb2eJu8AzGWB/PnzNkzpsyvyFiXl6YqyJPmZggZJMllXkBtx
CVmogVc0dyYKZMP4UOM1GQp7ZHaYnAEEWwOAVGqRuWxv8ZYyZRcJurSNtF+WmnCK
W+KG6ttc2x3R0rlQV/f6/FyKxqZ7pthahSQrrTiAjHTQSn/dGWRVqIHqTupgR9TD
2ZLhRFc2lfLcHBJVE+8Xe/qD9U9/01DvDnzf9COjRM/8gUOhOO9ypM4RB4K1Tbnl
SALf5vJ1v9FpcO42Z2jhxS7llIvAeAyjNLWNEXFRYcB60zBtbF4pcAKO+0rmDZGb
iS+r2bWDhBdiitZft/KM7ZdT37faBnCX+gGIhNEdhtG+AHzyK81LXZ5eht348mp1
qOGttRBMos2ydih7qkEJbG949o34JnxxA2aJOcHlMX+z4007IuxuW9xjeHoX1Gtw
/pzWSUI7dxEPbU31xvPR3xgjbU3Pt+ifrTcq/og7Eza2JKZNvasIteTOTbZLGagL
Gd8csDXpAwtu+opNb718bzv3szpRHDvFII74O0aNWKddteJt3QRa8scW6ZCfoARw
wy9CL7EjNZmf0Tcw9cknO8Olez9dr8muyFwi0XEBtp1QmS97LKNwNXKtIEcTTkQQ
q/JY2KUpHhFrlIK2KPDdBttFb/eh79YrSsQ3VtlrXigi0IuQnRuFFHtSgKwK6n6/
Qu/vvUQwAZ/aWjG2ObGWE71MeA7EDvO9Sr5iw5iCjh+e+Qnvp1aEYOuci+9g9Znk
IiaWsq3A5ZQYHUi1+Z7lQPgT6bvPN84jYWDw3SNwv1Y1XGgEAcsTZ1kxT3M1AX3m
EwDCuH4c4nYf8dbZTV4Vs/NMDtYUx7TBTOSAAvktdVft7j+LadElWIo0qWiU0uFy
R6D3ra4T+XlLzSThL4MYJhTSoVc7Vroq5BT4DlJCaf8W8EtU8I0L/1MJLW8RNijB
5dlvWk2YBS3UWh04uNIMTZv97CToRr6vgFgK6D98PuEb0cJmv/VY5BQ3wtGFCzWA
Ct1n+evRd1lbmlU5yiQO7H/ML6d6WBl9wmly+nEGYwriegQq7SPP6A6tlkJppGDl
1eGWQVy+it8fiTI6aBAHM5ZnevVWDIW4ZX7DRLEVO5tlJkJdGwN7+GQfSOBbvjOW
OH13dXAjGA7eTnnudfwX9mF0b5QVpIuXLhNJ68rTGrrm+lY7azBbOZ82/td8f0B3
B0J5C41FiKEbDkgdOkhbnqs37cWgfbr2HBNKOWVXq8bGyMJPSzF17h3WAb0Sf1V/
z96PwbFohU/UdOLtnrxkgv1Arn7CdmHRZ2hcfPIqKNxcbgoThv7vFkfbU2xp3xGZ
UpVsc3LfR8DfBjNPgGlnxRu9LhqqNm+8tfUUSC4F0ruCysRjDyXCUmmyp/FuKHo8
vd1bUTxLWQ9NX9ovkVbmt0K4jAZ2fDzml8fgZgsRHuWDgsYtxGuBcJGeWlGrhf0b
CnWUQeJdTGHdbW1rPgeb604YIDpSLC7sjkKQQXjs7y3H5WhoibmW4T/2EDpdAZf2
SiFLYtcDvI1X72iI12bAAoaDjwGPQKoa6YrlznsWtgj6/SObeBhGyQvK12KGFgvM
VfC0nQIiaoYud7RYi1Ckyr198Xem9YWIpOVh6Rm7xgnD4TY3GjmSafStlBaNRvar
NbCLH5W5xUYMoNlN+YMYsLQAqBHkrZ3UsByfEC2qsQu5gpL35wdDv2gqaDHxfFvj
hZPUhEhGS8Bwpx6oGIgfJST9b28pfoWQWnAokQ2OTRpBD+6b8FZ8RIH21uzPNeTJ
wdVe7XIdRMH2W1/eitDOBEPSXBCsYvMq4iGlg0ih2rf26W33FoP8tDUCVGflpr/F
Fdn0JbvBjpEQ93NQXMqPPT6sTChrnvDqOIp0S4PJ1MaF9tX/zYLz563iWjY/dwPR
Kcfn6d5oW29AIENNumRg3XwrB/llJ5vEtnanZp5bYLhnpz0fbSdPbOpLCzp8h9fr
hNLs+QBEgnG3M46AdQi+eF0MUCzvBO2Nolw+5ioYdgfHwOaVRwXKkde4SG5mFTRl
u9M4vORsLeNjeRcFbtIyPpdBke5r35abtaJr9CbYhLhDTS5tot2TmLi1UB5Ua/br
byVPmTS523rWebRqhkNl+BCjJb78fFEIYqbBqIU5Gqxs3SmiK6gUfzHaSQumjy2B
6EstYbNP99DFSPIXfA1dew6jvqY3nu1mYfoWVDIEUarwuPPJL8rViRkCFrIUrBTE
hUs8uei37LC9L3/0jP5WR6CeCYhJkFSm+mEaUknamcTfbo30g6I6FzgFnSJ2f0y3
0UFrv5c4+jwO0u37CuhEyZRPr8QM2fuP6LoJuLo2T0seQIf+9owND9ea2iJUwhC0
B4sdNSabSDACrUAoko1ojVV8zmQIjbyLAFxogfRRxT99KvT/QVB1skS1Hs8ZTwi0
X0mDkHdZe7hEgAZqx36OA8VHRZ/n+dyM82AwwpbnPzabrKwt8cY9RgTNMX9eIr00
gqSuYkQjXAWZ21/PcXehcG8VqeBsoBDqzCGz0HxQ2GdsJVeFZuyx4uS5yjv1rs5e
79OgaFA1gJeP+vzuCYiX6czNpo2UtsAgjNyhnbq8GeB4om+Z2SGzSEAsoK+os/y4
zv75RR4/a0zbX2EQOJ2CzVUL0FJRgrpy/vAIbWHFn+sbx1m/HLLhK7mUMVB1LDRj
rS0q8nAqKYK0VM5GaiqpZ20bJHDyMmfQeCpF0qOx/jbabO2L2x9kod17czPz0IFE
VBKZ4QLmQBhG02FHSPGfXFi5MNMtONr+Gfrw06DLfbuLn1ruBaryPd7OLjp1VSzb
NeFkjP0df7vqL+lwOFeBD4K8CCrReK0Y74bkF7BNvpHdFfJXK1Mh/F6e/8LtSYAU
rzTyGr+OyppKXOL7IgElA/+fLinDt6on6paCGQ/2yvnqmUSXdCioXFp4Xuu38rNl
86seNnuHn7RZQLr9Dv5H4bnQPb2D88Q6qycOEn2kFdp3SKN1jZC4eEzEUx9KmwXk
ZHvX4dHl369R/047tCxhzPnAXYc/FnHiFNPHML1BhYohd6UzwvH7OsI0Iw84baqb
mpoiZLQ+XAaigrkyV44Rv0+oFbHMcz+T7b0UnjgnduhLKOoTqwuzBtBpDzHZQao0
70UoUGDa9Kfexzu7kKRyon8tDCplgSeXuFL60QS45VHu1KaNj4g2GhTLCNirDS0V
gwfPH9Ju8fZSLEOfvjJ+oGUAt0SnaopgaFwa0YmBhWI+pA773I8d7wzaHBzOqBue
cZykgvgnfb0n173J1Fhov9A2KIE4xrqoM8zoz9L/0obrbsH/aaQajUj7FTsadRIQ
NsvA1cWeNZ3T0295Q5PA0oSVAOWDa1pDUonXEaGRPsEUr4EQ9B9Uy5lyjEtcGH23
SLbNZdcV5nfa/dv06A0TbAt2eDrUAhOot1GWMvyLPFONuQ6NxiRSQYWyHkWQFly+
sO5Yrqs+VWECx1p34vToT7NYLs0zztQO/IqYPxZhvDesgGrmtIV9qGOa30lVFhrr
Q6JPNWgKBalSqFC9seMGlcG0zb2EdqpSUsYfxTzcymTEeAV1ZU1upp4HdromC8Xy
G/A4uQz/dZo5JDPrXQjdoAiwKdp9NDFG5xMGMP8ve4f1YGqDawJnRM0k5noIbqsh
pGIsqA1aiP/Ms0QVbP2I2DOJOhuo5LQEPgiKu9HmpWNC6AzTJvg1OBzAhkXE+jTM
HA6SLj4Jk/M8DTJu1A3I2wcrolo69z47vxqJtN+cQ/JUtZI8d0MSNYuyr+Sx/twk
OlHj+75Dvk+vG5eAWtefOMkp0wxw/jwUlH26Hje4ZhatmHiXx6JJvFEMLQMP8SCy
cQjTvYis9dv6IZX1ddcqrwyxl3ZmaqW9uTkFhUPn5iMDi3Lg5BlrH003625n+XHS
DiNpcW5VnFpFR19UrwPh3gacONuwZ4AUdnoQ3yeiQkkLD0fCcfmLvc4WM47igFCa
kdYusDTXH9Mc3urCP+G0qk+6asFQmUfrn0BEBVFtLxwHLHm9vro+e2SFoSvLWUnj
f/Odv9c3q0Z2ljcp99POKkwpjJlaV7LmFDqin21np1JvUc1ZwdGVGgyZhMo6e0TD
iyoK6nmezJZR9lYXeyrdCmHTeGIRaFd5FT0Ef7OebHmv6A6T3w0YdcAakwuKr0mn
vbY8osz8ixJ/BkOAgRM8OZccKUS9jLyhWtmm//XgSxryHjtQd7lcLKOey+LcsEz9
byBlZc77K8kQ2B9TKtVgJk1IgfwiymwLiFX6MTpTViFZvwr2YFyvOHwgdhch4IJz
x62DoU2IL+jXhlSeRbLVshNKtb46qQtUJLNpCnJqOEqJGgHsslp7jI/MiGQK8sKR
pHdGBhy+m4kmOiJMFDstyCc6PFIZrjZzhbJEk6ZdMd4oCkQjnG3naQcpJfh90jSf
qXeJ4TerRWJ7wkImRCs6AK/RiH7BoRskicy96J5WuOMYACS0uYDGiUuYX3Zw9trL
Vm1s5GosTCR7I86+m4SbyP0zd2EXoI4LiwqoO9wJQ1PionxF2eg3NOAOG0Vh1V+K
sSw61OT2vW0K/VjrdZhEGFLafN2iFYlzBTmBrU3ZPWID9HTGTK3zktnEmqzgKsyO
81caltOdNGuzUut5dpETOXhlawhKnuvlos9qmB0Ui1EF1t+xLU9U718ACrLAHERG
26/21je1Slj/qYT4tsWYP6v4aqZGUI2h4Cly4G3A6WlB3NzlTPH0Z8vJ/1zdztrf
svKpUq4Ww+BP3A4vL10oyiE2vYGQGRtK1QNORTL2dOFVjmAxNSqSLLw85Fbl2jpg
mrEqtoKCSudZkIkvYn+UkNw6/oH4kAl8cskOBYLcCd0h/r0I2yj5K859t3mSYtWQ
a+Gjlcz+LqZvQKVz/DTpQsM9SOA9ZYbneu8mLHNBNZLBkmzto9Ln3ePWCivh+O4h
F8eDRVuXDMZqiF2L0pm8ZH9B2YB4FctSqN6FSiFNcROtcI43B+oM8Wbb1GvSMbms
9aAqRNr+A1WZPmsStmELxA3YU9ADeVFLwRWeVlnENlqK4nNhHy5q5qeJVTVORHTF
y6TJ0sdU0oGKUjUWCTFG1wrEGHjaRWZl3SmzTUFSa27WamzmRzYIATDNKyQpo3Xc
Mhzf69Zy32PSg86l4Y2dFV0JqFKveL/d59cB5Z7h6e7hvSqPBCHgOzRc+TSU8yIN
5s7h7kgDd4t7JEuu9FKy2aWpqU141/MdFBZ841uUeEC/13y6Y1/9kiT94KSv6DMs
uAz8FgU6BOOwSWKUMxiv6FM6nuQ9/43kr0293BKtgBbX+7yoX+i4+1lrCtyqYdaY
05j/s3Ii68GgJbQjPExbj2jmQB2pPSeDUFyzmScr13smWpxxzsHkaj1jDw848Nh2
gY5zZeSDrrMHANv9joHym0L/Bp5FYiPhb3mxjWrKk2eaLrPBVRLDSO8upM55lR+Z
GhbKY2Aav6n+Oj3LzlApnAq8qKAMQltGCWH2fGHNGvMXK1PE3TLNbQYy+CKwEWOx
t+g6jeNuPgyKwfaYGEfGSqn0eNeKi+ZQLmWHPTqeLx/5mdXYxT3UGsG+BVx9FTog
tiiQV4R+fX2Arabvf5jbA6mD90BsMLa1mJMMHcLhTetJbmV1OdAYuR0OgJuhYPJh
mkS20WIeo4U7Ee7K67xsvqMDyv4iwBLpBCcZ4CpDgZUKRJGwi5Yz22z0NSo9Vn1D
/O0X35DepQVFT2Iv4mJxByPCtJULZHuurVLCoHTjLit7t34rKnV7n1RQl3YW+eIZ
Sc+NPJXfy8QRSHQTUVMUyZx4njZb2Yzzo+uE5s4keRg3xysJ1Px3Kkf5IcdZhEu2
Xv3kUXwIHpGosmfmLnr4XBbckMjM2s5ABPUjhPGHR6PemxrQhP8+1AGpUzg0UZq1
srZNxpr2Op9SPCPMYZOn2nEvlJvWFFvk2aRYox1pP4Z+S+fzNZG8CSpvnZH8NkA8
e9XNyHfT+RZMV/Oi3iF0ajIhU7+EDQY/HAsStQH+1xu1Hot0cdNn7DJlpHaZQjCH
LpDiHwbZvmco/Jj7lnFhdNnR6z0SAXjfM5KLZbkSJo6Of09lE/2Zeyye6M1YryiI
c/ZwxC0qmQqT0Mhx+CZUwmCzoxCTBujSCdevW9N7C/v13wbILFw1RD9djhZs9pU/
rH9DRJhlyG2sMy2YYVa6bN/XFgicjFvMLi0xXS2lc2mWHEmOEeg6a+B6UgTsCLxj
iAT5YsfPSpoCFcL8gaB4U8vgml3/CGsgJyziqO0T56HOASiu7oEeOHS4Yzau8FT4
0MLyyCKtU0CrFd0Dx4yyiD5JJXjQctef2y+xeKBoF4osMtnUh45nCaaX9w+xp5zV
7PJ6tu0q/OsOh3xQIfbyWC0kx3GxMXPS78Me/zUWMqiUhHo/TfqpEyD11tyDqCWN
MRpM/+QmO7ddWuaRgWOwviQ1RejymZ5/jsRlhTN6cky3YeHijErUyt7vtvqQwDcq
1MQWAj1Oqbv1Fsg0avWtQWAeAClbWog2qfueRi3MwEsbn62/Xg9tITv1ZpVOP4a7
M0ax1P8hgV5s+YYOra8H70CBpikD9o2oOHh/CT/0KCX8GQgySOkq6+16uAI3X1Wd
JxNoqv2kP1TmjEFnIolbMfPNP7CMRtceaArGmzLFD6VBD4ln1pupCVxE1FkM7JXE
zOppDa+7DWdlI8q8MpABuS+OdZS9cbxZ1BQHNMkkGpQJ1yuTtrrmFMDCA43UCchQ
vfJCzOawyPFKD/8LcCW9aK9AMVATlO7LVlCRhxR304sCfwMq77DEtFz7w0ypKqbF
mt1mTfqfWdidOSA0wbZ4Mtr71FNyUxxAQcPhz6vcc7WHICSryrP6abmQ/u4s69RB
RljqbzE1u968PRGeUZKCuGo7H/MANEZaa4zrTVSAn9gnFdGh0y6ebGv9P5FL2k7c
6wzeA54tv8b05BS0LpRxjRNqD9Su9UytSl/H9puKagX3/0v7jhzR3ABgWp2miNjg
GhBWWGAtFZ+tCAC1GAwvHMetN4LfXEERfF9U5jPuBPgndIuaaVNi8HIrIjpJOl67
WTVStCYXR3DxJ3qQwHdf8GW4pzgAuuBTF0S+nZIqeYeZMN0GENw0167eQ3wX+wjO
65JnWHO3lI7B/WhPa0GIFtRQqlb8R7tBHqS8tTwcrkxHB/al8bqTvd+6YAA0VWE9
Yv8VXtBNQcJf3pvKWfuiZKFrWF4F2PAmY0e8fG5W5bk9xgossyQAqgm7PT94iLfz
FrKjJdVl/BgSh8tT9rRhlNKnvFlZ8wgstd/z8NmQ/KH/4Ppe3Qcly0Lc4Uzaev49
t4AupKVb7D+UIGgRtJS/4qKgrj21spTlT8UcBMpy+W7bltBLqA8Q+dlP8tkD4nc7
Pp+1KT3hxXrwIDcpSNcR8iyDtCK3IFjeI7zBfU2GDKct4gEg//aYiJNi1jEfmMmp
Oy3hY8rPvzVr+P1OYrWP2FzZM0aBZAySx0bAYY9+zdvqmxOvKwjtRtuGAzk4JSF1
hAqZcZT2iDF1gqk9IZfpyy1tZJxNZzhkj8EfJntnYnnkVJ7cctwK/y5YjhUd1Y2J
4C3TJ1T9wZbzcVm1ZJM+ll6j8IWpKEHPvNOEYKUBcw52MawRRYlIn7eXxdkWGwQC
wr1Sqcw24feP9jqjrplxz79urWDGLco8DLiIIOwY14kGzyvW/zQhqp/KTZt6w3eb
qugF0Ln/VrD9+TOZvB7PGNk1Mto+fL81Ei/+Or1kpI2jscQPydyYAalXrRcRaRi/
AcyVPCn5rpAZ++Bfuuqwwev/LJpOP/CT38FnHF6nH45FAO/uuj9z7tmRflNYMB5A
upMUQOHp81B4jhIIe32MitRh61Tox4ahP2G5kNExPYZYZebrHwNWLOLFSfuXtZyv
SHeb5VkOf1HqNwMIQOeOXZjUyHz9l57ruP0Gwe2X8rFHd6cKTpK8oNw6vQKzy+B1
lO3YlcOQTtZDJ5td9GwJ/j1JX1UGEwIXS5MF/SpAeVFcBfeRXo8s7ra1doIs8yo3
VKoaF76JuEJKfpwOD75AKA==
`protect END_PROTECTED
