`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCixRmvJaL8uA6qaVBshhnUxRCz9ZxHGFRJNT+bg8JKN
aKCyfhNzFTSfSLIkqrqUvvGKbzA1XSHwn3ZkaxtZMaCb27T8OqJvtAwfdxbYgE9S
/wO49AblTJ9ed7dOHmPaa5okLk03T4euYdvzKnsgXbeymOZFc0yY1iwfOtnWdW9G
lG/INYfd9eNYduRqn4BT2kPaaw+YUG0N7cP3mJzDL6zlP5BHXTW2seng+UE/8WND
hwZ7bYi9JCJl3li6qkKMX+A/OJQaxll6Fr0546/FDqTAu3W2pVpXLvj2A8nL/dQM
`protect END_PROTECTED
