`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
/Dxc6ip0P1wOibIjgjmJHIYSrSQDXfmO7ln/EHju4mWdBHwKXAxGe7VxJtnYzoBE
p5hQ2c1+p1o8oFTWLmNoioMhzsKk16TmAuMQtqYUa0B9RcjrT7RiHmai52YG4wgP
UmMkjt8KDr8UGJHwGl2WsR2DeRTCLiBIbv0sRsDEGsJRd7xs8Df2Vj395xT3RGTI
TR7ZKx6rgkqDV0XDmN8RYasm2DNZTp549QqZwHFlDPZOW0AFuEJR0DI/MzslA/Q4
bcrHeoAswpnJ8h1yuN+IqyP2wATtlwiM8iX4FAe5I8Y=
`protect END_PROTECTED
