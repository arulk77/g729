`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aQVqqGqsliHOg6LsZDbzveqqmyO46KvfKiJf4/9C7nTi
55tb60v7hP6VlxPMBhXBgc0vgZkqtIK3fGKqJ7ahZNdb279tUHAfFVVsnwiIEcwr
Uq1PCjtRKHkLS4MnXhDlmBCoUoLPV3f8iGm87no56tcppapl4PJn0iZ181WdHFKr
3Mz4D+wcFlX1zrBNqIV0LvxmLk2Kw2YrFnoHGJNOiLsYZw6D0VexLd3pAIkQJLuS
X0G0s0pKwP75F9Aj9Px1qBI4xbGKCveR+dq/ogrIlKJV7wM5gsL+kbCE8sBeM6W2
Zbwz2zRZGaI3108IfL1t4gsipqWBzCiYGtCmkn/VBOyvA/ngufYWExzFbIN6B+O0
iIhMdGvFhw+vq+fQb3WstTBPlAspO+a4R1USrZSH3A8ALIQsYQVtPvwKypPg9dPl
x3rxap8X2BG3fY09rhan4lK/UPckKXMsy6RkAk/lp+bwL3+oZI0NUVuyJKqybLl+
g4J8TGmIMY+vFldtCRGKbg6/xwCCOFrqds2CNADFwoatCKAQwqPorFze/4mJAbCJ
HnU91MTbCh5ekCfEJnjOS/jcfwPQQ0d7iNB6ZN6J0tBZrbF7Skg0K/xrnBWHI6Nl
LpnBXXkn6BhX1rjKCEXE6i80uFBjj6a1vDHLcg7loLHPv5cBwgmBtwckQJqjUgHb
E9DTIivZwkIL1pmOuGkNWGNh9WSn/Pr/Cx8zVqlxqNGl3x9kzphVJ2+ZiCk3lgPh
cV6L+OhRNOhbfCi8VcAhuRluOXtOVikayAqyzavRpXI/Wc6Nw3RBhuPeT4BV3RDS
chfH9jRfRBJbYGriiWGKOx5R70apit0XU5DuTCy/HBiZx+50F9dlDv1wzCmVBCAi
`protect END_PROTECTED
