`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49hYccW1s/9hY4iBF+v0mvyO5QgTIeBGX1miiXjQnMR7
yBsByZj0LFp0wSrRs7JxRRH0ZPbBJsgteoMBSJNb4rLS8f6OzEyOig+kulDS9gcA
HaGxrpVXwcBxaif6f1XxoZprdVmQW2aEB5fO0aYl241/iqbwZLN/P2PvkztuPqyG
hwZVN6T4DQMYYIVne7Ln8CSosplb8hXfRQynmOsjATictiSNJCw/iF2LrlrSx9kA
krQMK6QP220VY0BcYMCRBMoZ0+X4l8xuIMtn1N3qj/U=
`protect END_PROTECTED
