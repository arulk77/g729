`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43z59J1UD/XrDS9GFINXDdgDbA+V/+tJQz/QQ5/gVexu
TK6dL12jDyKgRZwZS2CcX/GRbuC8hY16Gnrls8UhLTKgmQiwnVc1/mfhLWofvDT0
P0LO9vqnJkJ0CymkpMVfI1r8Nr7swXUO7+n7epbnDHOz0g6sWZSuyUV+M2VKTiga
/XNc60bydC9qkWpG8rn9MseCUPwdAeSoFEHWvNZ7mN5f8RxBm32UGDcV+srq2zjN
QkGCP8b8Zgk6DwRRQdD5haxC7Cv8ShzNVdyjoaVFNRMHAiB+CfNHF/1VZrQzb8ds
D3vsLbQspotzY9a21noISQ==
`protect END_PROTECTED
