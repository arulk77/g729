`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkQDmYeYKO26/GZp/odfPnoWIs6MjAKtyh1yr1FD1t1PM
TKYp4O9EjER6FFcJx/bmAnXYKMgJxqkNNLbHTTLETuy/6dwO1SqmCWuxuwWCodiz
Me8LKGaPCOziKDGZdwv9h4YUHR81arY/FUTYlHrhbAawMAE5pTo8KHuNPmIQ3Vfb
5Bq7wymd4Lz/m7FJAfdm7TKsuUk6JCJJ2c1zX/3AGwSbnR3TIBHIgGzCBBWKid7G
NUrGbPf/QSMX9IxpionH9WPYYAhKMEuNKFvac0xFLxV2TurGNQIbmxA+/fZPnpLP
pjmYvnNb0p0SzI650HhZ+w==
`protect END_PROTECTED
