`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFY4Z60jrVBVvoY1E22CsncGovAtQwJs50M5HYCB+5P7
87Prv15G9LCdjPzu9o1hbZRrRuxnuXcvQ0cZF6rN+xgRZxuts3oKMTKclzXoaCsv
AOfLGz8MB0pniNQ+RyCdsDcb1wNiR7u7BaFPxGQGl70bo4P6nl2gjxAdIWPi6I97
D6o3PWsUz1X6RvkX4xsdSWZxDsBvhm6fv+mfaMDHRfbv83FTK/4os4dGkc/mHru4
`protect END_PROTECTED
