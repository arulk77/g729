`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SakcE53Bkx+jVMwAjG77vWnKjx5uj3nOO+5fJLrYEz6W
PU79qPY+HPpQBYQBYicyyG6U71ky+oo6KN0yinMO3GNyq8PFAyV3a82R8THz+C0Q
9l96Qu3NHYuakfQaV1e/z72XSd0ANMeWk9umUTWARapHOHPJADi7NIIM7p1L6q29
+sODddP7llUJx/tpL6HEUrcVbs7CTg5nB417gPLRIMLBFI+I1ROddOfgmlcE2O+S
`protect END_PROTECTED
