`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG8Zn53xbnd+MoLtUv+ib6UGmEAupWSPbOFTo4VHdTCy
SmgSywC0FkF2l58jB2INVC+ByEGFaBxQGP+xW3fxabbyeKOobyVX2uNovvPQsFLF
hFUQgljnvmLRw5j1SutoWGsl7gwXjTP/iyCwwBMcXLW7bMuCxq7JBMlMyyzftqgE
DMQXL59NFTr+YD8zcOvzod074FWsyHd5foYpkGpj9amTIvxjGgFsqDsOb2QqxUGK
AYZ2/Wf3tNT4oRp0InulVVez3syAzJAVS+1IQXxXYHL376fP7DIVLWKPf6fFlVqQ
M5+yClIqQRxKSW0GuAfCrOQtNeRvFYgXg2Et0lmudpQTDiXWurxSozQH2CbCid60
Gasuu8ibugX+xaS/5JAQGnEuhFZVtrCljTfaw8/BkUwEbEzGlntwWPsZWCjvE+q4
7ogdxVQ6LN4rfYkT8Flv50xrhM3RxClKgf/ud1r+SCx66dtekO6PPORwh/zxKnwi
Byhzo9cTE5VGtwfwj9qH8EXnRg8UlBX4nWsefFdl9bBGRL6KE6QUAQSbh0MxDrVL
`protect END_PROTECTED
