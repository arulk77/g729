`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveE/ptHJ6gFwPFp5a4LBZgUGIPEjLKwKnJDDkmAAJOTPA
AehxBmy6SOTL2XJ/K18rOuDsEXYri10w2WdJczCsSxonQ5nVmK10dDnA9NigrUxe
Pt/LqK67fi39/LR2cJ8XHQ68INbj9qm7/XJf+gcfNAYT+D/7bmsqpKCps7KDuUH0
dnGSNllC1089p97hTdwuIg==
`protect END_PROTECTED
