`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAeEvLqtBP7nUcTEzSBflIoB5/wp3QglUSc4iebwC5uKP
NqWX0qp+qlT1z5teqQKbXLIXD2V2lp92ynHeul88mpjCltu5j+v6KpeNbYuORvmz
iRZLS7ylLfYxbQR60m7iqCGm1gu1HU/RY9WHgqQ/xOs+NkbAcsvzD2eF1OiMOEFt
JnhjY4qPlrtUuovJEv2Wu2kMsgOmjFkunPAnRaK9r/LCNb21aez8adykbHN4z0et
O4N1qurIQZ5wv7DwBLwl27Yp9kkw4clKUyDmlyM4zTOU8tSrmffYlqAfM9FWVwpI
ASx+idXcsoYhPOZ80tBYrnOi7pqrJlUAT0r2W75xo75hR4qLbyAyVCZSM1WhXarI
5brL0dQVvRfmlBPNajYYFNFE38PMmT3ZMYNSc1IPLD9uirvxQHPccIf/lm9epRHK
6mBpMnNzZCkpEfnnZPAHybXXFt70hTuX8fZQ3WmDGZFPVDrDdwA5TgGcf3ukEl4O
KSOgFlY+d55rWu+mJJJ7OlK08t2N83/1Z7x5jC9/oakRJYUN0Vjs8T96EKVChljQ
sIsAQ+s1ylV6nhkW+TTguzfPpf5MpqU237LUPN0vpxPmbcM723ewXYWj4Ll30xIy
uceL/TAtxYt3EVHzWA4GYO/F+M976kBuzxMaIrn62oC6GJyvli/7/WkDVrZbbIeZ
KHffgV2j0OHVd+XuW7HlL72aVcaslMx2vXm8yO77dMYGPNj4gyHCchm24/SI9zed
PVZY/41D1plLnE/uB6GtAe10WuPAmu+J0Q6ge4rG5s1/kayJuScm3actquGCxfsy
SMKRrIhod1kMm+F9lU2lpTg4AdAK7Z7/FjeS+gBlFHM8sY5Llbii0BFdR7nZ9h2w
Fec7JK8KCRtRM4V3r16HRX8pHXV7G0QFIEFSBEX9JgW3brRK1Jwuo+1yT+Rg2Mo9
9y7plljF8D0s/uVPkXh19ayoe9edG3VkJexZQCPYEaRMvNnk2zaUSReS5k7/6QmK
w8qLTk9aWGVEgVl+/eUd3+MD6v8kPm3ibgQ6KZZkujJbdb2tlpJo4SE/j1qwpN8J
zMQFq4DNP4R4x34H2fiC8LEjbA/34BPjHb5uSQoj2io8WMJ1DBNeCshg1800h5+6
RYy9eecliH1pIBE99gbVNfJwyCYcfpPas2gucDE3l/CGQ3riwPeMZdRIERR/txAe
IWAl/Ht6QkNw9qmXPaux3nonW8mROHwgtyHpxmgnZZrCgegKn/H3yOUJuG90aK9n
bgI/z3/tDocJm95W/5l0D+Op8C0+HaoukxUslBOR7m2wmP7YZRRe+icfb1NtX3v6
3YXt70pZpqgVx6gC7XV80AQYfWCzrz7/zroj3xP6PduR46OjuHjEHpJiGdivSuu6
JkH6fXkmS3QzdZUYTRViEhE1w8qD7H1hFWnYYbkg/MBtj0npkqnIPHDmwvQpIAL4
qHX0WHyUOAKfgWkTvVtPDiZ37uJeog9s/Uu69EcGytLqrLEOoEwEF+SLJIqhoght
KudnRggYAqlZZvZMd9jjw7OM9cZ0RfIUBYP2U6EscEWP9yvQZJLDM3GIjPLnahqt
5WuBSJmVvyzzMQqSHy6LTyHGVq6QMTr00ambV4IfwWvctELRCiQq6Mjrk4amYzwu
sKl1xrTR/IG5QihasTsB+8fuCzqd+GFmGg+V7WCcUh5S5PWZEFOV/nAZQHzbJY3+
jMew38pfudFoUnOuG3oS1QEPmsRJaXnfW9/vshS/Zgd8oC5z7YRX8o5C3zKywMMX
5TITj/XxoqoWI1JZSY3DWaYP13lpXjAM3+m48mZX7e59OHKJe6caSQUVs3LexvLn
tob/7+8PL/J9W7eXvyyzfedW6mP4jyhTs43ZL+CQO2jqpe0FNmC6aae2Et0kNbZX
/w5OZSpSv/aRLF9h5Egp8t1mC22wr12LxXegfD/CI4JmM3Z/sJu7fj+fSOtZVziX
n68Q3FUjUUegS+fqyaahjCo86fsApG496QkGU1HUEhfBUhIW3ddlHVNu1Fh08KjY
SOi8MvwB5pCoE+efXnaFx7fpaX8Q1XW3dZBE7Y8/oG3XT+8ai1pXiTCkfir5u/aI
U8A+s27XWGFL7kGwrSrO3g5Xy/NsSH3HTcFeBK0mBOzdqI/9DBuZXDVn69FpexnF
oLItfa6n9H0Vp+KOQffq5DPwUH4HGS/UgrkuU4WBwVMnbv2sPF5x0u2+xPI32k7R
RDjcfSizKrPCxGgk/MpxMBeQMj4mmAQXsUuLutt5HTcPl5tC0un3x9X/PyW6aMeb
vnimsueRT5LVcn1y7TZ2VhEKqCRIG3VNyX/j35pB9gJhpZp1pluLj2OReyMThoBu
WzHJJMDFGjHN44qkgyEc+n/Dz9M9SRl9/RxDzsQTE2AyN+VbC6+oPrt5c9QMm7bw
KxNo9Qnb3YnUdVfNTrBRjaSt2kWqyYkUauuUfQHZ1wOSPH84VfnsyVaxXYAI7jkK
bP1Y+VLdguN/qKVpZzqtEa1TuvF79aPLVCeIPvqfNnAaybheMXEzcLLoj5ADoYmY
bRNAdN0qyyAPTMF5a5veus4prKa7OljK5VWQQRoPh01jhxJhienKijZ9oxMcQKPv
NYr2S9YFS8mzq5aiF6AA+9aY2eNr8VyvlNfcVfkiJtM=
`protect END_PROTECTED
