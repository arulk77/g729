`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePp8iAFerLvs+F4LPQ1TaXbr9zLdoU5ODQdMqdCHKHVm
Kjx4Ftdxywv6sfuouvBuu90A96LQtHkHStppJzhH/UBQfrKSvFOMgy65sgAIZaWj
aTP3C/37tZNtohK+SKeVXQ3FkYesGB/qhoI5yM8h6MJ2bLBkKibRUk9vyg72gfuP
G2dLDSTbTtEToTtyB6W4i6l9RZFIXcXl+5sZYKR5OtaxlIElHI78Lg3WKnpTSePk
GLsMxvWD0cOcdlw/eLih5/+u8MxDVCeHnwG9AG40vUGBrkDYG6lZzIC6zYUHEFjh
RlVBpoCUQaT19ZyLYbBsD6JHiDtW8HG3ZUxt45wRjJMBWVwOsmfDYQEiDwkcyCTm
3XdF2NT/FGXx98/k0NrHgP2ULryb2iZ4tlHlfzgnZG7D1JEbPlOEYAzi/DBqeMlh
xAC6J+lH/DqqVv/U8Hpfxw0hftR0st3bpZFVPQ1QBf4G6LhahlawghXSxK6zR6qE
`protect END_PROTECTED
