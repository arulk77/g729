`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Prgb+lMGK4ankHVaNnLDq9mOp7+5QOj9fEqACw8ACm/g3abbXkpx9EcP9G9ecO4b
58wtzS0RSX4IpnsnugSdSpqqrONUgbS2+ZWiusrl2k260ULlkkxxLJY76dNZPaOe
MbuzO9JfTwwS7ZLo7sfuo2TLoc/dItvSrhBicLB3Ia5jVyO80qlRHGn8fUicVD7+
3zvpfTIZC2BQx6Hz3dlYnQ==
`protect END_PROTECTED
