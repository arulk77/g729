`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEd2cwU+YLWwvHgatRzEb/QQztbwmB9Cl7W2Kxvoe4OZ
Pe4swvwcNjbxILBuQBB9Ee6BA5+hbnKaV94LvWjd4K86Br/SKpDuvWPQzDV8LeZI
zQHHEBp+QzC0f0HOG3cMYcs0+RVeRCSkShPl2kDD942yQkuxS4XTcu0OoLSEGuBS
1ziOLs7/0nBCNvbotlDeJ7EAbG5RtnE4yQZ64Dz8xRjGUQANRAJhwJ0W+Qrrre7y
`protect END_PROTECTED
