`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45z47xGBkAslooWhd9BYGGdlWFyY2r5noDfeC87fphDY
A4DRAhHwFpAfKCrdMRNiqnHORd8YkN7tpH+XQ788yCzP0jfLBqsXPJMXMpzgVB9H
nrvRtOxU2RyxAlqQj1XTKkrNnB0TjUhGc2/Dnm7fpdU2F7vgmj1W9ojgAf1yEVmu
Ol6EJxBHyQJWVMyTqh/OCiH4rDpn489hc19584M+0AY=
`protect END_PROTECTED
