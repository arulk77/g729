`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aQDHxc5AlU8Gvl7rUrpIgG2Fmnz+AqMelddHnKvAMP/R
LaulbUNVMMrsnwXjyEr4S5We6TurNCCR7F9HMm01ti71yv1lRAsn8mWuRlHFY3l0
lUQbjgHBMPMM1NLJBeDm+4SE6vV+WCKP7oG6jpnccQwxqNqRNhAU34xXPiLaqCzE
QDqzJfWFUTttkHGsB6WY/3QPySSInKFClU16sd/RRQWNf2KVVs+xkj2DYaBwuDFT
XwxYpQd6i2iH/34e+yHRhygzBdRw7Bz9JliVPVyb+vROl6iN5bqktmwTelu/1CCX
sELKoGdrj6jLd0Rjr9pAn5NxbSMPpDAVKJtV9+08K0qGr2P+TFucdjqpuxtPY4Ek
BrJJFW4lC2Armqi/y45VCZPTZUKymrguEHb7hdXTAKlbW1IG95rwbWEK8GQz+SP9
uRCj/ODP07rV22K7UHRoCfZ3+fC2lbr80MsZZeI+VBrYPxbug0mwMujYGLkTh/0T
AbohXgYSdzR4eUnCDPKEu4IPA1J3rBrfSZp6GUFNivs6zKFt3XyW6cpmKzViS4uo
BwG/G8/WyL/gkUCgfXbkJgtcCPmnojvUPZx65OEBcdAz1/uTHAedAqkPqtEgNilq
H5cKatLFJbMzWRBHL+plnWz55wrFzEx+bamwHDvHtNMQaePKgwNzB5cyqPvM0JTj
CJl6E8wWCAfYUJRQzOJVlD5BaJ1nDAr1rDBW0I7yO/IGfP4PoIOzLJhhYzFdMQQH
XHlfeMc2A9xj0sEoYXnjbkRp/0V295ie9dl1nPsIrV5dT50CthS+QyDS/P9WBEq/
tvLHsIk230QL8PGq/8kUxzucxPjRhB/I2d9dJ/gt9oDl3sCkbATgDbACO9L53Mfw
csz79yB7qyqv/qSOoVCKqaOKNwJlCTyZd/WyOrpn2o87u5BKIsPjkHTiJH3e7T3C
3CyFlD9TRy8WAm9rFmkGlLWv3OKsaCvV8JL3Q+rAgeEJV4u7kAGmT0TlWHs97TO2
HWXMwPc0TVouoAJcnHHYrovkDOAHfU9oTC5rwFlTvJLg7ADVzNuv3VyPbY3qFkVc
QliGUnMVvt4X6atEOpffU+Yy3pNur50Vsn2dSzp5JyGZ+Uqa38NIIjUsN1bStYzw
NsnnR5Df7eHbBE6248b6htO0dob+2ln88IDJDPSDpQ1UiKteFj0YKtaKB3vv7ylo
mJ2wW8X5Z8xoaA/iK/0sIlsx6PBWa5mWY2qKgs4xDp0A923MQxKLrTFVQ2RF3RoE
SAcB++L+y9EXcdJ2q7h5L20yqLzIXCoTH+TOXkM42Ts2QmdUZlAXzCFoWa6EKXax
PpMyAJNjLOUiush7wrCPaEHIkNB0Tt3L+w5Qv8jAgX0jbWalttxmOBWmz+a71Bqa
4GJfmM8LUxIQRZDSQhx2Lw8Mugo2Q37eAIaUZDKayJWMtBfjn1hzaVOqSZbZvham
aVX+4sfz3EXQVa0X/amWZOdaufBTb+5EvrT1X+eHD62aQ3t4b+XDQQFB3WRfwQqW
KyaHEMHHJeYVtlJ/ktn95XPaDMblloxJi8ec6BNdtzDzLaiU/4pCkB+DuxOzoi4z
Qc85gHAz1YUz1F2um/GTf3cllu7RtwgItQdxwAAPk/oi/KdisHKnAeph+amu7uP7
nBGTMuelwNZwm6aToglgjYqy2ZEMibNRn8sJjh8EVcLWOUTM18adqXGTGVNJUgde
0DYDSa+8Xea8+ZeLEKtmXQCSWJxOV38f3mNWHPnRKyV4bVfp9s9yW4U+5tYe6VT8
ItkWRMoJ8jyipRhh89KxRUhHvF+5w6nfwMMohOto2WmjXj0e7IkIBu2RXs3HY6LT
usSyBuFFYZgI71P+x2qUqOQqID3B5TjvjswKas5hGSSEtaSTjkTmmXmpb/4R0zNM
t6Meg7fRPN3Ee1lG+zG2S5SyP2abXUkbP1D7+F6eqSP/+SEls8Lk2g0D6oBy5BQR
qx2BHB2kj1iSFur+DRQeQ8WUHP9KPdgiggQ85ldtz4MbHf0uLZamT+HqI34sCKDg
VEmoSJaiApE0BX2+8sOYwjDefeLNQ2FY5/hYJusonlkaE1vr0pNwND4j/ZT6nnJT
oy1EpsWDcTgWMvxYfSyus54+txyPxDYpT/gFDnOEyt7YMDNpmle0urBtHVrtRQnZ
uVq1UWUwJdb186LHFOQUEKxM5PFoNzaxULR7g75OLMUiJ9tw/lfeXl/0XsalcyW4
DaGJMjziNAZa4oRYU69/FyaqBIVzVWBYxncld/lGHRvIv06myAiy7un3Cj/X8eC4
CMGMwpAwS7ywEDj7aS51GL3NStPcYyqF3LAIQvtssbYuK9LyDHGTTJJDtAsLj9c5
066jyeHg6v9icXqFsRNDMCSsjL3tgi54f4AHpABaCpjtcXtRnalrQv7Fc7u5Aj1p
eP3FF08YN/LeiB5nVOpMtdcvypdMm/MTZMuFySJxSh12EeDQr5DiJpCe7vwjUUGT
v6uIEIuiOAdieZAKI9BJBNgWuilylDWpHPUi7en2/RhqWsQUQ4UNJDO8QLcqEDo8
c+PbiiPq/qmsF0X6+m0NK5wqFPQwRzIZvwbXe2HyWUfczSFAOZ7GKl3Z2RU7SEEN
iGy609ANd1er3IGf15C5Q4tZ/3AnFuAMqAT5b93RuU8YXICcUTz/CTnozzbO01b5
f1nk4xsThVOE84UpOPuJmwXvpwaBxEB89gxYLeAHHIPhaQCUdwTnWoi2cDaxlfJ9
9mkkCrrV/t3eGuHk/fhaw2MrXwhTolvBse4QN5Jo7gHIT0MwQz3YU1CgqmMzIFwg
rMBlSESjY7H+kDnnid3K/u5z/vlyNfc36l5+9fCnTXOtIUc0YftXaCTlSIIBbs85
7A69hrUeJT582Eq9Mdi7NyQETAVKtHEUZNiA18Uo7TZK4pft6aqRtLQ1/Zq0gA5r
rJeYHiiKO83ybpwK3MfxS0TwqxOzIzSiiWDaxK3QBD0jtTAZfUtBDSl26YnCDUDK
atF6EgPrcaaGUocGFWseJoTkZngSEQrPBbR5pnn8+xLS7HIErHYRP7D0r97AwrWS
MSiopWvThumMeZ/VL6JiFfallcwLCxAWaJu+TqMeuWpFSvPtWbcior30sWM/DJAs
lDlmPRxUKMQ+iPBLe9rmWM5cyhbDAeea5s8oAZAJyjptlCntqG0sWiMSLHP9oKLh
XU3LDePk5qhCe0QFdZhSNqoeFilrI2DpMGznPSigc0ReoVOdPtGGy4rR3uxEkVHd
mkBn77mlyNT0K2sD0YW1afGw+KAqGNjROaWmJJvta60aqecD1RwV3mA2CU9sM0B9
xzC11D//5MsmrdROp/NIuaBaTEJBS4d0dTkjZ5iz5DQKhV5GdJqtPB4DAvb7d31v
MD89N6+r1FTqpb6Fe8YtiFarh6IOzan7nRjEPkWmow/kMEBwjX5X0tCT9RHWsabU
//HaxoTgl7dMKp0QgVzVWC1p3x1/UhYQ/5T4f0Z/Vwcjtkxqu+k9zL9CLspuXMht
p9+xxIGTmW4jDEYt/iGM+be5tqtA6VGXI0d5EYmC/Znp/7X6Ab6ptLh36wr7pJDL
W5YN1Vd/pAr8B3Bjq2Ht42y2BrknPNHSAOmWbc95ugZUj8HecEapHqf0CnBxwjJk
MdsukPiZa92IT+58IJI7TUMFtbJbS/9XquJ3z8mI/9tiCeoIQRO8gj8jfptIv7pC
uajjvFdSBgC/A8wIJ5ov+V3aIHdOSEo3nlRszIyOG5PFFF5T9jBMawVH5cq3KKvb
w0tQ9CiXOjAd0lxQyDoamy3obEXHpIC3CK2EtBM264sc/O0ux0KoGKFfjU3v19us
KkbthuO2n25nkuIJscVOHjgnSNSU35+akitmst9JR1PkPoIak5s5Cj05AfjBfYk8
rniRKVPgmm+tM5RYflJrvpSYQourCme5WWCsIDXRaXcWLSTAPITqimqglYHjk9E9
+Kllq7E/I9gRMThtIk6h9BD+LF7juYl4P7hXML3mCEPuqFWTQHgYk/X3G+mPg5zh
/nwIIQ7rqFc29LxR7AFPMdoXUQGygvr6MVFOon1Y6cDpnH9DchHR2zcVmXKx575b
vgnsucGC+ipYUG5JqOVH0BUsDTkhU7WxFMDnjcVeFMmRmc9hxHvdYsZ15EPM9ItT
4fDL02HkMjiVvHzR0Xc9XweiHosHSt5BWMU137a0ztItCJ/hymjo9gK3Znk3BoI6
yg6aCAP1SE1vGw1qu5j5HJd9PfXsS3WdPFk4MbVAtEac48O3VuMb6OjUTAWoR6aM
fzZsz/BD+Cr+u+Jtu0L5Y3e6Dv3eQGfWs1RzLvAvprI7XzaPPSE95j3uoPBFWzLO
ZyjkwCELJhBjw83SkWCkgZDWFIvBBbwIo+dvltUiBmbwkvFKG8hLUd5jhIJYU3ac
KozRZClzoBzlkFdaVZMNYPVmQwPRmocXPAqo8wdwlLZVQd0S5h5MdDPWJbX8XG68
g9EIcOj2p/1tMnjI5kDwVKAOnLINUtbN2FtpcLEXuBzq5vapr6lHDGfE/kWU7cX+
YRgql0RA5kKee0Va+wwomY3xEy6p5H7AehnPtlLI6pngIObSn7NWg76t812XD0Pq
e1GGDi7Wpt61XlrwriD898jA3nX++7TLMQB97Dmc1Rvy0fJ1oyt4c6dt7j52wMce
4atQELEQRNOEFdxMzky4E6uhrVZN5o62ua8tweyHLwI7ps2MBJYOKMQnlTsJe0u/
NA6qLwC9KGXXf8cBc4cqic0cn23EUgQdn3lSgI3XMWdKltgizmEs2B0AJ9uN4fJB
MSbatSyPw6vS32od2Hkq4lzsMtN1g6JiwCEN22Vblz5sRXlqpoqt9gIJ+9Ia6ZL8
JOEPIKkujj5utP1bBLc2UCM1cRusi5c3E9rr19tU9lpKN+QBLaifUc1thuM16p1H
27Ni6APoi22SyFN2EbBxwz2ASh2jwPtjhYIkuWxDOBDCwldGPLgZ6i495mMHpobW
tUbLSPK4E4M1Q7Aec66UBnW8I15+45wkm8yFHuY4wh7OECJRx3gVqZgExoTyiNyy
BKxWwNN63SQ3RyN8N2ZY3Yw3adHjwIAjfxWRS8zcOuChld+t6X5kQhYE2S2OBqSc
t1eilnGeoXWU6IGw34ZGchX4vdTrKmCk0D/kvQ+9yx0uscgUrc0GrIwaowS7CKMa
M1XjXqNCl3Z3PLyie0zL4xSSThnbL+BLCXT/mlPgxdwJVZ6jYydvFlG1FYStFEoi
Rjmfakt6rZU8aLfyZjqreo0LoHC/JB2x3BIaNmI0kc4X5+K74y29228KiwpySIo7
ijWN3Wvom1nJ+4IkuyDwEAnenQVqhZ8T+PdxaBqY06cSkwFDcJ9pHoQM292WAIXq
/zF+kxHckb8jgGmJGbZAI0fBMCciTMfH1+1KTSKMPPTJ8zy7bf7zqgKOgHkSwNof
uvY5p2HwgONCmgUZrw8ArXWSJOfzWbKH+RL+42Rm93/RuCbFgSIGaeFIdCSQjZ3q
QYDehsfrMBjAGllyF1fdVWkQF2iNcfXJ6qcIMp1PwwyQcY/XomBv/A6Hcz4hUQWH
Ol6duuD6RlJ0VoysVSrCzz5ocYNyOxbf3G5prULSlyhukDVLpwSbzQVmsQ3mWWkM
4pbFuxjBloltSehAQKTpldI08ERZezVtRoKpQo+tQf2JxOG7I1xD34JKdqg2kWtF
nPm8XYiFivaJ/7MFa0zKo0BAwemOQyTRXpmmv29O9idh0GNKYBMDgUzBC8D8Cobc
XRyfTi7RAcfljCiM1nYW+ylwmZpqvGB1H9k6VqL4Vzwh07bVoFhK7Ef0XOVXxaJH
mKJuVj2zJ3LwsU2ftZyu+WI3MkRuXIHzvFtVOhVDXhkmHUCA316sBGZBDVWaETtk
cNhtfNHNTM8A0AqPqr17Ss8ytF3dam32lkKDsdioUPKiUXl87xPYm4qn4XfHd8dQ
sWnl7dbfOMrEDrX7bKxVH7bkBsZvE9FC4kYiar+kFWLQ++YT6YQhPM0BBzJyT5pS
gjy09USsjKLfk6UEMXbTogO4boZKq6uPzmqXRcTSUNBqD+n3j+zDXkiUHUZT/HOS
W0ccDKM9G+zu2WTS3qt3nhnS3JyXB46FHkcmWrdbHO+Bo9CnheEQjzAUP4DTYl2c
Ewd+ZVaVJ162cr4Tqp+MLBAoGbhl84vS54pgb/f1Z3Xag9AOv9yu6kF9OzLqOLe3
WENvobpI+mnmiuuP1mrKt1g7ANIYphCB+JKToPjnSca71JjZxWaOK3vRUqCjEoAZ
9KtgZXgSh2RyvQf4ygiKiV7vovrZMh6I49fFkhxXKiBHCYUc5j87nRDw+qEPPCVb
1WzWabL8Plwtl0bpAFy6UVKnYZfZsUvwVfMOyMRkGt6rCnKi8d8+QtOskZdxPym1
eNTtOmyv/sZpSuCuYQl1TS91EG8hNstBnOZcf95CF8bx5uiDBbfdn6OzOxFNc3j2
8uMrzae2+mqhIOipj+A4tYVHHE+2S0FCQxkprd13BUvXcAdsF79j8gytk7OZ9xkh
rNCcL8FjvKGRso3/b+KuM/A3b3moKzz2cUFRk3WGJVfBzDM+xExkFe0EqVDk8ucn
baAjXmBQ2MEVs7vOR83P10yrEdicfv4jT3TTwRprPe1kl1p+lAzny2SVvRflxV8q
v/sdZiOgTs+3Sph0bXb751x6VBZistZfW8WQ1uac+YbqIc7bNaskCSJCWCMlg/rc
uLDGES6Dj9369v6OjdbRvU2bX+PnSOQJgEDxJ5IcskvasZnh3xqQrqPzTBXt6ecp
aYxyNvrPJcM/alMIoIIV/EJ/xqegrEEkXZQnUMymv9hXut992cQJJYwKIOctRtxn
KrZzPSwX7tJ3eWKpW06YygGNihVOndb7sWC3iAiFusKbU1I2gBbZXEYFX7QnCRKq
mXg4Behe8sVRz45ggsetu9MqXkNElmpoDrMINx7XabkZZ5BGxezPvCUmH0uyNsSv
G9nALErC5EbGW0219YrPoEyw8J0GnrWdWrA2Kp+mYNlCqNtrFAHPjYp7Tl4O8stC
mQQ7WD1Nn7KIDbCXFkGcgD2H7QQa3itmUseqWd/WuByVrwJHSfRo4FgNEMqLzfc1
arRL+O1EdVzLG+Hw6jkcBkAsIr3FHElDYq8rs4eHlkrqdNWkNe4h/OP6DjjpsZFT
Yp6eltHNxe8q+Jk2ISeVx6nAXx85fHvSQksUjWsrOHfjB8q2/4jUiy0QXJ2ytf5+
hW+nYL82qj3ndf8JSm00CRr3lRhHK5buHsvFyb22xjGTga2rqI7nr/HtZSGplOZp
Cx6NJg/fHsjwd1bX/d4y0o0LxTX8aYPYQMxLGGWGBIyCc6OGuINkFZNlpCfUdi19
oNNuQBwCjPOKNFJu+IiPczBcbav/tZxYigZ3nwzQEC7TeXWL5c9erXJKbv6CEL7x
v92lcx1s6A7GSmlky7IA905PXFJj91eop46K4r5vQugaqydtse7VuM2vA56N8/BN
fGlVBFvaJKvadn4J5QmDmvqxPH+Z41XEFer0IFOudMhhbN8AIC7Vhj4fCxsV3oY6
CEMwir/fZ5YxEBxGrNqXaZ8AhJ6f/3WV1l9P/Dj6xRd5e+htb1TkOInSJVvj8t6C
raY3l4GLlBTw9/oK4IDhygFgDzka6R/aJ7Ii59EGxFvlHhZe/xkZBhI/IOsfarBm
5gAGxybCLuvg1QzJD8GlVVRA7tboaP/lLrplRZzj1+DShR1qLxmraPptcp/1CYz+
NxyNCFnBXYnvzrry3iTVM0ZR5yZPvwJ9Cd3gLInVyQRzKDOOHH1fvpn3Dv8pYYU3
tBYNfBh7YbSRustCJqZsqgY06Sz8DU++MyS2xK65JGBs4VhTieyU7/6sked7mP1s
0FOeqHI/Z0GDFUpHygNjAXg/LSBLFgFZv75K/o28DShMRiMA6zR5UGej7qK54mcs
6rkiopyZ+h2tWn1vqIm10hNTB4FE4rQXK2TOR3iQ0/2nJE0i/Kr02OVVzquqfXxn
QngLo0zECfSmmMGoghoqsiD7iSPxglmErfLpd08VqQs/X3DBE6dzOY6sOrjTFhXd
BGpb19c74Qkc/8Zo+DRfkTRQDtcNTyTKqZE7jcr7uR2SGCH/1mkl2sXf07bDoy4k
96HMdTfJd+trpVJt1LV6lq3rogZqIiQEtUffJ5s9crT0+0aRRIHGQlTv3sdhbcSg
buz0AIMusm80kqamm+mvSsuRQqTdy0Wz1TKQhabwJiwbKqu8ZJUb9dR+dS2rTczg
dJTTi2aY08QQ5/sftD/YrTF1+QdQ8iisUIeWcPy1Eyn5r/uOgNANiQbVG70nWo6X
trhUMU+TnpWtk978566YvZY4m8J+oo6fvuMLrCMgjpJqABFuL/bMWPmySdsKEsT9
TCpXA13P/R2hl0RyqCJgV6pTvul6+ILGxSwbGNgS1xMRtiJhNZNlVtVgKlEtLXPS
S3FyenTkJ63pVYxnjd+ZBiZRzHO+S7ZfZmfa5Y7iTQoQfRbzzrAi+UMVSbwJd8l/
QeGBUQMdKHhwU3YCLZOfYkGhrjL/kgP2pQtydyl3tL1gVYzGxiN+T0VmU2J7ZKJH
w79Cg9E334BibxIY7nLOgSijFINykexCHdNz1UA8cAE9N2VpnbHiarmAMTLPaErS
Q5q7H7OYWzRpxKJw7y6fd+ODWPfCrtEbANsxAmb3LiXqK5xospBWVOfO1DmhAd9d
bOkbP/brjXxsFLfPrrPcEehJnWuSRoUrtTKqv/dmNatPVwweMQuRokAlFKLroVen
4OsnRU/9XbYE7Fsmud1M5qGLTap6p8LZtRt6f6nxQZ82FThVnwHmvg756qosnnGu
dS8LZip38/9DtikOb02gGQEAeviX76XupS9G2mvw1hVXcmJX21vl2pBKCZA3fnjp
F7/KiBeR9NiDPnxAKMIeW/OL+kBld60lwXtz5LktRk/5+COJPwmq3M3ty0QvPgmA
vX3PiIlNz9IHxBNsY+gbFrMUTW42oSpjeeHjH7MdQ4AHWeSnORs/ZeBIFk+GCLR5
PxsmzSmVa9PnEX0JsozoJu7qHNgmR56BOPdqMMJVBqe/AmEt7eVW7GsTWpjEYAhO
gjESgn6UCGCgOZeTRKDSSG3wy1Q0gpMbRIS3krlRoxXf0CnC3BOphB/oNSjEkVIn
X4v+2ByYFUtt3NfuCHrbQ/vM/5SklXlRSkBrWG7Awatjebc2sgDryttX5UJ1xWCw
td37ApRZ6qbQ/Z8eR81EdTFyZCeITnPrRMeaGcNMOQgPFLQEAXBKwocmvZqdHa1w
cY5oiukfzO9oSv66lgKC5cKzWE5EwO9FdSuF8JBMt6vldQE7IOLEK429i544X7Eg
IRSAW15T75BdYQD4gjSD9j+AF50I16R7QFDfKCYmkxrYNiNRTAXwxQAuiPMwN533
uMfqiISENY1iZm9Gus/Ts/fNTS9wwLRiK3Ropol8W2dCIgLDY9vacR84a5iwbvTZ
0txwk/KhZHO+big78aBiMPKZJY0CFbpH/9OSU9xlfr4JP1Vij8nTyqA5naB5SaGH
bbnC58dGetyD4IJSbB7pHEHTzLC59K9+48Ol3OtWwKDeazee35OCLlF/fdrmErEv
kyhPwFOhDsyZCY2IzQ036cSmTeREVYFF4aGftPqTlIt+pVbhHjed80WtMt3Mm7LZ
PvOESm+hUVoKeT/b3YvQDV6CEyy2kdPTzi+YwPCSRDwe1hj3dA8I0X9fSZAfPr8k
aIGKjiA65d0yd996hT6v2Kcqj5icTRDdG1SZ2Z4tpyevj8KJ07oPKipnhbtXE/1T
WPXtpG6umMV6kwxrg9NWMxpnG9bhCtgiDd2oROeajy0cApwzj5PDigLLmnG7Nw6c
9f2j9lRsXNPS/8FpVkVxtR3irV/cnaleEN9F/ZubmF0CUtX+OPbicy0JdyyPqelJ
Ugq9z7o9P5hasWwCR+flPgUKAG5Nz1979FAvWYdKpQGdEvqNayi0aRMccK7Gz/7t
uDmvoSqfzxJeKdMiPrZR4zNOmFQFOjnY2O8yZoenjkih8QaPwRDnIom5z7+1En/6
hBdRrmS8WUFE3xxdbH3JWg==
`protect END_PROTECTED
