`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SbYfJFPYvGMOgSXW/7nTk0zdUV0jXat6J+qyVAes6yGw
9Pg+ghCFK+eiVSIBsZVo3Kkh2DvtmkXWE8nEoPWWDBu6UxEfVrXh0r2dnQ9K78iQ
+5oAji7VB9pg3TPtjr/RvPjaWAZ/h6VrCyZMYkMGLAq/1S07PcnZu1oY6gt0VBYk
YwHVbCSHeATPIQ8n16K2LxD09swnC43F45RgmzqYhVEp2l5cU0/iWZg82S7kQNwQ
PmLg+WyTCWKoTe148TLtCIPfEzLqjcnP+S9F3LnRJUWlI2GHdTOmj0+KMAfRe4CF
47IRsHpmVCKXTxazQ/bTiMDmyHqlbVEiuVeN+Hz9NrsGM6a3OqdSHo4NWKcrnjJI
r0WPRt/kpGqSLGF49XhcOOeRb8iYP+KqKgKuXhQjimOxdhbrNZLUbcl5MjoQI6TP
KAjaJAkyR72vhgE/HfZCdDxcEcB44JKSBIRbQB1qOS/icoZqlLIo0RQkOLDq+ixO
acL91BMSdpMUyksC1/yR/2C1tCkivg0jnQx7YQpjclXXmejQCLXgDqfhG8LrSBXx
rJtXHt5qo4fPISupYhiy/9wQs9LJZj1fpy8NmRzRxSB3lPpaSsh5KAwxTx7f838+
1dokF3X4vQcLpTbf8iv76rSyvcihS1n1XKFZWGpVGLO1W+NUowoOyFZQrC34pfxX
ATdbMtERRHbv2QiVyDiYI0CARkSssO2YRXL0ctSQZl9LwHvaG/8p8qOEXsKy+mv3
912zYZoMbitgjRw3J30X94Sq0lOmLI24+fH+igj329jihgy4NIw5Tv9Uy/2wWfpc
w4J6jcwvD0wU90GolUDrdqcvwUH++R61VKt1tq3A8C7Tg+mHwLbiYA/+NYcmtKq3
uCmbDOnVdcRBnH0NdaOOe7P3vRsQ6YC+VhKEVOxM8L/BuV4Jkm0lefJeitGWkEvf
Y9DqTszyB3Nl0fB8ByPzoPx+kf71kn7SX7eBxLwwHvVOgF9rrnLn9hEZzcmzuePm
JNPUgdzDUiMwHgtmwHgSbVXj8dVSZwEA8+2OIpBAf1ZmwrzTetZPsioIu6PjmsWz
fAvomlROugZUxlL2B0TJXHemyfgK+OmCEMulyo5/A3q52Z9bca9W0EK+XwJW5CFk
WmqRWPzNShPs7YUxpkm/vSR4DY8xvQVJgSM8Kww1Be6UT5bUOxrxLf6GM9ScJrMB
Fic1mmGxDn7ib8dFgCQhOppqZk+CwnPao4M8hbzSbxrkvbIFoZ8gryTBRbySaWE1
e4CyK0v+/rPKuVdPpF5SyMFOdZIQjxhRpo/lX704cGtRDiBP+7eVHUhj/WPkliEr
cH/GJ66EvW+8FIHR9t9lD45MM4nWnOIPa+LYQSHvUk9Bcv9jjarzpL+215by4xF1
jmnU1Pm3JuU8UXas82wsXQn64+ZFrD6JL6pkb4VWu5WxWYCeEksW4aYZYKqQsAY1
wAVI1SsMmVxP2W/E0XrPLrJ/yPMC/0mePVRaic0pFT2vEj96RTrxmxuPMfov19J9
aVUmt0YMyRnRRRutYr7oxF00QZ6c5ffVkzZalJmL6rsDMUntLJKtrw15Uz2UprW3
f6X/q/66zyGnizDG0oUDhBVKj/095qjXyQJTzN4ys0evbRBs93ND/PW11ZZmHYKs
hyGzUGuFfqsJH19SfKOBbJehybm3dIfXZ3ZvMIW+MLcQEf7ynQg88e4Pkg/EsNQm
Y9oWAvwIoqi+sDy/zgrbbmNFOUGE7QaIs8pVhu736Z01PDI0cqg2wzf87EMFYfja
MdtZoboEGXIiIxaZc33qjjAcvhXjBVLzQiiI/ggULtOsGDwQ1tYo0/GSDNjDQNlD
bAKP0dRr0c4UnDs9v68g7dvNhC9kZ1HJnevImfUyCHsYR6DIadnh2gfOdlykA1Mj
2YjeJDOCDLf1736ON7iVXr2gxEqUR8drUJtBfFBVbsAZIarE/zOLqGqKTwL6mxH/
9zQYqU7tlhR52tTiHfN6C7j9D1g/kUhOK19wxv2avcgeJzZtEc4ZGSc1xz6J88UG
leuQi4+llouAPFgi2JGqECpRiJX7Az8M/OvvMgxQxCV6Qkcc8MMlCPoEEWsWoXVx
L/6hxD+pHjtfdoKNW2g4wbo2dJhVhJ2pm2W1jG8/wIpf8F3VXJitIruD2eMT6WpJ
dSqYaEdOIJKCTD4t0QmzalM+Q1onvAPbGumtsfEpX0j8f8IZzRUbKt90sLqJdO8A
KwhWtTXWUXI8gkx0QwyJwv6O53sEOYamnSDog3hK7ho9vV58ZtFcSseCTlY0Tthc
Hi5hMO3SBB5NUjkcmDVK963IUpivNoft1KAjwpFtCLQCMZv6ud5JOskN0BSLHZMV
pQhvQTjFMhf9K5n0Xl2r9F81tKTZJs6HOLYnPoLZL7mkeF0d+gisKaX40muTGY7S
8gXwVGxBN44G4TPsmMhiEo/55Duahd41pPvW6fiRoX/xF4njSV2VrYCAiJyZrp8P
EKqXb8MesUZwR5CH5WiUYC6LpsP0O1KMaDJZdhhpfbwmT+zq4K89o6hmZbbRfU2J
DTle/UtB6kNfQrEDnRMlHE1v2avDkBHKh6pVssDleRkdUEtxZzSDzIWQlOuIIa0n
keqQ4HdsSy94WOxyNUzB9/khmTVw55gaj8syDMk7ImGMjEl2EiobfaGKQCZPhKdU
c6/lQwRTnYiaQwg66ihaVXLNVN8OjUSO5XW3UafW+LN5xUMP5RpuJXf3XAbJEJx1
9LRYwhzFZL29tk3FlKMeuA9hV+7f7sZsCQ7lQ7tiqqtsVs93Z9d3k5/5X2otYRBb
UOiDK8sdHv3lpWdEQVLytgOV/XWQBuAu/lRQ559hQhiI9S32q0aORNOVvC4ISTvN
xmTakMqtxve/xvR0IZjFyFfJLwta70RibXg5oWgTe19BWhLVMDV1Xp26tFEd4GSY
Em9P3BW2LJPG4F2JtVB5ZURGFh3r+sqtn4xlE1cGntF/2lSiPF0v/tPV6tGcBLGh
McxXqeKyXfOPDF5I6oCl9DS3R639p6Nqmx0TMf2n9M+YXfjbSGxxPz7T5obrnNGi
4kEOqBDAHYyUvEj+dBkLipFA2BJT89lB5gJ9wXC24zyooNY6rQ0FMgKTRx92u5Ea
d6Q9t57E3EYRIEW1xtDjRIfO4BzMkACZmhm51UDxFvFozCeXmQUhl1qeyq92yGKF
DQawGrCDt5HKyq2ZtMMS4n9tZQUvW091G7Fy2azkOoWSDrMhHinzl38ts+DraHyG
i9pBf9bvfv/MpAdmpvr8vi1ez+uc35YK3niYnThxa/yl/8Id4eh9FkQN+0fQX1hO
SW3ojOTK8a9gyGkEtamOYY5Uw/9FXZto/OlOFsN0rZqNH9SmyJjEPeJpxFuAVtzE
6ywHa5by/8iP0PQLs/X7k4qmosd4oj7uPyx3Ny/KAQfnVfjg9r3uuBqy13YWalup
0VZtaiRoMyaE1xaPtXAW2lo4Qe8G8cAhH0EQg4yPn65/6ja23hyMqsP8iVP/WBbx
424rl3MceFxmwLRAt6V9zCWEUap8gP7+8VNSVXXzTuHnpSD72OyC/ceUVk6HPLab
Nzq+e1vjGp8m1IWHTXDDwC8epZGHzH204a9H16G7QldDi+dV44PZENX66tbSKSCl
7X6vv2XngIZsbzCKwP1jQ5qGzxmSuGUuDFgEKc+JXMMKOarLsvWxOdU7CLCuRaJc
zIRxLWWKkbFD4rNA53I6r+84P3m64G5CD51nnfk7B7lCPKSOc3rQT7udLsdkk8uG
gGk2g5O0oRTcsUR/ZUCvOyOCGkvvCzpy47i8DGNCyZXHjeXiMnu6Otgc1pVJzOVX
GvULO2fCIEGnZnqZrxN6n2NXI/jUZpZBPfN8Spnty14rwYNCCidr8aR7jeF4L2Dy
r1lbNtx4aTKgXGHrFTK8BQLmW5s8i6k4LpTtrfHzIOfgj5W5E+Q3wNKeUTUT+xsJ
o6OfV2BWUYGvIwXJ/55MvOkDlfWaC5ytMUYKyOCAC9n6uc/iLscbGIxyT+2kEUzt
IXngoBXRM/P2YnK1eq4gOKNnYSmfybd3C+DO2tHH4IZf6xPjiCKS9WsT+U/qSqXl
KrFDYD08zoq8Dy1oHJNLCNUTgCCmuytwvd2aiFMZ2wc4XCQPaqjUeDeCFtWe6aLo
b+lAZqA4Xsu5N6CPhUKDRPLk1p+Ciem4FhdVMiWrEraur04XP5yF0nfNVlfooJ1y
wfwr351RAjRx/9nWVp1VrvAH0ZSpDH/WgEq8BI0243f+HxXIqrBydiLFqFYqamjA
RyNz/nBOzNbLy78QBxsUoB69YrbLWYVT0IOIGIAph2B2hqwjwnTYaaolcAMNwERU
aNHGA6EM0J1+8HXb3vMiyzZlqa0sJW9MJJ3R0M9y7nPlTa70AreOXUZa4Bb3GUHk
ZgMofn6uhU89eXiZ9y+DLRkivoy/yZEj9SnLBmJ9hZzFq+SDRG+XgnyRVrJTf9Pe
38ALqQeC+u58mfQmC2TONCkI87/xcDkzOBP49eAS8lOHV+GDZt2bqXNwPijknJV9
TIHBvmchVQhdGCKy175sQjSKrIfE8RnbSykDz4KtUJmyLHMxhCHKF6RUUOCtMogb
vkgwaRz4Vzme2N8CQonmPtvdvlXMrFBVKOZZ5OfSKvkUr4UBT1j2Lw3e8f8dtbXA
x6c15vlM9L0wVSzXydciHrwsapk0hH+AwkGEyvz+jq3uUF8FvQrL6G3qlqy3266z
oNHeI8piHLH3cRmlqlvpG2cYb9+X9lT0fO8ffwfekaDr+dbs/TWlnYEFVS2Yw1DB
M/r5652s5vSlfQRJHOwuwO24sD3tY4LSbC9vztLzo9gD089wzggSut18NWhSm1Jz
wOg2DN1LpACT0CCQ/cPaUDsoGLWIk6Wc/lYNFddj+Hl012RVjpwDahbpgxVl77jg
/Q0plGIDHQy0M/YzcYBkRQDrG0tIOCvxfCk+5xjGUfscMyU+9aCrCzjsiroOTUjb
VdBvFVhPp0YEvbYzH+Qx2jZElEUa5Ya3rLtJ+uwuBLwolD4VxpsYgbcllZjZn47A
inREuZuYuFPMfPc5IrQPpWDKKxd1Zma5Ybai4cilRViTCdploKQNWqEYbc93TntX
xMED6+LKGVe2/JMXLldPK4Qw5gMoGwNE+MW0zw2A1YoPV3GKPU1U3yGuYaszCZ3L
x7atI+o3pnryXbhZl54o+pAVKhyWMpstdhWUsX1KXvUpARWc+qCsxKcQzGXRb1Kh
qT3jhfEOahp8Y0NC8LZJeue8h+llejQgq7XnwatDRWI9jGFqHBK+yGEZmJcDOnjX
IWTsKiBIEpRBkIAqAVRozidy4+drm5sUcksHNSB7IEObItqHfjRRqOnqlgIJcJX6
VG66vIHyyjOgtngDB7sI2VTavG5LfLqawDzory8cjB0oDVGr6QG6we29cxLR/cac
UaI6UyChHMnAkvSJmtgMmC80goIqV6SLi6VXbOl/E9CxgC2J7ZNx/2ex1SxXCwzu
1c5V1vECeL8vCacITRrYOzMdxfRsNtnRBGc0d98hhUCHloAOaqEb1U+PD/RboVlF
Sa1zYn6iepbTd/hZ721hTamTwiHhjuhhuOdPKGLZtVpgdx8Co0feCYEQCmgjpatK
3duOcuLoT01mC9wVjXp9vc7ACmdRcmEJJh4QUJkyWpYSf/vNYbHQTwa4PQCiMWWE
6/6HcPavQLXZX+ncL+ozUmRFQUF1mA30oRPp90mXkSyYqh2eIt+We5mCTZcf5Cb1
/cHCuf+YGCJ0QSrqktl3m7jPdOYl1PNpre6Q9SPjvTVaYvpdMOhqmi8Q/vgyq7in
7rpZu24zvSuATW200kIReYhhYqKLtDrHn39f1zd/plkQ6ymgMzE7trh+5FE7L2ge
kxyOTqt1ipbk4O3oqARHK4cvF+JjJHiXu74ctLJkXmvWrrhbS6uy0l+CZR8Rlinz
gOuWElwp0CBDdhFH5nlCwLW9mQA2vv+LQ1SRznzHFVhIqvRAY02Xx3IHvQUtwOaY
J9suQpif9m0AKmf8T1Rqk2gOuuRw8L6iSUXzvxS2JznvZrtEqWztMJMzVR/cXe6b
ppQk+jqwVl2hPgm26aGDl2j6apbYLxeDgoAQ8zAaDgoaQvRg2f2+q8F0XvC/YUQi
OOUBqVTPXbaISBIxF7Da7qz/tag+uXp7y++vH6an1rcyWWri9mFJSiU3Q8w+Rprt
z10qW2SkUjGxjuOKAWA4OqqjtyzXXfzniNg+9nZj9Q9/4OpjnaF+LM7hxYHv7FEQ
kO0L1TRmnf/y5ZmBWZLVJo+cyGWWLOGAEELBWsJusmdrVWZ+hEJKnK/fkkFGZHL5
2Aelb7sUEKni5rX1XiOtsFz8Boa06FFb8QcXCHDzwHqoyB+2ugF+LN0z2IwRVY1m
mfzUr/CyXepUCE7ITGJWnyL67c9JYCzPh7Juicgyq5xEtcL2vQumX2SUn2Woh1oA
+qXIsT2O4sNRN5V/D8j8o56keGppmPgU8asnzV45ey0DkmmoK7qSYLFjbOyrcuTx
LrI3AMAWXhoMVIf2RQE7vNWJfgrkMgqNNiRc489/hVHOXvUiPnsfx23tO+GyWTM2
1uVtOkmBQc2BLjGRgUBnMg7y2KbTKQGGXSngz5iByh0vPkZZN979DaYBWR6P61co
lRSA3oM5rDpagfTA7JhXApDtZN0Yf6KTvTBhys2p6gT9GcfJGAVUT3XaYGCJj0vs
6pnH/rQ5occRcRlh0PUbkc5beBB7LaojLUTz4sOI8OLrFb7tIzORNvlylkp0ov51
J2ZOQkhlFnO9RcRMXM1qj6NeJxjId01pK08jxriFfCSav1eGfgsaAqycsJ5Qy4QG
RJHyIOUWtvnaV0qbs5ULSCT5/4Csoagk+KTKdLymBZRuBLhWoKwLHa68qgndcjGN
O1Fa8j92jgl86jXjOPvs+Hdt1e5IfdovyfpMz6WubPAnExQj3+X9RIBm3zR7T7aj
TUlsCkgsXTixHrZAvDfL62KPtYRx2Zy+AfCtr3EhDtevU15YEocAwv2Lr/raCJj0
M5Wkz0dPhJYY+a39iA4uZxI2hg/OJAkgDp1lNuvW+AeRR+XEaILPiVHRI02OBykN
3yHZxtqmzJYryRxBiIl7BIFsAkgA3R3Ejthd3W8xuQeAo2FgIniaPDVRzJNk59Nb
bjyL0jkDfe+LbmeLKrEtG8oDTpZJsN8HWrEixXSmFhsVbMN7+FH6d8OUBVQvtfgX
dQEUt5fURzCyeXNXHD01zA781PVAG/3fWe8ERBvqhHw09IA7B2QVkVuZJREu9rc5
xr/rxE3zKP3qGxaEQRHt7SGmwyfNJsrzNpf8tYlCQ0ex7SRUZ0fmPQLhDlm4BIti
3pk1djHbOIv+WgiAuF/OGaBN6bYznYL6UFubndx9dY8S5OTXy6cYYKwEkfyG4dxy
nDuLnPpdFjK/xz/k21CXI11y9OTuYp8oHdMgmn72JB0I4TPHO1w/eQ8f6m9ZQF/x
Nto38d/JDMaVKYkokw7+77PNHDBKrMIqO7fsTc+QOyBbex0Z8FhXMbFwP036zjFV
vs4sODF+K6t7FVUBJdRa0nmdLaSnE9MCBeDa9XpfNdtmLWTw4rlznGLk7uI+qd7O
QJbuLPWZ9EQEZS/WeAcThnUj33Jr8Fx5pyvANdz6YbEISU+c4vGXhLSDL4qnQ9aC
Hg+dtp/hl8PVcN7wYummyV5fJ3Eyj/7xkih0OAF41gaiinFN/M/DVgx2/58gfPwL
tZ6q65OSTfcDJSMLSMgBb7rZ1Fs/jGqAXYTufaePsar6W485nODq+7OGuqRuKfo8
eYiatMIrXM5RNinsOrb3Rvvx9KPACm4Y+1/ZosKUhjMqjeuNt7WFSzLJosdhOFpA
JPPcIKUEo35tx+o04tEwFLrtQmOLIYFn7Rj/YRMZbOsZwI71YDX4yVbYGBcq37yF
AfDuIzMckUrfOkB1RoUCPVNEi63w5+TkTX+Ngfq/zVKkx7RzeltFw6Ce9Ckikv/Y
MkbNflcxoP0OoZepX92/3UmMoPLf5pWCmgm4Z/S/kON/zNlheitskBhRkdfrEp0W
27b5rnpoRqpFRZ+Xo3PPU6Mxhe2T24ImwE+IoR58G9tPPIXC4RUtKxQzoulOEjY8
JL/AC8COoxKHhOQvlTGyTXZ5loQvoLQb3mTIWDwcnqHHkZG+5GhP51r6PBxxlze4
EFIEmTs3tT+t22jEWEVRDvPGHGbKgcB5KU7pof6yNA7N2wA5Q9ORtFd6/RAEx0Qr
C+y9TwvTKtrgNWIQsZx/Qb3dPC/jvQs43rmycHgU5JCo6ppHF4Bu7hNYiG/584NH
8pk+MWtkgx4fI2xiwkNMFb4w8X4c4FvkrOxxMrOLfytpGmPHzV2FTDKQ3pw6jruB
s3504Ai52u8K1AvwifHwLU+VHZIhzG7ZUhIQyxUU9nJ/oXGAiHXcRdXgA94YTWdL
e6xTiutjmjBWzD86M3G5F8m8jskevCfHckCjRo3bYygUJ4vXCwZOb7gohXyzx14E
fXgPdrxsOhTx1dq3XK38Iz7vDJ5L0IP7twsXzeMm3Ndh0fE4dXWfhRoOZiMJUTCd
tHPgveQiofKEmdqEgqmHrrCYrxU0LxFV/BZNZdk7u0rkYxbUnglNVlzCfshboNyW
Xd1MQY6xNBBPXAEPAwg9VoPmoHVj3g/xaotfi1oowZHuAKf9Uzrkj6wYCw0pZQ9+
j7j9Lc5uGrIxQKzej9qOQHEmgB5AM6PD3aoZhq5R7uBrkinGi13sSblolchSI3oi
9VhANN7jgWSpDCq7Vl5JzL3iHKsPifCsbPkS8zIRDC+dkhfCieV346bQkaTohiw0
YoLwjxX9wO5/f9N6ZSPXWyrUGUS4QBmfXnaPKy9ic0U3STohZTdrXO10f5XNT5IH
BgWyqZKxFnWa82wDwFZmKvsAZC2nhwT06A0NwF8xOn1/2KrIO8obsHeMCknWyG6P
+vouJ7JvVaIdhzRveKLawoUCtAU/N+AmVPxA/MAk1Sf3RfXsojn+WZ+29paYe45T
uZpofRr/7JknrTq155F9x+DFlpjr+ClqhcHkF3QPTJUBj2dlJf6dCCBgAieVfMLJ
kqQrPgOzwuUlv0VOkFKuRNoJJXSOgAb7Qc+YH6ONJiPUwHalDLafi2o4awaNWVBS
qN7fQx1LXKKfPxCEjtwoaBIaClp9aHCrmvB999GwcIbcSSVgYnT7nTXRBpfCG9pH
wmSa84oZ+pkZltdPBCa5IOOqPiu4wcpZbH2LAxgyaC2aEMR1+Byo3pbDtIqgBScB
kp487nRMDLN47jn5ai45Ct/R8Se35TjXu5ZFBxulaWtjcX28TCBvDZv6aaoiKoDz
LhOnK7WzHQwzSdnv+xxEpxYGIQco7eoUn6cwK5Wt86+iIHOyFIxooGIpXpYspReC
5bCQzJVA++tVUOUe5kS3x12XxpQSVnUI+iNcUlA8s+Y3KzFWqlLhhneL3YuOG+LT
k8JHiW2k5QIFNTIu8wF1MzaAHDQ28SlrrRQtQABgP+ii3S0yTm43dw/bU4H/4LZc
VO3h5hl+E6Wi6YspVwcwI4yoQwn153+Y234pfUHfZuMkQSZI/ioDrwnojBGS9gWb
50iild96cHODqzz39d7o+n/Y5SCymp1xjYoDLkHWz39YIQySvp9u9rE70l8aR7yh
9vG36813eMTw2CPLnxwCQU03yc1IgAUGj1MYKsqz+V1KWRhN28H+sQ4ZTQwCt8KL
TCl4Ssfjnm9Q99Aj7UfU2PZFT13v0KU1uZqgGDIABSUFlL4sSvq6IoMTvJ5M6Yvf
SksXz6YeYpBxN+lPWcq69rPiqwMDS1U/s4zhd7NIOuBC9xmTFjhNwBPKuRckKmWi
Fx6O56NaJTLp//5lI9MMzYHiM3WkQw2BAqk+qRjdKm0Q4TxtO8BRhqMwk/RCLpI6
HMvkkAwIxZfAUGEAEctb4WXHHxa/njc/sw2HUDwazICF+iY7C7/EqTYPvwo7dqri
5OJ0NTqRZJkvvcux41kvQ2wj+kDcTxXwM84Pi03hKhd4SEXB9aJz3XSIDPyYZXMZ
weetRZwvEvIbN+A9b0jdAtvsorQgu+eDi/GrBqbdTrNtkUtg9QWisPI7WCM3P456
rLC+yc+zQ6ZtPf5iIOzpHN8MMFyB6JBhNjBcM21gXr1LwKNcnkOJXIradrjn7tN5
Thh2ny57jdcMta0nywmiu8gMaKbe5xckm5/VnhIjZNxFTRzDofC54QYVi8sfqGzQ
qGp2GpvT3myLXoZsEFgs7/YbaLSoa2cbuyFDQjA2zqh8+AzWInQUGhW3GL2/owzi
tG4zMVZwcE+D+1mfQxYLF0XKGbfBcqGRIKRKS1BWGXsAnvoNiqAReDnbEGmIXe+F
BplQpTuCtoJ5jdoTDSz34E4aIPh/pIMzFS4arleeAsZrmDqJ6NmuNOXDRB4VRYrR
/5fwC9LTsvitFf7uLfLsejowWHbW2aN9zV5euIzH2B3lR6vxeO2dLv2F62WhVIfU
AxKeBeQV9JKzFwRedD5eyHQ+t0H5yEkLQUxfpAn5J5bCRV9q77VvQtmNCSjzfdoF
SR+h4PWZNQ22eLT5YCxHfyTZnlTf478cjpZeAe6yO0N5vPyL6zPnKK0p0TsE20sX
2UVkL1j98q1kYUnqH+6rJ/4KECilXxU2gtO3QKua9YkpWF9wYd8xtC7QbI1Y1xdj
U+tFNucnMnfPL75eE3wf/XyI3JTnTxCVrHrblZnG56qUDqsrXtHsQhft/InZeeoV
JGNsa3Cyt2G+caOHKPg6vjGO4jM9VFKPa7asT6SO9RTpIhtmfVDa3A8sucIVGmej
thKRJ/r18qKwkAxD8VRn1RoQJbOcB9ln+W70qJLMfQm73pZqGu4EG6Gk/7KVmfTF
z/Mj8uq42jf/saFfrSlndi6UbIpsLk1nzVBTs4tzfWPi5BysP2HUEt1GhaYaQarH
ANNFR4tZaw30xECTQR9mjIRY4UCakjKm4YyAQkuCn7okdGVMC6eGRQbjS+S3kZDW
bnU+QzXr6a3RG6zcBzaHXswqwtif6soJz0eujlNSlylTZSimffglwFzH4Swz+S/6
hpBbFnHuyk9eXs8VBVqIL98uI5KHYizH1+xtl+bkblYTtfYWnQnkitt4ZCBbcrtX
KnVNq/fPRWafUHM0e5cNGorPf4gdg8Nxm0+rKTmJ71OyEUM2XZQgcJvOIqMlrz/U
CNe8CexcHYYxLnIraYUxHQEFH/JzqI5BUrBhddvQSWKe6UFcjlkgOZEJmD9Vh0FT
OxZdkhhU1lT7HgWN+3ncrSwT8C/SPW7YrSRpQ+WbbD3VJ8thPfutMJCqthfS+5Ns
GiZz6TNxca4REUP4whAG2bkpaA2hphnNTf9FaYyoJhU67/u/9wokXZ4Vtw/7Pu0E
qwVXBbWERgRzDXoiL7WPp8aWDiF2qXABA9zaV8JlBIqrZwQr37B98+paGObH9mc1
WleTto6eXorlwwFj2COYP2KAW//yZv1VBzj+TxbwdcuMtTTL6lhWkmkA5zW92PZh
D/2zYKKjjH+yqZZ6YMb3hZe6hlVQNN5FnDCqBOXCvsRr32Zm2nmkBafUsUTrzikx
PH49xsX5IV0sK5j5NSNx/hrFuXaen7EcO/13w1xwkSpFEmA6DMB49KNyXkOKDL7w
u89xbrjCMpBKCc8yPYdSEKsDnfBm3h0R2vVRHj//ByLgyvT4ugw/6HtT2uOqheGL
zO5mHVYsQIftBhGzxkrJlL/XNFqxO7ufvum7OFGrUsSrXme/EUFSOl3fGvMT3S29
Wph7hYtD53CSFj/u3WmfPatY0peHjfqSoBJ34oz2feRZwrYakDZIUHnvxF5WiQAG
Vnw/tIA8WijPebl7FJImOAdYCyBrypMFrEybJqLdsmOlkQuznQvQl6gRfPvLi8yK
+GQqz2xV878bKTfzZwVxqTd3LBAPqRczP3LPa0HHLSRZ42LhHkQzwKO96We+PyoU
NfXIBTUwmkif4KWOuEv4j0RX+VOVcg1HyE0nobx/4vsBFiZhY4Azxo43bBpGfUEC
rkalzmQYmDgWyrLhW4+1bTf4Dm9xQkqJhl/U6S44UIBmmHlvFXHfkQpTOIo4RZP9
vqVH5X9NCcyVVKheUjZrak1S/NXMPcgPIiz2ebRL+XSHjaxR+k3PAZ7jBB67pWS+
8/MMKnF4VWkq/ObGYx4jIAHECgS75EiO9+vCGiWqq3IDEkK2Xuf+HXWWfA2baTzi
JrO4ABQeDz+wKMZtpw+EqHGBttjyrqyYgOm1E734la6GKgCpn/eXBZj97Jx6w6Tk
34+9sEN78tVa4Co/E10aNaBSrBTFtN1pPfWm6iVeWbs2md5K2JgDbf49kUqkN7I6
Xurj3l8eLr+jOcRQ616HHS+p2nLfbYNGLymxl9x+Y2v3gL2nuQ1BIamx6rRjW9CM
rySCAJ9JopeCFe/I+F1LyglHumsTzP8rmRCHfMVs4gQXFwACfSfIV3TohcnW3r2d
sDcgE/Ez1ZJZzWkpdT+YRw2cBJjtQwkF0zblHiuq39VmVpo+D8su/+CDIBq0Td77
3BKq4Sbkx8lo2/oqywx8qyakaCbaUnNwGkg8OwCoHKNMIq7lnOofB9+0RY91iBz7
SvglFBwJrPfaCJJp/bCxf2o+07In2mTZR4Vl7fgrB3px+DDx6Lo2ONg+U/BMe1Ld
evcEIh7LAkaKsvMk2lKC30Ac0BP01Rh/fCizcEeLs+cr16PnreTBn1y7w9AvVXtj
cb0E/0uIWd/IohvMYvTwb1xuJbhA1CttCAVttipANkt88eKXhgdPbp0aDapGJmRi
5G4iBcdtOjbmob2NvP2ZBbIXkb9NyGY9gL+PAtIWkAPAqd/BJNCzgBdXP9ag/2UI
XzrucEi7ht3g7xclO2AS+vqlEEAHA46DUPz6M0IN0LBkKEtG44qx08ODire2mRRf
S0PdA5M8ztRodh79ktrNFOR2bmEvATm4U0TQhilnLjBTNBfcAVDUb/AkvR3RQf07
eWGN+2NOBT3jJY090n/238WbpSpvcnZvu9U7i6p7jnOdjjDdSWc0FjSIlPfKoOeM
hIKMdLW4c8B6M/lgBDlTU18pPp/cjV73pqDtIUmWkLFs+Im5dC/yAXjQiwWRPL1e
uGiUEbSIopzGKT6nCjNG+xLjpG91dmJUxmQy75fcK2NcBwCAVZ+Rk3L1OMvCo1I9
Uz3vZ/KtYQnu2xHBNY5tWkDqP4XIk+dIkjl01xAhMiVi7RTndzgigof8AVZdiqGy
88+W8Hkubb662bLykcN1JR6meuDav4ijFT6GtOzpjSWTrhGQwa5fUynuIXrOcvh6
/HIcLHv2EvmflgtL6hIpU1ePUBAEL4UiYBh+Fmo+8H/MZEvh8/ZEllL/Aziq2YGm
FsdiNdVH1G4pWyfR6pcN0qS6bXn1E5GOB8OA1ld7EfoA9FnMdjf7lVMKCdRYTteI
HU0Zue/t+slkPNpPtTIPlkLvJxsF8NSFH3v9tWfNTt69dkG8AIaOm/qjwAolne7d
mYN4i1dTrn4jIIg8PmItoiWH/m3DRwd0RAJ1LRbktKtXV0819MT+BSCOVGbfjc7z
twc0wcrV+3y/jqeZSeQYBAnlYjtlFRafyQBkjjJ3j7us4vfp4EXaucx2Uv40qMMM
/C4JHxPgBVgozsjdmLOmEou8Gjy7ufDYCH9MRGqg3usVL6FuEIONkMHUdftaisNT
FfvxG5mV3PDhpT8aK4fJ2ldezBSgPHbyAlpHy4TgpIyTBAhDJy4L2ULbeUpbLpf4
EAyLLlkYJwjTT2LrDWwW0uUlfK3hWnAmLwBb16wvPlgXOYPV9Zmdn41KkMgsSN1Q
4ObDYg0mNfKazhy+Y7qlzq3r49g7rXCHpwxpv+dBVppN7CVuaDdAzrAdSwayjMV/
25kOqtumZnYA0CzCW5jOSdwDRI9m3bzi+XT0QJMNrXdZCfIzr/dNPfI74RMxgm1L
yHDFP8u8r1lBazQWF+5/5OjAKRqUO31BVrS0Ck0xd14dVez2YJ45Z8PcYrgeKDaU
AA3B/dGeazv5RJiI/XWSxlF2+0o5bPuAoEEakEFHcDjom8Tz9q+z+ecYCmyqiU/i
GZl/eYyPVgzx5pQyRZAJ2PjgCzLwdKVgrCQlUIo5g8XWvWw+XmUDt/iJCbyRmkN6
jKNjlctkc9ACUOmBTJkgEAlwdEBBxRLhcEqZ1zd58FZ656MCZFzfRFBjaERGthS1
w7STmn8SRtZ2yW+rMybf66oHNd4nDc1IRgni9iCnXq/OwoWLGEXxXzwKxISa1IU3
eAc3Jg8MlCnBPdMMJs5WJIohwsR1j6/kgM4X9tnsVkmZecBogYH+RMIhsEQu4q07
8XUJBF7zZyJHo+nnWa6A1bKyPSHbDN3L1m8YfMfzDuA+CZyZbpNoaf9CBHteh3Xp
F+J0R36dL8JSYhlj8VFp/4yFeISdOnTfmwd5/y+07ka7yoPj//zYbuWfqJv5vjU0
bolKOvJA/t8fvUb6thsYG2c75oX4zH2Hv6H8CSExC5NilEjJ55thXxTcI3hU4tU5
rJDdXgwE3xV+TlH/PRWzbyLExHYIvoVxp8UHE1Bh4/HSp5tCYQdz4+pUApfUSLYo
wLT36E+KADYtCSSMAM4hAKAFqdPNasXJqIgNRYV7hqI4ei8FhW/DGsIA14BEMW3O
WYQkWumX4cWev5mYL8yjwQL+rrz+h3r8JVYci2fJ+o8syM3rW87lcnhhd93crQtz
dVYk5FFR+KvzYp1JVzTvmCRMpAtMp+0Zd7TkEpGewFKZYilDiR0EoC6DbnZUxYMx
ZP6hR4gpUVz0Cqem6oerKUz0BHwHHGwzuNVhH5W9qObpeKAn8W85haB8CIvIjLkp
nqLvhKJk41cJyu+OaTrlCz+21e5J9IcsTCaQWknIdLTxwQzP7dyG8pf26cGM6yYh
dqPPh289RyIZ8WwuW2gS8zeLu2e0iM5sPxJgUWyrEWwafAH2UpsnmdGWpe5uX1sM
Qy6dWLknenEKsY1AzmgSMMWO0Ry0FI2sMSu4JYXg+xbjhR+JdHQl7Tg8NWWHkMCQ
2i2hiMe6KQHkX+nexiLC3ib/JOcoWpxkb7RJg3Og67fXJLZL27vdq2tEKy7KZiXe
NtkreSExTE+/UWOHML94dyFA1BFKEzHTVtBSJ5ugCoJc1hA8S4k5u8PafYw9/wD7
w27z/Kgj5FBt6kfTv00ewGwtIhfxvbrsYlMnvaBFtYmPtcIVCPam24ELi2aIdXid
CcHYRf/WtKaXMMsvTKs4Bxg49rn94/jtWFfDLGaDjRf9vNeHJdYPmjcOain9s6Fb
RQNjBAuOZEh8+LavnU4wlkQ3JaB/WoWqpp7imT5YOgEWGCrlt5IvYHESkhl2IyfG
+1/5Sx7jyvi05l1m/AEL3TMU5D/bhY8if1ACG61DNlFd6432ch/sFGzfCabQYZop
K70RyEbEASUQxr1XHjbUUUhvzocM8grUXGjRSYzU89zGhiLZ47erD2NFU/1EsqKz
KnS1i0JHCIHAoZ9brzSU49pTfE10R5jmP/uzhgWM+YASqsjhJSiTyWAY8titQ/Vt
EYXDWh/OzNHK4pfFuAp8DcM/AeSyC292A+fN1SQhcP7hrEgsLgTatw9nw4ljak2+
tvxChlpVzjzYQcMucBf8bDfqgnpFauVug4r+egY4Dl9GffcN4e2kkh+OCUKfXMBi
7DyWIukzNIy7H3PFFgR4utESRdsaJQbQ5vUf9x3Ymf6neVo7Qp3rdvjXDeg+ht1l
QYLqHk0aOS8s14AA7csRhJ3vRaUm1bjJ+3kXtO3gUPibR/7XR8fJs8GNNSqT2etn
rKLYe0cG4swrrodSIZIM+CHp6A+rNb67JC32GmsDJB7kORXu6DNqHFYWsR7H1wpt
p91wM47ON2jduYb4tVnpd6ruxQz504oI0aUGwBDwS/CxdNB9b360HcLa7gowV7TW
4md0tEDJFXEwG7JDt50ZlrxUYoSrIIS93rFyxltP4j80M9g0qKdvdqhkV7kJ33yG
NJXtUgAQw9C7V52ZcIookTsxxZZZ8Zvv3e1yx37wb00ROQCrhu51Ec2DIr1EnZko
Hv67dr3BDw5sAK44KggGYVg8Xa+KfMhWtT6VPkPSP9s7/rPFr7yCXSrfApEwh72k
PNZXtXehOXVffovRYnEm4STngNcoJoVEH8RZIoxzCDArn95n4vk07ORj/GU0NgAr
1jrPdU5ezMbHeb85Df36MEdznJi70qgdFFuS5rH87Z1KzZeZ1amHumTzvl0sKf6+
Tb6rF8i8uebU3CPBEzvByiQU5NpuNBARDi3CXywIuYq7C/6mFWsZGg6VpimLmnb8
5ERiB54MDgILBBJSZQhN46cRFtq4cCB0o1j0WjT8kjvjMmeWBIPHN0qb4+n6Bq3j
G3EVyeSHPk541z07Zy7EWfssXFACcYCb8Zef8GTkeULIndWxhEoXxGlFGoEgtHxu
VSyLENyS7ybvTSM3sSCzQnj8UHmA1XdtefDK3khNCGf/usu+K1xFYpKDUMP/phr8
mK+aBhBRHNjTu7kzXGu8u/UPeSoKdkKoC2ysjMYUyfsas4X3plHSBOMpvsSAQUuP
CFF3jCuYTOGBeYUA/jH1zJWpsNRIpdp0fvCRVwZqonUzUvM23YiWK/C377Uj8/N8
c3Wvay53boGSiODuHciaLJccbdED2BWhnstwrQR6Ymm4/ty3koP+JdUDEAtCOkll
T5gKAaKe3Hl3cz+eMv6aY5GUevKRwm5JMhygVhGsmhg2R3iRnLE9JHBsmgfL8/n5
G0BkPE9UtWvMVMR7R+stjhYYVmXbsLWTB/C4yvx3M3PGpqttNqgBw1DOEbDJ7hxB
cRvtRHNHyr/ssV8w4IjSLeGggrnzXVGpRU4bMgGbDZ1vPn+DFkO7Tz1vc4D2g4Su
OYUZ8Seo9MTpP60NCNAHPIicj5V8KOlKFB1VlUUHY5pbt4PRbon6WHqLn/3aQdgn
FrUmAexFSW3IegG2cQ23x9nqYbFiSVtP+cY137wbNdG7++CvAtzqXlSO3JqypCQN
m33R7K+5mzbDDPoIYbO9CbaG6/f1zfSPyyZSZCpYSk+VOw8IjFCIWn53wH9/mLAw
AqYamrmst062VFsEEkINCYDhf3YmOu5HRCstB3q1wsHfXf7T/8pXk3EoRNrjiutK
YjKlwKeDVJLyyz9COoBUruhWkPWnE4iPDzdDBbjrEJmPRcAmi2c55EQwydZJ5fmG
`protect END_PROTECTED
