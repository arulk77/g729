`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB8Wc+WUFDG4e3zNq2LDmzOA0m3mkOvQw4JtTdy6WQzz
aZ5z0frhxqjwdEqOTLcM/W+r/UWcI4OsgVwIUwTCZ/dsf3ZT6Dztsi55QcGtACgj
cyke5gjmuqpb/C+1MzleFoWQwN9aCltbj+2WITc3Ygf9DTEblDBP6f4uIw8/L3GX
UVutaqqCbBuv/XV9sNYVYzgbf1u2WsQDKIZDajXkwL9rxwpZUTxM+gYelbWMHJmG
sJfWb0PjXxHK2c3y75qCi81Fq7BoPyJu6Gu0ZXnf+70pq58Y2BKx5leu8d6EiClR
4Zai9WLQoVcVkCU2QO92Dh1BamAMkg7M3eBSDPiBC/YGwq3ULScCQMxHXJdkBcPD
PDaaTUDOuxYLgM6S83LBn6dXclJs3iU68bk5Ai2uzrlmjzcNfpR+jFExsUneHfgW
IT0MED9fU2BvY/hdOBmG2okz9jZAEU4TErh+kK44hivxGrveavGVbtwlPnkYhEPQ
XcX50qEliCef29sWKTwj7qHwizJ+FW3vpottYVMvQs1eMSQ6YbAuRoadVcbaqS4D
GIHzPSeEyV3lAJ0IR3JwBWhFNI52QyFkgddokV9a38JHF1m88PKRFGEPiD53su1q
G7Y8bGjMJLu6nUVeXL3H5Q==
`protect END_PROTECTED
