`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIeft7VxJHeKRyqAZrv0dC5FJVBIEqlHUbtO56BoL66L
R4/9KtjnER8fwXstcXPQmsBw9E3TyrvXLQIE2WRs/SwsUsI9xSkVnrQcalog7Q9G
4lo/vietonx0vghT84wMGw8c9qxnTHX7OVAHIHcOi6JOPSw2cEFPPFH+PpATYvdG
LB/Z5tsjwfESxhZQAHkYMyMvJHSNhP5g8g6Tf3FID4D59nNVVP6Ookjui0U1s3Wd
esmuj8LmM5fNvrL/sxWa+FHHKJtbkGxsit0EwtHw7p3IzOi1arsl1roiyiwTrbcT
2isGuuKk/FQ1Cz1nTERYu+e677zyAJd7/PCBtTdlL1NWeY0ZqlmprJ5bJaCEOtRR
`protect END_PROTECTED
