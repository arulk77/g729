`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOcgLmP0afu+gIP+hHlLmWUBslk/PsBWQWmqO9Xjksl2
9DAjKDgAUtpuW7tPBvR2GkdD8diNueD2Ed7jgt69vg8BWL2OrqtANIc5kFh3ufen
19iMMKYNXWQBk4IJUWCOQjccUk0UIDWZBgkidHaYIdHXb0tabZURkMpVXCgwH6SI
1vaXxoz4YIfbT85ivnQaug==
`protect END_PROTECTED
