`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAErzXkNyM3K280VQU/w2JBc/ubHNxMRQe/h3HHo9m8O
PEXfPkL7nG+u8aTDaMLr0pPMr3CrVieFbyTsPxOKq7V+YLfv3ukxbmBk30hWlut5
PRSmeIGKoZDcjuUobpXkPa2CNks/Cn3gUqfmpq91AqmwxW+ra21Ak7SUb96WtN6L
ogy39Liw5QVha4lgt8MN77OdqHUAO9kf6p0U/FSDsf6VGaSv1bTbXp0gAf8nK+Yy
vbmPjTxCaCpWLClTX5bWCp0wyYbDZi9bURfA3Y6SkYf3g+dxs/Zy3TSvo1+d0d5L
Kqj17BIAcQ8o10WPV/JXC91Eg4i14IYoGInDHBE5UbvqZo9pREp8y9cqEPC8c86X
JlscWEab+i2EAbWMU2+KFu8m9n9nbVfL00gwDDfBA0zUKOIYhQLzHozJVjxf1zhC
AvPeDOVPk0nQAvr9Xb9oGeIYRu0uGQtupL38lIJzXk+rtMxcxw9ykbIJPC+OhmeC
AW21bLR7bZKA0ltgN0Hp2cwMT0Qs0S7W2KqbsFX7LYI9fKoiHWYNSktShqcfewx2
5vyAqG51QbI71lga2mEs7tXEN3Fo7l5jHFi2AD2c1mqB7RGzXRVQHn+FbJeP/JE4
kweRTYlVMojfyMoeXqjPv0UiSEJcy1cS5du6OsJmTpFs/YWc8zgbJ4XbP+N9yfK/
0NvMm59XmDOcwXGTngpp6JjWf5WbS4tjTHyrxuf8BP8dxG0eHzBCJKtz9CvbpbdR
pqJCY75L+fTQGNYmR3TM5OIlisw87Obuc+v6hNNxnP0u5dPIelQZgmK6idY+8jn8
z3U+DaPCFRbFwM22JvagIx3JRgZSDJG/dnq1HIEUdnU=
`protect END_PROTECTED
