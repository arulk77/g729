`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42NseJ/465epZNikbniOuHAy0qUKbajcnUMSNv0gcEeE
MBqQRSw/uouYzclp+WXXZ6r/Fs6LcS27b55G1ui0QVrypVM0xrOKBheLteifqdBZ
d2io0MwzT6zuMWAO9TVfsM8C1dVcqE+BpXb8oLrhjhnTvjArxpv/CLrx3YKV4wSS
jo74s68jENqSoiOV1GrwHQUvMmenQzuvia49mdp0x7kw/cARSrFhJAO62qqhYzaE
gH3ymXwE1pTsASVJCq0H3s6iLFruAQbDVW0SilDGjvAIDhlFBXCGoJ4iOGRXgJB5
zXRGY24s5K/y+7OiEAKSUx5ywKyC5QvIq6BHwcRZfEphvFogI2wvgJjdlpUyx79z
Gil58M3Qh+a/gwCtxyrKFg==
`protect END_PROTECTED
