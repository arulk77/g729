`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zXSLyG1R/gHSEAEikbGc00flCqM3FVlqnxZCmpqufTM
XIvwCUnio420v84Ct+iaBC/eUcP8Ces/sn+z5wpYORupH6GBwtiJQM44e7wao46H
irr7hlWBNzjLw70HXOEPB+B9jIQFb+QUnV0TV/hYXK01TYtsN+TXy977/cNkPHef
p7SeLM9L6WAykQwAOlElY9VtLzkdRADBBtQdMmIeHNnpIIfKSmnQlhemFf2HqipT
JilMTpLBvA87NV56IeQEC9Ppd8jr56oqEeOUrnRvbZHwXAmaBrFHRTThS/fDiagY
xcZ3pjsj2kHm41WI9ZKU4w==
`protect END_PROTECTED
