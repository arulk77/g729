`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4x2D0SX3D7QasNDvJaykxP/wbyH8CZlVFL3TlY0mFHVC
BUj+4Nzt5LzJh0GmiFH2lzpeLDj1O6LuRQEvu0nVzCzYXeYVte8a28qPDyEYpewH
pFMqJOsRy9chFcny62O28sfhiPkLT9KH29TjQ9HET2nllthwyXnqsN0Eh9ROfnO5
S2LF/3F377ecD3lqIdi74jMCC/l1T0i4+USuq/CFnyFv9T7BiKaTrc3nS3dqKoHZ
kCl5WqUDERudWjmeMqZUVOCSKL/RBHszY3bbp4HUBQ9rBdkn+sqYkeAHYyFITYSJ
IpWgZP405ZWAmeYADusqAg==
`protect END_PROTECTED
