`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAXDpSX24Zw7c9IUIDWgxKdhUsrLgcwncAti9E5dr0Ong
jsSFLJeVIyshIX5dUVpZyl8k2yVaRAE+ZwUOG9LCclsubys0GnXUU4nt0fUQsMzi
/5epBYMIJYTNi5VHyCudcqipDJvi2wjRj4/JVtkEZDfEQ+KGE7+27+ZAxKKZstDg
xZ9apegIe7qPlld6lJOPe3mgDQ0hgJkDArkqyO7Ig9CyZ+QTnR/ZZoJTlEDDnq+F
1E0PQINF4A9TGIkG66WPRK2rwpwsAVCai+r6vmwGEECTVItx5551Bj487FosX6Ii
1v3MJw/Yu2yFGxVIlwcOIe7q0uWxQb4B/eAHrMSSjCFPO+mkyCQ9FaINc7EYiT80
l5thnsdcHVei7+s/yGBsSgHPJoYUjV7WxEAssaFV3cwz6V1suV1s8fcGSVYvaOS8
b1IA31GU9wxR0ZsFO8EAbmGqyNHFZbnhGGJVyaTL0YBNaNsIBY7x0qln6hy72iLs
O/Fuqpqd3l2yI9UpW3B9NeFo9FFfInl4MyLMlDosHRI7ZuYsO0uYz5unFQZVy1i7
maK+i9z/KqEfFzw7YPbQ2CUJHL4R3FReGR9kijeAGM7wzGApdWB+nkUYG6Y6WT6f
aDa22OWBYwuRPX46Bw8Qs/OyLrYzHhOttERafPaqXtJn0fUUjT3VjmXFHnj/K0PF
MCJGBd+uqTeXn2KYglUYtitKhEcVE28ypMdMN05dO1o7azPFJYYXr+DmYJ/J5Csx
Aw5GPWZrPTKUsJGmgbM93WJoSZTqotqjhelCNKatMiqMHCuVLhn8QrGkF2YJPUz3
NinisW3xHsGx2CC0Cj9Z+xKARB1JdK8eonZaxYXDUgb/RLWsrL0otmUqwPcnXJB2
a/AlBv1Xtg0FlC+UtM0zHr9DbvhD7eiZeDwNTM3/YTCT9NuXWdkMPGRzMv5lg30p
CthM596HmZ+jeZ30bR4GmaflBR27Rz4D4wU+xFzmThhHzmaN1ea2y3DhAWBxxpWl
MgCgGN7lE9DkrwX2IM6XqWiDij2Vx6/HSeqNuruGUi+QG0hiO9iiRc0SRpq8VXxI
+UcYXJVQ19PRaA/6If3Ub39lIQQ7DpgGEwfPksqQkvEkSfqmJ5XqXxQRmPySNb87
lXEFTI77lpGCTL19xtKDYYmjAqEi1MyaIDKcM6GYVFHmZSaMQeujTTSL2/91QOch
KjxTaM4c8sRXxJpL0DE5uKw5/pjLWzlhz5Ab7yhK21sdgJ+Yk6K775EMbMLfwk2l
MbOsv9rkOT4DkFnRxMu/mBTSnKmlnStzmREsh6MPPt4UAxgbHrTZeZ1jzjEJoGBI
Nz19CbTZExzoVogjSoFzL6vjJnM/VRvserKblU+BAGISKKgm0p3lBrEXjuDPYTni
KJotH9+DxBxf1aiA/FaM6A==
`protect END_PROTECTED
