`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48gCXk/THgnLlLqJlCEIjgGO9J8ZSA9v0SaR4Z189xjc
Bavb/I/w9RpW6HCS0cPcbxmIpuhaPlDZOMQJI4T321LIJV2WprvFyO5HlmyoIYN1
6H9PHvrSyT9Jwm1lCwWX7exwtt3gfGo7vIGyQCmITO/fbQsoEylKaiLqMgHJquNw
pqhJYyE5JFoai1MQHlEbzxEZKoeacd3UsdjGKrvjvR8hfABxJ7DzBxxr9Qthyop2
w86CFrSjiPh1UGge0Ygb+ZX9l9ldbAZ3NNlxRnWilPWGeeis4Z27+fRnFEyiMIlg
UDqp40WzYBanxTjlI4/lxQ==
`protect END_PROTECTED
