`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM24QnDQz3DLw/FpXpGkmo51L6YgxT23dC+ybIOyAd8r
CGgPVXQDso3TCtX6MyPUE6E6r64XrI5zzZxdZXAKsW4LQH5KiUKeDB4zwXFl4Cw/
CyUjMagS1kRAC4VhuQEyT3X02/ct78oQC4Q/EjPAkji1AGETXSWKHX5FsLCnbnuR
V3rLz5beWzFO1zCGybefaSC05ddhixPXHMqgp3kE4NdZRAeMwQmlIUmI3qWC0chU
x+Vu//TuREuhz87fJzjS1DRU9YdylfpgpNCXTnBecszA1Z9pwYpWBxuR8Ua9u64P
Yl3U9puNANExogUz/VbomIs7znRKlzcS71CKXV8c35FQXKT8hZd6Rimdfplaaajn
lSbhP3GVg/gSCAxZ75JQV0KxEwpKa638hJV6eB1GD/u460JsINfGrPzhrCYTAWBS
b+coeG445goKsdAwxCW3Et+AkcCjbd6fiqo/pFa4u1Nj8a3CH3DT4EgbRwVRWcWH
`protect END_PROTECTED
