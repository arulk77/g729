`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGMg3HEf5LllOfmgvaR/R06ISW6ypNB1VSzC+vEtefNm
HoYFBRmRlpJmY7tAcrPVIhaNV/O08GPOWlPwPj0wTPoLLMx70vUaDlTAyWjMemkB
6yav0rihPR0zXNMN/Tu5wsnR7XX7W6c/bxa3qrUk1hCIrOJX35zkKyIoBF/tYhwh
dzxcDtspbYKMI34ZYoFRkwMyh1xK+fjANMarGOOw2mSuQv4/z0EIU1c1LkY/wZnc
`protect END_PROTECTED
