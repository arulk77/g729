`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu485pRCDMu+oLblJsRjSnxRCdU22P+dtwH/+4JJByjQab
LaMIyibHufiQoHSL0IMsDXIq9WEnTUfcMD205ifmrtwUeUuaUP0At3NtsO07ONbn
gFX3M32SY3rGhnHipVSUoNS7cVgrixBrcIQ4R6lKb29dQeG4W7toPeHQXiegmQ7f
ercy8nLZng8UGQ2aLcEi6Zon0WJ8CChmiTWCdIT0M/zy1EsXI7H+Rr+8LGiy8iuu
/mWIML4exZ5pdThFYUnfIoOsPtZ275/DeSsSFMd96n2Y7eX+lMHDZQj2LTgCj1tj
ZBgVPKXcYnSilTEMhJiV2A==
`protect END_PROTECTED
