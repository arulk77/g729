`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aYvxyxcMgDSLMzGZXQuEuL/BzjM+QizrYhAT+OEKta9g
3T+o6apipZZ2AfhAF/7bqtLi8oBdU1QVUy+USejl5JyME/bbIEmkVvHeMQT+69Al
GwU7OieNzOBkKXsvGYHSntjTYEc6HNIs95+KBn+BKi8SGUlP9hg4WHU5eILRHSig
gs9Ms4NyUUnrtmFozofXbGCUo8xhkQm7cN1xt4bmYm7UbQOpoLHcr2LmHETw13MI
Oi3AfCX3Gm7ozpKCXxWThaXJvbBt1P6AXzwyOi6jMBQlobl48ui3ar3/bYgFyNf7
MGIbxZ2dyvPGXZjVvVHmHXaAbJgy+zYKzrIJH2P5Dt9lkJcFnyBDHtwQ898X7wIR
`protect END_PROTECTED
