`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMj3utS2eQd2AEtVHYIDVDIkNVSDDAvKa8nUTFrqsIP9
3MXQdhbhsqKt0ZejmN+ZZBK9QCCOgKEQIdtgF8LcHObV6sAOpVqw4T3x1W13R/7x
t2fjPZxlmygnVRUOukbVO6M4H7yFfjX5G7FHbz4KW/aqbjLGks8VEtMo+/Be75DE
VuSZ89bPwNiGM3G1Gf1btw==
`protect END_PROTECTED
