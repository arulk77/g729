`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
RKs4q0QTLqrvYpr1SgXVaBy0aL9NSZn6QvhmVYhYsAP5T+y8R1CP4SPFvpTDynme
7WHlzlsWPa2sQ8b7VBxnfHJVmLBtF51fWJGDBlkaWlUEQqFU3oSbM00CqEtdP7Fp
pZmLCv8qQT4HbGVXyuWQnOMfqizmIj2Z1UWE+D/WAyIPC7yscL/RbXWpk44IZBfm
Q1pgxH5sYIPxIGmzdq0GDIn0M5QlQc4tamoU4Swq1pX3heoPEOKohA/3pC6WThal
sgjt7x+6WtrrOT3EqbIv5r7xaQu66u1sgNkbr2Zwl8W2EcSNav1+X2NhQbmho4cF
RN5vd+33jui9ez5QTGiAhUpAzLllUXoxrHnjmPsD/KOwXF6MZ9KL+Eo0U2oagdWh
SWrvfSO4Zh9OIW5cck9LUAg/c/psFJTULJUr4mkzPuk7h9y/sPckzMlGlCqoJUTg
RUY/ljxwtwxKVIeykRXd29/tfHmMNX3tGp3hPfJ+nyzHCpjG0hJSbB9sYCc27klE
gL7cwf/MJ5BqVV5c1LyKJpZaUo/7Ex5olZVoDG/cjORDaoU5nruMKNLhuH8HKb5i
Y5xSUhmLT7aGntJzc4biz+bqsZeVGtUUfkXcu26dVxBsqYZboy62qI5NW/aHv3zW
h/y17RiefEEo739IjuJm8cfIvwHKpHWZc/vor04ITsQh0SzqbXllarTJpOSse7/D
EXmMzMr0KIsSFPxMYZ1TvDn+uWdQVCE0u4FeyVt5QLZJZdlQR6b4fPrN+Je0iX2g
DDHe0XLbPUOT0f/F1V0d1OgEQCW9ocM1a4o0cTB+1zP5qRjVYPTetQDoMwUyeNDI
`protect END_PROTECTED
