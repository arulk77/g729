`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKXmAqMTc5EsqjhqmoAttJCLFieYy4ve5IHhCc1TgHK4
UgwiRc8aIN/il/vvdizM01tAo/VjrbCqG9NA+4f/v92Sa1LdRKSKDs91+GiQEU5h
XJsAr00jsj8xh9aB1qNta6T9En1s8MOaEJ/IamdhrXQxlDdMZq+FmgU8y6GmRJAz
n/eQzFDLOGYWCBZTyZVhvA==
`protect END_PROTECTED
