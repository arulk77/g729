`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOAMynqc9XBxy2IA6RlShdwo3Vcs77xZJmwlGZnBgF0E
RZehKbOC8W9RLMQyvBpXE8AWi8Ul5XKs66TElVvfzT0Ig+ykpTp+tFn3nvRRGIFX
6cYrl+PXoRA9Op5nib9SVKCvxkZVh8OJH2mXjZnpmkq59umaOVt1YLOovGCxq5gc
L2Ip78oRo9HAro+JHaWvokHRcZlKdJnAVnW/Y0LmSqBmkB0LhotPKi38zfCeABJN
epmv/55/L2I34eaCcX2z0gSI2bINZJieMMMtLCER5IuPWD4W3DyRJNX1z25mHL+n
mkhdq2WrM45deqEu1kCvKYbtobnKEnm2h2gzxKLhl8uyxjRipdkcFhwULE8twA9+
A7SQTL9dPVDsHMRUvStgWM+w4Sop+6xWFEthwy8uks+PhZb+T5kH4glAwxEtKVpw
vxDtR0UNu0VvrsDg2bDMxsNXqRg+itCpMy1c2eJ7m5ErgTbAfA472sO48KLGEmYx
UeEsuGb0wHUSN4qK7YOPsGmDmHiqcTJ2Gig+JAi4wTzfi4WV6nePzbVVxF7U+hkB
NKAJO1PoCHbC5fvfT2QHNvWmHtCDsU0fKeSYRoVvltYdb3WffR+hPZY+t6JAZTO6
WLlYB6aepTZ95cBpUrG3RA2stET2n0FjcSCmPG2xL1ozYAYMwP86veGumpxQx0aP
4sigro5qoTNq8tNEL9r0ay21b8oWH6fhSKq0p2VF9VwLazWYTZbmRUrW5yiyJuHT
b0oQNPa0ToLeEkxqiSxa/0UKX4to418Zft8VaYiq2/PnL5HkSzcY3laSAs8fdMiy
QXT2trbnVmlQX5HruSz4VGVJmtIy8ompxPvWVVhIREYeYkxNcsbXXHYwrth7Vzxz
FMyRB/e41AzhXMC8dOXlbDYDvH39DTOTfUi4Iul7SSVvfAcRWx7i/W6XyorQ2qGx
5JOS+pLk2Wv22D61WBK1jvFZegrZegAmX+4lM42jNELwL5Q+sgfQRqF+R+lKkBGn
p+wIrJpabvam6iXX9cp1k2Dq50E3kv9Jqk+K3YVsjRMcvAfHq0UuSMFEKSQX0uXi
WvYrvscKzYPJgLwbsUHmmOKmA+mk+d62NzDS2XtUtIht1TYn/zEGeFp0/JkiMT77
q/m8KhJct1Ij1KDuzBGJEbVnxcSTDnUxBLnnTHk9OJcj+UVYPwGPREn1cZ6ziWdp
bxcLWqwXbZtQnsbEJlbkbBGHHWG1y4LNLWC7yI/uDJVOZe3aMkYxN1oxtjQ9dBgU
`protect END_PROTECTED
