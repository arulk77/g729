`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAZS+TP57q2bUcaXdqTaOIkVvZf28QnP6vp58OcBFx75q
Wvm7xb2b8QhtG+/KWP2EGervf23BaKQGUSfa8buWZqO5XxrKgVMR+VVpR5riRq65
PZtobhY0IjKDI382UIqgRb3pvv8qnGSOUhbKZJBbKkxBljPlXqgCBMYfey+0vr6w
Ln+skFVZHNpP/JLDxKgKG5uNOL5Ejx9/jvh1N3MUzgxX5MUOEe4OigHdz88GzQNK
ZthxFL6vuWyVtUbNJF6HIY22JmOJGnjE8igMJ1OdLDUvI42Lg2Vs+Ayiih5zKBFw
DzUGI4u60zpz+6jE6hqqcyKVQ1YAW3OJhe/7g0rj3i82je5A5W1j3sECC6wMvAy+
E+bVnbULRkXwusswKx0htN1huN+nuyZxIAcW5mNcwhjuCcgTRAxNQ1doiGxYYUId
r/LTRBKvM0GgF93a2MUb1PhOjy8Pc6KvDHfiopwfJK2l30rbGbz/5Zc6v/LE2bgH
KGOFG7btF1sn8tjHWOCGw4WURY1X07JVlxSArHOLE6DvGfIgxNejGdQFMGTD6bkQ
ZuCc1ALYUX9C8IE/baWafNrz96utjbEe5Gkva51WRG6hsjwcMGlNZY3LfCU6nAh+
Gsc4A8d6OfGLMtvcp1cc8oAw7pLN0oak9aeRZvP3cxdbx1HCFetDkVRL17ILwFm1
MItgH8mgftmGOZFZJ5ofgRHlmA9U6pZkiApm8f6c0OzMpaOLPc+uZmyMnIaMe0c0
85lYhWuTkZ74C00SJfrh1GVXd3XYptT0AeP7ldLZZN78oohO76zlhDQCMrLvGDBR
H452PaXBuV/SI2AP12231vA5z+fVQKw9uEJ+T3iZAD3tlhI/B1A/SdJXBKYRSsow
wG1WhQpHsCvm7nCybmozVwDY1ROGp4ApsfHWlADrmgK8IrAqbeJ6+LH6q8lQqPBB
dKG8Ji5fqBwgx+30D1l5IfVIKHkyS/jmI6fYSOCUxNQfuu+fNj3/ASfFEV8RPY1I
RMZpwdx6gCl4fdM5NLrBUaXl1ma/B6btD2DRufeiE8be5pFm34BCHNtVcHtk2w3r
E0KIs0k59lxGvUI+RjJY0De0PeolHE723UrNu1Fd6ic=
`protect END_PROTECTED
