library verilog;
use verilog.vl_types.all;
entity SRLC16E is
    generic(
        INIT            : integer := 0
    );
    port(
        Q               : out    vl_logic;
        Q15             : out    vl_logic;
        A0              : in     vl_logic;
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        A3              : in     vl_logic;
        CE              : in     vl_logic;
        CLK             : in     vl_logic;
        D               : in     vl_logic
    );
end SRLC16E;
