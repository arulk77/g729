`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C5SlZ5FDrdxmyF88qeYJ43/Ai7BVUfWSYUkNUT1wWBFi
OrsCxlA7d3oLi1VGJeQDhcqHXOps8lAMRzgkrA77R5LihzhbT+ndmqryStjfu8rz
bGxG2qPS9s0QnTPiE59hJhNei/MpnZZIUy5pm+alojYQMAKxGJV/XiPmaG0bV+7U
46LWMkZ9t2Ji+YPzpWjKln0Wy1ekZdkc2AUEke4/5Kz2xyg7NC9lNb5Mac+yB50x
Tv93dFSuXtDlIUicN4cKjtE8Lao3TQrsfNpkiFlsWoCTnXGqPYWw9Md2BejI1BH3
s+KshpHJF+aSAljAXSZCVYNA+qwQQSt5XCB0J5Rmrlu4Nt84icxVs5wayMDGpA5x
iL9yPHjYCuMV4cpvqAysf2PHjP7Y1ZFfYigk5JCRBodqE9dm1nki61MVEzosYtOw
rWbew/xukt985atwtDCwoaAJfHK+2C01EABk/2x1kEEy6MzP4jc5Ji/EdCv3ULZi
7muMiDfSJD9OlyavP5p4NAKKDpnjmSPN718iBdSKF1+tC8V3AJrTak1bNXTEJ6zq
AW2qqZGmXEArA5PqrwQ3gfdDVLlifnkg/zuRQHXP00GU7j1CRsiimVvPcKMaeaRG
/3nxoH8YkfG07iPQHD7vLb4+pFKRWsNE64GH78zoJBpw1+enrWAYPMudd5arWcSU
wHdu7sAR+O6bSYOHQL3IWhxkgAE/TtjezLhyZIspWom6vUGqo664mIw7FzOnsuil
k/EUmV4x8p7UiOvFK7MWt1BS1asH+fQEOKwyYuzya4FDpXpfeeaAB2c2Nw/QrfZb
ADsbouUFImMuyz9VWGYSn2ZHEJi5Yi7HAnQSRTG1j1UJ7kGM+lRT0+wtS+m3EX1q
X6J0AFAVJPl/nCFCnXUccvcImi5qd8WqfURzkuUTftAnNQjYxMaMrYkU1osKxKIG
E/x87WQ1PxPPVUq2zKSV01ygRsCU3FvUmh4gWdANeht6/DGBHzdG8aFzHjoRF34Q
NMiMUd/SMGykg7xCV6r9ncVpJ6Vxn69LegwRhp2bN+I2L2cVgLx4XBfg23dsUxAB
x4vIFzhsFN3KJ/KX2XVAuhU5aG8JK+9pMMaWtp1Irlo1nMD3H1pUmH2dEUl3PZY8
GNcAowjZ/3/xjWYbHGbdh5Ane7b4WOc9E9ibTchluCn6n5aW9tcdAX/iUAA8lrY0
a+UGLZllrZcscfLLayYeeUN0Or0tszQ5JJ/JJnbwj4AjfQ9XKUxyKwQVRjCVhA8O
6bK0fFkINz4djOStjbEPO93vBEnRcSACTWC5YlMW6rHo6o3APRFqm/sUdOxGIjZm
2UcmcqSzgZRQ2FvhjynxBOY5Zpo1Kj88IoKviT6ci6dfE3QQosHn8WfaVCuvWJMw
mmQd2+osVgYuJQBZE4iHR5gnnCj5sHFmuk1slNI/7c7DYZLiiAkLtc/OhAqDCcVu
B1VEeNq+6CEJSdhx520T9t3ie+0V2ej6WQ3pBMQqKXlHPzx+rG/2n7zwDFK2nDk7
Nc1d5BebShHvZxSVbMRL9cDNMqffwjjuAtk6w+OorMccAi7hfvPytb2f38LviGjA
kRcsvnOihSK9QPggeKyPcG2RfJh63zcSZrTofiVH6M1Iaw5ImnU5SaSfS9o2WAUL
Usxgufc9rtkmNzguHC8DNeQ22HBM7dZGoQzulLRJvCnAo62B0Id1Ehac1YT312BI
E6gRiFGPj55fU6bvOfbE2Zc1dlews/wpDHlYKjXQ/NE53XJ8bNrtqoAUlby4Q2we
0fk1wky/KDufM5JYBNRkLf3PI8BPltUB/BJUVavr5SoOgm61+Sewlx/SHS3/JwmF
mqPcdrPquP3sqn3fkVaUtM7dUIZp9xTCc/PbKMB3GWjC3cmh8bV8c08HVn58uR+B
HSR+2A1QQ/GS9nZ3ujkPIycTxPmEaM+yN8M1FMEOKMOCIXZxuWYjYPgTBGU45XVV
mFkbJRJTJ7wKZKWB5c8JruffsZLHhV7xUpDkHgDGdIP1ciQ5Huvxg8jzY+r1QL7K
iR9qRTNtEo+wCdrzlIO4iwoOvyBTpAevVEIxX1N+1lJTOcxuxEVLoFaaZJZpnkQ6
jvpi+U5CoAVqWbtL7tNo93O7hxuszO5oB4Rd8nD+LKRVRArqj8phzelnV8fpQ1xP
7Btpj8xR8gFdf0ITdUj+7Q25yB9C/bGKFHybI5nyzjW11glesXgZnxaOPmsdqt2J
H36x+IX3RVVLR67I/JKmZrcfXqgQxPHU5oLW4N3sojF8jbL1xTf+edd/hXn/D5/x
C3QhjmYo+aKiMcxcgLZpRcRenNApoRS+km1+VYnJPc6/R0mZX61ZDvFWhc/MnclI
dx/VAdqbKDD0iIDHeopcILMifZ5/nLYHkInl8mbRpV1JWH7bILrCjiC9w0JofQZV
421H+YK+DDWyM5++UVJgHIVnN6lR1v+Cbnpea8+X+fADG+Y1dPAZqEE4HMBIVHXZ
3uE7cdTcAVPIQ0t7VGNtzyD87wOaPDN0ggNm4T/3UkFqNH785Z8C/FrVlbC+jW5+
2uy9D0SlFNEtasP7zs02N7KFNG8YU0QnvzHnjN0/s8Z3BySeCcyOXBvpVgKvFomJ
2X8kbGcg+I4Z3D4Dcb409mZWjiee7j2uMNsDM+40mVhezNq6YnrKKEIRr1bg8aSX
9/W3tjF5QmK3avnq578aO3LDK+di/W6vjJfW+Ezq5oLiHxDfUiUUzWKFdtr4kW9O
8YRitG+v4lgwkQeTeTUmobUgWfZ+bAz6+a7B7UOuHSdcANT9cApbK+9k7M3i/Cp7
bsIe8iPpfKcStG5eftaQFrUdZD1mxc18TCNTeGJasQH3DEG1/NdyzF1dq0VoLgr+
CK59DCCRsDhaLOD8UMwuaAwC/UlnL1mHSPBjTJlwdyiEfqWIqvqDkTFpIVv0o0+G
VTq6lpHq3TxUYNklTswa4/ipBys2IYfi3swJK+BtYkh3WW5kBvw9j+AuRU50l5Hp
oANAVLRf7IQ2PbWCpe5TpBFL/0wQqqIIxBLR+lIn0vtSq87Aa5S/s3fzEhsUlLG6
x0p94PaeMcQJ9QdtdYoSMP/emBwZv9es2OuH1vd8QMBw6UI3WSXVZoHh5Koi9FDn
BQ3R6DW0F+1Ajl0nFusht6piv3xy8a/EX+UKFDFbUp6MBBULe/1merbpV9HWVpSu
l8lcrwM7SsaG0OfYL7w1zQ+yGwBNUcniaQJPBCSgNIOmhfMsxVshQd9jjtBUqN0s
H7PUdcZamQbemaeOquwmFCFG3urb52PmxaTMVN8juoqQqlBl1jDmO1JI2GQ2Y9Rx
1o5vww4kGziyeqTCMVv/W0F0oswZTyu3PFscW5vAN/FKrKKzamHg4xJFPKu+ucAf
Br9NCGGwd88FkEkbjOGkEIy4fE231CRxkdrh0yeQjpKOgA74aYvBSzDVTj8R2dMa
7kEpd4kq4rahvaYUXxZhJM+ZQxD7GLZL5SVPRQnLlXHIMqmxLRp2XAXCOF/hh7hQ
+8wPQ6nZ9CY0Jy4Y9oOknmvRoGVcYalju0onzWlfuBF6qgIqHr+zVYHcG37hjiEX
gHCCdOH+SGxL2qxGkTgWgGW0zRrb4NSjYRdiTpXcZVhLlttdYZ89BT50n+5WVr+e
pfBOTr5yDEfO46IF8z7f3zldKZMugNaM1TUZu1CBqq4=
`protect END_PROTECTED
