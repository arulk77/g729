`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4jUYkdt5VjR8oFbu7ZiLklQMIyUW7D9uW943q3sw6bx6yoCSQwO/JCw53rQ8QW5s
lk2FiGHi0V/OhaQ+c7Oou2Ma3cFKNQKK0dz1RRtI27Srasstitzcy/4znGtr+GFU
AnzjD1pOLkKsMy1HPUDKlhAfZCkq8PUApbRfiaxE0iAJE+aOhcOXk0j2kDATd1u6
pFD9iPylRxeok0QSRiYCpYONZXBnFRCsY2KG4bXlIcxZo48hq+7XgmzlRBhs90B2
O4gcOaqB/kDQpSQ7ASTzfmL9HlEbE06GfXvlHMqSW46BI86Q1lcmB1hjv0bdFHhp
`protect END_PROTECTED
