`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDr1OIpqPTbcW8ReU2Bxg7A0SJsysOtdd3JmJZ6YOJZL
OwFI38mILWybdX2bVgzNuaIHWVk8YPW3q8Evhf7a7ie+6jZdNOzZn34v4+JQ1Ldg
7a9TI++2FMxqv98tGqdiNZ14frOSedkRosWb57GkCQZCwawyInxjcMI5m/9YQXOB
aon4gxHdAmYE92xUAfoZlsx0SGVPv4gl4UWXRHWrLasjPuzVKHEaOp5Y/M44oqsf
6aU5UCuVvpRP9XfQi9mPpb2AU4OqZUL0A/r7xiKklbHztcqMR/ThkeNQ7fO+GAPu
9StyMkdiwwAg0NFztKZz0QlhnGyvpx9mRn1letQJb0g=
`protect END_PROTECTED
