`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveE3Fgf3WU5149jWS/s6CPop/PJ/Xmn1tyGd2bSYXX/CW
ry7onN3Y/2hAWrbjaoNxbDPWIItwQQRwcsCxspB1KvrSveO/s5A4uSYOME9HcNZz
vWBzF9dWq8rstnE2UchveQZeEB2eCq8KiygTjThv2ABTc4tuC2WB5t12CicDPEqs
nhzGugvG9KfEtqLj/+HKrMnMTyrOuNuZ+HR6lhuTa4MJin//vTJHV90Z5KDoFGtO
`protect END_PROTECTED
