`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45qYDeOPRLYhr5Xm82qs/J+pVaxfl3RzRHfOO+HjA06R
AJAXMKcS8Mzhf7n4uuorFumk0PdoA0NO6TK49+Zi/ZTrihZDb7vxwgrRF9xI1on+
yfQvTDnrzbJAzkAVYP450ZDyofTWYEQ7QUg7om2iOx3j5x7T4F5w03lU7aKfkmfs
HWGNJ770nTW6b6ivQ3Qu8ohjhXo94liVHNhBeoJEhqD4TaxtOlgIyxyF0HBWcXni
RkX/AMNLPhw+nn0USRlgr/OrspsoJXeOq8K7s4W3lH3p8Q3t6AzMqWmd4tzl+BCn
G5esdwWl5NOs/xxFUyNF9IheK9YELRv2IcKhEMAQs5kgorH0v34oHKhbI2XmKpLa
Z/Yb2B2j8rVmnqmvXmnzGw==
`protect END_PROTECTED
