`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44s6leCuo/AoxlkkSl8qOdLJZ0n+edfiS2rjq5OW4UCU
nsEFppqJai76/0f8OWhdpL6jnJNdd6pzAoUvJx6mdRFaJdXft0V2i0ZWojbD4GMf
Dfw39D88K2V1mK/+zGN1JhjHvyp5iTsFedruVRN1Pm2upo8ftt4wM2HrSutibNaB
Uu5f04BvZMrzf9G0qoImO1lCDwU0YH0Q9AyNVSRtaFdH2JoygSAJiI+TRNJu8fAg
ZuwsZfuBIvXNz68SraqWdEwgsVapS5ZDVCZYyNjra05DK5x56WDytI2l7WL+k1p2
gTtEDj/CUhNxD2MAAOs6v8uufSe821c8apxS36H5p5ixz7ISMo+iK6SPkb8eZe2+
FrokLWzw1Efb7KKErlWYPQ==
`protect END_PROTECTED
