`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN6B99LN/l1UrXqkbNu7Pxrm6vYDeCe4ETq4WJfoqERd
Ke+F17Dblh43OINZgpWptpTYNY8HiV5B+ZmYPt1xNuA4msv59xJUI4Gj7h7gIxo+
pPxNW0h7iiNj1xRet/zUPflUTMf/0798NdxxCk5rKr6jd0gAOlmlKZFk0a8AaHpz
HuZ6ukHcul8QbVTA9YEDudUU4qh6sDfAf2+UlqdASdi506Zpd2chp1X35bU/5g6e
SX2kEsOpaz7t/+dURZcjafUfcuz9GIvUh1msTOjknxZgVBIOcFXVtAW5Y9pHx/3r
rVH5AeV5yycT38Rfi6tnZwek+QI3ExGq4R4os93dTLnekcRfiEiEfC2b905A3eip
`protect END_PROTECTED
