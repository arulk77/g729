`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Prgb+lMGK4ankHVaNnLDq07BJ3X+auzZeNaxnfG8sLUiGY2cekliFuUaOy3JfqJD
CuRlCP5o26IHlqZ9FIjauwCJ0lxT97Rnr29NqabOrAE0wl2uVIaJ7GEF3cvXYUmG
HqTYHCJr2fOcApW9DkEKdIwWLfAHc5ZyAPRBvI3TCsnteOGGw+b3BcuetKsAMJ4O
Tw4DWmNJibSCS5+LJaq+jF1yQ+BYUx4l0XXZcLMVyEg8TXpREsX0YyqYCsyFpG5g
up1gx/SntYo4U0NjIAnzlcdqeCcsXTYLuLt64X3J39c9V0niZN5+GsnPCxswVXiD
`protect END_PROTECTED
