`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL1VN9VvjHc/nHVuRxeiMo6KwtywWnj3030ji4VVWLu9
7jRTg2LLajnGGGZKC2Ivr0GOCgbduqUWs8H2VQkIR4kxFz54WofzHYhVpodHv4FY
/qQvYOkVFRgg6sWJ+t9jv0OHmDTCFpDmt4MiiUB3oEkSe7rpjorqMIjTttsTRO19
PpAhAb2hP7zlMx0th75thKXcAf/nS3bN4am5YkXJvNyYFsHeX7w8yiZaAE0eNfIw
3IRg4HY3tFXyG70gXwk+H/svFADuLj6vPOS878OQ74efLsmwfGr0WCYm83oyDoTA
bVWnrC3PNtx9+sayzzKRi/RWb6cC6fIMVM2E2C6bPEp8BrtoHxSf1hQB40LIC+Nb
C4ZoW3z+NeqMG5fVlDM424PQ+hSNgNaLSQRAatuS6P69BElyCkY1UcZcwceNkOFX
d1V5JHHeK9+4W7nlER4KheVsBicQf88ZTL40F2laYkVY2oYmGO9YsQG5d8VUeJTz
BD9D/oFYOOtqkTlgPrg8GAWZ0WA3ceDuwabEhdBiWeKxQlFayPwoi80R0G0xgGOO
POHYNhiS3zEclx3kkSC97g==
`protect END_PROTECTED
