`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C+WUdoY2Le3ZKDLM0zruTIn7/JY89z0I+JFHT044aNni
ZkljMu4vU/oTEQWAvhSRvAiJYtAF0vc1QGZEsKKZQMsTTzt9q6Kc3uGg24eo9MUT
FoZtwYadyCNu0pipYNhIo9K93arYAhk//p5VZHhY/TPSVuxuy2Q0I82Y+1CB9oax
vBIcOzgOmeq1bQv7MtsBC6BS9g0TudQL0dayRA/qpOz8rjbd/j0bWYYDQ5IBHsvr
YN7r4lvLdTuPSm31Vxydsw==
`protect END_PROTECTED
