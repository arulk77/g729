`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
nmLzVXiFEHkU7+pQ4s9IYsob0BSukRltyNe1sYm9528QHfAHjpMDGXpZdi6PLxVe
Odg3fO3bJKkQn+cn5QomRjmn4XUOXUuSqJCumXNeohQIqMmRoDLMaHEotZJvTnme
2ieAhwkZr1nDUkUZkviTlfrmIHncZdgBAcaVrfobhKnLARooHsDg2+5xOdQU1+Oa
ScYCoUSgdK3kcB/PWIH0RcHj5lofo5yFrCpLy6HS2sY7I8QR3H0Ir8yvPJ2NEDWw
PM6W8Ny+P4vjsOX6cJ2sMhBuSiDsFj9Sad6rSJjuk5uYvEsYj62AcYVEQH3HHn9z
xVxeXMdc9ufOqD7anL+/aBzbo+byVjW9tZhn4D0oVFvMP6hkoCAzcewZibtZPEzd
Nc0JZsP1TL7J7VURFrcipf2Hw469eYfNIsiCyt1dPzJ7Tzamm/XqR1SHV2AsozH5
7yVKxI32h3cpddh5XiFHUvBS5hFk7RTDUwmuY1JA0JDb6nVODbBCW8/bU1+lnXZd
G+VJ5h/GMx8JUv7LQRzGgF1HdPl6kTA1p2G8K+q+Cy2nMy/mRS+iTMTO4P4MRnBy
cU94FX8Oolly2modi5w7aCqdMo7bHsCoUXjuJkTis8y1FQUr1HuNfYw2i9LFjJET
i38tzjSKf6sGEjBDycTSkixIKy8xoUM6CmOA3yJIytHgIg0uhmiRShzXU9RLk6Dx
3ObTaKvEcxnmbwhEGdqyphcID0foSiVd4p0YYF7/5lv9xf89RoTAZjQFmk66tii5
uN8sUSS/Iq4JZlTxcwMpnduGey89pBu/byTeHMsbjPi7CTDajlUSL7goasoWV6bs
3svI6jYlEFMN4Cb10FYfrv0z2ku5VaxppMJDrIGI9Zybvako92R5AW3qLrbBy5+E
gBxRovXoTYMzjE9dtUNI1dG61IIIxR1eODXsj1qO0av0Sn7oEzs17Wgl7xjVHwUe
ULOeOp9cNKqXzMxP869o04MGXs9CPF0elExa20P0IjHNr8zvtWa1pk0O/D8OtIGf
ezeGJusKXHJhDniGgk1oYmWvURS42uUDMupCgHIeGnXlPJHN7g9tQk0pgZSSYQqS
XXX1qEI6lrbsyOekRddhGL4u/vqED9umPHaijCqn0MJ9CJ0O4aHyg/+gmVft7tD3
8U8jT8006Siwe3QVIkIOuUr8TAnKfFA+XD9s6aDhIc9cm4smwJwSeoFLQGzUYmOm
L9a59rG91JNsNwVmDuTbIpPCAfKwrOe5TlwPMmK7pSVgHgc3DlwcdXTv3BbUL3RF
ael/PzWzGCBtWCFKgh5a3hUIxid+Dm2x5ogtexPIm0xp60FgxW0dv2+Lhp9U6B+m
aqQmpuNj1CvzDEWs70jEe5G9BxS8M8u5nO73DpeAb2Ha/foVULPYY26VTN7Z1u8L
+fG9HRpXz9tqvT1kkHNAs4mFEvLLwAGLFgiRdbxO90tjSEHBM+eDFzhWHwMnJnjt
ZDG+Yyn2KHRX8JsarPb3UZjYjZY7AxzBu8798D+BdQlOdMjgEi3npDL3yAkDcCFk
Ehve0P22ch/3l+21wbmo/5IcBxqK9kO387M1wYnMhm6/Q57nwXXgNFXf7xVWCaM6
kVKmjVRKG+DPvTwRrJ9Hpa96aLfdOJwjTSJmSPw7mscZNXy/L2FLNPUJJLSn7kZB
Ej9utjAtvbdO9oKw7D5tg8CQi3afU5JS3tx3ehWJOSYFohg5GvlqLqF9c3UYkJMM
nrv5XUATkAxu772yL7WG5/EmpTvV3YqcTGcrE7nfTSuip7vdeBn56xWvS32dB5ZF
KqWdhfxN2JL9mgS34G/zqFyV3LV39DyEsM737qMEWJZfo/ZHpOakoHSNYJT4y5iX
xcitZepKmY8nv6m0Y6/cjDSw9y7gBue5aNSyY9niJdbTdqpmysvqLU9BrOyCvqtT
QJhjoEE4L1gwtviLw5TZRvxUeu7WaGnprbhJrYLKa9AxKqX1pRTm6vQOiUMtoQnH
uWYMb1uWGMSLRDbgyLIqywjE/HRSpe1218BiULnNQpGB0UCa6fq8d1Ak9rJnSAJk
32fENFxTHe3tZr0avuHDH0cgfE8jUlOALi9YdmP5qAMoCOUv4R5LC3yMy9dGJD9C
PGjJl8k2H0yjiPRCVPxPPSsE1ngCoyf91hR9nir0Gj4rlgi13yL/Ik1bjv6p2JL6
nfhoxNCHVMhu1Ivkik/TwlpTvOmLM7AhrFbFZf72YuhXxQomgb+WgrDq2KY76qWH
xRyQVrAl41103nx5yPZ3fX+9u8x6mIf6K/EVlwv8TQrj0B+AhWEMYGX/IXmXTSIa
7OOdRdbtESl2O3rrQGfo1ESybr1Jz9elZJcl+5b3H3fwrGzOWBQfqRmCwY9255Mt
/ooSKd8dH5IC0GP8K/Q9SbCJUyNbruQaiUJVxa1IiPO5CWKLxc3Y+kBxbE8UslbP
5B/6w6GNPm2rJsBTtx47yOX7rShAEIgyG2DjKvA4o9ASEWW9e2OPQMBuvY/MUEP2
QMqwQRaeNEhMJVTOYPhK6OZO3A3dI8ZIZHaB9M4E/q9nnc3fTStY0U+HvmRh2rOa
6DjzFvVgdN4rd87UqjOFAkt/1UXDpyh2BxGPDdfnVeHsKSdy5hsetKCYTcsnM0m6
eMFzdh1EQ0HSlqCS0xzC03FKvbDzaeAkP5kM3U1021qgUrUWK39TQiwzO+7zGaxU
j+GXdqFwb593xSUYJqRryF8SiT1QZEr4MCn3dUJ1y8FIXsWtin0bpTXwrgdkoL6/
1qD4XSAAfGduGJDT/BsBmSvUBIzk7mBynGK+BQ6tpgPw2LUSHVgIpWfUFcuL/7+p
9IpCO50PlBQKF2foiawykNJZ0gFKCEqeNSgZjDhTWoNfWMX3ObpUMx7aYOQZhJ5a
WhV3wrtazi0lObKivtHCLlz2fZb0r0AWnYs5nq1kuatQF44HxgXFj8MASq1cRIwi
ascJ7Ecir4QF8+14l4mVDEj1i2hUi//WyGaSL/wjsg9cofICpybSbEjoYuleS5Di
hbo0YqTGA5UoXUBKsRAhsxThhX8PkNJBTyzkZKp64OaOaGw43Yi3ndiSTopHtO3L
rGRsMPjA+KJLRG1Yrb6R299cuFYh9wLYhkVNlApKGBiEKoPtEgpggj+kzynY59Ua
vJisBJb10OSUu6lSPTtYG6lAT0UD2odXnDHEsR5KDar9ONyPH/7/LNmkBf/b8Jor
dP7ZzQCDP5wunDYGMll/uiC2OX81N+D/ukxcUH6n6CwJhoJqQXOXddCz++e3sgjW
zrqGfeGgkUcVt10wQiTbgLIvrWxr5WYQHQcJoMLRAY+tLSqspbotDabalUcbTrbQ
Y8IwS9FUJg+wcxTCT89UUA+9Y/MtHl0u/BP7Hf59ho4mhafH5PQh9j1mS1386AyV
lgl0h819pgNpcCF4nNuEOXfwJS5KAugIYUTGRDDzfBDza2t4nqiHXngDSN6Ahvyl
OFNjNkRK4vojdePw29ZtYZo7/amjT/P7NqzPfzVG1EqtOnIn9DgFdnoQy5n9sRm/
3/UeZzLfkCntVGbJySz4bLDrV2G3VyQuvrYyEVA0nAzyQJxoe1pWJUm1NBzk4AlK
NOdPKl550h3oe4q60HLsG9GB6tzM22yadeF58KqHIrB4h1zu60JzxHVDDHYqH8W0
YpFgEKFBw2pysJc8PTqLEKWAMtUD48XzcCdIJHfdOBk=
`protect END_PROTECTED
