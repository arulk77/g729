`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43HvbUWFVgD4FLtoSaIIzJ26CkXah09rZ/ipzLmu4V7+
MUhqN9/665a0cvjyHoeOBGtdo+xed64Ct1KS0l8/KPuOvB0z1Vgpa89A5gfA6SkI
RAQu6794OKKs8FJ2oku/ILnsYUoJIusGKY/Em1Q5rHAeko/2gPNMeAwibjFYoD8Q
KzOGxM2zgOTMGe1JBy8kgHxLgoyJy2mKMCXxMYQh0kI=
`protect END_PROTECTED
