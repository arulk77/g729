`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
w3h/3Wbq34V9zEHTdWn/pOsruqFRCVt5qh5sheQl/anXMnXtwaBuFZw80nhlS+pz
cdBUsnaX8ZWGPdSEYHeoJaPBReHeywzfAnY4InSc9bxYCq4qndMkG+Fbemgj2nyr
UQPf6YX3lUzee6RiBVIAB9JnFPiTm+Od16/dgkZA2xhfhpmsmBIot6snlk3LKXH0
Iz3w4br+BqkVSoGyPtmcJ4acTEHDMQsDKQsAr+ESpw6rGkVng+QrXXOBn8a3ZNlR
ETOhSumvzUISuozJBrNZetduBallV5wW2H1+VR0d3zKq9OJqthOQ2ARteHYinZww
WnL4AbnbyAp6t0z3C2Q1T7b/NBdq8D2qVrmlxbJje3JEGKX9BVXEp6WP77HR5qzt
2HaLMxKVvglwvgMrGpvSI/YpktOcJsVzZ9TlotATr7A=
`protect END_PROTECTED
