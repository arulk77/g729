`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43aeD1gWWxRW7AiSWfAmGWcfXNasfFxvM/eaAB7MXgQ8
uWYYxfSl8n40KVaVFZ8MbNuwF8ltqx39eYds8WzUm1SGi9juJLhE+uER2zJ+ddsW
qq1139ap0mfZWPxwSeIbFP4wCaYfyXgXjuhCwigx/HECT6iPrVfls61dsgTp/6fu
PZr2AUmfa7avWL6eTjCnCuuCyuJgofnz0CFmt93OWg+nLxxptH0SAC3eAkuWECws
Txl8027GP4/uITzb02LmqRJmtbntrMMe08H8WxmMoSE=
`protect END_PROTECTED
