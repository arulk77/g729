`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNyD5TdMXYoz81DMB+0xdemyr7CjPhAGkfFuKd1pbQlN0
ts02yeMHfKVwGeWVbvkg5o8E59ooDdl7kLm3fRREgwsaPYMCoFIz42iD71iFPFMo
bq/rlE/vmGXJD1oqa4KAeKNtiK6dsZbQ4ithvPbkcEHRCSZqTWh8KL6TFvf52S6E
zhUHvTO/tARKWWvF0b9FJx5438VKafHCIVHTX3x52mMNiP0AO8Cvph8Q7/3nKwU2
/Z6s6YBp2rY8GwzeYuXZpe2fkyalP70phS4Ec6s7H2D0MwiEKjMr69HQQQK/y1z+
W/GMEnlNrFQeAel0ts733U7B4DZyNHeQ0tuLqxXSka3sHI2uMB89FVVYJ4a4NW7W
/uvgyHNBMcZZj7FakwiUU6BA48vQqrR2qG/D9KG4l5Qt48Qp5FnavFTCHa7ae6g/
0jczvi22O/Xz5E8ZPs11O7cRrU8E1Ch2FcojzBBClcGsQoDd+adou/BoJ2izmatY
PxQt6uQPL3UZUu3Y1q07ldnh9w2D4V5XniQJTuyvtl7rSFHIpqIUvebYqfhVLCbR
v2Se8thKvEmhL7YUpkwmFWfV7u/xqJZD/78ZF3vYN3VEVqAWxXY82nBqSV/kC5Ww
kvr0PvaXyI6f1glM4u2+hHKcGLjc9taSLblpjRD5ueBoSC7CvVK62PeqosoxShl4
QrDZYeF0pc+pmSMvZcl8GtQWeP8cUV1i9JTinctPWPvAlLJoMy8RhSEhV7WwfXC/
LReX2UBa+1JZZnU6+P92rh0+CDsu4yIrht0eCnC3UxM2+uoKq+gLiFbwEZtaVrMA
Dv1COvuhNS5oGYUuyKjnTWfsqk+Y/E+b33hCfw/dwI+HOy9wlBJaD6xKUopdtN/t
MktfYleE+OACmeuWUewiYslxMn4fSL4MGbJ7ynBjDNRDvwJmdorH10DMdPhlEMIU
YZJMUK3raRmUvNrRVh8ud8u+zEzm+/blzZLwLHwcYXrZ1JDZkxvN9UTsWu66CTsM
44rXeYrEuJYY4wEVpXf9H2jAVVjFCz75kWdXsVPyjgAbxd4szwd2db9xbebv5yxA
Fv6CSNylS7Pmym318UffTz57J3Hpe5ikTgvHDYkTXLeHGswqAjriGlPpxDD+jnVB
mp3isZufvtwhWyIBKTaJl3cvC2bpM+hJgzOXl1E4kvS7xqOGNhpTqw1GHLR4hLOV
yxCB6AaOTMU2xcHY1GjHwQXVD8clCxJ1KAg2V2n0iAaVaW4g5H0ha0nir0hESrun
nKDVFwyqB/FAMY5qMk0IfRNof57WgrN2+TS0jLOl7UrgxPDY9oLBje0rS3F9Psty
z2/af3pStJaoGvmkfdNmeQB7ah5JXESMsqrPlH4BNidq1n6iXMkz27tZ4zYPXdGw
bqtlXkDHeQdxlH4q2TpIcGjxgVaSew7gDKnBL36vuXByt39++Pnl/+6Ij7jUY8gD
iGICgj1m0bklArIoGtq6prtGH14OVo0DbuExQIDnTVCZHc9O2vKcL+sa0ARwG8/U
y7Gi2HsY6aIOrvuzREWckn8UpgJf2WDvNYwkCtcBHvMfnvwG6u2HoggItvC9JmJ1
l0cqwz1Ju77034dDLGLHI+7zyIUvqxZjOt8nKqVKHA2xc+RiAPwpexVMGKG2XD6w
/G5uttvMjyRtmENctMl1+UIpPSwVYbWCMERY5RwhOSlRK3UO4QmsYlaFBxfjxHOW
l6ZOmIQolFFDxPYz45KASCuNRBiWmfpC4Gg7sabDocG0DX3GuBLpBXWRHzfuwD/q
5iZyopYRluKMKsQXuSt8Xydj2P1dZ+Ei69ZyrwXE5Hp3niLSloQxG2n0wHSMTdvT
q543U4ax/YscEWOnFVVYbqE9OwY3qgOvMGj8AkEzRTGU8NMO2AJdCrqe5hqtNgJo
KYKI2hQCVpFOzb+d0MVFVmyfHpHNR49DVHHVvOr0DOQCgbP4dqx+UznSHov7sUCs
eAMZF+3FEfWfhDAisdruYxHWLB95OWB+qe2ACjCVkv4pXTbNI6VXpPtVa/r7o/c6
+ca8hrTVXrZq8EXaYXlYp22YBzW1cd4h0RhRQSfwSMPJMY3WPSeEDeYlhqbz0Lyb
tQMciQY9QSNykMYRBmMwYSjeTJbYOyNtQSy6rzQ7mgzzSLj0rJVHrPxR9fErNt2A
lH5JTnTU3HedPKJqRju0A8dcv+/MwnGNGzkTSjNdm/IyLjoEdICXd9q7c2eA5+sV
xPBI2MxdGFI+fQc8JpMUgbtaTUGbsu0iG51iWN24EZxVLjJnrjCXyvwhdflOMl/d
Iy6DnqFl+aeUN3T8PxHMP/LhQOez43s4AF3jPbR85L0CD+10YOlT1Q2UQ2c+Ixo+
yreh+kCq2ePicVh4z4GNNssgmHiv/yUt+vL3ZKe2TXJ1qr4eZqNEu6Glh+5+Z54q
M2Hr49m63RgKeFpR+BYo/l2cEks5nU8flz1SzvNSY2sAQ4g61+9tyRRoQzeOOjVz
W/rn5egwfvjhcb4QaZojpxnCTq2aeX79sfhLwcH4KwrfzIEqPb/7fTczJGMrR/PP
1EQ3daw1ezsBuOCNMKqMy+3+tENQDz2hd8VIBjQyh6EPYNF+FI0JSm071Y6SkjSF
f3rQwodfRy0q70iYhOFFdXw6SfA/dMhPatmAM7Okyi99EE5/dfSREHDVsuQsR99d
pJnFRT3WTL0SQbj0KO2H3CsWArrJPxZALSp5iEYZV8Gi+IlSgNKYsq4Fsxe3v4Hd
PQOCNjTslDY6uVSFUB9YrYZzAs+iBu/ZMRH6owIN+NmC6kLid4TzYauFWsDjlEvf
B2NY6TtVgWnxpHFEMlKroNVaPjgNIyipONYnBKpwgljOrzoIpJC1WqH+g+P1Q3gp
yUf3WXBKN+yKxmyMLrMjtTl84Mys40mjddOgYhuxAf64i/USC1KOHzBpJnWftLcA
OF39qi4UI/iOSVsnqMPHod+ami6YSrvxcr1HWfh/HQdP1541EjfwRPTQ6R90Rzfq
mc6CWTfxUee4IwPNH8ZgVOvN0Pk1XBugtviR48F/xBINOsLXHz8U4s2HakgdFBzS
jKCQGlFT4+Mg/VeaasBvKZL/JLkthG/FhyGPNv8FwTh8IfowXzvghpCgPJtbRsBj
Yy8pT0bGXZd1R2Ua1dydJvx9rD90ccahdWjz4HAwLa2I37g9L5qO9TyODr/MLfhc
4DfKN/JkuCi802Sv0bktVYNqBGhZiyoOSOjGZHPPZPgRLbyAFKNQ4ZCxMAGFcogR
SmQF/jEddUg03DYyuAiKUApJ50SovwxJBmeCnks27M4/7voILP8Qo5IY9Gb4wkhj
buIcsezhua8exbgB0BupjwXzm5t5/I9mT0qKoO75eI7WSDHxKE7bR+9HznLA50ha
CJ14k6O4Xx7v/rkfy1zWysYi5hEIRN40QO3a+P0R0SY7fF+I1Ziy45rtcdD/muRH
2qZYsJt6jEQM74MbSYNXkK2r+Gf37pIgk+zcsi9MOW4z71IhTj12aDRwUj30cVA5
h5RIjzDDG2sqIKxKUZo0KjkGIEJTQtG/GEv8YKa+cgPHuMVJN8SxpwvvvKY7A95x
yLAF3qYwyJQ+jMqAcwy2BMnoCyMy9MWeIfs7wfaLKX+An4Utcm1VCQeywJB7mAO4
gTt7qeh5LyqN7M3sPLBv+tHwjs1BDKN6IpXyOj+0NaiMonY25C1BGsWKnhXkhzaT
3rT+DNc2shvZwwUTcYS/kLK2LtP6H35MMtWDs9s3NR2tT4+OD5NynvcUEIL7a711
oQ1G+nj+badjeAIoe3K3j1mw2hCCbz9ONocwb1YSK9iPg+GjhbwRjCEML3/mHvxF
sVmWEZasbRUVrNWV/LzdCgBeWw1Iru6GVXIonGB1VfDXniHDGbg520B4wfHYkis/
w9MnQezCQtxTxgVR/cBLZL58FM3dLwlVQ7P2GukFeSsTeDy8VK5FDw4361kydR5I
VITjyLdQJjJLW7I1ymBGIptZ+XCTfcRATf20sf6NqzmnSFRV9w+5krD2Z9HsZOoN
LhCwpYCiV/SkLG8HR50FGCv3tch4mHbTlgU4fX4pR7is1JGL2UXEgtYUDpdGW0Zw
osy0BKTRRSKKdSbI0kjjWgc8yrEB5k2CeG0lod5OhyqS4qufS8M6h0aBKGX3M3sO
xrJ1hymGQ3TxbDwAsf8cRhTeQcx1ywLcvmw/9c6Oq4M79EgCOQV8ehqafwrbN+tK
c43rPdvhE/l5Z5abR+78nFSx9qyWmnnEsf3HcrvPhmz/7+iyfBSOGNHxXi1cceFM
LOSsRP4nH2Wq576TrFs4/6J1C8MUXl+Q+xNGey67Bgv+QQeJirp5+M1X6OjzS3V4
eFXkgrWz6kqpfR3zR80RhOl2c3s077o9qj5n7mqXKYHetUqBoyqam8iGDytcOy+/
IompietaTwjtXO4FMq47WEsXX7QyGauTP5KN2Q6zDAX+Z1wmbD4J8Xn15jSHN0Jz
WOfM06ZKWfmk2jYXqq+0ctGUvHTylMNSZb3+6g8IjK2BEwlsKAtOcKdOVYSoFjjW
4pX25nZZwk5GFPjdWjyvjrTTWlA/xODdRPGjnzCMo30tTCFFzA+M05s3I6WfefYz
TET67Qn7KZOH+P1jvgv5FrH1VKXmggVYn6W+6A1rstt//LndCRcYzlvP7kleyJO6
L5yhQDLjXSUTlA6zJrk+JMTT4BvfVlcsH+chX83xPQBprFZVB2rcb/gk44IkxTD0
o4+jATgp0Rck1SXdQVfg2JqkHWyvJ2eTgPxO6v7lxudmbz8M8qzlA7KAXpwmxqEh
kZb/h3Mvu2GqwRkh3Mez5X0uGDQYH5IN0D7SGsHfJPYKPdnJZOx90XbvSbNrCeyu
yO3y5X/lLLbJvcrMe2ogu9WbZ/vkwgxbImz4Vntb9zSPbMjsqAx+b+4rXuYnMUPJ
pzBXVm1uTp6ZbtPzSESbvy2ABwQVRqwbfWw4RHTPnibMZgJBSImAFV7RYep2Ocpc
TzY9KBEWkv3PJFdlvLllgQexDtQeXNhHGFMr97D4AgHwrKBQ/Jb+sq8uru4c8va2
kJTVtKIMKYEL7BbnGa323LpdmVV6U7Swk/ldpeLvurq/2EyubQUUVMno2zgT4X6V
urgMO+wAl0p/PYjlvpTOYKeQkF4IM1Y79FIICCJdFiIrSMMejDzEeaoZg2/6UIkt
OdSYr/ntOg5RABk5X/oS8tksOZH5nyRbLkFO1jx+DgNTfgZfnR1w2tP49tyGFM/o
ojz5qXcn7MHNVYaMgF2VcWaNRKJYWwt7iknSjUls5EkcaGhhnvNjhmkoJ3ZA4Q2K
IbStzN+d21PwwC8py+/JIssFRcrbprU++iixvSjMJiUiSfaEjhQAMWnaDXZQhPPO
Ljgj7gaffvK9og/ibjSqU+AZw0CHLWd1SJTSokjTJGFDscBBQds82IyiJiihCjjV
lI/jUI0z+qtS2YlHNUXCd5jr+rpsbC68b8pRSLrWVHG/GUu0ggwMWdqZZORRhkv2
/2HDG/esf9ApTadmCZd4UWCRx5FNfcFEYuWBWqYVY3yT89ZhTs3ZEntbBO4vf+so
bh4knLIVfVTULPaPkViWmZJzAg9ztloFgOT9vaX8Ut0hnkBUcED4ldgY/fyx+jup
LTO/HUbe+urGKYwC420lHXLGON0X8wF5uFeEd2W3hB6fMd4Xl0bCrk1bFRAwptRU
H1YtX9meO1BN8nmENrkegJPSEIhNGLsKfcpdgTRvyvv+jUDuNda4dt8zGGeGNRMj
xcpkel600P+a5SWZJp7HBI6lc5Hr34RCgMB6zWbGNT777NEuUUi86tlg6rI6pdys
f4FIjH8IrSUr3a3NDltooEGfKb2vLPiAT24l2oC4fdh5ykXmadQ7VFUBxsauToS+
isCkoX098UOTme64sfRSlApfltELTXGHME4jsiJvnuyH+fHs0rK1FNHZE77g+iER
8McZdklatLaGdACEzYTC0Ouk1y/KOQRptyQ5TFiT24dEJheHnosKN1a5701GlZ5I
HLPv77x8IvN9Na9b79UwkHRDMst4+6wn0hSfynOlDjnKrvFhIeQz2vuc60+7z2L7
niy+b/L36xRByBnbU8Ps3TD3VAE4XcjOBR5DsvluvPwpBZ+SPQAA+ZkVSlaVrBR6
wT3M/FsZpeScTFMpIoybD4vW/aaHd5LCQbkgaInxpqkn5LDhUEiq7sISnSmRfRbX
HT3Rok3lx8A6WTJqtRWYWQw5lcagVEzpW4xACj8qSK3zmFi28zxLHCFrPxldmZxm
RkFy0F/o0zxAFm4C27ZvLt9QpmbgaHDYJ6EoYI7YlZ81/1bIPE5bczJSBwkIW25K
RGhOY+YWlFgEvOz/fZRHGaZ1NuxyPPku4CXOu9+Iiz/6Tg1LlTRCnc17i55bdtxJ
YqyfyxA9188Z8x81JxPQGUBCP8KZKCU1o6Cygpn0jihFErakIDm/uUki65SNnXX6
SavYwaer8cnS1JzUnfBmE2dZo6jbmDv0x5Ec8bivLTDZDOTixtyLD/UUc4Pw2U3o
mGFS/XdD/1MkFrmNX3oKW/7t01Ovi3fblsmLGXUc0Vb7fILxoDlXHPldjQUN3xn2
W3b5ABeGdGaq/EJuioYjoKzPcaP0EsQ0/CbizFcd1yw45+2axwE2m0vO5+X13YI4
Sg8NBMzn2DOgNNrfaAQUKbXG0YTQ2ROKRTiU6UmvormWcvxffAEo8dUcxaHBsNBH
7d8XWyMdvl5Sw8+06SbgK+Nc7uJY43Yv33GyBchG8IUs1dlLZpd/I0pwrebAr7o1
J76pTa6bYpYNkAf53YRFJauc2nJogDk5aJaKgyDHBdZ5TgG3c1xic90GGDrdU6jZ
isRhKp4ok3Pb9ILyWAq/sbEDp7mu22xx+VZ8tdQyT5ickZ/1Gfn1lpMvOA23itbN
yC1EXYUu4UabgYQpcyMmLaVD/H2FYIuc4AZ6rqR6/rm2q6d4tqavTTLGTcrSFYIW
iDmlJ7Sx8hpzxqREpkqX2h33CuSteQddl9KLGn5Qx0dMHqEFzkKmE8Jzxi14MkTn
fVLLM51S0UDPQobBEHjupKNcNzBiQTP7oRhK5g/yKols01nltLjVLX3oYIYhkwq9
t3h1DsWgJnUnANHQ4EQDpNvHBBEiJPDVmjKkiPeDVNwQuIZK3b9ZCznwe/ANlc7o
A91ZMls5tAFib7vONOBPOABwA/qTRKDOR3tac/BebzAGU9IzfLCqJ2fRdQzLvUu/
CeX+oINYmY9CV2yibdb0iuqgyNhJstTsY1zmfLuiyJ5xftvscqm9vYxSkioN4XwY
m5VUgn1qCRXUmkW/V4TytgfsoD/2DlxGzVsDENxYU65SN6KjakMWsOV7/EslLIbF
YFso4hkyoj44bReN6I2kUleED+jUqPtj0edLnX8A+Bopft7jupU2xvgPxsDA//C8
KTfxorOUkizpWbk39k6K5J9KDsIzZJJfAh4v0req9x1usFNFcRQmXHbsrTLECttr
8xnBiE9GtbP04yjSGJpT3fTXKud9aPDbq6eoQp/d3eTLj1TblHZshhv5x2YOQoqG
SdL20iI+KHj6XsbkduGtnfUBZVZO8f9npXs3JuDbm2g8FMagyhOFg5Y9YfXY1SnB
vq1dp4Q6xvsqd+LV20/nCbjGkcLq/nrEc3m4gcIiCpdfEhyatP7BqvcF9RMEGULQ
8olrVvkW0hHCZFOONxEySfzk3m3bkBA3Q5qcbvhGrYKQBsihzAE67SFCdNgFn1Hr
meRVS4sNDUqGxEr4lka6ABwmAloH0IZmTSun1EGTai6KvlmYHy87Z0cLgYs3tc4J
y4zkfU//cDHjV6GutTel9FfM2P1d40npfxVrmyL9NvABQ+vfQoeLojl9KrEU8aqO
g0mz3hwCjRB1cdj57aovp58gKo5Mzi00cy8vV/0ytwLrXsDQM/uHvP8P1fJBw6jj
SSBIUmvdc4ycTJrVAqr2huk3PCahPESheXKbZOQ9TabROJ6Q+nZeIHl3y3I80YCW
VS1pDj4HN9QCNkErFI+impKuD//zEAN2iamxavAl13UK30x3PJFSBLpadJpzXve/
326mxVoPZAtmMkpeAeUYb+DzCDfMrn/ukbtXhWQ6xlBU3UVUC3SlNw+yLMdzmC4H
W0KlqnzEtxh5BVOC+JKKQzBmLVReqrtLbY3ZxjWQZ45eXplsQkwZbosOQC7mDu1c
r+dqXOv3JSo4PFcz746fCiUsLC0PW6A0qXq2S31XyoH4DfUD78UfCu2M2KIk5Knn
8tP8pGWjW42xrhJOem5COys3DX+HuDoe2idHJRhGx+I0TbA3pEDCUrRs+fKSlTH0
dt5BVerXKViQi34aPnzZ0SQpGhb+7TMpgNGtiWepYsStpgwSpMj3qP8cKvwG3PSb
PD9OP4UenhiHcBA5SWiCiCf+JSFoEg8fZwN32+f5NrTbutGhWzmoS3b621NEPN+I
v1UkEQ+w7KrIY+7jRPIGGWihUqSqz8SIshs/pw2ZwoYSyEcUCN/X9ezzCM/ADE1d
4k5oHzhluH7chymRsIpJmitkNal9NUFPdqs14iNmIifVuD+IwI7+q5/jfyudfw3Y
onbwmY47E0AlcukazZrSxVYb6HnlPPucMGGo56ygBKKCwViIIdaeZX/KyO15bJ35
i9sD4bwifOSveGQqLqO1jYjvzQBibJsvOAL4wmfi3o5MilS/dy/kfh6PCgs4+jTC
+i0Zde2TdNbMMIpDMaLK3UKQGR33F8PP90MVhtOVoFAgm6P+4N2CM1onQydYD6Pl
MTC1hCMgua1ZUpAScN+QlmIsW+nKTz3JqHfmGQ/aU6Wec4ZF1fU9XGX0q5QK4o+R
sbPTuLOJ3Sk8HgSS4t/98LWqTinI0q2bePgNAvK8yPWI11wExQH6pdUEmbUieWwd
qtkABAl5QFttgrkYTcK14pTyYyvqoCYM6iWm33wQuTWb0/tNjbNhTKrKV5Jmn4g+
AX0CocmHUIRsTfhvwun6o2Ml7L8Za7jXIBZKUkrk+xiDLP+Xw22W6JQov4jtfa5A
gZk3+pMh65X9uB6+ASHU8sNjx0bCym+gePrX4shBQB4FR4zMa5eFyVIVcSMWfczA
JsPChVMX7CY1fOkWo+pMmgvVQE7u+IiPOy0FBsJsnJrSMIcIm9Kpc5lWbDR/zXFJ
vtdE3T2F4uH80vAMBvyuD0zJEw+r5sW9t5TldoRS4M1qCjSyBjlxg4YsnPEnmM5p
3wcnTS1DmVVJPq/vFSEBcZHKRQws/jSu1WjwG44vOWbjh4M187P9dygGU+32/+GN
RUe/HceR3GHY9D92WzEaI/o5sqIW9guoh5xERkaYIQ47X4kXHQTph93zJ4e9vUKe
zanQk2RmCyPtVUeJyvN27G3EeL67F4kSRPA7EthnAZV53HEW8fQ8chplbp1ScQ/a
aHeEp4/1tEhkORjAbGY4yRgmOwyGjuMWbCsr7LofcAJM5LC5jYFv3CBtIQILk8GZ
KMqzu2WhQDPQaf6/kbSzL26GCTHk6aDHORR7pbczwp8Fgx/C3D5LfWJeE72pcg1f
bxgRtY87Lljb+PdkTgObUjM09vFx8Hc85kaNCT1i+4Tjz2XVS1tdJlOB5JCOIrhe
daMy4hX+vSD/g/O2S+9P3Hr3qQdeT7s9BpeO4YSHwUD4bkqRE4IzSn/KZJGln8+q
UbpvmosHAEdKO9MsIAJk2izU2u4Rr+oDn6wuGwMqJ9UYDpbo0YVoaDqqbRbb/DGY
t9uS6vVyJyxDIu6wIicWN1EkHJz81P7/woNtthOrK4vCa6TdplGplPhBXWXY91PX
kXq0Ck9LD51RR1/W+jWDSgOYbW4R+NQE0IdISkArid9RyNCmIeX9BOWCNijfswhN
+UCo5FLSMib1JX3RYXg8vmS688eiHw1aJxF6hJAIkVb78KxU+fs5Fbk47nuDyAtV
TbEFCC/oei3FtvMfZA/1WH+U02AlvC5JZCJeOGkS4eHwgETY/BfbtlboiZCa+a9u
X9WhB+GTokVfWgM91xf1fT80lKxZdOfmVbWSEk1l9N2gnvXfjrSagL0Q37S5tTcs
il4UQjOb+n1wbAwuu4DWe8glmaaztB5c6gRp5IgGkdZCqMXcmCy3uiMmUQfGOO8v
kZ3XJJD9Cx8OUSRdJK5ZHJaytuzBrDbF4zj2lsWSsjFRCxS8PaXU/D+dxkEbkeZ1
Ub9A29YquJxPKnxIspLYWyrxB53M3yWfakzw14pp9moNgCWtgu+GvvR3d9lTb9b0
qZGc/uxWWossQ1kmsyjbJyWnWXQ7gsBMtZsH/haydfLLOKWMQ6FqzceKDzQBIMFJ
jPPFaHPl9NxrF4rwBiR8nw9ANq/HxLCSC6IlSedr/vscjVjHsPds4P5H27LtGPmE
WH4tA0kAtW/2Tg+lLEXjRjBl/p2qG2nZZq+AdrhssehtPsjbd0QgLXecP7Ytqh15
LzG8bcqyogbUTMZpcJg0Weo94DU449tZH4mSODq2vJ6JiGgkltS0LcgSbbRSOVJE
rmurL1WzCbFxZo1nS7Anu3cO3OQFDrof0ZwyHyzChj2HQXVdIPtFePzX0wvsR0Jp
uEiEwgABlB31hXVanZmFEJpmLtVkwy2Zh3gxf1G2xQdWyH6x7zaNE3IfS9KOsEWq
LKRKr6FQjGXPwfQybzs5rQHwFNmSg3NEtDSxjjBYE2cj37kb126YqfQfJlCeGuYn
AnyYFudb9qPARm6cNA7I1uGSOYzBSwaulGIFU76inoQgKidC7bbMsIr+uATDUkHT
7fYkDftoiNU4e9oJ+m9A8TFT09YEeJQlh72AoPdNkj8tF5XPGcAgpW7osTDk/Atx
nE9fA7pwRmPeRvViUwu0/SrDFS6GIp8H2d3ympsrRxS8ztLr+xliYA2zXuLTRrxw
4a6GdLJbYEF+3X0YkiZuMcvVJ++sBgrWLcKT4WLemjqc8Guze+wT+V2TC6cZdf6v
pk2kvDZX1zk2YNFqiQ7Utz/ERooD/HV4LO36OtMBZQ6jkTfBmCpE+GN/+65BTXU3
0OJJMKJNGNqEu5o88vITIyeoYxL3Q66nAiR1Mvc1T4r3xky/avqEk6uXDRc71+Ui
BZX8Ko6CZ2Pk40j9O7fByli3vsoiMZlZKbuXvaHkEKz93BtgX7yzMrV0qi2LQXdF
shPwE+zJ6fOv4eBa1ad+VsABzEyKX/mCm9Xu0SlD+26tol9KT9uE7pOuhtj80Z3e
YAmc8yOj7Fehk8SYkG8cJ6Yh0aBI8YppSWf1Avj3WOTFErRuqs4H/k96SCR0TkHW
CZf2CcAR9pgO4LCOE+rw/sskbDXBY5JeDnuy8kmyGnDKWsOqxx85tBPkrmEU6Fle
FsRU9qp9vx3I8tmkiGj5Np/zapMP/ZpJsVFsVd/WbYxLsujRlRuMewFCzVOPP2KJ
Mr9JUE+YWyc/l01Qy0gFEFqHgLqweE20Be5X5UE0/XGfh69/RrMcjNYDLY/W/NC5
ZKVOMxRQ6G/RAAvUjhvXBcf+mxS3rqoJtK4Pm5Zl7z901NWx3tNQeJ2lyqRtiMTo
uOQXlG6/DlFzmAjthpGsqL747CtET6ZW1uGIQissgiIe5eCnFC7vpeIomjsl+kmH
AaCbPITd0MYFp+FNdU+V+jk/Rx5M+Qte5fX+jK9Sw3GU8fChqdhEFIMsm2k4Jxhi
SAeSl6CRyZHxZ+N8Sv/lbWvevjpOt/RqlQTh3YpxLMkt+D8lezaLygj+VLioThuQ
IS5pT+3YQA93QS8PEo3LjnuTq+oeftz/FZzIgjdkdLQkoEAKbeZaSWYRJ/91CwTT
EsgD1KzKXqumJ9WXhyXC2yR3YYjUFlVF2Hafm0lJXwhj1ZHFVx58OMjz/7T6urxk
ttYyOTy8K4CQrl1G8u4vhld4FjSg+hxLUNAXkJ4+vU+C8Wt/u+/q6QFUC6TbU73Y
VaTWE3TwCKbxaHU60MUCp/GOoJonyV/BcjjCE4/aiRcgb0DfPKCuf8Momb1AWOYE
DY6Yao/CkE0LOCILJSU4w0CNnTVGz06dSH/loG4zazbOUhD870Iipa7lXIGs2vCF
zUlUPJasMkzibjKzxsawLNy4V6Nj0RCx4//lPgJMfX+SERxQfHj0bwnH9zA9FhZv
jtXkZtX61Rh3bvBVISp1TKV4vCNV3cxKb0xpE2vRd4jXjkhwkMy7xsLhslNSeOOk
0mFWnTseOjPDnNBaKc4Pn0msduFcjXh5uN+3PxHHdVOz1F5yNym7kMQw3/P+fxAN
oUB5Egge58EqabWpBcEv7Ljw9cOw8qKdZJ/WxjtHcSJLN121XJxxWV8ceVtKWT5Z
aEHLkCJLO6C4eYwwhFFkjlW6xki6QHDlRwt+5De6JYdF1C9Meq35ZUbVazV2RpYE
CadIzAPDfq4ve507wsZeeysLdXga2aB5H+e05zTyu8ha1DUm50UJAkpytq+DPruS
3tlNJGC+enoFTqIgl93Ru8E8tWukPGJlbaDa872AgnzCPbsHoRKrvR2Sj4l70aD5
gsekd26BNwA4IT2OZSdtqtzL9+smnxs0uD1WA8JRMUcPWspbbsQqBEzTFx7Jifjm
p+M0ux1hwCOqUHFbqjrKN6wblZv8sinAAIg95xDOz4+0FotzD/zwrryYGdUnNTjv
IK3dCuPoNGdHDkqlavnFV7f1wv9/8xX0XE4Qj0oJKHy1pxBGmX4rcA8BiNte1iyK
M5nC78kumhDZW9BgEcFhoj4WVLRrmcpwkLKz8cJ2kgU4Et2SGY6aBPZoBME0lqWm
IjBkePkXuY9R6rJwqz7fpoM4i2cVAOdHjDeNZo1hA6iZDhD385zKbT0rQFxkAtaR
OgiMDruY/PHtRcMlhPuDWmNcecjacz4Ym+H6mycWnW3/gs1ZtM5Iq1nxOcbnY1wo
aDCbFEj6lV0MUukAMZPyHHHBn5S1ogtlf/7h0QlKBcy1VKUQIEgdJUp7EkUeKQi9
cLzfTIl0xiZ+cklQYD7XP81Uvrp3qfnPCzXl1YMmN8T75lhNJ1X0LYOFLCMEynZy
d+jLJVv3777R/7KPczQfggnJVZQiyEKBfeascTaUZPQvs8NiCaaUqW6ifKT5ks/H
bkNIuVRpz+L7ga5Hh5dtxjLSVXIfMD1OdKLrTjwergkbc6VlcP1+Rf+V5EUcQMeZ
YmqnGyevCKrdgtn4m7GAvJ8OO9CYgaMAqHgxPxXqDBYj9oYcsfHVhZ39/yJmt4o1
507gVVfprBxV8QqMVFiNk4IHRMjJDOskcXuRQurbZiel8WYqhWw+LUUiOve0QOEt
jJaDTur1vRcAD7sSPmCeGBIWm4AJGEaidCWqTDCHRia/6WR1hCP/xl3RvxVXQMJD
oJhIlZnSISKBZVdcVzSTB2vDrKWQq50ypYBIPwrsiLIXt/ZxPHMf9qioMcAyUY36
8JORf44aXEcsBmgC9uODrTBR92yGW3vdfjxgwZkEWZEENoT/wY+dzFjRyP7W+Hir
D3vadHamBKwc11Y3qUCFWwLhicYmhCGAjgOVcef1RKWhuJAyNeFOFzx49NT8cfLI
0mHro96gA6huByxECbbjnC+pWd8WLs1ahR91zksBxgQHeW2OsLQnpBAzqSGzNk8d
TP4WRYJqJuTNOqkA/+QTsXtnUrXXkxz+tjdOaJilMrC8ctHB2e8MubN+v/dAQfEy
j060NYoIMnh6TXudqECq7+3x1cIoGWEt3N2KBLr8k11KedIn9a2TOTmj7afz9bc7
HRuUADz/YsCNeNwyHJAcCik4kgkxqsY/+upDd7d9FAWGvVqvLT9C8GwzfhkIvKfk
19aBmJoAhu6QP6vhR0nk2TRUNlnnVikOOZCkgRNd0AZzzeVONe38mhraYDCvnLQV
1x8mmUOrusibvSttOYgmsikNA9bB0axZgGrM5qFm/C9LaUgUMkOk9sqLbOjvBeNN
9cT0D90JjNmvb2unytqFwhHGqGKs7HZ0BMpPjYVCiZ7I/wUag1eMoeQBiADl7XKs
U72mTiE1Do6PMhomDcu3Jmfnl+ilXzAVs5KlYdrbcojKhNJmC/bWLCQ6myWv9OhA
4bF+fIT8At9DY6lFOZhbd265MO8dnxpXDsgTY+t0xjWTzT88z31hQ4I2vVFue6vp
`protect END_PROTECTED
