`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI2Fy+ed5JZJGT3SqjGRa/0HP0PNgbSsLJU9ScuBR11z
pAE8NBCe0f3O7qqg9RMjLSCTLiIqCzG7jgnnb34XiLpfk5W3yuK6Bn0fMfd6uNyw
RYd9HgTS7x+b7ASSx73QLHvzv+PfQw8gPxPqR14rcTsadFCxUdf+1szViKczPfLt
ndmg21TJclUOhRSaU5xN2zDXf6YS9vweHi/S7ocuR/b2Of7xy3G1G+tJWmq50Byu
`protect END_PROTECTED
