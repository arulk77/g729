`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SU0TMvMpZ03N4vRnycIXPr5sTnf0O4WeVjNb9z0R3RTv
uRWyD65SLRZAbgpgo+zLvOqvnwNib5CiXuXrdIp2XGnshdvNPdaGtuIFHCTfjl8W
zVxKJkbRtEM47Aw4mFwDS7d9YAWLpB8cdaIMr+kpCQVzIb+jE45bVeWouTyg08gu
qtdVI/L6sIjD9x62nq2tUXNraW36LrWO/uZZ3nJYD2NRyNcWFiFiyL1iFb2FVTnp
yuFQQ45rhPfN4mi0Eqy45iuPvasbnIqwK5s7YYI1snj4AErKmOZ8IlfpNHGlqW49
zWWQckW2oEVnBRlRtiEJuNr11kuimOUVEBO1AgDCrYHQUMxVOFL4r4yOoWVO1K2J
ve48O8SuqFAKwA3dp9ZPe9IGVERdIOfWfhqGs9qwlg+C0IUy4bXUT6hUsK6RVxY5
Z/hba84pgdiFFqRybRYnXtvJjxarV9BEl12SNjgG9pkeVAKlVlgL+7b65zqjR4aR
ZoGP6MTrkudpl1Z9zK5b9G2bSIGwYShYW0Ii4EMxBgr9EdBaBbJfXTPnCAkAG1pk
xspZWXve9ZYovk/6WGIKVDMA3++I+Krr2Ir6a9XdrBXAGHOdtKzQCbGA2/PvfUKH
zF9JbpnSg5iCgA0CxOujZlSIStSRTdnNknxX6LTX7u6vcAT0hjcEY+46vMnVV2lq
6Z10t7Byttuv6BlDfds1z0uV9D2xsgKMiPj2b1WlBXInjqT076Dregr208Afa5Z1
kY2rrQDRiu+2+AWn6chqequaOLGZlYykD4KYExWvt8yQYLMBAqEyjj5sSWcKi0Hy
pXp+6r+Gpa3UW+WUrVSDS26KaOF5sfxD4t0mS5hnYCgPvWLWEcAmgtDqQQaJt4Ij
TIGLLcFuyN7RfGVXdB1tXSIQ43x88SDmzrFOMAKul1kN785OvYAmUyE2XF9HTe30
`protect END_PROTECTED
