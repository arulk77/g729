`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLoCszoLYk6jZ4M7InycJGV+qI0DSRCUWnxsuVny3If3
PMFR2dkRscInF2vd5s4EIZCyg4UDjrJ2waOeTUjb8suB/pN5pT7nzpD2XLYscbrq
CYHiqv/hK99XEcNM7/ll8VPliWdOC/Vmi4YCeFxemEYKkzr63Xf8e7qZfwSufLoQ
kP6BS1dAlc8YOWx6xZdCYPEycmHF04FkgG7MAwpH8joX6JpHkOTMUswxrAw4NgLi
YRwlh8uZsihPlSCGCRVW2oD1pKwKGsBTvDQd1/tDHnlpedxiIEDuCw3POM8/egUn
rUOrEuU1Bd/BtbZCylnHnPm4LLe7fucz3AzqHLTpUTdmQtpW6Dtth3CjOQXstjlM
`protect END_PROTECTED
