`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDRcMTnkgI+Z+kCcec43UO0FfiBYMtZPs2n2Gvrdx9gb
yWyLz22k4a1B4jJMe1xK6n5QEI2ca/JuJr8kCtaSUEbc2EgYdnWjjW4/y7fapMEQ
CFgQgxtRG1CtS1nlXFiTs2CYmjrlWcHQcf5uIt+Ju0GwuAEOAvRxyFKVBQMoG/m9
D3EvRpTwYeLgrKb3vjkBa/vudhO5sv5OZHsaCfP+AtkfmoNHI9VokPnFCyvU9t8x
znwm2qsoWTFzlzNDCNY4ig==
`protect END_PROTECTED
