`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAxQ0KIwIx2zqrj3swG8NySvZNzYxlYVuBJiOUt+kmoa
PDnV6m0dryhP33FB9NUaomnMiWxOASkp/KpPp7PewoD+6CbbfFUK7+/Ubf8V+C2/
KxKqq9RjBP3Yb/SSX5FJARXFjpLFy0be2Czo7kELPa3WMhQqV1T4wOOSRPRKDX1H
`protect END_PROTECTED
