`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFktpu6lzoBultYlb5fCh2eQyiNexrWHpwB8r9F8KS90
bZTrdz1IOHYfbAw2zZjF7SDQHvCLaD3pN62rAC9RJJUihftmMhfMeX6o0x74AZaG
97tE15vCicz1bMbHD/t7qJ+OsUm1RlHkV0FyCU5VQv5TGcHKLcvTU0n74hF8E2TI
`protect END_PROTECTED
