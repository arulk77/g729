`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aUbcZFjLXirin5Cl+WK36KEeG8VTJyNu/OCKlGMt7gjG
NXObnLv6/SFq+s8mmVr8j0+e3ZY4TB/tIQP9w5drGyxDdQnnO23MmGQ9TxFNc5XB
EgeBK2IcXmIodPVdS8dvHbINWUZR1+5T9EsxHIuTS06hDKkzsdcy/vNc5uOltxID
WR7GlHf/abZQZTjWJiAzXRYcVTQpEWIayxuvI3zVl3k0/2Cp6p+M+vRPiuIMS0/A
julLengXzC5Fi/nwTjXJxE0pv5amddvkwx//2UVdK70=
`protect END_PROTECTED
