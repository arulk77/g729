`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
hTF0lQNpeswqu0MNaWp8rdxesK2XR6zYW4LhnJYblHk/1IlZGU6dnOT3Aup89LID
n7X2tSb5igSIztlaTNO7yAvBEaqIm08iQIuFyMv2SwiUdEuEDcqX5jNZ6s3I8MnN
Z3MG7MllGb9gXXn/RxIT4N+qFdoCpHUHnXKgYn1pScU9VCMZpcrk4+n0mX8PfQ3m
03J21NidWBfcm6BbLuwJfu/5jW6mF46iKYF/DZwag4KY19MNmSc0siP+Z7yOJ+pJ
ANY2+zYQykNicTu7l3Pb7QDWdhcH7PkIK8R3ynJrK2zyI35LDvBu6e3x8piwVsUr
ZVq3getdMBaVnpr5GUoEVwsBqfjb30ODBYFRwDrpNQr/0BDw0mCDB3rAzHInaIgj
oLXCZm75QRCv9VF47lM6kzjvgVVFAgR4oiQNB5auN3J3u6QgKsGIeeTByCGNivWL
jd6UYf0JY3lfutt0MNEYB6s15lMX1EXN3t20NIDMIwTEmLj1A+r3SLlusizLbGbL
CK4IxeqZTQfs/cIckMBprdeozlctiKz8B/hb+3JVPOnjnSj0RbkdIqZeCXi3C0FG
FLjZvV+d6QZv3VhtHqCCAz9I39PzlgXqK3o5kq1yvui1Oube9MVl4u4hUIP2ineL
RR3LE1p1Ps69bKvv9Cz9MaftePg6Fgdcu8oet/Ex93ZHAxZ+uLr7dfy52SoIfzmf
907B3hhfQEHrOmZTE82KH4Z7TmuQs9nirglbthElM//Ewe9WqbEqgbYAwpy/6zDy
lwKTqQ909BONMVneH/tsdzYMVz2X4Bjl1DW9vgc63yvx8gOvUnzVYKb8Oxnyb4LL
+yUZfZNWbkL0jYiFJfrX3lpDGRyp4KBXIQOA/WEXGczjG9Zl5uUCbaquOnFr2apl
yD5lqbhYvCccflcpmrSJ8QxkZizq2oNlKc64XtYZowy5XOLGfu62iuze04ymrT9L
TZaE0DHFu4ZIFdh1AEPYZrHW08RwUr++FXqM4DvIzzx3KNAU64iK54yh1g4vm3QO
YML6uND1PvHqBJt27/IPCMyIpeM13Lyp+ZUnKXeEObGGVxGF60PfSBwc9ezKpUhs
oRU7GcvyPP61xWVdPJFvcmhjLHupeaUnvkrvMssZ0xNhZhLspbkiApyvbyrZyNcV
I7AcG/Yp/PX1y7pdDSurWx0RHdkJDGORuy7k9Z0jgRkkMD8Abgq0qUv/UqFGi9Wi
ZBnYZY9eWPnQeWG2aBTFz2GGqRCWRIw5F804GWYvAcS4LF2NBFty5qlE1iK0sHp4
h4xUCN0bPyRIoxHTo4czH8HKE0dD4TEm7L4mb1ApwLr+8zK87yhJxDroRUrOWIr+
qUAMIXsgo9qm4U5qfLDiSZsknSqLnqYu8BVK6y2vArVwpPjz6nN4nG4dsM9+oUBd
X8+PQAwPylQk6a4i8GJsjDGjsd4QEClpXA4v1ui45gKJ4DTk7CanGWZWDQWsS9RT
026cc8VdaGfTFHgAUI0CGjAzPhDVKPcr2OceRAd+1pKA9Qs7LSto24EL44Vsy+80
HHQtgK1ckw5OUIZtswsaldXo3fROpQpeL6u67EA20vvSEbINjfpUgD5yJsrFOanx
pNGinYQCeVUAWYV+T4OoJtsqe7FVgbVMerOFi3m0WHMUpyF383AI/cc2tMdIkzOV
Tgpz4NzAYrEaBP+GA70G5aH+cWS0B7bzS25mSWxGE7xvmp7IHgiKx7jJGIrlF0Vl
peKZuIZi53fwH1yUv7fV6FIX3yWei7Xt+bSk0hKNIVWePSpn5gaibr5Q1fwFimfd
PFnz7nockQOiemSfYeAj4HK8Duw2hpK7zTMltyhqF+2bUPTUA/1fvP5WrSP3tnB2
16ruXNxwQr4gwjVToFYIQzIf2pA1HH73xc3G4wWNlQ1zOaJgNzXZqi6HUgq+1T2W
4ZrQD2URT4THhOmNcHJ3k4BnL9+RzMGZ899k2WnBdrpxDS8+KGcO8ufzayHXSVQC
`protect END_PROTECTED
