`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL0TtehT3p194KEFEb6fLoimXa506umFz6nB62TbC16x
D0nlzaJlGlgMA6ULhYrwlJkG6RWP5g/nmHYVfzqWtIEbhF/jalB1eGq09/Euw+yn
TNz+VkEu6VBtLDJfieg1FPMDQmq5ZapLXdm9DZ3XFDaPu8POsxup5iXF2Bv9CYlY
FZBUBZ6fvFDYSALG7n7rTASZ8Iuznioo+K0gP4BmFRlKIYQAszgNAF+JKo6kTGBQ
qt+nn7GUJgXYSLshe65dc9quPo1JhsdKrDLIVTHolVypQ9v28VtYcVQRaBAbhWBU
xuyjbgMPOlgihbcvEUDOFk4BXIC9CfBiLMgx33RZMZlTvdVwTS3PD0iaRDWB1Gks
h/HCGsN0/Rm0q7gVF+CL54CGrvMQCpy5xpoxwo8qF4MWGD37gkTw9/0jsjX543lS
ireCssCqTPq4aIAU8usS/kK029WLtzCtXM7UfBXjMTFEVJwy7T5WQGnkQDekBWTk
xZLIwxR3gLpKy3YpjC4hE5CCYW6EGI9yk549hFLsj6TnLyKUzRIY/AtABUjQvNEM
13XpQEfjEVzg4TOgqHG0OssH9KRr0Ptih87KwpD1piFbydhGl7t+5SrbyLLrumBp
nD3jqI4ub/miyWRPzCncROg599lx/zCeZlT8W3onGcNdsvenJJcmERK6qWN2mcXD
`protect END_PROTECTED
