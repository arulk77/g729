`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
K15/5zg2yz5wMadmUMgJMBtTtXzQFdD8PVvLyL/GcIksbgs6a4nNOFRC9b6kmxV2
/xMugRJCqys3qyR5CgSLpemJDilqbPbXCFW2Nr1N3JZ3jXUlokHOMq+mFwqWVFeo
YtympGxM066U/MdHOtXrWoFM+Li4G0IhS3ruK+VIny7BhkOMiTAtP0QOTjWcZkKj
EUg5QxMO6rX4zC/DmckTPm8f7IC8vxU87Z4dy6Hpbd7SXVSiCx28mblC4kNKunnc
GYsRdFJb4Pwu8+sywoyH3ghF3MtKi9McoT3mhRuU2NU2w/L3UwympKpUNDHT/l3w
7RolDkioTT+dWAX77aCEFvcaekqObhnCv3Va8ED4aTfZAL7bzPt+w9CaO/pJgW9a
ftMIKWxPFr/pXB1lC/6F/S1PurGC8mYYo9BXuK+Ss7xQWDgIW/ywI9eU6NQsNetG
zEr1P52BuLZK3dLgCYHAaIaP4qyaLFthQo+vhQE2Ig4UkiftK7PkKw8ZrcKfYgxB
/flR3wTsi1v0X2bbAgO7qjeZPOfkIzG3QdfPE51b/uL/qbrlrMZGvZI27d3GU6PP
nvj4rX3mk/7WV89+Atc1Uu1sG8brJQXseWu0NsmUBgfoARiCGc8raNKuh+lSGzgh
dej34gPm+ZTMFaXnGbJdraTRHCnotYq1HpsYAn4DUa4G0pQndfpHX1WmHLmIKq/P
`protect END_PROTECTED
