`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
cqr/NMfR0p5RUysmVawiy8grFw6ABkDxFhKcsewssmJuDP9KImBEnpznb+HZ6gMV
062D0wLRfGEp2iSgZvLnijqiXNMhPBbCxO2lTjEq1j/N/NaPy0ssjND0YarLdp/v
BZQiJINxQKivJM5L+pdFkLWHtg4SEEStOZD28+ZQPgxoyG/8veCJn6qMFinsGklr
UgE6ZXzP6hCMadje5lv9LK3EWKxdQ0hCfVx8DSv8FpU=
`protect END_PROTECTED
