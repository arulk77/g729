`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41IUlYiyiD6rr1IZtQdg0ksfJ13Mb1VSLOdgahbY5JO8
ypP6qQ/n1S+/sxkx6F18Ozfk1X7lVqL+tKXgH+0wPRn+jqRl9U8o7+RGXtis4M2X
Pl4FC8Eoob8c5ooXyylgmzkTERgZwvIhtSgSVIG5xXt5vx2XGImgObln7QRRbUPU
IZUOIu62cN1Ajy6MBkGtUl429Fi1S9HQxGbh0q6mAxix1f90QJllXTlWXEEZN61U
1ElKXshsIkxhiELGaKn+nM8pZDaPH5P/fpUNZMnwP6sxhZ0p3YIE1egKsoPCpH1y
ckuYule772Y8KJt6OZkshQ==
`protect END_PROTECTED
