`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePD73sLlPVREk3AR7+2u+xf0UHH22mhLZYeYY2znNoKr
FnCVhmN4gUm9dtrRBb9NQC/DNFRYldo28tlIXOz3aKFHscdbcampIsGnSMuesw5/
qWHPS7ase6GeSq4eyUGgJ7WQloG2l8qId3J352ohHLIpOVoxiAfV1vAYMrAirNQL
jQTdJbS0fhdiq3iqtqpqZpWbqjw2MpYuJ3q7PuSwWw8tUmnlPEm/fXo/y+R1VGpe
aFBbyWj9js3nbWCc4RbhvFmbG3azpUcKhTCkDJqqowRpKLud5GQxPdgkpimzh2sE
o3Qt828NvV7dDPflkJtR8RU8Khuujkcgo/xImlwX+S4KoiFop4eVEmmOQfqBYKy6
qGfGFH5cA9NY5xUr/+6vxztVzULMIRfd6/KJ/rfWwhfm4D7iMhfjEu++4ryoLLUs
2yzBqU/D6IyHi0dS1e6nXzPCsYK2u8EqKTGqQfmIgoi56zMlV2NyrmOA2RpJFX5/
fKxntFqdv3nCyTCyy1vPGsyu6wBjukU6sj/QtYDREOURzz+J2HOmiZS5E+352W1J
`protect END_PROTECTED
