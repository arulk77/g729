`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/sUE9/5nOBTyZ61RWZIMRDxAWCAv5sGzY85rFilNc7o
ngo1PVTADR8ug8hUJbi/RjKEPGmBZgXibuM6X+QxEYPNDgEADZaiiC7shWI+uerh
t6eVNi7gddrvM6uPHZyqEtkJVBYbdcALoLCSvO3bUubZQvj+/KMNwBA2/SaarRbd
xPasyHea16HfXBB8E8WHYzWgnjzo4kun4LTQhq3xFAo1Yi+OsSNI0liBGbF8O+t3
UqSiYR96hT2AH9kj0XMnOcJDb+Hi113wX0pk8Xe7pds=
`protect END_PROTECTED
