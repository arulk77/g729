`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveA97mUaXVENBcHwVmN/n/tOES/al1ksQy8U6K1v1eAzG
PX8TVu8p0B4fb34vG/1g9l6Yobbtn+y6L/2TNsK7CJXV7k5MuS6atbO83yHFnyof
CvFWkyivXRlEZ8OjuHqp4JMTkT144CaH3cz9BI38+THO1irnwI3cPlfLXtKb4WXV
PnFl8TN7Fvg6VcHa32UQX4e41S6tXqaslb4oXw4StwB8PgiJIaCV6cN2qbwixPLt
Mhui54dmwHgoTwxGNUrCayu6FizihI5H7H83+WKp2Fcx+dpzM0lb+6zl9O/syh2a
ZhQ4o4yb1gtIJfQ/4q4dWhanSLyq+WAhREFtHwd0eJmEzYdmeKzxz5oatBdXMut7
ZEC38W8xP2I8PJ9Y3lczGw==
`protect END_PROTECTED
