`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48CN1pRVd4UDp32Rxppbhxnd44zeT+slpJtJwMeazUWv
rtkeJWY7Ta7ecnZzpvAYuSjx20y27VvrV1r+qWM9vluOns3l7W8z12bbIwlsegUe
q4VSAp3v1eiTXaZKHI+DcC2S0fnTaDZDTR6S6ocOrGFR8zKfHg16sJV3cnLCM93z
gwRCc4HvVQQeum2JAEHkynlmdFWhvVZx+Mj36PVsJ/oS1xQUwUr9yue/CGYuISpq
3vQ8DKdOO+ftcMCmaHgvBMZuo9YHKtkeh9svsuNznPdLmdAxP0XUgbGoXseWGLbb
B4RuMWM6/lTcgZCLN5Yp9YDZswfZ5iI41PLHmLuxQuR+i530KhUGiHuFkebk8WIK
OVBzyF7m2EFWyAOIkh1Grw==
`protect END_PROTECTED
