`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCgdx+Eo1jkQMn3nj8TYynSIWvqsETvsaS5mBOXu1Twy
ymqIA3Sv9uTkAXZKCNjSSFxPzjwIRlqkPzaa7OIsbZjoPPebKcQLKKdJv5zf+FSg
sJt4yRzJz1PZO+vFzTJyiS+iluONb/5ChZZFgk3G5NOy/andLr5fF1CZgpAWY/2L
OtR3crZZlj/6UnVsWF8xjqGqbzsi8vPkXHVzPWDHZ5oNRUpp9Pe1XGE2flgJ2gV2
BUEFvkD8hvdya5UkjhDKLHbqdeO02o/y20c+Cfi/6OMMCK65IxVFmL2Aiz1hY2og
bt1mCiimMR1q1o9mYhL7LlKZDifUz4mBi08eMgsI3B4XrgdfEjfucdVqssHup9Vs
26kA5wBfU6nzDQrP0HOF8vEGbiB8YQoGQIOm+0KLMgjFnRA43/cW4fiv0YUIpAYs
82EbTiZwjBWRLIkYj0c/GH869snNEons3HIkU+30tKCDZ0K7bmofTK7FMjAoLQ5y
U0W1gbF+QQITXGci8oUUMYHNdsXLYOuOo/NSYnyEOR4VgI0KTKw7vUBQukfE0QfV
ZS94uj/dH5UjDtVOUTielJIlWw5+UJaq+r/iPTJevLJFETjUpV96h5wpvlO/956s
RMGIfQy9h+4hDhixfAmj+gPPQD0KTvjCMt78MNAbY8SPr4vD9aBAH5tnBK9d5dI/
`protect END_PROTECTED
