`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK/4dU8ycPNcWe1K3YXNcPYrbMHZe3YFD7ReP/x6z5FN
Hi5MKweR2G9m5TLKUhNX9inVRo9YgJ389xHTW7xnz7y18Mn/e4UgCyMzdcL1T/NW
DPL35scIra7YVfTlqkaZ/3kwWNL27HjlXbT34zbbG+y1ozvcjkzh/R5gsQs4vHg8
+7VNCtd6/qNkTKvBNUBlW/uEjxK5NYaZk4p42RX4VFIocaY07pCaea+ZjvTLlifp
6QtKLShWB29uPNa6vswSqU9H1yn03L9n7g5j+YRDbf1OijoLL2JVsMP8bV+QDnWO
+vvfizUV1D3pvM4eGSxnWydV5sHJxiqjfdYulek8D2LY4wg5X7A9P2IYVHAkFULG
PhRsk65rpKd/okurUZjR8GcI03TjGgqxaOq0mggkP9HR6BBDLKpeQ7DuTm00Hu9O
ccbpp7Xoz7tB+T0bePwr0e/o94zMPTtsypUpGw/lnB9ximiLwQON8hVkoN0DKfjO
eibFtvtstwvA4yhe1kHc4xGBO10B0e2FjmDgp4FFWxu91rq1kE6hEL1hShfCl2Br
`protect END_PROTECTED
