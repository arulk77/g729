`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
U3eFg4y590/kC2Iq8tmrpEP8nJvD8Ia0sVYmVG9iyRtyG5WHNDRcHV/eMFiQdik0
FZs+t50ibXz+b7s/uPgcyt1s533Ybx0lYWFFAynI8V2LjcEdTAORMgZos/EPjdxY
DmggIgwXJUZ2v9In6wjX1+UGzfsi7tog4vW+sQkA39K6x137rS1A0DCve1k2G8N1
YhXM5udJMg6kjkJs6Gdia4IecBddjjF9gvyT4iDzFNST7qcNzu3KUwpYXhXyWuO0
OrP4gqg0j39owk3w3RynMgPcWs9MLll2EEDNcizwmD6q2hPaMcs0kxJkP9tRCm6f
KETru20hRkGsVVYJqX8iPrQ2/zaWa+ou2olSv+c8xML5FYxTttkOR1iKpwADIjG/
nAmZvsSyNyneTDgIh7KvqoidL4yRCPqzL+YTjM5oZn96IsoXcD4GsYagx1dcpHEg
Zql0TZjAKfm06e5CO1rFrWbV0tsJwou8Z5+TtO9ol2hVcI+DdrujHRRTB+cH7hhv
xBrF4scK/C4AoHpS2VUMIRulVhZnGQWmk+vSNohyDl6NhUGxEHQfEqxxnLvYeAAT
I0wHQdq8nirOtGU/83yVkQzl6E5uw/YgUuIOP04FEMCT9U5fJUjs9rxe/ymaBTwt
JkyirQzTAvmAUoaS2hMAiadl3dImVl7j/5JVfn3TdqVBSCEL7yeFI29YSdzgq0VO
+rmapisgKXlxAii8F/KZ7Q==
`protect END_PROTECTED
