`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHJw5cTClz1QeW+4W3ScWb6Ozqo8aRmZ+BlwyaZNr9TO
g2vzNTVscfm5fnkUPVEDaAIvQB8t+TwE8InM/ejFP7ThikCIlFrwEUdAIWgD/RBB
PgKGLM96M6VOQ4U9rtpAmA2rrDiVGhu7YZCqJs5xwohNgI7mH5jl+yZiRP4O01kr
0yix9OUMrExKuuFA4EhyKI6xqqWqTMJJ2HBrNANPEC6Itc8XKsSCm+e4OuJ8wGG5
`protect END_PROTECTED
