`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePqkVvUcytp3rNjmtgDIBobAZXrhJb/04YKw0+2m8Ow1
J9omeIB3ZFwY3gryKsOmBI5Dc0tm8jK85QowshhD3b9M9IKvH9QnivXlJrJpS4q+
RuiSHaaWuwBuEpbDQaZ0ok53gPJ23SszzXUHLOJ7YbP1i93J1HoZSP1mF9B9+dHf
K8MdFmhcFGEOO98h6+2OtnyofUyVwHBPzvOSOnxdIUzOVyuq8/YKmDr/QyPdRM55
j+hVnbYmnb3SkomZ6aDNFQW0BqriC732obWKRaPIMfqwVMWWHYP9TaIOOMD2Pupp
5LWznh8J+O/Lk7SBHWQCwQ7HP6KXVRnN6yswzAR36VTupSsfMOSN1hml565BH6lO
ug4Cl9TMiIHyvVByi2zIY50EbmARn9MaQ+2S1wPRdDFZ2pEg+g2A9YYgrcg1laLb
t1l6+/W+LZDtMdJjBFJr1w==
`protect END_PROTECTED
