`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN/kr61SVcdR+6e0LRT6azCpUQAGhK55NhK6i1tZYqVDM
QoCBDziFen3kFw0d72iGebSx/Ygmx7aDMr+ku810pdrZXnpiVSrT2Z5/z2TI/3L/
PCjuq4BlY/idiNDaAmHKS9lxwBh5xrH+A5tDbnH8awemwSl5qN/rdSH+VoPdpPL6
3KCF7uO7icsENY8cBTwsDugCVIdCG0qTZiPXQFRtuwkN+dNF8hxAoxGQXiEyy8Eg
5rD+XmhgpjQOOxnJhTLKy/REFZ0Q0B3Z2nNeg+ffSxIX06d9wknYSv0+zHKcCfK/
vS1xRGf4YAIpfseeZZb92xO7Wljb/IecZVJsvLwM/3MUQijZDaDCpbG+yhly+O7z
9JXBUzb+Ry3VVlaiWOB48QJLysgd9g0Lu8tdzsOqMv1x2INBgkOatKbdbloC50a0
djlZ+Anprsph4u/oqTK0B59WAwUXRArHM3Aw/KQLPXs5+VY7GiJDvSU1zVeOQMOG
cHbGtTBELadjTxPkBdetMzdzf+e3jqQex1vldGosX3DwPlhkxDe3YsTcyEPOvpe/
2iICriFpIPQA+4TvmV9HI1H5LjIvpNdS41SlIF8WTa2NEKmdQi6zFrIKvmqHKrvG
Ht5Nin9YAdD4VU5B8t4EqUCKCj7uMTuvzJGwpj9Ll1oBR8qjaBtep3Odgo4IqpQT
0Va8jALvRI9pBKoDPMwMcCwArjus5Lw0CMsVWyuyQZlbnrZyX/ZWyp1Sx/0JJcg2
b668abQeZ+QotDD69vCn+MlS6JW2VDwJMiY/TeT96kWnnHrpgAsst7zdSztBpjI2
GVvT/bI9sr+3AWAPoAuzqZgyz4DoyIq4RhNKagE9w939d9JU1pNuUZ3sR1JSVeGT
4zij9Zi5HRdlfCvWFfhjfNRZBPfsZ8g3fKurNgqO9hRPB271WEsNtqxVGrh+Akyx
h+7O/YgTYZWmLq6sDXGjBQWPmCCto2dZckVHv9W+k+85C28hJuJr6qJYLE1k/PRu
TJfc6fUmgWMze+bfrY7q5pMvV/QjR7qmmCmfDWN8E0bDrSvdpbNZGhW9PLxyRESu
luh2JUxop75qk58R+qkv7CUDThYn+sK5q26OiA9qhRbG1WFWewrvikh0sWeCqejQ
uRxh3PuZT3rGK8+dqLLvr6HwxEG+e2t28ML1PY8zfpm26BJPXs3BYW05XWt+Fjtl
4Jpoh/oFRO9FznsWZm7BvnUKK0mwHYj1InKue+qL3KbuakEvpnOB0bXJrxbSx+Z+
b785zBLC2DzXcl6Jk2iDejBbeHyj2HB5XADsa1GyArDy69UeWA1mxTYMhbZUPqBk
oT+neOOFQAnYEs4cCdl6iHoiY431MDxLhcrDIKmMukUghMErQzWTELgVpzjpkoJ6
Fw8CbEnQ5egV2XcCDSKyMJPCmOEeWXJ1Rc3HqvG6CGdbuvW8aLqQbEUpzTVnjChp
sPO1fEjDD40ObGPfPusOaQezI8sKRpHH3Zhm3YE+B0QdMLItltxFSJkGOgN7as4u
8nkjyemxfb979iCosDjPSGItd4NOdG4MCtAy2UtXDWJ4iQ0Hx9XJI1usqaTBZFSc
9uFaZ7BefRliUQsk/E+qtOGCs0pS/IoYq2h6Tec+9+JnIyGqO67GGY5sR830odnl
WKPW5sh8Nw2C1WkexSZFIVICWma+AGbehgAbrRH+5CJh9FAb29KwtOta8Zn3AiY6
Jq+HizwoR6yCDiKpVcpzS4HHow+N32aCnxIcEiwAQtRtBkp8DPLclqykTr1izPKB
z+4/AaXaKojvQk8eEXM6Lj4687fPS5P6PcVFAcnx1SC4tc7AnI6cL709tTYifuiM
WPdgNPyI56pgVL5KWJ9pglGpXI1TYnkIPS7+2TTjFcKNe1H6F3pL/DVmWoXN5TXi
YNQ31DaxyKU1+iV/kFJCjSI7OrkFcouZzsIMg6iJlvc=
`protect END_PROTECTED
