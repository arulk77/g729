`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDcJ98Exi0Hn5OG6FAaxyJPHsbYa3odmF0btoO/H51A7
miJ4iIKIVBoqtOTrxhn8tLAqjUX/lrabsO+f8mohmYAx1w5TfqLjxUY6YT41oSGb
8LkMg8W9soB9Ijp1wOp8MEnehFllDN04Pxu8C4cviA7YxCUmb0E/IW2qC5T2XUlh
6HLfeIzuXiHKzrGimMXlrhbVa5YnrQA6fmj/7NTnBP0SUgry71jj+kXej/vxcMGP
RfDYsf57ATZ8OXRUiYOW7w==
`protect END_PROTECTED
