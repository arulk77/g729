`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEv6cmqzhwTbXUzIYwAqQHbR9g5HALKm4I482uxsDun7
AaHxh8z2uYn4vkkJua7+NMZr51zZb4mVqN9Rn5f3G+IGilgZSQ1aC4zWuokkIqPn
CKgxj+yTU94z+je+9YbcP7z6w4JAFLyo2ILrAc2V94HCBtXItGwOIpIi/oUBNy5/
kZ2+N7LI+abdm56PtzuRlAXamdQcGBSOuyLhSjNPCdtUqbyKAgcnVVbD5ugXlc8w
Xw8NvJTVFPgjP6Zb6dIKwbBbthmDMu1BJIxzCuoE0E8GrkBqA+ax8qtK8a0Y3E9B
eIChbC8WYvV/nzW3CFnM1HFOndlY+70pdwAa9vroOk6yLxQIK0n4b2uSyqltbFdp
Eq8tL6i5DIm9l1y99l8ar+jXwX8vJ2IJOj9miR0xsU07MduQFB4lsMY7eugiCBjl
T6mb8jRqde7IJVyzPe+DnkDpYqF3DjWEd0nc62FOk7wcK1zmxqRC/pizw6vHUHGL
`protect END_PROTECTED
