`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43YPOb+K4lT2ysLonhsn0f7uBU6UU//rlDtFTgTtuRXI
ZhYT+G+xAbSEjuo1JJ09q2ARwfFU5j4pfFGTnudicGpMfZvgQM7SqJL0VJjt0gbv
/qx1vGZioBuYJi4c8zkt6LF8AABiRE3ru9gpqpITbvY3NYkXTv36BXQ+Mfq0qN9H
r88QupVB95FcOqU/J11hvehdyYNl2R5Ti6zaAuxwW885g3TBQC8O4ZdKDy7KJZQa
JxZkDDFvgIgePm+H1uruezwUcWPxXO+IED/bf2DdyjbfYeneHu3iumiLbDFuL2ye
BPYTFMvqxj2Qukd1qHyNEA==
`protect END_PROTECTED
