`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMb3dPgHw+FHUYyVWeB3uA21/cHJOqLK+bgkxFn7uT/8
CTH3GgE40UW8Kggig2Gs+NBBSaRk/ylH4ph/fTGFuzx9qUOvFnd43c/DFcS8Ikoq
aCG8wUuOOLqsEfPIHqP8jo9A8I5K+BORhXCjXrxgxb/ubjUog8B9y0oaAp3uiPv4
6hXMp8Cn7EMWR6wSuzab/Fy24ZT93engx2h6d3XEHUcHWrydJFKhcdw7ZS2dpEUZ
Yh6+3cvIVBLPxArknm/PFzLWXz2w9bWzXxnE2PVKpXqMe+YsK5jSCEHEVT89ocHZ
pjVqyiyL0z5uHzmAwJa3Eg==
`protect END_PROTECTED
