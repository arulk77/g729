`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+Or3YrwFV4XvoCCZK7tbbT00alZ4Gy95P2T7+VxGfRcstt2TYLudhKr5eaKnjRlB
y/Zv/3fXW2FHVlnH8BZ43m5kOPldcgYLDZ2kX9R6Ak2P5/rRRufTNNJ53PeV2tOS
fRX5OZbEg1YVVz1cMMZphmOckRXZtgiJMe5TWfLYXhTeGBrA2LPzW1P10cLBInFL
6uEM6Fvu1nass2K6PtRjGAL7jC/l2WPMx4VVreyrTinnsgEHcNLb4MGQfrJPLOpy
Nv+SMKXe04B2198dmtuExfq0q6cTvCzggqLUlrdx2KPlgI5pQg3woBBtxfFwiq42
S8g72C+6bbpgoe+XIFfWVh9z1119+ew7+aLsnrgPd8Hup/V0GLOxanctav4Bv0bb
/jrpf7Io7GUIjvZklhLl9VSrr29a1dr76IMXG6VaP/Q=
`protect END_PROTECTED
