`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveC2PwwTJ98wsKW4lVCUUYn9JMOU8k49dm9PW10wFhAyJ
BrCR3B4riPSJuGBeLtmjgBbhq79BnxcDt9fP2yA+FFrqC8r38whpCtV0ue8pSY4A
kCntA1nzj+XbcbWnlk2vT+ixrtAC2i4KK16gVTRQD8gtLQs0i6z5DyxgInmkaeLK
PodGTSoUi/DS3d/EVUeUFnHgqQFct2dlNT9+2IhEUr9QXwzSp2xFcnkrNovqmF8k
xOiiFRt/3qNR79GDwcPYwiDIHSvEV/Slza2hfBA386k1O+kjtb/y3uYeh3P7XlSI
hYuvL9cNQruV5ImsgI3WQE6H79oKuxj75+KfT2p+RgMjwaugVdxZi2HqHD3IYvVu
9+d7TRrfDGDjY6NNO8g8GwKyesdG/pFXDxdSV+kLS/iWIlsdrFcSHcqH3QQhZ2aX
cjICnyTezYCPmnoCMyLW5TMuMbmce/4PQFu+RTm1z7EWoBTdgLZC4zKkN4jUYBet
5vvG4lxXH1Cy3U4kJNw0SqoX+IognSuQPnNDfPyRLeR2oBkt7AoHVaWCUuNou/Xh
LwNQKqwAwhy6W48zGLYDxp0Fvem04ccMCUOfIiyWx78BzX4XgiTHiC5QRErvNLwC
OWyQh1uGauBk2V356us9OQFF/J+gCRc5/NpXpFCVE60It/LI5PF0Eav7r9iqOjZI
`protect END_PROTECTED
