`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAW3Ya7ZUJIutuv60eoFUNQCqzJ2pGkb7N+vX4URQrws
e2s4jDl1vnb1doSQpwaOxLETtQUieeXHkriHZ2W2+qlDiDXPb5X5MV1DIp0gBJWJ
mA2uzivAwuzI/fhdm5wGkNDR2Ce7BYKDpIGf9Z1t+vjASNnIAwgNkhMWOcCwuPTC
3efRv++2+026G7p2Wy+sXLKQj7boQtlUfkTtMzguoCaDoAXUrua11egH9IGGovhk
sibCKQhbEplUrkhCQZbv6yv9UgnTKQ17ZXFv5NPM+shgaTuTUaRYErl+p8nPDEmn
1tQGvD025EVwt76gb6BdP3RDR1EINBVQMezn4lMVzDRd/sCmKc3QCo0kUUcyZ+JK
JM40UZX6GFsO++oY6QvrNg==
`protect END_PROTECTED
