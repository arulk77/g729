`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP1GG/zEthDQHXv+7GNooqpTj5XrijCPe+L8EzmU5zgB
YOzlenVRqtiB6cYpPZkqAoBIKEBeiRhw54Yx2isvJwVOVjjR53c+VmB/jaNnj1eZ
aKTyEMPIIbVNV9fy6x9GvKvCULhLf3DCe17gu7R75sTiLXMFrk2hZ7w1Ovn/CdXw
j+x9OFWUErQgFLcTrhvtzGjH2x/39bunTNt6t1P/0XKPKjEyse9pZpm6KJ5/XjhG
P0CfTVNNT4UVRG/Tk9kBVCwRozsZAB+AEygyI0UpKp2SnS6PmZeprvWaKsjnRiwF
2fJEfotViNZdLBmw2lOzf62BqgAstXTEIkSU0y+DaI+st6PzdbBewwT7IqIemv5W
ywTuGssnh2FHSTsmLlsylfsJMQ7LI750gTFlLXZFriTwEoyNlfmRKqfLDf9v9mFW
JQ8577HRU5V0ORJXS7Ok89NLQngmCSQnV1RxZXTLBBlqBEeLVio5cRer/5sfbDlW
KSpSiqcIoPutbq6N7Ku6mD9xZzCgKDKqVS23u6mbow+I3oYxV+yPcAFrVIYumPHa
`protect END_PROTECTED
