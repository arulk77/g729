`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL81brPGdUE6rKYuBe0mtsN0hM6O540M1HHEzKGzAnSFTi
TM+SV/hDIvEHQDS2WQ9K5QPjekIqSjIu/BOWe+x1Ss6cmFNnAocoeBzU1fR1PVJu
vFng74qdMkwjyztpnl5+NBjG2WQ6TDUKt5HFlzmJwrcIUFaLGjovLDJNceNNSNXJ
5crQPEN+DTKP/053V3ZmzS8D64+CZOTPquqQILNpc2+Q1kJ6Apz0lXHhWoBMqsiR
hYtN2sWGZiynRnEXnNFEjXuqMcOQ0rIQr52pAYnJ3+6NUMpVnRXOMsbkXYWgOD6f
Y7zo0Gq7fICvKjT0LMd+kfeLN3qpA/e2eKzFYsuI8hBDriOgRyNShEngzUHQEwFd
CCogkktIS6VPPm9M9OSBUC0G+duyzh3NkIHJ15S7mgE=
`protect END_PROTECTED
