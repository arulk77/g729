`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu417DXDYA2LdwXzkjT89mE4lK4Dc+vN+7J4tbqH4GKMe8
7tQLT1w8k87kVDj4hN+IIYeWKcT//R4f0TL9P5if0GGdgaGcyDKDQx8nEPBxLlpc
rLQTuUxUWIqhcEM8P5uI1tiQiA+c/auvyaXXoSrmwGi0/c2R+Kyp8YaJWaeTLzm4
gIgFTY58j3rCj/SH/e8ArBorcJc0G5ReN81xuCU0d6CFFDRKPs53BhHC8k0a7bX8
P5zC0WOgnT/nfeys6KJVJAzKI5RvWK9nw5LCdyH7s+0I/qGF6adf5sEcxZ37Pusj
XnEPSlkRO1ADeBfiORg6iA==
`protect END_PROTECTED
