`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkfPD2eHNcPwtsphQBqIKeufV/pm1ROOBFkZAvcPaR619
qlEXxpbWj2woJJE5enVlXDD0V0ECUaJGEUcW7YTZ3IOpGbhbqysCj9FEl18/GKKZ
zJEdI+aKFiNJDHvqk9olXthMct3wg8wAm3b1GrotwhFjjJR2DYNpRGFSuMMX8bFy
ZX5XGQlkwBU/AJ1S5onMl6Fi/trwVV1SvT6P9JvAuI97t7h89waqQqEQQwVyHivM
n5VrPmVDkAfMnU6o92kaCOkFLKQ6BfHawLZNDhe18PMMSmen7U/rFU7H+TmYW0OE
sHpC1OuCFxI/AxzGVEqBURUWAPevSH8zkO7lCQNQtv3RZRq5MnuF1/ClL83d9VW2
dym4vzTfaHq/ukE6CHnB4XEGFVE+t3k8fct0vj2tFFCvQyOIyp2yJSMt3ml2wLeX
UOyTAkGjuXXsBoFFpgiggvQ5EDKtyecTXXfRUXPhEtf230MN3u2/U86ajKWZWksC
F6lRvnHIB4DlkzSkmPVlAws8AIeVJf5HLuMT0PvKw/mu9iaGVdV3SgpOCBv/1BWx
`protect END_PROTECTED
