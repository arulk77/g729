`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
sSd38QaV9jsHeeHUAGmtrQTdHClHAFEvMcpPvJCydt60Uw+bpiizMeIxa6NomviT
98a1j10mcmH1UxQFTxbOZaIDsp9leYOX85WSHuicc/OdIPoNB3Swo/NLWgNuf0lg
6aoLP9xM8rHsKsmsi9fr8fXejd2c9ISwAu2oqWg+u6Iv/QbUgwzUQj06zDEQdv2P
hSnCDhp2t9fdk8n1+pc3qwNyF9GhqxHqOg6V4h5PdeX2p9JV2bA5XnWlWK7x2WX2
Fjyk/L9yutwIS8QA1zhJDkzekaHJHNK4zjk3hbNGyoNwGxB66vPadv8cePQCYYRt
PElcsprRGAPTYys3pq4mofs+XxDbTA8iHChHrck3uAI=
`protect END_PROTECTED
