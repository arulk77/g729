`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aUuyKt/CX1iPqn1pcIAmxFYa4WHLMydVdGIEIRyi5KJn
yN+t+Dl6eGeb/bckNwn06q2+REKKzSFmqM2PzwA3j/2ZikckMoHtUqwdDcCwXasu
BM+QIX4kJcMJaimkdc3MsyWlh0UQWJGwISVPyRhEsU7Nu6OXxhzqvY13PihB5CNI
AvTiu5jq+do6v495eXs2bP9ttmAyLB3/aJEqCYtLLRkoy7TGXMvweEqnLxFmFJt0
h3iqNJimvflHMifK+MrkfW7i2gSyW9ULqL7ZTfZcztRr1nkzykweJnyNvBzHvy0Q
/ksE45+xnluIfFOJta7OyziQt2eJUS+e82vIBfOLJ2/Cknr9GQTTr05ScLlG3YjN
S6Ca0FTXVj6T6xY+XFH7wR3gLh6idRQK2H5VZl67QZmg1rSht5yITEvGWSfB/68X
iRuzWWUGRQBhkFNAYz6P55MjWE7KXfPWt7pMXBq9c2MJUvF/UnYlHU7PWHuswwb7
seqM8BnQOo0NdtYsUx33EHYSaZLc5s3fOd0TTySpXBuROdWPKgB5bX4T8AeLyvBa
4NCXxPkrMOI8arPW/SZi1vkkLkbLI+Hd2Emzdy5F969glphFM84BwIfNwi5kWAmI
3v6y4AJeknfFa/zWyFdPiePlq2gdex1ge28TZzr+0zGuUmWJVG2Faptb/vFMhBv2
018PB4fTOnG5Mmvek4W33BgqCPxTDRIZ8epme19gpyoAIu0tMI9apPZNH8uyhLMr
xKLw//fgwjfB92X33Y9gsd//o6iIFo7X6/aJuOBKDjHezQ2So0zNXhZqhZ9+p5oI
qB2uXdHuwhTT7MQIns6Ssbgpk9Yi1cvaEhdVj3gtVkzBRW9RhhlhbXDy/4Zp8Aka
Xr2yte9jIj1/zhPb2IoqRmA2ncJ6YpSVrtU5bYhpbN9JqK+fUx8bWKBaHtNBvR96
X2hLsfuAl6510VKprSGYH3C7Z3Ky0IBY+Sv+/U4kA4OBoeo4bY/LOIA3jWe1A66J
dR4OZwSW0ZYtZcMIMmIzzN4xP/E9ej3cJ+1RrNPHcqVTXwfMQRrYP2K5DEe0ejD7
8tvOlcu0XKY+/vrthQKlxje+KKWZ6c/KsxTAPmbIZXSF79sdfmdYj370nnRPxfDw
Zua6tBf7CPCiOgVanzq2mwnNrrkOoIJlNsP0W9PsDL/YHEiqUZUqkLQMtjoCs4eW
8RJTKz+vTKsBU6mfAYBZVFlcBeE3MovfN3W+B/GjaQBo2fQih/HMSjB0fojwhmN/
SKldFX/iuYEkNRHMXEWG6125ismz61+kHl3FaEM3+8LQP/yV89TgYrXwNAqPWrwn
BIEc+kFH7Kz+nWn/wENjfty+HDTR5RKuEaMYtTQLWT8vbcqeZ9Tad05VaKZWZabo
1Xhwv1cpOx9wK4FcAcxJ+P3yW33pBBQkUoYHbUP94yl0dKvg0MfpO5abNXpTTwn+
yFkO4+yTI1oCIVKW7pVhPv5DxDiR0TfkmgUo2RvccS/IuYzA37Zvu5uInzQEHWu8
zoFG/p6QW0ZTxWG+cgAKPPPH64xPfFmf0JKxkjGSGg6o/hsW42V+LfK4wrZN6cl7
REYeDdRJDeVrXN5VdaVXm2PY9g+i0hGPRiz1KOTLyz2C0zlHQqbofIjXjK2Or30b
Ci+itOISTrt2Arxr2/WSUAA9y+ZcxecOnK7tFJkC4Mdomu1OV1VqiS6Xa/FnK7j0
UfGlRKTN9Q4QskdCDqAu3KfaNy46TDBzHoaxu3/a5r4+1r2jwBIwYPyf9hSfBCbf
QqnZ8oJMP2NZLUKp3sgMu4B25gc1rje8Yp20mODMeBt9qg44vdq76fQcF3Y84uRM
8cPnKfNyY9GAXVNDL8G0PHrtq7Nm44y4eFBZn5QlBrQrLNwE0CyP/Ex0/L+U/zDN
XQc48AIJcXL3BIcTsweRLVr5twO666xZa0Q97q6FFgIGbiIOrytVmF7tVUdBe01u
YZUNcw+M7I9qhlcK11lbNBmCcXgi02QKvdhaUrum1WnsI1kC4c8JbZsxupjSKa8U
GnR3+rqTltLIXwqti+c1gfbtzcTAmoe4ZK941NKETwPKnj9/SXue2k2E+xfwYk7J
DuFz+zjsFyVB5LQzBz2ziXlRauffEvH61T/5ZKO8Zt+LFJm/G4ZeqkGBn5lBCy6u
yvnAmHjsxC1XWq/+wQpFyjsyRt4tvF7VXTHhTel+Y4986jx0qgswdFi8op2721jP
CbtTof1AKvqb2jfLf5LVhACRteXyifKHeQPtDqSbloftg+rtJYhaAA/ctEoOmLbg
PP1LTPNtYTnTpli9lFJCz+TceqhZ3+ULzzFQVs9U1/9YtBeDQ9bNbjMDkiysz1EB
V/NXj5zxi9Igf6/byCJn7nwzRpQ9r6n7WWG8l+6UYKQDBc+4yt/PSek1jaBcktZG
oaQfecAsEqVAS+zO+HY0rZO/JqojNZbaTfS1rzvZ5BctrWjhkVjLhXdPK9fXpdHv
UnyBwZSdUFmXEiM8KGcbSOXsgfrb1gCK2wkNHTWAgC/LgvTZlHa95OdHBSdPXGo/
xKrOA+jzZRchbJg+C7kyjOeuOcO/5oTdwm9F9+7g4CzTQsBM3CXzbJOIVMx0Jllq
prBZIyufl0OLw1TwXJ+po0IiQskuvM2rqRbV2JgrNF00gbqSF9zDFn+OKknO+sWu
Q96+Rqz35AITtLDvVq9j/F22oL7hthz7+hJHGxZp6Utyl2qx4G7NhXO6LSe983Mc
HGAmbERPAhHXh4rJG3axEjPxuTFA7A8xid6KtZ4+q7zFd+0Q9rxoojcYsdcHjE8f
1FG7fZ/pq5s3v7Hpmf4Xfcbx3ebu1nZJPqY5gHw9u9sb4y2ihjZeB2ThIwUOwk6R
Elu1WwDs332YetOwBspV6UeD8qUFIINCZL66BQyFUaXFbb0N7gdyCIzupspFNy0x
AiLZ8FOepNS30PbT7gYvbHlx4QwWpt1ZP8RktTpNW92IHKzZviEuxEck5an01L7M
mDxKEsHXa2fQIdwh6cavk6WG8MEekn8627/mlic6sAEdGTdirxtZlpYGb4mslNX2
nqZngiFiwVGeuRmyCBF/YJI8R8reMue5DUzoaEC6rrkZcIZLmb1Zp8dWoa6N0VLc
ol7Ea268Y+qEo1KeoWBLzYr1LR4Dl0fl/6H8HRNW1IPBsFWMGbyUiqoKg1Mcwl6P
Te8j+9EG91DlOI2P1NLlNz3exoX5KCucf3u5wtlhcZbHUr+R2bhmsRVWZqo35yih
7yISJGsPozbe7jdOGkXWITC+OTbnd6e1JzC0dRtU8ctMv4gyYfbXarItjTVqBCnG
CiImFfwMmPYVdPGS5xUud58sVbTFnSe0oe/pBBC1lO/q+IOx34/ZSXPsD5SH/FPs
TXaioAA5qDV2NgOmNyQ38rGl6BtbZVLL7dOXvyzPrpl7Z6LHAcE3rGdH7+47EOgN
hzjMu+5G1nZMF5b6az8mp/fCKW2nU0wmUOnKIjPfWdsZcITxDt25RQeGDT7duU9I
Jd/QOYDo2RU31C7XqVjKwg9OM/pD2CDfSpko/I8T2mgR/ieediL0heffTYICdBvl
X75FaXgqjukNZ0Y8nTtXmXRJozuE4Ae01Sj5ELxqmE0xMcdkIVBTcvfubCgHDV4x
rfnPG9im21cox2xT4aAkKh42sp26L+Wxxqa/aqtS2ekn188G+re4qbZmXhPZI2FI
Fl15Z81hDZLSsq9sZmehjvDL5dZMVRvmdIjs1nES2VhvimS1+amcgxolbLk8ote2
HHTz24zz1CP6fnIvqABQxUidH0SLUHn0nTHChEUq2oHGY4Zr7ctB3hZ+GYBW+1QW
45Rkz0vWGDaqKS4pbTy+DQHFABkmSkPzVBdOpx3gB93YH8NsgpYMLk6mQ9osoqAz
UEsqhmKFUxIwdZxjYcIJdH2haMDgJPGd4hWcIb/1XLpm1L2BkzljKrMdKoP4wlkO
H7mGH3SRu8Au/9IC705vPqkYBUZL1a0Jxe7y+2VFiUPBe8qDzhEhOXWfyGGwmyVj
syiT/KYcT7IPkvZcyAxpOXsAj2Cj645327d/YpX/gH0lkGZ7UmP94HeHUrRfCN1m
KfYRjwT/JkVSrhmw8WWyfDuM2f8NjtgNZCCQrSCFbggu212bznDpzWAVQnuiUpEF
3L6oRlisEqi40SU1De/ifS4WSqA/Cs0FfG1fkgdxcoVL9c5FTWEbfwKohhavhN2t
nUQhv7CgPHfYVS+aKjjaCyAl1aQ96Ry9+IyvuSv698MzOBcJdK/O/f6WScFkq6BJ
UNXFCZl6OaCKHXMy7iN6v9FzHuLsH1AIJK5/Jgzm4lhGktQU9pNu2F5V/NarSQZW
K3M+D3dNULucl7UNJZKPKirIkn2Jvkix2fTqpnJFpiSvIvWsXPsv1f4AfWneA+CS
WM54MRbxMVeSAONezUzxWn66lSsF9Zcjj5E+VoahSqX+jDDJQj1CWYp83+Cig9K6
9tdomN5MjzwHZozpua4v5n4cpIxq9/IohyUbaLwpB12pQEO8gwWhSZcYI9qFf07R
s+nvLHocLBWCvnqU+wPBU/LhoyV+7Lq9Bhfw9d9VT9OO5XHI2mmt5wwjp9xTdTEG
`protect END_PROTECTED
