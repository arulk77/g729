`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1acd/lBG3RHwvD5/BaVhhB7lYI5lcZJVCSgSV1Jb3uAwh
DuWks76RRBC3VeOQi0fwcG1CDZmV1LYBUi+7VY7bVyydpziYbBcMkUXDZbzh8f1I
nksDFP2ekwxQblTdOdPFI3HyRxL9ZX3rsA7qzwOkUOWSHiOUpU9VI60gQPRX+J55
gVw4lDUR+/i4jVWr0Qz8Ny2QO05XDb2XuXcAika0PaRwJOGki91K8YcHDL8pUY3B
xfDAECmZULVrpwO3/IF/hlTvthXLC70Pg0xGdL0iS4Hdu7spQrz5BdC13qhOywyk
cDz89oyuuiKN+l9y+FD9G9e0sAg37gqWzUaKS48vqAGtlbJQRJUn4+v/6QKC+yDz
Xo+v73GRwnUZBMccYtaoFgCyQPVtcDk7vXElWyDvRKLhveZpO7GmisQXn8tUswdc
ozEyszxdD8OoL3txlrYvmi4P6TqElecIJ+hxAvAnOJhbolNWEveGFKGjNXdRsHZ4
kay1H2ApXo5xYRAAXLt9i9fXrOGmYcP9W9uHuaA4YEROM3FIG8RTMiyNOA+LwNJA
g1cYnphIM2Rr62xqpIcdih8iomYa9pKV9WcggiOOMhFgmB9DR6eiuEGhqWAFBPvV
r9suy+wOzagL4C0ZWuM8RMGZiRtqSOb9r6G8Uf5J5NwmlwKFmcHZD4wyK7qxKAPy
4GkHquYAXyYYRB/Gk86IGzUqIa93bHmwHiWK4hg31g9Ki6+R+KnId08EGXaEiF3Y
DExVJaL9L65ufSJdo81KRUAcAMJOko7kSRvKs5KCWoj7ONK9yv5fyAcA2AVYgwnf
acgaM/7fR1+LoaSkPiziQH5yQxitoBROp7/X35f6PO6C7LAc41xf6EIW/euMJysP
gPoos/yUhY3dfqkcdF6ZMdElqQ1BjT4GDfh96RjKdX4O09eAiSe2v7zdnBhkx1OY
y7WP2tL3jpHF/E4Na9hvlEJmZwFvr8pUxMz3lPlYAipRG7u2bQs3Bamcgc7fZm4H
E89Gbv7oCf/+AQAkJ9Wm01yrz3ut5OwraZB3BrSdmTfoSxwhJnchYW151SR1tU8j
udhVUylDNONeJwJ+1Bf0ZbDgb7AeFa85SWYHPOFzx3w/qkCX7XUjm6iRvJ3vKPRI
J5/iAv+eQPQt2X8UuDy9TWbcp8HYA5VVfb68DpsJEkg5v63QYZ3c7v+0KmWDgAcJ
Ovs/U1WDDDptyxrdx97Ze6wd/lUZeCRDRK0d1gEzIqZp9SllKIlsZ3ny9OGgs9OV
d0alufZI9KemqgWYrYleFP6Fak+2jWqgOxGjWL3NABlsVLDo1sgKZoaKaeSv499g
s85VO5Gc/HB8EsYnQB8hoU0HTX0I08H3paco2KVwC3UxFD/BF7x0CSh1pt6TYIpy
eQkPTHle7lZzAsd0ZzWSzoyPFuTxTVmzq0ouhA+6lsgoML7NchCNWPVq/lp30rrX
nyO7DrYBA0gFdaVxih835DqicXXpH3s7GOHy577vECJC0qM4cY0TX/b0VoQ0SaHs
Q/ifZR27ADmIdhG3+ZT9m7HVMZ+HkrkaAjjDbeAkaMlEeg3yoxFEPj+kC+WO68Jq
0501KWwNIsKYcZ7cGfzDW6heZlpTzNHrA1uBfzgd3lto5FglRElups6pPBAnT2lj
4yavMHJ1rBGa34UGMSQiEMBEfz3Xwu113hIQpxz1hssSr2GNoiYGWfHZ8R3uHW3c
lraZH6TDjmg9LKLd5cidtb/YE+1sokEnq/qvw/5KVQ5ii9cNJkXj4x0VkBaCHwZU
2+DpO6aOBDfvztynC5/bzYTOtWPPBST8ie+Bivg5I+U=
`protect END_PROTECTED
