`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveC849KSpo8/M5XzkpxY1n9KxPs3qSf7iT1oD+PaCsjj5
Xzf1hSccHohEJezyzs5aKzp3f+Se5/yz/S2KQ28srkuJiJrRkK2Of/7ZtXySs1J9
XcGu4VQIyKYtfsL8QSOaE0CD7h/v5d3/h4xp17drf921Eun5uZOeMZwAmxC61Pxp
JJX05o35ToE2pLWYx6dE/+XntFIgTih29cOhTsq752HXWF4snggt9inH03qT2l6H
fdjKCa10zoGIeitDZFe6fEwU+VYpLSzjLkv66UC4h0jbXM+vGil+bfQhJOQymR3a
jCRzds9djrxWKKbZYmfO9g==
`protect END_PROTECTED
