`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aRC2/jiiPGHNG2DZW1SBfr8mHjffUbFMWdhhnTkf3ADs
/Mv8wXIRoQukMowZCuHQ8eJB7xt3SAszwkq+0OF7cd+TFvkR+a/xPl8rFZAkYRmK
yT9GexiPTNyjmkLL/+xidx6LST4JOePjdQO+2exS+FyE+SGiMxitaDPli+q84Chd
ZeJ3HK/XCv2PhRHSO4V7rVxEwE58x/aXflQZn1XvbjNwoqJmOmwTsfsdud5LBBVp
6iLJ6Pd/9h+Yr9ulqJaIALg9eVQ1Yw82G/RKNHazK5gOY6xgc9y395c5dZpWHknk
7HwraCiU3k0hcnlmrhJxftfkAvUhX+M89GK9gbJ2jgc5KBBMORuGlCivyyIXNH7i
j5HojVTDnZKhfXR7XqKS6v80GbLjIU+Kt7s41mxTn3wwRAFrO3BSQIQToE1mhWKd
mLbu6w1i0NgeJ5rzwDmHGmVFsMBmsebEh3iW3j9xjuPxUcy65CR331Vv0tB48r6B
lYo0PdT8IWUV+5dJCqTtAH4LPPYbP6pOQCHQXbGb+IqPrfHNxa5oGgpTNOs37gxa
QflvUiGSX56uxKKGIQiHAp/yLKq2GSYUK5H4xmsJIKkaeSHThfXxq96sh1slZNIK
xzP49bdWfddiJ92Y6jYZW9zVeAjG4VqYP4JlnWKJ0leG0jXOUKK3lsmpW4Jpfq38
ATY2/v4lkFxB4LiNZmPVYUjN97S0K+nslVcNZyU8aaX2EPj9ju7+VmLPbwox00iD
5vquh86RrM7+VxahfG7jWMHZpugKGdClTfnvHH7UgobdEvJu30KL/yzqg+3pny5p
DD+r7D/S2IYLUxW9yNPMJxTX5wN26QTOp/eM6pN6GIS35PPtj4efAYRkQ4ik3t8s
N7imdCbE1NaUROj7XQfMorZxeF5sYZ/Ob8tnCo6mkMwOhnsbII18+8YDFAcg13yw
BFekUFE1d5xsbkRhgdvm4JTH0SAs19UoO+N9800TdSqy01Lyex23M2/tethWH84T
X27dIsd9JMqeInXu8HiRCEAAReUrvIge+eDLSh5ywUkiZdBta6RA2NYVeaxguH9Z
VeR24BbM2FDiZoai0EZ1P4F6kfx0EaxNyjc8tzoia0kq11nRUjVfyNt4Z1PvBNfl
YWRFYVRbJVg/DPNF1SFArA==
`protect END_PROTECTED
