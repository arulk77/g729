`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKIdy/B/BhiPRCETG6KN8MkkUshC5xj5fx52lcMOdEmp
FqUawTeem7cniYDCMTt3cMO9cT454UvM/t57RPvUS22eLFM0XfC+OGHCJRpU1J9n
mnGj2CtvhFTLfDCMW+HjaAHjA7ViJvBkuVft00vuFX00VCjYDMjueuRwFzFTgd3c
UrLATZqKTSC+VOW2VWn3NfkLIoYt/dIO0x0o05A6xOiVqFuYxm2m//hl3AUdDpRg
`protect END_PROTECTED
