`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveH+XJKn0CTa00fJWaOYUkdGr8sm0Y+DmGnqAjkdXqsxT
jcikAiEpd09LaDMfhibcBrGTZf9uih5NFLTE2dCUIO3FgHKtItUf2e/Tb26cX2jg
nPqAsyg7l6cbZKfVZudiROymy5PCStn1OsQSxeyRDxlcACnAGM2mSTrZOtiBz6Xq
cXXXAyjC1K/Im5GeHJzAvxIGm0pRS0L9N3Ws2Nu68oYV1XW1/9Oc6/3sR4HRixcg
10wEK1ZZMJUvy/YMa+i6M1zXr7QgxS9FguEJzTx6QUWTOYoXdsbKPLOmnKKRUVag
xh4ZkxPcZUeHhvK298qN9G4diXQ1AUNbj3I61Twec2FZDh8FR/g9Wi0IA+SJcaVd
IMlGSXd9b27FbRYZUSIbBJc5IDnTHIOc5s+edCPIpho09fjPO5NsDxlE9wb14VIR
c8XmLkSQQ1x2JPRB1j/EzlmSuOHOkGH8jNkAeBTyYWgXol4ZAm+qVY4MuiWh5ZN4
rZh18xSJbMlTo7WlO6zg0rZXenkMWyVnm1pYZnNkUX0uw6Eq+kK3oIzl0KEsdmOF
`protect END_PROTECTED
