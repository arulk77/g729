`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCIYB2n3c09Q1JVQ4V8k+TmdpTtKOkODFXInrK2DjUJ6
WaysqnPRbCv6u2F+fch1DYnPvJ9tmH2tqM3lv5xRRhD3caQ//wAHUtlaFWWq8yBY
H9JE8nepWZVNCLrRQCfF8648wV2Oho8GpDpi2at86hUaXAe3cgRwu3OSPgwLiPft
NPgeqYxl57ueKwtU6/7krQ==
`protect END_PROTECTED
