`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveE+MkiT80gib8gvNBEWjbJQ3fHj0GkWmw4QuXDiv7RWM
1K7ymMe/XrXtSyk/qdi7P3zkw7xUSMeILPyS06tuNwtbx8hg0ptzEKRHi32JWyYu
ijkFTuO5P5HC5KN2lSui/XMOen16/cUxQaxxWhrRJoSD61soUBPLtpXMq+ELkhlV
QxG2R/K9c6/AdA4ewmvYBJGAC9Hq926wZwZ3yOtnJmpLTpKkjkqdCsfCK76Bip+N
kihNzRX8qat8Om5ihZ3P0fe+Ky3ovchO+a2FBkXYGPyzjlYuyMM9M2z1y71zBVWH
W0dCNP+dD0dOdcguK6zrcQ==
`protect END_PROTECTED
