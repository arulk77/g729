`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAxpDIn6YYKtIMQEs4i2qm3DYaBrlDWyWslOYefbsbqJ
MFzuAx+TQ52hOBHs1LdGKh790fCoYgpJDfded+E2sCMpzDOPUlQ0ObH/JulZKFQ8
Gk7WZF9m4xAgwNLvLC3NOJIDjH0wWn0hVkPL1BVMFPB9DSEI+IsiACeE03SUpfzZ
d8xqXzLyuFeqpBSfAYUn9zmsQnFGiGKG/LNkegtlP3AM7QORLG2KYVSTOo2BWG8T
/fHzWvbecXx9dNFAA39DsEmDsSFK6DSohxP4Dhno2M8D2lssi02igJn6tJY7iUg5
B/Y54mtAHc6MIZHF2x8EWmIhcHNZDe3qRZxXZd+H9qJiQUloNMRSghaUaQrX465H
DVZA89vzkcoBco+vt2cM0isOIFiUPi4zn1es4lG99a+6Qzzxq/BI0kIH5NLmR4KS
RnYuKgGeVpL3KWFcmfn/nfwj9ZHVF9FCotLFTXnI92Jz35evPtIP3F7/uDjaPpXz
xDtxqoGevkr+laCAfS8u6YPuAkJRkdwcTsU8iC8//RKPWCnN78Uycyy+aBHlrgZz
oGL9jXppDSaSN1ULdOwAvylVFQWOMdv6vshwlWMuew0w4bLBlR1pcCe/JMM4ZLNx
Yl9TMblUtLChG/IDmElQLTnQcLubmyXE3YHZmW7cAvh2Z1E7HnQcI2TXcNzz0fdv
t4YE6fr2QzbZxqaUExIhfNJL49A69imSxfZIAM5Y4/oR6NkA22RY/zVM+Mjn9mEr
AQ1NaqJM4Odehw5n+apyP74qAxItFARvLl1gwfZ+xAxv8nE1Jt86MQXzxSAuCBe+
eAF42gngJLNeYXQVNqw7/H6SqzAYKNzYHvkmB8PsPms=
`protect END_PROTECTED
