`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+J2sRe1hrQ+m3RwgkZris31Hq1UacNguOBcRvVs3Uzy
8uMNjMLCwoEobqlsxNeE2Y++wkijPciSoM+6n313L0WGPkqgKRCtDj9WcfQ/5YT4
0QPfnX7RKC5FTOc6aEYjya5HDX/34RnCv5MaUJrFqS+83eaahav2d3y9dJvZ2iGx
lmoH0k3eKVKWORk8c8Lat1hz0hAC6Ng1CNmvgVmoID6/aCNUVoaO5ji2soV1al17
ZAtTCLP+HrqAD2Zdc2Uf4SkM48bk50t8ZSAie7dFw7oJoJu/iA1dkl5iaXe0AN8E
+175SPE9mwhe5UJ1ZWFFPQ==
`protect END_PROTECTED
