`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
++fQpixHJ0nmjLetCyhT2nXSK1pCuYWjHAAjxAma2B6gg7rFpzFSlzRaL8yz9Aa9
Zo0pMjQrJbKyzKSW/V/bo3VIhT7asLQXyynC5HNAmOfecc7nD35T6YmX3qoyO4aW
iq9yaxz7jIN36MAeh6g4ZWpjgA70SKhRsp7eo4VlBsYHH5IwYOVCQbI+tpsOSLR3
Lc1fiG0qze6jMXKM8OQ7oxfRVDNUt1AayeUiuB7TAxI1KNq1kNe16FwKGE6k1yT8
QofxCM8NyfTViI34zgeDRBA35S+bBCv6iv6YaQa7mBfQnSqlivyhi2AGYcKm2H4d
289o5edSxC6xu/XSB3/iWAWKQLeHSkkq0LuO79RaPUc8OKds1ohaBranbNtNcLHo
7I5JHNjYMcTuQr/XhX137tz03IYzJ7gNX9AIUIOpzPMff/WOz/fgD8UXUYWiuubF
VoJX8MSczvjUc9WZPhejBG7vjCay7vT3/KyzBpf4XsxoqA21fo/n8YG5foTGi1MP
c7cI046Sex+APANzF21wADmNjMfoM0izV3qTnvz9wtcL6kwXe9GJawvOJEeh6bU1
Vp2IfKR0mLqxFDRt5Wi+7Jo89IHgeqFhMxRPFBwL333xBVmHX8z1K3pfP2Aq+OcU
J4fr+Rb/xb/2CMeOtAZmPvB3clWvjlIJBxu4t3hZ/Ozb5WA3IK9u+5jqK9xszKvA
2YknzBIC4kMVuWPcnRvBbpkaM0ArV7bRroJF/6JDOv2H9ilbidjmNQewRUEn8AXP
JUh25Oym81H7Yh9YFxY46VSq4Yk4Wfg6LQ+9qxMNoSgTluBPGfj8sUEdW/IYHxoj
VduodKA5ImbVm9V7EUyOOBDhJ43Vxjhrv6XWrEfPz6jdeYtpyzBzx2uRCIYf+fhF
N3D0+LmaSj4k/AN6Y2iK0dAJaEMzs11Oq8FykSXGbeH3MhTzs6nGdPiDH7S4+wzG
DAVqoIbzHzfNp/hfZMqpdoHUJlC9RdN0+W4/ueVPu+XDiyX/858Eipa5eG7zR1w+
e4YDRSFlMA8U+hV3YMDyE1EKLSHCxYEtYhsPVBGbtbtKv/j1am6U0zyIEp1COHrY
4CZpY057Rv1UZgb7G0Llsd0Ia782OZJQHQMn2qsfXVGw+OT7xTkuH6/5HMuyZ3KR
KRSS5/GDPDtjSBUyrv8s7De/TlaH3Ro6EPCKmrZ7CQD8gLBZfJDPK5WfEGbsr0hF
L2OvOvLdLdCq/A4wFZttJoxShDSYp6tIYjtTGdXNhMhEam1yGnNPBneUxl1Yk9nB
2P83uVcwZFh48mOGt3LQtrdopbnASwEiyZbEzRc0W3k5FQEwhpk4iFIHITHGuKS1
VTQD867sq+DXFNyDTlp9z/gm5R3PDmcXiom/0YuYsgqdT9YBZtAA4AHXXVxGBf+J
TiOoYyBb3Up1CSmM/YT3+v58hUvNbic3q3MusbNtsUc53+9g6h2qZSgximIKxXuR
BB7c6CAGFeug0PJtasmeQdDD2JRv1+gbp7h9DKb5N+C9TptMnTl2DIG0KQjEgEzr
nVECUYlZ2SREDsJyLTEEIYNBlbkwVzHnd68Ev0cSdVLBQcdcla1Hpitp6kAffuMj
UF1O40/8R4D4T0VcGxMUa65R4koz0Z9BzEVC5SZS/xbacedu4A2RPsd0NZ4NgGr+
s8ecHA5Rs0rT6RwaLB5GeAeZ06NWuc0n1z1a6/3Nh9I7C3mt0Jud6WLUwRvZhelb
3vI0b0MJ6/b3+1FdMLdNygfSFNaBSWezhkRzEBb+fvsuQ0ZsqUQKUZ3EM+7VIVn9
7bREp/9sWPHtXX2CGB7mAwywqN9SYSgOtCavI8jMUF5fx8lt5Qb/69pMZk9ofAA/
V4DS5r5GUgade5ykKs/3cNJPPZTNNP29NrXcELz+2jmQ+YBQW9Q59a1XKGZ7fMjF
xDppaloy9mNQ8OG7Vty/kcwDI8PL/bOF4WPjWHteDZZx9iQ0+1ucaFvQD14LMRxG
LFO6UJKeYkGyHM/mQeHZtgAs4gVsFjL/PvghiPl3RM7Em7Fd/FhlHqdoXEz7Gl0Z
Z8+0vJETmS79U0lZGFQd9avFOT/5p5CkyNBhKtrVEIRhL9FxjWo6QyexFqMHo0GX
QWIU31sd7LRMHw0n22RhrOnK391MeI20uN2cW4F0DSF0nurh/LV6HWFZbrEHt6V2
CMqMIrAD3kT/mZtwQSHY72LshgFT+PzyfCEEJEGc76CrNsDRDCEp3YhQF0/RAijF
UHnzTzGg2nx2RmEBOdnXSL8C9oolNK/XJaFqdKQiPoselqLcHo4AcobzQ6oIELHt
AAo/M1vdzGFsgUW6++fZDNTdmVJjnPpxL34YVeQPQik7TxuKDkoGbRMMVY+IXdGz
YQ95gUWcf/WKNTmcLzLSCNCH3lsPb4IThjYhch7dNQFEwuM8yv1C7P3zXDggdRdP
`protect END_PROTECTED
