`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
BrG6aInmHyQbERk0nVApsfCQ4GFk1ma/QNgROAtuBypmuJqRtzU8PMi+Ywnms5ec
k3MhR5qN+Q+m+kjU7rttFQv26QzKxECpAs2ZFfoKrPCwfanFZTenGu67NySdEx6Y
gO6Zg2MPEtoQrq459Dhp0WlIYqfTTZxo+UJ/etiCTErLa0qVjS/F18frdo/VwnN2
sfiVFJYtOd5yty0vIjBTTXvcwq33RStsJrVCbTXuDZ0=
`protect END_PROTECTED
