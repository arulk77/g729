`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK9qLtUUqrEEieRPoBHJl1hLHGnWQ6/NKRMRjXOfSqQm
rEEU5UCBFVu0doh11lTQz7If9wNywU29HzCRsoojzTsSMNy6Dnw+jq7+rmtBAGT7
Z86rnYCIW/2krvOvuoQfjlELInN7QfR0d5AMzmP2+R4S6OgWKB6yhZL+KWBPGvkP
7SsBTF9SKkspuhFUY3/QXFos74TBGxpBFzJXQS/tyQ6KE40DP7E+u3FFQRMbBMxE
2tu9qwd1+75Gu8cVeGV+iFOLCJBmrAnWKlHBPK0kFxJHvR2eg5KIPBNetzgWypdY
J7aMhnXSQfFP2zw+7Dbw2xvrsoV31pWBBPZQ1cD5i5EyfFk4sucKT4fLqzt+RwCU
AC6Lc6ARyBUV1ucAuqW/zPTlV0SoxVz/kqT9Ilp/gyx2xcGiipWjYdDBr3uVo+ka
4vd6jyMreHfK+Dd8J0iW9oXL/+cAlGa35JP4vKr4tPAWOhw/H+XEJR8+ycweUmY9
7YAKmDwn14VxACaHPXgXzkn/1VGrtMqypu9gJq6Ix3axXu7viZkQtMaUsXCI5q5K
G4nlnSlHBJ7OUUmAj95WzZoVNiDm5P4KrQLvut4TZcWw41FTwS/FPRzzVVidMT3z
zwKgyaG2YhB98XsWLo4rbOgbpwXYCAn55le/aEtujpwSNExJ9KIKUyzSvzbRicN9
C56FBLhqoqXH3WBV/n06e8SX8dcnFV+yOnxkcpNFfkSjcv/TNEymIyrOdIMAffSR
sg5NtZ3yQqt4ZPxoAlOSA95FQ7jmZJhkrf7WjM0YC9teVNbqMdjEOCUieUHrqqaF
si3hU2w699XXA1d6Oiwd926AdmfdSKt+zbPg1ej9yyQkyG/ezjHQMNSCwR7PflUY
lYGO+uGOio2aAGmwXSSFYzNrDpGxdtFFQid7Qxu2VKam6sc1MGM4LnGzpBdOG5Ff
jmNklEsMKGeobDpNQn+85fhBICw1/cCVzrXwXXnivdbg7scb7lLc6WLKXTerxC3Z
hD12dNzso4zHKEhSBypSgql6F8k8YTgCxZngwqiM1tkWSE6q1uqaJ3qpW+062U4Y
+/RA8UjNKUCdNaVh6fNOYksKXQNPdzapTHDkc3VOx/zfSIGGWikUajSK5wBkfuuo
7yc4nwbFGBJkeA2c6iqsjBefpLnkDBDA+E4mtGtSYMvnDaPOwKZ+1k+aXU/RdKY1
7o2CZSLvROjKeNRS7OFF9dVbkZf1eR3nFXQcgXe6hPM8ASomCc0Ho7WjOD2pUTcz
WVL+ZGXPjQMmMAAMAJgRD49YHwoNjQ8alt9W21640nrpkjC1cFpTdYxLBrjRKam8
Imu1hvq6M37WEzHVVzQwGc5j3q8nZK5XzqpqDfJ6YIWvqSySKJme3F8M/uNQt+Sd
wMDqP9nxw4wYrrUXwpRZ1xjmEcJPIR000J7fuHvhz/XkipEVCucc4toHTkt2vjdp
xNmbUWtFqpdPB/WFjZr+61z1pPIjXaAU0XjjOJFC9xw4akwq3n0xgkQIXAnLaWBG
eKZCd6tlm0wtfwMErCX5eEK3pCd83j2vQEnLIofPZZDJnw0SI8VM0/jKmjvcF5R7
ahj5s8HbclsYeXWaJyGKtXloo0wVXHZWzHvB62l/DmGf9hyNS7SkKDUO+Qc+ZQS8
UPX3cFv2tDU7Ad15nePr9TBGaxKaYes00PK3HZOR9HipyHZ/LfEKQVv4VlmP7iKz
dcIpjedkFOjRIE8lmErQJwDNDMqpkseIinsYzmp3tQJ77sGM3YckV9VCLFxqjqcu
+yBELF/t4MYr8nUDzDh6J/hM6P6yykllDTYx+q95cddyC0aTn+bB4gvxuPjFQEMN
cVblkLmpW+5eS4Zx4jnEfOhVEHgPc3CKpwiAh/VXp4+ufYFEcMDccImSV2ax68vR
ksOJX6exbQrXdwlXUvyyKJbbNKSMpHLR3DDFl5eGo+vC9mhdSzzPPrtBYjQoUNCk
s5B4lES3uXEwV+m0d9IomTaeXlgOGHezQjLhr/mY/WLTvcPoYjP6WKEq8JAgl907
yO3tU6MDLHJLXLGBec7bBQmsn0XyLtJ3QT0VXUf/a05xAWjGJ8FxustrIij9l0fa
AWN6kYJzAaWhUadmIgvXth+ZE53q8jtyvwrJQi366s0/hk69xx6jh1CV9OqNleEk
OzWDrZTCPcJjjRjnapmXhHutUlMhp09a6rJaO1xIMyztPRzZVm/U5WBZMeQhRbXf
7lUv4oCygm0QUlyCOAWlP6fDcivaTX7xFFl00PIePnI3JORanaFq+AoKNEXxk+WW
QYfqs66NQHzgDrppaYfnGRVJE6GDXSPiXpfnCABKJaL8G8SAaIfRD+PhFnEtjx0b
Ms571PWZrI3wba+RJaUFLvlXAcorWZq5iXjI3t0rX2Z+IXZv4PkzGv3smr1cCZmn
VU0QBDBkIhYJMfqNkG51sRmDuvxub9WG62UprIGjhUIWh+GBF1/ibVHyWpWyvrCk
JCeYrmUGnhNgE8cwaW84/8KpBA/raO79WOYqWF33NCheYD22vWf5YTpMZsZWwL+n
EXYNpi+TVDwz+N8ajLzXxN34xZ4TVkUmwGP+CoPQr4a3QthSg6MQfiOuM0+I+pv2
/eU6be+uCMGWrlaWJF8T5jz0x2QRck+yi41Q8DtqQ46Eqo3KSTLqWH2O0POGi/0w
lILd5C8Sbuz1xHDgDruAilDubP2/i6pcSUXgw9OhiM4d/EEilSO7Or0h0F/UNvye
+Xr7uoMcDv07CiJx0cnLtxnqdZPJYWhuvCfDpDFDLGGykRDxtqJIzTlIKq42UmgR
H/fpZZf9mKe3oQwPnj+U3FqteG0dhqy0yLtkJKHEq/Et2T8nl38SEh6rhDA0NMOf
zskL0hZMeVfRKYFAfPoqVD/MDVb1yhclboNW3cb8G5pJIYgV2klAh6wK9EjBH1nU
KG3AEv/CFuVaKhv3GlXJykOhiumGwlmb6DYub3pzVmp6yNKdSPBSs+W0V7b/R0Pd
ZZujhO6DZEy5rQmt4JNlSwjSzTWFuXMKJAIXOwPwu4f+xlrdAAoMEWlkbVRZ2Dy9
9O5HScyaKfJJtGBnV25ft0KoiAMyx5OPP3nxhPzKdZY6X2Ynyx7GlVbX+Jo9dHCq
c7vh03lIsMp0iyANIrXWd6bIE1HfdScrQlecy+rRDhmH22PgDxCmt+h7QY1bv1d3
IQmEKZwcnenPkvtMMiMgZ/AeCN+Sp94RUgSfsGPA/wrLSi6MPrRVd5lS+dBS0zVI
whAf1dhs0mfDT5tYuR+VG0q6L50AQjrAcl6/SS1CuwdWwaohY+2ME3DFDJeHRipL
9OcaWGJb1L4h3lfxZCSWOr4ZtxY2l2BnX38SjQBUEt07HUk65Qp4CORUYPt4O3Z1
cStMZe9L1ImVuz3lm11sibgsIHkJe4PZFgjggY+DD2G17NPvHXeGcv7rV5E9cH9X
ZJUIkQ9gG3Y8r9GIzYt9FrpeJfoZdPP9kc/MJcwkk0E+vtg9oOpGM7wRw2231/ao
Ui38E8denOkeLXYlWYpvMeEMd1ZacdMoWDg4/R0ujHegrd8SUjPAjIycMVJLoIZg
cJyI9z0T4NrkLKDHR06kBj0SWXVlrpKky/U1v4Rk2yYMvvhcaT1x7vL5LSsBygAg
7+T2jX3xGsrscDVYn6o5LDlduNnVXIRem5CLrxv8zZsbm67/wPtvflKmim5AKG0K
4WQpJ2yNiBbMCPD+hH8v7iw7tkTvIbC9NBhuhHcUV1sIxgBMA42GzMT8/yQNlHKj
4XJ2DoW32y3eWXMtoYx4/7lNildELFjb2au5vhPNBRK8BSSpjN0aC1a6aDqNSm03
s1qLbsbRQea7yUUPrjlHJRXeXjltgbtw37jqozcnw+46mUkHhn3H79/TXbMg9HGJ
ybbaFNPjz7OMJHR1MeRGeTswjnn7WGaz8LS6jszsVTfJYPBH70cAc0VJfoTOYAZH
qUTrZdi9phrsnj/H7QF0R+w4J8f6MJJgsNT3uQiLB/XbBLM9nxyriLkhSmTxG5L2
2Ri+rswpntpDWqPEU/IOIqckls6WxR++m6794yWxRYTlDXqBmtBCmH97UOEKKQtH
ZhgDXCTvTyN52m7S6PJOtFJUBcZC86vcULIeCMX+W4cXYXtZp8KscCQ4dRLXB0S9
AyhxR+xzL8AtsTf5UFiA4/i+MivQ6TPGqm/Zf5nSX5nomKwv6x/Ra25QSRSdKl/k
8Af75lxpz9xJWAtjuElBw05uSDZAi/ANhN44+qBfOo1PlDs/fySgA9NwES5KztV4
DA7KCR/UdfzFbgPkPbPHGiu1A+jzcduyRcLg/xeLlgveJwK/SVo1LywITiH6JJSI
k2h4AJ98n/+Kri/t1Lh+bHE0yPCYTJNwX+s3mFByZwZe5uGtG68NVhk2QKgNr4eV
G9UHrb0ijIEEg45BP6RFOR4jLot2oiSCtYMWt8rcWj6xVB83qDQr+rqxNwWd9Ly1
Ft0rtbjUnlEDP6aJY6dNyfzR3jmt7fa6z8I3zDIdKF+d1a6teyzy9mN/7ghtPplt
yv8Ur3oRfhVQXb7EwpSTDv0s4xxkFAHqufuIuwKry2LGul+2JvFmNoRe0ThE2Ah0
5bRuuz+oyaipb+qrCqt+CC2UtLjakL/R0sL/NnqZMpLMqeVia5ltyDBSQmTCNxjn
0PmRfOJU4MoCIC8P9u+Y6TWY22zQfTT/CSY+wIB/fJYxQGIWcYvX2LM+w4zFCBcd
8i1Szp2SehP1auMH+WalqkVArHFyds88N2sOdzODJ3c9Yr7f3jG5kYJ9FLxsPkmq
LDy2xa1PRODWuFqKeRcTbODkC+B1afAGy5rTsybwMN4xPBMVSxK+VCsoZAmNVumn
Z4HqKdr2fS4ycDLak6ee9qfSDSzxUenGx+yYqUIuILbvuzYQn/lKixx7Ku59oaRO
8aiTJJHPi2Mpp8+nu+yaEXcQ0JonlvSSxVsmvq5rlgM3jzkVSJY/mUytAQZVxSQG
agEIlPXWR7Rqxf1d/PC/8tUoerfJkI0iEyZ/yKA7bU+igyjin+mJD/B1e7h/+Xes
J/Hw0BneE0FY4B5+0xBI9TDpI47+BJ1vvRLhP0VjeBbs59YrfpNvavVyFNJCnyQQ
Bp/eIwVsta282woUe4E9D9g4WuXLC1CCu5tGjuDXzIZjat2IudLn+EkfT22qTruw
umnbq0PbV+EHl7HgErdVz+XedtBcBJfd4WO8oZx1nHMmZnnMCDl3HkdYyBFnKxd/
2ynABz2InR9W0LYPTGKlRRlG8avLcnp+39QopCCtGWAaDUYzlK/x30ZE9Gj8Gr6Z
MyAaFsM9PSSLPIsDEh4jWZhNl5NnfQ3TnjfkadNawtZS9Rx1DR+pnBSrw1+w5Mnf
NYzX9RebFQoUd6aOL4McvSGePB8FzqWHu/Z1QM/pj3K969W5IMrTqFmp01sMcy5b
Tl2DOv2Cx8ahA84++qqc1ZDb3SZn0Lcc2q3HDrl1/uzpZN60bDAd+4eGe2vrabpZ
AgjOuaFF3bhnpinl67FLvnqt/waSsnOKctNqCZwhEkChRQTYSXrBh475+Qlsoe+k
7X1WL98eeebRSTU+OkAfxnbT9ugoJHyT1ItDyYILBk1pFv4Ee0ZT3UTAG5lKzLWD
7Cq29+hCFautURkmLCv727EogdLd2JmV/JbXwFS6Zk52FOBjlVUYRPAI6qnIP9Ua
MGtt2K4a/+6ZpYi79d8AFGYmjxPj1vyiBOxU7yOBWgIOaSbli31aNOFpJiK2DlCf
TcS1oRrZmILJsNp+hQdRQlVWVAII8A5l9S3m72HiihAqLqNDlTQgLQQ8G9Mb1WsK
o4GcZI9eqapz8UUMiMal2CDZbt6MnieND4Id6WzVPd8tRH7UYYrO3LB9AQ1v+4OX
EG9TM663wdvlVT8D6Obu65BF4xX1zErvF2Vc/9YwMrfs6FNlor8h3hvPkc9xsHzX
0D4BWeKJlVyAdsxfXEs30LHbvYowzFKL6moZu37c00qHXCEJaoIQ5a8msdJA0/uS
eefTlVVi+gRErBlMofCv0bQOu13y2IOeeK3N2cvKXa0kV6dcGX82v+ErMD2M5t8N
bZH5VgTc3G3SvP5tZ5LCJwHdsMuscA71PLaY63Ut7gnwSWde9qniJfV7NWZtq2j+
ALT6aYsjuci29oUJIznvNWQnyCzOH9bzwx809QydsyWWyMY9tTFjdoPEF7c6Euct
w6haFuMvPdmERW65XuuvltmGXFiLejrGs5zXIpTJ/KnlgU8/hTpCldYQ75rXacn9
RfnUptqa9eo/SS1sOxwn+ymQx1ZyQFhvpu24jp76mMLL933wcN6Db+UmxQyJa3Nh
YqnQp0NfE3VLdy0pbCk9/Ax+wb90SmwKPVoiLCtm79Jp5sEC8AjokWUyE7BWrjrP
5DRBXb+mX00LXwBJ3BWJSPqqMeeeTVKwB0cUliPIjVjbT94bAzdn4YMZxzJ/ico8
yhVM/wVEitQLM4RyFxGAOdHdhhE9Lq1OrwWZOEegZ+SC7ElaoSFW6xrtDCCambwB
H6oKmSr90CC1B1AonJoJA6WWLyy1Giga3aSueGCcouYXo2aELN59wOqin6yEFtHj
rug0+r5nhT/rOE4ghiz2MIW6+ivM2+HIQxlS55cfaAIWtIx1xkcz/ot+u9lPi/Af
dacxFXhXclSeyREwKozOg92pt9LqA9ggitWBexZlQmx66T67714B7vAdz3EQTFWY
J/EBG6SLyUi9KVmT6+sUHHFqwkWEFufqF6wIqJk3lG/U/N2t53Zs+rwmWoVrRLbO
wylb3irXUQ9NzE3sXxB0swTNHwAIBTXeZJzYGxKxOb6SfvisQqHFqzdzn5VbSBQ2
haRtKcQWEdCQOsuldVR+1XpM655/Gt3gDDxpSdBsyiLlQmZAShWaiSfr9AMp5LXj
HkyQG/ygddp6ivb/JF5f6T7m5qxZkProw8HfiTDdSS1apHOHIUz3qJUyzTa0c5S5
SiCuygsDBWQM8uiuZYU5/Arbl3Fo/6oohzsUfHqG0ldH7FM/mlPIJL+pBbGcUY8/
OT7/5LN6+IdIq9iEBCXH7WgXRcBtDf+l3oa1tPHrmlrRW6LtdVIYLgwFYMMt/BGf
M8KADG8t2c98eRqouhgbT+zLLVdZ8ovkgqQe/ILu+FsNIFpqOGmNcijJflCtyp4v
joVVi8tbNxHPjDHKE/Jj3Prn+SZUgr5/iRw4nEDF7JyktKcn3ZdtxqTho6OyLHhv
Pz8Iqh9oDvFC2kCQk0vSJE11IlrInTWYZTa7yc+3bSjbM5uEacbArhTDaOE768CG
RaaXQao4iyCoIhAWh5JTUxghK/iI065F4Qz4hHq/wS4oPjt1nV6+6o61vQhPKXE2
sqLQgrife38RjxYQut9jHWiZ2vz3Ty4CF+QNvgLxbztlaaJ9r6jg/eYN+tjmrghk
q2nN/YndbNnjkQElYXjWcdx5OqXAduG8Z2vEg2azxsVbQyrz6n7LPJ50X9heurp0
6xyovmoUzitJaV9hj9ntEz5H4J51bV1saERFG2Kfn7OZtw+pFu9AlxSwITQefZ8U
nWpcZG4va+sMZt9aDwaDO7Pvg50ii/ISR9C2jKmAMtj78kqNshfTUTiShxMi3GNZ
bU10zY/gvpy/x6FN7PSh606Ej/9j1yq8Ib5v14Hd77TEpn3fq6GxTBaxjdTBSH8t
gMppksV069PkrawYRURh+ZOO1KrK5USldSdiSs7Xj9e7xIkZp3Lvjp2uicGas9fI
+Dv8chkvO+pnmtLt5sBi+nxa8b0wqGNqjr9IvGmcRT+bDlgLbzo4qzdpmwVv9meh
HqLUqja45tFLWdsExDUSL+xEJDFw4iiefOcWbPzrBUsaLRvHSEHCqA1uUK2uKTvn
5GtdTBjUTEqNMARpMlLzXbbDnEsJhAvrN+K9B52r+GCPv5G4s7R+LCg/7QjVIsvr
2UvRx/n2djZ1lylUIYdapfgjyScbIFjvnqGp8w/VBeFy35x1gzrue4sbRwZY8tUU
j9iVk8Gs3lgCk0GlcrMhv5VaGUxhw9znymM2OKwZUgox9fyflOu+6U+Pck+3X2sl
3tZznDoXXjC3zS7FXIvrCpXSH7FUw2+2ZL7kJFMJ8kN4eQbfxKVGu9cTQNhXfKSi
0/Tm7lNcG2g76jx8j0shz7dhXiVqJnYv66YobZ15bO2QCfzBEoZUxxYWOEmzwhNE
i1FSzEJt7ID5CWC8unqA8iGM2vK6baSfO/QgAHv9HXCwEBao+oWmLgA/FlgR52nf
diCyiNniUvDSOr/UNM41pAVGEhncAkoO0MFYA7jvUnr/FHDXvEYrMewIH16O2i25
CQY7zSu4/Rs2tlIjm4vNfNBjebM3pHTAdARKrZW/RoYGquf2sjq1hYKqhxUlY4jD
iMGVfbmKetuWbsy6n1muInXfy/ArY6uBO+u082iArFQbiMkRhwxHyKBAGwO7+cFX
UN6mRiOeltK2wEBHsRhpkWLGSOsGhXDnnysQHjKs7N1l7DSe5XBF9NltJbKRdjrm
+vjUjb1YSB6ZhEOrh827eWHVk8mf9D4gS2fzXx8kt4ldM2gcL/fiK3++/VXXP0/A
l4TQ2riHpvBrxHR6gEOTU/DwyRMs/mhC8y1c/c+yYVaOoEYJ4vLpSdsMq0pu92qd
CuMlOUSUZXo35GFYhLcpFH7/nBjGnOZRTLCMAV7wYduCRUjM8Kn9n6PZrEkz190Q
LTELDISC3/awX/4bMaR/JpwC3yf2rK1Mp7GDA2ygOgq5XsCL86ezWhATHBlazfMT
IyAaUsFnrTLHn3nV5hpyBwy0mJiDcCgUVXYYgfvdvp4YfXnITx4ZM3MrYFVk6oOW
rth09++oZ8t+y0D6Lkt7N5oC2UzpxLGFJQjLCY/cHSqQ+kE3vfSk3TKG4nRFtHKZ
HAKYtQEzmh78Wc8Ksya8fcPq91l8+nR3Fp/ayRhGfb9Ogytj6PZtxMZCNktAFBc5
kTahr37pf3BLz1OpZ1rxGcXRc3t5OvLYWRH0/GwrYuuTWFuqEdTwBQzVy3vlCdA4
hJfNJ9fQlSNi03qzWQYV1mt1R1uHaEm8DmbhwnWOZygHhNqRJbCdSKY0XFHhgYEj
din7hD4ZV6Ou7zNJlF98hnD6uuWAbvZw67EIHpnnOaHOXTLM2cHs6KnQHkwCxOwE
jje89vC3cJeUdryhB291OuQxt/LLkuK1ul1pDqMGt/4zgl7q5no6ghCatWqCcOhS
qEgeU7Bb9m34oH2dcCPjdwOnDZBL5RWnvEZo7tZVHaFZCM8sp/umQnyRAcXgR96s
RGeqFmyb02iOE8qnGspKOyCVpAy/JySb2aT+E6lp0+/LQO2N1xPnedOpdgpglzq2
hbbbwBrnGP1ZGS4ttpecYOGcXbnO4MU7dRyfe99SuXJrHp0B7ld7BRsRTIs+A19M
YLtWYxyc4lCMUD1hW9ewO19TFpY1lDRhBFQuxkLzJDoHpOpnE7MocFH5wR1UIPc0
ZmLjNQK+B+A/rK66lmPKllKMTGlsvnTYqj4InkiUehwcM3GagdqvVSMy3HLeIArM
pv2Ka+toQyegC+Yo9EpXoOwT5rXCtmzrDH6uZfjGggD+wDvzxfYz4BRghsu9BKUq
eQYIZA392VrOJB3bEs1nOaeMCdFv+6L8N0twYCdh1aFAaFsctsjrhlGbRWVYqjYI
Av/+Po3URDXdRc97JlFwtli2dnGxVmBXLB/J6XWmVCbbE9i3ktFMKSElMOt/fZfF
R9Gst1ze7R6XhmsgYBeRTEpYt+Z06iSWaPrbCDI8/vH7LdQvEAQ8tIqql0t3nnUO
nVScPFbcVPw0stC2YWszmJH7INeOQWnuQrb2Me+AeCdoZ/uJJXrjWQ8i617aGV3t
OuCvsHsIW/e0+GjyR5b5SjGwxUfTzCStc72Q75ybBPJ7TELSYRH3EDPF7Zs3pHiB
yzrMJFTCqojiwTq9gtERqhAPtxbZ0Uu1Aun1khucI/BDWYnSke5JkIl5ux7faak3
0TgQRAmVFbcrSJUlMfFT0n2JsED5YZsdZ0+/kWwHznbSgjFp3GP+nh/vvb7LKcPH
Ot/vPVv+6+O+0v8qY2tcG0CfFKpSXtFgHRJtYe68QFCoJFW1wSgOwVVIfIF3DKAT
POSMJhZnhDsOD6bFbe6Nr1C+S0zhIYlyatjGvcoBY+OUT5wDNLCCk+6XVYR+Jbn3
qF9IeyOlO34d6+6zUQm4yZhiqgxDqlPxMIE76oPGAaDEANSAOmDgI3zuJE8/sVXC
eTNUNTusp2o+c19jteivXlF85ggWlIa46BpHZAcIqZ3y8l7ARkaKYEnYIzoMkpSl
s0lSbbDSfl8TUrQTxf4BYBWNVVV/DSJDdKXRHTupRTpXeCTic6AkVskE6GMj92VQ
fVSL+W2IQgORlbHzitawoBtwNlxZLfGMDQJsAV6TTUBSmix/BK6m8T9lwKsP7TN/
ByJa4mHe+xvlAgzaJUNbF6BjMtY4nXneZ8nBgp1ML0vHM3LUTLfbC9tcKVxw7E4z
cFPTmOtW6uRwFRIPEd39oxZRrHBhFNBdHbrn4pcbG7cEgCy/OHKKPdYBVIlalITa
HsPYCYZq/10Cbw4SvKUcszxm09EJF6gA/fttYYV/Rtiym4WUmf4c8Dn5QilQ9TnM
WdazOitCVHxkorLYuT8/S7nI5JWQ5xD8Ov3C5SFb83h37l/JC2IfZqojvsGZPrAV
3Lmg2/L0FFoKCVWxOBNYHRtfZ/CPFcJ11v61Oqr8FGAx1wS1LIj0ZaAMJ6/lunWr
vA9g+9LR/1KCMtSNoDjut/UHCHvkfQNKtfK4upFCtKTUBBddEhrbarUliQGM+wZ9
V2Un8fHWVWGaLJVyzKg4osswnZuDQF2fQb3lc6zut42jHTYJzQEfO7EgALVQtkYR
WP3HZqilOOLPUX1dXaQyQHJvVquhwwTV9LplplMd1an0c4JqVY5o9zksXk86ik2Y
ZfSyhFnSLXrx+zWuvpjnDJiGX/aKhuSyEuzdi7a+4FnsnL6kVfLbZ9PoMLMtK4LV
2l8Bf1qcTe/DKFrokZozSBojuoS1KOa8vSfWHEvOufV2h+PjAQzqxrlfNpGlEt8K
sFn/xwHF4DBc4BqSHQe/o51o1CE01/oWqixuJuGV96pPEfbHyx8oJhKL6HBm6ggH
CsTRpYKq/FidW/mvZ8Hv/FRx1W/9KN8w1dhqRyz+KjcV/ZtX066YQdeK5P/Slih3
CXWRgj/xxHopFq9JJAMB8cgMrzCFKmJUeJYNGfDEW0rxm9lwkhnwyA8+AM3iwUyT
s9C3XScJrWhCTGcCfMCsEdA9GDKo3+X2JTFurXg4W4oT1odfraghp6rDBkiS2iep
XMlTzcVLPvqRCG7QJ4SO1fgwsrEMZkGTPutDhj8uYbNtj4M28ohPplR/+eLdMknw
cRrJZzdn3/lrS043xG7938rATToKgpzZZkZGXEUYhEKykVXZjCPptqlWnjlznAUu
GgpiIZY5r1tHKSVBA3eSU3E40zQR4MAkiUcf2ENb5PTSHH6ziz1VPJ+7bsSMedL6
bANwE6ESyZIpbzdUlTJl//ZmEq30K7m1RuzM3eO0aPKIa+2UBjtZYwrQ9Pr5rGo7
/3cNBaEAJSDhKBa84mxEIV38PQxK3TEuLtVGShKOiOEq8oenN/FdL3huVNRnrTL7
a9oPps1ZWkJOvt7Dl8jLWEuMZMbOoJ9QQ5O4WsRw/wO/R/P95aWcafqm7fc7wK1W
3LXK6cOu5g6d9p6d6bpLYuJ900s2ad6jkhpsjNwU4/vvCFemGsMGYKYJ9wmrJ26w
flrUi8GZnQ+WOCfmafeKyDNRptChJRbzhRulhu+ytLAytXQZwwVnCg//TZikn4Ug
OGTO3j8Rs5Y/YfUWUstsleykV1UvJkphS9DQ2FeEQf5sb+uGyyYsRsO0DQEGMq+P
BUR49EcjFJ6vqdZ0vcVKqanc1s32jwP6w9nARzJSTht/ybA1rokrS8Js4933D5Nd
tj0AUm9hpjjFuZq40lPBJmQ7ji0ZMsOkz+V05UkF0KHzt15/ThnCXJ0MyWVvRKiK
wLMffMu5LCWLvDaB6KEcOPJNJ8WTw0Tyt5mHGI8qJzJmsOrsH+8BTeYLwcTk7zpz
ZxGtFfj6r++ghAeGwiJrnQsbOE3LyNvzXhUabZaE7RGmGybxaHtpIaqHItF2xAEc
OLVtwYCeuY8LcD/H0pv6BYSnQ/LfsDVnnxOlc6jFaGJDFe0MRJlVVD0DC9fSyJln
TnHKZLS1/GriCaNHSqgf9L8S7doZ6XsO2k5zDBtmFYm1A2WzyJKNYUvy4J6pHhs2
ig+AWPsKdvlzqRMHrFJdttgc7eaawJPSSkWAEuWS9pE7ds7FAzj5Fjcbr0xiCaSZ
MhmYM8ikvCoxPm5DKD6ayYB9YrjdURrWAhnG0d+rv+2mHfueCVoasc2pxCFf1T4O
xMGLVc4bh0Ajcuj4+yFEDSlBkgRPYo/mvXLepZ3EsiWWA1wyhRM1eKqvx4J0VcpU
0ttEolwylYFaQwPUFL7Hz+c+/h+tyG69dWXEd4zCuCdvl5gAWGA6ylfNbRpQUlGj
HwwA4p1XkFyYYzwx+q9gW7ZD1SzyfOs1ECUlzbaER/zkj7PAa0eYC60DkmlDDfWk
pVN4TisrHD3SNcyqazRXO3yc9e3e3kJkk5dCNv4/QYFE0KU/L0HAVPtbf9aOxoAK
lDSGA18G65XHpklgBK7/f+qic+6y143gKv1HpW70+9nphl5nYunVLfvxdQ07PriR
1qnGffo+nLSCODOfB/vIZs2Gr6loiOgaR4SFxPuVMZIsiadGEakmmI9o0HHJ+1A4
SQddXoj0sarqiZLjP71dtYu17MvdR8rq3hxyykIgvRRSDWaVeM6FVKPO0Ejl6XN1
sEK5577SEmG5EE7WQTYI8wFa80MmqBD/GLwTjcMrd3ty5JrSeD3f3wEGohAeuFDj
Eq3OQF/fx07mShhwtc/2kiiBzjkm/Vm3tYq2Jj2rB/sTckOtzPznwRAr0EvA2z+6
0z+KhWkaVFjUbvHHltBtjzI42k+0hJnbzP4SMqNhlc8OVg2SFe3APCVTceF/bMsT
2mDS26OQySP9/ROd0A691l9QKVljeRiRMOLlfUlgKvS8K0w/HDry+mihrovvzR0w
3idNYUXWeEIsDeobPLmQbaQ76wp7KserTu897pkFulLs7RK5c3DM5Br8ZaIT7OvC
O8euorU937yJNtV98Rt9LjdRP2y5OAoc1zdDWC9deAxcXGC0qbwHGcDpYSqrbTQF
CIW6gBi3Z+kSQS/Jgd7oIpIMQhJtHk1wiEKFBK/zrPy1whPsTXhsG+X91vYpmtLs
R1c2ywUFxMeRj7PcQPCAS4NZtO8CWnPvHGiLyatRdHh3PgHtWqjAOll9uhLeYjcA
xVfqlNgm0HD09TnwvRJJO/ZRjDm9LV3asSkULR2HF4mVKoew8QloXe9o7/ZFLnaI
R/zEG8iEyLxRnfBqyBkVZgB54MvtkNt3k6Y1wbO45zO+BMTJVyGCTZi9tmK7GIny
6a2RgJMukU5xVawCZz//GokW/Ra3BXWlMPuTzrqdtrIHeGxSmNSEOl3WIDdb7J31
iXKLbDhZtfxNlESmDtNPqavLdWVOnWe5EpTzyKUgO0ZxG6YxocbvF6e4lgokMKFH
5vm7aCwnXjGBhUdXWuM8MUjvuXnNDew7JGAyRfA9iRlz6cRW4nfZQ8MFfyr8unf9
gsf/ZM8HBVnvJPb7RThsFmW3PKKNuw1p44RHWzfWtM+y2PVWv5PRFZVrtNiarEIy
lq3DAh2/ojlUTK8CnBGPzG6cROwyPUQkKmrAiMCa1mX8LykkEC3+f8lDeSialgKK
LH8h+5789YiTFu1S0OV/LtO3SbIWBNkkQeb2+ZqMNE2g0z85H9oZS0lTU0Uxoa0O
OCM/db70SyvO736ny5Nrl2Fk7l956kWanFznmCAz+b0MqIRgj49U25mTPQFkWbus
1GMzPBMrZ9jZvYJJc2k07ZIp7yH6OTbaFmS/tD+QBSC1Zh5EjlyOx9vHWaXFpSVv
i78UPSR3ed6h+y1Y/KcOecqyhpwqGwRzwCOvVRoEgDhH1o4ImgWz0EcT0DjkkD/U
RmQ5uxttjct0V5TMYt66UE/4hglBuE4EhiNOExoxrnynPA1QTI9ISmkTQaXCUMGt
L0LIRXj3vbWJZO3ZaBFEn5DU4GN75StA8UjIWtHs6cuuKcQuzXJgOarAp0MkhNVU
rVhrK5p3jGqlLJ4Ch/TEPNakCI4NMjln5cMbmY9rso6YYiDHyUXoFpxuIRWxaRcf
IK73ypaPM4k/h2PYzyl1F//bd897Z9mBOrX9ZrGrvwtj7n3gLTEpqiR0hNijl4uV
Q+35N7OmzuCaZyzgVOLpB5Tfr8V3Y/xMKvV3akXK85yDp3ZqtyFGZk5c2KGkGPk8
DSgWpWjYy71XRbbK9frZLoeEy+YDdlcnxax7OJ9utDPDQomTyaDOkXRDt5ZNHiz3
FjatGuCICAWL4mA8hn8ATgT4FDAuIsrwa5NFxWX+cFRsrW9qQ9sn+WUGXbZ9RfO5
/iyVZ4A9Jt6bZspqsaKCGAAZZYhCc/05J+sXu2wNtg8eArRP4nE1+8+iszLJUM/e
1L2HA0Rnl5LxEP+CrcnXN6CP9PqzVoMvDW1FUm9zqLRRT3KI5fEdkOKcIb7PBTtb
0PnCkr5dCrwljN4bGo51vjBbFJyZMqVq1cCFk2KFi2VfqEPzmUea7v2WkDYp0BrG
YtLS+IVMHwRFeCxWpyN7ViDD4C9a3sogkLdyUOk+hOHD9V1we6o6v1YDYfmxSThp
BOyPCDpqD8Ct8MITsl+rLksqa/pnSoTWDDmVeHSBQ7nP9XaKcJCKZZ6rsYjD0Zx9
taj2ldSME1rKCd0tq1nm7dpYaZNfebJra6JcBuue3LdHrAloEdBGwGxtXaomDfr7
mXkIO4RenjDQyjvab1Qi3BZa5T0G3lAKMi2BYqlHUkZyUxbnt5KdM1GHZPTiAKp5
JbDqARM1S+w5DeJ+4sqQ7+hZ65kJdAkFujl0jOpGU4F1hz4RYRJmjdnYzuAlyXIN
MJdl/zEtcbu8k0xEyVZjXXeccCZGs/IlwsAuZOqx1qyFLBMWf2sPELOKzkdrPbiX
iueu4i2vf5G53eGmq8pgQpEXFsIhRYs1kiTVrwOAIG+Na8T64s+5ZLQSHoZGxQyV
221WEJBH/wvKbCJMpnFOB/C78Cc9W2/lYD2yUiBzjTcekUbvWBwaDk6nDZkhXDgH
on5RvEBDlt0nA3/nAJIaCxCg2cvc9YTDDVpwvuRxY3H/73NLtqOJ9XHRK3HJt+nC
EYhLEW57jGOehVi6L7PpGlNv5sRtdrycrcZyIXgKioIRiTteL/A50qoM0I8IRgKC
jfqoMqYbOriwr+BAwoc42pHOanzctWc+7GqWLdbcnDFEJPGK+Njh9L66p5YlFlWQ
b/+HLz0w4n2TzQPgnYeyJH1KdgwfvERt9WWM5ByCTy5Np2nEYOB/ynZphNKJdWp1
LUUfghqg42P9A49J7OlZ6Urr8WUAiQ3vjEPZ48l9++9ou7fOPinaZYGzuklGRJMX
Yl5TGo2FVoNabbCQb6LdILtIbxtBiJxnPtyfSQa/4jbp3l2dr20hPKodDgTM5HzW
UWBtN3F2QoeaalakJdbkci8VBxrd3zjOCPuPGXNiXTZ1sdBcJNJID5luH/BXpVVs
jol2vghUKNmMQlVQU99JwD36vcQD7V9wGBYebRJBJehJy18f4va9ivmiGXiPKvKx
w6jqgYVKR9J0US++jDa2IXCHJ/XTC6HTcdM6TIQ9NHCu50KADCpkZN7bgS038zZU
`protect END_PROTECTED
