`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45nLL8F8bDxDvwcpU23iB351HoKyDJbD92dUk+9P9J6h
cTgLEZ7sqWJSJQ1Msrd4JzsA0seiPfX5FOAn8BkgUWTF2GUn/gXnMPDuGq9kEThL
xbtp6L+3zqeKayIOdwherreUv2MyDz1Vr7rSAKpTWUgmHd/ROndW7V8Rsi2yV9hd
gb4iWOLENJ6YT8s/fSqfTUMkwWbYESQtIYwk4gSZWXQzDfbx+p1t8MD6RRYa34RR
G9VztfMhGEWunQAgr/LWteOlLqv+pAJDn23Qdyx+HM/pm6g9RNVsIMvtnY03yvvR
dkrywXgBHCciYyzzrfD5Qw==
`protect END_PROTECTED
