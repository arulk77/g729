`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
oxKdgxjLm47SHyCLqK4e0NcWbyF7dbwX5kl5sdBjt1sIMkNSt9eeQBBo2+5LLOm8
N2FB2VQF0xZ+qSCWkc/0X1oaW9bBt/gWfznez7KRvQmfJ3Re/b31mWV3IqMc7yxM
jXRmBisy1bEl19AZVaC10q93ERraq+abARhhJTdBHlFNghlIaT5RdQFr7T5cG4FA
7AfoFaAdJ8049wg0pLADWDOuX9kWxLvjBOL3JmvX0do=
`protect END_PROTECTED
