`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47KqYbOgSV7ag4XU82bmQA8AltP3yIAbRa2UOSc3UwJe
WKweTr2/LfXsgFNa3ePUB2qcEe9DpI0X80jjJiu5x+mmV3npQ9GnwU433cFcmnnX
Hyw9/SKPzyb7HpNo5CP46l8x7a7St1jAHDqCJDQtu7k9TyGHp4YVvm7FZ1jhFia8
7W8VnhHVWMFDjem8oTM1uI3ivESkoBuzuQCTGsSv8BWHybJ9PynSxMDwLXZS5Pwm
8bEaMNvZ6zs057rPtZSjcP/CdSm5nPBJ/hhakFQNTnLcgvR73L/4N3DZkrjKPHFx
TAOrX811jRswU7BHKyyOOEFRtM1bRaYH5dw70rxI3YxLLZcxHPkS7qzQj0TBDzfA
iS4rmzKmS2axJszPzE541aB1LljOBk0wHHjGvv7a7iwTFQmj2r1zRn4U78xzfCsZ
BK6I8HRy8t/ck/d49ZAA6A==
`protect END_PROTECTED
