`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFr4ujqyjWrqjgJQt7ataLyO6fNczNauqR3oQVUfQqx8
/XAn979mq4hx7FIUAY7hYUo8eqVvUGrPdM25Pfk+L4rMF7Eb2qr2HSxkpNMC6d6g
uxNdAZ7ZgWgkfDjTKdlB4koHBHe5fsimlnDz8dBs6aUZgLz/SG1enPn0EKS4mvSz
OJhhiLilefYoTALWdvHXxeKAnZbUDTpYMx8DAHGfJFGUW7Gidw94ECCJyXUcUmlh
`protect END_PROTECTED
