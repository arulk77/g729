`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNo2pNc/dBumgOEiK7q3bObL/4yqaFX05VX7m1I2FRce
KXCBoTjDN94anDiLzaQGyAagUhiVUz+nxrhWRceJl6ky4Mbk96ap/NHGULBl5II+
yWUs2bj33WPiroBzA8IwDzDi2v0Ni6H3kF5SADnNGFLlGK2HvM4HsTnucDev5FBI
V9u3aZ6Y+CDEETQVspWWVA==
`protect END_PROTECTED
