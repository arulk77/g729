`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGcWLbuiWXfoLSKcUoWrvPAGH7TlL+pzjst651K/m2vn
g2dIkxZWknisVgMyHXUc8ed9vG5iJYlJiVm2potG3DGZQ6SOkbKFF3GOgIEamgwm
PhR67H0YgYnyote085KYKfjdITAVg9SEmS14YNCwpnd6O3QAWKeKJ8A5lwLnHt6c
oBpvVyqyUWHwfiu8NaPLfoZhUb+/yyvoRzAhWWvIuu0hu2sQdP8JJdVo5lMl2UXe
`protect END_PROTECTED
