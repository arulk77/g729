`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xeyPVqq4g/w4Ky3NdIqL9gWzLuSzWrYbO2OzPL+R4Xw
h60S8RAzHJNUScIrvKRnYN8fL/mKz7O3Lr931RPBC0eT6YxYInzYwOMBzbQv5OCy
umia43+rDFKCJsAvQQDwwvDcxtr06DjoXmAYNcDQvaSD3hEAj1XHvM2byu+2D7aI
6LFkIt/0mDXtuFxPnmCk4pYZsEmSc6NKeqIg5R5A8+3ToajhY5bAdmq/T/NBiNnT
C200P5B5yxFQIvNIuQdlEKHg88oV93VLcyqOFY0SmzTANySq/6W46ha3Hs90Hp/k
8fe1Zu5YY+ygNis5sO5inn/uIxShJXME4l0wxFlQdSC/zEaV69pJT2NwUF225DhR
i/EYxh49RT4MKfrFEriPLaPfQRTlc/JsCgas9hUNCgDc0jpyGlQmfJcS8lG81AY6
HUidX8nOoqvn+f+JFjxN17/1Za3DBU99+RTQ0+FMQ5321JJUVJbWI17p5uu2uzHu
`protect END_PROTECTED
