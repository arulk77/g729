`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+pvvByY3Gc9xqpgIK6CAvI1yVXf6t8yVJbLCY8rElxboeEJ9YsqzIuHEOiLqKvbZ
Pvd7WmDDF5jKSNJ3Mhf3VZ0d2AHsDms9D/kf7OOA9UiiYOWXeZZlNESo4rplUFXO
eMK2OJSk0kMkH+eMZemCKwBe8lkNp/N7tAGfoMqdRF3sXadLLGnfaz7EHHBA6P9c
oymCpjS+vr8CGwx7LtEwfgXGq76eeQKWrW6Ck9OmYXVtyqXO4qk+wk1n0WS8v0W1
gQ9dd942+GyE5lbbb0W5zomz/dM4L123f12l5FXJjllvDsYrao60gXGWYyNJTf+v
yVrt/3hU/cM1c+CurcySCh20PZXeqSRamjPG1KMJxlQ7qcmqCmZYBhbXOwcWEBiM
BH6xcXq/zZygJSFcNb1yeu0VVe/oSyoEwnICjIRPt3felZygEONecWVFaNm4qnhh
R6ggs1Pdf4QiezidqF+fOMW4rXJfJ5DADwqmnKiCvgUyDC7m5nWQLnmDW+QkFkjd
Y8S954waQgw4I/6SwaVMQs8FTa0wgl75d0eWkpf6Bt3iDISdRgliIU4KTljnKBAx
JgnENEMNbQIJozcrAzH3PRgSSlLedoSYUm+J63gqZwtYwIPgW1KArGR14RhAzaM6
S59Hc3H/VPSqWOsQLO8emdcj+A/Cie63zHjYBJFgXwigNx0/y3tcf0UvWm2WYJ1+
eFloISftWCxMfo4xPCHw6qV7OgZaHgPQiHaVFAqB4c6c4Mb0ImFc1fGbaqHGzayp
yoBwZuhFFbZhbHb8FHIPH4eUQJPOdsXxM7w529fD42V5nFIXagJxn0M+VO54IeeB
5qaK5BDiMr6c0uRAH73ShS+WH+vvTqQc6a63jXoRLnH/34Daf5njlB5thuZSn8H4
uilSMFTXAlj+ZUvRnjcU6YDQHAG9E8hVzBBXEllu4QOKhqCqy66ugzYZ+dL7qLOl
KEDD45XJWlgK9F+AEoVEA2acH5K7zl1WmDgcKyiJQeExfNJayC1Knp7HBtix0Tml
t8O4rhRVqsVLvxlt0ODno9P+F6UCY0Hwqwm87D0sBTyV8h0HBw7T0dFyFuM7qwG7
`protect END_PROTECTED
