`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xkCiitGYPPo50gG+A8SFi0zfI1fTj+878rLkogKywOX
Ybt6A1/AAHtYVElpPfX/upDanK4GPYIXVx9+0bfC11Twtd4Ax9m3gqh6/dkfv//t
Cxi9F+TDC5bfNmNJ0uAxXG9tnsSznkTFXQaKqrkfGd38Mwk/Xb4YSs1u0Se8gbgx
UD0gWLPQTTCJaDhLDNth6tH0XePZHO6oL638tAay5noLfsRU/Bs5XIl7345W0W7S
v8kUXsTW4AcBrIWx+iFPLhwY/AXxj9ektJiat8sMNBQ=
`protect END_PROTECTED
