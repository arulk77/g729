`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKtitpvUuhT4TeMXXREcKTiw5j5XDV+44X2wiOo3PU4v
Em9ba3jhVpgUjsRBX9C9+k1zLJKETw/2yYWETHonad2WtIfgpyYYPuNljwjtEejj
sdvMZF1NK+b3NXRtzalXFzcMjlIyHYDG03At1xcU92+6fVVmxDJj9vjitRvOLZoX
`protect END_PROTECTED
