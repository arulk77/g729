`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCQMTx8qURXiA32B0U4HqSjwzoacJClgiuKWNrzOEa3i
mD2DXVSmRtOvsAanic2NEu1j6U83caD6X2YQBRRTKR1xyHjBjIXVpU0vLXvIIO9s
dLS1DKYMctU0lu3lcUbSRdLtekWIuch52tFleI5m+IenWIAqs22DiWRbmedfrMf5
XGBsdljVPbNB3enGZerO9mQVaHMh5fdY+yxfOKcvl8qxscOQ/xFRN+sPvyI6y+l6
weEovXGl//LQg3ahziI+50VMB5qnEF5DkbpaNoEuisdcl5LmHCTKMsq8XRji4bOR
CqZFMDhO1kXt2rH89VkKBY+jmVHWKrXoaePQBH1Pkp0Wz8ZnG5RANkda8ufxjQ6H
mSXfBkq3dZJ2pu2HdZpxUTVL34U5N//QTtUQ6SyIiXlkXSUTJDuwqsvsouDjj9LT
lty76FaBKx8wiG/JvCVr+kPnHUBJnLRRA/YDasgjbOWqV9g490HRBo8XqyW33x6F
OwCr9q4bNvV/TZrMLaYmVwCbecM47K9rd3Ma4R2Wp8Djn+zaJb1MeB6GrnswoAXj
`protect END_PROTECTED
