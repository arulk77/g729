`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNSWdGjrq56tSqB6SVFbEVS1Ui9+UpTo6pazC0oI7jVu
T3qc5dAyi47tjz0BRgl0Q39jlEHYaL9429MdLbqvhmtp14S0pKv27OFbOjz2C/J8
xn+Lcp4SNM0lbianvSbkXO+XAW7M66cs2QmsBHiiZTByLvSvDxMy+s8FQVfpYZ+1
JTVt7vKTLkV4gVJPwB3RmKUt2tR1xBI4yQ1+1JG7dBd48sixSfQ/R+cRuCqtHAyD
Ed6Z+EJTiun4RJd0ra9MvHUQpPrR8icr5nsyjZP9WfyWpXvopJ9dQxIt3JEqxBvn
Sh9tIRje810EdBCxO4yWgiweaVBPgMr/CgOSdNA8xfDSU70IwqMxnkH700x/ak4F
WJzd/GDDSBwr61xH5lMDWkdnrhwKakfXU9ITGIWShH6S0lasRQnrdgwrNldZbsYx
JbRNlYnp2xELGlQbWynDikmF9dgGufnQUsIDhNvVtE3UE9yLm67any6jOGXB82uT
u4KDIHYm1aLHutJtSWabDI0tJxfMacSeILxJNEznZFRYyDaxPrh+vmDQiQH9Cr2C
fdxt7CcOxcoADjoDPC3/jSEh4XvnXDVnGTivHjxtO2I1E/9W5HdVP6MUBcG7JOFo
6oaemXQs1Ml2yHwob4yi9OgMOqrc5dOW5uMh5nuHJV/fDHcrZ4MDqjcHN3/nz5N2
hapDlCXAbrIh1XSp14GTvo4leHgQ4ksCwcZ04zHH/CeD6q38sCKFaJOaH4tMfDwh
`protect END_PROTECTED
