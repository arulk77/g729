`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG+BGyWzXKx0fHRe7T6qjYCpTUF6SVxycTjHmYA61kv+
LlOYXZEFLMM1Ph/QzyCu9bnQuRdrh2YtbKlNFI8yelgZMDaMQB4NTkuGA3CwJbRM
8ksGiv9iLy1+PAPcolTyFcmxhkacCwu6hyxUhE0r+j/JkvZ/SbII9vi5DEJ3oarS
qvqsDSxRv0dOA493dBBEDbFiUulJ7wXEmJjEJDfv9t0Rz/uDEzghKYROyQsLA3w6
`protect END_PROTECTED
