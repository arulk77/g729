`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAKyFN6TX43oqzB6OvChOEIrp4Zs9G6eJU627iVoyH5L
q5L/efeDvb/oJA2EzS867FKHIwiDfK0Jb0KmuLj9As4nXvkDUVxWhjIJYaQnnBlk
PRLZ6ROLXH8sQufYvS/p+Q2taol1L5ZKGt5V68JEQxTCOwmjIdwylbFpsrpreV98
sB+Lf6g8uVGHb6u5+KDzNO+rXiX8KFXNxenZZ0FDP2ZIE86qelt7HFXR0yqbXtDg
polb4EF36yTcFpikb8R3GnGBU2e84iX47y08t9jIEo8tZoTjRedHJ9oQHkRO4gOs
Ab4/XkJj+0wxknhZG9V2ZdL9Tiv+H2vKEle8rC71AbwGzAPwt98toV7JPxhpEvzX
`protect END_PROTECTED
