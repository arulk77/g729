`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJb7j4YlMniDMt/doMp0zXEJxOnm1DltzFj/9GJOVVHe
16vKg5l8chkZSX1933rGiSE7JM2XAFX+DJIYw/UbwSLlt14BZcEzH+f2/BVpeqHK
+gEtO0T5/0nHQqjEBnHHZ4QjR0e/VAaGk3jogdOAn045F2ilvNySIhjIJ95bnYpE
`protect END_PROTECTED
