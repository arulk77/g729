`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN0D9qcVUJ5OLFNQM1GUabjHmKSApgVkJgYzFnDB8D85
41BgycFbFBlncL5W68Q8gdyQ6OZgYz3aoV76aHOK7qs8chknxbXSFh2uTs83Uby7
6Cgdp/YiwoR/bCsXTqo5Z+Sk+cXhl2iTHjNvHwwhOlqIITA7567VQf5+klIkXG0E
1uODB+ALjRzo7JoFOq3NqLt4KDBbmCLV2lJigdIdBVPmPjtZLXobKRUg99U5UD6P
SPBuUfb0WC5GofIoY8afoVhqM5P3biHSwKqULjmQE2GZ2y3NvWtQ816NGpiZfNld
k2lxZAuMri19XBKVyfGXYeF10xPSp8rGtqKTURhi0rsMLe5Qul+CuSXOmB6wtFKG
YRJkXE5If7JbJlgTriFTEs9YrSgTv8K8NANufZ5lDSAY4J11ROUBBomeduP9T/CV
Y1BxULSzakpx8XADAqdlGglQHkcb2maC19oBdjkotsKJAOCINj8Fp880Pl4Twx1o
Qq6dZsQTqgWNsCGkmWt+hxK69v/R/2bOfBkfHsU4KL7rJXio6PPN2UC6s+DyCWbp
`protect END_PROTECTED
