`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IRt6XJnkfGRdCWB9WjSDYiGd/sy/dWNNkqa2iYvYtbsgFrA/SJ/Zl2lgpjzWaFkp
aRvyADLEKleZs1jgwPyM+JzCZ4QT+OfDV22coHbG96An9I1jJOfoZLvatTCzSuQn
LwJRENUQp+KfKsE2RzLTQPKDkTZOijkcoq5iG/sH9Wg/O2D7mKhETpG33s9B/ZSz
lukYPhr8gt5veA7ZkncjuRumWTuSTBJmivUqCiHQJXtQsrtXLFhzDh7PJSpq+89s
qMVLzaM6uip50r9xg/buKvfjcwdLDPlHfNwiODlxostvORV9uKMKF3eMLyNL92xc
tCyZcdN+sx3Bbi94h1PWFw/e2vKrVgFBcwKW6t3zJjBf+W9i8fMsKMzJSoosTNc0
LCP3DY3IsOo3+Bj0Itzype1DWhUAIM+VxSB9WqiFJofqx2qWB1OrQ5lPYTYnYHaZ
UOg8pqfNLId+oR9an/wqIM8hHw9iGDFRrpBQqntx0Gtak69vHQYKRmM0DFAe444a
TNGZVmGEai7W57xm6Qr1aIC6amxCVoy/wwjJCKosAjEq2ySkVtwOtRBtAASJbBRG
0X6720/CB2AZWKWTMvPOINWa3mKDyFCCqtVvDOH0i/qHE5sfXNY4TckrCmxnF2p1
LyrJVad77IsiAr9DpR0/m6p5SpS7whZVd5au8Wt3dS4Lxhzsv/BF4cOaCVq4sr8g
5qMG6cVT33pNNaK0aBduWgYzIoKYHW8ID62HgJ+5UUMMT2Rdc3mBZuIGbrGKJ/M5
/WmsPU1uwqclYgTe/T+OSuGhvJsnL5KYSaZcCBmZOUS9VlwRZIA1VnoYiwyTE1VL
dnl6WX59UbyP45p3VrZu9tVx5bC6TAU7jXD9JJDKYILvBkGwFKTnTvytFi11jFyb
+dsXDf0N3uwYBtFafQIA0l2CX3GyqNG14ErGyGNgvFLaNFqOw1w6qp/PzYaV8PH2
xsyTxse6nfhV99jV9CtNduuyHIbuVWaY3B7/1+jFfR0c8QagiDcJeFF2Gb0EdqBu
dXAZciwMWsCEIveO41x3R7PT8GQ5cuGpE6VDVSmyzO3C+inlGqAWtw8GYbLIMfQe
BdjE3xscxYXEReT+FPAVr8XPvitAYC1z45NlxxyyHY/R02/zSiH8F5TrsZlWGgoT
pd9zOn3Az39e2TAW8MatqOGjm5xGeEJXGL60b2r/KLtyEjXTPS78WLjj8bMVgUHu
zYKcJZ85hW5zAayUirqrnzTTFq/Yu5+8i4zTV1jX9YhXhd71wQHnNCW3J03Dmdxm
tdK4XY3XtNjYbW5b9sYFzvGiwgfSHBlGBnQOqrtmlQzoPx39jueOn3mY3pboNMxZ
B1sUW3HpiLtN3zlpNOemg7zU2gC65909QG2NVBAgCXUxDTySBgM1MVgjvnYTGShw
n+7UbFk8Jnmf4wvrUFk6Ent6ujhOKLmeiUJTS59oLU1nJPpETexlCLyPkg+S4nIG
udULhe663rT5+9nKEXvbSqkv4wfg6oiXuqakPOyBsgcRWt817HakYwIYcwQE7G0V
avi1OmNI8deD7nAV+fM0zk1LjqrEn+YpawKdXGZi/yF7edVbAKEriQj2Lur9B+O3
bjCjVFEsysUfKYZKR0Cr9l//Nj/Hi2pdCcQ+Uv8KK1U0RqjK95MO5ko9ZausnRgz
3EcMs2F3bZOTHmd8WKFWmU2UteMe/vhs/NwLnVYtHmxSsNZLno2tt+pj+n2Fz3t7
NT/EKmmxlZBcaGCqCi9ZCQazwckj/aM2Jp/V7QhH/YiCMtg6J8XKSxMpDSokcptX
7hbQISB1bstMa5KMLgTlVMcJbb+jQvD3pNRBFbSDdT+ex/Uy3oJb/sF3XI5EKiP7
NMgknqhzkHnglEkQZ+aj8PKojgHI0Yofd1E3JMor1yNq/q0C6xm6NNCc9J9NDBWG
OIS6rwkSvWz5s0ZEfvkow208ytPqmv2mmDpCn1ugxqdJxOusV4Eu7Eb0Jm1E9Qab
v6qNwVlcU016WH56MQm+Y2QtmyGTWZD2NXcdwi+83lC+28uDvsZ8TzNamGVeHJYy
oTMgC9zrfowUoWWhBNkccD4OLrds5R98+RCJf1UuqzA4GEq66RWj8JU1oQ+KKYNR
7zo5W80BjT5ySGFTkF0SKQ53WmMtJaROZMdaP0+iGW+oH9UpbSP2T0pXXPhPPNDC
JWr1W46nlz4yLZHBySbNWsU/utgnZWdLD3MX16VYb1+FsNDOM7IbPGXevXp5PyGX
2ZsrqbKvTov4z2ssDywgNg/SLh/Og4wJMo0icHdqrJdsNpsRDjlZHWE4MnlAfNPE
s95Erb6Bx8ATBtRlqLzQjs+e7napmVkwFvSDf2GxOoBpqCjw2ZNWqLuKuenyKqcS
sPFEJcyhbzLUrb12fIhS4BtYgbf1Rj77Gx6m+Wo0LQcRwAlsilF/dVsJdg4ltPum
URzdGOclwtwlFY1asleYzYq2VdRegcq3D/7RZ+L76fqnOlrXxBngldpallZYpwdp
Fknnad3E5lpL8iBkna3Y9kHA6VBpuF5tjZgNVve11cgxZCu6TaerKP2E1NS5QEwL
I5sHGMMG7qWbQNu1xsy7rP6bKy9eHC/JK6XXm//suYAax4Lk45sMkyY+qBF4iZsB
AYZMpFrzMH3ZibHZlR2l+wfRNaToaWsJdOBNBLM4omr/YB1/vgl79dOZiE/vleH4
5i633dkiXMfacs+7FrlZUD6XJVh+mf5Ko4dXze9K2M9ryKiMIqlRBKj0v7BhMsJA
tgWO4DsyttbSYdZgTkYxMnz+FfGO+U+LpFU5gFDktCEczTgeNR9q/BZwo8lnGXLE
Dz0aiG0pyJGDaUDuRAk5nPQTAjjgmX0hjJ5eA4/nI7tRyVKyx1pAkxLr7zXu9pZk
WAs0sZ9mskjC88SeXAUI7L25yfYzJJm3YbjUc+6xK1M=
`protect END_PROTECTED
