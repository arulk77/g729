`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48KlNiEgX1AArSmK29IbzNPnKee50HBZS0EdleBitf7z
La1UzfP06cJJVI863oNhIIKGONeELYFh9IfE2UfFrkCNr8io4hZ5rQloEadaKR0T
LkuUKzQn27/vVvpNZJpFnweovqGdBAS0SwM/fwDJBrzuaNe9MO6pHySaQWby3nV+
mdSaLoTzH3vUebTiCjDBngXac0Rrec2KoUpEhxB9sKC00NstPjpheqnWnUGejAdX
o9seXEAMYiA5DYrZOyyGGLn0hMdqSWDNSU7AmXSx2mayoTHtnmdFJ/Vx8th2VrLw
UbMCJUHe3kfor7hRnCgqP/lhLPW43UYgnfk4GN+JiJLHPIYh8P4DWNgwaPMvSQmE
HHzz5IxIGucfWvNO6xlTdtpEwB4+Mk7wZXplBclkTlqTURdSbwuDP7rt/pTlSi4C
wsj7Rd0DT/ztUJzUzYDcYgrhr/PoFUp1T1WCBFQoYM+PkY6dR2Q6oigPrxq4R2cU
0u4Vkfdo6bw7oGJxAj4MQwsIcfDKC1QdsHywVI688pOrGGRegKRrknknTcpnBklh
pQw0t9d+gvZuKyiVWEo+WTMAHY/8NGSeAZzStgfyYZNBGkZcz/FsQgB6puBaNl0h
`protect END_PROTECTED
