`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
60QSG2IVIdr02Yqt7lup8pobgFO3CxvUu0xi873pDp9M3uQMip7UI9GGS70FZc3T
kivXMmXeIYtyeWUKyopSwv2f1RHEicQRa5OHf2QExCoPpZapxUcLHlpDFaeE+v+4
DBuxuQAko2j7o9lmcoNO48nrQCWiey3NnD3Isv+fpry/Gr0tjgfVanRq6VHiG/QI
`protect END_PROTECTED
