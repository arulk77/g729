`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4708nyzZDLZKEAPzEnxDwHLWygLBqB1dRfvAkieg+MrI
wpCyqNVJud4N4IKlk4Xkr/d84u9K0njIttZSesPOhKUvER4jhr1A4bzOw5W7Snjn
I61JJsXNKt89nyeAm1LE9p4/ePUd6fjYmFzOzTmppxuYCBsemYADMRHkQERsFIwT
Q/obN1+kp7z29DLBHPTxCC+bkaAA51tP+LqqAQZxWT4hVYYtj41+TbCRlV/UklQT
1shMwqtYuFBwVPg5nkuNwfx//QE2EWXwOGQGHr4va93CcOpA18FE/XpMaxHcc/FB
yetanqCfSDzwVkDMbca1wA==
`protect END_PROTECTED
