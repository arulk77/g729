`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8Sd45DC79UQUCuPT2TsEh5W3V5BPmEBBljFCPoFjVF8GQ
9Fcqlx+kG2J5okfACnBA1M0XgAwAUYmEbBgBUfxSGBs5BJahYWas9WglyRqCiDuJ
0vD7BSq4ykfv1p2jZ4gUu+e72GEVqvPwLkTEA1hz2E8BBwbNO5r8mHYH/q4pjfQP
`protect END_PROTECTED
