`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEyCZYKNDdVTDqeFStyvAL0DvFQ/SR0lagauXyyPxAaP
gifEUCcZkPDH2+uEdKjLSpeYKLfazuKWFccd3rR9UlV0jOcgegcyTT8CEwBE5NG6
CzsrverWqyNPNyPgwfYA6RQIsIvNstEQ6fLI5xPKFacyYWSwjZC1FDZI1cnm0gWv
ZUAVjvqBB8UH6m/0hnHvlw==
`protect END_PROTECTED
