`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP1jQp6qxReHx0ZwiCQgZTSJcjulfPtDq9aZk7o29cvl
PWhllMYcN94vXyd2cb8X2h10qtyaGhPgMRsjcY2MH62DmS9zmDc7BqVFsKSnBTQx
4mNoczNZ3oE2rOM+JA01k5CPT8GPa460g73BGWS7sDsLm4Mxiby9p6ti5a9VjwDZ
dye1kZS62l3xp2KQQqG1Kgjwu3CBZFQu1krhmiQ0Q2rcp2sQrOgzkQa/R3ColhO6
uZMGODzsLjJrEqJTI886wTMDp3L1ThrDLZqZKSnu1OlRa0C7bOGPriDRkgfN1cpm
NgQ9l4D84A46Xqmv1aW0x+G5cWwMVF0wUjr4EaGcqKqERnqsqcKUC6SwiqGbyJas
/mTXMZ13DJyr3RibEy8Fxty3UjCLC4H+Y9ttUvgs8hwe1JnEvYZqsg8W9UxIpjg2
qu7uiGTFw9hZYCnSYQ8tn96qbqs1FGdeEJPBiIUU/7uGDNO/TN/5JPHJcOPf6cXH
ZMcYmJkqU6sJ2g3A+9AAnScmmKmOhyEa2VDFi7XJAqqxI8DgrWCMP2UmT1T2qyTA
ojLpmJ1cHoyDgieiZNb2mL27tkzHkqSAPROlp/qGEnyCnhFgTLIPsJbMBTnkWUDs
5jL85Ps+Yx7p69TQACMsETdIitndq8zYIfiQq1yTlJNkmlNWjKYAbzvgrOPMvD6L
Bee9iatVIFcJOLcpZNGH32qWRsJ2rosdbJ2Rb2LGL3pUs8d7BGAo9o49QFyOjDjQ
N92ZeLLNlUIb+aYa8b1Nl2UDjHx24fe7rx9YgEtmXmfV7ThMfScqW0CQnzZ+s4TR
oHlEpPCPAsyzgh5YMga55pJz81M+FdJmIZcowQabUuk=
`protect END_PROTECTED
