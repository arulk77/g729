`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDASerf3uRhk74vegkWCblj8cSNXFQxU73EmC96aLjuggY
77yO1UYm3vKeQUGAZRXrfoqZXNojy4eeDpckCx/8cPQ4uKM3hVTpdi0EvDZduP3d
91P5l0x1SCrJSMF68Usj62MsCPKBmAoeNEptPCFDg4ZLbR2vyqFoK4ky0gRo/9Zw
8W1e5cPK64TUohOotBnft+XSoauu/T9QRraR5j/ymNuuJ8RD/wU7Zz4C6RpIBYIK
SV55/GLwyUdfJGaKJDpS7k6Eydwrc2g/ra3k5w7zGHX97jhvSAnc/JLcbJnuHNEd
hGWCRWFBMC+O7XR4XkW4u1lTWxOUarbDRdas1khrbTlIA5Z4oBrxYNyCatpV9VzV
h+QVHIzGO3iVlvk/qQ7srCBhRC44NcHRsfSSw+eV3j9E5UNsdzg524ZvV71S95VH
4iTWW8Ej68/bzZR6krZ4sqPSUGb1ZdhFwdTYJ/8CRUpxNMBXcrEx9W+nx05xtLCp
8FtHdtRVb9zmRxpgDknuIrgrq7xBEHGVh9cx8hBN+0OiDYfgJeeJj4dtCpqZMDpp
ZwDHP11fAhg7xN1Lb939GoSGsfh+609fYbrojtAl/DYTFl3TVJRtBSQ0kpSO6mWn
jt0JeOAJmyhJr6KgUgnz1292MKhZSkbCE6tFDF1CEOplQAEo55alY6t67zXL6Vr5
fBaLwBLCGAsLjW2S6Foos7axCh8U+pP1wCcypkRTVEQ=
`protect END_PROTECTED
