`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wKLQgSbEeHJE5rDnc0HgPvAuwFogeYmMS4dugLL5DEl
vO1ime6UcgNEc7uiizBgb6AxEx1wiUDKY34hQCHJEsfA6HtSG7hGx6XeYkMwsur2
QWLUl9y1KvOfrhktHQhjdiddkPNYcr0K2Fk6RJU73aykAoiXeI8kRcELZKuOKnql
+ZRVsV97Wrf2g/R2VkeDqBPM3Cjeta/GaiVxdOq+UB0ki5JCYhZ0BniCJFrluX7x
VTyHlZ7Mi2DhqE3CU6/smIwKflXPxxVLoHBgTkX67UZ4XTIxMooAFGmHatJs0sY2
05SEr07hw+nftTbzbnKgmA==
`protect END_PROTECTED
