`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QNw40IqJrFvY2E8HYWz+j0UNAeaQBSUMUMxd0u0rrVjXfkhrquHAiRj7h8Q3bAd+
rrbeCtY67+5zHubOtmgGZJCtvye/EAyTTDvXAaWm08H+hi2Oqp7zY6ZoPjOgPf28
KJ9Mg0RqKhDGqF39jLfeRweBkVuYzSawD6SAsfavbLvI0VvKd6az4qhZitliaNg9
+7TFXonWF5B0KSUlGcZY+KhriQLG5zhvHU2qf8dW99UdzP9uIYPnjTgq5GQb4tb3
NWK4ip7ivzoa2B1NxHq2cr4DPCxc1uMwcCpLR2AJQkpeBykWwVh4Vr3gN6gIHA/4
`protect END_PROTECTED
