`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDTrmiB7jcXIi/OIMJrE4228oIHUfEGG/3dzpJh7kGHp
AvFHSNM8i0ZDfTJqJc2LwdGGtQ7vNaoj3IJG8DBQZ3R9KcBURY9WOl+EtGFxPsWW
9Y2e0ifMzotopfMqcnzXALmLoTmQzRH7T6hibh1k6+wDwJGxdcOL6HBZVYPPnH0T
DwgLiHTEH0Pw0k1v5CXYbcvP7bbaUnbnDKgoStodgYyP5PeuMi3HG/c8/ZJA69Vq
sktocz8L44jwtwxH2SQUJI+34tMSDfKzjx+ZTKIClqLrIRl0elCzN8jz5ery3s5K
K+smgfOrOj3chybc1QYfjHIWkGwc9TstrcGy4S88Dr3DjlWY1QxPKsSdLlFXbpPb
WMwtxIlcb/Jlv0MVCaEzhBkR29y1DIzlHOAIuvc+5aigWCnHsDoqkpvNv9e9ejpG
0Jp6qFHBeDPB4/Rr7uirYkQDHGHgxaK0qpZEal5lKplZHUkyZhTdV8x2lKEKb279
6Ay6ZjWs/vPLEqoDX+bCvvKNW70qFvua6NBl8DrGs15F18dcMUPXxtgVLuFg3EHg
`protect END_PROTECTED
