`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C5gqlrphxMEJo4wDPeDUHYOcgW6WeqRADdT35CoNjRoY
++n8vaYLiz7keNoh5X/C0OFaQxgddcTPhnPjoJha7tG3LTmyipMLJ0AO0vqN4bAL
4E6LiKQrdhlOBrz7gji5/fpTwmtA1HUVg0yxhrD3VQyhVOSZn05xb96YrjU+1ft4
BPcx8cFVggHMr+kn+11RgDNkRbvNIWA1hjne9iHO6uGouYnUHk8HSqB3K31ME9nf
u1DNRAaIlBL5duUTS153uGlEND+rb/dLYmpVujg5eRQ0w1r75lECLW2CpzNppFn6
wm6RiNyjbhp0XAyinYW4RQMG7Rp7JJhEVqAQZuoc8bmRfO4robfWfoQq9mpq4m/X
agXK61/5WvyRo4Omu20kLSp6zx7xLV7AwxkUlvQnFCD5VuOhCSUzQgfqDYe9Z1nM
Rezgh+N12wNstGCdhtSC3IqGwVZ5Br95t+y609c8oqCuF+LdKIBTqgbkufa9Rtuy
KNAEXUjaa5gtMsYhkBO8+64QKZUhJxSqRlgsFn3fyh9EDUo5PIQ4XKHTxbQboAqV
GfIQNduRF6Ch0c8k+26iBd6IzTmjfRzqt73q4ZXBWysQNQUazU8nMEykVJ8nCDuQ
q3U+In+68rUa1b1mq+qIRhCNEEUSwNdbEsoJL5G7TYZ7FPYwVXU5Jq1BTIyB3nKZ
w2QlrbDfSfQjZ1fLvWxAVNcCeXNpZ4YQ0ZJKTQc0nG1oA2YUnSkQxwu91PerhNqK
emYrDhhn33jCMkv8erFwXp4nxaoT7Gc8KqClNM43T4cz01k/J6ymg9qDtRxs9Ds3
C7bLsbq9vIxHptVq63HWE2XX/QRvgztrV9QdKRu4NzT0uoA9UfCUR0Brzni3RgtX
jESL/rEcXQDtQVHmAgMYQeuEwxs17X+8+gXLwmoiK3ZCF6RrUS68LsHQa9w87lLy
1zbi3LtuXEnKOQBMUwHdBwS1RdF/vjZ7c9b9igHoPpIqPpXiR1d+pcDrWkH+M60P
IA0LDeDGG3wPVTREeCGfYif+Rx094/NR8WE6ur5ecs2vqsVS0+M5BnThpEXr9n02
l/PEKsoVhpoJMV0ybLtI5xThW6PakN8kQZWehs4EGyWsVSA4HL/E663q5gXxmr2l
DRzVtQpYxgmoDPfMxWTHlNPy57nCrzptULhkvj3HmgKKNGP6RQhlyS86/d34byCx
SLcyt9gl+BM2hSBMdUnQ9ISgowAkKwfdVSEpes7tXqyrXL5Axr3Ou2Fv3Xlb0g+n
K6xWpbAiiiMoCEfYhNk8+ztbhgBO40tt/U4C84LWCV9OGUU8438VeEILNxVcg83u
AB/+ww3GYnkvLm2QHCsw5/nRrs3HH2RGZylJ6BiG/aLYWprr5PExJID1/wNLnore
tpokt3VAhaYwRNM3XE8HqgQoRsxOfYoxKcW80EgStFR5sUmpsbGvebMj92LX6eLz
GXhhQvYMJRrbulNCA+DsbgaBO1EAsUPPl4O4eVczg8K31agdWkTCZqMB7yliiakI
UxpLRLbPb60z6dk93HOrfJ9GNK092O4CIFXbKpgY/jFwhrMWC6xQnPpI/xjjiiC8
MlsyIKyh21ayB2W0KC5NqNXGTyj0rra3N3t2SAKRJ+3Jpkn30X6zGsRpqfHhYBma
mvnHe8O/2TupLY4lYnM6Qw4C6In+/oVyC39jxdt40WoK/EFAoVjvTTxfKBMkkxMT
jVJoiMkqvXfBWtIYFeGjFpp47NsgV0hGR+1427wPSDPdDfCqgs5GM9yfwe4BObTQ
Mn1BEI7eNGkqX89Jn3aDgEKppm+cu8eycuZ6TyF/ijr8GoAz2Kc0co6EpT8urBpc
OeDeNAgDori5FB5DO/GNEjdKg68cDbzceC+wpUNfUJVACt1kkfIDRi6IT1kIS+bA
cshUmpTJSEF8/wz4uJsc+iDxFM4ipdCZWo+34caL5+apx/Plnw7ABqP9wZVlIAAD
HT85hGZxtWInfLMWOlH4EnNeo/UHk8ziwZJ/o+QToNGQ8g0ej1/C6CM7BCRRVOhY
WF0E5Tez6UJVniV2duIy0dgmBYtn28YhXdo6KpOocspnvVQ8F3iKkCLbr5jv/L7V
3YO355sy6jRlxSq9HDQHAG6WqPuEqQTBVfLylLC17XMCU25szXwut+HQD5kBOEqh
wsTS6LADNCBt+apJ3xFZ4wuegpEuemOmYl9Om0I5uppqIB9qQx81aoXVxX7D4FKq
IppZbsb6dK7/+do3MYk2K8XaCzGgXGxx4YRWmZBa+vBBgTkFxxRt+NRBuY07960A
FuXkbf1BaZ7DuOsX9qVY9EitSriJowJVH4xKTRe/zlnQ+XE5cRQNCDx5W7aLOWpq
RRazphsHg4BUKQmozC3Aa+w0x5f/ZZ8yT3l8V55QbTipUYsPvfafH1oS4NmhICCF
bxKupllOWKRYKOwys6aSomsOmtbuPwJeRCwz2qmbjyW/vvOyoQevtiZCu/gjBaR8
2gdb9l58q42z0fm5M84QlbxfvpdPKyHkW65r9k918hiufh70ywCDsaS4braHSm0v
cKInvDYGxheMbu1G5H75D8wqH4SE5+V0cnSVH47d8hnRS+sqydMDtTzmsn7nFuw1
s8AeQ85FazNUtX0twDyOPteMm7lo7ZAGiVuJD65HHEPwjzhDJrvgxiy5Qhdjj478
3mPkoMeSOZUrzUOEmj1cUHvRTI4h7kb2Iqmx2roa2O4+AnI/MUQ4FwZ3j2zflDBt
kWcSOTPSCc4CeDmsIHRHrE92SIoBpl6i4cWPWVrZCmfuc+4MJFskx20XFKOd9CCp
EbNwqGSLGA4Oihjtxmv1peWn3I+X6xhc/XekWW6hIBKXQxFUnL6p3z+eN1G/CH15
pTxpxFu+Vo4vWTF5JAmYqL5QPZqQk8J2R2FDTg3kEyHpUpZRgFJXJofqyvYVMn24
mkPqS+rIVT3ko3gVWOodJ+mXS4QFGdJagIYfUaK/Exu8gzcbGSgJbaCReaTrNcEn
A9q7kwoT4THW2aGtR1tfmh0ELc2B1LP+bSN9GkZ+dYgfLB10rq+Lmi2u/pHz4+YZ
MeapqV0NndxTf46RNQak/t/VVoP5GVaXUKz6GkJCt3PUM/BJKXdPpDQlhfsqy4yr
GfB5ZTuxX5j5gw6S7nmP6tpXJvdDtp6U8n0HO/YoRulF8/HpKEydhx/sgaxd2vkq
/70sV47VOwVSjZm1mnBQF+8JWrWYqmbNrHinjZsEVE0UXVdRvnjoJabK9TnXrYjT
TgCuT9APdQ/mDLcYS5gZdcCL/7/W6r0jbWifblmXK8B21lLYd/29MF6BbBxYs4L+
AOUKlJ7NKv3OPjaxlHzDl8K6gqaGDgAZ/HKa+/3/JLGT7rj7og+1IG5w4FVFS6sK
kkDzSq4gj3KzjP2cz314yT2zIyvecvqdWiswgMiCjn54xh16f5zhSW1QmGjmA2YD
bOT0S/dRw2xCw+S16R/akNvMqO60jev4yIkkSjwt3htKpK24mvBobtYE4BYDC95Q
/eckQhf7aJzMDJDOq7/9z0qtQBw6IUhyPNKA/m+Mu57Hia9HyDCznrKNTwN9PwtC
QNIk61f0rXJ4mItdeDmponoXrpeEcNGKBYB4WINfvQBicawASYUFgmESnQo+3szF
xD2hWubHz826Gzvwrx0LZrEdz/J0kr9LWSs9g0uwQ7rZvDCVh+kpS0f/3ZiNGa5P
XgFNMyUA8SzxqZpH4/GAYleYXjG9eLA0D4DcRG0vgzRABG13KzJwlBWsASoBJSsm
pda7tN1Z31rpR90rzMzmmKcrVyzKQ39QCjG8iuRVJGQ9PqK5yDf3dzUp0zgkUUun
2q5/sAJn6k4eDhoGVkHaa/VktTmxGPqHSpnwIhlO2zlXD4K0tEn8jzgUaTp00dEl
XiVS89NSi2IvPdYxv8W7akxvlIwZHsMnZzrMtcuKq0pqpLHk+ykyYs7to5C8DDMC
xm4gD8JmMGx1BHtC7kKJUMGsBjQCpYcPlBrNHtgVyXNp/RZanuaTK3TFyWrZAmgW
eYRRgr2+i2e6wWVYtjcvmxp8AdCKYZ55s0uhHqrQvI5roai8wd6KNFc5FyASWoVm
A8yW5rWVU5S32MZraI3myfwPSsDOtxM5ifu43zz/UY9TwvfCjY4Sk2vDgrymaz84
B8x+/I8wOJhWWwKDIb/bvsIy4S0NDVm5PZDCMcAdsF2PAlRje5TX3a+wielN8j9k
AWV5pXBZjgzDY2yF2oF3KFMc+0OuRewcsWIC6xdIBpcw5qQKY9KSe7B070ppWu8z
Dg+v50Cmnm6Y71olAkR8oM7ulRJbm3slCHu6aIn80Rjd3mynbpO6b4ILQ5JzJVxx
tbPVpQVUfpJxo2sZ+DMa2Kc5rOpHri4wzgNjgwsOdmsW7sBjwKp1BOB7Hz3svo2L
YGOvQbeT2VLi/x397dQnT+U/FCD1NuNrWBmxtmKOaCkQl8H/6YVglGAt6exwTd5v
KjoRF39cIFnzYIomXsrmkW21IbqLt6+3U33TRWgIqUIDnyacwGSQ/cwwZyCX29O8
cKKezopLl4HYM1KSSD7wMwa+QnBSn+WLmgjNcCDuFNcrIy9tY9RqcPrBYYz3NVwI
Y+ktQOv0Ahfm2M2mjPeoSlpHOjCzP8sM/qmwh1k7bTDoAALMeiH3f03Q4WcmmCHB
x4FYbf73JDXBranDYpbExadj6nmtYZOCpaUXryAR0WBNh2npbLaGrQk9TTmbpXTW
umAobxaI38oNN6teA512gEHn6Qf3cWbOLX+/uvZne7oyuosJcx5aYyz6WXXvJChG
lrkMcgg6yjs34kyE5jfqM/3B71X5HuPO0N2UlUtb9qHIfCd/05RClP5D7ln4I4ab
vvLXMglFtg48A06eq/DyrGf7fG9RWy4Yi4GpCXsKjofVpPTZssdDhCL20ye6zHop
/HypaKv8VJXWp4h6I0bAgRYGvrqWjtEoL7NRGvRDleQf0mKToilPxciQ+f4Zor89
Nqis9E5rR7zb+/tm268eBS0jWu7+skQaQkkvqIslzdxVBrJWdwDz/DXWGyXmTt6m
IliZzi/9CGjx2oR91spjD8lSzYZ+D0vQ2NRdCCKJmXGWC2lW4kfqK+LahruvSnbW
mQk6J7/aE2r28Jx9BEBKK40iLrUcmyJJftrziWS3ZNBO5+gvt0tO4e+H8e434wkz
SlICtmZFm4MrDk/tZM0SMyheTL6arYD3N1abm4Zp8MUvbtDW+5mbZiooU3plropB
MsNS7kgLNZnMBjHOBbY6Xd6ARASjMWF16hdFpRXEZS73WVkPSTclu29F5ayHpjvl
`protect END_PROTECTED
