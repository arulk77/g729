`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42KF+ss8Zs1rccp+enO3tv1Wr6xCAYJo+qcaHI405FRR
2S+787dlGKnU5bYiKN9mem0QdK7FhAzNV7qGHy2Xj7qlkvoPatKfCk2N0PVYiJVf
oNSdg5vMKxu6j1oeWDYBbb2U1y3yIUC2p4I6dhWqPx064sECIdkJRHQ7bAoH6iYv
q41/avMQR2zaHxUS8FhY5yOm1oPdkr29Yn2TC5dASnA=
`protect END_PROTECTED
