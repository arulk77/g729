`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMNB39inr38rHb/Kwh0c/BqOvBCdiuSPxG5+IznfsyOO
FXY7Cn+jrKl90OUdC5Z+EEyvmLImzU2k+kqh3Fqnfa8aBqClAeNLliIsh54i6fot
AYvjrQRrr0Ejcw6B16QV2eGKh+dfvY5HUFN4dchuXCzwe4yp7MKQXnrMyZSQgoC1
c50FhuxwZojCIiEBJZExLViTzA4jdRffJLcCZNh4qkq19VED9gEbiJNJKZcuZNxC
`protect END_PROTECTED
