`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMqq4+D9PQ/69P6uOZnQpp/2UuQhi3cDOI/AdCOR9Wl1
+HHMVhc+Aa0fas2pUxr6dOG37hObPeC6ugF9yPJkO9a+e7BfSjQiL+kFPdsB53el
8hCb/1h6E96DPVDBR0IvSI/cb06YFl4bNPF3mnTQMQGOF64jfE0vaJ+N3cCIaojH
kbEKUlGflsId+Y6kzpcI1zoZC0pehvfobmckKm7V5jyjhv8+ErPWDqW7RkU3sycl
hwI29WnW8snmArJWmawQjKP8/M/Rm+t6uPlmqXBJUFt6qKftxOnK2k8xxlEPYhDa
Q7GRjbzNEBSXFjBYZl533JQrA12fQ2vLlmf49vR9eueRQh3i/uQgtHqdrzvaueCC
ICuDFLCvNjM9nKR38EPi/eSdCySlFyc3DyYqi4p26v3NEeQ/grUnWCeMnekU17LU
UOcK7aRExHBxsu5DPOUxKXs9tzzGVxX6NPVOXSVMWCeBxQhHBFQIFvEKnilSjwA/
7lrpg2BzHfH0aqKTDSk+2rHQQObz8ls3vBy5rItDCemqY4/o0B/jjF+D/s3PM/pN
`protect END_PROTECTED
