`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveISarFlIGLZ5ecU+GuvMCwZaE3Z+125GKttQMGNswYo0
xFazc4CdD3OBqNdcVkesxrFXgiczqjFRqlt+SarfJVYkM4J+ZqrOPtQ0Rhp3yMDl
9eWmYExaK5b+r1EaEsuu0vU73u9YO35t+edTDB36IMHPJloilKm81jy/VfLO3b9k
/rVHGibn4nmdYaBx+jKCEiCVjK7ftt417ybNJ7xuozy9mUJTN+zxtX++Dlq1Pawy
QyxI9Lon2yqhNrl6xn0rU5P46qXS+Cn6cyQOheblWgFVLxH1qNWWdUDlvZLGWRoL
AHP3+d2nVuyCD0sUmXxwRqnDzi2TsAxjTzLiWMxPnFMU48+m26vRiujHETdyiVPT
fhY8+2+B2RuHQOimzH63/w==
`protect END_PROTECTED
