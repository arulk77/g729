`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLeZMrK7jmfJ74d3tI3PGj7FFlfXiYmZlmw5783BhJ6R
sZZbT3oJNOTJ7V9iVoLjpmlYOXCTNa11XUHjruDCYiyg0IQV7JR7AUbIr+faAAXn
5F9cR1jbSkekVctn7U0CC+BtNWVv42c3vsgcug5oQrJZqM8Ytvlht2UWkPs55zWb
aLp1/xTS689boAAbGP75IxIXuMzcbN2z0BfmpmXrCH/TvgbGFhLk/73+vlh+xKIE
kRcnWu9K9uWdNE1VJfOpukGwjMIVK3E8Eelgb9B+f7WdvmUoK3pxFAxdKx1lCX7H
awDtWIAcQcXmxJWBeC0FUaYk7KU1Wq8qNjdCOqbmMmRatd+PHQlHCfKIclteq5wO
DPKYN/TFRRMPGEcJpAyOOSMBAqvPGsaOlUcqoALFlI47/7bjkgxg5jbFrRSx68RZ
Bid0sONTxzbs32GOu9r8f5tDfEgdm9EPcnz8A3ZV/CRd3R05yqmxXIGiSdmeJQYM
73dH1ou13CugRSw8voCPcQ==
`protect END_PROTECTED
