`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/YbMo9iHDQoJtLLhjSQLE1Ik5FuYYKiOlmpQArV68cM
rsf5MuFkuG1xJ3zFwy4V27USCMGcpShfan39Lmbn3uOL0hQp/rUlhcMXgbdLmSo6
R+NNETv369FkOd1FLq2B4NZ1aMwtxlLgOJzM3t5u2OoAWGIANBNh53dUyNotZmoi
ZZycOVkXcqKqFF877Hm/qN6OyJEY44Y+pAufOnQEpL0oialBXAuQHNXLQrJbnvgh
q5JOJMy37nhfySIt2dPL/XnLUoepWgWKmvn+RkrA48Q=
`protect END_PROTECTED
