`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40+kGxzoK09ovoqIRRX0m1qoi3lPTep0dht0WvrZQicY
EKqU/XGsNaoF/YDDUNY418mYk5I9dM5qxpIf+Y/8rswkWBIKtgBZT5Pskrk0tPWA
1GcNQAa9wIpvq5KJI9Mczky97qrgEOCLQH5Nkkv9ki5u9GJ1MlROKpGkcHgqPaUQ
110gMMqx/1no4utiQQw+uccFXdatRb4UeGloWgT7wU3NTp10OMKWJgWZ2cb+y+iu
HqEZQsdU8vVhm+KHZOnPkALgWBA5OjIs+wVlpLiAjIKQKZ7vjHSCr9fW3dZHaQv3
uPOc8GbzLYbt0CzPxiAcczmMqQBzIUm6Rzib4dUZJXuJKIW2msvVJX+yRz/mk8hw
0UcaT3P5/bJedgifaA7/igun4KgqL3zh8knopQdwD66OO24VbXjWrq+OWxP8AJDS
W67P8oAhY7RHbr3l/s9kmQywTIfERch2mlDbYzEEKc92IwGTetuN23eruZJilpYP
v+1fOnXPi+VuGPvcOythSFUz4+hFpo9BUVMWmWFTxiRt/oyZora19vSC1yQ8iETi
DzQXTHFZ7fblol4yGJzwrI69nZsMrRVbJ+XTPJjM1aHIkB+rCfydceI/qi47MOpX
`protect END_PROTECTED
