`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
jQsbyFz12WjO3u76/T0s44dMHFOsfvUfQ9R309DFq2xsp7chqmoA24CpAOnjVKBK
DSPDitaL+N9sYbrCxQyea2vapgVZQpX6vXGitn2Kn40qmd8KyST5MvQXP1Q3Y2v8
i0Y06k53TLywdqfDPtbAVN2ezJF9HRssx8+uOT/PwPyFNUqLsbaXIY/tqTRK27d+
uXyaMtguXyFs2QMjU10uTDbdrkH90YoeaE5nElomUqGkH529vQY81pncKWHh/6dP
tIAds9f0vX1/Y9n5J3OMaWSImpaNYdhNBtoB3fNKary2BnXVEs2NLL2tbx1eamu8
x4UJdv0lLKgatB2egrDOePreX0S4uqQ+aQadtfINVUw=
`protect END_PROTECTED
