`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xy0droCyUQkWvqTfB6rJn/LWHBdySAXlw1sWi7g7ba5
B36AB9nOYj8ORs+ONjYTMYgtm62hXvfYdLYgAlBk7l/O9scysr4xTDybNoh3giem
m5vM5c+coxHDtSTN7e6U/3uP93DcZ0gKcSRy44hfsw9CbYzPJKG1AHNtNNHzx+WK
iKMJ1hobOWLitMqV62vq36Egk6hO7C+eCCkl2Tepg6kRs3cGQpvwA4vEbqZev+w+
fkwoBke6ZS+/QOHvXUhIWXDdWieAyDJugnHlToVEDJZdHyhvZH1QJPMUlnpgnx4w
CuvjjUPG6db0pW/ZKikH/PNZbT85BaDgKEm9F9VcLk3AA8+ge/LRCTsh3h8gLHHk
aXwrNMC+e6PY+dtiGNashmV9QSbcFPLRWMn4l/KF8rpAugd4Z/Ypt1I+YAFRKRGg
l1KcL96Ba+Cj5AOCcZFyZHKY25gGB0FdJrewLg7m9igE53FLHSoBvM+i1yS4/f7u
`protect END_PROTECTED
