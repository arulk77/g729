`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePjVz5egD26yyFSuooWOVJr5KtxgKkeHJznCA0DijTtR
uzHmJD70FBkj34i862rJJtTz1bZ9aW2RVnxd3tdiMGefzMA7bI8ZulTE2qRRMJ0l
cwzHlHHNH8pQPkTASoE/Kj9DDqUsdYn5A/j1qPghvVivWfqD7/FY1glF7Xwruxn4
KxDD00XUDka+YTy7g0A8HEwHf960CB9fHNdVhkmCFRT95DS+i8vGlYXhpKMKuKqq
`protect END_PROTECTED
