`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHLwGxsqnFG7+6JmoCgRrSCDdrAQnx/H13Jrr45JjX3l
v8DrXs7NCKGftT4FgeiKfprmj15uIP/OD/iSzpRVI+H7jwWDovgm8M5jIT3Acn/v
VmydLGlGqq5vNqwoelY4aWgKbxhH8uPzpZKcj37Mwq6yCXECJ2AAzTsgFa5rD3TW
J7rPgEum4LwkTQ3DVawSIshtbl2rk6jqTv3kSxj0NXrhRAA5f6UCJiRQyY9I2FUB
1q8F0WaDWXZGtD+3AK6qyYafP+aTjPAsx52IgSG7GyaCxep0LKghTFfPAhUDBh31
ftGM3tZMrkegtIqb9OXp7cOzr5x7QJ4GONmrWpn6gjY=
`protect END_PROTECTED
