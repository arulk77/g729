`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/w2dPh4HCJZzqQmE7A0GJTSMLawp/RxctC+7GEFmvLq
0/RRhLcVNgvb/Yu8uhSZf6JOuCVLl8zLkcKPnQVIduefYX2KFUyYHIILvcjflYGs
HSS4apnmZwPD31hCWzmJdADFahTZ8+2WIbYKwOTF2aftA5otKryTGDYtozDMOY3d
jcC8+Ch/l/yl3/DX2sGVc6A3CNszv4lNhAa05HauaRgrXEFGIdUQH8cw+rA+iIV5
ilfUtMxZfzyIovMS4lAUAjNBcoKgvGZJJphfiIuVSgm5jF55tIJJFdBUbSJTkkxO
B6JwZSUDVQ1E8ye2NaRMNlOjM+ofKPgbac77fxrk3f6mO3ufI5qdzuetp+G5ULA3
mE1SI1QPfRdGBNyN+o36mw==
`protect END_PROTECTED
