`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2nLc5REuo8sPXz1EHYd0mx6ag0AFk9wvtWlGOY3zs9KbNrz/aSA7W7azvvLMpBIu
0NgaaRbDQklbDd1mnY+t65VUTIdET/Qj3+/UKGT0Z2ZoYUm/XfFhy5lBVln1RROE
OB5s9ehWMjcUhxcOGIP+csJ0dm9luTQWt1+L2xXk2vCzs78wIuTkVhZxakba9KEu
oQ+4R0IKoDCQ3/imDdhIes+Xp4WUZwTz58YZDxfANnu0Iv1GpTLO3XdRgR2xkwRu
3GBWrNroiC21+Q4plwCJHimk7XcQLlxvSej3UIBR1l1EG8OQ5ZvCCCGyHQS46oE2
0Vuq1QE640yB7vEBCkKSfWdZvzvVonI7gH928LeXOvY=
`protect END_PROTECTED
