`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ14vD3aD258gmVQ8U30OrkniO6Ke3i8IsUS6PtihzTM
GVeSa5ephEFxVOr8zM6xl9RE/G6Q9KDIoi5vIuII/C+dU78SFfXaMewtpxUJDeT5
Mb0btYr0p53jdX9bgNbhqMfXGx/xsyKp+htxr/X0s04UdaVRqi/W2LWLR+mao04B
T31xYA5G5UdZ3KjFchGjyZlynEMUcZV1jDM/EqxO6WnfrMg6hs30/djoDgddSiHL
/yJW0X75fQDpwqs18nB8sjqdQnR4N8OIcT8WqCGx8mHCZbcoit+xoRR+JEiAItLK
qLSATngEA4vONtRE++7Hyw==
`protect END_PROTECTED
