`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Az3KDFWET6WM7BmeitXTSufqb0ssHjkHdTj2Dmgo9kUygLoHaNEoFDqkM47FlCKr
Gya+xrS/AdyG0zISQgz6EdfqxlSVE2tLNvQ7jRos0g1W5fs+fv6YWk/SABgPTeqH
Rx1EjFlOuifNQILCHrxRyEcpzBJcqNijqgmHNS59DOym/qZ3xnqMLWDie8B+6LH5
8YfKhqyLNV5uIgGaS4tR0LRqSWL+H42RPPosEys2IoGLmm5rkXgzYH+0HPme5BRu
OgbQ325gAuw2obVN1YmOASoOf7xmfSWFuRoHYTKs5x2oJ5bV5FceIChv/wB8p3La
POKhG2Bx7ERZmbhO39xSw5CSYQ/3DnHEdrRO/IhsMNT74fDlltHl/lN3jbPCbAeu
rG5Q010B1ncyhrjNlGF743P0ai+g9dndfOas0AN9H7byyF+zvJnU1iulqStzREFF
2mWKzI719Ccao06pRCMtlRAsSVg1j8GWZVJ2PvVFcwW41RVqeLrw+m5ErHIBz2+D
6xeRINWFvpq+oLN0CoyRUCYqOU+zZ6zRz/T1aqKcq35juCFnHTm+er03kC4xn2Vn
N0QwY5xS/fiEdODlJhN2dST765VbpR4eVrttaH39HAogtjmVkb55hO10ISx55ti7
YtF1VJ7cnOOviRrVLdbdwkCZwI0Qa0TEakNucZspgUKQrGdR92dcdCIACxYaPbzf
YfD1DN2aGL1PLi31Lu+qJjMxk1L4tlQdkyyjCXqUkSr66H3wzqfEyJv/vnzEYzGC
B83jzcaXY1WQJzhIujUWqBYmucswMnphH3NIPltgrDg7NAuMnnwK9k2YcuMvxJD0
2wjJnQs4TdTqU5JqvS3pTaGws8FPWq87qODXQQYNYIUM9ETtHokeL3QutfBesvEt
t60m0BkldpikiB8h+Z6aUUkyEu7Yn7zZAN6W/0BMBdMcXseK5AspCz77JhfE+sPT
exrf/6pvsZDv7UPNXE0Kbnhez0x2qpy5mwhD5LRfm6/m/iFzsqPZAr58CyfoL5aR
vri2A//gKctOdXhD3osO8jbV8Pjfoc7WqKAcsScYp+rD9Tud3KhoDWD2Nl2Hm4hO
pDR3b8VYyeUfOqj2rP9mcaChCwR6Is0zmwzpYmRS9JvoN2SLei7pu3npQfNCXy8t
vlpyTKKbZ9ll0Xd4CeZ3pM3jOOeS1DbTtoWvhPCw5zJcIxPkODz2Y2AYPq0pB8vC
JZI/hQwIGNgJlu8CsC8pXunNUmlXd9VcVdzfj3jgKQ9YhcZgnSq8052zDZmZj+DL
vckat7SFbaBRywTCk9kGQ1J1tQ7T44Q3e7tv1L109fM9eWSJ8D6jL7Ug5XuDxqAA
SaYn0CPIkOd6knNnYk4p/unmSFFnsI8d9LbSNJOwo46JUUBYQcq4p3mYRzp3w1L8
qecvNe3OopdKYqnVV4WQMi9iHHyciYGo/4lEXXTh0Su9/33ECoSfa/CleslcU+Qj
lLfC+5bUZxgXY8D9cJeatJCJWs9WgV9ye27Bj9IymuWOIvd4G7lguK0HQwDOzNrh
niHSRpcp4ZXgyBBkdGUsybEH5PktRm/TiotbBCEUfzy0ZJ/3clvnwt6XgmpBZrRk
`protect END_PROTECTED
