`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
VEnwEP6rhb1JENmvaM17URt0FgUP4AAelstPH0RzC/RxTmeN/TVOl5aCV0AM8aus
R86cnpmNUu4Vr4T8E/Tup5CEtIXdWupfcHK2dTHKAr5l489g6C7AjSZ0n+m6Ebzm
7GGKHvfxWXjL8fJgXrvmpCwEBeCXZdsd/FZjGhtGrwni284UrvtzlJvJPV180dSs
HUc1RRDjJmnbHZyqhsCieRTTAbjPaXwsdl/7iDsWhHiDeLyx2IzvwZGmPKIdqs9t
QCKEzRjioJ8k3rkIRqvDZ8GJZbjiU1VuGoDBY77txkPkM8yrkUFaLxx9SA6+A+d2
t57JHvXbFSfsHXZly65yqK2eDqOY+pR1kdSIjO9/9Og=
`protect END_PROTECTED
