`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDASAU2/E+S0+O7MJVVPzWjLbOUYPi3FPOSvtXwu6WCPMj
RJzLwW8/ozP0ht06YIVdHLiTurN3BCY+Irr9pYlcvVc2b91Y2jVCSu92BW/E1/iv
ItPOnD6KRbi9nstXZuTLnfsk5h2msRrMAyOXgwvpN2+kjp+S50qHo3TmMTH0nPFO
dCeK7TJ0sGxiKBrICgpFXKkuqEn3ysmpCRovTv6oVAutfU0Dsx3OIv/nsqcCkcOu
PmY4XJ/kKQNfaOAR7+YK+K5s3v8PATX4k10r0WfUG/1aapqJvc4829+zVV1eNfya
WoA27/7DDthHDYFhM8zqHcBs6aLW9YMqHX2G1M4MzDX3vuiYV/Of1jd4k9nbqsHg
QLh1gLaSZWpT8ynTu0fhWmAD1UqN/s5bsj73f49dI4RAIH81aRtvbZcB+ziH5qO7
JVUMTP2XPS4OP8Sz4M3L4HXGJUem9VDEdZO992VCWhoTjbk5PgKEioE6HamEt4FX
YUR/RZn+I4CWUtOmVrX4/HyM4aOlL+nwxLxkYuLu18qKcDGIkJaFznOZhfZPk88m
0rSY6esp/raU/ijYXwBX0/7q+bYA23LrkJDho04gCrbET264UsZO6o3jCjtoLf9p
T0a4y1bqKSF46KROoKpb2JnQX7EMAn3pUH8zGXEFg0IV3PNdR42Mg3KUllRYaY8p
S98i4YB1kVFN5hZrLz760CdgZEiOKMOlsrD36dkLHVvRR0QFHxTDk5s2vay0FXWG
7vDhkmzdnH0qtug8nvrzgLW2nhFzQDQBQjOIQj3b31XfeeEpaYOCjy6bCOsOGrMC
5Stsm9XVQDqC5IqPEgNwzqIjL5BabwBWO7Bln/EN8dxDm4dSccvuwM4ODB42V8A4
S4kzu00UpBVl/izza7lEeEgVsMvtPo7L1EsJ4KWSqb6x7C7gcgkjruKN1HGkoCu/
JiqFDzKeKVGG27XMXfnixS7LuH7Q4PurK16tLqfsffQQYo/dHwXOeEWgzFWhXIvQ
2Peaf4/phkTJTWT1amx8FNqS9iSXdRPK+5Sr163OGSkKMlu6lb5QlPvLYOdQWwRs
atESzXuFhXM3epr5bN38OgQ9feMoPiCM+gJOZ8yyPbbkr3wBuVIo9i3bhIMkxkix
NvO/jpYM2+yMGIq/RKl986Pjs3cmODFSg8L0p4iqQZD0tBeCHy39RwR7hcswoktT
hlUy376MWEU5wtZaHXFmnBVlgaEnCL2xZmca10XiqNMkhsI8X6WgOAO5HSubn+Gz
UV1bSMl0uqMeYUWKXMtGBnpeGoeftJHm1SNwtUxyn1EmhyzU1/+MFCSDh4gyx1OP
NPYpPM/WVYZou83TklVCK5E2uRUSKIWReg5+k08Pet4ozuMtbryzX428CaIqoeWN
QnJvt5BRrZuKTO+a4Wde1yaTkRybxbn6szC8fYpOaOiglUgO5LNbQWs6hkq0C2MO
USuoXit2M8/gJbbg4VXSC0FGkZaTOS8UrSF4nUHMegCM7G3Z83O3f60RjbrvKrXI
sVSiQgH1w0QMlb1h1aOTYmmWweYQGBNXEAZZLIptNTdMGTQL/l8DRpJQiU/UzYk6
oZS+0d6UatkGdYbxttleRFso+LkMQs2sEOVhHEkp1quMaa4GTem1EQ+y5JtmQHB8
rjTA+pwQ4nLmvF7H8bJyZOsXbFNx7w7uqPzALqX7amby4UztNpLMDefiGMWs1ppm
fSs1whnBNS4KjZBOVTDigJgUsPgFHUEVOxHTZ7gFIw/T3l+uz9vfCcX56uWJRGCS
4tvBZymdLxWvcK9cV8qDOnzG/GqRKBDsVdk8BeS+Z6lZAkgo2uQnOEUCqZeAEqGo
5JM6cIX/c0ejw1sZyF2CywTKu+9KZVH9AKGWX1djkOc81/8E6wU+E2lJLAx0oJ94
uIWyEslILh/8hc/FAUg5yZNDD1Ys/RjmSQuX3dZcIDOT6DgUGm9ehHrkXYECZqZO
2iPAb6ADMBhuBgdPX6CsmrQzI6O1QKvFqXykKtk61SjvC/JcXbNisRtQ0sGFHLZr
zUjsJhvXzPBtI70vxaNaNxtr2/1mxHwK0jJM8vex1iRvCKR/IQQmiwX0zqPlDE5V
Jn3IlmfkjWXHdqZXlHO0KOvz35/+p3qZTnabelqwuZN6KboKc48/HDA4Z5fudAZ6
r2sWiKi3byrf0q2KMzOmbXoAOXpsSB4AUbcLY+lFDY5me40xLrCJFUl6GA7DrZ/6
jf8oIoDCKUZUmL0hIvzXCaay154oE6t9e6CpUXsXFmfQ+VLrv4GNuzHaEGTYmrBx
di5+UfS460qvbbLxBhBiMXteZ1x57SApRCRMLvjrqoKGX8fnqOC6o8k5h2KzVy9K
mk9Rc4AzNI5eUr56ZLfRb4tss1POCYCLpa430ISpGZICY9aapRcDksrm8W3gfJxd
JroR0RHiVfb4L+RM2xhg0qDbk4gQc5j3G1gQYl/NIAu+Ci8n7vvPMjU0lJl4TNxO
Gp/uPyYuDA7/aYIUZJbq0XnQef2v40+uOV5Wgv6/vH/tcaxnJP1eUhRiAkXb6m1h
hVoX/a9OEwAVe0MxPgq2CzcAkc6tLMLIV5tYnqhk0ucx+t7Hpe/rkVeOxGivb0a5
aGS8EizhK1w0PtVroSUijlj6VNptqV4cDZKCgiHz7s194uTIhY5mtICzGHRo9ciy
sDdJTqCjcm21CtmGQw2Rnzia9e15K8ZFyX5Jjwgct0DUun+UeVI6fUOsSjKExTOd
jxGdvO/e1efBZlorO+uznq6SJCgElLBmiHb4ACWnN6cDhXlFhw2J32zHoTn5zRPh
MN0iRhqg2LZUDd7QzwV0iKmK4grvejXzoGcIRA0r5aHM+lgFgjq5NYtkqT8mlNt7
s2lKgxTr2XvRceL1wXcO6zgky80fvAsTjOMcEw5xl645HftQMB3nyRr3kmjjz0/F
6GpAZF9YcjyqdWOaj7/miP3Te9vFVcSuN/C889zgp2HSdVbc2sMWDi0eKPgK6BGZ
BssJnGcz5KP17JZsMyLMYGzVsSM1lzVV4iMlbiPWI4bc59ThNa0tJixBatUpKVQ7
SkgXA/MZohvkMqqt+T7o4d09jEfwgWgBft8hdT1rE7iZcsO+w5bFAaBkpLVWW3ax
YekQBW8Kol5w56FkBD8UG8kR/tqa3T86/crfLtuhKKS7ef5H933oLNQzkKpo1jZ9
CIAlSri7iDnXA0diTniB8eLXJgRZf4qt6ASzW7qlKNl09yDx54yeSmCqeQgpML4b
TLGUDB/CWplONf267Anbrq9Bjm9Abu+U/elUMmpdJBY37sUw50WMcXfpgAumemOI
IfZVqc7AC3wpBg79c2wchH084zI7E/n8zkqgsGfjF+MaeYmp3AOWXb561Lfte5nM
qf0ltk5ya3kzwhG/NORjdjrrAesPyaSI9Zk0XzkQFBV2ovVf72gAd2ihND46dPu5
ZGEM6S5XEnCNYqbAYx0lUf+RcX6l2sfSvuvmk3gkYHubDdJ8aXUnBvfJT2lDPPnS
cwZdNj+mIOIQ2nO198E7L+H3jl80Z+kygrJKSZ5kShJj81InGvVfzKbApzLdiCPj
LxNULO21bK5ayna+yKNEZraPRFz5Yvjyli4y8le/MJOMmRSuIeQc0am1IivqWdHR
NunhVzJcHXi1PfujPdKykkGP/mh9qzZOig4UP137PAJvPEUCkkQDarsqbBLL8c0N
OT5CxycCx1nK/7yGpzSUZuaYNVwOLd/4b2Xo/92sN7thse/xJ7/KVRpgcjmQyDx1
w4h5amEZBmz1oDW4135W1ZAJklPEKtDektwWiw5VIVKhDKjfCvAk2CinbJzMbAYa
rEWgIeuFbQjp7Rv2K+D/SPwhryT4OL/HhGfjWEFzr7UgXUCN8VYHoFKz8syCwroE
mSFBTy/B4fhRIHXHHPiRfWfqTTZKFh4hT0PyxSQ0dIOPWh8cWB1G56O10LS1TEL3
ElLBGfmCxhwHa5ebShmrabLTc103/4IUdhovQgDHS6cE8IxpAzCVkXdKe1Bwc3BT
sHW/xHmwQ0j9IQ/q0rGzD/MPqUKM+WBzNtXetRknA5c4YOcpdNMpRwqEsWy32Kfo
nOJIp+uL1awJ+g2rn5fEbcUuEccGvP+2rtJiw40DMyRl+gaqJAwIIjctMTXicmEa
wE29afayHILuvblIFQ+aI5Df8j34a8TWNeCRWbNDih0B37e9mglKUqIILWzsXZin
gdO5UMomk0usCB9EMWl8dLnSZ9h0NWhG+ekGVMa//W0IMLSxEkDVoXBkvDZaJhQr
IlisfwAgUkCVbAX1Tb96kX7iMAieMgiXe8jgDcM2I3LL6vm2Lnf4uOI+/QS0SPlL
n6c92UcI5s9IyH5Ir/5NH+zod+FnPZzqxvFGLAXmRzkG7+020CGjpKtEFOZwpcuv
RMLkkHxnm5+KCzV4GaK4ksViWaFGf5aYRWDSmXAivx83y6qG4K82U/Vg8GmM0onQ
2MhIhA7XGwssE/sfrdNW+BzWropv741SCSu0oi//78PrloBPHex52XnquCTJRjSV
HVCxRxoVU4WGQIb+eEVglwZubQzKRlulotN+BAmEq0yU4F7j10qnmWgMh4R9rfbh
oRirt3maEkbyU26TSlueoLuVxNCLpSIER2SVYh88hAvp4P+q9oJ8kfQCURNA5rm1
82+Aag0sdfMTGQb4srJq6wGLYey0YuKw0Pht9Y1FqY6R6AzKj4XL333uQJKB7iEj
VS0B3wmwQUGN0qKaAWP1ZD6vrJfR4zVxrvzH9xyrDDxJ8Em/qJ2tZaQpmP2FFGNl
8q3KlvqKgaG2ducgFXvO8+h+k8Tmw6bks8Bf9b4ZSBpZn87bHlVet5rIGVmRxGPk
ynFZVSx/uQzVZMMFVh78k4wTWUU7eE+4cxBSoeQr0PpwLG90tZyvHSsjwU9mYArw
WqljRA8W7tniXQ8Bwz0jrG8PgoBEFQevSkbs1COK4BAkViaHs8BBuMcIaLNo/man
xJtahv1txz+jMGK7Vd1PFkjPPu3PIMKr1bG69TnfRkaQkmzYnh9fiXiqHS8CBCGR
BsxKvMXYWk3ladV4MKH88Z2r9hc2Ro0liCtEb6eQGkREUtXDWV7GiAd4NgIwH6yJ
++IBxx3h+1PyZxnbiW3uzydYex0WwYBXYHM8AM3EcqoQtFzpylX0am5MxpazyW3A
VzBa9q9pjF8Kn2GdhuFzHHfA3jpjQdg3w1ONUNe5s/Nyrrx0Ff456ECAB/crsudh
HeIq1O5skUfAryLpvKt9mPesoTg8iBYLAL0MJh9Hto0Hjvey70iH/+UcjPrP7LLE
lsuxZd+FYHtsj9mCs9y1uBCG5J1mc8xGAaYSzYwAXGviwKBYweUKxyfpmgAT/bTq
a5rycRtihlSKSudga0dza2jVEjIyXbKS0tqPI4OvkIpw5T7ZMPYZSvODjnxAxBuV
oC1b5uHJ7NNMkk+6oyIDTrtBIQkwJ7JD+nNa1l+mmpv/OCW6WiBDnZUv8fzaAyAF
e3fPpO2duTPFExi4TDaek3VPigIOkJSLgDNkGMazSIwhWoUZuTnkBGzth73owBXz
t4VgVxYFJ+8MHOLcmvB0z3O0wjFfeIxZsJcbtZswRBsyufTegIGoK595DGLQRKW6
QBaUd6dwhXDITrjRFMaM9j4r7EEYoqnN0wiAqvkPhWgjsnsjfgqc0ohDZM2hBsgb
lFYS1xzWp3L5vllaASsYnQ/EzM//DjVJfkRuPoGXppVShLJ4nydFF0WIVnRfXJbK
e+0Zq1cWA0yOgtmZpfvKuFcW1/N4D50RyAD9fbJvzaP7rNTfJzBxJwnmBYt9httU
kWgIDpxzBzpUOVhda1RZ80jUIL5k0cBGFtVKFTSf8akPw8YrYskHwiycHdEWCi5G
5VTTq82Ko9PIk6NV6FDRAKLitWBcaw0pF2DPqt+CuNeB/Y4c/OsTNuO0XLFPy4rP
FjUc2IRa72q7oUGPIQy93W1SoEWlxWrfWMjyR0Tq8QYYNOk9/kvjMF1c7X9GY6JO
96dt/oSWgXVCn7XCvMkjD+oD7S7Ik3ykMX57YqLHniemVDCGrB7hOYUlidvCGJX+
9lvXWbUZmEoVgvL8Mkeblk6msE1rz1MczQZeX2gnDVtqdEIVaRisY9zx57ZrxtZI
MNhUveHPF4nHT5Ie5WImeZQtHNZzTCd79ibmfSR8bgjlM7ir0gXS1BhnR+RxFBu6
UJcHWN0sQRDTXBdVEB8YEQo/8PuXfqmjbt+BtQUCsk6aLgR71oiIrokJ8FghQFAb
pDm21tFNPF51m3aTh55ovkPhDtllhdfXfO1fsEwu+L1lUCuT/MsC642v9BSOSofn
n+6hVxTqHYpU6f/OXFLvGL8WEy2bEwhV2G24Lxz1/YU8S1xgpratZ6pcvgfYq3wq
qO89YrgmfIdiEY8muGUIuA==
`protect END_PROTECTED
