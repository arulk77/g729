`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLWufooga4ZsOwlZ47QoQCn3c18rqSs5XsmeEcqTZZOX
eu95zcsAIbYDwNMeea+HdsO2E00U7OZKD8Mia8Ww8R0ue5Rmn9kqdnhozlA10D38
sAzgJHk1LAHSbu+7eEkLWVGEe8HWcka+NkDb/1C4zXETckl/2+hTJDagkijYAlm2
plQuhM5Bl724fHOplE2IZWOdJHXeOfzNQrwQ+RDp6JH0UuoulsP0g4BclxuKpeFx
KLWoKw3EUlgzGtb198kTHkubVAc39GmGduc8gdO2Hpz3ADG/hhkulmrplk9hIw1x
NVPhBGSO9UnMajhSbD3TP8DEw+2aXC5Zg2DhoQN/WxDDIayMoFHysYz5g7axi5hE
mH/HekdhEVueF7eWLLRv8sHGx2lBqXdQxHUcTOKBAMuxjyYcSvzTd0cE++5+acZZ
0ayMQlD2uG73WJvcvBrdpj5J8lM3oQhIKUFTgXHBnckywQ9GeulCu+XqT4YebD4I
qQw2m82X6WTidB8SIoKLzB0I8TRxw3IuQ0CnxwdtpI5cEEQnY3y7bHZT0pzdZWOG
`protect END_PROTECTED
