`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCdRk0qxJ3dBpOK96jV8899uQozEs431EVusnYCQRQxe
MeQLJsNTeNCny2wkkepse6cMfg2P0vqDLwGzE+ApDXdsqxzHeoc2N3p5/vZNm2/y
BRoLvB5Qv6HEs06KauadgUrFyz496xYg+QM7SMe1aPpnxfD7Eem0RMCrbCFdcV4C
0hmoy/kbIf4/SbVgD1qKtSF3Xv3k+9Lhezkdn5USQl2uhoi3uaEiDGpY84gc4blb
e96nKWYDWu1KnSENUcfygRRNGdkPMK2nQalv6ZOU+dWboJgQGXbQOmPbnTCjmQBu
GAy3rjqbJqvp+cuTfc1AiNGxhXI4c/Gkzn4sfhcgfnrIrOiTIdTHvq1xPkzH4Akm
mlywDBCL2DNwnOnq+hPuFcvCeyGB7aU1cUGXCdurrRTnQrdHjfk4XVWRX6z5kZCE
cTdJ/KFS97tg6ZPwf6/AR3V1mAs//Ak7Gyqq+rwWqnXhPfHaB/cYkV8Ma53TA+gO
WcTMVvUB05mBZOT6C+Bb8AaVdfkzYnV2/raPOs4l37dVDB5aBmqz88k2XHsyaKo+
V1BV8y7HBaCQHAirPk+QATyMPLylV3ZHbAURVX2Ae+RRsRUxXkMMnecT7yClEdde
cPqKJDCC4lNiw2dP+jd0PRGXCizTKrNg5mkBs8BywJPO6iAIXSAG+5VOjk8dXfGN
vF3vmdRcpTu3KtFQN+4lIe4toTAkoMY5CCJAt4Di+ftJHeA7PG2+pNzbVSbUbYEY
0Wjxl8HBFz89J97djM8Ketl/zzISbUa+LRZLHSfcxBapEfDYrdWXJpcnXsP2n00k
gIZI/q+9u09OOOQ+g2qPtk6nTJLLdCt6DuSwEmRQj+l0mKSF/co2/Gb4OI30rIuW
RzVHraVrgkfdjHPMEMW6KPCXrZBjyFLQ/SS6C7Hz+C9+epsr2sANRNY3kmAfXFFu
CNqfpmBtlTxdViHN8YuJhuD1AOSWHbxD+MSDf0Ptjcta0cbTONXn6kgTRWI/dxex
Y8Tx7qOX2XAVEU6pYGElsKaAwpxYTChKn4R5DaH50VH+k6zySWwr5d2QECFuaUBO
p+BDZFATFsOAXTj7bP9Kl3U4Da8JZw7qsDAfkhZ3UpXzuD2d2QAkwyWgPB1fDcHM
vg+Dw1ao6pjhsexwRCUMF5PuSYm4JGk+om1HJ6aQiNDbO7TiMYogJ/Q2EnK4xpds
bxmC/2ysQuD0zYm/yxq0uGz5MaUeqo0btcNujRTLZfFSzbUC9KbQF2a86paUSowF
DhGGMih6Snfu39E34yexTIKgRi26cTiVXZOfKaqubQUs2mTY9NLR3tcffCnWKScg
0taA/L8vyD6FGxz0oY9tJYdxPPO+C/XSKylHD17pklcQqVt/ZUH0QxzRXGXx2s8C
b4ChzGTPEyq40rDvgwreT+zDIofo8OU00OJSDbPydmYg5QOYhWNeqcrHH5sRz7Xi
YCYIQzefG2BLE15prqoewMfEv7cL30RkdCLK9Ft7iWhRR68mnaUHGZPFXU4e1SY0
ar2tDkLuEvbXrRZlL2uMF46c1d+9HokbU51GD6naT9AY2mg71R4N2GAkk7s+7u8O
GZnNPY3S6sU6rnXNiWtq4+rQ3Zy6gI8omYSyd2L/HdyuAgE9kWSm7lSuVOUpLV+H
0g+JildOGeldYalJb32RS9t7rDVqbuLO7HsKSCAD+hKh8l1Z29CaT3KJGSJIiJ9X
yz8+bLNbNNJ1/ZR5UnPem5sOIxa560nmN8kyryKDfVOWQI7dIo9sKA/27bBx+cho
Nq9rKWUw60FR+xPuevD1oiSSf/E6frtMc5snUQAbWBDMb/Ra4F58LcfC/ZUiHJ0G
LdhfWbOIBjpwHfZZtjfvD63XFeewJt56bkZMfOu5TzpQCZbICYw0N61c5+Jqs9A7
XWlStMVr8cV2ApTyzwsLEeeq89jJXlAjDOBptzybAqQhzKcb53If13QXXkfAQNuK
qc2sZ25V4rlwTjcZFB58xCMjCeb/QdDhgwqWYPNtOWMbT6w6xkmPDZosWFJUaBJW
UWqxtT1TIzsgjmaBM2e02s1xcZgUNz6NfU8fACcL75sjuymF+YsinwPsAJtdv6Et
B7xVNGGxB4n5RgX0RD5Ba8+Z9v5rZskZbIwsqtdHgX1trzXW6wvRtI2BMFckhvqt
OA8j/3VlqAhrIHJgz4zKHAwaHB4iAZR2L3GLkoJq192xzUEr/jKdasB601RQ/h8b
UumPb988kDUBRLDzmFpAhYhdtLg4RyCydSaKRUL9GqwgWoQtziQmP6XBogSfjCor
EcmmnboXwfJl/4H3z9XXluvMLKYR2nu/tiOH83a7Dxsobbr50AeH6JaoEvvQHmrN
L2DER1P/aYBOV+KIMW1P4OHS2w1tANC+GVQZ4vO/yxQNmuAUMKDSEBjz495hKhia
orcQB0E73cza4LoJArFvPsH/CsjmXw0Wtwm6uxYu0N2OLec3U/Ye02Z9e1dDOkr3
9k+KRLb5d5R2lJWRvI8tfUDMHXu8SOUH2/NJn3lhgzYuoa0wvo5K3TYn5h9zdhhp
bYYMI8yqVAjqLKhyEHdH3VnnwsX9bYlvfKDG47yeOGSdMQTIgNg7wLzO4fk31ZVw
xh/0rPXe0mU8lMa8ZE72kdQJKeowdcVYhYDtXpKz1116sCYcS2l44MJXU5OVtZbx
0FuIJxDcUOH6D+4z1ZPJ3AgpM/6F3+Uvl6CwsY3VCQG2rWs2lQ20FsYluWh6cbyn
7KVy5S0k+YBY0jgaJi/5LLGx6wgP9EpfU/tbe2f61OE6TcsJVV8yYFbekzmbuTZS
vFC/4eVM0VqMPq/upAxYoh+005xzGaYg8+9PdxpeN+pl8LNIz8VGavXddcw3iY5I
R+kjJOPllUv2uV/Jk2MLMZOycVAxK9ZsgExgvGMhfbyKtpz+zFEfEYh33ZHP/Q77
VDmYlTHTsMhWfZzwDZsABaIL/ygj9HDDyJoknk2uLH+iFYr6T/SWxWvu/FuUEMAp
XpcYsqS9VpuTYPePxxGTdFO9c3Fiq0Aa5+YuPJz/5NgBb0uYnRA63TGMg8ZdoGmX
JDCsWeZsIBeKJiX3NUe+nVQ+1MiykDrY3REkOu4mNInBw54ffmwNdbuNJYxkb3Oa
KHaGsGcOPzHWNhSdzn6JujUrHuaTGduCwTrAwYhngnCCddIhXcr69IHDPbCSxyZj
ZjK7eTARLErZKYR5Dx0bol+KPDtTxgZzlx08KerUczYqcjSVDXqhZbiSbrFiKhJI
Kd0SYb7Nk9zDyV/VRP5RxIjW7E8+Z6gO4xNivfR3T5QuL6vIXXOT/PGXoQD9sTNc
uJqNKBxRdyxwq0+VhXbXQTq3UMJwpW7sBDmygCspS5AdgrooqPUeFHVu5PxdMIEP
vAetZxyxAHMqsRoYLpt989UnH5SgS5cnWiU8Ppaf4RUckd91/2H/W3U2EYfMlqtl
0AK/v6Y5PO76aT/mrl1zFrOd6JXb7zD7yrWkNsQbVREjf8xIkzOozVwIHR7dj0Ts
Q9T6C/nFwoWOcgOFRU9iTsgHHDbveNNNs3JIsM51N5uaCu301XE7fSMRUyuq+2jU
8nbocOi3t6cJHy87YDziaQFXADnjksA4jXWNVGgtlSbRFAslKrBRhNTTnh12Q8yf
8o3+kB3ljHVa8rvyvQ3jS1V0myaZZgj7KIMKJltoDMXOIWgJ/jroIPydDKNOrzMZ
bN7xr9Anf+hD//qo3Fx4IvrBkPYJXav1QBk7xzQre8kQnyscaGqoYKvqvIIFcUBF
J6zC2Kx+S/mESth4wuzGLBeW3QqtvNNeWmJC4CdUamUigbZGBjpbmyn5ipAQ/YVS
4kIavlI5jDkXhL0XkJ+iUdryxP1CsOCkiBGsEU70+XDEZs3cUNvEZTopcXOpYgjx
nkGHmuBhUHxFyJUu/ZojycuVQyhcIQY1yCo6ipiJZLayInH5lbJ9a5cpAnv1pLyv
4c6Uu/qB+OeZkLLhmELgv4qVFoKGPHdz2HT2sF0HKTufqsFbdc6iN68d8yX7UbKX
4XoAfPmA/VpgeABic2TC+9w3W+RZPYhrH2ZcIuDjB6BG1HYto0ZvUaoZJ56cgWSe
v7lXuzive3xvKYhw4PvkGf1/x200NrBq/ptuM3DFReHaV/9XmTjYjYruLfcLvys+
qprGrl9xATNL9BeoObJo+za5LOAdgGl664PaxGNqZaOhBnBiL6ft9w3Z17RzDrHu
443qSN0pp56eElVCa6Q3EfH1ztSz9FYifYDWRu738z5lCMLaa213JKdjpJaPonEG
BVYGUEUmZJq6xQI5MairmL9MOO0FqOE1KRtLPxQuvHNyyyuipcRQGVT30R3FTGin
dAJZRpDOhr1Gnxf2SVutxmawg0wstQidcrau6lOnDTr1h+yZCIBkQ9HFUui+pChO
ixEo2WaloNiqAx0bwhEbmWNXu25Jh/WiK9L/Z6v4Y/yvupJqGpOs9kMOWLFvXD9a
3/ETfMdaRvUKvYhlA3tXz6FmUhkPNKJJZc15BBh+V3qFJQfwjZW7/v9VxZMd92jc
M33lK6pe48HsDHUanwCIdKT9xyv00K5ygZgUDfpB4HqojrlPqyj+6UDAmU9PkjdI
RY32xL5+BR1rDIpAj4CGIU7QRIU98VX43NpxsNRB+YToAZk4PhaLITKUoytV/hUl
ZBIH/50Ppk+lQ5dyVXeRXJKr0uQepHtR1kydV6sTLywFNz2G3KHV4+y91GNMlYt+
5KDETW5YEl4yf4VR0TvMAnwpcchLgyqE7jY9J8upnDRFm2bsFwapxHD058YaOoKj
vF51SVA1ziCNtHmb9TImBAVcO/yW12HkmdIrtx8roDPPo9zXT/naBx5R2Dqb8cqG
KH7a0fH31PpJ1OuYOQS0Hs0pSIdUmTtqnZASOiY5DwlQAwoWlYs9i9Bul3qhiDeq
P3v759sLzejccRV3wu8MNhisYsz6kki8h7vI2sM5jTYP8nuEHrw7nQwWui7rvDIi
qUSCTNw9ONtvjXzjmag7UMSMW+NMrLY5F0lfIQBl02V6TXhBKVE8bhkyuq8/Fmnt
tZK05gtJ3NLYSSarRIGOssAPM/To1sVB8w/6RH6OT0CiKEVd/HzSVWSV+jtjvCfr
PDW2disvrsjHnCcdn6ik3HnzxznB8wGkPF4AfzxckMPXkjyD3fHKpPrVCQl0aYUF
qCgraf9KuM0tux7pDMihSNjUqYEtZqqQBJvtC8vuoQO4A8qU006QxEumL3MN08aX
qYzC17WLC0X39RNDk2E1CQJreozLLoNNgx6TgVvHKmBFJ9Gs6AWWtFkmsfsVjadX
bEwEL6MNEX9ood20i2VgRKi8mipJZ/uABK9OrtePZ+FnI9TimasfegdCgZVolSva
qftL4E6Uy4AZPb+DPPbvpTLQf2o0iMAbxf6l9NTgfBhGUFk6BLtkBFT3NNYbg7x5
ZCbHsjkxPjL0/RUdNZOrOEFdS+FxxDvr2y4a93T8KvqmzJdY5zY9p5tZ8tOgQBmW
Dew+9oeNH6Zkr7edJlRMRMbfyeXe2gq29oE5fwDA5Wm53thCh9Lsn1qesR9C/oL1
uFmfv1jz+RCx+Y8PMF1mAwYcrsZ030Tt9UmyBnEG6J9B71e0D8YrfHxXOJHIGPyO
vAisyfnALsLKuhCIxzsktj+vPj0KE4k2o78RNjVWWm0mjIoR6Kvpu2K4xrybdIki
Fl0H94PgF323xj8MDbAeYrY5veqQpNorAU25Ph2JxSD+LivLXL0TDNVLFbijDgXz
XbtdzA2YndpyyaNwVOZt5r5R23uHEVC7A0mIhEXUdyv5TY9uNYcQuiC172hOW/Fv
KDCC1cfvF7Qey/vPk1HyEqHg56N1zmQM62c+NkZ1vnSJVYilaQSC0OO6dVzjXcAJ
b8wa+vwWi99fyGLYEmrP1MWSsXYAsBhrjUn74tBOiv8+g2TzeFfyjV+9+hWzbO7N
chpnGsYoh+FZ2ZMJTqfRYuem5mifikwUdzhmr9vEbIHQE0SVi36Ud8OO0wpj/fWZ
FnMbbcAAF0Bag7ewNu5yJcu/6mTVyh+wBiMfuMqP8oC0ZwHTUf8AIOmsHd+Wrr0K
ftj3GB+ML2DBoBGb953Z993KLrcmSSWo6//KPCjWxX2FE0rDEpSCCTLohvglnlJk
ZcnlRhOI+Jm1TfLHONR9il9XKHjyXXwn3ktfSiRYcqpf0EP2akxF2JuIz6f3Ux2/
ND9DoUDDrkokV/bXWNoLkbEJ7bBln8DPw5RPUdVFKw4Iv2lInTUeRel0EVYyZ8SU
X011dklN1lpMCrdXEuEC2t0m9ofu1ShbqBqEaYXnnRrdvGeMv80yAarRzFjQXHb1
B+5WI2ty2GMROVLrkSerL21hRFnJ1ifW3cDVMf8bFm4Jx8h1JsfjJLCm1wBZr0wX
bdpTVY8DPAFEa2vFAidIjPrZ6iynQDZi3KnhrMyCVc9ne9cnX1J5Mq9FMQK/sxUG
WXOBLiV17qVQHxrdhc15R6URh89/bMPi+KRz6pey5q62H9Fa2VkoJ3M7XMk6Npbv
TpBlKIPluGINZ/sEzNZktrp8z/vVchBZVQ/+k6H4z68ojDNU03wKxIxvwzVf9tpD
T58bOocw/zifhab5eo1HJnjSfnZbyx6YSjkUFizHitKG4nnuMOPa4hFl0vgK+6j6
oZTuORRSA6df8rozCET0fburXQRw9G0d1YStm/LBlI+kjbMH8/VqlbvjV32kW4pB
bMpX17Iz+ANRN7V2Ll0hGXLYUH2YhTr5L9Wfv8m2y/F8HzmZFBVTQFGHWE+9RElu
t84B7TX/3x9ETPYTzquBRNgyBniOzTKU8KkfENATgvWLBloGEb5oPVOxEtKwnglP
rkJKgF9crKqQb4RJO55aRioj0ZNerSn5czD7M9DZwkewVgVAGRv+WBI0APVjIiGe
4wmK5o8ml8ctFeuHu85pTSUpeAZjEG/nI0b9U9zviXvWR9TDsA7/BrowLmgGPq42
AFjSD7ydceThn72k8kIMor4bnjxfnrHo/aYNKPkti5NKS6DzsiUrgJ6x1H2ojOVI
ij9LQ9t4pgkCw7mhYvGAFyyxJ29qDUsveid/4eq7JaFji0MG6udg38dkvhgkCrcm
l2xrMjz37NJivthIGQwiRd6/xUOhENZpiGF5L7/CbUOJiu/msxmEY6cVaTDFVnmI
W+ih0fG0ohJOhtvSw9gNhr2Z1V1tPPSrvdD87UWttjO0aReI+V2GZ2woYNnUAr/C
wPpflexPw62Yra6AOfDHGhkMU+OiIfc+7ys0a+CjkQ/O9FjWOTNrFhd1vttKH8+u
BhVDCZGVxkwUXTof84q2xaL7TP+Ynr25QbA2BdgiwZIr51aHL8Zrnc5CzJSCZliA
T1LKA7MODLyLGQ27Za1VrhmMRIrPzoU67lkWAGuz2snYZvjvSB2kb9z+AFBRLYwY
bctckl644pUI03rnC0PYZhCERMcHqOfx+kyjHmAXewMcx1Su/h8CXFVZaXC3VxRd
3mDuSG/KjmO9vtFmYFjxlk14IXKtJFpi31AlTKdhEp5WRI/FHI4gx6+Z5WzsNS64
nsOidfdW8cS2WdGYfefBYf+OzOckxYElmGgGaUDqSS77VpbthwZwuGI6u9Pk4oYQ
jCuCXuiyuk/cjF7tZJWMZhoRW3o1ksFQKfcPx3Sr+nliuJmSvSl6FVgf4773+n2V
K4vM6YhXCzTuzEEcPMyxVIfWpZuv7i6DO5osWtveDTu2OpJXi/hrCGCQRaslgSfO
/ZI8jWFbRlvEeX7Bhhb0hJkrWTLDLeXe9kIF/HuzrDigoqJzrVFqOvWUT6oRQ/GU
rRTYPwxgZwJxwNeVMELYpdyXqzDhC2WrSIJedJCkTeQcvxVel/+0+dz69L9IhlcT
wYS/HJ2hh+XL0MMbXk7hBNb6BhBrdXP8b88rcSlgTClaQjxvOA12gc/8tleXFynv
BDRQuUD4grhoSPtkHvdevS4ROWgok5Ja6TZN1n2YJrQLj9z4D35/2Qsts9z4cGs+
lD1tehIQVXfBPXYb/vDYaI7kal38vSRHABv/BV1NGkzZxAWLR4KRemkun2Drq3w5
1MZmxLr7iAW2YrKt1xYWVqCQXrfqoqPlgNhRz5pMnBpRasQsGD3Vnq2LCBFAhMoT
GBCPLY8YJ/Jx5lOCpkrh2gJ7PQ2OO8IouFPMz2jUETuSGsXXA4CkkekSVULXERnZ
xpT4+FGug0/1IRrW4MaElA2UfnvflR8aevGCPhwRu/eyZIKIloHd45GvunC172rU
iNx1o917uVWlK6viLmuoOj8eCm2GULGpp68kfwNB/Lm2G4R7OBvtN2SuWIfSoiIi
BWFC19CpmJ8tPSEM1Dlv6cI4/MP7BIR+iliJj3BwBRUxwL1ZFYx4LIHBwxjWHMUW
PjiI4/0siocwHpR0m6tftUIRYz+H0Xm8bxwUIgGDt5bKDcFOEAjDjsX8ESKDtSBp
Bn67OJKgjv3SKkZkPAdkvcJzw4JZsoV0Lj2qDKaY2aumTy8v1GWeqs0VQ0omkM5b
wDHPciwncHW9gYTdk45Tb1F+WPxz0PYcnaWkSQcqZnRh/siPkOc78xFfXRWD19mH
bBEaPRN5p+D5av7fmuOISWlOLtz1lzuegwU021PAN9B9WUAPFrvSIPQW9EBjyyNS
i2Zb5Z1qTuM7TSUIhjvKnyrIXgCkAUAwE9UOCinPwLBc+/Gshou3szC1vPQgFmHb
QtWy0EB0SRYSBXVT+irwpPvCFJJs4nF8Si6ioQFGHEFS27vTgyLSSW2Nb1OZCaCp
qlRqJ+PvjhnxogeLttBjNx7HL+bnh30eBXMOoFuLZvEOj1C97eaG5GESyc7DtjHR
YbrUCs1Z5MnGOzOe6jn8U5qo0NpVpkqBG4TjhBYq8B5bnyDWFuuVfFGvRJxLC0sf
CpTR8Bh1XE4HpTpWEkcoP2cQw5Ozwt69lN1NbRU8moH250bxCyANwqhiYQGlfkzf
d1cCuAzJXOu7Y/bLIHN8eGrHT/QoRfWLnvf+Omnbi3Hqp788VCps7wGE1aKKgkon
S9LnBmhiB1nxhifip7M5PnOi7i2+Tu3eZz+PdwFThBHW6enXa0DcnWNDwhjEUU5k
GJTMzTKDtPndoFSeGrDB73M4PpYvpRu6eHHBwQ9DdD6j55iCFrXOu/qWCEM0l+0M
UWOov7B3cOYFXstKu/HFt9SeXehwaUHVGGb82C57rjs0lqJWBOcooWQtmPJQ5AOv
MMfS8y9vAypMWboy6WXjfvjientfVvdObXMXA50G7khvfdi7hYmAQlBg4Vl/2t8z
a7W9253WFOedHlook6iYjg7vfgh2f5M0fZIJ4S3CC2ihCEYOOFWXqYkryXpkrFFV
ScQR8Xl/iouRSlBH4IcUpTIGDIlR9tIzBpIKRlDEbtCi/R7uTJASU9pD9YiP0qqz
wyeXcw1CaHaTOqwgLEhCV7ZwqFyZnzd3fG3HqfnucM7t327lDF4x4Hwy3BlebLD1
zi/P2RVNVkgNfcaKpidnHGPVmm5OCwKrNtX+ACHwBKfWJj78bWwhtpxQt37s0Vsf
xAkN0mPPpuDSvUE/fxu5nzKS3gSjnFZ6AIhiy6eXtucXZr5XlUmLDf49C8vqKWWi
V9ioTfxAsytE1KVUTiSQb0GHRQ7/wsr8Ek33gbnHju7K1SG7Uks06lcelnFfISrr
zNhub1u9EvyIYQz5jdX0qT+9eOUPrv5VY6gPRVFQmlSzv5xYtKNFDIGPyTcUF3PE
Om5TbpTv30uXZY5p9ut9Xx9BtBF7ltFiu2tnAWL+tigS26n26OEeXy+fIgOqM+F9
PR99sgABSlTO264yqRKiXqby9368oMBskKY1pAoyvzBTUyItzkPN/0u1O7ntqvot
ubAnaN26xGA990BOry0hffHxgK7ll4sBBcG5ZzFBEx+ImZtGysRJeZf1fnhgi+Qv
dKRWy7DeNrzlRdO+RbLwjkQU2iOps/ibW/16QGG4zYuM5oO+PXh2Nf4ZlTJDKRzn
327QAue8xuEK7+dOllKPXvVT8PX4ftqIKUQlOOdqDAGZENojF2DsScsCVQzmL1HX
oCnzF05T1iucehvpzvKguTUgebGdXdmLsL+3O8RdVyiG9QJ+c1vW8rPjfBPf9xYi
vxWkwykslizYm86ccCVGUXFImck0vcLhI+skfFZjcNFnUkogjw+EwLOXz2Bmpbfx
n+yBZELOa5w2laMDt7cLwbjNHz0JnLWs2ogis2sKUjt0SMRsmp8UYeRh2Pbr9Bzv
OwGofP48KshmID4KYpsZBnDKIwqiP5DNaQl+46x7VwN5h08ehfERdA81YN/qmrUv
Y3/oOP9Ur0cg2DiqqOrk1x0qDy1XrFohauOq+0ZRTEZF4WfNsCvOHfIgGtDyQgq9
Wdle3rxecQ8ORsNXo0OPlPkXO2BRRqxTHzNU9RfEwzFd1x4YD3/U1QH6/qhnSDlL
YC2AbmSjW5ZEEu28iSHfmXY66KNS85sLDOTahmEQsDRe3UC00uPCafb6GFt8qHnm
p85Rpf2FM6yU+CyROWVHOBrLapFdmvBFqHVHptWhBMDPcs6AIJsRy6uxt3bwfJq5
W7X9Kp0H5OVhOHSknQz4Rb7e0xAmptb500dT8PHTaMzW7FdSCebVo7K4Tfo9bAPi
RioOhyxl+vrmXeWhRQj0PcQB6LGBTI0hZrGt4qQF78Z9SJYzJS24JyIDQlb2Jjpv
VKn52dbDazAKx9Zfs/3UoYQ/rigXO2IizGbB6fKuDZjRIAghNpnriDR2efA3RV9/
3CEdpE1Qh8wCT4gfqAg34uIJG/NjnrriV1mVU3w9I0W08lp2CozJbb7DDOHVEDXZ
rVeOnMcpPYJPsyhHBlWuvGx+OqAf+WMvcGP5q9q9yHtvHb736eTvIq1hw3LwQXHI
rbd7tLrP0H5xuEpZcQ1sv+GWC40mxtySpPJHwD1WzruI3TSy8Ru25073D5Z5LVKi
uC6uzCNr5ERkcA6w+vdM5DA3zk8UJfTjVoF3YBREWq84+fjgY3rQBgiAPKEfERLU
7/Wj5BZryimwKulqgTBJcSSGdGHtpfdlX9aKDWhMdjQZHyNilvtC37VtbuyC1r/g
t/49xQTbCsj7sJjJRxQEyjEs8By15Bg0Fq+dm3PzSlfIX5V3PT/FNdiA5QDmkNzi
xfbMoaQIJNtstCRu90QZmjsqx0SQ8EVKUQ1WUe158U1LltmvbxHkWhU7JZq3ahpD
L2mEJyQgVqpVtKjbfGb6Ct4x7OfMN7nqe9kVa3bqk3x2wLGzHnJRUlCUJiAvm/U0
5tuiHIGre9Ayr9H1p0wT9xFCesKEVBBl/CGPmDHl7PmEJQW5K2mIQasSFqM9Gw66
QAOQvrM2LGbRN2Z6jt6w4Udw+vjJZtPAA8ny7Bjd48DMRvF037+c4kTLXiT2IsUG
ghxb35mv8B/5qcKaOV3vj+k8vQiRf5RzHK+ku7vIxqcXLHX4A4KnWQpI4FSVQ/ts
Z6tSU0L0PrH9hiCgmvT33rGlpkl5ksJ6Er5DU3wktd5Rr8FDvqIXUDWfjQNuBzRr
LXy7pQlTefAkiKINoVd1rzjJ3EMjpcmA8CQgvIAK/vF3yYw/pakeDNipDnLZDigX
GE7eBSihXXpv5UF15ry/81KnidiqA+3tMyPjhZI/1KmZjrqcI5WLKDf1SX4MTr3c
RPjgUAUbqfYA0cRKsGnnmFI0V0E9w3oYgCfxoSuvUA/fO10Xs4KY6CQJD0vlP/oR
zgAM9sFWkqPT/4u5Q9BvFxOn5vzJ1PAuon51Mtrg3g5Zw/9HSp0eItsmrPRgaRFS
1pPb90pK46UcIs9NnKYxesetqFWKag2AnidZGXd40gvl0fi0YqB7kpRFbO7V3Ltb
0apmHwS+PUAEy3ZWmzDOai0qrFam7S7BBMRMv0kRTVbsgE23ULMMCSmunDuqMzOE
rnc0jCfTWquJEHpYb910b1qEP47VWcdZ6C9foQxqC/J1dOzHLoqLfkORHXflsOj7
Er6Qa+y4nSoln+YySUI1DK5Xc0blywguM08E5iqCJRPbjAbRUcpkmhAamhSojjd3
8M6w+i/Hveildlx4PHssb2uw4JyITAWBZ9kNkdBRxV+ING+jQ3fd5bsCb+kVKnPl
1hGF8xSCH8jFnaPVG9XP19VE5YJ5hYuAR2DbZMAWGJWcyNrkW7qV1XHs/27ZvY9v
TK25YQbKfu0Puxl/D72d8FxrTSIObjYhd6XSXOvODIv/c9/+E1fi2IqplfO+LQWE
kpLqhOIDJJwFbXIH28tm3ON+X2M+CfqpKNFhQ8uK35KM5u8n3AMfGKeCCfnyU09V
CeZw5aRJ5S8qYRg/rcI9FDoPhdfn3QaDQEfVshikHs10IWDukRrTrjNUJtsQTyg/
IqWKkTLImt22Ppy2PyMLsuSvy0noTHBLA5RluUp0WMV5sbtSEeyQkvhdSgap8dWj
+p8GnwN9d+ZwYxaSDd4BHRBBEhED2IiLHpfmOOIioAxlaBR0GI8ADZKYq/oBTXhT
62yZ8OqDKqF7G2S3g4f1+9vL/DpYrChcKgVi5R7NfroSyS6GGffGMLbeXE9MxBSD
mJqAb+ddd/KJVHj2hsdsToffNFzm3/rNvTRRou21t4E1dBxg11HhSuZeCjwraquH
pCM0M3WDcLsoPciQS3l27wTDo18n01ySsPq71F02FwzHDEBQaB0MoUCHGSkkRTHM
yhKO4PrRPFWtSE2bNCRnawJgRKe77tEo+Gf+iiB+cX37AIl/Pv71qiLQmmXNDtTa
mIM0w/4hs2ATc+i8WpqQOOayv3zK+WhBiKkvP+gV6mUbM5MFHHnkURLsMcyr7N/Y
ueBnp5G7foUahgsXepCtodCvrPzPD1+NJJla/wk5dvRb62gb0y6Wo+YiD6iuxAfd
QmIp1NWVsB3fdnuzgaaIGLf/yRYbOCC6Q0PsdymNV+WrNK5MQ5+ACbZ6rH+eIuzI
MnCWlztqszNvGbETbF+A8HUibwwcvjEmaG6bxDtd0sUqjEjIjnRZZEr+IbnvLW/S
z0CVTK6zX9WVXom7yQhEWW9zbB0oEEpfx/VqZDbGMdJ19bvgckYZNfHbbVP8k25Z
vQDZ/IZASEb5cyQkvla2BULUfoF3Uyz7UMLv7xZbz7cFSajZlIhj47bDhvZQzqLb
fjX3reYaGk/6/mSVJpZ5Nv4zZs2YXCKB0XKLOm7H/5I3iFVmDx9KlUWNQwFH4+AS
GZOI4XIx7gAq1qLOnduUS5C+0h18931dm1gn+zu6g2j4RjucxWJJqsA1htjr5ltA
9yOSwuANskYYwbHipWKRkFjnoFS37EVKnaHYTf6UbW6qDX3nnx+YgwttgtYdJNB/
1xUo6QgseXehn9PKAWUMhwbdkbV348szehPbGT1FDkxGeR6dIdcY8ETKaar06rWU
pDnPUCZOeLpVNAiiBYnAhatWcb1wBxQebWyUx0cJ4edZHBPw/W3hb6UvRJcYTAJq
ce10xgiqE9ZK1QGSBMD/3ZIDb3XsYjhCvNJuKH0Y/mq4oDCUWXwBi/G1iN4H2MJ+
QKAYAaVBPk9iwdUdjo+Ncq+0wOdQDoY2mnRpYz8ElNzyjSOyV14SMAnTNXw3tf+t
SLy4e4p0mpp4hLcMMQttT7lQZHUH4ulHKxo1UtA3f90Xa01n7n4cmT6NOYC5bHHq
N9G3GkzXC6zazeecGf+5L3fgAh/PpldANrYsC9mXWCIXM5xPn+eOC4DlrZlVw8ao
HSqwsf8wSf8ye1w/suc+waacXGF07NMpfjRrwEkPot4ZjNmQ+L7G20l/oN/8ujyZ
hXUvJq1v8jcyjc4Hidkw67HzO4nrWqtwfQJSLKeehmS6I1lMrnm2rLToCHeQjIOV
wBY6O9zJlYOrRmKq4h0OJfyU3QEG+uA6OYrnx24pKxaNiLk9J8cH1FV+BYToClX0
F8IJok0bQDlnrbwJ/9ub71pShoimOOUBp2vfA8yw+Wp/R/6P50Y1a7Y5+D50zJ8I
C1IeHdaFvy7LTGZtWZNIar2t04dpZmQKZkcb624LQ4GjdDc/xBrsd3PYVpc3zSkm
hpGKyaee5pu1acYNWSa5MDl/UiZueodjaAn7H0CGGt01NFh+YhYF9bGFOf/PuKXd
FE2fkh7FjFCxPuy5vFWfnyUeOfL5npGVBRD02O4GwizNpzRl7B/Ab3zuFnwXLrKT
m0/DcEahCN4t6sMe8W9jql37REKAA/0/SotfKb1t930Dd03XD+ErHoQMUvaEUhp5
xK2HXL7XKXMt58eEaaY8QRpI+gRnlX3BNl3C5r+t6waxAxZdbMI2DttZfSM7NV+l
rNH7lyR9dCyetO/Tgddzjr3YVU0isccnw9kZGlCfDlKI1iob5dI4UM8KkjTBIVha
cg8ePAWIisxzvkCDjczuLjEFDeubKp75DRWbyeMim7SCpqrSfy5IcmluG+2aGZw/
1jiyDFjV7jQA7n02n+G65PnYX+ys0V/CZUkLAkjOdfnPOz8HuUH7jwrwCZePiWKQ
180Up1RZviqtlKkbU23MKqmpWyhQlnqqHNW1cvQrW1bb8aGVn2cENAOW9iEMCAgf
HQkEDNLzUcpwS/IYjdvwXt5Lord5Cb0P7LUUYEDPInNdeVBRYhIIuFDRPJNw9lO0
7eIJ1iCb12D0qn/xtoqwS4SEBOhzYR+MjkOg6YiuT0APLyli0xdGh8njwB6jnn2r
Bd737GeEw9LP9KTEcbEqbcIXdbBRn8LdWvscaoizaY8zTt+yw3D3xZfFmxozV4re
+++ZGKabWR9Gd2tDBT3g4owXaRchGoRCugS4Go3DJyzRpLAUemFxj9I9qE4aYvd9
POGCPBDxv4urNCVl2FyNqN608YnIsTMRWH8xNJjWFWA5QlN6toQLHOpKmZ/ZOKSm
N6hofCLFASJ+deeH0YHBK3y0T/vWmv4iHPZOHOGB/WIXUpCfTZKcClflSFoct8e5
7hPpemGzQTxd0l4I5wVOcBW6l6kb6kkVjeGI6g81QpYjJLZY112lmfYbzv3h1BhV
S93nFidHwV8yh5N1L6NrQ0PNAgqvaWJXqcarhkzLnHlbjrY9xBVrXD5aJOkWkJbW
oiRfbpudqtUTXhipzSoNS7p72j5iCn7DmNAGDcnogUxATmjHyvbMTwY8jkvQweuX
R6Xa1m287LPX9LzcYGBM5f2vGZzxAgFZGW9fLqid+AM43BMBNJ8LcU8Qc1tZx0q9
JEnvU6siZt0SqWn8B1/El7ELiRdQAL3tW7QNqEmwRQY/XjFwSGGcozhqbTbZHbNd
GNPXm3Ky57q3ADG/zoWdaRvcaaN5bC5/k1z9+pnzg6kzWdV/1Xuv/bQQ5M9/BO69
VolEIBeX2f9eQeV/AZmKAkjy0kCQjlil8aLY84Oe5cgH/xlsaNxC1aOtTh16fnCz
KfATxpOS+jLyABLQiwpUakZVbsKVgCw6VEbhv7pSBYKzbM2SvXfAgPzgJRGNPKD7
XSOJJzKj41EnwvxhovTwDhl5eNgf/dGj/vPyyVz1G7UjY1yB5LMg0OPnBdvqxjFv
+pLUZ5GgNschzC1xFm7ymPlnfimCRN9eqWuWfnEWzeN+J5DD2DnabsaZkY2WL0IF
XNh5cyCwluCsMEcS2KVyp9jSqPyICMsWpf+lsATgQwATnhwQrdKhE67I6fvsRLfd
WvVYZw4yTaVVGO5TWf3By5Z+0sNA0bSB6jShWU92bMMoV5A32JClOWEfn4AjY0pe
4mp2XE+B62yYsWB8kvV+o8ZryYadOD0057poF1bW83oXSPWUfk/zUscbJ+Vkggv8
TxXbm7O/DRikmOQIz3pa8GwQribOq4BCQQ2dHTgpMCDi0BhPuqLq/qwPKGSMW+wh
H77lsMNHjV6gTMkJPEoBpe1Z6ljbCpvpUGfvNkIBQ9uKB5axjzsdTiRrNJEvZm8f
hJVzhSf6pbcAM3JWF3clQxP5REU9JCxXX1hypKcPMnzavE8s3AhkHZJVmv1hKdck
nfrLxRNjCnZ6NVlrzs/PvmbHmCaZE9fQScWF+ABy6xqSJaMkCj0mf3xcGx68iNTp
SErQ/2Lojfi6rAgaC7gBCbEUtIW9XZJQVpc59Zo9RNeXPdIawoGEiuOYaD84ytPh
TyUmjtftcCHVgZ2+ElSTP/JYrMaffuhfa3xPIXIIxfqWW7jsi3k9kOCRuQzZoFfU
6HM6dl7PEua1Zip0WdY9xtaMmvmI8j3SCOih/2cpqfi7Lt94tNVINm6o92VtebD8
GooxVtRBUYBLRZVqlqnz2XXwkQvvnG2EbofLw7vMakA5ObsszHjWL+eEZo4xVgz+
EzDAV+8bBcqQhKtUvqYGtdCPOPOEtwdpKfQC9fdKi38o0M/xV1f4m9WqhAc6XkUz
TU91ggd7ZBrHVxnKoC1b9Syr9C1CeCbl2Cb4ieYhk08PlQmUG2CpX+2fLS5M3B06
7h4GwXMCI0wwHc7GnI25ABAcT+Z572w6M3o45gL3kpTiMqCoksxaLhCN8yVBY8QI
sx/ns1apCqMkBsoq3v/MgIbsTGdvpnIvE0eQEdM1fQgat/3vgzTiw7jwbDi2O/0g
ZIucu7/Crqv5T4PGcLR0cZ8QIxzH59I9v5hkz5Gl1+ioI2GsYFeHL73cB6WBJvzM
itU3HLPUgEGXSA6ML0P2GqBYAOgiqUCG3Kzn2T5dz69S4+pmojBYUcAOup+gQIaO
wgBmXn8qRePRgEY5h8IfQzI6Du6cwZ85kUaD5bueAY1tlmk8lVBqDlvC82W6cTke
cCHvNDVK2G7OJMrl6oIGbqPRIlv82QnwayPZmd+wOBy7e88vKoS6EkxWi4JMcH7w
HfWx4fDuvQT5e0fIaQz2EsIIGThW/SyB07p5RHGNdvbVEgHnO9BEfT1ne5XrLLyY
qdRLyYKG3uNwrElExZOUUeAkNhzgyfZeHujqi5lWi4ikA+dAGIdpQ6stqNZZnn67
XqP/vMMdpX/PLHDb54fHZlvopmnqvAueF6qi+gCYfxbJ3A3APsaXjlzbpewvV2Kq
02ksccewLtPgU97/l667qTZt5AhuBFFJ6wOts1rUXPCWmSjqo/RPB20cE1HGRLrq
nhE+bowsyd+mFRhjYGcsAdjsavk+AoA9E+KRGk0HoCv6AN0gmWXPIEEmtUfq3amR
rLL3doZDI679veD22iRtKAjQtYx1SN/uqWnPl69u+JUQfNP/ZCPeBUeAYW8PTRfg
s9V6IzFm6W8fgTYD9ifAjdPGzKUR2Plci2L6R2p72sKoxqti1hgJOujw1KB2fx6K
5gLLlqsjZHSg0Ohkz6QILAhA0lJ+IyRZ9cw/K1uOi2uTJ0wwCOQ6iihN37MJ/tiP
oGER9ewKVRJtGR+EmA2WTWKspuVYnoYSptRA8PIAGDP27+CwwMyYX1nvjIJiFcAZ
C4j0WM2vC36Frg1CH9Eod6l//LMGLouZVLilLVje9pNlEuFIYGiEYjWmgnex0wYD
PzLRhJa2xOAgO5EsJJuW7PGL7aGS+4KyvVj+QedayGAgSUGxhTaJui9YdFTEbybJ
8JszrnCOr1lhdkOU/arSKB4rPEhbUvks4wBrKRCYxouR/Kgka0rnAUWRbLjEV8G0
0tGYdv0ocdlo/P7XIbeNKuaLf3uLDjPHlyRfuxOZaeP7jFP97EstEQZBljoMoSrl
UyECRYqFF7rfy7mcZBxggUDhLkm/JJyt8oHXkIPzoQclZ8xuyKZP62ggVR4bBKy+
RigIW+pwUuQbOR/UVC7qhRhAUB+YwbLWdh6CkeFSqFyqJDfgBF1SRIgGEYCMKmkb
lQZC6DKRclHet7H/2NRt2WII4YU0zmrTUMeFHJPf3bOjirq6cLCEL81mtBeym3gJ
WNYKnuUorncpDb2kOySt/kuQAKYclMZ6zE/BdKtvDoVetnKyvL8XwKE7b8F9lPf0
nrUPLf+ub2ATlhA9rHebkUSsTN0uTS1GAFq9B+Cej3XTqDcqurDMLvBs1wVnDcDG
rGsaUKHXX+De8Z+Wrrvrl2tO1q1TYOUFMjliuSJExIR+Phppfh2AiTOEwcRwkUT2
f356WMUNDoyuSd0t61+tUqselsvTss1xA3wxqAmI/wkGc94b6JqJBrthFzZ5CGvP
UA0ITbEFLvozAaDU8OKO0JbE2v+ERUIyGrjyqcTCg+KD8pxUWtKuN0pA0h/GhtHU
bPCXt5bnScj4/PgsKnrSSf9HGnk1mydHAS5nDk93xH5dWNVCJTCbQL5iPYoSMlb4
X+PWMbigEOfIeLUP3GE3m0/qe/EwNAr3FtPRxLwmJk1DfehbwR8+SQSnCiEyRBLa
1DvC0uKErYdBAQXRFkbL3I6VRqqbjfiDP07YH4MMCPfJvOZ7a/dsre+XdR5ti5ok
pvMGUt1Budp45IKb2Uom49dgEoUES3dLKcIS7OCu+sHCe6OcpxSWX4c8+wc6wKY1
5VIiaktg83az0TrVk1p56zbFDJE1e0BQhtKPnqfM0oeBNI/hMfmmxPBVaLcTPKDM
UAgSN3fkuWPIHEwsxEy3NyR7y0ojErWF1Vwg2wj3drHTp74ttGifu9w3Ba2kr+4K
0LaRgIKlm25x69NwnVIZqzRkOWoXEpMK9aH+w6E69SiwY+QkbUh4o2L1atvKsiMx
1AVO0svMR84mq5CyJUMtYOT191PxelOjBHcQL49UOlg8uzbESqDcbjJmeIDpEXP1
7AWeDLb2UMYkOKzgXbKUK6GSrrQ1gID1UfupYVyJG4jfxEgObgL7y1tqQKYlGEFB
wDSJTvaj8wk+Qc0eXkRo4FWlrMRWBgCJV8rv6sVI1WHpF25soHygIdI0pDOA7aUC
gtwNiGhCyymi47gbrZbtKS+lFehiFgz3JoBjLDG+/+m2llpIHi7IJo+GHc//laOv
bT/mYk76hn6Q0sl9UHCddtW+Q4Z4PYL+0HxB2o42rCQk1FGuPe9wa0Uu9niVaw14
V41wGMDiem/5IPm9jrTuE8Z0k7t+K330J1YUk3ZFg2ArAYjIDzvN9XjDVCPGKvPt
4DxPHIKwH6+FZid0kihzHGqq7zzAZhupvJqhvxg+mGKuyXbjHt/eMstBYb++5+2X
Ep3oN0bjcMQ95XC8zGhS9vTWd/4R+e1lIQB7hhz7fwZNAwzIlCFfNV8ONq5Md7mw
byd9DMfv2ZciLeClWMCg1LzpBfO2y1CWt6yhOBG03wNP6Z9LhKfcU79navsiMC+e
DimGltfSTOdEKIS+UUSzwn3LOhFSIW6ZrEiudNY1GYH+hu7Adu4zne+4d1NxUbzv
/bP/xCSnGaSJjcm9wgb/SZ4IK5QiNJl2z7a1Y5BPW2ODYomgjdks5/rZeTb2gQb3
ZdmFwgYLsegBORFVisXSCl4E48w2ky1NZ5oNsP6BdXg1+NuwnC3mpUaY/JnJqtm7
4vdFCB+7QGrkdGX7o53lcK64csDy6sy3W33w2Amm00sf98IfjJdtnZ+MOD0D/jUp
yXVv4VmIhOFgk/Ot4hTHXi/u2Ie2GGqX4Kz3xn0PK14+ln1PhPnoHBGGw/7ejSom
YIm21zhw58spQzZtmgpVAPsQo63Y6pu1Ef1juLf9a+yF+xjyMRduoW6zdrCem+4k
1LnAmqiivgIK/JH+tAEk0wkL22yWnmTf/zdr8DbzcfqNTVt/NySC4i/7ulCf/wsX
4EgUq3SxYTae173p4I15VGHBiX3EXDHRxMhOnpfTLVrMXntop/mWbznGoH5+R15o
57W9BBvKK4pu4R4jb5rFIIdGKas1NtYtIFvC8TjWRwZZigMweadJLUyhzLqmsTkl
oJeMpf38+xVLVwshG0eECb71Uziwyz95n0OzUOPauLq1tErMQwowlLN6mgze75fZ
ZOE/wWyqr9AYlN+UcyN/8oBbwk/PWQSDbw2j6zRIHmj66DN/CORnF3KM+Jh1kpp3
5mLDL43jru6utAUZuFeLffovM9hVJ2t3sMJkYAcI8VvXYFjNclhaXCNR5S3P/M7D
dw9CFj5npM3yXS+p4GGoyvsRGjBQdfpOPSSbSyf2NtqWlPGmr4LN+wdIjXjRbGJ4
2vcIFY0eZ4PnLA09cjzCCHd8b8vaBy3w/3yxtAOG2/mU+qDiFDNtP9Z4j8A/h+ub
0PUt1hp3CXytzhP1hNy4JYRFOODOyr4XkGG3J/qDXkzYk8R8asctC3+om5KlZIbD
jAVFe5A/JZV92iEC+WWFY4ZIXP5DtqONdZMgPxvnkRsLRXls/sSOuK0V9B2HGtsD
UAtPCR53ZXSb8/96wY025GcrTnHfApbAoHmoKiSf91OCACyhDHyfFHuSPP54ZADt
TBQh2KAe36yfoh8XlUOklfApamJUxOrXnBm/45/GRDv828TsockpkmVjD/XzZrXC
AMMdXNQYu3KmQoE4HKbriU2eHPBPP1MlVePSQJbjeRyrycC2a4zqK+Lek/0QnoYJ
Voj72VMyQJrhZjX9B4h8eTRi3YnlztcRPt4Ccu9+y4/NcOeySzpLwlHdDUUvML5e
T8bf5JoK6J5PUN4b1KSd5O6F7KNnv52oB5RYxQYMxc+w3XhKmezElNS6niRVYHvz
I3sLH2WA+CNqHMhb2c4hkyvcwHXE//BQ31Z1859tjv025KhUfBgB84DVfB2Snksw
wxAVTKEfwTqKMgKLzSb0gLJc06q2VmYv4VWZjipF+SIDAiAY5aJ4Hi1SPVgiG0m1
iv1wzLfu5YbJjzs/AcHbyPezNssgnFbwYXQVHNz7hL+OdOrFi3VnasqPeCnVq70c
7EXREUt9JmRFQukVCOaKPHtu5f0EHBiKQU56J/eiIDI/zDw8cI6rjkcWk/095vCz
zEG0ckkgMZ6CzgI+00bg8kA0Nb/IO5FORezf6mN78/seNCOsRwaO2KHXshivqwyf
FDI6wLKF7goS8KoLsIQ5qK+k8QYOqbBjX262RBq3wndwWU7lpXYlwCqNCaXLlo+1
Uuj++APDSDyxV0mrzgxD/9ubnf4934DhkT0o5bHbcYs7nHMOiOnWp+l2x2abuWXy
Q/TYMhqYgvtzDqc6ASC/ui43VpVHPykV2WYijaqb+sh7Q9+D30U+pznr960X/I1h
JYFG32eHOayLDfs2a9Yyza+S5caKWM3slfgqYqOPJD1LCXe0C3548z9l6S8pu4iS
JghlcKv1a3QtJgZ9AFukdPgPu96WcnfEm6ZnzhJekVsQxnJMAL+f1k2KOWo/bUGf
SjLYyW4N1xqnWA+UemLqEKs7UZn5DqSklFxB/S2EmM2g/KxpkhXYTJ4jVbtN4DKH
eafTs9vPC9Cv0kGW5get9/qPiMuzbKf6hXcRqyBwD4YskP4pMApp2O1IMnqxUKhY
1/99ZknrDmlLljY5S4IdjDUFVMOTvz/nF5O5F1Pwy+GukS+B7AXWQYjnpXuoobQS
fFQIjPbgbV7VRbjEM3JWpxo+YhTDfwyyKCgstYRBhXI3/6rFkluXTFqR1HoSv2Zm
+KcQiour4aLGOFzSUkafPOebKCaP4mNUK1judw7KTIB7VWzE2exxlkV0Wglxt2sh
yYb5TRel1GLqg5Arv35iIBMjiHES0kHj2WDWGZvNhJaKnKzRtOb4NrIrsjmHPZ/W
sIUrkSKAszLebk1VfBcuGG4Rgc7d3KDJM2F2IpQ6VZ4k1HxxuVzlGvpT8/oB9rPu
36M6m/imoDuRL6mpN2jz2F1eFDc20KlBQMIz0aFDTq+xB2V4c8rKhWmJYM1yVxNO
VnwBCSlLAAoRHhv+HrSKy5jYOqIBH1zpkkVkVjQruSg8G9auxmtr+MBTyPVcIBAw
TOLIckhBrVYtsljVirQih+bSlZLo7oforopmFSaPHM/u2cWa2dWR8WXt1S4jszZF
ONcN3zK+2YX9WIIMz1zHHXWFYI5u4s5y7lfPYe8Vh4mo4HaZ17FikYcKen4Pd1zX
bRfnS9bSxDXK2Dvj6IHJG/pv/RbXCQKehCU+yAyI2ibbsFxuNUTlYmv/DzEfE7nX
y3IIInepLeJ/OUuZyf6a0dNQEf3KvdQ9uFKjkJafSNnuB7jFzjidkzWCPmdPI0T0
HfSLzBAUH4FI3CyxxjzcDTMxcEDaWIEm3JfoEiqx/jDtgGSaQgK8pWQOxthaGYsu
PE1dg+iv2zTkvP6Y/2dS3rgYdjGJfGwv4L4zVPJHHKMdRL43Jd3Opa8xJa1Qyp9Q
Z4uFuy7c2KeAr7pFkuDw3obLWxLVNIpxjQekZ7sywWioLis6U1W0ARfp/fCg+FPx
2MW1fZwjbJrbxMy49DMmMGWykwdsDwvk6K3iw1R3xhdvlhWUQ76xTHLQS6rZt0a1
vP8XwPpijPbtYqc+ThbHwRH2Tt+cnMzy6NAVJ0mdGnIshE5hf0w+qpVWTSVqBafY
4iE1OMSScuePIXwXY4gnoSYP0cnaT+Dc/sOLvFgYRog8xOcp/olohiE5snkwnW33
o0/EqZJdC49RxgJTXNM12dgSuEviXNKO8PPDSDDXHFZLij4iz8WwPV2gO67IymnK
nDk5NK4WtDvQ3pfhXLjEn5oZU1KvwZQY+pNlZFt7hQIt6qQAh6aIpbE/yFcsM8JG
V5Xutm8blGzwYEMXEyHmgxbXAZdaRPOE1YWP/q/JIy54GdgCXl3bELplK5Ako+bz
D8vmu2CKARaG/LFDQFyGdzkd6uqQLNj7nMR0DxkO633Roj6h3l7m08JCw9T7FA+h
Ixm2uFNSwEWYiR9rJ7QQvrKXR4NSo5f+LUZBVezWIDqMpaTWr3925SiEO77ad06M
aJzwHJUTVtYH375h3/2G+F2MO3Rnu5LwDRjxywPysN2Ly/mA8df8OjPCJszEmt5j
LxxvqU23r4525Ki2W2QG5K6ZqbuPl492Au0sCIaa23hIhyvlYWPp3QgR02YV2vot
7vzOWd1UKmgOI7Jeklw5GBsadW/9qORyZKHSQScOrjMS6+YkNPyfLCdHvgBDdmpy
QClx+NKQMGGQ533VwrKtw87uhNNPh3pakPxBbhNayJ5WxeiTv54cGFPQp629isYC
DoO4ZLHn1/hBrnEOBsXx8C7MPuaH77YKcHg2rNqcnLqk7R1oRj8luL+pkwXH6ve9
cuSqSHM4nM1zsdiTAGq+zFzGGMoNMyeiZ/8PhR1GushUGgbu/czHbVWxay3x8yC/
WvCtzy85VYa3x+jUIcr/ce9nGBexygNlbQqNWRmUYZz3aSyM7EZvqKoIJTSlvEG9
r/mjrsHDyvNZIa0w7/QxuzxcDdIXE1tfNgBOM57MTlyehK16/QscCXdZqIBJ3syj
HWIKpDRTYNCann2jCxvWX1GLKAmWpkHmZyVps7KmCPIeYWM1a8d61FGeMhcgWu3O
hya7oBCfZ1OTbB3ceeqra3sMzLJcLlutcBAsxJNpAHJKbJ7z8anWJNzl8sycC8dn
zgfJY967VF7l4HOm1Ph13L2eMpOJg7CdtzFQw1HxuLQvKwqsUrF1arKbMpauU5Ly
VSYpXwp/W6vlHWUO6HNCi4b6jh+m33F4mJ3rODFO8BfxM/wB3EE4sgd2wjxeemRQ
7aBh+MV/LeGNYzqQv0fnLdg3KXINx+Vw70DIOgEtFy1462r1203bUeCye8bX9CEk
HVfLrpiFBVn50Tv6H+N+eThOi5JIxHwlu1Wx24nw6ve/KhTXUhPweq+kyHkAPwTT
JmcimBHwxPGdbNZcftamHAqXWglNmTgn3WhrW6OImEy6sRBp5+K6RXJLhj0jqsH3
go9z4dMdAw87FQoJkNDTQuZnezDVpW9ZnYbZyVI0VJdAAi3gir12+EgXRwOFBArj
zc61xrapSdU6gD8YTBiVVeSeJolpgNlkKF7EbOP3F+UsoChx0DttDrFsPZo0uuqn
L9CuMSoOeo1ShnnbT/CiyUwEn4lQY/BWw0MA7hLRe1fyRYyEEmnstykNdLCveOMM
PksAAMOWN9R2FW9xvn8z+1N7fjweleucBbilxicXwoDBtt13CnMN4oWdntk/2m92
+nKsAx6i3daKVyluQI+IiryFHM4+OZxjzKa/+tycZQ+a/13IjTc8+na/VW3Q6756
YX18LIK/42/NLhsBlNJP/mLfN3RhN+AckFFR8HL81ldb4uwcEcg8H/D8ICuVWrx9
RyJ/Bqomv0Zk4hZobdyj6g54S40+RNh7YES2HNf9a7UDoP1skEH2Uhau4Usz5ICh
PMCNpICcm+3+dyI9SN/5f684J7oPs9dwnf9FkvY6p9d8lAROoulS+nMYtvfqdqNS
iXvrD4FKrlXNjH/GpYVWyxYQ0jVYaR5xtEy7mBU03jHAOzom2AkZDMeo8UDzfRsz
XDrRD5BRhKmcmxaiF165pODX0ZurEmoTG6YSxDbtF5pkcNXCpClVi1OAdSgwM03l
JL45umJnEQaxBU6UQ+T6SjzvGfNC4joBN+rOVa1FY5zqznt3uXcUbtzKxs9pHSxe
n0TSH+FnxUS9ywZeUpFo3YmaaIBFEHUrlh1+M2TM1QqrLOPpCUPqmambo4kRqTa3
wobXU1eF3H0xu+bXzedLMsBP3JuDVH905PwUZlIXXts3Jyo2/pTt1HelPSyRMe06
GKkgpUYWD0qfBoA/XkgMenfC22t4JMBHegHp0HDg/V4n9T4vvhLsjxzaFoTNIeOf
j+zjICvwwoWLgb8lN/EsNRmZexZZc8f5TsJ6HIowjCwWUQyUUpE1ASeIur0mpckK
OXpUckCcjv3TeW6WzrtBK7s0JedEH3U2+MpgpPlH2E9b9mVAHdUZ+uF4+Vbqw9MO
SmBZ+k02M9tbiIg051Su8WtrFoGgccCkEHnJ7YrDqaBGHN5VLJNooUWCTiuBPkSr
+hwss9b7JOgLKOBKTS5QNedr9ywtqQC7k9beE4IDb3bHdH4k2ST1ObZqT624a6ej
6JXXqDo3pAUidQPJP1z1SWPjJtCwffyH94qul7sOWn/ujHPsSrnOX3NIimQ9AGKI
PwQmGXbJQKRG0phhNL2wUgLOgi6zJ79FnIJSJHXqVczsmOkL9vE2LCDdlFuk1vNb
sij8qnM2NepmZOGgJTaUBNI73vCaCSePFRVJq3J3UAa3gOLraDuYUO7f6USl9hSU
vwIaHRT1OF52VDnDH3oBMVIViikc8pJ/psbLqq1wNLIVAtiVqeeDIGtIjk/y811N
EzvI4mCHzlE0reMLKmmy1Jgrv6d2i7o18LHunLnS9W5UWmOiewAkvRoDyTPyznZ1
abiXWeAlpOOYNBxAdUDjLszpOuegAAy6Ln8Wg9Zk73Drm/gRWhaIF/o75TV5r4Zy
V2I9FnHj8hDl1VJXjH6tvhq/uzoVdcs3iXCtQl7N0uwzwZMm3jlG9tmMNb9KpCU/
MCl/W6bOUN6FG8i1F/Cw3EPC356ricikojLH+4qQXDgRd4GA8sW9KVI5obg/61Zi
2BmpLHx7zxFo7m7UefcAixAPb2sVbl8jUXDIaCrj6e3kiHf+S5C6SY1QKb8ixf+U
PwRAIVo++0n8nTQoAuRMQRMEsM42Z8C7knBms6qP7t6euPrWCKI8JwMZlZ588ghR
lIHogMLuJlA8HD6HWDijW/QP3xn5eVUs6LtkgVTAvhw9Kni74q1/RF33baJPH3aE
pEmgUvfmigC9IZi8iPeugz67SIzU/qp69V83TL/sGi6grGC3VrUGUS9RVGBmMSZc
xI6nLNeLoD/hFGF3GnrpM1+gL4axicOCE7nZNl7R6cs+a/6Z/VBVHi6ay4GquT4f
LmJzhzdPvFj8YZc+ulT9jDggOKvNXl4+CXsitBdbwl0bmJq+13p39LGl1KOBvAUu
YuqNpjb3n4zv0RNnKAt/NkD8AAp8/q2xqYdjm4Djwr/aAP6jGOjg5xcTInadNLDh
zVlrWFBbahd5WRzlviCVAFaGp53Q3qTH4pWSPA48j+O9kfygxPf0uUA1AnKr4W3T
fJM/g850ucg+A9MpSP0uQF7rOSeIsB1APTWI3D5+VMtUJmlulVHfqHGnFQjzn912
E3Vn+Ia+jPgLoZ7t6MudMPG4k42Ahs9uH+nwQmW87D0zwhMQP+aKR/EuRQjSmp1L
HnbDG/w/hqfFlaZGWms8dKr9k22E2n/9Vd/r89T+yGCZVI58p5zt/I+dpOfoiYn6
FuEikGBaHu7cHhj1h1Q9YqXAglBS2fSvMJZjZ/HaVF/JGKafrJvFaQZzDjnfrl8g
5rVENRS7dre594EFnmche/tZh0Kbyb1FMRdNcYtcldxwMEhjH2+WGXqZ7lLLD0Ir
okKsXzp7oHWOhS5GOkXtDBNQq1WRCZ69JWH1sI/MvVCwsqLfgUwTpqUi1AdxmHPM
TtSI2UUsRf+DR+TwBdqvJBugwaIpjjsOht7GDv4PZ9eJeS9t/+i4E14ZMzsfJ1CL
F+CfcFVDGBxZFBqtEkGN9ndixuHymqtd+rmbFdoCsQ9dLAjKsiYEAKj/m6fR9HZl
2QKGuUh3dt86537TtWfjiMbAJEffZpfr9XRCdCaO6F1Qqbp7fMyqrMk9o0ypw/8J
WdDw1VYkRnlLrdUxu7T7IUYrvzbzJbvccLD+hxefE8e44rDn4bQJfnjjHpFbmlvY
U5Bcc6rJKEt354vmnPmsLB8uN5WAkmEo5vlMzDnfE96CMc+oVcteP5hns18UoYeO
Oa4DDduIxLYLGHKl+pa3tP4EGU3HE/pdRyTYDD/+S21z3jhVMCrqlFskJjuc8W1V
aMzuXDN8HBaVfu6PBCx9XBdnSUxr/Oyg0L5xSaY3f9bKr8Yp9wBGzQxd8NZwY4+9
IEo8dG9w4wt/H55GQntRXOlkziF30eF+O3XB3Lyq7AlzJEx95rXpAxuDAC7z2ZYW
2uK3Ht9lalBPXnTvkEBUucaS9p577e0cjc2OGAenpwCckkNQJwVmThVB3Q12CKGb
M2IeVGbgWWN8nT/uSxLXr2745dit/O6lDM0+VO24V3ZlZwvTa05YR3Us91GxddKt
f7gTkYImc5FhNEC3h2UYGB7PUgnXfJGvLt3+vjfUzO4nIGru1mInDi49BS2qpM6T
QZP5V/6Ut5RwTMYIDZ4WKMwrjp+ouOeJjgcq/sVFmbYDJCfvqqtlXRajYvn/pbdD
PIsTMTOx0dD4EanDrMtCYw1CkQc89fqpH891OKXowjtdEPf2+q9RrRT+IbLY94Kw
/i4rSNpFfl89bQ/+Jgy5DiPrgsWDplUud4ykyBRizpmgBD1E4Py99dMayMRJH9P9
TI5V5CxP7XGguDYGg7Abs5Xh31Dn4MwAntio8+9MV/fWF4cbZDvRnfjO1FPCXY7e
16yHuZPaFKnHdQ/0d5RpulGH+2OvCvYI9iCHNIiHUZF1tdrLgIjj4u0HNq/Itgr7
O0kUHXAy0pckuOR7Ks7xzm4K4lqWhFVJ4yPGQ1Skh/JYKlltWeaOSjmr41e/xu0i
aQu9nqOz0k6CdkFscdkF/WpcLxwh21RFlLccLtCGjEgS9S9Toj1Anz0RGEpHq1hR
qoqcX/e8r+6U/dTjW0bi1INbWzXlP+mlyZlxLkF/EkSKOCVofB4mWZHn5qT7zYKQ
+vxQBJSa5ZkrNDz17lvF+bg6Z1L1XMLT0R33/9CMpFTvXCYu3o6DezgkyRSfcnq3
PdtoQjeHAtYBVlTor3WGwY2dsmskyIyCQTcfDa4AmK9xkOSktiJOvKxK4zWJEz2D
evmW4JOP0gxTo5AlDl/UURu/bU8roH7tb7s4kD5S2RgUSQQaeZ0sIAY4oiHqQV6A
KDHfJ3tt4UtciZUtNP4XDg8aVkZLpfl8OOzglfOKfNSFooMgHNGQUWxyIbBvulxt
ekP9tPUK8CYJJ4LIMJPHg5k3uiX8FblL+i+FVksHYZKot0N5XEEt92k05Wmt8D+k
i1tWWEhPDAOfeilF9Nu5CO23iNZNymfInID6wGCByNFd5LpYtYGESuEszbwWc2JS
klrf5qAi0AiQIlvjYtMQKs91z8WrBpft+fspqBjTaAvriiH3ZCGCgv0F8c9JzMOG
JNwyaMzyHzoaX4abnb+mgkEzJWawVqUS/qNX62LhjJ8Rkt7aE91bFj/Yydezq7eZ
8eD6y+DPKut2HlOuA00+jbJVwOh+44ofrV3q4TPCZVzA7hq104V5Yh4LkKZEy85D
WG2ltnkY8qRaG+xF72cyU6f3kmhmFgl9zVvEL74hF4Q1ZlOzG0cSyNSZynyBjZMn
ifXo1X3M1xXsJZwAXvW9LcM66+R4McAw2f+XK6RiiljD/gT5AD64K/iI2SEtbL6r
2gd6sAH9ODteQX31fRnkA6qVtMrL6ribUW7VxDj2zof3OXKeZgA5gf3/Bkt6mIxe
qK/aqZTORNbNNI0en2nugRlPH6k9AXdIlrQ/dN4gK9i6LDWHdOUf6+S5ZMMH+epM
VvJI7AWoielw213bNgq7B1ioQCiEPf3ZcsB/4F6Xkq4nvAewLasmDx24seN0+gst
SuH/Dgb/qoOvMy0cicZs9tlzDEq04osErTfjWdx9GJFObjn/9YK42ZzBw/TOPEea
yqydfktVAM+eyORohT/dMw==
`protect END_PROTECTED
