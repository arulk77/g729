`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JtuH6pKUZ9/PnzMjzX+mw6bMtdScZsXZrZ4rFIsvdp33oj33yvLmUo1b5tjWRm12
3DNmRz7LbIyCEuTFt6ABSpMH+W6k4EUXECG8hRlQtZc068Nk5gsdcWiY5AXHsdaN
fdOqBEUnWKlBjHa1xUckF1VTeqqzR6opsEpKRBAyeIYZB5XALHDErUWFQ7EcS8Pr
RE/T+FO4WCzoWUABa2/VO/mFajiBOjt536aO5bJdxdkEJkCz22bmEYn3BQXuRzu/
HgXIYH785PWeHKzD9sT75T3ZvEN6EqT4MvUNxEGOgb/3UIeZemZvQISqVeoYOwS3
92VOgnZaIonwgCmtksYBwhtUWBzw6pa6S4+NY5Qn7kaJBvyLhSeinafTVL1xdex7
wNno2z58K9y7jtR8AVebmD3Wp48Yi4vpU6wxyeLvVeY5IVlm5CaEbTzfsiOBPZhm
DlxyGQmZHXTY26NWG0nlXI4VMt2Yaj/tgFSNztncc+NKjmGVLw30jcPIRSoBHGaC
kVEP6BvX+o0CamRqWWzqMH+FbNHbyUgznLMf8/CvKNMnE7jnj7JNlC9FjMCaECDy
xvHB9myqJuOShDLNooyvqyXNBDkNc8cLk8wEqJMUmXTNQKO0W3bAU+JPBKu59S3K
9sz1AX1wYqdzPVjY8d7W/ypCjT8Jadqr0/PGpzeZoUCxDtf7qVE4ByMXGgHMUmiX
fmtRofDXGbLLK0AYajInAXLjjvllkRhnl/h5zb/9pvd8u/pGgIYYQpjKkHduPirx
bP+b2SruqGLmogg8ixSpOb+oZHmYjZXCLFuaYDgHOd87G2+n+nTLgn+CrsBLCuMP
rwZBDrFR16MWFHBKOwUiJBQngR008JEvpOny/ddWruwL8859qQot0G+BitbadmpL
eO0vQzzVBCpQmElZvuvPgdOEZX3zRNjoYhPbFf+4bj+uLRLIDgoUjYYNUfisZfJs
mqg0+8giUiP9ui9cKMosYumE0qeaDJSYSlxEzcP/e91Ix6xYLLDJImroGHPE/i6d
JGwv/lFbuxvEmPx8LqLMfrBDAhRnuWE4qooIv4Dh1agR4ufA6F/B9Hk/AVew5BBr
Wvsi1HOi1bMBn8JW8ruHCE9Nk/z+GNf0VZHJs2yHSf3dAD8C000RU1DGmvh8Xa5m
nhOq1fzG1F/ATycMu3OEmOfKtGB+BCRNLvH+ZfHRtJogQWFcRKBHsY4G3fq0sgLt
CIArWFfznljl9g5lzgevBJJBUdTw8CR3iD+6Y1nyU7ugm0hHzhj1MVTzBh6T3llj
lDxd5FAHZZzSEGy7o42tZDTl1hHxP4ccBWYVQyglThjB8X6bfCA8ZVeZA2TBzgz1
PH6D/4np1YlW3Q2/Ck8VeCEr5+wVMo4g0QuvnScNMxrpKfVSCntP6s0pJwnNKF5x
WQOvg7YCxydvBBjpgA4Cn5fS8549wNwZgkNykuJYv0kzjnGEASlQfIQH5M0FMnQb
Q7OtzHQSaCgsz0jbWjxXABnDdIb5YhhInU3z7t5M9SEqKf1odMHUsiuTKJ+AG2mN
WdC6EFrT0KbUgr7LFzG87q7PiZyz8Tdmswx7jklxvxGoYOjmJpXI3L3WQ1mFMzzk
y1MBaFd+CDHOlzs8M9c/WHN0TeKbRpZEO7/0EHOOSF6wv291YIigspR2FSVyuLXP
osLW9i7FTvElLwTfEkLOUuOv1exoNR6ex6RIJABTgmuaqPdmC51qw4cwrY6p1OyZ
+zWQCAP2+GVLKxPGfq/m5G7y8ZzcLtNylgIlnffiThZno3n2Kp5Nwz879iIjnEiz
opLEDvjkyBha5gP3Y9/hJLRyqylwBV7jNdr1w8PwMZY=
`protect END_PROTECTED
