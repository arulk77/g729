`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49sYXKfpi/2lhmvgOSBPGAW/aq4MelL7TjcF1WLEsjwT
1R4hO9xCJAPX3i3jq7rMA+cQOX0de/7lScDPDX2cVJtHvVdIji4zZNMk1wHigu3Q
sjeqz3IssQcVpSGh7mMgZ/RVPAwRzo+sHrWyT8ueZXOSkZyTO3Na1pYkh88l/oRF
vbdLufWvqxHlY1GX5pe7muObVwym7k++CowTrhQz7J74VlA4LM/svHb7caumXRB/
AjDbXwGRKtYqy1+cJPy92NkAX1KyQZrauGE5AkkPU3RpXNcD5K92IqIFD1Z9Hzim
5SHlctMo31GlUF0DzS7qGAApi9eTaNQ3vMxwQzwQzc01Xju2qjMx+AHbxwAyQwTR
+mhkcySbASHKuiZWWBwpbsH1SxQK+/mwUTk3TFVviIi+amcP4yg1YDe1HXbywasU
DGhK73NXOiMP2u+8D3UYpETDVnhuYFyNY/cMNEDI/K6rVSj+XaNHpotrVLMtAzsZ
`protect END_PROTECTED
