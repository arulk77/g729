`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJLad3NvpKGO3F4ET/30BChjEwm/5PmUn4KEntD1/6Uk
0P5yY2Zfwn5Sm+63YYoioEPOtb7woAmZXThJCV3PMpDDf/tinoo05WG84bh9DlOL
sru4PX4yamg8b7BaYcyIR43gw6jtSCgcXk/ckt1Nph/oUjq57EH3XW4c7YSIejxI
+jlNtboCfFjDHX53aGhWtQ==
`protect END_PROTECTED
