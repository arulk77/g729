`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGGJHvTIQma88I8h/MnZVe/sllux8PInWFifewH9RRvn
C3U20HG1RTej01xyOqRsaAcRKl+eRCRP2ry2V35RGtjXS03xARuwhxKRk4OkqTqs
+MHQs2WfutXtoed2zWEbJyfuxbzYfuexviDiog/l+Lg6qXH9jzwuF9vAqKklo7O/
ctWjGU6h/npCwtaazizt9+5VPea/8egp/lOE06XCg8Kr1zdn/Kzn64NPcxmrijh7
XHxcxIXvWLyFiExD021yEtFT7A1MGLct48glnm6hviPJuDvpipMik8OHCnsx8s6u
jnRrFfClaFP83BTsb+qIew7YSfnHhixZRoZLbKfrOYCaEUgs2qIeKE+rsxCsAzoW
XmwtLhapbW0l/uiBUBFpJw7TLo4ABLF7DyhLY6HJzuze6rKSHfG8Npy4xzeethHc
SHfoyeNUGaCOmvdl+wKR5mOWSyLXLqyr7Ta76ngI+nhwVl/M+CV1wqzvPBq1lQak
wUJYrKO9Dm4GQDvVhA9OIDEJjQL8RdxytB7NdLhad4pm0Ccgqn8aUvZuMOFzoQAi
UIg20sNjoC/XvEmK86/U0Ii6t1IYR9jsK5NnXcx6VO+fBWHJ7KIw2iWIDQqEtf0d
qM2tleaKZ0lXxU+JCwQJaRLvpCGCzivUgxvNsLnz8IRB1b2FMEJOo8j6dENd9eFf
Cbhrd3R/xt1qRGs/CLxAvv9pE10ms++rHhOz3lZfObNf9quNItgJweHvdtYwa7TD
Q1hW9CWG87yC1r+1o+1C59/sP57zpc5yu1qOnxjWU+oXkeS5qhSO0aTggCkcJnj2
t9tAhu9rIwdJ7IF1kS0fvWC/SY/u9hyojNxGbVax+b8=
`protect END_PROTECTED
