`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu488BmO2BWqF/Uqc8r/+rUabLRPrELEo1LIcPiD/yY3/f
+ot4Yt4uJCOmBM0299t4DvNt1cGHBSkFSTxjQV5FV1AoElHpRAzGW2N/J5c3tZr+
PY5thMBvrY95ctve4TF6/J38aM5wJX+mbQHLA3rGCB8HIAhsC0pC/T5+X9lZKgXy
cOhgYJM9TjU5tbJlH3c9brgfwviLGO27vM61Uf9rfNZ1e1uDSi6HSynixtS6de5r
xKitXrs7Ed0exnSLriIuSMIIePmondv5IJrXd/H30RrUMxGnZTNdtGqsA1MjGXPB
+0ispUT7r+5DEtkh16dd+3c4NkLVAN8dX0Eo2zzXulMnt8HSmmEIwIp1Eg6Ap63Z
yOMw7zq5xJhrfYsCnIR9fQ==
`protect END_PROTECTED
