`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBN0aC9H6J3KTNkYwzg9vhH2w009FoMIYYHgu6vrP+ZH
9swQHZp32hCGEdpSkW3VCP1tVl/dLs4r+0kruVDHLh9YppCHgmiNl/bmB6eLHYF2
vV7UNCV/KOjKtmyH/XkXxRexbiL98vcSHc6hHDwfDU2sm1crmXLHgeUaypyHVyCv
kdRMHSd6i/jyZ0x8ZOit/viZlQABZ9/rcBvNnDGULGZGzB7w1wL0N2odhBVnqc1X
XJWBp1yR5CLsOnU7iWdtBITeXLB+hPtZsCawsYQAFDnhX/ykvM9ONHSk/Rhfp8VC
ZQlcr4j+4yrr50vWWvAH8Js+7v2yhQXfdj7JmmAOLnPxuqEvFDQAFj8BVxgfxlCY
Y9o+0yhtIKErv4J1MJWHVsl9U0+ChCmLgm1CyBxb4HqBlaNQV4hXSY3VePcmSE9w
Fb11sdl4JQ51AWjlVCXxtxsf3YzbWPETydDj3UfopL8GOuvd4BhxNwhWweOD+omi
q4JNujS5eGSi7ZF1k7jSzyEFJJriry5Hp8VTfGteQ30YS1nZM5m//4KVlpgpYaeu
gE7/N5USVVJq+gOLHbujg2fk2CXhMzfWftlyYt5ZD9efQr1xLOpxLGzvqnkG1eoJ
`protect END_PROTECTED
