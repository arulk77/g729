`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBgYJUKbDIQLw51cqGhorRJ3gRvwqRDgSfndsCukiohD
dhLVof2dcWT9OUUBedDW0RzMvg0sJp6BL6ujTpZz0e2W3oT0nhne16ATM1MIEJDS
rWAan6wRnhjhBiZR6I+Bbu38t0hpylNtvD+Vqd/KKO0eAuqzQmUOTSzh9hpp0GvL
J4Cq8ErQ8RdgYugPNh6PETx6onWKjtYUOwj+UTWBy6yGQK652ovRMm7WZTtFc+//
sWbHdJgXbcApmRuVUWnN85aDz+tuvQGc/CRdjRRr1/WZk3+ORTT8TYtUGxjJxF4y
ZRMyPBR/RilAH7KcFyHCf7a5XdyLCz+wCzHaHvTpvhQw+2GgpLuUK7QXUBr5s5aC
ivo8358XvJeGIFZdgXwZIoVGm+CkopC2rdXSjHIHzdpMvrD4FuSr87hSdrrssZJ/
kv2FqrvDda+grzbYfMvyReoIp468uj29Kf84fGfgogVuk7P6F2dKdwe/OVmNX623
`protect END_PROTECTED
