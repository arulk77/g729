`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBw+qQJss6vL38W17w8+sRdugyrrI4xeX8tZqBrsl8mx
//JrnoL4LSzPQQpl3AbAC4GhbDnsvtb0e59NQiJzykNivBDbyRq+ypKs/aaDUDDy
pwhfabWSbFW62w3LpCdaDonSGSSLmucEsmpk8Emq16yrQ2kTWAKjyIFNkDQhpu2i
4G2iSuNy1QWRncEzEQ4/6uAwD1eA2oaedeLBEh6UhBqSAI4azPZI4lGZJlzvgT0Y
`protect END_PROTECTED
