`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4ytpQ2xhKWkjzqPtdnEr+42j1ouYruZw3Atpe1Pgm5DO
iuZ67JZEXBWNCMaUymU65nL10xH2bUBpgaUGrmB0Hnrgc92JH2xyBPApEodPuIXg
VwnkpBSsL2s50V1pdSiGrLaRtmLdeIvv33avwVlf/pQXAGY4eMhYuQctauk8nJSJ
I8WTp0cKxaM4XbAqD4oHdicmviNN9um9yQiuw9DoIAZAAnfhHOiyYNXH2nwWLmDY
bwieCO41Ae/tFp8MPOLUUdQBnmglySPP+BuR+7Pvdxo=
`protect END_PROTECTED
