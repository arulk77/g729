`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKBia+m6KmdEpUFooM9Ug4JRqfvaS0XAil7LIa1vQnzF
C7t5qEaxq6sqq0R2AmgADv/IJ8jXwhnnYKGQKDwPoxtda3H6ViFPLiw0/JLbO8Cs
bwXmVqTur7oQuTWtOk19e3IDOT0plbDsrSfxutMrnHa0zKHBTetHiAeldCQJTilj
nn3GuNxYrxJ8Kd1YmHO7qgHimcQl4uroYwfVmoV/jp9LviBEHVPzkjycUBd4ZbP3
l/puJym9gPClxOWx5Bnr2E8aXLoltGyQOb31O5kmolr1IOOhEZcczt8N+/2/uXky
AmOf8+CgJRvWoXyLtUTB7+ZK9jnvEMaBavTJa40bqR18cRPeqIJtdQgTUCctp19S
9qVci38JRuL2wU+lGPKXLtQlIayLMYW76dCObjAcwGLvlF2sN/YvBkXI2l4w+vmR
6vNbyrZWfIvZ4Rkgjx9u6JeujLDlZFswBLXGhoiBlUzKknP9EfHaHv8moPIS8HLB
c7SMbUUEe7IakApC9nCYv/rA22pkK8rQgW6IJVwXKwxzcm1mbj4r776Cx3qv4wew
`protect END_PROTECTED
