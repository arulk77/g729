`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePP+jGCutmeFHwCU+5ZiUsDxwKU2vd3KjUYGyaL9rTaZ
jao5m+RHBeJq77ga6u5ZBjlEEyCwFGQ8hUY7ZVMJ+ecxvfujev8wZla8jxmbBg6T
264a0lLMHZ7QlRbhZgKLanNxxx960vpp9yZ0BNeaYxg6GK5i9QnkV9+yJeicMjBs
FWT/qvdzGSmdnDIB0LTy/Q==
`protect END_PROTECTED
