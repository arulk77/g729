`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKSAOp+un8cZWxWH7Rg6HmfK2RB/98YhXGVQIfUTzPMX
xVqjyzaISms/X/vTH8eaAzhxzjEQT/26wt9RVlNQlGpH41s0slo4q15FRiNo8ISx
PoomZYvlyxLDU5c6auoxfy6zEw4UIEl5Ws9cowpknDPNHDSiD1ikzTtmyN2uiOD4
t74zwAFhBQe7B2tOc2dO7OnK9GPfJfj+cr+va9Deq3OOLqNoaFYTXGKawTznjE3h
p+sodx7OEmKE+yz7q/knTqAW9if7WVge/Z0Z/1ACPupagqvmjHs+oKZaEVURnCez
fBwynnW/mX2d5K1g3HxDwcxa6GgbBMG6zeYaD7FomNGTYu5fMJVRF3DBhK0ggQMF
PigM6QvFKoDetm8VzBWbCWi0f11kqptw8dvtBMb8xC6FTHp5lw4CfcfcfxP+YxLU
JBH0CxXqGYYD0qHlXZOwQZ1mqBtdGHvPpgRtEaEMNUe66qLq6z0F1wiNozeIs2Ed
HOzJ8Sa3kAz9bZaGOUYAh6VoonfS4AKA3fsYQ41oKM6UxlEaqfB6X89hamt21Edn
`protect END_PROTECTED
