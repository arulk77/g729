`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
BUfcPb/PGcm2AIDUHpeSqBfAcU20v+CPCXYR+prfAl3Ru/YnCRpY3Kc8Egp0titm
AycWsaQkKmTNzwh9yd7TCSN/nJR3yhIQmKsOeKOR7iQrAPOUmvYkDS7SW1O3A31E
APpIdQfO7J2VOqoBfpO8gJyz4FblFeuUQi9fQg/Gvxk=
`protect END_PROTECTED
