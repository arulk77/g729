`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
1IkYiFYXomgUyjOGxpNKfboE889iGqp7963nfGi3906m4h21CXSIeQpB5I6x+wc4
K9kaLwi2jMsjsc9/m6nNnFI7+5pDq4FMj1hKRLY9ItM3Ox/N0hxts2F/xk9pHsJb
LkV1QGr0XmfmIdTj+wwS3DzZZqmR42MDdM7PxXOjzqyOA4mzCT+a43LEiIIHZK1S
nHE0DMiWwND3agV2vfAsYgMyjlKrfncHsWjNt3qE3/lwPQ5dMZCVIr06GRrs0n4A
jVNHdcMGBRQAHt9aA3eQxiFnD8qB7r3NPBTDPcT5YKQ1pnI428jLZxzznNcmREQa
6zybowmV3Ohso2Ai6A5450E8JqnfT+nssNeUMZsmjvO8d28CQmsoT/6hF4TPVtM1
nC/NLPR6sW7JbuSQVIMRAZH6AuusANdwMSIeq7ETYc0rSi3KzyQpc+R3F7noVV6U
B/Z2BXOMSzpjOyadx4EgpPwyVb2jL++HqB1Y5QLVnJHLeCRpV3o1B4cl9ZzloK9E
D/Lb86tbfq9ytRcDvHKiMcsPabIKuk7aq8mhSrFmETo=
`protect END_PROTECTED
