`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47ajirht28GyOLDTCjz4DAzpS42KkvmdQTHpp9GV2d/H
cA6IpX7RJxaP2HgIaK3hxbeYGa4QD73088XVqtuLeCKp1NJY2Q8p3XgCEsbRyf9t
Ip0c1yiGda6hfJ/Oi3mCUdnVROuidmS1zhelWPT6NwKd7V5sadeJDbOJ2A0ToUms
QQirnGuGM2Up3SGbSeZEyocT6jr6JHxtcoEZM09fPfBfz09ZTsVHbX+ib8d7/tW3
+5E2+cCrvq434UXr+LMgAq28Cw0w7PKELb9oubYL0jxK/mJcQRTmx7irrhBmYCQL
XGP1VA5b4bWcOReIpRlG2EmhcOv6I9dkMKtydis5uvykNmJL5Ejn9MHE3uYVLJjP
+m3IYH9bZNlfc1r6mcx1TKiJIoVSYH0piyjAy9IJtQaPdhkg0xnyminwh6paydW1
mIsnfN9zqqhVUinlVJ+0wA==
`protect END_PROTECTED
