`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ8SCwcicr8NJ/6z14CFig7YevsXyXU8g2ySDtT1C8lE
Jpl3fz+vtX29RazrD60B+mnXQQ/hNL3rt/kc1Tg28e1bJJ24e51q8vSEiuttU0w5
MMQxbPgDMUpyycS5w+V0rCq4L2qhYtnMfy191Ysooju6WDXxK/tfTU8QCNgnjJjg
F74r/l6OgXNEsSmEXCMr1BDoH+EAjcnJGx2RPHmZRjczASiNs7uQKZYjMO7j2U3W
G1oddeAqsluqszpr2PK+8t/nde7Arf1edm6mRFAM+JW0fruqUcdn+7/TDzc6dhvV
vl31iMoG9ABfLV8aoNMTawN7AIU9/oodFl/F/Y5QsG5TBR9cmO3ZTiRt+krY/9la
JMjmMg3oX9AuOX/cRzHQ83yzV8tMC0Fj2zyoR1CJ2EUYO0BjNMQBgOcKCVfTD1m8
KxNP7BricUIIo0FrLuj1+3EVNlYmYmXAol4X+n8LfcGyIc8uTU6Gd9zUg7RSyGAq
WnccBBPCKpDupWBbTlVQLT+3R9PAvsVjttniJLna8wKOZIcuxy1HRa1WJIRTOsqR
H5Y0Cd4q8iZxV/K3Y/GtDO5CHZ4LH+7HsNogRTnzp6AvX7bzeU01dStuTiQ9/77m
lzem866eHWPLSL7ZQcY/WiG8PZNXSiXR+tsULWb7K/vHBDwqMH2W2Y5YhCrHDUBr
ZvUuXhRzflfLs0zcCnIvGvoBt9ExdHzm2f9y6KgDXJl5Qz17mscgyhqofAJN7uO9
J9y9Q6Guh+Yzey7q16To3Q==
`protect END_PROTECTED
