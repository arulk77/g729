`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEMEjRNDC+OvVfZ+NHjj8ER0MihjOBwC7VLBku2caM8Y
+Kj4EJd80A3Ky13bRSVjsaukdkKT2dxNV6s25Wa4LQcnetvhNv8biaWgo9MACxLR
s11UC04NQrMobZoMC/PYXiQ3SA/UBoB6ZJ7Hv65cO/ptHMiyrgIAR8QCTdpnDs16
uxRk+nlVkChbjMr03z3NMQR/dUD18WWmOOQbHf7JFjLeMkQAzYQeWNHT06IB7AEr
cDaT9x6NyzwzLcygOGHXepaE2l6Q7F/tB4z0EBwUFJGW9/ynIFCu1gjxtR6kogfH
XIuQiz6CX1oy7S283mQnCUJOW3YPBexCONMll1cpEBtck+Kpvi8LXWCK34PFFYad
KEo3WD9oRJEhQ574TRBcQ65MmkX5WcEB/wr0DHdbETnjNPlVhsd6k3JeNDH9d/j0
ra7hz4EbXk7UkgUHbP5rHPtODPvXCqz+xB4rxlGrA8Di7WWugayurQiCajCoXF0c
WNWi0f7RzECGbAdWMP/tAA==
`protect END_PROTECTED
