`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGq4UHV9Z6VozVj4IIkv1Rj2kqf2JZ+tHAP7JV0kZraq
6GH7ZWALljI+LNNEwkU+yucK3H1WGc11L4RWBjvXoe5ofVq+lm4zUMeO9v4oe4uL
a2uumd1EvhmO/0aqLy2v9Bt8CqEYSz4I4+IAenLnqZ/uW+0ArCAKdDPh+qKOSNnQ
YajJm8w7T+1WCyl+wXHoianVLbIEmtFHc5dS405OEwuRu4NVEqMT3MISCj3Gwq7K
YEhzh88m3mMN3c/HJFxoCeZvUV9yKL6wrPn/4RoST4WR7mUwJRssIqiW0NFXVpju
rtQe2As3RncPxx550dnKcgdqRe49mvL+lht0PItsfX+388pEYch3rEOaK9qW6wOS
GnfbOvG/HeJYM9d5b5OJGFeIABMe/KpH87vJ219UaUR/jzB4Z2crT57ScCmfypTN
XnlPBwQHVe7dwhn/6/4OrC4lynzGX9hl8xxK+/uJf3COWq2RBfYjHqbKKJYqigrH
h7jeb+OT7xvhapTALeScYHJfbevkSxORcf5210y7cNClf2VAd/N5FR8AbSMzmkIi
3+oR2DZd4TfYbU3Ql8vsDrvbTy+87DdqxKKigEIYyZLGENGcljoAGAplN511Zdsl
99IEYnGHW0QzckJPri/AyNUY4Px13iGWMVvRHrGo0EL1oaa9evZLaac4sXu+HAvd
`protect END_PROTECTED
