`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zAmESeYIHtLsXhDbLpxBWMWvVP9NmUDN2NJuYMGW3ze
4vIzsMUopnDaBQt+hopNlzxtFBw/yopR4U+D1gtqoy6YEQWqxJ6xuzulo6K5s93l
WZg7JxS/WtwsC5/qsnEyOdfiGt1jel2cgZ5c3doauct8Og98OhgN/ys1aobk0+KS
CFhyfFR4AvdnoBkP+3V99313oHDi5UYb72dxtEzHzdvge/plWVW/jtcT48Cex58T
7ksRnPCizvdCU0zzI4/5CIWkPrMsc1r1Xj6rVH6ULS4=
`protect END_PROTECTED
