`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD3SP53oFaY3i3BDxYQN33IbOGOQryV5Kk9pKne7M73a
1V/17adglx3dxGJbzVPTAq9Hhob1e+cszDV5/6gksSjdqF9c8OihIoezeOJoMy9O
Tm1qBS1LE6TkITeJF8EuAxor5TFiP2CshSwyp/IgQSm7Hi+nacrMTJviZZeCFklN
77foWMrlI0Zjkyf28VB9ekxl50mgz/GGkeMmqpLhOem62zcAITo4LfCu7tAY1mU+
Pc4fTlQ4NQ6y2TheXnOfldjOat/SWdoIVAUG1zKWSU4sbc/bZX4UUWCgXdJHuS+R
tfHuRmXQTMlNuW6Rrjoo1l8XvdazGSrxxOCUiPkiaJo=
`protect END_PROTECTED
