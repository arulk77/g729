`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
rA2hBHSL51/AUtT6Im2oCgFoKjuMhVVdeWVesrtlLp9r3Z3UyOph2we3IEvQDPEd
Lb2tyGyBOFshLii+ERYkyLbnHgQzBUHAUHJSvVACUhT1kEqEL/5Ig5eJtzhIlfIf
RavBidZfNKzqwH8atx7ox70pxg2CtLaSW0x7W3t/rPM/5OTlIfG9yYHjzgjD+DxA
z4uQQ5GpQNBKcktiZ9Y4n9Hhcg4P+SdEYPinvJaqGRajREUoouerI22x+qHH7LwD
T2Rf8VEBrGnjmYb2X7RT16tjOM2ZLFSuWHgAF+Og47YtFewPOwvpEcloyycIWUmA
8JIO86lkfHfRw+cRh5DWdXFfLxwVQZIgmtG/pjRXbCk=
`protect END_PROTECTED
