`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mlFBzCyNIVABC0bhYTMiK43i5l2rUjwZlqbACUft7ti1wHRnN6qvUwtsfVgq9Rah
VWWhQL6kaTCLtBwFnjNPQys7fx/TUUk0ErqciJ4/HiHUslD4K7+eLHVhwl3luUZh
ljCV19jirPfzv8f4kQXvToM3Vd1RfyKTdvz29PX++bNjwRxLUuqE3OUA1B77qozd
ykFcGemdOhO8YDmwV0p10BvSDoiELB4FXcAu+/Z4ZX4RdRuB9e+YYIdZJXxV78pj
C4K+qACr+OzW4jH75eP7viOY+zkZlPvguLZ6q63MBeXKM7cL1MX64rKaVDASWemb
FCJaLxf//sKx0RrucHCqTWBb9rek9mWLbaTXCieTEp0GaPuTupcr0+GpxfkQ3lc8
JBv2C8HA/qupnDrEBWACWFPOceA1kWOR8Pd0LaWXWspFjEx/6CBp4Gty25dEVoL9
mjYkHIIXq3LByROm6HsQdwzKKQ6tN0Hq2NNtAyxZTLN9l7QEATRBb02wuf37Cp+j
CRAeGrueuma/yynXMl9IJddhkOVS3zEj5DoejIJ9qjXeua2qrudDxDfBW+VrExZp
+6FufIjnfF1o7bYQI8k9Xa5R0khyxG+hArDZ8wB0qejszmDbQPc7U073VoMCO8Ow
sH8iev0TkkpfvoP5PNkDurHC8R2gMHvvWF9avSC1un7n6vrkyIEWm1/tvJ7f46Tu
UWewrIvqV7y4CR0C6UZ5ebgLAO4JJsbv40hoWGCCYcxfZPIbV/kj3SraoVNVAZOk
ecPAc/C/vKJ44ioDxL7VLe/TSbGCDewrq/71taDOwi3ElPRuzcSjPgzQgzN+YDya
QIHsN3vuyo1XmhlPsUdh7l9ZVxVUhfhZl6tCgmUHxvACUbnFR31oubYozuuuUen8
uwjDNMZODAnYpRvYZMzQGiVvPzizAUjb5zzM/g/DLrFG9R5aF+QXff3kopkQ0DII
rUvEy4HFx7oPI/4/JD4ayc/16P40BhMl2zlXYFo2NIQIby6xHWNzNmQQQTnXOy8O
fWiszbYOvWtzGAaHOdhX6DgXtYUhpUmfY7wByRt1aRR/dcdOw90QNRv+2gfFlHez
uAMekEayI09FnobA+rtZTJ4C1uce+cUIP6Exj8aTbUKnCiwBCkJzuTPSYHL3YCaI
w6/KjBr0ksYjrvaspItWpkzpQRX16RCelmtqSAgkzfxgE5/NYEi6NRUoQOBiWgMH
CH3jzK9RX2okHqN6ZGMA6r7+R72cKgrbrUBJLfO56nKBosg6i2Vdbg7JVhtHHQmO
+6HZfKBpTONkGc3gmYSN4cuSaoOrQYFUPohrYNvB2z062LO4zzuhPK59pFHD8kMn
F3aJx8X5Y0DufRB5I/KJGaSpRF66LeTaFwdxNz5BayskCHmxlPL+JISerditpRcP
w46wD6UyQAErF8GoqDJ/T5iamDKxw8nKVa/dOuPB/zaJ/GCNkFco6FCCvciXvx1Y
zw14xsCaM81UBU7IVDtIxBGoWE2FyWYplDkZ35847jEV4PLyOzvEGvhSYH8hfCHv
1h52P0V0Sz7zmda1lCAKpmNEJ8auGsCvW+hhYVdMres=
`protect END_PROTECTED
