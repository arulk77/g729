`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAYU8yF/LAEc2eFIOc6uqhKqluWj5Ls3THQ/w8dr/XpKO
gEcgGA9rC9+svM8PIr5x/rgUEpZswW5anzz10SUK7ID13HDImNp8oYc1aYOWEq+I
dy1qmMPkfMwNGRzauKtcFLd7kUfcYOhtmGkc0VwYqKoS7egFZicajEUSz1EpV5ir
tcrIn0nbuJk2HLBalTvVSj3vBAl95wb/+E/TwHpdzKZJoiQBpQNTfzzyDw3sWWv0
5hyXimYqOgQO1nJJhcOy5MpW0Wx6O4a8Q7tGEwb8J5cOYzVFC0JDnAWKUW6j2+/T
L1dmcpsUupATaCIjJueYLU4fZFV778J6LjjpO/1yqsaK3S/wJDGqY2enaH715uNV
LQ+XuHrk6l1sMokr+nv+pKyLfYKzx/50d3Qspv/5EkuqzAnc1NaXAFtFOO6lHKas
D5GZDGZ/K/7C5MsjQYV+8Xje7yOFezpDSWlZ9fzmBiLOTXFPQdeN/RppZck0q9bi
LnC0g+Tc7VMTsDeyFKuBvh+Fng3np7u5/2hGchJ7PZhYChrlMCN3gIKGe3xbOX/v
7qYxdcahtICtPfW3zZZOc9KoOO4FmaNHfmmMye7dD3iG/1B6FvxMrESKgciF/P8H
6aY/ROFnjF7nyzJQR2eKqO1jHoZ2+fy6C6QPhQWJIA/nBqB6X2zPh2Lc75lRehli
3TzDdATSsvvDciijLYTHf+sfyGQhicLSN/P35VHUnuwN7KVJOBA9MK+Jdt6CjBBC
SY9IaD97b0Fnl2pZqCxGPLK3/Je1ZUqWrGYR1npejSwKbB4mmyqdxVWecop/cUNA
SSX9enheV0o6ItE9MN5/0+vctoSl+xjmyq6mvc0dLqcMWQZEO9fwYaLuesfZ+lEQ
kCSNuDeSJefMCET/7q9crTn3DXhlujiYchnxOYmtGGAMEnDCRVq7Gzcfm+VDJqNF
rquaNDeTticxqGYIHnLKZcS6YBCPoePMrAM7S9C9+F/HHb/jJTfKWUundR5n1xEb
guJvdwFi9XgfuE0kxq0JnVx14WvrZ9SgsUTwhRO701BNjNbcm38MwQRGlUtAQh/J
O+1lO8Lb4GYZ9Q2gVJEY+MxSAnDvAzMt3TSfLV+qAeZ9RBd3OmIfwNeZqRwlPHrk
b8Zh/C9rrxKrPuuU/NmVzIg7W+FVADZQBQiVcTYR02x68m+Wi/j8SpcsU3/duH3W
PZn4ZuFaiZrasIjA0tu8sluCUpiXL444Bkh2kEqGRWtwK8WewKjXzb5qel2oCRcl
s0KspZG571MQp9CiTwklQvvyWoX0hiTcaKpU9O9vCZBUVSm3qLlMPcWlA4kVW4Dm
LylIO2dOojPt9Yddi43e5esAphiKSvQ7SdJoIqwlsRyYFlWCfiOE8BtYk6Ag9IyS
RuqsMhVTbbiVP56tFhibN1qCbYs9PxkCofc3FsPWvl6vusclruR57HW8l3qb3vir
pXIrPdfLPFaO8q1v75D0JbAzZj3nYoxkw8jxOG2GdXBOVmgwh3ULALmL7FObRcBB
iWAulSFeis8l63GwtlRmzxx56IlrWbYjoYp8jjPmqnvuyIugZW7mShNKvwaoVqMq
bjMZbGqtCe9rBafGcZmrIA/mriotJFeCBNNzWRy84n7sQJASXYIN8z/PBvPTaatk
v0UxI/DRaWfSplBQzBQB0XumNHnf34SoJKxM2V6mbHBOy4wxtGGVVNheAh2DqrOu
k9nQAFPpcf39amca2Vyxag43GRx3t/khPt7bYW08/W9TcoVsQTBt8gLjB9YkBUSm
9rRS0ucmYoLDAeZ+SDtHBKzZpOBltyFTIJJ8WqvOWPUsWsXLnvHt3brI2x6m1f9+
zyp8NVdFjG4EvVmxcS+isZ2qyq6LB82Giw1Juv0BYpaLbyVCLqFwf5PRxhMmaTmE
ByIycflW3Yi1sRRPA47xN5atdWV3999C8TCA6r6LhiLPYk/+ofmMJc5uv/n3hn0i
cdPx1g/3bHVv0RxtJ8uau7W0MjGdiGiE22T6orkrzIjBQpDyArFycIIKUSkT5Ez3
Ih4eCyeYu/JChYGJo3UESAhGWC0heQam4bL/XpdSCyqq3rRG8RgrJCz+4BRLI8SD
cX1V08nRzlo2vTiZuhzUeNZ4ZyRyqEn3ae/x5d9B45PgTduTKEw96mPHXUQ7Eci+
1KrCS+ucN5oAMfKBvV5zQ07gAnqUc4OlMzh7c4vu5IM9lzHkXI2O7v4dWX9eq4tZ
7R2RqqdXcVnaUN191xJVPf29neDASs5hdNFkHppR1Eh7ZWVrRDcnUdYJzzWuzWWX
vrcHXWKN2a4qhHiPkd7fD4I8P+XwQAiYoW4NouWZmNEXBq/T7uiWjR7sSmvtLGGV
ETQtlAoQzm4cWWwdlenYZMNtTp2kfZUaWxyIruqzb78/7igu2kmLuQ8vRX2iAa80
FLCunvKwLLTca16nN3UeeLnXTwIPd1XWEBv6wMBWBVbHK2B2Z8iFAswxxcrARiPO
to5WCZzJiL94Ode9Uyv5u/hO9Cz70CwE3K1RG7UTuv5mu7q5oOSvHmmg5GJoz6sf
AaUJ6BC5NBeUCdMJdL/3oCo9iB8tA+Rw8fJYtDFCpa3hH5WNgN5c6lBWInywCire
bGSUNblfRkjGPz5CIkhVwncZRS1OIW3BDhsCO3+6d/5Xk/GyMqd26CyK9fnxumxX
GtkcMmfeicTe32x6kHu8fNo1B3MvlEXPp4miGYHlqC+evTx1FZoLNwPJ8LcH7B5a
bi/AIJlhaj10FJzj39RvFcONVyKPrI2nP+fXfUpM594lHqqI92tYsfMV6O2TbSf2
dCwmWO4ojzSuLtaToMC3yqjWht4a6AxkWJJ6q18AVRfJRRfGHelonLRuGvEVSXjI
7MnkKqwBRL5wwGI0anC4v6Bsyc8CFNV0aHhoD7pCpKUl9qsUuEKMH5gvM3XMhx8Q
uFFoK1hxU/FxcmTtSBJ7fagd5vjCNKkIEbo0twEZ40O0fF15+O1i0X9CyQIxr2q1
PLUR6NyCzsbsWFGvx7HBLJGZEqROhEWu75ad8/H2X2wYUF231+LKjCxRxjuaevgS
owrqnc4qTgW+rUzcFuGwXj1PWu7gnwEVwXmrqvvx0X4218m5BR0CYqCMiPKvitqB
xXI7mmOM3E8sHCbMWUHlqM0Lc4QETixnHQ73PH5tZB9Lrt3AmvGVNrI5KoHJgUpd
6zMSLWsRaq+JcBQ6CvY+oq5T7qOFyYB7om7xIH3d/Bdz+25gSv/2atWU/8q/Cjtc
3I6DdXECS6DB/5KTG0+DxV6fBLf+VmXFJEzBIDsShmLpx66tX0SjpZMUVLZDol0p
wozRO9GdDG/8mrE4knFg69nLePejPLF0MOOTETT/k7a+hUGimC8iIyRxAsSTyxO7
8LRRrNuFTXyAdIbPnVt/rIWEq3G6DL5W+BQ5YkE6p8CRqIejmuq/EbMwGUBApFLp
xdD54ipYB1w0XQzwQDUVHafIE8iqfjHyE0gl8G5KSjih6xyhCC0fRaLt94XMwWdu
N9OhHtV69o8OONNJTymKAWBXqdJXjjaxW2g6aNAlvcKCloIR5M7sKtw3SRHT63xi
wfOYOUOoxKqBSGTrlILVtT3jiiHWAiyDsCRN+aw42n+kuS31NyY8jgpiT3MSSN14
xqVBkW3rA7uuij/NzUURLoK9A4ZMZ6RjfPlVZt+Ba/zUq61r/NtVka4oBpd/dKFO
fC7VJlFcIKzR/oylrn8Entww6X1ww5ge6MqL1OfRRAKLi8fUC7XsexU1VT1bKAM0
nDaFEGUOGXgk8+pn9RhD8vIwfGPMblyXY+0JKB5yfQioqVffL4pnDnVq96YJAUs/
xcMBrhCmIleRqW7+NNeqRBtCllWXzvpMgHLlQe9Fzbg8uue7nPLIj+2Mgqz3Qc8S
+wQMc3QbewQfUVWazKwS4OFW1Gc9DNgBba+jgCwG1ZYQGe1eQvYs/UF2B4gssi/M
DL7pfmwAMTZ2WEHp1lSJVOEVV8hvuy/Omrdw8teGE1NmZ0fT4vRGEUuiZ3ENdtq3
7K2mckYf8u7b/vBeRdOaVX+ayHTpGu8cd2yagvg+KD83PsX6TKqMLFfT66uwN/Hf
1C+nVpXCF18I8bV78ZuHXnKkHoBPjCwpnDivxA3ep6f28SFmCOmWiLu+1TpoyQTl
T+Zm/cQFrDo92/kOx2CVvnm3hw+MZR/EQO8PZHNFSazY6h/CL9liwEDKu/cYR3KA
AHkXBjG974lrZlRZXxLb49fcIIAayI3tQzsBNYJPaX9xspb76EwqQG9vPKU3btxa
aeNEgC1Kl6AVj645pUTc/6wtNrf0ywyOrztUw+mvSOJrZxD3ymUdU24QyuIb0Yvq
eI3ODfDsKCfGEDzKEuIVNEh5kaA0uMO9UbotVUhUOEKMEbd5X8qzWHenku0jPuw3
6jurLVNiPz6z/SjMaz/PHJUU+qKVT33QXKodFCSz4gAUbfpfqpdvG4vimXba8W3G
oZqrBlHPOgyaTUn8Ocx3Po4+4znlE329xZpJPM1mSwsFk1QaeNtF6NakbaF+tMe2
I7UI5zICV5LQ+Dz1dNW/0b1G/fFP7tKNPs1MZ+MJLq5JYQEaiSW8Len7p1wuBV+A
GGTTMDzVMvAmcdW1D3sgiFh499nwJulS3RpH/xC+zgMJH71dhslfCSSsdnBR8CFk
wArhbcrnxL7v2JsamEQB5pdY9Iq4CLEVwpe2ZE7yGYc994P3HtsStXlWZ1zkYcPA
O+Ehm6+WaEyGtTjbXzdI8e1I9MyctWvxcMELvaHwtiOS/5WWMwv+dNi73PuCuJAn
3YCjmw/MlmesqztcJQOcKfOmaZz7e8Z2ld737F/Uz9KDgUjp956tCgRrlnQzbElk
Q+ntmiFRz2m4PrNBIhiXhNvgJv04pTaGCLknb74/hFnN8UowdOA8a0mieH01xVW+
acgF7vzlfjLds2NMH0r3bzh1umVGmNV/n3aSxw6cWflqiV84zJsmXoUdvEfAuQrt
X/vRyTtKnLyk72sLIfc76kfU+0E4Sj0TlFzf0Grst8wJhztNassifWaJ2tuHP+mj
NodqAQzT//utd5gGLh/Cv0SPZgJurgLgmhwFG9jOgnLEkNV2W97qnHbsnCwPa0iW
HhCgrctgay3evnu6NgvY4liw+l/jgr6xlSqh2UzvejxLxbJB29IJzAXvy2rV/oT8
HmnImEGxlcZGyA/azxa+b4r2zD3cZFw/f5RZndD6G+HkvU2oxLPZb084xd+TdAJE
RRUL1k5QvKdxvwp8vygjwG86m9bS7uld9n95XwbyoTlt6MqcMTl0pA2oJQOPqPBC
kTCJFYRGBbxLPWhT72+6Fegs8sTslu5QoJ0h+rKsyqK3RDL3qfYXYQxrUjPTshCv
euGJU9wM9y01uVA4KZxYYED7cQtzkWtu5ZwsiFh/arb5BRf/BCcgJBg9Ph4lGCuU
Ph5JZuORhGPV+hr9TlJ7Z/OLRflxbcJcf175O885hetR5mcRfeBDiPXYhvj0hn/M
dmy1rp1gaslPTV4dlHO8viQsUao4o53VefFeVI3X8/0LSg06YoSXJIu9mGpv8uSt
L50wSCtqQNq6vdLFMg3S9sOo/EJV6GBiMhD2Dy8UuSYC11I8g0vdWOYGno/Ye8ll
LRgc4NPjH+01Ds55bvo44h5iGUz1oqyZ7vfwU+1nzWWARKtG2RF0WQbxIq0H16W3
+ZT6dhlyOaFh9NseoVf1n2CD8tWdnCsTPDmCMPuh3FnojrlakuoSIY6CEXcoQjLW
3kRldbHSq8fXXJHpYL1nmn/fFjKH+/acQFDLzXHjMl6jhbnRu9VqnjmJzdemTl/I
zwdKWsOCMD6NwvZAhYNrERZtWKyqoW3Zz1xpYXE7ENIxQK5lwu0y7N4ZVVszCs6G
VRsrrdkieeprnfIEtUdwTs5F76jWz0yR88aYnjMhQvcUSfig0hrPfVJka57zRl+U
jZNqXwcLmeQpBBN7XWZ3cv679ayCvzwqgvqg9LSbfQQNkxaEHMr8eDHsLVL6e5WV
j0pkJwHXLff6FHsIi/fTBeIyQhd4n+7fHSkbsRiM9Is4eGxQ7+66eviSbMLB1gJj
A3GvMNVBzio6IpyE6P3e8A3IU74GCTLJuVpGIE1IQPpJGqliQNEeHuVawInlBCRd
SXYz0pjFYShkcz/NokprTavs2nsR7ApNiulse4v5oYAke59BgsQjmVWrTUDI9Wdx
86gOjUnXKEDtC823tCqTLnKwxv6z2QnBC6iImxv2zRzMUmDo36wzXMcwSvIvuGWH
W5YleyP1eq2PZmfLx1CsWk0TqbgP6/U3H5GFbyslB6+915ACtSBs93a0NnTycoJk
i9oSnGjn0inC8AtK9bZ0f2+NvZUkwQAx5sMRTXIxZz0kLbh8As7CwEbKZKjPCBGU
ZVw3n7d7VpMZVhrU16ICZy82EI0wE5Hj9QSwPLV/52bnH9uksTqdsl+fn3hK8VPf
/NmnLHGdDp85nDuvsrOUTixVSHmFdJ48dFYuJJJmdBjItonWnLPUqiBso9PPR3vm
k3l5/jeWElCJNh0pUVl/NXNNlQjpAqMFGj7UhZAY3Y+xz/S5BH+677WMVRkJWUA0
M2CTs+fU6+LA7z1DsFzrvRqSIJCV6PckEwMRDZqahxV3mlJ6a1ai+eA3EZGpCqaB
1ZV8YHBoic60kV3FFVMe3QhGddNIpEv5NplAlTBWbZ698xBR0WDfwCytIaIFIKn9
TkJ0XRgmtl+H5udP7AaaQYKQpw4g9BhNNpPkuYege+aOl3x8lOLtHeY7Vgraw5CL
psYax/e60ygt9ElrJQNIiPE/RegejRodtNvdldLg3vkSvZjBh8/OKbh34Z0w48Wc
Dig1CbQGFZKAIRY4B56L9tmd3it8Z0e1OJSy8vu3K069XpFbloS1yJrfFxj9F/2Y
QxAuQh3iQ2DmngHiw0cUt8SzH16JibyDV79WOX6HIFSJL4LWp/ivmksBbwbeClIH
JyMaZt9i5/yyeiW5upd5NyCkqV+z7rqAVi++k+Xqv9jYvCrYfKYbnJdO8afU4VQl
6HIV6/yDgZH0UID0onyynKfW1tkx65t9j+XIAcFxM0+DUn9H226T41XvUBY9AJg7
n9RbbRfgD0pNfWKfn08Grd7cbruqM4aSx65HmJ0zjlBIwXE1i12KttZHu8g8hyoT
6wqoKAc1qPYiLZn6pYp2CPzWztozlB3A98/wuMbvW7E4AUdTkJup6OZPN3iUn+Um
q/d0dw2QoJCRSau634HghCa52kdyYzMhwFMyjkxCLcKCumfFVyZcjTf38hzhH0LH
eOZQZParKPObiIyvACoTHw6u+g2uJ9wpuayf1iIo7GE2PANSMGM2+DezCBNrTtF2
P1z1dl3RorZSrJM8r+ZQFu0I45AayxgwkeNhtlRge0uZ4T+rv0XvDCA0auKIqqNN
ujLF/55g27N4X2ohKto1haKSvCoQBR4vRq4JoZJOI/uZBFQ9Tf6ArGXq/8nxlZJ0
4df0VdefXzJQ5LFfH5h7Nl4kx3K3C+Qvv2Oamzn+X/1tIeIC4zJ79A3p1yRUFFNk
RdNhi83Orqqy+28H2EQ1BDlgiwc7NvRr+JxiO2yi4Xamm8eTv+dZT+8sI3KkJ4X4
14qbdGyM42W1QJJcwoY0PQ/AjqEmbYL+lDRcKMpLYo1lNduIylJvG5xf0e6H/Ob/
xM9YktEU8aZJfecMCekft1Y1kHPgYYJuiDU5lZvT1Qouv7HqESqEtL10Ueh3ucqu
KWA31MZmuwNJHToKdVA/TutbgG/WzTQT8Ywc8XmTg/EcLAHwOS1FeCtVxRa5rtqQ
dTw8BTBuZ7UopJv+4JIfsc7VWxUpVpn41xFIjfF1vb9EXbx+EBpcTRx5LKByhEcZ
KIlWZsAsewVOy607yC2P5FxWLRF4ScrO75REoHgYZgnRzGje0jVDLDXUhY1rd112
RHAo/6owPsop+9IE561+J4CrUngXon36asixJ+i6n6ijJF9TqSmlKPTNBs3yjVrD
kdoZLoQKxyVZq9oiyEKtOLUfilxvzWIUac903eaWsKnl4o68s5bvBuw/W8qFk2bG
jtEB5WwnQq8PDd7aLfk+07WuSsltggIgX61lZHMNzYhWzdbe/IOTGd8hgxO6jKnp
Knd+EqnDj6MoQXgbE860xkDtId4ji5P02BcA7WKJ9ADF8Cq7ZalMwCFXoEyh2CHR
oAOBSfpJwZPn8DfUHh5mpauqHrDmq8CZBjRdZ0wpoHRAfcJocJcDwbcy8fMmA3F6
vslRxc6vSOFiY5yLNg8BC8epU1BgVx3YO9xTAdUJGmQJfkPxSAsqfjq5su/+vg8T
TzIDmxx0tm0CZIz7BfSO2k5VoUM2AFiTuNaFm/d7EBAV0qMl4cnRNIcRZrXZE65y
FQo7K4SFqb7jy0nrvVdXzDqCGSzvjEI0N0TAaq+G6ossOrnBz/0uH3PLtQgNO77S
WuU6kbbmYzFb1jRY/te6nMha0zihcP4OevLtkbXY8AIQwmSoPyL3LYcQparOiQrN
cdPIdB3hRybqKO6N3yIkyp+CNRLdcLaofxPJOkreaaOsQfi/XO6AmWjoxGieM0uG
4pMIkJfPUW0L29CmXX3XIVE4hBQ8nOWy5aBQ3y++7EL3nGPSeCvyWs9Lkj3Uq9rS
IAI2lBBDngIi+M2YHqQ6SMls2mOiRl7HTv0eblyYN0UDCeVKFtjnxbReA75N7nY+
6jQZ6eETIYzzWgG+jbRoGCajm9APTeFf58DuyeAPmYLOjz/2yQWYA6Wcdg5Ssm5u
dtHkucUrdOWA6bRB+FXBbtIwu1Qw7KplaC0D86OXuSdWCszaGKx1Iiu70o484Gzn
0be64jE7hJ2JBIFJUN1N3tGcOcXKJTpJBZ31CXVPeFIpqSXGJ/V0Al8DAlJnbqxz
g+8kU+uTIKdI0/FzftjVTov+dIqdzhy3FD2KppRuXTzMdj2JZnSadReGGSRQkgfz
/i1K5e78SxR8VGjdQzMAkguIhOsM36aETzlymzLeVPjSJ4Oc5s8uue3vMCLt+8Lj
3nSefkbOg0HbgAbyhAHgVXcwoFYJjRMEjBP+Tr6KBRLBuIaJXV2s2Yz90gv3Cvmp
07CFwWhzHJW4hwHs2GF0kkvCdPe42pKhAegVqGh7ckgBrn+Efab+nXjoKZpQZMKK
jWSKuoT+yn/C808xuJ8U7DEViLsi4Z0RbQd21Ih6M74lzmvTJRBQHAcoGm6+ohIx
hKJmnFLY8x5BIigiK9NdsRcmvWNRijq50R039iZGWBx+6mOTKm5EwqFIZqS5K2mQ
+5YRxtpROEmJkFxhNk8Q2aDJPa8RbNXjpYz5E3zgQI4L+PacJ9TafA+3H2s83697
VgAkioQ59le6djIxIZLwVW82wvcNfKQWS7K9CsjqCCb1w2l8O0eHefOzGMsZhDdG
d4ZBY0zRaDT9N2HAF5bwhX9KpxoAgd9th8RegYZRw2fzcsqzD3x8g9uSLB1EHK96
Qz0PGz664FR20Rjydp+idIhYH6b9oHfZxO6p+x/0VRNM689SZy8TX2BTw6zY1Uov
E1mE+NmGZ1b0IYXg6aOz3hS9YGL3nWVeEXSJIT0D+2Yw1vkdM9DXWrdC4aj2NY9B
V1ykg6Nu2bhxo8IA00VV1YErEwvtppkX5l80+3i8cjG0Moq1vjVpGxDqpmXEtFTJ
XnRvxYLzVFLSXCc/gAeUNXsk9lVz75TvrogF0agDD6vniB6cbqzO0G1GvOF0+IrE
gQPvGFhytvvAC2QWMoA3LecFG9lNh28LkY0GPIS1g9F76e7i9fnJZGMA6jvfKQsS
iW7PW5nay1xI5AdRf5U3Kxs04dUuCCS9oOtuaP6CPecaGhkWO5nYSWqH9jiITpAX
ERsm4e97v+jF6LG68Rn27O4RX2UdKvT9j7b38lEQzdLQnwyE3JSR7jfzu7U+F+RC
ygGXTwzATy8KJc74LiixXtFZ9f2xmT+bp2AjlYLQDmQdJVUwu/9e/MuAnZ7GJ1As
grR8vlcjqi+YZ83F+HIPP7Vp03fTOcTqY4zb8rgiOGru4MWAEnggcdUVDyq1GaBZ
p8bHKYA/DHevFGpz91ZaEiaEkRf+Zi+0FBFwwb/DEzmfuGyopOCT3ubNOtLLth1Z
1KXUyJ7Nr/QZjffyBrDLrvNlEUgph4oaqfaqXxvVaiaoqpa6uQ7JKsrFNDaqRgb9
TEgbZAjNpXjwm7BNFFadpcNxJlFNIIvkiZaCnvWYUO9LQ4p+AKzn0DYsLLBSsxTG
h/1yDsLYDKePHlYgV6i/x5NMSCnKYV5qINybJrOvpm1ImhYVCE41mtJZt4iQb8Nk
BkoF6cjuZhMiEE075FFNgfYy3Dt8oxGCOV1NzowlBHzQo5tG31jARP2YZCicbQ6d
kpt4rVgfOFNQvHYiCIpCXyi5As6tWJhW7xku+xO2jcWKzCcnucl7xIBTo1wZTeqa
VaSrINIWvKgIL6e98WqSUs/QgyOmiBPcdMVvgEs9yY5pZrhoZFxM3dWI89opsWOh
XG3zuRvmq/ugH0+a/uSzxqhMUtJcHunTfa912gODcAYc8JA6n+/LUlaZ38/zDspc
HX8XDDrI9n4NZvbJQljwHCbX+cwrqSQIwalY/fLSkrd4UW8jFnNPg+71ikpkxPhN
yzIS6a4TY43moYzTIwiO5xb4on6wQTdmUlZszjYC6oG2fIUEo453Onrjrkx59kH4
m5v+QqUhw7gYa6kkSzaHtK+rmDxIQjB5/O2HgvvEgANjNddSitSymJNR5mqsSOxf
RJ0I7V9haTHub0pyTVw6d+Lxjse2M9CAjHf+dV7fHq6koUYuVSuH6FCXL/1c7APi
+PM/88FvFI1YrFNo/KTzfFjCDkOgDmKxL5ZUmkfPEiFKRQ982Nt8iGs3zyOoQIbK
PIJ/UiUoMA1PdAsVeIHIVTjzmRXMF258H8Lj0Ar3P+xgebfyKaUS/Fvlt2nquril
OB0j4XgPXjBuhFc9sT/y42/wt328LmWJJNAGP3TRfJzVqGQz/fFe+ZFB9sFwMi8G
205b8+h17eSkb2MHf4ljf3F981wQlupq5cetA7RYIR6M+vmGrfUBXB/HVtHHB4LK
sYvIF04oOYbq76L2HjsZxW7d7i3hE6EUcEwAKmvLQEfluS4nUPzDNeilElGMcADq
RmBS0Vuv9xPI3/5xF3H5h/4UiasCzZrsf093pAObMlFVDbVvjf4wBDTqb107tCfI
dq9CnisHR1WnPPmDOUXPl2hkKTvzOQvuabpw2Zy4qwmzRX2OKYHayFh+DsaesYyq
C0j8mE3Fa4n7mR/I0oAayRXaqMt4zF40w8fe2CHn33NCmPQ2+mvRiBKeRWJxbiCC
cnM8UlubbeAmdPNs6d529Bp6ntZzzLlDiIhfFAEpT0Eo+lji/25j1Ar+EiIglsbJ
I7UBYRRCNEJU2rAOS8PNR5KGHMgbts6+TS8rSRaJ8XMPSP0vgB6/M/YvggRaT+in
8bTmMSkzV7F3CJXOwMzqsjBhjENjqqHDnrFI2qVooTN0KMdV3uzitY1Pn0Veiaka
XWGuwSz9wkqo070Qpgc8F/J54x3/rl7KE8eVAurznGd6UoDy+TZ+e3KJuzH7JeW7
vy7HoqKZz4DQYYwFV4R+zoPi5tPSFn9dDyKauBojCdiScFQVWdVjPkmpwsMSQ0as
M66FS6qD0QaGpMNX7jAZu5lZrseBzx/bEP6TzRD4LcfhlthbHJWpYUKQJDW3doOo
1zwZSiiUYb3vY9gM52kypQ8pHdFkdUWJqLS+v5ILEOXPRz03l5X52kCPL9AWA9EO
/vbZJRtErxgXkX87U5Z2SpEn8M69S1Rh8SJ9NAzFibYa1pbWIuyNaBLB82LKdMij
eWi04y+aT1Q+xVhigkn/4d/NWf27I2EQHRESF3Wy4e5Lhv8RO9C2YqIgbXe3tOGd
3BS+1zFB/8QDhmx44DgfL3epnyeeoRWI4hAzMSLwF/zHASnhlEO3hd9eEApvkTU9
T/xEnlqyGE7KCsYUBV+gkclWGpP0shXz2GsNuXBDrvaZm/4fgb8hC8WieajhT4Xh
NRcjcGx4eJmeqNugp1lUeWOB86twpO3okL/l67B05om64fyfTq+4zlaFRitRgNP7
261KTZjFOl05RLsKG+GAPDhAGtBHIMN1FibNdKdDY8opYU7GKvbaC9EVEZXuACul
Qhgqx5V9qD5lJl0alq3W6AQhIxyMCMGAyFfEM6QzwicCi80G4grwLe+hNfoWt2Mx
TXdtxsbzkbji9tVYcc643fmLEm90WzfGPEBrdmgdv2b42dMl89vWeTLlVuae9j+R
ARej6o6+sCEEuCGi/HFzSxht2crF+IwZ40TNQnNjUUMucELvto9DpjfI3uz2+zNi
AU4ZuoBjSgs4iLtH7JjhC38BGWjN4MHe1829mh/Mdj9c6T1ERE4eVR6zZeJ28jRL
/9yW9W6pKEId9FJFJ3TbfHU0wTW6JD/hOLQW2ciumWzV7opzu2YIsxk1lq1319pb
UmwXwYmKBD/8k4tjXhZObDbrHYswWYWSgaXpePU9P17nHzPlDYvWV1aPBTV77pmV
FhA1aA6Rdx36pcpFCXRDPBybBhHzDiTv5kH/a9WBs4Le93kN1fglUYFJIoHoTxJ2
T+eXAiULvbWreyK0Dj0fwpfwbgldJGlMjMokw86RfrTSuFyZK2fg78iPqlnw7sRC
IOkPFncd9h1AWmFJ5rVCHTjtnDweeB0qJp7Lc9evgspVahbC6x3Wskf35fidzuy2
kldnWx8g1EP3UZAQNuf7iR94swPnEuCzcliSIKhqwaRXPCsA0HFKayCK251p0GLt
UXqgChXF0ccXUIyRR+CoV9hcC2I5aFu5dmi3oYjr1tgp2iPUKG1sicjGNCfIIu9D
S2z1lzN8Yf2XYnP5ynu6MrbK90HaQTwdfbmMfEQR4MzIIrvZGDGgBp438SE5WvAD
ijlcQomphBwpo71Nu43DXVQVlJs0lK0iREOUHb3uCCSE3pXYMSLa1ExKAw7E19zO
xexEtCLswg3JCgkaUhbwi+4CuT0eHE/yFst5B9bhpVY211+5ynHS2bVDXzf/LvbI
mXSlIdZWUCpCYGuiYOsoYkx12SHgS/13So9ZnOsvuQaQEmr674HmCe7ZL6IygmOL
CV/TEqxgq52MwSuOXqRXzLmzlh0sYeeLRx0vTUtqSpGfYPIAmZwo/Hvvg2bSg3ZQ
S3tn78b1lho3HzLSErEvJAwvXfp7Yj+Qomb8PTuqydmsG/FF8XyqzQdFgEFYWyLP
Tw9cA8OmllU2JWFi3y2+hZuPJNox8s4qxhA+D2YT1rGG7/DpfEUex2ZDh8JrH7pq
liTsY1RQUm9ZzWRW6KSYJ0qM7nf7sqlfHM+76TRxbmH/QX6LKVCqxnIWInuk37+V
9lWmvAoruh+YYUlN9grm/NxXrVEB2twahj9B9u4cEaSZTRZDVB733Zn1jh3XeFEh
jeomnnMmTzFD7W8qOElt276LCqxh0NK3msdlpomDT8rPFEyp3A7EJRdncmQMQ7M7
He6ID1BhVWYtXpR41wfc0UHNkxw53yv5/gWJhgD+zBovSxJ6cVjNtR9nDBypUJyV
ZqbiL1JQDuTOgmdWa3+LNgADqFulBBFtHKpaUtNqTiKZQ5y9bNXGFe+pjmJQ+lI0
+qjLg/dqmw4sxqazHqI5BK+5KBbWaSjpOIu7dtZThlnQPJR1XqTNYoPNCygKWFBH
dKzjVP91g2e2nExZVnh2lgRy2N+BRYR/kjVY3OQxThUT6LuYNTCAeoO/ZyftA/dg
pUy2IuIYKoE7q3m+x/KGTnTUrRbJTFjSPjiPF4gFUHxmSBF/c7LRuoA3gxj4WDof
Sw8LIhwF1ExGqTO+vHLu86gKLokMYu1Kk1glfO4UGESqcb6KqVQfE+0fSmzxmM04
Fnbt4FimOGsSXQalKSGC5EYZu7+9OOP453/NLxT9VWJcCmLTDYsfGvKdeq04vQIi
dKqW2vzU1zeEwZod8CqCKniRwfrqP7Nx9Ah5ePkMzv4knM3vojODmgrJk2anQ85F
FDYuyyxSnA8g2j8hjyFRGXlJO4TGvkiaG6aAxhjL8CBVzZRKitD4gDvvWXQHMJlz
ZmJvbjCxiIgbkJcIN3qApdp3Yhg+MBOXt/41TMSeSquYJlOHb9jOTb6b/9O6pams
1P2KZH5a2K9yCHopEVKXkoOZ00lEhZCd/zOLMVbXsAFPGlrAI0T/JFJvzAwtMK3b
ir6+Kg4YJq1YcCzYac0KNGHPRyFkYvWWsjSKJJXk//WaVo50A3nLQV2RzX63/+2k
t3IFQUHA8kGpB+U0O+hIeLaXQe5ix6iTHcxJElIBkniC57XH9Lr2hKfiVI9TDHuw
XTVjf1WnUvX+e4mCsQo/JxE+xCm3PJ7l+qDkQhPGRrkn62CfmrmLhAGPXshVzk46
jVNlvOH8tBMjyfqdQgAUqg4VheGpbT/5uOL70cAhaFNcBJwlpCB8Wje+MUR0CT1I
d9ze0jK9vIxB1Ig/VR6O0AAG0cgDMmhYQYjXgDgLSY66VuL1OoC85DMEaDxn+LfA
1uU+mfO24d6Kin4xvEDRq+o+XQQ5/sJDQ7wBGylKwi+SoOt4V6yR4SAUR6HFYIC7
QCxPeRZ+QD0RoUfOq+oRaWjnhaWJXJCTjm/y3KKQMyCNkHNiPpWy+MJfZmZNf4nC
lm94pglCC3kprSyFoowfHAUPrSl4LrfTHdnT4NKO5f4If0c0wmgr3zelp+UlK5uF
l14b4rYCr3Svux6ITC67G3mEI7JaLwflJ8z6d2sADV3XyL4M6EuJ/0sSZV1By9uX
sdwwrmAGVcjYvFdnH+SA3U7nFgoIeBdPK1JK6T6fTn6UzSl5pX7JUuk/Va3+eo+x
0+2NfTlbRPPNiUPNSGhnVJqoBsR/H268mJdurwCuwRYE8cxpnSJNfyazqKNJCt0T
Hde/gAjGH9L0oD4i3Er8x9I+RExxNYwWViONhjA+2XOzjBkXWYPZ0SsjQB2Rna9O
y3G5kBRkKZc/kYfhYPrhhSC+pMk7UD1om5s5rpcTDqCohIMz6j4ZxHlQSnKE0Lc4
hRFGznOlkPdg5oq492Z9ittPiie3UcxKtncxPmMyVLnmbr1Q/OInmH8fAk+mFGdS
bFJA2iqTMDVEOy5hBY7yc24uHawqiouq8sYY+LN/FtGIsJvM/He7qnFVYQoO8E2M
NG3o95pQ/Sv3t1K+lZL7MOu7WVj7lEvFnutycBGGubntGZ8L8TQpG2iDEGrBH3aK
GbO9dfO6rPqt/ooXBKDx4QQLtZlioiguGhPizPtinvlefC4ut5H88pADEIUhj56z
S9jt3EsbkFJw2+TorY8RALvP0TvvjUjqPul/Q84ihZSlz+wmtJR0KSxuvxZ7aB90
z+G1bnS9ezfEbKmJC2GMc0bM+dqpVwqVkL1G7tVkVMWLFXAS/fkw2FXo241iYlpi
KI23kDVJfABNQH79Rl6dkWFMAgzNBqjvKc5IgBZgRgboend+AmC41XXA396rWV6w
WlQXsEoh40iAR6bdNMuT9ooz5aBvvX0sGrsXOHOA4vmiOZs/lEbKwMNY4up/u5la
3bx5oPNBQ8j4Iw0hM5M6y/N/sDbODln3UeZZPXqEYqPX1sh7aSjoDZrwB0GEfCRL
PXi/gHJuV293kE3tUXIkMtoV3uNZfqEt6NyP4+80cAMHQ38EHPiRLMg/788cPRqk
KXXbFiXVY7z700XYSurL62nooLvA18GXygW23DlPfrJARjGPG9kZ1bicr39pysNY
Sso8pLWdSGzAuZLC9bz3LFYFmTWued1rcdOHQ2IHdMbs+uNqQNVCuUACYAZ+rjva
pb1a2rjhQd7r0DBHpvyCZQ1Vc5Zq8GeAW/ZeeXiPPSApLiN/+MfcTYuEbeYZHC6N
glZgJwVop7AkGrnM8p8E4zQHBcVF0mGa0pEy2qnSE4UMMCFD54O1pbUnDW036T/m
Au0pUVnQok2mX7sXTXlnDUfSfnkn0d6hOB8fMfOPvrXIBkq0KHLuNiPL9gCDMGRa
R8u1Rz37Jn5K3eDV8s/jpT7HPtySigsSZb5P75iHKMuryf2sBjigVQCPXEZZDvNu
3oBK82yApBuN0ryvmMQ4HYZIlm2RGn4xwxxtSRVjpyBoyxcWKnEQUnP/5racIXRg
FaoB4/DXnlkgMEoqpFz8U4DAzA3yQVEcJmy+DZR8cyfAHP5KzHTKK4gTk8wbHvcM
4eZnt29Y7ATBhvwTsJOMnsnA0jQMkPfV8q+nIPqeVR4QkaZGgP247ALTBcfM3e1R
MPK6jSnzleiCxSe6WSoF6TzIgJkmDoBP7ANr6QTLmTKH+lUg9Pa9F7kCUdH58mb2
S5St2El2BOC2HsvubDZFwO7PYpszyRdjfi7npaNPMUlC3sMTvA+RCHfNcqLpvkf4
y+cqMI5ygqHf1Tnu3BXJApsnXT789wc/06yCXCneNNlg3H3YJymvM09GzCJ/Qlbu
nqqaHmFDj60w0JqzfFm8hnTCfiMC7Fy8gKS0s9tLQFDlOlEuk06U6O1curAVR5Cs
jy6LYxP0ybugVTN0sot/LtrhPmuTUoFpmfL6xpRWu+qR+qBnentyCJwpJFKAjoaO
cS7B/LpkBB6QjyJnxVzPzVYAR5/z7/v34FeWJKka1bS6u/enA/80XnRl60fZ6v2S
ZwLrgzU/+uO0TwgKfveUvpgdyrn89GrPf8KA1qQKbx4VLxtWz7Rhmv1KuTuNrSK3
rSsSkjmXQGAjU8pITL2qmeM8ncIglH2fN7923N0D1RR6wjxiCFTYzc32T3l0NlqW
izaLWkM3WQQ+GtyQIQxALOm0SuNgdJX8/J09b+/kjJ8NwrqKsEudPFGnU/zxog2f
unssxC8bQzm9fK8frULZ1nfab7zJiPChOrFRJAUXuXhfaCc2Kpmp51a54OoTyh/G
Ane3e16QIXRrELsT8ManyfrjReu3pGNCYBNu7pjaCRyAwF7AWVJ4/OSVmU0yweSB
zjE/YB2gJpeEe97qPcO5IylcSiIVWBEXtN3ZrFVYSS+BHt9NWXn4jun+XwNsMpxF
UuyZk/FahAgvu/n1Y5RIRueoFMeJWfJMJH9hMbdBwXG7c8E8slaSEbdvKFNhxPRK
6J4sowuxl0xuyDRRaYeyVn4t9sMr71EAKnh6FYzfnE5ygNLMreh9s5FK3ohhGkAu
KmYUw83arnkoMH0ym1up1mHawSDm8hW/AyowyG+LeO5ChiqbNhBEOTyai2BaLTF6
MWldyco+56rUssx2kICz+95pNm7S02J8JcefAWi3Sulb+a63Kvw3x3RKxng2+His
VsyP7jSW7KOoGV4SDYC/3QTOSx5phT9rysO1Jm8+08EtEe22PXKsIViiZPsQOe8+
FOLW08TeVPbaRK/eb2IITFPt9rUyy+Iz2CbCgMEeqiCVy0wX02fDd+Wvu7BF/sAU
ObF3qeLKP7bcc4BUHcFjDqkeYvvnzP1yzKlaKClulbM/i+57BjozUtqq500gIc4P
4wr2P5zHWyuIPdreAOCMgjyf2UpPs3xd6Z2MqoLwUnR2huxXYg3GapSGCcfbFvU3
XB5SfdNWUqz3pyJ2XhANFgZ4R1k5tx40Y/cM9nEDfhqdmJErQpwyuzvk00sB8sRu
KbozmsK8raYvJE71zwUXzKRvyC84QQQFPwZQD/8pG92ScimnyugKiZwuh0qtO1gt
UaBgvN8zYkgqM3a8jj1VyscmphAfd/yh8xR7w5eBTTWc7tdZNEOpV6VBcL2k32bZ
o74Wnz6+L2tFXawAcVLv66SbD9EBh/6n6InViBOVvxeeQv49JTTrH9jRwprtcL9z
fRWSJZsjqt66F6hTK9/P3PW1UWfGloSXhg7JDvFKt2Wqk1JSD/TMS7a2GVbzOZpR
xxffi5Rs/jvGrPYNlsMkLlQ1/avwppJS1eoGVEetldkcvnEMAy4PdyO4vYWFx6gZ
n/WxK8O8awsEHiaaWR+yI+q9kKjJwt51F/ODJ40SSU32kGW4XTU1B0Zy/JSkC7Jp
4g5v8iqyXTw3ZstikhNrSC9NZwkNuefutyUlS/IV05RIni+1/ssmOdZejjKRM0H8
TQCNk2r4xuS5hP2LyhCNqVyx/OdgdyRgfNP7/thanD4IznRRdA4x0w4pL+7M5cj0
oXvwChiDI05fJNNAPsOGf8hnxEn6aKdFCMqEcF3+oZlPZtjEJaWdndHUuD2UXvji
OI3FxdrIQObwhZaLUb78xKB8xQXMvETMmWo+av1yjU9ZHzr8i5GX3YDE6Xn8s4NF
Gyc6XTBIfoWnMYEOn2vEIcGXPTeVrbxTTR29qnki6cnwY81uF5E8vPnrk4oLHyz2
dUxm1j6fe1AohMhIFxcmvn9fsIQy0tOoTfCRuCp0s2Kkc8Fw/28t4l+Ffmvdhi4m
8vyd7hbJMK47Q/0Yoq3LatrznghBf1TL2b/Srko6HW/iewRTPCzRkKKkNRg72OC5
4v38Xjx9Auj+UEGOPENych7mRClkMIC+5ImRH0IDtgh6zd23aqHI1EORCHRVNIzV
KKe1dv9XRlKYuvNoWd/dD/Lm7RyaZIFxrq7cvtkKmY+DCJvB9Toi0mguVyvxjA0h
VHc0I7eVM0gvZzMCFrbq5ciLhZ1jPZHvbRFuU4vznWCjFCPqWaiUU+wI7jHgGjSt
K6f9/sShngXK1bHr4Ta92vtKnl/u1GGel1g5yD80fnZjKTZ572L3idbuMbmtRhnU
YJeqpK8hjrkGxO4roTXJ4cVnsKKTpvqdBn/tP4By7Ux47nmG95Cfbfpyva4WP/EQ
6igAVwq9c+oeW9gwt7ACLNnKE9zXEj2UcwknJZNMxeydeIWX8QZPuSUhhkmcHi6y
kEBHGbkFU04o3AS9pfI/uAsUwMkaLTRQXUncvmIk1GrtlJFP35WfNUzi4QlW1xvv
DEN2wHrl2Im3AkvOjBP61W9I7O00AD/oZhT4RBqDttSVicvVvyXm29/ierTji9og
JzbbGaKV/I9WTw9IjQjycgYNzMKWFnJXN1k/7r38mPQxJ3FB78C8NJ7ZaHExqqYX
TZnOaDPO1JsVBCz5Gbvyp9dU2s6uXem6Y8CI/S2wobjL2tepfTtJyJ3mSonPMw6A
xxqDJtDtZ/H2l3iuo0RAKNex4JUbCsrpLhemxez25bcI4cj14CFmDNDrun0Vqvzm
7n/BCJk9SXGw33b+uUQMxmR6u+bPOGcI820tFQv2Fc3p46jKpdUSUe/8Gz3NXaKy
V499mcaznUkAriVzK0pC/SSYN5ngZFj+gF4CNJsPSq9z2QdtFS+j8tcm/YOM9z6z
uPrx06ixRnv5YP9jYJ37a7Y8HaLYV9B/fH7YpGiaa2jZMjVJ22o4aJpY8ukJstTk
M5X3tJlYG0WtyLoivpm99U/egaUCn8wp8HGQHYEufn8kRtG22ZTVF1K3ggRV1im/
n/KN+rta5FSDLoGdHGab+x097wiotqRJLsVThuzSrX7ysjQITxDl0pQRQPhtEurp
mdmnKPkOrqIz5Bn1OaRuhdoeIFHMMjutc3OOAL+eiepEWoW6CBjrv1Ti8/v/whFe
FKj9mUBipLVBtqNuy8gmqnrdHO1c4ITTfcb+9NSx6sykFUPHSFvYDR5k74s/fFPa
/ix/ViwVNuFkJlekcjmedHdv8bYPzZyGa+Gpk/I5EWRUnMyY14epWT/nAq12ryTN
FSlvKWgN2vgO5u8KI/tPSqzi2PcyL3Of6ysV79Nfs7cj5ev+e/5jfkJu8LHWv71h
IXd3tWs58GOpdn2Ttj3YTGvr971vtFAwT8E74dawHx5jgHdHO/ijX9LXeqy7srjE
jo8XagXf73tSQXQzR9/4duIIovsF8qh7EMJsmJPewTaQvZhc57OOBR7oaNZ3xDwK
UFHQNeSEUpQyW3FYyy+yA+hyyUUouUQt2i0Aq4I6/xytyK4oUR6YanhiUXjcPu2N
BQm5wTg3d5FLaRK+WSDrsnlbQGexL9rGybRev0mzuK7Ph9ckXVsF6p4MGuCgCBMu
NE1IWBIol2XTFFmZNQzwbA==
`protect END_PROTECTED
