`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/UObQeOh+hxpFoXia+X95ITJ65YU9yCr0+5TcwXFvTY
RXW9KVc+zqkeP62hkyPNFBMbLlny3VCb9Ptvn1eXLkhypwmohjdjW0W6ROgCV9Qa
MoST30WrjyXkt6Inr4cORn5JpdRFMt3TbQhV3W7DLar7iKgIRv7LjCv7gPTx+hcn
XcMVS3fx6OFHPAnNMbcd7S5BhbxSjkl5p46I/Sknd9TE1xA/AZGIaPqc4zO8Fu4i
ufAVHyfuvG+BvRpeF7d/Yt6Zeff7qy6tcYtpMzHPkVY=
`protect END_PROTECTED
