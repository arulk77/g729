`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Vct6X93UXGNo2dZXjvVYgxrvDsfp1agxwjj5cXn1D9fUp2yzB37P1SvGTnmSiXvy
N5yfYDzEqpAvUoU4ucdZT/7S1aXxUwdrA4nn7dl7KIfyyT9trtco0TeMn6Rg+w0c
Lr3mR5xFZCqCRv2oZYFccKlfetjABhkNn6DsOoMgJX55wUm+Mqogy4w56wcuv7Z3
2cG0rB8LSU5ga33IQ6x4UbawVxgPKhev590k9foxjJRqMRESV4oYFTKtuLBTKYnd
V+oGNalcMyysY2DAX9oQU66439S51kbKXI+BgYhQLs2c/EAPGME7bhWClqY9lZJB
jaj180nDNdxR3vCA8C3HoiZzKM1cEX+EszdQj25Fh0t1JkxjJAdg9CvVDvm3USwf
MIzo6sq5/f27rl4o5Zvhoa5e7UzaNhuxLmTDLdK4v+EZipVyKTQpHmOCQvOMpeed
zqILMhTPAxssGR481SLRwEGkfzW2+rqR3mWv5wTyaiu5kcuiOglqMu1HCasrRxoX
KeXC3Q5Lp2TXQFp9Ch2trf2415jgF4mOEumJTxJhESaemtEMVOnIeiGQzpsaKLHp
LjWASqsSxGgupYrxyCkOnqUm9NeT81APHov211wwnwuf3RgFp1cXaWnlJHLkp//Z
1WRsMdA4W2OauKTC8prjEcI0oLeonw2OtXOvw96ioM1bn06sBdlhwSRa5kv0oCQP
1e2wL/SQDrzuD6Y8t4RmAw1otvOy667OFIlVn7MuUJNMIXWXeQ+4GUplR3NMEV56
NjfMXsCDPaA0oPv9JVEMxQ==
`protect END_PROTECTED
