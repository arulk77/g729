`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2RtTiaLwZbJSuPbraFO4dgl5M65v6GsZjxrVRh+/eZGIib/dm5tSaTPn1ey6jyJ5
+T8IXzs9aQduKF+hcF5ufj20UW+GEK9FUf/Xlgc6dvuJNJFA54NQdo89d7zOGlBo
LplPyaxmTru0ZV3f4ELFVaIDRTV5nbbjpC8wFh7Zhc8UdTpcpLtcADDIf/BBf1cW
`protect END_PROTECTED
