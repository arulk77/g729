`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+9iB9xSzq8G065HsDtnVQLkENDsgvBsr4lt84e2P2vl
NDDPmaNc/4ZTl2bwzu1Iz1w5Oa4X0bNIOeawXvkTZp7HC0hkks//SCV7lYmlVQfy
eq5g+R2kfwOBVEY+CuCebynR4XINWKM5w9EBLpxYq9XYs429SvcFGl6JxMdJsoLS
q8ilx23zzUVjHsaMh6NLqfv0H8jbN4i+WVmq1E6Qi49lusNXg3SqIo5I54PqL4js
214pkUZe7tzY6OG6a9N1Tw2DzqFB/I+ZFSS3Yr6Q9Sl4WIQHZ38s+OL7xfgsOaUi
JHPr/j2Opd+VkzYBxjsaPWlqEBVVHAYPrXSzKO0smWVpHaTMWP+paY34L504adX8
kkgpvAgLL8oUZY4JxP1f83XNRgY/VUMpsAhgkFVUKU0MWY8xc65H/y5fHazTatWt
Mbvu1S0ZOaxNCOkqFc1Qb4ldOUQy2q7LETPn5t57usJpdjLjZdrOefxLzl9G/mqn
`protect END_PROTECTED
