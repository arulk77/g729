`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePlUQmcjBHidfkQRMcCFK/aSWubFxP/st9fAE9ZMB+Vp
/8o1DioSfJ9yDoM5HxorNwHEhINELcds5JqGzTHFQD9LTf2dyC+YKuFWiXn0DxgO
c293TtENGQp9rjkfcOXbWV0X2hEOV1z5g3f+z2/1P9yAZ4jDkr2rfRFscNjTqF8e
mVhNLUbssotCcm63LB1flbaZYkaA1mgnCdFUzJUMLU+0nhoWg9At6s/0Mwn5TuhA
892wQc4Lmmj60q+hBU3fHsoRI5/W6YWpmvz/cVt9I+rklP5u6DNUVXO8a4K0OpEE
r9WNY9hmstfz+8CqFbgMo60MmuGDDfGCSlIbZHWlxj19DhqdCTA9ML/bAnoz0paZ
8E5MwK6bh/kQQGD0OF632SNy+ZAInR8neGbHVCgq+7xxb5JtYwcnqI3e+FJeVM7w
GxzqejQOYLRfC0g4Ub5JaQm8RCd3nsAznUIxG2JFouvidyFACIGcDkm0+3CuWhnN
SZu3OcSWG2fsNJaJeeXONBOm1dPJlhceZ7FyHxtu8TckGYKRy1Y1lO9O6Mh39hgi
`protect END_PROTECTED
