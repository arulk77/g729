`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
e/hYIPNUbQ4wn7NFLKWOtyTSs/Po2USYXhaRAsRXP18RASdhCkoR32y5Sqtpva41
ORzxuCBytNtrdPPHRK+0/lCfmjXsWXopSAux62q+vMu7a+3B1mg1idfN3ZmIDtpW
PuoEmLtrcsNYQphnfdzDiPBWtJbW1XT25D7lF8NZcrhrrRSdwePImMv8YXRzuHo3
S4723/ZTFrAn2cMWeRZ8Tt9vweB4bEPUUBMgQRUbzsS+ooBiaQwoFOEUwFwuagJv
Zb9y+MjxI/KZ8jhP4l06VDIxoB0ySdWei28O64wzS0U=
`protect END_PROTECTED
