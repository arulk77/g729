`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB/9Dk+utb3kVt4WwfNlE24keu/3XwNCGhMeanBGpi01
0O1ZGRhzTOa3sPPx30ykzXG/jVhhDJDH5t2xlWHBj8aBO5OvQ/vH3y6FknrUhMTK
DDB5Vr2fZp8TaANKGeRsFeGjGR6ZVJyvkmBfKQJjYZqqUDkKNg4upMILZ3825ZXS
mv6Q6Wr8X7I9X3E9wTnWAHOl18DjxUM11qqQCMhNAAkmJ2DINMj+U1AHilbLQs1e
`protect END_PROTECTED
