`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCSKTB3avWQEdGkKs9LLKiJSih/AqZFUoHiH+SC1mWL+
5pmOLVETpvuOU+/DWV/J281U2zdNjLEZ9oVKmXIMrl97P9mwdjmEWnlwgOF6WTkr
RYUkrwa63dFR1qzEmC0GnorbJ7Xt6P4LtBF73axc+AjXuunacx4Y9s5Ltx7wOs2o
XEldvhOzzJdkEJ5PgxPjMjlMFYaMyak3ioag/OzTug62vztp9WO4AhHqn/IcWAhG
1pSoVGVXFiGkzLzKNmqTtjIedGD6CoK/5bm2lnhLLePAEa6t0gbwqhhMsBI19H+7
F6A5xgA+N88p1X95eW54kqNTkiESAbSJHEzhVVc5xF2ph7jVO46uVTHnMmhSWrti
V0GiCa0onZaT1ta7ZQeKCtUXgh6aR+FH9H8FcSQPiiIhbFcLPRZxiN3z3ssjYflo
x9bCjN8edn1it4DZjYGMUA==
`protect END_PROTECTED
