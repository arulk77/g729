`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF01Jwat1EO1EVUn4Q/djWV66Ttn2zXc2g9W51CvQsd5
X5mK7VQR1I8S7Yvnszq40QTCQLop7ojoyucONJ/G/z4vkk5/hqIWv0pj6i1AWD4T
2STiROADGS6gJKHWrBnMOBy2MsFBinFKsNJlrNO7tN97GwhcMb6u+E9IteAEeE8u
r5azCCFPGmVkiD5heYLFcc147bEqqjXb8Iu1Mj8D0FY1Ii5+30tsBKUsgBIFSA8O
kjdmiHy9b22rYq01COX57GiYDAogdgvaHrzTWM8ANhKdD2t1iuKCHaUIEYScEFtV
7DFP75rHtrlD78Zjjpxypc0voT4roBo5OASIdoSv/DQGQyY+ZNr/V6JQkz/k4RXH
NTkVSSJJ06+cN5SyYHNdJIZsr8h4pBLoFbVSl2RkhhyENWxKxVqjgPF0CmujTtm/
C+730/xBYHjTcVSGpTkWExW+SiayyyxrduW0KEpcOooU+l8+ptupya2BBA0Cf6Lo
LSiJAaha/JqSiCQrpQMA8tqh2p2MKsx+sVJ8zyHstdiSS40F9FhYDxacBKPnN9IH
7oij8xJXsd3PPlgxZedFBA==
`protect END_PROTECTED
