`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAlESl8GttWOISeMW3hXFOc6lsen2vrjKUCeZ6RuXRdV
EG10yqXm2u7yBWqBClLUiIDRaD8BIYImg9LEDF42AgNvSixjYs471xWhKAKqhKrX
Ww8yQzlkYJhGE0K3opzKfw/lmxizqldhbiVT+PNCNTCGPVNxnnccvAptWVMJWJht
Mj6BppsHpSV1RdCoaVaQrCuSwyWYIJK4oWxq3q8z4QaVQpldIyOY6C4hCe0DzeYT
`protect END_PROTECTED
