`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKTbczoqK0e3M7TMX/CptG+a2sAFSGVmVZ9rMC+OFlaF
xK9BJYwNA9qHdf9pg9EMKjvc7XliFIc8FJIKw6WTr8XQq6blBzmJBijzCrfulsLh
O5dxC0nd0rM2x09lNVsRTjUGHQE/eD6UwnZlwvoknfHj28uHXYgr37vBXq8Thl/R
7UR13PytyQXr0KlHsKcDPg==
`protect END_PROTECTED
