`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJVnxtA5K9/QDEjz23A2EvMeURvjwrilQArAasK6Hgsu
3vczfxLqsdfk411OSFEZnMKXMYgtnVZOuKLSfUPCUcwtQS/p70whcT2PYmhDizli
hFKHoDvKV3UNUBb+OzMhEOgXHVStlfdf4PxEdg7qCoDxB+BpL9ghwVAuh1bHyxLA
BlsqqV/3V3dHNsqwuTGAR99swVTCtDlS379bO5f5gPaaE1AHtj6J6y+r+Dw+n8ED
aR87T/EW5jgCP0F5wFnn0FigTTVAv8295BFuBxnJwpp0KsoG3EtOPWMBmjX8YqjA
`protect END_PROTECTED
