`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNuyViMuIQT52qndOTL8njFKAaCwole2SvqiYbRglNoN
oPBnipiKXKekNJTFIaTQ44v0lHkFR8C8pGcWSvv6AzwYFGsscBabgcGK9J41rpie
vc5+5hFtBY8YvjXtzUAwvIopXvKHj317wvNP0ZtbfpN56MqqYON7xvKueQ9e+9Hh
JY9qPC/ATMmUxx8dCTFTajSLpZALg5+D1zBxFbIDha1boAM2t3yDtpcTib54W62g
ZOhfRjtvu9NrrHJeRMS56Np134SvUGb/lsHxX21puswdLzsyEOK8s9qpmjQJbFVA
yPP41pKJ/2nvLA1UY7lP5w==
`protect END_PROTECTED
