`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEnILVuaCqGJTIyz1iW2Yw0vzgZLokyTwBsC5nEhOIje
izZmootVC3QwarEjgATEyyMOYjsH9n+6JtsWl2BbK4BA/tFqQrA9e4cOwMxe4Az0
9uFY2rZkfSTE9NXC3nFdfUPYfmWEQZSd/FQ7+Ywt7qXwZ0vZZ+YR6ruycjlO50BE
h5inV6GPR4YmzwE3+jdd03RqedXAxRe6V+T4MimfS6TL+zk1ohxaFnka9+KE/lf4
SDveCgW8UMuiZZhgWB1nqatM8iFsNh+XWzaBbK+ckATpZH1hjrIgxcLM/J6enRKC
WYZCYQlNXaKT7EdomBxQQpuk1ZSaRsMKwlSVXl8RZ8m8BoGO3bECMatIXZ0RCTdX
dHRA4PfBpyJD1USpmiV7C5/hGs4NbOWigGFlu5oDah4GBQ9+OfuGBNGdKvC8k20I
weC0rgwt54XSjmIWLBny+Yfwj84jxnhjc5Se2GU/D77i/n6vhScnZzZZxZ35ipMv
7UzOeFUrjnrYMHipLugkoZu805XG8t8Mi6VqzT5+QWyMo9yPNK7E9A3TrapflENv
8ETQYCcbdpCPWsuZfFewew==
`protect END_PROTECTED
