`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFVrnouHVOApfXM4O7zlieQXGJl8IpQiZu/IwdhwMONQ
uvUboTg7X7EOtGOjRtyD5p7W9V9GQuWjRUoGkLmV3Ee2qhlx3dFd3QJv3Z6VbEjN
M51Eo+6P3m52vJ33nqaT3g1EfKHDUg40EQQqn5WWBF4OL4Bnjko2ws52YPTQlwxN
96wnlX8JO2LbMllYauyC+W7JXqXuwSUsppYJcyKhsbs1C/62Psil24gmmkX0cncC
IOU1qfasq9sY2K+U8xukMsVWBAvHlQAZYxAOTo0YUY3d8eDNa8AlO6IVUnJTwQcw
iqFBf0DsCbRyFWs3JnLMVLdYcsb7uwkqaJDyHR6hBo9dbL26q/U2klhGee/qPDou
Y31MvXt/rNCzKE/mGgWR5a12x0JhgNQS3jakthmIu4E3pWTobqSMmmN8DULPTuQO
AvGHt2wG0dCFJnkfF8wdnduLgHli4jtqYlu66NhLs/9mW0Vy8HVqynILT3/DQt8k
oNS2LtS89QRqNkIJOkHo1XWA+IO8wDB8pygrgNc2hRj3aHCgnl/E6zcEYczhdVqt
`protect END_PROTECTED
