`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGKYWfHFkcLMv960107K82GRIyRd4Nxm9zNP8PWusK/Y
u6TMSe1XOc8CyWwMxbZOw1nKhxaOyTNY5XKCNsG7/gcK2zjLEP5n/aVlaAeN/Wh2
E3Tc9ghxzjtO9nlrGpb08HAmDmmi9Vt0Tw5xthfiquJ7MTtpS8mGz2IUptf2NDmq
sQy0Bn7iAHlwbGdq3lwrVdhU21mMGglrzhMoSgOL7OQBZtH+YZ/z/BZuOasrZoET
xDMJwy5RimMOZ8tOty/FOmEiBpKxEwgyNhr7z5eAoSAlnYpXrLlcIJvYFtnZHRwu
QaqkdU/GTqur+8bM4jMqQA==
`protect END_PROTECTED
