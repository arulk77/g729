`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
nAsgBJeZJCxyVzILs3oBlLFUHcexnzdF4z1J86taF1bh0N2KNaxGAQ5Y8D/fOkhN
t6eKl9e0jnqJsUGFaixcPV9CpOeE/8Rm1LBXX4NN813KcXSILSEAwdm38JizzOgp
5/vELkOZUaLBIyIX2WjJekSFXjJitP8W0HDpRc9i/kydEyY813AuaZy6wssY6NUX
QVNiOzt7L8F4CfUu9H7S4hAxgNvWlvemqJbUb+AcyLdI9yBqjhP3L7i7yuZTz+MA
l/mB+5dposIwPB81K6jz0e0qDEDz0L6pzFx4wmFqAHtr42cJBdK0g88ckmK/x7Hk
s/7bb3l0NlasWAPU/VhqyEEq2gy1HzOqvoWvAqfisuqf+sDrntCJmL+Nx3Ll1qD1
KW54Rldcv2GQBsXHnFn7nQuPlCV0/fMtmiI5N564nQk=
`protect END_PROTECTED
