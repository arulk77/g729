`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ9wVT+CMKrUW1Sq3tM22T0cPIdgIVTYFVTusWIw+Fyf
TPekw5JOsO96RVtSIlrEH6tWCHDttYg6j4DAcbzSsqiV/1ZVCxu52JzylTVsFfJ0
5U1jah5ZG+u1lLomXbwgxsV/awT5totAXFdz+5lYsj8uISLPJIYx30E29v96cKL+
h3V+XUTQCkqDxzp3J9cETCxm3ylB7GP3MMz3Vgrp/AN3J1TiOQiOKwkEweVdGHEN
`protect END_PROTECTED
