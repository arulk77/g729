`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4xGTMl8f68Ivd+IZTfjP3J2BJ5kFcbrw423GOZE/HfKbwxFRsfAe5hIjAm4x+8GV
WzKilqVTXldEpf5zwTkt0577nq0UYq6sBYzKwnITOH/4bJ/6d5+KJZM/v4kCQ724
qEQ/DTMvFjfXDIa8wPZCbG7mXoA59F7rYDNsjmoK3CrA06tF5XkqYxu4udGbXeC1
LHGYOXnfSVVwGbU9Sp1pRSEqOQAJcg075TSLKfDGIrO+t/IepP8O2PBeWpzZTw89
c8q959rbCNumA3CPQg9RBQF5ZIHsBVMuKUr/t91N3dnwsCCdlL+CsqWouGfbE0R1
hbVCB730mXw5NVADQXXPf9XFzn+dPSP/fcjeqB0Gd3WZFTXkBP4gggjjsPGRh72d
eGukkbrUDIxxzo7QbA81guG4vOvbzPgT95ciWpxbLMqvH6gnjqDhOKaQdRziiywM
hXEKuwqGjAlRLqMhxhvOCf5sQPlVDsctsybFx1vcq+2QCKcBTKxg1lroDv9oRMc0
vTnOopHpe2+bIRHxUElzQva5TOELssE/r0HdqjwgpB21psMJsLesugf20VVs6fUM
zpl27211cUQZroRPGWHFkCVz+8KpifXStGpXrQLRdO24WWPWb/5T6mQ+Pa5x5duP
jUHhe2Emqm1uRmidT8K1jfhHEyLDbCSht9l9K6yPDnRYmQZKg6kvDTHddEJZX/b4
AXT8DS+APw9ef2lq+DpnxLynXW/bxBDvepvRqF0wr+s=
`protect END_PROTECTED
