`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49vBKxykGmAD8jr8NHHOrEoNuCXYk0wUTH+NYPaQuTEO
LdLlaUnJ2bQCb2i44QZs8+E8R04Re5WW8ZTlDoNzDbO7g28J5bba0pZrdp+EhtHK
JzjIaQVpwUAD5pBGiVv8VCjAq4tJQnlDep71D0DcyorPFl4WazWbPAJr1GLcU03r
pfCs52yvEfTTxN5tFtUFKiR5D9FGI/1aIP3uWhcZSCA=
`protect END_PROTECTED
