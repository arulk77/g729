`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMWV7IjfbU5L6vsUN8xZyNZd3wFsF05/KHCn3Epbk/0O
UwX/jHRIf8qSf2Jh0OtT6oeyQgP8gH6MySkX2IUJqeX0fCjNwiFoDyus1s6SpbOi
OBt3qnKguLOcyZ9MunA3PI9e22MY/lo5DO23BneJB27NcRQkugLDyIIl59TJIDXa
HLF3PZhxySQxE2N01ndYZVQGQQuvyZ6eLngh1Eqg6bfZVTD30zfYvA3rnHm3lgeJ
hrVpD0osMwfaBUugMAJ+pUcKfOkTnevaDwi39PR/Z7ZW3FHeDnKweeeaDBXzLN0o
EnZEburjmct5MFVQ+p+QttbK6l2XiBjmwHr+8BxEnUfaM0NzmFpbFaVkPYL6fA7k
Z4QpVG21q3lIWMWTAhLJi4E7WZZNUijBMfkPDLjN/KnBvtZGsJyUUJPcveKKhiVt
vLneYi6Lg0QKx8jbCjWfTjx/0leQaS8lB4ojdOi0XhRDFR3j0FSfYHejrbvLl8Gn
YaD6n86/8dbxZoiXQ1OIylYUrv8wiUHM2+29yG7+kBriO3iC2QQTfi67WqR5FQZg
a/hhwKYjF4PcFw1gmkC7yg==
`protect END_PROTECTED
