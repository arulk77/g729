`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
CXDo269tkFVLssJhCUcbkYma5Det8vQYIRx+F7E1vj08lLFfsywRCPWQaqYnQFke
9fv+Q0uVtXMA0EMeVqgoiTzwgyS+uvtizzTX21uGe5OuU5KI9mCRfGTvRK4q87tn
i5M8Tp10kZIZd+tKZ7X2T/Yc9KiWHJ84t/OJEz3W9kB7FwVwrZWESh+0TmPQoRCT
`protect END_PROTECTED
