`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkWqCxUE6aRVJ/dpxCFlXzYPGivGORSfxN0gTsT+FB6EY
nKgVNOkDH/IfhBoP8s72+UtXwX3N1+LwcMmVEhoeQQcq2YUdVkI0fO6Fe1TSgLZx
vG9vW8QrcdbOfxMzn2m5un8KDtrKNYigCpOo7I6TdEzRN/MhorlH4r2UaPJAYJdp
bKHKNXPTsi/JzcBKflvFOI7Nf3T6nm0TUQBI7iGG0d+qW/RoooCR/hKcRjVWCwgr
lAmXLus/EekRlWwsYHtvNsp3vOheiXpNnUx7qjDLhujTuWlldxH80Gptj/S1VrB3
VBNwRf6UMTpm5EFVadBfCOdXipBdRusBL8+QTSVH+XojtZBJmUvzyaHqN2jfwXID
4DZpfeLWb1GBldzS8L5KVLCywIsEIIRiNHmsk91C4JI=
`protect END_PROTECTED
