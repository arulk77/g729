`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveORQ2uczDA3x74iwueyNJLRHz3NqmXFFUZFEzL8JVH2C
No28xZC38Ns4C9YFdlinFtx2YLb28IZy5sCa4u4J+g7XjdDPsG345U/90T1mxjrW
d3KW97bJP51uixuVSAstYMykWCRpNbOW9kmtb2S2TVHsAlbUkLf+GQyuguJNh1P/
G8GoLTmaS3d+P3O49vQUOHI+BUKV++efeMt8pQVmpou5n7w7m0m7nizUa0pnBtK8
q4kFCuujRRdYMzpflkwgh6H2RIGqCRy5Od/0cyETCQjxcnO84RN3Mb0r1GU0aQsk
jpIDsgiAkSz/COECGj2+TnvH+VOIc4PNbq1btsEWTEUU/9tGum9snCTY6SP3wk+q
nR44deLaBy7D9MmSOT8XcO0EsnfaqY7GC4zt925EIz38y7P+TQxvFOr/lx4XbALJ
5iK9xXbIqFGIv7kQkE2X0N+KOUw+dKH24sqUNP5JSJJNFlxLSeqs1gFINVUODDgq
Rx6wRKgoIVp+ka9Mnqy4PaIuACvTGxOJ4HOusi1ok6XVn9Fy3uWF/chIZfUm6Mfq
BGVtCw8v0VUlR1CZ32LnCy4n5S3kOuh5olJXX44vxWvNlRLPP5GwAg0y6s9hioog
jJIoHiDZVD+31ACnt3FUDJNoxcz4lJLV8iiFmWX4MBw=
`protect END_PROTECTED
