`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C4j+b/UTo3nQJsVymDcVF29b9ERxn63LnIKQqcVKFuKV
LdwVqQUh3k+7foCfI0qUSvwThNZFLDwx5dPp7eLVTmQlkUERzrbBswGe4VvLqUc4
ZkFjxpJO6jqz56JiNHOcW3owv/3Pu/sCWGwSL9GJR+eHOO8g6PS0xJx5Hs8OGsYE
odKCB8KdIjHPpIbVokqll/loQE21mRXV/427q0xd0itnN+zMVzcuTDtEnGru942o
dTtvjk+5XUX4Vm2K4t9mVBiegLqzKHba7OJ7Jq9oiYUqiC4Y39fZgADYUPGKDOoD
gpCDCP8SJTtU0Aw7lUA58bJwvX/lqTcPcAxw5+xx20WJDtsC/e7uq+uO7Mw92iBq
feo6UllA1WZ9cu5aO7Be0EcUw74lXcecbc8dcdD5v3C/JAxSEoVVuhWMCfm8QN85
oTCNmmUoeIbPGTumaOLSmwm0YTmOxJS1icUk+UDv1+ScRv02JwWVnQGX0K7D5CWd
P85wSXAY2/vQ0/m5LRH/bCXQ8yzDQXJWcPqf1OWJuDA1uUqspIJ+nXL0+Cvi41sd
aPJWt21V8HVV7/bsiTXBRrU+kD9kKGFCaw1oUUhTXC9fM55PWhcurKSBOMFp9y+F
MBknnxPZeFKS+ydeHGQ16hMv/xepO5fa1UkjRbePbi14/z6bSh4MNjdGcteor397
oPE3fNvZ7Xp3J0+wLityfamKazhOUQhzWwRafV2pHomsQ1nV+OKNW6mM+DQW7WdK
eHNnAZz/ShnrvrlMIXkn+e3u0KjfhCDf0aHLIjNDWvfmfwQirJNUenuZq75/oQn6
cTlCSM3Dfbe3SQDCJ2aTPzCUJWsHft6tdO3emCIJT84eEQUHYvkHWJwG9ofIt4bL
SPNuQbn8UMyXlf1ISTcKqVEdJJ0oWMEXMxyV+9B0q5vSTB9pYJXGcNj1R2zV+ddZ
JXZwr7spFMZekZWECdasj6BaiMfUDZnryPNgxN6Nd3elUuCfMHPGvr8QAW5GNzQ0
XLxQmPmpwVKu+MYE9bNKaaD6RY5YWkdOnW5BpQHRkiHwgBvXAhWuvYfVHHJghCwF
gDKnQYrZCXjSgFXCgBfEMh8hBIw0eltr3LL+VC/ek98o8n87lG8WF9BDnX3NiVTM
W3DVUHP5QtAwT8A9KwuiUuRgB5g1CBTnuXokIy78m0bTAlKRbHsG2gW8HJEjXhal
8C93oxBYyY+pLfw+ilU8IGugJBSO0SLsejQpFSa739qdkTa7uoCiFBr0F4xy2qHF
tZwfWDkNo2LlCV00MHDt3hoYJqIBWyd9HxHz6VRNzQCB5c2bzUZnsxJTBauYgUOJ
52z/MOPs/FebypVESkH0ddrS6DDhbNkqqtQ9Da0sBde3z7G2BGjngPOR9qsAK0pT
no/RNqZnUF9ZqclY3zgHd9OWAB7jN9umHah7CcpRLklB+FA60H12v57XvsOllcwY
7h+mQq39PTSeGIZYntwHc8N/sqaYVB4y/Ffo+4i2Qsb+e9mQjB4XTu1FqwCWnLon
Dc+rmQY4mJ5+f1LEdC/zd1qlEdHgvlUfOYM6eVZsnGclxL486k6GBboHPIOmrBrP
h+8hjKe/zy92ccSfZPxGkkhCYs4yrDZUUZIKHukzGptmSIH55hTyVJwQCWr9BJZ5
KPIR+poa1lGMZuMx+n1cESOb1xHRgGJgyj2EvRYIgUTnQbv3hYNB7R5Og1PA91yx
Pd796i9QCuxpB//tSg9XdyhGMrloXeHFHXcgkRJN/VNXHf+fTVKcy4ayHL1R9W3T
Mp26M5fh70GvCQiY9EjnxIC7EH4WNF5jcXmFBes73Tv9lVZluwVuE+DYdgOibsta
egwgPoLwQDqGT9ifR1/tgd3XDZA1ZiRu052XQow4f+oecMAd4DEM05gIRJnZR+66
skCEmMD5bjGMM+IoE+34kwhX7MEUUn22MHt1nQQJ6sxP7Nkul3tI8O2LFdryLAee
pJ4OAY8reAHFRxA+I9LTe0n2HDRXSjgA/As0aJQ6aZL97oJSIDlp91KpSUSX0EpV
tPYzayKbOi84EHVKP4j0e07GYqV7Ue0nucBLuia2HJA1wDgVL6rTgxlZGSbeUjK8
9/071PUDtUeVH1GESxnYCcswcNXuJopvOHcMzcF1A3DrBFiEA7Nq9wArboqwO/Kb
6Zv0b5Emvm4Bm2smW9qcRTjqdQn1PcG85+yaImWyswVtY8hThX5dq7zY6lSpnKw+
OrUxapx7ZCMwa6C3KEG+cw==
`protect END_PROTECTED
