`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
7RWERbz/SCu29vx1yp3KRKWXr8bOMlCok/fkkwkGET+7GGOgWIJy4n5SeEcAJfky
PFtmpVPJRRffHP82ftClbRHluqp+BW3KVHPDV0jCTQq+owlbBwQS3OSw6sdcR2jY
dV7N+rwszZ7EophOslYrrtUdwQI6cty/XYI3eXZcgJwugjiRb71WjKJCzwpPbgY9
`protect END_PROTECTED
