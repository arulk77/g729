`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu465p9rDooHYiRFkdTQBzzt9ErF+S3jdZPNm9AKUCNhpY
GxPMS+o0/Xob0R0o18MiLZ4psj6yG4mdiEPuuCOHFwEyiUQnb3TkRTBsKq4OumoC
sMJGvAoQ5sFCDr9qzNWuE5nFHf3Yyg6dnwAQbtoHXEvdSu2kEmgdB7k93W0wzsoI
zXzJ1O9xEZN1qyV8MKfAU3gi+wWRJ3TFgPJSuna/VIiO0ZMMgn4SjWBLMUwUbJ7Z
mJKsPd5k4CGy4vFAqllhaHEr9u8M1yAyW9MM7wRlT8IGQwTDyDHQn/18ARSkuTLU
nqweFAx98RCb0gmFMnAQE/X6Thc5P5z2LBDh2HQWn7Ls/tpNCdOFo7gUHpXk3Esy
ygJlXuruG9oVOIBtNe7BFxJcUc4wgAR7wPiq0jgkud+O41cDU1xBYI6Gz60T3OOk
3A44vf2EVqA4SRqmtI+TJseWCpFerqCYnJRCMF/jBk+kLBN0MNjYP1JtKFCsEmah
`protect END_PROTECTED
