`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHm1KLySC7p/9YTp96K/l3n7SvyMkm/p0zlDLZsj85Xp
hkTDnaU8Jtm+2ucruqVloFpK5JcJwdwlmqJI2yy7BEH963FGWuNnp6eolYSP2DFU
aEjGeqT/yhvPmCJFjIceyxdY0fF1XBKcHXUmELLN3gOgUUUTzNNQV9apxgSvzSWl
93VqZv5/g9k5JGZn2pOvXcXREfgueFDLy4b+DlWVh78G7F+uNBjIn+WtnH+iYG7b
TBLm/mvddQsZcbvrP6+/hs1wMaiRvpnHQuD7aL+Uy1bYg3LveVjBNdvtId2+zLAJ
5qcvOrhOx49bSbgAqUxvUF/ca68WdxxxhJqYQfTz6tl5trNEPISj23zh1mTjwDYw
`protect END_PROTECTED
