`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAWHwxcMUY4N0ixgj3KJ+rVwaYaoOlwixxkaZEc7GQnAP
E0v0gQomStlLQbOzGl/HxKq1/t/Sr01s6EkOdPZRaXI5osTKAwjjWrpgnBH3WneT
dEgFbSVktX0lPXy+CRyQg/pWxFc72fyn9fz3mjr9DHGEryAovE985C1Xmig02nQY
Xc0hdCPwLrT6ej9Hp6icbe/w5baQh584ugJZWKbYJ+wTp42PlK51B8y+rKuKC6bs
HaA5myM342PfitxUAQn1gcVehMPhMGKNTzhJZguKzeQhB9xgsIjhfELH8q1C0hj4
0EI4epRBF7GHuUb4fPzyketsuoLF2ugZOBbQ09iRZ8IsNysrmWQFbn9xkt0tT0Qx
o0sujJJXjyczwt7m/CUFnTDlZ74Z5DjWccTd1d8nJnLM2lX0YIywNeuZ+VrLmokW
GYBET0tQem57rdFvZ1xn+HGkW5o4DMHOUosQxjWkkFIenhinw0UdrBhgwXVjiKfg
PLQ7yq1PZHcSxHXTCrz3wsKbcFrLuEqIfagcFHjMYy4dRkGuHGNRHeHscXAJM71S
vih74GK+4MUQUOIIBPnBgd3S1Ej0V8fKMPn8fVDjCsg9AxMXhnvEhteOR7ax/5Tt
S6T+KRJCa32uGhnS5tVxwocGqhE6/51H/DrESuT704zuhfbyS9ieUC3x+BRl6qJI
MuI5EPrnqoJGbI/OuRzjIm4Tq9e883l4yN8TnNN1pAmnv1wkXtOlyqXr4N6ib6Bs
zd+qTRp/FOxsChaFWVDhxuK8uKN5Xhp4UkF61v7LZBZz4CelPRK3bMlxIr01/xsX
coZ7LOcVsm4FrUbQlqr6GqrV7oTsfWT9WM1VamTVdsIWi1grONM2IaZKZ96ycqW1
OdzeoT2Ca1vmXJwR4p1grEf0rAtc66JXP9kAWcJaLeEu629m6CO68z9XcHaEmaBc
75MppQaw6Wd1RN18Jj+oYjeoLgakMLorfXU9Swdj0DcomwIycot2I4G6+9dzu3Id
y48E46d+s4IohkoRz7SGv7OHURjL9OuvK2dNKhvRC5Rvd1Lg7WfwJgfWKpTwQIQ7
3K2Hl1ajIG6ahO03IIHvJhgaxo7z8J3wek/F/msCAjHgaM9Ew5nkkMHEaxOf8uXP
9h+LrOJvOd3v5aED58ff77onfC0jlyCi0/La937ycz9ZGLvfCvMUguGcyVznIaVj
Vf7fZgn3druzkY4QhAo4kHjTHtv34OmgGUuUSw8B0CavOi4sGVITJnuoGcrdjUUS
zkz1/AzS+J6y1S+lEy6RZkEziZjVZB+4fujhwDIlhMvRTQSo71OWs8bXvA9s8Mjs
+W/cmnoZM6Ukd3vvPL4OBTzngjV2ZWEXJeIjhLOnV0Mgcg3iumiGfAxrlzT1ZUiR
COsv0GFEbOxaW4UoSOobv9p4VJXJI3LzING0PVQmG9zl8erSP3ewB0HXPzB3EdwD
YN5uoOPr0qbzydkIjT30zvwwMwHMBWiKBUMtpAaDI0ZhY9RYXXiBZ3HHMig0N4vm
QWnQla6sb0JT9rAP2rn5A/CdjFbniwW3iWfUyok/UKgUwUeRLY7xk9KETgCU9uRp
I/e1PFfVRIzp0dJttMg+w6+MjvVOvNr8aenh+ooWQE8da2im42efIQYPneRhY9wG
oac+2KlDPJrqvl3MwTPF7uQRipwk4cqR0EKsUkQBSxYGB95y9EGhWZh44Ri/4hav
kHF8u8Cqxq0z0K3+TLWuVW1sk2jFr1wf0fVeRBnT5X/lAT23WdRljKsz3fQmTWtf
uG/iKExorQsfV5/T2cr75e0PeOClKem6rYz40m2wRVWB/Z6xD31X4pgckpnvFj08
ds96G+EVWzBVyeBRwbsX5tpBf0U41LpxUU+DmW6OJD6t1TkXPGQcbGJWmDTwvAVK
SDH9taWqbaaVSfuZ09k94XzvcWFoeLcOOy8BPMC/HXOCb0WCFxyTnz96Ssp0xIyV
sxOQHPR+pbyF29BTa7l+IpnsFfr91ImoPi8LGEFwNlSk2leIZBD9wrOBvzJMZNUx
LUQ9nJlsCCi5OppTBAhW+K2dpCeuOfnWKlO1kh/gNiI9eUsCG0oRFDTBHwgjsE3y
pLTt1H0g/FVl0VEkka+S9rhTgLZt+nrjr1u0hySfklaPwPgL+lp51qRuVQZqVdFC
gek7UneRINsGOotzRmpKfjNaQDRgEiEufOIaylOeqmPyryUnz4utGYh6CMaoG/X3
mWTKfcBy0Maz/TczVC9TNmkthkhMWEqOgh8sCWUaVfDIHdmRbWxIF5rMJckeTDY8
ojbYMqIID6ZyYrBp4nK1m4mY8M8oSd8oyb7koYail7ZZUATitrckqet/ewAmYRww
`protect END_PROTECTED
