`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePdMzGO7hwYfvg6ezQ+BV3gYfwq46eS6hRTlGGoUFR1n
20iJJSoXLsB9ZDEDJZzQDThnv4ApSo89UxrZn/TvLafT8muu2dIBIseBLqgs/wQU
sJuC6LCxu4dw08rf8SXT3YrNJOm0ZZgt+e8ghTR1XiHzhgc3TFy5RcD/xqpMcwku
tLIvz5yhMfYa6opu/H7bi2Ex0zPgqTeoXuhcQ/5JtzDzG6Cr0G/8J0WeP8fTYYqY
`protect END_PROTECTED
