`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNw+IJxuBveJ9iiFBsTAkXv80xjsfXxzjaavgG+QdZXFY
AV88NffbqtbTd4bi7hI0iCf+wSO88vLfY29KbXRU5LCKQwKgv8juLL/LG0epqc+c
OO4GWAGoVSLxGU9MtWjluKVJl3wKFl31SmFNdIOEoVFOuRASREK6TI3/ULwvmXLd
wtVqRlRMh49d3ETIVzd05LncIRi0MoZTZzrmW9N9eeVdezIlJJG1oXZ8dtaTZDZF
XxdZoeCrA7ww8N6iiDl/YInXcPQSouKf8Vet6A07Pm3ZkihsOcM1AyB0Bb6ViReH
R1NeHu3ulKYMJ0964dkm4VYJ3Z9FYrQ2+juOznZEkRp1l/LzoW4736FWeMPGH7z7
vIWvPJMdzxeJoLAs1z58vCEZ9pjYX4Lz9xK8/tLzu18jOdBasNHNxeER3Sh9G58z
qirA89CNX7zknKCfdIloF79ADydfm2ZPgK6fCyxwCnP0xQcoptoZ90tZlMcQlOX2
rZcJrNsDe7dQZNwG4lgFr61bd82AKMgzhi4Y7ksSp89tRVg1knAwEDPlJGS0nUB6
3rUAXmawtygq8dX1WKYV1xNhB9/cKWOi7xbhzxWpebpUtHDNJXhKtfx3Dvy4vpwv
4GQE1evQFZrkR8mwuykwFRhvo6rlhDFxrPQwFJVypvSB9oK9aLHnLe6eEhcAHL2R
21NmBGp71lx60GX5dQpArQmIvchbWb3L/I/m3SxwaClyYC+O25s5UW6/qy+v7n3t
bfWnjYKqLEkT6u49nbu4pUACYMqALKlePThgaqnTKQbU1vGXxMosVkBK8brQZZhS
yvYdloyYO63K10HjVWN0uC3ecTTVlpkle9Briza23OO16JS/jQ9KHW8UPH9A4t0l
XzIIVXYsw7AWDNZZLetCVjL4i09sSdPhtSUyD2oXHkk2zLku6c/YxQkxfaqDY7H5
NPB8DxWw/GDx5JQB3+mhj1Tkm661un55cCcPh5DqUZpAoqT/b846PRZvrPj9uj+g
A6KhEwDxrIvN01pst9s20uxTVL+8QQQRRVI+0pJ0r2hIWPrAtce+GLoLINqMEPN5
ERe1u3dl/sc4cNKNOdM7eQg4IxDGVPMC6a1VMyQs1PEv0rFNxKvzEEhnQbekTUUt
IqxJUvTjjTEf8FCaVP7S2w4IMg0iXQOexuE4+aeGNSs+miYmK/RDfp8OfMH35zWO
6FDhX5H0lV3jsuDkRkLJuo+bRZe4CSeY+wbAO0YwTt4tukOGYFDMSuKxn2zWGytx
wsVjBmQoOnohklTp8yawU1ZXVxkQ9BgUKElYhc6XpWzzxwePakbiV405+rqVdhm8
lh39bjmhOMcwMwLtHtdWLWjSJ7+NknPOF1ez7JoZn2DBPgcQg+hO4mZVjHjMqDgq
Syts9yffL0EYUUrmmHjHMvBlhdoXclH9c2BbjSQBcoSUyLSiDpYlHoDA+apI++5g
rjL78cLZMmzRA1KRsddCMSEEsOB9zL1epl4RKwOcQpcburF17uGSYD/tmVBoqEVn
rY4r84EyG2CqlsB/avB6ez54lf1YOtFAXKzcbSv6xWWAaPqrAISQ0gOPOLd0K4Lu
X98JXFTM54z9HnmrqVytuO3Nflp6nWmdIsuoJXbV0f65T4X8a7N5jl0m0pWl1Yse
IvcW2CXL3DtWeo+KqixV2Yjhci4Umr/dAAuxfD6N8fRCu8pWqvOQl5qRRKojcFwG
pas0POo2VbkX05y67xbwGlUFfjhUCwya2EnWJmtV44F/OBoA76unQ7eJPfEgrAAY
0zQvTiay5Z+bD74n8cM2lyxRQfU+x4eMBoAVHMpRi0dNFPP8zPFhs9RNU+0IFllH
UtkCNbfHj92mcGVHLzNEL+I8tfbLlv3LHSJv0280wQe0+HmerOqeYUyruOzKkBaC
n0rrvo389pPocSz1J01u8QvTTuuqiQakxwfhQWjxuSFlbPUE0c9ctQEiE6xJqP0I
dalwCBbC287MeqJKGnNUIiqPHp9AQkOtQ+yxkMXcafxr8CFHyHozLGVGx1D7YR4s
LIw1LIu68CuehCyXCwnGtdw2wyzAV4Qxv3K7hncsuceR+WSrJzmdSll93r84mh0q
rx7n42bMz2v8uNcBpr9V+8h1IHRM7oSJG2GTM+vnY7rF69QDjrsT9A/amy9rhIFF
By6cUug5M27+nTJ7mFooj1yGLy8m8lXbp5mfN8iri1lIgGDtuoP22rnpqj0tT30c
xy+d7/6tuLrkmqGy9AlSUZ7AEF9nX2nXMOLIrxJO8gZabb9L3kl+WfnVdR7+MYfS
GSTsFemFtsx5QbFNP8rDU7JKPtf0BN07WjFvx/W1xJ5AFfBPASmEq6jWhwxGl4v/
xuyC3LKG5NYzGCG8dsxmUCrS+v+GXM/1v90+K0Ll29qx7lvqmddIjT9A0HMSt/XR
cq3tYsvlFfMjazfToQLYtB51Omw5RYzdz/N7s6RXPHvYYXi8z/K/XOMkRlGzyNl4
wElhOIxA8P+Jp7WYcIZJrm7jiHp3jNnalRuXq5JGm9K6JCbrmOXk7kzGJOoJ3pA7
+bXFN90w5yZRE7IZlcb4QYk/xNTxJx730Wrg3COq0p+B5kvmft3jOdaLARDoamcH
FrZdka8P6XAhX33bmIoEF60jdCvFZDgTsSz4dSLBzGmldILD51ZFOpLlxHAVGQJj
A2S/Yp8zy8uaUI3V2QOJJxtIkRZNTKCp+ev34dr8x4wfe7iylo7dFYnNOc3Mwm4j
wybMArFArDzu5J/IzX7g1lnholivJKuvgh5cAn8ZQ2dL9QhAG+uf/cdppgE8vg09
/rCBgG9j+08bgOXpJ1nGRSn7PyEy5wilJURdNbiLtPTMKgGJ6bU0IL98MFjrjFab
0uijaktPySnJqxvZCV3qxRmzBTOlt1R5Ys0aJpsB6Pbj3gvcKRf20/At6lNOQ8R5
+0KIMGgzyEhh06xleIt4Utg1/nZ+NSNkwsq13HsVymtg+4rxTwVtcu3UP2QgOWcP
wgU/r0WN7ATgZWAcfw6Chr6jxT0Gu7ODXk/GGVQ8B8KO0JzOH0JYtxpDT58X0CXy
C5/SC3CAtCkb8bRrHIYrnezXWjt+SmhZkDYPDWA5Ab7N1VKK4fAveF+4NGu34/K/
GnCoyjxozIDgTJvQA/65dG8LeQ+BtbnUpMYKZ2c9D6NlWkA/vTJ1uxCkvNub0Cza
S4F4QQw5LXv5vbIxOEKFDLpwX0h5EaMvNOjFKe1Lrbq9MlnmsZJssmdnHpvawlkz
UVVGbjN5wvKpTU0N1lD+/1nAHW5yiWrykK3NpP/cReDlkAefwM3epYXQUSroIkJS
eCRjJpk6J6MUMB3rxQKAQabt88+nVFdQxGfs33OK0sUTyx1A3QbXenQdIuVujgfw
SZ75X/Ow9kNeVsreNwgdS1Z0dzobkpOR2uD5mxJvN5OdjDCSXUGM5Wmow+jQ4INh
1qVAw8ATadPDxsdO/AdzZEC46NKZvxC2B/UEfeOdozb8oe4sBGfOewba/d4vDFPn
TbKzZiL9jQ9TL1Y7u24i5kmn2mIHQMXM59sSJEvYTLZZJcYhyC19bq7xnPhhjeKr
8XTVvr1g1e9dcrfM9UUJAV1AC9NvCmuTLuLGFJ98phvBvyjhZbGN8+r6mojA3OSB
BcTv4RTtH+LprxB6VFmJ7xUBcQOzJmb3/7cuxhuC77ntMyV6AvcvJACsInI3FGCF
xzAEziYyzjG5VoSPPEaRTNsKsuUBHYbWN7HQOlGJvC8oke5Y8zHaRmfRT0C34hV7
YxtONuiCf7uEOyvqdQ801EE6yWZQofR3y1J7ELoV36olPO135jIsDQ9fJX3sbT+u
IVK57FA45vt2am8RitQqql3GW5RIEAOYaPiJ2gkesI3YYGe+BHZaX7yutXtT7z2x
TvkvhKtWPpV6hhoVj4KvnJu93hh5wi8AwmUwNzocSmlzDLzw+3hQbc1v+fcwEa85
MI7cW87JAm8c1P0UuqC0kZ3kpHfaGPnesOL9zxXuBX79BBwr0fvUST6SP4ZfYaNi
0lnCd5BE6Snmoxl1ge4EWcTLhRqC8Lspq4zsqB4yukzcpzCMFNaPB0zEq19s5DGB
yXVFcMR7XfIJaX+msj3WvsL2Upl5zxdWMbm2Oz29zNuZO5dSCNFHEwEFOSP8nVaH
F+Qrwmz7vwBenjLuwLdaTkkpe37CF1rZSR565gLOa10HO65oZ3st4wZdonYtEEXl
tGCYucOPmvjmRlThlzMDQ8Z3j2mEBnK9XW8zJE+xrKuDBueu87w8gZKa36w1y6bb
2ZDgATuQeOsJQ72ST73ECenXdNtAu+Dybcv4G9o9AeEtBlOIvV6NWlHvlio4ikVV
c/GUFQCyhPuHEF8cj4EI1ovZq6hXScF5ZLGTYQHaJXB0PlfXPcl+IdU8wcWCCJVv
xGS1SkiIMVDeY8g8nPaxkRiFe0Wo+A6o0aN/mLy/UYhzITpHpiI0uCOVekHomW6P
kZl7wuNsjZlQrsb3ZpxXr6LOelGipa7TVFjdf0NYvGD0PfWTMnq5PKp+dOf39L/2
yQe89p+SH+o1KspN5ANvtnHHyG4KpqtjmQSx/8fS4WgKsWtTeAZCaMNaYRP257PD
xsPocAAtfraViDDknFIm0P15PK/u9aqaPXDJ965K5edgR/ZH8I2nqNt9lRA6ZnaZ
8foziRxzPZ0pDeIsG+q79/8GRdDJeug8F3zLDp+sxYcwOVHCCQ8zeoxuK+TGxwrg
P82ne8rknX3ZBXQ8/lhHLThQ6TkodCd8aZ0aGP+tGxd2Seg8EtmFjLAbbVIEgirP
YyIJvHSsRjiVysIdM7WuWYJNqD+jySf/H87SnGhXJ8gNExyaW0G9D8uNPIly0k9Q
UcVlua7fZqOlp2dBIBDhOp+K9g6OIcVulhSGS9vaBKC407LYeroBbQ/sWmpey/qT
TXJWWGfNHwIW+jBWLQtQ65/jse+IP06ZV1g3/sROi3X/DSZmdKigyQ5yvPRKSU82
3reeqT40m/7j4s2c/d4gvRpLx8l/dV6ue3OORdLcZ0GpxDqVFULAEdrdsWs5ccsZ
D6CyC9NxFsWRS3cTAKKvQqSuOJCxkoCmW1Nz5HFqz0mckdvY3ze7OhGoaCeZdz4U
s+5ZQMsJr7GrHYonnHAvE/qyw24VxnDmY0ryrsZE1q5HAeDEThj65k5uKU2byuaa
4vQVkjFS21UCZOTGDDOUQ5TeVt2P8TJP2J3sVnnXdzzHfaacU20m2qwE8VYCFpKj
3f0naaFXQDf5cx51ok6Uagn9p91+Fo6U5UOyugK71LztY+CHXMAZmnhMNCM1a3eC
KR5LAHhUyCEkZ7OoQHzeWvbWGNDaLeKps76tYrkS4IdunXCLonY3FaWr/y3nLTqN
pDq34i49/1gjdGE+J/SnY2VEsTfIIdqob2S0CGMQjT9kg+KtTldCocgFqUgrlXqU
3KAWQwHdwDUGaba61+GtIWS5Nwz2nNd/jMREyvTVWRBq58IOsOlMkr+KsXjUqJz4
L8lXXg/N13QYm5SnS+XK4nJJ6cn8IpBnd1WIzfwylYY7cWpG8YD5ocLRNNqvYKyd
LmMG1xC/yNeey8xr5QVvsDA2AB5gcMAxt3zkdum1ZdW6s4niGvxrVPCE9qkVM30K
2LNd/aNp0yKnS5BDY0RcOKBbt2y5Ma4UaUda7EtiBhNEtGj7Ev74VSOkFH94kNvj
ttaOiIsScXY+LLZvgs3KG2Jr36yR+WwA4gdxw0N0W+lFTwQTaezx+9F3ZzkkGpX2
Xuvu6do/UwoCmyWXx58w04siMpNvVJlxF3D57NosFTCbdZ3wxDi9KYcypZs6dQ/c
/N1D4yBzMdesjAVx3E/R1qO32q8NR6WG75jOTQse5e6AcgXQK7zN10uaNWNyj4Dz
ATlZ94cf4UaiQcTM3re/iiFctkW+2yiIGPAPFotPpss4V5zsxNskxQg1RyKPOJOj
/fjjP5vDY14l4jEpWLuExIiSsiyiV66mVWKt5aYF98w1/XVGaQDDcGN215QpinHt
NCYa2S6R7st2FM/tov1+SMfNAl2n5sPAlrXHw4irRStXlShHMCUTbzQ5HA//ROoT
YbbvCkviyabzEDgVYqDBRbSd3OYOioHYoXYEwTZDeVbxosUqvaiYBltPQBJu9KEs
8M8a2FHqxEPzHFoj6RBnc1Y0l6OIRPUfcQ6rlYN4CElc8gBmo6ZQOsaTvgT1Gpy+
zeUABjCaXPpEL1YGajyrH6XK4WVgM3fom4I1DU0ppP1ONbzqumR9fIs7Am8K4XKF
OUoAUGwtx2ituGewIYCSVIpBw3SGfLXhHjCcnPx0pDokW69hRgXRHYkD6bKsHVvZ
OeffX5fEL5EF9r4csReBUpiwY2XliXJjG0FMIbEDhu8JG7BKgtLiI10sGIsQfV0o
45aRf85LcvxKo8UBGn/yQJL+WwwBoIvOjdouE8VNq42DFbl/sap+H4KN4ubD0tcE
13GPv81y6bJVwa46hT/l3o/ttopZYb5Vynsurz0Dqn0JCY6GoEE1WqtZR9EwUazK
gnikIYaKReJFXRY2ujjpbHoYi1/Ar9OTSNxhsqrlZLToYNcD503c9ZNwi6q4gzfh
/eKupaOLYVDTt3d0wjIGEFpx7nKYgQmJsTQW8nPZhoL9aBihHQy29biNkEbuqr8S
9poobX4pQFkzoXsqMza2a4lS1r+qADZ2b558tECo3V0Fm8RhXbwRZK9ULR9hB3Hn
peAFjTQR5T18j8o4EutekX2nmHBx+3+rlQTzNfT9ZVVU3zOYQH8c4KDert0EyOXV
OYIa66eLEYm73k1kv7Y6nnlRHfaNgsFiuIVtGQrcv4gTwo/9St654qDUFb/P5Io8
BErSORNwlpokiVjbhgefKhnxe/W+MyKSgDm5yV/FfSFIrJ8bg7MBuPUbj63Zd3Qa
5pgVbhs9mCCUhRNTEl0eUscPg0Qi+Wbk4O+uAEmfRm8CaHvmvxbeJsJtkQiMRYLS
LlTWZKGxkHtbJhmwXJo4HKbzhDMzZbyQL//JmDE+PZL7C6ZLILoo7QbS3ilVi7TL
I0wzhanAh8BebSTkGFGLoJ2FEEA5nIu/w3qFsnfq7Og4LcpIKytnP/46FF30ZZ80
bg+iqN1Wfojr8XPWW5H9qi9KbQtAH01sdHr9RcV5VFze3N4V+X4jaosOdn4PxY/R
TZjT1Nkagj1IszmAEo0rtLWVloo3AYYLIDbg/FmbiD9V7oez4NSP5KhifhzZJTpD
xJvBB3wiSsRCPRLHB39McUtcW1z7VTEu4BDdQQGsgmsuD7OexOWSZyk4WyDHWP4d
gVxE5uOfXMsuMNvcHDNcNex3GzrhRRke8tCEyz12a9H6QGSXOpYAxb+Z75VLzBlz
1j7uaGnt4n0I8/US88VhHHf472MaK0FFHJucvzGL2iah38P+luivAJUF0dLY185g
9zpwBqJW6mEDWLnPCWmdSkPCmzjFc9ZDiU8j1uaPYGovdKvnbCuLVocQ9jBNeCFj
+2EMLBYg7s+ihCUSH3JSMB4akZkqbxlLCSJ2KXzrNtMWSZTzv/w1w369OlkmJinp
+vKgkfMw4dwQYQ7TJ8OH7Bhe2cbEpgpXTejHItmI7OQZ9Ttv2FHUVg+2mi/0Vj/I
MVkSn4VNm2jGJlqqpBrYBVxpQGt3dYmavoUEncgc8fawECUlPrxaDvlD6Z1qYrSP
0T7iY7tlC+8VehzOlctdHk+t3VTxZd5swmcOereArXu4/ahrgWDaytF9uRvmD81A
BjMFCr76qJjFGQ5LkusnT3sKrxUuPG/xYQJyZFq1zTZNFBMWou1jUzxbH64i5rhk
aYTlKe4/espUeQOPYP5Z/W9oBVkhwXucoIr4Jn/x5uyxW79W3jMLLYizzdblWYD2
PlZ/Sb8Rcoqp0Z/QSp2hLecqfav6yuTvAI5bbiNT5eE6J9BmzLpgs5EViWJxwr1G
1IgDJDn6oG4wv/lySLqdZGFwBiOUWJ34kVxbMUh3r3tYoZemI9oV/KE/EItlVRUh
LNgorHJbq4DlJMKuOniNnrphwA4JWhz8UX5zGunPW/kmwRdwlTptF8rKqlTx7URQ
ueHdT5xRMep4AT+h6rDifWwVSb5f9/YsvH0v3TFn5SimkHLhFFW0a1QIyMmQW+Wj
k9p6E3aHqlWMDKb5Cxqal4qbV1qD8aBo2jqewDtB1u/Ef63hAgMeCXagYtDPOEUL
6sXiOhJD/mYhzqPoZtJ3SuWAelR+KF7vMPApggKjB/JqArYRyQDnb2UvooZnjkpN
A1NzIoD0+Zey6XdpYD9bSaf1yNPjE2NDEqXkgtwfzv9h4tzDWcVvyqCora0cd7Da
e2y+R9f9G5RKg5KRoUwN/bmCOigpf9Nr7/qEYqW/wREiHxv1nTzFeSDQJRDSVh3Z
Y6mLjHnpzi6rLIuMFfnYDJwqbmTz1GASUvxwdEFF/B7S5UZHex6glRJqgSyQfAY/
SEUFJhZY/E2MJMN6ZE0shRuweXYHA6+Kx+uVBzZRKRMelegWJjXGr0uZFJMVhqhV
7morr9hDFLTmX0VW7LR+ks+9s5CV2DBDyuSTauUtwBl35n9aOtsJhys/K9jLowO6
rCXv65IDOuU4GnektVt7U4b5YUkN8NXgEgNFe1AWx2q2nVfxwddh3VpN7FHaiKZw
PxEyIXmWNDmtTm467i54yAUtXRTtbkEcPnQqYSOWepOspUuDgC3vba7rOno/a5Zb
FGh6KrALU3g2rKVHbjci9d2lh5AJxg/1FWfZKvgvSYN711eGGN6uterqJTNS9SO3
T8vN80WITbPSBFJid3TsvChfqaIbZv5cZJR85hwrNcDcwLaLPF2w5EAGdcp56mFJ
UNtewyYgK2MNBWLld1m5karLkicIP4wgh93u0PwrAR/6LGrC1PM4tkZmTEURNh1F
mpEeSf0TgS+CetxEJ90Jyjtys237XNB8RjR7BBEof0pHyzEEcBzeaBMc0auMfgdo
AaD0icnlfHxQ35ezPtYmPEvKgjbgtObMkrd/K56gwANpxaLcGj9zLx1j1mprMBDP
Bmljkj5vT6cjQG9/kzLGjy7Z9qOUlXcLdq0jgbSJc7Jhk8E/6gZXaM1d2RNIhv4o
9aMswyHvv2PN4TnOYuitj2tADxQT5x6AOLTmYikYXTqWekCmZBrAsjPL9e1pePXt
b+Mh2NjpVTx0+8q4I6fa+/LMSRL4VNXO5tLLK1rPBSH157T47vvsyqUh2f8UA7EW
0tRdSckNKG4XlAljmn0wcKBm8HiijKhbTlokPhAMisGcAwpPlfbEDre8nvPq6cot
ZFEIc92JriuM+lLdNj9ZZE7lNAaccHGctQYJkpbHT339HAibF8xD5lcMWNhMmPq+
yu/hO2mo85TyrOyADilPegEVKuFofZeCdVNdKlC/3LuLMvr3OU0jkPgHnpeZmSu0
KPZ5LH2iUeC5PzRfIDUozUekub5yvBbRLu8j7GBdKBGu6ti6q+X9/wZCrhKkeBqI
jPBNfY/Ldr2R7ekN3BMFn3a5Tj9z6VMiLoVMtv21RU8IcsNUYKkwxeH5acaLIeUl
mhfI24MqOOn/JNkltGN4+C21mhnTizz4bp/1OI8TKmW6sZ+6AMT/JFCWPpa4pnng
KiktvitfLSr15qEJcmKDDzb174pZWguaTnDis2DTwaMptKA4766Q5S5IYp7/WLQ7
HIzuIJDzeQ48Hs0QNVx3sKapoS5s+2T7Vokr4ibJTf9+/Wv6DYPKkOwN7Syq35d2
ZLVSPqBfuTsuUGTkcapuiH8vFPzsfVbVRl+Zuiqtmr9Qy9u/VVUuI/bxjwB4etma
Y+44Lol0FNrhyOG8VhSVIjAkNWap6Mt7J8iarJSsp3TvZ7xN35IODGjXCWYK9qQH
G0nslWU4lDD0ClF+wW2UsgxOYFDNqWVlOiUqumAYSa05jos7Ih5tvDzAObCo8qAd
BSL2TFQSL/rztMjUUuFEl6GOTyzEqparfT8EE1q2CzKKjEEPsFN5tbSFuV2MweaS
8wSBOgks2UKDFVeDGxJwcjMvbv20Qamk2hdyRVVCGO+Tw+HiCYTuwriyc9HIk48Z
xf5RBQLou0JYTOg2+Amz7CFx0XUh2N7bkoDNoe7fVTS/Rl1fxk0zZ9usCijDj/ex
2JmqKRnt+1U+e1DIgixjUizp5dWUPhmcpNmxMXd6aT2jOhjDIP/kv0zMOFi9ggrV
x0cVTT+Lpty/8epS4F6bSk28XycwC0ziZQxTkwwfVTvSS2S1AAYfCUxVTSdzP+Nr
6jgazU4v0OXynvNw9AQlnk6aeGpR75EdbO/ow6T2XcS05q5u+VXrWrxFx9WFBhxa
l4n4IPsbQrIWViQtmBY9BRZMrEUWY1KbhZ1tU5w3iLyB4SP/pCA9OZZPIQHhfoDq
7mX5aXkRFvLMbso0ewwF5I77ghWfwc13XT+SYSWXnUkrYRNXk4AJWeICJxzRIlQd
cNoUnKaMmA1hlPcSV4zCKEw1HGY8jZm7vPG8cqER7BO3fRBa0e+SGWPl7YBXDMBT
c0gD1SvENHYztCcmo9tYSy0BFEAOKmJzY0CDPTQh7YIjL13p5mLlJIPT3tuHCZzx
Ug0HZHbE9ERXfYr9+mrVP4e/xetb6PuRh/6lbo17iLRYgrpu08eF7qaE1KfbanUt
yCx3LuR7Wc8Z3fFG7Ch8dhFnmSLtGehi93BPNxpP6r+di/txFAsj9//x6qMoT8zz
anIKmRm1BHOHNL44YKXqD9tNcNLx54vFNWcQh7/zZk5pBo9KaDLnbJSEDDoedlw2
rXoemGvziRsqA76ClkALQ4ZTDZYyyDe4QzVA+kPuvKpV0v5rV2YnjXt2mboysu/c
lunfwcY97aL+9YqxXkjob6doz3OezQsVR4O1tuU/FdI2+QkpKlNlrL8XSXvRQMF6
vIVWiv5y0TvTlgjJeBYr6iNxsRx5QQBbqC6zCEVZ35+yw1Nb1flnHZ7F1cqTK8UN
kSR8VwIPdp+oQH46caONVFOqkjrNOAXhNEKm2a5nVarkMxZTk5axpNVCjND+5SJ2
WmmNaZPeUWUTQ/8q0nbSxPQCzvlGcUgk8IrMcs4kHp9y1z6XsPcGNQrGxvLrZm4w
cAViHHmk6jkp85abHNt2zUhVXFz20Sy1RZw5lnEeU6HsRnlpTDpfnnhLQwZqSkqs
EDArm5YiYKcSp20T3ufb1qkjGqxn5CgvRGRMkA+f/koz5nyIWsjRpc4tdJL6HIfJ
da8KUJZkaQgMe3RhVCk1CbjKoAvjzalXFQ65TvE6ffwk+SQAogRuEpkCeiMHcWSD
NnmXCNvsUerRa4eXntIEyWoeChF+7l8tBsm/HWA/QVm03FYerBNQdo9NjcICC3AG
vXp823S6lC38E0E2j6hKDcUyMFUUY3OQKh6KLiR2awMHOiC7hEbxzdYR9W28awcc
/kpdVSBx8TgPDpqxrQhJZ8aihGoaDEn5RHcofrwCqhXFgEHLvgdV7gMl3QQi7ItG
vaQ/i53mlWQTPgt6Pk8cdDmQynEH7fu/2KmeQuuoim9tzmW9AVC331Mou3+cIiec
2R8/WMiKLe+HKCLWYbcFFp3I1I0HUinkWnbJDH1dkgy49QT7W267ZqwJML4DJUmr
7iq47f7ThLDsqVmSlSm2DdyaO8Xdxd13FJiJ6CydQqVEYCl5qMtdm1qtwdfZsR7m
hF9g+QhfrFnEOl45Q5x3qGDxl3ww6071twKwFpTW0X2aGy2Ap8iIJKT67Sq8cFKl
rV3/RwixL+CnFyPw4sKK2vSQUVKOns6M7Y5wUumZfyX/LMK3DStBGziX/tljm+Y8
nNFw1aJ2kHdqixn19AzfcHLnjT4oFK7ojB55cU5z4lQ+p6A0YPamU9r2/kPlq9So
gCHkG9xSNPpo0Qgim1p3uwtCNVlIOanyszMlmgNdOMo2gUNYzd8B9rPe/PaFdptL
IKurO1IBS8n3Vd4DFRCAGAm43TA9W8E137nc/zYGQLBlxvlxPDk06KM0gN2l33OO
V1mupyIBEI3+fN9yYkQ8i7hLH+phpYXk4Y7JFstGx9aWViuAw9qGIWplbacKlej2
Hk3GecWJkRZhhgoLtnCePFN7bYb/WH/HKL0OZAAzWtLD7e/0POpBm5A5nqqhS/C4
Oz3e+8frBYw0N8Nir1HA39qjh+DdFG5NSbFfu++pvL7h5Gs+iIcRNO1hPITHbJ61
49HC5H/Jbrnxdz+RXnlUj99iXWdG7PT3mr+h+1Aj3i3Hgl01ZDNEC0xCswysMiDp
l6BG7N6YFReLyOAsH7IMJ7YzEOSzBb4L9vnOxd+g4qg6d2H3vqXv89JdEBYhOGIl
pBIL2Csqk5lw6Q/VtcVCx6U4LWnsxMo0ELTEsCcVOOtwJwVu97ZFZzUpQjoRKvVh
RMPkvNTr/HAkLCuYO0/tluXRQ9OUD/OCwmvChbSlG14lu6AUIWyHA0JIn+3frtjE
Qemjin4GWlP2xntt3kCauuIqvWokg1BKHiUtXrXXFqoEkrLbIbyc/wZn/LOVzyGF
7QJAf+MfOfKVtNVYak6qUZTld0NTZWlmQYmDAmFb6VcUFzaapFAR5hpUwGPxYl6e
U9yphPcY+g8hyxAbiPUTcotTOZhhAmRelwhgsTLNNJOj5Z9TAnNwTw81jF7MQZ5a
s08WIe1RLuPlKM4U/giFdFV+zvwpL8/LTt+BRUazKdjHTDCGnCX0NUmo4Kr5bR+R
i2KC5ZFwpUiGs+0uVVGtVsf4kzdupiRtn83t0RjexzcUL8XFniDaTW2Pd/emxndj
t700rwjEyDHy8WWC3iynKAMZPB35DG7xI8+aU9tc40cSBllAUHneMnSf3iwOMrF1
+1fPn56W9ivT7nKsR1/6l5ugrpdP4urBmnsBTOm3XdiuOddnKkKlShLlQH79r/oN
6foyJkXBxQOFKz1eUcTLZ/lMeFPWsuufIJ+DKfTPsrrm1QjVbaGyAMxX+r0aXCOI
K+8eWU37dumY1uodCoXo2h+sHFysmsSrMi01qzul+E4FqUpb3qs3uPva+eWa5VBp
L2gltLM3tsgcpVOVGxoq1sXze61hvEVJJOheOas2BI7EWcgwZ9Rmd9ev+VwdaCVu
d+MBFmywy/eCuJ7ARnW7DMK96O+AsGeFpJyqjuBhb8WV+LlbU2bgj26NBc3NOcxZ
ue6cA3S4TMqVSONvtJznPaX7DGkPIrLGrjP+1b/SQGJcmnaG1pd9P5JL4WP1+m6d
7PTD/oTpBvTOh8QMUMocP/2wgY1KIog/zM5MzFbnp0A6t6u2jl0qPIIhtjE1Unx2
jD5prXUapadXuqDLYyk8SB2cT681dpUX9ljU5MPhw6k0NsivXiYJG4XXJZF6jkB+
o9Mv/9Fmog9tUOPiYwLcCaHLWd+FNIw05mDdxYrwVTqZoMcVxlTguiOzhPsu54SB
pHVNI8cBoUU8cmjpkrX1IqUqpn30PqD1zNybWGNajgGJgDmZX35HIiQzyr6waoUl
4LB/f2JBRW61/gbG222om/ZsMZl5seaO0gpI6UcMuSCDLP1nETpdfa3aPH4cCRjt
DBZMRcCA7XRrzWzSLWbM1EB2hXN95l3uEUjNjepESqRnggFNQuFGrDpbbD6aEKVU
rhNFzO1F79TpyPO+y7qRqCRyY454zDJ8IeRJ2YC1gZUCiCCSFmjP0M7tKZri5AYk
AnEfMGLzW99hFv7j2/zCnYx2m8id1DBusyAsqOFLQ17ixH2Odp6zIcnj0MSv8tOG
CGB3i6CfVQFL81kJ8LVnjYUyK20R8RJTvIvcwdVG+6BgFaWbqiEDUJ9kBiiFgUGv
frPIPYH0IR53/H0dx3MrG6+DYb2dIz0IEEhhvCtwUV/LtD+82dlw6W/MFeYMkVvs
CWQ15CHLaUL5by95Vp95nXbClgM7RW3QVcfYuye1CQuvZcTQGh0vn2RA71yETf8D
78iOnNwMP5W0JSANKnu0MPp1CDJkpWA/IxvG4YaXXMx2fSkT+m/goCdjsV4nL8cm
+CddcLvP/yUsHUidtKo/41Sv7VYgAJdb+HtGa4jaCoimoMVm7Pn04ORBt3zDOrmY
cEnnaIYofVDKcagotxyH5Mqz8B/NPBzKitGDpTp8k1eL9eLS46qYanBezEfyuWla
CA3O9A2WojmtafOMgivFmsa90CJQh5+OWIoIfBkC1xEMTeA+0hV0oNcFNmO062i1
BeFS0evLLB5kn2kqw3Cj2ga4DwMWIU+vShhqXXrazGqKCetMXknLwWIxyu1ad2vk
fmQIZYB1W7taO9vHhuAByG2qMwC8mSNAnsaHjv8RkelXuB5gOO3nw+6iljfRdCRh
KdPxb0beFmZJ9rLWxdt4r+uCZNxRD0veTjfQ3V7u0AQkW6sv/mwRdW/t8Zl42Pd+
ZBuMUFu1IsE6EAPJ9MVP/+VM1v/syJApfacF8+qBkAacaUjYDDrNTQWb+R1k4EAs
d/zoImez7XINiWVKT0x1etWdWn+3Yu+KrKQSihXZEKEaFT+lCERGCW2+VPuQtdtj
j8jjacN5y7JM9Pgmji6ixeyUH+/Xo3P6q4xlaOCR87COlFthOAHAZsDq5oHtL0w6
4p2/oWLGainRluXxl2AFud5y8ME8wr9Vw8JQ40WGXvEKxbFqjftqK2U9X3DXVrPX
0vjASS/XkZXSn7y9nxbzhnz0bzDwhBGS9hS3OtXUlwhLlBscvemJ49m2A6SNU6I9
umNrouWEEsbthPXXwAg8+TCRr78L6xLoJ+n0CfxmrgXgs1PXtFSLeR5ovASdlZaP
b4TxczExlcx+TpGuf1R5Vr7sGhO1/eXvEQRudUioqe9USDIrID/Mr36mXiOrV4EJ
20FsJS//TB+VQVmTcq5ew3DMjZVg+/KBNs+SX+pF7ngIc7wUhbw0+fZo84HDOI/Q
l8YdGgPzxn3hmYCu+D1s1e6oJE4uYZbk6gCLvmoActsBA+fbA7Yvgp4e/IdxlWXV
COonvIFoTx2B2esXE5JdHackzZc0tmvBSgyV+25HOLS1/xxHsyDDVMmr/VKIoJ5Z
QyIvTGMCGaHae0sq1d9CU+SDwpFV9UwwatL/Ube1AbzAXdLwjMCGPIHBuAcffbqr
Xtc4Rd8mwAFp6sOkDts+d59wk9Opi3Lz9aMrC8gE8QxAaQE5EsHb+6XfU78Mk33C
d6Eo30k64YyQOeE9W2u2vGB/BMvP/QderYEIMFnBj7IFbhWbYK/K6UpzBOYJQuPh
qdfzTVf3saE0zauWedr8zedBVH67SsDEBMK7OfkyURIZWk+o9lRLuNoI++couyLQ
ILbh/LEJupFfQBitsBqw37mCRVJQiW0iecIdiYxygbs2cOITiMI7FDe3nTJZ0DMX
E/8hdY9S/ItbPIjCzr56wJ1/3q82nftfagn92Oc4d0Oue9DMNbX/Xh8FlqKuUPrY
wH9p3CcrN5/88ExL3fjCXysX5js5Wy3w4MPQEeDrGwc25h3vBFZ34zDSq+9A8VfP
zFUcMaGuUMK/dgiyqGL3Vre/p+b3aI6yyOP7I/Nx0M6VvTfnG3m7GW1Qs/olZaQQ
CWvU8H5MYbEkf/fry4Lh61X8TlGMYdoAW5GzTu9u20I4MAbKcSCE+dRGAiAAB23l
owOBMBVqivCKxJQyoK60/WiHHZAWrcE5UrcKPDnH4CcyPLyhWZFwQgf88HD5nT5e
jitChGMPoN5B4DYDSIfDGsStITzvIOrS0dM0pMvSfVCUmrLs1FTZDGl976OVu/VZ
m2lCIkk9MBpGuEHTj8ekDAP1EGLDNCohxViaEf0DQQGqKKRb6mPOMTig+4Dm3kAM
9EJk35XxoL6G7kg0RINo+oaQbhjDnL6a/HT6Yqmi7Oh5tipx/fjruunBYhq8B57x
+EEl9oM5tBI9DU1enE58Y3IYzyI3L3CLuBOOtgpEpiyj3ilZSZ1WYYegW25glrCz
Rb8Id0Z6PM2esBA5IrYFFOm1liYWbbygc3PkMpc/cevslgy5dLOYqV4GJFbTY8Tr
kqdKz92g5QYyH1zn8O35bntNIDeg6iS2igD0fpcMzeFe0J73VQ16H+5ebFNnYU6D
Ij7wrKBooQ6A9FYx22/+TJjqQd0S/Kf8diyLTy7OiqT//n7mahJozo80bTadgVUB
zKsqWwTt+EyegA9RPxADz5kpfowcVwrR51Jly/qWfmeSexPYRSkJKBE94uc3+VHv
41W8PlqMXvH6dZL9hqDOYXe2ph1yeM+1RBsGScHfJria/spQmZRxfLKtXiqC2YJp
YOhvzWO8yfEVFL52UA9mzT4MKDBERxB0nsK/Qvn9ZRJRcbKuyF81f25ryFg1vq6f
BRSyPJOyuI3h+/N2pj2RgOA/VCAqrDIkC5qgCul0RXM5Dl9xax5/1ULogktN81E/
RqnHkzNlzZOPabZXusrAVi79LfKtKVJdIAE0OwQsghKphSv/7hXIyDXKMwsV99bf
Ve3agQHRBQIyLGMzlgittKx/QP/jcXdsdFYCMVklUnr6/DGMBzlH9zXKJVkBfyhA
3oKQIVy3ypN9ZyA9QqVaGj+af1VK49FyP2VuLlVDvXCvXw4d0p6AY5o78GrReQc+
qMJkceFId7H+fg1cDx/AvPK2cwGk98PeC/zOnyORZyH9L/bgwn6m35e8lEFh3/B+
3qcgmHJIoriflp9MohOxvaNLmUKonfwBZ7w4lqgx1uvf1oJ3xEvkwyF/mZW73Jtw
0vZ0FJnx0STSr+U7Me07wHK5MeoJjARtuqyQHpKdbTLUb34PArxbhhyir68x4E8l
ous7E7tFdGT2yfeQlGbRWgE1jqOKVxcJg4oBwZKdQ+AexEig8H+cAQl2p/zFHH6r
jVSideGydVWkJKsxuI1ywSMAZDOrKbtya77EDEJGA0Cp1NqX6M9RV4kYxrdYmgS9
wlCvga6r8nsubpKC0bH/vA3faMa5NJ9FSky0QC5IeNYdH+8T5ELLuVK15mpcBWoz
rNij+mlm4xE9ng/aSUYtBEUGvU7W5cvPPmLtN7kFWg4j+NmcVNV5c7izZWGpHHZY
R3PwKoe14uW6iSC5qV8cY4MjeVtNchtuDnhTnPLrZWAyQ+jkvDgM9RY8LsHje2yj
s6nlwGHGoe6j+mqCVhGEfnk87RBqEpYwMJNoqXHluatSzX4xY7Tcw2b3n/pdSl1P
O4SidbWt3vO0ort4ELBGLPzMlW9fwdTl6bguVmT5VrF2fvlrCWaUSbOTIxD9yrjG
lBIUWko1mYQee9tiTSOyy+odqNmmogQtSeXrk2Z+HoPAzpEjuADAqima1PBS7Kiq
KwMuwWOUWgVAuxEN4Gi3vuubHVI1wLICt0+IUDN84ZvgzlcwtzP6UnyCyLyzuzql
kvRETiWLOFqo823GYPNF7Fi+FjtamGyWwoRezghVDch56g0zgolJXyTPeQguc4DN
6S7L1PyFZGi5SJP5jfJv+FsTXzF1FIe6A9sCZWqxEsk5Q0h/kGr+A+ENmQIMpyFl
9YOeGplPOBvuHITGV58OxD/XfGN3T7BSUcQnTQY9Qk/RK3X4XwvkdSjZLCgNIPRO
fWBC4feL3P/+Q57F62nxr7ZO/Bm35nqyRh9J9tHRc+5cTX8cYvtI99pAr3TKZtxS
m7d9rdczoZyVD9nndA/wlB3SJKcNeq/Hxgk6qbllKe5ZHAk7mV+sMjxlN63eI1cj
/hyDGyG2AcblXBPgYAwGiSqcZRfyxEq1r5FkxrhQ49wlYW4l797ehMpq1dxWKz60
gDtDvioSaZjLQ/r1ZJ3m0rPgrfS8rojY3HioQ/LgGbGEcDqZg6qeK7/OHKUsYrkq
55fhdiKDZB1Tuon0bAgDyQ+6S4tisDVmh31jeoSAQndHKQ7u/Fr1sM3rWsExgqpn
KJjgH8TTDMNgziw9ZQTFyXtyx/ftHXJ1w7nMXfSeaXvjx8FwA6A7S+MSba87cNyZ
lDl820jb04JWE7lSKjteEI63tSn212XEEF3v6xbv8g0exYAANJN84n+Uqi9vCPdf
wGFBSdN9JXJPuSCJEIRNKxx7XW29s72FFdD9l3LpgIQ8Of0WcwvBvt81AcyzpFlL
C3pdp53/hde0dwOLiHbH0Qd8okK57q8uFpCRCSQ3Jdi3V33xtaDB6HqfpW2WqZMY
5Eci9GLpQfmzEDOlGWyi4HabxTXvMZ3a5bqZpW3R7Uy2sJ1OmDxClfvKYyNdK4Yl
bgqFU+Dg0WavKCfkRNuq6Whn5my0kAG+OgSTXrmKTH4JCMd+ZTWMYJnY9UFwNcSr
Bv/ST7T1DS4SaI4g4NzyKyuqfa8kUDa4vxcqcHhc0VS6p1S6DBhJnnQFQbjM3Bp4
zMqyqIWCrGyGNTqpVgG/BW5g3I95tiiYW+Cb/u1sZ4t1EUEmIJf5d95bLboQL5zE
N0eoPQf2rL2M4/aoqjsqaP+3Tx+47Da+yGwzrU6AFAyqQ8p/HTRyzxImGsn57cUA
1OCBAn0dLI0wm1pbe68TLcpKZGzcwr/wATc5bbcy/oOytOGvVuM9IRhnGPl6O9M8
KjVEjh+ousCi8EAfFtqhzOvLruOHI8lovSMOnG4Acn9YEXHWnJC++TpYZV1PIQDC
GNbOqkOrC4XJozRK43ti8IFYCLR7KtIyHTROhQQAePkhb3VNZCl3LNSa9+MXxYrI
T8Lx9qEictVMr+47VCVW2R8vBI0aqaEZiVcxNdavcaffpR3urEP8o3Bpo97/xK7Y
JviKmYyC+aj7ZAqjG+P6MXA23INvDrYHVl+GVk4I3YNcC1pn/YjIsBQ0dfMNlXL4
RVtNA68XKRUFT4dJHeAiyGpkIYrgnVdXzACXnzAJ+2mtqqrJe9gBzI0iSNfk+LTJ
lmeNEDAqZL7Hizg+Hjsy1eNSg11sj0Q2JVaz8Z5u+fAF6FNp3r25e3EJEpf/H22O
rvsvzXzU/bYxhB2rTZkzkFEIa5rDxvDslE1AL+os2AEArE5z+iTzkaqUUIYMUMWX
IqeG1olS0Ivuy6VK6vKWhSBafROfCsPxhWDtUM54HAqdlcrKckojDpoHxAzw7tiN
Km8E+22wnuEpPISo7hwsov2ukEkGZXVKecJzzCgTUcLhiSSSm/VTY/KcUZ6q9Xqp
e8vAhI9ud/gsTPBeKCuFbXCOVQdCqw0hrkZF0z6yDX/3i9mK6sblHv3D//ouz5N7
FhAPiLOPpAZik4fSKlnR4bpkQG5kfTW0bDJZUEAPY6iqE0M8CtuXZbuJNTGaC/Qw
KVc/OReDOA16CyR8U1Vxv1xZhka4KQOzScgW9g91GqONIrklyOrXTgeXEqdKwRVi
rUWMUZ1q3h1ur9Eogk9PmRGMG4Fhe00sNdhNpuzFsmtFwRoFNQTmXbEi0lx7S/KH
APoPJTCMkiTyT+dsOX0V13T0hnztCG+T5G84eTcIEG1ywNUuAQVgnX0nELTgn61a
iw4ZIHxAkeZG0PNDVXcl7cFqb1bIxn5SKNaKV6DXvo43vtj2HZ4DKrBKHFvdgsTj
mlyYhUqVqNpul8dFLafZHNJ3G/ZSkCi2Rjyt7fyTRo/fZYPp7zabK8uHqJYWrlzJ
+X9v/BriMAYuk3pocp2qWBZP+s1pw1vtOBBPTO1KvrNO3RVya7+NMu5YUEck6hN+
ZFHoDWQGMIHKexavRw6/BN9d15MtwwccazTuXmWc/fLntAxKx/jZUtWaV6piOIGA
0fXsZaGTYyytCzxf0F7UAbM2CJdZH4omiA7CGJCoDLsdgC80PwbpM2paHTHNdKed
Ce0a/HpqCBmCXIkznQK6Buf5MMjAyceyWYkTXpTALNFq2eGLBj5GNLqnDoGazzq8
1+MAX87uq/0qM8z2PGFTNJUiJoRItKxtFgTfMZK4W8mRMpBJZwmAT3NvPcnxQea9
aYl3T3KHMhR9F10XRYINpEwpMbUod8cWS276DFLsm3qvxZm9g4Cls6rHQgn2FuJE
VfM14+kMD8tmH6IUkC+aQK8MSgmRK6ZyA/kQQL4FC7RyUgNd5lztdlfmBbwHIYeU
GCxzpi+KPGUvKgD228NHXt5RBJSPgU/9VOxamPFS5MxgnrIX9EsMsRXTMlqs4GYV
WQsaUasTturiLOF+y8IEpDAH2+7wic+YWyqEHevaOrKyZpKYe3PeF56USY8at5F1
47WDvhBdVW8FvVLGv/4fKWXHBOtqGyfSUD8qutAp21NnMr5DvkOibE0fQHTghl9T
wI4Q2epkfICz1e0rSIeIhwms5uOQBtEjcdTlg6iAIeCU/i14TEz7BtmpH8ss1VRv
GtM5kz2kThJVU9O85M2OiQu3YesU8hZ4VuUxZLfV9Cnauj4Qk928OvQkKohU7oPU
oe7qsxJetC4i++FNh7dGlHJs/6xkNEV2vqGyKGE3wiRywa1DEoQmgY29CyQcGRB/
Yzk4sv7+KKy25j63GgqHSHWjODq+EHuJvtq12RKSU1g0aiQJKUY1UeYGRgO43aQp
V1EIurUM+Rj9RuXFlQlp18BhWzTxJF22fUOO6vm7DjJ3OhQY+iYso0S5ltz5jhXd
7rJKjXf3teU41zxSnf9h9c4XbtAR4j9eNm0AsCMJqHRd/wXYYsMTak44/4T/BEJh
pB/3ejiDRzXsMx2LphSnRKyWbRL17sRs7awjrH6e2CWRPdBDpw1rUrLNGsDV4ocG
oFzlFNoIwxrbFG2mdnXfHCPN8ebnfw/W650ljIXDefP0642IUf+S/Y+syRWfT8bT
wL2JPF7XFODq3P+NpMGVE1j9ZKQqt6mcJmgAPqun/St5O0Uv3uYAfgr33W2el+0K
Eh3YOWImcK3zuaUDnWZF33lofqkAnn0tVPymC1Vrimo2MReEzj0WaxDlW71Lmnub
TgbUM1v+ciJ5/gcgitLo3D6VR6NCDvT1i+0kCY/IP1ojTl5CvK6sWCyhj04IGMH1
0AIpKF98rE9mJafVTLXUR7up8UxA/7ngJdXBfg9rCDGRWnfhpnBBXMXcgOxdApe4
z8+f4coCK7jMPaNssMNqo5ceg3Ycawju7sTyjWsiDa5O/hj7y5pCWqlLcjlEwdI7
Tot3Mv0e0W0byN8rRXIYKzOfczpCttucKQerSVU7+aYVeFb9w9Tb0BRN38N0cj9C
N/PfwzzkSDgyNnz3sIYP4jjP2cMbr/1Aj6a5fOx+M2TbGgnAgOsRTsXTZ4Mk8ysK
bdCNNdWraZ45FMGTimPwA0/fjfHtzdmDCMF/77Q8ZJGByirVO2feZBZXcpCO0Rg/
95SIldUlgWr0sdqJmw4N+ZVzMOW42Er8rpFhKvGBpaBIcZUjC1Th89Ln0N/PfgyT
K7PKnjbhNtnq9V1rtjX2yzF14tiZ9ZnjKlhlvki0PIUNU87YDzPAdGuAqO+JHxA8
Kz3bQYGMcaKjuEtQ5/LC4H51JZX5ktSPjeL2tx4e6Cji4byGHOZxwYgXbPDxCw4O
lUuCsdVCtAB30kQmPdWwo2CMVR7IHHG7FqoWp6qbydNh38RfqJX5iwX9jk6M1SkZ
pTIoxZzpvROj1/q7z/h6OiTNEmAV/1yYzHTnUmxp98D4un18yTathyAuPFhV7ZCx
oS2WoLGrU8RgfZfl/SHV00JYn/xZ9O/iwNwbP3qbC2ckkyqTgSW8T3YljPEr9ojJ
Y1saytPjQtxtuXwugvelH+7rthvwWUCUuAuMNUcitmTH73Mhzl+dOrxyQ4/82sRh
zHl8MJ/GXL6QvK7m5BnPx1lKq4Q2ZUNUmLiLEwr0TRz8X0NnS/U+d1txrjUqS8Ey
cwVmVmmGjht3saxu2KOAivEddA5nrlnFobpM7U2xq747SUqswUKumdRpTj14g12s
/KPaUxMevwWpvPGtzIZ/CDFqr1Flo5vFqUzzB+4itYuzcHIyFRzS4wYtHFomV7Sk
BwQXQv/VvQMA7p8uU6E9PNUVuEDoC7TNsnth8VVTH0BXo8a2FA1rW0Phpo5sRXeW
Y4Zppx8Xqv3WDN8bFwRTWUT5ipZfJc1UMzeI2DwxwPqfUMdLF0geZOcYe7xj1LI1
KfvidsKBKT0FmJdbixiD8e06dq/+/DUq8KsuhD/LpESFdSQwpNh0kWRS8MGQkufp
IV6YWBTRBimaOXFpWYgdZdclmmBe66OMekmoImU+J9qQJcM6wYESoIwKnU1489f/
EH93iOnbvXqXZCfrDMbGdYmqNXf/nAx4OJDOYo4Q5B4q7jEloreDcpA9Ke34ljQN
adTLxzLL77/v+66hMsmUf2jW7dEVIi0z/6zpyNoCgLZgSfa9H4AWhG7KwyZCF+lB
w6rCe9VyRfRNt5dRm1hHO/MJD1JLGB5WzNSG5sq+q+kiUw1tt8c+86nI6ZhEoYW2
73xEq7+djcMoFhKITAk1dJqZcKhnXLYe2SojyO/2jTOln5RPUebMDtvpg31FyGzt
J3O5suhs5g3+zeBs7zcYqibxwNWRbhjiJS1zQ4Kd+2Ku/p9nm6bV2d3ZKnE0yENy
QDlnTzMZoTPsXPYRsvu8g2BU6DxsYWCQikesNoEH9AmR0TsR01mwK67ZAUv7DDkK
gN9kpQIST1IQJUivdX8di6GxNHuv9/oN1R1wLecrbCV6TEJUplUCG/eR8mQ51Dao
lmyMtc9Qk+xyJItA1oB73bGP5Y74m+yby+jOpF07Vp6OLgwna2VWCvadnrzNeSBD
7i1dKAxeRrNd9DEHoqrt2Y6HVREkoxZrlkYZVIB77t5Ukms0eLEBLaVnzX7sa4sR
xv2REE+JCO/UxLki8NjcsuBJZJDUmW8SwImTtnUA6x2Ud+ZwyoviSWWEGdVmeaqP
yiRZH5y9ngSpE3VR5jOJ264NNhiHdejkeLVbMuxXGzdu2sTQtUoCYHJpDXGmZzTF
9YWjxjN3qcC6fPWuKeHxE9VFsabfdzYVfrAAA2n2pT/fwci+uMFG7NUz3Df8p8Iy
ZZMubKgjbn4ZaaN9nYEKWqLYbaDpfzIr3jVwKocuI+mngeRqjKH2B5ZTp0tYGSX0
JpE+xmNs2jd8/qHn/87v5V5N5do9ot3sL76h7T4ksoQajDgJqTmxtxJIJ+SPRzg7
YJSAuVMheU9XbbTktQwgOdF3dbgqN4pJaUPdcETqJ2jpuDltDIbUbn0If25qd5EU
XAlhcaweT+gURAmXxdADr+UVMAOuH7ZXlOsKrt+aL5pS2UMQOPXMHOdp+ISvzq8s
/uxXFYDXB4U7Ts0lYuuYvEgpUw3RJIeT4Q0EbRwanOE1zgbLN3e35hxKyoqjO/TG
6KJl0oTfoUO0BAkTVXbqqY5z/34w+Dx2ZWq8b/d6QdgYApdLsvRWNKoP4If5w+tL
9ql6DMTIyHoy7NLqDyR7V1++V+41Wfw3x4DQLTJDZIvC6jOHD8wvV0jYSh86eZS6
QL35fV+1LVawq8h7aGWe3IPtATLRjCWiohzT9SkcM4B+wK8MXing4HJDxmYDLd1/
1zGK9P2JOOdNHtCHI5sE3IlUAxwN+P8JVY8xg6tc+Q70RIR9wqXQaKqhHGlLvQv+
5SAx7xyZ596CZUivnCRlSa4oCdeCd24e1YS4YxPwA+0/esBy5Q8SO/+UqYM1p0Kp
HCrFZetrzfbjXPbVJOYNXpxIiQdupXbZ0yPDSaAvxKx1tz4/Cy/ZpRrwD7EOIyFv
j0iiaAKQEsrGPAy3O1Hj8e62fkqCiVYXkfSsRPKIptJWI1FBacmfsMbSc25vfrrF
t40QjG9sXnkvyZqYMCxmDKKn8tGvG8fMbEJh+Vktd1LUfWklmp7HTPLzdlf9RVBC
/Yfr7he3zrWpQ3C0foyxDg1Kx8wmclg3HTmhfssiBEmjWNc7BTal2YQYa/SaAIRo
IH2FE5KBi38OeVGMM50S8jW3iez0UcgjlaTGeaXF++YI6/rrLPU0OQpuwdjgIOCr
e1vZx3/pdR6WGAja3W7vVrn/P0er93iViZoXZwN7JpFLXGyFeewb31YUi/Q3u4GK
GriZ/FlARWX/0xw/mmd54AMBahgBPZ8Oz78WHggIrtF+t+MVDJ0I2pGXwFSR3med
li1MLh42Pqs/f6X08DDCKCnwaVuAHh1UwxpxqsyHLz5vtWyl5s1kQrRjqT4b20Bi
ebjRdcigUV19FTezyb6OJQoKQhs6NIHyjTizAnw25mI38sTmj9XszEg/HiCqYBcl
tVRt3fCghx0UTUhZY9u2ddybI+7LcApb4rRhkJXVq4RuDE6MyJwNJdg3K8u5QDSY
1EP+9wmh0Iyn5iz27WYPJfkYDPjGoUSFzarouxJ92uLibKkJ1LKIvp+uPd9Xhq/N
dQCw6DVpQrLulC2OMm3vImluA2JKa09H/bxijCij+6irEteSaL922oeo9xOCOqRc
8ynN2XZCs+HgowoXWr/wvXNSanDpFCb5pW7fK5xJdEfayCBPGI5z67Ar4UoK0xdL
U+w8UIze736B/fj8761vK5QUmNZc0BFYe7AOgFeG2mwJomBHKInRPNmCrCoCD284
cyWAAsmPC3Gl5oRJWY+kuKRb1gzPB7BPvtzCAk4EA7fKDOVHCyufGOweiqSNOvC4
PrMHtYonhWUADTCfocAETXNWu0BXQCGndclyY8pvcg52GgHqM8aLl2hSoYyjhHar
+nedQQcR9SWz/Yu4KnMGuEybn8aZsG956VcJZ4kbGIMLUIKoh8uVkD6zK9pGTsQ8
576Pl6aenld5YwpR3drjk1qsirhB5L5OgG+CVbWNjNe6uYfc4Qfklp5IMVclvW7m
cYA1dpVWSQNPmEAKyiZXfXs+a1HqF0eQUEIDlN8pBUidRkn7paqZic8W5X5/0pXJ
RBAU6f6J88dzbfNliqe3dVzJMz+OfENhqxTMMKcb0VAcimr08l6ucGgv/580ZzFL
MDJFfhG0L6YD9qKj85aeq6S+UBAA2AYz/VgTM+BZ/chfN67TtP/H0Qq2QOXDB/H3
P156rqxbQabUi2Btr6j+8h9gr41odtUiAzND3hGkB9LeKOVMtF1YYZP2JxpENVAX
tokFVFJ3D1PHDTYqOyYm1QKsYwBfdtDfpF0qlhKEIkB1M6bF6/1qvDh4DSWKkhJo
Hq9ziEtHNHtVbPdFIpB2tALfH3mBFdMyzRfoFFGQcBIupxlcKWbZ0o2Dj7rbJR/i
UxVIr9FWulcdlW/bslIZDc86uTVN+2Wk7Hq2/f5STB4bZRbdehkhm3CXgUoUDC4B
FWn3Lj94mq0rL9XCQL14hrjFS3+WGMA31Urjd8qLdNxds0BP1kR8k1RYO1jYGTSf
JeBDdQF/he6oJzvNA/aeYBnKPz0ZRpSzLRXrSQq8c3QYDKNKXU6HPlR00S4Fo7rQ
Cg4yNZA+8SopqiT8BfvfZ8SQwvhyUdFhTgWTmwjky7/FxzVW4pEHJkhp0JsWEIw1
0GcKJ8EQr6RqminKXhppcfLwELGJK/I/ebn9fH1IJgIXR/gBuMBRdDA82SfwiF0o
DCgNS0IJFFf/cHUAFHkSmrHUdHJuAF2rlYMf4eVmsJ6tYhvu5eIEyhaJ/YMV4VO+
V5eAdkaAHE5QnfNNpDYnTcyEHcl4vI6MfJE1XfR1nCDCgNTcMDEFAIptB3mUtXzi
3GHOX6r/6s27iFw9ndk0Z6cYvzlNtBE9/MjbARcOaKhx0G8BqK52TxW13z7zyVMj
yheNjKkGRjW+Z9j8gjJI2UVEvMcpS1A33k70xC2ezABJmJJAm3hIbD+1Tgr3SMmW
bP5iZjA+oYE2XLHWS4g+FALjglKUzc1OXMZ9WsPY9UgB2D6qRhf3s5sebheXrEtb
9mFs4TeRrVKQkIYQW5mRNt5nU/hP9UpSgZ6SFm24po3+FgIhXRnXAWR2P9YX9bKh
yHX9x2nTLPhz3UjWUvjMQC8BE+MMIGcB7R9DKXQe0S59TFv41fJPTHPGxpE31Ty6
6C23nHPsBBRDIymBKHuKRU+LhezZbFLhyWd7lWRX/7SWeh5SqJeYUBBLhkV5mb63
JlMHCmLvWwHU1OjwzvA7AoQC0aLOKJemw4xO8oF5K702wLo/C4X3SRrThXi7HUEW
8K+DOnekeyfTls0nJgZ+TsHQfc1BjCTu8f8PkM6kK2YyWH4YuZNcWrPxgkCXv7fC
VIrPHIhb/1ggfX4YthVQC2bQW6M4zidEqyYivZruhLJhq46dn1pLQcjF1hoV5PkB
zW0InaluJiogMBDoTnYEbJxWhHMH3f8rvm5jbnkbTQ60UjEuZ29dNKh+0ldjcnno
Ttz1g2vlpwd2gQLHoN5fAp/3oS0sNkaMP+hLjlHWzkrwW4lSFtVniQz5nAKF0myU
gAhEnxcYgjjR6p9p+eafhunxZgxiZ4wYbb1kGC8XfltGtKkOkTpZha0PyUlalAqt
D6NdeieV+qcJWBRRSKxOCFepLnqVoX8860ZcFzlhpr9W5TPpipObj7J6VpbJhvPo
n3uqtyzo4nfFEciKh9rp2X+ugShLKpbYqeF/Cc39dlyKXV0qsLrhatYIapTU6q+N
KujFYgNFHWE41n427JlXuKqufgC3nDSXskEKwIjViZtXX5M3S29mErUtLHPyCzXp
s+1QjlNMYkujnnLy2GSi4yDoX4clNvfKhgtinv6f862Hcfypy4OH88DAQnmP3Rqd
9cHpEO55sYWkfqa+Rq6GO0zWT+Ap7dUNkxa11d7zu04h6xrz6/CGk2te0wohjmYx
oyTSjcRn3w6KVnHOmDpZkbuaPzcQX9hmb81pvwUwSK9AG1wD9/FOsZc3/0/SzBbq
F7Nd2thrZywZJdzA0kZNEBnAuVr4x/CrYrR8Oki4foIRlTlZpzrEgrl+oVlPUSbE
HjjLGITEAZeNZrls8+w71dYjFNo4G+8fOcrm2LQnOwSPENtYQv0UpvDNYHk22oC2
dXDIRt+YamsNOR+/05NRf1XxgpdMntyyVnpT8PUBur3CCAYl8KDFA6JLtja/0l9l
o9+MdQicktCEA41uDnlUgE74eVeOnVpV0oOyvyXljmv5UqzwQRIOI3jkiR8IN9ay
ErQ4ih5Gc7TdHSZM61YkKFFlIdwuTYdqs4IPcsqYwQKkdcroCWt8575llhF/b1lM
76cYMSuQqj/iZdWQqqCRwv1GGq6/1WSmPlbuAOG7su95pk/+j945I2FNirMcehFp
IR2DBrzT6tI4tBKbq52WnNiU0odch4V3JbmXar8oau1SHOJRkwqtQjhhgptMA+u0
tDYAUn/3/1503BSGD04Cv89xLZ/bsv9iJ0aXnjPtvGxdiCX4UEIZXhCYw4b7AdZG
jvAAkELi5UTUmY9jYSVX7hlnQ2SvBRRNc/6r+yxYpDskvHXaN/ZWypFYgmXDEKJ/
CUmwE6iBEepbo28aiMAFWtnzGZ9FZIsV1+xeQVDs3O+MGar5GoIm0Vov0Eb3nZB7
oZbT10T2sLAhMzZ5/7lVh7+mdBriQJUxYDgmR8dwVT3Rqwbq7bk/Z1U5Ev2VZ7ka
lF2oh366BCLq7KM/uC9pZyNzZv5uFdUN7XTDmiRKvLHa5NNpQS+Y6OmnXQxEuBSL
DT1CyioKbJ8RqV/ha9F1jf+eiwspoDOeufqMSOvR9dySnqn+ZCc5GG062ckT5PsB
glGCo2EL41vA+vok0t8UWZOasEz7ybY/fqySSQC6sKnIWK5UW43dSqhVGRMN22bq
GKN5BM0fJj3yVol89Ls2xkQ2KUNhc5EGUaqCD9nYLEz9HtMXy3QY2EZA43HnsLBY
0LchFxFIyPi6GCpJgKUPIjjR0/bJY/tXgcaAFcH1yoq9qh+Pxo8sRGFL1FPr3BXA
pyY0/kwpxRFB64pDUmYvwJ36romVazRc+A3sQFGw/YvBPz7dlmymnkb2tI5aSNc3
uxA1bahKPIXMGUTfaHUZ1mzlRIgbI1Th2YuFT9jitvIqhxwryLSAVDvSfCELvPiT
nNnIaMgrT4cE7MAZKy33shJiS8vD/Dc87j+vnYHiC7TNviaehR/4I6GkZA/n4IiI
/TuEYT2WUrqqdG1UqhTIxFMHCvZEZCXGXptsv/pElrUxA+8dKRLHegbbYpsYLKXM
1jmvYk6V7fTgL2mGqP3eoIEZwB9bETKIqppDlfBDJXWkJSQhVi/kj7beCWAEHweI
TFE2E/tzhlZ3cIQVB3XRBU7czHq3LW7wAI8fwW3FlYF9nVq2+HYDRrmWJMeBy0Ti
1ipv5nakvgyrtImTOXxYlPO/GYDjhPxpoCIxdF2P7YC8koMbI0DTAP+XIR10WsTu
PBe3uaa4D7T3LlVr9/bQDboF0k3P/KYqo/Ecyq76q2EBGl9rc87Sq06C1KI8zi98
d1muGakHP2rjHvUsVSSVuJlzyEFEMfIGI6F3SYScPeJnr2Gev86oMZmBVdzmSgHG
HXP8SkndzTYqQRw8B+JM7EZeC9VGyA0FkFhAteVxPuX7suFikt4oG6J/hWTUxfHB
XUveRczMSKd3WJPnxKttkl5TTfQoSblwUDiR3Z+Qn8i3hgu/iA5JA9GmBJSH+hHE
rHZm+xv0cAlcwMDpCkAt4Lb0T3aJ2Ehv3o+cOt8CVpaOpzdM1gP+Ozeh013nniGa
nko1nYZQFeLPNkRh4iVUkklgOdvsXFRWSMqeCbUf4Twr4uzjQSkeqik0TcigRNJK
G6NMP833mmJuc1QuoKEEV56iZ2f6jq9Kx6w5jytuBTHloK8nKJKfmmYjewMcmEOu
R1NwB1s29gj6sNNk/647UhVCHI3lbYe75MAmAKAgNvBQL3F1S1oUYgu0LjEYR4sy
AtMfnsvvrlDyBnFreUZQBF8fANFgr2R1yl6ucK5ZEwu9uwm2TL1s+LjxwbTJvWOb
e/pJP5XYMm82A4g3oTij/PTnL/MF7uGZru/ylyFRXA3YBXdQN0+0+tiqSUanNwt3
383IkGCq84oH2S2VmcyLY4VD0KZMWamI3eGiIK1IYC0m+wwYI8D6BMbvf30RrKxR
GtLJ14r+cMTIaV/krGLWKPlA1Ya04yz5WfG3mpvVdtr2NKW2aU5YwY5C7zmj8T13
ghXmhguGZmjVOM++tI6QUfHK60v7RPbWw6zD4fTmV6ZEmWZfpOCshYWgUCAEq7HP
uYr3VpZmzWpQxrU+MEXWJXRnExIXsREYfe7G6aPW9n+pKNXBD+9HJCIMCjgUQr63
ADhD1HVFD5MPkDb7LhOYVtGZfpCO/7o2x22FX0n0GTG8c9DtClqBL0wAmIk7p74y
fih2QsDG+T1mvlMQ7npUEmg8MgiRMjG6V4W8uJ1QS6dFgzl+SIoZcSdymVGP9gW9
Fp/z8hKWwsmsk2FGhQ8aTfzDNkwB3boPAl5P3pBZgFjfg0dKBsRoknAUVuAFw6Cc
wHQsjgutf3zTNQOSLJ3fjcZcyxjBBgqEEDiP1qd3LUWBSlc8AhbhQko+AQ7PwtPK
m93FqVZmBoxCLAutmJ22ebN18W0pcu+WPYe/lTsIAKsrp33t0mPay/GNwErhtoAB
IMSQ6P8ffyG0jVEOhBYBlvq1LPp+94OFTyDS6R3MKBuBzOUVlv+V8hpNAM8zi1KP
vo+13wZihccw6aRfr5NAe+63bMRJpT2cq0rlTNz5PBl/Nwv7M4xiQd38F1OfnSKe
EqpXqdXyEoOWw7MOYwHTv/L2XciXEPsLoDFF7+Hi9SwcYDGl8OHelvK751BcZoVF
19uRWxyKswbBmphSCL1WbHjBn52Kqk/Ksy12MJjnbBFsO/4JACgl8MChXcmURtLG
ZGVo4HIA90FzWsxmecZ3Sg04mftNhh4MsCDss3K5J4WJq5fubcj0Fgx0m3I0irnn
D+rBCpD8Z6CN23CDVSNZQQ2jeSVklJMCj8uBM8l27voQZ1cPJ6hAz/qaTrPzJ5em
r//7Emk5R4wYW1lm5vTzbHZcoEIT971nuH9E9KuIsyfRy7gv36VUwcfIw1kj2Koz
4kYY3IMClgB9Bzvd070jB5u++ODODGIMUxVJVsKoHW3CrK76pbxdTe6He/nWE+IY
eMhGnB/IyDalVoo3rSh9J1siYt1FopzDBy9j+7wWEHbBKWlxsSqnRszBIEOwO46D
oatyjQxWoWLLBfNXVBiqcSzdYFRjMfw+DKwhpDT0SOAL+ctg3GDFuvCW09T8DIDa
dlD9fR1yIf/mPTOEXB/bhukRZDxTe+/qe0GL1vq/UH6RLpHkl7DLuoYEkfYW8PO9
k8avA5CbzT7Gb4JnwpZTRcQXckEt8CrlH/KUNliVAI+6VqvCtf9evCgyYPZ/Z57t
enTjMF7GVjEDwMYK9XO1MKwUN9pZ0ek5s5P7TmZwtbPM8zIaIGalinYMAt5zM/DL
0zf670gtGNDCNSaJebufm5LhxGKCz7kUKOlv1uvPfBKKLUlTnDNoFYs54WJHpMje
Wqea3CyTDw7QKjI+97zybeR73VhVmzzcarBE2vh1zVzlgAR1VZeChPXrjyXWePEE
Ink4gOJxg19Tbjzabhpk62WGtN43UldRyqFKswViNrRDCCUf98/WsSFRXs5m10jq
lhUdAnYmiwe6UmQJtUKVUdJ2C6/EECwZBUUIE29RhKB+cvouQrQE7NU5PgVP0fo4
WtnB2nbLAgpWxyKudcikafQ78nY7qceGJCf+K/EZaLxktSIB2jSWwEsrVu0mEHRm
Y1kf4TcEOM+y7bCMJTEkXA5K0vNt08MuEe7m6itBd3yf+rrDsHbSQze4+4LKv4ZW
3ePRwGIEQvY66CbiyiGfusO4R2h3b83F7dqsJsNxrHpyvs2P+RN5x7Qyk0wmYZCY
GxwKQm5wPvrFoJLiogRFNmv66fEkaHdkLHlmtIQ4Os22sjoeD2Vm8JCF4tw0ulYm
Xf3mlsGVYsW6JCHIfKVWL+/RE029yLZmrWemX20gVfAtWswQhAx8N5n9KpR5XhpK
wWN0Q6AjHkcVGcgYd8MNq28BryZmX/KDMy+KCbet+35U7B+1nxRUqPsci8d8rA39
MrhJxZlgnw7ta7y1og86o4KrONO6ebM02/6nyqhhKMfXHZ8LuJGAkXvd6TXDAp98
4WnK6DaJhf85SWYV22Di4WFCJAwXAOpw4nILzd78f3JfEMVvNrgb22TLCyguomLb
Y5uTj5WYuIIsNzQ//LFLMruuuvn+RibwqCxl/DMbNne3Q1Rvqg+1088Sco/IeHm0
8Sre5daxgj8YTLLyurLuCfZSVg8spt8PK+Y6Si96wSmU67lQcbGnB5tHIMw7LJ8A
FL57IPp544JE9Q3WriQBzsdUpfUklEfTA2fXOJhhATQhupu5fZfYoFwzOx07s3+t
94hf2n+uFrHx6Wk7WWvmNk6fHmTzn3ShzRGlZaWn/3+n0Vvfua1eIlAecfhcfVl4
qKyS8exwkrHXbTW4yko0WiTgU7QHes7y5G40yyLF0p7tsSUPGzPVKCPi2J0xIO5y
mSmYcxz0AmPn7IX5JohbXf6zM/k5wFUGDI9M/LfxEX+e3dEpDnT/wScZUlueMFRo
p0cqpTJ6Ma0fJrzckm9Zt/3QueZB15TSjXKVLWiFD+jmhMm6pmHRw26ehJtc0aWf
3QuJrwNdHNz2vfqEKdE54Su4psKV5qYRF1+jZv5Pp64GF5o/IXVrqH0ljSn+WHV5
cV05pAmJt0MeTfGr5mxB26tcrCoRfDIDmus0MhXJ6b0px3ZY/aSxTfyuMuopRRuF
ELsLWMwCLySCfmUu9H2+qDYHscAWLS6F4UcYRbAaffiVpp7Kl/oJF8hnvsSDDoTM
m2OZE1/R7gHRkL7eUFbmISalXVzm6DmNBOU1HwNP4EyAycwdnGTLovnxxHmXgxj6
eQWtKejv0vVIY7KfU/ecK6zzHbqIya1Z3OiwHDU5Q3C0TKcWvK/pmFvDhqHWzHDT
cTt0EKc2m7unJlZnEgzV/G3KZtK6nQOMBbH0l0OH3P3df59K45Q6OxdXpDLVXCEn
O4AFIQejJuVccVWoAk1mvBO/7DyIogOBVzFNtuPFFigVxgx4DcVUpl9t0sF5mTiy
OXYXEVzTAXLJFSK5BTd6/VZzaR5lXO2vhx/KDXhMc0s7g8XH5l24cVgnrU671cBI
YQLEf+GJ00mz1ih4+KApJjF69bKBfB1khYL4CHLNqUHduywNqk4uo4fUM89LLU41
d3TB46iz+yt98ucAi62qp9eWQ93fV0qOEwXkoMyXNSsMp7//fXRyo6bWsjmV/gPM
8yLwTw6evcvT4EFzqjhshP1oBxEJ3Ei0MjW7PJKI1SsUrabWkK0U9JGFGtyFBqMa
5PJjWovIGNCh7fJbFjFQdA5ji6xIJ/O9QP6j7UgQ8HZDw+SoeeUCHG+dzPAUqfaU
Y7ogMtRFgTB7kmcA2jN20nsIPwTzHaHvd90b2B12DHDewIMgVyYlNS+nwYXvukga
ZvRE+ymbjB7p27Kgh10yVbYCsFCN5aYWfx1i/A4V9JLE5TlujVcP5Z4fwTYYLEOy
w3HAyTW0ieSPEdYj+27aHpFLKbLAlfrV3xHNf0XVQ5YfvX4qh5bxcobP7zwyPnq0
gNg1vzeZ77JkvMFMOo2YkRJ83IX8KnM3app/e2gatiNNivLlIKNKqNuANsKoDpJY
aqArNjmUI6rRvB6hegpYLAgLR23g5hJVzF5ynKVrQ56q2y8V5B0FucXfGii/diw4
AetwBq1jI/+3tYYDcXsVPNr18xZZC6hPYym0OXGvOcc5LHaspGsWaQInTF5ymFmI
6fvDmdNLXs4Rptu8JnpFVsCK7wYD+AbzmFEiHmplkzxOe2QjiQaiCzEjCSY2U95l
TKTOVvf1E/GHOUJp7dCKLSTckLFH7WBvzta8YOQCQyVejjV1ipUR/GjNGVx1UQzV
VlJl/ymnJxISQrJ+IQGywrWvD6O+ND2iolzNzQU9QKqeV0AExvYh/XzUoG7J0gkr
OZ6e8x7/lvYtGXZn0eSCDc5eAyC5sV+OA9XecoeBfiFevXLmg+OZwMcmebKfpcJ5
vyvIjrRC1fRf8DEHB+wbs+PdKd2KAlAIndHuN+7kk0yW8gSPmSrRfQ+n4XPkM+Ok
ksEq49SefjBr3E2E6Q6pxFa7nxExH9I07toL5OULRrkHFQNeUSgxtr1y7HQLqOi3
Eoa+1Od+4Nsea2bAPZ4848vFyGqI+nKSvNrnNSs90GPoWS9qteu/wCtiwrGEJjge
xtuAi3MVnEcX7vJ0ZNPBtiKFwsjKGW9lBl8O61Q8xUPoGPoJt0vtNJUtBAnLULl9
3rdKEHQMxUUNtuC5Yn2+lys8IQrUEq34DKPwQ6eBIHkAgrOSVx7UsOPObo9l+GeT
XyRrht0mulE8m+F3iNnzxWbK6lA2DfIBIIhZzcZOwe353sZbQnCaTKihQUR+EvhY
biJ8wIDIC71VSNdFXUrcZ0Ee7Cv9TeD9PgP7EdGvYdvxhsNBx/42lSeR+A6zxueJ
uGGrXWT2WwMGgED5MKZayuEL+gZlGa79cX4ukFtqiIT0AzZkt8ny0Z1R/uD5KGYD
86nJH+Q2y1kTOBOUo8HoWjf+jS15ue0XKJitQNhaVHOCGbRt0HLMIL+FN7YdLl7Y
7v46tR5g9BlmzKDfXNEB+/OK1BKMbLA+B3WsmF1Kmgut+p+N57FW5Fc9KUm5O4Mu
Ysmy1Js1BiJmYRGDYWArl6cafQUEv7FgrickTBDweh35yDzeVqPl0HWuEwAzqXWA
`protect END_PROTECTED
