`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C26jI7cb7fEWaLeS57yxhUpnZVfGa/ylmDkIdPxAKLHc
mZbz81sJUwMXOvEn+7XbEyd6Br1FcayOWyFLnxnVMFojK20sLE+jOiJZde0yiA4K
/NG5NlOp/e3FF3rsZF8gOG7pky4X7/lLDfKYiKbg7CD4FcYRz0nGpoKcW83ocQ1v
AFXui7i0/Ho1EqZWpwQpuEvM+4/tt3KLT5cQEMWWOYI7Z06uhCTuGj4qVgUaI63m
Vq8PHWdibHq+xzodaEI7U3JYj59rT7XBSQGnKSfnGK8Vpy8Quzxrw164noTaGtrh
BCeMjH2HxX2RtvecaUSRWk55NXjUHsKnS94/3f1UwqgwMghkJ8oEVEwIVqs5ZYmf
euxaP4LaejI0VLOjNgtiLc6IZ9Z+GWoJ6UvmPPfvM20HJdDriIAEz0GcdE8qUrEY
2bso0uMtKNPIoxTNcyRNtiTkeJ7895FBmjehXxyL2+89C14dDJoCM1BpK8l1yCAy
EA8w9WoK+uAVJLvGXjWrd/vzcAv5cS7nRFiuccv8fvaAlowpAvYDz7LOSC9yeUrj
lFnrVxC4Ih9EcNkt2plkqw8CcvcC3tYeuhbkEJulgiDx/agpZWH2WPiFKZRVSVpR
GmCqYWLctFQIVsUHhy31zhqMLD1OgdQChdGcSrlr5nFURB/XZVhRJ2nnFPEMpFjn
tKTzbALLknuF8FY9GP/gwgTSVvRcsE3DzLefsfWFBEDirvsc4YVZmH9adTfAw2Tc
moLelfkgamsK2f/pzdnndP04e0Vimn1odUxAeL1K6JtvSbxeTXkAPaAHqnn3QR++
iDuoBz9/7utm3IEfOx+OxylbqeLRsQVyf4S4ieEr0bGzm0gxV+d7hZPhYFuYfV2W
sf76LBG//l1ZCgAIhO8zE8SbvvqIDIWzgKdolP52xqBF9TEdKtF7ohBgHWp4pBwM
ZUhw4ZoMZu0hzmIHbaN42De2pJcZG4/2jG3oaBU3uANHY5M68q7w4OrmJ3AUlESK
0ZQa/vZoqQMTL1ozGd0pMuPUpa4EngYwmnCWmCy9vBFf+lgU4gb9N153YO5vX+Pg
KJiRD/qBWljPKIEYgFXOoFuEElK13afsLEmjCNM4C+29wJLnTqyqkvwRKICigEKv
HeZBN+madbY6++3Du5fqmxVRPF/iU0KVBmOnjX3rVgHvmHdeoVIuOlJ83ydwljN4
69ttBuL3S6ZW/gPnNaQDD32hD/xthHjlPgQbJMUVknWqrBOCUhh3EQHzKeq4sdP9
+K+eQUtLGvVCkFR4u9X9pVDCK49H8EXV0vyRv1gBQIHbEMABh0eqmWQXrL6JXDt/
Fg+tv79f4uRD7tYGIWURBTFaXJcUNJruccOXuSx5UDbDRTJ9Qj5tsaPt/53x1fh7
W0GrGQy1moEPxcy/hUtTxErW9RpuXglKiqPHJWquK76or48j4JsKXPQZVyp+EYgT
WiO1VsEQYnG1qG74D65lAUSLTu/SETXwYT4tN/tr9htvekqi3Zi+CmNb2aiKaKK7
xADhV0npEiciWT7ysJHtbIu5eu9YlFu67YiqOIMyJpIJFMvnnNzh2yeR9aJP5NFu
`protect END_PROTECTED
