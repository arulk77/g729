`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveC+hlZaVkfETKvaEuBY0LAM5rwb3jeA8sYCGngz+a8eB
i2ToQpzMJZi6BNFfFiLTuGRffA3gHO4n6SfPAMaUblObtrDiJzygzU6yh6mZcUDJ
GRBcMTb23+/CV5dY3l8F7/3vTun3hI1m5LLts7jQ5wxroxy9clUgGs6MKpU8JOGn
rKyMhYxcfpW1HQScXjtL2LWguu1Ur50Iij4/O8JQOb/HhVr5EagngXyZS/KUBlDB
VOI4Jx/n93WWdCpOk2kWNDbOhAQrsvPPUjLgt5rU7jUvYzsSApA8/PLLbkaYj7i0
4hIP6HGtsxh/bzZknuTbOS2ZURl5nV+3O03dFR9L9lecmUzGJakV92wQ5015Zsvz
Frsg/QNbBZieP109SDVWU3JJYhBcO/24Tw4v3IwufDR78lv28EG76t6UMsagkzOK
F78Lz7t911KGt1FUsOAGBOmLD6NaOlJadWxrCr+wCWGhSzf/btCoHhDTMXv8aYll
jSpgXnInTJQCdNF9j+aWYM0wcJkNHazp6m5/YCdYlehs2m7noaj63lL9j2wSz8ej
v/mCCdiMcdl2BVXsb6afuelXP2BIq6+RGBv9qRKLlf7m/19RFJ1zEUl/+oKYNMe/
hCXhtaKK5cZCTa8XROjIzcLLe7ahgzPRDQPlGOtU0K4Bf43iL2c1gVAo5eRzwI1n
roNgOX8uaSkSb1LY6h95bnarfYsx0+VRQo74aQEeLcLqfxGHY24q7uCSD1ZOrZ3y
oEK4kEnp04HmBvJ9xFCkYPZh8sEpE/lk0tTZCz891kG6FGK25q1DkfRm2FSn0rCf
`protect END_PROTECTED
