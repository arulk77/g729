`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOx/8E2hO+1apLjgE40FNzBj0fkt1JNXY/DXLl9ssVta
XG32sGrex06f9HhFCGd/u4mNPjjVIvsyGaehFfozYOdl43j3mjP0PjlqM/QSzEKZ
FHQxVFxx23XOVrKv1cfAPKAhzSeGKdm/Sv2kDjcveqKwY+ITa+0gIYm7Y6eJn29k
eR7yM/nC6pkcbxaOCLnrvbdekbds3cWhN6cUcgp3SmRglLK/rBi/Hb7lpblkZX5l
WlNa8BSx223TuHl///S4uI2rydE76GmgtbhVPlp+6p+F22H3G03ZFoYMOLempCHv
Cz7voM1+8WSxAbhb8YF07ZMnkvWpVk7mOftMMpJw53UDeG16FR+Gw+MW68teANg/
VFjcc1CBDQnyznCNtODwG+2vctyZ1C6tW+aVxIabbOIcXEIKEgX67dtEnvhTjGTp
joahKiy95aicqDMyaFG1z1yvzKdT+mGzlHdUUM66fSVq7ZN20XkeSsuySF9PG2W7
jNH49OoKzqGKri/8sQEUTGHiRAmLYQ7aACfkK9O6c9LeFDzL9Xk/LVrhT/baWR1F
`protect END_PROTECTED
