`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDdcdvXp+MXkUP5zaWfquYsl7b9blxTKTocwb3ti4leE
+Sh2Q8Mj9r7OTKqmwKWmkuGeqpaoTYFTjMJIh0M0xl8pW+xwYRf9l6TlLDKAjQ6V
tRC5b+eVBP86sG0ivGRbVOLQDda+b0PK2PUKnMl9LJMUtT57pYHiZjU0+EprdKZK
QdT+w3iTPfEHSyonL1h13Zx/B4jZxtIl3KxvN4Dlt2pr+XdHpG9Ro2HZK9XAbWUf
`protect END_PROTECTED
