`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aQGoXfDkjaiHYGnNLWxk+Hhu461zt68Yeh4NK7K0Kil0
66nVH3JIEeB/Co08wy2UfRfkQd36kS/PwA0kTNXWrduFAqGqoJRrySqHrLRLBq4X
GJu3ewnjE8MDQN+Ze3Wa9llO2ktG+sZnJ0ILcFY3h8aHIXwXXgWv7aF7C1FaOjEt
pG86pm4xWJFV/ulAOwDB/DDHNdBKzv6GJnZxs4zY9mPGIXtcezPMxRKj/oN39hRN
+PCEuWZIOmhO36skKAgfWb/XubU9fkVSYC49RDxmwo9DdJCJ4bes6z7XNk30lKQ0
mlm0qciUJaW36p34DU8Dd+odKsNSEl1R8cte4rMU0LpNNx2JelOs4PZ/D6z5XtDn
XoTnDqQuJZNDNzD3K/D9AJDN0BB5OEbQHNgAJF8MT2hQAkzv5IoKncgW+WRfrW9C
47u6su5CzshFv7SdgR2avLwi3PxOe8sLpfqTdLrqLpAGmpgiUlr7SOI7ezAf6p94
Txoo9FlbeGw4BwHxaqk0QglVy9RZLwF1XWqIxa2Oj/1s+lufoqFlYt6y2tsTj+rf
O+cTsbDGFHxL7GQetnnGz6+/CI064hCmT4iaT/rHSMiA9y1QDOHAm/vGmEQgOXfq
1/k2tUnnMNKbFMJjIe+SdaQpgc9htNmuRKCc7OloW6/jDvFaACsejVUzDc/xVb6q
v0AwfZ1iuQ6fWbTWiISDUA==
`protect END_PROTECTED
