`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42t4ULfEM6h7JRiXTVsRXQdoCuuQHWMZHkIuwCEt/y8L
PTuAkhhIxAQ0kAzLKusq9KuogRND8p/iQig09rM9PLCYS5nuYOUi3VmeXUU4+7vF
YQJqiNCZunDaNyhmUSt/W7IClTvJqyv2otFSl9HsN/SvZk+GzlmISi1hVgCvy8Y0
2ZbnmNx+JsUBG/T7a5lk/8oLhRuJTHfNO31h118aq6iIil4dvoxzd7NbL4IsVxQe
21YoQ5lWFgjSLl5Y3IiSKFrdv2qpJcM5xq0nCqOK0Fqmy0NujOdwPU/xpRnZmTIp
HPPQ/VgXM1L/7xDyvbVGf2gqAV8Dr4ShVtUdPv4AYRdhQdRkxWjbtQrPnoc+1h7n
fJHOgZx88DP/bmWC0YulTOHwjGDnLOU08dS0DKqKDNeloBJrxU14c6HBJSdSVbj0
QjlEMXHlRokSorOHWHnsVJgW2vPTBRBz0KkU9NTsgkvEowVf5Jhvds4xPHDMibw5
dkk2+5hMXAGlvQOMEkrtNA==
`protect END_PROTECTED
