`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
e0k4/3dUb86vzCElKEVqCneGBQz7fIc0q+aWgZSq7nj92WkQz59nrvipjQ1QGkim
+yWDsi0a8qKCWhq17oiMtZrG3RVqRyHQvAb5Zi6t4lBmozZSJcgj8LNYO/bFcf5i
YPSUZgHUzgDhnx7x3ky9MfK1yHDGhIUwKUkuxAU6TgvN/WgHzTC+ch4/T9Y47x5L
Ui6Cy8GonMEJnP9kXUuNOcQ6S5xhFGbqbRFMItbvGxSgAlnDROwJ9AVJ+b2ZovhK
KyOL8ToKcWzzrV3kUdWuBlhEJNUc2S3qLKK7ndqbnsavVsiGrISOvyDYP4rC65Hs
f0SWKFZXs6wN9z9V73THMZGDmPWxvZWtM0UDLA9tMvQ=
`protect END_PROTECTED
