`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
9x/0HsEpq3D5jYbpbgLZXx0cmjiYiNGm6SMGaYwu/wOWEKLN9jZvVnZ3qae2NgiN
RHPcT3jJ0+N7EfUaYaA1VcfXZqt2uOdf+c14L9IkghDZk/+rY13/dEKjCWu7uYfM
`protect END_PROTECTED
