`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEwP15nry0CsG8jP+UPPOGH74Ih7ULJOg4x+iFPMOZCV
BNi5KHvMm/08HdFrLa8+8x4rjr5vbH2hn5ZbdkvcZQLBZZ33cbY/08fDNDWAp3hn
r4fZIBC54yATpoBp6nhtx+ak02Ipm5ZagYV4PVrkE77brZCvfQATIqkCmUo6AZui
vHcPNJGY8W5p1THIJjl19Q==
`protect END_PROTECTED
