`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePj2Cm/05c91ryF80nd0VaLcbtrtXOXH/2mjH8BzIWho
U5GEeSmZRkW/BQygPJFEOVCZxr4I5Yho5fX8l6TTtv2qYxrUWlPCiGYv+NmpjBrO
d6qiGhKdH5y7jHtb5lz28S0kby3iI+wdY7iBN2n5RND8s1aZttRUbgI50zCd4Z1F
tpsHIUt4zTm1YwM8w+w0U1Gu6gZq+HCAW5dtnxIA8/FBYNUVaaz7VOkPjAlY+ynG
`protect END_PROTECTED
