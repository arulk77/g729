`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkSsMp2ukHWqyUgN5p1jnLfE6y0asY8/QR/KJMOz7iLtA
SzcbJtpDud+GAPIBYRMAIVeSbCj5gUISo7YMt+rQcd4JKJOCO5RkhzAVRt3YZs/w
mB8b15PMEJw71IBxnObQgqNe0MKPgpGZL80556DJrNP+/OqqRRZHfCVnA9zgA22F
Qb75VJqxioVty01q2x4itAw2KgAeDa9whMJMC2VtLwn+3KB2wBPKExnKVs3dibnv
OkxfpdnhR/tqVv2fkYlmLK/+4F8ymCfHiUgINDwlO8PJ39rPV+UDIg0RQJCJWk4/
R9s/yg7XMhbhkpeGFxQD6b+BsgXuezOOlnyNV7rQcEfM5LaHUdBNiVmSP9s/9rNe
dikuOXZwm9iFcoPfuZKfZn4AWPih4HwXErkTv6fNy2oiXup6RpO1JCq2p5Mfvs2e
Wz3obVmwoTw/0IuJc6rLMJ9AZ0oYE+dLbR2LU57Iyxmo0+0RenzV+d0j2oRKJwNL
s+AEsZ+CTziguTAFAUTfETwOsjqrrXFl8brJJp3kVPJSZKxsaP+P8QGkeLjAwzA0
kZ5jg+erwtpIX8Q6Ig8QiHahGS+0jjjn4bZBglCxS8Z5sVT3cRLP4ib8k3OLhSf8
3tSMiJ+pnx7ZAefl2NLM7qvtw0mMV/Br5Ru3n7xWImjuxfmPsJxN75o2WOeeibtZ
SAtz4tf0RWp6YqaDP4RlIpY9OaW6up/C/wvZORHXLkc=
`protect END_PROTECTED
