`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ZfeT7st+ochF4JBHxT6ZDCa6D4/Cvu9D4mikK/3vdfst8xMRPbdCNADzdWhyBXzF
YyKFzB+HhymqjkJNOjgAtNli+aHsX9MomupgOu4UNtfZKH4+++R4W9xmJeT6X4iM
tE360wSZDk1LsXolISlPIUea8x3+dWOyRwGZe9r96Rg=
`protect END_PROTECTED
