`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C2pRhLZK5nPGotC0ThjB2aVD/NyBOXYyf59VCtoj+rE9
JxxjAJEAl9mRuLxdLvNHBpPDl9APbWXEqbmqviuKBZcfJ5LehWC+zVWkeEiUXqmo
2tCwoJPHOKCsIBHs3mVDSfLhpSHAJe4BB7LeYrwSI6MSV5hp1DSKacfs/MfjKFHl
hedjyBmS85K2SFp4B2hwEb6w2+9fxvY0Tgfqf555xtcNF37AP9gzTjtA0FhjTZ7k
kzs+aiOBOfsE8kILZ1IS2cyqsHp91X3lMbFI3DBsRP5QUNkkpvu09eLQbRjCNSDi
1pyHldP/2bOWKGZnwv6WyEH90RUqdVTgTRxnRGjZnx291rkVvX/mSkTcWAd4Rq7d
q9wB7CV5oTzxuEfDL6ak3b9srONFxhHzcYEYQoPBBhnve+A/GoQEMGZLgKvCbeAx
29+tJwdzAyUsPuhcM8ublgBRQABqtiWfLDPnEo7+hdbyLHYc9e6SZY6WhD0fP5u2
`protect END_PROTECTED
