`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFNG5FOGR3ZjYyXXhSL4UPaE7uRP4B81cdVX6d2lU6E8
QwjBic4uvynNPdASGnmP240ahh3NAQ7kRgdTHMv2Nc8hGk/T+n5cY8N+eEahQopW
vHzBsqf9uHGMCQCty4BKI9s+PfxZhbI4eUD7b8y+WyqD0U31wIumuH64vQyQI4qW
i2hTe+Y8aCMO4U1CM514ZU3HigrZN1YQCSydbp68UzD8+4bfYUbYjGwvpOfC5Osf
WkAnRwc3RLC2cmxCqxPO9up+VWAooNC6xrW37j4j7X4ELVvjbSb9HbBMgDAaKXZZ
IQlYx7NhvHH86ibxdDSwKWpJ6y4tCejh+5bLHfTCt2GHtZYlx5LzQxDLRD3Qy/k+
`protect END_PROTECTED
