`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL3V4yvll98zIkQaSsul9D/PGAk9tkoAB0te9Cku8Gia
wihjnp7NefkZCRJ/cbZHV/kJVEq+x53eLKxYQ+jw0GbRcqXHb3ZISjAAPcgKEF7O
+iaRRdAmnsJ4xlvbsOiVpQfYan7U6ii1XPTOAYErnhcMu7PzH0hBdIXQnIzaDalV
tDHhjrD9QuD71LeTZRUvXOnPpDZLYHvz5vWrRaLSIXtHGSWFR2Ib0TsdURfQjidn
ztJaO1o9HGawLSC6Jr8LCKCGD/1Q5sPg6QvohSES568P2lZXHnDjo5R80B/aHjAm
70DPQAYsQjAxwkP9SxSZ8A==
`protect END_PROTECTED
