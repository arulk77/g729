`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
9qWieJtKMByOne2AwkE3bKD0O1vQGi7TmKsdCgFU8HGhn980d4IxWAbahU1O7Dd2
tXutZw6iBN0YvvH792+m848c4S25HtWCQTvEPuBDlSb2k9PGCrcFVuTvhTxHJ6xD
KEwAUdpmBwgopQ7Puc3CktI+PHUc6VsJytmYX34zjyWOQ42ftw8tpQzFcTwysmVM
87a8VIoHMPXxZJVynKaldRJxhSvM0Ng4fV86uhmU/FRqilTiMKfYgFypcbS+NnIP
q37YqqBIwRn82an+bgGA0VdEx3rRRDUB9J1spNntnciLHD8Ov7737mzfCkPD9tIF
0lqLxi1HJq6pP5fplPVlEB+viFdUD+GHUC7/2wTIh3CUoc3WMFZ/oxKz58pdbE5U
EIgP4j0r9x6ABBl4/8tGIDDttfw4W7k81yOsVho3gQ4RWf6Pnvsj+Kt6bDetlnMd
kOQIFlL22+75XRNn6Pw9ZXTEa9gFjQjhFOrdrWA4LCVhYNoeD/nU+Nps3haNCGno
IIDoVVF/KEiroRbhg5yJrU2EzJAbpLTSdpDUhbCugHB8zqMUdl0u+dKUClnvq6Ay
YwBO3oMlb+J3upx+JdTC5eztXiZStPN0Ca3taF9n+rkaONm/rq7wf/COir90PHI8
cQxoqrjuivJWzqDjwxqGFc5d3iGvkQgNRvcNf7IEMdPn6r+E5cll7YABKoOXSzm+
IsdQugdPZobcsrzu/b1N0Yy9V1w1H37g7HwxL0RzJAHLcueHhGqI2T4icIiLGPZ2
ajXREJ9QTR8TINnaFt81vK447jhZRy9bYCu2KNSW+bxSyoJ63gBaPwFyNOL2phXJ
SYKYaNuLs5l9Rln/55GJRdgwvw4rJI4AOCOU41O9ny4UjCw8cJxlyiGUX4sVzyFg
2CmKq54i4MhGNTYpbDh79JL8Qte5ykIIqLIzFRKuWVBk1xVNvLT7KokoAMWniUr2
tamGtvIcAqYKF+/WixaLfGBblXEMhTnLFOwo2HM/IKedlylW2/3ysVUWHRAgF6M3
/JuyoaAJBDzgVqlYCBe+eZPoPrjB19BBTO1BrU2QvyL9LxIzN+nmMK1r26XxbgXC
UU9moVXPzh8fgoWsS5KObpZVfC54FcGKQ7B52ZTW4HFqtGF0x5FqVVVPnNouLdhJ
KnzG+a5C5m+I97cPZgYjtvBhMszN7KOe084Cu7wkzRl0gtZS9Dkv9OJeaVNoS2i1
k2SsiuADEGijGrG1yenu7qSKOr0pohZcFj7wJgNYHjQqMiQI8OXEm59q1jY3m017
EOCuC+oScvAV8ehhTWYL9TWZJeoIKGDKpkxMIKp3N4M6i1KsBCfyqTwtDsMow2R3
72UPGmHYXybOkLMi+8dGILEERRo5SAdR/Dd/Bvr6zyCEIhft4E17XVmLXQqhCnOh
HapkSHzeANIftsWRPQR9MYisAHkr1k6x1ZS7rueaKMJqKU1N+yRX64GijDQjZcHa
3JqM99kdrT+f1E2WqF8ryOTllHunYVfu7gW26xl3nQRKpDkfC4b9ct9LgCpqcyDA
66ZswVMxeIkJq+7GuXBZzAmh99GwzDsLWZ/MuDUjCt8i0bqwYhFf3NFiNdaIDY/h
uwpEWHAJ/9+MxcpsWUUMe+V2YsN7UYXRuHTUK838nUTd7vmdQ31QZcM+R/aIsdZF
aKKf+6kgah4hvLMa1megiuTNtycwHTAr4kF6hLMiAxYP9bPmMub5GvfwGcRL0yIW
PkEh8NzP0EaPeobjIAzZsfgHO4D4Bmk8fQM/4yb10wBN20DtpVX3W2Z5QWWNYoG9
AdLa+Mu/zq1TvrZl89OXTDsyeo+eVKh124qbz5Wk64piX4zhBDGWDXTW+NC0OXxk
lMk0+D/I1b4aOq6rHIijGvERa8t307vY4BAb/dKdVTAeWWaBT0u07sebGHwjeX6/
plxavOfvWN/u3JQzBKww3l9kNDC9+ynBU2OdfE3NeKEecZHRu6aZHdBdDH4TcGWS
52W8PnBygf/hXz02AVIE0/ijF9802i6vFtO7p6daIdeUb/TQHKK/hvwlDNfoS1oR
42QuTtoQaF2xzDZoXCRSBwphIYDo6MBhpAkZ1u/2dmJwx2DW/5KwuvKuroNqSS5n
xv0H2OTd+9hGUsyrdizqYeSI0Ob7fXJ976ta6n65Qq+oNED5kzUWbbXL80Z28mQ0
bUNIpNHi7A8tiTMf3Y17YtgG26OiPbAnKlM8GU0xluxydYSwIWKm5dDayM3kNY3y
kMY6kAI9cXcgLs9Cr/fINiAL6w5LnVv5WLSB2y9qK0V9hWJqkE0rv6X9JcN1d08W
bdNxUMcVtyC/Mz2IonlSiNoxAPSw191gRhjwAKviByuGMgVBsTd2Z62O9QsWg9bE
VD82U5Jj0N/LsJmL1Z65mZeJQ2oEDQP2QOwAUrthfrJxw76Sv1f4N3L/D1H5jkn/
D5Ds2XjPTi8QBC7Xs5zmqpoHsd6ybXiRDG2NE/7Z4BWi5FlY72DU5iws1+ckzr0O
teNg4Cob7T0T6F8N5i8CfXAKkrpup775MGIa0ZPAHAyNdcdXIy5h1YUnsl3nhwsS
xlnNW28c8OJSokBXdcIFE0cRyqCAkPm92znwzNpV0AQfzHLA6C4RcGIC3i4HjCIy
4DWVpnS9y8rExMKHQw7sct62/q9Z6ddSgSS7vXZt5OCXQcUrXi7KBbrGbWqvfRRF
Ep30AmqC82DP5L6wbQjBnP/8AQFnLBduysDtBb8Mcik=
`protect END_PROTECTED
