`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI6jSnuVCF7QCFxxNjW6r1wgyf8QgZkZjJ01EeYPbvjb
8sL6HJI77afBX0jr+PGHCEMhi/x0wZbxomVyzo+EdHwAfg2rqlDHzKyH56mo1s+B
+ctI4CSJFWzghz+ZTInqw0+eumNWh531iQi0FKQv2XUMhakDGJvaMrLeBBAmH9w3
X6C65j9UoH+JpV/kR/rDsOnox/JYzNDhBpTyMeI0gkAU3sgP38AvQTOKT0FWkm52
Vjb8p8OdkqMGNMdEZmfnP0iDWZqiMuCeqFYDdofNqXBUpoKyRY4PLJ4+6LW7TbBa
UomKAN4gcZqAl0G6pQXCTkj5HvlTd62CHwOoyABi2bevf/wBLOrsbFEZnklXYudx
d5vBLj8oUWWqYzjeVUsZ2kzJFtJjgh9hoW+95+jIl2wM2tpAzbSqVUDLCf5qO002
YVLxsCYnEOFNddPnD6Z51A==
`protect END_PROTECTED
