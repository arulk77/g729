`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOw/JvAtKSs7ln+bcmrZyM78jSJgTYjFnQrTxemRvqT2
y73z3FzZhhiszV638zloUfHXuF/m6U91s7DCCK4lT7Hl1be6BEBzIeTrjoQfRBVo
4EJvYF0jK/UBmuvxTiwDfOU6sy1ua3iGSZa1SQA7CzVcmHku1VrZYKr/2U/t3Z3C
B7+lqCYljHbkbNlvljCpjTxmtjTI1np3Wjct7Uce0KOpfbfplv522JwCt+JjIHTw
utKbJxKdJ5Rek0f06W1wLkTfb/3VlT5eF2sJ599Wb5Z+8mBD2OfwND6BrIGiGvUP
stIYfT3poVWBY9Ltz2UirlBWUoJTL0d6PTsc2vF9ugYsrpSO6RZv4hLtKCNAhcdl
s3f2Jp69c98ZbVDJQrMMnvpk+ho95FnXTTPMB4c/pzNLpjUJJoUcnxIEnNzhJvMg
jeS26K006MsPkVqc9Pd/bGCv/tSpTKcDE17gWjmttF1bmyOKzR9TG8WXwIlQoVGg
XNjJAa8o+xHiuPJ7yLq5SAwudRPGgKbDXXpYLyGlWdtefvYqqkZkxFaAhKz8oqu9
DFIjLjys7UvttpTICfCr6tPtoajawGBa3KokZVuzPsQ17iZHWZwjkvAfAqk8oa8Z
q/Ce10tsIEaqhTM8ejblkKOmUAa6hMAoVohUz0LWvqQPexiBePEwjL0TdR5JzhK6
xaBeJEqgUbKWEONqFt7hjP0iEsvD4xSpO8BNrYKOXek4X/lnWCdi/OxcySeiEiy4
BdW4QijxpC6vVHyD9yWt6YbtehhpneFOr9wj1G7XT8In3bgepNJ19nwVbFBC+R2d
cPDRoPpBwPJc1joXsWlAecvKKNmnoxzY0u/JACZgVkEo7n5djo7G/tm5iAVm7DWj
LbA5OWN0MUrKtL5o8zKJIeY+jAdDMnSXQdzZaIe0Rky0QqPXWBxLHZE7sL0cy9Az
llBKb4F24gHKyHVtUmfmkvbU7RQ0FrOOkbpYLHWGHFQKJhf7hHonfJqQkTgYlVw2
b71vpKBV63Giv8rkUg0IeYlEgMmNxohLixeOt1B0vGqvDrXX0aB2oLTVFri0l2ML
DUIWlotWfZNfwxk/L/P5z6ATZAl6/ayA2/miXxZ0QCig3nlfnBuY5PJFaS2rLifA
X0S4KwboxPLeIo5DSKUHhuK5yT4nTRy2xqu0HS3zar/eQ1DtASQB2jpqkuIkEJL5
QEt5YaOnWI8fUU8inN71yF5AEfbiOUdmQv7hmM5bjyiOO6QYzHRyvhpYYQUnS2ZR
/NpYNlf7+Qc3yv95UU5Ltwcro7oZhmNyAsh/dJ3TgvMq8KIwN9bX9hBJr+0cE2/G
ya+K/koGnvoA2uVaCdVtsN2tIhNOfvNX6Qe8WfPDGOAeKCfMTLMCTjD74jiPSmRb
KrZtrN4ldCPHBKcn9PwKDtGfBsZbzF7By43MQ3P6wTQyUpGgJqrU9G5BUAgPTzIi
3TacjnokzkJaOvdXeDr7lFERAiMUGbAIBLWY1sT6IhrtiX910W1kAs9vxJG92jLl
UnYGyfxB2bTkfEgb5J8qCk4A0IO/JO2CR5Oa/fIPvZXRFIZnZvZXtf0IyY7mb+b9
hKXtgIFfV+cp85h5IEhD9AjGudWm7Z4cWnA3Zp5JnNbeUtGR2qLz0CmwBW+MCr6o
r5kge60BezoU4B/BsvU9hfgatJQzDpmTDiTrLl78DEeZJaJprPh5ikdQA/2WTXhE
e4FNeESDLt/gxuMI2Usm/dR0M9s1OSvfkO7gP3PUyii9WzKFIv6mIhFXFx+u4SsM
zaa6V5SyY+OWa+vTWKIQVHsxgZCSP1ZkGZbXfZyd3CDPACNFsNaxXEBi+XOPsHWT
hFXhlG4l1tPYJ8MEif+vC1Ff9Te4mctfenHX0OdXbMiYPHP4ikfVoFyNM+tMNQO1
G1DyXdfwW6kihHce66eIQxMBhgqEAOiuQSVrUTLZB26Hmey2wvx9lJ0lH4jFeWS6
eGXJfbGdhi2xr/cq4QAUJoqJz+HsveX/vMM0L5VrXKgh5C0Mi9xKsfNWtTaNSIPV
4BdNfsxEHrKuUUyLHyo1ULXY1DWlSucU21GhFySEGJuSozjCDXjY9w960dhLJ5Wj
NxWpZEiVgQm3czW5TfrVZz5l7COwXW41R6DFrwjaEyFiLsmAhJr52hE+gMDFMjI7
hmVsqn7n2oOSJ6cisU/b+QCDFwZCx1xX9GYzsY9zydEaENGg6jTE0YFfXsjbCiah
kjkQ+ycYAqi2FDp59480LJ7EYnyNTUucunonQ3wmXU1jAgoGWPSb1NwxmlWu6I3j
1mOjePvyygp3IhsnxgaUsCbd4HWdDcf6cRn2EWINj2YXE98KyYuVGhoxAoq49pVy
QDY4ne2RWJgKRREy3Toyg9IcipVhF+I2FArbZQsBjRWdZ1iGMzziAIlJnNMVctvk
+yo8zbBxAo+JUrBwhVqXbIXO3C5WdWZ+2rilYDaAoZQF/WjK2tXDMgac9fUX+oTz
iXuBmgXunVV7FN6S1gn+0u8X9GjCf42DgLwD9D7S1qJ3TegRqEKUM9tmqvIjIVRa
Io2KpI+H27Tv83SQiLBr1bDpagKisqhhSzL1kGEmgKhn6pK8WUeU/TwKLrEmFztF
JQZwc87mqr4+t1+3vihIclmyxjAAUNEZN4ZuiMTgWoVd1pGEk6hkpDvRx0+l7lWq
IGLk9jDrSetgiexF66Hi5V3zPmvAVEXqXbPGHLBKPVJJXjSCuyFA7J8Qz8iqsr+0
/6WhaTkO6CIlbIV5ldHuRS/N7MWTIjgcDy6V8IoCAiLr1dbUtJhvrpVbvlqfRza4
T/n7dKz3NqPwWmsefn/NioT3wVaa0orSr7/pvec5WGSPp2PnMN46oiA2ffHW+COm
LBFZ39y0ylfzz9NWcrf/vXbYid8b6Yy/Ctwl33BG84jALMXq5PkypCJXx2mTly/L
fHomoUyn88VV/BWMjLQfxxBi75SSm9tX4jZDs0nzT8XC1XJ+7zaxo7ga9Ddadvmu
IAPbhzkkQ+ng4b9Hgnj429T0ZKHLbqMjk32FEDIEsTwykuIPch+gJfTU81d3yfeJ
nEMsuWhU86dKgte3mzSTlnbPrUQiq1ok9rYPenBWftaqcbQu1cb8aTACu3LmNlf1
mQh1RwcEcDwqMlZVfmmlnb2g+NjOKjs+SLMbHZw9VqQbYTEArYoYry3/gS68qh+R
A787/yudByJB3QSeT2wCtkf87j8gfT8pqg2mGxWghJbwoqgGw7WbzN/HxaX/rEAb
nNLijj2Khl8uCHynaxMUrHWRvYQGoqbonjPD+QbQLK9SLe86If3ooEyoCuCFI19S
sGs1MWVzuFFk+Pr/Q+up4jGou2thWzQVM4EuZ7R3JHeLzqfZJnxVLb0PanthoB7E
olJYOV8KN5Kk/uGE3oz/3+zHsPFsTRjmM5ZXamo4lK5qcDXZ60QFXgPO92xc8DWZ
apVDlvFgzV/hAx+d+YAPBoHame1J7EGMEYHl/YpO57BDjVdBErppWDqPU5uNiJbK
gTYTt08RSs8bQ1sTNlwvf/cr0InVlL+HGwB0y1cDYtZF0hBkf5ZnCC9Qc8RdOQ+S
2g3FR6uDbR/VtJ1TirG5PSKuvykCo9pP022AHvDj21VOXwBomMrz6pd9ka0/XSJl
RKdA27YL9gx1urJxQWVodU8sSPXscl1kElF/Ti89p1aPJasCI+dugghhd3vw631D
QSDsmrWLQ314RzN3nnm52woUr8XO+iLT3OavrD4AImAh5Cp3ACinQjfeF3H8kPao
hTTrderjEy+QMFhCorlngKwnDg5Atawb7OyXMRWsbTz+20v0lIn/6ePd7aD5sbf4
Bo7Mzn8Lotc1ahdixK8WD6M38BvJU5IwKsoqBlQwS48cRSMdDI7uA3g+Cy1l/NwL
vNqZZfcM2WPw9Q10GoRuyU6rzicwfjSGE7OGHiy8rp+sssm16PDURlA8UScG9Hgo
12zk82dvrarOkE4YnYFSxZOOjGpF3BEWRn5U0PTxo3WCTJXbZaWMkYtQOt47EQph
TYPuG6JGRCCM+9XeazuocKTJySc4ZoN2jlZ0oDoILqeJHkDtAWO9+iYApJ1LX3Iz
f89luw5zsI5KvexJOSi6MiKWj2FAPKpnsXOnBnn/pE1idwd+FwymFiUe9ZA/Bgh7
ZIgQxJDirBpsv7jyXxgw+u2qYQsRhtEn51Bhk4Xtz7/odV/b32aUXj/TDwX4vbQK
y6v9JX2ftDovp6hI6doB1HLSP1xezIcR7HwD2xpep2pWU/J2137Kfcg5wbfufuXi
dKhwG+1wnHbdjtDb91rWsIH2VMjgefmxYMGQOy/j1aV4NdQ6rEh556m8oR8puokE
z2RRUfdSQrhXeBuftHglrvrHINNfZpH3za84xSUTYKgEP3X80dJTOjKw5RD0kaHn
ipDx/oYDBaRUyyqUln7fAVDKw7yrjL1nk7hzpaMXk6orWjeMADFB/VSZyCiQjVoD
upuOg5YetxoaN6D1as/anWqhZr1kkOu+VFpeTKwT5aZpp1eOQHoOSu0H3phbCLZr
03shLblTWxJg0VBRJBYpMoy16h82u3rtshVMjlzGogTJ6cvH721DWf7SOUkyQ6Q8
W2x/BFyZwNcq0JyBFWeP8kATm5LMtbKqb/081qW1XyjE+qSrYLal9CiVjyGMUfFD
EaEymlNQz2ITPhaf/3rxe8LcKtFOXd/6CO0VGQWji4D1CstSeC8dwwF5FhbfX7uQ
FTWUqFfFfxIUOkiUCB8NYNCB5qb0QgcDcHza9OrV/UbxvEg9l9ZHVBCPeMeQEXLD
ny+Jq7SGC5m145NGhLZOhJfBXPcDwlP12JBG8dW/QXr7gWZEnUbN6wLK08/RdP2d
WKanhxbVEGp8akqXbm+7YRv8QR4xAO4gH2WP999aFV3B3nyM+rTHWNTYYC24lMv+
+2y5Eg9PCEYQb/jeXxXguE9jhjyfxvUc37hU7On6Yo+hg27CIRaie3WIshb/skhv
9x87mNSRxNzgEgWb1VvuD6fZFl1a8NMhfZ1Kw9XsJkH2DMu2uKeA0LzOjCmi02SG
OSMGPQ1iGhQiF5xd7rZylkER+9DL0PhPVq4vHh/iuWUdGpZ804LVWgfXiOkeGZez
ohtWoNn3AXRid8EY7RnUdr3dOtJouGc36EGZYbKF85PkglHUSzPC6sh2f2dSd1NT
SyVNxcVLwCKYGwJTZjLCXCCHDd9N0IKIPxF16mR0lj9+R7V9+6+mgpMRjn6cmu2i
S87u7d4fLZHOOvS7ds9o8RRp+VuAVuHpslcKM4S5Og8MOgvf61yY/ZwwH1WrkYrt
EbFjOu7Mk6uR7vgZ5BCd956TU4IJeyQ1U9dLiqDNtNuTjdTGXQF8zOzNXdE0tPE6
MHpRn43VrJ2IsrUN3a7mdJUehBnTQ3266Bh6KZQQ+1851Yevje59sUQivPi6zpbX
6comwIPatKsP4Ez3YNR5CLlZRQwmQuipBO+GIBjpcswSwwFvLcou0dgcqYnn2xuD
BXrQr2wd7c1yG6cmnxH3e4iUbXDkhxwc+j2+j574j5GVqxDJl3Fism27tpMdJ8A0
SA0MNXYJEleWPqNrbCBT+4ZJ3M0vLcwkxaeolRdJP8smQZJzTwGh9GJ3+L5tOmpk
EDR1bPaPHiDhJtYVEnGK9dHglFuk7CJ4i/8UxBzG3U+A5yVgnQx1aIN27s4S0gLb
DFrY3JpYwKGSYr1jt2gcKh5CvPyGbmtELQYqyCf61wTZdYD3AAwlsiUZFv87/HDm
SRdeXlTY4Ahvgak3wuwwgg6fcl4L/EWxzRimSE5tbB/qOVkkMrYZT+RCiQaK2hqr
xH5TJl0C3luu2MqcDpKNRZexaTR68Z/k70CVQl3TtDvxdqP/wuFYQhmXx6xt67Ab
xnzBvLOfXXaEPPGYPOOOucY5dKDOmNNREa7bqLwVExSWsLpObKZq6mzZ7ENIKyI1
SPvkA1G9xqPE5wBMw7iO3+h4Y1sV/bg/xG5U9pZOwS8sJVwi2597UhWhyQNRKBpO
q3D5IEYfAr0VK22FR6ij6fqe9L9DjPDwd6yO5mYf1XSt82AMfV44Vx5qvVlSKkve
ZRPyuaIdqZYpNiY0dYAXco7rb7pACOHR1B5HfRUAoaJtA05iFJJy//ykazp2r5wf
FGpi/wF/3NoBDdpdvTm0IQhugpVPBUT5r7uaknx9cBnhTNnHVAleNZAZ/F7moN+c
PwJrg8bUsE4efhNShMzoCQAjrxSp4kDijRdi1QAyv/dsxSHFhfKv5b5GusbPcVb+
w/XHg1rJv6bZi8LgP/ksXlquNY5Og/5Nz1Jweoaor3zhWJ0CYPEI268mp31XcVra
x0mnTq7LQfnlO4R0WZrSNDBhOVxmtYgSczt8ZzJXouv2V41xo4eC5uhS70C0aB3h
RZHkih5AsGzySkpZHLPZuw7USa43IPxOWUTiCtzu3pGUM98GZnLpmQfISDFMJqMG
tTLgo1ee0ruzTUVIblUgSCLOh8stDybz+29StcopW05B8eqvtzyGvNXfS8KjhVDZ
UflZlkHDXZMtYup1POC7yv9yJmLoodO21M4xynYDMqITNX+rmoKrmgn+s9oOZpcI
0sS0HydWR1hFTAEQsv0ztt8HnRx25kZUmMqM7Qj2y/Wowl8HvoqU6ykuuc74GVDV
uWQhqRvQi5cW/Ee6cp0EkZrT6fzikaVhHP/DS5vbPJ6/ianW2l5Ulc66pbHTzsNa
R+JCbT053sf8J0XGcT1g+9vdGY++sE8hbEfbQVau/GPghR6PvZHIkr6kvRegsvRF
ULaX2gevH1ocqJrqaplW+dIbGpNHK99HTCRQSQUzgjy14W43qJGhlEKURxvpDau+
tdgTpFH7XfGVeN+7zfqpFVk+lqtkPVGj5pAxtH8dOMyQUiOSNY+LObJqrNYkqEqG
1S0V4gOF93bPDO5NFfLLs4l+8O6sivIJCCcmDOUclxHi7sDSUOaWR7WJa63+Dspq
CiWm6NhQFNbyaY/g0NtF8vaSDDBome9ADID9PPZhxs5iKFZJ7OAUiVpfOwY4eoe9
weD9T+qkN2uRioLZjWbvfwAQ0WuXGaqryL9Ckkzdh2xioEbHy/QmcMqQ3HrKnf6l
Bs7m3sr/FxoNpOrptji28xGGRhwBwhW3GQngywiogN85us6RsvAw/0u72E2Jlc9j
IkAZcgHW8A1D/KXX3GBQaiONhhqOQhC3BAi5AO5Wf949+wSXYE+pQXPKhNowEl2I
JmC3BbqV/K7E96uH58xedPA46zCIa/SupAHACao9Ihp1t9SGoIGCJAym9APCyBpE
g1EEGejwK8ZxXUFJGBzVZl0Uw5M5wZy93Yj6VDbvyB1zg9jGhNY0i7+lAR8WCbUO
XEs1GMRV0ZK2Jk8RhUvKiJUcjyywxHP8ZNL2RYs7ilNg0T8vaAzcP3D23N6YuY9G
ncaJBvQN+EOMRlygZYxTV0B8fuBVZromEkveUel4vlT7kCq5lVARA4tG9xBBa9lU
SxZL6T9YHQhzIllvWMFQYuazVuWo4UeBZYat3ALGvkhwzLHAK1UxdwOGtxdntpno
maLj9vN6ZlysvH0eXu6lgoCDjLY8N4VOiZAjtkOOnxHbx8Fzg0OQ8NsKMGDPxQ2g
SBq3m1zQAhDJrjcJPVnMijXIScyqx2V5KIRHZPYC6AojkDVp0ruCKvpe3xWFxhf/
J5N1zqWbNdzhpVJFNSGl1UTY930568n08bx83IUgMDZFf9ukdWgUHY7SFF6TOhD6
lexrGHjvhDt1HqFOteWdf6scCVw/hvQBZho8Vk7pyE2avt5pHy0NqcgZlw6pIj8T
SROf3cyj1N5T41/r5Bf9mioNnKU/DyOb7VtN3B8zsWNbdxULxKlouzIYTtkkHMme
3EUxwcDczjLoNbkAQNNR71AWQQdaPSLB9fvUndIl4nay3mf2GSzYJuNdfXPKBk1s
At62g/Y7MEWQS6TEmxq7/GeaG46rO7/zHIwtvQiSt47/3ebXTXglnlKababPlrNb
du9fHh/bNsB4yYKj0/3npXvuDoZWVzci2NXVJIQ5/wCKa3zLdo7z4jZwB4Iwqd6O
MOr81jtEkzXGFGs+MGljnSrBPK7qQ7hbrkLvAHzwrbJj0CYwkJ6dcr2OvnpmURsv
QD/ZM+bJnCEHkWK1Mk1DD7wdmHnZMC1Lm/Rh3BjYZQi80Z88sKSQkthJaMqfbGYv
W7dqMLMY+anIGivLM5wIPcuY049jgqilP4KJEPZ/jXE4TOr60gTDx8v/eFGyHVzW
UprP634mNudw26QeQS3KVYiQByASShVT6dSyl8TLjhJiBnrMTLwZo/II+3xwUQCD
/1j05N2rebUMURqrdYtrBIzGpS4J7llL+DbnFMSuJ0s82tVrJDs+YhNmg6ecHf+B
ZmBjtZU3EE5IGcfdBwA2cgjtPEjLY80Xky6bsTl0b8z6TlFbM+NAnYy35CQAdajL
kMYxCu3K+Wg8ikkN2PtovRJT2v+Qu17K4wu2u57EoL8gHPMAQXqPobgCht1+Dnou
bn2MH+O+FR5qs95jSL5NIKEZXLCbuOvkX0wtC+N7KVvh/xsMuo232CUg64yW1xWu
FRtmqPYzaSu/MViLiX7k2jqtl3LcuRCSvkJEOz3zQnrewK/Yz6KBBpDRQOIG7ctb
6rlHLxH3SOSUD3tnqO05rA/sZKmcjWcJ796w1RU5OOssa+TrZUmoEqRGAXI4da9J
JA/itTq33RB+WZ/oKdbOI8gwGj67MM9TLj8wXLRDmSlhfdwgCP89Az0Ctol/Q037
a8ljkRWcW03P5P/d04QOYp+QCgDuF5wHs1jSdZJe1TmI2rOWvcIaHqPZ70KdTwCF
KvDSS1yUnLcPtmHIOW80oLeCzixz/BC1Mv5BYIWBK5oyiybPUkomu5G5xnrsB/Xl
w2RWkCvVUMqoRK83pww+U6Wv0qHP+7f6KwVRkTM8EaHODvSv0AD5Tk+jXFE1tZxT
yC9VGMGxoKCr+k1KScRyVsIbaGYmHFhnNPrqa0TjSkY7OyZ6C+w0WqLRf12FBT0u
Kf71LUNARSosczNpBx94g9uioaSe93SdpkYBEPKyMmVmnib3H6eqYS9KwoAtP0st
DWvt49f/7kJ9eEwpUYMrvSbMVYeTsAco1v3TuJRnwu4SDwuGK77UKOkj73Ibt3HC
JEJaJ421YbQFBCjhqAM8bA4x+4pkbZNny8Xn5AywYPwThVQMN5sjxkdPLtxCmqOt
6RjfbBhonmc6xcFj7K7Wfip2N60dL8fqJYhioPHDCeDzbhk2Day3sN6yH//UHY7y
gLyV/2rH32Tr5AbD+IfRUru926aRgrbgUVcfYmqnshN+XJCuOKjkRCBx5tsFKIst
pC9BpezDJMK2lHg6K43EaR0p33K0Qzh+p44J2lMiC430OETOObNcEidtWxCMssYP
TEzxAnqS/5bZetyQlek6/9Cp508OMX+mTZkMsghcrqQaHisej348UmOToXvUtYHY
DhIq/rkyU6pB7UzME8cHea1nxas3VPb0E0l0pHmQU4BW/JJ2u0S71FhXnXSxQ8eN
PMuOQjiZr5KYUuqlu2WiqZpsC6bIgj7OpcrjsaxEzJbobX4xd/ww2C29CEd52rtH
tTgHyQ84g9uw71WzWDagr2pg/TXa89Yf2UXFEEGvrDY1Cgfr9FnV2XITRPj6Cg7C
H/MStCOLHhkqrDqxEh734EEZ45aobTFGjU4u8XZJuilYufRpxzK2PcyJxG4jNzsz
+4FHXtcM/c0B3g+MdqoL+Z/1K59tesC7+YswuZmoGQScDuVxgZzai7xk+DEOA3yh
lV6rhhVylbvEQBTop3+yB6ESn+EOeR7x+fNQ6Ruw/BjzVzL4MuvyZ9Y6yio7wt7B
`protect END_PROTECTED
