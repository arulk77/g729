`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveC4hHRTqvBIGqPoNspVD1ON6Ig3M0LX5l4Za/R0nMnaQ
skxGu8LQplHDqOBvJNQuBgcE4KAxWnleddCFmMBI5UBbPbIsCRVvt4G98KWZfgsh
HBGHFv+6++++4kd6MsOc94xa7nhCzzIk5wxDP12D4qChsm82zcYsX+ssHJBcmjQX
4L/MCPcXciuD/PzIaukdxQ==
`protect END_PROTECTED
