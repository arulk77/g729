`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHt9EJ9jNsbKKcXvssEtgd3RrpcIisb36m207vBfof8B
m+eRBqCYrWtLITr9LOwptbBfqIjC+RF6LFqj+09bYE7h+S7kf0DFDiaMH4yqxHHQ
ZQqBnZBSAjg5M+tcFg4WLRCdAJZiViL++GStgfjdOSMzNQQLIvqf7qrJFfEIhHEh
gIQwJ/HqL4OV8VVk8D/i9PItftGik08uSpc9pbqJSN+5svcNvhKTJXIIfP7Q+qSz
AHzrVvhJ+amNxLMef0uaxA==
`protect END_PROTECTED
