`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C/8IcxtvcGRiKvGL/F++2BQHw1tEPyN2J/faF8ZJOpdV
u0ygHmMbbwv+RVWOVSJDNdYruRhSW1FchhRq2JjK2yByFwjkWCiXullZLrnPj/XW
UOuddmFu7axh08Ss2/hJ/A==
`protect END_PROTECTED
