`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFVM/SYqRIJvCJvwJfpFIca42DU5zuljYorQZzq1Ucup
nOr55ZLRKLkNzb2GhpoDxgKiULa/oBTK+UdTAkKQKDJNMXDQYjGZD+ZfoiUkOAdz
JaWRlVMwljA69AYfc1f3EC89+CIJP2aiXTZtfYGA4X6if7Ohup1m4xM4NwQR0SsW
qyaOjHhMb5uEbqINvlFFjnJjtYlVPKkfq/NBXN9xsIuKhNqezApkZkaiyN8rct+n
`protect END_PROTECTED
