`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/ryrNx5MMXksya/M9Ep6DvKs8x3JE1NS8Jcgq+lAkXy
zAHh1Kr2FY4mSwj++3DKSlxCnWGBlGfTsZ2CK7l8rIc+f6d3CkLDNjAl8gHZFcdb
QArCuwAFaZnOKkSNPU1NrPi+02wJT4ajTuWBI9Bfmq8BDa4OIb3z4jdPXaipyyxn
YDaYAWbl+pZXAuKRRTmoY+bGueAB27X47vglsTLJhOvhmL/S1VElhi/QdW/t3qyg
EKVzh4jEeJlc0u10jbMnAazDsJINxljS4fwPClT3wzvsyf+SHwbO/7fC6xijd8r3
b+0yZYxu4oL+MH3H8o5hacvEp2hNBIEUtnwlHw/xjXson97ELnjAQ2GsVHqxk1kj
EIVWM/dmte4Qs+5rgVeLQwKCmrLUs3n3Lxoh9Mbd+NN8K5KzB6qgjlImk9dfSP1N
z7hF8G7gK5bfC73DAQ/ADqO/Hl+BXutWJ7oETZ7N07Q4ogM1cv2knoQZ8uvU14O1
`protect END_PROTECTED
