`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNJcPksKgF+6aRz/AeFmGjcOS3t9+7dQdAbACOtYbw34
fgDACDt9zCNKjcQil+pao9vIqPFGJgbRMc6nYXnU7aWiD7TyFhQiLIoXUCPO4+IF
jUkqFx6m93QJkuGHefr8YcVHliq0viPOu9lbXo0Lap8piN6KLJTMbqpqwUWwiq9G
PNcPTzi1S52hV1tC+tI7OCyvrxzmJ0WWeM3i/+1OkjByewUeG2/daWE9OpNzFvD/
XSNS7H3sRyrpK2OgKdfKVIAgA821OGUHRqGIUO/Zb52fkLnqapLyrpnu79uQ2U5D
aJkfi8AQnP/q5IX4gzcwJsW8zJ9f6dManBlWGdnmEVuwbKIWAF+dyuJr9CR052cN
eY1Pvb2seNy10ldFO8RZRyGGTpxlmWqmoPptHvJb1bZP/BW6NEp74g3+4ztyueoY
fNeyZHzisf61xqkXw1IoDidzfqCn/tfXg53CAKW7cd+b0DxI84lcIXT7WgMoUTtv
l0/WD9Wfi0TM0tUBbfl6fAHzTUbjFATsa/w+D0pZHcG6Wn9KblWWdBeuKv2RpI6I
Od5dhwboPyFwxnxTtws+SFSkj6yU8RnXBnyAyRg87BMwrwgsvn4NnwXwUHTq3M9g
nfBI/4mfdyBPvN+ln8Kxi/eA3IHiWmTKC0KUNS2WQCboKd5O1pQk/Yz0bGA+DKlC
2sPgvVXX8jnMmgzs3/QZu497iTb2XUxLi2CAYGUe/lm3f5DIq4M4MiqgnOsHBNUS
`protect END_PROTECTED
