`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1abdplqALTQJk/JgvERdxs03TmDOERMv79hq7pRHQr7Uc
PJU8bg8QqNbv2wniqVrZNb3Qcxk3mVTRqNoT9FVXqI/z+JvBJ4LuD9UchgiQ0hli
IPqIdNcWR3ZfJ6odn7dn07HkEJghOS9SmgM3OpolAxHjG4SEJ+XkMwjg8spe33Xg
QyGLJUD1h8bjKBsoM/7jTZlnxoVhP2XTnRNiCxdet4QOB09O797HOFBrMv7iP1do
SeJgwJRxpxAa6GV3pEpJYfs9yUAzhnupaUaUkdgjUJ88AbxYGVKUyrlGOovy96Sr
499CquC2xRFDb0Jgq03v2zSB4r3TdYA4F/EwZdJ7nDVOSJUc2IEMDL2oJmzJJQPR
zNsPgSp51O1dXEEou1RCVTSGTcpvbdq44rCElaTdi8hvk3rt0kD4CvrW4VN9FPWG
kV4M1BOxeUntFxlGv4hpEmHVAmPnk0FvZFF/Zu39Xz12P1GupFNScfIDca3goXgZ
T6bITivtuR6jtTUAbii+mtR2qf5HM2CQe/BFBMGvhXm55HWgfBDMg8I5qIbkIGAq
JyLitBqYkPHzdKochx02dFBCZnL8wUStOIKr5U9qAfoKZCfcd5QCli+g9+7uFz51
JmIWnuWqk6N9970OV7iHHPxyqjHTZrl5m96OCCKy3m0RHb7ObbaWYlckYUeInWlN
FZ8ziwB838FC/uL99dHHepSesaZszU2LWO2HdtrOgGIEeHCtN6RZ71VayMjCkwaq
yJPEFG98AfgnnWrpGCj9tpGMHL/sj6GdnM6zlo07CQw9Omv3jmuhMoivOoqcANCL
Oc49BPuivDyBrowScEJg+mbjz7weckJARtvtbboOOIjy66B7JYiqQVa5HvaWfs2n
EGGcgY/X83TIefGy2gUeD9aGdQrG1a0kz3T6HKVc0l4X+jriwRnOUujep990JYJ0
J580AMaMdILa4oX5FyNo0bX7XCl4buNthatbcABQv3u6kRpw4zPAr2puG2erfo6I
D+z8o85GHTyvEWFbBtQz3TpPnUQU9RhYMtcKuYGguK1u/SEtubDavlCH+GCdRdXs
SLTyfUBFDJJ5P78L/sSHpb4FgelA94FLh7TPxbfldzGK6Iqssrp/zbB0V0PNRh5R
z0L2KYjsUd+1d7IBENzSyNHgU6dEWaGbsv1kR19YzuSIaEsbebFS0Bv1jC7Dy1U2
WHwZfQTEboVtAMeXeANEda+sag3TpVz4C7YByWnJ093YoVFL2i/VTJvspD/4GLdT
UE2XH7ucHin3kljgkLpUZ5dyJdlGbipSrs1/8cexZR5bvu0S66TP4kBW+YZUeMCz
aV1+WvfUyRfBTvwKC73I8l/Z7cPzqJOJ3b7cDYAahd45ERIbfjlyDmannJD4V9w2
rYc3Dy2SCegqHx8hZENkcY/GstxirVm10GXfZu5xomGSby81g88Xjs8tnMotNsRp
kcRnaDPFmxCF/LiaM1rRy98zpxKfy3bU4/1L5o81qXe2llbG+XyFXeHqFsAH1pDM
DINyOSg5XtsWBSsEWZmMBTuo0sh5CdSwOT7f37VQh91SQaDHvLgk7M1uh+D+eWq3
6SYil2MeheJpTqyfpQOPYaNytGS+ookJL+vpYhrSGX1+UIU5OoVwPQ4bS9EmJ6Ga
D07by28ShfiOQTzoOqafEoOLPCm6/FFaNFs1KXHVqs4HQWr8DrGRIiEfpdlEB8xn
iBwvHtRveCtkhEjemg+jIL7kOSnOrgdZhSIIO+hCvLu55QZO1chjYS/Wdvlf81ha
kw54MkPtjsGOSS+GihSfvlGQ0imiXNuEQ/fp7cJ9DhBuNVJggweUmVM6TcrMbZyH
NzuO/eZbudGbMecgIz4GvZ+rkzHHaw5JOCnyy1m6bQi0SWf60rY29gE1d753Twa5
raJ7Bn3F4iTo2qnmPkVRhG1acI+Mm12WWm+e/lEbATOnxTgMvaQwiDjwUVUcJuB4
9+Qjcp1Od9cNmbuEhV+7OW/L5Vg/HcTUsGOKjQjKJGDGV9cH47ki7FIR0ic3KqTc
+gDZO8Dt0Q7BpOyrSQt2a+xl1FpfKqgaiDZquEBFTvh7N8vvu02pCG8ibja3nUih
ReRNqsE+gnCb1dAR1dBE5Y42a0OivkzKk1DYWx7inZtTaWgxYrUEnWFqcepq4Cd5
KPrHIQQnKqsKTRj6bW9x0i18bU63NqQdhXxppO2t8M4CQ/lVXYoZsIjqtWaDvPVa
o7oXA9FlpIwd19mFYIv77SG2yjfcOhD8YOSrV+3nFJADQwiv2VrEohQoc3AdCsxt
/Sya0R2OjpWOnAZmXzMIUruW6F0IC0swlOo0h9UVw/8dbyL4rDHXsUc0LVPJIWvV
L/FNXUcFNwO8vuF76EQeYZp0CENoGAAIbvJwui7MGUta3fj6QnPFfXiOqpR18Zfz
RqrirZ/fx5zdIMRctEj9MYOYkBWmMOvlGux3SPH7zbbcbdRQqNBWJvMJThxylHVD
SfpHyKO2IrJvkR3VzhjyU1RlUM+uDx8Dq/ciGUb7ebpLxCMhSdeCxzer74vSgLEL
PR2UxBioU8T2OM6aAIeLhZbn9MwD41R/qoNntOy8A5wDhEJ7qCJMNWlt+Z/ty4lR
H5v/hrCQk+LK/HwSwmwQwZxk0eS4Pu5ILJvv7dFDVuFP0Kkke7n888RniY1ZNurO
kqM4hIwRB0N3fC+S3uooDKOgpGlwUSNiDpEv5SugXziQUh40tWjqMa54kHEE3KGc
pXQFC/sF+GH59Adfkm7pz6kN2AG5Q2y43hjz7RY9oJH/F09fwPA9fjtw4BpCYWCl
QNm1LY8tDG6SdG7z0bLb4gDDSXvH1LsmFnOAyiMLq/1932CMS7YLbm+0VruNJVQ2
UBX9q/HiZP85gCCSUhbr+GK7Ly3pumnkRiO9uxciO/gGv5sB0ZhIwBRl6LCfscCP
3yGjA/IRUFlGJocfkDO/eEHf7LIougH4dPzTM2+NgsalHDj3C0xPz7UsKpWnVfDA
/8VRhJcm05Zexatgi/O2MN1Bzr/fr3JmLvpBviosZqCUQ/XDMNPBpQ8aF7h8C91Y
+jDivGg4Y0z0FLcVo+2TrnUuoBkMwBkQUhO7rsNTBdyvOBJb/gWp9aDMkVhg22mZ
J6WpKnVIJkEpT27nJajvrrruoguGprrJPhb181QzS/qY+Dpx529ZhSuJxtdn9S/O
3rTPO5LEaOXmBQoiIcS72khPWuClLxsWxlzDWpPFIf59ItIj3n961bbxmHKJqHEf
j3wqxHrlqMV+qM+Ig7Tg4bhSBhNe3MwRcx81QFtQMChwUjDHTAS+a90r6eEqgYU/
UC8HiFG1pQMn8YvLUSswFxKUC9J5iUuUYY5kwaCFrSzpHVok0XIDpv4GfVeT9gD7
6QPJXfdtU7aqzflaDzfG94buwH/zD2dBTYgRYNnkpv58IFMIhmGGoLTFcRrVgExM
Gk2xRAt3YYa3MAlVn9CVX/YnLIlq38NrCS0rzc/AMWd4wcimpNeH1Sh77TJ1pCjr
3nbDiMeiRPP7Fr2+yz0jpqXw4UHxyJ2Cvnoq3afiVrE7AapxCoKvjYPbT1Wv9Z2v
aFfEBA4jMwqr6XHMfg5cuhPeTFqezx83h3gIwyM4rSqLFEpITsYGmArjyqSsSCbA
Jc+1OB3pZ0Wu18ePO6trBOytV8zPH/ZRhASfF28kxwkcShAjMe13hvN8zJNufm9j
sPEbHgjDTCZJhsSKHM7wbmcs6pjvaxcejcljw5xnNIh0HvS6BRrg81yolwx+ujyA
Swm5CFe0uJ8+JvzzAAW17ZWnl7Jt0nkgmTSnpOqcd1tkEnnwvEm1HNtRBnreh8zr
qPLHAljjLwsulxlIrYlrvxf78FgJaxqJc47uwHuHsRcT7kCwbyrq1IVq8AJEXIkS
1EV9S/1pkmcu7HzWSIKu1fZiavpf75pH37nZnHQGDDRgb27bWCTfoE9EhphgSzyT
j9z4+nAddhQ2H1WchrPwIobvZ4roLaBc9+D3bubjcmWzA9CSXZS4WWRx2sg8Oqnk
zRZy7YFOQbb1KQBRm2JD9HegkVEyFYd0qBAgFBmTf4xXtherNfg5fX/CxL0OqmBG
faoETwSqGkuoaaQFhc/bp2nhTEyhGncjdV4YaJmsUA1Vg2vvnOmvnzLky02inMWw
pVpBuCVLtJnz8obSYS19P1pDXxQV062yeP68+sPYdDWqK/u64IonLqxE7xYyOikY
GAfMKFFQWmQO6Mn9keN4ZjXbJ+rCykFUUWhJNbQeRU+XBE+s1pigUJdidpr61Arb
2CBFLqc8p1LTTxxsTzn3siO4/3GKCxiPKK4X2rfdfqSTVGDQYW7syNg4RuYzhYLD
QlPb0yXtOIjJBkzPNsMuKAcFyOsMu5IU0++PTA6kG6v7vpB7tGMO2y/uH5xJYELZ
Phym/Q3QyqgnjFMM9syjmi6Zf3wgiVP4B4lM7x1oHyp9PzsO6wb3LEyUXTfaRdZa
Ii6PBhinaczBg2Jtram2A4iFHCGJ1O05XeYcylmK04EBWqKU9VcuLETInp2o/fPW
nXJtrFX3c93YVLfMYphLXOQJtvy0xr5ZpQks+vXrqU9DgCD0e0Vo1LKRYL6hPmIG
vUVwqI7f9m3okrsJ+v8oD4zroheP5CfdUacz7kfEdWv0sxKKZ/as7diKe+JlyQ0v
n6CRJ9w5rfLhmZaTiQX8GB8PvTJzMG7JGPAD60EVsIZ4VS9VSTE7P3L0e8FW6IxV
cxs4c7G0YW+B8EtaaUQkjnt0lbvO4Oi+sd7/mt5HnHHcMHhuL4pU4F395bkDqKTf
FXys0Y2cBnV9cN2YAuEe4xRarwRI+jtYQOcUSmvTefe2MMAUdQoPofjo/7hvR1ct
ULnqAstrthVOZCe/BOE8SRMZSm22Za32OI47F0M8W0sQi8gkSO8VoPnR3jkHtv3e
q9iUUWjzQ2BNRUkVbIFcIlvGgnw+8dH0DD0H9S+ghLOocwuS0/QuFc6jm3Ks3LgY
2YWpxP3K6mMZl1K0PMJn8fUxdJTlAHRdjkXKtgAk0Txgt77CxA6WrcF8/3AhX91p
bRReqf2R0xtDi5uVbqKapnSa/xTt/iYHc0/OxKc8hIMUnJb+EvUiZNHyZrKvlOQc
pqIOnWbLVabRddya3jYFha7ugRTHKNIxeofkYpCLkG7Aq+M0G7GTwyUGQ3eUUkDm
10Mhx3zYa9QKwQmerv2y6ZgUwRW+E7xchRt2YteDEOnFYnu+vJRXb1iEi1l1DSXs
+P87cg8jh91IQovnST5DSQD3HOVZAfkP1x+wia1sRrnYub/mGgBGy4SCdvW21FmT
sIzWAu1w9QrMzOs3hT0t9IGUujITwXHpgEC4oI2zBnOgsWsHPdTXla4EJRnd28WQ
LXNWllb34jpK1GY2G/JUMLixSMryqKdnomZhu/4ruB8bkuOqO01yJGrES4dgnOoI
DeYVBgQavXpWYwWXSbUSu6RXrnRqCn057MC0metakwSgXRlLEkO+hVm4wTYen5YK
j7FOD4tG1Y6iMyB2v10UUlc/P25norhQDKpuf+5JXolo+2X+EBHu9xSPOYtORLZS
x9eREShrG844lcDmbWBAwTtgm2FvrSH4cFXdK+g0tTk5OPRy8W/wjnO+LhIPV/CG
7M6/3xEDlQArRQRa+AsV4vk3qJhcbFoOg2UoBehwZUYzoliXFNbG8P0oLoOjL4s1
Lb7SJlfplYByxN+5bkY+F2zUDDlythYrr+/4MfH2OEEkHA7uEGjFFAMajpZJidWf
wYb4w7e6QGRntEyi9lphw3fLYTTSj85CPkUPjEfNlZowV7NFnIqvtmmKFqVo+Ctg
RpkWneUDMtS6SN/0nmKtCTUaHDr14IddB1o5/iNrWc5zPTTOMFe4eu5gO9m++aU2
ivdNT855GTHDnzloCeSHpCV4KFtlqJTKMPs11JOlGtbfcqMUziUQ39nsVT6Kfc1/
byoOysFv4cQmDQXe9PuEweQ3llgtqfISSk09BndGvk6Gi1C7qD6daVsEQP87AcKu
EWZnGVhET0bGftkINmIv6pRuOUkouLfyyI7bSiJDwQNV0JDukVlKxpnR72ma5UFl
5Z0Rbj4CMN6pQfYoqhNmRaiaPG0OAKYzvIeKdSg3oWFLm5E7hAzC8R5eGj/qqbK9
Jdd12DAkcqisPgQliBx8Trzr9ffZNAiQ7lOQyVESolsrXHUYDIvyP5jg3KlvxrN+
vKzmWlQjadQxGbFuK16zOzxzZaVf+6iyrJpWvPA20W2bbghrU9ZX3TlTpCNJuCjX
EIJ8ZmQT8bTC1r+vclIfQ6ijxtctjplz79K+ceGgrhBeYV8om3bBa7wPwU7KbG72
e9hoJluDpaMRAZ+H9cOl7teNMZd99/u9G16QtYxsJi1JUBym2emyGxd9iJnuVM6C
zPY13Bb13OpXpzpgMeeMEViXK1+d/j5jxQRc8djBwa1bfBF/dQZnq6riUzCSqHID
n907rQmg+dxI6x2cEQ/DLLtqUqEwGz8fZq5ZmfeGkG295o4ayQmVRCO3GLW6Fyhv
aqndob8ohZz9XutOBfS8ymN5onip7nrpy7+02jTjrKjnedP5a/nif+PrIno+LJvh
P7EaDbHmtdObSxItxUi3oqRAAKQ033ramHivhX7lR9P7i588VRqCwP9fqgnrPIMU
BCLrHkYUv501zwIYbZ0cTyLI/itZNugdG/giJtrs2B2R+M6ZnnDcZCbTegXOyFHt
YxhkuNYzn4NiFVpydui3LXM3FQvSXLszaOnKV+HKtDVPqrCImPKQXYWeRdGFOawi
Jty2/pjeOefajVj05a0xcsi04aYTU4YaOqSorOd8IyR99VCIvk/5r41Q8eoF/ebK
oJhKjqNTkVn2t8DsnMEa7N7Y6PyQDS2qHDCYKvWoa7GuzYFJCEXTgFMeHO927Ygt
/Q83owoJqqTpOr9zYjJ5WYP0WE8CXl2eKN96llHdUAToLYZGhpLcNgzB0H3uuzVV
0xhFDZiRKqY28LvsvoH8ZFMoY9weqqhLDiPjnhslHm7mFULp+zZDUgd/O/RLw53R
25gHHFTYrXR0P/751qpi0LRlEPVQM2zZ8XyB+86fxnjnUwPP6pSZpv4jiZaMJMZI
zac2FISviBXj/y7uOrZpzuL8MRHWOV732TXVFtiIxpsFfV3nhPex38nKdtaQtW0p
vzHLG0XgjGybyDjjY58Zv0TeHV0Nty9zjsm/GlWP0oB+byEcOZuS3nHg4Cl1jH7R
twOZgMVQ5oqYRrLaL37S8lbwWcL1ZK+7ou/Kbk0CcKLaOch4/jI3KkilpA2CsbVU
cKFDC832M9WXh4aY52DHLxn9O2pfe6RAepmXDlMHLo60kfDJjCAsTHVrTRm/wpaI
1JhSzBgPzL7fZ5QM1o21Jc9r58fnmqnP5HrdGbRjOsXiac+KZXPhtBAn5CqX1EFK
y4ry1IjFgnYZj7Rxoe4SDRgc9ZegOyozIRMQlzQiYm0CDO1Srn7iH/5qj9ELrXkH
t7n7si+bLETkhxcmLk98IHrVNSdHq0Wv+KwGrtn40EKMU2Ztp0WuX2JREyN6SYXB
GqvWrJvUOCAl1CXJasJPEYCz+75RvVeSgRG7+cKcuPwAZl9IgWewQanWB36OPGf2
+a8+obd798HnF5yLo0T6qC9uQQoD+GljfUubws67qvWdSNN9FMOivZbYpS3rWKGT
jYhHbUEenqRhNvgmCr1cYGPugZaZ0lWnZ3DJzLtaQFWsHJkpcQGtmrjDqAp91kgK
T35LbxNbN4wlFPBS5Qw6NbfFZ3dSFgVElKwhOsEuKmbd7MQw9x8KRAv2KPhIU4pe
XvayY2nn2zErI2Z9dJU8uBJo5o7B6Zo/nD8nA1t8VMtckE2lV6hiWoiauqWywMCK
ehq9TYP+3yxxAPzQQFFc8RKCLxdNqkSejH2QC4U8mcW/ELDkWHQrJLfvwHoXkjbN
Ai4UKSee5Xr8SnWMJdjkqQZLT5Eu41jDWWv+R9frxzDjbfhqSBFW+414ehoNqHR8
NEtmi9+IbjbCFrY/uMatx4LX2WYD9eelymatfPqJhXjTofw2PbGY0AumlkBzj4y5
hzGIND4uerzdHa+EdVUpNdO5Qa2Z5l/PAuYW7fa6ovqlzqigYxZ1PUSTJ1NdWktt
g4i1JhIPjFA0peaCEbq6/y0j9DY0qcvnAVcYVCUQ4vKOM6GJd8xEEbsCaB+zMS5U
+nKv0B6tG4O/ku0GY3BRPyJODNZlcexhr4D5ycdIL/eMoszBox17Y3S9rkFTOw1H
9tj3V2M/j/dZH3Jc+ISmj5cE7Ye6LqnjQ5Q4cEtCzl33ogj4lWuRmauQYGhWOZl4
5IloI3ZK921oq5Ezg93EW67Lv/KXUXGJG1xi6rkuRIDo5NGXxpO9hwySWvXhSe59
k4GRvF9b0UF9kx0gfx9ZaiBeOIva+0ljBT2xaaA17d181iH5BJJoCK73mfMHyQ5L
LpchKc1ce5EvCeSWmQN+ypiKX/RUAPEsKCI2bC3WKa2Ijf9n7z/ApnwN20xsWXdl
TXnqlSLbYSr/7UTOE+QYlea8+BpAHN5jFmoxPNZLxyHFUIHLUP5+6VgR1G9DME3f
WcTdA2emfw9fGmF/TuUZkbj+ye7kihHOy22AwLstf6PgRi6YI4Ns8QLwRskH5D5M
ckECjXmpznS5/9X/W41q3HcI+LB1QogC/6B7YlHdxqR+kCq6kksUxti9ivsf4MVX
Lu/dBACuVl8eq6bBMLAYd5lHeWCbw4XzxdeS7mczeiNGSUEDYSovFEYPE5YnhCDs
a4bzsIAJa1QWohgd4L4ZbZpdglfQMH/h6LzblztdAKY9rRDM6XtvQ+X0JWUmlCi9
lmpgsbAnvGvAzzHkGR3JFZNqOnlK0VT+6rPlzQ2jG+D3WmFFIyYja5AKKxftwRcR
wI2sKGFTDzGFdP9jqbVHpfBmSJpGNfd5q25SsgMTOd9AFf68zG6r/8I0UQEGHvbE
11jkw89Xi5y3yVyzMamlFba0Pra3xFWBJtXZQfV4AOpe3Y0O8o8at4y79/c5G6X7
RXYyujGzz22ExgsCVXrEbhQ0LurpDiOzVygc8xHy3lUtyX5ZHsICqbVf4rubnMDL
BdjykVQGLJsIl6rSr3aRvzeo+JtE8/urrQme5SMiwe4IVNl34JO4KnIIfJfvHovG
pRhFcC92sY2pSFUtvxbx/Rp/auMPpQoyxP4jicxt9lss+UAzd5oSzQJ3gBwgKsrR
uATTiX6G4WBjkmxIALrUdsI1SWeExfOhwzjKMHa3T8l+v2gpdNZDDZoLE8kBDeMF
WivFHhlG6xFKpIqg+33pMSla16smgegxS2N5tdilXa+hFdbDbPsrmNgJufzM5Bdu
7EzsdpoeRNKKOuiLT6Z6HWWJWpk9stkx85oLWqIOwTIFzPU5aGu0d78UuqVa5tIX
Oz4VrMH+z+dFXtALK6BwryQhFBXs6I/7lqxBt8EbnWEjaQUZJJuBx8qjTq2Clusm
aFfEfymR9h988iVScqmgAlTQh9JGzhYF7KJluOwn4TQfBJdzs+xuPIRwdqaTdXBa
Uj7yf+gH/t1V3ZKLOpBTMtb49zObeSz6kUQ4FOXxIS1av/24+/s9j0R/C5N2Z7JY
CTX7EVg5jxPWVReu74HJZpjAf7/BglU7mxo2yxqaeTmdcNwaoHZ0ou3sZKlA9qtb
PVuaj6f2drs5cMX4VE1jDPuZHPhjlmq1WMnu7/QI1POm1VsRO70hNi3TDxHJjlVK
1u+35lDrLUljCNN7RdgBavWLa8NoP76MnPz8vNfR97d2ELmFU37gojvXXDXUy3EB
9J8skXGnNY6iWEAPAQrPbXbNjzeh38slgtqIRWZXeqwZ0eiycXSclZr5QEWa00wR
eBmdz6EgnLij9vJK/E2q/19bWT83KDG78R6vmdgvsfXPruEG8jG3uCmSF6AVxk7p
hlZkC2PKy2JjLk1Hte5XyX1GOTaPpnjUEycdWHbqZE2G77FEgdPvmdhi3RBtFGym
V61osdoQNJBXBCGopq4r+zfj8DRJEBFF3LC7JOS3Rrn+tpp88is5yBYX9OtJCUK2
qmpEeYfQKNuS6NUF3zXNi+PuZM2Uz/dXCIf2rEkevNSDnVNqupj9nJ2EzUc4M5RV
Rm5HXmxmYVlNI4p87iJVIJjCalyEkvIZB9am4O17mUMgy6l8IziXk3YzDIFn0Gbj
rwV27NiDNo3r52x8UIrJ5xfjw5RzeFb+ci8h3CxBcNtXFNhv+ZO5NknxA+bXeWTH
nArcDWU4xCUa4oKn98LopheJzmB7sT8sZuglGLr2tXn9vomh4EHb7OrtWrBJZeue
u5gugnBLXblqLL28WxMLzLZH2UChSM79sjh+Kn6O4V/Z7U8KI9itPaJc8ex/m7Kn
2Llogyw0Fp4TO4j7HUHk5O2Vd45KpCDvxaHgUJaMFr7hsL+9OHmYpqgTqoC8IZFB
JiF10kw3WEQZ5cT9+npi6QCirxC0O/4caDTUdRTlPkQ58GlQ5mmSD7tk+KZpEc5e
zqlO3CkgPHq3zaxSdeEmkbI2osyvyfy9928WdQNHj3LiBimu44KJl2lpwrhyeAqv
OPpTqMGefNa0IZnTXZEN5pUvDAK3xF34rkctVf4JDbNg3w/ssG/Ephu5XB0cvKZn
AtNYMyB+6+r0HSYESJN0mNFxNHK/EAgRVXBRNxycwK/1YZbD3VC0QDgn5J5w+GY4
iYxOOEPpnPUafglmLSy7Z7ddqwUxP2E/cAD7BEAf1mD+4UZkmW7733BTHpPF3cUP
cVjZjpsx1khukLdnGiwl+SAKD4a/QjD5qqYholRxtbIYOPxPJNot6xr6yha4bapc
NLR+1pG4q89F9JprdI6gX5uBnwzvBeWoJ9xbi53MdX2q6erjnuQazMb3MRXeWDUQ
l6SloQV9KvrkqpapeIOLIzND+q8JCm2nRdeGJzhmxcEaNk0B4Jz3GYka90d90QNG
zkLh08CiORR1JFk1QXLKcYAujFK01oybGpkeXryQkzewzNScvNA97o7pJ7aJA9oc
sAR9uzv8j8bMkzmf+JI3I6nIEYoc3+vOqNWgRXgBf/tW7R2KQJdcLsrFOvn7aPJd
sRquSo9BdwhsQXbyWmQK+UgANzKCGOmyQ3wQh8Iz03GedMPc8IoXjrvjL2wjEJrm
YWmcOHhMemvqfWeF1ur/0i7esFkJwGT847Zso3OiCq5l6Ok2BCyTu6PFae9Ba1BU
Ztjsx+/vUE/hxvSC+jIRhIQ3f1DgXMaisTSs9wL5KJoohZ42rgITlfSkRykjPNMh
ltKe67JB4nDD0y8mosKmNlvl95Xe3aZ32wI0LkkDtNXA1geOdaBSFtxvD20Almfo
0uL7lIWsmIiGYHaRyzDA/uID6jER7GO76IT6phue91pzL/F9uyiCUshazpjAjDoj
15RHwrgmp7QTh+1SsGp0kETKz1WBHhPEMpBLQiVeKptaRGZKbt9DCD5MXXaSJJRv
dToM4uir/L04mqQ6eOzV9CfULHa943NNx0pbw+Rh+Qa4V8qLzo/g+1ubCHmRicDO
+L9JJpBBsA1yPXCUuVkRdzE9w6blMC2bwbzLUP5laC1O0+qFeTxtBqIptZ0quO86
NVREs9m67VF8eFOOrfDFt/qMmAGjUWvlC+MOPP76LcPIuW+l3o1VDUlr8n59XAsX
B0RBRh8KLyuph4RNqyd6JMO1DUWM5ObIGCqfSNgCQgRlbUESSmHnLEMwSA9oL2Pq
nEjklbrn0+Gs2GgVInSMiPSDVNciX95t8QYAp3tAYxRmYlBYPKfZ4B5o3Ob0AJ8h
HZ1ZJtkjTvWyLpXcrmDM8I5f+TE03dS/1csT26SDRRlKeM2TicGzemccoxcmFzrT
u4dqdQ9U0KS98Ug4s9D3ngUxDahyP4B7ysVTkD6+eNKlJP0mehrEertdOGMh3/pp
ngDxH77zHDdXzeNb1ryfmN9S4q3cspYmjdoSrS8A3QULme1D9DpUlAuk5uInsp8d
qjntcc1dITQUbKoMpyqDYYRPHwl1JUz6GMWUz0b9Yku0O7Q0pzMszhokIJKwBOT+
EeIvKqvuZWwnSkggunW+hZ3uVciMJJFQRiCPX6iWtX1wmQ00mZVm3CDIshwMu4+j
gzYrY4ZuCHUxKuzVeQyBE57QLegtq/q+tqGv81a18WCn4PhEkSNHpCSddKN79DPd
4Wz9Frb+2qsycdNrkzGDEUzM7IIKqT8x8CSFog8IU8e+41zR7pW5RYA1U5RrvmT0
XzGlAUOjRqy1qoeW32eZZ7uTGDIKcnWes7lLrzj9bpQZuA8VI9Ea002XYvcj463n
hX8Eiw8YBPwmiAnRr/fspQLNtd7J5hN2KPB8gxI7b4Sg5TsYWYNgFYPB/uLBVfNf
WXNBiFC7toV40yOo9pa57zwt4cBkZe0iJwMDmmfuuikShx09lJ2efA4SbVfv+Dp9
sz59AV/I2K31OMKBK+UVbm7ezGOxQ3+siH63uXP0RHT+6TPMHdcIzzKxfkC3m26e
motrps2DUU59UoKAyVWsFn7iHXjo8GfZq7Vvi1iKXH8I7zIbpFgB9+zulCW1VB3D
qBuh0QD0XLNQKn5JEznPeCZcTylwZF7qAHKoqXwYIzW/SFTYr3AdOdFKhxRmTVrn
JsIe/Bo+tofjb5ZSr+jh57awwCjgePt2iU5pOJmr4qhXWEPHjWwjRtcrcmv/2HQA
tKbKBRath3/K/r9NzGkh2NMBHBf8XYuTdQDqLA/Qe50Y1uQnnNaPLmSgSPjgugM5
m2BsrMc+GXMuNZHJLg/p7d9NnP1f+wNtTb/LOuk0u2ZyuCKk1P9P+wkK5WB35lBI
vci6HpBWP1r+eK5YM5Jt0Mrld43664KNm3jqSFlE3WNWNcI47JbjGKitAJZrdJh/
JEV8tKHOUmjE2+e7XtXWHGV++cf9VmsTATV2pEvaQkJXMZhb/x50x8OHtm2kllMA
MiGAdvYnYiOHSRLyx61e7we8xpltQOi94NK0SYBJbQPS1kd5Gx5n2RlfErhlBEt0
d7v97c+ByY5F3YbF2oLI/kMxUQeGJMX8KYZkw6PxVXtNd7OrnPTS1CG7HCCJoTc3
AKB5asmbphM2lqqFcrKuOU62UeiECeeb9Xj5GPYMQEI+Yfut3k55hbKdjo/ISB+2
HNBGAwWtZrswGKKIas6mVeu62VB+kaPs0d9/Z1zCEQ3AZVZpaUfoTb+snwpZu6ao
/coT7AFzutc/6GXHmuAepK46pWdmi+XFyyI9F/7HABnzgJIG0cLdSRnqu8RiH+Xm
OrSc92qWUI/KAtFo+82mN8quIZX/6BiX0TslIqyfyeIqt8DTyKQTXXpYKv/EgEsa
MtcUSOpHdlgW6XL3nK0PTPA9yl462cmis6yFP8vWtwLuMkpquSmJ89w/51jEFLiV
QC8W/XI5vS3TIp3UlU4RCmYaz+lxdUTuMJmZQw+w3VRqo7y0NJJvqjDyTw9ihb5w
w43Edpo+pRZn5BXKokOXz8fW5wlf9A08R3JL1PUF/sYsOZmV15lIa02vpl0zrN2t
yxGYlr9kXsvBE6ZtYxZ+1GjKJ0zfixz8Cqb0S7JdXBR415VSAXwQboPeGbemRpi/
/VLJvO02deDVxzgwwMw/8CH3Unb+h88bwp89ujGwM4jvIKrgLsiyzS1aQ2Inqims
9OOMDGQGYI0hltoJelARyJdG4L2OFeea3yhsyurdvLuxaCzRFQt7Kyo9aJPNd3zl
md7qndxtDuQMWSt6brmKUpmIWlXL+YnhuyNaE4FhP7wpNBDsTtC53umPBLvaQFG6
0dGgAAZcbicCKT+vXE8rag2MKRYxj0WffTcqSiis7WPTlaSNCabdyqumSRdK2oz8
XijbVVuylmEjgRKw9LW7Ao3xUv0L9J/iuDKwmfTf/hfycpXe57Wfp5gCC2Ax1KVo
/b4nrh71lcu13K8TvOaHneROEuYFEEVJ0U0i1csu/z52ZIvfs2pDaLku9QRpJ2+e
cCix0rlgRwpD3Ltu3bfx+4KhrXUKrdiuL2E1BJbAqKbz/FXMitaGZilwtnYsdUq5
VSscGnRLs5lJ85LQB2bJ+BhqK337gRxdsJ58i6cNO2DbcuEC3227wDp2AC0/9U/P
mNvn8mE7cA/9wf/6V571Dxbe7hFIxmqETljOwJykhxVkV3HKTJs8N2JZbX4ZT43C
/tB+uMV0HEin7E/j4wFV9ds6z4m9sVzecHeaCqMM8snzFBcOIRzFpPqTaVMSkD3p
yXf/4dJQkx3mz2+J0XfApw9CjT9XizIdfinIe17BaFFrNGHVAJa6Bg2o0Gi8c0/k
VaD/bYS5fe6trpPRwzKknYqBCqS6beyFWR1JoplLmmMjeQ1561bM4IhekMeZrl0j
mwXw/9SLTmDl7+Kx2o682HEt39XqAAkENXPUlM7YU0SSgsToRa14zT/UbvtVhyKA
7yQL9yb4aTBuJxPl+0iiuXvi2sr0whQ6OWI+3dDNkpmwQJyW2VRs8b0nda1KO7q4
iXrJvICgcU18ub6Q8pVgmSCuiUnwTaESCe7eM6q+pwDFvVPUopRlFnKjNjleVtCC
YijlAS05T3vTORuGy0qYcD/OjkqgUdnJcX96Wvgy3sTzgO/F//TY6UtBd70fxjeL
h/4oNbps9c5quz/5sFeeXzG4DUjNVZf44SjPkRL0U8+b6iEqw0fLWtTQvhXSDzBB
aOiJwJD1QhAUkS/q1hIH1gYM9BIkh12LwgGIYYvwMwvQlaWE/YVK9C/baRNGsC6G
vIwF/9FvlkmtUV+xvLlcJGW/Pksln+twQpKJ27Gv8Ui0eeb775PjrOZaGcSDwt6E
RIj6mjXSnqqgCIkhp+LGlstpgW3z8SEKolFiGEKQdTbg6Txr54krHIVduUDdl9ZF
hwQh4A1xI/5Gkl8CqD8XgyoBk/pbckrRZ6RGGJK+5OTZADVASdm/QU1vNWRdEvcc
hvy3Pa/TkkHKOhTdHD2YQi5oFiOf2B3mB1N5VLWJFCzocH5DrXSoTmV4T8QxMJ5m
qlvx9qo6vVnHgGmGYMfVwS9dJx8mEGu7TmlrhlFxCuFe/WCu2+aw9rqy8myYnx3t
tzyH08o6HcRLBkTC5XBMZhIq70tsNKiFeTAqb/WM4ksZehtwnHqV/TMhZtICEJUg
EflYU6vE7ZbHNEshhiVLL3NgryuOg/suIg/8a5xSA1Xqeo/HvrIdDXRlVsNkUAad
ftbzzHyfgOAHDIduWWqKZw8SW/OSvBHGMhGr6ptqr2VqxLYL11AMSTGzC3B+R56Z
oAzIvARKL53Wi/+O57HqjmkPUowO27/87v4eeTSsnZq/wEyaggJCV9quQTsjLbgV
ihwMuUBvzDhqWz+brZz5GB4IEY0s1S3Is6fOzOnicQeVvsFifCSzPRJrpuATq3gr
pYhpW0SAEe/qPmVobFT8AyCStvvF3Xw+mXVwmVvuK1uiJkuLR9Y93Q+33GtSTnC+
XFLV4gHIcuA+ne6tnxC5c01cSx4M/QZahW/HcQchytD6R6ZrVbqCeGxPkFaHV1M4
+r8L0rLFmfJbHhGZ4FEAzHAKZVpr3fROe73uTs58O+iPtzNS/bshkXcisvjdAIIg
eF+BWsdDGAjTDssolu7k3RQ4BPxRS6zTu/lJDcQTFdPNfCbRqaHN073ipvx6ajLe
oCuwmPqD69jmwdqEtQmH1YZrfSGc/FFMchZnRxieM7pZBdk8wynFloFbwfZW6DOH
54wQ1LK0LUgNOES5gxrxbgBePo/fQ6TlBuzu2Pnw+7eogyeQJYyeHVQ+0FJzWR/b
ijwrt4kNJsTw5m/YHNtC4f1HeNQtDNeoitGdtbaVzr3/ucsV5wR6iRHLrJ50Qz7b
Zpb/0vcwiEmE/XfcIm/de9YZ42ZLD9IuB+y1UYEEO47wR/o80aSYS51IK2VCgRmW
3/S0fUDYC7PedbVWpFVJDbIlsKzoekFJugMKzXJSBw3Shs504zLflpto2GWKQlJs
3WcdsCwX5hWxLIWRR2gZz/g9H32oHBlX+ln6nYe2EzEA1+5ZdzQfwR00OVT2HEDA
Y34icoeh8deJjnAAoRCMeozwIHQr3eXyegVexPKUHqTVyP4rO6yJLnZNbXOm2Cl6
FuAVCglHiGdYiS73Y15eZQysUMQQOMpD4gmsEV4xNA96uD79DAsmbAR6y0ZzqzPq
RU2WGbXavZjPBg3FHrWhyPsE+LcitpfXX9r1NMUehWF/zTCodCu36p4pnW/XYje2
FYSh/6+JawBCp1QuNY0q4qbrORXZ7xLMslDdVUfpCYwNPRuXNow6tpI0vNexLUYF
GG/Wiz/XWIIsxYZ34NmI7gZ2z9TKR9f2CED8pGNkBZeiysmmG4eAPg5EYuthXyIC
XTPReP0qP3FI4GMRNhPYmmrcli5StPECVw/vMDrQbTPIickie4wQ2NEGMFcP5w5U
GauCzyrnJM6yYy2eVbk/esZR64N3eqjirAvfcTXyBcOAclYILMNWppm7F6wux3E1
p0UK5n5kwuMw9Mbl/rqGk7AumCC4KOEYoVEIWCMRpznL1v/EBBtA4swDn51FV38C
qLfe+eRqwuas8stkHcDmVjspbz5TA0sbPKSPcdyvBO+6APuVPCVPle+A64NbvRrD
vCetMh8BJBxFKciN5nKv9AB+vrwivrf2GxFNIJ+64DxlFBEgtMnisWsJRcZTG4Ot
VGuYY+81y7SY21VyXHVSm3WjUTZf4eIIB3CPxDiab3JtqInIF4/zIMlZJCiBgqbc
ykFDHNlzMjSZ+fJ/sCVmyV8nGOYOeAR6L9M/vCKqkHFz7E/rUgh0k7i+Z/fyJoba
8IPCVVaInwHCG9IJO9n+E+NjtXEhfZi0D758XgAgu0wSI4MReWS4uJ7F1lwxM6kj
0joNYeWzbFCtwntJjlXzVTbLfsLIT/NCLjtxmE2kNvNllcbBkRETijromyaD88Pm
tniF7+fHu4OFJPofEvLcOsovBlEy3ht2la5otWenzPlVkmzCMx+XA0bTOiQ8JMPL
ebcensAWrLq2lF/kxbdHhOCWyEf8P8DP57hCSv7aKKV02EqrW0IBI3ftv8n2WOBa
tE/9VKpLm3YcFv68rIMMTDDfbwkoIXpob/97mLtJ/FMbgTJTKdAP6u1UMTcillyi
p95TXCeGkzY/0kEASPEAFdqAl+rfm14SS7GIfpP6VPtlLBW7smutTJZkjygPSgtB
u1pHPwDnegJPgssYHRTzQXmgjXN8gJwNusBHZBZX8Dsw3GIbRtCDOOXpv2Ou1oDw
ONxEJszSW5b2LBoHH+ievbVlHCdKV7sI5ExRSdqvwGnm+gPGG3tbAw4CkQaoVOKH
zlK4kZamUDAIrMC5OvonBrwBzExr5psvbJYGsTHkC6GO1whx1S8Y1LG/GWZ4YGGf
dbh/HN/6obL6FP2Dsiw8Rke1KhPiBizCi8f85vUQ+7WiLWFxdMnIPDPA+oAlTnfI
/8sRYHVCK605Wy8uTVv1KlQz/5Tl3qLNSNK3bLX7k8SWtcby/bkH5s50cdB6P6cs
vLJkUkllNGZO2gB68dqdaOlpDjTGsTM8vc/YC0vdpUzk+tniEf9J4QaxbQNhDXx0
G7fJAXZM2l1tTkxVjebZCbVGPh7/emzQn7Hik5ZFy5nYFz1vYWe/Nsw9eZXhAxaR
rd37wS35NonAg0vtqmXpjNsUp5/tldfK6c81j7Dxy2uE1fod/RvnsifqICljsiut
8KgNq4Malaz/2HxcK8WE9EplQUlR+MQjzA0iOnckbkUVQI0KNt7duhKWryOYW5TD
viKoKo99uWlb2OWVGYvN8TcyL9N52O4jf0fc345Y+HiYaRcz+nTbcTU5zdjhVJV/
I3rTmKsHtHpoHZ5H2jr+YF3YGdJo80RhbtpL/FVlgWtn+S+FmCtRTRIYy4a+Sgk+
a2mdOMXkZT4oh5gTTrC0pP/nl5tVeIHGgHqUHwo4QJi8ULUGMfTjHDuNVf/rFBmu
+PHn1VA0CZaf35fF0YuPNrmUL2L2DBNybWhbSZTkfUGuq2FSz4lqjCMlrj7lnG/t
uKMr96rfRwUqUgkGkmfZKZbtLMNkD5NaPA2EtO1mAnaSH0qyUV9auAALOjdwa8+q
n4LxtbONrx6E+xndWS0AUTqEXzrcMDzPIZKb4GS4WtqtciXMZWXZeeHJCIb2BPXk
9TjdVsHJkZyeTot1T3ZZqjIi9omsEHKrgLe7tiRxHH6ybbxu9/z6o8EIB82HvYcY
`protect END_PROTECTED
