`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDi646rIEy7wn5uBy47hw+Yfs38RDlN9hEDvDICxYmgk
bwn4iDUd3W83EI72bKA66dOL5lSP9wCLtrhweNgjQM7lhixgq0NHpmKD51/mPPrX
dfYxcsVDDypnBvwCdErW/DxwIVxfvaoB8vLNR0HqKQJYr6sQlfja2ayJ6cIWbKbQ
Kt3c6drIhkoV1u+arAZCw/SxtQngkEZlEeLXJoAFE2cARaK8yEfxHIYPt8qNaM5/
`protect END_PROTECTED
