`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJeBPvCMIFUTZW+ZKyWrjc2FVCP7KrWsa5xHVITHYqyT
TNWmogc18+DS0DWhYzFGzdF9QiapsptLFE6wiQ/nOKHP1dOvXQ2X3M+7mgVXT87G
olop90bQhmWsgRaERX7QFXEK+UCNtWgG8Bdgu6woHhrCUE+VCwpcq8j9rkZ1x1Co
yJ1s/BA1G1d7x5k5RKe128TQjs6naRUo8/+C9E9EXbnQSg3BFxyPVDqipcLUiLBy
p8dX4UEu0XhRjGjm75miFmcXLPAZjwMMTZeZbPCaXyOybESP4raqb8J58G9fotcG
cHn5BikDFmYac9ytDmNmlpbV1HhOawCgWaSxeKwAizTXtl/JecG3F2V85c+4Xwyu
cheMeAsxdOj6HRARQNPHbQ==
`protect END_PROTECTED
