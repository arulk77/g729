`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40hGiaO3tONs5yBWKsCS6mbczELVD9jS7TMZGFMUnCCr
MQ4VsiHyv1KrL8wyEAhGtzLD+ypVPbLEkJTKLQ/E1lb5JPnHcEecsNXwvDPHgBiJ
zwG/nG9qHLKmCXZ7hMvtgiOV+OEvj5QZYwS5vIEQYcFKU1iIawah3JGOol01C4UJ
qt1oaVHlYIGzbE8BnIDxnJka9rGMN+ab8GJp6+FaK2bUNCUsmle18EuIm4E3HvZ0
8No3OLZ9Ct0TdYjT9G9ahyiLjpFwlcjZnGLwVtArYMnLzilmZ7i/IV4KHxotD4N0
3DLpn1CHRwB+/4qSuzNT1w==
`protect END_PROTECTED
