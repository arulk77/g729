`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAYK0pb6nI+a9zR4flq0Kl8NkEpGo2jaQrvVvU4f7vMK
bgbuG9OKWNr/c7iP8G3WQ7meVfIvs9AMG0M3UwGgWvaUecj8+NWNYqvAr0wEYHLX
J5nZ0flBzwt1sPvvPF8jf7cqQz0Q51XhPIYwckkaley317yVMgUhoTiay82XJ3hG
dxwri4dsgq0owmC64utQu5uBt/PeOPlq2Vpco8/Mu92flNDJ/UGnMW+JWb2qTiFi
SYdeivEF0RapLJ7kaPqGuUAplbm4gXaPHFyvPhRLZEMoAnOuGVZi9BsqrhFVv6LF
+2V6OoiAbBnTeP2gFbYBwIYcgTyYheMdK+bZOO+GD3qaeZP4DjBH76RcyHiD3jbo
S7PryJ9P9BPHylGg/XC9ag==
`protect END_PROTECTED
