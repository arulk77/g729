`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAoJVOuKH80pjwdFB86YK1Usdnu9VXT+cv1dmAHk47rz
Yh63iRI236X+S0UHVc2d3h+8V3PQc+wES9C9U7PF92oJsianCpVc0ewZLrO/cqui
WlCtuMCHcDS2hAJb2IWabbRQNZvrF5Hy6k5ACdwuBpI+P7p5sBtXNURV2w/vK+UB
0c/I7+CVe3pYqmZ8B18djaDrvp5u0xYdk65klSTokR2T5P5JSf7zKYpYomlrLJzd
Vtjo33nTk2SV1Eq/y57oHIyt3LhQreSqJ108EOTLJZo1mqSNh4PQ7AEvL9lpizWz
NzfHc7e3LdHjWyh32poVHhha8QSvEPVoOYmvR0vB51AGGNMIoM091if41Or0D49T
5FQ91iO1kushvejZrLUJyuNM/H7XhyrUK5gE8+hTZ7SBv2/Uk4psa3K/KElSY5Uj
JB3ST3gzbPtSRv76RksaG7+x1/GExDW8ViFOQBNIkaFkmPASDtCBXh2udkkEDJ4/
zGsjO7kSR5GDkoJpXKtAXTtIspOoOgN9c6LBCTrSbwBwBRHCRT1376m09HPqSzTX
`protect END_PROTECTED
