`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
kiQVmPJty2Y/g5VjyKurwtvPClqmmOkxHa5alkITW7ufU4j/SXv0khT1Ms2rOp5E
2bFdM850b6u/poAm7mByrH7JDeFFO20ZQA4Tjhs/iJLcJ/ERgxqR6cbAcL+SLKpe
prklLdqhP86tWyoRyoSz5F2J4fnoYXkiWv4tItLnO5wtr6Gb6H5XzRdCTk9ZVbl5
`protect END_PROTECTED
