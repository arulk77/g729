`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePoSg/2xaL2Y5v2F7jCfHzIcQTNIf5wTSb7K7wGjXeKl
dvve9+kWX7gOAUAQrUtjfHAAXbTsjiVwN9S9gxGx544UOponKv7afNo9lmR4LQv2
YBofz5uH4Z5LUZeZVNgHyPbsoFQWncMdHk3fqAv3+FhkJpqNQY8rXinTJ0J5sfIx
eKh7c31QEyYZ3eZKELhmLLR1YKiba7+Czs3zbZKnH7a+qTjDzcAKqJTIAYxClvGa
wGHCsauCjRVkJlWbJN0c9yhY6oTPS2dvzl1o/WNlgeQf15qt/2YL/LadShZGauLi
VVzO3JZbMfoUQIbirWemJPdVX2+rDoEgbeFCgG4F0+WwgLFZX3kACIsqbrXLQETB
ckI840x+SkMzn1x9d88DhmV3a4QvGVGV6gAwe+mBU26VMcsEElpLemJW3xYcI6LL
MCNf0bpFMylRAzPcPT/glp7jXta5sFAlp4XFJDsFzoeq4DTN5hFangHc2hru26zc
ojoCndDsIIV3ab0aeJQZ8HwLiaLySic0UgFWYeZXtnuMDN4dFF4WQfMi3W+V5Q+J
oFQNvzK0ZZtiDshf0k7CkuvBs/7wUWuye3V4NzHeGq4aU2Dgqip0SugQRQFylzqp
VD0IlwuwLUSo8hFdIvXKNFiwMpj2P5FPeHuuoorSMEjlmL5X2i/R3vWzkhott9fE
`protect END_PROTECTED
