`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveO3KCbcQRnFJS+jFbMLxDaMuEIHEf2QAiDnb3QLLfc4X
RWlfFJ5aZV+n14+wRoDxR+YsS1g6Feso2lnyoDd58dUnO4OH+EWlUVTMbalKvVJ4
lrFE63TCq8jWgI64LguTS0ht4GGAVDgRAh+sO1YYePe1GnIFwcesT7Ow13AeIKr1
GU9VYNOFj972zW8hOavPpn8TxTZK72bph1BnBvx6mnPMOC5jjntUqW2S0cNca5NZ
q8MKZuRTbfzWTW+5IKQyHE43ye0kxdtoX25daErjQMzjCRr8k7q2CgJ4R21J6ej2
jM1BuHNB6tefHey3dIgctiS537iWfyQU4vJDGlVodLEIV4SAfLtjS6Q/A9DAAtq3
DNo3mn7kvF+OiyH0Y1TkNYo8K9IKnvbUjy42xaCaDnv+qzPF4W+0oyqp2FiRTbVk
W9O/xidgECBnyB16EEZ1zW7P2m1QPQ+fBnx9923NAzuedtfh2hcVXyM9SWTytYj5
`protect END_PROTECTED
