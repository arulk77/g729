`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QDOGuLErBihCgglDGS6i61gZ9gt1qcuIglMejMYOrgnX1nUjGRrXMHVuGMyB6wb8
WIdXzl94OrVRX4XKK3YqSNIMWGVay8/peFeKBB52s2CLAhb8+kQnG/Bf1dgkRRD3
t4npIudSjuvEnA5e1msP2D83BbPR92B8AvSekVYiD6ZyVHoC2ALGg/jQNwz+0R6v
wcQUv+dEio+PIW2vv58mVRnAtjnzsw8tD1vV3A3hmJZuJ5TlRk6laB1sv56rcCIH
6tfYHtrho2wcNQz/57CNJmqK0z5eGzEPr7HkDnObTZGsVuVqGISkvSIaaQG2Jpqw
ITNmktg1saGuGp185kMGnsC786qR3qVz+i7GcfYC+0iuSJvPFkh76ivYVIg89z5m
hoQhXMoHM4YhmHw7m/xFymgCx3ZLWCRitnSYpJf0JUlGeNny+uKsteseJJ5+dvy2
W7dxXQXVtP2LXbFt/XTBqlnBUWIbeCpEec85Lkv1teI0mEB62pJkvbQM89YKDVOF
Bzxa8zlgNuX2ZHm2t9kasY/GU/2kvPQ1NLcGShKcv8SEgxuVQujYVLl2tCGZiEZK
KrvaO6+E2ziGXJZv/kH7YIUqI0nJWB3bH30efADiGoiYqb45ABpvBGyKGhFIYOWE
JR8mMDWQIFZv2XGJ+vmH2TlpEyEyR6mXO57BjOsgCF5e87KjqhQOEf5p0Ow+8D92
m3YTS83W7C15KgbZnUOMMQQ7ebgNwCFTRIejjVzrhtooJed9bVvwzzHu7lR7CDs1
n6dIX+jdUWOeX/QXYBc8D0y8+mL3mRWsA9NBwLEP3RCgAqKIkZxG8qvlIXoioRAR
g+6KQPQHUCg7Q6priRhEWFaOvDzHwZJpTAzV9zgaXIL+wmP49jgWo4JcicNWehHM
TAcmgpb07yMNcNTzY/4s9khKgryxHonI1vkkIbmIH7BEcMB8MDvXyr3/brVG5FyE
eewjXG13wDp5vC2Q7HumvDo7lRG5aqM6ps4Ru5IQahkFP0s14pUu29VFcX+QKf5m
LItBHl6ep5yCE1DnE5v9gXaL1o60B3i6CDFzgd7I8edwS2xi9l+KiC+HmW5qCXXz
YkGPpYhXQjKMGhKIKVw1MUgxGUDwaEXhhWapMzwTocdMSljvp2p0F4T/q+7Js5Y+
JTwF9s0nb9NRf+GiF2lU78j7WiTH2yrQ6SR99tDywHIlbOWnhqMpUnOTeFg45YxH
ffLgeU56dRmX5qE19fkpXSxVGNrJq1YLYqwxsCewyOnli8qC6j9goq2p+763iZ82
/RTLXCvF6i3QjQ6PVTizKKE0pCrc/XuGZWlTu6j/Y/xnzjn9qNGfOO+hoMCvAuw8
OjzwugPy9aJdj71KKz/jq3D2AnJ2gzNlHyaOAk9DkIFJTV8lOEA1DIdPkYst+g3C
1XB1iDrgBvxL3XtQ4yZYthn3t7NSv/K0qT/fH62+lTz1iX/hBcNPKSvkwVDcr3wO
+bedIcRjTbmgfISnSC+m0peKjo2ZqwtI1joD/21DINyj87a7Fwhe7Xyhc1L4ozo/
r9C+k+9s8eHs+VVI8tnsJsYRsMwaWEoubmTuv1tmqnHULjHa7ZVNKEGPRCANcApL
huEVICfjZorNStRJfc1BkTT1PPlu1AZMq5J1CSpt44JAwlAZhOBFFn683j1Tj8JZ
24pGYXVgWXMVnuhM1phlAqBWsO/LIfbPKnGFNzNPD8XPQKMkViY1/m3Eoguuux7h
/0AtMbClxDBQLPCW3HFk7TspFnq8N7N3TuhCo7Xy42haQwJbD01dj3PI23k1f5ER
YMRyjHAHhpnYNCa+0NoU/gs2mGyUJKJGLcLiG1+ser4YKEMJWc1UWBB+/rdl9cry
votJE09/QSqqH21ZxgTW5HcukcjmfFcKF7M+FuXefjrhfn0gBmZUyx/2CpA5nsMt
N6lXL3+4tAqhh6sZOfYeatJWFmq8HonwC0rbENi5G7kezPhBmxzalcl6KO9uF3qo
Y28/MfUkkErJ3o8+L1Y5QZ1BQT5zQbttr2K0zX83pHZXHYkwTznslEODuJAXpw1N
UTHtvq4l4zHE+3ogWacMn29tynZFSMOjoL6+S1eIBITa9GQxJm7i06X9afToUnRh
jT4EQHpNAUNaZXsjxcq0FoP5SFBRhLBOczsrfrseF5Iy1uqtvHExgGYCz/Rg56vw
CKSAalcIUJCVUcmzn5ofYawz+5bJ2wcjdNL0dfwbnAw/WjTeA52RJ922Pbt7k2eF
zoNom1Z1pn96Sja307cTGVRiZ4SpJo3RQpq4ig0JeRnBgf/Ul8BhJP5EXF1gmJu9
tjRFqAr7QO4s78n8Y1FK+dCDNOhOkFSeyBbWTUTTz59UHdlktahlnT5jqe1qs2te
gYSp4wbW8ytyvPbfqaw9miBHi+iYI3BfgVRWVW3KZO362rbaBOFbzNh+yRhAoNhi
Szx5XAAPgYetZXv1sSftmNdZ5J+2T9U8Br+rCJd3iGimT5z+XDLQh3DXadvwoqmw
1mO8CNo6OzSyWU8quFJONO3mXFNOhp1nPb+wz3kb/zddCLf0bwl/qZZa/mvNX+EW
mVONWyNHw/tt9/u6+vrGtll3eGj504W8kcSW3zis0Y70gwRRGCB/Twy4nY2r7KwI
OP9NmcS4muEJkCvuEcBFj597zZb4PBGBMlI+MNPpx/Ipf9YVtQJQyFAwfanAhulD
HX/TCMLUMIm/metsG/CLCfHgW7Zdeu0KhvNi5Cni0r3XFjUdWis7JGe7qSrDXu7H
LFkIFwals7GgpmxZIcEToFHn4QqCWSaOrf1r6bemVDlWDnV+xdr5iCaZClNV35Qo
8TZ9mb0oRxG2kGixDbcGrY8syH3WPfutDwTecF6+0Dw3fJMaXVleeTJmDTeDFeeq
X+IUT8z5N767UIMZy2Z0kOTcrnF0wSy+aWUuyxLUdXhPnLZk4G5w/LnUJ999W7LD
ERDufgHvCIt8bZVFMIljaRGFT0M1pdIbEHIpzeE7Ga5tbWjMEuWqtfccn/PLCxMb
sjLFRUx0yxnNtoFJLIAVg+p4pWs014GTg8gbT3NsdQHU9mVa2BmpgmNgfQto1e0c
1TQdOxCu4ZlGtopLhsCAVz8CFaV2rzdr4NEKVI5j4wOMZOusPejgj/bEdVuebkMp
QnU8fpAyKNJ4qIguxhBeeM4Gaa2yEcUab5mXu8Sb1MdcTmexAI/42+4667gGUkR6
hQmnuePZNTkXHIAPtLV3HEctVDC9Cn5uqzInmViOOl4gzMmXC0mWJnn4GjIAVwiL
yIdAG+me80LD9GZYzsnNSZkucQ8IwqtsmfRZmwHoga08yvvkpUbGkv/BlPOoWfar
sgazbMUupS4OwhUVLYUMW7noJ/bCj4dplZWLCAca1EkgtRMMlBaNX7utLneAXwzB
ab+AcDso/wA5Abbo638b72790Su5vwMQucL4Z4nFm9Wr0ObqI1xE8cIOVSBx5mYW
ZEjuuot5+22rSej+4/uqLjqBCp9+uTJvJj0+3tzLKat7Dcpbf/Z5Y83QUcBAVrxy
GCbyiTa9cDCaI30QeqiqJ1GANVbenbxIyoX8SKeEeouL499nVIQiZ3JPpab5+YGO
TbRi341uUWi/1GD3fuWZMw==
`protect END_PROTECTED
