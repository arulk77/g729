`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIrtf9R1HYAarNWpDJI0D8d6/vOAYORsAhVtq3LTDhv1
HbFhvn8A83ds8JnHX2Rm6UbRGT45vl15Eeuc3FP4TlEJUZ4LMykSMFS/GbcucJV+
swHBMCG2OrynOXTUkQRkCqGeP4kZHG3RXog1rrb0caG7Vb+Wy4OLwDNJYulzPxCW
Nne0+6wHVMWH1/XNwTk/jTQjw/gprVYSuHOVvI4HYjXjq0Zj4FSLjMqpmtwy2D1d
nFsJVXvboDCN1jpN2h7bGlCZAj87/PNliIfqtutPotZzidGIj15a11DohrJcA/P+
D9M2GGySiAnhGIWaJfS4be4P5D5liZxASkeGLr/EHbYI3bJ3U1Vb3gO4qnAv5Xf6
WEfJfM31EDVdTyRd8hW0MFghLZA3koDXRPe89LgG0OWKLFywYX+MzpoUJZq7QErP
bz/uYcwnnLvRXcR33PqGdW/9WJPAA9Tuw9D1JVQ39XSt0XFBbJJxD891ApjLreKh
ABTfSDfoSjYasdnGjl7r/0/Fcq/UrSJ9qCqTl9Ls1Gl6CIw8ALOG6clXIiBwkfRX
sWBTsTrqSX/ruNwIFqsptFEkVqU/BCkiGoAJE3QdSKFbifcU0N77VHHE0f+54iu0
u9h0DbNVLRAx+GTCmfanHx/j8uQtCgNvQlc+llPWKITaOIBpMrAQCw3GSkM8FP+f
V06z4xBoPQtKqLNQOl6AZ7+ab7uWyNk2ldDZsPrcXFeN416RvArV5/Czwtc6Ydez
J/zjaG8QzGevhMX5tytekOuBiXWszuuzMSw+DZHQ3ANQlqo6NOufCgwQ44U8PgVY
`protect END_PROTECTED
