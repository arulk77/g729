`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8ScFN5ufyrAGTrr848IGSJXZt3brmyzmvy9DNZ6HFs7hq
HsHqAdh7ncgPWMpJenwYNdjDPN/bTGAxbuoNtl2JPrvuYRA3qED6+MpHKeW+oK+P
m8OthvxQlWwq9Ruj7AuCFSaMbKOu8uF7AycHDatdgT9cXO2I71kWQV6IXc0pwfvn
jA3IxJV9b5YfLv5m7PnU9nlmel5xg8WmfU+GhMEgWC0jwV6PV+iMKs7ETQX/Y30d
LsEJbnVW475hF9ZTO18FnpQQ9ccrD+U5nFgWWaJGjEKZpe4C3Ajioy2YFaAvL6LD
9PzYZ1z6stLuZCkapSh4XM69Tiwcov+n7Fa5HaOtl1fForLjf9l9SGyafUbYdBdu
OFm7rV5dSUgj+aMTrmY5wmaFrbp5uDGpfnsYmAqAlUdpV2e5AsR5kp9SyjygsS/f
0aAYX4fQzW9UnmzhjxEBZFrozfI9L63txEdyW5SJSc03mKLPm9dVvw46ga4GL33h
DaRTSDVcAB1emNFSlc2Z5hgaxYjUqRP5QxrU3gVLVG6ZzfwB8onYjKW1dmCjj3El
ZS43l/LCyI1PJBBVAJGeEOZJzOpAMa3TY7IS1U83W/4kPuYD1eoqJokpLIX2LSMg
mXlZum1TtGQpXotOziPqS/W/r/O0fLDHdf+vqUg42F2lN0tFBgf3epwX9e6g3iKU
rU+gF2vA849HRqyQWXezB1jUi3XuLOrZkD3Ky2XZCbl5r9sZEFiOOPjrKdpAXGV4
wJu0zhyHGj0l1sE/OcxmTJ1wAPDHXs5eqUJitdbXCpPrwnoLC+Hy3y6bWp4JS4p0
CP+kQa0KBgPpYWgs3OJ3qeS9ZEd3Mykie7QF8m0ui4LXarbdbCtfFWyVGJafcsDJ
lS5jiyaKQvrrAY5KQsjtT/wUJbo+2WFw7B+u6O5GuhmAEzlZLeBZfUVPAHzEuV8U
pbIgz7+/iDfPUyP8aer3eugduTeNfOz1Z/Tx6MJ3f/9gYxNBkSgDH5U/1VrJaDsQ
AVT9oL8dHMQ5EKU8ITnsQNxyOQRfeFHnxVYV2oDHYp2WfFe0KPMm1gfJvqhbaFgh
gWmTFgLyZ/fIYdL848PibimBAoyUWvwK34NqXLGC1vapR1Ht0MSaVy7P+S5yeek0
42CXLq+6/9qitu+9HueHTXyJFfwPsMGPEGcLGLBug8lJ56W2LmuCw2AvhQiOvOLx
V3VVY5DPrhqaJecj1iQJt90WNP30vHyzckh/Tca2F6CU5Jb9Ls/bkCEkxWznUq94
5k0BdsaPqz1K1OUryq3iNurm+y0GfS4+ebfeviZWRhTxXTv6K5J3hslsNN7y7hQy
XOvRVAG4eQqRHYWSyeDCmi/p+NFXrzNfVcuoNbQqgOxRp5pv4bkVgf6CxMOp7QP/
gMRnZEmr1t83feR8hfijJ6s5Ic/5nitzbd5Ct0soK5asXJjq2H7qqrzWNd1vxgxo
n6Cdrhb1QWuyktXHbStcZeZXj9pE/Sf7jYFWnNx3kFYz4sFRR4d+bWbaGEa4bMKO
nHXlL6jEMJ1GNyq5N1cHSIGlYPCGhMAyLJscPTLSNOSCvy07gEJcBxDP1C9kPHGt
Ggu+HMjPPVygW0uky/bFlgF5EKreRZt63+IV3+corVTCeGkAFMJgykSp9lqvVGjA
dTdQPF2IB5cxwiNUyp/N4Hh2NUQHg7+3ASIrcsYWYl92Mxxy6WtOP6NcIB7N83+t
G3GT1f0HFZh6dlgoXr6Kak02JsOXRHjuMTEpWLL6aso6foz6Kpj1houWNZZ9Xlwi
9a6iBl3gtGbBKFq4SYOctSuavApzuV19mGkpaUBWDV2KAd4XQCT9CApHM3JbrDtz
9XAeBr64UVD0JLOfWeiDu6SEypa9kyLEzFEB6RnYqDRQfBAjlCuA6ngz4N1pAcIX
i0rlEFOrJggpth8hmZVeB6Gm/A74L1cMHTdyKmCyd7kew/XzivdF5vwdi2cpeuJL
d09b6XU/+1+jwowUbpUYmqk/+HHe2++Q3epsNaV1k89x3Po1ROIccU/4oEMdlx6d
WCQMuq7jwlcwxeQiuNcsDB7Hp6hjEaecmMSTqwZdKNVBazuYdrcMGJvCDU2WLDZM
D1JfPwfUtG46Z9ipgmTFzaKH7vKjvzBWyKPXULkyEC1+2Qg1xJrSbqEkl+8YYtmU
P6SYpfv10OFyiuHPd20ceOiHxgdjJNhjOfe3uZLMyBM=
`protect END_PROTECTED
