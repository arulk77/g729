`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFoI0r2aqH1aj8y2jLh939IJI521BLtEs0odsuERuZTE
clu8rrr2yWaqdGuUWyMs3t9Ye1vDcBPKDeXU17xthYmsOv+I4UkwbUI/PWVhi1Li
cipMTIxPEE3qfM2FKXwPRXIr4FeNf3DHSxmbZUfkpP80+9QcagcafnrcoskBPAne
O9Taj+c+aa9Xk0yOBfob/A==
`protect END_PROTECTED
