`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46seu0yVf6AumBMotEFQzPND652hKrwxKiRMqt9KerRD
CDHVWc9BsJP05GwG1UyTFO9+yh2fBcpxxSDVdN/2CsH8Kmzfm0n9NZJZdp9QkQ7w
V0VxhJua6sOMLTu1LHqxsqnAkdiSr5SPdFgZvAo7GclK7QZverltGe+L34Lt7I6k
3fTQ/qjVgo7k+ZLzft5ehiyC4DUh1/rO90RG4xr3Gua7sXnadhuB4IhjhIAoSxU7
veIgSMMHrjH/VB2GrpZTpGoynhc1CNJI5nk7sAamKmh+yC36JPBN9seOOKD4HGGG
8ecOfaOY9ptbY0AcQlaxlA==
`protect END_PROTECTED
