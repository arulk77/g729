`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
kzJMrtV5Y+N29nenpET20ht1Q2aqFd5yLVouk/HwtDJtm627UaXFxm1LNS6mfC4D
psTuIttIN7WC6ejk/ORaTMRhjJFQwuWrZ2U2T50E+aFb2EsUAtnzRKnlt97TGfLY
HebUkjfuhK9fx8LxSMEjWuwomUpO+Ih5O/PrtXDSTL3u+iEGg5adjEzPd2Y0Hr4R
wXGKOs9D6O5QJ8JwYy+hlt+3mpEzTdbtnUoB5TnXSU8el56FUYpmVfMwVXYG5jtA
gPOfz0E0vbfzLze4G/cxtOrU6prPGIK4PJntZ0wlC1R3ucWlV2loCmZrsuFRFjs1
sFvFr2+pOoWGPAGdQS+6JiEArlf5qUY2bfe0dEp7PwQ=
`protect END_PROTECTED
