`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNi5hqyGW0l/iH3I1Z6CDVuXOUM+1ZeZBLAyc6iT8mlH
dp0cZkG7/Xn/NNPSLePkcjT2f/6yuwQQVUWeVAUU40cvYvswFPgTvM+XKWTzIZQi
tsba3jVI/6iy1tPocoEbHN4kSyB0Q2uLZYVjZyo3SmqKy6C2QB2ixM3lwSDOzxVL
cU0yUgaqwKa1LamffVuHA7G1d4KqK39KLbtLGufRC28/oVIG5c7hubmqTTjSa7q7
cmqdGWI4k64aZfprq5kpf3pSa7TgipOmlDqv4duLRsNehCWpeihZzoU6LPIeJD8R
WyPy6FZTOXeu5s4R9b75NJHcCHOnbDIOo53d1fNhgsVfdBNJAquOdJn1nd2po4xL
fWPKDkORYaLuitWKo0K+Uw==
`protect END_PROTECTED
