`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SXmn2UCOobeXNndEFcRN3JCtE4zYNPBESBDHdEuXbcvC
Kpk4aBuOZ1ACdq1dkbkAsBSUAA3gIlguZFfZbvb1SW6zrezfauR2M/ht9mJVMGN4
RdBjE7LZ4czFsTIm4gOw8hArgEmUKr7UEDWCOS83X+a0LindLeYJ73CN9rQkxDwR
Mz1ZRjOQRpbAuzU9RWVIhG9TXZ7B4R30iPC5s4xX2aLRTyyhZVWG6vO13J43xiYU
JeVECLp9SsoA10IEjOyqNH9pFPm1KgNMC/1vRueCA/oxjlPxObQcgXaQfXGVsf5J
EyheexcDnMqJiJgs0YId5PuH2UJSgUenTWU7QpJ0GOYS22ReOJ0VHUJhST/B09pf
pVinAnr05zHIBxUQhN0Rub0D+7f8G8Os/S3qjjmbmprG59epERdjUJP2sLIaJYh8
pWrO5AxrZF61GA2hqnYNs16AffxFZOyIObK5dlLKo+DB594z1CBNMvcXnnCEJ+Nl
oOq3rfi2XUGyBVotZRbWqJC6gCGe2RSAWMCxBhkg/JZGoZXVM9yJmI5CCaNP66VS
dWG/1d90Wp/4HVpHOg/JDbleJsw2Xt0vNhrZOcDj/ucAzqhaTHU2D2aawYEM9qzx
8ws5aQRvIxAbWn2c0COCwL3bHpvxRH46ZrtRbwzasdCgYykBF5H1oRwc5lmwXe5z
865RLvxnaEd4jC3/Cofc3tuott8v4V7R9AdOG9+MEva2qPCY3z8vZjUaAKGWmHhn
IOxt+ibX6c6EXbL7Yqq7R8JC7r5Oy+aFJBaLleUCTGDPDTd/SJZ9Dxfvg/2tKmZT
qlD11k0Tn7HLYD4qHjATBFfuYnMQhkfQ+GFndBY8CdozmHGNGYCFuCZru7+F4/Yt
jDJfQaR6nLc+0KGIL0vbLvcHmnIPnus9j4fXN7OHYquNUhtda2HuhQ2kaevC3Zcf
6V6sDMdwzkZHUE2sBNRnjPa7ABJr09t1iG4og0G1C3Xt57iVURYhzvfWvOKIeoEh
KjwvEgycbQjhanZKvflU4hJZy0At5vBGyx+Ki9uQQniJa7KlNQk4tV5pBxCrjP5K
eadbYwwI5oAvMadfiszb6ajW+sfYLRoAotU037JciBX3KD6shoXIN1Wy4SZvlg0m
q61nUzNvNfObdxPqcyvxlkZFbQ6gP+s8AkOdlkR/+y6NG7C8y3lfn8GkdUpf9sop
HTVzxRqz8g5t4HelNvQL7tT8PC+kQSksNDk7C3oy1URdx8DLwhlcWF8s2HZe4eST
UDdFuXr+023m/9t4JQ5tE5jh6WJ57k0XaaMwljl5JG1sCuNks5Ml0mt7BZn0lCOZ
Wzeiza1f1EDmXhMyfWu4pchtF6AgM+IU0qvjReTWqmq/zTIjxsO023COThcSNU96
prh0ypugmdKQ+VC5qSiVsShgBYCdbIaEHPoBJmIZxxHaNB/2+OWSlOS51ljXpU+V
JIP1dATo8DpYKgih0U7aEo/mzXJ0K/L6UzI+eymo8gtj0ZngAc4Corfa7sa9dyQ6
h7Lgek7ZSXv6zp7XP6zlZ7YcSeMgv2iDwqyNTj4CJ5dECDF8gMUk4E0OpWdI6UIf
kHByGxegBhSkadEK3Fr9dJBNQZbrqavuMn5s6EpgbaPfbmd+6v5Nm1COp/Kus/wa
h+nRe8tSYIR53VSgyVCN84FD0WvvQjYgMv/kgIjRwbnVJRO6tQ+QS2mkzWBPJD5c
wGgSjlGSu8DXld736wTlMoCA18m5U/NRQFAG2B4MowXOBnCHD9Z6a3vdpihzksrC
xJhWMbtVHnnZ/0RIYxw7YnpRZNXPmJExt7x9CXh8B3q7E782ZvG/ehhGVw0Y5YMq
+WEBJ8iPtJfsDwHtal2TFAMkvW/DKzbCyP9h8ShM2CGrv+ihBKcCeB0CkeuBExQw
mV6aF9pSjT1Fi0WA0D1nA6qGWwsBcEq8pnPay9kXuy5JRJEmSva4FRg/rQfGSCO1
QNXAfbDJUq5uUmBkbnQ8XJCvjWKdtK0iAWK2o9L3q71kyA46RjG8DGl+v3/kGJiV
Afm1FK+gxve2OJrn/bcdvHRK21twTveoPRiSUOlydH3nbwE3aFJw+LDHzZig4A0L
RdT7GIplZGHZ/iFohD3zRPL89+Fcr+ZeJ4mZv3B7SVYhTiIjuQ/kAtgvyfkqbPWR
OyzXo4JqeQNYT9QyxiVZykJ5mjvVYgR7usvEly8BA3kOq49qsOom1sYuwuEEKeZN
w2eQ6RePAObjFZC8LkjyXf3d0AyH0jmEy50XnG+8fu9BjvMFH3UpmTnz8bZrRRG7
9pnvcnh4P1RO6BC2U54cTTgmFWNB1gQ7Ic1VppwdfLMTeqCicuJW0U8Wg3Ik69aP
/dHlIdJLymEXSppJIwQxxelpYMvGKaNcSvZBGrf6/HFiYYkwNdZVw6IhCqLMpqQ6
GsW+TzML5UdBcj+44vqpHbDUI+wv+/CwUdG50d+mq5lCzOi7jfyqKxJnn74wmuzN
jh2KKtrqbXllV/fmllorS0Hn3BYdAYsZMXLcxNNIp+sQjp6CwpoPPpINEvJGbLlP
EGdWie8HgUlWm/YuMCTeM766ds+8CPqaesUSqhkn5L31EeaAvvRy5anRyv4UttVg
bp03yKABKQUcUdj24Seq5CYcL7OsUiuY35WhGi/4oyxToqgd9/DqVrpZs+2kzqBm
2e47TWBA7A3iX4CGpxC6yzIwCLRf00gqq5MbfEhkudY89zYiAqmejSQGuxgiTawp
ilYEwgxKgGodZj/bseQ/mZqdO0J4wEojFjLHutz/77ZaTq/f0+ZimtU4oMQEjuy8
mA127Pc3+207V6YHN9eZFy2OzWZ24VTUraIQx9SJGFC+bewqsxWUzcHZKH88Rz9P
tlKduBncTAV62NkjKziEUE7M6ClL5F7qSc8TiNBo6yDIhiq7qBphiVyGEBz8ZRMK
xLlBSeIdqufx4h1y1JoZZIgO7UllQAK2nykKMlA2oncSo8zwdrB91+tNEl4gBmvy
ItQ4TJ8odZEf2rJmiJ+TyERPinL2c2lEZ/hV6SiLd2LbyQ12cKhWplRVcNzXYc5q
Rl5O0z/57dmD/KRKCvxjW9CqG66R1Ns8AqnZuVcAt90Az1G23nxGxXWgobMDORiv
oJuTWstC1BaIxQieiBD9GdBeFev0EjKY+S/HvPDjCIPSPvx7oOUbpZTr2DSL14vp
HEgjgIrB00LK3ii2gg++WCYvwSHYh42O7D1IDskrKEM=
`protect END_PROTECTED
