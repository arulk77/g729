`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
LWEvlzVbOOad+7FY6IaMcBveRORazrAozgPMNNnsPXCnegRijZDXQXkkeWlk6aKZ
0rVDtus1/cDZ2ExCaBzWL14HopiQ2ZwwSzBaDzTBAMQj/gfqVtziAzUYQ/r4j6R5
fWHDn5ocBh+WEnXFzymeReozRb3vKZW7clIcD5QN6MDoayiJRA3zRTziaqBES7jN
FfWX4xNSRbl+2ciQFL+GP/F4ouCv2caEfv4zb49VTuxiGevLHEaPIG8ZbzKOeh/G
s9GmO3aasiLD/MLKnxmIXxvI3MWjQJif5wHuw4SCX1s=
`protect END_PROTECTED
