`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFutPEsp/tzkrHHjOv2Hk2UCtNVj9XAQBZdiX4qOzYhD
4V3Js01VHrnjPdeVqV1lRuyyhsae3WGRlCJMNzqkR5DDzkW9l6S7RXsYoRWHs6oN
D8s2KWr5GsdOnvGFn2mUhYs1jbZo89o6NO0KFuVUtnTltme06Mdu3H7I3laZ5k8x
qKmUm/9QRHrpKFSFIbGxdLocN2TH3sWOSp4eUGAXGuZQNOGDI/XCBAwD2DvE7yOC
m1VuhsGVaTt0pmJDcdzdBfSStJFre6LvApW5ggwsQ9Zl6sPRkeMhEXunLFYXo3Fa
Ia1JXJ+wD1K0RpgAwKAXug==
`protect END_PROTECTED
