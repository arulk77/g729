`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42iFjURvnxkHfBBA8AbTtgwZZC2N5S1JfCbCFj7HysKO
MThVDWMOkwiZv5VfUJMWvGah6C/Uo+8Ev7KjOFQiQMOlXrrgoGY6N7Uhso7DpXDH
3XqVguhFBmQDni1qDPzvdTsMVivWEx2yozcKxel2fJrUH8kRuRYTAMnY0XmzqJcN
Ngj0WP387LqhK/dCqpdYRS8F9TT1h85rc2h+KKVkNySbcbQVxaZkXG0e6aD5w4+E
3pMegZtlKBVmWJm7pR8XTA==
`protect END_PROTECTED
