`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJzzUTKplb9y8qGSMQRTfX/FTGqcjdOydId9eERZkiDD
0OJKrYaZSy5WMnQDPBsi1ZZ7JNv+qaQ9dR2Eo5zWN6FeigKECc2py0yy1YOgunbU
SO5fF864/jTwd0Y55yRaA8zqQa8QHqH0gXiiExOTeXA3BJ9i07rljsgDBu4jVsuZ
pPTXB8NTk47mKeo7mr1g+WKtrljOBxlzbATgSbbCii1uOCrf6NCxa8/Aszzk1glP
iWrTbnycI7/DKBmsLAtVvV/oAyGlKwRsgX1DzvvgqyLTSK/uFlCNKETK86RzMwkh
bl+r4xOzj3GYyAE7kCQL9JJ7fKHVRkXngH96QKos4ig1gyLCw+fzei4E9fMu3X2N
EXFdMAXpOKihOxpTqXy6/BOV+ImWBFym4UwyX4NLS5pDn0+OFyUuvuX3GZEubAmE
/RxixUcXet5qY4IjQ1vYdw==
`protect END_PROTECTED
