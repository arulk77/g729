`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
OnEYI+xH8QkeGlgd/jn48Z15ncBVwUhnEy5OU0IPmzN+32WqgfrLca9jwH5yQJ76
xleRAyioevOrm1gmomXMB61su/qUXk+DVywvOsgPi5sD8pvCc0Zr9yI23ceQY4NG
7n+8RqQKbO/TLeKBNKZez8FdBjzDGzgdl3h+akeiYr75V6ucsjPmZ8nEKtdQVLJ3
A0vjV2DebmtIEKrmouzF3gGD4Wkmhx1I4C8TtC58hTCaocIRDFfYIfW7El9I0buq
KWAIKoDCx+WX2rTaAkK3Ir0oGvOAbz2BrvqS+b2m+p5GK2HoQOFsqiELiaW6EMSV
k0ljiO7a/kjkit9I+yOCNXj0XvbDfRAPpFsl5Wt81GNR2nWaNziYGlggROVLCmXt
lQIp0aGIrYKGXkoo9vKfgolabLNqDXFS3YMzs7Q79EiASjq4Mn/NAIe8ktttkDbU
tIMJaco6Mh6T8QYtj5gauwaJMrQNF1I4jgLCHJjsutvk+7b++0Gqhb90Fp0ZmwNU
IHG4zGpyt8RpZjVf/ZsQgBUGWDxmxpnUphGHtM/Td/c5CDVlmd5q5rYnH/IPUuvV
VbKEoDoKRCgvObgBe06n4sYROo+eXpwL8mZIFamSXnepmAD7Nx1CMhEn468anbua
GYxIRFuHqEFAmde41y8AMA==
`protect END_PROTECTED
