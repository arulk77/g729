`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
nxJgektPWNiSRvYtwqrp2SqtIZqMlJmqAEwfeurrxxM2bsSlRrnUao01uod4I9cO
0dkpOXJfoacNU5a+BzIALiiFW/Yn+gKGVDQo8dTWRLiWpADniRFppf3pdqi3F/RW
QwPyg4/8IR/+OyZ8BeVqnX9aI8+TudAtfimLXwy0beg=
`protect END_PROTECTED
