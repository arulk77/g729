`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
GSPkFGlT+/MXL+LylfJGqF3yIQIUVDJPU10SBXh2cmm1rIQURYs5DJPsN4R23pd5
aaf76IIvphZfv1hOAx4HZdQAXbs2w4GQ+UhXFy9w1Ww1jb1VhhJOur2mCBeVHFQ2
ScU3ZKXBKsKUhGFYEPXO7Rnyyg8BTb8c6s6O0ziQo5wcsovvsJWqHO9RBURlxThN
SLpt5tZLb75rEYpdwsnKRqeYbh7nHS8Cki5+GurymKS8+OFEKjGPJkgdrC2k2x8w
lapUYkRxoUzzVwuD236YF+JWX+8qDaSTPQ0CriQoD1DoItl3TXhFunawMSx2bC7q
C0MpDcGWIV4bdUAajQeN+Leih6H3s6hYdtRHx9AyFgc8/dWzFEjV526Wdv9cBNMm
U0YPjjEg031SHc+2AZoT+0SXuW0It3QRi85ME+QUoWQGJtSPoqdXTArrSJJ+VD8f
DkFoQ/aBhqhvE9noTLo58oPq9gP+wj1QHzXJ35tlpcROYzf5dOTCKHT/3Z7EfB15
92lbGLTGWWZXhvGWMM0Xmiy7x47f0U/m284kUBc/iO5jqDDOa6vhg3eX7XuehSDr
F37JMiikPGijA2y6thB2FBnYC9JvjoVyQZ4mcpzZyPNvjTT68NnFsad3eYZrld0h
4y/LIDPnrLYCiQ2cYOL9mhwvBBsoo5N7K1WiXvXNqSWfF4BkeYBxsVG0KGah6Mco
es14jCnblyOpDSo/UzlWvdsgBDGT1VOQTv6eYFOfO+jS0569QPKU2qDlo8hCmVyC
OjkpWj1x8oaFimIrUsTDdGEDX6Zv475JhJzMWZaTEFira8T0pGisFtUeaqZcohJr
NpEzgL62qOAggjfDOXW7vXTCM1CQ6Whc57T66DWjSs8fvvcXyfK0iK0dtu7uSg+N
t6vhytLyhp2H+XM19LtM/ql2d2MekFL7ab+T3HCmnuSFm4AG62DxvmCk6nXpbok2
UkFv/NXwLnGae/FX6cEJVS3CKX9knYfu3cbcO2nvyghRGGuxJuNszEk6uEU3Qz7k
M2ax2QYEzsS30Fgom6p0zdFl/ZxJ9XASaXa8QFmEzqbY5ASMrc4tzD/ppRUOTLri
CC/k2yAYglyfZ8ZEo5JAPhkpE1ijjAj8WQy62DLaS+DcxfFW2chFunuZTP9O7nGK
uFhOqYkKqZsLUd5+gNB+yklRfloUgsirfcCNDfaebqGRjxqu5S04sDdzV4RULZaH
XMQ/YSCH9m7hQdgSJpYnsvNm5YqstoTcCRZr/cHcZkQUoWQYVLDI63mM/zM6W0WC
oBet5/MP98VO+jZ9g/PrmQyLYSaaOO8jN51RfQEA4LQYXavhigvflMry9c8F5IUN
0unRUSwI7oArRgWl/1HZhG+QyKtenRMtFQqpaHOIkd+h866LLqxE+nslDiXu/Hqs
tEgrmA6FjLPJ8GBanuk0UA==
`protect END_PROTECTED
