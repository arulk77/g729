`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNc+HICpP5aWtTBl/Id10d4Qcqd01bPKa7ySMASbO4lo
0b+O7Ly2uZ/TULTHdBpSSTdT0j8bbBzss6fLZ8RtGi1FncXHmRPggewJ5iDlgJY+
3x5BlIR5i11SKi49eOZWNbQ7BM4FmIGRTa8am37ijwa5KifqQVIESFChYH0A8p23
WzLTOEWButNWX9BTtXkXYrt0GAIzRNFl1wRVfGC4JQuuWnLxe7pJYjUlsM2OB9+0
zNcap8AB3h6iEAVwknWixw==
`protect END_PROTECTED
