`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Wye0EOaX4JdPJ2gj20MjQle0djE0XpIVckyUX9B+mRqRDlAG/Yp2HqFSC843UNm0
nNUoyrd0dqv3eL+l9uS2rk3087vvEk+6hWH9zAedyyi6mqHYHyqp7EX9ig+X7TCq
innStm6SmE0imEkQTrSENfVELvfzR/+jxdDnPadjJcv0hik4kdWBAe3AgMMZVBL2
9IpBuWtUgoTjW/uhCxHTnT2fj4mlJFMJr49q/yeBjf0=
`protect END_PROTECTED
