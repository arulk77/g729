`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
54BCoiLGyoUYJNyZwlyfWk7sjyrOz+VCbkonQtc9dYwOcHuye43mvTTAKOfTet4d
8/dWCoaUyVICBr9MN08MczWVTIMkAfF7F949qUbrGm+G1r7toI8Ez/IUbp0IgL93
8jRIwFwBNNn1/DlMGoAgfBVQESLZpUlEodVn2XQW0tMtOMGbcIsdhn4n9Ct22ndt
Txb5wi44fZSKa9SO7V5OddP6gZ3yG2Zb9REeyUqHMr06tw/a8Pv8jVCXPu4AiHp6
w+stvmPedKx4Oh2RG4FIogly8A2tSmV+AhIh5jfveqdNvwx2PcsQ5L2bTh/x9t33
f8wR0dQJ1IO8BzkCwFClc4+RyAyrmXoeiNFKmwKfvqkSxfJm3LuFMzUct5Kk3QsC
wh9cDYZFhoaG4yxXiujPA3CPZHrCicHNX28mPfQ4iBA0j+Vh1c1pZAMtLfoCesxQ
EybEky/GvZcx5OwMwJMMbbakV7vHJ5FGGojo6SOrFr7y2qY39VeoCNhdiYkYHmtT
yvXNj3Yq5hkEdF/viDHKSE2gj8WzynqF8o3zEc7fbVxJd6Sx69pnc2k6n8gIqmp4
0vK5qL+zbuRerYic/zffDCaPaRsT/VIITDQYYJNCg7324vx2QeygjFoIKVkAKh14
t6GzC1PTuSjc2/HkFS6OcSZ++FWfIYHco9csFxc5GjTQcGKwxrrCVQ0P7Y46k7Lw
jvZxqWkxx0FHQHbPzgqRYxSDeYal4hhnrIwIPZu+nLUXsaTBpdu2itkqxVo9iqxC
5MpdtTUEb3z+K9aEK9yXO30crnfB927PVZ4UzVJcVBQHvudNg3B7r4yw0+dXpqoi
5CeYHxWrKcYnVdA4yfLvSWvCVcBjSgXI4x5wj2ROmozPEhriwK32jMhfwiyto+at
J+28pU5HYeahW9EIQy3Xc9TL1w8/p+8Jne9t/QcPJkFnLqnldtZWo1tX8yvwECWx
1llklEky84tyj6v04Vjyzx4/iWTW3F7M5JseeM+ELc4peoRboVkMy8LGlNcTGTSy
`protect END_PROTECTED
