`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN4v03lv1CU6xwNlZTKMnGJ4oNj7XorVjirGgU1/CDgBV
yuRx/pI5N9ymTn6VqqZAk01PSynw5gwA0Wf/uULNlks492D/9vFQXBP5hZBPr9m3
sYK5t+KfEe3M4hmMw3d19a0hH6h9qj7rD0/m76buNIf/e+UsSaAfBuvR/tX0FiYA
BuHnqsRmnN2/Q1WWDCey/K3o/TWhk6loLufzVF4/KQ9fBVQZXi1Hbe9dz/tW9EZY
+iAjWBTg7L0INwA24oiFsyF3BZ95ll1ad2l1ZgDEKjey8uIyf2tulETjsO7YmpAP
Zxf29v+7zLcIG6ciXUl5BvEf4nXTQxvJJGAFuHMJdnOj9NvfHY39Xnkht/NNs5gz
fHP2BqZVBvDdlWk7SpjiQ2OtGrwRrBL9c/zS5XJ7+ybxe1QgDhQ8NGUbaNdxsYe+
OUvmYrAyZbPcebGFq7zjrT0/LNX7NHGBNMnTj4NvehpuLJm+FVxQEicpgYAatXFE
+EA1Nw/4y5ahjkvV/beVQu6N+Q3XEj0fOtbwrG7VtzbjNoUj3SoFfW+Y1FGFF0h2
50aYlPr5NvSVA92ESjqqDdxnKi8z10iGoVyt/6IrNi81yswLOYz0eKKTgKuast65
kgOpbd521opJwgYpEqK1i0tWrAL5LZ5sFjFhuXwUvxwS2oEaPaPZe5YvI2Dm2Ix4
6MeiwXDfWXhU6nw4RcdkZo2IcWb4ooR5QdRgbDes6nUmm1PgrB7AuVoGdT7XRjwE
NGXTn/NNqBsfAbQz1C98S+KuE5JoHgP91pu26geR/gx1ABtytamYpiISXoujEQvy
DqcSUHfeU5zHRfT3I/NlZDnywzFCzmM5em6n/NfdjVKtCmpK88HbWIK/w8sFSzyF
uDNXEJmZoC8kYG3RtxQY3dzzLTzdC5FyJWkpxuMHJkDqmy18/FWsrd9D6Dwgw7kq
GDLLpHOvStTonMoWWru7yjCnOEndDdLwU2RM3yVSkQHyT2plxIbg9BVySLY3HFM8
Wj1CZWH1t5/nHyNTBoRb/Q/xyiOw+V5HqVTWyGCI4RdutwzJTs8yu3V1V8rRLh7d
kPzGcdukD28EpZ+X8mWsVKIp74WfT9c2NVZN23GsDpnIpsPC/kso+8V3Tj6gQsos
hP0fOexFWNK//UQ9/9/hR3YmmHJSg55AYVSCXdg5JVDYJD+8USuGGuLeO1/8ieQb
InRgKuiQ9tAGRSuAuSVdvzaetr8O285WaK1LqspxHP4ulXlHN0xBYu7t1KbNLxhw
ShoGae9h2J0dpyuAIEWBA9imzbcIYyb1DFOWh1F+taJd4uJ0X7rdSTnfceDGf16Q
xpcS7L5Vl1pHLsM/tYfdyiQIAa7HigbiQDyG+GmVLPJ6ew+AM+dfaftzgXi/RWcV
iUMzFli1xYBowb3/pZ3SsDswXSq0V0P85wmElCpHs4LZ8tIq/kFmK1fx/yOdCEY6
BUnbKITZRRpKjkLw6hELwkyXjgKiJOJel7osR85eRBQyQb6iPpm4Fwwa8iOyqkK6
2RvQMUg6WEdrYz64L5kw78/BaYYp7/37ZiStqmHpAaCxHCmTesbp/6lkXq8Fcdjm
U2JcYmnHcpnabmQjPn0gqNyaB+7tbExr93oX929muFc8LiJ46vyK8m2RXTxpxB4o
sTF1LmbR4xN6STO86hif7m6L+Rgwxe6JO6PJXGmFqjM/OQq1w3WsspHwXKwgER4n
FK1jj6GHRi7HXPbnIpbzn0J0UeoakFlcETHS44d3fNgKGj/P3+nnyHoHlTXWR3qw
BWHXWwZw78MPCsGV7QkuMvmkNY487DnPr9GTdAgVBdYXJRLVQUiZgtwx6gIEv/Lx
6JR9uZs28ZhOLsXjukHDOVTCGUl38gr/nOsOwiiKq034Q4rarWpWbkJGoMa3oTc2
+8U27pDi69wz3XplcGvfAd/Sjfb7gNFxGToEghWTJFk5hQST+wbmzV0gjWw/FvPD
dYBN5cv5IFQFf26AYpguGdCY9Eh77aMRKxFSYCVyrKn1HAXK+x8vyQELjKIzAdYM
OB0j3s+S+mlhXzycrSjssV/3WISTBZu5iiEFQlQmld20ir4pgfMH97N2gvBzGxAI
ZkwoFY/EqVxFwAwDHJ0FLShoxqR5KdqS5cMyrzXXTfGgdGwySjLJlzXo54O4y27Y
H3y1tNrqR2bDyN9AL3opm5odWIatDv3Z//J2JNlYCB4t/gZkYTiVknKNSZrEvsbt
+T3pUunIp3PwYB81DjrtNY/DlM6ah0gk3QH7/XNomZCQtiRJyqk9m3Gy1YeptLJ9
tmvuvq59cpVZDoBPluFtOqAOJs0QM7UmBR0PaPrJ5TxPVEk4e/bRUWWFo3rXn7LD
wWCLNW73jOC2xGKtj/vOhBuwI/R2q6zPZYJxO3pRqttxtA3BCOYNt8RuxvbUujCK
/5C9s3Ljp3ZATMz4g3odF0QZjG8E4yVOzPe1pCKG4ZMuNCUocgDYwU/HyNBpVRsk
7Lf4QQ4GMosJX0XRd68BREZ8fj87c2tvZ0yckws4v27O1x8GIdZ7w5FiD2cAb/Hf
i2FzXhDhMG0ctdc024ug3B3ykm7lCvaCYQQW/rqZ4LxNvN9noIgPSljHLKj8mjgW
yBK8ikjJv8p8+KDhSlBWp9pdCbpjuRsSWjE1j9yjkNYilvTgD9MztFZV9HG9L5o3
bHACX/lQD6uYx86jnIHptLKbxqAJbmuGZNJ4SCfrrvT1NyNbPqW4B4LCX9d7SZWW
SR/OLqjmU4me+vxRYB8F5zhJjr+uoLnv5ggPRfVuqtHkxbkfm6FbErhUzdLEtpet
hNl7kDuDrBnPZGmIh+ZxSC6+lXYcORUmO2e2bVZzpNYNjE7faVa1yLZR1I+j7l6n
K/HIJjLdUoU20JCzyc7ydKPOuUhnV4nxzFhYXCBDrCtz/qXXC8eCjmaa8po1IKou
Mja1HSKrMW3sOMpWFzXqqh99g1UyK3PnrlCzel2rUT3AT+Fo/y2sm752ja2RCJBh
3LCpM5rXVuZVJP3VtqD6R4P68ivFn6/y+9hMTp3dFGvt0ipJDixQd6LGKuiijl5V
RC4htJfkvuAtua5Mozzh7Keoz09wjXHTel26nqGCCuBehZtDfTdZGm/2Y8rgLu/j
tXZNWHgpowD0yhbac27HzxoD6kQj1Kpj1oo63EJ5eouhnBwdHadmCv4w75J1ZjXH
gfmjBMqH1qtp8lAswnKE8ZtkNM5HdyOge7nkp13YqeoIipKRwkOHBiMgMvM7x925
ElGaw22N+cjgHFw+813fZLaI96VdRY44FXMigYwk1wSkwsqgCfj1pEK97YJmb3Wt
g/XXsVdRNtgixeFFjVMtlKrvjpRIZ2Ue63Jc2qNKTJWrXwT5rQ9eYhaqGuTdUCUO
wOdvXEj52JWp47b0pmQGMCvINHekNR+PIG+PRSDzVLycLbNTfuT5A+5A7UQcyrfR
3kkchMp2wyj8oyZxac9FG6U15GvATp8wWtHyDbdSN+cCc58Yc/nMozE1AQMvCDW6
YGnuus9SU5NObNmYlTw+SAnENW/h7OrttRrbwdMU7SfIBbcDGXEaCCqKxwcFdudx
IEWBFIf+1mxAzxtyJpvv5xzitDzIintVolI87RY/xKF6+PEiQpNfnOTJaapnRqst
Bo/HF8a5QDXvlJ3sAF/lyJ0HCCzNN5yXC7NyrXck/sFuiemvzripqG5nBcGBCCC/
5DZgHCqWAkOo+2SL+31y3oHcYTQZP6eqisBqmvDrQk2g+5CfTykBUDdFimtJNfCl
NYhAa/8CqXXIa5bwyXWlMABlX/21362ikkOhbzBmKRGSamQTKMKmLDa4Fik/HR1I
veITF9curxLrNTAnj2SXv1E+K+hCU516kYcjE0PaV8wArOyMW1T7MRbenuyroArt
JWnGinc7Ff+SwGyrSmEzfT0zp20TP3zror7Eaucznxs541AYY+g9mubk1vCHMbI3
qi8q+O8B//8KYYDUxbznvJ69vZDZUdvdfJMWO3Ah7Fhlrw5j0nMSHwEa5Li/nJNc
qQkmSNQqYilf3JWAYCpuUMx5KeFhlhwQXzeWIzRKuq1hZAY96XqFWNYNvu2AFCtR
/3Lv+hQiOsvsnx3qzws0EMAYyI2t+qHATqSe38B+5mlolvvq1tDEknYaAsKw/kjU
VTODRgkS4vsY8qg9Z3MHOvf2YMDvvoaZTQlEoLXOb7XYZm0buuQ0fW4ZstBgxd6G
ZJBT4pXRUmkuG9D1CVwPFjSeY/P7Q/bbIenux9RGMyNJZ/WCIszJxQWu+NmJEvd6
EXCiJCENfEzudR0WvlmFuve/LykQu0gmFLeO++a/y6zT8FOABRjDw3Tcckui9NFO
5H0wvtHkEHs8kanZ8663fomr/kif99F6E6EG7bT7U22+VFmJgdnMdDx84BW2BIcK
d0P509TgWgWfz7QB3F4jOUUPYX23cKGGZvtDLIa0ryjWBDvD+uC1d1IFJMZxfEOg
I18f970/dAd4dwykpzzPtXAL030Ezo3MVOVCxDup7/JoM/IqxGj2/FtoXIeuemnh
7baQNJ+H6bo5wSTIMmRL8JtQz0SicAWGs0NVNF7oAVjHL2pYKSF65hphcJRQinyD
jYs5IibN/sOr6R3Js6oG0GpxC/NctUPF2/i7nH9V8Afot9IB7hZptWAfn8DhscEv
SfIVaQyBI5jDbjTSsylwUpXY8kFyWLVPwQspV31OxYInhdW20vAkrklh13BZcOvb
8tRJoT2RpGWvKhnO1gEwpa7b0Q2jC6uoRd96ouOdGB0CW1xU15XHlwD2r3zl4t7Z
yKEpTa+D4eMHZvjPrAZx3fdvljQYUfc+easEOKj/8AwaVgCg5++IbntScZXNt61v
JhW26DLzqqxhMAgYApoV8qSQAnLgenAkNU65P5iU+W3KmfEVEq9nhuQKMfstvCq2
m8M1dW1Vc8WR0wZDFOmf6Q7TLGkKYZxFuZ3Q6mNi0kW0fPpoQ4ZuuVLcnm8H3vXF
4asIJQjq5Gf4RvdlbQ9nEspVlMvzUTT1Ke3UOVaTT25do5w+7JbselYZcr92A6cS
0dDM6iYrb4CwwwrmKSAhiZeqEwUxrSyYSf4H7u2eewxLKKCEA7/rqyNfVaDULAwg
wZdZMxz93Y8Hiu/57gGdIfw8BzNtntg0Sh+WlZW09pphq7pwlwZdzTs6QAUg3/oi
AmUAvBvisR8E6/6O37WNZ/nWLi0lip35JWwyywKPEpJQegZyiIx3lMgL3qbGh/K4
2cEgYQT7LDG5wOgyRI0dbSagEO2LjSuUR5bSEzBt2ihLs7g5hWyyy3FsE6KkW5we
jC284fnNd5Ct8fct9a9rcDSW+WtiNIyf8rIDyBDQ92AuSvqRZDn/Efua0XcVzhWy
xTe1vUc7vLVKm3Hj/mipnpzl6edAilhirNiZP1mGUWgXQioIYqmhvaMTkvay0R9A
R0HwWb0ZVM95AWaV9UI//yMcDTY8JDnnHxV4s7kbnO4RON1pZEqwDsECi0iuz7Mk
j1fjE0Z4qcx8a8vWtFnztv6Twlqq9SjOEZnaxhqcNvjF6uMCKMTMOOKURlcZ9wUo
TBN4p1qEXl/RgpzkM16MYkYjhafKjB+sKynIcYmUWbtsPWEFibDAnWRP9afyezd0
ESBEoLP8KPAzNaYrTfDmFggWZdUhvhqbnToAgE9QOt0ZnyA/cGIWqrGtyP2YMYXg
UPdP2+EXwtj9s3zJVj0Ek9qAbKdIfmguBFKccow5CWPzovjPmMUm2WNjvMUlihSB
ceubOKUP7lVC2erc5mHD12DZZuP8+O5vGfST+00CyAuwtXMXxuROrzbRwxmTGALh
SHFGl28iGvY9JAXhIBR8rsfK80+122SwGP3tJ1XdCiQRILeMLLf/21V84SCj9HJS
cTO4aRXqdVoX2/lnjLAFQe3luGvdEJia+CkOXsZ+yNuoy0K8TsnXAVz48ftXYu/e
rLKQ2S24N9/cl7SiIrNQr07KpoWiStY5F2PGIGwTq6zHpradiEX3x1riFE6PJlwG
q/DJHt5OZiWcefpWLDO4LsmeGgL5/Uj3uYJ6Gyhdapkk+9pntHxQmS92ERfUVu/i
nBOnvlkDBJ+6fFcgg1BITnoEcIeweJeShMi2u1pkd5mCET6Q24Mb438wsMb+5Gi7
8MPdzDCiaFKF1kPEebBrtvVXxeTaW1hQQYFpjMOp2cDum3CZuGJFxzQ+QSRN0/ip
Qrso/OTQYr9nL2lt1eNgz0p3Ka/evDX8EiRkMfYTm3Sp79JP+cVC9+KsYnl81bv8
HEy1I/HlkYjdxJbHy0Vs5pXT7ISU6Php7TyyWvbzL0HwKb3IXc04UBVNxFZR9sgB
uVMthQsYkywHN+ra3Pb3l4ggKJqk91XR0Fbhu1fLKHfaTGnmIqBqUhTiFEajvsZx
yBaHPgmT2TABWn7C61oY8MDgQ9U6JhDFQlPbU+S3nLoZ2ztaKAhztaAWzZ+c2TVW
REISQZr0R+9bTxHIdUAHlFrLUWjk0eA1wgAUAkjgq/XVD4S6iidg1pBv73ru6+ad
N7oaqSrQntow9soMzrt7/Gq+LJtTQ2y67eafJW9++Zwcqd6Q4rw5yVYvWvQB4JMl
9nolxmwBJ6HwBTOIN4cbxiOeiTiCq8j3a+Q8fMJozxbx6Fs6lunSMl29VFjb/VYD
4S6ta94fPpU3w2UZCayhkPa5CQ4UVycZlPJUlhGIc8s1UR0/wAcHjaWk5rR0RuKn
eTAfLQajc/UJ76QyPffqyXhchHouoBIxX/zyk3E+G9NhMuVzsyiNyxy0x0u1e3qC
gSuf4XP094OLjPqf8u6BgCM4e5iNvicKBCCTZ7sC6ZL+ywOgNERj1wBoFBAokmPJ
KhMNJrZj1b+ChVl9m1OjifslOOFXI/5TjzZ2CuZGg+B+0fEjt81SLJTVmfPd46O0
qdqTZoaqv8AQuayF8lAVY3PsWdDc6VerBj2tlqLPA8xifFgJMtzMBis6//F7ffj2
6lsCvwGlb+de/jevPCw1ixJmoFxIHBsVn0MjgZleX8oDxtzhuyEhD59V/xIgyTTF
DfyFN06M4+I0HmMnwtewhrlv2rs0CvEKo7/AwWRRhI+GlZMvgFMFVmQaTd11yfmV
/wNgap1khBqy5T2r3/8QFSUppPBWlu+cDy2oaAw3mitNbGUzKMqevsfOGx0bGNF8
4pY95A4mpkFnLe5F6bH9PN/iNyYdUXHezM04oCfSz1Mb+FvVRg33lSnD/flu0+Eq
v8QRALFdc74ycCuPYTIq/Q2psfmYloqxaf+SpzCWxWE2+4/8yIxM9asGE9JrMg3v
97Mx2c3NbmT4yjhOTZOr416t51jHHv1QNKVUUkoEQ1iMNA7+xZP55s5qLi/bBnEF
cCiHCT3MhsgRCZaP9jrVE1+vBvUZr9EZPDsAihumE+QkRJCy5+vsAHEjljWVHzHw
Z4VfPQpKqiG0BKbgVFEdPDMHUxK4/xxez3Ae28SYTzJUw8C1p/JOy29TioIGg+DZ
7UdCHvZdCJ4xOnpZFIc7WADFKNv7PoBGx4qozWFMZ6jcZBG69ZVLbM7Z2YAIy2Zy
doHQGZhv6zNoYRsTYliYgf/uMqZ03EIOjumBY5HvTZLzq6S6ID4eTG4iWhmHJFKk
LwRnsC6vTaM6976fGG7XrLLh9wFm1enZJGWAbQjOvRu/vUvCpHPOoiI9pIeWZs9k
zvOQTAU5df0yEh8geC7GlOvW2CELXTTQ7iqAi7guvQTkw0ora90We4nez4z3t3L0
hZYPiBzwIeYx/RKqf8xjwcUd7oDJ/O8yoLV8Rb5imOgA22t1RriMA7GXJaS/hupu
xLvfKm+/XoJ0fu0l1N6iBtMaINkEDOMVneoyNdAxrG5JFXK8z3xOcFygoZhFMmI5
BvHeluB71m4EX/yh+9ObJo3fRq6XVYSi0Uvya0QMbDwMSHFLmWuVvt+ogyJIqczN
Hj6cPoX6fnutbL9Etl6co0xAhnGg3s3r8BLjEx0i4aCJRqth9jpmjIqOQJbdaK2X
MCTTVmdsRiM86BmNNonLSw0iaE188XR2bjFu6eG2vU8qq3CGr/LmEZ3EYtPhsvFT
6D3VxCBL0KsQ7A9J4YUocCHs8sVlG8rh2NBTP+XMp06aK4HakfxqipaM7AujAsyO
zna0ZeWA3+uWCTqLazzp4lk22hn2H8L6l6/i9VFqJnR+vKjxW1RsYzmkiFMvxOlx
003EEVA8mw1rbKFIXqJHKwMMqPZa24HkJSB9l2MumuwuE82ln17I0HsLXHZbgKsz
EhBx3Ofk0Tl1lDE+ccwQgh2PyCg90b/gAJBbpq4oc0hWkhS+8cyr7K6z2AAnvKKb
/BV3I/uCOD2SP+YrHX+1UH7WwaZnjabrR3SHT2K2fOoELCoXqOTv0QfgqwCLwczY
qwzq/iX4xpabIYm08tH09PDKTSLoWUoBZhUogXDj71ANsJoaJ/I45O2AADdGeTYD
HEBxrv6D/fuLCiqexuYSVLwVqs7nXQQg46+6F+M95iAtENH/g0wuFwdkpVjxb/AY
DmL4RfOgNn0b1F7R6V4h/+PgmGV4uW6YsA/H84ozWuFTf7VT80Q8qu4bzF+PAfo3
IyMs0/wps1r4MmgEshKrs4W9bVwkoduXsJxX/S59NWcmvzKDYhkOy1btBYnKgRnD
+xrZiytDAcqabt7WQONemsBp+WJAdPnZvcfRns3OG9J++DSdlmD9rGJ2j8Vxl2AS
I2a7VFcNJuuq0KD8r1iVcmkM5q9OqdbzFEVIsKrpo4BbQOXnb9zDy+Dy1k68ufyv
5u/R1kgjeCFhPknpw+t6KbILAQDxJlAjF/pfz0GAmsuu3xkURZcZ8rOkgeI3PdgA
FQkjkc6RSFT0c7NxaVNQ4g+gJrnIGUp0fKahgX74QCxxuoleKcCjAjuqAogXXbdd
EbBJEbSNAgNDzkd7KNRTEXGZOtI7Z+pKt5amzqUGi4FDLb1prBfRqAw9S6qMYmai
mZfyxhTLNkY/RGi6h+Zs21HWZv07/qzyf45zq4kteQeWg00jndaCaxogIs7j5IER
jfk9gsSv5SSobiM0LhKqiyW3llgPY2CSfOCJVp8Nq8n3CZPUVUc0tnilaTLKzA/H
3z8pVSdnaSZ4UmRwVwDp8QNHspfAPj+ZesYzcaVVENlzMxr0rNg5zf4ewQgi5euT
5QNRRRQq5IocHvZJPuSLt6cnsj/PGtF5rQY/uXRNn69Jq3rYlU8SjO3wXAEK1gr9
+RzkzTI4qmSbsgv5E9D4C3Mf8SrCjMfeAXNlrrzt63h6SxBexqmi5hPEWtRZq4Kf
OK9TSNbU947SRzGevZsw/ut9PC/V8DAcfb9+Rq0JpPxxdMWV8vj1EvF3Cqrg1VWB
z91PJwkCOV3NDESEOvP6vygYYFxTErmqKQNst3dmAWKY+D+dZ532TNneKf/SfTIL
r0m1iiIHK7diO+PUxAQ9ndulmhlFWpiYbqzI9ufHkSgBnxu9FvjeHlPHhbX2wxWR
Mbm6fGGsS9+whdpYY8qwxUqzlC+OQjN1CH93KGP7/mBnR5SJ+r54Po69ODYN0q6Z
s0rx989pzp4xHO9a/wR6oFxM+9DJyVgQW59JnfgAhaci80ySQ1p8POzBgshTgWJM
i9504cdJTeyNG9nu6/gQs5ulGI/eeZvthzHXw+C1F8yYnYqZeNChxZQ4zV90Kb1B
tJHaRkDkfTiQJ86foB/l8Vr2zJ8hKsK54N2pvQnxndzBP8NsUbtD+K03Bhi4LwP1
tFnpKEQ0F/i0hCLVpq3KWzscYG1RtYnfCSL7VkaX5Pl1MMOtz08D+aY0KjaByMxM
T3FFmE5BX89ABSDoNqUpREkEAKx42WT5m3umkjCddpVnjIe5XFrZoiT35bw0h97Q
FgKDSvssuPrPcOgFY8XRQWb7wvFj64FRCMROQEZSBWPaJMZV/gdNqfa6S56U1zfY
jBE6cYLPuLDn1eh4lkkP1mMcN2ToWMWxB2GhD5rqvj2McDKLl8EjQV0rq1jaPu4a
4GL6iTxcLNamBjWdXKfyonFAnORRUuQMupktfFy1XfuIFcyTjlxckAkJ3jebhDpT
TLKJwBhtneKpAwJVgdjuQHPwsDjOLmlibUx4jdQo8t0VeJfmFWZOMj1232Kaj1dW
GHduMMBHXM5cLuiDXtBnMfuGRjZB89yT9n+1n6oI/NocPuOu0fjuMv62xfOATi6l
Y6b/czlYflzMHAeB6AMGWzgIWrxFiVnPWpCZ4D2V9YlzbD9U7L1Wgtoa3ISZ0tuU
w5xwfEgCB5xpeGlPquBAbC+3wQj78mL0MAbE1yeNWCQ+5I6dnZLR2n1xnralbqw4
yeh91v6L7tRDTo8HZamrSbIZLg/tfx40CmTJaoW/J57+15nvIzlW8eKn/8kIkukB
BAiPvwQv925vFbJKcKhZotDgI9ohm+bExsK6xbA9ykrdfAaDY5gylfPUQMAhkW1O
nr7ItY5jCjFHJQCgIpsSToWdnb329TM1dGKaYQIehPj/LO3TtALlQ1w/jSD/GJGc
qUXuwkZLzDoZQH57cibpRlpgG9BLawtL9Rg2JqYK1fapAom1fxjWBhOj1v8XaZg5
ZOFWGqZNAYyLrt6jWV2py4IFBwhOxV3oGQhryHizPyw2etI33TgB6p85BjUJZdRO
E/IWtgvXlhP4CCiVPc+Uo7cNF9NDzWFT1rJZU3iT3WOIr3AT/jf6uAWtGj7V4kNv
nqY0NuP7Oc3wDDyKUq/CDFSx/oUD07WRWXVhi4IemNNhbUGv0MOts0BBoWygJKnP
+/cYXBAY/In3zJIOTh5sq5o26OMc35NYnHZWOgkI+ve8B1sK5Gg7YaHNtei11+th
OWmodd8zyZP6HQcie5U7hHVwyNQH9EXU4az34XKVtAXdtPBDOKV9AqnGFtsOrs5b
E66FKVSmf2Nyg440q86iC8PyNtOXqtJu9/fYthmFbdih2PSxlkV1xtUkF9FiJGzX
41ThAq7odwvONhnigvqwwlH2BEij1GL6B5Of10ljpsIeRzpriIGQvO7WJROWhUnK
WGylG2xi5ww3VMomAx/FhvecE3oGFGEL8bUgnpemFzXWr97zPHFxo7nfhCUsiXVx
8RrtoHEOTZQQVpZ8ZhYPuj3qE08PqmO5I7i5BkGzgCFDPDq1YOyZxVqScfxFKxYW
jtsulhGUbMnTBOBByBCGLwYr2cLOgRqlI3AjoWFSbryL3arUkETXPvwCCox5KoJh
A4f+p/o3m1fu5u+zHhz4nLCPR/YqCfciRShBcAqqbIlIJoDM0tAAuhBF5xQpOSx7
NUneRjhfBxE/Uyhjy3kdPAlL9S/BqCf+jve6jii/kPDny81LX+4l5Db70i/Rvoup
tGIIffSfTqovcACpmgPGVtH8YsKtv4uF6Nt2Xcriq3PsK7AFNxgVavAGCM6m0obZ
uZyIl2rbyh5bV83ETyKdmftG3S3wAoHaRZ6eIYejuFcj8js6vouWhgSKIUWmXn/j
0Pr9m/AeSCgesn61XLqDtZoOnxKKZP90jPKjYU13kfM3z5snfJ6gBD6OCTgdMDfB
jurXX0gWsUFII8TFt4wpQmubt8cNveoXW+f/g1rpz3Vm4+U/8Eypm0vOmCYczudS
H41tahDt4qa8kFTrSmbeJxyW+oZ7bXxyfZ+Ti+zDLOct5aOSGbUmO+ps1lZhCgDE
a0ee9ARiejiE1lNzJlwCom7u0TljqBz/ak9lexeVYUbmYAnYtHzEBbj8RY4X97aw
nzw7uRhmDFxiUQ3tac99ixUKI4G/5GyPszXiF3zUqPxgSJ0FChV5MwUDrJl7VuJU
h1LQVwv8FmSuV2Jh5XFs6vL7apGUZrUw0zEDx17c/lygJFIITYmE0rOSJ/D2cfLR
ps8mkxYBQc67Rb4Bh2acbuFiMcQs9Ep5xAXx4VO+jSA/AiDJ1xpLR4wcGt2+cinS
yZBgueBKAx3IZkQX4Q/1ShRWWHM+GVDAArml0edw+DYvMipnWIRWIfrOBZECTDRf
rOdzPrhEkXC4ZFBhBAXESig5VZCB7stymv6CDQ8R/uWrOl9KrsFjbb9ucQg/ygfh
aV1dTa2PRvvD7WdOPj5ozlIPoEpc8Rpd78JhCpJ2DPZGoc6XAyh+1yH0bEBHEE8V
5Fv9NUr0qXyYLKJJcua4PASS4tDdK/t5b5VQb6BMCrTnTJS5aQTRfr3fZjLbFVpu
lOew7Gm6AwMm0grWNoHJik53AG3K7A5hUYEeqTXM2YM++1zfn06SDcjbrde0yjqd
/82WKnstmgFmkZaanEzjLhEpbcS4jpG29t8T6u7ZfloQB7MANIWcaax7kuuSv4f+
UMMa6c3/QlNPGGrW2XBUEgqXEaTRfp79eWT8wyoIer4CHM2sbxlTB8I1zonRWli8
6pTj4eMkX3jdM6MOWFNO4D+nwi17qryFGwhZ0F+cwOcYd47fzoroXhWXUBx+wZ9l
muuiJ9DeKzVZHayeFkzUJs2X+oflp8ULO037MzLnRSTf9GDb0C8h2wGUT9vgnQmC
I/r1LcztzGvYSoirDI9CaMzxieLKVCtiZdCsloamH34gNgUTnjMMWkwN70ZWmlbf
EFaOvHLfeLYy6Qb/6HPYxbUs/I/EUQ7R40EAS7/py4zJfhS1OHiIrXemcSz3BMp/
l0pmvqRgk9wmtNEeqlnVvnxFXmCFTQaHZXZ+c1DgLuzHXS6CLKHKH1N+9yDjDPMy
x3Z8lS7rfmO2XScBml/pjCq2qqbqyQ9jNyLvGl2TYXG3+s0oxXc7n7fIFrEnpL/2
hnGnTg0lcxjyyeiYSG2D0CMwFHX/6x0H6nBkqo7fVzD6Vg/Uj1q6g7CsNTircLZ3
36HAVp97r0WtcunnoSU1odONlNP0lgAiTt2VKEvZb47UK5emyR/tSF6spuNRTJZQ
oeag4kr47poLD2Nk9UnMRS0O6bXKyH/bsaChhfq7wNo/gbvw0zUoG1FuSwJz10ZS
f9eB/yzPzrFFLJUSH8I8nLuuBG9dd6JGIJZgGtaEzUw26KN4lFF3J7L/o/QCHEDS
9QsZeG0cGq+rhMmwSs8PhQA05xS+Po6bkM/Crme+/yKrIEFo7fG6MqwxoYIluRnR
H6VZsOja11sfDYIlw3Ktz2Fe3W+ULULaTVgLBygKcsx16Jg+R2w84lw6BADjsoy0
UiIHcQuho3BdEb2WVGirusJ8KNWTrABt524HuHW0yFVltRWf3Y0KVsHQv5jKkcjF
c6Ukrp34lOeGH73iyIKjz1eIFodAUpukBlmZ8e0VpQeC+bGQLwnNO0GRMhnIFGLB
feXWq6qWeeJ/RQSCPMg+LYvdX1GmpZei/qD/AK9aXM84f4mUV68Z3DRI9b8fIcm+
b+dqW+gufKTNnug78eWCho/gk2Qcu3fXteiSfQZjolQFp/VVPxMW7iSpQo28OTgG
opk5e8zpp5GdN59YsmNxeUnuB/kK1w/L5c/ORcLYmK35nVxXD8zngHg8ICYPRb4f
RY/eE7J4k+R9ZwszsdzZ93dbuZqNZGXxN9bZqz18dOgmxoGUvMDv0Zu/6FZfVAPN
m1bz2fx+idsJRjtKGtBfsL/QDCYqsB69pi+GdAyJJBe9wZ6e5JL3w4zScKO4fOgz
gPuT2ze5IvXkG5z2SOXc4Z6r86QF01klYcSBUuKdIcQLMQkpGrSUAn28/KbG/egb
ZVCt3a7RPHEMDg9/dbQxaBPk2mQbQ4k6fvySJzfsVhLtTlt/KTLSaupZHRD9mVuQ
+Zp8H7e3yYooiJ/VuVNk5ApMZ2TVHQHgpwZp8N+gSGxlaXwHSTbJfj2VvjlDZcf0
XaJiTa2jQyjqSEIM4dieYuOM+4njBo86+1r1ukndoQe9fr7NC+SdEct0MZR/QydW
Tqk2n3p1WuBl2FlLp6fRxXskrgO3yCRqnDPJZVJeuYJYPS6woAZ18xVQuu7wEA0c
bVIFbdoIqWxkwonyEmMM1HjHtz07rXWp9BzlkXGbyahnZiHfgS0f44auVCk6DuLB
HX3qJlOLHJ07ZWK48EObQ0/zNbXkLKS0tno1FY/FND+Idn1h3dI5e+Hvk/26NiNz
X7hHWirZGs0k8M0F/tJtFhPq2ark3Api1E8CO7PZ5jNgdm2khMTZicjvC8I9G7kQ
fcDV34Mxrlb1pP13eE9TXjr+Q2awFrb/V+mfDs31f8JloM9ZSJEbCGMJs4esu1OI
LizIAzAkjsCLLHEXY/bMQT6T7/heD9AkJg2dQFlCxfrwP4RCG8OtNc0L3roLbRNo
6S8S5A/eq0qFSySUyCyyeAX1O48JlGOHLJk1TsF7nV18gBgC1mmRGImHbNbj50T1
TV8ABfTggis3JAsNrwucJXHCgHUQ4R/m/HqocwmPUUQetIB2VYDI2/2x0MkUI6Wg
oe1desnh6gJ0ry7zKgsfpQxwU1tUlhMHdq1P547r0TAPUH/0sEAXLLzPejmogtuG
ecJRGopj8VcCgoYmcYF4wAcidy3B/HQbhMOJzyiBO1ntJGTHAO2uxdrnU9Wa08Xk
RYI7O0d3QhWricmf0qnpzCGb20MBG7RlOn90oXt23CMXnD7af2o1/ss+TlwabCRr
GupTduWGgvQPn0JZwzPc1gjBgN5LXHTssFyyEPxCFOjkTNmDBKtMXuEVSURWgAcD
rYlUgMtN2/rRA0h7BoOsejcYU8xOk2H5rHFOSF/wZHDfxkZdClaKAvvTwgDn6mnn
IOGxss4ogBi2SnA/W7TtHuy0sazbGHczsZFOmlNtpBb8f5ecqOJWa1bPPnzS+5LT
oyHCQpDz5w50Slsw8rYuttKDHS67ansGYIZSxmqDYk7rQz6rywQZq9qn5GveiYsd
DXdaUf9weljwHSQK4PZ9wOKcNGHxODzZF1WGm827ZppcO8B3HvkMUIfSUc3EFKZs
M9S5YQokgD4g49AaxjGS3XXmuZGV8L1hP2gOTCCXUcSqLv5VqjWDeTIRcidJKX8u
OiVzOBW+K7TXJ+II75rS7Sb+wwqCCG7QrzjUjUIBYrVqK5A1g46HrEGlbN9JOSEC
cSqMLzIeXmZ8244qvZPUC14X1MAYXJcVZUw3C+gngYc6Ozh3VmX87t59QJG4cxIc
9EmesVU9PMr3EOwTQonfueVt555LCs1L3TbBRZyywXjRzmxNQrRrmd3VPR7ArCqF
mm6urAUl5l7tdrZ1+BavmQKOAdk0PuM+/ws6ymyeBFsMuXI33Uyeg/c6Ks+7pqYt
zofuSXsPAYKFih2d1JPeyr2fOF3RiGTNcuzwaTULuGO/TobX+CLsMg8YVBrbfQiV
ii8uZsAU/vdH9dBV5IXIR70r6EyEcSS1LAmGyD1q3C1E+R4zIOHxoxZGbk2MTLRv
kkVsr/QgtYPkVAqW2YrDpGALvnMAuRELV4U3U6B9DhHjTvzSTR4z30p7GgYP3RVV
r1MUnszJAaJfooiz5es0ZswdI+Q+age+nCzbN9i43AjBLNts1Fz78zEadN/pFEUQ
pUvScubNDzOM5ZqQxOOKWPGix20VWecMcT1bEDJWW+wEp10Qo4oyvHGLr8GQWjIv
pcyBPGoZPmKUUmQ0DM0O7h0D1Ec4DdXP7ul535USuEGVHKjUjOtoe1BKdwbqjeOb
7aG7lowdJbVE52YUqZuLmfqyfylPLOhtczdk27qZcJ2kHHD3N7Ix5QFRQG0lkc3T
P0Pxbfpi8vmPSUASXCwFBqi5/5zMDR9xcBTM5fmWRpG4iN5nzW70xXq+P5M05ywa
hrirZg+egbusBJKBIV3okolRyn8os26zJ8YH4aP5gpM8EbeqtQUznmfhlOoIv9zI
NQQfpejtiNA/0I/hLQQ7mukxNL6wUuWzse6wX/SJEHFGWKE2V/ICActVFdLWNT6U
h/Yz7ZSCpW9zdST5vu6AEPL5qnzGlVVdsrC2JYSO/jw/v7SCDKhhmoavU3qw22sL
5T+d7PP8hmD7ppSrmG5ffiJdA17UVqpNw0/fQ/J4mz4cy7Mw7n2oCtkLyqi4Wi5I
MstGMfIjHXOLeb6xz7juRbYwZlLnjumenpOX5slswVlHbQ7mAVZ9CQAwvVPo3PxB
3aSDHDurETf8e14078W9AqzHXLUh5ZuDNwlKo+rIB9AQdLJL8K8i7HuIr48WN/4B
n7domFnFYWMkSFhjSdl8JphDBiiy4K5WhmFzn0+gOsI83AukkIAgaSgZ+JCzNVLi
fpXur2KdnZkdCOAvLyyrxMsxOXvXJ4rlLa3yUhVsfjYJqPqxXoFLc9UvAQBJBauL
OEchfxfPRdVSbFfIDW/BT1EQfwXcbd45f16OXlPYh3uOvQuJEjOOkSimGgevZu9g
eQRg43fSFMJ+nlW+hbFadG8J3pj1Wap6vN4D71wc2AstkdopYt0wdq4CgN8qcm3Q
Woe7keqVN099HTC4f6i4CGh2xliltGr5ztl/EUyksq/eFEuPhEdclboRVak+Ft+M
NnK3HTnIh6wKb98Q2iVhy/3VkeZQhO+7dedOJWiEOlO7ITpmI6FVyyYCHLfBR6ZV
XsQiP8TM4FpIpKYqY4DWlCAMtlkE0VkEDt+99PJ9N3sz1dVhUB+W2620axdFH4KW
fm/vXPZRXofm6MSemkJCOQgR7sUTcm6ygBEOYcNZq9cinCYjNjW4z0FyPmaCS9I/
9o/CsVob0/HFt0IV4EvMIBy2KCrgouoZs0ZMnVPcRvIj0eqGiav14qwHkRJHObNJ
dEM8z6dB9rfioCaQtVGjBGXQaveY5jgMe0qMCwbqHmGP1PnA+3v/ifGJMXbVu0d/
VTp/MvOdvAba4IoJzGpEl2M6iSkXGFESbZZSiMTaPocSwQAOMwKLry8+oN8cLIR4
pVO+9fRhNPQU43c9IMe/j/Fk9VpFZCAYwlNIV6DdbWl1HtKoAC+z9UcMfeR+KBR7
BZCS4mpFSji3LTeiai4Rt3bV90bowLyGDKC8CHjdMs/Yc+qyO0MfS1AGR/wUQogS
vKDIQfZgBVzWRU4PBaXj+/0TNR56vwI3NTINcjnVDdjvomJCpbEPLnYimj8wf8mD
NxffPMaJ7HbpP7UstnToNZG+GjCP6m9umABlLCxIXRRYHYm+5iGpoIWcLBvwBH+1
Flkfe/3qXeTgM14IkEfk9fbNj/NQpUKts70jUK/KxJkd1MKFGEFKeOI4mczdg46F
BEULVs4Me7XQgn2WEQ0c56BTEeqkROqc1NClSM0umO2fvbGk3r/6rBqgOIXIEixN
JiSfwV2HzWKOD+q9ZlcygL/Mk/8RJWBn8XQIi2KA1Tw8cC3Z8yxrlWsYOdLipNQi
I395b6v5QNkdH6skNpkWHWXNsTjQoj3fTEh/PN7FXzGN3kvJZqmlPYHrB/hWg+ZE
oaLPaCKgwoJ3w5nABpvriRPIrkMOTtZdYHSE+7jhb1a+hZ1r0AFqizh435LWWBZ+
iMH4wmiVZBFZgZXOfAoWDWOGs7hV8+WuBOIyYq8hWfFy/ynh0MBZ4ywtm5X/KUG7
oSEt7QSahxYEi/PxOusgw7x+d1drAHKXYZ6gcHVfo8x0O1JS4LU/AQCj/4LH73pj
gJBJnxDLmV+HQ6RJd7odKCEmJ8fvcSf3KMK7YiuYfZ0GcUf3Ic1R4Zb/PhZUsMRu
vFkDt0WlQgJyXbw0dEPJmRr32bvAUwGyD4Zbz3guWySgtxQOROBVgx/BhaWPzLYk
svSOUytm+hewXBmSMK1bfxh6vdHwCRuFuRhdlAPgQY6nBStSMMY2ymXh/hPrk+CY
/BZuzHtWSft9IESh6Icorqrh5YrsavqmDySF4b/Fg1P64G55eLHxQPP/vAkcNdr7
/ByQ58I4RAj14iGHjPmxwFVQMFBHEknDWctFCiDOqfo5ER+9PMdYfY6DuvrjPLAJ
1rci77cH2hyfA4NEqAkMh6zDikeGhTJD1gC4Zak6GhpcbSWnVSH/R2b8m7r7n0Jn
Tq+2xTWVoA5lekRBc6cI1xXVEhRvE63n8ON2XKZXIG9bA3BmZXAhHyYhr7+kVPG4
XU3tANYS56RUtP6P2y165w5TE1N1ihVsHeB1gVO8fQ0aNKo1KxXeOB7LivE2RpBt
eVX7F/EhFnOd7ikrJeMyJ0P8wibGmWzseLt52GKBqKrfYhvplP4cSRa5XzpC5CFl
mmvjpFf0hAtqpHPBDimB2br+l5iY9QfJL/iFyd+a+yF7ZgZWhNJf71vO2jlnQMl6
zo/Bwnj7FC+Xxl+CqduaeHunXmxlrqYxBHjQP8UWDFZOyV+8j8fSY7I8iBZlFsIE
kDkUT/raVMQ4MxYGTOrfrgkii+bL4lUmIA9B1e5017Kh7yjV7j9ZxCuiLW4fy9Di
FPgou3XO2BKjiGW9JC+LWPhDdW99UCkwGp2y/UHvIDeuY9ZU8vHyG0Fue/uw4l4O
Ej/Th4ULE+hjrcHZt2KZHq8emq3hgrLOU3vvqxy6whdwB+47MEMWR7EIgI9TJMOn
kTrrpRZOuy4ORc9l7SY9PA1id3V07w1qEQqJ5Jvjkc37Msr5VA3gJ9fldW5RrtXU
ygMRvAYAJTfFCfk3TnFfqEM55fXD7Shy0I64i6p84nn/WH9Iv8EuRvaKKK/ttX5D
N+PjXAJFCoJ0SXoBVRMJ2maHbGRNDJk55VehqmoX8CW8VJJF69soMa51M+H5QsEh
+QsoVg35leFjU7PMR1h/6Gv22R4f5aAbMc2+PPxanX3nO9/jrMzD67w/kMosnebk
l3uDxYBlbpBBfSpMI8cAEatxfiwVTorK9KOqCAb6XTuuEb/qrwzXO0GgLTa1kNlj
XUHIU2w/J8LecPFReQgy1spLnIUTNDCDzoS3Y7/uD6sW9jNT5HXf5/aQ+eKpe8jq
E96ZO8UHu94Voz+5Y1iVQVuU+RnHmnLlxrldyNy/1XAfLvr/1s5uHyS2fEwTO9wT
7hM/KUCyKFN1j8kotfjj2zxAreb8tqyDbrkQPJ/bvizHeV8tUtTdXyLXrC0hDNwt
k2CsdI7Qt8yTZFHJJqrlNJHLtH90jh15uhcdj0P/6huKXDn5fSclgMFbpmEx2cDZ
NkNfjNGrGEsJXs5kT3lohP9loC9At/VYhZ8K9U00EqrRjCixsgMmNHJZzLTJFUf5
uXqBMTZNlKilmdfs8TFtS6/P/FYP8i8HtAllje3BYrsFwsZLtXvIeqyWB01WGoID
kJqVW6qb9O6XwIGSLdxk5WEbHidAvjaJEkuSTuGv60AXsqC+sU0qYX7LHsvSBHAV
OpJXn0DcC0jWA9S+YQbxDPPdLKlciAfbr9AUJUA8KsacmdiGv9FxIVxqmIUsWmgK
fvViRL9bPnEKTRtRkpu/JjTpyfqQxi9IH1qo0nNvyMks6u3qWiqbPoE045XEqk+E
PbSV2WPlYAfihpYoIfnjIPWNkqHygYlKjpPTjv6DbxWvdh95hbqhRqrzRv4ATSW7
hXdvSWLGtpT0I6Ex6bZzrCaIcYFiNxY0JyBEeW9GIBKAAVr8grcGudfJW/cXvu97
FCNBcrbFtyP4zkRU8cvjQOJgqRgQ7CafKEbNzyYkZoIuz/9zP4ETXMyGn1sJ9+ED
VVGezUDYVu1gjJNimuEaN0B2sXt7hFqPsL4NsXxpc1EQxsxDTNPYKSogfu1wsh0r
lC04PmZPX9iyh4gqAenLArmn7ocVuKHDusObNf3f1s+1haXuAsN3aO0DIq8oiQbF
6iOwSdus1LY76rA9um1IPvmoBuVbO7yripXLte1lLpPYc79vukQxBzwD79DfLdbE
UAmUYZyPEYcPBRRAB1a1WLqx0muzZA5N2Ld3+42pPuEjXinRj+nVoisqo5KYj9/g
Phc6zHH7LyyGk0DiVCkCAPrxilxs41FOUzwlsauy7eBXICcbvnj+OwPjlVR5M9/Q
+rGzv1NuaATyqEXk+YJXEdvYUdagSSARTgMYcK1aYG+iZUh8+WHJyPuA/vhvPGBC
3Q0inw3FKaWe9d2N9avrrGyo8ZI0i8Qf47XVlnODGHPmHav/Z+niz5sX+XlwXj6a
lzoOMDQ6VzPmIntapDbYio/I+prCcN2Rytx/GjNhj99eiLuD8kX3SHjmjzEl1XDr
wBULyixZDciFoTsffffZVHecJd2bck2H13EtFCqRFK3by7Q0uDfaLrsG/72bCix1
HyyMPrAepSe6H6vNj3lp5m0hhV7V0itnYMoz005XeLss8FIeAfgCDhwX5Gm1yrHz
fID7oxnhpNZQDz2PFCa3l3wQdE4BgmtJ5r2LSa6zfgqZ8FxmFNumNS3AHK/HUVXh
7wGWG+g1fsbSeEdWsXJ/R6HROpMkwimeh/jdheWOOs+g0WOmzLDl/HHRInjNQ92E
Gfwic28y7l+xi4DMGQwh9A6WlLvuXIgqY4TuInEE+a0jAUFuwTN2ynVgNcwKdH0M
VF8VSLxTsXjmRtipkuzTd/nC5ZXSrZIdPj6y/iuqXHmdMnpXWRFSPV0keDN2BWx2
tkuQDZ4lqJjveuXGChVefAV5uzTn094AZax1VkUk9F+soyUGkbGWevN43ojlPnXI
QZS6jkAxVS28Je5zb8Kd/+qx7BbF24PkfuI0XzeY+CaC56l97NpCgXqBpzRLSbNy
fWcBNPrc1QaihCZUmEdfrKuOb3/uJ94/mSL0wzePVlCd7L0Yfrf1G3xkHuJ5HKQf
G2BYhYGyr+1Ph22yNpij4FDdhsdGJ4kRRJZKcIH1zhupaalnx4CIiPsahIEADhtJ
ZHB3wqKjlJPVmEoYlQyzz91bvx4VQai4C7Kos5FmBq9o2WsAd7x6JEJ4US5Prnn/
XsKZbBbrUfTsda6GfbgWRog3oC0p3uO1GgmWNKFo/E8MH8/UU1MT8Mm96jtyKgzG
IfHEUtM0dCpWph/Wz/WpKS/BYhh+P5CA6KDruzh5gWjCljn0giv1IWT74iOcy2Zo
pHEZa5fpIPdGF6gJ1dp7A3Nd4J1s13xqqceY78Vy0iZNpD6GGOf0IIP574RAmDdZ
xskZZrLTJVcY2XM5rE6AfepXmsjSa4tyOtTHnXUoV+Vv9kGJW4OWVrIa1EWVsV5N
EP2uWPpT7FoL02T6uJavTB2ZDbpmCiQyvaYmjW7eXPDEmePwWaA9/kV2tN8h/4I/
2tf7X3SCkcnSHt0S9r/WLzSDILaeRi1Zy0JvGhIQ8j7sDzpkBjImGCZ+U6sLNoXZ
QVyP741ga7OjNx1HbMNfj2TpueX4xEzXpXdHiTH8IScjrAPTJVhycaVI9rqYbJlr
ArCGfz1UMD4UH/ANkmAgTw0phnwJr9Irb9R8yGLGXeQ+p8KOBNCpQgavELFdaIrb
ei4w0dMJOoh1k5LzmY2eGbqW+bPW/HOsADYqTRexG16HuxBhJI28XMyGQzaUFfi+
e3+PT5+emoCPbjxlJ5d2fzv8TrfE2L4srgcBuDgdcCgqlXoqzBYfqBR3rqEo6rET
0r9cyho8atMszlUAUzWe8O80easS0DBFkSFWpqmMurlRGCJNVcqZjT3RQ5ivXMiJ
BT67zvs/XnJlhj54sL2cwh7fiGi9YTQ+p03iGu+gqA/LLykMDBiD1H1zTh/GuZbK
QZyKIzsB+lg5wy652gIGTHFK4Efu9SU/GmW7S/PeLGqk+YAfmX0COAayowAvGhsQ
BWAHJ/7bTLKtEzdhNPLjjP1q2cKIEN2ogSkth3783marenwr11bXNjm9Q30LoJqf
3v1rFSNqphaKs/uwjBj1hEDpwiaJbT/cO5hminy+0wt57f+eWgScAJKVlwZjfbdN
WOuGQM7UuWdDuqZ/8dPR6S8yGFEhdU1Oyk/9l/t98tcHGPgDvbnCeIOU48pyIqc8
be4/H0bzTO33cdUkF2IMfA5+RQJMMn+Hc6ILCZJqKPpPEFSn0tJ2LorOrUmATxd3
lPkucrAQcuQ5TXZepRQnU+fIYiMjBAxgldiTkp/5QXcFPY0TTkzHCuOTjdXc42/r
4+s4DnwE8+KYG9eNK5zbfZCo5IdHijhGgu+hMmVt7Lw/vxh0IwT72X9oKve1fH8r
L+PIUJ17KGFUEkWT4HBrOg0eBkKJ35RFcd5uW+uZByzOUO8Zn3C2Ry0YNs6e9FRR
lZcUGgIOnf+aHT21L/O7EzHV+nIfNHsPjIp0x8qG3Z5x02BT8LezamowT4pXju65
6Kf49UZS2r4gHWRtzh+q82at8V2IvJzEbK1dlxV//IZRotGjaHDDcJw9SWGbu9By
OnElZ/uJFrAOjuS0nogWYx0bkHjr/XNy8JL5WNYPU0TnklP+KYUana5zCX7lFUbn
bWe8SEM0WgByYBZbNDuNpUqz3Z4oTYlwdjdCSnUl55tfCPWsRaK3Lnuo5j9Vuemo
6IMaWCbTQgS1GGZeyziJxNDvMihMpU2OSJYb6xz3K7Y6g7OxZXHh7dH+FhzV+GFw
v7oIU0ZE6CATNPY19EWOPp6yDIRgAAoCTaprjl+Chuyo7dPoHuVhuLpt15AjF6kc
Fkw0AWu1xVGPp66vZXY1k9ijnLkL+kyNLk505yOtBUFWvwYifntJe1Sq34GrEdgI
QD7KJcyjB1smkhO5yKIo4jpxPOmezMW98/RvrP+HonSVG5cl8oxt6LRuFIiPokKW
gTg3SJZSp/4PnxeoBaSFSkVX67dxAy6JXUrqYTbN4dmOA5wSzudticSaObFM+jm1
pWeYGdb+++2I9dj5SFkGASNtXxaHpwi9PIrcgSfCsbuiDbimMtK9ltVmhCJ712R1
lo18fGv4p84iAZGvXal37ehCe0nzlyxtL+Xa2Tf1WYlMcZRb8RzjMxAs8RMvhbMi
sweCeYeZ6P2JCbhx2utaAMCz3QDRKjPykyc7YFt2XcPg3jlIDQMscHHMZhMwD3/X
aD4x6ilZUFNgsbFJEDdnuCLvD3oS4NmWcB5IJE5GWGFHwZNbnQdz9DV4fm28qx6B
MOqzff+/uyX0LRdTqdbmlXow1Z/SRV7+5Go0ky3rYXK1rx/tAstfTHAxqzuSWorN
K4EN5zVVoSmqRabdtPpybDhKoIdcMSkT+I6UfW26zxiAwgL//uJGM5S/UehO/YoD
7VQir0VqVJe+v72TbWy+qy/P4egXg67WtMoPyt141GrWpba9Myx88WoYDW5+wtQf
7XtGITAlCr4ncS2Xp0o0whWm/LmwYIQYCOfuDo8y5OZsmJQRs4+aYmp5uBeVCz5G
biGhEQQwt0FO8Ewq9/n0pogwD9GMrTzlq3IIezqEKLFXHtmrs0cK7Wmxjusr+SB+
981P0cJ1hfeKbZULxEhMbUt0Wm2XRXWJGg5qtQc0sJvfQ+G3dnNTL349YCWJVyzL
ZgKMyDKupxIFoOxGB/sSXQ1md9/bGiJ5FE5TMyFiq/GpoewkYDXOh0XxbVWFVaQp
OrC2nATHLFEPFiDh9FIcFKF8VvQdCatLGKlkDShEDOVgW2W3qaKclT1bxBbKxPnh
+KeCrnDWcWzK9A0eQa+RFh5d8Ga3OY4B1wBmr87Iafx1KRcJllrxxNEv6Bo/Ox3L
7tIwRmdOic7mrByb33evFkUExffxdIfhlOyevTrUqsWMo6l5AwI4v/ef3Rkr3IfW
CQ7UQoz4XXUxOvLvLdYWXfRy+NIs9t5ewdGcrmZsVJFYO0iL/3ps2z8UwxszX0+l
MmikVeMwiwwaVerb3zoe8ZiArjH9VzgNsIcwQdsBvJNWk87RibgRX5WycL7v53J0
fTCFcgmrKkP2QS//olcDCDW9bNYuG7OD0iUSC18mDM8LgkLwODbRpVXXN0sy/q6J
gEV0gcXmKeYWuCKvC2h6FWf6Bx0XWcoEt9tuEEArSMK52B/yVKMiQlbIhjWYC/ww
Z1+iuPbaVS68blUGdygDjdRphhsvpTmo3+v3LH1KF93tQNK0wdU0B20tckEl3m1n
/ZLoTS2mbHqSwLcgXyHThC1EUl4xADf7JW/QR3K4vFJ7Ciz/OL7sZ9ex54o2/sgP
bmeBZVmNPXxU5Rh4LJkp8zvqjJ3IM9Kz3ZAicu/136tkJPXZ/IlG6o01FJxwCmhe
sLBPsUyowu3pw8ZCjnMZguTMuE9ldEo/Zu28srfs4T7t6pvuaSKsXeJMJn63MfRa
CqXw4pTWmYCdVe4su8RyTlFqycCarNVbH1leGGjbTHYxNBpzIVYspWNUmkgRGFxH
uZCICCo/ureSIKMUTnYz9b7sqKFqiqJpWFqux7d9HcpuClPS+gPuS6kyi0X+PI4Z
zwNoVsmJ9JouXSr/AMFS94i2JEP7nMnWGfpu2hBue5h23LFLlXitD1n06KKrFR0G
1ylhtmeYZpMQb9DEo0B61vJc3L/FCctfl52SuVP4/C7j214032iKH+M+QgCrD5lG
6RwCiyHdHvPAUuM2v2ChyRuZhNKRh+8roiPBciXCgvK76diaja3qLyDQ8/IRBpZM
CgE1jY2qPdrALpOM71UTVHKjkPG5dMA9B0sMr0pfqgsGXBIj72Ab4r5djW6fDy7Y
K+3FTagegSOq8FNFCWPwZH56+lvq0esJqL2sfkVl9JbdAJjBHopWzUEiKocEwB+F
AlwX2FicVnXd3eVuQ6mlxJND77d+tsZmi2A54fGxYqw/KZnq9zGgwPEJQN84gk8f
eZSD1D940l8gRaAP0LdeJzv0DWQWvtZ8VFoESzbyLu/DHwZnbVTlma6R4qaaV7+n
20Lqaifq2MrGrJnpzcr9DIZSW0gTWE4mjp3Pp7IXLIQ+RW7KnBISvlRwuxe06znp
jI4gFWwg+68UrwIPL+0I0ltcEzvob0cm2lyhETN0hzf7malAqcg0F9wfANB88ZnH
06JXS6qtJfOdMSEJVn0b5lBoknjI9V+zSqVNWh1iy5kMS+ZPLlmgHTlrZtkr/vqN
sWARMsQEGv2ohP5YRKjW1R4a6y8snVAxmtjtNFEiDveZePKsMq5tq7UewrYVxOHc
rPdcM2RxeOfZx4qyI7kN/CpP1kqWwThkJKOz+L+3WB+sUv0t8zAltIMVhF5fhLys
7hueeq+rYXSw2Uo0erF6Dn0aJYyplRC1XKwwOM6VMrSjp2f03YfonBVTTSc9EQn7
BM2OpsZrvghmruzndc6i1jFqpsqxWMZ4w62VlaiM2R65+kObGTH4WOEkRs5fuo84
6bAq5rXXWAedka0uzJXl8W/jGafuHaaW/bJOjAIzv+B0ImEyFH9SeFuYzHy4EysO
U8csCGuQg16o9m9rBN72DjfLMhs9SzbnSLtaITN8Veb66+v26VlP+VLQ9/ncqKL2
/mhj/BANWlD9uVtAftErvGHFUbOOcHAhBPUOn8JrAhDDxl660Xq5e3DrMWE9QW8t
6670Iwmy0b4t1xRaa54CAmFIAt+9Q5KjdbUQ28kVZ8+huAVm8QvuSJo8Vzocg21P
sobhf0c5AJn+PJ5GvSiYLxf4aNvBUb1V0ShyNkEB+cEIuSUPShmHyNuMUdJZ1wSw
iG2pTPTac8uiqgUC9GlTKoi5SW6gPwwiM41fg5dBfFQwe1hI6We6TZRGIyXLt3o2
yLMKXr/acmM8VdFPpCETGVHcl5BDgOVgZZTK5Yq9geYg7F4F9yk6X1MNWbF8fhfW
b3+nYssN0aZjR8x+8+RytvPFJ7eV6b3lD9kgGT8lI/bQXkZVy0ZECT1myv0Ce+hN
847HFTW5sfnQCLAlbS5R6rdr5/KmFIQK8GVyp0iYY1QAKaTx90Mk+0M9LSh4pI6v
OUab9KQipJydF4stJgeuvg==
`protect END_PROTECTED
