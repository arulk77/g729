`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB5TWVRBQk8uq0Ca+Q8vGe8DloC/2Z3GC0xLucS3nL92
xqkXkXn0JPevRs3f0S8LOVspIyxLyreUGwpUkcObL0l382/yq1NxMD1qFFF173J/
gzLsecK9ZT1hGwdaZ6Ho+okLQPHriD9J9Rp6f+Tn11Ke2k1mj/8YfTOR4IM1gbz1
MHKtpCfxgRp5uWEv4N5q0g==
`protect END_PROTECTED
