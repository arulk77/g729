`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAbFyGmSlQ8aO1nx/QKxb8hSv9eWNKS49/GPLofJV/io
26AJxvRZEuIMrRAiKvi83cL1GMsJm5kWoR/9a18F5JzuitwA0X7WEvH9r6383sJa
5TIWDfpz9TUv3GzAW8eaXSPayRTpSOcqWF3J+ArlH47PphyBJQN+P4+hPpRFZRYR
CkM/S17f26yrcGgUq864U3W6NHqUq6CCNX+NK+SnByZATB+S5gv2gl+nLBs+A0A7
elq3l8SpoRciEmjxgIt1t1IwvfY/UIpIblTIoZM3QYfDXcEZ3lwqw5Hyu+UFO33s
Cxz0T1PDspLm5b1LHIXk84wjncNpf32TRA0Qj0hizEgVDuZafnD2BCgx3qy2fpsq
25NKFrvaz4KWIa/C91ImJwAgf4Tze11rJgepSsgEAMI8sTuMr7JBRt2q2UmzhyP/
`protect END_PROTECTED
