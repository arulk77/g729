`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN2ggRoNELVRRtOtMGnP9WSojidnELr/T4ouH3ZiMfGzv
yuqHO4zTbMhOsg2ulS+Qstv+2Aa7/O/U9GitzODdr4Ob9rLxGz8Xm2f9FNdIFg84
WW4/tH0Wdh/AuBsxrVd92wHJKEZrtKABEhZzl4oAsRP7d+93fc/CSYaHjYExxgvp
MNRz7BjFSivkA58216TtKd+WhWzaRzoQ+4qexBkwxuRjwcGkXot9HgQwq4HEHemT
+jFIX937lKbRKdw27SBZx79PvA5FVMoU5NLy1BKrgQDS+nA2sYTLjRYPssRH/Oda
LlEtQWEU0C9hks+B1vxIv4eOgevewasSsOELDRRvXR+wj4+3DJbIUF01N9S/pupQ
8SiTSr/OueaxHr4cg9/FFlMLPRQ8t0Utoz9HkTrX7E6T/vxugqg1Lq0k3vzCGZPT
biWBC/jPHtJoYyUws8xO6ZgqoPf0jy2mWOwER8WArFtf6WC/dKBFei69tFQexgzQ
oS725JHEAcWv1CYg2zPvjgvuP9m09FIJ4GqAraT6IDiZ6ix6tv+QyZdMdFMX8fni
N/kSb3NGKn71XV+aH2BzG9Da5UJBFzf/oaNrU/iNCMf8+lY5SWP6rIVK2K/uunWQ
Vy6bYJYcriy2osf9m5nSWVif0JCcDFJOg4cH1y6IDamDzl6ZhyjjhEZwN2/2aPsZ
j8X39ZGhCDFnzhCyUKhSWxX/UxwTA6RciOSOEwbLqpLylN4vAO616JsdIBgnXbWi
sE0E2tZ9gZXlNQSXz3Hn5RspMXw5IeEnMON3FgHjgqvzJ9gz9pY3yeq03J3wssNr
Mxiy/Dk+bLNoYMHSrAyXHgbP6cPmvP9hJm5wJMh/kAh1gk9GmTImk49c4wbPtlT8
ua0noG9qShLOGEFNTUATo1qotRostOZdXCSVainEDE8BL7lGpGuDDFMtL7HdKkj9
tur5Ussr5OeRlqXn8wOV/P9zp2VBS2LD7Wh9NaDOZMJdg9fbxtPdJvsy7Co7iY7P
JCmt32gU66P0IB3laR444YB7hp6iO70Ga2veBUkwuNvnxKcOsesEMBNRV+QvrjBU
0BFChikAm/rbi/O7T5cQUgxpVY13LJPCR3ck4n8M4OcKJ+GCBhT7L6JcAyrjaiRh
nLUmPGGSBZ0HAvunAPt8DNskBhtRZxSJg4/vNnwVgfv24Mz73zrhjpVOsicxQZ2Q
IP9S8nIYf+NCsLcUzDWFwIdqY2l2IDYBiOChcFyB7g23FIXsV+ND4vwwrG64QMym
FnTjqZhQZzo6JDSaVom4lacdgokN3P3mSzMWcHmvNNWGSrwuFHnbtvKaEAeZALJn
J+LjBOm8a0wSsfOEZ6n3/ms3GZ9W1EzzKuOiz4Yf5T3whakjDOcB3S0Iz+JaJx9w
XIs96UVu25HBanV5j43gHKkmZXK04OBezqWtLMGfgPeIqm7LfraorewANmqGGDVP
3HGI9TFxJViskbXug942NiL3dQXXodlpnQK21T3+padQY7z2PZG4k1eWOzEUcuQj
BV1fld+H5ZnZkegRRiYSCbUTlO3b5jx0KF7iGTKjtppnLqJiPxNzTlFXWtY50igq
OQAKoojtQY9COs7v4jn5ObRwwFzrcOMSBVRQcbrmwmusTX3cwsI9IN2648sWiSpL
ZpJTdTVwyapdecBMuoBHfPKIo9SmFsyonWAX2NWSOYUZSE047dJLi9ww3nWTBKtA
1ruDe9BOfuxvvj8OIgIVFFpTS+YAToWBAzh2VmMhImOQZiPIPDvVFDBFDxWMjyea
qAP3dR8Dxnox+2cdGOYqV27rDK2p5Ffmj1n95VXAcUKOqR/yJtJYJ9gFfy69gFWi
T3UdsPCSDayqPuI/5rbDOgvj2flpHUIvNA5+hRAM7pU7YqAandqKSwvvtufjTEa/
cJ5tzlwe08FB3OY+pmspxfHmDuFSEkobZ29NJLKaENnlSF72Nv49x1Zkm3ukhqjs
ZrozM/BJWe/UStIfXtyFEJQCf+RpgtcAhqCQOKE4KC6f4UjEPf4+sjPN9ukykHoB
OqFR75VNgMW6xbTeOzPxkL4XDIQnf93J1kqNnp7xpV8J/leiG5HfqXcerFWL9Tlt
Bgoox0j8e77U043FDBkanY3/MdeyOfeeRkQhyZbBGlrKz2IsiWA7vEy3FjjYY8h4
rZ38cq/sC5vWbjh7yukV+/4Dj76o9MCZvgRpOAvhWO/CpieGxfQc9WikamVlnwU3
zi0+zsVfctR8gO7MQD2XUipmU67lwJLLN5J/A92wkMOg1XiXV2bmgPoc5y9HdR0U
3Ga8QJXZXnAnC93vaxUeRQcfW1WwoSgso5hSDiNW/EG/SOym03IRnu5iV0v9ulYu
SXXjxuL+ycxfEgw+KOXe1y203KR92Dp6VYJ9yACveGMCt5TcJ3t3K92Fdld1KIm9
PfLx6fiZe43YvquW461GwSAD/L2YHiYQsfzx9n7NLLkziYYhpWsYdsY6ExtPo6XE
LputWHkq1kvQjreM1svJqIqFYRFNsy5J0pHgWBUf/8QqViJJWLpDeUPzY2czVEDu
sLtk0E9B5fDun4JW+x8tGLh4kO6cRrUyB5SfSl0gVY7uXm/kChbtmObRAkhvyPKE
I+1vvgie6sExDAnhAaAqcfaoNKf8X6teTQ/aKgbdoKp/DMtnI88gYsTjeTKPSFdk
chHI1FUbT3gLm6S0E/5jRYDV0bo7FwH4LOftkDZZHYGjLZn//bpvcU8UOZYs2MOr
s1a4bOoaLA5PAzLgrj3/lLpOf5lSV3HrdGdAEg0fjc3Z2IjB9DpwG0wJOLKh7pOh
7NGpWR3QdkYsC3rt1cm25lnsbP0rHpgkwZ5eWrtURHTXkniZcX52P/M/GS1qP1gM
unbxoQm4UYyozvCjdlpmalWPGxmiHV8ev49+v7WAqwOqM98Ykm8a2A1lAJ8D/mwO
nEpJJ6bwp+e6D+UoAlA+Q4twLtzxymMDd2k0feZC/4WetsgjFxEV+g2OysMitEq4
NGXNsEgzmK5heEpgk2idScxpIjcoZiEQw9elVAPj3L+Fh8tCDJjDamRZF05Mf7jk
cUsv+ytSxbHQvuQMaB1gjcMef2rPzxJxyx4/ozRn1IT2Kjh29MUZs/VtSdAbIyoa
89rMQB30YnUrYilIgf3cfuytc0w6FApouMonE4CgkSSPIMNo4oOLrjSeMtXEL3Re
iwjv8a26rWJOgXT770qLcCn6LNqiuIw8HqdPohaWcQke+ZvWrbWzE6LAVKJW8zoK
/kfZub9kryDJLJP0L9BklWq9nuiOxhM38ygFkl9z1wrcrN4GUfMv86DScdLdwW/j
6MKnJbVt4Gfu77o9/o3JbYxJ7Ck/ye3lHTej6Xej4Dm63H1SsNDDEXUCz5Ytc+eC
DYkaeyAi/MGBHkc55rjx34gf1X4cJYK0KhxzoL+f7wtR+iJDrHDfbWweE+P0H7CK
KUXMmiYpedEEwIAlR7VJxifgo2/uGNfiCcVC9GB0otgR5MuOvnY9DJlJc4CTMhuP
WaxfsTUSdFiHVo5FhSC6mTyLK7xgWeF4AUSxZC6ZqHc+knLNAzfDOfJVcUDLZZKo
+INnV9KRgoufp/txaRnUOpZ/Kgou6Rnwn5JI2FOT/oG7GQOnmFm7qu/PHMGnAXl7
qwd+EI7JXsAIx76gNDKv2TMpaqXPU60NqheVtmZSKRcnoozx4sjKG6s5du8wcNRW
Baz8J3CL6gfHcZky/pbXHOkqkcu4L+idCfIVBJTZ9WGpODufEcYYFKuO00TOJf3C
WQhsrKG5o/lYZ/0usd1eqyQMH624m58GsXbJmc03+u1EGPE88h/+/Z00E2lCwwLL
5SQ/riJ+TTIm6nXsWJqC3vMQABPlz3LwK/zSbBoMV5825ARuTq+7eKO67wJvvpxe
6tNZk/EP8bfTvAbreU1rm1LL6c6c/70Es2s/RpjyxjM/BHRa2xpSGYRSH4vui9yF
Dkv+btWhYHpmmeqK0Fhe2ybE7aVgvXOgifJEuAkfmboz0GxdlCWIX7xVxL1Gvj3u
ffjQJ28wpwaCZstxLuw3DiyxWF0oLjQBx1XZzGjRy3+C8IWkJUaBxoiU/ncwhj1O
J98UAB7wJZkT0n/Y3jrz/UI4siCvlFy3CRWjCoDnUk54xnvWokxx3+YjjP1xFDJd
VwWHWVzAzgB/PaVBNkCI/KuXmKkxfSnKqXwZ9wDJ1NDMj+t614YP0WYRVDZA0+yT
mGwyR62P5UhEIPhZZ72cKXXAbd9ju5276CDHp8BNv8cjXxeNQbaBsu89WfspMH0N
6NTF850Ti3M7NdeWew+Q23/OZ+JA86Xey4kRIlPi5q4AuZ+NGkvH5Ed8LIsj3qOD
ZCM3Tajal4ajPsUeuuSiU0VPxiMeSXIl145Wg7qfBnNZ2o9JRa6iAnSjV7wW2Owl
52XMSOkA8oDirFKi/gBD2Q==
`protect END_PROTECTED
