`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveC8jPTYZDgXz+kvL3VGn2EK7ERAnk6Gzc8IafuVwP2YK
QWaY7rKAnm4YR6f/W8ctlWhQOMSabnALR/3kdyoewpPE+kmNHgtsscv51noM8yfI
uXqxe+WnchBhMchOE/yaBwxPyI7yd9NQUtPyirTXxM6KbrZ85DsFI4NeBgLnZnBP
fgevOuWwbKLYV579soV+ekDMkzHhNEXG47aXlJbS5jevoU3GRcWKdVLwdWGHPX8+
qAxsbGZCTu9ygWoWZTv/4DVSJEFQSHi0lC4PwrvcEY4suEJbvGXSha1PUpdP6Qru
+wki1TKWtrLj8/wloGCn3hSt+J0asMCW51miiy8BEQq5ZT0WD8pB+PvE6JoWu4BM
90BN9VIadDLKZ5iB6pN4pw==
`protect END_PROTECTED
