`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAUGE2kSXmpDERxUYa96LYUKPEwvzG5b58N4F6QHdhz6E
NulumRwLoKZy/OWrz8LVWWYhcOZlED+GhdzPeECVToT7/V2/g+oKwSMF1lekfS3n
vwijoss0cJ/0BXTHjdyES3yyLaOp6Q7B5hkZqd0SzlYJDkk2Xnm/0S7eNgY1qP+S
dS27qSLbcmOTMIXTshASv9wtqRXrK8lkst5OZfRS8WmC751a6Gy/Bd3fQnqHTxdB
WwD/qOexS2eqdmQNiZa3o5I2qvW2KB+iFuIBLgWo/buKYB3jImh7gNk6an3JpKpc
Zqd0TR/wCR9NGS/j7SuFsu49BPj0oxci9JzlK9NBWFriMvXz8S7F5E582/Rd4TDE
/4db2vJPdFh3rCGJVRbyUCpDZllvxE5kSOQ5+xClRQX9J+ABdAzWPactZT2XfB42
ROWWolbMWl8MqqAmC2MGZ6X4DuQwPRHHDFnopUaspZ3dCAMIrgnjiSFA1k3MVjhs
YBxs5he4xt84CqDi6f+VH1s3YRIoScA7Im7FOf2G8+VitgxID8+NKRbulqGFZ1u/
M8e1SBs8k5r9b9JhrhW2ksHRdVRm0XMhkwQ/fIWvgc+APR5KkxkUMvFr0X004Swq
aj8ninlYXJE2YOVhYLh7ZUaKyxLQgG7HBC1fx4K9NeE=
`protect END_PROTECTED
