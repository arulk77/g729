`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
7RWERbz/SCu29vx1yp3KRMXlOMQyR7hlFPPhxQ/qGYjkhJZgilR46mhbgGjRf7cA
EdWQKNQT8W2h0ioe0El+vEwGNLWZeynd9qQUee1nSAXqWhFgNxrVGnxzRtrcbfdL
a8GVYoQqbfsrqjQ4WhIgr7loBIQ1+cf0emegruycsyo6rZ+AvVfurOy/Zq/mfi0l
`protect END_PROTECTED
