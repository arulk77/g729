`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNwyvgWcAN4fz0I8cTsAa6hueELCUlReLdJC7pJT/rM5A
uuZXwpT7eEGa7tRPxqA7kobXjs2PrAEZZ2rjO9qjz9unTD5NYXRf+m7z7o54bIrn
NB7hCakgTuPGYyQd4QB6cwCJsBas59lohagaOAuhY1Q52Diwz7+/rhvdimJ9OlOI
OhV2VFjQ5319LIIDO3+X9kfNDYYxsH2OpVY4LtVjr5zQLbBV+bJGnbkc5Lvu5BQl
aK6PhFY9ULxM+x4UNa3fb4lLsOYVsw5Y5BI/b0Ur7ZhmbYVfpAlv3ox4IznnPWdu
dArJF2Mo8e96OIizy+m6jaDc2Lq66lQFN9b7WltXDq63K3QxS8KmOtX7SNGfkxnG
b62qGGlNFH+Esxi6vOr1c9m27xnn40fXi/567G/rEGOOQZilN6OdRj7S62Wbm0pE
cBD1bfRJhSRN2VCsTIqUEeps5LsnQfo1Ne1J/TiSdgfTsPZxv372Rm3KESO2WCle
2O0pu1AE/uQWAeTYROetUfHvHyzXYrat1IPIW3dY3Fnq/GR7J2tvVpesbsK6soQp
i4h3bxXiu29Ubot1qBP2A1Y5UQ/lSMzySLo5jTwvgWHV8tMP+ypQ613JDNOgSNJ/
/yQT+GI/5ZMBxvTWIybCyBD0rWehFCytw4XyndeS2nxkYDbtQWqZnvmECaToSwOL
uhSHlvBXTqyU6CGzR3QPEAYhojA47JXZ+sPwcwKROM2jwDhp1ICNql6evuSJ5wSI
R3dTNaiq1zOJlsQ+hlBgZcz5RMuV3XwGdKZiNrD+ls0zdLnzRcmXIXPmvYfgHJiv
d8gV+5KZZuu112Fu+rAdm8YDex03dhC/CfEHDgvcb1d9YDf84duEiLabDf8nOO7y
+N/W1EORhvhNRPBJEy9v76Kb/yCW5Zj2+Itqa/T1uGXu6vEwOYxyw6o8FxMj+xbX
/c45WX+srAUc+NtApABZYIZm53/XcbHny7hc2dLtbXqm/I08g5y2xhjvK1o2y3CG
8Rp7rEdFArjns600fgBzTAGYAauKIwknS57Gn//A9TzzhuZ45WcfhbEfSTawq8RL
EtqhGd5fG9WQ7bT5HfJ/vlc1MtwMEyrhdlqegt9A1YFN/nb8SaDxPjMzWrKE5GXT
Rkaflz/zrY/yuEP9ZmG5m3CCg7vbfMU94QhsyWjCG5nM3cL/GbQEkiGrH6vtrvkC
UEkhgnXjco1EevgMi/rl8MkmHZ0NyeLbsK367m5ImkJ75vFC03N/r3htbr+4Oat0
ek5YOgytLrztddzh7SXX6ffuVEDLxqmSMnSGbGtUT00vDgVxRfeXUh4IuY+Jzhtd
3bKgMTUMY5U10CsO6GS1fuBToJakx9XnmhBSQE1GtyeZxadOr4xhteF/j/vR+UOS
v3nbElpgjRHjxEVMNk1Uv6aj0M8xqkNQR8iLy+fWakXRt88ODMh1HO4EO/b25/Oa
j/b2xQrUy8WsY86BINSjcz8M0E1ZIhshCrmpaDuKSIA6ZxgAxGj0BYuic2brRK+7
brdU/OG4Jk+ov1iLdiyquNoCYx0bC0M076QpOHcr7eTHeVjXr8CYfqeHl6InI78D
gepY8l57MtD46821SlG8pb6MejEH0dVb2c+6dCKX6+zxpCibn2NTBtLTx2LNrrbV
2YVOBKOOeaTwxB74ovYdQYtp0mCId8DxPhzcIwUxEwa+bzsFwIo5U9IROS3tFkyO
W1z4xKf/Msm61FwJlbgeZW/npxV+OR5KJ20oy7dLeeZVP4cuNIMH11BsQydANu8p
7q43j675PiWAnT5TGIUi8RxOLstm/FnaiIRPKi8YmwFf9Esf/Cox02XGMID2YtpB
FMAgqedUBorDAn2ry2F5lh2X/lJ2/UhkUzDvELLIhREPy6cTfkhPQD+73r9GIZAR
gFCfhTiwoG1RDnQ9iNYOR1Tyr0ERGoLES9PWSTbKmyL0ffm+gT8Jf4jTeUw+s5bN
O9I0HQveVcvLsC6tJxF4CReTSPuxHqu0rXbNJuT3LX4PYQi6VnLQunA2LbEQ2nbB
kk/bfZ3rXvB3MohonksBwHUJDi9EsNtmCXuKXD3b312vuvuOppGPwuRa06xwLvZK
w5H+yNaVawIb3zGFWKbORZtbOn4Qh3OtVTut/EhrWiQFRrfxBiSvL5A+9H0X6uTd
56rXJW9Nip1TpEBwE239vvJZ4Du8dZ9SGQmaDfjl6AsAW7p6uT/Z0joNhtGnrLii
JmrpddWwz1RzMqUGkp99gzewor8IPSWKBoJtfv2QYJKrPAcRlPxf7P9wMPMqDLVt
SFk9FnEHWAY2xJR4yLHR516MWPN6Lv2peKBIynaYVnhd7HkPW5FUvKWLkNnUuCrE
Bc4s6s68Aggn8YWHyQUfDnTeg0A4xiXTahLMd43+94RqYQ7pZFfOrPOm2c8qLs0u
c4CQSMkrGHITQcjxwg3ay64dF6tmYESyRL6o0pNczPZoJpqj4U2kcR6Ntco4eRdz
uMHV6rpzZShmY5212WLoVwBLEyALauq9G/0agnMRK+AXxQYEcD9WppR6pLYVV1X2
KC90CnRTKFBO0zwnmoN03zJ26nhmA2JfjI6kEq+i21pMcl8P4C1Gozk1ucFwTFkA
gTV17Y7qlAvtJ4BUBp0Wloci4VtIfl1wOK3CqOBMu1zymyajUXNoopF45/Z/+OAo
lpDBN8eAVbH6bg/OwXttanuxee69vuyAAdOQy61XvSeruuMvZIoa1w3ACxKUhvAY
HU0i+bhazDzpIreAWo/levA+mKeRWpSbM92ZtEgiy0tQuJF+r/zqP06duzmrnYsO
KbP28QWY2MZkYtJlUjZiRAzzEJ6g5n3PsYlUF2qKN3Fg4jpHHfYhBUWzGV2FprAG
f5sDRIbkcrpj3q5vCjnLiu66MMe7M0cZAPLIhDnEBlQ+z9vyU/w8b6igGtl06Ak6
U2N28jFxcJWm6ohcKXYRY7BYHQRc75ncndBboG7etumPFFZgGzru9CxP7p4Avn6k
WQ1iDmQxmha7CKqI4bfhQpEZdD+OrwFvRtCw0lV3VhSPG21ej3x3OUk3bPtUe6BY
DZnozh4qhlntdA/Or9oTgogXsNVwfQma2lZTKnWZXPic45oG64Ze875Am6gg+gdF
zFXvpV/oeinjJibYcYlBvYgpaoJeEaKgehuS4lCc8YjvRSWyT7mSbsDD+SGnetkW
0gPBH3AUQHLssh/avceA7oS71bKuLsfF8Y3Btc/FYkoC/0zHF96qEK1xmgUy9MfJ
jMBwqbj5gmfjgjEXK5O7FveW5N7dDk5HxhEsrIb07w2MqZ4QmrvhheZzud0gujMX
w5BJHgpaoRB44NPs3LSndQ9pcuXL9JKwxrnF2RO7tapDa3fxaARtgE5EApIy77Mb
oCxC99BLa4oOKKuNL4IktSwogPRMpKgdcKaHmgbOIIsJU5TnJOnRQf2EpuyPJGbK
dV1iNxbcn+DAebKDtEAcUFEPUN8FSVAv83JR1teyQ6lnbpD/kRxve3jU4Wire9nl
ymkAF7x1a3BIr8rlyOQo3JpcRspxrtuZG2WxQUQK7TXiTNSL6dbjt/3e9zNslVrb
zTRg6IwWPQDwc4ECSgATJVjSZ6BxUklEDucR7I4cSheFLm06ZurChaZAEeNlT/m7
uwWPrv47P1U0H9wFYu6QQZQMTvhQJxRf4XQYkWm4ZGv/Ph1/ruP/Ex4EkRTJaF6t
9myTgTTM2OjmEYFlHLjGzPBQhXew9rWMMpi94Tm24ek2Ym9QjdLYwI/JSRteWnL8
0q2XacN5QoAQTBy6ySTBbBKXwaZPFI5gGARpW4T5fnQzPynUa5g0fO7HCnW0jb9e
sS3ySgWIoijwaeZakMgCbXhcy/4jopWjZxb2PXhVYPrGo6QpM6wjun5CjMusAn35
yb6f08/Lu25I+dU2NtcdiuqGLlU3XEWprGn15f3Hv9gRwp2IfvA7ZmKiEF2k6IAY
UVrSxx7w6UCLOu4WPYB8Rv+r75m/j4V0ePQTv9JPvcEGyqI0PIOpOToateuDgKI/
RL3cukW3WxTGLQmTbg0g117M0jZ3ElvjCbSJk7HTOcUudELHcmAs1b6Rr1FUp8NB
9z8ZjOR5Ts5vy8ZO+crs1KuqK2y/AhTzb/nir6usr3/sSdhDxp75ZA/Iu5bDmSoI
PsAvoruSow1J0yLZGaIQWNgjBqTxhCiV25cBtiyfa7ZL1BF+dLuE14/Dwr5no3JM
UPpxraSd/Njcu1g2fdR+j/ODFquNt8ohS5rzK0+f6IGNTAS9+CRVucbBy7axDey+
XB9n3dCJhbCfkUf9hjflmeeeKGlfmHfCuDC2vUgMm3wovsmC4rM7+NlovDgo2kq4
8wurl5D9HuSUcoLK43d8yZPn+8N+tQAzbx4mF9/VbFZGz6GcpkFsr1L2o+YkYx4h
i9HDYAAm2OC4nKwiYGyNb+uJOOKz4KNeJAeFYuU2blCy0X30G5+lBQx/jYzfQuvP
BWotcEX7EM9Dt/ZoKAsLPuXWzSwSEEu//Ec+HdARZ/+AmYj5lRPpIjW3WiAjTOV5
uP5CJeYD2xiQgAuU3VM8iWPahq9Riw/aH3wjDC5NUz4D01kwjrIEl+SLA2WBnn4P
Yab4I8Qr83vfwi4iRZKMreH3U4vmQHftHknE3psb1lft+cE+LtL2OZTAZA9ZQ3C/
XmKGAaw6hwjvsSeh+9g0uQ3KKTxbLtjhXPc5jqbm8+D9Sj1HMKNRhSa7zAAA42RW
2XEKZqI8wEv/e4lvrg0wz89m4IMhwRzeZxz+gnmfUMI/P0RobslrHuW0lmLuCHmM
GcsKI7Z3o4NjRqOK/P8H7NFXxXdKY64rFs+3JMWoUC2CpJDn8wvSPDEFAvHe1PYZ
WY/LfGIT7HmzJ47SqsL1LQuDII3SWxfzy7x0U/fA5MG/vG4OKY5Wa/L9tvrymm6I
F79QU1TUXtPDRoqSx5C6fTKy6qb+4xIvoovXqZTgjT2O2yP8VdMXfbWnxZJOqKNq
Ui1bDPLh+yCht05EL6c/rF0gddUmiYyNR13nLEQ4rEikiRrJA7/7HnI2Nj4aBMJ9
8Va7iiR8C+eHTC4qZvi+vw/p/PvJ64VBZ9hBi7p+jiLxY0Jlgvkai8LvhVe5NLCv
sr2XQy5apwT7aIXwuC1KJetPJS1jDL73TJVY7tV8m7GEKEDMBgsov6QlHH3066ki
+n1upf3rYMeOAWJCReirYLm+l8FGrHvETfeNAoleM59Gq3iifC2Kw94UgXIV2u+Q
ImDdpGJjPDN/lr5/uRwJmte9Qu3EkoTmoaxyNPp9yZT1rIkhbQ394W+sy0dU3qTn
SM055fpDFHZdYqLZu+OOuucd/ATsAQ1I7jFrBj7LNrAT1hjD5/GSR9FZUKaEsuY3
nBEzXh+QPoSXQcyIsBk7Nep5csIqg6fVuNyMggPfmb/rzE+4rZ1yONTlPbvruKbv
VBs9ziWus6Jq62Q3qgOxZ1TJwxXscanLjPn0uH+Byzjs/GEXL4bhN8YquP/JNJmY
cQbW5xwMxfecqEHl/nvKCdcVijvImmCNeoYcbTjdovpX2ziitmf8ced4dNf+aQ+w
4+fW3b0YilCTsLSbGUpXLyaeJ9Vp+9fELDijAfVsVX4Eqb91nT55+vtrRulERWC3
hM4PSTgnASbGq/nzFdfES+WvPQnpMjwnkvuZeDylkEUd6zDh5HaT7wBmkS9svBvv
atC9hDqKT3VbNCMkIIKZ88/isA1lCU8miJXakJxy/IQ+BwmDM/5BXCrYs/vgQWtG
vCbi3BS7MJDiu13Fs9dElWszcpr2ZEeG3RyVN9P1o/sAFDxMJ5cUyyO1aVwAW+56
bQ/x+tqeSXXapl2JsQv0tqclS4SSzjwpZifDrw9GNPHQ/1dYWa/aI4etd7AJGEf7
LxyGXdZP9S9LBhZsFzCWNOgIrhQHQDltgymnJ+Ls0psX9pVLnjna5XjVSwJ7Nvvk
gvn//+hbAuEPkVS38Q2Ku9hR6C0m1r4zAGBzK3oKz1k2rkjJskk0Rm0SOadC9sqI
Euy6ICckffnaxvN6blTLtEh9qEe+TKosfh6nV+UjfsqAoNvxKXlitOlZFHbsjHAS
kjoNWNKQAs/3s4TgTHkcqQyoV9IBz2qg7wZBKWm32U5MpKV96ZsuGX1AcU4VUKwE
wc3eOa4zHOrhzfKtRftQSwUIKcTb/2ZfGwnGTTK2de+vmWAoPNso5WKtvm7zT/Z9
mhbMwcl1agxo+VHBDgLETYrqc9inHyQiQqyhUXC1XDDDLTeA99I6AHbw2mefEQud
PKNdF7J/0SKhC8ubWfnq30sqmN8yJ9XoE8CjTVqvcjzMg/T0ymsX56wK6+6suOFp
n0RnL3SCo7Ozar6LonC1oEZqHXpBQwuSj/U5KKIf6NzJ0dHClFfKt2e/mNFWg0j4
ILShqLnf0a2L3lxtYnAmR1cRKisheJ6kjgQqqIpm2SWiv0BDbLnLjPDDCsxk41KR
ZWUyx+plAXYfvcDkjRazxqHG4AvKLWuwuhj6udyO+kbjn1k79VRRdolIoP6Quqqg
jGr96Nsf3WffvZkGQGB2PuRZ9dsumKpEDtdsGTRe/nYAJfShNH0ge0ccwePQxs9O
Esyl1ld/54KUq11DQKNt3gFsMGQ3o/ncK98LUaaz01trcZU+Yx1cIY+kysEdhnCP
rWsz8ieuY0YJSeoMppHU5HdEWK6tiTA+n9kQKdeuh9iGej7QK8vS7o/ofTEZT8/a
1OqqLtYrvSDbw08CyhhjY12OeaOpQ8kDGCOvO2y9TcKaVkJUCzA+mqGKiUHaoliu
hPaebS9eApncb1/92EXVgI0FUZ9/DcgtaFhtijuqoAmBc+h1zDfI3PtfAqzobTIr
1QSqgxosSMELK3Bx1bov1e+nUWaWdz2u/8lGlY+TepPMl4mw7v80bUk2xHQv/T/r
EFMKnp5VlrpzGKF5tLeUhK4hd1Yn8YEjXUXxeTvkGQuMTTVTHDFFehaHFPjzNVw3
hDvpJ3vnjdzfAoMBtdG0X9iqj5EDl4phOHEIWd7pPCsSEbf3zPE0Xbm337wAmRVJ
mz4tEXqH269FQS75fVOFUYnwEV9jur1bfxaTNnytb3mZxykvjj5LEIFtQmIdNW65
i3IzoZfo5Mls5dp+mNlU1vcbIfKbZwRKpgM4/4OfQFYrZ5lKfF0DHHBTnRVa/NzV
a3cj3A1Nz81ng1qLEF5yrJNYkHpUkJ4gQxmzOQrwk3cEJBwY2CzKeivRmKEzML3L
xh4/sn8ghUSO1FX1e6uSNOIXURxeuwGglWbHnqidzQfPS/KQtxsA/8Kc8mC3UTN9
Da114EIO5z0BmyXIzkkZBXwyvmo1nkV8OGeLy3PKN10sUVXWB/thx8zgmztEZU7G
U1j+ZqyVcDs8gsGz8fjVWg0Y9OEmmetNG/ZTGSvahxOWo5dnRScwHAezud9FKaHn
HIUn1nDj58Oqjf47BKPpdF8FgnnFVtRiyqu38RJefI19UR/+XwiKlz/yqtSZg1JI
YsYJ/Ia/oyPScLNDabOtz6xK1MNDRWEeshs6SpiajTj/xOf1IlWMzksX7tnsqLWI
NqvurgtSGvdlmxUTl/AvoUiDJVXZK+LbXAqmHsnya05t10vWHIRcs0/j0ofwgAUP
3cPQ2kfHvwPD22/EoJASAGy6PF1VekVKyKW+0wU3J4nYd9TDhlxjGwfvczLsjsuy
xg2kvfXIYT6fQM1qH4dTVufo1Io5t6bkglJbFDD04b6/CjTvTo5ls0mueeNwFY5U
PWGh3+S/+nbQ0fueMBuHuaIvBZHC9QvUl3SmWx1H+4cuxpq+iQfCOJzi2b4wfPUD
B8i0dL3/QxpLaVkkWuRCMNLIu52j9jjy/JbQVaPFt0TzAGbl/Js0C/+VPj4vq+nq
mAV5Mq/O5iRCGMgRb8wvDXwozhrRG7idQhq6DWQ+ctU9zRsG0aPJZM2zvOEsoY0D
t3Mu6t4sT9fFsF6Ekm/97gLU4rHgheKKyw2hzK0lBZGXQdOpFZEJpSF6ZTS659Ev
V+GhWDqVP8AkFoEYd45u+tt55FQ8BToxgtsj9ZjBXArhiqIljn0J/8LJ80ySjhIX
yb+I0EsF4JSgn3GFnpnaMU0UIBuqhaXg64pF8tysSv1eYiKf4ZZaopAi1xC64zeG
yCFtYLwwxjplUd4WCzEW2TrrlUwqe98ztgao7c4D426+8EThmygVegNEoFzB5ria
LKMJIQS/BHzIZZGNsHzyfdoVWiQAuBBU5lFlzi2kcXiSHHcrtfXSVtueev1YYsEB
yPknWHQe6X/Xy/fi/jz4h/tAcV5u+NB8o71E2h6j+/IO3wWBSovoGa7x6Ymor/pv
CKztXQdOJSpHV5GY0C40etiWi1zntzV/uZ7i8TXxwfCSGEuGdD6qUewNCmOko/z8
yc/1wq44HwpVBn/Gl3J6NqwfI0ErkFq5VvOAxMzEsug1O/l9yL8D7zmqwQj+mFHX
uTTgDVqCZKdLgaIuM0XurzqUx+sjxtacHlDVZFtps5dD1HayaklfjCD2xV0J9kx0
sHgA4dU2hIeQH947Mku2oK4Ev2SWU2sYM+e+7dwRmyZOcNKH8kBbN0HU/0bl8sya
FWDhAqmQs+28IFH66OoG68kUkGVK/FjboZWw+2D6neIWUI1i5tCbEsqjbU/qsrBd
q79MuIOQbPz6PBr9NDd5KXoy8AeuUOdjVroMgHzNArmDUVhYJGf1VvP645Mu0Nva
eSLENrI4hCZgq9u+baX6LUpiTTralVnVBuVqiagcTgd7xKygMKNDavWj8/WAvg1P
SsWbhzzqz2IyCPgU8ak1ettIMHIT4ORZi2+u/TpkVWp3PGON0isFMvedZpCoVbpM
6Q8f3t1dd4E5lrcqv2zCakM+5KwJchzaLOg1wC39no6RZHEhGzcnbbTQ2k7XDfDy
3Xo7eRf1ovsaPuMjy75EqLr33W2ZJQ/WPG/EuqnFM7K4CZ3SUaClLZyaBLtJvcuN
YS4qjD1BulPRL4MCCkagZv3yT+r2JBVqfD5hjvGcRyH58+2G0qUOOttGb3uCriql
1ccaIU1vbpxrAqGDaraF+GZVQoAG2c1r43ZeSf/sIEtJ8xrYt32AW6BsT1NakLYO
k5nEac0xDRxAaOc5Bc5OZi+PwVedoFbOy2VzdpaiWOYAnr5lOfStDFeQr2rvQprB
kv/0EPOk4NzeU503h6ROa9Gy4JIqQ+zPYTvjCusBSZsQId7fbWQSIkrqmWko8U6I
`protect END_PROTECTED
