`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wLRzNFvf8b7RTpGrjtGF1UOXcgaJAvPkoFbJ3lknvL4
VG0dSxtZw843+8eHQYUsGsyg2pJ0+x5qI4tXVjSFEmu0zj80H6mY7TSkyAfeAZbp
wslSmUhZmDSa+e2ALlEx8rZ6P8Bxa1pkNrpg5rNX7SvQfVOXZd8gk7WpW69T7c7z
nXp84zWSWZzKBnyaZXXoVdToaWn3HKEvM8633XJY5K0vRx7A9JBPtLBpV8p3/saq
Y3mGSYHb2KV7vXDSqSF1st0oUT11/5Fbw0rtO9kcWl4iwODvmVObFBrMPo1bpnZb
w2Jt0craBZBU4YOJYuSqmC4XBTccnPxLEz+gOXRGd5wJntHJJ8CEoukaCqPUrPSu
js75C1cg6qZb96XewA6tWw==
`protect END_PROTECTED
