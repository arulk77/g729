`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73CyXaYFLCdzdXxAK28aLwMvdkMVu5n+hNZ/M1QNN2bj0L
PdRuUrltWgRfQCT07UftNc5MuT9CknrCyG7BtzBQ8aLdBw8SHhjyv9MamReiim/g
iWDJBFPrD6tcuLFilJ6aST4XnZ1mOFSHUDnQCygskv/A0roEQyfLj6Ux2xlEqJfr
4b95NmUjXfyeVDDIVT7Wm5Hjb2uiZdtmzcxs2KM415J2Y91tRjo3Pz06ztOr7jCS
I1USyV91U6Zi0epocytFYnFoKCKNkQsmPITjhxy8jya/CnuxD2nQp5H82E+RB2vB
QJlRevXTMt4Ptq3CX+WGkWsW+myQNEHqLxB6yPXuQLzGFTuHHo3eof6hhXIrnbKG
WQx3GD0cXY2RrzZfy29iFt2QQnIOMyeCkg8k0UoI5ev4+snAhhSK0rUKAYHDp3C5
5PxNyXwsfKvGstNFgn/9n0VC0uX3mgtCY4a9EddVhx5Z/E9Nmvzz6n2QCyTDEF/m
7pRhL/q1NYd1IbGRwsn3I8CjliVk4Jc2rxOY/6RoeFKxhrc/JfEcfKqh7xF9ahCr
CFeKz5XZc2pZXHfGX0SE7emUIP/SMFawmZdOlnKJlLi9twa07z7lwVfxht7Q0u00
NPGkPwp0d+3cd7zbg/coKbO+lsS7xYGeklc1qCRSCs8L0Tj26cNBjL/1UNH7Etdt
NGfeL/b4Qkkmj+U4Tf/d/OSfs0hyx0iAYX2CEiqENIrTlgXlLg1euf/YdPfTJHG2
vvu9kWJT582FGnVXZkwDruuluziM1SkufSTkUtvizTFM9dX7EngtKEwLrThbBjeZ
fW5kUslCKvMUmMlyU2jQPep5dC+ABLVvJQSZZ8/ea7ULp/MQrXd++wgP6kTfdsPo
a0ETG2PeJRqv7m9+TO2XYazp8v/953xhIRUGO69bMKwu4YSLAgrstan7nnMoPapN
QMijXhR2v9C/lu5xYj3QUOLy22HkGYVxcDVxuMhbyf1G56UAOaib9twM/Z2Paqqe
dcQQPtBCcggPjOGba6sqjTC7dy3R9JUso+CkJ1L61czsZvClPhlAbm50Bp3Mq5FX
Qdky+odbRyJQqQIsk457LFOIVAEUdWYQ1iQnMuoGbaRJN/Ioyyk0dRmAUZQz9BK0
8eI64dA/gzniyJKVj+vFI19Sy/GAEQQcgBEONYFiKXFYTOzbtEcVPoWvnATJrivF
Q6E+J/rOSz91b/ro7eCNtDKV1jfUgVOTQMo24YREbXt4u0mt+36ol2KvN8FHy3Yh
aZJzWhGMPzlCrnksfOy3Md352zi4McOM5k/dDe1SkFp9q4RicRJwlzJPC18iJTCR
hH1Y85W+ZYTo99C+8l+AalhXuXEK9dpek7ZXRxql3emti5TO/1r7Q9lZjf7uGSS1
eVtsqXkILIEyGPMrtLZD/mEsHi6kqbWWBGjqNvzvoYaND1SE/DAe/K59fzmmMuRW
e4W4Qi4MStqIUmmFD8DD4QJu0MDPY2cfDwJq7oeGRwvl9C5dFObhOUWnq/uOGHRm
xc+83eB66WTik41Y70LE/znkGRFhFFV1xKBRV0NWSpESFEJGKZOLc0Min/TKVqNM
AcLNddpOjjWnH3OcjlwYn8+WTtJF1UeT3Cw0gGJiTL9LnC0r/BUx4SMCvEH/XBMH
Ey5bUye/hCxpRe6E+2gDTlDPY5cAQQk/0iBQ2crETZM/8g9U0ObPCF4f90leEKzb
/gJb1UK8o8O3TF0G+xkiQpnlahQhP0tWw5H1SYPVdLhmAzTSHBWJr0omvLanA8f+
c92m8MwToTM6WVs65zaPqkLAhpMXihJgFKUbkTBUEXhiW6uB+tvDuiz5fUwq5pHl
2B1KGaTPUiZylmhHc9gtthA8NDUDQgN8LCQwFi4n+pn3/koOxICx2tJ2Kz6OwMVf
zTqEkN+/8hzUyXeH4AC++90fj0P+I/7kHmNIHAWVfrX0Vwyqe7ZEshL76PGfv7/e
b+ktmEQCBp8nSTHXSMpxlv3nVKQJLWsDkRwtAd4n2C3NGUmJZBKuYzYTm5NnJFJG
R/F3qyUFK+Xbjev1NPbZITDad56c2rzF9ASV9cw50pSSlFZ4pBi9+tqQVM6K53OX
FwuW/1vH+W01HOzSzoNIjhKh+lJU6ZmJLXT/Lac9lua8belMaS9UvDcChpL9bj3V
EDxqbuqMo80p3J5n9nJMV92m3RW4f/yISndAW44tSTEZN6Fqe8V97vwLBt+1od8s
L0x4WLoAtjgcN4l37+5LaPjWnZfNE4/omqJ+L2aoCYmb5NG/Y3hM3HhhKrTRSIiz
CJbrVlZooRFIgXYa4YZ5A5LlhIMRnKXcfTjbRHXxjFQUUW1ybPahmJFEwLNokfOJ
VlKusMFzeNoJr7Xz9jrl/ZNyGZluoj8CuUGcUh7+5qjJZIjxAE9nmMC4V5o8TfnG
gkkUdxPe8dQgpt/SMYgsWGQdbFdIB7fdoNv6aievFDs+lfQEww/Ja2YW+yBJlVQx
AAUZMeabKKyyOp7Bmy8cFwVZ8D7iK24YZKB0GcKDJyLmIqrMcsb/zVlAgpjJxjwY
OaEeuXb3h7RGMKmYjc9lffIZUew0KNpWXG2ZHoFvN1borkVWp/slUQYD0JyVz0sT
WWClttm+IV6E2qQigig0mwF2Kkl33hpFPWCjsA8ipUHoF21od3o7LJkD8uk6W0zt
GADKhcZneDQSh/WHECgq5GfpAsvPo1suR9T6nkOSuolV05mGNkPHlhSFp7mvhDM0
kNtgSLcLBtD+YkNVRgF4YpQ28C9fxwC3lZY9KzUd4CKLGENx89ZEk+FOSFDjvZw1
G2fzsttWU5eRHn707AZYLa00HoeJhCmIYrIe6y40sVk6oHOH63nAq92nf7h54Tjd
ykiEe/hpHfg+8LTCNSNJstsvDAAb9Bt04EjhY+8CdTypPHT5gvQpFwKNVkZWr7FM
G69yrbdyJ26/rUHZYB5eGapPejfhJcfHdjHJPvZpTnxF21Aer6E+XcAF1jZWTwc4
u3ycn55rtTuXzdiwVvYHDm31gAcKBsBgK+jqzTp0CvBFQIT7u70o20syyHwXHs64
shbF7YWy7sjQb/EpV1DK4FwGB+TwUDNVZ9dlk68jm0W/fTStSiHsQb0VzSuLyNsq
DvXrNO4pPwHxzrhL5t+qG/INvQhXcGCOGaLtZQH93uKbrb1VIvLdd2ewpQZBz6qZ
zW/qi2KcWh3A/UnElIJomokrzHroBKjktcTrpOEeoi7Fk1gSMdKY82Eoc7oVVVPT
ane5+jBVei2ZXBCI4b8W9DcT9QoU4eYwiWAO/cbvsP1vPA7yxtpirqhm+qgoc14r
VeHChvOtgeMzN/VAI+k3EDKSbDGEK4ELPrKVha/PIqbrzxddsOT7xONIGIn3keyn
pnJokhnNhKtFhiqpAOwideVXM+VkOFYlwK/siFqovc8+DQ2t9aaWxgC0kaoIPITI
DXYd5EEGIvGgymWZWjyqy1mg0PSCv9QJ4715vFUWExH5N5EPH5FDZ66qQMkYRYgp
5SnrTF0HrvOdhZuwEpMyUo+AEV1tVLmsgTUuUcQ3TUTBcr0eFPzvJLNIEBA08vdA
hDyfibFHaoiXoMXtlXK1xTYZBhOMYqWVuvRUsdpTHepnbrIeqzvf5Kv4ftw8cZqQ
lokPufquIIWWK2ynPARvnGQSm2XbsaLyK0QPVL8e6LuL6iIpoyZ70zLBLwSjQ1rT
gnZjRlzmoJY94ggFwd9dFviNiNj95OkZE+ElmJSYrO+/VNLD0uMRJ9bCSbMejr0k
88HjcfNb6UOeg8g46ohIjVcVIP6EQJO2/LCOTRzOYs8efrm97zS3EoMGP+dMItBS
0o0zcMFCSVaguhyZV+VNsDRKHwtz7Vz1fhbSMdmUXNUEahkjy7liA21uutMNzHCT
Yq78NUZzoB2l/I1TzIxFYieCe0xhS2Spwba4eE/Ldw83E2zTVgHqs1uyZP+nJbiC
Vj67Ji5tRnAYLuaCKnZ2E3l3e3SATGXKKenEk3MkYjxiQDQF7NnzU7QzbGATsW47
xqYexusyjOYnNEodGj3yq9q0pQIvBiI88Wy38f0FG8H1hjN90arA7d4EAw4I/Pzp
ASSBaARJYBXGPrNqTcU7/7pC+NoNtfC70Q9Gb/rb3uvNhYIsy16HIpFtmIESnI2F
cP5NjElx8/ypBcl88rBLSf1tvLwG+6Q5rg4W/2BzIl6QGlFhPt3KL2zsO4U9lA2O
ESrDkOpoyJQ/c4Qp3JrJvZQAN4wl4p41QbXuK05tjbTa6Kz31P6SGQW7CDVChwHz
zg4mIFR18l0Cz/p34PS+D3JxT7oHwnpon0EYQm/maOsfq1kQJY68kG1QavkA6fAn
CRJKsq1Sl99swC/jEsBDL02DxH+N36LIxDiofz8Fgaw2H4pGIbWmjm5avjNaZNM7
Plrwfu5OkT6ePKeUdMgg6OzYcIVpMDXdPUG2kMGFlLc2oZxHp2H042PwNsnXmvNF
wDQRVcjW/eHQNPbvXxDxtLQenj1ebSFARp/+3Yl8OrC/8aAtwwKwxmmvQbIGcLyh
Xt7Q0KkYaznfnqGt0c1BPLqqIks68GodJc8wmeFr1+RM2BK365YncCha2MSVGshT
w30aI2MwcoZeGazxvAWwEHqM36rPWEWTRQdJHgzu5/AH8aJXvTdzP31owzvJxbva
/AZIXqvqOOjm1A3Ixvam72/o191+dDm+hLb0xWXlSKR4Z7uNSJ9sJRpE78SXrp9q
s7JP4f7KJUrkXSv44lsUsavjR5RxhIp8KWtUQX8PodAQ0CxrO5DrdjUJJn0A1eYi
/8PB/s1EFCi6Y9ZRZmI4xuP+TMSW9pvDP5il5qf+Cg06EGH7DI717SpxXueBlwFp
XXbth4v36alGFuK1RPnkKyOFWfZUJafnfQH6zSK0h4ZdK5+Nlj8erK5lVIVMJ+b+
lsitFuhnwXzTvE0OVz4bsurSUthx5b2MZlOKS20sox18r7t5gpvKP5iTgOd4L55Z
sTpbxhGZ983zV+5rio1JCl0DgnIWZ9m5gP9u6l7KY2YG7VT/fvvdtuLZYzR0kFdE
kIjBu8cP0FX+4V0rLzY+1iLDrPbtDygfZtFfTeTZynLhLuTKXSnUKd/WPtEHG3Ek
eeZrRvFDV16zWw6TKdaY2EwuGMxTB0rTa5Njq/8oGwa+8tzJ2HqqvB98YwRuROoH
gcV15l3Ht3NcITTt0RGtQtXAbzhXg11WdT+wTu5htdaC+zvx5ReuzuNUh2j2TexS
vWSe9QjaDKSrjLLdbueBMxGajfpzvABm2tvaPt44HbBz2ZIqxks8D6wKlMpkHPRy
9UHrAIgB7rncjlFRoxVh6ID4QqQPEG4vv5k4XLapBvg9tSJsz8UnoDkaEyXyeHby
fclOD0a4LquGrg2a7E/SscqkRhtb1F4Hvdqaf40ACIpVw/FGZJFzT6cs+rpbwMEd
aY5rWOErHe8obt9VQ/j1O5e3YKaAanjKotxPVC5CfVOKreRy/NMjmxtOI/ZUdArC
yFcPaVFMNKhGvIE8Zr4IlO2abjuYL0kWaKLvcMO4EwyrG2LXzSeOOp4aqHD0tIHi
uPqYAfNXVMAoylOchFlv4McB46KaMDT6zOehUs8TOOsiY39q0XDMUHO8XRfiYODT
kqd7Lp0VefLk/hV1LBLIn+eVIo3n8Cak5xvDJQSKzfV72ag/m3m+Prv+il4x076Q
8TLW6vuO9uvQDbboiwG6DDNv0curHKqPozvXRCCPtEIe+UkNhrRm46PX1ef7NKOG
s/mQImnAy4hNxGoQmXLgqxeL17B36Sbp6UuK2ibZNEwJ7qcJ96pKDpXqSUOGVorr
REe55CD7mcTupoesei9U+9bqUJVEhxadWDxkBBVPjcAvG/OCz1ReuFDAvYdljkoc
+cg0zdpTAJT+n2qVcIUB22RoGC5BIKpwDq5R+dDfd0DdbK1DvcsHu6XirEm6YVZh
0jPC6azjAPapFSQrOw0AWAoaIt7xheifOOjuuBxjSjBa86GeovNt4R5z1NeSIQed
LrOv4x72ISRVZn2htJrj1LcxOozvyMGsoUNgCug9wzfDOpnTNICVJzPUpqTByDGd
zf8xQ331ODGmTeN8trnwlstnbFyU2QOfEjsZ26Lx6fvqVcWx+Fd9Lj17NOba5bL0
dQ1RtY8nKEezGWvXhuQkaNx5vJn+T4wp1HMqvyx3n9eDX+CtCLo7aQtAgJ5ZkLmo
05yzT07jlMsl6K7VwgXgHs6WFJzJh0ZOQC6zvi1d/bv4HMYhvZ5R1fZ0zGmlciDR
bJl8wmrQAxWqG2uFpFg4lfJJj4T5uaT4+XKcNfgTHuB0Fx32U2QFQTTt/gQO4EtA
ok3S8MushEpYR1m/1CYXf6A9ocff76m4vhSiNn7CdYbX2/+226wwduQ9KI29xfhS
Usb7cZM/kltKFxDGHVs5Ybie1Srk7VnnsFrbjKI5zh0iwZIt60gqHYw4KDChwj4d
Dm29AOHnV0ci1ZKrrgDcWO7YmlcPSiuOX6k8qkBQGX6pLQldAs9I4QjMyOSUC5dt
ACxIDYXrmx2Np0x9Cg2cOecSmQsmGq1+ifxCYzg7mJxkdMNrTzdieCahaDRVQSzm
Ofzmb+My9Zn5MNdnBPJIg0YuEqpnOeSKH2scrXZcShuJtKuwdUMZWSZVE//iwk+i
rm560WIfI+V0yEkUqeEGMdmYbb5UweVisk8poFlD2MV6FMqI+/pApwenti8c6OSR
5lxdtWU1qEU7TUoVcIPlZjvV4dvjDyT1+IGNktQP9TS/LqoGxqx4377HALEQh6vk
5Y/CdAgtbnW4Cx0GSgNJZBl+nGxiq1ZAz7YatzUAM9Q4T01D2FixfUQkf4Cn9Rfv
J9SYKJlkhrc8+T7dbb6Mx+PqOGnfTJZJgOQKenqZJ4IIUnNToTOvIAMR9BB5sgmG
hK4kkk3P3bT9oTAOckrRVJ5ZzGmwFekA8IiCfxtkea8BsG3wK4vF0ymn6sAkyicQ
NNdHbMrkCmckSWnfzVurGwGrk0zL/JRRJZRg/5+smCtxQNiK3wdLmVl55ExuQmlH
2bNpzm5HotTqhAqNf1b4eTqyYS4M5d3VL5J+dU7/UuVwyoBRyoQmz8h1S755iFNL
UoNWO29PHz3SPoaXnHAqLgUf9ak2q0HEpuxDimQNSZgUVPRUtf+iwzK35CIK/Hmo
OSmEv7Ize7zdmYAX92jPUtb9QDvAada3vKF+cXQshnJdH4a99zAla0NQmNzfWBhN
HCEctAPOLdnQx2JyYStVlMbEjSpE8AiArGCOOyXBgEFYDnbQCLTfEO/WoZHrnItU
Us3W87G8LGxwlpocDlTrTIVcAhd0cDe0eClBsbto+nTERSHCDx8mKJz9k7O+onFF
ukVYyu7eEG0oZt0inyf0Q2Mf14a58ZHGm8YRR4iTe2/ewYP3QBvTqzXvnT3lMOOo
wlob4Aq39YG79M0M9r5nLhmExE60B9ShQG4gJUXfaGWvI7CpWLud/n+LZd8u2fsl
ihTcPf6Es0Ugb8+mWGoma3vRUcqmf6zm10frHL+T6Do0feYF/JLlvV4dffRuBr+C
y48zJnPvLb+3D76tp9wsMH5of17ZgiciBHzbb6r+YDT4iVvj2eReVdqxpM+iVhNt
+u8TeX3QIUD1R5RWxwEI9XfFhimlVF87tsCdR4BEMj5Wqzmu8k+2PWTb6wYb0rua
RiN1qAfSUKUneFwVuU5UEwHEKIIUH0bdE7g5wKmvuWvmO2HgbwdXDqmHjgTFCpq2
GkwlwxV13AL8V4j/rYWvVaxAEHo++N9W7cRqqZkRO3oXvBv992G0TgrfucB45A0k
naMPjM+uuksqkBoU1g1qqgqLtmFNOYl6IFDbOnDiN14lCfYVsJbdk/I9AU8Lu3ah
7iBhDcm2BCGHkefv7eV/3mQIbsfZBuiAHPr7T3jeQLghY53IrXncYeEDaOLBy5dN
whRDnF3YsGn+fUmgu+Aye/VNVu6F/UCdNeKS2Eh9FPyUMfy5jeTwQ0HjT6tDH9is
zNphE4ZaDJMTS/I3jWO9zlwKC9Dl0Be0Lroq7+ytBwCsjNq9zBsoG8fUN95lH94d
Hte6yCuj+V8UO+m2kCFSmwlPglTo4cPsxFn205pkvkGYur1f/kmbLtI4AXBLtcJ6
Rh0Dwy2TvumGoopECPGksI88cz0rNaBUJcl+6MTLbwkq0Tu2S+lI3OLifjL2UUyD
kYsAKb3nVTpxOXNyMDNzvTpQWL8b6581veNr4pWGNzVrjifKD2nphs3S4XOYtxtw
Pu7FCb2fAuO5EUXz6jy3Cv7UikQFMnQOTsp9JGbHSuxcu6DZgXyLZOiJRTvKbFbx
A69Ob6lafs2wKEuDYlFFdNaeHhtu3dzpThv0NN8EkFAm+/zi3TMf1EC5E/nei5x9
V6cZOoqpqsCMJm948JdOSwEPNf3if++l07EOHx1MRINvTI6YzjEFh+tej5lv359M
cWXpAg+vLnW8tiXhjMcQ++dYh/ybzCzzFKACYq2jF+IVMsAbfGkN7HkoEyq/KAtX
7E4+KoQMwzkqs4ObgRa6044p9K/D79KY44ri3QZkcwArXq9bYTzPi67nrzT89yxj
I6cg/e3K2dA7dh8X36rkzWQnSrP836TpXTXz1Q7SYkDPDQUZ4zUyqhWcHhScGea3
N23qpI2MpoN4FWeihzRUEtsKNZQFaZKw3Hw2Ty+S9D53FBHAcTJK4giG4bj8FFB/
R1OBJ2LzpHjRfzFfcCnbgGYYu4k3JLdPqlNXTPEg/ubS97z665tyOu1wYEowm8EC
U06E1UuEKUrH8Bn2R6vUyU/ARcZ1f5m/bdeGgb5mqtQq/DW2dHIDl8BZXUF94+BC
FFhpmKxrQGD4/vPevtDC5wyTr64LJrr9AtqJ1ec2UbpERifbtzph7PP6dhSLIV2s
FMNUwFBq4LcBeUhyFZjv+TsyGEVDbuUyVH3jJZ/825mgWmmUEHJjJm7DSyvB7BY4
BNR76u/zFfXkHd+2H/2WttJN3jfMkpjDnCp0jqcAmcdob0KDYuBh4gkOz+S03X5+
93qP2VSLZ8nYo9FrrG3MKkJZlTrxT6112P6NiiyiIKOqLx47Fo/Xvtg6hsQyN0tQ
YrYBJVlRMuFJqZn00iEzVDMISS2OV26J00vLuKIZJojmjwPz8rEyKEMIawfRwqLC
U0QlHdy9fyq2hap7zG2ZmE6V4YQCokbt/wupKZkroHdsCI2UTh0gfFa41dHcaDhl
myg7Kvd91Y+A1sCfX5f8/sCOY7E34RPh6JbBiVtdaIA6JKq2o/eh7iGUyK75gh0X
OsYQJKqIzPZuKPTk+MMOUeWKflpfMyOb/2QDhWu6NGHvAJAdfY8dqMRkDX1zIjkf
TKwL9ezXEC3hVR/ZfBRxCMqtxsBWPYo8vI5cy98wMRUdcnsXK27AP4IPHIkcHGtd
+nJHO1jmhegdf3sP/0YBFL0S64BTrOKUy2K+2RvgbCePbfVeMkkWAtmCq7mz4FL4
QV9xlXLAw35uf9CRMdDciARPupPYsY65jvmd4JmXMV5rqW6cyiT8H7uvny7FrCdY
HGnPhAsaW41lotGEzY1y+AC+9zrFfEhKlb9WI44ln7VW8r/GBSC6O5gwCowMg0M8
NyCfPOqHd2gH24I/UlhCPv4FX0Omf04dgqJbZcHnm+/DGUSCeY0W0VCamOZwzQUT
OZmwZu/DymIu9KZSAUGTeprl9o6xXYhNRv50D89JQsH7tZUFCmAek14BwIwZBbdd
iRsTMxYcakUmBoK0r9DfuzbDJlNYRl4w4n1+jMwLsadUETR6Nkfx8YjxCNwkyrf4
Usr471R0OefmdCppLwbK9Mn5+E5SivZN4QcelVFexN9SpOCPkNFaf1z1AiNMplLC
zrGrPc63VMdkSgndCWA4oF7u3OCq4JdquepHQrM14jFufdECUr9AVvNkXJ0Jppco
zKkR304ZJTxeku5ZDD0b3mlSEA+7utEj+n9YETHNU3DWzf0J5gQy7dTQB5SnSVS+
HlchryFgBINcAAUE/N6WB3k5y87HwFaEoXfhbqpqDFvNAkAOeCjtsfPZ3UhzHysc
I6zTYeVmI8mX+creCEHGy3wc/7B8U3SoNWclCvSfMyJa5zg0nkjR32DQDwNG8Gzo
B16YUHJxxR+vl4+UJmbBl2h6l4t+3AImK23wSYFTtukpwYWYvxsXGvNeEERspUi5
98uy2o/WdacY2YDIkKrueDj/JGp7Z3u7m7UE9NwLvEHLWDhBPdWvZGFhn8H8Qy+r
2zd/tsvs2NBWJOy+WnALFl6AONHSTgBZGKX+oZ/LmdQCVz9YvFCEttgsdLI8KVF+
Nf4M32i+NDh7U97hU3oF5SBk9EJUbwDlL9Qh4auQosC2tFsFMQt0GNlCQ01aChTE
KMGR9XnWsfZBWdugVFfyEGI8UiKhRYKrbFMFFGzNpwZgJC5YkOBKgQO2FG/v3zwU
rGNpQEv0XpeTGHOrELupjDOa5zkjfhhinD6MEJuZQE4KZkpxbQGpJU9wcEfHT3GB
aUUmlQTQ5SYdD8OfIc20MtRjRKmd2m42bd/9JAd31TVobZ8AjdyODvdW0cwFA3Ra
Nvj3wdfgvda7e8X3Tzewa0i2plj0iZ4V9nr/SsK+IfWCrbhnlzjNUNXK3FpndDje
L2PLAX2AYMlKpDZsxJRM2iNRxSYOOtjwI0vWcXOOY6JVpKT8n3e3n+r/tPvp3BJA
4rF+HMUoAnlEJApsEktQnnOmYqlqkfKyWvHZaBh+OVhQZClLBLZ159Mb7DyLissX
g9uL5SXhhljYfU6xbORjxM8X/fmsUqcluAhNn9FyBda/7JQ56ssduTd96kK2Rczr
9MnTw2XyykbeXQmuwYvQdE5Vf/8s84EE0A1+O826YldXRCPGVrAbMwda4moWIqkl
QKp7M0Msgc19NjjX1d2StuDS0ItoJE/077M5w8cB6mtLccZxJuh8KZqdTmob6fqj
6cMDQN3jK3BdIgaGeOZEtBd4vjzTAhgj/iYZFREt9lhz8Y8vG+joaz8Qfirkcj8z
PyIS5VLfSllg+7NkyjU/IWO0XwC9r6s/JxlmxES6zZJ15nnomy/zRo4Nvnb08Pgk
AWHiJF+AcOGk/XdHFjH1MjGyjNjIRv5Pa7cxiLleS5TiFMF0h9QGQWz5ClNZ9X9u
oGgamlpqnN+DodYolciKJ/wveKC5CTMy2UcHtHBp/fWSuHXT7SyFUzL2FL5Kd50I
u169dGAu4qtHHby3u9ihZAJ6mn2l6IFJQbjOZnrKscoXZ46WNYhaaF+X546droKw
e+Hk8JAa2OnbH6Vf9Co8BE6S4dTKY+86QobS+BVsDyNfXFggekukMKPMQ3BtvHxA
9+9xaTxocHj2NXq9oDPkMh6ge7AboBrNNIwhY6ZeMBHT/1+Z2wBKv4NX7kuwXOmR
o031EiZ6EP243/4vZo73V4pGzblk/ehhcByWPNGB/EaN1yDiYBBjyoy/k1+hbiDF
DlCoXsJZDMtmBVIMRmBgjI9SL+VcR8fbM/FS2RUJg2pBJ5PoCN4vUkgyQ3m5pehD
4PLcLRsO1KnNVJXQ9iqLEG6vf3jIyBfkq48+1/OGDLGJ6mCrIPVjYLeQ9TgQ9BcA
/L/aXAwHat7RA3pbnEbqgQoDqWh9iGTlLkTRsn2JBvaIXHzJ0pv+oCP5IBA1IqcY
EVuX2z6UcNcJXfwwduXQ+IDPBAs9KBtzWiSlw1PvCPSrtKDTR1FERQnAzlqx/EYP
Lxyveyj7+FAoUlj3aymVdWqbY2Tiq+ofjgwk6FqJFpwagTbfH+IS6mSSj36oOcYk
Mwlve1rCGqS1w+JK963poSezvgG55JMyS2Hl2pl2r6V4koPbL59GCAmXOkbaTcDP
xNfb2Mxw/dk43fEsMGvvdrrClByosAXwtwsWCkWSUMKgBSFb638JqiNUGwCO/gnU
epn4mllnVXd+Z0HD5JrxCfr4L1xicU/iEz8m6RPia7mQ14Li5CGDc65Lx8H/jdvc
BgcopIC4PdKWQ7/+x8lTTn87TDIPWgb19/XRjF7HhDz4yeOB+eyBb8nVy47PtDQL
FiE5giy3A0qJ51SHgg9r/8z80m6wwYxbUGthSDgMyAFwraHC9lp0JjF5p65mXZpG
iXmh/iDqC5jaLne3M13wwT+Ni2HoH69DW+WpDH+YP8RfqFIUYrj1uu5dl/BeneVS
S8u4Z2HImw0C1iYaHy4+pu4GcXJE1AUnz0Ba5m/94YmIwn5vADozbTNxtAttkUZ7
HDT0ZEcYvpxOgueScj40FF+U9q0zLe/90ZUwOFshxwq3rooEHm3Tf8eBOuGdYSWZ
YObwqLzPLi98BQ+/JLRZRnL7QElkv0nP5u0cPltwxiZEqy3ifv9gBQ7c1tj4xKZh
hTdzUHGY2acDriZYJ7+m22WxYM289f+ItIL9RD2Q9VVHcqjiIXlubbRcJG/4B9zx
Zdk4TFPtdgqXZW5iGf/wzsr2/wzupPxek53L5D73ocgfXr0m+Vhv1EmaJRsqhktj
Qx+trmm5LRa7v4QUepZn35L2/ZmhBLKbLUIfUF/qrdv/FX9bxvT9h7shGDYS23SB
H2YnK8CvBPDFiipFyJlyqRUyc6gjyPFHzaSHROkque8PFtDDYtDDhHZM/hof9s+F
o/2l5KNSbWz0Kwul2PKbheIPt0d+aUtnezRlyDq6p/Vn/gS58egIPxtPcO3cEa/F
TBf0AaKlka3C/sscuNNRQBE9qQkcfKMTqoxNOYBC9yNIvgCaIOlAkODlxmMcMDPm
y44dCBmgRzq/cHdpB2oad3zyF3ILm/HRQr6bOkaLJYjd4y5TP8r5wyRUZaPGNyao
sYbCCucPpHlWGB9B4B29R9iW4WWbzujwLeKlrRHEnXLWHr+jMsZKBS8oorFjLsN8
Tqob8nkVxxDuVaJakpvhyhmNaWaEbdZdz3R+sWH6GkV8EdtE9bUdjOEWdm/S6YUT
NqqvGTIh726kDX6HMTuBgMHe5H3PFm/+F/lqNBEFC1bi2QObV9xqG063UueutSmq
fHM990bIzFOGQ27P8ljo3Ek+5QfUy1926g0KYaHQk38LZWyzapnU/g6PjNWiNLiA
Zc+eFyNV0vjSSDli1XII26b5SNu8nVlRrXvGuMqTZ5nhM0Vd6OC4hf5yoRJeS4t+
2Y21ZgW0ld23rYhlbvCtG1UhrsQdcn5ArFF1WhQq9yHHlktEJkPuEpp8/+yJ+o4/
1KpZGoX+5jJhupbFwQ6HMT+u7S6sw8SN4NdBcP5CrOBLT3pkPl8ywlvCllyPcjk4
kIMFnU4JLupRyUyxUZ2BxSjbwskR/R4IJBkg9S8r6N4uFdaUUETydwbkcoDGJSKx
+c2RX2jo55ShxrUIn2EYJIulQvrIQNEsBRSig5OH0CVDaA2y3MGievKU9vYGEs3Q
ln/3emmRO/RZjT9be1WU1GybTb47+bIhjnvjeg8Bkiotpq2XuwvbRXA8vxRhljal
PryV+qDsaJEEjAoJ5MWqlFa3tGuLA1Cu98Tt9GpA84KLlpbnFvDLgT7CT3s+IUiB
YAndHblCXI1/Wg+v2igDLYiCPsLFXr3UaBZbGlPbM+WNX+6CZmDt58nAmonoEeh4
+A7p6Ie5g8tgCyWXSZ27GxzUOJwJrBufZJFM8B7WXE6gSIPp5Z2aPWJZ9XP0io5J
hztfn6WinFvtD3s2VEyx9sYU5CswvHwaJUsEhYggmZeqaIzZjjcQP4awgswCKbk8
Xv/RrLpGqhdFbu1TAwifLZJlHCcvBSLttxCkNP2nutlLVPRevxchOwJgi2p5c/FH
cx+By+IOfDKR3fVCpnxAma5OidpJN1/W9yPmt4MkbDZN7YDtugGdv+A9bwbzSFXE
Si3eGxjZmHl0GvYzSZK3WG/MTjdRNUMwoVqWB8DBuj3WgSjG2jDUMm8zelBUTwC2
GMQAcG7R1q5KeRJWDPjRGA==
`protect END_PROTECTED
