`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOmVAnEOfP7iMFrbtrKiKYvP9huF6+IFFE+U+gjWDGv6
oJS7yKEEiu1trEXBITde1Zq7p8DaugvXLUbV0XTnqerE6ax0pe5hAsavDTUVlzVy
MdXrW3xBeLJYkZqMEotM9rwxL04H/nhlmQ+LFFkfOdsPQPldpRT+Rhk8K9gwLczm
dDf6coytGTrQYQ3BpgmW+ddGdplxSvED0XOkuMHHlIm/nhzxmKL7mmz7QqqWOWcp
`protect END_PROTECTED
