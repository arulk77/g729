`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JS6Ee/OUguv3S0KjECptSMtBd2RF50EJljivspQTgddOLG/kIUf6HRPz9bcrz6Pj
xWi37w5BnoDg9v9Q3v7ZwJutooDnY/h3zyo5UETOJsCq6XT2yoF6vdKpc5nGQkqf
tbtN1iStR7OKdOpO15yAHFFrWFJ//b1wMwJ1BmW+eGiLizRGyQsVsptYhoFpgrU8
mgLhIOUfV63ku17u/SF7ff51ZIQ8ILng+bKe5EhO6/XyTWfjoBliM1RpqCn5/WOe
z31N2MQFLMn0wuE6ws97km3W9dINCb5q5CuPA8ISdOagSbbvKIx0kvcber2Cr16W
8JThVBx0Hh3dCrsIey0v4qwMMi2OpG6wqzxagKH2Rh9v4wp0WfVdgzg1cnOLyhbL
5B4nSnnAGam9Eby7uZVchUuL9RPF7sI82cJ9TEOVnsFnID/xdInfOF1uovIPaJAF
4pGRnrtk3VZuYJ/zsSS346Ri9hxUHWrjUt8DgtqEvNM=
`protect END_PROTECTED
