`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yuiRMVF/+YrvtlPsLTNgd6PKhTuLavbY9cmwPRCtkGj
5Q7e20t/3ekgQ5u6UECVlTVKc4VjDEZ3Ii3LFBcCMC0jXZHRlwhIoef1iIbcyQcm
nxw325RY+0uCQQwsl2k0qYB74f4dYg211fYjUGTisiWn4z6uGE/IEDpfBbf+bheE
ywEQ3WdT5qQcjGc1CLyctAnkN1YmLnBcZE5KQEMCAr3M6fCgmnsFA0vKz1h1WWT5
aPMocD9iMKYZPrB4BlH+8RvzZWrX3EuRJ0IpoSKlEmvrIlWBfdjC3I+7N17DULxH
48EyjqBuLOjqsIgcMJ4+OQ==
`protect END_PROTECTED
