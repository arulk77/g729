`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHblYZsxOHWvdPSpsR9mJb2ifolRM3+Zv8C9e/OmnxLy
1AHYDpcFdL5uShwo1DEVfzfi8V8brXXqDhee1VGwe2yJ4xvvlhzXn5wsQwrHGwtG
ntwNP5lklQ3NjnR+XxV69kRjOO7k8NIWP0IZ1kYOl3g9pYmRzsCthZW4LpkW+5xo
EB8IpFpg6pP5JvuzpkJjuQ==
`protect END_PROTECTED
