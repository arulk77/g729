`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4w5dw7LOcUvxeUQ32ZS7f/RqxiehuB/ASe60RQ63vKFZ
0aefNYvIqyzM+CRbB4wQr+y4Vq9lfH1AiGpd6tYknIBeYoXkoPtA0jL84m27U1Pt
W+gsTTSxN3TB8YWipSLfiUhi024PwpXqApZU2WPb7l37munjzy4UrbQTUqz+rr4o
VAx/fDgzkWmC6eUTid7RnZAbAE88hIv6kjBvaQDjnLMRnQhrKTpYp8/ycRP1pITD
1WQVOPVypRWKN5H4MXkKZ/t7p/CzNo114LSUv0r32mA=
`protect END_PROTECTED
