`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAeQPATC7ZOXYfrsGMBvpOZAu5EcG54H4hV2Zzkh2YA3
3uF4Yz2XCvbipTa6vRXz4JtqGDBZ3skAmAV6rHvoGU5bUmhn3pB3GXddPyA31qS0
u5o8n5tlKRH9aBwBRPxwzRnbPlYby2irj10y+GvlAbpLj0GsoytU/QYsrZvis+ci
CrkB43rKZ9E/WjfIXLst1eQKEqI7mBzr7p5IJ88apVObTdkCuyYYbC8Zo3bSBsGm
qwr+91NodqniIw1pOrR5DDHzn8O81bppYY2X096M3EDkTphArmX1xIy0k6Q9WshJ
UYIvcYBqlDvfHlr2LzpsTg==
`protect END_PROTECTED
