`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48PKLR6ukYCUBW+J8FGbKNtF5Bb0RcvqWlFZwvabLcAW
w6MWmaCuhXF0HmBqbmKFuW+4Ur15P9HE8LqJIe0cZVnrAo0LJco9zK5U2EIfy0J+
o+szlaKAxm9n7FACfar8voVwW4QyBe8tr6YLQlQFMoZ9d/jqIkY41bJ9IE2GlyGH
qX31PQK7ifZj2XH2mtrzCaWKaRsRj1X6QXe1OzipvoX5tgqoapjEqi63SSJVR0Aj
FEEgeF2rIQrGo6N2CezaBN8l4SBhglRFZrubLZLj0ktz0y31IVXQpV4kI7k89vPC
s1SrO91WDXs89wGYxPyZbw==
`protect END_PROTECTED
