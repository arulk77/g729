`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aa+SXuJ7Xd4V6J80BmZ/y+vdNBnOAsO2FV9CSi4Y/1Ga
AKkYoWNaCKGZjvr2fBzDRXXAGlKDG3KM6VIO0zDwEk/+u7bLKaQ0I8CIcxkakpMy
eSJ5Aevb4I/Wz0n8pYQtEZqnX40V4Msg6ZOXreE84bQHcnS+N+kcF7mei+pUwu6U
vQ4rYPJ0afyoDZZh1RvwRJh7TlxuhoGJ3HwJ82bbM9m7I3qqrLiOXXpwemDgEHMU
hyAmMEARMy6WCPeMOkbMIKZn12/vQVrvwjU7CT3senVfW/yYakZII4izG0QRGn+/
aj3Fs+v+NEJw6Sb4EzRV25AtVuO9/XxuL1784omdIV6Agjr6fh46ZrAdw1zVaXo9
pyR6NdDKn395PQsHv5TdwOvGadqVd/8jU4271UAZcaQLOSdm2wrDun1YzazHiEo5
GlJMvuLLprdFoQ3aHqSm3v0Xt8qg7lmyjqp2OuarnETSR+i63uZAe+Qaq1E5+9UP
NmzLSdvhjNEExErs/c4oS7wCPwmvoAVik38RRqlGFITDTkPlPuuTMgos74vZgbMP
h/K7dVi4vGRfYeh3URVP6bBdmsAHpAmbkkndqoJDdAs/hbzcB88EnCHWogI5l+fi
F5G0rWW2FzcBqzqagEynXWmn33skwjvxgbLcNAWuW+R4XzXB+5+IBwaas+W5lIjc
exwvbOGjquRYqaY8izTa1YqW2omODQBJ1fyCcBTq6sDvV2Vi7iSoCMrfL03TtQry
0f7fmhJTZjz/HAY7houig4BqQeVvmyWgUXRFO4nEocMDNSgUUkke4kk8w7bTJU74
HdxBAGLVHrYCcMAo2uSvmSTiwhEri53aAANHY5/AXrymHBdGC2bp+DFQHLGJsfdS
KuBREuQYh57qrQpIrVj1Jz/94SAN+0V2QhTjIhwgmimRLvOTah46+J0fD2xYCaff
QR6gzOJr3ZFPDwSbA0x+rHcGFAsWVVVKYvKq/zeRNHAHxo8DzGBdkQeJTByNqxoW
imSja5rtT2WaVIFDr+I1RD7gT+RfGMAuHTSX0oTnVEz+9sq1oM7GmhB4pQ8Iv6kT
7L3gCuSPodE1+X/O9vSdaO1VbmbLg1ty1tp+HPEXrY2j7KDmUpz3+KomPEVw+Ttu
GQ7JGfbTaF3nQXLV2dmefpVza3Vkr9rnqeG/w2TaUKPHka5AHBpkOSwSwEbRbvNd
mwQ3LEE1ghJ3BN1Yac1YEDHQ/PWHUkuNl2/IHqEKgMpXGaC2oNeM1h3wmPzKvNzJ
aLdq4Vwrw/+FUYVTpZzyvGaEVeE2ad3fT2EdxzVRGO/iSw1AwiSlMbaiFtWjJvTv
J4vIRQdVXo8ku4nD9jjSqmrOXUEN0mhuZu1yFqHH5T5duKms0qkKDCS3KAovmFLu
apfWgTIRtnH+FF+VwZWa3/JK/wKfvJ0s09/9GTLTy1QWr/4LYgTRuasYZPmdblop
URA8ZumFXItbR5PPcyCIjRaOB+wYJZ+/5n2SuCHaXoOx1x1Wuz4rLT8ImM0UbgQ1
tHlPEad3nKiR1fiAvthmS6J2yJddAx4/5RaSmwVl3Hba5SE6V1AA92eBuy4u2Zss
8qNHrjBRSL07AZ0t8Qxs4odl41NjDzDO20u8e98yCGo9FL1UHtKZ23RQ9NOwtK1i
GnOPP4kWGoTQ6ptJswyYRk6HI2tNntm901Ir45nPeMnOGN7/wJ/KKxOBVo4acW1X
cG3D/5Aa9UGyq0a6ISNjSvmbhWva7HgArJ+k9NcdbPUC5KBIbiTLWuEhgCeGDku3
Ypqb+GT9pCE0cyDInCmDcwNjhcRYNFCXgoxyNp4sYKnE8Y5+KD17GrnZXYUYjlYb
hnemvpnL4gle6NOPUoW80e59T8cqcgmDa+l2WJcQGlkGg0J8jqETMvSScvw2Zgzx
mcWTMxjXkGudlNc66xY4UQxEXF9rj6Q6uNPi1R1vLkMggPhD3XRDuBZb6+BFdWyH
kQML00juDyw2zwGBjlP+opcLWuOwcW9/plbtOY/uJkodHWBvv2eSTlKnHs5jcHUi
oDjD/DkhOmc0BkdZHZz87JwEpYQBjS5igdipAIuluJQGEuRWjUfgvq/oUqKCoO8F
hdhfK0jFStnIoqHLaSBm+/edrdhf4m3hqGqouy/F+44EDVWnskjFKm3Cx4QB85Nf
nCCCciaQw4ufnCG1N+Ag6ZDmlkfsxDEykCghflw58FBIaaM4BJ/wPyMI0uaK49fN
cJOnQxGOggs7yvmFlNkvYqaXKragrrgR5P3kNikWO/E6/D+bsi0rweiCkmxu6pLq
fC5q0BcLbVUxtEkOn340gQ6IuSuBWRtDzTvV53NWk6df7mkErlk1ZtbEEy1kB5Bl
bSY2VHXMQSpczvStUjYJnRsOHfTQ4La2CNOu5ZnT7XjB98sfq0PwifOq+K7fhE9h
jVlC3ehzk2SY0lxj+zl+t4cGkrwT8LXlgUFikXx6cOUZFagILMwkGr+z2fLEqn3/
LwOLQHdxgj9kr2xziqUpnvq6MXbFIkarYbKkSJ5kk5nv/AjDIt58Z8XKB/RWxN2c
L6l456uLQN9LrFs5lVtsSO5Hv+evBRNlWN408iaZiDy8Nb2WrPCFRV1TefxddjoR
DJH/cdfNnk5h2HUsOmJC9/9BIHEAQjZwTO5fXisNdDFgc9QrViTHpaIyMpCvJg0A
LBEqGyDShxeNld7fULjlvglvz8wG3OPQRelE01zeKXUiz9i6oMzNczyeeRSaCs9M
lTon0c2/vH3vElTzlmsGt8no5gGoLA5c6EqJthQJaFflWugefWkjgwKMDVkGL8Vq
WIqWn4EUDuNkEB7MbSvuNQQQTyClYz5NoFQYrae77+Yjp+obTecHAGcfvM2rTuo1
xfWxdjJWfUZi2Cfc0IRpSVC9WZtc8HtvtnJIqeBBWjJR5HXP1gEcZTZgRbFzjmK6
8UTpOAN4YkFvGZjILBWhBsIyQ3OSeAtpUqpsxCqksJUeOQ+hvgHzAJrZ6bFX6o0C
DNGc0tMNPQ/3FRWiYSxtSNLC2dVoWU4z+DL542D26GeEK83sAP58kcddgjeruqPM
a5V4wTIY7hLy2WjmacEmVMDa/5dypQRLUtvEi5k+2WwW9e5x1YVO4bBMVGI+a4Pk
GlXInh7kGImE1leUOycUIvwZgEHCw9+7pSZ3PTasJdVM8L5LdJItYMU895QqzfWF
TslJg47HJJ/XpW0GlJ0i13iJm74MJ9uBc+1Ed1Y32bYe8GA8SQT8dbmDKnmiYSRA
4JjryOBJCEFWZ49VypiVxky6jDQmewnbvrNspoR1udBrlwSk0hWFqwDoqQgRiiQF
rGsmGD2pv7n/mSY/JUWwx45A/Mo6d07rUv2H4QIPbXlKn2zW+ZwlRGuXNMILkstu
8JNdByx2IVwBVtymaeV33IiEYy6rz9s9P4/QUIMznCqbU3ZBQn4g+T1DOBxEWX37
dPGsEe1bmU34bclFlDQL0WiLnDrVzRJ/qZH4FdsJuo3SBxUjBP6jrVswLmACA822
mZV/uD4jRUq45F1SfPzsG6k7TOsv4lkHMPIpp0wym8pRGATequiu2vn+Y0SrCUyr
9YZR7DQVWNzTqSwRMSV1QWxwgQfQYhEckKDTGQSMX1VcWZpNZB6eHODkK01zFahR
P9P2N/XsXX8R6um0ZtCWBWmUPp7rCEq/RgHTF35r58p///xU3IzvaglWYkaoPux9
PqLjwdgOtfq4TyJ0uCeSImbu96b3rYrw2VgSkU269l9owmjVk5lvK+jRP1PpcAn0
6FaE9wVQtHgzSLbTUGTy+w7Q/Qv1gLLnUmSJ69Mdmyu2H9l9qgqr+mcvFCYlKhfY
9PWg84Lbhw8zHs78SNLDJvHvOraPq2H3TbExFMLIHFQvY98OwNkFPo8zqzFSMJnI
H7hHWbnLo7wOrmyvPI6FINvzSRY3J0mwJKc3Di40rZ9ezayEJ0lwsPbSevlLaOTu
5zQkHcYrOOYQuMZ23DawEMv86h0x2SQ3K3qJsbDFfdSLI+8uealSebu9KVxI8Cgf
5OLze0aTmKT3VeGhWsvDEqr38R/bN2rqeUicYIGZuBwph4sI9EKqCzBlbpT/XyAy
b0jheGnHwKFquedZs6lWAAeEBPE1cZr56NNJQbwMGXLqWOf5kp6xIkJS1x6kd88k
JA7wLHDRXiaTS9k3Uea6K0jE3zy+WtHu+olTYKOtEkTALx5N4VhA6iPAOoDHBgnn
`protect END_PROTECTED
