`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNyP9NsLTpAAcMpbLrnl4h8KckxPAGogaaM7nPtyl6Ale
NQW1uaj3oPiLsrwbKNNyiK0x8OKfTC9T9D3PXO0FLCyg8NFc17MI+f+momurWeFO
jgG72ff4eZbp3jERJbse/7PDg9oUdVPn2GnXBPw7ceJ5bKvPtQ6fvqvDqqnc3QvO
mh4EAkxv0QjrRbPfpM4lz8Nw/5u/Qt/8nW075FP95PqlofwXta2QvQmd6npDhC7o
V/TqOkxD4VhCiPOBdqTRUjMncqeQ27N4x7vXE9h0U2Ss8GnuVSo1Om5AbXJpQF1I
eY4iwh/D8aCdWpOS3VgCUQ==
`protect END_PROTECTED
