`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
26vRrpesDoxZjK46C1p9Y/o/B2Xz7DUSYfhZMSX7iael4+YS9dCkhWYFJdtZZTsN
xlYS8YUR4m0J2N9mofA0x8fAHCTIWXkWNOwAkfJiKp82rMxgoS3M3n85t0PvF1nl
aD2p4HSw2WS4oiHZkn6g2jT9KJJKmjtihrzXCb/yW3R7+5GmrRAMCPr2qjyB8cb/
WBIXvZXE/ZG3ORjsQuQYLSTEEPqkw/Z09/KjvG2l7XLWVVmjPzaIh7iV9DwG13kC
vDWePNBag+VMIgp15PTMpcm6AM4dH9IqrsUVpTOxa6O2mJX5OQ8ITH7htM05iMv8
80IyrVQJnapc/SCtDuaWhF3OAM8ze5eC+MJiNww6nIS02C4hnl5hBkgAGjAkq8Sr
QjLwD/Tt1ddO0ZUK9w3JrAYwJ0ZWuCHXNlh3dvAwLnfMH5koKqt1HytQA/QS2nEM
n8zfAyUXvqgfdYDsPeZ1uRVLgGKhWFUG7hS9szI7Ue3kW+A0ncIgpPKPO9W/yU+K
ehTHZ1tnMwmkmVNi/jkIrCZvHR3f7kujhJIyTiGGLtBEdYnnxu77HZhjc4/tN6Pl
uZ/hgjy+KZb5u7S4Wum3S/9p1q7WKUL/zScs+r0CqcbpHsx6N7d4eRSpRbxMYCtn
diAYezFZyymBEfhurxsCxf4tM6sBfMrQDUh+jgeiqGvT5Z98DUkQ29RkPhDrq5+l
MjeIWn7d0PEvlCevFjHv6JCGwHlMpwO2pmf7UapoMcYNatV8yQlTvxTQem8NJPKf
c/Vc0y71u66V3ySRewoPY52TFCprZN2tNNADlnX3e8Yazb9uexADP1nqIs94TF7R
5p5jTXr+kfMZpaTCD7G70Q==
`protect END_PROTECTED
