`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
CLXz534f6QdeQ/nwwM725wEegFjLi7SLhGujLrZyRfLZvniWA9J8b0dW1AQX805Q
/yGunFa6f+TajdtXxRdB6W31fOxWFEVbDzGxbkZGv129uD1/1CW96xAygOYsfrfk
IUNT48lvrwoi9YaxqL4b7sUpwz0R/87DlK8sdtQP0UdAHPOr8sWzUGgbIDygAFSg
jJ9uRfkP/dHRagO/Ns6tRk/E6eOL9Kni14+pgTVB2as=
`protect END_PROTECTED
