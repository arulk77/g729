`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Fkp2Hp+3/4vYIXq3LBuREOuZgd0xoSo3AM7gH1jPV1bOztXqwXOj6OitBWcIy5zt
SXqdL3LniUoNAzj1bRR3PTRnxjfzWiXVkYCS397R47hWLuHO9BmqOYgL7kbpHWw3
GQAP22Q5x2QxypNEkeQkHJR2o6Jj5bSJWz1NpQaeUcvNReblnxvS6LcKASFD8ZSP
2sj53atrUt8Hd5smbuPCSuNk1BFqyFziAHRPcol/xfSv3clMOUqYROwd3SUkVDnR
IDktnZYrIbFsRg4pVioZrAUWYmE+JHEicdziar2x4S/cssZYisRhR3AuYjQX/4JA
gcsAVsMiPGUi1t2y6IJMHCLzaUfP18KyZAwekL2nBWtTbDDdi2l5sZLxRCofQQwq
QIObIZncGQtp276EGutxE0S/m/yxVwXsvRIs02xGAQRy+8cl0Y3G0pUjQmOTN3Oo
eNrmpyXKQTW5DvkWHKt93OvNSfXttvgXhlSKXYLvxSFVFVPppGg78dQ08o2l9avn
weR4eT31iNw1sxOxw4jPemMonN4LD6oJJo8H2W3kq51ciQEsd6X0NYWDeAq1f37R
Uk7f6LvU97HZQM7wkaSFRqBojPCpLevam5lmDBo1LDk9X9iYWa/NomdijgkD57V4
`protect END_PROTECTED
