`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBMWzQLCr6XtYDwcmPGdP04zv7Y6l38ue3sFmIxy0tH9
rFj3FlHzi1t1DglrEOFzF0Ia/K+bx5fKvrfNE31UhdpKe+x39hETLn4TsSnAzvGr
LnQ2tCphN74Ctmq+tbZiwpzO1UthE4YrDFgK2RO1YwaS7n/qTwbzHAi9Ak3zgMSL
aLhwgSd/WN9lM1d5uHKXiBc15XD24vz1zk0OV5JFz9DjzF9C3pQsJ62JPlR0zJKz
`protect END_PROTECTED
