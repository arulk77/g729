`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C55Qw7wkfZFGeTQ/1lLaXPzESwTi1Bf7hWeNg449+KE+
0mpvmEjiGBc7Lk/JR5NYvkGrvFsaZ0YmSjERGvQYlgvahmfZybQn2j8hqKKQTW6Z
RZxKaDvYosrUhh3zSlPfF0B/uzAsjDi/mK6le2A2Sk5OqTeK97plcJCAjxVl/S97
WHrknKyjjrrmrITRtTv5JiVrsB1en6hg5jit3yq2Kt5N01PnOsqZkCgT/cINihaO
VHL4nNNKhrAxmB5K2NXCzVL4mREJmV93egvoCmrSmpSV3h+i00zSJNz9zSLirUDG
jgEIYj1DpdMxhR9guC9MgzqvaNz2Uv9tZhE2j1diW78I9J5yn24wSegkLAcOqh7o
80szhkkn3hywZUPZOd691xxsDbvLkFn8D070TabTvUeJ4e/SA8fKfKQO4Mo3wYvt
4yXzUTjcxGmU/ne4MwSa0y4NjglMaIe2PmDEK7PaOS2TQJ1PbLOoWmvfwZhQ9s9+
TAyBfg71ndX2a7g6erkq8pd9xLtBXan22jJdoIydocRhfCFE0M4qC7qWmU/SKVA6
st6WV9xenFn0R7NI8TGJbwFd9VSK0vYLCXz2ozf6QO3fzxogrIPQG3k0/Rifc/2r
8PWhfq0NumcGYEJ+NvSUEO6UrosQJ80QveVhXroFRneEj7beFmdR0JI8WDn0sFM6
TuBRE4J0V0IqqLr9cs6XsTTcr+h3r8UM2lgeGe4eL+En+OaoiOKxAj8eBz02JJYo
/cAgIMObzKKgN+ijSxvlvUtkF+l/KkCp9DYGmGgwXuiGq8wQuDSnZt6eBx0PbQKA
fTkM23gSF5sgxfM6gVCje+H1GaNY7EpkVvZaNKfqbM+fTpMHS2Oc3HfdjL/8dWB/
Ejcy7H/0afSXRK/TqXJnQjZ2lKzixUSHS+nLmnOTBE0ORZgj29FFR3nLUuFU1akQ
l9N4AWOYrqvXXygiFYYZP5EF+iObrwOVgI5sEE9fqyNJ6sgf/iN40cA8+ybk7tWK
FnIYfxctkaK6dq6TMlN5rGzTk1ijKB2tYTZQks4IYAowY+ywHCt1uZax7HANcONa
lZSxwekgakpn8VuDSf88MAiCSsIWNNwGQ1QOJCFRfblaGyoNQHJLQz99MSRHqam2
QSv1hWhQQF15FqqMU2J9Hw5u2qmQ1p0Ap4tSuG8yhbVMizVD6TBTJAGMe8EB+Rvj
qYJehp5HWvzaJqLKiqKZlsJJhVFhwur0lC2XscETUz0td7JzhCp4QcHnv3U9RFAZ
9PakKPTKEe0+ySfkuQfetoPPxf9fbEvoaMQpvOXwoBNcQ4M9+S5OXx4OnysDfQHC
Z33MQ2/wTBqPTN3q5W6STA==
`protect END_PROTECTED
