`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
kOp4GP6OVnvj7MbnGMbAlsnEr1gQnzRId5pTHUBzWIGDtO/umCYyKH0K+t/wnLfM
W6L5hP2npQ4XE8GPwkvC3enxgeP0RMyCEhjSzdcFy6XpPYyXUcqbLVamk6hOw/zV
J4QOD9frt8biqwRQ+IUh87zLrZMoAAVpzG8EEsdikM7iqHmA36fuJ2Ah/KwChznb
9X+Mg/YjSGJ+hpPpyTQdDGldTf/8c10IdW9pGc0TgS9WorwNljkHBpKSWSKjgApk
QUi2NOi5nkuLplLu6QC7niwFryjEahM57HM4yWNPcrs=
`protect END_PROTECTED
