`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGVwdmf3HtQgCduTT5lSn8tfVnRjS89GTzmwsPUMuU49
qb1hkHd9UekEaxsceZsS/U2nwk2tJH8WXO8sWt+zAbFHiD5PYV5HwqcO9W9sFXWm
NvN6D39G1JFB/ot0u7pIpbiYFi/Oe1nyNVidzn8IZLukl8Vxk6akHGJWt19I0YRf
iSCfleJYNCKuck/jMLD6VRawnSqctjnTraK2LcYewWIC8ZLFufADWk+S+Bhzc4ME
jOjx3esTVPEsPDC8S0Bfa49w0ubQHXmyIiFolgIqSfKIQreZPgCFSU8bilTqO5X1
Gr3eClm/IWL5IFg/Zv3x+vqkyaUc4EcyB2/eGOYrsXsu6/h8agOdw2trla/ETw52
GT7QbUtwElEOkbMKTH/eXgb/DdFTJrofgx/lqMWvUZDic5RqRdrabr/vfnjFaaEl
Qc6Bk41KBaswrrb8Z6HxPMZxjxyHcuEphTC/dMTtUyrSSkaX/9M/cOXovszK/kC2
rmyTN6IBmKvTjuu61K484aZpNq5Uq1ColM5oO2/cjyXNy/INaNyzvA7uFTirBbbk
`protect END_PROTECTED
