`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
8bswbivoCcIo6u2WA3yDqDh4ikfn/7tO2IsTGm7zzyg7JvIWFF0MfZfo4bHMaSq1
tzc6MJ1Rcl2FIXZ3N1BeeI0pB7Zt8GGixejB3rVZoKxykw8eScRqlYvmgH3sO0fg
1q4GB23XpeGp3zAK0apXU8KdNZf1B5yU2XvcNLcxD1cN2xYMmXxPMUQtl/hPQQR/
KqgB0Hr47cwBjGRfv8R2pZ3i2BF1ThHfnzcc/3lfo2gR35XqYRa7keNnb81JMJMf
SAmYulaH2JwkfnDAfQr9I/xD2qHijHodewYcm95rvwUKqbLhe+q+ZGQ9R7o/vwsz
MzbtBXvJA3IA+d+rlyWSlwqmahAGb0Q34Pu0nEQP4xUWiMcrnWvoJi2ZyujnGoCy
RO0CbCB5bk3AwBwZlaqZLC7f+xNpng6actMSzmd3fVQRHfii6Zd0rbclpHTfnSDv
CpxvSXo7hoCRFxbTl/IonOIkHHKokYXevnCDZqPxDQBPCEGvCAtsRSr0be34lKdm
AXIyrC4Y4K/Vtj07Be53x37Ze2l4EwjDZfOSL0/yayLd3uIV2EeWPZLQZUTobK6r
N5PgrSyUg0KUen7bTY9qxWKw9VGVcZr4+y3A/byGpUdhouQeNX7Y3JOrEUzgHGF1
gp6yXr99zyXWT6GLuoFEuAFwieGGrW2zzIj8Nu4Vsy+wF7dTjkg6/SqDYSObzX/k
ATsTJx2XuuP6RxXiG8RJmoSP22Ch5Ar7if0k3lNWEAQ2znzHLK2JHYiAntGlPcTp
+Wg6CATEgKS0O1A3DQQXa0bvF+e9i7RlgrUSUtyu6i+XwpMLQJ1BVctQkmnRrxJq
edKepcYfIrLPOjR5hVZL91Q65vyBi0I4ewdPeTdUC92Qs5irywxnH8u/DQ4F/wTs
xrFk5Mln/o8vyUgFxxMTpPS5PkjhuIHyZr5kRSN/te3F88NjLLrF4/E4b0AeQ95d
SOgVmVQbR6DGfn68OMiP8oZIcwZDagRMD8jRXBSQRoJZrVhPyAHV1m2oNDcTjMXV
kX46W/7ABqZ0PVA1uB4LPgj4QEUpByw7R18HbxmdhCXcQGkWxVfCpcHxnQUWWeLn
QYSUp1FMdqV+QTgWTTZvIpE1Zj6xZ5ds3V4L3cdxHxMG0L12NSehYO8wL+xn3hVO
tQcRZ8ljeLDSKHsfb+y2BwhErzhewx+4LX8WILVrk1UyLTJhRC9J1+p7RyoRNrCx
qkugYsP+EOI/87CldxTX9aFZtjjuqC2xUByB1qEtWh+2+K9RGHZCfnJWFM+vyzyZ
3mybI9W1aHLpBvPSq2yo3A1+6UiUnTbSn335xCSoXZvhVsNOYKUMuaO7WPNVDn0c
ilnmEufKZ/CL049EsHuUqoiAL1G+u4btDgV6S9KXxdciGaiuVXZ2/s1Jr+DuczwA
y7ptt9WoHrN7mL1kL5kSCcyUyRT0ryeE72UB0FfRURAcWamUOAetw8l64ET+EkUu
uR1yXO7VLV0EN/Li7rQj5xB9xvFhYJ/NeObrABmbbNJ/M9H0uG2IB/EdBhvqaKdj
SZeNoTcTudlJqsYpwgMyuDoSSyJjoRU6k1D8yP2pNQQFtVvRWYE5O+P7i3Pn4BD7
T8Nqakx98KmJjkqwAVgc6MJ+EAtLZeXoDofsM44T2zGkX+zu+EXLP5h3iX9TIXXa
d8TlHa4yZyGj4RgsiuCP+t65N5/16TYmxcdqA49RM3aFia1+d/fFksVf0CstUxAX
1YRn6Y0ZKlMsUuvNM+f0kVnRo51gyEh5l0tVZXz1R39Cfr/+D166FfEM1xHVs8NQ
yM8KOinxjJ9q2Rkfvr6nMjIgGo2j0uCbgnKqIc7oLAQuQw3Cqutw3mWCXbVz8k/Q
2WoFKIcRQxVhYz+burA9A3BvUula9zUACrINYLvLAejhQe39jaIDc1YP/csuVPEw
97VQ/FA6YxBlOGzxE2u86xuhVcURGQ7mGs21BkLOeUse8qRY0dQEH/Am0IHUdhFU
5qjehhZCjSfzM2ogYFO/Lnsjo5fa75Gu4s/N9m8tVQzu17bkdAklcrqR22MBloet
PPhsqqu5lZP6xXeUvVKn/x1mAPC8z2RaTArkHN1j448iPCBLGbVkXzvIKiAYPJ1i
nr/M9tmwWuBJVCQpHBu4zLL5MtG0MzCx/6Sg/WXSWVwKL8NtHJuXnfxKqoJD8BdC
tAya3eAQOKd+w3OwXmYl2qORdEiDbuin6X7XmD001lbvgtVm5sXMXpx+lJjTnDKe
uTEr98oNuji1BcWp8+w6v86NoHl5qwEAtXH8XFB7/q4=
`protect END_PROTECTED
