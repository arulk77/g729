`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
WyVMlJh1FGOJebGoKBzZDI4L5RApchLa7cxRe1Kd+RdzGnkj4lXYPducCY//PmwS
TkdAqeCi7/NP5FAF0XYAjS+18fvyTM5uLUtib/FRoVVMrgV2IZwhuMFT3ViQcQoS
isyI0ZvzrDJzUpAgP0PlF4IChC8Jf3cdGuE/vQz9U1+Bg07vibEkXqgUgVPpISTU
JIeF/6GPfkxNlAc6V4PgsjkE0x8XrCK0aMZCRZVQ+xHZkidwIYGdikLL5UEj92bB
hAP85wj//O90PdOtBwUS78WpYTwTsKe4zHy+GFSgq3/ANCXmgpDyj9rNkxDvnlFR
148vv7zVYQvJfqE5MBu4R/aanghJBLhA4LhU0qXTIGI9DTtf+t77tu0vtAJr8SbH
8ZJZBgW6xLKhvPkYDOllV9awMCil61Qh8yZoW549AlRXh8cwpKo/WCw3i2RtpBw2
N08DQD4K6KEhNbAB6BTRg78kIMcMPjGvX+7ichpNXlDUIUTwo/Hf3J6lQQefgec0
zVrSbWrAwy8cyuGWj7+SreyBJnOOl+MZIESbRdHt7GUWmC7kiv/jrI+NvUXxyESi
fQYcW0RMdhTZbHJRTfUA3L+/fsNJ/Z1zr/rKBOXMebtGRmTtetbYZSa1RJtJVep6
N68EbzCT9DIjihapeV/VKHS+wqo5wBoiqKZ6wgnxqkYJAQs4PE7HfF7I5ph07+Ys
kCqO1wsOogQbfEV+MvzTu23CBZ1WY/D5iBIuy3YLFhVXBoP8zrkeW80KY6hE8K9j
`protect END_PROTECTED
