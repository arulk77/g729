`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLbKGcGmdNH8SP1V8SOCCgbeyiw7kkmenbOcylyjWDI6
IActjB2s1I9ZvvVmauGTXgEQUXancJoF0t/NwuhRiuTO2DJ8LFed+in3nFH2NGWH
ij8vZvhXutIefaTaeyZAJijBdRS7E6crH7uiIoG3/Lt936YI8mnWJGA1Xl5xkMLJ
Iu8OiEe62+BAbxEn/yhuTXlhTf+iPmjbbkmgrjktbbaTrTs5reqEG56hurSTBf/P
d7yU/wAgFPBiMjXleKawTg==
`protect END_PROTECTED
