`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aS3YcDx1CNlMy6B9boS83n8A49HiI1BgDUATo3k6b7ee
c5MW6MU63JSJaYgKI1ULrIb0tvyZkdDfcrWV7/IVdAk0XH9pPU9Dnl2/hF5Bc2hY
t7Kf0VBvxCVKdqguZ6tjS9cHtRHNIyXyTw4V4w0KHrNQUlovwFLUcE0yQn8mdI7o
cltJyH5yZaKP1WdMDW+VxUTr9GiXGyU6TZC9MVW7Xo4w3DjWkj9IIbYT7Wnj372s
pQ08oClaT40InNuTeE11+JQJ87PwVieRCG/1qXPij2LK328WCKp96xBdWxjfiVE2
BurxdRWe9E97rWcp+fW1/zMRuw4ockzrxZLysCzHXb1YK7eYCCCu1it92D4RFYgS
9Qbe5p04Pe/Tw/x8iHENaQMi2J5Bke5bCfnAva2SjeuQT/ENXkj82Daq13xNdb3s
be+dddbrcaiy49E+nbEGwR590EQdkcW/aclvKsqxIsWy1PC/Vw9lKwcf44lchVyC
IE+fYFAoSvNMQAfAt0k56ONyB25B9xpwBrPCoFTPbpWA1COm8y265LFrcxNi60Qc
1He8dLvBTOaYsaYITYa9fYMhfYfhi5howc6cU0vZeLAfHd8mEEz4LxQ7dQE6eebe
3z+1fgg2aGpdTZWG7AUcBGrQ+GlgCBMGKKfglNhxZqZK/emZp8Pgs1/gX8S/R5jP
W3nHnD8FqgbQMIUMtBUW909hFraBoPd1LlhB6EhjYiP8Igu9gPDsOOKITJdXjt5D
AaXi1V8+lhcsZlKNOy9Y1R3jK2BQNyYYlI0/UUkuhg+5pdygywElY/FrQeTt+WA+
tFWOtHmfD/TrHJYc3EScqLZ8LjUxtDCnupBfdYi10lkghTQBUYIaHJn/HpzrdL1R
dq4dxinNmj1K3MZO+13hKwAzF9ZAQxQ7r0yTdtm/QhUrDOers1YVT/SGf3RJz+R9
J47EThyD0h3KNVq2qN4Z/SinfkfVVUTRtKngymfvTa4Ii5XBJ3jH+Ci3eIqrkAPK
k0QbZaPi3PWkX3R04DctUmAFHityFAOaq6PmF00j4wyrAm97dohcl6CyLsXBXxNw
rTRgpCHrO7Syby0m/Z3ywQdUeJqxL9WZ6BWwHhHv+aHP4ZKPdTyKemI/Qg0rFTa2
sFJRfihLJgye34e7RY04m1cEjbhIZc4Hs3hXrqJlnzKDW+wLUQJtUEZEuQYeuMnq
Cwe8gTMiHoLIWTrJ6UCGPUYokKBFAR8RIUrqDW/hvJcAxKMjosGM/cAoc03Nf4ZY
nRTiRpW65C4Im8ZW1FcUfx5i4Gtl3qXw+Mrl5Ekvp4aaqcNVXZz4g4YqK9hhN0+P
4pgr/TFR6ujGcyL42t1k9fXkBsRcjTxzpaX7hvJ/3nvlqovAhGRkpzGLAn3JmMyY
oDV8Fp0/MJRVpVSkEy3IDqx5LidqUqmjlhiVKEKJWRCPTYnvbFTjiavF1dzFKEIb
VGbZj3KSyE0X6lj/74CPGNuccswzhU5WtBfTWq6RVWe+Unt1/xFIKKoLIpU76rLf
xuEw+lJ+t7ogYeFovfdQilgezsZd/M2OxZjh64zloGA7IibwQHZni5uXOQrv0U0/
q7ruQ5a6LsfO18bwF4VlBDCxt7pI/uy110vZwBA0KISWskTTzNelnBEyUoRIOmSe
riXhkzG5mQ6l1QzF3seh9WuMMld2JdRXV63UYbnxl949v4M0vKbC26FXunpnxNOF
bE+K/lGgxfPRmy7JQWQTDRGPlMwtpvlniBTQBQlyH2Ra1GksU0Rae/SHZ561Ff2w
Jv7czDJ8Bt6jwqybyM57mP/jUZHpnUFikvx7mkF24yJraOqvzjvgjZ6j4FkAfT9U
83phspAz6kmeVgBj6t7oXq8v3HRFO6wSoByR4fs/dXapc0tgH5PrOa6KD5ahE0Kg
tzeG/l96WPJYpD2U1ziAhtWHVNPi1/1ZXAPelXWghDHWc+r1FSbA6IU3+ZEmzJ4m
9A045V+6UtWsHA/3naZphT5ajKflgiTP8gAvo7g2pPZwLnMQGhIJ2SHX7HZ3qcwF
VsR/my2q4ANTE+1ksjk/q608kpQI/H2pUIAB0FfqphKQFOl7XN7T9ZhcSJXUgbdn
zUTIohuSBfVMhAgK3KUMX6K12SMFC8R9nmf7hw9JW4D0j+f1uVAUmf5XqHWJczCb
nWZsjaGGSzlO/a14eNcYQ/c1Eecm1KAbLRydcdxuKscugKFZD8BhN4FgPEm+3smu
uZvkaQSYE5FAkEDT64GBSBbhWlTFJqM7toyWMrrWZh/8CpCopODWL8m7ww+cpI+h
M1hYcHqwnfRATQFonS+rtPSu08QH/e5PZjR6dt5VwZvsZk9q8tesix76oPheV22l
cIJH6uAi6DroNwDoInIkOjjMrjFsBbX2xyk1PQjWgW+dnWNi8kHlQonYB6Z+tMcS
MyyIGvvoEt3NdJzkyMIMbr9QUAjvTuVcajmbcO2CmICgRQse7kjv5/c1/CfixT4s
cyOitnkUXCSzx5lx4c5EN4FSZlgg4gClQAOEpL381UZMDjKkjgTYm+6R+uioJe43
x8jXvqqqKRpz/ucez4rmwWGCt/+INzZzjWFQ0vZvS+M=
`protect END_PROTECTED
