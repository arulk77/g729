`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMzGribrqanRtM9393uiZltNeYylzGdoNMEfiDPBdWKQ
q/MF++K5V85fgQ7+16PYVT3AVjLlrI0BYx+I6J4YEQF5NXZ2Cz+USVu4nZvMnsmH
Wu7xFoWFk4ODRsiCrC6lnB7zjUvP1GcZOemOFD6NeLXW2KRhK5B9SSZ8DfePzNKB
cLVKLrgkajcD09Ld72zQLmPkFhP5zAjm1dx2sheEJV/JL1w8trfRDjVqYxwmvUKu
`protect END_PROTECTED
