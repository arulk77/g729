`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wvVNAYHyGe8eWIUUri/kAxnyJpSUZNHsJ4xFIlJOADb
Z6CcWIGYCyOLtE3Ji/sCduEeDbbfTt4u4iB8NiycT1enB/bVHlnxjWg+cgZNAX+B
m26yy7SfaDRAP3DVe3wzcd8su2u+vS0ht25HfH2UuINmtBqPqLRCa/0TgfoZ22ZF
GEKLHUK77/QBNtoIsJZ60L5jbjGsneZsD7X44HDBcAvm6wmU7tJP0j53i+lyngNK
bYNXRstuxaD+l9kTkHFDkv1d4JbXHqidVwlfiSapue7UgE/6fuG2LbTQOeBsSv6c
jRws6VoyChaw+c0mVwIlfA==
`protect END_PROTECTED
