`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47Aew8ggTXEA9UAnOvbbUdbfYY22Ps6iuuSMKTh12hJr
nJ0yHS8Bu6xH/3IVN1fBPALnThqjXPUtopPBV/XiHZjWThgKelBPOSra1kaDL0TF
ddcFxabHw//XQ66O6/QQIAV1/oE3igM05QuZJqgQ9VrAb2cMqbVN8ZwgciY5xi8s
CgtPVJA9bdSWTLnAhL9r94z/+3iPJDg26x+BsLca5Z2lBa7V3wT7g2zEzwImzwfS
twCJK4qhNbQx1haL3UtS9N+Hcr0A3iSA2cLzdDq3BhU5954hGraoxHpvJ2tIWeHF
o6LSCt/m0tudArwmKwTMgH5oWycXg1CErMMMqoKSZJbovlVp6hp0WRYkkEPfgEtb
KINeCLH+UhPqL3mjSFO2tcwUbz3d7LVGUXfV0TKKWnKZGfDCqX2LYlyUqnDGWauA
mXfmVR1YgXujVzhtqqVSae2Zpt36U489qPbz1c3bWf4k5NByDN3ef561JCLCxmeN
5pRLp6zP3CRhYDaPzX81w9t7x+cpZV/HmRGNC/ZS3rhsWS1zpZEWQeGC7eS2B7GV
L2qgjafIzErDBB+zguEkK4URkQwSY2q3uS4mHelvWrniWIes1C+mnH6sr/Zqre6Y
`protect END_PROTECTED
