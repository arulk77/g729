`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAiP5NEYZXiwEiopmWDO1ofXu4DwwxZJWctrxMbSE0d8
y3XPjAkLu2P14WQ0uC0LDsxm6iv0uYpZJjRbJdtt0FEBeoHGy8SnIs2eImjjB1bv
G6qgL1kKkW/h0z/zOtb09mBvcOAglTGS8Pnhmf0NOJ6uocGUZYZ0SNX1h33bbOl6
AH7R0ZTtm03q7EjXcD6BB9bTm1eInOsfYALOPM9PbGif3/gu2f9y88ixnVtd92lT
+uDy13k5U6Cm2ZbtZmEAtHw+qfoZJHkZZVb6BEaawAKRA8+dCsC6Egs69Q8zAzCw
OGcVsHtY8FqrxtMh1sFOhJWz4pK6UOW1uaYgCPyuKnMBkik73YUnDbg2lOKLFjqT
hU/e+eI8x1r+FF/KfnLzY2tJTPo4X9nrdXdHfaDJNcS31JEL6YR4adZIxfXdLndM
luWLL1OkSFljaoSj36TpRY3Y+6FGFMQAFjSiRtog25BHArTjeVVJjr9VssWvG0K8
FrJR8kkpLUxbuAHRERaLkrEbI9yRQ0EPh/XLKPrixO6REw9xo9hDfYapPyILU1CN
+Yo8Pb5NlCTQMLQGNACnhjCRrl1VdAcDXyQpkmLQnB9zi4cw45FW27KEfRiRmOrY
`protect END_PROTECTED
