`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SVMgF+8Yx/1Br94BBLBMGJ/Q3yg0WB3pyi/4WL0J3FAc
KIeAYoe58WWgGVxgCkfVHb0xp5E4s+BBXjSKAoSUGoI7bqyYdk9Tp0IXBhgoVBst
OsBH5oG/1HcqFM+lwJZthYEE7xiA1ws1PnMTBJGgZuRQxOwkCMY7C0Ka/t70OcG/
kQy4G3pJLyDa+DKfY/3MH7nvj039TQMvigZBMkTNeneIcRaArHQDSDjv/eG2vllj
a5GnRk0W+paxcVy5MAHku142vtAKcTUY6E3hXO9wfRIIpbt/o4MG5oIol4Wr285G
l8Rh5Q3XETLBXmyAVNyG54+wQyZcOkFHLMKHQ8N2Da4gZnaTsKqBenUkKwAXk5zq
0+vpRPdpUTzjvu9klLB4JC5HgvF1aUuZxl7DseBWIHk0ZBE3V5jtdgu0m7pH/rdA
Uv2Y+DJjBSQ7b7/4chFTircIesDW1dQvlqmiHj3wxd/s/DK9Bf+BCdpAmP3D0Ow/
dcmwS77N8lEFz3TtiLqQqGITdPmPmRTyEZOw8nDrB6ItK03l5t9EPvbP2szF77bZ
iH7MYGVJtZLy1KzoZpRf0e6tjqWcVhOXkK8IGS2JnHs9T3OsLDN9o564DD0xNeat
orJaG5DHmT+zKXsj9m5Um4jnp0+hXvdvYeu+SOUPiwLa/CqGRLYpgb/VfVoiV+Tb
hcF3qJCrTe0OvEqrW1mfkUo3GGd7+QDWiozxY3Ukdi7FVY15OpHz3o/vn8rNERdx
TIJ/hDZ2phshpfhdvo6oD1qmiYgUcGBTFLDDn50Z+fB/zxQouNKwxROsKX6cqe48
8LkDwcn/CP/aco6V6oj8WqIyjZE6cmUykkKKGrhldi4f9LOI3h17VDgTUadYrh6j
JkCfRFF6gF7dD5XP/BtWOzkMtqsTzb7nKQs+vuEBy9J30tf0lIjfh9ZntvZHwcBG
bfd9Pw8kn8whRDe03qrTK+sepRKw28pgI5Wa7DFzybbC71u1Nz+GFbuHIV/sHnXZ
DnukLQSGe1VPhGNwARzXfBVbEKxnDM82tzeHsToklYF5mcZiURTsBvE41cdeIVZm
aQnwoY3bFzjqQ1cVoazOorrgHDiZc4apz5n4ISbhccY=
`protect END_PROTECTED
