`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN4rFOocwvR0cxuQRq24/hqPm5cgBjTYaVw/LkqC/uzf7
nrkkUvqkPjrMNICivvoIPyneN3o9rDo5jJN10wq3m1Xz1XyDSjcur5IXqdN+Vr48
c0K0pMG1UZPck7OtO49o2+zMFNv+pF0C9rytcgR4k7lExpQ5XoXjHRjMqqaZkpSk
B/Ez/odkJNfjvSL6odO9DH9VkKic7Sl+QCmugRFTTwtJ87+Z0yew9ap8OYk1Vgzv
D04j1wzyDIoxNWJLLh8vhPRIvD8q7Sm4xo69Hy+w2yNZBhDUH/JDGofg8Is4FE7V
XAmHl5InGbg99aSPNcOcVCy7gVn3XazfMfUk0IDWWolddCDnLmCIEX+mpZkYvPCm
`protect END_PROTECTED
