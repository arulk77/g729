`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41U6rHKtkFLxwHZm38a/PYm/OOK73AAu/SmP1eMT+Cxg
+oidWCmhaN1inpSXVBuEHKyAE1AfSNcJ1hvNvdrb/lsap8XVH0OfIYJn4O7KSC7G
PqLUQeGqEOlu5G7ZuID0fSvopuQ9qK61oW4oy2SZlxvti/9idq9Gm21sE04+UKvp
WVuW1HFDRTbtsBEx122fUo03bBlk5VKgDVmKq8cySR+StthwnxfsCjkxWLu+HINd
fFozGNz183Kprrhl8RQ+l9VrSs6hiVYalsiiA4nhh+gRGqHucjJOjqMk5KC2pX5o
aEaAbqj/nGwC9CIMuM18tw==
`protect END_PROTECTED
