library verilog;
use verilog.vl_types.all;
entity GTP_DUAL is
    generic(
        AC_CAP_DIS_0    : string  := "TRUE";
        AC_CAP_DIS_1    : string  := "TRUE";
        CHAN_BOND_MODE_0: string  := "OFF";
        CHAN_BOND_MODE_1: string  := "OFF";
        CHAN_BOND_SEQ_2_USE_0: string  := "TRUE";
        CHAN_BOND_SEQ_2_USE_1: string  := "TRUE";
        CLKINDC_B       : string  := "TRUE";
        CLK_CORRECT_USE_0: string  := "TRUE";
        CLK_CORRECT_USE_1: string  := "TRUE";
        CLK_COR_INSERT_IDLE_FLAG_0: string  := "FALSE";
        CLK_COR_INSERT_IDLE_FLAG_1: string  := "FALSE";
        CLK_COR_KEEP_IDLE_0: string  := "FALSE";
        CLK_COR_KEEP_IDLE_1: string  := "FALSE";
        CLK_COR_PRECEDENCE_0: string  := "TRUE";
        CLK_COR_PRECEDENCE_1: string  := "TRUE";
        CLK_COR_SEQ_2_USE_0: string  := "FALSE";
        CLK_COR_SEQ_2_USE_1: string  := "FALSE";
        COMMA_DOUBLE_0  : string  := "FALSE";
        COMMA_DOUBLE_1  : string  := "FALSE";
        DEC_MCOMMA_DETECT_0: string  := "TRUE";
        DEC_MCOMMA_DETECT_1: string  := "TRUE";
        DEC_PCOMMA_DETECT_0: string  := "TRUE";
        DEC_PCOMMA_DETECT_1: string  := "TRUE";
        DEC_VALID_COMMA_ONLY_0: string  := "TRUE";
        DEC_VALID_COMMA_ONLY_1: string  := "TRUE";
        MCOMMA_DETECT_0 : string  := "TRUE";
        MCOMMA_DETECT_1 : string  := "TRUE";
        OVERSAMPLE_MODE : string  := "FALSE";
        PCI_EXPRESS_MODE_0: string  := "TRUE";
        PCI_EXPRESS_MODE_1: string  := "TRUE";
        PCOMMA_DETECT_0 : string  := "TRUE";
        PCOMMA_DETECT_1 : string  := "TRUE";
        PLL_SATA_0      : string  := "FALSE";
        PLL_SATA_1      : string  := "FALSE";
        RCV_TERM_GND_0  : string  := "TRUE";
        RCV_TERM_GND_1  : string  := "TRUE";
        RCV_TERM_MID_0  : string  := "FALSE";
        RCV_TERM_MID_1  : string  := "FALSE";
        RCV_TERM_VTTRX_0: string  := "FALSE";
        RCV_TERM_VTTRX_1: string  := "FALSE";
        RX_BUFFER_USE_0 : string  := "TRUE";
        RX_BUFFER_USE_1 : string  := "TRUE";
        RX_DECODE_SEQ_MATCH_0: string  := "TRUE";
        RX_DECODE_SEQ_MATCH_1: string  := "TRUE";
        RX_LOSS_OF_SYNC_FSM_0: string  := "FALSE";
        RX_LOSS_OF_SYNC_FSM_1: string  := "FALSE";
        RX_SLIDE_MODE_0 : string  := "PCS";
        RX_SLIDE_MODE_1 : string  := "PCS";
        RX_STATUS_FMT_0 : string  := "PCIE";
        RX_STATUS_FMT_1 : string  := "PCIE";
        RX_XCLK_SEL_0   : string  := "RXREC";
        RX_XCLK_SEL_1   : string  := "RXREC";
        SIM_MODE        : string  := "FAST";
        SIM_PLL_PERDIV2 : integer := 400;
        SIM_RECEIVER_DETECT_PASS0: string  := "FALSE";
        SIM_RECEIVER_DETECT_PASS1: string  := "FALSE";
        TERMINATION_OVRD: string  := "FALSE";
        TX_BUFFER_USE_0 : string  := "TRUE";
        TX_BUFFER_USE_1 : string  := "TRUE";
        TX_DIFF_BOOST_0 : string  := "TRUE";
        TX_DIFF_BOOST_1 : string  := "TRUE";
        TX_XCLK_SEL_0   : string  := "TXUSR";
        TX_XCLK_SEL_1   : string  := "TXUSR";
        TRANS_TIME_FROM_P2_0: integer := 60;
        TRANS_TIME_FROM_P2_1: integer := 60;
        TRANS_TIME_NON_P2_0: integer := 25;
        TRANS_TIME_NON_P2_1: integer := 25;
        TRANS_TIME_TO_P2_0: integer := 100;
        TRANS_TIME_TO_P2_1: integer := 100;
        PMA_RX_CFG_0    : integer := 10420361;
        PMA_RX_CFG_1    : integer := 10420361;
        PMA_CDR_SCAN_0  : integer := 113276480;
        PMA_CDR_SCAN_1  : integer := 113276480;
        PCS_COM_CFG     : integer := 23595534;
        OOBDETECT_THRESHOLD_0: integer := 1;
        OOBDETECT_THRESHOLD_1: integer := 1;
        SATA_BURST_VAL_0: integer := 4;
        SATA_BURST_VAL_1: integer := 4;
        SATA_IDLE_VAL_0 : integer := 3;
        SATA_IDLE_VAL_1 : integer := 3;
        PRBS_ERR_THRESHOLD_0: integer := 1;
        PRBS_ERR_THRESHOLD_1: integer := 1;
        CHAN_BOND_SEQ_1_ENABLE_0: integer := 15;
        CHAN_BOND_SEQ_1_ENABLE_1: integer := 15;
        CHAN_BOND_SEQ_2_ENABLE_0: integer := 15;
        CHAN_BOND_SEQ_2_ENABLE_1: integer := 15;
        CLK_COR_SEQ_1_ENABLE_0: integer := 15;
        CLK_COR_SEQ_1_ENABLE_1: integer := 15;
        CLK_COR_SEQ_2_ENABLE_0: integer := 15;
        CLK_COR_SEQ_2_ENABLE_1: integer := 15;
        COM_BURST_VAL_0 : integer := 15;
        COM_BURST_VAL_1 : integer := 15;
        TERMINATION_CTRL: integer := 20;
        TXRX_INVERT_0   : integer := 0;
        TXRX_INVERT_1   : integer := 0;
        CHAN_BOND_SEQ_1_1_0: integer := 74;
        CHAN_BOND_SEQ_1_1_1: integer := 74;
        CHAN_BOND_SEQ_1_2_0: integer := 74;
        CHAN_BOND_SEQ_1_2_1: integer := 74;
        CHAN_BOND_SEQ_1_3_0: integer := 74;
        CHAN_BOND_SEQ_1_3_1: integer := 74;
        CHAN_BOND_SEQ_1_4_0: integer := 444;
        CHAN_BOND_SEQ_1_4_1: integer := 444;
        CHAN_BOND_SEQ_2_1_0: integer := 444;
        CHAN_BOND_SEQ_2_1_1: integer := 444;
        CHAN_BOND_SEQ_2_2_0: integer := 316;
        CHAN_BOND_SEQ_2_2_1: integer := 316;
        CHAN_BOND_SEQ_2_3_0: integer := 316;
        CHAN_BOND_SEQ_2_3_1: integer := 316;
        CHAN_BOND_SEQ_2_4_0: integer := 316;
        CHAN_BOND_SEQ_2_4_1: integer := 316;
        CLK_COR_SEQ_1_1_0: integer := 284;
        CLK_COR_SEQ_1_1_1: integer := 284;
        CLK_COR_SEQ_1_2_0: integer := 0;
        CLK_COR_SEQ_1_2_1: integer := 0;
        CLK_COR_SEQ_1_3_0: integer := 0;
        CLK_COR_SEQ_1_3_1: integer := 0;
        CLK_COR_SEQ_1_4_0: integer := 0;
        CLK_COR_SEQ_1_4_1: integer := 0;
        CLK_COR_SEQ_2_1_0: integer := 0;
        CLK_COR_SEQ_2_1_1: integer := 0;
        CLK_COR_SEQ_2_2_0: integer := 0;
        CLK_COR_SEQ_2_2_1: integer := 0;
        CLK_COR_SEQ_2_3_0: integer := 0;
        CLK_COR_SEQ_2_3_1: integer := 0;
        CLK_COR_SEQ_2_4_0: integer := 0;
        CLK_COR_SEQ_2_4_1: integer := 0;
        COMMA_10B_ENABLE_0: integer := 1023;
        COMMA_10B_ENABLE_1: integer := 1023;
        MCOMMA_10B_VALUE_0: integer := 643;
        MCOMMA_10B_VALUE_1: integer := 643;
        PCOMMA_10B_VALUE_0: integer := 380;
        PCOMMA_10B_VALUE_1: integer := 380;
        ALIGN_COMMA_WORD_0: integer := 1;
        ALIGN_COMMA_WORD_1: integer := 1;
        CHAN_BOND_1_MAX_SKEW_0: integer := 7;
        CHAN_BOND_1_MAX_SKEW_1: integer := 7;
        CHAN_BOND_2_MAX_SKEW_0: integer := 1;
        CHAN_BOND_2_MAX_SKEW_1: integer := 1;
        CHAN_BOND_LEVEL_0: integer := 0;
        CHAN_BOND_LEVEL_1: integer := 0;
        CHAN_BOND_SEQ_LEN_0: integer := 4;
        CHAN_BOND_SEQ_LEN_1: integer := 4;
        CLK25_DIVIDER   : integer := 4;
        CLK_COR_ADJ_LEN_0: integer := 1;
        CLK_COR_ADJ_LEN_1: integer := 1;
        CLK_COR_DET_LEN_0: integer := 1;
        CLK_COR_DET_LEN_1: integer := 1;
        CLK_COR_MAX_LAT_0: integer := 18;
        CLK_COR_MAX_LAT_1: integer := 18;
        CLK_COR_MIN_LAT_0: integer := 16;
        CLK_COR_MIN_LAT_1: integer := 16;
        CLK_COR_REPEAT_WAIT_0: integer := 5;
        CLK_COR_REPEAT_WAIT_1: integer := 5;
        OOB_CLK_DIVIDER : integer := 4;
        PLL_DIVSEL_FB   : integer := 5;
        PLL_DIVSEL_REF  : integer := 2;
        PLL_RXDIVSEL_OUT_0: integer := 1;
        PLL_RXDIVSEL_OUT_1: integer := 1;
        PLL_TXDIVSEL_COMM_OUT: integer := 1;
        PLL_TXDIVSEL_OUT_0: integer := 1;
        PLL_TXDIVSEL_OUT_1: integer := 1;
        RX_LOS_INVALID_INCR_0: integer := 8;
        RX_LOS_INVALID_INCR_1: integer := 8;
        RX_LOS_THRESHOLD_0: integer := 128;
        RX_LOS_THRESHOLD_1: integer := 128;
        SATA_MAX_BURST_0: integer := 7;
        SATA_MAX_BURST_1: integer := 7;
        SATA_MAX_INIT_0 : integer := 22;
        SATA_MAX_INIT_1 : integer := 22;
        SATA_MAX_WAKE_0 : integer := 7;
        SATA_MAX_WAKE_1 : integer := 7;
        SATA_MIN_BURST_0: integer := 4;
        SATA_MIN_BURST_1: integer := 4;
        SATA_MIN_INIT_0 : integer := 12;
        SATA_MIN_INIT_1 : integer := 12;
        SATA_MIN_WAKE_0 : integer := 4;
        SATA_MIN_WAKE_1 : integer := 4;
        SIM_GTPRESET_SPEEDUP: integer := 0;
        TERMINATION_IMP_0: integer := 50;
        TERMINATION_IMP_1: integer := 50;
        TX_SYNC_FILTERB : integer := 1
    );
    port(
        DO              : out    vl_logic_vector(15 downto 0);
        DRDY            : out    vl_logic;
        PHYSTATUS0      : out    vl_logic;
        PHYSTATUS1      : out    vl_logic;
        PLLLKDET        : out    vl_logic;
        REFCLKOUT       : out    vl_logic;
        RESETDONE0      : out    vl_logic;
        RESETDONE1      : out    vl_logic;
        RXBUFSTATUS0    : out    vl_logic_vector(2 downto 0);
        RXBUFSTATUS1    : out    vl_logic_vector(2 downto 0);
        RXBYTEISALIGNED0: out    vl_logic;
        RXBYTEISALIGNED1: out    vl_logic;
        RXBYTEREALIGN0  : out    vl_logic;
        RXBYTEREALIGN1  : out    vl_logic;
        RXCHANBONDSEQ0  : out    vl_logic;
        RXCHANBONDSEQ1  : out    vl_logic;
        RXCHANISALIGNED0: out    vl_logic;
        RXCHANISALIGNED1: out    vl_logic;
        RXCHANREALIGN0  : out    vl_logic;
        RXCHANREALIGN1  : out    vl_logic;
        RXCHARISCOMMA0  : out    vl_logic_vector(1 downto 0);
        RXCHARISCOMMA1  : out    vl_logic_vector(1 downto 0);
        RXCHARISK0      : out    vl_logic_vector(1 downto 0);
        RXCHARISK1      : out    vl_logic_vector(1 downto 0);
        RXCHBONDO0      : out    vl_logic_vector(2 downto 0);
        RXCHBONDO1      : out    vl_logic_vector(2 downto 0);
        RXCLKCORCNT0    : out    vl_logic_vector(2 downto 0);
        RXCLKCORCNT1    : out    vl_logic_vector(2 downto 0);
        RXCOMMADET0     : out    vl_logic;
        RXCOMMADET1     : out    vl_logic;
        RXDATA0         : out    vl_logic_vector(15 downto 0);
        RXDATA1         : out    vl_logic_vector(15 downto 0);
        RXDISPERR0      : out    vl_logic_vector(1 downto 0);
        RXDISPERR1      : out    vl_logic_vector(1 downto 0);
        RXELECIDLE0     : out    vl_logic;
        RXELECIDLE1     : out    vl_logic;
        RXLOSSOFSYNC0   : out    vl_logic_vector(1 downto 0);
        RXLOSSOFSYNC1   : out    vl_logic_vector(1 downto 0);
        RXNOTINTABLE0   : out    vl_logic_vector(1 downto 0);
        RXNOTINTABLE1   : out    vl_logic_vector(1 downto 0);
        RXOVERSAMPLEERR0: out    vl_logic;
        RXOVERSAMPLEERR1: out    vl_logic;
        RXPRBSERR0      : out    vl_logic;
        RXPRBSERR1      : out    vl_logic;
        RXRECCLK0       : out    vl_logic;
        RXRECCLK1       : out    vl_logic;
        RXRUNDISP0      : out    vl_logic_vector(1 downto 0);
        RXRUNDISP1      : out    vl_logic_vector(1 downto 0);
        RXSTATUS0       : out    vl_logic_vector(2 downto 0);
        RXSTATUS1       : out    vl_logic_vector(2 downto 0);
        RXVALID0        : out    vl_logic;
        RXVALID1        : out    vl_logic;
        TXBUFSTATUS0    : out    vl_logic_vector(1 downto 0);
        TXBUFSTATUS1    : out    vl_logic_vector(1 downto 0);
        TXKERR0         : out    vl_logic_vector(1 downto 0);
        TXKERR1         : out    vl_logic_vector(1 downto 0);
        TXN0            : out    vl_logic;
        TXN1            : out    vl_logic;
        TXOUTCLK0       : out    vl_logic;
        TXOUTCLK1       : out    vl_logic;
        TXP0            : out    vl_logic;
        TXP1            : out    vl_logic;
        TXRUNDISP0      : out    vl_logic_vector(1 downto 0);
        TXRUNDISP1      : out    vl_logic_vector(1 downto 0);
        CLKIN           : in     vl_logic;
        DADDR           : in     vl_logic_vector(6 downto 0);
        DCLK            : in     vl_logic;
        DEN             : in     vl_logic;
        DI              : in     vl_logic_vector(15 downto 0);
        DWE             : in     vl_logic;
        GTPRESET        : in     vl_logic;
        GTPTEST         : in     vl_logic_vector(3 downto 0);
        INTDATAWIDTH    : in     vl_logic;
        LOOPBACK0       : in     vl_logic_vector(2 downto 0);
        LOOPBACK1       : in     vl_logic_vector(2 downto 0);
        PLLLKDETEN      : in     vl_logic;
        PLLPOWERDOWN    : in     vl_logic;
        PRBSCNTRESET0   : in     vl_logic;
        PRBSCNTRESET1   : in     vl_logic;
        REFCLKPWRDNB    : in     vl_logic;
        RXBUFRESET0     : in     vl_logic;
        RXBUFRESET1     : in     vl_logic;
        RXCDRRESET0     : in     vl_logic;
        RXCDRRESET1     : in     vl_logic;
        RXCHBONDI0      : in     vl_logic_vector(2 downto 0);
        RXCHBONDI1      : in     vl_logic_vector(2 downto 0);
        RXCOMMADETUSE0  : in     vl_logic;
        RXCOMMADETUSE1  : in     vl_logic;
        RXDATAWIDTH0    : in     vl_logic;
        RXDATAWIDTH1    : in     vl_logic;
        RXDEC8B10BUSE0  : in     vl_logic;
        RXDEC8B10BUSE1  : in     vl_logic;
        RXELECIDLERESET0: in     vl_logic;
        RXELECIDLERESET1: in     vl_logic;
        RXENCHANSYNC0   : in     vl_logic;
        RXENCHANSYNC1   : in     vl_logic;
        RXENELECIDLERESETB: in     vl_logic;
        RXENEQB0        : in     vl_logic;
        RXENEQB1        : in     vl_logic;
        RXENMCOMMAALIGN0: in     vl_logic;
        RXENMCOMMAALIGN1: in     vl_logic;
        RXENPCOMMAALIGN0: in     vl_logic;
        RXENPCOMMAALIGN1: in     vl_logic;
        RXENPRBSTST0    : in     vl_logic_vector(1 downto 0);
        RXENPRBSTST1    : in     vl_logic_vector(1 downto 0);
        RXENSAMPLEALIGN0: in     vl_logic;
        RXENSAMPLEALIGN1: in     vl_logic;
        RXEQMIX0        : in     vl_logic_vector(1 downto 0);
        RXEQMIX1        : in     vl_logic_vector(1 downto 0);
        RXEQPOLE0       : in     vl_logic_vector(3 downto 0);
        RXEQPOLE1       : in     vl_logic_vector(3 downto 0);
        RXN0            : in     vl_logic;
        RXN1            : in     vl_logic;
        RXP0            : in     vl_logic;
        RXP1            : in     vl_logic;
        RXPMASETPHASE0  : in     vl_logic;
        RXPMASETPHASE1  : in     vl_logic;
        RXPOLARITY0     : in     vl_logic;
        RXPOLARITY1     : in     vl_logic;
        RXPOWERDOWN0    : in     vl_logic_vector(1 downto 0);
        RXPOWERDOWN1    : in     vl_logic_vector(1 downto 0);
        RXRESET0        : in     vl_logic;
        RXRESET1        : in     vl_logic;
        RXSLIDE0        : in     vl_logic;
        RXSLIDE1        : in     vl_logic;
        RXUSRCLK0       : in     vl_logic;
        RXUSRCLK1       : in     vl_logic;
        RXUSRCLK20      : in     vl_logic;
        RXUSRCLK21      : in     vl_logic;
        TXBUFDIFFCTRL0  : in     vl_logic_vector(2 downto 0);
        TXBUFDIFFCTRL1  : in     vl_logic_vector(2 downto 0);
        TXBYPASS8B10B0  : in     vl_logic_vector(1 downto 0);
        TXBYPASS8B10B1  : in     vl_logic_vector(1 downto 0);
        TXCHARDISPMODE0 : in     vl_logic_vector(1 downto 0);
        TXCHARDISPMODE1 : in     vl_logic_vector(1 downto 0);
        TXCHARDISPVAL0  : in     vl_logic_vector(1 downto 0);
        TXCHARDISPVAL1  : in     vl_logic_vector(1 downto 0);
        TXCHARISK0      : in     vl_logic_vector(1 downto 0);
        TXCHARISK1      : in     vl_logic_vector(1 downto 0);
        TXCOMSTART0     : in     vl_logic;
        TXCOMSTART1     : in     vl_logic;
        TXCOMTYPE0      : in     vl_logic;
        TXCOMTYPE1      : in     vl_logic;
        TXDATA0         : in     vl_logic_vector(15 downto 0);
        TXDATA1         : in     vl_logic_vector(15 downto 0);
        TXDATAWIDTH0    : in     vl_logic;
        TXDATAWIDTH1    : in     vl_logic;
        TXDETECTRX0     : in     vl_logic;
        TXDETECTRX1     : in     vl_logic;
        TXDIFFCTRL0     : in     vl_logic_vector(2 downto 0);
        TXDIFFCTRL1     : in     vl_logic_vector(2 downto 0);
        TXELECIDLE0     : in     vl_logic;
        TXELECIDLE1     : in     vl_logic;
        TXENC8B10BUSE0  : in     vl_logic;
        TXENC8B10BUSE1  : in     vl_logic;
        TXENPMAPHASEALIGN: in     vl_logic;
        TXENPRBSTST0    : in     vl_logic_vector(1 downto 0);
        TXENPRBSTST1    : in     vl_logic_vector(1 downto 0);
        TXINHIBIT0      : in     vl_logic;
        TXINHIBIT1      : in     vl_logic;
        TXPMASETPHASE   : in     vl_logic;
        TXPOLARITY0     : in     vl_logic;
        TXPOLARITY1     : in     vl_logic;
        TXPOWERDOWN0    : in     vl_logic_vector(1 downto 0);
        TXPOWERDOWN1    : in     vl_logic_vector(1 downto 0);
        TXPREEMPHASIS0  : in     vl_logic_vector(2 downto 0);
        TXPREEMPHASIS1  : in     vl_logic_vector(2 downto 0);
        TXRESET0        : in     vl_logic;
        TXRESET1        : in     vl_logic;
        TXUSRCLK0       : in     vl_logic;
        TXUSRCLK1       : in     vl_logic;
        TXUSRCLK20      : in     vl_logic;
        TXUSRCLK21      : in     vl_logic
    );
end GTP_DUAL;
