`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF1C8q/ZDW14b83bZZ+WaUDgEadVUPMgqtPPl5APWbk6
X4Pmp73/GWUZdHgXbpSUrNdcanVaJjLDBZmFd/xtpgBZRwXZ4nYLBXNVzFPK8XQ4
kA4FBsJJXjIW/fxub/oNwiYUpnGV++uTWewGlO5H7yk+nIchH1v05bb1sA/zV/ET
CsVnPKjgOD1MiA3GvF4sInNOAaHu2+JxT49a+fjqyghDxX4TqAfAa+Xm0Ux0Lm11
q2yqWf2DLfWdkCfrhOTsOB/OcmRbi82kqcA2W007B3XFR2zHAAkRjnURUmaXQsAC
QH+4rafHu/jdeZW2+uF+fgG5R5NzFETwBV547BR3FC7ddKmDJ2d7XaoQEyibwQbD
vabys7AG7gqMpCXl0w9rUg==
`protect END_PROTECTED
