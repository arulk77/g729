`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
AlGTupyDt0c9gPnMfI9dfWu9IlmawNe1KT4wvPoxbCW3KlqUwVqP5mIXqnLZhW0F
AA9zFlC4aMNDwMiCZsA8yVKVtHGCKRBvNqxwUbx3VBJ4VJ6U5/KHWj4/e9BGq9aw
e5Ps86vLzXHAaRZD0tSB7qg7NbMA+XKwACUzEP49+WB4RYhZxO++fW1Bl+cl6rOG
nIJMuxJou0hVCL8IqnOwJbjaNHbnBhGX3hln+7m1oBsPUWa78SmoQ0roySzbpBqy
0vw8mRxq+UfS57YoBin+Ts7ui1uZDBATYzRxerG0Q/AQn469CqwOIAH+uUxyH0M4
MQJCfxQa5byNJxgD5vFbsTCWAN9BIgkuAS92EBztdh0=
`protect END_PROTECTED
