`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
whfZdEhQhIVICrvn0VMg7jIoTgWyi78P68I30k/sR5D1jflmGWgyIboOlQZV+ee6
s/3gnMHF7il3Pd3SUQAyR0j93OSJl2KXDAn+eTkRn1vFrIaqBzcu5qPGOZ1/2lAL
jxazYaqXPVrKp9M2zhR5eq4zjl3Jzl9BQUCPSEzpPhV7v01r1X1lyu29ZAD0IZk6
PZTbTiITQz0sU7HIr2A67yLB8hvxcu8wOoR6E2VleuhPjEpmt3G9uC+IQElB8GaY
N/eeQjC0sUNz5/DWLEuxGcdtknePLRHbP1f6YpnC6ww/nEDZqG6hOS18qXgknVn1
Y5bZul5mbMBoSzO/Ow7KCDrPNSJVaLonnEJ85SE6Op0LDa3rx1U1Dv5rk0WCP4Po
`protect END_PROTECTED
