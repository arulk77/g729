`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46ZF0E+NKFEUtM8vhlfYIkBz4hUkuAYuypJjq16OkGyo
raK50kGHR4Nd7bQKTQ1klBn4moIegL5MvfhKVMX//irqvT+51DUKJUBpTvWcFOCB
HXp6P8RZIIygeuMmDyQ/N/04K66VoPNSykp/rF3a3BfpHKxGmR/Y6DuEqtGuidqQ
L9gyMIPrnu3My6vdxQ7w0SsCUXNA44h9C0bNG4ZXPDyie6kKBzrNS15eaEBi7mMR
HX1hGNgKKRs7Sbvxh6ABMvWakDWar2oma4M6Zl7nznFJmdnQR32dKWQxfI79MGtF
n87/Def0Xllw5kDiwD9zmbJXheJ/4UhzrSKVDdMReHKmiY6QuRDBQx8dZbOAkrKt
g4kbw5Q208eJBdN/JU5vqA==
`protect END_PROTECTED
