`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4z8f5zyvx+eW0svewf5eVNx2GvbjkfJnaKNIvoK5575R
pNkvEvlXJx00lJOcEqBv6A7XTV+mD48Kjr2wf0W3R2zQ+Pxypwyjst2jxep//Hbg
BMdefp1ttyt7DPVuGCUOKUVwq9TNnnkwLuETOSHqbLStChQWRkF/DQlRQaSmJGS3
ci50gLg+l8xsRQUZ9yPg2BnHxuyEJUTUcJOuyNCqQXhWoTJKKJqUj+6WxlsONvQN
amCnRnPxmobZPXtdtrvyuchryVQxUOeBKOSE9/6+B4yHqekzkpb7JVxxslFYClky
JWw0kSuKxVFahd7j22SWKQ==
`protect END_PROTECTED
