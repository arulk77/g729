`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJBZmOFPChaeHco2/sDBKUtCsUBY4tCLQ4LJfi4Gv3BT
CMbKtUoALAMR86xsWBe2I8FbSYRD0IRWv0oMYeW1h73oFqpwpkflRPlYMW7FirhO
pD0M4lHQlKrEACn8Qcq+xvY2iucHhNYmsSrrcFEnVIdW8AS+NbbZ9iCYu48/pZ4V
KZsmVcbV+WVFWoTNYsnh1IFGwkM9zr/9cRt8Yh+s+T97iGZAO+bYwSEh6Rwy6JzG
wayxnkFsVZmG0ow+5BoC0Lmp+EP2Awn+8Dn+PNDgN1dXqs+JJGMuT2h8SqrXBCHO
V+tOsd43w+IB67vsqFC71Z9HZpk0h4UcHsSbB+U90dNKOpHnwV2n4Y8fCK7ZkcP1
V3AbT4leT/Gk9F1/7oeEfb9FH2A1L68h2aScWkftGsgQnnZOI3YcpKLrGDCqnpkQ
Fm3TAJwXPjZXNdpGapXNS70osO2Nh31Z3w1shLVn4Ia+962qhg97CuG5Y7pffBVR
p6riE0YYVIm2Ad3IvEFVX9IhnSKxw9j9108mmQdTRYbdBorY6wSz/DiRdni8mkGU
`protect END_PROTECTED
