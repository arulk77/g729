`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
u2UyqOYzRsg93uSsEjvgAT1+RhmPOkojkvqq0GfZmAzCYZQG/t+8sUxCHNVqPONI
BI+f1WiMPq9T2J0YELlFgjkp+iyU0O8XUsqc6rBhZQeVWErYROM6579qFe+5maJC
PuVJ8xZjzU4Bvh2Gql0UOI/+TpXJ1kbXufAXProYFXln0qXixOaxiQOs9UYa1rur
UeEunZ0L7taTEAEU2NJZSkQYPEdX5TscS/dOb76LxIYWUX2ChxEjf3PstpbPgfbM
`protect END_PROTECTED
