`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNVKQjEupR+//GSJcY22p0CP5nyyLO0OLV1KcRn5BZXm
f7Pm+yjlyZCln1lZD2UvVqm/sjjKsYnboWtVrH7GZDef1cdhuMfv+Umu3T2HOpKR
ULn+eSN7TuUccPWj0E1NmxxP2Q6OGPz7tvk/DRodaUsDf9W1O0z+tsxXmBED+pGJ
2wE3992L8jn/oDAQ8T7sLmVPxlcoZhjghMxjEvE0+LlaNgducn44cIwgHOnLOpPA
3NZiy2FnZQhvrpehyRDZbnZdkdsTb7lOSiLXDYJmnCbkdy5b0Ay6p2bLP+lK8pmX
oGmBiJc01ngzgvnTNSDJSQ4cr9uUMGLo4dRwSZK4liotKsQFt3ZyLifxbaEhsR+6
hDmpOXghlfCn6Uu8uibPP62nUZFLyVYkS3Or+hsyJkogVJ6hRvNZq2b5SkB1YppR
VoTqa1qkxWsSPClIiEk1sscNI8QTsKux9H0W3LPPin0HZ8de+tbk/RtMPLxdAQln
`protect END_PROTECTED
