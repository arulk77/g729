`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
iCUpN7xiUHFIidYhDqzksZiKVolq4RCXSwWLB+jh/iY2Ro0Y+39fqwwDtguixKW6
/jllY1qaCWwIH90EuOv/5XCORg8jBljmBIS0p66UZdK9dQ04IU6SpfdDX+T8OkI4
ZbKi/rVvT0Ni1ISxcwqxXg/7H9CWpp4dOS2tmqyUv4VbgGf0TJhFZFiOLaZFKYj8
0v8xtjawVpTzie1mAE5Qqt6FO4nds0BW00iLc8DufYU+Vp55u0hZSpmZGipWFGLb
TL2eE6BL9+R+awzBHelQ9Di00ejwgDpFzk9PLujqRVjVJOtAjb1SFr/5DlRWEjT6
yyoHmv9mycTKR09XNtEMN/pqfQXtBiRWD4kpoeqpWt4=
`protect END_PROTECTED
