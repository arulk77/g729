`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aZ7GtscqD7vBfzs93U0lfxWmwSnh08zWQ5zVN0hjyHXt
7VbfA/PAY1fPwnkjJSpYQ/X5aurnesRxqAx/BbTYd1Qs29flCXzd9khagxSjNiuY
+vJVAeQncCoD7bwsC2Q2+3bmdFW1QgglxZ8atwI9FJ1/HJZioShXHnu5bt2fNDW8
BmVK9qG2JoJI8h0mza80vyL+oClkwbq7RXNH4Kp0T7Tmmygs/O+xE9/5ebD72nwI
P+NyurH+C1XqjtMq+xSOny/sZeww3ZzDDCwHO4NZb9/6mgmeOhJM6DqiH6MQoAEO
QCrRaBebMozg74BZA5Hzc9vm2NIcuIE6/uPnUEj1FAgEvANsrRtLcTrwow7giK4K
heg8G4/d241jFuNr7mBcRRei3kMAPK7vo06vA1NE76rrOVvqHVCejF8QJFSWDouO
t76usQk1p+GK9u8+ZtwyIcVU0VKEcNwtHFVi4hOAK9uks6mSPvo8TaGu+wbX0bmr
R1ByJRpwt1gtuT2uFetrK0iUuiRusP0XFp47dGgXFDFnyiOtyL8w6JEuD3vvuM2m
KAWoUXpv+1IzCNYU1/bWan09cD6JWILHXITjmgkxNGTteRajnV3ibuBgaPo6zdFw
R9cNRO0kZ9i+q7e/RP0O6+dE4zWIGfX8/pDyAzvN6DRLUhO5t++7vKyQCtppVkxM
IAPvu4zNuGrIk5z3eKAv2i/vJlGX2EVrJYl/HALT7WFS+SAxxUYd77HXVmx4dNeA
LTIzoZdVqUlzFtc6pjgnIUSXmAB/k4txfCwvK1BW6ZM4NuQcXdc9eTujKTTJzz42
Kr8wbLczI9TFkghDA9edit8554EA+OBAUrf7mzyK4+zeW/p1a63tLReKS20OV/zq
vi8UudSodtDP9gXB/6qqY+hi/xHV4NbEwpdxwdTdfUSV7rajPN65G84UmraUK6KJ
`protect END_PROTECTED
