`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkQlZFLXQkfoSodCbc0XGklmw5CtKSKrf23ASKswbAZnO
WO15PCmCrwVoe9yTQFQV55Ui2c8lJRpRDoB07gA/2ZmL5d+Ce1oFsLqxotocc6T2
SCkrTdzTXLHUKZcx/wtXSG68taGex1ASvJR+WTKQunboCIem/M+1Ugkv8VoiMqpq
oOnHG3X9ZD4kPmW4u2peVSNFCOiEMAqdKfQsLuOas5VE/T18Efj//PmdigTZ/CKT
335dRoSn9KlikriyYLaAdoFysPz4wKwI66xomijNdx/BjUN1/Zh9jYTLGpKOUNpt
F9czbUI5JvpmqJ118VerTUOe4hMTGkN5qwKO9kLL8ZIjVrSJDEr3dv+koG1K62e5
3GMAU5VFFrUpAs0fSwxttP1XDx7raEchDk2kYb3STK9MbP+mI5zohdCY3SXj0G5+
hI/N7gz76z+DcFch2xBztO8lxmenLPfovNmC7ZZH3yii8mIVyIoMrnNlkruZJCXv
J+eRC+I4HUtHNkGF4ByTo5xNwnWOdsySQc8laOwbCIrV//7rNgivAFL8DltyJodM
Y1q+/RzBT4C/n1en9QJrGlauzHQnUmi0Y1ZsGiW4q3JnDYOzhLno6cO+vZK8eJ9+
odzYCV62/FvfEfRKdDMG1Nx8WC8dEw2kjT0ZDU7z6zRA4gXdnSoBv3bKp78WwzOH
QXCHmcM/2VmVzn2ee2cypvO81YLQjV3XeqrJ+etw/c065bA1ACsgALncxZZtfDMI
oOdFisJiucIf0wKStn3yvC3OHld3BFPKls1+ifFHGlBtlExhibEcbbLpEexmhsDV
doAt7+LM5ocXXdByAA4JJhc1bzR31tKfGhdTboSu94YIZqpRdqoQ+d8r31TxUwhJ
Xs0Uvvimhd9Iq+VYxdpAMlnac9RMgnr7LlTLuKU440kqGoDNWkgf6iLW9f/h2QoI
/XHJQYPSJFSnYw7t0+f/aDOuylyzX7Vp4LUEqwDRflPE1h/wIQZw3p1AhsLODpwJ
xwGweHfmnA/CcoMKNRbV9YEhippBRMnKMJG9UJxBx0PzLfFDWyYGnQM2AMcK3YIt
oQupFklBieyfovzIikJUENNS//v66/TIIz7ccqxVvhD6bkZkkNgHd0PW40AEqhPj
cEWHTgcCAk5hGhY07Gq6a7c3/DT48X4DKGtauSp7FCunEoDrd9cf11TepQsus7Xv
`protect END_PROTECTED
