`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHXVl2yCjZoVM/whSajbY1I/u1mYRf4G+ghtN8yk2nG8
FRMvTMoxitl7k/x6qxokYaSZg3+UbHnC/z4OmLwon/7MZAfV10RVnfxA9SzAcFCF
GwIYqQtskuqYZy/QfsO6IFTiGppQaQkyp1nT6D+Qvpb3yplSH964P5zrr1wKusqW
Oj2BICOygs92iiqvrg0AiagDNOicPbViI3ywN0vXmCJr0RIPkFjB2iyMgq4rr0xK
t+nWx21KC6zgfkVaQYbrslGjUeiRzx1Ni4dYFo28zKgnfI1i2905a+Ne7vagq0KW
ayT0sxIw5+f8xc55ILba8kVvlw4xzjMHh0J3D+F0zW3dFzrAz8fdwWpW2ChkVcKR
qWysOT2cjWHxlwdil1cddbPP1pM3WUH0Frh2xHr2ojgNC+L/+U3xhhpb3qmE6nxT
+jkuPXf8UX+n+31gfks9rw==
`protect END_PROTECTED
