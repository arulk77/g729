`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveA0kUISzsPQsJfjrKMleSMTRANeu4mmLMN5CZDqM9alO
U+u/l6LMd8r8hRrnuMBAmiAqY50UxAM1Q1tTwFZ0jgPAh1rspD4MwV9eEbjNSQdy
KkVK4lwlI7S4Xyg6+RR8oUepiYA70SO9LtglxH4dGG/WQG+kH8dgzyHgzw14t6Uj
d+g9vpUMDkyInLEYKykCy3A2VKWax0ta0/1N/gaOTRm0ms+di+sAiiAqEtpMUNBm
z1Vt4Ysy1pgi6TM2eWZj+67ZD0L5+K45n5qmqBUkQOOMOBjiHXHQH2hMidvWQ0nu
K/v0HKgi0PnRP4cTKSmyuUhF7Wz68iqlk5Y5TZBLriPksosrGjIS2RscsnzOEQZl
Qk/0buWrzwjrmma8mYn4VK7sLDQLgZUOWN1wCc8DW3GDrGtUd1L+y3J9AWvBu3bw
bViEy8feU6NteW4tKhC4TBRKypx5fx452swxYQwh9oAzD0BYSZW8mA7xsIednIMD
uP3SLSjhMaUwzJe0M0eOPPVRZj8d7KB5mhbDVYuhu0LyOOVc2OCDogr1lwz3EpoE
`protect END_PROTECTED
