`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN0qK1ibjt+RKgcCTuAQm9as+E8lybQPYHYAmnw+ByY0a
PJiPkD6yfrd/xnlTklPGDdQY4VypJizc0KuO+xjze7yBhFCsU9qKeK6kosg8GUXO
fnEAiNxxy9e3OzE1w+ksyRVTImKM1Av28E7ritS0MlNUxSjACz2c/Uc07HuIq3fM
Ul4O18UnIx87biyVb0lod0eFw4TgQ+L0LtW8GxrVUi/yZeOay+0i95Gu0aK2hFef
GnTK84lxIqXPJtvJXdVxfkPb6m8FD6Qxv5amUwQoXhPeJIR9NO3EB2YocShafDfm
KB0h2iQp/LkeSrxiLA2izQkNLBUjVigFVlUWBe9N90R/ysyZP0Dk5i/ofNaHC6KN
ZHIf+9/A/8H5jPci44JVut+vObIXMvbBUV1g4HalfiSFJtbN8Q/63fUQBQFzost5
2f+JauTTaXSd0kHpz8CB9qVxw9Q63x48gkb3MplqhYahD8QemaOvYz6GWYm1ZBF5
HKu0Wm8eAkdaRhlzGa83P52KAfB57ZTgFAZuwPUofAaIlhZCs5MaMxJtl8kC7nCX
R4TudJ2nHYEfkYGxhlPvTxjetruw3tD1hepHHf7nG99nCZ3gQ3IBl1Mes0YcFdmZ
w373VOAr7t3nyNIdG+Ps9hzh+CtPuhDH33fRsYsXSNKChO2Tj64C/Onkh25ywU5D
3wNVLks/qt0o18rg1OGmSYx757rGwc8RETcfll9O/fW77YoRwPtvItFb4I8qmMkc
v3rUfOORTRItUTLCl0IgGA+Tqm2V3nxDEf1cV0e4vLx7Qa3gnO6JB7EUH5ed8qaH
qbBTaZDS6rtqK3YqMqEjiwzFNJvIB0rq6HVAoRSQOPMZTUJd+o3oS1bFNX5jhxbJ
qoWbgFlZc+aNfhF16hzdpvE1ll/8u5hTNb3OJahGVlYRbjZTMHH+5vEjnW4a2Bpk
8NtwZ3SWw82wq1ADcy3QM07bVpLviy/Tb0yY3s6n+c62OHHlMI6ZtW8Fd9OXRwDH
RCZBiMUZZn+tVVLkqCP028aoy/XdgalxhRbwHKm2yd6aKo6ChOYnMcLch8Ks60xo
AS7xdl20m8SzsdUk3Q+a6bE7f2Uu4mKehv4QuaBgFOUikbuExdwxBnP7ekO4IabI
fMZT130orN5KtAOdif7yh/ukv9B/81Sg4Sw98/rYlv64ntevJA1mUg/pxsyTWj0A
7ICAfDKfgWOTPujTISp6MiesBrfYWvbTEm+F+MGtsLkdIpI5byanLxinTkNyIgIB
Sxsj5xYhuKPs6A4q2kRW1SAEKswAy3S+ZGO90upZqA/qvp31WpDY3BoG2yX3rGAM
R+y7/nMUq2z5BNWmmpHZBZDRmeAjIOMRrTEKc1/C+iCbcGlPzZ9Xy2WKjEs2nOyG
lFC//oYRqyf8q4uhQfaFlu2KMrzj76oRHIvBgCSDzdIerRxIqTqZB2yafwR2Gc9I
xqIE16VzezBFKpUS7OkC84ggpJ0gIxxAfCpmK8nR6J4OHdwhMxNoHUjrqkVB+jsa
puxCdm5+gJg0Dgl+VfmLzemmoqzhc/ja3rf5sqAUnUFmOXhFBrDBUMkW8gUhUVgP
wc7NW1bu1mC+IocjugaiDHYCCM3VmpWG+uPI9pcM3D4WlsiaZnURJwKebx48OaHB
XeKgKtCu9RwYGrsmQP7iNxiEDJKbrvQw4ep3ilCiRiBHPf/XsCD9LUFM7XrF6tT5
NUfPPwEAqDjuQTGHwTXy8Q+vmSEnwFyJI0N6hkpUN7JfpJTyVA7XXb75vfPB6ALD
SorEj4um5zBi9uniFBUg/NJSGdX2EMnrkcMXjXWHCFdW04iVvW8DhuUrxfHENJ7X
VsvgQ93qCEO59lcmU9qkQSlOvEIk9Ido1knZkUDoynbVtmjfxwXyr7VFlPqCwfxP
lR5MhRFGgTclP4D9L++rh3r9g+dor+HPPXFWii/C4RFH2sPDX1l//AFOOdcpUD2i
8WEIrjfKu5CXZ8FBUd+kIWzuwG1QYy5V4LAou96MUQN3bO7oM0wVBA+P8WYD3MmE
aTRu1F82QDzQM5tPIEB/hB4hBM1nD9QL9VOT0uz0fJMW2VXo1dUOuTYi89bfJMv8
lw7I9Zr90SBqmt9t8F4kk/f2zqcWvb0VOyBKGNb/6i+bNU9PhZomX6d9Rchv9B65
C0QnquseZpbULAWlaj0mKLQxvw6k6AZt3VO6tzu+aN52OOF6LHzoULQtd3nIaYw0
F8CVMZhVCli+S1mQHdLmjmb3bQG81IRFQXTwpblnRokFFtp2tAR6fWLveaBQRQGJ
8vd8UnhFcfUuTx1SHT5kJHJpusmn4QL/6EpATUr7ZgiNRvY1E46qxYVlmh9lXAfG
m9T7HkImFmBMzFXU0bfCqx8lOi0XA76Lf+5RWCGrtCQ1T3IJI/jyNe2TAg67gUlU
nPhlTjy7fhHN8u7Zz2obeVjtuNasDtMnpaJMK72/3shkUiXwFbjfdFGf9xt287pF
LpmHh4eWGlgl5dlAWKtGxJPFUplXMjxKyitvRXGGlcaMu420USmO6iZ5tFp9G63K
8E+I1yEbRJN8v/Pyo6qK3Ns0hoo8AtjeRzXMP/BP0/wr4gOCLHRKICyYvgg0J1xN
KAIlKBeA1yAFHXMu5Oxyd3elsxmuUh12imrkvWoGnOJdI+KL1Go790f/vTcSMf1A
5w4mUsuzbedGAnzUV9oYagkPNGzJyDSRCzTHWk/rgFB7I9TZesXf3ielx03TG4yM
zflYHP1UGwBz/NfZj+4gCjFpjrD/TaIMPkc7idVNEcIJGK6D0KBKsQ0Ar7DpGXq3
7oGX1mNnNDevkb0OztbHBec3lN68Z/O2JX8NbvFg/bhdqsderbBHpGUjpvaA0QZq
q2L3eXk8Fm1WPWdBlvYJerWEsBbEILirpc7PTORgmHCqOBWUZoEJtA+2aEbbDnsJ
e5CYkNoEUHwXYQlmluP3Pj9Nfw6vKR/s1soJuvERsCItebcg+AuySpVtg+b1TlDn
nDs7kFUMtbKO+tDnQ4BKuxd8GVoG+8qCPdoqYb8TRL3lDZ1Y6JO8wBJXSPBbO1SZ
heocikatNh36HLyyDZuZ0Q7EjlGlkm7Bw10lA6nJojY4Q3/RHg/FKQqZy7TDOo0R
PgYujMT4qF539nEm+B6z8abk9bDvc5dV4FzMVWXcEE2CRwr9LpsVQLB5Kl2UX+wX
OOHB8x0/zOSwpAqRbI6IE4JK6dX5cuddEW4z9p+LwXGPb7O/Mv/1cwKqj/n4E9Xa
s9LYB15m5rgOZ6vx3gOdyA5WbA7R4CVQQ6/9f7jEsKIWLQ21husAapsqk0t3dzWJ
GBNLF8veQMd8RhoWFKVwj6wf7ceotl4zey/cclEXRVI4o0KX/ma5WMB9lwsR3YH0
NPggVicnTADDD5r9pblUVMB+fkzBOhysM7Q+woxukIix/ZCZfLa0TV7pkZ5Ae3qJ
/R8dZWbH6OBHMy3Tps5sqkSwY6ZlYoKRqMlFZokVVNUMWj4QKoxWabLDGnBbMTQ0
LsDOSEnPBsEoBsn4RhLKSkq9gcUK5GHk3YFzVzP6z15kMzDn+sZv4X4Cf7le3rr0
BOBHlMhP7piJcyS6bDkg5ZKHiFtCXn3dy06Tr6O7mOKCNFNoWxpZUKvFKcVN0zgP
Rw87mz0G6MTQhpynzRvOysBkW023zF/yZIhUuK3thnrXEtxbcRmpZrcj31EpDi1D
uEIS6DX1C3vvk9ADYauGORW0gzIFgEze73tmf3rVyoYYIbgwxVE5JGIEp/SE/kYs
vP3OEh9kra+uf3PgUR+yzsc8HYhUJjqkC4vt2GJL2bcjJIwfb7EInYGon/dko99u
RgXaZnNUfxQLF22tg43cjRwuZw6CMQTmv5fi69P3gG31D5lbY6/6x2cvoGLKwweC
ZjKUiymMjp1uj8q5A/OHqJrMUoUcFp6FiX+V15S91BdTFY9/UafzjOmNxs7hlMhX
xJwUR6hNsBd+wY5gCUvRI5e2DJbieXRYQ9rpLLolKaXWnMVj/FIpe99vNRVNFVX9
MI7F2/vvY3hi9jXWH/E7V0G2v/APGv7gWSH7G8d4I3OMaWj7lCIfowAS8+asVRMY
fQ/uVOTR0qsKCCcXo7+fB88PnAX7VramOvMy7/szaTwZ/gkGBj3/C91/2QfHxFx8
sAiiqjJFsPii/q5rHmuy8pdgguClVmzoSGSpsr49Yq5Ysz8V4S9NX/ajAC/CQY+x
YoIFOZxyDFd59LXwpTWcOzkft9CUxhUQ21KOf4Q1S9Ftt2o2HcE40BD4vcRcgrlT
oW3vAyQ5hOtCRb+h0DgOiJsHn8VHVsLeTWYYLHhlAeGTS8zohfAjMMBxzpHmHUZa
u6u7dBNgWCS4GbKu6vVsdHHx26wWJzlkhr+ZYxXt6+zoVtKCkqumHG6LxQPEZkvw
PsOH+0zmhchN2Ov2V4VjaynE1W9aM2vfSy0hSvUP7OytBFqCvFon0vZ3QphFRl4S
Zhd/0+vgU9o6FXaH1nog+i7p35JM/3OWe+K6O+zcGXFjKchWKb6J4UUxJJcAAJpg
Hkxc+Cj7+uxOtdSuMUsVAjmZRL7YM4HFVvbq8vAdfNe0UZIZlMk3ysJ8+j/au/LU
mNmBC1F0327ZxAoUQgp3HXfZGDfpdQq+nx5R9g8qHRA4Hsjt6SxXglbeHur4pQbC
SJl9CbQIY7WICu6b87h4Ugo+L9XW/BQIBU04UOUH0ry+FAxb8E5uel5FAISlG+C1
z3Qv17L0RGfdobYHXFSEuarSY+SXf/Eaf6tPx3z0ZsTyFcNdr/sZy4moD7U+6HVG
ja+4CJAz0tPrK3oyxKRIFWWQNGKvl/68l2aohi4TTWwCcd0vFRKacWxLpTHbcrRS
aIsMsBqBpvS9T4wSLfASouDOpa9JcrtpwaxovkXBpwWuM6isauPH5D1/IJTuzYMq
6jqFfMoLBsLhRAqO7BpyPAR0WlGyVBZvTKi0UadxvV7p0SkwA6K0gHFSe2mac9QW
jJ/9f3LBVf2ti+4IZGnmZ4y0TqrE7enZUDaj30w/Qd4kGFHwwrn7V9X9kdEGbSuI
kcJXDCmrpNR77VcsQ/P/E+UVSwqipRqWdeEXD1e5S5io4fvqaSOLfrLHNrM6MjDF
Q2m9Alo7XN0OjHPDSeQ9pqHSU45YLJfm9kY4ikIpxDfr8hbHnbPbYjlF5H0Ibfav
ycJUvrUorJ3hc5qYoimryHb++LPujEXLJ7ByvS8p9Y9CSQXNtieEdcY3SX+wAMrX
R1AwybAOLzc+5GhlXkYLduvlMwYMj3F7Lj3pRTGZov7fA+IMvXJHLdO9gcellKFb
0WfD/gYL+2dEWvGRoIeYYUDvwCP7P1od5WDyDiCeElFjlrDx3rHQ/5y4+vSepnei
q/w1BBlFZUq3dLBdwbAujPjTd6t5HiDiatbPKLYWkZ6QrgLLXTwryhumCGiMVvM5
aSVxYj8vtBHoO1r5gVti6ak8muTA/zhMiuUoCyPFo1+kXuic8ugcH20E7npP9AYh
2xKqEMqDRwL+XEPihRZIlcYigdHxq35qhXRltNSzCe6QajKR4NTeMqPUISG6Dc7H
u5Jd4iyaZGPHQ06TKzhqsArFPrXIJQYV/97o6VKzucGCCWE8CZND6wToVIlHt+hQ
vBhuuWiaTfUorbnDlmVrwkerdFXNk9AapVNI/W1ZVRMdbRU+LaNbo2mvBQ+WIqYk
LE7JRqIwRbZiLULvbHYxX2je8o5JjkhlbpLV4Ze3B/kf1pqwgq19UTjTUPbtVynA
UM5QefFUeJ6YzK5Woxl9aRyeX4lAE9kmHPyIn0wwIWVxYSLUOk3qa6KY/eNOA48B
eLx60J6Zl0deCifUhVGenWW/+LjN0p7aB47R7uz3cyPaSwXyKA0csFF8fdNhYCKi
9CkfgXKXv4asOhhIHTEfpAWXWyPotPzdLDRbDpbLiV3c0P/ODDanzerwtLdPSlwC
fYZRzyKfUENyUx/t3hHEzJUecSyTvIFfdhSIlo74uy3l/SLnKXzRUbXIDIOOfR7V
pMMFYvvlNAT4WFRev7SO7W6TNqgET+eloEMsI7xShZy5qUGdMzkHjU7O5iFuIykl
4QjpK4urmMScxG2jETmJQWVyHn0lcHPWEc+K6AgUv31NeAiXwSU4KPcKcYVB/TSX
78JWoe79sAUfOROfaCANoJhR3Xo4r9pCvwMJ2NJGx/Tka/1U9r7TpBcUaTOXEXqe
zGDKLU0gom6jlEebKbKf+RCpj+BODJT4/vl7o60/xAcq5tvkOsnxcov5zzuX8ZRX
BCuD1ThH5ET112VxhFlBZzDbW2FuzShsCpjZB8RKIaSLd0zVawGQyh2UZk+IZ9tD
wwWs/evkIv8SBr7TUmS87vB6ys6pAZDAhc+hGJFJBJCgU+wkBcvG/258Z+TjkgqD
kg40b4MauaxUciMqPsi3k929hASNYYWPa/+PFJ6/BkGgi4bIoVj39Wthxary5hqX
BO7zoZwSOrvJVwzWrfDES5FraxJpW7RyUK8T619/QQZX7YujubRXl6q/qmQd/kmP
pBvH/nEs94/Cz7adnkxZ26kCTNonP3DCcASSuJhExOMYZxpBXQZiCXbZD5PG1htO
cvBAHMatPKoOwXP7QeqOXJ1lPlgcqrbcExmvOTdtCvuTkfJQ57ckNbf6onEDPqg2
WN3tcYjo/MyalSXfK5BB7O33R8C3IruAFnLeLaSag4SMQZ+lIjWotGeeis8mLkCO
6xdLxRQ7iJ/GIafWEhXCLR8rkv/HTfmmMj6qY5+pkJiMfdBhpmBttn+9T0ZcvwF/
p1R995H3BWsBXbdJ71jIJVz+m9EszXvKWfV8JNw6Q6/P1+CDtqkow8seWZKuIgjS
mvmBVSZzRT0yUwAOkK8IbnNxQ007aLx/4y3tZ1fU3ll5U2pVC1wb61v0G2Hc49sW
ySoivuWugMlVo5+MH/BLE6kSivzwF+X33yWsc3ClsYT+Mve8I7U1MU7F1JX7mqD3
IjqCIGedQfM3ZlKRLmOUZWIbGd/zHcvtBpKkEgCfF6Lii2ffaH5mmyo/zEsbdeSg
YqOaI7R1ZkszPbmJFmada0rhPmeG/7Gixhb7POULWFd6HducDWbHwJKcnpCW3SmK
cn2hq4wBOsV8sLzZoBTGmYLKIA8smnVLoeEwRGShMxggNbiFuoJvaXq+6HcqulPA
347ETGlIHJi4kG0HmRFPHfNMt/GBSuU9AsM9D/aBlvBf0CNIEUcK39Jjqjwn2Tgr
UYmCuYnKfJSRvxPaCRqNnp0KjPOoiblYeYKhOMavVIgNmZBhYxOUxGTzEIQUrpYB
jB4sIiLFId7YGl+tkLKj9sELdl9QSWGWp1riCwLwhkEE86t7ccywdDKKLfwaMxyI
K/FEnkUtHzKVrdbjzdwPfmuPphLlJCeQSfsatfYDuyGKlAOEKTa4/zsmxN5duxCP
H+fnTYWCGjeyhUzkeJlDMxYzMPhDaswFVOpdUG1o90dPo7EyAxUjzd6Q8aTiTOcD
CWhqrulYu1u4gEX1eSx97A52pd4rlA8sLQHixzjHAfMRd2oTxr+2tdtQcNaSTmbX
nwUA5PysGgqhFoM550EP7VcBNlYalcixrWQJuqsFXpgK24LK49sBIyhb5aFLDdna
tpK+rJ2ZDLNrvjg/PjpIwqpU/2mRhhE+Tv9VOvou4u/8LldYuou7Aeee7ri3tqX5
WxYN/3v3ASxqmnTkTgUP1xEuAmBjZ9eWIpPc8A0y9YSsx/kEtWzGlOUc9i1vuXdR
e5LMdaLse3sEeLD+D5rqHBccznHdyi0qlnIGH+zeVRAu2X/pWdriqH+o9CskrRVz
+YwmUEtt1KzqxaU/JZZjP5kIKc5UYNwqkrGl0AfMZr95L+XcQskU6CgJmwd60VSX
N5Uik5ggyxXhHNOFbSDmEzQfSz8H5Dme1nIzmL6rsA1QK8ubUJDm0mwgddpQppoy
Yr9WuTbfsyYDpMzImmlwqpl7aM6MI4cQaoyBM50RlvIDZESHYnoUhQzXCOQzOUUa
z6dOPiupo73gegWjjCFegaQ1YL1hWnqyAi3+U2dnDalP1D/FOSADZGHJ6oh8WFjN
jbCiiFoX8xzpOyuxlO2KItNmEx8YisssbabRGhZlsxA228hg7K40z+Drk0a14S1/
j/L2hueGTEYgW2kj5inq29fMQ5YRUvsA6OVT68IhAaz6H6+ibgb3MWFaor2MSmEy
lg9+UaoPmlb+5lVqGZVyC2h86JQUEhZ/jf4Lyw+H3OdpUZn+dWKbcIKv7fWr82bY
OwV1CgAtJmCxRl7J4pc6iRN60MG5V7yeKx7oC0ey70bfexCnPaynY/dvZArqWliN
dNH6AqgtkYB1/3r5VftCdFraS3WQW5jIygyMISMVJ2JZ4iQs8UDpC2lrYJ/keQcr
vCJcnYFYFmGKNEgzp7jvD+vKoUxWCElgjkXnkxV2rKhk2NffTOnmRN/onBlODZBB
6o82AsTgBHqGVhNkPXBMLp1Cv7MoYWVurtBY9/RQDCuFiIzK1O0W7m3zliB4QPUZ
CGRlDLsM6pFhhJb7XLOmsN/hEmyNUZiCkeSxx3ZKXxoZtXrm61cfq31QmfjV/NZK
UZlpQM59uz9+8sJC5O8P3KcN0vBibGAp5wRXrpnq3Vrvn3R/eANlPWpgKy2nFsjK
sidZ+rSEE1H4p3BG39kYJrIEPTMWoMyrTklzleScvgTqKNtIiEtFMaPgpr8LyXRj
tKnExhmhln5nchye7DIqxJHb8l/z4spASl8DydIIczuZrUrPtN7hobP0V2LP9Zzp
bCoMOnKpc35YWtFDW87/gELNJi/B63xMUP4SEOWzkAgVAWAAGZUcCWhQyST2LcXG
c1NHe19ipClWU1hgUDypkKLGp6E4qqlCGQDnW9VvYxibYo7vMqmJxYdzXCtPRe3w
ynupJEvVYn+zZP0EFDFjNyx44sUtYpFR4OWYOP7W77FY6IbfEFs1J0xjy2ckmSD0
vaSQFuZo7AE5f7kc0vOuU28kIYyt/8duY7dsNJqfk3GWg8G4tixVNOp9GNWEwcdX
TBfVPJl/JghgDJGwUV4gmAbjjvuz+/sq0ZoM7MZ0S8hNrQrhftyt43PpRxncPNyd
z3JZ+NWE5/JJmdr26Sh+oiOqh5ayYtsTDqY6BLq2MDlKg3vnO9ud8+8aTgr80UuM
2zkrYVJ8mZT++ugj4AL/51gt44wgwpj70ITq+wIMXwD6lIwjJnN9SS58RWGBRcqv
NXVx9jgyeNOO7xUnWjN0kOB4nUTXu6s1g6SWtRbOfyTp8FxiWVPOB68CNuwnnEQZ
OfwFGzJrVBOCjdYf+3R49UlRiO0DRTivW2guqTAHEJRVKpXEJDZT4LD8dOgBl1WJ
Xji07tll64pH8e2Xeu9ecEMF/GGqBUWyg7Om+ExVpIbfjhBNQ+/w07QA1gXAcHmY
lo9ByGZk0lHFQ5WSZAz8W58LUBMf8bAXPP3RsPIAB2goo+wwq3E6VKWutQ9kapt6
TD2tBpUixRJfN6tIzk/WJaJF/t7Xl1URcNuSa2cGE9H9V1LEZmNoMSbrctBQSbGa
9O01R3PWmLSr9pug9hcIVOit8wvx3HhtSfGc/CAAnc7SJOuNkBTWsrmDFmzedkFo
2boiaRVICJ+coV8YXsn+wAoEFXxfeKquEb/NUytAkaXhahEL9G0e4HXlZhycWCGr
roP//rKzFjMGP1ekuBrMCM5Z3rGN4MyREoNg0DVDArsWTvbYRp2ADnr/dQxlVnYp
OD83JohnhMkz7t0SFA5ICY+DXQmMAEVHL8240WL6iy5gTAEaJRosc0SfFnAXYb5U
zP8UaKteNr8JqDPYYCQAwstI+80ZWf73j8b61TuTzUIzJIQyE3nUp+8NmaSN5kQa
L+UzVxBA7C965/hVrBdAmgPyjnl4suIjvC73cUlzLGdqWVV+3aPoYfzX1R5tnfiy
loFt0MypV0p+gaMwonTBMFh+c6+QMtpv/S3/xEu3vSNOAs3z5dLY3qCNANIY74d8
rX/T84tPylaXrnkjF5/GzdvRtSYwinkmGpZPdlUZy2eaYHG1ug+gkFtWScUbA4q8
8lvyzxuudFJcLllzKD17InXjhYKLiS0TbDp81fVHVKThkOd7PArNLHQi/BEVBdYj
Q+1llxBRN9X612kDqRxGUwXFdvg/WXUIhVpEx4SOe1EFbByNWagJ7xXam624hlkN
+7PTbqMzGDDwTlQDafghWl7DA44WFrUZoXPNMhZPq0spGG2QxneYTczQ2NDTBEOx
UsGtdD31DarGlEQFQT/QNkLbD7VgmdqfHl+4fQtV2ypmaZJmBPqLNc3lcGyVMK/J
4IhI/Qcvnaexyz0kRIrMhvcRpCHHcJh39WkRv3UW7fl9DTNZewxPrADz4dnDdPfy
Ks6HWmr6ueiOIGgyG7phwb/eRXh1/ihrcMk+tSYbWgnxwrsx3n/QVN3PgHJFOKt6
BI29UTkl4QiUE3pwTbLNifeA6kKNs3PO7r2pt2bCXgt5ix4o4UT2TLTA3Ym3Rmzo
rIFxpZXMM5eXyBMKJgpEy4Gf9R62knDWb52xNU19UYlkg2j7wLblIkUYnx7cUgr0
d9jY0OHfoMW3OtL9AM3zl4MHBG5j/8j/oxji7R35ylGHxU5zcSC8/2iy4LH8t8A2
E50rKr6XGe3vjaDjm1rlB5LIPgukAqqg5MtpbnR+RS6KHRkL/6K5Vq86yLqktazJ
X6OPC32+RynmMzAX+lAlCem4BTvIWJl1lDvzxOh6x3WmVm3d1oxaurgbEH4OMnsM
/Ol217wkW/X2uurD9QgA+eb8veHCsAkmPOR8J02d9rov68uVQFm7wdxDoc31JA86
ZBVL0t0rCPPbSxX5I6ncFQXQUbS6gC2hw/LNdpBcCwTyBr/Ya95W3A3cKRAuW++P
5V52FL5NUgLlr2kiLol7JHg9wR7T6lMTGiOtip5eEblm3t3q0aaJ55OL2cZ7B8kW
km7fRC3soIN9o+BkS1B6pEzocBVdXgny0Zxuuu01KkcLS80A6w5DkifZTWVOPyPh
vEUB3pvGqd6x9REEkd+duvtFgCpEyLGGO5mFGuqtwyexEahrBl/OF7H/toxTz5rL
0bu/VKwDx78RzO5ug/e7hq64l2hAZYuNcdy//OgDtVI10nE7HxUnbKar92k+afuK
peej6yo7/h8uhFziphZjdLZ1j+a5TdYngy7wUx1wzU718u9YAmAOCvVxgaJKQJBm
QPsMnexMdtA+GMsHjpg01hCD3k8r79hhszCMwqFLoYnLz4SxmfKDQXLngqd3dHg6
ucHscCYdX7XDikiU1DAIODzhnSbXRg1U1A/57aBBac63nxPHXuPYP/0tQCoY6MNQ
aEpZV4gt7E5vX08LLSsLIPuyDSQKXligoBEreDqGjykjKD7p6rNvdGs8l4WGO7B4
6UoaKiBudSys92rvIFLcygtH4GUOhfd5DcXgRLPZ8zzAsKo4psErzPlf1APncvFB
Nk5iuvN1fx8/LgYGuMHNCmgZmGB8cSQUdYGHsyLXPjQ1Q7+p8ZOhmnpxH0Y732E2
aTX1quCsB9xjtaBceKBp8992rZxDsQK/+EelOWtw/jxbTuEkMXkTJMNsO9Z7ESkW
r5li+YrkiqnYvlWnIhSoGYffzh0BVmSEHECBBJeyTUkzBV/le/bIZV1nlsYFqOyL
HbLwr6pStnsocmVy4DuRe0KAxRYnE3UX/bPP5UAg0V9EiulVFEi7iWS5e9gAslQY
L8KdRYURqR771FZDUHZebtl7OdCA34k4fYgjLfhWwrVltvAHfosJiUfXGcT39olt
8NFxTxPYyHXPM05wlMBJqMAg4hGIopgDIgxSNMkM5VY6K+D6M5qJ4ERVlNbVsTbk
KHbb9+vtKqfVX88hvHgl6e2nst0TB9rsCoi/2XRMnperVERlep1XDrx2YEalgi7a
neg+twCKQJEPV6djZ4NHH3KuQj2+Ffn926MV4+hXJwU8pRN2ZCGYDfvbMU9AVJBj
3DtyoxWxIkzauIxVkR+ZoXFTzru7XjjzLq9YVbQcql7MhLZHNNXkGa7F8s/Jsp6j
qK/aPnianOwh2nxXqyb4n5Z6JsWG6smQYrnmSNXc9+AoqYF/MtEByNd0V7MR0KGj
78nZo8uIK68cd+IbgHGv8ysc9R7v7ZV9BNtAixg/jAfl9nlrT2qEb1NZP6e9AFOF
DagXPlHH0F1EDXXLAPwMhPxpar+0VTdsM0e1PKd4mCKc9RDetj2kHtC0GCGQH7li
pYPVp/kOI+D1xb0sUOOucW3uqlmBrmU825Fa/qgZWR+VALFn/waf/ZY1CBG5obQg
7TRHwulIz4JO6g2P78uFtp8JVYIsLtHKHQ24MfCcXioJcDa3lSBbqvYO3EsAiq82
11JJt60puCRvYiAi64oe0dsxYQdnD5Fw+UOSYF8QJS3a5Dm6V+TEG8bEixF+k/y5
wZtITJiauJSi42n05TFQjdF01sIZX0P81aUkriKsSIn9iiawwGvuaHA3dDvibGQU
DZLmX8mMnnyq+IZo9P6L6t26b6q4gbBSX8vh+cGlSbIqzkiTDgZv3WA6QZZKNK9i
a7WF7ndKwITz18Dl2EVPzZI5to4LjqsNoyZpakBm4NWy0A19wHtunp75dkYNBH1q
Yy+suAbM/rMR03VkPL6TNyO/useyikiIISlLJ0+NVxkv5MWRqbmexUgn1pB/SxuW
W3DTLRAabMLuCAK5No5IYUtE6i/WrvA4STo7FlIAkXsyePJwhMKsOnJYdsuJAF8p
Ki2ryqCJA9tUqrb/FkIAItapx7aLGkFicMy40pVsBDej9foPZNV9iMSdaPykhMmt
THm0BxvyccNOOzH6Hqyz3fIGRc7zo1i8+1p++UYFFkGykECmphn0kAS4acDcs0Ft
w4+YVwlnvMN/zXxzJ4DJCHe9drWHQjOEo8MoE0yxfA4s5fn9qLIH9lc/sd5ch/ml
xZbs9BxJkwAbkI+R+XHoSlpReif4QJOMCj3XvUrJ42XImB4Pm20vyuwXLSXBpsR1
bNq3RiFJFdWmWtldbYlL9sDY1LD4HHYXW26wcHNzqvoJyR6Acdq2K9BmeUOAR3xg
2trp34y05TF9U7lZ7ZExeXTpxn6unkd9vL0QN7hptqQ19BkEUmzfPbjDbvRebP4T
5P9AO9C+gwFzuPkd+l3L3b2JBE3nTbMtj3FOA9ZdmUIrr5bxB5t2eghcrDEZaxge
UgkFCxd/oQi4653qR1ZHuRd1iAEIwH2xfayd9cp5qu9thw09FuzEn88sniiMyGYW
a2jCaHu/59iwUCvCQMQxu23Gwfr8SkYPI5fKHYhAKJMbqdXup1+EwUl8cuqFU80w
vAXu/4tFh5aX9p6x6WWwqaXLpA6JfaHSO2jxdIFP/xAT4fxiaR7Kd8SBZwCKAJLY
/uuBxaaDVyIVSH67SpWfovfKttRzBr2WEaaBYX0qVxzpWzlqInwD5dvS/NPiqpmW
gH1/uL5Cb6v4KRUJiTDLLoVoi9XWf+/I+L+RfAIUVIDoN0L5rd6i3OCWjNCozQOR
YrYVUsc09c2V/8q/4bkmOJv1n5qd4tEZQ7VEpIHzywapYmkt1ytXJRVGp0S8StbA
/y5xIYbG88N5l6gUzH5HUWw9exHHwwh6GpAFm3ETabV/m7vQp0qXcbIKVy8N+WtS
HPC3lbJ5rt3Ed0f5gkTqObyPG3dcdldwm52hF8GS5F+AYUZ0naiJWT3bZzIP/wIs
A9fg2iuq8Yqx7J0jSpZDYz6iav2Acr6N/LeKcC7llYUlkqI6tmc4xZAEYVeQfR9f
uGHI0TNBvfKL4qO/1qlCBDs6Oix7o2ZI/4vRZ+kG1JYZFYQ4WitEsofSfSJWhxlB
IrmAev1zhXia5SXrmdY4wJ98VOZRsJzkNMENAaICW4WdurkZqlFA3QpUcpAjDEhv
VPmnFVp3H9YJmu1g9txuMmWCjhk3saQfAXqrp7Khl8keUMwy6y08QquCkwomhqWR
zCJ0s8ahZf6RiTkb8Y8eksYAx1KNbecb0XDAGsGjDlKkRefUYzM+RNFvyWBOG59h
eif16drj2lHJQXQWK1rVGTU26ePqTeGpPc3psqCeKzlQg6heOXvCL67qtOAGtTIt
UDBKjkN3VoPRthH9drkSQbuayAEH7vIjKHRdL46ybAy9WPLm/pJ8MLXHEj8ZJytC
I+U6HIsGmlHMb9pVeuQDN4EZMqXiX3rVoMGBgrc2ZFCQvrVByWzD3OMo70CtmnOt
wKjvNRzwyH8iqkrB9e5i9Y/Qe94U34inOfVo5P/NPWx5ENgimLeF6MlLolmdXfa5
Y6+cS4DOAvmo3PEbSzF/x/zTZd05LC/sNerRPdJ1rq3qEsnuZ4wHzQ9zTzrH5Oif
NsraIVzPnLNTswkK6sX3tzrXb92Pql1u3KvChjFAyrMTQRYOXoVN07GFgC1/tO4y
z+Ss/LwgB+XxWyDiQnNsbwW04By/OFe+wmhLoAIDkUIVzvXVKIvuboHyyFwZJBzT
dwMd4FnxIswsikTtom5xnE59+rInhlsBiwzg3BJ/Q3Y/eq32vmmjBNUJltwdn3et
I7067CGbTYvGgVYMnYAl/GXwrRzaISnRddgFxHKdSn/mIfPwQlPIUPVzzMPBYQ7y
HftH9mHaQwn4B/Yx1m3IC161BO3H2RakHSzj1c1/Jm5eP9RRUW7QeEStC+/HWihW
V/j2psQbyPveUo8Q1PJDIgCLTg9dU4yFOdU3as3ifwjFjsLYnMhU8kDS3SRMlYtp
CDe1IaZtW1p8p+VxFySe3jH9l4puEm2Q+n/KwlJC0o2E6NpWu3B0xtnC2+cseL2W
EIQGtr9EQq8d7XYzQYymVnOLwrmxTAaL5DZF2g2E/os6kmjY4tm+NVo5rEc/EiKw
aVK7Tjdsl+3PBHDo7SGY0k6xjgFw2HAkl3EXAHR4d6Z1RH71voMY+JFDIr/6A/aH
l2rAJmD3yytw7nhWy26ouDoQDLP9JNjQynL9jmePWwlLjrSAteTFFrV171nXpxDZ
59q7xwGlt3r60Pba0+lRABCN+rhbRAfJgm7czFjPn7IXaXeLsQR0I95vX28YbM/4
W6wSQobgNn3JhBzIMNY8Wu4oYihaV+ODdAN2skebh36u9Ide1xdQm7GuvctI6L1j
VSPvYxDJTlZZEaiwiovldSFFfrpgzDBycOHcuQKnPEYTohnvqVG5D4Q23nhrk7sL
B2iT8OI8doLW+e/wb5jHd2AW4zfhplu9jmjuI545mvyIj8AAAOKKDB50cCcxMuJE
0j9qf6yudqzMCn9h+t8G2mq6OO4sl/IAVZtkDW1AqKAF16+ifgd1y/0MSXmeNpgL
nfXRHp9PR6w9DepDr4Br/IpOIuzz7BEBsyWALh4Gmx4DdEFsuJCPw+czBv4tq6X3
ulQ+hWgh7cq8S/hv9Q3gEO7Lfyzo21bS7h7hexBoK6YVNwsBLsTN/p8OYIDTV6rT
qmx3tjdwa/hdMeNgHnKWAfRYu7vNeC95xeOJ7g2+gINsyj+/imP8PIopnSP7I8kT
URbzHtjoRUcdhD7HKA+vPTgmxqNWvO/PeSHfkjUuQyy4KQ8vJqwBWpxPGOLPN+Cq
h8Plwtyp+30dJlP07n9J7+KALYTNdecM1rLl2hIK0o9u0h61uJ7ZH92bOjMhW9ga
9SYK85naN1WgGubp3IA1DtHHFhWq3/xIwYsFAomDciy/ikt26BfZNOHud6qfkSC2
y8W39mJ2bAdeGWWqCmpg69d1pX91dqpN6y6GNQDjYvQxs9m7zEs5GWgzT3MrDAgq
xpt9o6bSYlF4r+Axo0mZ3UNrzq3/qMyCAFuLbTz+/cdUloWjH7VBvgJzQnrpcdR8
6qpZm+GZENyLRbw++2EVLAUM5p/fxNisdv4k7zqiJbJq2iiGTUs35b0o8KCG47ep
/WJfY+cCUpl1L1w065CEAQjo7DmkOsE2CalDIKYi0A5mtn1WeAQurQy/RTjVr8VP
6r5LhTrV0fXpqG+T9AcB1yXNO6JDt6fwaOrNKzWAPVIkhD1/ZXBuuKTeOYiPHyY5
VSET1y6Ha1SPWKkdd4mG8T4tnvZA7Y+eK2W4F0vUEJCIT029C1OA/igWDS9RyGRO
2z8vfnHGEcQ94zt0/PhPcY1970U5USqdTFoa34YO6/IZ/XPDRFiK2OKNkUSLrPGm
QJuKKZR+S8u0y/GhOQpEqQaSmB/IqGKB6eNbmrdGdQmYqYKKO9S5ZgDnpm/qLaUU
Z5Rb2K4Gz0wuJLfrGfYzVohxIVwy9Cg3i92RfPA7EIUEdkszhs19MO4TCzHuw5iE
jIC2dFn+oOZ2aZQk4C02iRZZBd2vc6BI94jvlkZr5vt6stWM6ff0/C39MqGU4Kpj
g0yrQhqIm7lZQqriY4Tutj+6sZEUgHR1PPAWiUsVQXdeDb0gBYBSOECYeJb4m2la
QLgIyMHls1exzCIBPXhXa5UQkDDtmKW68/ouSZGkIqzHdbNtOed+qthAhOSqzZWB
wzuWvx8+MMQNeDQhM70hG0HwZ85qwOUNIsqlbMjVBgdUc/LSLAiMSIwg7ORr5vOI
rguxkdqlTBhgpCmWaJIL4M9Ea4my2FPeDZef1J46X1Y+e44Tb2UqJGEUIX1bfHP9
i/3ryplh9ZwlFWiarbQdTMjzZvDvN5GFKueDHQaWiYyDncZ95AumFShu/yoGxMtF
wMNgqgTSym4IY/c/dgwUUwlbhEiOqBz5TXl48bqeilrSA/ezo1QSYPBP4FY4tHkA
vFHSINvFJH4lIZiyl5ww93SU5WrVuL76rOz/78vaYSwSpvdCM8U2Cqp9TMXgIg8Z
CbwN2qzYp1ljgwyWCNjYnaFg5oUrCt9E3M6Zf6g6eFRZKX0r5ijwukexr6KG9//6
rh1kDnYs26LB+5FZC9HeBgwDXnw9z/7SRDylHIsYJhznwUl16NP9S6D6v7JT8fAG
OEAA7tNm0vFTsmsiv9ojC4dW/+ZGAK3t2Rv2WuQ6WesbWrE4JJAxaZxfOHgZ3ese
NCY1YlRRDh1QISUIqxAzwssAoZb4CXoOabVFWHicgYeubNZvDP7Cr4Gw5TQD1jh9
CipoSpw8zv88jgkNyjUTww0de4iXa7bfhA8JUi4nqaMDPtiF/FTHvDe34J5nQeYk
Rbc/guXBHdz2wGXPOLP4e723sKJdX6jXwE8Ic1gUHaYcDls5txzebRCAXQ56d0g0
JPrr0ZDQ7Yg5MQUmU67CapdqhjjNXwM89LcDFJ/mI67Dw+zqmvrBTiuC5wwde86/
sBtU7KIGmewvnTlCBcHbYPHxdHmhv45jjYEnZQQuRweOIwj3mnHxZl/U9lTq/5G2
NHQepHS/b4FZ6Be0bUHsierBchXFyM+HrzqdzROELdlRV564B0WdCmq/Xwp+3fAk
g11jRkix7KtOjSeIyfRaaDHXwBv7phVJT8Ayujs0kWjp0OHVHjMduX9AL0DJJWiN
3lJtbXvfNXZSXkOd+wKibcQLZIhGA3qdHHDMZNAj0hmdOjOadKNTHNz2ktSufkCI
RBoY52iatudhMzeDYAY0F9umUZJlhRBi4V/NDXOFOgTN8WZTYEKb4ajl/Kcrk1Ra
n1Xv31UWRhOpLUH0H6B13qKLnkDLYOTKgdaVTCNxKRZDqk+oEollASNE1YVClG41
yspxmZht6CopfCxvwWEdmbYwwCpyry35UpgRAhB6v/r5EuTd9+JX1jgaqncgsvab
wmM2YeUbApfuLl20KvJomweDY608l69s8WJpGUDiaRk=
`protect END_PROTECTED
