`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73CxgnlJ8lRSmf3aI2M6QsxUs9CExbnz8/YXQIobmrcHLN
a51t1FUOy522uCilM0X5gNL3OFP8UrbKXyhb1EF8cn+cIMIPKpQMmkAp+hKZY0wY
02j5+rrgjpPO803G/5crrxYBHsgQ593mC7rxGngclH713W/Flyhf3lM94Gob0JOq
VLsfVaQlTKE9yijIILwSVEpYq8Ix/sUB74HGL1/DHnEIv14NywUp8MiAXY26zfE9
uW/BwhGc3wCGGDA1H1+k8lb0+SB7sOm73YPHTKniSKPGKSSAGYEdYGplzb+IVcNB
hewgMdB0s10efOWDmlSg72ea+fckkiL4VWyTPFfBOVb8B6nfb/U0ejaWvGUp5X/s
cDzan72P/CiOiuJW2iBngBKmdm+VHcZEZikxoAYYeSg3CpkzsPBgCsBnPwBdlqWj
4uh1GOiYDaVb9IRC8LA90MYX1ansV521hMNYztaw2scZtwG/XIW6lhesP00NDMYf
rLS8tFohRH7OtRHT7t4U6ogvLy+e8L1VYO7dT06ORDjarhLgLqXLuiAZJ3tzUaRv
cE3eHNraWS9O3M9Tq/e3/aChUdsS3v9XF8VxDNOZe4KngLfO6S9GfAU8KMJkqGOF
AZNxAe8aELqTZVjVgPOiOCVYgzaDCrFNAgEu1I8xRGO0RvSS0dovzOUFxJn3pF3v
Ky+ZfrjicqAacwoJ5h+doUNPkOL04GaRuDiLN6wwCbGHF5Mcjy3sfTzZayATdcAx
0/37c37JzwmcsH80IM+mujXjVhc6KRuL99XTUiKjnPkXwgKBXfEStKgP48fmUFSQ
nz5WqEYtBIARxKc5rARxysKkcV2YyzQ26j2JlTJ4wrOZ6nFIvrWYEGPxQJ+/fdzH
rFSg7SNRBuTGS4tJ9wniYtFZ2opLJVTvA7bBmLc/X8xwbQ7v1LVow12GJ68jYmkL
fnBO68RLHDJkmMOon8BV5WIDv+HuLK0itJLmLb1rMBGxAwZ+LbaX5KaunT4P2Kml
jny3v+m8bGmXdC4viiUmmV6HIVimF3PdyRL7njBxwmnYoPQ6SVPps68KdDOSg8n7
gA+wVdbsM+r2BwrYcMpIm5OkHNCgdqtXGr9Ho5/l0I3umKajgltCBrKGcd6yhrYb
JL1IUh7JDNBIx+SUrRSuN20J494J6fDl+Td8tpk3WD9Nd6QCCgWtUX+CILrnf+sN
YLAyWlqrbNP2Sb9cfgpybDaT7IRXbJqRTvQie0KrBP0SbAlN2Xghz7akm/o+dm7c
IOSr4ZJbEfdX3zq9jzbrIr/wF07XjOXXGzoApqzyBSOqtzE1Z45pojWCpNCzY7ab
wEuMpcHp1mxrrkZiA8jLqoqn9jLwyl8VKpFpkFvlbPHIHEP4+sZYUP+o+DQSTscH
AFAATn/utgdikEqfmgzaCgUXsrEnR3X/QWctcidv5V8WZWiFKpCgJ6F13YXM1Zl9
kSXcC1zJ8LAEnOz+Lf/xBiyFz4ubjKln7O/ogtOZLr4hT2iXjxm/RWp7z/170+di
gReNzQsZBeMSpp8T5k1siays6xQTtq4YlkS3oAuvZ6eEGRYaXVKVOheLdLjLw1tC
PW0caB0L5C56fTIBYw/rNznc5r7b2O0rXiilp+qMlj0=
`protect END_PROTECTED
