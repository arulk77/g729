`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73CwahbYvWiOKMVIGgGTbK8zpxd98X8oB7HvCK3aGr/JPj
wNJRCErmTPdp2JEwoM0Cr136Q2EHr5fxoSs5hdt+j0TdBc5Yg8yCA2LCmUkPNKH8
aaxzIMV5Umr6WjOiyfjb0fYVdYPolLTuDJPriZ+necXRBsJjuGzqDxVqqT8cP/Iz
krinz8iYYgOzPTnUyKBbHX53y3ESFWubx7skNZT8Ansh/OPVxbEVom8geiB/asz9
aNpoPrmY+5X0L/hU76Km0Krj1PnMFCEgfqJIabbRvs+3GrgkNNQh0BCFQB3Dt7Fk
GEalyeS3lyoZGh0tc4tol/oGk0Df713QoiN31Bs7NIHXuCL8zkZUGOszzb7SUHXV
phClycYLBIE0aePzUKsqpl5Jvr2Ufb9BU4Hv2zA6uhYtre/pXDH2192UMduolJ46
OYuqBgY8J1G2S8YKuR8M7SFUE86WI3ueGKGfG3eiMDg=
`protect END_PROTECTED
