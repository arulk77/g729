`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL8xikxYYaw30LJ9z08lEkeyMr3lywu3Drchtr6P6dbxyL
IKjn1u4SrxlWl1scXGOkp/lhDcP9bTwFXq3fRz0UajxgfmaUfCCjHDZNG8Pi+rPM
IvcSAI45WLVkQBM0pNfxYkJFXeCr5yc5UG8VuMVc2Fb76/on/JDg31u5QFbZtfxX
NgkVPBXF77rz3O0GX5/h5gAPy9L3cAXdZ9snTZDg9zdyrmiKOsJXHzxjk7Ecv1Gy
zCou6ABMKZUceh2mzS0mSZdsd/g+DYJO/gNnhrO5etNMNMMRURVXRxOHZgpepnhm
+epv4vSmM/njnPgxzmCU+niq870Ddc/F0GF60i3pgiSGZZqZyTwm0bNvDHcfzc2T
6P60VlTFxmSpWFeHpM0GCDP/Dyqyf+c6wHC/hAUWNKoOXr4w3lZMK2as/Zkrpl1w
Q+h4liE6DuUGPGEZFz1sCsn/XByIMef92QW7/intEP69Olekxb3VRcH1+AALX9eK
Vt18y0Sl2PcNkY4zQdkNG2Ebttp4xI3vJXD4nQZEt8/Ht1pJK4+i+EHRc8pMxnuQ
sd79BFa5oFDyBbXAJATbwkAHVtDiKF4lIerHsKM2CRyvbxm1Zn4nuLdT7MxGZn79
FWcmZNsbfesH1NIFNlA8z17Jquo7Yiz0CCzyeXpJWfWrzH5W9WwRxarGDtGi0xgh
zf5hE1feiUrazS/B/tE/j0KuOh2VsPNRWx10tRBmwnr0lBYwZQBYFM3Vd5Gp69u6
7xVUFtKm8MsU6St5pyxIWdcaGSCshT+c83OpUk4OU84uuqtUbly227XN6N0rbli/
UFR2h9Od+PqwC8uatqPMlqQO15ExZriHEAN1MFdKROJf3UUqqx++yDgj0RmLvumV
zJf1l+QmhHJT6q2lvlLjsdNueutApu43jXRWP9g/Q3ldjWf4A7Nv2bOQ/YsZLIQ9
0GGAZBL0Maoc0sFKDvr2eVvQa+Mvr4Am8P7aYa0nhXjo9DYkjlpsKXj27gLHf0WY
e9U8dUqrAl8oZi6L/lyKXUM2I0S1CeChLXeI88N3nSZbiaTuXaCweuzJ7WvbByA7
cgEW1zhW3f9azqrI/YpzyK7PX66He+iXgljSRpLyfDUrG7NejRNoL3upwiMawjiM
ClgScNoqEQyghVix5H/wAGG/5uGlM1K3lpPmFnliffasMvbdAHu8MAGY2Mq7xzjD
9t5lkkFJysooImchRxUdn2NWj3k7ljDKgRYPgTpiW6m8KT16tq+IgTuaZ5mWWMPx
2MLm2TyNSZg8uDCOPdKF8ur3kyZKGlciwHJn0iu+OO0GUCt9RkUNXG0oiwO0iPEJ
/FIERcPh8amSOKR0vDKNGNn9IHI+Zf6E+qd95ONGxTq7uqFjGGkj/nbbFVocADBw
kzkYmX6/e3BEPYezMNLcz455ahDPP65u/2FouWdexZ/1AHcThwRVnHAjSvrkG/lP
sr51EOH56zb34ZClWcpfUSPCb2PTrpQ2uTCabJmb4z9Aq+emhwBjmGIvZq48QaBq
axz0FxzFKokv8kdTOtK+4f1bBzvSdiyELh6cTfxnK+Eozj1ulXyC8GEY/YbMJiEW
25EFhjgSX+LILlqAqfzHmn7SnHKS8lziHsTiYUAeOYOPmoAHP3yxjALf63VL5Yh8
pz2kims4IymVBg/AEjgutkiG4hJpg38F+K6zs77O4SiLfLgrCPVoII+eMge/4RoD
U+Yq8R3Jl4ALd7m/u/gaP/G7JghI107N3HM0epM405RQ5gHhSWM6yOXJPSStYnch
jnR0MJ6EueHUk1+xpsUyGvTuUuvcWdBaNspPf7sbcKzE0NclxV6HXd+VmTIxtIcW
cPUSUMVAafsC19ck/SKJdCu85jbu/MWhieyAtWndmqlHcFGowblcYXDZYrE2kkNW
lHZSCuhkjuKyB7GF0l98xjSNNfAf8v6qZnMkcFBt6BFpj1fV36xzs/ShzNNbbyFE
3LC2LZyJoiyf6JT70yzKQuI8zk2xJmqUZ6u+u4bQ9lbXzTjJUetz6aLobFie+4/T
RPr9G8xVlQz8CKRj29J2SVzqqhl0+jErpbsg35gBvwq1xR9EnmAzaI7BdoN/jxuL
pPUWT9zhtlBQ9u4Mdgd9Att1Wq7bWk0x5qf9gfay6p7MPh1jO7v5FtOuthBiTte1
t0O3Fwz8/ZRSEuEkimxB84mAf24Z0xegOsWVFmEEKJtI2dEpVhlNC1hhSCsW+Sks
9uDGZmJPeQjU0TZa/l15DLdQX+2XEx2farYeJCFp2V0iUVGemlTRAcqwMaSGad67
fbrcVpsFKMYajCsUSDdw2sjyJWq+XRs0ZzyXuUZxyhbuJDxsezRdJVO8L/HvB/0n
unN1B/X6/zZVy94rqmDNHAE/CUnHsjPhh/c3qVz9cM+jKKqRT5wQyBQFM3U1S2FF
18WhWAzoV5WRdrSqYasfUTFD5b+Dsp9kLlhfjrje6v4GM6ll5GctbHxOAsgvDKaw
GZ86LBo+abU7St8eTeKHRESZfX8Aoa3Z63DgnDPfa+3WKBkL7JamwPaUc0AEU7uM
DavTjZJdi7ZSEztF/9NSe99DOvXodjei+uqaR7m0KoMpto7RGmqQNNqPoGG7HK7c
SgRYz9wAmqZRuprnIKQFBurXJb8C4e5lkdA/gYlocX4b0tAhIXO3pok2syR7onBH
KuY1MR0oqysznz66SACefjdm0xBE5Rmpk2R//jP/ZP98sJazmwMbxzkmMOD6lzQ6
4neINopLFWnCe0VnFkMjHFl97Le7oNp7txUg6OTujcghOSQ7GE/4vdDazdoHalHm
mq85fzT0TMHlGUT1gHufeWM3CJ+CAg7yHRAXmhG+Ng15oyt2IGYDdin5YA3p+VS6
wLHsE/yNAzxlRVImgB8o7ovXcmQ8fZuea/sUdZS1BP2qaeWu2pxEhT+CArXCvIq+
RcbJ5LXiH+DdYskgcyYRYJL71sGWgxZGk49vtYKoa5WfMOiXkVx4eBH3aX+QFvwC
TGHmokV0VU+drZDp3oioI/Jbo8hURsKj+LmteAa19A64evOaRW74kT8KsQx3xtuh
MfbG6BPQQE1qaKr+u/n0ElmMhXOJZfaUCie8+8/cDwATtanKTAfvNkOC4xiMAvvh
FoguDxrIzShDIku/1Lg2KeWjhDARIGYTMIzrhx9HtalrHE9EXF6gCTahzWWne25/
MJZ+t974DDjZEuYZbzh7IDsgjQ/pr0fbP6CTlouT2e72BjbJ1TfUJoNLlFcPNN+M
mBA+dVkMUA2v+Cxh1IbkRVwrRm3KhB9J4Rm9tDMjY+UrYScN1rexPSe4GMg6ShEF
rSxivuxSAA0hWcldWA8fejZYfAJj81mnU5mfBQ0pmmK6juI+oAuYZyWdoYRpSIDi
eiTboCegLT3UNoH1pnrfhBz/7sLt+sUiU20p9OsFBNN25fL1NfnQbfwcMv2S5r90
HdTKQUCdAFx/O8ZmMprZltL1cMWk9E/HeEB4JQ6PrhdZ9PBPQJnYEAR2xo5Q/F8e
61BiCUgbuGYOPhN3NO88b8/bpcPgTGlnmAhKdnqHiOgb978Y1ngs0HPUpcr/2pO0
+ksILs9ySDE8NIWeIXiDwOdp997AcJ66j19VZepMc2loCNY2IJ1z72HyYlqA9Qq8
/Z/XVPlJUQp4CtFApVApT0E79xFhdzQpCwojRuvLmqzunAj6s6x7VN3U33c7OWbd
/lV3/8x5Qwmf5RGEQGzVYEi2a/UOy8ZDvOoSW89be1MzhRJBJrehHCsTaWoPimSo
nvPa9x1ZiaNWqkmK+dm/LqmiRhHNzDHGepPzS9r8sK7v0AZkv/VdBE+oswn8it+T
gaBEHnjF08cU4qALb6Exrt3UCmt93uq7d3PeqvrAeayWZeccxCTsxP0rrIaJgs7T
Tpk4U/TJiZoLq+IPquZRn+JYNFLtqwp7poVuQjYXt7GA+gglTtXXbr4gGrt6gTrX
VEBLsbr2Sc/TQFvx7pJ0N5xNwetaYLAT7fcF8K88V9Z9ANMPZUGTEcKGzA72Lb4e
2ezDRC6qzDZdiKzlolw/fO+Xq0Y5FuSBfUKpbhBEeWOZ+ism/1pltzQIx+i2vbyN
yK//+zC16L6jvHjmHOMMpwHgWq56BYnRrxrt5P1OLgBifVnl52ekHgn/STbkZApf
t0osnekZN1OLZZf7VMk8xLWDw6eMZBCOlvrg99OPR6KyOyPZak0CNYrmPmPWDWz9
pmX02zLgsNKh7pc3PIJCz1ChS9y4pI7JrgxFaYGiqhs/ejxxhLKLWlqC4wnutaMj
AV4fvyZuFKWXLoffBfFm04BhlnLGdrvUpvcZamx+AYnS5VHzHZTwZtOp0MZuy8Ye
ENeEPoNnvUb+iMgoLdDeSFEaRfzTt18DQl1+bqgTHWdJCPaPIJcDu7tcaxcx5Ab4
M48w0TLMlL3EAELkfa+Z3y+P9+pr+15+L2P/bz9OIe9cVCFM/P5C6QVkLAwdKlyU
A7fnqSh2sVCpbRGuBI4pZ+bEpzmNn9+pu6IFKeEHHrcRz04GEhHitCDRQjUUip7H
8BolYQFnpG2nSfSZoTm+I46v5rDadEbP3JQ2CJRqSM0OnikY7Obtvo0LgoOMMLeN
0eqRoc9b81jrNSim84NBfm2UQAm3xVydPxPiBYrkLkeJMPmn8Cm7Vv5/72wfx8FP
vclEYSMEIVO1RkcldAyIJcEVsTj9a0RRYl7xHjPyXIjX96ImBppek3RTyh7XeW+m
DwWfNH714Af1JVLjgZ0xS7eyfX19QdLhazGbRxc6A6VW6n2+zvQmAO+zIGrcCVgz
q+d9FLwC/zyDPSwffw/8Gs0do6T3TzCEQZJ/HoF+BBbodmLnogC030hP92uFzXyB
3cVengPAnu4VN4c3NzHc7p6ciOH4rslKPaYy3L/BpE5Da9YdRcsCKEg+TNORkihB
SWNsJoQ3XeXXW2whwv6krDMxr4srBm/LA/kBC/ejPIGzWn2JvnktgSpXi63jzd8F
3vmPt6FmCY5aBA8D5aogoiP/kDIFrzyQdfEoLBrqqxTALNqceudV9IQ+RvTu7S4g
j4e9G6XNQsiCwPk5CXvSOt0w16mQyVgpOhsvfdFkg9pqabdjToTVPh9kdi2OSboC
2jjFUjmzEMAOGBW1aNLQppkZUktGb7bzrne/5tomxOutThRMRwp/OyKaWYQsUq65
44C0YDj+PdszgwIGCZ5Be9i3zEMm0/SecubLTwslGH5KpInr88b0wpu1a/sndN9N
YVaWlqNpUJX0ZRz+AbZEsBSmct+x57vrKnPFpVsTeoNFKAxRfPfyp1rZYlAMjT3J
hTValpUZp1JtfpY7eEGJWNzZaMqnnicZaJGCn2gnEM4YGARP5rfWhxXE6dNQIzii
jfeIxwA+NC22fF5xIP+5FafJynqu8d6Ax8n7lCFUxvooG5ceF4hyO4rKlkVFri6o
eEhhZM6/fieCKPM93twTslW4zIudRPfy7MkPvs1lI/e2eg+IUeONh9d1TXyBl6ii
X6VpMIz/A8BoCjgOJI98J3hcLpjZoM4GT6Ny0WlPg8gzB2ceHZMS6A3S7u2qqAlu
o5h6F62M2J3/H7DDU/aPIREbrtlA1FyW7iOoofPjk7jaVawY95rE9aG/7PuV2l32
FtUsV1QUUdzuDSlFAl6DTT8ecJXfh+I+6ZA5UYX/3trjmcY9izGyfSYVQLWzJAPP
94zX2pgJzKgSI7t1AORwpTdS6r63c6ePp9+Wdfpz5jTZ/KlvRlcwrz4ru6sfg2P6
rUCSlQrRuBHjX/kWrsITeOfeJEafxMP2ZPiPK2CUHO+v8vrzbCRE3OzbQ6J359Ij
YQFGhjObO3y/OdpWGNYqbpIJy31MlFmabsMSc/IuhM5Hyjd+22vCGU0bazRuv+TK
6Y2PNMoXiArYHFTU9JBYmDbTsSm8cYIZssDAdYCbO+al44LHAkNXAIR+iV6ssuex
ZO9fXHvG4HYQm0WDaRWX7dS0oCGPBdrNpM2P/qosv3WsIRS9Lm0ZSLEzyJv0dWcL
RIDauR4h1PYmelsuObDquXnCVUovXtCW/Z9iVIfGKrVmiH1+2l9Qh/0TIayQo3Xg
W2zLsyhsrezCHalJSLT7f/EnXY/1PiuNLFmSMSF2GQB07wZ+9F6j3pBPEvpzYzHq
iziFzA7CEx4zJ+MOnxRGI+Au5O9gGIcH4PyYbKkXlRYr1rGekfEOgWxWqX5/Va1M
GeJ4qPlCiATT2Bgs9wMZWAKj5eWn6ycLl4ug0pKYxm4ojDvNSevxtjcCDgY7AJRb
luoMwh+cbAeEWi2OCjqZmJVqppHnMONdz7JFY5pUbn31Xh/gxA90yTfKybISmMPQ
AnUxwB3ZhXJ0BuegZJSOJ6w29vkM2OvRzg+tLGb9KnV0qkqOSSrCLHKczXH+r3Cf
rVvpF7vZztIgMNVTCfQ1Bj4/x8CLuwn6xZymH5fmFxF3045ulOD4BWKmZ2SU0+Wd
N7pjlhXQojEPCASjsQvibBlwlRNisCskKe0ZEa72Qp2FHPBmBZ2yji2qdp9GIPW+
Cdsq93etHx+WwI8j3hUaRg==
`protect END_PROTECTED
