`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFepnph9uFC1jLF7bnETmY7iMcaYcKYh4tB5d0YcKXOU
+EHCf/biLaUkaxF/fCwuhdtJbbMw8URNn91SfxQ9qMENaiLdakT+s4Kmk/12iakO
G+kIfVHEqCHBVTSiqzESvu7gQzU4KMB9aM1r+28RyyK8pwpASVCm6yxUIRk9GC7b
EIRD8sDPO+pvFUOh4POYFlUCVlFDm7w5eLYXTlPlDbGTnEJKzMT8FrxSUxLAGRYp
vpEVOl98AnHSdyIQQvleaA==
`protect END_PROTECTED
