`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLSCFtP8ukxXoSKTaMfsQ6AyqTTs2EL+xAHwjlmOh+YK
AkSLq5mUEAgT7wIqJYF4kyhrlFkfLZooOzQDnUnZq1twkFuNzQ5NwE8wiHAJqZvu
zobHk0CpA8iUetH0T6Ri7d5ZI4e+JhFGXFoXCbCqqy55P9qMnTc0v4NFlPlxYIhT
wJ5LCxpaE3NZWiEogbwET+zJVz0wOk6k853eIBdubL5asUYz61I6m2RmmZBpuQXV
`protect END_PROTECTED
