`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBb3pWko987WapdCQFgAfBjJBxSsLG9ziUffXVfoGL6j
lFCPThoHiMW2JBXk8zIJo/GnTm8EM6ILythzVIGOx81LGtubhznzaTAg8QIv3yLo
5QfWqxK3+ARuppCYb6RgjEwJJNVbdAxxMJbBerjuBf58KfLmYmdFBKiVWwN+T88c
bTg11HgP0cCyx0ZkcNP3ccfL3TFt+KAcRFjK2S2nBF7bNHQdOPlwb8vNPnP+xQHv
`protect END_PROTECTED
