`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAY6xEXw15/UcCdfur3+aiy/rhawrpM9xCTKmfN3wrdU
al4KsszfYyJ8hC+1WzUdGUJcAUrJDN8TYKAjNJJWov2oP+Ha43EKXjmzRlkjX36U
57aptmp+OdRQNrowO/Z59Mw7X4BGyHwJyRbdgKFwBKB4PZe7RVvCHemC0hZvyIAc
UQUkxCptnu08bVMMoZz/N0ytqDjfYucyA3lmBemKbnBYW3qZ+XwLDBAZ++FNeT2K
oWqEs1m4WyXNerN6s/3orn6CpRSrMPKBqjIWC7Y25XQB+jPFgjsLhDYQMjQxcULE
ENZWyijgRDtQWyzN2+oph9UyJv2o+uIQEAaWQ6b9LEnw7WVU+ScRaRDXrQd7OxRU
NohK3yNxuLy4gfETK9jbueR8HKfPQ5nJpM5RW2Oz2C51bBebJSjmWER10k+03rxa
IzRgqlneLiCBOXYpr4lZkPZPUSe9j/w3Zi6B7nyj1D+ZFULIzjCl8crAMRnKXoIK
`protect END_PROTECTED
