`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aTgX7oj/qre0cbid/yMRWitThqv69F3VGKaPC/d/L/5r
z4BYlwtUn14k7nuuOwvmYCspi4TirNUq4LudeNRh5NtQDmIiWwW9TQ7uXl7a8hPl
SL166uhAIMcoYlkfHfHP0ZEq6+ZWy/0wrroAKbW1r3P2cgQ5Qp/q03KqQ9ICIGHJ
nmNf9J6GrtI816RBXLiwoJxGval5svZ/5hnFfOTBZHXbwnui15N4ypAHrXif65zz
EIcfwGSuIRRTNVVUf/Eh5g+yQ6lVtu+2dhTTIFuGSGaxuyiKbK/J+OqGIiIoOTzb
H70V/csZTMmtEnflyVLMeMOQ7tn/Hivzoz6rgjlRhijSeDz0S13ZBaNb9WGjSdT+
pH0O87j7vwfhZiNpVhhjrxqKRktj11mC5l0GXZHitsf9DJ5YZdeb1SRXDXBumCvX
aa9bCSH2YY7j4X/jk8k8YSSxfZiBonmd2UFY5ZQRFpsRT6rUqmxqJvVrRsUj7fFO
V7NV5b5lGkOJnvg3Y7tJLEAuWIkRUjJ9sGyLPKOceSWVefI+F94f9sqaUNsrB+IK
Romwir/UpNevYJW5fNsfJJTix6+VsQJkDa9VXkBnV+L0p3fmupbXm/E/NrYSujAI
yxiM3w9g7INmehne8ILrtsdNBy925avYN982kkGEZxQ3PIl24GBQC9PAbKdE3+1d
6ZKEuBvHd4Ja8ZjxVBWIIcYM5jHV2PjOmQCcVEMywGYjOZ6RggzEusgMBnDA6P1k
m7rj39kVyItRd6jhEltv4HqhmaQ+YvhPhHmXf2cy5X6hJjKwMgWGWcKnNxYFVEoa
2eIgHkU4f6ZKpPLw2UIM2tz043L8ApLhq8VaI+vj2T6I5KKQT1j+DXRJcwKjiw2f
zOKdKmxYHaZXYx3QW01koBiBo76WHd+l6qd0ZLSK8Z0zbTanEv2QTNE7Bl9DlBaV
DtDVPVKAoVOr8bgJeFapH0+xIFidKFp1Ay4LtiuNGBRBix91+JDxwW3VHeDtpQVR
Azv4VVqUWKF+VsLullLB/i4UXgrpyliKSDiMOGls0d6l6SxdSuIakaMgtZ1X+fFE
ve1S7IGtgmU8qdW4fZaswnQCpy82A/Vf0s2atVPllwjBevYAjBXIb4w57+pN6JSh
YO6UNw79L0oAYHfxYLNLy0EIlXRpwwdJ076TSH4N6dfniRlAFStn06qr+qPYDhrQ
FuOgYVgLHBcaoxzlJpwzYwFXInVR3nK6Nj91daIrBDy7Cq9stsMoBC8DPgwKFXnZ
EAGdLOht0YcrQlJO2U2zrMZHrHTeHtg6Rctviwh8RKK6NeUHpKhOBx56cc/gdoGO
D5i5hpMepVJTCdT0Erhu8fEBMnDixtKqmo49uaIHOrATbyt7vH4LEu03boU/FdNJ
Bilq6lIyzLAiiYFFxNdztH/P8Pnt7lZnSIbAjxRXcKNtWghg83i68z6PkxnAJz8u
Z5PDuJTAFyghTT6OyWo6gf45u1OXIjjACh0s6+u33SekP9yo/7hVT3ggw2N66iD9
r9BFHte9n2QhuZjgyqRk0Tjfr0qhWAWCe7ax+PCPZ4R54tJVrq3DstGJc//bFj1z
deiNxUmfWUk0aWxr4ReVPiPfvO8owdmT23JwMovM0DchTw1s26PpVYzi+5p506Pb
o2yPJBa6Tc43btyEjI7Lf/ZI47DQsn65tXsemToNnDN8PuJSb8/GYeyWZzp7Gwl2
fUgLKw95ChOEV/VJYdxSAZNbhovHwQKOkUtkR2FcgR5+QuSgZKpLjaUrMrToOd6T
LDnKf0DLy5YJuNT68gm1CTqXCCsYLwhRA4825hrM5R2zxH3yESJ54XdkAtIb7zTR
5oW5cCjcPU/EFgf68ZevxWKLbXNhxrdbDXm2g9qRwejPGH8NQ907LHdTOB+lXElE
Zm/EQNR+SDdnKUDhybmD0jj5FryfXtrHYyxySq13Rpy8z9XwQ47tvJjtOJiKl6wZ
0iPKkSJv6hS+3W0y4pKPh26y7wayFUX5BpzpYseh8FSi1SiLwGoof9acI+Z12g3O
t5AJgJiG1lWb1IOp9VfFGBuFSf9sPVDHiY/lbXeu2hnEovK2V8igFzmC0w22wfBt
kymJzYthcIAqq9hUvDYSGVGZStnodrpiXVGc0kIqxnEALfQUqX++BUjwwGmZRrxK
Spl+/AqtyfPV3JbNkha0oBLsNYyFcFCRGgPsiNV1n2WP3skfNIay0euzezlVVAw9
DkD/l2gdEdMB346m3Y3favfFTn7mjpQFbgQ5TRtU5Tb+jYO8fQGJRw0/U6lIxH4L
il9WGkEbOlvLsE9gKHP8u6dBDSCkfbYeF22M8ezUWb3jYMHjBPndwvU5brypXHne
rtomo2hDI8mI+jjiN37bep7uCBUOraSrULvp/XA7GdO6Bpy+X1IArmmmd2u8BKBn
0BecaM+uHBpU5JKbQK+3Up41IXuOqowfVc2emVDEtcNchn9DVXAPD7hBh7qJJVGs
Kt7S80s8pnw7K1FwnvSC3/DLw5eK6fkaAKqbOiJXikUHAbbBGekGatGNFBQWNilk
LNHVSW0MOIxAXCxnBOWp9vG4NNffZQaaCIZntzaCSxyS4x7unTNaWpSLNnTCcg9U
16406u2Xfw2CvA3IJ2V2xuoEYSFPr19A00XyVhLyn419K9v8Afh6bQOsUChPHFjh
B4VQz1bZ/PS/7l52BdIyvtB0L9eW4hm3vm/ocrjtAiyZX/udl9XzGhuJjwyn6O8w
NY0YgDuLzi9JPI0BEcE5xvoKbHfxzMWAZveWqlupNBzVtoluk4FQZVhJn0S02RJy
DgkyfwX93u2CKyMg7tBXKvWUymfl/5AjwUDJ3qYq/LbDRGKdRcDfSa2FPdzZyZkb
7ZjCzpH9YrEl/nodC2TbTvbYUyRvSAlJVe3YmmxDK+1pCccbr0xvjEC+lhsQbXfH
dDGs6Ba6bLCfIhqt3K8jnOTMD0QcB4vaRohCaYz8lIz9m5fcZC9mnytC7UUxID11
Z2shiRkJFPThovw/mnG4+M42Ll5lvV5qvMe0ZLp9QAZLYyqQ5PkF6q7VB2vUzoU1
i4GXzMoYU/8D5iD5UYieZW8a/pasB6EdR56KfyjEe5NL0OnySmjizuWTXboTw+0k
+F2cqHK1Id2MmfeNriKSErmCrp0YU6XCcNUGZhMeUy6Qh+euEJQ2AY4rF3S2Uz30
TSahE3jZzBJuwxj6GyFCIGFYARvXoBcVRSuYKZqayZ5fUeIsrTEbNvATejFTZKDU
BIx2lEB7Rjwe7B4shLOhfxwsHQ8HPYPYOZ3N5v2CCnIqgedV76Kvs+t9byCcRQ8M
XCP77a02C67sYaoxA3VRmpUGJ02WHf2X1D6GiSFkdzkLUEoZE1pffj2eecsyFy+L
yqx3g9rq5kj217JsXPVG59sE/0ejBbxRMYD9ggwrI/zMzi4c8KL8wKEaTQz1vgtA
YH5/6fg7h5pzen9VjeybQ0AcBSHQZgMZflFrl2wOaf/RB2b7LkDrOr7L8cXKFrwG
pYCvFsgCe5fXGMQsI+3lo/0nHz3nlNL7qDcVZJmGdgK3/G0yqRUgTaBWjZ/fORoZ
2lRNtM7HRJygd/qNCeck3O2fI8SN7Po320vbbBANk0bHNNzAYSJeDklTTPjD8cX3
xZcuuS0dAVA+kuETkIsAVdmbZDtoYJo8Oy9/VWKu4mzGYXTzifEB0gDDYVjQM3JV
e1sSz1L0lCgN9bIQEN4A79kmU4ISOTdPdnj0hKoOIdL1j6LJJ0PHIuB+ROOaeKCe
jr8VMpHKOrPw63K6WfpwmeJKp3RRRmcIuH29i9lYsCyBlyWVtxHLfgKL+rxzPUMB
RoObuCKpUdVTeS/2yDOUXo83wE5fBnEDiYFxHhWf622sCCbt2wgVArKrtHDQSh8B
RSKlqWJ8ayfKOrFpY5WvNyt2waHDds1ztNDsf6/Qn6UfRVxbIZFAcOr5rVhy2D8g
jiY/kIorBZIWSVR4Ix9cQb9famHb38QO1h67760khvFCpx1D9sSrFeX4YKycrh8z
3eosSdY32ohewDwGMZVfk04+LrY3xcN4VkWzCArOOVL9MjR7kEKB/UNu3/1T6TLQ
kR1QaFNKremSacyqwucuJZDGHYQh4dS6NyvapXcXu1emxu36iGeWl4dAvqEtPvPl
CmmRLCtZwWS+Dogw0X89c9isQoUseVj8SCfO9L0FlqF4nZVNr8QIaTE7/M25/6e+
U01JedZh8S0pEc+1kmdlvIw6yKzsLAMr5EBapEkIqSZ4LZIDQUu53j7SMThFQzEG
Y4Vg3anjx02ck7behTcCFN4z+MQS2JzaLErjewl+dXAqRpKsHuzSFZcntiGPyQ5Z
YRffGgfQuthEZOl9iHBAa8J1G/+5L/0NI0HHpvEkk8mTX7J9Vi/gB93pOyZzWluH
dT21EmvlhCFPuFOE+lCit/Bqj27JmeU5XAIHZ8xtyfHlukoxiLZt5GhmQd2GmIrp
VMRkavLWaQjcF5Fxmzi0iyQ/yJi5/4uOOoOy8b+77SOpPm4W1FRb+5v6xnb3b1kF
InfU9ZUWqOGtp+ZMYJ7VURMogcz2TxRWDIuRd4fLJ9L/I7q0heJGG/clcYJ849e3
XgT1pxfCRK0XwJeUN4TbHvP87safo50SfIIRB2m/+eHH/OblPFB/cnff+sadXE3P
+kQtWsOkUKYo4jRMwiS0U+Radr8dZIJfJOS47ucw8jMveVZt7K7Scuevw+Get/kd
CYgf/brXdT94NwtM71Qsqj70XPaww5D6hZKUMbUakofWnnVuPL1Me47VzNcgGynr
86mc87YQUEbzgPXvDJdDeOBabGR9AfLpUVeoYNHg3alXZl1MmLma1K5+PCPObVnH
IM05tagvFIUibmDziDL/1jQpD2Qqgvx9Ms3BBbe+ynkijiRD2egwXlv2oFIiOTd1
QzuFchilWw/FoQq8qmohz45Gxs8TtOCI7hbFAY6anhr5FfuuJOmh8fRW53h1/MxG
ujCLhu9/UFu/it1qyMD2tsoDWg3lNKOal1kgAGI2TJ7b4NthZodf84xa5yk0cT3J
9TAGDxm3wCk2Aelr3KM8jg6mhzlPwNuqqoXwgVSExcC+cPK0Z2A9IoXnUK8gqjO2
WeS6wiowQ66zgeAECUDsSMoVZQq75lRO1MWbwjA8Rrm9VfjC1cfcOfaHjxr+IrjX
gP61S0APoCxVD5K9QBYGS/aEchm6LzSlyZMxMQjgbpKyYCjbQn2SqQHCoHZtr+8x
N2izNnDqIw/dc7jbLR8iF9ROBNDUnnIKKKVC4zQhlG7Oos9g9SSHMPC2XHkR2PtK
3hb+xAU7bxR0sAAWYBDcXseLuRwemmmUzCxlsKgZIeSNlha1G059WhtjEBq/x1Qe
K62EsrdpM0hASwPWO18VrH6Pc0c1oDpStCCwGsOaivrz5Xa2ZB2rYuOVHNoSg4iN
Lz/WRytCJvn9bBlZKO6oeR3xJpPsukwx+pt2kZbOiNOjgY6NexXaqK63Mbw71SyA
hqa2biLxPG1gyguJyBcAXQWJwtRbm+NL34ymvLOrXwNbQCF6mHzmjaiyZJaX2DO/
sW90S/lGQdZyOo2v+/tR760VykEwVWHwEYbBybEqltnWbF2nLMrZAdadMjN3rEFW
EYe9U9ueBkIUqwdxZDHELHpkeTzNcL/ZqRr3WV8d9vhjDMgFlxrp/dOPzJXdXgs8
PINTy7d4+EHRh/q1pRVjxEqLekzDlDZPF5rKxxMabspK1vyuifwr5lZXs8NGCwrg
lOCP+cONYDOyIoOUbeMaz1d8OfBCNp5A/X1pwreYOtGr7CfksaiKSE8ZbP45Ru4g
6ADuKWJHjDycxeYWO+uX8mAhFSTcWkE0VBNRE0rp9WCBjA32n6viaipSUPfCxUAU
XDnnWNrJr+Yq0GaC871HqBxNYTlPsjXARhYSgAFEXXh0ZXAD+q+C903z+0memQIs
fDghE/aSzeIVGaEvLUFMeCebZ6FV3Str4JxsNN2dj0IViQ/eW8r5pSJeSjfgWury
AyuHZAOCUZH2kpBVuWetk+9SAo4TlAjA5jRaGssv2K2cDP6jP1xFGZCHo65irZuL
FqotfeP3pK+YkBGfl2C+f4pSASzztCydYJKTt1kG2GRENSk1fCQAb+/7k+AqqYs4
3Jlr2ec0UfzF5bXQv+e1vHbNzSQHmT4C1WY+Ce4SnMvzXSz6YGUgw5hhiUUhCoTe
Bb1+MtTeXrulzl6ReG30fZuHODuX/DyI288a44ymv6upb6MXT7UF4/WC2wRPK7EV
LF9WeJxcI/OUteHjO0pszSHPPPUieGXv/gFOmkKC7hszt9soYgMahoaknX5rPzX4
NVtO592ZbDuNObfZA5yhsKr27oTjTHS+HFJ8OUW7h9WNk4Fav8+YMFesj0OQcwxp
EWFJbQ8Ww9Aa2yOGbtyjBMj8qCYS7WPevHQsI0ywdyPo0DfcJkKgb8J6zsrwISXO
16Wh6MNBEPe51z372zs7OtQoD+wPuACFyK+mS2G9yUz/kPOZjoHv2TTEPFfZNYs9
zKzLkNqvVD+GSJ4dUprvEcswBcf0v8rXE39m4tFEj4tiictNM/JxWS8ae2DEcP/1
NKDyGjKsSDc/oUTzpNmyDIdCbVNcpe4i/fLWFXIKDOapPfJWyY8I55SeR6BOr65i
CDt2l5kiN8jFGIP86Mmd7DcQT3hx4JhxMf4lYle+AzOPaZtyDYBLPj7ZDJSfRugz
dSPf+aQXyn+qEKdOGqrUgzpOTfjOsIUJviMNJCgFmDGRw1fo1HOmSvYJPppe2dO2
KA8U9ve6EPokgg9lkxjEsC+nfj2UkGLo6eq/fapE5kBQUaBP4orHBW+cGhL4eK8h
dDfAccI/fJZ9qHqWDuo0y8yUVv7wQJYGeIwxNhqhLL3AlavwhKZjzfSxKW6zmK6K
TxyILOT50iRmty5Itiq/heu1hjLzQ8UFnaddhLocHIVRh1jfFkXa5bFq1JcUNwtR
Zvk6ZN/MV+nWtSfRXoSRGp7tSgyGHWwK/ItBN4vqzcRQNDmo0bV3/dTvn/bYiytn
TktTyGzIktew4AAl2p2Ya+Sr4vLCHXCZVeOFOA6UepsgSIbWvOAwL5vXRAsuQCXv
yN5bz5tI+vEQKN4E+j0CTlLeIrA3KuMXrDwnNNLC6L5thw4zAluKii7zNnB5hh5V
Uo7Lz+nkUbvYEr9IlOQwVn1bKc/jy5OZPSMI2NTk7XU=
`protect END_PROTECTED
