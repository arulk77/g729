`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAEygCHlrDbl6hhFNKsw3RkqIq2CsgwMFnvWhCupgWHX
NsZbltJRMy9keXiIMCUrb4IsnifjFfSoiajslNrz2AAZZuDYL5jvO8+NBOfUbH7I
uqwa9vkqnwJYxRiH21IMsLVcuRbCa+cuJDNdl+UxZf15gfxJqz1wJNOFqz10ovBD
1oUgM8kBs/o13r/OqtWusasudkW392MobWi3TmFuTDgKxXto4YcUDhofnvuTV7Po
`protect END_PROTECTED
