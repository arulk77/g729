`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aSeKcpfmhdzX5ZuVzL6QYwiiTXqHvX34vgqnnoNmSN1a
Qzr1j4sNQJlcsekwhC44O63DuhIXqbheqXK/hAVggknhCKI1GKmJR8JEH7n5Y4tf
/xx9rXoNm+X4e0pba8jJ2LbW2vFJbOyd0X/swk7stII+GBIbST317e56FHYXr9s7
4cCSOeTH/r0qcNQuSzsfzvVo2fc6na4/DaaSO6zU7BIwLCjmOAtMdwMOLSVHmejE
1uGGf0qaCGCU2B96eaZQJAiXhH3+aJD2C0AR/O+PCPa4/aulop8ze+K+NcKUg4+2
hlnSG3wybpI71slqwNqxAZ6XoNehdXP2Br9KOV8nLjZUZXvcQvLJ6tN73eiSDmtp
cTBr+d9cicPd/taDmoybC6qRBZXpaevE+a9xBscXbMaPL7XoJp27SyucXCE8mS5A
r9htdyUPKxHsmyrorIf1Xdwq5Qtfkr+YGdygsb91Wqw/sSmDBMHShHyxHP+7eP1e
EwvsMGeu7b4Ta/JftugA5dXMUknWqLWQOK489kaKStgtes3b4z70b/JC/CnKy4/3
FRyy7gEmd/fmX+o/uz7Sig==
`protect END_PROTECTED
