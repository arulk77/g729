`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
vvJDfCfNGFliIOGDWPjtHCw1xuzPqADFwBtojzhPmJ8TCz8yjHOWwmc5u/M9IYHp
D4uXRa1OiiZnQfotAaoK8gqd4OdJaOtqWeOlfOzZVV438SPMhso+j1AzaewEb/Ez
e5NCLPDJ1CJ0b3HEyp9V7aH8FeAM0HlOONm5RRwRbvoTZbqEOJT4im1gxwkhqtES
vMTySpMCc/C65qNBy6S4T8X35vXlXXnFvHKuf1djEUUJ0llIc8oA18npZPwuyan0
`protect END_PROTECTED
