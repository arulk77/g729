`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu489cKM3mB4Xy795bb/acw+URJylO7GbUraBC8JnArs4B
2+lIGHCwO1WlDDyhjDYC6G9PCUdfFld/53AXplHhGZwFt934nSRPlQEhTuo/FllC
xamWleftqm+cifoI1FebT79bBGj3gR8/MF6DwL7rAxqS4pBKmBmpBNcZIoKeihqM
Jb2tAoGYXu+lLRnyiCsfFkMFcWhAz6R5XK4gOT45XHZlLgVrR3i+Y4eNokwmnffJ
q3jTxHpA9xpU3CkuTV8geC17pQ3nwtnaoDmspwNfAAu+u9kMfRdh+tg5wqoCJFD1
gQgarj4QZTCck0MV6CVLEw==
`protect END_PROTECTED
