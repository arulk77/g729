`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
sxVKNtypUR+XyzB2I1bIqtwWiYqWS9RAGnnaWoyYZDzRhq0eIT/KJ9ULzjCojDgW
kZgb+1NqOorxs4a3e4CaK5T8cJAxGQ3+6Ckc62+sUbMygIsRtYPJHlsjPFGdUSyz
lmMQJT4jGBAfwKJ9VpG4jUojHVN6D/o2l7d4BDTBltsMM/8aWXKnSApIf8t2zHcp
tiZ9EKZ5ErJ9DpMRy4XBF/hTq/Q3AErfCMAXfeKxKLb2ttfVPfYuZYlLXu8aGJI/
J240fl2H3VVQmU3Q6uZKOHAez3oHp2v2rFENWt0kPgxhPv/2eAHTNRkHSr5FAN3I
yiQqBOSTWIKe42VvMaCXB2i6/SvNOCxd8EG4Mi6MCj7iW9L7YK/8aliRKGwl6LuA
HOD0giPQlPacAvXUCW/11H8teJtvvLVZBuXkXGAmgeGfzDYwf2vwTZ0RrRJgFZKF
JZhmiYtFAgAHqjWy1MasjDlbBCfUFxxgJbY8jIFee1VxGtnD2o18Bxll+kDWuy2C
5BA26swQCOAE9HrVUpnkgvf61iEell3bHYi1r/FcpO82CzitoQWfNe7LhwOCDYuu
oTy5rEFKXg4+TjyG35QVjNqmjJ3/vU1GOIzsOFv8KqPP3zmts51KNdCWcN7PoHaW
nkscsWqsKkbnIuu3rTMZmR+i/k+UbrsdWLHgEnMlpE9c7veA1DEf99cfFlRy94XL
JPdgaUxBtNl0PDR4ZM7pwXM+2SSLPLyzjhNACcrcdPf92fGqgCCPWouSK3gR+v7x
oCZPf/r0XDC+OXKgJxgDn5WvNvC3ZujPAU8/uERzwRrBP9zLC4TB3WsrdL4fwTri
VoNqbv6eIY9nYeDTBkvA58HWXp1OJd1WtfHceQfKMsl8uihxcfUe5MURl6tb2s3Z
vBxWChdcnDAuJ65VV2iM1Wf9LM4Jijw4f7fZOjl6ogX8LZAGG5lUNWXl3+/vrFNq
GQgPBBHQUQ7WkFPXkBBVP2vjdf1hcbQHo2jI5K4NAbjMWMCaMoRgQlEIbWIPmbIn
auTEI5jf/EY80OktgcznktK/3ojr1E+9Q47Cr6tJFV21ZVqc/33o2olUfZftpJiP
p7ESZfS/6AYKkFSsyBWhnNg3CLqKMsxfGOxrF+bfVkWcMjn3J+NCXV96EjMk4lK1
2fN2cIpDdEgxtt5UZ3I9ZNN/y+ARUV64p/qEbYKAeJ1R7NUpufXJcmv4p2wM7KmP
+05lFfNnSO6vgRAR9gHJrThIL5Qj8L9j186VJ/hpOzd8yuC8cwqvp0pilkxfrVyj
sRuO6Z8HLVv2t93Kms4GXweTQ1upDHPQVosmx9rDaEh83hpMBAOqOwFjwMTL8TB4
UT75A+8PpFT6s/HxNe/p6dJlwBnJXExthZmqC7OvJly5rx1oiYNfDSXy0+DZJsZU
2SKdkNbpW3sIYDmqUo2+AKRPMwkslqqTwQcJg/XEReqZQIJqTw5BOY9Q/in8AAeQ
i0vL07UUiweEzs5h3liaiRuW/2aGhylceQhPxP3U7kohVFpuAXtRqpUi6H80VIu2
Csp5VaZerHchcjnf+vHVCa7Sfz2CiWDM0L2YV9jCjcT2uidJUBDbioXbyhBHX9oC
dyvqX6+qn8kFz7NHM4G0wQ+CGKTEbgmIQijHga6Yx1sd3gj8KZJcL0BDZhR5XxYV
Oj56yTRA+gMdux0WYt6ACOEohghEqI7gWvh7eli2LU16IvmuRsXO1Ne2F63BU/fR
xLUvJ70+L6eb1DTxa4Jw12rOI9A5b/oHWia1lG4ChFSc4gYw7Atq4Dk383z1vbgU
wM0tthd9bwCLhkfIwCA4yeMcfi13EzkQY1QHONmkdFWbeihBMIjUJW3tZ4BfUhyF
htK5WvZAThO3zbywOaRoJ2E/EunMkixJDFJFVoxGYAFlWi55ouGwsNNssUttxTCB
IW9P32KiFUSU35f9Zl5Wf1Yve25AogB6iyeHPcCvOAFwD9KscQubt+8MsxUfIZLj
ViMCyhrNbBzA9fcik/BIodTqwzwsQgalZyGQuxYp03nsOb0jvc6Xx9xa1y9gewlK
m+E28BqHMwM6dqmiDgLRWou0AxCq0FrX6LTB5GdFtautr4pLXQrsZ7RBh9BrAoNa
aOZpw1A4UICHdXq7LFjIN1ZfywS+h/ZiDPdH+n9M7SLMWyncQ0EWqx1GLRKnoERc
YljD7O6chN2ZTaX6UlrTxAskn99mW/bI9P7ZJTAvJ6imNAxx02TB0nt2aGQH0+mn
iL+1nUzG96jyQ3gbsaMp7zT0UUGpn7A9uVVDKmSPKX57WU4WqLIvCMBxkVT4uNC5
9WjSe8BBI+U1BUTjz/Wxp9jd5uIWdrgd6BWAB7ZKMUKWwmu1bGne5kQ0m6VpGitB
tX0zS+zAhtjTL3g3ztQy/GdX3GFeWcAvatFuOe/79Z9FVtiyBt8qDNh1EGXyfKw4
bdB17PC1AW7PJEB/fKoVc73jgkexxbZUsHemQinwlEVr2SqndoCmgzofl6P5wOGH
`protect END_PROTECTED
