`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveH94Ai3PGiT6jdFLtxE49pHBiN78OAvEpW7qYxiJySyW
3I42ZPibNHl80s7yQ91ycpYNa7ryS0l3sa9gooXZn18qQ0tW+ziMd1jWohbHo9ZJ
i1pQL53oJX5FaDjYE5ucfDslvN4F3dVsOnohHPhI/gnHb/T358lMWrVlJ33XBrIb
7t8xeTgbg1i42rb5Yf0UqOa9DhyzeXSsTMt0L5CfpaT+2z5PWdEZ4c6JfqZpVazB
5nCqg5bG+ljUnduIu99cFg==
`protect END_PROTECTED
