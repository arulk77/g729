`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Y24wXqYsfLLJtR1TIefdMsf8UIPdqprlgKYGF5Fk06/xJHpaOzmW42x8v9IllA54
FdnLJFl89OAtfQpT5h1hAmq6bAG2dmSYp+09uqgGlqNXMg3ceDDZla+lPg9/UFgc
ROYEV88xkBZwi1Rx5waotj9fXrjOWpBm6zDeE2W5eG5hRv/SGA+2DzFXRIrJmTBx
80D9HDA2TUGKRvpfJ4ndGV8t/rpvF4ENVe77pgVtSJSFhxuwy7big8qBTtQ0dSRe
ewlkUNKIL+5Y/tqrJUnj2Zl2X0ynyUZc2erU/Kx6kklxLiJucfupau6auhygYqDp
+UWhnqWGK5Xj1HqrFiTxVMprAPR4eFuRyYhme1Q6MYk=
`protect END_PROTECTED
