`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEEYIBfiwp66opaCe00yFTuaPz0k0pvNHReNI6ipLL+P
4SIyvzl3928daACE31ZBL12UauZzseHuSBejvCUkUNFq0CCsUGjDsn3800u6D80O
F986fJNVvQP6vMF/pYUK87W5NoFaVwyS1FUQmf6H58t2rtN59oPdBKdwlAwrGRsx
iLb2cFT+5bwg19qB0XOVvsyh4rj2uXoMVyTUujXkQlufqbQswK2bsWzfwSe/GKW8
`protect END_PROTECTED
