`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN5Mqp8MjZwuusQ+FxqQGFHU7l6HQdImICLYZ/Hx1Mwe
KDMRl1XFZMiRq95sYEX3wM7gdNVw2CaO9cFIibHj1JKxO9i6EY8WSZkJJ7eWpIDK
sSmRRUyiLaxAHQnLR5NytPZRDqMmRNxY7AcD8K4mtp2f35JdpwUsE+XBLN7RBjZr
STi3p9Uz1FbTOMFUZZgWSgFOHnO+cDmi/ixxCDeNPSZ735qGIIE42RDm2jzquvxE
PhV0vzpHTU49c2x0ZcsiVpYB/zq1LPW8i0CjLxG5FE+ln5g56Ftwx57lDzU7/tUe
n4A304GBBWRPl03c2IBNrxCH29ZRIQQZZ7km2YmbYjg=
`protect END_PROTECTED
