`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkWN2fKwjiOujreNHynd3SmGVTcVDEjDTnv+Vwr7vLQ1+
nVk/FDlpuU3wnFandeZOGqb+sT+gySFhTbLn0U0WRJHguxtIyvyh2pLt1KGH4tgW
90BKwIPbgjvMm8iHSm3ozqd3JabWbCZinTC2kLcNQ6HETW5yfwDBJLPxbU3FOfsV
3aLZwFICcxEBeMWnptsBtPTkWRK41mgLNCp+NVCAI2w3/rMueMe4CvNGsGrFUvw6
iYJiwN4bVfDrF5WP888LQWwpE+ALP3t/MbDo9HeZh7xVbT2M7blsA36MakT8UWFb
C+M9y7QB6ETQCuDJSQsHOA==
`protect END_PROTECTED
