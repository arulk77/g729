`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveINKjaUxmUMOn6wQftczdmmQ1z2GAKjl8sXCtKsvmApg
ojN1QkK5plIjYhC39++HfLdnkC6lma/yMcnd2InXOku5iUkmEWuP9gwexIjCYsmT
AoP5fH/vNLpkZEZQU1A/HEc3skdjyQpOjaAeRckqhb+isn1q5uZ8h+DBy/pA+0iI
lnn2J3qIBSdrmGkQJIoujfXozTA3hqjuz1RBbqEyaJV7993tGEfjfzYALTTS+QCp
POq7KlBo71XN//fr3pOLt3pFUiZwMqx59hjbP6M6xUw1RFGdPIf5kUZITbjYKQpp
/i6NrDtgkZK9j2jUJ0e7F+4gsQbNi/qs9vY/yEHAQIL88qx7ft56q5oTXZLVorpu
cYyOahY47h4bDDwwtQEev5C3iX5QJppirO+y4PcTUqU3Ro6f4PSqnO4zJUoh0Eh1
ou1uQSX9Of2C4B7zENWUxs1iv5Fz0IBwIhcHNwQ8YASdy0x9YDIzrHVNbqTyCRxe
JnjIR8zap8+faYl7eSYLTcfpxZkiRNTyyc434fx862IwRX6h73vsj3TJ8hc/u2dv
`protect END_PROTECTED
