`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDEw9vxLUVbpT+Ll2R6ay4XC12DEgKkHEWWzo99mIAXi
1efEDkHPH0YBleV2mNf4KflyoNASR+xdhrmWIBOJqXy17jZxlsGUGII8eyfLCgWW
7IDoHSvUowDRQ+U69a8H9FG/u6BuyYb/JFO9C4GXCjEWyDAK67E5acNu15TEFm5P
4/yP37QzrSQluPfJqt9bqeYU9cbZdtfYkWThrl+J+B5qMprFSjY6gmIDnr0Cx9yv
CodHnKkYcdWk5wJaxZuXbjxTMyMb2aF6/fRJqocSpLBMQcOpmRCd7PYkjQtgVWCt
M1jdcgDkf1PrQE800tEtCQ+m2KnuKXniXIdP85cKQ7o=
`protect END_PROTECTED
