`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP0QfnDu14tHjClkzV/ByO2irOlBpmbopfR4FTlCODhI
vnKStSZCuNzqvl5FqaFdVELEtG4AhKWDgGNfffvcxDby83lCD7NXsi+qABgVGcq3
YdnzEgm5wzCgbcoadmhkOCZVsiqtDnVz/QyWjLLF0T6FXj6OtYmN5sqnnPNZnxRO
4KscqFdBwuEMZ3gW3ItkC1DSgPeB9DKVhX1YPtDyJmA+oTTE+vnTbJ0wYztQ14/l
2cq6Whxkou6/LmRS1ny8WoEdSquMJIkTHcjRRO3PWP0kJ/hB27iDVAtW3HoLBE7b
2VBvz4Pat4wngDhD4r3bsvl0Fc8r4CzRdJOsAmPNNs3k+apswfQWTQb1VJvhCJta
42D627ENCwe+lipNz03o/ytPwlaJCgk3+xDZ7pn84hYqrhneBVxmSvwWeAAWz0QV
JjhrCUnNTSrDCuSZLvBUUBYqieJTSk/TksNxV00VikGgjsWGY1+XDBXzjUDRZr1S
9HGrwKe0gsRfdJQLpY0f77qJin3GcTtki/RvaiA0FhZgB3qtHljAMJ7m2BKmXhv2
`protect END_PROTECTED
