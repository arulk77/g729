`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SUn3QVYQadVUEtvMFQlzRb0cweQVHzx80J1yq8MGgMD2
HL961hZ6/Th2uja7xVqBvSlDKB8iJNTTYwzSxCyIguYdzA4OZsntnpZs3aWEgXo6
nxo4liOCO3pooIiPulSDjgdHtgYhKKpENnW63Prv+xwz38LmaPmXpGI2yq/tPOPt
tRhB2JVmhkInk+bs6pzOggA1SL+kgwdqYWc1BshRW4eNNKkE+2O6MsOTGKLyPrX1
X6N6Ve5OWjOCBS9z0pzoacTF0CQqXQYNkzPplUvTbLVc+MKUgfk0jv+Gsl7bb4dG
L1Lc5D0V1yovwFMBSuv0Xy+5wwKfmLHa9RzhUJPvE5XPR7uTM3zhevYnIRy5kYY/
oBY2pBQ17xrY/79oo4U7UOMwhbqa+9buwnChv/ohq0WC+tkPHJVjcGGB9wfZPFdu
qJyF6i8M9239d1nSbhGSkkH/ev6QYCyEzBtmPwFOkVXmM7WPEypH3T7gfVn0Pp5E
rcsOmmjYwdlYF0XfhCYsjvL/+nOXTAlkYkts8Fv/m26aqHzVYXoQfxsJhXpMDaLB
BzyEp3T4NnbzsaoJ0YmoyGuWMXTnSJmHskf4c0LCnVklrTUKSJFGi7MAoS72gQh2
mbowVPJbyYwG2yzJIGIguZ17u4M6mpKfk9CDs7Rq/2u58jz0g/b3VRQ9j6uhwFy+
CRVrEPDDO/y3Y+t0l5qCU5gK3rpb2HZ7VceohlitJHpgdZL8VT6gKrf/4fQCzGFR
1YF436kmcltdQnPoC4/R7tCmYGqekXozABjMQEm1AQnuHb/vc/UeykaoPfAMMxWd
Y/3/o8ZbVCsC7u5wvSQQ9AFl+S0R7Z9d+ZL9HY1qNL3oDhJ8hF6/3v4Q3siimM2L
5NwxEF0CGGIAV8lDzZatrwrx8zr/nR/7rblyR2FDxEgJaQBobhPAi3SOFcWSXMvr
UOQaedQhBLQ/ZWLn1uQe3+Kxhb5dPYiqYX7HF9ZgOAXWsxeoDwNyhwV3fboOPrtP
AlOqHTzHdn1hCoRPTpgFGiCoHVgurmkwI5VClIkMHE7OPj3/p+hZznfgEZbbJHhk
HjO8uGlIgUa4Oo3UZYCjyAaKdssqw3tQ5EJrFSaZb4oy7u4jQhJQ1nUrQRQCv3IT
aKvuVBt7kYUh4BJ1WraIaizGjlwdf8xFAq4bGAEFrokv+k/lZzbeXpt4/SYwMv6b
i289FDBVa8F187lAZY0anbM7xPqiG45zaTDFmT+01lUmUX19d5Dzz5e+dHnwqL5a
UIVprHWT9eG62daMvblGMniWaWob9b6Fwe0u1CZKMgKPZ08cx7EdZoA80vI/FsGv
4Yc4BLNQq7I93H+Mf7z99gK6hDvk/3yX3pZz8Ye9sloO3vfiIocnt8b/nsPp45en
mU/8Iw3LvUJrcYy5iBGHVA==
`protect END_PROTECTED
