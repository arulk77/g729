`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
J2JY5BXj798crJt98j+BOdINQWOrGiU+bmImzzgwJu7GGzx3+SaInZQMt66NW/Xv
zfiYDQf+50V00ImCsh+MruA1kwX5cgeV4g+5tPYwdYsv+O6QwqPLHa7HI3Qf5hBM
CHoB8wcnxmwnhsAGEYnKzKTCr6EfUMvhP8wgrmA7E3A78X+qf8VWovBGPgNuPOmZ
OtwrVbn2AgYdfByPkWsPjDRqy/ACmJhc6XCfYtomAM5ZruREkq40b2rAc2ZnnPxY
iAOIqLalBZMRhFcdaaC8LpXrjJnxgaEf6sR3FZfhYIMRgtI5BvTPtYZwY2C39Ek9
IUIkxmylJ4p5r90JOxsd9UHrrAWNP/2eSaHIJ0y5C6U=
`protect END_PROTECTED
