`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL54akVB/PC1Z121NgRuZEfTJV3MFZs+KNGEYTHwcU2A
N/rdEUfyK6S7rQLYQItM+4dBP0FUZpK18dJtiMDjC12VJB2iZ6afd3z+G/ZiTgdB
9+ke/zmOwvDHxdmqZmvO1yWOasu1YZlnU4EOWKZP87KfJ2O9rzVg87i90QLaTs4V
lvk9YhKZWQE7xevHMf/aqIAj1UDbexVj/gkEyA6zCC3/SS7NxdAK91jN6oVTF+5S
Bcqe1n6ah1vzuxtC2QisruEiOBrKZwb/xWlH1TyZCIh1XL6edhQTyXVQ9xpChKcK
RXlWvsv2eLqKbCq08nMH7g==
`protect END_PROTECTED
