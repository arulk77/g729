`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveALJSGKiWV6VMIgjKWUVJfx/45k4ib+DFhJDWVqp6qIL
VGiwNlJz5yEUD4NaWagWDuCNC6UnRreDZb3tGtAtFEZLeZtVGwagV0TCLhyivQIo
eeyTIcP4il2xJlxmZIkh/CNSxexsxCo4Ov/N2t355joBjXYeGdpPk2MjpOCtu+E5
z2RukUw9T/FvzelVzHxcwg==
`protect END_PROTECTED
