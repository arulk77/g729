`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFDwsmrwyHbdNxHsG+k7pB9osVfBy0g3dw1c0wkdJXnC
q/qhINb7E4D42rCTHou90I2zmaXMBkFbc+rsrUCxOURSYd4ZEH2ck2ZCVj9kSDqZ
bWol2NdFP/iYnYfAZXsCiPkRO629WA20MjyRxv+4sJV1sUJmQH6yjPRWYMfCBfVK
UHu9MFJkR2xXGJNY3WqlctIBU9b9DSesh/JueWi3lzo8oJvJ1J2z/DfnRCBv8GBI
`protect END_PROTECTED
