`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
my2j2SfQnu8w7vwXILtwhD+2WJapXS/+3pvCwREu0sLofEGWJ4w9BpPeo38bTzIr
g0JVitOu9/oe24n2zILUexd+iU6BPz144qH74XZQZRP1l8pzEIYw0lVG+l76YU/M
dxHZ7fYmurfuRRuPOZvnX3CCz0nkkMhK+YZ6BRIGh92tDOComnf7GpS67Tfz3MiY
JFiuYXyCVMzny1CK12V5Sq4n9LYbaMSFrEReramdBzB6BmSdEkYdTsbqxJso/pHj
5GqQ8TKSuxVp5pHB4Q5+rEqWczydn+/ihsNQAbF4Y66m4mEHG8idTEIVnRCvIW5o
7BQVuWAJ2wENTSgFzbokcO782p5TMYF5LesmtxHbPDPoBRecMUoWZkNMiMIQHJQY
0lOhDwr9H+z+lDwH+nGMJr/ArhZ+IneZyq/M+75PIECr+oLA4Y7MzsUIuZSKMbVM
M9inQoV7CBhXQcW7VtbW6GQ5KZ/YelQ7VsfmMrQ6Q2Q=
`protect END_PROTECTED
