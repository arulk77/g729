`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB2ashC+TAy43VILEIinN1h6QJBEXIE7ULkggoh4SnYx
ulRvQiTDwJJ8aA6zh3d5HfRRLk0AUcA4WRLtIfn0aEdMYbAs/9biYZ2ZQXPg03yi
XY0IiM+fw2Dk7nhDhLGxcYtzE2k7vv4+dRT5o5suc2KS7Gzem1dXNF6hLih5M3ZS
cWwSFe/GtRK/LU6iKGRtoOV/dn4fJ2q3mIAI7+UxucdOatB+dQ/lUq9V9RHLxBbW
g8amS0zXedmhGxzGryHMH9RHIffHbxFnOU/HIAAWyclyiSAj/PtHWBIeLI6bHg5y
`protect END_PROTECTED
