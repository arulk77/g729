library verilog;
use verilog.vl_types.all;
entity PLL_ADV is
    generic(
        BANDWIDTH       : string  := "OPTIMIZED";
        CLK_FEEDBACK    : string  := "CLKFBOUT";
        CLKFBOUT_DESKEW_ADJUST: string  := "NONE";
        CLKOUT0_DESKEW_ADJUST: string  := "NONE";
        CLKOUT1_DESKEW_ADJUST: string  := "NONE";
        CLKOUT2_DESKEW_ADJUST: string  := "NONE";
        CLKOUT3_DESKEW_ADJUST: string  := "NONE";
        CLKOUT4_DESKEW_ADJUST: string  := "NONE";
        CLKOUT5_DESKEW_ADJUST: string  := "NONE";
        CLKFBOUT_MULT   : integer := 1;
        CLKFBOUT_PHASE  : real    := 0.000000;
        CLKIN1_PERIOD   : real    := 0.000000;
        CLKIN2_PERIOD   : real    := 0.000000;
        CLKOUT0_DIVIDE  : integer := 1;
        CLKOUT0_DUTY_CYCLE: real    := 0.500000;
        CLKOUT0_PHASE   : real    := 0.000000;
        CLKOUT1_DIVIDE  : integer := 1;
        CLKOUT1_DUTY_CYCLE: real    := 0.500000;
        CLKOUT1_PHASE   : real    := 0.000000;
        CLKOUT2_DIVIDE  : integer := 1;
        CLKOUT2_DUTY_CYCLE: real    := 0.500000;
        CLKOUT2_PHASE   : real    := 0.000000;
        CLKOUT3_DIVIDE  : integer := 1;
        CLKOUT3_DUTY_CYCLE: real    := 0.500000;
        CLKOUT3_PHASE   : real    := 0.000000;
        CLKOUT4_DIVIDE  : integer := 1;
        CLKOUT4_DUTY_CYCLE: real    := 0.500000;
        CLKOUT4_PHASE   : real    := 0.000000;
        CLKOUT5_DIVIDE  : integer := 1;
        CLKOUT5_DUTY_CYCLE: real    := 0.500000;
        CLKOUT5_PHASE   : real    := 0.000000;
        COMPENSATION    : string  := "SYSTEM_SYNCHRONOUS";
        DIVCLK_DIVIDE   : integer := 1;
        EN_REL          : string  := "FALSE";
        PLL_PMCD_MODE   : string  := "FALSE";
        REF_JITTER      : real    := 0.100000;
        RESET_ON_LOSS_OF_LOCK: string  := "FALSE";
        RST_DEASSERT_CLK: string  := "CLKIN1";
        SIM_DEVICE      : string  := "VIRTEX5"
    );
    port(
        CLKFBDCM        : out    vl_logic;
        CLKFBOUT        : out    vl_logic;
        CLKOUT0         : out    vl_logic;
        CLKOUT1         : out    vl_logic;
        CLKOUT2         : out    vl_logic;
        CLKOUT3         : out    vl_logic;
        CLKOUT4         : out    vl_logic;
        CLKOUT5         : out    vl_logic;
        CLKOUTDCM0      : out    vl_logic;
        CLKOUTDCM1      : out    vl_logic;
        CLKOUTDCM2      : out    vl_logic;
        CLKOUTDCM3      : out    vl_logic;
        CLKOUTDCM4      : out    vl_logic;
        CLKOUTDCM5      : out    vl_logic;
        DO              : out    vl_logic_vector(15 downto 0);
        DRDY            : out    vl_logic;
        LOCKED          : out    vl_logic;
        CLKFBIN         : in     vl_logic;
        CLKIN1          : in     vl_logic;
        CLKIN2          : in     vl_logic;
        CLKINSEL        : in     vl_logic;
        DADDR           : in     vl_logic_vector(4 downto 0);
        DCLK            : in     vl_logic;
        DEN             : in     vl_logic;
        DI              : in     vl_logic_vector(15 downto 0);
        DWE             : in     vl_logic;
        REL             : in     vl_logic;
        RST             : in     vl_logic
    );
end PLL_ADV;
