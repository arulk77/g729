`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAZQgK/Rn4eHxwYMu5eQ5D9TRhFfMQWZR0J3SnEzY6H0
P70WDAgWoH4NKJ/rDlXRvl89rTp9Ui6OEzpGgW0b1CsOFbwwgSSUEzR9NI31iMfy
ZM6Ekqa1xxgLrPWcmUhBb0ClLATigVCIF/OQafXi5uO1Kc1jS85SVXnozJd96I1e
xm97kWA/mR/6dd2amF6XcEPRxDUWaM18AGQ1wuQmTxm+s+W9WARBTdRC2YfXDUXZ
94NEJ/E43wP7vsHlodPmWkTfAhn4XWrnZoclervUU8gdtxX3cy7WXv9dpzhqLvHH
7ncfG2CVH3ogEGN/Twrp4mjtoaOqzwqJhR4P6ED4GD2ITIeBPTAI30LU7Tp0wN7y
KOTRrLudELUMn7+vSSUNul0/EBe3X+15zWNA9QZ4Awk4FOZz5+SP5dsZsi0Tpi3D
JMlPjwh6dEOIwrLgllmXgaPGm5HwqcoyGEAKLCp4RUsUp3929hlHHx0i9LbTzJdY
ob0VwuE7NoHhLyq1tiIjT+eh5Wpht/em88G/s2NyVlabhnd9KORKGIRfLQiZ/1GW
n0oe63FNx9v5mJAeT3y+OK8kvrSuS3ajJmL2zPdKOGiunZntXt6sy80zStk2zQX+
FOTQeKaKDh4Kmvnvp423TFVJO3EIlOa+Nd7kPTS3H6qtSM4CnfFZFrvaanbSUmqf
cxaCACBjR1CyJtHjTj4vnh+ccy0fsh5DogbcI937+K3XabUvBNIlqoT1aaO7ewdk
4T29+jKnGVN7n+G0TutoyDoG0TtqPlHvUMnPKyss7nA=
`protect END_PROTECTED
