`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOadriG6fpPpchiv+6HjjT/Av4/SaVr4fSm7zoWazbT5
R/B0upbFn1VfHf8v6QBadZXZmR/j1pSFwm1/wTMSF9Zq+6heZhe/RA1Za9QlrCux
DpCz5mqkBMm2RsbACJdOeIS8uYF3CgLLmzBsLx1H/FSPo9cXSBXbve0d44/NgqhH
bj2iyXu1EIRwj/Zp9EPrV8Ao6Xpk6DJ7sYH2cDUiIsUb++Uv1Wvms0ib0UU/JrdA
CcZnvCq3WWsvlkXWjxQ7ECpsKCBUxGGpA0WqzXx0ayUAgjQwdARQTiOoAJFMbZmq
vCwqdA3XzmQEGr2vB9a/xs/bR6otL4M7tXKBiL3k33N+fbvdFpOf1CIqWb7oS289
JLdreE/Eu1Oh9Dey8EjSzwt+G2dQkKP943FjbRkNhBxhFcZsoUWsFqqCdA7cO0Oz
8N5Wo440/PFAVPGx/QCKnWJBNgaDqFqkJRt9rLg5k9YK9nDVyqh4i+/Behdhx19z
jvrMImyCFEfrG4y7xLlw7t0vf60hge77onqmmPMyuAcDxflv7s0YZGWb5ZON+FxY
DD/xumN48GQb96/k7eOWj9P/Cuqp05F2yF5GfFDLL3fWV2El3AYsghzJbendiCzh
F7m1y9qzVpnEFl7N3qKPHA==
`protect END_PROTECTED
