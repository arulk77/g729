`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1adBFA/+HFo0MKPfO3coGsM0bjK7KzZ8xVg/Xx29UnJLH
f4iGh0QXRYcLHxBPT8KOuekU81MsKKsCaDVcvoI05Bv+j1dYhd/QhJlSaS55oe0/
M1PzH8rKoMfDIfpI7kG6DWP+j3xkBTAIemgVSg7CqA5uqOZMu3Bvn6ZiqaGRIob6
3F5eQ2PeoT8nKxkNs2Sh62uCF4Q2aNVEvPPsKUO8AOyuzG+OVjqop2xm3McAEDCT
rRf6+cqE5rzrC+3+yU69601394gK8ObQhnHTrK18roCzr9memOoDoCj0QxQD2IjZ
WUva1MeI2x2JIYwLBh88jA1BH1cMYh3Kf8lrhkVi/dubYvzTF9D2Ubz3GLSJ29DW
ib5G5F/hWSZbsULNhoHxfcXJHB96OkFg7mxmpQIMJtXykS0irmvHMd+Z+K2hqeJT
`protect END_PROTECTED
