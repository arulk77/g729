`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73CyLW9huybtxoEB0IYMmrdyhiJH0Zy5IEFpGEvWRRH4hm
F6l0Unl/iDfzRZNQ/K/AnrigBtyGCEcCCpOxDnr7DHz8VHv3vFnwHU6OQOpeKqvm
oWW84l1u58piiN9Gc9VLPLO+f+XmuekH4xk+K9z29S4conZJZ0RtDb+P/z5j6fgc
UZ+hb3vOktZ8pAQLchTqpJUVTOjlDcJeQT8enyVYb+RUF7zdHa6wnSfJ69+1jSIu
ht7B86cCULMTxkrpISedMqc4f++aywumC4aBicM7aXQOg7dvG0a/0RULQ+I0tw5w
LodmwEaZuOHyv0zORMKtFmKIydVF2vKv6EMirrMlpssZjOHsdPV7P1EiPy7MiOoZ
WCH23Ltq2Iu8rD4tXTjHOXdnqAzM2+wwsjR0tVCAfOJ42BDjWn0CBpUGc4wa6I4m
I7gcHnNblg7005t6rUHzrUj/ZTq9jpPP7iy2bysZVTchdhbb5UivGMlIWbCjdT09
3ARTpViHHFhG/qQJ4GgPpQ5oLuNDSrLUM25Ut+wEZi8sirMyuvO536WthHaovxT+
Wu6CYCdUkn/T7u+7oYnqQ78nUhPnrlS/lSjw2aC79N67jKAViBM3O5ibt8kXJviK
7aWp96y/YSrRad3wuEprdB+DGS8xLKZmBbIcn+W4AQU1SD+Nv8UHfqiD8axtTcYN
s0j/q6+IH2hyLKat+ghmkJhks6XVbgWA36fdBR/3FA26ZRjEwZH/29/YWCDqjBiB
rU0S1O4RWwk/VGjNjkYD4aGuvbRTezPZOPqWn22tZSclTzrZHhw6hKOPWIl8jULB
gZFHQLZmL6iwF+nyal3I2jgsqeGSsfU4slZkhp8HKBYb9zNCxo1uv+VahMh56i0W
yI4L+fGgyqUjTPpLT/NSWLuWufZvloCPb6UqcTlxOWwagpEshBkDC5LM509XJuLJ
bUBP6pNMTbMmpUEWLnTHweYE57CXYdmiiSwVnrM2ItPbeAJT/ElmfX6PbEs79gXL
gmoGJun8Ls0C45SZowIUlqdES9573fpJEJudT0A8Zo3ALenLJ+hMyqPKPes5qtCr
U5Mqjomh66fE/qwGJAvldaUuPNl0vcD0Wnlc9sXDLf4GzNYtjrtSRsIAlnXE8dUU
ScdD66Ewb7/ToxDAi6+AeZz1cBoR7Iq8/3mf43stPGD9mdxM/PRxxoiMeaC/X5gW
etVzipmgajc4EJmHcOpdWKPELbGKKzCDKooIhsajQvfwMq26CVFQ8MLeHYsyMErn
L7r1P7vTma55dw9DpTS3b3lccEQPr1UTaZrCB3xu96LL2ehzeHtYMsEl/xsNDe/l
9OwLhynzxXLAQNv6dkHGMwiYkphclmAyEjdSSv6gHyoAtyFMyOEDJk5RNQJoBjZA
Des0RK700EOBwFvYVun6qJyN7ryDVdWa7193tJFF+dKCKGOTMvL10TQsPSzllovH
uxHF23bdX8hgdsoCV8/s0Qt4vpCPpk+JO0LlhqXzKsahjoZY8KFte8lhne1P9L6Q
KCWzKvLqbDgcqVdeMoDjmtx972vgMiWmrGNNw2XUZjX7iT9lD/1jG4YFzwyDiVQx
BxrvDYVuDQBQRI8Q7eRskQ6PKsNyelvh8iIBoleY4gfX/rNZz3WUAatwLh3kpHjm
NGtSF0bZp9UWajRyhRtcfkiMYjjC4j9tHsKl/+LwcOo973NjlQVN5US7TiuhevEN
xVCBSLSnRJ2+i139Loufv/N2wpB9Hnm5lfNDxDrbxerR7VyIq17E1KEZxtgfo8rM
4WW1Mc/La1NgShY4SLHvrMHNK7yiX6ig8e4nDeJUTJCMIUqPSGt/ekG8jSEpUzlR
f1xIH5loTJ0POB5uTmdqSt/opMsEhgIHPz2AO87pRNQXSnp0SaNM0/oJSjHi8WGD
ie+YdOWoEPdES8ZJtryT94+s05kY+LU8BnvDcCuIMVvw4WPn7EI03lrBtMhbNJVg
s0ItMI6VuXXwMzRBq1l0ZOk/2kOBCnYMsaB6OMtVCU07e/eZQtPmcJxuv8e+ezdu
xbj3L+zYSJF2qUGRtVTVKbmsGuGOBwvL4o6idkHWR157sTuOwRNX8Qm0AqcVUhgp
dgue9DhdEpc4JxRKngyEWBTrgiRAWaW+jY/FhhCZ5cc7F6AiRWUd27H/TKIGrTIG
RFHGnfJ/11rsAEasADJaOnFUxW2IQEzRWHNnrXgM2phOp/MnFGu1L6sofbdGhJTz
ho/AaoxcUjwyOu0QLY+g4e921A53FGQkMzjY9fN1ekp1SGJ2GVZYy4CZ5p75KFsc
eHdZhdsyaXUTPTIFtg5r12RTWm/CmLR5ivVr5kMgaKgwUrAjiqrt18ffH9HdqdxE
acu4ewQSm7sCOqW+4B2+s2FzAXIyJGiP5dSB8tF0mvjFr3OSVl8U2vMpmjjpeahY
8XOYWIFsAWC3nFSfrB1/pT23kiybnrsmumWIfIUklxJKe7gphjuhAyO5EKcTRYbc
5cYgXs0jEl4O7AfCQxLaIEMDVclf1bcCKBermakkFWFkhRjzFSW4lAf5NF+c9Ci5
MbJ4FZf6fT54UYpMNkqdbG0DCbCFyDSGMpL/8c4xoutXJNdvZqjxPSvH9JNH77Av
BnGaTAp3Xolmv/LEsiubqtYKl/heqKWKlw/xVQ6Gka5rZ/M4Exq6IETOnqnWd6VV
b8fwOI8hTYirAEPqXbQK9q41bw0ymnWZcJwoKipudS9VR0vV28SPLwPxGF4Ucyhq
xVNsyExO1k4B7MgabF4ePf4GNWMyRm1qdnnlV9zPUhz7osd7Qlm1g850WdESf7yi
Lv+FEeF/IE27pl9trPt2XMaEONeNNKDvsMQSD8hFjL+AioGZBQuuJKhXO7hFTYZ1
cYH0rBCnANQb+F/Px/zYs1X9m+Aa3MBi0avQx1XNzXfYzujHPPPEuehpKd24OGbR
hzoTztusGyJfJfFlnwbtN+0YcmpFBukgYE6wtrtImKt//bCg3Xbk5v3zSk6yTKk9
7mpae7G0vPyqALhMorxgHhEtQ9g4bCZUX90J6v24JmX1JYxW4tOz43Ff+5j5vr8j
wd+P+DjpSfP91EI3uqdRLWkBfGGCrsxAc+wfAnm0NN7P2OeoaKOmpdNx1J7B6WTz
Zk7NCPlPocVyMR4FTRxxtQTq8xhIWj8oViJxRIk8q1bn1G0V+27DjQUe3HzXOVZp
bZuxN+OI3THhuc59jwAaJe9ew7/q2Trzt2+ROrJvuNRk9lD+GxzsGlHII/CdaUxS
k7zbFpfWQ22eoC4w3x/iMwNz7mTkSOK4YxbpWPswCf/StaPzcmdDfISeLFvbPaU7
vYPvkyfu+JGVCwdyW75SWHBf4SxYNB2YQVGPjBmSBh8JPpg4FywB74EsCw4INfDp
Ahd0QNiEtKyi4hHvFul0/TYt9ugZkSfGueLbsRCc6pR+yMlZwlHKgbZpw4vs8ZoQ
l7AsS19PHJMF0U6XjW4bnc5sCLQpHxWl0w7SgfjPoQCVUKOw9B/DaI12fXMb7HTM
0h3B1L19oMuYMRa138GWcZ2yDDoua28uMsmi+3knAPFIw1CqFl6ASYvm0Ay6QsXG
hts6dUWbExVF8J4fx40sJhJpAnMIVisEgeTkjQvLL9mHaJwTgY5EbhUgEr43LtJL
QABRcGVEcsmV0ysw6HNZ14afeAPfhVUeJelH//VGPwKeE5qmr+fNo39G0CyGYiv4
23bCULcQ25vFzm3LQwBYTsl8qYtYnf/Uhw/GpcuTEhJ/uHn4tnjgYScrtsUwbt4k
QfpqIFCbdHALOWrkHaIJIktG2Nqw3rHTm2VOlDNrxb3ipaQCPlCw9fwBksiGVU6o
YD34a/N7zfiMIRo12yviuVtxa2ZChGMbrVCCzMiOTHDPIorjq79RRyOXxyPqxdhi
RzDsV0rRzRDyaUmbgDh4NiUnTElfQtc/yB0utiW1mq7zWLX2WpflaLgbe1nekDog
gfzVBk/8evhbb2zjL3eduy8sdlQz8i0h1D2nLPnYSMI=
`protect END_PROTECTED
