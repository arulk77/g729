`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42hthBvXYzI04Scfq538b3W77AlNDWVkdm4b5GXjVScJ
I2kTU82zUF3jeRDyNuf25KbOdCRhqhN59mgUuy+92P/Pt9CeP6QCEmS6k3V0+KxA
mQA00oT62n8JSK+as+Mk50L3BsRhk0GLJEn9u2vO+FqGbfBLwRAkAv9RPa8XJanS
MBlGY4HIlamNeH8ZIQnFsQUTvmdxh8lle9mvx7IthEe3X032ys4l94P70tKuUqRt
epcCE/6tBzTxj6otrqs3d11tALNKoTWCP+L1rX0JLiIyDyoeRAZJ9ohJtPqoX+Mm
66nft7r7OuESWgcaF02ymRMJiSFE+H3bwYz9Pr51YIijJUNZXc4ZsHH20o4AzEla
A8vZwA9jJYZSpR9GeaC/lswDvpDcjHQiM9V5gK+B0/uBVmvBmjwXxDUYT4VaEUwa
v7gNVInLZ2enYBSxHdQJro9+HtXOc2OXVRX5Ncd3RVfJ4PIF0i9E5WCFuAEhzE7K
`protect END_PROTECTED
