`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46RhFQnzlYIAQvC5dm5pcbzBVUpJQfsAfsaIo8vIF412
LPRsIXyVOv8Fz/s/Sh2vI3919fwkEgd+yP7JTXIPDHO3pi7qKY9gQUnEmZccH8hs
MQfCE8M908ggraVq3U1OIw7t5BopTuiCPjDiDRb1ystCK1T2IIz1TqAajSj8u1fh
fBv8DOHpq/0wbAY7HvI3+0dnOqVv8U2DuJiLA6g4cHwqqJAIZAKgBxauLBsjGIcy
kBNye0C1gdZQgBMLoCC5WXQdf+i06rUGjQ3qvHeCy8q8pJiaVVoO3N6LfDyhVN/M
Bo0Y4ZwO1H8+aRcH51QCeNHLSCp0RZsktrKte64YcaGhuU75LG6RtT9Cca49mEIF
QvXTxVzl5FRroAaxhfJsdg==
`protect END_PROTECTED
