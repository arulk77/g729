`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHxpDtaFUPQl2/UZDQLKemCEgprefsLdZ5BJAjzAf9wF
1qP9CqiiALijkoPj3jbrIRkZNqTjKZ08nKc3Xu9zkywDatgXsgkIkRIYLy8S9VhH
pE+50mGXDkCaJb34tEeD76reRdnuk29rCGX2pEJLkQ8gEQJ++fkabhvTlP9uMjaH
HQAfiFADLlOScnM7ALlqwIsTPyeOSVsn90fPYciFiYkBMydGyUWfCtjbbeUUtNmg
/tOoXN+SMY1wyI9J0d3ynByDoa4US/dES3bjUcrfEYrdNg7W77GREGSl58LPuZFH
rQZtXYUmyR5WVE1Iel0Rl1A1nAJNj/jvJcnqpjaLpiM3Y64EgWn0x938/impYaSo
oiDabwpExfn0t8UhhBeI5EcHdC0kXt1RcdZtMnWAS2842OjIr/zzPxRxK4ck8wzf
tvGyR7jbWkt9X3sb96gFJtF5W35Ekzp7kVJ5ga4y3wI7oWCUfzy4jo+e874Qz8hp
+njRi1GibpYNoSvfpnOannHJtGyh8mkXnENVhlAB3AODR/WxUywCCEXVsNEuZilw
ZbLRKqtLQKpZ5Wb0limIKi7GK2n7eOGbuUvL+eLyuTU=
`protect END_PROTECTED
