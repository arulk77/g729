`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLtReqIvB6TAR+QWdZcyZdK2ubmHSmQpdDSiOnqkZ2Kr
AqqAyyWSUYFG1e7h9BM6a/9+aahFiwP+xPjB7GlweJ4DHCy7scl4QSkndPnlfEsX
NdajMPy7WSspN9UPGWblfcdhWL6cxtW/9BtrsfcrhCFplQMzJfC/6TmtRs5lNhtn
`protect END_PROTECTED
