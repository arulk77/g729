`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
M96dk34m/wQzXRRTfb4UKgk/BjpcF14YlyGmj/wJmZJITxhPW1uXoKLMO3wD87iw
is0F35tdnegYx7WgIUy+ogIhtDWGfgg+fuhY6OAJWMhe52JFRu+e2gwxfD6KdlQ+
puCdCFZ2vHJQRhdS4xCu2ZsLhgMIGl6tVCosNU/OgLZfbcQII6uFUV2sSyduFkHT
3muw6DT1g/gw0WW59Ct1HxOQ9skGeayz45vC3ATlp+38mT6EOGjrZIB00WmXzpI4
nEoc4Wwj3Yq9LQHckbWga/XXZgTAEVAINf5IfAH4fEkr+GwIvYuiNNUDsdpZ/tt1
jeDXmM1gqjaDp0gcpLackJ6fCZDyRqzyZptMKWm7JBBQnDFUTxb+l8cCJHnhh7m9
24LDFVLGkYtE+0DC+IgmOeRRNwbIQd2izFuhAWkRPJkzus6G0AE2rDN3EwAhj1ZL
R5mSXQ34BTFD3geuRFT1EjwDjDc7fpDRcmFIFUAsH5QIPpNv+siZ3vSF53TZfa6Z
ZS2aLVFRI6yYV2qWHcsmmS7cH/J9Y2FAYEwZAQ03x4LsNdw+LoTpxapJXajXtEXQ
jB0Wn+DO1Ru0KHlSUpaxeyFqPVbE1P/BOzLbCZ21EomRPf1Cul8vaoZOzuOCgh02
gxMWYkrSEA3FqnV6+5u0h7iuFW+rP94Hwo9vHSzxgeE9yuS+wnzrwfGx89kMBszy
R67OVkKHH1svYoMAmRB/wEZjU9KXqmfBB1TXoYMI8QZPpg7gjzGdw7YMlgLJ3uNq
ZomABZV7rQim7rQD7rOLSQ/mzi8+1GjtzFWqM9r1fR3IMVpLBy//K2TXXtlJyufI
frT7Fjcg+9oiGft6zgmum7dpBh3Ug59998892L2unB3KFduxJOnBon8hKQDkOPso
EclSDap9M9sVTC8uIC2tWlKvb6isRcvU8PcRuOtwxv2nZmcYhd5Cf7w+E1TT7M7r
nr1T08XBm/4pnEl/cFQjkG4sRouYSlXILKvfosf9uSpT9FVORECugCc6wN+QQb0q
`protect END_PROTECTED
