`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJxWtKwYJZql98BIYeeLfemDZrZ51Knze48JNC9s1cxd
4tHAoWu/6opNNJ15GOVB8QbFJD+TfghLyOsI8JGFZhCBc1gFLziAw4FeVPbsJmA4
SQvb/NzCyXP+yVqSZ9rIU3TspbnPuzUBip4P7SOv0agQ2tA05gGZ7xcMdo819ZDS
ExWCBsN524YrKLa+DCvu6Q==
`protect END_PROTECTED
