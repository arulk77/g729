`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
d6ikNxCuFadzxp1pEkL0Tj/X/ZlxUnvn9Tp3B9rrkYX+D1v0jSZPIlztU6o9ER0x
QEGSUbepY5CVoT5+7XM7m8J2jHwwH5yAu0Jm4jGAiI9u61xHubsJPtuqstLoYM7s
yUAKgJZ3fpSYzlNi9TQAVYc/04gEg4ZetKtr6JizYmHyHSRre8eM9XcGovcdt5cr
EYb3LucGHnNQTW2v4mt8mX30Fsy3LnSzrKMyfi9b2TwPzEhvEZWKkZbp/eH0dOuh
hoHECuU1rgOgoVBYQxBp3z4kn3MatW9M5npuLF0BUnHPhPRa0G0HeBKmFskB+3HW
guZH2NxMul7wRoX/3vjrtC9N8sVa1+GKlSIPlnKsVKJ1Bt2DAUYAuxA7aiNeRGZA
G29Igdpcd1CWym5EC2GMKn2zcdeJEnIoMiUH4UqHItDlH1Bmx5FizRHaiJZ3APvv
`protect END_PROTECTED
