`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4ymLsRGrr96zZa5hzbTJD+AmbKbLfj84H/QJR4CViuPL
DRKFuJwbltH9GBfSo8ZsAeyPPRnplDJEvaedKjTKmOB2RqjIh0uOTNEn+ZlY+z/L
QRP4HVTSTeablpVsM/VpTEDowjLekjXafyHnMin4ipFS0oIk/ccFN2QypV5VVejl
/iQsBRkSYwQlO7bGiyPfea2KLSU9HrhZO9v23o7rfwANLob4zfSGMgtKFTwck16x
gXtmg1niyDJUtWCSg8tEbbI7AIzrGpazHjR8D6y8bouOMxrCc19BHODiJseyLpkr
H2AB5XWp6tbs1jFTvrShqjmuRhPB1oTxM9PYW09d3D9VyLGdeP08mJJOWves/j5W
UXz5sJOhRS/5EkyNPb6vWg==
`protect END_PROTECTED
