`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJyQgJEca1A49YlHo0bmtvUwx5xg1yiNZM0uysSjLTu2
MR15cMkrcAi6/cqHTPKbBwBg6Mtcl3MmXB3okOR0vdIIUdHUXMMunw6dpOG18Bkp
/RR0bLm6ywGoztH6D0DwCjIvfHxj6io28ZNrQCRSi6ZYfTNjYX3SaTSfuhCxgPWR
rAbnBfq7BvpoKv63lqu/ayppXskrcBY298mEXklHBRWB9s5slriNYQyUq7x26O6S
sbzVmXQcAim7ZNidyTtTsMm2oO1Rw5nM3AAFqbmZGcU4PTpQBhaSf0MLmwvywZR7
pzj9Zx2g+rX5ms7qO4ZdchJJGFPIDqZ09el+mzHxmvYY19YHPwH1KYfxGloJCipK
KthPdUhZROXFdUXUODH/7g==
`protect END_PROTECTED
