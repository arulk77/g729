`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
qG51CK73IlnTWC1No8AfNr90Ypoh9o4EVjalmFB7tQvPoImbJaXjPg0nSH/kHeXy
OQz/ZE4tc0EnJqzZpX5FwkltIxfps2ql/sPoOFWfOWRtDin0loKJCXm6FtZAXcW5
7UeWJuTIGhUIffZWh836HF4pHPjeOYu0SzlLMxFfvxTeu/0mC/tccIgGL+yHacsl
ypXDK3E4AS5a23MG80XwCAVeFsK23KriU+d91pcAGK/8ju36lLhFvtt7uMIgfi+c
QBn1f24KVAqb+emqWG1oQaVKsas74rzDgU8TSDM2DnAg0OJiwLT/cVuudEDcSQL8
8mSisTQsv0jkqhob6ciXHp8ScbMH27kXOcNsvkpp5o0=
`protect END_PROTECTED
