`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
uWs4fhNGDVQG3C0tDfp14921k3VNTxqnXS+Q3Exkznr2auYMQFDijiJdllDEnThV
WxWxJ+IqY7F5lpeUUa4Ql8Y1GG16WH/55tu8IXlNU7HCLK1nS4iBHvQMTG5yhWMI
ZKX4EnMHk3u1rBjM/F7yBFdIHndrzN3LQBrwbFr8Ac8pQXWt+X5YmLD60C0Jtear
+bVpS3mB0edOja3HWYlcx7mZBJFFUGQ4h14r0oR24iiwj64srOYvXi4iKbGDcF8J
83Y+zc9wn/8gvFv3JskbJ//96dwCnmkpwHrfqL+5CyNN6bOwuHhG0cfqEgmdaxcO
fy2yWKJQORCUiU/dK2emdI+isOvFz0cEvZ+x7qKmbEk=
`protect END_PROTECTED
