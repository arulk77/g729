`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN74iNPQtCAJqpkkODSCOX41DYq/72M729pAlF+Bn7AhS
7Fg0zduDNnQbbcxgQNKPqqZUEjaHdYCqjQN9XT0ojYmd/4cFR8mulIPrmmX91W2L
n2myCCoMKOK8hPguCtnszTtAshHMwQ/D7VHJ5Jz9+gLSOdA+yq8v2s2KZtgkz/U1
tcAWE1lhfMzpSomoxJxTpbnkajBJceHeHN1rlfTGnTEXfDyfJ1XeltNKkfJIijWb
Nye+pU1LlQ1weO6YRfx8s9t4n2InwkVaRQLnyrEqQHrL1AeisDsZvjNZr552j9qT
osJBVcMSoVaLwzoZ6L+h5bBGBsSHjaLcHOkw/Ghd/G9epXsVhQoKsWd6VsdFyGLi
1VDfSLev1czqdNCb0e5lj0zLtCKQZvxCamoVFzuno42KNLXQWXLehwHhP7L9dohU
LawAHGrdloHaIr8QSLshbfoN67e3dqGkYYxKZPjQP4QkFEuCnyOrA1qUcYdtO/KO
iiZns9VbP78dfAdOz1biuH1ZV3J+Wz6+mkkgfGDt+4eVf6s4L2uWAt5UjUZVXR/n
K8T4+gTQy/tsUAf7zaMXMCop+k55rUR4NF30Xt9UCWBR1v0oV554QYlEJ2/WZoHE
FTDs5svaI3EuTNZoacoLNVB3amXe2tz0QdCA07itOaSk/MS8Gqf3LVv00UXB7ad8
l0RArC/RYNU+HJKs9vPgPxcuyJB1pL2Hm1x8vsesCyqk/kvEtKT2qQev2Ek0mZ8F
VKFg8mBO3sZOL+XmAJ7X7j1GvgjJtNtiHxq9Jb4RyVM9tJWRmtbLsejvdx9Dl3hA
vM1xEld8XS3FXM2z+NTnxJu5OF+RDYY+CrCFPzUznRv1jw35YaGVx3XROtV4u52A
+Qf7w+lcpMzRQTiOf1bXdaNWI/oDVVdygr1zGC4zZ12wRp6GREJf+B7pjrz/PTyU
22zo88tL8QPdwyTxRfPI1g==
`protect END_PROTECTED
