`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEHaERZb0Bzks2a0Are+fiqAcvf1C67cqFxnI8eJbgL1
+BBIRhtN1QA08+XiBgzd5xWkACZyAjerJqb0MHt34wfJtnRqaicB1rp7PhH3OJY7
EyF2WUs2IjuIn+A/6//4URBx8j5Iz61U1yjnjCuYGJGL9q9ElB5JY/hr1ladz6Ci
zNNbo3cfaQux0Qzuu5Ud3hXsi79mbQq8eSkfD89mnK1k9cs82a+rT920nJEc2oV0
`protect END_PROTECTED
