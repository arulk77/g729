`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAfUX2qVRHS6kha3sSvDGx7ZmHE/OV5MKhawt/7LCb1gD
h5f4lYp7toi0xWYsA2n9Gbdd/ooYFjONrvMa42El6YK3U9Da7mr1b5YTBfDVW461
JMB0btrA57+i6A0iI69M1izqECpJlfIpSJwGDFYoBt1s59vORjEIXtfE4iqvxy/Y
1LmuQ/oiNzO1dfd6chw5loB9FLgi+2qzKeEfcnrqp12LQFoGpixe3gValQ/0sFLz
QcCjmzME3kzD9/rVjPGjdYTCRhMIiS//6ajAdMYMGYH8apiFxoYkGgACNFZjLlao
uCxugq4P5Ni1KlvAAah/uyrgVBGzin7IWnAjkMrFju2D8nBfjH0XQJyj3KmvRnf9
i0UjaCkb2sG+zz8OEgtM3+nrw/8D96QATJfLEaMSluf5NP7QPwOArllxcyvo/d1u
ofmWPPOaPxSVVP8omx3qWqpzXjZdWmG5gkK/kX1qi3jM/+oj11a8y1hfZTBDFn3X
3SozJIHP7+i895s64lJV4zd7omSN8+lFJ0X4lpREpNcCjcgCD806103ZatlyQcVK
pdv0OzrAW4/jXiwPyqa0rai9uVlI9V/RWJzz3F2w93bUJ4ebRxn7nQy+MQ1ev2Af
J8AqTmZqS4rmMHP8yAwh7FCMiPErYkitSHDIVm8bglt+RjdCQsx1L8dNHHe5f8/E
a0gTjEHkeTmPnkQTAAPewDJTvJsJkS7ozHN13omRadNVXOznvvEdJtgIoP+sSXYv
Va/vG0bMG84ulspiYetj9wAiu8msbqWIStgMiYt9dW8c22xIuuoldT3hnbFe6O1D
ysZUO5zjxzfnFAhqxR5lWSZbjhEJ3ok+U2D577U5ZVbgQWLBrYeL9urhL1xIUhNe
FM3lEtp4B3nuICbO74CgYGch2LjtIWx2hVQNKdmgZKzwf4BodsaUP6hjKUCTIFmU
bZjae9oFxvE5m3Xz96+0zfinyWmdIp2unr7+SMgkQeE/K3tPTwHw/L1c3aUYeFMF
xoAPjx6GgEqFQjlbIEkmcmifjfoh5ADTcCNXKTloZpoULwYbyW2TnfBskVj+n7Vp
KdcsqXvRlT3L5CcWKPtaJBcdNDfl3xX5YyCfvzDRM6lGjiogvT0MBFEWwbL1IVLb
+nJogqyz1p9jrDn4mtJaKihhTvqt4aklR499Htqdt4kg/5eklotKO2XBXI7zIE/t
K2jOpGFF8xaYQCwhCafky+trd2BSgHGu+ackwWE9FA/7D+0oxjJH2kIXF5mfnPUp
e4EA2ryQmphlKuAKDzvDotYj5vYNbhQjyUN2HwefuT96XrBpFXHLaXjqG50KG4y6
HUMo4UyYFqjzyyNOM9a/R/2n1CoWaSCa7bX5vlNHOXXtje28xCZMwuCmoEWtNb5P
X2j2HeNWK7IicY4dEBvEDb1dmu7+Zu4PSDVOP3yD2bDOEYm8tSzZuH26GLXqS3gz
iQanARVPFwtlPwpSj6fbSrRmA3QE+Ww/IwstsWVnd2kLAIwlSxH+w29d1vWpFPI5
iw38MNnet9cwA1S1eFSPD8UjwLKZXSzrSfmIbDJ4x+3Hd6SeQLZP+/IghzHIjcgZ
7/+5e/fBuwHGSYmAMzyGiw==
`protect END_PROTECTED
