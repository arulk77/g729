`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKH3KXAVZ3KAPBd2DonA9AmAhlq3tzCzoCDsET0+RStJ
AM0kCjUtVex/6GvEUST0sQ8KoNtuwDw/2mHAsqVUZyGPAJWPLnwedEy9X77k9ca6
iODmVinwSTY53ODS+XuxqmQ1mPOyaRnFC01fRs6L9CX/0j/nQxIOF7yUyD45UNOq
XEYA1RBhjx2aOiUFrvdh8LxLFCONlC30aJS241VOyuRd1KDjyKDMb22Wm5DtCTvH
`protect END_PROTECTED
