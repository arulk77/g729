`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IUPb0nku1fkhXru66Y7Vf+Ze/zwh2VCuVi5z6FYvV0l5IdoLllcehWcPVlC1l8y6
n63Wpx9fdzR6LNuXfmTZv2lf/oxpZoJFUUecnML/WNiQtljxYU9gl3tCScsYjc2u
zmDLK5QlMayC1BD0mXGhckAKg3IAWW8XzPJpZR+l6llpC0hKg2MQ8uBjqZvHCl60
UBICcRQy3cC+QDbvWrgf4zsI8riChIOIbCW/c/rA2pES8gcByalmfI1iQ67iGW0T
nh3uMT1UiqWdU2Gvxiek7RQQnIvl2bW4KT1fowZTpuIb9y9ZU5oELEEQgiOCFz9d
RZHGflX0RovmRfik60chdc8KXm2xjRonP0Z5CdFSmwU=
`protect END_PROTECTED
