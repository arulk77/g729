`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aXAs7Gg/Va9YZoI0W4ebws1JvUuoPMa2r5dxv23W3Jk6
vN+DrbpIRtrFvLBl0GOHgchT8vLfX5okLkbu7rvjfSiZ1EgwwRSFGshtojysok0I
dDQhEofsOI50se6bAoK6XwL55V7Q00mSiDQVWQzf0GgMcfLadb09FAEAPqcLbSz8
qrtqHr7DiUeASmqfdfJ+nKFsRw2h0oSKqZU4dxuqtic5rqGJgpk+9U2GRtn6BhAV
mD8E5//n/qjTVhSkGI2UqhsJTYaY+zGZfW1N3RlDERqFvehLt/tZTHyC5HPhzAQ0
z/40M+N0rCaiVlIgrA5oMDilwd8lMZDkRJ9z91y/ybd4z8pRyFierW3jnVhAw4CT
EOQMRd3ZFoKv5JsEt3qglW97bz22oIcYJNscEX3OcJ+3GgvcwSud0NR2y8XL/Dc3
gFRPf+YZSdJ9GMFydoN5UABXrDRIMNF4tJnOTrFGSvR6UpraVOttP1fJ1sBiIr8x
E48Tq4jcTeqghACAjBxzWErSTVGlKtQg9qGMeJPSAgLBgZYz4KN2EGRdQ+kfLhGN
GgMv8EA6t5Yohgrtm+mLAVz6FpsHozBZbxHnFMVQiD3/eHeXkBCaoePPqxRJoEqE
2sPMGLbUomsD+0/UxL8esHbr5Cx156J+fpJNRr7Y3Sq9n2YD4mxbQ8TfJQvEWrDz
QT6dHZTyPiJm8y3v1wfzQ7CsFzzl6ZDd9vPVdsZX+AgTQmh9ZjSFo0rXZcnX0KCD
7ZZxXEiPQf/MenSJiReOoz+/grjHZYBBWLTg/FYGpy3//pkfA8QInZPdbilumBlm
ZGuwqKhprIqRQYApzlwS+/BDUXtsR6pdckL3JIwZtF17sMQjuWpmBkeeqoOz8SVz
vDu6OrIW0UnY+l7v4d/xfGPVw14+LkdjHa9dpYWLN9/QdtnXW0od3plTJu/r1yZe
uZ/pUC1PMtPgcQBzEMUqUf1jjnhimiXbzBBe/T/Xjg9yVXL0IRuLxR0KOrWmTjeg
m19mwwNgw5ClsndedjANV4aZSBDw3PK6kPH6szuVz/yjOVx1nnkKjSccsYGdwqwm
FWhXOaG3cX4gewvnx0lfhIEMRH5SfovJLm4dP1TXCQadrpNyfuEaNgtGbkWAgdKr
utmdIEUsSjZA6I9s6XPwsKNB/4trA/shHD4OEzn3UpvgvuRE6u7oRt9K4NUScbfT
SllUmEnmwq13/jsjWRPzJfzxO3Fyl/BzpwfG/DHW+SI07/ioCQSMwtlWv7/ZiAOf
NbmUOIDAQaguElA5ivZRBNPfhbjZSdktDflXkKK97mB1fzeyh3YhLaFoF45ZwVVF
hYP1avjcn978xpUXjUaOE5D0uexB/8B3n5+Ki6lgXVfAVi6hJdj2w9nUsgb7KTgo
I4+sEfAzsx86srJpwbUPTW8e6km3fEQ1FpGfEdjwN1e0T6Su1z9ugqZg5OKMVel6
w2I/Gzff8Z2AOZBWnRE9EbEGQ+1HIKdPo2iEbH0DHv0zVHfTFDxkQ7SiOJuE6Pxv
ZKKgGymGGZ3g6SVrhKB3zMpYl5Fm+Tx1NkbQxeGzN4UvRbX1aHfCbYUc8b+ModYG
d8b0Y+bJgoQkMxSkfGRV+PAG/ApPDdxii0Iv85Q56nckfm2OxnIiqucQVxiJNwbC
O4zQ2Gn5IIyxTv1YZEBF1jp93bU3Hz7PsmLy72EZWnld48y0Rb+KTE+WlLOv7T3L
D75550ItdZ5AN7BVc8e2XKDew9qFKOeAS60Csa2RnqR4KgtDQUBXgdziRT64B8t9
KJZMjGjKFaQ/KNf15hcZjBJi7u3o4s/U65komzUnbyiSLRS/isw74VrMFlA2Wwh7
WZ4SqSGoI3FIPSJb5yElRwwmPzgjKdsRHBY2O/+1laLwcYk+4rkN5ZLuz//kr7Js
dnSequyNzx2b9Bx1mmYmjttptymKcxlGLEeWiasn7AYv6gZ4XXlXuzhqxbWEU9hk
D0cMe+l1j27MyEnKGa4iQfeOuEDfO1Pb9JhmNnu9Dj1eKjcYdF3Xv68Xsn/cN6sQ
+k55zz7WHH8oSgA0wd28XjNoSkLueQqgPr6cldrZXuQz3WEYsm4vkqfhmrok9cEo
lV+Eydx6ZCVKm2RmRegSJXU4SyJQO4J5oXUEcIf/xyZvsRafSfucI8OnnVrSyqVP
sGIFXv3VgwuNHLciSNxq4fpT97dS4n5GEYIvMLmTGHsvUZYKKsPsOYBusQmafm6G
ZWgW9uXy2N+YNz1X0PxrpHwVhK8afR85BCLqFVeZe6JjapJlKR1vn47GUB6ApevI
XEP4oIZ20DKQjY6HvuqfMbpVsRZHyia0FD4Up/v5uuR7C7PVOKMToYwWiYzURpLy
ldU5mToL18sacf+FFI0mPBAHMK6iLIwSdqKVLpAaH4CqoixZVZeSi3vqaTcvjXha
mgBZA1Fg/9etvzclS/LZ52Z++XO9/C8CDDKuI4DS7Qp/7g3/ic7ST45wPJY83b9C
uSEJ/J3N+08WiUltip2DT+YRAvXa4g+L3jUKo+1/h882IMdVwvLvEU5KKAUF/YNq
z/5KEZCA+CQs1V8xWo5lnL5xeB1ttNLnWnEzDG2EaqKsZo9Omn3FHBJM1o5OrxHq
cyQA1OuFshu93s2xpZ944kJP5KcgzVUCIndoD1ljh6I7U1seA8ytuWRAl4mHdByP
Lk/cCaEoGjgnnZv/l5WXxi9d9Z5Sex2GaHmIQZkcvQBSvmwmTzRAyvU2R2ttTAQ1
JeXqba4wEGjLj+wROZa5IlyroF96mTOdm+HpWBSBnjPErxwm0TUFeHmQa5K2PyPV
TEUu+wnnbPTHt8c4jlBKm/eLDzwC9a9MeWqB4wWu74d+zKhlsn4vDdhoyCVShYBR
FWsuMSDVL1BJV/CgCVi4ufZAZ2XSNYzs7HO8ZfT4kO9g3qhRFew/HZUkmjiFnNiy
arK+KAuWt34q8OuXbM1aJe2nYCuCxpmV3ySQWMMtogTJemwcZV2MqsTIMP761Buq
lhbxMV+exmpJ4hX25ORxv7Mx+HHwAL3PRboZIHLz6ySZY14Sr8IgK0FUiW79ou25
f9ya1Ig6V2P7iqIXS5Qe/X+hjF6a3CdW2Qmue3taxM4jCPOlGihBBpbCJu7u2VD8
tpVxdr75PaZbNpSWYv0MAV92X1K2UFsqZxE7Ui8x6mgSqOAXuoCIj8aSa2x7OnOs
YYH4jEvp4sfY+VIQnqFxu7qCEXw2xP5xx5ANS0ZIkmDWxk7I9uiXSEzkTECmcbWy
LMf4qjo5Rz6xQnuvAlBsGSVfaxinR92Et66SqZqdyvpPzHH5vm3GXVYqRLomkhY/
N2SBYEUcVTDPXV2fre895WA1S2YBqWxgYhbxhX/WusOTkcEzatMevdIZjovOHi8S
gg0Qga+Nt9nuStyEZ/THh263OFYWwy+uPRbFqvb4UEo3k6SS1KFuY1PlpgcTs+An
5n9xn1y1z2ygpVNK27wxORe5Q6Lwv7WmBtuJmy6w6z5Q/YcHUwY9owj+c3AiFZsa
8odp1/NT6yY6LOYPILG4kulUArt1jwZVQYLpSS1q6s2N2zzn0D+ZDeNywEX/AaX5
G5Fe4PmSylvdGDvgiiCrtvFgKTBRo8E3hbM1xCrBEP//igxo9gxmNYayfD/Z8riv
EsyYt4RcHScme/ZHU8xxq4O6iK27fKy+yXU4nypjsXaiY+cLch+iM1NP5LzYDqPm
aYcNdGIE7iw1ex/ABCioePoWx6qYRa/CsnrR1KwPd2ti8VMVlyXfeCTvCZEM2j7G
7dSPoN8R0rmKzOuICSgRYm1ATz7q1ZDFf4/Lw8+Yi41s6dIhdw69X8JkweRQEOiI
YEPQpzcnjh/Q6MOXNJJLusD4ORwT0ThWYtengji9SONC4DR0Xi8KW2E7xnIWbGQy
6sKT1XTXjlmjAII1OcFndtoUnYNlD85gV2km69s+Ww93ueH/0GIZh4cJATLsIPBY
0H1GVAyy9vgYZCh5CRvW2mU6FsHlHMlzcq4nrRUd1fo8A/5FldYJWkEmAlRaipsy
U6pbH1Ia20k5qYqqZHr31R5z92/4+hIazQqbPvGPhKReeIHnE+To7oN2CqmjDdWj
BuJdipk9/bagbgnGR9nZAr+Ao1z9yjFJPZumia16VkVnz6WzA2h8e7sImcZ53VJT
29JHuSYDlRv2SApvF/vZF1w9eIgBv3wOmMniV9YWii5mc0VGHhaLTl5lomqTklAy
rpQprO8dt88o6Ilz1b/xXQ==
`protect END_PROTECTED
