`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2al9Q9ZzTEACQoO+fa4cKA0idFGlTk/SIiAwIfwklSsfj00VeEWjCvo4FjhFAO1I
V0rwKQ82KGJoAzY2c8hXxS2X16yR97In2EkiZUHkshSTy+D1fiN8GtfmstwynFAh
RFCuF9pbudjcv2BkZ4B9ruYbeq/tQSgT4UhyyPGKIF8a9HBSW7oK7cd1Zxy4NgPk
Wto8kfAKDKezZShdns1iknyKx92c2by/6xAGSunF1MPEMFCTyLGt4MEmmYGTHzDU
Ex1AYEM6H+FyjsizEVqSFU0igdNVNVFQ7UaZeAf94tur69gFnFNfNib77yBjQhkQ
wN+bNKIrKU54bEBSAlZGtRO0/wDyFKWebMa0+XcQ7mEoXInjkjb9K5ts3mFp3nKL
HC6i93BdksUTsinrJZfdewWpzJ9Z5nzPFVIyP3Kb0FSHRpufe7xkVGBvf1Pezlpy
x4U2FX4qHA13rapX4MUk2PEAN9LzG3HK0X8rziPPqR9PMMBZjVWKBd4ewsGuw1Ou
7WAA+Rg/JQ48Pca+3wVRoTG+VBUdljdu78jzJB1UJ/bBUPyv8YE8v3ESiBGQ57GV
FQjez9x9R3wsN725OFJbwQ==
`protect END_PROTECTED
