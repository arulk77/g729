`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+wGL8FIwP5BTgVbQVNJbvFZaoLwSEgZpQ9rWSzDVsz2
ncgo/1bHLzJO7js1WIkk2N0WWpIfHsCu3Cztxh7dtSB6xrLKuGyDOP/9GSDLhX8G
SHDllYsmnOj8Axh3OfUv9T2yQPkI3nRFl65Ot7HxLPcgL7z6dwK1xY9h4DULAzAO
ZW4EKGpRCNWIZHlSJ3KzySJAh6qmlq6AcNpY0yjVkfYm329oBXkSNijJ8+LXEA1w
C3tdc/t+bKZcrZQI7pxLUvBsBAMlISoOETMt8GvbsLS8VjX7wZV53ECwoSEsfYZS
yvnFk5GuoZxiagHlAeGE3g==
`protect END_PROTECTED
