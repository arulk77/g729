`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNAY/X5LqwwnKA6RDo61EduZSvjcrU/ky/BzW1ko6T7g
58oTqUFgv+WqOY3oDSgFfmI1yWHJqrRe3zUB86W4IFODH179IZ6J0iDXDrNMVEe4
cqYv5mjX5WzCMvz9BRT4afrDLk2Py0Jyc/0od2zlnRNIFkFXanNoi89PnBa4EZO5
HGgOwE7l82j+pb5e7Sd7XmZJPtoN3/KwFqiuIKk9vaUsnCEEbzcf8sKsMn2TCLz+
J95ru4IGdojV8HOAMySLGhJHS1Mnscd4vHKIEVUkNT7bfWDv+2GZftPEF/KXMieq
9+53F4mkk621XGsDWyUsO7Hl905BR1WMrs6jnY5id1PavruZcMPGQQdlu7HKsMr1
FmV9QyJos3XDUzVJeKE69VMbIdeBlEO/f0VBQwLsoGLdoPI6oa80BypxfQy3N5gR
lSyTR3jH1Qmgm4UrPlpLbxE/NnJh31FljoQAB0UtSDRTqePjn4sp1/i4Jb7am/Sq
`protect END_PROTECTED
