`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEJl4JwmBurQt5umM4wQ9Q7RprdpPVSh/B3zyJC2ExKF
s1kNAGhSK746eXamB+B5SbnFRobKaXOg91lIj0AKCdlm39Pzt9aP8LV53N9GI1lz
0OaIexiZ5tXbv8ONswppfT7q8g+2xshpvlQoEwFb92KEJoefLCFMN1mHlDR+dAKZ
`protect END_PROTECTED
