`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCQqIQz+aLc56ANnPu57UfJMCr48j0HJ67AifEjB+HjQ
+wmZUpNri6BApNzHrtCZ5Q9EEoohHbAjZ3AOCcBvHxNg9V7UT7SO5Ia1xNpdscs/
t4CGT/3IEdHiRhABg6f9pemvWXRy9BXImbU1lsdOglrjAcyTq7p4aIZFh4ma1yzz
HchXG6yPjeTWXyn1P5kktxvGg1oo617XuQUc21t9MAryvlAPaYLWSkP0zmebdMR+
Q6vHvWFWwqxcUpc7uqc6pg==
`protect END_PROTECTED
