`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBMgBrt49HqaZP0CRhGgfbxoth4rU35f11Ia36jBuRTW
eYtZD8A7HOw7UkIof6JLpGTbDs222MwZnS0Sd36DsWa2BWDX0mJfaFi/NyuqksGz
6I1mm2DvmZXx1SzjphoNfQubWelesCsA/AgXiKNJeeRBY3VkQkFKofFO4EOUlum4
0QsQKX3+0rNk/S/YYMpEW7z+OJezyQKpfxQ4Hg99OG+j4NNlyvVQs/+URJTtAuSZ
dJhdpj30WDIfuMTXBtES9mgDIn5pY15URNhBsjpgxAz40Le5kXlH66daahW/6xzO
vaY2L5UpMvvaTlFc7Ux3G8ovAt2gY8qVgABZ6RbUyd35opKb7z7O6MF/2ItMDZgM
HG3ZMHU4XwXYp8DembSKHA==
`protect END_PROTECTED
