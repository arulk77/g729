`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJw2xCeEkkXs69Z815D5jc0PwsVHBNXxrse612mY41fM
dijs+8q7DNGzYNgRqvCRqzZMFQW/ZXErNA8n0sIIkcvm9YM3/XEZQ0Qd8WexCB+A
mXgFuoKi0BdFVD1kGWR+VRpWitkHOA4uaP7WwjfzWu3VWgz0JvttpSHCTuQLT1F/
/J9dCqMI1QHuYV36G7IO8zWcgEb9JwKXcZRq8EN4qSfMfQQvYh/p9b+sDzV4wsCP
9hXpPdhYpfKI1dKrGJkwDOjAIKuAwdGEViUpp/ElJP7iSSkANa3vabbR1OUGKrsg
A1ItnWNwXeH84goKuEAM18UgaElmIiYwASX2zKGTOrqdN63egvnOTb8BpqsSZwkH
1EF/8wx3QUKKsP4+B6JrgTv2Gpok3h5pdZaynt8ktUvWwlFz+FjBB82pDNt9MNQ5
U2ayhQSWefQrZ25eJVN3p/vsTeuE07biEO9i5fsAnTd9z9UvKi+Wdx19MAMQ0/TU
lFcYFy84loqdEJpdhYUfyTWNHqAkG98Zoj+NldnOdeBAISy7NXtV0yI8plxBPqWO
+WBca9czPeKxVVulN8MKf8CEAm2EW4K36aRALJQi3CER8fLYxJmODBMPRk5yojZB
SgSEWmuZEDpiugK4HB7MJwWCjHjrOCzfQz4cm+YlwB0sND5aFWWQv+ylvJGWXehI
1eSQTMkfRqsgnY9RUYmMEq3Kr6bH0OvfL1iI3lMHRqkf5ag3wINzcT3OWruj+f8f
XZErO8Wh76C9Ygm4Nhp3VGK7/jsH/HTM/6JKxXY1Z3IfESa2YbagkWsNaPwSfzqi
cZeDODuvubW0a98K/5BKS49mvwQeaizv5ie5QbMPiMI=
`protect END_PROTECTED
