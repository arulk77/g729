`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCvvkkyKWJtBqde1YW8zaepUMYBOW3vY3aLWo7HWpBDy
15RdqQiyTwiDmMlPEAcSJ5VVGbq37BihlKV4FFl2SBXJt70+DWdBjhja5T+dBcZT
0O794yao/+Tf3o7embHlfVMhHGTjQKE8LAzxiQ+g1YOyOW19PhsKougtSc7ubM+p
9tfSc6kDbZdnDOPKGQFb6IFJJdhjAmpE8eRSQzAzXmthMxjRkz+J7sEXQrXVp3hw
4nSNDd9INbD3GULygl2+Lx6i7EgfK/0+aFdYYlYKpyonVrLdvL7DG1+CTIZUgTNu
/9woX6EEpi3t3VckFTDR/HHH9KnrVhztkWeWqv/OY6iAHK4btLO6VqQGd/pU0MnW
h+ORMT7RJUSUTRkhi5iwztFC2IRLNAuJlNUH0oM4bzPoPR5UT640OWBdIvj6v4E/
gcLwOlLLQD0qPeekkDbO0oXI+vo9AAvQ1vNKJWErPbOiS87tWxHq3LH+p7BlzN2F
4e32t3Lqiye51FxTp/YYZGxgiOSHRvS2PM6O6zzpT3eXmX2ErRidtSSxhD5tg0d/
RhY0YnFeDpXUDkjJzemdWKEVAAeWu+xaOU3/mu+pFBfBV5sKmBz4iwxGcEiVMlem
IwXRmq4+s5pNawk7/ZoNFaKCIi9rK86lQxOO3qeoXzOwTANmpKsMwPdTB8RCaLUG
Pt2RRW08QcskEM2uyNfJLp/rYYCSQz7PhSYpXF+4cXUpXnz/bpGL5+eecvtjYger
NtKERl8+ZQcjR42lTbfCeqENN30+rdEQcK/bOhuZsdSgqRb3OKTtPaOoEaUWKIBc
9kWiiKig4oNZhzZJ2L1YJ3S2AC3aNus+UBAFqEgPr1g=
`protect END_PROTECTED
