`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAWl43IZCSfuH0fx2br+JSdYgtfV5R30ep9W0IbgxBYF5
+RBvZblWfyUMsg6X+QSLOaCxgnlaIMWK4+P052waShyPFpN3c4E2zlOlmDVDczxY
ME2TqljT9Rf80apqUdMqvFa0QL9rFQD8oGyu1sm9x6DkxqCsehLSVqMyk344V0bu
kX1E9VR4ZNl7jqFnPL5gckIZCc6ZVvZTs4DETQkpB4FXNJyO16cDQDW81qLg0ri9
sBf5M+C43enY0mry4Yd+suKH5/15D6/yD7AntaXpiUqkzmIKrzBNiOvxW0mSeu42
5dCu7abe26sRq5Vs08GmJiX8QjHodBXEvqwl0fOulV1VizoiO6IA/h/6HY5cwHzS
YIQGWQB50CGZPQk5F5o7AXq3/JCRFUkff3TwTt7oJhly7/gGbeWggj5hhiifqLdo
B1Jm8rIkuMyR65zS+0svdzEntDPfFvCniIt/t5Io1+HuoVtJLaPm99dsnJW9zoHf
paiEX7qgZBJvTNnSCo/xoUKoFUBJdCPpNaytzM0YrJIydXF8x0RTOD+MCrH2UIqP
tbUYizqzFJGr2gqwyD4KA9+QKhc6nM+56LER7q7vKmciH4WNB5DupNhK57ijaT0Z
IapDkhYeQH276UNlb8mqKp39s+4frBSZTzhFEvneU2Hl159efAj6MG+HG9xj3QMR
VeaPMLHEvpmxJ4wGYfRhQv2CSTsLhYfqp3tzGZee1uCABNAmSc2CWWQsyZpoRek4
vj7g2sR+/WfYwblbqgKOixy4TwOf07qvTp2x73uzRKuDnN/R75wL+YxciRsS1Xhq
ZrG1dshtGxXLd97YisDox4hjyqAvU2Mtlf8fkvIaET2E0pkdgIfEGPBdmCzZICxE
C3CktfSe6mWwk/3b5OtFcW7x0WMujZNK4hlxHWZ70uzg6QqtXUV6w62iw6+MvY7A
FCsCDIBPLFQGLgPTWCAKNWM+SL/xG6swwPoKp8ONke7xnqA69gqv541sdo9iaU7e
CEiATQ/7gmpmLA6AqF0LaFs/9o4cWatVVChz+dygdlnUJCQFLYuI7F9Mv6Km6eIL
HsvJVjDzVgsnL2f6+DmsMzxOseM3irL2N5DiPNINALs8uUEgXGkGzpsGsYVb8Y7w
6L62R+mtRRgj8lEbF3o6b1f0DHPTCWDIdGitVeZO7cr8BApzUF3R/nCUhpr1RcXk
LfIfck0tfkHO3kKhH9wEcRA6dE98kPloH6pDtsILldtem2xwXbtX7Qq54RR+FB+g
4zf274yguqOXv5EEe6XInxmNnYHX0QAbPHwyWqS4aGZksFcC801VJPhaznDRL7oi
tJER9pYPEtgoSM3UzvnR9YQPwVCcAS9nwtsgxSF4RPAjvBR6Ax488h+eBFh41bZZ
UV7cVUbiWdx+pgmxIzP8sTdwkVj9dXQrkds7mqmFW1COut9OvpP7/g/mc5x4reB6
SHnQCbv3XiP5rs/32YC+gGTfQlynjL2vz8BlVp8d6r9jABGoVqL+L7fDTh9+Mn0H
3iRzS9Qqhd9QbVsyaS/C4hgbDzU7nIdDrogfjEGDdhmBv6t7XLfWsEb1UzAqhnRe
oR+GKqchFATvemH7VCCsq9CelkobSDEf49OZ2b2CpavnoPWIFow9nQHmqCS18gXf
TU7vOqVFR8+0mXD0wIwYMA0DgrpsTvJn7hYj88wmV5CAQ5+/F61KwiWAxKTvyuew
9qKVkdJdhsZSvnWCxm960qjdA5HLyC0KCaGBU6Ivt9vhU12wn7EsBkIKPnAfiMna
jtHqFPzytqnzoeyQMV9buEKgVKGPsFhzVlu/unhIVpvU6exxZG4a6czFALSDWrCH
EKERX8db/Tb6klIdxCWcXH4wOvuXwyx4cvBVn04TZqTjzoXzyn5xCz7rZnuTOSDg
WeWX14AfvA76blX1bCbDK5yHj8Ew/4IdycIH4+p7fH3UuDvHWreE4VxhDWzZHQlh
TjrWD5bDkjZINuPvl1u5RVTXxrSyuqQ/hNJ1gNLfdaPYHVUPGKYCcVh81c+ICGcO
XCvUn1Sjw65LXOFjtwfsRaBe9I02CzfxlNo4/xvSUWFFJVYyi0aUfwL3SFFE6HvM
w9BhFyt+B7ZfD/jAPlJjP8c4TBNTWY9kmjVHzlOxL6MymukvKagiqI/WiocJ6UZG
K24rWcXxj68hZrj0FhgtH6WTGmuhAzZN9a1A8lpBQEiVGXGgw3EXnEPoz4klbagw
cjcBa/Xs7cegQI4dk2ETAQ48Sh/xE/EJS12drTNcYMLA3hefO+OBeYCS8k481I5Z
59mdWVd0vgZgEd0cKI3Q1rJZtAbWRCHpv+D4xSLkkFoii6P3G48oZ0dmioHUCcbD
riPgfxOB3Tks6o0tgWbNtD3TqbLTJKaMLAuaf0Y83tB/xfbTTRn8kiRouyoSMnF3
qq40BXaO+e5nB5X9Z8H4MdZQGQn+PE43dReBenSHLoFx9odVElPhHRtu2wf8G4K3
/UMBIddHPLD3Ptel98xLH1dkLMckSrXszdaeNDnW+N5so0wODIAonkmkXHgkI0gk
dPh5/hQZCrRHT1nX0xqKP9ueV3sPbZWVMLo2qmvdD1QIPx8iujzw8U3SaLLmMKtC
aJr9nY33ehy84+rRibVmbi7XbOSPZvXCKvVYPnGUn+3FfIvASU9A9zo+ySntxx8c
mXhL05mv1m82jRlEct73mFUBcbW8ueUxtkQlatfXGu9+ZLGMdQ/CUUyiTX1sANws
jWzioZRnHMvJtNoU8UOYNSgmnMCKFpFYWEJRNucI8nBThH/Elx8gBKK9jVMJGzNX
SMxOj87lhoEo/+OpfvL+QWW/jp4rwh/T14CzehJPeIVnJGW59T/x6RTYClFWgTud
4bbTRQbfEbbOUVxOV1syW7B9IDdhOVM8K8vTPEvBiLVc3X90f7XdmBtfaxEU0G47
iVGwvrG4aIgt+tD1PI9sF24pS+K38uM2IvIZmrr5ZayYpxA0yGXUlks+EbyyaaLM
Oayzve6aob+p3ZmrOi3upGNVih9JuSaSJbp9Ov7/6lyvj9gDur5WRct1Vk7KSJ8o
J1yJQcIww1tM0M2TEI6Pej/NV/WuCQXwfRwN0kOBuXFiqB/v8gWcSwWRLDVp4Zir
Q/BInp58moZqC2WSbXuVdD6EQ5a3aQzNI76t++YDU5I2Bb011F4+akvEszl6nvm8
Tmyv+mxaIesyoVAYejHnk7JAH+XFn/hm3wvafKZhjSJvmzWAyOqlRWbPI2etMV8h
cEsBmRpOloOyHMp5hJhh/KnV74JrevgBzOurmmYyymoCUa4xGX2BX0qenHESX1iq
jvrEzzvWeTQUsE2X2LkX8I6OYD+GqsW3qiWO8e/D+MxUPzbdcmCNH1T7ES8nFLTa
EAw4L1kZq/bNHzwKfRKlWD2TI/54ENQUvCC31YifZCQQOUfKVMd0lx0sFGIi2JYr
hXOXAhJB8XVGfX1Th/UHQlQhe+siCYtxSWwyHVHpZlNxHjTXMQcFjkCWUZZVme5G
w7jzSE1cR+dj0CClCCzd7xPyvVxKB8dChAS+zQ9W7IeiKC4JrbM1/jP+VlVoBoE5
kauZVN1jvfVSC0INJkTfAZX8VD+UkOK/e1EeKFAPMv2V22ScK+CcBbIaWPYUZKZw
q5/3w70fcc9Jud6BRmUYxsVWUDq9znQ9BOKigAgi5QBwmuZRnhaafvC945YWcPJZ
xUaHN6hFlCNIUB7PVMOFK2/H9vDWHlwdI3KkJHS0VE6zMO8eEG0BJ0FTUhUbgofq
Or96c/KvdwqpDJnPSd/vaW9x/n7a/zKb72iMsABFg2XGwZWYzqye4nx0iWZQmCC7
N68Jd00x01l4Sv8vXfKFwJPLDM6rzSnKQvdjU3aD6oOX2aCHXfOXgmoyP0sIsRYs
L/A5EPthGfdilYhNxJIyWzgfQmivFcMx/KtKdqRmQgPMqGfcuqWmJgJRA8Q6Xf1o
SgnOWcNvbtIjKK/eLubXEnRy2OgjtTdJPJaJZum4urT9GmqIOeO4nj8maG5UxFsi
VCe1FzAUJ/5pxfD2r9tkqr0GgWNTnQfhjBN7aa0lfFZlnpVy7N0DFEB9aHRCOv4J
yNgUZ3BaXhC2JaACi0vKNX5atcuB11mRINlhQkRXzcl5r/5rWEeO5vMbH+IY80SI
Frx11Gy+fsD/iGX/AgSWBBvGzQERvaLpnXbCN1M/cTZm4DF0OFfKmULq/ca5NTMQ
hqbYngsrZvlc+M+dJMC21YaGcn8Ycf9Am77drDz9wqxOIQhx0vLz/I3V2yirVGHR
6KKouE0cVlsw0GNWL3uFQdBSOqmFVF/+BLt5hwk5E/xjiivpEnPMjnoTANSTBcVw
BwJU2XL67kMeQzqxcm1HHTbMe/dxtj/9axBbEO++6yfwOvTfNsh1IiFb7E6GsXK7
vHlEfmuMOpM0GlN+JgSiR3ORgLKBk+YNuVNm0eztD+SPR7QkwubmVE/NDCK2phmI
3f0iGhOJsMjdjNKDskPEi0BSD7gcONNFOYq1ufEkpoFvokBhjenmELOGcW4jenw0
i8WjQo1ruIDDUmTpnc6p5maaUiAr+NFqA0NmK65eiRkipNYPWy0/6/+EaticCLt7
k2Rpp8+iyjQ928usG9RBpJAG58FbbsqyEayDJVkQU8gFCaVUWoZfl6pmm776gJjM
w7J74uWynBxKl2S601LB1xQzg/400aoqCIN3ka512nZCRBy9aFsFwft9G1IeNThJ
sf+OFdB2LuWB79nYonpJ8y5to1J02Yek6E+RkVjYLzILUCmZRwwXks795YxDP2EW
a699O1V50FFfpbiIOjqUQVyQ/8lPDEyyvdJD++3xWEW2FVrf+uUzRNAjmlqAG2wX
uXD8jfDiqTa4NB7alMNuB5lDRWvtXyKnnrRv/8FtVAENq3LoGNw5fcAy7EwIE1zS
IGPN/aAMhTdvQE8PupkKzUVf5AH6o0L7zSvjjO2irLry7hLwQdYIP6vnHL30WzpT
kctCYcVVsxgcdHvVUcqre4THgRtiJywND0vmbMf7uJAII5lm21dDbURqkYa7xMwr
a7gLUNb4lJDua1KP4BFjTkKysslU5l55oEhFzvBvf38Z/DEJJQuseovt7betNIKL
ict14Le8r/tj1Vb/U71caMCjkREn9w5lgDh9CtukM9+U+OxbbH3c+LNbpn9wa1QF
R/f34oR0HhSDiUcDKDCqnAeJTbbl44bTYJJ0ZpEtRL+kfkgeGPsUrSpwKHKo88gk
UqZ3rarOiy6Fe8IiZLgdzV3e21jlh7K3v3UOlCU/qIIy3se+wSK4Y3WuLFpWfSU/
1H9YxBfsGwwOdAAV5BopECaH0VRMQHLNJYc0uSipGF6yJJqcyTZismZ2Z39yVVVQ
XTujQOp7jl1sdkfK996WKlseE4pVqGotCQtW89JdQ7ttt12fGV0wuefipWNZtTnA
GGOgwzGvAPvHumqxiS7Eihw9YSAumIfogw8e89aXh99w0oz8kxhiCe45fgLSxj00
tkH8ToGWEv4ZcbcRrK0EORGT2HfS1Q2yNiJnlnsS9qh2KewOQJCnP2sOxvpdIDNL
IVPMZlAW/QfZbNPeGPJ9/31VON9JMv0nIDPHq3xH+LuzqoG9S4r4oQXhfvExRmqk
ElSF5VLk20D6y+4u5aaKtsVTM6rfHa6iBwzwk9tXDvhsKpdxtTea6MJbW/qxnrGX
zc2gTxlrF17pLDDKtMKdoczHHAh7Cs5ffngFAuFpxAMTMtuGC4j+VUDqQmpem1Iz
AGIeob5j5cQBp9JfCQ+QSWaucPH4HM+70LgTyDT/pUuEZ2gv9GSJPN672K2kcLPT
3OMZbMEsVveVm4JmN0QMXGD3fODKpU2UHgz6u1+9kP/eTugdIfBwqG2JDk9ueJ2t
TpiBKCdnXFKimA8XUv/aZxESBwThpl6+BkHQyocqKoFmE4hlhkfInmhpRCdWnrNT
w8WETAjhXGyQmZdCaw/7d2Ia32KZo5dheKF3lTarZYHsP/fIaCSRYFM4+8d7WiMy
brFLDKJH2+xHtyygBYj4A/zqUgChYzY4S9E4DCtlGS4yn7ynkIeITu9jZ8Hgy8nr
0pAY4ZNKQPSidVJksy9E3skouT35rIJCNWSOzovBQd2/VivS4huJpWYK6Nk5u+Ee
hpCXBDdAOyagkOFVmqJ2xoV96ZEoj8zlAng7HkyKJadvdwUJHymPiweOe3fOLIaQ
tZRHl48MDp/LOCOq+vakW7LRpQlhyJxbqUYVpT0hNpElUyp6luhX7FvJHxRcs6vi
kieQu+L1NN/VVTByVeZLuwz8v0bTzho0/0fr99AjrPnfbXPBiat3UyRg6D9ulY+z
Zhbbg0v3/GHTJLoVyzjFnpTb9zZMKDu8lTy3HrIt0GCEToSIglOCj1/65bTGa415
kfWuh9Ft8WdJZDCZMC2XFQFj1RMdgkn/ErhHimonGslhOPVWSGHWbXbAzpvpIigJ
/LaENWQxyMnrVx7tbo9dFMH5KmhIbhv+9SaeMNcL6p81A4OmOIYoK7Rqn9UZoh1r
lHQjDi3hlbIN3gHUzrvTvvqxutga6x5FeMoucsMKEo3BbVol5smoT1oSBogCTIfa
EqY4JoSONODPlOv4tAgI4ZoQY3f2UKDzyjuh7roCEpLSlTZIZI9bZvT1qNaiUet+
LP6tlRS9UEb/C+m0J/wShnWsDsjU3J1sM6qjZjDKwOb0RmCYCopu/WTNbhPs8xkr
KBwmQFdXxiRGwj0bRMm0HyK5yggGudN3l8QhhW+DmxDpHF9N8rXdv2Kxd7qGNJL6
Bzn5u95E80YtH8cRa/X95lvOwLkPKPtZhZfAQ398NPP6okR1pCxRqD7AKxyIzVv5
AOQzJ1U8Ppam7XbRy3OLoo5ENlpXw7Ajj/waI7CfMhYeBROaqY1jlELEoEMIfaNN
CMhI1uXTeGQWy9hstVk6QCv2D+xuzQZLUujgxwBSslRTU/bXf5jLhyvqgyUadtmj
MjgR1JRnZg0aZVhkFldjAl01B5kp03sxVux18iM9gep8hirG/96q671IHErFz1yb
6LVUu1nCzD+tn7BW2pKf9ixHm1IEFXj8F2NmJPv1HhHfrJD/Jr09Jsrl0ETB3cDt
6LlWT1BCgJrPablZe/7C1KDQZHzcScdTcP2VQGhXiZGAK5AWPgDa97QltP9mCvSj
7oH20GycHQap+pW0pvz/MuXctOsofZgOEeUMDf1KgGsC3wzztkexwsWIFRhzl6jF
YqUzd8QSbw238Qa/hYllfSlhoBe6olLxAPtpP8XVK2VC+zWfm3D38lMNPdb4B9wc
1bdIQvEfhtlqvP2Bbx2cNRmznDuaCHGXvA9Lky3LA+t4q7TnJI9t3X5CGiHaod9H
urMIYWH8v6WrceJiXuD0/J2Y/1tbqTE3Q2dSpLbDYtU6mqPI0Ds1sqvYZ3X5SK5Y
y4ghQolOgiLusmtIwlGU+pnz+mf4G6axwYQJB5FvtVtFC3ef59sPlsCt70FuGj/V
1KRKAsnbMO3TqI8Cb53ybbPadyQRrwgrRGPHiT+4OZrOipGNEJx10XLggpM1J/Xk
KyLUddxfuuqAulrrr/yLF9JVg9xmLbinNqYL7Z5UKY21yURAHlBC7hjOFLk9jPy3
0n9MeQysAy+Lalljcz1U58U5HD12W86IEYOyusl8hnQpJoMiivVpqc9MxwQQOrN7
Vv5tFJD6te8x7dPqLobGJ3efeHgDebvcsUskemQUOv95qY890BpW66TwjcNkPpMU
dtj0V9XVy9Lchi8/HWWsWR0Kf8UcBHFI62vIaDzqchs4zbP1hbQJY1IoGW5CS7om
iR0KZF5ZazE5qfBD3XrU8cpMYv3asbpZC3gS1KWaa+2m8TbSroaVSjInvPEWFMAM
1Gm86lw09o4QGdtrUVcxgPfVBjYEYMaO8kJNYVNjhyfhIElkZOLVxoph+IlGg+Ng
4H0GBYnnt99zQcrO8ltWCTZyu+kUVAtzA2JNlYVCFwPVzqoZoBHdr03r0DEettn1
A3cieaAe9aNmeIz8lwp0VIL6IISKzphjhPEotALXswLmN4rPQ2mAnohHqxVTKLEK
HHti0XTXaEhJhIdrkBAkEMp0602MbCAzrwniv0gOX9j+awU11z3sV3qFuc8ndHja
ge4H5yx2ptelZJYtW5xRzIqsVXbaeriP7J7fd0fXx8amBUz08ij7vRXuxvyKlm5a
qCNFxTUl4JnqtFF9g2ByuH7Vmvjw5VqNJqdG1EN/faGkK5opwlTlfVEu8hXvY2nt
9AQT3quHCj3dOZwRqE5JNNqD2u0w7kBIbPqLetxrIellt1ik6d97NzR53AQ6wmoL
5RzfkpfuFqgsapRlgdyjr9NQazytU0gUV+moln9kQQ5c2Ssf6usHZfg6JDzk5DDf
FcZP78KUYPOSslhO7cCsKOC8hlcAQK8as3MnH46qrlqem0H58sf16bATVq2QJm71
wVAdkPy1Ad+wD/za6RSwK0NuslpUmvWuxcAsF6WMTrfyhU3HzgqdqY5AmVl+m/9x
Cdvncw/RCPpNswWGPEcRBlQ4Cf2EkNeAsL1Zw4eVUjlZNP1kIlCeqTOxlfCmMsGk
0+2HliCZUMG2YJReS6t3OBaBIp41glg51GtcuBNC8HI4Ba6REDfGO9/8ajmqMwj5
CFOi+9zavtStR0qt76USH5YbduVFuZIxvuS7eWzgoZahsA8/MTeWL3IlYdR68vin
d0G0MZw2yT61AWp/B971uNvb2i7tkwQJr9vdUaAvUtGZg40j/S6PjFQ7PAmgyoqD
yO98mEpnzFUeZf1eyvJ5aGLBfaocChVrHZnLZZvxcfoQwlBWUzvF/DJFIxmO5Vj/
wGHeK9egIVsRO4RICpWLJ0i8Xn/Rxs/QODfwHGfGWVd19TZs/s+HwpDegvncRhnw
ChAz42z5Vc4HADiP+ruZizI1ekQ/RSO0hZeRRwpa50CipdJwtLfa6tpQN3Z76Zte
b0WcVzJ8aW2WBdcda3+0A4artlQDdEiM+nrdOC0rImT1W+zHyhYuMN/ooUwyPtup
6mGBJLeWz+7YtYnG5oRQNsWsZTvHooeQEB+N8EiC82FUqyqSaXJhiEorLoLQiHLR
aFjSvJtPt5dm18oZHtbLJ3/jDp9PT4kiF7BGdK0bpm4=
`protect END_PROTECTED
