`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SeYYVRu1407JIvzmcoi2FCNnllpH++kLbb62MNehagyI
3YCrQZ0Sgk61y32VwFQIattLpw84XnRTwc1f+e4qv4zlxT99mN9IC1lt2tIZ+RDu
jj9UwiwiskP2PROLkNOOCFjZ/U7wfCdzHQMpTiTqEqonU3uXCeI0HLcaHukkPuX2
31Sv7p3BFzGyDHb/D+vhkR1EJKnCot9UnpvRz18mb1KBuY80UNtvaRcm0kwX+4ws
7ROeZbZdjlvr3ImVwMX19sAqYMgTklnb2lgNausabpGX1zO4iS0XgpF6pe2sveVc
L1ivHFeL4a/nF0r4UT2KxMf3NkVRfkYKmhvA4vp6JgT2dGlMMxFISDFrNZiC/9vH
Ukb8bHm2z+5eRo4Qh021HqGAJUyIJxRIMZsQ/RxCSkDoAfaaaHuQUOZQhJHKivB+
HwAFfLXS9skfWK+UMWBnMdG6DgN/2A4+/uFMvvOxXIiIozO7lSbZ/huJ3VF2D2ka
OhOEax3eE5WFdvFvGTmKoROMImqu8xhosEkZuLPqUmdSEBmFInsfSrzAnc4vur0p
lqVmui2TB9ZbicHK29XCn52FrX0Xbd/mep5P9HHZrsbUVFV3DAv1+Hk0LQZaD1yW
8RCbt5GaZk5ZltBB9262w7hooNU+h9ZmCbEStoXvS4UACSleiDdc4jv0VlJA6Vmc
`protect END_PROTECTED
