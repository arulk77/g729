`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAghKy/5kCAnW6lzk6npZFZ+IcZ7Aw+1uo2bAu1x8mxL
H3kPoUdX6xUXVKifaKbttz7uFq5fzd0WQzvyQNRbNxx+30PAzfVpvbRgsVeQHyIF
DeU/qvJMahh3p1aGL+WLxA+csvDWxojBtfczLrx6BOTEEOO0xU+8QGIZyt2mTS9H
3qzbLoS8TgZePUk0B7P/M6FtyWIw30wKeXLiPFtS6h0V+54gRKbeYszqx3i0y7Kl
PVf5zsH3BQsHMB33R3AjRQNTPMC4n/7KpRE9lM25zR16H8Wabny7ZalzLwQEbX9h
egcgb9lbEHWMqgy5QcIOuY34NRCxEg+icWroBSG4dxZbCpgZtqCoMI6LaEtWXXaH
a1jxgp/11wLH/uFznV/Utc5gVdDL354NgVxpYOozZjD5UVZ8uhRxQqSfHI9+XReQ
v9RU1GmXUFqG9WT1I2b2dpU1yxBkCJi/SEa7La5ilkA6m4hsy5Px4joxICFwSV1E
1dlOAamrMxn7xpriiRUyui+Kxfda7ouvPeEXkZCySoxey+iMccQnI/KP+Tdn22+H
FepjJpStCU3VUb5wCvUoVlia8nm0Xqtgsn05d8/mnA2GNYdK7TZuZ1ik616RZHYP
l/k4l5RzY7yRpsY2lnpWHLqAcePbt3JcGPztEX+8Q0Z4fzh0ZllQLVhA7GWoUY7B
/HUefnALxVbD2YZJuAZwXiZmzoa2kDMPWcDdvz/6onIUVhD3zBLOJMALrG24bZsU
6WVHtGGW1I1uE0MClHS3wCIcwPIavZPEmrjIzugOZRcenhCw1gbGaCt6OSI9roXq
jf/RnO58zcUKreQl/BKU+mrFYmXrm7MZ23xE+/YA4Simoc8lJK6fQneg5C2ZgI5P
GnfZ4XrAUlIihrZgqbbhqlrmoXfYzLVyvER0d+aBm++U3ymwOpBkqwLWWlrc20S1
qaAFH6yuZIS4QXUL2O36aPXrznLDKQNVtFZp8xSx2f270Jk5ZLAIoznOQaJFy5LE
Wja7YsTiB1gxcBtiEK/+QrxGn2kA1vdIp8VC6nJ0JSgvNKb0FKJh3OEyC9Iq0s0C
RswIVLzCT8IhPizGmFYnH8L3v8OxgdDSoxm+2A1gf5XZJqbX5pkRzwQiqOLKZnBB
c+OfBYBMyXdWD6SL5NhCpARQgKJ4tMj/fdHQ02RfcOgzK7vhNO2UWpOTsLTpo//1
DqfYZD9UjJ8UU0qLT1LQMvyNOjm8eoPs2uGQIadDPWF5KPOfZNB+X5JPXRXpExqA
cgySld1ghL475XXNNq8vuHwIz4nY4D2dFPH7Ol4tgLdiU1qLIY3wareobywzUknP
yldA9UnsYbcFV7hc16EjBXnPBOjHatwyXoxq7zdeNKVVo0YT9S9kJNAETD7QnVBC
dXF2+cyTnog9QM0zSGhbYP+bVSgAl4AIwPQGhrKoiQWUH41Z86ak4v7hlHWbmqfb
PKRkdRwFsZn20ftO/f/cMifQWNfrFdR62HJbvj+pYuQN9DpJAliJAs++s76IWQzG
HYGxnfiJkhknS+/DN1C3QT+mKf8cBGQY8sBhhi7wJKrkcjMAVG+Ljxng+8VEi44v
5wjffdTD5PRstNC6Cj/J9xzYMV9C3/nbi4iMNRSGJoH5ZWGfGE0qVvQSNNKEjpEk
B6s2PvxpXCrFsuLooM+iL3yWwX/ArawYMzRhU8bszjpKD+f2Tc4SRq52rNnhRGS7
xjcat9rwDTxTmZlt9AeYZg==
`protect END_PROTECTED
