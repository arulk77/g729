`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+BfAI6Ip5R99J9+tDLFfRIGCv2JBKQPzTfgc5AVejmb
3x1aarZJzQhIu1O2I26EofZhD0g9DZvmkLJ8mkL1ZNob5gL4fdBnrGAXG9A6FAAd
wGyRH5JXUraajX/mBST4JJObffPRiKXQR1C9R2pispU=
`protect END_PROTECTED
