`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCAFFEzHpLfW1kNvN51BBbW/UP80lG9T4DlurUAlJRzo
8WPcJ4qtyfL6cq9NsSpqAezgO+s9mUvhsV/P1h8DTGzpVT9EjjTc0IxQw4SFYOlm
kcKIbv7KDPlJ3CimsctZibOwXOPQNzNfF+/6cNlGoAjBAotia164NuXVMIqFlJDp
JfIbt8d4abk5ZihExBKWyjFWL+z6d38O3ydf6/D+jjFmgqWs0hKZ2URkYVLWrCq5
zM56VULcjsUO5IBwFVvIdUZrDeGLKk5zuI5PzaQcryBGkb/lmDubPQikxA+PO5Yn
pBAzgWMCTidVBHydY0ecgcW6Wk/iuIVg2jQT+sSbQRIb+OTAAFzcgF/v28KMAncP
6Sjf0DFhpKSodh17PxZxOyOO7r0Ly60a3KXUmuv9FBI85S3DEIXcZOtSdt8p44ix
VTdZpZgh4TONb4vpG0b70r/vNxTfcVvo5iYjlAWNZaCppN8r00XEJdMJKyqnN1qy
8CDqVdK1j6Hu8IsCDKAT8JlW4uNsq5EOsaDsCOz6lJJQSFJe4lyKojzExNElB/PB
`protect END_PROTECTED
