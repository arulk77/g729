`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44HCKhchrzsABsUw1MdQIBWxOKZqMkF/kk6sbLxvAE9I
8850IhON3CFNpyxGN3KE0hnXyS/ZcGd8/IDFmr9DyNxVuIduPWWVBAn6Eo+amTRs
HZsG814KJZYZmzOlmARNOF6E7fUKjBucnYvvRGw0bBaUmQgBKXEWhi69qZNaXd//
3KRCU9nBmR0FjlKY7DSKBhopKZ8TzuXIgf5bojdesJ2cz+saU39jEbzABrYvPWyq
or1k58QmG9LzZUvwBmigrGZvaEGmQbb+VzQxzX1JySWe5N7TctP+539UGUHvjMle
+4z8nWoU6QIVRkuds4bMOQ==
`protect END_PROTECTED
