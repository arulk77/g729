`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLT2YegYxGSryfLTGmGkMbq3dTiX/ZlpwqAvHx0fkkwQ
o0feE4N+fpG23mTHlk7Z3hVJsWoV8xrbnKN1cZ0Hj/xnOAgxkB1u12aVNTYQYPN1
C8vdN4xGNjKRZZQ9KjRhHJ6lE/hkjuq6tz6d9rk5A356a9szvLJCx9BQOBApqwEv
1C+RKbN8UbuTEhINQeXWMDb+Z2uGA7lXdB1ZcKtKXGRZjfGYCM48ij49xeDr8lCZ
EyKmilf1b+XxUXVm6VTihBaOUh3WBh6cUTui2bptOTvnTn1RytqxmPNOoXTmFNjr
/HkdGzhoVWgCuCkdgTGdxK+5GD6iZ9xmCCZl/KxoydSN+lbx4KcSsU23OpqCO7X+
A4WBMsDAN9EhbkV4aWj6n8QBowcKjh/v6P+0C5N64HWqZ+vUGRIPyYVDGhknS8Kf
7UstMW3VfVXT5yV07EKxDDqMs6Q+zvPXvrEe9zNG9DCSc8Tgf4iuP5UQng3iFp5u
xzbWNJSw+I6pJu0bMwBKGwZtYATDUqwmAfQeV61HQM9dRDUL8G+HGFkXfjM5D0Ro
93whmSqtZ7C6c/f4UCXFITGSskZSzAPx+ZXf6IvHsfv69d4nqFkInfohJxrz6uiV
sNBw6RBcwnw8ZwmZWn08rQpjV4hOJLbhBjKJvTkTJkvK8JC23Iwndu9UcID3Qh+G
VFFqkYKTCqQueOAG4vucZ1JVTZR9qmOo8YxA2d7UMTCue4IkaU5+rfJ8t1ShH7s3
0WRrDaIvKCydCLOHo9N1GBSgKKRepwnb8c8NVHxxKsrNCta1MZBLROD6cX+elw9U
+O4t8mXdXuNDtUorty6BofvG8rmdHDhXgTv/RdczTis=
`protect END_PROTECTED
