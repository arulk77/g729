`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
TtzqOnb2bi773XQMOlzcferjlscjh6Mwm1t7A8r0JfMlF/ETIKrdwmS8tg71gel9
HLXG2cjZ7ebCX5p8aMRD498gPgirRg3O/8LChFgtuafzyuw1Ic62F211utqq/+Xs
p8Z91OjIb45GUHWVwUpTwjTG5e4BVXFCXdKal7+PhDaiQCNlATQawVvrfrDdX7Ab
JGcvuffsO8V5XKVLUi4mLra5QaaU7iBfWErD1dL/iX5u/KtflKk2kf0KqO8tmNXP
eEcWTm5E6HElODRRZF4GmWtcx+aDSxlEYA5XoCJeg068YYTrNb9JJd8QTYVJ4y+T
FWfgw757U3Yid8g6u8r4PFhcrlJ5ZRa9bLueDlW4Ee8byd73RTKxTl5CiNDEQ6R7
FOjvr/izpVkLwjcwCuQqrflPGOgJOqIakLq8i4DotFZHeKJ9n4yPW4Zy4Vy8gart
tGQo7Q+uYvcf5ZAYLR0Y2yPYNEAvrPt50T18aUw5v2X0OKJdqsIddISLaoUuvWdy
iw0UC9qovSMhH7RA3AdxbybbIwtR4SVlKFkbRYt2cULfgO5ql58cvDZE2zSivn8p
BHY8BpVRfjW8PCatsx6f+EfCj/zxFQIFeUzqahHBsKDt1kMDDxssfbaRWhv7BKkD
r1EhrMPDtv72FPXMEXTJVxcYnm0oykLb9lSep47wg9CBZOwNni5QOevSGeZBsbxK
T+bFdqI1ZHcBp8sTV6X114aiesWlMegqd8j/jpBbS4J0RwRWrRrk7rcPk0FCe6Yz
QxAQsB/Zu/PJ80cJw15jh3cou8ligB8/t0TVadKz5+MzCYDx/tbNQYGUWGWtuueZ
zz1Jdd1dUxlDAfzAkQPx+fUxkoCHk1HR5SzV72FMPAY6MMQs04dDMtLzDQtGgJaQ
jE9MFKcv8HETEhjNPW/sJtrsniz05DUbeROP7NFmC2GYXSpPLSweAR+bBo2/FTf6
Cgp74bUlOINlpL4GAm5isjpzdnsLVx8WVy3bBrTftpR+MTBg8nv8wZsE4+vIPold
sn8AqlzT3GyQnFevE97N8X8Bxq0c49faiRfYVHaCzX0A8cYRKphMhPg80+sIftyv
tNnR+/Fs1QqLRIJK9hPLmQJMRXayGRxjW7NrdLPGebR8aJh4rwFp4if5CnCAoMtC
wl4Y/vhKNVxE144gUKz1W6227YHwIasMlJnthpZcUDyMU/XNtYOgh1QKBEOj5qvT
ei6tpwIgzUkmVmQudFlt1rxl5fnQMEiQwfVbloNTW6BoYe77fQ3G1S5nQPNZbIXg
JeUhpOzU4nolW3PcMPY+2yBJ3QA4lQWyZPXORBQbXvNZjg8+Q3B19PWpKa8RgMFs
Qbz+O/UjUBWEfselMXYGHLc1scUJQchT2XTuaXqUG0GIFQecykvejzWQWdwA138Q
snl+erlkSDr4xy6/HRdpuqpfWSIjkTmlbNOMA6sEtzLRCpbmRbyBteMZyLkTlPrw
wwmrB9tBfHiEXbyIlxeDi0Jszb6kOM5GtMHrGWS+CC3Yjg9kO0H5v0H7z5ggcBGt
NZYZ1gjl/MjmWB/q9Brz/FduPW1NuvEOjW2+NeBSUAHAUpoExaeybme314/f6Ycd
A7N+GZBISp4HNk9gjG9urQ7L4/RpSL6Leionj9/9bbhXHlKOXGoonCBR5Fs9BRka
/nUTcfsTmdUX9MISQWjp8S/3Cc7jCIlxcnxp71oxP3Qsn7kzj+RAfOF8LyrdvP2p
24M7Ocnz0ZUHKE0WMM5FHMWfFFVjxYa48bCUGtFk/gDx1Y9gSVFVQTtWGqO0/yYn
SuXP7CdsOGIbtp9n+lhvwkjMwXX1/QUmn8GaMARDKRDsizIxbiOgogI7F77JKPTX
I3mp/toWlKsPHXNRqD9aohf62lJzLUTpZEieRI/UUNMuuxuPjO/6UGunT+as7iy+
UOvtx5KsE9Qj2b1w0Z0PuXZGRwRmrJ+V4wIHsm2X2JRN8mEJIeTsuMA380CV9V23
Q6JDzOJuwLdzMhs1kV/wakWRTA6/OSIml7ndNzzU0twMq0HDLnQL6rGFESfIV4NX
47CWge5NcWc5un6m3zQMLGWXOCJlRU9qCVNT2WGwi2nQ31cSYXH03BWgpaWvr9kS
IImK1qKnACjSUSe+nwA15MuSBV5+mYHWn4PbQS9ERHFdKXWC34Zm+ziH4kv7PyM9
pCTviZm+a0+CE1Jpu8aka4sfIye4qNsV58Tqi/dZta1IYcgw+OwQisZi8nAbKrCp
aWltvdO48YlSFHs9e/aLa/XD4CtMw/cP1qZMhyoSmhvvt4lmb30do4snX1gegkpI
inArA/5ng6R/jIM82N2yWR6HYBez3m2JI+L3sQEZmoWHUys5SoRtza//xuUy1MzL
wk+BgWho6m6h78S0KjbyOtQoDu8zvL/9sjPzN6fExZxSbi9YYkBDRfGCKqE+d075
v76D1XFzfHPPtIdpXYI8XPI1k3e4BZt37vx6NjxzXesJnqxtrW+/t2OWZPt4w0qL
GYAapQminhrNa9O7P9HGcA/MjLyU6rE/XFd2tgIxSy/R+ji7fng3tjB8ZtyjI13b
oe8BxCc2XVdeukdUTW1BJcLOkj5+j2dF5d54CPpLgVm/5ytD6+oO7vWh5wqH6gO1
3v8rwyQc0kcYcqZU90R/AnK4Y/Yf1KJgfCTRoWNqsjF/chxvLGnHUrP3RJ0t8bDw
5YZk8kapN73cizxLQU0R0A0cLRiKzZME0EyQz3uMyNMlScvswKivJ85/R3e2J5gZ
/fA2O87Ksw3z1jDtheYBTUqvL8lWOXyUfLmmMyg8maBfCFbsekHXYjKlvFXEGEXp
yQNgYRMqxHgAG+WKh8uVtr5cVSsOJs90seMaXWDG1/5nNREXNsRrhB0zwdt/R072
OHRgq33F+y5cu/PqlK9YxeD7PBUaxayxKmlJSC9TR2TAL8M6JsQ9g75LTeVi15Cz
tFKY97pnudisj6ovQT7kS3wo9DtlSveDKQCZU+pRTfpk6fkoDE1GtG52p9Celrij
YODDZTqZbcQkHeBQgylFsfsSATgOtAb2HmaxFU0Hrl3//rbUFAE7XuH4ekuEDokL
VMgUZQ9ykMpe2Ol5lslGgTS7LvzFJ087/Y1NCr0Npw0omz7TysJgP3Rk7LGs1jf5
g3udnRwjS7BpS4jI6LVCWVYaYLqKvw7Ovz+4tS7/loYaj4yBJEA+gCoXODWysvE1
CgQPBk81GAm+HuAtbP+pKFxe535/JRSIDSoPGO9yVHB1zbkRRWnx8eZpmIm+/tP2
uL8Dod0scu9k/lN3XAtg5ocLsov7GeGstNwqxkOkCzlgemEXzGQqlQKjqiA058Jt
o1L01l+qLJ3mKOcAY9hkev76xSzyrLPt/kJjAkZ6aqJX/Glh9aZALbBQ9GHBQB9u
a+49KxhvObcmyJUJcNVMYSHHa1aRGNl2A2bO8uEGlfXdU8JYfEA4u3UMFWw/CAfv
P08J2Q2ZR92eT5cRBC9W++DEaD0W+1HxalbYkcAbPmMXlNcXKDmDFbCVa5xTtBKa
GjwMpJ2oX4KAumyfoGuiLro5LBchiePMAZ0PGOTCcQO1qZfUFGRNO9pJZZmYuLZi
wMyeBM3zlNpewPzgp5ttPyNOVp+TnIuLA+4r3qBP+fOCpzgBc2MGDVbm92oJ07S5
CrLfkJEZN/4itO1F5NN12m36pbk9fJrLHkEqsCJf+5pt9bCDTx53F3UDqSwDYuxU
UPXXvHpUdXJ9A2FppkRRDAwHoQQ80KC3Q6ZaG2ZRSVwc8Up6Lgr14wmW82RN6rLu
W4HpXV2eSD9zwIC2kyde1MCudNl6qcb4VyvvfQbUufxdl1NNw/TimGSPweyBitnZ
nwbXEmygR/TQvX+iP3tBT8KsHgZYc06CfD/2vDDtVgHy19L8K0p3buVS7Am7DgoH
j6FJ9yBB/7+lxNi5I5/7GPeVTE6N1jLzPuG2Gj+lnNaLIXJh1tL3pex4yxHR+FZS
1I1yHBISrj2TnLJxROR1I8AT6iM3xnBjHvyXmvF9T7pZ34ueqJhM16PTPga1j8Rh
B1mKSW9wYKkOnmpkK1qMimco33fPjW9lZeJcUiQ47Ng1qDiXb1HDxNYLpDgZ8+7/
Jh+PG9u4C0vL576Cv4xSIZUjgG+aWwrYHfXdF+DAdIJ3MV8H4oaBz//wVDkSUUqX
GdSJU0JdGvnu8rbsY0t164ZF5zTVrLYtFJMfaRvWwx5q3cgphswKHw0yFb/sHQhq
Skuzs+u7uRKK3gLEYTWtnKb7aFeXtdL38za7YnxQIpo47Yfjpv3OEhCJaeQ6FRhp
rPmhiywaAPYEsfl38Ne4/XQl2cGDxBuZmNOPN74WRNev2Zska6SVityfqm6BI78g
/4+0YebVJs8xqPM4nr+PjCDtgR6AbIR4GBRnhp4Hgp3jqM6+kATdpggCg8zklj7B
+wdWYLar2kY3Xt3YkZi3huccdafFv6jyWhEUrUVOKu7bCnIEG9T6b4juARYIVqC8
acaRHirL01+mk3CjBLdGAOQwIgQIXIdifqkaHelLtJOlrvXshRnqPYC9zyvGySRP
aD2kpsAX/To6XQlNWLy6XS1FHQCLkH4pGfbkTsfKlirfe5TnE1j/Jiz9ugHFnp/S
dcbGb0138Z/1KTIK5Vsb+sgGLYygRdC+ZWNv/yvNOwYJZIutxGXzgBTnxwN0W171
EObgtw99FR1nV7izFpkuXRmbM0xwADAMXx5AvP0e4JhG5vks8K+wkUsDR0PBuv7E
H5iVvjrmo/Aro02UXp8qIsLuzcYWJbNZ0so7XyAZhZc2wDE5Zsn81ubkKr3KSbvn
R0qrx1pH1F6I1S2B9iZkAKQeFwvVtUKi6YAS2JQA1TtxGbktfVHySBdJKKpGILUr
KveXgPBe/G0RLFsiBrF+DP3a4sw9IxooGxSF+2VnpWb52ZE4uaGlG81nEz1M59xo
R+dSyBuVNUOwEARIbMz36sOKArlQqrn2M8cxMsuEg/r+fN/f/WwiPIVcZuLDhDod
gGez9qzYO6nkm+X5YyB76gw84UCS+XRZSZpz4DEdSxME3Nw559lhNQ7JSCqg/maK
Oi7XZjSbfhnPMaGnLogHcr1S3WBSrcqyfEPRoM3hnRK6RS6iPuqViIx1LdHVCwEC
wCQL/A9W8dMtqE6/RMqlpKYEz31E15gyKGT7q/GzxJ28bBP66Fqqof2OVtJ1ncxC
cH36Bn/PedkiDNfwvG2HBWfq/OT8D4qyZu5CaG81T4CbPA2RTSKgfNV6v8ieZMrj
f/cSkjKvIHUYVPGkcaCdF3niRljqwd0dJ21DBLWPRVqOrJzxdeMjf1fQCk6WI7c2
JOyGppDBwFWPrXv0MQzyxxr2gzl9t/104aUE1tSKvrk8WBH7bQf88zdEDHRYhggj
Ra8D/GAjVXTR9fzD42TPUpttUc2DNC6vNAmgmz3ioc1oym0/aquDMxbW5sTmJyFF
UGUd9wI7lJrDV6+XjNQNUUdx1Pxqd40dx3ZnQ/uomRjfGNtUe7MkqV7sdMX/EJrl
/cJ4vfIPNxNAyivvV/i7iA28gndQsFTPZpohXG0ecrnC0o3rtRiFPeAfHQRQD5Qa
FRC4Wt6KH5FO/za4FKuvcc91raaeg42c8FVOh8UvfYyr0kvH53I9MUohO3PNbkyx
0FFUoAHDpynDtacHty/H5B95RhVs1yauHUcQD6dorxKg9p4QC3cLdkUQBWtnacsw
FtFH08gUIAe+Riwg4NTtMG6n5YLQeLCdm0aqEZH8ONMRuH+QA9X/HGahqloqYcp3
BnFXUZmdr+m6fYPCLzh8yyGrohvZh/fHVJ+d66YOyevWpG46dOKyCvqE7oHjtUNJ
7fJtZACt4cx5CaP2mLEDBh7hnFDjW9PHAQ9vqxD4uRnavfzXaiVlNO3hl+h4azoH
DPfrop9k5m6gDid1Zj3XImHYx26UA82/RVyiMLbkLgzjCNArjVOwFtKGY320HJdD
sVq8MkIPTYq4HMobcECG0VwggyUk1b45uPx6a0F3+qhIgzk8Hy0lWjJFXaQW0um2
1cN/Kt5kICSdtDICFKRvuYI7593XopVmQe8Oq8z7yqhLJTCmVdAsw0u6OK8Cga8X
aQmpK5DD0Mb68n1rAq/7UkxQaKOaANhOES/ZMMIwSBbtKuq4bTe/j03l/6rXn2+o
O3M6aWNp0NZDxurOAxsdI5RXn3Ab2y8PVOdUA2zgWIXicUN9XpM3qcmxAnJEdjYP
qahqjCbbhmwn070/prpUqAuxYsypOneMW8PbUWDShYDYkOp9QkmPu8Oyuth9ia/V
yncW7wGrfPWeepduCYOrmQzTZu7xT6BUI9B7SWKoOjPw/emouJQCkk1FwXyBQZwV
/xZJsAHJm4M736YjQSp4Kr+9wgK4nf1P2PSuhx94tuuxr+FrvvZ5zauuZ7solCLY
JkhKtfN8RO1AeITLjhhiptZqAZf7XkuhXSvtGefhPPfHOQRVgmUe+ekF+fFlgtsd
F9aHblrtWATltTnT8GsTKmEIHgQ8dpIZcCz+KHXR/k9ebb5ZxH5UBCLBOYYk0yA9
DLYaM8UvJdZHjICHkn/T0SWApAm8jWFrElLTJpo/KQqN/L9pjvg///IgL7BiZ58t
5sDxthobVMpRp/HLWBJfo8NGVVBBBDkbpxQELur5JM6/GrtSCj44W48qDCeY5iwd
fbeuC8FXfAU6jFUY2Q7dpNVxSJqUvJkjRrH/5Yo+AzUOEilNeGjgpd4f5oaMj+FX
XtgL1qlaUcUaLmy64xiamzY9+6FXzjz4LwJH65rw+M1mrJIb+wm+GdIJGERIhDBi
uuXMf0UudKATfoS/eGbCrO9rufoulLK4zYFRE/0/k47V3EQsWEWlrjKa+UK70RQA
3RQEK7Zioyx1lN5MsafBhjHOfliHKn62ap78qU27cNoRf9+qynTtxX8tFkT98fKZ
iHeBAu8E4wqyNAKNkYMxdevvifvruLghtQHCd1xk6K4wYBpQglsuVRMOiAkVD2II
LsHTdYc4K7lC/EUSq5lp+zfgv0CVtPIBvnf1ZUcduW2FaEJYOi/T85ZKUrNmO1xe
f7nsWrq4/8rOpRDBcjln8bv9TmKD/x2VtSCHCCpIAvDc6PdQowKetNIzGTUoTjjF
ivNTRmaCxieZarP3HKETrcZkeCBbuGsYXqSuLf6t2NcxKVrvpBZXPcEmk0SGWSnU
yHQ21g+Mzk8Melm6jkyNR685yZoCkKObtAkL2X05YNt/q789nWPvoDyRKfhu3vL0
4u5R1UboUPTaM/HiuLakdcMqiOkAaKEZFbGmDFf6ojdtStC/ozoosuG/jLierz3i
sXQp7QZrxgX8CkQBGbjvcTQxPNnlpO6yHreWz+cq93Uxxx5+9yD8pRA8POP9cda1
CgRbsl22v/2wlgz2kr6+h+BlYduUvSCfKyjeYr0LHYptYoms52l4EYelf5MxNisn
uUVZyf00jsgNek75x10RX0L47HsGobZvU3UMSHrbA2DftlDa7ti4aVf9GFaIr6CY
cPQaEh/HY3vkVISfXNtg/xo8XjMLco/uV9CfRxPGtNfmT7ftiyPXhAB00Cl/fhpe
A/qkiFpdCsREqk7xKLCVpFibjntsWTXg6otlM2b9qzU2jzm0ldVmYqzGlIaYWcLh
zhh7TyyJUvkjKrx0Lsq+6vsTnuF27WxhE2F2Pj2rLj5y0piDjSoUQ82flKyRoF27
rWyzFOR2Py1zEiA9gP2de0PhkG2TWdEJ9Jz99W9+Q0+pztcb5jYPuxWiZz87Ut0P
WUlUjxh6hpafeMEpfGFNtVwHQWnzhmcLxZ33VgaxwDJq1I5fjafvQbWNGnysF+Ks
YZ3XQdxBThamLygV5DEXyvHKbxVmgumzdO/zhB2nbbdvJ9FhXReII4lUPxwftvLM
nB133rB0pybJtt3QZeSV+nSiM/87Pdtf8cdxttugLt8X1vf+Z6UlZ35VDWmfs/b2
mTJ8ueDoy7HDnUpdrN/UhaBJwo4GgP+xOJvehYuB40SLtwtlwPMmbCcPVApkF4Jo
rryOjaAqiWOfL/cLVWJpd4mk8FjEEKyEjFS5H4go3caoWtxrCLUindPyxogittCE
nJHwFY+ThKo4ph03AgIRRWTkuXU9pgbzpNyn1mijEiO7ob3skGcLIf+S1ul+QxlY
Ifz60+aSWOKAcUQd7Qw9cE95xKe8pLbSQ6XqLVUHaWyBoJYGxM0pCFDsyi3aVrTE
x2rMMGrfKQiGnY9vimtCqUtvjnau8gxfYSVs7kOWwPt8l2lFq94G7iq92EAMg4EJ
UDIFlCluWMFVG5GNzZG9U2oThFaWDVM4SdNzragBddRDSbrXbIpIDpx8NQlsLcRQ
1ZfXEcOe0p74cHlX3jd0WhcXxWSw6jfBJp40XCCsmyJrbLBOak/0jWkuN9YTOybx
hK02mdDudBi6nmxcaPmu/0bydvEdycUefkCMMX8OLmBvvjac7diaAyKpVnN/3EL3
D4JAdEa9KTPPn3V6/55PAcy+1h6W0RyjkmqhweaEd6fP3Jb9rPw+hHalnvxSVlR8
HBhqQL9i3TSDlS6a96p96HsiJc8382+hwJ8d0syMJOOi50L62P7x+isRM3WfpKWJ
aLMlXOt2aB0Ifkp5/c6O0+nWPGdJM2kLoUfbhLLyqdJSJiDIHgQtihtH1qWZWZgp
cM1Udnz+Jaf3cgDKCCwp0Gp9EeSJZC6xtHM8xsXv2UeQmygSwuYg7ywbK6PlMVaf
L9HvmhKbUWKfG+8r1FMXUA0sNxHxCNEm14v8lwCRMlxF6xI1ak+XaVMuLmRSjCKs
KdkoGui3vV8ED3lXvnT4JsTbSBMLp0sygTmzP4Byz2HbrM6zvI+4jYtGrgyxA+Mi
/T0jAp9gKpNLhYvM58XW6uJHTlpPNkd/19bxU4RP+X3mZxiX7DWjJYk+adUwzCKK
XnZnKVCzfr/IxxBqQEL5epOCalOsYd7MN5Wc3jVYJgz3sXBvcjHWBsvzswo9HqEt
bEfXJy9++5zY/Nn06IDdKc3PSEuUtmwslA9M2+wg0eLSoHQQ7eV3J6qVjTZAmXSv
p4yW6fmq6wMU/j2Hq0amG0HDFC9cn6TUgGp/CF6o2NK0xQcJiATqAbtCyjjz4lRU
SbzoSXYL5dDyuFrCyhcJ45OLm1/D4vG4DdrUEnKr5l2lDG6YGt2mby5KLJrr5jDm
/YFM58xiAeJ9gatm8KLLFrENXbfXZAQYPwokrIbX+odQd+KkHsTptgEUkVCq741i
rnGE32icLiZQH7bJRTk9cwNMieWQgYOBZ1uJbqTug/ORfdEbvtwHgxbM6cIst9I3
00GSPoCWKOzKY9WRoQ6l11es0zGxTquse1eCwY4mTD+26sz1zVGsqUL/1MDBOlzj
Heo13s++vRsmHjz+y5ES2bjyQM3zNVevNKT7I8uWO4idJh8eu27kiR7KT1Kszxn2
lpLpHvv55EDo0ACS0zsZIWYYqjpJkwM9GzXymxOd/vIFXsUqZCCaV807+v95MFWe
CeRokoyNoZLdTNmnAE8xToCe+gJMxjjiCBSDi1wAdU+tmYX45IY3oBuMT3cCitFO
z8YdWb+l0HQd+4kbgk/pCAVFUTAEaoI+cBho0Ykvgb6PqZCbIWRPTwLWqp9ty3jj
Xc9WXwpzWaGNUFcS0zZWFhwgqnjo01trBeuEQiy+UjkdOBRXQ/DvrnWsT+95G4E/
Kq3OfFxd84kosuHCcQ6tY0sfKjmU1+gFn/KJO/6XtGK8KsGZKsbuVYwbnbwnB28o
ISzSS5DWnikyTeHOJsQ0xjoSSnsymp0f0teDzgmRjxs4pkoW1rcBlFgbd86YeNyf
k3aU1AUTell2ZSFKbF1egOjzUenOmfsgkeFNe0+qYjtGWwZuD5g5xAMBBrKzWj6x
YQc89tOFZi7KSS1bvqb5+NnnXxM2bLr2xXjp9a2w8abwfSDubtj5zhc4YSiYJCnL
FocjmvTHoLep0bogblU8HhnSNGNhI6Af021pc2DAUdlkLm0CfL3g1qBAfnafcQrw
CDt1LyQPnfO3XLFd3caPJQ0LpR6VgbSQAfpD7xN7YunKQy4Uo8Z0bnFmCUpTWRjm
qZnO4m4/9SlJMNI7AdyJ2okIeYdMH4MbVrdLfjperQUy6HhaIHvxoYEeQQBd6a4N
cPUgyzO1K/rfdwQFjtOTdgVe3OgIbEpaESc14izbjWNmRB+uSQqE0bsUSMu2qaEE
/B+Rdq3Mkr2VB4VGZr36kzUEkO3Q34mGOUOtlJ7hO0c=
`protect END_PROTECTED
