`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAMugcxfV6rwEAHRkzt0XFbF8gxiUxxGOXicN2Qgdu4f
iVNLRgaGleNMaRnW73YO6w8biOg2hgyLh9UdcAgROBPXAcDpFReiyaAtp20KvBLX
3Kgxt30jOzbScUvZ4SBOhnVQVAnjdcmi8Buwn+xaVolXlQJJELwXZA2n+pj8QCVY
D9EcNWqE3U+ZKjjl4kJrrxDRx3yWopIf93CCdwqauV6QljWF5CmS7eTfSNVdmFw0
5J4FOb0s7/51/hSh7f9DUjaiYKfkShGTiamTlgpLva9Z5MnDm8VEO58OEZRnjKj2
hQ7V7/yuskds47hGAg7tow==
`protect END_PROTECTED
