`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46H/w+fWGOB7B6BmwuywhB7UXHzoBNeqZL9uc6JxhPwN
94mWEkVGSmw2fyuTC89ugmx3s72RxB3eM8PyUuHQNY8tufQBCxqwQFEONZIaikdP
CWY4qaIVfxqT3L1YsZu39DcLYPzT+4EpEWrv/2pSWCh3FfjgrN24bLMYCR3DvJqF
PXtUtB3JqRHDZjxRaAp9SeTNVHLE6iGONk3bO/JhZ6+B0uFnJ1Isv1FHHcLyxMof
kTfhjMFxuaxPHija5PgscYWE6Siqtkg08aJW0mbs+Z577okPan8adqQpM6guGvCZ
qHE7AccOU74m+HzCLWH6mA==
`protect END_PROTECTED
