`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C67LmM/q1CGNUbXB0qFvYlOt1GeoLK78Aujn8vQlHDEL
7o1FiRjoTqqekNzEjLRMWvIMVGU12eCTp9CpzQy+evdRa7YItHqcR/q2FICCYl7Q
PrI1s13+t1t/RzLEvG5LHaNq0yv5/i2Wm/cJMBcCRZpqUR2Y7olvgKKwXNlmKV6u
tUN2tHFuA7J5cXLBYqDNNfzeSHaMqeRofiMxsX5pqvYRSAoOacaZXofoq6ITJ56w
mKUAZdGbVeKSTIFx66Mo4wGdJEFmyd11CSYIHQwtz61cPq+YQ2RRT/p8z7J+tKBd
sAsa9oEn+voUIiti0ey+dA7W78YhBOMhH2yRT6NZm/8uwJZ7XredQRxc2vRIoMb9
2P6uhL2L0FaOZfypj0Ln68XcKnNegN5apuebplrZgsbhBtsyUi0K4wS4N55rRaE2
QJfmBNLftmmxplMM153rGhO6aLdjCpXQLQAeIHjYXdLGXRwQ+7PN9daz5gt9mCgA
9xSA766DA9cyzmJuostToQAEZVBmWsdKvvr7LI1oK5DoX1WzCUSNh/XOPezF8tfF
fBgWLTs9cd/yP/dmXGo11YUnsHXgGU24G40GRKBF34AIOi/vUAlEXpgYKl38Auqd
QcKvY90Zrc1txpX9dxLI1u87beQXa6gJcP6ajx8CVzQHl51j1NzEwmWCrOHDa7NV
VjAEC3Fd7YexKsKlVONGpWw05Kzox/v1CY4NwZiZ+DPMmr9U9M7eBqi99A+8MPtC
dr5QmSsBYIZ3/qOHSdelpvD7gFifzg+9o24D2Pk6lL3eGwxxhhfkukKlEwULcE4Y
C4R6TFKr45h6KB4c+aLjL+fNPm9rx10vXFEs33utbsePs4aky9VWIFQK10JoJkIC
M2ZQvLjghj1EaqQ1jq8J7q0E9ERgRJixrUENv//wSI7nGnk+GOWnGrZkb7e+GwAK
VtFF/ACD7EC31o6KrybwVloQqDCfx7nq2Y1PBu92zBBNnEEk9IVC+N+2CHe7HUGw
RZz/q1fbZHF+F+D7Lqw21ACEffsgFprrekUzvqvCSR0DStlyj2hyaRHxxREOhZNY
Zb83LeC8Dk9WkIoG5FG+MBdQAad7TnuXncq/vHdPIVVZio8E171bcY1TSKImT+YD
G3cyF/BXPwik/Cm6K0wUQcFuduPwOZWlOdEl9IMxbXDyBp/NPXIC4AK4tSb8uSd6
roaho7vKfOTCmKLWWLGnY5ZwgxrBM3356tRS76D9czCOaVIh/GAMXyxDWhsRC2ct
zR6/4RGIVk39kba/g1qs4JYBNfcVS4jzrfRCwkluw7PUU0BJ5969u+IgRw0e9vA1
r2zmN6Weegct6kPPHvbQBG+T/1xY80nrZt0s9sY5j7vEzvOXYhsivykVnDMWZiOI
+Cuzez/X7WV7qECC5IROjxGtiSs7ShoOQfxrzlHBlsJe5P9XzrRF+QOMp7HVdYn3
2OFmkvOPsovbpk+0TW3YxsLKm3BJaN0mm3Pgq88zf2qyS6tAqM++XnUbE4ubgsSi
JxC+F0Gm1lqM6My7qC9pCd3rWMzBm3kGB8y7pXFyTXczhIVYW2W4ox4EugLXuZTw
muFRjTsS2JaaTcbLmds6VOHDFJr8oOACo0kibM3jXOH2+zf7Wx80kidgGdEUf9Pq
amAlP4GPUf7L4VEYKYamRtzy4mVMXgSUjEio0jrwRZtCe16R8lED9rjivNrcIkGb
0I1eUkz8DN5r5L0SPtywz/Im7yiQ7+3ja6AW4peutrLPq7lZzb72VWTwHKya1ZdK
NwD3IPE19yN3ZjeFw0aoLK/BJ0LvUWa7+5tcuclpFRjvqagGL6M3u6eLd//SGAdE
ZG3gVd8oOkRtRmvxkrnjRtBlrfDELQ43yhhG/mVVwjHwJ6lLFSAtmAsqhk32Ghmp
TlM8GWF9Nt+4tqVXclpngTgajK0x1j1FSfwg2URsbtTLpFgI/E5c0qSREloqw/D2
oOazLecVH30yQuQNmdMWx1WKP3nXGkPY8HapdpNcnlYKHYEm1Cvpr1p5vB9F71yV
tbz9xS5oRrF7ks6JqAQ3mBvV5eFTYU14k8ZLgSzTc0CaAwcloyKIypqVYvgGQkBb
hjHP8Ydm+EWG6nkJ1XfZw0d0s4hvrx4ZF/5KThSqaUA7Mhcw8YnZE+aYCQ29HJeU
Rb6Zip7zxh/FisDQWrqnSGe1MjSBW+mhzUM/b3soT2y4ijEacyCIitSdAVe8SQr2
sAFJXfedkBh7kUsqaq/y3XEVH4MXtO60aeT4crRU/WoZ29agNCbJxMVFWiqoL72B
GU3WSSDqdeWl6rUW1Emd4GIN+IFnUw2AdNbuaXAzm2k=
`protect END_PROTECTED
