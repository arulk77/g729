`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEoN/tBqu+QetHQ0uEScY9pPOCh/XZfZvXrYho6xe0HO
8jt3GxaJhYM2V+40mgOO9aYoUxUvqCf7srahgHWc9FaRjjlsdQUPAy6Oy7vj9imR
TNrxzn52Em9qbzJFczzTlja8lNGncQsKO0hqHo7+Co3P3jwNwO/RWtx0RAFPybGn
zNppyH2Y+kiaQaJ4ys6coyg1KQpiFufxBrXa6wpHkrPVCxqbrTnN6cXX/Q1ht2o3
vT0rMJ3AUfiD3wxw7BSFEo1qZ/e3Xft30oke4TFOs1Hbg6XYGE682tn6Ysz7zid3
IC7zXLbuvQlFvYSMFaahgrimzdFIypkoXT2vvAmHE9+oeCf13wIKdtJd9bAQB3zH
I0k8JxnKtZugKgfmgAkMAMHbKdp6Ou3pUUd5RmXWc1yPYrADiZ3HZk8+I1fwALex
EirocRMTdsBTVQzOYu3Jhfr9n3rKle9xOSSN6ZDPfdomOOPE9MfWTHKBZBPEloZ4
`protect END_PROTECTED
