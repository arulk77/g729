`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Q77dS+QJNTc6qpU+n8RT+E+f9Hx7F9TbDclqwOtNYMKgTYGCAFSDOkZxBhPuCNgA
7sZD0B8tMo2y3SWn8+Sd73hyJrQFthmyeklEo60/ebDoCtmXsG0RXbYtei2jzzrT
Ljq3QC+v4S1HZOv2IzuSsQjrvhrnYiDBB+nBm3o229tHP33MriYFBJfitj5GaSoG
bmkJw4Ow794twMJWQj2XuoEUzRmQdg1zpOoIOpFgO9DlLQypmwAxl4hcMz7Glcik
`protect END_PROTECTED
