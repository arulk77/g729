`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zPeVO4HuoVDkYlp30yDjmKbvX58leXXUeAUmFvxggTD
MIbW9g8vGmpjiVrtB8UlMs+52PXw9LL88u40O2e6OUJYO9yXF8IgXB7KAmHMSb1d
XkbjB72k0gGlaHC6JmNBkZc1flm6b6Et8PFLXDjzLQ7O8sT51UErgulKLPKZb1mL
R1Z/j0pEgiLcTjqCX1ceQiGBxHTFE0rwBxE7e45clKIuWViiiS4zohTLpyugLbeN
LqUhG91JeJqxUzxZiKIM/EqoQ/Kysvhk+7kHSTyVaAL+txhKCh22+Op2sgzOf03n
V8xxXJ8W4YL2drevhHjCfw==
`protect END_PROTECTED
