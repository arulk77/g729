`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
YLM/ZKIYjcGeb3eZroqKE44UQ3zaKFMh3wmR+peXkGN65wUFedBM2Qg22iUPeRUA
Z8bVIZxzLpgLAUhDu8s4uNPO/NgEbWc7dY3nM/ShnSM64ED8ImPlYTCEmO2diCC9
vbCggy1BNkgLAftbhDczFX11nigqStuDZjobopYOPd8qvwXYLDPxwyyzZdADicgt
T5px9g2x3VQent1Ek1FSYcUVOuZkajDht9erLGiYjt99aBs1j5wB3LQ5/KAPMfrS
J3l5WkX9rmfUX5aJB1CzaHewp6PXf8rGKD0aBBB02T1iJw+ItTiqS5Oxb8cnueeh
ItfFRasnRctErpjASaEMpEqK/2oApsOQ7um7t8i9Qh0=
`protect END_PROTECTED
