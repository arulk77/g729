`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
lHf60Nd4CdEgafpJfoAxuojrXRPcE5B2HYrnlfii8/xBxF8tkURa8rt90CumI6cO
fFx6r+WIjFYnNm09LgI6X8oiG+wP4wJfQYBNCOr/lrgOf4L5cnyZkXVYyh3mpq45
Y3UcF+XfdERkR2SdpWwyve+k3BxATXCu9tE0g2xDgiyiw1fCeEFPolSOT3IaImKi
`protect END_PROTECTED
