`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCdrBRV5UUpBPFa5cuS1lg60/CZqC1iZ0U/E257injL9
lRCtsuYEN41dRYb93ms12FPfBWGJYbX4gxAGUnK8MWxeqjb93FsSxCHkFfZzBmDN
/ceMand3nvYgaCapzy0vt066MWytRRGJIcfoQtdRWXt0+ypzHkbEjEN/svMMFRBk
NnIXQEBtENgq2e4yaV/RwGrLmMp61AuRT4DF80cM9fZWZY7ojRf/4zu4ezCJRYmY
p3thGJQH+X6RW7lsRLMyi/ZzC3QDzJfa3te04RLBsWwv3h2cbFc2JkcqzAyCtacO
QU4bRM8szcG0uF57RUH8ByXZFrvRfN/S02EXWj2ogKNnGjqJ1UZgSVfKsiXW/tou
VsB8XKuFoZdOcM+4VyMMnWkCplBO4+RmEPeRU0huUHVz4JdFpzQfYz8Qoc4qsOkP
TdBEh1Zug1by5at43W9v9j8YPBhidMHMnnjrY5Y0x6ISvi42uyXeRey47qUXnw0I
7dDCBszHwdWjwDF+Fb0G4WRv35bqPoJ/r7KoGCHAPlsvh/6mQ+ruRcD4Ndnq0J9h
ecLPPDpACCoKBf958qrS8Q==
`protect END_PROTECTED
