`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOMMm6B02fucmTTipsDf7P948QAMR8kMbxO/9SZCTT6U
p+2VKPOoFKLeXOzu0Sdm/1ZJoewVREu+z0HQCYgRd0Oz796WMjbIQ32Ur582XUb2
0ZhhVg2ztNI8ZQ+X34BFYkkapSBrg/y+DZ6xV6HSBs/lOn6cgdpxUUWqtMne3AtS
WBl6JrP8nSGuw1pEN7OSFTOH7OSJ6EH2x9Y651lcA1IEcaJIAAwkVDxDKQtLdswL
K811/0/3hgJWg7X1DRgrzLflD28et0mnxuD2OEZ/MQoprEUA5otvHpp0wcuBfOOP
d71VG0e1OzljlQI8QtT5Ad7BQKYK9Wt4UBKRtXMEntNsHASeTuS5ingKGGcQquSg
3iq4/3nHwao78ZoIqvZf49rn2a/nm4CP/y6NKaSSrbdxIjn/vACZvzPsh6mK0Ev3
pwlwmkRYRH5o9Nf6YIp4dIXOhcPTx7JUgPXdLHL5BIcZO6LnmBAD7aND8Uobe6bJ
`protect END_PROTECTED
