`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
VN3cZiJB9f6xREOOK65F2vygTPNNKLU+fWf2xA4szITliwhhhSNlXGaog38FeulH
CBhHuF9rnZAMA+yQxrFD/8lbFfRe9ocobcUgFAMzwLqgZ/mZKVLyTYcAn12Y35Zt
xogJluCBMm8nT/hij2cnMhtNlhIUElBq+8phch60PqszBnyIYLgJO1N5dfJ9JquB
rLqwQAbAtSiCTmxfulOZBt3B1pN+kwSnzmMkcMoA3259kT+q6pgLzL6KlhX9bnMY
tx8ljHOc4H1Bf7V+VJylPOYqGrqXkxr8wjKnqz+zym0b1NQC1LvZklw72cUwNn1N
1V/ovHz32P4sVo5j1Id7AeZgdhBjUmVGtpI1JbJnRxTj8UAdqG+tzMDYrZw5XROb
iyz4PJP0T46J2iKKmtnop1rAnfHvHLN17KUK5QS2oDw=
`protect END_PROTECTED
