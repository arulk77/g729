`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73CyVmJgXCye+v4xqFkvLMUYJWrpijpJlITZP7fSNtoWL2
irNl7ViQYz0SulHol/NM85KYe7nsuno3HxbvvnjzERB+0SfZ/U0fpP61xww6P+X6
blp//j0sXFkXVJQxHnTz5I4K1/j+lSKxfvVIthDS20wO1wbWgUnpSUa8Ue0HDmlb
mNFgNbd8UdCjZv8hZyW8ImqQ7qVeJRzpiHuWWsiTWcCe/ETtwHVEoD+oIs5cC4jF
Pc10yOfqvrEZ796vIY28Jh6ptWs6NY6fwJ9+ByVr5AH+Vj41Sm1/+BDny3jVUtb2
CG6tFFT7gQIBZfwft8t9JagNeRsY58fVm2nGg3VSF+uhyXpPRMfopOz0SPdlk5xF
lEiKKcJ6JQUNI1ewBFyvC8TvsF+953oLQjfp6jv0xrIJW4t9yi8ZGqbqoWLxZoU0
a/daJTeWnxHUR48OKmzPXgh8cXQox8/ansdWFxLy5EfLM1VgnZICgJA4EzfufRG6
bfpSuKNv1wKjlS5KJgGHibh2Ij7tmsMfI6anlaM25622Zh2uaJrkdXsmPyE1uy5F
H63JM3ZdmR+e5F6SvqjHzHo461u6cJqG1Pue564VHDq8SS02uYPjilcjYOfukaVP
W+Cl47BFQDA7UsrN0ZG6LRqrXGlf1PmYiIKa53uEX6q8oROhOFZd9Z3i36V1rTdY
`protect END_PROTECTED
