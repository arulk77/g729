`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yvrGbk8gTaH/JqMUpyejhaTT/BN/IL/HxAAZuukNkII
5VmNCdMf1oxxLFOJMrBN3UwODcnv22B/4KaMH72QZOlZi5aEjwy9ypbNotdrxJ6N
mia3rubzcf6KILb+V792yVVPKsc7stqVT/aHg+HGs6PK2yaqRQR2hz0c5amJahL/
gmtrPImzyVXsHTkK94X13qiBtQX56OdhMurYAd8T26cc9KB8kKRU/oJWK9kNMy10
50Z+kGhTF8mklRoSz+XimMoYcrT3aOzUhAtwkWSid+/H5NNGpxK9vAS6aY3Qf7uV
bGvfEv2WBA24FXf3D+xrcL+tQbV4kx/oCMmNklNfd0Z0d6cuxyUtOvrzd3/tE4xO
yEGV9+R/aZBwgwcwSTs31g==
`protect END_PROTECTED
