`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAn99Q1t+J1Dt+4yfWcuodKLPJ0yRSKBShMzDRgKB64M
NIw+MMHlrLyVe9s0zqYhw5nV1KT/2wUVCYTZnzlaGgu+q0s1iinXmDOKt56YCmvi
YHtHnkSlLPZhDmblhwi/p/GrChwAr4Yg5bHNlxLaGcTNG+1Xx507FRhCcrk77uxb
lZSQAYVQc/gfUeV8Bup4I7j71gOALGbyr4SoXtEcTxa6y9w6DxT8VWn2N7HfNwRe
QgYSwtvO346dk7TUW/F58/DNaA+78rZfqKFwoXlrAZNbv4YsVolDlC9ytvl0R6tg
qbDY9GsnH5MUU79X3ire/SeXfD65/C6dztfGQedxWIuuENisZTIO+CmuRVRl5uAQ
fGsVJabfOPg0U7hAGocFRmDVs41ugvRytqsWhhYObQH8av+whYt0keqaNiRDFEVF
xS9On2Fvjw36ycdlMGkp8vcG8QpNbPrYGCESr0msKsnXCAAfee0fFNSl7jqpVLeU
6YgdKk87vgxQ7UklBJ7DnazFpNykxtKiV1XCA5eFGC43DgCNwtMtyRDqzvsM02H1
TyOkUZ2vyD+yXHEeCfiwrA==
`protect END_PROTECTED
