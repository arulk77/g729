`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
22Bv+Dk5PmBjPAHxXu6G3RB5l3/o5qkmgSoV7wKBB7F8Ii+qWlxtPpm7opO8UTCZ
ZUm0bJOZMe55TeO3ztkvVEBDYMdhpDC5KKt6B9aGF+yj6p5sdZNfmIjCLW09KM/1
3zXXOLILpUzIN6EU8Qw3kTaPd+yQXEnJ4sgQHbXcaeCzI2TDO1RfdyGo8v5mETD0
Zhnmvooo3VCgQnYv0rY1wEK1miWxjfsfHgp7F+K9F4g=
`protect END_PROTECTED
