`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAU14YzdXSuRm4LdFiWgfdPCZ5Bpqtzf8r2aYHBfLXt71
jnSMFonMqi+AbFOsAkWvv6CPdABvk/ZEdKOl164nHBPMpg7jMixDeOH3FcNXJigV
12oaqwx1wXamaXHnP4cA6s0jRnKZaaasLvPxrEdknlx5hG/Q1gGnsEKWESG1+OxG
R4pXaI2lO35jwt98ik+U/eO4qBXmjhdKwq02YPC7KZ1FLdjtdyFH3x8UtLkVkdYQ
GsxlkjMGsfH/7yCzyAf0MyoDcwwRkgUmWebMVUuJEGoFKxipPmMoLR2YPZovBlP/
P9sLrbBgWXK0aeQMivqCmmctZRONlyuCUTmNDKSXEDrtD8UXmgwWmJMqMeMKFzd0
vz4718w9s1vVv7IvTcRWMwCRT2x0rpsc3UDmXLlDMnhREfO5iWHg/Hk0/f9jCCpX
deW7s78KD7FPxmVq99lJBzwkZKorgGmZQRuZX3lTso0rCMCjgoc9WNXVAhTyjkB7
BzNLaqBxlLuMlR2ZLAxgaR4xXFJa3J53XMvQIdwN0h3YqiaMG8V3vTcMYZLYahbL
B+8KJPg6LBuMjMpXIcWy6PaH9zGXoeT/FPe6N0g93a/Y6F1opVPjbeSmx2T6pgG7
dfBXsrtm8Ab06aQkBZlcQFyCcZSAaFRZrTeg9x7JPl3IhzwqiMU21aLh6ZFXSgc1
ICqFCd6WvfNa4n0739QJWNsEWhdjsDnKESHd0k+bK26b8pNN0X33VLhePMWOI96t
sIXvbcETf1U1f3eIpgygeotObANOdJtRjDxZVz9pwO2IYxFUCXo+z0yqxQnoJO4U
xEtu0d+ivPi0LMg2pLiKjPZvltpOs02XWMKKVAgs8yoLvaJsKRm8uyYPzlqaX+0Q
YbpwmJBmfo5Cq/cVIaRhcqF18lzDSh+kvB4JDuOXBLnkzrwLzA7lXhMAFt9g4kw4
uaCSxWjP9pWnSpdIpGSfC/tKrFonNA2dqYB8DkAtOejU+1xODBcDEYC8ZeiexFMr
r44Wx3Y5Wk008ldHPWVQaW0vzW3HHaXw7ZXtn/On5JBMSiMlgaPxjnwr5fL4yOrh
OliHUytoJC1OYRWhr65SMTwq5/7jRoB92SAdsRCqesr+Wax4bz6DvaLeXINUcu5l
0tUgLfBU3XpsmcB9ozNoBtglT6lUMP7vbFqUt3CtiF53vHxSWaECQAk03qn9KCKw
6IXQPE1laZZNFLSg4BoQ1DSu3/2Ir4CwY1ifcIU90+72JNL0BTSsFjWQh0OUF8eH
HDpYi85Bho+cT8GYGzSULHwWy4K9XFsC5fhtqvRgFGlns8fC2c3qvVCABsjKgxOM
eLHvMh8fO6munVAxCjAiZ0FAL1mDA02pBKyC4TgMGOL4JVS8jT4SeXgN252yeFu8
kD6iWcNTbc6isu7516cJFPac612qhHIyGgH8GjDxMB2qeonABQDYEQihW64dwY8p
7TXNHz2jDsgFh1hEuFJvaJno5LjI1aG7Aaazkup58UBmVM84eZLNrN4lsBjNsRHX
f04II/HdsIxU82dFXxIgs/0CDfG7PFDuZ6EuGTg17gIaUJt8YG+86R3LOfc7PT7Y
EEAwLi9IX1G3r/ShyP8897cjXyph+fbrEfwRNCHqRlcX5qZ0RSKx431Ngh/fXI94
PoGfeGCtFmeSYPHu0omsKduof8HnrGEvvL8ZqPwUnZSEcIr7NuKuehK1dZLrr/cG
wsU9d5yx8Q1kszmosA2fLcGfgP+3gO0nsKV5Njf0x+6NiEE5kStarFtxW/2UU9uM
ONH2Rs6TWa7DN/kZr8qibUEwFp/UOedCZj04EzMT/zmhcjHzXRVUx+Hn44q7i0I+
6/v0xnOaU2E7SuPNmbiA1sWSFk2htQonEIEMsDhjpMxEpkYJE3zVDlASsa44gOVZ
rrIe755of0+OSOInZ1kWFGNxSMLseqcKn8/HM58LGtZahxlxdmjnqDEKd/5kIrkM
Ur42t/0TmyT1FZMp/Fi8Xs8VTgFe8wA/H1EzXheIWPHOwWLSgC/65PGNvNWQvtqi
v+TDYSVPrs5ga+Ps/GCIx3cZ7EOb20GT9XlamykUARGKFZzC6vJ+O8yj17tCC3fb
4uQG9XZlCwTUUmpuMVrUqrr8w6Ty1l1GLqAFvOv2NBQTdh0/8I7krcqHrPKyqfk0
x3fhThP1p4E9PDDjKuzoQaIs9YsbDRx7qrHuVbApTOYnKYxYKlf7kH76vgg9yKQH
+leTjhjn2P9zgbE6XC2KcP1eBmfgALlE0SWr7zlnuX4Lve8SRfbvEORL4MGmb3U9
NT///oMcNqgcW+DxErfQM7Po2Uw5MDv2QevM9QAemriCPWxv7i5Nhs51gL75BkVo
wygRa02SBTQwGO0X57GLOFJoxjMSwUbcoGbEWkWpYAgnOetZhOV9+IUyydh+DDkg
x4vztAUm0RQagQhMIRwhz2vb2xU+269uvAVsaaBUHm09viOB4dgmxLzgM1oH0e2a
SheJl0vwUXfDcOhE7zhas/t67V0p8QzYe7i6KrAutR5NQurabIaMNjrTcxQjON5h
ZU4/zD+RjHz6ZyM7Zyvhw6BDohLblK4Czv69cpBjzul6PHaNvudnJ2XdIlF7afOu
GpyCrPKbn8TWjM6yxhJv1W01j/DEZbER6G9DrW47PsfQF/M3hCKUrh5ckyjzv8IE
4Bgcdbk+wgPyI9YWmqmTGCUz+eQ96ZfjLSFqSQ0xiIXPlcAqYrS8TLye6eW6+Ps9
qmrn8LpMxcB8Kcngo4FxuyQdO6ad6AQkHrxdrOCJWoU0cciGKiYbHkAByhdaxUf5
Hfewf3/+5CvMuaqDZlk+Vfib+iFZ7lZDSodaOrRcR+1jrduWHgrZAClEEfPSGcYV
w3G85i9NrqozAY+Lhi42VxbH8xvrKTSYxvuWoZbDNqY6Ki8s10Hk5W0Au0fOislQ
doULc9E+Q/KjyvjKrwGmoLMybymrYoQ4uGQN1F4YKjDZbEvM33R1Jk7Q1UryjaKA
c/kN0f+0K+yaRr4OsBmxE4ZxpktRpMOF2JWfZ8eIppoPyZTxMQf3y8bKGTHkN7YF
Ehy0wRQANhReA7y/9MySa9do43Jw0jZLo3+4zbgc17LPajkN1weEntDqnv+z9U7O
YlY/+NEma/j7DRYVoxVr7opMwvy4vClOWzrCS5TchNzx1z0xAd+6SCxp9NLnyB4+
jGSFN6n0GO7E84+am4pTduDvTsj+V+dpHohZ+IOGsWIuwvPgGt8PTsdWb4q2iXzI
VCkbnz+YjCz51qcXsHhkfOV13uI1Wn0/Df7MwjODUE7XApc/0BLKnOnZoYVtUla4
TB/WnD6SuW4YIwpAMxjdll7osZUnl6RCwA/fzPty3L3vBzaBOEcD9JT9V6zwZDW7
yPlMdXmn7R7Oypb4UqHxkpV+RQehYIBnMveK6wAmY7+/5pdnNHUsarkKahI+WTZ7
wIP3PB89g6uMonhSrY02ew==
`protect END_PROTECTED
