`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
/L5JmTY5jr2gbjuyb2E0lj19m8uWHZBnhliNU/PL673vrY8ZCL0zY1lzyttSOvXr
CXKadutwdyTpSmWEh7TCAJ05R0f1MbiUlhtKSuQo4dgWZ0fV6Tl/73hyiUhCvxKK
lW7G0TNYyek7QBRZhZH/1cwG9fhn8lFnMyYWbQtm1GYnRdfeeqUu+5gD5Pw/7NRw
zIqU+apOTamvNH+urWLxfpouqqgApxLR/eSBp81uFWeE8BMzyYqhxen+m/2RktVe
9NbdZ6vP/t9M64puav39Z8xI4d8fXhmsfYYng39SZaa6ulUKTG/ilR8vgfE1aJKa
`protect END_PROTECTED
