`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aQ+vfcmYM8aqlh310edMgWlveiuq5b5gnd2YwsqyCLBv
XAxtiXNY3BPeZU5bmIWttqK9KGzLbDTzF4/CZElCtEyWRqboMOuHk4GYf8lgcYB7
Iu0NTw5MNReW4U0zo8b3mFAoYauAu1H08yJ/RRy2DyjAdJYFGEbq7LweIVhcZkWd
Tq9bBQegUYlSeZRqFZSMKPA8Dr6Ot1UJ5NQGxGab9cImLeS92QKmqNY3mCE/HBeq
nSzG8td1U1/gFBCHrgilpq1/hmHiG5v6w5rWz9r/rolL1msPQ7oO0GAsi0LBJYNg
P3pWZR/9VN7Ae5TVUppgnKpbdF/bAObeSWyCEf1w7E1iuiDht5eVwMaVPhxwRN7z
P/rBXRY8DRFJK1mE5zbXsDXQAQT9W/yKke7zWWH6XRHWouAtJa3/xzLWSTGRp4go
AljimLGc/OQ+Kz+qJHrubQ8cDrjLmlWm0oeRnFXp958vC9dmRJvGIDGS3C88ItwP
B0Kru7OQHOQXXkejeaKc0oucx5UgChq9WRucd/bvrGGqbn+2geGOaiscNagneqjF
Uj59MOdDCV9E2bXh6EfJjb6Td97Xi7tudxm7gX/2EVp45XVUf9pxNeVVS7v22TFO
TIXfqFXrt/rrr5zVJfRsYjV+0ypcYbQigAQW4mvwdsx4bmjYwL0o4KLK+mwPR3bp
d9h+WZaOgHy1pw1ouzul4NWIfd6IvMUcROwdJg7lyf5zsvFkqZTnNpzTMigv5UwW
yQo05RHvylFGijfUVFc+e63fbL6S814OSQkL4/0FW+HGXl95IMhjzveRVu6sbiD8
Sax+1MPXiXTye6PUkcVelP8gBqdmdNw3vINOzUk1zIwv+ttNPzqnDEaQ72rezy2a
ugucaNUCnxvHg1QZpoNQvDTkQQVZe+hgV8u8oWxD9OdJBB1+/tPCiPIJ6a4nZGcT
B0d0lkhU1ph6XC59G7VT1jjMHH4xkfKmmnyHEUaThVxsgvJPaNbL2Cqx9iFSZ4on
sPX8znNSEyTx0FcIBRwMSR8uDmKpjj0RPUixzK1SkgMppCSlxaCpdUKsv4UR09KC
hTq/qh8jNsS0mfsmbTaZO4J1TBhi7XS82uNxSpO2mxUeYWueaaOT8luZJVSylQnL
iU6W+Japb3rGc+WympTPO+URbEEsxmDEIMuQZzsO6V0AqYkare0SFu8e9Bia3umA
CgNY32fiIF93oXiWuIiJweVKtWDQMoNFo9xTmtRJaWTJzcXpje+w9Gez4oLofvA9
by0ulN1JDkg4XzKbnpSeu+RgUKbfwJyAJIvi6k27TD6asUQ++deu70kcGQU9SGiU
RMXhyzEmfQg23GImlK0vzHTTPGw+vTqnvrWW4UxZ5jO1mi5U7LmqwbxlKp4PZd8w
Dl0dTSbf71MgCrwkndpH0L8nlO0+qTB7lqYijWB4P2m5mbwm9tw0rAerDJmN4r6i
ForRFuDZp7rLtZjiIUKXzv4n3QsS7JlQxCg1OK5azZWSbplRANf4lgW1322YIzXS
RpcecSNhZqYdpVxYFYmbgKBtscxD52b7HtkQTOtT3imCX8tQ43lkH4fKJZ/76mw9
PHFHU1YVkw/3ZsMiJuUtD6n5dFGSscCtwvGPK0oXixLf2dg9t4jZ7nxQKq8FlC9R
IBO0Len5Ntd77xi9dNEAIYeVy+3ySMWzf/2T/jskd8uNQZHgk06yx5XSoIt2Dst/
WELQHaByDH1oCKI+b4wAtYQF74bPxuR0By2cX7uhkVwNXlOod5PiJTRuUxdHARqn
dtmA62R5D88UD2DEn6hAPiDkLeP3iwqsVSMF7qaVS5K/WgDLRq0ok1hcZ2kXlth+
Q6fviqat3QNK58RJ+qDmb45vWWHN6hyOYKKKX9aeaYWUH47o2Ig1ojP1naaQZl1l
5Fo+zQBsPR+kZgp2MiXs/5V9pjQGM4y1opG/fblnqwNr170esv3P/R5JXZAswika
3so4zxtggE9Ppmi7DqJ8JLJ3uI/RJhsEpou6Zo95QNS0+l5jYgdfKKoKKLTjrVR4
U/RKPsLp73Ntken0Pieh7ZWvbNbWFj5epMpHqBeVrH21cCjjcF54zarLEmwCDkE6
Tdqqv7XATo9upc7kWz/snuaGH68xHrEZFtvPf58tD1jHGuoG//d/ED+39+WDIt1P
/wHv6D+NAmsCyRbwU8XYRBmd5JFgcdQG10lWw3ISYHvYLo/BKtR89k72OSBtkOsh
Rs7Q4dDfkW3OAxWrNvFaB50fz+tj5Eay/Yibln9rEgxPWBPNdh1197ms8abnJGIM
VS/OdU3Pfx7icKNdKJ5nkW/tqq0p86JzQ+PL1+QtJv67wACWa4Bt9CyfdbhIfLC2
XVFb2/yS3VWFfYzg7ojh5WdA+DbKS8HYrVdaQmdQlBRZ6rtLub6yoRHNSe2Kw/fS
hzvD5B173eMBjCqblvJlEhN3aYRiJKzYNZ6thu+wXrpXoa7CvBm3U9wKz8DU8kQ/
Qyx/o3E4z0iFi7fyciPoJDbNzIhDC5ztKWYF1x2kF1NHtxPkwHdPKiSgM1neppiS
RxEdQ0pRnqeO07RH3GXMfyK/VlJtyPmuOxXw4OsG8lfDApwgo5xylNkuGMQxJlC+
PDGPCaKXxAp8GTVJMn7zq1s2ZlEnoreEm3mWxhmxeNJcNHFi3TXbLtwzgacJypCM
yglxjrJNHPhw3xTfHnrz3fTfc+NAjWV1kHQuDvvH1iQRO++MBtlUZcYYq1Cfr7kN
qZXJaInRe9GTELfWctO23LkasHWfjnbWj9WCYBPHSGJhMxi/RS4EYxbXqx7BO3t7
xbIKagFkMQB6LJcix+8N0icBijiH8Nmq5B8WIf6dh3AcTzDsaB/3iZmkTGAXgHNZ
sQnnmR/Dw7KuPeIIDhTmvIwteukT+iOEuGKPTdmPj9pc0fA9kTKC5iqJffDkaoM/
9tth6gaJO6p1cIZ7WGWzcc4NOkRqCnX061h4aQeRjZ2NPhX6vWh55neHLqwYI1xz
+JyRsB2wdn/fCxCm54aZxlgz3TwJSC4dq7GtfNUcsj0Yck8tnuU+NT/SJrAbCccO
iD4zPwElGf833h8E9AOs8AyhQv7rLfoMKFHJC+Ol7Q4NtDbrJjGSFcnlpS4MeptH
lYyCsWYCdVJ4Ab2VI5rmsDHVsRdZ/zbuNROfBs3HVlV7o8s/P9vvrWrNTZGbfjy/
VdvgMf2+SOLfwaELFVXs3t8yXuhkgf07eDtesq2LOgj/hfN5Hrr1VGRWZ4hCAKRw
eCOPJ/ylPJIuJCEURaKNP3GRWOlFNaPAonvuKPeIGxQCuqELX5L5DENKUb4BDkbn
cEGL1/uB9n6RWsShqgNAyzyAoTVARl/t/o7GxHD7+Ure3cqBA1oZ4dkqG0C3bf1w
9KLjR+d9ln5aNb5AqrNdMJG/4rcTp3+RzljqEwoUpwVdQ2wCxKub/VEzPFEL8dYv
0rGnqKj0lQq+n/R91dVFeIFNXcCT7ll8twRosuyERsMutfQgCyifmUj2wxiqXNcd
DqgjzzPRhZu0NK0OzQxy/vKzLrAEztx+AW/gq093xT2/KTKXc4LQn+soEJo/9CUj
iIB65j3N8tcCGAWhx2vKPU7ShgTYS2kX48Iy4Gk37ZkTofbbxHqwftFnrBsSO87j
/Y5SBlRZHoAPTDnY+DD0xD5sRsUsKOl1j4l364HWAMsLj8k8Zggyvlg4YdM8No6f
e4S0235C+cGVtGK9Pb7p4Ng6YyFGD9SNVw7xZDNPHCYkR9KIqmiuKiKgiOuR6wj5
PeC9+5tUlKob5rWB15NSKmfDWxQWU8F5yF2K65kdLNcnTrUU9nuNFEvDAC+AZFYT
HT+xy9i9Nq07O2sIMVyMR0wstZDWr6WzNifFVq+s1d7/3aZl9i95yJ5fkURVvH3w
434fcrJsjzNjUNClBhmv4EgdI7Vwp3JiSU6oER0lV7dejzc2B5SmkhFG3QWZN+Oa
oXmrqsvnCuvm1Qtpq3Vgok7mG9rpcGY+07WF6yz0TyfmGjD1bNp0i2ZUVReSBqjG
YEm0JK7i8kdW1bnZYcu+HaGU3LKZhdFbohswpTe7w52bNHfapX6QPlE1UMejb9nw
B1GpJquYWGzMSpbXrV/Ku4qzEblUeg3Mvg1tE9TFKsjunDrMhEFj0uk54/1AzcRR
EVFOjj8vgOKYVPpvc96f6cfGo9JGGMdqilorPnhX1bew+o8V2CsLs5FK3nqQcEeo
ibvxMPz8Dk4nJoZpUo8Tz76pCwgqZYOxJbegeU2twuYbeNXfmnKHL2u3aAJTerk3
z/QDW/zdThub+arTZL7FU3/IcP+HkJi1KaADLtDp+R8BJRySdDznDqb4Xd/8lYtT
zKfrFKrSVAMps8occ/27V4ZS4ZHMJKck/wO6/yjO+anGr4RxpaaMrx6jVQlfpKc1
GDRVzR1icmVX+Vor4iAi+SUBqJ8bhke28tbv7qWV4EupQFbRctPdBWFm08aPVZ3E
HghcDXTruGe/rV7yG6GxzRyhyyKvLei0lINM+ZBenJYUp9xmu8xLfW9TMF5ZoQwW
OxAvK8PvNBB0qH9JlGZiIXpI+nLPloP0I+SSym2sn4cv5pnN6mdWJLRSdBDtB8PB
6dtqFKQZuqXX179vJOsPaZRewbngLuaLrd8d9VCUZuS7C/J+0kbnjoO9BHaJCHpH
vBsQeuy3btQy8oF3VV5pyaa9UfLCgOOmIqHfEechPbfsNINCtIuqviyK8bWZB7sO
o+wJ+Vk39uPfLLycg8IFqnBiD4GTO1QO6yaRmuq/i6l+92IgWgtZRMl8YxYwZSmx
ykSym/ICeF3GWuvL+8/QaUXqNQXeSIg3pqBGnUEBjUyl2QwwavuMGAKZsa2bZtVC
RAQ3zvW3LZiz6TZao6fYD63xLrX9XbBgzOdWKLGTyBSZAIao1xNweEo58Ejz7DNW
0x7iTqBx6ElXrYER2r5RhyYIhpEmz/WmsLe3BQAxhdp33uNe55cadWZRtmqmLEpa
5hPRrTqfB1O4kzfonO0JoriezjedfLA01RQGhzo30ZgRaIGydSy5YRQ6lBfjpcnX
lL4QouwKJuNW/BoytH9lvcRy3cmn+WZpiVRwPS2WOwfkN6fI+m4SgwE+lI1BgSH9
fJohs67M4vKx1+mZCZRQAv3sgvpixiTA5iK3yY8eUGVtDVgo1r2E21nRpgCLUWRH
KjFY+IGVAcvJ0SSJ+T58Wq+GEgxFjD+kmsjnO1wtKmM8O8o2YezpDr7Mm/GtOiW4
/a5vEL0hKyXUvq2wvTHGstdMVVu+7i51gd4kupKH5squPV6du4rV+bEe39UJ/PUW
9jDo8dC0a/5HJSp6lNpzho5gRIpjzQKl/kP7vwYMc386DVNOfjeo5Ej4+kFgyxuQ
F6ciw33ZfRfMmo7wvJn+tcatwhJgdwVeuxCYHAD7dSIMRdlKLFhyMMJ8Jhv8tcoS
/Sw9cVRXGqwgrxOa0Z4bulU99RAlGAl5JK/TRyBGIll+HshDMSkkuA//+zODrQ4/
Yh57A1pW+hEEKfY1gD06rQnad8W772XMLUScDU6bcbFtfpeUk8mXtmybI59Pso/4
Xuh7DqktZmyVaMYQvlhbLQrp/8Jmlzyd2sOZ4wbTXgBwyle1brHJukti4kN1ybNQ
527+TtPtYkAqihFpvplEZkekgighbCc1h3CTXFqWfqhXOzzdJdNAbgceQw0AAlEb
YHy2mZxJUKrCNb0mTLgRTCFTgoVeha7rpdrRe1VnGwgul9NZlRPcD1X9hRPZruQZ
ro5Rka08MQcjCkT+imQs4QocteATqg1ujo3oKT6orOjA1+LQNLLrnaPdG6/+Doqj
cony3x83iXoTDxdApJPOoCaCUy6jF2knrjwwGAwUA6yUobKwXiVywd8eIqy/YVff
lnfCqC5yoALmMCzHtK4T2kn+bkz890J+dF5nW2YvRiJzmJzCfpskYCPEN6iyMSvv
YMSVnX1dFmNe6rnFYbk+/+UG8rCVS4HB1lRXp3kaT84QISgwqagKHdZF/yaig4mV
0/QzTVoONarHLWtBoJ/mTdtUHAj8b7+lrS9Z/50LqtjPYtq4Z9xV0mSUCBsVv1Kh
JOxkbnQd4Pwikuhcj7YBN38ucCN5/AjwZmno6ZFCbYvSxeKPOoGf2XvQr+0/szKt
gCDKY4Tw9FIhq4s1k05S2u7/Keg4BQK742zgV0ezXv8rjdYfA5fr/Bvt0n51q1J4
33zFSq7QSplUCtsqF35p48Mgp86KhzPM3N/XXVzrkb75SBvtWGZf0AsNcFxsZYzn
Tspwyi59ZXl+4dsNheRT1Z11qrVZP1xThOE0br1TqPTQb/xWTj7BBLWw+bFhRzSU
P3Dlb35pmIF9fSqcK6n3JXAhHF15QALGS6gIkFEgcgLibVSuZ+IDHGdM80PHGIo3
v3J0J7yDWT3plW9j/PAsJ6vZqw7xNtNJOiJLPVbRMPC+nMzYbV6JWF1GARe2PZbG
/vSBAcKqF+vl9DlJ+s50JKFmermwwBdro+GO0v3tQo9vFCsvD4aWxE4ZgUgK1aIy
IjO6njYKrgZ25TdGVwpydCaHxot/q04mLGbJANwV2Ms1nYwg4x2fgvnyJVkYm0tB
bWlVMbr1rT5EnHtzp6TV5mU7dwemBsXcIMQQG4SKQk6bGxiQ3LopzoIHFoqoNs4M
EpAcEajHoQ96Qd5ehthkwryBPwdPR2HdEvURB++9dBoHQIG1m0CHWCfRttnj8NkY
iJF6HGOVLgqHRtpmg+jlmoLb1pNQt20Y3ZU+cx7iRZHdVn4XL4lqI2U/PANhbipt
nF/2mg38e5ZJqO4Vov+THDYNjYdO077XQVZX5jJjJKLJWVYuGiIGkwgVxUxCw76j
TT+OCmIm1TFS5WabmdnUa3EBRDbs3uE2h3cnnswbfytiXVkXaJI8lJreARxbfOGG
pvuJ2LV5+j96CHpUWKUJDD+hUgTQZfRfiPYeVuEMXj1K3vKMl1RIo59Bk/2CqWUF
BRkeDbOYmohwRe3C7204YsYlo0VOeGaWUIg4H6hTDP2U9+ffqzyRuWv1Hf4ZeQrg
NBQtWGZa7irhIs6KYiDj9iiWk6jLXP03Ze03yZ4+dcAgaIAH7rlpgXWBzuQAgBAc
ulWfGtWCa35M4d+EiPSnOFiJ7NOOJRzxSovfFff5xqXWgcMN74UlTNFmRrndGjtv
RcA9EUeWyy4k55p5JRxJEWzpN/TCg9MbobgGeWAt47oBZMgH0pwPEXhlf63Lz5yT
DaMGqqZgDwbPX8ImG9lBDDs2RKlhIKN9CA3oqJnv1yXzlIPq/ndKuBZWTGV9cLT5
MYcPLD9w44or7saCehdEQlJ14LjIzQ/UgoWcM3j0XKDFdGrgWbBYo7+4w7h8lJMP
sYHkoOAVAX62S+l5wt9JDtFR4mRCzM4eyC4vPjLiw102fcf8LUV8rN0Cp5WG0EEU
uv00W2O5F/nyvC3R4VBXVMS0FXPuFvi/QaAvYOjIxxF6+78JwyVUt2VZ3zO/FebI
3rkve0SiTYeN/JU0LjVdjgtd7kxE6tSKnQSQOLrB4HZZU3+VcDIdT8Pfwss6nJIz
o0Ktkv2htiiy5vzrIK9qdDnAM/v9Vkh/B8j15E7TWuk14laKWc4UFuPxyQoQREU6
XqicrW3vvMd/zTtJsxrX254EflIfFhNEjBnvi0qq/AwbLPVir++kQJX5r3EnI8R6
TSy3CpkZ6RB8k0sWIdO+pdPACOxnwtAbbjwwRmMLqmisCP9CcuCU7/E80cvf7BVS
`protect END_PROTECTED
