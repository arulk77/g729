`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCpZpfC5tjNHRvVLc8kXwKLtvowK5+f/odgoVUuY0ORt
IvV94BL+Mho/RNXqiM2N7FPecWc+CR3Vblh0egqlbL0XV7w5+OivTdcYcX6LZo/+
Q3NQY4dycK9eCCFanUvfn5ZrwdSEcoku5i1QFJI1Q3gFwXvIIGT7EHnDya0tzG1Y
AV6WrJ9JC3FYcdGNFWJn/g==
`protect END_PROTECTED
