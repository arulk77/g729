`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCEXLCsSwB1ILQO1cZx8YAUOv1mlqU3H02K//MyPNlSb
rxHA4Vs7iXv7XNSpczllxWPl9wHMN7ezZN17ZSGgpRTR/BmSrH5OJiAqXUitKi5z
XzZOlL8AjmwYG9LqhDBwpFfUsCVghct5nxoechrb/AG7V77sGPuNeOXixQMgND9q
hNAXdPJ08DwgwN6Tpjr+DVE4SqIqJDfv9l1ukkpdCqQ5smypLLmVGZRq5LSVsSox
2t2ApaHYlcNaYP/yNKPuSGb413kfp++yLVAoYuPIzcMNm4BsfIYuuis1vhWZ1Jrv
NjGekQA2qFCkNdWqyfU1EYGSlmBwud9aZSOKwrHXtxHi7sp9bSAAuyFJcB2aZEH7
VoF2oYRyBwlC32sj9POdBONKAyOljhJTuC6In4ny0F3fkroa2iUfpIDFJzekI8Tl
AFZ6uAsySYRg3OvZz7Hl3HY+QTR8Y9F5sefTwvjp1h8aZEvmsCdHrGbNkjRUp1Uz
Bhx6bhlR+ViRpIXPBZonjg2+iBgphbbDgsA/zNxUEGKajxuCxl4MIURqZLNwu3CV
e3062cR3h3M4ICHhG57bnCjCuTyH68UAryoyUYsw8wA8BA8XAKh3ozUQAtgwyTld
ecfKZx3pNrhq1kbAFGs/CFEp1JqTHi9/kBD5i9J4fBJMiNMOu+LUxv4UHi694nKB
XXaIEZv06vdns2EwnvcpyHL9URkKr+Tc74QQUOancztE2HzCaFgIHUQ9I3cR971/
sSXnudFXZxIi2D0b1BpsFkrUBPM/ZWS3pY8Evkfux1PF0pEypipHQdfEhtUAG53I
/tzmWsbae+CGwswaX1/WldB5vVRfxQJjfoQNRC8TIp1/zqH7IrRS4FI4OOHFA3Ii
5ghiEJCjsuw7UUtKqvjaTiOMIVHLKdO9CJciR62FqQRsD6S2YEY9DIRjhuWqg60S
W0g+DzR7PsR0jA3+dzL3ivqE1d7tNFSpDh6ciQoEFYSGBiRVdsRQx99HSgfg8KY6
WQo8zSBV/giM8qQZqM4tnvM+0KJLq820z9KIIlfRrHqxtuOVv9+AgHvTCSs9VutD
ZhJTYhvnFTwYlnppzcpXziWm/Rq8z6Y0X5Ww5yx7LbQ3H+ONl+9yblyMvVTekhrH
f2mkbV8BvZ8dtup/RLJdKKAED8X/zf8G9KQpPwTY1MsKenUpftaCusipBTiNNhn7
nSqM8BX1g+H9kwLMz6UuLT7w0B1Tl2FGS2JhvCQfbUmQsBe4dl+RVRq9uVt8lsCK
aSbbaWM1Sk/mZOVR50ZHJimW9dBnLECHoEgcPfRNll/WhN2S49manBw4ms7Wfigu
8JN+DY3yw7lhuIomnCELfE/xADmQK4l5JWz8+JR0+BUDh1AGNXUlC9BbCr6qkVoh
yc4yW5hc+zxCKNd2Q+ys3QuAMeTK4onKyvlVBCGCpk0wFCP57oz/4lnklzZPQz6A
s2AiHZ+rQOMzDzKSVp2TJ8tXqG53qN0nZvvm9EOGXkAjsrM5KzDpoaPIr32H6xHy
3rzO90zvlLvqIYBhAvw3sXVf8dZ+6qLgy3laQDhQRi/rtmwYXIMUlztdtxjrCHax
0ruFcoeogWpTe46g3/CSDjQ6+8jhRQ7BPkkTAccmz0abCmnCHDaZ7GJHrjSIQ5Qo
7TXY17wZVwN/K61ezM1S8wpUrXD9Pi8EW8W1N0KcfGIECGPZJTaPNGIzCbD5PPCH
a8u6bljH5i2YtcFhSd2+WeFgLeITexIn7ThgU/BsYxa0ygMpkAqSmxX2RsvcSBwx
gJ2cVKLvdzNPMn2e/KTbROf1i6v4XH+ksEFR+2IG5KxPC9iNggDjehE8L0RrnAoH
t6I93+QcpsjJPEqHp5a/yrIdfVodx3tlWOqSC6pfLMnYC/cLZpgxQFbjqNpHxBJi
Uf7NboKS8vU/vgOsMpLgpUQAHTQCGf0vWAODrjgg9Lax1v0Gun7cEtGYsR4G3BiR
PHVAwgZK4IoOc+JaLx3jT+bKYV91DDU9k4dgw7uSlvPFHPfo+600RYtDVRZhSpWP
nuIftiCjqg+YerXZ1rmlADjss2jDAj8dT0+JUlz0qQ0XvAQN4zv00w3bk23r3ywJ
myXYUO4sZGAIrdksl1o6/a5X3leMlIXneYyhRqzT6Ucx2tecQSoZxm/txP8abvul
SrBAftyzwkY5ihCspP13LhOM+iIXe21hg9uRZ8w6Fnu7R7MlA4bWxhuA1/Guc62t
rANpCzb/VPbmFJh6ZD8J92dzMvtVlKg8cqxUmlsJ6vGOrYQcVqiZxI8KqYj16ENv
WcJ/Qk5eykoPbY17tLmCDEWaKpsTlGLNQOCi1EMFrnEt4lU1Zm9g8sctGUr7Y3H0
b++MRd7IzhLiu4mjEcwXvGYBedcLKtX8wDyZkKrhi7NfHENMy/L9qEA96BCJkzGs
K+H1EA2nLXdKwpCZL0J/vIM45ybJgkebNDbcAapr/NqRLAfIL59cVeTDyx3hrc/g
5yBJLFm+VGPA1F1syCzm9t2codPJEhsR15gpaIvKAcTAyzG7VeTa+5DgZe5IZ9FT
49N4o9cTlgFFehyv4McG6SThzPOSmcjfzasRNZFSs0RVOReywAZB7ydz5IlmytHH
Iuj7+XC56FcgtolH8ZrASuGJ4fE1EGjPAMJipRpR8IuLqEc479EU0QlOcevKTt3v
OS60+HdZBKYJBQUlYOngOBppxmanysBhGoEuv0Yc555653DRCnPHzpIIORm7UR1A
5Uswh+6NtvCTxPyQSiOO6Xj6nHrJxJGnMlLuFqIjhDWolVk+3vVvIYPT5zhDgvHW
jnovj1YFPFxRRT0nuSUsBA4QUy5OwRpRWPkA5jQtAOi8xfNg+95pz0o/MdcMPf73
1PJs074rD82jaxp+llO9LhX40TUbQftnAsMjtjcdqvCj1+idwx5EZT5+oNq8415+
vrf9Zk1yODalGwQtqe+bNOpdyRTmH1XcTQOes22QkuZHSMAJgkurFHA/E4FgyaBY
zgKj2PGSB6sttfmaOKgwhX0juftwm6YmR2dTaPZfVuLh6cePS9ZKJqIt96rVVpWn
jRb+eO62R32UvteqnfzbV43AjLH18Yfa2i9sTfSpNbFkgNg/3kF5UVjn5Yv0Lzft
0JtLOV99g1WM6+qVAdXTm9S2ZUc/bbf3mUkh0cai6RQ=
`protect END_PROTECTED
