`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePCeMPKYL3S0p0Gq34l7QofLnRnqnpxjK2bspYUCbeOF
iZOzLs/Oivn+aKT/ilAk3q1rJ4n2aoli7klWjrHR/ihvJ14a3oZiHXoQfNjzcRUD
SXPlH0sFt+u9NEOUiPzBeO80rJ7SMNurfoYwibK/5I0IEADp35FZZcz4iwWEYQQL
l7vyRoxlFAjQ8IQ6KHOe5F/L27B5B23yLUlj+/IiWOTDjY+BM4pcwm1yMlldQVtg
KLxw8XJj7d9m5TxDXxLGfQn/LfVTscsYq45GMLrKfGEWNpaZr2YLz2lP3Mlt7LkO
WuCTRYrTnDJb972yrh4AqYzAgN530uDwu1e5xDX1Oh0I/kd8Vp6ZfEkEv4A9TF7M
JEldJZvUXCg1JyH6gcc32ymhowdc5qRjKRNyag+Hh6nvVIY5kQKuZ+r3Efk2cSNQ
091WedHCBGtUAGCGOjmzcczi5OdVLTuBX2gFdelu0YjIAtFAvwslnFZ/TJQxknpR
K5x/I99/tXCGuwZafrh+wdpkUvQHTpZHUIOg53wzQ6w9imicNUTuSe0/QhZAteZ9
+mEAkLncnvH+DMv9bSFNxZYg6pufRYMLc7rmqvbZKMmtbV9QS+6ZDCnBbmlS3s8X
Q+6r/DPBKY7z9WnJ2G86pTKL+BxtJJNbeE66ywyfhKlrcdAqUfpQSgCwEUqEzJF2
2DTAVDjvKSXMB5Htkd2SPZm2xYLUEIcHjjJ2szH0dEP6rsLXe+dVMGhtMBto8Zw0
RO+4PNrbGK9+bxUWb/MGe/xKRWE+zXVx3kp0ZLR6bSti74otagJpdlw7/XGw6NLs
OTvYCVNPk2I8YzM19cerCy0Xl8Acdf+a5L0pabIiLhM=
`protect END_PROTECTED
