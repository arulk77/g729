`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIwv898SJw2HFbCM7TCXgiesc14VP1uuqLdBYPWaY0go
t1c2NpsZP2jicW/GghTScTSXFQ/Y7kveh7Y5+FZKaEvZB5vLfbcN0tgbUKDZhl53
S80v/yRLl0Fth+rY4ZovQynSy8OMOQj3mG6Isqh9OmcAint02XF5x4TuobBySdDD
dLde2m90KoqnlIW7bYp54jTOXwMJ8bhv9jEAvV24Ccfup+zkReGjEELJa6X0b5Ma
XL7PT4OKGS+Nla8dN+p/pUv+tHqRMWLxezGZkkuTeaMIFwZLQ4LNGB3XpyMJbIxg
dZI0GWG5JBjIsogDMYLuAg==
`protect END_PROTECTED
