`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
d2+PkhqYXchSlHZGyBT1JObCamzGhEHjM/2VMYT74IeMf/1MFMkxdUUpJfEAlJq8
nhlbrvOdvlFBaGc5XT5o/g/emHlGruClkBBcHPeiPYWxa6gqHD1csutfojBtwym1
UR6Rq5/nDhalZGkmqa2UOjN9lrrkhm1xJp7geDCbQlw=
`protect END_PROTECTED
