`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu496eGqeNno56pJcjpmJdmIv6jQf6FvyMGYaor2FvASve
c8gsr7UkuyiOrkpVRkP3UO2at1dtXkwCq8O7nXJsW+v0+Wi9J9V7znltq7Q+1aw3
DKQlAGIrb+9wor3ba3pQcl7Du3GC7cXFJ4UQUIdUbx/IzjvuHs2i5VzGT7VjezHz
7NNYlybhSIBujStCi1i4fwm8d6bNrZTgH06et5AybR+bX77P0Vyy8AQD8ACKfJEc
VxqLTY2z4JnSD6Mke0rWOWY0ZWPfojAg5i1LOgDo74A=
`protect END_PROTECTED
