`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aSd4MC05Lvq968tL3kNORWuLdXdnGpzr5FSF0XOg8C/3
82ovJmUUNT2L9yTmZUHGxnBjDJDimRTqfwggvFmPv0jJhKVFU53795MNh+MsnmhX
2ybiXgdyvnbEfeTz0CDUrq8oponvVcS3oeeBkR98iBTigeDkFgnaCJnkvfgqPbeu
5xDqtZY46FyeEBsdilAuVhe86IEikimPnHhH13PjVDNoNj/wmisXBrmQY46YZRxY
6Zsi+OnoCz11EWJBcs5x21nFSA/ny2S7FRh5sp6usRohiOAyM0lpHp9tabtzYVeA
TgDZoqvNJ58c9e2yUWmdxOSqPoxDe8ow4WLBB41VTcG4WP9UjozuvgtnUpLrSFbh
zG6QLxsh5vYYUjp3cZ6/K55i6JHBM9Z9eeaHp6pLa4tmBbyaTFS3EwRcFqVueLA5
hJD4EExD9BVSskzs3T17Ms/6I9N3ndilFAM4RTkQ5Qrn9x5H3vDM9eich8duwcZ8
K6htTFIvRTwGJjmgOHt2aR5fuZwO+PgZpYAqb2AiQDZCAcTFObSJLT2wsAF2id3u
gxJsDw6vpV7WY2i/h2uVsNTLdGqYNiOBf5YQQozn6U7/ZK9jMImmEnTwrFoXe+Ek
tGPCkQnN7Zd2JNgJgZMq4viR32gORfyrrx7PJPKiFN/7hnWBNCYwxxquNcIB+xA4
1SIBCukr54Agb7XEb4/thJIg7YplqDjj97fw6BJaxHizavhMHDsmC4acTm3jOThy
giwerfpwuwH6RHZiJM80DO+OxJhNdLg+jSi5tuZtgyeb7/fYoRmTJLXlGrsKqClh
sRLmt7RpvLvwCTWehS931H9snWWs3EwhHoBi7zXFiKR/54S81PIop0LNr3mDzfEj
Jpxe3yiA2jOgdQOyw9gZZ3UHR/Qje+MI5qmd9U+7vKEsuSHhoPJi99b81uXleSLC
dOkSZFCVFypYFaoDgAk5JsqJBbmtw1SHsKj1X3nUXuvQ3EY8siDrymU+TjUtP6p/
MnOfjCLyaDaJPbmwKdsnPABr06QbHjB7wVi8IH1WMpBVM/fW0bud8fWNOdOyjSby
RPTYZVgF092TCYEiHVzhZJCz8jcZG5mQS8aBiQvTOew/NBQcqGu71i5+CaJoqMbI
em+LescuXkNdVg0Gq4wMTlTj7cynB0g2uxFSQkJClo9HXE0EfRTRhA2tvt02Q2KL
rFJR2eTGWABTTccV6ykuhuJagpDMVfdHPYdIzvSTqZmLbs7xwvOzuXru2g5mMj7n
8lvvvMxPc4b2XWU7Ns4PUo7Og+dYebBVs9U/OpuqQVrDYY6cZx78QEpCguyV3rj9
hFcZUu37dUUtD1tDeIMuUM08obhqfyWvFOzdcZAluH1TwyQbFO2+jqztSTj5Cwna
iMx5fBzl02ecQK7DGM05ZyRX9BsuSzwNP66uW/9dWA80E01o/qyInAaeWcAd9/0z
SLtsUPPSOtD5jRvqGCWar8nonjQDI6/Wx4SXfqtRxfftQQQ40w7c6TTby9FAyY+4
0czj3/OsUhB7MPFgRxUNVz53AEOsAwy5nqkDCajZ3Z/8bPK0iEzVEF2iEK20yD7L
xnGp44Vnzlx1hFYQW1zoO+3JpK0Vt4h86WvtPrK7f45SZPouy4ROcszUG2hKn9jY
LEfIulFH8fFyCdUZ4cnBoECyuyfvdPiSt6BcusOTLuyzcYlPDfaEsrAuDH0Z4Z7o
VRK8vkNQNv/A/fXQyUtvuFvaZEz8N0SlPNRkvbpKRF6YeSMopPvUtmR0xFSIxgVH
ak1x6vTS7Hwt/9HSKT2kg5eLbPz6tISa1TBsc9aG4J21APkblWKlq2rs9NfcpqsQ
qAxVp3nIYSLOay+JX/YaB7tsdUGEXbSSM/1TBv3mrjufFWw4PKjYgJXG2mI0i38L
5iMEyiZzoAcRLlGsPIMVKxdAL5vXaKM7Liv1Thc/b37PkMoDty6KMrr0rSHzjyLG
vGBmOqyqsQ2eXemBm8Wu9P6uTNYFdMAjSxNBEaWi4MI5MLBjDoQ3t1ra97GYqA2A
fjEs6rmnzhUkkKAeIcev/GKWYiuShi1+qLpEBWBLCspY2nYDpGPSKFJt7P/sD/WR
vNwJ2JwPKBwUnmWUS8okoDg0fcW/AQctUDrFJ1bz0m26cnAuh/X98ABLuIo5agB0
SkdGqgP/vyfjX50oULKx5F6V2BlGhFEStV3adBTBf5yaHJnEv9qiQ13525DQ0tyH
EXjWgqJ4biDzeI/S4A0kWT2605qoPCdnD6f+F9xm3UEDDAgJJRXlHDyioqmBSzvr
B/j5633Sk0dDfoll3tx6yZj5MCQrKvvxFUUTwrJ0PZsYCRIIDQjvwLK/0/B27W6W
ZMFyMIOFEusWUHFRpadQHiMYaUJUx76Z5r46ExtTnvOd5BvrmUe9yXnGSzyYAQ6g
PENaO3v2mQdy2r1pIIKyXrXhi9Fu49t67/4Vab3eUq4TkffB5jCJG+2KU0wKqMIC
VKwZYegfLBOqqDLtRqNv9BpHVIwJwc2Qnb3WozPIyffHvpPHLU5gqPJWvNY/XJnH
O3VLT3Pu2xtLYJ1QzyrdB2wqi3wuR8ctaVHSM6lMJotfcce7Og7H2tU3tRhtJ6I8
bwN/0r9FHVz6svBvq8xL5e6F/dYe5eH4YuSli2qkRj1OTlBEwgtMcdY8semwM43s
n9FAUsxcCQBwsfY9qY1NiYzhXZGDpz7GKFu43st2jd0LcmY8d02h2uz7UO9FTx8q
/nA9L0iWJ5ZCtEO/AO1ZMCWNXuZJISk7vxConWMUjlYWpcYo1BBrHD9NIHKCKOBO
XxoooiMaaudXOFs94gq77ovcya+8SbCv4uq3mK+BfuBSdI+KNr1Ze8Z5z5L7JPZU
S95tvsEhRKRe0tEG2sKpDw/oG6gt90HV2ckVSdHq0HMT/V6X81FRT3uMncGLEare
/1LQsECfvlbPNUyAiV9FeX6uc+BC+rO1wB17ePABCEPuaznwZ7VMMYsOccqfjF42
V4Kwm999yRJ2oViOzA95iihQkiN4ldHmMAeXKSHinuyfXTlQHKbpcvzs4bqEb0St
PmusBUz57iROLfO6PgJWMob14oWHhJ+k10eKh2h74yNgxAvLidYzVyl/DXFvC40i
ypEE2CAEjBBhIZwdJ/xuBhucbp5gp/qbD9CiONY2xoal32ubcdX1S0iEKQ0UaGqN
4hLOvi2GhOeYwJsAkikTTIcdq9pkAY/FWXJ3i2MrYggtCs4qukfpQ+33lU/dhzco
BfT+3D2K23omKR0k+tG0beRbcrymCfkHfhKHuKKh2GxJixGunQgDWaReQPnhMFRm
6dtqszQgDt5h81fij2s4rCYvxhrYa0fK4ayZfxE7PO1bALjU69XlRdsjX92/G/t8
INieRPeVWaR88NhdZ5ukH3rwwqM7LTTftn7UJmY6TQR4M9W4tgARED5v9aQ0cAti
yylFS5BdgAG2fTN2PyH/V+s7ZIA6tjG80bqghfQq55kCRtOq4YzvLP/jzMSWlA/a
uv7rtSJLAe1SLzWy+g2pEZIzKOM0NsMxC6j/VgjkIRx6zfSx9yrvAlxkiDebYHxx
9NO0wLgjS1GFsR4V3FiWXfxWYz+Zvfe5Nz1PwSbATzM5phLIup1hu5+2EyMETt8J
H15nZhJRM5Wma9SjrYBcq5/R4c1qoQQPZfkstzEG/+CKlt310ZB3EM6QTOy8bqje
QAaQvd/onR6C4hzmat/RbxUGd7zTSMWXmS1B1GW9+zf4a1VSI/RCBGNwkvO4FGhv
j+nQQ1i6/JfZ0MmOLlRFILricpGrnMZDSSk3v14rgW69jG+U28pfZ5rViZ4/QYQu
l4bUV8VpGdaykdFDsN52T3Zsff2y9zYbAp0mR/afwi1OKlt2gs/qO9v3i0YNHksL
zvY8upAcM/ULMlQkPzdxxRAwCvh78b8I7xl7DwMLoGZFGZolqjERkEGhyYCIUc+v
puHg4Z84q+f9Vf9QD+Aw4ff8EEpFlCexAUzvgaaS1Sh6a6idZehohxD7qraeGu70
X6W9l/o8dbbu1xAcHZ/bdnPVj3paWxN19SbBg3rkvDM6bT5AdWOBCj9W8iRXSMWC
axkAI7GDPZmitRvaThu27O3103Eg0GEqdaXgj8bok9HEMMhlfU1dqrED83NEHWYU
sr93XtOiTXUhEInA/Qa9bPhS5BRQJ+e1GSMQlaV7rs6Cy2X0EiT3pk4E923IZN8O
Hxjan0cXasQILXbv7CWwXIJ5LtS6O1yFrSPyWsAnHA21cUQrIuD/XlliGNDuz8oJ
AXWYhuYWo5DJ1lH/mXGtxnvDy3muwKj5GE2+6yztERxG4a2IEOPi7X0mm1g2kc0F
HbO58un/GOIqM8BZbtPJR0vO1ch6SWboITT9CUArbmPFrYrwpIYUYYEyk2MqK9wu
p2+JPWx7QEpjJ1tTSAT8420+Yg96n9UExNFkxJLhP6LbWfqyFPlwwU0vFSN4SpPf
l0PFW1iKDvPXAVpwJOi10etMGw42I7rsjN9VB2TXfKuKvgMx8dMjos/5gwET7Deg
ytffudiZsnUn3TiH3A4f3iPwBnz8dZ8GhzE9zGk++CiAaGq3s377cMuuTT5JSCxS
LOabS1CBF7nqcr6qj9quLDU6o2LDl87/5FUXuh0ppqRAUL7wQGAXcZVKDqQMGXEo
jlxdW5LbjbLk0PrCJvUaMwAryu96+9QVmo6noIC5fkPIFtpuNO072gBHu8CXmYN6
GCWEz5iqrFrrTtbf6q4x22ObCae0rO2nLe4gKaqgM6kDQu8XQmegMVQaE3CIF0oz
RwngaD08eNCwSWq8yc8Hlnb1tQd24mypMIpdh0zVGCitS+h6hO7XVREyOm/lg1ol
M062FwE1hTvzNV7Rkmqr7GUAJydilP06rzTzOu40Plj7m/xfeyOGZvl16VUa88W3
XU70AjV+fhk+XswvW6RvsSwWSmf55rklnErARGW4kodSuaAj/CdV/IHGMonlHQb+
LCm/AaOse2RJYxlTy+QbVf8iQtOEgtgacn3tFju9YM45ZGuMd766FzDX5xPa/Qrk
S/eOqbCSKReX/fSF3an2XkSIn0tMtU/m/FAl+Sy7cTe50dfndfXlUCwF1c9/kGEZ
n0+CYkHw4X8e/hp6tCRmtS9La+U/F04ZLNXUhObty+U8Y5DFi9xg7VOgGRlENqNQ
suqLACc4ePxIQARnUZvQnd6oyKQmlRm0PYHpuPdWo5Gx9ylUB/rsL7LsiehJNO+h
f6Rl1GKeQ8uHQv53Nhgca+5VDijWPxGIRRyj6Jtk5KrUQr3iKRXOQMzzZDFjiU0L
1Avs9xOYRIO/TMsSt05g2wbjNj0s8ur4VXKDfbC+JIXfR6v473yCmMAcxXdolFK8
h9LP3PbzAW1cRl32nnHHhO/P8O7yNl8qQM7WcY2d2WEjgRHIrWEVJSQrnr/tVjRb
TN5Lq5WwWJwZBcHUPeiodpCp/SagqPQq8hJu/liPL3r9ssPdaGsQ9PwImq+Z0hPD
ciO0zZ/ioi7YdK8kYtAlLRKMxKonvRAayVRz4M8WjoHt5bDtYvbxfIpyzZIIPdtb
JBdb08ECet0YM/wpz+KoyJhufeJzL/U3jfmYToowUI390ZljO7Is6n22f/U4RULj
Z5HVvRWx/qA0mCKWUFXwmb6ytaGCd2rehvvME67vkCSUzxLI6brj4C1CUPmdCoST
vztQ86P9rLThfradoIBAfYOCKgH4UmDykXAqdjPG1WgnwDLUTTHs/yqz2Ug1MogX
46pnVTHOA5ruCHemg8v3ua/DOavOCoPd6MyiFqcuBK1l5CNMznxZiI0Ntpyn+VIo
IGFhvCtDr7wm8ND4gOuXv9234qsBcfWCH47SQn2IeinSOGEuToGu9asf1mZVT4Fs
OXscs06XIxLcDkSFzMXQo5+9rCHlaO/xWcY5vgYFdhOxolJCzcftGAtrr9//Dj1I
Mx74FJEb0LfcG8k53mZ5wJKeWUZe076acUL7rmqAB4Q24PCh4DsX0qkjZPB0hPpX
u9LsV3Jy7PQII6n15lPaUYLhTlBbtTIN3zJSHL8jKnT86xGFpaFgKjMIZ17UdPfT
971I8GeeqZLBtLKSKmbn9T152mT4UHGcv7pHCks19tedAtWmiVfpCkDbp3/38ztQ
R2BBGQV+wjMIfc5APuCz4E6AqTwPauDClJJ+P/+mmKtum78TaWBGro93kCRHwcpV
JInFDhsIpkOrld8jkhlBjrdmEDLthQEL2J09j5brE6Ex6O57c+RGw7/uV7rvxD65
N3g2L+htIWX1+0U1b1dL32/aFmMbgpLoReYCkrT+7oZUYmVzBXFE1VV2c433Dcmy
ibjIPe9Vg8ZJhOerVjQlBlIxll9a2hHvUTObNYd+YCXWaZ+dDGjoYV1HsrhBljl8
R7N2VdjHljrpcxBpJCXw+tbJCfdm4IbJlVne3guNNQ3Ri4veU0VXjU/c0DzCskwx
LlR5hljzhZFVWuOhuFJnl6TMrCcu56qnt897K5pXJDzZPpHv3JoZ3Iw4aXAIg2B6
qD7FHIjIvQ4LMW16AGkuIqv/MedITEUlr6WkQ/F0plB2XuFuLcZTzB7kXAFvhgU7
Q0KGLhkS+CG7b73APGyrzFBYG5Q/OBJiMBPsqWWCrOdqsknOflY6E8x+d9ceZzrF
zhHmB+F9AvyodFdYWDOGhxgVkTV0MZ8FweXIKlYgzckG7xWfVa9UFWGDvFRc0Ywt
IFhSnIdayXRzRdrIJ9ijqcwigVZzgsAq5BYM5P/ol/Nx/zQtP+CzJWvIIB2/1/oP
dmFOGGpIXvFY6MW6WEVuwMqNHy6jPrXb15IbZcsgY0o78/A53CJqftdTqSO5eUtn
iE+19D5YIdMvsaQLSKR6iaVz05lG1AuG4GvAF8sHAb1bxkMQJWz44TpkrIFGQKCO
IcP8vcHrcMPvRdZiFhF+T5QXnj338qZjoPz476WFqYfZQdMZls8S5dNZjTXpSovi
JSM85nTPpAqA0SB2Upg4gIbVFptjEYkNOm/0xT1K48jvbq2+TIGz4AT7xr/2JC83
mpWKhAz3kn/Eqe/Av1frxRFMM5EEP6aR9s/mK0y4DmGvv3DPBt6PWv4RmkIjR8/X
DYWe7601kURDp10TsdqhAN/126MyqXuLbNAiqa2wnUfTsxc1wk8X8I8/Q/BS8sLI
ba80ycc/LZWVse00UqAZBScQW2n8SDQdSJFzxLSWqb1K+JvAaEW3hMlLS9H2bolL
gGN98IytIO3WyDmHHi6R8MIxDHCrkUYu9Ply6twFNauji8vVIzbhMV+vlNg+jagY
gO0pAXVa9YN2Iui1Gsnx9JDFqbrUNpVLNQpTpxh42NIIkDJSzl1st6y+FX8ipAjr
E7mgwR5eHakVUnyu8EvzFr201fVvE0SZ2DeGAr8CESsrekY6RtNZo3oXOTnYWB08
sR7hSFwtOF37v+aueP0aalem39QWKdjnvi/40hB7f4O8ejvc+9uk1mXN6deJUSf7
xOdYF6JdIOXDvlrQT/3wSrrzWGs9XDBkuOkWd0mlwP7N14S74gfFilzTOoCDgWkJ
w95qyVg/DWe1C+OgcAkPBxxYsYr2X2Kgd0+S+2B0rp5tbeJGXMXDqK5mXA4GiQS4
WMoZU08V2Lf2vmEH+jCOouuVIc5DInGDSnr7cy1XMR3yPkfQbkTwHZV0+eNNpox3
FZtcBGdIVyobU4n6T11J6PjiNdr7F66ir6TzdI3mXxR6akeWn/S9+htE7AByhHzt
wz16CIayBhxrt9GGdEnF6aY6GApFZlNIYmayBhhbHacOYY7+Fua6KgIwICrtUgRW
08qGdp/emeWtQM3vVQpVVjW5dzKN0tQsfxdRA2D2tS3KS6kO0LISRQL3COTa018/
3iboF3fqDX0JE/DOiPcYSJ2E9O4PLUkTx4DmEDYSWoRqUxgH8OBiia6rfWcS0DpO
IOXzEnNZy+kjsJ+uROKyW4W12yNHj5/Ad/+ESCMfEWfR3qMqBTPqU/5qfqZ50nHJ
rWUduEnKOFzPjcaugsxDeRmjwcM8L8ZfSSNxFruSePnJU6O5Ypb3k75ADFdGv0Fp
jE0+/UpVJTO1ZIMgmOIf6+v9lj0r6FlwH2M5XsOj3IO2tJy4wLoHOLBUtwOjrJV0
J4N+anbRv051W9zk7d7AuHqxGM3t2akKIMgD5K1Cv1x4f7amBcOzZiG8xZPeGkwH
EoxXE30t3QuVCdjlbU/Xi34fx8VrCSE5+MYn3WnUM4fr7yZNtE0C+b5z09545dLD
1lzMw1VRVTyYMHdgKtNEKjh7GkYUe/g+SbumTc4rSpyj84QGbbk5b68MiUfYHQWs
srUbS4rn/d3Y+KCQ/mPj05C89J3to/qbFSPeU5aJkwsx4B367FE6TKrGe0A8Q0dE
KYlJ1rodeGnAn/1aMlNKlUn7xzq0VCyN+uOmrdY2f8Wq7BVV4xP9xC+Jfz+06TbI
wIiR5zuOU1/Bhx6wgVRTLfdqI+REUiAAZ1E7yNL3KIKBg33Wx7XIOoEN4q9fan1x
y3GJAkrKptyOHeAaLS9zhbYDeyhPcObC4JRw6nV0BTPFpd/5X2LLY8NIFZ4k5djG
vRs9XwbVuzh5awEe3pvzlu3rj2C/wJ8hG1wZTJCjbO2Ueo0fLVahJhZBjiYJfF6A
JhW5GQjkmKqDj1NVakcIZKHeqL4t012PUAv/kpHXrdE2jCPCX6fBGtDEWyxOSC7Y
98ENAQpilrtg1Hkv4sikg2SZDU49g4VQxdPZJfM8RyAafTxdO73D/opzgeMTaCRV
WCJ3SWfmDzdfM3whpONbxby/Ns3cwIrJLCOioMjiVzWh625Ev6e0ezCGBY5Tyc08
rvbXmb7i+by4E9I4qunoGU2LDEcdYlPXLq98y01exuw4q2ym3BAAjd2lmWloPd2n
eXOVw7Q25bN+7vw3wb+LJWBU0lx58HYNQ09GtVUDgQgENFdAIhEdJg4GNf5mR/Af
40t1ETgAqE+j/qgtrCLEaTOvKAhaoAI4tRpw82rG2fQxdGmPqLGO0Y8JC0rG7Iqj
eN3Z8qfx3YM8fJwFTzIzNcIj9rE3ApBowDh63oeSimS/wQSHtj9siXSqzRFSdoOv
tKDCA1b8LuASB/V+8jXXfzKBKUF/FAZ5WEwx8mSTZflS+exMLHCMkt8QOGuW/dUf
ZzypQTGx569voXcwuJEXJbT8rpYSXizA1kG+ZBr8Z8izw07n4e2SnCqO+u4alFJS
v9sVksXA/udWgHFI6dSQQVwQtZacAQUfTKLPV8XMKRkNnxqQ915aoX9wfmxRCW08
bLNpzqe21BfF47uWqMv+c16yJ3iotyB/LSG8ovBZQ4owbg8k2ly9yRaHiw5WjnmQ
a3CLx25QOunSzv37LEop/tR2uHChWYne2bQ5l3IPWX/gMm627WdQz93BJsiiVg1Y
3rftN+NKn0F4FWL8RS6IPdDEpUtxs+kwXmETqLu877PFOs2Oc8iSJMwAhbl5ZZC6
xmEbT1jkafQVzObjsDS2pdgJPS5PjIg+/9Dqc0WSg2b2cFQNCYQy4OGRlSHqcyY/
3FdSt5UNhRN5X3hiMaUjFNkb+5ReAgCZ4fv1Q0enj5VOhoeYmTC1lJSnDlHBry9I
WQFWzGGmJkAjCriMxCKV4qiznAFpe2bM7gw0dezlEr4N9Smom8JmIwaBS/Y/B9nB
y7TsipyS6Dv7inVt0MvbCM/twmoBNF1PhzWq9LqmurkOliJ+2pPH4U50VIGY0js1
cUKstNBvaHVMxBxcM6ZQJyLpTMvCNpU8WWJxDHWvUJD9xp+jUkSyk9LT75tJGiQ7
5rVW61Ja7OIAZShj6t0YY7uxKblhNSspN+0pKH80qTNcNY9ZRGzZgX26y7WYaTQp
Tr2lQ0scAJCLkjP5Ssh6dFiHxfVPoqXw8gCvkI/3tiBZbZivP3fV+7x5hR/xDADu
Sy88LMIBV/AD8wV7B3pg88Cti74tWrAfaCiAkYWpkyQ/lEgPk/VE8DgspXDm6EJn
Y1xzWV20e1xvqHJjtmBatGCtM9cN1dQV4w383gbnSMz8VDafSGtBOW4RcZX+87it
`protect END_PROTECTED
