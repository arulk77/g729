`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aW7lxg4Ftda2rP3oNVopicM5H28xZJZS1NDQfLo5X9DQ
x74ARr1y6aIVU/Uj9grOXa7CnB45RLCq2WUinX4H4SKLYCaRoCKX91kiw+anJ89w
M7zH0qJSa8OfzF3/OXjQsI8BRgmElMhbhRfmbNPi2HlAX7GLyfG7wz7g7OWOaEqi
U4Tk6zaByw1GarGwIrO38wa5HKohpq21vhTjpWnqW866MqGuuqIVJsMATU5PY33K
LFkY6/ziFXAinQpUvBtfuZtbe664QfbCfmxbwOPK+Rvgi4/zulefZx8GqQUq+WVb
qaVqq4AOxBKgYzCQ7FVdrVY6/7tpmDKmBxVkyUTeoE3mFhvjLjd8i5zjtMOS9v5D
6SKMtCYBPAF33sOO6+PCYgi2ApjRqdzAShSPGgaNrIukJg8fVl7f+hb5apmAHms8
qT+oTVllxvkihTMwoU/OInvnLn9e7va2vt/gF2tvNDhOlghhyu1x0bIn2qzcD4cl
`protect END_PROTECTED
