`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLiIqpuaOHxy+xRmCXWfOReYUmT7rURZmqRPvYSYTc1R
0svBJJ8iDE/yaTyW3bpJJX852uUX7mgui3fIJTg675b0uu3G8rliHRDE4rLOFVeH
XhK7f7eHQ2yKJ/3Cs1W95qcDKq+yR3XAmCmVMVtsslnYLK+aAH9/jHmPSHxNQy0b
a2Vlu2d3CBK20ukqcDDDfo5+O42+XbkDaoi0cGCnKRI2a4YUr1FLQcjTXlIuQfc5
`protect END_PROTECTED
