`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBhRIdAuUM+BkKleexCrLTinH0aWB4+kuxMG2/FySIh5
7xpKs7gWhseRCAABYRwK2PtadOAdK9tCjwpUGJwxWvARnDTeQufJScyM1xxalJWU
BA3igCzw9byt46w36mfoa89knsMae9WcIVxX1vL75UIkXBp4EcSQg5UZ1amXeQYx
iaE4M+xrL2kUtd92GubaIkaFv8AIX8W8SzqB2x2zOR9z3fgqiWKGcLu4lSPdkeC4
4MhJhg7juu1AcWiKJZ080wjZqrp4Ytb+WxxJDSWLfMzPJDpDUUGyI6sgTDnzPgRC
ueMuwqqqvo/pYL6Fbd7/suGKgFSzkw1/mT4slYyezD5knaDymVQ8io/2VSNn1M26
5PYGtdPy8vycVtMNIgZavN0VYOMsGaSSjmmx6R/HQNbBiqJUYU10s9Nfy2BfzvO6
ndFBIMWx0ga1U8M6UEw2uTR65rc20xj93DQYGiAf87HfEcs3l1lcTpKF33y5FNNT
Q7tBbj0hXuw+pQwnCy+PPA3HsmM2TM5C/iaQiNdYTnoCVJO4E5bXBwWMDzXstn+u
pwuPnx/WsMNoUMUbliidcZmT6bjTJFyBB+F84fmElPHkpmVT1TcmLBoLS8rR86Zk
`protect END_PROTECTED
