`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
BVAwhIDZDJI2i2gYvKkxLi+LQpkbke5WD3T+pqSBShxo8FUFbv8LSVaUe2FIOpVx
mzSwqwvYai1Ld6uu4DNIfVRy6iK4XsU8FdAzUYYqRa4Fq8lyx9Q9+dbzq4Uw+R99
c9wI23IodUpGRITDJh2fCixjKQQKPe81hKN6Kl+v5UY51k5zOmBSqOx0ij9uA3xu
+WzgmUFD/0q+gYFpH2+cvEjfKSN3KLlrRr2RsutQ8MSUlY6czQg3nLIPtZ6H3QEq
rLafH899L5mY1Nl/JKAHybFgbiDKFhrZmhem/VNgn7UfJcMolnnYtqZFiTNUBMWn
8sCxknp0UKvWp8SK5IbxaNfXr/qJLOdlGY4zLwwFY1VB9cN7Ci+0+maMDSt4cH4e
8Lrr5KmJGSUQFWvm2FZTJvDoB/q4AcYZALKG4oaOnbV9VaaGfldMWDd5YZ/Iq4KD
nCwe1MvdAK4iecVTQI4ZaS2PLb2KFwkyZxlpC8dy4KW3c59q9G426aV+tZxqP+q7
yq2Cnjpe5qJ1j8tbFef35enBXaUjCdFf/i0NrdQ3mibv+JT1jOhJO9efcU2xvDL+
OI9t/5ykUHuLqy7n/YlIqgMm9wigYGuDQ96U+rOYKOEJZopQntG88sLmvcw0f1yo
f6B4cNYxdTz8GGK42ah/h3udM+bE89Lll7cmnn0mucAR2tGjMdgVSzizHitVGOxf
EH3i+42QCvcFauN2eyPp0TXUJDqPy9YAtJ/g6l1bK+81tRQqmtZgbREcndjvl3Gn
SU3HnFncYcvaJZqnrnm6r/kVcFtM1lu/84A9ikeDtEPy5Pqi0ko9SEU3pngDM6aD
bC391gfNDz3T9uxjZZ4P9Ppb0jRhEjUnWbkUmogJ72NXyfIUGU0aITZEee2l7CBX
uBQLVfD6RfaEm+Mq1Q46Nyx2BkN9/p6g+hSZD+02GhlYaeyjXNOtilEXnPFp7DMj
SaR3wgz6vQHUIk3e0on4kKOnJIyrjRfO0WNZo+0BwhERS+/pi5DxvHGUGI2EBkar
PoOfl8bk5OLLw2E4aMz48cwrjb30qbv+tx8YQSY77WuJnaFU7KOvYqJR8jGgLSDe
Ls2SuSIum4gVF8Z7r18KhOi0GoNFgQ2AK080slC4NpoLA/a30gFbvHHo22qRubt0
lyNZBoY6Fz3J/Tq11X1EISyDS+0LJyUNFZzcC7B+vr2b+mQFmwDcFGVf5W2HQz4E
2c5h71nnPYszaAsUAkFwi1MxC01URupIQpvxn0R1uogOFBjbqlG4M7XYrk8l+Gtx
H5PP0JsbkKUCq/rNcYssydfVycR7Cg2tYnDQ6xowKYLq4kaqT/zl9aZGEiXe6QwV
bece2z3x0j4+x+QKLhh5MpeuQGQXT8m2tAnK2OclusUX48eROaaZ8TaGxacWQbqC
FADYGTE1knkZGsAEjyqQPrYLOgOv+QBc1d6r4K7hioBl6DMThJL5u3TTRuh9sCPs
uJUvI+hv3S63b9ICqniNFO4j3pz3ypEGLeimOSpkLtUlh42zodoFuoy58I8EYb2c
XSqpZSVH4KNdbUkbsTkQe2kUv8MzPg5bJdLEdHlO/TGm1Txkq2axAg5+OJevY9IS
jJTE6NE007pTOIQ7xNEKy2vHXTGvXeV3Cm7Oh4LIyeRDiQeidEqJ7ZPQHhbQYrX7
8DJBF7GxkRQodJaS461lM++8ye4nN9//kG6G7wDZWoKsWax86freG1xfx3HbVZxN
Aejn5w9tXMRWATI19zZfUcd5Y+ltE2ie+YfzrmDvCJYkEjCeuDI4IRqQVRWZWe1L
E5H4wnsc6PhzvOVHmWQq81ogHRoZoW2S2jtD1VCvEg+g+W4jo8WH4CA2NhemnC3Q
lukleabDPzEX473iX9gMSaL6gYuxsJC5EZVtcB5mLDYAtNavu5kUSnYuonxLUCVT
KoUnm2jHf+KxS8s9djjI5vTx8NJ71VAhRAy9zv8QsgujAFuAPnrMGCRwoQ7xTyZz
eoPExerDl9hfP8wL9ei+hPG6iHvOJ+XyhuVipZen1lpCBjfw6Y3mRb5ZkROgJ8Ie
LRl5/8S9lPatGAXQy0mw2G/o1gpO2t9K6M8Edth775V+a1RZXFza41799bcZLIK9
vuaAA1G0DYL3FdYqF0APyVyFYRLErNjZ1raE25YPkhjG2xGOBf7vwwFlR2iZ1U25
YZRHhpcKGlgFjA5neC0/IOJkPktdlPCxOO/YceEEfemyE8+RTY28gPFNzMC4jDWS
dybIUlK00Km6Iqtu89YgNPYzEQs/r9Mnez7Ni5n8FER+WqlygxYNCKr6A9y3oVWw
r4mQoO588WCp9GFsANwDPMbZ0VkkhCWvIduKbSV9n3/DqGSa0u4lUmP1XOTCGiWF
AliwINej/rRhQ+WxFkNduJ4QwPGvyVkyG489mIugW3TvJTy8tLMwZfGlIzNFl3Sc
HrZAyUSYkjg0z2e7/QRuh2hdgAeU7QRFoGI6mo3pI4HrTx5cdfTJJEGQTM/8FkU5
J6hMdzkwqjXs39QceughnICx+HA3rjU1cMvrJjSYbemTEK6/v/4y+UKlY689RG87
98A2FmK8w+AwdvzJGmLfOGx1GP3CRNAQaZcHWmykRzspJvaqXu+voAS2mv1WSpRI
sW4k1feuWocmYH2Xuw61g91rPzHw+2I6r1ZiULoNJEojEZ6g6DC11dvmVAX6hYLm
E1BLXzugsGp6Gk4X3RV+Tn5zRMRdLyvKBb3qTBFG8MV3jvfOcbkgCuFEMbFzdrv7
wBh3BJ3WY7xNaY6k9Dlnmiau/0XYn2GbruoRJKuPI42cJoWa+CLYcKg4qYDkrLoO
Xe503tgrr3SWWnDXahx4wY53awOf4Wh0f/twoyl8WdhDLyFDq9vf7hDVBJc/n+vU
xN6/m43/U/GBxUAZfIL9s017KHLS24XwrTrDAVfpqpvTjXAFAggkbnUgF1UbUxHX
jWTUZKyfDVZ1Lx1u6camnELGk+Dg3u7hWwuxyzNRMbvE50SILuZ2CLuOX7gkWSgG
gyF3aRxx5KXuJ8Sx5JDmVSauo/Ei3PY7FiP5J8XPgcQbzrhXZICcNpbM7KXz9/QQ
avIkzpgxfeof/YCv4toVFtKgpnbhsLh9TuB5M95Y7RX5fN+h/SXMOfyBkmvy9/RM
xmbxcyGKbrn9g0GpDqOWdsfck/5afwT7hrqoG0GV10sg3efFSZmCdt1vujAi5/+9
+4Wo0pLPm/ITk/8Adt8m3G1DV33fs6mFXhT4yaA0YiYu0/b3WTWf0vdNApHK4jtP
sTglmTE5V/546MZ4guWjouXD4+klrErWSyzSdC5TMCD4BrFicfW2TNllnc5YERYV
xg8SRATOrG4Ro3uZU0fWTAdrLUV3jFFol4gWkOw8b0ET0G8xI/UcuAYdCVX6eGz+
x7wsowdCm5B1Etc0Dpm87+DeK9IJdeWMqD8o0vGzETWazp3YLtkNNbnIWutcwlhs
NT/bTqJB10kDW1/5G3uxNXs8J8ri2FoLpmuu7J9lO050MgY0+lJSwpH5GsF3LMLb
LzxP4UqKZprqE6GdWEXidtyAiUqZjfmHA7vz9hNXjL53tJoiqqdAFPALDSVuwFRb
sgAB9kM3fnBjTQjMbaTdNWaaieMCUPEwuEMiGK+YozKu/SM8Xh1MRVRypsY7TT2A
6XXhDdhQQw1e5n2Uly6nFfLIdhesSwQIiDMdKIYSrvks4E3Z0+VBURqIp237wicl
xyGs2WDulZumP1MwfJpsJdzj0iq+EDhLeSPVDUQw04DOAGqlXcF4zQ4E5zj7zJjk
XoNYE1j0fsFB5CJ28qPzurzmBHDAebPOUQ+I5T5EcVNMr+wFNUqdcUGqhUdylmge
jVvLRexSR9PsEFsvysXyOe685EQxXc95f8wkc8VyVtyoYwM2tgpACcpwQ5o/QlCu
8H7mLSMVRy5Qa2n0bcygGTK8kmLfVfMAGJ+M/9vcL0eD403E/srw2GypNyzK+4td
h/zy2E4qKu+sN8IuQeYsRxfFqTnrik7Au1UxZhce8mssHULZ04zFjkf0AObis8GI
oavx/AhLKvj8ZqREMSuWdZoKghts6gB9umemUQqH6fSya4gvSziSKiaymdEtzEiF
8sv43vsQf86gK+QxgQwTOOKLvXHeqHbGsR8TP0shWTAyS+0ubqnxnsF5mCj9QFo8
5sq3jEXXHVkft114oQbtB1J2KYVMYkb70y/DyU4mxfv9s1PsEjeBcGrMF0oC0ztE
A+HBhcc6i0gff7C1GJX7aYUXitxhNPshpz7O68MJRh/hyU1d7e+OJdH3TxiPnJ5c
f73/Z+qjIQie5EjkFntPUhPIAYORZyDbzxj0Tj/bqXfG5S1Jop2yF8bS18GkTGOm
+UY5NlIajMLg14CXjLLXrEQ6g62sEH+A31btE5bpzOGYQgY1QZqhzgbrn8sm6Yzg
FECZhqdPQYRpBpvJqOJNeCzG5gzKPieekQSasn0eS6EN65KpgEDBgg85Yly6eDrz
WXIKedHHN0ryA7bXTyFgt1Qd5EY5e+OR/TDR5f/3xccvjoyPXhEWDjadQojtw4m3
tatPftVl6xvJnHMBb4WAXFjDclVN0RU2ydXpukLdYXz0wfbybWjHV4Ml+nxMfNYD
xV1Bo96+0VG+ZGgofhjYUMAvB/2+dIp6PJK1R7VrX1IirB5fBJgTOt+ny3oUKpka
xkILndO2+rhdMwgKhRs0+X20td+gKiYrMLq1KYmLKDTn2P2skqBUKIJPHfWsop38
LXjEcBdlt87wRFfkyg9qIO7MteRQ53z9es02QnqzEzUNM+wweg9/bEcbK3xFpWJm
sBk4tXq7vnCdtCt3Iz6tkCAqSrwEvgMtYC6hY+2uPvRBw1XNRwCT0kvwO7krc6SG
pBNV1UQnbBKMDQNGBbxmxqrJcxk6TrFp39VhqhNpUBA4BmDiRQV4VxM5CV0ki6IH
bnBm9GPM6BAedMaDQtZY9KJOkGLCGBLE8pkUk6UnZ3iHgBGKiLPn9U2nNmrga3aZ
rGUvEveFUSXZl4PgmmsJaFwvfqZym5ioMXLjvDFTHGTP1IYqXB5hEeyC48X9cNXl
98L9VWXo/7Q8VYfyK5rrU6T4AUmTVYD7nDPqQH+dIVoDLTvuBq7rf054ItV3lfPn
2e8bFFbx0L+vIBaqJUv6JTHdwLuhTc2s5SpZTnzYYXTpF5Aw3bs9HvjOOTIEr27O
s6AAUMTnB4GaKOGXgt4QjBDoN43vLv9N7Ixv+RzSLf55wBNcyJfn1Uba4V6pq7Ow
ycRwjdUYFk2MbEqZdaud/mFXQWBjstjb7GsuH2h0fIq+36CqG6KvH1nlTMBGmtZ9
GUheaV9KkkdDHmPRzRQCCVpM2bsR8Ww/u/E36XaB2pHBR7csftrO2f3NlRc5i4Zn
hGgdbgz9DgeB6Y8A9d3ZsvcbnG9SQUsEzLzq9XeZareXVZZVgMqi1F9OK6e52Ji4
VQv+3JTVpov4gNCDJC5PTHiLt1qLF3qj5i3jdStdqfVclwnv93+fwoJ1tLGKlVYQ
Bsu656eSrls0NL/W1cpOy6JskrJoMib29NGQ185TnqFhf8We3qJLjPdP+pk/Argo
lxGx1KZNHGg6O6URyo4NE+5YCPu8+wsyxZG8LrVktp+RhDE9s7/3WnuGaZFVqX0/
Xb2Hlft88pIoMYkT0zzlu40mssxBGKOLRcw2dPKyapRB+CoNLI6P8U5EOZZgrNXE
6KOGCXeq9yShEMStrizjV7OWJTjO1z7nkU82Qh1RNaYo27+MP4bB1e8Y4CFF++3i
FGKabPusAwmTMrzeMNa4wKH+O1n+SCjx6CiZIXb94GsxO9epWluuzZvv3fsgq3AH
n2ugukLlk8RF2F5b5DyUuHg3UW5r2hm35FIpP0cH1d97ngpjilNDscSp67ivQXCE
0alK2cX0TZFc9nn1gV50Nfcj+U0ZzsTu0ejBqhuN9XF67tCUHLsezgRxOoNwaOBw
26buPySXtT07uM6KKygr00UxgIdj5ZQbyki/jA2TZyro5K+gidQ5MrRkeO0C7qxR
E9YzbFfdn3egRuPdZowVubUUkNns4oJvMzp1MY/Y20ihQv1+Ia6s5Jj5WUXEDp/v
W/tEmMWWhSCDUB4Y7vXGO245kHWJ+RssbkLTC5TqXsHqwQvPpqtRAzUyP3mumkmR
lYy2Yw6LSr7Q00H7T16k7TbzTfo42UnLK8WupuAvhU44InG8h3hz2zrD/7fUblGc
U1+ao/n3M/ZYM/RCPKqEZptHYwoe3U4brEyP/PGkvROyVm1V/aicLD4V8E4rAOiy
AkuzYavmnhhOMDPdJVvE2G7P4ZCrbZGyWiH6rHVx4RRzNegBM13YaCegG8r7e9bu
grRfolQbE2ZIzyfsZUqhOKBagEiU9uYnJyTIJK+IGh//YBfhx2xouPy8q0drnOzi
gwW8daruIVi7ryjB9ROYLKhvHlWbn6MnM5P3BbJkW7R9VIzzJQWyNHvICHc3R+go
Z+QYoe15uO8Rj0yVzoZo9rrqyNHK14aJNgylD1sdkOLizZdfsVTlfRqCz+TRIFa2
hLJ2DcZuYwXCm/bHGEZqWrQXfGtE3/9U1u3MHMnG8gT9l8Sk1dEXip4ZO/pXHlqG
Q0uKAT6Ku7hYW++DQt6L1w5B9Z2RXSWJ+y5nRGBnw6a9eDIWQqMOyAhrbEaZRNq6
/Lo+NwK1Uq2fTiep2bi/+uvdLF1+xLofcbbgcvDm4IsfHzl2qQmViWwnBIslkZ2R
qRX2JTh7pJezQ9VeO2oIF6j95q9nCXQcveVx+7C5zqiELj2VxImTxL9nuNIE0ruu
YrXoB2WWDe1ZCtV1JkBakinuFsYcnz/RqGy8mhPEeuFdnqA6SMHPH2AcELCX262d
nmleVHBBt1DvIitXaMTjE+muT/5PeQbiAiH24srfnffB6Xtg8dp8MPndmxm/Gonm
w/BNaj8hLRiST0+rQdMACv5iQjACJVqKTHFi+o0+qAkVuJrHrkwsWLRA9+23gnKd
VE1rZeVe5MUVn/iXjlQPEGk1GL+XywyHn8xMkd3d8n/JsM8ShZ5aNlfKKoTOBp6n
JtggZmUii0c6J6Op132fnJCbfdWEeBgv8frBP5LT2FUxZdcvcJTcH4mMKyJs+Ump
w5IvbWlK6itpQWv8x2XcsYuZcJNF8ruZS1CFm/9uxlc6SU/jQCntxsKEbfzQNcM1
bvIpQQKcGTkoFn/uTjFxJX6UA3WK2/zyXoP3SNAaPwcYS1psNSY2hrt/aBUSOS0s
BOwPPNjPnRrcW9AGGK3CyBPS6IOyhKBukmNZ5497wNg5Q1TUscciMGd3/O0te1hE
+cz+rst100DWgyd/44WOUtPecghYohJgb6Pl2GVoTghu5quF/3dbOzwXWsZHcdkI
iT0Gncziqae3BFvsR1kXWRgkgjfH5tuX7pfFcpRm/IA3BYk0Euq31TEOY6/CbCVR
F9B2CqXn6cOD3zszEKcQ1eB2L7yhTI5jhjijytbyUip5KURsbG1CAedNEba2yZFf
id6DHdyvclp9wNRHjJciwOHVz5dQ+idOXW4yw6DDTD3P1Vwla6HM+tA4qKXuRtYR
TU4U8L7kh2+/fPATnFKYHcDNFd8WlHU0I8/iePAhAM4238JDRdqiPLa3coIfDwaQ
/tZhRd0ZP0MgiOUur6U2zNopN2KvxY8VN/vfBnp3f09ILPbEWLVIk/kA24LLMg7A
ykCE4XR/dXkVRM2s9/KtgxUIBOjYKnxMDf+XTQnBv41dtpFWOzP9oNiGw/L1rgyV
cftJR1jhoTU2IazG4YILdOT09LIpmEqRCUVZTdtWvfjkdeITWCLm3PbbVWzK7K4t
629Jhw8jowyAlbevXMIaAzgvOU+LoAnRWT2CYgYcLajc2wJKfapbtyFH/sb5KAoK
sEx3vAzLJ4kMeetrKFZ6gNx+2H6l1m35bt+4wKhE4lLeTm98e6FlEo/o6oGgVVcY
pTlOdjHXjUHHkmLMgpHQ7iI+xBBGErpuqaNQNnTIpOL1ggu0jPFHLH2sNtKyMyzi
gxXSikpG6OSoH0jjjROiOVQWAV7GBs3JWSwrhi6laf6ZyrFlOf/mZ5VEiuEFyVAX
JEOP57EI9isY3txbRT4+SwZpclvTfQD3rifslYhXi//fNvbfc0b4vm+ez4WdZgRK
nMkmiymTcCmlM2DWAPSCl1jAGoz/YgcHcz+ONdhf7q88Gc9Cr5Qbd+yGzsTNV2vc
BeBRXyx2YTbS2oxH7gKdQpHBx48Mvq+2JUx9mRXShsh3meBwAmvynxKpYUurAZ9i
MUZYDcFlUgoyD3mH92blW694KNlTD+DNLkG3915+GHJqXuMmsSk1cIaL0bUjZoxh
X820s8yLxrzjsz4coXJMrgMk5mf+6B2jVahSPS1GzmvtQnOtxrf1pXdGuAO6RpMz
0gELvSwk/zZSwDWPewsnZTt9J2k+1kXwft5tJ/QTflx6HKy/F6DHu5+u+2SBV7KK
R6pMXilyB9NdtKO0RRTBp96100l9nT4VHum7sca/Ycv7Ybr5kZ4AbVrcvDq+CF7T
VUQjCfm8f48IqQrcJC4HySaWTPQA8qOFpctiSdTfIe9CZE6lWKS8V7N0Ns3tSuoG
Ps2DaiDbsakRzqu2ncj2ZNmsaTIcY7Q5u4ph1RlAedB3GM9+5kzYpXj0HrRj2v/E
z/DRCrSYKaPdr/6tcWILb+C+Oj5wP/TNkyUI78FPUPmf6RHTlY8+/jnVQ8feWSgc
UOsQpgxr4c6bXGpktQM1FHvvJiohtAPKd0de1PSzcGQdo5tzln8TpSbXmuugG/C2
UE6Carzwyh/8Qvi2Wx/qud9uwGfxMdRSaBc8yPVjELLYPgHgasW2gOj+8C51zzHM
E0+CBt+w7Hmi1tBlMx6GkpncxgCCj/N9VdFm22mBH2W80HpqwXmqSgcWIvrCIwkj
wXFhW3SCbJjec8DJq7Rp04EfxIGDiWp93Q+loOifmHv3PpNJYHmNiHBMRmPvUIr5
XOScwrY/ilw4MYdbmoDq3tkENUFUsmd24vfUueUds18yTeB3tc4ghIv7nqJkzcQe
D6nQ3ko/ajwGBFCW+8irQJ6YntBWUS3JCQXdI10hk8VvcdcSuZPI4xd7Ho6/9gn4
NBc92I0V10gaY2Ksn6fKLlDtueq7d868A5ruftY9gauan9hE04zXQ61b0uYU4+aG
Rjh18W8jxxylar6svFQP9k+jDAV3yaY64th73IefjmHEMrx7xKQyea0Xif7zV45o
sihIPqeoYClfQwYwQxKtt8nUFDw3nbR+e15sF6uV/fCBchmSXKO3gJmtXhfFHatS
3C/dKxzXryK1uYmlpzZtdMcPmUfOjlCQuKFGmtoZfDflK/MVjgdGMlYN0hBGF0q3
Pqrde/OcGDfR7yfzEDfevI0TZrs31bxlI+8JLp5wMsuGpbyJuFM7+Si9npLfZDqZ
fwI0JY++BWWxFGrH0Yz7ZHZb9GLAZ3BnPWmPIlPXcrsFoS42//OK/IYAxblsc9j9
7KQadv5W+TwBNr+C+oPYa982iIm+ZYYfQaJuj2Mrr1DIklcMhbgsQWX38Xr9hG3E
W0yiZNGcF945cX2Zb6Gdu7H72Lfs73JZp5mzCOcAF4u+jGZkf6ah2BlFqsMxHlNF
yDm2Bhw3uIRxXq9HIZ8T8wBdy5huEaN5K5M2mNgV1nuak2MjFFwkOryPHkm6rv66
+1voXjue5/2xeIWulU3BKb3xzUQNGAy8chQx3M+Iwftqp5Ydqw3FZeVW2YJYDQMw
A+hdj1rPKkFkXP/9jBB96yh8nMKhf2e1XFN3rCNLM9LrtSSNG8bV318UgsZpuYmr
OEkBbw3NMGHBd/d+UBAc9LzOrp3BoJ/r4D7yxyEVDdVhMr//to5mhG77TtpvjrUs
HCH0NPI8NAPfOZIj9zWm47hDQ1H28MFsVrbnStAtCNeoxM4HvDGT+fRrQsEAgKh3
F7cpQiWR1Qt7FuK070i/n8151swBLlcl9cSckFd4HQcB0dERet7SDjZhxrlxdUab
ifO1aXiLW85MQkh3ezpmFg0+uYrV41o00PSeuYK0DS0ZeFwATwPwt1SrqGLFa3gK
aTty8eoVrojBwhnniWxJglH2I05Tw6XQGkBqMC6ae4QzvyzDj/LORN3trCBsCs+0
qzvxp+6uQJYMzzfp/LYbIkNSnLSLMivsZ886o8TD20o4ljR5UFciuoyXHMRCkANv
aIHew8UG7zrBNRwKXKT5Mxo/d3iDIUmh7HxacHuWG93Ua3LZ49PVphGZuvTZD8YQ
10I6PeNTyJ5WFHkUN04Wdatp1f+yq/DQ408AUWHWLOZJuwxClxSOMwxBuJb93XGn
YATpujJLVjYSS7j3HWyQbzi/x10RorxsBO3dAzoVgrqZ99mrmO1qxkcHI9YTBqZR
1eO4zBlKh6QxH3FEzArqXAYTUI3OJvydo/1u6kQ0ALWZB0aPv4bOIH7/jJiertFl
nEi6S+/VmhPdInQdeL1C4XIu/AmOqUIeSlrW/sYi2C0Bxiu9PDGowHQQKV4wMqss
8yZOv/ShLYMa6+jgmT/BiG63nd+AT6bTcSknWKqGU5sJZJ78vaQJ7uU+1SsJ6Y+t
TsGDD6dtKfvlm2LnoZk2UOy3MTI36Pxdw5d0Omq25KbS51PLaxFWjKSxcDUT2zQL
QS4xau++DvFCE7NT3Ad0UzuyR1SZUgLS88GPlhsCGuDnHCuwWYbJqBHaI7H4PrQD
lFJmg1irBTp6QwrPDSXXEsVAnwmPvz0z5zwVnK75FFaYS5L0OihXscX8Rv/ibwCZ
o3xuEusJTJg5pxxAEn1agilVWilsn8vjC0RYI6zIZl3zawFFnPaxrd8d/QBIQggV
6VwDzPVWx9Soq7oFzJ9tpgkqP+gyBk072s/aIzoLpUaZIcLdq0wUpzVUSjL01UjO
V97qQGSeO/ejkCOHmmvVsQ9wC+eFhwyaWBT+N9eVOUBqLJnpWOJfmW+tOHkf8C1D
mLdpDsR6CrVOFvPVHxnAqPS5CVvOI8aE4xPUlVPpJSzw7yX4F7bofjxkxCYbGYDj
UJu2fJpgwPXRuPcvu6hgxGLSOWM8b92yVQOF4pKLyVPq9ruwUMYhQmDzEDaoHQad
LHHk+aHEfLZlO6GdiyV5PrH2KUw91EpDUPBEZcrHy1JBVm6PsAFj2zKXdsJXTn2T
l29Ttwg3vtoDpVlb6CsJ6rJ1lOtiC3FoL1SFSsZaRchAMyicDEbgfjFPPJminBrw
R9WdnQZ2RJIgxCQOPSCTutr35cHyE77zpVk2c7AOwA2o8gVSOstl2J06Jh2RDZaA
Kv8Qq1JZpjazOV957h0xbzYi7s7Tev/HZfm8QxGadIvr8wt6Xfoz4PWZLjp+OzQM
2D+OH7Hf9/Dj0X9FGkqaUHbg8fh6DV39zAae3TQ9rzDc5xMZcB/gxvbNwmINrfIQ
YgEy/rJ9cQkxZYYbIg5tXD7NAIq0D2qb/pO8y2fgoLcMY1/5VPnDFWy9UUXhFj+k
od9RJ9l5Hpdb5bfA+FDkJaunXTjsOh3OtonEH9jNyFt+CWQo5QpauKGVNoC/MMN8
wnz6VxlD0zL7uZ5d+AcTsuN6KpRWsaiI9Iuv+OckUaV27pMth6izmVwgwtxNrJYw
3XoclkUZxJyYtJ5fDxoNsvCnz2vxHvq/AgO1ik1TpEXErbhdrsbGcbqz2yv0HT6f
PwijfE4VX8TAUbo8knpHjvFJTtlQcCF9/OIX/4NK/55shl5HM6pK1GWszimb2Rxe
sKGkooSKw9hGGGLQmwH0fmh2vbmTtSymq/A+6Ig1GGEai3QJ6EbRQR2lg4mBCmUk
iYGMt93NbIH6RXlRnmN3LEU4RG8Pi9xS+XigxeOY3QljsUfsy35g0Q2GPTRuEADA
R0uDPwQK/insYpDOaCR8ZM9T/pgW5if8hNxjZcRQufiMHdqWJCF/IBrpANV2wAwZ
S03Qzdqe4e4Vys1lBls2Y68ZbrElaGd1O+9+v0kHoUUE5JUTKITZc6dtnJruvxao
l9/hT54ne6EIrFxk7f7epOrJF8BzxqtroZqB8C1YqXtTGkVdAvwVSDVKwHDZckpI
TPHCd45yXFvtMgjskbcqE7elVVBH2Bkmd0aZi8nzBa64JcHl3/WT+I45WSi2MzKA
5xwQytmB4EdwgjUCF0thRg+Ns9SpQBdttr3SFcgM3FpZ52BXnh4HG6Sg7lgyGPMd
qWO3yHaPj2KrU+Bfk4zIsG5q4jzjVFK0CDZ6OmrLEauOpla4064LAYPx0dq5ROu7
RNahQmC7NeQKzceEly/6/+wWG6AYR/X/D0NTmZLUSbQASecf0CW+Xu2X5dHvLWDg
kQwu4DIoWdszIJHgjOuVmCQFdnpXguULJRZZ4yCDFdfXY6GyNUMc/XyRmhsRWLvI
gfoUoh7ObtAn+F57eirDG6+6j/k7VVzu/6hxQWaVSGBxLM6WU+opjKbsUmS5gdjN
DXqG+nZmMbKcUM6H6yPv/dr5t2LrRBZHuyPAPYwM0knYEV6FKABh8zqqa5Mc3r2G
CAZVUzjEMb7NyxXf21DSnSoB4nWDuFQ88gQh4i3Oy+tmm+fSfVANQeJLQAdZSeAs
Z2eIU+76hhz+O8f+ux3i7Irs2eqMGhzkGNDmuZiIMRAiRmeqtdmjdQeq/5cz3+Ny
nR4H+X+UnPQQ1Qe7EePVC8TrluOIWahG5bz6nk3IziGmvl+t4kqRftoTHEaMWCr/
qo7peTyM79Eg9zF8W8Zzy9xqZr79kpVdD1KmlFLojLNC4TSTQKNn28q1m2d+SZc+
mIbMugfYJsa0/jtfMCI4MeuyrRZ0JptkWl/BL6ikZmzpG55JiAc2lIOQmKlwjRgo
Ck00k5y0yJgqlh5fK4/o7NWzC99v12sQdwJCBPbKImUVv3ykozclWikJltL+h00M
+M7gcJW8Ak7Zo2sVxh9RyJL6AJ5sfgo91l8TtHVQJlp6LX4AUGsCs1IjIIEyS/JB
54fu/SA8YN/vVl8IAfPy9zHXOqRpfXiPGbiKEfzeIBxcM3TIibuPMy+joH3OS6wC
tqnzMUABdWU6jWz2jVQF13snA/0x1lAAJnd+nb/xiONWnZvf9PamcjtZ/Vs+ml29
MzkacvP/VgLCuZTVBSw6Doer78lek3lhxiV6vCqUNIo133Su6dOYYBTJ+J9yCkgy
Cs+8M/SI6IgyvzrMT1j3ypsj3LHTjKoWxbEq96tdQ90fEVPkHANyZFaah/sWphwY
s+l35oGujt86VSfgcvVYYA==
`protect END_PROTECTED
