`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEbjXp9PmY1NLsp6U2bdACCBpilKcZ1tPRN/nXG6QfOc
iCvQAMPGW6C5aXglVP8WmMt7HnYn6AhbRw+Ak/FMlErQWb7yMhFODXlyXncQuiq6
hegw4UqlTuXVXIamj6fUmye0554Im2hsofN3DJFU0C/xhjbfHvIMGTreu4cNSxZb
J16LRniaHs4yc4ylXRQ72tV0JW1ZlwF0qXYP9T5z0tUoDHxeJKsLOeffJuCmJclg
KGpMEN3vGXWNhjHrZLzASJ/2snd2IOMaS3DOq5U5awSvl/xPjJX9kbNhNFb9eEfp
Gvy/BhZSc7tJdpkP3RbnSTPqyQYyke465+YyqFQZAvt1RN9kIB2IjCar5qKdJpMb
`protect END_PROTECTED
