`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
lmay94B7QtBVEuUapwmGXYmPR6xaYt9gyK1qmIYPK+UADCSHjHuL9MzShJYMZhRH
I+vh4GK3p/QoEax5UyZwdgrLeNzXazLGAbVJWEqQoZTVsA/b0KgpBSBwll0mgCj4
XT/+cMN3T/zlKZf4SY+R6AIi42mpf4TLSJvutgszcXdmk3gCelMR35W6QiIRkZBC
18/VkJTextR3SzPi+qNI1tV/GKvSvGkfEJpYBEewefCcwDckxdzJBxuaWqWMdycn
g4vZR4QzGtLKhScBnYsqAVHThvKySlJUWB+wHF985J308Ahsk3Wz9NvmEPN3aAXQ
2R+C9OP5Qi8MDYgYShUjpeYYIPsBYHNH+xOEDvrcVH2zLI4bkM0lDFDj7292JhTl
f2gU1z/zN3oKW43aFF5C01N8JURoCsepLq2LSgeJwgJ9wIJQ6N1n8EnAIO5a/nb7
WJmDLm5oInou0efi9OAvnA==
`protect END_PROTECTED
