`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePig65q4CXw994g4eX4y1Gq7BFYsyZnSEvADYSJcFNco
z/dJmZXxODuIDIem/TdIbkfA9szFhXpzPhF3Obp6Ir12qys0ziwr8Qczi4i9z++J
y8TMIAdIrgBr3erwxXhkDVOz+QM8ykzWaXUtrSFdMb3DbUIPt1V/UWPJ9ZIDsmd0
hPTNUt4t1Ieyth5NI5oSxzSQJp2TaG99zPqjmZxeTbKj+l7n0nsAhnPubcI9WesK
uUzOmS8jgYiLgtfTnubzL0wVi+hOZGbAXOtiJL3U/x6sfps5t7JmWd2sNjOk1W9W
TSV8atfJgOyrhoI7YhPBtgDcWwPqhjzsjl+vZO+1/dCi9gXB1IociY3aMVNKwRQW
qWAwK5gXizSDz8s9Hj/J8fJY4VFLwoEMarGZEMDJTY0f2+SsMahHgGSsu+jeop8s
gUPGivTvgGJM6e3VQ9l1UdL0Zq+wIdO/qTTzGqSav8zonoYN9VrptRbOFcpvbNJp
`protect END_PROTECTED
