`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB7AwCIhqYwwSvBEmxA572XuxEGb4/s4XhMr1rrUjK2q
8q22YoqyPsOBp2HFH7CTVFU19yXOLWnmtdc8w7OTYNgBqTl/Jzzx/wz+/HPvGEaV
l2RcTNDoHTzn3LvO5+QA/Ci3D6tyZdWSV1MjrRi2vsa4woBvgD3lYHldbvxu5GBp
7fRvNr175rDBrblHZxStiA==
`protect END_PROTECTED
