`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKWdxQ5WfjrjM9Ex5/fC7ohYJo4mo7Gac8j5Qg5uB4H0
fuiu4Mws1fuYzh5eIgRuZtqLsi6+gmsJtBSXt8HOAfRcQaVfJyZ57Rwr/qcFJswE
f5tgPthbGA6URFnDKRi9psY/j0sqV3Z0ytCGKpOTTsDOYeWFKC0h9IreZnbM+Hhv
8qZJ1rnuqtANGMGetR2pT72/8ns+sQjG1QrsVpkHhm3pFl8S6u9bMFVHHzwpkNiR
gXYh2R0ZH2+seC0wzLAwxWffmSk/6N/ujWEpCWJ2iu++3O/vIxIJtmjXPGWR1XsC
+1NaUz9yRhNMGXS71hTlqw==
`protect END_PROTECTED
