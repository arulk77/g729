`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL9r3h2sUP3hickHYXbninyuPB+UN1Yp3CNJDNDvrdDZ
FM2/gGukZg6kUqrOIkBL63tYoYdWVijNXTN5aqcxQ03ugliMVvsvEiZosaVuhN7S
SlDa7iWskA8H8ldEYRWgwNEhpdMEqy5/+udkbl7Z90D2yEj3hDk4vh8t8KSHqTtS
a0ULZivgcybMqQva1SzNiyA9vuqkQvhtwwxyi1FpLmihmucplFHCONWdLUrf5G5c
ocrJZIpVZKm3JQpzoimXSw==
`protect END_PROTECTED
