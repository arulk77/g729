`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAeYQQn3m4BDWT39jhrxgz+60Wc7wGhuS8TFPyNx3WYG0
auKSaeIWxei/Ir9aRIPVKBJWUnoyL5xNeEDNPIXj0AuBYgx7VxFW8WMf6C/mv+AG
+WNlT6Z6NjVF3JB8ezncgaTDTBETxd22NvtwQWqMOVJ655GUBrL/igcuCHYLbmDe
zhwrQTJWbcuq8anxOQTDghmpF7r3TlA5xW8JEne7iVeNt7fChp98L/zgHEw1RQoq
oTYHxSYvpNGSufzr25/aAO4PGWigGxBWeP2jjes8oNJc6Q2JwqUBtgZBO8bzajAD
q/U7jU7Le2nYJhPCvF5YemIV68NDDvCg6xFBq96AFI6z4TfXKpkzD+gDTUw4p8Cb
J8JztB5lg2X2HMYCRLFEYTC79IQc0Ii6//n7az2CRgkmq4bxn2eGYZm1r7llTe4a
cCR15EJIsm1kp9rEgXbeDnyEQ4Cv4/IwxQwJBSpwQYLmimjlg0t3kTMgHcTTWIWJ
ATlYf61COngiET7p7idPdWG4yj2ZOjXJqaqU3UkRoQd71/77MD6lSFy2GnjR0fC0
B5OeacqeQz1Pab2e95AaBdFoCTnh2J3lzQNXj3RFwu2Cm3t/Oq+B7sdj3ztweluQ
7Dc5W+dl0qj+kQEGvYrWLjUGytmb2njVBEPDNJQy5swEj8Igb0T5z07mUtlafyHx
uT0pe9wFceX5JXLGNLTcKIwNEkwK8yZBxstHHQzVLSY8k4BhcZ3N2ailmdsvtUvw
L55PhZ54x0bIl1SHaV7AzQXSEnMtWdeME0pt9lHKk+hlI+5G8GCEbC/OIal2637e
Lz1g8PB8vUWdV0kH5syO59EMTVfyT+VY+VLm13MzKX6AEc/YJm72R+nE6EZCvzRw
fCcIiXIUgUCDf+m/2DJzLkfEbh/+K2eze9u/7DDQd8LG5tYmsO6nvZKVOhHcr/Zj
VI/JuPZUtggDqa4fehXauZVPtS/LpHb9OWclHe6VBHctZQIG9cIDN5iy0dLtcn/1
QZu0Jo850en/MDz0WvsnkviCDZm5dnFnMVNM72fb8EtJcn9yKckNtySedjJI+1Nn
2iYbQz92wVCu5s6o9DYOuPDq05yF/sCHo1ebf0yJzcj2UOQKz1m+nY5nAk1HyIxc
HHfHRg8SPvSLILW47KjL2mBOLSgBU1L5BMXRJt2SjSuRXXR58VPFv0z50aF6AWFh
Bcknka3QjmaXy3iqyaUWa7w/Re0Ck6zbHO/UxvseMoegrHFZQcp4AWX3alNdcsc5
EekWdfx9jCKAf6sugtWc2e6slbIHKxY60mi1pCgCoPZJlFH41E5XifABTiY3qkd6
yBfqkTd4kR8vBR9qOnOXdG+uCDC4TuJw7pGsAPvdlN3EYzfPKwIvjgkuOS6bCaO5
mP5cWCoQdfTQfk3q5TLM9XwnjL+c+iITh+H4adFKdiajIIsc1luGZBEI9wLY9+p0
xBeAI5PfZVPWDrJDfbYOV58/uYMslo7oogSPH/Xc18kssKP0RJkEzl72/35POJP7
8ZL2Kjb4G1h51XQ2pOW9ZB0Dw/cYgAZP5ZuAaCfDB8Sqgy/r9qKOCOsHCpLZySyC
K5FC0irusBn1js3ySntZwAYMS6hXZA3GsRV9BwuF/smThu0WomjLpEYZb+xAQQvZ
eDiX2oYp5L9Mykm6KdQE3OzdlK+a/h+p1edGAPBwN0JA2GdRRoj+e2ZRKHbz2KD/
sv5xv56q5yAFjMd5iDTMfYbtDXMYVtmd2NF1yRSl4HqGOoTvcU2Aq0FNQ7IbrO6C
Kehnvz9frMM5PtFWi6P35LsUoJG2Ox+Il87zTfV9XXe+Qv1dNa575lX+FGx+iMQe
IX8/U9pqrXLNe4SlTIYynI1el715pGLyIhd+MiBazMm4MGdpYIE4c/YD3DGcEBWv
YbzqS8jTMlEFe8MoOY2EnXVZhpDxozDviLs95TBak1CRO+qE0b4i2kxNtcWg/vZF
UyndWImmKz6U1FUGb9HDImpZf/d7yvNMmSceRWKaS9xJC56zZZ4lY69UxZX1j4QS
K5zyCRDEJdSWZK43/jKpZIyJ1ZXooxkVhfH45n4GqrNCVeSy0U1zpNi+7fzbDVOx
JMT88chgG1zCiDmYyFr7qoHbkT9p8aaltDt4LeLzkzS1AHvZAUcDohqz06WhgDT6
IVunDL+3pYngDFfjfemM8i+G0fPfy1DNaLyD5vvikz82BvnsVNYyVuVGxSqu3+kH
+gnCrUpq4qLPMWZnzFpQpbE4w0lIbrVfuB8Z59TNktT+o9E49wFzAle4qNn7lEl6
mM/UlStrW5EaaQ1zApv/hzcXVZ+4s3ldGzQRuOELtnIZwmLLa6vShOklN5r091rC
7kJyMJLgpyNdJKybKfhNOKLaU5pfhnAHXPQPs9eF3sBNbrbCX9Aingbxext2GL0x
S/5PbmvoZlpdFMf0cacI7SPWfXhlm2R1D9fB/AUtXdUJR4mVSuuRhVpfXWwK+bX3
26ds/oIy39r/0KjXtRgaRFGCN/bZA7CH4OJxIqjvArJFLefoVUNE2w+sVljwMpJB
+uiaRwWLtYqP+krYXibzj6ltce8/kv5mEimtYgho663q7RP22eg362fLSyFYA8C4
riE0mw/IEGaMvbdriLkKSDkVwXC8Qv3ZLBrIY8b/OiTVvEj3AJZEAozmRPY8lAQi
DGJssO3JmhHyQwk8vnNAwvPbnVNQDpmfAF6TpvgBzY7uPds/ojnNf0dCyHYjO5OZ
iPm3ADmZFK0IKYpau5kmtQaYYKZJCu0dcvPxwZfJI0tC1+JFV7tQfEOUFRKdrWXA
wtRmBG569Tb74rct2MN4UzD5OJ+BTvE8ytZm6ynIlp4aO6CFHXgT5DdYcJ9h1Djd
Tpk/B3V51Yes45zZ3FkZQ+k8lpDdec/sEpscMe0yXiT7/A3d97FPr4s+O9Px1xNM
r1BeSFRP0sriums8PFo9rurLA/HF7yY3kJx8qicKuGMk4C5lHLBEgb0+gfLGPDo1
FwiHV/v+lqPvcGnxGL6yrPjBallG18uRR3PBBzBdeHo73IO8enhg/Kh+UiFAS/Wx
9CyxN0yIr29VZ0HpWPWAclUsBmO5d21v3MfAUetoAyg+0ROnsPR5S+5/lZRg5WFZ
E6yzG9EGXJABBny2GyQKivcTJrPk2TDhn3q6qVzjgMx41pCsd9BWGDJqMHWAA7Rh
WQDdGCg6qmvBP67i4ffDRgoCqIyuWQXJ2yLkFnqOkSlow8QnCmXRAGsIuN5Vr0Qd
qXNTfl05C3ORDn5gVzlYuUSxEuJuYUrp4dnAakBnJkbe7NOo16NjhQSaoG8bCpY3
ahQqPPTTLDpAnOlV/I2MiuNpj7VJbmYoGoE23g6maI1bsws1ff2B3uHwNRj+HRMZ
Gdzs6UFkGqjwSmztrMmM1SEY8XeTzWr4+nz1feSZUCOKjQYCo4NlrmgwCQpXHXca
6FSCph80W1DSoHK9rXIz5Csvmkmd19Re2uTp2sbw6fuxxnmICIErxRoha3mr2Etp
803fznoIBf2cpiRz42CiEEa5vaCimJf9TzJcZvr8IaU3MYkfsWCnRo9yuBPd6fH/
Osw43XhNQJo9MM0YnnIjPe8nK+2KCe6I5JqVyLCIN/l/5J08uBUjQQoyhrT7knSl
SVhY57RhWX5vI9/q54wBQIfgDn8sjjZXC7kUmyeuhNTTkJGWiCnBUJGo+xsJ/xF6
C0Sxe5LlKjELJkdvlmO/GnEMqLoywaXUnENqmZVJbN3EyqMuPM/6YIUTxsi3m9Ps
lgFlAfZi2fzxK4DE49b0EAmI247mb2AZbqhgwOxlKHX97Cfqy8tfAUUeWyAad/SA
sr6bXmDa5MPmo/QI9jngFvj4thT7OF92tUrZ8L9GWfOo1Aokt3FDoepjBeabx00l
hlmhLGrkeFbE3kTkHFXZI8EAZVDaRqYr/igbheWzQvqDP/iDzEagEQZB1EWh6JGS
QFudIyosXOx70Sw+dM1OsmrivNxlo7f1OqEE57ndRQ9yj/3PDZK7qkbot1PEGm1F
088KIUdiNVWzU+J8q3RyLCvo7YB449kiMciz04Z9+zOU+ER4d+l3Uc6kkp7264IX
3CgpA8vS7t6/uzosXHXo5gG5CXScEOFSERgYq+G6fOfMLjw63KsZY30Q9jroRwNQ
eCmuUDhx/wD2Cj/rQCtPlT4GG4+da4G0RRRMk39ugFNsOUjk+ruY5GgVbIu/ztMq
4zO04fRW6w/kqEo6CnXikuqFrSoKfHX/tc51fgvnSgKY5vJ/pUbowllmkuCNATWb
/wTr0UrSqnDL+auaqge3mzRzhDYaz80muHlLQezZq0Oazcg4lnY12uPT9TKyh0wd
XEfEuVJU+qiCCPdXAUZBbiP5E44v3OgcHl5OBO79HXMdt+ddkpbkGJxby8rCmct+
5uB6Lr2GtXjFLd/ZhC1yYLzDUHr6npDnShaQea0a2QxTaDu4Foo+8bQxtO2QSEgy
Yx690c62Z2Olm4FVPWI0WSL2GrGCyab9nAdOkjKRDDnTDVjzx/hLCR6WfwFKbbyJ
aoI3YwfqkpcR4/wn/bZLucPVIbhw06BN0Ks4GNylTZPd3yvNtZwuyf1f8/GgVCvH
H3HnXNxRQhxY1fv6cKn4J41HAo0UaJloScAExYeKZIPdP35NPFfkKAfxtRw6dCS/
l3NErtv/20mr3YfuDzsl2MngU3vuAmTHVLYhKYxjuaHjWTgfaP1tWwXiFhs+H9Nu
PhlGaBAzFUu7Mrxt/9VV9GsN35YnOJjZjIsgkrtNEreLWqqjq0Yo4OuGRMKCr/Wm
CrXT4lHMQ7DjETMC41rPxadJEkZ7G5HIva82KjiISKM1PUyjk9h28HWMgNHfpWMV
GzD9QK2aQF+kF20XmANfA/3jG9hwMBAqUpX7kA5wDaokc0AerTv1uiX5U9KYpRba
lf7mINvS5oLkAsyI2wpKdAjN0vbFEJF08yppV7sXGQeWGeBW0mxUgIzt1/Dg/jEL
Z1sSKcXo50UvKXfvsssNs9MqrQUHoqimm7QFqEL0QmjMIcB04ldJitReAf6SbtEY
gZWIeXqXSMTEXeKIDzCM6VqYdAyr3O8eOy7E68ZSB25PrlQN5blQQLvAHDY3532m
eKXEy6qAr6/BskbszaQP7U89zn02mlIiD/rLFPkc8IkVivf5SgMdROmi2VY6i4jt
/sJHINn16Uuj7lncGvtCUB2iHB08cwuT4ACxfzmML8yvIlhLLyiCiMXjPKr8iBwR
/98WvjQsZRrqhxG7C9aQpzsGQgx9hzHiuAKIwJ0itTsc7c39OYL4Dqge0ebp2tqQ
4VWBgz9kqVHzDTIWK6Wr97ScEZhOxXqDAzLS1mghdgaPS3kZ5Voukb4d4qgsPuBi
NrLKZno07c8PwVbOOklH0ziB/GwQMVdrWC/eH39BNX+lvUydOcjqlqf8gEfO0Y50
nZfxo+x9XI2q8m+PWxWwoa22NsUOxjmndR6AZkX/HQwhmHU2wneLFJH9n3Qd/uAG
gRfolizmG7XhL4L9jKl0aqUDcjziQl8S0q06LBHiWLDCZO/chpeOIjHs2aw4irD8
SUEhEAl1EQwHGGsMhp5Gg8FRWCAmZEH0NWwSIv02K0kxqAOPOsswxyMzRFwxDmYN
PN+u5HCTDN2OimMaQHuBzQdqR/bfu226bdE8SJIqVY+zepfBWWJTUUrYmOSYWexG
r56LDlvW4yJvZhZIApf+5dSxqE1yYj5YmFW7llWkScEdL/eyKxWZgY0VaDPazZ45
ACmqUt6bEd0D3KdQ7CCYlxSUXwJKfVO0OQvPSwE1NpNIohmYjlwmeWbZVpeWlYez
kXAXA5Y9z8pxzzwGnyML98Cj3n6X1P8BgjOENDHWZq3cDZzVDpCT7eqOfnwcWTC0
zfVXuIq12sEY4V0Di8eeI6Oc9vmSe0UVlhbPwJ7owcN3efo9z4Xf23gROmCH8zY7
SRG/e9UukWQ7Zfmvjn8Lf4YGVAiof+PDO+m9oMSoC9RX32vrH17LqQhBrFKJnH4S
lxM0Ev+k4K+KkFPPFNxFXsanx3M9G6Rry6Lwyj8cS7I4I/Vv3dandzLbzT96sLOK
5xhUs8iD8JaN06kms0qo4IghQZ+fQ7NodOiL3L/nfCGBdv8bOkIhOsAhXhAy8o8z
U6ATw6yszA/UT7kyH/6gVHiPCCcIOz2VSLMo8iqneGQbKyV3M3IjbFHuZnpL94tg
/P44WPg8nnnZh6Z6WpfmjCMPdhvwmyrmT9+U+LbmsGsK4C6AvibsB8AevpFsHru3
r8VjarYB7IriO/A/3wujkUmnh06HeOVWa2o4AAi4F0NDruczuvm76vV/4mw84XOf
Jvy+086AYj/2b+jE0eHDqJuojzNbggnzgZsZ/pSD6jm3g19DxgTBfptrM9gZBaHp
t97Od92c336sjLxidGdEKkLBATCak1y3T+8zKx8OW+UKWjHxfK5rjheBVtF9kzo5
Udp7FVrtrjeiWhlAYAOLH74X46z6POcg8pbt500qs5SSBTuLZhwfYAYPCWk+GodR
eMJ9Z+Y9lY7a1cJyMloWPeeiN2SAcCCfb7DEB2o+/cNZIMRGVcwww00Ncg3EJ2Vl
4+K6Aw/jElV//8KNOuUO54KtgUmi8GHc3JThz2IGwHbS10q3YSoV/A6CJJYlm5qC
22D8atCC5k7e3gH49ZPcAgbxT3PAJ9MqDdAD73XRqELa9A1SI8Gv96r1r9y3a2g8
t003Z7aRIXcCuS1obfJKHMrJroZ+jn8V99nc8z1ENNFFkzzaR0EuKTVz6GBAw3Oi
49njODFhCGw53cCI56B/ED5UD2E7kr/4dkt+02o2724Bs23tMk4lcBM6k84vJH3/
RHsXiaL874K3lAZRIt5Njvf5uFlg/DAgBrJeH3YO20L01NhUcblasmFOHhCm8VPt
i1nn6WftAYplA9yXELl4/AMo/lSIPjYM09TpMBIvEThYmnW07nVZQEEhNHGaxDLA
1BJSrPmGdG6ZEeCHTqcl93580yzdOHSQ1vZS09SrvvY4x+UwrEgO6jgVQ1tSa7Px
sV5F8nJgk0TwcEpW8zLBoyGjobnyr3I3eQiW6i6Wvh4bBODW7O+/6vk8h9MbEtr4
0+7yCr/5qj8isClzttMV0db22WS6N43oI6VmG+jh+pPrWuBsbdvG6jLiTThau4tQ
KChbDc5fthap3UOcuflCh0jjlQ/tmEDqiL/vwFhc3P2MhlwzqeNyBHt9+Lm9V9Kk
+ntdXPvRYUcAcowqsDsp+3GscWuGjjUDXvUZG4j3Bfup2YNBydXWLFEzKmeKW2sY
LPMqlYpBREs48n7d/d+2oBgVOQY+2SxdziG7KrRKDlImWzl90febsToSLwEgo0tw
qV51U+zNgYoQY/C/FCJaMfR3vHYa72ZvZH3GSYOIqB9fhLBDSdvVi++tHNl2r1LI
HUadodKnfnt/ntcBOyozoRY7uweMBZSi0wYXWO9Xb7FqSMdEikhfhDfQF/X+Xc/e
fMF9sokIsh19SSoWqR7mjckO7dlp1DTM/IQ7DgeGQdiBGYLt4bhREPvD0ag8oHwk
9rigHffxT7XSsoFqKHFmmQC62fAQyCZuaWJTpnyzQwK4oovYVMWTqw7kBd6VsqRo
3thF2/4FPTGbdDTFET+3UWiQ1k2MTbaKgrg6TiZPD7ooq+yYhBjaiAhuPL3ZgBYr
82qPBdOyYZ/5hLlI4FVupNzJZKw94ui8ITI/zi3WnayFWB7fivhc5Bh6Xg7OhP4j
zjzU3qu3A8E9EVhrCr2WOHbYdTLoZDVwNQ/Qn6FLFHpiJQzIUw00lkmb6PMlELll
po4UP/aoMYJBEbD+LGWJ+dk1QPlA3dO1e66171gz+WzVv4guwtmTC2SFMuszbh8q
c4jC7X8pmv/aKh38qrTkzGr658ytXIQUIEw6gFNDcrmMjRWwBrniH5tEqaPlNmhy
l7G0D51vXNx09lcGx4WjE367QnXBTy0CJb83ZgyCEE7rIx662r4M1nKTyNDwzzvn
ryKXZFCAkAKoHbSz6NS81JsXWHTmSNusTH3fl8A1TkoTFW2wAW1JYP+YoAlWLzVZ
Mc3ERVz8iXwRl1Kn0HoWKOApb3Sw0eddg92iX2CvQ69aH6IjHZ7i0GEnT9z+uJ4i
VGa1Hc23wXyRRbPNLg9+nw5pDQIg9d2p0zuLsjh+bU931EOIpXRhtSXfwAEFplU9
qfi0hVKIIiDZdA7xuIQYr0Kma/Z8PkwptjhJsgC3Q/OnaFEBnjTklkFi6YuHBq2G
1PTyGNlWFfK9D9dihCtaB2AXm9uwjcQSfRm5bnIOt7EpjNY9tu/4pHcSiQffK5Cv
rIZDQIqBZHrT77rE/fT8V63FzdnubVtSe8Pouuirey5KMld97ZHDS04FSpRqMgFA
te5EexkIY32XaViIFQwClTUhhyceWpBfSdkF9V2HzxPvXAUzZbUxQTPKllPwva41
lrCkybLLOw+EfZSGNv3+5Q6Pm47yS010soirRVEWY08V7cj+nt4zJGIBlF2HvTaL
vRgn1GplUrn3FM4TN5FaFk5XAlIh8YR55JsjX3CcJB7afBZlfL91iJJDtgkw1lh7
6UQ5XhC2cWQc0k59qu6FcFP6RAr/rHiMGVs/Av1y+0gaVEnxnG/TKnyHpiRNe9F7
sUOzclYX3dsOH9mXFOqy6KOBF94XOPnuZ7OUCiz5i7tZR2GsiMFdem5CtIqv+BXU
CU8zhfIH/rGOZ2D/Qj0eNPKjtofSUDYPapexijA1PxFDWRuix/r5WuKAarBGUa8p
4GtzMXI7reLQcNmv369qtK5zxmavdHeR9BKu8VA9/fVdauRvGushKLk6bGFVh1EN
TRZlYrLYUXfQpDjACt2xYOAHrPLNmT2Jh0X1Qqh57OUObdORcbE261V8dL/T9f4U
i3o5Hw7Aon6Y/1/w0orrEq0uIrRpHIXRAFK32WC/8XqEZ0MTzGpE9Oy5WlniO019
9WSmmnQCX/BIEzCy0vlc2ktuZNGwYNemg708zTs7dJBooExyVZ7CJEzXLjdEdL+6
IVKEmt/U1HttcfCac2p3CyK5iLr2mP72pd52ZYJ7f5GTkTFWVtpBmoDVzH8qP1np
t/k7MgMdzIUefJ2aYqZim2zl70pg267ODe4TS9Q0O01vNpVV9YeneL/luZ/IeeV0
vNoE5pYYqkOj5n/+5hXisLyYfRVN9TzOcyW7I4DVMVrRqubi+qz9bxjcy1cyXAxo
LQCGJgvAT0KKX89vhNFdNnmHNL0wcPX+evPQctq+Q1E+wtKD1W/349U37NG80Zdd
tzZdNhh6QZV/+1hPmp0asZJn3uoVMxzszoYLuybTNo/5bEwlmhXdo+RdnGR1frdt
WL7ob9UgvvOIzUsodonhVPvHRHewgAfw4tH9VAW7rGOlrXYNJVqfYmJVJeuKBVMY
wSZCL2QJ/+SKbyHFAvMNsfbsvFR2x2zt6nlZqEEUlzEj/g8izxxrIfmRB8pHf5X6
PNkL8xWamrcHsqxcBNpQAhrL9pyYkfRFu2mYjxQkfkq6ST/BOuJyUjKOF+kwLfC6
Ur/N7bn99ml7ebIUtxqj5W22Om0Y4oUspgXwrLFBbpOCsExtF5EDq4Oe86ty6ZDr
4OCl2EHTbD7wWYXxylHy1WdHSDk8yfjOSkotjqLZ87awl7dsWU8syydpfbHFaF5S
vhJMTqnVRVqTZo7JQscTQOopSFEub9daM5HIUFyhy194mOsWB5WYeWIWV3edSsjd
U3gG4726cLN10ks7IrRrTMkkEPaH7xf0Kou4X5BKix/qoKvJCW7CD5PYeSNyN6Uk
az9Ply8rFbMcRmFPbwJbuEiUuTSrCPUmNKoBsZJaU904wZTTFFgxNfb2DPMvdKM2
izjjaQOtUvCJxrlhzojwOGtdXPUIc2lxJmDHDC0KVg602tS0AVXaxWG03kwLgOsH
ZPr6D1qUMVIeI7DjNzBYQMzFVRdym8dCH9u/DyeaWXd+4/4xMUq+vp1+EcaaguUF
V7x2+ePeqA2tArwou+E9r2zRwF3K+oMG9XBVhZ3nprfIzfZEjMtLZtYSuaskDCLn
vTmOEvL9RtcfaFr/GvWZqgLLuJ/f4bQLeF9aWmnf/VNqsPwlLgTLNMiGmWeXv6Lc
/XUay0EUnoBzQLkqUcorDbF4znkwlkp0iOZ8mn+3hl4J13dU2VXHH/naMKZAoGKB
oNiOGxbP6FVoARq1wY68LEIiv7aZ4YTxYlA8E+eNGsHwuawMd9b1zvxEnhMHBZG8
WqG+1nFvjDEvYxXdtGMh7X12VxNMbOs0cszksvULui37STpA3uxrNHFXkFnY1UKQ
9ZZiEzZhhYF/mVwKlr6p86R4elXzkpsdwGSpHzW+4r658YyETGvF7bAT+j3KtJRZ
AhkEBiIvQ7yUaYXFXUZzb4AI1Yn0vziusuxyR1V3CNNIfxzg5u8QN9yckr1wt+bW
jIDW2UuUk9hJe219FxM3NpWX3Ik0lTIZ/SseoGBn2PMMItOaAQdxHAaEZHORGr7c
A5Ic3YeumY4hEuDOWAmXCuIjBhuQByXX+cGxl0BocSKTnt09KMwYSBNsrKUYVofh
NjEgPF4DTWcBFHn1t+aV6EtrP3qNr1z1I+nUv760cZ2K5ikk3s3r0WVMrW4Mjf9u
3nxPCh60wS9LnACKB5CpndvB0rCZlm/JiQ+tSAN8E6VLg5dwpHMpStcaD1ZSz5rR
cpnlgVlLVJurvBJyV1SAUYnBuHvAcPjRKWln6AcgFD0tYtl0qsYMMcwiGJBzy6WJ
VpVY8UlgSKyFyf0OivCK8ATQEXlAA+n4jFcBx3X4fM0oJQsUnayizoDHnnW+iWtP
P8GdzvFC4gF/OGvdyVHTZ/Oh1wvdkwfVI2TVX9arl157AuV/q2fepUo7KpmPREue
seV9z9H1LK2ZhiKVA29prj8dGAC4XGJyF2SMDLqePTBS0Rh1DgWeWIInqX1xiCD3
qWElDnSwYgOPFHK/WMEHK+muyShpHbdLgLr/pQGXk4tAiDja9D/TacKi2ToaQTMF
YeI0nvgCRU2xJVGcsrpF9Li0Nd2FUo9XtRwGIaLfbc/6B2l/vYWbVYgdtDDcnWfx
lCfzeDK+VWPDWvf1pGGAWfJl4bjhd73ly3BeTzA/Xv7/axFF4fyhnz5+flDiO+11
WEbK8cnB9S6km+oruhUh2+vpb9pVTf6Y3rwGUEfW5uzK+qU4K1fK6hdH1f2hXK8W
2p75d8CZVxFX2JJgwFAfFKxP9uwFIMSogTqqMBhD3+G6WU5EaOtwmKBdXAe2Hv0c
IDY8ZbxpdEByYYI0heGu5OIs7qr9qb6e3k4fwY3Slt63T1WQXX9O+T34EwzEXE3h
tETf6vCqgHndnn+xmYqbSKHu8uGUPoncM51nBvwpmXQsQD+P1Hbppvh3AbYfI7jV
zoFWg3LhZO2LzereY/8FxSxFsxaUWB8qgk4ewxytCy7ZBtOoPSIJfHQ5YZ+OIYj7
guMdcDvoCoanrBnVPk2jUtsWomqKPshfpfvkZkxy551x0JPYcIGEi8m/mdo37wX/
7QbBmaFwihaFJCLLxlcwg0H4V/wsF5eMiv5hbnAfQUaeIaq28rCpFJPpiP84HRlh
VImgiXt1x4xbONukqWWo+rUvaQ2poVXEcpxw4KyeqInhPhOqimz6JQnxY8s2cJDj
HYjhfZYUNMyhS0xGZg08+I5o8cQ/W0L/tGt31G4SBgBe4eqGPh3s6QCEtmLR+X2X
66yA6YxWahnjZEjD8PFZqe5Jr+bfpN6SKMfxSMcLxiExX6+miLLn0a77OWnn4gTM
qaYDNg74JhZ34V9/ZDu06W+rbzLJGuXSR92W1aq00jO679XfGu2PmRs8I3N1ogVc
YGeM37xUp9hb2qezMi/mlCjyA2UD6aPSAB+ZZx1nl2sjmg6z7FRBYtV3tR6zA6al
0/FQVMxpqjdzc9fu8DEZ59ApM2j+Cs4e/TAd6a/cPBCG6SfkHTH587x4CxBWZp6H
NAQpMIrdoDl3Y4N2Q4NGFBU8lCmR7VcNT0BvPvnlkDM5Il230U7L33uS+FLkADvX
1CblU9npDsSCIIdba/ZQjI8PVHKP9W82CCOIF4RcobHHsTavVnmMEuM4Y9vALLV5
zBwuJXrW0MqGamI8vyywC4dhOz3zYl7RA/vEc4hEZMLq5mhmokBZzrzpkGoq7jjC
W/rMN6Ll0MPyw3MUQp8xei7VY/h1GPM3o3JazAj3Z3jjiMt3dwYP1Oa5xx3wOhgZ
5CiGxzO9v2K8uI4cZs3PzzlNKHdylJCuFmexPWBg1/4GisAxRPcnI4GM6sQN+w/e
tW1lYf3laYnKpCCO6HFTZNBX6waFE2Px1chUEH9PJsarDuxC3/70YV+YGQ6LjPEQ
FGImW9Heiw7ICzpQaHnr7k8p38slmJOcrLmzARXzIXo6bH1AnTuTpsVkEwlssbgH
udTEm1lKqJKmenkVCUb72c1qFOgjLfZJQFRUz2JTfVM48PmPdZSTH5jqGigNiHre
P0Bo36/b5bZF6TPanDOGje0GUTUMImR/EMvxrVvrIa/p5Boj/wzTM0BTzdExdIFn
uyTIAyGggcsafsudjJNPFUYIh4uwraFj3wQ9Wds8T2JlmbgQ5L9qFOO2gOjLD+5v
lnqQCTEUmhY3yy2kri0kgF2weSWb6yRSYiIMJ9CGgq8WK7Be0Sp8hM9Qcx1wx7AD
7zpYqWN+vKEoQsDFUViqOO3yaYE6+PH7MQN7XcQjZRLAwPr8Bzg3opR7x4d2SHZ5
86luArfEfD/QRQWIqgRfwWPQeKnM5whNvzJvZqx4Mj/hS5OxxeZDj9NIAtasdQD+
2dUuypPwr755NX1JtRO4xE5qmYkEP3zRkSCMR/ynDLsMHC1UId+MWpQUHNarwU8C
TqO3Ud9vk+OQtP4alnelft6+VmRJ4mdPfTEJgvo1gVIhWRw1ueMoFxKgIYuGY+/5
35NSmcQHKLWEJXzcGhAvxKOgeEGdGx9FyhXbOq+n38xzq5gsWHrW5As4+VV1zHHV
v7JdHnQlfmip9f5CCbiJ4xtDHrUDvB2GSfXi41Psv/rYzFw61wY46kFNhrVXZCHN
KznsrEkWXFATSGP7UZ65izLTJadn2yu4hnlIXBjagow+Qq3/yuy7X95BuzRVr2Q/
IXv0yj1OOPGXcN+d1Xfmg8XXjhlUAKSUlTTXfn6wzEG7n32gEQyjJzQhwKHcFbY0
Q7Fl15oUwmhHkTyr0PX+l6GAdSJ+7WeOMA6fRPVQDF8eDJxqWA4UndphInK39V1L
tzBAFfjVeQy62lII6aosqVwxLN6Mb+kcLBIL8Z6Mmv6Nhm2kRMcZ7be+tvpr0cZc
75HfIZkz8ibT9lTUrf3aPk+2ImBwwDpEnbUofdjWVTZmUxhggZm1Z65gtnxDZXm0
9eGMdyvGoRiYHs7T1+GgDMyPat93QbsQf+94hkEl4XaxrhMB3JwLjzvJivg+Mg17
oNyIzFEZYmb38zpavcyLQ8gn4Ixv3gXVolbqcYegQDyHIEmM60DaoLbH6ive10m9
pqJDx2dMjK/w/uFK+RKoU2zQOFv+7OW6xVwgSPh/Z0518or3iqtCsBkFirPycxyM
HwkCNUiWGS7D3Abxpcd8GS3kZ0D8O3kF3pA7FUkM0P89ownpNt8foipdZr4hqYey
x4lNstJYErpOJT2c73uHXiJiaKTOAXv6INlG8ZusrPAqiNCo5b8TJNam29i55i2A
zK4mHcre+Ij6CFdqiNBTbjZVHUnsJmW5SYjd9ASPkNKTE9qTjXWl6+D0NAXdxE4n
XVperRqkN2nEHhhKwKu1BKs5IApa6Ll5tph7hcoCjj/hordeeF8H2fe3vJkrAPFE
CG2vOb3msE3TNxiAMoNgWvvqBFCfEsvP2v9AIZZROIXbfbhNKxIs2B8EO8bYPNYp
uptQYQ8wzGTiygQXkwuGtfgDKsEF9AMVzzinmnzdkVfTiP8WYjumcrruBlWXVzpm
03pJ2xqCl55F9q/4cTgbG/mAvS/nWq0BqvH7mNxnS9HxuXPwHJoLxJsSb6yzjLC7
dAaDfKp1JUDTjkuBT44BHe1tPhvNDIhNXy7M0YOk8GH1EL1Ft0BC72nvyn/YCRtn
pbi1L7J0eXYYgSPNlyKhDJ63/Zn/QhD1NgktXoqG33RTUqyx46qMi3hFMjyVOCa6
r1YHEgQrkp8rELIhydrNQEm+e6YDNa1j3aM1Cn93KfaoEzlbCIfwS1YzuB1eH72M
b5n6tX/nCqrWxD6ZDget0yVApUQpP0NuMLNKTkzhe/lfbwgDxfo2vXtgkXTqR9rf
44qzO6OKHTKbaOfY9PBe5t3OxfQ5jxTJN7VsFbJKk2OChlWQUzELfdY+2pWPzjDG
VqMERmc+OY69M+uVKTaxjFWHvuuoe5juRVPld5vdC0PBZiazrs/PrxURWsysezOB
5Boe9viOIW9yDQn/0vqrPTiEj9ZripyXxIBIWNDYcmvkI/Pwa0f9TddNZZs3ysOe
zWLY/jqJEbU5dF6gSCjthlzPwjq7k6T/c2n/SkuZK0P1W9oKhoYBITmXcbKSM7F6
SI8ftCwAVLH5Fh62+VVb2VBqdXIe++1hmww9US1rqyjhkjqbkQ9kmx9IPZQh9MRE
bYGwobr/lWmYLYSmqxaAWIuj3ye5Ln6KDJyWKtkAsuCMVSpEI+Di1Eu+ZUGynU5Q
AOAxYt+96XgAaCHRZNgw8wqE93KEv2bCCaohLSrB2mXmCSoQJyCNdzg64qC1/WGC
fluK+n1SER4s2TDjDxCDkyKSkTDxXnqYmMjcvr+R/yb9AN5ieiOPB0BCPAvUFoF/
bg9TQG1Na+bhDjdLSwDaf7LEDGurJKJtKN/cKNvo4LHg5MwPeeE1ssH4W2t6EpQm
MNIbmQplqcqFpippW0lAVv0olZP4NqKs+kKRRAfGY4sn6lklW08jQl7FHLDWQsKl
9bHpqFdMjY6rJBlrDaNEAOhUn7MSwv6ugnTsJUrQ/md/ekWxMxBs6gDeMfehcSj4
DZ7aWeheAxtYm4kdhS5iHcgTKx3rTK3OR0Rkag0cD98BlweuJEQS0Jc7sJN+qyi0
/WkUntwrjbRTqnUhnRPLSBSDyLQ+y7vbdPeQqm2UoUuGoyhEgSzWMUenSBf1ctLk
02LCkjK+iL9nPkdJlEhO7lt728GKv7Y7kiRNXnIIU2x8cd7gdwPcpCCgkXP1PUpv
8/Sbc3gxQ4CArm1iMNfRWogf0mJP2vPR3SGJq4gWUwItCtkZHv/aU7q5ryc2YUh8
7Ni6RyQy7LWv6cx+i6XH+UuSit9RLcW3aoJCA+0m9tTlo/WDVSubfDxhUxGmpQad
dsIT405aDGtuanNakFqKlWxIpQ9z8z8IySwHK5CjhBxmJBq6wh4M+e/rAA4l5el+
apeyEzMmF4BhsMvKrcXgINPv+etCcgG7DCEiEZ53y3fi/bPPC9Ue4SQF97VmQ+eX
15zMw0ZL+J21zx2BIzSJ0eBT9IhL7+Qo7af7PevLBRoo2wEPgdatZbwDdhySpsDr
9i2X6tDoFCxIzehdQCZ3+FKTNePHiPfpw2kSKXC1sxRYfY5hQ3MMNiZE3QaSUSHq
4nlvPEmwbcHe5tC/32V+/iZhhxSZRKhAMV8RZPeomgGvB6DKpQppLVBOl7sdlj9u
etI8kOHhgavkKqc2uImMVdPcWfBDfngziJid26Qm9sjdo/hhd8lFGvxU7/XMgtnl
TXSicX8YkgxtG6Hg+4sc3+3Bx4+Q0ND8IXUDa2VXD3ORr01Mom/yNIle/zOf2tqV
1W+KUmEBAhE9i+NGqK5ETr2YP3OIxaXg742O1SBnYjG7mPvEOpGDZi+4tvmOz0UQ
UHkbF0Q1kXHDGDoyGwIGUz87X4qPHyLHi8jGL3RpWqE71hL9bgWozSLXobuvvOtS
x5Q0kusnnmnCytNw7O+rcRzgnCwGPJRR1ZnUABh2V4ycnt+sR1Sb/UfzX5TZNZrP
18z0YF2VvwpgnYveGsbuUHBCMEZf9ENc9P2I9AAVGwosPcTZqOgnSXw4ecD9/PWw
HmWKdpXrXEJmhaO4xHVZk9YOWP5VZM+blLErSTOmm3agWDpNSsaQaZ+0KsimW+Pg
lLkNhyFj5l7pA0KX1bfzldM4yr5ML3at61P5Vd7hOM0tssV6/jv4ReD/Rm7Tr+AR
rmLOeDiqDbisZetGeX8vJ2jYZIM636Gh2AF0HVU9ad1WGZutVFqYY1SWSPUATNUb
n39CiKHw8V0KpYWDbCaBUK/JpEn83rIVUXGraJCSYmqzlyLUMP8DZbpyCfSsEwaz
9aV0NiJuusA0gOViAOSOJE+RN9ail2fRf9eDsXbC2l+go8ZWP/G5pVMkjco6IfMb
MdTSNVX3cFY3UwDtRz13eZySsqgEoCFilrDV4gtf7JJ+xfGpjOOg0OlV5TNTYtOL
5Hv9iTwOixIQ7wVeqpIDi/jr/16yqTM20+PKkptXcZ9CccOKwYyRn6sNUaEIsf1J
st15Pf7MQAPhe0HhrwpyDv4WTyo8a+LNe1CLtkRM18f0rJ03BWcAe/k8LCeHU1X8
Td6xKNJ+bJyNIiW2vaK/mRoPHx6diq5L2G6Kz3ZLP0LnoWlSqtyDKaKT8XPn1yuX
VUnW7a6gmgj3utk4lwL1cndh2JayvWpdnS30uyTHokgyIUNaib2fetCF1Ik/NL0E
puQ+3i3W4PtolT7AMD2+OnJxuS+2x+K6mQHetIIUZlTfF1FTPzjWib37RmSWI0U8
hXHcQYpGRbu1sMduEG0UZVcnT50/qpI0HDJXyC0P6221QHiBGWqXmD0OFfm7eOs2
CNNolC/3EWfaxgmRItqSKFNMNAfptIMiarY4p9cNPAe7C2aBXdhjoHRlDYXdptdN
6E5+aAr4/0/gbxEYlyiXASbK3FbEZsskz/XEVgNlHqWG3HpNcAMu3SJ4tTjft594
cqG5pkwlxddx4B/P6woF29aKjbxHSMJGw4ZWEYn3CAMLB5VClaJ8KsXORdORU0Eh
3b5zmGdX39swqMjF6vxyr80K2uCyt+OBq+V+SnPqzqhkqfO419yl5xkdA1gUABE3
iCHrmK1v8vTHLqJiDb94w0RBB53Haz2XmerpZE9N+jTXibmsYGH4a1jNdeDrCdJt
s/9sjN+9o9ZfMF/mMA/xxKJEsWDAd+2m+9okoLgultO4VOVFq8E2bo+dHqCbzLeY
0j2TGv2qdwJitGnB0CSqsSacTEvG2Z8uB1LCsSM9fYQ8J5Tu/l2+hYDR69p0UjKz
aUs9vsaIQRav3ZW+GgGLs1cGoCpxn8CNcVqeWaAmQYM1dCcwUPw0KCYja5qvvj55
dGsJK1ie8+te08PHKT3cWGV3A0ZJ46KWozppTZBNjSf5kuYeZ0R6RnDdBwpvCnrs
wW5ItxWhiNYv9jqLF8oM/lkcmghmShlxPeJr2/2KJfrPKCw7orlfhH/uKf86vHLd
mqlkr4+1O3zusTHGVHWWzfwIwJG8GcKFykFeiOQ2xoG4jOe0ecLUTzzNxMTN5Bc5
SzzOWJv3NNVAYSUtPaynaELugS4JTpOvVihQHoCtEfzxl7UFQf37xMtEJ23p6pMH
nJOrmtqHp2OuCQ7rs2Ncs1EEM4hjAmv4vSiGCGVx4iQCFAMxcJRtF7hd2hrjh1GJ
1QXK4G++WjexCNLLf15ZM15Ec8eawW3HK676nQCO4xmTAVYn2qCBFteaCyY62RnG
FPAe/oca8yPUwlTRvnYLyxQuZqb8ga9E/vrfKQ7KK+URwXCIYyhGLiLbrMRBOmGl
MB9rdHorLb78AhQPfROSiJvxj/x0PfbRNlC0VtMPE3O1tnSVqIhFPunHEcftmUPu
AKmOqht6hTajmI991Wne8FW4fU9ef54ULua9vzLXJi/0Q/e5xEeaSFUIO1n2NVHV
ONc7Y6T5S8y953troQ96AzNMPrt3BXhlhSi2ZYv8wkWeHT3s0xdNeprSCSWRgB/f
M4V9ziV7rYtV7+S5OsAmRivGZDcA8A2A7Ovf+qegc+GpVzPNbPbuZL8d36+gsWBf
T2JYkOENKwzZ11Zr1z6TejFSA85F8I6BaQ9aNnblNISQJydpWPq8Gw/s/a0w0hDE
PjT4zroVWHBXqv0bXk5y4KQc4okhcyewVPdj5FaGJCl9hfKIfKp9FM3wrvstZZAp
yb9QSOoSO3LyCI0fmmJOyeQ+mvIkvnNfwUsRCMCYWY5WK879B7n3pqSyvbweWVXV
Cc67oyHBYKuAAf8FjmomZZQAwDmG2NglzZgduV6KfDnrA4xp0BcK9xHnmslBrawu
Ay25S41aqu6asjtpXf8Uu6hMXjQ+qQzt+bJSCI4FJr0jlPhJC7AAefd9Igi7Awmg
7V72I+hzxJ1v+iS7RP2TEvyfWyiFXEIYpI3Ke/+bdOkNSEqyAvjVwlpHQPwDtCUa
lOXvQC2MLB5cyGDb9JrqaRQWP0r1fTXwLwgAvvib2HOy2lq186I0wFwP4DdVmAWn
zUpIy+dNwjV8UbTB5bTjFacEBvqKoAuCxwtKhHoQ4kDAecTGAPmhgubMOwrZSE3I
+GjAAE5vUgY3e19u229mh+bwUFyTL/7XMuCOCiDxsQCsu/pJEK50rfSoH4oRremY
OfwADODjteipYLpThO81XCh4ejEi2oNWN0UA/af6yN7hwDB6cC6gKKMzgYR6TOdF
xVjzuCJp3cQRyfqe6dW7f/tWIhjjCkCARViflnWK6kyvCySBYwhXydjpXD5mKmnV
svxn47Z8oKKAXZTC5M6Xyf34iBQoVHPBOe1VytZ8L06iyHqBOQdoiEFqJCD+Jey3
Vp5FqmJKCy54OhFMIPm/QNuGlKCkyjCufCiHE00wgH5sLLi/oIc20fu5vAL5PRzW
5Dnsg1UlQqCSdO/GsmoVK1MKmo9gPuT49zBavechCFNPQ2v3nYfNpTyRC7jXGHjr
S4az3MPE0269ANmTMsydiPXhCkS6lqltJJyv4d/uD6ODQDC1vbCqvt9M4AImGvXP
ZEDznVoyuum86RDrA3LyeFYgIRaWr5H+Fj4iPzByaRaDHCtFyZCKuBGrfRQRYGFl
SPCaGINW9/u7K4Db0LGgsYRZ9YSEp25snUnH2mKc1bDNynXi1UhKMxUk2BruZH35
YsXNuBZ0MMhdc3815gXGhOkPSs1mT5Fc0xn5YFYALIzWb5INCNokCAuYgN14Dtp2
lesBWmA4Jvcz8+qvkikav1+LwV9LnWE6D9gBQYqoec7pB06P17nmiGW0VTQitbv2
GW3yRw3phLbKos5z+tl5MmriS2BP6aslC1536YfWdP0LGwwfsrv1J04IGBRZJYf+
1oUP+byivUbYXhn+UrJfAmfln6NcN8YXet2MK/wGhu+JmssLgsa/uhBapXMvaQlz
QR84r8KsTpw4egjICIvh/Ib0dGaKSsZ/9Fr2ajvbhkWI4xrsCSVbygsBjQXSqE9h
NoxXmYXTbgcOyV8X/ZdGEhmzYVwIthpvzulAahE066cgg6mQ29EhdW9EpNzAmfov
UMPj3b3urkhh0ZUB6cM2zgFnYoLGQRz8gCkbH3xt3PJhj9ZvNQmb8xBxLswwrbne
XzAh8oxiwEmNnEHAb1G+Vo3avHWYwf3BhGxgfkkEWwPI/PF0IW/6u6oS1mbmXSMk
fgtzaC2PPO612l7Zjwdm2kfpbydVxfPrQJ6nfZEHDXTxxHroEsTmFZsb2e/KcbTr
RzkokohfLZqPR+3ZraEszL1E0vspM1O3LjEQr5E8c5judOcZ2UfErrKOv6RHSlvQ
JyPnaCeuzyu9PVbLkv7EHqEgStpQEbkiVQIKPPSzLwVpgVy6SKZzM0AINg0k5pxt
TIV6lDCMYcM4SWGLCr19ZwRNatNhGPL9W8CeTWe+BdteGeKI4dwdRjFF3lsxC7Zp
pETCnHB6jlkNAej7pmCQnn3OnPEna8PB7igh7AfCOuXfqF7ugcmyJPU/zCIwzMSY
E44RJQ3JAtJb3RLDkYstzy95ZfQe7IDsg5ytnThKiRfuffESJULGKN/YWD2KkbG5
y+/NhKEf3i3J0zfFoHfdDg3yswvPXbSRyWV2IAR9mJTg95HRnttOx9Mw7EFsVKiN
2mK8NKAOUrFSh0yAOgIcdihcblC9vK8Ju3mnqeBF+r0MHQnEC0B2sHXYutqnBqzI
PzoP0Hp808K8pVPkicQf7+8CD6rf88EQdM5c0t2ViHVno+72lxkOmx0Vk/EmE7g1
nn0iiQXAL53MKV0MNvS2mLsVCPKrRp3Bp/YmB+ESHXM/5BglbZzY3GFjwImqeKRH
s4lgW4AVycqmF2R3Vzc3hBDApT47B1So+VvmbOyTV8xK0tbgKoRUOXmBxVIgsYou
bRJa6gvR6lyc8hxgC1ZFy/R+OZGdXBSo/T10rrrTP+GUDWrKEwWMw0cmMDmFqXbz
aQoUl+pYZxIaGVfWlWNOKRr6AQVQGwTd+HsCj7DpUUuY9Qirvx7BDyCp4fW+pxnu
jwneFpwSkCSyxkzyIxIlyXETZpHcoaY1fsThZ3VjTvpOXAfZSd9ldn4IVj/GQfT0
yahDEO017AzPI9hOW7OKtMFrkOCKS9aHsLWdgZapY5iTCIyEc72ioCYpHBFlb1uH
4nT4XaRnRA6lZl/5JVwl74MTVOdOLE4PpjYNRNlfhxv1SQ93md/G00A6T1q9bH0e
1s8Dy9xT5c0aQbXXFymMjRX8cc0FNUAKHcx/R0zpCG7HHB5e/8HJ5WSPRs4MvoJT
b2CR1/Rh1D5da/l/xveiYnXPESH/LnTLuF30dxZ4uxlH7tZNzO+UOZnYhW5BAYML
+8XBoZLVi1rMnB6AXRNGXyCZaWzBZ/ol7hiLS7tmUhWja0whs1LVpbZwhbBgKsPb
U7NhNjeA1zfAlrodWeEbg5jeBlBzOufrqxrzGrVngFACyJmi4C3hxJtt3O1D/qdW
Zn1FkwrUfF5SYbbHAZNODQip56h+u87I67k5PcHydqSvbLr0/2+2R5gptGIeoSKO
zzNuKgg03UFIAmgz76XYFOZGL5VDCocyStWkjd9syrdelbSDHWAT70Mk2p1pD0e/
CkwGlRDpZLkAjDYzMoMtp1WU7XeWZbQGaIEOOUgISKim6wYLkpjwLEgr/Hx0mNZh
pR9x875q9tTYLd5Wjz4V4SItJu9e9IBkcMA7XobiTXL/2xdCiCDvq+PfhspfayyB
z3aRqNC/+uOW24MGWbGfIktrBClGoIA2xFi+Ii2xTHu4g0FskS8SLuubNYw4D/vv
4dHD3T9/mjKEU2x0rUhuAQnMdFtJRzQNYcaZFxb3emWgyNSC1qJKvRCWvRymqFNy
0jANiSsty5wSrdE7ykNUL8lMvD6TpyFLNZYODWt6a02epsh9k8nFoRCJll8mo9Vx
30gJATuYx/NbNfYLdQs7PGwuI1FbZhX4q8BRHMZezD98IehPcAJVsNpOL26aefIs
fsPg3JuVDdtUQnIFdXhFB2WPQ/twb2jjYLbrJ0RBZDvZ8000l9Ks6tkJ/opkomvp
MKYj4D0UMgPuWG6Jn71TkdL3qmkVosvGCYtxR2N9Enbp1V+13uGm8CA9Sy4Sp+RC
DBNQGEdMgaWEF65BLKiFSGXJWWsnn5LMi50Tf0Bsnr/c66eFm4n+Y+yNIkdb3d32
6MedYmrQDZOYwlkwvhEG0BruknY6OcgoFeiZiJuEt6TCrBGo9wPvfSsNZ8g5S8lD
dK1EKm9m0t/brXayHY4Kvi0Zdi7RxKPn9xRyXbVV/SLCLrEiCYLQZHQO2rreo3tx
hFgom+C0CSFKKw/vJRi4dZ0H8skiLDv/raZ27r1XDICa1rO9cFUgjbTOa1bxHML2
4hVc2GeIUU0L6tRttrhRt0f22dhdeyDZuTKvXe5/xCc3gF6tfRmXcREiUKhB6CCL
Ayby/NEcwEa+puKB5byyOFSR++EOC20N4uaK4VF2rWIARrMHSv3/CLug7W2hTD1a
4HHGxu7LyTQaLqZQsvfXR8dICl1U2Lvevya8Z9R5nWo4EnM3MXB6A+82bNLQSO2i
D5WIDB93a6gzWrJTfv2CPB0cP9989zN0wBt7HDSCoRM0InifX0/eP809HMedEauf
aa/V0yiqoqZmtrSgS2Dj/S/f6EvUjFKUPYWG13TLP93m1PquI42FhAJ7fS3aJSDR
P/NOTSN6DhGPGKVhnU4pKhfSzrTppMfUZyOWhWeVLewGva7im3YKL5+YGVCiJ3kV
48dM7GbiUEAuGIOCRG3HVpRgIsDcLCuE9x2T1117t9Q57Z68/tcIt7Dily9zqU10
/8S+5IvdR5t6CKtdFqXXOZRYR+LK588XOcl1WrgkFIwCJNii633a3i1J+Gxiei0b
+oSZjuhdbrx6gzi63BJrodN1O+T17uJVZR/dA4tf3/vy4TNvnx5qWdYbEVphfm3L
1mifuV3IC4RG1bWobZgxwqIvVYwIb/m4ErGncT45X28yZMwY179lRh+OlqJlxyWW
+ATj/OT0dQbzxAdgYLsYoYUAKUNiof8q25OjeQmwcCqz1et+2eUSe8zlqPadNBAz
d7rGJUJH9S1XUbK7rysd/ArJ9rEO05ES9hlVMuT+CxOKFaNHRe4dfymT0ul+rGvw
SkYzmIctD+R4HPw1Q6IgHr2QKG321lTWtM7xNJio/0v/TSFZsQADITw8TB4BnRRy
gVSnN83stF2D6y9jErEMMTCaU0OSgIeKBHXDPa+xVyWelDSGV2W/w1sauFB1njFv
DSuOlKNmL2ua04/jiqwfpRZ/qR9j6brBONX7V3CRHg/PtHtA2RhyvvnFiZsHcjFk
o2fuP+Wi9XRoJZdbnMKhm03xecTOL73R9UVnjvO8ssFaxXjykZ+Wt/mQCODbqjtN
tg2Ag2q9W2OaPBCPHSZOah7FKM5uIBXuxAbBkIyjrbfsYRUAzQ0SaB2i0mmFkR//
2Mi+WF8Gt4l9MUuN0aV2jkXoXzncUcBUbf1y2tOKpDwZut07YCco1YHmD5Yv8olK
JaBOrBXRrUSk6SeZuz5Xk/L6Kr6DiYQc4gL0pFRtENsKsRE6beafx26njP2pVhyI
KxSpuTW/hO06iwfVzBCnChq42RpZ0rCCQ7hjdYaFAGgoPOJQae/wvrkrUktqzb8M
OELyg2loUtTW7DP6UKFXRKPRtdcpBrZh/0wg/rXVIfqGOliXdCgXDCNDTnwrKGOY
oEeaDqArr6GKJiuONhTH5KmhbODVmNe5Y/ONy/c9MWCM7srkpFOCHHh+/FN6Qe2d
K5uzZg7Z+ZZAT8B0LKt99QnAIKaRERpfUOBILUriyXqkLAqW9ZghKLzxuKEezWtw
jZd4RuWH5u9PV46aF5lf4DdqE5946vVO+y2pXe4qHDzBuYGnkdsDy3tZpT/trfNf
B9zYNk9O6fdsWh3qPjbOcjo13lWNXI4Pq0J0XxNB4lqwBklGljh78O4NUbN0N7ZF
koV+W1ggdkSsAGb140GBMPLXdWXeXwCjbd7qN8fL+YRMipoqBs4GiCqmmwsRsw32
T9lO0OldfPQaQOdehdUE9uE37dw+/cQWYXyO1a1zI+S10+X2YL1qFwu6Z5i4Y4mt
dEjwnwb6TER+xV9X3OzfE2KNG8WRdnMCWVSAZbRqtctihrrCQSuML53N8kbIzoQn
Z+50Wb/+fVfTcksDg0FljL0AjWP54Nj9pZDoCDS5rCPsbryjhXTU8zxRk2ptpFm/
zbulykdgUX4UtYv+GYhO2TBUkvY55OV+xIFFuC/KrArE0PDVQG+uauyUxvARcwbe
WdsuvWBBlaNFrloFhjqiVOJp+KCbdhnS8qqC+ybZ/+r2ahh/JZ2UkOk7+BXA29M6
7xvsNucx7pJ8Yu1QoKfHH88GNSuejnYUHpkM40TiPGWfmtl4K+MoOV1+qTjoNuhb
EbUQv9OVSPYP86bU9gGEgVLNvRAfmLzKKmqKQKroQyh6VybjCaqbOVh6FbW9zVIT
9qCVo9gL/0bekH+jfse8K7flr5PYEiarRoggXszUcSLt0PIG4/wbM2lACxlEYahP
AugHxENyN/GKxBFiAqLWQWSiGM6oqcrAIFE6SsMdkeTWlhi1PnL16FwQZJL94vse
eXMsFgK3lwLfKEDQmmQ4W+oBoHcgLq5ZJtEtj5iV89o3S0TmhrcbzdUvQzHE8cCr
ppWRpecXTRb2gA+7O49qbLUQgiwh2VHgRKpfzTUPmT2qnY4icAD4AcXUm2gHFnyF
AxGzvLf0qOI8A04ZYdV1Ocyb+yIjp4JRvtxhXnm4aKZ/PiWLR7/5TM0LiwkUgZbi
3r+xdQJgcIhcmVkjv2k9vqYoQwIduZcIhZDmPrC/WSfdnrAboYmTIWI4wroE5acY
rAjf/0BYc9txfNa70z1261+vm2oHGXNGPUg1zAFLPNT+ELqesKzYEdgAGjmK2BLW
yevd4BuolfUmjxP/1cJO9upJTHqrhn3rKfDIVdJDccr+rFU7JWzW69wjd3WSh76A
2W+jSiuIJ6+bwnm8Sc4+swvfbF25zGB6OMiZWcIJ95xBO575qP5tugM6IoW0RgQZ
blIYOAzVPiu0CLMuRo9oR1CPrsudugYbJOOop6ujfu51mou+VV/SADSfB8XwGY0a
bTxWpjtQ11jJad47aDxknw0KNee+wavLStnF8e2GfvH6ZfhcoiO7LeooabrS5yev
HGNQKp7+metlWAQ5+x/dvl/g+v8jspP1bcCNB92Qi6b+LH/drnjQATmWJGR2SekF
PfeqErQYtJegkvaUXveNifgnlI6xr2Q+MQ51z4DdfO4+6b1uZEkGioHRflOB9d1E
cJdcjpYJuodIez5NTm4zwPnwXFjT2AABhfGPYlFDNNRdT+lf8WAJf49OlAX+2tlS
LX55q2TGagPS/bL5A4SkKYQYbNfj0Vyb47SLuPEl5BBircwymn+Pi9hMSazhY7y4
/D+YyfNhmYtNMeViIRsbfHjbK7BWkErpLt0ydLeID90l2sDKtEe+1pVxh74JmJf6
hlgGUS3KHIp8cU/lbsypEk56m3Xx1C35o3Q3FXBk572ewEzWxneZ6tmWQm1K6Yrl
UW0e9yTJtoZB2NCyUkGqohNecb4sTBDiDcAhBgD6k2aDy+XV+NWGhLUl7g+PapuM
n57ZVQg2Si0OhiPEyVzIoFRa6c2vby/j3RxXXyBu70e9wtj+JeWW5dfJI4JOmYYV
puc5jKwNUlRkkYI/3fNM1RlK2mFgI3cq3zAlHjug7wuo58eRWnlcuEAFZVTJ06Mf
ZRSvbVLDDv+Ie0GGDIHV16FjqnBb3KfzHzCWA63sKyMHHyy4rFJEecP8xgDIo/Ih
KOz0XgwCgRbYlWzsnwnp6dLPH1p/2dO1HRB44I0XZHleTblpDwwi0QVvsLoRmDHe
6PQUDVRFrVXA0Bj/lgQHiLEcN+kA/f+IXbVEUTDu9cDm6cirYNwazywFhdTu/F0R
MVznyDSiEuv0BO+Vb2WFtaZTnquEThyuxODgMPkqnECZIarVk2cNpo9LcljTsIUK
lotzxTok+BS1inqaUGcy9m2zzEf2je8qF1DDMhvcuaAxPFJtx59zRXeRpzc2fNQl
/CTKEwxL3JHHX1PYiDJCivpX33/0GT8AUZhdEE8RrK/2xZ2ywT9rQnxMJVQAgeFA
96JWNO4Xl6+sanj+B9txnI2gEOEvX4feoOaKp86/1A9+1Tkf5U6TBjuyy6vnzbE6
lqv411FXO3GNYEjyzD8CMLLmM8+km1eeN77FqhGEvjAkq8htbvx/y3675ic4KhnB
xriZRNZ4WUmEhCngJO/ceE2Zicw4RbsqfFZnhOHNP0VYytrZiFMXUTwsh6INLwvW
JQNvVjv4Dxpzunbt2rzp5jRxDCFW1liB2OZBgcG7d/ZFLMe7w6WVB7tB4Cnr7rU+
Q7dRkgKXYqpi1NdNbZVF8ZuJ0Zqdm/RHb1tvqXSORPrMM9hJ770muL8xMO+Mgg1V
h3PZOhvV/hpBZe7MTRcl/6mPN6S1ADa69nhglXZam1ZLc5ADbO51SRk5YzIDHWnT
PfGI6Rf1TAaiO8Q5uzGo/8obp2NY0gobEVSi5ngSTAHpyH4s/yBdeVt0J29od3H7
7B5V6/6JmuSIs8RGiuJlyijxSoXz3fVpj9NnrPEW931sHwxPHcDyhIsOgNMl+whm
7nIAqBkXQDYiV5YXu7Ao30dBkpEA95aab2VyX2cm0GOEV2pHaLNj+ohAfOl1D20t
S2Qobhf0RGhyeQvQ7ibDtvKkCl8b1VHZlQZkvcrD+qXuilEMsL9FlHV+undcEHQA
YcjR1C+fW5AU4HM6L8cyKuc8vBX0ZOIe6lQoUS/94DaMM0xHWJp9i076vLY6/fXc
avMRbfiS5paccqconrNhrq3MIIXHK92Mvy0pVXl7WFj+KNesLxYEfRAMao6sAJUZ
hjcN9ecePrhrtIVUEdtIYRQAbPr+8Cc2GasuRkoUUW6VuCgsKKQEGxw5hAVu2UaB
MHloqGcyqM0GXw/xUK1yle12FjzbMhR0ZVY18yQSQA5mSNY6AAho9tTekxFEqeEU
jZIPlR+nGXPo/b5FK0MVIvIawNL2OiMnXV0WE1gyV2YhJz3IB380ZNgdWhLQpYQO
UQakHmQzIBDcKgy6MAgDQv4okDs7BSuMUaeUWzV5MXB05x+u8FRmrdFE0+2bDnEr
swHfehPRluhkkK7z+ZC29P5GOzdWp7VYOV1WX/Ma5XI4L4rUgWA0xM9B3A+EsTVu
1io+j0sKNAwRxij7xPVs+xGOaYvHqhxOuGXJEeEz9pBqonEwDihciUgfnpKDawE1
5mMpMwMlNKsrKsGdmwctK3Ii/5I5HV8L3eZOx8IvSKn6RdaWz121JTFEqfsbDE4o
N7ttwtg0OuKh30R2dxzGKAov5JHA9SP8YVUmDmiwLLBoUqXY7FIoau868NAgEv24
W9N5jQ4CtzhJXSlErgyDbM27e/MEy9TOtmsulMytLPZsB0QwrSHVDM2iG+DUTVj5
3c5NuZe18DdDLfC/BMXZvayYhzjOCuAAwgNhj48Yzl8QwyEDpUymTkJb2LuCb7YI
p8yDOzcj3Ox+vlX5NbEWNTMEKDLRQEbpElqhbWwDoiEco2CdLVhVfxh+murwfFow
sbzhjrK4YBRSpl/oNvmxH/xq8pi4MjkDW//VKdhdpxiwUAZ6vCoLOrzHrdaA9D2d
g2Fmn0v+p50rHSksbJ3JKyNLh0vHUaukoB0zIfRari6FdU56o+aSvmIUfTB76To2
oFwQ1+Ahjm2SHCl6nC40Oha2cLXQ4JWKfcgp785UQvZaJ3PSOX5OpUPl1AtIVwsN
004xZ56wOVZHMzgf4Wj+ELjM7LHikdGZECUiSf57rUHRfyXA++ieOLD4LpFK/CHU
kCCZGAcGDynaiGc6jTUxOdePaJN9uN7ZJY3c7Gql7OSY+Omwe0KNF4WIxsmlG4+A
2e3L2Lys8ITaTcZ1uSbqGBWF7rN+IklZ7JCRJ7AKZpaO99W71mRxev/RKnJR4XuP
3xHaHQS89bFxe2ilf/f9EdI/rn/hjWAOwhVfBBIHgO4uYkWRr54Edp/HoKiWBP31
xgur/7ql1znUsaEjg28sy1vkzxoyPoXpVBFGTwCsaQy/FHOi13/QD+RV3GiGydIs
mUSwuD1oHXVNztPOUfyrPjgVTMuReFbVjh8rIkVWVWx7hgGLkpjzaP3vNl0YSRrO
000kkXWEoeCeTcrUi8L3PPHuRkHxBLsYTZFpZqsTqq0cQWS0UrebB18sG10C/Nrn
kxwmbV0jt8H5+kM7TTwm66Ui6XwA9nKRgd02xa/Dulb9jGo87hMPafkewLMNwWR0
odcUyq2uEnIi5qp2sNrh2aQ/aBuvCCis+qG0Sxveo6hiGjGpsura65wO90nZbFhb
HOiJhjenxYVBLoR0sT8yt6UKQOl3jCgoEuLdMsP8ESH/w3rt5Y323xFsGXMlX6/5
bNFFvpE86+uF/jWcTQqrxJ29WHW2CgYXRgIxqag9Um0pgLvjChaFbbAyUosW60PA
d1TJxc3PZD1pIP9+EmLw1Fz4R4waTK6WKTTAdQIj5U0a7C8kJwTv6zwACIy06Seg
CA8NwQEzp+P21lZRMuvLjCusiJd7NWMAQeKLqbRqxTEPua+T973ehRQkWJZ3Guqo
0FvbDHjgSIRsF1h9ubdjfhxbmP0eUxSgBuD7Ojd2OaxT/HoauRaiErvGyRw2fAWz
SoZSv24OJ7pbcnYu9744c1giQPtNLYg4J1R0bsPSaMWBikr/Dpw1geelSTooScyp
I/cL2c5DdcZyBkf48E8QMWCwnN5O+AOQTwmHKiDV+ONfBhE1ZwebAE/ucdfCWoRa
OUudCtk3fiJQFeK1/qnu65IVBV6a6YwlrZO1LZMeCleHlLKCwlIbE+/R+cAUjKv0
VU7BV4yLBGO7mHfNGkcCsHjkyhJe1IU7k2Ir0AzQyKayErTTk8vaSkN84OLWHCMv
52jf5LgLKZkU6cYwPxcEd3uLBk50fmRluRqjlCq8HsD8Z6McRtspFmqK187Px0QK
dOsHB4NHT/hJlWlXbovd+p2WJ2Kb7t71vG0N039JHun3X/KWY2UYXIQGs0kpKvTX
sdk4ZAH8ZNACWi8zQ67EXNNs88OJRwi9xuzIWECimNmvxCZP9VBR+Vey9DF99pbS
m3dlg1Mv7DS/9XUu7OsbROSi2nzLC9vfzR+T8PYX4I2gtCMM1hJVkLNI2JiUpndr
O3q0o/M1JCFxudABKhbbdCpl05tT+KffANh37aL9rS+2fykZQc0aaIF7JevhoqGa
m6xDcsimI4emBS/Jfawi7My1uS7Ps6pytu+R392kgQnQ9COGp7gdxOHgS+q3rLNt
Q/pHptNOyuoTQE3M8mcrfcGOKXE+JKJkgPjNbRN43V+yaZdiCHlLmANe9ccJGTkR
lU5cAPQWMXDSgoZH6LAGXi1lveX6+kUJuC987pjqnMy+Yrnr1rbUsFZeoYrYi2RA
ZQxbTcYaOrcK3iqSwrLZd0ig4fnQulVGwuIDkfEx1vd9C/sNk/FmoVPAtqEs2e1l
ardaKY6dIge0fVbr37G6Fb/2nazJN2je8tEi7NGUPtEaoni0evbpzs9Kj+cmemdx
kxaIr9RttzcHuf8BOVv3ZAYKKvRS6z1eJ0dzGQ3ePb52igw2CehMorRbfovKsQ/5
/slUHJRUSfFQXKcT1sLFbGCi90SWpfOoHg5eFzN7XhEXc58aqOGB99thI0kOqRJC
NNiRHFYY20COGxx1+uVTzgU3DFuYhycf9P/oXRGSrurQ9i44qBPTdJStJZdaTz2B
pVIg0URvt205VwhPgPjRXeC5sW/i4lSQlNTBanYTPhOMXn8XECSnkBFLaj5QMN82
5C7ENZNIy77EmcR20TvMV2154I+9H8RNNoBKzpwf2gaimY9D6GUmm5uml30RsTOz
YucC+XXf9eUyeYEIiODVBADSX8N4x4FeQFmTLAQePaeR7bdWezXbK5zSKjdiKy0Z
d61VoThi8FbEsq1ZE1u8CzsdRIUUD5GAUWxu7obYYQyjNr/JgP0pQHDl4r26ChPe
Gb/QvF4w4CH3ac4urBR6mTlqa4gPjcqt7SHiUWV9FQcQIoEs2g4jSrcgpGwMtXqR
DvcLsIqqWfhGHwbkC3V+x9ED6ZfbTqrPEPABy6xu2+D7hR34eiKz6RcrLCM16uap
ZN83iR4O9m5mG89x9uZWLfCtnE8vjFFVhdGrWJGcmub09XcWbDjhWhkEFRYRI5YX
k7O0IH6yqDWlDT0p1flXY1v+V+VPRH/yFPN1tU2GvA9TcMnXUapj9pKLGNP202+R
Q6odRD4nQ2bdoODcL733CRiC6Hdz6XRk7ykhUUa60l7gEFtMxVzPIQrNEboTQakT
kEQ692egAf7vu/ToXw5Tfn/RzvoqMcoXuQ42q9kJod8Rqnr0O6UqFeM3MFdeWz45
B0VaHOuSEGSja6oqlU1F1lOqO6dyOcoSb5W8OLTUmA33juvOvgcAggPiU76OrQ3R
vuMGmeN2oyqTSBdfdZiBhYGicphhBudo7mewa6XDk9y1RQSUYkdPE9Kl+ZP3mtG6
vcPkVElqa0vRQIo+edAULJApXBqzyaTvjHA7X1VdiT0h5dN/laiZV8tXQfF+5N/L
TeoG/KO3PTkds0h+IAy/74ZA+7zJC+SpTRJGFMJDLcTSQ/hZspz0g9gPc91YT9Mh
8smkpsEUQ7DshQiJCaMEpF3hfzRjTdDKtgO9dEPz0SHeFXpQZ6XZtga7uBz1G0tJ
sIpPPklaR5BOGrdo16/MX+U8BEnHQNTaoXbASHTF9FIgjvhw0oPkCCwGyOo8P4qp
1aIuvjuNQ60dmDuH2QM35vzQGxwY+TbY/pagSlu/fGmCDLDpmxAb/SrTODmC9YB4
//m5yhmosPe9JOgF3bfMyayc+GCkWXvt43/2ZunZaqIjWWlANOf8HLZSzRCpBQYa
jMnt465CiUcX50n03EQSOtUrJw+FO/BPic03Dt71m/EWuSgJ5/oI7YiGJHfGWpn1
wCnQHwidWTrOT6drWQEh2ZuujsrmfLv2CAFtBtFOKEPyNp4rQ3k7aGPyGxtDkvrW
2bDQxna1QBGjb8kZxLbrdMTCRjlZS5ePJMlp3nTSeXQyL2SkEELTto+sTInrdiRA
wGs7JT/8yANwkXMQRsrqUj6BEMcVZg5fmEYhtnLjYKG3aN6xni1+40G/NUl+DB8C
uAMUpTBwLOYE8YwO9kygkR7yasUabeWFlRMkuJYDFAz4iok0/d6gWwZOuRCEv2TQ
XLgZ/BIUAVzrqt3OLHAaUkEGWfph4GiAgvouPVTlGWW9q27iTfxL6pni3h9YdxzN
z2ZOC3fiVp8Ov20ULZV2QUEHq21S+93OmcLOXzTQeCGp2Q4oU3zdv+PdhVWxYrWs
byk8O1Lg0a3RfGiDvx6Bu/BGfg6j7xEAnTO8zhDK3EvKjbc0mTmJ8gs41CYpm/7g
WuHZBeS2feoXJOphq2BRno2WS0ExE/56qNxul3sqT0fEUVVihWfmUdiow7DDyJsP
uJMSmD5S56/P4HfMtf4cJOmdgShSW0kSuA/Nc7A3f2g128dQIFlrS3PbsscTTcGS
nUnbgi355CTkBWAkr6xRyCQJREoFmX6nSWKI40yiujywQhXQBL4rImjaAuszO5em
EPnkV3yuBW3UZqPhWixHYqv3s1Yem4T4xEr9btTyD5VczvuvywFgEVx0Cu16Ybdk
cF6nAZLgIHf5OIV2AKclGzWfF76cNrmIs1Jo8LLH51xNglRZ2kBk1sgpjgD0gD8x
UUhXkrAUXd5UJcEVaI83F66AOXrXvLiXUKCNNmxnkTKswOwEYG1I1Urwcv3xr/si
CCokF16DGQ/xwYIOhI5ZsT/qTPMcZw6NAFA/7wZda2w3OQu/+M7xziA8N6nQr/UM
EH+YeQyUkVsI+M88OmLco3Tt+o0D9rUW0rkE/IFgEmm93wn8JBLtR0prY6VoJ4eF
MPCfsMG0TiKO24zcfr/u+V+hC7M43h4nTdtmtDjIjXz7L+Moz4jjdiuXwbJ3EBUm
5sYNrdhou00c+lSrMV41esOQBHHQp6MCF/x2ceES9+lHlGIx22l/JZhDniMvT0Uw
FMJm/KWEDzmdDZrlT0PNAruRYj7098DiXzbgMPZGTjKqTFcHzJgkx1tt4A4sZ3Ay
IQiCBzEJSAh/9nAZVMdPTy6N8H5VEVEi+eGKPy/rpWl79fYIIQXWL7iXMzIBEFVQ
VqCz8owp9ltKKDzLPAFxNmvwUGHedr3kU9pK/zjNg+qxXbdgKBmY2y4fe94e5J5p
qfiasUnStiUQtxiDaJTBUk9aZXLd58do4r0dwWadulgDTTyJmzmQCHF/BNOjauzx
KRj/HXsT9NHL6kZ2n2Kx6FWG5bIjEY7glWQQRbJfPMoUbsvSwAFIzcikIP3hiKnp
qEetO6hctKkxyK9PRW4zLxhyacP8TuuWnl+bMmJgCldK+AToJwPxaMyvbiGjazyc
shDxwFonbELNRGjFw79FUwCwn/iSjnPS90DbJs8xHz5oHkK1qPGqnag1yfJDJ5c8
rlRbiGgGs+0+achhApN7nEXoZWDJHe9gmabglWHmCCCq1sH3tsyriI8G23rn5oxj
sgF38ub969z8xqjZllhC2DLl+Y+5XWmx1Jl/4CA9flQkZYJeBpUE6R/9zJxJ6CVt
VdiqOc1n687i/H5HFyY8GTjO93v2Z2cbUaK2C76MBTnxhU5Z3HTOeEICKdAhh4Yt
P2hwi3hysq8NTQgPsnJfNaAXIrsRIt+0DMQroPVNrhBtbOcGTfjsuO8gMlmI+8ro
qyiRQamfy/sTzF4TTUJ8HeFjuzT7WX25GfDbpUlgAJbvZMbUy7dbJV7Kzi/lONTC
Mw8bZXnAr4Zyx/f1FT4OYoGknm71gyv+FTE/rhxjb7jOOC+z6e1ElsvdXRsusjxk
VVx0S143TDdRuntT9NJb12g1rG7wxBydWHdjtW3CvSbyfGf9Mj5Nz7LU9hObtnc9
GggIX59Z1A6vjje7IOIf4L3dDL2eBRPqdglWnZXkhX63HFBkJZ6dFUYNH7m9bc7t
2WlI+jj6eH7Rc9E9xweWOzps1s8Mo6pzXu2VAF265FRMitbBD7EHOfMcEOuYtaFQ
Rk7b0HiZLKv105Kg/eaR61L4T8OSPBvgF3VBumT7pqmzQ7aGM02PNetv8csPJo2h
3JhVhUQjpyNZ2X/S4S6f66Nunojq/6kTR0ut1D0w8IwxbQGoQuTf1iEmFf+QwY4B
Pup1B8dSUQkMJZBuz4SRILqLuFOHJnvirI1Da4kAu5paIR/qKKyCUFjk7n29WkCW
yUKl6GLzG/ukbzm5OaevZyrBlSeSVVWcMcDpogJt8fohhBvQ0YhOcZji9OE+gY6b
qqgZ44jA/dDDRZkeSWCNhaERqUwUiZj2H7JdikrHuKyqqo2SeIRbxJHRInuIC1bk
+mGM4jpwjAtt5yvxcZtEfwl0Q/4rqP+3ErWc14SxU1706fa0/HlWhsiaMS/QQoWu
chZGeIzr9G2/INgxrsRYWtbaTDe2LvuUTfpNA7DH+838hp/iSoK8ku2SsKVQ4iPt
29uM8ubNoO85gamO9ebAjSJFm/dEtOMB9ZQZYgE53zSWm+EhYY8OUbWDNlSni3kI
sZ9vTgeg8WoYP3NeDmyK0xZgfx9qe6sEfUqfyMtNyC67nqYdkHovcWASuFTL79Yc
R/4PCMvlvWEr69TgNLIW1TmLyYcL6aPKGEg9lge8sytjNqVg0J+7RbRehJIyv0he
wgJopDWqO/CzMPzLULqRpK+7ZCcVSPj2ijwcLoEP6aad/i2A3XiSHBb1GtAALtHx
Idf15IxDCr6j0xAJfHSflT57YVv+CbvjMmx4JXJd/rqj6f02p8rR/PQloLhq6Ix1
OmEiyjIRJFveS2JJgRQPyd8E1XTv1IWJQauSJaW3nzYof3wexeXZAMLX0teR8VsF
0y7KhrkJlxQg+DZEB9+7Ktj+74/9H7zeHeMBdP4y0GVSd6/SEYn1/FqZIRMRNxW6
f9nYBmFbAWhwZorjuLsgZzz3OjnTNNTRBje3VLocjcftE53Y2TQswD5mfh7sOKT8
nlSLOOYzc3l2vKOLY3+tuI9dLPeKOgDdB0R6/U62/9unZb6wfJZ5amEMQg0Wp7Ny
Wylfxr4j+oUCtTQKTxYvIlFb/qnctAn4bViPBybppJwM+VHRQ9giXz02/UTT+ynm
SFpEPKmp+uN5eQJhFvNz6HX9FHuFGIZtjtOZP8ixPrwz7othIcE1LPCScdINhvU3
UVa7etMztqefox67XQuKAcq4VYfBDVDcWmpb8rU1Wk4JB96vxFOP0kZb5i1yRarV
8vw7kRZBdUZiup06SdEp7G59IbJm/7ol2iqQiobrkZ63tz0IPg+WTFNh0qPAaOmf
5/p6UocuZkutoYAqW68B7ebcnp+1zNHtMiiI74wWrJfHZlFqX0lzwN9adK189aYE
B+b8mE+ZVQBecwmVkhK9NqPA/1SLEC7s1/FWrqOLeeqC0+7fXHhunzqiwNhQhkQq
RgjlyZ03pe6ctY0xi0uyCwbyqqO9l6orud2sO7CbxHy9RkfPpCQogRgd2aALr7wO
gD3DDrAY/+DKluDQ9zE0zj1ieUIWmYbLf4ouRF9ope9H5S1tpFY6Bs0nL8DVj6Vn
Cp3Yy1yUPrsQ0QMMe5QDtunOLJkw9CMxMgNbPY7xmfsuKM5TspvNopJBQJEHuvGv
nX0KBncP2ZzBzaPy13sEoxqC6cHrOTesmtiP8tnAtUyxPSbtaEPERfmtE5taGayV
OQPEJR6M9Nd1vYSd8TKDK796Ao2Z0aAy7jR/rvbZr+9ScT1F+AQgYN142Xo7yAim
xNfChVFd2c8KxRpikw5zl216wNs5lSX6+KIW9DoHxES/34y6sPOp9qcUnAjuRHwN
BR2aUTD4TEnRdtkSKSI/VZQ3QyvyF3AQShV3wDAt58utXyf8aZxqOf0JuhoL8YvU
iDkX5TUQo+A4SDo/rkzJdnPq0Uao4sJ5cREsw8Q3JD754S/xtXkqEeb1zl6rp8Ga
sr5J5tsbfrG7L9ykFlInvBJDIFmnKxjscJT4/LHvEYVJLyDMpMdTbs8chu2dJeU4
VP7D2QCe0EpVz9S1PU0ZD37Rh8dCUpmMbyU3iLsu32r3K3BdtjDkuNB38l8p4O/1
T9ulOQaroUbb9MOQkyE4sbz1u5ECWVKk1JvAdws7dUly29xJ2+nXB9Ta4zo6S0CU
1hzU5DlH5n16OYwcHVHy3n7q8soj22Td1z0pfqIQU8D/M9eVTQZr2QR7PX1U1bcF
dGk4S/C/BZyMHvEvrUu1K+6ibDmHS0BlUNisMB/0Yba+mvX0ylir1d6dvwA8teA6
OIaFT+Z7a8EZCg5szZwSjnRXg2Zc8LFtOa8TOAbmy5aTbB9RmcevgbCtTQ4C73Tp
57scBPSis+Bbvld5Cad0/FwnAn00v8vQdqItFCJYpxMxc0z+O/6UHndKFzB+eZeT
3frbevy0rgzzhPyq6cS2lVdd9If0dcyYR528GvClaJiW7oPEny74dSQFiN5TkPUu
xR/K5o/vh4hxxXBbbGm/RkwAFCgO8Ax0TSpa9BxFZnshLs7RadNCKNnC+BLxko+m
2zuPRIrLRncy0n4ohlg3avsp95H5Z4EGPZdHa1Zt460EALN9VKw9zkh0qIrQglHo
CalUHWlazEGT17mdRGE1gEZ5RCDNdVVSG3/x27OyfOZlg6ece3w7p2P4j3K62VuQ
2OsAgJ7kAGZO//C5qHGMWbKIpSNC8KbL9FcxlKoV0UDsjC5ngPqXjBYb3bfm9t3/
mnAsboWWhclLJeQEoa6gk0YAQOU36F6G0nv6jzCpGsEJpyb9a5Xz4bGNob6LA7fO
2gcfRXizzonbGZa/qCZLFenrhbNZcqobbaXCo1J85vpndRP2v/oxVhREsWbo9OhR
qs1Sa44wrtkj7ZwztsumFS6WG8/ABhGPVB4CZ2WoGYvKVkaZvMd2Add8xlcQng7H
jhD44AWFTiXRnCaYMPrxXopUdgGWWNLBt4bssYOx6hr7BDy9SG2tyUaGDKWxN9KS
nLIVxHNRmzmqVvBzqo8tSjXKU9pHjxKSZshM5udy0RYKfS+Dt1xv5Xs62iOzF0LV
MyZkDBlnwpCg0iwQ5KQhd/YDnhVCrbghWt6VkAVn3vsmMh18DACy8LKbdLnxwJVI
4TO2AtbmqlxyhLIHQrh6jGfsdP2qXaASivkIMPejPHu/4hc0MfRUutBqXr6ETV3g
TJImohdbi6RrKMX/LfFN9w4PlEFuYANAo3MXrJDJcniNgY12E/CmHjo31hgqSrPu
/QcWi2NGJ3u2ivH4+mrY9NdxTKELX/W+TZZgzJDyz5TRBKtRntDm39SYvcJ8Aawr
7inDJtRgFSHr394uYOz6UfSV0PsLYH98fd44ii4i567WdZ272GAX/5mW8LaIFGfQ
GVSSR3lZg7TuxEgF8t8/7B94AFcKnL9Huc317zT0cAk8+ES1BS3caW1tVowZQqzs
IJZlh/iyvUZ+MbYKIBr2qeze5xWlFSNslFPgNOFbB7JJBp2/BQqAPNonLByz6w+n
yVZxXAWgUFJ0w6p/8NrJ1s5R57HKyqc/kqQYmdIFYVWKd93JocAye+nHWDZHeOWn
9QIVE3zz3KBXAaRJVdgHy2nXOXOIvHle76p+v+wXUWDfkcP2kEADKSbmsocp5kIP
BUHcYoJCfJBoipRfRiwVZjS329h+EaFCr6caetOCp+dlL7fxcvv89Et6w0YFJ8zO
XVx5qtZaoBm0/1vFuroQ8sSIeAUNKGyH5l6u46E6cCrQAe1hYeEg3X02CJoEamMV
r0fOSRQLWAcn4vrWDnnBrtV/5mjIbguTzDsawUfhutU5tmccDul+ADkTWnTLPOfr
UzNe1EQHAwxbHC/CD/U2LtAhwc0wm6MA/RKAgewsu6YoHCrLsXJqXp+nq4PeDbOL
mmYndH1OemGl+8FAtiK7thKxAAj/x36zRYgocFyobewp2Bl0fjdHx36JSs3U/3kU
IhNtwX6rFzkDvr/xZrSu9hGFLnOY+U8P3RxrqgXU77Ets5mXjSKwIQYuG+MiQkLL
aVztQJqdO+g2y+E7thPuYUA2GI0ka6YUav+vq2ZL2ij8m7e2YshTP0pA33jjABnK
sOc+cxds0pY1t0my+ClJRPcXOmsy/XEOWG88tarn9RKPqm4ZPxhPZOKS4B24WdSE
UKA28MG1CqAldFV9dPIIH8BYVoS/Uq+uA2txWn1gLZ1R8VxXP/Zoq8p25Yw/GXNk
WgS7cfKG9fYrLOnyH8PSQ5xON/D+c7v58nbDVV9EvJ0VXNVnT8rmt3ErfIyZ3ycj
aEcMgOv9jrRWXNfYqBGo1HyBmeQaj9orxxT5zS8DdvvzdMsA0hPGAP5XVMAdBXrg
lE9/uvfSXha9ZVdJnMXzlfW3hjIq6pa1HqG20WLpAJbMmBzqURQj4qHU3nuD/MFF
jf2tERg4OaGTNAD2ddy5KfVNCIg9bPXbspDSM5hIIg2eezFDnnTysV/KkuE5g1um
Xvl+8qMV06CqhHBY69Y2IrKBgbSCp0XbciR/TOhBI6Y9rxwtuYji5i2SQBI6QQsq
AqoOdiJWPTWo23v5ESPRM/kL/xqhIUcufIKphCU+O3PEdMo60C0j2/SbZxkb987c
H2h4tMykmP+GSbZdjwhcL3ZM/zJwEVyOd2XaMYL9NsVSoPi6vpVx++CMXjPjzrez
7aBySgvsecsQyTfqGZve4kIxFv9yN8pJZuVkhBmQ2Yyabvkf1GrON/PBMuN4U9Ft
5w0xjNhfrzwenmXTN9N+z0T8wpVBhEzGy2fqNirP3pBr1hGZORsirWxwy+YzEbX1
UFLgw1vBfEo6AZZ5pleh5J/E6Zp3dCmZFq/A67rUnxcGziv/WOEDTdKt/VfPGpfZ
pXbVDSfdJvdlNr5Q9xFwz8bWnf2DjG1zvz17gcpGMk6DjIMdPxp+a3QbuvH40B4s
SDmb++aoUteCdNtJua0oaFLAEk+zgsWIi+7RNz5JcQwsfdKWbyKP2xaHA4xwaQzk
t4FhgV6P/3Ut5MWmBjjhbRNnX+0aX3D0TkMH+yT6gsipuT5b1XzogInbdrcPEPFc
5VZ8TBATiw9zVJIhQTWBS9+SgWpdsTO9U60dTIN3uUQn4gOh281ewJZ3GpAAxi3r
k1JYArLoUKgzkQwHvZV6UJN4fAD+xhOJtFlgD7jg/ETXOX69Y/LfHHgX/Mcuvkn5
jfJ8CGXkNy4l4oTz6X14WOLlu5h2R9Q5UeIM98pn94s8jX/2lqJ8mmUvo4pmdTJO
3xqXeZ+JXN22nRT/7/f7v4D5lBHU44f2dxMdeEKHUJPeVOwze+vm/ySlUWrabqlq
TGtMyOQSPlGRVzAZnPqLvGsRk0LaYyLE9xel8xGFuSodPaoiK5m5E4Bmre7MN0Ni
fkQZFFCqJ7YXCcFHylQTRVhG5+r4/ZOAUQjNjuUzFvG/4896mmzQ/857FLu/hG3x
yWbDBbrPko+KH2VbFmDk6HrxfUcSqRMa2olSrdtHtyFilBsK5wl0LGo2HiiRBef+
l6VGaKWBJrnXpU2pixg7PT7V5MQqE50/FWxpID5O+HWtUQlAgYJPXOowqsfzyP7q
OGDOUe1MrfFKVt95AmRFJOOM9zIrBkXtnO+cm84c1ECn42/ZBDYUWqfcxtpe1TpJ
XbOw8SLiqmZvKemuEsA5tgrGWfwfLSDajkaM9Rw3rkS/WgprsezZWrFNZ1wPUZbd
6A7NO0VTkwAWyk2A2l2wEZCRoaxceoKcG44ty4bu/iIAPs2OUVVPGev5zv4FEnX9
oMajYpNfumPtyM+HqUQoHbeZfs68PkN0usFnMe+7ofHCTw5+8mYAYJ+IHkxiC7nj
3YJzc50wBve7uCA/rztLuXletXJt2Sty0rx4OUWz/gk/jYlc25WNUkqm2GGkg1Mq
ewEOlX0/vKeo+R4FWhj6e6ogWFqFU0eGnMjCCEUE1FiAfzU/gMZloBs1df/lAiHD
iKUm+QJUTLQH+FXEdAl2q4JhnPlZeF2/Kxy75ySbQj/AlTrmVCJHz5/SRi2QsX/u
k6y1LWVNAUc9CiI1ugPrbkPVKdu3pITX11PYIryuOBlzlb9aG4IbAFQFm+e00YmU
YUp9HdGKD/4fJoaYe5dpBUVKyq0WOJGyR/9Zu+BiEvEHX/XEDAa17FOOokRo+nQT
k0a8RmDNAau3TNJG9cQdJb+E4aDw/7Ex6vNXIb6dpKqTUpVKh4xEVQKDqoC9Wjpg
WpcbfwW3IOZUZAavLqDNqCO7JDzROADIzA9cYxjMv0nmK+dPyPjFkWhPQMLoppbV
AW3i/hQ2D8aDaCOZ9X89somLDyziwWvAUFE/oGvMStMQVO3BoOvPAWIfFv5jtX8u
iwehHQW3BlHac2zsd7C8p7gRBT83SzFgI49XYBc9ZWDzNG4kdf/OxC8zv1h8qD+z
4nyt5+S4FjMVW1y9JCRpvcq6RzAmqqPmkXbci9VLwA+5ij7EA4P3410mi2N6zbaI
lvp492tNj2CLP7wsMpW67f4U5PhplvQb9ugkxRXQEofvAXxo7Ml4aZg7Utrcl79N
HZqic/e0+edPONcavOaxB4SN0+8EdhORTIAo7+BqQsgie0GNO+9aLBa7gE+gpOgn
hIvQqJhpxuPHbHM53v/jp6PZSOPj74CiAPh669PqbnGmyt1v2eunmQPLRJpxzbvu
EoedYzMNcTykzhdV1Z0AQmGyC75QiLnM83EGVn+O6c2d8ibKfHeZD3jsSwbjLJzW
zOxTp5Uyc5aeNUNLpsazoqAjSrroCPdepdZfhmHwDJvYQPJaVG+yQXAer2Mfa+g0
2DO9/tiTcahVmiNb2aPduu3+4CsAVwFEMPUQqnLzMGDidvMvZJIeFpbeZY70acWu
MWowzvYqN1+j24hNJrNATVEAaO+4jvW1R7ObLo10FQaHcHHI1pwKZtEwmDtrgw5a
cVTZ5UoVeex/FqJRXzZZ3yP0AZw1vAW0p5VRnFH8UO0gZSM0dxHsjEECon6qIVsu
Tc6AnSsvFtSSyI3o8KOTPCWuO2mdaY9k4nXpGcHRVRGd74rDABqqU3Wpia4pU6Tk
R+KmlZiKFVXqbkKlNUAFiV/FtTTO2bvWxAydONDzkUU27qNbrEVdZ8fdsIJmwbZ8
Ha0rOvbHcZc0vKal5svjKKmgxvbN4YTSZj8RTUIxpNOCMNch+Mea72ls6fy4/rxp
LXpLS5u11S+TNvoHZhOHlw+hAgVs32BQH+NiE49STcxyxzy2SqFeN6pUyF2dFgKb
693izKPDM7/FaBHIbWnwlCHILrnK28wphAxlXEzQrOY05pib2+xHSiCMCDT6IWpD
BpDBFuo8OPTnS97ueTkjprcYkwvP93t+7XXVtIpjCG0LN/iDXQjx6iIE1MunpElU
llHqKDHWO5Ti6HAO7Wf3r8R++maw0qR2IyfMUQtxXv5qbpwa8vqmbBBT7GbIw+yq
oMHibCEYbfiluiT1jTxsHvzrSfaHCDIw7XY//ryK2lP3lByrEWSAdqHRVeQLqPRS
wbb7TJEhS2LQ+nZ97UKa7WRv6VbX+0VJXfytyyFY2JSUszS7dZjOFtM3by2jKKc5
/b3c5S3x8Udoyj4RNj+eDzbP0ZGgqQGEVoMPuorUygerrM2rtAxU9BOkFIai/vuz
p/2pfdb7VlTVkcHBxGJbiPTDPdZNUKNqE23UBbzkETrpV2hbwn20U3WgXxtRQIjr
l0HrSh79Av5AxflKYyB2HnP8QF0H7VVurKQ9MvSJhyU6CrhyP5w/GVtyiqEkE/+6
K2PUekSsdYj3S2SoD2VVNK+HCpWqChGPNKZfX46kqf3MSiBUGWKe/yIrycl69kMX
27q+S7KiQ7Zp6y7Pu4Z3BgZfQpUb7V6g/dAvTCKX22VigNh8eZkMYFnSg04zf2P9
5tmbSwKIXU3NTMKRhVdxbrOmMz8Y7m3O7HYaZnX89qMQim8rdd/4zqgLRAsZXyc8
sZhpUlMhuqLXwJ007W5E1TeG/2I77BZDsMGKKnCvGCMkX/RAK8Q4UbQpIB6A/ieX
bRcw+0Bmz4qt3KgF0y6/QelkuqAyP0118jxjWgPUu4t+V7IM4gvQxxNN0xErhn4C
P+L933/CFkn/GxdTss0YQbfFISEUU7XLIOA6rrpbO5ARXjXukYKrrvIOqq2p9Xb4
+A+cMLcFH3p/tKcj4qs7nX8zWVjmrMkfxQLMZ9AE+Fbqcma0TJg+xjgMxZSMT5ec
Qvs0Bi7xqfqXf73UssdxCgjER5Gs3g3sdbKZ34sVuxbcE8JlCFzXeEPqipaE+GRa
RoSs8aULuxKxBzNoQHz4L078dlzQ44v3LG6DsJ0yH91sTfgPDQlZ//PPsfqjkhF0
RMWW/T23A12UtQNZoA86nlbHy35w4iaK/B9Rku5Ty6wlNy9XSIjiFW61iU0p7eKf
oV9c2Xj+oK202+HnWVkaa4JVfJ3g5WuCPSEEkDvLLhe14eg/9HdCY5IB9YyKNfQb
X7/75t5z83npVfog3yfTeDDjvNSrt0wextSKT9fQhVgfw5vhGsR0uVCI5e83JCxI
OFC12XOv8g2uvs5sUEdjPxF9tZmtaqacpcTkKnlXTpWy/BmSNdloSP7lnmwsy9WA
zw+3dHgUKWaootPJZrDCfowIEzSXr06Y0JdZPi4jh2ZjVW1gVBFo92LjUFr12hC7
s7dq3hGP49lTTYhBS3Snggw2bWaydXpo+WptkzDTWlyiuoidXyswDjy4yTYctUDp
3mpLxA3VwAMZHGfs08fVWoT2qADKDuT9bctU0EfszjV9DT+KQ24X2ETLrK8Xg7Z9
M22+h87J1djktn2mhozBuX5fGzz7KNYHrEIfJN99f7w1pw/hGUkMVoLMSH4CwL5h
N5fWg6saRYPjq7q8TEobyVejLcsq+IQxaeHFnsXER+712GydPiLMRqzcQx9fPQuo
BcLKfW/7YBVfScyiohWiD/YljUPag9zUuT4Zq7gWpY4ObYr1cQWkBacXQzEUT7q3
6R6SFRnj6Wq5Ff94h6V+7jB7fitobucUIjZh9eAA2pXYv/lbh8REMAutcdqfroJQ
eQhUrZPg7SOz4MWYE6wh6AAtv6STbXX8XZri+7YXxwx3HMPbisywtUOhjCRkcWfG
+O3ZQNuOdVLw0dd3dykoORCDhz63B9W3MNMPkNa8A9Z3w9HPP5/GFJSR/AXdkry/
nhX5+oOw6jlRBFu+5SJ0XjTKD2JbzZ9iSkp3nQK6A5XuMTwovI739gZHX8g2mrii
Pc5E6cqLrzEfuQlzJ03Qz/DhWSdmt6kF+EOEWMEz+lITtY8HAcyVWG1inrsWuk5m
SJSwoQr11ctdU+a9JTBXFqC3cYLNtEf2uU+YcbSram7qQPJJagftkmRUG8kKvCrt
/xdXDN0L1QkhfOMMO6fNYdSOobjYZsDlSyZwRimJYN/QoUAf9SiJzzKFlO87Whsr
ROtBNBgwzkzA84ws72TK3GpMSmaMnDnIr/ybp0NfDhJkfTtN+0pjTbrTPltSleeA
HJeMEtfwk1QOKuvyXpVRziaiyxNQjlBkL42KjI2I5qIYikm0+9k3sYq06ii8bLr7
4cUJcm5qHnYD7vdlSuxPvRMnFdpnzXW1jDMwZet2pzkBfv3PNvJUcYJ9amPwbp1/
hl5Ptzee6fYv0scvrs/xWcjqmSo8SqTLdYFchck3ssZ25xrPJCi/9HlPp4QkQPmi
AutUuSZw4YCvjHdtNbHoVGAe7A9GizH6GIXCA4esCUO4M5vo0HKsp4S5fwJrbNYp
BxcSDHAzNi7m8niJmi+Dxsu2FScoh6v9kEW3sIyQMTYmWiBCGhSey7UvSDdzPRUs
H2aHGnBtPg9ed7KgVZkqy4LqiDbKnPKWtswrRoz5XDAZGO9fjHIrj5SDQ0rmf55H
h7ke2CzE1X7AFMswsG1UoNt2bUfeKipR4muwOsXr2Ga34ZvqIW9mfqBHJplcfUx2
D1xsiJGJcC7KyQ6WBflLHgPzFNyozGhfYQ16cl50MXKHj3G6qMBA2pztn/X5nB1+
IB+vIyOAWdB0By7LZwhQXaaXXlyaLGrWoAgPhE7EzyuQeK2WAYDkNZC2FMDiq8Iw
ztuld4vRwW/Z9jRcKND3wTjLqntY/2OUKLiIa5dKh/45UciNYC6yWyKCwhWAyVbH
uP7onbNPeVeaZGMTdWFBGvtpf/bUDTkkIOY1aj6wVJMRAthcEuODAJJNlATpgcHL
/mM5vh76mwwQEltPNDX6+o9NfBU5YWV15L1b8MdwguzqyFm0dd20kPNu9HePr/Vb
N/3QQmxhGWH2xfJIy55l7mF7mGV+X3GWMC+I7NwXgQwDBq1D4ViTKNGVwdXKHQY6
iOepJWoTs6RrxBubqDIQ5a78c4+ctp6Zdgq0DP4Kt3iNHUruLsshuzhgidN8hpea
R/RQxjSawra+LKk7hxUfojyo6VVdK1Il7YjGFlLwUImFOx8O8YE+um5EuU5IP7OZ
VIWXU8OguSgx/CdW21TTvCGizXN31BSWPZDt9NfU/5MWxA1dIWGkFPBz6XNXNm0i
6AWpcn7bBulnrWpq2pz5C7kCFAd8ROcal6sYHfI4wAVPN9su+Rroqnj4wc7bujJg
/rHXsFGW/pudMfhyRDnccXQwOaD6b+W7qrn1W/clTSLSjLyOk9bEwNaj7T2X9JmZ
BDBQogMvv0esiaPsivI4Yco39o64h2OyR4CRUu/t3Un76UdnqUo1QrvhD3WEFEQT
x0fP/ttzy5vJUt6Jbzyn6HThlzHybhn/BwG8EnQkrexx2pxfBPT0xpmiie7y3VlU
bedLz1d3OkPBxmC8hHId1wQyms18BeQn70iAmk+ntUac0DCbofg1hzLxdXBrug0T
34IT8WfRIjnJRQKQzi5naV51fxgSuUddqq0Z6b+2VhAWwvycz+imSXbS1GIXiP20
L3KyjRCAtZ8N8Plt5GKcwj27sSFc3OM8+Uyer8fIqKtXkOhmWAQnRKfwTRWIsS/B
6oPwYCwb9lsJ42BuMF0MKy3+9AsqO9jcckMM7SKE+2eSpfa4gVyGfiJBpvGaBkFn
LU+dQ8UhXq5MWEM8y0vl5ZJxJF6+KIV+Mc5+2T1q92EMPuNOSfeXCck5MdwgwZRC
8IsgtQL4pYdEZKrPPcGisXQ1UFPVB0y/Qdsf7gZf4reFJJZ4LMK7dK7SXDOBPzGm
ji+ZoX3Y/M2tPJJmU9+et7oNVP/4PIQEGlYklU0Y+/cPSYopXZSZD+MnVuNoU7Rv
8lrVT+FKikfwj0qETq5YwBiEMirHd/ljpLnZ5FOiQPpqfqGGCI07yvN5lpjye+lh
I+OwT7OTjRvNYwwzx6dmNRmZlGYq+/IE/YCItEi64QwBqTbMTRw7tqbAXv9OrcvI
i/1Vn6ugJFqK3kaJI4qbXR2ojaqBUN8M5F2oQp5ssh+XZJSbaCzPuHNlR2JGu9lH
0zp81nnpXTSMHQJxREH3qsvNG94jfeNLV9EyepJezHtE2dhcjc8vJQSw99RZCg3i
VGpsOPTtS98G1Fr/lGB6wytux10dQNv6AlqwH/p/aA/Jgt+fc6q3qT0fIXudkWv+
wBw/tzxzmopI08T3klCL544uiWnmR7qSpIiOIsltnXp5+v3blMruYsV/WOZXGcCW
piX12DN4acUxjhkzUQq2eu48/ObMTGl30KfZnUIlbF4ohbKTl4mKiyfWOWNTNI3W
N1PvnQNQCoGqHONaVoHIm6PjyvMKhhBcildy5UAF8KNa5RvWi5Rf+xqQdMbMhzXY
Z2MFrPPVaqRRkO4QHbfrbm1AxS28cYpKXRKwQ6iN/VPF1WRzeUO2w+B9Ty/KgFu6
Yedwe9Mpsq0J/+Z1U/emrkBz6+qcFKxPinDkZ4wyD4cW/TMYfQxdFBfZ2NkH3UIt
ZetLRy1j59RnGwn8d5Q3I2+NhKJlNWtB0Mln6jPh+Yq45FHYLUkKEEh5L2WoZj25
6OJIK1OqkByHtbh3bvPn3vTBTaXYpHUgmqq/ik6j2SL4FFv446mLu3ENBvobZEyw
/yQURSPFaASg9+7yF/kRalplbxquOvZi/3wkg2N5xgEqNRW+tgkyYFlqAodyZejW
TfQnlVY1C92rXAhK72k8PZxYabURrWFj0T6QQfyzeyilHygCPyZT5TorvMnNUFap
Ey2WZy3I3I77NuFJAQLzDFy2z3FipfK7AaohYlcKUA7reQQGsE77cE6XhHtB90xf
vmmUM+Hig3Jo6d30Ei55TMlzelREM65q26N2cYIElpulfkT4e63BLg9pwLgyidKr
Q71OT7ynUdY9lEUuCu4UlfuOrghWexs7DnS+mVhyB78wn6j4EsVSQK8Qtv0bS9HC
kp/nMTwxAGBVsHPI5xewhFTwxhREobcrOQuBi2H3roFqxZSwLhqCcQEjUkzU5N2/
WTuZD42s5hPV19sClRQKOBTQmkZcMEgn5QigEjIJZ4B+qE54znT1pw3pYU5Whz4k
AlMjsaheg1EePY1K6THh33USJM2Fh/gR+yALxPlcX1qzE2L7E/v/fJdvwHUJb0JR
yLOV7gsfUJhRuqInoEvgrSnW4FvkIF1GjCztYSdZeZY0I5K/x5RzYLwaJ0XogUTR
Mp4hhskw7Cg2McwZfNMwGD16dvND84oLRHdP6NlWh740jEfmxMjCiAzNrk5f3Vql
69eiN8tvkZU8ClKIKMcBTiQIIY/tqZl+k5rNnHupRS002Veu7Q9InwSkENSbQDxJ
w6TdKO/HVBbCJkBN/8HpaJEyFF0SjM6fK6H/jmdNlNJoJD/cGo2Q4qIzdcqMOGM2
FK4gh4qOPALiLxR2rV7jwv9JYdxAORVzEYZ1mb/8ttAZ4LvxH8ZRurhoe01PbTn2
lm0tO0qJj69UsJaTzEFWRRJp5Gf5UulZkz0ahQZuMFRzUH9nvlArQpQI0EumX17Y
7c3baDe+wk5CQ0cYhI9+lK8DLf9X+3byDWTvl9GaIBVvSZs8Wm2YKNU+FrO/Nu7/
efjA1KAcuSkRUKJKtIXBm3BiBdo5Xf8F2Mijq2LjgakEmIRzvd3xMA9s5EspSXA2
MlTGdwIhxF7I9ugIJlgSt/M/f2TNHjHqTVEcVBxlDhgYnd0AVYYw7lVyGoUmBSL3
zquoPPV59tDgd4j9ojtHiK96o7zpMQQl4G3SRBFz+XwG/Yu9xJfWWFF11Pu95O0/
eshT0GaiIU5AwY3092oL34G1k6gfMcWJ4yOKbxd4Ztjswk6cRubYeGZhMfQ5Z63H
O2iSjNc6PBtAx64SwyNwS1W0uD2UmaCvc3Uxxy87zyrIsQctsW+I+CDP+ef3uGqu
GAqBaFbd1PXXT/rF0Hg0KumkVjh2mkmg5opMFG8LN6WIpmTgL6O6QVXM6iu8/vBq
pfB9eIxZskp2meDPbFQsBhwuA3RvfDZaMJgJHf+H8LNHpywdz5hjD6WbgSqWUH4L
c7tDYX0YMPlqXds09iiISYUlY/W8MaosljadULuCfS5YsMmcTWzwQKftOmSf2Dz4
531lyzFQXU1O1ACDrfG/Ur1jS4ntdogH7NCh6o6nKmWuAxwXW+ffJiBMc6ZaYUhG
lgq0s9AGHCsYb+zt+PQ3XFYhaCQ2d9x2pnS1DlqWps5Dhf4Vyp85KGOrnXZYL3hs
qBioYQQSY+eagQUJuj9yR2R3eLUldXvCxFjDMM5CABfkwn8O0dpZwng5E6klNEuP
PbcH8AEsgLlX+bHFMG0BXAwmvG7nhCnAHDmsXaQR8Wz2Eiv/6spztjGndWY5Q3BF
R1un9vQHLVOLjdIH10+gbqsOERlENX6AS3GWZXs+SR2+Xjy5vEmiU/vYCvjEHu97
BUX7L7Vg35tRJuNia2gzPusAlY6TvsjI/VJuaPP4MuM3r2tBvr75cjV0G/gUXM2P
Zz+yQCrMHXAwblfvR/oJC+JZekZzY702nxS07HGWzJyCiWX5fcCuQrGi4PYQWeRZ
QR47RfiN7Dqtsm2uXbI18fEPlB3YEG2a2kTkcRA7oRX2q5amRtw5/OdDMVsTm5r2
XLIMZAxZ44y/Z8i9d7qn7QM6XwMjZJgN2NC+LImhX+ZbVXl3mVsZi+VQ1mxUEIB4
iC56eVj60Wj8QnAEThXQ2uoNTQ4ltkaPgnkBEM9RZtvo694amvySURP7n31hMPCl
mq60Cydh318lWET5R48oEXpaTJeTjpE0yFzv1NuCFjTjaXA27SVyabtQNLRVAQnI
OtzAvLPrRYtn5/bgL6SBqvgxznixVzU6ITTv9WrJbW6Mk/didBuDg3hMcXc9pD4c
ZoD9m8mOy5Jzl+f1sJ1+Nk3aAhGPAJ4Gsmcbmpqr22gfuExW/I6GoVsI7X3HIwQ6
Gd0Mkl8lGHImBJZttDboXRvxRD10lBVZ45xLRcWRWFkpptn0O6G2Xvq9CoD8pZz/
NJ/KOctZJRAgxbMwMFfZQ6QxkvREpUn/slMlBL7cbLFOm6+nVjsGyrg0lTd9mvsF
QYJLeHDs9A0dibd7GGUccoagAjBVBF7E5lPoDzM7NVoFQjodalKt6E42z+M1f9ki
dqxcoN3D1qjhdSGvRnLtUgAQm8FOR0sgiigO3uBad413B8RRSCRYlhLS9jv0A75c
DZWGpfH1Z+tGdE7++RQ003Z4gcwJXpTRUyr6otdDAJ/fA7Bn0UjEhE+CEArk1Ri2
D9JxjPiFkO4b+aDwNXTmG1CbxIxf2cyTmJu7R8CsBbOmyb7P1pcruCXG9Se02TPv
PDK8BlPvpnmHl6lmga2sqSK1LY/NcQyibKRmCVIoxGc94gQwyGXMLLdYKawnrKDl
kO7X93SE8t8jd6YM3kM1a+QmyZxnyelPYdpJ5CYk9YgC31619AxAiw5/8otc2hqN
HpgwGop1DskeHf8OMRLap33evySfprr/3gkPCdev6phX5tVGQwos4cQl7VQhIohu
m5IJ9ecSTFsHFw5aXNsyua6EO+SN9eesxHF20d2DoSD6v6UwfQCO7ZORfPQ9w9Zh
hp83awej8QctWqGDZZAMlLP5GXLmdJxswvylcX8ROIsEbgd708tpBWp30lTifr4h
SmE1pNld9T+6JT9LNyQRXRN3KNizcGzgNtc2qmxWhfx2HyuBa7XIa7LRHKzEAPqW
JhEvhX4+V3WpKfPUSpEedPnF2mwIBIwE99JxevRBWJa8cjjeQjjJl7D8TjSrqUck
Q3DiQPQKgbB1cIWEJisqjgiyjfz48dmTuvoILaU7UsSqvKlNAo+yDkogoAK1y5wJ
FK2mSrxU8woyoB94bN3PcRx0DsRfQcrIhCJNjY8TOJuD6L+QCg8SiwvnTqkbmIbD
P3/MQdxCI1hKiuXf2j6hfTRUAgJ5bUswawbiHXe2Va3UQ9MWSMhFaoumbhkjVp0t
N8Tcwevk8l9GzFe0y9XM/tGScuHRW07nJVbKDPpMx5zjOWS9CJsa55SlY0QQBzG4
hug5ThS6w+muoAHL4Bi4GWt/M6BSd1RB8bYsRqRz/rwIY77rV1nWCxQQvY/N48BP
5MH4c1PnUcft6mQf6C/tHTsH8cdWFcjVerQdHIt3jGTDHGRnRsRA8CWENprN4XrV
G4L2vy/F7fFjcRxhcIPRlhLTUBk4Ga+JWcxlm10pPkj+rDkTzrRHkCPr68xJPMlH
C10nPsIYPtLFz9o4AdzoQ5+KumKKYytPXgsNiced8nP9cp+w8iPzusgOOQ1JbF38
iMRYrj62r2ICkgTXAT3q/rjA8p5dZFVEvFtLBUEtpDinbGc5bSGSZGLtlkjABzco
s3JzUCf2n5nBqSFSyEV28ZHR6fxFqss1/ycSnZhdXpRoAqeeqQw2p6Er7EswmR5N
W0H49wB56X/YlhM0b3C3vlmFkBqfkRJhbXX2Q5x2J6TP5RyuZRXO+2j5tLpq7CtC
1Og+rfH0ZX5w7QcHq1LLcGAzWHcDAgX9oy5dJUsM950nzRZuoCREfeqrsPS1y/g9
X993g2egyv8zbV/J7PVU5G1faDJ8Rbf5bIpjaz9v7xbRLUhzu9CkaTr8lpS9QkQs
SOp4UaOHgbBga1KQX2qoD8+20vdSvzwwRywE+dV8z2JlZdeyAOxmzOZ7UQra9aQW
QyuC3WOra0HKxwEhHM8ZlIB2qwACxQRh8zcOfVszIef5GtbvgHR4qQn+8sJzIidU
xxAyiccjf30PK0O/n53YPmltV9rax0+iwfSj8lK9nk8=
`protect END_PROTECTED
