`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mWvu9Ipb0oWlv6dk+lnNzfsPI4lZsvXM5NXWYxVTUViwgl7B3FCHq3vRlLLtCYMF
r3SkOoSzhZ6EtL3+UtgkORitvDwzUsartraUOGcU8nYQffqB4W6MjPGS5OBy6JwO
Vmn1ui1drUt3FfrbFF4M+OcayJfE46nPWLW/MY5lzVzjPc4JXoudKHJ43nKw/AGM
`protect END_PROTECTED
