`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN/4LnIRHhUeP859EHcZ7kLUeHd07FFAQMB1EaEVeTay
SoBhBteNkXQN3t/LtGpXYLilfbVe9kVMyFORE2tenIqpJ8+xcy6Kvvmr2V+g25K5
vBWFaL47E3jSkLeLMkfkFsTORsP/B3YuojRfVGiFn6aBw5BqVKkbQuE8CHiAl1gc
4pOfmTOfJPSn0evZfS/UIWyaLxvwOldoFv0UAuoS6FdXghtcwaZH2Z6d4lIj9Wbv
CUJlysmushjhF4pKwbgFGxtqv5yhdD99kEBTK0Kf/c79khBaEsRx5iQ6ZKjjgk4S
byl/jAl4oXg+bFldyfoGBLoFDb3vUeN1NyKFH4vcjnnCWIPzcbWhph4aMmoW2uCH
4JI1LU2Nq+w+aig1XomeEGt4jKwaVKTMoluAWeU3c8EOWoCS4bB94d1DqSAaUI2s
opi8/LiTGjJD791vFAvtuSR1Bp15VY/9DhQxIWbDrRETEZKOx5+Rq6+KQBYXHb3P
Da4clT9gSPFME+BiSvZJjOUfko/K4c2QLq7CWBM2Nhh0Tp8x8aSQ8pxvqkCzuR0m
`protect END_PROTECTED
