`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
PepsihenQm3vzdDxlx2USQDZF1NKGy8ObfXi2ZsYeGih5v8xGStKqgKzwqTmroRW
Xe3OTQOpsede9FKOaLLvYRII6y8d1p7/Z1UNAlc5HFHiumzb5X2hkvEI01T9YpT8
zPTWnfDa6X54DwRH08GL5tizbmknnGTmwS2a1zElQd+oxVWgpkPVc6nCEs3kzyw2
+xdzH/ItIhNVGOhn1Q3FqMjXACNJ2+FfiJ2I7ej59vHaVncWySrmFLpYJBPRhcA3
b03Qn2rvWdekMzKNjceJKC7JE/hixOS85yYqZAQaEcNnXFtqLIzMYEtARrwQ5UcC
ZkyZMsoW+fS62phbQdyEJrk6Qr8Xr0wkluWKz9Gjz5NdU7WkIBND1i2GiMaFZf7g
T1zVEZrHdmiZxisUYVWWEsl1lYFJmvtL5zF/GEh2fr2qBGCegRRJ+u9IY8X/NgTw
X+cBwYIPQieRJgCSAN8TGuDpWFyxD0GMZ57plcy/WjJHg1kjLvLCN7EE4TJOWYnf
YWJU/Xv27ok8hWmYbAbhLFtG/HWTxfJj0CIjsY/W1iAd4jsR+0JpbJz+JfFLsIOU
sG9osLkJYUpujDvOHRFBSjn7wY2FYcxxQr/WVj+bch9ajsz9HDGQizUZxqiPLwSB
Wvyw2ZJyCkGHeCgcndd/PvjjG19VTGjcVANZVI7w/ZdB9Rir0dhxLpYOFUWWlDDn
psyBPyk4F0IY9b7N7sZeRs8EgJPj6vo6NtQQ8gilqJmCSzrnRYeC3gKUIQeOohcf
CnVA1jBK01KRdni2wzZKT2Ub4UHxqiWBC3921A2Wt1t1N73228FNSt0A2867F3aL
Isl046l1NM+PDjRiWdWRIZaZAyDbGHKNwAqUTKK1azi/Ikk3uEkxggF5Yy9T3ffc
NT2cpiytjtgBMsDCUjxauoBO0+3/Hk+0X/coNGOPJLv0yC/PZAF+Nmw7WI2RBofj
j0y0jKldC3tSXvAc5ldze/sr/WqtvLj9mYY1kI7t/WB2hBdhx8ct8L3MG8pCqIMU
LpNSD4fGkjFwTpT9n5J8ix2wDPGsYkXmhzCB7cVLTZoCFJpFyINS3i9Y9zP0LwnY
0ARmn2DKEHpYSSIizGRsyWbtJXBHCSV4UOncRca05TMgx0H6qmbQ6qqMkpZL5AhY
o2tq5vhQNBJKJ0/SPCWbDBmVcrYPMNvG2UneSCeTYw179nqwgRtRRNGyPG8WEc+5
YKMophg0N+Gb8q3jYblnxqvxG5qEDqWUBS2KIfGHkJeuG+x6yUSy/Yju7tYmBLy3
`protect END_PROTECTED
