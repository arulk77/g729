`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFlfeuhaMCsaISw+PHP2kOQzIRtwe0Lcm+3oneYc9AS2
r/lpnmoJzeqj5/7DJ6y1V7E+lAlRpO6qtjHI2ResuSKjnl4PDddAV4o69RTR4i9S
2/ziZcFA5Itvm0o5VJPeV2GjauTFjRUDPfxNdWhsA5MfxOTCSJ+89S2wQxON9YZu
3OU1qqUPMonrSe7itbsHAEYE5cOXP9yQM3TheMT13rLFLBvIXLGebZPsoRiMRHGq
DfLs9XQC7lYlThqQdMPMxz+fcOOXYKiNyLL8YDcCNUmuMP6XV6PUIvkYWs9yaenM
uQC9v1xL4Kozi47uCUQAKUgb8Jt8e/VFermiTLJ0wAZNAQMLqJc95Nc+WLlmptaD
xniQ0WCrA37V9vpOPw85HA0UnXo6e+kizVmm3WZiIsIlP4l0xBY12QN2zz3XeJ8g
d2uv5EAdhy53HAMnc2Gtby6D+TR7peAK+xKhSZv+9rRynzeoiT+N2MWbQtnlYKzH
sfuDtFP3ij0+/eyvALfOFJDUGCdIQOECvalEDcX/lt++kIoDJ5CPYivgfjWmTpm7
sguCv5s8JScAWEdVfRhXj0rjBdunfrdkKCugPNuarPBZijk60ySb/T5X2jR0+twf
U/TNjFm+M9/U1GN12MxmlO68nUdHWOTnKXMGyip8dYTlZBfYDlRTgowg63wVePJ6
`protect END_PROTECTED
