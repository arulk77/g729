`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKudqdPVWzWs8l+52HEuOF97sAaPfbIT4r/Gjd7L9h5v
WOU3wzbMIVwKnzlFocUsG28l9zc2aa+TGy3/t9hqgq7X615FTx+hcrxVIefGYbN1
r1r7GIrEnLYsjGu+ITHLaXmUpzVuZjog/SK+lRjAqCEW1gtphdcinKeFIf4C6gwT
FHYMpmerbcf70zbw6d/n9/TPVfh6Qvowhy7dtGnwpYmojICEBbdVqmE9z82cowtw
PBCA+6ItbM6rmPzk/9GjqJq52IqBzg4N/P1pqCEA97k86h0wTf+tQ97A9nSODphM
Dm4IjCbVzze2vf7Pl54susNRyQvoc5kwypKZaJDj9fY56g1HQ2Lup48/oAdY1uK4
k8MZcU7ppqIRKjc3KkZ3SY/k2JuIhZh9RFcR2LMTo1ieaIQ4elxQiO9B7JHtlo6C
4N4yP/ESMqu4qZ5upAQnPud4AtrMiDD2/eJpMxKXHrJXQeqhoOjU21nxrrAEoyto
VZrHYYvwxP/O+QYM+UcSRb0k5oY4ZogH5xr0qd0mDWQdDxKVOQFqZbht7W9vbidZ
NHCON2+qRFTsvn2sc/k7oCSV3e0Mcle+2qGKoVJzyKJc4x2jaX81M3KyWFyzmP2o
`protect END_PROTECTED
