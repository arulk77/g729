`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMUHN1UPBuMFXf96A258nl5qDUX4iaGueA3EkC89KQAC
VE2eOr8TFSf6K26+hR752MKc4JhU14VjS8GRehIS2KhdjvDS3zP8IMnWs9OhxP0Z
zKhezNf8HTmewB18GaIC9cNIQSF6RsSt/M1F5b+I6+UTk9ONFdC7Pnaw8hn+bGKP
`protect END_PROTECTED
