`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
39P8mWpkFgF6JUyeFYe6PCPXWEvq+bmrodPebtswsB/FO4KLHrwp2rj0pqej8Euc
J7fJ6aEChtiqS6Ljl0crqBcJdOXhR74rVeVHM+k9tpWtvG09cazpJ2WIi7ZqmrFG
L49upuXfqlQMIOxyYcbSglzWxeYbW0Yf8lCrnJf1DntpExkWdMuH4XHP1eU4mgbi
pijeBn8flVZyU32U59ZI4uNCY7rxyOkzcKZ179mEjwM=
`protect END_PROTECTED
