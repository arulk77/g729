`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
a8H5OPZEoTtjmDtz5AkocVlFiR9yMNWHtT6as4J7GqY56IrKm5E/U+F0riyPO6o4
ch9iXpsWe8RkoveBNnadWlsFk/lJyMX1EhXhJENeMo5mNBnC5cLsOwhe2hnoBEGq
CIX9IUJVOLoxIciP//qFFURkmrzyDzK6L+nB7YyXOzAALeanNj7UgmRwnoEtE4Jb
`protect END_PROTECTED
