`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
whfZdEhQhIVICrvn0VMg7jLXoi9FgQQhrHfMC9Y1vkdFCFQZA0XC+Ue2pMHQnWvi
pLVLXMnrhiCn/hlLThGaojTWHUsIruU25gkh0Ys2cG1fQ84g0gOnpqeDdOh2WNWk
+aNM6KnXGQecZmmbPrsze2XA9PFRbh9c9ugcr7cpuhVuxtQ+WPdeDoWQfJW6suJD
PWfOfpCz6/OOfSsekRnjtuitHSzIIkljwBIGJhhPPLCZ9i8uptRcpHOthhr2nlVv
PeuChvJJmWMME5edWpyWFSQfHL4XTjh79uPmj6RxgKf/OwZ6JJ6zOviLOkDv40XY
`protect END_PROTECTED
