`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP9c7eMN9zWcrDkPD7xD3eaD853kSrakU+f5eCGI8ZY4
iA0MJKCjWcH5qa3tz09RguzeeE/CfliMjA9cY53l+Drat7Z4Ck6GamAOJJVFYvwP
9EaOgdgwePxISNaD4bVPksiSVntbEqF9UFGod8QSEDuwJzOoENO4+QcMI2AqCMX9
Lmf6iDEvXL3AOfTao61CpI9drt6tWnJs2R+HkBoxsdqWoHWCbK0eV5JTZXbY9vse
g0EyVac9Svzrd1R6/a50yOvwS4ql+wnAc3u7yczorxppbN2gHiBLICcvK4+NoI8u
0Zr25qxFgobGJuabILGKdGhhX7+RfI/E+lk5YzcS1kVvS8UZjbMo+RJGBWvYYIpm
uQIjuAxpOlJ/e1nFRpnnrQ==
`protect END_PROTECTED
