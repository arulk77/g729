`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveASMDMFgt0ZLFsveNLXSNcH72TflA2n6m79l+xbtFNSz
jtCM+E7WcQ3SZzIn9INM3UbvleiWr+y7IanLCy7BFe++KxA81+34e2DGcTCHgi4B
KIvmrBBnpstC95eVgkhZsZgpjZ0d9UAmj01kKJCBZ5Nza2JUjpy+GFhaOlTHttOy
nnoKCokUkvrKMxDSRgSq/A2M6YR37/yBZVrMm/Xp+LZo9/Zo4+oRIpOjSVcFjoem
CoantN9uKBZnUt+2OqlnBUX876Ph2y1MIXZms9HTW6zVScbuMKIj3JY4VJGIBrqR
voZ6A4POJc42UbQBmkTfCg==
`protect END_PROTECTED
