`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGwFuV3tBbTRmgBM5GeD9ZNkoWPYs89LfLCpmsck0IOx
qeozJ2Z/M+u6+jSDcxWPqfWFs4OPAUwcO4Vd+2lTA4DQ9s4XS6KEAYbMkp1sX1G6
z5hQ0YIlUoLLn6eCfOZFybr1QWu9oGKlC1rNl+RmJ+AoGaT83dROo9eanw4q91nF
hS4M8F2Ejb1MEnKpboE841pmwnfqp9PDMaX8XrPm8RJg4fh1OQ4pEEPYC+/lajuE
`protect END_PROTECTED
