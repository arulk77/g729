`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCbACUNgAfwvqWLyIa+c5oLTxSzEqUYwbrzH7WpcEWQ8
q9pEb5+xgP28CkMK/xiRMvVI70wkenWOdPlSFLrPtt+dKDTdxZh74ejMCJFlehMG
Fe8kvUW5jzfjCr+G1lU+4seocvkxU8Lj80mSiBLD2S1qVwG2N3w7w7vz96pXdyvY
LZcI2b57Kq9zN0+jd0lYVgdvAsGWGPl26+FHRaLng0dWUhGrdfOCFSl3sHHmL0f5
J0aTzTMw0t9T9OQp2gFskwgaY0mdgFneqKRvfk0+uYr9hchdLzTbt7ypWzdPmgPT
HSr9hC3Fx1Qc31jx8+kUAc22IpoHj8T8RpkxeokBCpkNKOXWFVxmjc+CYOw/HpED
OPpah+ZJr9/bNuMYGynFLSxrigVOVqHSQdgNImP8gOaS++8t+9CcY570wUCP0Wc/
hKv3ZMlmOLIdjwRgDRf3JNkE7KUucFJbE0D+6nRrGtIA/+7dVL9IZlKK18FCbLqO
aZkv6+k1nvQY11Iz+4CqndN959qwTNe10Y3EiVR/vbFj9W4OIdy64/mWWkeEqh2H
OAaLR7ghUx08W5mw1ia1bA==
`protect END_PROTECTED
