`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wy2JAL6piEF4UM1BWxbkdMkKk3XbYchqndLuegeq7S3
x+03sHtE+nSnBVZn4p06tLsUmJAP2K+6m83WAu3eWThAblFeF/jLEalcnyGMXrx8
6YGUjwAI+exgUOndpjyK4bDhJ8PZ8EFYwk3z+4TfmfWNHtVsIBhqrJFrcaHBtUJQ
XIRaupsa3VOz+48S67OYC6YREektJVECFVi0yMyJEZ//AM1nKd6MW5TL9BtNlCYJ
5NwaGBSPhMhGuRE923LjUjwol59ysfGucUN/oDGzTql9CQa/ZKO0v919C/nu5Pw4
LjUrAmg1O28idum+hRlDGQ==
`protect END_PROTECTED
