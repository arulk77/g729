`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJlSQJywr4NhASUxGX7W5xcCGf+N9agAFZUj5furpLmG
NL/T3ri13QpZ6KK1nvVjOZtclc+AUkn8/eOVVVPOeYGb+ZnPU2UQq+mojfQmOIek
HHswAk6Fh4KQearMoeWi/cklO2AUGj4eX0wOnfsF2wVpETKVs7l3pFBN6bFiuKKk
eqzWW6U7cdmGo6HNoRWXIg==
`protect END_PROTECTED
