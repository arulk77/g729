`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB7Ly+d+m+JoDDPkUGX+TpfO8Vo9M/GXhzvVU+lRuZGY
Pwvjtn6m2BTzjJwW1h1gvY+x48RZ4M2tjb2uToPjdi5F3oBf54h/WPaZJ2vywc0z
YFDGif/jsvaLJNj3DVIFpztEdULPvl+1QiLQukzylwkelFdGb7WDWHAlEwVAKcKb
71FLGKsPdTszyDaKe2b+HjHG56PJJge1N3GoJA+jlWTMhMQV+l5DOrU7XlcyoYr7
BrZNKZDde3ynD8vxcXpXqcpdohmGzW8kEaK/uMo0CUWrUskrCmQ/jLbv0B5XlY9K
ho1HTx3zJoFekI+9W/4soB4EBKTTkYUe05AL81xlNA0+YryU18wht77r1W5ccaPO
HxLs+whv3MeSQP43YgJiIOJi2BoFsyZDC5k5cua1vEvvOTP6w18Vgjft+ugWkM/w
ENITwuJ0a8g1JHpJxvQ2phj0+n4TPmgLHQfB8uVy70RHloJK1zeRiU5DghQT9X4M
xOGZSSfNSpukmykTAXMO6/kQHecyIPE9P2o/9coXJjLzu4CDAoSllsaB/N6i/fgU
`protect END_PROTECTED
