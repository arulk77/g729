`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIDLDRWyBwMDjLmV+2jpwQFJl7zilSFCLF63cqq/z2Ef
Tv7Jmj4H9GcWNr3EpbD206oHLv/MGMVugRZub0Wj35xS64IWxvJzCasok/gzPZta
0oxBk0oD3+xGfbdvwdgQNc53Edm05se4JaqJgdGDuTazG9BG8ofCuCr51X6jKACU
NBcpTBhpOMBF2eaAmjpfTxQfs1sQCxRrthqLFhMcDQQWjYHlUkpQZy/oIpOfE85y
7Ks6pLLQZBzp3OVPDlEmusQ6YkgD109tNSdsLUgqsYiBCo1gmhWdOAmNWsmqz0EZ
UWjzH2dB7YKB3S9nDKSEFKc/heepIpovs/yW5jjTwgLWqlOjQgHqbwuB/Qpczg8s
7f9aXVWesZjM45I068VbtQHm+QimKsk/dC7bV3oHNJVhRiuiZ4/dCpm77q+ypi8g
`protect END_PROTECTED
