`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJwnJkC+f/bi3/2fzWt3Qpmb1fyTJbdOGmJ0BoqFUVNO
nTui2x8CgbkiWM4ILHSN+AO2oKVHmUEOT2/ZLXtq2RkMysEocQlkNcFburTnW4aK
vDphoqC8p2bjOmvThpwie7e/8XuO/5cEYX9xCMC7RuG5hVA5GtMhyuwOL1gQeMSG
cHUdi6u/CnQ/b8u10+0b1GWFgWDIduWwtVzynXtBAahmtlPK/enw0xzUk4fAaT7+
qHape8w+RTivfXD9XbofZ6QHEHOWoEY5ILVdGVWAapbSc5vYjgczrlbzZNMnl3vX
Ywp9/UurKQmPvEszHxKsywcqadA+D3CDohpYzgBe21ZvN+jEL90FZ0mhMyyRAnFg
Pak6swwnlYYWEE/r+pIt679Te3wUDmga7rwfkrEovyxz/Wjhq9uFKDc/Dl8A2aEV
v9nYv0iEbASrSkLL/yjSFEk9ypGopm67xIicZkmP9EoRZQaQmQUnSHgYlYWtz7LX
q7wsPKX+ZjxFPLzuXyTKMZuDd2DmQ7Np+vHPEDZJK/L7Ia2g74gyp+8Uk5HJCc8C
`protect END_PROTECTED
