`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAw4mncA5TVFsSZ40cQCVGf6nxd5cfIWI9Y4rKdIeTxa
8h4J4+eispOreF39kZJivs5zAxCKiY9fG2iwPDniI7JtDzB5IzaemsHIzz21GBMg
NPB9P2dvW86K/7GexomQeGB5SOnAVwFf5YfhwfmMxd9YJ34+4EWxlbmNLpISYtu3
2qMX6bS7PU6SNwA6tPDX3nqtWc7ThqCfil5hsd6n1WVwnmcxtJQw3bZ/DRHupDDM
G2sIsE9zXg91NnoNq8i0b/tupYEDX6YUZdqozHpMs+l4/Xtf6mHMmXvPX5toFQbt
luNl003Z0xy6/VuDXbcEUbLiNoMWeWz+/DFQlQf6rf+7lyvvGUwzYRF7keg/o3JB
6Rkjs+MJthXGdrFYabILh3jhjTz8xsCfkZ2cLIu5sFCe6WpBZq6aDeVG0fGuGfKf
4BRiwDIr2uXzxBm3r/brlvVRYuSTK8rEQZCNt77UuiFbzSgWAvrwUnNickavmoRP
T9szrH+MlMK9+9y8sHwj4A==
`protect END_PROTECTED
