`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43HN5kJ3I7cK0WLrLNVyrX683MsxMDe7CAwKuBgNYp1A
M1GV11NO3aWQi47wLIHTXo0NQPRQTE2Wgl5gsUznpydE+7RWLIYLtmPx0GQR+CYj
YG6neioKes9BiA4b5EZaoc7oUuC8nPyjU+gUvM2sbfJRmfO2c8KjwcXetxlugKb+
n81oE8uKoBxzJQbvWXC2VKaROoya04ghgGJ3TYQoqv3nN5uiVGUqD3GMYwWkCKYQ
C+FdLa4UDPWpcgqhqH40ghYZTVy77VYOfz2dRfD4kSofd2PuDRWJT1dwHB4aUqNV
qB4dm95Qvb5m/ugzs4AwCA==
`protect END_PROTECTED
