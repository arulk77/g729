`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDAP3nopac6+aJT4ArgxUR2bOJO+uVEzz0uWDTGkKkvx
5C0sEAmB414+KKWuAEu5nyoFqQoLiVE9u0M3J5xAoDr4LTIhF03jKDyF873Vspn3
x5Zav91TWAf8TSzeFDS1K2CaNrA6FcU3xoYumGikxM8xtm0R7FTLD8AnX5UzKxvi
4T2xxBQ3Fnt9Hwd6cUWR2Qam29tlTEW9g0W14boJ9I1Xr1FTLBKKTk+RQk2yw0bb
Z1pqBGc9I1eUij2wt994BfChAvd3FiBRuHAlof1aZCzrYo/duRr9dR655eF4BXLb
UEj4YUWxue0DUqOVeYZibfqMNb+XTprQcUhzY24pKuksFkaDFvtIBTvFEVbeul0f
LUUUHY82ObvK5JXAI8dyXv3tefK+nIXZpjco58ZqHHpQzkY+qFgIgfsaXELEx1Zd
deUubZ4XGpGPPtNl+s8neGpiF5at3dCmcjrj8YQSBRE=
`protect END_PROTECTED
