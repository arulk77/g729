`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42B2zyYFrSRAyJRlXradD0Eo6SGVr13l01aaRdhx1zDM
+tBDSJfoNJx3q6Cn+RQ1J8ZcSjpEKAeb/QwXvVxpcPsWkz0qr5f3slFlKa/9h20d
v9MT+0q2uM+ResTrJelS9hnLEgVJVmOVhM/hhZjcUATyAcdcGYXGMTEbuqDWTcKx
LKlfjcr46YdbJQU4xBtc++ddlC8mgulnJL6/w2LbI343SPxcyIBRxdeVLt3QbgYX
PyEdh0xUSXqc3p9L0tPMLjhZ/Ai8j/fR9vMqp1G8cQv/Wlq2ac2HHrT1NJ3nd/4f
kwJI05diL3ukdtZTAafZNyugu5iJNFDFR7niX9mAyDrKF63p0JnLz6l6lt++RYPi
yIGRe4EZwraSQ9tgzxs5oA==
`protect END_PROTECTED
