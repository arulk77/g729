`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu439b3H8dY9NScInDNypt1YMiJDHlRSti3YuZGKCi8b/z
Cr1Lwmslb1MsIN47qt63mQKzefiXJCU99Rf9A53lx55jtse+DnUuT/J/+XiTTpIS
9cN6sfgNWpqpEvSSH1L3BMpKLWpWUe7ya9jpB1QDYh7YEBvfiJM1/petYo50cgd/
rp9eYs4af5riCP897stwW7DwToT/KFruuGWWLDgp+7Po8HyrL8qfHf2Uu2t2lPMS
Xiq2Lgwu+381RsMWq/SghxeIXtk6LTQEKk3OjQIM5MQ=
`protect END_PROTECTED
