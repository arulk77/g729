`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QNw40IqJrFvY2E8HYWz+j29lkt9/ertpAlzka7MwLhKYrA/bASvWVdVBwI60IFxn
O96aNEW+iGkZJnU4x8omGIrG+oh68YpbHN4YXpA7l4yIycvG6GFYuc+OZIP35fTB
hweA/p6S1Q2DJ57V7BM6f61piAimHFhtTPZLPycJLmuijZCA4HfoScY9mxBR3n2d
`protect END_PROTECTED
