`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL8xE8q0CykDkphT2o/2/ZD1GDDgnoWJqepvq/HjmCGpkZ
t8DAY3XK1+566uYo6tGW2h7iu/4cXqe+oPghNvfxqh4F1KLps6niL4bA5D0D2YMX
bLgYlBJzMHOHUzQIwjCRYEhxwhfD/tmTCim2JIrfLaUJyn88p6W6H/XWrsKigFIL
BK16BnpHukqJZyVI5sv6gJsHgdaTrxajZCeLsS4gZugWBjP7RC3VfpJzcwyUeHDc
XYMqlbHi1u1i5WsNmLYeMgPZ9lpo8k4ebqq/toKUt/hDY4Rt3mu9nNy1LxXbQwS4
wjacn0+dblYpucIWs6N9bns7Lyek/Oq28SUeHcKkOl1rHR8tjF5GMgjnUcNeTHBl
Lvgrr0Oj3yPFNZmBbwdtEqlSLI+X0bWK3uUmjL0TxJc=
`protect END_PROTECTED
