`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLevy2i++6vkEvwZ1fjR3YEAKijryZPhEnjce3GhmGx2
/O6SOdvNs+gJoT3qLRDiqBqzqVUDaYRh/taIBb/mHnKY0a0Ue9Qu8htVxLmZpBp/
AglnLfRawkb4edAfiwW1ohiLnWIdlmzoIAWRCrlOR0mQa4ZCu3EFqP3aktsthy4N
N5eWxJ0zM2pOQFSmEDfbUeB645rcM+mheO0Co551w6L431mJWpOh6dI0NpH/IxBO
9Fpz1fByM5mpcUlPwz9eKLUDqVGDMzZ0TwhYWD7R9wvE/sFQ0zTW6qxCFqPS6kOs
9lEyGPvQQte+h1Xe/3SqpmOayKZq2llKXGLWjMCEDeQQuYpRHLIdCsk23z9jszuh
hwvyCoJv8+SJ1/dB7cicFg==
`protect END_PROTECTED
