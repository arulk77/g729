`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
RPTmcnCipoYoJ8G1tSseRL2PsjlgecejgI+WeY3JVN42kR44mgFV2N99ojcsLbOw
sXNmbR4H3VYbFo5QkCHcSZnLqZqUIaeAjbxQEZOSas8HV5E44ZAxJZnHnk4d63q3
Dof0P02WrVmn88r3Su3SUqJWDBmVBO3049GLVJ0lo8Evrz2QK37fsW1+v0knnEN8
xxYUoNo3LreKK6fdAk3R/p9Y5Do4fQCK+lo0J0hnxGOOOWaAg1fFu9CkMP1AUYgJ
7K7S+pRDategVmF+9le79k/vCGagvghXkEPTm2sY1idnwO0WSfMY9jJEk2cTRaP0
flu0gzcXA0E4cxo+9sJyXrY76sRMbiozwKtgVQkXM4Gt/rBEyxEUOM2FB5dvvm28
0ZWPwhInWlo1S3x85b6BMfwRt1Oyb5wOjYI0Bi5xPiIbzZeukEUOsUt/nOWBpDsk
/GVAwJCafcyEwKlMYfrlZMK/LIwFY3VUOZKNnQDjtfOhtw/Oy+JFJuuMHzZERBcw
vHlKhpHdCUxM32yPfef6smasG6uOJuf1PO1UwAvUaUlDB5XEezhfCaRNViG9Jm8S
yOfZ1E26ab7POvznB3+viFLIbEBNvq78dGVjInVraEZ5VYFeEc4KudKhCmxx0yox
ZnYNZkTfrtp/t4HSDfHM6RcNaCvLmR9eglOQTCJtzhXHYvmn3Yqx2qdTcvdcI4qG
nm9yUz8UiXqtcV65iQUsQgps1MYa5J84YLJtB3QTD0Vyt5AeQrA5Vc/bouLIfaOy
PNPcCdhVT2LdQ7DUMdeg/7SYnjzPPzWRKbnZh/4H4TKQ7hOQot4o0n5Vq00nl+Tt
DC1jPMdbE3ricoYXGadec/FADTkSpuBgQv0tEPt5BVBb66acdzvEhESCl+F0mRpJ
sYdssa0OYffplIdBHRAhngr/2fycTgRsVT7Ru8nZAgQN/I2kdcQqs8mkmflyh5k1
CcUwIrtkazIXVq8n3RouMoCIUQdtuaEWyzAYVgC8FJj65855zPXJZ0WHnOJioBJD
iM48rOp3jf43R59AezbVMcPJ+zramcbYCTOL2QEFIzehuhoIwLlRhv+gCU6Fl3e/
DTL8uRI8i1g9/kjNLg91pOFdonp7OcUt6fmbgKsfXC1ooz6gGjvIblxRckmAkcT5
6/iVIXdhrcTz6sw+eLMkUcF4x4wnTVIOsK7zxRnquhRrL0eKkroqj66ebUKPlYms
ZuqLAWXQglyiQvfNr87ooz1y7EOI8clSfJm2pEFqRl/mj5Lv8mYp4i9fZCHrfR7v
+DU7ZAeOdxOoZWx41GwUUXM9ioz7XKEH6hmRu/WKTJD0yD1+q8YT1Nr/aAxooeST
89f9PHB0sJO1SP97PLpuwjVVaAhMNcg3VZnrKoa9fYkC6wIhCo6YvlZUrkzg81rL
xE4OGnC/oxmdfAWSak9Ax8T9vOoN20GIezgmFWVmP3AjBv4HM1H6dOBVAURt47pJ
GqYRkLKBwSOBBA1KaBIoCviaWpanXgC3w77Dj08nh1eCzAkj2cow1eL8P3OPTtEt
AY+JVr5nhkr9zPnDiXrpWsOAJEacoSJV4oPby7iMNa1Ezwd9REvAOJl80fSXrgGk
O2cx8jv+5PnsrSAwtOCPTWdqBcLBkY2KasNUjSM2iQl8+dLSDayRgMrW3MT64mwT
8CjvfD4BS/xUXx67ZS/kTE/gaD0AkOWnD8EnfLiN+yFcNagBwTNAtHCJ3T1ifaWR
ybn9d2//BFFDz9cecWCYl9oU0RbqiyCe+eHSxFBYRkC9plTqhZdGb1UJUSQris4p
Up3yzfsSeiioLB1z76dd0ikbJwrULYSKPjrlkj2hdCjRw+9gCd5NRvyus3OqairW
gJkSa+vrc6dWTm3YvVQTMBbvmkhpPGY7Z4ldmV44oPtZj4fLweOMpp5zz823Tj2O
YGF2JZF5ewYDunImr5+vdUroyiOjDUwyBySeZq0CPzsPcGHSUVefmr/TB/c0hEnV
5FyF2hru0BewCfbFiivNQRV/fEDFudIbcGObRLFNKlMwkPScwrboDkKKnA3g35cQ
BzrOSm/GiBsdZONg+jYpVqhe9S41dd9ic91x77KVbks4XNoBsBlN08j6DsSbto2x
XKr15LMI4k5jzxtDDrhYqoZEpW/LY1H8I1d45AYHlQ4jMu2s2POnEreOiUwjUCb8
W76O8rU41FIePgOh1LdZWoGC8X/tFo6peUEsABQV49FnU8h0PRrLvhZuHx6S3SaX
P2a6DEtVG1c4ZxEtL6PT2Y78BS1H1AY5AWBJFQA3GcDuM/j/UTVE0AG5EqLZD6al
eXLEqGSA2YoGX6AoZCINRmgpt+1fEZUjhTxs0UN1JtuSfuv3Qn/SgTBjBY427SJU
S2QteSR9fazD2UMboGKV7J/x2RLMLIkbL/ahxWwaK6xXCN9XQoBnS8NPktEjcRNo
z/KfPOtW0cy2waduFaEg3xwMqYqXWD1L07ccd1f30qbYwVRQ6+yQSvq5plF46WdZ
Tvh74aE58Kus6Wgn+wFoR9WVAP1uVLmHFvoI7jKeKP1ODJSGt0cVGCWInmJ9jOpd
Eiht4T4MtkJDJndUN14toumKfXzBkThG6qFPk35NOAzpPqVSyibvvH2H7Y4gjWUt
/OWnyyZ2vvVHHckgnYSvMeTjAqkqobpCnPXp7462EuLf8EXVrnzydbdUQla90boe
CDnNwSLUbi38pAPiuuXLNj9POOtgtbP3utjjzzNIuID/x5qUPbkrtnfwQQtE/Olf
EvW0jSfJtwabQoj882PQM6mVCOGUkZXpAkv0e7cN3/wdgMM11CsSEGPqKEgzycSX
eZjC3YWvniT+6OWM3pHgtiLo/kQiQloF/yaXah9zgzNv0a49etMKXb1jPT5MTxWT
XSSF3dwEJAtunww7ht0GQCaMQC6LnPRX6poDSDl6q+Cuu03IImbsHhOqTIjAtlFs
F9tbzh7113y4a7+DM13ZjtmNN2e5oVEQGP0auuIKIi+/rfTbO5O0N03wUqidiZO5
bMQ/eMlkbkFR0ERunf5UZ8l3HLCJoudcAfRrmzemNvknMCy39GMohy9WkGq910Tx
azy8hzKgkrBfb3b++0be/KdVM5XDu1QQDDD0o3W8XEysnFouTGIWF7U3nj1RJYbQ
hVN6JYxGrCmdwknvZDvDnk8qt9jeRAs7OtqiWR+AriAb02zVqfJDazVp+Eeqkpvg
O+vapXZsGIQa5Pv4vCVB3w4w9SsUYL2kWXMxY3QWyH/CPaJqhG0V/VM6oosmRnP0
jQyVNNXbGq5iC2wdApXXiVU/4/efVOJVZs6F7G2noEsTBnubeGvkHpEMIWIiBsz2
wU5r7pTBc1Qc/ezsw632gpR+oYhUTtnJEo50zOf706wu20WL9d9mLDhcz1/6a7RO
AA9xc5BhUfnl5KVMofTTFLV30t8cTLYO5KyNNG1jrUFcvFp9Vp+3udd4KNPCBRfA
LKP+XIexdCq8uj2ADFSbhlljqPShpFoXUjyYqz/hijCAP686vxE6N85Q0EC3qN4w
v+OLEUUpMIELiw4mCpRNahxToGejSM4I/4slT5GXo/6Qf/yqRi0ZqclUfiqDG/X6
/FJoyOvOQlzmT3vn74OZkCftHBRZMZBYt4iAPEaMX+9ncP4pnwz/x/A9Ly408Znl
aHVN5IigB3yCuDD1p70c1E2k5DvHemkITr52Qzx0T8obiA/cJ8pKXOMBABlKSkoP
ebhpc/gktWNdnqbl6g6vJxDI+Hz4VnABjRHGtNXLaKD+6WKMQG1nVo997tgs99/a
NpAdDtJpz7UE6sMLIvmCCbwsYiaeD3A9Zk+o8hfhr+FSX/HOibGvE3KSgdumNCro
iEmMkyjai88USemWPpsrbisp74Eo4m6k3ZAaqfeLMbTm8I1jAJyaEFkHxMzUB9+T
UTz+5JG3xzeJQWlZUw0BIc/qPDe5BaaS0ODhf+FEV0ziaLh4QT5w/IBTjZxk1F0c
tGG9XZZkjB+1GAuRFnwEfoYSiIcW6W+lueaJG4xhsv+CMMfkUgyHVkV5QMQ1xX+y
kQk3GVTvPLKBQREqSLaRdFKMw5P3gpmdetp/oB/enqgSEiAojAd1axE6BFOF6jYI
64i9TAIVF1KIfzgqoeEXq/ArB4kjQvd1Ed51xnjbHlgCpMeBez1bnn3baYeIshin
jZjre/I9RkyjpYi13BeycEFg2Mv97TapZPK2et8WzCq3zqJqY+0IuAxSxmukPla1
SrEMiBz2Dn2CcckEjc7+0QYVl+wJNvM9KDloC98FGi1Vo4phh93wmfd7DKLj0egu
Ev1cFG4G73u5F5weDoBfhG5IefJoKsNcuAn319+wqlXPGfqTFDYLLmggUZE0hE6z
19WjH35rAy/RThIa/mCzCowT3YddtO9/mySA6VM4f7W5J0Tr3IFU1mpPh94z4SUd
nj6TaX130AmMU6Xx+a3j0GjNy4pYXAVV1m/UL8/iFU05SFZ3EGRRxiP2jwaZoQgm
9zREvm/6ieXB0Fp0x/2EHt7pELHs6Q4w6eHTj8gAKpo5tjiCLWy53xBQ57P+7jhO
/c+S7P+OISH5IaOrCGCm7FK5Ipl4sgiacdYJMclrYeXihMAj8HqdXWDcKhVYzoY7
BdnDHbZW9Y8FuDAdG7neeElxLceJaRGweYS0iQhNZAiGwJa9HZbbyBwSevO/Q6dd
v9TAivjq03Mz1kc5f8w+/0il97F1OGVrrcuXBXbdn0F3lNIdufDaxqqUIj4Sbu3R
0EL5FUfKdByJjG15X8eJ4H7kdvGNtZyH13lTxxRjna2olOr/C5wcR1z37DAohSAh
Ovvd7Sd3730QkKb0qmFe9RzHYAnpLIMZlAKXOQQaP4H9E1H5WOrgALahFMBFkhiV
u4qynHj2GX48VV3bOAH8kUeEwLZ484WXAJ7NY5cglpDEH3uQkift3UqSdCtiZmFs
T4GxN/CwijvhdavvBv5hO6ihZKZg8AWUI6eG1dJHxem8BGirp6rvZD2iUMi9a/j9
cLE90leMy8qIy6Q7AcNimmf38gZC/caDHkcbEky5fzgD84JorbjB+9CLplrqY3fF
m6Avf440SHorgxG0+wtAL5X+8S8ana45GjxQPf60n+FUuVHuwUWIV8fscWs8opAR
aewkndrqPI/+dd8UybkaXM9dK62LswGJhxC2qM72c/0sgrJzdTBMI6gDT/RHKcxE
p7HI71T+i90HCS8jpaQP8xE9fGVyT2cqO9YTBbiXrAw=
`protect END_PROTECTED
