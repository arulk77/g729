`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QrZgJKp6KduQAzFIyCyoK/mwwUOkoKbdr7DiQYnTpUj4m49ltd/tS8i3vwrWz3wh
Gbusb9bgS0K6uA8ZQHWyG+RSl7bxvMVhIDDavbw1QNBwW5QIkGgLmWJ8wyKCoVlK
+wyXFCpNkrUQbddiObzTzntRgzDhZRryThcxjq5O+7oZagwYcrIEiMq9yD4XsKug
qJYa1kRTmV5TeBLtnYTh1SuM/6KoM28HHhkrtNGp11GptrUs6ymGWHujoFeOkmrY
YhwJ7CwvkahhoudvN7MCav4VFkdw3/0KVi+F2HPb/WEQit33mbzdDlVQd0U5u56E
kuBkOWAFhpeR3v/UqpBfIsgZ/0YyjN5BIxt6TJcN+5ab+8PVmFnJuf8xNuVRgJbo
NOPvWwEKT9JdISDWLu/9OvJo+DXio1dCoSUzJ3ruGyqRDqkolUDZwkyunpwB6bhd
DmuYbNxoLd3ac6NCLISauzBjmLeV6MjPbtn0b62xaj+lr5jXpSgoHP1ehWQE5Mma
nUvm9flezmlklTes0NY7OR32tWMhScMyLquZzEjXKWWdHLpXR8hq53y4RQ3Jk7pt
ohFq/eKiof4VhfDAo6QkUXkMmCQC1Z0uGyTTGcaGeVYZxI2GlLdh1kcLTGgicgB8
S6fUzVPlHLt1XAaqpLYyIX09p7sDA1rqsjn6eVkKiY1QoY/QywO3ZTzA4JvL5y0W
MIgJzCN+cEkup2GZK9sw0bgfQYhdBKgB2xXcXnLDU9cSJSYRZUNKdw6aM+RGVpyY
f2ef+0HANbzPcZkUZHBAPA+71JkwnmMib6IvB9Cuq6aAeHOK7CWVrefL4UcnEY3Y
wPGqxTV8ngj7VnfDo5heiOGDOMn7o5j3lpYEmqnKflU=
`protect END_PROTECTED
