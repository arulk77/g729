`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJzRmnB/tFV2MFRxLrDLqQ6keJMgz+KOQL4QXNMY6gdK
Zp3z1itqNtttQiaKwcXTUWK3m8soqHDGfQC2K1VKE/eO0zlg1NN/uEgNcFivchcm
enqk/sH95G7nbNu/O32wYXA+tAKtVavaEZKA0CQdkW4z/S3FKwBeBeuoKuur0Ccg
rmT5Fs0QxXQBvk0rk/ulxw==
`protect END_PROTECTED
