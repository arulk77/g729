`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4z5iLUz03Lek8x9v3BdKB0O2I90/FwKPyodX6MwkSRRg
Y3TBVmpIg5cKnIuzgLtHKJsruCAyk6lABkKiTzkuSYQT4wdguZcV7J5ZpJRH+s9e
iPjzkrP+DoVUjpOYhZErUYPOFb/+DM0ZB5+hS1MscIw8J183J0VqnACwtazqa9pX
kVUrbVoZfm6WqfJL60+YmVsApaUHM66F2bxJOQnpcyuYHLOHRPZ69nNoDvR9o262
que9FaI4LxP7jOwQ05bUy4yvoPTSMxK60b3p69LDeXVOrO/i3meO31PHes4nGnXP
zwZt+/+NeRVkRjl1IBYhGw==
`protect END_PROTECTED
