`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yfFMHa+j62inm2yX5VuTrTXC0YkVS+79IRScyGbTTBN
GpXJQEES5A5ApBDTIS1xzXWvWJHLagyIilw4I/cOEoOdBJiEUO/INWKq8TSeKNRr
nblyRtRy2/fbfuHPoMojhfI7A50MF8dPrxDVWgAuXfadNr4nVJ1l1aJt9TT8XXL6
Lx6dXw4A3k46EzfKCPLx+dwgXo1KZNbTdcrhHJZJx3Y=
`protect END_PROTECTED
