`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu461TRulUa5U3RLyMbaoLKYYDQc8rDxk3AgXON/XPxeaz
uP0ZiJYjnIAgjLOptADNLQ2cZAjnFspAbEqTs03idkZrj5CqOCnz0c69S8rNA/3s
S40Cg/qG0Uy30LdhiO2gIOjHQmCknuE2RPyv8onK2M+1iCSOD1uMW8znaD4Ae9SY
ImQ6OnsGuOMS2XQ2kB1M6VjPtvJ0kEtrj2hYMC6AaN5ZkGs3v+QwdokcA5LQ9H4o
xyFgkC8hWu+6jay/QcPGOYsZ0k2RQRWuAhx9nDdwt9jBRLcutMb4lRi7OxTryva0
+OWzmSBG9/9PfFvJAwY/AEnP1Fi6zBY6JPR1HHYC+ZPnb857nOMfaCoMgmOh2KOW
pZ5VgXJh11zRtp+D53V2LGAM7l4wA4Z0b02o57POVYbldoqTyUnVaXzxl4+gj/ma
OtbVCguWwNlYyPkzy9WYTyzhTXBg+Uio73B6wRFFZV+20OEPIMz2WOL3V6JRrYDb
`protect END_PROTECTED
