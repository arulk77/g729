`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHJaF0dWBhT+9R731RszRG/VNJIEc2mp/rEL4aJf9VVV
nIiM/vh9+BXZ0sa+xTT1PmsALUjYsBAp3pnLsTqQx21ea8U72Wz2KSaUZ5tU9O+x
+Uy1hdQlBN745mNJ+ONbmFo5gH6CYPOh/rQDrJiTXNw96nnrJWFjqMFL+pYUq6Sr
7ZSXf1yz962kFV7SvQzg8pZnjFaGoh5NpKUwzZ92FJeWIaxVl0Qt9cpEp+x7lj5c
8ky6uajK4Gj/rL/7CAsNzB41u/dnL3XyATDoOhKQk8dPXqAw3nKuUG1k/YSNFIU/
XY78x/lxISSp53NvoPhGZ2y25EnHDBmiUS3ka0PIjcsoscy4KIPw4Uu3g8U3WbuO
ekTcZpMdugnAnyTgFCpzDJCjFHovCmi3X7lq/lQZxBZRsxxQvV2/zuSe5pjjhmhL
l7tRB3shOmdAnzAE/T7cED1Ndw87jgTPHcuMj+z34yD564MP24Lh94V9hhvbI5So
gY1Fdq05D0MhTd+pSta/jhjPKae8eF6dD/RQkExMDSxn9gQHsopiNYHaI11R7ZjW
RUo9aSvX3wd1Jvrlcn3uhw==
`protect END_PROTECTED
