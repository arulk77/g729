`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yqHTjIDx5RP66yYm9gF7m9rfcuHOMrFfihnJE8WRzzX
llQd9MixL+LEouMV9a+UoeWiEqzKNYFvWZJ9guwJNXZrbmO2cESi6ziLIjwsqaqf
kX/L8bvNbohYL3+X/gwsXurDAuDwqHrsak1pFf747YUNKovVNe7NmbglgEdOKoSm
K7JTMQK75MipioaZkkoQE9DC2cjZ0QmXtF9CrMvcsuLGb10XKvsSncnPGSeQ41Uf
51HPBN1fIm/Wz42rImUP9jrrArOLJ1hD6hDi7hHQ+AA=
`protect END_PROTECTED
