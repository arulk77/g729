`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN2kHzIMy+NMDut7oPdmD/9kxs/ojDk9nlTCVmNcQuyLu
pf2xxQ4SxK5TU11vJvFLKWObftk3axKDgBl6rYaS9ZRFMUtiSl9ecwqHaeJIZe55
A/VGd8d89LpxM+M4xNC5XwgDo+MzGhQPHIn0emyQWjGB2y85aQhQpfjIhF1kueC0
lz2B/qiVOu32/yOcN7eh3lUd83LEhczbtlOmMZW9VK8gdZ5zTwO0XRtG08C/IHK6
jWkz4+Q+DxFFaydIrcxN5KBaAtz/ciAIayPCwirPRfF23tbLmh/8XG8jVeK/yq2A
VLyyHZx6YNo2+gtpBmgkvzKy89NDPoqGVIR/zKlb0Hjik96XcyzxXvWslrX2xHGE
irCep+cF2bJgFDGuIZ81pERMUmkYTrGO6+v/mJvHvhxdrJtK0RQhtwJ2eBF0CDFg
r3V/SzAieccspm9XCYBK2n0sNKvaf0lmfTLeJY0WzWu5FYz+YNe+iUock6lAQEo7
pVhbMKMo20cxd6HBohGSobURIGf8xoUsdo5JSoYSCfkF3IlyChvkJG6R1AFZvTkU
/Bi9laGWqSViooHtXUdIpHBV2n0TwE2asZ4lFI/zVJbEzC+pZbGwT50Q5LHbo8qo
UbiVXw3EDHN+wt200jxnOAoumh/ZM0WOu4AFq4mZrBt/UEItaVxywhqrGpjh/E7M
tZ5W2h9TEpDoFHOKsLv0dGCC9q2v8oo/MDagXUsGjtE8wy8+DfarzAwnyU9BV32E
+xEk0vLvXl6TtuWUqlSAVjMixTFDFCArHqwMl0iGapIqwinR7igyEeRv8HlOwbsJ
9mdo7K85yUWAZPQ1YOvzqO1sdWHgA5w6QGdAuOq0hE9gAUOiE+iRhzK6g/hsoXgH
1UVhrrZEVOzIMGrmOkQfQVjS6fgVz2+nZzsAtgLNggFS+nQicWMKOYk2l6JBUt0U
gFiEnIOP2sBkpV8MJPAC6qNdiR3a9hLIPfDRUYocMlzDGXAu9E+J9719dEtFCzZt
4/QwIIgh9QQ4DQwqO/NMTA/TNZq8Co+d7h6iw2OuNsQ=
`protect END_PROTECTED
