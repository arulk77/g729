`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHb4vzZt/rppNhRPvuV1CTIHNrySI2lRCdn7cRP1wu/d
o/H/4KRE3EpK0CYY7uk2OtrrOQ2Aq/R4w7U911MWmT4F7k4gH+9O4Eh77BeB12hX
woh/4T4Atn3U2MyMknupi9RQFMDu/68jCD2gtBnkdCX3dm2ybkVZxwffsuyDdPe0
fEm5Ttx7ViAQgw9vPqha3bd02o0/zlY/n95O06ZnZdNtAFE1i0C0i3UkYTawLOmN
POZI+k+kgenhTS6IsE148VeWI3isovzxAlOIofK1opaELi0u7CBGOP1moDb0kI03
TIONMBvflXv9iMMymydr9rEsVlglNvgmstqvpz/CiOav4J+R1Pllc1Vxv1MJqTCx
xoyn3cAdP1WByNUnjSjIlhjxzcX7FXoRNFdbSgVKXnbdjs6b5aNh8YN32YgH8fIv
g8EovDRPcroOb1OCX+OOhA==
`protect END_PROTECTED
