`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+tpJMNsycz2JOK0Ljl1xelcrx7BK8TDIpEQ8oZ6cgDj
F97nEBl4e3J/hSmno9JH6Q6NmVQpnYivbR3Rb0q54V1Yo9tQaO5jsl/c19TQO3Gp
NDK9/gdoAycFNBGSTxhUK93AT3ty1g7ggprsB0HJt76XwoCzjtBwxEJVx302ydzy
yf2D7xxC3zxMjJkmxcpGRSAmGMFwlIbl55sk8e8xN2g+bhZVfbuGksQlOFzInANW
zDibLPIgWXq4FLGFmKQMN4J9Zkyjy6h//yymxIuqCcs=
`protect END_PROTECTED
