`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAe2akJwRRlEAEOXmLRvddT051jTpy3ryOwamqQAjEPyt
itq6VebnUI6e9z/BFAzQkcJScr/rjiJGDWWKkICwgT/IpLP5gxaI+8yfAdnHCoD+
tBysDUaVfWWRdb0qNJKfQK54UVEqk+FcJcMpzgNHT5uQ3qssHgsxejYOKdtXW4nl
5fYjEHSm+bB8UCOmi6RAFyXxoYwcq99Rr5Jg/xEBfUzDHSlLGtTLtzv7q7j1c/Nd
jdmNA8s12iDD8o609t0YwtC/eIKUQ1BnEGwS3v252muYYAoTUkAp5SDeFcLyzT0N
GIAKCKPAqzPUFTZnalO0mlnmrXPip8MEO1x9k8DZOByvlAOWdApsXnFoLZ9gp8Sk
09BzM6fJoAykgCXz4X+QRoEraY+hr3DvW4HBSUuip7LdvvIuWHtAN3NxIkflJ5ug
qg8DM9UL973M1VWhk+yQv5p2AXBAb/DrvV/G1A+j2PDTt2XJNJYxSMXqn/5OrQWs
/5y4volDvdZcTiWZldiTXvg64q6X/Mr2cZtHVeC7QnIPdJKmbceE5kURfo9wvyrp
chAcADtqVSFInCBePUKRMkfILANap2bBTrInNS8KUsgK+L3zZ34As6y7QokQg9s1
ahCPo4zknRNoCmguPNqyV1r2fJKa1sAD0ukLv5T1zSRqyTwxQY16JjW4MaikVH+Y
SA41yzOnh4WoOST70zp91w+yg7T1lNRUREYy5E9m44kbSATCiS68Op86rK3o6URf
Yq/JOwvSe4CQsaHc1/Q22QP4k1D/dli6GxZfKqtfWpFGmNuUBOPD/ekWEtz5NnEJ
ZIep/qmKvqRUdF3x95zJY0/S8xwXmb/3e2fRUidCDF/DWqQ+Ub0GuRKpvXYWwArW
iZBwqbVFlpUqIwXgYLkwzMgis1LErD8Zk68klQSlv2R6soqrtRRp/ulSHuZmmghi
lRYoThCUtOCANesP89PQtOmhQFrpbl/R5NHwS0j3v6LxoOIZT+pRGqXj/SA4xQjn
NpV69x6G7T/BG7AxU9Q6fB9UxgnXkspJvUJo7LZ7A9xRdxGoemMtEDALI89OXZ8F
CJ1SM2zKqm/m/IC8aauc4V5anzmf3XkGWTSfPgVEe9u6ESR+HGRD6J+PJvmt5CJ6
G9PJPiMSd2yAaej0Oi5QFSnMufqPpJSdv9DDH0MXisCq5YGJLfROPuC8Qlv1+jxt
CdiqYVEgFx3kK0ZB5UWp2AhD2eZLle880D1xWvqYhIidzsbJHHLyAeWcDwX5r8K4
OMOfyApVBH02yx058OGiis+enR/mOvylrDok2SbkmWdm1ve93X/Iz60V5ONRzQ80
sETz/o7HUR/5akVT7DNsYkaXI57MzBSXDsxlNRHvmY7DaF7Z7Pewq9ynceuvnth6
OsKU+Ed/XEn7GjlCYCY2XynLm/dYM+iS1P6GbWY1u7uyJB8ol1/BwB/HY2ICh7E2
zblAsJQVcQpBqwgXDwqts9cNx876EEJUXSB0x9ghaGj8kTlgbsKTX2JtI/jY8FP2
O/CkYnQVgI7SeVcwO/XqCqVN9P+AoYvbpdvSMiuxO15rgGfuBNWbMYtc+FDW4B6X
YYd/KBNjDErk5Jt2JLebt9Gl58zOd4NJysZ99cS6W+Uls+fc3B8+NCWvdniScsay
tghyftlESzatg5MvRnx/W1IfXQEC85YJIw6njMU3sxlhBCwL9PkrsE7f5l3p/XV/
75vG68nkbUijUPnjUxv3KPTgH4knadi75n3Y/lYOAMcm4Fe28QpnSboJv/7nShEa
7O9IU9V+WN6bPk/3aRvFFwevtayunaLARhWxsXqooqIqUq7hUnHy6AcW/ORiHROi
Hl63l1ZK4YQxyRql6fKH1KENStOPWYra/UlYk/AjgNfNx9rON4BOpueh9S3y1t5U
3i1PzeJLhKqdaMd7VtvU6YtaIvFHN8vuzLkvyzn6MEhgGoYX8/u0o6QQLpEsfZA0
rKaVkmV63BB2xDVXMNNxfQMi6UXaiS418oi8IYK9odtD0pKiZgkAOZdLUZwgzmij
7Wy6qTLFD3919ATHIao/1KbUZccAl8Y5OJaKVTML+8BRy18zAdGF+HFDt8IAnC1N
iew0NZyiGtDPdC4//t/0gOeQ75GLwa3s9ku1LXTbi0MNEaiwMTl3N50kLYqhpUnM
OJuNJFPCwXxLkHGeSrVISmywFJtQK5KyVjGqzNfcxWqr/2bvFvrkHCMmgYzyJG54
pg8DoCCaSLPhzGwz+bA9v1fbcj2pnrzzAIbO0swtEUfKPIKCdk68lQ8vcxIWWffG
InQGdwfbY9DK4TYF3LIp5HSDezzumqNEwpmsOHXd3Y5mzfI+ntPcTy1/4d23WM7z
ZJJDT4DGO9mzmNEU2QepzOF6cYv9Cb/qVJ01lL2WXylSf+4DaUsWAKgAgjlw4qNs
nyftKFN1HF54YMONVBUd4eqLksPDmnxBJNWeUCuiFO4G3UmIPM87V66CgCrVUTlt
iPI4dEjIvVU7y/C7+jXcPMA3DDSb2vZaAfvKZ2baEpuPJBStxsBX67VFFkApr6kK
ffYyIXXpgmRJN9BnKfxeomhExENZLBySh1Q+tS+AA88QLS3vdz5fBJleJe3DYedD
wUmYjjDnAbJJFZfDgsCWsaKu8gcVrWRT7LeLKRQZyRYlWJysBwxCquQaTKk/CwF2
l2RU5RJoXBXOifPXE5JNwgAknJVT0zVP2jil9OuUV+YRhcUvSLCiZ2mYk1vqiNYD
AEvU+bBsW21AXkGvAu0JGawlv4MM87idF0fUdir3gdwFOorQpG1ntIJda36Y2eur
Gz5dU3+J9YAi/Y7ZyyUyWl8Pnjh8PUY28f5e69rrAqphc5nLytODvzKzKxd/2Eos
UBSVLwbOtPgSRK5HSTlIE462K+6eRZGqDYIiMpTUbozQIHGM16jylMeXmG3lbnr9
3EgeHoDLF/kXOqo5twH2sXwG1oaib5QBs5IVg68ijiuHw5QhhcgdVq5dAKEoI2yJ
6DBi4g8ktOXGnlXxiMgff6r4WsdoV65XP1ZI2FQxjCICh+XL08/Ko+kuh4Wrn6IC
lmtl9SKXwvPC8Frn7Zj69icUDEo1bBD9h8rzYwuzi3AyC4mfglKhKpmUlMaILsBb
diKVkFZkAewpENuvBPBG8Di7Kw+asxyqKbzhxCQAS0RJLp+v+ur9wuMfCOBqzk0M
jnFCxLvmn80WKS1MxNouqaeMv5yBxrFYIdi7zJ5fx4/Xq7xZz1gR/GZQFn+1bl8Z
3dpoTopyQ0yV/P9YgqTq6rfdbvSsLRroHPzjZddoa6JgDXdP26lDiEl0DGqwjhfl
pWtvxHHiNe8Hha5kFE/8UdWVST69Y2sckJGrlue88OnizMmRpjBlYF0d64RT4mq8
HfdDIXIl/UZ6/rfYOEZrwK6gdXk2HIWGhoCsi4/k026gXvDiWFShi7FTB676YVMw
F62bDsALAa0IpgoBExX/nL5IKWZAbXIDxbTNYOFKkOPE7aBjy6nFUjdGcb8f4cth
`protect END_PROTECTED
