`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJOA23K4vMeDUZMhPRi92VhGQqkN48UwsUkloppde0rQ
tqnxvPsHX8x4LfLohOVc+Gv8Lu5s7KhYqfyQ4O7SPLy6MlklZ4QKQIbJCOK3QjED
CZaFs2dLgezXQohUV/utcbOrDo+LG69mtj1TH2fByZqQhixzZ4Yct6zx7Szc/qFi
cCUV6wzvUwMdE73i882XwfsY9lWgi7UG/k3zs7tyT4eVuH+S546ObK4tdf+Mu1Qq
`protect END_PROTECTED
