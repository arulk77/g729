`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveO+2JJPomYO0i27/sWVMui5hyACCqoyv7y2gmyz2rf82
FJiJ2DarcuhY76NgAQFIOyrwahVCFGdnKWrYelM0fT48yBBnzXtQw/wEEACzq1Hk
sfGIlQZyVSuJ7E9x9z/OJsu7kAf7O6pRF8R5DwHYIQ9g4ZhCsAAJMe9U6L/tmjWG
2wAx8n34AXfBRPq1vF+VxTkwZI6ddHjFfJY+kFLOn4OKy0lUymkAeZAtaRrdETCG
`protect END_PROTECTED
