`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
f6g9dNvZfV1RXfzD6AbWWVmBUr3+dHDNODMRZS8cHSVBL60n6GcUwl5rnHdkw6OS
1H1DPAsLaSgkq14WS76IOJ96z3nxeinYSdBkypkOw43+ff3vS1Sn0XVcJhTT09Rv
FWlbpBTD/oZybChpM/CzdtVaSzgZYVPOytO+l3SlBzf4NmnpXkUaH4fvrfoXUk8g
In7az2fDAtEyyLU78ieHbAcIFBqLUWt2YWWfcClhAeXQ1tlr8s1RVXfi9ftyWKiX
Jt5cxYLykV8707Qzp5TqACDu7MQ1qDoroVEIZTpbGjjiQNKP6RiYk+RU3ZwxKfTL
5xw82UsE2HAPica8L6H6BgekEgkL1Vo6DayVpHmPW5f6OatB/21lw+8pv5yuBS8G
h1M1MI3k3ix9M/9QC6GfxG+23eRMgcNje9B/xbgPnlKwFdiLTTqk2o0vaVEjwbCV
fq1zXOTe1+mx0r5kS0HjoY2z/hmK4mpu7CE9MXtCxr7Y6poCoR3l+XQAkN8h1qrv
io2GLohCA8vDskfwaJe0+xV3SjHdANpC8dIyntF/HTScBmJRg3+6r2vpm6qy5X3w
NaTAm7Cuh/ySiI5Ln1kao8Vi7/YeCybZymM0fxySV+TnyWui0k5C7/Q64P5UQRrO
PPVrNwxf0T1H+UrYYdebnHsgGmgxi+YPAyZE6XNd/mgw0MSfae4MYo+MENul5Rfn
sPe3i1Lv4knZ/1stYqyiXNLDh2jqD41GVYxsibOIBykcF9RCne83W16NicwKoJvp
PyLUKgmzdre5Smrn8D9ZEa1oBN7hPiXWhd1Bp087nD9wVCS8AZY+KQO++4mpMBma
+EsxoLoL5+tpdiVdf0PyS9f1fo94qk0InyRtNK2eIoyD1ZfuutM7KvYr/ST4BVZ1
xWaQaEEEKiEP0crOYdbvGwlvUn4oEeo99e1uaND98IpRT8Ht8Rgthcb1YfT7kX1l
zU7Gjdo7L3VSV7AM84UGacPK+0Op2LVIVdrgfszLYsvgDt3QaV/u5IxTlrAZckgO
rJtvrDwGzG2DKx9yGC09wjp2whFQuvdjIR3H82vtkwlrFVh4GrsUlNSybdXMCM/s
g+8Ai5h1GfXoMMqTj/l6LqeFUnXgwlsf/AjPWfRq+Z5xiqTezTHtwggHdaRn06T0
2GuIEnddRLPBR4KIEaKQhT2xy7bKqXBf025LKQGzwO5s37EDqqy7CiCq63VJ7OLP
4FwX3of5P6QFS3ORi+NAZSpp+kYyRo0ofhStRMkvmiTyzaS6ryQK7I5BvAIpO9rg
GaIkSw2JqG9dp1Y6GuJ4TXDclmknAHven6tRw3Ik1x1BxrexTJuHNg6o0BooJlm7
HhQkAtvMZmjCS1mWjWpm0+XoaQXAPAPl+yV1p9f/zzM=
`protect END_PROTECTED
