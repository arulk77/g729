`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBLgJiyzIiosQrJn4OXAd9100+DftkiX8i9Nwoob07AQ
/OCCmimvTCmok9x49iE7qN4XbbW64+fubcRpcT4Io50FhNs3zt2uLR695ril+HKI
okoEE+q3bWFtXOC8Zn6acolXu5+YkWbUsNxHWzbhI5jiRRKx1xRkA0OnVi2dX1QM
28/KcJBPXmjQDe0iNkbeDwmUjnTu++jK6XLiGvrRMG0dTy2GuPhLN3J9wdzeYJ1y
DAGi4R1XVe7HQM0u2IvgvEvOALJ7lpRXhwzNVHV/anj+0YXOiaPszbjnR+rt3tZv
R8w9fmX3IpDxYzbkwxFUXgJ72Q1NWK9nYcpNx698RWtY1AQ8v36gJC0SCadqVrZr
b7O1AG0KEQbWRpHp5rXKui2bfmDQzaJIAVJgJ/Y59x7C1591glIM1UbIQ/n+UC8Z
g6qb8gOdqHaIi2L74gaj3Ej+SZQg/iAOEE0l91ai0QE48euehKvEG3vF/WIxDbsC
52zs4suzMwYAF8u3F9yGC5u2i9hM8CK4J0EpJVif1yYPZdqDbME691BGwqpxxxPI
a/YV6bbXwv5YhuvMh1Ux0UVDq0Ij4zinfc7k49BPjDd7O/7E0pgahb4iEMsyTXdf
9X4I6IlW9v7kN3pwNPhW2EkQ90bnndALCiXvbPXrQNZ+L3YmHrsD4ocWn6v8jMrt
E+DgA/E7t87X86AmYRKKKpKbNLsgmk5Qx1ad38RpHzLwNu43t/TgefO8+NCQ2SRN
JNyC+EfBGqDXDtl25N0g6IT3Hvbi2C1AG3kLBVa/VW12etuTAwxFEiIgaSO0Kl+F
RxhHsJIhj5IOqNeXwO13dAA6sFFrbrTI37fFLYT+KPcXUWgulvELuM7X9JHCspfU
nskDFBmCYAlQyjCfiLMPpq7FZorakOIZx193wOo62XbPIZawCAbg0Y3FwbztNP9I
U/GyrrjtpmSUY2CZxCqO9x1vJ42GrwuPizdjuH3qWOEdY07SUfkOQUB7Xr/bWze1
3AmVIPlJCViHhwvop+PFKM/v31qD2mh+QAejj4uPUvtYHhtoJkY2hh98YM7r6+kZ
ypNdVI+Rx48kCbdc9ELNXSgaRM3Eqok/bzOXyYjNu75ZhqaNtOIqa6IIvQU3Cker
bzE8SBN8PtkAvuXB/lypscbV4+8BPUv2XtmkS7ceicNUvhW1i4r3JbLUGGBfJ0H8
eQSre1ybF3RoEXgrd+Q28Vgou9WI/l/qR01h0QOvUqGQBqHXyHueZOD0qcXRkgW4
hdhZBSVw4OMQx5gD9+D4sz33RA7ASLSlbnKzY1Ah34amggKNu446V/Xj4Ox0RBjf
v9uygEGR+I9FGBFy13Fgp431HTCovMtki7tXLcdvbUUEjOxtaA+C8C4gnpwNiwKp
li3r42BLT56DDepe2UrrltlAPTAG1hE9nR3o1SN+os9YFLgpN3Fmvr1tMmYV2pK7
vsLoWCnN9p9lomdh2rFdeWrvBzFDF26QS8JHc6whpNyTIjNzTda+dq7qG/6dLT7H
4+F/pQeTMF1HkOjeyCPZyTf1V1goOIqh9x1Zh/rHQQ6sezCGUoJvMO3f+NB+eTsP
EF69/YxX7J/wFQzVZxnAIBr9dinH4hTF6vyfqIegJeI/TRwB8IkynqPpqdXVHvvg
hv7JC/p6xjy3nH/nZ9rfxT+tiwqAXLJJwoG9mj+3eF8Mq9GklAZIHpaZ2aIljlx9
+ABh4/exMHdRWO0LhUV6tnuwQXdmTIjC0YhNLM+fiPDg+n5xa1Fo/HKOvHogpwj2
c5BwNdQffxcO/xbJjj7pPrF/GvH0+F6B8gdyBmNYHPiQpoovJXAMpeGGJMo7M8Zo
QH0rPevPKCcjv1E1ppET3FirEl76mVZi0Hsm2eYyY+fcYorXOPgu+93zhAuZ93z/
gIqvD9aqyjeW0LyGswAIIC63DpXb5sHgDC1SYC89BoMuDVpQWo1+ozxjy+9J0R6F
gYE2YmzMaDG6mZgOFrxF3ESdO9UgF3s0PTVkV57d6G7DCMKOZeu/b+zT6tm39ktY
5N465imd2RjM/5DBgHGkSKLQVBlaaHOjrubhT/YKfzESHcZMbccD3/1kH21+UUID
xkwWt47zBXvPBny03yVbQrSSkmsHspTVgzQioO/eWZ2bPcgH47B3NQ5C6QlrTZRZ
0VoLmi3CQ0fbJ5yf7U0l/N66lceIbFx5zIfKckVYxUpa9YrVhJDMH3lD8nHnQqWS
7FzUD7usU9zhB8JWG28kLjYd0vqAQQyuj19+6oUyVLfR4Gy8xgKyxG6jeaAok28X
cYSs193lVmgt5IPiCuzCqKJUr2pn2ch5sGaUzGfZQ+TJNnsbqRtJiSYVSoGyCWtU
10U7UF2pAFQBtjz4S+ppYbAANop8VVRoY8v+ZrQndlSG7Gi00UZ3its2EDwtRkwr
6/XUzN+qkoN228/kJJJx7cBqIXZmxgsd65b85iVhiyQs/xhchQG1/cwB1NkMyJ97
GRVA2MgTr11FkXZw5ItAT9Vbia3ylm2mWlJX8gPRrKJ7G2PaLyQQFYqejgxrjUKu
dTsy7YG1VTlaoobvCk7nhoHec+X/V6aCCwgOky5jx4CSWx1E2/Khg/It7EMZmylR
qUPQRGv/Imj9pM4Ths7Ua6i1CYFW0GILz26jbC0QBZ0hm4cNHLJxlLcnwBid/ydr
WF+vgO2aXM+Kif92XQKN48SSHuL3tcWyURv33tWzZozjAOwUptzqSD7FcDMruTjC
Wcnrhfi6UuCyZQOqr7Snq7i7l3TdHWv4F+NJ0uO/oh7okdu+52VYNFZGAH5o6QHs
evqEvghXsSJVQGF4ym9MUSouOUv41J2h4RHQkzqRIVyTiJcYXnGj71VUOaZGBTT1
sEbFJdptiWtR5TDq4a2yNa53Vgl4fCJt+tndYxXNpnzfFBTNKFlWWOLHPOmb854i
+aBYhMtvZQCvhU7xkvL2m/XZyy0swjXxzgIKBFmDTGSn8vzPvZRJF9gVBekLewSy
vjhowzdmLAN7QA4OKaJ0lSsqv0S6zHPl8XYWMHFgDp4NeKd8pH69wcASShkLsbrl
cDaac4Xi6FgfgspR9Yav8XfrRcC5TMvpE28IHjR0MlevJPKPb5kHDOpQnZxX9MpT
o5unyJ3RgKKoROA8Di6A6cFEDW7osAnpXCm/bKSWD3kHyAxNtYEW08+6dLRpjq0J
J5f4Al+fnwg+4uGYIbWDgi1WARneppQfN1f62FPp+zNKHzIZGmk5iEo8KSeuHVFy
m1tJN7jKQL7hX0oYeOflF9ySD+0bIxMuwNIStCipKH3KKAVC6BRur27UaN19ZSqM
FEBVa1dnRH1N/UD/aDPo7Y6Ev6bSN72ag5Q5iER+kB8=
`protect END_PROTECTED
