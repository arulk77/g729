`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
9twiOy/OGlehx1Yk9XQ8PFi5q4XF4aZ5Up2DEghjInH2Jw2gEoQkCpDEQI9u6I+7
ikGiLpBpScoPLV5U/ejcvIcZNVHbsPQLMakuVtmEJpeBPjLDEGrZn4b3PeTUIT1u
asYURTWMTJzq4R+LflIdm1j90aWRnjMaMPtZ9/jlFdyaxH8otR7HaRH7SnZY/k7F
`protect END_PROTECTED
