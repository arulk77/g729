`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIDoK1N40OZs3hZJAEZQioaRlNzi4exD0gXYwaMurPGi
Lsqtu4FyXgtpik2CHXVMrA1ng3j+9/we8CcQ3kLF9Y/MDkz2ii9jE+TeYSNK9fjg
zziR1lwDe/BZq3VlVAPIp7b3/KtK4CW1wgfNQ7XcX5ZBiGbaofmNkKqpNoPBDMJR
hulsyoUa1hwomLuEeXP6zueoNbDsC+xddL6/VhkTsPOtFFp6aSJm6Zfzd3zPI9FX
`protect END_PROTECTED
