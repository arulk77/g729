`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHzQ53c1KONh4QbGcPRxfy2bieG2wqNlCEHpYMbx8SiT
DR5VcylaygHDycJ+2ppIW7HAXjTbpermEv8jfkuufCmrV2fnXx1zQXoHndksqjxl
I0RrFmcnsao9/CtfuRNvayL+oXeoQQAgDSNT6TrZnSEOImP3cO7B/E77JOkWe0wg
rFF13Q7GPCGqWMUjrCpw4LC12dM9LPe1D0g5/PklyQfOUWRhiqSIDRybHsa/xMl2
`protect END_PROTECTED
