`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48fDCWa5Fce7jE9QVb6H4FsM0g1GknXu6xiWOXWZ1VBd
furLKJQF8ojAJMqHxBLjcvgR7woEWEHMRcc8s1C39iXhHtNvuB1c82KtEGFppXel
mLLhcIBEoEe0sQ050UpqTFWo3L8ecsoMHJzBFi5y9NeUvY6tmzAaauNSM0UEvZ7I
cqiOotp3TMl6YMgXjw8fjWFP1ALY8+aJuDzpOYgESpY1+w2NuKAh1bdrmpC4k+7z
Pg0sv0SKLnXux9lTcf8GHhr4hXV6QLurfGe5iyaXebA=
`protect END_PROTECTED
