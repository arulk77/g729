`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
72DKe5MEZSH9IT4s+0rFcNte3wQw08K3UcYuj7+RYDhtCzBV3B7gSzbn/7qGAPXZ
apigDDcxubyAX2Bn12GJEXqIY2ham9nnwTE6daEL5o/t5Y8C7lRZpLrqZMlsS90q
Wi7Kfl1Q625zMcM5PSRm6QUZ7Ht3T54JCBDI141GJsJZeTtydpp3u77bjkzg56qv
tRcAjlxVAm44VOlEz5hPHljCCpdDdLq89JaGQK4CA7qCObDE1M/KhzIskTGsZUZt
lopzBSztyP89J/iUPACpQw8nTRoY6zqc4wv4zIUt89hHBgQmrLm08O5G9c6XjCUy
XAqxky6gViSZ3zVUJvBN73M+AoFYNJXOQYBVpzipZRaTjPjL6tLOoMhOV1wMjuZr
NpxG/Ph0b0+9pnc6OxoQl/alOqfhgWorABmBjCm7V2EggFIRcq/nE8FUL9h5+SQE
x9eV0cl9CocVG6fI04XN7TgYgVqw/h0yY7kDYjR1ISZB8Wr1AbBF35q+Y9gHQoKy
zByHA9EJIq4xdXI6Ln6UAFrouFOHDSns31Mj2hGkbyX+Xt65wpfLiRWua7beI1Gt
IukD5OpGQwv8HUfl2/JFuXjk30RJ7UgQQKJDtqP468USlEFeiY9UW0lWoNNPLzFE
0fNcGBDwu/xz5ZLAOClys5YttaYAJmiQkhSS3HnFRFXM+R2o2jYJzjHN9AsfJzik
2plyzVKl0zz10J6yO5WBHxBRIujeo/Y9RpEYPTfxt6digJjvU9bP2BIhmJEbKiNK
eo9r/V0BwRt8tOkieV4GDNKP+f6bjwsjI4Ys2mUSoWVJ2gCv3QjoDn1IXYI9FFEi
PBfsvRMfE+59DnpDztT6/xn8SikVjCbiiiY/F+zr4S+StUwcArg4Q++BdffwuaQS
TBkvS0wBG561Q9miCilPjg9Dk4y9YoYC9i1x764F7glWwNY6I8nsKeHkVIaB5kab
x0cOI1fTm/IwMdbwxjhtJ6PqyOv6mLdpspwNIFCan4hUhpUU6VvU7Wx0rlYyKpb0
Ll2RufwgHisPxyBKM02lnWw9jUEopTR3rr7zGTKQU23BwMS26XKU6w8m3yN1+FRO
+wLsWGllyJXpfJftGbdmrpdGQT7zvttadlnG2pKMabsgF4NsipR0czxIiIov0RYp
vkRwtkdzlXkOxyAijwGWZk/h7OrOnVsAzyHSMgBjvXFv043jxTLvTfHB0PtDa2eX
99nPe+gnW392k0Z9pbzQm6PjQF4tsfvr3MbMXNttbzBuSrqxJAxdBkDDleata34x
Y2CLSj/R5qzxS1aAP0CZdgh+3C9Kp1dyt5moGQQe6j2ieAhi0Sk9MzjYHvqrE8Oh
Vg21HFSucebhDyananFBtDa651SEKtDJr+ksrW1nuOHGryq7d8mnNXhl2/xZhSW9
AMZ4yMr8B9BZ5pZtoKCg/eOmV9IpFiHSaI0C8oMhZOtX+POJcK2OHj9w/34CK58y
tGmcfgeQfzAnjkDn+/2tCRE/gM8e1tLEY4GKpze+j+sUyrak8jC1EpNOLOr85WMF
Ee7X+Y/+0wM0TIRRsetxH+nIKbNFjaw/5ftIZlLfLQcVpodo4W00FK/49YOIUWIV
5UaRiQ/AQzBQ32NhC6hi2yRSmyOqnUe0kDjJqS+j66vqnJP/iigF8QEzwo/alau5
PI5HSkkuiKqJzKks8QJdnqNHHI/yM5WOlEwP9wItaE+l46fPSvsiZbqdp5wpEZE8
D8asfyKITRvUB6VMAIgMq96oogeneWXN9+8zuGAyn9a3BL/MAdGk7DXJzAvB2pRB
w+oyczQM3fb/AYuDAomRPzvozG/O1CpQtXrwS895uiYsZBtMZCNhS4VOnDdMY3jS
bLkSu/AFQ4NlxkFtrqPzF/baY7M2z2oF3ayxX256IXYngn0TPu3408XLNtoIM5no
OHV7UaDu0lou6Lu5bYkBK2ewPBMK1+bOnWEeTRxPyx6/OWpjIQ7MlIK04vqtvLWX
2HxlAAFAScVXSZHeNnoBMChXvrFIMni2d2ykhxyx1ZsjyO+a26SlNZFSEJrVuiMl
9iPM4d0nRjsm9pzSiZCGDVl6rqt8DaXMR9QNLv+KK+LCTIRDfYZ6sWe6cOM7LA/Q
5Ozq0uf6L2d6Syow56ou25uMHsKSb+PJVl1VJMna8dl4NoIHKbYV6Zk7GqyNPctU
5/2lvP6PUyw+WIONKNbRI3Y9S7BmzGIw0T+H1eCReMaWzDOE40JkcU3V8ePkNRF7
xJTTLWuPN7ZaRDRQJ8M/fE5SAfMfi43NJINdvq7tXwhXp04oe23TwnN480qsV4BY
y53325Z/WdfQlWEsZbr9Sdt0nda6POSk8lIyfZ6Ji+5E2+csc+831IcMMKjRYPkr
MdvK6ZjY6yBtGi//a7bmBfQCQQCa2ysF51HgHPsEv4kGUNEHgVWzhDX9IV2ErIPC
M6T4IK6XL60WWA6us6TSCtsz1ErpN2qjxp0JBDwY2eGLjidx8P3QyK+xaogwhau+
yxqjc+q8yNG6CE0f2klhdh3L0fy/ikUZVxrH7djSvl41VMIfjisrRSGRXlf2riwT
URVsN0YaazK3AE3GDG+bT0aFA/r3GLjoaQcrXQX40YU9qxpIOpxhVQMnewIuIHLM
49Gt2XU44Lb4h+CDuY/wy6nfnKaz4jtwiH3E0fD32vhspOcFtOEmwcsVZIbsQv//
muK8cSnfU5vXTCvfxAIZmX+aLfTMKsmf+e6KcFy56jYkhOzafd64Y5Xcl2SXFeNI
Qs9gz0qnWDLJNjkaVJFR0hyIkvq2B1xNvPuPmfCvjvl4f7eUWpsPVaYzX3U3Fi2v
S/3YDoMkRXbVtYnzsFG1ik0+OauopzlkboC7hYddMRGB16AEB8nQgNyK9YDNSAQg
lAleoUaBgp5p6Ch28oW+udCl0zuF0ccVTwv1kdJWTfEA/c6K9s7uiUollL0rJdWt
errMb2GJpMEhOH9RaMeoPP2JagtyN9RVUooKlJ5pQjjOfzoI52mRLvO9UtjJqCM3
AfdkuX25ya6DCh7XSGtbeQIqIw5EBBgY1nZxXOUEr+cBBZogow/9ZNxlEHA5W01b
PuGIvPB1GznC6yMFWSiFusOfa2dlo5uYJ97dDRBaVdTC240NNmcLXx6Xj7C2A7SR
ZL623h9vWSS+5xIoCFJtTwkQwa2bLKdxiOI+tDzVQDbc6/P5GveOhRJ6JmXaDjcE
ETVBTZJzbRUXKSowK7ZzKdJZxoFe8GXjQ5Dsl0LJ2defh7Z1lPZmycfAPTla74Od
ISMwNdybKPGWESCLk5km2EtwrU0+TWagDsK2pogUZoeW9StDzSeEcpiXsC2G0rJ1
ItnlAo/Vu1P4Ip+Etpzk7Nx57DcnESquUaExxRp/oFAizMEK40WDMEXyUZX5Le6y
COInWBOt4vKcAVr1BcCX5nwTaC9awtRqljHwuL3XjelNH3htuC0sx5WDs0P9Nu9F
jrSZ1Gchm1w8ZRg3jcmosAnJgtGG/xEJU2BnR+D2a0dMktWA4f6+fIF3xFuxNNLu
dlnVk1vbVSAZWXSPTzHcikX3xDuFzHLXKA7o7DX3xfKQ4xJQngtLxM60MZY+H9MI
+bTxBcL8CCr6JrdUCxtz2IgNRt+twClK9c79pH8mjh64SvP5UCVVW/JnKX3oG++D
AMMMRzkEXhfGgZkuIoBzT+dUi+WCuBy+2ZZMB2tQyA0Z31wn9OsbTY9Plo5gMzgy
iJetMRn1xH2aSOJKimZqZMPhw5gIoxddNe3JsublgV1bSJ5kqJGKsgzVkejDCr6W
Lr6tTw1qKIdYHWRkuBXzk8ywhH+eySVJc8pPVehM0qWGTFcV2zlGp6EeP/zkacD+
AH3h573gnDy6dqMH/pgtVXnktv4azBTYrI67AeyRC4LzgX/DKx5mVOpZHzh7bHfQ
oBC027kHV8cxCjCc66vjpQgBfFoXBPJEcstd/1X42e07xlvK8UoXhNZEQdyOOWY3
GatE2ea+0s25ibGo7onrFwZ0elw6rfKcXrdPs79tyGati5g+KE81Ks/64bK7YzzU
7M6SYdlO+NggYv7pWbfImAyrbfb5qNKfBe+xKlF/HzmDeGLGD5qjoFriisvqjWJw
5RGwuueon5/UXrdkrBFasYoN2Kky7IwHhmU1VVG1By6tMoEs5hDzWa7wVh1/ycPP
YeLit1hMPJMsZpwkwncuiZc6CTbVNwkA5RXxeknGUnIx6HlZyS/lQ7Ay+97baCzN
2C62gmpPV6SdWClqZR2sQRJ7N4ovh+T1+k5scS/hexaoqwMORAjigs2mJnrOILB8
4+PdTtOKjEKDKX6vDaY9Xh5KGaRQ/7oILs48j6wzte07GtuT8w7mhU2NGSYiHB9V
Oz3SfKQw0Gca9sU+6Xcrg7xpQs8w6dl9v78rxNRIrs5ftjJo4WOHNp6hMyqq5IYs
xRBQpJmPUawch/HaxjmNQfa0NgeMsRHaqRdpZnqmeENXqhGe9fJOBsRlAV+HFAtA
Zg9CP7q1Rx2wqMoKi7AylfScqDFxqBsuRguypxicCl3QVTA2yIRp4FYXHen32G1n
Aab9bFIXeUX2/yVloJIf0RkgR+lfhkho3qclQRRIUvKD1xoPToRtyTgy0HBaluLB
eSpHAeiAEulxM+3ZW0K1zeSiayrV4F965v73BooVrhO4EKn0//l0ROApWRuqPtSz
INZvvc7CEgBoEIAREdU2yCCU+Hs8rHLGCv5TcGMw3VePzaQKfnVF0YEsn5ujcgpo
+ziRO6NFdbqwmwprAW+5WT5SHUeldpTuGw6/KhAQrqTT/Vs0Su3jzwQu0rwBvrCG
vax41mJMyVkysy7Ek/HiVK3eUwayp8IdFU7EcMTVLs4umr7+68vh0cU44pv1HGio
3wq3wLi6cLMdp0pUOU1SO9HR+B0d0FYQeS2TgrSvQOt4Ct1Yy1Dk+nMEG40xEZCI
Hh9C73+ShT6m+qmlGAbgaGhiRD5wwR9NSvV0hqCPDhlUlep0vd2HffjvT6RVANAJ
8NVWJpIihzCYwxX4pVfFBBNnCcJzg9ewRQMmQfDLO4+5T69lRFVB0f/Rj+QMveCS
asnVZjFRkYc7opZ5R0DfkOOSc5VpyO3DAKM235NnVnAp8R+5fs0qidTYYMRc+GeY
529gqX94lq0f7ouL94a7ZeePERpxJAZW8MfycyGRCErBJTmP+PKynV6XRWgaBS8v
dGLTjnwV4JIW/kLjVYZKUM3f6eLU/JcV2U4duvuJVD4YL3VkyS4DfTjhmq/eu2TR
aC+SkclNydupmoG8zWecuGwh22g6tT8EHZLOgKO9yPaJmS7lmJvsvwL6rZSbyI/P
06hwmSl0OOroe7CBe9+3Xhf7l9KvU/qw54VxQNiMQvo0Wggb7hHuAOfrj8QOSuGa
E3rY1dxxtbg770kca3lWjaKabKFErBzUuvjKfnzU0fVwsI92lJAMgGE2wtMAT/wl
5pJ2p2mosYZAV4M6449ef2YOzpNeWulqOvbf4jPOrFetA3N245POHD3SvdEoFird
U918IDzdhm6LtHYmCPe2nBAnD0N/PyaZexXFmosOZt3muNkNpRTFwbEoUgF7eXeg
UF7tM/jc9aUigS5anv2VppH9+cluR3YaMWnKJxWjOwhGYjhyRehrY1Jog44M7J24
kCvTq5s6ljlPoJXaUXhUoL1z7e6+dC3RUIwdIgPn/E52Oq721Z94Bh2Y3spGhxSU
MvtKe8w31qC/lzZ3yAa6o6s7VdeMRyyw3kym+nhIYAOctV86dB4oUVZ4HUK1SOA1
SmCwyLyZwkpNbhEaA55vjCi/ktf/n5fjNGHEvEPxMhf/HDvUX8f1H0lxfFiIy69h
5EQi4+Ngvt2zkvHHxHiN/1dW7u3DgrsYoA7n9Qiz7tCvqsgJhh4zVh5dyd04EZOh
ZClZaTYVr3JNkwpPGeIuFHuZPzDeNnlT6BhryCWF/GHp49jLGQXXylcbKzZaWGHz
r7YQn8O4iL02n0FEdeYTQrNrds2xeM+erm0BoJRWJNUSrF9218XCjHSnP3uYPtmK
Ny4sJvFwrcsqp5xSmMWK9GdDp2QKfJGHM+wX0bXnz2tGZJjGh5I2Mh+YJQWRqkyc
I9fVGSTDei8TSbyyvjQKvRuLNv62y1Cw6iAjKlBsNktTv0YccbPBIOOtf0s0NbAY
oIcaVYqijkJbwbdrdj1mtN/dfcwMZLSDk3XUTZEy0L8v/DF9tYYBqqI4y1xNvcUY
/oqXrewqNOe7ab/aOHRt+PQVDLVpeLsd9ZHbem/oE4nmsCZF9HmY/qPUgVwkkZMW
7yv7WojYc9lZPDltnpn/zFtWcmSQDcSgSojDhcEckhS7yamR2JNjFxycoG9W7aDi
nZ8Ax9CDJi674Y1FLbY2dIFS9hyWON9IlmBiQI9oeVdGzyPg03EFVGAAeekNRclK
ic/yTQNvG77CGogoJpkzuRvCSrU+e10+l+XbdCTiCW0LfrnWVYdr+/cq3VK+QdXJ
IAKNPSZD4SWojX8I3FkGWgbrPggIEwzEyYzicpQu6ZTXqwiXmbCx/OXZMuryCX0T
aEeIEI/UidShMKBnS6GttZMDGmy2nYAKRVdVN+NNt6TgCS0eFJt+j8o3lyO/xDPY
hjBwYyw5SftNlyfa1JHkD98Vc/KCiDdsj+KGIFPTVz3oV+ZufNrU09ZdMCCTIqHu
tm8qJkVof+3NptX9Jryfg6Hm/p8fv1nwinQohiY+/M5Idw87Z7iUHqBxat1ccnBV
sUMHO0/sSzSEdOO+WNttD1mlc9ftLH/zgXAbO6aOsTMNqo3RPQCUuEoXP0AEOrfT
rZ7A6IgH1qa/ykhZ5M5i7PVckz3QEs+D2ME1G2ys7Z5rUdBhzeKLISxmWizH50y3
5HynS0IkNRZO5MXVyLtqGdbEgX5crPC/aNIqYcI5kZPluPwiMcPf0zZWImVDFh/F
NiH9ZoB+2DgDyLCV71rQIIdHU529c1hyW00zkU2hWVhpBrOcn+nNxzsddIYyG5Y2
XpqJOVjweBTUCzUNi6/iZ6WsaPvFS2uJCR0xKmCUlDlE1m1SjTpUhGXxiPQedtpo
9kfvLNyyXmKvtWXATNkplXKbqkWLRz8yZy8b2J+Z7yxNsbefJ/P5uCkxeMfuYW/q
z3kG+LH/VI88DvRjJfG4TvGJgA6iEPir2kE7gwBc6xXvrZmA2Avnkspy3KiRUhc8
7lRFhfIqhroIhD/LfmzLeZflFj+QKGJF0d61z/HMNr7WXwpJLR6ZuPUvofXsgHrr
CTe7FV78IKgjgTkJjAseI1V7uVd3O7xfhNRGewazLHR8g21n6bv7zxMjpOqWXlfs
rS12VLLs1nL92+tq4ish35X6V5MELwAjltV+ugyWWfdUEcgQ5eRPzdecigAroSZH
YJfxkPnFvyyfcw0fQMj4cD+zIGxc0Z9EEX2e/4RwQCrR7gIArzHwrHzCSdjgdzBm
tiEGylfMCKmnZoRO2FP1VPgG54gWhBse2NdxKdtRecH0CkZu8oegavqkiFI4HClN
JUGZlzHiMqFkyM3mf7SgjsbOzzA6qFgdOVhirVe2zyNdfX3ZzAky5Gy+8YleJjEL
RZdA8UZnmhzd8wHjrRsLCjGBDMhOcKWpi33uXnbyax3ip7Ga99/6Nauok5+orrts
EwHvA0FX5KI0GV/pckC5I3h5GIfce0nh2jvCJlw9THglA1GTFHbu9NX1+Ii+toj3
GLc7fLLN5X7BSkKxtzoL2gWMEnn7VI0MY8AUVcmYKo3lIYiiysWTRRXtppz756Zp
/VXVN9MyWZkuI/rDwjlivmZvpy9HhyniAAbzUJ23Zpp6AurUzKd6ETeinQWSJcaP
F2dVLegN39XCykv0isSU2SCsWGiUttv8wMmTJuYi5+BUVUwVb65ywFo4Lnjv3RJE
Kr8bgOVgD5YNsRwpdSva1AHObHvoQcRv7MaQinASxZm2/q1XJf6gwzbw4esDlT0h
r7BxRmrLD3O4o3Z5hf0S6z2Lb4CBYt+Dcm9zs/gCaCWLwGTRdEtplIcQfBV2muqX
H+sY3eAMkt4fPNF7XmyYmea1a8K/Ve18cU8XB2Oh1Yz6myuABiTGnxJYqAyMbrHp
dfStQ2BFr/XAxymrGNQYowY885bModmNjXvfwjfwhqhrQ+isqviFJ7xDw4Q1Eekt
y/Pm5yMV+jhf+YFutFn5aIG8qwPU1P72ocYjtEyOCcbDdNGtZn0ck9YIq01jFjLo
fgeyGPlti4IVMXKwsjNwPIBaWtv0XpRJcaQ9A51sL2qnl9+n7+kV/tdsWtwQ4lft
7bKPCfhRoOSYtKzxrYQllvVDhXqZywxeXfFgaTvRWTsd25PBfVi+7LLwJQZEOvRZ
3jt1gIWGhhj7J5/+Qt6uIbLNFejMZ34zzSpxi2GbXRw5kc31tsvlbPb2b7RomGx5
n2XGceMwNAUozQ/mw8rULNGJbpuPMkteWkQ/rb7kxxwczY3AFRWXKxI5ZUgQ/Coc
X1thZ/Mk+cTKCiIoRjgFCN0/ke+M1M6eS1IwOMrIW2GQjmjilRyRqnJL0bpzKggw
ftWaN3vXNGKODmfz/kJrPo4iGH91344YryovI3wfTAGm6vYv1jb0e1kWVIIreF41
kWtGMYjgJ5IkS07Y65hz62u2W2Ogy9M2DN5Ei1xWLPSpBJh9Itp03LAeuQAyePtM
aF3SUubxjIm1nU/GdzuVXAvWj3EabZmxv/B25Wz778bJ6Xjhc3R0NI2kMByhkcEo
6Q53I7PElQNZnt4u3TX6zPkzzJhXN49K/BQJQCSuFMpCnsJkuP8gWZZuGQtEc91O
B1gNAwwtLi5mDIcccATJhNE0MWUIMCYxNgc3ELH1Jzc+f2XjBXRuFwRrEL1KK2e+
LA7rX7s6fpHsn0tfhwvMP75wXXK5jNmApLmBk+pRWGfiJlpzCPgfn8K+QtqqmgvZ
F7zqjZejXa8MQClgug6ll01RyGwg8B5xEWe3LWIbrCNdFnwyDuFD5X6YQNyV5lHm
qyv9IDPDXzWAJQlve7uFlFsTRkEk7CveD/R9FDrWY/EIltQd5HfNDBYsvxlh4fzM
VHrr929pFx6Ss3D6ysNb1zMojGFi0FmPa2vIHvUz+vBNJWy9PCLoqV5dsvkr6OYE
FpsrPQtA+rwrV+tndsnxnk0VVKtItvaeavbs8TWFDrVh7FV7SBosf1dAuHAuaOVw
OXIXFlUZ79ikwAqEXGYQRbzv3p83512m7o+6FAfW/1K6DsDfSviTiwQBbh2oVbjc
uahq1Q0Vi442hhwlWo9X2rAD5FGpyV0vykgQpaNHqJX1di7K2bpzjvfxx8UvpGbH
T5dCIFNzirVNT49iYT80nancP0IReloA78qDBme5w9F2DIfTnhmqLY+Jc5EwOjEX
Ovq8wCGIsaf5xJOv2ChfeQDbXlOyCYnulvithsfredyxBXlh7px+mF5PLqyxTMyh
DGfnZRF4LjMs60wbr9QcKYDQ58ZCMiDWMtH5/LPicquRIVptLNAImuP+F/F7wWA6
DqXROASTMkrrbZKx8xGZbZbrsJdPeMidKKC+sH4YiEeN6U4h0yaa3G5SmCrHCp+g
e4Uv0mQthLV+0XeQtVx7K+4bdJ8x8CGvHsm04CSnVxwgqMgli2M8a36yPmZkqJ/m
65rCeUzgobSAlWemapuyRBSjyRxJcWgfOYEDjzQtQt4mWp4VcdCEQAyzTSkHj9wM
LBpUiVUh8BOKjiznQoqFv5ftRuWkFrI7jhLrYAyil0+Yt5OMTKZ1t+ZIDub8jx7o
rW5bRi9ZnDgrP/VKyo7uf1du8RcKPQNuNww2aq6DihacPzwLy2cB0/2/EzJyEHYA
YXa6XpGiE/OUT3O6XM2+LKGExbLTJ2sblbRVXe+NV/4+TmT7xPdyDghQdriLX3iN
Gc0qFCrblQoncmZOB6pNaJDy4GD8EfW4A+QyEy2jr1m0+0C4hI5mAx0bXtBrPk3w
1KqWz5AUlXFGOKXMcb97gghmAGbdEZuTF8uS0TDnF6QNVGElv6C9NekXkWz4xU5o
xAac4uu+O7htqRcT7RIQ9O1nqy9Edx1HOVBxpS6YHQQOzRaOlKBsqrK8/suVJwqB
bX6dB/afqIpHdu5sDCDpb5T93VUPEI8peWFlvOgfy9JKfO3Ma27qkKLtjWFKKkyN
pt9tZOgC/abbob5kAMPfw1HdY2nK44Oximm5BUBf7/2w/SuoGKWu7yrTFelu/qtt
hBH8FtQ/DezyaSII9qNAJn6q/pt4g9rkwgxciIBwNod7O3BrtcM7EDVJpI7945YA
kLFcy33uPT9R7wGo9OZLBQtvDJ5wqx6uzya47//GcK6EraOz42pqepIixxilNurD
YMDHn/v+32uS6BLcqxj1ttlPjPbl+Qx6lw88/GNV9xWVZ9fIaOmd+H0+fw4jUqwN
Vzf/e7HVyN2Do23xlXbtqdkUNUvyEzvmLP+fbJjkf9d0hK/s3xFM3S7hiEXuzL/O
q1Xp8ANka0tt3wNaW8HgXDcCbLLV3uE/e26iQiws+LTPQqedqqCceMwvzqDY4ntL
L1OOZnEld9tKiluRm+O6BE/CCv+lC5MOdb9eGbWBfHzo8SJichsmIiHpUhoO/B2m
+47Y72ZEugixoP2V36+n9S3F04l/ASLcLeEpO3apcRvaJwKqNMGgtMxp+iqi25rz
eT3Nr6cbaO+EXE5KcB/6FZ7L8YyZHoh0Mz8CflW0/ftfp2myaIoAQmqeRnHHCaVL
0sxxI0qZCQM4NhdTMLS2evxYqZcmM4nIdd6tHi9vDKdzqwrPFJywgqKJ11vCstb0
e52jc6wn17czNkVBLeyrt6hO6+O2X/iFqw37XHsnZMIYjra/j5iCMFvKklvW8rhb
CaihIKRlOa9slLoAWeNChGmBtHhLlgoVptnjb3pfX/pgl7ilXjTutPkGGzB5PNTM
ibE2FAnuqI6DA8YbNE6+XKvFL/8URPHvm2z/CsmKP0UhoDh/LIB5tMV+oFg3yDLd
MfqZGpVKEThwA+ITMfvcLv7uhBhqAJKVBNY5LprkeziSebMxPJcfNT+5k7Snvvpg
j96ha6yp2VR0EkdQhOGbSLj1pon2ElzzTU4wHX8bVlluAn6eKBpECnMF+f9K8cvc
sAFO6NfUGdojGg8lSjsaiyVZ346Ri4x3utkZLbm3He2FV4wxesCnv5Wfmmazj65r
ubf/472jSs8VZah7DUIWt3NIK1P2i38I62I9ryHS5MFiAswa1wGn7SunOiJ4aY0r
1tHsmloXHTcHCb8CwjY3CcpntKrXNkdR4nxKJfoYkvrFmqPGTmkNctNbFMD/B68n
NfJ2DqZiQqiGbVxZgFsB7J6vOIoSrBOBgt9ST+iEUWo5P5GVnF5fhaKJczo/eirO
/eIR0E0KBYMJyZQ1PHqm+xS3HxUi5AXLeHiR/8viI/5Qc9GsERUYuPFMYF6RYbS2
ZqTV+BYxzamMjWoJWf257UxtfHFYp3Abg+BvbDbTlmQSp8IqcFyLoZ0b3uI+6SId
iH0+OLmEd+dS9b/iceteqGISVBsvf8VwvWIaoxGsnYX296D7g1yd0ROcf894xpLr
QbZiUZOrCaNrGkN7v6ppu2KbD0e3Lj2dsEG9Tr8d+SbBzYW00vR3U6dKEDT5/bAg
DlG22R49sgjwf6g/RuQJfQ==
`protect END_PROTECTED
