`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNJtOAFSu2W3q+d1U0xvIBqRBp67cLLfk0NBXc4rTRVu
wAz8tS3MqTES+LW/LJM1V/yEb/SLTM0cdWko2fULsp3H51EeeLECs5su/Ft7txQh
TWHgGnuTloJJ49wI7i/poKfpBQ84oE++hAuPByOcnOhzLjw8Y7IouMhpm3m7mwvp
/hDnr/HK7KR4Y9Hs6i5C/QCq/bXqpW2k+4PJb4LPAsaXBKhEZS5mEBPDPpuS+8Hv
3KdKgPFWA8oYkN/NMyrsvb0FcTGVQadbZKZlGsJl6PsqdcuWy/Ay0qWszNI9EVu5
mDu8PYt6guZP801kP0cVwrumhg+IQyYtfjY4z7IGSdzcE5vjzVUQve+dm15AFERS
VLuNfjMaH2Aw8yvPBt6QtW5MM8xlp4qcIaNyIaQ1d3CjvrcxnbuhelzzRdeKMuY2
uZLz8pxcGsbg4wB8XkwhpszPMdJe8xLLfOEnKHdWJPk98gqDKwTllmkiDFREbCr5
srvoR8kQ9DRSzFL6XYD2/4fqTlC7WaSxQCCdXQRSr4j6ewXqSWDWtDtIrABD/TjL
9F5LQvX7wrxaweHeAbdfJQamuo2LLKaPxGYMKtzBdv1MNnWxFfYeJUiOLtuBTdwq
VZKo5sMxrlX4vSW64WF31BPi3r2dxYsN81x/6IsaLSPKtekM6ibUcvdAQGEmN2ga
xnk8vbYxaqYU1PlmexG0XAOqr/ULVoqGosi+s4jz3UIB5wx2zzFELEGcOcHpxu3T
y/IEFCKjVGQpqAEG1JpJrtytZooqrYojo53rwwJA5AG7ej/JRuFCKD+pdUuVLNqI
`protect END_PROTECTED
