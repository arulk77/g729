`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAd61+5q+6NG9Kpdfj4V5mwo9VmW+qQqfMIvMju2w5POH
wNgYLhGPdpGS3PzIEe/xJB3mCa1j+4bYTouUV/9p9EOPQv/JWYWygjf+oPuLXL98
WWl+RjNzHYEz3yeUBPe9R3dH2LIBeVVPWP+7+Mdpn3D8zhE7ovQIDNcqCUzIqayE
vV0Ff1YYR+6M9Vrliea9BpcMzaD2qsfNutliZyQGsXyj9pL7LusLU8y71iVY6hIe
hYW0X76JfgcvQYqRNS9WtBtmNdGr5IPu7YX4SJPB0+Eq7huQNJ9/fz9zwWjr5naH
8+kvsQOKz8FfdZHvPYhLM+Dhp5czfVn2SDxgCp/ISsOKV9aBXJrAcWjc9yRKQK/+
dKUAKbBrf8WGwbt6Z9ALI5MdG8urKDiwfwmOP/8ROgahMjRFg/4yDcMmwbfiFgqS
32H0mmFZiu3vlV8jf7RKNtJ7oyBcjbkNgErldNI8B6lvKKHaBKIgEE9beiAPmzvc
4oTMHIG4yFFD0vz9I+Cjnc5w6LwQVhqEY/IxtA6hS+Y/dJtv2nfS0TmLm3p/Jrml
LgyJWZm+GO3qJruS9M1Ovudb1XLK5zJCfAokIJjji4TmhaTgR8LbAML2ZjnC5ntY
4c9gHhPuVqRNittaCOYNqO2p2QcfC4YQfTLC/u0syr8zbA1K4ZvbG7v5R1HmezB8
ydbdb+BcoM6MHxA9zzzwA5ByDVS3qiTv17WLVj4rUswpmr2S8oC3FOqVF8xSA1MO
46LGwoQSjQjw1IZ/XCD6RA2B7zNgD7ATC+d7KPGAGst/ej8uQCBRE7BRJmFUbpRR
hpmFqg4vOisuTx4ZYZqdvq7p4Xl3UruKHg0P987MZxOJRtWGiDokaPOC+uxZIAra
QXr5aPU3I7YXUvzoSJaByhQLhEJm+aTWhhVYv6AxUra+I4cpS5vSfOKgJ/JUv+64
2kQSK0BGeX5zScxCXSvqxirQ3CxKa8t6LjS6l2MTrkIH/WdZLH3xl2851eKJYP6R
u+SJDmVs+CKOzevInAtUJZFiCC3CfnL0+cSpeEKuSAMDEXUtJKYhPrA13ljHM3Fj
KGfO92ys/Ad8z6yGqSFKXAdKUKIGKFO4y2i7EfgqK8U5vK2KkrnkJZCUvzsZYfu/
OjDJnHbGtEjlE1o6585z11BMHKpZBnQtLiRj96fw6ZgNlwzrE4ZnV+mQoIAo3336
pTgWw1bXli2EPSFbRAXlhAfZWhzxEuhXRuyCMqyn0qXSDXzePgT7IwrtFGNw8wMj
TSh46ajgbyM++WdKV9m+AzqJ9DMh7GLGUhVKnF3yt0CRA8b6BULe7pC4IcZCPdv6
WmlMTL+6LrIRixxd2MIkFP8IcupJBJEGywpCU542j8lJjgfcv19E7rBc8xmzQOmD
8IenHKX42hXe2rhpApPQyppr5eNmpI2TfYM1HdtpXAbZCxLae7R75ckEAYd8LRtu
611+fAZ5R+rWuA8gSqKDATKsw7VaanNcYkPCegAUF0MImb7lXtTt0jKmRLHwX2sZ
rYmWhHfyRrwcicYMGYPr7cYG4RyWQESh1gSJjHU2dh0epEj91KTIwGfHK8hU2gLv
zyWOpo5MULftJw7hbFQUZWrNGNL6gc414bd44vx+falttfSNw2XgCDCwV5YSWeuL
CVHMZBsUhrjEwoBmJT00nOI//zWLQmRqoO9vNu7wgsiM7n7rNATdSsQ79KijvYKR
nnsdXMWWKGNjfvMklksmCDld6znqVIkZueGvQjgRQ/TlwjtYH7v35utm1ERIFkxS
aNahluOyOIwUHYhQy161mM/eyHoWxDWR4aCzaZEpf9b2rBA6N0o6CdJ1lBnxo9cN
INnHhdLkIWfv4GBA0gsC6tVe2dzxYbLEv90bm+YpkwrP+j7FBPNqacOM6tKn7xVt
5sObruQYQI24ILSH5A4B/UJf1mT+SDC00wYknP+1jaxS7o2PWs/Z8YP84bK+CY7G
FrA7eJnTmFtlHN7Um0xuBo4KtBq4SnHghUZx/vK+kWFqCX7P3yb+GlVWoWQquPR3
FURBCYd9Z/LQZJ0+GI0kSOvwFyszac7qhW/sUEtokyiPUgoD/ysjpQeFak8hzqiy
dQpXsKDYDx3FKZptFIkUVScW3lfG+/izj74NArUp5omgVntfiR4ev4i4F6HO6423
Gk+0sY+iF3eX1IZgKQ30L7EOMocN6nVTPf/0pBKtgL1QpEReGByECclWozjQVEA2
i7m7qX+Z9xxBt8K3ZZ09+/dPf10pIlUVHWghzgDfug+hgqFCzB4Xiyb5RUBErS5W
bMQPfN/JfO9yoTaH2miuvbMQz8CyobBHJKfPZ1aDccUC2tuELT18XiaVV4OdsicN
ddjxLI2FT+cvgornXgVakvSo7R/FT3BNdngwDHU0zj2X6zNG0bck22PL1v1lvwwS
1LuXyV+twfuaCwLUzCwLNJZlRcxoMs75JtplqJ6m21uSMzPTzLJT7oNXzi9Bl2If
4431wYQ4bizarQSCRMGDPEKcQh78EZwzKceByqV3VcmeYUJO6mZOqTuVXpFhxH0Y
FeIjl2oWZpzo8aP6jRaBqUZKNFPTuVoBFFaVtHgnGPwXJP28LHjFE23VqrsSPKz5
Fo+MfNcthlcpNZdNEexZcWIHhzXyZTqlq0dn9BW3QZBnhPp43YSw8ZGoJantCtEO
livCsO70daPZ0ohlZ7Yi5A/mOMLcSWD4j6PrS9tOAh36qfsgnYIfUc2ZhW2lfPtM
19u8Rgmhev3cXI6K/kSyYAmU+MddldrDORPRoLQxDjd54qIP8uCRPmdUa4FdOoz9
ev7Rh8INFO+jDUtyAXdChWzUr1czDfcLSGrUiFWo+8CBLu1HYoiTkVw07Bnlvx31
PR3Fs4rFFCOf5eoD48hueJzL1SMw4ehBJT1gAufO8rPmOEoQc/l6CE1hciufbokp
zH+yMT0OLqvPaiwPovMCcwmMJxfl02gT+rU06xBwF9SyqE1hGXhKKzdreOcCIsG5
4bdKbmdW+K//Aa7jwGTVayqaVaoL53i/OD3fG8GuYWlJP8lzKDIjJzKJas3zgOpL
f+AUxl4QGeO8inYEteVEVQtP3MU4MJQDZmcats6ltrLzZ6BQah6+MKZFUkxF7kjy
Xxd4Z7xhy/WQ92ohua9itUXKjr6nhmRJ6WCo3t0wL6mgsf2xZuKeLAt4gsAlBk/1
h31In7QxmZiN96yYCM7ocPmTN9JiX/LUZZp/JAg6WRqEI0huq7KdSuRtE3nBTxNU
40ATuLh6+L3R6N13jkCGb8Jis7MNHGMTk05ZL3l6ba4F38GFAQsLYsTMLrAtinli
k9ae7iQt3cDAHQ30BndWAFOKlAXR4jSPvCL9ChL/jyoziqFscJtja+1Rtr/wr097
I5T5TkeLPj7e2EwPDYiqQ44UloUuYlOaSQWz8KP+IrVTHHNL9nK2NTJEuRuMBmGs
35JcGrOWplmsYbUx1F/PikEHbJoXb9pABbC5Mnf6TksYy4ylbacDvL8YjKaeVCAR
b6oFLRjtd6dVqhmA1wfmXPA+NNt3gM5ppgyhJRADmy2y0b4NRbMcLtQiTUz34DsX
iVnCiAhvsNom3l4g6lu8muq/Uw70IoQEhyDPTDXFeizKGdCgr1lsRJhND6LhN9+/
uGhxUTrSF1Rs80GHpbIrXhYmCxs1732VUlUnxe8FS1CeNihxg4VPdCccRzia9E2C
bVkNLw3xm0xkofxunlHZpHOK+47+0ygmBwaFkv/+imvoC71nDKnbtFuN+tdG5Ur9
q9spUy0oOr9Bw+x0ZRk5nCmmwz2/2AM4FLB5pX/eX74ZrI8B1mZ8ziMVn8KSghHz
frkyBSAlUMm7AFztgLnpZuw7+Jy2D8N9F763Lmu8tYWqRYfnx/tOlt8xYJonD9ml
/NtOPHecPTakzyAOskfNa5OQGZU5L+8Uo952p637h8IawHUgpaQHX8oasxbGtw17
/UlbQI8pTO1wSF+CCdHsXbMLjMbpjo4IIYgjYjtg0cEsLXBtWRHZgqla1QptQH2U
Mj6wPYwe9XKYlbNRjkZhsqfeLtFA3cCuWrb4CJpacCG5xM4Pfm5aGYhpB8QXQz6D
LIIUIE8XtRc1+0aBNP6UdZzYwNs6qtoyDicLQ9kisEuDnGWWBMPlnM2XdU9AlBYp
ySLiQbkck9ApF86xg2Qt9mWjdP5y57rHHwcCB6cYEZdZB8NLGbXlBDONJP9GJr+U
EFofld1k7bMbQ135BsyP13ZlzKsGuR1jsPJ77d+gK0vrLqKZXFX2FiVhBe6I+ddg
BGVsDcjV4fNh2QIpe6X+6eDg1p3ZHF/Jlg6RU068VUh060Bou2HSFSyj+v4gGl31
wFyHCpmIiF7WKm4FymyqTiVLJ1T46YymvOuE6H8kUEMFr963yFnYsbIVfoMhTIDL
hjp/w830Ona2+vBwswXzPpOMXzOUIuqEH0xl6SEv/CFhnKPGvrdtzfqcmerOpHdG
wuF0WQsZxV6Q81JMZxytVj7AKI10KEQFhpkYLlJH6TT+X/fNqtEBzIXcUcIwWI9e
AQ+rw5oilQ19aSK9abrtxfDEMKQnKi5w11voNt6zBcM+u45tnlP68j3BGiWrC6Zg
xq1AXE1+bQyiDIdOGPqQmaSfXau4XUv9DIm1Ll13F5jSePOMpEYiIFPUrb6WNt7i
gnG7NzE8l3kgiv8pDBQCGVhNdEnzx9vPxZZrF2RGpY7Tw/nmNBByww9gwqAgjfWf
2EkVCrBYC4Ci+rk7rFaqsBGgpehLigc49qv6oEKDz4eAjpd0PHQEgEaXNzzNNHNr
946jgtkD0TO9umXOPb6epkBrnwa3v+b8OyZMLB9ikVturp8FMPPndTiSh5wHaMow
ZAq960t91RujhSZ9gtIgPxDtpmAc7ExTjDqO1AqLvaW6Vc8FkZic+0gdYU32/f+A
RM9LrIiqeti2mMTYD8lW/lAZkn73cUP921VYiQhrg/FEAfxbRmZIGXoGUKibRjLw
RPqNfFRYTV5IuHUJdprFerCDCdQSDXoMmbol0aAeCSPYbsL4N6hpsfUxQKzlk85z
MhDsgTK/VAR9edMZLmiB8Pd1Z6x/6yKtWbwQ05n4LZQ2cRpre4JDMxnd6wReJUUK
ZvmlSDrPTEHgnyP7yVDckO/X3RCRwfiYgAwlYtixtoLxCbXlQ18sNpCJr7thJUx3
ekD+G5+tudyAylrBx0Ob8iCMjuHnB5CAKhR4XAPdwIGFPeTN11qf5dM3iQhjCIYY
gKq7FVCygNhANAr3+UPcL9EdfpOa86tS4UqWYYgIrlMA32hk8C3qrS5UmqP6m2A3
kwrGxE5b5l0TMBaZs6KTr44w9+eJ1cZBdp50oL83IzWt8MmjCOcUV2glZLixxYf+
dSKre+Tl0I23RhiM8nvyopphrYNoMyd3zXB7dMAhyTnJgwzMnis3zpXcSPxj0YNK
aGAxaSGdku0daKppF5mW9Wl41MTK2jW6RwmTvkzflKfSjVaYrdn+2QCnPYGBy4Ee
lnKm+PjhAG191rwwEDP2FBHDV4FxbaWfLUjlz49+NHoaXrs+h+RnGrZelKLeQ+Nw
ASBqJwDYXQgKrIYpDfY6d+cMJGq5vS4E8LOw/AXjYZx9M5MzZa3dpuwv4zE0ShOz
2f6BE4rV1safZ8rT+ic0Nd1TejP717EKl61i+R18qi9LO/xEkKRY6+6QBcmFI380
c7VaaIIzgqKEwu3rlJ33P/hrw+sw7qySSQFN1FO+t1Y=
`protect END_PROTECTED
