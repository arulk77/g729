`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDrXNDxofmOCL27hZ9c6+ggy5769bPKUsq0oFFB8jNLe
oyjFSk5aiaCB/v1zgRxW0Y8BDupSq6KgL1PxLmLueMNOk31xlqB8636/sZOPzdKJ
E6VtqqkQGgQ95TlYmFAQujJyGH+XDQ5XBJBo46oPdex39etnZkS7bn2DdyLgtffD
yVzl1Olgtc+b5gkXH0i4DpLpgOgP1iZWXu3w9/GZsXji5AD9DUgWj5zlRq1yGfRZ
BueccmjO+Nfs3NqauWZY6CF3oZAfvV1S/P8gGEWAHnI7M0JtOe7nLrJ2jXxVs6JZ
lAi5PEo+pHog7OBNU3FHXA==
`protect END_PROTECTED
