`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2EBoZu9tBf8wFLCnm6xiM+jmsEaCkkJgN/rvMPycesCJPlS4kXCvI5gVIBLdezik
u7ROOHk7dcFCAQUoffoVX1p//715NT4V1a0NzG3S5eifctH2gqMBOY9qRUyuHBGR
DECTrgKP7+hnG4/7eIEekF+ZnZmFU7K1zkoWqLLyfossuUShNKt/Ndn/lgLQFS5J
9mIYQQjp0jeMsDtzCERztMz+nOwI7IUf1yRvnSD+4KuOsykwJsTdqK5DcvQcCEMd
/GosAmzCwcSJlHAYXS5Qgd3FxlYsk0zWC7XglpHnPZOY1ShUCswKOW/zopQFOcl2
`protect END_PROTECTED
