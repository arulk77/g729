`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEISU62koiNUJBkAwQ2oAiTsTdb7ryY13XZtDQbX0k/W
q24t9zFOBtcR7TWEQqc29GQQ8HJQjKwOpmHisJOwejd53G8+zduKqs47DbxkBUct
y6L2Ht9h+wbsVilUq3OdWDRy2hSE9k853JdTpjIWpC9llnUJv8JHU9ncEzJCUYtB
S0Wbd/7WwthqIcsCU/p4bZ8iLxR1bJKNyF0CjQRTe85vxd83UvMJ167ZPrVOHQgO
lsGLBBaGY+Ysew/GJzZLJGVBABXzbuhPtt7DAYHJYCGQjGOu4Ml5XocnwAsqSiRB
C+wohBqx/WXaZI0dQw199rSXU0EEmKZbfiU7Rmb5mZv7CRIKdqXAlC6rob3+qrQy
mAX9f6ojZ8/xahLzWesfoA==
`protect END_PROTECTED
