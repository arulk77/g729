`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ZAaJ7QzJ6woicFnQfAn5xTchXaPXaweIQrWEXgaQ3+UkyK71gW8kQeVOZhDpnEvo
sZXyL+Rlk+VxNhWkLHJlPzj8syCLwLMINqVBvfLRMkE3mTAm/yqThKn5CKnCxh5n
tyj+70sBKzYtt4Kxnwm0wyoUhPeCo39+oxN9dBl0S1ajm0ulnkawBsyDLbVO6ijz
raeFDNUNRJR3Jt1SmIn3ohhj6lhxCyihNyCNgeLJLbLfCBuAJqvkthSC95HkQb/E
U89xbUwsV4/RT7ZDUIjMKsMcZFu4FIU5VsRWwJfd6ww=
`protect END_PROTECTED
