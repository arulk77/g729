`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C6EJBx5J5JF1Om09ZazeWfabPPylF/d+1108IleP9A21
7qw+eW4Sl1NWRAEUR6B4UTVtN8bgZjkIqrmqHzQtL/ihuhMXhgNhC3mY6GlgjRxv
VIWg+xg799JuwmYRMsAYO+QrlFMnR0OunF/zWM4GYv5jbmePj83VKqwUDwN+vRjB
8VTmPvEjF8eva9HPbsT7Jb5+/RBqRnf3yVYdSvRNSkmfeieJBCZKPXXrvhjWeuC9
bR9obNdLOf0zEj7vhVQjNf7wKRnf3wFpvF8cgf2adMJaRUo6uNkb/FfKynQZkB5p
CbeFOFnRP75XxZfC/dA7nL2+kb/Tk12mhrUn85Or3gntbTnzxyzxKGXpPKdYPeTn
8woV+cakXQQkf+t9uLGHvsAbj7fMwdHkaFbB8+KhEoV/s6TKiN5njDcQCDqzJXH8
0IkNCqo1N55SQEEhFXVA7I/RpChEBh0PGqHE85rPLMJ+It5gN7o+AesNCJhc3ngm
uHlGJT7/LNdN0b11Dho6Ry00fciUD66fOEVbw6SeTxW1z6H3zuQILZxepny7mcHB
PhzTnGrtC3pg8qBRzrt1pJlazpl/cd5diZf+5Nae+pAddpLgBSxWxGJW6+6x9Ob8
BuSK3cl7s4v40av2bAqeMHUmXbqgd4uq8DRk5FDxGdHI7hr2+88hyhPmgHOjLJEI
/RSZKITwkTT68gOgsHbe5/rt19v1wD0qGGMDGaJuMo6/suYtv9LIXWWRQGk4kPuI
O6g2+ZIeCNU/E36h4b7u2cvJN3xKm0IfU1pfNKmoZws06DtvZvuvSsCCHLUAHB79
Vpw4nBxcdb/fOXmKM0Z5bXQ5NR4SqzB2ooXZ24mexOr2ZmbM8/xQ1QSQUjcKLac+
1DkOnssWiPxi3HS60k+VApnCS5+Kn/omlRHfYOLRDnhnEtHfg/fn+5M+QGK48u+O
eAeAsshMOAvzoxCNV013cBTFDuAB8PWNtNgLmTXSzSFjfL+1TniL+jFbHqcsVApb
0IefA7lbA7My00hfZaqbkNgsOMtN/dfP+vG7kvip2nS0JWVbaXETZJzkDmLTvAGk
oYpsbvucgPvk1Vtq8iePflalJ5ifozJvnyEicPvkg7HQ4jmrgVoKqjcar5MvRaoU
k0tJNu6TfytrTL5b9PFyGfAT2jpAKupPHrxP2/2lBN7v5GzveivnJU9gdeiS2Hbk
JhIeQxgYuAVrja7BF1UsYsR3/qC7+IGGvTZ2Qq1q877SW0BOod8OJX/WcpOBNVBX
mQ0L+CBvRwHKPD/EZIqF1QsiyHQEjy0J8C/X/U+7irSkX4IwQORPQX566GVE1FXf
Lqy7sFbGWBvDYcF7gpsmi6nYNp9XlQex3Sz/MRmRBYbJtV9BYxxKP4vuUbKA03sf
Ca0MFCdjX9F+bwM+rOwfaYhvn6mhNKulJ1uIiLy4jACwBAlJrMmLWGLtLHOK3oYc
3QZzPs2tDanNGEWj+5/RbxVmEvsP2xAabxUnbKIvz4qbw4E90Yj9y6QEZqbr4uFu
IbjgP+5VjPOwaXXI+Hox2wP82cOtDTUhphXcGlwcno4hR/YScTcGiE2S7W7RT2Rd
VrTjvIXYId3ltIDBJfRWgP4gHDSNDSGgeLfvrGb/oBsXtMtcdXUQmFeyYS8xmZzS
2UA52WareC+RQfzhpsOcEQ==
`protect END_PROTECTED
