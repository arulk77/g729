`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
hqVnk55XAzNkkP0fK2hROZaTy5KG81S7cZZRib4AHASgdE+70VAN9UNOIvl/j3Qn
cUtYx5yxVFBfZdK5TjFRViF7NAwGQpwCEsfJDGI907BCZQMJI49RhslkI0GUgCEw
/3Ph4d0E7raksKR/G3f6ZPcaKd8shLDPE7EK4fr76//IjBMdcnP+OeKJCj3gM4As
xk/r1LMZEJ9xMk9VS4ZkWdSs7wzkOdxEYZXhMWd8igsxdEOU09sL3cSQUgZqZvya
6tUHTi9BDIfCeLD3s4RiwRghCgJkUImoTBgf7XM3jJhaYbWRPGb8XYjH2lGoSx0s
89M11tlO8WSmd6kXp/xRgnyScZUlJgTaa3x1a/535RNRJvDCbYqc0HjJ8DAAUPI4
LhcsNnzh7CLYgzJ0rH+MfRxCI1uDQXCXCweHnYjD7JMrLEmqKc30xsqyXDV/xNOO
1XAU7KUF/x+NxtBUHC/LuKJqw66xlfkKziO79DZLT7xKLvlCnmTtSW3udzWxJwta
Sf6ayzQvVPinmvIfPM4edP6jFidBDBwhsxr9RkuI42SRaeTfH3TDtbJJoZeUFLex
a07wBL83ytcOEdpaZk1FbEZqy0dQyq8xBfHsAljkIM1f2KAaiAUFbmrLWDadHEjf
InEUJoGttD1Q4zAFvj7e0rnCewFOoXFDiUM9enYTikyBth8UhEfuHQKtXP/RWiK4
FkQkweO1kyuCZkyYMPBoUBMiFXVCplpvFAfu8exOZTBH9GqgmNts0hPNxZ779a+i
BC7fIsy9rq7MYO23P+BP/MLoYQt+TujH+eLKFjyJayFj5Rk+9UIZiM1Jz0ZY0nqy
CpbWeoOwggTWGPCMbBYEyntKgVhokCbCrX/4R9HRAZ7o2vog42KGHl2s3hD4Upe6
sFCBjYlo50cWQMxEhfUgJp4Ur2ebCSDv7AqDBtROhC3YbBbZ2GpPxAUHJpzqUpRM
UIeQ7Ujmcc8m8kNBvCglFEGdBCmYLFeqxiECKk+PFMFZwKtHxkUe4c5PpoazZedD
3fqF/RAGgxUFTdRFogWcMkeol1ePSOqYirCiQEIeOUj7K84GbOaXJdjrJgNIDRm5
BqkrZXaLLfzSMuhAme16ChRFp/hNN7PlSeCZesnu+1GyDxjNr9ig78Rqk3v6naG3
vJs3QALHIUr8/4dJEOnRWNVkF3ml79apPxoNZjpKo/Kh4+KMc83Nq0sEjDgv5sQs
2UTYTFI8C4gxQYBwqTkAa85gqTUS+ozGlsCGHgpkjwGzYwL47cKUzNQi1xrccycI
teGMNXxHZtd1lwYYuKd3rkn+XWlQ1ikWjwTRQrURa5BfqHy3H/1d4/KTShtMEmr+
Y4iLZ1VZDZCWWPHP1TbChteqz+4tS0nIlc5hNzmmK82i/4BZfR1FfIAIR06cjqSk
rPgIIt5d9NAJuLxHVYFrBxjhNjo4Mdni9KTVSnt3kAxl4Dud4h7y11CGa4xSQFSA
kr8fNdyqcafDKvPFq3PIiq+DUCccB1MFlse0gufCkcGED0dJl8uzhM0F1YpSgeFi
ohL1uLYxysoZcBYFd8lbHgadeF+6CwJ8FHYgAWGqJloxWS22czFQM1gGptX4UwNu
azf3NnD9f144zdK4GUOWOeJymPuECZ/LLkH4zmEDN55tfDUJnpA1qwMtZfp0n/bT
WZvZh8PeQ5k1dP7cule2+Wv3jm0xBSvwDlgLFv1k3G8/VC37a/GxFKFNXOQiCT6Y
7gkbeZ6VIs2x23wVTWjaWsB9LJwFyVMzH/3BlLHSf2vBd25AXCoq14yYHN6PozhU
G5cvu342InX7PBhlSigte6cCh+Rua2Lpd6vutYAdLjgdQQNHLEm5ovXwHPbb00I4
`protect END_PROTECTED
