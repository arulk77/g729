`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
HKVMKNqUPZ9cMwzku2iUG17qBAl+kT/TM/2+dGpq4dVIqRpvZdrP5x0l7i7AxThB
c+DqTLfy0Q3QVTMa/L5ajSec4dyzouChgoSGjHM0thlHV1Z6inhN0m9Ub7Y+ZVnk
yADbX9eG58pECs+KJ8KL1IG1ZbPXMUmuPaF25Pwr3sY09Ko3c2dFkpgtkpdaYtqV
5+5UD2ET2XzU/sMh+tWyj4mzPKRGWw2Ahv4oQP1TsGk0GP9i0OtMbjmmKGQIyJ0K
rcUPtoVP/y+THT0v1XNZAfTtjtaxT5gvXWRYfLWdn0YAkGX3iqAYNfaN9XobX6Ny
P54mYAl8DToMzVqhm38w0U9X7VCdSIxeJbZpjDE9qnMfNZwkqpFoJuQp+BqRSiJA
VkySUhkg6Ia++ExfPdV7gdSdJh+TfXa71AKwU/9wpXE=
`protect END_PROTECTED
