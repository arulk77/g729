`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C5PpxKZgAZA4n5/jizBQJHfzN46hcPbxOZ0Xni5RJV7x
HHKjc5AJ9Z3bw+kRxIpIHC89GTVp1v21dQr4Zx6d1VMEKw2tFimeKUNTYA9DdzF5
rnvFid+FG/mdhzRMG7grWjCAtDweWIgC4Z93HrFmGcLgYwmFqEwG/6jSOWwlI8cJ
Ne97wiULV+kGHlHQrCoTajrZgLKCNwLxk/6O8D6xW9agnuAT0wo+7NMYOgfLXo6N
lbD++GeohsqICZyFb5co1BB/k5EWcuS8ahOkU/DXi+pmN/C/ipjsee5ws/Rkg8c1
NQOue4rNKloRlFABjp0VvhY1EisMQwgO+zrxpRdW9cgmAOWKJf/0sp1Gs/gptOpr
Xe1pFWJylGMoyoUz1AJscvb2xyBmS+xsPKcsgRtqRUN1cfQsqUMwdItCVTc0UZnA
x3VWj/u5lvkZN68dDLnuMJDmIWh6V90yPE3DkrQi3WKI32FIirTAbpCGWZS1istD
WLiVmS72FKvzkYkXnXgD93L0DChWFcQc5RgLZdo4HGhhooqI1oLdIfbYSBAFeS0D
fMAdEPbU5ry+6cRi8+uYU9yVOguLlRgnifsTXA9UvHmVPJgMY54AJJSxRac6/1e3
jFvPNbA1sta2tYV7XoXTEwW2DBuXgCoBC1NsXPE2IqLdNyFsXOY7v0nfeKvbfHc8
YXWpJMRNYUCHfEod7I9DWmFcQn/T8U87L+wGwNRIu9c+9vXGEIG2EgRjLlepuH7S
wGTfvV4xsPuZ7OTkFHhZK2Oeb9SvazXz3S0x4db3uSZ+Kri+ms/u4T7LFs3DKs80
TZUfgIE7v984hqtVftJ71p206aYbSp00v8FRPVFMA9kAXyTO3+B9lbYTcJcAYZTb
5vEiT/LK5OXES4k6GeGvnzE7BlzEv3VContBFWsufXJBvtR0sMZX7FEtWps4jJ63
XAQrVBK+zkaKtbjESeF9B62DL6q5vuJsuldc/2GBLdgZDPuee37FXmslHtN419bZ
O38pBBPSfp7GhuJIj58t+jHMCBJy4CG3fEKWOL1vCiHxRkLwgkOBsHuOen2ABQeN
d1FmV4qmQaU+SbbDKW6++AlW+kD/P4Wt9AaIkCxQKgcZ8BWcAiidKTAn/yQEjVin
DAjLqllBCzLBN3eZtRLlbkC8rZ6PRsdht1SdMSaMG/8K7WqAZ4eydtug2QX1vTyx
D/e5FVXquIerB4fwUzu48ZU5FmbGdvQSzcjh6WBZ+dEgLQUQR4kbELShNo+r1Bcc
SVzXluRHSr9OfDK+dCoJkgrw9HdLD5RYOrmBHuiJ3fB6RjIBEXxCi70Ka19+zVZO
/HN0KyUoODKqwI7DD3xLDVLORs3bNiomq4LEaRh9V+jTw1N8Mm63QwRMJrSSVDeP
JczupiWlYrJo3Ibmpvbi8BHzG7hkf+xibbzt/NvzP512/XLeQtkb1QNQGNEieulG
tM+6MEGWeYnmRBoEkrg/LIhtjLlSKNQNWfU44Ji0IjJwEX8fdrbfwpieaU0XqPro
sEWx7B3NSqGFnd3TKkgzubhQOrhDdG1UNgKo1LVM0J37s6DHNb6H+lMFU8yHKDTZ
ibqm2frP2XXEHP7357Ov2L6lmJajfPG2fr2z2OLwv7VRruZokHTwvEQXf/vzBZbF
XQ6TCdkNNeOAzlGAr/6emKoI898yBlCd1HTCZSWAHALd7X4KEtApIFxPyXa5YYxX
dQ9d5F0Zo4/FDV93jh+ZidsiBHVK888nziKxf035rKQ2fjjH3apwxBkHOyKH7PCZ
k7pMETA1HlTtNNd6YLjcN1nSLL29KmdG5Fqe6j2nx7DBl/YGSX5tEntefWn66ifI
UOC/haA2heQvN/2Pu9Affi13cK4YBpuDkeTzyE8043DhVLcuD/KrmbSbBnau7qey
vVVCZ2T8afGZPnFaskEdLi5nYY5w07vHC0UNuZ4x1LUXxNPM3J7O+4ymg1QlhTyr
ijxdk5FSbOWDXrAw3Lhw0VCJNcR/BeaKHjWF+eOsow6O+73o4cLq7Ej5hGqQYn8P
Wnu3CfwO2NzGwEoLbXZyBgVFHsjzL3Y2uuYdS1Untop06gjiyA6Gor3L45SvlWqL
i24MhXVLzdpqOc873gQa4pxL3BIrOIyNxESJNmFcHMvc458r7SK/AkI7UQvKRzrb
r7KUJ9QIiqM5iuwrNrAzrgO2y4/W/qZNw/WlZUJUzo13RzbUkJ7XKeE0nZYFl7nF
ziV+XWnL04cz3ntQSM/6aceP3E7bk2l4ulJeaefZDnSaQ2p+8JNXNYAsuMiuCC9A
2/FxMcz61ksoeOpgFphwaYE1ek49JpkLaFWVq7BP2iGYZKZNKx5aZClstqhHf5Vh
CRGxB2Futl5v+cRqbRe3qo6Us3lAXX0cpcp/rprXzJUDIq8NjAT79KL5RneuDck/
IByC4FIig7cB6t47rt4Yy6NX22Rve5/KmyuxQpB8rtRw0RZkB+gUnIkYU5cvEbXh
Y3SIAz6XKmonLDYZQ8CBDHiYNkXH00ltrErT6hQ2F+jDU8uk28dHJkxpSCdMuep8
wK2FB6Q5wx6bvbTvNZF6n9X83w9N1CS57gNV2cDND9/agOAYvDjfYwGGduUBLTtc
a/CzUUnsgs5wzvJZynpFrTmouY6pFHhvYKN5DSCbwPbkQOvkvfVVRMCOnYBFhpXp
Myohn8CwVdV4fmC/rXtKGDU4qx645TcHHkMB93q2KRCfa+EknOCLMYJDzOi6oaEU
qgiZVTrsH/Rw4hTeIFpsDU44Tsh6fcRbTxHmEbr7d6qmFfrLoPihtf8kmHYLMgQb
yp8mRF9jgcB5fRbvG5pa1xxwos5LOffwmoSm0j+pCOPlMbif2US7vWKGDPxk7tLx
ZMSv+i0CTD1gR4m2ZzGS0Wr5mFrNqkjLz6BKMLlzTOzFAL4kUiyLpZ1OY3gUy6RE
phivaNHsL8OyweeS6EHjUTKT1ekbp/JAsFD+aK74LIj46p+tjEsKJSBuUW23FItP
/n01WTn5XKagkjlZORYkDxR5N/6XEI7XKyUaJHEDhtKJ0EfJlyOr2t2GKFHADhNt
PzX5qlYG18otiy8shwsh4+kzhhOmF5MzT3ehQN1EWwbTRMqaFGS/00cXTQdhw6ZV
QSw0bYIdOFTzsXg6Qqc2Lpq0iaNXdj8IpIhtO2+z44h2LkpGtGFIsRPImzjZSSMk
lwSNl6RZ6hr58+3tMZF4GA==
`protect END_PROTECTED
