`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveE3Pt7zQxe2Pm4/4cZmohxvaAjJqADJDWoEjw4BXXHL9
DM7q5K84Se4DyEOSO+vKtGN4S7qVOBCFNmbE4g4FktPRo43yzhkL1AtQw+2eWTLP
dGn5vZi3CWTS/cYpB6rKn2hAAXb5QgYMyWeNbg399xYR1pwNXTGeVYmPcOkB+Wkz
hWol/CAbdDIn5bq/z7LHGEGB1C8VcRsME02zIlUKvijP3hj86eNAzgNWEXABZMXh
f2F/z9mB1YR7Zpgb3JUC/OY6mJz12/48L2vDABmjmQ8DDXIJTuDVcpe2zVFEX8BU
QrE5TMddKuBlKbjJFRYVaY3LWn262xR5HprhJiZAzEr1qRPPhg5wtjnfkqGMsS+z
xsiQhXDZK6HJTp02B/kMbOymGSVh+Me1KKAtKlyKZ54/NPKIN0XwMf9Xdn/biDPe
qVSfhaVqWBXuHqyOxYYJ8Ltna5mdOU5GN2FrYMtiYDjE4vmkpj9AyRAOgKmHRlHH
hKKPNVfhz18sV2nwj5JAIxihxspcp7r5kgKW3gdyi35BoGJY5KkQIblgCUJJRDh+
`protect END_PROTECTED
