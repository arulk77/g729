`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SUNl1aPvpiN20BaVLTwVX6PEIwgaqepXZMTeUCFukLfe
lodznznP3DfH0lvhEsfh201WTuxyPkxfBR4pxqkEdS+23c+YMiqTOGDDUXWwOqIj
Z1z8n/PQMgYJED4xGUO5H6I6UOcv+3pbVv8UA0O/VPYiFRRC5YTxGIQBfJhZqGQA
F2fj2kG+USKKpQ2R9ZFgnXaRcaiO+isHjSxlW0rx3bxl98EvJpeEHzBIufD2feAZ
qAstF3i156SGY49SDjqAhtUIJ0o3G0xh3Cr4s1LFNqsvCqO8mq0PmIJc2WNk3t5D
mqTlaWebtTjg+bk0Ia06FRnz5Ecf/LA2xwqDrcKVuJk7PJ9bMjYAqljo/QkVslNy
JJi0yLFxWPIRubLCdWYPCjd1GVM+wEsQULIiXrU9v6hrerRHl5DZrq4CFIfE+A+3
Ed/mSP74250IHgbbsuK7C/mHrd/yMrSWwrhNrtz/mwoL+757ZYW7Vy2k41EVzDhu
1ZiEVr13fAZK9/YmfLfp/A6A7oKDbL1POKAOqoaytgO5jVZiQykzpR1G4W9wHu6i
9wPFbG3cQcoG3H5KUqj/IoXgmdoVkslJIXLdDhwaXW/lYfaygbZutcilV9qwGZeh
z7XfYL6EVkQxQb6FAT+veK4BVnZqZSuoXanTkVgTM0m+UfYjxHK16//mPTybPssE
PM0xx5ZBZzvAMc/sw6lsfNJiu/aEgel5Q3M5Sg4QGkGbTnsBEpEaqXq+fvx4VMgU
2P+jw0AbZoYeYl+GmNrRtvFjY1Bi1r6Zad53gifZ6QqID0Cqn/8ST4BmBPagWFgt
+vkloPd7ln/2ZV3L2PqdaPNLvouWgt23sq3zYxGPvH3CkTI+HQ4Du0b/o4LR53Q0
E0zTb/SmfS0ca9LyZCWWBgnQivr8odDi0GbUk3MdtdxVVmy8y0XztxebajfDGLjc
`protect END_PROTECTED
