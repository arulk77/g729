`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJyaqtMQfi3uCybH716YJb+bQSa9fJZpSmCPVKEKpEmW
xCCNU9Xz2HoCQz15AraCYimX2xB2HA0/G9DKP0OwlS7Pn9u9BSt8OHJllzpJoj9i
zQ1QqZChk/2vffVhqxG71KCTFYPSY1v1Hvm0pSRysw8t8Zu2p4u30yHj3MykMajp
siGvCyyz8DYyxQ4chEC6eq3wMLBUzSw0kRteI07OOGzI0V+VnM6YT8JDS1Ty53Dj
TCDXC2vZG5zzjucjq2XoRNX/fTMuW0zTNl9SvmvCJsJwDSGlnLAieeekPdszKrlT
47EyFPaYKYLVYCALD44V8AChQuLOAp1Hqh6m/HOeegBKvbXd4xBxfJwd4ktwdyaP
xkjxkcYxhB8GYVmPeeGlzQZbo5SrHJal+pxwSlfKtInxeLOhPNbsi+9cHniC4VCk
`protect END_PROTECTED
