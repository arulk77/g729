`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45LyOd4i3blNssq30/902s7S0Hc1QJLUDDP5nBcu/Ud4
bnf+BL7a1+lX4uz8Z2kh3LWzUO/m52LAtsMJTipKnSOneVxA5J32XWF94o7FaG/V
cMaPc7gQQie7VbAhZpgp7/MdcC8HBaP27xulEnVgBe5zvsSgzhAZ+5N4i0FbHbzG
7seMLx5xB/DZe1ofip3zKhrkUSwyzoauEa3MuywcG3JCrbX2C5eh/JSaWsQNVr/c
kHl9Qfz1mLeR/TZ9pd80DJT35nEfrvM6e3Gf1e7E3ZOQneATvQAIpQ5adTRK51dS
To3/VpGuPok4eLz74uKx3JlL/45mDzeurNtRCRsXlAQdIJYAp6Hb2u2f4+Z+MQJl
99gGAO/Np5wr//hgZ3qUaI3dao+qq+s/bXI+nHaxRhOnvvBruSxlsdldh0U9yXlL
154tIhQRnBlzF3jq983WHg==
`protect END_PROTECTED
