`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAYk4eUayZ1zl7J208hJ8MtxfI9sKZ0P6AdfhjmbElysS
jEE5hIzeeW0l6qLJmKticBJ+HlfHEI7UqWt01MQ9pyZoxmU/rOD6GoePmKJvlBr6
6hX2BSzvi5S2gdX/PThie/xxyRdz56i870ZDRD0l+62O8+bCnmZTWQPQcQ1qPc0k
Tz9DW7YWwSR3Z/7ZCxVKjC8QysGuU6hKrMOwQekU2EBDpJ05An/qGXW/RCaj+cdW
CRP1LVXpeOOCUup6RD3Xrb9UNzHJcT0gmMFuqLEyezI0purWW+vBVWMJFfh6epfI
0DuEO7myUHK9Grh14MYlaoM4fipL5q82NHT1V/vgMs8O6pAm9WrQsTWcri1Za8hG
p/4DutQnVulZqjMQTBD213bJUaH+GI6D8rX8VmF4RRw7zmeKpQGjBgCNLUMBgIGi
QsKZWsmJflJii2t6ILVmpbyqP51JppJ9iZ8ygJLIgVf6Pu2eucpcb0JZbEyTxLIZ
mLkgpq7Ciui83DvQzNxkL3rVCcxbfTNcoBB5jeQZ9mlZ9lKkDcGJCUCfHKlI1K0b
aOcArz5ujYCQYLqu8kpXgShxV8Pq1rqgxKbv4ecrGjI9SRv+uYM4no9le4LlUl+E
m9AeLbyz8qdFDobJZlRcYapl9xX5ANIdPhrbGfRuBvYMYBWEkHSfxM6/sFyU0aQz
OYCAJdImexK+Rp8vxWeDYlKkX4PvkUcfcANjZMjpvMSKW57b/2Jr1WNEs1nt66mS
oJswFJX5WTwPITs47dDwOdGYocs2C9Iu7S00f7ZtqR9OBGiYzA9ecLSvE4RhaL51
xNKeWikh5fkd2e9r7QMdkzzSNp9qgWseYKIStmApkuD8yfbxStJJG0D0TcgEwJwT
xDd07IKgk+2TvPUNF8bDDMF06a3OM/LA28nFTAIwJxIhLofEWz7M4Y2SZiGuEGcH
BZpRtG3AMCjXc0tDUu52IVH5UEPNfJMhi8NcbFCeDqPcOQ0vrJEgoTvp5UJqAN6+
YDpv8YW+TNpO3cbx3Q7Swj7Zb8BrlQ2DJzHbNg/MBjfZN/DIj6yxOHymVDxpjnae
aq59Bhb4armCGROn7JQGQlFCLwx72H2PqdPhrbzbVV22AUXxk8wqoZ4m0wRrhWvP
PXrrv7QFFO1d6c05ZkMPkZHe0xEGUgRE5o6R14OZPCjROtVcryMc/3BYUwZ/fQnk
CU/u4YeT3w2q2OXkApnm5QiWVKw1ntMa4+q0g5of0XkbcM2TIe1z/EEbhcOHmg+2
NCa0mDueIML0Onx8SBvbRj/cUFNiIALgN/pG2X2w3lCo00uDjUbqW3psz4cwTL5G
5X2OwqZt9KdazrtmcnTLpjSQ2viLqlf+1v91QgIsWl3YhcNthU/U5UuALCugBjka
xrILc2gc+suMGX5n6ETAQ+zeO6bGQ0ZX11h9S1KvxWASY4Ct8ruvn/zovOafPQXf
D327wrTT+TsN1LCh91IxTR4I526BFvxkcIykYxRtM9uXX0fao9k9yshx6kBxE90G
RrmS0b1J51uZ8sfgh4mZdq4fWjkLmQcHi+Gilf7DBX1h+aAWqn+hGcGroGX47CfW
tLz9XJreI47SVPVB8pgjC1/fVoQL5lu5a2y3/nbVTugvZfUy/IX65cOFg8Xe9QUO
ZBj8VKvvTzvSKw7KS+58PsXvOZBjQfm4igY1x5OhgwrrVtUfBfdCvGWW5+9Q1vZK
muIP1hgUHAlZoFwoRl0rGlyy3ovJbEdQ0SgNHRUszkmKkiSijDGiEsDjFhed7t3x
U6V0o7TU8Xl9FXkAaNRSACvcms25nqOQj/b44vdpvVuxvALtZJw73o3ZxzG4s9Q8
TYQIhCtxiImWsOl9phxNJqnhH/YPtY0EKrbJKYqdFHHyuh7yWHpWNf7SjcGSeasZ
94UEaFt/58VfzdurNXNaGTuU5KmDOYRniwHcnhrUCNGhT+4VTU/vtc9ax+r08ztH
rzjNCbau76qOoE/kxMxYo1bOHrJydqf830FLe1QyMa4CAjgkVVu6VDVQiqUg7qbb
T5r8LbzL+/Znv2pbeJ39CTL67fp4ITTn1P8YzybeuslB7lN/eaLIguMvtGb6bFOl
DeGXASv29sWDKIgvwCHF2mgpSYcIUtCXsVh0pj8Xt4fI3x0xOhdOlphw8+Wl34yy
QildaA2pCOWd0td2sI7uueVQbpbUBppDaHXvtnStBB8LZcOd+DV3wf5zPoRnI5Ei
IN7cor/Es61WE7u2wRYbC6/fkbrTmM3OdcH7tZzHBcO9VPd+Mu/9FSwYTJHeKREa
Z9NpykHy0i+b72tbJl3IxtdxurjuWa2+rviDNI+R1OE1IS8gEIqsj8XF3h1c2D1e
Dr9mRXyLOL/odtj7Z3bA+T7JyEc9OCg3hNtopLH89MkVt1Cjdo5kTC6x36kJfYnm
R8BEnPCHFwJbdIqUwmC0+wE8bht0rKo16zJy+q+EAfKq7XnkFrUuzsUMQgN7lODt
lXeW1OlU/DIIzv4Ml+03i9+2wczXFNO4Cw3B7q8b4tQ1wZMLTwDebcPuU8gvS+3y
Et8vqFy63A1S7JqOsqRSHALErHG61h3euTl6nJ8V+/nLY0ECpE+0WsKJKaHZzhH0
auMsfExzm0QkecORCXMHRbPlYe7U63cYknFD1BCNDjcTBZsxApzwMUhO42rd9/1b
2kKxs/GeHUBNJzqxeP79V7nH61ARSrBw4d6Pt4iEA9OWb34RCzUBl0UphYqbxjC+
UFs3rsbp8ap2SMGAgkLk+2gxlKwQMlvIEqGXA5pQtZ5fxrW3ZNqSxAcJrBAA9UJ2
beJB8Czsnb9sLYBQk8KjogIt9CIQ3ILdaMv+bn08DhNo4hReH2DUN25iMlDZmxRv
CTvLhJr2ETiuLe492YQsG+DDOtIHqAoibS5Q4mcbQPzPQAFu4dpNSewvcxWnWFZF
WeoMRp8v7yZysNKorqQ99ZGal2h4rEtfHszcG/rKM9yukjbcFS8QrX85ghX4Svx5
t7sntGO7h7rcxYkFHL0oiq5dvkA2dCQ33l1MxZt0ks5I4lPfNx3ZEEOWI2hicy+n
we2ryYWwR9bbUPY+LnP3nRI9T5QUyP0OhMI2mjVFqkU/fmwbflbH5azFzSDhCt6+
leJwicoPdBMkAJoW4ERuToBPLFFp8jXf8hh7LXPjjgL669uAkLvu/wNao2GFDvwk
mJM6/FiUJU9oNpvVmamygFwKT4cn4aQyaEn38W70G6P8mInl+H5KJbohPmDPqx59
8th5eAo/OhyNzlZzhNIgOD0jd+sWgKOxVamIm0D3mo+oxebE/OtSb631YOUvPVNQ
KqldlKHAEE386LPeaEijbAbrWCXCVVoilgSrhoGCQOcPQGC/hMeeKOWgBG/dTe4B
3JXk9PhewLRvhDcc8nGYFMha6Bb3EFyXcRy90oqFLCtc0nJK8Q18QyWFxL/De58q
0hjIf5ipxmoqOx+5a9QiwrXsNe8N6ZxgJUV9s0vrW2PWHyKwLftMX3XQ69tKz8f1
SojCZ8ZBFXwyb9wd6hwrDp/Mob+8RcjsQ3QYb98rTlB17+YQx+NOuugGrq4gzrAC
pEzog5CAYwW4IajIWIo1w4UJz0oljZk/CPM1bJzyvBTtrafwVI4sF/lt/yu+jpbA
Wz0yFyADzPCLdemyVTWdR/PsPl92GAtS168vYXUmucRVgbicbSbBA4OCxzmWoJnK
OLJXM3nQkGFc6JoKz3NPu2QAN0G0NRtsgpOTkvLeg707izUo3iieOcaEZGoJpfY1
d7GtjWgC3obja9Ntzo1kzg2uTmAvuhroHiC/z1Fq4wGbTJj6S5YeDCRJ9Prbg1CX
8m6IDQeyBTV6+unZXSbAZZuPZknjcFN++YDJNwZuB5GsB9vqL7Y8j5MNQaa1i4Ha
uTdfTTabnjCKn0bnY1ScTIpzvZlOqVctrxvO6+HU+Yv81aAfXjrhNbDNu9mPNWaB
YJpc26qGn1AtzD54K7Dl1lzb/J8+3sn3t+aEzQpQZ+otWF2T3q1QczRWfHhR13W+
63VnCrsBug7eHehSbn7mcxVYPB/jGwhNw2BO6CmNBoJe2L2h4tz4JW1NC643s+YA
f2aUPgWyqvBnKOa/owqPLYaAexzXWFehnJW48bvmlJ6p/pHR4J+/oORc4sBSB9gd
arR9YfbtWkvhGlPAF2m6VIS+p6cJ4CiJLmKs+KtaeWAkpiDk1Ye1rNMWrafqLCs3
Ew3/PifSNn1gi91oG3ePL1Dk0qxj04ihxLwg+ZY9rxCpSZJhNCqgd8vEsJoQr/Wu
aqOgqTEd09rdTmv7HUGeIMX3w2onwSx87DLuYIJ4VOCpbweohBGXRl3q6JvQ6P2F
61iT0sP7Y/s84SCmq7TAEKfbjMjVlU5DbcHqntaYrdV7dhoVnp910v5f9tjRm2Ew
pqCDuXOGmPFuqdkG9jdiKKa5xCqoQy7rxe4tO1xDbqwh2DuNE8PhOpDpuKXjyZPZ
6lm6lN+fEZAs980HDxGeNO7FUR3EHV6saW6txrGysZp5/wOp0cSggXptGTQSRa/8
C5pWEOvgCHUaHYpX6byiRlpXr91BjFpUoopzOuuUeVQLuXl5SV7Nwc/b6yA288Zz
Dbm9AyMOCmRj99/bNBAg5twQGtzHGGygWBGqRs2MLJIsdMuG+oJRx5wyTrEBKFJm
1pVPC7aVcVZabApLeFpiARCDe3nqobuzEwL7x3WTiGQnOsD/t0QjZmUqWk6dGSnc
m/BAbUmuNIGHkaP84N1//QBLQIqgTpkZewcqgWb2+F1IYasJxG7TXqU5AalEqxpt
JgeUF67durI7OiMeZA4Bl9y72xafk3AHkJHS2jf3eO09zxSmWUiZ9xqZX7HtfBdG
TZO1HTU+fBy4vBvzGtKdfZ0BBQ7bOkhqgUZyDx3Z88wm8oAVwktqV7MkxQQkNuFQ
1+Dioq+T3WvxksOpZCvpbhKj0qd5gkyWTX/OEq7Kf2tEnz59iTlSD3xMIMmMXRTG
3Q3TefoZIJxK/nhEH80sZOMIbNq8oN6bqBHpKTrMvKHSVHYeq7XES3kXnnRd9pNd
iKrZlQIS2dFAWO7f9SD+F7bWbErUz7ahB3zBDnOv/ifdTvL1HCPRNB+R0wmMs873
FPqTy7X6zLjpJ4/bM7BW4oCHUqT+bYyc3b9g+1wqpkkqHmhc6ImhKl2/T15O8f1N
g7vogPXDmdtaqHWtawAqz4Dy1jljN+E1SpVw/unN4C8r18Dsa0sBGqdKgdg1lqu/
SWtBaDAB+Fa9wCW7taua6nzGZCMSFXZovcq/Q8oukKUw1WItggOBjogFj646GFm8
5Y+AeBjAxidjUnVe8L9gWW4q+U96s/hrlNKHYdryI/AP7bila7mA/3zhhJrTRlEz
lUvO0cp+kdxa78wP+3pLz+8Hjy4eo6y3m2FbEKMvweuDHlZE/g7GSBJrUeaf/+Wv
eVsDMrgJhxMMo4cduFS/Pklq3i7jGKvvgMA9uatPrWgso1mxK8ddQI/nnYW23Fyr
rtQ/LXE+9brEmjCyXokwaPpw3t/KOGlFqplB/K8frfa3YSMASLTSWYGspK3l93Gj
v8QGGtbrOcOtSv/f/tMYvLMDbPPQkwPoQ0FRAkXkrlFGFUQz98VNKuzubYlG2Mn1
0pDc+cHbGpqnpdFx6/LU354axWqfdpTA2gRohLfQN55JR7FLbQAqS7N2Vl+O4G+B
UIccAOyTp8OmYbAo0kJdyGgSUu8v/oraXlOJZvzoIXSI+eHZbdlPqDiu1HZnX+0i
LhZwXHiRgxuJUSDiDvgjUgtOBJzI3pH5ZUis5+rxAriYRPhkn62yNzsEwyA8JL2z
ZI0kLhD09sEJjmcsESqDWBjlULvZ4wdZ7QBidHmWHpAV2Ow8RXL6X4z8IWJIoGyl
dFbU0mZtAMHefUVTQlvS7qg5Vadt1OXb/vck0Ha0bGNwkY42/gSgB0djkiMmQ4Hq
glUHLfjMI5L0vRiEVWi+neAJU4UejArRtlrP5T9dRVNkf2Z4vVEDJpLjER86uotd
CboSsBAKZmlxibca6FaWmw1Q+bE0Ct//5JQdSqZrnGxsQDvGa8nNcghDJIsj5c+L
kxxbS4mqXTXBjjmKsqApvJw8ub61Ys3k//rOLxB7S0x8xmX4js3SaR7tVER/JmIo
vwZMGgj5Pr1JwF8ONtCDn1TVs3Tmw6vB8p3KZcx68qnk+H4tVz7f05rjzxiKmegV
bIgiCb1bEne0x+rrIr7Rzh130mNsnp2ogZ3FwPcMfglrB0sfTkQDxXxrn47FSp7I
B/eeyu43qo2U7YNewHf+MTxleTN/r7s+T2qdOXfqDVg+kwtjERDvDHSpjqzUPLW7
t3xURf/8nLtXbmyeWJatVOL6rDcXkUlYnszSMkCGfqST1n/CViE13F9cvSnQOF+7
1V/EgE1vt0ss8CLEYgvutV5uFBjfzhy0baOQrei0zPqhf2qnfdPF4748sQFJjXjW
2ZSSQhz+11SnHzE56nrEw8EuZphEhxKLwLP/WEhXDvt/5e2vVmpUgi8N45GMj3ZD
cshOemrd9idQN86w9o1t8xYZNBbsz5MnPArlNvji/X2BfqCCAcoaY+FwX22uiUvH
QUeESwvNdFLB2MWgE+WyojuoGyjBrI7/AQqNH24h6RQVBzJ3BM8VDzp2MKu6PJIZ
F4IbPhC118W83v/2McWzplNB+aQ310PITBFMAV5C8hywuRMmxRsF+C1oc4ufV6Vr
o8iMUdwhXxP66ybgH8E4ORYmoiU7/9n4K6g5V9gC8Q5VMMZd4qOAKWHfTGLf11Do
/s1s4Y0RHMUjPMWyDJLY1/0ZEu2lCk9QGr99IlqlKLRl0UdV2yyDemzy+zMU1Cf0
4YSbl8zSEd9ZUPnuYjvXHgAtXe8mTqYtaL68ARbb8NW+qya6dqcxc0guWbzlfPbs
pmCQkHRpUkEGPYUK8rGKXSVGk/UcGtOvkUGlYqu+jdUOpeskWigSPIIvCvj3kuvu
tgodNIK+ytkUVGW6I6xN/KbWLLDdYD4qh/Xh2jqHo26sFUiDOdEyLGKomVL67xXP
tZwo6Q++r+Ymk/9snMttwpqzXiKUfE91jEeJToY0jpiicR8q/rGqicGUGWZLkKu0
i61QytxVMVgJb6qVBf/bpyLl9YqXXWH93KhqYyqAj+ku25ZCqtLNG4lPN3HwYWWl
HVwivQU5zaQN3SqLvtY97/M93MOnBDombsJ19HPcQpr0ik56ZwkwBTFmoDTC+sO0
6O2F07j9CukYpXuAAKsQPrWRSau521cbKYSgcd/UJc8bMvIF34aCHT92SyF24BmF
zqlj92WFyJQ0tbtO72ITZMNdf9tD0or/uUgSRWWO8qX2qOHq10YElmtqxfQ+oVI3
3ogwytjc+VYM3HgmP67UXM88y5ehL/1zcv7zIGwZZJU6GKbpGy6eFiZfeda/VtjR
viV2mZ3++lrwc8KqGJ81rwNCmOwJeamrWAxHQ3RwuHHWAi8Oe6pSyeEsV7LS1gNg
Boigv3onC2X8WjBs34Zym/ihPGSX0L8+fbhD0PTuTwPhwW10FqddmSWN/Idxs+4s
UGQFdZFc+qq97Ih4xxmkRArsZ6Qkle8yirZtYWG7J8VGXjO91oPp/l7W24/vO4nC
0rhqeg+rAVAE/E+Ogz2SWTyHkJkYDG2YyCv74e8VCzPpdDFLorS8Ikx5xNPY+1/w
SDDJWyjxDqludBW+HVbGcI+mwr8RDxosvDGJQUGdxyV8zKzBzvvgA5Xxl9GKX35z
S/Wsb8s6E0vrlHcE8e7oar2dLuyeOY1ibaRt4u+oPrTAsKxnrstZ0rr6zG7uZA/7
i5ij+nb+7Geq5Xmjnd62Zz7qVPkrk4y1wxkB9YBuyEYOtFoEpS7B+6Oi2+Xq7WlT
rjfUzLmXnwhcLqhIvRnUikso6+tjGd0k3RCC1vkjcEeCCTSCq3t1k6rvYqM6JIcM
s0f9lPRPH4OfD+BbNpYGeWxFg2+AOPEAX4Z7FH/Q5kc7eGTLlyQZptmC6pQRR4wl
EK/YaxRsqijV48HRYVThKpWyBn8zCzece4gNPv32cTtRWMLTOUTrleKykVicaL7F
xNEqV7R74IDV/65nbrOrQ9p+l3Ty9fs3X4WT2tLAe1OQalp/4fM3P5FrSxN01JZx
74vvABBnl8kjQzxkLNvbFfC9SiSecqny93kENcvnPIVtVmUGYjW/4iLXU/ADKNy4
6Cte6U4654HAe9niec4klDcUBUFEtS19mv3bAPfsP/YISOwOpigZt+REumTcdmga
OBxUecYzgojyzvISFPOsmJXg3kfOqQIp42faLPcZUpbXFkwCSrfkXDtF0aWcXfOo
0h1TAGW4uTh8SJQ6nQ/vv/kgKBPobzHdPikpsMlx5P2DezE1G4BBepfmy/8NUfpY
3Svr2YtmLOyZzAlBEzQekYL4YAdH+PHQdSjNfGkH5JQtcj2MHDqQAUuo57+9utNi
SMwldbf9oWRVcIygDQUpqEvb4pC9LbEVsx50TSe2oXWtVXkvnto3MXVmAO6hNmKz
PlZzh5+d0Rxnnb7THJoO2EK58iP5RTwFWr6tfQrWAdvONRGRWTJ6R2N/l16+pSSu
twIdJPVEnaRnPgoO22vW4P9tTxmvbUmV7Dr68tLur45BUGjj0pnVs5R33GPevZE4
qupVB1/tIa35YBqykMlInwAK3S7urhs1wMbR/Yb4QdW4SdnM5CPkd2sb5HFvFDFZ
L4MFb94o/7UphKAsDS/uwQcas1N6CSg252/KPPqLjS+f8TF/mo+btTmqYvBODrzN
ZnSA23dC8/tA5PSaRAiiV+xFXEDZJQQUxUER4m5+bzjx3+KhYuUpY7fJ2xM3aNeb
55O9LYgwlhxffVOnJ9S4CYOXLT5OcuAWFkgg16xf/Ou05NoeON8orTY4aVDtU0ZM
h7rgKCTKyfJFIXMQdfoTTG6lNXKZZojxjBhlGfzVWFYNWu8qRNnKgHVvSEVCZNPt
OpE3CHYtWEeEDP/e5AuChnAMgPy/5iZ3SmLqF9HWmLsn7aJPwUGE/vO+Y+/qJ+EE
gjYv2V5LEJ1+qbJ/DpPZnm3UQhbL8qZbaN9DTGlqVkHeWiWImlb9OTaQK+J1fIxm
2lUz4+VeW6YtK7oMFBGHNXc6pipmbTQn/kuopvOVEgsF+0hyMuMrjhUTrIGOdVvc
UH3dLcwDDXL/Y9ToWRSPc1kOkMTJcdQlnxhtH2A78gwJii6Mt9SJFFJeJtL93A5T
q1gQQtTy1bMPdzW0nVUTEK4mKCMU7AIwYv1j3kITNbaW2sl6fOr0g98KENhJoz7A
MtL4jys2g2Er6wQG9TYYrsNg3GHsZz3suYn2lVRQEaWvwJP9e1ORs62O7J7L0MU7
IN2g6Bgv/IjU6Qi/KyoWd7sTkTLboUz5ZnGqQyvlB5jE+DDyPxPR4er4l7RaME6q
VRphllPlCm7pvPmqFlFwNcoSUaXiPyQQtUR8q+OEHZ6MYoU26sQ/DP1xfZV4Sf4y
nqyRPn5KmQcRFVh3JIkWZWt08LqP+mvN7SWmnELWPmXfihxJPtowJT5bRKW/OjQ8
Xm4Qz4zUnlY/XnTVB2jmiMUqpWOiG6Jo9WQHipyrfqeJ4ynIgslgv4Wi+Nzwcuxp
t24Y8aW2FM+QAf82trCgaoDDKXtN262s1o4LgAURWUUWqyuMXmfblRrHJWvWsESb
Xw5Z54J1+vP9c8UeTWAZpRbXfeByh5zXH3IBi4wmV3OzYFdTlAqqSH1SiLdYyPQ8
OyMs/KMsyxawP2AdAWnPWdv0njCW3namwnflhUnYVOO03H1xiy9VAz9jJB/uGa9Q
SVyQV8r0UWlWDAWqitoGBXLVQZlk5KNkNJB1D6Jnfj1EbSy3yACZxCrN8zln9vKR
bROIvCDSG5X+A9BpCE0KfHyyPx4vTnsKDiEkJbg2E1sip/dgvRAwXks1FYypiaai
z1Mq2e8HjipU/8tDaUxzFPoGWitXHq3sgC0JmWSmNjhkMCOwYTkBgQQJ9Ph4Ct6A
UGZHBDGIPIkIBmhJDdyAx1UVtzVj5m6KGXUrTqge/8rXWSSxq0qQrP1wPp3tOp53
iNy4MFT7/rojrnjKZcdA96qQSCAa/ANrghgFT3IDyD8fHeIwV8Pnaz3rpMwpZ2XE
7fgp6WWaxobaZqtbVuD5FIqc13pwML0+hN5Qmx4T6m1caDwCocgmiaFsRWNisaG5
RKKdzf2ULmMhTdmqL32hO9x8TT2Gwu359UeqbF3VzdLBucng12xoy8vQrxiaZJ7b
YpUEFWaUEsbQNgVBwj6HjSo63ZAf7DkbX0tYp7ss0QGnkauaojqXg5Hp0YaaZ2wG
KgcgN2aNF0dw6xOwSZbW1MKsbkLORBfj8wKgtG3t54heKim6HI4l3dbMc/BYFmph
v4tjqKGWLfvTylvKpEsfPp9WbxRnNu3MLfqMa2bliN4VA2rm9TgwB4fdomYfCi96
sNh0NI/cbSe3sj68nN/QIZij9n8NfAX3k4Nnj6/K1LqgZkFK1HuxDZKAiFmy2V5v
yLXzpzWk6kv0s0PjtL435+G8dWt659we7VQPOVEA91n8i3nyENi9V0bQWwc6uCFm
IBYVDCFbJgjgQBcwE5oysGw8cKBqehWzQ4Al5bUVJl/6KN1vIu/W6YnrXvmzwF5S
0xVUgQgnGaoLlbSHXOIKj4UgzvGTX3SFC8TXlEsuDyEmMEPHSlGrf4AKRShq+Olh
zkdPfAn2GbFbGHVqwt9lfdTuMrWHHgEQVwO8bM++BuzIUpZPJZVgR0li3gxWtAjb
V9JGcZLeGmpgW73CD6Dh3YlYGjHjzL7kBI3ISy4ZdNyLKK0gfACID7UvrOhvoyew
yX1AQEtuTKZbQgHODD6axUq0Xsb33QuYWnwxFDMEAcklP5H15A659hUB2FgPhEYy
uJGAh8p7wWOfypYruT0ZZ0aTZvBPXaXwzF3xKKs23SgaV+v2gxp1AAGIUTUMq/+b
NIeX0Vf33KkvuSQEpN/TA/kQKO57a+JknSrzcK+LJDAsKc7Zf+yDCtdvA8QsSpyz
02HrXbjkie8NpslNX8R1+QqYfgwDtnizfMrTNccBqCqtzIT6ydAPfCdjRAYBlv/J
sjpA0OBWpbwBZC/e6xN7om1fzZMGhlvdsi0WxS9vzYjfgpSKRmcoJ5Qx5wMAP01s
O2UA2xMvnbJCQDNLcvQl8kGGmrEb7eEqe6yqDvzEuUftFarSVdpkvQXv71+HQzLE
cLGjvlUuqIcmP9GHNYT19ugrQfgSeFh+afaWyIn2/oJ/X2R400/gK1m4tTiQPXOp
WDBHGL05qSRnWIsqtgBFkh9viHQEvzUfx+pSLjXd74nwvreIh+f45H6vk0nfcC1z
Wz1NMKhKz3gRMhAfE3CoGl3ZbJEGmLAFnYEgPA1okiEZXCJP0v0Pvr/M8jfqqSr/
ge76t0W9Eb7ZYBZHtxV0Xle2LEAGbBy763gGmXn9J6jRIv79H6x2ybrkZqIxQcQq
dsvWCritPTzu1x7jGAphoVVvPaUHZfb9t6eJZp/zA6LQTZRCVmdbAf3yiMcdUDWL
dFSqJMXqb+QVV7GKLpdPQBQzdYulhcI4lKeF9nL3CDshOB0Z4wE7+Lmb11DBlrT0
b+klUu19nc/4HaT7ob4pCwJqahkqmoORI5ujq1T8nK+y82Yx0C+QZvNKvsT8iT/V
09fn5SBAWrs2BBRR4wi93unoKiHVnhLWl+1LHiHD82IC0HkeHd96i43j+v1cPOPq
cgs5KimAm2AV/xSHDrM0g1DGhOyjatT4gySgL8YIOnE8eXqJSHmBVf1K0hefT7Qy
AaXVvJe4d+oFr7UyIvaAmiTKnFx5//C74ujq6K5gFYmME9rhcvf9aS/1W7qes3wF
JYW2iTOVWEHDwB+KLAdNPdK6m0LkvkCsr3UQwv6Kb5s3Cvtbii3z8cbfA6sTjgye
BlUdb0PRL9DqiwM43/T2MEbub8A9iHhmsZ4/DCk9tx+Xiv0EklIOgpWqyoj+Nqdd
Zgi1pSq3pJ44jqRP6QQxraKiwBw2xhAeWnaDlS/vx0RbTrXG3vYYPtnMYlzLof7Z
lwm7iDn8xqQ3ABKGOnYBD+aGSXJvswR731j0+ijNMv7srtA17j2jBdlQDUP+uHyG
ikFNG4fIp7vQQQ6oIOXzL4fKKjCGpYtgyfaYL0OFtZ+iOaSW9hjK1A7cWzK7LIZW
F6z8z4FtvNMqKwT9i0kBmAx+7RyohHSdc477auMdhyjoD8b/PDUFGIZ03xoB6pNx
V5taBRDMATyCiDbcWMwxd4wONb5Okqm+wfqZxlSL4iQBxOqka7Eh4gxgM6jjNmmp
hOtLbP5pqfEPZ8BUkfQA+/PlepWwVQmC9U/8+sSky6WAR30jdUITPqmRniJp+kPZ
iL7RiUxYzvCZ0/CNneST7lG9fetd0OyIz+M4OIajSOKDAittMMNjTWzFYfqSKU2S
1KrRw9O3q5JIH0QVUKB+/lTh+iHRSNG8gU25x9gGxIEO4UppqkIw93UyMr9enPeV
G30epjq2O7LoSKhOp+glzucjHG+XuzqrDEIJrdcEFwRket/2iNkYd5pdf+lLtBzR
X69jKXyr9gDohkAGs0j5ndrhqWQmDK6zJqIwxOBzkQvTFP50qitYZ+JSCra8U0Vj
ZK6vVlBnL3PzqlUSZd/+HLKLJFhTrJ/RaMTAfoSBTywNsCOYDRF9KxHdriX/kEw+
LkMg6E9Xt2LgHq8InYmaw224xPeKDpMfnZRvBcA564qDVUQvdjvPJFf2SGIGAb3S
AvaQjKuLWEKNEZxbvqUS2QMw0grXcBJmvwOJrWBxroKfnLTJXXTFM/cFwbCkBx1d
f7RlH/7IF36mce0UezvvOeoskIjmwiHeWuH4bIC7Z4o5K1d7Otn+xG2xixdfbMfM
LgOeSkeBhAHAHS0g5mq36pPH/tAk0ptDB/ohJFUXi/yguq32v3drE6EWmImdFoYE
Kqo8Ss2IBY1tvtjcfCmFuw/2mkDE4oiNvZ8ssVDMKqCBpvyex6Z5e66TnvwkBggP
P/2KUZ5JqcwNpjvDogi76EBaHpf5Anb6+RlV43qjjLb4rt3cck9tJkNowkjDGEE5
ILhLjJJ4tnh3NmzWTIUqIan7cE1ROeanfKl/7sYW4cqy21EcIbvsY2Tqs/9X+ig+
FJDSThdyt6Bnq0Xuco0+00yLU+3ED+mwpt7r5WDOtDifoBHQXP7R6YhI7gIsCwTu
nUoroVfhgKIm6UFFHY3ivBiK/v436f8ZiHRaIfo8t1imWavTpQAFCUiX3OqME6mu
3UwI2sAVNUQ9Qv6R8SsjAnEPyz9cb8+25ZwskPFDK6plsyM/m4oXr8EgtiaZ43gt
cS+2jM1eIF+03qecTygjVl5CLGV+DiPrKgryHhRpabCRheZ+XlH4H5zYUMG4qrix
20AuAS3kJX2uzSKnflkwpIWmuLereifAaQwFHicKO5TPp1frJnGWkbwipFdUf1a8
qqM4N7sIKc796sGZatplhZXZxilXXsCr0AChqbAVR98wged7nW2PEUqo5W/Ai+Il
o+uT8YUiCUcO6fwrj5otWJ9XHbm0jVnJH6cZ9azmVJcluQjsMGZRw3vpbDnljy2E
OWmZnHGaKhTg0cGBT3EWQ4JWhhrSjJ6Fd+Yvab1V1mSiYqaD1/fmspLgtZ8twgPD
oI94gJN2ARk09vdtt0CZsHxRSYsTGWGafCFgrp3uXPcwLpR3/GbJ9tPhivTHUcMm
AJynzUDJKIhreF6luDsbU0ec+FvBTsSm7ds+rxBSnX/ibM09QhpOA7epY+bJ59Ma
tlcg+UfUBpprWrS90bbeXMVBTtiy7Pft3xCSyG2xlbY51OIOThpDZ0lQqnKv3pKs
0WDLfwsiy7PRjix/sqISUNaqe79IKnDNMOLwZr668nAdQCifFX/AqRB488wt2Gb+
sd8tPnXRmdkLaMJEBaAs2l+6X18S8wvut+DnL8HCNQf9nLN3ggwIqmLSPGS4e7fP
FRFnRh65BVIEzymX9Y/WX061S5xyzO5T5aNbDwPFh2yyCI6I1ZrI4SgnRzaVonRP
4Q7ZVQZ5hDmhSAVsKkKqfgb8yNivuPfhT9vOZQAE+HO4WlV2+ex84TeoK1FuCpx3
cNsySmxj3WO4kaDVnQQdQBA5C6Ccc2tHlHkneLXLZ70xWHU5pvtXAdE2hGbnBOx/
GusV7Yuzz0E4UOBGZQHEDxL4QzsPvB2NNJAxNVeRfztsMChBhhIadl2Qdx8x71t5
lBvU9O8WQbOTn0JPmuym9h7PnP++aNYzikR0/novGr9pTCyqMWsPGbBTRkpiK3ar
Tx0/9OJ8+RimNL7czTTHO1EoLynIpVqtp4tRRTRxUtjcufbwdEOEH2OUzZ7/QkpI
7JJ3/fpFiz0WnZHP19Sl5TfH2mHn7tsvBqb5t8fJkRUhZqr6fDWTw6Y3htpdHUCg
BZKdXXY1UpzYqgN5N38B0JTB/MTO3c2rIbHyBSOnJhgvFDVscpiV2lo4oATUN9vI
KpOIM1xODYDWBoXNQ8ApRwRpVrYw0VxCTlPcdKau23uvgTG++VDfYJGEFCWDFcJu
uMGDWRwAEd2wqvEQGCKLYnAxh4EhtsoBsU93/hAGKhYP1Eznz7shiUeGJEDio+p6
1WgcpCGTozq0zhj+E7hXK9qT/V8+zlEwN6WtkCjLD4+RkybTJaXzDEpTdQUVxhC8
KfAZ2oGzEh2/V4us/Mu2biBC0uL4GaPDaPQSd1ZaJhVb3JN65sC7/dq9bEiKKVdj
vUuxFKr6WIiKjq1b5qSzoq/cpwLVhl4ANXbwCosZr2e2/Wm+cUNB86zShotOepih
URqa5Iy2ONf806oHqA3P4oOSH2kX+cvl41v0BnzrfN+1tpkjde7hjz2a18MalIBB
Q4fpo7OHSjZt6I/XjR8JGrGqRobYxBd+BtzNuS+ZcQiV+nIYxi/Xiv3sYaxh6ckK
Ghbz6NNsqZvkOl12FkpbkOF0UOUpjLSGxdQrrVhe7mAWaBYUzbYNdWgVvbCEU+6I
eLXUVu9pjT8wo8vOivjchz+4cS9J2iutzOxARynpbxG57rv+5rONqC/MeoT+uXsf
xOldCieuHh89fwbUR5IPT6XaEnoFIj6vYaKekhc/FDLE1Ejar1/S3BOUv/SCJI7U
4dmGWYWU4h9huXK6bhn9zZsG39nZugKzh9cK7BgG42jjzE0cwCHXP6Lcnh7X/Kld
6DyDVVV9rUIkgbdssUWRn7tuQATV/PJTlz6QhsVlv4Nf0OTCIXKwk5GcBaQnrjmX
c3EMFxZ6cTQlZ3HQaPITwuuEQlkPmFMAiLhsvChufMEJZSfdV77HRdwX4Ow7r7M7
Z8ZJB4tRKvXF+/hGgY46oRAa3R3i9ql8syCxurbM8A0oAtIJmfPP/gq9oMkb5V5S
WKMo69nEMNdCf9vbhh9yWxbs9yc/GhQAMYigVg7aaVJtab5UlOcL4HGSWyrOtFv0
/8q0qENG88S1kRkVDgI0Ui82Khlc1VsnLNqu+OnmtVnJFkxpYN+PDuG6ccoThn2p
buuNuTSVBC9lXVOGARXgCsxMxBFGSRLCcm4Z3TQRL4hbqO9Ezou90H1SDHaAerqN
2qZmjt3pm3OK1hzGQ226m7+coOXd4dgit76B2s9QCY19+IbGby0R8WeU8oE2kXv7
GEc4wyYS3KN7zyi9C0W2ItcQY5V3d1rSZeHA6VsEW5raTWbZZzvWLbF71iPHPvch
dPxL1onjOHVoirGPGm+2tzZi7NYGE20cJNYN6dbFCQ8/m3DdFtaN5k9tkurwsD10
sj6IArq87vDZkGE+W41PDUUWEYBO6bY1zv8mYrTOK3JcRig4dcnsd5QlWe8LT51O
GsiLgI7AqMa3aBO658vNhPyKYaCKPU2LSa++cMOR/9d9e3Ts8rF8kUOVQ2L11Wi2
iSQxoHxIGvrX5b8U2CobvwqadrIxYwQHjqy5kzAj6TmAFQ09HlrkuV/9rg41mGZ3
hzuBYHkWqefS2ZOm5AAMesWoJ6ot2UD2WUJ3l7ue0gE3Q3FRUaOdXuPMG912EU82
DcFv3Pa5ML9Po1gJamHcl2FFcIWOY/53OqlBBfWt6w9dYvRI0wQy62OTirEg9shI
wLI+mcaqjx0RfXVrT9SdixFUITjqsOLSBcY2R4DJj6r8qRbFNIm1qaQSmvtW1mi0
NpJAIYcWgQxCGEwSiITaz+w41ekMDN5LrCIe0vwUisj1zCcdCb1Enqq5ekwutnnH
h070KmtOIXWGhVl9FIvggknCVGnUoVnkWHsO/FkM/M18CC2nhGSC8Ar89qfidIPJ
4OHR4vj8G8jkLbV8cGRQAc3qcz24SGHopelhB5MaZAx0VW6Yfdbq7XCD7rqjqU3X
RzCkC0LHJJl/3+JZ9dADCwzccpCOXSHtcTa1jsfy2i7M5wU6tif2L7p/J+dH86sl
mIHOjuthuRmP9b5R+iPi3agZWClk9lEauNOASR4Yt6ScN3Xs+2EBURZfzLIGjLKB
MryrNDXsvfKkjGYBgTRnViNpPK9CyLabk810ftlYSj3+Vr8R+P9xCcbIO8p6C/mT
OUrDEy77NtlLZEiy5jtc6ZnP58PJLzArKEVrKWZZJfxs0hjDmTnI5/HQxo0Ij5gw
uiYpzZjsA7Byc9zvXVtGY1wnL8k9ewy//gpvoJOd6/kSThM77FeR1Db5oCSU6Xgf
95FRnPI6tGGqGldFKIiwSZOLUVqfdEpC1k8nCJRCIx+2wFDRODLxmJVa2ZbSnwn0
7I39UXKKl/VpX7RC+xZ5gXeHbizzfiBxMb1q7N7/gAw/PkWFDjIf1XsJfvojHuTP
2vk5pLJeM/+82fwSzju9+DReocIc2oQECL1luHbJ3alOpMEs7fJsxEESm/1Si6Hx
t2qBBwu3bsgeGTdRtqMTrE0kI9B1mzHgwkghKlFk8pYPnVbwwmS51qVfyjZS1QCz
oFXywJikWxblH4eBTFu3Vb1/U2qyPuNOM1SkPWpHVkp1ehXoqhiC0T/JfwAuhlzS
Yu9UifFZ1PjJwtbRVtVBnAG89w7usZZ2IxZqGX0xrJUiXWU+hebGY+9GMyUIikOB
Tlvl1tBR/L2izUZyCAUYhXdwcvUYkCWKV6qIhppXH96yUOZF6O/+TWzPncZXNBXD
DnxR5UoJZf3k2yPetzc6E8FzXJxPS7uJ8FBu3EaaWfcF+xlwIewKmv45ZRQbBXMC
vQeLHHDp+O1uzF9TSa9JPjqFAU3K1djwnjO8Elk1Gaz6y+Hi6Ij4eNOFidUqLrWn
tXQ+itgXzB0A7sQ7QJdkGaW+hdP2SWBd1CndYY3JIh3W8opicKNqvA/2yGwlqacU
4s+Ny5k3MIoGz9bKlah7A+fk1o2mFE4Goc2aBXpaQRUhPB1jyyfcnsOpsyQrc4/X
fDMkDZrzhu3dVfGgpzL9wx9Xi985QlteR+uq5EHC5oP/qkkegHXUZo1/pOSVYT5l
KnjbxCcnuAHENPEDtbDFccMBphX24BUWWG4EyQ1y9s8NfUkLPD/pwsaPs3OJzFbQ
injeNh+GdkaZw5cZPWA42f2YoNf6xYvdLMuSF3Lry1hheXySmspvnH/n2bCA5J1n
NtYA3cIWJt31DcZIjQvrfm6eYlobMgHyo94ijFIabHSj949LJXJYImkAv5dlOQJR
iGC8GlDUdmk+lfgQ1X7d91U38h58J2DBQB0kXBwm4O0lGaWA4qF+p80J7F4QkEWe
qFpHEvNJRl7XWL46JCqdY1eLQrxbtorLbgxMKW601CiLJ1smFVrKAXb25ExS1LbV
SpoL5fTsGX0OEyILHmuhwexT5zrat0vX4sKnf81LJavYLW1g3+nCRtNJYb5Xtduc
Xc+UO7kty7vje5dF+x/g10jFcjb9jkaPLMF6i7pKZUFzCblr8CoLCsz2DnQEz79e
jFeNgfS1yIc+ekcioqnuAHo3JjGnpKKm5qGJrHBOh41kSWQGdmMQZv6KM7y3bSF6
kosnXDJ3Ir4AXYew8tEt43q9yjcbZDLSgZ8kXeuOdQkVyuQNorvFJacLE+9arwbB
N1scZVI60kYlHCI2E3EOk8dSiC1C6Qbz1N/mVshgn/7VJKd8mexE3RGTpd0mZ2Rb
v/caZ/xCTxNSf/NMIWhj0HL0KewVWT5S5YuYow3xXkjkdgKTfbHcvzi+e7db3p2U
JD7yhqwR2OlAFtNpt8/5Q3FE6n8B9mBPwrnQDmpsxoc70MpmEnFda6Hk8gkwVAJ3
gEQPDMnSSg4ZeQPOPnPFGKGXg3B+CVvCScDDpy8LukAdg9EBW7BNB+pkvZH0w2rs
NdhScSufYGOYEWq3NTayaK4ZQQO1nwS6xtg6pmSjDd1DfwlvlHKNN7tBjgmLe3IT
qmmxbT8iTH+T0Jv4PYzTvNaKoFjTDDa/xhktu42b4xjosOJJ9KlJjYyYM6OFuKfm
BeKZIF9Qvqx7nr1ERnEcu5Ue2svuvcduWprlU94FSVYhBKcLSYQb3ep+FiU+rWfv
93BHxWAfRYTXGA+P6b5ZiIjjJJoLjrjc5+jhIk+10ZaG7pluAI1cYZj5scC0ywj0
iqfA5DdP3lvUZ5H53ZqFoWJzIvg3Dsv3KPxQErQKNhvgdfDGuTQIOGYyX9GaZ+kx
A9h4JnCUjibKZ+ggKsMK6xOoRfcVWCnad2z0ZUwMkcKEztwKZgD7Q4a0t3vlcJO/
exovM07RwhL1R7gThPEOR2wYzzGRwJ4His8yv6WWY/aHr86klgMNoYI2LTiWc5hX
mgHS/U5eYwnRhCfSQOZPP5VDksgK9sjQJhL+WOCauXt3kk9OVlOMkmOLtWV1h2yA
CcKVFedykRmlrfI9/ipf0laKIQyRG8gZqpUJpMSsRzvV+HlBbtRfHCpFAoxTH3Ka
BBhYblnsJziUC4ejL5vlg9HErBUyaaIesc6mqd1pw3uNVI/kPxO8E6/mmbwnGwrd
8FkrggTPNjsTMatfswww8hQma5tMB67I5P/ExEFhBidiSrJKkLN6nCvOaDR6dSca
6avP05rDdgU1nkiFyrRNN6jGBO1ZmxD118cdxpuJmSlvSDaZSU/d1WTevXDi4kDO
oam/6ucEPka84L7tTXIo4AGnc8x1H/yFfQubUJ2m9gKO9bmRmKXg10hYKcPY0LtR
AdX5b5ReyplrFPwv9+R1s0qk9KMZpz3uIAbrTVJ3oGbOiwJPs4HT5hIKLySBrJzk
O61GflDc07vGZcMXTalI16MQvIw/GxESTsC/Vxz1NkBo7YMesvq1hPswn598norN
d0T7iWUIxfe0mZ6YuylQkAxwr1i5tKX7fph7h3VByOUanz3Kr7Jr1gIxgs2Ql1cq
zw95IjSZtAZvqcBoodHI7n8iFzn8wdr7mEKY7ahdaouGDdY3wYzcswFgn42+guEN
zQ5/MPqTgmILTdGx1Mk9+tuS+Ngs176Dwx74PKJmKd6MNhMDYO9iDpXCTwJL/A+c
igv/5JPDjt0h8PHBDie+8rnrQBpBjWXH3++1Ko4bbDNyIn64dhiHQJFL3JDOZx6A
dP8tGz6NIpSccj96M2znHXu7UPNSi6J3Ekxy2DdCIgy1fZ9JJZNKt4UlGuT72myl
8Sm2PkZC0kPufizPAfoDmEbqaFHIfpg0P8ltZhPv7XxtS3kH8M66xXyY0q78sca+
S3lxuS+Hca38s3UdGBkh0nhd0NGal6rfvlIUUlJkEF6Al6tR9u2zPQ9IL3c9Gj4G
rMCfwvlTUN8NHtJ6swFBnuUF9Z9Umf2pjtqHMhkumAN0eSioh+tkWnfhqF3y8QOu
WlpZC6/2bC98ukunnAcwq99p4dQ83mIN9NlHmo/VM9M+aywSVQ0kyN4sep8kf/+R
c/+tqDIqg0ib4VDo+ck4Bbizw2AFKEp1+S/N/XCK4rks66pdOkuQot/ffHaOSxfN
pOR9YTR8IBhJ1O/owayKwFIasOvxGrraAq3XPtBBi9jlFzY3mxiTOCTF3T/clWpl
N3kS9ekoJtZWn3t8vRpaQ4ylYAxmPh0YoKzOahJ8UpFcBq8LKGAqq3GJOvjYhbdO
H5NfNidLIuWdW7VssOlrFtxeNfhStr9cEA98ycCF6X/c8zh+4y+UaSUzzGfcHRfc
dfPPUbFbnX9cGmveB+vruqqccH0SnyvFr3J7ExpvtGY70WHwn/ApXAqkQGWVfFr8
d5HUHH0WdXkH3901TkzQ4DYAUCfin4E9sbjc+ZCglc9yF27Q2xGtnvmASZTbbtsq
pfEUU7l9UNVA0uGMBDoBJEr4erZVIGS9PDKBByEuThx+Kk9QvdOpQl9Uwh97BrP9
52zoOeSSqkdF8ZpjWLkE9qshhnmoZSZK7P4KDUAHJygUpsYHEVA/dRBXls/MdbSp
jK8m2iixB+mfvM8eooq2hMbWB41i9Wrv4KNaWRX1jrmKUIc1aSe56erEZ5NIEJk6
M37zRX8Qke/fLU4xjTozf+OJQMWKvPAXD80TwUAfBlrt2Qc74+Oz6aIcoyoF2htK
y/GfseAwBJ2DOJVa1XvImHq9oaJtM4kcbyY8oGBy+Oko+kpLiVGvqgaqCrM3BnqY
eV+wNyn/9OV8aAl31R+K9ZxZCcSVizGeR5bE4+wmRyxbl3pAt1jrcfBjseRdSQY6
mV5+N997t4ZBddZYuoas+wq/rDtJF4OW9vhgqcBrHeeFPQ57U9caXPARlPbLfh6J
d90ZAnVqke5ufRe2nYiawuU6kfqG4x0I0GwgIE4fCG1ypsILy44ZTmWIEXHNECO7
2mz0U9TQFFz3/fKZrDinFG390hK5fnysMTMbKpqnRWxUKbchGiANEQYuzyeVQAQ2
xqm2vgznDPNyu5OV9L6eo7LqCZRFGmgF57iGU3sy/9t44h5P1myq9n35YedDjaiW
X2lw7JT6BYan0w+hgo+7rA1MNvliQwu3Dtml88sDR44H6j9D8JYSFTDk9h6hrbF8
affl0m1n1xNEBxWAk/nz3eWfR9SeoJMQLdsphEb3TaXkv7jTbZ/6o8XJyEf9CxIH
2JTElqf9Yzr5PmOObupUiE98zBCW94aCHGJva0zGPuK75ZqcAvkgYMBKXbPw3YqM
UlPKvPl5NamMo/NFVuTogiNoy9tO7B2yG04MjOE9Cz1gP0awslQgIMFewNEU19Ah
1OyYXuyH/mL5eCohNMBwlvhZzpnNvRv/GCTW31ZYUwa0HZgi7nm9dWEUrPuywZRS
A3GDeJ0WEDI6xTWMrXDhxFoKmuwfswGw0MNy8AKh5A+UTzMZLkb6PPQcSJWuzlFo
TYi9VhQxP8fltQ0jMjPkn02xb+8+64q2kPE37Y7CImzlbySvygEwOWfRKWZVhQtQ
VAeq8elBAPjhlHsfrEqfDtUarCT5BDR2cFdS2sQHYA8rxJFGL9X15z1Dde6TGip0
pfioDMglTfCneimrfqWIo25eSUaGCRUI88bCxABdcReVgr6oot1zi2KGRdxMv2Ts
4CSqiZ+BONdsBxekL0zHyPjOKgVUnQSmPvFxtSrjFf6qRpZPpQWT22hGe1ayIG6T
QlVlDP5NtaBKW4s2NmijGWF82ofMEp2KMUyLbtAmb+cfq9po3bK6Ipiu+NhTyAJV
sI5/KoXokrk/uGsRw7GPrsXHbs86Ui0ug5/QBQzespvRzPHuK0VXgm3+VTx6/Hh9
FMU5R1EqtUt25zcl+ciOf1h+cp+WxLv9bZIITJK5XNjcXkA+in4Y6qp5kssL0yvE
nqJzZ2n2FapZYqJjCvpd7Gh3boVPUL8h6GeajgpdDo7K/GKNKv+wI0slkmrPjoVh
ZswRPO3xwybZYjd0Z+6r7WT56esPNEL3WbyZ3LRMQi9i9Pz/NytPQyaI3CAYzWFz
MVB8uvfgSLeoc2Nn37ewgO8tPkRp985UsyZq0eJYYXQ4xlhBK25ay7vz1YFUJC0L
W8DDgvVQIYaj43rExTEcd6kW+KowM0e2jEu8fPRsgjReRGGD1lf7V5FyfBfBxPMa
vFEhM40c57EUPpfXM0d+IFqm+7uefQRcY3oBohHkwq0NI5yGHsOq4sR5c58t4LJt
KgvZK9SXf5rgkoUgTKtoo1ZM51Y+X3BAjbCWcuT0ilDVjQ/o+tbNEXvwI3yHkuJj
ZImjHrMZjkXpTPx4uGlqeA43Fb+10Zd1xIfolCVzaIT6mPidGVfJyGE/dcGYCEiG
kL0ZSQhXlh9+PNzjA59U35KSk8U5u985yVnr7ImlMTh1yeVOtExxkfi+g1x7jzwI
nGKO+ccZsdz0PY5dzR3DJr6ESE9oAWyV/PqdUrJKmEiuVFlnH9DUAk32DPUQP42q
t0qVukFYrZ8XBOEB08DXrddq6V30ItW0HLyk/dfrTyg0yXrb3iRarv2yUYgJc69X
lMiIsQqlvf134BAzadcWMtM6wB5i/dF3mDcvWA61Lvz1TFweTDim+g3dwNXp3HCj
sxqG8w7HxSzzxDLh9Bwx1mBpkijZvyPl3NDvCCgS6ZGBoxvDUdjMsANeRhb6Fcwr
pTBtJdSIMd3XGQv7m5lwRyMNfldp12GyGVB1PhGkNOzsojNQuC9t69iH0SRYfHQJ
wCRSpjsGbThvpSfI9M0nJb1XedLobd45m+NndHmSH5QQdV8ospMjiZSvlRQNAmMv
Rbi+xrTBmhoAEr4qpKPu3hsqIlUKmXV5/pR2Wiyd8Uyy5S9zzWXshKM8xLH0TjY8
UYQpQYuDcq+1A6iByq+rf2pEhPFToY3gzxMGnUWVp4j2AqG1qMoXqXueYJsPiWom
EwsGyubnrFkZQuQGq47SJtIp2IG/H0p37173WOH8L9vDcYN5Hue+qvKHlj6vGwaJ
fDVxredT1ibEnFRfbsyl2AkH7IuPmFgsl9Lhwg6aKASV/TUylSByOtLtdFy/Fwdz
dJF4e16gWMNQpysb7VnZHJPXDTm6Yxu8XqubYPvDJul97xBjfUvjPYuLSu1C1vEt
oYLHzQVOTv8fdFYU5vR/DU5AkUehIBOAiuWZe8c+4LP9sxKntPIlimxLfw+ANG1Z
JvSr9fkJ81ZsL3ALmnObNRJKqg9ABvZw5x40nZ4sX9MD6cd6qEaesDmbYRD7EolK
oUITIexo68Pcsyzk6KE3FEXZOivW6HLdqU5hkDkMyFG20KA6tfQoVEPAMn7ohYVt
EGiF4XdFn8cGs5BU4Q3cBnXMK5ns5cRnYZpNiEkYSy4f7J2b+W0ViFVleAm1FXSp
6WD8UaTu4ygjgngj4chTw1V/ZujFZWH12vM2ICEk4bibQmWz+bsTMx46xI84lqlH
w4PslCgL+jR2CVoT+iO7UuvYF8dI0YwHB+eP8eoKScn1+E76pIojsMRh6uNtcK4l
Hc9tbabMu+ALXkgkPK12d5BLP3CAzozOND0H5aeAjKONzHiUHL2BgTGImyZECs26
+bXl5agg6/nVYL3zc2ca9t+Y4j6lUQ0qZFh7IBF1jdRdcmkD6Qwk1AhIHRoiwhXQ
gP/LLZobVglxitHjVOwjFwZTKulRVIjmquzS5TMwhz5iytCCcxL9TzY1JySmP4l1
ibG++7XXcB8fx4g+G7niUTbktpJ82DqorLhAXMcs/arhNyoNaTTe19F8A3bkcUfj
e2+ggcboXoktgsaZJZlXvf4HNzbSZgGwvggVdodxjPBB0FLYi26Yj6IerfABipTW
la/beM1fWh3jsaxxO6oQmOu7+ddXgxPA0zn8OVhK9b/mg7s2YfqMaAvKzXLIpUZB
jaTqjDSD4Nzelcz+wT/FlqhIHTYufFH1XqT1WSb7CtH0FvLruS5Tez199v4j9UK8
+MXfVD3tlVebJQZNjIpt6PeOhEfd5LNhz/nYO5HUgmQ69dKDuLYbK2JQ2yCOvjY3
d5OlojzXgF+AwMbzFbB0cA338A5VPg2O45hmW6ft3oFC3FYui6K96ZtCNsn+1Ejt
ZTLWy4f1qPbeivZmndSgNV3YuyCDewkG/Hl5bLIwqJIZMEpsSJDCBx1wXmKlyqq5
1erFl5dPltVjQkwbjj51yY3DZn5aSADYsPQcJOK1epxt0hTBsMU64y6xpqAAUWCr
2vhEinc9xEbnOyTu9Ku624bbAT48mH3i1O5Ek+HBTAPG2K71Je4LCrXGNwRxXTIE
CNHh9NCroIKH5XLb5S3OM2GBXU63omQUFAEiUhG82FQA5qdSwxJnds8h0eEttz/C
JMYn9b2vfRYe0+pvGjABaUmYaNlfKR4ShDk1EjPTYHKYjWplBBttVGcbiMzZfgKT
8HJF0r3YB6nqVf3TR94okj9hKZFofcOLDl2tOwksuusORGZrNk06J5wYWKqg2BDS
syZTOuBhXDvu8fsnlfhml4M+pRiY1N49cJxSstRsJPqQaa8GN8v0NZIxzDgWphYX
ET9juEfSmDFT3LWKjH2l6qKkI4ho24AE2P1cXAz7h39pxJu2ZqclX4zzaFyR1nmn
KfZCkfpNkjTowRtYblKI7uDb0ARr3D/FRbpQVso+iB7P96fJO8BOdkVNjKx9m2UM
G90EMx4Zp98zYcEze2UZcwAc+CaclUp/FsVAINd4SIYL+7mhitp1gx//8+96KHQM
C3ICwuQchcwF4K1wgFEtPYUUhhbh7fr1efiF5lhI9PO9L32kF1+5qL6uRIhZdHlC
xlGGkb9VPMgpKeMr7KNlHeYzL6lH/FzYW3AuDAtD+OpF59lm88j6OeX83CvMNIbU
AW99WcRajFi5NEOa052rYOnLmii1/17UV5QFBhwTk9/M8lW1fMjFG7wIWmP8Ako8
89QSSuHAO06jdwylX+6qWSfgH6c1QqxtLbNjmX20UH7pCg/WfGxNY3JmMYhzQPaE
MSf2SOIFJ3kQzdClqmx8/CYGmWs7+Q7lx4YD8HidoFO5dHy09Rijx8+NBKY9f6VV
S+HS8j4nUJWTyCov0vKPmGCY16HCFTulPmrTgoJs09IoO1HJS0vHMJCJ+cBScNRc
2SuomFRS/uHZJdw2ZABp35ux1b0VfVM6qJ8wuEy5rxKxy5FwvgOV+kU9Ulyi+DOc
fLeQGiCSnwT0nBl/aQRYHWB3j+LCcA6/eAb/DFe5M5RN3xvgFgC7DkshputgQjrs
f3XpIiR8Jw5a/KDykHXUQdpYoEH7lup/wYBoZftXM6ajeVcPYaN8Flaz2YH5CW9k
A8SkPDRmHsFDqgJ8pqnexHZiKXGmJ0pEcpH2ajyrnnBmoM+QXnOqtb6TFafsFUfY
qRqh5G/pawK7SO3dWwaAdinN/sx5m1kUngPrH34sKt47SYES+ECwLOEM7Fth9f58
je3gmwRWV4DyGW1l5MbxH3MU686FLh1NEmHDDwxoCvP86Sb6ZXbQ2exEyFz7Ei46
3hB1hBXBhH5PeCelChxNie3eKgPz6Yco5hR+FdUudBWKky5QpzF8MMueC4yOUnCq
9X1E8AP1g20kVZArCo8n78dvwsDAMj86t6NMfcy8bIlfboLP6FAjMETto2bJ7+eg
TXkLjYkqdJMuPGFNxy7oK4/TLjftvjtdU+03jgffMOsg4oaC792guQ/av8JN7Bgn
eNFILW3ZJao4yEqX5VM01vZI74YKen0QBvnQPWCa0h1nt9/0gHNuRA7fUSs8e5LZ
+uI9BbCXIHebXE8C20aMlqi7j8MyS+LcksVcBGPIk2l8XvFtznEEz2srS2LPUp1/
kIZyuIhJ9qU3EFhIFomGVSnrjCToS73FsdP7AKhHNv8A1xqwUVE38snsyx7iB7X0
hENpTWP5ept9pJReUxd4pgKkLpkaBTl8+h2zuyWXx14KS9ktmbOdWpwuIr835JPq
l58ywQtf6CL/q+rpJKyznR3GUfgUVSLMvS2esH6S/ihjUCks+lALP/vHpRD17kH4
FMMvBzUQv80pydGQawljR/nMrL3qMMGalj7JPoPaZvcZWDrKrxfba8CR/CO3W7Oh
Wg0LtWkXCAXnt7TO6cf1feFRYuUMxlMvlCwVD9zcDCSkw9qoRCAP4rsCOvTwsx6Q
DUC7i81JBUrK34Dg+q0ddixMgtTv+Wx+TwZeY5bVPWqbVgYLDSB68o0RAVmrRN9j
42/tt+CFMbxtbTSwD8Ui0XwypjweOtNnLxV0LRuf/BxpiTR9cFKuHyhLD6pOVi4q
1acHBl1hGjuRg+V/7cJegXGrpquOgtpcLPDF+8i66IBU+4V+W20B3N6qqVXZsLAl
NCZeaFqCs43n0Qi9py3cZ0TBoqBLPq9bwuDhPLEwICWN1xWaU6dBXF1W2VRsuUwe
t/PjeERSbkDsgLC5kEq5uZH51KUG/BAVabcgHHPrPfpNR9lId5lcyXdOkwJn9myG
LDrPcpEjFPQ9n80UI+V/srZFuPe6PHdTCc8S7+098Il35b/mpHrj0SEcRsbjA1LI
PmOQV98O13msGwZ9em16pb8reXZnpMUykhkDUGFeWAJSVy5VmJSRFSLypwNNcsNS
KvMsV5oW8JBR3XaAh9DXr5mH32h7DqUSEcD34rCcnVN0f++jLXldH5Q3KBm9/0aX
Z9SQ8InIWYibyXpDTobvEKLrLHrlVjlXvsC43Aa2nro7DRX+eztvizMFurpTxWwX
UGdFDf4ozWZNCrTjPhtrXTnGgGrv2LAvwJ+eAxhh+NUif1uoN149kf2WC/uNMNQC
NUrX2OjM4q4hTYlBQCOZjRGVQqRtsr/fCmSpBvxTgxkU71i/6ntDXhVVNNAzk9cA
y9dkwnOMHvQ0eEQQBaQi2h7xkEYRM3Oh0OhngTKkcu6S3RAZxMqxxjuRXKlsJwSG
gLVZEO0OGNBdPuytFAUWnAsagx1K7dzVI1kLY4SednaNm6m9pchjHycboOww17dc
84ZDX5W7sOUj+0Y+2GmgHKphnGSxRHENTA9dwxllZ+ILTxU8cv1J4b4s3Z24NngZ
pS7NUxxfDsr6tYabZpep7AwXZ9FmN8JVKo8QBifOR/6akF5uMii2oG1Ktruqfnx6
fxABO8hBJepGtJ486SaXMaCiAfZl7Ox9Ugp7//LBPHqRlVRv3GVlGEu2p8+fQBhY
E/0cAdJfRvVOsrgIdAhx34sHCf4UFAoHUN2msFXJXhJu7OyvXni7pXh06EIhhdXT
DVDfzjjP8VzU70EEcEHSCPAV3fIw4BA8m1EvmoPxjCdVkgEz4qfBX31p+zXSXwdG
4BwCFB6JkY1asA7yytw5n3fq68NqFhTuOeQ/Kd+f5kmJtpR8vpL4kyWocgUDgsc9
9MZv8zSRGUrhw41wLOeMHk1eh3kfKIWE+zEgnI+crqfg2og1n0SRiyd12ttIVM46
bk4TAkocELSV1SjmdMgYW+h+1uHdcob0Ms4OIuxsbcEPiJmTpS1yc9ElZh5tq6wI
8y0HQvuycpLcqzWfDMuMlRlP0UnhegCbLl4ZKpxymgxaDB8QeZzuptrfT9aBK3BL
8wiRphKnJGD+uGkKuaaycDvZB8eFoM0RwbX6RooNuL3QaF0gjiUzY4OqehZ/YO1X
hs/EI/E2TYLbQz8H8bgDKIrQr90dRf3UkrOmZ6+a4FUIFVaB24PtzYSS9DtmuWPw
sKAY+PwiW3IeJwRCv6h7s5+e1Rk7Df+k3IclJ1sZJXDJvvO3S74wxHCM9T3n/Uw2
VdLLDNDKnKVBw5kKTasICchH1cAQQD1vyO81l0bBEV29zkN0zMLFLhF+MzfAP9Dj
5kraeBKh8yXzhrQbCWHIBYeKZMBVgsZVTSPHmBiUaNQhlqGLXXCwRvq98EDOupb9
r7Ecf+xOd6f+dJxnCjN6FO0gHInHAQlQZ/duklVvTgwoeD3K4Q1NK2dN9TxqsGNa
xDRPjqEh6+VRdqueMv7eKZw7suP3JbZoYxgfOWWUgsjw3s4rkffOwt86eaqqGdz9
QyB06iIHV/9kBPuLK6A6oJBDyB90GpScWsoDySp9tcpKA/bfkr6nv+1KbO3XCkcI
zxaHaXXW20VKy12AjK48W8HxsG3G80g2rDGU3Op5fH1wEsg2VQff02tXemrXRip/
4SgsPDdwGWjfMXplwrRGpPyOaS+ggoN/Og9X9PxsWQwi9BLWNOyGiJ3+3IL9xre3
47LupfJpEV8J/h56b92tYs9cb8J0voFw6j396ZwcYwPuXDDBMnQjpW3FD1jSdvaE
ppACFQ5GgAM6YQZauMBNROMr8qnEZXikGUMp7X0xyqhpkSJ6rFMn6ujFFY71OCJI
ptKRCn6BNTDzOOsmjtImrVlh/pmitVDHmXT6QNXC7iGdhxv8D3I5DItxFn4hcvtw
3sf+swz8Y2ArGYu7WH23OBHBTX+fw3PvoI+O8zJ4GSyzEmu0lSG4WgLAGYEixVRT
lo+AYhJN5CI3voghI+o3g3PhS2VbqHme4g5i97Sg/fSNB6PwH2MIwmPwghcFdxkq
HKRpFmOUojPJvEY1ENHyw11/5hUc5oToa23WvQ023DOplFMs+zElM25GpPgoF2mY
p+RH/sVDiEWMIUEV17GQefoHVKiKhAu9t3D0II00aD1GcB5mhMk6ZmGu1iPdFfGb
JNdbRzO6Aq+Erj2zFfLib8XIsaLKqPAZZ70Pbvap6zPCWdaoiEc4CKhCSl0VJM/9
8iIS6thRYILHvnULK/T+U3fHB4TrWmeeZ+fZur/jnz3NoV2+aKpymPqczqjh1GA9
DRgLyqaAbQCNEPkG3OGTOMP+AFt0Ldb+avpDAygyfiv/wwtnAE0w0bwpi4bJ1egM
SXbAvJedV/7lQreBRCIjcxMnVqeeYEAcpbP4LxkH0eUZugI7jYSDqEeZfGXdySOx
wpqexWkJGLoK+qKHUt7/0fjN5ZEF+bC+fpV4d4Qd6PtqrwoqCnbvqdNUbgDJObng
6T2q4JDxL+ByOBRlu8B2cVFvPKig0C4dm6B483Paw38+SO2QXuB5ep6aezWE8bPG
BCNUezkczniMcJrqsvVilk35OECN2k6dTadjwf1MrugZsQULfj4Z31xByAlxIsEq
PIZ/b7r1TLfuqkacRjAPUHNeBUQavCw1E/7wHHTB1q0Ml6GVJLpqE+qRUeKMMw7c
LlRMXxylHSBjC50ausD6Lae0JggPzxk0Z3v8VHNAc9e7fbSl/dP1MbQ+vn/Kw169
nUm1VFXbtXyC+wClhZcb6s21fdLmvw3MrMWqflAKGuvrT4DBpg1B2wrGcS6C+Qee
w2jJ8Uc9blcyBX5djb7ydXQhK/OCiy1KRMzCgXJnIEm4Gyg0J1HEPuHbDa8sxQJM
ol/c5D7455nqnMsN6YYHmiHqbPTGcGio+YIuPhLK7/a7/PTV7Crji9m6Kk5omyyl
fQJTd1+X98S/1gaj9OzupamXq21lJLDkOnur4c23o8PACTgECIQe5szNWdlAdIrq
3YIuHzO2kPT5QhkBHkPV3+tmrrQ3np/lKMeC4HJ8YQOsraglPeDEH7IgOPl7G6g6
QmtoEXbJNu6JdMuf62UkmrdbHYgtefaqDJ42eJjoM1MaUDKpliwygjTye43QT0sx
/T2uhx1m5ikoEpvaMJ17AjtVNtP3W/cftywGUJJDqpadIE5v12+1YlgBY+GIQk/y
f4++fu9Dgg3viSc9wVJLDWFkc2JJGQJiGbCYpy6UqWLMO5FA1jrpIM36efxr4a+1
+QBHVvWtVArbDFgthYq/Dn3mt8de6t3ut/jXHmKmjKpmcWP00ooXNPOc97xyYP2Q
FYWoDysjVj/ChgBKAv3SPbfsoY4EC1dJt0wpw93suXhNM53wd6jhF0vJRTLDcXKv
/+ObYH2jzxLj/fCr2DS8qsDSnMONItRYTqlq07yFDIWsCXHQhysAutsuFFtr1S/L
lu3Twcr/MF/j2vtLyhECqKPmWbH2etUTJohr2QPyAQ0qvsG9w1Fkp0CWFKDSJ3P2
idV1FQVxcD48NvESxn0isjFvs2V34NUwm0S3ptZvT4Ir9N2r5js9bqQVDd9e3V6A
rJClA5dbSB56DjJ0pQqlYPrtW/FCj91AFAkfi1w7ufqVG9TpSUAf1EqHtLNY9DJn
N1KNdhN/daw65NEDsPwemV3CS1dmIvvp/Upc2n34U3aPFewdnuaTuzF6lB8lafFz
UNKrBkLHIYsgGO6BAy9CQWnp4cciSHsVUZEmdk7LYIT/4G45QutVHYR5+2bgh30F
bDp4zEBe5zDVfOnN54QV5n3db1cHxxfKS5i7FC6WI3TmfGYaN4fCnNL0+GyocXQb
iBrtsn8M8Ij2d4TnQJ2/79sTS4Dtc//aVK2h1TB7RcshxumFyYYnkfI0JYqHqYvi
7meulgg+pZx5ZZUZzpNrOjcWRP7nvwkBW/5BdD9bntnvEIt+bUhxcxUOL7OAsXTh
9Cyv002Q6u2uG8HJtq9kkk21UtzoLxVAW2zBLInqLthA5yEHlK+ljgghoEssG/ux
XEbsMZXwKkzX3hC4eKOz/l5ND9v42dmhdNzv8F7Ao0q4VNAGvSYGvK/FK9aWuPuC
+fTATG/QsHDq3WTNYKqSCn5w88JZ78/91CXA1oBAsbJDdtjrDDrhGE9+Npuv7gQm
NhrQQcXCVjhGhKa3yHcGTX8k4Xkuxphq4gxZKpX5pzLn7ngS6QWiairnDoZiEc9R
uv2rd3RuOoMBKfX/5prVZL7ubUOAKkLCLPVUGh0w9QQ/2OjPDxIYYeB4bXB22fM3
F7nXzsr0E3QxLf8ZqI5IsSdSJg6sK7l3VkIrOEpROjrB1ssltoT88AHMoR8K4LOh
Doa9oioLIe1aZLDDNZbYkLbjxRqAXrNT2c3TnWoZOD+asQW/zP1Fc+sAoDI8EDol
NzXyMydHoBzOg1ilARhxbYTKO3VfJciv7NAyc6sRxUlT+N74cwcawOeKrZOD5y7U
fYPeIAZbpeeUyVGBfnlrPSlch6OyTDJZQVDffzvQnZyZWgiNn5iTXUV4wJ4dvSDn
ALeXXlAIPfI25PpapY6ZE961VtR2rqb9TkNCQ9TNY953FqHNVdF+fTYY2jLN6yD6
GxoZ4u4UbUGZhwtzTv/p2QgqNMYv65fHS8nmLDeFVOpVmii6Jd7qzNMhMtd84zYG
KCMGAYiaF8SY+3b9+bGAgMubpQCEjEhAvuIpJD6/z1UaYWrmzpfNR2NShXPoK9Mo
7zAgkCcOHTVuIc62jqquiEr2+1wRKe+Nc6Su7UQStzAB/zyF386U6/0XGf5wvvUe
JC146vAch6zYJzgMaiABR5y5p8k4ZPkPQ+K2y5lTStqIyQvM9xX7h6h6cQE77P2u
QX4dxlPbCvbBNxlML0PZhh1KdLX5R4nYFtmGSP8zLZ5lJOe0W89AA7itu9/CvV0u
OcviD3HY+nJtNjR1X0W82ZYqXmgB12bPymWaWLwBqX6cpf9cgoFeWgydyoDGCWDM
Fu90TU6+aVtsKchu61gqnvrY15P89YyzIe8e+QCuEzWuzGFEeE5HQkZnmK4AU3Kv
+ItPWCnJfrzdVXtcm599BPp50c224wPxo2pDjTi3a3UHGPwcaLqoYho60dlPoBqD
VwHUq6Dq7IGQqp092GbYOEiUQAtbbYP1O+VXD4EFc8RRrmu4DDVDl6c6sDWTpUZX
MN4AUr+HxBK8jG9JqOKa4d/AjkYqxJvq5GtBa0fdho4UVetEgnj/KLXJLUTflebJ
arl2rDSr4N85YUziLt8y1ltZBaUSk6hKYYLuccsVcUi3GAHyRi4u/u25Abo7WCKY
Aa97W6Y8PQq79tpfuQqqekS5e8Ii6Xs8Mr0v7J6usQQWatmazi8cB3x0VGZnLRm5
feT95h29Cti57jNb6Kycfy/S0JruHPp6rV7xrquyK47y0XWV2VIO1aCtVVr9fac3
vVEVB+b8LZPM93QoIyEWNICAGBBtQ50ISGi0rqgWtivEp2fdRA5AkALVD8JRNinB
GeOVeAyIQkTPwqCmM69g7FMXxN/1VYyHraRHQiXegBQeUNZjS66NE2p2tnwryz9m
XyXBKtjiXQYyqV6f4XhgG9c9i5CsRsWLH8P5lJMQZmUf8SpdK8MPzk0zYNDMqJ4k
FOZTRIj6kchhR4mSmaPqvAM1cMcQRGYSZSydMUC0sx5yxr5p+lNXVXmwJrawnwAE
BNvnIC+nMqVD3xYkeqk+DEj2bUNEf8Zni5+g18c7kS7EIBDReYRYXRhU6LLBapVe
b87168gJC4rXDIm8VE0og2dH7eWaJGPlGk/InuP11gPP/ayLYJJUbNGxupppu02Z
UeslWcUdtZ7NGsp1v7ADwOxPefRAL/6epHxWYAbN8YmdEB7u2czxGxMF1QursUPT
fXPIn6r6TBGOZaviX78kIa03eO0HzSnIMeeBhXD5mzzZ2963Dzd4PzuhI26xC7TD
ngMd9zHFVzjFG3HzTUYOYH1jMMZm/p57aLDCDlKEao/oPjhvoAJm51tNawgdmOi/
Oi7BzTLgvwMu2WBXJG6n/btf01pfR/GvSEVCumrTIWJIaybMFT6BHKTMn0J6l0eg
GT1VjeodqvYCLuoW8hI7uuPNK+PLyIBmub1TNell/VzMkgmDD/L5hP2DH0xYYHvY
cqFIfBHDN4+l//54YyJaSk6w1X0mN7vTRmJEGXOP92v60yjGqX9WBhQ6MLOrc5hA
fo5fpj1op60VB0fZFZaPAps0CmJRDZqOB/YhYy/+ubRg/R84Yrt71eLZcyOavhzg
73fxWE8r5/2PIj1VlB70sQiFhmmNsVdNxUUaXrVLt77Tn8Y8e/+oYQ1yMYMiEQ3N
ox4qHeMgcfscHx5BVWZEOJVlGk+5XVGESoXX8JPmyQU2HkBGmmfXNGBwkVq+jQyM
Ga/OTV4KOmLpFuPltXEdOrwNaue1Pg4lagz4E/sv5b6hDUhlk5dBIEXNC8/T1Gxh
UJBEgDiiwDK7peEPqrjyTa2Vsq+3zKQM8ue0y3b/Uc6G1NYa2+fwAgGmO+u8Hdbr
nQrAzpSHQHpHGUJzf9WB4BxnPE6qwGFvdJX30aMo3E/d9st5xB5zeKS1mlaxrhG0
YITisaXlCYRHJcKvQrhTA/bUs7OpqgcxfwHynIX+dzl8Rs4x4yuWFatsmoxnliEQ
XZIw1ZU92P0Tv32hOrfWfz3U/+EBKQAiBRJzqvdSNhvaDS9zJCt9Y20v7t2hA2q9
fOYueoyWapH9vFWNlod1Hg+cI4wUBamNuDnrxyj8Z25ln47RKQD2goCeLUi4ej/b
jKeeaoiyrRffewjMNm+IDKVo9FNy475GQtgii5mjX6slgdR3612HHEPHZ5mzFw2U
I4LRRrY12xDXKnPXHjdQbkxt60RZwTP9OUeRPcOUCjzIdOePhXMX9srPbsyIoDWV
EVTjGTnr9GxMTGzRzjmUkYUGToDoWLeiLical4e2ne2xPkgk4J0islEdu+dHgOqB
xfvHwLayZdz3aHRQp+hcmIrSRSc5RrYgj2rI++wOl+6kOpP+NIwSS/T4VXTH1tZ6
KFmxtBoQpJvA3D8vF92RcBdudW+U5+bI/FXKniMRRczJXJLqLj8KRdnyUQeU9IN6
IqzbXYy5O8fj6iSApj/0C0r0ZfraHKYFRCcX54Fj/4ZaH3Aq+863Ee7VLeI+anIT
4PNzM5VshzSOtAd2/6GRbjgpoWdKAZLvzNxkcYAD5DBKBc8iiOwRwzWE/MwYuTxf
RDWh786i4J6VgpoC/qkqex7LsLfqW0ptzGBzNjvQWbohD8CjrGRCTkkiAR03FBfU
W3ecpS3fbWNpTH20Mnx/3fXEocHrZBh4Y7QDP58QggUTtPFxjwP9ecbKa8wm7R5L
vgjTYFxBKK0InAtJ5UNYtKbymdAi3GDby9gZ7ePVAWRfnzN9elNFTZldwkAfQHrg
WYxZxxyolqeAV8M+3JvcQdfVVUxKjKCwJ9Lbviz+ntE/THmtk6y7ZWRA2H9yasTA
Gf6w+3rzOf0yFVdY2JxJGwCkeylp7sJ+6d1TUUElGxmeFmHm+Pq7ggYXDnpuYWMN
vuNaR1hDpC/ss/epvSPBkSv61GTpdKO9MD/ItY1i418VTP/1JNy72Krp2q8IgIIA
C08+ncrEbLkR+UekYgLe3bjRkRokunMWw5tpycOSw3iFBNxn3smfOnEfuzqJLUbR
CBhh326/8HuclL4KV1vXJ5Wm1I4GY+jJMS3c4IL9L3BHecgxS3GclT47b9FB86z5
jjskrbTAOcOTliYPg/GHyzphzZH1k5YIxeSeiGoFmp14BICLwDVnBkzj+jSVlriL
/OiT23bxORYZGfXCSDNKQ/rGOvgbekFcfdSyS13OhTY/RBEhCriz34+NRFFP5qCL
9OCrX/QQJzk7N2uh5/WBgjS7jy4VdImvPI6f/mBbEiPfJt7DkQWFJ4wodh3tf91B
DJ68ZoO1kySG1mozv8+OEL/VjnfbTlH5ColWRG18wZQuI3/WkUp6r/q0j/WduVWn
TNhuUpJMNbshOHo17cqiT5L4hLHYm3JxFtWWqTn/mfTZ5WPgt9Lir64+ZtBLGEVY
rcFbJv7d2f1LBiiE70SoQiemOTsxW+JYFyctKE8+7YJ9ntOfdl9FQlJabW1RTffS
8qWQXkgfg1Fhc3azUL8pdzMLgdV1Lp3/b5B5Eh2iM8eLXBOwWyxFRayAtV9UzA9N
cpcZz39HzvLBIPwN7f/bSrcxK2hw6a5KPBnMOoEVKoADekI0Ns4Ab8kglI60n9Xt
fXi7ffQNws9b7P6s+qxYbDwWqI1C+NrbbFY4nSaE7wN/YCUHFA60FwlaYyjGUYQM
q1i6/qofQyYM5eF8j8zBaMKGPZcZyEIDLLlPmk6nW8SJYaT0yUWfgTfLeyHnp/Ic
acwscse3fvaPMGix+rWnK5+Qbjz3YRBseDAF4OLrlTDS0sZyUGlvfi5X2rFCefqt
7V+n6vZQxChNjKLbIGJ5L9SL4ojXne5dXy5TWrgamZ26g3aOqjyCCjuT/Q3IRwtP
FXCYjEvoustb8YBCAJIp5OPzf7ZJIGF5Rl1SXMgjtbRqT5RYZq1ne5mpua1PHWrd
qloKgKEeD5oX+xZC7O+hRYac/SeEfic++grWFOG2psQUbFreA/oV+z5OR/Rpv4GO
LrgQ1M4CGFdyG6UdOp4YY1Dm+dwZDbmMLTd17PbZBJxYnbtb/uNaiMd2mmEjVX4u
qMK5PXpzhejgM8y6gyVPh8/WES4hJRXb7DJhYCr+MhISDQ0a8f03UVeodtnb47kw
BxdCfkxMdu4Ed73HFGXcJrsu7iEG0mp9fSygXrGR1649S38tJVQ/wGwj4dswdVYj
VVM6+aEizwhEAo/nj70eZb9G3ZYI2h9yyDMeyncU545Nyd/6srYqlWir9tW++ijE
AfO/3pUu6Cves/m+xC3rHjSD3LblsAtwB/269/hgJ+9Jq3EB5FXn7dTfFkSfumuA
XW59Bf51BVBNwFdeRFZOzL6SJ29lQ749Qy16HEv+wQh0fx2+9WBes9H3W/r2ohNm
4McPO9hSn6KqLFuEYymclhqpg1SXr6iUqucfnZw4vXCz2lc8ca3Pb1jDqVUtmhKj
+Pqapw6sc1fn7tl1P8xRD17oeyLpCEtd3WfnaIhqepyJ1zQqIfl/Hj8KwIr5RM/C
kNoVlLG1NxGiYbujR++P/CzFDfacznp86Ky9/3ObSJ+5fiphJlazR6+x5VcmQde1
1n/zx8BCLMQC43v5tvS9E6Q9wPc32le7OKyYz6s4BckL53WPrEXpEOIli36Ooih0
d+FtbxjGr5F4dhT7e+v+pAnqgNekMarZ27H8mn6EjWawjO3mK2cDnzmgk++WfXtM
FQebOpNWb5sg5Fzp913HXMnsJh0C6xDNnaAE2yq7Ny+WemcV56nGOUkM0owXf5za
Omrf8sQdbk8WhATFyzdCKCZCQnWAQdzd6dusHemRKasHByzce6DtEO+Typsq+I7t
vObL+tiW372eYaxXU2jsobmSWHPHyDx48DzsilS+L5AAuMzZazJtdiREOEb64eVW
ynp/gqzf8O0omBnB543cJKdBT4FEXp9T/1Y5GkkPEmiHneZSY33TOIOMZ57iT4QP
GNKswhsZ2kTaKCjMCRfNoLo1/JZLZv2dSYcjYeMR6Rtf4JTGIemi/DQCy9Jt15NF
AYmMTcCsztJTjcW2axncYgpp/d5vLQxyg/jmAczKEnbm7wKr2V6KYJG3zyepMvR8
i4HxiD5m2wfRH11pc0Zp4AZPaGkFEFsp2hc1Zc8joeui3Wef2xYfH6Ej2jUYowB6
tDyt8VRZdnOpLqwqM8RCMFRlGfv9JK8E+MB3Qmw+8uMWKCsMyluvAQhItwmSXIrB
5agcoIDwGuXf9Cfa4yPOGKgpTo20sdZWlS4hZLhoGhqGUqr0pOkLOGMvnZJqyTMI
ca4HPNmqZMS84EmFxQ88q21aXcIPaDv/d83GPrTrZM78uyUww1UGkHAKRZEboveY
RHfKfC6w0t5hkJUrcB5lL22HjPvoubMA1VTJKWtFezaB6DwPhaTF0a7rpsen5LOQ
+95F/KX+wrekon8OWC/HII6l++2VTeK+oyatZP+HZ+MTWokEV7RjXZxVdLw+rJ1Y
OxBZ03Kr957PHaZ9Q4yrLf9Btnmi/oNjJxTz3NcSQIvQ8FLmFCtOQypyV3BF2CEQ
e16phSFUCaQuXdT51F3hfWcqWmCF8VX5iPCsQLqaTUMcflx5QCtEBdsFSmiys7cc
uYCVExskFZtkyuPCY/MxneNyAOSERMam82sG/5pw1RrPX4l1KLAoWcU6F1DCfL4i
PPQQvKM5kIg9e6SfPHYnC4SOzGCwmOv9RUnL5greIAkC5LTDM3Lrv3Qv3g8+P/M7
CRdvwEn4/40yZlkHuLxrWBLXANDNiuHv/6q8Gvktcop/mwoVsXBO6Xw0RxEvVyV4
W3DNu8QCUFg4eOgJOZoGc6hHU4T2kx1s77nRIAQUWbKcKUgllODQ6mjOhioPGpFP
9ldq0dWgX8a36oVwnkmcHyB2H7RFo46oL5XH03K5pkQ9bv6KyLCj7es8SzKDkaW6
iE3u+1Ob4igvOFLF+2nDPpT/Np3O0ZI7yujTJh85W4+zfniQygGzzfgzVl8H3dK5
BvBRTiIy6cGGNeUFFyee7cY873gsw95NjhgIHcEajVsarHgZlmbkoWKMr2qMgZSi
vgxen/N9bjUIt60qlR/mcUCKJVcu9u73b1UCwmnsEhuAcHuSCtZoAl+uXwq18oIP
LLCt4yTVmpSPkkVjYYXsTpMe23bohIO3MUa4LRCod1x5CFmZWdSBlN81edDTbBeN
dw1YXg/BPa6WnTJvzExHd5AqnHcUTSRo2czrD318Pn8CaMag4EnowMmwdkL+pNLd
3QIDfxeTKjXYZzGLfUuqX1NAp2qT9cpIM+ThAW+I5Q4UaKcAvPKeGhwGfNYO7+ZD
wZ0oguNeQYeJ9LHH1ymFthidhu74KkyPb0upAm/8Jl/uf8xMw6nMjSj6GbrR/ZVA
Lpr1d997L3XNyke9tIFvGRln1PXIgKcpu3Ww6fLg2czqObCdLU+ytEJL1GYauifj
/bGs2qaWMDmoeCvypv8hMKC3f98MoX8rhYn/P/IDUgoaGGtX+m7Nklmam4zmHF1Z
qqf0Az8wxRP8jGGuE5MEpOBnvI5+QOdqNInROPoRa/E7z8Zhn6XjrwHomlEjaTDt
ufmrAOl3B0wMysBAkd+PRI1otLGQsqpir4HJpeTR8TSwlZivxTN4ehgGMtdN6xr3
+v6MGFbfaYP1CC5LCq81PdA19R6SXMxirqz9bgbT1DSJ9OBP9IAjMt25ZqZug8Fc
n51CgUumVUrllZkDEOzQIq+oqBBcEd/vTSMx1SsnSzsDYU9foNX/swsaBJlviUhH
j9AKt3CCRzLmxeYHP9kocZIxcgv6Q+EbNPsVwCXvMK5clGnBDAOhM2ddd+V6c+Bv
YuAj7ZI5XvfDHbbPyD76IKdzpbExz3SLex4R16X+MFYVuAg182qHPrD21YUXkNs9
0Vy3z/1CQwuZyehg7HLLsdhlMZwgdz99JIvZ3ZyK0oMEgr5Ew3giaG8mlxiwYVQE
7KyPb5QjpI655eBVdE3w/H0rh5pa8wyFOwbWoERONSw8Yi46bsibobAgVp8TqWCV
cLeTdBYjsEeA8BWCwcOwFxYGs89fAvnKYECDBv5OJ4gzWQ1pMpfF7AIFypnJ3NPM
4NvwWmbgl0NBk22y1LySbVJ+bjYvmJpWDPWxRUcKRynGADAW+ml0HAh1T5F4jISk
jfItrnDscYIotm9wWorsHdT8zy+lxB6Hr4kXphEm3eG0JCNgAxRj4VenDCCUFxjZ
IhQs5OXhD5GBjXeCGFYOGhCDLT31RO/tiLyqym2Q37ufFPfD9AH+PwQNoDYQpDo5
TkSDxgiQ6AhogAetSrvelCZpt/JxTL4X38MtfQ2BSCl+YbvSfDfqWLnwiPNag1OK
ttmLlg5Sen+Jlavn01boebo/gJPz9Vgeqkrxn8Phi5f2lDoxx1vTXkJgp7lrQrZI
ZTErXgSti6t6M5/KGPKd8Stfwr8pCVQomOzkLxivNpAC/ZC0E0kpWD5okwx3woAb
JC2cBTeoeUke6DErjykDGpiZPXlIVPgp4gyxSiZBGd/7Htbt/OcWrpuNROSfiY30
/9NjDLsuyB68WauGjk7GHWUdheJZxnN61v8NniqHerWBnpSXfdUIeOsfDwV82g9Z
OYV83NAyFp37iDqI5L4f7E6EW2U9EsLa3OGTFCLsDRjNERwsl+xQCNGyd06OH9sP
FDhFuksglUf5DpuerEbx+lEfwOTxzmZ/9kuamDJNwK4EoUNYtMGWw6I7pj4I4fIR
RZZw+OKFXomtVU1HR9lTKMT0zmxYNQQw197NNSMV+3PnRkMCu9xNxYRSC32WyVTg
dsfc3WQn7U66aIAgmU2tTLno6qQIOzSWzLQ6/HjLfwrS/i/dIyEyIjhJz39CVs2i
R7tfvtT8p0hhsb5kGwgaYvKwJqo8JFFNuzpdOTnUBxAnBlYwhy+gaUyD38FzIZYM
mx3fSjmpOMLxRJS3xwWz/KoArQ7o9sFC60sdPE0dfw3kam1EwolsAVIszSnyh579
+JGmADPr85PoMRJ3UijZvkuVJCEOwL3P7L/I9DEP0ptyjU7vD/5+oi3JMWV9p1GL
K/LsU+kFPiFJ5x40vWCB2Xc5EYOwFfhkZcxzBN93v5ay7VFZx4xjI9QTmPX3pYhc
sugTOuikrewYuXoHnm3z1p9UHppbU264Wf249NslRgV3FleWKF0wG2YHrqxjBeXw
d+5grXcx5tEbiYyH+HOG8VWVfk/oHzbeGh05w5WlEuSyl9TmyI3tJ39IMyRop+eO
7BycI9szjkQ6UyATT430G5SEI6TdGS5q5FpwRsJ3wzvkFSk4FKAygLdGFUD+yLa4
LcUolLR6kErmJicxwtKjEfYlPv3vBYOQ4hJerwjFXtI7RIgA+7aAgwDwGvI4uFhy
+DzEnS/i1o4RRTTCn09gfSvi8drNRyVY5bRWPmpJ/ImPXnjERWmYAH85S3C0gSAu
e8HRgwhofAyzeRkMmOTrERxrFtVuhKAzQHxwiC/hJ+kKKymcRn3lKBSfAouULfXL
T53pFBPZ3B9rd01Ux4R8TWFw1rRUpA3e8c09w35hjQKYVy4JaswVhcu1ru39CQuG
vlNbSxZTdMHq1+J9JjFeKjY+zGoR5LSXMn5pRfe+RZW9JN+6pQx9d96NliZNxTss
VTikgwymgiynWZXkdUEtEBLlwHvAYQ/XlWg6DL42QZVdPZaaowdksFg1wq2G5ULe
J5wyChSPqFi5NiAuwT6pzwxSIKcFdDKIeIr6y2LUacR54Gn6AsGSlBGnTOj7Gtt1
dxnjYoIkHMsnlg1CfgTHVHpbmwsiINJqUrvsq28izBC/ZBgPgYYIDZMO62nlCiR7
3zEL5lrzEyPILgRDGxPKiEzTW9L7KYsLaBl91n26j+5X2/AZ3p9xtJtwLH8uAKX3
wP47NdZ7PTMhGMuyXGtp3I/Xu7s2lpM1FG/J3FtHssurFWSFXirhQRoxkrTWVxla
+xp4zlIJDGgIEtP002EacApkegnb5aUH3CKRbRHm2abNKL/G5Xwv0kd84xsXjh6t
ur6NZQ06yp2gTVNJC+Mz5L+uWO9xc0VE+cZ4wtGixBpA/8VcWxQ8mONpSjlR0HBh
qzlU4m6Y+wIno/4JXZMzlWjBqCZieysGdF8JEQtzcGZOk/0p6fRT4JQyQ5DA4B4N
iyJdJZnzskPAHEjijia/mawl50GtHSFT2NjS5aj8NCvSDWGkSkonzTpHAKJGSkHr
V7JJtINPikFzeVrfWGbf/IIer49e7Fi46RM4aih4Uha3sg3Xv04xiZWH/pdv7wLm
XXRvnB3brvuxQtgVEyyJOxkc9RlUKGyjNtFIthRjhL81n47H6dp0MgQh/a+Cr4oS
GKjoORkCJaqZr3O9bpDIfzcRlyaQX7jAg0APT2Ku5Gqr6JsEaz7kPNjM6tHj6vHI
1lKFITNyDjNGn7JhK6lq4ZfOBVBCxH579Ouuz9QV49SxTILz0cWlRaA0t5lX9JaE
oyFGLjXWBiWK0o36IGiGdMSA6DubXFzrQSBPs97NALpJGUvW0eIdPSLmerJj3Gvj
I3MXCjcht2tOhrcGXfqx8t7NeNywERwI+eoU55Z6wxtliVYychYL/R5AoLvVKLuo
Y2ePqGjkgsjuZrLzp6884TlrTVZtBRLft9pOXFftCVXjU7QIR2meKKbEwLhJuvNY
immctfD54lDU/1aTxiCCYuznDDzfHkoIvz48hh1y/07pqGd2kUBXa9vO7rhpokIE
PFNt3KKJqc29+zIqlKlIQDmnefF0EVG3iYOqMPf6onlsxjVcWFOswEXUMrLH8iRH
R1dlKwGAfWdq6O1ZIbgEX1YZhs7KtRgSA5qh2wbdwAwH5hS7evdQEl7e5VXczQvq
g1i9Vtc0i9zy9MxmoPp95r5iHk4jX6bFWWXGUT0k9/KNznWfg6JxsSymDce3G22h
zs2IeHbIoK1DjselDs+gRqsV9u1iC3OiY/NdgxEG/LNAqDt1Ro56gIBWVqC82wp0
JcG6OQ5b2GLmoorEfvOg3BBv2lmUgGzJavyKmeegSG8XiB1g/ApbOtgSeeD7ehvF
pPMfPNMDH2ino0VKIDx7qdI9eL4u41Cy2o482O7liuRMD+60FrCHaJ2TxMVgAV+6
tJvWmstkt2qgakzikudWUBTsGoM1+YHpPgdpmz26Cf4yr5IyxPMoNrY/lFHo7zNf
qQLc3Ntvs+J0G+nrTVwJgd0qt3Wg9ICQBfYKlPzYt9MuDV9+GgWSLsjLreQ++FGE
c8ghRBlCAqoOgcg0i5OEoc8H2G5k9mta+e9foDIXR/+mwXZQ2JSqeWochcb+GJxh
2+hAvDFUL6HIp7GYM62MOpr7RvAyP4hM6m5RE1Q8QtC6mcYY0K/1BsSrlL7C8d+8
8j1fEZgt7lMfiEn6DMb0Z0dUCT8QCbJ9QYLSdAnOTWCRS/pn4cF+OA0mzBx85CND
bbYxhWOMqJrrG/2u8X2ykXZJm+X/glBCAko7JgXFFRZMqdbwDNgTWXk/2j5MKh/7
NVXtcv9imAi7e/gbSghvKOslnZ7uRGivtxQoZoQKCNqZEQMBBuy53ByjXUzjPU3i
Ut1ZAPkWf/j5ZjQc6mcDwOM0P0e5T/RRfJriey0tqykNxsrXSMAm7E40KQi3V+vI
jtUyvtrfOIjn87K0DiS72lTKOKp/OOw9XAyB1Gzyy2Esw2krs2dFNhgNPQST4BVT
95zUmwY+P0ALwc15FvIq8rcrk6ZTjxEEl06oVzbm0EGLOtGVM2HgbJtRxr2wU5BJ
x1Vlg9FU8y5Un4EpyU+C6qg/Pbx84qd/v0VJ/o14jH9YRIijzxnWBFORNL5uA0MF
1LwEuRlw6sN1LQnzmq6tAAXSsowWSfVEKSYWvDDK4SEoWnUAkl4IWy2wohMeEFU1
hJzaPG3zEBxy7MmXL2l/n2NR1DiZ17d6T6KsrbyizpJi+XAwMECgeTFq4j0FqF+1
Ia2CURK8L566WmNdjJrlBvTQhM20NcksV/p2b1chTxCBumhxTLM3GFdD/szqg2bX
4Bw3LgCYDVZI4m6N8cz5E2qBgTbZl3cuvbMc2klHvZnq9D0bD4qPDtPQkXzYSN1H
7N+JAcRnDHfLD+F6BiSUlpvj2W2h8LZamKze2Nzce0f7LLsoIvDUxpmZHfcjUXBl
a1LExnO5fB5uNJuNbn7DGJVCozXOsq8q46jHtcKji8MCt7aorGcSw7FXocwIfeZa
2G9hKUy+nNvIA0zSSI+jEMxO0Vk8Q85Zifju/nTkkow5yAWMV+Us5YSpssEG6IV5
P5wLqKoGcd3xwcXzl9ZGXZvfylzWOpNGAAjs6KJMGc/qQi4fpDUW5kJ7ObkMT1YY
ZTblpJYypIkD0t+DrIiJ1HsvKIkl6ktU7NSE/wF7oLe3JzwtJ64VFNzpXtlzX+yZ
jg5Bz3QE565TA7WvXkRK7Nx/PQFOq2pKJNK/wiMHc5v+HbXPA8OxyCFUVRE/WV4x
yo8/zAO0Tpun22HPmUOAWhXMw/Th47sXSPCiiHWP3Rj6UtdyRWkq+pxcM8ryhoRd
u0XFNqXtAZV/pL7oMXwKzy8VlqtdqSssg18Jaiwk4Cwn14xC0Wi+QhqdFN/cBReI
Z/ZovnLBlBl4e4PXJFxngSHURbwu4mN6E3CZtOLxgeBMD3fpW40GTSIPUtxbRGlQ
eIEQFyKUBEj/k6wy+XLr5hmjq9aI+h7sZCBEEFomXrJE4B5fUgNOlSsMb11SS+Gn
+nxEfW6luE7806QYXqlXgpOnU5/5ocx+D8EFuU4/Qn7+Y9KB4ND14TzL/8OYo4Sv
/ZRTPub/TvcyO92yBj+tzgGCFj9+Zks19u5vFApXx6EdZQ164cEbrli7bz9B3uy4
p7tb+kTyQK4o1ItiLQUgZpKhQCU6nH/Kg85Mo7L/CRgHdJlBuBN9TfTfwcqennaG
o77Xkgpvgv1rF6aG0NzT8VexsYiKMPjIUURJtOLVFO0LrrLfUruWRZa8VnLtmqom
J3SXXLl+8+nM7JoO6qgn8pipOF+QE5td9IqldbD6E5UbJTDUXcVTfSrgdLsVMJP7
2l2Pcyus+dYDLQo2EWOzkcD01ZbZKP1ZUPmGtqEVjsm4YvyNO7NsxBkCJOMKHIas
6Wgc0/ejAFgJEG3P4EGztKXrZjRqIWjnUyVjxJNnXeF/IFhm6BxzVHyGhqSUHZHh
RNPr0uqU5crfDyJDEAaH1gG8tg81u3p7AOont2uxAvqktf8q8Zu0tb6pO5SBVd31
7TgsnIlGodQkb9pYVSFzWTpx3BEcFXaTy/+KJRnWvSlhiej1r835jX8euQfZMxzw
RG45uU1ha+FeuCedOT5lphzTmD5sO9u1wYkto61KxJlksZDP1oIPx++M3iWtXjm+
WG+i4w4TaMt8mgvepHnYe1DpNxF+Km7+VQ18b2sx4DTbBBDMM0UG8cGXcjA/9HAD
f4dnMylLFyy+6vT+9KqBcUfHtQ7AITXzv0oBw+JXEZqLP5eLJmCRsBdakj7v6BMq
9thqyecjevEjfjorYqUfOvcA+pbEfIr6ELdQxxw3W97uMuYwZ4lJxpyTGkcbHEwL
EmZOp6I+txVkVKgZPNJiZ83Uz9R2/h1G6PmLELHVSuYeKfe/w6Ar9VH34C8Lhstb
Ya2rQ+TZGF+Jj/TqjXlbsmSpgpBOYLA9nt+njic/0+UqI0Sq5gjD7NWILtHwh6YM
onFSys+Xdt9pnxaIp2I0dwd5J33ib2+SBxA9AT/oLk2lDefH+0CIIEPlTwaPT9xG
NJMa2nGjRyWrASHHjKL+8TsbI+Pd1A7lNpZbuFFsRnKZJ1Hqwub/sUEgQKg4j10i
ECkAp7pNezcxzBt26D8f2sWeM7sKFdhqd2B+K3gxwWTMoLUDxIPPHhZivhzeJOr8
rkZTSoPeG4JYc7iyYz+1VgEy0bKsL/0+cIeZI2J1bqbhgXP1mfuhu1BCD4Zm8IEI
8UGzAjqr+0295M3MN4Hu0cMGC+fmRg8jz0sVN+IjyQwCJS00B0wBWhkjhfEYpFBQ
PAEInUpPL26mNe3KVuyGr0gGqhl5HkGbtCD6/XB5bytG6c+HlKxYhY9MkhJqv/c2
xBnbx4cnaOisVIYhttywn2tIc6LbKnN47VNgljCzUvwvjysTz/6L129A/st16hUy
Wa1A6GmxKcnUZKOADJE6yAByZRFHgaBXxlpNhhvF024QyUfn0XkjjT6XpqOmiV/r
MuDCMqnj67AUJQ6rMd7MykfsNn2f6ZXbweD5CbNnJkdkw8OR5SrHV8l6D3HRVhv+
aW9EHlgDgqFmh5FLv7LZLo0ALTnXc19UYBlOHz7CEz6olokfTG1ffXO8b4LpYHwh
2nW5IN8mNZszhwefTWPyfEkf7kN5xSxf6vuzEHMLk14tN9nL/Rq88/EvOuZWqIDb
JwzT3RXuw/PPrWvBuactbIySo1ISdTzSlN/sxTP4flx6+RW6Vi1ZmHhX5gCLchP8
nCT6zCKxniAaVoy/f9Olug+ReIRe5lD/V4tmW2upUbdy57dTOXOiWknzVyZzf8oP
ZU0wWsD24SQaMWrxUmPCYv/TJtbBEoipCb/cdCqLsNQHtxsOUZ+R9mwbIWLJufH4
A/gZApYJRoAGaG5mcF8ChgRd8UhG0TbA8+LC9m21m8VLn2HfJbUvAd/ugReaJ8TM
qH9+GgtQccvosHkBYPIY7iI2ryteLqNgpvIORQla83P7WkOK8o5P+c5xHvsImW68
BlvO7ouugHkNP9VwDXIjJsWTtfp1YC44tKuQ7NkX+D5SFV0Loq9QNpwqS34gCq2I
bvbIrwJlWeS6Wp4ldPMWR6GZrrvQc+NAWwLJO1mmtR7HzsDZDg4cLOm0mduxqRmH
+g8g6kkB3Ft9JBgCxO1IcE9AjQre0FlPfW6K9eUtgUnaCkQJ/yAcr7G2fIHBxyOn
kmr4EAqgYrYW81pVTSpmd9e6ABB3UPLiXe1PZR7M0JnKOlVR9mQN6wq/FJ+nH8+B
+4q8OoptYJOMe0HkCozj4pFSpA3VYh0/QY2eMTZqMjtyX+sIJTiIrrmjr/IhDskc
rHm9BPOEDskRA2LH+QYaSp8XYiaVHu+UyNdAkp60c/p+bmwgmjD46afXNo+Kj+fm
VuzEzlDAHxxWLS3dRPexSu8JKGkgvRHJo2Kso05Z7H1bCyOHHX5tGcHpdfULAJXu
8TZxLtlVTWoo12QrWmNsgfmzQ8W4cvuYIySAwdnUEQxO+LvSWE0ztgzDtBoZ4FUw
MFs1qik96KurhFztlhWrIIJZtb1mK2lSq6NRXG+ctlQOFX1oVZmF0B/3oCxM8k51
xtDvhoZnFUwQO+7Zdyq2qnKNRkmvJTRrIgMGJNZfv8/pJEx68RmIqIdXw0vbjRqU
Bdn936QRqiaAjrtRmZf2ZT0xzToKb4azcKzNtDkZBMrLeS9EYeLqGszg0ZuSX4G/
SYVPYTUPzORx4RfMg5PI13p7K+g1YUNeQqb+LldVvlB9vJ+Wgvh0DvGzl+8CmbrN
skn0DFHSQTAMrNPPA3Q4USBOaNjR/VNQ0HZycBxWUK59IKQMy7wpwJFhYuA1Ffov
/x/bGyM7cv0JwdEk3T/SPjDHjc3BbOxgUNO/SHd681vAkyxHsYeHIfw8LvLqFzQG
Lthxz2uvrnto++AS/pU+8dh+eyi3UyFyT3aCDY764xd3RHZLee0ZMI5wWfWffR5h
nyU4CClmAawZZ+GAnzEuofGNImtR99alvzUwows4EFLI04bVNxDSoWCi8iDpfHYd
rPMzcqlzWZ5F6oGIM/pP6NgxpJnOKoyXnq0+ZpdvqY/xs8/0TC33+HLkoASK0I1w
e5812/0ttWUPWqxYpAMToCFfdyBQ5RIpt11IYFta9TIrxmMorr77Se3oKQAUzgVf
B18OKO3aYzRf6UVS4/Qj0vFSifI60l2VStYyt/RfWbySaCKvWXLdiz1xVtSq632o
xOQaDr1UDOIcwPfqr9jL4ttzf4L7IMluQvdvyhun7OpKfcOHJvABgz8FOpJb/vmQ
1E9wbkHxuYcKDBasJHabd4E1WQ/+hWtVV3iXFYsqEFOBbTUliZaA+A5hnCGTJCFe
6b57MwQsC6ZluBz57zXd+g/n84tpCLNrmCnQsJ34jhOtL+qvM/9ogNB0hHMKC590
TcXZQTnRQQaYCBDYrVHg2XXrmVZJ8V8MNeRTI+jDEC8tPpyfmkOSvqXfvv/pHYDV
p+KE6Qyg4w3mhyY55w8kY/c+J+1SzMUK5y5i+91ykCYUai5cpYqgw2lhCnbcN5gC
VSsUU17G/VvPIqoMarYC1x+arHAp4q4p7qWpH90OhEGpenKJFj1gMIyvYfGtR2Sn
yvP2t6NFmRnlMFPkhGlqRl15PMIyVbF30Zxbo6rNBOCqaLb6D6tzg7tia31bilyg
HV+VMDzAuiNqnSZs5toRM7oVP2RbNmdI7rZLupbebLD8FA0EYERWJ1U39J9WC0g1
XNb0MUaQo26/irqHuRAmxG/PgPYDnVz+GXUzT/XKTldGf62ebC2xxTtAO47AbKbH
PVilIsNIsQcFIuQsuQTPPQXQkHdR9l0HD/78hzxFN1HpHhQ00qoiqZVDZSFqNfq2
EygbLUa8YIhNGDuFKO8qxiAAsgYPD/bKU8+44fFr7318540tpsFIZw6BA4qTK37Z
O/ABVRWrRMKCxDz46RaclWPGrrbIOw6RRmUt1j0afDc4Ye9vW0LkJ597sjhftYYh
I/kbcvjN38sdcRIFzneNCT/lv83X/yW3dDc8IQqAwwk5DwFbpSFTy6BeqEOtupgK
q6dzYp5MTnz+gzNwteRkmjJ5RdtUEM0ISQckx6aslopA0J3sMDfxWP/A9FVSw5E/
RWxjx46LDEYGjFFQdUM0Z2rOthOQNegZnP/D8AaxW2tFkwHG+LawPnWmHYTY6/Qx
dNGKfAL0g14xyALcF4rTH9NOcl/tQMGMk5TXqvIYvwYb/7004fkxjY10MN9QoLNZ
1FefcWDeHpdMh0QjreXDBvXEGcfB5D5c9gBhmg/KpZWh0/HJO/itqwmSBrWPmmGP
/ovAM6J3d9XTEVi2jv8MzfIgpkt5QYfZcTxVpBhyJFh581qnzkvtFcKQ/Zkt8JLY
xefrgw6FNDamxh7Sq1KNrqWxPq+lxSsx4F1SW1TU3az5EsyYVmD5kmk9FFnD7oT2
OlXtKxEsYGbijxYCUcYMPL2bjlbF9zojS0MYlZCI/ZHw/InaqyDax11t2SclUoVb
QsrrK5JesoP5R9YVUS/eAWT/g9XYIQVKWWWj4PHMli8XKIRkt29wtKIjywPCywkp
lxNL2/rG7Aq6uZRPu1Z/qPyBvhFB6+EQyFklHN4ZHX8DVyMHc1poFgpHICwFIUMe
faO3jfCW62zIXewk7EiySrgtchfPIgPYo0bgJibvsIWlKGJ8qvTAocnZc7edqi4V
6bMX+5Kn/oHFwljTK1GjhCfHtLKam3XxFBHyXaLDVgTZHVwT5GbIpQexauZGMO0Z
lfQnZpVylogQ4tM/6pKZGNOGM2qM4Kh3AmnukQWcRWfOaCqZ4FXm1PAvFlydVmJ0
A580itbpGo/5obcuKQH2wPkRDEHobStQjjyHzgS4wztEOHVksGw4VgEvcpLqyHzf
I6gujvly4/pWPHlFXc0uwulOZS5bcCJt2yDNKSc4sImp/5XvLZLOgPyRfez0NvKD
r7iMU/kgcq+dqG/m/HGAwkOjX5b657XNB49Uoy1lQGUAvFPacEHAAUgDgBt9YTLD
sWIQfoSktGCX7t6cBt6fazPfkE+m1almGtVohQncJdFJ0WlerVlvYU9504/izhRQ
rSqFczViRUTO6j+2mk5PJXHk0D65hdgGif9MBv+QuRzZJzNBnxFT/SCKgA8UEnXP
rrpysO8CwqvcNfCiEDJatKjYoLEnBoQt/kBg9gcwTEzKhVVZyyATpZHVbxcyEXgY
tyJKRd0AdSzE+q23cHV8rJ70UGnZOIL2VldJq2I2EU+kWnlAL5FJ+/CgTRwUCl7q
QbBoEVgckUMeNvfTYmkf5rbC0nk3lxmceuD/MuI1b18P3klB/+S5dp2/y5+6alGM
A4iSHd7o9lfWnfnG18Nrkdr7yL+p0PRTFFwZoTLSd+zs4TZ+eAVCGRCtkQ1LN9a+
f1HC7hjHuva86u7L/Xc8xiBe5YddOdDSevlxjHnkiWOSOdnP8hS7OYdaxnkatP11
YRkn3lS8/1KECcB0OgNeHTuQsAMsgKHhBl45+RCfJCPFy9jJkUF76Tcl7a+akhf/
fxpI+uX4A56P6w83rNv5Hk77ExG1ACVn0DPxiqhCvEWpzQM5u62AYuJoE7Cees+l
Fhqb9+m9M8UZkNlwQVMED3vot83r0EGnr3RxaBKTr7KeNbBqz/iW0RwQlpD43iXw
uva1nsjWV/R4MNYMFyZIT3QydUGdSk7Z5oIwvVZ5xF3wIq9Nonc9VjTqjcpbqwpb
wSA+9Jgu4P4PQC1ZiboYPvVzumRh2xP9buqEE03QkecElRRHvHkSt7zy5fJ+kGbg
UsF2qKXVdOQsnV6XMcFATz2esRzelTySh/IC8QDbITzsFZaKeLargYWBlZVX2Zcb
hwVGJBGuopeo3nsS/HQRPrdLqXnrWiiQK8eRLbc0qY+7nK1H/3lfXxbERqQehDi/
wbmEhi5hmMj1LKNFvIWv5m/rb+iDQY52vzTZcc8jkqQWdpN8cjn/AeIbX9XJxoDA
VDRLc0XLUMyk85j7ijKwjZd0FokUA1gYeR337LqeCoigj2DR/9Yy+nxYpSvsmL75
BP4itl1C2HXg3ykBy5kM40tnmOe6hD307hrGs4cUbJ4YqyTduCWPWBLpuxBq5d5l
YyBJ6ZcoctcEJAiJPxI51l8gHnzVEPlRNkdx9D+9CNwbPCHSK4q97ImqGs27Aml6
tLP6smCcaIlIv1rP/VkImAwr2t9eW2q6usIyHC90+r9AYgu56ggD3plIBPVAB2oT
PjK+iK8FwEkgEzagzEAwOunk376DNKvAg8UJVWhdZ5lkPqZ6bc2h2L/Te9y5QRcv
/iJMnM2OGgHaeTzHz80V5YIBQRViQOaLGM1nq5WxD1/LNVMqxbfD0mF3TUSFaKOa
VXQgK/LLHNbUMiriiuF0iedE6CNQIkuZSX4y6E/tNl5LNnl5Wa9JjbPt/XF0LOsf
xyg1iKBnWX7aeq7UGUJwn3/V18GvYxxDxqPUkjiyOA4ff+HMNiCQb8DVLL0dITAP
o4fRYoiCK8A3EXRO1FBCYfYRKwAxThMzcmflXlj7rQxx4DANjCBUCBll2PRkjrLE
UTKokS0XDPO+5zLTclSStoF7RBk/0i5M0iFr5j+3bqw85RQzbjkqGMwbji45gCeT
BjTQZY5x+fVmPpcYvlXuY1PuO8C9yo5LPycVOUW9H6f3kNifvYjRv0b/t6DV8vi8
wX+HbMD1KnSxCdEe+45qKvhTzbWqKFme86xTEZiH38HhfYj3l787ulNUudQAyvk4
yuzEnd6h30BGMBGS2gVi9PcweB/IZdxX693tRkmU8hQoaoGSKmebNuU/hu0FYw3T
Cdx9Q+NFtmeESgZ9FwhardXuSgeLqt4f9FnViPaL5ICdlW2WM4kUgQkZkNOkyw8G
AXjdDWK3DbU7940ofag8Vjgg9EKAxNu2ghyxvCQB3YArZm1GwSYk37nQwX2LMP3K
xjvXexYf6TL857GMmoMprJnO0NAIkD73gs9H/avSEMEcQdaoJs63kr8aVJt19PNm
JIZ6wuKE/RfVAETJO7qTkG7EJZeGOcqw0Kc4sN6x0CfuWKQmeldtNhpwhX5SCo2H
NRHA1XaabmZEIiLHBZPCWJmGDorSbFFANIS0NHZr7tAZ4sj390OMFZtkRF7Gl5iU
/79EW6gWXuE1Ihhl8mqA47FkV1c5joL3yg7tQIBG3aTGnU9heO3AnQW4bULAQQ0I
Cm5I5oHVpSrG/Nexfj6X56Jjz5pRSPMcBXZ35HtGE6xg4uqjtoPkjaKXrsIr6cNX
9WYiirbgzqfoHaTW/miXSCFgN+oEjIerB/uP1gp1WiIS1kKDGqMXhOP2CoyJ9bv3
osd1zOipkDPrSsVaPGI/75npfuKlK1amGAp9nsCrTVctVZki8AzhToxNh5j9o6nb
h8DBVYHabgeUlyr3WyKa3eT+K37fQG4bcBHD2iI0obyUl5fxVlBs73aRy5tHR7Tn
maZ9C5emLfJ8iDzEwmYtNgqZPlSX6s9K1NGKl0jatveFZMn7c7zaKzlBhkW1/4vR
drImbzoOMQONZcHEDDOClonAbiLQCrEwWTO2m2l/hoe+4QjW35XxuZJEsuMOLqr5
1+mDt3KYLkfhc+llOdW+OLgE4c44rhaSg5GoKOgT5W6M8c0UDjabLiKemWdO4v4E
n52GU5vROuFFXX4Mep4V81rhRjn2rMzNVQlVsdU1BlIdyuOwf6Ms64dJA8jc35I9
PZJuDDocLHW/Z5NBYJl9bNBZGFv5/SWaegfWTCGlDsLNR7GGcgV7lAYFF9qKpZnF
TfGGZtQ/4/1fhlsp1tFtMlVHApMUnXWRoyK3lDMx7viDKUWuUgZ6OHnPCpARaNgH
3u3RJQDw0/coYvfNQPu4Gyp1b5WcpgKSgKJMU2LBAIzgm5rXM+dCcfSIrCTpDNHL
V6CeY1CdDgEMg9csMSpdYGXisSN97qNchZp+2ncQZm0ej/2WgUDpwnkkGVjVAxuF
fC93A4qhgLIiQebFVEVNoecfWqrcyVeYKLFixkJz3LTK0DJ0gwZNv9TYe/UO17S6
LxJSdK5ATftk4F4/bF9/Q7eeW4eJzH9169BijzzErKcL1kCmt9/gTwH7YDqWjuHX
iBtpglHWd/odUPJDbTTle4w063Ke1AtV0k2ewQbWHyRcSI3Ye5iV+A5v4OFdf2md
jvS2UgCCDEPfb48tWCdSabTJsFI85j7YB+RYCeadZExveBttaWe/pDd65Fnujtjh
+OSHUIzTmurFGA5Azedex4TCTP+FJiq3uvXxl9opYnmPceOcXCE98rj5rdrHtaKK
sA7IjPPudCsUoktYinoI+i9IKyZBZ73ygT5jdrhO5meMfRVTb5ILvrODCLhdAg1G
WHBsoLPFW5JdRVdMLWrAbJ8bn4nb3ppEMfVU+ie9BRGOY5tSxb0I4im/rpxbouKD
Tsi9VQ/LA+Jk/yKxDaH7MNV7jHluyzq/SaZtJFfbEw1ePAMuibXwptyntx3EvhJ/
pjKoFn4H5v0TosoJKvYCSpc4Gqg9v6oa1XwTWSr8FfkX39XxYlkLAJrDiLxDjspf
r/2Jl4dopc2NqNX9xloZ5VnC6bvLP1kWf86fm3L3307odN9Qku6w58+4LMH0Q7Rf
qOZXoUVM884riVcEAjSnSQgq+YGBX053bfcLJ8tL4ZCE5Nin6lK10q/VX7gb6Bkr
RHwi4RLRUjSa3gKg2Kq8BlOGY9qGzQqC+Vjol2wZTGclBUPxGprAS2oBIlqQRTl/
u+ccDCnjaJTmrOc8zzrMDdSd+vOxSU1reu2E6aWb1soolzwlSsmvYTVbmVYfwNat
J+XC7OuTEQrb3gAAvKpMi4fAPiqb/VASR3t0NSUfaIi9HhS9118/j57FQtRe4Pew
zEXULPiVpBMd3lDTXte/+ofwp9/NO1pj2wGt/YCVKXib1nG77HQ4FRgmwqIwDtWh
rMmKjIq+i+fFKbsD/1ip84g4XB2tsnvBEwWSQ1r7xn2I5obTgD3yJLH/JDReTtpO
Y7A6Mg5Hjg/mD+cbWm+MclBLHFQLqMwguA2bjbx0PzTwrfxnEfmUG5VepbMgCQbt
VFxoWM8U/V6aNrKZj56wZliL6nzPQBopKUuBGHf+6rVHXj0G5U2c8TGBDp1h6sxG
aUaw0VCHHXHTJ4zKVd/OZ9vURKnWn5b0CpvK7vMaKej7MONRS85w3+z6ZFtZ2sCu
t+QLx25iEUsScgOpXQpVbh8uxJVjhEEqwyjxdHqIQgmXQKgSth4sSt2ZyPM4bLAR
ghGrDygfFFljQ5cvSPx7U2ZGbgFqgAxT2fJgzRWmpL43i+W4GsTcRUKaeaUO5dUU
jIDL92EQ5T6JaDy5S/E688wqKIkbE6LpeIePrcsPkFxPGyZ65cxMnyJUU4niFb7x
5VH0/7FtoA1iSxOpmVCaK68aVllHotvM58vP/4kpmO7Pd9tZBnWgA78keYftZIJS
Q4hFX3zhOKjc2NSb6zCPzrd9A74U80xF+zEkQNTNWPVdKD4fhylA35VQ7ldor5yT
kyJELjquxh6LqqR0xAGVqyJ+voMyWEQrB+EPKNKXoq0IrO0faL7TWmLNWPbsqS4m
mpXKwTnO2mRUhKOv+Mod8loeJY+wE98yMuNKLYT7Nkzs3WhGAUXHOr1wPCTrpF0g
4lPpWMrnkf8EdH9fkKEhcGRFvu9Vi5RMQn1QuMjy/Y6/q74+Mh/jcSkdqv/yLAKs
+Bv5qCyk9+BOh3zGnAiZdBd1xCV5+JPytQLXXGSw30qGG1ZFfyhg2lftLBJQk1Jn
g88qtim93LTOdJb20+B2UVlbOKS93Mxh52gqy76oRkMAaDjzQOV1OkihK1yLUKTL
5L0/th8AraEAtizftCLCwnH++S5/oiEc1+Knx8ngklQeaqHq9Cm0jJ4uKyI10TO9
Im8HCTUsWQ/wTjOiQdhkmYmyeIfuMJekiEqCVSuZ7tp7ViDLh+GHMY9xDKG2EpF5
dk5idyKeFufF7sCMme+l45DTvzCpB3NAUTrxx4GJ8iIiGidbuuxOL8mEy4+tDad+
s2AZAMNu65sSHt0Ss731XijtnvIJou2TYZmtogZfyTgv5WsnZ31Kub72kyYoDSxZ
GohCvD4bMZEZj83KwIJD+5fNZK/4vARl8sFVZaWbqohd5NQL1d5Z4o4Z8MdZT+df
Zl1po8XTzgO0Upusau2zk1f2UZTLzPgGp5tU4Kt5o+st6mA/77e7eV5hc0sGG0FY
gu1QKQRmNbL1ODGyu+KLARSLTUPeYAbC6o5YnVdx5B4UmFyWWTtRG/KPrlGAHEKs
Bz+oWJHj8uwUkK0qN0MRJNgHZjaiPew8nnUrg/0pl8mCr5EOX7J4zTYQirsKv0m6
KGs61kHd+6zr1wr8Vtji+NAetyAyn4YvkekT7muXM49iTKxNf8v5dM985Ivt0iuK
V9TA6OYFpSFK0KIT+Mp041TjsWEPmM2EMK1Z+GvFx/04nBr/9AOhtVOPRJmfc2gX
JSeCj7yzMq54wtR1d84YdEK31qJHjfV4cvKFXo+IxI8pzRoHv9Be9K193qzLSpBt
CB0a+HX6F7PHeDyd/z0fsQ7VjeZxxKBqTq8waVHwLNr01iPmnDY478sQxzjALotX
LrfqP8Obqw0x85n1Xt3PkbA2OHr2HM4qSOnfGm6eTR1Ha8FTQOqtu1RvX3apb82b
oPgqZz+kqbt1UEAfk8HYpBFVZgSXyphy3MTDaHQSxXf3G3omkXwqWF8t2zLgt1l0
TM8eZ3+gLUmKzavBt+AtXxJj6RKMwqZocNDcAxsBvPBQGeJgo0MrmVjLWdxSHNQC
4Q5sPBQdizQqoPtc0tN8xeXBDeCgyjyJS+vNy9HiEGUwX6MXqWt+Uv110gjB3fO5
R5CU3K0gJAvpLXrd8mU3uY8PBHlf5U/1lZQWKo3pGiQg1tt+Hu2GqJ8oLIHgQF6r
Q3VUNA5PR52Ifsvh7ZVQ+vwaQgTOKuGsDj+r7Tb2S3W2AcFVZrnBj2sPzonDBrMV
x78EZpyyam1laTnm/L9zJ+TW21LATzUSJeEv3fo9+Ud9CXjO5L+vjTOLZy46hzXl
+Qoky8aaSIWz5d59ahEdQ52i4NPcL0g0WYFxVlm4rkMm8lQK6Quqp1SyV4Pp4TLC
k5LUINFqJwy0gGhhlHuLMxPo6ULeT3RWGJTXvt7Hb1tEIRXsX68GSHvMdKuwYTSv
lfusn64wuTu4NrR1HMorI2Pqg80DKlKvfa32wr59guhgo6cu75ZE9PZUTjdj6xsI
O21WCdvVwTHDfGQ2Q76X5GdVnbmHZJmA2zgl19gUuNt1HrRjx4+oD8SqpEN+9eQt
8rgi99PNlWKj4olfqj8QHBIJ49gGC44/IFKRO6gCZoWKfo06OWr4o3KybLVzakwN
6GexFrW8WIx1LyC07p+IXJec9K8pDEngnSXv5C1ieCjTXq6p9QpnCzR8tqR8Lwnt
uzJiFI+DNkkWpmgmYy1LxdBkOtHkO2vX0dbnTFwCTYPvlx6QqvOLoVwtYjehRMJC
+tW9+2PHoKOC/ksCtDhJ4G+KGJQQ2pflpXprHe9etpaC5wXcNGN8J/BhCaCwWXKt
UVnZ302wYmEhUp+ke3HiTRD9C87OZYM2N6DZf6tLHI8ZwiDOj5lukYShqXA4XpIz
Uq67BDPMxC4K/f+zWUsiYer9xL3DrceMQvgu0DLOkcXV/l2y7QaMMBTfEy83+BPR
vZ3sddKmgDWsc6LNQ1+N4sfdhGUr+TnrqLzn/XIlxgE98oZ5Dxo5YiRInHjUQb5m
TmuXj6b1sAWOoFX8VrKbFOGhQn3RQl0iYV8Gi5TOoFzuw9VPkwoDP4NBitW42R2Q
rOAj3SnT4JBo7cPukMA874l5eoDu5hFAqbioZFBdP+q6e4n5njT0ZxXvgdE3ADgX
M8RVTYPM6tcKEgimhT0D5FFwcrUBeWuHf0YdxZPozYJ0cksXalfkwqE2bGSXuntt
4rMh4X6i7wYO+VSQ4O+Oy4che278LyJqRdtQZyX24N7MWQ/XVkHiwsCWR8htt8yB
LLVepjHNuom2h/UoS8QOjhrXuabu0AtumPjvwTcSQyqDpm+Px6qVyBazuuwMutd6
TyGQWjmnxvV/2CVgPaAdNexKdnixgYOXq/GapOEZse2kkIdIV3HVHUIA31/qqdY/
akQYQ6LFmWdluzejHhLt6HWH208Fxp/W2bBOpitncdPAqYy+ZFfoTiYZbeAzSmam
shKCnOaR3pmbUvMRhAKouuvsugp/WMRIP5nVIGt9huOGZM9Xcm1CTeV5SbkDSBFo
U5DC6tfSXAERq6kicrLGK1vXBsf+Tqfk39KfmqWY9pGkvE0idl44OktMjzpJkreU
9SDGAQcezO0cXOTIDkFZtXYZyERVcF6A4RUiINVrEH4STprvhpzd3YiBjNezeKOZ
nmqppeeno0DQV3/XzRfOqYhWkc5SCpgh4FgqKmvTUMr9gjcV/utXh8uS2mXJLXrW
nYY2yDYEJ9QuMt4fqjQzAwLt/0WB5Rj1z45rfojaqNK2uD9uMigqBHMPVq908Kp8
7/u0SgGWmPpQuopQnf+i38zWQ696g7hvdjBvkCfpWLNK/Gcqap3LumZNqCrts884
6AjC+9CUUA0FscrFc6yK6Jdqmqz2senkBio4t+Pycs+lzZBpA61H/KCcYj6nO/bh
7mGcMUDNDsGYkaD8ZUnpBUht/lvD7CNXKOT94eP9r2po0Zz/+jt2YaNMkw1Vg7tt
YfWamusKPl8p/iDZar0vBKjkzM1vYWaS1MwXQm+ica9UFZ/kYS5lUoGs6jeVJ9oy
pq1jbTCvNimsNlkABE9p5Onl51WfGIeO62TifaiKqcq3ddNrT6khyIuW3WtA/qLC
aJepUosGt225RVNX4dEWu/zThNFvtR+64IrYHZc9gJOaqePxwehEocfoU0qwGZCr
/3uHCRSasRbc/NPrTd31GeFonp3PCH3intvtA70DQvNuYjsbuyCVIIywDBSzqKNG
kpJhEaG1rWGWuZPjYLBfsTEJStoUd+x9xCeaDrkdstB+Oj0Vx8GswhOPIyf4web/
sBT28RyQ2fdyZPqG4I/LN0kybQ5jESQFibs78utz95X4Vz9E3dYanTIxVC+sXMzF
qqebcOTOAnDuegYR0P3Xzqwt4DAm5Ydj3KCAloTnoOJwbdvtzi3HopNsJZqEZGMJ
3EhOqvc8V0sAR3a3IkIdnjC/QVrIU7JkwMB3v4O1ATOAB6dSkqd/HDhYgT8c8WMb
5NlHKuI6uQpw9S0uxfta6JrfqvmSOu5GouL7MIShrKSb+8JvmcagLuaBjqkDDrWC
DH9FTCd7bHhc4T8dl/jyrR/G4nbnbxondmlVLjVft3yEA/0m1TFUlNQBM/m92Jk/
P7t6jbScNJoY/x6Yxeit2cUnQpG0U4OYLkGqXOakONc9USvwtWoE17C+3QrkIocn
o5YDavlEmu6lAFXEvIrwjQmmqmq787NzjnbNFXxHzumE6q6wcs1XwFmi+o3q+ReP
IxHDRg8Wk/PV+l2SbKxk+s1WINscnHkpVJvM4qRJOPOd+ICjZYz0YVu1yIdk+z8G
0m7OcQLyBEU2qfqDK9av/PyEmhOHlll51iJEYP7G+ZT0CRTCJ7zpCRNwfQWaw+LZ
iCpJ0cGnfqpMhaDhIm+K6AIe0tdi9kivLRJgVcreROsNLaZdJ5pPhQR0GyT4nOPx
vDJUuqsncqOpOoBGf7vQ4KhKgMRvb8cUmLNiMe9vBQNgbolx0fm9xjPW6viBa+s6
P0bWnMMjmrBslKeTDCIWKXllwTySZmxwRAk0JlhIer8VW3dynpV68oYkRwA9AweS
6q7UKduR1ugFRhxw1JVJrVjxgv+fZ4mHxc2rU7c+RgsvDohHoxiVzr04fanyQpCW
2BK0d8n4ZfIBgW5herucNeuu7uh2iQsXI9CkhnSzQE0/31z73/jj3oQh9ghpfBhP
Ya6QNUQUU2kO0EJHfbTAsi5nXHGFZwh1j1qwRZcIOKA4eFX03G6qcmAzp0sfBQx/
EwR8mUELqo9xipqeLa309RB3/z6ZQo82hG6CULMHl7e23ci/n5aWN5c24KR5AM5u
3ad5DV9OAVAPVfhOI2qaLc+jBmWUNzczjcfv2Ro3Kuj3yzslJomWC6hL2ujn2qId
egKEL6FGvZttHRQG/ljDUIgBUTh2NveEkitmGXO/joX8c/ZZSWVwJ8TXgmYxihsw
rR70EvkDBQ94pdtMWdWCldLxF46CMnUPKBhrrKXQM6aVv2qu3WfU2yHxP7PUvAOm
XGqBg4gUcxvtu/FVTy6Pxbnp74+85cNF7Xauig/BkRS434BDfYLfPl+RWWAbgV39
5xSbfXGkAo3snX84xEsCzHCwjx5Kca4dH8YOGmt/7+EAgdqk4dyp/sOaV1r2SUwt
qRlWIGEGqUclOoJhIbCwyuCDccYam+yVJqXDNwAD3RqiR3KAjzjrwoFIppP6Yk2l
eZg3KOg5NV7GB9iRHuEky6V/P4AJ4BcmT6dqQD5o1IaAHvDSjp/uXMR3t0ZM/7+e
DZRcPpyHWl2NXW0z+h11xXNRy7jRcO8rCXfJ7PzzJqE4GFglaRxkSvdB6n4vo2w1
7pDX60fkN5RU/Bi4f9NSomQnA9gHEN6ZGQeqbzZw/dc2qgVHiw+baIuSvygfk5zt
HU6cPOao3VXN8l9jGf2Dne7tN8SECealMk2t/AuRI2z3XIo2csZ3+1Rs1DbyeHw/
QBq9h7a2PuUL/tnkbhvbzM8FtZqqzuhrzafHQAppx7J1KWDITlzTGmBNHY1OqJ3w
H/v/IjgJA1SVTPuid7Z5HOuDKl0dKyw0zT1o7Hda09coy6C5Rv4IsBGXNXIN9p6w
2Uw3np/HUxZZWYQSqqx5a2xAyoXLXCWm3pihV4bPZ1r2DvgYoc1lTZcRa+JQzfGB
IPzE4ir8ms1Pu3EkWkRbfE/XLJ5p3SDjj35zcvE4xhmqM6crbSz4D6IwFY2V7450
jRxS1cw02u2/0rHxCoDJG0JPPY+HNPD4HCmwzs0tslYBNW+YyrCediPLYm1w/P3Q
fFuQsBGy3k5qFWwKSWbviFYPgxaOXDCykjh90bSk5t95s1zfsHOEWLT0T4MAbe/j
9cAmkgscPXET+LG/YViGl8UvM/L/3ogtKNGdgyfWejeQPNPwMgIZPxvgX7EUsZwu
TawILQ5QtaUeEoy1S6pQ2nqfFR2/3sUJrYW/rDiIbeIQG4NG8Jg0q1KLbrgXxUX3
KZVVVf+1FQZqu1C6Yf6ZD8Wi1T7fuBacY5I+LfFGQ4LVSJ3Hk96SnMvBTzwWFJ08
G4U11ME7xaJEbJGbJVGU4MbXSo8GoE69Em2f1oCjzsCDDa3jTG6RtBFyYkZvB48Q
GoxTbc+nExzLKKG9cOlMMMShOHdtP3NcCA0/YgdPoJSGFlBIyClQBZ1WSkGaqfS1
5eIMRK0b3XndlG6ORXwF4Xlb5/t/oab6JIN4xosWIoX8Ptw6KDRo1/HZYI77v0oA
xCKIHByVxlBbtsgNA6a1TzmoeBvsslQ9OuW9dK9YURmIHEtwAMC1IwvOUbGt659A
bFcFapShQH0MpORp6gCRNwQOFN/nZZAhdSgOfheI1pm41ICQk2DwreFxLj4/D4Ow
b71A1+chp3JKk5N4gjKcm9ToK3FQDVDU67VQVFLCtdOqi3Uh85780T8NERsh2Go8
5JVIA9xHADp81EH+hCjlaPB99anxiIAAsgjXlSWEzgIsedHUwE/X/B/oCB2n731a
tFgLM5O7g8NDqVm6t3Agj3ZTs7N7hdC3LjUB8JHmvX1aE2iNIxyeYZ3jApfFXsvR
paBIpo5N7cCop9zHAf/Roj1tdV9cs6eSfrHmF/u6e6VskEajI+3MfJTmbTw6O2tB
Z3mFuQVjCawEAjL1M/VoSj7pqyJ3LKH93nUqHUf3Ly7cfTeMGoml/PA/m5Zh+NHE
XJqScxHOwoHPnDtw5E6R0s5z+AMGlPwux4vs2O939TOBk7hVoHzv7ZceghsHLNhG
ZVCOxfQxqMgVUvBbcRksTPT6EOyvdetxbkEhAk59PmBYafLX8V6KUZ5XkQrlPoqP
kF7RA5o+Bw3obvMs+MEBAtvumacHKvPHRX0JXeW5juLJRBU6McXQ43D+/9RfU0ef
hiTsnQEMPJHkxjppNI3eVoE8EzCp6PsJ2BX/aIuSebMPVxqjyzKB9/oLSVcquXeq
U097p781g3UkG4N6Gh8xymYgt9LTOe6Ymbzu4IrdeEsZKE2qd2C1VP3wSaMT045m
00p7vvDR/bjhMzwLNMzJEl3Q4PLudFK3qtLpDjOVEYmasgIkxbN0ZPTMDiS/cawW
RHNFFMuI6wsycwhPeCcGqcts/S1N0W9faHyyK3aHg2dnLhO5In6R6w76p+tSwq8v
m97i3rdR76EcouPrDcoBmtlPsaKcrVhRfKWY/aDXOD+/Ts3Z4rBl/YFYB0rVkEKs
eyuBKt9cOqXS4/wWddh7eL0GLKEGen9i86bZdKZkaVUgKAuVPYp6C8bkhFW4sYmM
N1Fl0QoQxbQdB2joHBoAlNPQzLsi3w/Rmj54cv652rsEvFfR8ZeEj7/67obnjj2t
iV5d2CAxNGdRXojpYnm9E4wijSwVnx3f4wRs3MvM9zPWXLTz8VD3hJOb7STp0ydY
BHPXeeR7RdU06ZyqQH80+aEVqvrlN7zq17ndevDOnNwEPXdUy6nu/cIU+1/zXWI+
HenBlRNSxlIhkhRsfkyGs7+QOrND6x7RMqMkHSbRPvDMPY8TIUBbgqjiFyDNjy+H
MQeb1rG0jNPnWpxf18xDHFbmKAuyP+ZwHYfUcGazwUzKWENtrWxq9CL/2lY5U9SA
gHxlT61zrcIwjD/wIXt/ELCsRbMtI6cTHHQ6AaEC6ZqZorYMWLVk8Km9MQvRNOMX
+T69ur268ZaIz20B8QW+lcPJf/5/LmjJXNovCy4w1ziGy/7HznOl2kqeu4ekkKUv
EITzBui3grPsErNV0PyILaPtxQB7ktnAdbL7WtS0T0lsaQkpST0F7IMUtt/pbH1e
FeM43V6nCOlLsOBNYxgU9oM+B9smTQfQpjJ1ZGtTk3GIxVYNdySLgA6M5GMZ/vzG
z43EcAtHQTPe0RwB0krhFseI6A2iPlt7bGCd2AuDBqLvtWq26eaoOk1TNyxdptlp
I/RynbXuvdvRyjxqSaDZv839NVmmimuPG7Zm4MBeRePkH4JqyS93n3W6pmOU1ZlC
69t+lVxbRorhR9PFs7W1CCDaUt+nNztjdVqiRFW29VHaLisZhI5giOQZAXvjqfUO
IEWDZguC1yxE87L1+PR7EpCGHioyx6kPLLsE5rgUPh+yWHxfVOPyRUtj45dM6odP
c+XdSSoYJyqvt78pbGl5V0EEYgVWvbRLFHVKtLHuf1IZJnNgxaQTDQcBbgfJ58Bm
ljZ3Rfc5a+6/Fe/yjYzCEzdTrjN6uz1BTgoxEKfkHuWF/tCixdOEJ4pCOIAe1BHQ
0IMzcaD+j8cVD3YIIbMI5i7IIoc/3lR1s8JHPOsrodP9qnS39so/f5tpKalz7F+j
YVp3p8OHtw6pZSt5GrWHwQmrTigJZbScBHE05ffboiLSEaadLAVeDLCy+kwvDfhk
l65bNrcQlmu7rNDWcb0H2KvRacBODGdppIsV12CA07gXGReUILZJ//XRDzvEI/+r
EtI2Rk4pyM0VOBOqrvns2ha7uZfTYJKA/+FAvmOkojBtgjfh7qsGkjqejqNhGFtB
ALqb133SWw2hNp8U23Qf0nE4dRZQ2leFDK0HRG+j10HYUb4dUBkJct0CH+VEPc7n
GnLfbTumEKyjjOBLeH6Jc9jCEqoLKEEam1fjofBDsuQGvYJMQok47lnlcGUU9sXc
+E6FfsjzjuXXOm3v/9GddfXjTtsC/uRclhF80Wu6XFncfe6zI1TgGjq146fwanuZ
A3v6QjHVCH/OOxZwE8ONYA8QOSt1obcl2PiMIvGXKgbTfRpTXflgrTj/wXwURG5b
Li04KezfimBnhxx2i3j6BqQQO8QEJhUD7hW/RSwb7DCh+hkZgLFZseOWvGc7k/wE
iDttgoyupcG0Nf9z/wuIwcCVSJoH25jwdju4hAE+PV1feyFFMkGVPgLKoRMCIFq8
cF2cq7sxioA1Tk/LeGbTOD/1Lvhq3G+WoiS0enB4CqW9QBcFjNwGjt/GveCPBet7
DXyfOIP6E/L/zwXmJ5H2OdN3x9p3zuyTsTUrUfW/RB4fnjpVakAjp/yFrGu5MmxV
Ofi4WXqw8ep2JK8jD+DsyLG1TTLwavwZnvLGAYFjG2z4TcLvJoYNFFAIGKdIOiYv
OdYaSUregzmDyoYBrDUv1jNbaifqWRwpPDMn5nveYgFXoVbb/Zwp03JO1GeVshIz
4OH42HdQM5dl19UwQrgTky8DPIB3lQ2n1S6NLyqhATYuWNlaZlIUfl+tRDsri/mg
YIC5Z1MVcWKGTVkoYeQQDhs8Ed3YSP01kSxgxGr0h5Tv5vfNHG3a0x4BjMt177f4
WTXUqS1PXCn/YUrjSSIu+0zSMfuPVCx62V6tHTkTpjGrAZSA51wE6cd9gcY7A9ZL
jKx4qM5TYfl/K54jtE0DeqiKhKcCTfcJtlklZuJXIzW3lunpqzz2qvWjKq4+67I0
L2s9HLMfEn5V0UJRyk+0NYdHqwHeYWWrrpQr38V3MkSSxaEKM6tqL2S4Rl37fKvC
Dbnh+uRxkrMckv5uc03fd8snUusQzFzWNQXbFvOim1IY6T3qQnTktlL+ouiNlrEZ
lNVdITCSnDHPi+0m/Awut2lkG8Z4sSe5VxCH+uKvy6V02iyqjncjZ44UPtc2K/hF
RvA+HQYEqr4aCfti6y7cTdKRdp9Jg/AleQwkk4pUSdgOLPrdIFhOmzbkAEOB1Hd6
WDnaIjF+F5y1dUtQq5itlgrg4MB0ogKAh0NqVAts915fVFGEb2NvTx23P9AM23JL
hAsc7goD94dHh8kPruRZHVhCK62bSD3tTifykyU/nRBk7ZBQER8ggoSmQw+JtR9f
WBi0WxtaoLeZTv6AvOujdGHJRCtKczdNetzqAv/icQ1pTCZrx7b6u2JjYTemUu8v
Z+Wu5EDs+rS3Du6S79P/Dj7tFgQhTJNDDjnNnkbhOUEZXw5UkDEevOnVHyfRM3e5
86RRv2YuB/U1JPaHpvwro39S3QWQiN+rNc1X3PflcyaDa86iDlqhq70ptkvicAeX
mBXGLXfFZLobjtk4o2yTwaTmLT4uOfsB045jEmHv8tIL+m1KnBtiR4TlB0w2BIts
HGx1nXcMlvIvlCk/jvtHqhVasy8flMI3/zeTUjbP7BVGX5TSCYPo/W9uUc5Y76iu
z80UlihDeDO0SmAIMG/u+LGYoU1Ys9vK9dFeRM7AZg1QLOhahjW0qCg4oJ6lEbhV
45RbK1Ssxdk1d4sscgV5t2uIJd4qCcX97SimwxuipPlQqbaIOkAc8Thwe9AdOUaS
79m5NgTQGRRF7TQek5fvioJc2T5LbMg6KKlPha1hdbX4leuy8jSvDkB1CnrMzCSn
JtdGFY7aEMwzocEsoRQCv5QJOUqUwTvDbz5/SmnYUGIWM4kbzUQ3UNQwhGL/xbAh
9VxlBczdEYH2Q+vb0FzySPs+YSYMotHXRKn6x4Op7IHJBxEwfcZudzbS1IMwTRbM
CtJliwcUQTSuQCkbYMj5AFEq0De2g8AoEZxs8LZSBZvTaK3YKD4W9WoyzBpBfVp3
0QwFa9R+GvLXoNYcdc9e4tKR/PxvpS62vqS6QaIIF2q/NYLKoii40hDZL+X5t65t
HyNYy4O4F9MNKlTi0Hja2Ps9iBGHXHLnJCC3Qb1cDK6byAGmrpzOBkEcL9JYmRfZ
iz41/ve6oMh92WSBoNZPQUWiqAnDrdgESh++hsie2Gew7qkLDy0vN1QXpJJ5NYby
OOKpIrBfyojhJgkNwYS2rnnEc8IbBLx9TdDnqvm0aXa/Fyn3x4OyuRrjGfbai84y
p7yOV6Oxnfrh0kPu2QB5qk1TaI5Qv9phKuTZhHW2b8KkPMj+kdueqd8pwvmmK9zU
BruK7H+S8zF/Faan9GUDxmIuR51kyX31RoU+ZISB6Rylpt+bReiZ3MK3j4EOiC/N
KaguXlB/AO4ZdbQ6Yq8x4smAM/6Fkxu4QLaCGIfreQRhk6bRTmFmAAXb+SjhCPNt
uKbtHm9/OY6xkbkHaF8GwydwYEf6S89MyJxpNPonvxJHrTkthTxkSKjcOJHZ9h4F
0az3fhMUCD3L4Ew87kc/rYkG39vIADDS7gu+Um6a3LutZxhH/MUSi/Pqp3WM7W/7
bFUub36S4YMlnSOoTOoInRX3RdqS1xfztAGEBNmVlF+gysho7E8ZhPmgQf7YdzGR
sjnQZ2VMDLUs5MqgikhFMHnht8h6F2NI50qIle0127AKEr0eEl9p9Bt0qOzZ3MVG
3tUugAFoM92OuoIF+44f8J1WCIqCZswuykRYmM8F16rShJ/6GPdwVpzqVgYe/ixh
VM8nJ/VdPXKD/Vk7Imcyv2EHErwWcjVVxm1tHkcc8A50ZxyCD61eUiuCPPEYuoLF
dmyZD+lQ3mPTXOgYH8QP3ncAr8ecLI/83WkTe8W9RKBYkTxOw0KUQdtIPULJhkW8
ZnS88Zj9GkA+JlLGTf4OX/gWVyWmgrc23GSFHFUQohL7VaeJmhIdSi63Kord2yUe
FqB5IboYJDnt+XakdeAsBdAR7nVVDerHlkgFYHFZJreu/IJsILFFW3hHqBLdEN6Z
sMZcHPp53WaNcOZV+mxDVcV5Y4eMzv5CQNjgPoh7lqE66+QN2krVTLe6DTTxBa0J
9op9D3BYARuQE9Svq4400bBm7C811/s0JhkczFLVh16a9PaU2bgARO36u5P+MFta
J5yl3D6juJ57lnh9Nt4pJvYVrKhzb+xnmzjU1sIb8IzYzczXge+Mc4647pdytvxG
gBQjT5lgvRv42i33miFhlcfifGtwrISbMuQE/zyE6DQq0Vm/cOLQiNqlbKWn5FEU
6TNo5395g2VJS98pae+24X7Qy/pqhOhS7uHP9eN5MAQ9/JSJ4F3+dBuQFmUMTWwg
kGmcEx9hS+PXdCWSHXbxczzwJnfNW9KPDkXbZA17Oi2J5TnfIFGiamYWcFyu0dx7
6VS6v6p9dYqqvb9j1T8Mn6MGnhFiJ7NVj77I25PfCoOrw/giUc2wGiMoFIvQJLc6
otlg2f8K7A12FWQLP2CXalkAFIiIuWZP8eC4jqdgb/iNbQV+xLg074Wzlw3UB26n
6xR8g2neD7YGjyKiJhACQDedraQxyzbw3xGnwgw7pV3UBRP34LRYhy6y+jnlaCRX
tJsMHCDIkYGTj9J9i3x/mo7F6xPjMouS+WPj3G5Wg3lrH+rGFJ61nQU3xjRx9Hw6
m+xzUA5tYPjq0SYSnTRPswdZxrYIJ/eIz2No+fhzOU0IgR+K3t4dIBqWUJpN88Cm
4wO/fClwJeVx3RJhfDF0dx3brkIB16aUvUMNZgs5sZS4znJKxKwkbC488OgypK6m
9SFWiwAWJtxMlUphcXgBZw0h71rCDzhPlFrzVU2v1OQie5bdTAr357wQ7RQ99aSy
Ccyax66T65mrJbMQaBA/f9rqschEgvz1QQfgUk+O5bpdxzlN8a7va/ZPMopOLkqr
8QGdw8ZHbKTIru2u3KEpIuqGfCNsie63AB7gEwL3dspUgwKV5VWNuOsPVWQV3+bQ
mZfYc4IBwzG+CrxJMdJ0+4eAODM9GiOZo/uMDKPQs1ftzTs5y9z2R/hOiGOyxlt5
ZgGQnsnsTjIY7accrkMPLMDwjMif8W7VJI5nR+XHw3pbqqDlpe+GOSW0hfNN7GJC
ay6WpGDRJjgMLJ5HIN2/mxmKUKBVVY9IY4B/NDCEexbhDgrRZuTTHMhGpd7B73YH
qs5HzxKtNCYXurKtREB/wj3c2WxB0P3to5pXvSmoPP8/m3zJh7DjMsEaZWRYossK
Brh7mGtAMVRqPSOKGaOE8YrOiUi2ks3WOjz0VfHuM/OvR5KsSeJgQDoBpeOrBExD
QOdkQDvK/9jTEKrNmr7+BDA9+6brYTyAY5VK4iXNxtaZ8IBqMN78PAFqaZPFnkIy
cKseX3Wl9VXajKyYBTG88oVEF4+jMg2glHZLLKLFaMyefbqFZRhFMNNtA7YjPNG2
Qzg4gRuYHPx4/StN4QLLG6fRhw6/goKokfJ9uXeX97DhlTTO3jUSfPvx2KVAOOBB
Yug5BPS+baruGENcViNlD66P+zA6KarbPUgFYfEFyCn6z7Tb2NjsS9CDeDB6YOY4
QFFsnaS+jHlwttP42wKPgKAJN7wnKSSVSQ0100ngO4BvZLlH5EEIerize3gCZ6UE
8CJi9rsFIZ/z0X021Sknv7VRCBJTYxs6XV4UY04aRa83IUXSBUsKwafG42V1bRtj
r6lAnV7wz0mpusJ+dqKaxPyGWDEiZOPqvXN2bsChJ6M9g6ftI0zE/b8StEtDJJeX
qK0M9D/kDccWYR8XrtNIIpdnL9VH6kdBWDo7mtpHU8iv8bFmOjlRkeSoke6Q6Vlr
DN0InZPivphu2tfHRBeCKlTcuAXWJR58gyaB+nyozJTnd/F3Y94uFy7Oi9/rseg0
8ak6a4fVI09vs1bFWbdY4+VDMWRCCZ+3J2lBo3dPORqQGHzRuqJjQjiKn7UycYLK
JTzMGW0EBz04/FZdpDD3rKuR9yXJ3X4fz2JqwwoOAoH40VXqfmKqE9MPt+A6zucm
SC2ea7MlhWME9hakGso0LL65LTSGtZEEvC7AU0EdQos4osWC65FavD+TZNPkZTbH
xrokcIMIWrxDhxIT8tSK5/RnDEwm2jZqyu59bniuszNcjmIFss99b0O71wuW6+5d
cqzgtXrj6uZ2J9oy5WkMFZV6HAbKDYFcwAC6NUxPSi4lXjQXx/ZZnSTwRw/qDaFq
bbmwvLu05X1W5Hus1hWRZRtdUcKy9bpJOVbYQJBsj4NL4TqwvRisMJ4H+iUhkngK
mesRYzmm+1/+YDp1NUK5h9mBE/4lSVSVjeEPilWE6/HT4CEEUKY9eq5OwKHpL+BE
23AsL1SuNfsvdhHjhXc/CT5QEJ37k6d+6IdCYhfA/6WZvKYjddrMvUPuDgiYGXH/
JgvW+8oK9oHF+YIHgekqY1UzokIRFvFrXOfCDabuEx+w45QSpN2nxKj1QIzVJNn+
sPGkR4zj5kYSjvyLQeGeR6CuFDuPiSYLg8KcalrPx7my7mgbksl78yrUdGPwiuZL
PJpmrH9B+wMcDPQAO+g7CqxyAtZikf9A7Wa8aSKKXlqkzahq+dpy+VV2HDM9Kgsn
RpqwNrAlMZ6+2RqeeNoeLk2LiRe4wZxbe4nu5YjaM4LAf1xGDWXcYiOOT4vm7GuF
d1AvkCdHcDwX1YOk1wN5j081RHkVaBxIY9zKCVlSvuxbFen9x76pV2kmOvADOC87
JYwWy223gtfCl1/Ll8naLGg5KAAyw4iJusf8QBiu3aiprzqF10z6bxZTp8ZzCz6o
twbk6XwiLlbYsF35eN619TnjUitfK5a8+iORQLkYCFxtNSw8KQvIg+kCSN8J/7Gd
081Ep1WseTAp6XqSjmK1WgMbvCZzfQUc9VSxgrgtcZqTaeccqFU0Q1Rht6hWo1Dt
gKVaKwmyDXmzYAU6EzKU47y/g4tkjr5YwsS8eeBik/nB/GMRSaXDtXL8sf09w1Af
NvfKc4teEofVxpKdvl3eEEUXL3aJLUr8dh1JiIBsKW4WFIS3Bd9kmdZ7fW6CjnJ1
xzxfAr4b6OUKRvGkhfm+5XTWVQMui6uMuB0WzO+17Pi9QQadD+wdmasAwPc+AiYY
5EBgbGluMc0Xxqea1fcoFsmFSB13XRzCT+3TsUbqpXEWYcYeddih2Daxbnuo9h/B
4+GX8pJwiejWK9JLieiLLtQ7Xzo+9QNUElMZLR/DuMZJV5l72YhL3R4PnkzWhJDP
iHlVyPNU2oQ19Kl7ju6+3PKoCPIBlvxHOf4rkMorXR/6ouIBZaFt0eHNwHIt8MAa
9RtQJYMkG0Bm6UskyQLcATmgaeLIj5iel7mEtsiMhSEFxoDxICPHxo5DB4tV8cPD
Ok9BQdFf6Yu5WAP/qS/tGdfcu+Ad655gN3nbjIyfqfwfezNvoK7FghNSBsBpfNL6
zB0fRRPbyU9A5pPhsUxha12oB6ZzZOdLesy/aE31qiX2Bzqb1/bjBbjcffp0TDL6
BkiWn03WeDAUaenvdw3XIvrqkyjIsUzh74cWycrnp3eH9iTpr40xOSF3I6SIJRzZ
NuU+q2g5CY2C9x84pej9ICzuvSfDKWWyfLoLwi+Cad/CcMErOhmVlINWTHJembys
7fL0JJag6dxURBd3/HgN80D70f8Dnsm812SthYtIGgaovL7gP2J+l3HZ9VznGNTy
CCxLUmXPQp9zvVXVCzPum/ctC+DiqhoqV5WKycfjj9ha2B51i4+39oXTK0PPmN64
AWGB4xcxTV3PXzHGUfNkjxWhU8ImyRBeAmI62OxY6a//H4dIeJru3IIYWRT5kOQy
6qd01P95izJ6FK1YyGl8j40ULfBxjwo9UVi27ezuW5vjFkLkgYtH+VYyu8jTszKz
vHhegIrttVuAtkMT/1cjytX0RbiG4uXQm80mrPIgeM1cyIA2hP6TXWEExhaGN6T3
abFEAEXw2A3tzC6A3cpWW2dTu7wq4zaCvmuTGwuCbH2LPfbcM75Ob5puX1Q76Br4
O1HbLAgLlibvRTk9Z+ZYuxLCYz/7wTx0d3kFyCX6L6AayCAD+1rQHqmXYg1T5G4p
8rMBtWwPiRQFerokpb+v5gX2TKKHPoQhXVwqgr8n7up1fQPTw8IJQLkw4Olvtyh1
37CBGpU85o9srtWlAn4QcWnssTmfXvNb+6C2NyBiIm70i/QCpflFl+ts6OU5Jj0D
Cm9P4ggp2ovj1xF3OHP7cGtuXK1+bt7P5hRr3E32ZvZdmFDI3Y0YknpgISY6s5mC
YsOxyDQzU7mJcW69yDQkvqV5gLWiypEiypJIaMvQNnJt2WvDIVLnLF5Y2QZEzVEM
AgpemWH0MsAfrcj5/R2xv9jSFolvK90Ij09ZQN0503n182vlFu1zIBppDibno5c5
o5chhG+BLxb7InvE8oD2mNg3a2DFiX4qtMdPEaALr0HqJGicGnHM0JPmo/rk7Bzw
Hh6zZnoy/q6O1mg2zTUdegmLjry4IPJjEIH9/DNLrENcZaMS+FZcyqiJSiFRhl80
ULhd+1VfxhwPyQ8dVLHRfNB9CWl0ZNmm4FE0AxERIFME6fcTW+bpb9byI/gXPWQN
EgrE9SnrNxcfqKIU5n5wr4W5reyZN3yscb+4mNw1tsux6sy4Wzgp5P7hIt0paueW
HlTshenaCYbOqk9qwPBzGhBurOFXWgcmJHJDPMN8MsbK7t36g6Wb99cYdGLkF7ck
04GgZoVptVwtbNUPdkl43STqW/t5PDrBZyvQsKp3/a2obwkvwoGopVaObM+FR5Vx
01+WedF+JmwsExNmyXOKP9OffATKlxdhHNw3U9unsW/xUIewT3sLmljLjqqVpIMe
sanaBqCWNcElkBsXnIsN62DRxxLoJNcuwwJfFSuTCzjV3nV6E6mQ+9R/wd2A1kUY
HuVOy9GnsxigZCu6qySEpD1YHnFsqjfidTfHUsg9W2Ckd4g+y+D3IoXgvjdNPTLT
x72IUBD7ZYCG/WL/0HfSMGS3WIUEhDtzrIIpixYF6URGhtrpJo7q9O5nPPDntlDk
hvHVNqgXsgxcJ2A5+6VztI9ji//SZ3F+KWE/wCFn9ujeHo4zZt6VaLwR4XQpvdra
iV+VKs8HQnb7wBdpew12MoHjFvA89DcTrW8cdK1Ne7xrG7/h/ia3f96P7YTibwTu
QAlrZVrB531xq8LA38t95CfRE3IzR1RKZss+AUnMZtsuCqadvqIyxyVuImu/JgeR
fDaZT4acNq/hQpiQ2SuhCQ9svAnOsN2p9SHfqBOgiXIvWPtZWdmbqUWktL27IQfX
SM0JyhFPDxmi1zUW741M36UiaA6ky/L/0uJ3vN5BpSdhGSeFqr4QzsgSIlfm6hcb
Hg1Mi4lIP+dnSW+6qNZlIuNO9rK6x/EAvHrjzxRo7+24N26h2jyS1kMhZxd81wWG
Uta3vZtKDGi3oUkGw5b2el0WCGACjBwDy28mcPqY73j0eiKJGzFBcy1NPvH9UnBY
5621sN6efyd5eGGWFHu+8vfwNiU9lCczsYPdU0Pf2zvW35ERMA/xzb3UacmvwkiU
uERars9hFpACWViHelIOzgvfKdSFe4bM/Y+6A87C5MCrETwp6oDQ9Ao232IV+L4o
rbHL/iVsA9cNi86iC6EnEd/TzvrzxBq95h8pPIE6PZIjfKbnrMCjjPSYjlGNZi2y
vWWHwf6BImzeKQIcPkPRTPx6COfhY7bpi2nbz9ur9BFeNhWug+ESQN1/QeSG1h04
r0RBzqNE2oIBBQBtpQEvSghQ/vHkEKUG+TTomKz3T0FUESq8R/R9vA9a6ge4+ArL
S/UzOTz8kUIa3VWvE9tZaj4tWymSH22ANZXkVxpjWiMLYZqzQWM6zDcPhnZcPjb+
RD7aAGJBMI5/y+vkvHhQgbHd2U2QldcKH7IsJdOt7oOqQM7RuboEi7BUdelhGsz1
jYqaSqBd7FICISXzDVmrUnEmjx9HIpQ7EU+ySxR3PWfbAb8g6AeWYSW7YFXJvUjm
oJtBl0KiKC1lpPQTCl9c+7Uw+ac+mZ1nhnnIMp3n44V+Jpwtu4RxiF3+wgTJDMGL
E5+l9ZDonvJG1XlvyhYpxLWZb4T1PT1x8ZCiGdbibNDdtLLsJzkiNzZxRUTmhOOz
hZolAOIXiGryNg7g3LYp5Nslo9pe8S7f9UjaakAk/uvkOWODU4PFsehnHxcN8Uxg
t81XUooTh7i2CyqwN25M0KPUUNOWW6B+Nqh1UFzW2EMZrZu+CDNDOgGTutoe+bS5
B2u7aFUYi88MUS/l6mdA4IXbJk2wDIYYeGlZU6YJ4Zf/5orDb9m4jp+lgC+7tQpd
txrt9nmumLYZUeC+GUgSs6uDpLFUJiq9o1sFoB2WsGyv55ImKm+er9lVjuWE+UCw
4sAE4YrU79fyhJU0XeohTDpsQdFsYsfuzwh5HTLUXT0nCDont5XIrSQminu7NZuu
iHnxILLQSJsFi6UGnUfGN1Jd7ukz+tv00LqONkt5rVMSbRepWY8T6tXxDMyAtFb6
lTxPiLpMjZM2uRaiYaXcvsuL81/6UdlEtRELRyE2rqLJ39oASmJNBJdA+BeTK93h
B2tY8F2EOqt7v+thW0Rs3eNlZwejSalF1VX/ODhZfMxFgEDbbSaXzAT+v9XVboS6
QMtN7cmfGeAUg9jkqgNwV0icouLFc/KiRupL/OVngXm9NlYRC0Ib/LYusZfbnEFQ
CFt3szblfYw6mdC2PuA5MY6jzG4WJ66ST+yogS1roLptMHhAL45kAtyxG0oU0Cre
94O2Y7fcoJx8pnRuyDiqr2etjDWn4sCz+Q3UmoQQTmeFkxyPvgjK/4YoYaexwwb7
jgdc7AEcJt+MAEeVSTaU9MAzjvgRqPS+WSnf4IaFQIslD23HRlw9LnXWDD1w8oxj
sbB5n+kWdd78c+WsOsgFdNQWyY1eVaxak++2Ax9IguBLx7Bnv8bG2WQ+1TQ0VGA4
mA5F7hil6DNpFiQbCPIB+p5rEnKP3Nl3mX0hefJy0iT7u/CmvCkNPxi3dzVd6BNo
7i0KQhRDUIbJCnSfZGFjdKvO8xwNTLe7WIG/9zyQcIHNk50rXLlJNFK55dPxltQH
O6FTLromOBl3+k9aOhgRM/P/hEeLpmboR7VsvkN6tmN5dBwDICPwhDQ5c+46x9q7
DXJ7q5DsBCyn+TFttILHErCxwJ7/D145xESxctECF4qlEjJ+fJ3MXfkqyOvw0fJ7
61XgQwm8r3R+aXvCvGhpZxCTdexSArfq5one3xglGyQDuD6HBruwjTl5GEEGpfux
jKyn+7jaruq4RSyW2VuMG+B68FIusPI+ZqLG+AMMtMzmQ2mhhDS7sxH1xW3zCJ6A
DGR97zh5K0zuPZskpo1N/AMhCkW4tCKrqJwxw2Qu0gd/cd5qlioxqrRA+ckPBENQ
uFlcwRtEfdmQSvGA0qaw9ZitE880sBMCAm8TJZ41A469cr32bWnOGk7XPkSDIcTZ
F+3QG9bG4QbMV39B1shSJtaU776Pmom3S8m8IZraBVAnYgmlF1Fbeps3W3PvYUTU
AtYV6IOwEx2Df/rEawbmda2aABeEKmknrOKzGns8REwmFvoJGEyXjAkEPJT9AtDu
FhrKkJTVEbWBNTnVlk78Aiy6HbcVgcnByNg5ox4uopy/eqDQGYJ1i3EUaiEAZmXV
J2Az4jMSb+gvs7KBKOBAhSiNoWlTm69MYCIV3cIO0zCO7osp4fBbMzDRG1gS9nZk
2GOXy/EXcRHQvIPm8cQd3jMnYieyvbDjBNedjlBZDujAmktgkU2Paw7CLbHhvUmh
LZSJiadYk/N/9plpN8DegCQPsztX9V3qNX0Vl463UDIASMNN/kIgTFIub19zRwxY
6xtB0O5AkaHTK4bpAOyZXNqhlBU4iHeSq1w1hjpCS5empV9pG6XHkxVp8PV1LJRI
Sg3wjQftexh24Wgwn8uPqgQKwVMREhJWPg8fvxJafyFrSstDWrhAsgaCyI3g+ESK
35gTMMY7S0l+FxxDHfCBmM6XyFTC4rhYLudvGa5QT32CKlQRnlSThaNo+tDkGxON
FGm61u5n/PDP42KoVVPANpJ0hlYCNPMZ4XpTucYiKDG0PzH7l9qaLRL7yXBYyozR
DjEiycxryD5YvoKEIoIAdwyYSYyqlVLu1+ov9YdFWShr/ZGG/hVeXIRjEVfXxCnQ
wrlZUizyEqV7Td7+qw+1Cvig/qVzRTVRZSJuD6D2E7iaLECBT1RWX8cFsZIEldDO
2xD2kMXGYtyGcKJ9XFAJHdJL2hxIDULQxZSQx+ENpEl0WnFkHON8Ck08l1SvQ8U9
V4MLJuRXZVfCm/yrXcyj26ltO7IfAA9plm0R+Hrxwqd+HPrf5sMJie+mXyDZngJu
yknFCe9FAbc5i06woKnuhmJK8q6XEWjRBccv03fa+KE3szaMFrraysq3r3cvjSrA
Pn6EEXv18D9eZ4Jj27RXDcKIpThAM3dVhCb5JkMoZcuH9ECzcawypoWc6i/bM+WQ
5pucBgzUleyBYV2aFvCuqKLK2x/o5ox5OXFKQeT8Lvg4lzHdIGefLS6MSHJCcM/6
qDE+Z6yCRyR+Ev1JIykBoqWFyUZ+/izNtKz6soL1m4Up8T+H61mgdLNzeb1eHTAQ
kL7UAifFvUfkt4Vobw5ZH0DL80bKW7Ri40WKzEt8riEGqlwBvSfDhRJid5aIN+B5
pDC6vzZDVmyO1OSWiQ2nGGkbrbuhq4N5QEQ0fpA9cV/wnQrlx0q2OZZxyDRv7yDU
XWC+SH+GErTu/vkvBv73RoHMtPpbWUfwDWSjSfbbzdhGFidFXN8D29FcKpFOS4iL
f7gY50xjAQypghDj7CWp1gPy2QhkB3puNFTIad19EP5nsMAKLDkQ0zDae4YcQZye
rgScQYYCnJRdsaxqrAhY0NOi/wgaSoX+GBP6oD/8k9Bssup3gZUrR0Dz7yPaL7U0
QbO/L//mG3Ww1EE/8eDoZLSUq7g8wL7bAbZhk2Rm+mERnHrwGADoaRpIGshvVOmX
daVbHJQodeCdZCiawjqgGm5oqJCOKcTAVyIRG7/ITA4D990PrHikZrdtkd8e7C0W
+p7Nq+BGWuhayPOQ075a+Gvc/njx1R1LfaG9ODMfhQTcW/HN6WU/Y1UKIEH1FSJa
elKft6U7gcmxDOaWcHC9nebOKTTiTqs+GF5Z3+6byl8EEabdWvWrtlq7o1tXL6ik
Yytg2yqvl+CD7nfbnZ7PjxHCtMRSXfXQALDwP7CZdtkdL3mNIjrumCpR97X3Qo/g
ZtHa3BgvtxHmwJNTHTJY+i06YsRq9wgJpuaQ6zFw3wS069qsyVW49whcZG//pkTY
FinQKPt6cZ0fcEsPzsbT72P3YrU4+mQUQwnTRpFBYz0JNKLdm4Q7PA9pHhUnJvn3
RJydqwqSyVeQ31ql1oiqyhdY+1t0FjgAPsfzy/STV/BRPMjVsrv65g+SNCqz9Wd1
1CZQwIvfDbZ085nBH+TqVBn9Pnk9rX80iDatDEQ1AsjC2QrcLXQmglu3CiosCKKu
Tvkle++qdtnCDyKZJylIiCv28sJFXNzxDyWEPsdz9AOLiYpx+3PDQ2DHqZKYhLJP
gqGMzI6y4O3/OXuWY6z6BVU5+Bdd9h/jR5IlVa+d8xVW2ExGGK2FnFihpBSVFznr
Y8qtAWCVZoAx570ezhIDslY92FUo7Fbqif6ub1XPsq8RNTja7XwwBKByCNpBG2LI
KKQgsrAvTDb6OHfki6fotwlSgs/aFC90+C604eOSglfSsGoliGKUgBogdSDREedj
VgQXlf5y1tfakq/DmBTeqj0K39M/UcNxmQSvNMXNdCXtfY91BlSgjd9o4JwNdvPb
omg7O24RSpQNFfkw4ilogNQCefjCnLRhiGRawRXZpDGw3trKmwfx8n4RkAhhP13U
LLXenCM6TI0nkAHxKaUm2Bu3gbwJvDPLM+TRb0u3of3xZ3HH/5NEoqtZ7TK1J4Gg
WDTLF2wqEcNh0VYtDpzsLYItudp35tRZS4QjtFpyD85W6CNkNXErolm8KkvNfF9N
C3EebxxjVef+k1uExpLCYqSLsUNCjB1impIxONiEJuSqS15VymcgPLUvgWCADJwW
dm1RBNXcQVUC8+h5UFHIgukRDGQYtg2Xf7L2Fxcg8YSDwAr8gdWKFDNujFYOW4dj
rKHuCaMoLNZt2TLsDbnISkoEUxlJLqKsiWjI7V2gpoSZnp8V3zODlIBEPWVWZMLi
hLaeckab2hP14Zbef0lYx02itxyzcQg3MvcZWzC2v5k8TftQliJ4eXrn9Vu5mQ/p
cJjE3hq6cIopmPQsKBjrphQTwSQ4IjPP7K5O8ToVvcXxfpWOiZSV3DgC/OQSJcbC
Mdc8TrP0fqkSvnC5A57xp7nC8pA6JyrbvBEVA6h/vewLLTLX7SEXoItIiqRaz8oR
btk//uQOD2ccri2rb2OtWRPr/QFKigEHylvEK1Ry8bsuE8BeyA8bi7AkxHmXm8f7
+EHivNoiMEkmMURFQeiBdG6DkNOpD9YBe5PGqNiVHpTcwxDklBcgApvy+pAM+TYi
DaqDacfDlxjblTYRSq6J6M1L8GMXo/UimaNJ/8XHG24tjRGKvDy0INm30NMwBEVL
zCJ7vdkqD0xDSBeD5kireEnjVhkxktV7niOOTzjwI1hQch4nReXRIYB/k+P7XOgg
vJiV8dE88Wls+T5DheCy4EUX/3wKGS/mPeUgr0KXpo3JSYrLrBOYp7URS/Tz1OrT
qLjBSzro7Q4NtEkJez1+cv/xAVi5xNNN0Ho7tzvONX5FEui7RWLvOnjA6exWWLjo
N6a/q3LzkWQ/7mwgZfUOcccSNrJTNtFtgMjeoLV8c2JeA3Q+CPO1bDJ1HKVxvnHI
rqxrJGVpEK6TdVZuMRGju6gqAYrna/1fu1sJviPcO095g23UPqxx3BaSWv1PCbt7
B/8kdZHcx3tuwiU+Rhanby5m75W2bC1N4fGHjudD535GaJCG1hPx4MAoox5Kytt3
oWtrUpNyqYWHQfYF6MiE5Y48C0kV5Ie3iGW6Jc4EDhAHbkWg7Bo9jQ0XCqdAI/Eo
sWaSLN+gEG10e8N72rpd3CzZAyYnx2tBq5LrWrgacogA/pnYj/QXDukMfRrRzRMc
mc2DlPNXPRLzmdfyfzJWAdFyfsjwzOs6HJMUeiZsDD/woPpXKiPMphN8pLDGT2zc
44K9PG60eYS5JxvaRsmnM5UCDWOAtz9T+kDk+7N34e0IzfdHOgwQRN391QY+Dbjm
TTHom9QKEUvJhBHcW+pcd9XKtvihWdkMxH6tcPs6qnSzRHHRC4QW9RfUcrim//SJ
WmclZ7m4Ba1YEeoutA0PNRgg095ojB/goSksM7I0Gu29ywFXlGjrPJpwQo95f9H5
7wvkyaHzVoE0aQ6VTzJltYIVed/Xpwk7AsfnPRM+8EJm7I9nWitgsYT97Uxs01m1
sPK4mWze2iQJIvzfWGrK4feIo8O8miHJ3Yk6Er9M8x5ui1xkuSFMTGp/S6Rkls/0
w7PISlvoy0LlYcmDP7ZzgNShmkxnsCh95bnBa/gLD+uJ67q1E0IQVprJNnr6D5lG
OVNBU6VCNUymRxM0wp/aVl6erImAlAUjV5icOQNjqBn4LUqL74zRjcBF5O5KzfxD
4RzVPI1MFsyHwJjh49+Hffc0aBySwvjpyuE0MgS1yTbQKXNA0SDF/Yi9+Xkmr9e0
QuWdPZ8mmpsGS1CBvOeD91BYTOKpQ3vvtvvBfOiFlPjv7RyK90EK7AFGq3ZY3Qfo
9D6SkkS1+tPwq7I7tGuJeFRpo/FOP/FifKubIdnDW5aSMWkolNehiLw20w6RBIXZ
GRQo6wEQIVbRk4QUJYLLQIeyIgQUPPlCg7m9pX+fTxF84RAgc2YA8GHt28T/YtvQ
8/rpz1GJ+99kzF7CV6E6c04nZk2Y+y/6j01xujPZCC9f1BKdzbtbz7KP3i5cCm+6
FIKd2kZhWlmsllpjFPy94k5G8OEZFuZV2G86+Iu+gfNOvsSbOlPEi99R5AxXKp+Z
feIU40p9qZ+qRr+uUUR4xQdSLIcz2UQLvUDL7VVfFTEBNMepO0rMnnPFWx5LdA11
vus5G0u2DhfvpDxCZD71WRjYFv+CjowuCLRhmkVWSONiUd5EIQW70N4MChhFcPQ/
6fwfAZ05wua7QgIGaY4bhQnu3mD/QROaqBMnvrqJ+EaF/HC50Rv2S8cTljwIlCzg
Far+c33FslG4oNaOXyo8wzlID2hD5Sp+vq5uLjqara268xFvc36kY6OzckG3hMCy
WOiMaeaJVZUWIiIxMg3gP5jEyEXLgzaYM5RwJF1GJQCDZQmX1rYWbEjG0b84qEDM
mip0Cwh0Rg4dSpZDHm0gD5ivLl7XTEZ7K78s/LDqdR828etGLvojfpfelT2sInY6
uvCD2quRRH2xk60AvIKgCrKeWTXReYE73KaouQ9xXW0bvJWSlQD6RZEpNeUhHgDe
rjznsZvaZ2z8jK5PKr3lQebkKnvSpzZokKY/VxQvE2dDGUisW3x0dUKWHj9uoRgo
1fy3fpPgDgn+BV5oVzXi4vQkoXeVn13IeJG8SCPG1/FAm8a0lBlb/40EdME8yw7j
Hrn0mvTOzVIXGN5lOLrPy95dwN1PD5lvgLwko/WbxeZeIhVPE4oaI5HKQPnjj6gz
TsM51+m+sXsLGyuYl4YA1c9tM+H3HekXt8lBg3iEOFEb4iXjpzfuSpPAZzrlSZe9
IlaaVBV8d07+rukyWJxXzqfgH9Pml0ZXSfW54f3rLIXUDZ9bv8CNJbh3RtbFbbNx
CeT+pz+i34AE7+MxHmoBKj02NBFuGdcJVTolzo5RjgRknvLjz8cbghW+RQ54213O
PYby5sT5++wNYSVqsLBA1eZtCewVlWY/LxZXkibl3HC6hk8gGepp39EghF1j4lN5
iH0fHYHqXSE4N6REyAL8G9GpEejnGGh1UrxwmqAAQGGTAdMIV3KdExJBKzBwD/ke
7ja88Bx8pCKj2tHphMRBCXUElVRarzJkWJOFd8FIl0eeYj2wb9NfKjeBaUAPYSJ1
n/a3aiT8um9GDeigvL0c932Idlb5Esk8qJBG2fp4L91k3HmI9vyLxVO8Et8Z3Ziq
1J+Ye4OVhTSxQSx0Muv0dz3AsgvidPbCXsHsBxZp4HUXjzXQf6L21thF7asC/GE+
6KWG4Q06V1CTtlNCGKmdkSd3LooEgSkhJEP9pbmJGz/4zzSoOO+HYyxeovcf3/9U
YmJojGCrZbq2VPJyZRhBySH4/zW6pGE7AbsJbHkXiPiMIxV+ib6OM/sFBfON/MXQ
mbdr6yAtuapVQ6hDLHun8DvSYF7ExBBlLjTigwHBeLJRjTe3li6rJiyRvziJeIiu
0Ygpn5/Kbns6v2DE6HpEUF8SN4hLmpXs3kQIQ4oyDcIvGkV5mnsrhuNgHJ6kVMkU
qclfR5J1ISgBeem5HKz27Zg2cRoN5Fq31WiOScEkqodHECpBRv3Kb4ZrVO1iNUVP
5rd6JJ1bQyV4l2+h1ft42wUTanQ5zcJ2UhzZ4wkK8H0Rq3lzwFoiiVlRm2qVxzEp
of2rac9nsRN3Ql7bJKPe2Ff2AvrEe5MtIAzWcdhvgLC2y8EPsjdlnREOQuoxdAx9
Q9TymRWb7w1YtiRZ3eHTkPpNFjNH6I3fYe0mjOA9E2CxXIOxaLI3li7Wcle6kt5m
9W/uorgiMfq6a6El28wWkO703wwF6sKnAI6VCfBnc0RxXI4wai7lZob02sMsx2eS
/D+0Bf3McHaHE4oNP0YxPVUuPF1NYSkMlZIJX/snpeee37dGUOZZ1M8HjndWGupS
NCp9LroGciFUyl8joPQxQX+Ie7tj+9iEXgpPz+qbhusja9tOFw39xX3izlUmtO1X
iaGJN1wuBVRAL8QaCi8whYbHehpbCLV/IiaXaYiSgFoDb8j9+8XiKesq/9gQRpL3
o9dNH/0YoYP6ASqGy84uknj3Mp6Zu847Jispi0gQDwYo3VkzoPRjbXgs+zCwLTvq
TpWCHDTEvfRg25Yl6IPtVs6Qj7W6M+/xceG79k2cZkiFAGmkKEyYyBAL4WkXs1AI
J0GnCa91Sq2CBRJEXcLTwtUzAaagq7r/kDKHmjLn6YopU7TeDC/whVKDmxvn8wdD
rT9s+VeMHU17xgfqPfud4SFQvoUarXQwrovmHyrX6atf4SxIONMJFuUKGX/qJYym
fEsrfjQeaJMtjka/2/MV0X1zFcO7Yzmjk72yZX2lIGy2srEV3RBtBRXfILb0HUPl
S1ePZWhiN2cdQYyk27eHNT1fP6t+ro3we63ycpo34KP//GFAPKffyawmB/l0rL0S
1pWr9fhdU+m0D4S6GQt3RmCZViwJ3k3VoRJRoZ5VMvKOsKGiGDtdod0gP7AKG4mD
eL6jrNj8Hwjanp6Yi9stlGb89DhM/LToP9VBLJpm6cDOEAQFJ8qb60MndujSs7Yb
WM4s7V4Mo/kHqIZnTQPkPFccFHt6FEod8hqMhRvDYAwyvczcls2FE1b+WcCs2y2J
Som7MoPcPZiWsnOu7/NTwNpNsmIF1rVzw1A7oem93L10NuK5ZozW6PaG/msxQsXt
n/vYMzFS3mCCeex0Vnuub5VTbNu22cFKbNER09mnXN237x5xhf9GnPno46LsMKZA
4LPClAwKsLCO2Ap4mBoozZAAwpimGTgn9GaCg/TRfqqE0lz+CFBDqwBD2plCDhTk
bGzUG3H/Mz8zBsGXSIWeQMMkCaBLMTonaGOthvIJNbI4JLxXF7clqiwyF4b8a1Io
hcCeRWjVNl2Yt3b+7BoxdIrHFWeg8SHcEYLIuu6NhOoXiwXruSKfbw0C0MBxsagS
2chj00tnHana6HWRSTWBL127qXcFJ5SUtzGkCK1EiAyF+lXkWPOa5EezeIWncORX
3BRjhexLuFZ2fAFTFCaqjb2EcziNpD5WiqM8RJLFd8k43jMK0rzKQw4dr7QQCWgj
k+UvvP563dGbAsZiofycX+YD9y3l8tKrBeSOfncHKxxTEQ67Mmp9khFGueVidSZ/
YKHlIZvyPcANSHvDPvfz00OHchnf+z4yXHeZeb9yiNMSnY/BpeuEiTquEqLw0MKM
CU7NPm9NqZieU8Xx/r9pFmbndNkwRjFwynNdmg/uaJnRNZZ+aAlwBdGKxIfUlSX6
pPT6MNi0CBmNFY9SjD4WPBBQWMdRIaJQ7ULo63f4Ft0hZddwupmtqJ6RB5ckTi8O
enAl8mr1FfIY4VV13Ig3lcVX2sciAPPow/M3X39C/Wp+q43FgUmb75OY3S9YdO70
kGXRqY5/v1ohLArpBUcmQsWjUxeWHUgxxyIEaFGwjpxiu9k5VujmzCMbfeEnhUte
ZupwAiQNfEC/G3dISesjK9h+yG0jpMN4uVSi1cVq91x9iR9RtwIfGmpSv7k2jar2
9ApfThLOjwpBM0kVAJpT6dV7V9vDZYRy8CxbGbxqEaYWtKTlbZHt6NSQTrG8b8sc
XSRklEvMo9nx4cDH2Fh9tV8Wi8jWHEDd1aBnzkk1iUOCSN5M2zoh77DC+IB+pAzj
RnJyBRwFWYvLyHKrALm3u2yoSfz9aN+UBjvBQC+ZQ5sBEGFFkO91txp+5WdMGtaW
GNDoDNyjUJfvK0i2/VGouR9R0X6dLEyxDCJFjYYqEQZUxosZiuLfzUSijJXxKGqa
a8jZdoIbFwDCwvkYsaSCMdw1asM6B66L7tFQw5yzomYFQ1YnWU6mUwFzpG296uVx
86+j8f+h5AmhspIVWmFfO/tx+qLNIMFZJcbZR0doVnSpCnXEF98DOT9q4pGAfSBI
4FtD6zT9Z099htWCb5USWBkhp/OkIicVPWPoVKrN4KZq0rD9lJvmMYSKEdXQ+E31
ymo9zyDTwpptBipCnPgTE2DhrM3hUDXsdiUcVUMqlITzw4qzlNVYjm47z6F4Pue4
9ScoaozjBGmRZDaLlHMc8F1PmxrMoc/MndPjAAR0U81pkgNs5/4gSEDkbsCFlgQt
gM+LfVjLuCr5u+YZ96xwM/gegA28j5qh6Mtc5mdlPT4M4AiFyXiWiJPWn5hHqMun
U0Wwkf9vob7Sx5cGAAKZCj6/AFI5YKooETjpu0BFvkZ3Uc/w84a9xfj29ldTNmqh
qy/vn1vDvHYYmvWLSBGKS8jxShLmeS6f6FPeIF2aOA/Knys2U4qunPqt+X+l1XGB
mRM0IZj4OjHUOxMXPAdXToU074q4LCrdPAOnIPjQFgfERMga7Ya4fvTwRy094+H7
0b90UBOYt3mRdb3ZedSJgQbKlbzh1Ecw10CR7GmTQ33Vvgk54SZI9e49JM3Pqwoh
ZyaXLtgO3gAVlozcICatrp4XjnYDGoxU/NT2Is/ceRZWDUwGMvzpQyeZrhMV74Jc
nt1wylTIfL2xqOinkkNGMf6cMHRgj2lE0Cjuh/WuQVVxfZarxQpMC9kWe1alGuTs
JnrRScsn8nWnbKfl/dTrJ3jSsIqlDWAEIsBlG4N854zbc8jhn9x3npQrihdyj3EL
bDgJJecixRujpG3HOf2pAIGJvcXwYjcjpCyaG06nzIfAVzVtekYhIaulzaS3n2wg
0bkXoVGamzDkLEBQAdiYsAsnbKswhBlf9WGkp+ZiMmyjz4KFBoajMdfOrNmrIGcG
Uq4m4khU5xbu0Qna5xFAVbsNuh0y2PJKjcg6Q2EUhr+MiPBwo1hMYjxkCoK9+MUp
WXKV5LgLXlkfUP2rdXIdvddYM5ZCpNWKZtY3Z0wIRhDij/Ffs6vfQCnFyaUWV8gD
vkXENLWXOHiNeRIjUWh45gqLSvJC8RwpXC0G9rg13MG2wan+53pRO2Qb5KrfrkML
HEMSv5ZTCAFH+QCZF0gJ3N/GaoSPpuSqxYsygWT0VjLsQO12bSEoI9qOjmCgwUsU
59mRpKnitqd2Z2WCyZbbC+PQ1tzFOxijluoDaKWRK7E7tJqSxijm4jogppKdC1Oq
OP7nQ4WmkEuPuIoAIFauqzo8hVsMcTR2KmRTWxpGsQWeDEigvMzrGOtDfWALizlJ
TkTHxB/SwxPVvV7Sc3Tin0in76BIMXa64220F/oN+MWxTyyTS+wg2Si+hUeuToK3
leAF47OQ+PihezAVhIUWsM69kETlRGbBiKBWjeRsJsMjexbEyJ+lYYGpFEYeCIXy
5fH49pi9HsugjJfgcSXeUF4lbLZ+pPmXcCcdo+pgtwQvfiPqhOm1v4ahkWc+P9qK
RVoczVC8l4ZXEbpOrhujOxO6l49qMb4ncN35vAibo8p1YycUC68Ej87tvmzVEqJE
v6WY6J7znpcdFTZ4ovGhhvdqS2kw5yLHFncAIoFYV5/fFMNDl2l3ml7RlmKG/P2Y
uKelIVWVyJXPH9phwBEY+QsM/S441txyeVd1axCpJtTgwn4eupth56afXAIsPpaV
nbQhcBgee1u1bLz9Ik+N3BrcLKVWCY2h/8eDaA1Npllg7Jqo7dqsk0RdOoGbN84B
X6ooSF9matQqmrotvQN6E22fqy4lw3eNnOfq6BgbPKUS7zKOHJ2Ahp2LTLoNVa7b
LVSfJJaruSJxcHMaQoo1tZjNb3s3mWd4u3fTomNJRrm9YsmnDPt3X7bep8n9f1XK
22ntChlzLMQrWYIP9alxl24CuWlFUHsXEEsWuWfSUK5fL5cmhKsfxHJg3Go8yPEb
1PVYklIJnM9NPq+/09zSrteVJgr+9JIVflmCH8i0vjRHk6gZ+205yKFJ9el8+fXO
BefdL3V5dfSnb/AH2P8FprA76T0Ob3IyW8NTZTs2QvFM1wvebTyRmdlZwiuUYvYc
iUiMosYituBWBZOEfFLlrkGvy3uoxAdl9wSWkICiZWgRX0nasczy9HOn9umvii6M
A5ITTp5lcqGUgRhUJWgmATw/Ir6KYYxqHlbMQOFkvl5Pfy+udlOBkcKJcjr4nkcX
3S2+bdY3CWQLzXrkf3kXf57tNy5gwJzrk8iqe3vA2STm+Za7SGjErVRhyvlQ6oBn
0niYkb2TIjub1aBFIi4TXOTJ6dUxIPJM3MfYrxT5vgKfl+fQO7DFdGS9P6JRALrt
zJbPIn+ZdHfYhz45I8/DfrkWA/3nN+1AegiSsNKWo7DPTN9dRS1j2LpwBwKTV1lr
FNaEnzuHTVsdj/isbtEW8chU8OSmuIs4o6/IKjf2KtN6J4zr9kOrBAHfchZNNMY2
VhB0/pSrnIIq3lM/ysu6LXUeN/gFATGsB24o/9mUBc8GpffGjEMKLChk8/38kTYH
0tET/ZxiZTBTrxxr/a8Ou/cf5zm00ZOa4rWivypZ8ii0j0ghNCsivqe7YCvWBxIq
7rwL1q9gWoq1vjjGgT5xr0c4nSroTFBwqb/vO9t6mYDYXqMqM1l+hCVahBOu/Vkb
xLm8IfJrxcy2c0RGkQaQ9RPAZyKbntQ9ZUAXdAR2ZN+4/gNvNsSKOziWlU1XS8Uf
sS29xMvg4xGfPfKSxyMpeLX1465VfOxYooPNnYw3EgofSGyVql4u9ngUzmesLZrz
Vyin1vZyqsd79Vs8ed9/fgRNT7KZmpKnxlEb+q/kLfZZcLO8EPPVUWN1NyhJSnNV
JhbrHkXAlUagdj3AeuW9jzpkpDN7pasYQRA+BAZjMfqMiKcb6NDzxDlmFeZC0/6z
XKoB4KCiv7kyILjPBr3UltekVscqPg9KhbF4vbZQI5XmMbgM+HVtCOVRci7OdxZU
SdMbhUICHrQQBvSpAcp+SpDqcDM6DEvXG6ut88ISonuV8nWIgAEN9BeOJezBLyZY
te9kctSTKrB7cR84pTjaD+2As8WKwYb3S+5t6/0oMmAGKPdIHlSTqsd3qVXIzMNJ
3feLIUXo2KHOvlAyi2uiwxcsO4mKGwkO1B2XZSpCPWn+8ZyE719IjtctGa29rdwh
xmnIyxIeRCil0gKXYxywTPi+H1XeO53vU/vGBrXJQe7UZkF3bDFBg4LJaG4GQLmk
U+dRFwnmqiqszpdIVuUu6MMB+3BcysC2G2rcRgKwvVwRKUMxPe65nMd5WwWi/i/B
2zebbtooFURdWkXVUR89phdPpAJIreEUAcGI6cSmEpEsJyHMqKQQLMjNdhMv3HSi
kFeGwxlap7p1/Z/zsBAchl1SRY1sX6dmSQ3Po6Fv+yOJwLq11hn/uin6pJ5bPbNu
41z6nbPPoa811dBH7gDr/WHtC3BITojLVrGJwt2Jvkx4VgVNGoEQN0wZJVPahSqZ
1NAi/IGazLohdOi68lFIZJEkzlpHecj+7QKG+jq9LZ/yfHi+lMR+RQ8M6RSdhXWD
1hqYu4j+laoMbjMpQpGBj6Ek1xh0+asKIQBjD2oyfFFE3Sz4+Gv0eluxarF5QC4f
2zo0G24LJqFygkAiYJxRLAnDU/kt5Fi1yX/xOR+n1vVNHJPDWpebnnyG9gIZvJ18
wCgB/bXPoe5CzT8ZjUXB6lk/oO+JoEmZ5TfaFm2dhbs4BztJekKXy3DEbuAkNi09
kunXZR2QcAWnRaKKusX+ZEXoeSwaMBnXK5q9S7MF/KjtzWQumL3MhBzhSKOy4IMD
HrFneWeUV+mnLyF16bA+QqxwM8kLaH4yn6/1JTZKS2mJBvIeF1iqqxFQke3mE9TW
WAbOsB4CSCxhkhkJDNZIIIaMPE5+lfVRGLRvKD9fjRdnuCEhRCP+c31YoZj6XBfE
EeIfpPrwkxTf3dzi1eBygjhWqHvQ5HN4qfEyQLIr+Rym9kEOX4TuuIqwtN1af/cM
lAzV+GJPiLcw6SaBJ3JBv1r6AMiAJb2nyLNRw0ghPNF3ZhIbd7Tzb+h5vjmlP6wn
zTJ6vy6bnWzGNpktQi4oEuge8lsBNAHW45Esu4l2FFCi4L5f1vkRt3WWzvho9hWN
s6AIRHJXxQ4bB81JeLAJ7YFiuEXeElMqJzYN6B9RR3xta8AP/da6P/RmU88X956d
0oDVi/IPrF/waPc6ZuSIqDqXXveRdZuJoe9MrVVofRzh0/2CKXAgMDcUq9oR05Y8
tptUZJRTI1xsFPmQMF/zdw2N8ZhALn1dZZoDTujjS+ySni58PnKF3C9dkoWrNKKX
Ss20xfrVJ0Vf39aIzYHkp0NdEdMM1KDIu/+0T0hVUhU2rpUpb3IQN+fXDbBsCUxN
4g7SRx8Fg1CffrDfrFAD2xNBEGVQj5jh42ZelOXumwA5oW99eJYyUGfWlv2S4IBv
SHa5GksyhEz010m4QerGOg5qT2Hz6JIJXO4ebku3h+PetR4mx9l2dmbirN+D/maf
6fedsZd4cXAQLEZqAIEd5LwPoPNNtS//WfsB0KbBbPvRM5QE2jRmY+DLzpj+EGSt
JVrOlJ1w9B4a7Xr2HTioycdWhHNUALrYDrn7mdpOwmw79d4WrfQszASRAR926rg9
4nVVZGocyczK4BOhnMQiENepugffz8NDPQ6QGqEYIjcYnoVioCMRR3WfAm8+rZcj
Rnb39d+vOecEfCbQh95M3A5ue+f9Ou5XgsyywaKAA6x5xy2R0ETDH68bRXwwQ0DI
EwNcwb1y4HZ2KDWh+9XArolUuZ3UuJCqPnWJza74OvRetYHP1bQXnesuPUxSwdeu
p56X4e/9uOa8SNy/K+29SOifKoNLQCA1zAZptOzMvJ2+Cbookuw+4cqrB9c4fFTX
GIJhyXJt18LEzlHljjW/AFIUDVExA3+tAuS/MCdvAGlubJBgb2L5m7JNtIUnAVUX
ViuNGw1W1oA75eY6zej6XlqTZfP/KW9Gu1+PfpV44feYyqQ5Tmh22aOyahEm2YYT
8fXw1dI3bN791zSJDJFdSsoFoodrkoM7GQn3dGOkMPUA5p2mV8FJuOJu0cSE4Z8o
3zUCeDePlXQpcy3L8KS6KMp4sMAXK1Xc0NWXBWbBxW5Wp87wxQdRToZyKKfrurD6
4wzxX1PUw+3ZevhCGH03HJ9R75vmKiWcKOVF3G5++QNJEYW1JfDCMP4UmfHiUaSR
7z+igy5G7zHPfl+1DNgEmi4VKuDjmwlqBY0x/rbVvDB3bV8Xs0ifRk86/ohD3DEr
fA/NVEqJ2NEoekkfALJx8wMsqP1qosh7J4xzjeItwu8i1Y223H0jjVXuy7Pd2DBb
yICzEzqMN8mitgY1bB2L7biaWptKNdDxHkRHBRYi7BJpGBZ4SFuLHTWvd9keBPc/
zOmfYlTyhoHO2vjLwoa477BiBPxNn0jPcn2XtAuIX2Dxq60nsivHaPrsTfxl1VV9
FBstXx70ihv03XJjpYSyixRSxamQRU2AhrKObx5HdBfQqlWSuGNqMTIBoufFVvpL
3DURckdALWF5z0pjsobzPpI6RbwfBJQjW+Q8yZ6YjQ5PdgBTIQcDpDQrIJUnoxYR
yo/dJ3uhUx/w2EgZlE9XeQ3AX7tc+JSQOO1z7Mxl2KfB5hs8P4SZNBrzbkXya1va
jBD2t4wWl0SC6ENad3C1PsUdtxQLFB3J8MGug8xdzpLsU0bhCLC4Z86dGyIhcex1
ur68c+/jfSO/gQUsEzBCVaU/D1LZo+tmN0kpUKvd6yti9bLKxqQmyZllcJ0YGqKW
18AOozdBTijJbSfWq2CxV8IBBSIPnl5xfY3iGpLfyjKfOEZvP/D2coYEnaz6jdk9
yPuTGOBAY/h984wPJPhzvq3YAePhkv9lAOSuR3ird54u4pHS0M0yMxjeutus/gf1
Nz8fZuNcm0IB01gDJp7T6x+WG+gzQGlzXGgC4XkyD0ceT0lDLxlA+41FI8aRqS3B
BKRDzGhvSUW8+EQ1mULEIZNEyn8dgf5Bx0xSomj91doc4frBf3BSlCGVtnNL9gcw
cZ3O14ZKCL0dYeuOX/nqsjTtVksjQviPG3YeLnJzjGrFfvbS1Mwn/0hUKAidFe+M
qkTly/2suSyL/CgZENtYcIS6UlkMhhDSv+Ei/Nb4Al5NI8GYr3H3RL0b56ZnYWWJ
8S6m9SyL4Pd/Xy7SvMalTAiRYydO4wGfER7GFtFc88Mel60zbI/Ac4gksOWWAz1U
5rMhz0/xWXAn7Iw4R17KS/JMLlTH4nlZm9rcTRxXZqaBm9Ecr5teeAxqkJTKuA3j
UwpklkeHL1dd7aoFeHsTSOuuK20M8NfMQ/CPUDaay9KdJXuDs9BCUXL3ZKjmVjaO
Nn63bhHwZb9LbkjEi22FtJ2V6GcpXOAkav/dp9jjTzuz2DIS8LSJ+zv6TxfoRtL1
T/FUmvwxxjQSFJzUhOT+0JoFE55AlZ6sm8IQOn587XcvytnwLwMRWQUgkPl0MN57
Pod/gHwliHTRsoDt2z9XkLt8C8xhc1grepLPLHiQArHqj0RyaSLQNuNPygLY+OCh
LmnUCTHYz254y6IFJ97vu+hIB6crBv0QlFw1BP9n08ZpyqXCLb+BikFuk024K3ui
nNbebnHjljrwr/useLcw7vbxxzuh12a+BaOWaglMrfUG0evNTf+4CEODiMOiPbYu
T/rm7+A84pqs5WnDmnJbHGXxOYEWvkoHwZsrIBL2JsSVjRKf/awAtylhRYz651ZM
XHa4VtRuLqybnpF8oppXx/7mCXRoEi1m8CoBx3bKJnooVdsGGpxgtoUioHS+C677
hU7tlAvIs2EATrH9q5v36WjFyPReGT5B0f2VkFUl5RB2pwkpzRDt8boqRe9paiSf
FRffrNxbu6//G3G3iw4pfwMtbIgFgwrdv9Xo2MYIPxTWWdd32UwzFQ7dOrRK1SGU
IHp1aHjnZXwYFfXPqKKpF4TzSWIFzfTC9imkTfU0rWYcSR1ijHcsL+7x0VAu7goV
EC7ItKtT4U7qQOPHW/CzQvC5+nGjSm1O3hDzPYmDFTA7OSuWEwpKBg5DYFI52TP2
xdK6koqOKJdHNPhMQL1qN4aRobnRZ9WKtlvxfvLS6FnSzXAlFPkiCYnV3gPkk3XN
T/YP5gpKxChP7dmpfYFIY+1+x01148lOLBblQzGCMoWJm8lAt+Y0fby28dGIeBBY
Nbe9fJ/pXbue1VMNkmj4qCKLD2X/O15rtHEgVXzvD5TdcUHoNuoUQlCwFNvujJC1
YJyIHF9mrS6gkzksGvggu5hp1G7VafBpDaxSODZY7hO0FIlPSwH8T4aDZ713effb
DrSX8droF98BpEZEeIIbMF8bD/r2SrrDd66xABa3VLzMQRL4+Z5+x0y4JJ9yJn/a
sQJQ1gyjg48/wCa4IcwfnbjzdhXghn/O0lQUOf5Eh26nXA5IhIoWgZURHeanViOt
0x9j7TPLxK46QDMJ6EoP8UgmoGn3IcFFO22rFKuc9jaHXig/CNbrv01/Um/1vuPl
6CsASVVkPM9yFP4feIR5LjbfJ+9YP6GSR+Ic5ddb4dKnS3qHSH+rOlMRGWVBMGZh
lDQYNH82BGZ1j5vzHWKWdwzn3oU05rnZy4MupPsdcGj3Gfu/9T51Oc9K1sd/M+RU
VIHC8Hi79e6PtlBivBjzVAlv+or2wUS2Yl7gVcUk7NAPlh4QTMiB20JPGMhAQSC8
hzuvghrqhu7vhbRcy68LiRPu6Rzhyudkod76/F8jgY0ol8qRM/VOafQNEvFPGDRw
9pz/0vqlQxPGfMVNZFAKsKJhIuSAGCYEab1RP0yMoKMvQD55s0ZvZ/fSI1xLr/xW
xSZhKS29UVyMxq+IUT4hBX388r1G0Z3QFUQ8aRjeE/++VPYOcPrNECcVXuoLFO2Q
FC0d+NsKo45LZIqYXmwwdpV8jN4SqQ0TQGmr2uoCm7eDDd54culc+phxn6ohwdNj
x8vrqTk4za6DHGMF9tFIWMx4qEL1JPftVNeMFW2QUJgZBD/MOVOfp4Dlxt2G3zv1
mh5ydTMHjNSwD8Z0mycUkQ6yrwsY0CHDM0gIIvi8gai5TuALD0eigDLvoIQgXrnJ
07Eg3j0sf7eYEwxYt+wy9qcBbS6XPK3adx8Kj5bnw4DaZauTelyyIqjwnPG9SSXm
38c+9F+plTC75jsHW3vvft0Fz8pasx0Fe7kE6B/cf/uzkXPni7hnOyHUwb3BuAxU
vTxnnRffL1qiqwImTJ3gL+DhNKIPJluy+tMU754y44j6w+2NFcNymr7QbAEkLK2s
o/oSU8xy4SbLk2k2YCrDmNk7MCzM5fyDl5cDwHP0y00EzIxRKcK3Yw/W6Su9zRgu
d9x73ktCzfVlP/EpFPsTN1xdk4PrUH+3qvfKT3EuAnlFZjbx5Opk3/K/Wscgec2E
Uv/IyAvFp4TiE3Wn5/5XcevXGQ40VqMk2Ch9bTt4JI/Oq3XAcY/fykKJUPsiqhC5
HPJj4x8wlDekNIX/qm32+ZMQIEwuZzIMVi6SwFXi7fV63rMW2Xiv2z5uK7cFFewJ
PX2DzMEFMaNCi67yPhOooL+mDPxpAqfhu6tJruRwCRK0cjlJvB2Qsg1RRn2rnYx4
T6kI3CuyiK9epPTM9nzQRq77NsrLVQf7vPnO2K+5nl1Q81YuFFJh1OdgIeyinJiu
yJqBuIYPo9JeHdEFdO+pE8o71Z4sOuFMI1agy5G1yHHwxuMRD6VlOO5ju2cT9nuw
3fFVt3Xkp9Gz1emC3hkqsu9Um0Qv1Aq4o87BxvoyDhPzJj9ffGqCnWlkP/vZyedi
lkzeziVFZmmusmrnXUrqgheLjtLRuh+5kuN4w4G++Zi41FDOitSadUNHYOEkBSX8
3ULwJNIJYZdKN03undPAxBqf2qIXpJ/05pqxQwAAhHepf6y8xTvJk+m4XTgZOTVp
jsFGinAA6qsF7xz3XypmpNaOmak5OPG0PVvPhSjMCLLbNYZeCeOuf184iJ0hD7kf
mvKuCI75r2O+vaOxLdarc6KeH4gMKdGyrR7p1FKr8nsiMflViq2rj+cofIIbxNHY
NKQAw3YkoZwAm8+SNcw0KxoT++cAudvmJ/dXdnv8fA60nlIrz2ZcS2+8Mr8ibm4s
LGWWjWPcLc8WDZ36EkUhuSypQMk+vrYTvtUpXkDfl2wHbTQO72j0UQGXlAy/4xIx
krsycWXmCorICas5XBDxcWpBOR39moDEe1rjnkEhDGIAsqzfOdoUZmVukl+OF6YE
3W+sm7rvONOFqLq4/P9pik4e01eWah2zf2XpROCr2XXskt2cdre/qxbe7NbGF/eB
URYFMipa1lwNTBC5Hz0tLVY4aXx9v5VXICoOmJl/ir/sAL2xcpoZQn3xF7njukSd
GVWJid15L2MqttB/k5znSe4cSRuBlNmmbnxwaP0gbqU5Ba94yaAMgjhXVrcPKeTU
BkpQKtBSpK28QHWaCG/sFdu6WmL90s/zMvxENtcsP7OZdgPXs+Q3NAunB6456Awb
g0zlrNmO6XF/OGoaSvZxT12t5X8v2RCFOV3nl28wZwkSkQr+OHtdUEWxwNV28+5F
0TZTCuvtfYNpS/3SxiiH5sKtt9p1KtXi5CEdpftTmojbUsxdLfNSiE459ba3ahbu
P192V+HdAhJI51KDwZ4vBmtex9KYdNWzknRpqEeUx0s28YbD3OUfbfef+IN6AEyQ
PVCI9bt5Ot0GAs36qQwSfde6MO+pG3/vWGdDzFib6lKEcXmDIIdvzUnzi1lpyT/g
ASCiCjiQUjO5wyZkUZvnndMkNRA54xlUzwPSY17HgJj4yuWCdxKEXSh5e6VigJ0x
1aP4RJNzKX1HvAZLBu/4/rcwZwdBGl5yt/mjCm1GCDBliYWbloQrg0ZJhH35tGRL
ubedDXUUerJz8VFN7T5/PwRWo3fy6jRbN3G9txC2F/Zd4k7NFCOpJkEOcW9S35Iv
HuZN2qUVftJEDh9987999QBTkuEUHCVsC9EdBYQYzWSXAn4szHHp/KSsmOW8v3Xt
9qpkIjhJOUtW/hFyi92juUEk/CevxDjfq3YwUocd5aEYNtwrdD1KhHGs8Au3Vwqr
yyPsM4ZPeGa+/TyO2jSokC2XQpO1TSxnoPcMPdoJcihDllE35hefJWWRfpDBYm53
sOFMqMoMVPzi+PHb1V7aKm3wsuYUAasqli1j4+q8W5Y7vIs0UTjahvhBGtTp0muv
+aEYvCUsBKBNCpyHNUcw+CPIswk8gi7QnyF15KUtCX4sX10VPnbLRG+pLqgCTm0s
68Rarcl9pdBJV4jDUbCOtjb6KAmf64ryJOkIFKmqQ/dSq9XHMUykyoaco1mTED7j
Ed8U+X+x+Ob5BS4S5s9W+AA3Yb0b89B+iBZJFkVeiwaQDXF4W2VfEF1CCTy9KtNm
k0psMR0FLyC5qx6DqqGNgFZSPW4kbp3eFkW7KZQ5GaVlzW7SRyynYP4GGB3wIrJg
mRiu78gDfUMOqjNdp/9njCo0kjIwbp/5w6mlndjkycc7LjSc+isfOJHwNCUNzSuF
/ONGHimo12WOdYudO/qZZ7zmUY1rsxVjsqp94FTDj59/czE9Scw6B93lrf51liPO
KBz5d1+YsjNSybPCltnhvM9UBSayokEzKx1OsarNZNoKCJpbMfJOchMjgWpAUK/g
kU7uwocMR8efxSLwqknSmxVdVtN72JBQRWXBRh8uG99NqldWjUBr6UaOf9ursYIF
u1b0ybM7xCUP2DBNpWsCHBTKJKuQ76X7IS/30xiWZTRXP0oW12lR2ldv8tZDcbLG
J8giayMQzeJo7uOg2UQi2v7H6K9R26idWl4F8Vbt5upc4bra73ixDqQiUL7fsOyz
usKB7WbU1DIBQrSaf2sJc4PCUmxcumUIzdTrIgdy5dM1afIcithXV6K8biFL3HG4
rS7aOfjwN0PqhrcPZ9kXPH0MeO1anZLgTLBDTE+eVQZy0P7tv2OyfJJ48uw8gGME
sL8XriE8Y9KZcMEoAx5ynZnp1csVuOYv0TNqRdXd+JGh+og2ytDyIl3rbp7rF/ul
gn1jTOcb/VMCpjubNBHzZM5mF1XsfRjNu/HGg8Vcj7z/2JgwZ+ExC2DGNyFsGV/s
eGak1ssODNL4nI2n3bY5BBWYQLF6eRJQyEcv3Fw6KS7J+5+E37evrhAuHzWwaxVi
RAHSlA0MCNDxVfAoO16vrfhZH1xfBqOpHsHwgG3dbDdi3yJ7m7gFvIs67M6ZhDtx
7xT0uNRKBY2c4zn7j5osQC6IrOtmgZiM40vWQlO5jEp1ZR13mYZM9zRY/AiU5CAc
l78kBaYKFKCFCyvz7pzvuAZh5fSZaLzW8Tz4DeDvL6lUUL2lBG7l5eKpOFv8F210
1EP3n+Uk9QNi1DTFOnRzN3RXmJj7qzOjfdSh3IUQ9o8qAA6OTyasS2MBsnX0TAP1
xxpei5FSulGwuulZVVxLRH26jrY5IrqzKzlM+nKmTVTJVrtDvurs1eirDkD0/xVD
ZKrn9W6koqoh3+qmFsuanHujh2mlgDVRD4GDJtw3U6wZxZQ3IjLqM33cfBIwk/GE
DkB/WuAFTPYzL6UmEX0+dSNpnCAY9RGRoX03xzxUEbg0SiLOH7U7eLr8KcIU9wZt
1g/cZAyRTz5FdOqSILXzoOQz1sHeVkC5+1jXR8IrB48hrU4y5CGP1VvszUdna+Kg
PmgerwpSU9ZsoVnNcvMyG1mqvZI1BmwPhuIlWmviK4Rnb3dq1sUFcDSbG+BnTcFJ
1pDCV5zPylgrceC/ikv8KCE2+E3K3Ize2qDb2MPGekP93UVPze4YYncTC+XvYnAc
FSdqW6xNyNB0SUaUdUwZBJ2LCRQ7v+D3aqZTgkNflIJqUAh4kkXRkbggixp8o1YV
QwjVUofHR12AkVne0cufrAYQS/JCLrtQ/SS10PdFHOg93ca25tztUa1Wjc84c9ho
x78l/DiE6g3lLES9XuP7x+0GQnqkr+nuhZEYVQ0Dc9Cl4UpCUOIl0/roAE7zsbSi
FdeNkwAnIg0RcHkH5RAdgMhP8R4CHieDsbEnLVZUBz/Ap1tSjEic1YjUPyCeMnaA
ENVgZgpTk5bxglvvohOTAUKXTRHvDNfbtY34GGjL16zweZfT/ehgtuahzb+RW5gR
2IHUQTm/Vg6Ei+hrIsf0l+hbsGVwZFgHHitMSFIoIyTMHCPNDRYWNzNknCGgc5T1
rJzkn9FsqAjn5YOwN9qFEMq7I7CkYw2k8390VBJtyQfI90m77wETMukB2q73/lMP
W40tMKLo4DpeQRITN+W7hAjd61bopI1O1FZpG4EIcr9MCWPxX3R671LrfU+ykVxz
59vZdzOf7LhvADxXuclt48GJcveCT7glNPlTHH0t5kN6wZzkm4E9TYyrnzHu5+L8
EXoYbkBiYwJhAy1mp6zU/mtJRW9/HF7Eoj/rh6POyVhOCW9184G5qNYdW1Wuu4qE
VZZDE1IaMHErx+LYK0tEathZODgKosIS1QAUbeTMdyChiZdVyTI4htJMOE+FTXH0
yJGo9ZMCEsQOMzlYZtMh/tKq1naR2Yk8+4McSrPXIPND23W9zXo7ZLl4eK1UnQ/Z
AzpXi2jz5WVmfh+LlvoWCJBepM0Fg0KFG8jAna/IbKeDnKzIsL7S+Ai7vpW4/mTc
GHcorL/dlAx9wGCUGpugBH/bcYBaHM9P2z6u29C+58fRm74HZjrHaG65jbpwtIOA
jE71hCZJVBIDdO6d+H9rN0wP2B0/QlFCOlVBGsvFwWr9ASVBXcwzUyOeSFdTPVua
RzWgqDAobBgSKr+4x5qNhwm1L1bx6rrkU5qdISHEx6/Y6u/O9QJLSo6aiO9xfYve
XDIt3+kljASzCtAmgVh34myy/lH8Cu4fUnZrDuEEO8BIGOQPW60g4KETi4/JVUKk
3VB9B9n8ebZo3eWyBJ1PQB4/Fna4vZRJqQ2Bdb1SKjo/eWXvbLFsn29fMQS6r7Fg
22/+yMAJJAgRMUr2kTeagKuWjMsKgrB8CVwrAaffP1BZgNuJLh9rTUqM02p3OFn7
smWIka/p+x/Vl1OLQuLuP6HaCUOW1zso9fBEAgF5Pp1kHY5R0YbLHqtdrxKX7UBu
HTzhcfbT43BhS42DztSBwOsAwoyAfi10bgde4XWlPz1i/9cQOwwcIbOiBAWsVPDh
9R1/erGWTOHRAJebI88pG1EO+lusxhaW1JSnoJYVggJ/LrEJvVGB7WA1TdFtrwzT
7VZkpjQHyJH5ehwSf0Zgxuhk3zgy0S6kbjKVq9WYrCS0U7o9x4OIO6B+iSmOV6+F
Ok3x/HrMTdPY3dICUSCAaZY1G+RwDXM0hCMwTqHitEpNLGvntCS6g36dEVC6Q5Zr
d19KSeN6z1Vgwegkq2Ug4aD0dRx3LNQK6J/KIHh6AgAw3lj1U9lY4wP//zKTAi3Q
V9hCtlLZSgO1aOg46aI7XnvG1kYQ34RXhTiIjsWNu5dcVB/7XBiUiKOkmGgQqnGt
o26SsI6xgiZZEY3QUIANgcG3ln0NspaHP/i++yYImv91id51egxT6n8e/uq/ahHH
J4vZWFSPGdaXJnxK/IB3HHMSD9hlZ6X7WQuQKsUiHx35nDNsupsBDUQPzQBx1qm4
EDc/ZNqvTH42a3mzW+hhTQFhUbieUef18VPMgr1UA4mp84mE1RP9ZHzfAL64X9JD
mBjipxohfGa9AaYyn8hzw2KaRXvKJxWFua3ZiTvxec7rsA7ObilXtSJKQVOB8WaY
Of1SYUmZc9VpbQ90TZ40uCHWzpmCuB2dWREOT9/Vq2Xe0Gzxs+yN8IcaoV/FC92G
khEStFSsoMehbnASB3AIiyz+PfXpl5EP8c81Jr/NrdoyWcddZR1hO+t5SzcHKdgB
J7NzQBifW0IuilIf877oze+ZO4zTvg98lsxIxLrBNFz6XdmTASLmUwCA5eRZz5i3
YfP6S84JaA/yhYPW2jeA0PesavbGDNO3WNYPBkoDdLuxG8KYLqTURfKklpEfjBuA
looEziQAmEX/FFML2jusV7BDi5dW2q1gRSjr9G3ieo2NV644EN5q+B3omoaMSK79
q4Wfan40BJBpmXEoXNhiORyT+hrXLU6NSJLoOKJ4WFhs4RCJXOjb2CN1Wt5yg0OH
E8Jpl2mVvZW2QGNG3lEp3Z82KqR70Q+tb76xi6TreBke2WjNusSVu5DGATKcV07U
OAZeMaBajdDtnJiB39e3xcfNCoIh2wDGBSy51JhKPUVf+DS6TdcRP1n7eH5d2Ezu
3IONdY+a+JqNmBroqMuQg3WJE7PDv/LEo6IP2s9f9NaK4JJtn7JpILlbkEZs2Vva
JPiCr916PwmxmGk/3HxgUqgQbrQMcklwHtq5WC8I1yzht40aJVPPFP1sod1knAIS
O+Yu9kjvSoq360gOTV5s9EC0Hvg4noOkkEAg+vV1H1cTMsickeI3CJ9kgI1GBWwX
3CzbKly78Jnx9/a407U+yopBp54OLBEPdeu0+qxkhsr9DSYMOi8y5mqFvoeoOnhH
3HbkZco/I/Xm3tXYk0wpkrUc52H5a6h3plVQf56INY+Shzxn6572XDcY1sK9YgoB
jTsWcvUQgtixMu9kmCImRGvmDFWg5HeDgHWZtZ2OyK+B3beyDIA/vsTn9CN/dgV5
wAQ34Ci93ddr8Ju1UAXp1cW0/x6y6nhyp5viXGnmzyRtFQL4cPamT4zMYaj9/UVK
cCTwN8CQe+Sny2Mqw8QAH+iZI/R4OeQ4w3iK1wTAug+AgDFWPmMdNRHY8ttZyZjE
WxnCz/PjWZsEev6TksMIqOG60/gKB3ZrC5Z7/CeESL2B7sTnJp9byAaqX+StSS0r
O4yutb1/M3PN2OKIt/wcqZ+GQrYHI5IJuwEocO0zPdd82rK3otAqEvkIe7MAIYC1
S1pC9UzYGT/9XFk28k6dkEXxXKlzhdY2mDfECbCnFCEa1bWF7+RxJiath+0hOkrG
8K0XmQkEL4HNVBdDzc5hFSMS7U8GKRFvHFIcwGHPin1xGF0zrfAN31jT1YUVhnAa
xuNqKlnSTH5cFAVoDH6B0R69f5es9KSfKZ78p4ryMPgiborbAKVbMWXAS/VhNVKV
Ts0JLgExjzQIJCw7FWDjOTASti2KLhVs5rbfo0Pw7+zsnCXk/VzmggLIWu7JcLP8
hrX1qPbr1Gv1WQPMuytRQXBkpTv5TjZyNngYOiV4e3W82G7NsIf/vj8XTlW+vBgC
7gN16Y2rqbzotP7q4bHavqfuvqTtlu24pX9PwTihVGjzQGStcA9StDsVlovnUPZf
p9XbwcfWauTcqVzeJLMWoW3X164DBD4EVZ8QvlwTEr8nc9be0HO6but8QQHAcd36
P5Cg2BDm44HffxETvlOIwHwjZMahLvjA1DYl5j2WB6I5Hsoi7JFt2wQ2ytHhc+em
BWgNSl7p/EWbZUIUkoLeHY91PXhKOAw3xiOefCmhKI3KNMgs+19+e7HNQPOscEaJ
9sZu56lNNjbEuXfMUO6h5abOjNxJ3r6mlbMmJrq9jSEogmY+PzHANMWXgct67xZj
Hj06DofdtRRhxdYmVNkPUPAEzerE1hI5JywLHG5ljlMz8uplHys5iYVDC/hsuI6G
nY8L/6QG0hFIJrXxkQsUrGWz3inCkaKgKhgx3Ueg9d9gg5RSCKSNn2lMVgrQtR8w
NyhAvXo6Iok1DsYnaJIgIUgqUSaFAZRHQeTK99pW/v+BKgGXwNUWspkevm0DaN45
DMvz1GuSGUkNhdz8Vf/Pf6UO53UA1xgx/TXVSATtCj+nYBCJvmrQsW0hvYIEXKlr
VbFWfMLP58eCMgB4kzWpfg7capE7KslKa74IGXarmmLRuvph1LF7VyETkVDB5CDC
lj9Vb9KljA/2FCb8hg5SUFYoTAd9lszdsXemNhkK4g96LFH/f96lPbdbNmVnBnzc
Ggsr5mffrmRlmbPAdSi/YCNVI9jgjN6LkH4CXfa60e23PuuoxQGECyq6dwVwhwab
n+k3fQJTDVqyQA7MnjuccyIxz7imeYgVbAv4F/FPzDzhqutYP7TzVeqKzMqFmk7v
RlR+mqv2bA4n1mIrejcfjlJM5XQUfEF0+bB/NtZngVmNMmtV88gTVj+HoQcTgdOL
adjp66LBUVolex8BOm/yfAOGvX42VYoyWtnYPYgQveS8Cu66oo1UjiPxHFKXdFwm
4CdLV/NlwcOJodt3QpWExIbYDvFKIOl6Klslbu7vxdNgkY3iUhj0wuHqIRJHHcXU
QTDZArO6I2bNvlCj9iHnFmCEZm8005ViYCtDi8c55l8PkNsxO80BgHYesGkbU1ur
+MHay0+/m+datWMcM4Ubkur75UVetPqCzgv+0QoUME/1jrJlPFApVV0QtA9aMiiY
NSD0uVEuF720yr6jUM5LJuMuDGujRTozpH+MI75bS2QEJucBp7LhG3fUNDfRpgIm
U1fqMgyyAvVLhqFn5heZFvPjh5We4wHLV4qXVqaBT5eRWxxFckqX8m1ldjj4fx30
AoWpwwEAuGtEaAxeDXtyuAoZLe0hKKUwkHYbRzPKOEeYt7hql0Y/PzdgiTQCe/L4
khcZ0wE5Cpz6Jjf+eK8iOxx9T+R2ZGt4i6KSPRW4eEkfNEIcY5na/obfLp6gsc1E
JNgCXM4Jx4S7mULMEr3ffm0q12SSWb6HKQo+9TwBQ34sH1mwFh0FtOsw+yUslE9O
uFjscMBxhaHe9dwmZOTd4KlPmY25x4/ppWMROePKcCZnuarHdgMz8QGWTAWHwJIZ
B+O7d3W+4zE9650+npwfWoT1Hpy/7ivNfJUjMPlsM165GP2mUeuVkQGCGR/uaU5J
fuJ7KXqWYtoOT+jdSloBZvSRlxXLfivwtqkpBJQ3DCX7MSlHAouAY9hru97helKg
DbB/39vTC9pQXqb/9Tk/JBp2J51UCqg/D9r0EYYA7eGg/QtPhl3UdnqoABKMbHso
+4XL3aKB5qTR/PO+SnhFx/BVYL9Eo7nE4zlgSMal12/jSEhVSCuqeXH8Jb7VIi2a
Gdi+3Ve3+Jq3siBgh1BtR0aFaCrsYOoavzNntPq80M9Gp1j0yd1gNhNIpT6eHx+z
DPJRlt7/X+JSKjTmgTDpIT2OOwMjh2vNllmM7TDiMTicDw0s6vsXkkImL+BwiOcB
Ls2Scxi1LZNHUJLq9Lf1xoM8iIMeY0Uz0oeuz9N48WGPsdKzTCrN/hwSaEB80Xh4
WPXxLMUP7S6Wya6nlN3Adb6As9tSiqQCY+O1wYDmSt73ZP3tGaC44Rg3vjHg1qiT
7NVcH6kEz0lfSB1m0rd4A2pQdBTMu5LtZ/Jwwu3qeJs3zwMMQQ3ijh0hOznV/vAl
FX8mQcqpmtQ8Anb7OwkUesbPJw5dW35wxZJ3xksS88fDmlfbaI6DI7p/Lg969qpX
9t2CUG94WzQ6U93jSaj8433IypGfXZuUZj4jvDQcCqDzyTFEYAaoHMemy0lGThnr
kXbifYqx3eBYf5jpLp3Zmt75lPMNbbspN2Kx/f+OsRSGQrCBU74g837RaZb7IZkC
zszRbTHNaJ9IHG1YW9H0aNuzV9uEA6lHN6RS9+MKuHR+imNgR486fX6vxIrISTZ7
1eZ5lTRniePe2oJi899P9W8vIltyd+9IG0nH3gcDkXseGeZbkqtzZx9unccf4ais
IBRIh3EX5SobhOowVyr9L7FYG2Peg+sMI93pbUncu3wTZwIoS5tBLKMzK+Fahine
7IEIQxf/n/N5yrSpFuZtuFl5JgWy7p3VjJVDCIzoaSJyi7XMmImY6gVylWvasi3i
6hbWOgpUa/aJFY+mIWJkCBZWphDluxoLonwFyCufDkup6fTMk0HWRBNXeyQprM27
4NvwuKs0h1wy6/Y7ReHuxadr2Avm6Z70e5fwTKZ3gm+VtobxzYO1cj2r4a3dL+by
oe358DQtXTCtzPRGdMb8OTxUyV4X4WaXYBcyf8UAszJ9xlrxoGhkjouQxOkxtiP1
b1bD5dhjYbTMctDZgDWz0GQCO8OXzJwN7azPnsiRQu1LqUQjtCsqlYOHDlH+TuMt
PjJ0mAH9m8PKvPcHAZn7oOBxCltgXzoEBnYAHYCRaogipCNRIRw1/vaxKMPvxndC
FsDF1RNf0T9VqvTeuTuLznzQnE8ECjDIAxuJjUmoPH41/k+4XpjDPJRyUYq7asZj
9BJDY0bPS2+1Fb69Pfn42BCigvDRcfsmQJPpa0AnZYydJroq7QEx5kaO8ReWfgmm
6Cciur+7V30eqQGv2hvvhYEsipDfzL9f2icLtIPPrBlSrf7pYapNdqXFvIVRwNsK
L8hU+ItTzhC9B71QLJr8O7/cUiDUw+owMYhYV7YSx79Zut6t6kMJQdKvee2YyP2e
U7fMRX/fT+cKdlniesRtBBd970P7XPeJzO2kZHqtr9/pAMzAEe1QDojLDQ/tFYNk
X/w9Rwdk9b1PeJNYqoZQIQ91UbICVdcSXPodipZ6NGkydUq4t2a/c7Hw5DNR9LbO
6wNzOL3ZsUDQ4cpHSUOE3wuOzqVK02w/rjm1jaQzqLssmD7frocLKyvg/R0hyd14
lDVaTXUKPn7889Yo2XsTDbkB1MgI40vfH/3s6gnbzt5+/RxtDOlxTK0NTjIfW61d
gAbzUbmpbHoHX2AFpuAxORBBkZNINFj3hV1SvIKBHipbNpkWLvzm6zYcNA1D80LP
TdHUZthot+1txW6jsciTHFYiVN9Si/Y9EE5wvf5gqPLKRCy8xmqHRDVpfk/H+dm7
Wd+s+U9fwRVbu0SRP4zoCgJkBu52mLPnQgHuUyBNl9spfkd/n2hjU7fOK8BbRKzT
fxIF0Pmc2CUcdf0cs7sHYRFnN8z+Vo38YEPsPQkEQKFlWi9PbolsyCymgfel3+95
DHw3AxUx+aLpS9UnAj4KGO+QbboBQjbx1Wb03parKxya+Ce0y0pHNhBPiz6vBtZG
Kqs0A7H96Y/elX6hfXZtSVJ4Yc/2IGvkd/MQvtbtPj/9uhJhwwpIMAYC0SemaBCl
+GNO/KbbxGP9C8hk6Ki/UqnfEaFwfwrXTodpjjTQ0679vBoHXyAmxB18a51wmJ5u
jaChe4PJDIi/nvPyZjtY7cP3G51LHnig9NHjvjJ+0ZE1zSg7VuqWOv0MM6WZ62mZ
Ck0uzJgBbrYSKZrHc4ZHk3Ca272SCjXNPFVKscbbmWxwiUKjqKlJWDsKlQejUZD9
KUgB/qJYdewW9jG7x2gilcE+tWZiQtGULx1jA7XSSwB4lQZZ0qI4Wk6JRjtvGBku
4DIKAXMlgnV+caBnKaL7liNZY2yRDdlMAHvScyrsgKYODPXfHodS7M0pxz9DiywU
CD8wr1b4b5jCif7MrQKvwFBF2X2BX+XBLKjPGz7kvAjmtyptpD0iZmKIXfQozM19
kkU318WSD3Prk1ZUAj+fkfJLgLMtoGRn3Kue/DVHQb1tSnUYjiWprstrewnZLThT
qLexXH02kQAOU+pvWvGkVbnERfeaKu3JK+of6soykfqJPkut+0LQaKGzK4HKd3hT
PtczZbFj0SkfOUwAPhADsUSNOpOLnjIV3tq8eGUc28C1eDPsgx75Uz1EvNgy5vJ/
10wNsEmTVshDfhH6RoMybIx2p93zF5apGS6K11NYzd20EsibkSxJfA9qoXCf33eh
tzFTqQT9m0UD+OxYBv5x8+55ar/pAhuxkpvlwBKziGexVZvcwnW0Nx0QRUd2BvYa
xvNQicPTRFzWzkVZcRg1Y+TnLvgzoDFMP/5pIhLzJOFLQ79Q5ansYpw2x049UB7o
ngOnFLWR1qJDrz699Yti0L7ywOzmVO0T/HE0T4PbTjhP48+o0bcU6JYaIEdKhJih
5fODxqpQcoLNKydVnOnmBUxZ1mlUiNvxcZnDDfj4bg8WkTxQkhI1lenmxWDkEcAS
3zhHWCJTFi3NzECGYqA9PzbdQKlsHWxZfykr5dS0DkLYIDU1xilebmgdaF+gX7Ex
V9Bm037BmJNIZjLIOKwlSo1rOx0h23FwJa579eFyDer78aHC7R9Ntfaqg+HQmmOJ
DJvzDKhW4ki5F4H5RPFd3/aJdkgLYHAI6YxsTRYnYJtHw//Ez80UGbX3b/dpnHG6
DvoSO7JGfg0Wl9NiGbTDG6HenUadd2r4lx2C6kx8Jvo2wZwrtmIVRqB/H+xLgQuR
O1GnBfOqnm0jrxS9U+AHcW4DCtnLHi/niOwWF6JI8J1CyZYhoEksRPS53M8BDu+z
0mwqPy7GKwZPXmPgLouLadjOZsElDy6jUGDjgm+OFnRXAkTiVB63erAzarbXDJXC
3xocVUcInV7KLMrlOq6x6MbuwrSTJUX9RW0OeWgmMLlf1Bq2vYTPJxCFLkVoFD98
PF1Hb21lSrpYGGm7hS5UIQzGQO5amj/aAaBnVhelfMfHyRHDQgRc4XyYkzP1JJfy
+PeS8b5NHN/QDKZCLXxdX7jooMzv9G8MLa9jcA8/MwzeDoUowTluctO4smVjTJdZ
+NSMPvXAiaDp+kGeB5XFBZPYMxSu4l7migTfeZ3I8tu7BCVUD4eBknU6OfgPmuCq
8g9COyiTaMwI0ByK7a8oDLV9VoYzp9X4rWU4IgvtMUwynCF2/V/X8wjar+LElmns
5xKaraP3+CZviCRH5T5FBkzZYhH4d6nmZK0u6iwoZRxqllLbev2PHbD3LXG3XhVE
H63UxNvTdcm6Qp0JqkgzajFr5EbV8Fls5qu2NSyUGAShp1yA7nMMdjIkCODHTksJ
p0uESortNYgUjo0qCMTvqdi+Jbhm5GJZto3H5fIQew4WSzxizwDjtifbPJqlBG8x
iOCXEreaGq2Grhn2SQbIjVM9BDzgXnz4YAhRpqsOWoDC0C0fTTDtC3yrLB4qKYsl
yyr9Ovm4TB6AGUJ+YgScZ/NjplJ9EHRYrbSQpzAyi+JsSFhBQB20N/fsGV1iovcE
JSRtsA+jEeLJ83YnfUKIF4e9Xq/LElbbdLlkGXJAvtPt+j4yTpT0kjm/nIIaccxJ
Qk3kcyPOKbPQc1tGsTZaVgmswTFJA3XfXawuSWRXtTJ0HqI4IQsSb4psKPhdVBYV
ysdj2OkGw/iI2hgnrgssn9PsTKCFtIA/WuCOI65W7EfdM13Zoc4+Y78Yb4sUo2gU
EbzoBWEVA1NipCtfSJe4YyhKfLaPu7iVn4IgEm1BCgKHaiT74B+S3yOhiZcAn1an
sg0NHR513hnL2Qy4sjbeKQdaj+5BwTvPKIen3lLOaOJy/aAj3dwmZMW1RVK0Mg6e
HfVXMzmNBznT1TTRskVUGyNlKGiGXJ3fLmVlZDXK+lywImDMb38sgdQ8ESjECzdA
bouGM7WkC8ccJHWpterdqx9TzNMHgppkC9aBCPyJ8omhepltxmRgA7E9OGtWQ3CW
Kr8RbvS2V6CRL06pHJkbewVZ2mQlTiXvLK6nQG2CS3aoh+UeGzWRKKIvEUPi7Eqj
4/APVkn5vbshGH3WMMr5yqo6X99JG1+wP0AITYneGrpXRaVZFrG+KpbQbMKsTUoJ
tADdwFYOLn7i+NjQV3GpwzW10gK1zL1W17MXOlvNbomXGei2pkdi7mJa9w7GQjba
yNuaXBsJ0MH8gnquVq+UKLk4vkudbrTbfbDAsx+LRPfIlBpQYjplC4dwdN6arTYz
IrM80LOJroKjcHO/5/yY3zeHKLCG25UigXmja54GWFCRjJ3PP/HPQIoThGTVYKPl
wGGERrg6SHoLHoy1sJ6jGSiHJXJmNEIj8hJizf1IH7LZECbcAG4jeZA07lw5vup1
Q4HQ6AHhfQnaql5UWtQqHZ0aNUbZyXUVllikAmmGLLpnEb41qwooPJ6Fx+/P2AFK
CunXO+irfE6dcTkRWcjPoUR0xiNeLDWPTIS4XGzPuxArkbVPCnUyKBJWDf+Yq/sT
ku0zbni8I02igNT2/WiIRVDOENzsCwUqjNcUUtAYUPRefyKlrnPF2pdqfgcobnW8
TVKN6UgGSbCh8yIl+I+kcFRFgK0Ln/9poMfpZX5CVkE6fuTz0clZTDTHHRVaLa+s
g3T7mrLLMvlmwi2WYP1wGhh5NC29T52FFR+3qsyMADz9f+dtSV2LOuvePG/OoEv5
oj3Zoci2P511tEcByxkzPF5FtdPo2lqZ/WSW7IjVsdoMO5WCDEW4ArsWXCKEkwOS
VufP3kmlutLxsHtkNihBGDmfa50bL9ZIucafg4uGYFf6jz0zh9fG7NZdSdyq2fzZ
+OZGkSQbAfMxDDEJba1j+Ef2gOmv0Jg+7Am24ik0Aa93GfgKPDZDBJOtuZUngR8A
1DHq25byfWcOrEZuf2DCotSuVkwRv7FK0McOSYZWJ8cOAo+I+wSsnm+Ou3voah96
/pZoIoyCITlv2xDHCK/g5Skn/c5ukX4ll4UH5waLeulYLQT5CkFxYB75F2yQEhPh
wOUo7KSReA1e23aI0M8oqiyCiEa6C1SYDY5IIRkV7jQo8+gd4vIAHYiYHBW21g9o
TpULw7fhijzw2Mfst0r/AevnPFk4wMpPBJ4nFlfQGbjnGHCDIfEIF3Ueks9IE4sw
rwC8I6jHSNLzAYLK9W4GYMSr8SoNP7xX+gZZoiyJqg09NB2d1RNGmtKBkW0GXlJ6
/HbINb29oOjKfXe/HmBLoWJxuuq8+B38gLGyWZpfdc0Gyx9AiSvzkXybTQcAS45i
dpPciJadqDkG09s8LInC1WQEHMQ3XpElp7QskcqA2xw6NezHrF1wM5YTMUe1BXCU
mDEx9YxuZb2UpPLWRkPM1TdycbTftEenKQe0BHi1K5loTBc+lreBgtIgJWH0QYt5
TlXiHqW15nSRnpDRXShvq8P2uH1dbN3W76iKFQ3C+2t8Up8/RXhlSempQr55VhhV
fd32ozPswYUstDg9WLutnkUr+VWvAVqyj7oULLLiu7nxy6izxScfxutgTs1yRfZr
txFZbI+mWJhChdufagfhJAxjdABCTR+sb0nk99mK38DcmOfzv48F+rSWUAe6giVB
xiDU9rn6LJzW4zU3BtNapVuLOxZw4CEE97BmtGfe8P97DXQGOEFCFa5agHummx6x
mDUHd9JfpIFMPupxnx7HE9gwUcJWtHyTjN+PiVHp2HKoyEXxbUmz7CuxlRIxnDgV
wYg0GkhjGZPwau0v3pESIMtqsHgeg+IGrylm8kV1H6Km1mYUn72hKH8H6JsaJ7GW
4HP3JW7tjenOFAXh0WZKuD8oAoUY2D7JWABR9L9Qw6k602W/eQwDuEb6FIELcWuS
4Whk3/3zGwj+GSWsIUHccqoxdwkysMwkMl8QTwPD8xVTHZissSRY8X6ziGM49kly
NXRrVt3Z/PmemL3e2hcrinINb+5D8nEON22beBHyDpBZuTirDfnnJgwU3Mc5ZR0G
rk6wf8W+Pb5YQTzIgc2Q8L+krknalfKxVsPzO7r+tpiZWkwHoceSzIr1koSNo5UM
p3NF3juIUu1jSKoxLA98zglcrV2tlIcLTzINV6FOFWBC46fF81mfzzrvFVCIBceg
wa3wztb73UwsdpAR715HjXT//zcYiH5JlwE0WIZ4n2rGQ5xKT95oPjcPc+l8ndn+
KfbME4orNfsxE1AgnKdOjR5da8pA6sntzDSMAiOIjag30+sSQ1QLeJVQTn1Jr8ti
Pmt4z7GqetQ3xNTQ/g57ftiFO55L3RS42zWAwSH6htAmHQWwAFvlBF4fHSRa2Ezw
Tdkta6rA7U8FsNsHpMikxgdlrrm7gnMVGl7IYVY0CHzvTLDzGggQMbNjffMD/Kyj
8K0huB3+cAUdGjL38fLPmfpsTJPS0ygsji8Wpt+7kwa755/vB9uQj1q1Z/X7ZwRq
ei49hVPi/qH5IlydB574J1McQZkaCm1Egq7q0fA0BCFjrahI4xGOzZKGr9RDjC67
Rb6jyoc4jQV7g3mXIC7hxCSzF+XpeGceUimCtUwhc9KXQ8n0F7n1C8vRH2bn/HIW
7OvovgxvgOUKIaJAaj08JmVnCCJWMNzuqhiOu6eeOXedh0iao8zQryOIOQy/Oj02
oQc0bG+xjkuL3ZLS58tYSI3ctHw5da/Y8NocsWFR+Bbxv1qtlbuoH7lbEMV00zYP
xx3OdU+R/6axRCv8oumb9WQZKwD+hjBDfwYnWs7FPRNUyVUGfDhdPmBozTLTcI4O
e4SNrbw9NohxM4/NIlKrWCQ8BkeHJYH02JXjx+SqGbK9dlVXVxOYpe2zvGrVapSN
S6ZE5nGzV2fO4teGrG4Or/nWS9laJ6D5tQHZLGiVecTR4cV6c8EUYIpmspb8qjDL
xDAV5x/r+3bKhWU/pMcSwpGXLdoraBWdXNfT7Fk4QLNAt2S/+uD94BLNC5fbdD/n
gQMIe1A2dY2jdsIG6e6hQ39/Pd8YTCbqfSzEH2ambcnnq5A9RYS/yof7IIjM/oC+
/duvi7HxwE7o/obSm1IcEH28xb3lcBcf/ZvsfY2Mfeql0Sk9KQ2rk/oOQZJj6NTT
jm93V2JDcgx40DISNbEs3sDak8AdO7iv1M6Dc/z8fto0ecK6+9JxvbKXftlOAXgX
+ylb6/B69AwAbYykw9JfbgyH95BKXqc1zVvgcRKHVIZHA3FBGHP4KZdNSOcErjN6
5n4MqN2vE7cFrDeYTj2X8NUX5QCJmlYIzd/832bGdUNUZV/pMU9VFY312fgGFugy
iCmsnZ3irs90+zdxtvW6HQrJh5eNOpfCaiqSPEdE6a3mFKu8w3dc99RzCgoGyZ5N
H5v7if0FsxngRUpvInIVwznFPhJb23ohbxPgU+AfJ5+JBpStFoA4PI/PcFzZsh4m
PuoE5QdKlbZ4yI0eBx7ZwauRb6BKFBDYybtBbWUtvk+f1iOz7WkzCt4RIB64ysc0
P21KqDDSzDsexi95jTGiyCYB9fc/XyqAIOYjO7J/CkxmVy9XHG8b3ku4peCTekEC
A9AdBtuAXKjEXbcbeu4Be4Yyjyq3FJvo83HkUbg+Fx3Jv0II7JuJFQq5sbtn4bID
YZJoXolTmBZyu8H3NAwhsIS9BiSeTPS4GYTWL9qQXoI76y9tSkGOhwK50zMvtNcK
jypRyinyI9OqN8z30DBD3suENLc1uD9OY+SeWqXPTijHEy7PycOxY5uqA1urJPyr
kf0jbkP9X8BiwwqgStYfVtabf0BPpXHXB8Zi5kW9HyUHSvx0kQtsgiQujBk5TLv4
zgF9u7mQJ3q/9oKXGYG/tyfnhsCxQMz1l+TlOMESsbvuAzF++OJWOUGUzx6m7EXU
eB09qMx/5M5aMVA/RRoV7paAHYbSU5WR5N/LZ1jjED2S561O2sgZHuGG/EVUA8bq
AnOmmMZxXYSDm89KLa53DuXukjwL1SuABrYHHzoPIBtJYXCIn5Arh++04cAIK9iQ
LH7zFNelZqugrhy0BVtpYm1IDn7v7+iec0Ui6p+/nGK7r3ELcQbXa3tZVv780HOS
mGChFFxeCYcPRXjTZvZF6XtOicbCF3Y75XXJk13gj/0zscW7E1XDHs0OtFJ4keab
H2xp+JJrxg3BTtRC7Y/AUxGPmZISF2T/vq+pBlesHcBpH3tMNKrLNPPYhgcuZqxh
0mWZfwKzIQepmfQlK8ZAGXHocEQHdOk6nIPGKhokFe8Uf2FVhku4XDr/q1eWKWoY
DsPoMytmRuvxPB0MQXevMFLcAQRClqfOWdIFF6I4bZVyXNfRkiQZlgr1/z+FQHbc
gULHD6Fzxdencj68+XDk3z2J3vv0TlTF6G+Fc3kTSKIch0Yntq48yB7kzzGy11H6
wsalf2Vx4fdsCRx+FMDOAKuFFXUeWG/YJJms5Q526vHNBxxELkFAExnJI7ceT4w6
qN5WygIBtXRtbre/AqwGTmPU5UhpVOxyvZQEFtSB+Ey12XfX4pSgcLaQqgz0mGYd
3JjDqXpTVzDR2J9xoZ6DqxOu0pXXUMQDpdzIXVVkpQYLU6gXDczwkVTTe/8ulnRm
2A2ND5f/1lo9nfJjFamppusdZN9zaZhhOTjEiAgnAiHB0DF+qjEbW28PxaLXHKwf
h9GWdVWPx7NeZEHbzY9gK+eIW8YMxra86rSV0uLkgCmvlzNyDk7jd2sa0MXsl4pn
SxL+qY9PN7/AfRmFEUR4gmPj5lqNacjFpfawzVcOfTUD7LfkCdEny2TyWjVmppI/
EhPWPVKYkL+OHvbBDsRdNxXfluap3lPsXVe97ny1f+ZojDaJeu70LCXB+beRgbKa
XbdfezlWOk2FuodWPe4/ed26lN690YWwHcbDErVVPbCgpJ3Z/wJqLgAD+GQY2x/K
W9Lh7maxfDY0OCJuD5yybIJoerA2Vt+B4Bk11pYQwRfj//ARWVjT4yGU3JwIGO3W
/J2MgFVxsC8UP2gMqwJBLPHsr4zY0O4L9P4Rkwg4NkpFqkatc3qlyOQzhbauL5Cu
8RU1qS3E79BcJY+S8j0FkM0WbF3QIx7I2+uAf34LmwhUiu7/ETyzIJ8SzAl3ukZ5
D8TKkXtduZRn3RFnR9FCdKFYpRddQHVXphkQq0BupsX3iE0S/bCJnnFyXLFyy0Je
qn9ZvLlFTe7uYaexMopg3CLcDwseWipWxCknG0kXGldjEC61PLtIlJocxivT7WfI
V0R0bk1uOTM9Z86FfweFpvQMG+2dTqGSTbqGLVO6ECu6dHwq1e9mWAzfi6DXg6lz
FrzG6YhCK64p1HvnT8u5HHOn1hWFjw6t349nfgxGSpXGxfSNiCYzxJ7EiqjsM2oR
VDwSJXMo/8A2kdg+uY31G+tqJPlbxyLRMx/HYp/bdrT7pgMiGbJfXIJ4gELhm7Z4
hinNFv3wDtTnAktSIdzACpKddlwWp23/KG0MJw3TEkYqmn3Vw7jmfeB2XJ13qjRD
qht+HPnApQrx9DvDImG4eGsNICpsmY4bDigmZ9hwmt+wPUERXV2i3RqfRcWSYnt2
qv9XrYwp91HUbyvVLhxzgKdAJ6NKUAXuYni0W1JTp+GwESQNtUfEcXWds9MH2fEr
Zszmr2+OFvI7F8rdDWgjDv1s+vovXHSB5x/muIdoPQbdl6xlrAfELLUtV50cWVdZ
6CjWkFGnJWX+gtOjHuwIf4C65swkv0IDXrkkwy2R4lsifJpmPPHTWP1hXmDf/0Ou
g7OgtQU/ZVBwSZTrCpq4C0mXbt6dlRAndf2nOX65NXuZ3ZMqQZDguZJY1YtHJyQC
Fer05TXkgkcAc1lDkJLiA6EWCQTqStHOFBr3c9S34zBCeygednNEesiFPPqAAY8z
JXgvGydyZChdMQ6lZwFVItwcgKO/P22zDIpeKD255Lhe5dTXNuQGSKcpWc8h3uG9
Kv8CQqSHRXUnicBCKe5PJZUWmQ+zp6ummtV5zXijHZduwpy3ACqdvLhK/xc8pn2r
EMqWGg4WzfYNJWw4bHUGA0y6vrqVq+/MhF/LVui3JwreyEYVl8GaDKCWl7UV0o/j
GFuA9TUP5Z1XClZeEoEnt5cHf/JdgKET9ciPA5iihFsTI6pB1yNfkGgTx9XUVbjF
7Yo77MDS0qoJ1KbEPQ9CRCSwAirktftpHPiXU7HWF+QbzpNtrtgfnye3D+36E7W5
y9gZmO4JzjlYHeKwBGFDlnQXqrF9AOpgsh4Tuuc7aY9OI9CnVa8r7sxtp+rnYAvP
NnV77VChPos4Xpv6qYuy6XoH0l0DAxjnuRXASxo6Y/4GqY4FqzzDujhOaA+Y2HTR
UVQi6GacjWi19Je0fo8mVHAkPePMR+AhccgV9g62/Gtj8n8yic2dR12IXu3g8SvR
qlghN/RRZYl0iYxJkHTL+bvQ/TFCyd5b4Uq3V5p9XhlxfbhZrLSLvItd4tz4tqUf
F0e0iunCQKR6LRxvG3Y/eKCCw/Lz37VXB8oX/MRFFfNiGVUzpHIPfAtO7XvHlECR
Sq0cvdRPJEVg17sL/EZTr8aJbXpPAJEIS4ZXUsvloK+nhe6Gw9aaTABP6vyg4LX8
btBntUHN2PqZnxkZyX5TJn/Ed/6wB4vrzIivPA4j0O+cD+7iBV59+MoQEcSvLfOh
ee+Oj1+hqvlUBsRqbnqrbLpcZtmDXP68CQtvmXHMPtsrJe5slVPll1i2tBw0en6m
iBxUiK8IZfjshHREbcG/iwStlWmmNHvizE2Tx+DkLap64NwywoMETVWeVcaS2jUT
IOkJCPDyKQj+q65+ckdXiFCxm9fLXfljAs0n0s7XMT8w02tMSTGF+dfNxfXuNxqw
9plH21f9cB0TiDOcK+ysGaQKgoiMkLi0vWmA3fOPNUbBW2tppQbJwW3LAn+x5Y+N
yr5v4gnm4baKaXuVGOgrQNidJ9toNxi2am+Xw2NQLJleldssWcDWiqhNjk56G3Bn
XUBEv1JlPLkhLB+tgXEmVRx2z6Bry1ZHEqdhngkXVr+30ls/s9zl48SEHt+oxCtI
rKdnPzYB1eqTtXGezrE4ui+VADxw1bUklVfEUhnDG7Q/ICCDlkC45diKGbi6PAD2
0lM9k//EyqcNTrdsWPZhIXDXa4PCkF6UuGx76TX4/7aEm+qsh7hXI6bYxyE4l23L
I5drqITnvTrWQiRrzdhPqhZyXJKSHaVTxa5halT9fh7352U0jlf9+R1RkN0g9hCj
6g6LOYk592zTe3fmysjq+0zz0F9+Hnx+Y9M4nYxs5pPxrxs0Ylr9A/oZwHbsXvHY
3TIPSsWglBeCbeKnhcZecE4sh6ejWHc4mIe4dngNSHWmB1utFwIAqM7r3r5/ugtb
Cn1QaolLVQ41xkjbkqM60JeGAev9qTrIyOWpdkYtzdN0b1kYBb1SrTAomSEh1MIG
W8mt98ZhLHy68D4IC2PN+xcspydETOuEE7pf6P4Y4jEmYF2UBzwQCXYAiJxXuAcu
bd2p1T1Z7gUII2rvjKxKu+zrGdvygCKVMcJ//MNSYNa9yBjPMOvJom45CuOhhvWH
eO847C0bbBuR+FJVwl1UQWyujYx2IM1adRGD3rBOLQ5nHdgX+zcbq5DAlhhBlKPU
8Nq/q+RSgYYni+SslXI5C3gG+lRXhqdsw2yKO68eAfs8GRjZzir1eWxyq3mbhWiE
BWcMxqVdkMvGjOxQ9ScnJMODh5rEBlrnjkXPoCqLxmN0VwzCEoMLrcHEsd6PxSJw
kuFJgb84Vl7XonDap+fGqSqliwkwE7vzdBGM1D7CH2KCEkeM3gylV4GbUCdA93qg
XNEkGt9vADydYGn5dsXO7M7LsW7jiXiYfJ9yKXy8tL4nikZupCJ95gV9DBei9Dr+
hVgDvrLgHpQjM13iuZ2q/HZqN6hgRweeJsMpxydyYZykveFJtkX3aLn3GUIrhSDz
ttbu7J0BjY1mLawrqZoeeX/EKvih5ekXZ9Qy3/vZPE8vC/JIjN7MvUywErjsXjIG
+jDJ8MiZB1xyFPC/lg9hmhiX4uqULQk0sU+PUWHLb9+X5L7DCWMxeFYLcWf3l4/K
U26JX4kIP2mI0MkCAXKarwrUvVJIcpVSLfhYNPnZ6wb3nfK7DaKVmnOc+IvTop0F
RmSKmeJaWuihzw2NZSVDtwfkFqDNyKyQC2S14pP2wRNTU2HoKAPV0JMs34SOGPih
VdXz8PVV0srRDWMZDgAqqMhVnoxbHYgrUMGiJnTWTNBgAVhEo0uHvtfIpYRH0xyu
cN05qD/Cm70c5orZ8sozHatqxTokoCCzK6ZmewziTIIIthiuQSxLl0JyFcuopJBn
PsSP9Ghog+ujIOcsqs9q3kJXYBNFiVN+IffFAQsC4yw7VePM7h8wotLfMM9GLMhm
xbPyFdpsIOu58RjWR/ufpg8poSGPqqZcGEA4d2kvvul6BbGc7fU8HIsJR8mYWIvu
tzOTZU/w5c6AckL1g7tjxkHRyquwni5FmipGAiIfJRVepOec0eCC3D29chQxzhn/
XvljccpC88yrvpIY88ylJavCxMjMjbOzufi0KVRP7vtiVH5ROBWIKn78ZnH56xSL
xMc2rwG0h+eeqU+oYOPas9NDF7nPlPayuKWG7kMVGHVCfYcpvqhRtkPus8xKBxi9
gW9o+iati9WQMAcgaa1TIzmZwMpPGgRm+vSEtL5mQbIJJRTifMVFqXPXqWdcPCTl
nclYWw+V6tfviDiCBGG+v4NMIECwQbT8++9Yf2eDvCuwm5QTq/om4s1Tm7WDtC8H
So5/KMhHX0WksaqEvczpL5RJWoGfSqYXXq+OUj+wrMjIA/NISBM+KPwx9AnzhF8F
qJbX5nujZe5AxwVpBGuZyCzCi29RwgXbZPm4IuXEDtft5/R4OPV9K8JDVnukMj22
xQzaYvQsP9zkj3/84+lawT6ThJRTw7O3kxG1lsa3/pGkGT4K7FqIPhWQg8AXYDGU
tga/2mj+Hs2ZGjIk2tsbbcSvsaTvJ+YsmpTL9eVuhErmmUzf4P+hB/Q7fvG0XHh/
5a0M9tzpdWTLr/Nx4lRnYDRtlneprMemLDqk4s13SfSYrJaVSoueYavp+DjRChjI
5D3fSBwG3aehcswaCmeKKbQ1DndUNKebZPu+5em7SYN+RiHo5R7mx1HOxwSVakky
pO/o42i8A5ZI+reLqOgZ7am3JfjZPisblZDaEPLfMKx39FnBzPr0lc/rXSpP4tnH
j2agWw4k9QH92nMv4JKZbVd94Rc9AH0M1f90n/+VPZxcjqpJrmkvQqJUaf7Ljp5J
8+qpo/y7Y9K+xHz0AZMBCrUCye9uvDMYcLnMnnDzGgNXkRSbHgiQK+9WuI1lL1sz
Kolc3Dr6tRkU7P3HNV7615ljLBE9Y0VTcBjZnBvddQDPw9NO6u2+4x3Tsb/LX+Rd
F0uBgwl9c6rhCeZ12VAWwZ3OaO29PjlS3Z6u3J9rUy6MVd3xFQ/CtDjG/uOhDkXC
J+ZIzv8BQNy4axo+JYW+QXJv2eWW9jXMqqZ3eIshVneQ5RMrZslafhwHvnaOtBlE
6TGJfKW54PGgT+8NsvM7wO3M9pomXpN10f7Y/S7vk/lUFuVJqbwq9/ismF5Bdqfj
RAB+wo5KnIaVCgEF1IL1kVwnREAICfWqZw8wXCBmXLPaKr54P+u2j7dZHo3wtGzG
UPS/CDCjlj/gwBwB+UhMkvuqa9AZWyyE380ReEIcAk0Cq7mj4GRpqx/Dr7643wgG
z958xVWU/ATQaG98qaadKWlNAiuZVySUC6sspe232DvGbb9J3F2fmKpn5PNBfBBx
BMCZOE9+2ElCiWExeAHgcVhxdj5IxT/wMgGrnFte9nhPP/J4/V71SkAqhfVtdByo
NQvQSI9YkfreCH2joOcWf/ePwtOeh0uBFAYBZWZEtIJEqoUnZMtko+K90NUbf1Wq
b8uDsK73SOeLhrTdJPpYOvUdUiRbap11NX+AAauoprli8X5yHmeePiqyVoSH+1Pz
O/ReHfgixsezzpEEZHpPa0R0tq69UoXLFghlb4wF0eLeEZCL79VBgnsTn3CESXp9
f71W/z3Fx5Xy8HiFTmZKRByOrFhM9P6+gi8JJVGzUeeT9GCRvAZT37r5wYnEQL6q
AaJ/zHq+16odQ1qT45i0Qbt/7tDqrShlD0rrx/lze1rST+PL0wTK56hG+s0mbVhI
0yD99dmIkEImL3s4kpiUqWXCE7iiv86Md9vUq67uOD8l687o9O6N6M8//ERN6XnG
L8uySLMKrf/GZj4Lvu4qGLCG4MI7caTXcG/R0CeYIqLK4RDl3GBtl2JJOwiWh4iz
aqMRe0faDKOvgytReAvbIbI+XTr4Y6+CDuBRrREyDOJtvTxHrpNRYTl9ZNjLliKN
Exd1fRirUS3XXfxzCORYhfxZxdYDX3mrcCXdzsRApGgVsfEtuG034Jo7wqOat3ys
dYtMiRA907oRptnv3DNRXQE8My5i8d3NUc5SBNFek0Bm0CEC58VKPEmuRb6HlRJk
Gan04xQ90RwVDuQx1/UOeDj2rMUuFf21PrFUEmKdCABs/xc2oxkPms8mAXO9u8HM
7y6GNSeLVphNWbIwi05JrAa+Yrfmd2GeKHpDl4NxYCFWFCrpI/TABYSOil82oZ8e
vNsmdSjetFI2/ubpNojYlKrqYUbqwG+yhRQFPEWOt6KtF5/imZAv9Qika4Rkbh/X
wcJnAoLZBSPICm1NQ4lQrlkSw070dc6kfKePqxXymeySi0gCC0F/cWI7bqUWoNOY
xD4UUjNexEnaZhVhX6iKkA2Pk+TSjTDlg2OXt3CuAGR2MqidB2spaQssaLh9gnDp
AkBUUQEjgZ3VgJ5NzF0NoWFt+d6FhYhlQbJhq4zfkYJdlpvLdMbFmj+kKUCIlewG
d31lx+AG1uaiwcwTzlF+CtfVxdK2+dRddhZpF4CfUAFBXOCuXoR+UtH3aSh1G16M
306ZZWqIc2VntIE98mWOhOpGoZzAnd9vzfYsCR8+Ii8XhPtGnj1ICFn+QOby1yum
UaBbiFTEd627J2jYwlfaUMGci6tHVt4wxyILMXEmPmeZYuPH1sfToMEwD/x8ENwH
l/cQYuviWvmA5hBL1LzK9ZHux/lCVGfMKh+RNuN47dEEwrOh7azJW12913/fF8ov
qWaa0aq3PBWTRhCXeCsgrvRomcQ/1xWynIKNIfIFOGJV1MmHkxjYkG4/xZQODQdI
Dcb5R60xIqgHCF0h1JI0TG7WoxaM7hq6YGWOFhgnSqB8pnLlNjsALlhOp7g16rcC
wFNPv/vBUP5myG5u76Tz/bHRBA6ZyTsk6o5yz/Pl2JDZltN6rvhtZh7TVNhNWEst
+DaberLQHKoWkSPFMwc3Vr1Hz/eRFSFO8VZXPS1776GZOaWuCjkcOjYr46aEQgyQ
SNEbHLuee+ZHgM5eTexEcZdTrBhgBAYh+v/9jDMl7iqlFq/zN83o6r/b2ZCDx27J
dCvbDDIHTSTb6yFhtYHQ1Sz6Mpqnw4OD+n3z9qk1ApQotj61/l/gQfSCN006vjte
kXzaiMGXTzE2Aqm53qoqtajmqYSQj0kOH1P9AcYyJ2U+ZWIfKRZHqMavJMxgSBVz
H0jvAsC57dX/kJdvftYmu8G1+9rZzbMcc67NfYMxwDXmPrvq5loRtV79hasZRQ2y
qORZfHiEvqW02xA8bJwpTI8lstjjlybGKMyu5GhT52RchBsFu0ZzCHQnm3wPT48Q
Wo6VzgViEufHGKaorW+kGeaLhEp7M69sU/9p6dxKWeoU+a2gQii/zNS4gCpk3LGB
5J4yu78zcnA/nGp9/FppLaYGnaLt+nV+dO+hP8fnMkuUnTXpi0O0QYk20GQPJcBt
4O0zV9uMlC6MLY2hAWi4PGZ82ScwAPVEUiHeN8U7Cn3ZVV9Vh7FYzZAARYT19QQ2
Vmd+TfgzMzwF3pHQsEG7CFtGIx3Yd1UfC/5iBfmCJnoNP9keTsNaqdu/2Wuw2dJk
ZG2YHWA/oV1SMRXIGGbq3MApGysp/Eaj5jVyfS00QpG3QY7KRvyBiyU8esBbHo2s
1LFj1Mzzq/PhNLAj3iVKGrTWQYgaMAcugEDxORj41epeawHuI0A/z+aN/Nhe0HK2
R8MR0m+ps6mthYe49vJF8IljB8l1J1Uy4Bfy8F2hXpmzFJYnEx2KaSuu8mFCP6YX
+dU2Z2RATk/2aaVYjVIPfM6LvMYwbNoJrzd/GpjKh19t0wu7DAqsr8ziZ2dFqJD1
2Jh2+umQ9/elm4suCYbXPcgjsPTCHoYI6jVIPR1csAnMrFIF7hzUpcJZbhfRySt/
hkyZasTGtbO2bz30w2h2NcFoN4hoq9E2iXWbYitrIjSkLUCF65jkActmhFRNLe0B
mN8wW+7xY4vXAdBbji7xxvBLYxwYDIYejZ3+OTS9QF7+RhzSr7h6XXXQ6XrNUxEY
Aff5NYSkG/FuaiTJ04ZCmelrHPGKN/o3jKPmSdYK4DcxfhbOovojNAX+0CuON1HX
sJ6Mbwdvjx3Q0Xcc3nH/65+tOT3D8XywH/zRBqvW3ijiFAgucBKf0COMX3DmnguI
lzqZksN8ymgZ4LRlnQpL9YBCD6osjzapPIthNiIRh/uCRYwJWuUlqXtAYAcqwlun
wT8MticBZg2Vle8MjbQyWKTx4NHc3EqV8GDJBNNDKCkreCpUW/903WPNR56U5Fg5
RGekAV0zLZifwZ7ZhcZi9nJWHmTZThpMDnQMYaI57nGoU6HAzYA/NWHAbmjdNCir
C5DHln1muhEwsOOZ/qYcZ9ztz7f5Z+vHMvFyaMgbc2oS4cSRGGqx9alFMBvpGPwU
iuIwnhr8AVMeVUtdju8omz75oMgkruYjbHohNaRFhNTxS9zrSBD24rODb2JNA3b9
H0gnDINsjYLfIvIh1lmzTPMpZjABq5qBErnnlRe+p+gZpxiMjS6FuJ4EvafPy4em
o3+qUnasKHxd0JhsqXZQaNRgxZgEMTGXoNQ0ffWgYyhV9oOXsYXwnWHybgzMPb6v
gBWBm9LseE/uTp7+XoIuiKEwgDlFJP25rSgKjSswqA3kM6pwSg0f3OvN9Hv3h1hl
o5sQw60eg8rC1qlwt4vz36kkNPOHdP9mmrm9RIM0vCjLt2q9SI+np4ONAQC+/EdB
G3L11Ju2DNYKBRTNo0aczedaEsR5RqVqNSlqysF4oQs0EO81Q+NLvR2ZXhGjWiPj
HIOm3zIUjstmizc7FfNIRb15KHC+9XDd3bLkesq8sk0I8ezwyqlpPNioXxUh5BMZ
bzlnpj9AfljS0RZN3HRtK0t3k9MLX/V2F9qx8V9BHrf2QIOOKcO75SmKiurgsmtf
qfbIeICAnOQDKjsXJHpZ1OFcV443P8NfVmXCL37BMENSG5WZGKcp4CYC00sLMVwl
oSklHEJ04H59MBl41LRoWFWgI9ERHtV8x0YE5Mj9BRDiG9ashgt0Qno/fT3g+aOf
EC6Os6v66gon5Z18HJNvdwl79ylL3BxxN+V1mDYTgGdyiqnGDB3CYPKoEQmYF6YW
pahBniMWXqeshkfbIOwzfjDq1INuYg8GJHEEnmv+DgrY79tQ4RzY0N1VymI+K6b7
5TvunYrTkMpzbj40VOm80fcGLaKuHfEhuW62wYSGJh5DQOQiQOKSX9J4Xgr1JI9R
3mik9gJ7Vhg4r8irbNEiitv/rRkqU3qfaUJoxgIecFwqYo0oBC2IDlMzCSfAM/tb
ao6G/HNy7eK3KjgIAKcsE9athHuHTAl3EYEm85eeOYuVtviBLS/0TIgcu6uKw3d+
wUiA/EdExM9hvD7n7hhNBjd+5Wa71dUTZ2Yg6XVQDhTaR3pgvFADeFA0qZQjrWFq
tcJ01O6JFUwVrmRs+lDbU5/9o75WA/vRAlJ/UwUBPkgZsgVEntgi/96IHr+zKyDL
cbGEiMb9sahMbbusE1+Pc6ZeNR6Cxg73ISrn7bTAGb/ZyqJb5/PtUWQxM2PPmCIk
jUBUNaFwHGB3ARBdf3SbezeK80N8nazNdDAZmu60zZoRrCYg0I2/LWOv9ghJWMK0
GAy5/d0IeEqPXlsw+7BYWGI03PRAHI77lx6UEva6HZD280yo9REdtXrZSm/ga96C
x2tWqHEaZErtPTeIw9jE9z1BjHPG5d4uO2DyafZ8+M0iW8j/zgM5P+el7H8o6lY3
bs8f1/qmpTcf1swkZB4xuRoshU/QrSMpHMGB0VvzYmQYwvZPRrBG6aYRI0QDPjTt
aog2rqcxUBgH6UO5+Ki2HG8bz7+Lzr7hGkqu5hYJ30wWoHUaMW25wljJiVwZVNho
Y9VTLw3Cj+arvMW1JsiKW8Dy9m+LDjDTcTNyG4COkbsyVbwlwwClsUpQHRsZsASp
UfXmzConcUUbtIplomWIXWK1nyygNWVUH8W398k1cMfzwD9GDBdSocm6Yo27vBPz
Ulqr5ebJiQY6ZgJrYetGx8aw8keoC2uTbMqwfuWUX1srBqn+7HhgLp/dRjMBRPbR
HHtalHDcb0g7yt2OR0/mLhCRHfNq6Tu2+arhDW89pdUbkuncHau+lYwmGUKyIaBd
aLQhPcHV1PVarpmUYX5zDhvHvqkl76dc4wMFowY0HDZWQkdP2F6z2zPW3CatP0rV
ltB0LnsvD1Yl1fFUcH31Qs5A4mx4t6X0uos+omLWgCOx1wiN19K2ZxI8LenR48RL
GT4OIFGksNFH9gCSxWIlA2myUgLvfzAD5+3JeujdSOoDggPbEwXtzptVBxWxaRhL
T09Uy7GERZlxWcF4dLwqrwd3ldJxN9IyzR4b7nf96+CtEQzo+D84YTSFtvdcKAV8
cCP7yIDEEzNbXO1m4ocdfWiayqQmMB0b4vdn5WBjl38Ub/W1xZ+zN+8QYIsmT0nO
Licl3328r6thK0dgckmAeIYzUaSBTs2DkNDYjFR21T8QOUvJ/tzAlusrFBatVmYs
WrH0alo0cJsAJuElGbUB5K6vtUErdvbHIYk/9Lu6lRCbepi7dMoHRpkEZVCCBc/d
VZ3vPp+GlsX2lLKxgoVUHsURMYRVVSwdtdL7iDTWmgVobByeyLO1glYiXzoqf4IG
fiSi0Tt6100FDvpJlvNmMA/R7lvYXpfj5HGy+aeyw/xpAAtIzGyy2sJV2IV0ol62
1lEf5snNWNfViEBE0cRDbTlFa2EvsHSWq8elArlgloBOOUQatF0lf/+qKx5aIU4v
6Z3oF3w/QucgtRnDInlmsdRKJ0uTOgcuv6Tl/zw4k3to40jMJWIlps+j5pBgWQ9a
HYXOcHtAIl/aclPGSNQ7snv+mh/1OYyQIDUzDmMLzinS1Sgt6b4BKi53kah0ICV7
qe0FenyIlUEfA3IyTBhxaBpb5e+/Opycf5kCXpixjSx40VAYgzohTlIRhQgXNZ0m
jiYUI4TMk5gqgjwgsL3/iiUYFAt18Y33ed/t/Gj36+cexR6jJiNfj7AtCBw/7a/7
GqAQ2y2Hm1cR94IvPzJCGclpHZvsqvVVX5CoqQvGf79krd2e3g3Blrjvsxqu8ox2
iKLiHZmhP3hg9WeiTYpkToFN6VVJDb/KgBZb17uG7ouDSLNGUhcFMYaW9lekROQw
Pd5AtDkOIKdGEbgtepBnPmNul7KWxpQg5hqmwEB6r7bcuCQZwda2qIEsy5dVVoDJ
KQnpaDb9xy7HH56YI+pgmm7T0/j9ppC6NulcoWRtHAdn9k3T0Ci2CLzoQTXOVI4t
TOziqlQstnPRkOU6cXTF1OuEG9tVQj5E/U+NNrZQF98B3neEDab3N1/FxAO6ZaC9
T+ag6F3zl00SltVRZXdPTsUMizHSWtB2aK0u7wDMtusUpi8S3XGdOVKPdN2R8Qya
uiteGnRZifs0oj9ndbJxosm8W761JBTTIzs868LLBpBg++uqzJdSmL5CSx4NItBm
HxcRaAAsy4RRKOvNjwj+X4yUUvgMHLtxj85mCe7rUQn/ra/nMcQiLIVlICkzingO
VdI4kZfXL9jhfDwR7bvO0H6z5nTKpDSe4uv73Pe4/nqkcXewFylgXQBm1QUx8wR6
/9oXMQLhkCLbxP/z9Mv2Rftk7Sk2kEMvr0Sf1CE4YxVK7ER3Rzo2JxX5SJym520n
8MbYQ79c3L2VhPYbddkIRnZF6LBZby8csIHm0sDkR/zkyArGJprq5VQlCiw8e1qJ
WsOLFPhkoWMea08Um7+sdZZaPg/NXXAEp+l7W96pO7qV+9PkvCYe876WKpSCftFB
PO3noYhsNqMmAFYvck6V9YkD6norKO0Jr9LfEfFAo37YIQeIVlEZFAaCzFOVgaqi
c73gDOeTp64WO3CylxH0nbHh0SqolU5BSY9tpeKsg25DEYiEZGL8phlBUWsZZK/p
mcVcakirZ2lejLgXNwc7NVB1okzvUQH8X729c+XvEFy8lcfK2o3isGuBVQo+tSed
xkkSo5nIiCSPaM/kZ21ZFWtUKvh0dzgTl48UucImb2LAhI4ha+E8GtlUqpVIb/70
4dRCj8wposQvO+hZfG5NvM4+81t37oUHzqYmp612mbri5DLfVzAHSns6oKp16Tbi
G58xcQcL0JJqWK8iuMFCqIBE1osnuGta9+pKnYgtZ/HxtDp+0iJqIhIf/UcpMf6C
W26k8d6NhWMrimfQ1ME4oGF5jy68VbXbFy+SMp54ty3h+hg+QZB+NDMVqP0NZkB9
kZ53P0N+dFrLqpG8jD5Z2ccpQ3zt6yFyincl6aGO1VONRKfqzoTBw77WHxCK6WIz
AEnm3o3vIl4AN1SRPcyeWBHRfweUiGBOPPHHpYLOC4Puf7XvpykA+fKqX3Fwd/N/
JBe2BGF9mtSG/VOGzf9NdwxMvA/NemKmi0an66NO8Z11ChuC5i90F+tw3tQu3WE8
vTmZTt2gsY5cOBXJ66wXTPQ83/zoKdhoKLdqEYod0jmq+Vc3Wks+BSRgwQG8aKFX
dVqGmt7ktSlMR+YXwDbAmYNI58XGwiDnAjQW3WVIHcVY8sz+CVdpO0MXVyyvR5lA
VPccK4cTf5Z3X6tJtc2czDl9lyaJJrl0SnpIdYs33LJQhZ5cSyB+GlFYf644awMj
4ch2r5rsftuwdfJQxvHWUxZOp4V8OhnRq/rKmfrxSL5w1zNGBjsW9+lyuef3eXHT
baQkJ0RGYSRHCNriRgBr+SM7lQffza958Ee1rYuZw6rYj4YFvm2p7Gm/2lOXAmU5
z+K0clhxGf4KwcBEk1iSsBzOAFXtCWWS7be0zqiL0+8Uh9lj0sOCzospRCfeFqTG
6rqZaBeyz/xDq2ZQa+Nf3MvwY6/pqkkv9RYhouhfHXbf0hxMvObWlqnvlga8T9W1
15c1U7OscYlk9Mik0IMDbTZhOwR2fGHydfTlHOZYtwsQ6bDoZBiYWUhJEX9nT46D
DVIhDa75AHBsyXI19gcGMuOjBfC7W1u+48Euc4VpvMImP3i/ycMfgNyvH41evHFj
G3oy9u9mnd44nvLZZBrK0ioZFH19VOkoQfr4Jr8P5z0E4vu8r1wrWVIFzjX7hFHQ
xUkU0PpeyggNWLFl1Fbrr7bJV3e0E3OEaNLtfnIhcSroTqyO04803PKiCloU8V5J
pK+eWsSsdTJMjKXb+1REvnVfGRZLrcIH1z6wj5r1OgEGAQGgmtnwxzWYq59xzF7J
bjH8+VJCaY0z11TsoRMAYuOm31eBv2ucU1FrgP619Z7sjDazl/tSXPeVweiVgjya
zv7OelZh455m2Fg0r++ko3nsF+6axn7YWRhfTVcALEon6fWEgOQm9/saaeY9Fr+j
H+CvPPWNHSm+buqhLbAYAYMN1uMb+wHEX7w1UA6BoHjrvvY0iKk7Jkn89kUPp/Yu
e4ltpfmHA341d783jj55bPHT2lGt3kB04lAecVQUwW1jOSDAn6xSSbrMnsMs0Npy
Nd7U2C9egHOSurjtkJg5c8fEetOHgUzd3S14vlXCW9wqLbZ9i11Q/C3Oy1qZ9CMT
Ww9HnCKWBPGk28icjj5b5zI0CE/575wEiOZLKM06I1xc150u8Rn/hc/9ziqP19aR
FI3WuMHkj+mqSpADuYldHXs/71qJpHGTT4xgKMctYJvEUOPkW55BfkPbPFwUfa77
fyiTMMusOR6iqkgd+2wCpaouvjbWI3zDUxZtx3MytIzB945UgcaRHjjXzMBlcMBp
5BPcTJBXj0eJdoam8Lw3Zh0eNLJEYxF15hL8iVqng8mE8t7v3PFhfgpLpQaaHAcE
J0JILlT8VEMB+Xnpa/EETzMAqK1HNJC9gOD/yygBRVwAinhwHk+pleHc26R2vriS
JYQVjkF2A5SzfRMs+HQwQ97l/p/HK8C24YcInP/V+C3eD1MTZ2kPiqSzcj7k0J1+
deIHrJgdVNHnQ0yXNQPYJp6SabN1VBm5kX9jbzRkrOurtIGM6pYifdexQPFxZYpy
RmC4ZSsJdEw+zxn0H8F2Vu/TekOTAsvfxvcOJcSsPw8lZqyjlpFTAPzFQGRSFPlc
vLAzldiNR0Y7Xby1S0Tn+1Bxn5q2BEVUHTJH/iDuifzNtbeuKQvUIUtBTxj6EZ/M
UsuXr5Lb8gcqhRJpAppRbFCWJvgvlYUdKz4ihtM0xyvyPm1ayXpkhESVu7nExeOi
OMJ8ohioFXlaZ/nBq74Tilmj2x3xeaWELTuEjss+gun5D+7+/2puCOaY/Croi7ex
nV8HL7nLhngAihTc3OLiE2HZK04zwdDps0mAyoUrwvMZr+feAtwq9tbfBNRDmAcY
8ONA7XPfuRTfKKoD63mTDREQXgJXT5OTI9JDe4ZBuse3bJP26wEJx2G47Pivvi6Y
s95uyXNK4laTa+mnqPJIsRLNMv6Pv35gKbgAXGdbUw7q6zQ1eoCVh23BoDAo7MHB
UnigqJssy/xcQNaVNMW/OJb8rJ5BFssKVc3FdaoGaLuLveFBkeVoDwY9qS8rbIjD
QKiTbu9Kkz3cI/Lt0R/lPVhJyI/itk4m+rU/6gBR+RpB0pD8zvOg6yW8iM6RIb7a
c7vNXQcuSh/23vA88vVfmiM15abeyvLuWQ+p24fWkwlOkbxvsksxqzOfvyVN7l4x
sj19ioSaimZS47hM4DR2a1SXnPJfwWhrMaADOsTh2km7dXIBHBQhYW6ZQaq/iAUs
T+FQuvHGXtt/PDgvP96awcrkWum6Y/zNhoBe2n7akiV/Xxrv9OiQtYQFbDUW+94O
CRGEUhj7X6QqS8B03VnDGxzXZLCrx+4S4MHBxb5iiKJnTWQz16YjMSnpc6/m0HpF
lat8vmse5u0v3nOd8bP8uBxINlPaCmGfTez5EBiPGrq6v1DIrTM4cyXxi1rZvGn1
pCPylGUU24YFGyBKS+zGkUJ44kfNJ3Ow5DZraf8cPaLXK1RNNJg0alrgvLh6xwjf
fBqUNlu4XsMzkfMUCotJg8pZ6NjjEP8r6QBSkrBTyHR4OSecL5oy07Q37zhZh6jE
IXEWfatjGYWD31uTNwc9WQwU3VRNYQKew0/hElVQ4xilCl78usaQovaQvmxeBdku
KInKLtwBzlcGFFDQa/RBqaQNSzPO6FOeBqfbWlCT9aVkPc5VGsT+dLDLpGrVcks3
//bVI6iLurweOV/t1YMXhDuhCTvd3zaKteKa7/NLkEcgUO9PzQZOlH6UpcL7UbmC
DDbutAWKhuoN4Ba47nPJn4owkoG4weTSZhfel3u+ycvJ5laL8zFZ4jm5jRJzsvI/
4yhNJyVxEgfttTsI+oq9yZCgy1MQfutSI7xILXZbLdpgYg/dDSVVbV0FTyKFB7cv
tWGfojSKQaf+wDC1FJl+gOVwUM2hz1kyKUhu/xeG3yXaTYXZo/7xppcoIHCwboZM
ivk92aJ62YwoA/dS5Y4imZ/eEFmcUBr8uGX8bN00PurPACa8D7Zrnoog1oVtx/dX
V8qMnhWgllsdBnxpVaPvAXH5P+3wKZeQznBhCqH3zzfJmlYr/tNUyW43+aZK0+6F
X5GtG5hz78ZaVRGEpa8iuKhsw06WpWNGwZc8ti7bWGNedcNnsiaXzasibhlVU23V
DRhNrYKluW9SgV6ErbP8oE269X9b5BhikHdGg0gVl7v2bhLuYdwlcqYeHEdD2vnt
Jb2sE6tSuYyrR8YWXHSGiEmta4aEQaKyKIgzIdhOO1UZQ8xB1Qy3Uq199+0Jvm2e
A+P58PKvt1tA+AFgiaioUOnJDASWTG+GoJbtqATKlEU1nVDo/n19kvWYQkSD33rJ
Cci86PAkpctPuHc/tEKc1+u8u2YBevUK27uXl1nO/NWv/HIPUpOji7fryPOKsq+Q
+q5tN26CE0noZcZjQ+7k1CkECx1XRu+1o2ey2qwWjqxLe05hmwfe5604jBt3jJEi
6nLsRWz46Kccm9bzl3sSaWR1Odx+do6p+0YJLNsYQcssNuzgDywtYvyxDTxfmfLO
sbx9w+ChtsBPfHw8vFuLUQryzdny0tpUTKQ/HuEiPDziFOuYgCtV6G70Eag203+R
7ofRXuscUwnAF9QF3qBjU4BAmRVY2MEURTcOSjkciUCglShNnNdiWVh686l9RtRU
2aB07G4glP7odLg6G1Yp6vt0LxJQPgXKeY6UoVV3nmQAwR8nBOj+j5yl/Yy60ldU
wrEafEPfmorbeJBWYr3g34L2SbGif62wLlBsAGppKCDQXVoxJ6pkC4TyFrOayN6f
Mvk3Keb+auGtY+C5S1IumYzN3vlZx2YecFTbQeJc6Z52g/i03rBJz5hcUQe4aDAU
PVdvQn49ALEE2R+UW6eRpLjt9/pJQmm1B+B+og/pLNGqjrLBTR0JIZx34sGxj+6f
uV9Y36/5cMGYTzbXw3k9NKujEimZ+q70FJn9176j4dEDn0dEbx/3px7Solf4fnGS
lI3Xxe4d8cGqSaE4uQ18ry92cT5WXLava5Ylp2KbKQWSIhJEifftaZbhYOVmNAUb
5eFtdgfcNrb8E7dh4Fr0yiKmjOtrlVCP8B8vaz0DkES4LGfTZelMvZlWdSLGZEK6
3Qbihd4jTZpM92c49aFPTGFANu/63s2vj4UR9kssmn9YG53Xkya/y8IwQYLprYSf
n3ykyskmFQbG/rOPkv5Glq5uzjhBNdHwUVfcky+NmU/EfuKX7WRJ2EgCxeiLV6bw
aCpGxbKROuOoCJVKHSpkCQUKkQoItaHShmeuEUefhR4qFd5DRvja6mgH8C+JgQ/I
rw5e1zWvU8h5FHYHhMIZYyUDnhEInGN3pbgeLlZUH07VNUdG0+hiR3ndgWMoLu4A
s4lPsZWuROT5XKcUMuLgyL380LQRKS99/5G3OCRf4Tsm0Za5+J8NsgujhWUnv+LU
fQldYLM6hlMjcCioyc6g85wqfaMe4sSDB6N2HNEnbC7IczkQWc5v11Mxv3WPAzc6
2VGhdpzE8KVGaWzdxuqqGzehQBjrIOPvbmcryzTIlZOo/N94+0LtEprquFg9gabg
1xso2VmAc8xTvsJEkscRsXLY/oL5jMTS4SokOK1lVQWYvnqEXrRBMib6E8KKbXEc
ahuzEldo+xKQZTxkGQ7KnYx9H9rI4/MSjdHv0nxph5lWQ5sabBzfpn32KuqmcSvQ
caxwPLEY+ii/sppuiCU2Si/n9ob5NbWFQtF/rZawCRM9FDBtZuuE/4Ws2bI6v4OW
mIClrBsGreykMjO0sRY4ZSvpabuUBc0lOfvw3cgMsIHkWzYIoOJsLuKbmuImp4Jz
BC27e0LqAzck/HmquZn8lKxhIeI5zbhvWKUPPQDtIz0WPrv0Q0Rf4ZHTbFzGVzQO
uW4qr/es+k9eCEyCfWFLH4jvlXvUmyD6esgik1zgXkRfkfYxVyooDTc2FKTD0l8x
rKdt9YzzzFp1bnt9oxWqo7VUR8TsgH9XE1c1KUaRFxdQCARDqLwp5guMJvV+SSQJ
Y0Cc6fKU+9JcOxg1VPevcfpcOjK0AtM3QqW/946sIkrwTDYVMlUNuH/3LXlM0FoO
tGeTTZ9otITd27FWzGh84VgmM8O2RtRlFUc5HqoqJjclSwl98OmLOde9xxnOYLFs
S6K2f4Y7O+rg4VIfVH6IrU+pn/QsJDFtHV54X4qa31/0IaNudvPql1IgXi5jWC1C
xSPJ1c19cxuMLrrvpwWMK3ij9scd5p49joMrw2vKy6+0APhc9/qc6E2omWGWfy8M
P9SNU6AYYWzPq6th6WJ6Oi3iu7igA2+ihgXCbBq9uFDBcEUUpYQ2FyBdzXcI4zbA
he0i2At3h3/jYv761y+W2pAL6o866BJYYSgclDtYjlKcoPRH0YnOiEnahh838QEG
+EKJrJVO9hgGvtiLoE1hQVVemT4vieUiGdN2tmArLmFItCx4zVXnnS+/w7vNYBub
VDNSFVAhz3YVkn+zDc+Zs8iS4lnrlhNlpz0ax+SgO/MfOAtoaNBs9Z6Ii+cz8NSW
ZAdRQpvLVH8U1Lk94Ap1YrgS1F3VqLLHlEVBTkmeY8nLim6iLWBX9chNUeLEGFj1
3LaH0QWjobxbRmRCgftlT2/Ro2ERVR//1bPU2isN1YRAlf7gk8CyaIF2KSYq5hN/
hYVwFkTFn1wqbIUIhwXFZKq+4acJloD4a7rPtiYN2SG/+yGEKxTYueD/mKIESvrD
7cX/gpFbQz0BMXSMAPe5kv34V050mtyORuaoucXzF5py9W/uFeMj9vMZcvVjh2+D
TYk+30NoCgt+9Tp2vfQrcA5jMwUDnLytqup21zm63c2qXNkboC2zaTjnNr7syH+6
TPaYrfCe9aDIyfdulu0diQ0TecE9s1H3DwaCc37htrr0y/XFEL1C5NJAFONGGM+w
AS3W9AqYYya+ZbwoPugUOi97qw1tc7FoF3zI2DM9n4GRf85fO+WplrUZ2nFzkmn5
YyWsTBRlt+1/0k5bjKpqTMKDQIqfX/cF/rEKEwBQyysxxmnvnqUVIpiR0V9AJgnv
X9gCGaUqit+UWC6K//Y70Z4ZbkGk61PqVS/gfQPkrGLmcUcGPx4O44kwPA8BXeHC
sdoDKBAkcgFdXyFHruBKOUNKmUntDdV/39xXFTs4jYk3Xv2v+mglelxTUzztEcl/
y3ijEm6woAHiv1IUe6Gj59j7HMTJUa+6rsVmC5Lf2UR/RAT04+J8qtg8CM8txPfU
DjNbWd3E7AyWhz2VG2JVn3f++vzlyzG/wfJTFPDRCFRBM4xw9/2mYGo3LLOryt5d
W/mwkKeC7nwk/2uzOhSWmbYdUBx080oDPg8Xle2clUY0e0HxT20xd6w0emizCsIR
Uv7LFtiLxV51HznVnwXdNSPNl75V+6CvWHuUPCGSOp5kHrnoKmf1pJ57f+wca9A7
tdrxyDzkF0OxwAGbPIKdhu5cDf52EFsQdygHOLQoqBDJOUwH/EpB5uJJ3cH/FmdH
Q5D1ZIQ27kW180k/0vEkcxTsiO+AJaNfOGsyKQ9/f2fs9uxCvddwPCDP/g3X1vE9
BCZWzfa+Tc9yMZgrgKKIzyiGjSV9oNcW32fwuY9KLK+PE/Av4PgEEpIYe2R+g0JE
pe33XmD1sGkD1qxyi93vxsGZ+cWIVidx6sWzbWqXJCbiGKaHETCIQ70zLS734Fol
EDW459LbJCQct8Bpl6xFMsjv6vdE+hp3MQhM8pWnWY2PkXAEx8THjTE5lstoPFl3
CdLohnw3vJ0pJ8lixJEZzE/r2bgX9S+ULaDrU9fTFrOxapnokKLiqQGtZl/DEJU0
RqSoG5fxEwtm4Y04DPbDkcV19LosNm5/dYgsJblcgSy9oOLbyTed33H1wQFao+e3
Ix7MGP78J5mGi20uvU9Qgt0God0mk+jBSe3Lu6A2XzUjn42Kbc2E14r/86jzeOjY
wpoUoOyTeBRm2C7qFIvzERUIWvHffO3T9GRNi+AfP8dtGdcacrx8u6XRgrKSpbUh
wG1/X3DwO1Sh0wXOJ7NX6tMN0IY9tH37RJe0tPPrF7LDxxSEkynOmyMXj4/uDjkw
nRM81/6GBp8Fc5vDaP4siGA7Fapjfc7+/5tLeYERUWMQZ3n78gNqY44qQ7br97Z8
F15L4Q9Gvl17u6Db1v8xEHNnrWTm9br5cqv90MFxc4Uar8pS23XJjn4qi/I5aHlq
I91MJnQYwkk5uyCGQd5R9A6hQWGq9Mbmq2v7Wny7hjBqs66ubG7PPoh6S6C+D7QT
sYya3NN6ltic826rRNjo91SqsdFusQdRPsda3L1XRdFn/XpozNNJgA39WnwVZQtl
Yjl8dFueBX7qcr71nLF48U33S0rCoLF0zVPO6AWMLe2HtWr0sJoC1K2Cpx4uHoge
dC4xosn4idnf/YFIkhZN0t3ZNsaxhABsbgHJ40mhPW19SLFv9cBNQnxQOjGaBYVc
ALjU+r0+O5yaflty6m6DrYyhseWWlleSZti+jkzx46xvWjfwmGr5SsGjce+57MMV
//d+gKSL/BjfL72mHDINHtjcGyOn6EshWBCP8ElGWHPTYY0bqk+Jtow894tU7Ab1
gU10/XzNEggcBU6NDkxKd2Fh4msrE7Bxm2SFfXlT2p/dkHlePX/bns3hvd3r/Pfn
+ktqV8++EJjnK2PIHee2Tt4IIaul57CZf9AIIopJ4eiQ9wz+/XhILmaa7QyJXHsD
/s57C/emFGtlo+XFqTrLPg6Mdhosk+qxW2ERjG7bdpHY5mxMxGonCx24n9HvT4UZ
14kAoxun4B/sgXCdhtmM9H/Xj0Fa23Wt4v4aXr549ZRkURCnN4LSpuliNnVl20Yv
3MDmOW16cLq9w2WdVC/ZOyWGjEcXiw6MFZG8nW289e3fq974yGNkZ0dIL11ykLY/
+cH7Jgpbat/GhAGQuU4w9bXhUifkhtBfwKfvxoLUy4Qy7JfeWCTBULA9XVeuz+ne
B89xHQRpIS95DpiQ50csYQTHuavzKx3KQjHn6TZ10/o44o3rFaSjvyM/ng1MdcPZ
Pj7iHuCM8h9InA9PE8p8JIvAg/hZvdz4Ty7Bk4oFknbCLIvWtBvzzF++UUXlf6O9
K8X73A79AuUTBR5BAOCoCFmOxNb9yNYyafx5HoyyMICuav0/1LXPSvtA2Y4swmNI
6rypOdGY/lT7OwfPTGayk0dzmTO7hM02a+F6zalrA3q3HEM4ct9Uf8BYPXzyt68r
k96q0OmNsANcTGJp9WuMa+VnrMVvUT42D+CaqSM5AK5plDE+gNS4V0nwKZpv8Ewx
2aUqV67pHbEGKFOdX9V/oLMVfl751zQgjOr2gOuCWyG+atTE4zSmU89fmB6iiFl/
1c4PE493j6s9vCk8kxLSshWUPHz4Fp1R8+p2clqUKeR0NFm34WtUOgvQdUHVmX7V
m+88rwGns0aQyTUs/L8E+GHj2R/Sbp3VDjKmfcysWq8+m0jJpzEiBWiHPOG1HTeo
mwclokFKZQ0IZJSvb0DLXIsuzAG/YZcEKHFdUpI2Lt0bTH8sBT8v2C87JzgNhd9x
M701hVVtqpPUD0vOBgFDxTudg4IOYMEcH1SK5Bm8cLKi6vvSIzP5k1gjjfyRlZGi
zXzUEnpCo8UJKoDj/tV9hcZL0fe2JtL2gXAkyIaCZSzGPuqZ7PVtnjVjEDjsBZlP
szvAqJHAVjxl6B2q95LXn+r4qSry++d8wDo+OKuFqrVzJDVWqWYXOMTxqXjUusb3
XtvDjgNeV0IGWYbXW1a5b4sJ9VV/T1DA+dAjHw+ozlpc/yKTNoBM+gto7sBH92/U
94P3Mmlhbq8M4ISqK4u6olHpXWkEAARxtJLIsFIhfeSiLc7HPh0ZP33T50I412Es
H8He4OgjoMw6i2c/1OztzOY2yNzYXdsigGK1S2dHGP9du7+SWsECBOjsPxb0XnYK
zJWy2QAJC3S95RARUzH0cChcJsxGDxra0AD2cFaWIC0GpbGE4mLFG40sUhCt+3f3
ixlIcuMSZSdOjH8jGwU/WFfE811NzmoGODTMeh06SXJeu/nDXX7+C72DpdvLD9uh
pS3lcVDMhAVCyDTThndVEt8P0NVR1ix4dLTrupVSwzhrjNo0mTyKvDD1iKZajqT3
haRkh/x9BNfwllp35wuZbcV+oqG/0ZbJrG9Bkv1tqpZuiKNN9jig1fQXCnvLPzK0
UXWJNVdoJIIav9ER+vHsdf7xfmj2IoU4irwN7j1S1aaIYCX3M/s83nRhhkdkTPU8
OaAv8kNDkM3bxp7NXFG4hTJLFR6X0MBh8CcB9FzOFRazPy9GG7Yaa1Q7Q92q3/vr
/WuM7J61NSJ6oTIBjJiE9T2XQ2Rp0YbLV4eJiIUFwhQTzzZrX7Hy3zYV9RhYbbot
mRnwD58UrWnDS3cP6XHF1nPf6ZDvFts7oyd5TNp+AZ0oE1Zm3BRLVBvzw9veiEb+
2dHzPXsJc+P3+lTVaoJ8uQKKWb4tlvMJA44kA/rkWf0nmn1C5gJrNIMiAeKmeu2O
H3WnjEyZ9zduBhnhpAYABS5BRPXDcKX6ih+mUG3ni2sCmsWrRWMzyoZ/woTpZLMS
/EZUHMpdKbD5MmUw6wi8CAdFkZHZ30jgn95MAuoXBe8ZJP5S7DHzJtlaAhHZsND7
r/XeFsTXaZBSe6jN5rSSrrJR31AAqb5UJj6PMM4j8jOaORAGGxVdfs1UWeZlNWqp
otjKSqs3S230TCR5zFvFtGix69EFkHFHKAcbhG74ET8h746Pqtxo+uKAP/igZwBq
HFlJJOSoy5xr+nlHIhALfKr9pBkZUaNwoM7R9chBWvmy+D1sfCYUY2NR8sSAz9tX
jzYkZ2rXn58fQ7Pg22JiLovq/nW9KOiQAx6SSWVMkzE+CXaZBA/qZiyVpFWgBBVG
ZcOs1dv6HDD9k0AFHr+d1DqkjEBdLZLuAKefP6+oZeehqQ2Aiocij7pAarAen3q2
VEno98w7ADfwb4/4P7LokgFmC/DYSqB0/1hEqPZEwi+NNowNkmnQ0RSqJaDtCz+f
HrvrXHNWLPV+XQ4uqiY6JDnJuTzkrP2RriCbaTWYna/urbX348L5OXDyGeR7I+yy
pHxWBNnLTi+84DFEitx0ZOQ7ejv/cTnMHkVHPFi/Yu8Tv/NZdxnDNiXoICfX/X8K
THVsXc0FMZgVwBoVL9MmdiWsRjqUNrEsPiDxvE5x+dMhAvivVtMrxYYQrGLh8axn
B0it9tkBK8eNdm+Qex7s0hUtWCv56oPsezvZr2yeTBK53Y0t+z5GuHW7rO9oB+A0
a/UROthIsY9f+heINOrUWJMS2MpgRNYI7EI7StIJadXg8JnUyDvVCFYf2PoOx7Xr
Kz7r/o1Q7CXWr/KJIWA0o0zRqHGI0e/bB9qlE1zFjg1dwbNBLmMcpiztxZyOJCE+
i6ljs7b4ikAOz4SeBLug1Jqr5GY+XsDmSmxbs046ISwvcigKFbyn8ZYx5UKr/mnQ
GYAvFUnJP/P6NkA54GUFqX5POsqebwZxbvbKS3M1qsnzggmKEEpiTq8brMKCNE/M
ak3kcJdyP/VB4/xxt1qt2+rG19GUYW9doF8WLByqUDjHs2MFtlGVGgYOivVquJkG
rNUcZ7snKa/o3d/jwvRzPQ57qPV+AnVUtweqzXMkiQj+dTdNsMXuMGRPPVI2EVzg
upzF+HzxaiDTbBSFR9+NA72+wysD5vg1x1N/mIGMgxuOUsdZFra0XMbdox2nJQd4
nKO+kbrbsRUTpiSufUxIP4zDw3kbnNaA3ORMwwDAPU+leaftV4MkuY3Ru84Ws3OW
DHYHdULSNgw3abO3GUUovhMu0agC6zNqTKAiJ4p7xDYescWBm4O54kOJCUJnzFRf
4WVEs194TaO35sAeeBAixBLpIK1oY4S/jrzXugkZgxPZEg6UIlx3l5ZA1Vb93wB9
RvuVxU6DoiXYr6FtFnQ/m3gYf/+Ajwbw8i3pTKiebPwWY6vARhaYvcc6mzyApRUI
A7XjGWkxnICQ9qafSvxRa30FpVx6ADuaYFj0qr4bZqXLtHPz5OyJMejO9eEAd1D8
EBvwWWQl9a6QV59gaZ8VBdisBfPPqfs35kDGmRYIWDtj0fxHPMM9KBagI/7UTzpZ
Sy7LcTNmhtVP7weeDu8rt58tTnRPaNjIexwiPWzF40/sW46740OvQQPJr9Xq59J3
8z0O6Eu345+FL7NGKjDR4QMUt5GzinRkknL0LUQod3ogAAAOh7dex6+GvSgYdEmL
dwLfJYZWngbY/mvDGgYinww4YocNP+pJvcUyIi6NUhLJKCHFaDp3AnaCFQMa59P3
lfVPjjlQTfBPWUc7ndoqbTW8bl5jD2oFmStuu8lCUbziixanf6W+lOsV70W6kdZv
6JwP/D74rzTldaQiT/Z3cShYpo3VghSsB0Zm7sr6M2vQrV1TV6rxbb1Dzg+7hEIU
+5vaf2V/hm9veAakgWoKG+RmQA+xhO7ZgQWchZSjI5yiHPlpttXwYmh4Ehuii9nW
UTjARezY28Kz3SCPUUXn97ldJL0maIG898MUuWLnGME9P6Soa5gR8/SPIFEySDcu
1K/BtLPZC5urQk17j92+FhAZnjhFyiuOpbhyvZ/aR3YybZowdwsn4k21Zvm1BsJX
yDP6WpNLpQXqURTlH2vL14BuVLc3jC1S7olrMKoKpHtJ6QsI0SZISeH6Fj6nlqdi
0d4IFLhyF0VLzS5AdP/BGVSGPYPdbFggsN4gw4R+A75X1EHboYY5OqOSYJc8eTcY
xmVa2baIFlq8POUqGiCNPdNNEoZ+Zjgn4E8y1Bt3bueE/gulHVR/x5wRaA6zybqU
WgyYOsC/S2TzRzwo9Fkk9R/Nuq1rOJyQkTLT6H2NLH0/1SrGkqWzkx9SPtVUk2sw
9BOQP3oOsbfhz+Jgd/IDlXo28gDCUVkmBNrUMCI9LmAn6KafRbhL5U1HITDgCg9B
uEmedbenIzfeCjIwEK0elSNxvjFW62qmXydXpUoi/xhkQ0IaIHJiyT+yFGJWOwxp
mdEgG4udGPbxoW7jcUSfZqg+PS5Q+Dc7Mw5Z89366+wEDBQUvRPQYo2gioBgBCU0
SR8NRtzj3lX9rMCWletPlxBBbtmdddvubxKKppRriiH2jxiVH2/gXiudHxPeS8Z6
6y2EKk/8y55iTtw5LZfzXKRhRMuxJOjRWQFPiu2ul5XzVbpjN8Z53Om2UEadadpD
Wwuk1RbGbiGHUjBOQdviunVfy/+SWJrY1N7K5B8AA1eC2oaHVAej/McKOTr4UxM0
OK1VUYHze8LdRPdgU+ZwQ1M8N+J4gb1X3OcfRU8m2oAC2iNB/zIPqEM7oA7NBODn
+R133bIPr6QVm+N5G6f8EgpJSi1Qi00n4wZILYwP7eoSuNzgfrt1NoKRVeArACOZ
p6qKJBU6IhSmxVYe7s32LlNKy417JRwefmRBVNZSApNScgzd9YRoI7oC29vqesAt
w+PqvxvFTKPhzoTtNTvPWn3HnEzlbr1flgF8EEtFmevnWlnq0/WMk3xhdLvRoElT
MuUg7STi2sgKJDuAzmepedxyBWYoXrhut9MIpJSQI2GrSs2bSoeWwTAKL9OuNLpc
F9dYi7yXMHqLMioQP8x2/QCiuiekGqWx3gV1QuuZgOXApRmcslr0HWsVa79z2KdU
7NlUHVSqu+Yo8keMndMRvuc8pYO7aMNRdImMp754b517nmwIGqPCJXBijqt1NzhL
lgx5DelRoimb9EIW3hr/h1e9Y82eGgRh/Ortw6TCGxN2zFGPCXQjWHl27pMWxaAl
BR6jPND6E0kciQiPcH0kmN6EoN+UhASYB5Nv/RHkTDqBuzb2xeYguJkbHU1W/dRF
85Z7IbyIRVC9xXMDe9KPyC34WzPBLa92T2mWfS3FPuUuQBNSOobxY4KzQ/6boIxD
2rqP7yTzuY01mwpMYRFO1a+VWOzu26FYAat8maeV1/pTs5UG5uy+SYsQh6ZxRcbo
gQCcTGLRmTimo7CkCaDcXirDcrbgkMsrF7TZzbI4iORMruVcOrQKoryIpNJ1/ryZ
pwH0c6bsT9pNT+UwIHCZp5Pi64w+8DIqo/p9xHElBz6rXWUT50XDg3VscwItyjLT
v5CekJ3plrwI/4Z4Kv+eexAmo1ea+s5LE0r268Za3NjxuKlw9s6bNs5T4TWU1aTX
O+Pnn93el899Cu9LZd5POF9SFMnYxjVf/m/aaJn5Umb9iMQQuBXOYkrWU/AsyfUo
nyXOtemLfg81HIOzFpKAF3Wwa5b1P8A7nkTQcAIOP30HYegoX0zUAuIcBujaKGNX
KmjgelgL8cFg4ooLG7C3hTHbohVfIyxM9nDPVoMrozyb6AAQtfWHfUOAET0/YmxQ
IOqas+9U/TC+7yRcaNlq99HULNBR/X3D9hVD68rs+MMBvzFRGLjySFBi+eB691jS
SJX7jSL+bTQuTfNeSJvTdS7yCWH0Nq9NOGs87hzWTysHEQLxoa8L1syygybx4pEm
Bn1klyrlRskt7knPQdmphO2tq0nJhwV67aTBcjKx2xaKaFjtBi6dSH+6bN0JhNir
34zLzXgY4o6WMJzhYKG1tCRA9DdcM0uqoyqo0enx3ohGXCZOL+3cMV5a/OmY2FAf
k3IDznOPBHK7rU58L/8fxCYs/luFgeS5Xu4fm8nEiRDc4cPTHs+1coiGuBqP5C8C
thCq5T6+3FjGlZhUyP5EYz3q0RDLXclScfHXfLGcMbMiPY7lKD05I/X52bTov0PR
Ak6vkVO/AhFAuf5MJwsuMbYdwyTJhwGvwClkMtWxe1o8gvqTKI1u9N5yR2n0npeR
qhdOcThVyv5Gq7WuzZjbIJl1WHwPmYbJFilQNFvfK7ihklxEwsVbmDAbbRVmJech
MuA2TYLiz95O+EvSeEtied/NJMutdICNTkQtjLC2IPTx+ZIKVJo6bubesvfCdYTj
SZ+inFBqWfS5imHUic2YQUkkSTQwIJM9mZGpAvMfhPmF/CgnlIOuRntPIW9xYpy7
XtVs33nznEbqqZNMd0mjL+cxtcnR1NQbmhQaN8m96DlN7ipwwhAGyV59jQRnz7z9
ZZ9HZeQGw1dz6SH2Rh1NVZJiDIv35mLQhf5iSx9Jz/FjM2+TYlL7pfEwwiGC5+I5
3VaNlpivwNXVrbL7Qumi8eTVcIK6v/UBa+vkRCGcTdQwVkkPxuBu1/QztY8/auf6
S4h2Euj8OQZEyV82tzNsHzgpYXm1WtwaAd4jb2G6HXy39u73peCzopbe3eUM2X1j
5RyiTVmSWh78mXBYo1atTya5fKO9B/+cgcJaamps3Ewmf+cf8TZvEqidFY7GjlQW
PpHnW+v+i/HriPQf7Np7g2Us2MryD9F73XEYGPFiCKRIFIvOig5OWEgHyrRQy21O
iQ+nNY3+zMc+WB3W3+AzQvNtf3rzhLWOF8sLl7rul/3Sc8aA2fV6famVrhVTPB38
UQpQ3vGG/vmkgESOZxMkV81j5sTy5tGHIBwBb+cODNujFuJehxeSLR1bzKkIbXNp
k9BADdGYwtRfMlpkXj5uvRBfXVLjIp2IknoZzPs2CxTnlHTWpGsI7dugFDhOz0Ue
8HZ+YnVcgrYk+wbTGB8iGHcaiD9iY/qQEuGqDxm5qtVABRPVWQsVBlZsJKFcVVGl
tOriy/pX0kVtePN7xEU3qw6kk8yaqmVBxdLBb2xlBE0NMHiQ8p3EtMi78fyYu8hG
vFaatTERoqCRgJrVRAeO+82vtzCD22NgIN4H1bgQkUDJ7HCyZBS0n7MjmEdFV9NS
dZCYQ5rnbmZ1UockkcPlBTrnNF1PlZxmFZqntWg1liCmkougU3OLJESvpa5uvY7A
N58Y8B/L+xrMi2LpSOG0i5jeZ7cv+D5HDziEgl/adYvmwBXGwwxuck2HTRDBgVrk
jpoShZgJLSQGmmeCHYfbYF332cUpqu1aD1qesDKuKmKE9c30fnmf/f7FmE30QkTs
3ZlhymwRYJyAIhR9/4DMH00fh8+X3kAIwGrfMErkf1jSrymiYxvWYJDL3VA5oGaR
IjNLVJl7lD2XNCN9AZ2K39AUNxpkmsEm3PM6qCLAkmZMVdLna/Vmwbny1blIZzm2
GGnsVTy/a3ZHEAbsGew114fFZiVgQAUHdmCIoteYHscp8bFgyF7H7ma488oeZxK/
QJ+z3lISJ8hl9EWXF9mfOlmrl3PRojxypzcPxpVRv/ozi8blCBb5v4M7VXlNQzZL
Bo4GC4GcUG6eRUjSpOKZtvnUZAOgpWGdIUzTMWUlTTIykGUjuDyVM69ePvIMb+AI
bZrvjBG/4zAiFZD72Z8cSWyr89I0R7azgZiGRPjcweFpAwnAv5h9TW3lBUHmBWhS
fzpKnuPgzy/oOPUvnVlw+lSFmmFc7nd7rbubcyQDWsOFPT4gu5XOAkKKGYrQJ1uV
SLQCLO2N4GwxTQmqVwfVWHk8YXwkoFSj5/pUPlYzjsb0RwJDKX07qMB0towGoUyp
yQKk9yYBiFLcxZWqZ8JTfoQinpXKaX7ndBnTC94Cffhy4z6437e3MjUqNzy+QxuW
47rjvRiRaObwAkK67+eETEKOwgGejdEO0HLzSz5+JH1ukdoiYYcFqke4qmwd3D8k
bpUgzPq2pda62lYM9k2cY8iYsHVzmVhS4OFggQJA/c5UZM02v8Ksa6ILjQtTlVE0
HqL6OU21qzXVENs4zhKiOqirZFFApf+sJ3LSEMBEgonBMHoMlR1WXA4fMhcuB0AR
3uwh+keY97eIn7/Ud5ZI/E6Yo66SzgkOza3+xXx5AWpuJyEHtQi7uzJSkhZ4k3Me
qFsIUHxX0cygAbbBKUMGZInF2mzrDp8Xi4xpVwb8uAL9NVILhQpHEwM5qJfp8jmY
3o3gFgTyd50DKOPKJfk8zJ0tXqocWEDyYfINy2X8tjbdYDMuLf8GBsOPO5VyZpgX
28S7UyheHX/5KXvA5NnIodslQ19JCHoy6HtbhZsagjvJZueWHGW+9yYxoanGcnb6
FeWoZ/63sFUK1lJzX/zf7VhqxdjvOGBQCaLKnESEST8W5Ckpv8Pw7UufjOKNzNiP
j/S378lqTkPENbuTsHFi5rzce0NnN9cX7jRNHNKSJm1oWOOoKy6bRK3Gm3E7LihV
XLpZ9beL5PBinasUleQw33ArmtqOxNae10XUJ6RRCZvdzOnmTBy6bEZ+hNA0UuJB
oGqcSSfkm0BNyk82XnDjXXR/mO37Q4R1V7wkhi45wD3LetE9rR1isn0pVX/m8Nld
CINAx9Hpe1noio/ocr2K27h4zfLUuh2wh27X245XWHKFSh80BmlVpUlcFDCZdMA3
bOskkXej94V7U2CgWldsTnMsQWiefACT6NjzzzkVA6q62VJsFNINOM4ODC84H0fl
UgV7xZ/+Pc/Sh8bbnZsUlII7Bn40+dnfIuPiy5R/VPdscodx2Qqk3/8NSRjiLQXH
nBJuPs305Xw+evpgdnSABHiglR8Z6YwVuIqErWyBsLXXYsV/QBxApP8M5PLeOfmY
AsZb92lIB26iARvIAR/G+LMmQVlvndSLRxtQAujzLHplA0FRTZg9XOIUgtKIakMT
HwA3QkceXgsP/y7zYH/CJhHJmK/TOmUVGnIRQcKnLIoSIUPs+PUgkLcxj/xVMjIf
QUqj5/Ja6lJJnQTgU3NNcVfiIA3XfCa0j+DA6teupzTEsk2fMMAvOEpnT5LtTrxG
iJrz9s9UB1SipTmjKvvq9CMbtRGpI8l8ycmrqeK8QQIhyBN25zmwRBMpSXSNITVf
c1e9vDsaKKrkpm9xIkREv8lAj3jKu0WlJsiH1CrKPU7VErd8jGNP77U+Hflj2jWR
fRK40GeJSPy8aHLA19VqqybPhn6PLFXOU2R6sYFik5hY+pUZmhEF+irM9U3hvmp0
6jqq7ykBsacLLoD80byCerhowErkRplnK48VUZFRSpoi4rIoFlDqnX8epir7M/v8
rTFQbeFLzFRQB46IIiRzdEsK6DkvDtsTm0hi8bP2ct2iDwsAXSjxaolYdHQs9uy8
Vr1Qq1f12ZbgTJrqLYNmB3lri4Ba4iTJINbz1Rw1B9Irflc2WTMrDp6T4iXBrPdV
5QajstvZNvRrVavocFh4unts8feKQwgLUAwzzXhMV2YUC43sExWiZ0Vsw4/iu1mj
vSh6XP4LuKReUvgHfF2YAE1zSjHhnFjI7T4K2u6qCY2OBWSmWl3ij0CYJtB/jxEm
FLfRA27rxxh4OrJsVhWwLFG/Qjmum4cUEjvrMIH0ZhbmpObfxpOhWiFxa9N1gniD
4+q7s5Cd552semNEPz1uqyOo1dG0CCOtVieIWSAo8i7g3Bs5UuskmP3lGPUsHGnS
3PBJa3JyZNXsKqJwNIL3wtngkmTQGTMvt/fG6vwX8Dh6s1QdLzp4sp7e5Mj7Jl9n
NrcxAHWJ+P29JRKWISUDacopa2NGcRnZBC2gACM5P3eYdWgu1+EuPPbHs1U1T4mQ
wVEBmvH/TCj9yFNvpsLOHWb1SmOXwPWF7K/rm2NtbIPhggOJpmEjNxeEMue4y8bq
S9nF/I9HbPShMhtFwO0SKbicogx/X1cWbPrMZmV0iPDKMSYW+zfYMcGrnpeWvpxO
Ja44LzdI1tXXqJkReeeIeV62ZPjHpKp+utX5JvuaAx5gC59iauNVezCGt/62L4gT
/xyUDTEnfxiLLm4lKsY5HMwlD/H6700xRyPDmpr512jRb1iAqCU5nme4mmJ4XpGX
BHaLaUaotHrBWC+Tz89CWPLMnCAFuPR10KyGVjW2u4nwSkovJiGe1cuuU1uTO4Ey
+IVYKr0DGRk0fS5MggyxVi81TtwdGLQ1hu440gf+xUu1gAoGXaHXVoVHnvjXs5Iy
JI1mvlGUSU7KxYt8nFtPjcDc3ZMKZaQxebgWH6bPmpLUqFPK2E0pVeaX9Zu/OTD1
Km67yy1fNfejOTJjEYUdByWa4PCrJn/u7BmwJvy9fefz+gVXzpt/EwvXM7HkALEY
mzVVaCikugypMZt+DT3ONGWLzL78nxof4r87BMnDLWyuXWEwZ/2zn8UPc2TCEdDg
J8ofkvIxbKc3ATPpBeeGhdeT/3Sv9oc5zI4YW/WEuzOfvWx5nyw7nWjRbd54AbpQ
XZ83QqUnIy/XY+P2O5j47xXOs5RJ1jESj4MckXAv/vy7SHCGW5sHv+tsq0W9F+pf
4SvU+yELNgv41O56pWDcPXReiK2wtip1ZEtNbtqKNYm1Nhd6AIJNUYv70iNUCJ0l
d0mxKs3WyI24kqFXO1yJwzRStU1udx+IR6xchLz+NmSsWR1LntFZ3yFid5RDdOVU
kwjMITnoixsNYDuGB+nCukjx5rbb6n+2LfjlLNKq161cEysYHVm8t/ZkgmdUeVho
boTb+H/G0McoVlwruBtwmaVLGjQc/2/ZfJBe4vRsv62zQkqUWdBtG9EhkS3S4L4R
8/N9Qrf+GbhvmivWZFpXc0oHD8/6hFzKOy5yda7WDRaNLrsBbgfwnkMGoOXNKIZn
eCw4ERko0hzhvoMcRwacsXTFgP2Fixo+jlihyeqmZh3fLqMyFElB2vPFSVsMeM/I
5hVNNEts+X9rl/gwbbrN0lz/plbl6zle774LSd6T+zO1ATC5GEzuf36if95GcZtX
JLIC2jI4X9jopthVmkj9Kb74GIKFXX3+qCqZCrePBpWNZQEIbZn1Yh06AxPFq5DY
Co3qrv+EaQUN2/6RjFBJVD5HT3689Y44mGXm4/On0jY5a0k/M0o8qt4e5fbFOUdG
+iIomRZHJndnUl3wF75W0M2jqbTLAAAGqyhrxQi7WMaN0zdVmwKwsj3k9+IBzzSl
NOEaQlrQYpteryCAqXW6Ty4MWtO7k2f9jZtC0p8bpZkjZ/aaKBEkytzbIryjRz9Z
z1fHqzgOhJSpRwrfc2JX6vtuWGWmkIail9HnY3NAjuurHNtBx9+IYF8mz0OIflMY
qQYhtolxZ8Kduz2JQE1R2eUbqn9Bs72wWzuf0qXxrIZG0AT39kHri7loufOYKlBQ
WFuw4kQnbKZnV0zd2lBoIpXu4MeoV3YWCye+l9yz2XWzZlQ3QpjuWXqwQ2dSknbl
8W0GT70g1T4EUHBT8ROzddA60EdlqcwH2A5lpo9/0Mget9jee8GC2C1y/u8qMbc1
0Zb/TSFsoZEIWBzpYiqCMZMG/IvavuAAvw5RRlHSsCjonUSCFFxyh/iQ+X3r47d7
SxCT5eThSI9nvYx2mFAMB1DpyIEuvCJRrx7jd9eZiXSLEn2YmXcg6dCp6VZAo5Cq
lOu6mXYfz+ZteApjKqomV2fwl48FPavkbBx1aF911g4j+WXKO7RC2BDIxguL4+Da
eC6EwfSrQegoOEcXf/hOWPKrsZuoYOy8FeIdf2Og2yC7MHzKqvaSh0gANn3Q2TdY
CyQlnFCM9/kvCbiLscGGK3QJ+po0LrNBtv7d6FhYFqng7Waouw/guCisHOs6+uaw
cpCWaQyIhY6upTDEmtvbcNVssMJ3uIpQ5rw9G62ayPs6NiUiDHSGnbmWC6GUSpcg
8r+dv+iya1L+KSX/ljAJo8Hzf7o8dCHZ856E1JfLIV2c6S42AiRGjo2ZDsa2pi6N
Ogudt+h2mdh/yfQhpLnyxp1HUJpX0z3D2xnms7lwx5xwF2IiWWro3xwYDZHNIcYL
WfSn9+lUzL0EAnIcVWTmiOEVtXw2Oy30eANn+xMRMJYMkxX/I4lIvfdQx1Yc2TUq
JZaJwS5lyua6F2dn1INMJ4W/+GEzw/udkwc+S2u7CPvaKz0VDDoFEWQ2eIao0IIt
6a/51TxZVsaliZ5LxDtSkdEg64VR9+XCnxvDgeNM+L8THy/gRggZOYE8pmJij/5s
e0jpE600p5vvdf8ms+zHLYJWegQRRnasucMK3s3ZPmj642h9vKJpnM1z1kXYYLwR
jbbDuTwlVqkI+UwReJnNo7A7MGUk58yCWaWwdfVive1o9v4f/bq5EulgwoxhXY53
zCPndSukzDNqSHcZjo+0+Q8BQSybldg5rLR0a19Al5e70z9AIeQGr7BjHdjk1nOb
B5Z5396UI6knC5QsTV8xlAVULcmpDYkaIWQwkaNcQMfxwc4rR9td/lBKH/GB12H8
PPNup7TqfhpijCoKZVbV/TriKhyvYCcE9MkFVWn9e2N0g7cnVc5vwwrmxW2rljuy
kUD5apI1qfOUE3sN/2LsaXQcne5lXD72fLOJg9cF2h9cjzjoQ4PyKXtTiqY38bY9
E3bnCQu2NNA1Hi7PmB9Wn3LdhOdJXQsB4TGCk6dMRqoCIeIDV/yDe6ZSiDoXm0Gs
1VOlz4rL3qM215+8XZLjYfsR4ceS8BUm5slHiqgf+3r3tpGY2bjxwFpxquul7BJH
nIHBhPrhC41dx10WI74wYE8JmSU+6cau6IpuCQyuq8SOa+GnTt+hROnHngTVBiiT
nDfKQrBG0xa66F/tRnMgcUSizJ5xof+APt0eFClkOD50zCkzPCAxmyHjaXu13hBQ
E3/x0yU2QLoRGkKf8DvERvzlurbfHAUx4tNVEhNnlhfO5TldQCknqRCc527tEmC7
7J/VEKA76to0NE7Wcrlqgj/USoki/DP0zXQnQWsvSkuMs3uorOF5CIFPxNOVB6lH
i/6zeBBJmx8+kpxVESJlD3UOCT3EEXHtksdAcepipa3020H1dPQvpZmiu9+jgJlt
i1B0lVRpLv5k7laBIm12BJelrUZh4PGFqyX37/4SYgcC8O/xt7UpMflFJoKXAzjz
EoFJzqnrgfx95w1hO9kfyoVYpXFH/rnywqZgMncwGD1Ia5KkhflFnXSqJiyWFipu
f1aXy1O+DgH0SqwfreBubMq9ObpyRShihe/tdZaemcq7KpcFbI9VVtvwo/wNZRGp
bOvyXQrRVf+HqF2ghhHJrCjEV3lQn33Sc9LE8XVZs6Nhd2kxZlEeE2DnxMhgRNGn
+lqDOHoNThfHtxLgMzcnFepnoOF1tKnEtNayqTj9fVCcM1PMQsc+HoaneZdZkFpy
AJRsOBShqpjJNDIKFMdttpGUJiSPgj6WcM2QZJjorYI5NN1VeTYb1HWQUJhpRMco
Booq18VA46rEsuwM9a+avDf65Tzs+EXQjGIqfujZWDg8XZvFUb77+rVDYDsGKUvH
PfWj9YnX32wS+K6Hwdn0x4Pkgt8ocw9KSOVJgQYJgmS8RppJhNmrxfWmMBiCxcM/
06Zq/JYX//9tr9CL97PxH1Sqgi2dYs6XYWexNtxv0bt7VycK5YDuSHB1H5XSnDLx
sdLPz0W2UBCArwzHeJAL9aOkBp8Hq5cDJj3kig2pMzhkyVpSqBRJuC9BZOgUhrMK
QTdX5v44c98QaqK3ZsWM406+eoPug5oeq/sr2YlCQllqnFmWi/A6DDNiP/Zamiqv
6C6RrkxbJjgQleANU5iJ3DiI2DPF/9BhewQBZpE0VgtzlUK426cQR6LJNtTZWdY/
jUSEySCHnLjp9yGK6Fn98WMjSYFddcZjHVwGwKTSWYIGf/Ik25F05dvT4pMD1y0u
8VQqW58U004Spw5T9z+4kxA/hJNnFGmU0KRiuBuU8uNgAmNTz+9fjF0LeMAhGvOz
ZU/YaOQ+tCJcmhPaQrl26lsCXsxZmZRk0LjsVmGXCbx+khDgpw4Auvk0gzUpfcVJ
SCZRw0f+nPkthWTFyPUD+zb9xzhHPWuzYhE7lts599VW1OH/4+sogw50ldi/YFHI
H6lNMeS3k3T3DDJUnsWKWHejqwH8jHnWOHOfFy9rcfEqr3IgYERNmzkoMZuLA9g9
gJdMDVrxM3ryxCB3JpQEtxWTgAFtEU9NKZUyuuhRbsZk9Ny8UEuZCyxqQ0756Y4L
UgTg95HUL9XgV0Y8yePuSmnfd2YiSwziQVwXa9uohJxyMvA+x3PaoOKGBTyFuXPg
nQ/2rB19TMrq4+04KbTrrFnUKLkxYJcrzC0OrEp+R11NK9eg3ETlFp3mGnm1JTUp
SNpounx6VmdXnpLb2YpITmB4zyupr4vH5+DfSLnzmbcuKmw9FaImG2rinVr2KACP
EnQPWxdTvgsprFMn6nSkkxlP5RYZ7laycPSdm0yUiRyZM1QonCL8eX3Dv4Xy5nDw
iKQURQaki+qa5TuLpP282NPHNd8UNiNWmXd+aL4SVu4z3s/RdHBcudyMS4VNElKX
Ir+OgKbF8EwrCpRwHckbTua/ELmcGK3di27jt4vwVGRJlH54JiloduV+LoNjQjXN
20JTqyJaLew9JL40mEM03bIF6t2YB/fENaAQMfT60MEFShkr7KgtBgCGlezASiho
euUps8r9E8ZntnjnEl38Mllg4ZnrZbrjDkRFPFpfpdTptvdMYeNmbH3V06CUdAy5
qFk6oL65B//1Lp2eNSuOKPYFPNmJZR+/Cvm8SYWXNsjrTdoRhaiWTQMBhlbj3YIZ
TNh0oFCXoQBxsn4oSUVprr+4OpOfpKdfESB/TkWc2iMSO6ENHW9QWz+kE1QIaOSZ
7rtz7aTQaiMhtoE5WtB0e5whNsuee2m2p8UO645eNJy4F7bDznglA1a0dzG1i5OW
Ok6aQrtK3RDTI0L8RHUaeXiqqtCoHXBFD+PEx9e/4OgMGoswnAxNizzqlTxMhDzi
s7NakCcqmUcSxNgAYx9wXASHBmDYFwXjOL2QNChWqZuyjuz8LPgINwRfS6ZkBJy3
rN5uj8NzMFt9f7K98XaMxUbPpIzGyGYpjCkwFTtDs4eOtoxDankvDi/doYpavATw
jXVaBPMbYqmQQWmJL6MPP3kjAMK1BaC7H+vKTKhkE+azDgY06gBZFOJ41u1H70nT
oz0KatxUrS8U539ZfEIcc3Dx9r3TurzAYsk9skNT48usOyC62hwYPeqMZHDNK1e8
gY2PITd3M0Z0mm51cxCoMK/6WYT9JDaA2RLXsCro08oP5k6V27tVfXGv8AN6+ISm
qtI2bAQgN5F13PmMKw4b7N/BVCK1uvXr8TRpxagfvFZzPwJkfcOMq/EwGl7wxb4o
rqcAYAlhF0wwGSroDo4VsqPvgPoRXXYWN8Kq4Tidnho+fWvVUZN139GN5IcvkvBz
xL3wB6SNpRAFTEhg9zJXZVUrNuy7VxoQVpeGNeTXFLj0l127YjYrzIiAZfdkDbR3
MPvDE2TIe8qAtjm1ckBL2V/4nu9rOU5zaZkwTyPmHBev6hxI326j2LDx9GwDrIb9
gcdiredsqaNcfVmSAhXTYGCgtbt+JCJZmulQDSrQq9Yh1Srhl37TY6cw81Uc/H4h
hgBX1ydoRIECBuz8t0Azf8fjLr5no+SMtHaUa/VuRrhVQBZ5b/qlZho/j9xSiJNs
Z6fBZ6Ulruv6CWy/trphjGD2OX37osHTDnzhmN8hSacAwRy9QgVud30q2sv1uSib
9Kl3Um/rudWrH9EvEq4rTjOd46D7rTS2sZmA/hOj7ZeC1KI9JE+ssTbiLsNNRKdf
CjQH1LSBmnzpr6A4R31pzv8JcDBOI8Qq4QywIYWDPA/+Z1a9kFlxKx9zPu3cXDsy
JGG0G2nVNzwxDUqBCImKp5Q9HmvjTAfoX0Y6RfiybVYzPnrw7qY4WFeGIMKlJfVV
u8Sw2hmtN8FeuFMM/vw2pc7jpgjZ6sFUPgM2nrhKC7VojqZk+04GN7++y7jujKI9
RPR1ZU0OCLbqVSlFQncPLiEcwLAVSKAxmOlYmM1A+Y2QkSLqSxSusXToPlA17Lb+
E1uwR3lEjgxCpqt0TOxJHS3RjbhRgFGkZPgs/0Y8RBiLRm/vnUfKPmXrD7Ibxipg
inUHeTt2cVraJ1YxS5PmubsgMCAR94Put5BJ15+v39rcDMP80j0QeQzCQjDFs8WB
eto7TyQGfg8Q1kNwaaH2j56UN232SETjwsjqO8kbQnfmEvrXjtgdw9GHuX/rWdX1
aDu+0bhOFH++PsC4iprxyJMFvzmj0+V0nN+kSlaEnGrCSBwgj6vtjNVZsFBZpt90
cCzauftXtT+XR/BWOXZiRBSeydJ+/LeLbWay6qWm7alDhJOoN60nDh200nJrSYFL
SkJViTpYotMU6OeKMAV0QjATsGdyFv9TlGqIlUj8dx1Dx5X1OrBrUlZifvAiWlJi
c98ybm5FWdg1jr0yEPT1AZRklT4tqOO74JEBLdLQZceW13Ct7VN0dl8Chhyjn64+
VskevpBDFCoedskXilqHMA+mjNMYpuMcLHmRFY1/4JaYQ+2x09L8+s0oANsL9YUs
U3/PqJQQPSjlj6ST7UBtd5CYLZlbg1SWEwjPU9MXPwd/SqnhhPki1DbPNyUPy6p9
FuStyIxpSAsEIYIvsbUa03rIGYzkERyNypAyY+dsPFB5nvhgU9IlvXz1OmECfX/a
FOSq6jr8ICB+vdbEYC82tWv46FVChtfA8i1UI+42HqydrM4fkNutg9qi+jIFDXli
4SNcnEp2nizWBswb9q5LPP/dXQjbVEAkwJqmGJgsvilvFopw5NFFuDmE1q2/zim6
v1MW5CimybOwGPACMfGGr5HBdlKdv+UFbncQZKf3NYYxuiETonAvAuP+PamtQSG+
Tps6LJplMQ5kGWVgnQ3Jg/cUu3feTt3LRQ2TVyIg6x+3QdOR+TzoWBrphv0jXXqU
SvQ36zsbXfE+4uT21u4aaEmARtdFoVCcC75VlnEoOyi9RHzvFLJAE+qH+eRDD3VS
7QkR1o65cOTGiJdd8EAlcabTC0v7zC9Ed/h5W3WwkVSAx8pQf2BbubnUedn/NlJ8
qe2Y73MSTe/5djWWKAuRUVYF/AQWG6JcvPTVz+VOyupea8EsDlffJ5hu4iRSQTr9
kzGN9Gf5geZr7cl1cmQ6SzG7RPxl/+cjkxJOEqC0ss7s5D+VuEmL6lcNPjUdCgk6
2Fkg02wtJJJenuCmy1KTexT4B6SMqKZLfnu+TED5Ozj+mVmAPf7yzPlP5CTGKVZf
Agufo0LHWpRg7jQM9in8qv7sx3mXEOVw0Ph14MdpmZES9usupup8V64IsnmMYEhV
GA8opnyAcmNl6/wBs8jxtplF5/HLLKFkQYOFOSKBtk2RTxcHgWY2ghUBmKPVh3hK
8S66s5kLzrZvumHv6P6XLGBkWHhXvNKz18Ka471Rg82FNrEHt5M+c857xT+DSywB
4B7jU1ZL9RskGdbd5dtKSE8wG4DKbixOmC6lLQAJ/2MXSxoJN7OhD+A1BjCgNJHD
FpmRK2ogvfXV0M+uMox/Lz5ke590N6LsD8kXWjxTGQcUN9xc0XiiBwKCmqHNykLr
WQxgTD8P4W7KH3ZJegx5UrfrQ/jhkvTu+I8zfRvuOKwDwWnvbHyQAgAYBQCkz8RD
UdgQ8AKjXXGVR4XBmM/xHeAsUmWGKesUObfWQcqzHUUC7TalqbEVDDFpoC9VizyZ
VcAl4evtmphdyoj2NZzcjv2Gg4xbenBSPDmTidPKz3lPI+XSOir2culyp4PFR5d0
/JFSqJDVAVxoZ5xoDj3I01MDnXWYZQd1JAk+DKuekWv4RCj7gPsuycAN0FUId39f
IseL0/qpDRjmVUP1kphAZGv2JjBtL3CLHYJwft0udvJO4E0K0qJ97hAtVbX+gDij
KArj0t5FdgbkXYq/m8G4ZyOU48G11N5Xqt3FYJAYAk8DfDgMa3KGEZmTM8z+aAzR
V0/HAOs27zHUPY1KkDj0L/KlkJWaO/WmxEYW/d616CE5okDUDcdu6YvLTc0NXZRB
pYvJT+GfH1jRjcLlmsBrDlMPOQwd+ZQIkDKf/fTfKouoT7+RoevnbKzm2JgmQdjC
PtD/kPFUc5Ammo1RYniMemas4Jq0tFwHxTbqUEuYp9iQXpA97Pqe5iXzRO7yoC8U
AkQv14Ip+q1WgG6BEzlBG+vc+26rJqtAcDBdggX7QEvp1MoUBWoNXff+tTJ2nSmw
+foaGFx6LQJPUYqrXEVG2LTby1jdaQSOjjPH9LwXU2Zss993gyouE7RmcREVlQfZ
N7YveEpXKOK+cf7tAkBWuENtO882C/VUP6Mj4noefceHNQZ9onymqSuEaOkIHcb4
KV/PDQF+q/DZ2oFb4dsVaURZ9226nPn0TVBGn6LL+WZCSTx/dfzk53cAlTQa6/jU
1UQ0x4NVREZXZPpcRHL05w3Cw3+0CvKQbwi/I5BFZW3fV0RoW3Xg1A61ZNmUB7UP
v2PlLy3hc4oJqlWx0RgzwSaDakApbW9gJsiqgbTiHDRYpR8kiuL9qmGfARgytN4a
t/ZGlh7N4NzWHYkMIKRmjFN8GRwF+LFwB1mfy7/h8cJQ87MAzKtUgd7P2Pw0beXo
knEKZN01C6NIWCrWDiGWYf5VjP3LE/Os7wStsboig3bngx63rXm/ln2hJ5Q18sAg
vcXemH6lNy1GEZ46NkUv3MpHzOIETrluEdhy3tn1L1pPNsDzbamLM1EtANj5aDJg
t0VjvAKxoAKwrMltwohwH98wnZ5eP9rb7Y8ukcgI6pJZSH1faMg4Mdhxx1xbIZkE
XnNQ2PChF8v811yu5SfVF0o7I9On8WqQY2f6/3W4ABv2iCkYusjRkS+Juw6Lo1ZP
/Y/+DztiGZ698kN1Tp3aS9jIxRvFTwYuP+kR2LgldsJS3r6h6honGgJ/klnXflNK
hcsCrEAkUfLSrbpIEDbbvMEqFRqK7b4lvEujba63xWV1ybXiNOLFtY4eF2HHZ3k5
rW2IQNExD3s0QHnR07GimWwZtBMStZDJCn+2tiUNggQ5JgKC1yynQ/eKdIbmBrpm
j+Ced2qQTo+yEUnTlT/oZj3EwRmjIndB9boMZPyqmKn7sOo5B5gEPT/UQzn7kNGX
hRM0k8iWHJJuT5KJEBNkz+TkSpEKND0yloh1fMz5b2b7vNcBmNe2+KhbRYBm+nH4
jnMGdHio1lfnaeAzZN6fAfsV91xusVtNs+/2mP97dENoAOHxK6hJ4ecrssKmVxxg
/BtdFkXDISHKt4OQ7fG9BYAT90ghxrOOyz0RgI7jCPwc9tas6F1nFEtQ/3UfnACd
HKWr9tSDRitwgTxAgMMQB2BEe7ooN6t0qTRX6Q3exusuM6f3uHionoPKpjKm4Gj4
qCn1h8kCz87fy+6N4FCLVb+Y6qZtnaz5WyBUP1NfikWLq5Y7Y0Fsae3DrZZME0PA
Z1BUIe+jV1RdtP8FYiB3aVDFsItzQkHCxPDGbF1Xfy3bDFskQ4l/uN+VpZEhgImS
q2ObSt0Z7Wwyr6p97xkPOK2sFhrjtH2tIClhcKoeU4dkmzuPiJfalIs2Hi88IFDn
tyM6wyFAb4VDhAe7nbwnsUYNZpOoYB3EbyywT4cuY9r9gfxDIZX2bVBp5+gVhcuT
wCoV1nL9Du+/JnmKIs3RGojDl8HuK2a08YkAfMzWtyMEKgs71hJnU8moFOzE9D6X
MXcEH0TVAuqtXfSK3GadD8kcRVDayZDDpCmXI/sksgzl5iTTXM/hchoXWdVnlI3p
LIPR7AIuL5FjaxaqsVgY/+OgBGOQW++wWscC27lWSOn9iXEqGbS4jw11PM3SxKMS
Qc33WPF+9/Fo3jHie2I63W2bRTsNTdG3y5ujqe3gvljilFbXymcnZpUV9q+Xct3r
gj4A/kAfrO4OLt+VAznhBkYBTMjHjC+Sgyu4ULk7MqiI93nwSQ9V84NtuM5vwBFK
a93ZFx+7v8VKNbA3jEdGvFmBLJ6T17LqShiYI4OvyhPQxZ7/AA7K2U7RJslZnwyd
0bxpMmBXdhdMd8CjIoeY5I92b2Z12CHp5sXxC0OUwKcOnC7E2Tm3DF8290+PQIIa
8cU0i0fhBeUuemnhSouNGdjDYKYwMhjbh6D85EG5KCkWvwa7dv1xXAfF2mB3zoTU
AC8e5p7ozgTIaQKZ7hdtcvHIFuanXrSmc71RLFHDTmAB8XWJ6hsyVu3sr+bwoA6C
DsbjlvCbC+5oVhgfbQG7gKOCBj1l7HAanEsqFzwphZqQg+eViRtL47l+G0Xi0PRv
xdcoXzSZow4YMR+dwfsVTLeYiGdYBRD16txdh8b+e3sl35wwo4+bhMzW/AWsqgD9
lD+s8IfC0SSTpfeQ7zP2TpCSVqJDHPprwklCiguflaQZD0l+/f/4t3vwpoKisQaZ
VEsnzPb8Ewx+eqVu6tDQmOy6YkwLCI0GhT3XMMmxrqx3e65aDpRy5kvd8Koj3NrP
wCFX6l+XqGLENvIK5Qt4KOrJ+Ay9AIJxJpSfVeEyx7vgFi4roDovu3yp8nvzyBm7
q4fgTNzrRoDbbmicJESizIyYEUgHDMsj9vczIGiAPPgy5qSNRQIixNLSw+eeh8dS
3WreZxme6rZ19HXcScFQuS76NxTo66lemNW6rcJCtUqrg18XChOZg1xr/v7Az1px
aJ9SIK03QsoMIYb3VFNJzT4tZ1Wehspk30g/IuWWCCOO9rhSA0Ra4k0fG/WnTSB4
R8RGhvcFHqHxOo6C9H6qZgzRsT0X0dvhqvR6X9ko8hTKOEujFWAh1e3hbUyGcDY4
9KZCz5bzqwIqqZjSZHxDMbSk1WNGV5BOHOzQ1RVEpRD/+CLO8/b1WoWci3u4OBTu
/8bBfSYdubpP2brZplWbGRJeCazhAOmlQw2A0wxkz7uvYySKH+iyW0MyKybcg/xc
OkRlPyj6+b9KeqBWlKpIbzJQpw1lR4kSTv3pWXx3IuCQ4zLpuAlhNbAuoeF38pWK
avXY81s1Dvo1MazGAGfdswZ/hjJUMWOSLKigD2Lg5VBsqg8w1ZD7wsQd/T1Tuo7L
mAEbN2+pEfqpC0N/gg2TdS53JKwiurno8RV4TN5pQlxMMXXRYZo8nyPRhZShNTU+
o/5ay7WdI80MoPiAqgXGnBBcAgL7e/eSaeZzMEpLSt1EzZfcCibKqGIBGgFnE0aS
Dj6q4oo34R9aeakZnkg7T5nsfdNgHMqfRhsqeumEFdWF4+1L+4fB1pABztMAs50D
QtPXYXJ8wJT9BZRI8SIV9fYqSeIrK8JqevsZbO7YTT0BqxUiCL7celHiXwpsdiWV
FQCiMUBSf8nucFD5haOdQzv9g8clPO2z1i6cqHD70M6qpOoG5/wVsyWLo+13xBmR
jVj0/D4HjHz5Elok9qOcidtlFwCEIzn7s2f2LlrbhJtfDlLyrZUiN+48Fik2i6ei
/VUqB5fgJDzPvkKeNiDfzKhxJt+f6CNyI7gM2w9S9ALiXecq8CssVUSsIu+QQaV9
d7m1VWMoZjzGxmjiKpFlyCiU4ADSQrwc+iyHOP1XuZGxa2T20TH1vH6F1vTwoS19
Zy0D0wpjTF7U9TMWcAutoD7dmJ/1q3Wxy/svMidirTbeVhFRwryyotfvi0Rs3wEn
gQ0SkYK/2ClgyMtTfb++HALeU6G/p2NE1ry/kRiQczgmszHoIEBxgCwL0nWuc4zw
/LilJKigm7weOxyNXAbNWwSo0KBUW+DYh5z+eW+XrMxLm3xF/zOvq+HjkzDZw1kl
fkUkjBzRfa3R8DH1Ei7jGbchVyJOTnRKps7e5+M0TkywWmfLAQN04dRlLEStguv7
4rIVvjxI2Q+PU/oY/a0/FLGFQmQl5xWBOg7A5scjLavFDARxURhqe4GVNYXvk59b
xUAcznyjc5oh3cADxnSiiv44vWqegAXvpuMaWMRMsWM0ZIpfeaaVgRA4TdtfX5AY
/UjP5watzk/uUUfaJ+G1t/xbdilXt1B+Cih2K61H3b+fgKnDwrj3rYbj31QYJxe7
Tasgdwgp7lKPEtRMsCQbq09HqYBj0aFbNKDo8bGKpOJZTj//yhP/83JaQ4W8rYYC
MWBmpDmNsXW4GgXsrvcujCDdmib19g2TSlfCZb++hLdi4UQJk00/EsnZwZZ+KiXD
Qf3OwaKIripaul4uV8yLq8wJY5ohzJ53vla4igAmQ0xdiKSOMKaL/kLg6Gtmjr5z
2rdDIHfh5XKIZxiMttEi3AWPlYLyUo+X4gHx/xaF4VM0yXu57Rh3pFEPdclWvOBD
lQSiwJrmGMTLrozKVqgJGOkcgQh4G2HQxv+cC2gFgfQCz1uTyJveb6KXTDi07Odq
eNIooJlIeNN3oZR+58VZ54pkYENV9+WF5Pf1GbtgczgovC0xXYDEAS8eHrLTV3AT
TJ5eG+bPiYnPImtioo/G4wBb7Ygmo6/4n+/c+facli70MC/ShbkUXDJCnMfv2uDy
BZ5vMPhOgsXDKDUxgzZLJnn0KYaJUKb1Kkv7rQf1moHW5jDgDtfKa6t/uYU2Dd2d
fDlDDwKudgqCH206aP3ijTdONV/lqGofpGGGHxXg1VIywKstZX01Suq3ez/U1UzG
/kGdu03FHpMRKxgWsop4fBBRC6/C/BuCX0rGzUOQ4OCNu9lsZQauvX2AEWWgAyGw
q27BITVEy9tv09JwPcBLJ34rlWdjEHBNW54e7El+zgHn3kHbnF4Jc0EIuVCHpPDo
NHiJBB7pVk1442D3291keaGEP1gQtnKfFz0Z12YXLpo4txehOD2FiW9rkJU1JpO8
YKQQFGvyUiEusGOM9pnm+VZ1ucl+3FUgk4Pqe8vsaVFAm4gygp1MXEGrG/Ge/yBV
TOYYlRwiWC85hi0J6W2h3QBAQ0xmZAD7nx3Fian2v1ANdV8Kf/U9XRmkOzwPkrYX
4KVqNUFNry8T3HAWIeq2O4DkqOwzawUQfEEncScvTRgycqb3gzWIT+3+CQa4+BNP
2pgIjAQs1oEMqDGTShNBW//9Srlop8ZdvgXiYwyzoxwIfGkd/oLmRw7yAKSOCTtR
0c2KiwEPoO1hyQK1uwHR9FLXgefmojwirSslg43MSPdmWq6G4V9GwbbZ+O/jgvIt
FGqXFGAjRf8CIycQ4OMzsPSmwRBM1TGgS7cfoG+gVOXrEWK6qCJQCR8SkLHvG4Ku
cDmyylN9O5gHKPlMa+50dS7N4kIjpqTiJO7Sfr4JpMKzTBauN7bmI6P6+Do37/OB
lp+q3Qdxy4EeXZINFKl5ZWfoA8QBMNUYY2o9eAQpHKzf7T+xhWhHAEDXC5ow62rw
eg7QQd27vcdU3ce3kQfDU2WrGpfkP1Awt6QUPW30y04ZTjcswv91Ul8LjStznDNw
bFd8NtR+8V4FenOP+dVL4CViwZ7HowPwWY21Ug7ukg7VhWKKtXr7qy+y6rqtRhct
LrO1kgguPe/TlAtKvddToJmUcS43dH6qMQF2jcYOhQ+yDOY6IB78LnLOxyuqDrvu
lJ+0qfewSXev5UMldSPKkjznoCblOIJJv9BHpDJyyTkvT2P5DA53TLtqGWWxgOLv
2Gf7NXUyabIED/RCH1yl1aqoQFhi1F0YXXw4/S74dG3fzzNzZ2l0sByaSjGtsYJ+
I8TI/eOzdE09IrJHk5nwlxr5hmy0kQedrkLFBRMepxT3RvH+u1CMmaVpZYMShuGV
Tyd2rqofxQqazg48X+iFyXJDLjyleFCAFa1zb4uHTwsZbGXhouc8cAYTASsY74Ck
s9/VtEtREuxuz2OoN9or9rQhjhIToPsaVx38ExV30k69qCPi6dRRNfkBW+KMA4g9
9fUJ+q0HoXKLBCToOBWRYvkZwHDuGhGvPWWzBTvHi6Aks+Avm/RXEU4YaUgyXv8h
pMYB4fYUwZH9r6yUpNUivbaEjsUNuMuBRl7vjzx9VuPX6HHdffrL1IyRMk8ggFH8
cCUYktLqPqGQeMoVmg9LEogGQyfDldZpMU7BUdZqWY9g0aleTCxjSPQmjyXmj6rl
nwJWYAhRzWRHNL4E+0LpJuoyM2CVyMXAJdlnwER1VWmy0ZDJt6WzXoLADec1YK2Y
mGQehUMB5KFZJIeAGRbP94gOzxVKe0FXTQc/RciY0NfST1pmQmD1mjXaqwdrRHMN
JKqokpoyKBufB5N/obuMaUc1zGU3PTqG+Jjm/9PXItFBaFLVocKQ1uaVfaFxvNva
3aoaCpjLLZOgzZHygoEr1ya1LdHPumkGEB+B9seyEw964xbTqObJufVDmBmdYOpQ
EPM1n0v+LR+xUWgrmB+pI4l3EBvC/a1wSvi7vOiQVcB3vju7ZwMR31BnYienn6/3
+yJmgl7UJp55SBKG6RL9YkUVw3aWCUI+woCjdPRbgMmDoIhw+x157IzJ/knSeDYL
8q8h65Y+jo8W/Tjn/m+VNDMpfO8j9p9oZI244rK6edy5ETMOpCeqbbFUNlM8ROlF
HVSkg43UP3bXezxV0BBH30JKcHEuiMiu9WvSwMhUiZi29miEKRMish8J452yVVqR
hhvtlgB/TjhEtejQjpDHIifAZ4lGC5gdoJNQYneStOj2Lz5c4e+o/UJLr80jLIhy
cS3yagswhPEDHowW+8mZyTMWpMrzckmY1x9BTDU6NQNw3tXV1FIOI5PdCvJ4gBYu
zZBCXpNKTyyMBTR/uyjYOBc+sCnTY6fehmyLBXL92+f+DWg6j/+wsA/9ZvXfdbcf
Fj4itZoINiF99QM2nJiRmjA4jUNBTEzuakwuMT5vo3cpml39Ync2Y/UtWy6Vi5PU
we5r5u1ArnBibJZyp+pJUrXfdTT2yRWYltfbBd6JFCM+CXWnsgyONHnSQzPIA8we
djgmMpXXScJgNA57TJf5nkM7/Rv5D+DgcPKVukTRiFMf/wYBSDNw+/vbSkXTEghQ
kUJEGGyTgci0JYRXl8Rnmvr1wN/BmAByrOQePTroEdMwrMIECKbJdmd5U1IBBUUr
EebMJKzbzOVwFV5yIXgAr9hx1C1F5Vrqvl+BCJ5GXcASAmCqkCcklA+x8HBg0Z+v
HRp0wOBQeNj177cU4+FhPkoauA+4unnnRGp9LTyrYvd7/axQvpQzkpI4XPxlM3MO
fgHTc73V6OKb/PoPyzu0dlcMEbmeB2gpnYkcegj9zJ+ZNtI46OAtZ+Yh7nZ2+fD8
ScxCJB5pEZ8O5DkjFqhar9BQRR+IXwp19SuVWColmcETgI/WqKda+rflS0dbOEIN
hjXoAfIwM2oSqSD0G8D3nx0O6SWCNzDU4+4nF93ZT5x4WOtBS98nIU7ux5SXa5v+
8BuzU4/k9XFO5gQ5BjEoOkYBjPmdLHmUw9iqxYQexQGtHVzFb0C77cbuX40jJSs4
iujwmkIkpiteGAaKopCfOtzirwm+Yy4tUPNQicV/33+2pvyVH7VBU33Vp0kZUgeQ
zh4ryRXUQkDU5lIOeZZJau12lTsQpufdvvUYXZh31c6OvS+2OJCPJ93RUK5gBZer
mdoOTDmdE67axj8VttfEy8aqELqxbpo4SLNXNmzfNkTm9T4UaYMAT7ZP9D7GwYzP
wXp04OmVvST/0zm/CGZTLXxeLq9pmetmXP/zVOIzxJGv5NPlTuOPZzZho5HnF/MK
WJ17ad2wRAvEb22rOnqZSA+YDIZllM+qUUfxtzIcHFWrPoMxR6RI3RGt8cwjHsv/
vDPXj6oqZMwNnygWK3Jinszq47XS9m+F5dvHz02/jAJWwvE9DxxbHhqoFhI3TPjB
7baIahx4pntGpkSzGxwNrelf7v0mlRAVNocbEpVlAyEcXbhMR1EoIHO6kp4+g8rK
QWhjMcPVjj5kK0uYDtFVk8SCVdEjVs6w3nRhP3fA8xc=
`protect END_PROTECTED
