`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKwzVefqS+UdsdNX61KYI/kUC0E+WSLl44nJU5IBWPyZ
Jcwr5MF1/mWTr6u0xgy6Ld9zw7pPVH5DcIQHkLASrpYNm7hdypn76dxKNYleDxXW
5hMydqwmhkdKam6RIzcM/IH5uiexAlpu4udd746hUdj5jnQ+BEUBInD+iJO9Rhr5
`protect END_PROTECTED
