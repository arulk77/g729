`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
CfWexObW+liD/sJzXSjWsZvXmK//MNwPifHWo/9K1f+IGq1LPaRps5WAVsF/b+Kn
hu2/ZkAUf1X8ZwSXHG08jkeJMFErBSze0cfJb5TAzn3ab9wSSDC1gcYL6yEdt0R/
KHJ9MKv8Un74iX9d5rzCZGvwGscQJPs5JGmtXPBsYtO3n41R3N8ZUIE/rc88hwFk
3JduxVIFkeMkskpRDxXpSSqVofFHMPaFIIq8rFpttWZuQyhLVMqoFx5B2GuxP0R/
nF783tWZdGxkirJ4F9dbDcuvrwzwtlf/nj8CqJhOHKPpEG+Gx6238aFXt1cgzyb6
DDcunp2s1EBubW9L9rmrPANP2xkhuLnr9hLcazvFtZxpC9D7YGrTqincXnbGvGFx
qoMnQN5TXbskf7KdRNAjJQ==
`protect END_PROTECTED
