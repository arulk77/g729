`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Imzst/GhOv264eflPy3U1X4cd0wxLg0oPBjHNdYspik9sxDGCsnX/fCPPaLCMk0s
SSCUaTooZKZX4jDvQQu254evUu09L3PMMqaAgBl/hKG+ft+EXWl47P10KRDa4wVH
lvB8W5PSnHsN/EAqbSqsVmVhOimDomaqwzossFCpNa9y8flU8989w6WA7C42hrlo
PXw088E+LM/HNfIlZYiVKxMwHjXHI6/S4cXyceE0EWj6lBmCjjGG2dEIYUOVqIy6
Dy5Cm1ihhd2U7cRDQF9j4PjhvBXJ/8koP/FmfDc5rD/GQRFLaiN0HrD0DTn5K3SD
sMU+AChNn60ca9EhsZcSMIENMzXnBRZAXIjAUDzJogg=
`protect END_PROTECTED
