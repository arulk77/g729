`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNxSWTN0En0H0hEobhsJAaTQWgicgMv3ulwneuEfeCkmC
SU7Vk47Zgz1ebu0SvCRcbcVkrUeZ86rp5eXHMepC0NXRw8TVh7F9xcIicRUcntH9
3EFt5Y/uoNWbjWU6v5ufe4Wkd2hyCDVH1D0MV2tJXNiCs43ButOm+9vzXVSd8fvb
WcZwrihYGFNVPvucwZ+yPCdAG+kJx0iOwa+Uz5ru26BiT8urVxFgIryEPOjA4Fom
Xaw2/wibqFzleJGj8Yyf1Azm221KdmhfboxO1TZ7dC1P/kvRjMEayq2qW1lPcH+g
OgqqpnGCqJCj9EX8+3NyIpvczgy35FodKzbaeVsJHh6jH5a5dxRfuYHOT5+FSTCu
U6FFwRXNmnIaqfLXYEw2uLyAdRznXLyP5SpFJ/Gj9ggGoK+rHsdjZax7APvD5twd
N0z/tcMz47sNT1wriceV9YJRM9+jn5pbYrwGdllgM0BYqpLNDw+9P0/DHBIeZan1
AsUvDfQchs06JP2liBEsaU2fpz5e+pBnga/aTJyeK2szFUPOifRI0ZR5ugDegdH1
dFXmhzcI8Hh/VnhQdbL5nSRLJadZh4xTPX5byZDUDqpgXbP8SuRVEq2avXKAr5N1
fVVhWeUcHNOaacltjDN9CtyLx2y3HhB/S0dth6x0YIVB1ChGtWEwoM00Q61xTdOj
iKwQz84/kaAQq1md76rFC/ovavjl+di20aYQnyOR/7UYb9FHN/87kc/cgXQXtTWM
gsw2YRvKHBSrXUtluNV1RimZv4BN6otssGmGJXx2DKn3rN1xDt5OW+2u2KDw2hTR
kmXnJQmGkaZwBp57AZZijfg28wItGB9B6qExvtEdz8LtfhthpCVbUbzZrl628vT6
Aw4IwdxxS4Lfyh3041sGS+akQPYEkzhdJRrlN3ocFpsCYrvFnU8vRA/kNxbDJDJF
zhoucS0DKy5B5L9bGnwbmyG8CvWrsHoaepQtYjMdrZ8IsFxe/pvSOD4c3sfii3xQ
PlH0ygFJY8FORxEm80CJ6lTLyv70RxacG5Zyk9BinKkmVTVRMhBXXl4NzGutRZKB
86dd16zF52H6is0sM/rF6OalTN+1Q3su6Td2RsRc/UsUxzhPElvTp3leAsKBDSW2
E+smOx7IeBsDc//t66GTGf0idH5NBNLPEuyJvRmhI6uTOik8a4+8Koo/ULaDtw7N
dlclWKy5EnxI9vmC0KMvp6Tur10viwg/BtnuEqFc2CEoYgvw9Xe0eSd9MXpKD9XC
WtOd5rJu/SjT77B96Sf7MsfRau8f5ihoJaN1KiZCwovmcruMTaOQFG8TokA36Tj8
9eLcWZIqhIeP1JmdRqQ6LHMWNdzjV6Rs5nUYMP6lqezNAIyJh+bSpnglvp1peGwj
gzWrlXUbdSCzvdr+63go+HFks2moA04bn0Zi7kO9vTkz3MzAnvasT+l1lhjwbFxI
iGpmy409z/udl/WlaHAiLlJ2x2YjKNMUL+qD2tkv6kpeyq8CgF86b5xTJg21KeQ1
puxEZ/tKP1CJ2Tmehc4jQ5+oBxMN4IPde/GT8X22v8MmgaS8na7p96vcVQJydCGr
8WJQZd3ikZV1ny/HGaDsJZLGHFMPpQbgKRWkOKsVuU/cppMLOs5jnElbVXa+cSDY
OVmbCwBBgGAi24RMQo5Bm4BhEMgixyQqfg+e1CRSGiHcTdLsw3T8Eur2VQLl/o+L
l2Uhpjbkeimi3K1Xw70/2XYWn0cemYDTkCdxKB4gcT2OLqaLyZzdtxFExFV3ugP4
ST5sv+tWGglCBUS3hMefYY42hwog6vxe8KIZPYZmF15xYsS8LoW4C2nZlHizWj0B
dXsIBF93m5s5igaEvY98Az1/m/DDFaF5kRKMpW6Zt5/Nme7jDRwOE01fgue9X9qA
P+WTgOyWuS35iGNJhwO4YFY7aMqDlVT80GX3RWAco0bL2DAmmni0gkq/29mJAnfA
+yO4i5NZSl4e6xoZOh5GVDS5lR1D/+9V/ZW0NAfI+tyD9pJnN6TAwmpWJj6iXTF2
XO/BzBCgW0AezNaHyh8aPFdSZP4fsiiC7zdofTH8/hqZQVePGs8eIFp4x7hsbQHz
fcc32oo/hKzduofOy/p44GaHGG1+an4SHURzfde7YnRQsnRKr8ZezRGH4DodbxxX
sVWSvfmEarS+ir0wRnHleTAK0GbTlUUYdR+Vl39Q81QWVEl2KWwF7pNkVXtiNf+U
9iNmi30Uj/vhT5rhErUfOCZPTcqvsKFDk7HkEM4c+SauAq+uw2uUq7vbdowNPcrb
E/92Srilbh29YFmzztCfaBzdhLYCaja5oRm5hh+iEzOQG9ihXNd17pGUUOx2ODOL
1H4sLszVzFyAGHg9cRvZIZs7Eoe/0VXzt4Tj/Vc1GxRjSgyM5us4xHgmDdr5wWIn
lpIVzM/2d50LS2+tWq9qXY3CNb/LNTXC9l3WpjtnLNePy3JvtbRE/xd/m03snohY
UKlVU63TkN7bqFsoNfSwcqa2et4+CtAvtK7xZ220S1YvtFHq04q15BSuEqRts+c6
FH9xYdlda5EPRQuKCmaZl8Awxhyn3RpU1l20X9R9+kUfVi/4WZYRklgPH2vlmzVK
xOJQbbgbXwGWbkMdtmLXZH5LE+aYThR6aEy/9jgxtGgoHzOXU8RagaRFkdkCDTxm
dgGKW7YFGxlLgmywqFV+f8vF7SptZECdEaZIHleTh1JhbS1HQiKgL5WwS6tAq0H0
k6tIE927KEllOA1zPtIueM95mp8HZ+Rc/kv414iMMgoZq9oebBJa+jJFuHLoVHT0
8fCVkV3jjtxr3J5zkjNlGN6QOWaO4ITf/wI02MmTWl1+lubl/B/oqjdG8RokDiXb
iddSgSVGcZhE7jWR5Ey02dny8mxlxlWEIvryqwwQ++LoPyM+P0JcoFV9EnpN4PwW
9nAqzPN6q/gwj4BKFFxA/VPNJ58l9jg1SMffkETj2f8NdFObEGQQZHcMjlNOcAzR
X+y5f4Qhj1Iwk1iKWExbTehQkorMd1c90awKX3UWEwBDk5EkLaNXYs+Oh4CN8+HM
DInDqiLc5r/mYYJzTTQSkD2KRCuH/24g+NCM5hgp1q3hkSBwIZgCw3IBXZV6sd0d
X7XgpZcELhc00DD9aIaABXAFnYuGmCql+Bm6mTt86K3ff1wF3nZLq16eKIYlssPW
9RLx6+cRR9YKptsHCQ477ICxeNmsIT1mulb+ljr8qdAHGaKT+JqFArvJrPF7lrhy
yyqxNXDJOO2x2rOj9STKSY5x8h+/cN4d/jDG6hawpkPNfQUq0yayF+Untwl1en34
anp6y300e2ZpZTGRmLV+1UEc/9n6vBo5owayWydIos6SR8ia5qFWjK9BD0IqF8Ey
d7g/nrQ0tampsL8zPWJuIDMKysSCvYVhigWF3NXBWTmKIV9c8+zir7fsfsD1bqSU
Zpvx3s5UFbgus0exgrROJnej0nRmqDqvrLNpdd9aNCNH0+jU+Op2FMLb2B6Htz40
XRGO2gU8lsGr5ci9dZsn97E0i0V16PI9KdFYA8WmBNqIwdSGUiRjIS59fFU4NXER
+2ty6we0ncd8jAfzvcT+EeqjKEVRue3zdSvvL/PxLR2dusvB8rfzHd6NI+yNSA2F
lwpxwjPnNPSwxIgqho/QkkB/6Fo8rBFvycKSRqNSXyVJSRhYrbNK6irHt1zDXr77
2GvE9PKM4fmCk1tPKAr0OUz+QI6yLaMNANIQm5o2qHWw/iT60uM4iSycJ6NzK0K3
DofF/r/YobBmfQkSLemcCu4c0bjUm8os2X2AEldUhZe+GiU8o1y4NRNilIfXHViy
ozKUJxeKgUBTKDoUZ0ElwqqdcgEBt8i1CMzeSrFUmygQrBS5XjSFkjvr2YwoCFhc
5x/OEzKWyC+3g1iqT3ffQrk2xerh+E1ElfAAW/LUXGzZrNcIElOsYVh7AhOpqyWW
DcWTY/5mu3nsRrNzexocHzwCuq2Y7W+FgN+5NOtBuVvJKgeVtvOpLNA/TI7NgMHJ
BskO3PHfIUTh5G4VQyY6aq4N93d5h8aCtYL/WbMx++HdLO6SsvMc3v65/Aor4c0v
tykKt9Y+/h8CUk3VciKCt4i2q7dUWydSL+tl6Sha2xjPY7eSplUEy2mEAwPxhrBV
9Xq2hqBZyhqyxj0QsAbINGDZpnwDg4e94IkWtAp0+XC7bsMGkGKoGuJ+EdDzRiiy
sajPnby3mDA+kC5VG0sYsrVuRhx7eF6xvpcoPxgq5Mq5UFJreFcw8C3opZWe6Rc7
EV6OTBzya14rnCAUAjwNXMMYCpnpmtLrTPZ8Z6c5k/D77hmg81inyihj8dhI0AZT
3zHyzthrQxx/GSem0lX8OgnA75G9mPRxc9XjonaBdrPxxk0MainTMQ+gktWxJadh
4FNJ3xLMbUOAPJteBbWQl57MbqlA2bu3mTKH//Jk6c3hgGztRFza3VXUhFVeTb2N
5wbPbsCIJLbME0fIhDWHW0dhwDDhcjbIchy5YjxsFk96iOe/IERvjZjlDagAZTJ2
fD6umwEh7WVy9BVGKiThitcHNIU4doPacCGSLFHxOGm3+hEmfY2DFOWm4yXkVdBI
uSOdnkCsj/50MBFWb2WsppfT3hUYfc2GD8qHbjqeCWHgejESGCkLW8wALudq+Mur
FnUNsRHYmXK+RLpKwMaWOPC/3yxK6Xona8gNA0Ry10/ouZ7LhGAGwe2E0CU4XSbZ
v/1IBEf1pHEqN6NY9igg7xRfGM42eCcWVf6+AOrnELg/gfp8tm5SO33V1HqfvBWZ
`protect END_PROTECTED
