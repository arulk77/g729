`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJBO49t/2duoG2xKXUeZ/AHo3fw5mB3mOaMRVKR+BLGs
E3dMXNr5jnAW0OgsMwbHdg/gkpubqipIgDXF8TlpAuYGHRtUKbeO0kPZF2mbIl41
F7BlL8q8tSkgB14pdbBv/KKBeieHWNa97UZVWfmfIwm14xxr5qH/CtVjWUFssF7w
SgEzdzB9KWCq1QeWWnZL44aoKKsqk2ZX+bV+FLwwviRakbBjpirprDAZMtnXldeC
`protect END_PROTECTED
