`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNxBtb+uWdCYXAF05g5tAG9C5N6cgav4M/uObxZm0OafH
vg+z97c4tBEQ4hdXWgJPewq/7slhuGWSgwHqaSZDUZvSzHWHnBm2aCeRaCKYJSmy
lUoBrHHulLHw9aYL0Cv9PD3adOzhrMnsFOCtYVnGHlLaF6RAgwbJW/4IPEeZNqYn
4t42gn4rMkyfyWWkq1UVedJxbTAJHyNbJMDwtiVKVfd4az34u/OQuAUaL88WJfxS
yiYSd2TEEjYJ843UG6rdxa3MyIUe5zoI971nwDgyUYaWbXN2pGw6lXliMyVqY6x6
MdNk2azT8BD+qAIKcwyWViJU+XRR8uH9n+kvjYvLRQEvdkE4H8m1ubQjPG8ancQU
rq5PN569pSqcbJ9yK5YZ43L2qQyup1cD9wg59NCNcL9/ckWb1d9OL8uMO5rod6Ls
gEd6ss9uhiQc0JHn6fW6IFP4ObDuHzqpMtKVjtc2Tp8ChRAeOFod6WlKYgQGelm0
Fmp7cTDlSytA1Ru9eHsybStXsaxdK4hkFesnY9YaX55NjDMC+sucfFIXVLNxey6I
lgnvK5Dc6GynvKXH3LJXj5iVFWFaoZu4vcBJSZTbG92OuAgwHGVZKS8n/RTgdff7
kSWa+Dz/ISCUYSpW5M3Gsp4YHgkTrgXlsVLyx1KjTomps7XhB2PWvCqM8h7WN9UT
qWMFvYhlnm+JRsr0VSHFM32ckeKYOz1V165ybR7Not2hRFzdznguNHejZCHEh1jC
2wuH18jBvXgUQMJaLRmhczDYvWAULzkBUg4iFyN6HD68OFdxp/fYwzP47yv4wtXg
5Zq9B3TMRlta2aCIOwUSbyAp4OwgdMwxFysiScE8SeNZd7Ddl6lK2+XWtSN0fWaN
NmvskVa4PSnvTJo7eL00sR31r6UbavEhsWQ8cUEC47AJFW7VosW1ZsfqjajSkJVT
Jbnhh75raEr3G0m/GkCtnKuZ7pSCjThQJ59VWJagKxrNYX1LyU1IoF3xihEc+7i7
4kW8eu/W61JQUBQ4MzcxOcNXFZ2LAkezjaxx5ZdVTnk5dCv5VdKAZ95QmIODWqZ6
68h4Q8Vu08yikO8VQ3jL0+I2EPSPLEbO98HeOcwqzm5Opb5+KN0qewVLmubvbjNv
wDEYxiY6aPUDFfjMQBffSUMEUfKj+3cKC1hIkkbF/PZOCxvsPHgOBbXslyfO3O6F
GPjuWXkz8cAh5yzjdwL0knF9y8VVpfPtB/76gp1IuFi4PHJdhvLkaXzO/Fpp1Jzu
L1jAci1TAptv4n5ktRzHusPfOwpapdcHKQen2ugOuSDPwxg0qoqfOb2iBw2HHC9h
MT4QJTguNInetJPlJs1Z/UnvHlSERvZeF1ibXjxmx+eBFsQE1rmRrp77Pf8xtN4u
SiemrAp9UjyFxRpgEsz1zvqMKumdmKgpvCaSJaoOj/Y2LD+sqqJNpzvkHKT7nm4X
pbgXMpz756L5f7h+WQ5whCqLvWXMDN+GNx5QuoF1PyW5+as5sk7byttVy36B/FSc
XR29goXCJSkxs0tXIcJZiBwWDzoHslAzLO7tnfgDBRZ6io0U0cTfLKGi58zynsnh
4hM/Nq4fapgM5Hw9+azFUvcrb4d0XOUPYxQgTC4IocZuAgnYyazdv1VYolZIXygA
ILY7CIM5hpU8ZJRsRsdUDPCDGbJvmXlD31722YVZbb+i9VGvl1zIQTTIdTdylyb/
LvUZGXru3uBL/w0R2Acia5B4pEEaDHx2UrwFojBvrdM/wAasxl8UWNmTSdGcVwXD
B6slLzQeDWxSDX9aQg0feSrFHBapJmSQJwTVXIWeJS5aPnxwGDJ9a8sh92mPU7B2
Q0xcrNKGG1V6AVSJJcsNVkkTg6Cf3OvPh2AskqC9My5W6fvON+NeQkTXIeb4XNj7
rxX7y2bnKifoHpG8fBiTSzZ8AMtyAS4v1FBq2283ee1Qx8o6ImGq1+Hx4DmTIfyN
Jo8xd4lnLxv7CK4ao1ctMneIB8Z9BFOxMszMowHwTAqm0HFs8RmzWM++6TLsMr+P
gs+nSU5ZE6eitz2eq7wXgZpg7HIzMvs6n32g91xqn48YUrCt0vFLgYo9IxidqKfH
qjwcuZQzgiV7xXuhWOsUMELzzEWQGh8joohpLOMNLl87OmL8U64tL1Dp0xxe6VHu
luQUBv1n8IIRw6Prxb0abCqB6dH/s2mV7KUWlTMQyef5HVdAQTIS+iveoPiIFG5j
Cka93nTvfAvtKVqF//+y4p23C0MODUXDhqgzqVucUEI3fnXEOCCvn6SPomy7NCDT
DFEqJy8V6R6niweVo995RInRMIqzcXAhjyf8d2yns+f4pt1uigd4AqC0UDbsHhLg
2LAeS+GjlS5YyWA2FDHym+9twEdtug7IC74IUjVoQGwm6+jlmnLqcA+MML/gU2Yo
xTdfq9Q7Zjip02ZcUmh2D0sFJryWjn0Y0XYvM8fxvURuUkMztDm3+b4KxjdY9Etl
Z+QhEBmeNuff0q4Syo5tkudUSpmjztqn4xsRQDrxjJihhkhk3mAzUiIlCa4MHsza
BeAS6A7REYtXF51XYISapjcFxWh/gb3/g+CKl8lG56schRHa/+jyWik+RIdXTYlO
AAFHoHk9TXbqZc1ueOMzZRy6m/tJH+NGD+DjxPLmfdxk90wwiyn+VATJ6oqblQkq
g8JLL6ropgz+CmJBc650q04fUPi7BZ9wq4Bx9htVLMiscq43oC3urHjURgpJFJ/O
HFxyTRTh0KXBsFZedW9nWQC6hBqBHw7MmrSP8g4Uj2Q4KYXPd6dv56v5gUHHpgVK
uMP1Ow08ZIB2cpBFWAlwSiosgm6pTEy9g00ooqYyGRMMzfBN/MEJI8uZLy6vWTM0
RKWtp93PPGKONIcmcG2C5alOMX3ZAaeEfdFDipYEO7eNxRHsZtI904gPwAXg/2Id
8WzMYbiclWnN71m27ivx1Xnb++gOZw2a7XTcBqS4Koq9od/3VL+k0EGeNhLO5U6f
5d2Fruk6+VKn4lYi3vjRk33BvWDY7VPJF3i3aqmOSpCMgJoAymhbVym7OGONja6m
eSIUUfLlr+UpnE+MV3GjpHC0xcmoFuniHOu3gavkshoqJ6dMhE+3sG4DmBiqr+Pq
`protect END_PROTECTED
