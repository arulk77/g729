`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGIZq41k16igKj1y+U8FgqDGW/ev1I8hGncys0bMSDXN
HSKfHzyS628XrPL7iyCQDvrjURb/ZbzBEba3+04yGk7oVMg8oFrYEV3oUqJCkdo6
z1UnVfzMkEyqvD7NRHKuc8O3vWBp23CEFXxrfwwBX8GFtD8eqnYTpi0ubzIPWAzI
0TJ/RdVFy16MBF6qyLFHTdcindqfHiEhxDGTELHZ8BGDlTix96kC4R9KlKr2iDr9
`protect END_PROTECTED
