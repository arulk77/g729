`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
V3yNEgI5jsjveH7laAmP/rtu7rAKRMugOcuBALIeFctnzMcraAxVhkfQfCZUxKRU
g3YFPzwsLjAc9jmiaJN+kQJZCQLTZtVMag0n+naRhnmkfCB2NJEdZ1GdZraXzbpL
SuXgcguiZ3oVTSgExbOQwAj9MnSv2GXwLAO+a0432T23FoC/r0wSBgOiclPSRfXo
QIRdiiqLiFZdnr7lKrw+aNVpFU3x7FlGn/o/18wK7bmNmLFAHJ3NGtKn/ktPHSye
gPXtOGWM8n/DY/iPYy5aRPKZ0SC0VDbL44e5Tm8bm7E+3J1oUfLBNNrB+OHigIet
tGCapZdrC+KnU3xMZU9/fza3labKM4BgIoNoWWfaNYY=
`protect END_PROTECTED
