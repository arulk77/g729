`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
hopz/UeX2LidUfB2bbQ8IXl6qLfFS3rceLjgHVgUA3Cu13bV0iUSXhhE1Fmh/mjW
2oJ3v4dgWoclJLkULWR0C1lJlmSUD5awdBc0C/uyJAXUqNEtiGO3Q/gk5Mrta+Io
CFh/3xDqjj9iEvPy98ka3Uo0KRE2811K4bj1VqtZT/5Nslo7LbDoQMGwOgWdd90l
bqdW8lihAzGGks8M1oaA6IjG/H5hfd0HKHs2s83p12u51Yt6sRNUm1fXFC1CfnJo
PqBN/vaLrIPgAopBwOV5mbzEOijrKKCbuIfnRVjx2wCpBKXWfrpPivcoDcAizP0f
HNwrMD0j0tDGdmUrvRbYj/HWeQOiGPtizsMX1XAMhkVN+U7NI0UmrlP6II7wjD+E
qyVojozLNd6BQeh/0u2kdcDKqs//8yc/rti7fREeYO70YYetuG11Mh0rvGRkziZJ
153At77HpV/g4sCMOkDYuHwt3J5LLXFOn0crKu2d9zQarG4DOM0cJDoj0KYLX824
sjdqiaAWSrHsB5EEdZrOR6iTJUpzgzUwjmWSIxo4HWypt9QeBVbHuWViqE953N2U
SRoTJbZ4e5G8SRk6hJX2Q28DZzbP7r6Mkbkm8BNood+ptvwVPPc1w5xtY3JTVDBl
NiOEG6HiQKKapl3PFKGnq0cHQH/j8+QiQUNPzM7S4TD5c9l9AMNEk4VTXVf3EuvQ
SO8GIqXLUS4b8tHo/wSYSKktpuzfRDezJkjpnNV3TgIVWEP7BvxH3M7Fsg+DOq4G
1oRG123wNVST2YodCzc5LcVspthLENAPC3+tG8o6yD3Kng1HEN1lVeq3Zz++j9N8
zN3B8z4O5UN735IcgZUJjiTtoPV+8EnNdHSRpvhnqHW5DfaDqWQoBqOgVXYn7dmg
AQwkKYXen5lLr4+2cKA/oR1/VhNhuTGi98fEAFXTmZdvqHWPVRHhBuEuB0pItv+f
bzjrS6RVxV8kf0HKGZ+PaW4+vhqQyowsuOXxVCYX3MxPuBbA9aJjgXcjYW6+faRY
isrOdF+J3M+/OWVBNhKLBlO7mz1+NT8NyPEWiD0i739d27juXBxbNYBDOkKFaw8+
tYUog8lhOXVDTR2F99X6MEs5EgbX6g7Yj7C1ldhp3Gl/MIkldF7p953q/zxQsAs2
ROoe/ijVtEMlnH/bI2gHLYuCkEwWf+llaHt9fg9JTQBnYmIOiPcolGLY7pTOPWiX
iuArfj4TXeHGJHF8NsJq5G51ab9/uCXaNqYHr7fw28STuOPKKdvqqEfDRK0iBCNr
ZMYj9ZiU6XiBtMzh7g/ioakSghzpCfXvSpPdCFwuakKOFc+KWSu4Amfo/vwpXINB
ehBDb4kSju1Gy2dtUSnwn0yMBy+Z7GofRdK66VOs0oWrZoS4jZDqF0tWojCGnMpT
52NchUPKHhbZ7cFVbjCQcBWxeqBdipHUGRBsSREaGw7RHZhwT/oNl8I7541EQPfv
T0UJJOP986C5vXP5ihOaObEbSisTdBwOS8tAFstsBIsfVlzKyukAWPjrBNBC6gTw
z+bhDHz+s+NOuTSH5WAgJ61ghRJ3qSioBXg1YMIjMXpwQGZyLnvp2OaNtaNhK0kM
5DQC65iMhzbv7/Emn+G8pJ2/URMalHbjQ8aWO+QmddLhvP63jrmlAPd81gtdKRJR
Jecf60C9fPmLUA3UMGFfjPVNpD0g91JJdgJ0KoqQsRtJyqkoYmLrQ13qfbCLgCzX
M7BIQ8V7j80jVcAky+n1wVbpRifo6elJVqyoKuXG6pJN7gHy2IW5N/ZOHZWD3lbb
3YlLtRVSwD8qsTwYTxxwo1qjhc7jyFZbmlTKfydgA4e6C3NHA8cPGboCumVEkMv7
t5Y2DCPxFGQbS0OGjPg0NsrD8g8awzTPrYFx4xFST0CHqGUu8hZTsSEYKn0e4gxP
SoZWOwt+Q/sqyHu4627uSKXKkmPoX1hSsL/1wnU5I4R/N6DAhUURTti4MiXtYLaz
hYttPU93fAKUs3e1yjXS2Rvw/tc9xd7BT/eMZeF5xQC4mnPj9KGwwnzrEx6PRVjK
T6YgN61CZ4kDhqZZu8Uc5LxRyfv+Ro26ujvskAO5nzlzt3KmVHrM24WIj1SBIcKz
i3qykn/+noy2jeZm524yseZV+Pzylzke4VAfM/8TRWlx7gOZVMjqOR6zyjRZ5kOM
oMsHkCy3+FpD3fQm9VPmERJKbf/xQonanIQlW3DXy3xfhu6HhA1H+JVt6IM7pxI6
dpK0/i//QlqCKi+xNBwtT008PPEGjvIIaVkJacLEgpyXag5D42YdmwcQ8+tVISWH
NGQqygxs8q/JmGqx0cP1IpIEinYc/quXFwBJNN41iIqmpGyYBavmoUCerIUU5F2h
capoeGRBjZkueTJqfHkNzndoq08KW0RFJBqLBZ6O0PmRoRz9H7VkPqOgLgk6U1u0
aSIeFDJqra0kN9g1IkIA6fC7jTCCIcSWlSj7/yvo0BcCaHGGJsi3w7wGhR8pJ8Zs
bO60bbJh0GQAU3+O1fV8YRUxiRMygkHhQfIIXNrEBrOqw8gvGws/9CM5CLTUa0Ti
RWWT2MyPAryfDjNoZ9X1qCNiSXkvQ/fpMXdCAlSQWs2N48XR48ck7wkg5+NWs3Et
DmXaVn2wl/gRuZ81Wb1sy1+BkhiJD1xINA/79xUEmk1o8l9eN0K1NzLd3MxTkouO
tCUAON3Uy6TBHR/0K9Hp/lS9wLd0WXHEQI/a134pzdaiCKOWwhrNVfUcK4M0Q3ot
XmKm8E/NQ55/NCNVrzHlLvChNsOgYGFW+PROLy0NZ0NEyUQCqjuebYZPemDma2I1
fs/jQ7FaIndYrQSnjMHQhFVd5NdmhBzGGpYMgfqOXvQKZ9mWu0swYFFJh1J0DM9B
h5K2SA3mMaf+d1pmBSUW1mFr2SRLEQb+HVp5Hx94HEexC0piusm1uTg3uIDaVkKv
9lrT8pixzzRm/NUg46OwC7rTUqLNlx/y9WL0lETLiQPP/lzcWGrOXoG7vhNhlZeY
ULBQc8Jhlh0p16AfuZplkJSw6gmSMQHVAGcgwe0xBGUUvCZO6a300pI3lZ7sIdhH
kbSWqNNSQsaB6uYTQbJwRn/ltifd6+yfYHF02BEYN90xYCJfHr6JNEO0dXJHSZmA
o4wy2KirB/pkF2O0xW9AUlh2Kde9IOGivdVNe+XS91hBSKX77dV5CY5veUqST6Gj
SiTmpCWhsl56oHJN1zwbZA==
`protect END_PROTECTED
