`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1adScbN3IsSrhpSu9GOkI1QV5IAtN8TEvRMWB5TvonK1A
/xNiDbRV0jwMIvKpQVG7zrw6uEn8bfs5l4Ig3XGJaC196zrf7dDnr2rfIBdg7loa
E+iUNrPR4zC4AB3ujYdpxV4SeYjXnID5VVQ48yBhaWGPYwLc/3VS2/Wara5Rrs0v
4UxFIyopz7f4zgjypCmQBXf9Cwrb7iAbz43gg3lfoR3/C7r3TD8Z7Ehr9/zlWFjk
K7YdOAo5Ej4z7YLMNYh2i6+KZn6MSP8AU5UONnz2LW199oylkJPHnD8MaPstQLsb
D8VK1CqUnoXV5sMRnZeDwcUlZCzHDfEu/jP3fG1eQxVFuDQvxAbGWx0wsKSvwEiu
r6lcP7dW8WyYzmefgQIPnm7XhnPpUB0rhxExE64s5ZKb/HJT9I6Fi6hR1HDvDSGk
595M8DTvQOTPGonRbWryQInGFx5gpYkTRTpbRHtEkAAYXUfZdRVFxHxW0YprREET
Oaae5zGwXdfyO0iphzREVcMtdqo77NCS24x74Ox0H4ykHvhmZspFxPHU5kDIFVYt
LDOUT6o8qoP5ASRID6LGnqb71gu/IOSNATG6PJW7sTbu6qVco2QnzIP1vxTS/U4d
t27HFUdIt8C0uOVh0BjDDyek1/ws2/v5BmLQI7E/Ho5qyGdHtGKKI4qDZAseDLEs
qbPfUUDxYetPi+UogLFV6L+mAsMOG0vxO1uvE1T36+Fki4jFg9GcN8PRYmRdmwwZ
7EQt8gnDrHTOc8w1mZEcyV0y+dciRcQYUInJnEa89MQKs8A+cTNvOug1Z9LROuen
ksZtwb9U97D/RVeiyi8GIH5umBu8rEA9fJ1W9BXVD+2U+NGJgl52dUlZpI090Fvo
bKgmQDm8maN5C7KjZwQXvh79NSZh90nmprt6j+kW3s6TsyCWivDF4TkHBkGz3d1U
RRYEUqY22Tm/91pf9RMTrMV8D5QilJqSNuZ6zApl1CKEaKAb0hG9lt2TQtoYY6Fw
bpHccdxmUW6UbtXHH+Z/P+WY7LElfVdko2bbCJjAx9pSJ4vJgREe4txTBXBCeEib
rE6mMAZejRVHj1XIk8HdB3lzT8NBUwsWmqpHhVYhYjYIvLUuVtvPoZVXC8IRYgEg
3ehb2B9lZvfWuwwS7FN9ZhgfOZePWK9LS2/YwxfHaWTPvDWZZhVfHGf1fFa2M6LW
UXwHJjd6gJPbm3B/EBf/NQkDqitFJ6stQfB7ca4QX/g1m+xygpvSA8nXn6ADUXk8
/YDV1npcqwbhTVxiDcpbvW+/owrS6LpY2P3kHZHVPFx9QSRrAIcrZEPuF3bs6puB
NimkXJEd7XwTUTL6Mx70heCiDVm6KD/Wt40FfBLAyfHoYJxtGKrLJleYsZ+8taM4
N4Acl4hJdwuJoxqi7VkEs3Kvk17eH02ztcnnO/tUg91svUco4JPGC8tMK3rZdNzg
kYv5rn42zc7P//GrUVni0B2i7f1O+lPl8+dxfmZo0/zmwcJsGHcQh6LYsxMyozkc
8rRn/yYYgsIZntTCYtXUSjRZ4MfG0GsCs7TXK46mXCwI+yNKkENyuLg1Gpr1C15o
Ve5H0N33TbpiL7d3/7QhDChYQewHUa3fHMx5w+wHlofSgefdCE1pm9SKaa4RGD5f
dOAr3BV7qieNyGl57xcEDjuNzBPK+3Lq7PcOwaTI8MPvmln446WAO8uKa8DqnLej
zCRanOvm/ZZUGVJ27mQbGSy+IwtaOfUwVyqi/TOYjAOtAzEA7dyT1JrrTQN6NKGQ
MHt98bEzWQ4cA2qFnqzuEr9bim7uamgXGUdd4E0Jhdmj4qAOxS1L9ujO+xIBoDVW
P0Xdx20r7sMyqxQ2oHBDCbEnWoYo1/HD4P5GOfAKp/Ytmk7gD/1lRyxiLfnXO2nC
14CWXPo0z7QJHA1GMWpPbSF1qxJM/dACB5sO+LHPobB2Rkax90QFQPHDg08TcQ6M
OpN+EitfNTnlfirzCSBoMU2dQF96AdCpB4UDpQDSv6QRT70iaft6v/TdXGOw6PiW
AaGXA2UrCCuR51+gCPRU/1xq6lHRrKT9F1iSQ5oMfQWH86xscVPSQ/GOII/92GQR
JKYhZOaQDuMIZf0T7ZIrioLWImq/CeDgk4M7PGhCHXe2HorytPgSIZRDis8MAjD6
sJBfOGpgEIn5PyVB7LRjjSUlocFb7jse5lALdqieRyuGHYCkNVvRdMw6uA/PFVjX
mcUciH8nqLJAwXScJE4T2nNvDlLqSUi/b+zdUMldPAe+pkBzMs6iaT8hoh1Vs8Uy
AibnMXuXy4hg9U29fcT0IS9XWx5Qqa+ZcUPk+4e1oVEq5pXVG0SPfkmU7cdR8azg
Nxdcg8bJJLtkDCCQ2qq94EmDjYRI497jRGglJ7K63xa4eKfGynG8wTFXrHCfaK8P
KBoATpqXOkCXN3w7Cb18m5A3j0HpxaARivuoYJnCUizq3VCm0JazYB3OHk5UDVqx
cIF1SsNlJcl8A5BIQOnTUeWxDiha7fqslrqjJbY/c9BTV2fRtDCibwz5gAyFzU/B
SAOzRU3r2h4qkzhxtadJ4pMj3x4hYvqwQwy1LUqTvzi6kkMpWTfGWW8ENmucacWq
U74gOid1rnhhnWcOjTDW40+GJ3uEzN4ClZ6NEWNwJHfobAVVMopUX9OgQ+nFbTYQ
+WDgzkY8KJi2+SwZv2SIZCy+YKPsFXU69sK7Ajlx0XE6jhwdsHuWTBFka3+QSrMr
FtShWtjnLTCtE4QNhiEnrlmxBatumInxLjHP5acOllvZr47bDl/Hv2/C43O70NZT
YjrNCl618i8RNn2TNKKgcSDItAjlNrkQz5pGcux6wLZivmmRIOnnnPI2/BLUDIrD
pYDXuwyIJPUGv9OdPurLxoGSPcyKDKiqC4msqMFHpOmW2yOcKqjyMZT8U4/bvczk
kHwg/Bp+HnMpQeCPyjHGgKqk8OUQ3znRpM/hUAdluz/JedFeOzd5Oxrvoj40rrME
n9JD3UzReeCrAZrafID+UmfpFAc8ITV+Wudxw7SeqiLINaIeeuU+Pba/3e61/i6z
6sqNWQW+rbxwG6T1Ulw0dBjeBHTGhqlEejsEO7B+C0/dufmjGyTKgXJsUlqJNwny
uAbFL3O2Jnjhqi2QJKjHPTbFioQfNQhAXsK8YucDdhSj3S6YsUe5Z6ujgpKqWo9h
w5KRdNd60c1hikc3uFMX1mofgEqZYQy8JSR/LzSni94qGiTp5fGhJr2eANd2Otsv
Fs0cpDKFYqUfsGomg1I9ZjY56+olsWFQ9E9WDI7xHZFGkXF8kgJL2KO6uqFBymPm
bA+0sKvj4teEcPa0cbr6xxinqHvSVfpPNmB8J2ZEYnV4OOjchCroJGOy+gN1FAf4
urowchd569r6E8fyUZSRCakhcWh1htiX9ebRlGQXZBY9E4oyCgMcEkAbwSUKZbFq
f5NpE8YdTeN4nph2/RZAOw4URFuhTxIoLihr4sovVv25PtKdti8NwxKJ4i0cFY4U
uDOKhVTj2SoMB+T4D1xS2ssnvlW6n3lAlwXQ73p2jIAj20NM8Cyb34fEmQ8bCpVI
X2u4sy7ujlEA0FhhFtVmB3qbh/2lA6fjrEdb+za7tfP9R5zdTTJWp+yuwLemZCoM
BL8TS7n3hlsz5BSptovKtDDwbmE1bTn3Qt5GifKOlBEpesczYF5GagBCfQyi/ftH
tBl6Dd1JwOvzIF1bm5p7jGjy1B9yOPUt0VhBkcX7AUiU6RhndCLcpzB0IYYyHdAr
tPUmVoiQ/KUSo5gLvq3LSpirvLRYAot6hns8KENID16gNEeorsxEAubY/3fWqhWG
mkgvtHIA9fvdP5/ohiWFOJcEVXsIrYrlKgiao0OMdwc4AReav2/fvJSXQm+y4S2v
LXlcvfXubp/86Nl+H6P6UE4/eZ23gaU5LatovSbqZc8GsUSv9lZwkoTfP1Vhx07O
QQNfsTccs0nIxIDPiS4yfIpfKnJzpbQ3Bar89teHPG1m+LidXivt0HqXww/bKQzN
Y6sZbif3e8cC4yNJux31NYXl/xz7rEUwo3BVaZX/rkE7WBNp+YBFgeK1o6vhDeLy
L4Tal5ZeUNInk8Jvjl+ZlojYvlMUTdMvfny2O0So+cBbZDiAtltSRLBWqXkKiXMq
300+6wN8rrXgoLUVBV/nF9nl8zHpCcdbw3PUA2ola9n2G1IQjT5Idg0BKMxkZoxY
tMusKjT8H9VO5CExK0Ggx2fgTj4jbAkLvmDZFxxYgsR6MiG0dRJUEQAEwKcrHWZ6
o/M0oKGkxpv4FI4IqQ1v9ocAB3PaSwI5s0Fb3qpRVsT/jC3+5u3CO+vXDJ5/9XAY
m6EDMr+qtXGQn+lbMl39TteARz5a8FXp9lS8ALaLBERfGWAvd3M5vQ9Du5ZG8R3H
nkAU4WE35WbtcgX6q9gDtQJertqQKlCJfmndkxd6npwm7m+lOID/dwhY4lmrr7MN
7Mal8WTvkOuIzQhLzog/swZmnEmMSlI26gtSMUgVBRxspvHQbqdWePUty7d5WX9m
vYsNYHED8bckUEqmK+PLm2OoUHNx3rubSrpIHm9H0Iij9pGtqYC2MXezm6NLmOuZ
rWOfTWh92ze6M9XNLc+XZPZ3+vtA7NHlW3BAIa25mhpJm4K2C7mVxvSOHFbPp1nk
JRGaK7RJ7Px7yOmdkJ5xywViHf5c9ZhsVDdD/FUiGezSyDGjRLT6gdyoFBYTee8R
+DQkygexi86WMsLk+hRPa7EyTM7InIRJeZGjdJN21tHMG/O9vFQ2kgfgBQ0pOcw8
qR//nVH3f8d1GxSGYot3tY3AanB6zXa8BOGLa3lIsAUTfO8QIRKlT8Tey5zTTWVZ
bZYPNXM0Ja5LRQzn/Ea940xkAeif4yIW7FSixMTP0Nr233er4Qyz5CfBOSS9vMHJ
zW/5FGvPqw4DoRrq7xjP4fur6nr10GYmv/eELBkku5DWpr+WiAskXndTmeRpoCJO
Krf1vty8g5CRr6Qr37QDd4c8jTtFX4bMKc12xqz7AoBdceU3NOk0S/5GEXYYPRJE
yF/4XHW4HigtJyyNSdt8+xcAZO/KannfgWHUgSAxPlVGbuQMkEtf5Bm1KqZv+O2d
4CyOKI3Vcgm5NhCEhg7226qsfa8AdFOOzwflgRJM0CXxXNtkHeZU33m2PPDLpel2
4QvoEn167CBazmVoobrM3oTLSi9JRvbqGw61exjQ6z6cj2hDBmfQEokfhDV7p1nK
6hSHJEiBstoIT9gUr2cDzYh4BVLQYdtufpX3+2ObRcKwT5AxmqOj41BHvajTZq/C
TZS4WvMSs2DcCDPL86+1DRxFUvypPV0Ga6T5I0sUzWdP8gE1SDWKji7xJSiXWyDz
TgTsNcGQPvpBKjV1aDJiSuM9pC1sdQUg3cdZ4vNim0UjX8BT5LjZ/u4cJuEBmMVw
QDFWIL/vmMjGoeUQXBddCuydLoC1z1GmMg//IHTojIcCR13GXwGlNIvUNMFVlzy2
pytSoFm8uKpA4nqvt3LWoeN58e6bdV+tRxTF0Ew36/Sbri/dRxv/ACXTTdoj4t9z
WCWd7ohs+MfKL6aYbpWV16AeWyJD6THuIYVM5FCKNnzNc7gzKJL76C8SEaUTrRZM
yPy7+EVmaovC8gZYYvMj0ppcLs4O7/mPjyj+vdDAZ2BlidRlyoIfKLnIARw5taUB
EIqJ3pY+XqPeIymPDPdqBFUtRmTPyTPQOT/TXuk9DCqYwUQxkpW+vN80xo0YSVEV
MFKDMClWKOa2JPIUAy8I6kmoNYBCGEdEDVXhVEF65uLWP5Vl+6Z57enW2sSIRLly
hkmViLly5bl6F5ENZYSODeIHz76FpFWD7rZsOBKSSj6cCWVhckDhmS8pRw0Kg4YV
F8YoqNBL6vstbTPil5htH+1noj9SStw9D1VIrZAAZIZOxZR2q4Lobf0B8R81sPXv
lYL+bc2oEbOQwmDMfM+2loRReZ6hUk3PXHn5iFd1UcGfi9jTjoml9KAyLPf9vzj/
iRGPoJxetDPBnc9BZgjLcUTvDls/xX49qHuSqZVn8Ofoi/ZzhARgR5AlfQk5ArNx
GmtDrHJ/VgNFxxIO2UMFJnoHrfA2rHGTTAloEcxQ6ooeHtt6En++uTmVlRI2jBoH
/N0JlvJFzNER08vzoqfQrWu3OitTXdba9sA8+HAeKv11C6rbZJ//LtYWYTx6MKiz
mFz5z3OqihB61sjDr8bIaVWtXnDhPmVvEYtxwE3Ighir/Yw66Fd41bGfw/LnlAMo
3AmE/rKORZMGm04DIGIh6JAuTKwx+4JuXmRhxHPGuQdMsccvTEbOX6lZMQCuoj87
wkFr+ylFgLwFtHzPLqM64QKuT/AGFxWW3jnYQUW1hG31SNSIkmGupPMfTWjUmiU2
SMqir5X6V6j0PQziV2aVaSs921pIW/ijQdEwJN8H6LMaYBECKzvnH5n/3n1v4LJW
H1o6ZfmPWkuUsq1UdVLvQtB5DxiX5MjNd7twbcaUWRh9J/JZfXVNjvdMNSe3OG8t
KUIVDg9nprbDyBbwiwik62cakoF+1m16YjQs0afsxkkr9Ll+egaeYMNsz93T6Vcv
1cdlDZEgzoKWaPlp4/qnA46OjwXX58RVxrJg/nlgWx1wHA3scYL4Vvu6DudpIrba
NOg0E4m7C6/5v4DiVWeXrDM32T0juSJoeOqmzIQFKxu1foERfkg+tlqZpG/0Cu8A
6pvl32rE/w42P9eCPSasCapFsdub8DMI8rovvShDkkEOEME84ve0I1YGKlNMEuRv
FNZxh87Xli330Zglo7jefWKbrdt6XqWA06WI8XpP2m5I4m+sDco6L1q4jvZRMmYa
xFraCs8TylzsaA8sSsqDIJPnU3lfmF1vT74GmNF1xGEaYJ0LmTUKGwwz3TNKUp81
v0U3nM90wiO1flBYnNze2hd7EEsHQKzogN5SyNv6cHPvvxI+sVKr2bKTz1xZ4Z6p
BfqgaA5Xy7hh2L85XOBop4iWFDcpsjQxlkKPx/V+QlHR7+VoxYdAcCu0AsFfALxv
Kyr8G6u1qrgwoM2AbmyJfTXN9WSPQEUCbsXeYTjR4U5QW07XMuKh49rzS7OuJTwA
jQxcKuHhy5j7Ipwcxv4rXAu8vFZ1eLrtzJ2gbrkrR5zKh02uBat0oNzgpc28Z6e0
WgAX3lWIn7U7WpdwSNikXlWjra0b76Li6cj1NE9bz2I0IeYenkNTal2NIB+ZSM2t
VoYc5L5AmyE84Y8PTujB+GtT9SPXwqFMSY29Tth/DHld8CBdHtHxfEWxIpozszHR
Ano6DBkMRE3jNCM/I54+ZiqwYtXoj0JPoOT4HfZcB0TWJXy47oGGuXh+L0fFfcZo
sFHHBFNG562VJlDbd3ifNW0HOQATwG6ChWekdd+LluRTVPBmNTmYoqaYN+HHc7n7
pI7hlKc03Lfoz7xo9LKnSKFzDGZ0luAUJwvVMxhjMjYf31ARADo3H8PCEDqPbh4F
bsvsBtB9P3WUTVL5otmzbhHMgbpEI7Bt9lHx8qMdTM2Dx+//tvWuRmNfvJS5/mEi
O8vtf+/M1tNERUp0TmRy6s7Acwr5mUEAvjvQjXg66CQl8qz7v7Oi0nP2TwgsDYXy
AN3g0MargkKTnqs6xn8y58PC4dLj7H1NFA9uhpFTsiNXBjjvJZ/kv4a3w44JkX2L
tMoqI8aQasMiyZJDm7S742ILNoYE1bJ67qnMBbdSYM7n6q+C1LrShtrni6zrFhKS
MnNfThmW5cqsw99A6BP+UVgYqix/GYoYqzBsrjLHfbOX5gj6iK+yomv1MG7snqPp
hJuqYVkbzEzbaLZjotvChC1Z541VYYiIYB/E9BeaAL0arJVfVL5e5WQjo7dG9LK7
loFYbfSwQuZ1qLsjZ0u63Gh+UVkJ8VS4VTkZmnqBwYr7hY6NoUfQf/MafMCdY+5l
0WMjNnC57DAQhCwn77CfT/q67Bh9F+4q+HEM4kyfsa6K69mY11zEF4qYvVxfe50q
eMXjjLCoO5WWX+Pueo/uDfJaF6kpVR/gzjTK1hf73kKtG0Goc7AvmMbpq0ghNR/F
kZZtw7PSVtcFhAIFuV/Ua1vxp43gWTm/kHEpc4zz8peKzKygLU/l1ms1PMrr5lx+
AGm0Mun6zSWpFwssV8ytimm7h/ADP1/r5ara/33pHKrL33gm0AH/dvw4zLLqZi6+
vrM8ITjJTomVIjnCIASPJgIPahCszE6SxtAlIVqCzbtCBKXTRJ43KipmHcgjCD55
IRm9f8Hwr1yiknQPDr/7xkRtXsLnOeuqfUF3B9+rvV4UshA59iy8EmfKYiBh/SI8
0SvjMNGvDzLmdnJ/A5+NACnTLSxxruzNHexYtpdeWKg019uYoz2CKw8AkaF4G2fh
eWh0as0MOVBwfVZRr4Ip20trFxIijHi8Qio4J3W3z2ALrtwExXAU0c2mFWr+LvAv
WT4ag/M7sCqO8h4F5Mq0cz5cM4/JTNileFKcN3IywviIxuVIpyFmdtnXcp3lQ5Jd
0DJey1C8CyPZzgWL+2nwQk+hAY+v97ZVgGpeNWPe7klvUQtK64xgE2S7qoFTvafN
RMEN7e5E3xxFu7LebqHQFjEAhdRByBd6MfaEp0bERGG4DAWi4iZP8J4epmtO+HUV
/UNzSa7h5Pxw3FlA31MFKTbs9/NVSR9x0IqwYc6PXj7T9rFxmTAzQYfR91I8Iag4
v/2XrONYga3wTtN4cIrBow354EhB48WR3AkLOcjZJpbmnGjmlpl/A5ciPLGXFfjH
YHx8rFPwRPYbbfTeDmB9/FKLvnGg9giYhxWEFdsoGKewNRfRxNwaZYEp/wYBnOue
1k12f5ON516gDbXEMvKcwmC2TyOQCvq0Y6N6Q+yTAHjf5tbvGHIuSuKTaC/hAGES
nxUKqzV6qVxgZR/XtzKKzWLz7of+F4Dq27wPzS6riJzqQ7GX+7Pmk/ANO7TxxGGK
Hl5b/QSiRkkH0/1r9jC3/SB7UUF+AmwVKmmWwLLsIppsO+iEa0TFK3ETXTVwKl9s
2O6GqBrJyEE9VtsPn3ytUq5/ZXZdggB09NW5NvEu6jFskZSrvQFfdHdNQrLdyv/V
dI0fM5xNKU9m3OMiSdvPiVrBRrQ++WFE+m7HCAt9JXLevJv58SGBlF4LUlfVkXJK
Y/AqWdWYxhbv78+pti731BlJPjPekbEXnlCiGNKJBf4TBJ85UtTg2CK6WefoYoIX
FISFmLnLSAHdOgmyYT32wcNALlT44Zzhof90Qm/Hl9eHbir4I+CAmOVM1tS6cjjh
P0g09LbFWfJPwTWkQL6lGiimumCLq/qd2j02ojP4TeeRFyTA77tYwseUGL6LYDDH
VWGDLXybl1Wq5d3ZsegqBNLJXPIITMNxLNq2dgwbUBBHvZKsyngw3grNs31E9HoR
kZA3VIMXBIC3i+B+L8b/wBpIpNNYhBPlIAVQ14uGKlOiT6PQwpoELwRL5ic4b21S
5T7fIIDW0iuAFY1a374nSlPLVu2F7UETxr79QnP91iReB2GtVqybOXdc3Yhe5Jfg
Lr03xPJvpFNWcjGYiqSCLuz3bLyaR9Wjc5FHLN8YZOdFDQNW2r6dr0zuhnX/ssxA
zmnXiyDYiF3G21wrh0s599Uy7jd/+/yeJHBDxTW8+tHVxixEgbJJd7Xl3PBFWO6l
EpRxkHRyF+Vp/apBp5OCRBO07lsJaIgcIuoBBcOMXwr5XIEmQ7ZZRRtei6mYXR+W
yEYLku75RUOIFKKMpR0kvROne0EhFfg20BKex6uAjHotnbfISA8cTVuqQhf0p2WN
ULAPBxOelEyoRSZD7JjInPm18wcuKh1Z1/UdSDZg1JVeKN2Bi/VkowkUC8JcfTYJ
TVV3xXsbgnONkcGf0DKfseODN5P21f4WpF8iAZiN8bSGDuSCXwZrrPjG7lj8EZhN
LYXX7Og3Y5Nk6T9xoutn+3GwXWHJ4foZUHaVDHmxSE6Xw6sgLOvMC8rRsKGtQ56G
JFru9Sdwa5vCN9PUgt9p1vrL+Ac8MRRtx4a/ZKWhcG+wyBe7CJ8iZ9HfLLBcbIKz
cOrB4/JCxOaiMbDkUKsV/7P95MgKzbIjtZodXr4gdjYkahX61TEp6A+6BVkGF0d0
u+j9+e4ZDCottVLHVk9TszIbgDQ/D1Qjb53CjJa8XMnQHWbpt7ISwT0Jmy56pl+E
kduJtLOHrorlAmuK1TtLx7lQXOAh70PR2Ssyb6er+EZuMJWw5X8u0MommiYEn538
8oDGpYy3dRn0p+jwQ3YfoHl5dXCXxpQAbSzyQzcE+9l5zdq3seFAWY+km3kIBiaa
Ji6W6Kei6Y6mMI/FiN6ihNLk3KAipGCFvGKPux+Xg+YIELSOtsj+w4oN72vqPLjV
1V8qjmOlcC1nOqLBmnhdU5qI7wI2ebczqu1EGPoXX8BUglFM211Gh+Y7fs1hNVZ7
oJDZ1HPGny6LL3YfIc8nJf6jF+VISUS+UBSoo2I6j13YMZdm6/e+sOOnd9dBDHIZ
YtmybM3E60gpdiJ3qyGuPCKssfFxvObLw5Vp4G3ufaZwuWIXXfM3yJpFlxvzf1Wh
t91ugKv+P6wOa12V8rufqAswGbOS64683I0N+vpWeo2sOj5L9zTJelJeprEC111I
ImNeSLoQh0khLj77bnErq2vv81s3QAG/GxwR2CX51CbU502RftB29yEqkY0AzFFm
V3JrFbiJ8DCOZGsp80mCXo7JeySixRhHstXJbJj+Tn1SmaX6xnreYBGyh6kBJSsm
MIM0mrbSGLV23WRsOcytyZMmh7qtVZobNSBNoDA1UO3kMCNvImU9DntMboMj9pmh
52AOjOTuqKUGqF0qghMISEcU+ZVxkrbokVtGscF+Ie2jDFdhto4JKNFWyNc4IMEe
K1mw69RjgyXwhn+as/gPIoZYXZ22VxbJIb9Cw4g6Ex8qCaEViP+gd6D02e5g79aP
+C3Ut4ZoRErXm9N0GNheITrEnE86nY5pSMonERbnbVIwl+SOTW508CiGGRObN1dr
FDTlUzbAFozLDfXPB7wvOBFJjnttaMbZxPZEiE8Fl50dPtK6AMAEKeLme/0eJgs5
jqyPRt/VgcGUmdAwuLPTb283jTpYzdX9EndevbOfCMhILX4fdVpAHXXU0JpXxWHq
JM99OtnWFQna0/oLMOjjsETK298BSvXftDaNtJnvKPUag46BKHrvjqzV0dJ4qfE/
ANA/9B9/rYWR16Ywpcctbv1rVub46ANvqAAaK4T2KtpWSbgQG8hU9vZxV3CJCRhT
Q/+e0ISJ4JKeukpgb6jR2cn7JmtoKIiey90M0peHV9sY9IF7MCGXrKiJ0uiqRD3K
FLxaaDRF94ZYw5oCUh5x6SPZ8TBBGWKBpO3hc/yd3gyiXgvyWF6sVn+IlNReUXz2
hmwkepw28asmKY1WvioYKM6zggyOQ2g4x3Phw9zqBIvQCdN0TZ6OG6gJblxqeLLH
JPJyNJHfIk6odEq58osCnTHpWhlNGaOj/m1OFQoN7S+giuAoHuKb6hCJ92omaoRA
nsHufmKVKo0ggtBPBijnnz50JVlITWKMSdP6SBLHaRFxmqL6K3WZHzzE/wWUNZ+N
xJCvu0nJWHimpeYKpBdflIxIc3IEXHWuEjeCQRmxpjD+VYO/+jrHxv0bOqym3DHc
8SuO9ZgOv4VnzJiRagjf+HHh2EJZjaqUI2I+abt1q+eJbAWWI3utpn0S96GR8ILl
Eq+Lf8bMyg6ngS22uPpT+rNGtSaBbDeEsxH44W3gjZnvcIdLXPTq42FRlX5z822Z
RliGLTkVmS8pr4OIWd4kf1KBh6qEDL4Bhgewv32ImkKq7UppbEK150JTjvHbXdVY
VhBIW0LkcZJ9KLxNh4CCNuSDMs2WtmThBRq4iLIS5q6HdySFk3wBLBCOmkOj235F
tLYrXlgLb2x6ujpN7mwY/4maEv6PZQoRCgBnxKGTf+Xi1znlqllJxGbJocP9VoJh
Oy/WKrjkPpVB7a6m2nuqHfJk6JdGhCgnezaAfSb+aygctErcs4C47HxWIl0mydoy
99fwgRHN8Fy/QWtoctnnaUvieDvnJcBcmk9qqtYHNYJtdLt0cyCcq+c2EH2VtM1Y
9aUua8rmo+ZqlXUVMC6dIzpzrOVSC29n89jMT84KH2PlQJXQU/NuI0QLvunuf0IF
g6CsCTHDLJ/Qq1cfZgdz7dTpbFahm1RXdqRagdnCVVClvr95VRrtLxUGSO/53+qW
Xmss6xuYy6KkQtc12mLduuT214GFn5HtQXTO6a405jbjyrLhRnKDQo5qw8QokqnA
AyuUTi47Y5vEpkDsErKdT+gBDCs18r4XiIOr6aW0jV5tmEkgz7/E2AHjM+03LtYd
xAsfRH8dGh2c+9zEGqHChqyKB9rUYKoK8hUklNI9YpoegdJl1LmRGFswzxJrwth2
d6FWZyG1+c3DWtDz+rL3c9yDwpDBpHqXuKZHAY9/aZj95BLJ6frrbJtN3I8YJGa3
uEMtybMqZusaZS7X2sLsvMHfeVNInC7AkhykfvsJr7nGE/CQazo/ccWgZP44HSDW
RYC8FImmU6u+taaJgQ84Dm5TaiI7Fqq0xlI3t7i/KOkwpy7fhshUcAz/VjYwOkRZ
N/pTrO22goE23gelmPv8EyzoygOfreLxh6d8UsSvGhhmbfTrpHYJMXa7OWT7Fm15
UzN0XHkWq/BausuM+4qt/MmLKANw7wk7MxdqZ3/6KQtSwFyOx8v92AHUOenucaGg
6mhRN7q+5eldH8HzW4ZpLD5QTfMtGfoRt4x06SJnKGQioBqnUINM27wxKgnBdhGi
u10dYgGKpOjq63GR4wFwYuI5dc9HlQoUQgC/ID2q9llj43F+m+XYwWl0y86vZpCZ
cHu5toFCUxqpif1C3n8FCDEzbyU5vkkOk07ac1G4KxR4Pka3GwXN82KPfu8Pg6sz
snZcVKMbpy5anLc3p3mGTwgCotCr4XdVouFGvnpepRYlVXNcaCvOmSxUbR+dM5Fz
4fYulVLPmyYWeo4KQr5mbY2VvXH0KYaE1eVspfLJfkTy/0e//DgWSXDEB7KNwcXt
FGbn8jSb25LVNxHCPhYaUs17pbO9kk1K72cLpdEvV+hMR9aImA3q8LZ+TLkzH/9H
oqepHj0PwqYLJXheYpR5iiKbFdO39oyDEJgRRNsZKC06kzDLhofhWyFiRafB2VqJ
IpFzCWMm907CFXINWtmfFE8jsa2g/inLZgvgtfSDRgiKkCTEj0r1nHZPpK65IwdQ
dp6nMum/Uy4uX+4gs04sqIC9t4Enbmv06BJcjpdl4qOjqMdonraqXkHwtfmEPKAU
84rasVEYcGKseEeROdLGIi2eHVLF+TiA4twIeMH35n22/HJuPjLR1YhFO+RCecIT
02EfhBwuEqI4df8IgrAeJz/bPpcddL4joQaaCZHFCdSMhkpuSgapa9zrIgBRZf4b
3wqj6NnYDZI90P+aCyEoHQWuvGDA6M6DhAoOyFCbk9HIGFstaZUe1i4/dorDLM9q
pNQp2N12XsFVPj/SO4R4DeEM6LY5cmOYaAT81hHIm1aE8gOVcqqXgKbwd1zUFM/d
ybRcxucFKh05iH8spjCry1dnf29j7ig/J7eOXQPL/8ZB5uP8Uart0ZsFGRs0bX2Q
y9DwbOLpLE28X/iP1LanYdRUnmzz3IUnMCpHwbZ8zgFtu7lR3suc32MW5gyQ665t
VOGodep64IpGC9Fs8sz935ssHjzBscoaNfmh7j154ZVsKIIpGrr8Ka8a5IWEgAi1
iD1VAC8/yUIIAwsqvyYxvV0B40jKM1oIwB+6F9+dPMjmplzMM5U9sSWTQrDLtU48
xi792oDq5oP6E/9w5J1dhX2QQi35BDYIKQTiYV/v34g7so0iHXMdhx9c5X8jiu76
GFVJEc3CTt7aBNKW9xDCzSvJOiadU2owc6GUMo8lO0xuvcVZ4fOID5bEJZkeLbvo
PyG9+GNsddwxmdo8pIesiRPlw1yaBx+q7KAYnvbjX0KfLrWlbV9oVnmZCz4QQNT5
lOsmcbkdbjSdfumnU0wE+/JEORGVcbrdGKbI2P6lfnoG0JpMZdzmnULU+zKKow2F
SARR2xSHvnm+gKFJ8sTHDLRQuiS9Z/5nNbvuqf19zoBLzC+PJ1mBBpJZvoeWy1q+
3gab19pfSATJ6gu0TW2fXzVY1atvXgm+h5/T4ovPrMIH1yWvi69zgCIbSlHmEbb3
mclmCv/UJ2FL7R3R2ljOFKbJ8VjyT5Iq5aeBpzcQTmPB2RbHnkOw9fVBT+YJBpiQ
7IUB72PWSCWIHwBFZpyjdryxqPddPacfxEc/5sRRE1wjlLqm0NQ/1R0SFJ3df451
zsoE2VRNlVwm3uzfLllVR4jWWofm9p2c+JZsdJiHLC8rakP23w5zqduvqy9M4i7A
PcLVzUlpGgxaTPCnujFCzdfMlGTvff8qQH4vpIyRGrhlucryFmxGsN8fNKZTNbXy
oClAyZJuSGzp7HxGVNe57/wGWQljNFjmTmeoNeTc/i+CMofiVsuPwB+WxEtmb8/Z
G4glfiqua1AOM+dwiQcz/5UrJlPLCjlxw3+cZ34G/HbZCDs1OfHlEIfqQqsQiSdh
ePgx08cMphUtf5Zc9oUcXYML11el8MMYZ0IrvOhNaNvLUWYNQ1D7jd2pggI3qXmA
KU7AR6tWZ9Xsjkf9BSoIrUZfDJRrG6btWCzAWN50y1zITXV1DN0nmTNfVS5iluPy
WW9aEDo4Yk8ARzUa9R8ZOtf9R0PQlywCUuhh2P9Ly+/W3HqryA0hunIMALbcEAY1
ZxcqB4N5owp9z/fqN067/9C2Ggc2JFCmSRaPbSj6egF7fVkLjQmAkhnC1SynqFat
s0S2Kco4KY+R8ARYFnRnMyyV8r4TOwMlpt6V1e7qosNTJo2YRwCe+vFDRI2TaZgK
EP+Uao5ow7nafE+w737pWXE7Avpvaxpj6do/EQdX4eFG6Pw8WftMrCQ9kkT9EEji
F5mLNRZOg1YlYkEEHlpKuR3jntvSe6uO5cSu85g8mu2s7ey0I8p+XNmBjEpr4mSY
eLDbPcmO+Wjbtdluf0pNT15yvwIqJL1pAAMZfTf029u2HhZY0XjNSwvjYPT10eA+
7FVrm6/TQC1GZMPwIx4eYPUihNUpyaRvSSgZmsQuYut8XqWL7uQttJEAOJX2+naT
lUrf1m8aP64lebpBj5GckUqzkoIiEJqObvx1uFW64gR3Ym2DWj12sth4wZw7SgXj
HJhJOgr9x89cpbj3qj+7buncTcdFi8a1e3e2j+JyyUoFZmDRUOuliCn3Na5qQpMI
qIX7w9g+SAiPsBF/3V4lpWFVhoOQS22B6SpqCZHn2y3a4iDspCj9SGvb1DPG9do9
BajNS4fKoKNkU1NNEe0Gayus8G20Gz0m5cJMk0H1aT15PnoIQJJ2wps8wtB4VRwD
zOVlhfdlWn/gOp7TOeU8IxURQ2CxUaAEN8CMee/2wv5SGzDFcajv7d8q3K9se/xL
plj84Hf089N/V49bT12Jqw/2IIl/dKsh/qfcJqTl3KAfd+qauOzZEfEi/W2yCsiL
xvbyeZgYNNQhPODSrmMWiAbZgixAH3TUF83x8/BKgF37WS9orl41j5K5AvsXPMSF
hGgIGY1NmUWU54i+9UPZf5fgOnGhzZajNZLK/XKG05fWqCjje8FkrYqrysEK345N
H/zeq9ugkEuISJRq9MbMu1SL9ma5cUDtYzvxHXltyUjW8iqU+Pq3nGt91ETdVxZH
6xg7gXBv6i2lsAX67P3JqeP2A7RCmzQStueE0DseMJdj5tsAUCxBhn9YWBd2tANp
F6/1BaW+1CvsnwTG7WTG+rXlwK4ZU0dNqck7TiL69ZHdPfhj/7Vmb+b2T5UhbSJp
fR5Wv1puQeo8+bFXgs3BIEdYQSZt/EWeMaca1b3CPEwfPaENpvbVX6EXBwTFghi5
GQozdaiVU8RbAWCtfAgHFQB6gGK6XNRXk2pPkru5wsJnJjLYE7+ytKeqJI7ENhoj
LckIUb7PtxoxErD4hWUVVdCSJlZNPhC+JQ2vHVgj5qlL3Rw4Dk0z4xJdfHDc1IFi
yGlPgblF1cp+g8M+GDmZwLbFTUV3yXXp5ZstI79GX78x0Kr1isB+X9piTz7hX8Hs
2BumIXQeX/TqBvXEy7wZkHiB3ELYGjyq601sUvzV7GisFcuxGbi53J4QzCfy2FIC
8fEZB++CqvT4s/X89pLFLfpLCgKFmXE0vXKu+/5Y1scC4MEnKGMvUn/mA0puTeEh
CEJKa5f1fdb2frKT7ztfhO/Z3hU4Kpe5IBYa9vw1BiWf5o/fzsYTuD42wP6vceps
En5ZzFmhB42cqdSrr8sMDwoFdeR7k8Gq0Fn3sHdKN9D2WBs5gjRzxDlzu+2K7R2K
Z2ziOEJvuaYy8sCXcToAPZkEeClndicFMIaTndQ1g0eRiYvNVmZ2Y2uQkZVW1j30
XnBrbcUX5jiSMTqlUzE7eH+lMuQ/dt0uNovceJ1hivwsx41jlq7x65R2WnWMnvnG
lbSXbWefEQ5jDE8o1tb8evTbVZ5ZAg8iIsKRdlNROyeNqk8PJPGRk8VyROgSk6QN
LoIlnFQGCvAT/CDhwR7yY9n5FbOs6d50LMYEkB0wvbKu5i35Sw/HbRqtpkp8iu6i
qQFXqBaAkkZZ0L/K+Saz3ngDamyLpqvQgInp/Ltjh9mp9n6uGLhgGGZ/jKUxF1bS
5q0ZuBw4jaKIz5d1iK6UBDbBuZEoaiEqtQFnvsrmKMal2iTkuG7REHcQpBjnOlYm
ONISqjHJCuxBgyuuTRqHIxA1gLMWrqsAjSdrAuRxTIG8YIdfM+m8d4gE+FGzFAXv
W5wJ3Wck+9ZW4DGo9ZtrxQeLwv8ECDAjqn0l31IsyLfJtAsQuEt5kmCRxHtTQQww
YvBY9IkEVBPj8DLHQD+K5QvJuST58T6o54Ve1hhUhahMueFUm0Np0cZ5Nu3PbaCj
ChMX4XlBV4kYqwTTDkrXyqZC6JfX6YpOGywJcGetiiJTHGXPO5YCNJOiJNw1sjhq
ZEKfk4CtdJlIuz/+1XfTmyRmQbGqIapo4bQb6yURMIqq0tX/SNaDk3wFSzGWZRuJ
Fft4jwjew00x0FgLZrJK4XDJYW1wAIkFDrmXwgHJNreTBtX1K49YLBR1i80sab4b
9yy03E9mSJC7dZI1SMixgWUeTrlHwC2BE3qch0AhHK9aDtRJ8ENoEtzZku+9iO/k
557xGpUYBa4SoBMl78/oH3Z8dk/+9CcbN9WnvbUVbvGu51lVZtdyx8v5P/GfWFaQ
hKIvWVqYwb6302J+lzc0Avf6OqLXoMJiH3qcrq5bmAEEjrsaWWMmYCpVoJUZ6PiL
dB0xOkH+53UqOdxE7TARqQqPDkajWqo0VCsDg7HDVBcLpWFVrV5KJ+n+cpf47aOn
pXDOE4AvgKwOXJJOq1fFFCrZiMZ1aGaAKUWGFZ/t+SO7u6K+LhbPBOkoaLYbuhR6
XgAbAMtKNKSJG7YbFA/YcLKRZt6lAukOdX+5aDJq+oCN4Q2m7tinQHmCu244gSaF
LUbaVDc3pCYtuojvCYKNUW28oVKhAgxopr3Z2HpBxxit6yJQXfAWVP15oPeksP4C
8GtjZwsCcew75B5BQNoUhisGomrwgO7NzcDyZpVgESNYVFnOusZ+j52tjcD/qkwl
14Ms+ty/k0IOiG61r05PoM421Nz7AVUSI8SY/uXi7HNIZEK4a8WxPb5H39Fwon1Z
Q8JpjHK2Zv98fQIZa06czVZ+wK2xgpoubAVGA/QpZ1/TFhrlcd1H+uAPlumAud55
CP0mOfBVuvDDHXggUyVSMWd5r9OuJx3ZdVOYCllYygQLBxhqi8sJYv4ee+z3aqre
i2fUdW/zTXQFZE1BB9lkqAIxClQXJ5aXpz9MOQ49x+Ymrg3n0BFnSlBz6i46LESn
fmmpFtWPtrPwqpqMyWG6WXHHoPPcWJzWIR1VgRrtgSQKr7nZPqrdiV+vWe5CpdAW
ybGXdS7rHwytplhSVNnBo6HfoKc1Cwqos6DtBJOIfdw4coEnrJ/JU2fRLmZCX9mo
TWPsWd2KBDODdyedj7jL+j5DuAwo1PCD9kO6hkD/oE+WzBrr5njmm+dZ7Ma9YfG9
6Lbjud6ofbXj2NI+RxSd/y24SH19n+51XjwQYTA/dvIRF1/AAyM/nlTFg5wKe8LK
iOypdiZi95ZUy93qD84DVhFZNFqmmJe3rcad+wIGU3qLVZF0J2+732yBkf4x/Xn7
A7dKtiR6aqFGh9GIKEq3rdIkLXe69kq/W/s3M2i1qJWpRPaPx9ucvWwdfRx1UfCD
3FxZJqgR69M83Rk13BgZSui2uh54heRflBkq9HP6cJSgc38TymYoSEODlaacxzTF
B1jYCvFNsH3DraRGDORc9L7DkuutwHv6XMmscYLJ1LJQJtnwPX5gSpcLbFaspc7J
FynyDdQM5cJoex1Vj+rRZG+yZFfXlLSVLua+0tZ8E3TpfbnqlWjMyrWdX1JFvK5y
Ba7p4qIxn7VByLg729hod6oO9nUdsWpYtelOvMr0My0OomW8AqyzoGOBYykHxgWB
3zvnqzK/deU7lDfuPvU4XyKrCRJ6CR48TFn/aEfP0L4TpKguDwYmK3eB14Kv1Y/w
3UBJCAlNrmRz5kqJFLogl/0Hsrz5qHYEvFQ4rOuSzJz2jTjZq3NkDmJaBjURNA5e
vqE3Yb4XtwCTKfN+jfTfJJC1soGDi0JugOiN0KOQLmXrZxKUTqnJtpDLgWYPj9cG
DydIenQVvpe1uk4oOhJ6fNh1Q8fNfrQAekQZvsCvZjqzXvD2/apv64KNRIVlOHDl
2X9dA+uSXB7vqV07CApLl4eyRW5SXHdVXRv2CzFlNDcowe8Z/iueUR/ykR3yHh5I
mXm93s8W372L1DmJmom8iyVDlrm+TsX7xHHW6w2+3XUFa0e0jmhNk0o8tF/bHdh9
G9vyipWg/GCgZsMc7Y5Q7DOK5ovW0mGdqzOoDo0XSLPdbrklcAskoXwyLHlB/sYJ
LQyGF1p/HUEAqpNQnahHnOeYgt5ill3K13191P9+/aV9p9WW4X4K547h+mleyQN1
1PdlnWhjc9Ez3ROMdoJuQGroitMFMqQhuqlhl+6pAQ4VVlZD2/cEhNGyLdYmTAC/
XfLOQUiCIjPtz9iX8D31P44k1uQiffQNQ1CV7vuR+iLe7JLjXnkpKLe8JSml5qWg
/j1xjegTzMSnwgcocPQTqyRYA7C4X37z9qVC3PQUtDzuLk1UrRPxvc0b5l6ORUE1
ZpeNd+NURzLXW0fgRnvVe8rdn1A2qdbWVxZHYh8dz6o+Byil6QXYMRqkewEKetWd
z3tkQHhNfEmDh8yYGqSvYFVjh45GizOwJGSd0V28w+6IS3uXnDSBMsb5J9Uc5GWd
wkXVuYAQcJFBc9l48HAoOSYBa7HF618VUMgS4Bn4jPeCwYPQ9aDFkfM+pRWHQTl3
nC4op+TCRm+ya53+9eaLDtRSGHguOmsHdowcK22eCEmz5W/7PmyvjrM9AJgn/Ldu
BYGhBNhvsHPM16BnVLYUkdMvG64tffjB/Yfqhva7+IBuIu+Y6CMEJuW68bk0zVPQ
MksL6N005c0qdOgpbSCM8/kSxzy54ESxWiIE8PWvH1DWk/IzoPOT6/pyVuhiV6LL
tAAcVN5icvRgZ1u0ahrI14D9moeNyjTi8A4XRqip/d756P5EzkvMbZEJP0pUprON
FbmwYxtOSKHYYWCKZzEx8kQ0YfO9HcWn1DKBIjetMGkW2BWmIDeb3Fr1MUQYRfHA
sdc8zfosxM8MybXmXlHGncNN0ErPzw8kzQq/RJ2dSxQXZG74EsoUBdOBKWReLsZp
IEqkcTJaGBULNHTJhe9VlemYaY0GuSMLzf3rn9z6EEXtbYCOw0cVD4bjB8hfOI5m
oaQGVK3kcmKuoc6jImO9JxAyyyCcLApuWbRoyykcwUSL04hAoeGwpBEyTdEAQXMR
5ASgKeyR+a5WfsGLXrolOICmdJLWiVgeCOPssbUXEqrS+hQEt/ziOaVnMvi4+eir
CAsxjBqprs/8q890mVUFNKdHoXhkIi7kecNY+SpHfx1g8cuwmW9jZjGv+8KmH5b1
yg0eL2x5Nm4ND8SgkbLwGMmRxkAfsDUVwO13rSUvjrZqe2Z6MVle6W5GWFLrOij7
rM5m7LGkrZDJh82AQ4q1awCyY1ApxxIe99IEqDR4LoVe/NBPqMIJJLQQA64FybDC
vAtZ0Hob73uj9TLIfg73SmE/5LxNKQg8AMVXdvPvke66/YUrVNL2lFOfyqHqWomq
+e7N8qcb3OMp+lUC8WS/mn9XmUlQQCzFrzNh9cUadwNwpjPN1pF0WIRgAIj6J3kY
G20LzBRQiHljVtw9C9r0o0Uz+qVRa6aUtr3rYkbU5dOvoX5W9sQWzP0d6XSTwu/g
ARn9SBhMwImpZkB2Q2A2LJyQQDW7QNpZTe6Nun+oZEyoWchQWNTDzye98wgrDM7Z
ihv1UBLP6l02beKNre9iZaamjR908ez3EVvctRL/GHrhuHSTDpR+SARZmVT2WnkO
dXYojDrYaKIauOZQLLboyhovcrPJ/cKI2JMS5EGiuq8ts0IzV7gTfR4Zm5N9uM0U
E+GqsOPvFtpnxpKqSpUieI6+fn8jz1lxk67VZgrMWBmyrfLTHRUN7TKyfnW4wlyA
m59FueQYhx+UKuDW2/G/dtiJHU8aPoL26/nzRIzTzKjREaezq4/p4Ws+3o7Ruyy4
FaJDJdmrJ+flgNmAtieNDjelAZOqRW6QxWqMNDIF5fqD3Kpx/3i/ewM7Av9lMKQl
kseHWI9XL1gCaAcAs7jrG2P1YOnp16z+Pju3YADGarOwxb4I+6NdqX+h7r0eg1IP
K+t8Dy1+I3X40xd8nCAJ1bAGTwO5SPnDx9jhTBU6x0sRdXWmzjo7izLIAIkUHGGd
rCdbl6jZ/X9TZd16QOrCTMFJvWe840i0FPjj5AxJrLVnMidI9lgMFJTp6fthB9no
PSP6M4neGHd9V1pYVfJIpkZC4sKeBCx8wR4RiJqQgEySLcFPC9aakac75NpUW3vP
RX7wiFP/Og10vmGIgZNPjxuxpmZvqPp3PBWBQa9ISrhmEZwN2XkCi0eiGRlwwFZ0
peKDiMHIU80OCUZp7MKToDFrq08zVkBFG+/Kf9ey0Hb9nDnnuFzdZ6QOn8mHYKNK
tAYzd98FrHQSdQIRfE+eIIbZ8xXmby16ctQtjJwq1cD/X17lfq/bG9kkFzWy5pwX
cax3s4/yWCt88EwjunVXKUkUaaIWcqO+ZlU1P4ZDrLbPvc3f0ZSyyd7CFm1NmB9C
bmmqpWvR4p0ppTMjVduk7stgX6lxsWP9SdnblDUrVji72hC2of5pMQsG5INlLngn
z7IAb7aJEGt+f4kgjKQaZX1MUnSHhICLnHxy4/VneZxW5AEsNN+4RlN1f+Gqa8CA
7k44s2qahTKIJgYi01oJA6onCuFvTCYDH9tGFSHITeCDvUgqQFtfndjVQqwn7rVw
4q7+CK83kSXsDGKbA2uFanxU1Eckq8v841zDQwG8ZC02hCVD29nDJcyzs6rdqnqX
frW/hz7yA++tTgvn4a6f6S2iDKDR3Tz/gXaJjohSjEoygMM4hyumcfswv0CUiKJy
2aQ+nooUFDGdejkad3D2ONCp3SbTwMQtMSYKWryiIcA73zBQKmHNMKpI1ECgMNaK
NweUps1wk01MzC/rR0b4GFtSNQ70nmh9HebY5qknXq0Wqjaa/KhmCFlMc5lZqxwR
1Ef4e33UzNkzqud4J9U9TbQLddJ5/porYt9HKUf0FvvH5kwn+EUZkbuUB4awAThH
QSckAiDUaLXhwxYYVO74KMyTlsqqicWgy8kIKb1sSupROHFn5O6JWW3t8vO40JjE
r8fX7+RzKrro83ntd+XJKzzpF4xctoDS4QDZSE0bHE/FyqNnaRz4+5pa+6hGmVrG
6dxonAp9Emg2L/vMy74A+m4Mpv5yV6kSgq6Pfgik/gNSTGMRHY+xHZJWMbGLATXy
/fjE6QiX/0HtI0zHQPL5S9WXjKgaxSKJl22nttWwyfpn9JLGM5p2hLuS4eWHqTs5
Ei75bp65az7/ZNsCirMrB5nq5WRSgZRzLtrKJJ1MbfhGyxKj4D/PIyyfsgVwwAmF
t4E3hpdh16CN5qaTPnOZnDSLiU4SCjAOblHSGnZ2IE2A5/N4zBk1A0OZNUxBoiqb
j1YHaD7L3FVEPoS418HvqDw+9xHvswOWw6KR5YffMC7WI/EnG7G0LkFm3X/3A1Z+
7lBhH5pzpBSyGTDP77vBbkOqtMM+8qKaitro3PJg5zgIS1XWFD7FUP+gbfLDr9T8
Pks0+JsquloR59XPF0qL7MAWCt+LLxm+y80Hn7NwuSd+dYVHz1HL7VgTvga5BtcV
lxOanAp/PuBMWUX9Z6U3kfLjPMWU3GQIeg5+L/8n/HDu34TH+S4nEhgOJFqeKL0t
Jo+FZgtXmUUkLVeWPQi57tiyFTreI2f4qr8A4QSzT6bTrXp8BQcXx2EsZicCHjQJ
AAef0+Xsk+q1arrcgX9zvavbB4v+012jgarb7KPKerFmnxLk899qH6Cz6afdea2g
/44VC1o3t1pbBWz1/Efwf6ZXBhRqrMQk6brdj75Cn40Ow4AKoqfVHrTz9XYnVMCP
Q+Rtn5MLogL5trhKv0ct/OHNdsvLVUQi8Iab00PDZ0dJFI/k8i3FuYpezQ5oGyMG
IGcRqrNCSW7VpoG3fH7uJK7pc/ymjmhNcNyx0rGlGmSJsyjpHoD5YLXZMrcjD8HP
Yc3RakKxEV9CPRj6lEsYqxtp3nI3xcSeVeLOKdKt01IWcXQnjxA1ZqiOOWF0g3lC
r84VZjMkStnhSvu7qMRFIOzhd44GbeKqHX2X6w4Ts6YdS2Q+yjKkrWuRBIdc1oei
OXnHOhZIbbhz+f0XBhkNMeAm7o7Nx+aRE7Qbb867iPPDQ9QNdANsoaiLhNNwUW5H
5anqJznPNGPO7tWhXUa49O/WQdM63WVylj8uLy1uGt49f8ZlUdvPSt5FdBVegnm/
GORX5ycauwl5kFpZz2S9Q9t4Zfr+RM2NL6Xol7sBAX6VTmfu1VqPVUctUpGnrhzA
LsofB5uRimvEmZYnYJaUms9rYfUihzsBTjkIkamwFOVG/OQ/KzkVkuSGmuA0MORi
IgNrEBJdzWQq0ZIXzA8jqh5wHgHsfnFJ3BA1vGnAup2zjraAWseZWDYTEEnN+8Km
5uVK/LfVfwQ0V72mRcRwOajwIdKYNqlyYQexeWQRRmcDeIJXXn/deTkI9Pty3rMw
YDo977P4jqiGRsihfcHdgdvg3zPXrS/AOsTXb1r390oToKmWkcwpYMLfUUaSDb+1
zto4sWNkhTFKI/O6eEuhzwIJIQcnpjkRne72dMndhs91XFvUrad7808PZVSssOpA
LW68v6Csw8ln0YUqyqqJfxHbKWjAYRvEbYlPUFStzCQe0h9bscqVukxrpmG26Y3V
Oi/1xXVB+4wblXPt8X404PN8vWd97gDNuBOH0gVFv/tssihNZwbBhPa74BgviOG0
rlqcXPsaojADn0lxdjxjUBC451ILBzhGTq2Zf7mqjUDHXejibx9kDn6YdTBjjgxc
MXwaXag7evpUF4g6zDh3G1F2Va9R5YUPxhgJhsflEsMYM7qgityIuNhbvvxc6Akz
epoD5xjm5594hNodJ1Vp2jGtieTvWM1j7RzONwGuDLjwAYzogtq0eKltHi5q+m3U
tu6+kuFx8bgKCON40yzYkCkT88ZCYrEPk4WnXM7FUciZIKuhPiqtU72H/oEsuDVk
Pfq6ybJCokuOnFjDs9UqnEOsbM8t96uxM12eYxn/KgNw5P94SI5kjK8ypuHsyoWk
FlY1pWvS3Ozwtx+iBpILXXoBGIXjVBtaiQrKzbIPIvUQMS5tk1P+2Z6BfxktqcU3
rVJv2UyBPuqTTuumNPbM7qnGxOTbkLnQSVmp+QQkb+H0eYEEO24XKd6jXU5LO+A2
+lDHYwLcsuFZxOnpASHZMV0jVKw/fPu0p3XWty6Ro7ZdZWO0RDN74f4DD3vmFJLH
++H166fs+jnqipgdZvRQnyDzNmbUCgEg9Kn/TwD6oI/VUVbvk7tnYXh8/mX52zi1
8yYMPOSsA7XEMGYocW+Bg7JXYAbu7zh+aww75Kff6KwsLpnX/lBQMVBG3Y4vT6Nc
hTVVIftBlCLxBu1gmwPwA5aJPMwygNUafIe+6kXFH+tmtY/y5qEupXVUmB8vU5uN
72I79MGyoGcRatdTT16jlV8oTp32WO8vNziN5NsRSrrbdzlQg8JKdn3mK/BxJcvt
uIW6nqvZFvtB4MJEF9X9JPWBY1HoxROS+/KARZ4Yb5lfBArMNy0sZCeywcqqbAs0
5pYoUkI3XsfYGveh2ed0AqtF3jOFUbp2fa7adgFxjFVYbBG2mcBmZL1BLxSoU9X3
xtEfhZn8/naGT8t55vI6H/JYLuTW7SmI/Mu/ZX/ADtObWX5j6Vcul5SHCGCJIH+q
u46Yc70wm1O2fxYsyOKIwCkeQ/osiDDdUfL1GAkjeYAd0IoyHwtU3g6KYv+wT3nK
KjmBTYJGw6MiL2P6ho/aUEK7lOVt6jmWRDdkZ1EKNFZDor2k50L3cpsWOpj8pEZr
GGq6oSFSYqxvRRs1Eu4o+mzWDEq8fRbFpo8XX/vM1qD49IMY5I2cUyzq/TnOhNAl
dbj5Xi/tq/YnNmRIfAn4zVIDdSSk50ebZ/TpElRnzl1SMPH73svv3co0W7VX3ETJ
AZaOMuuPzlQ+61gFbTckN4cFLAabkaGfSMZ8oDOsSVjCfngVhAVYUPS2Sne/WeX9
lpp2gMWDoV4Y0yvk2+0WkaZBizdt/xQnG8d7FMRN9djTG66oNyHBVVA59LYUnHzJ
FQnPm0lQ4Xrpx7PuUPxGcBbDPoZPKERZULicZ5iLAr62irt3TTxQ9pwfyM/1oKoM
b4Mgd2+Wh0gB7Gu0LnDxMklfb43iRlN54BP63uwrg9xmHSWgs0rtwMZQH2C18biP
FYg3XLgWLmC5pFHEtJ5CeFp4L/W+l6naYLcL9zHl5r6e++TX61nhxo82uDNMnNlc
tTUztqdgBZ6zIxEbgYn0BLhMMZHxoABOIbC6tPs9wK0owlTzbq2UtA0wytFb2Sfa
kiInJh+ciB3X90xWiOxuR5NzusXcuri/dYVxryS0/gOL/1bE0qeG/tTicBC05qBH
Peaz95C2rp61BIrNfbXmUzkg1xDzG0AflV6hVjCMRD3SDmon8Bty4TTVTsXqJa7m
PN7U0dWT4gpvNKh7JzgqhvdVuE9xMVU4gz8AhReCTFo3P+NnqZ+OWe3e5MMgJFEQ
foshcS2ZEYEGg6GAbF9QXFSNoDb/2FkW9NsPjwKxYjcu88C5soF0PCoqhXxoVqmt
DfMlSSW3/NBwGP+Ch9W52n/OpugoiMr0PwlVq0UVQ8boqtY9kxAuce1yxp3qJyYp
IlyFh7hTFsDbHZX1yudkt8V8o6LLPaoFqYwzoI8X0Cqu2mv2C0abm1FETHaL/RxD
IgYVa4Kj27B7vRo4F4q7j1MwWoW5vlDE9Frjbtl7DxRdxqgXSkrVlUhdKilb2MwQ
RPk++mswT45l6K3+LVR6uNMPdxWXUlAPojJ883V2Ni0qwhvJHqlqMDqD7tjhJ7OF
tQhAuD7SSRSpAk2z8a7RS8/4HKRJ9oQjpSoj5V7dagycojy66/7TiUMmdSz1/uLS
m/FEJ8q9QPrU2DOZOGmnm/EZoXzcjksdCkUypYIasLWgUtBa6Cq6u6PR2FCEWsEX
UxQwichJBNqBLM/3qO2p28/J6Bb1PoGMCwaAUJP6u9cgKil68WFpdpL808zupePW
rQ3ICbSGeV5L0LWzEcyR0p2R75RWrdK9Bhhyt3e0Hp8j+4JB1sgFApWVV8JW85GB
0XWtafnhydB/CcR1FlvEwz5tqRDMIXIgldddQRLYOP2+hA6TJxaKscVX4HYFSTXZ
FRnESTh7YHtlArYeIFHuqxINkcaIcWhDBQ3z9SLyBYDR3C/OdwY/OrVXpxAy5ImK
0t/QrGxz0jmQvBvlkBQWfUDcBNqaqQtJcErxQZYHfqXYMCgiDxJcHxKK0Z6tI+9I
TXfWzIn7oVLah3oA8A4Ckf91yI1E5EeWbrW3O71znJfIgtOnzkYyH4QZaDReLX2n
N03s/iOJTOL+Qw8NGnRkYpcmdCO6Vr/axNqfn4K+yeO9gmYO/f0Z0PDyoM6NxUNq
I0PXvZvF30g4rb43uxRiEPn303TAvs4/7ttc5n1VhZbQEGUy1TjfmxbhTdBKDiIc
Pjy6wvhCJTsVT5qIYwHhiDnNytPCzpZL4Jx0Ov2KKQb7vqReqQ08PxzosxhUqNko
GVBCGg2uxJYNeyXDbpkcAbFcfV+uQOFOFpl0ZX9ae2Yc1mhqAWaNU/qC6rky7Kif
pHlJl7K07/xqGpSH1AsgQ/m6JsROjnZljkTsSd64YN8ejzw1LDo7W7eshXOW+y8G
afXCkfioPp+FBwASCA/x7g52HEgNkF3xZolCFDB1rSYoEdbN2BeB0zjetUg0E/gk
2qKhtV/n86It/rFzmUMkyoVKrLfxFkaC9WAaXN7g5bVFr+76gCgr0A090zCF9aLx
Hz46/KabYJxJgRkAkMdcpxSnoaQzPyJZokkNAdYjBe2D0J4znMDN+gi4UW1BZ6yr
fuKKZyla5Ubest4JJuUXqtn+jSJZRvZiyJWhLbnbQZay8A/IY/GJ4MICXCaLSSM8
iWyBMTEJQrV5jVrWd34oZJ0YXoRXg6ZTIDG4Ko6NCo3QV1/r9xczLoFQZoszozZO
p5tlu/G4dYw4RitL73dOB9HU52LyD8wzrFEzMANWfakdu3lfYhVZnL5xIDRNSK4K
ORXBm41rt9Y3B7LvqifDIvsZ+lqdOHxQ+pc/5U0PutijAhDDv69a3Ejhu1WaDhz7
91E4CNCHq1wITJ1MLDECYdj2oLKCTL9bzNbaSL3oMz9xxVHfG/ZqBhZYRUCzBCtj
Zk/2Idjtu6BPc3UsaPWeLdOyuQnp6PjyKBbN2QmkFYjDD7IGBmIPy4pVruyqenHi
bHmqAQ1OjvU8I9iGUe8+HdPQzASqU0TijTxMJzJ2sZHqd+aRQZzf0YYpwiZx3Nq3
ZzRfSYtQsUH0E7hFHRhuadeuni4UGIBba4CHUa5/nqcDr8TzxPV8Ue5dfHMdNfeg
s3G/mKD2PwexoN1OVq+sMjXYIUDqNbv7/ac2ZHTNb3zUsIrSJ9GFyhPU9EC7ASTV
npmO0FlwsJpBseJrNGEbsfimRAmuzuPejmsi7vljQn9y+m3A84gdZIKa2J2Ie8XA
YXulVvX4njklluh3+vzmJY++R7xB8ghzMc1XM3JMsdAo+Z28mLMVlBrpdXew26QA
QptRZ6gxHyIXdzPfr+cKI5wDU+nlVv8rtMu76W0+d53cU0e0PP5cwvAyl4QXf/yF
rO4ITHmlUSLcXVBXo4qjeo1LGOLpmG2aM7YH9OkOYL8EhR16Rn94T7gW5BBQauuy
Tkpsi2cn2LBbB5RuzbZXc0r0llxqYC08TSqMRY4am3y2rDlVKCQezebvUmX+lFwC
eSJuWOaBzgQ79cxknx4P+kqsQghgRzW5B/OS5GuE100JDu7fQuLYxSjyN5FjKiAZ
O2fcgEzD1RwQHpOnwGN/VzE7cXj1FN0fQ5fFUwQzrhdwxYZlFZNkCMU4bXxoHeky
Uoxslog93fAjxUFqP68gnxgrBGiSNEvNHH+0KMvMjFDw5dHRSxGZz4NBPmCGTzMU
h0Sc5tMrncA54BEqDBN2Gy6GUY4jPdfWQQtNDY5lJX1MU1G72cVf5YuN7d+rFKRY
YA6f9yQgCo//wSgTNK8udNOUOct1nTL2/vf8MJon3u2fOfqEQ4QuWsWMzcRWZfsp
J1C7spZmgISXEW6Eaxr1LrkV/pPebtL+GTTtVnXbSJQWkkmNz4zY7sv4HxAb0dLY
yeJudBZcRYGDA0EdZmKqsUgccV0AoFaijtqM79q6TwtdxS+AmVbE3OSqVX+Ku8zl
nUMxkoJRzW/tpd3htFOxsW6HHhfaKVaMwiOQmoikFLxggAjqfxtnVSmHaxkDewab
V9BQ5mNs9iQtP0j4WDFt9hMTBaEKj2QkdwOHzVRM6tSjKjsSSXlKduEXJC0tl68w
Tw0OVqwHhrRtEfmHsxE8yShIa1gWGYJVcm8NnGvvRxbKhUeU4dbotBRJiuxjqgq9
0G6HYO7T/YehbdTrUP2M0guuM9Ugsa3k9O4Mxz6SdhEKCKKl6iXgQa9p7b6C2NH+
c2YMpS6PAisVJMyEB/zKhf77tL3a7L/Y4+SvlFxY7ZJD4GaIdPJzNN9Lx2jIzNPJ
/Wtlrx7osJrwHn+hCiJGcZkIvXJrHZx1E7VBVlonDJrmaddx6gIV1Ziu3pio1yKI
qE8tC/4eYDq6j6Mf6oA3dY8pWY+l69kRy2iBtI++yQcsfHzlqa3jJO/4Ep+rGpbT
uIKCrVQ7LUn3akHan65bMimp2TF3d2M0g4Smzt0APJYOJqYr4GNCNEcjQd8S2L0O
SvSPP5+r0f/+B2lkfFfZ/cxGta0E3U3j/fVA+E2tfZYrkwIGD2VGQVyGCAHJ6PDi
6MwIcuxD3LceqqUS88duP38v1m5G1LQmDZZdXwZ1RNTD18ats6+XCVrSzAQR5D8F
nF5ofPK+6WmINCPJ6yO/ZIIhd7YVjpnoF/IQEluaUUEqNrwkkXv98bEMHMhQWylE
Fs6K0m+IoVIeggNjcxl34iLUl6orBMi/ZXTz/IFmetWkTsbMY33BDfQYM1vkKSYd
wIpNhu7/bUtlc7VGS6aYKlhCOoZ5FlrE6X6WeCDV2Y8J3TO/oAj8o7O1rRTPxirD
KgytvesMU212v9RywpHNNcbX5PwYF9y8q8I8oSi05ROTG6GuQuqulUXWf9xKFXzs
Lo/Ad266OLcX3G2akScVFEsx4w6DMfIhB8NDMStCuf/wiIwRmxSQZFCQl+aekDsM
lzkDl2x6VAPVUumpfX8x24EeJnUDn1dvPlO3NN6IUauicEfyS/axI6qh8DuqOr1d
qGg3eK1sHW4hHwy/J3YjXfNtoBmuf+HHfP9p8ZFvJbSZtw1+81ErtYoiN8dnIYTu
6EsgX8FBZq8L0Pl1e/vAu5kFwK2m8EzQBVIZy4uyH4CleRlqHh08ySw1GvZhQCH/
9yMEo3g6SIZDWw5oLH0GYYMXPzo8xC6rq0JeU/rU/I8ho/uJVjLD4z67tpb95vUF
nCVESPxtlZdti98VDK0iQR8VYjTFgUmBnPaoxV66RhmNBK7z3l65AhukBJJJd7qA
+pbBzRKVZCJIPTyyFpk9X2I6aPUYoXGXCpfjL7MMCsUR49uyOWVJ0g4bYW/YXKYo
46DF+66HhVLuaQQSIfSNSqOj5wTc7HDX/8dTmHhP0uBUmRpqYCJxAUSIX2Gc7kGG
WhIPSqRvNg9gBzfIT2TvKgADHyUvGpz4d5SLX/KEsumBJ3tM+JMmBleDQ6v99MvH
rMDsJFpff/JFvaD0UBPtLBsa0JXgPAS1fM2aKCV8s5MBYApBL6SGIaEv8HC85kXX
Fhnr6jVahTIdTItIwICWJagSf8Kq3wqErBfirwo8Je2R0vc7zq32YpSOeMM9KZE5
Bzp+E6ctp+49QR4dY3iKDBvqDaKAocs74XqRuI+NhOrdeX/3TlpI+0kQD7SkgBCh
A7+QofYVefihhgQ8iDop/rcbvpCvitDwe74Rx3R/Mo2fsarOOZ2ertvZsSwBAxvH
49lduQQRVB77mFjMfwCpMTLufLUZGl0YQOXJ4gIvp3XVHWl0jbwOeh3iU8KBoyrO
49JfUkLwDzWVyumJ8iHRTFCh5PB94XtMGoVZfTkaLMhdpbx7j7EP82GQhcPUHraK
FKNqG1fyXmQmQcih2bOzBjUjEcf39wSFntz+i5b6fH2jQQyCDFUIZdGLsE6G7e9h
m+/APjtuY0EqiVSgoyBO7B8qZ9+W6B1xI8bnTuk+kFJr/oHjs1ASVYk4mkbKEafV
tqkTFD+CoLPEZp9v4xHfOGq7HxDc61PPqkikBSFS9qO7n3C/WTU/Dp/u8XLVMlYN
Yrq+QJu+v84/EtNNEYm3slQWKhOL+fX08a4p2H99wYZjIQ/W5ZOEMSU03fGIweuQ
pb0FaGEyILn8mRMSo3rgI0j+Kwk5uvazF7y4N2p6DwNhAVEHEHx1v5bK/XeSbG66
tLiF2hbrnEVys2v5XWpSZC0gysfWcpqSjOU/lC65H5++/VHnYAWZMDLRH0+aoTFE
AZiM9mqgZveJl8ADdu2xpkq67Ok4bb+LDZJ8p7GkFYLdP0k2NpRClyP0zgfZlOLA
hVFIn0/BtoNU6Ln2NqfhKk8TmSJgEuTW2Z7WJLPzDfGGp2kVX8Novd4T451xkjsX
W1MLpAlkSnDvwenKk38MT5f3HBA6yiPMMFPuxizAkxBeaTYodXA/huC9+72yWrAU
9pm6DX3GJETzb4Ybg8HOjqOqOcIiDu/QLN20quOVOTi5VFvE262oRo9Y2w0n/E20
nMdDyR9ym7l/sVwUUjZgoXJqIFYc2KDouPtQPLOGSzBywOiHQQPkTuNQs+qbqPlQ
Ugbmed8cD4FiSATPFd7wdr5MkEL5xXdlO4NiXjUBVZyk4cm31Emz+RKA/dX/c7lm
G78VMgaxAJKgE5T95mo+p6lE3goS9mI0B0YBbAkl2Ql649ObaFQcFR4lc8fXm3nK
bW3ix2lUrRLVVgs4tIbaao/rBkk/qX8C8KQOTmqHc+rKDm8PwAtoXq6MCTJIa7gV
g28GHStUjCG4ujyNMUNS5xSjobZf+6j/Xx+fCnEsHLzAsxFXuOVkgTmIoshwxeoS
lqJ/xomLYKRUSErWxAArX6kW4sJtUgAfd6p26CqZWyhgqLP7ROHaBn2u3j+MGv35
xlVCrotv6KHQwTWKxpou+5Mwm9jn8FlttVKv+HjOUZSXkcTtoI9/o3ZGct4GYTml
bIAYrra3u75zzXQyAVe3twT51BXfN2nlfQNDsjUpfTLkqIbxhttR6qsfQc7IIGvE
p68G6DHGwMjsP9sWnkA2UzkXK858GXLB9BSHQ4HM4f/BSDy/C6d1cnwPF+LvdIdz
`protect END_PROTECTED
