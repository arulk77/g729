`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN/l2c6b9g196hZ6QdlNPbQMFOk3NQdmdMTEOjnuRnqs
TloH8BX9YB87llM3U7A7whPq4th3zoZl/JvJuFTTJAC3IYmKfAOuYKr78YrBzIMk
g0QUvF97cYolLZ7Jgaq7ufhlnY891lGCUi7mE6Y4G4p/iZwDd3/pOuRt/vaQuCCt
kaIdODJS0cm4bN0LWN6NgFgkCkwI84zxuGTd6E4C7tg+yEUDI1fNRjzOprTBCjyX
+P9UHsth6wGm3CERBZBrAV6OWpA88Jm0t4iPDyntBqaHGzBeAJ1KduzXIKxxnvM1
7jFR9rQe6gRVuLUxi3zzyU492bBuScxyAwpyaZQHwKdewEqZz+g8EXKydiI08SC7
PgIjEkmwYZChTnqQEY0utg==
`protect END_PROTECTED
