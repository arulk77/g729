`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wfHUdU2rrazwLlSzlX0iYbOsdrYQs4XNIGdx+awaOg5
WY8EQuwp+HKOzq1kf0R1YLesa3iIP6nulFiF20vu2MxE6ZlYAO3C6jtilDO55lay
D5cy6irNL1DtB5bSDHsHWy727BB0vyRKb75Aasly2bSn+EJPBCD7Fwxf49vNpWQC
4StH8zDr9QrcxJYgORcxCTg0NZu0J8htFeFZcKf7S/39OT6aV9Am+mlmrzJLOXnH
82i3GAcplCuMR+X6JQRxgUWREsyA8EBTJ9I6ooSI2xE=
`protect END_PROTECTED
