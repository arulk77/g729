`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C5TgiAOwHydS480E06A0r8tZRmdOPXKNXimHSHsMH43y
xgGk+bBC4+0V3pkcQBP4bFMZ9ks2/wGQWJIdQ0UCHtovc/PySqmGfFVytb66tQHx
aATlofNs0WWribwtzruzpT5CYrvEI65skW/ZNRACoSkrEff7FNWCsMVfQMYedTsJ
XMZ0jpL/AaPBYT+MzgO8aLuKW8fP336CbmaWKf8/jTDBjopTbGbP4cUGC3wEIO7J
5psQGS9pkiH+b+CAHMKICuQ2jrBiTct6Q1ymHtlc7Pkyuwmf4rmqImA0FhVLXNKg
SV03hS0Gx1qvEloTEVW+LSWYHKJAM5AvtsUgPOsyXLC30kp39o/xY9u/9fhPgoEg
ogLvp/y2ptAKNOvnqIVXu1w7hmC/anwOKOj97+a3PddXUVbtzDf+vGYSLnSg4vBV
EgZHtnKIfO77r1RobfGjllsfk/EoqEJ0AwcS4ZqRBB11UaCz9eob2MfAcMTSQEvX
I7v3uDifOJLydWvOBO1Uh2jaYIDAvxC16hEU/xgMdmBZsMWB6i+2uqY82ldFGA4D
Tk5G7zYc8QCn/XVDoP4eIWIUISZIUzxkoCeHFPg2l5eKy1oNxQNRzEaGcBmL7jeA
s0SRlhuNIBgdXyMbIOfAdgu5vytljDZR3ueqpJ/R/J/j05zjrYR+ZbEY+mEVK+I2
tSks5FQKfOjBRFNWwVjKnQ==
`protect END_PROTECTED
