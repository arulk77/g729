`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
72DKe5MEZSH9IT4s+0rFcLcyL6swMd2AqHKtDvupzBXzYoAK4YnbgvFPUgS76OwF
qsyQFQ9DZFwhn7VKT3EpxkMxjDjpC61X7RfoTFwD+yM2X2xF7Gk1tf2KaNfRtJ3F
XuiV3aZ0IC7vhwWGQC1k9LuHA1fGfER4J4cZFPZi7JQgVmP59XC918r/JrdfV0z/
tIsz8D2KNXaEVjzjKo+fZ2nBUJjjQ1DfwD9HXcefE+u7C/UVkY0O0o0q5vTEtMtr
ijBxz7jgJYZp24v8HsQ/38/irgFWThXIVq/uFNi4q7FUGA71Z4WX58dCEVkxty03
yeSo37lVaFWwBtWfTJAnrBIjBqFcTYrhd6BwYWbJm603Btu8qMVSzHMvUOnXs29J
`protect END_PROTECTED
