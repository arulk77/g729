`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKai9suMb5eUBk3+NHdzSdgG8gMLj426pM2necgV90wx
qHC1iZ5Ue6cspQerj7Xu034f7ddqE0skcZMh8vRIQiuoUPDM+j8r5wbeZXtExf+F
E5RsCOF6PlKxueoWxzhMACfnwl1vyxjwc8Bg5TsYAx6N8TCsm+Ch3eKUldNakvPO
CQ4lddhC3quIrtGWgIVUhZT1BcsklPoRGY6sLgtk7Ajuz4GyiaaTK7llFNX806xP
NCo6TtvAV8K4dktqDXmKG/99nyFgBaXfJvM4/nV9WJCJT9pXtF3nWnfpWY6wx/i0
Ja1Bx8Rb9QIJ+Pberwdup5VFl81DL5jJnEjo9WXkF56djmQavZtwyc3zBR2feszx
A7p1e2RoSOrtYkNundPusfgsIuyZhxOcmYHHW65JwpvrvCeQGKFOwO2nXqv/a2aa
Iy4DzwWTs2ujBKejDY3G7mYMlyfLkJDeIxJOp90T5MAfdkWaM/EthaC7xb3LPNME
X914FuxuAqc+mns5SffGeq2xowTBRCVj8LvwVaI/QdPIvs1XcQR5ODbOwNk1vPqU
PDBFWgqFIwOT4C297fEGdHl6bZU2iV01QaJ/0U7wPsOaz1H3ajxLVtMLzi7FuK9U
9Gr68S24+aWhY596xCZHW3j6wsJ51fmFvYcGcTMWcMevClVOxOwpYulIPGBkRBj+
zFjf0rzn9QFDbGXbE2TYHShYPlpStM9SOPRxT6d93Oydu6X6WJt3VeIwWtPqAIUE
GsLmaoAQcCI6u+Sxak0pr58fpfvLERpk/PCTF9XP9P/gO0GO/DNX+PIjf4o1AhHx
0bQp4EImTP7gA4pVdv5eLhIN2Xm4glwz/Lk0LewDRD1dQUqHmTWs8rTOPOKCNZcA
N+EtzzbEpuR8Q84HgfxGUE9IF0SJc0YeRUh9JIb+ftOCuAUuzkTb9HHcAPKUIwP/
aeg9KEEbEr69vxlaEBervA==
`protect END_PROTECTED
