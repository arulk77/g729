`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBcLeovOff1qD2IM2UsXbnqsQHlGlFUurGwPaTyYX1ET
GGq0L2o0tqbNeIEHgHZZO8zHmxpdFh+BL6m1KpbTr8vwnG7+ylPWNhlwIhqUE5iC
DjtKijAB00RVzKuSlBrWyYLpUkafiOx5scEK3AAy0CCbs0CfDosWBHiQ9lWR9WSr
vKK0m3J12xWN9NYe972mdXk7CIDTaUyTy9vtug1wmIBfZGp1nVp+fk/BJII1oBNE
`protect END_PROTECTED
