`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wnBnMRKkB6k39P9fb5k7IwU7oR9fEZnxsgljSBVQtdP
K+9u1H6Cl/N58FXHYsivoOtSkkOQLfBxEMwgtp5NoN4+S5pSVc1DtoF2C8enyBkH
pB6NyTOUOOsSe+yS4SMOyTdsYDY7j9P3Bf1Psv+hgY4oEWh6uzGlZfmPFvvYk+2Q
2Ku/iQBWjuut9+Us688tXZ6kLr+b8TjW7IACpoISRUJNi0CH5zgNd7oZygyXEJUN
ie4hs+7re4sD2q/NbeG5qY+uCzr/hq2Rhol6nFRf3RbhLAgVnHbb3O85gcd95RcK
tFcMWhQ3ogHmYSTOO6Rovw==
`protect END_PROTECTED
