`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SbGJN62/IplqqqkqUgjEJ7OsWEuzO6qkdE9tG3dA/SFy
XyGioYLjJLdR0OFweiZJSfhMSgdwfK6ZRQ6XAy09F9/J7y9rMzFUM1ghwnOTvCrg
ZCc2y8eMz4psoPSeXJ6tUPeZ/7sW1R5NJvRG7GSb10k/w0cFlRQqp/0GHcet8EUZ
`protect END_PROTECTED
