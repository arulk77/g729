`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFy7oCX3hmhqg0rkzl5su0rNg7kKI2PZjSPmqz7hYesF
0H5ifpzcybHI7eKMhN9HCQhiOLIv+94RZjJ5zbpu/0tgVD/8xDPnPQP/99IGZ9yF
XhAoDhPMVgjGnaA1EEJer0TuYlybbjm87KCxCTqXQ0P+69x1GhBgCsdZa+2i0VYA
JDzR9Ea7MehiYwYoKzVKDFu5kTAeY6kr8FktP990PgqZcZoS7GHTIPG08yq7L4WI
lpxnyQvB/S/iu73Ei9+pjqgQFLRyg0D+djrC+Q4fI4A9gNr48yO7a2+56miDRalQ
eHpI7Tya2qnt5eYv9BCWRDY5/Qzp6JdrJiEkQuEdXdVXdSqvOu1pAhtgDXPET7s7
wPJkUx3VSb9w5xNdjBxcYnAZ+fXKWlglLVq7CJrrs7bk208Hn20yApVAIjk/lSn/
`protect END_PROTECTED
