`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNgO41fobN+tZZnG1opxshkQpy9ADqeXN3KuYXNUY3iz
+TwWjiUkVb1PxJSSMQvpNWmCBybQnVyzT9QtAtBrfdvFXVCX2hFohjUr5itHV75F
m3jkinWs5q6zrJqXJYbhKp0vb9svVJ/RA6d3BWA+XHl7z1p+Ql/KjFO9ySFqkay+
e1q28IW5SY8tIj4I9ksH/12m8nTsdRp8kSlWLRkJKaRzLMvcCwnFsiIqhYqYND5/
OzWPar4usXssufooyIGeqw==
`protect END_PROTECTED
