`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePn7zcCA4v2M//9lBmjWOpihpVRxPak2cV6jKC6PBkQK
ZZco8FDU/v0Xev4TJzIal8s/hANl9mokpXivPbrBl+YTfz3ub/jkY+k2b650dKEV
RGH/aAzuQ2HMt3ps9WuiAkRdrpeVR1sFAbwxf6J0kfyTwyap8hmQxTqk5bOEA4mQ
uOwrVXmOomWn4PDI/nsgZZXKPOsyXvmLaTFLOEQcFAACRwoeyqB3bGNmHQRoW5SU
12edbwvMCbwdPH1J1k09XgXcB6aPodtuIJ39PFConzjsU0BAf6g14MJAkdEhotsv
BJ38P4cU6Em5tueQ7OG2ng==
`protect END_PROTECTED
