`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aSzDBC0xiT6X4JHzED7Q+fNDjEOtyoY3wD7huVpFrFKx
wun2Ck2o0+gS7BBu9eF/y1eCbNPX3UkdxcVZG5F1xhZfkx9JmOP3C4An8oeBjOXl
sFl5E4KTJ+bIKEh1K2hupBXPeOGx+LcAH3aYpYDSbEQwRNOYYqXKC92xL1fA/HmQ
O0u53F8eAmdhzSA+FkuxGQs/wbkDI699yBIduQKJ+mhHYAYfUtrL/PhdDqgzGIsO
uDyjUToUCOB8gDGuyUF9gpij0+D/wdqOk79A68wS5Jho+2uLMykdDkzUylnabfzq
guM8tBtKq68ktluPuNDYbqV+5MRbIzkb5hTVrqsODx8alBPw4+Z3XerOalLRQwe/
AvPAKI0XAydHi9eK+BgqBQ==
`protect END_PROTECTED
