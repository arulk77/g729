`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SRnJaTDBle0/tYT5HDHZ4Mvm4ZHfv1yzEIIpc0igC9Gm
eDBLJImXBqAT9sJOBefxkl1UJyTnQ0VetpYfHCUxgx+HvkrYowG0eR1duCxo4o78
5VGU6Th9qZyozFeHn7nM4Tr6X1RwWvUA9DpOsuZqhg/j3rC6FX4wRT98JA74rm4L
b7c8NDgNtIArWV8QTzsoJXKANZmURLKAORBu+jBCxIH44R4hUvbHt/QTxSxEPOFt
g3nmfnmstxDAQx8tTFKTror/YPrpHf2fpE7kyDo28WDlR+wzx7hXAg9VAs5Ti6nS
68PR9FXzqhybj14KVRWTWo6nKh5YknoDHa7TVwjFJC0cUGdrfgz5Ajrx+luA3ZLp
9SkFlutpnIMvP2uDOIfQQh1deSqsTEWsC0HQBQAAlaA=
`protect END_PROTECTED
