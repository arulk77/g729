`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73Cz73pQZuw5vwOmWqJ4RiZGPpg/tiLybktvNuzuQaWIxO
Y3WMG2uDv5k5uSHLhR2e5Y+UOboqkXQR8QvDIHzZIkjBTuy1+kSb3I2qyCUZIjt/
WOP/aT4TUYtCveOJMhB7xXPqbb95FbnwdBZ9l/UDeZhrj63VmG9yC5GT58RAIuAa
41gkwDG+FIAXuSCNhhC8xc+4tvB+c1XVedqx+jJjjoITjSfaKwGUAudXUgJYgtcY
KAoGng8Qtrg9EwAtCfwL5Vgj4EX7DLBicdQrOfV+8QbYLov6JZts5Otwj/yJdIy9
Vf2j8fhm1pjCElR3srPXXVmztWpS5OPO3mx76QJq2pgnfLBAvSqpwUYQsl+8tJ2w
TY0/PlTuZw9C4eJr5sgOv7CbvVjVGxbjQXqcPXK8os9h9eLicSi3GRRNAackuJVp
IG7ShoUfk+OHzg7fIN8ia6IWT75RjRnsoZge7FmD7FYkJQ8Lvh3Kkgygx2ksMBpm
2eSNUuHMqo/SCdw7Hk/SeQhmqJgabx4anVaDpfN8ZfE=
`protect END_PROTECTED
