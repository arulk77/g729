`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB0zc0N9g32ixo4fAJj1ZStz02rPWFLfvkANABZKe9rh
f0MUjI8B+KTQH0eFhHjONQiJ6Rw6xqgcKu48k/dWXyulZJgGwVN5ehArt6Vhagpu
Y/vUVGFKC3XC3/hsuy/DlxXtIV8w7Gahnagm++PiLnxAyYSGxUZTQFzzZN7Z0yWV
ejW/a/evNFpOWNS0XXQXAUOter2mH5mFkK0ifh7GV1f+pNZ3I5jlRP1+x7sqpChq
1QytdKEbDrpBNU4BIsy6GQ==
`protect END_PROTECTED
