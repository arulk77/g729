`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j5Hl7YkddKwfkRgfRyvr1HcR21490sUKvIkanKO0lN3ws99lMheKBunqN4sKl8gX
25zF2V70Cp9Gb5oysSAkbRpDaGSE7Bf0m7gw9/Ap+XvNicy7PkcbgKNm/+zsbQok
RJaQ0W+W+3Chaj3qxME97WS5A/1chLfiAfrU6vc/ql3O3M9atpSf4nEiRLWQmp85
9kPkhd9B27n+kpRhpul8ejrvbwhcvUUIyS5yNCK2yEFaYGZ4baLFU6GkRdU6PkrY
Mw5EUDCS9ZlV5KHvCTMzdcrVZf0lyAp5EyBgllnO7UwJFoCPDwpolnLghWBGt/7S
saFY0FEC+ptsGXjKyCm4Ljrx6l0AufyvOU2UgegmNYA=
`protect END_PROTECTED
