`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAA1vbwzPtNn4oH+4DtpEBFbnMvb0qRvnRXv+NBA0GBy
DB4vBZGFNk9kcJteI7Jm6/+Gy5Xdp86T80UlhqP4Sb1NlrhCBeGSLu1txAYJuUnC
epO1nrzA5uSKs9cG6JwqQ7a+23Zf2ltr6uUHTJGkE2WTouwYDoVeVE7YRHbE2jbr
imeT8xjKFMUwDN2U3MxN3jTHKddsh54N1FSI4U4kMsSd32+UUzB4+HfkQ4N0etkT
ZfPGZ6oAFbkxukFjNThrN8+IkqyBbiOzIfniZWLhVXkXh55o4vwi2kdbtN4G8kSe
DATaxupJ9/cXFH723hvfoNFoQLQo1rNxnAEp3/luQnNcVtkN3WKY/56WK/qaH3bo
LS4LwP5PAI/UAbzAZ78TYr0ZidrhmyCmzSBAUK5undz5Mzds8v1sSwdbWaLvhJWB
QOrb5tng4uMAUCN/gmCHX7rTRn8UlMGFeuOic7BFkCp5V7DYsxhiFHEdP25sd4Fr
hhjSAvX77y+4t1fUm27N8fzVJTeYBnJ84bFj1kwHxAK+OTEp1SkTRhBMU6rn430r
3lZde0kU2Zp0MQ5Uigdn9nBsSkQCEGEoc5WRxjN2iLmMrs1jVyZZQ0qRh/0cBZ+v
z4NoNfw73HSt7cHS/gUOlZyBBVakmztzdXIfhgpyTPOB6+ZbQf8avsE8M+1LLNx4
TP0lSM40aZaHO684OgZxTrxNUTwLFkC7WebGDys3Jsb6DnyLe6ihROHUuezAvmCs
Oj1RiUE0aboH2KAEx5Feuv6Qft9xmbAioaAHXchg2/j7RLK+dZ5mKoiArR0dUk4L
8KYavJUfzwvkbRSi87Zp+E/sQjuVtlqOpIUcsQeVSzw=
`protect END_PROTECTED
