`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAxghzOy7x32BIQcUTtjVjliFoHKDKPf4yzen+SSBO98
mIlQkTjniJW2xSCMsKLS0OcsTdrHkU7IaBE2LVtI6TVfiKPRCgmeBHR9hUc3O0Tv
OB1H3bTRmmAdWPh3Z6pSNuYGu9DJQVTXP1vkJjcD6wBBNkBfVjHyEcZvXS9LGHMz
A9Vf6QQHmf0wPv6spyjE3DoOy6FN/3/Jkxx9sjeeOygzZM/r2KHzODMT8Fomcegf
DLR1FxWSBgHaMmlhJjsF8RG/rPFSGzrMsOI3OvUidivcTwgcWIdQSQ8deSpBwx3+
klYZxv6GX3+nvVNQXpHX9ojpPDfcfBeXhOSPw/neBTOSBGp+x41iQZvcgDp/y7Xe
nqPAtQYszp692kTENGxbaw==
`protect END_PROTECTED
