`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
92f/CVDLePXooKLrD6yhXZ6MJzRPEOf1mp9tUAG87eaa1+KzQTYYoep4fW/FbsOk
5Qh0Ca5fsmi6Ovz/ysEyfnuDPweJgwIdLxEvq0EG3mLLdCjugS132fh2uibVWjVd
g+DA9fRBFcYdld7K5RzqXLnqqdh1tmNtprL1FwlKs0MyhHSRjGiiwS3CFNJAa8F3
F1XSfoaDj1CJ1Ayl9a8K25PWmpU3smkvbOdv0KNsPSb0ufnzBl3K40lgv7Y3gorG
27Dox5T6aF0sNLDqck+pjbflDnvf0vprN/E0lF9Wdu3p1VSE7A1Th4eXsyUiEHYB
W54u9oXBMQz41pImm7px5mKuK4MNQUjRLGu+4aS1HIY=
`protect END_PROTECTED
