`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48H1t2BqX3yZb4h9m/hVPvv7QgVjliQxhDBUfawoAObA
M9u3Qy/yirNW7O0gJqOrfX5QtyHtinsT5qiXMygLqxjuU4GWU7MdMu6/9dKr2SmZ
cKuCEz12NgpLnbTNvaX76/SrN64G6BIbfFbM4v4x96JTzpgbExxSGSP3Gkj7XDZ0
WpmvU3A9Az0j+TCFnT/QO6PKzd/aJCnptgHVqYlY9619pPXF3+UUNctQuQtNpm+i
US1k2A4NzUGwVsJl6HI+OGTFTBiU05LPpfG8dyJ4aVG59xXYgG9W8eisojWVU1jT
Y332FYiNeOL3z+K4BSSU6Q==
`protect END_PROTECTED
