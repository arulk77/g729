`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKgZ4J82+izwtS74T7N/tGrWC32j2Ya42+vDuP/yIcAx
k53qSVkdioGvqs9o1ijjHUeYXjbwqk13DzY6FEZVezWAxdfKytJPe+qKPYPffiSr
4un6Xt/3taTLa9hvxEtVAd3ikL7wooJAG0o/s5JwDFUlvABElqbJ/sMA0Q2md3gD
2nJbSfhdDLMylv4W21l+2OaIZbg+yJkw8eqVZNuuAsw9iECXnrpk1Up4siqNSUOG
HPqTDO0tTRh/ygw1WUt5eTIl59dYEU/l92HyISLRfx6ZAvoVO77RGC1QFelbauMx
xgRbPdBJMNlAe8oWgtMrPA==
`protect END_PROTECTED
