`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveChPrs8i11un0tcJqrlp2LidXgY4+IwL4etf/vqmzKgc
TPzDf7nt+LJGeiOIqcYI7fGwzj6VwlHvQMV2/kHjqlRjnxPwKLYBmQd2kwzAMjgP
2n8/cCCM5+ztUZdRKvrNmprVY2sArqjYRDrtEYwVfp4TD60cdy6DZRWJ4VFBp9Qi
eNg4/YeFOk4swzrbwdsLZA==
`protect END_PROTECTED
