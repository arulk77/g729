`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yVpBGI/ha5ZoW9q3RtVNxRfZz9L6OS8JurxJgophNCc
yi+iQJbaXLXkw0IgPVl9rDYkI9zLW0rr2ybo8xqw+gu6XiooGC7q58ddNK5yE+4O
do+vrf9Fk/nI7wV+VhJN+vzE4KDI6GRyfHO0bSFQYn34Vsn3JdukXBQMg1vOz/5q
jBHhzPd16ai9wG89yPczYUk6KEoACT/rzvnGajRMpTEaRxXV2FpG1tUUndP4wlWg
M1XpEO/+2rpCnNoxGmePTVGmyrZYDRSS+X0oyAiCBrNmCVS1P5xd5ZTl55Tg07/P
m3mg+YOpplaJsNM1VXyzl2rYT403ZaZJbwipDkcot9h+nS9ZYY90+T8LY/OvaJUX
B0NT1SDiKGClCL0UI0oCFQ==
`protect END_PROTECTED
