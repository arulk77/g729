`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
rGrmqmpdFmPKkaXHWrRU1m8zvSRzvGphtn7gUoMzZ/twRkZg3+MWkQwY4pe9Md9d
s7DxAKDopP/Nfq2cyh7SuxdIhdaJc1+q8EJmmCtgBo4+3fR2TfX5RrIJk5z+87IH
9cmTeBhWZ0gkVlmMA3utvjcJTfmT3x/H3movzAbvVrU=
`protect END_PROTECTED
