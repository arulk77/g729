`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDDjfKOCjfW08pmmpThcXXomqwJcpjApQOF5tC69+Pdy
wBJBeSyRdy6StwTyaaPC6uALHN88nGJtnmJl2ERkz7lXEk0cf4+eKGYzxVcvyQ1e
TnqNUc/ondVu/O8tMzko44trM3YzbQf8vVglt4gPlo8UeQBUMb1T/Ry+PqHUixw8
gOA6aFyvVun8xcMLuAHByDuWNrMUF0xkKhGDVM/snR2Du1fPwin+E6qD6zHEMHJa
sgIBpH2jr0p3RMoz/XAhfjYBPo7/fjl9MKYRJvuPvtjkZFHYZd3/vMZYHpJAqTio
+1qUUk/d/p9qMAT3+fFu/+sdVjxH+YffbqIstCP0I25Iks1GQkaVaibnhYCBzOlW
HnjU5HrMioUumomziNCFZIj4Cw7ESYfBswvxvaX62U3r3g9x9NDQGe988URTL4Gn
upI6HimdlNHYJSiKiAId5CwZy2djHuG9g8pgbWtg3hzrm69DPEjKHEpARbq14C4t
liqcRQpSWC/rAd7AAquSVQ59GtOHZlJDgg7hLsBwAE39QVWtfff2pYIH7YoNrg+b
T2O+NoYSAV9DoflDKfiwXqxczV/CRUqJa6GRRbFB11Os9TGlAyWEHHFtL7Fh5TH4
vmgXTqT6CNFDWsnMFZdzkvRi+O46rhv+/ZQb89kJpqUimHtD5viUkJKK3K8j6M+J
avRZZgox4VW+JoT4B1ZmfiNNCjEWtFVSmaMS/4u/UDiBdzg0+XcRXCW5vMVxI5R4
vlFtMP3kB03uTQI7ARmGf1W3vemu5WeclUaytOpqtb+r7XjzIQzXqlbpLsb7VHDc
4m4U724LgIS4hJ3G0nKSdN34EWNGHUhikb2pf6sqWLU31eFjrghOV42wircvq5yM
Ww/MTqIrZtSkOPvwBnH/X72xIs5d907mq7eyPilqt0bIWfWy3Bziocn9Tqd3zc4i
2hV1l/U3SpKWflHSYNU98b3oFyTteN2MS0ICZjfFvIVqFdc2VOwm/jXfujf/gIyf
vzPNeMn411VHd/tRNoDxB0Nth0cEuI3l0Yr/ciMZhVB61juaxy9kJcQwqVIoqHJW
xgtCkaojFuT4GE128cXzm9U78hZNrQnm782dmZwzJCrCkE32lXV5HpMO1QeeUO8+
eXHh85Pwsg5AF8GquO7dIy+NSBEF1uVVvn80n8gY6MvgZhPf7EeEqnT2tlXbkYwA
0z8W0/wt8PMWj1Cg8lO16QwmNMb50JAlc5wl/f5Wv3JD7tmJMEqRcVxeKIHhT5Kh
Iw1XCdPUdGruY3CC4aoHrZeSMGJexbaS0sJmMtibZOER9/TWs0UtPIDNk/X6TLza
S3vJp4gZeHPaQhL86apG6xLxnv3IVUFIdbB6xmOECg0RD6G4cWlg5qB9bmQm0Vzo
ebJwoCaF/49FkZ30unOPZKStFQV01MlctllU5zvSz6FLIRDJFEv7V6N7fjJ8suHC
p7hUlHH1qnsssIt8wnZdFa6KPp66sZ+2JHVw/vxWZktTxud0N9DI0/0ggYWm8XtW
O9xdHf+oNfntsXwbZrWLhSyuv84VGsUaCTdd0TF9NpDhQPhayqmTmE0w66VMX1vG
iDDH5unVzrWoU6i8GiIaB7+bVG6SznmxcTwHs0CSiMKNJP2Rx82Vnh7QRRHRQeax
fL5IzE/p1zgKCTfOnumP+ZflTzlDRmC2aK1uxPF9zXEYntFI9X/mWWhZJ0094Oeq
8DCs922RwMjfBPfhdqCFhY0KiGD9r1OvgYu6+V7G+RRX0e8AMdMeXewsMJzdTyXV
gee/VThkVmFR7sxNUQY1LIUMlu+Y//1eBMsTCwHb+Lxd/aMx8aMm18s0sRmbk9cx
5/1OFfvEZVhCUd/FlHnN8FMUpmnwg0vGNEJTc0TP/djkkIuYtafVfqy7GpUhJ24F
wwJVH9iGHB09DodhefI6YRVVYb/ZZitat/fHTk13PWSLUOg9vK/xq13X6DMjSl6J
hVdgLB5F3LBJWneGgru6Qx8vOc1J8DCqX+f8Kxqm4QBXV7WSOGaT11FhAqu4RUEZ
Q6e3LefZeJDHm24sItKTtERx3yxpkI0fEF+RAFD8ZkLyuS5h2AIyyQ8iYsV6T9OH
um6s8kKI+s3TFJfY9HHEms4ikcMpmf3Ee6hm5g9q84czyDkdd1huB6mCI/oYyyck
EH9VDlaVLB5MHR0IZxmGUr1pW3uqGovyo835wjVug9tmBPwq5v8biCMrpDJq/4kO
wztLuAr10QiGdzC/1UYrsUcPylHvaFb0xAm6MbREYHJ7+oOm3Biu8ih39gHwWWue
VWJc/DeTFPSDZLs7C3UmHgp97WxhBqopewoz3UOV+SeEbVChmj8r1LMuQrNZVWy0
a9HTymppcaXp8LWNa8I6rOqNbMv4OGfDsGkRbGaJZOYqlKip5Guue44++9BYOrDT
InZPg4tq04uOqEM4tDolbg==
`protect END_PROTECTED
