`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
V8gqUBneAaig4Tw6oDtRlkqWM0L3TC2dO5gz06PbERlFiZZoZindXU+vaHsctjRN
goH1LDCoyZdvV1tOe22SXcBDbUAXEJ06jlZnCn/gBtLuAjpLT/dpyjb8UU0oZ7ub
Fp7weuWui3P5nL32VAxsiJ5tPyHS0X8ic04dLCPMuUOnNFREVD9MFq9OhYML+7DZ
oWhVkwi5nPesuBt3nWgHuo2h6BDIKEkKHTlABIgZ3VMqpN2XK5IANUalMqtLnxek
l/5Ynsh5FMhUhzuV5wI7/R/qbSgSpaPltjP2Fu0vUGW0BK5n50AmeqWpiH6QeKVD
50umi6RaHTHj6KQO/mrjyml1ViZfjzjYetdc4arFT/q6eISyHSLeA4kDaYqMCoat
sr9Q6ytWcFqZsHPVvvugK0hV7L+YbTsrbfmgtkMwHEc=
`protect END_PROTECTED
