`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBcvTflKGoi1oTr6HahURjV5wGtkqnXgPItB65OdzAGR
7v1rnOoto4Kaa0DFCpBL0MkWvwtpXKNnqYPctHvq2iLzn3FEvgZfcgnM7WT6eii5
gw+9IzHnnGQgc1sY2VFWS704yMpoKfhmyw7eOxBBAWgy595q3nukz8mYJux4CqGQ
/ThLmsiq1yKPzNNm2gDOBbmbhft1eV7cpK8uu6ViEfMHGIghKi9erwTHkj+ldWbd
oN+4MfF7IlizUXI06H56V0byZK1tSUNKJxzz4wntlJcvG4mbO2E4kklui7BPQvZb
MYGwRYUpzmdQitMR141h89bCEOjkG2sBDGxb1CXSeFW19iU8UDfzvDUSJbJkVQ7L
y4yBwaiyzURlcoLy5G268ImgY2qOkuhsHuM4WRspS1SKxVMpwzQXWS6U4Q2xaxM2
Ym71jcC3kMhdAKfuLu04EOjtOF2clTzYgsrQr9rVta/b7tx2BPyY7K+3GVHG9hQ9
tipzGUvUb0x5JgmPm6M3eKjGyEXdt1jLtpeRCGO1i4aQluai65Gg9A+j8ytwYo/3
`protect END_PROTECTED
