`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aemdCKb1vJe1OHx+HDITCKyrVMVaki3uMSTKBaEOcpUh
LAoHmzep6eSCBCwFTtYd0Qi0uJbO94ZUOix7lAcBXuZ3RF9Zawy84aMkMiYBvB6l
4t+hvWINAE+XL42my+5YBFiKTnpzdR1vF80rC742zkk42TcC3B57VkYdHSkQbAu9
bLThavDQAyP3q3DE8s+o6JScMjWdnR2advzAMUl54cXnMzxuSp4DBVTHmdb+Koi7
VS9SAvbwtUJwfXdhfc6C+fwWMQaTOGf3FcZz8ag5DwIjRCvb7KlVqyTOV9PpgAnP
0SHu/gmKwf7NVOFQPdAsLWnKMunkg60lpHMPrjOFpxTFBf+AwYnOgSnBIN3W3T9e
7ixcxulbnUnm4E/td10/MM0Qbps8IfxRmpVvWdj/RZTUnojJpEIRrhrkZlOESjz3
mKqmWjkJDlpjBhJ6MLDNxz9s5uwWGBgv4ApMaBj3QenIAU1++0eJDtDTheNlvyaP
8D3xiR2SPtxkX1yQyV/Ilxg20wv6khFbiicL9V4hIPvOEAxWVyyn2pjvxWoO++kw
ZOz7s4JT3GtvEKTwWjUjLDNw3SxMwqefBizKtYBv1wdGRZLUV3CkzQFOaGVPqvOq
ONNUrZ8QKsSkKDDYJjvaPzavJ43Mm78qGsVjAXaPU64=
`protect END_PROTECTED
