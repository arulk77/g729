`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBhnurjxM16Of2lfWgAgW1kbjpm+D1quKp4ZrZo7x/nt
8w6sqo5AY+flWhS/lWmdFLympXDC++qg1UQI56cDKOlNLuCYT5mUUGi1Dobt93ve
miLB6sf/KQGreiRB4yn2DTIB9PFkvYJwqW4gEFE/urWvCqp2q838FE+oUblTEdZw
iQi6pbjtPwB5xj2yMR72rwmEaYO0Dj74bTFgE21/70pxVaFfEGKZ+jIciaOVRNFE
SwS9hOcvHzQQPqQNm4P4yvxeScoLv8OkjhFisybqiGPUAT0WYs0QC85FiGBuCD6a
uIIp+nEdJjr6drvmEPlD4sJd2fcqfupqc5qFuy+irBdWGkLctXQTY8OI0pUmc425
VA3pDKKwABQdfKuexds5fA==
`protect END_PROTECTED
