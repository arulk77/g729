`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN0JEdJj3wGsRlSNlcuiXddoXzXSqUXxG4aruY/0kpKEK
zw3cAmM9ObgBJetX2tTLZlBAOvZf92TAG6O1w9jlg50DN+eIiM6LY1yI+qPxNYLN
AIzvq7JLSlJ4PwadzBbkWQ715xzQsiUl4WQbnBS78/7WdHzN2dxLTaTYwvw4TPNH
S8tfkPpYAgWHZ35TlO22w+eEcGDYJoqtws33a5bpY30CxO+UAYSCWU2keKNNYKrU
icIR13YE6Adp76eDRkvVgJL7Ewb3NV5radR6gLGiAD1dkAjFBgu56cYPtt/zl7Hb
A4ZPPjm3YPwIoOye1Kf1enPX8muFUbu5dTR37hiKwK8rOXzf1Mtx6qjZz8qD2Fdn
l0fTVELCZY7xximsx3A4fcSakPShP2ni2wojl0Sb9/hHuFBlj4eD8vzVYph3WK+5
SHS2kAgUObqxDPtNi9Q8hOKYNH2E4HaaqTgFLRS3piiyyuIkzSDeFSll8CRX4XBi
1y+9pV3kHTZUjP+V+ZCl8LWUE1Kh+V9mqZTcJs9w5Mgh43e82kVm4fjRu2EEaYJ+
vR95SfbPyBSsZoB27aRgyrcq30GtkD81OqN1axZwBFLRt0sKYryGbl7x6Ijn0IJG
0RwuTpt+893GVSTuAKSvMpDuApdPVVbZX4DjStxUA63FETXXozbm/C9AhRxRZfnz
6XPLvD8sqM+enUVLXbTketgPtXnr6w0BOL+kbKRBpfsAj0tX19Muro3E8+h7i2Yh
izRfNnAjRHrHe7RM4xcGV6qYOqrxFtkUksrGK1R0mflEAoHXupm6P3qI3/4ASpfg
ua/mTh4hSSdf/1qlC3wSGC4gNrXU7fSf/Wjqdef9L1ggAvH7OtabbF0d6q7h8P8U
RdyBcKxuChIZ+AWMYpHemWScGkc8GgY52cH4n8tXRfdDkDIUHeGNyamaVdwZtioF
SNlTMMVXIIXBFtv37yNjlQkLlR1G2uu0pkJt2ME+IjLfDndyj8Dqz3c3Tt4cPrUr
sw/wyFGAoUnbFnmeOJdixcvLVG8pkFmg1lXfPMgkX9UoKD9k6dNafqsdmMr/Zes8
1x63ZDImwZez44ywJm4jWXOP2Du84uJB2Q1BJtr9B87r9QkRDBFO4+L3WHtp+6O0
pcsXGvA+M4d8ShJACi9urhUgx40p9+sERG5EZRL2gWZPRL5gHq151CLLP2fNmLMz
hRE2e/K+FUhtwzBkkV9IbhRas/8/N48AANvOCYYtYnYolWDyn2PrbQB+ZkiUGmOH
bT3IOsrbqCzULfAue91v3V8SlnR1ycJf0fGDlnAbWW8pjf7oCq872DnzzxoojIBe
YUGIqPxV1tTcnWOICzIxHGHkCfFdu7knnUQSRQ1RYeP3EmwA01UgiQ5UIlh71Uho
EEeFfqQERIz+n2UsxVP6o/iCBeVodgOD46lnvXftA5U9yexDh0ILC5NfPOeirZCB
XNfpZUjQqvowbGmnoEsDJN0gsTcpWEbbRN6xdd7iylr4ooHDVSweASk5gYsUO8V+
ttwWKYbxBtfBybk2mZ2QA657obOM53uxNVPojvfQJCk0npAeeF5qs7PynLkS5dcf
QjYSOPCj+hYRR0q0HypEDmES3DToBGyR4tm1OiqkBWfJEvn+f0jPp9RzvpwXyY/S
0qTs6Iy9nMSopS0SdlswrjqM0iK3680GNh1iP3KR6y5H/ncZqxbe8qEesi9WEmaD
N2lscYuR83BzxtoKVIXQw52ecOOw1lhYK2r2kIHvTMiupPo6SbzO11ZF+m8eqp3n
GhhT8AteopfyuQDL4/EJx5K6FGZHng5zmSdQIl0kDRAHVktcLT6NpPIBv3ys7VF1
cXDXyk7xgkiVWEhRKF3Pb4klJGP+T6oDOI1I2sj2C4kmXSVWAcxBd3rjsrWY6tVL
aezG/Z7eeJg8gbHr82ZSb/FhUn2NqAvU/j++eb+rOFXwymW2WkyKBW3VGUlHWOQh
95tRR7tri0PIoHKKli8VULkfie+zDkffAhIm94OloOiAE155klEZvAQCcEZh95wZ
B3dDUUogemRBJ7FysSxH7q6/tFD2DvNfosxE7TZ1ITpZJ0aYIApZPKo8lvE1R6E9
og1PPdGVXZj4TOBIXFealX9ARddxMOumTyTXPva+u9zN6steFbjQZjZ484RHf6ca
VxCnjRDwrun2QE56uac378cWg7iV5TqqdJVTJca+QBvaCTaNSapxh1chFDtNyxk4
+ZrKF8M5ENBPfF7MFk4iveLeHMMyQEx2neUZde1WjvGxtIIz4j1p4ybMiiqyRKgx
tp8H62PGheOd+JbdFhMm0dbUn0JkSknEfe+wir0k255RGOxUUFILQTx9ymG3e006
iAYnCoXzrFcROLAOCXG1sE4OiBJj1/bdunOxnZmLCNW8dE2kcWQk8nYAvyrDGN0D
jY44MYAmvQhmuVZa/icAHA5tvk6kKK86shkwKS5Aylh1i0GQ6QvGmM8qqgPAyZzQ
QVVycNDz/eBvmmS7dA8W4uiGoSahClwzK9bmuKkrsUCWiNfcX22o2Gt7YI5c1iZC
b3jQ9l2KPZefI84q57i+p12GQY35DdVCGjqxc8kIuSnJH7na1dBEuwKCBiR5rO8f
jsAaO9Z7M0dlTpEJtRQi5MxsZrvBD1CKtlB93g81Mcgt8n3JsCM8njLp/2b+0s1c
uoI1w0iyRKwzaeeRF8JieJBIexBk+G3XuSj8KQg4yBQ1HT0+HAsfBphyh8oXqVkv
Pe/vF/6i9GFVv5npbpvb3l1rP0Sx7NcOnGuRusI4/oQVkGshCKo7FDUZ3LkSLA1H
IiJdqtctxpUirZT7U/ltqbrxL7LLpACN+6JXXu3jC/rR7JQBDE2/IIYwJMgdgyn7
PyL6rYgyLekXk2q50rU2bAEi2v30VuidXg+80fjXa7jew9ozEAIM/dWJS4wSp4dw
PzEENj63PiD1jo0o8Z2d2Ub+tVHD0YgGpweIU9UW1iwidU6qCofn9znxL89edvB8
MNDuPUkw6q/vbfPb9U0ffHbONuYvg7bg5rpJXAfR8AoAubWcqv5DTaX8viwIjJvo
byo4UoixQNdpn8z3YBNjlcklLAk7n+NtZjSTjlWhuwqs/OYQsJUBXhwcHuU5kRYr
1ZufGhP9w2dtBRiwjgAgOrG8URPaiuCSfaP0VZxZ6SgUGSjkrK1aKPI9XyKXgvIT
z6PF+DG0ZKvXZdIr2Qv+u3fkBWfFPsFsmriCLCKiQm3BnFVtX91yfdEeHt5n1lV1
02XqmoOwRczJSo1B4lPZBvt24LdJKwwguY9UfagkkNeGoZCVoRpzCNd06SNRX6C3
`protect END_PROTECTED
