`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
DL4tUTUf/0c3SpsRjJRRmYLyHTHLrsWVVOmyU4pxhF/C+p2KHN/3e3NQUy3Vg8vg
jgae6G51P+9IIccFw7+aAPG1rRnhaPfj5u3MZX2rCBBg19DivEXAFQ5T6sC8g8yR
TcqpwOpsZa5mAymXKhihmRc56A8kdiR2adEilaHn9pKCVWl4UTNO8EOVJ0HtVB1k
JSYM45sYDR7BOEg3PkPnAb0p05isQ6UFtkrTwnuLIXgEE2dqKcSAQw9eb/2gik9j
qJgZdIUKMr4lUAjyO8hDE0GVB3PC1PDdZ+EI5wcCVRUNtNsfeMh3F7ngF+QLjW32
gxteOSsK3qRiypTK0mKk/XQNLUnZuAReWwo3Ji7en0xbOIzoqpqWCyHBdkiUebOn
7VtpeJ5xEfVvLAKdJX6F4PvZK0DI1JN4nYZT72QFeKJne88gNpWo/aEPzm/mdKoT
UFnYPszHiFcn7YSw+B7u1zziGgzuIAMGF+E67q6zwYrWvgGE4eZ6ri2VPonfzZRt
iGOvp1tqZ9UPoXTUjQ6g1sluIlhFWddo1V4TfaGoWj9Vwoi7BXITAc0G6898R2Lm
W1VMExQ6t2oGdkPQVzdA8AJQAvLQxUziIM4GWcZTcuZpfsQF6xmPYFUHs+bnSBcq
oyA0Iw8D/DjombX4ka/uC+Lvh5r2a9LLYKTDDrxATqLA7CQAIpNcmhsw/mAj9iSH
EvnHnV/HoETPYsLWBXgq/tddWFNDxKTnTOzMKmerd+lF0rZBmAYvh+/D4DHIHaE6
Ls41Ikysuc69OtNeZX0D4RMzBYqmW7ElNF/hfBACgzSp0wQ1TQAB1Yy6tKVCJBVA
Esfv4LYbsg6coz61SNO/MfH+CK7g+JuZC4hm0naSu1ELtsD3D/WfYF85Hu6JzDW6
U7fQwTJ7UesAGr0gu3eqCLpcPQj/pd5MhWobSooaM/G3iVRlf1Hrs4QVX+Ljh3fM
ZMj2NmQxL2kSchSX2XQh9wKozLmBYPCvkmhXLJw3wNbWvJVrnwCw1ZmUanURv4ZG
GduH+1v42hZnwZtoZXdhmNZzK3oCFBQekuEDnN7qfEA=
`protect END_PROTECTED
