`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAdEdbq9p+y6nkHSne0fb/klT/BK1ey3TKY/reaqmvFku
UIuKpSR5DBuqL9+fa3Jc2iOGxa0fuZo0uFEJ0qt/hXVt7yxpcmwFB6wfF+18MeOQ
63XbD6IBgq6frye1b/j9H42F3No68a5okRtGpeoZ5uBh0kedAnEQ2o+Fg/laxeoR
WX7BvIIZeubkvSe7Z3dqbWEZ/+rNwFjBb1Yi3qU4QPWGNsG2N5fLB35YHss1FP73
nok9ApRFGX+oprphQmwv4zltFgZWX0icZSrG4XYfFsE8td1PFrxefTi5z5EH82BJ
d2ajXD0zPIZYzkITQBkj5kwsEUzouhDX7YQ3NPsZG/CQ0ot6zMXnDfFmSTagd9r7
R2hmXFRt0EkU3uYugca94aV9y4i8rDLaW3MvHeG81x6/giIJMtMvojlDM/1lQQlP
J56Rm/xgYzA6k9wRJFeOim/2lV513LaGdglDeLsS8XaCXfDT4ykkq8hXk4KxSk36
tbwZUIO6j/ccoKxTNLmfmg+EoiPvHj8JxCiEm27sE0WF6hEWTX/hs/55Wfgk/n8f
aexSyuGCnfnNEtS7WB2Y4g/ORakEExooNFDziTqF4X1svfLqc5Nl5Lax76e210Cq
KPEP9XMO9yRkNIKo0Dd6oNyBeOj/FA3zL0dAGLnNYf3y6o9U6tptzmlEymEcM9i5
TjblAugHwo4zQ8D8KryLSV/a0AcFELsIVKMgL/kk19lCqDkEqgVY8QJEUaevKZsV
`protect END_PROTECTED
