`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAU4o2QjYsSh7S0wySLi4Vr/NHnQAarMuUr5D8rRyZlo+
TGhtVYNJ+Xnhi0tiM5pHdcS0bNJ/vQXlUB4AVzefNIcvMGRh0K3Io0mO+umYDGb2
1fuqUSGTMCgSzqmDq5kXUh0yJdymABIh8Lo/QZZCHlalCUeqOaDi+owC+Q6+hqz8
NRkDfKe3vrjPoVjKRsVRWL5bQbJ0agEjICnHn+FvzP1obFkYx9l5DQ1fyeCzr6Rn
C4DUquAYxDegT5XreRUXBVTeD6dR8Vj3+OZo9LvhVs2RwviBjUsfle7/fq0WFYQ0
0xcOKcXTin/EcBLyKyuAh9t2TayuYH6Zv96SXMtMFqnmAkN5Bb9/WKUmlvMKiRIC
6TDsZt0l+cQEbd0o9eX5zpMyup/3YBkryzwXapX3FnR6JqXXLJeZMXXlKtYCcdLl
TpXOWpmOvMmhBKNUb0qY2/UJMkQm6RbplA/r3qd5OxvwkEgBxtowe0aP/0c48a+x
MliQhDMslQiGz1eY23KuhKUBZJWXET2TsmqgX5GhB68N4Tce2MQgLqOeH0Wd6dC0
gQur0nHLlitdQQI7vFMZn7IPdBRm3PTwhQDHyyxAG9gHVV5cpdIeVP6IHAKUh8Me
i7AZ5sGUQqr5Hfg9Er03MDzr69Cs6SKa5Djrf506sp/eCJmphwQVjKkDRq+hVmUU
VyDBzvTtu/3PlmgFR82AGV0m2O0e6TurFPRkl9WuTkGM7RX6mGQOsue6An1D6OKB
V+VJNWqn9LyZIfrE9WSGQHvW2IwkHFRL2HVgO6WgQKp/q+1PusqhJiVWJt89oSsO
s7raQvAo7HPqdIoTzm7f9N6rC94kHbRrU8Mty6xZgoyqfylCO7jp3MKUJkTb6Hc+
tRfKtjzumkC9c4EBTrDsSz4a8myt2EG33cxXJbZ2a/n1d2mTRxWEFIj+psumNnub
M7iX2LpAEzUCpPawxT1Nr6BRNRY2vQYbU3wklAoLSiMDm9ZBDHC7zCaCPy7VgDZ9
/peOtN7utwgLxGFYr2tShWFxaQ0zuKSmxvMqP+nRBmXundID7wVl7MAFbwFfawxs
g0NR750SaILxdxIsBhL08J6fI9PLsZv0riahQuDn4/a3xM5d5Kj3+gpSOQsStjIJ
DJLVGusGP/J32RRkTgnzAskOaxbYis7I1Jd9gLWhykg+9yRkdd8VSf9dekrDd4k3
577ZHVt0mgesk9eo+moDi7doNWY9BG/0/to43H+M7McyEZcl2AkWIlxPy0+qLHxY
HGMKZ7qyxTXxBbm0rj0lwh5OjJup6xdcTXOwD7iUZ3rzpWce98rpcrFPFtIcT/3R
aUMSTyPhHlx/sgAAihiBczukuRgXnJELom+851QjxKlka/3wNVEeoBtE5T0hiVVS
1AB/DUHnXS2MhGpPEXa/oK18kOLiEEsd+URBCtr/HQ8vGJgaX5tokaufonPKt9/b
QXHcM0ZvUh5CFAChLswy8G+cxUcYMqICdBw4GydRfAvKCSjh0Fhosun4DWBI+aep
hDBcoM1FdRCCUeqegele7T7hEozzw9eBJ13tsKBuNEhDNTlK14sQmoI70eMfe2xs
YXZrSrIu2lRCnzw9JOMHeNj5Yv8SBgXLwEmA1zpLKm6bG6WbwEDliLC74u7HQ0Ka
B4ht2EmPZa4uuc+Th+sAopQJ4Cu96Ag30JMhq5zY1KSxeu86FQuH67FZSZMZigie
JrpurLtOAJHCC5nQs/94Gx97pMrQ/1pBfuLMN98u/l12rQ8sok/JFiEhcamJuc6p
rUJmVz4LV1z54I0icWUh5GgyrbrQcIoBhu/a2bPeK2JudIbDryS5EaYDa9TAXi1F
finwz4G4OTcVFG6BhHdBZ52EbTuA2U+RVM9+qjjU0JsG9dUmDX6kHWyvLmnxqxXK
WCrCUa13kxp4kvwSSGvZMs3JsHZGCC8srYHv+Q46n7AkFJAfkPoilXeiWoUAjNJ0
CdnlpcnX77Bb2PEvAQqiwZGCI2TfQ07uHy1wzfEahuVnYhjOGAqriYhEL0rLLBE/
hO8p03P8kbvh+pTddlnPyW6VMSDJO0RXVHFzSrbA3Q4ZsOMQqeHGJZ7NE4/sv6jU
sLAccIDqB+ZFE0EXr1pNhGM8fUmIgjfJma2Lso/1UQ5Fat2MqDvz1um1QR/JipjA
K68rde3do35ZO9AxVBp7Q2RjW7hl778Z4dIqRTHBzCpu3g/l+uPTaLCFr4pz8ZQO
+eAnfKyEfVTnW0gAnbdLR+xMDNm5DqDumMNn0ZPrtJekFAHYZ4tTLTdwmXsPCFaz
lniRIn6mMDIA00JVQXDLUz9xdSY4Yv1aXBkMtzZYO6uqsF+nOxExKXMjup4JTE09
T1btYBU0upBMUp428XswHdoqPFJ5+qYOVE7Qxr7wTt32x6i1ZsufiXOgpO8Fi99u
bmLM6SpewMd8oxJAkqvNvfYIjQFJF2O+5QHYgHjZJP+p+QbgKUiLT4+gRxM9hJF6
2OZdeOgnO8GYQLmsKlbOWj8S1EmF8YkJp+GqcBTAE4f3I+FCefyAXOMtAdlHn9wV
r0FmRwQ36kTNDkq0BwY3okGKg7eGpnNv37g1CzW1ngU+8zgzoQGYFAd+BoNIT3se
SYp/FNu1Mj5ySvBlSOjUFKbt11Oo6UXc7pX3j9mY/pOT988+Jx7IiRRdTeMmQaQx
H0oKkCHycji+BEPrkQVHzMrOsuyVfkp8g37mBp35tBk7TjbHZF81MFa8gRhw4UnA
3jvarMOwDOs1iA1a9p0CLAus5eTI6JQXzQUCMYiq+N1sOEVOiIJv80d7SGzEyIX0
BufsLsfJhV6ix3P1eT1dzvKUAxA1+XWnfcw6qvq/Yvl6NnN5+WUVJ5rOvvGtwJNp
iR+eTJ4Rq5Z/jeo4h4wi6Iu5LNgsDs1lgh+LV9XjfQjj74G0U6fgNLdizLI+aMoG
lQ0GroPjvQ6fMVwoloR1/AhKrgVdx96djxLxFg5Qube/GBxrtK+X+vgAu1A7+fWK
PyCSfiGOXSlB1DLC1qPFiZ6Pstv09THsyzGltrtlzYrfG+eaWNZgazUyCNu6q+Ub
p5+N7ztfWVpazkAXTieo6s81Ou2Uf9npI3BDOwuzfHueUqIN9XCd4F3yjnsqTXHb
v3J8tq1RinZXUL0IDEiskTmwnIxoXjyjKF3sFLS4JOSC4zc6u9vmCBNtrarBL2tg
MRgfDE/1dEgfH/XfiPZXRwzVQNc6xLg+elA2qZ6OQIWOkKLnzP4/sgLlVBVxNQQ6
MtjrUd6wvYA2dHSnK5kvlR7J4FPC3yN0yVsVUOTH8/1HunqqB4fFRq8xLqayxzp4
xVPtcy9HHTb9sTiLVVcijn0qqUVNTcnw6CaQAyjq5rq63LtUyYVBezvRG9bDGk9r
HrDCDMmidtVwIIyd+riBsrIdE/PdcwTAjS7CZfWVKvI+ghRjnRZ/YESCJQO0g6Um
6QQmQALdtY7wz8TWmtzrYghdAGaz4/rlmh+Gvs3WFCsxa6wGDTQk+mZOZUPNBNom
1DJYdrribKM54z59FYvaP/ZpEQqvE0r+Xhl9BheF9LOfj9MhwZZvaziVc84sQQ/z
BxuFie+0ntwc/VrDLkm2hwIMCik0y6K4ZbAxtPa4HjJca6b/rpFp6V+aCPjLtjEw
aDbS/Uh9/47D6YjYTh1To6GQgwO/75Z+ezRMzx5lhaNUhwJSKNh9SWw8DuEZgk9o
KtrjbXefFV/TEI5avIlvC/Iia338tH4mLTdtCKAnn6Oiyk/I+lr7A4wE8Y6o5dvM
qYDZP8EvHKPcM/wEl8TiunBGIXfTC0nQxL+0e33SkBQr2QS1A99xcPbhF+Xj9k+e
LzLdsjwS36rPlaEvoLF9s4u5mDXIf4HJOlFbNqV6YsXujn+uJ6Fqpe+LRjJDtivx
H4klVcaKFifpoLSUPegqvaC0D9CUSl7okncFbwJ+2VyDwcWHwfOguiXiUZIx5Q1D
OA4vQX48EoqaYvGcnZ8yEZyx8y0aX6o9/xiRxumyqKCwr2S6KCHrfEubO1ro6v6t
GzX2rg8hkJUtQcRGApd9J3DV9cHoW3b++ZBvUuB4IUi7ZeusNhYAvAgpSnfw4dI0
grLR+5q8uHBkyW1SOrY4j35vOhCDxHutjhS+kq4uCbDQA8gSxsCqMlufkZQG1QWL
d9BexbVs4brktlRyzTibixCqajDF1jqmaS9BLzVYECr7NBSb4LwYdCvbQ4Vfhjzp
Gog7YzI/R/cswF/WukMX46M5ocrAGwuZShB0YjXrwU08vauuTPNiiu3cXi7s0qld
/NHnGS4U8c+Mn3IhuXCT72CGYkO564AdZXJtoZ1gWoYHkvDJp+5RbJaFWoOYf3pt
u2QBZ0Uw0faB/Rg2bkuNfLN5JwERYuRaqL5JTPeasHQKyA9chk6hjQD45eJK5Wh3
+NTYXg4VHHqXFE6oTIub/UGHOyMuJEJL+9wVE56eMDfQNG4U6mgWWgfGieXgJlF9
3sceVUmSbDmXTzSawyceLNvIDupAZWjv3dyJc2sXQ7S6qGw3b1XXj1J87rKgNIoe
8yDpca1WL6R1ExcioHAUdIXQ26NzmRjIDWfQZj7ydXs5oILg9lpF8gEHsiIaJcws
8XiCXjALoBdeGiAk85a6Ee1O9av5CKEzezCna+YXixZuUg44XUpQLmlwggcKxutx
BWBUjiVsTo8ae9umaTF0qhrMeLUM3hX1mcd6d7NvqESkrqk5d3i8sIsSGLFLPAX6
lcb+TDHCyrmEsI80JRWUk6OlZMevlvLpvxlb55MMhWgeQUxD7N7u62N51TOqPjCN
OXdEmwKmZ93rKP1HvMUpUUSNhuP4R9AGMdQDfNO4nAs/DKEiwE0qar48tQSQb4qp
NGyZ1LSJvZfYTLkZLV8YJ1E/fDnlWdRWTk7N/TTr4VTyJtCM8KcaWVXigAXmki14
rxkeZRfB14NBMeSVXmjeTTOcN3cclweVY+78Wr+5gcXwrxHn/8RnDHa2ZxzcG+lA
H4XpOIZ922RdXJht4GdQ0Vp+egoNWo8tNNzEz08m6wBktY5oXBVnfCn8opYlAU5l
H4SdwK81fFQli5WqSWsVFiUuRPyscjEZlUz3NTODxtf6sy5U1v7f9s6FmPq93/wu
H+wECZaBv4s0k+D4dIORnwwEH8ucq8dKoEH53QlSeubEvj5X2Ymqt+5QwUAi3sXn
+8TC2dFsMquipP1qc2vjtTQdIcR096Eq1tYkTaGRfdLqlpdaadHQSk5+v55a3fs5
tzVFfaxcEKXcx1QqJMRENLKAqZCWRA3jzY6tromlawo6c5fMb5IRTfwdphgs0rz/
Xb+0XkXPjystYVIDB9odkowk6Iwfy8QlYEzh7gwOrgO5jYOyAXEUlJZAOKAi8w3u
OKP1jotdxKAj3z7sjDr9IEJFIMU+B29XQraVZiomSwIMujF/uMDVGurt3+Nnqy+C
Yl2UG5bFYWs0eu5Y4/cGVUjH5zTTwFx4d4VlmvwTtiIr7A1JWKZdP3cDL5hnQP24
/8E4QdD+t5Yd0ssY8kril6RvBQ85hLU+KOf3zcSfY/YX5psnmug6gSFr6JSdS8wb
2lGIYPVmOKYt6ZxUZS6LxDDiPkmjDAfNkTAJi+3fGEISVDpNwWDGTvUfcNBMW9zc
PD4ixWr+bcDp0Ubk8RWyUnjZYJoFRNqe194s6Vl4HIoPECbVrWW8e2Ywp5GTcCHE
v46RvQ3oUWI9TrjyhiRByZEjGbaHjrU2eVDnCRVw/FSiyu2XhOv0gPe7x6IPgq88
0M7lBVPd5SAhC+6FstJE7XWQ7O+9Z1Pk5J30JHn7HJaP3zoQqq7C+UquMiFkiAuc
MxrZsXJ/3yGmyvjpLBZ8NNXO+nXpUaBIv8JCDwyaZimEMKtoBMhsJUO6Htcgq2zK
19m5xD//SWsz77CF8adccBkKGNQmeTEyTRnf0yn8Rqn9vFaQ3BMqcvUB0k1X8pvt
F2ytynsZQzBh/0qivo58myKQRaWMmWPsUdQicvtM6pAb6yu0Lgpyk7Fav1oTgHiM
zLU97xKae/ObQzXa/9y42w==
`protect END_PROTECTED
