`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMHbk4RwXYwKu6snTmGXuPdlj3J6QQa+ntR1RFiJQBHA
B8/8ruD7ku9qtX5Kf1k2yVpIZrxRBdMo3qjH5DQgMtc4bYMD6AbeFu9bju9XiW1X
685YTaBxzJ9fFMHfIRsW1xc86f2ihI86Yya4pHYbYlpvM36oSLnEKHDoP+zZITgS
G/nZP7jyDR46AxUEt7lQXd6V1TRIxt9VauqoBeUFt6/j6ylCcmpsyKDI4fpb6dV4
mbCO6fWTpbVcOQI6Bm/uHGtUxpqbHHfsAE8eSY6GbTPpiK4+acQq4dqUXPHvtlwS
20GSGhCAtf6DkNUeSK57vVF8cJgTe9F6AePIaILKsJEbXyOzG9sZ28vLK6X60SQq
c31b9N50Tk/bea95R2Y4pNraQgud3YINGmE8xU+dtxPLdfMg1jkGOo6sNkwprJX9
UbUtfJjy1xyLxuBDduJHLjX3ufbTF4a55bDThRuSICOWB93IKpqMh5eVrwWrURO1
qixmz3Z5UMSTH4rrgLsGdv77gaejY/+PKlWKcScMnVYaN1FcvZpUTdRvX3l7GVgC
ZPM50Tv5kilOrzRyV7WC88NGk7JSLRen0cPlaL0Ct8vEzqo+2JZSwQqaswFf7xct
OMOPRVHeJbv0w+/6rQyPpO0Io4tcgYYHGx/p7qmLN5JiCbnXBJpqE0W6s9q6TRFL
`protect END_PROTECTED
