`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JS6Ee/OUguv3S0KjECptSPwLXcNf84qpbimX2OFsrdXIIrtgvw8YlC5TnF/Twvwq
Q29ypVZglRezoaP5ab7ksHkNSGW7++rC5DzWJBaUD1/0kpyhZJdBMetNOHfG5aLP
+FI1Wd6FwsaecL3BjJbJlroqcNqsSNfJ8xsp+YY/3/wp665jdnJW7GAtjdDmDfJq
JT/9/WrtwgiFgKAsPDIUMG0z80mzFHvFYUh7WeQ6Y22W0yMGWJFbzbPUJ0sl0CGK
uK0WfnX1N/TSlBZg0ib8AJJU+0k3cmSDOzsm6OeoABoGmM0e11RnrachfmGmamj4
SFvJ+Z7ELVXfP5zYFzi3nKwHzbIsqn3R6eSt3sqhJD367Z3nfoorywpQl1+TFINd
HRuQ48HfzNhv/MbHDuwIm5qRyqTwtbxZnCPYg9HhsUo=
`protect END_PROTECTED
