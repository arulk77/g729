`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDGuxPgcjWWq7MVT9u6jxapCG8KpZxstn8WsAx/g25e0
xobdHQYKtCzKRIL9Bp3LDQeqvECiR260JR5wd3RDyFqV3l200+TcvqcVhMQ4mE9p
1pQ3jjjeoJLncosjqR2Q2ad0MQwnTAkFITwqpzYOTYAcwvgK80yW95C84PLIl+Z4
UcR17A9bsTpDm/hXCKJHvQ==
`protect END_PROTECTED
