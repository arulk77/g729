`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHjWH3Oef3rDYOcjZFDXGzTZcsyGW8crG0xnKui2dR2p
yyF61jSGOsKEfOxDnakPPzNPjb6pOW/4sYoeUvXLnIJ/p8/7InArbAAWn5TBfxDv
fky+4jFdFfc5dNl3Z2EsKFsNWBI6rsC+UG5P2l/EBlTF+VylrwVin/qy1hYsNlvx
jTtNYNGqCObf3MZbHB2ePjt4r//G9ZiQhxcfVuMA53cII4j+CqhGiOd4SEpXIJJD
jvwS88+77Nh1BYO2d7Yifg==
`protect END_PROTECTED
