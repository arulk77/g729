`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4y7jqWJYSyvBxOqD2jLzWdl9gMt4sMLhSx1xChL4I38F
lrsVEEwy0Vy2q6hWTSS+zdA8hFgNA/0twYETVGhlfAcaPIdNR7TWUWqEr1GJK2ev
zRxQrvIpZ8S/Vpnu0SbVWVJw0dwVw5jRdJ8b5adBcC2sl9jtdnNZgIsD9jbCoVq1
AZ8ApwpnCbMBc1mHlq08S77C9lmZbrV+tykJJaJC0WjxYxdk566RlWQCLI5sGqma
CMGvMzVV+22QtIwAytf5txVs1YV8ml6/4++0b3V/rN0=
`protect END_PROTECTED
