`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJvHdiNmyX8nCaYCkt1LOWpJ9wnUBNoFBVCh7D3wKB/c
X+KIYLMOrwlSAWxmfY+BcZO/58zwF7G03r4PPmU5YT5bMc0kZ2Mm55W8EcR/tbaf
n26fJFdqTJnWRro6hbmNvx2i/3e52dkUiDy+1sSHmW9sIkcDVzieb0lWcpx9Todm
vHXlkX5UwdXNbvNBpRijaQ==
`protect END_PROTECTED
