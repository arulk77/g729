`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNcXsjI7y05hazWrV/+wpMYhxSFAEae0kK/Trj0VK2IU
XfQ7RPE7RDYkWApV1Q+4N+yc3WGrW8ITvQ4e+rFnjNZe7uWzUai+FXlAXzKo9HPc
kZvPwkoNS+87dkXWKOC3CwrLr2db/AaFJgrHtwf1ltfkPLVMDJBkLHeZEDkOZOu/
XG41Iq8e0dfvrNcHiZg7L4OKmmx62OlK620/Pqg7gDlOUP7uZ23aOpwOswPP+Sea
N4W34MmeRBHNlTfY4zQ9ixljCjaaajrpsahSP2Dq75pOzGATwQIiYZhcmkw5rYb/
0evw76yCXeGn1r8fbnt2q0QYXnvG10Io7HbCErgjGFmsBbN/sjIOZbrykR/PkNxW
iPGu6V1T+w9c8atm4YNmSkrf7gvn9PGo02y2FnyC272ycvZelrjAn1zJeugFTYWF
ftSLPhSRlewBQVZEaiEvezdT9OdsCM/VqUjjeZM0nBwcmB4SjpuTN3VftCQ1Jlab
`protect END_PROTECTED
