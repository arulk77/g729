`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAbvZwQaC0tKIcFOxajmj7EmkxTVxB8j7TKYbrGEtnGFv
Zd2IBC6O2+pC3IT8ggDK+41IIqu31cKmtoqw9gJfXCeGwOGiObAIP+D2dszdJFOX
6Uv9X393PMUidB7+xjYaM71BKjrOd1PuVBsyLNceBUWFOvyDTalCTO/XtBxhgSS0
GLLuC9cx226o0g/IbPzq/OLd5MMoS1BOEmDb++qbYHmZnApktAq05k/n9a8DISUg
P0HCS7wPOjMzMaX5u0dV7bohKMBu4SZI9HID1I2CzeyQVTBocv5RKvW6WlkFWo6k
KfhOHL7pDD9WTgmYH2qKECjGkPLmjr4DaiBDEK9tdM4TTTXZQN+x8kPPUxOpi/UV
U69dxVxVagyWMEsvkloFYtdevYbik8rK53Im6Xpu8u/1qxM/bmVHAbO3otBkyki0
n5aURgkMiNJfiAT8pq9PswNper02/P+S6WcVQDF0t8gpR87eynMkOBEBJpywIFKz
DcN44oJ3UuI6Isbfm/oFkUBTs8qhnqiJpc2PXLcO8J57+t+0kZqS+bTqRzdOuJuR
1j5WDOxxNumn3yoLBbzU+ZTAzjV7WVNMRmny9DQi/d/vFKMWivlESI6DYXuhTyDU
r2coz10OOyiwOm07iLlNzg==
`protect END_PROTECTED
