`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKnVFStg+ERgFfEqxMZrTuE2bv9xLeYpSIbf4NN/8R23
gIK2poXJU0A+ko/VLRR4iW7x2ZzzVoXDPFhctZ+3mHnET4EwDDTrmAQQ87QqiY5M
L2tamOJGSQ/1KEow7tG226yLphdO3qiuqW0bZRpYwPMq/k1E9OhPqK+Ul6vlbmaf
0sTbMvg/kpYpMK1I9fZZFfDYgtWWtEtv2tAz4+O+Bdy6S6e5oQRmPovAjxFxEEY+
BITiXTk5j16DnvPDexpzfw==
`protect END_PROTECTED
