`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAWCjxU76qpB6gb8ClHKdlsqFriLi54SIaJgvBivviZc
fHr4FuLz6SLvTonTP3Rj2ggVzpgCaeaKeyGkQAUozoPe4HDpDdOwCD0jlRtm2pkr
NOJEgR0apveOqWbRoIT+SewQlyO6AFH9qDPPqvG1UrYHlxIZNXtDdIOwjwOIIvzb
fcBrpVM7RJXqPvKSHHz8plHSaQWx+QDINmMa+mnXZiM8TKcz0xMtgCtkiac5s+BO
0+90csfYK/ZY2v9IJBeBoWIKP0NHK90sJc+56EiUU6tbjTARLnM9A51YUcZHVP51
JupebvIBHdFvm4vBfdGLmI/JuloRuRePOHuLZJyZinfHut5WZgvBYZCReY5bDpS6
0uLjcQ26KYMjXLtz3c0OnmGDK5n8du+c8u5yy1xwol5bEoGnPJ1OsTQj5miwbFXK
ZiCJ/Fb+6NRIPTSiUF8JO4+Hm9l+QV0elolR9hdofXR06/G7bC3OMrvwnXVlzixO
`protect END_PROTECTED
