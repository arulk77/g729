`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44LnZj+aln5hxf2wMf9qRFtnY5q73DmfdkYYhlLmF7Qs
8CPs3wv0IKn08aYoRKejtN9kEmXn7KgLV6PO/YpJLbcNCylHoF4iW5uyPxnQ+qTx
Lpu2PUDy88nwyfVmwLi7QQzuGeJTrdruV/U0LZ1YzbXKI2fhX3wEOV1R5PNS2ML6
5s8Sd+3jGtD30r8m+tyldy8QTTRZ/8YVbox97/TMf9t/Z12Pta6YkiXTOLpvKs+G
GjVKXTnJsD0Xb7ClO3/73vZ66V9pL3OWgRDcUT/Xbe36lv8pjvpcy0/LMX1jp1lj
7VEA+Wg/hvp1RXhUOGw1/pypk5sbMcZiFoP7oMBejH2WA+ISyJxabC2ObvRVRVrR
WcEde07HkHD+0vYUlj3c3w==
`protect END_PROTECTED
