`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
p954hZceMfP2n08vaiccxU8fvMzNL6xSZLHO/PKNsPKCvuOqs5+MX/wQb/F+Rxll
+oA2nyNMJOsV3OC71m6mLjQ4GAEj8XB5ifxSjLnb2ThdbxqKLBTYMLqh6q5l65zs
ywLk5Q9QTci5NgAZoNsh9w5wBZIUWOHL7rcFTz0HOkcY7FMB029pv0ZiWnDDU9o0
/bFkAHHVYcsUvYf7ikDCS0L2KVqXJ3Gu9vkWBPWTyQ7bTm5SulOogPXde+B041GU
dig3u+nvnI0g2HT3IwTwiU6M0dEbmYZJw2PknKRyDZjK4rniNlY2KqYjnVBeTNfg
X4gBHriiRGn6ebSA2n/Ye8Ke1yT1pyWmMsnGvxepymTsQaE0x/sHswSezO2yB9fW
972dPTd0Q6u/Lri3ANxbXA4OL0h5Gr8cf8ehqR4VF1wghcXv1Tg2UM6HaKPemqoo
fgx2Lz8htZUVBXZraBHztw==
`protect END_PROTECTED
