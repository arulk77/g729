`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aQrPL8uo589wR3py0aQmlHquChQzgg2Wr1p3hpu/v3pf
FXf16M99RhIpoyTtbLTGUwIaLHTPEdSrrj0ztCmLRWc51Kof8tAluC4bLt22t2OD
o3uTO0SPcOXh6ZAyVfcDwxSZE1UUKj2BcwENLuyovAqfqLkD4OPe4V0pDr5gMp7V
Dtn/yjAm02yKbxsL8Xkpb9xGaY9oYK+knJn5dZMX49ziAjPxCbBOJuSNCSpaLzXV
F3WyGe1Fo5gS70NXHNV2q9fhUxpfqQVUFZRMC1aGN/D/8UioM42KyelZyQg9m39e
8fyNhIPm0FPjFSUO5KHVzn1nuyf5KS/LNgEQb9tzrWix8WTHFH87Y4X6m5DqIUuj
ALtKTuZSJjJ5r5e23jXuCantPeFN8GboKF2GrISKh4KlSGb0vWE3ocqWd3zRNfWp
6QEjG9NGEIZENqUhiGVWhS2u9/zmvjKrd/jvLWkq4C1CsP9NriDphFP07XNXTTDQ
jgnNnJeFpyQmG7GYZlt/6vxt4bUP+CWn/ekjDua/acKfA4tShhkvo71BPL12D60K
kQ01UqLea/6TTL4VHQPrUDUJ/azxMYyH1R+9bey2ywLZpe8tIMT2wsOpR2b6PLOO
vUpAlY/3A5H5tBKlVxFJAyPiqRZ6ATvn4TZqSbRPwrC3oaGY24Doyt83vPHvHA0M
Wp+YPs2sA7O8IB/gDla1jmPcEDah4OFMEkWp+fqf4Y2K/CbjrT+oClGRMV785m/q
EwCPHRXJrtv8bnIAsvTVgah8/hnMag6HeG0XMAqauqxVlbgqLmqS3zhOxk3WBvRw
4tvZ/9qfFCdew7Dk9rsH/OHN+rxEn6isy9ndX+XBfJ3r8QDUGi2dCtHNebKFEDfV
+LRokJonYvalbicdI5p9/5DHyHnTyuy5g09ezlcQgLZRlcg/OCKgOCU+S0oIL1Z9
QdVcboUSUlSdjyhsb+nGHPp7CMKrmjhiWM1swxgCq4mvXAqAha2hQBsM0EDTTDyD
3xRgJCH0UrRC8Cv6vRd+AdfqnGr/3gbJ9lOCVyaV80nu95hbUxGIzsILN4HoS4VX
dLKT1ocbHOUI/c2xdWPm2YTxNifWfJjFk4hlMgZlZvw07ATvMUddgD297ARYsNqQ
if823XKos0BfkkSNVYq2B95AgLXD3YWGyrKszGg9/ab0osrnyEHJi+tM+vk5ZVWN
os+dcPTjuSj1BvhdjsSX0MeijV3irtgszQbJhM9YUppIJyVf4TnSUl7expkAkQxn
M/r1siFsStCTNNdzAm66ODfk/uwjnsOUby7UKEgkWlcOF8Bw1sMjLfJrEnEuDlwl
P8vImCqVMGpZr9eaprtXe/9IJLIlfqhWVEnx9jNI/Fdl/OsEnzID2U0UKp8cDGqc
lMy9RdJSccvI8Mpsr0mwcrTcOtnZmDHwGAATW+/1DVUCwI3yejlss0hCdMHiBsbi
UO2kYGaIRHnIk41fFfnbGkRtUeZGWPb5kYJqE40CVifYMGHHaBiggR8sXgp0GPxW
g7F3wIHxcY0o3DVIHlpZYQR3IyJ0Rhld0QbJUANT+lVl4oOBopILOoWJquS1a6Ef
+jNLcRSqRFguH0B//rKnDffgdjlNWpv0mATFMexb6V8FM2TJjYCYLsLfkE1i1WIE
depgS6gHmENl2O2JE1h6OE/9cNfCfnmEs8Oh49YghUzaE+wm/gEHtRP4w89QWdi4
PDovmSajQ7ppoCBvWniSRTyNZL878MaVZ7cuGUB3JOIdGmssuoxuoEzsS4F2QoLy
S+6ZKuTK71YMqhg4xSUGqjzc1yxQCEIw5pJ8ixSo8ei/GByn2zFOwTqyfss9ssB1
Lqd+SAFXrAoAACpJL+VJCG/EB2GdYyTG81n6EATIwIHkqyMDahB1+nja70mYmxg1
cMyLr7huheTfl/CfAJFxLp9w1MqMOIvhehYrRB0M5KUTxZnVPg5Yk5L9XMpdsJlm
24oNNAxxJ+GWz2ELj1j1F+eC/m9Is4B6ua/phaHDQ3n35Zh9ZfQrzsgJZrj7qTQm
dPyPeCjTFM7jQ7mhXc+6YiLxoo9SBzJCRNoDWhtHl5hhgqoIGWS+kUjePePxzzS9
I1O24/uZuwZTtPMvTWebIB+0axd5qf1E4zjVQmVSn9mBC71IguqxQnDR6RTR2Ae8
SeLIyNe1o+lXoiFJjqkdjFH5ySQWgrG7J4AX1P/BlpL8Wl1exr5P+Ut5mTd3w13t
1po2uDrG0pY7GjFi4tdPPn9bmKtDAY2ESmDr6J2qtK1KxpbOZEIrbOgM5FW5KjWI
xVATVQjmOkkumJhpK7poYUuNvrCyR5kxs6gjtJQyYa5PAJj3Sh3JLsUdAPlq+IWs
9RKjonCmeAEl0xKUWs5k0irQfmlTnPm4BryhKwpblIhWGbX26d7wTLGdTWOtW4qR
uRxmfcpZl6ZdcIxhmM80DkCUlsnit2/G6u2NS9ULUPZu9vyc/M+VYcjoMw0VKmnI
eygTRYsk1YUEPMx6aHp3tw84IpW8wUzT32fHuU/4jif5xDgZP8geiHR+DSyvOATN
xrf+cGsPn6COxMHXxbcfBeBOQLE9+SmEijV6aR43aLNZMddG9QIwAZeLuiz3LS51
3bVvJjVx4hYIFQZnmgaNZRTsWtgfcvj1m6tAr0tOJy/9s7KfzPE+H1Qa9JS7xraP
tmMFy9Rvh7mLBGj0vEDElg/l2RPO8k+/CWuaD3IvLf0VR4EknuUs1+xFZ9R/V4P4
iOe9p9bcWFzYb1AwvNPfIJeI5uUu2/W/7jyKQE2UfBOHGxjK92TBgNTssVyPsTN2
7rMk3piBi5f5wb5Ikp+bq9mAgxXkPXzRLto1wRpoaRhSu80i1XDCcQ2xvI4hmikb
9T/jT3594aS/ZOe/RwLqhOgrxvbzS/cCD2zthPsi5yNZZRfuTSKQ2S73/Ff6ISk1
L8cEe87/i5uEGIRuk4Z0y+dmP3asNsEl//ROeDNOOD7W7JW43q0NmOC2KV6IsdFG
4SAPBGIEsDGckCwppWFixKVKD7PZwvb89NUU3fgeGwz5Jf5pTn5PsY9B0XjTrAFl
YZOq/4pxgUNyRa+ooTfj0GueOZrEpO19NUEOBj1JEsTy2+XecZB2kjEjetf3yvI8
JLvogB/8AIWCPKQQCMrepog7PPyuvs218g6/xXqNHqyL2iuR0NUkuf+7rlm3CqEa
wPfmwcNk1Sz36SIgTIgVI7I3GN/ZToI0c4+zS253koA9blM54RjqGKcVY95PPWvl
xcW/LlitbycJP9YsT9gMVtF+nZ7spu2OWKRNAuoIytvbZHPQr0/2leogv6jWxJM5
DQLEnfkPmBWx/MsJTrGe0Ld4BvE0xWsZxO2ekrNNlfFkLJDdcrtsZFdolee6eDbZ
zuLJQOcfY+OFPmMACjzYs/SPfTWei07d+kjjOj8G683FtII+NcOMzcwprgy6slid
znn3bfr4FnTMl196RL96A3UStICkP6HWMCa7cOaV2dD+s1uJwI24ghoMq1oFOK5U
hO7vrhygmz5ar3emW3Z608gytEtYTG8iklh7rZYovrdg/eKBH8eGlyoe1BQ9oZom
dh2pqi2gRUXrkK9vDymtPUgZVd6MA2/CX7JZJWtlTdLlKyR15xF2wbeGYeoJUPqx
mruiBwRRrxcAmFc6LuOhuqdC9JhKZU83MM6DT/D0A+anJof88fKsvjwYREscQ8pm
e2ElhUrfzyH7VDdBBwMuB7wSu8agjtw3V/SArN3PvV42fpQCqI6VowDxKp7SGFy3
fsHUS57RQhegYZIlpM3Ona9hlzxFNG7HYCnAkIdCMKSIuzrBh7IgbdKS4trupj22
AVB3ZbbxHq2LhOyzJiv62tkiG3xnTvmfApyj4w2P6jZfbIuplSjBVY6Xhm2em09s
`protect END_PROTECTED
