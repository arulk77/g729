`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGNz/XCpYQNc/g/IM01TnI83kLD8z1t0XM7fNpUhq5mG
+Rwgkgw94IN/7avP0mtyzbCGGkMdRRPW0E0Y7N1BhhJvWjvZ4lVMJlG0vnxsyWDw
2FyydT+D0qoKmfWNevxjSds70AKgpwKysLlR08tLAi7Mw2HjbwiGXbw/7KZM25qM
uE4e2AFjeay9KkXyWymf2ANiK458qiiUUjEA+4yqrBnGVe18EQJZwH37j2+rZYeS
hHRkYrM9f25FsbseaDmdYbncUTuP8hCtVkJ/wG2p0K5A3ZDTISmMfSH3Ya05IckA
GF9KipfC6Z6MVmjNBGa/YD5dAnH7Z+P2nQX/lYMu2JmkhSum6lDPb3eWR/DfpyxI
eD0GNu2KqZdgljxKvHKEFpwPR8HObvAe/Mmv1P0KXXjQnBhbRtUzp3wtERL61oho
1sZJtypYjwP8q/fUfSFpjHX9REki5uIOFodXDlpkE0P5mMiRCTkMatN1BD3ndVQh
4+u9k/A1GjWSG/DtVIs1gl6iwhJZ8kaI/QTbzFf8jiSEtOozsiK2yoNH+bCxJIas
qoqcz95+SjbVFHsDQhiPvl4vJ/oIIX7kP3+VIIEN169Y+a12X7X9PEDtCsbRRnDR
4u0PJxraS46wYL8epkclkNBvIDct+mmXmxQzVNUmK/LmZdFqtsM2NHFLQZwd6Jma
`protect END_PROTECTED
