`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJZ0peUhcdYrthXMzmt+DoYTifBratKqOoA8t5EjZJls
k/eqxKEV/0edVRhes8AEC20TZaWIvzaBVevVFQO0LlDJjOovGpfyridqaShAldQn
N1MKj9YYU+eAX+411k0QQy4jTuB7R62OF+1ry9e9h2J5XUdUzTmkA4dIsXmbKSGR
joBb0sxBOrtByg7Qm24wP5BRZe/ju5mt2Dk1OMEbMJG5BDEnC7kWYHFsorXEQL0p
`protect END_PROTECTED
