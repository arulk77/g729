`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+dq9OIX7eGaVIiAywhKWafsMllNMLSI6bS+46/UCj2J
+d1ZisqXHCC2QJ7nkEewX7iEYXOikXVHNTfZMzSibAViO5XWEXfwxK0FTpHPQBGg
niRHP7CGxoJ7Pf0DeyMx0fO8ZvRRrkTa8nOVcMnGicOrce7StjaS6IXRXOj06MS7
zklwKsUrTZWp+IYpEnGs5s9nWabLSBiRuG3S2VSVWac=
`protect END_PROTECTED
