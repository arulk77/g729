`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ph8nMHTH3eHtJ5O3c+HaqsNgq97za8U7ym2X1I8gFEKmpPaN1kYLOJJZoa8FCkD1
+/stFT9GvGk04NdOh2VjrMnH+/4av4eAsCfxmOSJJHEOlMg8GsOTM+VJDLxlnbew
jXBMmzwGwmMcVtOLWYalHE4WvjqffPF5wiZBKOAoRMACHrqbNz4N93ufoqyBmyTX
IhRftaMIJnxQExXfKeP0vnFI4nEcIZDqYXNHb4XLxH3OK3KZtGgGWWtqqbRlWCZT
5osxSINbKULvQSHphLgu8TIuDhhJbId4vIhLorseibahH8v7HLj0k/yNHrNLL/bz
6+07rGjsqtUWyloRK/68hApMxspZzVqw1MnB9E0WS6X1h/ohQgD5pPxlIPP5VdjC
CnEe+a6uuiYnoFbyTnNaCReWPjGU1xBemLel6cX67gvOb2DuvYz/cfe65zabZpJu
OFCLML0hACZbqnP8BVvkGOt9dIZwme3qk4g8JbbTV7eCf1lmS3eyHuZrUXNMh7B8
wq+S7BeWu21M+PJaXfxdIuuDBasR1aBsrTQvi4X08ZSKpFc/4shhBLJKDmOdgI2p
Zs6YB7Z51UU5BVF7JTVfF6VNNB/6D+Z4m7PKcj1FBuDD1S9NdpYlpdbVK5UZO8B/
yPUkTplcfIu7CiYEbX3bnIHLM5gqTIMr46Mz8rGBJDoQmJb4ow7BC2lt12S/U7sx
pEJhBjaak5shTKGqCvbeaQgGQlMiNKPCSld8/Ly9I31XWfnQ9Eq3YPEBIRT63KGV
LoDqPNWJ2lDzmY4EXwtC8G243IMsSkV8L6D6MgRuch/0O6B1Z10Vn1/LYXYzk6mj
6tOIQtBpoyYCkGG9u+U2U8zw1fL3Q5Bs+JLByq471k8/RuXc0fd+xgfkHNz+YH2f
c0R0NG+H9rNKVHx9RkSoj3UGGQi0V5ge8Xz9cIg9sVZUQZms+SRDxcHXUQMRD8Bd
9sd8702Fe4zhoIqz4Om0REQ45qXa6HKyxOMpacTyt9q/ocIo1+S6tXjzIXkKBhET
DM9JXAfG3CDgVo7aI8E/AT3VmikhUqV7xaAn/OUq5/pzoMqbnY0S4DEVy27i5uVD
Ht1IURlKpHmxD0UHv2Lw0Zu21DzEWtU5WcVaUMpZVrDXfMyVfB+JN09QeyMqJ+Z9
cDmV1ZOwqJGMwReBElrMbNDpNuO2ywSGIBk+Jz82Bg56RjP82VEKI1i1TE53xHyg
QY32G57R9AvOJ/hUYcbHKM7t+K5k4mXEnsr/47Cdnyq6agRR5IJzm38ZLo6w96Hj
ejw3uvsoXDFsauqafKP5p9rc7rA9HxVs6olYeUlMNpeSQhQobJivu0mj3t/kV5Hy
YUKP6QvmIxx8iuEdtVvug/z7ZW5P6XmIkWizqaFx6sQonfqvBUdCY6macc1cx3YA
v7qPwjt8Iy6oU8t24Tlxr3RzBofrVahNTCRNMst8GH2+64o9cvgl10JlFzIAx/v8
q4nQfzf7rTzqG3Xq+MAeDMIYFqjkpFV5/rhFC1+1Lx1+TvcxovqXuAF6cx41CKyT
l9tP4uTP2ttnoEI2F3xvaApE0iuYdll00uXN/Upy8WjMY+oXJbBaxKM3cJKsvXjk
kdfsDKBhSbZ71Fi2pyCmVqGHfkIXVcvnadh5I33mzStpVuAHrvQOcIyAO7YKT95N
EM4nwRqgSfCruGS/1oFFkJwr68IPwIwJgMoBjEj2xubaGsn3Nk60rRPR3uqRYNWx
+iAio3rgpKrP6T45da8VDBSBukPof6C/CsfCHA78MZ8RMWVkETa5sYHq/JO23n7Y
b8rK371ip8LsEhBDUaOkmYSInYdb3ED2ai+V0itdOeGagZtKlo+dtiFjQ22dDZOQ
U9fuZ6vLwsQgdxP3uB4TYsUcesK8zgex9gXfneBSSlmRstAvZ7AV5MalWBAsKj16
CwdR0jAWFQmxCKTQAJUMU7GwTV7lFezn6T1S0/yQU1H/r29H17fkQd90zNBtiFqE
PQYy3aM6eEnzxdY3T01gylUcynwk6yz0dRWyJRVMkX8TNw7CelBVboFri51jIsVu
RKx2kT1Jmyt4H1dbZtwTHblZqkDvhEJCkqf+Q8ZEuurSIS1cRABZBjWrdl7kbb62
jLIisSMoGvOmwKWllOn7cxJm7IsDuzxxxocQ96WoSwDcRvdr2GGYMm4jQTAtQlcu
xkmWSEgvdsQxvz3bZJk1m08KUG0fRPt3Ab6ABjY8X1IHvJWOCjqEkqBx/FgoGX4p
hPfkaNPFw43vLsOfomDEP9eA10EoqlWyyr7i0O8QFEqvEUXoybCu6AZ3MbidlR4z
+Gr+CUrxnX3QuAUt4Kk9yJk2PfXMKo7DguPtBi7QIlIOH4uqGtUiszErUF/g0VSI
U2+t4vLWslO75gYigh2timKQg0Ej3EVw3qM6DH8qJ/8MB1nuv4YyrHoKmFe4oiMz
3qMGnpvr9MwTgMqNrJ+3Yd8hS/OdaX58dJFUs8u+cUGF1aCGtFua4CmT+8KKICR1
mvtIFDMKzfBiOWYcKzv/hun7wvOZoPzrem/0bR9hOd25xbvBGg9xNr5ZbLZsiycq
ezpsQ0ygubEUhhTdXZg9SzZhhYJLU5uAk5RvmuENZVCSDbaAWDtxhb3Mah9KylP8
Pc3tKTrbRHQ0MoN/92qBUeplKqdSEPpxJPPeGCKz0To52CRq3MwsZ13NjjGsZiPa
j1upKRitzpoV9OKp3ZOWpDlwU6YCtrob1QROSVrlRzpLteuY90AhLwuCYT2XxYVn
3+wOOpEeU+D9lhqUtBgN2wr6wQUhmLqwJIoYVvdKuvJoF/ZosMKzo2PZUrvOJuc4
tLAoi2qRFL41XHvZwOgshioPDeTx9H/u4SCWSlXDyDgrgDAPLWWg/aTYLeYkOlPC
pfGeIDSwPK9RkuEkO97Wu6CZa56dox83zI4LrPgC3WfA1n/Hrxk763ipfPL1oXed
YYVKHp6edcXhGQKbpnFS1J8TAxeo/CLE3/uC21b0zMTtJG+LXhBeEw6ubdmB3KVW
ycnpICzFY2oJx7OY8xu9Ne6qUT54/+GzX7ZwGj1BAPwhFjGulGEgy4r8i8U+lFmq
OmCdSJLRfWSvi8xQ0N54vMC0CdMfnwLwP1YdFZMb3czhJYMeItKGQcQ3zOl+1jBi
m53kF1WP/4o0z6jCanlPkNIbylaKrNPjkzy7P4vWeZsgJIF0v7u357L+bvH4QZW3
UICoQYmjXyblefE9S5mtNFZtgx6nB07qkjaQvEpy7MhYkv3KTzJDGNUQFOAUjKkn
bMLCpmsiGsPjKk/JWdfuaPEK8DDjACCtynXjb1rhMSD5sQpJJLNHOymllnESnUBa
z0vKnMivA38BZKtN1Is3czjLd1zb/ODRPzx5TYKib9aHFa900tVQ7YvUmo4of95z
NhYGZcVlDtEio9LAuG5MvnrL45y8xvomsexv7cxD/xmdxoPpE3789v0L8Iz3c4YF
U20rh7kJyT0DJtWEXDUmygETmh6tAugg4rksFyp+hbmw0foAmL0/kx5UkFrmjEB/
1GObbCE/lCugO4T3Uq5VkDpVxXZh8OrMvKHqZOGEjmyYdhKwt4sRU+Pb79zIN9k9
zAWPuDHe+NxEY42CJMK/aOuvaI2Oz5N7RXU44rwbXBcFB6vyg+FqQCjAG+o7oGw6
LzIfm5nAPGXag4zWltkF5WceWNo+Uzr45Yq5Cu9rX3774eN7oHTW2471U95RYncB
elO8nckxr6UWCtlUe7NAerTISwMcG/XDGnD0b7tFQ/R/uKxVnCN1fxxDXU8/F40w
PQRH806ZJNyDs3tzknFUtLZ1zrrXJBkeb2VIRXsL5domK+3mVXKUx0Fm+5L0mLur
9rY4Jz6QZUuzJN87rHJ8gt+/Xjf0WF8UOnKaVTUSvOJRlrOBBQhsWudmIWmbFKTg
Nf6UtcjFa8kKDCEZD0W0Vg6sDEznSTP05jT9lzrTDMnxVAnnhuMYZQzXJMHf2l3g
Eri70ygsn68iAd7P4zZaQ1XLxOh0eZkAsURB0W3Vd4RPfMUK0buDUd7dW30EjTuF
xG5uJNOw0i0WILufLnBZq28OC2DGcHs7YosmoiFj++PhGagj2naKsE/B38OHjEWF
9XvYLvf1AFVFBYbVkkmcooIGYQrboQ6Y1vnOdBGnHFgPJLw3oZE37Knujt6TDo28
xffcrp9H/jmj3uJ/uUe7igcxLFVUCnt8CDNSCpZbGfEn3v+g00Q1eS7avRWUeAqg
a4iU62bVcwb0vZ2gi6XQ59T6aQsjSbP2eTghb//WeXTsdGRPvVVqGTzBa3YCUtBK
Si6psnICjnjffU+02sxHRCw+Xb/4MFP4SbW9FOgcWTLckx18rwYSGC0R/edNrakk
9umTf12jGpxjHeV+ogumDzZOzakzonhMmfNq9U1Ts/u7KZepjhNPEWVPXIwWGJcP
D7urasY01gHZy/jWkFfAECyM3r0SUlGxDSfUDq48f0I/pDOWv6SLCRUN0xOwi42z
oCXzw2w2KBE+MsYkTI6ABXNRmI0TZ/JFQQC1WcKQcktcE6F6NNeFRPWUp+F41MYT
nVIT4pI/U9GEeZeb8XT67LpfwFw6GmcLzxEAWwPiQlcuN4hxyxNcHTO619T4ZXK8
/ni5LQz4wXW/4ghOq+PFls4T2JrV6asVtWvGiSnXvOJ9iU29JI15HcWGzKk3AXbU
pjuZzPRrXSnP+LGPPb/N60Sub42Q8fTbApQiL40Y0zXkogkpvSrSdK7Ww1KLd/e6
JAC0iY/DM4AXiPUG/cZdm4bVI1CV7g9+s2J2OWYti/IC19fiVq9LBJVnkHIWCPar
v6P87aM7LyOUnDsLPKIDJ5CgnubUkc79WQwaeFdVdlC022g0pwdIeaRg0/rzjYw0
pCA2rv1EtM71WO/AD1jgYcrutyv/0b9iZBRIMsw42bI4Hietk0NAuVIsjpveMfXL
K/6UJl0Zi6wJwdlxGENgzPUlLjgScIeiWZ+XxmkEb6SmVRssHtjzsP/+0fdbmVxw
UmIKUITNOZbwzYxjH+ofKnQA96CwC2Okgh0XONfX0wNMfd37r2WBo6wkHbhgs8wm
yufxw7/Mi9QcVdUoOv/V3EyETyxye7uw8nRggNaN20yr9bx4bRaKgNvQyzt/xaPj
+nHcW2y+79tm7HYMJ00A9eV6gseNKfaaiJ5JUHmqeAacHUTVHGpoOqqxQIaut5X/
LIx/LArRGWff7VmSKET70oWVEVqz4wPLZTgmQU7faaDhBc2gkZtUxHiVjMI1mvFB
m1mGETBtGGtMCA97T9lXr3sbNrcpslRFtgZ5OkDN+bfC4lPIheSy9ZCS1JcDhlCp
ccLLbYuHv9/eTwVTz+O2hoa7rPXNQ/6HhvpfylQ2lhijqpdQrSI2jp5NCA1thRTX
JG2uPmOjHk3pQFrmbq+4VdeQkoflPWvhwcIJyr7jwpIoVsTpLWZQC/fkoAQXll8g
uNh6i/ard6f7jbZB5eCVpYbmVho36nGLQlta2UpiPoGr57G73SPdXabenyuNJH3M
nzBuuSxvi5R2rfQgQlcEo2Lv2qLOuo4jvt8Cys1NjRocON1XxymrUdGMrZPKVUnM
C5nAKYTrxJrHev4ls6N+gGbbwTURuZAXMoFFLxZfuPmkL6FW2J1SlwwE8Yl4R4+b
fYHsbAMu3BvnIR/tb/XryAo1gBCHnnNNCUN3nsJSb1PmAWe9xTSn28DxJ1xvcryw
K307fjOmfNnu39ARkt3gkeBJFeSAEYMH41pQ/LpkoxoeUFsMliGTTUDiYFWbHBht
eTbc2Nhg6FS1nRB+HvgHAcNPjRCmhHU5xZCbuVuZoOFfJdzigX3ddrcZLI8wKweC
/6p4qQfys46/rJIUDtLU+k9zYBSq2VT6/6TiZ8GZtfmLVCJZAwcSk2QwfUva3Sd2
SEO9gGnPUSeFOZLt/rR9eUlRWfg78PKbpAmno1ar0yGEVrRfMxPu48G6KUdMtoj9
VBEAJXeRuN9yUPivie9ZRLyTe+ioJ4rt2Pk1t1MCBx35CJ+mmgcsg1GQ3d2Fyhyq
bvjSUxXhWwibNnX1YVuUHu14dEjdAEvh0x7lBrK7zCLaYqXN0gAB8cGe7ley16hb
+Tzs7EOCKuOhugS74RTO+zUmLfU+SkezH1BuTO+5DFvg/lx+1/MShUbJm2MTpRQE
hPmTVHxY2kWAGMh0ocBfjeaUCiYZHakQ7cnCIiZkOK9rF4QwHAxtkrTqMkeCoQDi
0OGoTvRqzFxX60Qlt5xCpikPTfJkrv7jZ/niUvwGB5pgAF9JZvAgUSVWO3U7Kyvr
mkk2M1R43vB1PsPoGKaG554X8iZz+I1YruIV+aUyEFVgpEdQdI8viUlt0vKhqYNO
aq01mIaaDdArYtanEyDNXsqzPdxrPKBirVN6L7Zd8Cq/YxNAovkLs3MJjvFGvntE
JDOcsIUkAso4xBirgUw8HYp4g3PfUG0v/PAXUlMcihot+D2a2QthBVvcgn/Kgy82
X2mfuCDBRO2r9tpRXZHdLr4inybsDKezuano2FPaTgnPnA8/lCD9JcHiIad7zhMF
trxvYsbIHXbp8aBd0rylwlZsdqMCIsKMxBfil362XKLaEyppbAEh+ThCqPUGsZ2r
ZxQov9twTe/bwwWaWVVuX80bjY3iPGsSQIlT5bJ/c4T6qmhOaU95B5lzRJ8CNcSu
DriuMaiJfN6snYGii/mb5TF52jbTGUgW1lYHsAljDz4a+EQYK3JXu+kV/eZrRUCc
QNFqGnD/wQAYqsNrK6E9EbwNx6ZEUU6/HgBGNSvytuyIQyU4gK74AgMmcXBXNs+J
uTTGNjOud/xSK8HBwP4Nbs560VOAKfTE55nsRXB+GOx9aJ5jUdmSHUPUqWhM0WZZ
Ltc43r7wsZYL1BJBiO0Ihv+rmxnj1qXsrdg49cgJIKNj4Zgz4D4n4na9Csi/FbQw
JkivP3f12dsCuVoWuTcjyBq2GZAhzlMpQ15hQZKF9vPBM0N/1Foa5OmtZf9Yg4ws
66s2UtQw/k/CSSHqhbrwNml/MpskWyr9d11fm76dITIF+tXpIF21oPMijOAt5y4Y
vwbNfXVU8aRGowle1tzxgKyZufH0jpkU7Zj8fd6MV9ZtiAoAwPWaNdZASf7BBHsg
jl8+kn1MM2E59t7q0tJih2EnZ2R350yBk9ivmOzLRcjQ2IaY//zfxOedn9tyDvi3
SUfSD1+9A74XGOksJcNuI3mlQLjqMUuw94+qGJCB3gUi9qKv5hpe0X8KfxIZTdBh
7Ilwl38eucK9/PVOl/j7aIizBfMXsoKz95QqYwZXGAPhOmpMswO2yO975FMNUVj5
+GnXpYuOfedKOO05ZJzAezXm1+OVBRroBiX0ldu2Fxk6zDNHR4IqSho44AtpWzLG
dtrcyHdnqnZ3Wov70niT6xkPWBjtuIHaJCnTfwesqpzRVH+Pl3g2qGc+BJrUNaBW
naiSlCGk68AqCZSxl29SvIGHp4GQbxey8z6mg9KGwYOhZ0blo6vVVBStESF5DocO
Ccvb69U+KbuUIi4eCJBVvJv05tuyOYLlhROUS2E1AT49S5WF6TzKf7asfgeUZMlV
4zD2E5kRxOFREfb3NXmdhHqUFEwwigEHen2nf50iYyEMM/Yz1Z3GKwQwhLHWQgcs
K4HT9XLTnZRdaXDXflDbYlxIAi0kDW+h6nyTdNJVzLtRBQqSoc6uVB1typRPx8/M
dv37b6hAgBf5EUrvBoKSoZblLXlvmUmiEY7dmLWdsgMoF4+UUjGF54yPpmA2a2dW
MbKQ7ccz7Bx2Jfj0/fzxZO/jCPR7oF9e0oyV0SgttwKoLh6iNbFjK3d+1wJN2Y9l
3jdw4mfNAj+KIC4xbOEDYtTsk8CdFd0PCd1uTgMbOnbfFQyqhXz8nrLYeukFSA+h
ZIz3EadhL4kkskqOdQJRvx3SyRH4AzsJTUh6E2eM8i645i0e22eJd8anFGCPEcLg
dFFE3lol7Ymfz89n+nqMG7i48c/IYE1XumDaV6rlU4lHrhhw079Ox5978hliVS/0
SJpJmNyXnihjTQ26LvP7N2yA2ooM+0fZNhH+yrZ9u9D81I2ze9MdlDCnov/Spf5M
pa4uMmsxd4cko4hDoGRJmjyuKqpjT/Vx+3s1Dh3QcXiqqf+1+dQXVOp8P10vUi8G
diDUn1oYxl1ATE2sMwwEsDvHcWvLHg+k57mnPNcwYTH/PKg1uvi5oSB9HCmXGLGZ
iy+WszAiVmbzbkI5GD9/c+xS+SLqyvYLo4o166xP4MjE80DO8vhtxb4YOWhO5yKt
u+Nx/2zbxCICfXAhBlWKZ9LE+dNlJ+uBzUJHgoHXOr2upatHEzHpKDcL6PSKXUJ6
/GgqLxrUXV+P+QhSVQRx3m6TKWYCXVaNcqN58TBhe9zgzI9TqlYoYS8xfissYTDA
NTWn9XWxMUVpG3QdEeGGFMO0X0gdRDDGgWs6OKsGsXOlNLpwjTLoxGDvAU07GpVU
NQh9CXwzfg/S1NiY4iocyITbsTP0z0tG5733qL7g5lHNheBdf1/WccenzbfigOcs
y5B0d/HEbLJAkMxaAhcoFffgRKR0VD5rwcvMghl/Y962nv1zuS9+z6XDL7A3XCR1
E9bC8Zq473L/+trYptzqDhbMtp5ovHLsa+3ykxTfiS/N/sV8cb+3QRQjGJq9AnWp
fONiVvF/0KCV1U5u/vDFCyTseywdYXBALRbIx1EkpVhyD9gAquhCfYBftzjvFe+x
6O167wIMdV4RioGHEvltqnAuPSKdAmE+DqO33D5P4hx210d4rPeWeoTlCTNXm7OU
JkmkK3J/0/KTu04UtNfeF7ifqDww3On6lRww9DtB9hu+CB7PeUa1LQwPz5WHSgu0
a8RJYacvUMKr47XRGb07YpFiVDQ6NkmoD9r/pJula3iOG7Rh1JSoCQFFfxCZYhq7
0taAo3rVy4wp9g7PRx6fGJPhjTQmb2Ex6tJvG1Pxf+RRtrIQ/ZN+uknVG+kZ2ViE
n7iOEkLVzPpQPtj/Qu8v3CnpPPm3r63K2l0tsZF9Kj8NGVWe+v73muS+g0828rV1
Pc86R3Yd7nZ0HfjvaOTk/yiActW78NSuV3P+phnjKvWn0JaXPHnL6ACyum5+9fKI
pWJtBXUvViEsisPKy5mtjShCaMtAUsgQfdETghZMnfawPT5efmb8giYYJ2BNGU6r
uCNIcx632mloYBoO3rotqNUMC/H9tWN7lVc8uqdXOFYux9eXwWET1S1yMlvnmB8S
ZmCqgRlb1Tl5DJJjRygvOPHBufySiqkiv+z24OXvQ9a8Dl41lOfk7YU71LUh2uRx
C8Jinm5BF0IXbrYWT3HhAqX+ZoX9eR1jG6r5y1eJIXIXJ3rQ1egD4+xhkWWde24L
eMc7Wy02YksxFXyaA0chAA5gM6Y2g+qztzDpMoUFmjtx0SzXJrtYyX55REKmeUBn
75hO4vwzvc5aXDvzW3HxBHonJ3xeEGh765Ygm/ugF4en+sQvS1G196AATEYbOF+d
u9kkYc4Mh7XjwyCfWzkZaXwHSMNbKox/dq2ZPYD/cixFF2hgOL11r2NjOxPyjCQC
Q55rv3yp39O0Ayu2QiC5EaG/1txMmK8TGu8HfA0Gz7T7aAeYLg3b/d+hsScBBS/3
kdWJf/NV2yt8Og0cyyLxe57nyJ7ye+WZu+HFd0YMnJqOOVWjxueHRQ4C8vWbfZnV
KZTTe5hJKWDHk2vGEvQn+O6kAzzp27GZdY0aUrhYgXhta9NSxu3o+p2tzcbOh3/E
AWmTsYdtp3udFf8bFCK10ZlqD/Zip8ekpN9LsfiZON8mwbqskcv0TfFVNQmA2w6d
9+7n38hYZ96suwozsydk+Zm807DIqsOcxsDRW0eGMeyb/fH0rTgsLMvitCYrYyfd
GsLtaiLGdHwHieVA8BV+HpLfAykJCLfYTWYY+4OQ1mbuAv6onT8fZXha5jdY/Lkt
3sroI0YIFurH6XV2DUu7HaTAFF3nkiexzR3oNVS5NA9yyHLBkj20/JcCeT+GHuql
cMWvxz78zNIGDB9aACIgkIGGZR9Vajm17kTkif63i2yFl1CaULCp6N5lC/hFaI04
J3q8u17d+fjD54xz6dcWqWQy3yaDRzqxl9BVrzByUlCSC7C8kSvrzk11+TTlOL7G
lKayz8iP/NnpOHlu4n3Q887PHl+CjAzYj0L7Bg0HUlZrEzcWOLJGU2rnWa7qqzl9
36N+XzV5LOYJ16XZPngGA3zQxqhxKL0mWYn5qvsZO33jCgXgVjkBBoushEmd0Y5D
Rrr8Jv4Cm1Ves0ILuI3gs1XGOMtL2KQxBncVl6qUzTfXb4pBNJp9oOU7dF+rUaTB
0j9XDDOLibzXeWMo48k69VglnPpewtwCUaJT5IlzPdig7Wzx+ZW0TcOGzVB/Hfoc
k7RRZsUkAVfbcLmA60acuLhEbIGq+DoYw5WEDupVFEH3b/ipcGBCPfXNe+E8McUY
NX2m0u7VMaO32LdD+iAGZEchZm0WEAKIjKXTw+FLUhIywLPlVJXFLNbLAttOei9E
ZDve1AnQTS8AKN1z6DuLHUL4ksxrKVAvvt6DPG0BaOMJODOva38/ySDxJ9/MVgo7
rbW0XXTH2SVPrR5EqpHmffqi+/kocooGvm76vpH8LXdpuhE9LTeO0OrTI9h315TU
+18QaJgi403qbuFZrtqgT+7TF5OnPzgEu+cNTC3aQpX9mvwP+IdSykKwttN9/1a2
AEdfPI9euWLpgCcJKCc8/eO0MKh6cAYY6Pf6KJg9GTdm/a2WJlyfUB/gR0f8xy6y
PjjUsl6mGADiSQxpCrjb0dpk5JWtPqIR69lJxx00ZzjICygYizgt9KAjOHqhHVn4
jxDpxYz6zrPD+4o+UNNUJd9CbGiE+bCpkmiEuMbH/RNvtjC16mKacqMmwciNg/BB
u8p+PxcyJbmQtJtdV7Mr8lYEh+MqgzwI4Vupna/Xp39KMFWXKTQori2Jt/piWyQD
FotZjtZ41GQqihod4OvQiuTcZ/04zIQxld77zR8pX+a7HO7olABTk3T9TklghFAX
dwd7K34Y36c+b9LbDqATIqjLarQnj0/rpIssuO/8mZaH6OQYSilxMOrzUkMHWqH3
8gaPaIWXFaNYNLnqVaUcE53ljljcofFlfPOVzuCFsLOa2feWnxxHtxEaFUwkF+m7
PdahKn2Urc7vL4aN8RxUKcm3hSs+sf7Zi6E13xh31hhzFtTcKCbHBNGqurVGZU57
jfOxEoW4c34YcBcKBXuA4VSnHawYUe+Fud11h0mYtsw9EEDUh4mP3oQFAXpYSEZE
0NGjaph4LML3cMHr6cv+LlccRZ171pkaN3sYxy57+jWtmK1fyix4AC82nlEOZSJN
DNAN+CBKruyzYYILpSYRDK9z8Ek5pKtjyefBa406l2rq5GKO7XX6+4FiC8QpFXr9
7B8CeRFqODPEaFq9SZTRMVuzZXCxHHEzAgL8AkteZIRpc6kMKCODJh93zHUVl3yz
jj/hBB86Kd67w6Y08KoD2xu1ZHzNbGhcPhnLYECkWOLE/RKzOuwKcdMxbZFfYbGs
oSSjBNR6XPK/vJ06KF3lcM1Z5mh9rkECGnOkQattvH3D1Wm2rsQfqQ2gi1JEPzFb
eCBPpYJO7MPSRwDoNKyuQ36vNC5wcV3bs3wAG08RtIiPewcFSDDWvmjYRH5JwAg2
vj9NDC7ZztK8szLOubGaroKD6w4yvzFQACEiLUxg39HxR4+piQ7qE6zXcuQtthbE
afDvO9TdrknGBGavWQAFcW0QiX7t9KCz3ZBPr/EMLeXBwAW/qjh8PNtULMfJNfSV
f3XZEpZKAXOxrRfr6zBntTEG6uSqD0O+yi5T52GWAN/EQVMZY7IgVmFnvqDOefFl
WqCeGeh8UGuQgloPDfp/KwLjoy/bksCIxJCHTOJWaH5ZKej1Dy0+j7hz919U82E2
pQbbnvLhrQmxkXNqyxTMouYmizkcVlTgY5poNYuNhkskQfjKd+q91XVRg9TjGE65
bZgLwuJKhPEoqBMWM1ayfViHHIIqkW3hzOqlRVgFLTR9torrC4yp7cmbhEQIrFyj
qBREaDYp1TkDc7+7nx3YrWHS8VLaOpxF3h6OexZ0QpnYZC7Lvoew0y9VqWZRHssf
AsySASq9N20RcJs4j4YNGEZqRzHdMxwZjaJNf5TVECQJT43XE9ZytJ7c5teTKxeJ
+ccqnbdmY7/o1F1ankQfR+WKmUxmQ6npEa3tUujW2IoDe/3XRscm6LNey5n2Dvwr
vTJS0EEmjWHDfcp79kCYdkgRjKL26h302jzE4xOFUtS1XOru8RA+RfvuXknA8Dwb
PA0mGq4jUjcz7K3MBZzjQQBnD4/lISfDVOyncPhvO1RUSOWUo+Mh7rzH3duTTLLc
EY3DK6kcMfLNXIB1i/5NqRq+8xCrw4Zd8brBRmR69wH9yK7V4hJb0661YhvDXWdg
MNJjpM4zog3WEOplqakvpHTxe7iSrTrccSCXdQVZ5/UgQtMKltSjB7G8EjcyVTsp
Ywd+6yt8f6OPBx0PI5bL2dWb1jxeFv8uT++eXrFPwv94mUdgRZBX2OKDroM5pZO1
rH6pU3xN//1Ms/2BvoVrG4fG0+vG6dQfNva0OnmA4C+jX4q3+s6I5mm6xSQ5NyWv
ICXohLOx4vIWR7pWHGqF0azwZ2IVjmsTJVAKxyRng4a1h1yvZ7PrKzN12HMlnBQB
+dFPWaEmkKruydVnPDSvzOEc4vyR3wNboS7APNw/hwGcwuFe5/wEvuUBFz4U1meS
B6pB4GLT+TxJy5f8luiB6+9b8B1KhhHJGAY4Z2x3xr8FFRwbmG9jMxDN7vQ29GCn
Ba3AVyynPC/tWr7QbF6fyqtmgtcadItuvVZzmZr/8gaFGYMAFWXRK0YTCLD1a9Bi
waCBcW3zUPUjWPo7RqApwv4BTWb9oTz3AHglsrXXarkHGxf56OvGy2dO3DrqlS8b
f4X8fpbjQNdU9U8+W5aRdZ893fmZJIanB7f8hpL7zxOH7SMc1yJaPy8nYDw/S+Xr
lxjA5sEaq4tLdpkVjPF1WMgDWEWl5+Y+A5UR61/WpWOhJ9ug+bcoBLesCfyseosj
UJIv3t6ze+UKoMJ3kTSnmbZT7gpwb+ZDAXPG39GQ9e0wYAkhhhtgUDIA8xjmbsgh
o28BpNqzZ9XgUKkn5VMJ9En4MYnC/TW6Tb0O8PSUAuesMAiu+1sFvtbFj0A76Cpt
a6ur8LpDiZ6vEBVypuTj+orjU/dfGbcWs5IpF0DGMz+8ibj+jfcLhU4tFgr4veic
5m0vynSUczTSxbI5bS0nP6qZO0iS5/qR83zrM5yA4H4M2wxvlJ+z4GMJb09KwkEF
eNLRBnSQuPU3CZoPEuIyf4bPaPMHvJWNbP8OO/Rgd09MdtogdCefibpvNt8wmypF
tFcK46dsFj7OVu1xqS6/p95YF/M/7f26qSW93EYW2M5fL8Xe7IzHJhVX2kl08nou
ucYfzAdq+L8VWxxCqEiyJEzHLlrXwxy/0PPccUa9KL3tu0d0QNPFsnGYFKiFa2fk
7ZfUrdmnr6d0nZQitk0fw9U96rINTvkhkGjbZ9uzGTYGmlmPi52mA5Z5wD5nUpTJ
3WvYnGva5e+JLQWJjyoGg3uEUf++QRj8goQAPbLUy29m7OTxH+Gsu7a+yX/WWEYS
cEb4VZmqQDnNcizvoBLSxqwrJEianGofJZTudnUbrOJjj3BRT6buJNdSI9B301PA
I5FTPrT7SWiOY8/GlNsnI1TmLzCDCc3AbOw3F+uyi2PLcqkJvmLivWA9bV3K2+5X
LkdEmPI67v5beT6Ll1BXnyHO5vGiHVHdIu9l+48QULJi4YyvL4qUBXXbWsAsbAtF
ykE/9Hdvky2sPxuvptFDgIvxi85OKKNAH4EKkYkTy7R6AdSoMIU5NNApypoG8thT
nRCCbROBLAv5BzEweHvneyRFPCgAdiLi2qq+VnpBPICG6Y5XQIHqcq0cXN9cWgTn
cs+6sTGfBnbVWJuvTmFi9fNKTa9siSXTuwNm5PZKAmOebdhHqDFzKtnc6/eEGyEi
g/i+EdEzqFRkf/lmWlUs1rqdnz7e/LUqxcciPdp/MvjY6RJERkH3dBFqbx+S35oh
QQlRQhEH4RO4TaeyWwdRXfSGPPFbem1EsUkHb80f/mRHxDVi3Ddo0K0Fl6BkZyox
Ko3D2MeyzJJ+gobIEhLRfOtVTI6ht9VFZ3jk9a+VaikzT+q/6BzS4AxtPPH9yme/
FHgmarL7UMb73MaRWTrHj5CAVMmf16mPSub7TtRGyBcYHCWc58neLev83jLzaprC
218ZIKWm85hNucAXBlVBEx4ozw9Ut+djcD6AH2+kjxQdE3lknDC/8P1o/DLXdglU
onpKsc8aTcSacmdOZCKDugQT0ZVPeLdoy/kpgWS+svnYtTq3cCNWUkIXFD4oykhh
JcjC/Gs4kASHDICU4PTyYxAYszHAEaXFCFcEPoL/S7S08BT4kl3maQq+/dmIplLa
BPppvqteX+rIjsX+AD+EbuZyMFu9kNF5hFMujDVL7jSifiP1IKi3zXqPDxiy3Df3
PrNu4eyGD22x1BpvaMHQDEqqkjte97nnn2uoWyXqRpHfwxEakE/sgQFhcuEMnK/z
Z3F2mKwbief82WiOz7BcekUD3+N4JpTW5UUH3jDONIcKU01a4RKIfx/PYtXOvT8y
63842io8MkTQkmnYgTYgOyd3QzCHNyvvOCyJK9WXATKN408cTRKPDhU/GsTrnFmc
bNL9IOklDR6oawK7+wj8HBnn7oLb6fNs4/ndXVmk2icrT0oqKe8CHIBOm7XxwAie
s/vPi4I0vmcqa2mJjkmWgsLTnlZlnIuFhNYBmcC8Us1PkPDf7pjtlp5MzcdQW3H9
0CWE80iejKm65Lkcifi6O2gqhbu2soK0aet+3rf/8dizmDvLeVcgeQmWq1QUpQeq
xlWupXHuRyldGLkS5gp0hbG9q9CUEEr7e0FU+zhGIxgt0FQRYrlK1PC0WcMH2x2V
qXOAmkkwi09ps7R83OkZMnfsLSaTiySqJCsmrKHPQXeqt2FxFIizrS8L40CfSZx6
KTBOwHTBpa2BLCL5V+VEab1k29T0Qr0K5v+yKQo8sZHXDEUOQK7fG/rtu9/8dxDL
XuZXfUCODDOeTSqFSdS+9kMoRrbhA3h+IIARvJoaBfIkk1+5ZzoXQvt/YHku3HhK
9TJnaV4nbIZQ0l03RZqjOuBlo7meehnlcquwtza5MMDRaAM9j0kZrvFBaEdzKZ19
x8Wje0b0IpshoeYl+pynNFZUJbNLQSvhBpTxwpg1sbfP6eBr/ERfyDE5H3r6nIwX
dq9oOpyCRmZY4shotGaA8cfV0WVk7XRUo0ca37+TsgWZsLKP5IO3qyQbz5j/2SsT
bd02kiWrmRRNQebD3l9MkYJalSANeQ0Nf/2NS05ImxhFOlXJUbL1s0XhR38xfsVw
MCLZuFgp66t/Be1JppYVgaN1gFtLUtT6rUDwWHLmSTo3ohiRMLI9cw8oFHwc+IMR
Lh4KU2ec1MF901i6hDOKIOhqfxcjxJfOdWgwcQluU1mDAkIMcV0Rr8tZRYKaYnXo
tbSQbIIpDapyIVZWEe9O2H4iXiJcTYhRsbOFOBJ6KZmOJ4Hypjj6Hb7R3vP1VED7
XwrsdnZI4LuYnd1aYO5gAas1U3M5lg5t/Nce6ROTy4b22Elis2Umq+nBGNF94ZO9
OorFb7GQiDzq7MyLwc/XP1rFBLqy7WwFUuuokxK0qTk9GEfk0X239RvBuay0wWTw
1js+Kfn0f56/zepPz/937wfg61aCERq8s8DYrOt4NQ0iIo5Q2qah6CwkL28vq9Lc
UQKRsvQ9klFMlWRXnHynVptykSmDOJn+U2M31BvOWg3zprMN7wkHUGuPpKzUyx8I
`protect END_PROTECTED
