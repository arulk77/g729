`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2un54ZIhnxaxw+N5ol9ELdBhKa9faXDHcM23LtdygsryFULW/B1yV+2KsEsU/dbu
EvfIBz0pyCUJhLLXGE/URH5mfPYjlGibFVr+os13nlsEZv+xfPOwwR+aFxKKkqyU
kV02Bqb91g4E89M5+6l+X0+WbzUEQtMbVUANWwXamLYz07CM1Vz1zVzgUQGD8y3i
5G12Jpz5qpifaEJAb3d3BxXCkCO+xpeamrgiYLY12D0/VIaR1hVEelhxqlO3D6po
boLjwNtUVFfyfuMJPJFOQAR41FybwO7kYW0iFwNXfz7X8CfSgJACvob8/yWAvOjR
3atDdEizqHCoqezD+eaZiGvYtPcAd8ulX/vn80iftHpVQFKHhxMwXix4gSz65fFE
aXuceQfl/VKuiHndpaWkOjj6HparNxzv3kkxqHn6YAsplHW/ecCl0dLFjDGsUVfN
AD4VEl1/SXpJvKgxg2nnOuKw4onGJ0Z/ZojE4KF2iOw=
`protect END_PROTECTED
