`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN3If/fsWsePBKBonCRgizhVyKWvnFr+uRADMadK2pllD
3/4YY1+ZYwzekN8IaW5tFF2DKof/QABSDAmPjMWm+H5m9rSyjZRLzjjXZvwZ9tLw
1UBrA6Sq/LOSvKmBGWYoLHEhlaiXV8EJtZNNA/ZelYqBiqtnVBplEluxIsHQHgna
kJY+zyPOVH89KSn0DvXhNgouo5si+NVE7MNA2OIbmXOPbLDkCNTFQzpeiMZbhjQe
nkdp38jksG3yi41wbOSZ5Aoj/qs0zesASm0A9cbE4vTvWGkrwuFIUMrr5Yddbb86
Otzpb4mMQ6abr9eCDxxk5pBlKaB5D62UAEvTic7eDkz/kDsdyGbTcky4YQFYQHrD
7Xnd0aKhM9zAqgZjn5czbhzNKJDKnh7RtUXoGybJQasyVP8TQ9eZjiTj3mYwRgTI
Q7SlG1OYQt6OIOQQU7WSzNmhpjquPFjcTaBm5/6+XGRL9hIVkSCxPyQgIsZUK434
EV5lLPMQbv0Uw5Dvz3oUupMxqja3pCWmIePtEWch21KRtJ+1UfeG4YXw1Bxbmxyk
cJtPLQ9xmSQu6CAB5+BGLPkgUsk65ENoAlVF0muyZx+ZDErFo6IhmslAZducRXF1
daD5Mszli5HIQjBki/xPFbtIWrvF/Z3QV645Tp1QKTwL0fq2Bap6C6IeCydF9ipT
EFnQGXnwgGhfog3y31K7W054E20bDSTfQJCMKPvFAprptq1Sy+1iTM9zDFVaNBqL
npj+08YQ2TD0p8H020GgbmUftT2d4tNbjGNw1KeuVAufUmZLtq4kHQoH6+bVYpBA
nv1fk6y49uAB+9iSzj/8dKzABVTXRL9R6K+kbLn/AsOzo77oKPXuel+gOqDIH5Kx
6PLZdFyogqNMXuPjXYdeIkYfWb9JSGn92jTydJp8GQFxVvtzANVjXvjFa5c3mWm9
FF+hFeJGXhi176T1WAXp3W6QYWlw4wt0NPMGs1rFTOEvtfr2GwvfypwzWeIBsMSY
ABWJuAJVC9EIfXI3Uo3O3JhtulTym/3/4nh/Ibk40RsqDtXni1BRUD7Zwz/vF1TB
2AeiI0mjETc9yOIP3UUf/4JFSw8ZGLpt/rhc62KRYqgloNutYC2EK6/DUdIvvW6r
dcdXaXgXlG5Y9lKzfQmCF89lOpyRu67h+Q+6sBTPwadnw4eiJtSZ1AokqjgTyefZ
fM+1g6LPzGSDZegEnf29LEn0lXWGvj7bZZEiLzA7+PmKY1ypDoCS+DbZFiezb2kP
qC+ohi3C5iepVWwjOdxy31S78CmKM6Q3+6WHaOTePL5OlfV195TwBdhRRAeQEjmG
7kToVpLmGgvoc2G5fMeLmexBryPLX3Zj+Pd6UgRvtiZxvP/ZBgFacSIefntP4ZQF
SWs3k9Y4q4WvIUkf/blV+l8njllYaWn9xaJ1Z+J3M+ru2Dek9Tl5uf/YiMm2qvlE
+l+PQnVhWY1YAP3U96C8VlxZwx2yO5X0rnb2OyunUvm6UGV0Zbr/pCwL4QJVW04f
Cb2FrHQJKNgho4KRC27fN6FAPXkto0M0/mdK5HdzxksfHoqjOZT607r2ZsREC7az
Wz70DXP3PAZQZbDSRuIPEAZafeYmz6GfL/bLEsfng1zghEzKXGjCeWgCpm/6tEUj
9JlEAn0+rnZZUHs57h6LGy6LJ0Kji7qhLXdA6CcdPPj63sqmSY80IijBbt9R03Ba
zLxhoGoVX/PzScSSn9nyAjgMNQXm7dF7WlASXsHQjPKRGGypUpMFc0DvRY04/89D
ikmzsvbyCA52q90f16d7qtuPHLmZr2/KUaSlnkzHc8wFNoNYgsOCJGhMk6GwvTeZ
h62m5TMqpE2n4bdaVA27ei48SV/WeFZmt/pqynWgzQ7S6gZpYerEvkeKWRVsuwv/
nhkgcxOPwz1QSWf89ulvxoioaR/l76d8LD3MRRdEPyvS4tPCrjf+nOyM87QIgnQE
qNrX7RLtKrhCS57DzguJ7UElbBvA6NnJqVmeAWkSwIPq9EtP37sRssfBnoU+4RZI
nX4oFrL0eZqbJ1irH7i39P3xfRjMb83Qv9KP8YJ4PzrwHHBIXdbHEvRDKBfGgt4N
0nqscWsX8LcNy4c9Ap2PdaEvJfcZXkApRfmKyFizSOyXMgcJSBq2x1cQeYxiGr5W
KkMxzD4etixJrUHbyjJrbKfrofFP1lxN9aClGKcCLfE8YEbnZCtkDM1azc0oxOgx
b4NyRDlYdqWS6fuG4pj/mJjsrxTGMVWit9x/1Tb8MmwnQp0Ez3e2rPZRBJDVWpOn
Jq/BsYtmY27jCtEDzk5OLxBebwwBBVokhejiOwZT50BTR0TyEsaD5M2RQ2DNYXGt
eK5qS1Xxjpf0AsbHbYPdlwkAjea5eKmTReA2OYuO7QyHurv7OjCvWeIKvnIbCtav
1U9QL4CpXCJxEpryJGYjIKfoO4ttqPvx4k4qyRKyTWDvg1GukUoTlFoyutFdZqS1
TqlCcK/vuigulQxIyqqLUv9tR7/8S9rCl9ebrE9zxDokXvri0xOxHMlSe6jaOKzb
SHJiO19+paCIoEMtHQ5tq1v/Hw29DQVWA68vyxRXfFYr0fTLZqKWL8FzecOqkKbL
tqU980lJO3zGsiVAP+1JIgncIZKqrNYjS0zUKHRgmgSuGGzJMyovnK0RWBtA4Ktb
2kYJwp4Rxj0hVqGyW48gzjgLhrSA70xv5qKFiXB6JiwOipbZ91DiE/J+28NMBNKx
WjamAAoKUbcaiDujPH044AOnel0pqWFv3vvtVCCA5tKevavKQlObnwXzGhbleMCm
lsCbDAO6MWbEhyJBbpYKppCitE3Of+K/lAr4x/DxD0i7HmPbbq+M3k7Qyj4X+506
L7H88SbawAbZT6C1VGai+ZnVHXR3eHg5FkLqgbJ5XGRh3tQhDsL5eUS7xEy5QYYy
80fT19FjfUk0mrP4ZD7J9E/t+4SaJM49AdvNo/NWSbwD8VXeANYKPjDySTR5jJyo
d1DtAPVKWJiwaPdW/T4w/w4eF9i8qhlZuPMtJhVCaA3WvbsNdOyQ9FG1NaKCW1E2
h5Q3IgHB0h2Ui4dsaRyc8CbB1FbyJKzC5xl9PE4gzEXOgmjdswkJpMwHqQeXOaq5
xrSdnYGy4qtuOIKQixerfKnQrGGCLjg7mLItfljiMuz+ehJk6gGdTNK8FlV0AGGB
xBb1KrfboyY9P8GRQt4Z6gISoIrzWlgCMH71mpu5aDOh2L0typdSVfQyya4EM621
Er7yWVQs5adrav7968MO4WTG2PYPwvG7aMlKQXMD1fIDwxf7ekab8yeCH3KDAUDK
3p+0qjBdW10ZPKo1xln8Hxiab3WefewkEkhOagaKp8+jSToW3nzTqlYoxnGL0JEb
3PKd/62+G9dattERREuisL+AjgYm+QCssl3QmLLTjt/yNvCm3ctrH34EffKFzctP
NNDqy/PyiPIM8p9RDPsCQzx2d9GWyAi27wMNjS94BJprT4immPOt9aVPwXKkbCdC
gBSfCdtDkJJ6RaGsT6nG5jVkTi3vvqe8j52ZRv4Zo56+Fit26oIx6i+fYMF66VmD
cwdwbCwUbzd8l8Wowiin2FHCU1rtbK9L19zI8WEiyDmhWslEfU2l09TIv8fj+UUc
4jLEl5c9jCfNngAaksEVokj816HFoHrhUY9Kdxxe50H/NUqjwx6TJPHklRSycHR+
amuqjyybZ9238xfED3sC40mJ6VU21afvzda7Uyuogk65VZYgBVHvu7gtpZ0u+dhv
fsRvCSIEfNLgGkUVn/03zoQDRpUYwSAPGb/YJImch+yp0kY8UHN9w3OsBN13oZ8E
h5DrHtVxK+5tPeJ7eCWSsqoOxHlFKWBwyOsXh7XMnck6vccbZLX5jTuowE8ksRvy
G61RJoSj7avbqWy0ptJaOtULfNqCl8aTGZV+vL3cel+KPRri8WN6oSvvIEAxFPxG
pM4/BPvfEwiyrPZBTCe0Dy9YpqfPeR7n32uy2A/hdNkcXR7pU/XP4jpM/hAvTmN6
Rk6UNTk75rnq4u/ZgCcA2tx9z7a40zAPQkx0hQ4OW2ibE8mWkdRxvlYTC9tepDJu
cUQVQdm/Q8j7WWSIZg3GhWSwCCP7s3ado0rAqjm+mT6fw3FRAOcemCV5WPkTjduQ
Sc1LP4ivitj8s8VHQeidpu2BPZDpGA+e2wJoYQkxPLYqIidlOzFIbEjB3qHE0sTQ
PYpOYMaKX/l7AaK3jLRmFJ8SAR7GZRRICJ8V8ZdaM+7/hlK34ync2JbN9ZQph6Qe
6mtAwhacxvQ1qMUo6yEoYz6OYYKYapYxoU/O7e8ri0Q93qWoOqeDpgUI2wHzIS7s
7YHbOG9HOcwZDdnWErxWFhx82bF7G171kypPduh7oKjyN8GUeZSlBUSGbNPoH/2V
Ac4CeKpRnNppTAcM0IefYLEKch9h81AeTgZzknXLIOJa2EE/zrFE+kAw5WemiwCY
tO8mtRf0m6Z7DjWA3iALWfzUHeMgRWve5X7EHNdSgrpuqB8t33lEBvZslooaIIYo
/wtzU19wTcmQbC9vXjkjRO/YK6pA+J0lrk9v3GZk3Yhdo1zs9713DRtr+z6eEwNE
Luk/bkxukW1SyrY75C7a4bU/f+LKQHufpsYQCUDAmNlUMnLvXjWPhF0pGuGZbLMf
XfQFkX+g6wAyKNSDINmD+KdXdDSB4XQpRoplzCoCV5l8pDKUmIM2pUoDQT4UZ6Rv
tHRn9MeujD5G9kJm/0lVh1/UDKet3L/Uk497LdeKzyjE0Qgfq4ERfOtRy+GEOD9C
t+nNti4D1lmGjXIJcwtzsaXOUb6G3poQQJXIw4ZxmKa2bgcM/2Sz4esxyeKPeb0/
vqI1QtTC1baVoRGtiUeZ9AxP6JkM1tFGmcJcrXLvUut/w2uhghxIkLptpK1jVfaA
PysSbyKuyZGOv0Dy5CnIZa6cs30Po2AjqHCl29yNqKtwz9SHSuv026FUu9IZnITx
oVg8pjQtSB9+GLS9mW+Ln5KrkQNhytKtfY9FQVnK1QLdH0QJL4YD7FyD9jFOt6vr
zx29LYAwbS4AZHYudLlgO7W0l8MLbqnuGZA/qcttPzTA56pzo0o2+Sgnj6ULcFUP
rrYdxtXztlk6o+B+iUT7Y7FF7UKGuIDqOS5MThKgN3MVamdiuiCSPgibPhkQ6JjK
WxXtWgSSBW31Y3dxDoSkauLdS1u4I/MbxkwxVJjhYRyGq6tImuS/JTebaOx76y69
4n3YMmg7uKyucSwawYfZLXfZWSZAi14puCeH8m2OjDk6WUT8NYj4cMDt9AbZEeeD
F05XTLVWyt++9AIwJTl9NgOvxmjE1ZDQabHQjvmD5SXHhQrBMmCqfqrJVxSO1AWE
6pfVWqibA/ltaId+KSYMXIYCJ7voeyzNcV4W88qZWw0xkzS3fizOB62KlEbyjzzj
bMPmNo7mXh2Mc96vFLX96YROn9Jk4d6tNV9D+Rcm9Am9IYlHXMblmkCtWe8D66l9
FjdiZ2tVxyZBcg17MwtTDe7LORCJRD1wXQzlPaCoYkvbsX3kwY5Zt0bsItlq0jLw
lR8b9dCxeK9+QWjMCMWFJSquQi47/s5I+XGXJTFn0fWUd6Gr2cQn8LJvxGsabfeK
i2kCdb8C0k0oIZU6+Ke+yiaXNtQHEaF9biWV1K1HFWd1TRICs11Hyw9D3LpSCivY
qix0j8qstZoErTaTpfr+2UxvH+YCH59fmDtAKxQxRgKGsS99xYB70YnO25bD2kCP
mEiOgGXc64XqyKStLoGVEyyPpM/AI/UEh94fOY7Sjf1SxH/988cwIHNg0viPBzOj
X7mXv9SWo6JRK9Vw8Z2oJnpOTlbGv6TC0nuj43yQbrELFVHVgCFbfNR2Eis48bgX
O3gADaaRV1H1V7tNrjTchorM6VxU3iLxQZBxgQN7I345zpvtw6ew9WVsWYKx0gKI
Tm5q5sJmDtELLavqRB8AkzjKibEqSvNLx8nuMfSl9iKGp9jlW/qQJvxM1/oF/hZn
2XWNwJPoQV5VKgyXLMolncKvjChhWmXLSQmF+m+P+MkYYz7ihL/ju7mol9rva7Nw
likOVLfGRSPRvfhSrx8zGqC4s76kNNGTK7sPV63hP3t+kIla66ldtS2j/G2g1lDj
D9+YiY4maQBOVZXvzsPzNWL0IRlpCVJI2HqBMBp3Iwxg72XsX7t32EyttG2Phnp/
hL+MZ7wMKPzWFmd0+eSDB/qw0l0BGspuPXFc2kqBsFEET1iD3BH+xYH/JgN5V1cH
oqJ34YTTRkj5EdY+skrpuBSyTh/lbUHAPjz4UEpW7tkByiXkEDN8rhYseZV1Ho0O
DsuxNzypnVd1NGvwG7qssdS5AJGdq4lYrqrHScEDupCsUrYaEnsUsXn3XF3jdRas
3RuwJD0IQt287B7TNGmWm1gw3Qlt/banhGZQ91yd5/8A2XDsSWLrpOsrK1ibTknI
hDElAUxhhbV/QRP2HopZuUBXjLs1cirhoVa0iwRmGcR8z93FVBSgH/w0gtlViRK9
WZNCtW4dB1npYx10LNFQeqBJPqdbURKv2L97XWCvUrsAFUD/xzT0JzA0A6s3vQGD
MUGyo+8PS6WAzeCvIjjfHL0owyOGAbFAaYtbVqPj7NUkMLOuEVpLsWUHhP3Hp+aW
ASawULcRLUyr1dh/V3u/4BlwPARs9bfN6QjybnnzYqivMVidzW+0q3LdJ96uq2xx
qlAIklr5itHf7s+ib3RZf75vcbkq3T02hS+cizpf2pvpYZEf3TMyqU10nqz06e7v
P9CH8kKsQkOoLQT9ixlbvxIzU2iC4mwOwHxxbhHxZOsrtlfpBXIZPLTxUUGnzYFL
SutEelexcpbeFVEZPVbZs7mQLyaKG2P08+b3f8xnBxVLhop5tKwVAfsmBmlpneZw
GwcSR4gJwohccB5N2+kCW7adwlOzNhr+x3zcTvROGx4zGX0wYNS1XvyP7b4ddRqf
ZG2zsU/QOVhADB9WeT+xXidSJGyRvlxh9AVAcT8Omela5bABACT4rHkWbJ3xMCit
peRi+AXVc0b+6rJ+zUzi4R7uM9C4Zjw0D3HX04qdheCoKZcqKnsYripFwMjTPAlV
cPVsO2VG3UT8JqegomEqIZDHpiKid5rUrfHj5eCCFU9frEnmwDdV7bsYxe2uSi//
vRfocNbEXNCgPtdiUoOYEQsSxA/iHeIZxyCB722MRRcepiJsnw9mfKKf0iq4yvBP
wYc7ghOiK7A6olhiWocoPqCFoANZg9UayksJt+WyKugXvYo2oZfcyOEdq3yvOGPP
q9JiVD9zUp2KNX/pWMTMLSvyNM1NuHZmz/MDqNMpkyEN56EeQwZ6O9MNLtJcldH0
FRiUIeO/NsPquixLQ5+BZ7az4bV80LjdrOZxMU48+rZufEMzYQn5jJ8NKOZkodnT
UqqknT2Lm6wGStZNVZVma+b4vCefHGg63i9l6H6whCNZyl6J6lqTxGWxFJDcgdrC
eq8QHgWu8/nMStbF+iSjgRzsE0wFlSfY7YcYFXSsSDU4KWlhmAjRqDUtxBGiefXZ
pNMxfBTiLNeUu3EArwgKbbtgDb1XQbo8fqxw827ZFErRKMgNaUr7EJEwu8mvjjn0
03F/DvaaFLbpjBCcC8EC0776XA77hZui1P9A2Lz64FiEvt0I7LgkaIRtREy9LDxo
GQAvypgnR+iSPxi5YnExs8gUwiqyGmwoDA2i8OHv8xiJsRYy85xJDobewsMmJ7Fs
05+GxquuxBCk14iJStucFSYWZT7wDxzDXBGOxJnL/6Zw7zCOii9iaXxQ5jSRvFCa
KpfvLUdm8WUlYQ4oJ5Yvr3dq/wYysfL5HWG6sDi2s/8AWxuxSp3JzvmKxqEZaXug
V2K4a82E6QnqYekbaXzcqey9k0yJ4QgPXEbnDfKsrfnWHCNVCkylmD0iltLT2V7c
JkNQzTRNzK/wg+R4tUkcFBjJ+cnW5ETxvbSI/qhGUE9+M4agIBApHpmdS57n3F7H
JxTUD1gBzC/hOXiEUzlhi2dujmdR12wmC1Ubcrg/5BJKVak3GwjHA68dZVaqmQSK
PlqsM01rmalySY3ZeunVQYOYLd9heiRH6lWu3fBzbqvnkj8QVNGZiRXFGSSSWLc3
FgUVmM9HVknbqyo4xp5mVqbkyJwOf+P2gU7aqwMLN75smC7bzf9dPLhPBfUO4O7f
pQeW+QZDlAyNbg/otQc0JadlBdjWokK6gxVAVtB2nzqSwefwKlSSMpaR5muyAyb8
Bb1qs+U8zw48aBkmsBfKuYQa8UTw4Gw19txdewtqF8JPKB5+YTlKKUi3Hfe4oZd4
FSsRmEb1wzqdFyIrXHwoVRE+UTzZx2rxytXqXHLmyNM=
`protect END_PROTECTED
