`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+opibvcdYxk4UlpgJbqGfT0WEfXi8o+wwChXdM6uV8B
r0dg1QPjql55ntjbDK+zPfsgsFPHK1nZxSmS9F+lM3AGq8Bm1MqMLTKwOAxSMLFI
9GOYwL0YItM0ijSijBEWbLSSb4BqMiWZuTAPCMcD7ReqsspBnYuJ3MNJ0O5LyxiG
0PaRjuRnQ8JgiWE/5GjfCTRAdTlQ7wEq3sap5Xs4mDiWGuhW5tu1wNWQMOFtpt1c
WIbF9/La7H2o259RCXAENdMIk/G27Z0Y5ib8Xrsh9E0=
`protect END_PROTECTED
