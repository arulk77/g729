`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePf0GaZgQ0EhnVvfi/d8tf5D5zBCj6HBLvqMYReK/MhO
svwJxDhem4HEadaN3Vlm/1NFnSfVdhsmQ0llfHLmHazuYl4PoBGdJAQ7ggzOeIAT
knFQ4oemV1JB2V/Dpsd9f6uSiZwpjaXEGD9VHimSARXyaPtancrXvSAVjTj5NWwl
vUr4vE/8aCnswRMQY7i+5T5y1tPmGV0O/LuXrRvu1cJg0okwELTeGxGY+aVedgCv
h+nc3pTPjSvUi+VVu3IDTlZTa+dOltNRGlJn+yc8KwqdTsugkuGawYGOVt0Gs2dP
7zHHPb9LWmZqWHU5sEZsBMdEsUsFnjQjpe4fdayxoA2f18hdm6e+bpdyxWjtNyUp
wPHqbbGf6Os58jZGfibfsb63NKZ+HwKcNblOfeyOXJzTUoxyXFKeD7jt1DEknl/W
7N/B8ebK7RC4tWxzIE/ZKzTjfQQx2tFrDwCkx9h07/lpSpACqfhQcEVb2XxJ8DNP
yZ4boZ9pF8ZFMU7E4XJb6BtGWXijFy2Yc1ODGPao2Z9fgC/26kSWRzpPLQeMAJWo
l8gnhuVINpxTf8UTb8vU3qF+CILF5DXIoRN/sLm4adtNY+phig3iMacsKHoOiocx
q+amCDoc6sZl++VcrcyAiYQq14KDoP18ziVeyxV21LGYzbYLvjOIA6dZJJXzPkR1
/Gv0gr4Sy8lyJs54LNN3jmfEpfZc2zn6AAVTHdYVKTIpo/ATmh2INz5FnJkcAPMP
pKSynVF6oxjxVG6pBNwAGDyNQ3ihwrUe0CWIZZLRUlR/i3Dhs11xhsGHKck66SuR
THf2P6elmNngRzE9+hqxxCtbzmE6v74aFWugc6toYh38Ls+gwMmAEv93DWhszkqb
1Nf54q74lx5uRbGmSbI1E40WkOLxyMC6QjSfyF+v5/ESAFSijUYe38oFtWghz4uf
46jpjkohZuFKr2JNHszzDwmdk9K6jySFEZXN3Y2OE+oNNZfjmyfbsis7+MfWy5WJ
vQfz1bOaTPhvuObEfLiLVCNptuwtMRDo+yn2g3mtDYbH9f+rKwebGgrmvEjSETK2
so9dGWo/2oVU9lo2xGrsiynptx8GeLTMQz7N6QVP2wBMAckBqOr6FvfC/+QAUIBY
wcyyLrKKHVX97LTcciyk6URAyKPhwY9wxqkFpIW/HzrOWWtDfHx4k4xe+lSCfG1p
x/nXSz4164Y9QyG+8NJHsgcbvIKus8hQZIKKbB/dFTIGVXLnY9h31Kp/B1qNHWzT
0vrM0d9t9wMfOV3WdrhY3g==
`protect END_PROTECTED
