`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF2DBDnb2vODZoyR5PWmfy2BR/CrulXFil6af9maQsn/
eNAJb5y4/+vAAzMFY4dtrjNEgm2gcSDQI/CabQDLZU3ZObD8SzkVUyd1FoUkrere
IAys2wXl8cP83Vk8K6JwNKD9KXcH0eDraoKbS6vVw+JqDtj6VDX3rg9UVM0cIhVE
wGOrTU5l3qNrYKxTaS3JmayLRCIx0oZQHXAuvFnDvR9aIFMX0QUhUs8l64rHoyNd
aTvNb1/x7XT2IFoGpD17ytsyAFTtmhLjAyJe2vobOVYCYFj9wsx2OzuubA3zBAJ/
0d2pHdP5euWPyt1QT4562WPnl1FYhnyKS8QC2jv6K/ictTz9Lk8ACYPSA4b3N2TY
`protect END_PROTECTED
