`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIVDWtDzqR6BzZY1MGR5KkXUMpK/3vBeUyQcnvMz9LZh
ea7Bw+xvoJ05H0AgYdJh9AqEJ1LFX/rCqzqvMi/BdMtE0zdlQmXM/XCm0qIAFABj
YWqXc/1Xb891WArMxgKzoaKyzOJiDX00WGmG+LBbcjENnEijuAWonplXjEeP6wVf
mwePS6ApVMFEe2sX7N8x6g1ngAzsdvh6wSpMVObIzK6BqBtor/L+GRvUtf30QgKL
`protect END_PROTECTED
