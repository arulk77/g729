`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMqfdwQXb3jlatn+fAgQZQSa5Qb+iGw/uzW5SWLOClSL
fnRZpYsCwdV48LsHAg8nhPg6yJ3G6zq3RXMbi8BmuRWty5A0z/E9cxbyR1P65UAg
KaP0crjuPX7s9qeexMoGqbQjXncIbXxk+4MJ0hij4YF/8jW8T07Iu7FDAJWfgMkB
56cUUAd1R7p910Uj+i+IxOk6tPPyKx+dgsoYUc4SwyIyXbP0NudR/vlqPrvzC6rG
`protect END_PROTECTED
