`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C4WuWrAYPOAXRtcRx09Kw/Y10CxGO8HbXEGF5Ln5X2TR
+HVPq994TEbvKkjXnfyDg4z7xwRby7SgxA7sC9lSfPD0YKnyNvEss0nOpLBGUXEO
PQ1EBtS+c90EPkjw5cgl5oGmj4QV5aVMjYpNESyFWkSgSByWR9g8MiZP5dPxTBDv
B1YKUOWK6LgfzFbKl08Z8gPbOwPtM3SrAV/hTHGjEIh234kWxa2VW+BoTt0GNCOA
RKr803/ForNTXS1ltIAhKXk2gcHpPKIdMglb16GVzzhtCJeE6C2tdnepLuW+7OV6
rtvunF3Obe1zHnOkD5g+zKixzk7X7yQE0XGqR6AusZbVzLERfX88fnbCBezgGeTQ
8j+F3AhVKn531MTIp7y2rNgepeqog3sR51t3bWvypveTCRfu6/68fmGUE2GQqmV2
7QwNsMSk3898ShNOGQOkCf6UU+ROT4bC7lgNcpz3qDwrNyJhkeWMs4L+QbJDjT0x
flvNd2kifHEoW3zlt23CIWq8w8pDc71FgJ7myohhC4s75/gMKl1iI6+juFDdVkgq
Xn6D1TyosEOBGxC9NmQKIcde8+qLQOZRWAa7AwSR99wxbhdl+JUn3bS5trUtv8XY
UYUkcOJKkAsXoVFCikEdEOvQtSmNSOk9o//VHDYpHlx75K7GefiqcIp7h5QtUNZH
63UjZUKDhLe2I2/10p6fDdpkwVKLghenru3eoNZAg53YMV4ySlVRXgvJyaxjgw56
iLM9CM08R2naDfxDojCUPIG25HbN3suhhknJINTNAhPvZXL3Jna+pBC1sBPZC8v6
kCPIw7XUZM9v8aqoLNv7kvcObziX47dpkAA7AF9CwCA/UIa8X3gGrgyOT4TixVCa
cWDy5XKBoI2rJAtO01v8FfQHBCBlxCvy0ZDDqc1YJivdYiSNkPvfF2vgZxePXOqQ
ZB+myUHT+u+pysLd+SzssvCebJ+A4NNnZQ3udw7Q7rlFnqPC9TK2WE+1VTUU9dkl
hIq6U1VCKhj6U5vOn5iAkkI1I03HYDv6kT8ZLwtsCcZEzmpFaCCZnDpCw2i4QXjo
fSog9kAsXHcR4YFb1xUL3ef4nqymRaRlO/KcMAoV5osYunfZf7E3DVsI6rpS3RpR
CMY26eqnlZlXaKuV4H171DiJkyRMbBiMKek3fOLqwmm6rZPS8yEWk2MUFbNxVltE
a7Q/8rKywWXBHs1CpXUVwZB7zK52c+mypU+6Ho40yZ7xVfi3v3yBpFZPAijOhNG3
63pN927ZqMJOtC2XcS9AGDzYxaiksZRDLLJpfOYdpXRU+FAoWyfxitlF/2KHHLf8
8xhsI4ojduGS8TiusuTmwh5/YC6ejIgVufUgHQ/Y26yP7gUAGGbRFA77K0kYmDmc
LS4C/V5ZxQRv6HvxcF0el4nfo2QiIq6G93L2x5xesOyk9kCrDbynudMO3NtP5LiC
Aav2KO15mfNhiinXrkjT1c0sAR3E4NUmK7hWuOwaj8zCllWhn1rVKvhFIjUnraw8
sE0ch+nw7aIAg2+ZUThnTTKXDtWZBc3pSE/w1pkfRSphdiV00C52icYfWvXg3SMV
4Z0uOHIPFVbTMrF3KJoMtyZcLxX1PZPgJ4LwNox6T+fpwbPxN2US7Zjt9/leCfRP
hmDY3Rrj2RoowBHfW9EpSeWEOxftO6ZBM/S3mXUfcA4+nKFuPslL0/PxKIIg9Er4
d5+bKyWcsHr+XmIMqtHHVUQ7ipDbIJTvVsxLsFG3MU1wxKfUB5d3zPme3W7R7xEE
H4SK4Dmk4OVYG8VIZmosxtJzDW4zTM1ZpPXjh7Iv3d22iIC54Y3bKYO8pbKRTS7C
wiilAUbzd6upII8bSqvXY6gu3JEMPDm4Zr1l70XEOO5t7xQ4lwgDSxEq9zR9I6bk
KEYJ1IqM1UXI0ssP9BT0CXNAXURe5zdJbp2IEybOWzbZ/8XmXEX9S20OKBAqQz70
sHKeZgRTXk4RujOo8EAR3ndRlrcfXbXgYV/4i2RMHGI=
`protect END_PROTECTED
