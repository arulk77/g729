`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
nrIbazP1EYTBe4Dh1zCOwck+22Dt9+EYHJ9b88ZoNMwVIZlfNN9C75aBL0HURgCP
5RBLQChtHNhBqY4077CsZMhoKE00vHqUuVDsY3O4OiIdA27TK28RGdYVSAfLtsxY
uT+Il0fyuisDBaiXHU2iXMMJpo4EFnDxDC4/teG78KpAyeeYdRiHNL8HwUy7aG+7
`protect END_PROTECTED
