`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLNZ8mXuszNr3Y5xIX7ZD7Ohe7m5EPGkrz+JxjfVTnrE
C/hMIKznjtHgS/TrbgGJx1b75l5JS34yZuXvDfjUtM5fpzT0ZXdzBPdIC/bn74sM
8Cf1/nkv8+ceU0xynxMgriBL0ztIYfF0Sss6qMEQ3HneFibnsjnEm3KJ80sZg00h
2t8QQAm5tmZzWpUE8mf7P9xfQxkMcl/R16S41YzdMaCPSXzvQkAYKV95rPaprJQ7
fTRqbIc2296OLkwCnBpVYUuw7NZqa29iYneYERDgnbaxkn9nWJIKc6KeDo3AZPpN
YK6uziFMFKda7m+c40B+R0DBjD7sRbbfPKP8EyLSe2XJIPga8lJw+yjTdzMr0vSY
a1tvWAZRCsoYg+fFHYv4wvfamLu39KMXp0Rj1A7YlCWYkfJX4VXQlzKEH8QhdzUF
FfPJxJo5ngLydVeY/f+InwIF2DrnqZhyMhsFoaieTr06QZOXW/LGCBMeBm4HY4D5
KgWhOeGreRlwYcnKlwQ5p2qUgjDCOYMOeoGPZ16TkEWHV4h9n/HNeMh8hyuE2P+R
CiZHxCkJ0XA9cE9KOvqtcKgNZC7SceIo0zW/fvzJqMu5wH9swq6VQnNhMsoX/soF
6NJsuHiySxlFri6U7VoceCd2psdOuMolVLlqPxBV9noIRZ0kY4IIbMQ2WPQP0DTT
FyNhxFwY0v00D52JSZuBkcffQpvP95QU0DS5pWcs2HJxbNknl5mliWqPEs0G2sDo
kyorbQRpOww5sSNnYLU1wnto1NW0IydXbqSayP5krS77E0c+Od5XCWXd0dsRJYXv
+sjMXvvy98fY8hFGCW8bn7JnDfwLnJZIhwLTLOIdVDGB1ilDCZoCmiodJeVR9SlY
O95+e8f7AN1cuF/ob6kPInKUTHBzmX9QHNDKx9GA8kfGEO0xc/8LKuinUWNNKRUg
bXcw0P9Nvr61tiY2ZisP5g==
`protect END_PROTECTED
