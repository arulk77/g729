`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C9aDPES5+AFe67jasyJv0peM/ImnmYOroLxUwcsg4kAQ
3uQH0ILFUb37isqnEvsiN4fT9UGhg8kKI9hglmBTetfgCtcMm+z0wxoPyx3/puns
NxvF5Lg1yHwycQ+YJgT/yHdXSTEESk3Bwa+rxBCtmji8CM7Sr5ZMranPIBJQO+XD
Y8V/aGi7zReGaKaafJ/CQkHShQdOLiG7V1+Dzw86uzrtCyv5IQTONropr2dU+1D3
J6o3JqzebK7XznpXpLkCuQOdpe9JsP7kUP9tntWgavOUboZda/TpwdfrbJDnlQDh
HVJDHB2YNRkyoSEjIfll5+3zwliVLMPj0l0361JrOJ/He9yM3zSS4zZYQ+ge6ZiR
`protect END_PROTECTED
