`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBhfLm2HMsvPX57H98xVCQLQ7YB39/IG4RF/xU7OgkwD
B7WgU2ggvpc4qF4JhvGztV0Nx41xVegmXeQMqBhqpc52ow2nxwwAgWukgD0jx9ws
oXkpFNXT5zOYGN+1HlJ+uiR2zUMwSHGbfbnni0DSEgQshEEaClZK+kgwrngAWBli
f7xMszWk1b0bR5pK0j38zM0s/MDcp4a7XjoI/NcIfI9uCtyaDjfG8eNR23v56GBG
91IpRjbn46ezulEvCCKSXal+6O/Awn6Jj/2Vycfu+K6PoWy3WoM6CPF1TtKX8OY9
bEOxeQcv1NKbHV1DWUoZFw==
`protect END_PROTECTED
