`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAf3TRSWTJNEzl18EetrnLJXN4TWN867GY7ePRW7rntk1
h2vG9mDBQEk/x5uF/qNbQje82vnjwPybNSX/SLvoKj1o/v2IC2RbxiQ1zcMu/epp
RiijwHbGkijUvJ65MnkoptRTKbvGV8k0NcWxJsoVt/2O+JOqn07GFaI+hIA+IJvH
KA0dFW/uh5wMiWsuT4C7pDZYOTOIx+WxHDvznRWAPYn0OSiCywXvBMkl21PpV+jq
ZgarVG/gayhAZgZmoF8jRXQYMU3Dffpj1n26UC9TcXMzXHMqsnGZ37PPG6y6xpuy
44W5LmkpOW00GlM6EVsw+fQjS+ABC48uaTIF/OF+Auvp3/woTp0v2MKFotsqFBN/
C9liOZnhY8N3euWpSPZAbsHYUJ/xBkBasz7ZU3La4qw2ALKrCedfhSpvEfsLeE6b
WmuD3fFmpwtNPcnUB7Y1PDDZ2Mviw5GqY3y9ZMGhjbtJ2vZY8fCZ//lRfMMaROaS
a9pLvN9kJeQ2GoHQcdEi1V+nE2lshyScMmjgnsaZu1XCDhaZZgg0Fc1Q8zPrSp/C
Xkzjb4kZjrYbw/8tf05yFdSQjiqMhNPrSTvF1BX8AV+15Z/5Ixd2MPMylr9O+Uii
Jiz8A1MD/979i3VWx+2DjWb75GGhrJaLVplzvzynkY4emQewCoUJnEV8l2lMUuLO
hpXhS+cM5OGmbk6NENPtjc8fJfaKoEFapzbPa1+BYbjFDAZjo8K2ZbWJjA2w8M4M
wKEs8dz6oKq8to8YoT4kbbio9YQ+fMXGsmVZfaz0Z61imW/l4z6y5RpfJ0RBWOS+
TaW8lpuWrLh94lTdH3n9jS9KWYcxOW5vls5BMXfDn8rHbZEOxDwTkuRFN5I97Uxg
m7lp+k5Xr4bik75zfKSo+mCyHduxCuAiZPBnzLcGFjMi5hKdbRnhS3yRohyGKHwt
rjkhc+/UwsDhCkwv7fxdcd3ncZNFcbsZU6VY+3lqTFdLyGOLlAjxt3KgN3bRBtRr
zUZHWBizo+QKtWNoKXJtqyMuucMqi4fhXEbOS+hwtUJ787rb4YfSf2DRv0ZJ+BjT
mUlmY+9akwrI0rROcedtUjmjALoFGq2ntxqdFP8o9j0OPaWxrhSSqfamhjXxVqTF
fhTYJq6NuCBmqfySiJQ0rZpwrybTrHnXj475qvG9/g+es/jJUbvf2YO65+VD4gyl
0OiHQ9JZtr0I7jo2Pyy8HfvMjif8GVPulVQtoMMgWesR1wDCeJ3NVmwUJuaL1iS3
3eLEHEWFzVqX9ZZ7qFuRBzOU3eGJ907Gqu6UOznv9l3//8pyZkrjTos2v58AdbiP
ltELp8tKQCaHwffIX1hk1W+qU8tAR3v4NpfCSkKoThej+T4Yg0xoy3CN1p5Ylc8x
x485bnyzvgDidIAHziYs5FEqYCxpeAwlihxICcBFDf0ha1eEGEl8cFBVzDnw88XV
JbxFerC6Kj4VLhjFd+mSq3Jl8rITTd4nmzgCGUJNHbWD6hOpablCMDwcTPv6P8HT
+1kwNiI4Y15jCMS3h+Xvb1X5Vry8y10vo1iejBlyBK8+0jPjoitL1cj0f9TRwhWr
Cbf+zcFqHYYeYWEMu3bKolTtP2o7C0r+O3QO53X5YL4eFJVsENNfwzLIlROpNOb+
jI6g6vkW0GKKxK5vbHi5A8EUdg+6cKwMRdq+wmge5nSIiKnTLb+tbL31TImqosx1
MsRHSjqgqm3iaq1Ushk8iw==
`protect END_PROTECTED
