`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Ri5CbAoge3yTtlCQ7uVYNmK6hMuCnMgHMMOy7S1BwG+Vdixlsugu8aY03P9d+8l6
n/1ez7Fz5zx4mnsCdQ90wb0Mlj9xPYKLhAf9gS6D1GmcCqlFTt2VT54hU8HpA0Sv
SJS0XOi+CzkawEihIFTRm6uNXv/X6oN4v7wWDTGoCvNqtY8vh0HoYeuZ553vSXJp
PiwB9b42X+wFIk5bbZCMtdX7w6cV3P0yvK2eoy7H8jRBFEhs/OblAk77cejl/DFW
vsksxQQrwHN4Qx5wHqNPOV/3HzWRQiIXPbGz+MVs/QU=
`protect END_PROTECTED
