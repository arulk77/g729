`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Bb/QUcm5QWVNPM3+fb/7XGNmGgFMoWHmGUKkTTsHWtDiJm+VGw2ailNxt8s8xxwd
3lyXgzoxFSnaxc+S9u5fDDFSUnIRNVzAjQW5UeTfcf71YrIGxbi/gFMy36pRFWHn
fY7SaH8gc5nMleBoZPftI1n0jN80vZwIR8gRZCcpKSB6PZQwkmXPqYhoC5xUF64o
+h0Hf4xrHywDiLokOoZwLL8Z8uGfpXHo+sN3Cx66f9e8ud/SSG5VOKmJ4tjtIvWz
DjkXtqOvFJrzIMnE0MvZHPBTWFFxslkQNNnRSNNpCEIKoTvOBSV8cLjXQXo+CZzs
`protect END_PROTECTED
