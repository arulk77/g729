`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
/3gERs1zVpV9UCMFp51BNR+sU7FxKSB7mvrzzoToQbcTGXhTOL0c/J/W4XLRnLsO
Y0S1V06g0KCNl7LzGkBfVMyN6qyx73R9OrG7yc0Eg6bkVOX2ePgCogwP6DtZyCgY
LW4AIXQumn3y4YESBAki0U18dj/fKg7u8Y1Qj2o5ZexwOIkDjenKC1lPL9sazI+p
Rd6eAmf81izgvLhNmHqgmOt9rT5lY7FBQjeZBK2JZkx/UjHjNYao9p/nuroGSmhm
K6eN+DBEUQKMzCwNaQf0d3NNpC75SnPkkbt48DWJcsLJqL0pUDcl/DoJ0ePuSsZC
/lzOtKZxHr+CvLleOISEO6vKJQ4t9+0uHS3+bNyhiPa0vqGrDybZiL9dek4UUHvR
u5cr3uLWV6SDoU3ag7gObwEABYS+y246JhIlXuUsr8g4rhzehrM3mURUp+rvQm4m
ginHDbfQHL/sxsahiqOQ+VhrBURV12UmRgzDKQ9k+o3f4Yq408bF5jbgTzOTQUsQ
aTOUQoRNHJOdTuZHtiHqSY5kzu5UmtISvkbv4jm2Nk35u7qRBZD0fkmKYm8zLnuD
Uh6i023p+VRgoezF+GskMcIMngJ+OjZHXEeuDHs/q5B+WKVbnoYzBXqApq3BmjkN
9D0ufXxA9j0UqnADEiFGb1tmPS0P0bdlFr53blzHOUP+Carv5AkVmIqhtsHRz8sU
kCSQZygYP/DbajHNH0iUW8LLtlMKZOmiBFneRbeNgbunbPysnLiWMEcU+nokrZ/R
0d+t3xB/HyhTkmngyadaW4fl2iye9Flsko1InZQwxY2aAPW8pDL2sbxMAsH49tkW
OHCshdwakby0PtMI+I4asezdWURyvbal+71/7qw46cXZvFpHsUIkWaxzW0HgmVAU
dWVm9zMtStZD/Yp+FdFyWjVqvTjQjxi78kGvzusVju7lgoF1sotgjfEayoX8KR/s
2ykeUS7El27jlx04iDI4ttbNoaaJiWi38Mh6n0fblQ6rIOqfroj4XLSUe4DQTCne
41EYw5Lm+9gqL0cnusyp8mSc1AnhFfYvEx1UBGiq4vJZYwQUvDcfhVo2RpPwdUfF
4KVOK3jiFoUxbqjPCLTHXNwDoNSAw2ETCe+Ztv7pWGnRKUjlTmDHLSeLADeJmiIW
QJDUdfw7G1AwCOYE/Rkyzb6n4b2pq88TcR57xyuCPn2VT0APLHPp8aqZqcSJrQz5
ZxVLZL0fQjoK5tXZCfOfqmnFMRWZFjAgIdPfVC3mWZ1TkSRX/x2v6GDV4zb/poVI
jTkQ+I/U/uvS1vBeXTrCQxzxKxXf4Iw/NWCdNY7a4tVnPgK0k3r2/q/zjRj5rKxn
82XesDSq95W7TSshVH0KVGkMuDIGv3m9do8JAc1MAHpq9HfBwGKbSd7tqVz7ylBe
YK24VolZ/Pn4DTEXC5M3AiYpPgEatTzkOxxNloTIDZa4yDDy580U9H7RLe59E42x
HhEBXappU4O1arKVo/UK4JHOiBiR2h+t2a/55Val+RZ5MDXVMuzR+WbB/U1ceRuo
4+OTctnln3ocbAiIMLVJWYMbqcCAsB9jqmG/g25svJmDVtRuDd76IbKwhbeoqDsb
efcYTzvyW3SkCwoHtPWCjtKATw254wIcL4o2KUIpeK/yaVZzeR4rntQcJE7XE4+Q
RgFbhZIjHcPIi6o2592B2jluv9nEWJzPx2jy62bJePTFjij9s6QwLIkh/UmH1o6h
2gMeHQ1EGeJm8pu+rnrs0zIf+8v2qS18w2GmoPtq2QbGFoBks7eWIQ+DUEq03PqI
GW73HPa8oc2uU48ZUTIpCw==
`protect END_PROTECTED
