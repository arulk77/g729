`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+OvrK2+u/ggRgor/OCF7D+Bb0kifAQNbf9qZDBkGVM9
YM65OEzeGjUKvoYptVjeyE9jasqlqaPfpg5JITrenM21eI84LcPtuoXToHLMV/A9
C2ZqE56Kzx58K9zvqShr3vsNUnp0C3JkudjYK6n3NW5fk6/QC2SnCV3HCOGYz/zH
fl8iD530bX4WDk1Rtjm5d1Sc/IObbhHHqzhba4poFq0ecc1ImNnYKj+RiZKCzGxS
4YelduH4Dr58Xlesrbg/UtPdUuseAzeFURcTcqa+rPe/TRPMjznNxZgDMIVV8zTO
VPpIGiVOoyDKgr15DX1sLw==
`protect END_PROTECTED
