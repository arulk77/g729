`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePWwbYq4VXZ+RS5bSV60T8GyRnKABi6v2HmGeIfQbLV2
mUwzu5v6zR0lGV7aL9ToScU4GavyYbuTlNhoW/GhyebSoqTVQ/zItvO10eb4eZe3
0I/GDwtaFk3Sb7TTV2ZiigGhL+IVAKfxEfuyCqdkKPN7Yt+WqmPdsuqSYG6FuTk3
gxMkp0KqMGI3kVmP4DQMDw==
`protect END_PROTECTED
