`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
cFzKFPL7CqumbBAEGUPSzbumSVM7VtOt2JqZpOJJ2B8EnF2ltzGU97aJytS9gzmK
ShKS94AWXW1kvgbq6IT5PIjeJJx4aViYt6qlwFHRIaDvTKklFNkGkIvrGaMZujRs
pOZGtetUrEBa4FpwzedZZVYvDHpbLqv9f2XSUY2tKbE=
`protect END_PROTECTED
