`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
9Fa1UshCV4O/JE5GZKFzCoV1DfBqUd33RgUE5ZJ9mFglpY/HWwfuWKruUoC+XB8U
nn64rnUDr+dCBLqkE9yJ7NcUI6AStd/lv/CISYJXNYHKultW4dPpJP6PhaxScJri
MfneZ5ecfpysS8DuE0ECLRpJ6BMo1scFiNeUGzkO02rvaLvgXwgPFXRZUAvsNoVg
939Gq/qh5OkH+SnFvJlkaOoJWYpakmkY2PsjaOSEAy7S4WuNuC+lcXYTB5UPl8+C
UAQglMODZvZPf8K6l0+bl5QdDWgwl/0AnFTa7qYmWK8oX/Wb15FtuRKyTBY4cjXB
C6sKTrLP+JMFLpsYkHQJV1rtJ1NoZkbMauomGKty0hb6xuxlZhLMZpuSMAWcwSsS
rjzEBRMGuxRCOZaqbebRdDqdOTcSV8zb8855h1N95YQmh2tGlLw3l7ntnx1/Dwmk
WMUzK6PH7ZJDyEB8/MJErC5viFMkdxSdqqjKwrF/mHjuMseNRpU0a3o6AVPPqlTn
f9ar1Hj3Z+CHcYyHn0mIcoru13uR7xjK6wPOwpoGX2kKRZ4m3TTaPGyIluurL2Wl
`protect END_PROTECTED
