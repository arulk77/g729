`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDIRsKwW74dhkyMx+AEz117Q5mePOSJedF3dNh4aWL8c
THVaCdBRDw2EJjEQZBgJkofk/M4xd0LYBKcprOOgBdzLfMKwuMo5ITHPleH+eIF7
jh/ChzoQ8n9/yIvNgCF6ZHuToBF7KyCG3NSqjSymHubavd2Jv8UG4K7NiqruMqdN
KtoUi7jbmH0QqS4PSVbQRQ==
`protect END_PROTECTED
