`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
eOtbRhv7WTNruIwTDwhlbQFP+9iTYYsNJzkAPn/8uyCrwlaXlsdI1nfgrVhAK9/C
7KLPASiBNTPCk6yIM548tEsfuKgClsOAdQMJtfpQK792dL6JcToreCaonzWy1T2u
rEHKcBr8k8I+dkpTqiIk2G0Yn/+TOimPifvEcZo8i+yJhXOwQVrx10rSoCgoeWEw
Clrk32VgSVOVUyZ6LgYORyjBi9j1XtZO5mRX+8nfVEnDLgpM/J5HQwSiGJARUCIp
I3CYMs9qa71k2W67p4x13Hdr+Aly7rOokaS/WKesAkHP3rPUo9ebnVT6aaRUp2vH
zqNkQxKpd1d5q/uncTZPz4I0OMVo1f7ayDLpodTKGpTJi3jyLOa1T6s2KapAta4I
4RkU6Thi+ihL/xinJZ3iPcZScyA4R4KmVxpDJyC3A6s=
`protect END_PROTECTED
