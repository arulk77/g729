`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCX0Zux7SiJRf6N5VcugykKfM3BuQagMMnuuFbmA0Dq9
V0x+vpLZqQbGkfkaOFxgHbDJhrMtXejuuoiJWOHA9+NoC1JL9BSMWlsyP8pi+ZDE
/XgDjcw3nsySSMGUG4Hq4KGu3CRtZOTVxpWaBqAPh22fKnboXabx27srAFxX+r3C
FYqaifCbxIQASL9MMlb2qHMJwqYhmN8fegkNh4bu6Q5YOgf1tYgmQVw2NDpaeR6A
6DebmuVD06iZXBwfGUyuUQ8pC7Nztb214MqUMis8vcI9xaEvdDxieZFDQu5+94m9
sqcVp6FJSB0rJE9KGXNNEqZux2anWj5r3oRbUU6QaWhCLtCWWPZS+PwfH0s+9fMG
`protect END_PROTECTED
