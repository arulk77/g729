`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBaLqj6liLDTesmxyHvZDYtGFu6vQsoYGfaJlN0BA/86
sS9JNdmI4Sit9t41FEFT/8eefqkwDx2nh3vho5zjwzTflt17amclcatrdfNptFaz
nefjhYSBxY/WAGAE618s8R+qviEWFRaMWAOGZ1+ZLUC7Q5fzgnX8SzPTPH5S4X3g
ChHfGCQ6db0OYjxVsN9OFRw3DO3dltXeQG5263W7e9lhawKfPZun3g060wOHCq0w
k8kIJPEAT8GW42qDYnevOII/6Xi5QH1jlN6XwrERTEnXgtsth663v8NvipFvcHZW
9J/wMfhABMh4921g5/6knQ==
`protect END_PROTECTED
