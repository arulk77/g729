`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePhoG8RwjuNIRT/FWmH0OUNXQQx3QbwZPIZPzzNlWOPi
mghRtkRBuhp7VA/lHhC71ugUtRlal3pDybLNAuv/vkPst4ID7F3kcdudbpeJ7FsS
QRFFjgfsLmC4oLwkMgcDvrAGsGfnYBd/C+L1iO27C8frzAyQ44QacTPd8lnr8cGV
5MTT+uh1wDMF93G3dfkQJ5P8wM6UEybBwjjFb7tUFw39pIwgTl9ACdusnPQkgrDq
g+eo69XvPb9Oiq3RFWA4bw2PZaJ2XoECb47Gfv1rAi60rgzlb/zP5nIZHBWH35Nw
qEuY/F5tlQhtfj3XIVxvRVRpVivVgFqtgvr5aq08+wTimZcYHiujUPNcu0oR3si6
e3w6aHeLGFzZL21LVpzAbg==
`protect END_PROTECTED
