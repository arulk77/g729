`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
vF3Va9EbPdacsBwCk2z/Ms3JHkr2nRmdlkU6xEIimxsWO/RNvC5YPh2KYU8bEmER
Y0fofJBJ8XkZ8JimpfvAEFuYIb2Hp1iH6CnBERezKBbxzrBGJ8KFCEv5mm9zCHVB
TU3IQBYRFKey4o6xDn+OCAPE8KtblIir4nqkz069aTE7226MJD5Z9Dbg/fyAB8T0
HLCnSkhX9vkJxxqMb5bApkhZ5uABBFqsGXMzfCzAt0SKrgySI+MnbcnfKurVS5o1
GKZEsaaAHMYE7gtGKbONCEocX6t30oKt7MskYcWzE6PfOXBLmEAFRajL/enZ2QtY
Mt4bUHnhRqn6SWnGzU+IV/3V/ZUukaGfbNAeoM8a41RShvusc2mZ5/W/iIeZem7H
zPG5RRdhQiFqTLs6D+Ipri869deOWEc5i2K6XyOwWYjANKhfb+2c9fWzqFLcrt1L
l9WHu59QCU39UrG5W99HAu+SmbxGZrfsBcGVhOJkmJTlMEliSbjKD7BQmJD2wbFM
DIG7z6EtimnEfr8w1U/RD0yU0GgAKQIUsxj4RYplBZIJ2TA6HDH1U1FHJw5o7bTo
ohtcjNlOZ+DsXDdmOXsm9wJbWL3NCPO5na2kArV/6BlVZARc7vDuA3+CYV1GVSCw
UCPT8TGDmfHoxGmRU+bYMWqWrBdkNpCyHXP9/xcE5+B0Ade0LZIxY6H9wFOA9zbT
HrR+B6tFqyyjC0uJFn5nYDOFuN5QdNoXPT4pW8TSXBJgK7KqT0yJVOirqKm240ZD
lkjvcDoF5sb90fXr70Osj9QBBTNNb39LQ+R2OsOh9ckIm073RrBuRzUwZDORZvEb
jG/SLGhOdD9Jk1N3tmxztu8o64BLDSlCvt1gxyxV2cazfQeLbcQIjjFFI2lPvN2V
sB6DwL9+tEmSkYEkIK5ym7nzPZQ6mz++LAy3bDsAfaq/ToTl1JOiCXXY1vIkBRJX
m+lXjAcH0pJo/yju/lnI6K6IeW0P4gifZpkieif/nRfYnAS7LgHWpxOlJL1xoXne
GU9fBO7HH1kmPxINfQN+/n/s+Kt/VyAq0KVBVpcrlsA4Mlpwsm6dsUnQtT3G8F99
kCsVYVUE1mjmTaya86g0BkPcQKWGGz8ONxQtL/HbDaLmG1uYbrVwHCGizggCd/6R
6S0XTxS0WTJJ9vAzJnAY8WoxxuBoBlC6dVRkBd80sk76QO2bHsytOt1DKv4S0GOZ
5g+B2CIS8vBwrMcywRzs5ShwD+LyEqCBUrR3tP7XJ/JTCpadcBk1U712nPdMHjgk
76hURxVuriiJ3m4gUPdgRu6etw5dwQSajGcTJW18oboLDgkI/L4JzZgzkxlXyM8g
F9n7dIG3AHuGPxVmqzUMVBsjg+qHzuDQhpnm3ugisudvRXzY4sTD2IZky/N8xYct
QltDlPRlGPXMcsLruo88zO2qSFVJf1tyXr7rmaY+hh3H656AzzSNZARGoFRptPhN
gwv9RLFWzMctVu2Ge+7N5324g5GzcjcOYHPZYh/s8nkT8+Nr5V6UzaeKqqKLGrMp
xgRfGf5EJcad9cagPAQFNOgr+D6ygChXj0amrVDEyVFemosp95R32Bjh00TXFZs1
JJlJgyqeOMHfrhP3/EE56ifE0Yn1oRzaLNqvwZgD7g1oElG8m3jrVqBkUSAgglcB
XI4lNbAmQrHu7tjQ2O5hKWtEZGRtOlNJrsclVw2ENJwGZbzjnea0Zitef0KqYSP4
iezVSo5RzEsl8+3iD9xWdv9u1iVcnG/GeYGyRs+dHOe2eg0iqwTb5PjMlmd8m0UQ
wGhE2bQUpExt5pxrr0bP9A6mK0t9KSr/4ZaA9HOrbjHRNP1w05ZzMsparfZeru1H
0iiHFgQ7rsfce7h0CREe01l0yjQdFXNhE45C0311SzITy/rNRkyHcfdFVe0+7MUY
t18pvNGnOFlN4C+efd1knTi5GfH0uG9dG0ZElqIeNoiFPFrEnFH1CYJst8Pr25wu
AA62YoZCH5LURBJdNOiURp6NyJ72GexjmLquBqRYhpYvyxrFTuBBGLEnt0liRrE7
W0S2CLVyWD7bG0O0QGpNdwSmCcCbrAotmB5YtVdl39FDTyUdgh2oYS5D+Mh4Oy2+
x/GYKpaVdMuLgBsaAkZjY0VU9utKjYWhQD6EnRcWaaJYpFIUT5PqAeazFPCL+NRA
bxesyswMkdnwri8d967ZC8PuP17hOuHsMdJVgOnKP/Nlso8SptncRtUaGGxAmKfz
4LbDAOHrZcViQLbxQn29qsaUvuvMrE07QvZlynTws0h3mabR44nvhrY8dB/bYzjB
U0xk7u/7+6TVmXf6FTBJpRJNvtjT0JuSkSLzz6aR0u8uUAWau80NAnlWIClJ5+I+
UpU8zyOC1E5W0kvhjQOITq9b1W6H95qpjB6+MRKHI8sZIjMnHBZVK0YaqnCctpNJ
jq3a33+AMTsw5YUXnRFSN2jlgzaol5n5Jd1Wn2qPIV6b31smj5EI9r+nUUeTt6JD
vUBoh7mZq7kc2/EP6v9D6Lp2QKeXIFzYvk5Gi/wXCet1kIcEC9VPdbxs8Rr8cqkG
GsLE61mSpLFgtw4gJi0+E2OCV0hFmsjZVqAHPR7cyc8HFy8Tmb513/V5+v60ANiF
z3JoyIlRkSsDZgoI3U3142XpMPax1z23MI4syaM6EcJ8qcJXxQvQIJmEagZ8xVCA
WmSgvuk7l+gdW4Aqzac2Uk9DLq0GaBjsWamSOhzWYAgd9BDMjHoNmVxsgOqHxUCt
GE0ttRXwAj6PKSkLO5cgtbqjKZdKTOt/aO2O9AjVzgbLuWYdniSaCPq5AMdZwoAE
pG8sQl+QBLewIOhbT5r96vYkrhJikwrC+FRh/0rtvu0nJ57LY2qNmkh8BPSCJXMf
uC7Nm98W7CE+w4q1JfXnCSDTWRY5VAuRfbNIjKo7Slgi+BnCmSPjqAOj0639r1kM
33CwXl8AbOdSz1s67hAkPEUCIJu7vW1SSkpFtbFuqZDDLUto78B+A6ZDyQKb/2HV
tceln3HOpKyjkCnZ8+1CITw8ZUNKLQzSfBGkSJOxUbq+Gh4OMj+My5n4TAl68DCQ
uRISMGRsPuQ7j3lNmOLzx68uabhW+ZHZqmtTE8VD4FFvJPM8AxCVg49SVDJq0JJ+
sJQe61r3612Oc+kQenS9ahv1lRYuHsPq+tICUTtx5VWdX4H/wHZiGFNoUVDw8wgx
RV0zBgrYtobusD6RBGDVidXNKCVMPyO1Xz6h0rh5zeDzsfv4dxe1Yrb0bU+khj73
uKrko5PLVYY0hwl8RtCZzt117cB770gAjUHcySjq5dyEnYBfDhyZyJYNkv3byVYZ
vCv6+np+ojFdEd8PY/5Zh5CeyZaJKRBodEQxaO9nOQmDHlVPisPMfdQD5YG57E9P
3Cp7n9XCZKXycUj2NfuOMlHB/v65cdjEo3i+L9t3Z/I4gItVxz7tvowJCVYaMnyH
JFESikGa5XKN5bBlgDk2CwIJl8c0cSQ4oiYWC7VdvMCf2Mi+/4g9pZdqupsqHiqO
jGSxddGXourxalE60AoS6lzgk/Zx+xX+t30YHTwTNa258zjiU/6QUhkLw55xKkzF
UMu1EgjGBldIQc2maWxgY255ExpQZJeGDYadqlXPDvohuZMW0Lv2/4LqySFqDt/r
0cDblUuJwwXJpjMNNQPbrhlVCfW51iNm9wubUpMNdGDYlNcf6kgCB+fefEDwDyPp
S7wWTszTzqmOcih9SZvj18ZkGKOAZFiERb2n9jp96U25F4G0ha7XCD991ivRjcdf
jZUvE2gQBfpHCKwJwnMh1veDJkU1krO3Z4TlYHRHkJRK/pThP+GUMjByzCHD/CSG
ibljYfuCYJbuGWWUH0Jbq9VqDEx9KRZCKWjAg+mchqQUKdQ/6aiTwUnQtRFm+tbJ
vIawZDu2T4uuAWYwEufZoBA6xtHoxx+XKlgMW2I6a/3z12o5+hC8KNuDnVqQ4IFQ
yJxx2mCvObJIFHsSoEkf6AbyyH1DCbtGZ1JlBu+iCL/xrHhlf2jUnZOiQIDmgjKh
vlkeb/GRv2LzEqzqwF+yomV9aO23yEuy/qrZdQXFIlIH12MDPkkOR/b3ZkRx25cO
Ubyx3slTA4vpeeRzH7KKrmS7QvNEMx+ELFBakwgrZ3cwQtQ3rvmiXTMz1zo+gIQ7
MnomAJ6F7W3jnR9PcYBGJf2DmSoWIwpOuN8c4N6T+0C30f4bJz23TQt5sF0ZiFDu
ktI6daCcsJuUgVDwtOvCmZHd8KnFqntaLwCiHuAe6tWlr4g4jV+y5+TIDLpG9QLv
nQI71N0ggs621fCdFAQl6GHOIqlaeH7b6ityt1y9HhhcKahBz+fDUL/f+GIFS4if
rveXq6vG33AzzKp/i/bwSxi/nAV/KpBLyBXohl2vtRb7mUg49gFNTL4ODtqY0Xw2
s4h2LYO9tEOvVFZwQqQcFnhx6LXRXy6/TV+Bcj0t+NW7bTEtAdqNps3lUFeUiayV
5xm1MrNFGU37+3/wo6QsOJOWVVqM3gBKAJ6UzmNQUb15yBo+NqUNTeWg83Vgdoj9
nQ+2Wuo8oJi3Elx4y7dGgpjmZCmvOvYW+LKVclvOQyVJEhlRu+RierYJxTQuXcjW
JHjQ067gkuRdv33/4dN0TMmWpzYrJ4mAMUO5udfShq0dTBFD7PMu0tTNnlBP035e
7hmvOWi54IHaFXoqgewBA50KoEKIWeQ0BBzrnKLl56QvF4+aK89+XwCVjHpsyZpd
1VqEjR3vh8oGACVlVoqREbfw9PD0jptb7NnUrrqpcXvl4XRsCiao6X7tapcJkQAy
VIY0/awMJnCaX2uKel7S8TvjRiJnycyZOJRVghi5PcbB/MPole00vqCC2d1AwPW8
oaiTe2EZw8dfHdMyNN9W7mzKeMF+iV47fIpuwfbu0o1PIj77+kXTfXmC0H1w8MCK
k9Oxu6b02qLN7sBYVw8LnNKacOtBMK0ggdkZnnC71itB6lSxKejVGcRNvBj+EEzN
ZFk3DbkGL+Oh3tuqjk7BsVmLbtPNT0qt8ottOKDQDl4SkMyRs5rB/wZvpdUhZVOi
iyTP+Q5j2fwD6Ctl04F1JHW8QiG2NLIHhzwlkIJRm7OPhAhnEfJ8D5+iQDKJGfvd
Us8pBgxt5GFjNfg5bxaArLY42f97PSL0vwIfczRHbr+Ck9Fym5OM8gG5nh47NDaa
+/rK8udWawxx0FpS8wa2oesCUtyCMPMNvULOLiKyBCQZpAvlncYhEsKuw++FnxFU
+qEZvoU8inTxiOzyWyVWR8lFqkpg8agcaU0CYIs+PbfzQv5cBqsZpumSWTygwMD/
ceJDnq/HjEn2YENrPQXVNLhZ43eEK2Ll3eka7ulKU3ahqkCh3MLcQkoLxNIMpSRm
eXUKPyv0M9NH3mFeiOq2tAWtsMX0/z1sfVK4n8ESFQgxQmDf/xyZUbQaYOf6JT9N
FyezjwNFj0NQFQj/G/Qs/Nn0GDvMlVrA8KkBmoZ4JE9J/Kd/9klCC4xiH4DAv1na
WIcKEUjkCwzpRgEe3lRxndm6ITViQzENsQopBAt8ycGr3QBicvQ4QLtY5Wlpn7/w
1DqfzQWYvqNh81eafs7dovTUZac+IrUSJrYQUx8qnPHghxz7U12NMPfYmIJYb5Xs
PeDRQ2JXL3LPIYjVzKU7MedAoh9CPXoh4tkcOUQgF7A4Yi5MXs8wqsDW9yhpXcij
1lmu/XTKP3bKODsYon1sGidi63qnU8gXfQ5fbwP3BgplKQiPsI9cca+MUFyCNAGT
YLRB0tWprbDcgwRkiZgRFeVwlYjBA3TyWVi4L/2guPEQwbheULrx+3YpvlGqjhcG
OJAuh/kJTcJvx2S6Ltp4H9kLu1ORKMlPtjI0t8Yz0gfCwAz3aW7trNfOP/hlZDMH
x1DZZkAY4kAeQGxlVju2XQHTR1u1SsCytPMncTao4KhIQZAC464ZWPC9lFIaWpEu
ZG6Dwytw0b7oUed5BveTfb3UlifsFr1AsZZfz1GdNpPZ0b5IjBf1XuxLD3NUZ+3u
cYIIGm0SliCJmP0y2iNWl7ZRBig7pkNfhJqLGZIvsP56hRGdWFUTpXRm9RG3amzq
SYyPjPglEzKrT9tTpfDM8z32eZ3969yPYw6wjlOSTNNEIUPOv1XUcndA2xsaPXIz
5ZPVJbz0qN70V9oX6WI7PB1g6ngKBi+VCtwsOqhzb6+UuI6m3NLdK1S/6ez4knGJ
cV82VAgG3EeXLvHHrqvd73nqZncxgcrzHj7cI5AquvivAyyrercP5NRXZ7gX0Tke
N+4pdVxFXDmcs0IWXUYJOTFYxRpisPqh1fBrSdJrH/kxntKwwr4aDfBaa9XOwd7R
BFPRbDrXlEYfEvrbOW4uuLTeRfT+70aYsbWV43y2NVJqOU3IFZ+7gNv7ZLZsBAZe
YJj1ZSqWl2+NSZC/nPlzpObYATl5fDw8Bkb8jIQeKWt4KtXs+oK3Gd+aky/eLH60
Dc2rwvx3H1GpUZBoFoNGiv9uOqsaP0s0Ca4XPo9dyNJ/5K1Dk85KFzlkKKhVN3PK
+HaDYxvyxh/baZwxp0tKnowieJxTMlmHr5E6NERZOzJhx90mVePtvszA7wlQuwOD
U47MEG97qfjG1lLfRPjNrh/Zebk1eHE6MiZtKZpByUTe3N5j6QmEaEaPCN3Ad772
+sultPgCF+uaxwOu130txdP2yQ8MN+j1ErA9rQy7mJwXgGEBFwJr0V1ibMYGWQwN
DhIIrgLIW18M6B3vR6AV8XCHJTTEZ2qtYDBh2MzyHKiXYyxSCeDy1MwlAODzzwth
GqvpikAhXkmVlwOWJA6RcTHCASnJiIkol3HplBz8Sfp9NZ96LXxb3EItdHx/vjfw
axp+sZAVB+Q0sqSVesaC9eMf+R/n17cMAuorGWqjRVqpbiT4vtPYQvSHMwkVk96l
V+5LcNXC2JFkWHBg06QSEZyHZfEQT5I85uHwIU/i83nvReAZYcQAKMQl0fRnTH2U
vmhLDqrKJZZWItfTtI/yxcFL/xFXpjFYswhCXsqG22muNH7aZEkrWNZNJVX/dw1R
OwqO1ELNqprUft1RsLSdgmDxMOBzcqvdaQq5DnfajpNpARZaxx8GXQrjl7KhjuM8
rihePms/nr/xifFwPVao52twa8SNRMx1qPLpLPRWId5RDTztLh5+qUmQjiBn+CMj
L4hno4oM52gWkr8jks5niaLWCR7hIpGIPGQrvgV6cWNL4dcsffduI2v7r1vLi2f/
RDfToGUmjO81e+x7gkphOd5uE6fhCz2FoP2eQV0k3NlME08qeszUMiA0TxZoQw98
+8tBekG6LpZWiluaS1lYeo+PW/Cq6NM39CSCFj6b3gobUc8qimVAod/ovZ5im3HT
C5cX+BWScwDZOLZ8VDdfnjNiyVZCLlFI2KFuRcFWFTwTQHjy52MQb6cy+r6BfWw0
+rL3RZdh7Qn0Oooudl+etENP2RIyni86Uz/LN2qmWw6jjW1S6bINX5Iv51igGM2s
gulCTIY9c2hZ4SlHp21OvGQC5ybRPKsVCZ45tLIIMVcxw5D/l4sii9eAG6NNWRiO
/EpSp7ASrorIbpKv8nsGWkwUzXeUFK86IN4Zsc6szeiinnwHk2M3P/KC36LMwxOR
C48xvj7yDmgk5mSA0qicW2rsjTSBU702tvQBrZjtwUPcJkFx/7V+HKP4hhOU541K
EqJkeNTy/8W47sTPehSsh75O6JXh+AGKioCljs3Z1Tv4NCWl+H8MbvoJD5qdHvrC
qljEtvgfyo9ZJiA5GzTAyxLfNroas/xVx5rRHhuZZ8uuxl5c2qJ6w3GTZs8ZY+CX
nq+gy/R3+pSNUIBbo6cPpxmL2oZ8lK7eiWjqkMoos9t/fUw5VCcW6uThBgOmbctg
Sd3whW84qdmLVow5KBtOTmYvXJs09LT7vkRb5VH/DesARd1mNDRgo+krf5Lc8Ghy
r3a4vaiHoKz1V3Jikh5b0aMJ6tJ72Wvm4/BjWzMQBrJZjJB6DbAotSy22hvRu0VA
q/dgVC4sru/8zHuGpuK/UlyLhLoABgyXKdc20wYw8X9AbFjpSEEGF8O3y2zJhm5e
LJZQqMC03F4Qwt13PcAYsU9Vbpn+99TVuIP/avhyvIa5PnuI6Z8dMg7oUq7PEkwr
SLmHyyuONgoCA9AsbqRQvwqY6SUXIOjKMkkxtxBwoY/r4E0Xa4627b6XUqXKlHAF
/VPyMwInGCPUXO/2NV/agWvUDS48bftCpPAksTq/RotvAPfhc0cTIDA0VKJiw8sv
LUcXXaDDbAJLRJW8n+7fGkXZGM5mJJXdpd+j++3FclDhKwXknx85hEiIJtEuZoar
+NvfIK3h0eDeVKxFCmy1Lxhqr53XIx36GTIKv05BqwFD2FKhJ4WefI7hMJFAcN1P
Y7cZ/2SKZV5Gqhb8JEI/vWvZK+aWsg0lomFTICxg8PKYDs2rckTtgyTSMsYQjBy6
GXlddETRVkHpaBxKyTvEAl4Jx5FuQLqE+QYw0ECzqWaQnLafMEu8z1vkRECU0vWL
SVO4JT2SetsRCMOhTlAcurY/CzM5w/s8CiMIz8cPhXoC/Zp9yuz3G8/hjBY1ayvf
a9s/jMBHJV7lOaOjzfSDxRC8HGDQ3Bou/m8dx8xAoosOfDR/ca6zHT1VPMM8y8ck
p+q21QQrkTLivFhpyTInsiOIE/kF8FeZDhbm1SR6UazzsRAbwiKXprkqdWs2vFk/
6g67iE9HPeLpIcIITkp0WwfPZ0W6V2j8g+7YrqpJO/A4sfb0YsrV5FMJSur2vWIY
WwWvF9eMnXhpmN/u3C2cX5/1gly2VjNj99JOeu3q4QWeUgEMD910IM6d+hA3SULW
3ybNcKELviIgnbCJhQmXndQBUtOIaDwONaqZDMGQKTqQrJFT/XGS1E/YvDHcVQo8
V4FJK4dugs+ycaHGAHE9uPSaIWYU30Qu7BsotTbEYFYuy262zNz4NdatsziLa7Ug
pw7O9vp7XXn6K11bmxLTqoDSC8cWbZ3OP+jsX/GHgaNv5wd21183/t7H9oLxZREV
nx0x29T/RDNYwiUBJBO/Mx71cN1x3sBHHXfGrJwBb7Eh1jE01G1yVPut/bgN0crf
qaWfOqHjA/0iv7r4QAwZYoYrDZkmNXiWrxiNufZMQPe5xHJ3G/MsefwqKyJy4Jzp
tnVKVzUUsQlaSXg+so/PgQzsQxJTJBgTJBz0GGvhBu+xRkLU0iuBwYe3SAF3f/JJ
CGXLZTES2n2DPHxV64vlqmC7aZlxHwV/DnyTcfgMY2YmiovpEibfPkjCwVeb2JhI
jZk/oXm0ThIXNIoubfEHv6J8S3iLmKhJmzfjSl8iK1ySUCfgnX4qLW/prcI32aS5
luaLQQ5vTjMwf1fUd1Yx+0ZBeVaDMT1YDy9cQ4tKW0/L8b+QSwKkUDSf/nQ46wfE
Xg7m26WQsfk/uNSpjrQYCUs2EmfANcs0z8hwZrrOKj4HEZ8WQpuz1mtiHn/4yDLm
kQytL8xZ86Dg1MjibwfxHxCJ7erP5atrc5r9EVWkZTqpDTOuII/J0Z60vxTPHNxV
SnAIbuJbt6xVOWjeZuz1axG2ldUsT+SvEstH7nsOgRJxLv84oJSojTp0JJFo/7ZA
wJpDanOZwuEsuA+0+olDvtkLM0K4dB07655zQOb1Oh9qKc9rbmuke2U4FTNzTEEl
p+nm75BVFU4hNnusmEk0U66GoTd1676ZBCyVYLc8gtDueIDMEn8U2ECh3OHEZHXi
PysBLew5R/okobZpa9RI/wmk+UTuDmNhOV2IFIEVpqtHpD6xLGyQoB7bkJT64h+i
2qt7WO4nYLteFB/xBN6mKgvunCMdS+lDaVzVEfq7tJJ8lNJ/+Fl4Ar6sIf+OgpIk
8p5Lcx/eXHZt2PL4mrBXUDOIAU3rOy+DDMUdYEZN3HHL3VN+DCOG6I9tWOs5RPWH
X8BBgSsQ6e0lKUbSz1kFXTZaUFDSidYWVBI+D0hRWo8zk1EIz/bMHAp4T+S7oKDQ
QrcTgvX/beBXIQdUwsCo/9mGZ93f3RNk+qrb6EV5cLHGC4ogbnrTH5SonfLyAGj6
2RC2QiFidbQhb7++MHyJ3mCXOjY23aYg66St8FdOjoa/ZvVRfXqPiU0vujTTdIvo
Pwj+GFyxvvrSwdT5AXtD3Eu7E4unciqxE/M+8fUfxxt7EqBmBsPY89c4J2k233R1
6wVsSLGndWq6dGtBXYTjZjy9CAvGsb/QCq4G2AobOwfqrhxEcYyS5aZA38lG9F41
C9/iaIFC75E0GgVy4TlBMLM4P94/DBxHq8YOugmCSN/N6yDdtXWQVYxeu0+zYK5Z
XSb1U7KqD0Wim1Vj2cyH6l/qjVsfyvvfvad0o3guRFroGvIZON/CX36owYZEU4rR
xae8g5//TCLO8pJk+9hYn01vYnZEELrh39zOEWsZI+DBbjOqSnv3+cYAxYJWevy4
/8AF7iNlomcdKjuhl4OffC/iqiQHtU1prU2AcyNTUsvkPmfiYpGH9dZvzsUsDKjE
Rk2coTKwsuR6FycQp5MarUtpCpj7om7Wt4g4g8EaI34Ndv8dc2L/zrKK8hxTi+Lx
QxCj6caALdjt6HXvBMFcI6sJr5UO8LbFN7ioy2UqohNHcg20GouIbHBiFMi4n5e8
bkDP4AQeHnimTe8+Ui9ewmhYFRFI34glqXIDBijOdBfeL9vtDAsuo0NipnVl2Mw3
0QFBQ/dfvzFMMJmn3qSvJPh6JyJa4UP5nZ6YBEGPYt3PAEtiY3qu4HgAkPBlWQY9
kSnMyYv7MGZ80vqSs0uiZ1N5HB5bRq1qS4yqyb7zmAOcohhV7f4iW0qDbFumFbjA
IdoSLymJSUClNL1Y6ycigJ3OnUZkZrI09fIe3yt7byGKEI3O8/jl7aVchyVXJfg9
L/JRNxx8leEk9yfphXIU9V9Ezwh7Su/IACFWSYs2/46z/yGnJIB3eHfcrioX76tK
XRF7HBFe2lqIn+7guEDqNI4u4MgfrFV3k49TBWTqbjOWBRnG3kWv1aQdP7WYLOCP
Vots3Vs1b/TJ+/8ROER00XsNl9bUIaU6sbgkpqzw72O3BffQIrbpe1kdv9jYe7Wl
sUVosuK+gZBOUG+UjsEk1aXGKmsl2Ky0rGi06DpR18RJjUWi6kG2VRP64ovksWOK
EvY+6/ASbc6ulHjvlG2mQEmGfJ4B5pqVRYIAVUPMpjmylUwbCck0VFM0/DK95H6b
S4YoWr5d96JN2/EaKGJAKrikf/ZxnAOitZsIsvIX7afHrj3LPXal81uKEu/SZmd/
JcCAe9uXrz8iECl5hEyWFnpYzQ2YFJQC9831qGHXJpqNqgZPN/1wspehraC2gyBg
QoCWAIj1jcWnnKHOqi5kurb+q/NbpKI7QqYAnoxjOafs+e7QOZjIZNHZxi/m5TID
ZN14OKQDaHSP+m1mrY31B+VIl0dX9M6k864HfeZBUzHKA/iWRWUOFT7CXl3mLmRe
G7M+1BGe0N0X4ckqsj8zUQ1lbb/wHsrk6SEI/rwXn3fNav+KM0yVIoaF7Eck0CXK
rQs5zj0j+orQJqYV90jyIREgfH83w1bJ/cBN97FgngGUPQCC1/vJP2Axszj/ljV5
GImrnZlypXCFnJZjVPp7/OzY14MsDlm+zvduH1qX7C6vF42+gE6DHcmEzaDVNYH2
zhXQzbmi7FK145muhmobMKdxoxPTqkkj/YzWCZlTXu6xHafD7M3VBrt0GjpbBeZa
cOmdQR+qUCxZ4BkK4EiMKYw2LFhUKBGKDqrl8zEKyYPazORkQhGFwQobWy9tegLJ
yQJO+iPnt0/g7gZ/xMNV6uqe8OLnr9HOrCiak+5L6VBLfxYYONqapVUpmY6a3ciS
FbjqM5h7/Oi1IAMOCtHStNsWYKUC5TwmXoZ9BWU9gh2wqRHU30CD8FNZrQ7hOSUQ
nS9l6R9BqOMPS1cUWlkEAuMZperFE2BLwGPsg+fYRuvND5arcigL3tygdneAkf+K
y1O0+4G2wC2qZ5409vXYkFEyUfu8rlrwYxxw/96cRA9qukCYKuBxGuaZoMeuYPa3
GkrojiAYJv/r98J1Z63NhwwvaZ+H2gbKLaR9l+dDaAiPAn7slGJKxe6rE5nGeofK
yjJWzLCCypHRiD3roOx2RiW2RxKsCJAiUAhnrMXfeG7tZp/YcmDlkcba865IyrG5
46/0c77YDorkYUPn7Vd56lEB4R+9Vcux3n6QRCdOaYK5FqivBxGSVcKh9StGSLRc
Za2UKBHLtzdc9BZU/aAmXWM50gUF9LQ1gvPCXYVSwt0fUitH6UQZogM/9bd3DDTu
1Rt9tltHwDVmSxXmoqc8LHgXQhojj/Mrn6UYcbaH3qdM/ratZHL6/9aMkgA2r4BV
qkrO9mfZq/7fprA49tH0ts2m2Tj8BE4yluCcF0WuPCcaaVUtdPFVSu2+7Igl2nNr
XtF10X5g809lU+ebClP52BqFVUIsBjvK6Dljk6DeIBdd1mFeow6WMEH8qdmG0k+T
wcC/c+TtZ1TZOiNzgPmgPTxnGzeN8zcrLBOhzNyY+AD7iPMMXRVOqbF7AniBPX38
5lNkA77GXJO72tVrRv02XXTgEh6asibtLKG/ALtkKRXl9TQEI5T99cf4gHGrL9gw
55mGzeSXoR5fLcfm0enFKYopQcadY0AXqVwPbfiU8jsGa/26uj3jREUH387H0Myu
yn/graD40s7sl3Xnbkv23vrJ1mavnwVff/8xVM3SraNdvtwqGSMuinEiKYsu6jdw
Z294Tbg782MBga3xt/AkFSNpU6XPymCevWnQ2lvKtbCxGOk1QEqteV5K17tc1GaM
WZw4jMGIprhll5dpsFHRxXBqjaGow6QJOP+MA900w+Pw61Knv+TWQlJOmeBTeAY/
kA6Aj/awsDUatoh9UT99uJTc67qdoAmFCB9ta7TkLFGWbZ9UaOZmwCTM0QipEc6I
l6+lFwFYtX0m8A+xDC2C6pYkbeK2FmjUupjZP938SEpAk/55TXhk+cDbr67Cjpf+
Cop3s4fA84+l9dMtA51eeo68s0RMUeh0z5sEG02BDQLmk/LixKH8ffl05iB+TAoW
8jF2sS3NHr93V67RHD2Hq2M1ZIBnCPy1tWxNWZs7RqKsnrDGe40/vGkmVKF5H896
Y6Ds+wHr71R703iO2cz+/AvdklQH+tI973SvL8dNSPEdSNu19tUHrkyOvL/KNJz1
qhWC3WizWKGdHjMPc7pUMlwUjaxUID8vfMDVLfNHV3QUHRK562zTGVjYznLnYt03
fkGiZAv1ORbYXP4qVOwapmGqejUHmOCQVYXiDTqUricHj9Kb64/HRb/s2JxdKc0M
NNGM0ejZQBWVT8sPW9Oo1OnMJeIyhN8qp8YAaJDmVYqW+VRk6vvrF7dhXq67qekX
0yIVi91hi8hWOS2cXB7KW58KMRYx7P3HwpH7CaL8C4fbbhYwMB+k/SoavbnMjmkE
dha/NRBoHJ6J0lIxVz91TnZ0ldpLfU1NvKiCcWa2IBU8wlZFQQQ4NiVIzbXmxxSC
WFGd1oNSb5GrIXrO8ydmfTjXjLUnwnTGQPZOkyq7CE+ju8YgPymwF7A13Y7zs4vl
C8QtFK5TBlbt3bogmIymCyAUKXLVwUS244zS9tZc79tQQQhvkhxxUXemTnizTcLg
tDR5laK4/BuwWHConv/ozy9ntVnYSlijHROUyKozf4pAtPpoWGwq/5d88Vjufzyc
8HvVwANU4aIwxCHn8r0byJDcRODY1g+11QnJAPosCRBnrDQirYFdCKwxmRmZM0qX
q0Rd4ncp9USopqy7sJ+z506X/z3Ev+S9G1m4Op7F8/W8EHQHcAFH7luzog/HlqPL
cTLKJKEbQEyKKmYJ7QdYnt3PW3Qt4DoxGwssDVjMpvSO1keOGpxc7bvaAe8pu+P2
/hHznp91H30YwepTb7V+5ShbpgCebFwG6peudLZkObxfDUsYmwu4EL5aTd7lvmcC
q/7LRPYwTq199PL2+UtoNKXcuP5beTfkYCe6p/I1LBCvEgMQvFyhYX8IsUI+07MC
ekFUdq2vv8Z7WcepLprZou2qT00H2+GYBvvxC1apoPUzMS+HQbgyekRjNujdVyKJ
2vLjxnocKAl0rNhXtWjQK0QvhZjRmyyerBWNiM+0fMwxe+/TtOwgJDmLJgPrZoO1
mh9ArWxfZSWKsHF5H1LTMfA6xQVh2MFyqE2J3o69Zx+kpqNT7qY4meST1XN1k+FS
+6JlV3voVDw6t7DBdZWZGZJewi91Q5hWWiNGWYVLyZSfTLYuayzgmUH9OGfF9N+V
eapowPDgnreV9WbQV9xfg6GSk8WGvA5EGxmmsxl7irgeotil0ET6R0UvcGnul+PL
/uvWmL/4zAvG5t3jg2W9DuT4Fm1fX8lOm/1Z/r71RDzU14OCjlUctnd3HVxa6NoD
U8fl5NCll/vHDSh/j3djPVCKIuoplwq/0dh4hRg+lXxORcFC5cUl7dGC+/r8hy7z
tbHyddkEci3cHKL6cq5OEgJmk597q9XEeTS45DIPg7B2u8O/T21wUVTpRwyAqNBT
Y9OPxpPh1UxJG3wSeVQF4msvUk8o0sezRtD9tivy3P7FjyU3B45FLJftUHubu3uK
U95LXLvjm+bxI0Ktm9lKQbLzM4yIN1ND8AhMmMZP4IgR7wLa6Ve+xq2kyYY/VZ+J
3leIepZhSgH9Uk+VgVotsqK8wlY43RnZhY2jRrdfYuAEXEx9ZJdM52UrYbexjNhJ
NzpWZj0o6HFY3EEHOki/5J4qCSkcz3A/zNGQPmB1ASA9LRCFrSDNoDEHWB2RL+KS
VWP/1E9FTHnNvKVWsWse2PbJ0K5QugIPRsmaEKSjREFsTcQVPyeBPoXxa9Lj3ZFI
3yaweOZaL06CsxMRdv8NbVHXWVO5HtkgHoBWkoCjO8LakFDTKrAo14KwyscL+vW0
yLJgijFO3edy6cIA7B7nZE1QyLWu+CffeZHwgEndllH+mpgl4jjNo0IN4S33Zuqq
xO6wdsQY9NBB4VkqpgJuHK5YpVEH951C/2LkS4xUbXnB3PvuIGJbUFxOJ0Kh+Lx2
bSB1mwSxR7HOIv3N6KUuD3RSWNVoafJNOAVQNNfC2d5HiR7nP8vNPgVBJem2FaKH
JoQIWM8SaonZfr9M55F1bds3qSxUIhmQeuUVGjhVvd/rQ2Wz7sNmMA9H4wbnkZNB
GevyxQy3WLukqARm+9fKrNlcKu6T6/jM1EqsjGvhjipBEcuhT30lgylkLW9y/qaO
MsTUTfPZCAeqmg2waPzC+U6QXIoo5G5TXTDow3OE0/kc8KfG2TYE3T/d2fQU0VF/
bdESN5WY7oG5BeCa6k6DEew+lOkSKnHIx48oi7bGONqKXu1MJD3eBC6FiquMvWOm
aSXaDcvuJcHv8XInWNRNRdHLTs5zLuZgm3CdhIq3KBmQjG+qbUV8Whoxh0jzFmbL
smntIq3/Ij43ZMS3+otun4nv1k/2z4ab9rjUPnXV6N0QDZWdjYJWsNaF+iRMdvnO
XUqK2BItf1qOUv7mk8TATWPEywGhvl6BA4oATLAMxuI7rp8ZsnkaMo10WQVrmwkR
4pcZ/6VjDC++VD1iFVYPaqYl/aLOpDOeJnCSoHJUbU8iMIOOBBPGp+jGG7T7a4pM
KKzQfMnuUaICoMRU59pNuflBjkpyq88s+zxrS5ZNgwSgGc+jSjn4aev7dd8Cnalh
9+aQRm6TudM7TWU1z2CREO+P3RNzfbm6UlfJStF9X6OhsgSwrfpCXxg7JONthbOT
AA5VIgOyAm9Z99UnqEn0Tj4fnPozqZGWMdshzzEfZYw3be2CO80qQiRw5x6BXmX7
aBR3yojsFdT7Ubu02HYf0gmdtUHN6YtklbiR4cCForniybD+yiL9oBOb9jrv88pV
0PqI/nOO6Kq5xPn779ATw3HOZVOW7jZ4d0CL6vWrfmzujiEXwaZQDfje+hWa4HgW
AG1JEDZahh+2g1PA2Pk1mcqU+Z+Q7Z+rzBmb3W23uPLKVQhjCugAGDdndDDA5wnY
yjbSiWJZp2A+en6XaFe7gOMBJqpXO5bw+9hWtQIlIMW14UMiswWX27QM2juNDcwK
J92kKw+ZokW+FzDo1F9OXbQ9CnezF6rCq813abAp4aohtYRbS4eOMtTcbMivzmLw
YBjMIB9aQadQzEyri7+9Ao6MCfttSA4tj3+UEQHFDINIIu7YgQ1+tRR8KRJDobVP
28X6cvavq5PlblTjUID0mOC6S7trdxyXS+/S8LKjbIHfALGESO0UO0cGIWHn7+F/
kQxZyy1tl9drARulWBHEEtxuSbUhjQM74odFBplDCG7KVzM7FwoXx6LUFWC/7wAc
K4zi1zPsEQHIHN8DcjCmr+9TUqEJmEe5ZF+1D57yzY8DylrTZG0NZfPLswqoTk+s
Q8GKm/IfTyWI/RV8RCPH2as5Dtixv3NYiQD6ZWEFcxS3O2tqZkc5RavRGdlu8IW6
6Q1h03UTH/KYLUeknFNV0aJ2vBs81EwSHBymits2FuMNaLhy/TLw3n6gnqAbntdR
9afoXuIoflzF8aNvGUfH2EQnsXGjqnyO+CDaeCACsVU6Kj9t2tllmwdYA+mNSRtH
vrMm7UemAorq51LeAZyfU6IdTRYt5uW73dy2SuV0IoYvbo0wtKRjJFX1CwZjLSYX
iRVfY4Noxp3oZwF4IHYjAR+TWI37ECe1cu8Dbs/i9GWoraH/of5hpZ0RMWiDsmW8
wbndgHQB2rzxpcyP8Zj1koUh/OTxCCVpHfD2cjGS2vZYAZAYgcbRsyIO/cSaPkf3
7GJV3A2KNTAllPf/U/26Dy6PQARKQIgJW2NfCbCpih8BwQ0hNyKdVw7FcsetanSE
Xd3ZKOG2LOK02rmKftJ3oGKI9WJJpvyDk8/AYuRBflqtGQtU6Qbu3s67cZtltun5
tn5OBf7su3pvkFMHNpI7J81w2HQz+lq5Wy8CSCbMQ7nnvtld19O7EN0I8H8e/6K0
P0yJC9v2gKR7VjAYBMSB1TlFKXNT6qwL9Lxgg0zOGy/18jUZQoxxEGMEmztAeFk4
wP9bjXZjuLoMBVZ/wlJLfExugFPPW30hQnpFrm4Lwk6X7wYH3DzVOPLyjAM2P8Z8
8ZLPVvyjuvXqB7/dEjAupvxgSDevqPw25McYLSwr1yUpn6JqaYmYiOCZenCR4k/l
yl5amx1C7aGYWt/ZlCKuIfjtT/Ua+XH4EZvchc+nFBoMcJYxO1dUBaauUK1j2+ah
gY54wwJ4CU+ZfhrUuuUCeaNZnqMBYSH2RmQ8MFEQwnfEhN8f23xrfS8CS2xT/vit
uyBY6WQoqcabGTWt43FRMd4cAyMSrRAPYiiW2crM+uOLGmlUpUIwzMjxH8q/DSy2
hU2HSTGI46do1oilDQrut6bLtB0/YUY5FX35RtdyMk8pE9NW/Z15yZ++WkMUfedl
/sBW/kT/M4jEuck41O8lvbFtrrTwEVaEPJ+hzOhaTh4G8SG1u5IXy1A4oDvHD4/W
Rh6b9ziRPx3x/3M1uHYltfpIeejejofGdZqAbn2CcqCyKvs086AERtjernwN5byN
lKfQbjKKz48MTgjAqluOi5gJ1KneuOBtASfJYrLx3SmlU6kxETLaqKRYoDXrFWRY
ohBJdqkHs9YhN7naT/Qz8/XG/p4B/kZnpmaSzy7+c27a/z/q/IUyJdgLclNNIBVY
pARxh2shKyWq9Bn4NE7gnQWiKarFBQ/ImAhWDrb7DJHJyjCg5Q+W3cf3to/m1nvl
5BUQd58obfvuQc3byT2k6/vwLmXCOr0hc08uKTVTJqFbYR7CXZPgpX32gyK2HI9c
q3YNNY3257XjmaQdNjm1XtU1BRKoq8xS9us6m8cafipyh3cxJK80Qpu6pp4k9tmX
p1QelEvkxZznTtEBRyuUmpSflexGozgFtW3lCwQKGkQ+0ins8WJxQ+rxPcH5kakV
8tRb/nu3DD/REfAP0u2rvAvm2KXMHzi4IVWE4NL/1ZsvT5IVHQmz6yyEH9fVYCDj
GD17ilqTZqY3dzg4rbW83NxKTim2BaOqRZWWHYvKWVPpBsEIqyntZEszJAfzkSBf
kwIY89k0bFQQGC/F38Jf4iMrclYGsTKT5B2EGsaMoZQsQ2rl5Q6enDn1AF2o/U6l
oEKloQI3ioZL+ZJOLKJ/uQ3n9h9fhBiiaRmACGyaX1j81HtD/hV1vq5ZmKJhoGm0
9D7PJpynn/QmLnzR56AAyrDiBRREX2+g9GD754v3/neKcAoaqJdk2tk5WHcxwMDW
LKWgiLSVQePIRIwHEZf3uVKlCnN/arZANfK00n2GeSoo+/4/yRk4e8RHdBiwr++7
g8PhoIIkwF55Wb9raGeKYsnB3hhgloiErp0F3PDgcJibBwolxoaFWXqSwkxtsOYX
ua5XHLyrWWV7uqjAAqXPJrc/e/3GfnjPi14WdMU1Jaqz5WBok++sd3YQdgAJY8hH
Eud0gOJePxp3VozP9wVga0Sk6BuZwbf0brpM6xyye6DUAJGZM4JKyl/euLWg35Zk
SxOMjXILb+SuDyC4c122yHmI5stlKk1LF4Z4QdOdAf2A3N2hUyp3Tu4QkcMiSva2
G+uz6oSu31VOl2sv2sKzS6+T9lK4Gutp2nQzICiD3JRva8xiHdUyZ3L1LfWqL9Ah
fqgteUg5UNsrnzx1x+6QarX9xyoR6GGFZs6gwLzqFlO0p1N6o9WsorxYL68zT2K2
wOfMlXCjcXDmZzDn3gZPlEJWG6Cx2Z/LEP7ONRvIq6n6ZQEnOkpzbIScktS4+cqQ
OEum/xFZ9KSUveMbXbr/7bsbfhaSOkRak19sUZRWLNRxRdBzEMamJdaj/2iQ7ULf
yKY6ZlJAdVnXfaeuJmvtMNvX478/EFTlWLWzQMQH9000pedmJdrxFwNmplOdDk1B
BWJXTdsFhvJf3JGcX4ctT6FA+9Ec7ajtUGyIe8iXRmBTsrwxxyuYTVsl440iCZYT
zCqTyY3CaMqpCRACSWOJXeWYAqXO/inkAwCkStTwL1IoYBElz/+K+kHv6WVVghzU
yXmHsruMelwo5ixjG4+Nz85ZhBKlk779wZvMRwJLDJLUsyIWQM3VfOGgtTVdVxxR
1nJMcS7xxTc58jkRNRWXgV55e07MGdwYvUJuCssePxO/G/A5luaKH156ytcleoO4
NIgKn9YoayWTYRbnWt+DdhyIuVyBn9PZ8DmH6eaxzhSyYFSGasbL/6z1kSq7GvqJ
Ap4A7wDZlUXYMVPMd/8i3L3pXUsuEz7PPDjevhjVfUQIAFtZ6wTMpvCfNfEMqB+Q
dR95rtu25++4NKiBJD787929Fh0BXGWS+2NyFtkrDG0Bo67QfiAkesjXLN+9Jd4/
zbW7rxA4pIFxeV/gpVnCb72JyfLeGmF3sEfnj0IYDebdVF3DmWm91LwQs+yXNEfi
6ogUK5JBxUf6+6aHTnJm0zEKXTalMtFfiCpd8OFzN0dnENh4gh7I+nWoDyIS6vhc
CFpKJqzZeEoebBgTP47RwNcJZakDapYzO7+0yQNvXDmYGHq5t6qy08Ax5RqEiKnW
AbTtkXOiOmK/SZ351YBfQsnx5PoIzFC8Ndf6WBZqxR+C6Y0HU3c3c0N0N5Kr1iyv
XwGy0qH7IoLC6vNRCobeoKujATcj8yaRFXDf8/QWj6sR5DsNc3MHf3UzjixAMDgZ
zvpo+MGtq6e90DuPK7bz7dvt6r2XbKrQ9MGXNVsdrMLl6Kb6fPfvnS9oTThWq2fT
ehgTxgvAZPVDnE943ylKsBJXp34vUOGSVBysZIC5IZFOjry8GJPO9zNnlf8kKXIL
JaO4+kY4A3HPB0OEs7Z66uvj4pDjJNs0w8VfF8CeLJHKAXsUhFSsQzTfepBiCLFm
/hCEUSQyuxyng9x4zXZJcexBV8nAPderND8fMVLLIGFRqG8iYn4i0HipYMvY9eaf
FkKogySnk2AsFwoiya00XHlEJk0aekXMq9SeAAqrEEFqqFzliLZpxBROGqPQumkX
hvkv7h5EReKRU6BEeimoOqgvJCPPrXCWOjrYVwa8q7thsLPPk6ucyHw8At/Wxx41
73q9w3yzuXDEfv1ZWjroe96WNxral09HVXpqibg/iqWVFhpkGj27M5eE6fq61R32
+BSNJqU4mHFxxaf5h5ID8l4lLxjRxuP4+rBtZ7G2s2MDAqHhUy1ObygoIYyR9nMa
iTZVCKUJSaJOUji5asNlDJIW71XFrJz1VBpJ/AeO665xVl9ZWcNO9bw/GOdVb2ma
ZQ6Pi+MprLT8k+5+haTZwySf3CjirGxhSmVn0aWFpUQ51k4LOcWhDR5myEZB1n2g
iQqTSzH9v36vGV9O8o/geFJzG1bUAXMgJo9Xc6V8A+Lu3cCNT+BYowvHYPJ3SzVA
GsKMOgRIVdnLMqdYJeQ3+cfpyOodvb92jXKwGrTNWtRJPEscaffbaPvTzRo8odfi
B2B0RjzACoYBUxXne2jbA3tvUGbnx4eSzp97PkDhuAKVCRcx2fAhaDNqklEJAadL
RNxKP30Y5t0OigbQU2PzyN34OZQWbc/MoQYooeYepvNGHsvmhl27Kjv20AgMFJ/y
t5a2bFw47bk3oAmbjx3ajresPeGpJF8BGTCtz8mZnO6nUBpbYN4cKmUmP+1jXQno
gcnQ7drtkEA8EgDqh1U3eIRzb0VlIZtPvHzn2ZCkIzUMDqjzqoJCBdx8UC481U0O
Z9wUwteWbPdXz/Q823zgLKtk0H7OEJmiiqIxQwWDdZ+lhkKyJnovDUZDXIE4F4nT
KdSaJ63UWQg1VPhbiV5EL55SwP4mI1SfDwD8rWSHYbU87R8VJs98bIahd/xcrTv4
+PAc++yukORmvy5S0++snENHpZwM27JE79/qnygYJERw8HQt0JZmaeJIhkKirP2Q
yKSXKoGRzaw3jTO4Z2LyvkTSY6/jYE6mQRpAtzDmSrOmkdACDVkZqTG/2FQK0ss3
3EvObWiGNlfldwVOnuQju7NSq5QgBvb4JVMY6JejXeOdz9LY57iViy4SaE/pE0BL
LtWUhR0aFJKp4VEGQGJ6x+rshRibCTbACv7InIin5ru6bTN1a/tYZRitRJzIxAjt
L222KCXoSx3IZjAH4vmoKDT21GynRYBjRFL7KCrnU3hdt8ENkXo8rPWbEUyy9qge
N1acHMyI7fNW6yw3OpwvbuuCB9pDSNhicoxXLq6t/5c8XoxHfZXLHrCbsNBbfjZp
GE8fbB2417ij4hPDffXR/SrRXU9VNh1YcQFqLPWItm5a2CBwYvrEfcXewN4Jhku5
tUI/+dr9j29mtQp2YDJu4h9QWhPtsI8trGlLRP4r0mv6ortkCx2f6/BZyi2hLsmu
835mPilyVidxd9JcQFGpG6JqlffXmdlBCNu3idGEesg5Gk8mlni3ikgfWHSri9uS
sj5iU6jlC6wkmW8lCKw5glwqUMZp1hoxzNANhtJWRVgw1kaTkZNF9kufrD06Euag
Gs90hLTP/Y9MJRFkly6OQQiHhyoTmD0LQm899d0HbArL5mRFJEw4HRg3DmOpVbMc
7bv97iq8TIfI2gn1gCVC0vxhsEJHLEOH2fHhNW/Juzi7gnj8z6u8wwL4brpH4UIZ
Q9SE2no+wGPF2oq9+eKTkWHc6msS7wqZUT/mnSi22ZTJIbH2Ymdyjn0DcusJ+S1u
IjOQLlwdfiKZb31Uu8flynEwbAW6ECB8G2cuMPIedIGp8q24oU9IR3gi3DcHF0YD
JQ4wbVMLqmZU+wgeKkRVoUr4LWO1o+T+M9qwT5Hc7xbkBzjPjtjsybg0HgppezdW
1XVAufmIkCfFNMtXyx81KeyWuVljtZmeWdQAb5MdchyZ5y+wgq1FESjcBBvfo0UV
aJHZHfSKuvx2V+BP1kdS374zR+SOLkHArh0fL3T6r/DmymofzWvAWPWo8wdNriq4
NAMXoyXgaSofumX42d/vJnSQgraNpxg4cAoZaOBpCG/w9EFe7Ry42ubQI4lXmCml
OwFvSfWGhF/xaUz1CP4CBOy523SRT0UeyaBpREnjIuG9HyAFUK6lHB/6n6BPT04x
aZNJgwErbOXn1YzNjmif+L854l3W6tJ3bHo7LRzCZqi4vWbFjB9UFt8Qj1nI9TCG
GMheaa0I5xxM9AmRkF1b+6gpr9O3zvq37Px2dfqH1xx2g2QQuHwbk9URSJDVWM/e
hdT6BXVsmWyyLFxLhNWGkPA7PmkoMe5S31bfDJOeO3o/T4geGRhmQWS06KSG21Yw
eOLVeZagDIExo3zQ1J5F3AFDmMIodMIaue0LbUU/3FoToATxpqNI+eqJnEIfWKLn
TIDfCSYw0Rad8NEpQyvWiqHFAc7Lqjde3/pSaUfJHARisEGJq1c9yaQANq1Ta2Xd
uaFT/0Vm/AfGEIX4F7M5RkTL2vAo/rd7wY8CbDmvzECMsFtzDzwPmbsliq2SoPMJ
lfo5PBQ/gr739KNa3tqdiSjN/yQ8LM2LAWZlxIbV4ce+w0xs+s5DcjyVPuJgpxHG
HzuqDJuSpNc4RM0yTwrd0FrGQuYWB70Aakc47YCAcahKZEIyU5+vSsNGaLi6ojdP
Sjy1iKNhxkFytRP58toBlY9fjbbRIzfpmKqfD7pVszBx7QnvPLGa3AVIhAJTTLcG
l6gNMFE8aSQmsS0PzYpo88Tr+eSDrlWlafJ3fTwCqRHGqBOpKctNrgA2orxYBilF
UZA2mZ+pyXGUiwVmpHRyRqx83GHpC1hktWKNdCei2OG03tPBv9qUXanhPpME6vnW
6gO4A5+TDIcPMBbT6MXNG0jllGX2oy4btgQRbE0l8o2PTGaXPtdCTWsbCrxv2wpZ
OBGzhBtHSNx9Yomza9CEhr/xn7bAHeLlvPZVqFDJ/NMlWsA9kZbgjIH7jdjavTK5
gBD7CEXKtUs4uaTL/imyY6p7Jsoi9Bc8i8tF71yC1ZIMTSdYoEp4lvnOumJ2WYH5
SGo3A7wRpDskYwwYRvpcHaak5UIBiVWQhDrP4qyzo4fuuSfBkmMZvA6+H87MIf6x
vYJe8UV4QZiVXUum+PuQ3BkUGwa7xjagk1sU4gdCD/gjqcwBylmlnxF4T1wO0PH3
QdBX9dsovrTTHBACRHO7blKs7i5gAC+ykLlyjGJkFJvzxbaqkv9EHiirV59Zqjr5
4hOk31zBB3qi1uwjKe83sjl4sEAm+TEaKouKcS7be7IKgJeNhWnr77IAyZNm6jBX
MVrT5utwXF73i+H5zrOdl1pQuaPU+J6KJq9c53rVGLKi/bGx5sAZyqZ7WvplSASu
0p4U12QhGWE68BccXQzcgC5u6csU/YwBp/HPPxZcYo4vMbsfV803FjBsZh29JX5+
79pLyMUUiCQMOaak3v6c8puYPbx6Gjaj+HJY4DGmpM4GG+XEvYs4Nql3QoUL/4ZI
kXJPk9ZS1VLrM9COhrNZDRNnOG44e0twXonv52Yd89doW15die0Uf3p/uTyP0rt6
UJZhR19sCICvWUhLtHtdwEgbqb91kTm9O8pvrBls1SQ5NgIc8yKx7VvEthAmW7M/
9OEjKxQy1jFwPc2s6D+6EZDV2gf8QXtmG8vfKMSv8xzWFghDj3jIFpA5FfIzGIiB
wCCPbfrjyUG2VIhMMfb4le6sCS3ULAj9FxGf29eleK1JpFdAuTH01yemmRzcz0V7
WKVugE68W9oLOFzZnsjctWRQQ0h4k/DoT789okhPsxt2oXeWAqH532nh4vq2KVjH
986YbaQTMRqOt2iQdLFRuR3YoFhgcYotmoYFNimQgVrhcj509zE4RQydjzvhOhtk
Dzf1pf8uNylfKUMrt7wJm1fM4axBm6V5AHXuDk4Y/bNNEEypTTlfVtuh0uEGQi51
CBW7BD0LxIp1j18l2whzC/CkXwHeMRvPnDlfjjuzp0hX+8RJzeODNEUzVUfoK6CI
H8hMc561hOrbI5uYMCncIS3jyw1M3ZDSy7pWn3Taj4LRudiEjRQsegk6sfYNcVJo
aRpDK8ClDyYD4PsHVdWOkfiDSoints/h3Hsp0x2EUbyd5DlEUohKngWLHOmZ1wWW
3BP4AjQOWQ5ak+Jro5XEeQNTlr5DbCfaVnE3VdW6Im6XQsHhejF+aH2AH6F9gwkQ
YwJk2NP/QhNlUS9mCZhuFcz5KbQ9ZtSi79Pe3RYHCpLwhaaBSj/cN7l02FbPUEiM
1zq4GUxho3a4CCNw2uz0hmfM1Dl4YZA5bFLN8PKpjda5PWuGCAntL/aj+9xQDZEa
AnsPRzupIJdca/0kZNXS9SltEM3zRyX58D9nwm8iPB9LnWiCvRvaKzjTl3aqrD8U
USoRQJwYCn8mjdGZ0t+Cub8jPzHWzIUxEs/9z2PkjDFYOGhuIzI1lOIIXUz6sZfv
32IdIiienF4TQ+nB6ygzi/BXTlUMosQHfsSaGgq5NvK6jsTsAQs3p6JfkZmsXvej
guuCiUwkQbgroMqd8yZJTcp2QX2r3y8eOwPscZiKDctK7op4D/1oRdBL00mnWsAp
R0IyrIbJAAswi7Ex8I5/HOuuNt7CCRTlzrWbWQL90gsj1CIqLllZFIg3b5+gHx1g
QZn6ddZClFH4YuREKbePTmwF7B2wKUJMj/ySEAComvATrIDj2chXzY/7iaOJzVPT
1ujAdlhjLzmnix/pE+PPWAH7V3eCndfsSB6zDX1XKTVDKPuXo3Kx12rIdsPiBl9F
axQLr3lJfiBtRwsH6gHrxb+bfhkgg5JZ7zhA3zuXj36td3ZGdIAVWW5gKAFhsQTA
GWZO2ZXGl3wI00GMawNyHd76KIh4Qw3tsoNM3bACv7UX9PJntBmqamlONqs4yHk2
JwdQKr5lUzVMEWE6PMc8gDwai8dRNzq5mp4/aO1Y2kdYdy4S+V6dGxtPMRWd3C2K
srX0021tCwnLCSAtf/WNJlaArHF3X4iIfmUZFBJ5NotBUQS55ihXeiQTKoN1dJ/x
eCVTyZDDfQ+uTw96zcURYe23DYKeiZ2wNSmHOPUzSHbaGA1UOOYLKAuBTHKJ5xoI
wtlZGo3YmDpRHLqYuu3W7V9VFmpVG2kMLJKv0gdeDi3v8kI02qee8QwRMM/+LXQ3
dOHc0FzVrVZ9ay0dgpSHDDPvLFmKRMjfguCV3EULQCD9znhDp5oPhRZ43Ifo4NaY
k2nEuEw785YAi+Du/OH4aPjuFi/yTd5k74UOFw3uU+aVWdnBrxC3w9kqx7YRhwM+
ivqBEKOgcRSp62H+JXtnvRwwMwvRwISjl6cs6TahjO7UO+fVMhzlzRP29Ln/doA8
+CdHHfO3Nqm1j2V72hZhdSlrex6EoSD7pE6QGNhIOcYsVsuLQldtnD7D+v3qRr4l
U0Cl+iKwcIZdDid5MLnAh22wk+OdmXqBy/+eySazVpaDxEYakJjg1WFitLbD5af/
knMs5OfZYd4IuJof3JSpWy+y7g2aVgfk5NiLAaddW8xYzBmFHJSlO2zqyU77QeYv
3daJuqKrWkMDxLLeJkqZ97D/V8Gnj0ScwmJtw9mSTIzk+d2MjJNMI41BnJPkpBZC
9a40yxy5efWVxkvRvPaUg//ZVg0ES+syMF3Gd3kyEFzuuj/FgMeYUHZzhHLx5ri9
72BIdhuXJm4UFXj7n+gxCpe+8Qs2PX5Ig7B9BaqJ7NuD60lsd6hCLka++0bYnfQV
WFMs9lQMWZ2w6DY1wWTKpQ3uSvoWPzAW7/TqtgjmPo/D/r3oqo87LUAhyx4U/JRE
SKzX/M8DwkHVJTKHd6Woh31VibE640a5uhtsYWiGYDDi3i3ZBYVqMo1eYwffGq3i
XAqxzbxVYaRZ8gglfQvG6BrvWlyV+3xoo0ZWJpWZ2VmzkybYBf5hiI6ca3o2o/Jk
iYxiDyEoWAgG+HRMUfobNCo0+A1ZlYczHjjeXjNmIFhAeZHUHctJLRpHUo9KCk4f
u3ZC1ZIx6Hu7QuCWb7DUu0k94HD7RpPd0Km1cJmSEr93aCD4Tco380HRP0a/TDfw
KcWiLDEYe4mvYe+x5wiAeZjmj9sj4tErN1yyaGhkN5gLpLG37P3OUOKSzHCeWw1l
hib83x4o+7bBE7403QYecC1irAnYsbSUtlYOyLa0bE8Ar3aIdJUZ5GlQLyKV84QP
PeJvbrYbYMvUjX76t55FuPunfwC103CoaOydBPj/wJ9U/z/T1gzZQIuDbZ6cD1tT
T/Y3QeGuTYOFCkMrSGRF1/3BLFJInzIqimSKEG1gEt62CF6MZS2CfpHHOdNHRJOW
+ZQFwP799/dnljkgJOCWskdsFEMzjEZCehDTB9942xLginTxfbI+WR3L15BzY2Eu
cRx3SVoAPc4mxOaM6SZc+2cYSEfBy7vLVbxYxvKjJnYD4LxXhjolF7tRNXFgvh4+
T6EXtONZIVmM0jwksFtphUSpdNoCgApTblomVnaMQauRJVr4UHpw/mFa2lQ6RL2C
/we8anjGuYIGxJGTwQbApESxwKNkBisQssZFCUsSlQRgSAchX/1gEpRCx4rupaOv
wLEp/FzfAhyxEY9MlT0Uf788hWnCJwdQEhN2Zc27zGJJQuyIO/gMNeQcaeYG7vcf
K40lKkvTqHSJfU6+9HwjTXeisoZCJsXsKQmcw2TWfIRBXNLkEEqjemPSdSzZ7JTG
+iBHF6pLl93W1haft/5I/HVI0gvLvdA22rMy5ddrr03DB1siqB5TDJszkYc2eS82
1ZkItjYqjx9N2AosQjhBs3Ne4maNmc4wiqIcnThQuwIPuAX+7Gu894p2S6ePucA1
UPXO/gHcQpJC+mNQj0v0BvklzRqpNw4A05MeNkCPJIKdjULEPBAKHQoVvxgMHg9S
DP2olrBIvX4DozMipCfR2Y4dbG1D+MeW8SCmWi45emJd7ZTN7Xa3sA+1o4O8ECPa
h6bD3WF5raPpEmOUjiKDpMR7rMigh2XFd/LVz6oKLziSkTD3neSTE6jOMWVR7tLm
vq8qu61UlLPq5PJFe1Z6FiTRRCJNXIO1457I7zaBAoxqY7GBcyWU3RMDhvTKTUgE
bF8GJBWklECbgYZaSqErz9VDZcDNxqj+g1pF5WnAAX4ID5zBwS0lgJAZ3iABwZLD
HE9Db2SqKmIRFcc8Q/jg8NOqY3jj4xf2FSgnWVrk4CdfOskgFLe9IZFMcbjKomtl
SKB0D0i2cPR0Wh3m3sgWyRuvx4+BMewtzRfSL1b7bDkrAREr8Xbu/G2ecwTtVuXR
Vyf7xbBQ5r6aamPh2KeILVcgzKbPVwNQ/Rwx3nMWNF3uJSWlIygus2S3Fzc7ELDI
AcM+BBvyf2DZIdOPnd4zTiAGmFDLDPENhTNKmn/lXwL/qThbRj6qYqsGp6UFeEnu
fi55lAUp4Xq4GKNBPgppnO+1oC0HtXCdiUI/KLdDE7BT2PIjpMdS5K/12uOeM6w3
YKYVOn5iAwOiZnhMKihSxEoU5SzqPklwWR4Hdqbx0g45idayH2/4nlyffaWiMJ9h
0+1EhHdzMQNG8LsSZPv77HBP5CrBAGYxKxnTwURYu47AE+SES10L1UgUSfXsx6wG
aVbpzFiRHW8HIZKUwv56K4mMpJPXxGoZ8mWDkShXFqYqCC/89/k31XOWg2A0ODsR
6i5xh5yEFqTxT2yseFqYfArYq1zHRIlj/W4VKYIUDarvFEKzFlcUO2WNK/Q1Xuzn
L9RgPd+AYF6XXhvrqaq5joMJ9wibdTHK8b9ubQDOE2Ry7sh+wSB2+db4kYD8rCAo
fMUbDna1g6YAv+5EqAhy1f6rczQeVwnPDEO9zjIvASxqrpQpTNGrKrAC6u+CAbWe
p5nf5Tq9rP8I+2KqNeLOlBnrLEkAJvJcvVhwgThoJ24Alm8+4oUby9sI6WFfiHhN
P9PCsbcdpz+Bb/hgDkUvRcXAU+VsnDJ2Mr4zhbkahNhFczpG5jae9c4HHE6b6/yS
erWqDIkLh7mBy2N/VlcNoA3sOUT6CsPmNXfvias8M+QGfku/ifH/QRnpEOyaDxi1
`protect END_PROTECTED
