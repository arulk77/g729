`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEMT1IRdpoxdRuxWTfWuieiGQNEDIfTcbG9FTrGLo97k
j3r16OoD89AVr/B6qJAM399229/yiegVRRjANiJrSJR1kQZLe6w+bj4Kpzr6C7gK
ncJE0batREw/a80UZGDnPI+3XvXqYPSrW1/pKsp+aLA48Iu2YuIPJF+9kolZ+HV2
ynJmP1pdBzmtQ3q7bwgVIlBO6GNzhI+SbbLy5k81NAKS3GVIW+jbpeA01rU5y6te
tTN5mPmuZ/QQyXe7nYCTdyHYgZwwiH7ct+ErWnFJeStA6INl4QyCsC/4WoKvC47d
bu0ULLDz4kHhbO+13tQeO2p3dhDOk5rFNvdCDeyh1x/vhy7C/8nUgg/LWzMe6Re1
Kf33jeG1fVxvumeXTwB70XKLr8fmeSJRmzF0PwB6iWEbnFuYjfdeP5xxtj5GEkBt
+9iI6G/kd/uu8QyC74nWFoav4R27CpAUqe9aApAAa0z5x/Pfr4xUTSZyXrW6ilvZ
`protect END_PROTECTED
