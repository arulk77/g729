`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
FkXxhfR7Pzbw3iaw4t+qi+zO/sY4vAPWuU7Nyv1mVeA9iYloxLibEmgebin2dHZW
CRi4AjQG3nFPdVLh4J3nSXriN4YfYgDvfWLm+Yl3TL6qPB0MxUwjZrY55J4aDT08
wLY42HVFOkJissw3OzKxRJKAX+7JXsYLcIAqPA07cSHFL2EZKYaAxkGEcn5Oq+gC
nZ5BG1XEeiDmVXq4RqCvv6iNp+cyVGxWaI0ypkYpINBZUSY+nJw/jXWuJ8/Mud35
oqDynY0cWGs0M+cvzS3Ro/KpXBywLO471z2EvM295zX/ull0gl6JA+AFmmwD8fEL
bMfKfvFsBjAY1EKysWvlSynk0uZqXXCOQRYWU7Z2kvk=
`protect END_PROTECTED
