`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
0ajqx7GXT6PXYzUZrqS2WGLCNIDuj5w9H/UcsJrgOmKLxFI8BkPPVOGMM6+5JFOK
Yx9QMLnKihV1TVlU5x+eh9l/ezLrxMt821httt4COtvytbFj+TYUhxnk/PbzN1Kj
mSdmfBSWghFR8JudJ5HxrNC5Wa9Ef5ILoTQ47vPKfVtqWLCOZG5IYFZBGDPL13wv
zfvANFJf8aw0A/ppc57ejIQAdI5Bw6o8/27C5Ff0OgOEyjRBIIDvn+5KidbRa93g
vsNFEGoAbJOnJQIqK0cUZ9teJh82cn4spBFQY2MJSKf5Lf6k6zv4zEBeTWKeYcXG
9b8t3WptpfRDvN3dIQd5u7lL6NFRotKbjPj1zmWH5ys=
`protect END_PROTECTED
