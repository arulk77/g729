`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePRYmZ8kEbo5hzfUkIDgi8/j6MW5TowxdpJbvfjOKtEw
fDGHtsmLCiCHlibhOnW/Qsf6y6N/j5LOZdANVlrGihfVzpaDfTZDKOfuBsdvP5Eb
0SPoHubn36f8X6ZhLfDdJNEEiOB4gfG3R4fx59gHgkGmaSE9YTjIApjiXKbCRdvL
NoDdBHOGOh0GaZNjzsP5Nc2JDwBOAK+qLwOW6LJRxwRy9GxJseiHCp6Comcqt83h
fjZ9VU6IC7KmUf524FTiPNhc8WtQc0C17Vv8X2PXfOhxRxgxBVBrfAmTL4eDqUEB
AQm1f5bL0biPpZmp234faX+VVwSTFWS2KYVCG6ts6xceV1xlmuUKDMyJ8s0cm0UC
qgdIOJW6nlCUJ5HWbwQDYib/yrmDRh1HpsB6dFAp0QTox/5utZHMt+B97aJptXkP
KhlTDa5RFmxw1WqfRrzhGU2J0DbZrKOUvmn/P7clLOSU50yxkTUJPS3Lmf90TxBT
ZSbsysRhz28LZbQ5udTBJcgCROOwHNAZ1v1spWPSiokNErTf3rEdPQubkGWlZYX4
`protect END_PROTECTED
