`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDID7x4NybP5v7RS4p4CQLmZJKJvteSudvMX2B+NC95Z
jJ/+IKcSyXEBqJAh+oROi2PitAUGnG44wNHIB0gfuzSBKSBIv3d5yDndmrjiXRUk
xeKOAncxP0CPOmsXv3bB2bG18arPJp3YZJ86GmuZ/5sOOUC1wJGhAG1eOu/owT/A
t/mKXpVfgV3w5/kKtqm017nIbUyD5gp3aR2BtgAuzLz0Jxl5iZ6p1VQRkVd02Bbo
TkUxTDrTxVv1jI8dRKgbBRGb7bUgUDv324/mxKuBBROWd1q9mMdYwb39A4ptL7yg
RstPAIHsu6eSUtxBWF8nChuRNY7VnCEFsFjH0Zcx4KfxqmozreMXz1jq52YeWzTh
ZJ496yjOT4L9yzDxMyaXX0gS74avzBFFwMeurXt725ldd+xN2uMOJgfPv3g+X/WM
`protect END_PROTECTED
