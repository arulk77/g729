`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
xyh4ebcoKCLz6Tk9xGIV8AKpriQcmzXt45hs/G3eY6h+7EKlPO2/F3gjCkwDg8x8
F5CNyEBU9eFT8duPdubZ6guagCxnGogrwCln05ytWBe7QQCW0/mF8oZok/AYBT1p
msMHnPYmlePoZ/fUuQ4j3EIU7qMjkuf0J3YbkLAG5SPSaZuAk9B5CAg/wrY+jK4I
qLJBh9RhsIzMOKndielE/24uSUhG9m8N7izvFGQnyXHbWPydF5hSgclSWlUcel3q
fp1gtQDjsUDsxZflOXh22k3iTg/dd4lQn2IZqqAggqWXBwPTeOG8x3QW/Ipcjfqq
/Wu/+G1LkMEXRdARiudPbBjW53sRIZNm1dQS+yJD6hVEt39ugNtVyREzRh1RVPvu
JZ4JSv/vHl5yMAWEyJ59fJAkUeFIvmweIooFnifrYrr5nT/I2jXj6LHtKRxX5h+r
l3nvFLXTb2e44F0wv1aVDzDaxPd8v+XZ4PV1NKgmLz8e0YeewVnKXwjs4t5fBU9l
oEBskBnAJjZIFDfbGskERw==
`protect END_PROTECTED
