`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP7aRhQmNJUwPed/cRvHf1NBzHTwPE7eisNMm1OS74Nw
Y1Qfnuho2aRK2jhqe9IKa7ZdC/+cD0wCR4NXfXRmXN7NCWTKA5CBUElaVu7UieLy
PXQ2C8Jt1zgwBqs13LcFyNDBVsE/2e1m5F094wSfjYyxLpYx92ZWLvi/iFtoQFfQ
Rh41BUfOgSSZ9YHmIu4BfRHp/XTLRUvuwFJqJc/X1dd9Z7EbRNemDT0awp+x8qev
pSUBHSbZljq2s8vQmf3eJ1DxTaUkp4r9GVId3z9Def8ymNvjS5n59GqiTkHelYJh
C0aKuY2nmhq/I5t2wuhbiw==
`protect END_PROTECTED
