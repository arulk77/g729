`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAV0eG9uZwkentQEhZ5undwqAPaE5jHOx6U36BwV+fGa6
99OhN1gEvCZ7qe2TToCZNQB06owdbZWoBZR8OkcOXRB9BZslTp8PZhFENIJc8K/u
r7vTKpDzjK6U4pLCnssErh7YwSqW4FAO0MIjim/Kk1eBR5GAzrCjQIBw2dcye9qZ
lJJUxDoRIOmJLZQ514/86UCxNfmKe5wlYaSXqhrtnVTw7rtnH+YRxYbV2PnBwppN
Pefe9PTSqQhVFPg8nFKOFLuC3yOuOwhnz42FgrK3iEdb2RqJqj3WHu7meXLgfMs/
XpFFQVsMQeDb16gmr1Vd5QXvxLMtoyBVXqSNV1iSTKo8x+pklBFhPcllI/PHlSuW
ZQsMJSYt/bNI6BqOZUeHD2SAMfEGgWHH/MDoVbZlhcjecN8nu88uGVzPFeAhHvnT
fI7ai5qTuN6dl1cmCM7FcA5hoPdciui9REqy9ALJ+pMceucNQJyOdk+Wm9I1nVi+
wGwS6zlWFNMQlK+w+f+3SWvdAr5UahRKwtPFz81aPyem7Rl0B6JpSNfFlJ0sPR8k
0+59GmZTTm3UbgCI2px7NAY4MGqr9ihpFWuc+Jh6UF84t6uhe528QKXhH7hve+Ia
/NXqofHiqaadiIXgMb7iO73DvKv3CKyQcbcymGuJrNfcAZd8NlQX0NdBtX8F2EKq
J9qftN3uLNIeVHrXPswTAiF7JfKxU4f6Wc1UrcvXUT5IzHeFPxlJ0hzjmxi8+3oG
nD5D1y0eLY/ESj2Bu2/MhvYSLqhdlfEM/nmvBS3JG8kjQvPFNhDtNiABYVPK4799
hB9ZGJbzrh7o1ZnuWTMFNU8NIsQCeKMpwJriEG3Xv3PtvCo4gVpcwy7rhAYtZnTL
o9IKLgimq7uuDIhmxpHnO+mfaXG3IXkLWk/qcOuFo+Alaxxdvxoa5Y7nH4rqeZQG
M+9aKVYbTKKWP75rFlrk9LS74A13sqzjVY3mB2Husl4PtHYmrtjqwnbPAQeg2WIc
bupkRDz7T5U0WVGMupSOUlmCrWCJ6UbNTEW9erD8PnZBQF2erHXCM9PVP7unUvsR
zdrmnoYYO17/PuA3LtayTytKdUvtlAIDUp1nBRi7wx6Ogu2zIaXCjq7WxEhaGUFI
QTsvC5wjt3lu13I1q2uXd7D4de3f/gIAb1cwPtSw1hkzt5CKDalktE0MRv9kKTZA
OeXwbSLuRV3fP7ycnm2sq9gcRAu1a95AwUytDgDisSXp+gFtHuT0InpF3275teS5
1RHWFNnlCTWAih8V0qHKwSE757B95tMOCaAVP7iQRY4dmNsnMD3wQMaUHoXSu2q9
xhRLop/SfOU7EaXihsEvkkRTOc3kqjdL8MEbZ6pBX0vCmRzyfDuwA9RmHvyyeG5B
mZHlcmsSkS5+hn3A/R4DZb5MuOUUDZbDTqOVQpiMFMi/WRlLZOOnPus/+pYLoWfB
g7RrzOYcjYOIkVXnIWrSfCM6ZSGbJV8BfamCFhu8u0sXAvA8y2r4xo3IvPurh5yC
48blVdT8OBb4ue4jZfvWFPerRHcWwhFIWb6rKI0olEJX1cqN8h7lKgVvxAl9eD9r
1mXbBwpMJx10Dpws/6dstO6zt8DY/EwFWg8OPDUTa+m5qvhiPaKueEDpfI7G0xon
SWwBeSA+roTkyufUrHjQVOPNVEmjxRyWsQKzJwZAd4K2Ore/lFUO1SPbuUVjXw8W
KdCfIX7sGeLlyi5ZZ8vJD7aw7TiYgEs0xxt+J8QOq/8Cr9iTd2a9/yMQxDDMbeFE
nd6pL0Eh4dxj8Woqlk0B1CQUDVbDo2yF5bvQn87Am4o46TaFlqQrVZInm7zgtZYy
ZRO6tye3diJkbQ8+rakV66djvnPyuxdZCWXYlXPk7SOUeINe/9uddgqT+zth43XI
7xLdFkTAekUkVKAYcytJYSre/xgiZOAT5Cly9hC9SRcU7/0wlQtE2Cvcdocg4QFv
vfzAH15o9JG6G59l2p+EcXa/UeYVA9jZvtVSgBbq1qp+guG8D3sShDoC3iEaTJXj
Gu7ILfUvxJ0fngpR2XaDBRreju3/+HA0pbr487EwKoM2B6+7HEisqfDGtARyKciM
V0w+blGysQFrb/YVto6yCNLK5BqjcRbPFXMiLNRD9KmxJHTYvQzgc88aNFRwzJ0s
H7wIGosZTDOoFPoNYPE0AsIJQHhjgh2K99vdwmwv6i4+S1YQhxk4zUzeWSnFrqpp
`protect END_PROTECTED
