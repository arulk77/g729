`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBggREjjPfLfhe03YKvBcbbXmrxm2OIQRxzDt5EDi0Lx
xvohHiTV5MqwVsWR4w0oyrOxrvZpVgvH292ooHh0OBk63AiytqnbthBnPZmMHKY6
7S6o4B3gYGzumeQ9rsj5wZPYJkqbkXEzTQHAxNQ/rcxvZon43u+phYbr/5CkR0yK
fKghmozxhwdhZU4Nrv1eFx1tzg4qYzgVk1LdDRM3GjKTYWwNpl5aXqsVjJgf4a0o
n7rcoo7kQ5EulwFB1gvN2Q==
`protect END_PROTECTED
