`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNiBxN5VawkPxvI8lWk7tmc5lA6M9p744q8DfrsSC573
kx5lbocHBiqcLVMuAYJdOcxdxZ11Egxeaxr+Jv6PzIPIWLs6bXefwLSmlaSnugXA
iAbfpv6RdC/yzAOamndeIVVuQPUoVt/uTQoZUcRfOGNZvVRZx0kD8GUWfh0VLRqG
xcl7J1mXNegKglzxtn2DTCNND8VSboTfyhvo2MTJEVuqfZ9rAyHCcGV4Y/6Ga+yd
`protect END_PROTECTED
