`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKxTI/nmlBiTf38E3U0dICfV3DxgnhtsWDdQG7i0S6en
sptH/xMhGrhbRE3eRl3GisVBNQaBgxR+IQQeQ8SS0JXrVcUOVnlqUrSKc1kzKch1
lm1zcWsjsTtjuUSksJeVjHfQASNCT6jo2KcjhyUMucYngwGmvgN2i9W8rJHU2/hY
tamzPMXu0A8CXAvzGM1fbWyU31cAPhg2TSeBs+BpRciS2z+o5rvDrusbSEaaaP5R
RR1Oia7lnEOpQDuL5PeZYXIYNtc04bxRpU7EcJcAhDthbLEZPKWerJ0vyAnvMtoF
riAzderMbU1v465SiekE4FyD+BcILFptpGkjaYSOvLfuVXwf/amcc9PKNcPy+2vb
wH56lH2PY1kFgaZuC1+X+ZGbGcWXbBtu6o349ZVUGYCpYhofU3rRGnRO7IA8fjyr
mRz82oKwAjA+x+ruNChY9e1VgL6TKc3ArSREfjhf+RPl6VCbop9K6b5AEi9k32yX
4yMSd2Ihyx2CP7XKX2Xp4DnqVLeIxvgitP0QgW9wl9a44XaO9ajgF/K2kmLvCi2u
oE+yqLUhG/M0BL5s9jtoMdBxg/qTMfNTVIKy7g/Ja0L7kDbKAdKOj1h+kKCguacH
LWS3LVxh8jrpkrktDdlJM2zmVhdnjL279xSTHuoF7BqDI8o1tm+imuaycZ/9hGAd
bC0fdJZ96edIiGPKjJ+/pV0kLoQVBn7Bot3VLwS4oMsTtqufCoE6enuMJ6KhfBWD
s3lYR5A0dlWivZ3kehGmFwQVh9Pp2rvGtItmWLj5RX3NtiGfoFoZMT3zr/bSkBTh
cHjUtWbtYWo2Odx9qyOQmBT7R0iwnlE9ymrGS/KbPsE=
`protect END_PROTECTED
