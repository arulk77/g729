`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG/L5MSV7uFaRfCMyRyxZWK1bNhjkUCdKM0cc6nll7Qh
emZVt42gMExUC0qz0l4KtZUTd126L3gTz6T9VkagIkCYFBSB2Pd7+KIh54H43cIW
HRPnQEklqZzge43lJtMoRcYfzWOx9dkXyIlt+sLjY+GEdEA9kRjHV3khGufz9JkQ
KPpBhe3fL1QFC/a/ZhcNg5wGlkfwtg8/FkfOLEFq70Di6jlaq85cIEfpBmHY2x+P
X6Ri++94c4qdP3jKonIZdP43rwKRz/6xSEruNIK44lOQ9uphNMOyNgtbjYIB7c0f
US7uoblpzVwqFP64GJGY7UTMxcVfXSOw4blqzedMLjYAR/WNLMRMveL8jgZoe6QN
qylA2GhPQIhjAYmVB9vVtS8VUVyUlmq+q0wDIIemVT7mYkDn0mrrJpxKzjdibgQt
uIDr8ND1dW1WvMpzMGBw2dpJ18g6ZSHOr4aospabCX33k2Lh833cmIjY9QSRScNl
zZb27Eq1BJ8RxN4g4x/JvDFnb5UqS1eF8Xf14/Q0htsMy/JVEIREAdjK9X/dD29F
W/KrLfb2pG4ssV7coo/ovEd13XgO+nN9cZLrkoRY9w0fgnrSQ7drvGD2my/LBwf5
YkFbj5N88c8ZZeYo6HxyxQQlOWcRir4KY+lAOqiHeW6Icl3Z2Jj7huPjSu+UmZcX
`protect END_PROTECTED
