`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGntPy3Rn3QwMygZ/QH5rQvD/s17FlKZriQphIjHRUF4
RplkCshi8TBUxyU23jQAASE4YtEOqTVwOevNSOGZ77jF2XoEY5KS7zXK4++nyoMZ
DTBA1N/NcsWV/BBThEYSF3QlwB2XrYrMjojf/TH5XvKhluHZX4w6YLcTnxL791AU
ADDqCcVmGGHCCDzOj7S9PGPwMfAZZSWd+lMI23kWyZ7WRnHHdI1jxqjfDJqjIL4T
KesnErD6VaDs606XzUyUCA==
`protect END_PROTECTED
