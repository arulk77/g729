`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
wlkN//Scmd98V47qTC5OZktGLlxsKVRmcOO1u1RR1wa4IuW5hX7/66H3JlJE1D/n
xifLr7qbg1p4F7xN4Wat6gm2nIG2edEyZ2Sfr/CdPIuqIGaFV30Gqph2Waq5fGLK
H4efAwQB39I4jJuIcs68Cg3Jm7iPC/QI1m7p9khqCGewpsPqRg6kH6NMrTDKYwOQ
LIEyZ0HNum/SA4iEcJZXmO/6SatCyDTx2zxIcABSOEo=
`protect END_PROTECTED
