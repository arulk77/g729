`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF+NklHVm4VPtqpoztD3DdvyIUpdWiGdRUejtSvFKE1U
BwHv0VagoKvYzTJMvPOsE+YT5HnJT0K5C0KHi20k6fQkWG8uhaU+XTEzJmrSvyY4
jOTDjckDZ0k/FMxpXerEuZuaTWhuX9/apTOaQJ25/T1ODfcwwXLCI+BQbvlzB/qD
36OszKgD2GqHWXX7J4GOQysi7RQX1zhcldaj3PlnWtrAjyQS2hoQdRhZEIntPDen
nkFq/WNVsQF9e7Z6qPwizZtrltUsCNGBpiwVij6LYsnGoH9/jrGDi3ckyEWQcQE7
3kIy6XtdnjOngZJgJ/JJvshcJIDT04r5UJD9lHXUtqoj+wwHz0zH64W5jt27CJjx
3/c2zvJp9SvmGGoxUky8NsTfJo0774amObtq43apXLvrqDV5yYq+m8I6ITxQmvFi
MSmoXUlRTQvFOzFfn6gjxA==
`protect END_PROTECTED
