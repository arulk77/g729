`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIV+hfZ25Ma+fOwjkyYXeCKLaj0V6uLVDlymukRHPnAd
MxyoHnWWvuEKk/f5M2InbVKLh0gH/5vmUnaj9ShqyR1sCFeUpn8RD/RTYs/Od7uf
wsDEeRkrTQUX7d32MEvxFFVPLNvdvsyMI9SvDvvLfiYP6c/nRbIQC+74gyDe+w5q
12IWQxcvm8MJlrPU9NXGrfFEHyH9EQCOem64qdM5Gp473pO8TeoitIyR+kZq0BjN
UxoJ7Fdt2wpLqCKmPprDjI0Xe+71s1pXtY1is6vw+edM+WZyevod78eL52jWGLnd
hgc3YeirMLExyZ4bXUKFUrsQ1MiyFK2R7BFCXAnFKwCpHlUEPrxAarkWbS5te8/r
lhJH+UifwoYHa/ywD3rk6jWV/81j9QMXRdUXF18BAu9ctnmD+UlRJ9vyjDIPH9mk
7+0WHfLNSIsOmYp7hnvqTkXLqD0PTu+dPQks2ZfJCqMqRVWrwWUumTyJVA4bVI+D
MD4sJWfcUoSafImhaBvKk0eAtehIvlCtBVWTCV76TmmGIJb8p6UiRjympLKnbMAj
`protect END_PROTECTED
