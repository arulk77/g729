`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
fOYstXs7br0/ZQxRCCpUIlkX/7TDkBsNcYniMjm2BMQzLllVl4VJZKB0YRoRcYB3
/CV2yJ8NT3n9YOr5zbn4V6/v3dACs5FvbRaKlaBlJ2Gpx3uzCwM4EpS4wdr0Xm4U
5NXLRV6JqAjSlKxXDTyeCvgeG9hLKVgj5inoC/gmgkk1eKNgOLwKyhYP9SzFFMmw
FGKn098gi3mdGVJMBG4tqCMlAYY54vM5uTyze6K2izon2eK8HUZqgaOlXAs5xdV3
BIRWl+B8llRF6VLNcDhCzMS+Y2VUqbzVysWHZn2kgcc=
`protect END_PROTECTED
