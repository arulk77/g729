`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePJs6GrV5tEYY1kXyHyE1O0yye8jn7hnH6aQh227fyPl
42TfyR9Ra8vK9t8obu9LYcYmiYHmp+pJdxaJG3vwGXwFyXt5tqnRPYmeAk9FHLES
UdsvGotyU7MWZfduS8S7Nw8Bc8aL+KVj/xPCKBkFczUAh4RGebJRx77H7nLTUdPg
tUOBCfWippT4Sv8DoKePCbEYWsMdnbl0Eu4T3r+FIcc8j20IPxV1LPa57Zfp4HCj
`protect END_PROTECTED
