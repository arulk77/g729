`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAUUOQKsvieaoiIYhKZHTjFfGi0z6Kq6czYKZuc7Dk8bP
QIXxo9XUfLd35ZzEw9Dj9lCoC/RSlCMC/ZAwT6ob01oqnMWm6aTfc5Noymlfi6c7
3FnVmceFJ0IWBcYiuum0Ejqg37Uvt8asWttdMmxXQp9oUdDh8f0MuVx6mfshaTL1
c2DATtYN+3pwUGaC559J11Zw8Rc8PJ7i+OkqKn9YDBcmbQEjwmSQlMmn751kiSHV
clPw5IAyWD9mjSQI5yvAMVPZH3m7Kk0VTIO+IbvuEkoDin63MzK8TRfuPaFdSGTv
jSYaFsP78gZ8g5P/WbrjFkB+AMNJPD5yvZfhQXhYGJjpoRnCy06zxfS6H4dmEtRo
F16AXqLMAx+YXnOxWhhVr7vrhAIEDkVo3ajzyg47EhyXWNwS8oukW+tuX2wiP7nX
vDoVogjb7GomTjGTuw6ZfSmjcSx8DdBkstH0A8SDDVY5KpsnxD6+RNlz23eFRsH9
1Cf37WmgtcTiQLeKOSfm/D4p7wmFYwUjf5O3MCu6bSk7Th7HuCWR4q0BiGtdXclD
aGLfkImiYzbVjwZVP0IUsqRUb42yXSl8s2qXaHt4D1HhNXSgEfOxVg386hWF8PRM
zgqOTV0DW5mxEXBtzE2PfaNahiRh43LgClx3G0+gNSU7NUloW6xo+B62tfzJ+7Kg
0U49wUHzrIovRnaMEB3337fJKrpyTajRlV9QqfOHwW/0oFOtDKZ4BwNRbwzhhDZK
/xYYLlxy07v1vpDYTfWYzHgnakzWbcI454Y/falbuJoLPacx+/eLb+9/lmNRlzrY
TYyAnmQ66F0SbOrBw2fBt2lypTKgWfRAGwraekCYjS+afMLdSNBS95cclwKur1V7
USncnI6zSnjQP8mYeHYkNAxe8XHa/IFXXwXPTaJcRVP06rAHgeXvJKkM/CkS9ENY
0XxZvpK+Dm0nSrgFq2QGZUDJfOKFsUyUJMV2YbDexcPq6KpXCTnAIUQQE5g8SJNf
20XB8giZm4OrXBrlYGyWFJyzibv/qNkmQb/xOj99q1JwhLSwwg9rZrzVfaudTzlM
8R5ykCjhX33DHqzfIg49GngJqqZMKSDZoFZi2uY6S2UAEMuBxYJ1/Y/fwygnSNPo
8F+42mUPK6uv62jVYalmIBIZ28TEUoaiv8c1e2lGiMA8cJC2WyC7tuP0ifUwoD1a
AQHkHEfP0022JGDu8RvMWMAFlVIpPHXpV2fSfu4KRJ7Mskwxe7/Lj/RctgVKE36a
q2eFsMMp9LwM03/CxhDS/3r9p+N1oKjUg97NdYjivoEck8rtL1jlSKsNC41jzDrj
zV8TSAb8Lk8HFLELd9eEg2gkmKi5WY1MgF/jwILueBpJK1G3McuDI3Jh+fxuB7pM
ClNsctDMpugTCBYPOLh3TW7l6CY3Am3vfciOsCxhtA1HAu3vaHR6hyOZnm+a+Qu3
UK4Y7Hx7GMR6xenVFpaFPYC5V21GE5ZFQnEKYsplrO/oKgyBwfeS99Dm0Iu+jabd
k20GZZXkx+Yp9IvKU+jD+xxqbXib1QdTst62QYqbVr8fEMyX/RIHnhBXLlgFn5yH
OqiFkSvO1L+lgAwtexzwGk9rT7nII0EzrGiL1bg9QqHZy5NsImeMmLmxdMSB72tz
54ra1alCPBUAIyCRPpvsbjh9XJtsZBv0Tyr5KEXC7T/BBlFaepynCECp+vq7VDBE
Y0vebok7rvxR3j7meCtmLM4Gdq0WBCYmFzLfbQjSFDrP8eUzVYXhC5Oe31oT+hIt
bdMTZH4WYKVYMVMov2dpaxSQlVABdmdb3yEg/mrBRLZjkNQzCGn0Wo9Gjj3J3Bhl
VQqFSfMam7eqwY+goeMmdwdhREKLfWHc0p0yvarNtSyiA7q2B6zAFcnAIH2Bm6JO
8ya9fNKXlzrgbYp8+BfR0rovaMSf/cbPqVcRKW3PZRfMuwCJUdRa/4clw1tI5Md7
tzG19QVmEa92qqLcXfX0AFGHO8PoXfjoTN9R5dq3KoxBUAZYEu/0fCbO2NHl3/pH
1zGo7k38mrMyF+uLIptZgzikZhLTjj7t1BTWyE7rgL3T4Ajfqeh7z7HwROf2mrHK
iph2bBFw4zwcR1ODzzOaO0GOK4QXANz53EiVfkVAXVtf5YmW7EmVgyf0LOLVFtwJ
ArVCWb0zHbJVTsTXf35w45XhfpkcOC9R2vKlG+CfCe+MypxrQ++2BKA9atOVog84
jmpTReR2yRRIfDiYojKPPNBEcxdynWcYnGpBnylhiUpU77iv7GEfWkYI3fnuEgKI
ZDazsf0EHUcwpjeLCJ/v4sAw/LWY7vo60DCpeqajII4vOb1JuVgZYukPb+ikc2mH
58ezzTix3dBaW6uwx/ChMWiwW6uTqt3NNYrb5EhDLrpxKZoAj9+B+Z29RjIwLvAC
Bu8ZuPIuSHgUlzNBpfkre2j4Rsc2CnDYwgbzx1MI8fd2Y9UDuQ8Aux/ClUOkNSJU
trvZQOCyCmvI3xwlxAkcs2VN6aD6ldLtIson5q1oePSR/KXxvXA2E+p6nViaWmP2
o2U7aH3mlaprqNzWFOz9jJMIDwp/ydMO/oJSWaQESFCY6afBHKX27TI69Yt9/Wxd
x1gBJrFMpKTRzpYC/mv3ePt7h1lNiIss06tseLJRULAVdy9Q+5xve4897fZHVshe
zNiv3ULjewdEWuWSdX1VGwM+soeHbq8pHERSJ2QCYlohWaDlf298Ot6nz375+N+0
kfy5pdc3SMiRXD0Djqpq/0rVuWlNz3f/A8j+EK5A+HP4jjsCbiLSKe9WDInh9eh+
2VjJPZYkxX1jckR6V7Y1bA2WoxA13NthVkHT5t6/NDuUrj+XLCdli6/IQJd4bF7r
vrZKa163iuJ675hLOwdEIxQlIUSbvx6jEajgbUxmH/uvwGnogPtoCxAuFw/aQB0L
6ZUGtxqC6md7hx3LeyWSX76iuhryG6gTWJ1VFsQ5ilccgkfOjkZs+qH/EGKs/eij
4zgVi+fMmYdQKvu454xxC+Tuox4klEWEfW4KzP5cYl9O8WxdEjZZ2kxZuYEmebQG
G7AFZoSCEsZOYqcba+n9cAgYodsxAA0xAl5EDmElIYsdQayw7AFnDv8OO5/T+RAV
mCBexKaTndWNUlHnye4IX3tBRTwnOdMKCKmaW9JhLCIDxwsVyg4FB4lP6LGotVT1
92Zmvv9/hSlt3xuP48q5DM4jaGvwuh01+97QdqnDI17kqXth8V//JIq/y/Ma8LvD
uh6ISf8d/BspyJP7kzb+Yab2+ynlcGPfwgSr2EYw006jwi1T8KFf4LwpltbVV23P
DobehEPKHjltkNOO6JtaEx+HYttOopQAFCwHDmJ/HT904Aopa3UYYGmJZs3I11iv
7m24nYsUarideVdESvPbcNADMZ1Zh6XQnYg4jF27eK3juhGSU5s9uhSrg1cy6hee
pz1gnG+Ew60PIlEewkb26QgC219TWrUmy7AjJkpiLWVkT1wBNw1lyWPDzEFKXzAX
k5WyrOa319S430PZGsiWUyO88SY9E29OxsgJx7PjiHr2XByzbUk/1bbDR8DaHjn/
mVd9vPt7aDc2LRKOUT+S0VFvZdU9xcF5rg9VIjWJfp8YuGQYln2uA6/P7wAUSJyj
Glvl4ZhIQiBP2vR+6Zc9tNP+auWyOP9e1udaywPqmHBS0VAj6XOVDptTpzWqKpi9
re0xf37lRaTeDBl/YUBs9WLefUniUV2Pdr+RslnD0SeirPeLsxkehrSUw4K8gBgl
/wFeN/toUhsP6bPNoW8uae6pmQctvvLoH+K/bp0ZpamtssQ7JgkMNPyC5xsjRG/U
/Gj4hvObfIyK7RBSc1XzsO6L86HohVPek3pMxTZBV54ysIhPPccsK5IokmJ2hsDV
AUlqpx6BgcM4QArlwcNyB2yitntkz95UiANES2TGuOa/jN4lVG9GpXHKe5BcGQgV
h6F+ktFOB1gLJdD0/3OvSk+bEqu2u1WW/esVuOYapFGYZHaNQ0cy6qLLjdQgkTaA
2aDhUGr1HMOYBeu+v9BeO5ECznKKkCyxSmxNfDIEcgXFjygnbUhvn+OhZy/Ua/qD
bbn6gxCL/Jpe/m/cYsopgUdzr0Dg8CirXXwJFuoX0DdNP6tGpdimt8BhyedkkPID
2FPoF5eDf/MlH+ky2IUNeX2udX6ifyQIO4/5cmgm+TqqNmWHgTFq4ouEO7NfrG+U
SN/Ksp9kZfi1hTZjfYm/sZ48T+/nP8eTpkjLfVFirvktP6ZOhGtOFdxIWi39RnRd
pjOi/mP4PmBxiVPxctYMtbRXobEwo/OEsLs0VdhpTpVAXMW6of1PlZAhCchLqNoB
TbmDc2Oxk0xyRK/tps3/VYvDKbCPNvhxBTEXvcT4SxEbsvd/yvcQfB7ST1CjAMCt
FMJ+H6Khjzz+55yyAdJORbpIVJSZWUhoy4D9AIKofVlY7gLrr0rMK3htTPZpGm5D
aqXdif/Y5twc4GzpjFExSZK7RQOy7ybzCl24OoTNCAIe5XlNoQgpi8WpQjlWYi7+
CnJaL13iBrPq+aci/aIIKJ/AdcGvsYAzP1X6M51QIwbamFMNuPrtlowhkSlbx7XQ
MKrnc2X9+A0Fu4TslxHbmrLXEGWEy49sxyTDwMpiGDsJP1p193yMTafjmrNrSAus
i3+DiZ7OKw4+WtOVV/4Y1PfMvd8Yf+UXa8HM/aFSyta4uF7w8v0bH/R/2cet257u
t1G4Yz+/YfpjEPcSg7etMNThAYqYINOjjTbK6/24WDnEiY0vbv2CAkY2TB10JOjL
wyqKLgOBdE+/zFke+pDJ6DaNWsbyiO2OiwfjR0Wj2U/1huIhKUPsfAjVveA/5rCc
oqfBRbOboaSPvP/nomNJeNr5RD9AoxeXwZJMSrIaA9V1sTxkY7CMq8ZGWlPAG6mw
vHEaGaIXUOh240EzNT9CiUxxIIq71B4h1BZx9cFG1KK2FAsYgxqQVh3pv5uKiZZc
7imAQOglPKycxLr3Oh4Bz4B1nyOc/24cPIlTv4YneLhIoVhg560Q2ddIff6Aydik
W+B4olXhzXqRSyiTn0EOWPSw4VluFhda4y3+QJunvGv8S80j82TrVE6OLEHSVaJn
BBSRs4OAD+c6YWpVG8mT0oVEErB++gmtstRX6eBlYSfQCbLqBDYpVJjDCz9Uy0De
nHt3NIPg9DrSwnKDUZt1/8tbmzpTCWPNk2S/Z2MZOL4HKPYAUkZ5mev8gRnN/XUR
HEm5ABoOKm/s+eRR1ecSrncpFn6KRWzg7IpKWvfzac4LHi4Fng5UMvKoUt3qGtOZ
5nxJFGz9Khb10oXJ5O2AEySZTMSwpp9+kS8Glz4E5/zHCDLTUEdBlZTWj1lq2CNM
VVNTyboFY8eQxmP6W22lF2DaNpA/4tP1pEG9LyRQwkZBvEZR962JKl1L+vF8bA0e
ZOpjiRfGZG7pyJ07SAU1QOPfWjJh0nAmBPH0vekZ4yz4PaUnm6Siltowalf2IkTW
kG+s0JfaSx6zUZbqJ3F4QjYgYiC6i/ZRwO/NFLFzZHproG4+dhTv7i/euE4MBouh
2E2TvgkHidk8N3juktZvokDwkSI+ogd+0I6NYfWGFhy30gxsiu4x0s6o0BjZxJ5T
N/9Sank7TWZ6cFmM/M4unINuUSxo6uUnAFCkDBTUlOpFm0GnBS+dlvqmMyuhHdkd
j6eE4pK/GWkLF7JZxshrNKaod377jLhejPBoWjGF9OygLtRky8rH67c5CShiTi5C
0cJIzlI/FcH94/CM8w1aO3pGjJwTr+MPOtB2BhbF/C6OPF/XJxeplXXrgXNRGrgh
qUt7LiDx2VRW3bByJrbVM4ib3+iNJlIKY5Y/yhSBLFPqoDT8S2uv50D8bqges+4H
PGbcLxB61XN7DFCmk/UiqEOcEFN/HrdGN7TP/BRdgbzYrPfBzvFdosLCUBmc3Cw6
dnaYVVECzeEk4l+wk4PNiW0QwWdHd1gYR6+WyNrF4c4vmmHWzuGO3wYK8idZIyfM
XV52/ysnkBfH+VoX6r5Ww7yP0Py7EI+Fv7FwaHqWwlSclkoGADMpP/0q5VHeF7vE
RqzvIPP49YpAZre4Dfe4Ji51wVyusUfTLY8l8uVh9GJv/FZl2LHJvuvLKoa4ETtg
wMxJGyZDUfD1voWsXnftfA0uS/CEs+03mliRw/h8Jwzx7OwRrMcnrbsUAlWDRSJM
jIQhCjaOZDVcvgaKNmYihZsL8m7uqA8pRr/9MLKdVc9bLx88vbctmFS5hlLrXceK
dOzae8QHqy2FppyjtgCY8VGA71+RG5WG4p9BRCIvuQyPi9jyi570/upfKgyZGx5c
tFzrqY3a8yrV/8Qi771RyDGa3PPnrgIOVYqfOqIGbr/wPq56ronKRLfvYHqcXJm8
FR4amsucnMSqF196Sbs8657IrFSAixARomK3uVuC0j5hTHveDzYlbxSPJA/413v+
X7A28wq7guOVO6eFLGKvz2kOW5pooeTCocp0tH1NFaRhLcXuKlx8xUobUWLt+LWq
qhiuxW2RiprdRDGIj3lMyYL9a8N19giHIder3LYSpDNHsUMq/ZLCiUkq0ipL4O4n
TClzOLnKy9Dm/GTcx57Hs8vgCspn8o5vWCafm5DsBHlKLMVJcyv/ZTjItwks5twR
ShwhEjbZSdTwo1z6DQJvG1WVP1Ez2gTWl2Wi+zmj1cSJoHq4otIPay4pkUlb4ep1
S5Bc58ScX3gtbq9feaStnxaLru9hbHmCFtQ9egaDUY7fhrzoUvIHomuO1VmplLRC
l+S8FoZgCVsaXI1YhFXbJ1aYjT1nTIzKb0h/ZsRkeF2Wm9euJb7hq4Tz7d1SQ5uJ
pA0ItOQFq4bZsFtxZQqsUDkC6BVP/96/D3Kpohfpfqc0hSpk2VFbwZ2eY9bBsqjD
zGZmPuyEbwyedPiL9vFL+DFRHucb4hM8wN/f3IBKBNHpjMUpcHkeqUhWDlFqomsm
+2UGj4QMqwl8f+cFl9sTgLG+Y7OH+5aXl8X8OwYvIP1v4tGhXzhy8c+6wdSwlZW1
kC8cuq/hKjSPT/sa+6/h7f5xRvk8vLiyWCEcwR2pYQoEIWVjQ0VDiZf3XiwDqZKS
9klHxvrH0vk3lRiGTSkCNXGMzwQlXTjxgtEc0thaFueSaTaMjDjS4Ed2QJTtI7X7
dJRd6tOYVjdht00bR2a2KeUmvlZviitla7HwIHw/rdHqmVDCMsfr4IY35V/8eh4Y
kn/Y2gYuUCDMnN9ksjlbs8KRXhvj5dVUr/QkaIgpyy6EI3Mivlt5SY7xD4TXO2fI
0RvXqt4B313LylP4aNiaAK8gSBZfQE6FTE7YwiKn6O4jyACuFURvhjnTHI0SxQFB
P88MMkCWf6kDk7JeLmSHrLIGZZ21zxpcNc83FcL5ua8cKilpqorARNNwLYZ6R701
TsXjndbjWsekpevimRkcF7Fr2psPF/pWrYFKnC7y09oalMnoLCIZhb317x1pNHpi
yyEKob81QDFqfryt0kFViXR7OOhHaGILXwicwEWcmBK8utQzTrV++8KOu0IsKJX8
H43PlKNPjcCh6mPVYfqKkenkYFDpe8XMwGw54voqUsxIocSD8b5IFn3vYzZBkEFJ
XU0t2ovJCdU6UNZXvZeQUkxLjPjHdpV1eSWW+WKdmN361aNNaItFvJiokmHNByMA
4rMh3gs1Nsx94YRpzK70T7HM8g/Do3kJC12Hegfug9uetwzi+lvdmBEysnl5CBw7
c0dS39uQE8INFX24NZj5sKbQ/yXwKSYlTcBhpV/p7pMsNx1Qast0u38Z+9JAXKZQ
Ubzb79MSF0z+O2QXTQVHz99Zf+f81JxVA1cXSYbfcHfGDdC3NLq6SYGyfiDpH/CU
6gsLy83niTqbhrrxJyF6+9MqOhgEXlZcG4erX4NDVF8+PHKqlWPYfTxJKQSzpXrX
u4nVoExt9F2gQEqGwtPHQwcpfU4hfqD2UiqRHZOiJvDSYjsPs3vad0gkTZMxEG4t
iY65hJ0ROz0lh0VVgZhoA04r1jMsW7acF+WClQMtF0OUcAUpkTP6F/5DunqTJOnt
RYSngVRsQOpVMK2DainBp0TxOFMdrz9GL967CV3a2sdXEFiq6VRl6dDLPx6sOgwe
57RlaI7gnGkuJ3Vkfk5s6swaSnMyWIjl0PenfifbkBKr9Yb/YH7sEPEJ8RCgcYZS
E5manyCIOCd8g18+WK2OnUF07mG9f85Ic9ZKruTQ12W1V0+R3aQuCyTIGWn5mG+6
B4XpiSKvPPiYixf2Bngzh91LlMxI0vOYchE06+TVONMaZwRzr+J+ccTU0OMWp/gM
XkNA0A6+g46nzE9nevZZG86CFHnZ2Vjp5AZusOWdaIllCjT3wSGea9+3Mv0rs59T
TBWDDc9+R6sRjjyjZZCEPnd9MlRHaPrpFN+HKpuz/pK2NW4KcZzS7veSJrlO8Hl8
HGlWAa77ruxPjXxM/frWArMsU61ixxLLiofK3pIUpX03c/gZa4tLHoqS+OXXXVlB
RfR5SurESjZP4y65IRoe3YlVgKOf9GvuMW/WjnC6W/TlQYCvyW0myQ6qKYUjWdp8
9HygoZPk1Ys7Fwzyke7aqdqKt6+lEBQNEpzcISloAk5hdQtH2xOVxDYXUgfVNEwX
Ov7Vcye5Rl6nJWF3nHyCbl6hQCP6+mEUPVmmBOjf3UnBU6e4XQoas45nSBSP8vN+
1Kl1wZaXSUtC6lnPgfySO8NVpplf9oqdaDlu2q0wUkm3W+VLnPnkuVdRq5wsBUMy
FukzGKwFBSalgyqA0awi69Vfxfy6TiA4VVFrqfe/YG607JS2/eJ1xV6ujK2AxpBd
bGFrh96MU8k0vQTMzeqDeOhWA2tgg/zziB3Z6MZdowyT9lZQ4DA7ec64nO2xsPUI
dJvD8X6n+5JQ5o6Eh9fA1h7S3qlyvVtcewJUHQnqvj+YUdUaxIfAOeuwje8Etute
+e7lRxTll0XYjHtIpJUYu+niSHVtkltoxnZbaf9tFxX73pGdPfIWTe9Ve0oNgddp
BGJ4qRvW0o5gjaXDkDDQ9hTUFbUke2X3PHROF1NA9U2TWY3FoT7bPZLbKljw9y5i
Z/AGvEWAl/ymNTZxVLk8lcERBWRBh3yJBCKlkfNmJJpOTVJdIL7IkoivhaJqpLbT
UiSeH/p0tuVPhuIfLl6u9WUCqFjTZt24rJFOcB5ETaoPaPuLk+dgpQsq3uTLNVOQ
j2/h9bqxtchrkyQFS1W2dK+iY8RVPBvpofdAo9an3yRkYNbvD97Ki7tGi/W4ZEy1
Nm9gsn5tTqJQ+0CKrdp/sq1THQ0+SB0sSZhlNDFDQ/rErKTxAfca5V6c6tSRhzQw
73oZiroW9C/JFmaaVegE6ihg/bbT7zSrnfCnQxpwbeMoZ8f19R/AA+AqJfzPjLgJ
+7opD6EU8+2lxZcq2JqA9TcZPKhWBy0B5U4s3Dk5+W/A0pxWPgJgqO3GgBgUXmzJ
2p60k351U/YEqhy3Zwvhzi1/6EcJc8Dp63EoBVk75TWMBmzx79K+3u+/uOGk3FTc
/MNU/cR4xTbZyDDyYEkE5BMGE09udgix208JN5kztYfNwXKmz4wvOat4plPNBzjv
JJLSjJ0UEtYOVUGg8G9+6QaNQ4T+USpYgPXtsKXAL7WH0FfhpRJfeSwO1PV3+LQM
Jd78SPlonE+KFMx7psXlp5vZnQwdOEYdIy50xgO+AFRAB0U9pnvlhZN+BdDL0qrT
0fkCt2jykZPokrGY4YEx5wu067kL8rbGO3Y0Z04+sko0y818pG9+ajr30KtV8kJE
HhH7bJRtUWwD5m/gS4mWdF+QOXXIpjzM10JKxHZ0SCkywOi4xTWxIvc28fhrwPL7
X4aLm0y1zIgS4irjElTW0A/4poLUAzeIuQLgvCd1zJaKZ8WqUeqDvRCy8cbiMvEg
5Wg6+UTCH6sCKQfd9egREOL4ZI5aHQ46iSkTIszzQr6sP2EMTrlHniWMolcSCtXV
LGSx/gG1fDviOcMoQNCdZbqUVBr/ku19PALIFeIVLESwyMIN2JWKMyUU0bvERbrl
nARU7OYN113vz4KFjME3yOKQ8tmEcEcGZYiYIbqsXhLZE09hjadYfZHw5TCYOMFH
osktFzCDJC/jxX/EVH6dew3CVBC7qzKC0IBP0EXN5YIe6SGMz3+NJYeaTVycXiJd
eGGTDYwOATuPfKt/af8uj2YmQ0nchpNFfFy3r4JZzjbwaVT7sMbrq8I2kesV/rS7
Sjasurnhtjlj4OFHtqPs5TUqSn0v0ZOdkFICYhZjSedzcBCCDQ5d5tBC4Vt2T0Ti
q9SM2x1msgP4Q/3hw7DVLrXTIvTSMGz4FemaAB5w+fXoqkftiZe9/xhKkItABoMa
3e7AuPRIqvApY6RXY+o7ej0IEKAaiHev/EumDGO9aCfQQ+Gh6SzeSLb1ihefsrAL
J4jh6sfimAbOIMQKaxTnlO+vSKV9ZXtbEvAGGuqzATqVTSr0JtOofjRdKb8YiOUT
1G/TzmTNwHwXctChPuEaQ6a106ig+xIp4vuGB5E5jitU+iaYQJOnhCJ2g1CudMse
3VDB1O3I7me6yXmm4QqFInlpgdu8vNkCIxE94C7pRBcZG6SAzeZ01dZZqmOGGy5p
4Wff1fOPoGRc8G7eckOAMYvtgRohtoJwP+g1rhPTsgqqJT96M+5Av1XZEm7Dd4Lf
44W013W4A/JHqnLCVa/TcAa7Ofz72IXhFIZoVuydGndlJtG9Vbez8aN5tB/UBWTd
0GJVsTVibyWUUgZa561cZtFkuPrJ6XJ5+hY9mibIao2p31hj2LRDgJHAsUd7ai0t
6SvBrkh0wYxh2AHERcBtrSOZtvmdyFyV8OxSU1Vf5PxPW0i92MMJo2Jr5yJh5kov
Ci6dU05rupxg6yb2tdj5XpxCvP64fg47S36K19OOy8JmeP0g2xKE7pp8zViuEYn4
owgLSFMliGyiy+x8C0ysIc3CnCo+TooVilE18uTlp8tL1rYcsUJW6D8Ty3AO0TS/
88L+Rbd2TAMs0WufOJqOmOm1N3cLSWEwuuZy93eEQpABR66xmp3FjCLZRodc7RqC
hx4oI2pD9iIcgxAkOHAykN2Nrhoix2dVKABGUQNF6u9UYDLEuobZYRUkHrxmlIGL
fwIiwu+RJhxhfiGqEJDnfhYFMv1sJ6VUgfjw1S0KUd9CcRyDa0pjt2h3D6rx/ujV
FqzD8MuWyhrY2fBCSKgc3uu1mBAWQPUBUSh+88z1fBNhmf8mPIAODVuruuiojaO9
ETW2XgQlh2pZvOrroqKai6jdNGFv8gbAX7srh0y1AwJdps6eQhpbuMu/Hk932Vf+
fVkOPWLPGqil/G/udz3PbFJjnaN/Rg7RB/LYveA9Qxs2DCF+GbCpCTd2NWWbgisn
Jv3PLULyZ1m/R7lGrsg14uayeHjZO3Xc/ZqOHN1WTZAyTYNofwTLG+p55h/fc3mm
obg3SJKHFby+uDuud6gAXT0kJKtaUTajlXJPPN1Phq2jJVeLx5ilWXNGsw0GpNxl
PIIoqCXKGO/lDcD+yXdJL0J2WGxvrZvHTmwXvd09PMwD68xeeaSwgCo02hWdVoWz
okJfN/J3Fh3qAfnDsZnz8cZoADX20XhP56P7JT4j7lYEz6EOsqS/4x6C369QzZyX
6/SibiqdbTwQeQLa6C4/0n6idObm6JKwRCPgvVyE6utzDB/YPs6qLVHk57JeJfFr
jBlBzAnG0J6D3p6UXad8N2s/Mg5wOsbN+MBY5+ScNn4z+OnsLTkHHqTt5DYR2IJ+
EbvEM44QRFtrHYYA6S4spbN4f8xjbkifqwqpImc3ZjhIzc5nzCZ8UcxQzVMSMzFk
f7zOtdk9aDpejs+gT4h7p1/84oD+l10MYQRB1U1bOC5QBf6sx/3nbKbkFLS866xR
Bh9VFY+qhKW8alxBLstCmPTJnrD0eeI25uo+EQEmXkq5E77FJ0q+kwD1WrYmxyJw
jTCc4hmswtI69X6z5yuU+gikhm56y1Wrsb3On1SnRiquuje4G6uqmhmFyIxpZDV/
QzbXqyL0iAhhOqD3wH/4OJpM1LXi3rzaS89cCCqi42nR/1YXQzTDJf7ggr0TkTNK
yGbpFvzlOdjeJ61/mEAH0M60LUw0IYFQ9vyfw8TeeAGL8S4Ph/HMkE07gvJU86rI
HNROXVhnvVSnTl0JkwcVHZDk55M9ZgNKJQ6xL3xRvwZE3755C7FZTXi3KI/0bGAe
s/ROOOELTqb02MmudI3NDkVEgIiyYiyuedMq8YlS6DeP/Fb776mstLC5A/UBiNEy
qKjqu85KFnLrDWCf8rZwQVyaGYoLVAdL5mIuO1sMXlStk4MDcuApeiTfYyENEUxX
yLai2q8Bpr4nF/pKYUbaIGheym6dmQgHezp4Z+ihdXsPnVflK3fLHaAuZbuKxQR3
WQoGlA0gpvKLpP1VFaQr2VLtW8jdN3FcYpKThtyyvzIPUzLPU6wWfJQdlAjzfdnG
QvCcIUL86iZYtxap2QTOScK225JNTe9E8/H3DFhIqqRBZBtCEZAEEhCeUe/H9vKr
/6ye0y/4RET2F12/efl0gMXiVKIzNrUESnVBmBR34rAtMLU/zlnuRkFPVG1pxGXz
hUNkmfVGyLRczAjl3aNjmu38Sk4P65DE00H4Wa6JZ+7doln7b/nn7nQZn3qs75W1
23u7rnEBJOtvnV70Y0I7sPBUXKD0fah9jtmB/7t2OspD19NQjfYck0TEYsqFt1Vs
X8z4e2WsrTXx8O6YTh3t8Sku8DUdx9RieXNq0i+uB/c32qpHc11jhCZ/3T79GnIX
qm9HFGyh+BHIpBswOhdNL1xjghbK31LhKl0btd6ssCX3YrwKJg+Wf4ftz81XTiu0
hUEijNN0zaTCDepwwR9r61AEMtcrI/12ZtHtY44brM34ft8xR+IBc7fTvYHvfDKD
+VSuwShaB8z70NWXi77vz/ydiNrO7FWwBGb+kGzgLz7sb86+S4Fzo4KehnqIyQJ8
ypLQKs1mjXHSmegzWnf8FE5sdoH9G3LYwD3ERTFHYb/hmLFW4vhdezevLHEVr+Wl
wSMfkQgu2ZzIjtNj8RCOO2/VTnUYk3Vs/HeV2oTpSVrbCUJmdwMYP1yq54cl8snC
2N5vBi1liO0syd8l55cwBpdG4ab7SMoaUA+ktyjbgZADGZDq0o6frlvptth9lIdY
K3y1FB7/1V43H7lAwitoGu4nfRs0fSqSsnQ2S1Fm19a5oes7GpYUthYW5U5Dc7yu
l3OoDBgb6TWbO8aVBQRwglvDFDV9zmNzUocjuGXygIBIohApcL01hhT1OhRIhh22
PIJRt6ZyQ7VYVPsuaoWuws+jvFBPbgivjQ2f+iJq2CRhyM1inA6J+Bew+sQCiW2f
ZowWOz0SjhE+1IXsb1CTbrS+SULY0knlpeRG92QGGZyY2iiSouGNsEtIykm4oXwO
ME9jHpqlBae6Xw+zz7xnPom5PEQrHT9MmN4W+jGX8DcJqSqOUDpZwMcEuDQODYdC
e1lIzBoZE1lHkl0oAr7CYWmUA2VPd+GW9gAkZL8QmieVmTtOl+1PlzHh0GlrE/fc
eJHfzsTf67jg6HBiXdwkF/6CkYsZZnj7dR+VO4QODwPU7ALMEkledvwBswpAeOkj
yoPYD4PfQuxq3k7V2DVeJWNwFteVkm2XbKwZdCy19JdrXhX+nVtj3O/m/LLrx2vo
zeoVxuluLd0PC2eh7ImfCS6hPjQaOdQz68VTfp66Q17/QN8An8rhLGA6g+Ofphax
5i02tL+jM6D2FFWrul7s4/sXdY7rEoP1p3U6OtmYJ5gXbApLcH1qyw5XNfVRdhaN
X5PcXl0TLSXNR22yVRVzWsXumM/68njkXgo975MPAKewOtzyZpteEAshqUdhnf1E
jLYtipJ/ANFcsz8fsaEun0H3bVQRvg4vVTGOfR8HOCzxC1vlzQ8zZSam5UrPfWMN
nYt0R1SHPszO9uJThpJF7J1DfgGaqVZawDh9ShW8+juTMj/JTUtYzKVM4dfUfmUC
yVwYsBEOY7E4q4qwnlLXAxdI2wVYO5SQZV3xpr2rk0t0OsikHTPJ1rTbn+vxV9Rv
+Fxzru9p5TBVGYhVSnRhUhQKaAT/93GtUWuQO47neo5H4bN4sP5CUdh/vn80Q9Sp
4mImmMdiHHq/a/hEe3kpkCG97GMqV4dLKAXwze96l6FNVtwFnk+flNiGOtbVHG/q
xQ/5baKkHxmhzbbzlIUKwDPYe56ldjdKCHyhhtNPFafsgwHTg3eAffWZ+MYDtSXv
9R2+BHSDWbJNbampqGWYa00U3HdXxYsPUKskY+bTOL3NoFmRESCo0qHDWUMkJU+X
TAX1qLDaEZoe0o9zsHgn6itgiPKFGpLJ+ndSsAs1RDvfB9V6Ez1Az3y7O79/c4xB
uDDd1/VEJoAGn1Dti0M3Hw8q4vADFyh8urQxMvBMGwfFvj7j2akb++PJkqWCj3jg
vM/8sfWTlAOm3/+fS1bfFXyowhgbqMHCFNANq0Oh0nNhuZsiCcfYWCPPOkafCVhr
J46RT2Q+zlRckFv/BJEz2fBJPkBGQPTgyCsov8VtG4nMwPEs1CimlzeEBfHe/fvV
jkci5xzZ6HoehrzzWhzwB5PqOlIT8BkbH1aMUm4raafu6wOkfTi1R41hIxIAwmHu
ChtkxgRtaGzNdX/JValnzIr1fREqnJPLth7HoFS5pey3zkXVBPxrX+GMb2TIWK7N
iMhzOCzex7H7Y0KQqcPR8IYe/dCnA0hi/+IEEaZhtwbjflTeKBNTpZoYuf0Rcelt
o2RSA5wH3DLNAJ63lwfD7MouG6aQi/w9qW0QLttrQEkPHpTvtr43oNtUSx7BDehg
JQFwRxN08ON980OaCVlL8ENhZ1Wbn8Z93sarInaAYcuS105sJ6+AJICfl1vvZ1Kb
HiTg006U4YCm8R4xkSorAAuFyms4By7Z87gg9gFOCcWkkOwsmRa/Ajs15qKhKi/T
9QUdz5bWzCR0D5cpBYxk+0klEB7qsmGIEtxMz1b4AS4VrOPasIHo4maBRdj5THE9
hNj+XmCezGQsq8dOydzysghJw/PDcaBD4lESLcttxwEclG9Wr3XYo7ABgvF6nrS1
wwraL6ZsWJX1Tg1OYI+2GXlBDm8xUQrvEcAGjtvQinOU6p2KAstIma3DzO6BHk2D
D58QI7twEigASe/efwyUbfED9vZC8EqFCydtljPrM48hAV/snf/wjLokP2NenV1w
knHCravHRv8Wlo4uswfhzhQIJPgSXuSG2g7ctm/8PmVKDHYepaiSEp2rgDEd3I/k
h3jNUwSItD4S+TOqtIyCOG+Psv5DmUvKYr+GdRDr3fD9dc3wdUdu0xeJ6ajYAQQr
IvVe4kUeOnf0jI+htlOSGApfmjlcnkhu9iQYNqVslk9LqUejMifqi9Mpd6XUI8aB
HkePXKwg5Amf4nE7mprVhy8mn0533864ixcmPD9JHmvj2b3KWRaGUom7o3+qnlFQ
FtAWokXUxRJgVpbjntST4/kHESnrXrgX88+JFn0YLrOQH+fIuGn9G8ArpoG9m5BS
NzBlIe8DcI7/0jZ8ODL6lwoGDfEAkxC3gbwepu4NYGQA9Unj81bREu7cJ7mzg+tB
tvTb+NN3iEv8WotTl1YJsAYUHgJYHkJz/BVKm9GJHdMSajQQIrLgLbvtaKdckSrq
LuWJ56WgWMN+mjlz3lyswnjrGKdNyIDermpH3fkX/x5r4l79aZ9QeOXGQhMmpZuB
96X8x/fJa+yVOQSv0m36lGvltc5kkpaCDrgj2yXaYZeaF8AP2k43YxXY9U7IoVze
1Ed4CUU0pR0phcU1X/2M2Rtf314HBTQZgWMkTyj+92m9y+Jn2NmUmLfOxnsUiibN
YUlKUQcv0pjQtnO+cVrSpc0Sw1C4TE3BtrycXHyCNr0DdqTwCtEGvQ4Di6bCoT0T
iQLixvzFSQ20dSWrJMRHIWgVCSN3tehF0O7xJ/y0suXqHeSjBCrrhYJRJuJrOZgv
sUa5NrRRuR+OP8HKYNoXH72C8DFMGRAy2lfWHVgAhEwt8O38EJyMQa9OMBSiXsCV
EqgjnbqGn2Cc6XiUz0ATucErmg3vz7NgiySJ3XACOYx5QQgVJJFpaJAC/KCKvC5U
hCX21g1nQsam+hf46v6u3D59YKHG3zytGfdiWd/fDCUfoYquiaPw6qGNZDcKqCfP
rj6JgpaOBd70e0BStfGhyDhJsINI7kdPji3Zb37fRMg1q5Nyf1TbO72jMLuwyxH8
Y0fneAuTZGXr6Gu4+NkEy7xtyj3nEUKyJR4ux1a+rPSp1zUoIyKrJ5k73z3VlcLm
eUDZi2Us/nJbRFmjlIjHfZtnyN5MFMtFN+Wo7yS6b31TxLX7WDEhLUPm32GZt9gE
X8AUUPhEsdXv5/ad6RrTbCokhaZ8vUu+6KE89kEqJrpkQpAB3FtH42BF7y+k8nT5
61+qcLiZA5gCd8grjsGkT7inC0ckW3cKmndh1UdFNpog3Fgu4ShyzWxVUueQn4kU
qkVFzMbg/W7KCXg+MvHVRJweuELbXuXyu5pAAgGlC5bYdM+jWpdyiCraLw3trvbc
gR20OM2pVzQiznUzpleOKVWaHRSsRXIbDdn5PeQMfx6xxAvIlW+6AgacHaFhbQSf
4geyH7Q4hGoQEyrlyN1OIY/UTyZpD/Pqu3tHWKwLsZwPBKvjtsjrGa2V61riFPUN
nG6DUD/LxqWMUTkiUqJ9s/oMXknr236vMpsSGn6v50SDwd1Ig2YvoKGRUr4f4hZa
AFW3Xp4Erw2RxGPOm9tT6B5Y0VxgZQ6pvKOD3xqWN7Ve4thnh7vGbi8Ca9lsd/zm
M+6ogyjDNAxxiNnip2oQocBADvzat2hkTCF/eydwLWIkLyVNLgM2ayw9sb0NYd5a
Hk8pxa6xS8gMaCjbCUc40P2zlt6KQ+CMtPe2Rhp95HB1/F4J+DWDx7PjCVW+n0Hs
e9+XaG8tQ4BDBBihM9MSk4l70uTwEUc1fznCTXSZHQ5XfPTpNJtBQiehrtG6u36+
xekwK6rJA5VZA/JyJ9Y4mcvKh0sBnFREO8upVQcEywAtNvO6Fm0+QHhPzN4iyaIi
EpVwxjSR6vKMwmseJe0xgrNPTs9su56TtuzG1UYJM4g592nX3D6V43oG8/S5N7JI
Ac7+A0tSL7TD8a0QC+bIC2Ldg/0PvPnbb0RJ6CH4+Se4mR1sMgIQUfxIWQip4khD
4w146qgJbxrywnoMyh2W540AxYutsCIQHjfL6BGfWLFtQWQfMap/6uiYPARi+CW/
BwvMXG/J3akrA01Uk7QHVvou8jLGPMd4UslXiPqoMYzHrDnMNIL+Er6k+QZbA1Y7
n7y4WAImXQaOb2lUD06vyaQsDPFVdGd/QxSm9p5wvohONNX+LtP/KgjJNXHv/M4Q
gmAtpeyo6Hw1CjOWMyxleCGwvn99t2p39fltYVnfvkCHWJxaHjglGje4Wu7baSar
5Lfhrhp2JTTtmg0fo1JuDTf4PHppPqxUl8m2sFkZRl1myMsDmo9IrAFqiK03yRoU
RMNw8b/LTVm2i1BAMSmyUzw9m/5BXqTu2DRewURoX5kFjWalghnO1SEhiqiqqjNU
P/BBEPxwFpKeiTOiGeNVBfFFADZOdRp7/t6P3DeHqmvGjA3Vu5cpnylOodlBOWVt
fZS5efT86Gn77PYBM+uRxRdXleRny3y8UCwEnPiSjnlqz/UajcEWWh4zLU4lkIAe
kW50A2UjBUO0Ke5tsrfeX7B+EOFFmiiayQMyAggk4+MFm21w9ewXkPPsgCaoI8FF
7pncUaaSrw3wrSKCm3dygWa9omENQEXhSoFQjN6JAimefqRd2k/rSsX9oRamYTb3
cNr86fkQ3v3rg5d3zfX5h1YYrQ2qqQNLDaK7kaTo15IUFmbjXlKbdVMZZsdH1CJ1
kxK6if1qZRL1HjuB3cQHLlV6eWPfqHCHpyiWa7XgAjxk5l1n6E7vezojlNIq8kfT
5jKWTpdVTcGV/8PovXiQLLth22aDdbaozgf8cf7vErniSmPHBnR+19eyCz8mCXE5
uj4SXCSgWyP3zuj1uE/Ug/mkXdED7HC9tr9iJ0Qdg7IumehrsC9uZ2MicVwCWZP9
aIaAQ2swVvvvWFp64atWPkeFI5lHmN2YgA+XiGDb8QaIFeftJnZZkTPFjbGITGho
x14ifvW+BxeylPAUnJSQtyWEEz2q9r9UujBVn1dOV+oD2ko7UQCSugWW5GFGBBtW
Dz/J3phGhDJEe9H3yXDVo0kTxdy1FqNJg7asAB3wo6Tfhb9V2DBG+hRFXh5swTtq
6cqcKy1ZlAwjr6TRLsenrdEbcWhFaRdIv+K2kSHIwGXugEiYY4lo2OqVsemdtMJd
Fjj+tZ22gXqTbsFtVMf14BJqLYIwnjR4necAE6YsiEKY7JPStv2qL+eL6Vaa1V3r
7aYynoX907UlR/fiN4OzFpcAOLO29Z6A/sDqFcqTmrlveQSpd3qS1B7qORlDfeQO
dvM2Wgv7oyOO6gBUbCoOGg28cemq1Oa4UIBFxmEufHbe5izEaZcSihQAzduz83Vl
PEozL7QIbfAu90FePYzIn2NhBUCqqLv/x7OovNV9Mm80CGszIETOmFgVbBw5rq78
fEM/H9WQP60or3KVa8skviN0r6RoFMUdr4uvAe9J6Ih0tJYUOq5thvf9a3EzrA6c
dHAxB9+tukij7OKawZGMSRhyHsNKAFHFletvGKOWsUhruoN9pirdUjDlKh9hA+7E
CyJuyTtE/bm3ZY1AMEIowB9dDbjpyvnA3tMqL5aMCSY7q0pmnCUHSeBIGaqaklLs
xivmkpS6cifO3rDRFPk5iM22sbsYCKSIQLRNSFyl9fvl1nVhTcllb4JU60MBQsXT
fGQuon0H0WpLxvqUNB189qw29eAedSh+0aE+dpbPRXCkZQG/gHfop8qeF5AkaHGr
Q67eezIFMUSkLPB8iuwaIi0C6lxZ7TkuO9FYdx9puDedUgHA7FbptaLgiKfBJMPc
LLRegDg75jB0blKNlabRoBA3DyM4GU+fcm0WLOk1AGkHnEfM6YSMkhzoTDe/bpS3
YH+va1/ls2t4v/noijoSQjBdtyph2FHQ6XbV4lWMCpizm7m7v4AvHaByPD17cl/L
i8eMqxI6PkMycshRc8tkr9PftgBF/NxuoCLKt2/p8ESCwgoa7ZaBKIhFjHv+dL2z
QtREfdjyy6xtT2aI15rBC7EL6LUhV9pT6QpgJF77mcle4LcmJb7MLyvnOreB7sQB
RyMe8BV2RDEDiC3b7iLPk7PDrRgvpvGGJbDBsHmh5G6JPRVBI/nILSbksyMpSQVN
cQxnMLbqHCnPETryJLK8+GYLqjqDsI6XDfbBM1pPF5aSk4TYhwSdsILZrM7AQt7g
8HFC46O1qIUnMd+D8wgrah/cReP7kxOtucDUGyckeXvTHCFSK2N21172EqCD7gXm
ZPNe+lJ+yZI6yh9TYAumQgzVCsCA1nZ5lJKgybdlqwZry3Wzr8uKDdD1H8RAe/bv
6lze6jI64daWiMmpQAAg1UNWVChz20Pr/ejf0LiCZf+aIj3JLCEG6vRGgl6yq5t6
UerqzzOmahh+/1u4DLKN4QPZAbYvfHJTInQlbHRykjNnWtj2nvjERozXQ01DGkDf
3JhlHS39TEC33+EyZ7YmWh/V1sN9J6dmOv1QZ4tRxdovDtqZTRpcqK6SEU89OSrD
QF9biXtYOouyNjya0iWYLVmeakt6XfmeCIeHEzrS1WhSO908GK+RpHO55nveh9Sa
L9YZRks+ZOAWM2Pvaj2suW5hC8mWIRpeoHXMsuDJNZIIBnAoCByZkrQEMvELgFU9
rQSwB+YGK/0LkBuHH2nirRmP1t1Cix917okf5jv6X5bAa47UBx1PLM5XWkv6+LaK
RVbKK8lEplsTSQiFx57pIYL3XPfZBj9RFglr7VFYjzJRQVP+7uJDABvaoL4lks2p
sDw9ST3D2UXk9wVL7msAxbuYFE6eADy9c8BxbwpXIe/8A83kHvTCfTlpVUAsoANl
EPCbuZj3DAvs1JYKVCFRRzDvmouX+ZMNkBLsJfVSDBAQN+1GHhihdw5Yz+eIWld0
BzpB+JXtDdwUfhXg9ctO6ykszXpzbDBPqHe3v/WZXcq4tBhDSrAPQyzkNsLh9Fgm
3JsXHXA5mzD1e6iuso3HjGJGdxdnnfZx9gEzFMkXCd3zFSGaSKRfw58WBRGX20c1
o208uPKvIMHiN1BjMsDxZbr4vbZLv3kk+lGVZVBdsT2GD1URh+M93aRwgQR5WLz6
y3iUtKlbB2xh9kanH06nYOXrp0nXXE7VHOspXcWj4Try8n+aUnmlX1G7wFSkJhkA
GR32xDnKSFyx7r/uOcVGV6u42RO1pVRm8Y9cVqqC3+bMgIZvLh7XvG9R9rNBxSDv
ew9SPoxXebtONCN9G6z10Uwax7vJVuCSt/VNtSLEfje1Eb2/K22/0WjJz2j4B3Ih
sKKdH1ymdArdMG7N/nRh8OfgFsnDtazCFVqx5cjHWdxIXTSbucWbDLqHa10msrII
rdX9HXu+SwAHxTD7+9jBSaqncpznUUe5CYxzSCERkSaFr9/zI7xD7hgZ/CEcN3Mi
38dsrviGaTgTVfd0r16CihWHY6tz0HOaSIeP+HbCxFu2bBcdGKDg2pAF8pKk4Imd
noUF6J0CS7JuFDq2s4W2BBkKr4yCfJd6SWO4Ett1QAUyozNIVbxOcCg5LURqb3Uz
yCNx4xdEa+pDmeHrugrm5zT9k74rQtOIleDBuSGaapi5ndnn9ErLfYvurM+/XxBB
bErYY31L5QXt27ZwBV911tZPRAzVRhK4phsRCh5WHnSk/9K+8wq4CLdQ6Kb64C3f
FwYytVfhRIR1Q9niBlAj2/FQBPDH1YHqDjBHsIyThTfiF7DuWQiKrVVpV3B13NtJ
PIVgxu7/6r/aGGMGaIf3CSQspzaltbf0KKKw+uJGVODF7CPte3SOx2sv4Gx/p890
25GfwdhxhzdzQPaP8Qc8K2fTuy3ywplo5UhXqo0H0cAMuYFsOuKx8+gclivoq0ti
1ouVvm4srTeiRA2Zaj7MM9cmishBC2xJkiIsTBGi4REPeZ7oatmQpE8PQGdYruBA
0GnTjMUTbdC8B/Rg6d9GJlpB2P9zLshiG5PGVh9OGAXwDUwpXJsMeG3jg8nh2Wn2
R6szYm5kY9qimCUbuU5OHHzmf6dUdM9+spNFSSC13Ok7zIBlztrQ28lw5L9FABNu
Epj/tuX99viR3hdWfWTcrZuA2DF2hrN2dMr0PG2OZ5reL9wX0nBwN4a8eORjxzS0
pyShuXrGRumKiaeixbTiP2DGHu9LFjK2Bl3TrvRZlzyyPU6hgN90jf6nZOD4E//R
2PQBNgtxuHXUXjN9oQpbusLv9ldyqJhwxvBOl1Wu3CHj2IsGLsRfk4m5GiawPmrk
5ij3U5RJGeV8t+0GXrwb1Mk7F/z/azEd+WOR50FlXgOvMZgPY3zFBS9XHPQdpP2N
VSCott6esN7sQXQzUvUP0Z68c40LsOL4xFQSJC2zaQFXnXR+UlimE6f2lTdenq6U
cyDrNQIvW1yd8ObbLadG3Qjqb/ro0Xit3rp58IUFBwkre79U5feh1/wZ4nQzPNHt
YuZNFIQW3DrkYxKBuaBlN8RKDy6Mn7DKpeoYJtBITznWAQqpAhWLpY6po1gDlFh7
u3PcivoMMAVkenaQGaBzPML6nLptMQRDTmXzZT8srbPHrN6iQ+NuPh7aYrpBxAWp
Oet2wOT3QVugXJPsLu62FSidKxI7XLeXHWbbgy5hcCXQ+nQqI9gqXkxEzJKeLtYV
ntN8bhh3jZZX1mVPx/1+DTToPqilijx4/1iuEGKxuZmTllLbHCPf4DucsvSz2eDx
th5Ydsi6suZfIg4xVgLpXQKp5aNQjO1Pd/+76rj+DPnT7zpI1NhMxllGRpAsc/nd
0mkpQv7DKJ93EDXpy9vlahzXCOuZISeRnCR/ZdY0vD5OHAVj17o90KkTfOzM+oUk
EVvtkj68QW2WHikEOQVGC6vbD5ozXDePyXhBtAiPAknwHGgBA3TzNAR+QZ4clHR1
AMy9y4qBa67pfiZCCEhmENRCkSrYDjTM5NwAUup8UXwL0nfAHUQJw4TmNPi3rHmZ
LyyU/4k+qZZsUAx2JApqL+94AgyaemLSdYmEY0nJzvG7FZgslG4Ejr9I5bk1NCWr
wkpjigIkN6RXkLMKfR8QXFHWvWVbrwFqlW64RBnII6IuqhfmWFOm6yJYIqJ9HGoQ
tJLjcBOzaBgtlZcFxJbnpHL9yz1TqFG/DDIp7DePbps2yt3eRd8Zov2q4lQCtDjc
GrW/+hzpy81g/IA9dhtaNG6HSi2Wq1Aw/lcWvBFuJe9WzUJzNaP/BeiuhlYjRnaL
BiacytCYb3nyHr2pu3F5sPpR1lw1CiDwv/Niky975dewrXPmtfcMejIMGiVoHFeP
va5/1w5QwmxSo2PdGhM5sXXStQ1MuXbNDuT3KYl/hvc1VRbFuNab4Bx+NGrhuwbo
VbqccKWtL7wTXcW+sGB3r/p3yIoCsnkqh7SX5BMuVgUxB3rGu8Rg4PEu/QZ3G9xb
BgmHsmOC2Z2gVOKRVRCrmD8uJA4g8sYNdDZnkMVSUN69niw+mjTzkHt2/5lpteWy
GDtACktmGSue83I0r2Ps6aeS/FfMqB8NxLqMrHTiiw2uSWT9BDaf7FYhixIrMsaX
HplX1+dRZ+W8WPzDf6tJjQ2/dxgJIscv7hv8lyXfFdUBx49GSND5Eggcd7iuYOYQ
qyimWFmClN5fqMt2iFnmfIVzevtyicptVgxndxXYJQY2vWAcj3JG0qKabOxUdbvn
vgAeluZCOpY3oRAxL/Qe5m4WCf+LMIl7Lb9q5pHBxr9z/CrNubkSDozwgVEAY2M+
r9UdqA+i0kDezy8P29nmR4j/muxO2zmbFNwiLQSc++KtKZ0ZKSX5N5bwnDa1lzBi
GVudCQOLu6Fp4QfN0F/pVBTOopYEoQlrU5aHbLiYqphCzFCo7vk3In3UMv+SPgl2
0jIsdKvbl/zr2k++5ivMZPxFGmRnIa2qwtg8rpAioUJqjHuugOJBAAXelqRlygHq
Wl0O2GRR0mS2VA+4+WAuhRU3sXzsJoqmLThJCUGA7b/qjJKO31Cgc93Vh5a2ftEz
E7aHOgSihTPsVyOA3VsgVEHoTOSOd81yZrEtgnuxNugqM123STWgKt5Q2iVs75Gq
9OtdOIJB/v4htLX08b159ReJG20ug4SehRjXNFZwUJoBCHlpED2p9/4hyFWP0YL3
p9ZmYlw8muZ2Jx4mKpFphOCMJFX8P6hL4O5TppF0QkxAGkhnfVD/SXGig4pz4kJD
6ZrngXHDwC9mTOdIuf09v+nzQKy3KJKofJ9hVowLRa8lNuoJFetfeFOcNFZpI1tV
px0QYk+2gFIA+6KIxqKB6IsCtTtgYQddajp/AHaJq8qNEq6vy8LnLp5DKSkuLwQN
hcrfoz58ZGeKMV4Mw94aS5HP8Abyj5UUfCtgQGDj1CpvEYeomSFfnWJOBZGzF86Y
IeIbIhKfXDRennVTeCLiHxomw4Z+BldGoA8YckD1C4/Z/EY0TTiiZNxW6VPteqHU
rHm3uLHUBsO8hl2/BJxRZQ3gbr2GpOkpctm8cr/coNlv77WpfQStQHOOXsmKiWyC
Oz2fX/qi5nrBo62prWZTCJiDSKu86wzvr0kybtHce6sG79cwMqzmE/2TnQS3uikC
r5MVq0L8XPlKs6g+ya7UBd4sswVtPHkEQngGjIBaJ+u5BrTjtnCYQ13tNzBLNJV1
sB/dEcX2sacZnSsO/W/HVbWJhmT5x9UBX57LA7vnWsThuIoKTXG+p84orBjqizOW
a/IeAmrSAZhKS3n+8SsTxs0msNqFHEoFJNGctvRZIzKFLblZENdmoccQKZ9Txp9A
uN5RlyobXXjW3Oh1p28hd0Ja7kUJjAr5UyjUdGfHjeaFIh+AjROIryYrMnKK0kKS
4ivUkOFIwmK9KGLktBN1sBpNta5If5Kbc3vRlZ6e6Onl/tBQ2RfBf+55ucRthrEx
k4IEZ6cxaNTBiNFY1EoGOpPGbeS+xiPeEu8Pp6x/VNbGpB6zyDGmom4H0Rs/hTng
PGHbuJf1K6YoxNcHaopZ+gR198wqiEbOxF24if6hQsxNhpcZwuE4nubvRPnBujTI
FC22u5keLBzCZGuF+vIIUpOFy6gq6U80v+Z5ntuz/HgSM0sNt+6Uo2RXPQczdxaf
fMf6G9zDFDK4Hsps/EdbjqsDdLAoUM/WfWPf1B7053b7c69J2TtvEgqxaif3tp0J
H8y30yI8TdYHQJnnRoYhaIVmGLZPE04o4NC/ViAPIvJViQjpsM+iKJTSU6b7WGMC
iN1mUjNJBicqXzgt2MeROtPshJYMa/wrP7sCB0y2D6+AZcXVvXgGd83TGeHjEXG2
OS9RSVnKuHTKc1izxYApqccL36xc/A8R4h4KixnYE158kMCsnzZldktbVKvtFvBY
osr8wayX+kAHc1u+mL91bh+RZS2V/q8rI1/CV+nmKbEqtEliD8ZtHQlLEEeALQPm
N7ur8DJaAuHuI26UDCZmgsRZR4a2Hae3Po9tpHFabVIMB1O9MTXrZB4gCJsY96y0
EC47WIyRAuzmYTSTHtoNLcKHsyjx/v1T94nSTJNV3SX6IaxVjzTM2JhgycW7VL75
tCttPZUVQ1QMfn8Eh4H3wCFdIYuvDzxZt6/hahilbJPwdclbKC+17V19mRN1WU4K
XwrFf9k7UpsOYB9MjlrcqESKBk0IZ6+1AEXcrMQ5+3sl4AxsD6lDi7rmondqzc0f
weaCEgZYdXieNCr7s9qXPm4Xba4xTzjlggdeLD//wwtJ51RMy53V7szO3DXrcEro
ee4jo98XJcgc4d9JDNeHOjxBXva8Jz67H3ChemV87is3mCi4VzOJAkJiAM3tZhsu
J7hz/KA040Tk/fLkmIBz26Xw7RQRChADTQLS5bMcQlzya5N8AhPH7RB/qzcAH+VS
by32Y3w/ojdFJiw/jGIF7Ch38+KI6B1aS7wRdY0DXcK0XTVwrGMLodJMExtvkP8e
B0wmbV3n4/Sv97XjfPSegOxscODjHu155KmsoAtRuMJ1pt1IhwfMfc5+bwRYf+hC
/l4x0J2LHFkRPL1MdjEnERgVaSf38GHeJpFNfGDJobITLhwwqeArObsVOOj4KyH7
k4CE/ZCCdf652sSCwo5EngAjahBiLp/wIQNneK6UXaqgtzxPh53KCs0x4ssdmqIg
nVQ+zKyOGVX5r9HesHmqFMAF7iDVLrwEJHavYrbRZXFQBLD1qHrNUB6wUPGfUnbD
8Gu5VpfCjoORlafx6Cl3vwL0vl8vSnUmT6EXf2NEs30ugCDb3+1mX8OoLFn4NQ0D
YLyM7y+rwPTq0PMkeUDivU3yLxwZ9HXmc0Y9y42oS6NpgrLo5gc/LQPMX8wMAIft
7q3GJKnWvvR7YFQBl4/lleOj6EoumD2I/I2IXbc7ilFpgxU1kIFqiLj6uuuki6Su
cXH5/EihhrAHFZvJ9PWJCnKxk/e+Nhc5eaGzyn/ekc6xlEZaw6qujdbMlSoWf/zo
ukXs1C0funomBXYJHhf01++PuxuzgSKqiwnHhULRO7DFlsXqWCxzVQft40EZC9P+
+llAjeosUViUXkNE/5B63pSMtm752A/ya7QbXpT1dGDX2t2QrTh5bgpg1xwW59DO
GbTTcXtTWB92ucJlW/cMBkHaYktH9/JfvYC6AS9lcut67Kln95yBNulSKHZ/Of7J
7x2x32SDSztH9puRbILJCT3/3ax3MCVWFuHOXE1UidM7UgikSZ/j22m250oS2KXc
jyNuS06lVFJm++mN+TQaYGJEkaZnFsxLMc843rFLfvakjFX82kqcvxRNHDStQob4
DYPiuLiv+hOEDkSvVeRF0cU5KUXU6G1E+VT1MX9z9mr6X5yK/6JJTGdcOszAz34Z
mSLJhxNjWzPDRwozOG3cri4rZFPcbes7LWuG4WHvpvsda291lS85Jvd6DvAiMNDX
A8YCrhdPy3rzRIKPLtw0aVmRI0rr/dGtxl3XbCHQQuqZ+NRiM+ZoIUA31J42Rz1h
n4lTzB1huodlDK6yWYe0XKuEZqNbGpL6QH6hzv9fV1vuMAsMel49aURc+WPH/N7C
uiVCDpfpQGMZKtbZ1RB0aJhcX1lD3qBlkgPIzK2OfDLJTEmPjfnymdWnSbTWPLqV
4AA5P+5thsUVSL1ZJxIkSAeQn7UhGJNtjS0lXsLOztFML5JYMW2BzUY6Y/L9sdS5
QfodWkZSGANfm7NHy7nklMhXJ38s1bbznYuLEEwEt7XRu62P8a9sKjYEBiB4cMGy
CIcFtyaap9tRcobaQymJTDgsjjlYQr6C2n5dIvF6Yv5eQtoKj7ltDJVOvKnpI+mh
2WCwaveM8y8x9nyrAjM88Rjrc3qjqDRU54tNTTp45T2zBrxJp8JgUIOrMQzHIuBL
awYBKTJD2x8dEde4vqWksXQl10j2a8iOcF4AiRSC5ZEwLskF57/teTQyHsUqibe0
eEPx8zJs6eYrLHtkB5C4AC0XS3l6tLTsFXYzBwmuS+piIkNnwE3scz3Lm2O3OO4U
3wlkDMCSyFLfEdQ++Wylu6bOKa/wZPeuCHhJ84lYJZ67qL1wMYmj2zSaSFdG6e6E
HmL5vS93Rbvcp0tQ5HjeNDsRZc3/xib4A2VEXQ/Bq08hTXL2UO2mLf0SQg1sy3Zx
TT+IoZPWRX7/m8McvbeHPtAb1LlPKe4eGTdYXMd86CMf8excMhGsDHrOqRsZsjgU
krVE32cGPuQGFhtLEXsTiudj2jtpI5tPc1tS8iSr9A/ZhPUNdrkNKwc/2/8EB0qo
Ryo3VN8DEcO1+87TSE9mM8iEVHO/4rtIZQjHVMJlyC4X6thilHjsZHOG+YFP0K1r
CJMpQxZ8jBJ7hB0B03FY3/wrOeH4JY0WoOSX8UMLXiwu1zN9emhHAY8HQBNdC/HV
Hvy4nu2wwLd79OIDgr1c9aROzdA/wAO/an3klPxWKf1lgyAJ4yHYfFZZQvenJDCF
QIrTwqMSgHsE/CMbN9B0ycAuW7kfrupKTY013MvtFW5LlodvtJ9YHEt7M1On0sAT
HurgshPleNMQ2Ww3A3VQNFqao/PpAv852S3EOzBw03TLVSK2URhGzQ0Qx/pBMiCA
BvuVPBkRU83ZXrBzX4qNeSHhX4D078em8XeNmUXDK2Js/FLxDj7EDnZSWqkAaGtc
wNCIDv7+qZfOIhGrYT4K65QK917/ugg0FYPgIb2mVwjqA3YtWwzkXOFeC+8+LKpQ
/x0EybsfOygyKKpfZ+tTIbm6dPAbd66WrFkYAnSj9/3GzH8QQrHHkUQGnTL81jEh
WZuiSt5fUngWA9osD8+Pb81GKSmv7ZAuRufc3wXK3MkPn6NMI1o0jrhYtQzS1DON
5+WyIxXqc6TcnFl82bWJyns0i5nDOpQxpTcwo5jt/uEixzixMnuW1I46N6EjH1/Q
+p4EF7l6tY0c3quAQYLNC1WfXhWSNKd27UXTYPTfc9pGf6DO4Ox5wexR/JboYOme
XYvutshR9AqgShSHwo/hB3ybWYJqR1/bEi49KeRI94kzUP2PcPiKcgodB57bmFxU
UDegxfPNyQIIYaZNvj2mNCMHRYE/eNqyDWiXx2jRpxEOiiX0ZMqtzVo9kyMJv2ON
JIrbKdBGJRCHEVUdzen0GAdW2BBNnv9N1XEUVygfQIlzY2dproHsmYpFv6yzukaf
IFWi2gG+mCUQzudOp/8ib7aCIOHZOP5Or5nk2Q2iw7IkcfZLUMN1NRaWfwnYzW/v
2ADwPKGzII47IK1ZHbnAHkX2mfUtiZNFIjIHc9EtUBSulP5fgCA3yFxNcsV9gs0c
bpkhAaKVhsgygsCRPLjtyoJuJy99IM3nxHuV50GgPzwAObKg8eBdVQpIl4677pkk
k/XeLq6W8aMjLYWdELRpAQWVVxirwgGGA6+yp5cuyKm/JlKrte+Bjnqy/08oOwog
UMD/Ak5cKsy0CBYyvXv0Nuy6VWEIPO9nVkR7xMRhkt8eAfjfaEWKXDk/8vMDkwKa
t5pgJOOQ/5EMW0W+gXIh0A4U+oFhTr1NvyUiNoJ0F5ewtwaJeH6da0NDKDt5U01K
MqQ3k+vrSkxFpg4rC3FXN8WwP6XVKgEiumZm5Xpa9KOavLv1wP84yTVBDQM4hT2a
swsanf6DLqVDd7meLbHyRd1Q0jZv6PcPV64lXTJPRa8nz1RlVcvb0/3ruUG6D3QK
c0OlF+wtx3e6BTzD4KtqsrO/MROr5bOEPAakqLAcvbcYEfh7T1ssRV5fB3hQqOSo
Sk90JDKxi6/YV5cskB6EZ+SVStxlLgvBO3GsyN9gazRLK+UpNh8I3U8//1FAeIFX
xj34494MXm7fz9QaW3XijIgVWetWaVGb+yREsu1WP/K7wN6wSWRN7eT7bSRCQnc4
hsn+fGOiOzxnkx8EBAXd2bJEBLWX37PoEvgI860LMnmpC5jnIF3J6Oad4b1yf4gf
4fw4l6AX7TttQoAE7tyut3W0u2rRmO+VFBiwJzYElTlXTtJZtmJmsESicB3WUvl6
yBc+FdGYSCIfsWxG4bQhbu+/MG4lI+jVGwPH6HEDaFh84g+jnvtrShtrr32g2wgj
eW9GHTV0oN6bYEcnuk1X9+QAfRFWYQkSkRt8iBnFD4wMprSRMbqzaBElEl5/MPPP
c7T1Qdl6S0os8o6MXVxpVnEHy6mgNRkJERnhsjLPdj1CH1EKv3wmvP8/rlCkLXTZ
lI6VUnMNLQcc8sXQtQVUF6qqVDNda3B3TAxGn00pcGcZx0RDTgovpkF1t2CFowYf
1urekZb+DabyUik0w5pPw24gsrqru3LKcUAm2uMWC537cNxk4FKIZpT/ZhW0CMGx
x4WL8SwKrU/bOy3XYGBMNt9ene2WVk6fwOBLMDajoDX9fKAuF46BCMuosnELuv1Q
KYchE68uAjbaEsrhsVhrtIXGcBU2+DfPbDk4r243DKaZcACxNWsrKe22ZMGfNhD+
a4w2uPZUNRWFp5TGatij5hAfpK0aprixd5Y8hru2rgCCUv5vVJRS/OZvIlCfe2Eu
e7gN0NA27xIbGNWn+Ccrw3QYrvO45uAE6ba9SGAI7K5CEJb7UrkHp6RqVnVYKO1Y
d6UMPOxh1Z9imk10CN4J7+8ukcJ8gqCE/tx1Qe3KSqOmPigGbptXYNWHEzoQuIWi
BNOUm2ZbaXg4V81ulXMflgobkOXWs3w7IPN7Np+4cowcsyESIpOzCzvBDaTh6dJ9
nnyLYSES4Xd/iAnmyS/g+QJZwS3oGTfE/WqGr67vRTTVdTFPqatavSTCn4/SfWYT
7TjdjMRLmG8Ptf8F61Txe4NGrPXRmvtikKziJMUxLdZB39RbzSxNHKVEwhMwEhSp
L6bCUItXWRs6HmW11PXNmQa7ll1O0LZDl0MOasjVGR2hhSlyGXy4dGQcy34HuSPs
gEDG0KKRtk+03g90bQENSUrNzIvfWXVg8NoiM0H35IV1F7w1Xck47bm5N3oYSARl
ivEyenVNpUMc3LWOH3b4mlfetf5IPy/RqBUr5od99CZg6Mw9kEkZgFQwzz1bnkmk
UpgKWjAHhycL0yGUjGDZ7JfMdFgN6wz3jzgvgFt96/IEZ8Z/HdTK8KHwbAcDT8tQ
jWLWC4I/yoJcLXj0CCR3WMh7V/+04EUHkBk9O8ExChxYVZA4yVQLqr4f8s/JMjNm
m/0m5Q81XJh4zwEio9p/Xkcgelku76ir4/8H1UApkKUYStwAJkEWvW7biLIoluj1
yquNaAxAjf0D+TFp5QXfksvVhcfppCdDGm/hVfa4H+jF5hmkZrsLxmck9wE6C10x
ia0DgNFlZ/giwrpQHXiBqu6uK1wYLJk8M0qJogzSsluzEd647N/McxmoLQLJEQaQ
+SYeRYD8Qpceg788mmzlkd0bL0AXuLKyewq7deqM5iO5s8fP7Nivcg/p0odmPhyZ
GDNIgcAcQy3BvmOZlA1DolCz5neDvmJC02z8alrZ8OFEpT64QAtNbbRApeIfnvmt
5SxAjpzCqpDWph9lNSgTB3d/iWNEUbQ0xrezHLc9mWJGf61+eKsXhQaXeTHj0jVZ
T9IuiCqVy6YQTfgHpTQ5vdCQU+deFp5YtBWGWGsmPb1+2Vaj2AWAjMH17ZNdxsJ8
NC+jRDBwIjXYD4h/NANZ1BS9/Nwx99nIMtOHCwr5aLvMz6Rxw6/Mic2X0tjRwX/k
yogmutZcX6RtBGRxEQS/zIRthAzFYUX73NyctE16Fqy3TypuL5a2Z1E2V09dcH1s
hfnTUU9PFu4we+uDsp5vOj4+FhwV0PzyFR0LXL9a766wDaRpps4GEuJpNiJ3/y1r
Xl73OBEZajDqpumfoj+yoGM2G4pTlt2tIPyItVMzdVAXLixYGdlLCLvFpNr+3YrC
KFMapBFkmlbjKaTj1h57SvbUMkvMf1q3RqM9W4TsoC1O0a2EoPzUV/SCSGD4Lcsr
5IexGjaKluwSZqh5hg14XN0c45Qq6qa8H0/rxrl1M5qaCZCThl8krD1F//GPF0Ao
T+67qwXIOvXC+dsAnEt9coa5k2EHdhpIFCS1rUXGN+Q1kN6AHcn9bGbDnVgh+6Nk
d0H0jKtzY/SjoeGi7gdN/4vUy0cr+qxWQLMPSLtp+dhRQOE6u/isat+JHiH/LWjw
B2Eh9ec9WCi9pIxaCgkSFLSMxcm2E4rJ3M0psEoKPuEfnmbJmkvbjmhuHg2MB/Lo
SEvc2OvG3tFyLVWuIiuDgWglUquUuUPOAfWtGTOIvWmmoqpPFFoa19C1V/HOKE4Z
wNugnl/eExsLUboXFtJjE3B1dcIHDSJtsR4RUX3z18npyRpsalux9VTUZ6RpzLT3
dnVLD43at5rOwGLrSRva7aZag6PPxTeHvYwxglj6yoFLCKkhQTAWR0MjbUk2Rcru
lGk9h11tTI8LSF/QxoK4My1I6Bnk7aKCG+h8yr4ha+zMwRdnXnqob151mTvqQ5Cx
Rby1HWjW8M6sNio1WkSPCTRomGfzfJID3AAaNDK3gF1nUVQpKLl+EIhmzHQ1cyYC
d5NO41FWs28QP99lS2ty43KfbrplJvdcqzHbgV+c0PpbK38q82HwK3SPlIsQGu31
SLH6Wy2PzWrwEc4WQeledLg6Ex6eNDTrGKm1SwDul3mFiMLJyo8HrNDU48MGRpfX
eDxXp30VP4Yq2JEjxS07ZdyCqGbKQ4nr/XbzR2Q7PwxbQJ6ZIPSjFByVQ3jCCjiB
L8Jl+y/GsX5N0nXK/hp46Q2vfn/KDmitDtb+hJ+3yFyjSLGG+sTYtOvEjSnv9bCg
DX8d5TQ6Wx1VE0Btum/iOy6VEJ01cnrkn6j23c53zaUx+KNkxF/QOI0ftJBKESkR
aHmtKx5agd1ndFISRmZCrgz2BwkpZ2K8vt2e1fry5Wm5aahbig6wrpe46wnbnrYF
KZrKdynS/lfY016WZgK1lR9CsHKeLAbEW9Tk+WW5FLDsnqOzCd9BsXpzl0tNeI0b
2oI0FsaUNAqTMwR8srrtTFZJ8bbEEVaBCHpoibPedU+Q1zon193IMWHNzfmp2asO
nAXYVQDRkofbC3Mn+x95Zr8wb8sC2V7onHVzdWwbUsPTOfEmEvVHR5cuPwdx1klK
1kYklbBEva/6QxX7xFjJOXNDimt6AGZBjLDkSmMgXnQjlD3c7IpAHk8MM9GormI3
RIIm2r+aFXbGa4jFSPb8Mn/2WAmjWr0xhIXB0mnriMgYTmB0pDuBEYSWUcIs/0Mr
1tuHnnK9LC8FnxktwG3wS9B9aHBzulaQ8lnMjMmyeuxrZYEqYlkfwM2JRXHnMcqT
x15Mtgjjp8mwk14E5rNlm+BlDl8E5t+De436xtm0ozGb2BO887bzN/r3GK1Apg4I
7U2XtvmFFk/IUkAldtbtyS7mVLb0qRO9y5rTuiUOr6LYA0ODheFIrhcwjy8auX2Q
4i/EbJdib+tgqlI2lKvzox4/dTnGvD+e0ha2amncnqADvzPmoCjvuKRgT+sr/ZW5
FQo9UZ0XOsPtxda/0SKorVKDY5RtgWMOZMFcMuBPYQJjTSSdU2lD37BaYXWiP/ms
yI33nvzpxiPe9oPr3EJof7aIoW9X0bqN/FRhL/N4b3bA1q/WzxXWzSRYGwp0Q5Hg
f4CN1DoynQSwRFfBtXd9USFb+fNsVlk0nFbLLa66ODqjVd/4wr5f78toquoItdqZ
FzXXwMg9wD8h8jwL2PJ/IvqIYUKGu3GOyLf+cPrSxKCopuHPysjhTRR99PV/i1FX
cuKX8a5I12VKDlX4EhJjMv2y0SobWzGfyCnfDRM9Z7Li4Kh/JGW+2JdsrEOZ9Ymz
rNZPGlrhWcjL3bTYPcm5lgQFQmuqS8NSCGW1FuifElVBfHiJRVFuV/TdXYVEvMq5
WlYvjrCh1GoFkzryhX+iJPvnJLM6JAtdtgS6+fufStesRKmENLVpuB8+/vL3DpH8
qkLXcvyNwrVl3LYrh0mmL7Yf5UXsUR9opNr0KDWZtHC1KHAjxzhe3hsnTf4wivs8
BY2uYEn/35bvk2I87DRCHwdOjvoFivRjCyb96dZvDuj6jXyv/nNAZLb+iph0aeEu
PwJhH2qmLieUqkIf4FffbVq4nLHoY95POVZDWtVgmBNs3y9oB+qwYZO1u2RNkHms
3FN/PvMGLiSjQVqObR27q7hR3kPZ9+Nh8ZXWnY6Z1XQu2vpVKNNN2dMmS7pz1fVs
xL3KzZYxd4hG007jQsfhfI1+9V4sacPRAtJ2YXqog2PcPYdbLOn7kWXUIyVDoHpW
G2FrASVMHamyL6fNl8Akoz2tqqZhlI24xwvzBtzgP7DyH5z7Xm/QAekbBCd9mouY
xLb0sGAbZ7Z7sVlGYzUVSf+5aONIbMKhhJkvV+bsaWfMjAM3+TYsTffQs9OxBSHz
3y3BvWUidzhYAYRDhqiTMacQ0yTk891KkeTZJWjM/CV92SaVMebWwlmtjwCD8Pih
8yBXV+wWh4zrZ4UXVAV+rWRw+/UtceBPYBquNF/wHMzkxb5ppRnHFFgAleNuv63d
Tj3j2z0jfbeml5oqMP97JBJayk6UEScgj0HThL8ld0oMlvZB8GGp6p9y2z56Xw/P
ZadxQoZODutPkCNkPuvk7GEVvCL2AhXbQW6A/g5e1LR0xrYdS3lYjtrlgJ9HkWRP
+E4tvR2RlB6rTCn4RWs6S+dJuobdr9VikqvQIGp0YYHli4L7ci1z3gBcBm3J7UyQ
DRWage2rIUeKLsvSzTV6U8T7JI2jzMgDGUc//WvFYHrvASAH+urQzFwW9GFFKtbb
0wudWFGXqN+ZTZfsA0EMDldfwoeKqJywIqmKxZqMjFf3vKJO6cG8ydLS9Gr0TioM
/BZ4WZBnCPFwadDW9+xfFeVR0yP4BV9hAQSc47xrMzn1uL9jd6MgtSAn9l0oufgs
9ui+sXfDiX6HdWxrgf5RJxeI+pYlDloBcy9erhTqja7Y9dzmQdnUNUp4Mu4s5JIA
dFl+Zodw4jblAPP9G4v7lCyLPs7QgQ0gSLbzmDLc1V7poaoGqO61dFZvAflB1FNP
60I7su/4tVwz53JROXANlal0i/H/1PII/8Sj2PYpgsa29VUnmv2a5ojZKIsj/hR0
qrUO1nGzoI3WH31RveDoGeAns8KuxKnlfLBUiXqPcylCT1U7hjPkCXHb/mtqktWM
3dRi16vZlJuwA6KIHvxLRm4Sz7ml/AvZihsxiLVG6Gvb240y97gyqi5/dIeZ0oP5
yONWnlqYlw7HPH8d1wWNdUMQXqn/HtXkwV9bjVGoMeapS77O2JJNUBEi+juinkuR
6rohIBjz0JHPPqRlDk7R9eqKDGLrfGSKNIUY+jIa/ePw2aDbkpOTov0d6GkIBQSl
v3iu3KtBaGpltFXWu5N6xlmllt3HDYk1UekuV4b4i7j3htGFsLSK20HMOCE4jzZm
zNiAYfMdkoEi6SpvsM4oC98YqMgWgXGybxX45IgMp14L4XBL5XcuHzhxNHiATJmA
4uIudazylOzFtFe/mOy+8TeIl2mvbZcJEF3h+UKptc1isfSCkaoVaa73jPkm5hkJ
NrTZ//AmJWe/2HPBKknUHn+Uw4i5wMmMMXQJ7YJ5aQaaHXRwSoTWToZIgAGhkTbm
RZ7FzqrmzoPxglcjgVNn6MPGnDP71rt1qbtrer2JLw7+HT7ka+cTAHOt+pjXK2f0
8IAwmXqyoy22lN4B1rQK43R+m8exrWS7MDHhEM+cERKSkg76xZ9WaHwHEF1DL3hD
Myu+NIkmZVH8ApTYhiSgWjv4HBtud/wayMjUG+OjLgtw+yTzDbLGL3BAFuC5DZH2
qEaL3ygVZDJ6d7RfTY1ePPunLQ5wHHC3lR6udhalI7t81zNibowKCohkKceV4PG2
yUDCxO7Sf8eb7ECPJfJkKEmqFZwa1kqJO5vtzaJXrFvLYN0YLUnbCZ8FKp0HGfH4
sioI0DP/vDIwJS/Eqx5zNfwKsqblBg32EQVjhH6GA3FyY7Zjf5OA3CiXP9kHT539
vstjTA78Nz5J4Bsm+MZIpuiu7MldYb31CAzDmAZH4kmnsYVrNxSNTuPtG6unlAdI
XsdNHokJLIftUYIp1Jqhzw3WKdUsGGGKtXuz2U27jP/sr/4lBHL+7/7gdlb/5V+j
M4fh35uuJhZYX9xlo8WIYbMzJAtG+2HilK3tC3yZEwMbHTG9oshR6IXTOFZy1Z1Z
Svd6HqgHNBwWzDhbo446p/dB3keUyMQJluysIL1Lz3lq2BrdhRouK0p94gRwbljd
aGV7Qph5kzugt03a5WGgy4FGGZb3Qrlna1qvPtvXfy0HMkImu8wHXm3usp8awBQI
qbpRROKgOAPGA3vK+WOp0XIMCEvjHXHeb3jRQ9rNfMGxtjVnomBzkKBlje2kz/Ln
Heh1BBYhQiJbCY2a8SOpuWANCHfmaZgR0idykT3RbnW3uktohjWKkfquYlYORVZx
aEnk2eYahxISkLngOL9pOLCcuWapwFgq4qCma9ewB/K6M9b8Zt3IsJQtDS6cJ5p0
p1cMKXUY+QvOtsj8s7uVuW4wf7GP+5/HUXCvLTJnEfn4YTaNktPPIfVCKJsGtdT4
e1+DuhRGJhLKVSLnI3OuPt+rtZ8TYnzeX61vOeqHd2DdLCCAOje9IlxgyHhtZol3
rk/P65ps25BDSitfv1Duzw3/qUmCEifZRBw5jZ1S+j5DVASDlFhiEtN21/fB+LCc
4u05q5ROVey8FRTaTquWg0s09sLTOOlX8dlnBguTBiln5KM+lQFxSw16iIwzk2DE
Z0LGmYpmbfNwZgSDcPgM00BdwJJKchR2IZEIM6eVSiU4mVtTZwKpOXUx6CUobZXC
9hS5BQHKunU1MNOOe4FUOHLKZ9ngRpj4GILfz2XCxnMjgGFPrnyjPFFlM7XaNAn2
PMrg77Z+p4njQZFqnKZr5HawNBzq2XvLpRuKUVTTun+9yTGqwjdClFsOZuq1jHGP
JkV2CB/EVrHIqrSVofCIq0Me8Ff21loHULM0+R9WK3BKNWiGF3GnvoNQzCB++pI1
cTGJCIHIFDTQKpr4aEq+arJkCnTZaEnHYwBHikEWqx3JtFud+g9YkEjrCLu96xTp
nIYdlvtgqUxXHe7P76NbAS6GNjFUGlZ6nY6HgURhcK/8CdB5rU2udllwNB+rQOIJ
DcWNIqK8eXrPx66cuzVK63pbQh8SAz020MiWLvbpkbjoL9RD6siA/H2AZ1+HEqla
H65c9EU00hKDjTiEaYABKJvH5SiAHTxRfeKQd0vpvyhX/zxT2Fy2u91FFCdfDS2O
fk9LiTMrpK92Bp+6oGNkkd6E2WH/KvrxPg7c0zk9kH6IZoaopNxd2d3Y1iYconzl
4i+dMUB96WhSoUo7OeJssD5jCFBJUQd4Y7SClTZxA1rAb//OmhxgT+hyMcwL6CA4
eqzCuJnTh3RRUFiHGig0tsoXhloxTvmHk+XHEb1MEb2B8TeqBcO320Xk5Lckp4Al
k5wS8nwmcd/t8JRQyDSXQgjG7bvM4lYdCGE49qfkaZQ/Vvix5PJBpGQWNYq5d4va
Opg6sIk556xvdLC6OeAEzYawvbw2E9JRYfS0kGI9noriLnIxZilYMHlL6IkU94Jz
Zqui7x/qVqBkaZ/TjF8922hpbRbYHbK6+6WQKKdyVI1e2w0vMPPPk2uXYWrqYsp3
19awXzFTBelXfnzXsPOj2vX54z8jAYKKeWls2B3vv1oYLilhNoIRWteqOPb0LmhC
1IOsSQY2jbXOZ0rbJOAjRjIFc+Bb5npOFoGNHWAOd4sekfpjmWWxT7UzA5nz9TQs
P0NVadJczj3qpYinokWSvCkpwrzRkgfzZ2kBlnmgzT4Lu5gYEOV13V9BdZGnNYYf
PD7zjTBCsNTdH/TMrwztOo9yBWbZu9Te9UTM8SIhmEx1jBmn4vcpfMscVardmJr0
EXc9ziRoMorxuynADBhl5BzFssdY1hG3+2apsccbddgq232niqLt7IANlw/4osqN
fvHvWbH7ow3n8at3EUVNBUpOfJOZLyUNrKh79PuMtyYFuWpZiWjQqlq9xP0ekDQw
y4dTSex4pyNfSdt6m6iIe3aar0MfA+PPQS8OyW1om3czpxRBBgYNbuaFeEnogdKu
lO8ss2KdRI3cqv6FfO2ggJjKv4gty5tUyX6/beMDgcvgtoxT1uFW8qra0M0sJTcx
6fwZXtSMFezXsaiis8BhZBg9hV38XjZCOvo6LqEvU+x9Wo+7/5HQ7J72n3luBHpz
Ws3RbAGRhO6cACPWbbhGU0oZQxZqdAyJVFKFNizLgGGN77C+qn1dOUiQjH0PKSlf
ayAAv94h6vxca6Q/XnO6E38I6LJggyewXRuzmOXe+dq6u7R6Xw9lXaVZN6jgGZ0I
ldsz/ls1nF+7MdHcQ+QQjlH3+3jbWjH+C/9LUmRr+U51B1Bn2HjzV4TYHkcH86gu
GB96cca2tSiEMPo2vwMaLhB6x12KHKBD+PkDLXX9wZYgce3J+DwfLDRRln3Mubaw
nldZLiy3GF+Nb/Am6qc3LM6Lel93dr7K6c/GiMkwC05c+9lQx86GkWzT5KT0d1Cz
avGNZt3ERQhs2YfzmV1tTo0pS8CGbp5an1AhrHY1hyy2mLiyIS44LFRpuO0LSviz
D/bnmqwheHd84MshzWmxUJBKrtcvl04NMwnVCvYov2JzYdvXNnlt5V2YvqTFwmG6
jABeMcwjzVEy5eWrIRuuC+bEluNzUbL1Fp2sheyzZXTISSJxt6q3Rl6gR0CVWr1e
MqlwYrCfOXZm3Ha9ojWv/nsgdqhHuLHg8lSTxC1Uz8fAdlN+HooXO8zpoAyHt9de
lP72wC4W+o62FWfqeOUhJLcFFtBZIzxIjrRIO6900lnmEJv6tjKWM1V/37cS2q9J
j9PiGqzVP9Zx18fwZqFhhXNmMUUKtne3+YdzY1RIpjWsH3OuSDI/MV+gTVF6ISNX
a0zVc2Y6NEc+H4P2XWehagabm52uoVKylO80/ZhkdHvlZbWg43K3rFaAI38iMbcj
kk/Crln73IPQtbbb62sBH+rt3oSbagNZxSUoWYD9VrB9lIvAEAhTamMCpLOh3zHe
QEf9xO0yQ+0h818tEcPjSwUtZWUo9PEg+/tgBPSAhCPixPv2rdz+Wskx+JR57E0H
1zzsHZPa5Zuunghep6dGU4xI3bCCtQ/Wq2SKHiMGaq6vG7yLFCmLKhGHlyI5bfbj
ExzJjmELFBMxhQS4o67nJO+tPq96pP6IB52pom3o9+jlaaO0Cfb19g8cSelzd8+G
MxRrIz9IpUcQtfQswkyfiyjYZFIplIwWCwVxqNKHAq9AYyrVtRcaYLGHS7zEL7rj
WxATeFXkUw34AKWZeiHinFOoltgdEl1BssSLsrQObZhXt4+hcoYeJQMdmM1zXDfs
MKWCChvtIq0tZeoFEsaRLDA/BzYJ6fh7lR8TKcRgOOI5Ewlkfy4P7xDzTZoRzA8s
qaNtBa5yYvdbkvTo8J9DNunE2Ii9ZWSO/TLOTJCLMrOiKxGEcdRF5rYeKl78etYf
yglWlYeYi/T2a/hXxMC1nFtudYBNHDrLwa6b573nuAoMppAE7UdjzkrHo8tNBmQk
QmTFEQfzRwWPTi3pVmaVE/14uvpMj4BTv1HHSqzm2DMg0oqhGmUNA1Lwxxlm/yXv
xDP6qxzb/auicXqg2Yix8fg/lmq2akQMn9BODcyJNM/uyCYl6Iw849ipNyVmtpaX
BVnTzdFRtQqp8FdVMjgxzFq6Nhq76C2IIRzkZ7qBO4+OHY+Z3ss4NgYUPMNRH/DB
prb+dPsOSHtSKUyp5U8oQJvnO4APZMCaOCG+bWKJMZOf4rr4BlXnPF6ydNvLsKbQ
Yb3l7tnfYnlfJBaQGWyspH260Y6WkPnRlA8HXgO8p/jlufzQh1MSBM+XfAfbHbcM
I/5Ks5hWniJ0tu8qFSgwQo7MEjPwpTcekmE9ie/Y8COr4lwBcZxMlWnABcBs3XE+
4OMAfdZJqcxTPCoSESXdOfo2j78SFYrV24ZCTF8K1RK4m3Q0kHmAYHxpRaVDY44w
+biMZKUrAulxKqXc2bhkGDtk7EIhMG83xXURpuhlSpOGmQKRrbZFYZZHf/tHZInh
YBwbY+jJBGUIkfWVhPkg3tYuq6GVHNhzA4M6+Cmh3O9NwWYXXHbRfsEVLm/hnpqP
e/cLdAGPsr6JcgqgoT9vgS31SJCTxKHFZKFXVKbywWkX9d04CI8do41xfpFuAlp1
1RV/QKH7CnLecO+nzuDkZDoApFjXysLq/AhzmLh+hSIqmrqtfk5ovlbShPZjPOmY
kcQMoPYj968uStkzo3LV2PKHql+U9FP4KM29zMMKNgsRcxdEluLmugc575USP9k4
RygA79rkk/hYh2pmey050ceKrfNR71TIMidMHaL9JzgjZq5pkTuZos5PFr/YfNp9
EKRp6qPSPU4VPwzS9gxHSGXhwA+vMKWcx+JNbDQ9ChhD9DoOLZvSiBIZN4MOM/Y/
Y18W14+YkLBH5Y8H6vTecUv4KbE6O0eb1UwABkkkorbXsLZqeWNqBUUD6CfNDTor
Kgmp446yzj8ZRi2Zc5EoH/PZHakquMZhmgpStlUAsBlrP18eDwIuf30vzbzwBauY
mKyS0o8WTtnWz9wLWRgew/wJJkFdh7MSPe6gl6KwAqZlSyYBfakZWZHDabrzCUXR
5izHTwHl7McGqD+DFlHcvJ7VYeshpDohwkxRreAZEXZwIDtHd2hj00VtYLgZWjiS
NcunJTPDC50gFPrwsRLCFXN3rHM2SpK8Kn80B4KTb07y9TKgOP/nWmDAMwNVKxNH
KxLgO6ovuIbaTGmz4ptpMV0KfWX5K0EDLzZqKvxKI5nuq/ktx7klmlwvhMg5XBj2
+qOvwexetMJLnW6sjBLkDrXBPlZWR44RUDayRlx/BZ4vsVprdor6BmDQMenLCmzd
gBIp9n40vO9fdpAbEXNcWDHwufTQBmTAO543D1IB3Y8YAL8a8zngRAVGsD3aU2VT
WeyJJAqT/gOoRljzkcmVVtcSRytDOBkmwmXnxN3QifNdgYfS/m8vMnGXEySainnI
j4uRHUyL4Mk+W+wT6U5iHBz8HPiU1Xhmy77Oux8jHEV6toUtAbIA6hK5Bp94SKc4
Kmaa1IOH4Uf+P/1g4j1MhgRyV7U18omCMrtzZAX39rwWwT1hf+tC2Yrs77jkTQOF
MYB9Pun25lVV4Z2Kz1+tDYdiiUKH08dZr2n0kV1BH7JKIL60CkRAnMWaYEr5UuW+
QkxFur6r/gk0ElHL16CrukbAaFTAukXIjLv/n49Wpy34R9yfHcmROXzt2jbv2h4y
xgq4r8+8hwjaMNtCWPIFlJyYbi8vIXnXrSwJquzwwf3BX3Y/uGySY6USp7pZSy9Z
2BZBsrAH7CdEVaC5cn1wb0RCI94rp/iUKCTaYpuTVtzhHXOYDOUQTSDT2WyzgQDo
MiOOeAt4a2W3RZewtrCwiE/dNevqM7x7IiCGWVHpg7si6nP5TS4DHZMbn06D3q6v
OlXNe6TpdKsgO70oxKcS+qGqaOlQeP+d9+iCMOB2pKR0ISTq8fVluBpTu4X/HB6K
E82g3Knoa53HSDw9S/NOAcRO7CFv4aXWUwkFfUqJZna3Jn9sxTCIrRzbjGp1owyD
LRrw7ebbJ5xnFWlJOEH8KDkrdLhlaahW4geV2yUZ2YhNH2r72rWzbY/GaG5FFpB0
Du7Hy0WroIyJF40m/hibAlZS97g4EolrihhoLShvAakg12ovxub+jhxdotd3C8mh
J+91/pePCf8mX+O9bUO6BIoYX5N4YcRXuBZp73i1sPTzBux58Byk7U2/gKt69Kq0
dfDiPiQaRcX0E4Cyk566BwPLF+5+Ea5evgr3Es7bIcCGgsewL1SYiUTO9mB8AOzT
ITQ8wzCjcALp81szVkIlCxvIYQZJT8VJtZASzsC/nAWypok5bYpc97MT3paU2pWk
RAX5BZkgG2JeH+3vJXqG4zZOMjTdd9T5kxhjEE/Tsv2eq+RVn5qU5pZ1P0rzAJHI
AsoKFlp5BqdiahGoeTMtO0wOHkHGBN9nIp0OeFhAcPQzTUXRwEYJkKSy534BJyRk
ABikxk1UwzZbjDfeVWRi0UBRt1pviismWKCV6cwJJTDkkeInwdUVsDkmn5FYjvOG
Jlpdt/wtTSjEzhRERT5YR5FzkIF2YS9nfI+yMyuhP5PYCU8zuyb2V0jvDgG3yRlg
pV9Nk85YXZu8YbETrk0R139ByCiq5YKO2j3HkpapUqZRNMMtSi4VJe95bNZj6CXb
spFn6Kbo0QSQCVDvcdGvc0e/7XRWu6jxdOV6g2SCkOgdcueTTp89DxrOdUYVnRzF
Gt4riXS3L/kYiHa16viW8wcA0lnIk7I+iAjvkoEEFpLi62XRSMdBnGmfcJe2I90a
MaLfwAa4cOKL3j5J/dcvBfBkh5gi3Nssjvp3MlRatSskZ/UbAxGqy9l9PMuwFMCF
LpdMVyI8SRPrFCXMkhAdPFO2XJ9u0Q5zW6/OZCL5Z6Kr94gCfeMKkVb5r7yjx+P2
Yk0Y2AzPCs6NxMH5UmjiSsjztyLaSwnM0COitvfF6Y06FFWaoYynHcVhra5n3WfL
CIf8NnHHB9dla/GFgnaKk5khhUTgIwcmOom+L2M4oI0iDXQ0g/UU5OweeeO9nD/4
2sBVcXitKuk93qEzo+tFWmmIM7PGQoQyMiFGys4jF++KfZRSff8Ce5DQ1FvB8pt9
YfSYannABVr5Fj6i6ZrVHGZTFmLy2j1i3VXPnSyB6BdlsHozGJLIwUoyId8oY8KN
1WREVb25s3ee2p/OXVy6SBPNxU5zP/H+RkD9qLNjEuvxzXphCJHFonVgY3F337UQ
IC0MEEmvf0ccfaj9E0LSbQLCJuQ8UeirHRqToUvBS4aC0JghstEnDk3RUtrBhd31
xpflGqeT2oEny2U6pCnynWYiRU9UCDzA/WvgXAoUqACyF600r+Plyam+RYpqBbuG
nLpwaLxIxMg/2+0CWt7ukGr0Rg1oSBUKm5KTPatgsu30O7lqGUE/TN+/FMPGNDKi
sjPkrPUFTYBXeucQ6Zo4lndMomil8RhL2rN1Hqy1+spYiWY9R574weSB2wwQsbsv
H4NKxPbUuYTiFEcAmX9Acrwtqn2bgqeS1zqxE+2BJgOdhuKVpcLgvs/Tb0ysAb8G
y1F6irSZaHbDQ+fOjQGLzJCpxx7kzU1qBFZegIMlfCYCX5UaPM1pxanH4LQ7ZvgV
QPL3HDnhogCxO+Y/8ps6bleuVEWAaDtGU7C9dPFMYqL5xbHbiYmR8GVWiYaSymXo
uGEn4inim5chYatxYhVfgCf+eAB7bA4cxHdNs9t8QaCB2IbCDFufgoki/4lhoVaO
4uPIjGO4bnpnKAG2U17JL4Cdp7AQnpAvdpXEY3CAUuFZ8XioN8rMVOl7/0cXyFS4
Xr/8jdWdLAKvxuLQvFOpHyWQZ92pzzmusaiRBgwu2iaZaiKqvxTRQL7xq5c2Tusd
GglPcxtOXyYXzdhOR4g5JmPMOz8ggoQeT7CGgE5KtwBS0+x3ykERL0ZPw/5A3foi
BOYtHqaXERl2kgnp+HxMxIap8b1mcdcZW4TZTjh2MReCrS384VvfwLlFnA4PPfAa
7SPLxGLZJaK+oIFYRf19sAiYP/Ss24wzKHwTxkd9n5sNIAcYlHPni4rvWZ/0zxRU
KgSCzxk4ZqjUQ8GGFijv04Kp5bUYHze0xejtNmFPAWJK3K6PDjPDaMbTZNeyrLyN
WqypX5dVgvUuoKWfztThnI05Zq5xQRtLDuhLN1LpVEcYApS3KwPfR06Wf9cBfv6X
BYW9sVC3zKhPfXR8vDU1L77K6WCFlk3v51LS/d1uGSaYJFD1N9MBK01kFJcQkToT
mhYNN/X5KSPC+gPmXbKe3O3xDfpvw5HyHEZ/VBwq59EAr7NPrGnd2TEtLL1S24bM
FX/y3aoLQr2LqcQEl9/CKFAKY8vTSxrOWIt0btlZUQBn6TphMWQ2ezKvvX9/Hfr7
fyB7XXw+3SP2jX8OT+q75b4Y/3b7QQJeen9I/zsNrzS8WVuBVp729vOlGuf3czLg
qo8lLiDojf/UkmSkRz8xUr22aFOU38Q5tJS/I5QEhCfme6mX5IMJuHmU5dXpMQCK
2zG2DlFcWs+gpHIEeB4X1H+bdBzx4oUIGeMUOugnoKue4AOxZwcB+A6K4SiOSojr
4ZSI7eKc18j/hhejWerry2SSa6N9bSLW0Yx9Y7rx5v9BeQ2VD7dxOH4pUTKnb/nJ
MRALB9LOTFE/71JHxLOFjlUw3DJdQ4odvP5aQeZpnjzmsY+C12mCGMUnSzSM5Ect
4mgpLIMX6fuYnlCjNg6OfnsRLlygNsY/RQV1s4NwD8pZQ6Lt3hZLazwUGnkXSif5
XT+X47EdQwJjH9VxUV1bZeqUIAwLf02RpfjRsr1hWuDZhHa24TT3Ev3ASkiPN/ah
/b8Hva0jqWGDer42S20yAmJHu0RK4EVSqPNWMe5cP3XpdYsMPJB2RElS6TpMFcID
DqPFbwAZX1s5oSUMLnwOPAvqo8lyyndCH1LXo2Ijw2O/DZ+oQZ6s793FLScH/ZPK
W0RfE4p3hLcuJ9uhdxB80Aka3RHGB4iGhA2T6dqDcGsgMMzjluhQ4Bf/E6c6vUqO
MPv2srO9FuprHUwp1oyP8Q8Sa8YCvx9c6Wq8/BqGs9lvNKraVEDmCVybOd2UC5Le
x4XCmJYrUUdrvQY8WqZiiBNyhnNkuR5TQGJ4ciZeB2yiOUU9tnaDE04L2WmuPWsO
Dz1gato7JN0SSxKbnFWcz7PPtUuEH6ZBEIgzgBjtKg8UPo1NW/y7bPKuA1/1Owu8
06tcj3oHV3N1QWY4M7ovcsh9AvOCrlm10kiRPxXr8X+8w7eE6yHGen/PFc4m9EiZ
E4tLoLUMrvuKrf9kCUh8Oz3HMUXFepC+ln25Xq1ElTW78duxOjXcmbENOFgVo4ZW
rNjW5cSgPZTTcnT0DOUxi4tEeM2kfVx61bttABfG27UvKvX+6kx17qou0g0bKYF9
ZAyh29ybWERK1w+APFz0FKMome0RyNLMCvJxUUIJQBVMuNeRJ7aHeCXMxxEtYum7
vcDQnuLmElDMFIEoFHUI06IH2CkKT77MGPVXOvQs1XR1u8A1PBxCrxAfxUhA5TTh
AtPZWw/FjR95SCP281KrKsBDIqBDdlv+J+c+3/oI//PLc5sfbWmF3en8+U1jZ2pa
iTaUaq0V8NsRUsG7FiDDX9IXvLfADz79fsDwrMhr37nKHwyWRFFMnq0DHnFikDJX
N7zgMFVjRP5qNSXApcR/nTi0J1ph25QFO4zgI3v2YeyZdQ1XyUKIlfC4DhafhWUr
ib0CezPwmzEISFgKssH38AYqn8OSPrCvEJQXyk+hjX4xtOSB9IjGFirxsQuJcO+K
jx9Vtanm8tCuYHXCbb8g5Y6xpUqqCmxrMJsLQyV5iwTQIZd2C4Z1bsbU2m6zRc/s
YqHQRsFqQ5TM1tStN36XuIpuENw9mZXe49HuJoaDv7VrQt3DdEsbNMerSNQXm0lr
9TxD2oRZMN4j5XBEej/1+sL2/wf4GC5HQvvH2XzXr8Zuk/e+pd/VaGADabA2HAek
j/HTqlTKLw/57qEYhRrEl6ei55BzpHM6GUkW6HDtT+D/T9ZByqFwLFGibCL1TG+w
0Oyne1dhYqgkgtARD8C+ta9RiQhOtJdRgILGlDdwiRbSSVZMAhE7AHdmVOsNA48c
vMskc3e2R7rWvvcgYBei1iWWbvVS8UPwTAmE6FvR3NrttFEW4bTXIf340I3zqYf0
1GXWxkUIc3+ySeLf2CKRLL343D3nio90bIGYDWyEMOBMXsjE4aeJsh+iZ1LFLZvc
6GOEiwOAf8Nu5EqwjwpSGLrSuCNxO5j2SnADfh4/nVBfQ61IAQupjpeIEPotwz4T
H9W2dCLkiYbNCiE33UavzF2gQOdUGNu/HFOPNjZ1grHvVCtT98lFhXU587Qb0KjC
QCT44BLiwjQeIVIclRWRr1v82pLzJ/qPESJOvTkoxU3ajyg5cqdWRFn0MORhy8MW
UNX4Iz3RjdEMLxeefu/yERD+i96re/Uqg4fY/FW+K1aQW1yWyB+OXf3p4F/7zPvo
7cMyWtRwfLVeB1SUts07dFRkI954djFWBa7nEOlgkGkZh4Lwe1tAL8maxudJuA6Y
GjpHiIn/5zOBdMlcnSP3giI95eJbWI0b1MXL1K0NQa/pvBPejAGjZFsQcfXi5RFI
60Cp+LHyr9CDGvGugxhejVjdkRckh0O5JLBsr8bdjztFhd8mm63WIJiKch9wLoe0
rZINVp97G1TpGoPJo2Vt/z5z2o8HhyU7bP5wLmcnMFZbVV3VLUVPWg/v61EkPRyT
G0TgSw4tsI4K2bH2K5sf74NK95nKR1OGCG6g4XLwaviMZFOoMeRPKA8pHk0OWhWB
sHOSuch5uf/xaVHJPMAlXE0b3Hxoa07ccbhmKmmKgrKhjfVHuO1pVe0IN4wrfazQ
qImsKFv9dJnm4JhOp1gxBagOVaZ82W9b1l8834WfRO+zz/UFZ+cWijZyhuhc08st
/iPx5PDakf3rcYnb8D8kGvtipvmR1+gpCj1l7rg/ZQ8V15dh6202414iTKsBBsuv
ohSB5QJHX6n0SLCjQ3kmza56Ozbs3/JmfW2yGWG969fXfQ2HJ7lnBywYiSFCFFFr
ukR4G2wOARSg9Ohy6+TG3r4ycxj9OOOTTcJ/Zy27ftry/sGf7IuWeES23xhJeG2N
t2BxSjghENT2KrBICiXaO0YfPUlGQMX8An+HbSU5NW91o17naRLG+An7Cdg0woVK
u3VdynZ/63hC387WJNa0MXBOrpQ/iKc1SJn8Q9xp/xaVS/HYHCGKza/83X1aRohT
Rvuc8eWPHfCaSFSsoFzzpeXvTELxblO+v43ZyEXsYoBJtInNIAVE0h0d0KBmCKQT
9lbxRGfcfO5Cip5FZE/qhtXbXmzr2QK0B/mG+NRKj9qbGDJa8P217qvHmDJRpvZF
vsxguiY3/WBmIRMsEYq4ze/IpLhPvDxkmgs88gRo/1l6i+p6FfhiRC/t6skF2Hde
4DxT4dFSlrrttO3LKzWjzT8Yn1tb2tna9eNGg/6AUg0zNu39zs257DFku3vaPsmG
bfjjSnJcAQrRIfSOjKqE/9UNOApnOX2Tcd4YGTNh46WzXlU5JsBB06emNRAGIW8o
/1upAX4Hrmjq3elQPWMumF4HBmtRyBS/dlOJe26kicqhlAdqTzZFkW/OjJSBLdYw
nUhjB6raziNoQpukOXinMXICP9vNU9lrPXNxK+Qom8R17qOZjp3DB2y/k05DpuMq
7PxEr9pm68v+lIW6excs7rDu6URPXEa4r9P+Km5wwdiPjs9lE6lSM061ELHZEwHf
AXp1vG8O8w2Nmt2sVsQQ8lkT56nSIGeBp47bW2gSnH0sduAFrM1LOHNgmFh+cuN1
N2v2/m3S824V0Wzzp0V/tL+IghakoYuR3qOImmc7rV+gCkIEs1FtqP949w9CG7Tv
43BP5CuaNZeo5qZEuT02q076/PmhSBnJ67IKr5K6xILtLvqUpde7sK/Q9lr7NBVw
VG4SuBM8GFJGExo528GeI4Ts/ivQapjBwfV8J44xjFLt1ga/HIjhNFA8u2ddPnJp
CQFNrztNWAKp5b0WEHzZn2a6BqjIf4aT5YdiQe6SLaWWo/o5Pav2faWAPeJ7dmqp
2whGieMa8yJhGdbLySU5xDJW5uBpUio1HF8jwsU6neemtOg5SwgcFu2i3US9JthW
LIDEmm8wTFcOVoWbkiA+YptEUWBx3opbmRy8YH4JG34mjuFzbzqnM21QhmXKnM3U
XqRZI7lvaEem0b4kcM3zccYlRHby0cHqgW7bO4yiEGgDT+C1Fy4bgEsWA0uIQHcm
blYMaTAEz10QnjWOd2kDfNkeeGmpZWFLD7SP2PA72ikmzIp3meLMy6qjFPI4eAke
y1iaxorOxEiM6OoupKE+bN32uNwjBu3h5+6ddq7sbgRMHwG7ypBog0rzVpAlFD3A
gL61cnDTQhLzA0VeZzw84wARR4wcPLAKG9TJen0+K6lfNsX37nPiXEAOTXUkZs/Q
kiAIatVi5Z38c7cKIojBPIrCS9ZcS2Uq2ZWzDCb3DY6Xf+oHy224umeHhOcFFaWY
PZB5CIpWwzVAw9kV0GUq+J8c4NTn4gGTA3IEREcc4XeEjzyHE/jNRRiAKSx37vyf
IPoLsnPqmFAXG3fE5cMHI2idCocdH5VcipWtI3HBcE7wrNragXR5lUcYY0CKGXP/
NlLHSx++ICQtXfzLDbF2dDsXB0DX5flGdkCu5aBRB6wuBceLsqiUZv4z6K38mN6M
/ovyepUSr2+hQdGBW/PI157JDyI/dXJcelxDP/yZv29rHKTtReiJud/Ah9c4wUkf
zlgqD6Eq7jY+yqRIGd9GuTyRw3fwvraTrf6zRgEL60PftIuLfaVtmKwxAbfVaAEJ
qGYoV+BYCdjy1zBoFabJnd2GSG+mmop9B4aDAl1mutiDmiwsXT5sBnw7XCiv8Leo
AwK9XvZ/7Dh2D5QkDzjYNG7b4DGVapAUPPkLE9FwvlCCqBqrXrgRCNXPktVap6xM
LaHUTu74M1DBJKb/iPv8W+2sBCYuRNIqK+xrVZxWZ19arvAdf5Y00Xe1vI3am2RQ
NIhte5SOY1HFbjISTGgG8Fxrw/dJT8jZsSLWGjixh+X4LNgYi/YtD+wZpbMm06Nk
YT9lwRenrmVklSbvcO16J/3Fjovrszm+4DH643W/VKUzzheFiZ1NRl0Y1lQv2Qlz
+DUU39qx0+JTECbkzsA3y+46WDbksZpwztQnpv1Axe0eIAiVaCnkQYGLOrIrZUph
fjsY2GStNNHNQreydMupdr7MhSep6pPBoY83AsEgvU6dvQb0O8gd0oBbUPz/sV3r
ZToNVdg1yLvQ4rKLp2BojjjhmYz9Yp7uchZil8lgWVV2O06lNNSCsyalla34txTw
byadNdwBARTfptAbzM8jfG3G8o+ytuLYdsLovSJDI68ntuuJ43Bbrlz5ZtpTkxC3
t/g/axUfoS29Zvz6dN92+c1cPTBCt+I/7MUVsU6xofYLYRbl1sZXK6RpJYULPcVj
IIbWhM81sWupKhdR43VRO3rLW1CkOw67zpDG5/aaSn0wZUvQ40hyonrIsJHPDPVW
1uSniJt6vzkmnshNvmBYSlCKLXYyqe7Y8Q0MLp3U+eJNSPqK4iePVWijpQ4Qz+6S
ZufqdKsZ9pUaiefZuzuTc2ZXzGAHAY5eIgWuYO7+3mbdWNv/w5kntO6ScE68ToeI
Sz0ZwtE2uJCMLymgI1aR8jkSLTvCZA50L2IQFV8/7PebFT9EEEHlydg4rqDM5ZOw
8LpbCYHm3kxoph/dLIE4MWKWv7OdwCcgDjnIAhssYz7zTZHgOh6/VIa3+tDbw9Oa
MjEwkhfaoWSB1oB9lWXQRHO7sftN2l9pccWYuD2uVOpsHh+UaleUxel6gctBun1U
u+qpJBf4FYI0O2E9rJlW0m4SlMZka42m3Reodu4OTsxO1af+Yg1U74Wi+2/ppxD1
DJJivt/QVMV4uVMsKNOHCJ8rzs+HoYRLzvL5ogxvoz6uDWEx91MITmR4cda+wWoW
2VQsYlX/jfAO1KY1O05eesep2y2v1Tuz0iG/oMxeTSz0/BFXDs8bOEbDxREWOEQU
cYkIS/TSs7/+qwGJG6JBrD/EFN16L8h7qOO7IYBy9DXQrysdLRqwPMlhqODznZG4
cB/cShTMWVpIFGFtSyU9DsC/A2kMEHbTNrAEZ9dvjFDAceB0pe7H3EOkOItu4YE5
2TkACx1fy160b4HPRP1UodIbZAcMPH4t982v3CBInWItpatel2ABtI/A3+iuyKED
eR6FnN1RR9EF3V2qxhl2zIlrYrPAtCAt7JwGihU2F876RcePvGonADJavSHQNlD/
zFpjH664nKE21ZrPzM8Mzq4djtB2SMiVMh+cqZozfrW6rsRPdBteU3IZ8AqmNNfo
L/xavwKL6PLfFGfAZGLga55w632lw1F1p9fJwavarBISpdHnNZuL9SGSd5DYay7L
sjPEi5hebVcfFoEO/6bsZe6TMSezzAMBGAk7imPG5bVSDvEjDGZV1a6l/UeuGzCG
BK+4s9kuiQXMa3QblJxjmUiFxpGYz743xOBUaahkc9WkYIKeCh8M3VOQ25kIX0eO
d8EufKy4mkYy4FMDLs0T7aviT2rDTgcRgYrwiaIrt6Yg1rlradRGXVRij1rc0o0L
yn+HFSST1nYdaCEehSLcZLPFi4eO5hHKw2Wd/O6K6PlpA2XNjhrNjl6+7F5zZL61
Sq2ojFU82S2Cyur8jXzFAp/6hwdK6avP4pu8ykpa57MsAwOVT6W2LwUbDD+f2unN
doWZcUunsbie+UIhTD6V25/PkvyX9b1oMYv8kfkSgsyM3wcXcFVdQAiXwWUMl7vh
41Lvgp2HhUDcFEkQwUYG9en8okFO80PsBEwU1JvuORdZNYRMcdlRWaRimz4ROnsN
KnNDfzoy+7ub7IAHVUmW9KsYCBNcUy/4cUMq4OsswSCsVE4J2vihgZamcsimpNtA
676Rwjju9z/Ryhlp7a3tQaP7LKNuTsSzoBEvlR9tNAD70xzfl9llSrh/m9XzcfSZ
wIC0UNKcx/xsJNNTSfIJu4KW+7ubYEa+ewBFjE02pP4NvNclTTVIc7bOPJFHWZBs
2ImxyR/6RVae1UCaviWk73y2zTbT4KZKUfgwsaXnJ/+txQw46+MEEJIjN82rXyFa
7HBYbXokIPk95RvIV1+MUnnEFtr4MFryuCaLKIbMZa8eTDLcGFGfa2a8OyppbvCC
Dt811Di8Qof66SI9znIR+0QD+ZdNpFV/rEM6+DyadPFeaILf2mcRTqu2QPH/xcqg
FxqsmUCLMvcsWArt34DKON5G0zkUMvyj52tiCHOetANpxpEjYm+ZvUVqPxvyxe6k
ZBx1VMARVis8JzLcppIdBOzAwg1fcTr3Wt5E1eLVJcHc8ZEzp3eoYjhlspp481e4
JWTA5QhhG3N/ufE9A4wZf2PqbwsSNeNvMqqhNyr2ojxJEOWbmOqmev5vxm2R6Vcf
1Qf9eyffVy9Ajpqy88/7UGCJmkvk3YQ2tzOXAbXkke//ODasvZNq+wgDQqvrisGe
G2rNrdzol0qjE0BDReeW49t0JYLNtIJp4qeb6R/ohcuAGN0BtsVTHhB/KlDsnL5O
J004M1My0N9xdxOx7MG3SzttPNRaU7JToMZcOCA+Zjnb6mc1u8oMzykT9SToeVfy
Rg/ZUtght8nSjpYfVPLOMGE9PgDCbZCQ8U2yJ+x+MLJWUzmZfXvwlN3GBM8XyQS8
A7pkjyl6BF3qnSny6XZyzYVWWj6CJAnL1bDguiVRde0avcfAZqBFdOU/NEO0LSJA
wwkI4t86ci4BMxCVkje/kxcQn/DsrZwguM0VzFS1O9fxXzlcLHJyII4P1QD/IuQj
xiy3ZBmYn4WEfGvWeb1LmH/h0z5rSbMJWR6JZAsRM24ItYOWmOA+RcofrHjAMDS7
mUTRgEYk6ioxzShcv2dcMocvxufjj7Z/vjVUAtjIlLXa7NNlVs+2j7UhOUnSgfsp
blEqSDLrpTozIsZIX8ShrKHicy77bM7+meCIfyafYh7HMwPCS3JLyGQyai1scZb7
m0sADF2dpThk5ZS+MMQ7Qf/i7W8vb1/moOjP29xzoY+24jbZ1QOhyd/f1mhXDKyZ
SXuKEFR0TwQldIwbwse9D31AfeXwQfrwO/3iwLr3PbBuPndz+M2Z0hSqcFDlYOJz
utvipXVOdyGz03Wtiq3ZSqycHTXyxPo5/PMXjEhNnTauo+bq/yRczFv8ugCBuQY7
AExBGuHgTnXjyGgeg3nbmVzxZxeqz+zOfv3zIaycYj4ytQVrjI54TdTeDdbCaoPz
bmAzloiazSWqDYg3cfMW+8MXpEQNqEkk0qJjuOTArxnREA6rqLuTuD6BkVPxDcBG
fsNUdzC+vO0T9toyfKGTV4Qh7rzMJZaAKhEIQo92F2ozCa7tNtbKv8LCzAFC2LeM
ZuePWUlESCkGRoUrwhVMPAobXrhr68h5TnhtZJZH2bzcH8LLmmIqLe5rQwlnywF1
8Yi7PISDKvBBkWVbdzTn6JZdjTYHfxhcLt7BFY3q6j8jPCcsPHLKSJEZyNMC1IU2
j23p9UBqpenuUgPiQIJWdT3ve1YfZwUuKMf/xE7ikvWb7THdq0xiW7cc06qQKAFy
wpHUDX1N8zWuNadX8Q2JEAK2VXkE2De9ZZbW0+0UzKSW9Yk89zXsFwQJwfLLRgEa
PSKvEazIAItR2F5jBlJE2PAkcCujisXC87mYeOdTBoN2sAM36qlovtMZucw9MGW5
LMq0eRcqgo62Jfk1+1gNZAUJdBXQ41Pz5e08A68qE63GaS9msAxVABLERiWJXUeA
zLvW7tUOPbni4yDpRdsbRTS2+QgkZve5xzxkZZ+2/eW6DtiHn6FqEa0u1tIc4bse
btERRebAx53KdRXpeRcNPppDw0YoI7ZSMLfnUiS7E/Dj6vOo/g1rh4bbS6CmWbP9
bGKS205mm2bFvTfSwuJOI5T+tH4OlLm/Rb0tenOIYsRCuH6/I44GYeU5SQuxM34h
D5YTxQilu4uxabOLmTKimK1vKcywS3XvW8UZwAIjr8FQF8EdMwHi0/yjoldLaHWj
i5QhAHLIyxGhxtflZ7R9EMsprsYBPWwGuuZ/FaxdDK5xEmMuvQIALcr46guYiUgb
vdMSuitNava47YTmEdSWQeT/twbC3D7JjTL51gEm1xpqp0LV6I+rIX8S+fTb+e9n
abOVXFGllY7HcIURQ1dd3p32sWUWg22XqV9PfjmkeecFeVI6glQCDLJi7qj3coKD
Oof4B24GOgClAgUIVwkbeubEz2ltI9ub2HYOHoTBZqaRIXrt+zHI9gSSVyIA/1cn
Ma1gzpY5ivRDzgYUfsiAu20JCR2T6euuGDEtmM6iSJfmd+37BOK2ib8ckp6HmYUO
nO/SnHmcHNB+Qe6RJXxacTZ/P/j/8EhnI4BRhkuamC/FgWyo5sNcl1BaE3bQjHBb
23yOozWlh5muWpMJd44zQ9K6abpU6ZjYdtVtEXOfKd5G0U7uBktRZsZS9eCTTugK
FgBCqZ9uVLk1lW04fYKMgEAk6YxQP+rx69ppUVtjPpUWsiahrONeh1C/F+YFTMJh
64cjLARw11k+kf80uC5xuhuBSgCFDNdGAYvAWR02cy35KJGsu439T5+1fyvXxlok
5Wr3xxULl0gBV3i7Ja97zl3gTaodt55uOTs0kpErgyG9JA6jhncTdfHZbghOegjg
pNOpMSrFlF2BiujyD/3aRRHgjf4AmnHOtKRWeibIkPJhdxVPL2EnCOm9A07Tq3Jn
J/+whsfBBDVvm+Ze8IpBmISR3jCNYPYzxPuvnxujDWUinffX6yoMhX9U4jQg2Znj
wB30boQ2PMP9Y6B+iPqzP/deyRpKgGmtQ+4+dYU35zFA4hhnaA/atIZJC/7DuOUi
9BPYNXl7ejQ1rHxVWmkvc4lWebBo4RcF5y3rmxURjnyXBx7FDVlIqKNgA7c0H161
0nSQCR5cbMw5MjRoS1E4W/t+NB0N3aOISCbQ2eUIyNycvPtMfDSjiakXwhB7X+vG
iMGteuR0uPg1NFhu2yxVLRU+3D321qfnMCxc8lx+sJ8JqNYrK44J7Cpac4StZe+X
Vkwo3L4T6B888tCbo77HGdvZvw7wa+EA+HUmyqTy0qlNP5DvRfeIs6zP8KsHtUzi
zPkNiPUG2xlC4xQrP2T05gy1tqSXx4T65G86B7pAj3jFmqfsEygOzCIsgL4w/dNm
JfFyC19KkF6K7IvOSnwWugkdccV6CkD5VvYtTzVBtpWTjfgGJfGK2RMYIgtWxYOD
qJtVRssI/OOnVlo+7L+XmMFS+bgPG6a5iG9Bs4i9FACma/Q66qygD6Y9JUEcZ3ZS
BcvNajcegiDdF8dQ4pqB6+PX7Dopqaq03R9HIPVKQp/0R9hT1Fmsi4334QWeOX2C
LAf/DFPFTnL9dQqC4sYTNNzJx5d44T3OCaqw8mav+ieGeNACk9uiBleRMVE/9aXz
FO3K1UvvG5axZRfeEmUIgKb82VTI5bhhrRHkp2/XAhyNeyZU6x9/zwP9kknvKfjT
aDS770/seLNoEC5anbyXAVF1XyMSDpUGCDugbN/FJuliFAjkqRTN869xoMSJPbBw
UflNl6BUhDVzBhtLuwcB4wesnNxCsCviDIgPhU7nm6L9c8Rwcfk9S8msRT0Qj/AM
y87PpBkghLhHpxNtfV7OCPIIeVbBTz9vFrjsUBwbiolL45RB9+J+HLJh8w3ARuvz
1uvcRyl6kvKEqJxsx5m/psW0cUeJ/aqQcmZR9fH5+i56s62VQTfZwreU/6ww2Z1u
4ysOwuSlu5Df2VJi+DuUEHYbM+SoNZrF1YQ7+IVnN1TSf/yrKnGHxnoKC0Oc7Vng
iwOFPhRFeND0fLoNHVGmLZQEwU90NwUazk3+NKjizXHpK5tEi9enFvqXQq8Ql86H
y8KYT9A5SGUXHuDUPmUs7keKymQOFtGy2ZS8Z4nrkksmydtW50lpq5CRb8/G4/Of
CO/R3HY6EB4EiT6tMpVVEpGoAZ1NzhsvzdZDc+j9ZjSD0MiYGmgyAb1AbBWnphu/
qGhqjrO4ZqnLL60K0wkbrOxPG+xpSV93FwG5FwA20vJGGK/X5U8gsASMbS6G3xvF
56dmzWMhin8CghPJ7f99uE8Lo7yvRy3WaZ/hDs/nZuwcWaOYWoMwgasE+8ppw2VH
uq6ieCX839qHG9GIKGRVCUIlROi8FQzTd00AZcCXMRHV+IKdxB+6/CNfg8MZQ+6w
AwIFVUEhxp+Ki1R1nS/28bmKTKelzTkfS3cjOXw9Tlu7eovX1GGMMncM++88tKzz
NcPLbdFcGruF6BOwRWoSFvCGBokgEnlbRSoC4Wgy1txfR5TixT714r4BtN6KL7lq
lT3fHw0fcov5Sm8nlucORBklBLjMqz8ZEsXzbXfDzoj7MrPYWNsz0Xie6iLgGzT8
TC7gRmeXXKWocJYrHRT7U30l9clbfLzRh1/8BIjtoViYXVglTnIfHyn1SpZu5As0
YV4ai6cyh/QIMtDWzQ/RG3R1NPqg+Zz3phD/ES/LqQdFe9xrJsBfb4PWca/4jyYU
qJCork53PR8mqB0HORI3F0oZ/lTeamB7GfF5TatzCHq6s04fO6JnOikKLuiQMomN
RV2uUytQpvzr13s8Am0kSOoaLajttlXBoi8EZeG3U3E1KxPi1/3MT8BQsznxPAni
J299+b0D9/P8foXjIm47kvoVjNvmsbOY2PghVcqLuNqnEi/fWV9CRW0QoPvsYtRi
GI5EpH/hUre01+qxl36lq0IXL10y5oQdemQNyGF5e9/FbKgEYSP/DQf+9rNxOkfv
rkaY6JiZt0/L3pr5yGgrlRp4xa5/hbmxYE/B/su7cYWPomcicqpqevwb6iKaOP9y
VVETeuIV8XaoT5lWO60ha72cQZXn8+lQXSuxPaHzwOvJ/Bsgg+W3w9Q/VcsLC1gu
h4Xf1ZpMgKyYNqPbYaqy0613VorFLCeBcHXsdYtojfBUCI4C+/syKg55KsxJBz/7
XLw1LLpCOi3F+Tz5lIln85UBewE8ptnCf6Di6D/4yuu5gPPJy8N6qz/Y1VA8GSiW
a58ozTngsfr8Iu7CXPLC+qAxxZkaaq582+IepAuhxv8Xy3zO1KAtI/d33kNaOBSO
BPkE1djJC4ApXqpojEBJQIoZPoueISfFUJI7H8ALwViyI8hizSWeU6X6V5QvOjnN
jbPqnQIvIKCkbVyY+dGvb6EyXPz5PAiW8JlsJeB163fdgf5WeA6fya9pXmvh45QL
ZguDH3CgXYRdCQbaBIrVkyjNZDtsJZ8y0Uef7ERF7UCeyl77iPuba/YLiW8H5/iX
FfWnkPxTvyEKBDC+Wz2Xzk5lMgjK32SZfdWyYgTdzvgn4igxtBkVyehrlDGI7UmX
U++7YCUSmMbiCTjoJi9sD3No8qXE1roSGsNYMRtriecq8e+XSKJNezBVzKumEdY3
iQHcucbDkC68MfP+oDv5LPEBbIqOxKKzjqlGPe0K+FZRPPlb1qRS4eGwPDsD1E5Z
GDqxdT65s8HAXUVdoPKozw==
`protect END_PROTECTED
