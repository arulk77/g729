`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJWCOrk8YF/6p5+Zi8ktOABV1d4FyXYxXMiiEtSu+V05
XGZL/rGpGsi79t0R0yJGDl9o3rW6QsISJdnfxzYEp9bwQ5TnQyu6tMgsQlKMI6cn
KcGHBdI9tZddVl5ieUMR0jdsbHIhPOVnoAbp3DhcyGv/HKm4rCZtpyl2FJIupkuf
/fdJqRidFF/b7SUZphflp51ji39wl3wZlMjunc1Y06eAdWrCmVfuyABjn3hi6oPE
VWWf3KcQ+rE5FLOJWn0ghxDVcJFB9LDZjaA1VIfDsIlNApX/ofjxqM/OIa+I9r7b
Zr8qq4ELB+Qc7uiVtHviBOsdLFegar4eyQZdyNOjOcLsGXhnJ83Nr5Z6goVO6apW
yZdgpRjOPVdVAs1EqYfN7nCe62OdKmu9a9+574729JCS+zOQ+9LpdBiYf8OB9rhy
/qWjG5ngqPY0v0pV57P4TIS++JYpzGZYhdqhtdwyeP+yxzb6Ke29K9UxJ9VjIj00
R+jPNgd+IaSQQO1MsWWsRg==
`protect END_PROTECTED
