`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLhg/235wZZ6gLDIQji5kHcvoAwXa+zEwClMOgqpDpqP
FZN3XUAd7zvxjBSNgJIvRPtGP1hzMZ7+au4aNpSWUwpYasXll5oAiFqXOVPJULgU
akjVyBegQAi0M5wWBiCsNnMO5DPVtGCCzqE6Mw7YbDeBqPH38Rh8kaAulaHuEron
NL5kq3ZKy+QzaBx9PvmWB2c6qhJfi86GVKlSWSSw8Wc2RRLiZXyVsZOvZ9YdXQxS
MazxIvMT9ZDVzEYOWBcazEUz11CrWeajxXOFRIqN7NasF0FweTpDrxRm4Lft+XNi
Tc4NxoPpnrB1j68nA/UPyGwsIn6KNOatZWZCWqzBOp7Zqd6f2K07uBzS4a8teoY8
ow9ThGkMZ3sBz5d7FDkDvm8T6d3/0/LjkJdQygXagO/TW7KyhGP8UqXTBuirKrQ7
MvlPQN44qDCaqRzEXyVpwQJp7amknlN75WbUyCXa0Wo87Hbm8cdZW20haIWkJ78m
YASThUXSG96pW7N9WIDyZnUULuQSsZ/IJ2UzX8Vukybva9+/eZaD6fExxLN4Q82O
`protect END_PROTECTED
