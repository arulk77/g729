`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73CzsMOyOwYONEGj21Dx33qN7JlgjpqQqMkvugcWYLHSkY
Nv7C5MPD1OZI3pvm4wd3t3CXWmjndrWhw/2XWVaR6ZY2RkljCm3vEpOSp2yTR0vZ
JVLtRjWicI1GzbULmnLpQYTZ60IHSAP/Xx/HHm5jBSK1KPHLLpjBbeTiF8q8sb58
ZcU7I9QYh7zSnL5pS89dGVPLVaRGoDCCBLu/vtztKo4vpIrR8Sm32wYMpxNs8UMO
E+aVL+E3CTlDrYozm+/PRwcHhQD1bwXPV5+7MbQftbC6s0AzWP28om3eJ5RAdynR
vOufEUNiactEmkrpzFBWik3fQRSTGiRMibwlyUB3vucQ3tCMajb58v5vVP6ocfPS
NdYbB7q682NZaJgMSglADxb87+msreCniDsn6Dhea73XKkX2cGv4FwlKRv35JrqG
UMdPQ3OdLkGwB28vJGMdouX/ijVWZ90Gp19Wi/JyVv7S4GiRCQ66rwSJGdUS39Tt
JlCvRI2Jp2t4M4TASK4SNj2+6jsmTJ0v6i+DkY8yLUOyzuJgh3hLUyd7nQTePUVo
imSJ+fh6GW3d2gN6AzNEMFVxQ1F+HfPd0VROIQvvcRAm3mJWKLUWBKiRG89b0cvh
DBxn9mjaBIrVQcwfNLPyMWPPeUllmAWOQCccrVVo+Zafi22m1zLhosoZIZQ09rDG
nfDmWV5VHv+fKk8uXwGnl3qkbrDHHIFA48xTMH/+PooEddBio3ZbNJg+OrVM9I9v
E9+HdrE0LireNVRRfWEG1k4elEhQW45y+LQMGHulZpWEo1M4Gi1mOsbljm1V2wts
0HOVfwFUKJu1tLDl57H+WcWHr0Kk4KSlG7EBpL8pM/Pykz9Hk8cCzgR762L8NYNJ
ytw2lnMSdJU/rJKSxVhYevq7x/SPiud6+E5tSuvrpXg4gkuPZbyU/ds1BJBzUBOv
DdWnjqy51qK/OtOw8aFHM16tMjrX+bz0kAqegWBYoIy0o3zjXnFid22bhGCA5SfP
DHp1N5P6d5PdsFd6G5CAhA1VPG53jj9OqZvIEZHkw6aMtyPy5Cg5vPbJqjkuwXdk
jVsUeskbw7McWMHkU0vZqvGaSEL4Hcantk4CuGcgu8QtWJ1KMKi6HP9CkpgL0Edg
tQRZruWZTcddbx6QzRzrBVz3YUi2C/D69JqtWbyna/5NyZnwF0WPr1A1U9HfthjA
F9cL4vlfTkWcAhYFDWs/gLpo0fFN9njxWAomf6eFxYKSbtw1xD6HkRF7FWZ525J1
8JhQshZL5dJy+QXfb8U8erF8Oh3nFz699r5Q/TsUnH0kgUbPMQbomkbM5qBy4QWi
Wa/uoKGt/Siy3c1iWiF/Jgj+gYRxgs8XartpSnXZXS1QaIVreaHDAFphkUXk3I9j
UUQxqpG2mRScWuol6c5NsqKgsgbCZsgFRKF28l1f66KaiRrHA5CjtlU/P915kPpQ
S9J5C+lXswcpSKhHq6z7dJvkqigIwSg8LUVn+4awejFY7KzMvoEAEKj2XmWDbFkW
VJkWSN7urKtkSYPmdvfmYl2a/W2fTzuYEIB8lg68BdIPgi/5U6pcsog6amMJWM5L
DZ839jC5sx+jl2V/tVNymHNudGFhKlcXZwkeh98gKwwpqCsvnvDGWUqU4NX1HFYA
cWQz3YfPmUazD2U196YhfteGC5GgKaq7GboT/t0BLqR4xgTCkEF4hd4jkUUWBfHi
1vuyI292bcXYjJojMX88L/OVBekkUWSKzEq2MpdxmMnv0Ak3OoLMEM4lqD+dp7iz
Ly2k6HLbsqxvUJTM/guV5YC52LD7pOMXzSHH9gthF14yCD9jCnvQcZGQaDcczVtc
Cn3tHsjcTrfYYHRK3dMLB0gkB7Dn9ErNRr22zJYVrC5j+Lmxgw0MNQB/QUwcFXC5
mpc3SEeyDNCGze1sbyt5sANFpP9bmmUUsBRygbfnuGKLUujZhT68g76GySyRB6uf
GUh0MYGLf7xNVDfvw1GGSCw9vp1LmLOzEl/Sl0bL2n6UpcdLS94VqdQG3AepQhj5
t0iPL8Da4O+XyUmIIwesSgqDYmHoloqD8o+GuVbxBbLtecYJce1eaForjAGEuTNk
n9pVqY5yMhdNZc+7kYjLdJqESdBCWLuY5RzVCLNlxGAMNuuH3G21UcqfGPwWqYeG
68Ye5mdSrVEE2WmitV6vQJigACutEoiHFOGEDSL+etA=
`protect END_PROTECTED
