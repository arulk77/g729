`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveARk5ARGymwz/RLaXaynIbm/II1/fnbsg9ns7C6+oojK
nx3UGYhxfaN9lTjsIaRVDkLUCjK0hIvf7I1JcwLKU7Y4EREW+287b7K6HzFZ7X4i
ET7zuHk5YBu1+yB3INXZxZKX3yCHw66WWBQY1urymb2th5XE53wBeEaVA0YkA8CX
yL/LdAfh3zGTckiNfLXEPQ==
`protect END_PROTECTED
