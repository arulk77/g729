`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46WBG9l3BqQkkGr8igQSH2LTdRYmJXNATjFcMKf2IJdb
BYNKT0YjXh8ncbuNBBSFal8ekfTuei3DWvQak/H/2H14dwvyiD6YzDxJ5aeKft1F
+KB3G1fiJJ2L5bmcdYy/uc0IRTQzqzHt7PmI1NY6Xli//xFPQ+WW7Mylw6Yaxdy5
C/ETIx3k+xiX9P0abIKa9t0IZITYDC6pmvtBIsW9nuufwDeCru9BuiXwGaPs8pV9
hiI2a33WHUCVPXOkWxhvq9uWVGROsHpnxZbz3PdgrM1p3D2o6UUIQVfmCKCPvXoN
dXaPzxjyUS83uEIjeAmhIQ==
`protect END_PROTECTED
