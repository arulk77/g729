`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42Wivd0t9Uraux/eWHOj4ZDO2Rp+Ld8nWsd1nbspZ/Qz
dFv8ChEb79r6hbN5LTLjtkpCvlC881XHF3GubDyk9kNtpFOLDlRtw+AthCYZ27PI
2o+dmWOgs9pQgnnzyQPvwh+Qlw2iQ61+28ZyyUAzmTyk/yoUrj5SP0pEN1LuOvJc
IjXY0fn21ixTrLMMzLdzXTj/15dgaNMbDqm3e2xk62Dy8zxYqvvI2MG0BkOu1IZ6
T4H/4AT5NxR5Fj2gO8o1oPRiQqdSS4k+fmLm6O9S0YMEfgAJQBgjl+GPpxZU851i
UU/jyoJxf6qdMi98DdAh9Jnci0mz7YR0kWIDPYG8fMIbwsfssV6e2pQJXjLchvxW
fe/VBjw/Tb5oKO7Ydm7fmw==
`protect END_PROTECTED
