`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
AGi1C5uEEF86YnHyYhOCpehkkkXXHRKWOIpFALzo+EpMVId1LWfcKUdI9+doYc8J
KiJa+4wegzleNi8LiiWepCBlzn4XLvA+vTqQhd9H571A7xtB1RMzsibOPAoAbdPk
pRN0v405VJlPT+3OEAnOwFSodfSOBbx4/wnbni0hUMcs40tkmi4G8A//VZe5S0OP
1o43HHH7CIGUnQNHmLnt3xqOkQNm4RAPi7AgvzrIb4gvMAqNCYn91kvpJSPLLraH
YALtCdY5qzzrGYWs92oU/R9T2q8Ww/PJR8/VA65jCH/vLRdDHkJkWwBlruUlHWQm
tunJ0Q6ctmmzDlvXdifXRGMLA+r0li/cSpY+Xm6APAMbM+tiegvfhZmzmAvbX5Ir
GpCRAQIhELedmdRHuse+sTJhMVXrwg8JtsqkuOW/HCITujGbCuJGxuw+gswjtb0q
qMLJgDelfgquxFX2FQ4cw6hiMcH63FTI9FhKfsPtC+lg6ldci4rY9dPbKHVWDg/I
oXqfSNJPkzI9jtvVmd9WOgMCFaz2iop2hmRV+Zpcz20EO3OI0mt2KxCenCFDu1bi
vY7Hyribboiuon8L8ijc4S6Vpj5kIsb0dvRO4WPhBDXLtPK71yFMivGZm3kTzHar
lOhKCVvqyfgitay4X81DKMj5SR1Ytnda1AplpYXqKHTK0fH8D98P3U/Qj8ZQOl7W
KiiEOVGeoTg3uUlC58ZIU8i5S8QTw4mH7z3DgDqTGOI/HWuGx9pfKWgHlMeZu3ch
vH7YfE0hGArVP+wg4+LmdDwYwlLtsJSwN+QRbUoHNYw=
`protect END_PROTECTED
