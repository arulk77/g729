`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73CyNQH4N7T/55cz74naRk3ANuaxTdQPIpAyso/nl+niP4
UIJ7jzdaZETf1eveMQ5jFF3ee0ibeV5S51RF/Z1eHhMpl5Vyl5TbMNCZyxy3IX6C
OcnjDDdXdHK/tPehM8R5UAOTj7C06ybleqMp0Q8fQicJCIXs+TIM4ADZp3A2FhLU
sTnKDOLo3n2yjXctiCi6CFUXXxX/9GQwhkuG2Q8KARXcDv6FjdF3HBKt8usPJKD7
BUfxn1nFAfdh48XBcIw8chPu3+6kaKA0lf3S6e2mnDUv2g09npb5QwgcYUCtKx4v
bkcBN2WuUNiMtVDKrImIj/tKnkgZXsBmqXpKzOZ7+ooh+r57jgy0P84zqi14QVgR
uV6AzhN06g3rlVSoP1ZqjQKmavNOvw6qX+XWMNnm5RSiDWwYXl6LcrWoV0R9hn/c
0rS+cy7MSJODO/3QSCo1gEJzl8/q2sz3ZZIz2Kwp2FiMzwE9Fm3AKtiRK6/5S3mi
9as3r3BgE9Wm//irzjPAWhfg9hTilcLSbuyPvMxANoGeeP16fvgfu5XEZEzMD+pl
+rOWL0oXVk2qH+7eIW6kLWRxPWgUFtQB5LPLn9d14KBHNecUs66eytCLz5tcIz3K
YbNvM+uFlIxCvnGMb+g8yhi0ZA+Urz7webd6FHNvhGK6m69vSmwjDNipWby6CORD
hUuEA01Gz6whZ1uEdqLgazLY0hOhfATSNrk3vhinNlpXt4KgvU3WInZ/0jLkj6h6
+7fk6HlS2fXfHL7Ii4HLJTtkFrc6G3guEslbO5xf4vT7dsBwcM6+cDuwM0uio+pN
foxf3jOw6GQ7dYdzi7lvIMr/TDHCZVD+21EFyeVHmXDHyW848JLm+V876vFX05cK
edT6QU1XF9/IQK/LWGYU+XlNh+7sfbzDMiIzSukGyoAuseiPsQa5+uxfZqtmQ0L9
GWjFVip3ArdAuZlfCiPPTH7Yn3VVY8w9p9M6e1+KS/MZQKa0dOpQtzMAeonNjI0q
jHfpCX/lGFYd/RFsjugVx7UR8jq+HdQP/xUEAXeVPqifUQOLvEacWvnarNwso7sc
NEzJ0e7x046S+elE+DslPtLRfvUlv5QgY+pDwvuo1iMH9g50k2NrCPIkz0mQ+ms0
oX2MK9S2gxxQCF6kPfiQD43rLlvHQAVof0ECsBH1EI751tAmqCZ7Yr5WrkNDMHPF
iQeFWQ8p3IqEi+sixwlpMloZa/YeLAdOUQoNradkIHvHx/amUNjxzb+CkGcpEAcf
QNaOGxSdP1ri9g+6yD8aFI7QVosfKvWQlJVDV6EbcPfbWOc5H0VbpIU3NQ17ts8T
W4z+rv0/9sr/yezYsmsHRMxLKCUzeVZahQzPJV7Hl2Ej5dku4+G1eIxU7KzMiune
6KPFQ4FUQroQhj32zs24ZkEmNifRt7FYfOwx62jQgDasH5mpGT50LRpGHgi1XFQx
tRNeci8idpVxOKyKFddMwxZtsNg7qjAPrk7tsUVZYfXvKM7kQcHQgzIOhn2o1r/j
rH0I+o4Lh1oeOD4zJUZoO0WzbDf+eDButTS+bvW1HT9/n68M4N88pRA1kBDTsBJz
ZH1+GHgiOu0sQncuDwNa6CnBy6oU3DqCqREy+7ZmDA7bGQiCAOaFSYFDmaOtiZkQ
oiFXFYID66gvoib2TAOeKipJdROkzf0Bt0ExlXYWrUk=
`protect END_PROTECTED
