`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEtqCiAlDSAbC25I4m2qWKm5dRptSTDuVmx2A9CQzgMC
OZY/KPa/QG7uQqdeISiV7GxtJbgvLZV2H5FQxdlmwY8mXc7Koz4adAFyQeSsXajM
mmOy5mFs/QOutq0AjSxjWsrDs+yxAiRXIZAuuCr/uVJRhLbYXZReVk9sOPqAL5so
ZQts77gwpNhKFlE4r3iK+d+NE94xfEHwrI6/CikJYTNG91QjSRKAJHSjzadtGaeQ
nrXNbG0Wq5z1nK7Hwn5SkWKhmeiPL3Pp+Iy11V5PVKjA9KpgXcqQJJrH5xjQ4iwB
Ybh8lT3Xvb8AikrR+noZkmAlC4ZQCiJ8+fFlyc0KVA4usIbpkEoCvNUFavp0S4l2
/jpeHXCVQP2b96wLFfkOfRQ/Gq4dE4TmqMoCStWltthde/ZoYNcxKeC/SGzutFOe
+8eSOLD3jJI5qnCPVSO4HSyI3IxwzCC36/Rzq1WLguvoS10NRsHbOn9XBfjLpqhf
s6Pi9WgVDL2KC0SaQR+vLKQzKmYlBvXar6xelGjJh3qV+XWfYDsYEMQDMnovC/+0
ywUY1nK6dBWiHKG2Gu3e0krT1Scc8iZAuVbd60actNXCz+9YjktllxLbJDhQFoaI
26VF/UGeByB2qkCwBP1IFskzM5a/mI6f2msQ0+FX54x7mqzDSjllPy3e3YHd3E6W
XJDs2RZ+hulrYco3H7snMWiKIzoYR4Z6Vmzms8khlNjtKycg6qcu5MOC7QUhWOZu
amU59jKAU4fy5uvQ1Nji77RvaPz/qi4nV1nkeT3w13WqvUkzxnVnp+7cAX7q0rUl
u7ycyZqPPq+4PfumY4GoURRmJR3LOxq5J2fqCk/ETHJ4RMRjz1yX7udHXRo4MdxH
SuIf3VXzT3Y8rabgvCsPPhYvouTauNf1EhN/zONUVcCMnGPx4v3jY034FIJSrbpy
L1FFXBPrzJA00R72KDm64yuwvmqNUwsWxr0xRkUStaDW6Obn423yvh7WAJyccnHe
gQS2q8nxI2JXa14HgUhMnU6QOXNSSw6FvS2+lc6RVCGy/2TdHvJf29uPh+Up/hUF
nL8hQhVBk+/O0zPmqTJ2VV8853Nx0gK6TpZuO5g/v581mPXRaikaLbdEefCaa93n
dFxr+gACqIsguYPSyXc73V0kSOlgTlEgOESPkUmvMR/rY6XUvb6U6MzlaTSZVVbA
Qvo3iJgZoEBO4XMxbGHLPQUENCg3Ev5053CnHb60RL8X1Z9/S/HWcfc3jGF8ncKv
dYgtJbuxNqI5MAvsCNq4mxd0RmAbS2kL6v1w1Bf7a5buVfPlM4JIPznVZVcCZ5qD
77mYoDHWPMT1nZwpfrXB7G3LniVm9kVMorG28cPy9RewKSwNiF+z+N7yt16Fo46q
0U0XQYu3JYFc3pFhq1YIA0zo8WKM+124HGXSdXJXHZhcx0b7GA3k20DnCkiXoUQy
2iF11B8zIgsoqv6FdPB05srKiEZuvEnIVBWKcm4TNCX1XUDLENRrmBi720UWtNso
23u3fEubqv3F04ET067d4GEmrr7otZT77SwIAS17LVRW73tUIrT9/AtOWUPX3hmB
0hbLBYYsnNKhVDCm0XvpD2FAKfLspIw+LS61cVeeA2y2lsl3P14yYnPi8sn5oPQk
6UTz5oNa/At3JREO6N/FqATMR1QgxGUvvtP0uPuDaP22wIm6uBYocDsziQ+2BpR9
wHfwzJGi6gGEkEgdRQLKn7aZgzrgeT64SdX8Z14PMnBTjOfhRNcUMuw2OtF7Ompq
6htSvU6ytwhaSsEjzIZ5HLMpzUlm6ysdSmtOhbw+ka+0KutY+xvuS1tuiPngNUpX
ug6k91U6kvb6taEF3Nbp1S7imyZeLvXusZWW6YqtpujqhXrZ4gdZ1zt28+QcL7aD
vM4/5it3WvIHKwn5aoTaOFbkprR9csMQ+5yyMCZrFQSsilY8yP/h3JY2wmtqRS9D
y3b0GrOqX+y6TiWdJaPJm6+xE1PCfL0GCxldek/NMPbYjDPg8QnxY1U7zZYkCJUX
90hTBeiHTJ8EVYeF3/AJWBX7ngjZFn4DdWROZSS6UekGJSMWtCL4+NAI99ghkkDI
L/AoqSt0UjsaKGVmjBbnlkbG+XIvIBEFDqALxEqPxXsbIm3i+8rkarwx6FoG7nqY
u158x3oKVua/R8d/8VY//XMPulKtzBzjqIwQ/oeW5mUSng+NylqlJtLmAVdrOPaO
ckEbiWcU6JcZfQT0lVJDTA5W2S8FtIjTgzjWRkmSPUMD3RmJSLwZzx4o6GXl3QVf
5yyTOAVkfeP501iFQW+PYz7WjJpPzFr1IpC2f0StT2hlYs7Eadw5ja/YHDowVMlO
yjezM66XF4n4eEWhKbcM78F97PuP6jFOFdFhoKqGj37M5KBsi1NeVkTAdTUZn/Wq
nQIoNYB2ase1ihSRnB6IyKGXib6NIHA4/zyZuTtgZwPhNntfapGZt7ea1MXQ4qTc
1FXRRQBI7bEPiRYNs02utzUOxCaf7I+pw1AkMpqC1oMtsVSot+UIXVfxHHqWrmDU
a9m21YZfyO3TGtw6Ha7wJF4V5QlPXsVfRQY6/0dmp4sop+kBpHoKNLr7uOgvDl+4
PKW0e0Jt4HD1pWCjWKIoS0nTJXGfvlRQvUHeNyMKZMghNdTFZNeXfeSvzdavbsdu
Ek0MD5oI4WpE/Kpz59Oh/M2X/piyNpuWfod9PiEoeu65oqwqn8EvkWe3RmewHRaO
zFsqZmhO7uATD4IWkGB0OO4+4y92R6lvkLlelN2lNQ0K/T8SCUWPMmFWpobFK5gw
hFoJmhFyu5Wtog5wzSqoOn+hbt1+YVsdwzfRJmgRgLYFJyK/Vu1s66dGpScAu9gy
DiRHPJTOiXoxPRTGlfDFqC9DqOS75iJNAh1kf5fefF9gPUdpaoF6ngt3mpJfU86B
DsOkjQF/kdDlccmRKvnobtTgVPbRLZLrtitSfKkA3hbMG0LQy+glI/73LU6jKp5T
71J3GzAcWWC/GIEmifTrBv5XP5BQGWP1TQrg7ATOfj6lVJfcNPEzh+Yo7rOp2x80
iy5zbd/asdhYPV7quHnCdQVeY2HYX0rCQDpfBLHd/Dt8R7iAiTPRMO4B+iM0zjex
P9CPX3cx9zfkZ5PcaOLSAFjGdrBx97jJk0FAXqbje6e7bQsPdcM2x4Kj3Fkr45G9
TfiKrR8RxPpfjLxFsibsUPQmjuVmi1m/2j6+j5V83NKo+I2pdtvsI9B0JcccoDFq
OpH1bNF2VYukddmHaGqm3U99+bM0xf9S+kIQF2RJ/FgXvljPsLJN41jLgUgusXrR
zjLS7s+bKSX7YZ0zq3Zbp9RfsL9t6d6dVKuVWxQ4TQ4Jk5pf3CaZ9n8AiaeHsepO
yqy0Hzj2vmI71GOwujOLDd93aRh+sRZxYKRj0zr1kjvr2QBrgQevBG3eNdWHm4vt
2it5NYqPbOQAAuNsUe+/+MlJBTaneHfZC+Ix9ht4zt6AHtTuY7kjU731hHCvtVrh
DgetZGpTMv/E6BVkz/CsYGqvrVWY67BI7AzNPE46v4OQv55PEzyY3DMsJLK6wgFY
bJVRppY1dAv30PnSMYp+S0CDRTcmMG4KXT/GyiuBpZTH5Q6Y7djdHZT2Quc9C/3z
BXxzLvSVOPB3KfPtRp0R7oNYSG0wnw6iEbLcYTDFhd410sr7+SgsTivyvp9qBkbK
86Z3X5hY+kn+Fpg6EMKHtX/XQI87rHIGOr5XF7dMv7sIQObVxAPHOgrxQI8gRD5e
83t4ndKknCE3YHLPkOirm2oWtbTx3Y5R4T3EA92mLdJOXHmZNvR6j2HHFXOQf5n9
tpYlvLXpDVmkoXMkbnulM1o+R3INPEqo1SG4KVXCuCVakZYRpTGro7DOLC7bICQY
ZyIRzxXqKm5dEVeP5Cid+yKwI29GY/hvEj1v+ChQGvQx1RnQ5Vqjf93OZkE85AlC
jwT/xCFVi7+uzil2jFXdZMW1TpLikJ+n/t7KF7ZPratQKQ7XGccuzWi5XQmVFjiD
qV+T4HcpHKKK89AqdsalLkld1XXtclzxt3UFvqh5wBvZxx9zV+CnGjoLzfqMfWms
AIyZswPDeRi42bWPBOjYn3xvBQG99PrvVRaxJaLMB+M5KZ/3j6uVXqIeIJrErcNv
CLbGJzvoAcC7DBQZKDuc6LZOgNJBV5vO0xxW06sLwY18jYF9N+x5fW5cj/E4K20H
QCAHYTsX6NZB3TbFWlxbrJBLC4XW3devjuMVE4CUYE+aucbCMopwAwtQx+AEtDTp
P5zzRwp3KdHF1y8aXVbB6Fpzx+rufRwByolrDZTmS7b7uIzE0dHtcXW+HWkxFqkP
VrWot1aA5kojYNxvgh4fgQwXyWmQTJ18j+dlSwfX7tc4c7Vl+scz0GiwHoLAF6wZ
Hsy3IBdFGbZAx6xcIWLTg4Z1cIYbBQ4fjtkSqggLC8m9GXFsGnNubm3FKzHZqgz4
Bz2CraLyx8WqP3KBxnSKyNuNk/Juv+I3DR8aZRDENkZwp9UhUI7a8q+CKpP6/CL+
7ZD2CQAVaBDgh+hS/21JPU6ko/a56jVqcXHXvB5jt3NShgEpWhs1VwVpcVd7X62y
i0TWdd8Olcn3baSFdFevQ7XQnpKE69GW7FGke7IroGEcegeeLeClTfLwSbTLIgGn
D0owpuhcUmjRyzVPZhZJaM4fXkYfIkN016ZC7I8kVYW6Ka7JsFMo8OUmNkyirkzJ
kEysrwbUn1dDdV9QlJR6QM2id3dHW99ACu4HBVXACQcMacUCg96+ghQ0dfcXg8wm
nVB7UL8n7k+e8geeZFG+10sVF1JfuRv/n4zZxpwELVL/32TJ4suf4YjcjnPtjhA3
JO0MTT/OwE5ftEPetEUCsbg7AFpXh+6BsxvzyjNwBi30H14k049xwRmi+MGEFkrG
NrfJumYJH0dX8WUKZNqDR1Ziqx37qFufpApZyhnHli5rCWUqSwgMZ28f8RYFpifA
uE1CQsa6We7CfQc9nUuWGBsJjqrAG4JM0uYiXUcc9XFe4uWiC23MnaPRnmfp/t2I
J8vUmvDiatiQEbAu415e6UCg1T81OF3NNUkxNoGM7m5BZii/YTPr7UEiTtDIgf4g
hj0BFrHrv2La0X3G4sY3QM9ETNcrWMupOLMbCOmGmHPqqRPp+52z/yIzoDJdM6m7
3War8bv9jOpg53KkaGiOiHG3F4mbbJH4+EpfsLN1EXKgyr73NvWPBhZixwxui3Zu
BMWKzaSY1Mmr8CObl8TMhJXUJYQKuC4x43KMni4hl2rKd7ReYicyW0Yvlb1LiZSH
Zm77F6VoQgYrnT7W5iioeNPGuAZ5lEV85LT/jOzzRGY0/7Zw6WbhhTx/L18Z4zS8
cZtMPekLQDOnlKjpqMxQhibPEpyEKwOqQrzDR67z4SgfLfq5Addc3zX3yv3ZuSeA
PVN5oG961hYMVFiVcSwIyIFRtkB2RCvs77ICRs5uW7AI1u8HkqcVvr0VEULrr68I
Eg6/8Rt7Fj1SlDV2X0KE/p0djoAYtYJRlO/TMSnTMOjy7Xy/aLNSzUSKxlOXWUjB
47hfyYwIsfGKUx0d6NFOYk9dGWhRYUC9QKN9vF/V1wWzb5xeMwb6fPZo/k8afOgp
jAkV6e/2SjvZWn4N2XdsfuXn9Wv7upWL6x/dGybkNegveDMj9rcdVATsuEgdXe/O
WUXg+g3d1B2XcUWwU0/5uo5XWmI1pXlIC10Cc8+eaYX+eEF8Hcfth3kVf/X7X11J
tPNAKozGKWwBkbvIC9IZwvbKGPW4mFELvY2NaJCwh6TaevBwJG8U8UfOZtTs+Su0
IZ8sB7eHuF8CfkUduhQlbUWQ9a866jOBmhrK2e2QpxHu1ldPWa38wf0eVlKdnz73
LsxFtXF85xIADFF1jkbsqLR9CrCuP+4yIuD/ptNnCI812mnN2ORUm7RJ80cyOkgS
uIDUGgy7c5YJ1RxvlneXMI0Hwb/N8rqtYT8JvhRjQsUMj521g3OEc57idE8n2UQk
Px6PJRBmUIgcVKoOPbTl4CfewWUtJbmN6a284IEgrXw8qHirWWDutRP1pm5n9Dxi
OKCXT2+u9dHeMqI1ahJTihViASTLxJNnXnu1qe00qdSZa1c9kgtaIBwIdX47Igoj
Ed1XCTQ34qtL9YNA9sB6Mc3KSarUixL0GK9fsOW3rGNx+Jduow260XzoU8sb/5SJ
IN8OVXR0e4X675POE7nqSkt9NKljIQ5VElPLoi0oNrN0EYLlybR7dGD2ZUUtcPm+
aPcLsguLeKrLah4LOP53tLsAq0Mx33/1VyyI7/odjgIFVNAH7Dwz83pB6wZIZzwp
/RX5i9beFVsQmpPw/PqpGnyF5hU91QIN0DWI83wSYTC2HWsCp4V2jGDStnVyJFgA
/x3DooUCOxGgNkq5LKME7tw0EbJKsPdGujJDRZmYt1vrvvnsZFwMAVaWZuZFsPeX
flOe/TSBPZoG2Jxp+66BKfwjnSJzEQNKWuRqmEBbe861+N5cmGYv/ERWVjnieRwp
SpUrFyLPhyZNFewPzjHNAK4t5E3cx2einWPEtXHjFwV/LdyotPJ6i+0GF//HNdVm
8P5fOEs72D1FzxlJ64IOLRKgWS01E6uZxA9/Mxnay4fVbZg2NVqrkAKAo//CkNgE
eq275a2ydZLbj4xa+Ai0TqG4OIbCAkiTTCsNr9Zoe+5f+igQuTLmeH3xk5qJPeb9
gXrisP1I9zE2F9o50TjVOGsduDkdhvMTfGoFme+2ioG7BTNNDDV44O6EaMVo287O
hUzR+2tWyGG/SZrznaBzfzWbgCZ/lcsJwrPPZpofS7pUe64maI5vyq7VpLgZwmMy
zWCZPVwZiHZPZpYOnIEvatGxmKltdnXkSnjFwMnu+PyaSVSNGRt3gkFDVfFDmYjP
X8jfIBuB6Piw6sWJhQmdV1XYiT3h1JWrrkaSq048cOxiTqZpowJZhk2ohIrP7FAP
+TAqYhWx6BQ2pxTKO8ZRis3eQhw94/Ui5YQvuN7qH8mu3IvT942Tt844CMv990y3
L5dXavvghnhf63W26LFPYoakuJKkJc9BMztfPstHPCROKXxT+p8IxgtC+O7BOFW6
Xl4YGDovxMH2g6oFEY5DyujNft5mV6621xIAD3m6NkZkELmQa417R/EhZ0Unwq5y
dbinrqCuyKVxd6EI40u6gygE6XStsNO0Kki+bmSQjxa5IZn/AJFISknCl5JbrniP
zpRw75TKRRGoIkXaw9rBrgqYxuSaQFnSoR+dxUui3J8/RZbDg360GnizaLfuuqdH
7wRv8EBtJhuwiawHHFmNzpRi55syR6C610g6FZko94tDD+EhQaMey6heZZT4w7lj
B48XYuSlxba5vYZtknSRhBb0gpEgf3Bu+m7TFbLVMs1vnboqLKccBSNWQwRxDtIe
CHfwFs2zUW/w/LxS+tujjLgfnAhky6jT0hqmK0bvXYHMAciug6MSCem3HXdxQ4kL
iNsbO4+N/KyYs086keEWBxKMJ6WXvXwQvfLVJEJ2LwrkbedIcfi+246GL2a1F5QU
zGC38IVV/NPRFnhw7g3LWRl7ea16PJz5lFpZxbwi9LPfUxl5H/RkUE5uC/s/h6m3
eta0EQsA/Y0/Yv5y6R/9xGb9MzDUIsVunVGqv/f06laeteim7f2XyICE49hCESdD
6pTbviF6mKVdPWnciiUO17lfNZfO83oKZgRPzeFqO4C+xZdmB7+LKbl4iPRmV+VD
nQCz1TcCu8MmwmdZkt42D7i0wSxESkRNAZHpCESD55AosU1AgZXtbs+2zZ2rZuyW
QEUFNFOvfamfEHLcClVAcpK3Py5QjUZvpCKDisMCgOkzAKyXauGfMl2+HmtvCf20
KztEhaZMlmW+2zGlt2+4GKAMkA6ZC6XoyTncsGkI8ozzD0IkQ2awtiKR09YeqbsZ
M4UTObDBY6ghLJHKN2LrOxpT7g0H4fcv6NmP8HgDVzzAikZWKr2n+DorfGF7sdA3
FzbC8+Qp1c4lhTcFW0vNJ/CnLCggGCA+u+s3125lt56qLrsSnO08+du2CIkAS/7d
4GJuqp43RBT+9R2oiktgM7YN9weLF3vZS0UOPPXOEV1EvKvk7aEobvkQVsDnZCOR
7aK+P/BopQxeJm/snmUBc4LJcTTnDSLkneC2pooVFHXrFrrVZy1UELFUh9C0MKRx
JlS7sqsCbwv7jg/xbqa3fpRoVNcB2EvuXaoxtPHMWTIlqmrpdg548q3sr3plWurt
+5VUJlixg59hBQFwED1VBeldL17F0RzouUm+spz2vkA50g21kSvWCB0D5hiZHDjY
xOd0/lCcRo2BXheb4XqlM2rXw2xz1EfLIV7bH1m3oW97pgfX+lJP4gMAbE3G3fJg
Jx7dWAOpiQI5hX1vm3cU6NS01f4AV4UhnPg30eSn9WE6R6H3ulFm6loH3JovUnTy
PWO9tjeDWMBIoS2vEIwL+QO77GoP+zAcEw29v2D79S2B+ddeVuLEaIbQOGstMaWB
lNqy8oyBHGm6F84F/F9qfiN32yyzbX6SkZke1B91bdEtiJil9AnQVvbmUzkw/TlQ
gfdWLYI12S0O+9bLbsd/Lbh7sZveNsLlS4/4VEsz3NEQK1AGEKhTrOEKDblSqY+d
XEPn/FYJFXDhXClxU/WVml5N2z9MDsUCmAchF8dnYRUyihjIdmgoXmtERkT91EtQ
kxbaBCVv92xRD4KOOgSkch/7wU83FuutJbeSX8AmD98w43V4RjV6om77KlO7t0Ld
4imNkglTJsXaGqkjWoqtwINd8qRIlSCfnNZoSlaLGfRXjMHIbVBxXKKshDZgVMq2
Dz5M8zQZ+SjymjRGptgF48CRVRMYe5rQJblVrj2Vx1WNgOS5LUVG2zsPlfjAee+k
K4HQBza3QYfBt//4duBHYF1/nW2tuOBV1HVRq+L24MUV9CYAZPDR/Fj1LjcWifbI
BqzJsHhn6+AoK+69AX5SvD0BCl0olUMkQ4NCQsAWsJrPlz3kFkm/gO57SPf2bkpa
beFqvPDfrgJ/W8FWyHUEzv90yKE19X2xB2X9h04V8Ei48kJeJtmMDydWCEUA1Ish
hfoXxbNBhSsbdu/Ubhn1kygasmlhzBJsZh5fp2h3QDC3NVy1DbipfQKSeiaQ46sD
sBYxNBhS77pYgK/QHpkXa8Hr2pG4INdejNstvD6Ps+Ba57b+KxhEX3ZU/c5OWWFB
qpDCFqFVJyAPUdicNABuHfKYp2rOOWZem/Wq8c7hSh61psrVPBZYi9o9s+XVSW8u
wSrigJxZBbwD7XzzZwgqy/2jTkNTk9nsVZ5A8aSp/ybuCrmNoUqlSEjcZtchN7vi
j8fQ5Odka6vo6jY8xUrNn0cTGpu8mSJSVgs5eYMwkcb+UCUrGvxyUOjXT78NOsvH
fnzQdxaMIQ7yJxmUUrDPMfv3U6SRSewGO6xeYCtver4kLZKRQ5t8sOhmNuZJM0Gk
iTRxkmtuVw3uEiZE6e5XAr7bVXd4W7IGvDaZpB14kfejgeL+kc2VFULwlpAzXNfK
fqH5HrJk0CWYM/s1kDSlCE96eFKM500sbXwe5TDMmnQnivay0kV5QJFT2XwhrHia
q0tD0ChiHhDaD04MnJ8Opy1cLTXV2B0cTvXGmMiSEp+V6tSZjB4Br0RX+pxnvIJv
HKqVmL3598rRuNw4I63aKGba4O46ofmxUXI6wXlm/f+/LDbaOGLH+dQ+3NwaNCu0
08mjZ/9eTXuXC2XXaFjEvATLxDpkfABtR+HEWuBbIOg7QY9O0PpXVKsU7L/haVzx
eLyOmGHX9OwK2+lRr5wR3rvYSleNGSvnUlhyCoI4t6GPBHWMQaUp5P++V7nEbrXr
C3a1gdePFPeOPevtVkTPkEPK2Ss62fLy1okgYITlODIEwLRM9JhYkE124AHRXB/e
p8RhOQUswub1BBytfDIixcVuGV/dchWcuPj2EeVp0mVLvJFfXsd7u6+97SlUKsyQ
GA/nTnCROcTH9jfw+U5caSLwdzUIXZy8ysZXbJRKqu8uRWccHPQgq8c8nOlQkBU3
uDYHFpmdVdeQ1x1Qn4WE5ODGKxj5ETIA8GuIRlyOW4rTLq+GJEabtD3reID9fXzL
p3RiyDP50mC9zfl6rvNtF+xVhTTLuV9B97KYh6cK1ZAQOKkeEr83G13BR4GrVmp5
1DlXGGZtUoMWv1UmamWtjQ6QSP/VRMru1TMf8d6OkohmCwdMhpzeUnSpWV5KTZIp
3W0XsiBhGw1b7UGVt/YrW7X8F70yKjyP8dH6wCntENtog0nuLufTyI2n39/jOicB
A52JaTd/v+kotiZWV0SbRvAwarjBWM9lkeojGDoJ+RjN2xBrFKB7kEat1/tBOsza
b22oGxu/wHT+QyhONs6LWTv+0dptQ2+I7fvL5d9XlyKbgP2zh0pD6SwkC9lwAOxl
OLeSkCT9W1IqA64uX4fbNu4p+UwcvBUkS/GiAbqjI5MB4oHM7Z2gEyRx2WO8adkL
aPc2ne2+C8PqqfzXgOwWlvXTvuIYcq0cMXMcgznXorm2pqDSTVNi57DaCrbKFWwc
YBB2g0wpEmi7woeoZYMoluRSEycyM42ZucFlc1fr3REWqXWB4DxftZi3H9E4DBNk
sz48W0QSDRj3Yzm2NplWBg==
`protect END_PROTECTED
