`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
iOWJCtV9Pg5cPQ6ZTAk34L4O13/4t19F5ug7J6OixEMLqNntajAv15wqtsL6BhaQ
onHUUae7aOgXclgh/IFMqhOXCPkha7hvlizUONWonuoYwaXretlCdvNi2ECW42ea
CdiZ2PIxGRJOuLd8rhIRmzfybnV8EUpEUO7xOL0gfa5d4zPGDQQfegXeT98GvBkb
g6EeGAGHtYce5wU73fnN0R+8rWRB3+ZFamklY9fJhlVlJixLYSYUo2qHSwf6g0aW
T60ulhZG9u7tOCInu0DUURUzG8JwjTOFtU3muOwMhdUm5yHGHYL/dZuMiWYSaofh
cntQAiEjZiQadFjlLh5tPH1uygnTn2x9o7rKkLaeZgs=
`protect END_PROTECTED
