`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu499D9x5GIdziPY5ShbOqnKEzDqx2JIRZx0D2TNA38Y+D
TGr61N8+qCVBM0XLs3oboK5YsmCQ0wEHy2mfLK2SFf9H9tvm0jSmaMvXMB82NPFV
2HR5zc9w31KiyWEbuuJCirgDvC75zl6NUJ9thY3ACbVk+sxB1l5yXgQiSpNnudGC
GXkEiR2B05v16ol7h6VR680bR1KLYijd3d3VQxrfBNy0j+EklI+gjrAg3CseQEKl
IkCnPcJ227jEy2ipSdED+WFOgc2JBdTPMHFCbxo6tRFuRRfVVGgleWiat58qjiE+
6US40mlfi2xOFsMJ+YJXGQ==
`protect END_PROTECTED
