`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xIgd6Ad4lPXdZmLr+bsxMPqf53ZqttVu99RsSZeN7s1
V9GrfZgYfZAC65q/IWyJQPkWHx8cj2X5UL44047UK8Bc6ZtzkKVYszKFoeZaikPu
ME2n4iG16eEeErwPmM/cDieFB/Y7gQSBEwE9nTXasDJqcajtVMKMZqDwVmDU2ZQE
C9DYtcUGOi9jSpYTt/23696NPftVqE6K8AzJ79B8TErK/KVnNoz6XXxW+8aWLRaw
hjlw1IsETmZFvl37ShXprDbUKB0c53MwrRFiXgg8MVk=
`protect END_PROTECTED
