`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
eAse3CytsydE5WrL12Eu3FBzSYE38icquybN4vSIPO+QHPNrMOe3TU7oFS/Ft4y1
j7cB0z5zHJc3oUQcEiui/oTgBaKcod57Yelqcxs+jg9bK3bt/unXrMNi1QdSkhgE
mJmxTk6vGcUo2o2wkUb6KjYLn60igEMGOKmEe+zi78Q=
`protect END_PROTECTED
