`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMBMVx4PccRFG8pccZbsiFV/mSUi1UBEP594YMUPuS5M
zY+mjC1pZo1KxRN8h6FoQTAxmbkDGcSrUOBGJouDd3vikIh8jiyC1lgjcXYzam3O
aoQWa9YnDO9E1OLClZbQ89aFUtq8QWReMSUO4OhJYSCxcmYn5+f+/IYPiEXGS7f2
3G2w9/YhYfbIHZUsgi2da/hhoRUBRDl0gs3OsgmttymgPFfd1Lq81B20Yo6keDIi
0EP/wV82QxDI6EUnZ1SIBh9bX6L44RqUEKTkWmPL9wY4GCGxBRyll8zV6Fv/isAl
JlIEjsQAG+ONtWAzBgZl1QBqJiPQZb1CCf1AxUKS5mOhjUnS1c7o4jy8eXwF8VSd
vYotBVMwVJ8BRnB7UIrngYwsr+H5QdSyiZZuX5CqPHa1FnAbpztEjUp2qywIui8a
ghuBKFCRvahfoOH/G5qNkytakI7eRUQf3Ywkf6j1u0rtoJdNpLU6WIdNUWSNzI2l
pc078Gn7D1IbcJysLL5MivC+YlAKqtx3hh+z/a4osk2anYNx8Z6H8Zkap82iCnux
ML8BdclKZy0LD9nzPaUBX5I8+Rnd0bEWYV4/3lNmnL12C8gIOe4xA4NVa8awmtq6
/NMYuYhFblXDXvPnrkbKphUnemG/Gf3oxD2gIdRNzLG5jzJ/Hicbcvnajz3t0H6k
vf61ryaDyJJXmvtIXAGk+svp8I3QUzhli4R4QtUbXHT26sTiSwTeSsxir74ZPXw1
NNCRZf0d8/PR5enWp4Zu08OUrH2pshzVS4HvSqIbTn3uWEULh+ezm1PA2KfcnjGs
kvl7yQLFdQMwNifo46x3IMSCalICnTSNBreARGK/4P+m0qaMgGaH86CTOIVB6HkH
amOGL4WA1e4fzNXM+S5xpOAYDSqCq5SuFrnV+rNcbhxt7W3qJNY3POaBuf6pj+6k
xKvCKltbcj5gXMaF9d/uMt9Ezv6fTVLj2xnGFrlnD9OS89ESNte5+KQM6RTFZmhZ
R+QFR/RM5vu2rX04+au+6RHZGfw65xe9IrVladFdkzMTi2WzGWn96uG+6+TjYoX2
j5879jVv58b3gVmC2vfVkrY4jj7GPIsPobGcLOVdkSYz28TOERKcmEP91q/1LCne
opfPNm/CSxfXbqKhsTZPkDuZoRHeNVNH+4Bptk2g5Ar7oMb+78eS/OhYKbz6XCTh
p+kK0HdvDKUqcR/TH67j8/y9MN49AzAVpN+5HRZqs5Re8jURe82nNQPLGffDSuz9
cSSvglBd/7SdW3ooaikA/qfH3lfSk0j5yyuMtUy8Fys+2W9w0FuVihMzlm6zliAB
wbiNmNWlyCR/wMcenJufYUxcLFG8uCtt2jVMT/IwbvK9dwjcpF8yLTjD6vP/hFMt
Msgke7VJQ7zreZEa33AKBtAmFIFJMXHZJZGiZVPtf0PU+EWL5lrRdfWx6Lzt8yld
4CEUU4mH2odLHsKVyuVXkjYGBRJiqCtX/TsY5/RC2XCt1E6Rf9UkX5TsP/hR5uwR
T+zoxjkevsoZRPleHluXVBTnnumM31aKPp3Rr8E+RYzKYFMRUyeFlgRo6JgsPXfl
TXWz2Lie8pLH+9WY0aMTywoC5/JBEGnozN8BPE0uF8C+ZYsjnT+gZu6AlXu2rU8z
WwVWNHXFLlmXRCDTOQclmH9mV7x8nwOQ3l9QVYepIxmC9dsU+X0Yp9yYuC19HYyp
gMxMMVb/AfjO1hnkxg8HtnbKbboKkPiY/KmXCXNIwoyyk6Qe2I/l6nVExwXWY3vU
lMGlC3ynABVJlIBunAjNc1iBW5Mt2rYGw3zP//4uVTBzpKVMiDGJ0Cige/l4+ICI
XDnsxM9e/DKuWg1jipvEYP8nnHnhM4IhgLpWQ4GX5PRAHf2QIBdxIJXdO00aZ0Iv
tOlwCAuHDaAIOsOFXbmiZrI1IKUM98CUuVGa/KefJutvP58C7jk4wtcyFpysjRqk
J1ZX34+yKhn9RgwfdWsNoeL3I5tqOCs3gb0R83Gs/Fd6S+yELoKC8dG8SMLNu9P9
kNyD4pezDdR7lyKn1vAd2//xyLuiq9KhsrZsnwdMwVLJSNS+QSLSd3RCBDJnk2ul
k/Qs8B9AphnNzjLHIBrq0Y+PzRzQRcrfxsWTJG9hFlXgBkWc9mFkCLDptO6Y+z5Z
ldOlxClOVX22ejMdMSkm1X1C6bAzIAsG8N5aUqHGn+8=
`protect END_PROTECTED
