`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHAGyhRlFserWFJKWXNCBcEyA/lnpxtBDFgfSwCy4KJm
GwGMG7Z86aEv21BL/1KgT65R6VBz6V4my+6oyGoXGA9jKMiDwx6P6VWV++m7LmVi
CokcCNxrpoH/MlvjOPnp2RztP3Am0zlQ5Zp04lnBtMUsxXuAJZo0uX6oNfLvECSp
jBlVcWciPbZfrgu4ewMEX+B1Gvgxck8tzFvYCl8U5YqOioChpzCy1nbIqf1b/5Yw
e5RlHWM6Ta/Rsk3CYTPfS88/AQ12L0uJM1SOae6jm2UbY7hNamwJGYgmm/S6pMtD
+O3SEMwVo7LmK2/2NHeQWMZ1IIL1dP8V2ZenNlRvjSZfaU4Ufj718auo1IUKun/r
BuDy5RyVVHbQJIqY21NwodaJES4NbZPj/kfzG3kJdn1Ue69bBGxjWohh0k0SpB2w
s3Y/2FN7Cln/WxBKa9eitQ==
`protect END_PROTECTED
