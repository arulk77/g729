`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNxiA7pYaNIF9CYjgDuMfEjNwy+72pwuq5dozCikzuA3D
/5Q+4swNeNoJcxfvVrBDwiqCk6221FT7QNEfX84/S7A3zafGIlqNInBIijM0s+7F
9W47/LXfrtABw7i8dIivk8lMByFH8rUOhvvL3i9DaOxxMMp9eMBkN/45FrG7dZ+G
MMyeYg35uFuGuUYxez5DBWuFeS0j4UPU95S+6NNTHjJqz/7xZ8lYfv9IWUfO53hR
57cue4RuLwabAApGV7FBCJotVyo0qG8f89K7J9x61LM/jqq3cQ1ArfH0+TRlrN8p
CcjiZY8Ov/f5TVc69w/9L4SJJL/FLjIbxSumA5sz8L+PNn5qbbkM6X/hpzS2m22y
jaZewYJ65vRw8+4/r0XikhNN879MeOl9Uh0fwk5dEYcbtjfihWjf4oIAlGLrB5p8
rNa44M8KrrkH3vzJYXp9V8QSjRUpwdn2bajpTCbcxFnV8WqZ1o5Qb7BwpWNsRlH0
e65X4qKaoIQP1fCAAV7+ta6tsdi5lMtoM4E90G1JpNUGvP49NQ8WjWeodBB39XCI
tPWp5Str9Ucwpke7eeBt9M9cRizR/v077X6d0pCDKnzGLbwDKmuCDVpe00y+dGMX
TQwr0xoXBw802mEBF/XkEO3SCj8adtC+ThTCgSDqeq5d9qPDZr8+a957vNZ3slsU
Yd55UnvChR7AQvWoNnNZOWBS8dkfT8w7yW1dOxVhUkEE3byiJZWWgUo7Td9SNXb+
GqwyXRmgNyOvp80fgIbcY0aMyZhsMG9jsfsxjRmqyFznD7Q9j+s2BHMzUlBTqpzQ
pVUZNgk2ROVw77v8Kkv2WN3HIq8UNY4avcNb+2BhkMgLx/Wn5FT2El5qD4ARv946
jE2VAXvy7jpUbhquGvl2p4lVcDz0yt3LgKbtVn5TcOTIYTZVtG3ldRLcclQvXCLM
`protect END_PROTECTED
