`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveA0OaP+mfr+91pJuSclmhTDnGeRLIxzdj7+Htb0t9Mf9
ubgBfuV8i56n4DgknMIvSwuSQQlbY5GNlUYjCNNYnaEWYtH9kddxWiqPpsyBzfLs
x+sHd28WntDJhOSZnHFl9cSR4ERPpgwD4BzioAyzbKJcCJ192QKTK84C+c849DtR
my+dLAd9QCx4DjLtYUwWjzhFb2VeIB77pQinhg2sUteVp2R2r7qhPQz24iooYGMz
WhkDlngO0HBZiyR9W3L8FmQuONrMPAE8moLt/ravWCuQhI3scynoNc6lfh5vGXgh
vyj50osyb3J5Cz/W9Xv4Dg==
`protect END_PROTECTED
