`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIkun2Lw2P2L/7Gkr6yk9uEt8q7V6o6TI5mHpIJy4I8W
yUorNrq1A+xoUMws1d8lI9RyIcIoImpTDb5VQZQtoa5KeDo0nssYIcbJxAyJVbQx
7shpe3+yE8TmVbesOqYJ1H/dAYAJICgoGMUqjz32gLXUPxGn//wZ/jZrSyX5jHlF
sgJWyf7QpPKuIIaMMECqg5ey8ujN7+nOxtbGYE2zr84kkYF/E6DNv3sSOBpKcjvY
3sVRGogAjsMF/98l9boIlRaHSitZ75t+kNkNFHWzlrm82lpS5SSw8c4vvG+GXYAp
+YKa4ju05zOR7okOhQCHBlAd/2WF16vm42SnsGS0FfBbsviG6hQTvFoq3YnHRwI3
RWNGB5kMp4KPcFAUotimVtygFLxpszhqiQN1UsY9AyQiaUoWSh93OpFcgkR+iVgV
swRnWXEPd4Dv8mZtlQgcjot3tK4m5JwEdQKeA/tQnn29HzgIXyhYh7tu6BVGRFfT
Kdra5LPX1mSDE9DvLUGHV3qZcb7B9Ywu3//qTlFhDoPPzr3kZ+fDGjmO65m2PT2P
h9NIKrHY98PvqKfRqu414l8iOblOZUXVt51ZPfpF9PEwOH8qb46BmhHocXjevaLT
4p/cNTs9So4suwknT24/3JhOAAIQCg9NMDrmcBxiqOij7HJy9KF7KGLZwDDYJTuC
nvQoTBNG7W1ozVXWodjukvnJgWX70CZtef7CmmrTeOvdderJRRjDPO7nZQDSC3Q9
WDn7VpXazzK2zYrrC+Kct9LG4cKufZeBb2xkjFQiuuEgnTdr3Fq+TYoW9WYNaiSC
uVYNzs6x5RQ2Ey74+SKxuN2YYmbEmymbOFaYwc1mixzlcws0X88r7T3uxr+is5Us
UTihBjashh4vGnjnPMCt0TBTHEjrzcLyrw9RHo7WHhcDg3UUFBXAwRUJKxJ5g0IW
RDl2jAwLh/adEdTmhSVMUgvis6DYX9TA6EXskkD4jjl9d9ZI8ATXfM2Y7rSnLZhe
znvvO8IWArmlOob8dCT8048bSLlqJUQs8twp+ysB9IHWSbw6k8L4ovZ7/lXEo8f1
ylYJvhyp0x/3GpaZmAM2lLlkiXsPImcaDPOmRINSEOVqVJ+x6QMOi2k4m0oBAyXn
Uefzr4+eLB9FdOwdAyIvqwEjdoeqUQxr6qGcfPEXzJQXeDVP53L/bcDMRe5DNEty
7mwUh2bQAh9ky1EoQSOZU/Qsp3xfVrhdYie3v1wKmdjWg5sDJJ+AlRjtykCoT0dz
nQa31ykIx76h0U1+1Na9VlJ94vmBHUBpKe+5VvLMQguUTsxygM2cSSd/Wt2IT1ze
91qaCwj3oa1dq2yzhx9cpJ5zP6XNT7uZjDZQ/KLHS7QcSJ98h7lOmA77E0HtPhbA
noZBv1Sx5z7suybc5aI3c95tBLM4q+0LOIIsUm1y2087sPEv0jkanR4uu7Yjeq1Q
4vO7U+/WQbUQKeJ28i2r0KlUcWhxia8lD3jLAs9baw8unzfN1/9Fy31V8+ouZWVC
B5X9t65ShY23MCCxsJ/HiimmEJUU5DTAm6KwEFIfQVskchB0VnR8QlPUtxH8spNg
KZ9Eas1i3gMyeJEZyTHPoXPJie47jzsUBtDf1jvAdNlIlFICIwhxyhixo/uOwBrW
rXPUc7lP88WB64Htn/j+IVr412NGBdjoZA6kMmjILx1Qs12xAIBFUJfPa6eFXCTJ
O0k2SGME8umOWT0PBDJMgT9J+qqt95s33Zy6TbqmRlNQH2hY7mGVfaTw67/jLdNz
0ezqBd9ZD9N5SXPA+39F/vOWELzLrXknQkMBYyOnb6Dz9pjtNUWiu/NYrT2398tq
3EMoNdplYKatySIGrYqauz4s4LtF7joKrOAz38S6ypxIO2OeAXRixbqTxOSFVRKP
MUwI/V1ujC+GTMLvKkGkwmZYqKiR8x9I5FqpaLgMPDkSPecIRv4OEvJTeH5uUnUB
tg1yduFuJow9ByHdWWuRKqkqsNZAPdJbMvBf/RMt4MDNydWhHmuXVsAJ3LoYuIoO
oQFEZKR7QRI51Y9JkajUGwLKrtLSMMqfRD28KWBRr+0=
`protect END_PROTECTED
