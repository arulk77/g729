`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ae0zGaUQPf2eqbR7BaYMH7eFu5yJCrOjaJsFznxHFiXUBU/hf0Fs/Px2FMW896zB
gI8m51/LqnRK6KIeW5moGDQBKDNwqJ5euJDy9h7SWipdGPmkj4u6hqNOA5NzSTyt
P4XEP4I4361lKbwkHbViZv0tfo0MxRkZDWZ5FaDPO8BFm/LEKT+itjsI0Q2FRgBH
q4AovdOMR8hDoVBcpK27sZQBSkqvCTBCesgheUm0qTV366XNGmItTq39ExQaeVnX
6c3NpjQtlwIouDafG/BZaSJQXmu8rHJSYkJMpMkbdR0=
`protect END_PROTECTED
