`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN8i1LeBHezknNtpRUSSuAfcU/HZdY8UWY4r9Ow2D3Qi
zghCihi59ArTuEt6EMrnYgVRxHzdoRzRzRPThAB73CiPqxTnmS1XpoiRRh0W2yTj
7nbsUFp6lCYqsAok5wcRb6r1fPwY3TbDFVvj+ejsSB7yQbwh16bWEdfSF8jRD6Aw
q+aJtZtA86kTId4g2m+ZTRVX+5L7kK2SogQPiKvmPiToHIgdFirdfhid7r6PLx7b
S4wdR1R5S6DSYz20KTqqLTfjb5yEhdNmILI727A4Cmg6q6MayYAGWurEqunR5PZK
NH1GDknsfPu6cwObHPf+/7ywmdLH3dVTT+fodubfGKnsRVIyGVp2wonEmR90dkpm
nEMbvyL45TWdpJ1C13y8xw==
`protect END_PROTECTED
