`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAdm+412YSpN3hc95TCXjAx667jNw604URmjqN61adyoA
AVYeVT/l9WE/jjMgySUhSc8/8AzNSBAMc/5M4ZWXQb/6X5+YejazI9mda+iBFG/Z
FZIBERMyi67sWHwFw061Kd1+pCi2+Ctv6MFIEo0UNrP0L9C6CYkEe6fz0ijQvVNT
eJv7daLFh2j4Sd/qYJYt8NtX3sbkYrpehd98xCe76JZp24mrjpdsTxyFJGfgiJ1G
qNbOU+q/GZNC+KoTuxi/0CoAN4DmJOc5s/5/npdBdSP40stJdtI7ARa3bIU7yaUf
Twvr+DNr77hL4HgPPeRAtxxVKppsGX0OaKViuD0zwt773gPPpk37k3+cLFCANCn/
WlLTyfhzC1aXt2rY/VxX7JjeJ7uLwWI8fbsawN4Rlt/U/Ovkdig7z0Knmz8wX8a0
qI6wG4xMSKdZy4+yqYqVnRC+H4QCqNt85b+mvxiuq+GV2zgv2OFwWrVqW/RnzvTV
M8bYOgM8cyj2WtqKEYoAEzo6FYgtRj8GBgkqLRDKTvdL2Gkj6wkowEmiks69F7KC
JBvKlGH0Gwoeyq5NWUwSYIGGjF9R0Y6FoDWaoYxfzQeHma4jifDG45R9jdsYyNSE
tfmWpnAzEU+ISwm7h1DquUnxd7t3w1rq7pghZ72wevFVxtM2TYyqKRoVCCw3O89j
oLlBr+uHQFE6IYHMDIeG4Wz51zvAYh2nNLcbzFvEhNB4daQNYPO4/g2hYXRaZk3X
n7BIHo48UjBmqHzYOAwT/EhPfFEsrPiPJ6UGg7Ve1t5wJQffSg/LuYGcan42ZVUn
D5mkXunM+JHfpatRcoqEXhRomwvC//rVgfM8vrMd8qGSohzCNDlBLTyKr0YHZqLM
4Bw419nwJUPvfSK66F+lKaNeWlEnvaH1d7Cvf599kA2TiWdSL2GA2WImvHbkI4x6
ASF4hpUbGcSOh77TZkSkP3vsXeB6VjPi9WofM2mDy26YU+/F3szvQ4nE1OcnBaWE
0rmVoa6cGDccktX8Kwx3GnXwK/v4leI1UWCg4hS+ROs4+ojsOiILlw6q3w2rctfp
479v/xRfiz1kfrKu3cM1kIP0yFPMtgM7fbb6YafLg/3dkSQrWT2NVP+zDYWMHii4
izlZdGQ3jT1H+mcc5QZ6Gs5yflRsvJkQhgpT89rAuKK9Xky7uwcqoN0NI/SXMOyi
94Xu0rnBsaexggckZhpYdJxArOeewSUIDm16SGMiH4IeOFisOrtXcOg+nMkNrqST
1fjLKAkBy6Nm8VpcQ8fAU63V6e2a4Zk3U1iCk96pKRys/9DVJ7IFkkCB7r4ts2YX
rMDjJODpHNvl4ZVPpr1CY1T+EomuUddKBaHElmS/5yXx54cMBB/jlEFhTxXyPgcr
bi6TVWHrAFVNYxeouKRh3RYnmCfPlOalY2/b3E2aI5O8RQPnu1Fdi1R82lEIMAbI
eKuwTQDjpY0xGyDypy9G/oDn0+BrX9mLu9s9GeVlfz6wmYr1c53lk0q+VfzZo7Kg
SI52yS+NWkeV6/ujYEH0C+rZZUsTVWwBxilht1jJSIKjoeyHaXgAjlihS0MlQODK
vOovU78QxezlEu5yuJ7P56CFsQjSRh0nWRstg08C3sfU7lLu+d3MMi0ob0eZfLl1
x3GgOs4rcLDRERx7T0max4TAOb+rPhQHv9oJkYfpj+f61YG3gdpZoUyxYGetHPwY
M9s2jExx3vC/43glReDF1FNkEiCq1Fo34brBKNENq1ZizR+GpydLavfiZBHMV43p
sclKh0R7M9jDYU/4ceXbYJR4vOj+fMrzE50dZcw22YRlYmGXmybyZenJK55w6tG2
4o1V63fj5QFG1v9PbBZ8AGwxuP6990XSGt9WXzs7jog/rCkFYwixyyLCjIU1LD8r
4aIeauk9OpSw4qs0RdfoVLm6Ymt9jK0mOEGYiqPG9PP8Xqw4W8j2TL5w33dmmrZd
VEKndQ1dCZ+QD9wV10nbV9z/fsirZiJi8gTq+GPcNx5SJ7Dfz8yUCAQiy4CyTQcR
C4m7JK7Aw263O7lH1oaoSmG/rrG+5+5c3TZplxGjU4/j/ePlsttZtYv5N7UxSpvN
lqaicq+26E3mNx6qWYBgmqac0DGyaCyH5YHUGPXuTE6RH5QAefGL/3R9JxLSqjJb
poXq2x2VKTOJWILaUure3KwqBPVfm3NgZ0twAvEPCC8rYxraKUoV33fGK+BJY/2E
WcH35oU4kq/6rNDQoFIig/pwL/H26nzxV9c404JaUPo1/zbWJmZAuWf71xcz0wlq
DFZy3C3zLHrP7Id2UEbGGnfQxn4bUMIvMe8JYUwRAEuam88ZJvglFbMYQF9p+7WV
bWvl1bDqda5f3TWapXtLHSl9S/FBP+Dmm/wDvVh36tg6A5Y3fIkq3VCiDWgoC9Zh
k6/WVwdcKK9XqPvapIVUealfZmEri/TpziuiTONe3+CKURbE+vcETTwqAfF8CXax
6h2n8NzrjpMiIfVSnLPEudhH/gpBCmKzHPi6tm6IdsakiIQjJyqY69cmAOdSDIC4
7Wve9rGPHZGYkzbctHFSP5tApvQZ9Z6DLyv803xdJdr9blOHQsdHfkBGjsxNH3Wa
5baQSxIGjKvXRl7hORVHwMllHyT4XrMvkEPwQgDi+ljVBNJpS1Wc3ra9OWykhRLU
yXq0iAKRSj3OXUf4AO424wzVHask7LAgSJlHMnZsJlZXty7CqO53A6lCbbU0h+hV
FxSNVCFFw7o98+Ld4pgcT5SL8vxmTTF7OEFMsiB2g1vuAOMvsfSa1Nr2eK1lfU/K
0/B+2dEXDwK681Eya5QfBo4ccgOUK9rLmdI9L3EeAQiEetPOfPldjX3oQMRcImpI
SjtmfYBSBXvbbP0hyVqQ3sE13YrA2LkrDBGuIprli15XVbhrFYwgf2p2BioM5KsE
1YlU8j5GPcYB1dyGi0V1/O7Zox5pvBkYS1g5O6Wi1rMPF5+WKuEPateY/DP8RyIw
YW1FFVXbQut6/6Aq7MCdI3QnniyskCF0+fo16cySFR/h4EIT3qSK7E1LWFYqHY1I
speTHlF33C9CMQ4o9rwp12F24cwxWPKCXBnkFxtv1k0KqBqk8epL+aycqvd8pWRo
Seb0o0NUivtjM/hiyuN6WZUqffTiNyyPpSbjHDTuLvypUZIXV4eZfCxTZ6wy/c1d
WenOOL2FRaekawAiHXmY+wNUzRLglqacJJwRMp4Sw7z2eZ1IXWGCvlvTrp4jfdBq
qhxvXJKeohlIQ+oy7G7temJZucd58Gs/0GbVloCoJjwkjIJzdd9yMtNAuNiQU9pI
OkXLO+nzWROwcFB9c9lvgYJeAublkfsFb4b/UBvXW04yI1u/HEIdsmRNOGyIusGg
kIT+l401Ro2lZGTxzZE3a9bmvIZfndg5Fo8Du3YhROo/iVosLTHIzj4Z1V2xsynC
0CvH/CVPLAtDxVwzy3zA9kgNTXSFNoUeV8dSAmzyh34oDnfzs5iuCixp201hJM+9
+JfItUHBT+7joEtAC7LTHKWKBdCJtQGlPevwxuJAnM5mKd/cpJZmmdzfamzcJq/w
70pcm14voVjcdfqe43V//Hp5ipynDg6yTgRSLu7tMuCjfUX4tJP0soMGBLLBlVz3
SPVp9bk8x9YXO28RaeGm2C6FqfjHlLN4zF/jYDA/vEtGf3zB5YIRY5BTfAePEsXV
Pl4bwAB+jHzVOT7Cb6HAhLCLWIRZaPeA9CIE2XIIZn733sP1ke1BMPbz/gXcsd5D
JXsxObecJzRjF7krPujBuTxuY0T9cnv1YZxpW57s9cpbvFcan4gbDF2Ih+5n6ywN
GG1nbR/TSDeD8SjKjEynndpbjlmim13osHrxBG8t3CLpVF+oemltOFJ73/GGVWGN
2HWDskz9QYc88f4KxS9kvYeis/wGFH/eQ5jYr7baplmXvlpenfHBeIp5pptNQd8A
EOfjArxpd0DtumN1UEhWrZXGUbm2OxhNLfSSGcD8++y1uYWIZSME0Q/kQdQlZeVt
n7C6I5AQAxQRg+IvCl3uFsfc2VG0063XG8PSTskFukUL7SsRG5QTSNsNcZCVA9g/
2xkioKzuGMHDIpgRxMuBOAzXQZ2Uw0o8Cg2HKFKbUT5r3tYYFLr8EgEdcKwzU8FK
jJTOziPtxqyFjpFvMEo23VZeTrXU2XDuynezvi4fFr5apq4ma/qDvojbGeQA1/Ht
mrJzJc9CvcDSqkTd3L3PrRxZj3Js+ltaHqd3cEYpvL/uH9NQEPe+HSE/NbsD7evW
iEtKe7b7e4eQ8Q1hOwuXNLPFDY+4On67xFSaPAi+M51yBh9lUs606bzehFZk2ePS
sTSLtzdUlb1fwmL2Ql4Sg+korLUDJG/gForhwhJwPAPvXMDzc551iibNTUukPQRm
utMPZyQwIdiod0TUgpe3ot95POUIUZCzm6fzfTYLlHxGEl9NMoS7pf/7/NNTTzR+
ER8vvtHz8bmN+mr7H96iMvQL0NeAYMWknXYM/9ALCZE/gGWAG6HPJlfufPtzC6m/
25wl7VmKa2GcTw5kKnClcMPma/POt467u479GMqjyu67zmVsRbZESVU6brQvVhpE
l4l8gl/xasANg9EwyEGM35GEKJUCg4Uc1n+9HnrNeur6+p/2OSvvVkrTg1HflhgU
pQ+5ZoTa45SB2Nmstx1EIGHwa5iQ56Fs8n4LVFJU7ESh6HbTBkkFIJqBRzWqmnXi
/hAygp+nL4tjmwRqCVXTh6wR3SALyTLkDO0KzV+9QPiH7URuJWKkz+jCPZcMkU4a
65B+gI87/PNdCQFvuY36CzKmg/j/XGujxFZxQYNIXafQOo8I7pIQZ9glu0DNzefP
2ElGomLO8Qf2SDxvAGuFgtBgzWhKKVH0uXw4CB1/XUO3SKprTJZ4G8VOBx/fVwvE
VS3fY4iTJRnvwsRjUtP0bbVm2bVrTxDPVFRXq3WCUZ6tJif3UDkmlPLNazz5gscE
fHNySxc3+Q0k6CdHzWie48298S3l7vh2OzdIw2UurPKMnhFzIub88+dy5Jok5Yq3
QM9zx8rVIvjibAeqUkBvDIGODgrk+X4uBXd3kF2of30XNDn3HHltSnTl9xraO963
G6O7iitL6W3VryUht/JyOLVLW6V8V17WHB/LLDXkpApACGmHQ8TW9aVGO9Fs4pXR
eQ++9Y0KCpRviu9REpt5Ouve3ys2eD5I2PxD7uqiT62KKLirJT0VllaPXh3fGnmV
R/jcbAuWRZC6IGzomdJnsNy3mKZg3S76hACy2mABO643tuthVxMTKxCTwQMuh/iG
RT8uF+ixPlhbOrwAgFPFlop5JXM+OfxDms9IBmVfknxhRiiAxXUXSM5/aA/Ipxm/
V50pMjih7yLys1xTUtke5qfsJbbInqB0xqzwA/TEIG9W9F1+rgw/Ly8ND0fpA3pC
lE9UgWfkDsfnW9Eq/FH6MpZvfaqdo1Zq3lGuDDerIgMwC5q5XF80FlYqXVBC7QUi
gTyEZrBHDbyqWVptvmy8/T0xW815xtCmZZPx4IEHsQCq0pvUYOFbQQzk2lmqrvDA
20x1rQHZsL80lEdwAoL9dTg9ANDcv11B73JvIPx/hTzESKuVMb//ZDZ+3PVrLP56
nf6rLv8pSlN9T5KPgrXpit5DVFJW6fIDTvz5gyAMPPmkyUk3gcfTBSwiIANo1ZDZ
FJSKQ3dsQYTVb0jj7ZqGVDxG6gieszxdwIJ6UkvQoECfE3DhV//W8/7DW1tikb/P
yQUB0UyrTjwhCrg0a8lrHfe6zalg6Bmr2UlBpM/+abwTJ7rVP+aKvwEFKGoIUjF3
2BgGpqwBME5guG3TiVj4TRkKR/pJsQFcd53yKnYxhsaoRef2W7HlRbpbEJV8zDkN
+L4c3gKPWI/vUNZX4qB3r/8qVsNqayw6Ye+Yfq0uO9R3cVR7pt/oN2S6YOqdijfG
R2Kz2VZBeKa6gxx2O/uy1iW++QTfE2CPyYklfgGzKJPPVix6aoGBLs8/VQwbZLC/
SpJHx15CWGwwJcGjGD7B+Umt8GmRteyFVvckGWJe+rtvvHPqQXMYvwnaUw0gebos
FSSUB5hlIBK09lMvqaCSRkkEIzoS4CDuixfqnpBtLFuWhSLCklLqUt3Qify1lyT/
SlkagtPcuyLcOB63l3xqjMfgZt6oCK3fzVoQdY1dHBLIDc6zC0dxlun2cikFnF6q
kxCYP7GuxrbmKReuMrTEuSMorSO8NuS3b3RZ4W59msUzUWQAzdC/bp8wfELYRrRq
awNLcHYADIx1VJZ91PqE1mbmz5aZu+PxxQNHaKJohrlnI68ztVXhPNmjAV6//Bez
CpiRNkF6AvDpyDWSKgFp9LQ2GP0SZy0GyY7hZc/lVJQhO/nJqjJ+mAizi8krP/39
ldjhQYICsOTdy0Fn+q/eIw6uN/ZmFyev+XsVzuY9bMRpLha9ZRQ5KO4eBQKw5/yo
nBomw3g/PS2rkdxHxmE13p4bgqjkf39yJaWrGZlzxtAmQa7irSfIeOs25LoVkFOr
Bu+3nPQakeVhVfOFvGVNmdXnfegkVlNmjZ+NoqtHzK3tcn8PizJ6g0pbW+Ty3ZAA
FwpO+ZxXEQLxTeAQNPgNWizLJrgtP+UruqtJWxnt2Vtn+9cjOcnI8BfhvzBsTwP0
6U+HnRIY4hj1ojnpDxAzVp9YZrVLdqnKul+TClWjKYrD71OKM+4/wynHfPOHmCpF
cruukVFmxRfOMWxbFK/F4V6PIE2u0T4FmBWr+bkHFRm+NW7E6aG90axfaTxY3gEp
RfTk0ENI91v/Z3AL4GUgA+9XM68oHihgl1Vip8izTvt3ZiRnC/It81z/e4dg3m9p
ulPGktuTFpkzHCK5Bl0+MqlKEHo8qsf0/49o+1xWBulSPQxDMREVL6osQWNFvQ+W
lKY6THkbNeFf12EmpEeyfbU3Rqmwc4bzkZWkmNiTEZY1ryQTj6veWa3ju4iAT2tL
cC3DE7z/1MrWxWvIOTpFIDEC+tixzXh+FQeJQydgSweR0mIdZDMWCQCLg4k+5fEC
7KZYqcmy1oZ0MNKrKd6UvQfAHYv+Tg/py+nZZpi+NvSLU9Mlxv5RmEqugYjVpr51
Z/WaB97QaqU56mXmZLdPEOTMokjOWxEWstcgSnb2Guvbn2EPSR841WeEIfuKdjZF
M+pTpmbRDJ25qzYA1+RjQMXzfkjZZvf68emati4i3kLDt2C2njLZPSgkXel8UagD
8qUKZQ74bhGlrldop8WU8E0KABNwVi5d+yoE2iubn3o0g05JiIPsPLPNi9QqA+7K
Hv8/ZxOT5l6nv2qUr+e/zkHlgB2CmHzWbVSLj4prMmNIDmmNXCYoXUk1jilXt5Xq
lLJ0dJrePU2hX1mY2DT969iEbij0WaAinkodfrMkxByk2ml2YFrjvBPYPbtAZcI2
ZPDiQOmo3O0iSBhP9+l6VWT3ZQfTFB1fidlVxEjj1kn5Ix+fdVu+GP9Oec0Om0xA
4GU1piP4/3vksbbbG8PvuzTkdVQw7yIQ4EYZG/AItfmGCw0YDVykEThE3IPr1gJx
DKorr3mkbUMf40gVrqKwXicPb7pfNj2QZk6Hz6DG3xqLSbUHbx+ZqONPIKVq3BjS
IU3IKsV9hVPTKNp5BlPkXt5Bkzlgqc+vAjcn+3FlYMTJhY9hZJcVHQ5dCMSihJiI
FI4yxy5XlLFjH+6l2HNGlbWOmOp5/ZdbKnx9xUs5SmfHN+meucsCMwUEJMt2a5SZ
Ev1B32tMFC+GfvTIA9GgLMhmQU618rI6xzz4ha4lrM9KyfPOhIkQRtPXlcFCzdfu
Icr3UpUtZFGf1GiXAzhgUJ6ayH6gq72SmJlBhtISWW1DjLC69yvJ0asdeQkMdtI4
C+IJgld/qIqlQNlWM86A1BYACzhq86igrf/lv7K7LfeW7UyRpjGxxqVrha9yxAlj
WJse2oJIBVWwHu/WLVfLHgOzkrYg5B6zgLF+O1eGFH4VOJ2EfkT2Slgjuni2gWER
ASYU9/Drm5oKRDhi1gUH1YThGeYHw/TdLgOGzn2YAc86treAxGx6lxBb5W61Rfig
QX3hf768o3mvhTCNYd9xNJ3XQa5eXSdfekEAnM8D10YeLLQN/9t1l7ezGRLF4eh1
ATzzFtx4dAvhWsx929L7C5paQcNTTIeGtF5jRyGIEQq+gjrOfeHb/HzA1DrmXYCp
clprKqL0AdVi9qrAPUKN4yJPjslP53sbns6WYE+8QcINqAKlgyXZAfcApAJ2JCCa
QIx/2uwao9meUtHAs2Xq6/KYjK/6skUCVNWrNxj7ACPl4oi0BwYorSK6LdkpaEEf
cBfNrxukHJ4YPzeNfV4AtQc9A96ocFUA8bc+VNt/6ZAiFVxOmbPRPUWYWSPHorP9
bHE0NBwcoycd0+QYjwgY+YY/4jkkh7WhwXDbI1m0I7uw4P20Du/4IBNas1MBQitj
nO3JlxorSmjsxsckIbaaIVzgeNvOcrsx4a7Kr4dT5OIQ+ShK6fNqA5oP9byxC3yG
PUhwNYQMBZpzbDU5fYz3lgW3HxYRETxxKNNOIFvAAsqWmWVKLmlofIFmu4LbIHMM
ocLVanBq3BmCe8YVtF46a0JMBCfweEj8dZdIZQcWoPocVHMgcONeQt3eJX9VlF7T
pBx9/Jr/rg2qBJ6w3nMOyFM9CIxPvTvyexJZiUY9f3FYB5/tmQ9hm1ASJ8hG9rlJ
0RAg/CZovdmHoEMn32gFsDiinwGp2NCHn6x2fObUIFL2TclHPjNdSSBgmpl3nAeB
CGndj7DaZhlOgmgzrnR+wYT8x5058oFKy2yZ8eIHSSbKaajxdL1zFoR3DZ2J4/dk
l/TFoJochN9fK3h26tRrGt62lWj52dpGlnRKIvj/IpTHgUjwfD9rtMPKVycsHAb4
YtsBds8tvwFYT5/j0bUQeusrLoCF6TwTHzt15ZXn7WiOKm715fGjqXEhPNuhzC1z
TKjktEBAq5o7Z+JU9j1VxL+EZ+dhJxAL5y7TrfrFIAunsytBXyADFePo8RjTbjak
EyN2QnUjMbTx+Dr3vvp+HiLEd1jYx6W4Yx5BH3PP5B9apk2pR6YJBAj1BTI9D9KG
mqtNqxq7IElfC1CG/U+Y4C65j9fZTxZGbcSEBumKih63lNJ1ZaEGSt9fwjd2S8IU
2ehSOvaL5jfy9hQFTZcE+pUcVPqrD9GVr+8T0iOMBSy2MXP1fszbqf7T5rrcXsfY
1QoncPL22w5whqoDzCVdB+PmVxRasTa1yNVMrEDHkgdeHGcBqJGk+I/EOxnlE37n
l8rXNzRSLZ+7kcrjQ1Ab9KvxfFDm8/IrUGK2BL4C+iEskNshrTK8arco/uAQlHQW
lgzgihT36vWXLsNrVr1ZdlHzRv5yjJghONHJVYmtuOa0xF7nsokfrmIC5103Qalx
0VIGI6MYlG3FSxzHneX66hVTr/MDx2HKXSe3ksbFBXgZKeLjoPWh+S7i94Hm8P2L
nN4KAd238Wi43iKxj3+pW645TBiKD4bcbh4XE/l0vXQY2y4b7gji+qEhQ9HLIkjS
/55IlBNsiKezMLS2WLLMEMYzb4jUNihlDMlwwyvj25k3kl5hVe5qekrgWNSfbyu0
6zIxYnjFrLHMLiIlduly5SopqPd8nsat51p3Cnyj61ZM8HpK9FnR9pxmVdm+XzIw
865fPJ2qQgiTLJJcFYFdwFxFXgUoRUqNBQSreNZjUmVPe2XM+xzfH4ZAgN7b9k0I
fHZhV5FZjqGx2dPZSosymR1QjebMrO0uchWgcTMT6gcpF5GRyABNGh6E6cVb4OnD
DP+tQZSM5XXiDs5KFOV3XzlrNm0OiadC8+jrg9lsOlqGUCRQsJcctHEdgQ4gsfky
Pjm0+BjR64lSk3P1a1Q19bJYdqeN+pXxDxuPFT6OSVGRKQQloYhKWgn4CPYc8k53
13Kq9fJS1no50yShvdL0X7G8t+uw40EARoT8/NBcwtcW+oBhC4X9d9CC6uyHBHcy
Xeze8KWWX2cDvXKKcBCpB6nIfekYR4vZLZ5pdAjQzjVnOP6n2MaCHGaJkSX0Hp35
dUV8X2TU/W7t8gedJTirBoieOKjHKombMscJWKyuhl5OHcIsxPmxnsjKA2ZdMh/z
DdZu+7kqDikO7IoQJTpZY6U+0TeXgSQ88T5+K0jcvXsmVJOHK67M9EFWqvUzIuNw
xQkLGdG6Z+0aWO+MaI1j/Sln2gH7yiPSVtl5TIq4X8zZLMZjeXluRHJr0J4nL6+o
EofcIeH2wRWCdZi7wBBXI64CmwxDhRiLm55PO01f3jNRY7DVfMRFjtkWa6GQ2O5r
yKSAKb7isFX2gp2MKq2J5ot0FisDi+Aquw/YHv1UiI6KMARnyZwvHTkmLTuNJoyh
+hs0c6+CRg8f4yl6tiS6sS1f7oDVdgkcvybCYqbpgfPEdP3gskc3ErG1DvEvEiub
SWW4QII9Utj5+Oto0bH9aMUgPFavtdBa//A8jp2noSpXxJ6tKTA3BvhP+al3zdFk
IGjxX5KI8XOBLQ9exjvL5uEgGpZZSIHiWEfOpzvofqc7H8GpLG7MAK+iallfg/xP
uFE+RwSLWp8DJwKdeozoBn5aIqdIzJP/C3g0MEpmz6pqm0qDonMSWhKs0cloTL9x
pO/qdlQjrMdFLxxCi918fL5NmA1I133X40CKOrRP763BjGHkEJl2Mh60nMBj8miB
8813C+AaiumCmuW5S87SgP4U6SZGeFKm+7a1SmrpJBAnJn67yylpjC3sYq8NOVRH
s3E2A3BFBFE94kWp5g4aDr9GqhbNqOtOksEx6/wbSk7xG9vaZsG+t910cGBG8w9v
kT8QrABoUchZVEllcKef+lHBu7AYaAK0ok7gXyTPJ+WFXkHMgFmPGLj/vPsHF519
c4T8EN7T6bWA+jdrvN7FR922jIs0hf1tnVj0vbtyPFZDgqj18tKQG1fTwKK4b62L
qp9sqMbWnDdBwKdpVIBUIXMUL/ydVopDCMmN6yii3mVNT93pqNigsBKGnnIszVWy
AwNVm2oKYqRDcYqaHoEXZVi6+x3dohBy7Ouh2KuwdhvB/L3s3EJllAB+GrG60q0+
Ea2izK1bp1FwQUUzLsyZfUCn6uVtHq1ymfPC7d48U75TCYWvlqy7ZpFvbDLRkHYq
uxvO7IliYU22iPKAwgxQO9Ir9s/iaUSV03E5AddCroonFqun2i2uyZYeeAVaKayo
hF9kK2o1zALtDG4NJ0KQJ6vWTeo8uKxO7zh2aXxSUhyFXKCFo0Z4x6Sfisx/5z53
bN8sJdnQAi1vmX7+LSO3bf9qhvWyPdRsSlR9dOjGF3wJGDSZqIwXzt5BMHmJs3Ok
R6A+xEQptbB5kw7pVi53dmJQki5kRH12O3yiEg4c+9ZsS83YHgOtpk9ez/topEfb
Jfbycyfas8yDY3TjDd082rdhWJYf1QTeu94QFCW/F+ZbaQdjTvMh6w6wUdVxuq76
Xnf8ieSApr2HXRyI0FQYgMwrocbtAol921jM44VafMimx6lNvcUq6F8KbYfHY5EI
SFW5UMxBYzbUT4SacAHfld74l36EMsqZiTxLFpkA0M0a2jCsHhI42AZ/YlHmJPlc
1QvLD1S789GI/NVKzrdU7z12/vePB6loOmmbW0t/cfIRw/rEiDxgAXHie7/RfnZp
Fy/D7rLAG2cW72verke38ARkp/4H81CoVyAkJ5FrWU4yAJ4HOXV6Rjs5kspRGiL/
XKNK8NcsKO7r7c/AFYgLXGREUIq3gpEWnCc0GMGaaw/TG+V+clEZbDN3oty7fxPX
3zlSFWu3Dj61/U6XmjWyPt2ApZydxXZa/CEDTB+ABvdcg5GrXNUACA2WARDWuc7s
2H4u5EYoBrNglqfSwLW7nyAV2PbmX9GDEVIB5Z65WFU7OtTT9xLKDqb09fQcLSHl
QQwObp3U+lsUaLzukyr/PudtQ+Yil+3vpJv12vxtSXzWWsBu+AWautm3wSvonAwk
auIot//Lh7lctlDiT9R03dF7f3MkxI/bKB0UgvsOGbFWtAMOY+lPNLP0Sl/JoSPG
4pQPUvC1NMyyzRNZ3oFqL4GlDVwjuAp/xKvYy4raDtcuO9wngTQKXAD9CxV6LnVQ
HLfOGwv6pk7uuizvpl8tt7mz9wRGhYt716wWE0Y0rQXpbW+/C3IelLerbIa58C3B
QGRwDBqhR0+GQfzSnKIdruGp2j7iywflZCoP6L7Bm6cIdumSRS0Shn8T++qH5L3Q
nzgPF47ky2Z61iM0PaoKbMfvA4j5piNgRFIn1QaAhx08JKPfjuncje5HK/OZb52w
ReNhShMExTXxgS6PZbiS6rMDX+qigsDhoHvr1ptOjS0n43lNl3+te/q85H6qhEjc
D1q6D5PNN8Y/MlBuRZpgCdzPUPY0zDjdLEs29mSV6syWfJSL+Ev8htzCrSCmD2b4
0kTgpCsi0kKeOq7KWYqEyGFEKCwWyahsy7KOfuZ8b+CAFq/JZIh3FUpQDBFJBGie
7wKVTTCdggOs7RtU2FquyPbFXGoKTZdRIJW0Lqi5ZQRr+02fEJh510C5Ob5dQjdf
vt+9lBOdPNQbIRMuaN8NNI75TWimCn3jZ/BhoKvlJuR5xwqZowNWuB3nN5ElpQQN
+Tf88/p25cLh3mGl16lil7o8znFO45SPPKwPgHxa3PHB34X3tjUrMTdd5EJsxyHk
rQF6Abm2ZBZGAZQKE1ZLk13mR+E0Tpqvly7HhAdqmPAu5mChQHIAXRun6zLJg0bb
YkFRQo3qfpqzevCqxxB8U+JFuk6YNSR3XIZJMo7J3Wec3bJW8+gOsqeOjKJ2OYO4
gBs68r44wmUjlOPUjm62dl6TYUIzjAkPReJj3I6UxgC8sTxejsph+XEFYIRyGzqW
D+v4FHWnX34VrKVZpAVX7EXt9z8uX+7s7Wb7+ZRaAlXId6yduSo4uHBpu9JWWRii
3qLQqQoHNSs66UNTgth6uylYO9cxcLRTT8D+EGdeH9vuoMlSV8Eocd3RuOlk3A+J
KyoyUdGyJqrRyb6HOyiliGSUoZXQqU7jxFUc41O5811nM1kD1JYh3Q+xtgUgx/XJ
BUqQPamCu95Kv8BgRWtXNj/8nlZrRTl69XBS8sxcXFct7nqrfpTIBAgjLI3hr+Vu
78bdUL9AFV03hnJK3zMjE69ZEuM3AcvQuzvBuVKoyOpV0qDUQYnlTizRh2YQw+VG
cywyr9csx9qbVx5fLMIoBFqHHC3U04unOQEI7PYeCpE+YArfmhOt49Pj07e9ZC/r
1Cq0Y24IhC/0rLMSKI5hYcRA+LK5DtuJC8O8aR43EQdg7ZiD1gadX31Y/QtYpO0H
sc7zN8l3SKDSXnQ8KeeFROyE6mM/liVpYV0tgGdV50P40yXON9dLRIYy0V/1u610
EsOCBQkt/u1gLyKmtXQb59jB7mIutmkEccpGBVPy6GySS43jCEvWblcGL2EZY2oe
Yu040synjxtM8zitA5I/MgjGDsJOMoGWmiB/u04M1W3X+LpgcNb6+3UUOzsnJ6p3
w8xxh5UjL6oJBhYlerWO7d/7ytGB91G3M9wfOfCIwCLPoR7VXJ1xjEA2++F/kGed
2DEJSzSBRC3SjSY4d9fzmqkXfX0JxdMU4UkjKutLEv7Pd+nqu6Ab81ihz+3yg+U4
nvLq4Hsbq1qv+MOHLsv746k/zviOalzCf6p22M5Kf63YOSxjhFuId5qrO3No1cne
l9WxaZCcI8ydGqYeFSpGpbHnI4qoXn1Fwk4lR/kJLlethT+eeI+nfNyOHn9ljGOE
q9WdpLYFLz+sRQj+neOIA25KWoMY9Vq2nsM3hYJdclSsyINZbpgPEicOV96SK7h/
pqwqS7G+i0BwasOlJ5DLz6cYRuHau7w5on0Toap0V5ui7VZ4FBRO+Aq08JFiqjXJ
jeirX2hWuCPwST6XXYEOitoLBZbIVo+2vi/SBU79LSCYOLS34zU7PhRw9zoP/K8U
4HPzdX2s63gw4SHBZgu1GH3k5oCR2nq8Qvo21X/5RBJp2a4I9Dx/2IZEgLDLulWE
Nl/uJUj7EHxNjLx0KB/hpxQ6Fzn2V89o+9QNZBNWvbLAoZC+BblDbbW9UJTct3N5
iTpzSvCBT4Gv9bFM5beW4xyzeS7qwdi6YGMi1u2WyDPWhg++hlXL50zqMNCgUkqG
+qb9TUhk2+KaJPXlM3P7WAW4vlkiez4PRsyhCgxSOrb7LJSzh9Y1/LbblzSJ5ydM
g6oE123zu79kYztRPlVvdqjh6CTgtH9p2PI8QrMdbp1xOLzF9zutxS0ThBN7nNIT
ppY/toFBqhAoglgK1aVf4g0DJZzn5ULZcKhuLfrUrj4u/X0mnmN7eUtNfne/dU9C
qNfUFY7B1gZEIfy1vtXZUQGDFuv3X0bquMXWWNMZuTGXiQfllJdU1ljdKt1A4Ang
dKW+5DCEfi+gVeiqGofRDJLOg2LqOslBMppCgHLcko4vJxGLvfnGUUfgGb2KaIwa
pnmLSBuJNPx5FE+JC5+0R7BM37spDxFFBuYL8lwmKzN/Md0fZBtUPBbqEbBqf0qn
qRU5JdPWJ5xJqin3ZTgPCkHk1a5A5RFvRiPxEFJQsp5cLz1LGC4FNglVvxC9Lnuh
Qlt+8cfA4RnZr7aeUpRoPY2jsnpj2/inrLpPIsm0wZ53Lx8vY5iEY9DeU8AQyrLp
xGUtwmilFeqDFFHnq/tc1K56of5SY4TszCEzjtQLtQrmiM2Mh4PXgPCjdO8e1Qki
/nLWpxj7SJeB87snDr99v8+Sr7SO6UpBuhoPOfJIj37qY8DlunfsvUsK6ec+vx47
8ZSVD93ESIDrrJ2NQQ1lSUo2ZCoq6fv4G3SGEWvPXWJuu/9VsrRWkmJ/JX9Nlepw
uzh4r+Y4HDYh4cboYWiWFVBliTXh4fONS2YxNVz3whw7sLq9hVXmbHGK0dGFfIwA
S+xCdt8uPCuNS7DQZhXBwTuoTaxCUPvzWYaZL2Qmb+vUOlzZlxClyy5xoGuKUU6k
0iLjs8WMKahJ+VdbhqY2+fZVEsuY1SYH2pjPmDX1qyt8YjEHkQWOKBfO9S1b+x6j
XjxO6E/rdS5xKMUqJXkqMn6393WcR+gAgdfnKYbGvXcUpHYDYgMC+IbNOyfwlXuU
R2s3GTMBm7EcikzlN2+I9LJLMwVrLcRKFxEFg7W3h1+UA/XcuN25xPgGmkoSJQ6g
ZLqoZVpHQwZ4Qlxa5E8Ru+4DhBiomPurC280tLVOyCsxuW4GVlvpM5dgy8Pb35GC
Qest4lGOnTD24RvvFXVZn+iLk0dXeYWnDwBoTP+OZbDoXOAQAOdf0BzVSx+sUjLm
YCv/8p0MRwczuxOLPi0O8OZFKb9iBz3yp+PCOat27pMo0J8Ecp9FyQpXxkW2vUGJ
LNYN5AgmIAIYFglelf0/jhXT2ggNWAyHoItjiGrCuPUcAcLYf6JxssAEfhmjHdX9
Q+p7DZt6dZI2Th54SLEVVdficljAzOY88CJswfxixSrGIC0QuixhFTH4+a3o1oqi
w4ceU8vYRvKxrLECvFREJt6aMaPGRg/sP8qJXjjGnIhcXtQV21fMoay0y6k7azp9
nGvdxDPutmST3jTuHxvtGzQEe1JJndycttvgYjtZk09i+hvS1xame3v917MxuMFM
YNPHpAQTSQ0EZb4rhg7NCUxYIyxkom60D2UGwjfOpeahq4gCsf1T227ye2GrVb4K
HtKUkQxKsKYxHlWiUaeH98DgYUnOoQQf5VGCGSpOYXbt/jbzmqwG8XGSpf1nerBd
YPrNNNau7qHAfCYBGpYKUjmT+fjycjIH1UtOmCPRoP8I9H13czOJ/1Wx5i90woyf
OM3HEQ7Vn3nplCBOdfu+s3d6CP4hJdZVkzFaTXWKtInbDI5u7lLDewE6Bvt51Glp
gCd4c3xUUY4rVK/qlaDgXdakhrO2y1lTDFHOxk8LvpohuAcRG5/sUvnQPMOQB1OX
dkNXm96LZwDnf9zlfPJxm1x4FlZJF6+JftAYGJJ4GQle2+uMT25OBLP0tuUN+B3e
Mh2Gj6GOlkYT+VSMLaa1rm9fe5W/eb0cxuhmZBrXFzuCN53HEoqwq25mIUTEZU59
KxrFzDP+AV8WdKp7xgZ3hWdBcQwlFW8wzApJ9ERErUQdGTBpyXkcmLvC6Fw25uX1
NqJd8dUJT8vJGuOMTCKwQ4+1r517wGqMLlKQy2C5nyHe6YGxNa/soen5qSUwT1G4
+nyPZO1jZLG4gHGFCNfCyvGNZYYv7Dks4A60fogIESPYWXlBOCjjYyA4lY7y5iez
hiSl5qrHslxm8E1p/XPyBSGRY6nluv3SRt/t/cR4PYG6sbT0Fsej/qbX0XlMcmHh
TxwPDKwpmqkvyZjCjnMDDMLXmLE/Cqv0y5HF3CpU3cj0abGgV2dj1LA9t3I9bF1p
wPqN+xd+eW0N3v0f3FxtvL3YRotfUAdSv0aYBcTyeGDeuSFZNng58ONxrwpJlZx0
niBychdaVEkWgGpRUULpUmVNOaTeFRuctmoYF25p7FLnh0HzLqhOegBIhdu1O2YH
tbkgx2794byQGIAS22T8Igo9Hn3FKWBR04/hQcARrYYa6Q2fatgwDjDIy0v1Bnid
WyYPbS8kIjxqA+hxTZzdrWkJA3PlYzNPsQUe13gngmPCWFdLrPSEpfZu5cLXg6NX
MNevPz2vE1bPithgDLZRRR039Ed9Uhl5mZHeiAVq+cOZCqXyoDjkoYj5W57Uuix7
b7oK/H2/KJdsh/y1HlaK9U27Uau7l9pU7KgT4LAwAY4uJNcyl1tAx3J/IF9QaoR8
u1l329kOxMtwEH2wUVpBOTX5RmtFMrMhoQBQncd/86VWDSItp5a+b1yCId/GzRlq
b6ZpY3dwOhFRl/AHG4Tr5RiSx6FxSiPSJotd61sNbrvJN+NetPkmzOQdXoxtwLup
xDvgJrSXOI15KcTBRdeo8dCBAFaHOzmmstFgK7CbS2yfuGeEIys9UKwsOzkWZURc
BvWNTFsjIRqn30rVQoGvnoYHN/dJ+KVgP0duyue48dZb9WzSoznVe8t7DYKqFiL8
SMZgVOm0hX8agda68+lNr2r/nmbE1zzx56ibvzjpa8W57hKYTbSHZa3vNWsfFcxJ
FOeVZVm6Pd21AlfKjAKZ9PYuiJG/PDzc3rssCCx+qYeQU+HGzQjzNlWQscWoyZWG
va39bVVqTQq3srbMQSndz9400x0dxDdupM7pQQSJ7LSsnPLcJ8H5ft2FEKpEiD7Q
uAcZyUSF6Jf+TgZMQKeg7LWA9OWebDjPsdLKfnI4ISAZvWKrrO0pSrVrdquioEon
wU5s8aHEWIplkVvVoSjIX/6YWQbR+BvAQ1DIhk4MtY5BzwOIlBoQsXQTRrRfQQ2f
2rP32t5+ULIDjKb7580jiaCYo3ANz6dzT+D+REeBk6/nAJ/aKWjoiLuN1CPFrCO3
xepxDWCgpCvuwjRdR4yDa3n51Xlf3kyBCQSr4fr++XOlqg9QnBqZ5AxQrkMWl67A
/PWo6czdERZFgytvQTIyZXLcXt0qwndLce73c0C11JK5bNj4oOQy7zF/oLbzyW9T
MQj0pUZ+j+3lATLvleehsN5hmoyl0MQob1gMK2tkUb5jfeRhn3s0a0GzpZZUOloq
8A84di8UBMLelvsMMAlUyPrNwgIO1O7PB2VJFRu9ZFUzjSEdoLmwiJ9pkOMXpmE7
18ReslDjkWoAQdO5mk1jdPUhxrg+VWjKZ4vex+O6zNWMaotNi0WO6BM/0kKQNITJ
LxPjfmZgmfhIEegHT/+dbJOha/p558QkFPBgD8cr1nrMLV7lN1hiuwXPjczDMLKc
kngXeL4eSrNzvMW0XJf5NJxraV438eVfF0oTuifjUtEDJG4Erpd5Bt7kpDzoTy4f
u25Q7Ftp5tjF0CzA9oMPXLxSFzCRfu0BWtcMclS6JQ1QR3hJE28xQYvXNyAl4Bay
VPzo/XV0OOoyKkIYiFFOHe7Evt/ujSYrmryJE5vDeAa8IHLeRAprsIF/TSF95ey+
S8XkSPhZKA6EuHdmcygkp9PuB5UqOleOcqjnNRUA4yTXab4EFa8nrjPUXZzDeeYE
dQOePwxARtQUDRCY7nuaIXOI0wC83hvlPc16nT5j9HtqQWQj5A/H+fkgkVl4yIyC
fAJEW/qVImsXR3lEyskB3Udx18syMj2VRXGfit6kJWbuqiIkZ11PvTqmIMnkURAc
Nn+RV78mltWEoJhRcd9owhVACJ59skxKEUBDNQbKv7ctBKnRN56Q5JZEoxKOxgcW
JS8M3Gg30tcMuphnQhGNgqiqKbmG8UKYNCG2DRkNgxWeKaMcSJJUxtrykvnLLuqx
FoiJc/auos5MQ5vjgSg1Q4Wnp8OjKZOirr5OXUiWhIxEAqZjb7XH7rCGM24MylMm
F3RDlGj8G1xXdUlMKVTKc8XOwjJzAA1/Brs0U/2SEotMZbPkS6W7OI7uO07bJDoH
SbMEdyxqkPDj8xnhz/9Y+UdHoJMHvI+Z6azp0uiVdgAqrfjRFZ/CqkNHYeXGQMpl
bPjCqvKrndv06BtNGgsBv/BSQ+fWxQj62x4ZUbE8HsQQe+OZhgsf3Q5V63h4N7qa
sQc6ruLCuo6XrdRyJSw3kH35PG7k2OKIUOt9gq+mzFHl7foZnTrpoNg/DVG2Lubp
fY1celbmPuYln4VPX9/+ZVF3DjOv3xbii99VTcvm8S7gxmRG0UlMZs5kjLs3hlnY
ZUQCCCTLtOiO4IXpP5Uq95Y0tz7BizlbqAEu98SmgFJgML93IFxAS1Ng6d5xBV8n
VylhSxVcX8SuYclCIRsxGxLTQr0HQUAwlHM1UTqxG0e4U9Vj3PjCz6UF/TKOFJ2O
AO3D+b5hpeA+KXZtiUggMCnd9AakD4Ip3vkebiOiMEvjZWP6APezeJzpxtd6a1FM
ltCZgFkj20pN2tEuvRFT0x4mVGz2RddiaqyZHJcLcfcpm7XEQ/rtolh/gOV6cf/n
DTT9clvr9/ugvO/a97atd/1+1kXWQUDxaeejkfIcmdJ04b/t5wdrWMmm71sHlgFF
QDoIUbc4L3Kc0zZTcEgFtAAfh7EAbqFBFQU5tqM93o8sX0QOTvmkmOZrHdB6Q6WW
9/E8X3iEPmVRKpbsZo2QepeeYTgfVp6Plj8eATql10i7sh14gyChCDkYBgJ6PBs8
bnZPKanOQzCXeD/xVuVFRBlN6k8IebkuxlEIpO9jR+FIaVIFCtiNkh900y9B7RNr
aD8LLyUCgYbUFUfuG4snWuGcfS2Y26CVoOG1aXtp/8aCYtB8lWkH/tn+K/+geYGX
2JBspfMbZmDttk264zXJHJdbiiv2LWZLwVZpv2dPbe2PGyoTM7Kxz5w2HxX8XCk3
SEds/0C4O0kk66aLWgwDmdV0bdB2WcxqIQ28xYOje2tSCoWvmuRYgHIbV4t/VxhU
kRuhDPwftmp4awvnGQ5u3kgYZjZUP6cHsdjXFrWzK7vK8gsOMm9GACvgfGiTUq/1
g1DGdGGD1TsIR41XmnZtBCJyJxXdkcxtuZlPvgJ9HKoJ1YdoCM7HLokGYolbkSVV
K8Q2ity6pGCHc8tcVdh831sIc54zLJUDxWtqNSqYal9YusDmuyPTK6xTMjnYmAc7
vFT3f1RqBxu5KNbHI0MwiuoTYKfU+GKkTQj8/b3lJmWEV8MqDgTyEdsjdlwxdB0T
KrPYlhTBufvwpx5c/fKZgdS6u00057ZjTNGNFniyv3r2fOOvBnoMNIObJJFcdcWr
OiWJnfBV2viBTJB7bC72ETyRC8ONgdPDhr7evJ2a3ao/7h0gOxANUM2H1kyR64K7
w1PZ8QVDwnyF6RpWZIaMMqtStatNw5XeHs+tN9PGJIFZmvx+OaQZMbZBEKPm3GlS
JRq1UWtGXDccRN1GqTXu1LeDQTHYkuppIGmVoLo0pl1dfAI2t1mdADfZ6tw0aZGj
oZBavXjRTOPhG4e1Cl+NhRia4jwVA2zRnVRzYYQwjc0m2o9uMAHguuCFDhMU4DUf
oaTEV81cfY59KjFAABmr77+Y+6BFVaMS/xNeQhxI6ipiHdxJGgVEoD2miug8MEyJ
N4m4x3ySe0ZKOsK5UL3A2G78VXx/cLuW7TD8qRzD4Vpgkfsgg2WWBBw6EKzs/qvi
NLxg3/XyunbflcDLSAwGMrYqisO8gHnzBUQ7xd30oJ1kUCG9nFzIoOpzDnRmhtun
3LCLb7tKU6Adh48a9DVYX63OpVkT08hUzbIohmdy5SpSiiMLvpkiz/nMdUcLUbuF
3pVvCacyh7r011Lqa8zQRtFVUMdwuuD9vhnGrqG6sGO4LkJxdNd64/4bSarj3Zpb
gE6/4J8WcDNRafCdSkLa54EAQ2YLqiY+86M/SqUMp++t0/EFPpzIrJpTcXjtuyUO
xNgS38H0llb1AzKEAzlduoKmiklhgGzkC9FPJoq05WdGDBV772S1+8j68ARIKTga
C36cp/Sri2T2vV+jL94NFnQFMg5RY64ZWJYhjlpR7lXU5jcde9cXn5OlW6EY9WZK
+oaNE9f4v27PUCcKHGqE7ZtsT0sn0JKmnfsxy72GFv15vcRBARXBRtKvIgMZVKjU
0Ew4u2KgvcUmLPyean2AXbGDTWJpX/ch6atjz7Von5cVE0HFm7hR1MuZx2mlisEt
4Ks1xDQ2hBfXTzjua6SypGnyi3mND4GypWCed63fWoRF41QrdTJ9USdHV7s3G1P4
N4sBiOGCMDZEmFs+wkctZ53iFBvfGroBFEc1PzzQimyuPvBs/2IW6GUZjgbB9Vws
Ay3fU2rVbnZS+dchWSCNxWh8/a6iCLDXWq+TMalTo8aIjMKuvSajTeE18CignYsd
LNcxpmGxOjPPMS8VL371BzjvcB3rYBfIUkrOF24j882xxyqqHl/NuPDjmh1ukLMV
VWUeUtBIK5pbcX8Pd87IXef8idQqQbUHiVYAEL5RIO0kKN/3xkAMRlBfswFAYB0V
DiKEZIpLdhFwbeY2pVjogCxfUgtQZs1MPRqTQmtyRLMJZGl6Oe1vCGnVnFO4bU89
2B3xdEBl95WJrFOdQOpYVJwUFH4NqbrvCxbjLd3tNkxvHwmeYhCoD1sbIbrmnJA6
robcuf2LuowyxqxICwueRkDFI4UCYmE2ZJn/7azKznGgGBszQ5nrE0plXOJAfPTJ
GRtr8qWGTtw9MqX0i0OOmXQrNceuWq1e1fwembT8H2klIIvSlIn/kQsuouIiaNV+
vncC3dNWct/dtAqJ1V90uwFW9DBUOncoIDVpKBvRFunmUvIAMXUlP5mssc9HRTZx
OvB9gBeOk87pK4fnonNKM+IRkcmlqkIxtCKcWQ4U8WX5sznXDHdQqcNmfLlbpQ+f
I0Dk65f/gVazG6LVPWUs9XpcxokE9h9U27ilHtIZkGnKwdpTLMnK3yCYOW0rByRd
IwDt4cIS+aNfqKOiI/0+QCS3O1TOJGS9DOscTVfEYWXK1+9UWGQLhNuKDLIXcviL
JuIXiEer4lD/XeiHkUlnCGIjfBAUx/guHiPZjs8Iklu13k9FTBsWdxvRHfAeJ2la
ZrYvDZffDTJyZivwXXKM40C/YIOrHz2qRaSzZ0WoSNj44gtSz2Xv0JN5o3XDSAX9
wMrd2ZIh8hpQZer+s3Q3HBE6SrRK5LHsce/3sO6hJf8GlmFM/Huv1pbTZBg2lb8X
hyA30QeK00xKzvANeq9niwdX8XI68pWHsW0o3keHfqaigkiIJG0Uxx1b6w5PSDTF
sZamhzT+OSrZZCGLXlfbIqZii0neBJJ7XTrTwGJWS6YT9k+ZUpvyrMN749miwlro
1gz3Fduw8sUgZdG8b+KhZHHAiKDw6XuoNFJlVaOQCtTjXk6FpDzWhGKk/DxO6Vg0
MOvbCtYocL7sBOhwAeYviA3Ph9cFuFw83xzMlWqqoJGgMyzWctqd3n0Wtj2Yu3iy
ukHicRgkvlnCnQYJYuGlrorXuRHXmZVwAQy5Yxwu8P/vYzZ/vpd3cbpe/2xdltlG
6jVhPSSJ+zjVdTirIjjMPYhi1PINhmK2sZ5fVyOf8tL3aZ7JkiottBFSBXjV1Mkj
vxaGysx7k8GssLOgqXZucd9+UvkZyQdYfkMt2nKYZh5JYUvYWh8Hy15NBTkLoLRn
t1rubMG9xK0sy8kOmiWsT0NP+NJSR2jhxCXc3h8r+EDGwBldQzcaKViwzgUhVXyG
ft61j3pNdO/xULaCfgjPJF9tIHk5j+MH7drlDgeSSK1qRtbHuo1Sk1nbEeoQM2Ol
sj61gF+mVoNw6uwpaxe7NlN+a1x3VNsiNNDgtceAzzKApaSegPOBrYe7PUBkpR0v
tWw0QcUKXhq/Do0rmhhZ3VLVPj6dCrqXZws7+K0jrL26Erxj6JDy7eaJ2LC2EsyB
0nqp7MTGji29/cj+PiP+fMit34EJVUjgbYxk2G+ZFNZvWlVRKveA1LqTF+U1ELot
yVY3eVYbtlnelfjo6qbVGmqyf5RGdSc4mHame8UVsIXqGB+X3UL/bgt7V+k2BFwy
B8Y9oh56AfETuVeZQ5ldO68yzFpESxqzAEmAfybtz+0rIfxZH9t2unaVva3KOgkp
DhdHnSbno45ytLJz/eHzC4i03X4F8ZT3RKj0oXlb0w1cBMXY+PW3dpkC0Xgl8+wN
pgw+sB6jWGrxS9VkrSJtm2770vqIncf9HFkqJ+tK2GiA8tWkrweGmFKcW5zlN+46
vL7+G4b/bbTu6BPe0yuRiUdc3cAG9cVnVpq1R1GZPEFBxXCiqEGWq9tv4lwojF94
EkmU4fn8BfVw9O6KF5it860VsLWUKyZJFvW15X3m5PkASJXI/useT3nBESqxGs4f
pUUKLyDsKO90wvq1KMDW6XdFRAWA8hIYPyJwd9yLkIPto4k0E3X4leszlncZe6A+
srnCvftUb73mdPKB0xFSf8IuF+Ps4ZXJLKA0POV0qWe4rcH6hYjP9ntlNvIqf9Zg
PWqWL8bFVklGCVx6AA4nDbtuvQ7pvBbBHIBzBZGhDSFgnr2BfuCoqc3mLIsahHF+
JAU9AoHPAB9uULWR0fWOKiQAmKOphCxCMdk7eCcrfn0NWAgUnmjszVnr4qUKgURz
33eGteShME4v1JBllhwE1TL2CFg+cZaLvRID4Fum/s6hTP2GYWr3xqCMn9RJ2j2l
I0iw02xWgxnoe/ovo2gAaivCuwRzuXqNxO44U6MTkrVdn6CSYVnNVvS7S4/i47zg
cO4VrsTDpguQZgCsjmpZcfh6RT0IF5kWsfIo/yHLW6WIxGtiHZ5AMIw3cWXxjKZZ
U9qZngVfmSJlx9BxZE5CfUFZhp6CVxSncBtWZHhWJrSUNElkSvDOqx8AwQFUckSi
fm6gKgta3CZSHcdS4/OQJpivPk9gmUG7Wz7lRk/3NhCMdVx2OAqpPO6ubJBmYLR/
JfRB6GT0JwRSboSLMeLlg5Q+BTgxBygprAnoYKfxZZnQLSm0d/EnLN/ip/Ozrjbr
CXpA4Ywh78R9e4N/fXO4ZsfaFBgWILZDLQeHJcJRtroj+wOOq1p4E+Fn40Y+ZyVM
41zf1unoZIsfDLILhjkceMH8PJ8h1u1iOe/cks0yJZxYCfxTokbWU0cfL4KtY0eI
VvczJMt7mi2ltk6DUcVq10DZ52pHyVmENapaSNFTPcjwb+X+cbVxYO1mUfXMraEs
vLGEgY7PQP9xg+0M+u+7b84OIIi/3Abk8riqPQ4QwfsyzR0JpNWOJASJp8bEo77A
oroIx7axBXWbyPizzYSLTfdyvRcgror9TkhYZ9SwNhqwqeY2UNI+Y5ASusHqDN1U
GraVvgLp2Wq3M2m8gyfH39TDPHH+TQJoOF0BVnNqqJOZ33cfKAzy141V7dKgaItw
UlzgrQmGR5geYqSs9NHGf7hyvIFQD/4mVPBBwPpMh/0OXdd6b+L2BIhyEzOLLhUZ
ag+ALFzj24nbQ8zuCSVPJT5CpCttKjmF0t85tal3b1II8nsefTCHLzFO21loBxTa
ADoL1eHDXxXGPzH1grYqRXb9whczQeCHR9fqP5VRBA0ikYi5YlKObp4246sqI1je
eRbnWNKj6wm/v0TnCh4vBuvWTYTa0iKtvgeNEvJGe6/1QtL+rowTgqNVe0XZJu0I
BrDbFAhntat9zCxkyzilrbChzA4vDEjLS423fnZFt4HSrxhux5JGpvR2o/5FIHvO
D0Bz/Ji+FRVKVhkI1TeY61VjezrgWX6p8Durzyir3SPLbdPKYaEeMXqDX1UViyJg
j9f/Egy7Nx95vWlWU1U5Mgd8XWampzg8NMPG1D7LEEpERncTEV/3ZGAhufHan7vJ
xDGAY9GmR0ZRveHieKJea2E/e1u/te5jtFmhEyqfBx8bTf/xD49qevW4u/y4ry4E
fB3fxaf9f5uukA+dMYxB4GddtPmi9akhRecelvhPtUdi3xohxeBadeNNM3WwIybh
xaMvYSTAqwAqAwbbv6VdlQ3CkAeNpdBNY21raWaRPDiruB3SuUiMom0pVZpiIGqu
Vt4cfOy1AoaP3kscpqcwJrK6mjieUjojJyULCGevMm0inzvDAG3MmPBUFJ2hYey+
9g1ywXUf7YrwScXH3Ema1xCZYQtLZ/4BNWUS9n+KoaYYDAo0pIZ/Mj0Q7IiyS1Kv
deA2A9Nq/oMrV1QxcY4Rk/4Cw+YKgkM1JC6I5n1DAt5/g2fOIJyfCgOOjgdyA+zr
qcPa65YECYJLvPxYl5BbeAaMprsCg2h43cOzybiu+RphZ+bk8ZuQU3DcViVZSgx5
UGDk6mSvEfKqlmYqUwPeanmpF1RHxG+KhcevgrXW1iSoAZttxsXHe6nz9uUYlYZF
4qogXFSyjVoE4KGQYAZDfcQOtx5nfzoTwcmM8tbjUDiKKVWvYqtUB4tA4vJzT91c
PxckDFcIipW5Z5F6SRrvibuxnn7ym8xBHJoFQzAWQKU3iHdLVIqYVMyX6a8Gbqh7
I5bZvSNtAdpSdJSpqcygDMWTbVPwjiuGqo9Xn80y78c7QL9BeZI3QCv3AlMck/Sm
ZMUSLxG8Wa6m0ve5awzgockPCssMDpCpwdXoYspnRrY2CcBmZTXN6Q3V1rMB0ltd
8wO7uKPzl9rGQJ2rM8tCYdD2JyXqfErhSOnw8NZUojYWiqAaxWK9BDdUgZLu/1Wj
lIttwpurIuDd3SsHqmp+XOEDENIzF5P9DBj/mpk2on1e5z8i0dsOE/1RB2NOgqjg
lniyBzlma0Y/DXTHAuHfTrmqWlDvfK7FT1hgLyXqJkR0Vr6LKpE3/xEio9J9BgbH
DA3Zb7x3J/zG+yloaoR7WMoU0M7fVs3Vyx1TXO76HNnOPHrYsonNaKoKAEZ5NQfR
69eJPUwIcLZsY61N8zu1y9fn07QdK0X5wnDPhWjCSABxUeG+rbyNWico85vxbHJM
UlW1mk7LQmB7Gd3grndcmOvYIiI6lKwXqVNWpvjy97eGVuVT43Wp9so43ZUnB9cA
NjpwE3ndwthoMcfHwHp872XhCZUl+q6teB6O6sSv+qNP9CvYKdpTlVMG0OMFM2/e
gafu1xKd24EtPREoK9DA8Gj9xgrFi+u2BaH57uX5s5eVysiWmG2oVeMYBgc9s02H
/ulJEO3Qw2B4RUiTcn2ARxaAcA4LiDNsjXpXR4G3OqtZ/ZXVtcGSVUmyTC/42kO5
vghzFjZVgnuYWJr8lwakxT9LxREBzLT8bvD19WqXWEJ+Hzpqyi+U0jis4epB/dd6
W8ngINGXNQBWxk7wM0/acy86XOzNGhngWXpdmu2hSBgwInqMQ/Yd4LVPwKQEGfXp
+xdrVA+woIRmyFpX3clto7HQpVLdjI1Pd3Ls1blW/qPrD3Z3diZNpD7Yk96X3hBk
DtBFEBKgS16BzZZ7yssKlxzlvaEoXB5Y6lQ5LWSwJ+AGyf2JOWL5DmYYbtE4CoVO
CvYf6Miz2GI8vARbm1HinG8Q5nM3Pm76iQYuVEcKnvMzCT+L4MFsSRYbK9tkZh+z
tj7rcAjil9TXstiKHuxf6Tooklfbh8MUg/dIX0C+pyKs01MfSXigBFtHrsC3QUQC
BvnA2cS9x68UJsbTW1OIUFJlDC3evqdLIo8NJw5B6oaS7/68wnj8DMPx4wUPkxIc
s9rZHj9L2I2NkgtCkVzW2cEjtG6jPrZH9+0wyD1Yvq9P2DgImLjAiG2v/hyJ/7kO
OY8MOwanZsmEhh2WCzIy99ka8ueJG8kij/0x14las83td7582wLsdy/keMTkVW6M
C5wBCV4G/qN6Ncsn2liM+PHuYjFHwsFGJyXJNYudSd9roBeJXHcCo42LHeVKQpA3
oPj0fRlvN1Z6G/gG0QM+XKE6FjJDc40S+V+t1gozqdfTf9BVAcMNnhXdILQcSu59
cj/UPLRE61zA4JuCuWfvdgtFmTP8w2yzd54m13d2nkElNwArX4lhmWNyLF8ROw3r
kjPFKLw3HG8HJGJWTm5ef5kKWM5pNLv61Y/4khoyX8PQ0mVGa9YD3NKuPTDCwYaN
CR62BuQd0EY38SRvF8qfP7BGEZQ4LG0LFOPnbY1rWnYg+K7vOwKRTFTZqbzNvMXF
qQAlbIyJFwg2jg/vKm1BdyuBVi28s0UZXXHq07NCOywcxmU8jsr279fCXUoIvK9f
HJOX+67FWS/WFMVZDZ0v+gfMHmykFGPKZB6Fb8IFID9s3NcJ628Gt1Uj4Z5wmTl9
9NOq885a6ow1AEgJRrKCFNFWb7zJpLAWfiugAF1IKU+UKOQ4TEFvAMsC4UUS/Asq
A+98DUoDB6MaR+XB+kxch8aG9j70JnxtfetOdStsDblSq1KA2KHdh8ShnaCDk1MX
DxsaIiaRVlcnuV7w+98eASBlBRxs4n85Kd0XfLsauuyJy1+cEH5ix3Exz0J7FZc1
IcYPSHaAr/mWHdRcnGpNTNmjGmHCisqx9+LM8joXigcZua2Veoxb/iF4HA5/o4xT
/zF5hG/M5rq0fZRNVHzr/4Cs5Go2pPHD/YN94O1MXsnbtO85FjIwJzyhFuK2NwaU
ZlBlA9J/w2n/SOHGNcJVDAdYfnFGS+BJ1bU1hiBnHPs1zc4ZhvxpCIDrALyjyOwO
862sTUqGigY2JP2ZcHWDw/Z96rWMrQXUMKvvaRfzc8yuVm0GPxvMV5CCUi6U7zJc
yN+wBbwPDT8XKWRAlO0lz0SwAVoS4I5EFYPgIdN4R35cb7OzUOVqsG0G+xAp6Mr/
90gwkBNYnm3Ch30CG47B4SqAKxnf+towY1h89Hrybw81n/jpSpQhzhJTNZjC21qS
v8Xy41begAVKBGzYsNrCwxHgCH5g1ndvFZrPngktGLlmAcKi25KttLS0H75GNgj7
CAoqD7jeWBLkFI/T4Mxd4sqPsclD6M+xxtccuji9lhagQrf/Umy+aghB/fOieS9q
5xYXHDmC3k9lH+OrJbhEJQkkekRSZw7LLcIJE5Oq02nIjxEzdOd/z4M9/z/UH22V
7NhPLSggBPmZJ8X3irPUfnhhBw23LI3m2+Jl4tA1zFIw3JuDx7zkJSzSsZ1n7SHF
qevUN1/22kWpRJ/ZLay4go1YRhJ2KRnIn8YuPCxCnLPjMwJV4anu9UmXIVtqHdiA
zjo6t/ACbELJsN5M0OhTbZTGszNPGoMFTywDLHSiDB3gqeozCU1yJ6DINy2HJ7zr
FaNt1Qe8ZqaGfVM5Fszfw1Uhio0il9IZyU6PJUcMCMspROKDc4VXDn9fiW1NBeYS
onwX2ZTyrQt5e8WMO3HjDwgF9QBnuoUogFQqjwJ9JXgZ7zBsGOyKcAz6HXLxD49w
qeGzJO6+M1ftSnyBcC4VlSwRGIVWfOukEW3wyWIu+3mH3cFpJ/slMBpgX8aHmZo+
Jj1u2gf3/rRI6NhD3FrGL+Umi7uGyl0uAURCkuF4pk9w+/GWQr8ckmv4NJG+/e2H
cf+Uh4ovnmRdu6JV2evdUZov8x3qCIAchfC0Z1zeXyTK3aQ5jWzN8nuW8lRwJ12q
n2Vgk31yZNV1e9Kl1sU10xK+ZlyzINF5eZpLiF1drSvCjItdUNW8KTxHwNPuAshr
Ze1s12TW3IQ7ZnOyu5NtaucMPcIwZ7Dlfj4q3AMlyaKlvJE5JEWue24U1r33pkX4
K/aqMZ2S3PouZTPOGvTo9phIlth8jaCu6KnnqdAMGzTSD23lVQbFeh6IUTTsb8OD
U9bwgjOxmy0HMtV6LA7/H8c6MhumKQwQ6Kw4PfptMHeZkhDRtX1fti3c/RXAPirb
3LYq7Xb4rogVnJjINP4AvrterT0rWi94ZLa9ATLGpZvIdDB+3ZcVKW3ZBinvzXPt
XOsbkHva/VE0Z7qOP/g2xcaFEmTeGpeQqLBjojy0BUNeE11VA75Zmi1z/BOwesb5
OJvmRVZc8NJ3zg8DeRoLdAckXPSllX10Tg+5BaklvijpGUq/3wOQx5x0Dh4t7U5G
hU64JEc2O9Kpzd9YhcYXi+iiASpbsjAcvvgZrrmPqVw+BvQZVafBb7X76xQ5tkLo
+dybLpAHsUhUVaZwavwirseScY+WgTpAfezZ0Ue3a8woG9+/kG8dlgI2ucRt9YNP
Pw8595+tgAIhz9ov2RKg8BW1OEnfv7qnlN0Vzm8n5fIBLWKoZ+6IZXfk7kAvo67S
lAyQs8ilexlm6WiHi6fGIOc1iwIbSCjMeaTntN4R9cb71g9oDX+p9L/tQt6z99Ie
CLg4d/K5hfuNW07zP3WWip+Y1QLvzdo2o8GcSKMg2fkKtrLrlJEx6IGvF6Ne5d3P
0iLVjS7p7oApb+DzRIDZEzmti2Hn+dZrM0HNVGDnkxfWOc+7b0J4C6odCEXa4bv3
501pHA+s+Qf/jbiNKCslh+LIXA+EnGGsYj1tUOBkrLzXNwdjdQscIiXsg7lYz+v4
ZkSaxbi/YEOPYlfkWF5f5ZupFLAooiPuMxNEEhqsiAuYqtVjbKYqZTbs/Nh/Nhw9
semng69nf011QQim1xSpn0cuPyV1dhCez/ZpAGG5MfavEWKy7xwfj16oY62lQZgC
R5i39P6O8w63JPAIQXmEoY0TIZgkvIhtS6T+uey2unqu6zUexF8ASheLzwMrP0gb
eIK8wz1QJ/0RIONPICD7lN8fMLLov+0QNMRNyf4ll03P32cD0oE5CFzvACYHIpu9
0UM+8YEDH6n4Vsp+01tiQkrx6W92/2FF5LRp/tTQMayoIGixxKRDfXOXgfEyBFD8
H/NmF9kC9sabtJs1bGWCkc89x3jQrWPqQg7Rk/d+dq+CrzCBkPjCoJn44xHFptoz
S+7Uz+zPhauQr4gqMjDB5AT8RxVeGVeYJozrtXP+sAHtQxLVzeKvLLE51lvR6SGw
V2S+M+L614m7VU67YuewSywo8n9ArmmT+WiZE7MHs1YpjpJmiC9eXwolqTDVnGNX
EAXWZO0GFhQRqI86nFsJv5Ds14UcsKbxowPWsdMYrx+Kom8996yMblKgM5D0xWEO
o78Wraj4zL3tN8f+n5/eSrIcMtebx2V81n9RDtQDs+vPxKFkDxniaCXn+XOZISpn
1pRi5Y3FoTk0RhLIjS2lU5huuj+mRn9aLCa87wTSnIQrhpJobcSA3ZLTRTsMRB3d
ZVJBmvqG8PKFDuYdQlbt7KzM+vm42rbqOKnEA6K0YzlstfM1gYb9WRa7F28tADvq
yBEZiyqO2Sj5eLScMGuj+tCCdAbv/pxXCclnzxwoH5QX6A9POSNAuOX+oSK/pqzi
sgAktKn+DsfX0mdvx/sMmI+noasdrQFzk0msdkQ06D0KiVEXhxtx7Y6gLKFNoeaE
ikvkJp1mih6UbSRy05k8rHZJV3oOY2ZlEv3wpOGD0/kXuCI7bWi8oB7LoZR/4Yb/
ohgh+PSiNkv7RFu5Gi1oiG9KGyGB7bW9V3I+z0Q1iX8y1SPbQWkliqFY52dt11NW
zEQBuGrurxDS5nJon9Grc2zorQgZK2/XmWoadkcl8jdpfNFZE/bhOgtFHO6ShyiR
Y1UViXuzIIVgE5so5jIJsf/XTytWx1KQLKjD6GMCMCan2grvSEql+YHfFVa5GI0Q
biwAVRTdgivJ0nvfm/OLWkjuZ5btJOSZxgFQJCzCN+4U3et0P5Cy0Q7cfoONGlv5
zMxsHZtxbo+WvgsV+wPgEEN2qQNT+SOjW2Vg9GB72ruJ3NGBjhGz4xJ9G8cB6Vti
bFbZSlPXcQOFyXtYbMkVavRP04cEnLfE9aA4HBuhWx+7h9N28x1x7s/b1izPYLdD
azru5AX0aCN3p1okyS02SfAxfoMoErejy6pa12RQU8hASW2T88RxNkUaeEQ3ab3y
hVpazwiJMlgyBvhnKd2Q5Nn7gbFcNbv4CQnJSfpjXyPkTkwOolw431JguA+9t8mT
UCqvJHob8/kuyOcQ0RsFgnU3dhB+ie1K6vKz0WhvMEw+PW0UOWoLA6EUYYxAbTHk
eOYNn6lQCKYhH1pTb0WwRzWs1NXxVnJgoP5a1DmkEMSSqIpsJlyFo85ECBBBZvXe
eIDWmxaYZhW6LDJn20wsLt5A9k9vW8GTlWI3d6nvluOkuHWWgR/eyZNGCH07k+Li
lgm068UUdvJQeYWOzESPJmS1GyPKiH1Oxnywerc+oEYC8KeRrzAUYN9qlzhcRoRG
xvVg+gYXGyKRi/XFfMwrwssRKSCza+ZwIcRdUNQXoVlaiLKahm6VnxEIvBb23PsT
KQvxP6o2FgwAD4Fi/mhW8f44FvPo0Lhq3TfyMIuSmFUq6c+k/MbbMNADXKncTeJg
CGbYpIwbzIMwqhF0AlKJQO+ALDxoTvL/n5w8UVF0xcx4M/TEm4pkVIAqcEWzrG4/
Jb/uGTXp00pK/56IV3HsCYrYpJ6+L88JfZhsBzNhtQ2ZP7ux+s7Af6/86NsdkDUE
/pHmXOnqAzQ4lF4Ta8KjZ9H7iiZ8yCO4ScXWkvN4SW6zd8/qLTE4QWr8UnOqwtPw
ZvJMULDXiytlLWhEpnjjeGpWm1jtEiKZwbq3RrKSC5ypPXTDTgnRne2/WA2p4os3
NmocLTByhB0DIsvgaVT43qjcOYnJJ4aN19Xm+Y+rg7geBVX0MbyxWokyKVVCdm1L
98P/Kbh5M62MCloXCHmh40ZUqYDLEZsBLw42WUruTQ4kFDf3m1/kmiak7Uywi/Oi
yK+MlSvlm+PeytaGNvSWTHf4j4vkSAtBuC8NA5t5TIWZfg5ZdyixO9HaudK/Kio1
6Mvqmy5/XLz71tvQ0VJ52A3p5GGaz7ETG2iy+an8sqPb/7qZpNnYlq1RpvAJ7RYY
CYtrSCZbSv/xc0ap9udXUcb2BokrCQanPSehszV+zRKDYXZRcvUyMe7DyB1PdJ1o
sqNDQFHYHS5XPKhOmSpjIMmPwjvpjB59UQLubEF+k2xSKT7cci/iMvYTnwrC1jIh
v9Mz/Siahoq/ln8uhaEUELFUQkxFbcnsoji72Awj9HgeCXPf/pfJrl4n2HCLkenI
B6IbxzaIsV5Jc4ORiNsAQbwN8r7tEhEsEbYTvuJhjruFns/EhbcsPPSHjEOIVs1c
L7WEiZR4/wZg8QCL/vfI6TMq7KBVV/sedPwhsmnDu2SFuDy7YU9Ki6EGiuUrSmA8
Lg56uHmGg3/m6Q1IkFmSeKy4OfnuZEKmp/3hC1jDtxV0xRz5GzZ3wP6t/hl/C3Q3
Izbu6gl/EI+4xWlqpGj+LkU2DZdRZPHSoGQR3eWqM6VAViV9HCNwITm3imLeIDhU
bujt3u6Wx1s0YL9IZKTKYPZ9R/fFnSzP1KUHQT3bvX3nxr1jKsnx2CdXnKGOg3fB
JZk7q0pgVM/EvCsjFEgeuZElTBAboRHgMxdyZleo81v4bdD5Emqj8JzXUjDE6pyD
jZ3dSjN5PwnCkjmhXYRhcGs2npYASmdhK0gu8yaCOAgLyywkxVnZBT1XhdIi9ehB
08httbuQnE6aMHQnLBACgi2vPwguWdsjIcrbeqr94+HuVUDWn0qrOthCxFgcPgER
f186IaVppa6XklJhfsjV660xDqCi12kA4JllxK9ZCzpo9/fZaaqaZlkcW7gNuRq5
4y8cPqA81s+zppRBcuQQauvvo/LkrT/RmpiHYC5Qjq9/R6lwPW1HXcwEjG9tMpru
0QZDxAp/GchMUOsG573hJ8mMElS/4MUV1z+6oIO06DK0VKwDBvy9/342h7EjxSBk
IR2X2+GaowN1oA0xOL154v/2ZjaLEro8GWkAK7tpWcgpgVo035ka+y/gkY6E0qUn
Isl0A3ENYo7jKS8Q4W5xtSFtcYl9ck64SMNWAHWkVyTO7hIQKuzraS64MZyL2lHs
MH1Gbtv5JMBVQatOVARcRXzn7QdAEXFIzihe3GculqVLljI8ZwECBGVQmru5vyyx
aOJRYRxnuaDtCboS61jnvvkvqEFWUHFZkWo6uZWyx9aFoYqPhfRGTUDIrb5tgb6a
5FFHCT3rA/S0VLYx6JchohoOvj67rM0Ml7mHR4A+ZW+76uwrf8IYxUWiCm2xVKsO
P/ceu/njatWjD7h+8pmhJYyf9W6C8A84ItpduLfR6o+on/7G1iUdawt0qkrOWlPz
3JG3TLuyJGwJ/CFepe3C4i3w+lH8MBojgEBk3IDEWGTIf9mqufH+3tIPoH/PkFbv
nMDTN4lc5Uc/AbCsl2UL+KBCKo41LQzd4Z5nKd0NVek7xB1+KNglXQ+cCNuQ5TwZ
GFnBVooMWVkj1uO7UdBpY24eXfANxN8F3kTudEDfNfJAf9BjPoIfQo7ff0CCPo0y
fqw3zVx3jygwsU2phtUBd5E27ho2WEMdJhNpfHYg6JoMZIMipDdloKUWl9II1qj5
0evEyzKqeWMXmqOymoBTKzVv3viEJeN9UTS1FCDJp1qh4XjH12BBwNobDu0w7P95
RvJpXQIaND+p0jth7YmKJEnLrCcpPX1FV9rjE1G9P7SVoaCyCunE04VLBp1Kf+hV
hZrP/g3AlOkdV1ui8wt4pLcTlWVFiQKQFNSbKBSBUWaX0E0FIHP/7sLwODXNAX8T
Ekg3kQkuXWkud7ji7e4k/phPxjWnyIykAMTg+5BlPaO01LjmTCRYPfwJW6dspjkq
GEwNyjYd/bOyfjmRKNEszdI1o99VplqZbsg/96paEqcIF5fNcv6HRts7VaS6gPUv
TGtY0J/MAAnurroiCtVmoCOQxevkyQW/aioFqjfUtmcG/EpPUT6UMCTi/HLoHnQb
+6xHsgiTVczSXI+qnES+L9MTCYFYE9+ovbUgJUbwAevk2tubxtq7ZKjgfswbU4/6
g3gGqgUZolaxO7DKFfb+9ldi6NR5kODiCrBGsiWaSV2PmmTPzDZvun9VD/wHk8mx
zq5Ed6yG+TYnndWWyL1UCz0xx7a34NMybWRggCn1UP4LfXYJgeW5kRgcQFyhB4uU
FYb/LxQe24KiwNEqeLcMHhnDrLwVdLHuskk5LmvaCiyw03ztSJvDUFkWklmjsNKK
9lZHPeep5SBbfsWmG+QsIPhyKmpNtaDgZJ0WZNvReKrWGAX4YSkw4du8vha90rTD
2349EIEcM5JuEC7l6ZtqXTd0YoI0w5/qOPiA43Xcr7txeATfklkLmBV3l5NyULxE
3xNhmLfHFlDmfBKBEKy9O4WXIXVDlT/k1i2tUHPMNtO/Q1SXBTD4AMRZOd4du1/j
uoV83fmow//m/T26eXNqNtvwydER66BdZPRCgXjqCHcPFUqibcvPDnEtybrsCGmd
Co+xgONEFVY7LHI1oPa4FfeaHwvZk924caO1EXWYrQa4pOTiRIgJMPkJ5dRaKrQC
chtUThhWMoB9ZlbnWajLPyGZp8AGb3b0YMEPSBKIYIcw5Cf4iKiPtcgi4/4r2jfi
+sh4YhAjqgeQbAF2dcLTMc+aIFQBgLBWKrdm4tIEYaV0pn+ZSMbNcxA+RnZ7iXtA
b9q98TEURh9btjMAnp67QpNmq/lDJxyyvrkimluHxrUtT9X1tPap2l9m6wQjj7SX
H/DIQ/UkaD1e/dffUU+CNWu6j+0/tne/nTXDH27BGbr4T/kwviI8xGmjkT4clvhG
6o70VTWSH/N9o3cqPCk10YQh/sVD+ggBZpf4UdsPog4QSyUjg4nzWmYTv44J9AFU
Avk+d9btdzTIrkBUVQy+ii8RuqdmH1JCtv2PCURlmaA4REckAqes+PpCT4U3Ninb
9letwy0qiOr82szxr3VLMo8VrYpg3M0Sxbz2YXfw5d3wpURHfduUhJjLc1eeWCBk
7WjTR15cT/Lh2bK22V7ZY6rnmAy1Q/I0TgsJGJOMOF/uX/zKfgbMLFd9Ivp63OJT
jon9vQFd19VAfkPvJoOtzFYmERhqhqKRILhOeVCsU4Ks5JHp8Ex/oE4p0xltp2a+
zACkMfQFCmy6OGDQdPJNfwbEKEjxaf2CyV2j6X4CDJ0nZTNU88lCnC9zmxro8PuA
zl2RwDBcNoUKUsiKhFcu6QaSs+NYWRQ60+uGSOQWY8HZtm62f2L6XrLk3lrkcPc/
E5y6KsUkmQlJbc7BYJo8aeykgdHkvhuYnmIlGM/4VEM362v74dTeJyqVQMrp7Q74
lQHDxK8l/pKnIcwn3j5R3zj44o6vgMDcOhGL6EsUiASZv58nlE/Cm4Ib5iwMT2OP
k9e6JFryQGgijLF8NasctrEdHRPNA9/LpDq2nhL5ZnrWdIXbWONag9oXxTNl9Ikl
yEVeTaHd8FWcPjcOoNCRlk269KU5F1HBdfn6iLGNFqLc+GhjMGQRktvacrEdZSAw
2gr/x9aUWD/tCxeAFC2bXEKMefX7ozK6ezcl7OUr652Co5U2U0X6Lb93va7j40Vm
xuLkjaQ6jBFJEFjbVHMUy2f2GdIMGmn0tNQ/6sAxLtO6G4YaeYWeK9Wfp0IaYH2K
wHdnbblVAYaFwkDNvBM6vW/wO8smkJ/JdWxHVWILtwvtwgn4hMCHux9uW4M3MqbY
/mRgQF/Np92hc4wTk3fAndiyLrN3IBcEsAos5muOTC1+Y71LmOsfJ7g1WolEKkpC
xNOA7Wl18Z1puVSyDnfpc60ggN8OA5qH7KqZp3F/6Gad/J6n0KgHJ0IyPA8fX08H
p9Hi1B/MH022uS/Vj0cVnnG39PVrxmHk1tv6ugcv8Yq3fDZLARRRWC4ACckc3C5j
6F+mbK42I5rgxCteg9HrpAWrjVuXoTjZ+OiWNsYUh6YR7C3C/kS4sZ8ntl2pJzGs
XKtK0kS0uZyq/SS7D6gq9u2ZkzspOA9wDwhG0F+mo+rypJ1VlrTLnNSsy2YkIwKV
w35R+uedO9arQsUCcdX5GNGxTlrGtuF83rjqph920P7VALkoZuCSfB6QwYYLgz4f
X45Ff5t2sZnnvpBiiqYnzskZvTh5pMrGF7/+ua1tLuNvibG/SE3cpj0Jeemgwlt9
m7zPxzDZeCSciZlNc5lRQZI7mOsgKCv26nJoKWwlVfDttYY5+VZ2CfCFqwjfAvLc
koFO/d9EOa6WGN+ayOJ+s+I7GEBfM4mxv1IxcFKAljhF7OriqF9Wi1g5b0Vh2fp5
s83/LDahlON8B1z3GsyZiOqB6rFZ0pCINbSnpZTIgTiWRaNeJwaWJ8/P6VFHGVcX
+yOXyvj0Ib0+/aGOoeUTaw6dhuOvfIw7ShJ6pUxmbh4fw4/llw7d0EJ3YCPQitqq
RSy55MpQr910ucKMw273vCOHSSpQwxbuK3qbSilPz8m2MRMRr9HUkFBJ5wP8vLM7
hr1kAqPVK3/u5BaGuWpibtJH4rzRWTzUD+q6jIgmPZ7sFoKDkNoOu5KLjMPR3wRs
i5RXtywKCDhwt6d1qU4YiNCxIjdYCtlo9AnI8meLJU1BpFlmvYcVlo9KELCflNHH
9mQkwRezt3hNZK8x2yfs/3Lj2uDPLK/X9TMYkkhzRplafBAq1b+UjZ+366SxFbnT
mi0Sq/wKz4fjNe2iUNPtbxUWSrwk5omeStPCRJ0QF7QwTyWeCKSVX6bZnHBQ3LwB
WOA9wCUbuYx9JPrZaQPx3Fm4t12JsNfh1qxFRu4wKaE0wN9OSHU0OLlZGJ+nQKuh
uFNvKvPQUkAsCkYra0Tv3bayaIyIBRpapaRt74eZzpTee0/76D3mkYKKajdtF+cl
ABsmv24aJYnuMzLn1sLv1Fox9FA0k5RTaL1WXWqdvDN9EiMe8x/SV2LFyu75E8tc
+sXlShFkhk/joQGempVBfYM303LEAZvxCKlRXnUkhUP76oFC+u8xMa2vkitV+KiG
gULh66MBHkKGKUt45sXhr2wG2akMD5QTG9TvOnYvMSBMR/M1oEQI5VfQjXRu6JKL
Wuq8qDB3qQDSH3rVTPiZSGZkRnhQOmaIXKX9OGzCTvNHF740M0cq45tM5emZcVym
/sMU/DOeGz5DbBbF3rgH8rx2K8JO9XwtaMyjspMxydNSGv5YFo1EOqgViIBox5vr
hXWyHsQKdEVLj19kexDO92spluXT+4oLmDkbuHR1hZRW+8j78fVIfsGccemzaHo8
h68WVgkmA9H3UG1Rl/x+UWtFOzKGIDRaw0EDc9towtPEpyc1GhIrPgEf/oW9mpB9
/MsXngTVukjUqaBUlUoW2KF6m/6hISnkvSvR2wZcIYT5699QmlyXg5YejBhquB9j
FGZ+lbg8PIHUm1EfBGBzQ6ZWV92XgWAdtT2nDqCaoHCc+RmN0Tx5Oj0zJeezLrxP
PROrq1c0uIOr4ZN5GB+cjzAMexH8jaiUwfHiX5ofHK+WqVqU1JiP/xMkXAhl6Rlm
Wsy2FD+eUVCup4V72B5shQeruBYQ1mUCB56EpdKNRvAAPH4vdLQaWhe7eFN6ezjf
SpCqpCJh0kcK99aq2VwwOJqKVYW1fw/6NrjYVvrhsvS6YbQPi5VvTnbkpY188J8A
PgMA2MoAKxtEH50YIVPGFP3Z3mDFwXmqVecUK1IrwX1QADvA9O/eSuzkCQcpp0lu
1vLEGX+GLR9fMI4RajfXrltDTh9eI47Sca3T6W7u/2YPkAXITRhmxepOO6Ov8A9o
+isv634espCOVSRqilSRA8jp1kW1o/FmZael9FRJn0E2iIOJaxsmL/opReMfpXQN
58kOjlZVBEXa3cSaQ/kGHki0sE8xf523Cqf6ydzO5D8pWP54rVeDMOplrPSraC7E
0tkWXPVIxi45lxQ3Ij5wz3lnglN92+J8/DK7X+mgPbPqi3S577kZrdJEC1IkUIMa
maL1o1bMJF5wKwJOvRevMgr3uSiy1Oi2xpkeESHH7kXCUJT2mYAbCSmm8UgpNsix
zloqVVMe+nbIDweOM9JzzFO/cFgVhznmy09XT1PY6P1DXK1wjOBb6vDnQPVamIcC
vzSzQxg87dLJQlThm1+XUlWYkxEVCFqN0EbfYOWOW+0utopxFoC7kBaDT0GwFfEn
CjNV4sI7ZEPMumQ8HQVd8F5StwQdoiZtrISitFz0P5B6kZMaMsCvDEPrV0svqPu2
VKMxm/88Dl9b3dbS/ynmKgTdHZyt4JT2TTNxOaX4P+5cYnjhXBRKqZm3j/lQAwGr
6+ALl76yq7WaQhJyWBe8r7Ql1rUdZQTFdGbaRoJp/WV5kDn0HZz5fIzk/oBdVVIc
A95PTYvDYukw21AXxBIOhzcy5udIGXB3DvpZHQonBl+xKsCZFuDBdOKIU1v90EBY
BcwBlcRaCpHiV6sUncPnaqc3+/fnwxIKlmkBuMGplvxvOyYk+OdQJyEGTxEatX3W
gs2RXl8LBWyCIZooxpmUjS3Pg67fRV3kQKu7nFxGf4Ns9mFjrjNMOdMeYHgl+G15
4zBLblqcYs69wrjBoLhOn4M4YfAxFgdlVikrcs+pTY5sKQePjOqJvKoX0pQNekbK
bA/ok/4L1THaYCK0qvgNdJb6QQUFNDV+LVjTA8f+gOeOzfbDMiq1TJcip8APSYXr
fdlXVnW0LVHI9Q0poSuY+s3nogLeVAzcKYUUgKi1Cr3FQkhJEbuwxJJKqzqXFgUd
6JibWcVPHEjOnE3H69xEr75t2kCIU817JrlwElYMbStNnNuRWy2VStcYFZik6erR
TvvZOccO54ux3H24zbrQ9MCZBver7f5XcDpL2Gm0JwMYIdyD35fa4luvLAvPiZoK
mfKP2+CgAd0M8seTFT7MhYfCnqSGWs0Oqa1GhGvdx9WsjXNkGrFCMiqLGaQ5lq4w
fWv3Esp3mhBX7/fAgi0NC/ETTBHmDx2fdF1gy8caWqhpZaEO5NIv0yFVSAgmtjBb
wuqmcqiAZ40XoTI+MACZyImNbmRrC1mNODVem8obwsBjgzwb9mV2epvQAI7XlDYM
+dVEyUZE8FA8Kl70TtVdJoOfmpjfTMyLmppukmahUM+4ckTAQTJqPLaK9sNqUWxq
nww6e4Pwnc+XTEcpAHMy0VkpG2RgHIRbOez9TCIvdJK6ZeRcmqTxAFmhGqRwPDFG
8huoeEcFy0QS7oDao9fc3VhRoFKcgQZDIjBhA2Qzsa9vaVKk5Unv64ScOko9On95
PdVj358GX4qr3W2Y58b/kp8aFiT0W/2eRk7d9YMNyKJNWp3VctoOHfaZw4MWwmf3
gVk5qFQPz1eVVewYnwfn/OUVZhJ0ihYJ95Tdx2DqJzZ224EOHlRUAM3YRi06Ke/i
9bIVxwNpLUSAK3vQAdi1Jr90RxgijjBx7tchFHpLfErFRaSHVTn9tYHYJpHJzOnb
xkkMXo+ssDBrM/lapN3L8lEeI6QnrQJebOopPiYvi0rnKgisiHiZCrkPMCUDNokr
IadOmdaFmht4HqpT02VDjY+rWBu6vFrRaH3ms2a9YvyuWUx970vTv6LfepUbLFaR
JAEbj279RVZ9s0IPDCONgtWsUym8MgqdkJBupVr1oGMG/2hZ5FKitd1z6pfhFgbi
LsM1FkjUJcRw+IXjZIf88Y4vP0m9/JR+SVqphUFaaWRhT8fMGzprPJ6Un/JEw9GR
3voMGyIo4X+47GuyAQliVEYDVb/1FCfpuM3dGZDleOqQKyA5/RISACUvK8YHcEPL
aSSxMEH5wpLYDrLdn7OCqImY+z8MgUYd/VAuj5Pf1J1ngNA1Glyg0JKQFzKPxEKZ
RIIlLBSiZsXw5tFtEifoW4xAM9ellOexPb702b6PwJKTeBzNpF/kzhc8qWn6wU6i
PnHmRJVwrCSj+cb9Uqaf5eGcmsbcShIxATPhlP6ohiDdmWVRLc/Ahhbg0KoG2hrf
ep2FtfMHV7wX5KphIt0La98fj1TowuTcyvCBQ2vY4okwitWUedQL36uCoqcVOdv5
SreXze/8sRTRYV1/+VNfdSRckKufvlVUPJXPPrFbJ4Mdh95fy0rjBUwN6HF8uWbm
JrHS08v4JnOqrWeTe3XbKlsvCd99cInQx9b7AD5z/OjjQZTjwyA6fX0EgmNVDy+4
TjBmIwBmCK44tRV9Ls/7oJoWg5tBlb3m5zehLvpUHAJdQ671FlK9NYgEfXcA9Nne
MrOMfYKoGZ6avfCKKu8iLIZzjIXA60lFQGUfLb3GrfJyZmh1+7bgNP62aBcNHsmU
N2QPKx1dcr7vA1law55J+w0YrVYmGdaexDbdHyvcN/1houSsVM2rmz8KTUmeUcwf
bVt7MUM8VhsnqE+E00o0m7IR2Ba5G3ChdCXIQjL4MLOhv8g8rzQHoZHZF8s3l933
+wVCxGh/0tZn4UbykQPh0qcPJBloYgB7g4oHxnUAGchf5XI1L5CpLqA743sJdsuU
A3v31ousUJbzf2IRGR4c8Mi/AdXjR3ufqtuTZ4WNIkCLVmzu8u9YgNDdSpaLgNbp
StIBIfqONmdIrTiMiLJzU6PQW4oaz8jvnTXncDQ3wcT1JFAZOu3Yz7HaR0g6EXPQ
DaoN72M0RHUpl2GWKdIuUc2TogwJmCeKYgk3s+gwC+JIUBHMBLfSHz+Pyw0lk8kR
Id49CRC1RlY4Nn9DftabD54qTWyvDlF5k4NUAWDuLxfkuGsTt51aK/GgeE5CdR1e
hUGSLwcaf8BEj9y6GLslnmohsydbiTPD7Oz2t97vYOyotoqQO0l8sjidOgm/P1r3
jPWFEDpQXn+zYxPf4I05bBPs6IWd0f/XMGNGABRXNyrI3SikcT/bFYnKhuXA3dJ8
34lUECkd9CL/JPPeICllpjRz5yxIsNdGPn5+zy0BZts3/NJ3bPLO56fxlNRXAAiO
FYXrixCp+p5pGfBVEyeKgkXGTyT/vrQ0k+WTtGiKzJPB4kVW3iYtVtVbQeW1GXbV
VXrwpQbPDxs79v4J4OoUy5KZWCJKVsb/oEKVbyW+Q062oHoVYLxAtR93bHuux46o
dBI++jIhZf1/5X8CHNsklLsorqW+4fQrgQqwBz2BJBBbAKwETZvKs/s6HHeAiy+u
8T4n9Ep11lfgCPo8cghZmtkvpPO9tSsyutQ5C/KQbhaeJms/PHhlgd9v+iHpwCeS
jGQPcWu7EMbq0gmUqjpEKnpFp6SNuUVxPe73KiDHSlkHrYjwvrT+bWuSh/rahtgY
kKq9G4nl0wGhiNNn0RmSynz91H35qfwspvYNqXkmVB1Nx6nMkdt5ytrBFFTttx0o
++DfJ0nz57lP4/2orGfKJcBivbhddXHxMX/22UM1FS97Qp+J4nrcozPqBCxKcTBR
5NVWlQNZ5e+bl2i8csvkvdvBjMgLxpBfGWKwLTlxNPVw2mzqL3/Igp8Zlz6ur4IM
p4kWRmegeS+iP0KJK5PRKwVUadP1SDxg3kXvvz6dTTSI3ueiMPGD3DtRNJW2NgOv
gnXzHf+Iuo+4TCUPg56nwPXUJ04QC6T4/LcOS7ePghKTfRyixKFrNHgXka2hbneT
VB564+leYyMpYte2Q9yJdfofWC71lilu+9Me5uW0+33Oa+oM8QWCmih++mav6XFs
4qEquCTbNFdQjy+Iz0O4zaQTjivRUeCo4GgmtUX+B9ApJo2LCSFw0hNJpdi9TSUL
hKBzN1KTRKAUp+pdaIFgkTBDgXZwLVvL2iD2yhPxwr+UuzA+t7uaq+jLjYTEk4FI
/zMzRXWPJkZRoamK0pWqtfreKv0UvU0UyHleQ/A8VePsgCVt0E2OolwGUNQX7olQ
EVSntNJeDNPdx/8sovaeWJgB3+ZOE+TXbUmS7XjJqIarITOvubAkefa3IThMEscm
4Q4mWaFtkFyCEifqsPV58jYcT4ObDSeSf7ncEPZQHfiPOi6O/YTRnxGeWB9aV7MY
11ypB4P+Gbcz2ikubJOhliUd2TU/WBu9XGa36WF+R+rr1bs1o1vFcdTDOUlEd386
4KTLSTotrAyvUpbjP1X8FmcAtQIMvwmX2ipUXh3BPKcbJlSvvyAXDDuzegXcwrA8
CiidriDIzFrqbP7B31ZkzsQfx5yaZAp9r0N6KTXJhHOLLFxLbR842ZhUfr8xDvBW
bUqFOnKDzPb1QRuVOqNudth50DHoH2CaC8J19NJ/tMR6LPu+JUqIxlLXVJJHTuwf
ypMQ+Chtf6uyC0OozZge6zafoX9R1o7gESOVE8LQwu8DL+JbWZib52Du2njwrbwi
zO5x8O1HMnQAqWZGVmgtJV20O+q83aVMVmweIE/keFCkkNUN3uo/6AAVUBT0Otjz
/74XxukzSIHdDv2sSLjNg+vSgwC1nZqs0xrZsuanUBBlAEUAZ4Zo5p3hWxfL8hns
0Yrm+TK0bEMrf5KilxpJO23iKa6cd6gmHskRLok/SLwep7+NtbFeda10fomclPm3
SH5d53gaZSRdZTVZpA/Mv4YdgHvyq74XAm8WRSnqjQbVj6IJ1xK5IStHaL9ZMFvT
3J739bedQeaCGA4vJtyWDTz9euUZXKwpYvO8xxfLhmhxxVKZneBSKc/J7CLrTNEi
CMR61ILr3d7Y/Z8xBwW9oVvkrR7uBYdGtSKDZ2H6zdgr2mKnT2lBn43E6ZcPSbSi
M3AhBqbVKrYvKUDUr5cxNYV7GuMVxoo1hILV2wRxumH1BenvR/ol1fpmRFY0pcVA
ieWv0Njhj0W/6C1fsSyBcSv+OdwWKSyClcGna7LSm4XvFN/MG0+4dMMDWzyqX6+X
vGHua63ekFw2sdE4tm6dcyWRJM4hrbVHZ4l61BB4S7iNVB9gz52P3/m1SO31vfLn
pRT4wt7RywHJHvOIpobf18d8Dxue5mvoQXKIChSWaCnha4Nn6iA+4PqM6v3i73st
OmQtUgl46Nyhx8XPSwWOaQoxuNlS/sH4Xi3MvMcVdDr0zRvq76rQtFfVmkaZynL0
y4P7/nbsDb2Wjm3uq/g9UIlp9pgMWgvc5xSE5YwB6O8lTUYb/ffbD4r7S3SYLLJW
rvHimyOowHAamw/sKOU5IBj/K/X/DXZByzbnpIAg2uIJwSFlh5D7S5glg6WZGWaL
UH8SyDCdflNf2LYmHz5s37awqWwzmlKJsh3KIswHnwhygIw827gD92k9+y9lkDzk
43XP65L5PcC7p2N29dx0pqySRMqp21KB0nwyPqObCzxyJmNgVr6vJ7aHfV25A1sm
q0EgTsOVEom4acuxPlOo7htigcmRiyoW1fRwoKkkMjosV5yPhLT6fkuviFL2/Sqp
kT6tD6mFeOctCGeD0IimSxlO81MyE5oL2p5+rOgMu7d/4BYnadvmwui1o8Jf/kob
fV6oXo3URl9UUdR8Q+bprG8P2jgyaDW9IsNp1oH/vlQBpINSE7OV/QgBn45ltPp8
wvJXcbV0n5o2m/wzESE+NMyFpk6QF/39b3WbiyiAhzvEbiEoYVg/qFMFPAxi9mcx
m3LV5KwpaxYNwyN4qNpH99T+H1LsXUPsXtYb+RVeZf0B1KbFq+mLKi1ArRQglVeq
okPjqTxItdI7o/u1//oUTf9HdFu2UKISnOnFCrB83vfkELdK91D5MIBDiSv64BWT
MClj60SziegqDrD1M7UkmDmy1bjaWyTxPRg+adK3Pui654p10DwZgDknu0y7I+dI
yvIKfKmzRlc+KoNmmlzjhObpRUydRpoInUhX/6yVj3PypGrCON8fJYblhNuPb8yZ
1pIuPfS85luzApPHzT4I7ZX+AE/VrPgKRRwW18kIYcEKDgCuzXLLhvkpm8epJ6AT
FYH8X16Yw/EnmAI4XkcieM5kJYissSGgOF/P3MKchUyThZ0c3uVKoRlUdwlw49Pb
H+WVA7P9THkwtKL1weKAkZOAwGvK2klalWeN7wubWp/bX7Mqdz5b8mYrnY/lFRgm
1tqrP4N1lskF7l8M3l7wahV+XmKe0wzC9dmzU4kuu516eK4gRKUNSGLONWuYQJ2M
rCtQ1YhtCrV7wklw6Du7DsvMBfydCxnqq3dT0Lm2yPYBrd97wk7cX3dRXQVzCPIP
MetqDMqSbM7541ufNlo/Ces/B0MGhByCreKYkAkCRZUmiCYw0vOq7H+Og03mSd1Y
yjDMrhuOlZcDee/vraNNAe86zEa98a2bqEhSZ8yNGAqsjFXvPlO7ixMTzDpdrwat
hCg2huuAqQrrlwoCJbwiWat2JqGmKOIl9h7w7wwdCg9qC+/ANjgIxoBE/IvrTli7
AwRL7Wp38A3POLePMO3ZFWkgpg6/sA2hYS8pRljwtZy2bjEMJIeS1nzKN+EaXYv9
lnynm8DSlRqc+v8OHjKmybIDfiH6o6/VWfnaUue8YVV+tp2i5FWQflJkIR60Q967
DCGBWILEiQynbPQeKOFC21acSjcsTFM+ObYv9YNPS6a06UKqzWXfHG67XIu1GiWp
vcrB7NYJyikquCTMnuyzm+CZBQhOn0h+Lz9suqzXtYalpUxA/loRnibqXJSIIFk3
Eq3lhZgHCdHH78ApR4XOxrSEA2oyLWlvVWLfN1n8F+yOv8dTiUc3Fh7LFwa0k2GH
9aYOA/CZu/zolU3lmDCDKEECsyJQrrYcmK3bkOruhUtSsEZY4Rv639AdmQPBeMjd
A2JzvPhsvPDeHD7p0tvQgzmzWhMnlO2sNjpFZxPnJmcCF400Vzclwcw4I5w3brfl
9nV3ddt03ayGOktQmd7IzBC2l/xwMrsvA0FKR0uIKoC4YeetYx1COAD5dozHdoEN
mII+rQ/bp/zBFENj4ourEKTaSJFuKPPGbXGm/kPuhjBvNWfKzXXJjn+SgzJ6izUE
D+ZKweOpxA8fHknauGzp7/JQGo7Gwodkp6+WRxfM7p8ipFgawyi/Mlw0WEIVAzN6
hoWHJX7gzwf0B709ONZGnjuRh6si1KlfCTJQAZGDn9iCdS5+WR0QE9b8FbOD3Dim
nSHm3zgFCNPFhxjXJfL5X0RM/HvixHz4o6JgzoCS6gcMQhcg/dUDTnxiAov8HWAj
0XlG6lMo4tlY60Q6hTDZZpm93v59kCngtNoDHkbNW1ERxkOrwjK3HgqQUiRWh3UU
I608853FTDh+1VrnOWPpdB/wK/gqelzSzAcqZQH5k+J242jmfGez7RC0ZFRUjyW4
T2/WpT+JwALaMVvpqXFayVuTg5FPrRZv6aGT8Ehf9hT5ADRUfwwVD6s3fpcTnBsh
XL5xO4p+IcC2d3Xu7VaxjYW1hEm0kM2HAuDXtU5uxvyQh7otBBRjMwSV0dJms8c9
wLOtkxdrnwaU9uFuYgoI17b48oDmc4DkElAECkWA/l4J8A0H6e+R0edt30T44abw
5ye/0qZb3gxXNHvY21F5PeSJmv7PXn0C0fgdLyzpnaOJUkwnsk90TG3XOO98DuV/
VHI5rI/aDBUSV5pKsVqFiGPbx0DGZ4UtCdBqkzkv/RsKdmWnmzpBatRTe9L/PIX5
I+mxmDMcKS9UmRBCTXrHsTK73+NZ6o2PvSCIVjyWg1CfI9gOsnyLr/fJYDX8CkpQ
kHGqyGpLYNuyrmYuR9F3X6jNCNeFBJQ/xTYNI5XBtjsrcLvBcycOmL1rvrZ7CLMp
M+bZM4myedUzX9RdS0PpQ0ixLPWSykHCujl2A50vsdcVy/I8lL3ffcLl6Zgs9SNj
8/a16A+wPKNr3FZDbDRHsPufgpPgIDCzFjxNGr621ohhmLlEhStTMBrTi/MqulMn
5v9PSXVdOnQDQPX6KJPzk6VJz08lKyHlejCeDqepkKRCVUm3C2jWxa9EZRciFPmz
Dkmj8U6e9IquQNBYeGmTiQFJbx6TYfzg62BWdosjiQfmXCN4wftG3Yb2D327diM2
C7y6wH4Etl5kq0rNJrXh6kHea360w1mgb24VZGzIHHhOEy0nUTx3Gqk3wDDOwXUq
G23bOr7yMXiXqEpCSIk3hLIRjFqS3aiIg47CboUmPhWDMdkw6vjy4apYS9YQtItL
txCkpYNoDD+WhJJzNYdfvzRJYPF2n8CCOcPpux/sLqt9IO8We0FeQ92TZsk4DWEZ
VbRUM1OsNciTmGf5/UDgs/9UMxOZtXJiWl0df6M4lFH5kLwdyTIMN16FWK0M7TNW
vJy/vsNJm2sN9zhcTOR+0T+iIoWBnEf4LNP95tBYjZfAYHHOu+lOWs5rJsVZOaSX
Of53y+IErfdVDuqNEc2p1Mbh/0j29pM4/3tEyLr2m56GplBFUM9bAHXuVXqH+Kld
qrfJ6jWufz1O3NgmDQE09n/izYc4BgSSX+1CS/fVYMUBJHLjJikHUknAt9aPMYPS
PAaLNPuKR2PQE/SlS88wCxxO6K8B+dq7YL88WTBK7b950OBvaIND1s37sMVQKsKQ
ZCVwW+8zULhhNmFoOA+cKk+J2Z+j9+vNDa6lUZtIYnGnokkp+aswM8L3nA/Hdjkl
MNv0eQSxTYBg2+dHe6tBujB2yGQs0mhubgL3T0yJc2DH+5CwJCZtpbyqeaQvFjIE
GpXuo8rQjGSWBm5gLQ3x77KPudB7PsqTs7zuZetVQcdVAoJRGMMKu5/3hJjJCiDG
WqpR81ULud0UjRMjw4DGS3t8Cuzd/wdT38yXRewmh4x1W2Z72TCBfQ8z5jSZxQ3Z
gi/UJBM7s3mdYSXVY5+sTJTe6+kFblfyLnJv7TFHbAJLQxXrrYZUlt001Q6CIP1w
ISNPKPZv32zXCZCnyvZ5BbEnS4xQ7ikBUQ+CUK3eo3NSkc6OKI+I2sK0iEyyO7Yn
Jpm/N9/B1dXs4/0PN+9xsXbwz5QhkY54iN5rP+wmgGERpvYtyex6Sn/WgoXRbUrh
VLKnh2iIQuO+7tytHLC17cZJbyCNDPqQjodCSbCzQ8yq6i+uXke8CYG7oCrAZyxK
lsbL/S4XOWgZ267N/l6gore9LRGdaF/Pl/U4cf3MqxZHhbUbcwS7KBdUjr9Eatnr
NB4WH34yaGWWr7YTuIbyDtJzOt5Wj025HRJABIQSOcQJx8TrolXlemRRv8xIAnnp
PcbYZzwfQ6Ufsr4qmsmZRNGXOMM+YRBkVVptszm7IDE6UiXLrlMgPWBAQ3Pb7POd
WzuYSKX3k6c3EtGxJ1ldGW9iWG/LtzaxaSin4ilPWOq+z/hrp4CUkNnInRCJRdiE
fId0PvBrg9XzVeZkIkAy/CH5aDKke/U6Z6u1wSF8hrakEPRsLeXyLuhZpo6IJj6p
WDBfbBrr53QeQAhAZvp3g20wpqWxLYHJTsXpUh5JfqPH/mXoFQT/HhiHwr1zOrmG
kTEZ7CQnVigyZrpUf3Szb2Hobc3kaazVV/6uTn7kNaOgx2wgRjf+CEDmEY3lxZZ4
n4nQaDLY6e5vrcpXFxtX8BghBnxNzVKAgQ7xE5Egr5THL3pqI1mIzg0dcN1PBl9t
mG3GPRHa/pZS7zJAHNYBnQFGE9Y7C+8Ic9M+nQlbLWCE1GpZJKQSVCaaGHmDYncD
OQyPoBSQ0rkFTTrdrKbboCNSnFGBkx60yG0mWgf8ytcem1tkUAkxAkg+3Dd7NLgM
oHve6T0REEp8F8XzXEjeml8XvXFvwyT17b2frtIHjM2CbIL5GjzOZWRCikkm0sdW
FzpSpvMBxj9oKvJPSrClXvKRZrEGA5d7H7E7T+0VMevi5JhzFW/j7czDi1mHJD35
kY8gEMVuwxmvNF6rmToy3L7WKSWVHvSZ2ZxRUK48F/R0SdRJHfy6ZFToNOjNKZwA
Z6RD6BH03MXbmXBjeRACn8Fdpoz97NV+3pGtMReSoMM3hflyAx0nZKTMKQicIszJ
NQm1Yf5sjmekeHBJ1HQxhdkPLgQy/NovR0QP55+3ySAG69XV2cyK2yBa94aqQXCD
IOisqKeSZCJkJN7/vNZgRucA6juHcGeuWb27F3p9JBqfIJuBfwZqIReqTJ918Jo2
iKClsoshO1RqzLyldlbh442V/ZVoaUZhTLQvUdewrfh2JvbltyAh7IVoyRYehg0t
zNVndKRQrZUXVO3eJ2EjwAhBauzrlhBXeXCcF2/M/rUanJADRhq4CEeRGJTISPNE
KUa/fZ1M8CWbMnDXMCqOR/MWquNq/ejWCMUkDAHSY9a+Ia1vSLHLRo3xdsXAm3tH
3w+qPERU+zJ3QaZolVzuJcrAibBLBJRS8ym1Upk5atiBmHXCTj5NG861Iv9d0NRM
PgfDsQ5XD/SPypq44fc+vqNgDvy/QcpsSXaOFRuNT4di3awoRcadXDbQxSYfiydm
NkCuJ5plgG2OfcZeLkLd9SjKvS9ZdEjbTZynPJ8LYOmn/i13Fo5hcg3cukdvNlam
WdTbcQ4rB5HUzxmALfsO1T6qkReQZNMdYLBk+ibhYEI+z/w/OWfpLKoc2l1gI6Nb
/hfcQ+q294LKfE8lVHIkZ42AFuXTnsVcKI+5OOZprwACrGehVpchNw+yeUCFetNp
a6zXfVyc75AJaEG2hKRJFQS3Iif1T4zdM8SaHxujdb8gc5YRCnT7E9Bzsfyu9Hu5
/yRBOrmKiG3V3Cra91miW/1zBSYGd/D1veXQuTAYbHxA+4IIeI5hjDhZ8eOXrgzu
evJLnACR9jf21I5dnR98e3iCoYC2ie6VQ8Lv65x06h8Jj2iQNNIBOmCDQH5t8eZq
M0Zij1xCnbWlkyt4jNq53DxfK5GuT5vD6+PjVTcMip2/IlqnBpXGog134pfBhzzE
9WbxdAHAIA1Mte39QWF2CDATBBzn8/c1rb3vRL7/k9r2708MBN81Ujr/PWCB47qF
iYmcydN06AGmlp+kBo9u9PgV+XfEXL+o5pq5GkxiblR5hIKemiru1G4yW4Rb+Woj
Wo8bOWifhEy99OD48Sfqiph+BJOUEt2hynrmIwUpM1slAsFRirdCEfQH34NVc5k6
vThBctFbetmnZxFvEzyvy/pkEBdw4PKVvwGDZipa4OJo4BFMk6EQbmVQlVHzIAQL
ZIEItvSVYWA7OU+WuRGFcg7B8Nt/6jAk9W5ZAdMHLfkWLVXLxT3OYPdt9cpe0AnU
w6g16+VsZInygE3uht/OGzTZ9qlnQWZy60J3Q4ji9GpvWGzNV5dWdNXq2CFw8AIA
OGV/0pKRXzTxid3fokySpaGp8CezWiheK8DqGaTG018wZIhkEzjrMmOlgAbi356u
kgjHjRVN2WNwAecp92F0PMSfYKlHsfKM7pIFleKatNn1d+b9guwptXH/xvteI3l5
Ucd0awidgfu8XWCOgMn+Rlb0yq91NoT+nRNz9jM32oTCMKecsVK8Xn2Nl2otxtYZ
4z3Z4PqCvwBwcDQlGeYCJEGyvQPxY2pjUP+L4WNQUCY6ZRYEwyGR8F8mAib2jKH3
HzjXEIUAm37TLXWHiR9ced8qgkbLWeRTwkOA0GS1aRDJBFwVMSPsZFFbGA20SMjW
rEd6R5nq/UuotrG2WFFxGHPjS/d3USnDv3JqZ5R878Wn9AKl0LQx+hZt8F4iYGri
EMrpzPXkuluOgyZ7yOMQutzbMxMShGl5jzCN0Uoh/AGlOIIdBlQKbiH1D+zbbsPz
IacZuvKO0J8/1W0/zxAQjDErMmg+kQ7fWl3qey/ymB8upAPcxUZqT+Ove3GQcp/t
KMZDAmJpdRYKwelPHI6ECrglrNXCPRLkkxIk7E++053C4GgiO6D0ve3CV8zzs071
CNuHGUBDy7LjOdKplDnUSoyDqm92kaMdYzNoKVOoT56XF599J1aQ9az2SSTVigxt
73x2OXM7xjSNSwOW0++BaFdyc51SOsk1zHysB1d7Ilmd0219m22evZpvJt/kL0pU
jmeoiXWE3XijqOX58G9BNJHUlz59vp0J/M6WzDSQVehWrhcb2a0LYPvefrraOOgQ
5U9v1XFOsRav7uQU5St9lqhp91qn1Op8d/aSpxPbQjLMlTyUVK5OwvIT9zzOOz9S
YOunUTDpH+WO4WF5/WbADVNYz2SoGaxl0Wc3sG9HtQKTIDQASTJ8w5owM7TpldRm
8D9rnd810fAIKVPkjrRBs0obnNuqFz3Hr6DZu5B2qaftyjonD1XjPKkLo2EOcCL/
/jzpDcM7PhBHx5n87GnYE8LjJtFHFnieqXtwJxoKwBmgmVU+gHdsT4wzZDprQ+wn
uHhxu2bhxR1+SgW0gTs3YFC12Jkd9YgTrH/h+HVpnVMM63sQUtX4taXMm3hqF7Y6
zbzUUA7kJvgTOlfMTW/9zVu0qzKPtgzNIXkE+EFl4Ex1/ag6DP0bwuMasXw2RW1v
TTZVkODV5hEuPz/OjMc0eUrsG3oUMtQ5rwwqwn9PCtUgXb2iTZsEIHOuUC5yFrIp
tcwgjrasyjSkOmUcA/LGre4RJAWI42FtrJ1X7gPTuF4SG61J4Qzn+bt8gf4GfvbB
I560m5AH+0jmY8yZXBpXIpZCqVYFe8FjFKl0TSFjocz/OlOkbPrKdanrSMKE2L0O
79Rub0fiR1uweG2RrCDG7ME0Wg+s/g1xEA7UL+wvOril2/j8RPvn8Y4el/uaeMXL
4gOfYv+uIMHPpYbK+g1FpMcPplQrZfCpiICRwqnKkOYxXRsparengB9Z3bBgzurO
Wdu2F/hI99NnxTgGhJq+emLG4rBiZAimnbVFY2xjnpldSrthA+Njye/O9tdPy40O
0dTIVoF4JSs9hfD71v1lXeS10X84vvJafb1yVzc2OS/MoVOXOYW0DVsUvg6LQ9j2
apMDxFzLTgWk6zV6tMroo+150GeUOL1YXSoYqKKwS+lMPpFuZjhUcu60o+2LBovx
SCItzJ/2D/GrdjfZWZZZM18dGz/1DpV7WUmmJcwxu3jLzMQlHb37kx+z9bSSaRPu
xSdMF2VDv4vfccvtzQHDOCTIEuVRhTM1zMqDyD9nBQ4wMWnexcHX3gakRy97lGyz
953iUMticIgNwoFbAq/CB4TbyBgy/sY6U1T03z7rbVeWx6vMHzLYIL1T2ukYGA5F
Fhx8tH6pjtp+Cx6eNLlomVF3dp01HVEBeDbINrzyc/ouBxzE8XICW/4dTGzFEqv5
1HdimKFe9mcJaJwQWGWb+DduMoR1kL3T3ejSHGGTLygOMNfU6APMl0QtS9kU0YyA
yzgWaxaFKR3bk35wVJOGFNUyk3EhV44ou4fowHJjVVoEaTxdWoQo9iW5s8g0kYRU
H/rH39eu2fWjw52be4K33GmSYOi03+BONn44YOcjoCvaQEJzplptuzBi6+IUIFXt
/KzTmMdkySviQBoFU90Bld49Ha1cKAo829W6JEjBGkP/PzHwRWsg7Tr7wJY8toul
bn2Jj6SMp/pmCJQSNwuI73s/JWPq5etX7tUx3rxc320Y6c1y+PbgJ9aldLcb1syn
ofmMbM6WBp/f+Qv5H/XR3qbb+5zY3HFzqvQt8vjzQUWuXWjmyTrB8gtZr8WGSPaG
Kein3MnUFiAhZTagcKBhef9wKuqOOoA9Qqdcr9aVwZWQgjdKOj5ZkVhgfGWeFS4l
Qcpgwb0r7dnus6jA5opX25rk48BoM1Jyzu1+HRc1pqOedeMfJ0ud5xXGIgOXqcyP
1hHFAxBbweaPrtCgugYbXwzlhQY9SIRBt61crmVLkEnNcdw2M/TcT8Jc731mCHQ7
boS/YV4SAGc0HOT0E+FK/3BvLBKJFbNckjRvOFNhHSQPEKG9MffF+cdYAwv+w5cE
1zw9bDMLntrxyGs3F7AFzeP6vidHnEUd48fbpdwvvRYq2k8uuwKl6c7r/qIj7k1c
2kmVeKrmW6tblqlrS+OQHEBTzBZkUJnyLSeYakMUVO/PvGTsJ8PNsV502Z+Jcj/d
acw5xiczttujq4bvCfGgTv0unX4I5MsSxzuhyrZO2YE+qbJHzpWf16NMM/JI53nz
b2ZKczl8ofjn5GD1Xl8ZsospDsvZUgSmu+lloNV7qrVZdFz9G8XdT4jNfIQZXjmO
S1vV2ihR02+RD5g2HXnE9OQ6xm38ml3eit/LlIV2Q8ra3kFmMIC5o0XFcc2KRc37
4tAa90FrX4xmnouYT1A+3NUk7ywNZflhkeAZh6bbpoVt5JUG+YftqZhilwnTQmdk
YkZ6BYZiD3LjitC9UZRqlPnh083nJ1t5GB0rvJtRDfL7pM6IL9jKJw+y9KQo75c3
kcAVLHEGIyOY9uTQr3j00ueqQTar8UqhFARjwpGrrb08gs/o2R0FQd0EVcxK+tAG
Wgu/W4agJo2Bb8Hl80luWD4CPLg1ODaSh4u7AbA6GBL6KVL+RWFX2CtYe+L+FbwJ
POQZ5SrvWygwKcfKRRNaSEWs+gIZl6wCD+XGQPU1ff8vvgc9YS6zPvQWFxbOs1FO
H/Sma2I7TgJi/6wDGoMCEaX+XozMC1s8EXeD9hVdBLn3A4baKxhyCjeo94AnVw7R
nO0aEguQ6bxiIGDasH985YTKoc+5agcaLLMMvXnFUVl6A0GObtr/VYkTpwJA/jR/
kT5yumYmMapEunBsQDt5ZwwiVZj4d0qq6csTOUjQIpL8Ohm46ux/LKrZHKpmFKsO
w88V1mTjuBVvyi6GOffR1dwOOV3B39R/C9tTeJwCJW8TSWbAY6PViXnoKV7cBaKO
wDz2EoDbjv0uzFFiF2wzK6FDwrsVfKEh1pZ6iS63z2wGyBi+e7jYt5oi207Tj6PK
So0lBDze+RCHJf60Z5skKc8tffDBguMDcrUNyeAEWuHGC+L4FLzdFT2glUMnBdpV
85a+bePYWEgMQV/GWyXmMwnawGgdbpyHt62GPOIEGc74BmBjY3W7xsU1j3XnYJme
Nmo2ep1cAVRN7/qKKnnXOuckl2NsFvhHkFl8yRLLiGD9/mt1pFwiF1dOl7jx4HTM
X2Or0AEWREPoQgruxAWEqLdMi9g5xlsp1HagMASkiJQYJhqlPfyAn8aNEVjbCrNF
yIeaCFlB0QjRzl+O2NdK6K9VNC7vkDTHGtChlh2ZWEiqhDiWCrV+uN1mIzh7tuuR
rg5e+uRjDL+wNJUQW07WlBJskNxiK1XRVkdtbgCnUxcJuVFxKZlx4x0iUtnSNst0
dLY2C2TN/G69HSjgXWvso9FzmkvVCZMzk1qCPDAilfvfhQfxo0qDR/8QmWo+NVsi
KrsucZnbxaNRjQHlvrLpWMYCU8P8bKpGTSb+QgJJuI+4SAGRPzJBGgCy87p+jsEh
zXaxA2dZaPDfsYEycntlqCmmVAoWS70FwtVPIAJQGxmK1Gg3fV8OKQCLFPS/cxoU
B3RwBIfFh/jnWOBstDYrYxCsLgzjORxmX84PhYWoafKv1TcxHpc76u03mlKhrbtL
2KCadk4qJjdSbww7mqo5TuTiLrkR1TPcpPOUakOlHTTdK7dFZIRjacDdy4hCyfOL
+V0EZMBw2ptUl59gwFwXG+ZJY4MenFQtpK2BOmxVBCiCZ4dGFWDDF2E/qGc02scN
a4A66sMHahvKV8iqOxQWI01w0IKpBOM78Akm183s16880+5cYPZQDNtn1mYTAvyU
Y63FV86eq2ueMvNGCnr+ctveE/anRNjF8lLd3ernnMT3Ai/e0Cwg8pKaEHuaPeeJ
2C8ior0feQeYebqcE6B+b/mKYhU9Lfy7hRV3QsW57PCOm9BEtZGypyH61bmopzuL
lDr7SFMM1ptOZiAtz3zFIGVIv9uc4UhUdZKfLi7VwBdaEVVSIvczgG4CizN9EUKk
1WvW917jAh15u36COG6bEFz70b0tVPTASqNE9zYIgi0N3eFUBVGXw1CDK6K39ke5
yl2peD83B6SlkY1seUalRbxYkmS5XsFWNf5UUL5HFr6F6YJEfds25AjL+g3ZQke2
0LugrjliH5et8tRV/twP5Xa3xEXCsu9Q20ojTg8vy/8zqLWbKkyCsjpEcGjqvsC2
o62eYZKuwayBcBD6ObLUmI4mBsGaFcqAg0l4cBnnnCr+8+zsW1k6CmIFtkVXW4oS
0k2Zr2ARHEEM1JMWT4VwCu+auaGhv1ze6+0cuDo/mZWKkcqqFLoyejd7viQ+f+b8
HcZXeskEHn1mHVWWDqKvJdWqTWrd6v8jWr5D92q8F19Ojo+Ozz5w+k2sDd1M+9FE
yUAj3EMRjd4yfnmCk7roD+GBphAzjjVWz680juXjDnIM0LatoGVqbD7KLbnfh3cI
swx2O2/GbU7iTye3n20UqLh0vgxS6VNXGvDqlMWyI5cc4NSOI5O9Q9LzIY1+TQRC
z8uLJ+RHRYHCyLQ10QzDm463C7Ci728qZ+xlS3Lf4qEaqJFJoticKV8S3gwzH2p7
epX7WpzrQulVqKUADps3HwYg5/5um8r4HDa1I6dUwgzzEHCgtGe2Bmt1k7bW3aXg
/kPIkTZ1A9DEzc1Oagv0EqaI277Bp/BNCApxldIUEICan74q06X9xcGOgnPF1NM5
yU/7OwhDPiNwVx4mxkLdH6LPEAiCzn+VbZDymbmd0yQwRrZPgfAJLHHb3oJx3eHG
jDsv82tvh3Da1zLTlsMAvTV7rUVuTv1+h3vN32zVf8wdonLMsbuE92u8vWlWuUbA
ojxGa2Cth1Q9skynS9j4DfIQvmIWPwtCgsaFH9rj9uYNFLcBUapqONaApSsSglsO
aJw2tPL8VPAA8REbrDZ6wrB+VpLKvxz/F4Y33xqmbVvNjDVTRDy4QYlC2s9YCCb7
nkPG7fKuBIIZo2fV7roRcrq4+fvZi/MbNqLFR1pCjxvbIMgL6mig2rFxjfCZjG8J
QboitVSNW1jSx264pA5QXj4/1wQtNbK6uEzACfBd0bMWuVdtvUEu9GhpZ9ZxNjHj
24N3qS2c+ET0A2wr60SUAvrb4JWAnsh1beyvPHi0Fm6KIA1RcIK1j1m8Z6jwXMZ6
MGJyysV+/25+llLlUNjP4uvbH+6Tafwml1OTOYad14EgIOoVym2d652a0WUW9BJr
7kUi70DyqE3H+uYZeepvsaa8Ns/ZYJ6Wi4hSviHuxKAvTaDZQUgCyoy14ftpCXNg
21o9gNgKzYzg/LC47ybg9gefQM8nfejAnQNllthPzqqMCTGzWCq+QDf9W2OwQ8eW
8OTVBEl+pZFHs9MYM6h7fUnazxNlIvGCMaaxaBrv5r9e3KZw3df/cgIRUtIf2tCg
rMWKZlHJqrkDPW1l9lnVXAMJSp5pTdgubtGvEaJcxRxYND0wuZYJG6epqcXqqfeL
3AYulJTCynrfoccEMgdzi/LBwNtxd6I/4s/3TBU2Y4nxOt6gtT6UTuw2lVWGqZ8w
xAOiK/O3h/RjnVXgRrilx/w8b0nJMO7xUxEYki2jR6ybGRjWa5j/TSEDlLvZB/VE
uBJx33m0zRmCJDUpPTzE/v3jFXvQ/izzrMrGFeSMlyyTAu+jmVBmXTn4pNevdf7E
tWIaCiQQiGsV/NQE9DmoN1oMG+W6GawJ+EaTo3jSTVLMGU8NLAcKF50EWDopjWiU
DBP4VM9TGAOKYjtutOam/XViCb5x9Mj+Ad+0JpCgeNT1WQ/KCzQyuzNDOQqEXjM7
u1jKdnn4ueCaLXlR0Hax/OUSRvDZFcR3U1D+1YLkAkggem3Rk6QCRhsvpLT6LBEr
O8ypd5hi5MHLH0UhqUpai6mpL4LU2Eh929NvrQ++RZcwGhyIpP3qM7Q3PqeXJsbt
iUDkG1/cIla/gle1vrRhoJnOyKaG8Q/rdumwBV8rWvN73Lpp84AyRgVBBv1X8Py7
piE8aDZHhISJIu9QGu+bSKS7yjxitHK5/IfsHD76p6btOW3PFKOLJbHNyo+v8ahh
1aZtWKDosnYsNNFxhjr18V08NWSn30yzrt+vGoqbXktTwHZy9TMq/4OXPF0bWeIl
WZxxm4mLTm2U+fX2y3NKdXKcmMeAthzZ6obUFdqzrFKv/1fYDe4dFuJFtfjF3biW
F/s6b0zPA7bQuQKxHEuIqm8u2DfWIwPOqyJfW+d8949D5hCDXhbTe5Dx3LTr2pP/
3Oa6F/EsYg3zAWlAn2CcCaW0pgw5LtuPOj9vPtntOne0W7cT7w7q+dT4/xqKiT+0
5eWDqtR4j9k3fzxq2MvtEKte/G0w18MtTwfa9GV/Llu+o//m5ldi1aH5p0j1CTBk
vu4MVVmEBQJ5XgmBDrKlHY9UDO0sR3Qgcowo9IadNtRY7R/glW4FsJF+4MJUO4mS
gxUI7l402shc69nIkn92o8pMOwG/V1hrum3pQXNikb8lZ2LPv4BCn05Mk6vDqf8y
VvIq/Eqk0eskDsFBOMzBxkWqDICiBptndmfa8Xu6RGvtXOXXCP+jYDLqTRCYawT8
fu8cUjhJhp8SDXtYGI7jkDFWmG54L9mGALk9xC/HB/Cw88TeLapZycUYQQ3tXahf
fNujvRD0bJBRxpZZjENVZDc0g5+ddpsrPN6AP6ylrtkJrT9s5Gcqw7rY16U2hyuS
g6WKXqTga/gf1248K3q3Vu8MdV+eWN0wAIRoWyn64iCsL1sTDAl1vsSGiUYKOfpb
gHs572b3BUgoXgOXLQAtxx2uCQ2hlMJt08pt1Gip2o2mSPMXj8sb0ptUOaZ5wgd9
hPc5iJOTCg328d7ElgtesZKiFP0ej2W4Ym3CIuKcyywTnvIfI4fI1AdNoy2JuaIh
U1JuJsIJSxjehTHh2br+w985g4JcN3nD+/rIh4OVt8o4mK9G7OVZx1kXtnbkNGvu
AXnH6iaBLW1yMweyFe0b1g417ZV2R+/ymjOCMfjl6d9IbUpfxJRUmsakLzYYgfII
Xj9Vy3cik9v9Gx0D33DzqornO7jZBIMv2+yOKevN8hvSritswisRUxNDCEUySAwt
ExUWzSyDY5HKNVgA0Drw+4TJbukNNYfX0O/rN3fOOeZSG/dTL2ossK22H7ray96p
fhImJhV2nH6ymMSwv2Wvm0Z2HUP/oS1TgVMxAQlg/t1WR2KiSYiDSV0csGz9CHbK
xxVCk/p+5m1Z220ekPvWiHlK1u+sZKpIfH+28l6k+hUWV8L8/ZBAsEhJVJ3fsp5l
4a+61kWLwLj1jN/3TgegEqeI/x2R4RI2CkbUEbQo16eK+1rdOqk2e0tb1g/gf5uA
2QGZ7vI87T76oPoCePnTYuKuRlIEJUKnX6vJ4FLs1zgbWW2eUd1X9c6JZ2MurSh6
0ePqPwjtXu4GMef7L2U0jAZ4fj8Iw4eSiEFTpU8dGdMJu9HWoS00LBVSA/MewSFY
lt1AFj5DJYKJgJfELDFEg4ii2yFLGgi7L7k/6o3MziVQJOSmCakwi6wE0Rkmt0y1
KkAaXh1VZyBaABmAwN1uuvMpswa2ZsH81v7pu8jJbDOCNtoe2zTgNK0rlJqgAmvD
PKPINmn88Wt2WU1UP4qYxKkwwZrzWHZYDk9Zl7U1IFs7Z4UrRf+P4GN4TGDVg5oE
Bd5a0nQvvaxy5t+LZEWXVg3dUfn4MG0QyMt0IGeLqtJBWSrkZZc3DXxBE2tTlis1
GhWaSBW/02vGO3OqNJPKCzIw1aZB8+TooLhlXcXcopABANjaTimbZf9W4r1d5vvD
T67J2UKYdVYrKy2RGIK/ykZqQhCBh+nQ2TZ4cPreAlpjGUdDfhQIDO4A7BsvWoUS
o0tIbEprGNabnHs7JVMsM1bXQcCGJCuiKyfDanP4YL67Q3pAuhlifryeBYkozBDw
rIQ2KcqAeEzduK7/wWwhN0KbogfSDsRbTp5C5RbikIN2SKx9V3LMR2w+16wpccnl
k7lShJeGiK4uPWAg/Fq+iaqitUtGLc3yU+NuP9DHTXSah9L7My3AyCH37dDKbSLB
dH5k2YgG9B/Qb9uGlNv/dA1PQeS8+QNKV4hpCyjbhCRvjMOKtLWIUpx37PrzK9Z6
vBIo4+b5HsyO9dwx0MhAYKZQrhfyCb7vBjVAIKtDEOf+XiG7i6JdMu8fDIA5fDWa
Mq0S+MHmhCh76QtnYpvFR8chO0RF5qYnIiX2mrmV7IrDRuto6AVfMU0r09s399PP
K000rcihKfeIedKo8ufS4YZ9x1ffeAsZ1lM8niK6B6Od24oJG1S3HlWOOIGA940U
rXvXNPlbt8r+u8ht/8UnawkW5m/LKm7P9GoynDKkbwJK4v+VMfIxsmO2UmVZXvPA
xCZmPU+gaHlzR3sWkxgYptOvXyTc9MjPX2IMJZEC66mqcK66SZwnwNqs9stJkhIm
HAOSdzAiUG7Y/F3VB2KZuh9DdbtS7Ame25/TX1bNfNG2WysHSQfIMNkfc6jjYGVh
xBpJB3+Qzfrce7jmjgHfl64Gn6+uip3nesNF+KNsmcP4O35Ryq8S4/OHHT3lxyz9
kxdqYxf1CzSHc8hTB8x8rEn76rflfuESvc25/ur4j9Ox+5rGy6p9Vp0BFhGAmv21
ifDuo84xKS2JNSVkp+Z4yOL19JGfx/Zdu+s1Tq1iSsLREsYfhOKKsJCsuRU5sgNo
anUWo8gh42Jn3X0hKQN7/V0gmeXl+Y/iEQRM4mSIF4u8Ot7Ns/Rz1HlGLh31Pg1+
trRwXhxYVFlTpX+fNcOVduakNdcLddUXSg586dKGOR8vnD11RDqfBgVEHkJXX8iy
qMZMZxhPPzGOoWqb//d0ENRiCVKk2stE+iQAfV3hgz65UiBioOmXffb4gOglmf8a
pOU3UkkNoAHVNobAquN2qtjC8Z8rh/rCKdsKFimO2L2aUB/WsyP3QlQCZI0jJBxj
YdD63Er6rqM3da8R20tiTJcscu03UEpjrgEy+2T4/S3Ek2iL4Jw5qUjWbo7bnod9
ojqZO537j+mYhTt8vX6h2NR/lZq2nskqQKNvp6pQO8qeN5WCiCHwlBMBNqmnRyZr
Bx2fh0QZJUzEhSIXIvuvTjPyvxjfhVS2qNyx72CQokEQ9zDj3sb86I8OWD/5haxp
fQJVWBZx+mw8pz05NCW12iT2PJcOSTZUKdfVfI1Jl9at7V2GvAHjNvQgrap/bH7b
qz457ZOXFXm96RFQcLEP2WNstLyUl8aKKi+WTiXTOH01myl11FLlrtUWqJU6i7gz
ntMBmq3ldlqlsaz6OcfKuryCXs4BsNw+nXTci0Z2d7ctOnMFYvMA66o2mjDM05pY
12k0mUVpfo3OGeWl1YbfSquEaSAHT/yp9akOCAoKMDmZzwoOZjV5uQd9z9gV0yEq
GT543fnmV9os1mO9dI58x1tPBr1MLry/3sMqhNPqFVGWBiD+4cXBCg7EB6oR1efW
TbOO1yxLxnpAkRFIedvuCXnStnnv0KCiFM5Q7lbKvg0dctP8yB36pucg8kIYyVSk
FCeaXg4knX2OWDnKFRk4E2JpUAbdZcXy2WUG2+iQf/TClESTdjnzLXz/euBOUvQW
QVF+F5EG8ZSV6QvZ0CYkv8+y3FXlJ3IIiizpvQ3E8EoXSZWNHIepooS4JJeCwLsE
cYDsr7Fxd6E2AcAw4SBCBYFUPd3pNSxzsn7AzFMeXvwbuXKVpkPEi4mpFwTVXAez
HNDZ6Ygy/e8bj0wb9w+AyIKW7lMlGwBE/kL/1TviQd0X61uloQRNvIVxG3iRhJXr
RymU6d3NVCL4DIcCq0hY+sY9tPuRQ0XISKI0gIyVriFFcAwdaXH9xW6JSEvVAlWO
1p84vKbrlKwf2+zJuGelw6nTfXV/yvooULj8r3Z2zZvnCGkliqyfglEql7dNmKME
WIqF38XO3uJk7Wp9H9JiQssU/S56pQe/U0KAEt0V3fpOG24tppfqdkKSDS1ATtDL
Or+bGuVmOI3y1CUH9wghc7lAfV6kQdeEgqVzAFe5i77eqvkDgHOo/FLFD02kcRGV
iXcX26r7vejef64uBsotWVW41iGvPKve8zwFF/aBDF6fvhCYdrq7KksQgWjA+s3+
UjvHcVMPVN1sTavRSMSOEcIiqivHkodoQaP7FQiSrn3aJOlqmtXcK9UVl6T5V3MS
XWzRqZFHgDKbjUV1MqUwzunW/adcy5Sy0g8Te2bvqT91fqih94ctbmYBKV8lkeVK
QXGvB3o6Gy7sx96RE7SDp6Vzhf8r8LguwPXNQhGIG1iRLwwdGkhPAQ3MxBWrZYI6
PSioGOfx17ezqqIRcQczZnbvLlpRQgxcNC4C33Z9enzF/kkP9L02GNwZh4sV05Aq
qiWGWi6tnI0NYJ4vCfg62e6kZTsckg/32XDnSwY4E4M9omjdTksKckL3dq2mJC9+
y4JKU+6oLLQU8pJu+gYxC9LSNdNp2FrZSx9ue0bqRasd6MBtHI0wyOSMoGpDsrq4
Vq57PnPH9DM0xpK5a4znMzI+Aw/45rF0NkB2VYMh95gk5eNvNBfORhZrRx/RtyvB
m6A1j2EWGaH50H3+xe/aV9UWVy38mvOzMiSiJNTYYVTTfTcIhtUyiGBePBxiAaCF
Zf4GQjAXwYHYsrJUTIxuuD/++FkOmR2xFUEBSdZR4j7U0y2thZLFtuRGgAIdvPeW
Fbe40Pf4XWVjzgPSLP5TPK52SgY2bnRo47JGnl1AtPPBsYN4g3LWeRQG6407Lf6T
Ss3tYsW4zg3dRAQlDXEP1+GVB3bpaMxsDMSaY4LVtCMrVVEheTJSpuu8QfG8pcog
/xlwUyK5EG//jfcZETQQSc5wgZZ96Kf1YWlMNrhJfn7o8IF6xBHzlmtFb6bPk0bV
+1eX30wcT135lRZu1f+Jy1VAW3w9rBWxEfRyIuz4rtKVyymYbJUvypRIpv+AoNxM
jjj4NcfyVi4hnN2kBGTx+rxW85Yz6a/BnhLNORPohNH7Bx3DHPW7phuahrcTE/9v
BHNbOyL2SoKF6Yx9W+fkURTV1PIzeKDh+4XoB3dEYJv5pXjfDbeC6055tjvmQmfA
aAzS9J4yo2+QgMg8mRZsP5xpXdeZBabteQpLxtJNfGr+073O/nsQHCuXrBpT7L8l
vsIOy/7JYnIl4yIqB+qlrWuWGaudSYQV6Do0JhzxwegFOKEmIzeIHlF9obx7WXxu
upgnmZY1UflouxMnJxB4E2Xsx3AgslgpZ6e6DP5ws7i0MS5Gi75tWpyXVErjazCV
nPIlfBqYtAfdbCEyWIgrqxOWRmTgB68GvHC4fCQjJ6ik8s+W1/EVcJ97J+D6Sx1L
bQp+hmNnrukshgoAMaXegS9b8QgqWpgCfoxddBbhwt5cxLZ9o6Bhz0Zs7eDYqMWC
CEo2YcwLfpM0cRCAvZGRhgcFw5q/CBon91yPAZqrrcR/CQh6bu9bPwG56TkSFdri
Pq1KLU6iw+VVnrOIzYVnvbOr+pApAEz/xJm42WvKgTsUci6aF9GUbTYxcuY4LnUC
0wm9ZXE/1ld+hCer3tJHx4WA9VzTH85drAssNZugW2apYyeRYpXQNsWz6WzUbYz/
z1dMtVMhwGambdDz3UYDbF2vv+cBKZaaxX8TG31xwSjoqsI+C5rAAMOATAKhxkBX
KsPkxrlSFrPwejZUYhDgxjPUjZbulebY4YG+sq2lScTAS+NgF/HSYQ3Mi7ZYhnwk
nobsPzgSAw5eAKj1LCSJ32KgrubrkRqeYB9qHbrEcA0lLVGEA/BhKljOwSbBm+l3
rOzZPA9M26He+fNH/JFGFVMc9LZ+KIsSd6s4LL9ORTLJqj82FNPw1qi15dQ9SDMI
cjXSMuswdFYL16rPVB/kaUer8ixcSgJzFrSXdQOIlOGVx68oMayKwVS5y8j8S4Ef
ETUoxGwXpow8rtu8gjEUR/2HHbDTdZTbp1tGPANNXjhxiAX2gRh0KAfiJ0oUeCOo
n6QnssyEOjP4kY6Jj8ci+ekRDa1MAT/pWdvAl59NIrEFkMWuOxw5uEcyOiXTMtSu
f3/U+4JJ5b57Fqbd79uo105oO4vyEZpEPiwUoNY3GAd+b0NqZjwSzsxmImELHLk7
BfV05oVVbUDl4a2PwVpTRB/35udbN1xd4oJse85JFekm1/rXE1WlwwD1ZQf4Mv3i
rFT5f6ct6XI+NlBYXUK4ve4AUpVOHaeQTgMnAw9RimkjXPgxSiyNvthpXbmbQI75
gvLBx0nOa4KfuYiVT0llXA/hO1z81gAg3P/ba8NfQtn+Ppq62i+hu5EjxfnxVAUI
JiD3CKoKwakELHk2c77RuwnKt+eDJdY9YjkCMugA61hvvhtJJeViYHju1ZKJPR6g
q+Sgo1yc0X9WP2ZvaDi5aw+tjfynEmer+4rjKjKStoTuuZmtA4ds9adlZ/NVCGG3
IUXCXxJFifWfSL4BCyxzfdmGU03VAOMMF+8WLuixgSvT1CVJ/TNiSroF68wqpuQA
5jdZmeShkt+Uqr6MAY6Uu89z6M8YVBuqX9AFMn1SkIpAnBnpWwhBXn38UTQE2I+p
liQ8j2av89yffLyeMtuiQ8v0eVzNMn25HzHAyWpRk5GJwM0ICFA0Db/evr2U0WA2
Lr4Qmiy18knL9ROWy06taU+CbJQZPISsTA9Tt48mBQL3+nEdmsyTpDzRnFMQk7E/
5a5sMwkkH/s1OKIfZqYVmS5jXUcgV68w9XhvwwM8cEUbLU6SGDhjRfilmVzv3G1o
FqiCkBNO/vrghVbvpquu1YEgOJ8VexKBGTyqkdqyyZIlCA0hTiHvxuvTVchgKGE+
1GiOwXtDtQy9YC16+R417MBmHCoQGcUFvmHK4u9wq71B/5A0IM2OxEGTSv1uEYRj
aCFjhJIxJ+YEQoePM6DnZfsByQF1pQEbzre+FYM4MagmK7kbSFQs3ox2GIPWU/qS
YrqYa7V9tqPi8RCoC0JoZxjC1lPyIqqclAbJm675Z2br5j1tAsC/gVEJfe982TZX
jOnNtYyM8YBIiyxuLxoK+hfb9c2ckjLmAE8kONCeXXyysg5ZHzuK6LfOkMUCWzja
jN1FFKRoBoZMfbhNRs1JPsOR5ucoB+mJlxivax7lEgszV1WI823v8ggsvEzs4ib9
empn2h1xwq7htDhjb9HW0WP+7jxtuOCu/EEwCrDU0te6Ic1uLJj5kVOO2rhFqiyj
laOmS2gnq9/BV09pb+MSDoO4Ryu5j8uArCEM26jzT9CdxfYXDqlAiAIgBdBN1TZC
CeEOVl6uWQBdNOdjYRyvv2zlDDPhUjFEBW7cElniJXW5VEuy5hSIvmNTe5RbrAJG
QoHuZOCZP7iAdeJeG5i95neANXSxcfbHcbvOdsFIiZ0rHt9fAQUQSds2o8+emmqx
uPqSVF56JOYJRYGfNV7KUK75dn9DNBH7iUlr7yz4djFH3jF4ShHyFsKtDaoWk8ZR
4++VK2fEeyVlxMC5VDqdxOvDhTjM/pE5l21LVkK4ebEie8GZcMXiWSkIHRoluxrx
gXCSiomV5MaG9j7xEf/rFO5btw3fLwxeGvpEjQCciudqvte6RP0H3k8GEPbeLhzH
QW0qi2CH0bu0QR6PZLIEcIee9GtCKKHIv/iT05r2dlHHL0vA5791uiETu5kouweA
Ck9hlSYsz6UCOI28ep23pMDsGf2t30TVBaYYbTgiyoS48lbapyvJwOtbaO3RPTYv
JjuVhKyxfMkc5nuR23rwAqzzPgAQHlAojIUXgJS+kiyK/ZKFghzRqwf6ZO+oiptU
DfpcXd0Llt+PlCeGDILHS2L+YTP4/Pd1dmpndOWMwiE0Kh/Q+PaDBGUtAw2rTstQ
4To9pvd+TpzVbaMRSuiPPyIA2SyxpDF64fICAdGWLSG132mK6qyJ9Qm/khRT2hdE
ED0m2dFTWYYMtv8ugCS2jLdpoNZgprjmuU5XAoSRske2CC07dckn0y4p/nZgw3Yr
wPVZkx4r2JEmKASpKZdx8A3YhLaNzmkmanO14q3rOlfns00TGn6sJKUmr6DzZ2cr
Y1faQ4hDLOWECECr7gBC5fju9y9Lr1AT256A7SBUJYeVw5CDZ676k658tZsvR+Bn
/bhTvBlJszWElfjTRSUFatjCozZsjqbEv/re20qvJLDnXMzmpL2Xxbyjdcde0jQx
MvVcFstUaQil4fI41QOeJBDRZKpZVP4qrxZ8ZPM0U+Kl7GvBLsGgIhq8pgxeeAWN
HUoA/1GIXbTustr6BFw7iP/I7ZbjIOZq3cYvQFSNGQpHagZBjRm/WxNJvunUsnF1
kUocU/o14ncMcehmtlRktDhgKLEynfUtdpiSAN723KXdW5gAB4K2RRw7v94AV9IN
1sFv4WfTcp6+ZR2nH6u0J9CmkxB+TTyMWH6N2q/Ako+0UX7VbdHCMzYjhj0OHTXW
Fc/NIFp3JGMr4zcvydhxFymNrSqJOnRx6QBL8qeQmwA9ptX4gVRxjuPN0RuUKymA
vOVk3NekfNQigmc2weaN2pzaMASvfrhIbKlixLv5lH3B+VEOr8sASqBeKVbhPMaf
dVNkd17rLY1lBVsX5SkbFZAjPu0d3YhkyQEzfh1MCWqbcm/azFvTQPdq5DonzyTS
17jOpkHBfGkW1uwgBFnbiU8cBirugKhNG/OpL5Bhh3xb8kjpvxGIflSE6fCD+cMA
+iaezv0H05dLxNM9cWOwXw+ViWls8lBfDOehuLNYQy7z04OKnX9gaOBoD21+/1b1
uoVY9aBjVDPa0MRspU2SReKKLESQ5gBY6xufncwZ8W/5syeuLQcr+9jum/YqeBnE
lkyRMOXwNs5K7F7i/2OVIfVplUXYz9wLCfiCOQqQhVv+8dHpHwMD5iuH3WyAN/nz
i8fboT54ZdCFyC/DUMQ3aMGqqile7zlgoBZGX+I4V29IOuAod24K5QPMyaredxgt
gNX72DRd4ehAT+PGaDegcGzGrhf+kEVWm3pooY32fYu5Nvppiva0vacZbEbn0aED
+juix1gSa8I4I1scsAuS/pGBzwAXL9ErV2T3r1vREYl4gvQX+w9YCCwp/JsLuEPD
5VCcFeqkdvzrfe69w1eUy8OF5UocmYTkLJMilazPEq1Ur4ZJ1lxTibmHom9KC796
30XlVEXGQueg9EEkn662qxbfRM6TyZJ4CvC7Zx1Lsz4lMvTaH/YDvh6IRIUI2a0U
rdtSzOwy022PZ3rzoN7A2ZsHHK5BQK2a4AlNE+o6btngvZI+np5J3+iZSlJa3Kyz
xlomqmWYLp/eM2x8w8mT6EPvEheLPXImLzSp/m3MSmSJDph6ck+hV5ZWPxlTrZct
aN/6X9BNxQCoc6kVoSVM9PPUmT1UdC69zHfXa/SCtm/qFRoi31ClLaXRT+6WPidg
18QfdzP/PQbgG4O8zb1GyvrNDXfOQkhh2yUjIjVG36XDjJhtzFBP6pZeIel8/EBT
46u+0nu1mZAYn5N0Dgr3UawQnB5cFUxHarTV3fi9RRAx7jpDseuj4PUs9H0U3wLe
lejLccuLv6fopilrT4Z3C+6fzIwRne/uGvbBl/+9XPPZ0NPOMR/Xgmg40ri8/Vqa
H/NAcz7F6fulQj0CW945YEmxjvuKxmS0hOjCtwDoCl3R7MPkb3HPiAESH/KVomDw
5Cq5rzjjgGzWra3Z35p+dmKRpvDO6pwFwxQgXj6b/j5nOGl+1kwq+1pLEC+ZxZKg
BdRyHyS8U6NisduMQUvIKUG1s7FONpSW5pu1TTTUTLun4Es90ma06RTSqXvzhwpu
Ih+7IdoOQrjIkF70sVhIyduwcZXO0R0aZq9J6iNCh1wQhBjjr3z2aUJkHMRaKV64
3nWb/XPZLdUN958Y/weEATEWHgbjUclKhr68z7rwpSkMQ3jza4I3RImzZ/c8KQP3
CWKrS1fu0+d9sLSR9y490feqb2pXmrU9UQRcRrNBvZEFb15dKT5KfEQkC+RF8KSo
7nx/CW/sJLo3m2uTzo6eaJxi49qtJ/k0wuobvloxhx7rW4NvzsvIA1DJhAC1DjGA
TiuBowTcTOTBpBHvRgAJuuvbqW0zGFYraIlLLrWPHt2AD9uwU4EDeqBO57gh86ln
/IZGRn1TfGh583uGkYfBUwHP1tQq2zM7G5/kVKkkTubVAGuJHJEgvj7VARY2f+rc
jlpbMYXKWTFmG7doItM9/zZKSupNqQ/K6I8KrfpSN6z0xxGZ8m0F3+skWf2RTqTk
3rcpN6i/MD+ABSR4tpgyB9D//Mj+Z1LcBTJ8QvQydnChARvH2EiHcAQmhDeA1vi4
ABCbDeNwfbRkYD1pFUOiB1kBN5fpxxDk8TUk2fY7D1Ke9okIdXvFbAYRk5jfFMLY
DZ7pWJk7jbl7d0r1NlGbZfjfkv5SodQdxrB98z08VnU+fq8K+IYZPM5yCpJjVbgO
4cgg8O94d6zqQhcu62IcfzNexSH8eNn83aW9YQJh+AX75cIqXPogPwnLrcDM0yd7
ucthU8Wn2P2HCl4yH3NyRtppQMb7SrGZRLQ+V4xroEA1QnJGJ/9VasjicFmOV+RK
xWp6I1ZntNLDgi5DYVWv/fVBcu1NQevxxfMNY/KvOPxqLtkvzQg5SYgmeZAF4eJp
OVhVTveQqFaOKmqyo1v8qKJpCSxFcQee2tJM8Xz65y0Do8HuxN1B63midD8qpYXB
Un6Md+8P7dlSWSE5KsZaENudNgOPqnPrIYLHkgYiAZvDzv5no24ZVrOOxgj9OG99
ovqQTWxcYtpz/kvkWtKFOkRIYkyKuIzh46VWrFuHUOjktrAU7r3NRfQENVlf1MF5
sxKDhseeKpgoeoRGGe1mTZ7U39EnRnsM+/24GFw/3sGITn3hlITkDhlMfwdPmSCM
fQvSdDY7RMl9Z0KQ1eADOLfGV5wUpjW9HmejwP/gdCeujknme//NHZpS8x+fEF5N
Ad0svAinWdj4b5xn/JPv4Nh1IvyBJMKqo4G1wzKjczWxDMiX1vOd4K/T/fcyeXb2
mkH1WqAUR/dsU0TmoHjk3jAz6IJwSf9E4HFEi97LmTo4k0GQfc9vtAikQ7RHkGO9
pimW3D+NPMxQTEsP3bcFGNHM6dpabvA7ZjHaILMFvgHE0K6+jBNOymuNgOsE6muH
+sc+ayvuyw8u9U5vheOhzQNyzaQFj59WQ2nkVAUe9MU2KWNw33ubGE4Fxrdv9Gna
Z5I+umVkils2lKlfJO4ayfQFC4hl9nMnIErBYglY9h/NC3+mM5wDzeqFF06QGgMv
WmBLaa1SCXi5EmxAC/oW+/5kegTzJBkSYLVu7oJxJRIeuqHShKLiDNhZSivChr8m
gB6JfldZLGRblAX0PhiXNjke6oEcE5GF5IHJE/7ZUlfBN34CecDaMxcaJWF5H9xG
0FoGb2vXGF1+A3u1zd0Lqn9x4X7QQKw9DARqOh8s/E92/aLSz1xl8XOpEV/4AR0F
UWXBZ/EBKtgWfk43mDIHaQoeGbBXzoxUN3SNNxff+qw45lMHJ+wQr8oRADOTKWy8
vLy9u0jV9mqd4actLyEmIjpDwzwqX9LMmABSut1OSzpgTIT6kvTkJUHX0mk/xws5
dYsfBiU1xsm9dwPxcjaulvG5hcTZ4wwC8k6pD8SdkeKh3NU727l7UqzRwZJ9vh2x
tbhQLw5z4dtuCDny4ZT3fBb9G2S4hZKUyyHfpU/C56RfEeEWP5t9Q3ibkNC/+o0y
KxYSmzhQ2c7x6V1Yfy/cwFdDcr6I7D/M6sKvYFOEf/EC1vkybgA7EjQxkvSoI1JZ
f33CMCjmKp0/+U3pqX6MkZGGm8sZwvALj5A7H2MgKAV5BRcBU6SqTQyjiul0JOe0
p8iDHoFwpkbBqcDa0DWWhLRIzryCAfU3zK3c08RwkagQ9Z4tCDOzyRdCEHpDQv7i
ES3mkZs9tQnmUKkpbcok6go2B8oJBwlDcz12gxaUjnC8YusU7B6P+mkjgMlS4qg4
klWzXYQrov8shHz6j7CX7Vwj15AB4zTKLulMjk7Im5mdpdsmDpo5mUF7B0l3O4/K
JDQXPxprqOOqYwA0jiEbIsoS6l610nQWKG8cMU92NedUEFMP07wJ9FRCzueE1eh0
GW6M87ntuZNIpfAZKn1zNwedw5b9frJSd4qzBek7jfeThDNMKEUvQTPyDPUia7XF
83WeU5kj/1+gTVD0Rzm7RFToAU1S/KoJ93qhUQEz7mphP9/UINJLcIv5J3OuCFNb
vpb1ztJQpZEaIjqE+k7puUPiDNtzV/8AyZqm/GG4I5gZm5L73Nz7CKLTNUlvVOZF
hyVjrzgV/fQ41UrbUkep825z1cM+zDg5WgS//sDoGyJI+2QMV7DiJ8BPQTQgo0V5
KSvofUoD5Q1DiE/M3elBrzskz7dRYA78XTyFRzvmo4MSwK9eQQTW/YJ3IB9pK5IQ
N2cnmEIeLtHnLDf7uX+ika0oTDiImSw6yEFGxjYUpsoPs2mNcK2mdJlSF/uuLySi
/qgdjHKznzH1BwWQ/WCnetcwE6mDfdoNugiEal5aGzeeTBNXqd5RelogtLy4frks
6pCnFxcuYhuyh0dEYrbrOYZhNy7SrbuRUe3qTtXfdXEn1hYIuqPizolTK0nzuD0F
gSAXZKnzajxNaedHGDmYSRrn+4JpycTWDFlvW1iSrSx6G9g7dpuWFA6aF7OeshlU
r3iNiL+cAbFHIqwldAns/Vc/ArZUOzjhcmpObLcHUPn6WFXFBRK/UuGmuWtARx9F
Jngp+Of4LdFDE7KMNwgSBD8WSxTrijy+8Tq0CEY0x2smvps7MTpK5OFlp+N7tXPI
ocYZ/KCEVXJOTZJbZBQ1xRUzoyeOnNP/xXR3PEzq5wvBdx0Pg2ORxl5XOWHYWkyl
QzJtXlH8nzrEU3Vz6cr4uHnH9ZF/k+Tzg6THuq91l825cukzCE8f1Ln4luzoEdH9
x58++te4quTczaQoAvcQQwSN3BPgp5RHFff8UsKrbt1uu2JiDj5PhVtS1LVmAYDV
CyhSHHkZDOLwszQPV+1a8wmvOKRijAs5IuL+Uz4wCNdXTwVmVwnL20cO+yLlzQwm
hQHgC1T5aGK8rxOGO3RXBQ05kEC2Ct36dqYOVFCdGyQW/2ttEDF56yEPm09FtipE
w6DW8c4PN0Kbo7HZyBZaqYIkry9AJ3ijMKEYgM9+C//NNCt0ht/joRzLaq/oBW7F
+/OGQ0633wY9Ztu/OnmL8XKi89lML9LiAijjoEN9W/bml+YEylK7BcpatigGHBLt
uMBz02WqE/u5BZWYOt23jfIkIZHH8U/n7Ku7yoYwOqRvuVx06yCU8CaJeYnBlnNW
+PJ90feiUfOSPNoJ7WSWto+/CX0INC6vUUC7OhzoY6k1aAHUyf0CmvJqbgFz8wtA
h/6dPiDnAhgKltt6O7Iqe/Op2Oa32b1gOWSLkpa/oZPfYGQfuTEUk5rdjLM5ohVp
Wz/WAaG52mOo4tY35GvLN7nQvddmjtll2nC+WHXloKJeEvuijh/q7yOUpmiuq4ux
/cy86GxVfoviNpnCSLwv4S+fqRBQaQ33Pq4JPedHDXUGSBrpha39LJE3AQh4rKTT
JIo6PKPAhL2yk93bg8eV+tbdxmU6Js6xCk3skIObv1FBRhEyFbbaush2FrC4SSmp
KTT2Lvyyqf6SjxmAsr3UVLu15YRjcpAzZal7iGrQVR6PNqWT2Qb9UGn8gTwm0UDE
9Qi0rFugD1wX6Z5k5HNfeZ3ZkD2L33kBZ8olcVSvUr6JV9RTb7p4sxDGIqk5YhmY
6JmzGHG5pwlQ5nSrH61OpYz8DV7OCpjpobxqA9EBmn9jYy/h9tfeqFyBhz9oaFkY
fOdC3pLtlcTc6JtutMoPNrTBT351hC4J0+YItNYOBoPd7617X2/LpPa2ACGn4DAo
5FRF/ClaslqCVubqqcwi9r/XaqfCRHdzcpMNwE+WNChbwTViPxBNhn8ZBsV3jVhm
sUnykvIz7YAE2inXW1JzAkMDWv86UVZYEyBd+w+qn8OOyKOq+RFkkKYia8RIIcUZ
9Uh7mECHVYlA3BTBoYINQtfDnFEIv36HxlzKAvJMoQN/8BaA6rJS+y+YSysAb8fP
2q4GKutiO+CrOUaKiOebYzxdoYW+l+xXbCXVzz5PPC+qQZw9Dbqa1sTt8b3kL4P5
DDWPSODpGwN8mun1tDakZM9SMFw/HYwi5Petx0FLFEKgpRiMj0i/A1e2TSCAp1No
kSt1V8CZCU2Ic8mkgdRdTR1Q1C/sSqJDPD8eH8APGEMfu6RwcsxeuppwlK9ZzOdX
UYdoDx6Azck/tWQrw/qJo8j0fx3drxcSldxdqG4RRGw81RvBLqRBdiFTxOlTkh/D
G1a6b/0sps2OSMn5iJV3xppV+0kVrsCl4kAC0nWwT1mgaBewdFJ37BV2fHWr3epV
4c7juMqX8m47mz6/uSE52qZXL61E9vz/8FVGRaR6vYu+m8gPWVkrl/QFnEbbfV7g
+qpJaTNgq+r11K11I/qVGgcq5mC7/UN7P6Il77dRciUGyB6Hz5QDTk219xHX4tOG
QAGTznuMBoXCjd5XRskVzG9R8A4cuiNdDMrdkHfVRTV0cillTLSgVxq0BRTnlEAJ
vIWhmWsaYwe2nEN+muda8NHoDlyg2lYtfQVXHfxOiXOwAJu07l7B9Wf5mc+GgOkD
LyvE6vIH55IM2syqiwbnRn7No7f34pg/Ke9eoilY1QpKNgm+JCYWyPVQXhD5vBv1
3YTeiEgPxAPDRDjdPQK3NzZw3c5D8qjsrSwtM4mFriuDmubk9hNy5VWfGMIpa8k4
zZ+aboiBsUm4QQ8lng/BePNbBzoG1wb1Ps2hVNr0NBhjjoUrLPzWEJjQuaYuwoZn
rWuhkpNcDGX8QyCwC/NFx81yNeKQNZgKuHBUb75hHQnDw1eObTt/b6Lv4oq7wG+N
bLi+551kc98bU/DvRZhTiU20VVQZJBEnoj/593aM01GroE5mgKhQP7v0cr0JOg2x
B96TRKBt6W14vGgzt3ZNttUBHAF8uYTpW1ac+eF5iIWFWrIomD0RnsOabONHMIhi
mOCPAyO41oVJYRdHxmNKHCChmq5ruRcwN4jrkdAhSEzbTaPegeteZEI64JOW62z7
yILXdLAXhcZHVFxKpw+WI4hgKqvKLU/WJNDte/opIBbgu0B72EVdtJ+B2Hk4moNj
tZ1ZgoiLk6pwPaiioBabQLERYsfuZGjV2SzGuS3ot3DS7NjlRkSDKEiJOC5Nq74A
OefLtdmSri3eaUMA8Ho8bEU+oB2HqorkD0eu8k/uLShlOrB3iCsOF7K3r/J48wMY
e0gdItEPmUOW6f5Envd4O9Cxk6MUznDpVwckgWPf8DHnXTb9Z+tZcqpB83bdZQPH
6Ns6rP57cAiavwdyoTvNytAnbDbiEmwUTBPkgJdorqAMYmt4fn2czhx+N2Wwpi+M
kpuXtPSRUZbCX00oWft5JLGCMNRgOJJ/KxPF2JFXCJAVcjCeI1Y67WuXYedbf5jT
MJhn67YWjnQ2oFGWgNvxrSZI8fqPBL8IqpQQzmdHY0BHRSTNFjcBJj+ZWQVMAYj7
TSpolLMFjYgb8qEjW1O5ZouwgswfFWbzqh3xufSHu3hpCTk6GXMqGaLgpoug3ngD
cPQXP9jLauLBGirJLRV6Ns6bhTNosgizS9n2Sq+rDsWHiQ0R/12jox3bTfHVIE66
0+wKh20srm90DSQeHeV9xxJXzcn6JkxJkVGW+i6A4V8xxSvLKKKzi8hIs3Jo9AC/
jMepodJN37+XQutuCvYUsXgKDVEAx3LGkvdtBdqO4uTaonQUHa4Ggzfpw5Tzvefe
4M1MTixF/Mq0r1f5C6rn6iSKsUKGhOGNXqlF03ZTX4a/q8JF7jbIDOLOwAbLONpi
lsrOD6VimHbA4eU674AXi73Cb6zR7F6dCjNiJtP0p8WAe1VzktfTZOeyxDjQzUUg
JZ40ef8vOsPgO85PvQ3ir+biqC3apzpS3p3dxw4yciT7nsminoK3Tyn/TETw26Ap
eGjKzFcVOt2yfW9xOGKfswTRL6WjTtl+4lAwhybBkR17U/S5Y29U2FxsXySyU5vN
X0ILfuqq5j/sXIBedPawMAjGUo2deizP6vykDrx7cjR8us1YNGIq8tk66YhiPpYZ
VFSROUdUbSXd+FsZja9i9tnG4fx4m9mBxwM5NsI74i7V2fibc+o3+JqHsIufuCDa
BDywWo6c8zGBpKboD9R2SeZpfaiLVrM/7/69RZ1SAQR9srzFpUGWLHqxsjdBF6q7
9+EdJTPxxZ/+m/JeCzNnQ8F9B51LzKwG41xkf/rBZ0iQ/kr9lSqwcUJNiEbN0aIm
UAFszPy8Gs5M5r8j3+xwv+mCUCU+U3nr9F3/xe70t0yJchQYr1VLN44taM8GZicv
dlF3Eizypa8d5rK9Fsm4ZaztTgO2K0++3EIohIS1fjWPDouJsKuzJf85ww2s99fi
5ONjk7hXYGRw2VOFIfPiQXtbeXCRsPChA0EiAM+7Ox9DAMugarxInfeSJUwKYArj
/Di81+0VG190hX5EvPUM42Als79HYfDp4pXOXGMZWqI8x7btcU/uo0oV4GMz5TOn
zRVjRErbF3L9p+3yArQaH86xUCcx3utUh/OtIrSjT9biqQoV6i4pDj8aCqO07zlA
GZqqU0SPLw/m0KOc5x8xa14SqSSDeN8CuQJVGUS2f6BrGtu8dnCfECNQ4AXIUqSD
eVHUeQPNKO2qlE8WoMa2hDG6Ed+Fi9c1Wb/EQhkyAKZYgUQaK2E7xaXGtJ+9vsP9
dCtwaw5TF19AlRotf4wzvy0V0Iimb/76VtQba7LJ9ZUnDmZcvwpXZDTTVan3dcum
WRLMO4yVOE0BsNQJZ93FsWWVO08lvyvhP3VBOS7hNHINAKfjZlTHyrr87VFIne9Q
nD4dyl3b9inCbqdnRXXBhWcVJ/uE42uCZKobUcx2S1N4K9CYgZhkC/v/g8/ufEGe
p/V34Kq2ks/mfRrsrC3MI4LtXXTzyKylQyP+0SnLCWCWhVeROywnCUYbAuQNGpNb
i0nApwc2cZTFjsoXXLU4oXRmGgkeabEKbKfZDMub0IZw3MHvAmObmLJ7uk9nZOdV
mmE+gvFSLiUUgzYRsr9GTVnv1H0tFFjN6ZhBVnMw1p+yS9usTLaA0QH5KHGqV4Di
ityEFWOmQ/tHEK9Ex3yEjjWpQ5pncRehI2TJm6GPjNq868nhG/QJIHUgqx7LMEul
WDRE3BuPm5Nw3UutEhZrZVf0jFfIF2TNlI2NX18xHFoUoDJU1Mw/v51yUhZ80CcW
jfAVu1vEvKfac6fGqOk/EI46jhlGjeVlRuPiykd+UvOnmyWBl6pidFdcAztxuM3E
KrykVCUUQeMrcJkP7/rHa9ogvieDTjf4jy/A1NrRC1PM5mAZsVexEwvrby73Xxlz
bLSFvuS9RY+B0IueOYz6OtIzSrc/uUk4R5nC1gCM3o25IT6Bh5xrCQdyRVRlU9zb
rZgAGQuHOtmbjCqVRdtYogrDfQtcyH4vuti0GUgGJeLGmvwTT+kFyw1cH0tb3C/c
wVNwkU9ZJ4JHcR6q9LTzcv9f8vuZs5pe21sJEfFaFVtD5gA+xNreqz4sM8b2h7Zb
eHBLZRDMdb3neJh6m+dGC6IZ0YztOJ3iqZE/R20L3SYwy19Rwwm/yXo1BQ7vYKHK
471LlH3wpnlSUyce/unZ4G6ln6FNRyjcCTpLqTfNmBw7A/H45sLMasGOcybYBhKn
S9b9V2KGKtN7Vtx61+8wKV+1Te7uRib4bSAFAuy2wgTISLFA2Phl+rP+MhGvTkSd
sRrSa/H6H2E8dnb0GSu04mlyyUG4jx4FDjsZcJ3D7A8mE6Amngne/VHCrgvMgjB1
OixFSZ34JxfmPwDPfuXtfwTqzACI6kFfHyKg43M3EevwssnL6c7MG+ECWUFBeGoa
xRS/K+oMfzRX1QmGlikJOAjHBlWIxguJi0fjDIf7JQ+MNuW454hMe1B9WSaJ+0ol
d+VZcFCvDqZTBhdoXptFjxgUZArdF/QxrY0HDiL0rap1gYtO19k/G8/csWNHMz5R
vJUoFA4jKrWVEhXMv6+G+y3IUfSeqBTjmBInL/Z2MMYaUy3YVDXqDcukJfAfvCsg
ufY5T3bWsNrXb8HWd4E4Aa85ZmQM2JffKm46JwhxD2Y+y5IjdcHQhrsthjlcEjip
gtXSWJhQ1eC4ziOcApZmlOocvvVdrNyCGJxfbU4BhUC+Neo8CDztEsrEpDnaYk4t
5cul+CbGqtac34Dzq5yQojzqC7zTc+Q5Q2Hwxg6x/tmkqaw6xqVJcI69JEY52L85
zwuAtKO94sJJCx05auVhy9f022buapSZfX+MAbSngDDpAdRjvmJkLoz/TN1p8lj7
O2iGx5buqDU4RtvKXwYkQFMapb8qrekwk/NWgpp4vs06KH+Adr2PMBZEbfdOLPSQ
Dfvb2gQMDAq/IKChhHYu94VHBtnA3IzA2YMW9QaFgxHZgzj7WH/QbBMkj3M01kiw
V3buRL2xZzagfJt0Oj9L2tljJxdvmSHfuBHnHD9Oc4eMPqiubzaFE0N9ooxUU68B
X555E8GBCN0Quju51eFk2FQpJ92t9cVPVYLBZxTgLrfarwy4xNyk6ZkXwngjt2Xk
mYY8uX+FDx3heqjsGAW9tFNRbzmP564rI4aXBS9FrscVSDzWdXMi8/uYx/jnEez8
ncr9hZJyuD7ZzL6WBsAnhZFf6JfZejXk8Bw1fhMynPVQCKbpbjK4rbPBFMp8TiJk
zl2m/dvxaWJtnvLNxhQ0kSXgGfstuvU/uJNIFiyH8bPYhRIV+MToXOrwtDhqnAHG
l17lZOH/GgFSM2V1bpCaOVynue0yxIb6t98XhS1fvjKVDarSekDrdHukSxbRehAo
6M3YCY3tPDAKYgoTbrmpiogTlXeZk2MAKBSAEtJVPK3RBpEME5Z9yyq9BYPdXW5X
3LVdk8cFAGtgVnAIu7VUH/05ypBJoerTYXQVU5p3NduMh80uznZnWz5tz7xbK/mx
Kz8GL2A3nHn7owG43ZqBAEHr6UNT47Euf659Egxk0nva+RbxOhfMQZLVIdaIDL4C
7/4FMODtVPWgoH+0YH4K0NfYpOCDM0dlsZ3NjbINUcZ+mTfaeNFOwckcAp+Ft4ps
aUiESLtLwRzLiUplVvka2Ja/D1vpg/v0vmKzUTxUQrGZUYIu82mGynDBe+ySSGdF
gDtKlOWNT5k2k5inNxzKHvU3G8x+q7LR6R6Io5OioJxhQDKaH2YS6VQpo0D5HtzA
5tRKxc1FR4O0XwuR4OXYYK7M/D/IhbyhvvSiBnNPAJG2ArqId2lh4dEliO2aKxZ7
cfpHe6dkCTnXy62GUDQ+Try2Wz72/bwyrU1UsVdOu+zD7L+W/HJv3CG9lKdBhGi8
v3j22VUYFL8aO5iDH3MU/qfC5MvphLiq8/9lABIctWZQ2AYaTKAVhYlYVgtrGC+O
17G+Gel1wGnGvz7PyYrGmO86gVeATpMu/3t63KnCEwmtC5koqwiFvEBF/w+xgMuM
+WhtSK6x0s8uF8k1IBzr8y6yammiMct5GkDzr9Y3+rEVfRk3mGhXwUDjvvzR7G2P
2ZLK67iE28FXjPTYwSi5QXbomwddsCtQVj2cIq4NOeIr8pBY4gDksXsJRvGcogbH
i944/coV683givecPnfPNC1/vNwX8ygX4mWM56Sxk5eWtd8Za5FvC7JpXK79D7wi
YQwcn1CJ1ygB1kpuZg53ZemrD7l1U3rmzsqFtY5Kz6UoWKTIdL+FXtUmNOOHnDe1
bybaRu6i9yblHxpi6T8VsVnEoIZAwidM70ntMQ9wA4mYEXJntBW7T63Ma7DVaRMr
vK50dA80SS+RQ2CIyDPzB5LWDt2HT0LAjDCdCdYHieFVku3d1zMiPnLMXtXrY5yy
IfwskHAnVR85Fj64vQk7AMZg1uNgwfBJvrwYeXpBJAeOde733fNxvAK7uEKe6UVV
QyIDiy9yw/eQ2xuptTKITFihn6LTQ4BwWd2UVWMqZMMHhVUYhvrckv7MAud/N2si
xyzeWCCXbmNOAVO68nqMr6L2lsjvbShzbuZCnP0eVDuUW6tIOA2SFC2QAJK8d8PA
QSigy/N94FcKGpiApzEMpBFdPSPcVeofpXR9STc2oF6qhAwUgmxAzAb0kmvgSQG6
MPebFzhPkV/Rg2o3T9ikjgxyRVl+wxNfJYcpGBZbZ/K+2/F289Tmm11lIJM5IyoS
ofVpJvenjeIwS1DcJ81LbLtJ1BXS9+mAxSLZLZzEnMMoip6y1kn4pvznMrR2Pi7p
6QUi6Sbu70zq9XKF1jkUMzDUPixNOblDVm7aV0qsdNx0cja9SwxENpMtpjxUL3eO
ozAPFVlT4cSAN31pyC0PCtNgKVK20Zy8Tol1O97L8K0h5nux9ndUtA2QUjQc94ib
pT29lUn6gc3xZxrpSjLZnh6rm9MtFr5dW/Dbl8O+cfH2rzSiwWH7j8BqZ5ebrX91
nCj0/5X6kHD1p8LCC6+kcTrV37HX+Lea1zTHGgbOlkQeIk7v8qbpMeURaV/5cUIv
j7ONPw6lEnHdQ9rcd6zwfKv2tsm2JMt7/sE8N7+MdFfNR0/tJVhFZRq0PFKcHxRy
n0tDk+LBoasdtsc43jq9bS5dfaUqeRSjvKHI2wAehorb7yC4qQ3XesLtZ9kl6Z9o
6I+fvU6/Lrc46oxd2ziHTx1KEMnto0Y62ZGV26MIWjttotLbE1JLtLMwaf8wbxbl
rsXPklpHsbk4kItDxIkLygZWMQnOXEuc893xtD387sAJCXVl0jUnLaaX44GyORz+
lILUS+p3SnTW8WKYKT7yx9gxlAnqJVdPdrfs8ekuu2etDPovbuPsRzgNoDztAnMB
sTzmdGbz8MSp9JpvQtbaRQdY1c3qc2HCnDcD1EQOhscKhbyj5lzlORdWLRe/l//I
X+dadwoiJQj3DMvIs1lsf/tpTDKmvVEvDOOayruH93XK6sQijUIc9lsLjRHXx38i
PsrgwT9o2BfDCMuTdA2kOcMdcbIxxUiDMA/1kuhSHxOmC3MIAdElFCCdU1BbwQT/
VH9ZUwV/0tT2xn94rbOBwJ1JTjDD2POg2wMJcPdzKKcJ+Ohqo1wVjp6ICSAg/MDX
H1bNmLHuF/yBd9r2JkF48dV+swm6zOM5rZYPo9LheC4dFfwFIjo/CenHE771u63a
M6bRk5VhVV8kS4vIvmHaWDtBz06Hjd8wKS1IfXtvv2gqj67Y9Rf7fWRCpnWlneQ5
Lg3ohz8wrwN1PDb8jIjdwNvxRXhEYzKdwioXqY3pqaNAw5RcfoqNfq79b49GvlU7
NCKZ/R07VrD8oV+KCUzuaeoGTOCGLLsd6Xi4zggvWyz3wzALsvXzdKXKRxPBfg8e
r+eHbgRw+yhJRpZQym7ViNwYZTjXtqX97cng+5ovlB0/dHm5t2npVE51SOOrGyeE
CkAsqg9WIH3JQTf2mTsa2uNe6c9eCBhPyJNNT9S/H2ij5ZGdNioLkokaQECNSkwt
P51oHI7jm9DAlnYyPNiO0mIilmrWwh9FFQz493LYiGolS9uah9Rpz14P1K0aaBv8
t3iSqZdq1bbGX9V7Pp/Va0CeXVlE86dMiAf6hMy7rvWtjDUNA6GxQAXrrEfP68dx
4eJq5DvPnfOvWnkIeN7fPe678QmBrwWpsrPuZOvrABqeBVJ8aFJBOPsaVMPQgnQg
OWZWxrvIRTZmCMq0YdWjgxEN9ajCtz9s+e211wGUnce/5eEegJ9roajrX9rIIB2v
ek2IdQlfEHHgeQsiLAM+8R8WFkhTU3MRJrvDdtViHFdGamrwGpcviGBOQCUdxUlv
4zrgblQHXsFSfSJN+bLIxZnIw439smU1DYdXedBaOeRXneob0duao9vrCQDobRaH
gjtwiP8wPdStkOTBCajw5/K6QXlNWkIYjmbVlg+tbDGBJUlisXhs2/jkHR14k7QD
q8iyVqOFA/JTyxIjyhvOF142VwvV1esdz91V+73FVZT0b632lzFsK+fF/d8m/WCS
H+FLIl7Q9xA2riGQ8HlcQLnaqtUHfcXFftl98CkZRtmVSwHS/uoNR6LXQJcBn6rm
CzNHr84BxhqkR4FvuFxQqUtehOY+VfcaBN8jvZyM8hw/jx+xmvA3+V9vMBULsMHu
rYjpP/v/DwX/T05zYL/kgVbo+baWZ6ZlC3YRJGTpVXoLJVy+hiTOylVE/Kb/l2xA
mVhvvo7lIFqbADJROGRw6JV2FxWt8kmAXf1mekMIEWvZIGfFQ6lYC2x3sw01fIyF
Pjr16x/mBaSC5lAK98Zt30NOiI1j2LPcmZvRO6g+aBnyTzRml77ITA3Hsi68AmK+
L435XjPNW1+pxNVeHiA88RX4HfSFTXH6DeJYKQFIYeiyID3s2CT4HOk2AxMlIAqC
rBEcLeVgV9WvlWImw0eldkZNv1XLYkOW0jtOsvH/aVq6qm4rjhROu6Qpiy37HHoQ
jcZ+bqKCR+qDOTrCGrpstlczliKUmGgGM1Ir1VHOz232o+cVN3x0681JG4sixtMC
KeqrwuGPKauA+cXMJkFlA70JjVxvKc/okRLjRbaQoXQ3g9VhrVZPn+mXU+dC+Syj
fySw7CVU+gYMPHAXMpU/xJf3/7sPUIBSVQIlMxUFQ2YGfoXaB5umc9GVpWA7LNKi
U/JSCxNTjvyfkieQbV9Kk3DqMpU51u93lGohw1eTjeErTwWZAGmBUrw/NgzYg7wS
q80+dvQhOQRjrs3x84ER2l4RTle2bhnF3X2cxRSoguLP9DWHAbkhOEzXnSJHJ5dh
c76Bz/YR6k9IvDblMLSg+Q+QI9B6HeDaag0mvtWmL23kTwbRz7KhVozYEg497Oa8
Z3A9uowqDBD3srRSvzI7PRl3Bn3pfTJHbrOuTJM8UI5YgAZ03ndRMi4qApzv71do
hmgdP4VcmHwMAj2xJWXqk0J7jVOPLSVQfcFbWevoL+GC0WSig9slJBEBJfF4wwWG
BWoKML1HDb6Zg2ih7Ow5w9atMjfWLaGUvAgR12FCR+rOVbcf1q9aWjGI2Kwpgq+t
yWdjQaX8pQPeOUJV0p+i6sjpAOlYHvPV7LnWqM6kkWjsbCXk5PL24kGXgc2CkGKN
6ZvTnb6SACuUkYcIkK2l+HSzkFrLsBMx+5n91J64pF0T9vIVtv/SpXmcFaDNU9/U
R6UpHLujtQ+LJjqjCV6HRmZxxFWrt28Z+c72IoeYFvVTc17hYMwI05FiRkyFyHJu
FXQYZa3PE+z4/9m34mqM5rlH4sK7xPubDX0rcMQx/wfH8/LN7sd3w7y6SZo3bj+q
a9uChyWuSjeT3ufoH5Ypy/fVBfiHCsC3nJBiYlnfYPoPBNJ+Xz04o7S3qSERSXgl
Xn12yIjrLy6nZMRCFEQIx8z5PCqWcbN0OEYR5YZks6wxp3xmyOvYtQJCrMJKQ7Ey
HbMIgFAJyf8vLTeRLKbshFwjNk2OOBDoS73fDlo24D4AVI4JTY/LOXFvMOzQW42z
hO+F5HQ3d1nxgkPLZ/hNj0K3f/M53FL8BbsQ63V96Lh82Sumsj+wKYkBg/g2orlE
REIaSl8DbrbLofQi/1YghOrU/RB7VI5eBkuMivM5aK45jdRVU0+DcKz0tOmLzsxs
/FVw6Pr5b5AhWghQeyJTopO5hDpFSV75Szm/GGcN1QhjhA2nXOKJ83cTGSQEQ3Pj
6b5Gpy44Bg/x8Hs3r+o44Ka89mAZtMQpCLefUNzRL/UYbqhSIvKE4/yqKp/2kv5G
d6bJcdGAWVwSNEwQuSQe9n1i5IkrsoZ1DmipsED4Fybjg9G91S+pX8d+KE3Rxd60
uZTEOSyjXKHgi677Gxz0YdJL8KdcgwLKGbuGCcGDmOVgs8BEbnL6oqhyeDWkz564
kk4ItblnGs1S//HRWXU2kUJcg9NRDc3TSYd/F3deBUoG9ibMAzGfVC4x/UFdJTqZ
Z/3mqTkwkZPA/tPL8aMhs+7tOVoTHEdGM70NSDA5ejwJ1VkhvD74Bcw1My2Ztge/
QRRIlnU34k7Uo3W2qjZvdNVBSxUR5874XQWTL6uY3Q7itxtzR2RJsablI/WkQ9BN
F+rv9o1J4X1zi8fygP19z9KfUv3vwh0+bTqPGD4fmfTJJfE3zcKhGt61AI+ZmlVg
JcavnMjbP0jiT9KdN5BpdDGWgrGA7hHe5Fx/3qJrAFsxcknHZiW+RA7mLBeq9hwS
7x4cGeHlvzjhDfSi+3L3t3ehvXapD0d7uujWTV9z1hjW/6mkPc3oiq6NJHsIi+WW
sd/o//Y9BTNnQEf1gxXcJbgbEgQ6c5W2pwTbaKz4qvXCHHPxEuly6YkRi+oySJ3a
GophQDPo4Mpxw6YovjOWTblwfZUCH7HGMfKr9RpPaW46/do4PhTCzWK8sij6NMMg
LObKw12OTyaLvCZIxlBkkxjaMeM4FYkbjW/4nUtgkST3YAxuhrkHry4IwCttgPOg
QYf1dge6jeErDbSTayfFrzZlCyicbYcQmTeO7B0LqsMw6ypyAqdsDKTiXeCqFf2r
IQJBA1r4bPxPB/SA5TJpLUOST+26D5L9d7GSJXs/5XF/gt7qN3Px+FFr7WdLqka0
RVsHsOfhL63uRb9lDQUjzHm9Sr1cjj2AkWoJsl8WBnlWttfdHbBNhQ8ImXB75TFK
hJLe7eHBJfAKvny8C2nNrGIB6WsSRqFXiD/k+0x/zEMum8XntQ3V4ZDdK+DLIBhU
oDbGBEbhxqH83ceLV+YTBZr5myxi3bFXCW+cBN4DebgGf6lTn+M8MbOuOCGVXrS0
grN2g1iPVYDKEtLwE05PEiuLV4EaTGO/HdedMBrjUIKMBYCldYrLmCWLIGGA4DrS
2/2e8QUARCE5Heve47koEanzZBIxGV0Ey0exEao+8udZdbWcm5vITRrIwUlSvMcl
mBz0RHETUnmfBwJCdVEb8K/UzKEyCJnaij3SLqlIrOTvX6zTJQYvlL0Y7x8VkS5u
d5zjQ4GdHPhm7AmAf6aMB66Noy/yUhGyrH8GwMOpJ30ih0hEKEbOZ3w0WCIu5GyG
w/EbuIXnCoWAeWKRB2eQ52Swi4yXrLaE/m5yBc8Um8X0L+PlcVUF0o0+sEEj3XKr
uKb75qo9DJhuJRYOSg+eLyObVJ+Fo8cBqauhg9y0jQsOeyiRxTqj8lemMmDqGkkh
JrC6YeVtYQ9PXVB+qKwfeQgqPRk+3KOMcPPJwkILNqqmporVF/ulIBoN/MyfUgPb
EjgoieoFfzXFVPvNlBP4kriWSBsI03dmNY9DOb2cPfLuitPIESxt+2ZtSaVIdmlp
vC8JGeXWq+JcNBdM+C4+hfN5a7FS71SCcikP/zQvr5wTATqP6PTHyfN5Dqh4TACw
rbV9VzpZYtTOz0EgirHyVy0/8nhI24RPZy07UUEDiFVfew9HO4mZ8c59AgL3jrCL
xPMUBzwjRzcvxSIx9CYbQixgbUtZ4dyEDpk8yN8hLIg0gRcAqAMeBVOc8fltGVbN
vOqUutXi078Hkm++PdZoduxDIdiz6rWflaPdcyBVwujJ/5G95S2zyq/AUI05pxqI
gGVm6pVBv60urjQcEf8D6hwFj3WkRui7hMSoKVcLD+VF3w966SbSR5ZobipqNIej
LD16y7g7tnCLDZnmGLBUmhIeBmSg1rc7qPAgHMq6BKzia+EXbD6RvtFr00SPOCg9
7rThDX5W93IYdzSE7TJVySEA/Djr5vmgo1rVHTtzeqmcHbTcZYAhOJ/BCGLOQRco
0pEa/0QT+IF7nRSe97X5glCujAu45OxqEqS3dIYhXsghRi3zgIsZ4dIMnc0RYneC
Dr40jWspTwfvQEsq+8SRt/8woUwVC2dT9yNjhHe47kUO96aNzV77c2tbTx14B0aj
WSuamHspwJl5uUtMLH4ZVryL+TrYQrrcmFad1p2AIYlDEMu2ZcsIOSaVGmp7v92L
3PCZN3nilWeZcBdFwJepYWFqI1qPV0F5EqZtJpQ/W9fbPY/MLTFCqXxngC+UsSJq
yGokyy5LyX3vsZg3AxQUlrbiN4m0iGaZA1ksygjFCej3Jt6e+k1qKIAqbDdVZR2/
ADQ1e+sBQoS46XC2MyfVMJYmtQGqpkUQ0Ui8DQ85aHpcmezVZDmtSmac+3yoU/iJ
QLb6PbxA7IebB9BCaMXHfq4OrtirPy72IGyGWYQsrPpFkHL9rzgELHR2ADDc6PT4
uPKl0BxgyMTnNNKDMDqhZaGq26XAZJxb30YF0U7HlOf1ovmfCyPdGQGBYadu4orZ
Bi6dNrKaV1yM1dkwrZBwSyPqQWXOPfeHlPRxa7kvYBTLmMa3twx1hoL4tjY9uXuO
89nPCY8fYTKSt3lXHN/xylG7tyoClMWcdKQreWZrZJiak92sikekMqxqX1CzMXFT
jVe5lCvNQ0fWPl1tvh3Bb44w+rm71I0nofojrx5mPzIX/Y+b17ynHLkfXvXxmy58
8MyedDBS9UHwOyaYv4SyAzJ6WzgiS2AHnlWOZz8RKFRMbGekIc2NBxPDy0fhSaSc
PauVoazA1mGi2oLumEt+q44e7pIaeZnpC4X4AmhwRRNt5LGesuVElon2eEWiUxFO
Lz+dcN9O7QngRXue9SViO21A2KDIzL12ynjtaA8hP9BlciRdPDPU+pQVgIzN/M3d
sqftogloHRuf1vJaItsO1+h+yz9FP1Rd6QN74uJijcdzc90NkjHa/eoLxuvgQKiY
37GXWEr8RnZk6180NXsoQZ32qm2nqFhigviotRPcaqP9IjkI7tPOdKNUVVSugKxY
ujkKfzFJm6LujnGCLAzwx6sYE/lm/aHf43+6ec2TXZAbSvIWz0IuMzZb9lAq9RYd
i+/XetNd9C0AFHVnGiC5Uia5l/O9yOXsVoBilOGiRM1smk+heeiYOW7qHQURSFRe
oN2oZyy79HFOWExqRymdPI719dRbGD8Ueai9cdJEFZ/iSCmph84Zogr1pd19SXEt
RBykKfOPlvHL3aEoSussO7uOcAOxq0qDUljE0iJ8VWREe7wde7iNSyUcdlw90pxj
ImkYTSklK+UcMs5Klfg37DTa7aBBnuQBD/LPUNFnm7gjnHDYPcYOHcbTgTAxcHtB
AOJPmsCGGfXtmNPN804ZR3FyhSvmHYGhXcmAbc9ZtxFWT7x4LYBjTTEpeD3Vt+Xa
3uyyfiBa2SYXSljkyX7PuZoXMjmwie7iuSZUIzwr7nojLbxMFr5a3sV/pAz382dB
TEJPaj3IvM/rYkm5v1/Ya7LWzX++AJARpeZ1ffml6FWWigJwOKJGynyQPVR5+I0d
lzElRnTtDH0OAiqYZ1doXrj4Mv+snwa8to9hQJDFv25ZVHPHzlXMmFtgcmQz1ctN
4QhKa4eFEdrTJBVQTJ+glil/tUEKOVCoaAMlqmm7+3Ct7I2/fVwg2lc6LI57/2aA
Uq2WnlZQaFljuVQ7uIiDPj4/+i5b3tMdRIAitxPCH+ve6R1A8lF2qdNPgJ3+cxQ5
chCar23PbyO/B8G2+av30tBTdMw/VqB7hdbbuhSZelzuxKOFvcgZjiGpHqacQC5c
6DHledOsVamwp+RFwpUq5cC57zN3A/ONWhs4VZTqK1IGdirPJN4v+po4TwGd8AGT
Gq3iHM335+ywVQlfLm+9+xs8MmmrMOu5XdoANTr64XwV9ZdI+Tc6YMlSpHG+lXTR
b8Wz76Qn9EQoGQZOWJgBb5DOr9gS03KInqzslBSS84wYkeSSlo0O/Z0B4jXzZYpn
xsIOeLvcmTKzvkZ6h3Zgdsi4bNxqt7fNxZ1hToBqNdrMW+dKcFEeX/jL2HjHWy9h
bevse1q/ThN0KcbCnw9g/h3e1XZ01RyOzWuFvsLVQSftHLuWaOPCKHIO6EyT8rR/
1pYYUk5iErlS9wWjRQCQW0/f4bG5lvE7wVAXavnfXtbbV9JdiOTLNjDrnA4T43Dm
aCC11KDm4PQJtK/iFqV9htNN5YsYErCThUNdTlxYfz6A7w7/DlAQ8abFromJpHB4
jRc6PsqH5/QY+/jG+gwWqduYcH/u0HZpP9pfB8+e0ZjuYyGlnPXRY5CkK6rvlBLM
CdEzG+LPYUdw+kVtTw5Px9GGaLAAZi0h6lFWRBy+l5hGAohJU282iXxJhUjyE/VT
Ew/UGUnDZquLnqeTCKlj4HNTbtgc1LQtsIyaOGKzQULl7Do975+6DNapXBS1NShn
SZF4tq5UdB0Je30NQFSDniJaQzQRfbMXjY/A2w7A1uqNQ0O/uI2k9LpTU43j0r94
kJI5UCARvtv5K1LtTj62XYIqLt1mml7j9jq6giSdxP6nMr4K744qsKsG7ubqMGn2
RoeHaEf27W4dhdT+6O1x/zLZWxDFfTFCTu+Hqc5qP2aiCV5auyg+sEPUY0FDdAPI
TwjnJodPL7OF+Z3GBZPgsQb8nk40xrTVqNwfMwFMbksfScFpHu4Nec26WR3tCXCW
CTbi0mmXAghYFJ0zLOmoaN7WH8JpyeopL/Pv1Q0l9uB5VJSzgh4qegUp69fv/GfY
3OBdBUUs7IhnOnTKF0F5l92DbH4w6/xwQ41GNrhOgI/9nnGyLO+jl9gncC+1E1hE
oQ6K05dsrzJUDKWBYCOT/cc5IY2S48T3B2HUCamqyG9zYYqFTTnlbEPdPe0e/oZK
nw6O+YXbhEfQlsyPRwptc4/awaXVk60QM/ypAIa4AUBVQoA0oe/2AAZ93OmkKJbQ
GgKTNKjEgJIdsj9j2JukhAN1a1R/QQIUVXrS2mQ+1QxFicLuH6Pk8mHW8a8xJrCZ
s1SZ9DVQS5o/OCxE9eqp8UAk6Tau4dB9RIErFnapIhvSoIWrFluu+qnu9xRNtayb
J6XjLgTCU97w4/XkeCbQbweUs0rHsAzQRIXXHM8y4jAvOcTq+Bk9vqOsEWaOZCW2
5G5PQAZQ/dMCALSF7ZOwNd/qi0bUhoA8lO4qusia8i3GMFlbg3y8HEPTyMEnyPg2
nO1K3CUs5iInfVpEf9addiY/Biz9ZC+zfbA08hcPtT7ngpz1LGo5zsxthNl8LXTD
ukZDWHbNh21KuPKp7cCP8lmt1PYXicTjoUp5l0qtES6dSacSmWsid31aSHMHFD3A
kSH63y3b/BrAZ5gMmsi9lGkK4vwO9E2FGS+NZz8pQeLH6FFzbATyyvYJAkoi0i6y
SLSMlURw93Y8qM/uVmdPgmwVx4fuR20gvx7qFv1F+zWYwxo5xD9FX2M1LA1w17Eb
Yg5wXak8vsvE84wn+2VeHT5vJfXd2lUWrRdnkWDeix/GoHECNvMrEb0SZHzYwN03
imUOcSdsgdBqCLdxxkD2pYef6ryI4Yq5wOGIg27QG0+xbW6Lq+/WoJpX7e/h6FTH
7/HaDeHYDdDkoJH/2tl4ylxZmd5Z0VoG1vasvcE7ROvefJZNQqtM+TPcnHhyvtuC
HAhPzwwkhzvXJKj4RlaLqE+IZoQFOJHBt6IQ/CB05m3SyqbKXrKxMB+lNG6jchQw
dZrvntHCi88htE9WCOZ+OT8eze0MLNSPatu1gLQO32Lh+FMiUq3S6fAsRKY4xAp9
OWykjcQjqBbpuKLmQeLyfJaZLSWx+XFyXE8vbgQG+/lzmxFK5IO3LdekStBBs2J9
+vdgL+2o+g3Y3c7jcXRKTk0IS/RGi4kuk1aENPe4+g05gYRGNyfe19xp0M5ZisD9
BeORxo3fAacTd/9VhcqwyGb/sAC6kFpC0tYv8u4T2HBnI5k4cZhsOxOw9BPStCUS
J1sbn6hfai61jO4VSZreQVS5X6wM1jER7kM+btEW5YIV9SHjAqBEh2qx9pCbSx1+
66bKIdvfxpUD5y+pAJCp0pqdaVmdFX3dbKXZPCGGG0d27EWbqsapZbNQlFn98O5/
AjnM21ffqqBYQvzZppQujztBtl6KwwT5vZidKZoFcoRb3UzE1mw8aWP2GIWQ+mTx
UOm/UBbHSpnecLqzWj2PvkgYYtMtx8N909IouDoD+YKGWbVhZ7di3BUcrubJoXTd
zhkgUgzGyfy6qiBfVlfApKvJKlQKGmAOqmEQ44qGTeMIEiHDbUPI0HJyTvG3FR4o
w/OuCv/14fv8tKaXroIEtzNwU+hYPXlVrcBKOLjzExzTaL2mXu/AcN/H+5EyR10W
MKeQwnsrfkS196RjaQCw+XCvLa0K4YpASul+eyRqX/fO+7P5Uiu2vrVNGANxZSav
gZd18DJTUSaO7Yi+q36MiovwLlIFQoDW7golcPutfYD+4pILuyOhHSU/asoLLG2o
J6wD5CTLFd42xXXdVdT4bF8hZJFSrdRQn7oOUTKxrK9K2sglybKGNLA7FBgk1Mwa
S3jcH7XqHgp3WBm+AMx6p1VnFWv3S4e2K2txkoeF+IMPuIFcRkW/4PxsgsqvdqoO
NqjvIIdC5XjwqIk/PcR51Eb6thr8YS8xoeeKeUOEcKBi3s+Fu9DIorgome4Db1w7
3a2OHSWphfB01W019DccGo6F6ow8NlY+fPZu1JF+PfxNQgQUfufKyuQE+glytqtQ
5zggKiWIvInlb3aOchOtpEJkyN6oz8PBKcjNmn1IJocZklkbpd9EjqtD3oROskQo
P77QN/xELwA3KdVG0FFyv42X2vch9rcvNx3d/awf5K+LqBk+T38hPAaYWVCaMShN
JjX78Xl4papmbYDQHnEJGdD7z+i/UD15DFS7kNLBUO9FR5xqG3mZhuYtxDHoyszl
KHWKWBC/cratTaTFwMyRDi8+s1V2CsNP2cbuBvYwlKFMjdFYAUazD5p9RTOKszRA
3JPjCFPJZNXASAbArJo3F+YjZ8m7kIAxF1YAkswmfcEylavPPvl50POFrKMN6cDF
mGcPtDyE6DTIsgEVhdMw4hWJBPPf5UP0BvrGnldFNqMy80SYHChPjWRXOTrukahE
Ph+goTwyfoMrjAjxdMqSCPI1C391GBzNElh+GgjCayWiXsHxU3JN8i4T3qw8xO8t
+8xZ1wWZXqq9+JlqBrrwgiZWMRn2IDTBPmRYndBaEcsK+WN2pRIdrgVPLa/x/Q8I
95XOxNRWbbLZqRbS7KgOKu2QUdoE6TdhEHbFqaFA5421/UdOVZ8a/cZM0DaCq1rD
NMIuQEVuk9BH48qeDoCHW8i/nBuxFxjIjdtMJ/R1lfdF0BaxX9Z1U/e+ximtMQ1s
j9IN719UA1SoFH08adbU713YFLlR7iKPXflSZ22ftiYocle9N8gtSuAPuo6/zyWl
BFa2Srln7NAvMGx8QXqlCnI8kztcdb1aKlStBATRZuX1K6onSKZ/FTTq4wj8n82b
AvtNEQcXOMKhfKDbUUJ1pjfq2gH7Yp0kCoO+8DlX1OD8s0rUofHgOmkFm5ah1lLw
td1d9+ONym893W685585qsjkkXspdUNKIhL+djgCBfk2va59aS81D5wWYJGLQTHr
eu1cFj4QvNMhNztyux7yTjvy6AIm0Jfn8EzjpNdeWRPbfD/UsY+Cqnm+JturABd4
2ce1QhTyyYTlujShx4528iGR3oZxbbjjWXz99K/2jyKo2jQpw4omhim8R7mhVJXz
kjOj7szaRfVXT94xrBC7HX6Y9V0riuY0cLEy+wQRE7eu0FEWjTLz2Dg9vudD1+kU
eGUODRV1U6qNZ2IjKpIvxO5ZzSmUYvN/fN35sYBKEpCrZZ05Lh63aJ29NJlQKJAF
2Mk4RBIMRaXjMFJGtxrWwO+1c5ChPwx8Iv2O94KKdZY3PRQvb2wnd75F33sypaSr
oIW/iWzOzuuAxw14UDDNmSjWFl8AMRRz3+POTzlxiofHA1CcvigZVx149+TeLoBf
5QBPhZvQRYAY/txqJYVvzo2HyVyxh9Brmem0MbD6p5sEEGXfgLYZSnnQGghvMTZ+
r/fdAwsNeKyf8oOx5Ig9S6GLABoV1sSwbqpoKvoDYS4NPqyvhZelPjxX9oPJzz+u
Y+qJmPoQ1FEr65RoByWtbzjiUQYVsCcDdF+/l3s9lluimYAnFwNOS3VT6umoWunW
6dxAIX8s6jRyepuY73mTdw/pZrhAEJq5RjjlneIJFXFYi4v1UuB54Rpe4AxDGAmL
SMCY6iNKfCPQRP6UVMhLa2MaHUfj5bH+Zj1vp0EI4QVE1MQ9YBl+fszg+/Q2/xku
C83zixWAzsam2WiEXB0W7ZymxPVjmn8RvYC0vpUnnZaas1KYFDZG3pQLjA+1pmNQ
rEaQeXob5d89r41qljqb0Sn4/YLTAZteIriXkzTafF76ERCSrMxITdLR8HUf47+z
q2Y6kERTSZOhBICFyHBShVOe7HDS4/CqEtHTmiQh7VXlMEsmnZEKOfEVnjWvRkpz
QZuSM/Z35LCpat47OVctjNPQe7iQ3w2vMO7BrNo2o4uTbISrYiRKtTuSUBYCBAzI
fI4JnloOkejSePctyvyCiDwcohD/g9kJX2Ekq7FpANp1CcUXEbc2bVxZi8XBEPPK
62SuPxFr4Vkk50+ixTLA9bIWoADkzz5pOelilgGV9uUeYy8wa+OHbcziw7/gocuG
ICeE4WE+b3pGLy2EIZ3YPXuLv0teb9+79Tq+2cginv1NRHODuki71K02r0VFHpcE
8wYksQ/4/QaBev38LFh7QowSSRMDiafJDLfOKCLNOyrRnP6Jx9/tueAVuX9KVm+U
hIDvS8k09x7anx6pktIqsF5w3U6IYP78yJpu9n4Pbc6NJ1PKXeFNXZ/SwVONqfCf
/ZQWGgTnFG6F6R6xh30iwgL2PORwVyerqiGeoH9/ZHRv5ZJFO62YiOgs7bp9DLVI
UXrY5+rYFmajhLBaifhpTQporOrZX6U0RbeQ1WK8FKYxIF/5dS3Myq/t9NEk+Q1U
8MBE2Zqa93cT+jyQHBsSajdfZ2iH3zUnpsfs76VBEl8Tu2pGg591GOto05uC3mTd
ROqJDmqcef/utNjySQtZf9iA1k9KQcvHdWOq0CjEg4tkMCMohAWhqJGSFweqVqes
jHv8uYM7G7kJKjuknUiWi0HJDSY1Mzo/K1X9+ypEuQGYann9k6xcOp/wWEcSS4dK
XGxy4Nyc0azFTprrsGwD/V0lw8FV5uDzofZaURzBKN1fWjWMeiTrxLcB+5BeaKpq
nEPF4IKZrqsYZF/4S3NwRCRyBIIbPfIVPEkvYd+vW7Ju1xc9yIzKiOOmqzdwrGpb
MsECZ0orqOYksGXBcAUcuepFCDZbSho0KCEFpjRTv3CPL4XtQx5RKF5/vXBU/Ljx
/xMKs58BxmhPEfrCpiL/FxMOD1r63AhG7Kq3UTzWlkQdluBHDUFkH8mLcDkjRRvg
EklsnuK8fHy2lVOhr2BbLfGArjYN3bBiol7Z8gvz75WKz3mVX6ICt05Nngrmog9r
9nB4hvDODeBfZYjnOaP/29QGP5fBbPJtMVTTEPvYw5x2hmGmjWLyHfVeJeARnxy+
WI56r7c4B41q6SawR8duPWTcWw1+cm41+sRQ20Z891FsbN6QNRp4wpxEjMqIB0Xt
MQOa1z/aEabnxkNviCetTfB0d15BgAusmjyLKnkF9s+ivHmoAqGjf/dQ3RQnx7iY
pd6jCtE0p3G/MLQSLZ/uh6PBD9gosmuRCB74T27sDbd0o1DdJmqv9feSl73YsIsm
DKbUrb2rCnHoMqvfBGBLfefJqkgHS46UKLPjcwf/6x3IFCHAp22s+N+hdZkcdpVI
mk5vmGLLP4xvNHKv1NzChI+zKuBcDCl8Oru0NpazaL0ZZXwjk3tD+f0FtS9ek1dz
nSkG23geJaNCnGb3lIrL97bNEU2rxxKal4tBvlPp8qo/P1MTxDK8vQVdp1YnR+X6
nanlKeHs0k8A2CbRk57gfqbiA3rX3ptUi4+DdutIRMM7iL6mnJmCQcGljTggCXxM
tbyIRPt4h/xjpGyFEy3kIZqQV+4627ZST3EbOOnkbp6Vsr56Mx+zOoiWU2Azn6np
rdLI/8+DHjPCXA+IKJuNz+1oRm5bSR/pkEowxDB62IpAQJykN8m1qLcrZ02ELMm/
Dve4RCIyPk6ygc/Wo8PCL9U7aj2Douf4+htZYvDC2hEQ41ja2mhCCtcQ0ufulmef
zqITrGWCmyOCeP7+gsFY0/vKpCfYxPCr2IVIOKU0LGwZgavCDD+1e58+ZeBnRcgj
7IdJL6wSUcy7PkGc5Xd9Ug1BT/fTOLGslJFTBUv5OOi009HHmF2Aes/5ZZInbtO6
LX5HmXHmkEE7uYHKlVitxIddCXqshWfBRNQEixWFugdLhWqbS7jnDyvYagu/aqx2
XpB6YjrQJ8duYfzhAkLmN0kY2szq3EDSmKVGxd0dPlOKFG6DJjrtzlUscjqTQzEC
1X/P163Si62DYO3OxeyLo9xfLSOak16UGqkRwu6xPGCtmpWreCSOgfqsLWUqWSa0
gvZ7SkXDa58yyTixgTTYBZPgty3eVLcOIsppHUWLPlnsbQJHM0WnXWp6mCqSs5U4
KqwTkd1qlPibZdvpOfviOHUJE3CSDg5je3naZt2pWBErJ2CkOzUErF1PzfrjW6sM
B0JUa96oGa+kr0hMZKuU+1XeGgApILFQ2VrIcyukxHR+xNhwUiFhDgjFYgpZM8Cg
Xt3yOG4CKaLjORtJB/Z0q0/gkVsTbos4zoDKIBikOgZn7VdXNRhzzzfXjWsKEYkd
XrCGwMe4dGzxKEmK8h1+ZnnkzrLpg00C+lEXh+0u7r3Qad4XeAf0ObGF7lrUyi+G
F3YZhmDPLvECPTh4jJMgUHfBNduIPqJdMwh3a3BEmk+pFAH0iQ+nPwFC9EeKG7w5
hcEeijceh8F+61uEq3iDB/BqfbNVlmLwTgYE/t55SKyfojAGjuU4Te9dzU20qj5J
HrfKH5WM+t2WILEm4Cj6pkqlltLjIXvb3PL7h0atqadr6qF0u5uU82zP3Op4nJZw
OxqoLhJrgALqrnL8pizYVnzV03f526E4y1evsFR2dehoLYaZkKW82cu34JNRYc1Z
u0aYdecrH3uXYm4mt9WiabOde5ftDjmCBx10F7JeaxBwk9mArWRuu95w4MwkljVk
Il/SPS/lDuPWTMVR3txO3PIFfSUcnTtrE4iTyu6xu/rCMiPlK8qsSDqeXyvIZbue
Q0j/O8+kLSHYF/+OeUesoemATkJTr/dkpcMBoj7wGkWED8vWWdqqAv22q+Y/w3gb
lod82VZCEPlIOQLsiAAH07Q7yWrw4hetl1o8kZnE3MCiyC3wiAmuqeytps40uM2R
LPzm4rrsuXsVQiIdL0KCeTW1NL2JsR+wdnDmLvdYxVrj+wNmo05mxX0lk9TRoTnB
+Vt6v3tpL+smU9AUv/a56eZmuCyuoXIUd7ZMM/2XMJlw+lCpwMLLca+PuglE4RNc
sAdBHdUIxGMCMkPhRcjEHVz+yhPDiWO+JhqODN6BLVJd/rpJ5GONECc24Uts8mpp
RsGojs/80R9i4IRVQjcsUETkfgA2PzxO/wyucAAPGM1CI4W/JOOzZJ8zwN+RE/HN
6uzBaTkk2EolZHRAp+ec1L1q0xXq7YRNDvCjHwKQ2YZNBWcAq015857bJDz/O3G8
YTUfKQL9mM5tMTAhxLxXk4wGqsvIFLMCPUv0JfvFPLtY2Feq9phnzWdu7AVbGSQ2
F35PhCFb/7PB8VUr8dJmg08kWsEMd4tyS+ewHnDEQOmHoTGCTF42uHSmZ+Pe8SDZ
ouqo7lJA9SeGDrfVQAacVDsuskTtr4mbFgKVFeI/ynzQnrXL0zLcbtHp3O52yE+U
yQD3hC0n4aG0JmtJ+S3wRTw4QhA7shH9yvOIT+UoJdsJH1DJMxp/fXYfBG7xSp4I
rCVrY1TIDlemm9KCBW7f8MQl1LBI8OQIj84AbOjRUBDBdnHg2p/c2ze6R6cRpHII
97yAfpIPcWAKrJNROzI6evfP7RVUWUQ7URILnAi74SWHgPBFRadmCCfXB75y9vX9
yzJ4Koafcer4bM5daLuU7JSzCfhEpOaaVG77FqKFDBOsflW/+/zXXCGQvMSStz6m
btkHDAz/y5iVleeBpmZ9S8a49pHy7H89DKQn2REvGeLWizopEMAIvVVmHBqJj4JI
phfq/aG3kFkw+oWNn7qMJP7w5GIvNM2v8RHwHflpc17XBKdECDve9Bo3P77ShVMI
iIw21PJymCvodtwzFxTLptMWUfhiX6WPLBUNJxQnDl1k67W4uEcBeNn7efKpqO/M
7p31/PEhEHh4A7rNJAMoEAEkYEwYUEjeLA2r5Zs1FcgtdKA0z07T4VAjUTEQNFKE
pQJIBxontTKQjza0qa5yWOfu48LEf+ktZ8ApoAAJOQcwavVbxry45Mb7G+ZIPeEK
ztsGdQDoZuSs3eM2PWgVG0wb+b+PokKkZktfxQtUH5iUxiWe3UaGXBUvpyDeNXeG
4mqEc3dHK44eGFFcbMiuYiiUHtYSnYLzUttxzmiL2qN9IRvQ76lojREeCruwAqT6
J6pA9qjGhF/VUidz6Z5qgerHzMDz+x78ffSVxv2O/wiBJ5j8ZHpio3OZqWB03V8t
n/XsK0idlNSzo5fy7r3l6CmFKo4d4AZY1Bw9XESMvGseev4eWRvjhj7HsliWytSW
u+cdN1RK7Uy8BManHEFpcIcjASe7mpCoq/wTjpWQT2BEq8lfFUenCvIM3TzM5mCw
6kcgQ3ycuJYidiE66scseyGV6rlApm7dkI+ILLH3PLqUuDDrEqQU+wfefxcImFJj
HyWryiBqD8dstYkeao1mkZTvKc4AjWagwYe1UkDPDnxGHc3ywoFQg0rqTnSru/0V
/Q870VF/VJByfzwdHHNAhtVhsjggjhvn+5irMMucsRF8YDUzRTsF5DLQa4ryjXi4
AJjeEMVEEsLKnxn3nycOWVcslfZQIYTGUBJ3f7w981nFrRooOk6+dBlZeBmXgCNy
HMEhvSj8EQrSWmoo1B1kNwNZKevRcCRiIz2dxQTRfIbt4bJBMBDYBmYzof9jS2Z2
3vigArS3/qclv/hAPoKhjy/qTCX8jq+AF0rwf3xoXyKjjnsBK69q+xj91Q9KoDD0
NEEO5WKv6CE74YyOzs8NHghNoAKAQQlZriEA65OPC5olEYlZwI4PMxsS9g8dYeQi
592do9CxT2NPLTZsHSFjnvglVs2HL4anTMMjcP502xXYeRw0gLtAtDRSVXQMK9UL
ecOOeIRcjemGv6E/JC56iuHkjLJ+5FFC3vwssyZW8IuZz1w1sePgRED5G98iUmlF
9gFZTZ/Lrx8YCPzHR5eHtJc97S39WVrDpvlaE9edE3djPnw66ePl3yWhsCdGTTC6
ZMEsMXs4/vMOj312oi4IpGwqgujt3ClMaKGPOOZeLP9yvkv3nMFOGLbNIcNBiQFl
Fvsg0ihG/1yh37jx6Q77uKmR/pepXUdnkLGe4bzOyP4guuutC0dKMa+jphp6st66
IZIdeBBu43X85p0tOduJKRbfVPtcCgehic+UmdVLELgsbmxvn1FaEntPPi5pj9mQ
SwKaveBPTj+cv2VKouLyQue34nM79JoYx20lsi7EmIXvCXP092Qk/XCRcQ1cKGsR
A0+S/1HQvKPtp14sHnH64uAdTr9VPDqAUQ26uQVebxchJ3SnzrylGZDy5htSpGXN
tEyUZaSwN/D3SCdoLXoOQjSnxvqwQr83vMPbjkKi7mGskdE6tOn/DCesPPjo7Bn1
s2DE/Ebs25jvNB/TLnez8E07JMRM7mWjDr1fBT8iFJdVt3TAUVV4q+H9VIoQMFsQ
kTflgWbypEAfuTnpaZwbav57JFybWxNatapwxjGJ6YoFIBwAp7IyMg3vHK99Osde
9+h+jgvPniR00+IaYs1ujgfe4u9Gvih1BCk+S3B4eDiR/olSr5RdRp0hZsqQLUda
uhAe4mvF50TTxL4rk2rOEf1w2AqL5aZRbCeJtV6wHQblQFM+4C7q72dsgBQi4ALk
7uYtHLbzTIq499xzh4Vo2Jh0MtphNH/Vw1k+Kq3OYfPll7iYv2xAmY+qOonSsozS
kEU3NZ4I8vxsFZZw+nTZjIEbZsV7gVZ9pVXEspTGPuFWM6RW9ZHGT1qdUlAYhyd7
Hy+YoDydx743jyXzVBjZx2qKULQmY6NSTAatBAq9ZIVvABluVmD3IfL87wl68YN+
uHmQspBP54jKDwx116O5rjjO/93URralptlr8Xs1p9/qif6rKY224Rm8K1yGjGoU
QuQM4MeOcFOzhoLBqjyV5+9oCI/b5Pkqc952xND5lVZWRI0NA9Tq+8PZlSBXFvU9
yUMaU3h6sEIKq8pGsZaZT5fi+i3mfAU2GCGMfg8FNklPuR78X/iKrfWlPURIgpgU
bXvRSrLd49qj48FyJntluSNEa01RJt4ryjEOzONHaVzsL047mWPzNQ68MvXOaRIb
//5LRwDc4qp/L+odzUyU+d+JFltfC4LoagzHL1nLadKO/kwqjj1UNv+qRN0OYhuQ
p43Sqb05FozH4V4OlVmi1zl3I/gTDSew2/T5uIdnxPboOOx6A1ruMgNCrh6Jws4F
rikwM8fxoyUnF7QYHRPMLl5eefVA2/KGtNzeKbsCd/nqDZ4kuAT24kk7OIVH8OZh
BA7IEr5BCJiUyOVg8ngbaLMgahtOeJcsqlDRPlawi0iX0bhz2s5AAicbGdBGpF8o
MaJszbDUXZ2rd+kgEZ4WXSHNwO2gl9l8h06syIQRzgHEdeA/dL1ptyIwI06aMaIs
ERJatiqj17l8aP8cv9/X7cKysYszcLhEVnCUunnLnIBZ254NJgKnWN4smWqZmsnx
iQinawKE1YpCW4q2YAJWxfgNugAFH6OGPhonNHyG572E6hIF7dQeu5wyWGIDEGXO
AxaFw0XywhKrLmSkAh+spZpdK+Od5EYeomE5aAdVGOV2shFVoR2HhMrJtwvABOmi
XA7w2yce+0FmG2lF0it2eQEkUM9sXxvaXrH7si7OC8NaXzrNSPKj8WRWckQl+zp4
zta7sNzOxLaDlDXbnY+F7VMT+KgwooRpgTemLEAlrp7aRPbFo0XGnh9OAVuWdbIf
JNFgUiFTp4enBXrXJKFNIPupFgn6hC0rd6lRAwqH0n7qz/eRbiF+dLLReDHSrOC0
5v8FvYJCDf1aD8LDAfKXZ0OXcKA2811CBgPUpCsLm+pPVk+sDEho+vmUA4oOXkJ7
LTYaaVltVNI61hYfiPhlfTRZF0cL2ceegFD1J/aAg8oXsaDY0k4tRQoT68Bat33e
fN/E91PJXke3IjRNHVbfRjhMbX33ee08PBLUPrrySFukL5iaVwiPe4oByejePF7Y
3KIC48IvGiJZOFU6XsHgp5PLpL2pxrd/+DD50GOoaslggHw6ax1Yz9zGBHvP4Lbj
DBORxQds+nsjK3U40f6hYqwGUsHoBn52+7bYBwDxyWml7UipA+HvAuoX+Z4Q+0Xu
AfgdTCGImBA/6xzll6z6OWq5nJliAmq+wFqUnD42SVvyeYE5rwTRu8BpGKQmc1Mu
dqKrI6UhB32kL9lQnw9LiL3TC3lI4AHZfb6bgLN1+LTzjP59e/UHjnimATRKNrLj
CS8kF+JgZYM2+HQ1E1zxhLmUr3YtGXiHxq7xtNgOnDYrSPO6HDGrpfBD6XKzDG3o
Ojf2RCRPzj1Zr+x2WsDVbybgCwI1gZ3YOs1ijNMkVP7R2+0KDVt/XLiVPNm3d9ng
JjkIiW58qyJect7pK/UZo3J3FpU3MxQd1fSDyxFLKuiDfE2b6T+H/v9WqbhH/X0W
DFusNHql7tMX3lAhHNpzWZqLO+U7Nc3hYlk2nurJZuzEgjq82cPns0eoumRM+h18
vpijL5L/qqjo1pnzGGMpV7zTB2ddDE8vCDzbiMY89ati7kebdLwb9MLfznSMG8nD
cu0yrNzSCsqoAJ6IGDbDu9bGr1vlqQ+lVarFBlymo501bRw4TO/rdCfdZ3kt99zh
SSQD1yiYM7thBur26hx2drixikWl83TvD/aLZuffZQdiBYQGQg4EXTq7kvNVelYN
O67HR5mRSGggWeKBu74BITLMqtFSRZV33guMUeOA0S/Il/rWM3RZFo6bklZ34bd3
nKYg5GnvyiVG+wSJ98dlwH9n/+gAJenu2RoHBXv1YMyKV7Y4nr6eYNMe3neG30QH
1ioq+8pNt8Z2X1iA3v1fu4lOLvqwlNdRC0ion+eHc29gviZm6fownQvea0YjMEXu
ByMpwKVSVILmE45k9+6VKVLYmNg3OvCePJ8XVyWBwxuQuBpJ0DxmyovC3mJ43LjG
p0exzcMqSum1lhJDCZO/QTcAqgP5gjCnxziIGtUR1uQHb8LCqmDjRzTTbBylMUgA
+TxdPE/nbECVMTIWjwO1ATATQvnGJV4k/iqC9dWbDSADNCSdd4nlUnMxxR5dyLmO
qVNJJF5ZslbE5b1gAfTJEJFtxDLfNaMnAIqK6djiaRnHYWBAPG044+1gmJN4n/G7
UmZgzlBDvPahgWZzAtP+SXowRx0WpStPT9DBYSgusxSfD5KimUFO1jWaB7ruNM6M
3RX7krPs1aUQEY1NVsuLDmmQWGtbHiRSROAvEpAOey8/HOLFZkRJLFQo4quL4bGY
quEOBi4s09Pjdom4VsiOVKgpOH2xpoutyQVcHQV3dEnlJuPbbsIxn6ElIEhFi9vu
AvE9PIgzEyWGDHWzG+KL3PW9Dp6UOCH2D0bwCS/DIC3cso1a7N8bzosaM0P6Zrjq
t+A4ucbr399L+NloLzLHIrVyz7K0HkjjlpbO80SN8MTylTS/B0Y1Uw61bLvbIsES
vfckPwIZOQRSOfLR5EFLVKSHUJsubeml5GiUaS+oS1NP61rUJpo5B5WjzGbHs2HT
HomdO9FUiQT0S/Ut6JYk6Ttk0PY/amOQWkH4hwQDkR4ZxC1DtDcJ4sEDgZrWZrPk
W4o/pbPkHihtkrLk5mbvXWaBMbzj5WmDPkwkGPwT9KHoeOGRRmx865miNrne0RAo
nbrwpcwfLabfR/9Zdf16i581Oa9GRR2mH5EDahauWiogMIW7ldOAtCj4U3K9rOPV
DhF3g2dWWrfmsElOJ0Ji7zwvCmUhLetBJo5MIHYqenDFCoDchEa6OJ+7OXHaNMZd
wFZXbM8dgMzxQ1G+MwDS0SA8FQceP4ry2vfVGvuV7dGN9cjVeolDvAOnhUH4kKCk
qCEn+VMKHAncqx+zfjwOSq2BEvzvEMGVpQnQ0BMLoGihgiWUtHuAModae/ndPIgz
lfs4x508+K1we008rJr+wiG1/ntMf5wGnOWWYdENZEm3cc0dh9YDl8XvXH7aKvQl
ou6S7i+2AQTR7xOU7JHHD2vaDb7nASbdvvh7S1MXAeSOLSUwnLs4+2wlOWtAgSop
wn0EakBYamaFiX0kbqeW7G7cgu2BG/oZ10+iOrxgOUwOFDwxSRHzp2x5ljlokPr9
HYJZfz8RhfdBoL+wmuGsnX5IuR7epIHXJJTioZtIbeCJpwmlvFvx9oqMrM0xPphv
mAMOotZ0WBCTtVLCW4ENDfAKLqzJKg+WHH6uUuAmXt1l5iVp1Zsz81Z2F1Uzy8t5
bwreLe2DWQWove1P6DAvRaxAjz1AA6UV1hqtQGPDMt5FdRrl0R1O+xS7NthJ7k14
/IApgMmaWE+bIiTnGaE9rdssr0j7LogXYJ7II9zrPzMPtqq2eIz8mxS6nyh0blEu
Nuzodt2Ev3elLXOmvMbl1BrlD0NmK+xFVLh6seOjjo38CTwB1kT0Yj22ZnaE/4ND
vhd/epVBGPTFwhkUeVpBP2RI6mkdzT5je5FGXQ/zrcMkpRdZKECt33PL44JHXjan
0z6If7JxuHXSK8mxqeYH7G1zWglLfc+LKN/+KzBxJ3vekj7s1o6sTuKAapliBzar
Bzwqch8PtukMuG0sDSkJGWcFLfCPNuhg4BwLLyZg7LBoF9ggVApcRtUE8iTlC0cN
5KT4NTSvyB00LXXFSWtpwpU2z0zXz1Wqb13887Mkb7jF3KSLL1oiXAJP3JoWQpZT
Q3k8Ha+6plr+vUvdihvO9v3HUgJt0Q08YAWOB7R9H2sBTcJzIcCwNn7oFclTMpBL
esVvE7Vv2XGxKmpiZ5Nga+67v6feBtPvoP7+SkQSD47yXgC/Dolmx6eEFzZrwIA2
Bu23vQmkZ58oFIpCO0p3agA59eu9dLWluB2xqrr1L6UFCVYhiWnl1d8sryJM3m3A
TDK0AhKRoLnDTtZqd9Hyo1Zqi2+oqBlfZ2WineNLTjuz5K9BAzA0c5/wkyGcy7p4
hS7zDz8qIqNH+DF/m7eIaVnHex4jxHHKrwyGznoe+CzX7kzIpvdgeOFoz5u58xuZ
UUgfN7Yu4a2i5LhnaLcBdbUDNPXfvq0D6Xkt4LJ1XwiWHa1MngIGmkBqjYqgmU23
5n1nUJfJL/AIKoe+5VvoapG+uQRpMVPSNEDcqMkge1HfjACe9P+bYcrmojC1wXDI
8lbR5/xGdMaCVYLFIv1hVwP8cG3jUfJviWiwiqXwcNj+isViEnJuU2VkApH62bjv
LVbCnILRj5mxLnC8wEUjwWq+tlzE/vEBLjzqW2o44CZAm5M7sBij230AXJ51hdNi
ZxQw9zXSrEswExl4vRp61NnMcCL/T+eTnG54VZgzAbXIVVFBA7ahr2Ouk25pooZE
4IlIZgKCgLEjSC+ZesTIw6J6D0Mht+YD9g8hstL6fQl0NKdZPrBDn+K3geYq7DTb
8swT3WGgsX+TbI/cjtssAR+JvAIxeE1RPVyv63gDU/PviGaV1iYBqU53NJmHjGEp
TMfDoGuw9/DpW1VgWw2g78UH+XNqsoKe60hlyVdbmFPcJjfHkzFLy+gA4SziiEgE
SGhXoRI+R1LeJTbAzpezElA84LIDIEIMxiMn28HG+DKTsN0zArJnFo82LCx5Ptmc
9wQkl7liuIMy/mAYYNUHe1LJyNntsL+nVAveMuG/CK4a+yMayWjvX6ZU/nQ4j6+5
IPk8XPa1CzQOvx2yNnTRXFSZo+hAY1DZnVlh6MJiSSuQlZV/i0U3c+POuMA/hyrx
gufwfULwhTYflkWYNPc6/4jTkdal8oZd4TtZyKszCLgG9RA2PEpmyEiJUYnHY5V/
cRjNQEkM3grtmX8RoZIxAO46aK/rkW/wQ5qljjMmEj0lPXDRXpJbi7pJN5ZojOjP
ny+6HbQp08l2bIneOEFn2O5+mJLYh+9+byWUGD4JBzWf5a0ySnh3GPEjbK8UbyFM
PaTEzNxp+0WugsYKvam4/x01UqMOsq3vjBOhelZaASs+4qhTx2k7tKUn7lJS3R1l
otViK0zftPPrqZV370Z5bcorqqaYkj9b3QgUOtSfoCB/+mKAslKh09V1LrO7DP40
gR0xGrvRQyFqptopwgb8bKghcFmb1ldVPv7KV/JkEo6a7AcMwFRXY/Gt8lYTCctn
hKXT64/zSTHD9Abm21hcF+HJQYqC3lum/TZ1j6KzJ9MsOtOuNWi5369qkWkQwfAo
+13yEPFtnP4GxbDHSQuk4lCEu2ueetHHzsTdx1T2XuxgwyFmxH1wSKc1PeMWBI1s
CiumYyqtfN18C9Ni0xU08rAwoEi4k3evDU4lSHgLRkHX+dU/PbtN1LKRCBjXKKEU
Z83XXtn5HiQvf8IFXqewHKw8kzHOF7/dVA1fkMNXLcC8yJCh7njZ05TYV56Aw9YA
v8+c7Xx76bwAwHOKnrT4pfjndK0SQoC15/rTWDxJ/aVN51pDrY6RNGV86fYj6FtC
+LFKbXdYzmXdvPybh0IPQbLdXBv88yO3nEJBYGLtVF4Pa/z9EDN+aURzMAK9d+wV
LRyZ48cyhoTSW7MrbggQsm1oEjS0YHSE+ofDJAxxR6dbZnV7DEeFwubdOZyXUz25
iDwkuJRogR4PaKkTyMNhh13iTR6mrplwum1BO273UF/yGNmiUKQlcD+aBn/kIFGq
ymYL38DMtdLOwlKDTse3fhgbFcoxg+KXuthvQ08/Dgc+6EoKy5AiTO9GQPo7V/vm
FnoZXi+0SVKD4Xjz7M1r5VaWjiz8L6SYRfd0hJB7TQplM844MygcwI/DIUDxj4z7
vk2y/8xJ4Mhse7lHioGvbpMyZ4xVa5YhhufS+pOcGTUwXJrvtWPpZ+pvPQ7U9Vpn
AtCpUaTf86ZRJ4Hwsqx4ArmFEdHgJk77+hiAPO2cbX2MI7D+phMCwHo2i5vftgkw
KHfPa43eEe2JovJnRK4QIirDanmGX+1kDwqERifsfxg6oydwAldOqT4krEMLPH/6
TCDUaNQI3GEaSCVOcQEfCCJz0FaLxUwiVfRGxgxPgcndKM/pvU5gO74wVqGithfT
KlGoJKAB7UZx6919eFzMP6bK24PBrjWMB+e2jJEe8znSL2I8gR5qwmKl9N7fVZ0O
cWlFvgVdUS/8aneHfJ6eLRgUYL5MnDjNO6QMqMc8C/1LuHVrcyo5gJejbcZ/o48K
J4hISBeoWwsJ71Ngiej+1vjyGgdlwUWI4oaWBp6r7fKMep56HZ0zQut7GFho7C9u
J2z6tBdXvcDEUP0S5ILDSXaMQTeSvZodeJiD7cGogsEbgRIiwg0q8K9JnbjmFX/t
vsohb5fN6ktncHVu44oHicbFDuS3NewnNYr8jfh07ng9+HVGhCOVIqrKCOCTlMGi
d19mBBtVkxdxeZAj3iu1H72yQ/uaJp7nDkltzcHa+fpuGARPsDNoNxjI0aM9EKb6
zTiivk5te1TOzPnX98Aww/1wKQfGxNZ8/rmzg+IgBp9CApBrNExmp9ePvqyEXFk5
0r65nlQwuTbNqseCWSQWztzfnl+OULFTl4KNyTog3mdgKGX5KAJzfoihxqaoQq4a
foMUf8YtSNYrKblszeX/UpYjX26gAYhrjb1rTb280PBOsBTQsDWERzSa71VxqCMC
EiAqJrSsFQOvT/60smq3SteWW8UAXiQ0LdeCSGoo3yD+50wkUtvmh/uNMtLmUqx7
R5Sn9Oj2JjIzwoIXA7KMpjz7IFWt6jkk7QHzTbBdEE/ss4YGUqz7/WKYAO74Ox6g
duGcqCWW/bdxSb8bOqO4wDEtizA1FM7AzW270h7eRuGpxkSnhUeemj8YPobaFcst
kT72iixahU8H6B80hHCkjQyktF4A6jfkh7EZJvGj7cdsm6JWJODImOT5AGiPE2R2
ozrCgmdyh+eUjNubI/BpZp5Kb0PgKnjdHQlzs9DP7iAxZRNvjvAcEHQOqpQUj/60
tATs6ARG0XHnDgyIC59zkPNDiPNGSzgc47+/8O2PlNwukgZf0DSclFVI+aChX2V3
6f02Af8JgGE4nVZyhaLQrp7hxyKfsaUhrPZcndmQ7v3Pf0lFGK55xhMsNqQR3L4h
k1r6amEF6/8LnmEd80mFFlM4roeZo7fnanfATQ7CnKMo8JTPbh31Y5uLVoZu3Wn0
Uj7E7n+C0cLI9nw3Ee1KAwMSHbsRRYYtondSg/4IlABwE5iINmkx4E9Lnw0DXH/Y
BiDJyTiDc7Z/PqP1/guZi/568/TEsKAGJDb9eBubcHlyRzk0k9ablYIhMQaYhBS4
4Jk23Ez5YHaUIUx9qRQLBkFFt8XWJK8w9wOwdTIdvu8gQCXXog3V8y4lu/dD64W2
6OYNPHyz4te153kSRkbbVs+343BzwumnSCnQ9gDPVgic7jOOoVnOxVXxDtjDw9r4
Xow+zhU54GfbNHJtHZa5FB+uIMYkp8C0cB74QrEUSkDkP9gAw6yOON3s4BzfqEZB
Zi5Cp7Ulj6sjG4UeZhNgpD+kGG+myAeFYXgpeVce8RsZWgycGV9LPXk3PnKaYLmM
wTF0Hc32OiBGOfazlEV/T5//PxGlMSCXP0WgFR1eR2Od8xKZLVVuqAxlNaBQKvYz
Zh6CBE7PTlzlIcyONNJDZUBLk2DndGSupbV7rvB6Pb405Z8PS2QMFYYYSGOyGJdR
oaBLVIcAPd1bofg5uBLcfHxQhw12h+sQwWhuPd4ZKL47QqV7G+EfotqxkeusR6MF
G+FKiG1QOJsmZ+OH4V2ularBKsqD/HMWCRpJ82QsnqPrLtn0YvY8HlFfggsk7FFE
3LpOB+rCgDJMLFGv65ApXNwMESOCt93YlqrteQmaTFtbRXPWelWJLohY8S1T1TPW
9iPxoRkeLtEUHjlTIqFimFXMOIYtJvLKYSzrJN4r+yQZKEcbQqmxAOPGq9jCvmEs
AKu7Rpz80TSr3Bma1mGWBBq0KQoGMWSQ8gztqMM+sd/MqwOLkAG+f1ON4dy+hgRp
V1HBBFpHdoM//PofN2FePuGMpUuSdvE5BccBS3oWvv0JZKg2frRADmSC94Iw+ia7
Xopy3cO5NUUcnxzLFVmgPI6PvshEep1vx8A9fYfMyfwDWPP3sYJ0Y14dMrCgzTvc
sjyra/bEv/wGyeZSmrBKGSgYzYeKTMshPkZb+/HkhrYJdyKjgBW7E1DsekREtecP
ELzHx4arqzd1dlane5EdZCv1OR8pXsJSZ1dYCehlBdHyYLw0LoqIWD+dVUh9/lmc
ZN6koY7YFJUMUpCOJKf0u0dY8DtfI2BqNvOU+H12Tha00zdug7vrvF2LBPBVpCTf
6v6lyRwC6XTDp1qV9nBeDY33Xo3r2fPtMuCmruBSliSukJF1feOaBOV7lh7t8RfV
6WFGrlIXzuSXx5XRAODKB4nIjSF0XUbiD4bo4RZmR++bk7kSdA6nhO6zvPNzvibG
+3N9aYsywZdIIzNvrPY8KWtnhTKhpTdfHsGcTazzU2Dy3XxJOZRINZ9LO2D/uxwP
uem5vPnph6+/tIfOFmAl3tQ/wqiALceeZ4CtrY3LHSUPDrY2j4A8QauHX0wBZaJO
VU82iMJ1nMk4w3/n0ZB4Ml+4lTnLeD7k7nezj3KxgUf+zUHxa9ASJ8aiquuFvYbj
N6bOnzeqTXqD3ZUQmj4PJBHsTD5vPGC6O3r10FeSCWwtPY8z+iYEVLmn4OJ028vz
C5zQoKmF5Ww9HY8utRRITMVoqFdM9OjW2xpOvJo25jqjaiJYlq29/9+uaLSaIIxM
EcWIp/h3Q5AX1kquY7qgh1dFvXefz7Me2+1zPDpY/uCnr7i583JbnCXeI2N63NBI
XbCqTRn5gFPKzTEJ0egLiYez9tCGu41Sh5bwRiXvT2gbMasrJxSg2tGxGViz5bHf
iqtUHdrvihYfvrlwKGeDR29/r8Rzap+B2ogI5rYBZtuj8ncmbOtr07HGQ9VFxgrA
gmFNoDgyONNHmIEtK5JFn8Zkrle1ZykrDhOtDqndftjIaTG7CdSIMFqvjmwtkYpw
fiuZLvhCJUsH7YBo2/kFlOea6sqpblFQJg2+jCi4WmhvaYkPcxqOEFp2Fq2bgVU8
W4+J+f6UViEgIkTtB3c2qZvjXT+/reFsHOdcDUuH8A1LMBfKqqR4aKN2IWRl2p76
EP72SJghr8D4YtNDDN5f7mEH/zOCYl9qja0oXaElYNheuvaK8UN+Y0RKI96L8FE9
YQK5d1LW44QhtTKizVVsmCrxao+5N6vpCct78SW+7KhV3abObpVnZ4wrulqx36/O
dZPYS7RgZbLQYm7YzjOt+13MuwjuOFmJplCO5QUpnRWAvpw5vUUNwT1uYckpjvnv
c2gagz6zxrNZFjEt4VPunoH7NSjHGohhU/sOIxf29kOIncypjb4yhgTveRtBOndf
z2Uj4Dops2sh/coQUcqRx3gckSq/lxK0EE0YRNWeM7mcH1lJqy0FF2q3omgUrFfL
Woq9SB3Y3jA53iqHdgGqCcrft61qcA5Or5gw/L+gQTMeYxO6WC9Pkaq8+4actOf6
quMwUYwAdBIX1827LhHaxIyc745+0ptp12ZgOIkT0zt2iasz7gmzCjywdgnqLfLZ
sTPBMbpoV8VlulXZ/zvH09z1i+gi3vTKlle4gPlzyhnQr9LeZrAteEKaKtlkjus7
OIDggQi2PMh9JQywkAoyIUGMIeYyV1uCIl/9KpjJEomQrk8uCYDN4T4xwd2Lf+YO
2XTlmd53fDAo75PKl9rUbQEzcXwgvKHCKp4jaGPpz0NHV1WKenit2yXa/0Skr4hB
+tvyqUaH9TzZfzuVPz6nFO+bG9rc3WcgheDWsH4dFgKGWfIHYSWzN21B4rU7jVZa
OpzfpqRWi1Y3VYCSAGesy+0mfL8vxEhD4ITbEwX972Vkbusdr/jfcuPBzlHGeVeg
y/uLouFGFQNvbIZqgkTbsM3hmBShwiPkYDTcAr7bpS1gzrxPs3TyMgNbB4zg9v9t
UqhcXRYygZe+KlQq0KlB29FlT4SopQp4DmxflOhGETKv2gxh/655URGODu9b9vYv
ciTq3HVbgNPyC8Qbev8uq0pQ+ELqCIlhWGpa924vs+87an3xiua7YjK724WzPg9H
ChGnroUq7V1k51Cm2n2DJdlfP5GR9gCo+SW7JkbpKzTpJws47BQYlt7dCP5CSnfP
ij184HO22zvpF7m5fh2I5Cq4wycnSxgan2ixqCH7uoil6DCHSjXjzhtKJyRQd3p0
nqeKvwbGFkai2UTlAbE2gce7E9lR/Zm4NGFDyzp/oBgvfomHb9jnX63VdXOtFa0g
hgUWy5GtRuSHklPondoV6gR3DUsblM3pBpw2Ur52QYtcNSwd0ez3SQoG0rft11d+
0CYJ1teuhOdOveKiLsu7nsfDVCJ9qdYMLi68Zc6yuM3FQRn71f0UW52e1It18XMe
DCfCIx4zzc5Zpa7brWBiGqs6p7doODgQCAAZNKGAITZ55PxtwwGINnT4ZSXJ0dO7
cRvPLb7uqEJDH+OXXSndy1Oza96OyS3tEa/IvBmwVUR9E389nA8U1xjUgBAEkf8s
HGbybmWbptKydFgNmP0i+En2fSWPhotFSuYQtrZOWiNLZxcxaXbX2CMMXM0UQZTK
MENJ3V7+8ErXezB9r7kdX86yLst/EiTqHoAypp3qZ9xjBF5+7ylDnP2BQBYX5XKv
EYmmrTjzafsbR/LiF8x2VlRBL2AdGy3NmOJK7cjqATTNGPTjh7qpihdLHHG9J5cA
AHeRlSubyRqncDe8vqYJEMy3F/xMCZmcXikAqjnwOoSKZ4WEQhhPZ/bxF+xiwBV5
L5QN+UUbXJKv5r7IcrcyQifM9oIh2cm2E4VSQ5LH3rNsVf0inNWE4c9ZAOV3F9QE
9vGIUkAbMf2DEq+Zatz4NgoMY3IXxAEfaYN7cTSky/lNsFaftSbhJN6+uKR/XEje
TVj1L9ONkb7ydAbYqpf1HJLQsbR3q+Gu4rdDs2WCYgnoDgNpYy6Q4K7jFDyUhnSa
r3ovpDyCtfIOI8j8ctkPvEedDj1nfmyKib1ioJT2a7qZmGj9fMh719BZka1EecGg
tPDJcBntxjZ5UqAI30FaOPZt0+KBUH6MyIkgGXGSsuWEoJ0alp+XbMqb4pp0UsJE
ThIcYcc8AHCkHid+QQ5JB+El336SSG/K7xy5gXzSgU6GqCg4pfPdY4LMuZ2V3Iv2
rxx2ZFdN88fhP9AvpXgQHnGxoKgvDSvuZcVbXmSOp8NfL6AQSzYu0DHrjqZAx+vl
sPlbhgdquHYOlGBD9wsjB0ePhtxRCZ943CRd4ezfcGDY05KKtTXVFypSxYiWOYK8
jRZ7Fru8UV7NeI9GHARPRlza5Je0EilrPkFMaNgpsDBFhWZzjM9fm8uXtq2gjEEa
a8psg6mz7jHMzaZBT6Tg4dORbNJziV5JZHskRr+Vgx5AwOWx45/uNmJ3qOaypwtx
4Rxn0yG+xCxEx1d8kuN0Y+J38HTg9JuVCtoRvLPv/YYMWnr9aQkwDN8Oc9vcikHc
VA5rikYnk3wCFxl70peO2mbEb7+MttHfyjN1m8DAL2vOeYzxewkP7EaXdXT4jidZ
RQdWZnsSW/MD4Awz45+45GhzlHksLrg6+CugqSyEf1whrKpbXsJ6ijWBqeL1q1vj
sSJ9b1B2xT57Tv7AypuiJcnSGYJxyn7yfReehqm3/tsrWeZcrfJy7oL9RO62GNvU
o86kXBhWTCGdsSbgReBWh8qvQZDWXA+syZ7HsPpF7F6ILYJOoQGMEwN2iGeCNEkq
TepIVmr4e6jV4cehm+QRkMtiK+9rxpBkBmruMVuRbELX82xg7GbWZ8C5HN81kPYx
nWSkXCK9IOggE4mjXE2HS5xYAOraTId9ouFnm3DoIWvIoyEkp1nGGdBq+u8A0sql
NmJfLpJTBAiE3xOb99+/4Dw9mhwqAfeNITZG9xA0Yz3hwgQkWGAjZqPlkfw5Cpf0
jhGF8XCOLABdZvp4+77BenYb7r6lrAcAhPbx0gOshlbbJZk2B8S96GngWURffDQK
o/rIokc7BUqKZXSRsOaQjbEXVdI9oEFLCsj9B3j49IOBFKDlbZ3m3Gf9RxdxB6PZ
k0f+uQ2iLlSOZd2G9TmYSmACnSGZGEXDteXDIxVZgtudhAkM9LXkldKG8dWV7z/P
WAOjFmm7kc+NMuHFAGzLl/8YsibS77ZS16U8CSWL7fNyLzJP22ctzq1OFvNZmwfK
mlt6hqtvaozaVAhyMRT6KmqQYJ0ux1ADrWVjPt6gCg0+zd9+KBrro3rHDzV0iB7j
XV9uDsJ7vFSXaWvEdCGs9LG33yCEio/TJW9wZ3Kj1DhzT8ot77KEN/HRk03V6reI
20Cnai73WV8+cwfKi6XEehQOm3DabTXMHaYaAlFFrfU6dDkeENtJPvFFoEO/m+dg
LGm6HsBtCKWXi5hQVW2dSMn/L4ec3XIY4cUMjsNMWM5BZwbm+8ktxIoo6TTG4m5D
3fBqKcNob8fntdkOQogPpWxznCXXnA9wB/oYqoQ/b1i6oDq95rB4fUrUVt9E6FpH
Rxu9jB9qjVAuFSdQOQl+2sFEU3IvzGbcEwxYXlp/fMmXVH+JqcuQDDUEZK2apaPT
zF52VNJM1LkUfKEjhjyP+eqBk2VN/NEE+fgtO1g/OqQXcXDZ/Ln8FUvkfTuUqnYP
xdZmgenGMfcF/kCKWhf/5ygVoQESPiIqpPAwqjWJ5s3P3eMhcCY4j+s1lnVAHasJ
yuTQ9G05QMvjzgj5oXTVn4MbkENMbmAQr+b8/VkAUa6qPuhMshJ3hxJ5kvqsduMc
v66uZsYhrb4shqRORWYFJPysmYkttNnQeRXByXkBmpcTUK+1ewEOQCryaSlmTlOi
wQ2vsfRlvu26dKXAWjT9DT9yssZ6HKHg+y4n1c9CmWboY5WKE0jJ0QCol5qr4Egh
uS2T60Za34OYJsACRmMW6MqlekOqWXrB/WVqvGEEN5dYZE5+uqbcORH0o4RnIsrH
wrrEm5mnN5zwRPagkY7vB6ioHHLz8xDrLrF5LwzsOK7LQZFQVsf/FhQAuyF04uwt
Bur2/LY+g+6k8oMX0xdV1pisKHNwhONKsYdo9Wu4ZslG0RVhwhB8Nw0ZR70ZKGXa
jVQ1lRHn63dqWSIGr1+BWe92My4HbhLgNyy3Jnl6uYQFNMEH2N7JwdygQvou7LFr
oqBAaWDBUM7rE5rZzbdW+lQ7Cw8Iilktp1SOwHMG7wTU+DHrjkrd9H2ClS5WVPxW
zt+75kvYEyN/070M/GI5cR2TKfGbfXPkMB5m55nst20X2MDGj5SpRAnx+tcIQzM7
F7e1EyVOXDtuTLMCMTxm6rYOxQz1iZq3ZM3K11JzBKFHA2kwJjo49xOMU6JuPUTr
kNlZQDMtX2tIDAG6QoNV6V/mFQv3mi1h0r4b8sCxTl05LJCm9l37dRd58U3PPFpb
A8hC118N22JjD+o4OTWmiz+kEMdt1nLroORYOeLKErbupi8C3Ke0LTtMQrFucCgX
tLdwIqRsPkJTbX7xBVUl+O/N0ug/DaV09tp+6J295rr4nUMnZwlD3URDFmw2Muzw
g22X/055R1OEcxxtDlZt2zu7yoeJ8uPgGyjH6iz5AllSxNcJss/bovVgtk0OmjtC
4z9d6NfiLE7Rndg+5mHE5mGoQ52puD65+RBxuhsSNGeCk1LuulRDd5V/iLWI2J8S
MrxV9Vd+cQkr5hLZc1Rek81pyRPmrCS2zloBijvFB0qgnbSWLsy52aXHU/nleP5f
4xiO4e/K85JtU89QaKxHIBrh2sPfHQaSV+2Dg0Tnsb5HN8HZqsZUirhvOZk8esW/
ks2Zlg5BCb9VsU6z4lD279dH9IhX1v7Yl7n+GbKHzv0iO4zXGfjIFYfyr17izuBW
YuIg3T2ybLFZHPBZBac/UP1fuxaabPpQ4KtlDbkhDUjYOBzTXjoU8j3P16Wjdst2
ZAQpfniHQ4xlhcWVvQpXsueZKY7uMgo2GfHczQC0mpqSUYMyvTczGr9OG5EMBR/b
NR2PvrY88gAn8LWR0Zq1eqjX1mso876CSsUn6Omvt81hrwIohdHC2L5vz2W8QeUG
6cqSZ3Zndu7FhKpsx4Yk19wqh5vxrBf6Z7rFSy8ZZAZJ5iwQDUEGW5kSmrd3KJK7
urep9udTb6aEBrKFoQWsijlgGMDXFcnhlKXOqMqC8DeJ68sP1/G3VM+lOAFerUfS
TUMNbR2A7sxHoV1Ridyt9sXWFTqQIcCZqY3YeEpJJm0I27V338ommFrl8ibMw3i1
H/6kknyIlMWLdhq+C7Pm96i+ItMg1tuo8dNHzrSWLTz59HrfZhNI3dmFsYOAUe8f
iBqI075459c6tYAOv3nyYzioO1d3yFGYIKBNs0/Vv5sy8DRWUWGjp27lUZ+txRlp
rdmJp4k72S8Fn5l3NmB+8t3znWToO5wXqYgLOV6qwQnPgVptlgmDmQ5CsATUxIbZ
nbi1Bx52fLjxKBO9phbHwWofYpcThuDRVZoHSbjfJ3Imv7fdTlppu9h/SO1Z/txj
OW2tP/wJs5AoNVo3VKp0d05UksYsoBSOExR5fr2QrFDI8VK116KzumKgcjAS8/S8
f+xNySHL/XlySeKTmvq426eW3deULgF1urIBOAWZWYlG8RI7CIzcVT7zPPlahYdu
8X9BAzvvGJB1TKuGYVfibamg9rFh7iO+m5RDV6ovdDQSACsSmmV5ItMv7hGb3CxK
r+2s+n3fVfNBm9mrcxY7b/K8H0QgY8z+wlYamDDdt5axlCSwVOQEdVHakWaJTdGS
9MEz5FAh5PhrNq9yrapqSAs7rEl5dt5U+IjmVa0XjbW4e0rg3/GnvBM8rcw7zmcW
DxgakB945fgcn0erHSf0U01ja24UHapXL64YPXXM3bpEvil0ZpyJ+rHGBEY/EuUq
tdUUF74BVJrm6Tv5JSISUedJ8/tHjsOAx1Gw9E8xpRqg3mxKl594oZheQ0qa/lom
iPXTfiSeb2amC/G62eJDa0RlqtpfakYTIcUg/sBs3olGdr4gpahwdDBTpOJjJG+a
FntU15WAfrsO48WzEmK4AVGuglKHNxJtTjYp9/ZOz9mI/+KG4SO5hpEidxVKg/4I
ULWmLyXpI1xnwsWCiuaB+r7nkhDvwajOLiWZQf5SpjmphAjU+P38RP95dADb9kWq
BWumm+L932VrpYsXNwLrkjYbG5yyQu7Vqp4KDEVmRmDyjqk247/LO0JudLh4WeuJ
fW69MlBf9xS6CmIsbI++Nd2gdYQjM5Sg4feYWZjuN+ZKaeozNy70+RXlQyTi0XPS
qkGarNyzuB4KDuKSqgNM3Fll6MXgPVgqdOtMB4Ydc/xzkhTQPpaKOgNUNvd9tFVF
KTrlFxhX2wnmyeRps9HWhPe8FG53W6+kR0HuvrB4A0JXtXCrK2WqrHDxBp1P13vU
M/unLOCzqFHNhuUx8BXcewVImI8XUoHX4xfDaHIp6X8ErpR94Lnnc9vWgp3MZfUR
DrvWoz4n8eGzj0lloayzac6SxMsFjAdXnfTG7yGwusKvXDJaJBJvPOtq1/5Jj4HX
F5zlYIu/z/ffs52ipc+9kUXW500Z1HyN0nLzkgNVKavWXXgy7t4AZ4wZIoKnYfus
J1thFA1S0B+2bixxg11wx1Pkjd3ysNSoC9rzsAlC8hMb9oAh3CoR2zekIVwBbOxH
CExu6ENskCEV+ysJQHdBiGMZtZxbH3m1T0wO7CsQj0ag7le8MWM5JqUAfaTqXQXd
SzhA02dO203wyJmArNVF6cEPU+hnhUfdBo0TOxyvPHukf59Fz6va7vjvdJJ2Yzsb
pjNVm8ijIK6Uv1jFzXXS1ZkxyLgi58dNYfdsPk+fapV7aQsELamIHZGh+c4DXHS+
woA8WbPZmihwyzraiM2TTTxxyGX+McrQEQYON/tCdymhLh9Nxi3GMjjuviCkuQp/
J4/Q7ctqd5x+e+owV37Kszmw8+TUe5tg1Z3JhnZ+ZObUAEg+wLFkRhjNuULBjjFf
fWvcnes8l3FJZ/apdx594aHHZLp/Oi4/FyufX2i032OH3BQnjVENwmt/YDspqe/E
CLRdVPRs12ehPf03/MpQE/IXtrVHTipztHPQQLAfC81nxN6wPEUp0SPTn2RHxMun
Jhib9qQSZX8rRxlafFRPnDHiPsF5wKGjKYRnLITLyCtb8wgNROtfuk33fnwP3KJH
xSKdOPxqBlYwvBYyP9OABvWgTHLwwTJEtHPDG2pNrqk2Yv0JjUqYOhqFBTNOh6Bo
m5yPTtxV8q/VI7ie7mzanwpo/1kSCZTMfV+OMZUbvI2XCv0DS08GmOIQB5ToDKy2
HgOMh3ecEiXPPSUVAWTnO3OS9zO//fVter4lIkwld8mLBigZy8xe78RiooE6MReR
/kHRneNZCNnp8L7MSt/HFUbbmtsg3iwyAVvQEw9tsBdByOOWxTNTcju6VEIzDL9Z
yzzyk+EguUCNuHHZrzVI1ZaXRmtG8Pb9+zcE/rEP1zkugRTur/lfMyvnHv35bnRb
2nacnMD6/Z8RHBrhFXMXgnsIDBHS1zGjfdG7QNpaN5eENtUVzhJ1IL+yKKKtrCD1
hFnhED86B5SXCZ2iSGWJ5dUcVmQ+eTufZv1+nvUJzPGaKSCmAWTFNkAfqNey8CCz
frGv5ShFLRq6+6SiLwFLWNoqC1ep7ONqU7hYOhhYdJVUUyZrOTxYx9tNa3mU9llo
8kotj2+CIf+XqWojmDwgYnaKuPAYR6k+M2iXHgdf2BGSGTcvuQspm4WAueT1eTqD
xn42OsOxbhZLVKm7N4OecOv3ZwV816q1RDL6+ibwwJnx0HrKPJxJ4oxztNFZr1+s
mzRyD5TFPzHBN0OkzYBajNvWQFPY6PC14I2rUzKOaU0KaL+iFKZ9V9zvGZ26Fvyf
fZHlyf7xBpyt+9JPl1YvwxwqTcBZMVd2P5ZJWE+9IW3X5shO4Iq6fLWRb06ynOZW
UoA3za9/qG1kifIs37hdntTjhCwXGaOY4Ib0uiX3cXUUdb/FvA5wrR4Mia1ovicO
Bc42kdASMQ39dgcNk3NFtvaeIH0ZyhGPvljEeofgx4QOQp10WWhtjlr2Qq11PXpM
ZlcLm/JuPDlGwueZt+bmBKrwcjAwXkLgP8B+papqFV94prI+t4HXqeM5GLnJ+K53
Drhk4yJJlztdzGwvNwDDKIBQWsbiknbSyqlBGZHCuCLJMo1AEzj/cCYdDNzVL8i8
HiGd2b3pgN/jumm9uJob1t7UJBPL1F/rkqkT/lCNZVUE008bq/7hIS3YV87gJdKz
IdVZfLVy0En/JNcZDBuG1jk+Kyv5PfppqYn9mRgWbjzJikHs2DtaNuycbqkaP0oR
Qb9wNkMPgHqLKRvuvZvE6eznauJzkLBOSJyu1zyMB63Jr4VFfkm1Lgmz3YfwbmXg
xetTbB2pNcbPzB2L+ArfI9O3msLORflTMyEbTD4dD8M8XayB6dxznX/h+Z78DuyC
fYxErAAhBAXxfXAO4YvNuQdi66ApZUdi6agAc4nEbMxgVWiZRPV819/8eKZWt9UI
n8SaJb7j5rQ8ck/Bvf30BViNZSaMTsC7I6b/cPxpwICOZErXtxj4BaStTCa0ONCV
hsqz13zMU+aoLOQIFRV17nNC8XpRkS5XpqyjSGcokZyk6EjJVFEUyne95m+1w7nA
RVVoiZkQHXkNnJKYCryXj1BogEq6ZxnlLUYaUGY39Joonq3/M/puATWRBR8FkSFr
fjZjhruLAmXjSyjkVv3B5bOt4ztqHarFtW7F/IkLss778/ycsfdx4dJmiY/2lWoB
7agFpvNaKOM56LiLsClF1tYy7nkyRyNG9jiAWgayZiZ/gOCUXhEC/7NSKsvji5bD
u7BZzhUJAAqAJ5zjj2nb3pjrRTVrLP4rwSH72vQ8SvdoADMGzimzH9mItDlYKucr
9lcoydIUc6THqCFLMYe+z2/jOqlPr9fo6DORHrRgEBJaO0XdYSI6Dg9yZIHtoBPS
GIwyF5gIhf7TpqGEiGXuIvHF9GbKutRdD8qhCX8n89ZT02YH0ad3NZb/6HUdEWo7
OO1j5Gpf9KTiqrFmiDNf+q7CbYFVcaegB8y22UEqGL+bRl4QZKrz2qZrtZm/6nJV
9AyIll31MWmEFDul+N9dvUrY0y/G0MFaESazT5SjnAKwoxMciCAHEvN9B3mDHmtk
Zxl27ksp9y1Fob4zaCoNOo7M9yUAnrXFCQMAq4J1YTJILIJKyfbDj/2JxcSI9ytQ
s+v8SmEYaNnROOd4iasCLqDU9iQKRxlCNydN6BH2M+PdPKNfgGsI+UHFydTsg4Ye
pPtllRxskYhE8lKWkrQpqOYyWD9QP9KE5nsEENCLH7EdPbpFoJxx8kaemNqQsV10
Zw3z7F2SKWlAtn7uurbAneQeY4CD2aqPakUqWJ/YH06yfgZn7w4GCzxiu3As46br
nNy1I/QOBMr955vegO9Z9rMORLE8UxoMrH/8x0XQuU5s3wVZg5ydLz2ezHrogK+G
73OQEfnLicMG5rn5FnkqT3LBh72dnTsp27DXqFcCx4R0ict1BdBo8ch4AkCNZXcr
xgMgs3qvvF7dSiw0ufTp2ZkG/wkT6bdrgR5erDkhuD2e/uoKjux+ehU+JE99zofa
iFe/GltLpZps/FCT+WxWPgb+WA5r6Hedkfy7tsjKyxGNb4HB5q/m2NPS6xiwjhby
qzxBAmF7UfwrtUHnlaxU0rrQ7GUBKwCvYrWvDRxIMZOckqiC+Y+ENup1bOi9Bd/4
2AVJPwophnFogmL6ig6GsMBHRILpu6G2Rv1feD9ldIz4bQaO+RnrKhVLYxpEzVwn
XD7uaLvjToiZwCVezH0JBcxB2DWlUoUwZFRBHVLabVQ0AbmO5PxfCjZle7/arygK
1QW4F/h62Q0HtnpQxsN2BvGIMVW9JIxnlOOo5LvA5i/TfYTZY0Xw2C0jjpO4uWlM
hkns0Iou37KLbbZR34hk4F95fxEC7kvqAEjrqm+NBAJZox1wPblNS3+3j0KwaLlf
QaOYVadmt99nar4wZFgDjQ5Wnquy6A/p9gj5flzyWEC45igenA0e1XrETGgeruns
omOOQuYQWoj9BRpGMHx5JmY3B3IQfdrt/xmSzIklqWx7kTB0W5nmignsg1/mT47j
h21taEWTynb9E8Q1Oyn64TEr7ej3XBq2cCCTSx35B+zMu++OibDS8fJe5ON3/HY8
cKJObfVUnXmTdyKBJWMhLK2h28RKcBfvKWcT/Ai2Q32aJp/28wEQ7Xev3taAI4rY
g0qx8EzCkpK9HZn5IwhNT6/+t1iRPqR7ei3lLK7JRMkb/Si6o0q5b/SfVebg1Ntq
zt6Ve26piJnILZogT8hR7KU0WCFEbk3QLJHWfwfkoTL5YE/E0yIGNvuyYWKa5061
f7myX5Gz4c0uemc3Tit9xmP4IUnXiiZlKOfaKhvJq1dTGdKiN/+L5M8t13USdpwD
K7iWo/alZxDilvqQ5X5ubIoEvNPscDtabJUHqVDTQoRJ2Y6lw37mhUsJUTnlK0cb
O2DGFSOHTcmEbczpQR6o9ei9w8qnBSG/mfxOwvXiWPfclkB0P/C5yi+FlppV1LyM
MfdrHUzk6yPQLN3kTSbQWMcUBC/q2cEgY7G/ac7I+UwUk6fnZ8ILqI4vj/8AtReN
awquZDlABDk9B/Ko4y4CzBXoTH97W45DI1g55bG9EK8mkKgDi0dGA6d2Lh4n19g6
Vleu8mhOb36Bq77bhBfzU1DfECqoSx2K5cAUlHnHXeqQudmRSHUPOv/gniVlQjkM
oJQXENK0S+OLHWF+vrf+w6biGhYUpFKsQTeYEgGNy9C4h4fIkCGaoskonpK9CWLW
zFJVU/7iwOn0xkfCbP5rufPKx0OxTwYdXB+93OkKn3kOzSVY3bV9pM0MROZp9hWw
iMXihKH/QvmvcFroAlD2yyRQxJDWuBndeXcZrySYxx3ZhxjEFuQI9tQ1NXwaXfGK
5l+Wy1UlCF3scArYc4JD0cjb/pQO2iCMbcfQUi3Q2xSrLsjLdByXyzK+7v9RiFOW
5OwZ0ni/VPGzdaoiWWJj90H9lmlsdF2ycmrFZiW9MVtuSRQDBoAjjRdWVg3BL/hg
Lzdye0nG4OLzuZ4HaC3krE+5q03GcIbf3QNWlMQBhboJjoDVxRaygoZ+ewtG/TeV
EIgg+RH5L5Dyj7rAnzhCbKCkbNBOd2vI00WD157JOpTHOXMWo8K7FiINAB2sJMMl
yCcMPcRhk64MasAuOANYq9lzrvcnX2PVjNVEfvn7BdwcGDAXiY8EeIH/7a26/R82
+apiA4Qrv7v5YrsnnCcakMANxy8lFn7EV4IpASQYD9DUA2Ki3jZLF7C0ZBVmIJFJ
T0QoxIJuFAeW2GETQaU5U5ITcMyuXHPqW41ALEOEmb3l4alBOUXd9ach+yVGlHEx
ZiWfEwYnp470Bi31F/dSQWzIdb2jFuggtsEn2yIjzqXaAyaG/PvzAn9Xn/vIjGoF
qcwyJd0YpFirTb3rRu9zJuyI+nK6MMuLJYw4K5s56rgT7MgrmTiQQORkgz0Y9NCs
WYxU8ZB8fWJeBiIHVf+2Eb6nrCXxjebXr39pIPDg9+xkHEnH4QSceLRhbEr435pV
TZXWxgdsSKU+OIli8n0KuhR3evT1ha6tCvqBZp5gKEF9hksRofO0igb1tCwHV0BQ
jklBhyulTo0De2OkXlb/ghcSTrhLyMF5YHLHczScj2w5qnhmU+799wBA4MK8OT/F
UxPju5wxYqCVYaam3h+CH9RkbJysdfuT04kE2AadUvcqIRaUBVP1BbYfBRo9o2xC
1CoIfqyLsImWmDQalg/Lftg7+KznbAljiiGzxk48fHlYrmMvOxPk0mm5OAqlZvBn
g+Vpvp7NsjFYRz/YYOlEU1OCpPZoQyMLSaFd6gHMVjs82Gt50RBrQjJ7CdvLGCgn
P7Xpuu9mgOykFHSxG0omi/R3GaQy7qlYVK7R2PwyeQhjr+1CINcRl/JyqBZ37ZqO
FPQjrIEIrEWcsxhSxhewCOsBA7wDvpcpKlVbhcYfjoQ38nK41RCSi6gWkiukoXpa
vfHs6ZRCDrUqVXuFrhg2DAC+HzIF13Wy91NQ7MTY/OiycF1tjKStgrgIVr7rTcqD
5RIMZKfnuoo93JggA8hw4LWXJPplXeuLilCw5wILZaagfGPpA8mMfTQTIU0ucBHd
sqCyeE8ERc6P9zqcQ9i+TBMguKtSde+P63tYUUF4X86svNopW8X2K9dF/hSHukem
Psbdy5Esmwlm4h+0Db/F4nwZg//jxdZGg2VEG1OtL5wTiZ4StuSUwHgzeepDJX1h
IHk1L/S7Ii0oZh0U29NaRJnmXLzBpXQGthseO69Ms7bi6GvdI2iqfeCKqZCS54rS
zfwg0gB9M28aMISUHpZC+Vq4xx7S8b7Vj4L8hgseHJpoDGZmcjYbbi8NAGiiWtoH
2M9jP0ap32RiNE0BxZaDS/UjPzfxcp52Gs8o23fl/mtVHJxA3lJAF9HZi4/2IJqw
YUkGX3yWAN3wVncSPblzwQl9GgEl9gkvCgG798ywWivjulsTY9DQLms1qHERz1ND
acuKDTQwL5Hx8eGS7xECUEk32+VY3llbaW0mqiFn+j1YJZnxqUWjtMD9fokTHRVH
8HzjqZiSoIzXbcj/sBM4vG7CM7CObSNzunnb5gnvbunNfaFpvW2UlbiWPjyUIELd
69QsRPCQZbDiLO4B14T0wtwsZxtUm6GqdwdXoEO15muukgXbK3roboVRhA2YcUu0
3bFUsTs9l0zelBgj4WUIBm/0CJXwIOeCwuDtx9cfyYcI3bIJ4/ZpCsr+CZqy5WFR
pPXaP2Y1LPhVKzBHKHg0KFMrOtdqH27aAiL/MAybmg8vj0bpixw8UfNFlYtcS7Fy
KAAo+J8fOFD7ypIGDPjYh8smizEgKW7DjueTr1JrAknEItLMT8D1TfapU6bEsK4c
EI16eWERH750ZijPUiIdXP1q5dGdNEfDPxX2LShwIeyzt4CDlWzmS//0g+yUs1ES
Qmy9OwcryKkU65ypmhHgJjdFwfPRQaOu9aklrjCUVLP0haNz7ChMK7Ce0WgVcqeD
5Z61zsLuo4k08UZ6h3N9bmrP8kDFdXLz+lJLd8CXczm2dY03AMumhi+uKK6xv2yY
R438Ejy5cdXSLch7BGTODHlcoqT18kODw+tz062adFMpzV5YPsLl3uprRLJ/pDWE
qSSRmJEhn9dzhW3g0dtixSi2KhbnsQ76IxKnRxhvkrHqS9TbYpkcIkv1IZjN2EIn
ZExZa95iu782xjHZ/TYjCen9TlLJZ/porrWz1BQkcbmVFXsbwaTirALFs3lDX0Dh
2FrLOMUzfw1ef0XplBMcMcakz4RKRmN/+48BCJXHbpObONwV7suJtaZXdRBPYuya
bEJYTVT/Ho8VKC/yD8/Hi8GBe4m+SaDzBPo9e1PkxBUtxzOteD+0TSrv3uPAGRQE
tDFdVnwNpeblyGrpLyQcxkc5RA+vS/MD/DvS/8067pMq3Oj+pNHEqM70ie8dmtZ6
jpmlUsH3ydm2QDyuYzasYQrFkr0inCXL//uaexeqy7xQyfd05NOLe7DDpJwaXkyG
28cPTJ0H9KjRVMndJOjBbc2pkl1c3RdgYoVTBvuxcQ0A3JeKOgrnGBzS0kdhWBlB
sy9VV1/qM/KYVWWsupPzsJeT9BtjNab2ZS8hTqLXFGqxRsmOphe0VDEiMtZI0Ibu
lbXTyd8HN4C6lqrgoRLjKR7+KHGQKrrxv4z0gk8yY35dXaCBZtsOfCnZNUOVdJ3b
KRvkbyHX/hjxCu9pM6NcBbS4BInjPTJa6eDN20NJfNMjS0bCZOFxTwljDJ0XzXvs
hS6x6wP+AKLrZVyLEdOirImz4Dfaqx4au/rHWCHkNL+E02FlqDisgyCkOJjd+cmX
3Eb2aLOk+eIrGUVdddCckEKwRjmrebA/lWp3MnxzJKAgcvXDLy2l2QKvjZSQ0DkZ
C+0nJGC2bWn0S4C+MhSlifMfkurABO+9adRP709Rw3pEw2kutqI1DvmTxvJxtseL
Ezz5GHaEAXCAJGDewHO2aaKcYQKN4if//o8FDSlLEMCKsE95YOnl2WpPdAOSy0gk
bngdg57IDJrGTPeEtUGg5E5Us5sc9NbTMWIhp6XNXg8BSlOaNm6EKBidKegEs/yG
u3B5w5AlsIZLBGzXBvruBV21PQslcZqSEG5n/aIWLLK7E9By8NgTz9ujl+7LUyTl
Oyo5H3XXk/D/01537X4IpLaCOInPP4w7HzXocBe9MXqdyHIy4cMBlW5X6L/l4Miy
jlpiQ2QFknD9pZv27ghpy+qA7g00DE2GQ3ANmCdO0ZOq2N6hCT0hicdWAon95myZ
VleUUhYRTqxTTiatsPA0Rvbayp/lSN2pG+1xi6YjSpoGFHNWqEGbgDC5WDDfWEth
DocLxvZIWjz0itvMeiqHNOhr2GxvI19SUzgHCwkR9qn8igMywb85gjWt28XNJDzN
Y03WX9UyL50Nctv+y7tkNDcW2k7f4ks77hUv9YG64pIMgvzsohLtB6vbcih0Nzb9
5V/s6KutsB7eG0eoFCLVL6r2L8rNY3563/YrJ4+BuB/pr975fVBTiqMr19Kq27Ti
NRPiTS0g8SN/RXiF8c3HgRNDQDdsJY3Z0BZ/FQ+0Q1oRVDRjfEHqVL6kg28eLWye
jlx/9eeROKMy5UtI5OwXgGq0bhrbRDzxCQBFdQff+y82GZBbtJiaHBcpWAr2LeHB
VuLFdn7DucyGKugKDqGRvLeVlBLHWdqQWN9L5FQh9o9OA7AYJKvXsiauONfZsCEK
OF3VD2EGygqKIMhRBE11D7fyVtOvTHdTYe1WMkvIa2SbBxaD4L5oj8btHX7gUEzn
d4uZsxDAL31ZH5om6uKSL/MYUIAHmeBD/FBHJyNI8ojvHGdXO6XqwKI1l8nL72qO
oyrlAakgSBOs3AGNmNrhSLLabxBjBD0xamybc0Wj1AIReS9JhpeQx/IT0CLRHZ+l
VbfxUu06DckMjx+s8kqzVN4Aui1ce8sipSsch+DVDsg34xvNyYdQKWzGPhgRkgMo
wtMc6/9oirCMU2+barpfFoS/jGee+yweUmYNs5KLz3z0jUlWJ1Gcernp8enY2lIW
dZcPECNIVX+6mi2TVPdfDzf/PN0gYRfXwGHe1160uUI7MzhYhY6pluPmVmkxKlzf
mJ1LmdxY27AL63RIPCpUo4Is3Xvsj3Dx7YeoQvmK7uxqEhwFiqoy3y++ChIXN1UC
vp55G9tqmz3sX4Lnd/4xapAVZkykSaeGWzOteKkypPEcMvfpAJPJx/m1CZB8jxBX
BrSipDnr/N2N4ZMtX0hD5a8s57jtjEFHAe1lUv+ksHEm1crxImVS2qL4Vw3Oy2tT
kVih72mhCAcp5uqvJOWs7m6QLBgm9+euzrVSvoKI2QJ5iLDufEfflnrXLTf6ASPA
6xpTCRrzdxVARaV3nvt3PCU9Wt65lps9+FEOEn2J4xIrfWKQTNmjR64VdsQmh4M/
O0NoA/fUwIBDcxPADM/LuKieL+7tX0NiiWKtG0390AkGOAnKI45t2xoL/Xjpuqq5
8stcV3WDQ+cg0h1rdK+Lro9caKh6iZ3jOHL5uqs+51QAfzGXTc4kWb7f69NSlVoj
VBvSAdGgppeoz2lCRcYwSg6SCjZrCIFjlkwACLTTceHXzhxRdKY+VT+5LBi7ISOe
pV0WwIx5Hr8eDcCsJPI0SY3xCV/shaEKM/usNqCOWcxkFspVh5b8PjoBfhGmEh1e
nUEL60rb0L1P2hQx8Gp9CK7FmZOni1iUZyjQnp+5fX5Jl/hMF3BGpEnVjjYprO6v
UW9CEKkO1/Wr+CD7OHJMdGNzd7rbl4V1Fwx+tuGMoSABakCFNe6ARzZtXBUsawlC
Kkl+JKl0WHGVHWRrRnpU1LhQDaN9qWjbwslw8vfHakahbGaPcLrtH1JGPcd2IyBX
AG8nFQYHyxYWCqutqn00gCNtUYIKTjU9Glnrh9PO9RhXs7qWNXliPoW1lHmVDpg9
ug3fNiMf+vho/DCJi77FC6qcHpf6kBXQSyaM7DmYmPm0FSoHkdipD2gb/jPuUDq2
bL9tApEE82vukWXt2n6xPowgr6YVh28/q4Gz/8cw5pOjPfCR4/fD1zxT8v93CGy5
bl6w3/+hIqM9mr8o8ZkcsE1zk0SJqSAMVouTUIJ+enTa3kgwLUReYDhZXcMfad8k
PPZaISOF3nd52dtWicOa8BEODazLwVFwesrHJ08hQYSsk0zmJx/pfph2WwAMJPAm
RBnRVry1xmPmpXEOKSzbfTxKO04LlqzHOr20DAyuz6OvZHeLhOXyxp0iQw5mRJ64
yM8Yfaf1zYpAepkA2Fdpe/xBK9mDnJwZB2Tg2/ZFN4VTFle7osXBWNyW5bd3cRUQ
ol/x2ga+K/AUp+VptxAI3TpGB2bcym4xbYj0B5KOak9TOQIsT6w0GMKQrYGG9d5U
B0rlhw55dLf5lwnVyiZfFRD0Ip9udNyhdgsCi42eU2M8TVPf7RYpucK/IcruLYic
PcsX8JnHWBTv9+a+/WILMKe7RNieNBAy9ZzKFH5EUYja54uhHlker9CWekLaUcsd
kX46oCtsIT8jFngl7yXsnFpYrqByNXBP61Bb8A9ZtYF5DjpTsJHCQfdLJSkkGYao
idUt0/kUtCmFqSob8YLLGBuOHwW7yj3dwLKk0eHANNWklfXmRtbq3d/qVGSZNeBm
lX0AKzsRMItjFXYvCTRtp/2z7C8yRi8+yO/NowTzGGM4LQ0Oh7vi0Tcao8tzPe+U
QDFsM/oy+Fzco8Dcka3OJSHV7ggrFtk7JiZx4b0JJmeQHsz9uVcCz93qoTgTsDbh
qv7jA/7P4QbpZntxQgqkrzzbzrHIof67SfqrIEwUb9QffCteEk+qW6sMhguKpdS5
t+rTGi13iAsYKQecC2dhfV+R7X8OsqB2kHNBBf72XitF2xmA8X4K/Tyu5TSdJgwL
IB9RETaJJPQmy5xsc66qLUw7VJf1pgiyihFhhZ0i3YWswV1tYG+lFUl9dwuxk1eF
FPP69VN81nk2ee41wRUA6pfYViWVWaTY1TvVLonPQHsMBxqZHGXHFPwO4A6wtm+j
gm/tOT1IViBhxMl+2xpE9OMmlmgtKatwH3FeHtKCcztf5YJOYD5wGFyJp7e2i9vK
MMMTA5AgVr603EqYMzw2nWaFqrzgpKihJ57Pe3dOK7szSJ5HW7qPOog7E5trMIXr
mHVratC2h3uqQMNSWaCkeq9ThyA1v0wYFTMi+fA8wuV3ZDXn+r5BvAwbbEuZbTxs
rhwVTUTVoeca6FUqid0A5wUsvQkTobJOFZPJKIbngu3pml0OmxOdJcSp4krUVsoD
6OiNOJw9ZjzSXf0gjBYF9KHSKhiONqdckWEh7qXVfLiT/T7rIvPmhRgISaIFOZOY
HJXLyjylGEPYDSfWldOzrmXxzbhlmFaTHrUf1tZ8ON5RkFuJflTdQTiCTRaT1sj3
15iichintLOmjAJz5fh/r97aPscz44pIkxFGLzE8+RpmEgiW1kiWBolYvrNb2d4C
/4LZ6Pw92lCFCEF4nhoJqZuoIj5rZuN1jY/oHPV2+QLHMyWRXdo56TTp3epBRli+
yLlF7ovVP6AwMj/Vt78caBSkuL5zDubbcRSRGrN5yzaw3htm3ntiTSzqV5MYSzy4
yUawckqBBlP6S8dv0qCV27TYI02gQFNxKsx1ZAJx/KfsY6NG9IEkHW3HrvA/TxqY
vIST+3MM6YpzDNAQSo6tJuZFtBLTYHYC4E0+/05Cr7pWfeYMHkEuOL1v5bu7V96V
NceaMDvVnV92X5iTYJIawn3+U+dy3WbIK9gMpUze0Hr+sFTju/Ytt9peSKNWlRnc
8HUNRE8+YKan0JLPnpviTX3QHQ+EmzcR2zWPVtuB8q7Vw0J+8SXuwyrqSiBB4Liu
TdFEbFI/OOEjlAl6qPUaJhrYeoxQ+ri+DzcaA5LxqFjlrguhHFZ0m2NcrXpEclwy
Mq69isGQOijPQVCGUeRca4nJUaeJQ9oUugS0bFjYl4gTXAjNq2Xzj4aMbCSEFFc4
SrVStAwJb+0SiLuQjabNobaWEUFJeU6RT/vTbFeztiREeUlSsU4ekc3cjly18IQ3
gLBuVnNAbFovqaf2Wl7MEq3rhKJiOIQeJaNGBVgO7OIRiugt7tOop5LSHRfrsKrT
x7TCdxQvgDjOR9D1mowABZR02qAXbDaxrcQwCp3KXrNrDVyaCuJeTF1GJDITgx1+
HqyT3bkobcWvCgu0p8r9Bs4sU41koDO42gWkyvS7f8Sm0JUpy/AeNjNm5BKdZayq
f+pi6+4eZf1NnNsBL0ycxYKlOpjvCBVas0sOp7tQcPIRMB92M14HXsuLO6VmNYky
D1jKTQmNb+3sSEMy4VX6yfMjs2dlhl2uLWR4bl51dV8FO/pMRSGINhenuVK/rNKN
RPSvqcbghT/nV0d3vjcsyoBVsiKDCJ+jRnDaAoEKvxkGo/Ud+D3F+f9YBaYidJ4/
W3fRvs3gw+yz4JzfZ9rZINoCZDgBdikk65UCGDG15pqdh03UL6BulTupXv6tnf7M
Au24tSih1T323TtzVDahQxS2Mutep7xyKeYFc64gpcgslPgy09Zb/GfT3jRjWE0C
UgPETdzrcshjr9JUEAOw7Wa3YJ1BrtSYpT8Qft7uwgOkglDl6iuWUlO6OVnj4sg3
1dM0ZZSAXLGMyDY935UYflABAQ5Bn6BcyFBNdQwrKWa/OUefVMliv+3uGyXCOYEj
kGjiAmk2ZCFT9GK0R+OY8SHEHmwXH4YlSdBCFdWjy8Ry6pWHToX6zvxRLofeLCw9
5kgwC6OL3MIMsVzFRn4V5UNA1ZToR+nLGumJfS47njU6vdbeNrD+i4mzvKXCwTWq
zFctV5J3wogTpVh/WE6StmM7xGKVEoJDc9WUVOtzuZuS85pS2FeS8Z1UFbLLDcWz
+5eHVWDTFQpYbYg1K6pJBBNjYA+UdGAAWSHcpV3+BtdPVvcfkekJX/ZiRv6sf134
TUkD2N5he/aS0fWzzsS9/4uLMH6PiZC4TrBZ52dhGzp1Ug4mViUPu5e+qacFFTZp
QJAuTt1Q4KGpgcdgbtZc6eM4835UFyzcNDJbV1q2mgSMnfekuktY9thBlkSNTVo1
MkJHBINRJ79ISV5Dk1nCX+baAByK1NrqiyznSb1PHpXecT5DmAK8j29EYnZJrpFk
Oj5pvIFI9AAJVDJ+a2AvhVoUKL3P8jgMqevXz9Hu64CQHQSif+uXeXYqXvHfgJlj
CH1S5D41KzeTD3/3Y51PRZQUEi2beY2cs/X6lO9HRVnx4lXwjkl+OLLpgdYKShrQ
icDbelnHEuoKDZ15qq+AeGhhb/oXSf1pTuYualSQ2ZAcAIyCeOMYTaaMWrtHQr9k
opGGR/kVJlUXylmPiDmcGw2OPHpj8cm8kLn2s0LgZdgVVOfJDeqQ+aVM4e3fvlDR
O3tg6iMBZvYo/HCNV+qpJMRXHV5rdYSOZcwqTrtwisyxlwd2a9QqKbe8pLygOB/u
P1tBlclogToNlatghUcCPbb8BDxpFDyAq8EWTc1/NHopmDJxJJlMI36l7QJds5+z
Vo+0QVQ2AJGMyQ/NpMrgokZg8LZctOmI04mpFPkzUdBBvSOEIVnHUO0zuOm0d29z
fl0AK22BY+Zg37nF5rekaryna/HG6pvLTE45fTY9rp5Q/f4uUWf0Xj+cTk2DFIPK
cqqZvHp+miF8eIAVueClbB+bfA6pfgNTLG40RU+0AfPYXn0iDBBjURUY5T4iqz8D
PMVp62APaZasPrCdmq22UCKDXpfJ3bGhliAbhQgdZwynEYcvntrS7LSlpfekXjer
7l2t3D1ldvGJQWNHFfwig04I8iOHe/6+hDALKCQDnil4iScL7hUlF7YSL1BaTnS2
xcZRokLHTE+5NygUAIent9zeGfutULsDcjWfccy6VXR0rD1PSVniPlGrwQn2s2Hx
QxE63/4XMrra69DHpstey4E6McVLPYmo0Y49AoQmzgcXfqm+BDL4ksSj6mUEPp3u
7+XzaBPU7zL7sjGmy9imktlPG7PVfiPBAug8yLjar2r8f9MXv/NZkmMss4CYNprR
N2aEtk/7ALzVRGofb2D8FYfSV0AKpvpdjG4ok4/rnH6gQiDJfI+Kgyoj5VmISkBl
EDum0eaCr8dWcprKaFXm1f8mldX6kUrBBWNbW3CE/rNILPi9yDDdy2VdGm/48W63
Dt5KBVftml99Hr4z3akz3/HUVg1f1Vu2EHe7ZAWH4bkClaqHd1e3XLVca9LIjpBW
mp9pnhm/350aDik5UeJOs9EgzJyy6fildmcEw5szgNJkKlLoSw0a1efNt2O8sYPM
21VHEM0MsKMm5lZwQOS/gUmFAIp+497ZlrajhfBYzPRQHVrOPh9TGVir2k9E+7o9
e0KLtCaIlKQ2kxaIh8mK+vQ0IenZz5wqfWi1z+1e9vqmUxiZQFaSzCulPnNZ6gLl
8B35uZyaP7QxAR74aO8zn9kufiwpIrVNFUrVdgkyu/RNCdBFB+kUUdqkeUi/BIXK
JwouF4nVFmFGedRIt6R/p6U+OEPrbsaKP6vG9f1bDH4Y3xvHifwB2NYkvRxuiL4W
9Eesn55B0/+/TuFywuqDC+sPswAe1ZTTB/Xv7XxGunla+Bln3AhSDiqjThWAe58m
hBLRP55aQuE1Ue2UTdRq9hWjP2GmUusPvg+2aYL6kMPc3FKGmjIOW/nCnYwFZ55o
DXUl3s6VdgNogPxuI0+WtjyelDtQZRBo34Ir4ho06wMng5GpIoXfgJP81y9jpIix
/Tji7Am7OiKrjEtO1KSHHXffp6nPB7etbPrfFrLPewcucnn77CRooa8CeHSZbcvm
8LDkBMjkqNnuJkzHdmWO2HHLD9alRfv+p5QzXpacOsrdvLFDVwS1bcwyz8Snqr5s
gieMeJKA85xPmMItWSTASnh98cBsh/pzAO0QaMwWgRsfoQ/1XRgC4q2e9A++3bOP
42CU/VuginPcZQFkHeEwnOsmzhmeRAci6XLskbOy4ceeuGehuJSLnLIPGMQ1tO7m
IIY5peJER6200zl4OjrWW45tby/sBo+wwandDYTy5lECJqpccWKqjYebZu/vIlRS
vZeXV59fj5llLd/xpQL7v4ASgWPnMqNxRL8+4Xu/BvzdDvFH3FISsdOYuEhOrq0O
iSpyVSwpKmU923Ai+5QnmGTLxAhzSLLCS/yCVgyMN6QLeX2VZajTkp8fMaCcSgFP
zyHk+nt1K3VredmQk7HxSQXKTrtvAOIGHUYljzB1BPwbsYAHGc2j05A6M7gRKvXS
WvkFGQ524bwf9zoR08F0CkH1lL+ak8Dq0GNGduNR/+p196Q8rIEo/9gFTvPweoIJ
RJtW0M4BD4qyPGfRfU0jQ+U/23Dna1O8Tpy7h96pfMl6TXcRTp0fPgQzU59lCzrl
TuJdfYF7XyrjazdMmXbV5LKhGjfhtFkBE2Qks/hpeQJvVF4ZK4AWFJ3GDTJq1cNz
o9JGVysJrUOPiaMboo2viMhnSxXDKaoEa2ThKM4d/YTyYhiAUqGWFyppbUAdCLoH
LV6Bz/lOdTs8ElgZke7dcIWufwdZTQXqOfF5nVuVnVDmC0ey1sCtxRssVrjOQHvv
Zze4Xjf6VLemkowtK52pgeDMx+B9b9gqN6toq6Za9gb2fd4zWJL/0OBLumdbaXVv
ehThRnS8e9qBVKeEPd5/zZzYeNYeqkZcCl4LCJ6aJ1fJvrqpbNMGkZqJXz0k8/a5
LhlcWTqyr5z5BduQQwx8r+RzVLeq5v1lLZbaTBh+aiedq7En96NTuAf9asdEtImI
jeB4ENRpPdvX9b9MKFW2ROeKJnvruMqRpLV8DN8y3HYcmcG/NSpU8KR5s/zAoDou
iYs/JSLok07Sx0YOrxAqFN4tFIGYiLoEi2kOIJRT0mUyiWH+1TGfqXh/znaTtMtf
p2AAiBj40m+DL60AW20jMNDLwfrC6uFHbMsHkl2byN7prp/4qjWHjIF76w8EWdnT
J8IfXP4gkhgXrozy0xwLbHAvFthjrtN1FvxROmwWBC0CjPCRuPQOh2KE4zZxkTWh
spKlmNokX5QQWM6Tm8Ve5oF3emjclF/uLI3IebbhG3jzvApCItirr2OJNxsIudEQ
HCGjZdujMyKSTM92QjR5RTcYWciPNLray0dmWeZ0Nc9KsXIH5LTUrBzBHnsTvLM2
KxCUr2ZkRoRjw8RuOIQEX8Q+4ZRqSU8DkTd/zS7dzmHbJOCo+CI1ce7bPUPByz6E
dYiD1ha4q2FKs5VcgyHzl0rsKRw5/jgHNfDnyWQ5Z9nIHunI5/fCXXLq2NFh+YF/
9PsUJfdMmQpBCsA3Dca7eWlu1yOZ9LJ8J4m2Ky/l9wiabkFu8er307TLHuusOBQ6
tS8K5+h8JCZTqCsJlKIVIvvwnLBeV3LbNkFVJE6f6KwgjiLev82+/kKR1ZFVQZjz
sY8EMbiYIupT9tN5PPg0epZEnzibAWXLgW0fuLXKUC7UYvnJa21dXrXYxT2NphXh
v/L8pYojiYu/5dqCNtIiudjQM1EYJkhhKssU0aJ3l8STMURT5LRLqMGRijPDjZww
jk8eVNZ0eNGL7Q+d+VD3IJmnhAEtF/g4wQ0w1CwZxZlilU5ymEtHO1g4Hh1d/25/
ihnMQnv7hjREfN3Cmkbyfk3p4QKcKggmlTCAvrYA8aUEUvID7GoUlyeDs/Bd1ddS
2rUkPkqVLo+MovNPKsQt5aLZYqsHP2gbW1TGCTWvALPGv67pigIdP+C3MbCbGhPS
7GjMbwx6BcpAIaETiEPithyftgmrYTdzA1RPKGfOXSeXHHrG+GjmjF08i4K5TirQ
CQXwetWApeqlVBxQtTOZ6eCzpqlCoencRreMPDH9ZgYVBoAMDbeUueQyBuTVqNfO
E2Slib5VX2lkV86lmamzw6DoWItBxI4BDMD2AVfXyCIJY1m5mybsl78sbK69aWv/
SeMcREzeQajZrDqGyNms/toNHUV6r4j0YtWnen/QKWtxOuyjOig/GEU7qRJHQ4Ur
c2FDajSVbWAk/y9YreNpLU4N6yCrm8J9TRTRSSikg8t0WtRNvEZjfSnKUKNlS/5F
yXEj6iRqrvbloe8RvaZ6InL4JqXI+n6/nWN0c4lyQ5sZQhUnacVCO744YCsLMBg0
0/f5FN2zvEcvYLNhnT7pNaYaUUj9XzKq8RTGxzslVzljFeP7B641Et09+MXDZ+JI
34LcUj+CscZwQbzTB305n8wMFzoM/fedOfkwZz9RKs+EX/7UvowkCpwnP0Zd5z4W
Gg8aFzQIaGiU44eaqes/CGUSlJpag8gVlBT43KPw8/I4fjLE5wMxoPRxyNAE8EtE
YDVw2AoLH3JmF0dH0JprLWsauta6kDCdBgA4/NwCqXhuYttdZfLyGJiGuETxkBKs
9A0W6faGApzd9uqb1jAudGvHDmHCmLUMjeyFgUayLffPMfeFJXZQZMMD8LMtMemS
tIcb3TvmwyL4AxPMAO6i2BAKyetMxssjFxgWkgSCM0+JfKdbOYyKBy/PZFVqrvvX
Ux5CpGn7wdQB+USem9bNHQhy64LlBrJXylMFAIbZzetO1nelxSZWofqiIExUa+9B
h0gm/Hq0m06OP6ksnqokwLYy2gjWlCuFp5vdweq+aCx8EqeeYQd8Rw0DyvvP6UqB
cy5/F3SV0l0avrKXqnJd2+2rnbtt8oEt3v8RkTbkpCldEBN5kPRAV3GVzxFHqq3k
sUdTp2FPUrpu7fGzHC4UMB4cO4IxZIeRNs1DnzCOhyYycagBnOu/9LoDQwLhrK48
GKpQcIBOLVM3Q9I4jh/jNuaNwgtOG4MPvMA23Otc4aa9XkNY6I527AU2AgEHY2YP
Z1Fk1fl4/UvdayywWAid2Ff++8JarfqRGz9u1Tezm6IDcZNMJXqdPgL9ZaZOJe62
+anTi0SrXwdjta+5twYs/pZDX3UXtcDcBbDQl3ZbpONvVZvcDh+Kfa5CAj/Ku1fo
mrR4lF/abEze31sN6duLTlQ8+EWFLtDgf97H6Q9ib3IVMUp5ooyoDP4yX70F/XBk
b4HrqLaduKGBA1Ir4/Mm7/yKkYSQBjAlUJPi5+s3Eqb7SXa5qSVULDIktSQTAbyE
i5SmaoWQPiCjnM4IqGgeTVBm93LCUACrejxip9VIzkZk1sDkJVBNuE5UGhdxx/W8
vueboWewu6joVhxLjHST4edNppboI1v0JJDcK61P9tHnepyXTESIZzkLuAErbDHq
s2sTplZHJ0iBch6eKMdlxc2DEQTOJe86I2bDXPoF5eCTYUDc6Vc/HtbWMEMDKKYq
1t6ZxJkEx3GIREt1QZ7Z4NWlBDf6YWJbhc2hOMCbI8P1nqX7jaR6wCxGVuZl1S5O
ZeKQhvWGIw1sTZvBVMzxqypAFCfI6rai42SSCL1dN6MVmPykKEPFLNUMpOg9+jTK
OGtSSa+mUPDdtM9h2BosFXtV3lXv4i3LEGkdmMpyID0iAO4uIzd5iIMkZf/Qd3pn
Ia5FXOGnfjBp2S+OQ4rtXs7GLTOBnd3oC8WEVtpoNmM9YIZ/km4ndwuAJEImvpCV
EwoJXVtDueThKOHMKvcMUDBiYk3O1rqm4Lv6bnJJhdlMBnuxBO9tGkh5TnL9Ahs1
z0DTjsEJCWqLxpp6Nsvu/K44EOA73KeLxxvH2wEVMuOS7f4bP789iAZ8eWKZDvUD
b2EQbN+cXDPHxY7E6ZcQ3u0EsfiZJP0n/j1oK8ADyRiJXrvBMOeZLto23mIhjiKk
2IKqARo0TYcQ4zHg023197eB/kqm9+BACZ6DIe0+Ov8nBEBf7NxfG7zJafbxEoHR
qgv1uob8X42bQK32XEujTkrdmjGh6i8Pc15roc4gpsw/XnI/OoBVm06P/vPnbobZ
v5s9HYl+nQENbf32wo/vXp5F2KE38Docf7VtEwwCLpZkUaLtD6R03KzJQgxeu5zU
k8gRj4l2jdLqWLJCgOpSgbFof0JgE5iO2PdP3moxWKVOVBkfVawF2tp+HrR88yIS
Om3w7CeWZSsq4CkpC6dm42J0X4QT3v9wECD5Vy92T+ZdiblssRf5Y5FbAuMRehfv
rLaha6zM4PmyeCGffzw8DkLpUke6pAn8pbOeuOF2Ff8Kn9p5dw1wIk+14EBBXy/J
UNz9Ysh/NnXfKlwtonOusEAjAZ6iGDorHElBOS6PR2POttqY/5AeqLR12fsAhxNV
nvRfND2sEH8bUvmvCK+02ITBcYZ8B/FJ8rUI8uA5SGsbjZ4fas0GwXL7VogSxILo
/N5GoxiR7wSkR5UiRqOfbTmmUSDGZ+mPEcANPuZUlnNqyBqmwb46AI5xhI028L0l
kaQYYOe3XrOOHa34yqq7KRGuDumBV20vbqrloJEEsfAK6IiKT/XaCbKfDhckLbAv
LqsFnXKIq6LxRHRHkoGs/a0CBALlbikA0mR/nMeqafnI1dzwy0wjoMtehsfA98sm
ayTzZTKiJ8255LvSXH//1aDbObixlAr09fUldqw2zjCDuCYIH+jUrI3yEsPsAUJe
aTTsONZQecnOhu+UQ/zx/XBBBuhkZVTO9I3v1wxGq6GwtqmvMC7dKhRjqJHRTTRs
zeNa7wtwKlqId4DwA4MCxida8TrL9Ak19TNJReKB6uX/xKogRqV5ld+iBGCnrM1R
OuAG0UFNJoc6/DXUJEphv6yngIU/Odf0Lr2SE5O7z5KHmqoZWRRqHcY5MY4UogVe
tfkyGR/VEN9ImUoLJUyKcpdu2tBCkSKdFqSDHYpAj++Lg0DF+7/dH3Bu3ZwoH5UL
shcr+QEhqVIZKAfVx71diVEzVxqRG9l2Br3yev8ulh+8acceEg6ScRQ6i1ikS05K
GXHZYp8bBRro0GVTG13heglpjy2KPqaEk8QhpV2LtwYQbV6PA19eq0PSS975nD/p
WxK7qV3SSVMfM/tQAYljlQCylfpIBW2AsCSHeZBnpNxyZf8qfOwBH6vkEqUGmtbT
bmVaXjzZnCizeJGItttqnB5uwZpyu7NRKPZBTpJ28kg3067RkXDZQpyY45DEV36A
B4jyKtMyX9fM+twhfbQR5WK+iSKQ0FpJO1VCxRiY4HyxHzyW7AxnAtT2XIzJde9D
W0c53hm0fpBMJ97DyrBTRGrVNtyooOnJie6RvFurhp2YslqGI4uwvlADzBefIyrA
lmp63sCYlMMvdJkwR5ArASj1Csaf3PhDtKDDTJI25+2v8qJfufLT3yVa+lvbGvus
W5nplI66VZNwrwuDLSsyAg3ForOzR4fYpH5h/siXKgQfixRm6De1O3wRVLdg2lB1
GB5BrSFjeTlzWij7m/Q8xwqa22ifVeE6rrHPzkXBM5jndvO4gQUyQVq/ykH9clMh
vEAMUmdDeslSE3DQJxrn6CcX0+BDPLrNIrg6JLngqNO3MBjbYDN+1myGFM5tzeIY
xx66yCRevxaE+31UcJGlmpHoZyJE1MbQYfTDCnV8XAMS+XrPbg4d3N3P0hDBYNAg
1nrkPGJKHXrdlTxkAsP7Sg9jB0k/dp2a68fDRNs5IyC15eUuu0l1NvrpyHTTbui0
Q/fZUbYku6Wa72PDOdsczn+M0KWSBnSJdJQVrtTYNUUm6Q4kQEDVEYTrLfs6J0/a
Tw4vSjbea/5sWMUNN4/KTXBOHYwuj8cb0yZvgMNokLM2k+UP/Gdc+xA3CqF+6ooY
I07guUFPNFiSX4bHv8VWYh/GVRW3+z/iZAwMJ9aYq2DwFnH+kcCCNo2y1w2hB54d
l2NSllgDVQ6iEitvAnaLhpjvxKBlmgHSaFeFo6Zdg6tWIFrXMOutgSNHmLHqcsEs
st6DSiwRNnW0+Mh0XhQNw/gu0mudYpnz0e0w6aOd7uyGFTbzx4iK1l/fusUqxfeu
m4Xn5K/psMnR6lckj4NgVhXs0KwUReCVWquw7XNguWObv7lc8r38ehYdSWC7tllc
lJurq8Zc4GaxhmwRScYTGUzlM1kfIIzJH7xSBtuOIS44YTJyix+cQiyrCtnn93Hg
rqZyJsLWSpI4YwC/8iCt69jsM9PP9kk7e5hEN/P/QOtyu9Nzz3o2jNpwLa7qM1gw
Z+U3ICVO5dFVXp1II8uQ1J7pAmwlh7dw+iaAdXV4+1g511rcL2T0mWUx57hIDPvi
d8kxVUnaHWY6XSkfRDu4f8CPZBDMiZ0csYKfaCF8nAQJeXPKfwQ3Rd1R5/3CGKxB
4hFUaCR5w++Ar3gSjL+XbWcZChmotC5RI+5lR/u46GQzvLbTkfwiZYQbuaRhkBpx
AObhlg93GwKO86xBcMKDuOpdu9O2sycZV9OhGPAZQxX/1KBn0ekYG33JSNmt7Kje
1IW3havYhGYz8WE8CzwwbIE3Mqv193pdBP2EL87lnF4onPT9qpYSjsQcjkQoAIHB
T33LrRnZSfqzCVGsXmnLwxeeQvCKYnL3IBtLcdF/f/dBVlYU5kFH4R1wKXYPgHh5
rO8O4denkH18Y0JMqc146L+TsbXltD6zX+PBCGDpJAHIyb32xw3lE3jDNwKo+6A1
DV8jWHgC2grctSee5qIBJ82vK7jtASIKxzHXcdzqLI1Zs7oBGHEK+SvBoBmLOHFz
g48D5BntPpjZ0++g1cG2jYUXlU9In+6MCyjoDwGxDQj/xFhwms3PkkkYWfv76Nl8
yxFfA8kldPIj3IvW11+P+fvEW7bf0xE+ItE4qLRwFdLEY/gVeP0i7R1XmJn0MFqz
CTSnhq2o9nUl3ZIyVMgRMTxCgpUZS1P/DrehdPmwMSuQ2JWE9fdgCoFO8JQzzpSB
ZjzRbN30W4HbCcYeQqT9PbbWe/4lnwZkV/qk9rBXWwRW++666PPWEYa9MafFWV4r
+4DW5PbxuOqbfs4lD7Lh+Mde1RZ1Ke0J6T1d6dR/Jz692cUtAXxcIto8R01H5Pr+
WG/IOsA4zOZOsiNagOCPa4oaSGgUPKrHILVSHNWozbfWtCv9WFtyK2lfJsb/kPry
tRxjbOdliFeaqxiSilhOAGpU3NaJPNgPT2Zv6YzQrpRkgxY05SKvCL3q/rFcZ9Vr
5eqpZp9ycDumlzlw3qsNyN+6pVgdHLs+bS3Wy6h3ZiQukjk4MJmrRErzPPL1UqEo
fEC/1IcayK7/euqcAkBZoJS4l/UUrvi9NQHL7XfoSlXSWh/O1eBB0TuYt2qPfs9D
chDszDCVgnn6oGaQ5ZgMVQ0OtxP0PJDqJ4ul8wATdCrVCwY4x29Xu+sEmGE405bL
b1cay0tge/juXtFpk9eSxyfYhQ7+hkrKrq07JCSjn0S/4y5kJvqpm13zrJmD/OhO
vDxmR+SawuP9zeJ/so6g7oLFKo9o7utgx5FLusAKdiiu5cbU0vfrcmouWzCo558T
bwcwn3bO/lkcWyvFbk3RIAML9MFuIYMDP9nvYmiGsSJiUYmltoS1hNw6puGQa708
dPmAn9mF/1fcVIuSBh0bB84qQ9pzZfo3p5rTQRj8QKLmAUW70uXFXjInf5PQw4v+
oN4W+aomZ/7gNVuI0oCHn1l0nMQdh/DVC+TUreyqljdfqt4tTz079wnd+pLLUvv9
vuadNUeSdDkj5S4UBLzdmkD5EkVHa9PRKBL9lMH5fwVEocG7v0Tx+07vudw7Wick
+QKC+oRxjRuTuQKRZcJDzXa7VAVxQfpc+4woqjDD5TWrNpoNUCX+rpn6vKZfXZ2F
iIE+Sj0RiAUTTE5qbuZ+/hBmt7rnTyIFtVmvBd5GtkpFXGCLZ+Z/TL4vVAsZzJWq
68I38aYVJLCFhrvnV45oCHkvLAtMFX+744/TeXaYWE6puG67jwpjgWtfYhuQL/yD
aQony5t751j//MbMEYkAHeYgSywMZ6DJARt6WtQx2kSnyVt/AZbKWaL0jh/QYkF3
mNfZ/OKYm+t12P4FTwto20zfl9QqrUwLhIgoRUEOd0TS7S62ACrvIVryC3HDk7g/
EcTNhZq2YrOWszrYW34sEGrR+5AaYiridrloIziwgajDyJcMsQ94cnybZ0Gd3PiZ
S2Kn/MxorDoQGAPmsAvKNOZI1jFWPWQs02Rp862syAU63IFIfuDQYxgwra2Qt4DN
Z85f2hJZnDyduBE424X90DECMLp4fIT9Zjb7KUFdaqy5F91DZM9hGysru/w2s6NX
/PFdHA/Aq7m4q24UC2NcwydjESMdTJ2EBG8lMMPhV0a/eaOzm2AePFK4He7cn79o
sReD377k6XOLv+lJqyzXrgLsNl/FSQyfTfaQp7gJOw8Pn2kWq7W8Bt/4dNQdMSxc
RbETCMRFiNb12DO+FnLgloBGKqGcNqzugTUF0WlRQFRgH+esvdvViazy2SMsI949
igJyY7HntYs3A4gaH6kEVe2/R/M7svbjl/fHAZPYaHY3ioMA863cxaZQnxbMkE46
mtbF49wqq9Ynj4cco6h0IAq7qanXD/D7njKNwjUrVPSOFSe4ZoOFBw3dWxuyv874
yNtJOvYr6m5skIuNX+3z36/f4DR3I5OQZF3V4V3hqMSSAL264SM3EQO9/IT8i9bv
57IoH4qi6Z9k57CWv21GiXe4epiTve2MX5aPkhvx+VHDDiwC7D67aq6EW1HX1wqz
VIU4FDzQEoyIbve1gG6STu4FPkDw3rlXhyr8aCQfviFHAg7qpv+qP1yqmBceaPy5
vAVKJjljtklzzaOxmLIykA9F3cWJWBJcAYZn9GuhyWWIOlsNH85WUHzmfdrOUSGq
g5sWWjRZKiHBFRag0PikIxbmRjX0V1qdakpzNK5g5MX0yspG6hPndtkHQZ/K7QcY
IZvKRQUR5Qgmd6AfYl7UjkD27SGRj/V7UnsEQTZbX2i4aUr/3Ztb8OQlUAcTcz1V
HZK078X9vqA0DLimG1ocHy6BjX0ze9ZG1WkVUMyUfkQMHkyqAYql07r0KfVeSlCY
4SnzBIN7qPhHvOvwmkj91ArDoJN5+gV2FupHO3NQa+IU2yx833z9meHm777mSwUp
YWXBaEj6HIUKNrjrTR7NJcLeyKst4DJIqP/OezGUhv6aYDZdGaByhne1ooDIedfn
Usl0S8ZK2dh5naZ+ZXT6qsER3W0MAjGh5oR/oH3n3M0Ud7Fakx8sZBxPAtX8nG4x
xVdulenYHVqnGC9VXLRvv7xprEHwY2y714wMOKSoZYy0JNv9Yuzj1w0Ey9Rrj5yh
d94E/L9okvhyJZkMcyiiLaaShQKhtiLh/sEA2rAjTvFCPpd2pT2PSOk2kUTbjUXq
TZfGvb9LgLR8hW0j3qvziOjGNQt9N97xmlzSoWHThPqwDbaLSK7Zxx06J/thVQOm
ylUEb9MSP3dPt64S5V+1x1AKn7STV7x313XmoJ0xD5Vn0eQKJNMoCTHxOaCiahC3
BL1hP2M0884LCwPzPtz2CtFv6NwbSYrLGsfu28FGvvfog4rVgBHJptd/mfu0+RON
pMEXzB6S57fNRNpMvcjPZXpu8CeJjwDulWVukWZw6sZZCvjzUfEqAy2tk5qGKYZp
jbaC3R9vW6gLF5aNojwVMO0eN/zFrvwlTGdJoLzaHNmo/OvAsOduq2GlnAUuEJ+g
fWDeY9wzV0SD2eS1nUXFJUj5QN7wPtFNHjOD3cI6j9F3MdpiOt1l3I2tBjG4BpAD
iIlR335PPkNld79zB6ngXZRncV6lkZfD2cD4cF1C5KDLTdlLEP0seFa+yhCpxdTl
qDUNAqhxT6jEmYe/A0V0mOe2SjI+LRuBskVhxkj6QmRq8wF5xtM3BeJxsqWFpvsV
rJGYo1YfhE/uNC4xxqA9ZXBySXSX+U1vdReugAmksuj5PZoWLP5SGbcw6hgZimCb
g91mSW+wnHOuXEYwiS9WPLRo1O+lM+WF7k1wm7KlKWJ6yLg7olzbDcpTJVIbuMr8
iKudBR0Hlo2qinYaarBIuBO6fn/NzLk6Lw1UCkwv7HxcqZWPFW/LD8H0llsAaSAr
C6HbvnHn7ObjpYXGf/X5FQfVZbMmvY06Fbk91NtVfUSTgRAjzhNhcgDIIiIjleoY
d/xEFeKIju/G9i29MpPRM42+Ton1pPIs3FM9D7dzCxvvaxwKLo7+WanY1fcWsVQJ
Yegw9sSLl20CxjjsVU1Pk2yZ+RupdTesbxKFkmTEkZiByUDKZVgYh82+VXUDiDK3
t0EqkjBbHYFeJidBRyaHfqrqs7ygBjIHucCXKrhRdCbyjSu40eScRPwE4kMY4O+Z
a7VttRLbNRIm9wiVTrAfi5zq5+i0aeF996T0k+Hm8MBQcgVa2VYTShBBQs7y8gN5
frdWJNHipmviGDzMV05ehUbb1dj5LQNJ5+RwTgnWezXFq2E2SUGZSQTuU1Z+7ddA
LGDBNhxWbhDESUVyp60xGbaeqjF/9MCnIK/BxHTIreMEes0aNNKhdZU/0z1k8Hiu
zpdApPSU/842gQoWKT6nhiFg3w1nrw7ALDEc2+MHUJ8cwWMA/VBgzXuBcMyGUPhM
4ZKtyWRSsLk9M4kdv8Oh9tLVzBkxPaGUzHXUOVsjmtht2zI11KcxOVWxYOGu1sMM
qsH6s8TO2uZ3N+PgytYIXN7esMiRI9g6GqMZFQolAwTHa/JYntgaECpMxEcd0JZS
4/Cqf3uLNnOXoCEjqI5p0IQalJuzAGKSY4acb3MCJApUY4oHIwisS2475Ayvw/IP
Pfyw+/d8Bc9FtUmX233bdEcmm6wycjrHT+sqvzr9NHU6AENqdL+fX9Rl2HgfzOwh
VmNJnQMq4lMsGFJwI5ugLZutVE5DU+01M6bLqdQ+/f5xKBpd48W8KrGhfOrtxvAq
svS6Krieex5ixgBO7nvVnCl0N6lVzZX7tjw9M4Kyalq6OJTgU6keNdGhvDt9J+N2
wuEoGTRypDHl4PHnM5sNaaIj9BxMtQlAzX7a2Zo9I9RkhRp4Zld/hL6E3m+Giplx
GiUgcQqzKh7SGCL2k8k19ugYcGi/A8yW//as5zM3EAyPXwEFAqN+5w+T6kL79Bfi
ggC0/OFOQL4HwQpv14GJsL6eITLt4PAiuC1bB06OeHSkfDWQ1v/U0rBln14N4/ft
j97lDSx+ITwIhop5lqt1Bi1ZU6OXJse3HhY4E8ZDIEhyHndNKXbTL+cIDC4fZ9ne
N3omxHKy3hdRpfCm9DfL0BqVulmYb1tehUBasHVDcDXQeBb2mPeJtARno4lwAaxC
RdxVIq7i4d7hkciR5gbwGJp19b7ioyN8648D5rBnF1yiWu4uNXVW0RaTUvzWtxBK
U1ioBjKDcibTLXlxsQu9dIfy6WgRqq61RqwJid2ZhH23SrIUSjg5BkpAMrts6ksw
9Gn+lzQBQv9M8mm1XkF+GKQKja3oRKy8l62/D3z9bAaPXW5zeLKcyb+rQsaorSiH
h8RYZg0Ft397tTofcXAfL2kuRkH4GbzlKIoipBQUy2L6V24DyXs0n+XAb3aNuvFw
JrV0wAQ0ZHvHo2yp+P+YDBI9H7IXL2rg6JOdXugDz+7u6FaCHRNkHEeImWSuPWvn
kDW5VBjWt4sEsFbOhCbgZkDZwR4UmyzRTaA59OqePAzNHLbjl2CvWyiyhpp/dR37
TLinQmcjJ7yjWBkK+ROnh6fkVaJoHNqnXI9C7LfC6Jojl2ts2LHNoRmOZZ/4p9Ot
sozlTwDOBJ+buI1BH4CJyGzFQhhq3xhwWWyKubD9vY6hcWiU1hx+lopb7egsqjhg
/v3D8a7J2+QsLC7jf6X0oV+59JQXavv8nZPQoLtY6s6X/CkG3yTbW2I8KMbWwmoA
Kra0gIBYdLc3/FZqRowoK1zutGWIv47q+ufHnyO9RPNB/l1f2tOYzzTu8/Se6Qrc
pstobFu7aOnR8AiqB12XchUrKZThhMOKDK8AH0ILQ4n1JH0swdNUJxVHtWZqmvds
z9pwjfFfQAOij2KivHuJA5UvBBmlZQ1h9RWoNzm+blRtYm70IIg7d+f9dD99WqU2
FzQ92KzeIdC3w7Pp+ASDPSOolpcWAYdIiZ3oVkwpF+DZQ25f1Rvg9l0HH0S177s5
RzqyKXdpUnnx1XtMh2fmEcSG++DX28Kce1ty0xlqRnBYbBuNCx9YO9qPOiy2rJLD
AAC5UDgmYUhsL2TNICdnuZBf8pwnPNZ5jD+C110hWH7S7bu/zljCyQ0AuFhZZ74o
oueBHO28X+0T5qoc4XzsI2rljXj/O/G9Anlf79Ydilb3TXOENCz49GxGLWLZODge
CXAIEdQ2JQznINitqHMEfYqrP3WFK6RCA6rpX5k02pY5ycQQGt1SWVS8/V7hFXSA
VL//7pitZbeM6UaVhNe/jHH6yqhDF51LdHh5D1r3giv9syDbVMGCmBXWf/VuDG+0
ikvzZ9Dj6mU/X97DSylOWrKG4GefY3uG2pywp6/3WrbvCc6cnLzprHQ7LQ5ohqwS
rUaR2Geor6u/18DfbhmeGlrmnwwZbp6SBKA9iQ4wJLmMmpYXgp0+F+D7b/q2aKTG
Hv1xfoNXpVgwggXZ+267+WhebgctUgiceH9lbM++Rx0pE8GRE/a4gbHczhca1eX1
qj2DbA2hnvUl+UYXxGVD1Tx68scdd7Hz3+3RzPeNUhGR1Yub/Kt7IA35QSW+lHSt
yz8RGo5KdI8/+qVgyZE+ASb/vwWZ7+pl6O2H3qdIyz2zpo0dWpGE2sZuJgEaRLme
wOwBWvEgoRv8W9UQE0ohO+Sz7DPyN3beuFIDEanOKcTlIYBMJCZjnAz4SfD6w3qh
51IkpH48L2AmbzVg8hUFJ3wehNPdzu7SWbc0y/Wvq5FcunuWq0qHwkC27n2R/srT
RVMg8FGrTSIvjgJcKV+bubK2Lx+Xgz0sm2AaPpYxDnLYLtm1QbKS8KC7lmRvPHVh
ghhQvnu+k43M7vYKZrXnXTRe6B7qeX5+xzX/o+tDd/IMTDdgAfE1dAjX06CBQwEo
sii9UTLFFs/Qj/vSgzOLfZzZt+PQihCwBDC/oeYlc6xCNuYbNg8eSqopSR3cKrs4
gXXx9p/+L2lJ5n2ZMYZRSWdrm8J2ZnuW7U6JmKWCr6r7Q/GNVY0KGPUgrqrdRbcf
yulZWb3Z2lAU3Doxv21xemZ6VE0KV+89zx7Lmc/87hyZ8fw6taZ9fJv5LMUfzCi8
Cr2RWvWGEee9TC3fMrUSh46kW9vV12PzHKa8ZtogkFDFt+YGVbGRSixWRHmp8KAN
o4SxUzjG16d9QvFCbmFPsu+Fc9Xi/zzXYg2MqAYqFUs9/Y2mrQ16fDuWVYi2fOnd
dWi20hCQbcnhu1w6hzrvK7kqWkrZaPnVv1RGsJOK9p0e4JRX4WPjZAlr+e/bAo+Z
JcT7bXmc603FNpdnc3EIAE68BYrnX/q1F+18lD88MlE5VdCEaJPAp0uPmfcKxsx1
c3X2eYHTthaZez+gVF8cBRvBT0xgrZrWYZnNz86vex5MONRtZKXE4WBPG3EqU9Xh
4tpUG0rLDlRrEJBDur3ZjfDfYYdzmbcK7vQKgMAhC/e/AnGki3NBVCiuCFhu2833
AFt5+zKxqyR3jNKwGml/v4v8bFIX+jQseyb+EVhMJNoVid5eQdbzYwOrrv9bfP3S
Dz4L85GsjbnfccCuVz4N38fQ113XiA+Yx07p+yqQYZ62XZsweyp66uMXTYp/i2Cl
LT4somA2wRhnXp0qvyCsqb/LtjVteU0slGrM7N2ybinM0r3ByQwJ8wiKMDapXUTS
1iukwK9MotthO7HgraANRPnA0NpcYj3TdZpaj6wCNQj+hftG5TNUgrQyeAeztUwc
swCeuT3p5+F3LJ/Uo4Yf2WXUhx/wyhM+8rT2AHgGm/m/Sf7gPBd6q+x5ukTirA2n
+ZCqtbLS8ff0o6DLHd1j/LJ6XJP3I9+Fl8H697UYJ/gJrWbuhpqiolV80NyzNmgs
HY4m/Imkwk09fG8s0+o+lDYxFOW4dME2+w++0t/UBYrjvs6csZ1YyTB3jKG5rXLY
tIxLquyhI4/WKYYN3dF50wit7tW3nZtzS4Wl3hibrVNBV5zn0C3PZcS4RjZaPfdz
rBv/V0MGotTy8s3dxEYL7Ptva6kwbnWAicJivHoG6HNERrDSc7Pesyv7ZYNKA/Ms
1VS+zi+K5DINkk5lIWrDPzEASPPetwRD62K+v5X01IKzmpF36yCOI06tzV4jruE5
TbmK2ZIOPJmR8alcCfLVx53NWSHBybErr3wpmObKcpMQztyBtgCqxUMPhilxgb6q
7PnrWgioERD3NqJCu0Q3e++UFX/OkQmjUqMZFC989Xks0Ukiv4NtX/dRyzOEwVyE
0eB+4BGHn4jBWLVRMhXc1asBCdZcJCCniEAGvr6N2DfxSTvJ0g+bAQPO4JLf/G7l
vYQYPIgO4DvdmGHT0TsBPABXUmRmZpKEOnNzZjH/kjBFyPhB3QXdz4uKD0w9cEbv
WY4wTeRpAW3NoKYgBy4W1K9pHIN5fS0DquUhj9JbmJjucTBWe2zdML+uNCMNRPvv
zI7rjtdvF28hEUpjWJQNR5OH8X7mCrbxHSQxPFLixwmit0e9hi8E9C9fdhPcRb7L
bwt2jFqlBM2K1sHLTcvldaPRYa2u3aFDR0XZGKjDQWD6EZuddrRSOTDgmJUQ+jhu
c2MSlyFxD4PBHvO1PTBADYD+hNskLVPzmc6v7AQglquOw4ouUIRzwxaWHNIZilaa
40kbP9LhalbW1bz7BquO4TvX1jYa/zmuP2YY9PY0vu7f9kxxO5OmvAfLkoiK8N74
L7LsdRIkwo9E+TnnfoF1crM8RROJWVJpz1dK1Sho/7SLiEJcDNc3RAWNspcq5aYG
dO9FrPeaQXDPwO8gJGfXArCWVwpWQEM5A1tMNJ1u79TzCe9PG3b1M0FC2JiaPn3Z
yPn8xSz+vxn74Ji8cSaat+Ef4jzV0tgtZygqH/TATXQ+tRJ0qLmBfgVYXjCwm9/7
vXXWrQeFpS7ynFFkW1dNfuxXOPFe1tU1Qv3ouw9zD/VUBXOOWcv35Y/PTNQBR398
O4s0Ym/fkmdc8zT/6RDH9X0bDF9hW6p0JOuwCNKnu3HBD/Nu+AoqlDnBSzUSRick
YbNOYZ9IHKMxgA7831qn+GuYHWm7Qe+aES7bKP5yIJIHqGNgGWyGEiwmmapf9g4x
JSszs2YzSxnuYZwPPl2X9lb7G9zUl3FNk0Yk+fE9RrNMuibLitCFxm5zoqTUuxyn
NYIvV0sswW6Bs+TidDmojxGRbUOpZoR3ZFZJ+3OuUF016poBebXB83w3GEPoVheM
LjVJzzoYDuta5ZzxK+VtslVAXo7i+sC9vrGFEDm1xpfn9JGcrTm9FO7pElzPk3vM
Gt8frmQQQTzmZ9I3XCqw5HgfkTwif1KR+tGe0jsSDgz9nMe6ISJICAvQSoOU2i9p
kHNu7Ti6tA/ZwTIEaV+XJJqf4lnZ2ZUzTcLZwBKGxY+6spL0Tf6iI/hkzT2x1ZOb
jWV99QYWrlRb6BCtjbfRJdRbGLT+I1tKBt2MUiPcWEFFRqataeQ+vjbIwBZ/xOvm
+V7Jl9FNcCaa/zIkOuYde7xWfRQTxAntiNpw/Z1+zr5sgZ1izm9DvNSGHikO+lcz
4+siu8tfcHF5ztG+ASU0cIi+OxXY39OQwg8cuT5/5eZ/ruawy5ZHWctOIaBJwWJC
6+AWn6z+yM1oHeowhhOvKqUIsSTzKXe0JUP5v0fspepcJpwsF/7CpHTw0FM5oGjM
ifANWnN8r55kXjz8HIVX7hdC54BBuzmfEf1rym5ucxh9XXUQMP8DNx42hjtltJJr
HxNzWbYo2Pd/p3DTxXZVjH0litfkIGlI7uX9ytJ6Ezrlj3CyX1E1aXUZQQN/ceqJ
7WNOYTxSMbakvACys5ll164SN2LfmWhPF37fIQisiYYvgXR5OBbvaA4MnsEbvQdZ
Ly5HdTk/wSy450jIJQfvReNig9rTdR3LBZACh04zGkUapxLancIN/+P+ZpMe28X8
CZjP8or9YF20vxTfCZZu0f7w99aFalGg2ULaBmvpWA+2n9j9xo8pKIN9tT8aeyV0
raXfl1Kdjh8B1E7NUytQQohsiTROHREDzF2b3DBPXAD1I6bflHR4zDSu3ntH6je2
8hctWhMI4q6161MsdbRlNgqIpWxKE44O8V9IZzl6u0zikGOL7HCLi14KIo39/NK8
H87Ks2ZxzAnlkvX14N1D/jLdy1IKcBsQ9c2N0w3BWbqd6SApMG67N4nn2GS7dQb+
WlsOVh0MGkGmFj+9M3xmQhYjocFJWm9KXyE0ZjC/UaBY6yCjTt874I8pezOActXY
vwIhMUpFRtCAtCXmgHLl25SDXHRye2qBWLHyZdbbLHg4Q5g6SB91mSf7OnxMETRg
Ju5H3GG1sE48gwXbN1UeL9IXk2R1RB/UoopXFoKiOfbCPeMfrYW3ucArVSjHbCSZ
QHZ2aEz3F5zYp2q9lKvzdBHnSoCqHCHLQW2AV0zPJ2vbQkU0tq4CJ55em95v2UlC
IQVuW+RfeP5ywzSBS1HeAhLgPrJkVtXsK3WlUXhAGVXqWeAN8YtNLAg/vbyP1Xbj
3lty/omj4B0j73EzJB/nK0XoQWUYRbvjAT4N56q0Z9+uMmMPCuQS5Kpt6s1kQRP3
pma9iEw/LbuDoFBntrEqdr5Cl8N4qppkj30nABkWoIq6H8x5iOPV+ewzCWKz1vNR
5xUEHPOzy+w3AiQAKOReO2DNfi+WS9Ecf+peKpbAmYjXIRmt+cC+LpxI/Uj+gIj2
Z1PyAwOfFSa8fibmev5aeyUerIAgY1Off/IFKh0Jv/h/HzNCVEnFLBRcxJA+3kTv
ZyzZhB8VMHFiD7GiKOqlbX17L+zimXdnp5FKJKYn2j9NtiLOYzLFK3PIX7wkMITC
baaVSV2N+JyR5MiZythnvJusWhdODQyKu/yLeovRVYZFtv2biTwWSYTVbQiKcUfP
7444FawxJSi90oPtxNe/bX9o2o+n/dctObL/1MUt9CEki7T+JdfEQzeg87JxDbZL
/tADD9HW1iCESelRiGikdZYUl8RjtyALpqiFVE3zOD16bDEAkZEjCgwyx53pP9B0
fIVKlMds/GDQc1GDQQYV9DHUtrhaIitHyxYxiW7hrHOj3bqttUOXyVZU6KOmj/T4
MPJbF5tOsB5L4Iy3gtzagWbYzld1Wgvo5I38syI1Kz2FmIiOk+F+Azt9OZwAWaI2
siBBaQBJ09xT3lALVGHQui/C8JInunAGAEAICaLxCMQv6bpI0XwefbJSJfwbhCUs
ThZxxx6aHLnv8XbEAqJ6GwLas/W97It9O5BGmOFOYwSlW28AGp2GyWkCf9Ua19pV
4KK7WHzIa03dYxfPS9q/0EZjvYN0mo2LR4APSf55uFuaJJfiw+DLj8qEwhQ971E+
L/BeWRKXM2BcvKwoBC3XMFYPAl/SsANwiGBtGXKdxUzmy3lxDocdnDLjXiUNAnvB
GQ6/tT5zm0G2gEykMhSfRVBVS40nS9+WhBbAFK4vKq92sNl+xVWZwTyVU8vnUb4S
G/JyXqHHgvkI7nRM50O+nlhlu1WxlAfU+SyMtg74ZyMbMMGNAZRFauUXPdpbgrbY
uBmK4WTG/4mAO27mTKA+ets9gyVThuNyTL9gsDVmXIh86D6JN2/mKfyditTCyMcE
dc9Gnf7XQfzMHlS2z+ni56GLJIW8ru8tywZI9v7vryEWFI4DJjYsNKDmxcPPje8w
+oNxBCDawE0D4VXJGJ6zSs03NUk+tDooXYk2qlJxQjV+DWe4kVwE54sugN2y9q8K
Uq5nWTDZODc/g+Nn0Mvm9v9yHA986KDPifCMyXygOU+34ZQZdlhobW2uC75gNY2z
4Y9meWhysZHZQVWI+JoGvwBrMI7LFUxnNNrB9+7hfX08Cu65tUnvYS7dlz31T+oF
2z/iIiPOxO6fdEfzkIJdyj6mdTcYy66ZoCnYjnNIms2t2u/VVd1lSwb0FzOIRPHy
52+NNkiCj+41SAOZE7utu7JlaFrjn7/BDUBkV6iysrZ4N0Dtddt0DxjFdNL89mbd
BHuUykYRt8PWjbESKq88q6LI0jWfdRLhFV+ASMTEsfPt+Gd1c5OdLxv8ZCcImnsF
/ASKYApJYtj/nIdrwzxmEaYmnQy8D5ZjydmVy0RUVuIjoL2k0u5GHfCpE7wxGi/X
N6J57DKHeYUl4T/4FOIJa1DwQsSQuzOfgry2QRMZE6w7IabbWlYBsv2rCmN9TCbW
6Op4XIhpNgQAyFL/ldr8S2i3YZIjXyyYhKQGt4WVq4DZHfNd9pX5sRP4+A/k2uS2
FN3eSiETniAw5csrOk9QIYt9wjb3bsoQd4xoOEecVXRi06HPnpm82fmPsxfZjsCz
MoR5G2d0ZyQhgxLpgU3f6y8HTyH9heQZFpmSKgnI2XqJsWxf4GfeH1FR0DewSWxa
gS73O5zFwmfR7NcxQgiifAW05/bo1RFv/pXPP3Mmzgb34JTz8IAixgyl3eueHtZQ
JBMkBLpuSZnT3ns31HdAcHc5W17ILDKWXsOGHu1+t3HfU1fc2WQttxhxs5bRdVHy
n4Vex+mObw4Hh6c8Ja6wuz/gzfWzglBKvQnjnpHqPHf6Q3Uzgm4NjZ+jFc4XRiWF
Z/pxA6RxUyU/di+CPpI7ujNfngdbLiLk30+HXlLXidI2aSRgW8wHfuEQ6cK3MIO+
2XTHQACV1hcwZqnZuFyliNJHIHZDvemFnJoboBTmJiaaBkmcroRtKNIuW2Epo0H4
GMOQV0ciqi6Sc/duzqpPdN5YI8j8dcC7IgE8R8wJ6hxnM6t3EJToZaOkB5CKxtI5
cfxHd7IyCozJgyZD8mAoyP/0gz3czuiuqRSB/Mt5pAOhJv4XryN3iqQ4ieiCSgqp
KtjH8hh0QNbSXCJeRB72UhqQLE5nTeTpNBBpSO6flmM6ukVbhG00AmXRAXpbHtam
qGtoZdFi3sYXC3ogEv3nma9ML/+dF21uVfUx5ypCh6PKq2OSYQ9Jd2XBg+9Gu+0L
s52i+IVcsumm9DwWWHlrVuD/ixl+XYYZ2jfkNdMtDdA1ZMZahR1z1fpWg7YuW5Ac
fjKAeOifioFvIFMO3TtMMtLxE4ij0pUWIxqyfLh7f03ShFUatgbQosB9pexIQj+/
35b9mRlKLbS/45BZ5LHUb0LMWwagBtLgJtgTqx4NgwlmcjQmiolhE8+aJCgl0L8C
fH56YImI2lPWfblYGl0jHGFsHFtL0St0SSDodA1Lu651Iq7FUiyAQobIijM/kgkJ
ok+wXB/jKXv8JJ7dmF0DkcO4z3jhBWSftIlmUkmuPJLygqA4rQWusYZC0Jkv4qgr
eID9Wi5caD1whX4xKyQg47dsH+C3jBj5ZElRm+wrRwYVK9V4xYq1wVQZ2RVbWSeg
fwFcKjq/0BjWN6ruvTkMEOAQno+2neXyNnW+XabBiszYd/Al9rVFpt5BdBLWnsij
hwiPfDDkFrhfaIBz1hZlAHKcpg/HQzDL8x9UJFmk7WmrfDlhMa2zB86JDnSroToE
HBMLR6MZMMV/yxNXGbh7fkPxgZyHCRvGdN1Q7AlOmWRD1SkX80la8+S4xUrU3Usf
KKHspTIJVlJJ0utjHeSiHn6caBCCnsDnEJ7twrCcCD63MQraiWgEKgSCok/JZjy9
Kd7Po+2qV0tEk6rF0A/Fvu1UI0ohDC51K0go08xPJ5jPuKx0YVTBQoZeRwnf+bJv
oYSD6FCscFiCeAH1Z50UTgSx2ZMXWGgfrPFSdcgp3/gfpmui0FwQbc0rqcy4dFLK
PGXCnER8Dh0wHtcHXobizyIHjJutXXVe4xoRtjuSqFGbQScbBJLOz+tmiPlULiRl
AD+yW7LO64t00bHY/gkV4eBwAHGisr+3r2blyNwGscf95w7UU18DWxX2aKRpi9Cz
ps+Lb+bHQqL5K8PDFHWaNmif/yOuk62DLiTZTqGdDjh2JcpOvhxQ047/L+5ljEsh
DhFk7w8jdZBKl+VfBVmhoF1uUPU1EF5GZhGMeKDJFG3jm7jPdXnp4lv2jlp2qLTZ
Yfr8XyWHPzUNwvBv4keX6dX3JIxzCB3hSKALxsZMGn1dfuYZZMJScaWH18VtT3ey
SUVtcJpvfQqkaWDoZU+vw9Sna0DCADjgPLI0Uc7b3rGcwsjQqetvfSSrB2AZRQiB
6mDK1PtqUOeVE57dwU2ZomY9v6j3FI8B1JHhq0tUsZ77P8+eZTQOLgxVZrdqm8xz
v9uRXDfW/ZeNux/oJpFsRUeOlcLHLiCPzh9V405ENHr92zGu8JDzV2O0uW+FQeoG
qpPBem2ptQpkRM6G8WQ53gleFfcAAmJdlwlxaRBtyFTw6S+EK1D3TuQWyB0LDrNK
xnLosL8QlJDVyQ2dmZqNJcFb1O1Q2eA5tEc5/x8+1X3ndh9WLv1F+yxLgPb0sHSH
iPhXv0xpjubpVALhaSAYbMDcK30aFZr/6vodHxONk9oNFnd+6lpab7LXiGe5PWIC
eYLPqBuTuWvYmZL3jKN22E5YYwfz2IYHX4sIZbbtUvM8QVKGuZhNO94Y77QcUePv
AanRM/QyyPQ5wN32nAFpF9NTxNVhnMw4FBHPDCsjyQERpAgw4RP8hshr2Yp4RdB5
7hJZCOQQywYOXX8AVvhJ8QlZL1gStonFqe6vc92dKU1lc+FBmTYz0nGjc6G9/E0f
DRbHsHLtGcSyQPntRwxqRlXfjwnQj0d/MoEiXCvh2VYoQR5jO9n2N8P9LOdrXwx9
QFERV+Ga4HWNmvQGDtvvZh0aCZPrBeDAFhl0rnL8i4joNDjaAx/WkEzfG4jgLV8C
rQvSASuxhOO60Wo5SJq8KwO/bMuUTTNsUlGgcKdvKG14U3ZeAmo6RQN5M2sVnVvn
PKFhFyOhL84gPGjlpyyIvr9ym63GNg/1VbieavvjkxmyE5exgDQMFgk70rKNriO+
eUUzxhx9daYl3ekzD3+L3nEYqX+DUa6iJuVQC4gIAVXAhF+k1XxLEa2xy4wLFZvO
I3pl5EPazEBIA8F3gU1UyB47GXf91OKBgXao2kpEdXRPFZ9t4XowqLnrvoqtskVW
8nSq7qJvnmJHiBdWbUjBFbYcQ2atZLFW/VUVVb51QUNA1+bylXPP0PjBbrzeAm8h
5gvUIBJFR2mpWPih4C2y6kGFyyA4FT/isj/4UGNRSKILbUYL4c9EZsn5BNoCQR3J
ouDCGc1RShYubkf+qruixNYGJYPuUViowVcPeRzjfLYhhWOWd5XFfBsxbwPfJ6nf
UBPtQAcCNCTBVrE+n/7k1tIS6ti18Q9tV5hALLfFttUYPDWSpzDq+do/9+Q2TVhI
Tu+10db7fWM5TdXMR3O5iijKl8cZj/1UaODvmL6Ot0XImY6QEkcqxabczjI4JuBg
4BilrX/JXyLMB/VHNMdlfnLbwxqrU0QLa9eCkHmb/WKGcoKmIWb7qdLleb7UbNba
NgKM6+He6M2Xqonw4+GUiBGTDWdGXbXWzSrTKB4wSO6x2MPcZFxAj3jmH00WLTVC
NwCQjJPQSwn4ejUUWDdIn5aaSDmjw8gBVUiX/r3gnm3g+nMuOk2HpI7oFLP2A8kn
i/tjwxcgRO/J7nW4od0hhrer1rbWECtMG7zqkVTzrb56rIBf9e/FmGUpZn1WCi6O
S01sNBlDhUrInIp7ciIiepfmdsQSUBOLjYR9C6kG7E3x6w9LFZSPuHeLPsR2Knul
aCRMvn6LQR+nIQObiJyj1yqa6/mBzwjEhB5Gn7a6JFAS96kvDWX0MGPn6ajveoo7
ysI6sCk59dRXjZrxshbIG8gavjq0Wf7vFEDw3LZ5FU78sFylAniEl99gpjPh+uQj
JLnH994DJuv3UI0Oh6n897NgpJImaHwaL9UrJn5Lw2sy/8JXt6VX/reG7p3j/+7B
hk/SNkNMe6qjNKFJkR7WmbaFijuz8L4uzUYd6DwVjXDh11r1Wws0I0RDk7dV8XR5
Gnms7av0GmYqVYMkM+W1V/9ez0KcMSuaNYAvgQdI20QJ1gMKHiLhOy53aEzm/QR7
rla7PVCPpvWfiOkWmkxD6ROTv4a+JLbkd+YTGLX/hND8t0pFEClq71Hqr4QUQUDz
YD8ar91z7uEMYWqoGD6+6mIYH0nVWn2iJuF9svH0Jutd0i8ca2+98dUQnTu6TA0I
NTYNr6XtGdThxQjBOdU/kULA6RuQLDa8/8mq0eTGXuP2osUPpQq+pOdBQZQ83Qzo
akx25aM/Clk5fjXv7eKg7MkkjjMqjjpqDGSHSYOSajPdkMzBDhLDC3AZTwqrwaeh
ROSEuzx9u2Ea8o9CZXEM2O0eNFkv33uPzdG3vHa5YkZLplapCB839I4zQuA7BAsb
9yWVrL3TjYXkg/+8lXObmIMfJe0x8xRdKDRnlws9QnQmXTKw9G7BFeexoq6J8JoZ
HErVh6PmDMUdh7e5CkPuPyfxMmnk+P0F+smlv5BaEPe/lCnqY+bszE3uAzsTyIaZ
vTEcmZ7TYZCda7BHZ/oYKMEUZiWTQ5pGqfgaF0rZt0eG/NAMscAnhhfJQ+xj4sh2
nKkiBBtcvABLR7+/3s9sWq+5rg9fS9jc+vD8+t7coQodpSp4eH/M61LpUCD6TlLU
g8+HnkL3QNtjD13pQ9osEr3i1cfFc5CG1tKvbvnT8WXTJ0N772vRIqcj+ziXFpRU
758cI/S7rozMuPxvrvbxzVpfjQ6ZpIfCoKbQPMSK5etrySZi/+SKvu0VndBjeUv7
nc5kI+5B65dveXgjg3DtERh6VRD4ys4pOf7nUSQEOCBqdljq6uuzKt/ZGJDtXPOr
ZQ1ZBIwWvGj7LCmLtTOw5FTCASPDqpWPzh9xAQ65UiEMRmz9f+P+anAWSMrMzPI4
miAfvQEQchTm1eKPJ6M5fB48Ppb+cSqlCSN9nSFKs9/l7pcdF5JAsl+8jwLeXcs7
IHZK9/EfePn/Y0Od56ny52AV6eymNNVr8L1jaUDcXXfYQ86TgX4z7f/Jl32VVRnO
Vp9kVyZWQW5SR9UruAnKbNbCdDte9FkRVaV/KZUWaiYVW9baTfADn3H+8ff2RGID
ZrHkqntQEY1s0bXdKaCnehM8Zl/V+zKvwqnVc7ROZmujDnRdIVdWvReJ5Jz3+iOJ
WGOCdKn4tMMkzrPV9npn/iXX4rRoKE/dscFvC/91RhQqQ4Cr/AkFMPrthSO3232L
A3jyR5Vu+Jb7Lz27MlPdxDfCIwsGV1/eLnP9fh1eFT1ogMxZjVxuNHEbGLpBRK74
R3dgnkvXDbppAV5iDZNCf3ea/Fg03SXG3mmVHD6JUGD1zGRRCkmEUrbZSPE1Kq4c
B7SGOMoCWAEDVg8b7Z6ZNHedc4ZBebqKsv5brX088iCKCoh6fCAhMVNxDd5QBh3z
ryNwC1essGJOGjQpjpmVXSjaKx3yoEZj1JH4Bp48cgZ+jALoG3/sY9jUFqjp3Vg8
6/vbKETMMMjW2O2ogy00mFvLaicUJf/hJYfAswmhA+lqM7lBdGUYpSVjj4PAW47R
pOHf5KOHm2Rf/5oKTfe05UY48XvlyeB3gOdGO60cOLnN0WU2ZY8BBBiPoWtWS2cN
1c26C3emHL4d+PloxSnonshEyRroflpH+VP/DARGbXMLemP7vMxg6zRyoQ2FoYpS
Q5O4OvxhPve+6DoA8ByKXnHsgK+HpfIyOm0wO9YjBNeJUJwF81zCszp+cb9Epx6g
eXJ4KNV4rnbktOZdfRJpDTIUeZXVY6ZrTtCKjcc/8YfO2ZxBlOS5xw+2LbfLo/Zt
whsAal2pkVPKY4twFETSlXOPLAV4zRyd7mLQVFMw2WkVlHKvLuEfQ4V5S0y7ihZE
IQkZDbNW2BM179c663VJD/X5HHTA92LRfzUyuP3/uvo7V8gmiF/jrdoAszWRuGNa
dDJhzek13TnlNM+nUQgAXVpXxGOZlu7ML5huAMI+HIHrrdCHofnt2ANn1B1DI99a
9HE9R4eJBuiNdrKKwZf5RFXXmEiXibTTt5ApHpj761CZYlsrl5mHnmxidMGp46bn
rm2YA9icQaBUooUxbSYudpfM4iXGkydQqaEv033R7xu870Sv/skc+TlW7Z7giVFm
v4eyx5bsgFCjevm+zBOgo5WCXAcg4wD9L5v6YFLJOeCFYo+ZePaHCr9ex9sbx3rW
uSL7Mif4dRP8w5jfUs45JOnKcCrFWP8B/9bP/x4VMrZlFDtnUSIZUk1dNksreass
W8n0ECWjPg5MzDVQE/KSYwy9Zv9Clwt43G0JjrzRvqzKw7GJvpKvhUg+9KOdQbkb
gt8++9geJmVYuvq53mMWPBQIhS0HZIoC8dYm3lArUjDewjMaIlTkun0xHZPR/566
PyTCGlEZ2TbNrlANCB55gkTGohap7L35dSjfkJZRkXFHpbmQSnv9RfPD8jGPLDAi
WDVVIpQhz0qKfSiax4JOWBGQ0knnQ/vJzAE3QHZj9XBYDgbCvZiJwc2miJLu713n
NAiiqqI08GFpH+Iv1JcThvgVYAMml+DfpJ2c9XIPl0Ba5xhh00GH1/Eqxq05Z0f4
mle3qABIXOao21fU1h/g33fxIYlfA3utWCWeIHMydzVZlwR6AWWcbmUa54Vg+UHs
l+JIacVQprIJd581c3tMEUcCiyIILz3OkRHIjxsp4zhoN1V7gSEGh9goFIN2y7++
S2BzFYT0zeKM8Ht4RCYBMQv9JVBfNpcqo6wmPYmtZpzgwSESb/GxdDipMt7zoqmB
eGM5IeSBos/4RR2ypjwC2XrV11ilTIflymQIvCQvyn/TqWveTteBH9qrlp0isM0d
Uhda6045ufs+bccDNup0Z3vSsE0cf7Bm7ngIPdm0RRiN3JK3eteeoqwBVewbOduM
+M6mNI6UQGFNTWAQ/HWDq8KE7QKR78XedXzyInGUSMrt0tRsfNKDTbtYngbrgHOS
THDeuDthwR8Kry6EZWMWA9qVA4eI7EiooQCpdpTRfQXqK+7W/CsKKV5gAgP24ir/
cfTPN6SV1sHrWJIUWr405ZpLbkvMmZlZFhlzKtt0LCqwEbpy3vx1lfCbnSGKdTZg
L+vUDqizDkyjUdzwYk7W8gwuKJcvbieFAmZJaHXkiiRV1etjYAnuRYPz1f7NjaN4
LD67vsi2K6zgfhCCcmlUy98mdACDg65BG+1AGc2uQXX6xTe254XSiapUQB73E5y2
eZlNnQJTBjajB82LFcISmBPnYYYeQNhNSNPj37mfgk0jEAcB3Eg5ORK6N99gtmmX
+gx+yl3K6Uqe75X16qJd1Ln7/Dzea7jUDMfG74SvOffbZI586B+6Q0UgjgljIojN
hdapO8j5gbVlVpHF9cI5iuaDb51UrSZ1zkDOx7VqCl/wsc0IIQRMYnxaxEZ1KT3k
81133gOSzDqBLzNchXA2KhGqSbx028mzM+Dg6aPThElmD14uhG8mweaSS4pgXXik
UobuTEn7XRSkVG2uJSIeleD45Hl90L0JgkQutLlZWmv7Bc2T6sc9nuVslVkgYUZl
Nkcl/ESWVQrbYN2bQM5yrBVkDiPkYHdVJBHHRMfy9PA0UIZQ83s5gNZi0/44GDCA
A7i15QgvzgKETnSqsW7SFzyfc505Dcfm/Sz0jFgQU244vm0lkgIkLiRxy0ZEgt5j
umnCxTXcbgUiOx6V1O3uZ9El/VYVm2Bt3Pz9HbQi79CXQ6QuvrvB8gZjmYNxKjno
X0bgFw+TOfqvQhCVJpz44E7QNy/udxuUpc3Jk+dTVxKW6gHh34aOf37sdkSmqLLs
p0rVasaFqL6+V50vid9B5Bvune9LhF4PqfUnONAbEm5bBsKCGA63WpWMA6dGeRJ8
w6tfi1tX405ZZqh+jSEMz2ZLzEXEWhhInml8RoqRvxESyHKjc0T+UkS8fDtGCg3U
xby9hl0HZ3ew2dpG0JjQMTfYFYZERWOcKkGK8nikd+jlZrqJVdjOShv7IB7Ubx3L
czrcpzhlOzRoTw1xECGY/Po9WYh238AIml6hWqy/sV7M+U69tnKwjJNv06I7VC0T
bp7KF61LoLny7Xl6N5rv5fQDt/d/zfXzknPA+O/YXJI3y5rog4XYgayRcDNfabcI
vkYt5cwBjfjv/raQqui3PxmqXcjACJGVoNPLXmrBi59RviANe4uoh2x9sgiMn88O
VqbSlZjwoDfLrIQw5CvRc46MtZw63lz9cmZHDmf9Nkn22ILI2u9ZKYAeI1Y62IAw
lGold05cqQpiHmomql3lS6Cp7sePRl6kMkkmqtKf7UFpZLuz58JIFZoUmVikF6NQ
vBk0QSKmBsACoDOtxxkxjP1CtP3N1flDurVdn6zifn3RU3VAC11eYSGpwTiNghSm
FkgHFBIwnrWDnwducdUz17S+F/Mo5hyQsTGRODPmDA2LAgzFPZTAMnpEpVKIUMpb
xiLsKy9IR4d8TlviU6NPEC9fxOVX/7UkdF0xWs93+QSzFB9vXb5Gspx9BVhgzORx
jgvc6LCQZ4M3Azi9X7YiFroZ9smzZjzMMwNNHMB0c62u/JmxOtHPugXz3HtCRaVU
7byNhra66Lw/IFxWxj89uXBuxwqGcpnMVCaNuQ/niiOnsVVWEmJ3Yc4iX++3IbGo
ccOfO1SPO9rjxrHv6t1WDLskxCdeT8t+h5tD+z4jcRzbW6mtBW1Qwyzb1Zr9yj+A
M3vCK1OSnVXkyadOfdevV+/n/Zj1mJZYpQJE5scKTuGzRqhCIP2OVIPA1jrrTJKn
wV+0zeITXW6y49HSfmw7iLKA0kUV6Cc/Sh20YviXULklSbVEMn3kuWP0P0iIp7+p
5S430o7gJ1ZS6wzb4PqUwqmTSpKEyxRh6IKQeJt7duvCeDoqWDuzzxns0jQfMMSW
S2oAn91qRUky7sP74kCUSr0K2GBTy3IMTHsTcksEVaToTNdKjsfOJNKKfvkwaxTq
Z5D1lzXcQoEKrTJispFzFDzOCzc1/Qbc3UI/5sq92EmpGbyw6ZDrbRVUYUHIHyVs
sPIDLPj5g2UX9vLtoF+pakQRkKXrFjJIttZRuQoU4WlUkxQkn7wiV2lg1jzJbwRY
tBOpQJSd/c6DCjDAJSNDYzEzuJMWjBCfmI8JXq2/h76P4iddIYvAKj2vLZDOVZih
J0BOO5xbekOLFTo0tJ217+azQRW0/Bi7gJPMhnzYdVigRtsiN0vmLNG5yPqXHtE3
AHaWp3AHNm3NzMqJ/ry5SC3Do1ROczBrRHas+hNOZGibaYPqy10+rkzGtLWYeXlG
PhrNSrIoYs4mFMxDpfhYe3BcuNU6XS8hTPt59XvAlzwjAfYVEdziGcwceP57eZCP
scZPwe3uvdDIqYU5una+7jfRhBf/z9obz0FMZTbURnhJIY072QxRXUqmjnHOQoK5
ShfBdvNy54tJv9CVslH+cnxOFHAUGPWXIgYYc2LuHtrh7lpU7IP5faniKigQsvAq
uBKiTp3S7F1X+NTUUO+7UuO/kCJQhayt+U01U/azQGJdAKx/Wpwm4ZaBByBVYyvf
556NMhIaRXDjImypCpnzPlqFoLGLtjgFT4jjHqwfNqAre1PIuZVhVbbLV34Nb7v8
BH+TgjTPQUx8jY0IPqdghj8hth0eNsRPziDc7wdTxNLrHf5eBRHvamguBPMdEBHU
qw5Dv1NyRVLdQ/EzVBL1eJdXePPiJ2K/jP/3bZCeJ3fFG2A78Lo6AfUbVRiw99wo
YjtRHQ3JrKf3rqWUB2sSG7lbaLb9Cxou4UZbqItZbRC58mpj+tBBMr25P3MpAhO7
G94hYtO+srzHvNgAPQ2g8b0gUULHCL21eVA9R+pAYFUkH3/BmafJm27du+N6NrMv
08OP6G4DhdFSK7m3P6s3ZryVbpdULADi1eHtxGskvQg+QJDg2i1t9ZAbhu5zuMCu
41hFOXyNxuMIVEG26UjUZKYJHOaa54gyrE3xZR9JTqESD8akRNJMAeZ2aE+U4Gzr
a33DjMbTaaonQg0gcjVR9NLecosIPNXHD12HLV4upSBX6Xz6DchTtaQ/WhdehV3m
L4Mfe/aT3Na9JGuaTV9JCdQGpZ4NUurYxwwYvHi42fjKpN59/boy7BvKee8nPjx9
sZZPIFi7fpFe8iguu3pBdDjjE43LDh32MFxPpgX31EduCQKbZ2uLeYit2Js+rtiN
zhQEsRSC5eDyeDoWDrTx702f+R4MBUK/k7VL/1HoczpmR/RCr38fxEldDn3reAQt
RjdXjcbvWKmkSJElvtiDCIMaTyonzsNswB+UjccdN8nNceCAkYwm7DR8AgijWtfv
j6trSPG4jeWVBzL4fUrEi5tb0hphIx66bch45gJK17FFLXC7sFBu+XCESyr0Yag3
RSQHiNIzG7DdJ1B7uPUUH/VOyireyXSc5VNtBa7PEaHx2P8XXT+gaaOwA4CArKEf
plqnD3YbMgt9DPo9Q1BgxKKPkWai1153Gatvl3ZkpZsNEJj4HpjsYt3ZMvp5kMwL
VEIrVXkJNHlVMUHM09Ty7ITtKfkAXK+WLwkUbnVhyXFE67IAkc1qHC7tCIhs/Su8
Ag5dXQLA/PiKIJ1kcB/DayEPkJocr+Nz8a3Bc4jNsdsYlFsNrChvFos01SEFeCh6
GcHMdvy10S62wyicOndqZ9fVTKtXplp3ZMai+4ww0/6rOH4vrVrQJyClOP7guiT6
85PwmZf7g35xJehdVrkgUBmtIGd9b3JSsRo6V9tst0FqMAO07k+HBL5TE6oYDleM
i9g4pqvQ2rHgFIjpd+S+yQhR4vgTR84MMQsx+2bpNYe4+qbNVwEiRcMSmAyS4kFi
eq3Kp0WmLS7hkg2z7HaXA+LBSb34+C+OUWVJHqKE8sJMoSI/MzYd5FrsYPJw42u3
X13ThZ645WPbUpowTzdy9mIJH583ZIsogqq+aQBtBXlje0I52zhLoUsrx7XUTKPR
82ax4Czcrad3W+R83x0dh2o33EPzsRDCURWm3pqtoBMJJG1yH9wF0vYBx8ljPbiQ
aiXxlVfQ9xgzc3MY+7whmeoFj+hQ5wYS5cEFJY8iI6ONaJ0PqSYbDsHsNwnFdANy
ER7UFth8N9qHIOLoMS2Y9IrNIL5CKJiMlBanzmNlhJZn8KaEsakX3oZ7RJoZ9uXJ
ayD7UPFD+vWHJO3f4Z6h+5i7Gj4jgOZifTuaDanr+eP5qGUSM+2uo8EOz0GmvEpr
1dAWH0Kw2n0zD65GDfZQFprSr1rVFgExkexyHdjEJI2cuHxm/pG/2bFscNOvuNcG
lNO3e4g5d7ta6wYXPKEQsGehSaMNSDYycTKWSL0KUSahO5+T378xWCjTtSJOFks5
Czisj6HQ299m7TmM1rb1u2JjDY3dMCaUXkIt5AmVlVhC1ssSSjoSDvhwhbjoSOEi
sFLs6vboHEKwObrgpTsEHn8QFzHG1arlHby3X6rQGvoBJtIksHaorVvVLqhkvSf4
2QsHgSmQfq6jQA4Tpj3vQUDOBKUtSmQFRmO+SECDNj4gzXbv6i23lK62fRtAvjvd
s4hhucvm2dBBMasT6GAdv7JG2fiOFzpAQyHW/AfH0dZijKs0pQI4QUIRnRdlwKQT
raG+/0JUhyoKwcseMk/jEt0K/dFd7ID1Uyki8zVV6I+2H8mSJvvbcitpuoKYnF5h
Vq1o4qFChuvyyELcc61HVnq0bCeFZ1b2AT7CsA9+vLka+FUDYCHrfXC6VPmbrecO
So9yksjqLpA/sZR5qRx+Bh5A96jC5PAa9ZznhMncnJ9kPkh2twIG+t4vuQx2y8qk
2VPCTbA0vvNRTwzDaD8lf5q+UHYIEZ2BBc2dUsPpqHJ4TUkkvNcAcZiwGUY9R5er
xbjD0NDk8aK01lG1U+tB3yyoKJGeIPpcsdfTwD1wD3UVOtDSTAIXrOzYMRns5+I4
W1Ez9oraG71lIxTEX1iomTgPxvc1IQ2cnOyZbA3orc8Y72lZj2Y+j2J3+XEDdAIC
vLbztU8xK9zoLodnYGgszWpEmuVAo1edyRJlEfSiXthPBsnaiRsi6ttQoqy33q0B
ejrW/VJSo47nR2YTCgJ2RMAn4zAOaWZQ6FXn/04j7//8g+YoVOtgbSyRjroKnSQ0
z9KFU9FstBC4qJi3lyrTJdMEZL2a/1uX/8OYhkVlqzkbrJEUNrj0AUXMUVWdpzl8
uo7lSQdWGJDEgN3RWp3wUp9ZfhV/knPtt5470s8YHciDK/N7u6DxryM3oO+WwQsW
2uhNctXZWGUB2i1iMdSZ61HFGWqoyNMW/K7za4EInuCq43f0tyFYHazjVrnruZq0
tU7u0uw8CzHXJB5ICLmOjW+uPJf4tvlirR6QEJO10WKgvNFmfCdNmb9wj7w4+9Bf
FfYblCOzfO8r+E5F9lBbPUX+YlGDT8N0YCnvJQINKoii4PK54fd03t1gVMsOtkXl
6yANM2E1+2iyCNLn9hBLGAohZwBSNDKK9R77aXQvgXB0Bd2j6LGZSlADFBmoMUgZ
vjsa7j2QKLCi7gRIWULaC69Wy/s7I81sSY6ZBJgJ80EcwQn9/CPMaV7yWHJLLDSU
P4qSrE8q31QA0zQ1tP0W+Hb9d1fTwP0zUXACiwWjPbKQg4uT9ulYucLLOZo9g1ld
x+/d6AGYihxOr9OlwTZ9ecujWWAN4zz5IB3jN+VlnRRUxRxOaQyqtiLmxy9jd1nW
EPdD8P5zFTyU2/RCvSLRTntq30KnOm40uzeh4wWfEm8S8RUMKp6KdLB7IzYNp0+2
hSlbrYexUAYhaUEwSm28WZNEoEQG+abSd2Efa/oTiqfiS9IoAJ8agJ/HNv1C6dk6
SfCST0nMI4IhyLIM1gJ7PSlOW2igWptNMMC1iXdr02GaXLvqJGlCRB7PdMivhLQ3
2LXbqCVk5dnepzQbdFE05RULiFU90HxPVjXteH+f7vdnX+npGGaRk+XFARBZr6/c
iH4dPACOJ/CyiplA20vTglQp7P8RkXy9sCirgAIiLHH9t4D04ViXkmhl9o29kXK+
Y+iKrgExAa9awDi+F8B+oMIXx99NQ3bpvwKI20aIJQs8hx2eQ/2LHv1XZ9WDw3NX
2phpbfEg2hFsuRFh6ZyPyPQJr73RvYS+OuHhgQ3CP95H4g7mJK8d6oA8jBZwp8o8
X8JLBDXGNZ9iIPzPjXelabBdszXTiwkwShNK2ePlgKbeq8oxkq4HeRLBpp7ain+5
s1GXzWr1e9er0Eg3BrC8f/2q9G2Zl1MApdNZW/Q7+1XU5u7mQ9KWpVYugbdmUXGs
j8P0qK560ewSpyEACo7Zs6I5x4xjIyfy2dwm0CjCSTxm9KYEkfETlFAUDWrxJhcu
rUECyr3FJseCQdAI2EDphNG/1yZbSfQGEA9L2o88iy/hZXD7HZT6oDD5BwEXGY73
ixLw/+nhmuVMysQ3Dr6IlLZRY0jSLBY3SX/FDuBn2z6WMjlPrM39czJ8E6qdU8+u
RHitXBdbidMANKzgdGsHfuZLt5t/xBbTQISnTLM5bvRia5RxeVtHmqMgHYh+GmE7
hHsxhOuDedypuH1pRNXV29gH/zNGUYC2lBqMduPVVBV7N0Rkdns+CmYx+wgN097f
Wo/i1WZCTXKaJP89J0+0qNL/15xtIH/5q1+eWGZvL/cBSe2oOfQzCQsN7kcicOcH
uyLcu4TzaBkZlTTbLynRBjjjVpvPp/zvA9SHG6NhQ/1i2ekuhoY/a0Ced3ahg1fV
AXv/pr8HBp4z7gP4XbhRcfgPrvBgVxgI/jxywDlaFBqw2jjwrEuL6T9jlxXB1Ga4
pUkEKrUfSAAZMf4n/rKW4d7XQF4ZoD5lzA4yH3waLpGBtEBQqUFDAFZiosVuAyB7
8oySi45EuZMSrweqFilxI3FLj9cmsKZXliDeLd99I0PRB3gqPQxmDhscDKzSO0Eh
/4KkYDlkvYDzTxQqXfEyaXs3TU1dht7+150wtf8DBtjTCmgvN/uCdkEcaa33Ukis
VPg0X1JU7QS/HhMtEzUxL+0MO9EzQUhjjxBo8QgsLa9MGy5GizdjuanxGWj6/HJM
ErXE4VEmMGsYwZT5SC+3G8Q5ICgjXn/mZg1zwwWYp5Ex1ANgP1BYjDb13pu69zRT
RgCatHgplyRtvjsKhk+FuZASuAUpdOUAKE15s2NYMiMEgjTUtASfoqJMhHEtFWjy
0mYZsbYRWflxWiB2kSw7n5TFLh5U21VJX2U3fz3kURLh1nKjo/KqjcOpLCMlpE5n
H7VWccWxMjlqPh82ihiIEA4CxvNxkCMzkCjyVW/XwyK6wdktazph0yVx+HBCluSB
DcjdnYSD5Ed1mXoA6I+8rB+YYY4ZYW+i1mI9P8UechOUry24y1prn7k6tteNWWrr
TDAIDC0C5NhKmymE3TVPqnmkkugKi/RI23FS8AvjZEvpy4MEpBJdN+0kiIRC5rXR
rrFEAIxnV7AFeFDiT3VHj66aVCrlU3sUWwkT1TeiSI86a/CWm7bC87/Ium8t8wr4
erSfBXvGLK9WNtVxE+mnHLEZluXzA0vA/i52DBTGfX2V6JbkzCNpDo2wVYYkBvK4
6jRnPH4CoCoZ6rdbXuL7H5ETlJC6IcexemLbrECJI2D6cSHGAOJiy57MnGNXOXFz
9Hec3zTNyXFGAqIgh0MnpKJ/i1yXwEcKzB2zv7tXUyNwN+RLM/yxlpIyUaK7eCQJ
mZDWlG9Fb8yFU88QGOCJjFrtoI8uGt4NHAuIf5law5ReSU9xTxqEo+MDMkVBfQr9
DsN6uGudrVXpkHNdcLzLURJB9mAr0704LUAvSYUd65dDRmPCZFortRs85t1Wq+xT
U9bb1OI+sDOwVLLulbucJ7lLgpmYTt8+MgYV6DfA0GAt/8AQUiQVdtw7qckSUL1x
651B7dJPshPr1K3mnPu+fswWa4KaqvK4q7iTj8BSQ6ggSwTP4eNC2/W4OlltVPvV
VoRZRkBtu3YfHsFy9N9+LlghCXX/U3JwWzeqvrMmKIFK+vlDh4cOGmVdeqEmNrcv
RVDdDGz1WtDAaSA9VKxHmFoe0FaqwtzKsjkI+DQR6pkUfTAwPb3UyOq/e+N40VK3
m6/yfUQ7yHYsVLFvsp4i6Qe9XHubXXbavdEci+l/29iF3Ts1T2bYDQkL2j8JC/+A
aXgMcpeQiS/ZzKx8vfwt8L+mlH+pHPxFv+7Mo9oGLLBBUIYo5OTwH0/l2V50IvPt
mpVFc6Snaj7RT/9yN3fT9KmeM0yus+jHNWNEepX6acOzEYPM0ybieYQiVpRSUtHg
fcYdJ8sS/kIyXu+1+Zq/1ipq5lxJ3/7tHRGRpQiW6nkJynDRWoGXtkr4hOIHND2k
uHZI9ylqA0WMHYYkGVRaGSoD9OUzHbVGY/jh71wDU4QUOuqACnHNYZM5hvwZsJUg
+XTX74e+HjucqK+nZYL7HXYihCQ2XiE/STAdyKSdhriW5XqVdU/NXWfpCiYgV236
dXCtTEK7TgqBgr8x5B06yUAj9QF68n31y3Upvllm6pKvFNFPlCqYsMKAhPcXdfqh
hQJtznqUjpZMYCwO7F2XHQ9xGV8x9gmWfdWPbFYCkVhpWv0jGKHIVTLc8IPrQlEt
3QbCklkQ2+4orIUJwX7txGx8UKzULiofL0mUUyLAl8trjm5JgczIUWi6IvuZesmO
PV5CDdTeDio+9wXiTCgmXW2lnVAorjOqMbjARyCfZ+qOOBLAJxWUm29qyn4T3neY
n6lVH18Lt2oCc/yM+CKqCRUiNXO93CRZUNHXM4BHCFKMJgPTK5bQCVR8D0D2MDFN
Yi09cWhPpX9/d/tXGLaQ7r01l2IhbTEw/UnAcFQ8rcGse5tkbQ69IbVSJ6KAJXNX
kfVb2xM/kN+bmEbBybjlZrV5rdVqjyJGag2nYgys8tJVoP9fTv0PF6lxjJIE6xtX
gGtr8RTuzLj7Tg4WyRdFW1aVK88zo1Wj2tAU3oF0bS2MlJY2ySuSSBAg5l2lOjG3
TX8crwz3CAwUcdcKhiM14/ty0sxHmiVKm2dRXKjUtyblyHw5mG/SuS9gW10sxK2y
TTsGrMd1MJLIVMqPKBp++BPr7DRuwr5JG49AyOUHxqMSTehhkyWCAQhLL47Wn55s
w4F8co6cm2oe6KbLHHasYOj/RupIp9auKAeUiM8f3lFEctHrc2esMLBoKXl6OCKr
XwNdN985tVPi1ZrZRPNleBvaBLI10XDJoV39NXVXxGezg2+k2EOT9s7eVma9DFt0
XriP8eTUmM1wVMUmgfjNQueKRqVmNtjJYE9cVse3th6lWTAJpyraC9b4hhnW7Xc9
WrFhMXY1qWyEs/uAgK7ZUoeoeHMl4Bkz5yB7mGo07eMscHS5wMyX9oJ7RO/qHndn
VXhQ8xw68X7myt4dy9FmV7Zzc8mH0gGbrBw1/N48t1P7RUt8OWLTKO7FiAq+jXq4
ig4vLagNMfRUIw1EgpML/gcq3JPD15FrDNlJr1sMAcAHB9ygCl580n3OqZjPmISs
8vbfn4v7u5a2L6leMXXATEaAbEtSvPYKdBCWnyJ27JkXMkJ/xnKgsoqPFtssP+9k
x7S0BoH62oB9Rw2Myzx5fb3yyJSDDnjZpRP6w5fRDkM4f72tHoEMG7uuds6vA/Gv
PKI4GzpFQKfpbvbuF9Xw7yc1zi7re2K8vkzWdTC+QEOkZkcPFo14YpddyH424twT
8XFY5Wgn7b4NlyHiBf2RkIlBAwhikrHmRzCnrvg43EERPWhBkA+DtvBQWbi4gG15
98nIf1jsiVHzKhUCvIdpYXl4DxFwnial75s8v53orobDUU0tXXATvg7+kWQi5SEj
JGxFWzgWl6z/c+885WmxSXT37/N2UruxibyhVhPDTqIdFhzJTjUGvmz0uZ1rXChJ
nE6XRFoPWTAGEskwGHsYVsrYThyxWiWq/xcPuTn6ViQWCg9P7fhwqpVQ8xtnNJpm
cIZ28H6RVK78LxN7qtUp1SCHxnkn1W3hU0IauHhZgJ3mvlbgdvMvXOltsUsg41l0
3fyroDiDi0s20nbN5IFp6D7ZN0t8BWXpg/es8jVhp4pGKWW3VHcA5ZxyI4N7CptL
0i1mWbvs1/r7d+w7Ze9ZOC1U2Xa2M1P+uMqgS4vnSukP9ooGcypZx5nZ8zK4rKSF
WdUXhAWF67eYofANEXY04DPCDSYS/4YgNJfdTPHanZ2Ks9l+vTL+EzFzKliJ4AMn
Bn1EVePi/omYHxXJfracikYYjTwPTC7eRz+jEBfbBKIxfpJssp1URYIfGyMpsPVp
jVsuEcHD60n+A5dMb61ytZVczCxb58jdrDIdppGJsNbBjp/VxnfeCymyNnnIkCIx
ZBbvsBdCrViKHC/AOpNAhQDuN7QrpKsphBrWYCT5dTmGZWaNtMGPunY9C0/9tNkd
3ogYkYKOvKum1p01/JmAbL2XSmDT4RzPscq5hBF202zQWrauRWvH2qPJApyXX6r/
/woLMD/zbCL4vPOO3dnpO6aSt8uFtxciYVv0k8aiA/QxV8kkn/M80/uwyM58uI3D
0l4UcCzujhDaWObSj0QfXbYRlaMb3AXvrdkJ6/cBR+BpK42NsCZm9GkOmoEEOx3/
eG0ilUPNOnj+0Yxacw8Vj6rWWk73ta6K/HcKfYc7LhCDXGY+MWaabCq6kymmHqC2
b5mqEsbyoO8+wJcNzdSY8TK6ZLuLpH5HKSrmUTSEkHnOchjoaElaKhWyVOqh7j0J
xClEJrMgTeV2/qvrUJSuO+RhVUDJN/CFrNZ+17Dh3NDTCiG8xGepJRAY7NAObN1B
wfoK8fE0IW030MiXLrsV7OAMrMP1hN8M2oKU66CLe3jyEOQlzYVNCLQJKm4ApEET
g0Y1tqXuNUqhdh5z/kUonu4UgVU6jxvPq+hYD9hccU1kMUvZca7ufCJKPTfHmPkE
DDfaxtYn0QsRwrMZ/ALBu5t8qXqr/jE52s9dRbGbkT3Evt0cYaLBjlaS83HxH6id
zI1rPViH0ZPCMCUAu5QKhV1jQLVZUeEIceUsLcIhEIV/kU0KTKrAhQ2TKxC4Cx1f
UpYh5/McgJC1hhHvfYtqZ5Y0BYX/pk+j0/hrl4+hIvlNSYP+CtpP+jyoB/jGoSJF
7VKyfc7PxwwnmfckkEF0lV/ZSKXlRkXhlvprOeFxOOQgpWZPm1wCShdWG//BFRUr
gXBSi1DyV1wRKcJBvayxst1kgI51EQnTPqo0cbs02+5RyanW3UrKbbFVpLvxSlez
FIiEMn/TQ8AuerUwmFbOt9WoJG0Erf8LVDKL5/YofUUvVH6GOEWUc8vyH3ffPsn+
nXStqNQpkUr6DACYXKeOGxz4nopHZ+9mG+UWr6xQ7dGR3afeGUvHH6XibHhsmqMy
vmOgzmYYKEiVH+HtIqpkYnIkCC+S2pwxKQdO1uhQoGIRYTUNh4z7ljaVO4DylWDa
gSggei4NItKV3e9FpAnGRtATkGw10bnWvyX36RTnk5ML/SRvjsgn123GTPoDlKFq
PU1mRC8jpqxB+DZBj6N46s8qH5lKi0TQclwq9Iuc5Y7YXqXuKQblifQQkyBEPN6F
SG63XkK9hoYBZ9IOfE21SV4WGw9N5xi3ugmsw8xBnYFhQEO2yNuYMk6ZDqkgMeoP
NTHrRjVEtUuvEa37SifmXUD+7iNSnGrGC/hzFCRc/jCFV8Mdnoh5dyB+qn366cGa
WEhKuAQiaI1umtsXSCnJWZxE2nIEjzM4Z71xfzAIS8ES7KAlb3dJ3juCyqM3MoC0
ymUMOqhUVNewkeLVYSzzxV6Q/kQcIXJeBZ6njyh/rhL5VBmoHXymC33z9KnI2bsE
UaMf21+sZSQ73blLE7Hi6KocblweHVqxS+ZZF+GzDh5l06AWN18vvdRMDR00A1Ki
9tVT56/kMvmW1XZQm0OD/bThARScDtzFXGMI8jl389wyG1+PjdrLGRZ0SYN0hfe3
cxnN1tNVxCv+kFRUBM91V4dER8sGaEFB4Nt+SWWCPVj1ZlJ0SGwUW/waCHr3QETF
1FyuddcWdud7aRAXfZ0yL8DDfpl6A0SFpCS19FFRdPXZbPCX86w9B9OjUrQNyP/4
I0RgVz3/kXH84yCAql01Upb2NazGxIV+wLR/FYVOib24KqMEsdq6Lv+SSJOu7wWj
bkT0bWhTQuSzIkcZwnlQ+H1nXWM25YSoK6pZeQ5HB0gQozD07HtcMY+JDdOBxYMP
Ap3vb9iH61UorbJTbNA2pQZLKBOOJ8b3aZluBeq7AhBDUzrOviqQtEpnoaBTw7+K
RzNWjbLKQcCyYKlXOduM9tXYwCmjAdFjh1Bnugvz8bshf1xkquNR/aMVth2WVydj
ufXq62opngdhefib8JxgAjDXLsgeWzhM0ma6MjaNVetVi+OS81QiAGZuEmjtaHbE
3QXi3dDkiYTA2wk9FTwJj2mLAr4TisvtzQ5oZoII+123ZK3SpFrKmHY6P0xOfvKz
pOSrOKwt38rK3xrCuZSdYsvPxJN3w0mwSxiN/AdwCc7nddrR/3uKFhpN9twsmj3N
UbXSSZypufFNPVEPPwqCewVRuyOMIAPkkxXo7a6HysutJuQvjQzS/UY8GISf1Bza
fTWqEJAG4w/AkYQqmsfl8DhtpFENTvyUIX9+KB3MrtU+8HNJtbPMj2DFqFpixbC8
QdIoZnB7sBbpQHKgkfElPm05u7qDvkC4p2h/Nu7HkKhnxFclN1MOKjfPEBM9K9Ux
q7m2mREQ0++c6w0U43S+MVSKVFVnDr9savAxItcjEZCcKjVNOhwKvLM+5aN1Qrmb
WUCSfQnsV0gD3wsbvcwKtzAtY/X2gNYrf3wVGViHDb8uZkg5/muMLCBTs+7uIIPm
hb/18N+G0AkA7uLw61v+bdmBadMziQ7vnnnz8f9a/4CuKKimMgBUO5uVKNLvzD3K
+MoGLcN/425+Uw0J2nPj9UFGlLcW5zm1YGeBkkhviO6fzjd1bGJkmoRv0Ezh9lO2
hXVE1V2bM/W8lDAkV/5Y/bcNvh+Mr/Ol7K38xkjkXUxK59Mad9EHS1PltFDKWXv9
CBiV/8RDnXmyN05k0urAb26XU0RPkCbAYpkf12/1/5U6esaZFDplaCAwrDP2o9tk
9pKR0pQqdcwNIFEy+F864CrYPQt4iBM3jde+lsj/6NTCaMn4i+Koni1t8h7T9FOJ
VemfyC/jcIcctl7otBK056rT3+GinSOnsu7VM1Et74DpSB7eiqboaUtzchObukJ7
cUz6xAhj0moVJfuwbPCB104Qvb49omwjkS8M27K7ELNtsadlpSmzNsW39Q7J4+Dk
KsGtYqQTfSmEUVrskiBucqSWIeO4EzRBE0ITKP4nk6ce6GbM2C06lr/pNXQzXQzP
3mu2S7LCgNyUE5GW4Z7gFiOeUbbZPnYs8ELvTq/8auqwSZ3C7GCVb7Iz1zgIo2yB
hobZcDtn6i/Jlx7GyGekGO0if1aBJ1Iriyx1l2eB6Y6qslOHjybx11cG0ZyDqDKp
5E/N2WP56P3H//5vetfBhznCkGIt+vCsIvUWzyFCjIn+a9bsGA5GkjOq0A9POdTo
Lr+HTDW+7pJJF58nS8qHVUjgmHmadBekZVLoW3F747yHvyqLMqFIqH5Rcqfj+Pn5
M1ztUbVVI5nuzApK5fqhBGYvfvCyEz0+ebhoU8ztH5HWRevyV3GxeM+JXhKsg9Nw
VtWoHcYYEzW+YK7E76o8Q00WRIYqBTDbeob4/bc/fI82g0dIRw+vo68Tk1kdob0N
GOq5uMs1vHPwPaiq73K4X6kj0ew1BXczZrT06qEWfscFc05ExOEtAIjVNRXIpI8N
gRcQnoVG8vQ8lxvNWEEtq2HObOd9CiTl06r/1HBvOI3kLrQCY0/pQ6MQ/XE2jTYr
kxEUAAkXOSknpFd/VvutF1xNH3MhMqFSBVk6Khi5oePi4AjvlaxI1i8nnpyx92Xw
WOIzs/9UMCVfkn7MEDK7GgSrrqiQk9gA6nfGhmc15bCpPn3R9hVlKqRto7ErS+QY
KobgE+WA+JdQsWbV0qocH+dGi4zjGiKv0KUTcSUyH9p8T7T39ObhKqEzGsMckWse
mj/umk3dBC9oBUvBhK74GsYkILHWEx0jpSc8txeGXi9F1MF29vGzJInB+m86M5Xp
sJHVIfFyEbejxQVXE49Yc5kejeT0bZBvH9fzriY93wT/xS20m0gYaoHuGU8Ndcfi
pGOcQJW9waEfuqHucm/nxkeANL8lrYZgG12BQkZKcHXii+/bnnTMtmKYMiqaKZ4t
O8MGWZ9tEa2xA/1vmBM9O8qoeNh4CkQd5CiZSdk8cBlj7AtYWxwGsa7wl4h7Wpn9
DQ2GZNEfNK6cpNqEInmf1/nULpXqmVeEysuq8B74V606Q3J9xHLEzCysAdZjxlJL
0sxs1xMm7TrjLwn/hC06Y/BkcwV/GL/NT7sRhkAGYoYqh4wx+LSOEsQh8KcjD/u7
HeXuZOjACiTUlzeD25NaM0dXB6FYlZdz26YOKOKIXP5RWiEV1BgKTjyePtwjNOYI
08xma+Ejrw7pBg4ewekyqZsCX9pW4Bk079QDXtvUJIdJ8BBtHq5mVrjVag35g4tW
BFQ877l3hhHPMyXaRzc7Uaz3J0lNHbaybC9JY+htfD+eFTdHWWODE/lLDon7Kl0l
ksgxWTt2AUJ1JGTCvt9+UUuqtIjelneoKf3hAzlnCvyqxNYHOET4aK+i/KYRz5UD
6177iPXdyxrn8XPA/CZ2tpAF65hNfbYJOIL6zljdc/IbP504TFlu6CcFltV9+Gn0
5XIUgecoWX6as4KFkDTygjARJDA4cFu/+e7sEsdU7EXLMFjwVpzXqtY771FWcXJF
8GWfHUJd2WG2XdhRZTE7opeBAp9+0UciuNiDS8CqHt0X62DZzTfsMM2dK6wfLv5/
dsBKhuPZDD75yG+yAs1JE8CM9VBe1el0E3mHebOj8ZnuMq2SKJwPmmjwkCFd7PVi
voScv63Ntml7BNDMKJHVxHDEt0GmoiKMssgHsQm81F/Y/xe5x01HLHG41SmhoWI/
asWV9ka4jHn/he7d6cTHV61eKGK4Zlxc2OJ7JDi80lhflKMFOxU+/fw6pz6tRI0O
WkVgwIr52+/ECjdu9LQ/NsmoK5eMhvF0afQ5m6OKyN5DAJGMlO8iS1v0Z0RZ/RIY
RCHgBKtIxkB3iXIbk4tlZqWHTg2WrmPZ8+OeJHnUlMiOVHt0lvI5Cz9JiUqgyciX
sdbfFd72ypGR998NBklyI6vhZ5XbtRr1EFDKYtcwTUOPo454cJ8DVW6O0d5BDXFv
t84aqU073jnl+p673ZQ6Owf6mZ7YAyN27TtPQda6oXViw5Ev14ANhxyYBso367M0
i13E/KLHWol5VMB1dkjgQQQJxPxk9lBWgG4rOuJc7IkifjfFCre38Quo+zScgM4b
FAnirxMzZgEDOUW+S90jCZtGDUf2uODfbxNgsiRtvhiPGhSU4eLZoxejc2P561ov
aRt5pNaU0oNLq61kYuDAEBjKasgKGqtrIgWENx+RPNp1qRs9hSpq/hrpEZKtE0VO
K3vavN4saVasSDgijj8u3oaWXP7hNvye4EZo6fjaLzE4UwNeTBcCvDxo+Fv8Knd+
MnfT2HljI0q7u2Ui0rppVCYFDrWU0+vOQ3vcrXX2OPtnsE4t4fRZj5i2BB61IvJy
cpBr+Fad+bOmPOTsOgMPpuC6v16rnX8PZgY8aB+GdIe+07nQhL3J4de8z5+sDTZC
U6HxMm8k2xbMlyz8Nq6bb4hK5lmuEQBV6BEJCGatryvLu2FV+7HuPK11mLrqeNcg
O6/KXX+HZ2w943W9vUZ9a9b6ewioKN7/DBKL++bgBDPhp7KGAwgfLlhD5PvDk2IO
rHO3SpeoKj4poWJmEO6P/8PYFQSTj34ULY2rasCs2MvfBTaFDbQT07RP6k64nEuP
2vNZ7m6cuAXUg0+L7IrevxWTjh6j8isF5hPJpNSzA1uVYqQ41LPAg1hTR7/SqwtB
b4JiOXD3N6ibHIjD2yjxqAUIg5IEwe0JZF8hQh9QvK95h2jnQAph+0NzVRV4kC2U
Mi4x285Xue4TFlx5HZT191XbI0+Y9UFaN+rt7RXR7xGL466MKyOcsf4NAC67uN94
eMz8f3+qWjmT0t/EdPSwEAj03KoIV3vvZKfH51WU/591Bl/JsfGwwxw5SQKed9EU
P8kQF1BIdHOMeOpDFAtNf8X8Xw72SGX5ESr1YUAz+UbDyRlBQ4x46wR6wVTsfyDk
Vq1HhtQEyc5i+xVdFJnRb1atwZVyogA8MUdcp9MM6OZ3wI0zCuz0BcsS+EF7CPcp
oE7mdC1y1rR6r6ZD7niDn1CETv2Nc+mgc4+gsacmhkqxmJfyRt65m2goKkSA9HlG
tQQ51l9Fj3VsXJdvHilphZyCgdymcr7mrg04ac9BQiRSz5V6JceV5hZ+S6csmpWX
M2kAKCQKaifTjJcI+HxZMdpvBh66A+GNSbUYKxTdAP9Whxrpf1MviCRbkfExExyQ
BQV71WfL6QENw7uFzOAj4InFRr2oPiL7XUl5rYCgLp2cmozKXvyQWEJXwMs8BF1A
hZxhUFtKyDgW60UiPvGPg2RlDiqlSKqnPHNziB6g3p5qXR1T8NUdnCrocacQi99h
zzmCxW8RJ0jYXUYJiJYRQm8h2REST1uJK8Wkd+KRhMEF+noOY+dv7R0cyZsLbjBt
mBo1zZ+6bdXX8IWhZiijxdVkdxfGq8dIdu+vmupgHZ9psQ3wgT8MK0I30Ug03BiC
UzHaMJ3f4McVNcjakotNoC7WsT5lm8Pua5dSws4f6YkL6nQ8h6ASa3WWK9HEoeRl
yh7mIyrnuodoXgZ5I6uGWwMCYLL0CeAChRd0ckxF9w5ewUeaTetYr3pt1ESzlAS4
rfKsGYxMtIG5+M/uri6dZzRJ5xS51VqEeVz+IFZGD5hh2KN9dItTCMN6O2a3RzEq
2QW+8yTuWgWj4wz4xug7haVwrDnbwLj/D/E/cySawRrYdxweaXm9XoIWFYQf/xFJ
GTG1fBYlzpK60/7dzrIsPHfz8WnqYVZtQ8buhBX/8NsqqFVQJs32i4yfF1bu3A3y
OLbB1AiShHu1Fn3GscqvmcHVjqZhaeDqRXEiT5xJ7qIdY12b43ytlnJgPqHCYVcY
nwUL1Cmaxwq45qaqKcep3L9OAXu/djg0jGe67ZDaJd6eL8vzS0ijgL/NBk/xG5yU
81WkfCxDnaAuCTE9M6cmceRoRr8stz8/evq5dAlqUotWAGh5oQfIdJv/uUlk/vGu
BKaTEZITxJ1c/Tf9JuheHhvgRFFy5WJghh+CRYS3nbFwIjkIG6gVlQMtOrUcMBou
h0naLVmrS4alQ+JAOi8xUPfWSr3iU8Zl0MvDNroit+30hHLtNRaMQgPaVe0MjLja
uastaQHiYdD26QrdWP4GYk66FL9iJ0ij8f/AGa2zh9dQnFXbnAS4YLodWovVidSi
8XjkGaIKtClV2xNWOYa/0VBzMSWzpsoTzVyJ0qiB7/dofvFavRnsdaWbUCzLxItD
6otgQkKJHaMqi/7TbyvgttBoWPmpygAs+Hr2pcCSBf93zwd+BUjZFevivLlGXCIv
FWJg3RBmUHY8wIsh2fn+aiSm/krODLVxlbCcAoHhi6tpWnLVJR/hnLxswAFj0VKJ
z/f28m9kovQdFa0r/U83ggD3woKYvnrz3jECZTP4d/x6J7nClixhMPQ23gubu5/W
ke3Hv4rXdwZuMSnq56MXlOS05XKR8M9gOafQHMShijOp22eZduLyvcwJyVSA4tiK
NT8IJylGMwsWmtyWxCW82zUZC1/Ard703YGEG2CGIbOEiT4vG67uWmFdqheE2wir
qbFAbbWBGV7BNlkU8w8jTG4AW2jV5dfe9F6uDdiazAvpGOSq8ls8swuREKXuDL82
V9IO2sE6UwWBiK+e6bKWpk5ewPhKDgU6sQKUscHVCM8eSPYjf8WaE9ZCIz/wgsdN
BuSLMNb1Z4Y5i4AlgMQu36zZ3k8ZQpfHIRAaQoBbWgG6ihU3rN8h7Ao1mNS9b/EC
yUx3V/x0JGLmWRjgeQe2Dc196Hj4hGHiASvt4OteXYleuxFwYxwtlJOgUO/m/11O
e3QQzxSXB/F7lLcQAOjE9va9CtUqwMJ6LZhaR8ytp9ErPlimBeXQSJcmjtWNS6Yh
wgtPNQz0MK2DaFoRsu5q+ipPXCKJknQSta37w+/4csSm7s9AO9M47FJ9w1qDTwz6
62EPXbhUfQ0vs19p7tPtDByt9t6jhzDX5in9jRtHt3VrkvZJlOByo89DxY4XwhEJ
jozAvNIVIIoqEry3Nc1AScDXjs/Yl3KAhxcxHT2qW96stsjv4nAO8krfRaau70BT
s2xV1uuXt4Qh1b+vSTEJC/U0/SuPSzrSin2UCaLpoPSoQz/ogL2/0rJ2smcigi/x
97M3ZBfLuj56euQXEV9Fbee6HCZtaf55SS+irQ/TdDQ4K9XJNOPR4b6AW7AtQJLs
/CkkpwlCGXDtGtYRTbdKWSfmdbaS/SFFzUKKzx4Ro/S6r4bU0OHdMVC3ykKv5/KA
jOCcEBPcM86ldInqqFZM9cnqZus8G4WYJ+GYhpV5KU8xGZNYrvVko98rhVC46wwH
2wVW5nqc7nyvjkBuSLaJnY6V6i7Z4a5FRUD9vu29YKg8zdH6inwgwTJA58vn2d0u
nTuccavYWL8NJi+cngmTReb1a/3ZfSbCdrt5+effhA04BmXE9XtGJYPz6XLRBtrR
67CGlPHJkZ8SKNYRH8ryD1Xhm+Rv5RPA9kECA5w6PKCyNayZnNDGHtxlzDsKT3Ag
hLvvfQwVtYkkwqbkQ0OmUVU/I2DnJK0ftjlLzqUH2NwZZzadSU/ej5dbGH7TLgTl
CbJLeHN0CW8h1K3YxzRnrlqpvQ8rGfyfJt4xqhaPccclCfUT4E+BBtjwZ/S2i5di
Nix65fUDPgpbwisvCaIywhkhOgmngm0YVSrZgFZ3vH0qPtM3e67uj3/famjlHDvD
MDhZ17FQcEXAuaognzsApDS3FyX05ucBUaMQJlOwUDYOIrtTR0ocBbvHyZ0jm0KO
TPOzDUC3GGj3g5sKB5LEoU19VDDVscPjsZrjO2cHYK+3+wug5eWWqyJ+kxamoy1O
TE8BTxK+1vYMgkr7mlLwqWFW+MP/Fm/w1Ntf93TzKrzSlYexiYqE5YP+oBb6FOuK
LR+8h13l5fHeUXBfcSdjC3qT1yiubyVYTlYbO+3i9shPmg3K84N/9TkFutQMjtnn
q6a+XEZbKoWUGBRtEBKHScrG6Gs3WhBUlUY9gk+AAGNdkw7A0BXE4xUBcErQVmpl
Iqvyt9BJlJmSGg3zUhKOgVl6MbebJq2Xr3jHKGXUv5CBVQPpByHRWZ8ZaiNlKUwH
urq8f82s8a5FF2BNwTIK0RZi3lUUZV1fggrz+JWkOVdx1mGr6viSmnnyXE2CdByn
UaFQAOLcBmzBtXokEAxcBYHiLwmidOv4csQkmj3mKwiZDKqLAFeYHhFyXfnGL0At
PrcONZeT4EcgWkr5Ss74W+wop2MhfQxa7AdXkxOmN7LdI4RsqjTmOA4vp7N8JG7Y
/JR3wipLw03gvqZUDv7k71NC7mAoYuQU3SdxkCn8SrAc/Y9a32UCdwuQ/Y0kykgO
Ci0g5CMfMsguzYHEu32XmXG7SMmAfHRl05x12UCph0E2tjhwBRs7Mf2V9uA3Vye2
GERAsLN8hlRW9zx21lsFUJ48CH0pdM2FLmef++0xHtCubn+eNEKZZZY8GL26G4DG
I5XzJXqdS45oo4AAan1c2tkWJ1JcWOd3zRgQoJoNX0YD+qnUXbPUIyXIsnuFsS2P
VCMN9/6VFJ0/z50YLuZUarwi6qNok2okNcJHXUAR7208nAFZHBu/ol4IuKVAiIxO
sMawhPkBnyo+uxlGDjImeUyGSMZK/oSTC2JtW7ZFrpla2oTSH1EflcMPDcwmWP96
M+DIXexAbsLof65lMWDNO2ZXKGY13F3OS5qCXXyb5TVIvjFfTjfQZCGPt0lAQRdW
QKJjJi7cyBOQNBpA0IMT5HSieZefDHKghyLsiKAa+SVSuMHTyj1qOoaQc5wfbAmH
HIn74dKY1VuJB4b7AYXXBxQYnK4Jboy2ZyvvSLARdCEhQNgaRftnynPraxTZ//j0
pUwfFf2gcfUkEF4nupRzW7RexC+DHO3nRZwtjSlNTSYlzADUFP/WlcPm7Q+jkMVq
t4Mkeyr9xx+VDXEPktdoI1PXLpBKNSUDXS4o/j4W5TfH4plthCG0yCvVz9QaWQow
lulEE/7sYOSGIdRwxf9R/1F0267D3mNo1f4YYR8sW+ax/6SEk2D8/uBADD9v237h
hBDdCk7cMHJzeGhD6wFNegIaUWNBBfamBKs+YQJr/7DGOGjPFOA2fflIcAQe46PO
Dtn6UxljhRa0krYbCxHWW+1GSln5HEMEVfKDea+lLQCMvhGKhfuYv8R38VvkxILB
qxabwmMexkWXAKiThfLvLIUBjPUAVyk9BLQWQwwga6IsCD05xPwdhdlKiD9nnpuH
Lj8mSmdxaSiHVGTG47s+dgLfTXrcpTl/REx3yk+4MpiKg7BG0CB66QeGvTp8mngl
oQ+TM56jWC+UeumceLzd6J1ijbBqjWsGX+DYPe5BvexTc/kiC8p+ZUR8ecdZfi8/
Jtf/ulD7w5f4vggPQgUOa7dL4jAp/u8zz67MOYnfXzTrEjvpkz9q1uKa/LVSlO+3
7nwNdtwvUqnfHuvi2rlnaLvcCrsaQXT2noIt+S/m6I3EeQ3xSkQjxh7n2xc/FFw9
7qTCo+CCs1tg178Qll1kVXAKe8os18S4SG5lm6ivCECDCkBGv/uGM2n9S/uTbIVy
nxBgtjsr9VxB4/N46sr3YzQepcBY3rL/V9W1yqN+Zv9IMKYfs5uJOLbn8QTVbP/T
F+Ly8wzQcuz1+8SO0liU47VXzgK0sGnZ6u2T4KHovUuJF7pEnbigwQFSlej7A+EU
19WA3Tox4OTPgdsZwEWG0SbJ78frOZqaNECKqqjT0KPIRQwiDPihamKlK8pPfVra
tKSfRsJ/yyv3kKcNaBDJiZSvqSTau7fJRY+CKKGGZikUIKmeI72LFUZdaICzj7z1
DtLAJD56bcu1EeoUMWchG+VNtwuspH5LGzDcY3vFLnqU2z5gvPTeOhvmqcEc1jkZ
7FiJFGtTWBhVIDF/IXyTztFKQ9YBnlsWT+xJFoTCwFtq9rRBKbzXVKhal0OmZ7TH
TOUwkD1G2AfjgaycLjFHtZLOPNMGn/JHxpsuHehYabviY1DAs4W578NjQlT4lYSS
J2O3hRp2aBOalh4iYaXXh1BC4oV9aNMg3/9fk3oOTdDbcelRpDE1So+Yxujsq2mf
208PVs7BeDgo1atymEJw+JNUMCH8iexJx7/SD2crOB5JQakj6oS90MhV/B0L78bJ
NwF1ng2sGJdkAD4G0om2zxDh61ome8/vVae7ceWAw/P/wL3YLfxSkJAhtTlm259b
B3JtXGWxw9xGtzhvCuL9hnpmsiCZ79W8xv4miu8O/fR0HgA8CNuTeM8LttaUkNJw
3aJl1zL1WrUxDhb/BdUhM9WegSsT3POCH5rfZ+2rwqh2WU0KqSdLsP/bWgNKg1Si
gEI51ojoEmaOGOmfsSvmzJmazjaT+N99CDPVXB4PVeDs/DGjx5G6ZsrE+dJpvaUs
DfThFyeHyYXXU0hJRTsBlAzY34pu0XRDj2G3O5P6EwQUdHQyFFSYDz6ux/pGZY1z
s88i3kbKB+bPdOFhdXt/SBCxP/6/099aQZaGYSXcyfM8F4usjFrlbCZeH0Wzno+u
SD9NHsxpR+rOGFAFF138B2pbdh1blCz9fh7lmRhGi/k1CWdp/WCGtrjbTl0fUVlV
3cr+CEzaFWD5VmIgByOlj/rTcb3cpHfrCFRlxD5bPE+JWtcaWjaShc0pdxeF5YqK
8idxLwB8JQSRm+gZd1RSc1enASXrIvTQ89BUDqTn03u6r68G0v9Pglf57coh6Io9
pd0m5sZyIZVNbIiuMyruR767rEchd1TKX99K8XbjyQMehuI6kiGjYcUHcKk9Xc3n
Kqj7AlSS7uCSLKq6ZUR8cFY8Ao0xNyQ+0xwx+qKA/Mo1Ajx5/Jjo1ZcnAv2db6n7
Xk5JgXEjzgSYfPh83UCxnLzBR43vCg47ii9MAfOpUxgs3IeVjb1vuxmHvLbMY6Vn
0R+Utn3F715yc5Yvew5sw1pvfngq62uOxw23FNBTd8J5MhjbbwstqZhf6SOf5cD0
7ZoUG+53g9wfJDpF1poFW1le9gS/Ggww78DKWeS9or6K9qtNV9zGr44m5X81im5z
0dJAsu8u4zXIr44y4WqTyOb64TC0ZqoDHSGO8xuMRzNv8bSLQTx1QK3wSFpz0ZyP
jO+B8i6KONIZhiWkFr/TwN7VObLWhkSoHxXJBzjjwg06WKRqeEqdkYZHuebF/IKp
Q4ShYLIeFsdbrlqwep/Q/DNJ2roaE19CEF5AfFM/fu1Odnvyxp4TgIFq7n/aEUPm
9CJh85W9BqbSMtvdy5/bH0AxQr10HLbGYqY48aTU7srn0wP2nZOTHqOADZLa/JvU
Odr7PFEwqoZ2P0ccwEdntJs2SCHiBNXxfX8MR4tdgLSPSU+RhFoM1hcpu6I45K56
MURhykJhvMx3UIuD80Qo8AGyyWdf1sGUCirmJN7444TcWpGyMIQAnIiszlxrvBFt
W9m6imIOH3PYvhwOmLitj+1rZ5zXoWNmDA603rOpbHYpXEtXk7aDe/appj+MeFX1
QoBleBfC9VoVGT4ov756dNEJjyYTi5IuMLREv0DKFALM1wyme2oZT5AfVHv5sFqG
UJaxHl+czhd6HW7SCabH2C8sWYxYm7EtUFHDg3nCaGQFDGC55u6oa6/g1/vxELgm
N+TDH1YusDD+CEB1iGupyfF1IaKOvLdSpLdd13IFfezo/g1MG+3diNW7fjbWaX4S
IKchTvCfDiNxfGTyc+VcyHXKcyUeiFB+SzARrM4BCGmR5QkgyM+BLJNgHiKhMJ/e
FYVCXHpH5la6WgPgbLR9Vcr4IF20eoKvMspp99iT+EEVWBJFkKLCTiRE6g+xWApJ
NpWSe7IJrAyayEOzu2HgBvbr1oSTU7DiI5sqZkMlPlzduczcZmUoX0x6pLC1L0Yt
rPRdxz0u4NKQZZo1+nqH4GqhmVsCM0RbcuYdavVEXC+XbgC4CEVD3tbK/64B0kdg
yXuHUbytP/+vKc+HKHLCGWCxIA3Nb0D+bskfU+AshmEzmER4UxZOE3HnOdh7fOl9
rcJvRLz0Vlms4v0r/3l+LArkjpGO8mn9exPEh3dVQrVvLbMxKwRrRDTQjoFfrNLV
0Eo+bbcZYaeioJAH9JRBX85NKq5nHmCYsYxXHSA6w67O8qF2qR4yzh99ce4JibhE
auV0FBhcNNY/BaC9XHOLzf5csINmDzQhjpRQTQa7bXvBXM/V29jmkFN0jNGqBDRc
NfQE47ZYmQ/k9Cmx0349/JYi2Zf3vPxYp1xDimhgBvESbovhQ5U/4YAlRZ5eFZf4
D4O3xIAJ/cHTIQ4FYoopGHOyadZHu4SKMbGnA94UJtyPfuYys73k5af2w/L1yPwX
88VNKZZSY6kN4MktGO2GU5sb71DrsPKh5oqUWY/uunQFDOdjpoUozQ0GredcMrns
wbzQBJvJeVwdLTEjXQtv93Ju1xiqr2rXHoX02MmvoAJKOr1YdDivWgrFTnnGyTOp
1p9XpxSol18HtkqEDT6FZVPlY7LhAdoV0vgI37BsyQ2WMRWo1h+wFYMZoTG8GYac
yvRq7DouShED4ZZhxhyZcr8i2qWPqbqFQcq2dRZHIUanghKs2gWTliKtqodPVK19
NTPsvVZjlGE7uIcUw9C3kzFb553fglv1i353vn3rilc7LISFw/szm00Nz8d0ya+o
6rDm/z2atVMWstdVcEQh0DRM2eB6MuYjc1m1d9BjR4PXSGp+E+1pQJdAOow7M2xh
FjB0b0VHM8GBrapw0tib9QX0CCN1VdgnZq2HQ0zge85pMT80rKQM1kCNTMqnjwer
TzEEJWc6C4xPMmHiEUISKy00AE8ntCIsQOX/+S+JrFsZKUE+lc4Us5KtfUmuLrME
RJxZgRjw0BuTeR62Mqw5q+Quix/KzICsF1sczljravWkHi7AB3YvblKOgrOouxb+
BaZ+9M1YkexBOb0yY5UevRpf9loe8nmPugjWVGdC4LAhDFQZAgkBJizqRq9up6VR
kjD8UCn8d21+FV4edQ1jtZni1skf27wGPvUdnhQT7qUapgDe8B6DnvyyYecWJtoV
+yHSl7V5dLRhU1xh6sWm0rwA6p+zrr2ua/9KJz5Itr7D7OAKimCI/RSiADkSG5Q7
z0sWeuYQScN9A2W1PbZxW84ye+G3WUtul53EsXqUmCDtgThgzcyXjCmRPwMr3KlR
T0psp4Thhv7/u/1Vo50MiXntpboR4tEBn8HDT9Vo39mFaGmQfd2+VdvYLg3XTsKY
azbZ72Bd8av9JonoDjil8M833v0KtSJJ50i9t9Ney7FYdkDBwkdnhazP4i5DIzt+
u8+IPY49V15ykI1qdqEvefOUYvOdyXeFJKwC/3dNl34bGhzn/fTqpFg247Mg490C
Uea1fKb0NmSkeJ1FEPxzVJL+V/ITS6tpWm/9bg588RhzDWEDvFIMOY3elLZzvdQk
LXK0SNt7UmR3kpvTRlDsuR1pHIBHcfcYUiAwrAvisvtA6wYoTco1XuOAsmeKgcO7
bEGBXJsBX8egDrwxBebj91ni5h31x6F6A6073OrQ3EU4OtPl4kBlOlwsEoi7isfI
kpNj8V8je8uoRmuxDEGsLryyD0cAhDvJmapfxnDALsK5OvYc0Sd86KQAir7zQRoX
gsohuUyCcuRDPX2cJHNxS5uOKYKSlbPKTsGnmIgdTrQkjYy1COZb/dNEcU8URv+S
FOD6UWa3zoahDZ1nEdEuNOW8jhs8YnLZ/pclPUqeYr0LobFLzLlfbs5sUi3Epuar
LI+DVn5IqslAJgnNDVZ7QBJxM4b1pCYsExcHK7Cl68oRbvMZzfi60WEX9wJvga1V
2zNo31oNOHfj4BeXnlVOPiu/4IheHUxoegSnCTyvbX/0/5Wb5+0MZT8jLNJP3UGX
FKlQZiVraN+MaBMSoGVXEpLLX7QSAxXiRxaz//FiWGIZnhJz26mQa+0EINqFfLQa
ZAfVMPdgF9/hClmo38knvyFbKiivq3AWPJaN89PNUNuTg+yo4ImZ+jHENuy2C/hz
IZ+dbNj2vE9BbgqBZdlSnKBrNQzUivyJkdUc2Ok6nZ8G1DvSIl86cac5QuDDO1PS
IZ6EtbtMAwXo2ZLrPuZzTFxxbwKA/7AdsRF+gPqhjorHlm6ihCDr0pfPyTPsp1Pf
i8voPTiwT2GF4yAuzlatjV9kLS76hGXKERXIqZGpeQiCZ2fLPi5C1cH7VKGXNtKu
J6ZUzLfDfw9rp5AJGCpzXyj8Y12cHNLvlwQSmdSWKuNQOnZa99aV3HZU55zJI3Hq
QU4u5qu1mAPN295uk0WXqb5Q8ttnY9L0LDJ115ebHiSp08M0uZOY67cmz5dAMEvc
U0ajZGNEhFdEtgmk6qe/LcsQthOokWPJW8RcWyjOEPbgP9kV6hsxMqucYYAWzWv9
yt9WZ0LDIIJyLZFSDiIOjZsrYciSOSxjX0zdVBeqkt4VYly+HShKV3lav1jQs4lk
KJppt5lLrNfyvF/a1oAkUBwamsCgGP3+zz/9axaaupx76SvoFPfUi86UOQmSyzrc
3s1To3sxbk5Jj9YLqEYNK0BBIzm4WQcekwe+zIoKtHGll39MfVP6a1CWnjCnv3Ms
bmIFrLl9kmIHljNRRTon3aw/5pxrcCUt2tZSxpRVQ8AnH37GdXIc6WuGIrq6imvi
yqHc/kaj/giw88+V0vRuiBPrCrroEouftbvBn94mjcpduREO1qYCe3hkwtLIFnfs
u7VchUfROROoZxgFDxzeWfbkYZr04SvIBmMg3wElU3YbYdh9GUXsV0nI/yyBKwm9
LGrHWnZNNuyR0MOx9ocfUP/MS6wN/HrLr5jtwSbL1d02ohKy6Km1yiQUDoke66iD
i2f4PuWyjhWAGkWq49uvUkQjTuoGKD+TnRyPP8HYWG/dWd9PXoa2PGI9LUNk/WxR
YDaXyy2SzoVcRby6w8sECG91iST7fRawKkes5OiZoFfXwLRYfNFsI3WI68uukIoy
dNWEHi2RS5JWkFfdInbjoEzgIkZVXxQxavAicWoD8X3iylieq1X9U2moD3sBlECg
JIDEDh6lVuy5tAQ/eC3kppjr2ahhFU3bxuxhfwbvJC9w3z2yAYrKlp7VxMnUEGEF
rJjqlX09FjwY61BIlt+dztmBL8ShL/6H1CayDmcWNHif5cLp3FY+dNgYd83G9PXH
fkc2tcIvcA+31mFSV1ZrzYDZFnE/+DsuAefpx5CCUMOF+cZBcNOPUSIDFDSvTcyw
jCr5ZkDuoVI/Om3/LaSsQtTluC5KjhTCBAx2+eZdE8tRJYLLn3rG7tf8eEWDszw/
CaFANUciu9+tNl/BKljeJlij4r3ZXqM3XpWKbXLEiOBucp1fNX66cqH4DgG0H76e
nUNnOONk1baqH54S4NkIXRwSPhf7DhOH5nqSP0wpcD0rFnS3sgD2+DjSoIkgTJjh
tv5muVbEHtVCJLx7IURCAkwnWVdUDvgGcWuM4ML4kPtXV3qmtljpI/VuRe+cyEoc
3bolldOmARxVmTRObhtUOSBrd+uYEEqpM84/Q8Lbbjgz7S3wszdyvF/V0NPCbn0O
KQ15nCm79p8x9pHALcNjpDpfR/aLUyie0hl9rUj7EEIXYqdDacCMFuvUjvwzJFS3
Me5NR37scJhj7LnZw/iyrFkrQuVEqmXcdFUu+1hIBGqj9D7011xhykakFdoMZ5kK
nvNv2pbbS9SkKpUpDIqPLB7NOnKbNdM1bMw92hdx6mroTHiBXxUX6T07ydOkgYeR
SdsId8X9b0P3Ds65Wd+bRkUdNuM1ph9Hzp330grEKTNEhFRN+Tp79N+BOxJ3MJ6Y
OA0eMiLlZgLJwCUSJeO7y86jEh2kYJOgDbJpmWZK77l02ubU6jMJ2UEcBWwO5GbW
GyjpOufmsItBRRlS6UpTBQZUi4QlI5cDrvn+XbOdfiBIhhmtPQ7ziEYkuaKJQbeZ
b4brIw3O+2dBbwLOCHcoetnq9xbqGfCa610BKjcgO8aZYekxolBfbHbV4iiaG2zg
OITEvFtuUBNjMf/uPS7Nvmk1RWPmLhAG+rbE5V2Ec17WohZZHYDNIXN+S6V5bUip
lSd0XotrKYi11ZuJ2cmnFp7P94RSaKR2/Pamdfb+FbV6SiNRQ4tgAQlBKPEAzmqi
dE89I9np1r/jK329DJGlrwQPlWFG57xL5sul4ll8bD1xuq1iBmBzATKflxig2/Hc
mKIJGkqLTPoqP69BLfnkGqA6zJUAd2PxQvCGUbk4vxZIJ06FjhGme9u6IRpDeJoZ
kZ10BCD5QKBWTziT4q5jJO68M4Ntqkepn0dr8mIdB3HNLWeVMmA57mc3ahNltzFj
wfT0AXG+K688+bjgydgB5ev8clEiI+C8zAaKTq2S9ngd7DYTB+TdqAVkyweQYQKZ
XXmlzeue3lhNj0hi+aIcX3ibuWqchXcCj5isJGCOGLg702aEfj26hbGVApvh9nK/
HO/IpPbhl3lNl2omeA9a0rxnEPUmO9+41SOsvbRS6BLwhFiT0LGQQyB5ez2kJXMG
AlIAlA3bCxggfdNpv3AmBwpGSF8ve6Z1YNrM8V4x4XOLOJyvD2MLcl8g7i66wv2a
O3Qk0FivhVtUpDtNJ072P4sXDJkafoAtjKYTI6bnwRbmuHUbYuWxUGSfK6/pSweb
Sh8k0l57JuhPHUqZMXNlpwuSZJKL0A3Gn1e7zjK3KCX26NQ7AmAaAzzCeRd3PaIq
G+O9KMCe6zNFwjdzchhdzt2rskX0D/NC521mFY7gedCv3OvzpyYjdJTEcw/9kh61
ozYlu8DiEb16w1rnPjhF+JTH4xzR5WjcDL+aWShzqqnWHafSMeRPGAL9lgJaGh+/
kodd+nHR5NyoNsx4F9EYcQ4cQ/NfTmrf2hcpvUIhHMBmhC+zrb98wXGLcFtP6dkS
16im0tPs6U1FqAS7a0zB3hs6Mvp59+6ntetxu3wmFW/FTt2kRnMTZ88sFCu895xk
uTqJSX3SnTt3UZFgfMZfLyEkJmfuM/MyZI024yj85TqN9qNFq10s9btGdf8VC746
7Q8Vx277a/trWeLmcak7d9QBqyF/IKynyWC2Y4DjssV+L9obgZILltHSyBGR9w8S
cVHTu8D7AsQpPQw0s+T8GCullvI9yPM+dBZi/50pxhIRRi8Ow9DBCGYvuw8uxhKD
TGMa7W9D12T1DyeUtl6zAIguCc/0OvPWxzLT3W4Yak3Jnu/SuSbOi2jNT+99E3hL
Upoz9qOFSKc7q2dcSHCHakI53xurc7jfiUKJR/Bt/YygSHpeLSqET/riSilynh/2
boFy+TmYm3m4n4nKkYJFw0/e2XZhgv4YnB7CtLzd/rzH3pcC1e7RFGc2S1BUbOG8
4Qu3i7OuxsKPkHTtUlVdfLRABORLQoG3JnOdfjDrWHBiro/PR3F9yI2/I2XaYa/W
wYQHREDImyUhlnMH+IfPuniPRr5YVPBogNqXkynwL2xt+eGnQasxgGskBDyy6pdE
MzHku90XBNOxoh3Ibtcojqi+mkQgMIz4wI79PwKzGobncBiv5QnJ1LSHpvehRAnw
QhELHRIgaP79fsVH4Q14E5jAGwJ3MPq/JT0TV/u9YmiDRfr6mqzE8v8A1wAd9jrU
Uro3bkSRr3mMrCkstVf529/1R+viyDzRECzXUf7BSY/DTUZPlZijwNDv1jaEYWGw
CLz6C2v4OJMt2XXTnvTQYfeTBSznR+yy5aU7Kk+Mo9x8vso4+eriII4IaEelrfXf
dFNOrcu6y64qzI2RoHwronFSKBUy0jMxGKMZNrnxfZtdqu5uYbj+/qquBjt+4aWd
wCRpN7jS8fdUglKbyA3nnexZer+bgXaRnH1zVrK8zw6f/n4w9Cn+8xakLQAiIrwF
4N4NEKYuZMVZ6w4ayoyjS3dq6gX/OlqBQW4uF1BpC6cq1bqMAW6UsvTUwxHSEPGM
4VQh9XgAjnWoV6vg2Yh+wK4miz6lwQarTfu7ZoEcKWx++nrdkOmeCiQy2pQBQjem
boVvtgeqZ8NNIiIQEqac9TJYS4VWE0H2DcvO8NJG6JRwlzY2vFISHaB6ml8xUa1i
qOgJNpPt1/C3OzHRYPgrB7zos0MTq+kKj0YUWE/6ZvlAV50dyQJmnKTqufmckEgd
ITic87xccyaQW8XkZscbKvmrt5Yyuye8JNDoquOzSp/m/Z2v2gEVki2AUB0GIZsw
n0edXRQWVzMYocH5HtUZsZlpN4+wxaAUmwbhVriOfRds6d8OaXbExx8V+tOqvZdj
2S6pPBbFMf6f5nkM8uejC65tVlnLSAIsFK9umSMvS10rrrVoAE0EMqYp13wbhEuZ
OZseZQvkOSb040QeBiOSyoLkHw1hIDDLnMZ8vMUt2dHUlKbJbsSkyl5uFmngTWkg
XO2TOItrZ14go2J+Mrz1HBRKGZCOyTChOBr1HoUnx43jSZVbp2MOe2jxj0bjfoyn
NarHWMwzKnSnkNd6QebiIdARvXseDjXNynvBBzV4M0lgObtuxJWUjO1N9kUTvUUp
BlWM2VdOk11W1LIM1pNpFgwCaXc5LdxJUFHwggXRH14RG1/NpXKXi2YiLF00Rx5K
iWpbqSl5DDt/qpfdE/ThquKQc1tes2vR7UPAtRvzMtLyBPKXO4dYhytIJLBhaS96
F/Krg+4RO83hmKb0fy19eGCZpqdqU3u1LkGMOrn6RgIDdjpxr0032eXVmAXPBOgN
uZ1FV1mviGj83JRYRKXDWy7kTZ1AX2EcTTsF1QBMGLIvinAfmakPfRY2VYESG7Q/
HYMVBbJD8Rolo7FfW39RoOfz0Paf4hI1AdV092SZE2NffiZy9r31zPX/m7ke26LQ
koM9G+wGLClE4uffXAliUzqK/tg9NhCcQXr0w1Y0V/8NWrQ6UZs9anSCg2oQn2RE
Tv8hlEVxBejt6dgDF8h2HnBIRB0AtwAQrwVuUJpJVJ+0xPzQLgoIlVO5W3M2Q0H8
Cv/bpc65y439dUJI2qLIeIXNKtODdZCagVBj2nD5KxRQRXcTBEaj36vcE/grhVtl
EYZqH98l8b05gtEA2afPFOeJ4T7avhhXDzGSEf0N4H/B23bzxjhzi82zzCNpnXbq
WR5hJWIe3zDfPUJwU9IXeHLB2iy7mexds89cwssItFmjYA0F6ZcqzMXlgd5QoUdb
ai56Eq+hTG5lriULcogbu/HYGSn7vscpHpaDU1/HOSgfVQbXdknNpg68A7u3pMhN
PIEIGy5UNS/4NWsWaiWvIsos9XbE4/JdeMHNJrcKZLZpUcmlHSziAdds0K2OsM2+
BdQKe7emNWWlwUKE2J/863CPqhF/KEjMCc2G9eLKTSwM4WaBd9hD2+ZB3xf089FE
q1L+WRY5MKnNyncK/N+5+3iOkSAwUWVPZ/nFrZoVsp3yr4Y7g+3KCtv7yINLmTe9
qXsvTOAQ5NW9PyySmgHv3ISVH+Ekt1y1PnexZA/at7wRW7mx5Fqp9OcZF+z8un2h
P6w/L7lQ9ELs7+kektAZ6hNookXqIctNCzm8i9wtWta4QWkzKTaH3RNmxyLCDtNJ
xdYidZM8iDRuzzrMltX9hbx+WJl0Ua7L6BjVhBaVSOV9XVRpPqPTk5K3zLvGFkv6
Xz5Mx0y2wMo/gV6zT01/1ybWPHVUlhpebyP88776ZPf4aPGO5Yu/42kQ2WODKiav
uAf4bB9feiIrmnaFiYwwF+I74yrX4Y/M2LPxSxoINhU7Ep6i6OfKrausGunoMsdx
c7wmBNOSuZCmf99LpiGwMcV3PCaziTq5w5r4G68HLCeBJ9orKmlaA/x8whu4AFvH
V6Q9yxbkY5is4HH3uDmKMgfU7Zw0yjbgY+2PRt5nm1l1VIQwPnwHeGkduGdGv0Ba
qWkvD50Je5nIjJtYme1MQFG/ICPSyxRIFzC5edbdD5gymfHbyWyvwPq7dfIoJYCJ
LMPtlzQ9wrddpPrfJP6K2qr8L3X8F+1ILP4Cf9idtuOX0Lcz/NHLksVGLEGZ27mg
JFcLjo95Ac+2p79z4o/MCY52bB7M3wgCn3HokReH40ifPFedaw8zzEEnkNC8rPGa
uDfCPsEb6t/nPIXU0fILh1ZtQeSiSlUq+Sz1v5MsjRB5W1Yvqhy/DT5OpW4ecn8D
a0kevFTczTxcceB6etrqBqBCICuHL/1FqRw/6BAPraDRKUv0jwnoTqntp1UsDrh0
CBOhko1y2M7LHJCzeP3BNmOeyJOQyj+dKzdkeTzxD23dzR8brmn3QBByAY9Wimu4
CO5BCYynlTWNxubskVuOGQvYAHPXpYRL5R2L1NNX0TKMY1StoQ0TaRX3ZCmZ0588
APgQLhUKAIGxN3ou6gAp8+jQBNV09/BKbTB/lnSefpOepuqWDS68qhAloYtvKGAd
tJyMesjHwP6DY+mDt0CdDrEF4OaCiT6lHVdb2FR6EPh702M9v//wlzhcQMgQeYBV
MFVigkYF88rIC3lVdOcTXR41J0Xs5OPlXThRBX/xWOoRIBJlP4+RcvVrp+QhyGFh
qLgzYkws2GVeS8VXbPOutWVVJZ97GWm5Hrk2zeXZeQiQSFLZmO7GL3sMcOBshq2x
p/3QtvoDulks+8Ct7vEZPhMGDerYxakomlxYRDfhgcIdtO2Ws7WyXkUh+cRWZ+c7
0iRf+mIZVIqGkx+AwJhhgbHTHSUnJ7V6Xa3TF0YJfX+VvGzYuiD5TlQ7MKRVfhRj
4cl3w6qOnq68RA8aaPoGzHuBXHM/XIZrgUFlq/MfHWnnOvhTNdpdCN2rqi9/4onH
pAtFYOxcxu4Wu63KlqcyJo+mp4g0kd6WKsE0U7Ggrz5FofYi2cp93f1l4z3x/2wb
oCQtIDXgDwTihThH4rd/hCII+tsTgWkyu+G6SG37ZU+aV/i0lUu0xBvIH/LgBWxf
p0e1oyybswuBfAkMJs3lLd39BCddy4JCL5BVftZcO0lstoUYySkDV59+cNJalxsu
Lc5h0Kzvpdyq2+ntrzF3IVhATrLCse72OWsR26lgLeJ+GSuLTpov8TTdFJZ7S+vS
jzV2acyRhRo2jNE1gveub/OVidiLPX7MbqFkyfghotZLib9oHFTkPuQMnOAVHn7S
Jru74AK2fSoF08S98suBcsWMNmnUIUOwAcG2gUcqGGTggbJ4lbsXBWBGLXSH2+Ye
h8I/xh/yNAA/Rmp5pWTVE9s21tdRmqRQXXUUsUL6k5k54UmppXDc+JN8hWNJuxv+
79ONXTdLf41H5ZWVq5A50UoLOkL/KGOho7jrmRI4ko+Mqu3XNIGYO6NwcJzHxVDq
5Amy1Y/89jW7jR5XdVdmzxM+hen8LZ8nUOgUKmbmwK+NbkNMAqgnV9Pfvuj+7Xd1
sgPcFqmie7t4VH7jFo+N0JxtPNJkBKiqDlIrAFb3N1xY9G3hCX0aHNMppvwCCkKv
9mOlRAxnh007PYxA/vxcMgorY7rSDmvAfs2SSPx3+nfnadaJvP0a7ycSeE3ibIve
esG38Kn/ZvwjeyT1811piJsq7f0bzseQNhc7k0qGuPufKM9/q1WbQS36SSg/DcPU
Y0zXXKS6p9aPyqOW+Mp00V0W7IZ1uhX4oJDecaJnrCjL7RgMvaE03H/ywxaukPBj
FvVRQaFttJaTT62NQzcJvtwwI3GK0zrUWqy0HMKEWFltYHepVM3FaJ0itvAaOlc6
JbM5iBYsDrEG//DqvT51eX2d2FgJjwtnr4OSZiZukOqrFn2s7kPi7TLMvM51wo0E
EMVdITuEZ6eJFJX2RoFmgVYeD/F1gvZgjfn8l++7EQGQpRXCj2Amdj+iwu33kBNx
wR3EYJGaECEGe2XQsL5w8ukK4vSBLpXW7FScuGrcZcHa0Svgbu+ZNdNbhWRsXkVS
+D0RLrcXlShW8GDUMktSsf6bhNthCWCORxYo3XpOrk4GuTh8T15HiKi6Q9WkKwR6
TnjNjRLOaaebx/KyLKRjO7vp4XLr0r1GNOcLnxz7JK3v39e0AKHA4TJEfwrxo2wK
sgMHQOLKbrsC3Z5lbB90EQeOiUP0J4c5Z772txtLKU5UruKdEqfQlnaD1UmL+uY5
swnw6lsPKvH8sxHpqtAVDt7CIe4rVE6HYc5cVMR9Vq4cy1AAW9ahiyJvlNWXxMOj
AD/APv3GxPDpGTXBpZ0kOelpAdv3mxI1OKPdRhnZLL7XUgZfRvVFj+CcQXtqmdeF
nMmovv2lK0/yhlWwzF0JH/klke/3bBJ7MMiX8RwmKKiihcG7/f/URhbI0xbLZBDf
RFgMd1uGKE+nflsTpDP7YPyd1UNp7lzfJrqnWdtRLphewjh3duyk/3CnuySedtra
VrEq6SLTbMxyA9JAmLtzv8frow4B7p20qt5cIiVKwkBceRdZ4u4G5nwCHAa/LsIN
OSCSRsZyTkieJI8aRyrV5dWEpHHMWJ4YlQamRiq7icq8R7BQ7/hjeOk+uu7okh8V
xexDw0MYL2JlZwurxTxsaIxndeZXIV4NRElkUoJThmzAMr/Wo5rs3hnXOYj6hme/
Qtd//nUyF7coQNxeWIuPQUdGjZXWIsWaWb/dYksHkLHr+o8PDenbQYnXoDq24DLP
gTXXoqSV60M3doKrUz68NpOyTJMz4MOyZBqts+DDwjUSqA8pVtEMbOMxqbJQGSxM
Sx/OQ1sGiRPNqUTgeeBJMnCTHRxh0rNRH7Yp+j5bzDi5Y9SeLW7Ce0WJ1UagVTHF
59maarQMM8Ows5P8i66NxhJZTP9m10Q0q1/rq/CerZAMASQP7brhTxVftV8P43/h
W3Kq+6+CCb2B4zCUTylxDDwQISm8KO//+tX6DQ1dFu2Gy5q0lfCnR5roJtWX4ZR2
pL4z0UVi5abFqENY28v3Mu/z9C0mEwVt8Se95OcewV42NnKKtC5nVQhzTHLpoXxZ
9+93a826jn3YwEGH2m6lxiaImIP5HOGh6sHdlAEnkgGXTdl00TQmby/DAw/TShmJ
k4fnzJiC9DrEFffYzucqKj2IVNCtFasYCyZluZYVAy2RwgD3Cs8ONMU6DUHLZGQW
A7mlletOFSAmaLnp+miFbhzzWkKa82w5eCZh8+FYaxk9cq4/P4yH305ID7F+GqAR
FVGGMl+3I2m+E9dYRHgvpub0NRvD1gYRGQ2yIZqp+5i6J+WsSWWGzURGqU0OkkUF
QALWs9nV3akjPpn7t9X+VYjjPKf240+IAm6XRzGmBzLdesjL9k4pHLbb40cvU1Gw
5V+mhOVacTgRJsXwBd6XNdLPf4VcfmCSzT110Ph06pdupcdbNSZoKSDXU0jHL/yi
kraKusKfbd7euRzdA41BQ2anVR69IzOkdrn82swfaODzRrXIDaH7zditNZKRD3JI
EydRoRJbdwFrtMGqaxF5dS5bHxllS/Gdq528eFgmuayC0TBReDhkutMw4Ci0Hudl
mfwFBnYxL5wQ75PFVzQfA12gOFAg5jOHRd8+JbaXwSeuj+BzdX5oMIvGRW+LXzKQ
NFq8a4EtKkfs5QFDwopYCJ9I0hJwsMDNYIzEvj/GhpK9cvfsfLOUKo+eHPdPjoos
jrLKejH6wpYIPHtE7k/+l1WMoTsabSFQ7c9WhbdxhMH+ySNXRzsNZqMcs1MzkcP6
duPdueErlJDo9jMzWjT6hkaDSV4yFwQ9nJbinW2XLmwPC8HjMhGeKuAAadMQloBl
6IgTFGwBklykiCH2R5HCTA0AUgDpm2OtAcoN4AiCo9oSP5W3rzOJBemHDh7Bm9zW
BHSO8TKGvfQ7lyaqIu2oCfa2nHHKOutfWuYbM7EpuU1m4EWHkaKM3+OmSLeS3D67
/ZsXvogaEuiQQud1iAmA9alI1kORaybQ5fMoPhDZwS1m4x94Ve4O/ohXiNxcXpsg
9O9hhzmJdUGXkhJKYlB6CQficl5pa7J7nNGAPZWWcXW4VsjA+he1eC7sR5smIcFl
8eoM3mzO7DLwYt3QymzyftOEK1i/qKftihS18nU9/bLB5ctkMCYdDDcouT25uBco
xGQfAX301H3LFXf9sSHe0HzTpitavbM8wl8cZnXcfiV6TD+PfqSbJTg7iO65dToY
WW2XA6bhV2D2dyXAGvH8JVK/dbxNK4xhWcu/hAwysgXTmHNhQnHvLPyOnZybQ9nB
IFAetC9uwkMPCERdKB1Lxmb0sMuqBMfj1DzC8Ia6sARflBOkdxSxq39OL0BBZSXm
aMoHiyWIRE68mmZ07YdJOcQk/B/ay+Nd67zQo7XUDaVMLiuNxJlM/KXOKLeqL4Mp
JYTKZSFm0jkl9jkO3nWp4n915Qkl2iZfYm6DjoAghxsxnsDCVO01zc6svaAlnP0b
wAf/3L46JXdFf7E8UCQknXPVwVBr0s6NrwTjqY2nt1TZpQMYkh7G31QWeuZLdyOn
tgBw8zBJtzNXHH3gv1DhJiShM+YpmdOQCfePHG2xvXdwKFX+FqxAax3W0o3nOHle
QXtKwi3X9C+0gzwJeCAwOvUNtbCKnFrbXzeovc9Q7WEmGkEPjOE3E8Zxc5bsN4L3
Jq0VeywmgLHpmGt8a2ZBVQyRsd/y7bfFZ2D4TzABsDPNKbYkPdmIhTtAtTtXKAtP
eL7yupGGjYdoHmnUEAvKdVjcRqnhA5s7Tp/1NyaLm10ukxcBOyxOXPsAPu2CUa8i
XH8W1qPG5WcjqK3YySd54Tv2Ph1vMK/PuiFD2NObg9E0baLPLv+TFLkg1q8TqK+7
BoiyMkr9/JyD0umxLM2mGBaWZjnkvfhVdjwLGVbIBkEkldmmYKPzyFMJYuqjFyZr
M8fG4NUu+psAHRIbY9+/TI0PGfd35OpbAUHrPNjY8XobSywit/QkwjnFUvBBrsJf
HWC26OsR9xtPP5dPrrhC2J18Jn8a5V45nlsYO+2iFltkilKBOEWqPhXisAExLpnG
xyF8kkofsbMaOmfqIU3gyD/Z3Y1QRmkfe/GTgTlcv/TIeb9j3DrR7ygaMMZ7PelH
fEBfX9/hZ8kki9i/L4dAzsugc24cEfc4jWBMK3wk44ryN95GuO3AkCAsHfTJdgoa
6zYBIW+j6vA8A700Uttpsy52qZWmcAvW5QjSGk5GamSRWZi3RJdbVNGb1/q1OkOT
cZDTYcEFRw2rynDiYrgTSZ0ShqDRxRD/O4YpW0fp/QHjbl0M8SIubldxI6skdOP9
YsNWuGT0PG8y15hv9mQsPIOWJAFez7KmCTNEzrTXrtbMpE0rncvHmL6Rqddpwn0k
oNsG+K3YShC24htrxcQKkkOVClRixat8yCN0IGltzI9AL01gmHiW2DXTOF6e7jvA
LzXyt+VWkKVLOMk64oDycvMfWLnr1H9e52z+hwn0VIZSAbaPCN9KairAlYn2nlir
b0FG4A1wEeJsEi+vzy7akzFOJQVj2+3Ci5dgw7Xs/60rzX4urvC4/jvTnzIKfHVh
EWISOIVBAvFVZPpH8A2Axhb/BiLWBsmB3cKPl1SrosiGMJAAMZkyym/BUcTeVLi7
WeSh0y3uKdPYWas3uP62VF5hFIic17VGvPYrG//ZrW94tFVMeyGaflZbEHdpmvAJ
rM4PBKO88cQYG+r+HfM2l3LoedAmt2aaY+H63S9RpSgYzq+GiDUpk/SqRfYLwzVw
pDOCoVcY/nrqekA5VIDTS41/zzeDPtZ/GdAChe3tjG1z3uwxf6FbekZF/PhXpmd3
1ovzgw6CnNFM4WmziBYxYFj64+57WofIMspQolTwzKnroWqRXmjz/BCcLOh2hgP9
sFff/vGJxKdLe7oKKv+8Yp2p+LcX07mdQNQavBKqdwSlV9gUbofxX5vJ7K1cYZ+P
IkUILleqIRekTCy3+PkagOVaz16Phusvyr7cSQvFmWfcuEM8hJ9WN2fqvSQMmFqg
7YXyVgyv2dAu80OUhv78Z/aZxAwcLHFhHo0flDbdYqj4OJnnZOkvv2PnUOroZKir
+PZTZNjaTCEaG2mTg1zo8bvnmlfqDc7sf1tIy2+lVVhceVYxQNQYsVozoSem4154
y1tISK8EEVUGqaPQoo9v0VLneGTp7dupu/1l+Ea5wMR3aQElZZK50w4pGbbC8uOY
yjsp59yu7O7+P0p/JZ6t/zA2T1/x7ckNx6K9R/x1OrKlxo+AlejB5EOzxoFbOE06
daf/dhGKCWIfb6V//MlbJuqbkQtzWvzp6bhlzdmDr0WEQ7W3NgG/jZwykYgULyW2
GTF2wqapI8UeNsVPV8U4yAvuNmdMPHyG8JTBhvPf0tTkO5i1hwyNSIVFNPyLdfhC
oUpOxHn/GumR6mbbZCYl8JL+ZsDOaADNkIvlhOaOQeuR0GrZXekfhSdnjELTsj18
tI8O1wAjY7KyABahoM2esLryw76eZ+Vx8+bBHm+JhIUfUkmK78meE491rU+psGZ6
qvVR5//Qj1kxXi2nuwsFzgWNyOz8cSLw3Ezx3emgaadSBg1a6XYd+DpnvRR4GN8B
2xIXzF2OQJqIhTzCnE7CY+Z+uG9XbxFSkzDgKVQp6ve2FMDM5CaZBusGNy7t8XH1
2E6HjE75GIUgpH7HhMg2ruOiZyTE9Zc1ci3JO9u1bLUSUjeLOKRnJlb1l8rmWStb
u5N+BkAuxTX12mNk+QhoSkujDCFS8r4Lo7x7VD1tzicZJGTAHvwlNS7OBRhGuoRw
7MC7XvhEyZMZT5fFoeByyHnp7u6LPQLrA/DwuHkNC6ygxcfm94zRSEjeSmyr1PIi
XCmw+HUg5QpWMTQyC5d7PSmasRZAAEurDiKuEbCkpHD+P1XSTkK8Af6D20niOUXk
1G01QbxJ6e6iQn3+OhiHgpLk/42ppmvsAWHW/Hvkh1FbVsOQMNuMBa68z3otxsuk
IO/i1yjewW1fxziPKeyzMLjVj80D743gf6CIjT0yNmmccH8VimCu13DCohfj2w6k
dWVRkdeSkANNhPwpUaSxMYEVa9EZclxOrZyLMQ9BF9XHHGBo/i539KHSE4uWy/OQ
z5cedWMDA/OG5xm95B6L2kI7hAjv4oZgNSPA82CCxLnclqa8VHX7ZWljw14OqPTw
gu7VQErC5F1npcmilskUwzraNLsc2O98DBvFAg+9zyr+cd8Urv13avxMHpRBBNMd
RTGRNquPe3heh0q/eXkqPMA3YeomuwydsFPqvmYKokw9r2WAwk8W4MBYuG0WHOk6
3SwVivXoXP9T+fvTnJlalq+SZDXWN6yI7Tc5QVO9GYwpFEK32X6/OX2Mw4EibEg0
Q96sP5+HHr0HixA/ZmmPjNqEcOzFcnwv3z7psP7ei2kLFG9TLawdCvF+6HovCqCe
9fQaeTP7J8cbE8h6uTFLP4k+2vj1p6bZr40Kw7+dRW2i/6B0V6NEWht55Ppn/jQ+
YVIOoyD3/Sf89ie18jQfqb9BcD7VPoh/FWFJmAMT67aYi89JbvaGjtAraRg0skMh
rliIIjU+FSNjwBuX64jRBmZ7wSXI6zEp1agsUv4/J4kKG7alriq8kMEHN/SVsnbq
wX3tqL6uAnw0NbUFFBSLT8ui+FB8Zl5GWrcyY8padbX5cyKZDtX1+MocjEGZ5bAV
4JcpeHjQs6tnU7qFwrRClbhu+Ue+4K1HunwsJqITTVSyLefE+gb7oqkBWRLl04He
oFa+u40rez2mQCFuKYhjB3ydzIR9pQdDmEI576D3LSDwBOjOdYEHgV4mbxW84eaq
oajydnleOfv6e49JivSOCIKj65OIy9XACglIKQ01mN5QYar3lkGaearLCOCNarFc
SjpFPHQIFS5OVFTxNsyuepAZrzxgu0IcUmoj0q4oFP3kig4MvbxGmxvyny8gfVb6
bepdoU+xh6rLAzHRYb2LQiF9Qowbhw7mAXprk3mEb0msZtvp3Kpyo+ofUnOxxokr
0r0nKBRi2++gak5HqOIpslPSSkTyuTkt8THhr+kgVLMCd31Qa3Ly78MhqvjONHbU
0g/G48CT6xtwi1+HrntE4ihGCnK3JZ6QLUuwvcMIc7pzrUwD0zy2HPV65F7KJOPK
fKTIuzMrnMsHFRpMGRj1HxdbOMY0Kdejz0iJQuVTRs6xqdanaaXnw5mOReZh4c6N
ytnCxTKl+Hh59UZLyGZKZVB9tKTutvLKEG4o3DT2JpRd+v0pJYiEhGbh4TEtH9/d
shgkAzaXEi+yLDmYKcojCNKGdfsv5eX++xG27y/b/xRG9GTqzVx7wlmR+3uyjEY2
6hh9xd3eFSPN/V6RuoJXDpJbFKu/Ad9XB4cPuE0ZC5m7V/LLyUyFP3A2khyVyu6z
Y8Yi4b1X43pewwvqsIs8K9DhotE1yFkV8LgL4EJwm2Bb0iiW2M5HjdbYCEAdspOJ
Vy0jb3TJWv3ipPRt1GIrc/VgMMU68tT7EMUYtKVf+1/D2q/g1nPuXJRub6VPL7ot
LgpFm3g+6KSZJZL+xzogdtVqzDe/nsFXyPY9Up1mLBocIqZomu0aC1UrCMuPw9tn
CaveTozAVVbxq488BchgD9QYygNu3jc9pBLsSnlWCBVsUDEkRWfRNFFAwobmCmDR
iBL/VqPBQpyoIHkprq3FcTaGNONN470omBclHQKAFTt2cuX0xTwfEnmERqD/n3ZO
umh8H2QV6n6CQ0R37x0o2gGSrf+H/BrNrZIyEJJY8T/fz4VPWrUyaNtRVqH12Qt6
QfgkQq1kiqc0XVaOaAL0FV3k2aaU/6+282kibEpMN05MVzsgSsOWkHMGjIZDasRd
qtfLFLgEdTYTtB9J/SPGLdLX+kYkhY5fPuFYMAWI9i83kTfA7d13dDVypA8vbcRB
5T1YoZ69vvAHPAhfibyz0///a7AH/d3zMxpm9j+elvtb0gKCiW4WrPVt5EqTPlar
gI73nD5yY4q41wAqB5DP9S8/6mCBcqyhnQdJrevihcVTr7MRjzdtdb5DDkSKoaiW
aCD7TBRv/nmkc1cAuh6xvh1M1LPwcsHqO3D3IrGNCmGnn50UHGeW1OCkhenyMxCH
ECJ7NzmDG+TdSF/16N1Oc/LX1cQGDVapJRA6ttGDgQ+17RWAOJ5jnN9/4+QB6Q82
O39G2HPr8WveCulnCMsJGdQIVIhGd/tXjIho+E76HSZpU+JUAGoLj+HdT0YiXMOK
1EDxtKxl/ytiEyFnQ+tEEU4g0gVjI4cLcfD7JhlsVO8W2+gosmr3/DJleB2zdppA
0u5BmhIM7oq9eEctmZXRlLgZnTwnUHAvRBw0zPuxcSP2KBoSG3GogGMXTK7oISRt
MUGv5ldveZ/hst+bKmGhzQq1H/Jjk2P3JSytA8E5C+fXzlIgl+d/TSWZWrCrKdEb
0RarJiG/IEC3aSglOrUOZ7zCj0V8Mb3Os73+WOWcw08oyVzuPitINnbySpJmdZBs
QXDTcBP1LJ+crgyyM3J64CwzZCima6ruRwnHizJl+IXelch3F0iexuh2lXYmFFZu
8f7SnK5dktCaXaiifSAbj0o/dIPopveiDeR+iiT9JzRZm3PHVc3NPC6DFBnCKrwj
AD0C0q89RfpkmTWkJ54vL3nCFLO3NOVTkLJ5FRCAAxzQNrywGDK5+ufR8rUS4Shh
fhHUS0Ad2jpfdhoBarxWkd8rp1FdKb1DnNGTgyidEiykfVqaVnQ+z2x+tYROmxqK
FOEKdM3RxYJVlaoqatBemIfC3VqiSMCUF6TxEbLmAKJfEWD0Ttuy1ZHkwcO087FP
kzfteT5mkEV3J0xOHxEBRnlK0GYV3TYuvMZeFAT6GVIkWBBsMAId55cuZt3pqDTz
z1w9ELuArvBdbKZZIUGZx1AuExiRFMEsPzP55LEKrS1oe+pEO9Cp8dy+Km0h3eCI
RWdNbVrBInOrrnaiwwBO1O2fxu3zfxhMB0ZvTf28XzrqoovhGO5Hpt0q0qxkNB0v
EFnxlMPZSoeM10aCb6Ak+bdcH/g8zfsiP0xMOgaPBOAEtYbfR3fv0UlbJrMMqy6c
qMORZcn98MA4NQVBvlxH/KCvjRTFG/Fens+81Pmxop/CheN3YLLgYWXM3+ctALVR
VrRN1K4HRq9nZfIFbA6Of7kwkYkXr6B9jQHO9ngriVLLoxh0FHrGWHUhYgpkCZWr
l7Mm78h3Avqp/a7VOH70EB0gsvyli2La2P4YyDrjfWIcNNXRGRUeXLvEGw8hRTil
sLyXWpuv9JfyO1M3HUujg5nxrOeKwzzy2fYndGjyLStLNxOqZa28DX+uywURV6dY
H/B8xQIqR0yoCNe8zu6dfaHgmPYJsM9qPEW6RlDp9gR6ehQtUkW55/9iFUuFJmPe
7xg/+RES+Rw99TUFFQmJtaa+HIGLL34h2lTRapypmgkEXuEa6fE1XGeuKbu3UK+A
Jf9pGQjxR3yqEV3o/NzXBW29hhFctHBpYfdpufQU8AzudgVof4B03gUVA9tRrCYE
9pIYXVemjoAuAfW/8IEIb49c+j24D/NcZaWFhWcANjA3X7QexbePrRi5mZBTM7AM
JCStyZvUeqFinObTCDbVXt5tkG1uBoMy24+bdWAsXDQQiuBTBWqEwYqEkpeXJlSV
pVa4/j1eUjRr8EJ1QtKWvxYVI8KJbU8ukqJ/wcraRZlWGpOfSanrZbZg6jgwPElk
qwCZbV7xRW/ncR+ChXqOQ7dfAforNquVo3uiLoZfu3tzcUvBOOtR8sd8GL2vtpls
uJWHmubKqucHBGi5MIKar9FGXdEkF9/jzwML5UBKRRju4277dHWmAElLLXpUlUVm
Zh9fknJZBmwQFRBmVkT0RPvqO4W0sQl2tsGEkpGqez3rtspq2hiaJnjRIak/q6Vp
8WUP7tkD2l5ldjYpI6ROIH2F8tgAOLgotatIqvGY0PCsKeaLNrCm+WSfdK/OZW8N
78aCYSEVEHlQi520NbGghvSf5Gb0lgBLzfuHvzf9tlBpfh9tj5agnJHGhzlwegsL
vZ/KiYP2L9Sm0+y1Bjr3IzvxMC0E5VINxi1+YvuTxNJetm6yF7JAWbjo5++OQvrd
k2XmnVJOWKxR+2Azes/PdM1/BYgtfNn3HXr4VbIodUGqFCysWrPk6x14fDcqAKUC
Wmw0ub8QqUCqNGDK+mU6W1ihsD6mBK+SmSVHeOmJofWGRTcFEJ08xgqPEsCJFyl3
ie2YgMiznK8rDhBdYSChxaD85gUjBETS/NYc9+Q2s+SeBBAkH//xhlls6a3UT+CX
0glivRyZlzQP+FRC04Grr4Vk8l8cSPjqF4zJJ9oVygZoYLpjpVU/ArjDewQDjQOQ
dNqJ4HTakFuLhvPZwqdur243mcVxERqjRea/3b0is7s2vNI7i+zGrbiVTnGqwpz8
sDzT5u2VWUEbHqdFVMj/YZIMW6Q0L0WBKcbT4Ti0X7RmRi7xgDnPHZD3UOwrQj9r
SvADpVjZn1yFne3yU/H5o2dO8zQz76mIcFAp8ns7jlNQ/dVYYdEHU9Py4TGcjLOK
CELWNZM7byvtawZUQN5RIk8XjEuf8L7TJEK7MmZf4z4ZVN9V5p2TQ1ohRiLHPVtl
LN5hbG90z37vOOzEhCkCIcNZCd6OJcJuZOm+zPz6pC7n+Ml+564ZZNok4bWkoqcv
XJdg5Bsc9RUC//Bl5WiXgbgD5eO2D7RIuQ9bP5gDPyl9PkSgoQF7lApcvfm/Ue+t
H+PpE19QvcOc4Bep2R6ywulVf+QGtQuuTv3M5TNIozJ3HyolXpLV++zaPM/rtmHu
43Lotci5MG2TeaVNoptHO7JC1lCyjB2NW4klERIGiU1iWdhCztgDzdvPF+0Tiwc2
IaEM4rrMZ2W4CYXWhNLCAyl46X/1ifZQ7LYQB7LmZih3DE075XgQiPBnP9iJOArO
YbyARC2qVwJ33sDYVanPdT119rCR1dOgSX/JLI/w0V+fLarAyUCBDb+FYIE0+Y+t
3M5ZlEn+GS9AJr5LiOpDsByRxPhNgDLnG1nKd3zBi8WFPnDc9qkMLq1WSIyqXf34
/4RjV29WWAi6X7XuDoZ5SjHWHjHszpnBaLFVTaFj7dfceV6JafpKJQXaUEscc9k/
cMZoGXv9SPN4N/MCOFEfBiw924sijG/6JcuTnNedctoCnyugaMqIE+rkYSlmooUj
pdYCV2zsOMZOh5svkX/8Wp8yl84Jcx3/3bSTeroFYyUCo3F60bE7NjW7rFhcXlEu
hL0QLGtB6YN2trnbeEiDbnRizdHBEIdgiRNi4gAvmT3RQ/PoMf5dWYkXMeMoz2Sx
7dAxqSv0DCsy0/D++eolhTN057jYdx6z2vrXWa5D5d9CWGMffaFrXFS3sEHGUhxc
+qbO3xfHyu6zIBoo94Kc23CZuNyKdvRK1KJuoy3y+OFqyAAio5XecnVoygHKRUok
k6+soMGJREWcGD1D6s6N5X8pWywoY3JFldqdcS/inBQob443URkIDeV4tr2NAM8w
lzLFClOcVwe+sAOOVjwnHLhj6gp0OfDTyR4pwzwhMt1GuKOcbzkT/MyANePXsnKu
z+S7orLUvQOLERSREDjRSwdLeFTCaJvf5AeagNcQSkwnPpaxdqr8Mux8B6uv95SC
tAH1Xi5zJL3rikUUX+Xj8eWB4IqAHDVWqE++i1TiAp5EzsYthdJGuMoTmiN5MYrZ
TcT5+Wyw5pxl9Ppsh7NY7eb+UI3gMhpDt76rdxed/BpbemiJPZ7btJIkEZkNgRv5
7af/kIlyM2zBt381zyTDIcUVh4cvK+YFNlzqWPizjggYwbMVMm7p6MWm+yYLJc2F
sKeToOP6scGFrc3V2z1lbb4rqT0XpCfebuQNLnzcvzyARim1HvrW08lKsb/iKP9e
GJ+5uyEgW1MzUf1RunD2JWw9GyQ3fAozPEEUhq22Rlp+m8mu5vpOjFs9y9+LTX2+
KMIZ32HsRt+46pt/Z+yjuXXaXNji3OYb6tD4semWm1zC3bSuhCOxpZNlKCg4mwqx
Aotbe18YDHtnkbE7CEp0exxm5p91DHQp1mjBpxJ2aKmTw/VObD4OrZEL9+RPNfx4
Q8syeKBEp0TjiYtD4lTNxZkp/mujkq6B/W/T+f8Q+Gbyhh5rXXPOwuYfw8tg176i
AjCGj9+xjADf7g4b2ysdTAMlZxxCPpcXY+JujrT9tGcjFFKYjjcLnjDZLEM15gyP
tPCBcyKAYkLyM607hvryDSH0Tk7NTQ1a9KWjYDUJWx2D0YzWY20odqeHmb4Dz+Uu
tn/jmKlID27MjdUYiBV7MaooY34ixiRpZbXPW3ZqThwmYOM36bd2nAc33GTYncgL
hmnQdP7qpMs4thVzuiu6MbnXPDAvsdtic3iJbc2ArMDA0ca5lMHij9MB0yonWM8A
dubJlAp2Yxobzb+6U83jOaAKhJRQvm95urMKwvFPVIGRTD0dtYPgTXedK5q6BzMe
Z5T6bEc+zhtLtHjVtI6fexmQ7Kt+RSUW0ESy9rCNg8y3U256q5DIRyCxfMNy+d9b
AMMfzSM0pGrRxjlXMTVON+LEdzy+t5KvKDnm6xfsWzAzhe2L+TX8CsRkx61f8PMm
+5SgwsbmA2MGG2Tol1swiWteNcBW30zrT2JVBcaBpqAsXvbqhlh4jtIie40zT46i
vtAoOyUCXpaOC2clPG/nkqxgBJPsCABL6ByLCwE5DnQo34hozdJT8XSq+Ycc3qAS
38AozcY5wjUK+lb05nwPUfpvTzcr2+gSHfYxwybvrqWtQ3gkaHApxtKv8u4LKoG4
+DwdXsoftzgWJoIa/OJbCMaaY9dStNEu4dZEgtTdxRd4D2DMhbpHrtF7Ti/pTwdz
u094IXVCVHgnBVDcRiaBWiQne6rrvVLUeIiKbjWAAXR3+ScNO4DZ5vt5iSi0ig9s
q1fJ3Mr1D28CktRGlZCsVHkxSUW+6iGp6lTCEJRW3aML5haZhoC3PVfm2M0WrUw/
8do+hNaaKk76RzUP69iRZlyrEahxW1ApzIG9b5m8kFvc6S+4PXx2IB75NMSsWv6K
fOnx5JI8U3QRh6J/Ik1350RmK1Rg6EM303BZ1L0q9F5UrkDjcGpVdnGc1MyazM4Y
/Mfheo4xW2EzVMnNVh7qlSCSTuvw6rUjPxf7n4DAJ4KRn6nto1go561fayjR29p2
WOxHRzbetFQEWyptT/rato87zZnONwb0WpM7jhnS8wcEcmlWRBeUBUP0yY+CEr8/
y/cVZ0/LZV4+nvvulfLH4fzLo1SxSx2oXSvd6pq1tOAAAlkaLyAOnehUW73eR/wl
aRKxmNUNsYa9FAXr8m68BUiSDmnQuTktpSi1S0K92gexTXbhcsOmlSqv62uvaTtQ
/rvkqz3nXfgOictF7D7IZ1+Z2uuWyEXgrMqHhhSE0il2BBfAbHQOMAdonpE7i3sJ
82ChgQoBS7gPvauxP6BMUpATFBgc7AYgghSgQCn8zSXRgtFGnyUElLmU4fDWNx4X
zZDkX5ZTqt0oDr3uI7yBVBBW7HpD4LNTMW4x3Du9ljmBYK5Uxx5OO39XtBg4ahlJ
kd29qVCZRVUtskWscuy1Iqz3p5FvZNmUf+og86esUBOWB8Dd3qJQ1guPVfPXy5V0
+GS3Q5etVbZU0Y231hv33OETS7APBTVry8btljwwdcujr2XD1eyJP7S/QULLbzjF
EW+7uxi705QxkQUuSDZvKbxo8E9k3qH4MRKjL/ntIr31fr8He7+vZTd8TDNuVunn
1KO7ftlOaNqS8ltcqlOnEbcezKQ7khXBgMNTaXgfLQlzpC6Tqu+TuwAInYQyOyG4
rlzURCmo+JThQm/oJ/MBwtEovibZRbE3eja/+rvKZ5tOU/HZK+BQCF+78lpCc/OW
QZ/JsntCwIjSb5r9c8XcCe3qZFGsATnTRzWkVEHwnQ8B0Me+tw2sWBxDMtdyN0wB
ayR2ZqaA2M9fTaa4Iz/xROBFDxE713wCZvPWT7R+PWEIjnzFxygP5EbviBk1Oew6
2aUdaKSV2FtBCt1kPkQMl7416F13bu70dUybSs+cjYdIzCkZZfbMcETaZDhWalpb
EHGpv/UBuG7lmC0K/7BWchV/GLg4zUS6YyoHFoLmOyNonsG50iMTX7pSQr0SFTbx
4lYTZ0uqkMjq3pBtJTow/FQAbKbgW4x9BJHx6IeAekiHC9F5bAiXgBUk5Y7kzlLO
4LD8KpcWw4oVdv1IrWfiKUssBOBPvTBRlKicALrMQc+7lIizzg0rL3/OckvDqZkI
+MEIA3IZqLxF8qiyVy0LRTbfwJaSBIfhdEhzANMAnCtm/mBELYhwdEiRs623wspH
4W3HgL62Ze6azu5aqDWght96SGoFzMghjatJiVU3I3+yreiLHGy8x2aGvzxfVGK3
KWOz9//1Wwfvg0ddpVoA7LeHJFSvFD2+bnkG/CAZLCDwnYONykHVTCgKKGbgrcSu
QtlbIpW6mNkqcWt0rosIPh3ZR2teV3G4H5KUzRSrn1MlECAiasn+S0Vvk3JRKgMI
PhZG3+wLEOZCqLEL0LmUW0WXOOvwXqdOZxvofduu3A2syzi2Xa+VzSjbasvrCEcw
3PnLvb6csVr5XSp7C29T4P7hYYSR7zR098AEDkimIwaQ02fg+TF0tFFmICkoD3JS
i9anEE5WYsuj1sc4X2W0ODfBwnexwXspG+wQgOElPltBK0iIEcfYlJALyA1F84EB
gzEpI0pqke8lzhD55+GmQxWLVkbpTPlUOOKOwyiS7TOi9hszq9aARV8+YvLazJDL
vouN9rAQiVCtbtXKNuPN+MvoQkA/Vm2scAjmL9N4qElqrJ1xul7+l9ecLT8wvIvW
9/1K1OhXrHkSo5qLqM069+f9BmZxsEH+P7Yba0OtSCLZEJyPrCNzZOFImFwqxppj
g8w95Hz167DOCXt9/RICKPhdi9jOx2qoFL1AZ/ra8klpmo3V47jRLpsDTW9sKk+V
0YBB+/p7nT31z4wUZejsHXn60iiM+6/DUYpm1cVZnPpIF/0RGhnXO2f+al+XcCtb
V83zypLTcTEv9yrK3FAhyHlDIUfKWKEWmnMCoEakU2usIwQrkc42ZSVU96U7GLyp
MZydUtyfkb2U74EnPteQHmnnCBPiIBZ3FIpEjre2TsLd7KFPsxoAXU6oyHxit6j4
A3PqyIc2dCW5baXms6mTb55Iu2JGW9wcW4xebUGfjHEGd4r7tyq3y7jnq7lNC81F
AfLWSd0vh+TAvdUUTwitBbF9KHfNqEw7tT/YFELd9JUxskKqYg3Wuy7DU7kyiMYf
1RCLh6GdHcrxxrh5pwaupI+M7hOdKHpNPoCOa7BsfokzaIPFQgAXa51FRA0pXp6L
oWoAwPw7VazwLGTRzHdm6HGxgUi1JTSV1O5wQk8ihkv9g3iWYyH5q3I2QodKG757
jtA9rH8cg81948zsaq9pax9viaeiTw2XafB6i/IUCx41S1H5hKJoA42k9wKPz26e
AzoTNDq88RrdInZWDEV62pftj8dFmDEMIjDVDGwkOKiciNcy57lCxGDCQF6NiF+Y
pa3/AcdjNz37jZfV2PcCdSETjPXjsnYCZ1Wm5fwp80XVs95Uj0ibwDbhxH5t2fPL
GpKvcvjtD239Danqs7pc7RE6EH8L1n+KpYn2qIBmd8ogeG6klp5Hbqqs6L/ODgCK
7HHTMUpZzMABGJibz2GorWwhwa7PPMEm3gbijJDz7cY8iV1AkO5E2Ay0oLjeWJ66
pQ8xCK4pPs+CG0obQUUCIoMWKrM7fPlbyqGzR3rKWtPaF0m/EpCRWxJ79CaXDDY7
Z45QlitqCvcYONvZ2QEYvtu/PrwFvpYRLNdE4lssEIfnN8x2OOLt1Q9tSpWCP805
jAUn7CU4Mh9+zbMDZef4eotS0a6TCh8lDjl7Wlxf5358Mx6JsaZcAQxFk13F0+nk
9QfVaZBf/Ak+H8X8J9J71xBbC1G8makx52WR2pYj7JIGA1ILF5axOaZCpzgYpPmF
fTkqQN61ERaM2oguIKptK7HQUBCu0Yu3187ksnuuz+/PuShKLmoYCIFjGwy/XsZA
5TIeunMq2XcseOYB0i2Wc09DvLnQrshjmR7TwSPOnNRlPUKNTDbMfheD/36As2lY
OIRG6WXU9ndfVRz+nxzY80DNgk9oVIvHLmEISEms7TN3dwVGZrZQQW04U20TQRe0
IQFpCZ/yR66rkHP8t4/Qcj+6kj/Hbnd8niACPBK7L90Wq5u9SxtJd7RC3tLRqGGR
mmJyUZgEmznBk9Ue030Ubs06j0PkSCuCxgmNJObUJiowE1UYdZVqvcELv1/AXKHT
pcG/4Vkb5z9dKk0Uz/348bq+PC0VPa5EfVpqrJAcoFYeK4HT2os55SePbFDHa9Km
QsAXHUzZ921aNNodwnGGW4BgME5j7X9T0fhgILOL4nkd5Rp6xtPbd2+9AwR/IdTN
jidoLLratVLkgGQawK5rLvaSs60ho3aufQ6FjHL5Am2ZhHrhxKN7EXczs6i6+bfp
Zvpy76MDBeqoUY/wezQYrCJ6cg56zfShjcB2lrJlUmINLLJW7O4LN1GpR8+DfKHW
cHqY6zNsuhomRazzQJHdowQKqc5W3QDSsbtKLhXKwAlccXwXs2qJI6MXA9rxyHAX
HVBDwOL070E2FQEWZnsbel+zIg/7oqjanGOO/x0lScpWPmZbq1ENOSanbDt1RTOT
DreZO+BsfSgEpNad0kXbH5gKCwSa1Pbezkda+fMTScOqoT8vy3cS2dNjKuTCzZE5
9X68+KZO2S2fHQt+eTWIj6t/DNAjFhxR+BP9fRMbm3QhipKiZWJRy3F4sysqAZFI
6Yq3bqh46vWv2wb13uawJI9mIcgJCNBHB2h8oVjPTy9pGcr200i0lCmEw+Qdpofn
0zyA8CEkpy/cP2meJjy++1tCeSdbHrtlwaZcdtZ25RG74Q+2QEhK1dNotWjae1fI
9499C811TkZp9mxKVN1GmHQ1wdOxhqE2eqBKUa65PpM7EhVqp/1EzwsIJ5ZBSyWy
NNZSy1GZ8K+WA2OuUES5z3sqC9/B5uKCjOIjbZpoS35viEMvzdbfrjDgRF0J8Jth
r191hgV9ZNWaaXARfLlUnznNh7uaOh2fji5UwWQadmh5NQRlHp/i/NZYJLC3BzYs
o61QppDDcNptG/jAMY9U7fRpkm2PLEgd37QHSLr0076C4a2y4YgmEJVVp8gl5zYQ
F+TZhNJs126xpsQzf8ZaW1xNqt7NdtFuhLOkbvzr/+2xOGyoHpiyBoX2aI7BYyrW
xt/HdfRWOaIOUfnFqBxdfq/deaSwSTY7kQfTLe5S3YQU0yig4VO4q722TxUo1fnt
TMuJ8fRX51oxzryRxF4IrkoI8pvJUcOFLRxK8VYRX5f3qYKwJ7PlGO/VKiSC/vnH
M5OTBI8ZZxNHRd0b7pbjPsQwORVszMkM2O55PIGNJuMh+fZTbxENLT4VUV0Zs45o
tFRFNL15v+KIovggqny7dn+QZC4yD1rLhuDWRr8t9qm6ggBkyRZTPJlBVDRgdldR
A7gHs6vuGI2TpYSP3wa6VFjndtL/ZZocP8kcGiQajunnHBjYC/AgVklBM3yCH4lV
h3RWJA0iH2Qnw0R2HA1YYFo44Ly5FC9fFg6RqDTiKOrabXjcmjzm4+aBeMwzsnkW
9vTMa/UwC+maCicO27eQ75+H6L9ip+nOjJReL9vrGJm4VjQwTViHNUj1Kr1XNDmn
QDqMsL5nyY6Cp4lPwfHWPWISUXtXufNgrAoeDJJWXwLl69UBWbMsrg6jeNUeHVp3
A89Bf+wS8PlF+qvuLGwHuomjUBCWYATTHhCK4NGBjzn9Fglt1y3tWcPTO08sANWA
zW7Baao9Im6CaQ41Lpa4lvsppxyYfO9z2pfYLAK9QSJq8Jem6mJIV6CBtMKOA9lb
DUUYU5tPe4WQ0I/QQ0nl2Z8US2fiWJz8KtWmzIiqB4FmHnj7lB800CnUU1DbAxwS
JK1aooai8sWfRgDjltFYJFSyGI0bT7PQ6RW32TVRyBfUDKWNDFkWXO3WuGEX8uPC
KLoAhQCoCIT0b9246+kg3g1ui5wggEcHocCTSrG9eB8HJMb6BgeCiqdcGh2bmi+z
CyLq+jr437Q/Nh+eUTzMwF40bhL2Caeb9Iq1kqWAp+pZJXCKhy9N4I8tmXcfZ2NP
8GjFc/m1YT02tMGRGoCjrS81LKJRIakUoYk435UHpaHuRynqwkVc4fUnbxp3jVvG
eCFSY7bshvnUIAXeiMPlHM074Y5GXeM2GohPsDhC5dkgTxdeTYeA634NTEEsfocH
xuB2Rvz2CaK5j/AdhqKZAWgzJJeFIEdHwI/dmmRVFhpCYF9bKKzcl45/tXg+dn+2
ow7uUHVwld2y1FU8k1+DMZB5JqAynS49VfXm6qYPKMmuVeAMTJgcmc6qBHB9Ofdh
5184I2cEo7TOsLo323qjdDuf9m8OYpI/tZdoq9m6U006PoDkDGjRZafEae5et/1t
XmRoooOgR/PnmqN68YKxkO2FaUvlCV6NyKY1CU74IVSzcCTpAcudz9rdZN9SP6sE
UIva61VAd8cPRzapTNvSathxAw/8jFlCHBmW+Mhnh8ZJKEfGStX648E0EXgEoX6q
rqdP6b08Bhff/EwnYIcWGpTH85OZaxl0+x+IEcgudHhD7Oh4eBHumozG7jDAiAxM
9yDJXgmLiI9iN3C/DRTkp9Lr7XpyhkQOMxTye7CJ2sXcIlQkBUgjlfF7bOgqIN2q
p2Cy622w2st0Y1QwQ+RYPb34ensf8UHrabk1oZCLI+u2mbx3TeD3pzufZh/HniVa
QP4QXp5n032HwJH8ODIEcuO9wZjSCHi2trT7yoN0O3GYczwQAI9W04flEY+h4Dff
TzgHgsTcpeLo017TrXufbkl4AuQUYhAo2bdQwhQwNACyvzsAywtU5nYjxEhQW8UR
p5CbBVV0QZdKfZB/ewQqjgnjALWZxJ6aNnbLOxFLRNw5vmLM7X5Z6jjxMdb5Ja58
jXr69VHUErX058/Eyie638oCgG5d9FHWVIFi2ssfWVdbLSOkPjTrJD7rq4pQdO8z
8oUNnq8IkM/ECtlLo0PVv+fK11cP4oJwepL708LSqnwRMf+4ikQt4KZtHG08X3rm
TGfxAN1iFUzdofAWeXbjtYdwRUZz2kx9SQf6osd6sUHbjoMdVCdpg96xwIvZB7x4
kuU5wTAYUDikMvJwHkozkjP9EgxDL3A4Y25imDasxAsHuXEaJMGp1fRaixJDLa1Z
zfddWSR6JI91PSohwSAo89vHhMGYNZqhyqBW2vRAIEPmGGcQE1KM4xYTH8wMz3Pw
MBM+p8emMNC4l2FPy9UIO5c/IOVJ6yrYA6QzQkxlfcYtm6v9UUc5ANVdCeW6a7Hy
msuvHP/oFtJkWyx0yM1Cgmbq/z6eDKKWYunwDmcApZ+3hwUcdANl0lgvx2CC34E/
0lNwTjOZqR8mba710kD+N+EelI2mQTKp1/aOkzPo9ybmpoKo4ODHowLJQzNjhQK3
/ACs6/cWH47QcLSE3anmm+1XVvdInonKkF9DQWdmxUF1DiNccw6LgZj7P6SG2ZNH
huNq54pe8JaifydtjFpZiMx9fXxWpffNDNFjvffXAwK4O/J1DGqYYvwtQQ8UqBZ6
2c6LlergV8PAMiIIgREzqSg5S8eqssikxmTz2o6q5P3GA3TPvWhQQkMdp2Vtu1k3
ZEILRmhscE2V5vqf8AdMN5JQeRVUNP+XgMLFkSIExIsk3G4hKp544CZl5CNRIiaQ
4YKMfV75BhYDOPFCm12AE78k7dg2eNHY0yJUET2xLPEHJSqaC8s6FQNeJ1UY5wdB
TYakL7a4Yvq8ALGnB266vPdHeQeRnL9jQ8MzqBmL6VqmL8fzlT5Sf6m4D6SknXuf
lIS112k7vmjXHqrCohOWVN+w6MN0WNHMangKFIq36opsjnGfHzEutZqL10ZQmLx1
EdyRq4cho+eFhKGeMNVu1vWGQbTC9lLpSrxeWsc1OyWr136scrZC2D0oPmppqu9F
GEEprPzgbAYbpPwfKND5iVjpz3vy86PYgGGIeQ7EfoJzWPCf0GE4RUj4InEm5B1V
6Zb2vk4MQ1ZEygTR22C0ote1L6uN0E6n3sy6I/hhFDXVG2c1OY/xTJYGfTcIQXTB
+T5PW/cC9PL9OZSZnXXIn74X02UutzAJg3A0JPIydqB9Vski+hzd5+SPwY9lEpHy
4z+kXfJcDMCClQLxV4mgBYPB/W0BySLODY2VqQm+lt6AX9AjihlCAcKNTpPoVG92
PE6j00nNm4WNTrhEixw++4bAa0B4L3bUcY/GZkXA2Lo/NJqxXqbgRsYcCY8adB8W
dbdMTwzPugfv0nBLYED+uYpa6JA++s7EwMkzeBiq5i5v33A9dioQCe1JHnuZmyig
59fzlgR1qxX5SnBR3G/EzPQEXIuj166tRPGfKETwuMvDeMYlz/iFHHxM74qaiaJJ
HD+zyYlEzNuOGP0l6Gu94/X7K0NvrlgXK0zPw9vzkqjR6vjmLLuIfxMw5AwZLLhc
/pHjUvTTsuadLFRuMvpuq52PQnR/fT1kbcuzGu4H2C4Y7BlmmamWqNse9cXIuM0I
IIFims9l/5IXC5bBLlijKGhGq+9B2TBU1WYo5kbf8HtpTuyUIvaOj0bRo2EmQQ4x
Ox/8cIFy0UePFg0+jzswpOGhdWM5N0vHm253sAVhEh5QJmBQ3Qe60/a0kvk2xMVH
Y/dcCn/QdJ44n4SP2ZO23l09DHbmkWNhYNWmpaOQutgHZo48qGsHuOagGDogaEX4
G9Zdr+dLrhQY4g1bsGTBn1fit7zqnH93TKInIkcoTnYC2DhfcUy9VuM8+mwNbr/c
pWtBmxasbVpDTJJEa+vUjLXfLxDSUQWZWOGcUGtx80jLMdUPA8+qRmmYOX4dggtF
n70VwZkN9tB/l9xprgCl0brwdyaWZrzKISzCAjrudAulQN3q4t1dBDbANaD7pydo
rofXSRVjKSd6ZL7uS2JhMU7hPHIsr7UTf90CzfYmMyY6uLmSOn44w9XvWIMH8TbO
7gq4AiLjvOiiIqVKAvzDZyMXkq6plSLub0xjLNXEX6Mql/rHYtjNcrUzVgidgoyi
/rQGWJjyrVtoc+f3JivWle58LGZgZWUPnTTg1x9ektoLQYbSUdSDPa32JcKSoJKw
qrmpcqYJOqUcNNSCnwNSjBPtFR79DdGzr83/4mn//JHpDYCX5THbibVWA5fHpByn
xFt0L+dMPkgWA3KW1SMuTSqKkJQ0OemNyT+At+ILl470sRL8vQ1s42H8uEY0we8l
QIJySrtq0KAtPh9LJ5jOXz0xx/m0TsA8jNY9QsdH3yt/DRZEiQWZ8RFBvRQbc6ZW
exA8RrIgGh02eTr5bIG2YAIyFcHX/5IbSU6y4d59o4eVu16VF57PywuWzUFg6AKt
eW5gPo20q/3sxpJrtK/sdcUHeGjbInaEk+hDpFLjmObN6sHrM8KomBFDruaJxDWd
ULh11wAojFrkuACZKmXWVuoKORSnbvds3IL0JVvBr9LOgsfon7KkoTzJ1Fclfmd9
lTK0BiiLJx4jhuKoGxpFoOhpszAvH41y6KzbOXWgRxWSJzx+klO0rJiF4nhRE/w2
aTyinIRLOFTvNSrKslh+jwPQIg/oQ8D6nwJu7sk41QDvXOHJRpiD6VHNEIQ+L/wR
4kraNN1hDzS8jb+XL/vrPf4Myn21srKMaLtPVhm8AeGsYeDvGPd9RXlSQguVfuo2
4ae13ua45T81BZbwFdOVrWIUn9dtwuBbycGtJghBsg+d1F0VmUfBSG1xj08jEveM
JHjPF0yxODFJBwN9atc3IQ9cQVAn13TZnHZa1Mh5588JL/7vjjN4Zn9aZFBM+02F
+pu8rsdQI4CzsBU++4Y7xsTfUH+T8Yyn/8/a24BzDTVEMSeAfr1G89vPbBQpku/2
nJYfLl4sBK9uvJKShjq9VPKT8QZ7cOrX6ptVkr+CoZn7oUYWyYCCdXnySebagCOy
KkvItcRyizMvdlmN0gT56fb7beXidLtmJmfahGyRT/j7n/vj8YBfWDpaTn3gVT/z
accQlA3iyt4GPFpXABnSp99nES1oDRKX67UW8EXZ3Z5ROdi/2BRbX7/98Q7sCMqV
V8Y0oexky/yV6RWBExg830kQy/Y0Tn0HDogcjisF3Hpu70LKMpNAp2ICX9d5h8yX
8czLrc3ttI9Hcgd+PavCS+dBLlsgCY1Lee00NarKGTjZFRc4s4Yx9DaaemPbcOpN
eBENisbD0dBUKmMaVn9Zal645SO5GIKk9SCMCXic1eizHkaAsYCay+2TFvzpC9tR
ShuPDCX5RslVy4mwcYCPzVwxNizU4+jHS6eWSIqh34Myj7bn8Svi1gtbUQVo+Pd+
8QWKrc2st4v6sIrdu8zrSJaLS7OHJC+tZnJUq0zunMvTKu7ErrRl0NnSE7K9ZT49
snzd1EwP5quVSaCNMAh8mSgA2pNynYrUVxTxPAl+k7ZWA791XdLmfoHDTCsFoZjO
Am14k1UOl7jJnaAX2OWZKMgPhwuxciFwml21+IxQpi8w03r1lfY9ZqRE49MQ6xCM
/MPgTS1zE9juECrbN7ZIDBFDWwLrehP3QG0PgJBrQs+nD86meOisjYxVAIBX3MiR
KKgy1s7Wf8niS9aG1G6EXmJ5u2z6+FOdSdrSQ9t24oEs2RLB33RXUC/ALjkKCqOE
WfW/C4j6Nd92szbRsUbVvwrcNz8f48fn4RHHmoP/U6PYvf7x3cq2cepaf6yqmVSR
bfH43pVAqKqpOA9+/5ihLvkjQQzcje1KNsD1davRJvyI94zwmIsIp9lu8bmJgTtL
b3Tc4SxpRsCiT+q8Hu3ZdL4VFv3i+Qb/3Am6hCFtmyY9MlZGQNlGi0s1jLVJiNwd
muvJvXoVGWBta2VQNEjNAnoHEhF8KY4nNR+FqUe1q2oWO+mkz0DW+OYHniBzNqq7
O+Yhrcx5ceseSfspwvsoEltp6wfQ9hpjPnlznyTC+2JcQJ42Loryrmcg11auPL7g
sB/MBCrOd5FWklGk5UIzNKzGLAH7ghdxDLNnYDV24HbQ5FjLwFUQxV6VcQdsogOt
Z/O+SjauPyhfVo6wTw2hT8R26M6JeHPXIqF0Es5ZoRPaYyvRfRvhzIhnLYDWh5DP
96kaj9JWO3Gs6DpDvfiyT68tf7yLoK9P0j0sGme/DOPNxeuQjpivzK8GSO2v9vmn
5+FArq/38JcemN11YiDlBxFVUKs2Q39E88Tol7FPCXXM3h0dnuHELeF+QJIiY/ky
zsCRNQTWISLCNKR6Atz+ilpmhBLu227CkD0UUIY3yHrhglXTGrjSvrwGdZ2LQ6JV
1eh4ljc/EKgu5WaLucWjiibBLidoxnykuECGosgfw+RxmpUts85bjWHSvdi2Fhij
xhsgWrCaIugGGqVPo+o++PhJ4jgUef4my5Nt6aFFB0ajp58tfso4Ny6uHR0rJMeT
Va7i6lauE46NXdJ1582O4havR8ONJUj53lrQCcJHQ5idNzxS7nBgVmEh9W2jwdWp
mf5KXuN70v3cKBv6tIaKQAkZveND4BFjz1ENZBifG5yc5eQQK56ZOaF6WW9C9Omd
eAptwSdVQwn3VNXO8CkbcpG3YXURLBv4X74VDKCOScHo3eMN3nwGp4JEOBhw6dVN
F7vMyyLV1FF2tYnFyegd3N0EqTUiqUcudS8wdMMIUssrKTiSb9qCEpD0sSoVXvqZ
T6Sq+6sTrDpMGqYtycnhFC1ML0oUiO3Krn5DbmAAkS+L1w6dCPSlYUdDRX62xKjl
r9KgKkp2l5TbLmAiIDEo4jl2shfmHGiskAcSpo4+NRud41yFhDTTdqnXm0C+fwEv
nVqsipWIhCFklRGURA7j2hobmZaftJrhnt6SKKuhhMW2umC/6zmRF+YH0hwEG4L0
cGQknmKUVG7shuwr02MBZxQtvLvaTYUF+wmUobdJrYmzjpru2U1TG15SsDgFuaOZ
lQWkGNO+x/KoQKOhyPUCy6+sJIKs2E6XQINxaBhNmjhzIrcQ6voWSwb5ll0yu94z
9FpP1YIE+ZqEtXLoqE+cKAWVejeOKvchtiQfPI9ibIpGycX/iT0/kKMrA7YySVQM
7vs7Pd4jK2hGwzY7WiFNx2hbkaxSb2qHfumPPu0pDW5Yh13+dmt3oWTbYVKkdq2T
rghEBn7C50N67R4GmQ3a7Q9DVQBMYvJhLf9XqnQo7zPScb4fzGaXV7k0EYe2Mw9P
26Pt7CPezMXhi8wOVXFq4O5o6foh8poqJfM/munlkJILoG5RE8LhHHR51tQ1Tqqh
LVt/D619eyHqkxQ1b8M2kU2jjSGjFmd6qWCPIRSGvPUnP/ow0UAh1hY1DlslSsPs
SHPfs3BR5qJyNDljiCmwoMUqDmRRix2wFnph7/AbC8iW6WJO8qD7gHGTRFP8aI2+
Pg/hgxGabA1HY6ADxgxNTnxNxhRpw6bZhlgwCiPYw8MroWa58NHWaM8gzsiFwuDZ
H94rpP5vvB7L7nYQV9BJiJDtAWuHaDWB9eGaYze5XFBI29JYxYmbzl70Ccgvw/SM
Y6Ksn1nV+DPqN8F+Mba3QHFcCZEbCRUZJeO+WKyLZuWgh2eh+YEqxx0ffq495rls
XxetNY+ii7zRcjgXLJ8Sbb4vw0JeO1WIkvyXEpn6tvZ+anUMxBHOQkgxTVcWYVgo
2eaSg2fCz53JgYGYsVUA9beZU9vsIuFmGtcXFru/Acr/Ii438kZillsvb7FF32Li
oa7b6DfYDxoPvQfq9JjvZgO3dnU8k8HF3NnMDCNv3ZzWB5pFIcCwH+jL/pAWYZyp
MmZoVzKQyESXMpB/PfGyusVRSN7oFwpDVUG25SOX0w/o6+srXtVdwNtBXDgLzDws
RFlZ/K7/qWtOkZdO+YzuSBtPbSvb9bzwrkUjUv5UQtF9LLCWb9ZkBVxE/bPWHfnH
cXbRtlz2voODYdnEhxYh6Jt/TAI4nvkVsp+AUxizt6jvgQx08CLjAayv+0QImmVk
pvE6+lXF3+4E3FzbQfJ2c4KHOvlEQlpruaLzYZEKN20FEU9eL9+TkLsg9Aew90Rn
eIq/wIgClOL+/zJ+R3W03u/v+YEOp8V2SibdIInCT21ASTxQjM8iIl/2yKl/BnOD
kCIJWQRT4GKgAjAahzYEdS+aIZdV3pQl/TT9KBK518CphyHSDiecp/spdWsko3Sg
bpMz6WA7VGmwR33v6CFSbD0m5nhLkFrz6ObkQwYJBr249uJW0CzTHPDcw7WBwl/H
+HxFDKlTJEbPQ1CLChnn/Uk0QO3B24j6urqgKPBMzkNXldIs/ig0EKgkZjDqwHKc
tqXOXsu/cGZsNM8my/9sEzX3pB2Uk6Rc68jinik0INPaGIh6cZngqeww2bXPMlUt
vVGMJhWmvtco7yBJK7s7hclJI3O66mmX1ozNTucD7IkNnoHSrD1tBOLNnYVqQvLM
X6GXZs9gvXyeiBnXmK23t6/o4102TyOsKriFAd+aTCPkRajMLj52XI2eKLVVnV0H
i5ryR+J2wecb/AdtgczYtxYHflogS4BXqGznedr5nFkECGpM61CkO3eXGfZqawwK
zZ9bsDqDHHZkM2PfXJviHcPJlrrhasES31NZZAE9T9nQ/uZIB9Qrnjkojnyt8Ljp
EL1UIYrV7DVOH2ukOee3ujceKZ385e7byayEgreGiMNARQTIzG1dyaLZBVyUsUbO
mrkpn1h6LxwN+/eQiA+YKR2BeVkeu5x9G83vzjtrUb3Q/ijx5QYdD6UGt3s3Wxtj
Ir5hCkrj/AVnFYZEyOYV/GUB/MEnH8pOxBLevZFU1BMY/qlxtBH4pU2zP9ywObxE
O4GFZygHXigPTbyaQhLk2vFQgbMe7WxzKGJU2HXUTln2Jm3gCu1QNJlat4NqIaap
mHiZE17l0BUf5DLYs8+CEn4qIV7J2EfRIg41vctcpum8To7w7AzjxBIb+yQMXIXs
NLZSkVKIN76+wKnj5daHVsMTfryElK2urp3UVQ505D0PSRjuxMDn+5w/r0yMyyaj
jUgs4kcsElTenM7J4eeEhLA7Y4+DpyUYc30a3EqPBn/X5HbFepU4KJDbQnffLChh
sXq7KwAeNFhzk10UlLTrUq814XoD9jC0mf11NZnnHmVVTzE+8ELykQ0rTkgbyBSj
zwyfO+rIb61G1G+YqPZqikJDkxZucc3V5QnP+j1gEFF/S7B5kwUvs7A2JvhhqkyC
+Lv4rRmE8FIUKNpz7RC/jJZidNm+Xp2bExVGO0Ec1kEyDs4Vo+qwiYf6dLaZEWug
xvQdfMQcx07SJlxS3gwPxuQGwvg8JKXn3fDTnXpLpmC5HFuCuYSmzzYdruZmUteu
WdRo4L361SZKI68arExzodVASnFU6FPqlMPYa4nH261Glfc2/kODrLHZXG5kossJ
RjhaMAosBeG2dLpTFXSyIWTgeK2GXauPX4cNwUWqJ/zmFt/wx1jqcF3uWrh5iMXN
FP/S3tghp5J3a5RM9fkpHXn3Sx1uVrg/TtMqAZGlySA8UgOAK++Kzg6XApf3CZht
7hdxkbHFySjAbQvrh8PuKa67ZOOBhXcej9qpU0c4FRL02os5W4jxvVtk/fMPep3N
jkoR36XN53T4e02AF9PdZINXBwmY7/7T/PBhUqFY9Otsdqj6ZO2Thbh5EFVoMYB7
jwrUsgN5FuEU8XOXl4XKuO8pzOR4wQ0JAyuStyruXfQ/yXDkQi0uOIUmEpLiiYw7
PiioHG/RgyOlbBXrF7sHuxqerh+OxIe/a6mY26UMv010jedRGaXqv3GAiAIkW9rG
7RJuqkWh+ZgegHLCDh3L3usBEu+sPBqLrmsQECHxIaEb0xvVqTtx/Glw8Gc1ShLw
vZuLJj9rSg2uynHafD7PRgSSnwo0S+5EHwjK8g60znmurKc3Jn+W4xv0w29XXoJI
waGBH6UOk8d1NsSBi7XM5erfgvD60Yo+2uuNLXZdnXO7tZkAIQTqkiFyXXw3N4+n
s7NcBqawjepG4lC0E90PxCyNes0Ex6I1YSoEq0Zs1IVgy23OtvF7nw/HU7HYZ/Ob
vUZT7X9cQ2HaTzieKaq7FJWT82nFtgO7oHLk/JzEoVh7cT3wt8jGam4Wzet0hzHn
QN5uxf4GIXZ+VoUuD+YS0sBG48qSsh3nmVEM2Du7kUXmPxLEjS925kFan3psUTVm
9t9dxX6ow1cLIU3we7C/yiV5yBbq8QUSovdumh4aX0YyDylfBXmcTd0gYPWzIvCD
BjwO9EY+Pot9MLZqvvh7FKtgTytSC0k86EgvmIKzhs5icp1qXhwHRov+dFcom8EA
cArBHI2avLpaCE1XSigTpujf/DnkzeptzylvBZKC07ZIg8f+qVTrqrKBYOIGNxXT
RU7mOhDaeasTyfnV9CufOoEyTOQkj/fiU0BIyGsSiJfa1vhzYDG53LsI+qdvCfrS
DBv3433d4IoIpPHqqx3fzDUQBp6St/t7PAotEtriOtiKot34+MKz02ksZ6S9OSas
JZyeGYffGtX5UHNlxdibUrayZYskfRCex24dCTYGn/dpddwONpXlI9Sk1S9vpDth
+ERufje9SeKSqsvvSFaYAofY0a7vb3/YjEaW2RzjweGTZCLvK4OpA3Sro9FhvCmX
VwBFK+wciC0zBP+kf/rRSMLlumLbzUYIW2cH9cdAsxMOyXpdg4RXJekItVV1NAZ0
HU6l6pTuLJGGSEgLmut1l0JGnhVaVz+CAWe0A588AnqLxcLsfj6jP+aVqt1LEtYI
iV8WnYTEvOAtdFnHlhl5h5JtQ7lZc4GLvEs5dujJAPYyZAaVJKVQgtavClBMXJYU
xKHLSD82lKx+5mhTzYX2IVEmd6TNZSDEf+tWlItBTec7MtFr5QnMbtGHBmAhgsDj
nGHysIwTe4dH5zLJNnrwvosEYUxK5HP9hxI+9+882GBVHbN2lEU6LH8TOrM23SUi
gysmeFY14mH1U+le3dnk0GtyqzDKkmZ3vWpIwKrS/imHiZeYNNobM4PVnXe5NJnI
vsBP7uUkEiOdvFlXZlPTfQ0702fohuDJL4cnmT3FGwbcEJketbyHWMw42CS+yQkF
16b4sp+3HRilqnGxD7HVAeTop7JI4ICTz1cpTHemrmDVd0kzv8om//jXThG1VFRr
okOnWCMGVdlutoDJDwbKVbwq+JwnAMmXcMt29VQjWvuBRZKsDaAL/o6/GSih/+zr
CGQ/AMhkeW7+o8s+Wndd9Pnl0P5mbY3bS860jwcDF2BzH9jj0N8Xge9hIIBQeo5p
3K0Wo4lR0nGL6spP4KDV44fsROQjpLeveayPGGRIOu2OH18WiALGmIZtTdqSaV2x
iqTVM+AwNb3KF2I78uVF5GSymGzaPQsG4qSELYLcIU9rVDYBd1wWX8sfbB1v5QBK
9vDnolx1VSFo/AhVbvXacrZ2igtJ5srqpKK8snKPRIEe6I429xO2fMpyzvl9eHOd
/6x+KSmA1tzL7iBJMSX6wlpBKrmc67N+ek8jxCmtbnCclDhmrzHhPlWfrcnsda94
wIrLE9JJStArUwCY0PsDqQSVUPfr3LGAkvURF4DhMCPYRPHPtXN3HHtR1icV62Ju
YZ3MXAxzZuoIxBDvrE0SiNVB3Ahttibaid8r9UUviW7iyMr2Zx8g5EUyXA7XYAy6
YIjGT7xVhbSz9FmUhLFG+F/9hhY9MiwOL8OjyYi7rElpLOCYuBwDlcTUmOxcs6JE
xhyA8aUAdrvK9AbBc5aqaJCLFNnfLMHx3s+X2b+GGLxbm0KDDpKePdK8Qr8nMy8g
huQnCo71P3GIHRkN7TqNf59r28hdSn1Idv9fCZwDJoHd5qHdhPbLplMKFKRZOd6g
ibmzQys0mlKniPOI45n1pYqUfqTkZfXJwYmHn76TB9u1fr86YBvDUOiL2XcGYhau
okyDc7SSgTukiu0Pej0xRmTFngAyhoRK88548kR4B1Ok6t6ovS9P7kF7dfkl2tY9
I6V/YM0XH+oBXUyUgibRbu2nfPRDvJwOKYc3LZTCXDqBvaSlI2+eS9SqFZMu3tLg
sj7K5Y+HBi1MLg88Wuh8E6C1fOHjH39iMrWPmmRTj2Slosk/o2AamnsJbWYN3D1w
SV0h3Bt+9AJzltVB8N0yRkGn3dJTb8OmnKzRO/GT1u+tUFWgw4Xbx56Bvw1SjzFf
7C0FMsZRzKSybVQj4bcEj18N0wcf0fm0O7uJL/YbbbRnv64f+LOjt+0CeDMj0QY0
kQDS4TkexcbzAG3c9kxkyCU/sB/YQMn/j5C6EKqC7duw5EFGXyMkSNiqK4+fUla/
WOwT319Jhoss2S0OpCnSk4GuQeHE4j/keUVKe/DX1KWJcEaTGHbzgQozdoB1HuGn
ZpOM9wFecIm7GmrZyoYybdIFwh4q7LhuyToh3IR3a+0S6DvpFARCfg9yi/dIHKzz
dNf/pMBkoSDAJujJNtvSfEavUHEOufkczZ8HiSSXvBYzT99l9XQdcQONBNHA28Yq
2VSiNsclKHJ6H+Fg83ODfarKmi3mjxxJ0LliMVs58IrCYNMxxX9l4dwfSLN1RZPg
3E/Q7M6eSc6lJbn61q4k+qjQ+l7Gik8cIJ9/eYG7EBsrt7V4ukhMCISHcJoHinW6
D6KiQzia/Gl0rwJkyZScuktJ+S/IIxiHxHLhAQX/EV28UTTKbcRv4MipnUaON+/J
f2BaL5mUmwSmzc67zgSaHGYeg52g+/Gzthc4IiZsmjTeZfyBK4m8VIq092z4Tbvd
QA+jCFEycUTn99gjZJR7+qsJRHrgkrk3eSAyWjs+mI4lbsjMpZ4SpUh2Z/iRnvXp
auMr0mJcXRH9UiDoKgsx/YvabbzzCCK5AyaJwYB9TWdWHtftS6oWevAs/WZOqOa8
ekJS6PFqIStZ/XwU8TrwbUAibL8RHApbepzlT/63v211TJBaH/rXbVIhPLpKB2vC
eysuBv3w74rysPM6fkXZVJ7CQRyL5Q1xoYJhuKqVZBUmWpZAFuwTS6TzpOJoUNKg
/wmY0FayJXVwKq3GhfCWNi9KUnTJs0ZWa4KNozN4YjHy6HHo4OCu2MbrgKkb2457
m4wJrihqpE1Rn4rJXhpWVlM95+bdU3Xr9CXTbBEvMcX26q9OH7FR7ehp3d/MMwX7
oeW9virxOMd+KyWPWrbb7kmopUQb7PL/uvHxUIo96y0lVwvXxjwRzNqlHnV0DzNh
8Yo51Y8J3MrRanr1wg2fitcYZL3XZ4mF+eolj29hOu0+j6bTbiwPIji1enpQfXvE
mR6d72OyKrYEWF6Xu4fXNBBaXp1Pq2YfHHyqYYlBNdCZibIl3eEk2nEGjvpXS604
H8Tm/Mw8nkKymmw89zLUEq7Xjs88fbnq+uRKOBTeU3gxuhLA6+wqeAUrmJTcpAfK
/PVZBcW7esOS4RSp0mODYSEGqbM4iQtZ7YlJh5+2iQ7kfYPe/SGcGjTE5WFm1oVl
UcOFdZGfQ2TCRMkxkIJyc2kQzWrklGvnim8GzqiuJiWM8mFEDOsRCzKx6YUgyETR
j4tX5dJIdOFELdB6SHlibXtPeepVHEeYVOvxsucsXXdHpOopNPb95XoUHl5833Gs
1ao4hK2DyvKUYlxB9Woa+3TMpIkNsTCvnIgYPC581u7KooKpNlL5ix9IE2Hl6Uix
IDAJizZllR31ZhqW/l+AdTXrKCfC+jQSCVhMHH8Lve+RAH9LGtBcY50LWd7KyOeC
oR3q2HyMOA+pEk9KNj+WCdI6PEyE49wKj5/4H+D/zcsoCy8x17WtfewgOyzCqFIw
dehBfZ53A0a0s3vWGLILoPs33HYOO9KvLyXjUGi0mGCyaV9boNCDJiE1jdBScxtp
49Ay427QvXnIyW8Kl1uGTwtPIz3prwHmrvtkK7Iz+aQDvlWUmeFRl9dvSxBpNzIk
FGwrRD8sQ4bowcscLXGBE4IR6UVCez03IKzTHvoV8ONOj6UAWkb9ZhEdOxWUMCYY
CiD781u39sOStShW2XbLu97ebeVtjsOsNmy0V2wb5fkeZLW169ssu4RriyanpAyP
PtvXRRYhrtje8RKOjI3DsmFoTnDcWW2OGscrUyoLtn+4Ce5OCyJaEhV5wic97gn0
9ZuMZVJkVPVInjEkszqNdIhMduj/znUsJ5k0eVnaiRTkJfOcXMRtnYX9yaF39x4j
EDwT4NwrU2VZOh26ZDtlWX3Zl5ept6ioT5u7/rDsaCRZcrGASmMp7I9tHdabdeHx
I/pGVhg2EoURjeEQF7vG1ghxk25XlkSZEaX7Q0dgxhyYyL/CigPIcW3/mPwJxvhQ
D5c5BfF0HopRdYiU3pmy8//8mkG0qxcqWWLSx3/nCJF1SsUoy7UKttDQ4QgIplqk
wQ6AoanJOVA1CsKP7bMfjWsm6voyKkuSb1tkxIGuG/nK+yDpBhh9ooJ6JEW5b5q1
kA8bRzqkRmCk3xXG5UZ/Pfm8s9WIegBfT8vhhOfmX0FMOEzP8bxjbB8Bo6muUra+
se9rcIueIpMahnuVvnueKW8hF506laKF3yM9YCUQjYKZYoyqAeaSz9wLQcb0tWFe
nVptYRaSqMd2/nVBgqUPEj1NxYgiGfVqU5lTvCv9EFQxVAC60SruIfMNxUzRXG30
VUvZz712bT5teLZqqd+mLmN8Q8Zs0adIyBE+t+1T2zecgL4glh2ATNtQGZWV1A5g
OdhkWd9u+NtEFjwsQt+08YFRjFPhjBaQbbmH4WgLvP/wWq53boJcApZvEe2Q3wjU
R1B+j67x4QrVMNhQvcBZT43xyMBNOeqvbKctM8hgsj8Ha7UuiEnTWA2kB2D0qEO3
VihUAT1vqU0bbcyAbbuCZ6uhlpwaG2/lN9n3ThDXIARPwT96i1AI4yT9yNAEZMeF
bjIglqAfosOuCr4e/69Zw9UYVipvQBbeAJAXJROABsoifPJmGvkPiIzHyAnNdPya
VwnaI7PsWZE6JTEBf9fKhRGadvGF35Ck3zAROR5lHLBktJkPZYMNv5F/4n/nfleR
Co07YmbHZ0VVYtXwaqQdjBwKhD2ZYEh50g++UyvZkGh6fInCqZ5qhPLVxtl/6qK+
t4qUQ+bcooWG03IanmQB6I5Evuw/kxVE0BOQ9Yeiofu6lYg+/HbxxoqUHUN+vXG5
g0liu3nEO7ExhX8A6qF++Zq9OXfZF6CkDFqey4UFHKsbbV9QKEJi72F5dr09h0En
PaUDOdJMQnkHJFw/2FoXFQLpmtqUle09tpoTcci9zKFnaR+Omf7YCX/jDqyD+QWQ
qLts4A9O2jwG2GgWkChp7AuSBpG1lJEX/Katan+6miAIiez8pzUFu5JO6+Dj9d8i
FkJPD8qinVcLvHKpkCVOp2eHyEtwsCJ9Lm+h0vwbrXAMYhCkpSlbUWbedvKpNhgp
Kv7l3MR7/psgowmX7bJ/hkYfmvlzoaum/ESa3nNHBJijJ9j64xWCXmpS8s9wxKIo
Hx6V+5/hcSVz1WccjYn93Q6RMnxvCnkt/QkT1qs59i8qCbEhVZKOkEQpG2wUj5M+
/lR3zSmAWheD65gBpMRFdnTYvnNeyZLxNVEmaRvNv/6SIk7MUQXIXbjY5CNAqM1J
Kn6DbDr5ZmStZh3LncqF2FTWl1Rl5Fz2E6ue6kE2a3qXqF/PNmXjXj9OaqSsagf3
BW8cCsgOMBTerBQVrchieGt+g/q8D4tCUOCbvnjDwugnpi9q5h11OGEe7jgf+G95
yJkx3A6vxlzvJ2vJ53vdWV9atOezw/hvCTa4IgH2dOy7xoimae6o3qJk5EoATsXl
67q1Retqh86jgrXESTX+LBJtESoj7vhVbTod9/PZXYTF1Ni9c/LiEFNgRzUBkMgi
DHQ2wi6j2hSmt+87XGWfiWkc+Xr0MA7ZLA00wZbJaVnJF2ySYIJUJybl6i6hn+t9
00WAoIj7qcjO0wIb/7wyunuaFb218WLsnTg4pXfSzXDGoAG4M0Ywo6v/rwa9VY25
DRhvxa2pw5utCDmvyJrE6kTzh5AJ14IFDmw49DggUwUyKNdleFEQdU6BOvCKGJRs
CbARSWjxo7b7S086+zSsygE8Vf+lAI7265RK8cnUZ3Ms3Jk4UUeS3ufrwKtH3qrK
r7YP6p45rcLetgleReeMGrOHRka7uJeupYI9OwnBY/GUjoiDApKFvzURhXsTgPn5
qGHmmijGiN1u85p37T65NBWT7eGiDhjVDbw4qIqIaNMKdFAk4XF7oU471u65WbZg
pLKMHNapfXW8HQ0DwOloelncbBvYqsSFjTJ6Cl7zPxDTm6DfdDhV66vJXNi2l5n+
LbSJL3p6coVN4xFBfUhATXt5m01fJqpJDuYIPVjAacWrFxzUj4xA2cgy6R4BMX5Z
AN5tnn3Bgor8Dyv/7TBH8XdjWo9hdiMgn1rx18/2wy1U+pgm//qgyfO2ga6tbFLV
JC3tuQinTQZunhfjRWVZtbRrYjz1Odjt241Yo+syP08rzwfIvhecYWJCMrHz+UiT
I1laaD32jKfsjAdzBD9ZuIC6F/Q0ghJQEL3eZwF4zzYCD45152hFu1CAxKVgw5TK
44Vy2dygfAkgvnAQqBZ/sKlfAWyejcDaHDGpeDnQCIro2EL6OW+55j0yDtYMt2uY
fEZQD2XRNip4KATyDuxW3argmZrSaZ2BiqogaChZHIA1S13foEoJKBt+DGphlavD
v04UNwOCcnVhJyDppIamMzNhZCXl+I9MEQnnpWU+EJs2ZYA7bIIWJJbxxmeuYuwn
kULknzjJj/Dqez7bQoVpN0kGu/eDfC9fJXJ7h6hHWwu1dQkb86nS7QZpBiBuyG4S
KDyyWc4CGaO13lqr+ibAUNZkNhQyClRU6JkrnSzjXgggajuWyT4ygtUtiVUEDdTf
bm4tl1mojePTPzPgPUF7HPH/ECj3OCIeuueKd2m8Mb0Fxjd5I7oHEG2onsCeuJVg
r0Uvr/rzGdAWLRB09PTrPxh6w/GfpIjIYPfLtNm48jTlCQJbBi1Sk4Ea8z+ysMS8
hLQcIG21pyF41w1GFuG1s+/KGlh5nUiPOopSEFlURUrRNoyKXn5EUjeedJkf+hVT
wmM1Pa4Xfiu4Va0chQWJahKII74diM1cEjKioLL9cIpdzhCeNYKX4Wcne84ywDNU
mwAEYn/3fNLTcbI5YbH2QFwPlFz5Uui0ANrHVpJBSW3u04td6D/exlYD7i5DX+O2
fvOFrXjekFTqm/YstqjF8Se5t0eArGb8Z89Jx/qCmgFUV1pp7VM8zBEN3NV0Chxh
IWKtwb2uL7sAtt/QIWFlyguFqXcPkjaOcy5mGlvh5CXa+aObEabbgwnoskTA7uhI
VC2UY6m6rnTKHim+hiAsk+DAneGX2jJFr1oswwnkj43yE+uM6RXm82HYZ25i11k3
UWFbaQgeAH9CgUoDheY10LI6GULznj+TDH8SBmISxHQWeWI08Swcc2bcK76GU+DJ
HEtpjJDf3lVb7jD7OIVFFjoXiEMCUhBr0uVvclcL63KYNNebOAJFD6qZjTOjwMvV
ZGwSjcm4wb0cyF5fddyxTiDh6e3ZMt/0ql8mMgTe5U+kCKVRne7S889Fu6QB9aeB
kxYEqlnKi6VT0czLbWtfWMKcid9N8+J/RlcUEhXJX1awQwkroPqEkbCV47Dwo6I+
PzhDTG+csTax7z0tjIFaShKdmVnnAvHUGBXs81TI8LPyFJMluOvQgDc4xYnExBJY
aUQEPptkzegW+8UmTGDtF3BSQfvSfh4ihGSDH3uFTK6OKY9QJuAyaGWcYgxrQ3S6
xmu0L9hxhj4nxaXPrYqRZx6zFfuDHH4Ja6T4b20nDtzzT14utANdArY4qmMopQnH
+WC6thbAIpJq99dWEJbSdo84FGr2BRDis/o7xLvapqn+BweYtO8JJQzoBSEY+sjw
oY839jLnIONgpa/ji2wdVElSXQM2dAadVkk7Xhq1NoM+JJ9jfmfgjajCkvio8VO2
CPf5bU9Ud469PLIp2BFMYkC50tH2wCChVNBZGnYzwnduMzd4+RoQwb7jSe/qF4R4
JKoLIctxGLMmKmjr43HE742yhIbbG/ya15OHojg+ZAm/H0R1qbwYu7oSWweyu9H2
v909UFzh+pzU0uL4XEyQOy7KSWdOWNHilc7l4TDfvqO5iXRL5L5SP2ZByFf8+SQl
jwv543xxDXseTCOg0LIuC/pIcD596Oadt7E0js0EjA+lYMVn6UQBlY0JIvzX5Dwd
CJ35asZEPmDkntn5BC2vACHiyJPaZyjqVVnn5r4Dy0maDESEJjLRwrpsqVp1Gn8G
mcRMNRs1TZb4LpUbCaU6dCAl7wyoWrEfu0mO9WApRpbvOoJE6hKQmwYlonKOsJT2
4DCs/f2vwsraMDwLlgJLpNSnJcxQ10dusMpuzN1lA+U43lNG2Fsnnmh9gKJzDgcx
DSuQWTUFec96/U9p1ObCHnKyzzSk/9CUTJwpbxztdnuOMGwysMX9/lYehWNFezcK
gRhpABKaozzinDQCv1Me4KB+3iAv2Cv/45v+51atP9oVv+9Jovk+xD58Lp1Y+8rH
aUkNjTU+UUJ1tiuNa6+ETFuHzVpsJ+5wlSb63UTr2pXE5/5z3gYZYRqS34b8za0n
0NjvKc5ACvDG8ER0Wl6jJcloaObp2YlPfG6fjzl9KHxIL638QvLVKdc/6+CIZD7q
KFENBqrTJlM6dkv8hA+s2nGYry8bjnO/UxnnxDi/lgs69vV9Ed9Us3BeYlQ5Ctbt
DX6AZjJYg0K6eJ5vFyiInkI1bcV/jkjRVPkZixxS27/Mv/zIwkScKWzchqko4rBa
no7SAY/eHKgU6yYKSI5f5nvSejWal+VbZtsDsTMReiZYgI49Aw9hUpeVaCM9fDxu
JwdyVlagrprLzXcmqul/Qv3/1gBa9xmdSd8Td7cdf3u2HqOLYaFmbIYUu6f2l/Yo
xk1lM59kwnT2WQHX5ImBpsmL4iRMNg7qRjBJs54VZVmDsWmUJfnAScQfdRw9Bugk
9TFz73OmoK6SfEhGA0DAlctunk25dsgsZrEw24qOSufubksAmzq+P4wpHs/AWgPr
od7LW4ADcL0GIHsVk660OX9vqc7bhdS2jUdaQOfYDT4sp4hT0bESsZ07lrBQRbrd
qlS/ZfK6rdZIxEz9vAyMPgoM2QUzZHujh7F/CRDfCuM8fFzTnEhVzAH2ueEWAWr6
w76mzvbA9Hjvhqq4bysT9UwdwcILtO7ueOzOowGESZRJF59BmDE/W8yQqOP/22X7
OV3urGMn4x52W48PSDOB1W/C3Xpq3Meti6oMaJ+wEUb1rdgGgt/4CScXYEk/LQ1B
4qW83hKtYVN8lVL0JapWtwxa9gF6pQxzwUL3CKS4ScjyvqJKjKfoqUY8xM7Zy647
aTkeJSEtkeesUb/Pvhtw5KMuow3sYU0E4Fw+vVFwp3RP7VZDFjJ0gIPMSOViI0GA
nJP1bhJNlrJZkgVjiJUWkVUhzgJNaFMHbAbGdL3wi2VIEnzbWvVtObv86qNWfuTw
DkNeUVQ1ttF2czAfu1F0Ibd9bLTDuBrcJbMMsKtDKYOrB4Yqrr31WDZq4Ipe0ott
5mPV902d6WouuilGsRmjYeHG/ZgZohKWLRJGOga6z4B3G+KMbIeK5+zcGX5grN+j
QCcSb6k/H2b7vQ6CsZ3pg6RloVlSAwpXFAEmFDrtMZKWrPjas/ZROQ4vsFtMWVQo
eIEHy0MLszGgIH3gKGy0Q+wIZgQJGI4sUcBvTvQ1hqPlEKsqcdVDUP8drh9BT/TW
Zvrmp9coWc3wc9UOLBnc1fDI8viCynCwgJlVBnMUkfid1n//sh+mFAI6iqhvH1oD
IFYz11K6gDttl41LiwYJcItWDTnQmhZ54tiwOFt9ERzOmke0OmTd8A+yjkrUh2t0
26XJEXqbF7N4w8NOHQIcoF+aUMMPeyYXXHFZe870XsTDUHxCu09bbUlDIzMlME2g
3xjtfU+iQzTh9F+GiZiimnX4b2VIByN3Ob+JfEPnmjcR+PMlzt5QAFVkAWPg2yVS
ZPL6a1YabGO5csmOW/t321UGMPimJQRYSHez61XUEGV+TkPocJLJ/qS5Y3McbApL
9UEpRdHuRAvFMThrSNU8Y53YQscT68vp7XAAdUoNtFK6nC9QlNPr0SwNyDHyjmn5
7+tUnd3YQJd4TcLpg3mvt4UDA5GZL7dOZ2ZFRdwueFnbcDo0Tom5j4ThBTv97NEz
r35UvVfpPUTQskgo3A1MUzTQxBglI1/fhGNFtFTpMSVl+nRgrni1Qbk877d9vb6M
6IIc5KkfgvuXcUIUS6ys7bLw39LArVs1tQA5h7l3lWabfbt9G5f25EmIcT6GGhRI
aDdRCADY1KI4JiyjH54jJiscE9lInm7bkFn3mS372KgCxH29qZKYqnzAYKpUw0W5
G+Yu1iH+fJTVSCSwNrglQCro3gN1KCG1xEA1Ewbo1E8/nRAKzqRReNNy4Rui3xqe
WckqMM8V7hFZVu9j2G8vRV7SE0aM6tbad0gU/F3ifWy1k72md6hcnzLDSZwZ308w
tPt/iE16Kh21wIcITbUCKyfORgr3tROvaSrNUNBNZJN8dUPgICZVTi2XSByCkfq7
W6p2VVQjNhdf09fenkPqXxX2YSiSz8jKIaOfo1ilPjI5X6hbN7VwuI1PO+QyQwko
MtxME2bP+Ne9AqxvFB0SFz7PiCEq7bimUSkn3YcK1ZfTOR4BZfBXwIYIzmWnQeC2
Pnm871eCnm+2aNyS9fFJjyb9MHeMawJnT+xVKi0DbiK1Kl8AaMTPOgSQNVzUH1L1
WQxhWGY0tyvHTNVACjsxvWyCXRlH0OH6yYWdRfKec8j8moRGkyuz1kEKHb/gZQg2
4XNBfTHW79g8o/FoUxuP+yn3L9j06Grm0K+x/VddNsbNEvgE6rJmp5ny02x2m8av
boG+eXvqC4Ro8NaqPG6p5foo2PnTZhxhOot89inpZ2J+vn1y95L7bT/AC5ayNMKY
AgxVknL2Em6EeautbfWDA54gAsOvNxkCytdS8BWoxWULG0FJf8DJwu3zmWsnZ79c
PkTLyzpiYon/8ciNwrL7j/UBv2MEltPsvkbCEHqL6oEQL4JyJgZ6ofkpbvh+nIyd
L6poXGvouKH3IcBR+p7u/50+73tQgQpI+vPtFnjYTBeCP2O2blTVq6UzMZi/BE8m
WzaGTc/SYjZqlRoG/yrPI+jrycoEvygF3joZrUxx8m8GCj+BEVWSxRXTxocOKRMO
cCLdQvoj4oKpvxuJ6ZotZ6LXkcSgELQCtCT8EFzBjVU2C59dMzPgqvJQOeIPvZJq
US7aC6ZETSIPP2hEptEEGuowcJPTH9yMs8sKftWfhjkRBRVHfQawQp4YvEwO7pBh
e0I/+x0KJHLdqLjjF6i5AQ94e+8wEij11cdJjWCnPatLfc5o3D8dK3/HaQJ7CQ03
tFDvOfnShKOBgtBIu6Bpz6ljGrdvgbKfQJdKozl2ddCZxXchQjnoIH2Ir/iwc9hs
za7xar7NBp0i05CTh+LyuXCJkgo9VaQbJFFIOets4HQLrRHrQNeQjse3RMIcy9Iv
roj1JKmdl4KjRoQI/oE/fv5Xrq7QSNbP4Z7GXRpU72WNchuWtmoR44vwov6YsRm9
/Ne3Ne156WAPRnWBH1ya+OemtGrh75HQ/QJ4TRsHcJLseRcVQ0mz6WiXgZotMQAp
oSVlxgPKqKZFvqfvz4UQdkF+HTxodBBnKn/hShehe9Xk/YmCDYEIDbIeFYf7PSIW
7Kqj0EVcT1/Ocn9Xx7krNlTPdeDd8Tus6yPX9IYZhURJhQ5bmG2CWNp7IHjVcwWo
y9k5+Q07qWbrda6/wZ4iqEAQLaqMiZZaDklkoLqJXCWxXlbMPTnNDyoqfqgU0/jx
CsWbSV4fMjEZDiYennEbXptyr9LY28+7qTVUAu0Rpx7B8F4H2EdpIpZj1DfxzSsG
H6HPQ4Mp7smZWugo2VV0fzbwx8SiDbrjW2fn+vh2J5rDX1rKzu6IyBHz4u6Hahgt
ZjwceV+D/RLFbLG1xDbVotY6vCYVEneKgKmCaV50FwN3SB1v46b6XDqxvPihUn6w
vLCXnN4xuM02EjPilqZv+vIG7Mzsd+t7F+kVkvlK3leVhCbumq2sUVKZLRq+zZvG
vYBCFkaqlllTctl88WHBns86sVpyEtkJ7k4JyDBXCfgFr4pTWQT6hsOCSoTW5Qpz
T11mP1vFSai9PPadjwcMBG5WzmJGYztdBeF3JszWWGsKc7KuaLAvhg1N8zgNCWGu
EO4rIVimLBuWdqsn23xt5Yli5TvRZ2qNw2WmzimeBZ8qqjYLOTqNSytLVtDxUyKe
Egmk/OTjOYJoOxn7nxMzARt3x1hN6dlxhM4fYOWKhuf/k2RVWh0KKhYf1pzCcdLl
emsaUqnB4tJgzeopd89/pErjfPsOjPvvkHZ1ylMD3nhOAkxAoAiIxw5oMZe/WT8M
UZuHwHok31gZuoMz7V03E5btpayR94c3L5FXKb2umV2i2O16sR8/azns5G+hjXIF
pf9h7fThuLcrj7+lmZEkiUniGA7AgkRwbznni6BXmBkkIn+Wf5ScyLElChRFh+c8
vlKxCuljiexxo0NMkFYt5NUEQaFUJ1nhyeuZtljTaxXEXBPu3ucb/Vn5WyYjcJa8
r0gH6WvYlyPrJVmgIqHCIPHumdGdRZOt81mM+2RDfDZQms+KokSzgm2KNQO+hkX1
ipAiqfOyiDFsGmMK9uAFugfHLgyOa/DY/k6YxWHbxbpLBGKo3Jt8Ekr1H8cNgDDC
rZZ3hjWQSg98aEJKSJNmFgVVhTXkUxDi+/5ypOll4Qctx9qyVN4BpGXaZ2+XiGv9
EssgKSzeNVPm3/wX3gYXmiJ9lM0drlYN7GowkRExp9UWNwmBtqc1HXOniS1BkMoF
AAPzcTyd826YI9M9ZQIKpUfEy4SAv3wqBS98DR8t5DaN5MEtMHWlDFlEwogP+KmI
T2ukRmjaQwYvaBc0EK36bPlyD3H/1YnsqH8IH5JHuqV4wdy4sj9WoKijXlqy8QrM
7wcukYZMLYFikxEnq57fhIV8QOJZL9uOhdzg9VRQnjXuBSxkpO7z7SVGgPOTdxeM
JhjeI9Qq44okmtOYUjhxeKL/UT5jMCTz7goXcFUmF9gav3onduknwJg0AVJQvKwl
Wed6KH352Y+o+dZRjbAqywJ0x+4GxToJuJNVXqinekWz+3faBDozPtD0F3jAumUk
htRlLOmlmBc0W8mf26ffmYO/aDOfYX61PvRTpNoJ2gLDrCHMQl2TUj9/j9NldGn+
VBK7KnGoL/TkRPdnFxfpgemcLytpcxik2EzPnXnlLz6OqU7Bvl/1RKXl8PxwvOhu
VnOsljkgCpwQUkIz99NSZXKclFx9zW0n+kD8akFqHR5TRelG0LRlcIojgIiznna0
n2gQNGcIG6oPUHvEnbUDFOvKaqsh8Tzl5N3jMuyuNLWrLdEryGymCtqhCPfCcsse
KqmlpFNwOMXk9943LLq7Yb/Cc5oF3y6UPi85OP6J1Bl8ZpnOB8lD/edVpOgHAQ/4
CpNcG7tG379F2zEh1tvKg1qLsvVnuVkfrsPgjCLXIKiy2pUUBKXs4pxJD8TkSGFn
qgjoL5QQGnXc7rBdvRClh0hHHtD6ofofMAG2MZ2UU5GsraIgvZEjg/0mUPLJHwIf
ChDWzM/l+qSEOzuMkxNidfK4vSa8qhRGrM1r7BkWMB9Ap732ZVMZEsPzS4ixPrtp
qLBqwDdojGn367tcHudU8R9pissX/WQpTErHmJd5OW0J1kAi4GVnKmWF/iTYqsMv
nw3MYkDixxlX8wCvnmveYxT/5f8SW+jGA4w8Jr7pPFDK3LZgRidW04i2dqg3o5RV
Cgcs8UmdWP2WG4QUcux7Gc0ONPtor/15Vtu7M1XfkOX0bjGByVTUC9eBlTyX0xdG
iiKSTP6agp0FldhAvz5hMUNFHRyA2j7qT4lCbwJMvvHdOo0Q9PBTRdiLgurnHHch
Lc6hkC2cyFc4W4SghhOUsr8rwLi1SRmlL9HLMCo74yq6c6mWfMMF+FqGPxrX0rxV
c7pMTreojlpz1rJfpFdnrSlB0N4S2gkvPCvUkbEwSr6AzP9lrPWCAPw9DnteGoD5
rm59fZCP8gauHuiB9vAHW7kZ+KAsUM08T0CJOnnB108dVO+msfS4/EhbtAYWHHjb
ZcjcwVfPxoP65VOK3MWr0hyr4az8Z9pUZdeDY+viTTJfioQSrAxlKZQlJFIEmp65
XX7MaYyYG06WfqJ+LXjvU+Ytgw94oXfi90nI4F5WhO3BI8btIu8xQ3OA1zq2CWQb
b8Bc1eiKcrfY8mQbHc0wPGFxA2HqR21qy/32gQE3iAy5prFmFhS7jycOBC08ifCo
FPajZIC2aSXGMRnv3SM+QYuY+IXPhB0FvR+noWMdusWfnH0F/JiSVS/nevvVH6v9
aOeVYkPHRAFHdoLiHV31Gtx5viNCioujeX8azYv2ltT7bCXZnwLU/MntAWO9vfUR
6scNwkC6Darhx0WzK5tSKgxw4AHLzXKAEBayDTPDbzZU97pxIKCB99sqA2r2HX6m
iUqRmhIrJatrsZNCvmGq3d0Yhc/foZLE3jYIKD4HDjRlM5abwP0u54EdAJ55Pv0m
Eye+7wozMu51001UoynePpgFmDuwr4EXPvEMhBZYMvIvuc1peF6EsWNHKBmZmZKg
Zzr2Hp2uBRH7+WHCED29oXGxHpKmNreQ6MMaD3xZE/wTLA5kFQBsEWM/8TnevnLU
DuVOxv0hFVvrzLxFcERNN4UeA1tAPm97/+b2GFUN+qNW4It3lAMl7TviKHyBp5SL
R5U4aNLzcDIptCMS/Zc528q6YrCqz4Qvri0RTyamLhIaoMddH722sKThHjmGgbY0
gw3pp2pG7+Y9zLyA+40ihNf/DwR4+lO7bEkGdyedtAFi2cjE3ODd/Gx26tDosK2e
bjBBV2p+D8B6+9WQJlQMbY4pmzKq1WvrcCN3jP+ypLkH9OUjVXIOdA0nsZTSCyBx
x+5gIjRPeKtIW7uMDU5/PovgphCDNCQ3TlbXKQWrS+XOwnZ+geC289Xm8RQYFnYZ
24sRusmd5S6ejqilSvAp78kB0p8pfpdaVt5nGOPjbTdnnSZZEXCLjpl0CIzBjvlH
rb8G1lvBeJgxg9K5UY/zpEIvL+pMG9TDBBX06/zIYJeXlgG/ZAEeUC7KMjd47E8i
fAn4f2PMT9gpkC8d/sdoAzGM+aXzBTPjrKMynjXLubb1YJ3nZVVHZF40v4OJi22A
IgYPOAsRvl8adWNrz8MpIcmwhiKVMveH8u5ES4s4qsXs4B+WALGjDy0sbzGyWkUW
2hWGznF4yD8coDuuCBSI+m0MGzGgYinKbo6i+4D/UPIcyI+BDVJDj/uoLqcJvQxw
z53Hj0zH9PZkEHwzyu+aimhgztXgUGpnO4pdISKD/hhqjofi84ssxFpj6+FFBbpS
aw1j8bBDrOQ5RsSnFO8kGdJeS+2laWY3lI4ySY5kST6kF+PAzd9k6FQ72q9V8pdX
vWSkIz+5OGykwvnNCYv3yvBmEeI65EuinMDGM6WBRZJMxlhjFq4aA1cRMW02BLxv
KQIthnEpxr1aEjbIenmvD5WPsU1wljdMbS0rfGP6N/N8YplhX0GqEnBO5HMCtYO0
wgxYiHqC1MmYWoKoTmHgoDaNcTdhTet9Rc2UmENLSsbUX7UVeQsjehIspeSOM+fb
aDAMT+XiITfddgMQGuZHKF5slDPzA68825lFBotWOLQ1vUXwBePM9t0QAqreWkG3
FFgF7pINmdm3dMBaWZ8PI8UcZW5/IV0EP6DksdniFarT4fWKb3moaz1ssfpr4SVO
QDe8t86SE29UFIhOIGFO8tz1770vi/tKyWJCs20PfHtt04xqNzqhUHG1JeycNIPz
jL5F7CuhxzBQLzHRlvpB8pv+xl+691Es8Bhdq/ZEggvymw2xHbSRKC9Z2iuUzxVS
nEhL2YcYXCDVNiOF8rKzb3lIITxeT2r+phosakRTo8DHC1+pwfkf3/2QQxwqK5EV
Ko4cyH17NgQyJecXDIpmMvU3dPYArwjvmllyssEjO2TYqcv7hGx61jZDq7VqiAk5
4J2fYQn/txrBT4L6i+j8KjBUj16nkXGBBx+Ysvqfkn9t7VMMMj7tGOqvccpo4cVb
sAPuRsYlUnMsYGVEs43RFi8cfXt79jxg+POYHcbsLtnWpYLWmZIepMt+P71me43d
H/Bz/XK3qeXdPZFtZyJnN+Qz63Q3UxItAeO6halMkgVcTWYxZ0QVYC4gjthblMwa
vxAswATVZyeOVhnRnItn1iKyzipWuleV9xBhX08gmYOWOFhFbVqfrZWJ5uSD2dHC
zB19B52UOOBpDqj3P5HXxFk+4QX/Iez8M1LfjFlN7xoYWTVhImS+wa1uoZvVh3ZM
V3qJI0BlRJPhBhcxPnd042X3r3auymw08ZXctlnJbLsMkf6AhBCGTLMWiBfX8XQw
iYXmbtotC8IMPoVMtaIevLjTNcCGZTwf/npibVp3s6j+QiLxmaCJZHbUDtYL5VjG
mBwlXoKxM6+4kT+iI8XC97PxTrmnfj6HQmFOvPjSCfn+rhifh3JYX+oLV95Tn6gx
9rrmn4LuM8Wuqn9OyoaUjysIgCJ3j3ULRKQzUPMc2K4EsWvy7OoMMckPxmm1eNmG
R5fVazY0WZK6fJG077WF67Z2n61Tw39c7BKvZ7kJiWb7A8pL+sXh7CbQhE3/vcaj
1nSeBw0jGkoLWmLJZVdE+Vlr003799vWluNDmxLlEgsQYEoEjiZYS+nZyyziLb/V
O22zUC3f19YJBqEVTW0VPOzk+TpIzWTOljV82OGsGZhxxCqHTefe8LdwxdSm/d+M
CAV1LJWbjBiRYshGuBeWKz8JzrP/GcEaCvK/IEiZX6P6P3Pyv3RuX9wmH3RCBfAC
gJ3L8agndjc+C+9EvAL/gYWWxVdKuasxDBEsJtZcnDNYNGKBxayd+MqPQzDntDPD
C6ZjNtEWH3LaaOUZieVGQwOdHXD0Clfow4mExMYYe+RwoAY0YbpgZNTMLd9CIUZF
Hw2QLf9mTTWbdMfxxepatDyMaoQ0gkbhB4xk/hGPCDbLoaQdMxGj8+p1I0V+GXKK
FN1YiB7Ks5Q1TsPqXtMBKZaGssFcnTX6kuoLEE8iccVVNYNcCGXYkdm+roidSaXi
FuIzDfHPMaAQuUZgJVdthldCAd74ar1Y+nbi3u0qrcEvklegmifT8c+JG0PPXkG4
bwwt1znU8P4e33nLP1nRzlHibQYRwy6/dfzTbdy038/1D/Mt0/aCN5+TkDn29ATY
BMBZBInzK7WGbqqqaQx4HmyZvqC2zpTyC+QIiRDC9r9uO8NZbMuORD0E3krPiQYF
r2Vlap98o2hzGDTjpxrtEiNSftaV51cinc31OY2UqrqPATnuSDxscr1XQaYWA4Zf
407hmB1rV6QOc0HUZiIVOmE0aJi3noTv2GNHitMr8yT3hKYbAytgttY1YnFG70Xe
kV06y+N6dF34adz94wt+pLkdyEkfaO7LbxzYvE2X6PQTyai0El7vmKRL+V2libGi
QA7W5t2Fk12tw2Ph2Y9a/+QHYRTEYx5z44SHTCExOW9t7nFI4PO9qp7JtjBSajJ9
RGQcErMJcxA1KKVXWLes8Bfkk5/sDCZ3OkOIM+AUEfFdjoT2jFqT1RRGpS52A0M9
YA/vg3hinYSLfnNj4wx05dmNZkouCynUwRf0JZ0Cjco9bnHMBKKE0S260BUheRLA
26JW/E3wiiRN/ycnqPbpjof1xEo3WlQOuT0jtwzgZ/JFsNqpiKqAIey8LXtE7jtt
Gy1l454w8mPyQmw1Yt/pd9k4AuLb+2vNKwf3+Z87Iahp9EFe9cEXN5y56ZAKs6JA
E+CgLhP3UzIoaDVQ3qtqFAsijwHgD+NuGiWo+8tGyKSTgPmIm4CVbqNy8B7ZT3KB
2fB8dmndyMryn/EkMpleP9vCHqx7wqozNhfrphMA8XWaLMFiR89jzvkUYEj3Qos9
ttHeWOrqrYYYD7saght7coE52OA8dCCmCIco3lz0V3UUwwNWjXivgf26VyyVfJHX
HiUrsyKRzRM3fSO+j9TvoEcxju1IYPescfBBCHutdF+xZ9pGv2FrSXHFgr2kIA6D
bNUjiIc8ZiewUVpVcXu4iMAdAdB5m3ogYzZTk4pwhIBEcZEB2IQP49bJUz4lrnXj
kzH97V930GVquZoUKSXvev9sjmNx09HVXPCNJBFSmympIkZaxeSORFBmD3kK16Tv
LZ/kkwiG7XtaZWb4x+jxOVEboeW1bHNJrj0Hh6ggZ4UyjvQCTlPN9XfSEen+Whso
RprCGBCAEF4qyBIw0+ny7Yjp1t9ra0thEqA/08QB1+l+VFHVHKK/HXj9O9OO2Dvy
1kdlXNjUyTrwNhvScFCROtwjc+fccqiHLKXtm8C78RNViRJids/cFfAxRfGG7HNM
Ls2ONz+5TnqjhCkFnpJcMrAkw0OYqrPur/w7uINJp+Z8jhJvNNqM7h1L7ifYlup4
O1tpp/wvlW7yBsBFMCQ0S0SqzBavY+q7q4Hxvz2dtQ5S3qca+hFfypK+Iz6RFd4e
cHg6rcJCRXXdzM94Nkpr4v0ptveyQZd0bc2xRAIKn1UD7D8vSEfiVSWyRzdg/J+t
64jI3lqeTOCCmJdSpRHR1uaq1IjgRGqZm5E6dmDQSju0XJQyzrg+dAv0Ntvk3FER
EN1952gXoFMzRsclgqsnjhg+pzSZLJfVfath44obYXtF/2EubMg8AnQZ/QxGe1+T
5w+zY7ocLk9SiDRZXh9wK92xQvkZnfbusRye5LkRjPjbo9/jKQOqW7MMVO5wXwIt
951U7r6x1FqqQQEXbaVF9EoogvX0RVMjOnLt1Q2+lRBtU/TzfrFBneDPrz4tq3Ud
8yB1fwmFQWykMYTcDxj1dk1OeDCL8Fxs5BjopaIZtdGTK5WpLMpmYHEf3w54jp0X
l69QuuNqcHXQ4LCmXbx7tNHCACPjNmN37rXPf7WnRjv7FYTU8+AQcQXphWPk4kUO
o88wkExLGohX3kT23ojF/R6NE+Nz7w6OZhF3dqAS4cRg6iYpP/ccEP1yS9im/Ard
MpXBGI/JK+xmp9GLTVf81HUXBCKlLJ170FQ1M1JyZ/bZNj2hfIO3fXNUpV+nOF1N
qLdJyhWvQlKNz/1BdON80yB0tPmOOW1X/0OWKxxzu+y2a102r4Kz0S42ykUPlY43
c+AOhGdJIY5dGQJbrdcOYnffZB6uagfIKWyUZI15xiJPdzv/G0di7O6z3onYk1sO
lPIXEgmOP1ScLKEkxOvuxPQI1DZ/ud9M41qgFnDN7H70MrGA8eyNBey0CvBldSjQ
gc6HjBAypTc21TaPYaD0yqM1mxT9935Dzlu9j/CB7cPtxrC6XIkyTP9+2lsKcfZ6
8SU6YORoTjuFO7lgttfmP7iPsBAV1oPPB5Mf1T69WZKu4zFDxHiwIdxT8G4w/Bjb
VayaaqJFTeijCtN1Dxc5Fu5ocV0x9obNoDQ5vuKGPgFtsjkwgdusOW1x8oP72opu
pdoF8olW+TIlXRrRMuAFR2NcFeq8iQR2p+oKOodX8N6QWyP+Y1ZlWF3PQhy69nEH
o+Gs9JmLaodyvI/s3OeOc6sOA6/IiPM5X1eobvtctoALYieudM5hMe0FaziDsCEM
5BYXzNcEsc20/W32+6901iFdSHyuvgqI5DFROJKzLQFoQD8t3YjPwTjwXZobIMdc
wkuXM2sWNCuHl9++jmyDWVXJCFysPtpnswbGtxWm+JK/9eLoYepxHavcvFRtkljb
Hiu77GCi94e+kApCxj4ZmC+4hrKkUaxiNWQAun5qIjQSW306GLhQQy14R9g5+8O5
JCR8vqK5uI4uZrXb4G5shZxz4haazLB6VWH5f03m5bcctKdcRTWgskGhiPqcETNg
q6MLOl79aYwKnon+emt/iQJuts1HG3xErgHw2i/JJauzxE4Php46dEYEGWz9K59E
QNud/TiMNLwsM5P8qx9Nk9/b4sVc4nBc97m3xQkC2Xrh/hZxVsqcE/UOOnWEjm02
JPgSgT3HRSlnR7Wu7P47UVm8irEpY3RBTpGb9YUOv1sC2rp9yygOsyWS+xDE//FR
bjcl/prXlfv+4pqBEr1f50oTS3lLB7E1qABVF8jo7RJkaudg8S5FeZLe4P4X6E7j
7Q5cHE74/ztV3yyW2bJMvhuCyOni5n8EzI5A6FtbVCmN/terp+pxTw4MufxraYr3
+xGbz/zVx3hwxCDcWl2qOIB7qq3njv90PavtAWxdQgT3mhyTYIFoSp1z57fbhgAT
cEWz7+IaH57/h7HBOfCaPRxi8+q1ygugE5fp9dIfKgGaHtqNGzbPGvqCd2o3CPyH
tPaDSAAgqMu7ngEMb1W5M7aWgKbnyU7FgJY8CLucjMr/o7C8I1NcsI5FIRlua62d
I8+sc1rPvD/XIgNrdNWgM2rPvPXhn/3i5lPMuv8XdBI1kYXCdeAuTG8bfgOJW4Iz
B8MHAxOgDLI6Jz6OsmIHu830UUzdT8cUTPr3jBlKMGXf4wr8ez/o7cjYbjX/zN5N
c/LelUSHSTDxJPetWVq2Vye6tk9kTKpSgw08Q1LBSmu609a5/cC2jhOLW2sCCpRP
eH9cEpzM8lO/qpAirqJgp8tBLcvNs8sfOFkYCj1vCpP26AkewDuWcAvWbri6iiWa
cFO1f1+0DMYEWvo44gb93BeGESBI4SmY7U+2wjiGDAJ/AVJp+Eh1OFc5XzMXhB9e
+faEli7IM6H2bLOMVoV1SOj0oivjnsNk84hiOCuoQeAN4GDr8WLQkjAgDDM9sCGC
NCr6D1t8BtShAgZ7jk63nhoJQI+O+p4Gsip0QVIFaZsjR6xRx3hEp7nfVxlbNH5V
ySZCD9al2o9Y4uZWMoFOucPducSuZxRK/4eYN7r1WnT+AMLBvddIiQtIYu7E0FD5
tCJP9DflkId2ikcMNeLcpVvRepBkwXKUwU6Zi7FuSwN0lmjcEu1aOsJ/RMXsLK/9
9zZpmSjh9G6CfgHQTLo/P1RuZckoFogIIcHGVs+nVO4AXdLtweKRs4iLyU+35k5x
Ww5uAaAPnCfrocsaegOkjv33Bjsijs1Qev0QN7BEYMCCtJbIPYk7HjZwHOuX4dLX
E9JQWLDENA2Ejk7JlsP5Jj+/aPgzUiZFXaJqUKYp1Uym89BHqXl3/jRfvDzJcoZV
Dh2CO3e84cGx6IvRC1OEprrE3wzSNrBXoZaqOKcjStA3jWeIrC5jw0CmGTm7i+fq
c4uQQD9Nb65+Yh888TwTglYTDY79Xtogn5k17LmOLsV2WcZTO5qf7mPgdtYEUGqF
C21rRHDjp8oG7O5heZoXC7qhYjSY6y8Qi85SSDK7XTGBB1Oy6xD8uqQjGRqSvKJq
DrU3EfdyPY3Aq0ZzKCSohSrqLiJicM5lIhtGtEENAVuOm7OE+4zXaxdO2RnQaAvG
247uHqyrIO/mqhB/mo0liG1h5JemYFDGLHF3cZTppVsgXKPlLkBeYHhWnKPc+QXC
jhg0eI4ciqeFSS3do3eS2sYDME5vfwZV+W6Jn1xfTMfRV+OcDczYM71CLcCi99Rn
xY5Wpgmg0PYzDMd25xT44OiB2RKThvDtwPt6WkHoHdtqx7vOu4qjQ+DcdV5TxsL8
hejYO2OVaXNTWJFf7TQd3Mjrrqk354ptq2Q8hZMXuq1gS5BdWtavHx9ZPedyR9Y0
lC7upTVlROcyJhk4fyS6z5EwkRyWIcOxhgJ+np3jHd6S3QmvpPqVS8ZBlN5hXUdk
T2eFoRNxLGXJmlkryby/Kjuh/oDVKnmW82Cip3EELTZupor8BpMQ6d3p0rJp1itc
pw1l4XKDfGtGzALhNB+6S019EoSImNL1+SovroOBpcIoMeaiQvl6X5zwuMHNzThe
gSoH6Uw8kmgErdWk02+X/oP25Zf4Uv6L5JqbMrFDmQj4VJn/xh7+ZIGNFfN+LUyD
jmLHpjxnuQ/X1hp/QGIO8jE4nPs53YZoRlLba1gKX2pqKNjjJeNy8weN0lHTSVdK
QkCV1iGkmcUhXlsWm16yL49HHx0YnKmn1OqW94vsug4x542FvtsBEPxSrz6XolGm
/mAPrbyw5a3nUrIibvDE1pLaTSK9gX/QAfxV47dEPH+ta45M2QwPgjjZfZw8lFQC
04JVnK/9HnnvMQlVfjFjL2jpg09WtjWIG1aRE3gK3V1OBxs9UJ1Uz5kfmz5hrZBr
VPiPvlvyfJQoa9HaWI5bVo4V1EMdD/s8kVI+tom1oxmAOzM3KhaUZKv4q6Uporl+
yXEgyklvDpN9XvW142RO/QDP0sgmWmWhozh0UEFarbKTOgXASVES5olqfMlw/qu2
9rkabxUIgQnLT+nEDCDII47G3rMvMRmB4rr1fHxfaMuDmWGLuMf5swl50Mc/alRE
dyjAyKjoNoIi/3ljjCSkOCSMkS2CHPJHt+26rBH2Nl+WX+ao49j6Uc3aCDEQA08q
RT0zFpefi0t5IHKvNH9sVVzs5UlU70MdsaKof1onP3d0CTPI6andQcfjz2seZVOB
JO2VBfNZjQr0vw8bthGibbV5FZ/czTB2dor99GGaQA66Me0ZcYXiBmfNTMLZI4Bx
Ab3BxM/ZTFLL79eyEfUj0k5AqBF2mqiUsezyK6vzGC/SgeDJp4AVhcf68RhUwIj6
sxWZWamyDo3IFam4TZW0tR2jp+vIfKuPNLVN+iSb39vacOj0sq7eok7xSGPf2xCa
5O8bbViPIfBurCQsVb5dJDNdrXIsNnzkes7y4rbR/8V1qEtVUBFkyv9mez1aDGI4
lUBGr/49LTEKBkPXVuquA8i2h/Tgw5ywBJODCq6A7KilTQA95mXyijIgZnMr00no
BV+vlu9//vjlLa9Qs1dlQDA2b9gIaU6psl5URqgFMwUAb8j5GryfFY1TrUTuY73j
h5Ai3oiraDXiKU7bTYmPWFABoiVn0QFOgS4mFl3WoqBgSNSANVYk81D7GqIsVlZS
K630ZBXrGTAGJskqJhdsvnQPqt3/aSnKUUgJiMdfhdCozQOpWm5/hiWxuhwHuCL/
XLi9kcMmW/BzB9pAsUPArncBaI9GccobXIYEqpd+bfBp2yhZHi5DgBCz5aH4JqSq
ADOXgTIdAICbUeyvncmBY9XoONMzGJ6TZ411R47WT40D4/GLTI1tMTTnEOyfEsFm
Is+QsPCuHhu7r+ecyO2MIIEaEYkzXs63hW9w5mNxTt5BJFpgSF3AVLAbwIc3A/dP
IuC0orsWauLVxFhmhaftLEp3q9Sh3NGZnLQ57bDHeXaMTkk7tJAj8fs3cMXn0NLW
blIJTtRoSzEENREdAHcehjZPWr7IehOpQFS/dAFR+ExAPhMfF5d2vlusislvJ249
WXTLwby8S9i+Rx0Ox76eFOuI5K6996MXbDSWuRm4YKNO6FchLgamLVOsOt4IOuZ6
cXdVX0+5vhZddHFunjtVQJrtahGSXx1H1PIClBlQrtbAIc8vAhVat6YIDs+jvy0K
NJTvlPsPd6GhCLQ9M8YqFh/Cady1YEUBuF+mgb0zXjRlMbYk6jP/BGZnASmCOJPM
nkpG8zmSSjFa7lhw6POSfm2qRMOnGm9OvAq14gViT7FS0KK08ufmUAAHWr2X6HbO
EF2swLOmPHEZyJP2NIV9vJPcv0ZFYyOJQ0qV0Br+WwDosHWg3Kiqt5SO8vsi6ksj
LjCNHtg+QQQVjW9z//UuutY6DrkWwTFnq6ctG7aD1o6t3dMsKf5K0MMjLBu4C53c
KNGzKTeVsluErfivr1kHgKu9vDYU7bSP4ur54Fj2Ikgy8TjuFWAw6Yus5w5QYwnR
u7h+jDifp0h5YHih0HLybNcwgS8DcFW4hQYVTnkVE+0kaEfrCYgRKa1m1J867MOJ
8n1QAUFtPa/rz6yNaFp63s8xEiL45VwrABqxwWbkLp4TaTVc92jwdiBj+j/Wxl20
0LeX74OSn8hAjsetyq7BzywYaOLSGrajTXVU1UW2W02qw/+0yvpM09p/KTmAdZ1K
arJ2Gifi4HPmwfLq6AMwvYwqmos3EBJVBGdmCBeWViuqVwNJv5mCSzAAHrS0JiD4
VZhpsZPFAgqmXNSwQI/pOC0BMAuBiqH5hmj/Id5T0G7TD/5VvTwAI3OioxNp6dIY
pGaTIAhNSDuFuL/3gGOzZxSjMIx7AAcUmaRzTZyuysP1AByOyOkFMvaoMlDbqs5g
S6tbvGvxQEoSuEprznGrro+n+eqr0UupBmJmz4niuPJ7BwpU3grioaBiSxgb/zdj
OEk71s3l9/H7JLR11E4VTijd7S+tUgl+ZfczBfFVxc4j+Va/oqBFzEZb0ctoeSaq
GgQxjWfuMvKsZvi11mzR9OY2jZhqz/aAxxWD7Ui5xu9LyvEMHTIxBsk4BTVvyVpz
jSGY5SG882OARHNYgoDT1NGzg+GVviC6cDvqNY9W9mzzBAkYJ8covZS43ED8xnM0
TXh+MtcQTgiFYGXwHB+uRifkI3v7mDOFLIYDvJAqYUNaF53ah0z3v5DqcGGN9Q/U
TA/s86L7ohAp6JdV/kQTF3OICVcPjC/3GTmdYKmXfNh+iFs9FWiOzc3t1D4a6QwY
4plVFh2tMJHycRM96Gy/xsXU/+FHpw0hNq7E7lgOixhpQnAJSJTVOVYuE/9LGD9+
CjiUIKZEaIoYd0gIi3biVAhF/KMHNFe1ebBdvbzV0IF65ne8g4LZKS9d/HrdKzaM
5O1HrcguWEGkqFKHuIBta6zQFb2hc8C4SwxVkr7zeAqjAdWNpS6PZ8erlRAq+RLd
garljI7A2O/tXxFZ5yq9uCrrd/5da0BS+E9ofZSqcfap8YZSXQ0JtdCAKAkSAfXI
wgkAn1knIoxKBzAvNJDvX8X3dpIyhJ8hTAwU/0JEGmFKmrH+OCUqa6SzJAi4hJEP
GGcSzv10zok5CA8TnVprAECCCjZjlBbUcze18MwKET/4L1Q0RS9iJmWWZSOV/UmP
Fp4PavzITOvyhuQXDwO3iWepkOyfBjK1DvSUkeMTEPoPEa6AfOGeY5wMSY2Otk2K
VCimWVfkwjEeW/5smP3HDUkZnxmNYjqFG8yqX/gBd1eqwuataUhPZyGhEhnw7WQL
c75pMFWlv721Hqav7VKGy6bwlb7TjcbH847xVzAcK4x2MVnYLQ9/jh0Ee6O7osNh
l9IIVYVUF+7v/dqC4RgYjjvqVAlvNPKRpxhapPckYB0/JGz6arnUEV/3IoDwNObH
hhBvPFshhkvL51QYuu0O6Co7nskFmzyOss1BbFSqJbdmX+AyK+WY1rx8i+pUbr8G
k5Zi8d8vnescuFiozLjxoSXd/Ir0g64xp2CaXSIlKXaiNOj108skWhUjWDbeSsOE
0kz3LWnJSaidNKGCSfZvkrgeG/kWjGpcejKa2r1uZDBTsQSnUjEBr6rbUbTj9A/F
6vdTHhk45a+gKaHMPmWhRKot8TWKS0o7evGROWHeZA71+hSDYsSZmwXeh1RIZ9/G
OGG5M3OGymLhZY5E61pKhDtAuZew3D2KtLisRkmxkEMDC0LV34YMzJhL15CMbfyT
g1E70BcSYdIudLA2d0hCVb8HMK8HP3CN8rL7+JB5grFwvaWKsRlq1f7S9jMNPoB3
q/HwuIjMax/9boHW61NhzNkxoE39WYD/k1Kx0lOiMR+jV1sTbQabdQP7nhOrGyAx
RyVyIzEc86loPxaQBhFSXa8N5MOmFkUMF4LY23Amu1a8gTw3D0UnmBkNyMURT18h
yc9G65GGT48qAl5WkLTCu+1Yg2YeLjxKxxbw8kuh1GcSJe1/F4XaFCT/Uxuv2+tE
P167UYZf3Ewyc2gZh3MWM4KUHn5Sn9dch1sYyaEAEqjt7XSwQR65jnvWjH+px7DD
zX5j9zqrN0xwXLxS32xxGEFb2YCpzZEypDmRlrhIi8OuEU6jeEyV6wKoyy55RZKB
B6+TnwKKuBaxMRDA5n4YPXxzvVeqvHHNj4SAEx/WIkutue0UxxBbxqyBhaZlmJpq
AtIbjKHET82THkP8Y3yGaaOMc0I43UeFpr3n4LxN0IAfgFmOr/eVOeotYQkum1OG
KU/bDlLILV/lQTovzH4KFA9mmMmcx25bEDUJdnorAR4a8EDfjsL6Elf8+5DXh/7i
1zvTBGyEz0L2btiXRFjLxvEZGMkk/lW+hZzaLBl4v4OZh7qJvdfs0wE72pUa1Sbb
kHbaHDmnAXitcQYKvLCPij9PEYt4/cwCCv8+h6fSOpuJwkJy2Ipb7+hMrzjBuUEI
Us311n5Mv7AvgqHiwu6hOYvKBSg9m/V3bXPYRbSMcv/G0+y9bkFEg2qYH8P0lNkp
pnEg01BEXyZU8hkulXSkOaL8oB2FZxX/q+T+j8le2i8JtInstLk1YLWN0cQ4Gq5W
9NN5yGMb7+rW12A8n7d5l7TdAgDQQUgcBpqUEg2B1K359VXNCwmlCiNm3+zyZ6B9
hTcq59aiUpMgW3L+CpH+5B7KvZFMTaXGqn/IFFAduyiCgYd4UPGfN8YUh84m0fim
5NKfX7IMrDIgH/QF7PSDNqt0O+DF2Ul2B2+c7NpP7CD6oL8YWldOF/LU+tej6omO
CKVOQIPfCVWSJd4ZdSgKlQxBorprZDnWLJKOHDIvp0uOuxN0qSY1ki4iH97SlFad
dhS+Hjf+tlVygSpvpJ04flmz8KpgA39neCcfiZ/HgkLmgsHOm7iJbW1po1EKMol/
PXuUIid3PgOhOEylR7FMh+bUYMHFifeGh6cG7kjMUZVLEaLC9aMmf3WxSt6Q1h0n
zHnD1VeImImJrOmb4666nVg5w+9FdGXxZxL/rG/l3PUSDy/1S3Xi/KxvLCL/R2A9
sElnzK4SGb+KzU87M8Oe0R+YaoHTU7YwthWFv2A42+Rz5QzGpIyFqFuBv5+Km79j
Qid7NhIoLyNXjmj6M15wTdpVONqk/Otto6bDWPaPw/W6L+nFhQB5V5nxWUR9yISI
/eGGGRzJtzA3l0sb4I3YyOIchmpoqCCkyODo9SOb3xmSPSAzsC+u6lQjV4c9WF6x
oZ4LBrFxXzLInxjlrFBbpCuiLPBYBcQGe8OvHEVhotn1xyvVPQ5mQ6YVglI07YTV
6uFy0nGzROv8y2NhU1+DVQTicOdtDPSDd6a63+9ZcmhqDfRQtXwTEfLBz1/UQyYK
phfcJ7aiCfu4t3F4jJPiYxUV+iOg+/eXa4TMRBaFIYg3HLYd8FvH51IbPTm7DKRF
88eoU9Eo0rA4/q2zawtMmajtEkDLVNlA3tlaA0G49UR4u7SLSe2hKfU5Wcryu/S9
aSATCfpI98Yy+pvwOG774i2FZYGwuUd7Jq09lu0lg4+5hfpmlb4asG2dS1q1n3HV
JwNlOu9e9vjAV+6BArFlcRbQf30uqVIdx7po3U5TsNqt13jOYqHEOF8Eo/DpuBDp
2M9+SWcAhKGQbKd9CIR1nVuPXru5amOaZKL5/IArt7O3vjIAX6AnemH2eKGJixsD
3gLBl2mEO15kWVc2WC039OVsvFSkhMBmIXFPOzNiSuc3uNyYBw+snUvBVZzpqJW8
0AmyStknkjt3qZz2xCFlhq2geHQpO+JqFMY3ZUrq7WmtGPvml/mEOg/H3iLKNnu4
VhCozEjTalCpOUiIfFksJbU21lpWv8Ag2GZAwOqsYpwUKZliB2Ewslh1IUuAPxo9
WxDTjKvZ4RRByOK2s/ukJ+J7S6e6hbqTCdsiUYkuauL09z4HF6arfZScf9TROkte
s75gPI9HCL3tjiHZ66XR+khfPKE82YWsZQ1pyzQiYUAPcAbq+BPBbyEfUJpksWUF
TjrPXKR01aMh968ksySDN6s/nsCR0mTCwLtrJ1EQcs6/EfrOefBEe9yeE4UZezbX
FBVbsxF/NMXspzSwaY85ozjB0j7b9oMi71y2KbaURlaPxuDVUkXKndKqecmAPkwd
XtaQ6WKooqWzZScJzKic7ICjt4gJkYbbLQT3P0GjP6dPl23o5FwKh9WcaZymS86e
G5cbrHexdX0rPjt41WMgF8BTzMnG3bFrwM1ZFkYqmAhNONyp0k1wAF34oF+KNlA3
cZVR7mCFxOFkNtYxSzHBS889kSefZUwOZ3QZVWYD96ksYWO1hFeK+V/CB742tQUq
9zddMv73BRi1FokFRZzPmE8wwiwVBBNPydLYO5RWXJozczFSNv2PijXzvLawSOnA
2ZyUrbfo9k9MNmPXcHvVoYyfy4J9Ra904kmHZXvNqsnUTtrUE9WrXIwRT6OP1vt9
qtW5ECgMrverl+HYpdBjdc2qbADLCx7p228sJJStUObYjk5+9SqQc/zEnm45seSC
0fJXk02Fk9O0d0qZU63+/dpAH339m2w/1xYwtu/GaA1qOwZT5KHS3wzx9P/d0c6Q
HKv9kmTy3vkUERJR0ntc3NripST+zPK2Mv5Bi7tzLkhxYgStmO+HLSAAb8DxCCEn
Bsj0dLGbt+RGSfd7HNZS+neEDdlyxsBudFQj1pwwLX3EYyUc0XKNStPEa/ghKi14
p16JC2+atn/GO1AE19iAEsLorGKRxGF90OaQ6HwkSjO4CHRIzYTkeTScIqs5fl8G
RQg5nNvMABMDqXD6j/VvDnL0+PDrwDS1sAGYlI8IxYwWF6LdydWP3CUCJRXuzYiF
LU6tpSn45//Uor1If/QmhasTsOprmaGMbMarp7uh3PKu8qWTsYi5WBj37pluc6qz
TgifFMsnF0yiokNFQOQNF3waqyNcnGzP9Xe1ufKLNJ8RHOHiHBXOan+RUyGqfcVp
NjzbjW79sLfkbajqMrzTIbNJ21s/JG//WpNFJO9Ux1Onje7ISkCoRFsOLk2JYv6d
FVK3O24L6mcIiA0IityA4Eu1CDLlWhzvwav40f3WuG52pHZkf/N6zTnXMdO7yGNk
YK0ff1DOkP+8g3ePoVmxeWvI/xki08vf831cF0hR67dWgVkeJCQosZDDvig+HsM0
BKiltJp5TxGh5Jq4xBK4tTFz+eSvpWDm/uZIp2k6dYU5ErbRMmKxwJFDb8y09YfA
WR0sCHyRDiSmfKFyV2tmATptQyZIpQVF4dJGHCoDM+FW/LnZHbkOiG9bPhgUwcck
lBrkqjZusooYyAvDyn6rIGLC96Q5jn/8k4oleB0rrDqTqpqpK6zeKZJanSnjnEo3
kRJFbGLUDtSXnwS/LxK/pYzSHV24EOdj5YnSz9gjZT8uj5P8biiUBcNJfwx1TXIa
fDfqoze6n4X84JIU6bqJ6ysQdMgA/1S85/9nUQz6gPOZP4/i/MaQu9aaxsFyIRFp
/IphYj42UA7z5CvCZC3nDbhlBzkK1b3NqUxmWJW6v3zJQ4dx7wtexIqzUQh50Ab8
Vr/6glCVGz0Nib2n/6Ak2ZX3BTfVw5x+J3jj5Y237FRKjAFpPVO1OSZQ3ToODq3E
b1CtZeesIhseSC557CcT0ZBY6jusaE/3M4MVw62XHJrVfgbVwdLes3oOIqf7ugE4
t6g8dd/xc1LuekOBb10GdNHq6ru8rDEvZp54Oa3ElSIvEbJw7qsWxToVTFikLldM
zBGcdMaqpirKjVgN/sXAaWXARTIAbYBh14juin/1dsyt7/1M2HSgmkiSusme8F0Y
OymQtw4djBT2cKPq69yVpc8uEqsZ4mF9wrWjoPqyIs7WHpSl5WWcqCevQBJDUMvm
+3ZLVLvbTOCqYNCGodZRlZo39n6tDla0zBciydIkEOR8z5bQVWl73PL0WCRbS+DI
zJ01XznpakUTa0y2mM0EU/JSclxJ2HumaYUgO2JjvVleCL0f6GxijFMLX7azu9xF
x1aEVy3VS/h9FSjqUt+3rbjlbAHMHxdvoySpgX0nInJ6zfWT4e36uPCMLC1AWRY9
q1OgzNXIWL8OECZIohUnS1Nef6lQyWdRTtJDqliQeNEYpZv6VCoLD8D1HwTw11Ka
JB4xXPrwr+Sf2o5SJNK+Xjbwsod7FH4gmmgsZekN81CS1uNjZN1a6/cjTaM2S//9
0bSusIWScQac5KrjSuMczNniKE3TzfyreUq2QHEEd1UAd4TBf8ravoG7Tkm+IIIC
Uwe65w97NADFxj0lk7oPg6BSy9S8J678zKqEdOI0dXXS7WiRcmkLPGa73JbMF81R
GLLUtb/P6MtEKfA94sEXahs99OndeeXpR88hM0U3/ageaIwGj3ysBmKG+g9lgKTO
u3sgaJkNcHPvkE1gNWnJSvhKubdX4iIHfdK0ThVv3inb28S5bvcBk+aEXjpOPg5e
mttoCIAvRBzemfZHOOeLcB7Ed0pWLX4BuDSFUu35X2aAyh9dHEq9Q5q6l7hq1gQ6
fBGBYfQc+UxNydId1lJBaRfWv6BQVizc5vzpaOp3GZ1TzCx8U88zz2K5RmhV0SS5
qExqzed5xEHfWNqT9BDJPs6mMlF5OgpVlx63ZFpJpteqVD+6gYZQqqkw3QeWma7n
icy4n+AIIEyFOspsTgLKrVNFzdhe1tVM05EbUwqJ7rip4ACQiDD7MgB7GuVLQuEX
be97kytNJj9Z5C5eOz4zwdzzFBpYaFzIry2CzAqxb9jSYT8XA6n1vNBj+SXrD72b
7MoE2Ix6OBKGolNp/gLjFxoBAAEumLh26s7GBv0kA8J4glC/lNPWAjlEuBlTGlVf
k22YRAFM2SjjLVU+TmQVlBjnfJt5Twf5ZRXPEbTAljGC17oNpfIBXNofmByLw+ll
iIVSBi1QHT7pSs8vLmA98rzRBzCaXisEWkjhoh8dvH2WopSrsilgvQ8lWCEeSzuM
gxSFMwc9twOZuMClDBfZf/OmqiEH+RMP+qnBQKrs2IKqVzDSg+csuYiOtjwWMo84
0TbqYiwP2oA9lQ/U7B6d1Gumjqq6n33DpBW8lIOIlukCU0hyPRZoBddBlzTUrzee
zjPjDwRKDmzV6NpVvmrSMfMzgWXa0kHKWJK0mTL8Me121INiXPo76UOSLejSFHst
upCCGFVsV7O/Tv31/OkZrxxLpX+BLkHOsCosYPjT5mGj2rlL1/wsTCOdOzcWRzPv
W8A6W3CHmXMgxcoxe1gdlQN2SMe+7/l/2j3aKqG/bgZj3VxDqgKsfji5FDduKMCI
4ORY+eVa4yd8gq6+kZirzg/hvQFp9t1t0BzWqW3E/JsXXaS/tqB1dEF3PPOoiVif
yA7aj+K6MRa8zT2RY5f8hbM1ZfhSOuB5LrrEtbY0L9dqaREp2nvuG78bixNvxhdN
F7+bHf5xGQK+lF5nfHRpTS0G19iXKYN4qyLASuHUA+LdEwixKgcyPtXRKdFvO89T
2C0ARhF6C72Y9VFAbVbmM4ZYv46c2yqEAa8E7vk04FVV6gsCsDygmDn4W2aQZPUY
yuYzPg4ebPgkGoNveWsFTwP2o6gbSvld4GxKDK7ZwpUlTIbduK8YZV7UB1BpFfqz
im1c1FhX/YHvAk0JoIlPsugWtOJ6dABX2sSNWFmp381KL6jqHAg2X8I/JqzFJswQ
qsu8PJZBrM8XLzy0BcSffjabBFYOcA0TyLnxsz8Ysaj04tgXp+wHuAGOO4sCopQ5
eswXENVpg26b9tfmst2CkdI2WAHNggIuxHUaxTzoel1YOBPHjkIUWUW96Nthomvo
UwTxTKhWG8FpgZvHpFY6l2ILaSlMMAiYYXIquYtp8/QTgG+LRqF4uModGYM7hd/O
Of9QilAJJjSYBDgZgz7U01YGUXcrMP3wkkVnivBJFRPo99OBtTRc5yKo6/J+SGoL
NoWeTy58pHVDbUkuPWWiK0GnpaDqQcggjtrm5Q3UAOBq+hhrqLU9zYpgLqU6T2Bc
F3NKvOxQDy7Ng5YNmyG5ofR/IlZ6idBqUojKr+dgVh5z8RrpMZcL5srXVjfaz/Fw
CaOihvKPTz2Y95G7JLjbEoukUJgzrsxpNlfgRcdu+2HYN7q5UenKThvk6PEDUZ+Q
JgujkAHy5ANEGRcicQcPJXPgJpO0mYYdgqJN1zpfBoTmYnGnFh3zivu9ASahMW9A
Nxdinsv19i5/77KTL0RRa/Cmd6NDj3o08Bp60RTl2LCqU8OpajhMdQ4Ezdek0d0W
SKgJDiFgqr2CBPtvbYYt3j8UuI/scNmlM6rQRV/K1Oyo05xZvTbTjGh83dLEfOK5
5sBoJKwJiCZ/EkDlTmZRnIR4cSXvelrjHPzz4Q4pAIstHnscCdsFJoYlVGxacboc
1DN+G8YRc9cxOL4eFWDT/p48a5q6HHmIoLckyn1VBzXYwI8knqLXkMbQUSZCkvyP
grKaUtYsYOYP+BokWdi4d0X3IARnk7qKZIlv/FJEiM835UHU+GUMUI/sRqyTj8YX
MVQPLPVCW7zoQaiHxzKDi24WAHElvFWxnO5p/2dLZyWCZubSP+7R70lS/YAli2mi
vB9RiRJEc27RgTH6+qGiLW/o66i+oxppC3gZU4dC/FOHJ46SxV2WQVpGhvwTc7n1
vunYjyHmCvZXP1dC8L5xFo/zLnhMBBOiFZoF/wFhG0hYqmUm6cweaxARYwm4ACQ3
/6QmUduUCEvv7TfmqB1vsHBMUvpVHbu+OkbweYpfXJVKdUDrplC4i44Fei7+soe6
Ku0/B2F80ginfRoGyjQTEqCHq2QyYPGh6zrubdbTF9onFcWxiyKkSGYxNO0EQ8ZK
0qLZYma2fLb7y0xwPP/GHfBk2ta+ceVP7IyZcB0DGtHc4VWtT4K+BW4u0yfp0tkg
eMSdcnSGVTeT3fjI9mKE1IDBg/3FkmuValNr5s+hnoa3NSwOef4UjZ0SFjeNG/2J
EoXFBedYOKT/1/etBb+rA5ergk3RkJ5KBka6rYtjC+YfyeWDIYqmAp04IH6jyqO7
UYqFvSPJqNMZXn+rtFKct5eCJTSC3x4L446EXgXlhDkSnAvvy/TpRFnOhKQQBZNs
5Qpkd9W5dKCI82X63qrQfRaykglGQLaoQxxnAYNPfsHSO36RwzguoSjTQrd982jE
zIalPZi6e2XIvUgiqx7LQmTE8OOW4l6Iyz2cSy8qvQh4zf6Auh06O9JsR4Lbkwx3
1c3BbCXHwe3NEEnDRh5+BFjwW6faZrJtHQpiYxeZyOOukIuLcRM3pbvzKrzkAqOi
23NJi/e5rUHpzPHaVuXmngOoY2IbyYK1r+qwwQOa9+R5xpU/QL8afSCZmpFCjIWW
Yl4TSMdFmsF5SCJut5eVEORzbgoqkkTwKonh/730og1MpRoAGnq2VOIV9z0fIVwX
XKOAQ2ds/aPMRLjYHCtomJqz6NuyeDU7U1lqyUIbKGnnpWfPsE2RoE7AdpGs1u47
1mvVs/Epzt7zOz2H6tk1mnjreGqA5TxiQBcBEWOUO3aCPIMlfu1dUzYIVb9Xw7pk
1vARMcXbeIkYTtHOsUz1C/hWWhMeKUV7w2pdu8Y+Qko2JW+WIaekGJT6xwVK7pX/
vxklBXQ1L5ZIQRpjLApA6pzGDcDXVuHZyb8fZ8XFdCbqYWIaBH3wW5u7EDbYYuYw
lp7fkUoPeaUKD5R65UlfAdZrQRH4PRPS6wv0Tlmj8zKABv8t+T/FgUyGR1sUKNI/
JMA4HhtR1mHBsfrwJjNjbelUZMN0M2ewSJAum1hoysGyVtzspf4JcP4wXsT7DLlm
gkNAzyfTHBq4SKRqAhF5gccooEc4vy4xvmHxXak9znQbABF+lIL638SNH+HujotW
8mzNO0Q1WJy4oqlj3fyk8NuQK0gDrYQdK2wDTas57Qp/g3WzpuQY1SuP3jiZHEjf
1OdMbXJCKMvz508Jfs4DjpJ8w7UlAyq5MjGM//LHm+ChFq1fa/DKIu9WjtVcl542
dcRIMA3osi2BSlSD8D6A9v5jDGcabtX4JAD+deKSj2HPnVBNljbHPIz6MbJ7K8nt
1jYJGbtKR4kHsIq/V1aqDA8VC0bAedPuIYvqiBq7K8FC0RmarwB9jz5t1HyG9jMI
Gc5UBndXROIsF8bzXzA8A7a2ni6ZuCG1C4Qgyuyz/7yaK4L1LuPmzQuqZkDsgV2v
VhVrsmfySvWKKyEmo0+k7L9IBiCwdbz09Uifg4Zc9j/sG/r+i6cG9C+0qe1XI6aa
+I/Km6gj37c5dwImTfOMCob3ki379t7OumTryGTAR6LZYGTp7443zN4tVGZvu8Xu
bu6IN7I7jTRMh/ev4aGoy4XSwQSmB2zXwJoZaSQ9S8CsLflJw0cj/dh/fdaKqNRx
QtuFm2vR7gOPiOBrhgeVy3GhbLMFRUHPNPggc2mg8Y3FhrGeDoDjpNijUuMx9xfp
9fqo7rXVSH4znK27pGcypnZllXeMUc94DQl1tuY7BWzzJEmcgtd5JwjltecfNaUT
nQBD/XmvedYwjmGmXXWg8nKZjOUkWPBMKroNVoVbTwmfu0dxgGDMa1tsiD4yFyrY
5/54bRWiEYx/1MmtYSQ19Dfsh3vag43zvCxQKPkWsZHcS8rAaUD7U3uRbu/Dqjpu
MY8o0eyHsf7/gQu3YDcGCCa9hGNLYTrn3ahSV21Q4ZZrXgI37UY4aKOLAJK2fpSb
PaVl6d8yVqpNFvJMDociSCJB+cQwibVhUVlvy4xibEDeqRW6beWK4SvHkMqWwruB
7DvJG4C1WP7aia/S+YM02MXo3nzi3exqT7rAEXjx7OCxS5gQ5yG3KS74cnCAi8Cl
/BWp1dzhtwiEWa6k9/Th2Ud2eHSQ43akEPf8cNA2HVL179R58CbqHekB9htfouOW
oT1KBWWtC1t5BbgjekAof5mFmqAUATFmvOcxZOmYEU4ISuAcuiQVzWD9H66Ph83A
u2hfjNcnrB1lXLq8L0gz/isgSjyZxtvUkVRQWnNz7ILjXiglJzRzGl91p87BmWbC
nN1xg5V2xd7c2jvm0ErlCXKbPWqmWfFVi9gWPnsLwyYjTCPCtAoG8YeoEw1vSTSW
a0yzlbQK8t23vUM0rOjddv8fo3M0JbjVgitG5PZy/OssdXEIuL4nBeV5pm+hJvUh
RoougckLzGjvI5O7w485ITHpB+w3SgeEUlR2vI+GzqA5AM/vfxM9DB2XoA7f2wEC
I5xAWOEhy6/PCOe2Vm1aAfC+ZHl/NxzcE9mAgrVUPk67Kn7fsm47v6j4fBJIWhKM
G7JdHO130cnSe4psJb16XvtiDXptY55Q9Ph2Ue7zOOdHb7gHc0w2TqXD1kyJI0Ui
WY/t+8Ya8yBxLVEL9xI4qaisFQ4mNs71QXjra/P2vmfK3EjWqIvZpC5mli+RsLk1
WRTsVSqvkc0pI6d3qv41+/PWZSE6BiGRb/IvWeOTG4n33nc5EX77O5/JkTA9dCf9
GWVe+RfzFORwpNzd4VEKjZWEFW2oQLo7e49Ym64m0xuTZiFKhqrP8WlJrSrycWpP
fDBB/ME6crsdsmfEWNmAt4oRQX42Bo/+mw9OxV7yH79P5RowK07fQxtrPhIWN+nw
mBiC+0R0X3oZaRRNmgywOsjn8uNyicnuggpd9oIQkdFFH+aqYCNqzubakZ+P6hXj
uKhBUdqtTN3HIuDFr0HWkeExkKn5ARyqBph1dvvgQJ28B2UvsGGM2CIbIQYUTjum
aAByPX55wmkIo0T5iwcPlZ7pXcsmoKyBssdUJwUE7XWUQHlCy4CLiW1BZMQvXR7q
P1uMGNFmJGwm+zUPmZ54FV7PwGCbkAxczhWq0D1m3+PLJrgzvKJyLWI5uWRi2wPE
zpwM4J55dAQZ4E2DtPDCqHJ0yNQNYdvSiQDV2ysMyRMVb+PLhCeCxtOiGCrqLUWe
uDxApqNHE02KApg/zI851a6kYK8cZvXYOnwluiGq6tqkzByvw76DM480FdlZUh0R
NPgw8IzqSssu7h8aiZJGQQERRffzYDjLshEPW+oKLWtYoDPYjxHuZSV2ZsADTiN6
oWdXBcUtK9ahy/w6JXA7cdfbfWKa4abiIiKTKhcQ0C7FAj1FZ4rpEtRjCep7jrtK
PY138YqvinxtDz0NzJQOwgocLxtDzfTfr1M+sjHf/ZeXzChOddQZonh9boCVrzvv
YbHxW3kZTdB90rJ6bH66vNbfALN/7B5tNKaGNb2YEc1kl3rLC8ldbMOwAx3RmMTP
0l8yQ3KwxbBkYLxK12osBKAFrocKA9lTl4EuLKQWsOTBOhtAH2In/zZAE2OmBdhS
z8eOTO/emNB5JPxTPAUjkxKxshf8hoseGgoiBRQrDndQ0rFRS2e9D+/oeZ3Mzdwl
O+9DXnqKvtlHOX7rxFpmAyr4mWNSLjQCMIE5YgUicRPX/MHVhg8SR89qRPTnP/3G
pas+sqaJ9sT+Nxofz5fyTvwIOHwabem+53U9byGfSxpNi1IkZVxe2aoJAj9+8rMe
mHy2G1amLWaD9qvN/ud9K9BT2MLkg4bdIC7LJ8sWhPP0RYTlFFZpNcigStdCuYoU
4kjTQYmGY+jm7NQGAHimD7N9ze0LxQOGWcuiSQbD10x9ipIUuvHDUtRrqBJ9fK2I
bLq03l7Ev975QzCQpYq3A2mrKmgm+rr8/3EdHDsUzI0sqCGEfmrqtK/sv1IdKLC0
nSSvG7RciQS4UY49EsL6Q+KRnuckYGgmhZfGTfOnM+1qce0LUa4J4Q16YsT2JS+T
/F6EKHz9wBleVcEU4OEyITO0S2XpEpuOHgSMSQiuUngCCHm1jk7aT4nezjhF1K+f
PAmHmO9dE8MV4WJAxe4psaJuj8Ondt+U8AhAB+agxpcTE7W7UikFE7S8rl9W0KO5
LkEY8RfaKbvubOsX7dyGJ9Z3HCQimlTHuTDEfrLD+Nj0SeiuOyUuD+JEsF5hlO10
UzEJYrZY3QzfD4O8ho9kZTDprWvpy13aHDr+UHVnOZsPqwJUDL0FXgvmOJ/584vx
karIKCEq47+m95k98w99MS3n5Rm73Lwj83QodzqPSMsjX9DSTMHqUKTpVE+Nx8jH
o+fzAz8WaoK1A5FPg2HyWqNSFPgnxIl5LuqYljArRLRuKvUSSPl8a/3iM6mBUf4C
WujiD0dZ7mtKl0LOJtI8sJhbuoAjvgrhWm7Vmtmw1Zg1/yXybDEE2bAJVOB9dFfA
znEfxNgMNSSh0s+dPFwBuJlyOH53GJMVnYL+vboc9BWHysOCDSwPZbpUYM9lscvv
340NoNE22siGw8gjAeKFYuQztsRlnHkl6GwAex20FnabKMZSUlJYWSW0O9n2f2E2
jN92ThZcN5nxbSjvMOMtEy9SMaIoRXIdh5DexGByaoRH53X7pRY7/kMmQHgzjst7
J+vmZkVNtSqFXcA/vbnn3IAIoSIdlv0ZGmiZ+zAwjf2A5dQ92q6o4tmz6BdwZj21
jhmH15ZrQoNiCyMJNt1BnXIdAsDa46IgiMt97Y73gCWheJBHNBPECr8hiSctKk8V
xADVDfKrbHAlZRo47LgmQRP23WIKN5vcoMF1oqQPlWjVUYJJ+wpNmWOh8b8peFDG
AIoFvrEaqsXyygSCZTM2cPGGIs+a++gs7T0hoqLNhMxwVW4CsMFFFQQHkyXmmILL
eJUIu6+jw0Yjn6tNoxXMQx2eiQGt08/d94uTrytZ5yD6SqwzZtt2X6SAnFJ5EN6t
7IScWSZrytp7/JQzQaoVEpl/HmjkerM3lrwtw6C+hW2cPhrs+qOdMKPoyBiXP9cD
ANgGKg5kZPJ89T00ZMLwqswvgh3J1P5umAEGPI/9sL3vF20Dxzslsed9twAGFEs0
8WbOX5lSjXE0UKdsoW9Ds8F7zfyiFjUdnWB5f/pZBclZbbe1Nd+27KC68reJqYmU
id9WHwnYcOXQ+++QChHXjlnOxGUJgIUeE5UMoLPmOjNMorJJpcKTtgIPdcLQS8B2
DJ9i5pgTOulFofyCICOMkkKTlmkyG5ylmxwwHbCt1P7DaF3fWHu983y8emqzlhgc
cGM4H+4/VWZ3tlLpi+rWOj1FXpuvLATnVSzFNGLuqb/rhhzGRUJLO/+O2QjzZUk7
f5aS0zPpehJQnWxAr8KwaPu6hpR+MWC5/1pbv1xNl62qGwn5fq2Qzm066K313oWa
g/+0JvCFGv8I14+u7G16Q//M6AVu4kYM2Ke+sOfzvW4UPnD/mYWuWZkXJLJ7Je1t
5ZIwb0WauibsFEy+cg//m4EJ+xjQ2B08uQz5szIRukMuBGd77jS84Bbk2j+ABsFo
Q1X6Y/TbzUi0HvyqXXOHMRup6R8slKkixzmCDbiaGCAX/y9lICJuS838wMBBrrgn
5AByGzaNjr44QoiWQ8oJ7Ao+0BFMsbZTrZp3jO621aKAbJ9kV/wK8CmKgXi1Ri4w
NP1Pt2UF9PV+962EAweon6EYo4OYG8DxWjCdaE1Em+HZwm0o0TxXnN1IDe1BPHgJ
4p/wbeWNd4W81N0lNkgLqcseivuM/dvghCAtUVIavRI/AFV6R+ZjlZUbqVVIQjEK
Gwgp66OOVNEwDiP1nTPgsYub4gKApyzYae6c3Q8mNVqP3deWM79UUBst4mCqsbOb
yK2wCJz83v+JJfK2nGQlJVbBExwdD3fbl/YBGiYZL9joIMdyBIzjcH5qJV1n3AMr
2pi2+KjsFgRX5qpnHSE+5N2MAuCKrMEFJO6QQcrk1MqlIgK5aRMrfZxdZjMZ7iNp
R/3dWTz1oT5gPKYLmmwEkpuFtDDXH95ZkBYFdgZ+Ckqpbngo8rkJoAq01m8odOPY
J+q0epaPPbg2aAo2BQvUCRlq0lnpc9bDizFBm44yxkwz98pueI3SQwJQ9MVTLDbc
S1VqoQY2OupVGJfY0qzH7qR0o+5n0jkFUFWXIx90AJLG76onHRclo9yvgcAgQu/P
gYaEAGKj6RXT+hDYjSVcVpl70BsFe+O7UU8TcMpLjWR2oVzOKPIzFgMikYmNbMMe
31q2ROUfjHvn1uzb2gsfaXw6lH/rwlWjCZAjS5M0SL59Hxn6B/3iy3LLjGp9Suh7
PdtURcceOrD7M/DqaMLSJBk+dMrgkxPds/z6PN6egM1WLWh4LFFd574S7Lj/jDPD
FFtykLFaUQIWdzhDaO33GsAQ5jL5C+iwqp6LhFMdtLRC4BayK+aGnwiZug1+lyzi
jUIzpt7InCNBO3cvkpidPEpnA/s37i/35exSXInk4HTzjWXgZscbELH4GHy8w3+M
jc4J9/KQ2U5EAbjoXkH1dLj1Vzn5+iDqvxAOLh6YMMKgEm4nuWit2llchEyOL6Y/
TuBrSRcj9nThbZBH1PAZBk4M7cP3inftpE5Zp8t9O8HZT7gT3HFtb1JW2khvjGgB
6JUzcHd2R+7qUK7OJNZfZwQ+KKOnVkPPoxc/Y6vB6UO87w4GIEdXnXdv0nG2lGPi
cbJMYNLJxEA3DGhs37DT7356pvNMWio0KzzpxTrYn2mA2ivehBzxXcoTTcKIMf2g
+lkUXnn/MuSBS3DQsVsj6EgiLypwPaxThJbkjlDxV+YdrsbTkPLX9fkJZ7mI0y1q
GmxrOavNPhfYN49/ZpDWVZgk9SA4gDC461STCiTDRLPBZ0NnY5ZIVvO0e6EamjvZ
AnON0kCVVHAyaRLON1ilJYzJNKJjtefGSu6j76wu5H0B/IE6wYMDQl0oCPt+9FIz
btk7vuTsZE+CrzbMWceeRSVSO6rccbMwK/l6HxwavA+CISYjSvEpLH5lVg7gSQ7S
fxxD7bjh65XyHP0w/YrjfDTLCyHM5W7k8hKy1LsyfieULAxzWZ1ZMmvETHkdDLtT
rs256e8Y+GNTWCmoV9CzKHwEg0XDLYFFIAw5XjLJQCPyVP/kNciH7Y8nVRfLxPwX
H/yLt0nKyJS1BxIHfECfuR40cdmjXvOociUDz6Y6y7cp1tM6sO1P6XIN8iss86aw
wYLxG7fwvCBtxS2Pmq5KHI8YlMwtENMvV/wQO4ogSWmCh4kzL7oNYK6tp67ZnfZa
LmQeIfMomWdwQzqTzNwaFbOrThUOUoYMNWkdpJI3S4PzhfaJF2zibqVw4OJnI6+e
rYlIYoRhnoCDoMQCYm2LipzwXPd1wVaI5vyN1Hou/uyTTyCi/4ljbYMRa2aFKDY+
KWj/H7YKi54+6bEvKfRBUT7x88RbNea2mAlgZa1ev73ofTIcxAd+ycMc4Vb54nh2
RYQwAllvWx80NILhpQ1YXSuVazPq9jiMGFrJi+rhApat9sx9musmBO5B9ippI8Tt
AtLZSUqpM07/RziDrybKTnq0xL+ocqTmTHbpiSxuutS10OJmY/Fa+xgyDknaNpuk
Yc/7/c6JBuIVxUgQDii1jXBvj2DoDLxSgbOXjmNLIsGV8L+QGJPjKeAFG2AQrN3R
Dv2Pfd7ypm4fYIN4stJDh3enI0Ly4egRvQgj+S6g4nuGFdqJjexjDF0WJYHuLmGv
xzowm2JzKJcRe5UHvl2jaunH0igVdbO20dl+VZmHecGwPiQDUv4C6HLS9hiymm4q
xW/5W95+fOSxPxJXRH/PIcMX4JdCltr3C2l1rZEwp/8Y4RWgplZcbJHvZv8rOGZf
q4VjFblDLMfju8P1XPt50+vazep2lPCdtOXfrhMRQlDNqmqpxhGlTfeoANiYX/j8
gHs3N+T3wdit/7pihwjf8Y2uNrctB1so2WSvNqq/wlW+4K74rGbQZkN9hQ223ge2
spaRBjdTZxcPW6JaviOiPD8BCNkPWMeKcUDzjaaBbmwQAA03peqCuxivuKfkUiCO
bgTMYCGRm2hjGc2S+fnrj81fo7nLkbvOt9uaT8BR/ZitEazdqtsh3mr6fFE0hvo1
kADKMghUls8eRV4Wl8JPD0aiQTlczZXb28W0kQht3LHXlrI+v6Trn6ft49J0CgVW
9i4w4Aq5CQ5GNm44/vrcUOVze3o5s/XgMaQHVd4YZd+MeARdb9xmnzCKxH05N17Y
S7jnb8qYVrH6QOFWdrW4hCtTG/ph6P+076Ak9FBTpuedsZGb8WolSXB5W4YJkusP
qv3DA0Yq6qM4hiQggH2SsBd17A1lf5XydVbeXXz289Q+nk4RneTsA4bOD9Guf5P8
+9xVYucu8ExlD4D3ZuTPUR3WYDXnyyillKH7ndST3Z6U8ahgy1jhSLM25h/1DmOX
CAqe2wrXbfog+vcKCXSg2EgdrwXI7mvIPNZxq9zgwXRkxpLEDLA8jrU0JMk09qK8
Siavm5c8SBe5SyUen9pJ0HJehBXN1RXtnuubXHzvePyDTi8D9g3bFlch8d9SGANi
9SqMts6iVFlmZkXdaNSTb1IHa8bSGIbcur3EyQGWbcMMU6Cb5ByUyPUvsTLibU+4
3lN3KVmsdiUiPS+z5EQxssMWEZU6f+wSexD8+gOh9g/LzxVATt9sKZpVYZ1IFvGK
mVY6vsgOBYW1CuvjWn1FnDtpFL1aAlJgRi52uDfmVKMGpL2MeAENSneGJcEz3gE2
0xmQXm1rPlyo8O/ciad0572Z8gP4R8Y8A9gKh/oEPvgSxiz96YP8jF3GD9ktRWAp
BZUFH5enR9kFMxidoXfbrcC6PdF5oZTQVsn/zUUKfqnlkaV9ZoeWZOW+H6kgNMY9
QMVbs/D68eP1lGtfzjiGHAh0xdVYmE8VOBSxfin8qK8yFm0hY9O97/WrIBNPc3FP
qBcV3AeajsIGIRsbCen+a44Gms1qha5UdkkuUpzA/8uZ5Rf+I3x9eQPUfjah/30z
OrPUWTmnPW03A2qnkC5//ZBNalRQObO3uC8DsaQywcgI22Sqps9hDookn0xiHOup
5DYJAEV4pSLUnLO7UAvQXHVnsrYH17aGM3bueqizp6NjsU8teYG51rFsQQnhxltb
Fvidpn7AeWaf5y2f8y5t7Xz/v/SwrQsqQ9I6phe1jHDJggpQiqIhFQYItQu+KTkl
DOHJiyHd/irByUP3ftbkV8itnzaa9uFIvx+Iz1IxEeKjayQkzDexXYbnWFfH98hK
JY7BSmdoYjL/RSaiCgR2wqf5wj/Ucv6or3X2qc7tkubxEmD1QAa9yw/vpwtYhd1O
w3IG4ShxXBM4EqN5K5QIgHhnRrROSYUSAEDlaPL7G6fzuMlbYhs4AnBXBXVyOx1/
zHjCtiEUPzfZFcnTJq0J5p7ERMUZPdgnh2dS4bE/uOrh+InM/ZOjDTgx5bgJPOx2
Mflhe90+VbL/DcFQZHBKJFF6egBemQhsuSi9K1RrFfZhJ4vOt1ZUa2idBH3KToXu
LgnAz9J2Cleo9sHCi6lV5p5gnPwi5FqJ5S6kdsGHD7UuRHWKbi2CmLbF24NGq4Um
9jUBj3zt/sfM0PQkjsUiQHgRmh5B2a3UCRs4/mswGlMw/LtmpFk/Zz/b2hyA8dT9
eyGR0g7agFmG6+Xdmh93l836Rqo7fDtAvz5iEZcOazym4OB0X+hiQsctLq1cBWn3
TFDqAENXPsbPVefb4qtu7o1tXhnQIANyQsxmXPM6fIJeiadERHeclKnUnNw6lFkE
2icMaQ3v9m4Gsx5yjbNvXEf//FbcR7si/ytZ8fKINeHU0Ss3uA93dWW/3fKHtkkU
OtEPWPTVJk3XE7EJvJhBlQSVPKHSqOdiL5Bc1g0lJNm3DBpJof0j+wExP1M+p9FW
cLFD2NydToSCAn6lXgswo0KAtyolgzaic5YmkQT0d/RcZYb9edvbOdLwWU96Z/HC
6CIWGPzJSeXAraXaJWAwmsoep+CvpwMp4RQJWVrmqlx7P9nh8ngHC/B7vzZXgq9O
h7SJNh14HWevRvxTDexzIUSDkcLSa6Dx/dbZfFEFfBtyf8D0wVjv6X9rKvhpPEqe
631aXDQE+yqaLL1RlS1WxJQ0ILFEbS2I8GaY3QZMTOFmkzr5q/4oY9R/S9fD/ikD
SAvsC1aOMz1dwDwnFTD1MGGgiNNI9pz9a0kw0r4FPy8JOOxVSPrUG8sY1yaJ0291
V0KFL3CgPy4WNNfQBJYJ42yx8x3oTCXf+y8BRKTlVnxcoQS8JTBeyf7Fh6qfAXqy
NyxscUBhT/F5rabpK1YJy0PlD2vHPK3V4PcTC83JZSgOWBx8d48u/LMBoT2ckYQe
Ffw2+gp7b6VdMLpGaLsaJyiDgjQDgup/tZYAa6zrXejP/xigi1sur0wNOAXDueOs
5iHL0bM544AkSBD/TZvR8mNvZ/xmeVpflBcDUqnCt8aq6fR0D/nihFU+ejryXqb5
vHzXBa0DdjYXMP+/dTFhcQct0BFQxICzTfprpcX7OVzDwJq2lg9yJK8UQSj8vdTZ
Qvi5t9Qedb1JFVrVK+wKPBABcLY/2QVZ4f5Hv3EA44g7AoAP1h8eqa/9ixbyts9v
QqU+lHF8M8zx4Oh+TDuXVBheG55YxdmktHiDuIDK1J+CsOcDaMuUA6ceylgyUiYa
DcYjd5fEgLKnmvIUBo1t7JDE404WHuj48xuK9Yz8i4y5j+X5037QQQQDvB1hjNxl
r8iyEtjcGuv7VrZr+MpfRg1eK4wQqP/xeeNzFMhz7LVCMdHnf8sHvLXpNnEbGGJ7
TVdtaUQEu8JPLGk+NXdaYx7Dq8rA+EvdRDgNgDcObw0I4CrttnUpUmkjh+dF+kGd
UjYEBdnqzr1GhxR862E+M7pSRnCPsFHTlRQUDPXs3pPrIrD/5ryiBADwRovcw+zm
+1AVyu4GBHvVJeASlM6yd9wqFQ8aJHwmbmts7fE6e+JFsMlK/bpnWt8XyZ8A7lZ4
gZpmS7ljBnyGfn2ntjR7Cg+w83iAfSFY88KhG3ja9XdeMAq5TfSig4ZmboilpVTV
hI0dNVmCVqk50Zsh1woYiuXnwiBirAeCJYM2UDfZPeawbwDYe1PyJFUcNrJeSmJO
YA2HZTL5Sz39YJj/JsZZd5hgaxD6Fg9dEg1mkd0ef69K38SeG9ebM4ZWjhjP+OeK
oUucea1ADwOJkO6bt797iXlE+o0Ak4qPUtYoX7C+7sjTyfvchf0c6XIBjcj9Q/JF
FEUuLY/Fe2gDrtQRi60jJIG9CvuwlhLPnYbEW0RNcxRZGdQif+aL2Mu1FLdVWvTz
DB9FaKfzDhJQRIZ+m9nB9b7+ObRtZGspNgX33CvrsTmALjE90tUnfIt6V/m9IQO4
ofZ2XE3TiYD/J+GbPDVVGfvViS27lftMQTjx3GxLe3TNe0+TKDRfBYSgUbPBq1+r
h6YtWdyKgdFJRXEk7lzPrgywVF5qnJn1Gw8AZGUE+l2gc49JDhLLhec/A81iIf43
3bq8XWGXRMdrCFImnRxBgSToB18DEpqz2oqh2/gSC33fwpE9Jxu39OeKM60Hh0A5
3jP6aqW1dMenABJ3nNNXnTomOK4AdbnyHePILL4XTSj6mLF5YxQ6wsBgUmCZUWrx
4HTzUfbXPGy3du5SPQklLlqm2Z1Ds9KmTOJtOE4Njs0/lfRnZ+m9tQVsDCG0Ah8+
AjIwDlsVVEfbhafHhV7nBr8AHeNHKYVBtdTS5LNs+DTfgUgTyzYj5VXh3jH2gVin
GKva3rT5FeHXmHsLF//IYy/Q2GRYIhbH4uiou8qAVP2r0PUHmbZxpvgoIGaV6ntB
nlXCNq1prmu8KK+HNcRTC/mdghjVbkZRJD6imPJK0CkNOkt+Uv9ToqlAjRrIaom3
EO2dA2kweWMChz20rs8QJIK8QWMxdd4QNxyc8u9B9dPs5uVUkxPHjn6AQgGc0xGj
pXLEm7Ia1iU59POYhnATVgp7OlapSycmus4MJTx0qWfS3g6fuxhuURKSlTESkCpy
w2oWtlwhsGx3yCZY2FF05EWum8cgKgXzj9W8Nnl4zzG5+eQwitYVI1kCaUzKlGTC
6WzZkhhQdmPKfNXqepPa5BPN1Vw8Pbs6tlOkT6XCCAZDMQLQVqWpH161jpHghNvX
J0u7xwv6t1CFppmf3A8Zvv/Kjusw4EoMSS4FqQNzfa6GmiHz4o6yDMz2o0uiX3pj
xIZpnm2eea10bwtGk4EupRM6av0bP8UNHLPkL4M32LW3780Mwze2PngDu2sqlgdj
6y1wlm45+smDUasCJJTuv+M8tLv8N26nmFOBRYQVmx5/pDUeH+8dFCusecovw67E
f70H2BldIpGVLD3CTU3yFT7rPQm8gMi5GK/rbGCZK0Ej3lxM1kqXI+6I/JTfNHsT
xMnNVaU+eLY53niaxiN+oOW8KRSeCO4Io8saXcvX1n4WSnFHA/EAYUcL6NioUF+e
UhTwTbED8tnY6DodN2UBCxafP7QMpvUrnVWE1elVI3uXDdHH0NpCRjRioQeqm/R1
ulvd1QQQKm6yJawIl8jNDOh89q0lcvxemOsRtQ2jLcfqGN09x2+DAIY6VKVShzZi
l4YnyQsm0cHpEk1DBPpFrP2viXTRsDWrbTHCDvp5A2ur6rKl4KnRjDqLW9nBvU2m
yoYOS9yvTzn8TKDdR7fee4usR6x+L1oRwdETYGxMGpqCCiWv6qsoYmmBa8htat/2
OF4vIvKYd3yvltiSyCd6Evp5P9t45JtLa1KE43EC2BtkGbBJz9TqxvQfie9Eo0CN
Dhn6dbuFrVbqTD4BuZHZCkFxN2FYzG6rmcsfJteYajXfOqMH1bxgpW3l0mo0gWW7
PffHBmFUNMuQGFPiG6iaf1J3TVdu4vAmDETiKPAAgW+fvb3hiwVUeiDs1jABZgfP
/nlCIayi5o/SRPGXlIDUk2hA4rIN+WFL/+ce/9LgpxMLkxcquvrdh5iFLSImoXEx
s3R6X5utNayQ4+9bXdLwGgrXrF7wqx9KTa8rPgo+e75XbpLLs2xhoQY+T3xSIJje
WrkEVjFeZD080W35Vlp186UzvMjpBhnlfUk+kh3cvCp8cojlFQ3zDMDDCXYcoD54
e9CS3yh8RWHL6X4WiIbKST8fJf19UH/xIPA6qAn/YQregSavHtHkLLs36FWrnHO3
Bpl+WkKa+dnl+nhuJsn+CzHvv72iTK2jBhN8ma4shDwtRz8iKL8I08DWvF3tQtDJ
Y4/bSfWWLfN6SHQLbwEiZcipUOiOL/pquRx46r8vWIp/u4cPw6Uzuu7y3YLpZ0mn
DC91/eVzzTOunkJYKwtmdrmQGE5teMT7PeiSvpB6tgKlzSIUI2HtKI9WP+wbgf72
iRLbeDFhRKcsb8WLg1UhOwVsuYLqBIIrUqqNqsluu/Mn2X4j3PvAbvadnlXagvZA
qEkaIQT6ETjyYn/o/1YxTOgyJ27vKuTbAsnAtbq/2z/y0cr2j+uarYopeCUxRCvj
m4T/PrWyFHZ8ufgOPzNifC9UtbdK0rDs7GTt8ldK22nB6v19M0iKxBZcnwYn5O6M
cWhrCY+qWTYqaw8wN97Vy21wVYMTdPVZ5lZv2HHCAlPplKlBMAYUEOtty/e5nP+g
JqDgEULctE8srQrLXjeuVWsl0G7eVjIeJf+tNEOM37W9UiiqhjQtp+/DL4wC4SPv
WSCzhXGdq8uODQGOIpQ5myxLsrIuLO9Dho7OjoFQVJ6PqVYycGJ7tjZFR8H74YOq
pP8v/xSPdlG26VFjRPk3knlRxKt8WT7szeE0maPEcUETqWsth+bcINKwJ1HELDo0
PC2WE8XHsP3O7+Tb5uyr0oqCHg/id+2nhfh3KpHR91xYJFEj3qnWmvhwv/Hnd9gq
guEG0ZO7Zhg2XZC4/fPE9vCB6k6Z5rQUm+SNNHYmGX588ixM9kKNMYi3tI+zSiB2
k5y0Buy0wD0DmPkMWDxpHTYlJuvjiJEyz2j4+LIRPYGfgSTgwtk7BHXo1fgxhxXU
592YZYhvyY6OETRFoBzJhQS+fsZ/foS/qUNezzbfuP5G5cTYoRQl9419qr81aDPl
FdpFos4dp+/pXCtMZ/KAH2xfoa8wZ7o+KqhPCNEb9QZ4a6nFtUSWebjGCE4UAQkQ
L5huO96uiOdLOLlqL93eP1UodPrh0hT9BrgPrbSA3gGlrStCa/UerQujT7uV0o34
j5ZQOn1ia5wgYCaS9dP4py2NyS0GQS7pvRvt4Bijz5zLZpmxjnWorkDF429gXefz
g0j+gs5gt4eL6dVZLIXTGVB66EmamrAQkI+YPzRXjiuKOx+lsbDbhk1mPX8w/eiM
CAaEPeffqGuDT/NOmzvAMYHcDxG4RTvHaa9jmtKKA/FKTyZ0vqb+rdnVCMWOGGzq
BJeDjzikMAZt9uLaE/pzvzfnTZj4Emm2q1POleH3fy0xItQL6TL1//sVe0HUOzp4
2uEKHY4jDOSg71EtwerFPQJc2ctgNjTsn/pGxUpuLviIr4AARghm24AbZuS6qHXx
yrRRF/xOPjAS5nXAhsNIYLDBW1QLg61qLJ9RdDJrk5oo7LUtQh+r68YbajmkeGEo
cjeAcKv+p3hAzaft949ewdlznEZLkRrWyN9DrwmZi3SjWM5bZALWTDWuNIgUbxpK
mCsfQItwPphBB8HCg1r4W5fb439nrCM6u8WKHy+wO069wmkFo9PwwX5b9PKNBrK8
7qp2UrpVy6evDlvmLVZGTJbNQudOO+gf2aQdeAt2ELdUXT0AakaZhoEAyrHsKNGA
LAUI7dH+UC6xs7nZ06OdZGUoOMktlRo0uKVySMPwltz+mtkUrF1kBqN5vsIFntik
94V3Wp50n0gj0LbUd7zqg4a6yuKsnzns77VFRp5yjNbrJXVb4OYOvelYCmlr4VuK
vnefvqahdm+hUGaokcBeezZPP5ejSfdEL5BcJH2TOgBd9glBr6lS5SbmtnWaEipE
YBO4kNPck7BvwYQgMVJoegyLZt7m9otd83q6DXXf5xqMPcWXcnTsqaMu54NHlayG
DANIj++bWOIi+Lk4OFDaPgt5Fs4l2Vdw4OGilD/L3MhnuL8gW+No1Cr74TIe5Ler
9olDkY6nmMH1b5JTVNFEPB0SGuXOtFG6uuO2AxNcPo3C8e84EDVejj3WEUy4j9e9
zg/3gt9Hd7pKKKY3p3FjzTP8rcdtj3N31LdafehBd21tqg9ctx1Tc0P2+Ceuytp4
sdI117B0wMqoncgRocgI+saay3sl6vJ/WVJlYxPPSVfsDFUegx0iQVnFU7Du5WIl
mYDWLis7E1BavtIRv/pviSymO9nurxFqfAcOg+qVMXw0nDDzfynGKeao+kOCLgHo
19NAckOOkO9lvPeJQy6mkd0lXHwBarbWMtyhO5MhhSmOw6GMbqj+Kf6UZa53sM2P
U6hm9ZH1mVkj/DTjWz4TRfS9WiPTSr3BIARMPCCkd2tov6je6E+//0fa3vamMcoj
4DraVosYJd+xC2H2q2r2kWhk0ytS1jevWEBbbqTxP145GMxI4Kl6bUVcP7OsYazu
pC0skmJ5dtScOV8mV3eLy7EdWkJfJLj6lU8N72aiDZG+k0QcdI5u4IOwtVNPqym5
3N1XbuJLHnE3UjwdFaAvtZJuJrqLCO4Muh7hkXIN5WlhJo/OMsT/pHBuvezBWhuE
nCCFz0ojNNPApCzRJ6iBnCP9SCGEbNyj/9MM1/jVM0/oxO+UetkLUQ1d1f19o1sh
WMQUIcMBjtZbR+eZzLmpO3H4IF151ArtLVz3v6g4tJ6szFaf2wj79t4HR9PA2LAJ
bKSF8PFmor6JatzmCDI9nkGq3fZEm+MR1V0P9qFq5StKLic4Tz8l3kARQj1DFIgT
HP4/xVDY1YLRp46WFPDaMaMRXk7xpBatu1XLfq15Y9ca+LigkCpyqWEDIq6Hf2cf
lkKToRhR4QByKQ9wus8AXHJPmzr/tyIkqajZKoRlrDsrqCT2tsPpVk9yINiIVfzD
nbA+SsUvp3FYOjgzMv9041MNMgtKWCrQtw4Jq1pdTmN73C2T29TAFYYaparnDNHB
7zTdvQx8jdXBG0xgDyU/L+6OI8Ea4OtPr+OdS8ikcU6te8GdEEaCeTwP+nrOzBTI
UwkNtg4trn8xC7MKNpNV1uwV4P0nyQ4i4BMYWSuq93I0W4f7JdYHNCQ1lc0fcenp
e9otzt8wok8Mgvz2BpE6H1E9WdDY2/WuelPS/vD9NlhsAEQa0DbGieL/MC9mzrt1
cImDyHipkW1ZYlQ+WnTWyYgo9fWwu8Cd8+I3VxiQgCbx+lc/r5sT+oMmwbIeOR5y
kgCV3dmxbBdlhA+XdVpIkGiu4+hQe1CfT3TQZodyteqgX4uIzz6hzsLG7So3Qd3w
GmDz1U+ro+8d+HL5B2mRKt7x8P5EeNzJ0+nIosFrFeQqp+NMML9CFuH9L3Dxnh5D
CqxQZFXdrzW7aRG3ziivbeOfxRgwwJmZRqQwV1C8bICVqmpk4bZApTYJ9k9m6R99
Kqm4FNVYce2U4WGgcTqUtaqGkc1orKPB8W9NAqLjntrbjFQRbmus6HxyWwNrJVpN
nHZksApJhAcrNDoMJd6ddtAmzwe4SxbC7z9QS4q3L2AdrWXC09b9Ewj3woBcVuv4
hYh7PHdHMjCKhvXkdWJrgupJRFZSFmEpgvzH+p1i3zM3vKWPhaOrG7bAe1jKg1CS
LNtSEZD88wtiwEXc1fXkZVEOB8In+hzEI+CalximJidBgLYFzDIJ8I/Cdw23eQ2p
HJQ8ouIEnPzJUFHz7qHeC6NYdiEnD9Cc/lkyPNY+3eZk/yA4EDf+Mh77EeYophmP
+hoCY1r2DgujFGQ8Kr3TDrfdw+BQFOfwNS5D3z/gHwvazH7x5KCKovBCVo9qnmuq
U8Pd323l2gSCKvX7UqlaeUvSa9YYgVTKXmxo6COCWjPO0pdfCFPQJppjJQvUzAVF
b/UCLnmxJjU7agYwxKQB2h/HTUWJ40FNLKDnqto/vZH1bj7ZO5leoQ6+hXrtlP6k
OZdWlQx5JgrhzMH7il+cj6W0q1PX0edcQ+w5KFzdBRHsHqQYaYfJX3mOqbcU+wXD
TN2InPkGPjn+l1+HOtEO4JfD/akovdpZoRq1mqrQ2lSe1oLV+DLgD2UL+UMbNAq4
xlNPvV6nnnKJ0OaHIAwkQcX7BpSnEzPKa5KJ3kPsT29rqmgzsijCL4mh9V1B6Yjc
xK0XpP3lkuIrVJPULdlmPNGl5F+uF0f8FcDuS8l1SaIZruwaU6AqcXkXz5/h/GuN
Q+fwy37KMCUH2TjlsWO9OlB+yCV+mf5Dvm4ivMtjL5rAjnw6ml5u1Rgex/L+5GYy
8Wkbm6hk1l1Q4JM4Er1FZYrZ76TlUsragJaDVJUh/xSo2JD/iksUr2MmAZKNka3J
dMIxH+6YVufbbENPXHtrg6qz/pRvLiV1zSGUPjunB25lWvMMdx/OQylmNceMCRB0
A0yS1g1PWIS77Cp50pap9VoXa5n9u6HjxYk2I7RsmrV7cnzcOb9N6EfPOLNDcJm8
zFGt++/k+knELluDG4ehgrBHafOk8iuSKK/+hZ4DOyLt5resEoE/e1xUzGEGdSfP
qmDRrABfRk25PjQdacuQvaWcDD3kJFlXFk9PqKrql7T1lklZdPLhslrX2Ys9KEIF
Y8gBa9lGzEHdhXtkN0XFzx5PIhl+lRKsngXhjCEDZNJLHOMA0/G3NO1vrTLTpu5z
lQTSFxM/yQB6UzionzF6/nXF5nMY1ShgiH1CLYtvz+u9zYVRAiumT5lLtTpPJx4c
R+hDvGoSNPPrBrV852pOXkdRmr5mlrziVZzpYFcjjdabKqeiZiupFutdim75jM8V
svNNpn4l3+qtDk+59rhguPJUmm6nDni2RRFFWElhLpK+ByLT+IzxZtDtzfMMUbuD
ySyB6Yjo8RlJ045Zt7wAUaQql/A4nDwXmCzkHI91j3RnlvIuMzlI3cg5Z5VbVbR6
iZwtrLCGbCd4AH+Dx8G6i04lK9QqSWJ4fpMNuAVI/5NSIlDM2kE/U16hPYK7ruCj
mdY4lKxRKTIeo/5MmWWJ8Pr0woc61Wf5P4CAMK/b21BSmOKwal36ko/pqxbkk3G0
U3Bzd/HqW9uitUujc5B9hcxuCRCKEj6eKJl6d4DD7NYHyvilXYz4i9495BLoFOU5
thxqAx9StKXinW9ZRypXrtQ/cDdRD3bQfVtFHddXt1zUHbsq2eTwj23CGyu2VTRZ
GBh9aBtR3gl88/VOw2Gy1GM8hKKlJOiwlgcA7FwG+i1s0c1bumdcfKQNgvHAxnac
idRSnKWZs13R1K6KIXgsa8CZ55P/NN+uH6/7YNkeVmxDAC54yj3xKQQ+JjkAVdpr
pMl5pmoQHAS1HYvjP8S3R8JUipvNNMwL8abShAp0Ola73FmdHl9FqnVFXy3K0IY/
sxF9gJxAcFGhNEsB5ZgWrd8TuhFCoFSGvI9nDbZy5kcfYrSL2HM1mSCHRXg1Hh7/
EfyzAQ6CnbSZgwvKXdJ1oa08WqdT6V1KcD/A62JXAxrI0g8LxjbKCvzxQt1+EYmb
s6WednODlwWlBO7dZaZdH3gyNqcknpFm6a1/KTqVRi9sm6NRFZIwelbTMNSA5lgi
d7BOUS556UUGeSmMleE0HwcWfimZREAhjYR6yfVCN/n3f31Opd+JkbRCYnLPhsFz
AibwtDduD0EICff6JraXag5JL+dA/+Q3TPi0d1y03dQTmKUhEuA2xbEu64K/DcHE
/tO23kAhRQwrtePm4Vf7szOwEkp/SJo4218ADrBZIAJ5pBMv0jq/R08lEbBsSgCD
tefR5jVZ/93Tgd3mKgiRXXuyHY2e+5b5cEd1yTcbkCKHWPCJRg7YW2wTYA+lEfR+
CjJivDfeoC94q7hJcoEdViGTk/y/4y1hmozg/rf9hodpqpzh4rvUTGrf3la2W7mV
sM7zYA2EktgJE27luZkpCFQWFnsvbhz2DmN7SglQEfVQVsaBTUW98dfUpV0jtjFD
fXaNXeevXiCcKh77CwqtZNY39egk76X7PTTQsbufX3HgeErwib49cDIkCj3jL7dJ
ITGEHqtK/AKvjfD8XCNew9i1HtwdZFDHF5HZiGAYwA3y6YFeigFRj2gql6ZAEYV/
OcVyU5tYHe36fKaphgr31FHoOB7kqL4v4iBKlR8UCu2b9cgj9cEDEH2eDcfAa5jl
FLB9dIZxsgb1l3Sbe+qTLrqvzU6OWpmwvjBcuNGxCW6qLv0j3l0jSPnvCJ9K13CH
uKwoCtWdZ1GtTAVJjmr80FMkQSmQSpaeEDEHQvjzsLyV7mKewcSBTPHAL2rfR+mh
nu74cISa+aZZGeUBq/fmFKmbJ3HiQpUF2nSb1X1z0W/ErUL03w1EwWeFYx6bz+EJ
F0t7u1xx5daO/dnbst/wTZpVrBQH0hXBmlaMT4c+Lb2srUEwcDlchFMfMuoBOwN8
EGWXATH9dp8hdRpNL8x0kBKuVHZvZT8VcFJ/L1VhbyIlRLxt8HKOx+HNs/3RiZuj
QpklU2z7Ax9G1KcZceDWgERqOoAYS9Lmks+SjSSyUmCVJcL3RhfiwK7pw2HSFiXi
7LsWVm6EdoOUbqI183I/4ho2FBqrPmqcMkqkTIgOt6X+CsOsWD4QVxEN+K83MjHk
WpqEU/hch4iyhCRfH5D8r5zDT1xY5eNUuYld2xx5L9TrF6U3rb5CwIPPIFrR2n74
x+tnuXQatnf+QoPEtk2+ymbfXS2J59lCOSJuSJ4zy5KS1gTkITGf60Sm/sI/5zqv
CTcRq1QWFhkhuc7NNzte8ob8wt+AjsOWbx9huPZ/rouomipIIYSIMPZmZVtYKEar
xlWX6pKAYBvdHPhtpNPZuTxGICI0a60pNvaQXhiYfRDKavgy5pkIup3RNAvfZtcF
KulsMG5CfCNNbDJLreOZDC5R92uT5gB5d5+o2pyOqDXANSByrBl5Ew6Q545nbT5F
OLU1448NNE7DSPefgUMaxp8J/8PjGg3fLv2OGn721o4YGi4MMbzVo8ZG8McVEJB0
01i3xgod381ERbyaZz3Uh5nvvK5DQJbNj+f3s55OsKp7yj8u0zO1i8y+7N2tBnVM
lMrGjDEsBPs40HvhkuKI0YXXGEMDsU7aP+1hvCfg7k04+eOBqTKFRDyzR/9A8VJ3
uJFWgXSo3Nbcu9N0/VBgr0FDhOTgXEcF4NL/zxuQQSHu59aLvoPbXhhZLnHYEapZ
2A5vK7fHncbg5dF/b6C2PeEKPAES8DGm6D126t94APQ3Q7OlmY1YofxUHcLlTR2Y
pQd2HJ8Ky/dHW53DnABHwcEAQTTsrH57y9pFBFhMmpgjd/MuVxiL9E/GkOHV8f5a
OUOMKL6Nx9W2iEwF4YAU62oePzI+AIqQgiFbT1N7RmopzUi0kJkgOvhNmv4y8EA7
6nStKI2JFWpV6/tkcQet385NJnDjVwBsAcH3TVRuXTR1WtD98HWMl4ACp5CUUoeu
SdKS2D7D48pStZWuswsm9Y1mEeQwUdA/3msPcfYBRDwO7eTx+SWuO6UOdFJ/hdP2
HmEXVjCR1Aciq8gNtDUld2zrgxbsT+IfiATmvpLv1QYC4E/Fx3OQmVdRAi5T0lG3
NNIGpZDNmqAW0k/V9lSDgg1wAbomWd8FvFij7vatYHl+mk6i6IPRQQKGVibp8pF0
L5wGWVLbU/UKlnhgzC6vbgf1XSdQ/pueTN+1DT3TA1AIsam5scLBtfocTAOQsUfC
MC4F917lyIBM6klMVGr2hpSpbLmCO85BIA+22HoB/uXp0gXjZ/tV1fjLxzUBYi78
wPQP46xpr63JKEXZncHWHEw/cn2DMx17YAtiEcJ/EX9eUVo0563ebvfDeJVP/UJJ
mvvqpu0vygJvjD2z9Wv+t9r6oA95Q4PhMq80ZPwkos+EiFMiY5j95ylcBWDB+Dc9
yA8U0r8z7RvFTzPwFCD7U3hcihnusKvjiEGL7YHwB7SbvQKgqKAytck0Jsribh94
edZ+HlrvRzCnUghq3HcGp9lzxnmWM0rH0PBHefNgc34E6JACFwmK3MVQ2zLTNmX+
PRLy2cVTeN6oBO3/amReEMremKbvmquSq8/RWxq3+M46ZIN6+CeOEdRScFuB4xih
iFLGJFlsPQ8sunDYDDhlptUfLBhF3BENaIqXKvXIo/3sWPCELZUQk5mogXIzx/Kq
EV//2s6CW94/1P7Zy3BQLyslu2ei0iQUfShUv/7QHXeI99ZhnHjmZdFGAmieoGgF
epyeLrPPFRYDRAUPQzX+6vgFITyJolQNi9clpgVN80YIAHYejWjqne6BxszMUglG
UxTZ+9yIrmNyOJab4/Ec19PIldySPtjF5HPVD5znRIZc4dW4bH35tnm52dL51CYd
HnW21wgM/DWm02Eww0H+qFBJ6tPj3xhfo4DbKeuCvn2IKvuffrTkgoGfmxA/GyoI
DfrmX8MwwgKLzm93X5dN3BVuH+dUv/c9RcMzFdzeEXpsW04q56F69MWXkkw9I4Lt
rprw1akaoQOiXHQYUYlKgEeCSu3r1VG+nx3wkN+TlsdUUvQ2AEGPQYWJCaoC7yBD
ja/qOTr5w7A/shOlmUkaHpLM8EQOMTusu+pmEbMr0j5R3NJOjchhDW9V0mcPiMfp
GGGzHz16CePECFMW3zG6E5HA/87OctVbP2NpzZlJw6TMhpplJ8za75KTL+SyAynB
gmTp0b2Tjqw7wR//eY9KGBfrgWIw+IsXAoGoXwZpOCmtxsEwmKnMAHjRZq5Srw/B
C+oVjTU/jNGy00Xo5GS0oexjWQmV9thzY+sOv6f+ATWoIH+h7PZuWuxOTJ3dEUz9
1Y3f2BXBx1bgLO8utY3aFryy+BtlpGw0612ph+LsOCGeBLdHY6YOidGkBGHGysr+
xEkA6ddL1lXrlUUv0i9n88Yt0THYVzObWgd+BlfW+z7GgUWngW8weL4M6maoKTsy
NiNgmC1TLBuo4qahY9oWZe2JSiixSS3hNF7i54g9geyMk3dn4s6MboL4YWaVyUSf
SHYtpVvRDNn3hhWvaYKdqm/JAt8PuF1dxwBRAprXIJ5/haf7jdDYUmw3JrZ0Ih5a
0n9mtGBfeU75wyX2FJOmkUe7CODVP6g7wrf+I+iVeUX5zuyLnyyrpRuDlXDPmBak
6xYg0y9FuTgmgz8NHcn3GTNr3O4kku0B2ZaT9a1WU7GqVxMUciGPHi6WIKW48mnK
hj7NuectvgTnxHVvswlX5tH8CWdQkY6UWCer9JQhrKThyZGjLmm1WMCG2/VSsrde
0RlgC0r+y/vEZOZwZziLjTepKj5OuIAt2XV4BHNM3HJAA4BbwyWYrE1ZNKsl0hCl
MA7stdxMyFuLlActKPJDfqMwFT+hIkW/VLThNP+VLUuYwJuYpovqBtI0AX0qO8es
h96i8j/ggH/GrSAGNFhTOGa2t6/caWGo136ibG2P3xLoUN/sADTm6W0kCu7fyPO0
DEIf023TSsWCI9kRZzYbqgAjFz2q7kkg+Yu9hQIFr8Qs6qSKZ/51moAtBXwjm1Z4
iK+6h4q5t/e6Lc6cnGiZCktTY0Nlik2K7XGme8FMDJ5NQvnPZiHqqOhFqwHTJoRb
0SMfm6LKT47MAQeno57j3xCaMXHqGDiifPZuanTzOj0u8AckTTOH/E2sop1/UP6T
j+gihBZp0cEHHzwaIHFwhwwainhfdQ7hjdE6SvPShx0pb40aZ5bJTU8GzlQpyU8c
dlxM1kLw3mwm2XXHspEDTuVq2MflVOBvYc1CqwGASeYDDp88iKEFtR4TDLnks/1o
+haMzkvH+ecPoptMhiC8gO/amSrO8FVKmYmpJoBKUEFvNIdBGqRCkJKVh1bUkdY3
uQNZItwE9hyegx/qLlftgcpgj7ttWmxyqzc6d5Zw/ED4/LY6sbeNZlmnjEO02UJA
49F7SNOJZ6cNi8I7QLyanVG7UMeXUtemy9KQytTjY6pXh8zdu/I3e36VL3HuDmhf
l1VtwG+DqYMEjNMe/dp1+gj5WPAmcLwWyYvmNivBETSt8H+TT06jXS694VAXT5HA
hm1CcCAw7Y1NnKSCO/L3iLVdwQ2VyXW91iRcdZHOfbjXF+rzC0OzCrEc5dwwPQQd
jbUQJOcX7nAkFUkx4rbljpKi4ZqGkOLlzAdLDcP9u7ZT8zZwy5sykBPlpP+Vgoef
jfB27fAtIVBVVSWxovKxKpsCsAo6e6aCommNnrtHqBuAFMcOwTktwNTRYqM7duLq
CG821iWKBUDpPiWXnB1gper7WiVQc19w2UNBUc4svaEsdFy5HafgivmF08cS7DDg
prYWFS/YbwmQXcpOnhhOIu3oH8RDCWwCfHPae0vf7J6oBmEVUhm+BrWgEephu6Ip
tQ/OHn4z5S8zQzbWqUpLk1691MOaZTuAlOO9Qsoe+9cSEYpxblZ/KcDoFqPCE68X
7TgEUSNYwUdX8rX4DCkoUi1/azdagxD98NOlz0WlQgbO6HUEGbU+kfqOdCkJiAuL
VUo9wieUxroF/21c5rJqcSHDbEap4Tl/Yc91bWmTwvdsNoYUfDdhhAHTbAWJlbH/
QfhBGheCsv5lt4mwWqo9nEgm366+IIxGSRbCwks1VvJIR8hI7ZDHqPyw9/jsy4zA
d+7iEUcdEJ3vUO3XH/ZCoVq/z9pMrjSRfMA2az+ATllsRaV7FT+e7q3HVfopvPPh
1PpckdL4w680kP1qpuU6kI+e1A6FbJlG75kvHa7fBHGtQuqZ9JchhuCJYY8pBp1M
PWAufBfLuDmSTUb6s4gwKwuaeEYId0P/vMOJISgjfxlUhazeQVCi5Z3iNiklrQw7
6oZRSPiIWdQRHpNWAN6nR/5okYl4bXiLeDPAiFtPR/qbtf+33VjQQ17qkJl4K6tW
s4J3xUkH2mKc7BLA0kb5oWy0osmE0bAEc99I8rMw83Sx50G6rzK5zbILFd9d6rhW
XeAgmwhIx8E3mvoebS4DObEuoEzeTO5L7aBiiKGprd3a2YzW3GYsK2cUl1JKMMe7
ZP/bzSVb3lniKxDjCbtmL7aQmiTZbg4YR44Qjscs50hCC8shmS1ZrqNR4XoBt1hl
V3CaDgHHXit7guKVDFHnbxjwMRyRjd0ZpPn/joPR6WXd+6WXYhl2o3vuCm1XKMkS
0yeoLT7YYjDc5cfXXE6FJrs5j+CK9IVQJVZAnDoeRPjTOPrRbUvRpCl1Ur9SImvY
7IK33n11L/UNFsezOnubc56DePSUTWB4caUTSRUhi7CyB25iuagfTOd1HNYGTFQa
Ovy36f/54XHIcKnFsyxqN87ukyBrHz1wIfnNyyBf09BQRX1gfwYWcKtdwoABpEhJ
/CXedM1sC3gIM3cwtyXf9/85bLyhHPqMOEuGv2UbyXVbF9eR7RU/rDiKTbeXK3jO
LLJkydBIJWjIdq3Nb+IrS9NT5sdfDtRDlA0s847KXaoOju3wJ0MBjKmWssyNIfjS
7NI2hl0M4H/n0RrJSmRXtMXGXGQzJK2pNy9sn3NDv5CmiNEstRC+jlE/5akz8tlZ
KT/yuK+ZpKUFQWNoX+afgn4iNLoa2yw86hg8slmH2GUvgvX+X1JsX2RZ7cUxu/5G
dyPYVaATP6SWHcna2WVaS8+mcZWv8FHYwpB4d0suGLCdF308JBG2kJ+JH1vOxjke
YgZL+4dGXOP9/k2dHX2Lgo1zoqGFUUV6CWtmJ2qtTsOw+yzV1c/vo+Bz3zQqRuD9
IV1D5IVPWHQg4DNBPI3z7ECE713x8yVM8MXoBTWT+bH9JhzDlYSlEHc6A8oz7V07
h8ZPTJ8FI73IrJ0jdGeQjW6qXBI19p4REQA0RHd5nBQlOQU9oeWUgaMW2hiAmHjW
I/+rbseXOn/AlLdV1jxu+UwMC/WDMvUUbWIp3H4I0xrNt2B+VrQmHrzaZ2ItO8iR
HvfWwIiL7NwZRiHFdd/txkMGK4nie2w60380TCYroJdcN27B5yti3YmjARTUnjIR
CfRaw/YwiuW5MOCJX5uBimB4fEE48guqw3m6kyx1cdbHBxJEl0W1qowz2+WDn9KV
H4ZSr9EYpLZH63uNcwCsh2P6yInXRRFTRjS29wZEV2GOUY1WlRos17IPZg2ckz8W
jwYKMVaJHkKEX9129NWKravpoRV/E6uvHwsKV7weIL1Rs8cbtQFTpJtTKZJlHl1K
9XzR5k5xm/tQ8FuVr3hdx56s/Ef7gy7OejYTvvlmaGqHxhkcmgyevfDcvzc+9IHR
U0yLI0xXt7osMrFD0dOjfUxEzlKfRRASLY65lhmqZ0CsJD0u8rYixEF8+1ucNhRa
4EjThLYrcdLz6OyuEtOjBlSadVqsCGj/k8cYe8CAdoXLJfD38ZmHW/0JepInkAaV
MQrvLRSbTEpzSr65S0w20D+fDf8ybV/lLAt6dKp8sAjVKOseRomwTRP2JRW3+8wm
RDt50EO5Aeqd6zUUVeyVitACQlA1BQw0IZQycV/sLnuYjGJ7hmDs4yfX+9659NIi
LGexapfnMjjbw7jDMACcLaPMOI+PRxumCI8zu5D/n1hjpWD8UQQSATWRtnUWYybl
g8uBSEU/oqmj5rUCBDbSQIGkIQ68tPYmRTsoaIiMn14IGqJU/0929ysjIB0X8/Z/
Zeuecmm4jQ3as2urrrWTV2XN7u31+X5P1sK6dO5FQxR5Adhv9IrxSWFKi8lYq+jl
N942ITTe07MEdHA77zT+IFlxYOficgpFv2CWU6EDoaZlP25W98xoyWZgKbrfpAgr
nBaKLs9Q8osUFgkgJkw4cdVFnT0qbqCwfXvgqOrNp34XcIEPcKic89Ni/fU7RDOR
hEg7JHr97ZeEB64XqyuYPsHj2jJDXMyohFK03IcziBg+RtQQxcwGyTgmiMtyIN8i
z9FhNSKt0fZl42SXGfASdReVeAVuuhsOGX8U0s3PfpOO/Vz9CDXqoVSLdMTG7iRH
WxjlBqGK7w14sSE6XMh6q5JXnAS7lWBGfVYVUTPEQHeRC+ia6B9bBj9tgQt9cfKT
/rY1PHamHqQpdvxVOgSn65Xf4gDhlU8oayHT2xFivmJ4SXDOiqDe+vvnEj3i19Ge
ksmN1TpDsbUWQGD48XhnAfxT7EEpb/tkXCDbxFPN0XLeoKiMDJbMpwqoCjc26K8L
YUNso5AThh5g0LtLe82L3yHqrWXxnnBQ98nwtM2KJmCgmk6rM2/YlX0neBTPP2oy
5FAAzxMd69eC6AglNekNEz2jzgC7NZoCeb8F0eEt3blcCeOpQH2xJMl3oy51ZcS8
27RBxkNyXlThKqdRvLPljTRvtkuURP1N6mpKnYl1lbYM85RkyOQdIsYZr/d1hd8H
YrvSmG6ZbgTq9XEASpFdRfYqa6/mwQLn0TFXQKC5x2ryc/4PasPPquEOBkp51Uzn
5us/oA+oWIZnwsn0Kc+dVPag5d13sIuiHX8782dX2rUAwM7obhlTCKYgyiwJUFPZ
/rysXhMNcWJqJRab2E+22eiyBdEY/Z36VwOCO7z84VPu4FmSLC2Karadzio1UMza
nIT54ZbHdFCD9maZ1SlbXHp5acuUld0MdG9r/UCTCB8exAx76r22h/+a1sliprwK
KTpoi/wBKU2v/QLVPmrU9cBQfCbLqHI4z/NKQuEGLkWrpNLDB0DOpm1h5TfYliJa
2WB3RjkrVWtvTXf4kW10aMf26Uhmm7Vbu+GomBL/VteYFn8TWjbuLHKuf9UOSw2L
6NohDhvuyMqsDsMGgWE45akMNP+0icornadbLI+ky1K5DcPj29heldJ9fgOVByp4
DRxjhhRrVV6gGzBjCaUJOSjcrmyeJV5rcUtqPAMZQGmYUsQtM9jIOqf4hn6m/Otp
5juIDYN9CtMbaihobEnBhfDl6reoaPQ21ZRMl4C1ju//cRzDulwEAm/1XLIKNf8Q
8rHyzhpGljDabTq1dPkVmktSR8aQmZpwzzYU/93s7kUAKHoJealqOa1JMCI5nWAW
CvX3OWl9gNpCtgsAmWMdtkBccCNnrnTMUwKwx8OWZ/6fK3obFPGQfh3GeU3FaZqW
fSAVOPgN8dqJMDyID7umv/1w0g6799mEtmNuodU+ld7Bhtx1BQ/GHfzQjWbydTuz
pXvB1KaSWQJww32IwCuNjAYEWZzXWnP+fxxf+5DpYV7iB1MvZnGu33DZdiCgiF28
sKHMAP94KKHr3MHai858+SAo1qbv3KG4UMKbd6D3L7gWSSFZDauJFtFaR1vYnxOE
av5jifw7hu6v7DvuOaSSheYSD3HN/vP/jutoryFlLFDfLBvMFFbVjrdIyWTiYCdQ
q0hwd5Kb/xrYXulohtL+1vM4cIjSHmj8kt0tnHZT9sstfxemqsQgpqp2ppqpY7dV
5MXvjtf0UJstx2ZNDM/UIt9bxx7XKdGygmJ6KQSjjbYAdVBXPnub2UArRqWo6bJN
o8qhq+7I4jtdiGKARAWQSDkqxviGt2LinNKpLXTC2I4xhI/46JCJmH5pQ8cJV3Ou
b+5RSy4tVu1RcLMo8enjzUlSQh0D/VoNPmxP9gyJIsP0NenXXhndvD1iUOhlueNh
z1mOOPXID1qaQ0buHDnJgyD/3sk+PG4HkQWu2M6OvodnYauwGpPgtl7PsrxAp6IM
Qk4VRgvzpn029Ik1YxmsW3Rw1m8JFoPvsbbZANoiRfw7x9sNyRj/ascplIiFDSQA
0J9gjYSzq3mz9tUltMreRAry/UeWhuFqSZbkM14lj3ERguGOcMm1wfBI90hE0NIm
D6bDppLl4sEH73nqKHfwjVmJ/FWzybYc1R4suvDgd409435RWvjOnXGzx7KlGzAP
JC7Bc74aOH4aQBJanCHikO7eyesSB221P99+m7ApLGc81EN2qKm1HnGxweTHxso+
joXgkIjyO5Amt8v81zRDRwVIBG2wgjRHsEtU2Ufnxw255xlYf2SX70LmfCxy3xZP
YQKM7z5PHIi+3jAcm0e2bd+Dch4MsN+fUdcR2xsFg4MVdmvq1vKx2DW+TgLsQojt
cCj3nomRmZKbPlt+7rXR/kZoK7Aj/IarfVBjhBSd32QK4o9YErfDnfN84/lJkPYR
3ok6s77c/oQFkNp/jRZkSWNMGW5Ne3OmU0sUzsoZ8GopYlYu6kGEeRtBX+ZlEqd5
JBe0kLGz2LVNvS2tyLgk0JsHuK4C/rtQ4gWIE1HCJKcK+PIIZe2L8wTfzmHA3n46
d4LOmr8bSPeD77bJLo4o1hYJ4Idd6GPlKdNTNPHwZdIoOdm0ZW1Mr2loNjtNon3a
fEj1zwGCK6DDIYJYmsUAcplZHuQt63PvKx2gKX8+VCwJ4qL+uAgioFBLkPwZqguj
iFnMhIwWKbsL/q720i4XLsdM+6XZ3MaMmNWEUnEYygILQ8oJcJIFLWfaBkReBPwj
jmyiU1eyhm9HXP8SHSoAFohhtASvbBK2+BToDjXJrawh+xewx0IHXuHWwnwvKZNd
oDvQqmkDuKtcuCSxhf2gnWVbP6ayzHArtXTwbRIgKEH4J1F1Jh9/CfNZp4g4LMTR
13kcieMu9spHdWCFZ4Bpr4GLR8eJbPFbefo7bkytGmh+uiYhfYApijiMPkZpD8xH
shdzR/qZwlPN0yP04tBOk6bIVj7+LXGLJX+6gYp48tPnWzQxVXfXOnPgOEc8+zz9
2Md2aQWYdNM3MA1jzgaAYcLtNOv/2aIM03pP7ggIqhY+VfdyAR4MkF7l+ZMpi43F
d+1wZ4VxoOw9LVcz+oW53ZkxgkZPrAhwweIMGLJ16Z0HLEfvumorz3WO9CmtCAHG
3ICNBM4yrwTcXdZPvB84n8YlfFV3O59g9tzK2zLMGjiew+AAWooYrS+hiav08DRt
q4lDghnKQh4HI6B4oG179LQCVBmJ+y6QVpInY5UlmtPYagkBz/pPbVfpyUZSX/co
2aPGqQGKeS0Ui/0AvHHGnukI7+7WrqgW+UhFVVlaucep0QQJc17cMh58VtJepghP
xjxDU2TZlhEnbBqbZwX2vuBDyZvFECyK/e88L/Ex9v5SZ0OnyVPFWsWYCOo37C/B
yTJIzCQQL/v7D3qK3GmHY2IECTXwoY7FkKPTS81PTalvI4P8kp+y7cqBhSrhA9g9
f++bPpmq/O4g88pGh+Sebh4FlBBFDg0+1UEx1yQWcccmespsp7H4+WWxBC/VKeQI
9G7yaOB0ntc8nYOBVlsZKEkhV5OH1h++QSMmlfdF259FVtNyl1BfSGooyNFT6E3M
dSnPFsVq1KIrMclSk77nFti4MoflePTaS/2lU+z7SWyHwSjEL0ktGo+psbn2fWIq
zIN+mkO6nmpO7vlVZqd6XurEsgJiJYp9flS6wfCGwgrpTMQWQdDFj3EaCzk4qD8n
yNGBAlX99AzJHEOZ7y3mxG4jDJO9YVnO/Bu2D8vqz8JHCUQe5gj/wzDER6HePqC2
g0B/Z9+CJYG6jsZkdoDZx2S7b+aNTEZc5MesnARQgZ9SUvLUd3R39DLzBSLHw5mF
EOD53cRXuKHVtRYC80a7io8eo2Xh0/hlCubvb9hpUNjxbPXx+iRyUXEbrrpz10ZE
ws+fklOONkimV4h8+3XBcSPWF20XtH32xG3F3JZW01qg13Wm8CpOE8+ECWa+emc7
l0ihASsqOjXLSdJMTCRio8T3rrsNvl3KvrS6VjzaQ9F1kjS+E1VbaKWOSheVewnX
pcwtX7KlMvETLFNAxfuE2FmICGQdGRyYk2+Ib2Nc3VqDdX6BIEEEZfpnhKEm4V7F
P6SdrNl1H2zSyUT7SBkfqq23in3ODRB5Ac3BAF/4a+jreyL5AxQVt3fvnmywHmfb
QX6E9p9rPueruc1nLtPALxlXUP6E7qo6CT2JLaLtubmfAdGbKh2RUOKxU0ynMlNv
3wKvg2pA5peDC1bRtfzvtL+OEVgcoGJrFTBSluecoKQLwJhW0XXgXVZEVWZBL6iF
eGfUcrFtZIiINjcA7k0HFpkGYxTIsqD7zIvyMEBmoydftEUfI3ziaNh2aeZXoRgk
FJOHgdczG6KRfpY78JN4vNSQIrhgq4qaXJukBRwRO38JbhJl5s5c8Vp1S1YNWiDn
bQaDwa/tW8u9DnQ1L9F9BYb7nUgktPd4poBvVOZL+JgjV5h+q4uJarNtLBhHoWax
2ydsaXTn6nhfgJP1QV83iJnUHH2zgvyHGsZ95qws5aJ7G4eEivrbG0+k8m8+X8Xe
fPANM8cHOldIUduNO4TS0LRF6SRKdlmVQzsWqKqqmb1i2CAtImpL/gRp/u2NKdiJ
QVXs7lkAVtrEN9d13rTR5bnrFAMWspu+mxjmYT2T4JQpH37xdcY+qrKw7cNHS4Sx
ok5uavLJbiOed2RgdQFh7tHysoW1W/2iQFhBvPnFKjDsq5sB//b4RiYB8qBB8735
qbRjBeNkUgJ9Xqc2V6eHij17hYL86d8F681uub37E43Z5365HCtiOjp2AJnPB61X
HXw6QkvLy69ROQoyMy9jGv8lOsOgEi/r+sveraGy5xWkODuH2RcBE/UJDifgBOsK
392AFm8Q95ai7EkCRZYQ3q2oHRlO3qDIOYWTBmlaq7cAbJ/AEk2uZBxZaOKI2Xg5
/kCTY2man4FjP5sz1onc+pqiyvgdiH8DHWIJIRW6/DuG8HVu+grkto8ZE7awDw9k
axWi/iU/1JFPPpPCnvwssXhILI/boxFU02W2F1UCSci1NTGbC683TpxRhv8PB9Vg
OEMJL9lWey50GssZ2FVsCZ+P8Sn6qz46It9BPJYINKPd8kwZ88Cosf63TEdXtdrN
pWIi//l/PofRNmBJM5hy72pHS57c5kxHy0lRmRwN6VXvzYf05AEZMQgeZXOWROPC
cuP35Qgnl/NrTK/NxZpAx9KRq0C567rqZ7m7OeOjpglTU789p3Fn5kMAwUDQYfTB
jtj3Bbeg/JYEWrTEOtMB6LqBPoNvcNO17katpzvoTryYNMSm5QPlnz6yd2ggxYuV
LixGvFuPvsDBhOf+fiyMc18KpmkgmkefLvQftHlVXjzACxmb9jvdxbYV1le7lrbb
/LALyeLDhrjslHDr6HuPbKLJXKLoVgdVCW5+KIRwiwi2cGzfAAczAWusB3GCJ7gX
ExdrOfRH7J0naDlU5eLPVeh8oioNHNLqRym1rsw81nxA4ixS68Z1giYFTpX8onwQ
M1BXtKxjCGgv0IU7KFXChm97Oh94DeHUGlZTszmnJiyadv9GYr53Fhdvp0U3XxEz
7T+lU+6mtWAO19zOqCXt7dnKOg/FtOejdvOYHu+71M9tI/PqwtGfnGqKMk2OuDdw
QrdNG6KKM5jyRbjk8agWW3aYssfv4jck5y2Crt/c6Hw9B03tYO6ulSdRgzfqe83R
cF8nHnFzFLws8nTJ2O6YMBr/Dr4vUFXEnBD5bj1IWgV+qYdG5gI8PYUVOVQTnYS5
2XUpmewddHBhb+4+WsOv0gdzRBikqWpAPfYlsdZBolwa1PY5MUTvrrxEmcwmhS64
INjLFtwcUn+GNoYcyN/79iaMOpe/eb4oaodD2Jx5xRCX9xGqKU98sM0ktp54x3sh
9mW2FcRJqsPt8/OEfrzrwb1nYbqQmF0/BzDMCCM/kzxQ8Gvhi3mRM7brzUlfIa4B
6agPsan9Avu9kRYZj4NSv1USDVgiTDxh9J0wcKzwQnciHUb9o10sUq77SPpf2voB
st6bcykuUSfgezADD32HVUXOaXD5qslJXp/7TpevumqrDklhzSkMCtmbueyOxAUQ
JJe5Vnh1HLPLiTYPFRXCUUcmJVHGCwwKZR/2fTAwRPsX/I5ljl135+u83JAaHnoG
anZgWVKUJNMZq+qEPtDrjA2b5SqlSrvaEpnIcbXDjPVDaeP3KNBMjMI30/k8mtUm
tWCqEWW2dHOChW08G23tb5qQkDh5A5CRdlVzX0rq5vGSrrtWP9U3mZ/drnfBm7lW
S+2eMCb7JI2Y1I2fI1+8Z4QXBgzBlzL8BAiQdyWfbVFqw+ydczZbyJ4BdWsemOud
NJgwzPGgtEgjxWzF85NsYZktyZZ9dm2s364Jxg9Z/g6fo8BvAC/w0UkPkY09hkJK
CyZvt1nY11VRrXXWgtaShkugUHuu+lwtYgGwhaftoxB5jyV+wnGzQeCuB0HAdhgY
dhnLF86jD8BB0n95YUgRsDrsyhxGrG8e/sjNz9GNQ3kT/12Qz4vlhRhKnaE2Y4Fe
UUtIwU9/nIAYtOqeiSiVlWKm7LbclKW6sjkAkEQyVQBTbpyQRMjua/63tbDitn2H
Swy++enHBajXSKTrn7W0Ps75jx4CnUJjTAjxG379GcpCq0b5LU70us55z2PLjmXW
dirMN5YXfhPg5/UDaunq8Op0uH57L8DcJeiPG2pi5+4XP6CEUdKcLJnQlr+f8umJ
Kzoi1xv0XcIDAsO7ASoR3c4O+7V4OQijML8gRzOXGWWdLNW7ySDlCbALYIINGAtO
Iioskgac77mIn2wuBY/Ttv/ZGV/5/5WeSa9y9MyTrUjf9plyPsQKTdP/zwp7T9z2
xWorG8AkEc8A/cvZ6Vvt70BxUjHW7nWlBv+MFbUdn39TVDCThj7Z9Dbax7GXIa0O
j8qi2fTB/zkMdteLsC+Z9dR3EOSML09+IraYg1W6AAAj+Lw4ac8sQtTAloM8ylka
uTfkNZlRwUtSUB2APKAlVvrx1u48DXdP5rlp2qdqlphQz8us2LC5ArG5687Wsi/0
quxeB2I3r1OpS7cN7qtw/o6U+nIH8/BxwPZBfqL72DxQlAYz86PVduKBt3tr1uvy
kx0QB3YPtFjXFka/POmEUGjfZIoE7XGhdltWRpTY3vWVuEInSfvEFtkqk7UVcdaN
45m/44YbG8RjiMhC/AEiT+jBU8D3TvPVxiGMhubam+6nrdCZLCYHTAcERuP8NNEO
hCRSq11nKA0T/DxWxeK0IfPLMVZw0oaFT7nIz9L23s0gnPBUQBWTVYRVcQuE6dPB
Vq60YoX7r01vU3BxoY8v0SwMXiyPeQxGTeM9mh86FNCt3yZL4aTUtgk+Jw8hVrVc
5pGrq7dbjnNPUfAJHC8E/XFBQ+WSNKq+bxzMfkTUB8sRCB6Xv35XoQlWex37VaWO
kp8bquun7M/mv0tNj8NrFmS3/y9YwZYomnkeo36vE8DGRyxRJEhggfOZhugOSz4i
g78VXBnB2D7SA5H6S2As66C6iKdLw8yKx/oHormjem+csrKrDqEJ3mtKCgfZOoaR
Co5Qyl8yCgkczDUvtKSXgWN/BIY+3L+A/soEHocOz/jgeS0xwyDD8K0tbd7iOuqY
WG4KFczAsu3GpG3cXsTFvRW6tu/eYia5FSokGLFxAFriHfX4VtWD6VwjoNXqe7zW
4OLcvFB4EOUHFGEp32o+uCcsD3Kbgif+5Bb9twBewZ0/JYHM8oHTQkKfnmQF5J/n
0yKpiVHtZSETTGVQ7CTepaxtvfv4rcLW8jJ0JHIUSpk/cPmSLG0iGRsevBhliJYj
L3DTqGjEoORwCROcunohabyc1a8pvgTkLdxXGuiNagzUrF3aYP3pE+eiauiGjcC4
2cXLc4d9uAw9xyyXErER5oP5RR88BKf28jUuMSdaVfNzmUkjyL0szWjb4mbq6GBz
prbotLy1rH8aBtcfZKUMY27KxxFw6hPDlz09YMD3V2XDztRZ+UhtM29AyUVWqwoS
9yj1BysOCDnFT5B4g5rHm52TigBF+5DKteFKiX3b1h4jKA/wWHnT3swbYxQHKlfG
T1Y1vkGkUUXbEqmy/9r5M9bZI0pOYBdeDu4Zd0hJRF8yMAyESvCER+hm01ZO2kS5
sIvzS5eFm6TK2KLB4zKF8WyPutlxY7SbaEsKcClREEBCmRYoElzDrtjMUQCHADOd
fQNEyBkk6sberKUA54tthyzQPnbtGIzS5ucyFLdX13dX/1NnqinnL3y4mbevjScJ
j90IFwxDndFmH8TAJXHF8ptnR8rD2ruey6NZF9YvJRyjJAd6Xqsjipu7gzFFHW1s
+Gi+LRNuJ7tBSPOMFHOPeWk4N0HgTC7TZP/6oeP6Ln5C/gju2YQLJEOhMIMWyZoV
vUX0qYhpqkKVhvxcJUqzoxbpWSryaFg5BahWnWRINvbufTgc7pX/SSZ5OBVHgKbJ
0UsKCUBlcul3+qh3BUKygMYxwqTS+FKmx/4c5zn4aYtx4X8uBpf8itWrW45no+g8
URht5MD7rcaBNWxdMALanUw1HUFejHfn95eARkTy+88vz1hpf0wpw5Hgk3GBBWJO
uCr4Ud6qdZ46mm5zprNz1gRnnsGxrZ+a6qcahhcS6fLwxfpcUjmxDnjw8TkXOXV1
D4aJRr0zb0AXkPF5QLAXQKBuw633NSU4tSzaPPkR7NqTt27znpYFKr0LlctrUTBx
e0QOyASBmVVLQYNL4+eds+70V4j12ld3+ShVe/tj7y0b7CELUFMu0/lJ0LGZ6Est
r98tG06MXsVBJA2a2zyUzw9fhWI2SmypM2RCBobHoq+kJQFzuqKoCTjgA9tlxXND
qN0NbLCGjfDCuaRN15GsyQYvN7IT7sp921Isv/tKKhBb+UQxfvlzE8gFY0SoAVEO
Fi0UQKVZ48HV0NnSxPBT7XxcmtSbZ5G4ZjDUo71Bji4q0YSHsmEfvxmZfVciYp8C
nhjYn7J/C14/qOb2rDHFxFrdqIg+ah33W0wj3TpVNd5l8lihC65Q2ZMT5+OqcQNp
kByDcpWI2Q3rdSXLjc0xTiPLoLuoVIDVdepb7RPquA/mMNprIUGT2mudF2PjncGZ
xL94bHGpwrDAhObG9WGgjXgNOEa60HbQtqnaMkm5xcYzOyS+Koum5iocQln1orpR
UB/vdIK+0VwSmf5vE96Ng8VKm+n8IyOEVYFwzLkvPr2M0OTW0wrHI+vcNycrndWg
FT/URrjcttNT39XixQ5YRcm4F93UwEtVZNsfxXKhkddB08MAM7KbgVDjd4vZ1MjB
fmFJ7a6MyfcbQT5qnK8WW9MS+oBDZDsULic3/+6tlzO8hVy2Oj4C/fkqG8ZeZ+IZ
6kX3VgfzpeN2wx5FBp5Ycuih1hs85LWNw48Nqy22CleUL/CmghF2WdhsuzqpBqMh
m6KZZtRQChlQl1iekt3oLmhsOnIaLhMfsoP++QN3JRKYnauP1xldG1ni+c7dTcQM
0IDqadWo66kSVooLwBj+t08aQ3H91p+tjQLj9kwKjJXoQh4nElYrIN5/oZ+PjUm/
Uilh7ZiXe/WiO8g7g/6XWV77MQuKHg0WUR73SHIrIocmbRlCDH1WFmxbfuhsp0Vt
rfGxT3UFQo4US3+R/mWTnYEp+pdId3EgNyUkT6/C4A/s2bO+BVOnSogTvFSHx1iy
Shbp0TRzA6zCyWwkIP1YCuv18CTCKYhocRgtWg6rxb76EGQchMt9sdKiII4lJEwP
bkBqStPcChI1rGWrS59a256HJT/pHadGJ2FYvmD+/y5LEMxyErZVZIDjNiPhrECG
gOtRnVgOy8uJDqYlHxPL7IOCCG8vZoxh0T7t8C8htIkMyeutZ8JnxFdtFb5yyRN8
Vt9bzegN8I+1SLpboRTXbVg3GDzXuIsbr0E0PjCEaYSt5d6nKfiyOAseukvBivrx
g8b1KtwanDRmAdE/j80uEJ9z4yAeQmP+hdQE4gdsg0MD2rT0ko5vInRzy2piWAM+
mYl4lLm+AvgSf4iz4Vu29Ryi5NPUyURyFpNZHLc/+Ro3beic5Yqh2hh07thqJJ65
EcgCOjCPvgAqAzY/kxzugPwDz8NuqJWP/y5PhMwUuTJDeEa6X8ao+g+S9ZTS/ONE
sJnokIS+dWSlyqBAPYnt74njphnAxhTUcnKN32godkzI2/sxe3TCd3RV7bUY4wqh
hknRJY1h3+xt09o4Zhy0Jp6fVgjqyMPeLBmkQOEtsEBVjKe1CtweXOPU1UFVqqPn
T9W4uEkgCjZiAWGdqdNb5TNCVPu/IH1V9+tAGLVHGtKnTfjri5k9RZYLyn5lHsI5
UzXCgskdmVZ6Q5WVVQUGgKaN6VIQ1SaVy6gKqp8do4wTIlX1sMp68SCwfH1Lpc9u
fNzvReMOMLYuYDn3Lfm0VDnjU9rrRwhgvGYQzTnrNu8qz063vcOG06W3/N5cgLa3
ptmspyhuuVxSKZ/FrkbQZgBCkte34yS1fuV2N6ke9Nytf2Q6r8ub034xnQ3yifoo
q6iYsfJNiH1JQXkbKjPrYwNHXhUJ5hjDwtDMzi84ebHZ9SAa1T74MgLl16JNkI1T
GXrZapY0yOYsyi7wzkEVDvVBv4lWvWVrPNgTFF7SOq+RHQ4RHtXKHJs1p+3z0TIG
IkOng/6b+0uupwQuBu06SlpLZwPynuvZU1zjxW9DeziOwbAro3wlUoYTSVPVihdI
0+/orusKTSGKCI3rBXN2Y6+NLzfAC/M5gd4MRuLpejZ9XsJR3cQjsn+LkdVTAu4J
87tS1gehT/8JAT8MhJNeySjnTsPtnLiRzBKi63pwk0lyhSxN+EOrOBIpzlnqwFCl
ohHEMmOdpjLp7KTVAHUgoFi9nnBfGv3ciYeE/jVU7K01lqqnKEBjz+k4ORAHrAV+
v/Ek8hBuJ7BEleFppJegLkZIsme+JXixX06D0ZaXqZZXEV8BzTFqneklEp6dQQ5l
sbfHlsU8XKZA2IucO+iciznviOICkl3JW6ywyuEQW3OArZBbRGxgbxBTowjDaN3i
ZRxM/RLdBr8ZW5A1ot5KKcdIuRlo9NiKvxj9YQEu6HOMrum7TiOTmUZ+WBQ4joDe
Q/D7HOFv6lvck10sM9MjN/HqaCAzpIel0h4I4p6sS87nLivWD10H/byMa0qLreQD
jkQdQ486TneF3H3OYkvKvUR26e7Fj1Dk8hcVaEH7lw6w6a/bdiVErhreoG4m4Y1f
OAMHxxi60F9W46oDU8bZSngJKmp59za8qM6JDMLfXVYQRoprLGn0BZ3EAdzGdEcr
eb84jHnGFL7yu03LIKtRUznidNjBZkwYTeaMAcOc+r4+S5TSbkee6wgbKX7UTxv5
U/6R0/VErtTIwUOXkdJKnFFwL6y8kxF7VcCG7nzxr1lWoLg+4+eU8bFGcSDjmhpY
vAiHMpnuotS83FvwxI1j4n+1UD/oh7B+wY7LUXY7mLZlj9dRD8j+rMwwCzgbi+Rd
4l+vPHsbKBvdNBZ4706djiJVob8dYVnydtzfktvGc7mgapmw65GB4VsNx0kAH5Ki
/oUG4QmXh4qR7l1OQho3LjT9N6Ir84BhdukzCwkxk7BWi7ulSuuhVL4djHOIpmVo
4rJCNQ9nOBK71idBMO3lBpHqBLp93jbGhJB5yRjOxdC5oQU56fH/HUb+63I4rd/e
U+n0Ib0Fk2iLdVoHlMFzI6Gz0TY5qbct/x5AAKBXQDjAIBKfacRLFXvIx2IOQ9Sf
lKzzdr0VgTbAWYdsmkDA7GdaoXrlrSivJp0zKZJ0d/xCu+7+W7T9hXs1JJYggKia
jnEFNwlPTXDdoVhMy/xMQRD9WGkV+bBdwhYpTR8pqDftwg9ytb5S+lPpwZYLibXl
3Bk9CLxi7sRcjllFMiNxpHusuxllyEm2N72yHDcI6ES9MDCeJJNlPSWBjJ7NqxiB
anDW3aj+aB/ISyNO5PIDH9tKjYK89UgGi7b3dRytlz1bd+y1gfyT3gJknacThW39
SQFmc0KB45kzz37mOvAjNhLRe21bs0eOPfoUBKMqzliQcVhMVSEXNC20NbVzsPKf
gXC0i0D/M+gK9BtEPff4SJCQZa9bypztTrCWYZp5JdDaaJDEtAr8EMmOyhJdZhy1
MM6B+Q/HLaQpHevsdQz7kuuUHxdfDvul5dsibFOauHe42Q/2OHuMlzicW96TcvCn
o7u4ZvRlcSgZoq4CTSVJxoQfx5rFM2pjqwhYkIW6AT0HWg+Ntk0thu1g51zhHmnh
zDFHm+6sBGECkedAhwZXWVjN9JQ76sFsLj6GPTgiTyP3fklZMTpLP1j6tAlmKDmd
SLoVFivQQi4Of3pnkfFxt+NhAKCRuPlC7ZSUBpfKKd3LfojoRdLSalnIaPEZ/Zzq
mkZXinI7FJ2XGqvpSYX4YAf81fROovctohrBmJxKpfpBrEuiyy61J0s9t3UY+Igp
OAQ8jCw/C61Aaylu1pvw6rf5GyNvNvhgo8yw6mPCVSuOjHqsoSOFRMy+sXFY+CTS
G39x+EBqHzWEZEijUhjCmrVBwy3+tqEEMWOVPh85x56NlewamZicUvyivaEW7NGf
Rtuiv7T3SiBoc4q+NwfpJ09dIwLjl+7DawUMVm55rRoEZm6tiHR1OokA0dYkMfLJ
50VhkYr38JHeQ+xHEYdILoZy/5hhf5kFR04jkT+Ulmrmyzz+nVXUhpnIBif5FjPg
rYfijFd6Y7FVeqwtnLJrJmekaszD4x63PPCtMWwcO7i+3gQzXETQU2cqq/k15nGG
JQVv4D4xD4YJlWcLHn3TXzm1LB23xxBQDGqDel0agzrTXzeEluvERb6FvPlZzeL7
E1j5Hy0lVXlYpfNS9Ctq77d8QbhEaXG7dAi4gYTbJ3oj4RYWSYR98j8Vdd+unMi/
UdAvsNF4mGiAnXI/B49iPeHeeWWvlsEKx4swAeqWyzHmTamra+u8sSs90QRUTTFT
rd/ASLlEsFuqGXv+tWHeA7lyDA8aP23sHH8YR12TdVQxiJE5RPgOpow1w/AsrwZI
m8K4jh6aqauU69qeshHKkZYkl0ueP9+53spLuepBODij3M7fBy76JgCW1ECpWBsl
DbZ9H0786NKM3EcMWTXdsil4kwtH0qnAkMWwRB4LTbsrEFcpv8dY8N2+AVVmWZbN
+/aVnsUE+OHS1SzgkVCD+cF37smgZkrpb+/t9kJwf3jDBnCAKnIMWhuyIZntYKRs
igBHXCdbl8fL8x9u4EdPA4geZyv6eEcCfJxawEQJ/Lo4dAYyl9Q+fXVGyMugvdUh
KWyDn7UlSwJ9Ye1Kfu4h39tIQL5sPEY7i0RMuDgs5QjSYNVPUXdN+lhU54RcBEru
p7i6p7GKs05R9zH4qnSan6gTFKAColX8YzVU6a3kvZ69LE2xFQiZ2e2g93GDfS+C
G7pF41kV1OCeF0jUOEyjEfsE2dHDXqwZml6gVd71ZB3e5LVJ242537R0LHKH3Rr/
wdkloLEenydVw+LmSxhYfXxmdGVwZ0cGakx6FqoNBTpaOjHWiwejAkqK6ysJ8wmb
usRumtXFy/Xk2FMpWUvR0x7Ll5HV6fnuW+O5Chk70kMxnv8uo/i1Q7Dz7zp261N1
8YChaoBXHpaGOzF2rVdodyqXUhaPUIvtYYb/W9R2vH8k5ohRKhNUHZtaDjUsS37G
QtFilHabEbbvJ6OiHYWAz5Jq7hMUOYO4DwXPA9qvYCkEM4q9s10l3tPQEqYWnJc/
N0p8laFgge5uf+d4BUPO2EDdAJx9fY4YQPmmT4JoyUC88ldooN1YJ3uXa7WZXqgf
qsB8XZfLk14ZVPn9X+pc0a/Ixc/CNy4oShlru/6UVZqOypeLp1X70udSzBkFlQM2
819DAXAG/3pQBlru6BLqqDStP3RemK5QzbwAlYDjr88oYDe7pO86+bheYtDDNI8e
GUVsZ60Dl2zCFtA+MyeOoLmb8rVp5nZnX6mbFEeFBc3cCnnJWa7ZbV57fVHfYXgt
DVj//9JW2Ro5vlhlxrZDYKSC7tqt0afXEt+uf/ps9saogyWM5Togi5Z5wQ2FFkKT
8WwhR8gvNBN4r6/n7NLt8PzJTcEuRGUQ1copSf3lVqf3YMN7TN2nti8sS7n6IPPf
L9Zz8rwzSTmssBqcByhXRHWnchN458snweYydioMPpu+tZ+7d0lfPZ4uZ2827oAq
1Y8IOzvBrD/1on48iitV8BNSe+fSQpRRQTYKtL3MyEOTmn31+6X9BH0iRSZpdnKz
mOftmsw6UZMFwGYEaawkkvwFQWztsCTE5gVfJAaxoi7XD6VpoWW1bvo2zeJUmzdZ
nF1+Vc07DxweT0w2td78KZqgFpcySKMsv4vboIpdkyzf3WnUnPH3YbkxFiKr6YRz
Mn8HbdpgPbOeG727uA+ZKl7IMUsfEeRHYKi4FNtkJMELU0I1nKp0gtby46XT9VY9
s3Re0+4iam47/P35ddgwGunt7OWU/ESkqS/jzfXO5VL3oKrfgYMkE3uzIMD1y5Us
TDn59xz4+tKv1zLcyZ0blhKObWyzw8PJc30O6bqygviZOeMO/wkivNlNfuftZhb/
g3u/yLRBDHjpBs/KKzZSZ/QOt1Y+QXk70gGGbcnyIbf1TXziTVNhd+zuvw5ac4aK
xR1QghBIY07oPtivrYfFZS2nVbA25stmgubuiv09oFwKPQdCOSKCz+UmVlmqAD5g
vy+FkFqwMGkCs0QYVmkfy96NpEXVDybloP6cFw0dxIkDpaisqCx0FOcAPfY2v2NE
gBIiZbI9/2Mwwi2nCHSdLc7MnRBE2WF74L9qxpmdC3u4Zw8qpuqVuOArFFVwqzOw
7VYMxAhLFkAMZ91Htj4gzql/4SuBVlWkSN+Bv8CxTnOAEDAEdxwN8FQuIFyzxCum
8j7yfDqM1uHgcsZXTQA5OHfLYpJ6oBJi6P1hROjB8iC/5Q2ZvYWa0GD3bR2OnQLr
okI0x8M1QhR2i3GjhFtNwHFopKNNW8RCn2abJRtgZvcZraKhzK01mFUIy6JHMOIM
Yit6OGZMUI5EfGjHtWNlYanLR1EPPz+yrp0RN7ISANRxFNIubaURnQccTeZLB8RS
+mtubcwPj1y93DVqhKhwcN6PBRrL/atjaeGg9PgvnlrKjHg+NvC/2zgKVucBPdXl
fi/X5MWPXMl1buhxv0UG0sjlIEg3+ZOyFIIQzdTXKqmZoQio0A3iqRh5eBxgk8vk
4nv21GqylvQyUxTzJ6JfM5KP4HlY+wjBNRXnWiToKByVf2QQarLKans5t/R89PVr
KiftOy5qFphq0D4Z8erfYRLSe64uWPCx/uhGEOCKxS4+/AKdMDnKycf7IMO7bF/F
ACYxf0VcP7wVxWbuTQuk6q5MLgN73Np6NfM2FUWKgR+4AxxN+RLkYuMJXE/Nqvo1
LyqJtvoC2p52cJidHiCbW7C1OVmFNUuqID42ewWUIGvV64Fhj61KBufJgkklSkxB
7/eXd8RNMbZJnb1EREcJJ79vRUXQJLpqucm7/jsYIMmlyfNR7/gt1CGZyb4QKTw6
MhzM25cZ4eH+fT7kWGkOBVUZXGaID22/y94dOXxqeOm0ophHzbHceiKt/kN0BP/D
iq4ZO9QhkXkNg0Flxw0JVIsPO70CGiFKlICkf4zRe/XRYwDPSEfaB6DtNCxOq4/8
0YBD2w/J4cL2vmcnFKah3yLvcBsoJpwHtN7ORpz1LRnK5yLlyFIPAn3VgXlLg7Ni
+WUs9JbD1NloI97NoDrbyQt+mzhfWP5e7kn22Z+bO+FRib0OFY4KdHyR9CRfec+l
T2Z3RK/VEK8DsifQ0symRfwvjhpqt7GPxj93KrRBpRDNYaPIoIU9FA74p3wVnRIZ
hczvU4flGJF7jQ9oW1ved+GmACPdMVYku/cBLgftsqRlaKHgq2Lf3EX9uTTJEWmK
Y6ou0w1QYZhBa3RJhOdnGe7j1jP+MopPa1DsEMa8h+/hoZ6cJeWYvWVBRyJKBXll
aNssT3cZRYkID40N6ynA/R1VexzeQ+6XWCYd5DTUa8K7HDMp+SuKAErc5keVILwG
BrIWoojq3IXQdcfPklHRv0YstIQbkfU6J2UEP55sTmjHG7r1B+pRARp/4th8AFsO
N66XgaxboaNDB5o+rknVVw1KH6tMsxSV6J5OSpy8Rw25Hwesago0EAJc4XLCsMPD
OrQwLlcjNSCgGfXxQkdkzvq8c+S/2fT1Xo/MTbLtjUDqgOi5FgYTbxWIm8JhAklc
Q4RgjmqESPRKnVqPdAp3GVQiC7qq1gyntpTKpOK5d0gZix4kO1VrdmYPMGqyAAcj
wTfwWKL+XyFdemVPdg7tqCWewlPvq6pdWL8j8TiB4mcFZaUVXWH7yhFQJDNv5WcG
8RLFevQ/bIkZRNvZFiUokNaOZBX+7mMOS+JR/00tFqZa+54OK+5MerIKF3KMy9Zx
vaN7bxvGOFjjDyzWZQJFNNBBbQ5MZlVA1M4WFMPj5ij8fp9NKuzev6miwn7pWOej
8l1BpNZn8Ve3iqSiC423tgoTfT7trRDjTWeeWCVHlVfocgkZlr+nvwlTRBgsrghu
VHN77khhAowu77mVaU2yedC5xQUIWnBL30hY1rG1KNPAZ0Evxb0q+IG9gM8H5jhK
VgtLFhKu8VgYdjjG86GZYSEv8+9KhBauZ2qs6fxgT6FFb9cc/TwhvZRc0zaaIkJY
oDV3v++Z5+bcoP7OvumKf/yfgS7g80SEGy6PhvZOSXv3DuUZ8kbfLUnsmeJSsdEd
rCLiEL7Oh3cKMzb6uPYwus5vEFGEDheUhaghkl5NDDFBzkg6wrmz31w5v0d6Cifn
v1+nGRjo+C7NcYMArbbI9A1gASrQ56czmeAZ/FpcDJUeeBeOa6nbOs+U9L1HUsmN
BchAd4brSzk4VJW15MOGZjtIpa1uss5ab3ZiHQF7Z0E3pIJZWtNIur/HvbFTzdmH
gRibkaHn8wwtdfK4JWlDAqkgh18YzR9VQuxqgJvleMK4y/S8uc2zvdb/gX8AwZMP
sXZOst/9wTH7HBYztSh9AAU/4fFfgnAZrN8G7TDrkOg8TnEK1fSPdHKig8YjLy+v
ysiYLwx6FF5lZ+cOENBFSJyqXT6lMItxXzojxGAInswRwp8YIZEzeinkC2QxhLxe
xxMO+s/HFZ0f//ttq4rgeapXq82mnHTB+gtzdDk74flbqV/EYsswjV1ZH712NLM8
KSGt0p8aedCrTQ+WEjwut8cTxLVVWXYWk51SJgl7Pt80cTahEJ4EVexKcLaPyFIT
7EJyC1DVCDqqqCVoHN0KH1YgMxCFSOl0RYVh+Fcwpivh1M+9ddgTwX1u/73EUmHf
whxGgoy+AE0KLLh5oRfqGA29Wh0IjHHIOpje8xB+aLOZ2AYuxTMlp/XKEm3VsMBs
h4T3slsmzrXtM2jR2vanPTDET0Wyg+nYH177QRE9ah7Qse3CQ5puvLFXBS54Wo/B
3sV+9yk+gUykwSOoBXDtWmxL/nDnLViMYEhwnPgIYIOUvfDugLcRl875XeaKz0C9
UBvWEubfOxXYeQGgCy314hz7ogZVKWr/h0vyPdcdfMZRnqFRXIpkwrqrq9FbiBke
BM/F4GYV1N3OUflPPBkwii/Z7wnRZR+AVwp8UZGwsQlgn69ughxCHTWxxxRAB6uE
dR2GBUt5D9lzm649K2tNSHt+EnQzI0KAEaxJV0+COcSfBf13tmYZp0M1/d/YOsS6
WNDTxTifmzjWaNtGMz2YAoY5Y1Pr3O9rOHP6j+bEcV+yWfruPSdDA+kJ+rIUuAXr
LPiIXxaz3bjwvJ2EZTzCQRXHX/NI7rC+LHOig0Aebv8hZJB+PunRU9+TW2fWh2Aw
HuMQ5GWcDupmoO0KZ4I5IyJm1EEDWZSasqYts/64T/wLaMldZyvKYena25F/2gIr
ogUR3vpj8rQZEILlOK9d2ZoGyYoRKQ+W0syG5mcKMrLgr1aFzvGjmrQ9oajpaj+1
+Q5F/KfYr/jTc8wUruTOxDRNw+Ce6H1TMav2b7uKuVLhUH/J+I2e1JPd3hUjQ1YE
eoaq3uS/w2an4ZJ1tZwhHMjcBB1K+d3WQ9yGhznzE36CS+673yUYh2iCg0fCob15
GR7iA50rvSvYQtVZNvNGd+ytM1BK6RQt2upvG1TFM6piBZy5i5xB+edcuxtBE3rZ
O32ZOqcJ6Z/JH0LgwZgmlHV9CuwZFcMsLS1JtNueqQcr/YKWI1WF7pIMr1QeVkuc
kw2niG+kHnl/mBgMdV2Rwwemff/V6m+ro6/WxPqZcx4SIfADNJWgbIyjQa64Q6tz
Bt8bZk7JQHV4GHmrWMsGfaMa09UtTaoMscf2pYrPH4QqLsuYEGLi8MztvdmQyi+7
udhr5w8SDlkHb5CeDWFtYaVRA2oZI5rYbaTQUeWEbE56GLNAgCoKOYCMQ/sHhDNE
sl1JlxTa0H1fiJKD0cvjlu9JZLxp7T5EUqE3w2AAM08+i2XGirOJAkEC0icuxx6B
HNniJC7ofV4EJlhVc+UQKBuLZVTnxUGXkn+jX49aJIjx6vaKJ+eg9wZhu2GYJIwn
0LrsgdXCM2YjuvaSMjlNK5UcSUig5DnlN3oa6w8IEMMIYKJ4rmuosW0UV/yX21Le
9lStwg+uWxjBVZV36F6k/epBzBN8mQWhRmGtjlI9fQ9RhJQDd72azENlY/IKuGRo
AMTvRs24JEmMDAO+U89yKw4KMY+FQEG7BGDzvCUzIu3B/2BEArX+sKeo/NDTBaya
fmCVn1xA8M+q+GZYeFbdhjedmJRXe6rkN6cUT/sOx45ymlEnkQBoAF60WlTIu/6U
tT4Jlehwh+YkP0xZj3WekcXi94qQIiJ6dHXqpw/kAUBMjxRZWDreZmM9XEyHod8z
eEXvXmsvx/+d1jBdDKQIdrZIeYHYX9BKo+MB0Qtk+uKUny9VGAqETjdRX48vSIuT
a6bGRZYbnaOpeUKYsaG3lD2Y0L15hrcxdEm5NS6aS8LDwuUrj7A8YfqaJeYEvjAC
3YRw0CX48Mwss1+X5SAE1is6XFfK1WdPaxpVBFPV+lUwuhebGeC+Z2yAmwsY9TQT
n8RW6C219A2EF1MfeJhORuGgllQTcKiR0DIIqhNErhYyrWextwPRhMi746pptxOK
vyi97dqz+SRbYXd3xq2bvgz9Oy6y/GqgB9NQrAUFbO0MMAdG1vjXCxV4GJpcFE9a
axMFLWtay2MJvhkymiEBcd7uiXq9NBQhjbnEGRn+YEVH4ld2Z6ZgXw5nnRXEJ23J
m9eacclAgli7mItbuE20+5l19czhpgC9J5ULfEBOPMt4n0u8gDQKbgIgTdxiieS3
lEz52kQrSo7hBf+ahlg2ec2KLiI4kv31LA6ZCmtUZBzSYd6djgeC6BwSNAsfG7H2
yf9s5VaFjCPqImtiWnyVyAW/+Caod1s47rNb6C8yBePitZfMxC866RddGo8dRMor
Aq73e7SIiXh9tjxuYa21O4z4nsSAj/IZx95EzznJ/95c6X6of6DRl/a/Vt1TlYIe
pL39WCPx8Gog1Rdo1GlTutwiBDwNhfjSwgULnaNopEu+yfveQLrq96wSzQzuOJjX
TGmaK5WthzS5wLOx4H2P/ooIPA6rhobKwk+wHqGSab2QioPNv+BLPjJvEA7B8fRG
iL2nVkiO79KqkGAWjMP3efraD/BO7R55zJbD3XMwOx2ZiIMPQyMblqBEI+fBpozt
6hn85GsOp3EQcqbTcR4aPmMHwLlE4C4buTyO9bQJ09UHeU5WaLvIH5/9vazF3s4K
pQXJZhUVPBAd2bUmjhcmCp8LKkFBC+QKGZsIbzKvh0O07miOiIYTzS+7fj4Bfzz8
uOPhnuQZut1Lt6bpXgqK/g17JTc+uXo0p42XShgLum7TkX1Q8n+oat1zJzm7auBF
FcCuzeca+yZnEhs+pbuw9O4s64GxJQ/lVjpshTiZrCHZGN8+aSQ29F+bCaAf70NS
17t6n0GoiQEFJo4z3VmyebatKgFjJMX61zvnXxo4PYqEvAt3n6wXGguRxcOO4bQO
+lT2N/YCdEvcF3ttXbWPEfuRCY5yTQ1OVSQA/DFEdLlX7DK/ON4jmvQhlNVc0nG9
kL/H6ObheB+dFTBPi/IhygV86D+dg62Luk20WQvmV7KNTqRduObOtjLsU8SA14Ii
T/OUtdB0Bbx+X4TsGRohtHkj6sqlbkyAzvXWJ0aHFEqJp4P3EdQsHuSCZxjkb9A9
PpEwljitLLsl3Fe8MY/SxrPCNzindTG3p1/rj8Js5zb2g3eWVmStDlHTvz0hE6UY
ptb1jgZiXtFeUDa+ThCi8klcCkMUUHhQGT9U8fkaMBXI402FyVi+79F42wgx1N2l
NIFGw0rUzof0TpYal7LQ5ANj8vGNN+NNiU6mCTNqukVc4OReK4Ua3FLitgyjIaxU
dfJrogPllYIieCsd0j6XvR9o7iSMRzq8cDpp/yK69OPFc8QVVNYJ2muUm8oCIF9d
AglAKEsn0NbfmajpZ+WVN0/uzo0xbP2m4ctBp5+45K71gy71dqDnJtKVQm/nN/Rr
oWfLDYDMpdJcM6WXt1XVp4bKYzb0j/bGjVOXcfdwbGMDbHo+T3FaSmpWUiPrzS5p
AsFRJkUZbitPPU+HbbZ0cUusYP5jByVr2mRfoQs502MHsgEVy7kaEI9Q9XcDn+TX
PsUPf2D/44H3tVQ0R40EnqEMXl5Raypep5+I5Txxg93lNnYxNo5vZcBO2Lft72F2
zqAYmev6uLP3iBBt+vshfS0XdaPp5ldLdT8LVS3XvPzit3rfI0NvnSVdYvrhZB+/
7qBROPp2qR7UwjOVpfcfuPoUM94OdzzYbqLb98/XQk3Z2pGRVC+OFrzSD7JoVLGP
F4YYdayU6dQO6Em3ztyJaZSxpdQUNWAuV1MTq5T5kii7RhsUkuY6UAkpg01NQud4
w/di8z2nPS/kbXks3JfipIe9qN0owi4wqkVAbwEzhqyIzt20LOGsJj8s8pR7jtxw
RSdZSn8d5QQ+LyBGpLFdnbjFlJCo//Bjwv68qEZJYR7/lsl1La5gL1Qkn4J4oV8B
nzMffL62ymC3k/sqCfVqqjhRDtM3x3qR29dY1VjyMKdmQTzo6VL8gIf+YmJWJQTK
oraV0HMsXuuHx1kcFzUsSgWP23LpW5zUIgLGfxzizEue5EZ7haOqyxts1KGwZy3F
gASieCkLtZbv+EHfd9h22B2SKUPHNne9H/GL1tby2uxE87APt5EwQKNrp3CR47lS
MkU/w/Mm5v272qSEQrwSjIFgA+z0gMOr0Ubkvu4749LwBZScL+ucaYp1veT10D9K
kTq4WGQDTxiFLvMwn70hZRCoDdHKbEwXbrkR1qqyyqWuusWfDyDVY6Ieffgo81hi
i0mEArl+7kpThkjs6VZLB/DExVwoxq+eEC5fmPDQyjy6UaDWLcLPF+HerEnZeqnB
FnGAjR94t6H3d9+uiP/1BoRiR0/K9TaFoKhqvywyUqRmJl81mEfaI7ypOIpoSCyd
smW/WR8ia/hwiwAMp3QpK4HOAgsBC93GWfVVb0vaq9hRDsiZLjobd+IcidXad1K9
/yJKGXfVwyEfvFrHsndwQ6BbXyg0x/JiBMAthKC/qYxzbCwqtC8YBFODqkg6E260
gkzub3pCGyAhb0nK36NitWz/ch9PX7Oa51uDfR2zPARpRRiMLg9WrsFOjlJDM7Ep
xNcXxIJpkq1/N9HJhuqco+ZCmp5gv5awFf5v2S21RddSuLz66hTC/SGNVOoKtVy/
TB8dl2QyakrzrWjP2gPq71Eh6P6gqiYIOXl6VAACjj8YSXkKXcOrbjMsCgD4UM15
eOqm4zp91cVoA9SesKgIcoMcdXMCCaRN5/AJQGxEFR4yGWRxoRQXizAtW7OIatrJ
4b7ok+/zZQ3+JzPtfXMLQDodtMws2Ue742BLz+Vxn/RJ1isC0cmKUZbmevoPixxJ
SLUBgdOOPt114XSkHLWFG8WnL3q51KwBfbNebpiX2yRzNetjHtCJDHGe7S334pjf
8epH1YaP4MJ7zz3aaNTqIi83HEhPuK+3akCfSUn+++be3sbUEpaaM26HkkIvNp0X
VozegorK5vR//6suj3JlUKz7i7dVS506v9lQMhmETSBhnMKld/PF5Dz+uk5KT8Y5
DBab+8iHVoXroe7VWvbVEKw4WO2pd0yrPKqRHYqRS761WunS+iFDXHkmgt5oJFPJ
Cqjr2EI53Q4gi6FsvU/soI940XqT3+kia/moT+xesOCakQzmSNSeM9QjdS7yOLNT
rwW0heJCi9hiH7o8ND38vIdWELkUKri3UoELH0hGkHUhDu8EhibvYm1dazL5WsaQ
1E9rIjR08XPn0HYb3Vw6F3EgtKV6vys/jjO99/LH/KfSHn+Fi2FZ4BfKymDr+mvu
gljfSpBlD1aIflUprZxns6DH949eJhMx7vlEu187A56rLGLiwhq3/ied/md5uYt7
BXP0LohvJAG1Rwpra3/X6+LR3qCDmlYoFO8qhwhQbZG1TQS8wbML1i+zYUm3XXmS
jD0Mx+bvKErQkc0sSmoiMe5/86runQalG39vxBF3vkIoYvBO1BOCL0Ntt+xrNRuT
gHlXsCGNOybVPn1A/2pX4WVda6DmOb2maTuhGkA37Qv7RRz68wynKk4x1cRdXc4r
rR5D41MmYt5CtFRKQNhdfR3Unm9pl3HuP/44QBTD4HPjKGe3j9IUm8j8PA90V1ty
zfQ5q8fmCY6YQKVDb87+hONCOUBy0alHnosZAy9aKzFd0N63qcwDG/qd9Yd0M98q
/UTp/KVSpLa9SQziKdT/cbYF6HsTVE8ewUjzsAJ/+B/nKokVSB8fTKCwXUwNXoAo
nWehE38eYEoa4A7fKrPV+FqSrvme0OD9L26FtWeNuNGGFIRz6h1ezCm/Ou75CyjI
m4ZvGcj1OsOwE08c6ERtZRb/c++pvcI8a4VG0XxFT+nGB9plTEfV2qK3ltYIJfcJ
SThZuj5LuSRgKRZe3W1EJCGdIvcySbX9jFxuDD1UuYif0/DK2NGy55VQQW53fZsW
3RjY/tGc2nRR5WGWnepEQNWKipH6C/u2ITEetm9fsHDKK1haiyBojvH9vI0PA/6N
pfIu5U2piIUG0smzrnAK8BN4fNN2djZCiyolH4oIewj5W0qpd3HB2SW4mgCvEihy
3F7aLnTeX8cjc/gUYmcOGfGYAH2i0KnPcYe/I27ksDuFQRmPeJXhho6Fyk+o6O4R
MPngzRObj4/F+XXMFE6M5xPj3fZaR3DaRg8G0OMzawbHjssCzwp75qCkZyDKIgc5
l0xK7cLhllEHSKkBidYxOP9pioYhiPWXz1/IYB4qLCtpZVDr9glSw1Rq8B76Rr2J
cTGytY+e8yNr41hj7aD8dZb6qKTfxPjkluxV0L6h8e8/Scn1RPIIc5aTrQxr2Ddp
S9BPdZfoA6OzBmaxWDBfU3waLyeO0R1yxQBulr42lws5/5icq8qp1WTJ59Mv6rR5
k6Wj3lkGTJFqOtoYgtqB7M1Iz16d7NR4avc0IWtYBenpHv4yIBCMC/hdjyhYv+B0
5hDhtKD+xDCB/W7vvN0UyRy0Ohu4b1TORJ7tPa7jPa+R3CYUTZ0ipUgPBlZfoBwL
QeN8S9sohTGIQQM9llg/E61bvx/DdTES4Lb/L2lrWAgPTzMlHRpTO3l/2EUnhT8e
DehdicssDS0EzbNP3FBijqty7UrUUI4a6OR13ws18CvxXT7Ese2w8BRRxkON1/4z
5O6IbwKCytyygWEyyCJQtRZ1aEn1jI+XmpJz4V8/BNQnozIPCA/Oeuc/ZT7LKMP9
BW2IIR0dfDAPs9hWbA8yZYziFkqqfDQdYXNLQhWGPTXdbPO6e4Le2nnBDsLpsIV1
06hEDKnv7BE36U/T51suSYsNzQBMNTC8CgKP6u4OSs3cEraEpmkDIGiem40cEdW6
YVJ26RIusEsqVY0xhVmOFc84o3kPWXL0erMbNdeQjtlpE8Xj7A5ZYzAHOcY3bT8O
Jb/ntpsMegHUVSbcn2HA9nJ8yjR50HaXisfI1DIL4+JEo+uYrLvs/ZP+jm6EkmD5
T/aO6qoCp+zRfT8kKfQYHmo+XU1Ju6XZ7mt/f0G53psIq9htjMTUoZ/bZMjL8cO5
8QBBQ+FAop+mnwAaGCQeEYSZSC498oSSWBNtsykS4MVTb4e5RQTz8iKqdJjY7VBU
DBb96h5FHz/th34Mgol68EdegkbLxe8Tp+sFCyqFNvvJi16ezDRv4qWBzmh4/sOM
M78zGmHlM4Us26E6jpWrlXVE1E4yvAZZdnOZB7V+ZXDgcBc5r+WjZ8tqxYnMdVX6
5kWb9KGmP784Okwe4Vv27OHPBV0q9BAoFq+7IFKWgIJ8ti4EC3MzMDxmVrW+khC3
F6pD30dVwYbI9DkfURrdBi4znN/DWpRG+UBh86cxj6m0zuw0a1PUc1ns0yPpUbDE
ETJV1I1jjFpXnBrtnLvuArB+fhoifT9/WVEqKy8xOlxzAeaBBETe2ls3QBvZAewm
C+ziLOEiNQaEChf2eC3qNOH5nyDIRCC2EaEG6B3hL6f/GvVoQ1AbBlcpoal1G4u7
3T4Ncn+GOr5+3EOE7AfisMh+sD3rri6NtnqBj0t4WiS0VMKnmP0w2RhoZV12lhuP
0SAGVKNgxy5/BajwipFsXhlCPxV4fY7mP9fDdZ1P5l3iewkY3TY1F6d/XD3az85b
J7EOqdZWE/zEVY3UXJQkT9h8kRepXIzBBHdvAasTCgdUQLk3/i69kUNBmb1a/Te9
heCXj8y+Bj7CFIRhRPBbq0pe5Q9NQvqXJ1GqVfUuRbx8GNM9B3sKPmbjPCq2Syb2
9lMjf4/noXo6Bu3qy9e38wHdE9IXz4StY/znHwxIChTpqrbqMCSSNHUpaZ/kvm0W
QxG3weqCVUKpV/AF8Ee94DpriGU3u2yMA9d2jfGegTr6jLFdv5yXoaqfnEGYJ/FO
RMtGIYkuhJOk1nubCp01kX0kD4LPM+Heizs8ORFvWTNSsG7WRvLebYgkECpC1Jmb
Fq387+3PApN9DMezBK2L+xSPjY0OCtyItdHmqrrMXwxR8AzzMTSPrUneepqb0bc/
Vd+Dh29+2Oxg8IA+E0VkWwTxUZ6ua4waGGsv4k72QJK7mTfOxiYHUizx7+uthdu0
LW/euux6ilYZCBuRH19greYDPs0gpvonu9XkL+qYvrKzVci5Spce6K1k6VkCmsQ5
vXt+H21XVsGywGYfgkK3W2S2XypUcCqlaNz7DWYHQ69WFk9p2zQYt2/NGoN2/smc
vKPjAtGWfeQymdzIqWCOt+ekNPFSXMsrmEkOF7HlvZZ7AjVdzfwu5uwQjWQI/hqP
bgSkPbFX7E9x9TuRCdjTA3uw3eu4qqGsc5WtONlsStso1tSF0HWG2BRJKdFLA8eF
+ezfC9v9uMyL7j4aL9JzTJqfaN8WaE4KXfO7xUN34AKCH0DA8BNFnXxWgQzh2aaR
Na2tXyldvzVHgMt0jQHwtH03D8XUC+urT/Jce98s7peGWS4v4x8XrYIaKkHr0Dmi
RUeLvecM8xnUGNqv5K8IJKUUSkgbSOmwBWy26Y2m174YQiyWTSxm6yIX/wk4YJtV
las7oAyFXYTKWQocl0U7D+z/1ufdXHa4m39nZy2jM0aXlkFA6fE7jZ2meSTRlbjT
CD7FJs7lg1KLDitRqqWIABXa27kiUuOhX3Lg5oMhqYJm8YDYkE56ZwSo7H9AeU9E
2J2HHXsYLBAdYhYl5WjRaXP642R+irnNGZFAuJ73j6KAZ5JuquF43NCdHcN8xAcq
jUlYpwL9MwPJlZZn177NXUFg42BnhfnvElDwxyT1qVJOOi4wga6HBH6ieyn7U+oI
0PLRCSnCqxLlrOe33NIU1Nqh+EgKkwQnfQ+2HsqSQoWdPISi9+pStfN153kTa753
L05sGtMg8E2Gziw79p5IpCp+NxMYiqVPRr1ZRZzH6ja83YAPjDY33qkoGJe1XfSH
YUOAK9gb1Xz9s91nzQ1LwWsr8bYxepursLC5bKcMtDK07yZtmqHAgYDKODV1UnkI
n38Ce5cgSdrbRNaKGwEzYH8XveABo+5Pj7OpG+bIXio5MTwbW5ADC3sNfDGYgAbf
DZ2AZGtICeRpilh/Uf5p6sbVWLc8kdl4zg2WaAt/GPvkuIQMq5awx5t0YFxPkEa5
gFjXOYi5w42jbmFRVd08m9hl0sVsiET/U2EK3MSVwZiNf0zCdj+sbrNatAeTK4gs
2toJ/aeRWDYyBkkA9alqIFSF9vmHQ2sDoi6bu/1KOWhOXv2R0W07lE2bnmnhegTh
pVMjntI2yiyoInWqsHNtq8o+ubJMu3/ZtfH/ldE5uyHCJtbg72iqIPdwrSUwqAvK
xjyBlXc+/oi+KGqL/pKOT/T87sH/YXECjh9x8+2wXAqG4kO0kRpy3OEn59AbkALB
L7NI4gK3M/+3D5JgeIa1vKcGIltfF+Vl6+WdMJRLgJaY6fHcNyYR0fpRBdGSLCHB
hoCp+K0fQnk1ecp5Wb/Dv+rq1MebNu3Z11P8pcisrMMZQNiUGdABKbnbGZMJS2ML
gkgSlrhZ/O4GiIQRSvAXiIO43Op69sbUqsUkscMlehTrrKgUcLk9sCqPuVFO1aGz
aUXX7JjGES2bGfBOfm0upSgB/+xmGnZv6un+6Z6Y9Y6re6ZyyV4na9wRrTGK53+t
UVKX2e4etBWBtvcqOIf5AB5Nij0WGetU3HlvFJuuQegOah9/qg3AbQfWkxaNqfnv
TYDFUNqvCNu8Wm3waJRPNUYn2ajNbUfVXOl0ERc1Qyjin6Sx7k4KFGEY5E6ShizE
WrkFE4TGuaHolxsY93weaQuBhrOT14THsSj6hskmxTxcapp8C9G/PwRMdEStj5rH
Fys8ubPvHjfcldtk4FqWIU7SCZLyzTVCaH/3bvrvLdoxJNZxTGf+jukWELX4Z6BK
NRgxWDW9lgWbtjgvIzYbAHJO4HLRIHR6xpPZapKUCX5UFl4BLDrqMNbbKzii0ABc
KK/L5cZVoHVBvW3BY5SxAp+RaFwkzzIZYFwGr1dwHHgbe+mcxy3t+d4thP71OEfp
lyheb48VSkoDImzHsN76f4Iih7L6nT5gCfjLLIkrDroEAiZCR6CEu4YjSq/pr+eg
qGuXThqydkwAKOEDtrWbuDPtuRLGigcrXTc7p4xxZ8MK2mzJkZ57A9VF5PkXndXP
3yQKLBqWM5FRCbiWjsmO1aKF9oC7wnSBR0owuH5vpU5BtPXdmCgFDcwNgvIOB2ig
Cbrmn6J/BcUjrcSYDybu6L9jcuUR9mAEjOLhzqCn+VyBuGXhgww8ahw1133a6kFC
ozvtmMY89xR6cHPJvRc11L88CMCuC3/cBUXJIMw/XX9hO13JWTsvS01h1SOxrD8/
nmm+GvNOR4i+11hF8JnU6mbHykhlnqlGrpdwNkdpkS+wqMReSuG3CAPVv9cAPRTz
h5aIOZNhd6/RGuqeJOFM864bxC5GTy8ghww0amDOyLohHpypDscPIY6DzTznftE6
90R4Jqt7B9Uat1SUsUyt3SLxzN6IXI85/WxbaqG92gKNwODcKbP4y7jQ8d3Nn/un
LJ00NbWREg5Zlsd32WyUUZqXpd/2hPJmhgCCXmwNX/1znLbBewu+XuCSZUIFGMuR
KlsZ+6EeNFmJ68IMkdBQOQXt+7KVP7Sw+EGgfSyfz6p94HOyf2uUtzD1KmOB4mjX
GjfkWbLUGtYL3CypLEHwMo/IHYY4Adff5eETWI8WUJZV6KyOlG7KDQyeLBhVnUDf
6+bZJnXdbYnfFPiNab2gCyzl8H6tCz2Mup/8JwmpFBP5DPajDSOloRHNlWfjUgnf
cO0YVyoBnYXE4qaYbBiGuSMHkKEu+sk5uij78tgLXxx4I018Pc+pYMfE2RzRAVch
EPvllhgEkbTnxhIEsXu41gJ0fFmXYhRfX1znMB4f6+mjKY1Zd+6+lu1dMx6LQs4D
tcVJemAL27BILb4Oyv50W6pkoEjfFV4spfB2rpu+2+Hl2YtP462yoh5E4xFPlLbk
Jaz2P4/TPyadVs+oNppqjes++FcUDOt5OpWn/HKPc4qr2a/YwdghoGeiwmYa6K/M
tzaUSqvmkkZ3X+H3TaIZoG/lskszt+KXqe7XX1ZIteCJZ1scqXfHLRKA6nVbZ/Z7
1vjGZMcg8nqe5YA454Dt8576bxOwNl+UOfc3hS614qrH+2JuJ05ouPf+8P6ZQDzi
g6dd15LD7ESZFuG8LnRfsMDhHJeGP9XaJrnL/3ISKOGiClSR3d61L3O+s3QuaAeM
YZTYA0GDvPwkRUa75LOHvbGq6Sjk07N9nIzVybadcoSY6JIReObwTh84PguZ5MbO
Y23kKjMqM6cadGA0njDJ2lT2OdU81bWnIWA8UEYvEDUUdzVIFgGwzfo1WfATmsEd
sEh/cwhDBYm4xVNhUQQ8iKwyZLbyz4+aC9m/r2zShzNdotgcmbQUdotQBiNO3ezX
16hhOLBV4OeFY+mRkXH070DP5PZdCF6Zbs/4Ovy6NoivZlwwUtTYiT8JrRvCnjJl
W+HmJp8g78xE3+QRP8CjsS72XHvp/C0iqc9Uuf8Uj7yhHnkNQv09GjRCP8HpQwG4
lfUOknqq3XhGBxbuoDaR5EYiEpq7hzfsKtDXUTStmlXeL1Ie1z0dlo0IXHhfauKi
+gSrEAd4hDpwNNZTlRUR2PYBm8vATJ33RLWOww7bXvgZEWK580nFeJLM5P40FY7e
ghPnnT9AzgVm75KpAf/tmnLX8oMo2+1F4FcuGIxVc9Nl48RUXLvQpTzgPKH5+IUa
jZo9K6MFcbeECRq9jDHs+xGI0clp+vi8V00WcWzeLd4t2HMk2yzm7IMk+n9MCyJX
rBeHNKNOVvp0f6so7qIezg07jjOmgn5mKYqRLoqGYksxsDLozgEcNzURpb2HsCcF
WWZKkRA4s9Rq0KKTjzL0btoTs4u/83ZLI8lw+YBPOBccMpbD91Odc9TWp9rh6FZ0
9MEZKwAqKlEuIOytkY2hK2Q4NzZ3WAJ5BLItyx1h+YasPld1VbNtFZf2hD7pfBJW
5Qi3JUj+teAyf50ogn5feooIlpxLcXoFN8OSvlYKV1yBNGAhD1r23JOG6qsasluy
vlCxR09GRu595djJuvNyAb60xmD5xKPmw9iu5MKClXHPsb0MCln8VvufQ8BYurhV
xh+muwFCDnlSUHoRT0FFRPpjBnQ6ltfvjHp1rXNjLn1Hd80IUAZXwtH/qw9vdvqi
GXhXqV+LCk9rYliuu6OTSHQfEUOLBStWi/855SfJxQnC/tUC7dFMKCNmleEDrdkt
JIu/wlGYDBRLa4sG4PeVxAkACXNvhGnp9NrX966gI0+t2MWd/TiDQT8qKLR5gszU
fvYBwcw2EgmPQl4D9eeas05eLkKTLpSEKq6GTQcCuyHWyjd0pb9sNORjjE4VBXMM
g8FCU+F5cvL1NgFn/C630PaASBPBGkH7phJW16ps2cmXVln/5MtFkYOjJd2jkOUS
2bY2fColWu2HuiVxzF0OC9+bDqQhMFgsyYwf6MMx7GB3tKoJRnpybiLWymvIAJU+
hCpKMJTItBECi3g4KnqyxtAGhAaIBO8XkR3ofTr1sbexyW+qb8DRgt4YsSgLegha
nfmBLZcEVx1jRjDcGgNimX59CkfVV9JcHRKXdUDfM0yx+DeUNuvQURTLASVdJg3n
vrX3qd9jGxxqGLAX4w5tKq2AqyYei4IEFbkfKUC8hVCAfizSdtttzqCJJh7+ND+J
svPb+oUHP8M9LjzbJbW+wB1CsOMNQ4ZXdK+6CplNI5j5PYcCr96v29T3ToSKg83b
sUspMl0yK6anb11QyxnE/OGr1Z21IJtQFPUuoS1RZtxZcAO3Kh4kFeq6VWK9n9ns
/OCOY1IDVJv1Iuy7rkF5aI4c/8F0cm4nFm/qwFNuTqPXPkrj4paUAZub+jSVzXuX
G6y9od1mDXAZwhBHHBFcv8Zza94715q1PEO+wVy7F7OrVqMydzYL+z+xDLRUMKcb
iBi1KwoLLpCnfntUpLt+e3EjQG1k1dhV5x6AkLu9cteySWupR6sy+2r48I/YHspl
yNOL2N3mzi6OqSDXBfIAWo4Si4r8XxGTUs3uqApNNa33yfuxibHDTyzyqgikg1sp
dB8EbjbbTtgrUn47crZGVfXhO6GoVixfwm+TUTQAQVxNxS41VXoG2IS+PRb6cHrK
iOJPp+xYl4O9Kk2KoaFuxvFXZlF+ZLWrIiWuuPOibyC4CV98orYcgja8NFrEzYRy
Rog3TrLYTw2iGFmgMObXLwR4IMbtRgZZIKlG5z0pbwTFMT3Lng6cEOnkRvoiiuJn
ij2845LHeF5+M90Ybsv3uCaQmp4y8s48O7kF/1QHU/t5a+kxYjs3bne8dvEUULOs
En1dsCVyfFY0n6UV7HYYwsVaaq0yTjfq9LKzJikaD9SehUvZdJSwhDn8WV9m6kpU
UP/vQz6v+al94XpVEIBz2TgQbntwS1gJyrqgtpqfgdIezfF7WzbpzadAbq4OMnCV
Jg0phoqwA6ZT1mbzTpkw623yNJZ1gRWdHUVk4SXH8sb/jRVij94kSRsBJ2+jPQ/g
4hptNbIl0kjgiUMj/Wvd5JluLdRjFE4flZsh6kAo47h/aeg0a/RSDC+rSKD1PskL
4iK1kglDQ7HfnOOQ0I8OZJiliZlekI/WrwxjnUmJWAkVloHt2mq6Rppv9Q6q4LK4
VMaFAEm0WbVivtCkUKwNLUd9HtR/gPMKcnvjhiPmotUJEvTdMmp0WYPtQI/5lB/t
M1jQnmBvN2ejw05RaWw/hSMdMVfaMsJNIM7onhyaZppEzeTCaecf+atRd5XynnZQ
m6e7Y2C/ReGhhTgWGX63S0bgrOcovYY6qoPeQvQWvNCdauTTkYVV9rV/4qpOsel7
iZzWbCB/fanqsvksQsJEQdax+tlqo90eHkNsl/+s3W3KBu5fX1BcUpORy9Jp4IfQ
HtmjK96kGXvXz3tCPQZWSCC8mnADvqaRXXI3gBpPGYNLu3fs9o8jB0TN7cd5yq9O
7nLVsx8lgrxR1uUPa19VN7w9BijtgsaiUnHpFNQYIIOh6wa12naso8VtS02FKA7D
Wd3AuHUDqUaa6ZtTq42l3IahO+wxTztVC3FjF04EcJXn61QC7wWpcCveZWO1r5uF
w0aKAjf/n287VKQZTG8yX0p/tA8Uy51auBEQDRTUf5F5YUSAvnvnW+7WH+OIp3Pl
8iurGgGA727IhmVUrqit/IGQ5R9LCy0813iRUwVbHwc8UqQqsj3Awq6j9ge8vYtE
PnUOlbXCA7RowRMJX8Irn9KReqNDbQL2LPfAcy7IvuTP+AvjyfCyewqX6MAIUW2c
4jNJ8bJASAcmSKxZtyOX3YkoR3OxxLukFXCWyI8Xfo5HSuZsmyaYPeVNvLTT3Qbw
BuenHj27ouI/oRurLqsH6GB22hLwLSompsLU0OXuy8SFKtJGR6CrWQjfGE1QWNan
/SIoWGGS/NVT+IOCdnz98WtN9vDMXYvE+hKEjtegZe0Ex24WkmJ2uAMzy7ggEzZ7
wVtA2A1Zkew3K4z+0d8eMnupekXSpAmYw4ezpvoGxS2iGCxIDm9AF+i13kgaggSO
Z3Q6TZemGnI4hqZ/DBXRZHgdy/8WbY1l87cfVArUF35UIuwRkZf+KfbBCsA8S08r
AHcLDhDtSz/jM1V1PpljIozgggr0oBcGUIlj4JGvXF3N6IGm7tjcQO3uBWvD3r5e
IVS9ezq+pk0Aqz2/Py7HMschpr8pRNAh2Nie8z35sJ1lsP6p6CcJSTzMIITBrnOH
1Heyug1kv1fbFz9bSqXa209sMpxbiS2aod7HIyiCwm9m08NCxNkoxH4AOAid3sS1
GQ8cS5zdkwW5Trbb8NytivWTDKeLA0bgILSOV9lPu7Lt4RZfRvoTph4Bj51Y+gAM
Kdt4L2/ObKp6buVISBo7daAVkoWyvr3jyFeVhj4YeLEE9jJ5kyCt4QfZ92z1tcjP
O2pPfpv2FaTNwpdyMGHjUrQDQSsuhs7pMy88II39Q+z5mImmZypGasjMKVRS//zz
zMzbScve5BNRWGJIsgXZPydyHoHbuL/XMNP9CUHPt4Z3SD8r75ypVdWE6i8yA06n
Z10Vtc1GWRMaap4gEQmWz9wPiNh/VMnz/Or9lkmFtTUxnHX7QUjHm3w07+koBTg0
eIGb4fJYWfH5lENkcG1AErshm4hJE1aMqd95dUqcWWcGLsIV2TbejJGXRxgUEf6y
r0xJZ5QgJmBk9JM7+ZqiNwMUZ3HCr60UMjnahSo7NSNLFSoXZGSpP+4vHlTG42E7
r+f6kTEDNPugvNxpO2Tk9XGto+dj+6+Bw2aF5zbrqvp3XHez/QzPm/1j+qy8qANr
7COGg5lOfC3BO5Pcd/pUw8QB5pkMJKxqs0DBGdc4gY8wouRsD4MuI0s7f8gv6xRr
LJF2fePHErHOWK9PH8Mphc/Zc/nBdNn0rjhpCrOnJ4SNLPe84LV6RwggGwC5YJpy
MeHJnomiYD6slut0alDm7/MF3Ec1NtG9s8Kix9ELVpDVxaaBEme0VWhNTz0hiqob
/rBsl7hCJAbMi1EoliQatxKeTgypaB7SwSGrZZBcXSBvJDfZn38x9bmE6pJd4kNX
yLQBeMk1fHLitHQ/VS7ml8sbxOMbSQLGr7S4ymbMBHVZWnvF6SLuo1a7eMNO9ABm
bwJ+9hGXOo4BEe+NfY+xL/GEY9NrpI+Zq9tI/itPkMPKVAthMdBN+eJX5syEiwnI
3JckArszc/BPuFQhpGw3JI0auLPPnoAweE/l1sKNjG7GryLqTO8r/xE7U0bF3fqq
TAbY4x+ucZ0Zk6rVVnV1dhj2ABoclrZ9h+SasxVqaSDJOWtDB0JFBb/1HMtSD5Pi
t5nx/LsjfOhrqA0GDBdGctDRqS3XgrRn5THFpp8AWsLjJPBTyZrV/1iItHNyCvan
9zf+TJ3hNEJbBSok3x0Hyp9HukdhOrbIERdNGMtm8HHSEA9NYF1TONTaz6G4qKlx
mxpGhBpE0FzKyg78QMrgP30jGBv+ht3QPxCIH9xQEjDo/Uq5rF8XnMGiVb+yK1m7
pWDNXSUkgpMSDMU+2tcdlP7aHQ42rTz8yjSpGIQLHnG3TUOQs89mt+O5xCeaex9v
b/R39ByqEwguycY1Vuz8eXVqGMZbbISFcSDWKbayMdILW93roC781O6VgME+epdN
bNGg+TJrqNUvVvZy1su92bJnPOooDd6HLcJ4REgvj9A6OVPf1zvWpHwWKKu5CL1M
yr/sHjOLcR2DCRZsgUMk4k6wEMA+hk0ZdWYI6VzpwWfATuj0C3WGIQN8Pbp1iCk1
tXWp5Yu9N7jxxHsFfDwmtB8vNUNZGL7jtSQ32TfmKsHflo9WrpX/phO7BPOpQ7DH
/H3p1uHsJayk1OePTUw490bOzaJ/1Bv1bl8hB2Qk29YJp2SIlBkTLq07lNS/70Iq
MriDgL9z2MLKl1jX9r+Ft9iityvM7+ADcitrVtAqE7SnzUecP6ZQMAtWWbUY8LvQ
Y+P1r2q58uv7Gzew+ndvguOppqg3Y6wja006G2lnufUzD4oc6DUpLRd5Mf4+jRRv
2cL3bOmBiOcuF6G9KfaWSD3mwrD8scJCJveWr2OuuIdKzMal3yFksdhVPh59h+wB
w8oJWUlY6HOvRC1IcE4XH/WRkiqo0GBcmm62U9xX4ojauu8ttatJkPDRqsFrR9zR
K/uwVvec6MKVR3e8ZW+u/cAcKUD8h8P/i9UEoFa8BanKWyCJuqcdswgRLuwaxeTn
Tf5CPBmWhQSYOJzjcXfHUYPwbvj0jKt6Jm35Y9HeFv3uL1e1fQ7xLqruC1GbsltY
g3ajcrSuBi2tZkzplD9/GEtQGOL1fZnJY86WdmVuIilqbUhgVIdHEhBOmxOTA0uF
KIT7ChILdtFjAO3a1kzj99DluPwCbkMZHVGrWKYn3SdJCqkXE7GafQIL/qn0Dbko
kCLtcv2rAlPtVsmua6RcpM3ev5r99Ma5s96iHJCXTeQg2hTBrAtNVF16k/5BHrz5
qyH9sG/9Vc5X2rGw/tdihHayWsurhMj74so0x9j3gW6gYNkighqY3gNiR9WcdJqm
Dgwo2QRFsDZJjol8dKxzrMJ/QuQmlKamWvwSGOj7A5nIsjTq0ACX/K7xlGvXW+jx
L0y7nP9QqdPWS3ngNbHuX2u8OJP0gD/80mLKgHxZnos6VLvgF4rBoXuk4JUWxe84
nrBx3sijOIDvPjwEOQ5Gy7DSHaAzXCgXPR1XZJ8MOGt5rfgX9LpmYwfewYRb6vYp
DsMSFfTn0VG2IMz1GiqZ3B4ZK3T55C25Z82stbhKDWW0fI58EUqmwMh1OqfShXZz
TuKdbDXQ3z8dw7JX/DHXAWLwCcqsjntVLdhxCARHZRZGPOPpW0My6QKEiod4SKGf
6FovDBCDlKsaKiNj6ihskszyBLq/gic2BP64eu07hc8GWXTRjxa8iQ6F2FDldYXe
/7QasH/PEYap19K+AF+ak2bWczgqtyrK3MfZ1ucPECBYr3yOnu4zc3qfie4QKKRN
S2CwKAZtBmiCXPA65i89vJZshx0ugTgn4xoSxggUUFJfyjymUTEPzjrz7KJUAdan
xxzKHlQIq0ldXLE+UCPi48uUFyxBbhm97waY2L9hY2e+bImQKYDQRqK+oTDM8Z0v
WV2gsMkaBSWkPMRRQMwFH4v39rxkLfFXJWe9hA/xlnwUi7BDFKi8ZHW+ohORKGfb
GAsHVWD9wZ2ebaVCo/irtGr+Y7utbCghECA8eDfhCCj7becK6atSR7ka07HkDv5V
AldScp7bvL5TVXzrmocc5ySeIyPptUfYFtI2MUIu7+zZmm4WBg7nk0NpkL8HFhXb
ZBzo/dhQkdN+GO7eACX55MrD4AgA47UZSXxxqe+iBCKdxrNmoJYVIQxwOHNNsZyj
QMgBwQB1GePsuYWg/u3k0+GqBFzki7M9YUeD57q/vsz4Uq3DES6m5zOD7VzKV6jj
AzgM8WmRqsI+dNUN+JHHb7R0DxFoGr8J/AShtv/wcHbjTuSZxglIfNQKksqstq6D
3X0DVoSwVJtNYGDa6y8/sChrcQf+pWj/HFUSN7D89fo3vNamQR4RXTdcrFCojQtL
PflcRXFDfcDRjEx7AWbgraFKiwADfOrj5/yEDlREnBwIMTAAepmjTlF8SuXeCmku
wfPhkEHfsKZrY4VjUmMjGo6XOztbpgjid/E4Djnc9+mL3yCOHgtTKo9bs1PgQpDZ
bvFpwKVDnmEkJtxf/eTb+vkfqnAz5jDK2wuZ1GHXM7Y4AAPoJHFSfXyrY+JuBobv
jCNWGsUQkhAkBlj1AVz7bPZkZC6njOSVshmAQOfozK6DkPXoCeez0LLQaUTYWDaN
lTyN2SuH7Vw5hvgSCBokHSGHLm5sQaRt+AdGibcVkgKLDrQ+sLofVe7IK/AzcdMN
B6gQKGAtEU27GxdkRvqbPSBTQKEUoU74Sy0zv1pp7qiHn84q1CUVEiWYCoesdyI5
N4W8KKaGMovxLMAJmixsiazXb1MyqhVTsXX9AP/zWWnWqd0Lf2WIos2vTViehYg/
J4K3AGqFj8rx+CQur3WK6y8cuSM9XmepxSZEF6iSotHw4SdPN7PdBV46/Q5ksCs+
LoY3kVb8X25zVeOM+WpTtxmvYVOw2ktBZ+YHWo+mcV/i6DkwWj6Dwo7GdL8YfGvD
erAJCq63xSAihrR1tSU8GXpm+Oim1Te8lBMubsFOrdOJsaH9yI0CdrDu+WqQUOZM
ckuKaxP+lDcWPZQnZAruL+1Mjj59jbkwvckDfzacYO6uQpP/8TFn3LVxIDvo/Q21
OUDb5NtlCW5eP6yNZa0bGsZlWCE9SjiD3hJcONkBzemRbyUBFeejWK0umx6kBMQ3
KnT60PJEsw3RHhk9MHToE2MaksZyO+DHbV711pZ5XCwPxyfab0/LgRspSXICx0H2
OcFy0UYB/sLo8iAzZzH8qLaVsG1N2CdrVOKX3inIf0NKgGN0nYNBo8pFZuQzRqR8
TLpLB4/tuHwnijmJrRPQbiqg+2qfqhrw9IP+5YRlGZ8aBayBqfe16mrM2EOwaVhJ
OLFZLgxZtAe7ADyo8cM06CfgMqHAgGtrSkq2dz5s4cPQdDrPqR2QVt/is1OYMoYi
N2rR1UV0Ir1Hm9HtIc2zDlZtqZ5b1945BVvv0+o4DDQfcGG72I+kN+oHjwISJLVU
m1ip1fCxw71dZ0fmD9PxrDyrVE6NRv9soXgwNxoCE/4CFTgEoFbPRLYnxvFD6yJz
NicXMSf2TTG908DXhfyKoOJTebZDii4GUvCCawKhYR7sot7dX6pKa0+f3NjfMg6Z
igAbp1GjWJuHOF/ECOP8k6GYHs6A+kpjQbunfSYmQiQcfJMdZnlraY69tq2bwlJ9
v9NzLT79F2Fe9swCxww5CDNAZcrUD530SsMNvGYOrVVVlmFPhpzFoKISg/IrYfUS
1I2UfFPQKztsWzEyM4bZteM6M3I7h++aUKGUqTdv2KyfGqkoFjqEJSolIrnQAMCX
XNEHtj/ruyqrkvAiZBg7UPwbhsVLHlSHWZ0tMAkcgShV9gOG3Eo7/WzZrzYvXtpm
4eyw7FutKtotOGI/yFTiTm4yuJM5cLcL8H0MvHukzAgTxfE29Ua3j3X8K4Vl20+z
RvxfMY9QX2TzsvpToak+DKLoTTBTDDhBVwNgalsZjYA2WmDjevt5KzBCBQEvdDLU
CoAb+6AFfiLPmGkFquMglH5+elFJJlnwjmtlf1/JMrJ2SoLabrYzjVCKg7/xpIvO
Q9TLHRG5CBmPulAHxDOZTQUShsy1pjv5NcSS7D5CP6nFjFjvIOOuILq2Bg1JnfLl
4VVCtwJq+Gn3DZOpzsqhhu4op7XBjp09jBAhO8YSqFVkJJSzG6sBZW9ydyyrEZzP
OtQOwudtwc1JKbF6Xe0K1a9bTLZdTuJCsRxoeqZRTF1oLEGxWdfmq0VBqAMRbFbq
K1n/0pdb3ukVJd9zHBKytJ14MJ/amuUVNeGPJEcF5klNsaYcWsS5m4kg/2Ryjt8A
dvZEO7g8sBgE4VVPIJK0R10n7HVHr+WSSssFNIQc4EoVMqYEbpH8cHQyUwKdGlLm
qovdUqYNx3enRxZR29eqrhJ1IPmwBq9c/eLlpGeIADnIejF9rem5ZFMOK8hsXrML
0NVp7WGxjC+QM5jVef58P9n0RL4BnfshLvpEXOKwQnBk6MZnyZt1T3BcT32yxDhi
R3nKLDjwWtKR4nNI4ajeq1uVU2SDozFnN607HFZQIKkHAJ+CNTUUolPbwt2FhTqM
shGHtZx4ieFaCRHJm43TLSCpuMUHLefzjxNn7T5mWwa1S/SgJoloKzaip5pLd5xX
Sg8zBRm2MGzFw7sotRrGHLn/8NEh1jvl3U2F9u7Y+yxmafW4loki8CXNW2hDXEuJ
O3xUOyVeOfFnh61bBGITlNYC5128GgtiqGpj5M8iluUxQo6kzrqocPhkJA0zBxw1
NMG034Rz2+faRZ1RhU+0uRAs3nhe39Pnb0SVfek/q90O5f3v6d3upbi/ZYwmLx19
9FzOFat7xOYekqusz3uI07WGD8Yqz/t8fJ7z1E+V2pfWASMQiBEBSslY5FTeDrsV
9rpXmukzZ9J+jaHGZkjg9Iqv3e18FvkW43KJfhA/yQI/HdMWi2VYb4bYij4XBbhw
ugjnW1GVMCo84OnPi/fzk7ZW9XbTp43D0qUWlfEwO6mfXLfD89LJK0JpT21QIRcl
1hj2GXwFVOA4w7eu0IUPnmGz9ysWi77lTf4ZRJnmDuyNRN/UgzY4O0UZG07mPUvu
z0xKVzqId102NRyn7tJzMzO8TSxJhnDHPBj9Y10Q5A2oIS73SuuMV/RGo9C89gLD
P61a+7YVrWexA3NvDG1abyKenefNRk/LvVXnPOj0externX2xxOBWaYYTaLcSLWw
hYw6JztD1VTg2l0RjzE+//Jbe2ujPk5crplYmGPytNux6dwTvJIWiyou8+FwT4rn
0HL27MuP7swEvUOvXkR+OqjY+Ro6sVF+ArAP9o+q7kKTfmQbfYs2LRH2QgJFmme1
dJhv1nsWDtcbgvyGrJe50t8EJrHToJ+3yIOdwiMp7qv9F31kxzwtd7UIzOCus2Z3
Q1nxYyM98VgX7RILMJ8PJu0QiU1pLxwtnNLzF4kFFeG6DYwQROU/kC8HYVS9O9J7
IetsFwzb3k1SubXd30HbA7xmfQTZDUeMaXKjj0L9Z/sxk+K2agr6bxE8y60T6HBQ
7/qy/T6hHeCZbEXyJMpO2u3/c/C0hAYx5AvedLOkQeqSkE5GGauUk9b8L7mCCiUs
fhLi7v2gE22k3vxgZwBuCAxy0Wn06pjo7TKCEbvKZ70zIsGZaOdiNj1bP9CMwR59
lhGlhGvWLeL2IV4E+G6eKnzMR9rPeYWaKWyXnY9+oBJE9mH6dlUiykO0l6mprjMs
I1SlAD8Hh9P7Sv44NdX2wOApvZM51yyGwetn1YgFs/D/Tja1QnY4FY2Te6f7RQOR
VeAPzJCwZEJNIdkpavF4owm0W/xll4d6EkvuoQS3Q1bSZUhCEx92EEEB5/UXvyTH
l+uMB0NNMAr8UI6R/bN4Nv5FGZIoxoxMusmLJk2vUPsgC83xZAlStqE/CJh8P/Vo
7iOJxDhmVZX4fh9vJD8X1xshhaSjJDTG7HH5HvDG2DYz5XnEdPta1zEF2Q8yLHih
2YCkOJsUlqR3W2HYdWVrwpXrws1zPWEfq+z0SZNEgBm+7KZoZJTtp4NWI0dwo81p
f9VH18VRQv3atz7K4fjK00mMCYbX0GMh0791kEwj2NtuDUuEGY8hkCGuVg/ftg78
P01P6KPNNfwMapc9E91H8XoB0XetzfGV9Afny4sHeH5OSbiiuYkdG840ymPytV7W
BqvqKgoQD8tfERiKCImCTi3n4tUqsXNAyTxkpa1xqdERxrCYVDSDDPSwWGc7NSEX
uyTbnqLwuFSNR98NYyPjExmfWmvQtv91Sy+YBnTX4OFPVKmrwNeess9JJKzMDoSq
uPSqpXb5UzVFGx4MfT8VFrX/+cgcNOueIgcGA5l0roS7uVmPYXoaEu9zB7LPrlHl
BUWtRKPk09zkZ41Um3iDOv/k1PsREVX1DU7GQfrC9aHQ13SJzrg/rAPknRFd5tT/
0M8sGXXHLwKMahoeMfhsVfntlOGHSVhmqzPcsZgIy/qL0zW3sKV89iWWqasuV4Hc
l2N81bfbEblkMQCd+b1oTyp2pihvLoQnzp8tiF0BPDJ+jpTjqzHfSVEFdKOmiqU5
adKIzljb8qslxiXPgEapkm3Dt5ln+yJaa2MiggP0vifPAgG/J04axPhl+FRt6O49
lR9UCRInwRzEImt0/aXYddk+Q7YpTfRRgv69tvfRBgWzdM4YWjLjCiLGQ9rPkk0L
cRRXS8B4S2osu18MOKtq54JxpSiRVsy2J7IsLvXFzo34b5wmJQAsD9RJYqDeSzMR
RIDc8xwyMVn0YnYvhwq+Denbyu7Q4CKX9OVWPcjRXs14rNA2nPIOwYdMFl8j3qyK
eAa/Itn5YsvsAbZltSker7zPSg27CVl0unjwtraI/McgoJT9uIOPQo9UeEBOnjSy
rf/pCRIcdo4j4nWYhEu45ShdiQ2GJm/0Bc0LuTExFdRRjDVkG0F9GFxYaWLSbO6K
/8yGC87JglKYCOcGbzQyCFaW9izv82uzKezVzmosV5gnNf+wu1b7zIVg8kqKcPGL
tua1g+wGa+Eo08VKy1yhf/OFXTdMEDwfMhjJHy2orvwHDA1JM5KnYz+Jh2bbs1wY
vwhecvZ0LnhSqGFBDGDm7LKda5TZT1nNvQLZwBeGDHTGBz4lh/KDrd9kvUjhPWcI
ltBBGLFqzCcvoqsC6ZTJPQ8o67fQJ+wqtd66OE0WWKOfHHqVDJwUdk20G61o4343
phTWajFpKqJMBelC8N1Hl4DVdenUxBBtVZRmyTENdfJtCfOnO2RHf4ytoPDa8Coi
ADz12vA0A/3o1ABwW9oGr5iobC5aSlK+PAkvJh6cddiI7HOkxLwR/hfH3gEA3K/d
9NoPUotX1P82niDa275LquKAGAigB7XLQlB+HWxGVtpCRsRAeXgaawZQMAv5aFC7
tSuVzTGfUDqVpWRGC3NfVLXuxjy89B65LaQBswd5YA8+zwrHeDcB1x0q+QLSPdcl
OOFybY9LbUwY7bvy4MQBxn4GBXnQ4Px8IgCh5tD2wFAqFdLJmtAmiA8j7ONcoFPi
22lfpOWCps7RjbWr+7LEAM9Zs1838bChWrIbfYnHdW9bM/Xci/OrjmpxHYRgLVmv
kN0d581pcAt+IFvpIsgaiKNubjPFVYo5FNmkczf4VZB7MJNB415for8na4aYP/kw
Fwarpow4dv5RKwvKU/sgvmGfnZu9hRgKe9F1qi8fHbhpi12Xkps05CxncEZp3OmJ
+yaoFHy1kv7YYDp19j8KFTAucgPlz8ZXiXRlT6wsILKu7PGETQeG3pW2u7D9nMGs
K26LpA+HQL1/sp75N+soIhJpNsFXz8uN+pGaBv8axm88OFVt89w3LPW2TJSzj+Vv
DPp5hscEnUaZ8XydZGRPcT3N7AK1Ju+duw7VcjJFSmj7QrDvNQKlz7f1xUngC+sN
Y67Q18pp6TIyHfZpBwrO2Y98iGAIKRyqH4UbvkvGkOaFuJyjjpI89qT8W/9OW7Rk
xJDRWyjhywVMCLDPJUTDwWMxPYdWoQXB0Rhx2SlyHtePb+6taxbo7/+XNM2Wu6wc
4gdmbKogU95va2YLFzMS56cLJ150cpjhuNCmN/QQCU+cl4fhS3o9kPguhpQ4yXx6
ZGZZ9iRbsgBz+rjMKefNQNPau4xDu+HE4HxunyzW+PtbxvZ27I0OGp/LH+Kbh6Iu
hRIJLrXbk5Qe7/7jw6NfwGafkPbLLlzDzlgdiPsSmviEm6ewVJ1P5/PJI+GR7nbq
ddBZk4dTZFIMFtn/Msm4et4JlpSbM31u1ZTQLKlgCKy2xgwulFvaLt1Y9KT6igGe
dNyqq5LRPQSAKqPmtRpFvmfu1vW9/1OoNlMp5SPPEAs+NTWbJWx2+eTESoMJhO57
nbMdVWIVz1sfb93lKpX0zLUJFuOLTzMAK98pWKa8PFS3Mvg2YJkqPuCwrion8dfm
y/W1P69Pwne82fGewfNiokV/NuY6Gtvkv2VcZFgIYV1mzR7N4gxJjUFYv8duabB1
dBcU2GU7FCrvzy5xXvpyqWAQgiAn8atcui9AAfSaXBEFjv8t7nPROgIRGEbwB9//
kglQKxyqZVWoizL9veineWGYdX5o4LckXBYkK8OYhcQB+wd1wWjUI0Lix237TLg/
CCP4nbHL8JyOn3lxG6vFOKiebyunVaFcKAaZ9rUJ/tcOcXuBgyy+A7dlLgf7vAaw
5NGS3U7BpsCFYLTuRUVzQ1VWXPX+2IqxnuvGkGTuBJzM3blqAs7zzp2B8m+dUTuZ
NbYLxBdjeFBk3DIeZnwkVRo3pkQc/kcKHI37I8QePVb6PnyNkBSl0k6Qgs1GnRmE
wy7q3sME+v5I0+WWV91LdZZhysp/fmF2RHa8Z7a/50cL6avSri8F7Xe2GfNaN2H6
vY56OfYOHdnXquYgk6WTHdjtRYug6PvMxT9SKVNMdn8VyV2SS8vOKfaHKlWGmLX3
SJj64FsC8kaq6t+6CLS6ofXOm3SkZAwNdhZwdYbmDNVp7d2F+SfUK1xd2JobRuzw
Ik1ERAL229+GO0jmSs4GQMFjnd1yLUmRQ0ucQRFRNjSWjrJSOrpf9THZM0HWctMn
HW1wJVmXgQUgOtVq9hNqKhf8f9n+PZUbdWcCp/+XLX339vhbnvwFhuY96aBrcm+P
aEzYoampy+NAsqNpOkar2eAJ+IiKEEg4iGcUhlOhNA650n66RR+6HPGG1e0dN79S
568piUkPltRYGiSkqChpW5+CES0nHDMwCnSJxw+ZGh9MhacneHmD8Vw14ToCUU6d
ytvK/y00MP8NGyLIAd/mVJaJ6yYj9cuTqHdqZjvdfdhzSxiVWUQV6PDGVhs4/vzD
5gqzzZ36gGJesTqH39cGrjEotvr7bMvcf9jmsrqJZ9ssOPaTZC0f2HCJtWeVvEHq
bma19XATFohle2JnhB8+hoiB1MIEb7MTE4TzIbTcu8d9wyIJi69IsuOqeD/lgC9k
eFFfY0JNEf7+LO3G+6B4WEp+TnrYEv0qggITAQCC/+73TYL5j93ucrSM15NAXEVG
fAnMmyb43N5KfLl6y/UBGdnyWh1PiKwSfIwzcl9vhJ1nMR7khsVgQcn5/nxAvHw5
dp4Fxu2iZ8wZ5mpIePEWl0eJDrlpk5yYt1RI3X+6JuoLsgxbnFQXkUzY6ZIbrIya
BF94spxfNmZ4/oBU4P4/ZHI0GFpzK56sdKEB5fUpDe8KsvXUFY55n6H/9KFUpdqR
hOBEMeojx2agR0RHOp8JFvMwjN5JiQtVsU2OttRGlgckbKtpY00Z0n+WZ55LZweQ
QDJ5TLezQhisDhNbBGLHz2b68PMHXe6HqhVDYZ8LO5CruaYPPpJv2/d1Js336VKk
evM7+5GzcxmnyweswxNqPJmVXXyn6fn0r3BAOHu+DfTU7PLAMZk65I7WBtjIjFPO
ewqKrGLTn+m35nXvUTRAaorcp/mx6Xsln/fHFMmB662OyIseKuvDm6yfwPhMCUH3
5tKDL3l3i/AnZ3GgJMHQJmx3i36wtVnxemp45h1iZWiTFrKyzHMf6E2+ybhxhMFw
DUNHC8eCPSxxR39WCP9vMM6Yes5XhR1AmuoDAb9HWbC3nrXxKkYrbb54G0iFMOS4
CXazz2JiMaDJOyXbCQj9Ew35mHKC9BNlL+jkpebw4+TeHn9ZOYwfHXqwjYK4deZF
pzstMjI1Lygk3hxvfx/4aPlcuWmfyzu1Lju48KuoWva6xId3ptO7Uig62eSQq3RR
0hzEevJoeipMqATKyQWz3l5dPCef28ASV754zSwUXUzUOMJMh/hxxbSUtAxFhyvJ
pCZ2ZSMzAdVwwOdiZgKGPnD+BLL5dAZvweSMYAdM2d2rBhJa6KGuJqLysC1gSS6E
32OCPAHjiReHIEqoV9Vc9YOKZG5tvgZ+e1t2s6kX2OkA4ZSm2kB8WjqD7JyHGb6u
QmgPk19M0Tpv5gScI3sOqkZnLAXyE2p8ysRuXqeWNOj7pGqIhiGSoNM3hZokbDWJ
qiEEyYoMquIAABe/pFcPK5w0K6/ckNv2dGTqvBheN2J9YQnwYYN2K8wQC/bYlQca
Fa+uLQggLpB76lMK1UfzPOvOky8/cnbEtWk1/z6BjezbpqiXiHtYZewSiIBXYRyg
YRBwzD1ppfrBda3BbgQ/taqWzYX3s094iXOw9Wcol/8xZJpHq6nKXIU5J1lWmlUM
LhtR47yLMfBp9jERlNCxNr+QwGKlIWNqXE/03bCjdz9ACuTdfgiN4OAul284+eAZ
OHe15dEzw7FQZKj+A3Od83TYESQIq9Twbrwazxmim+icHgmCoRF3G2X/bE2/gpy4
ARlVvYlOCsxg6XMcBnPumLqRiI0dhf3tHmz+BXWEFVQ53rliJelU1ZDpj9BKGA8D
tA4M2EYo4Yce2lBlWGeq+92JhRf6ICEjq1wtNvsXvdghLW3sOIWLnUqgAAYk7Pk/
J/KVbF0Kh0GtZdkZw1e2NcwWxHbxAOE2ZhZA/ZSFde7h2B5Qkat9JSmwM2BjlI6Z
+SIwjSv2pmVQ4OyX9xreMuhPyPQvwVmHh7fT3IPPsixPI3rf7/a2mbHpT9WUqG8O
Kz6x47mbs0CLaGC4YhDsY7qFDT2cWFogWNArhPOAlgjnvmujEoaxn1d9Il88yybF
0M9sgdXvRaQzc55LCLOnswU2X+PAKaFjCTWKAMWBe6t7czX5uYxnvJniEsl+WDeP
uyNR25Ct8RZqithBR0OpxMVhX8XfAzq+w3OBlqhCln3+Ssm2LlmZksFZ/kZyU+qc
Yt8sRr2CuF88LNvVqhCCB0DsNIWgyCWQVubKubfnWiDEnsOIGkqSr5+fgPXCT9fa
cb3Qx+cruFNfLO3FNn9ZEQ59QEaa4DUvvUljj1CJ0h97p8lW9FA9KXBod8EEb8Ua
rQrYVFSZNLmYVawJBXFHBjpokTI+7yW+7+h+XSl7Cwf7yTYDlmBAlT75e/NhKfEq
9Fpb4meXDduGqzolf5aoC/UUKYzK37QR33RY780ciFcjF1xCMhZreyvKi2dftCc3
3cyao3ls3C5jvp2Fm/JvNiyTLJNLNC32298EXySvLJnrIXOnVFbXE364+NPaeK9U
XObT2Ea84FZo+OL3/F2yeQkkBOJigcsCE17uNCMyDFbpbk76vrn3pxXrAKcqLqC4
WCYwxFsPbo2d+HzTq2Ww7XaY4KGShIlsXnXxM7vLtw9awYsnA1Rgv5tiVXbH9Cbd
DN89fRQ22+NG7cjswNoONj4SMNp0cGeAnIfiumav3ZiE7fGtSYdizVCLeF3aT9Bb
4K1zneTd4TWQokclgnzxivm0VYxVOef8IcnIurUbgnjCe74tQXiPHp9r4gUqLgV6
iGPXua6U+Os4xRri2Trwyx03nFLENP2wLWfAaVddVD9dTPxzdCt/KWwPwtUlYoNJ
ysAOPuf339hzTMhkycMAcxwW/AR2yydZJZ2TKeR5vr/F2V4oarWrkgVJ3BUXJ3Wh
p6Qo0i/ruCe7tWvAR0ztG6nSAfSiXHvdTKCAMGFEGhUAzRmmN87N/5bil1LXKaik
qg2S9lCH3AaOxiOGv4x5UsSFtY4bLS2P3NMbyADzJzrBtpejOUFBDQcvMNjZu3wA
wOtjZWcX/Zmzk5wHEe058QqsxXEtpBr8V1jVKSx9JzbNde1nTp07yqDfEpqX5I0v
GcPQjGzMf1BGXu21QLQeJXHVnosddhC/0LaiGTa1RF3G+vlZxM4dLEdjvq3Qo8GB
iJ/bEZo4h/qtdWVVGIRVmSrI7iSOqFC4O6DoSw+rfHh7+x891tvEj7NNXag+jRNz
yCSj+GYXYpb2Tbvcvwoj0wVlDyALPJnu5iSCAPOhGLc4UzfuQ571+rHJlppWyxRu
mDwYVsxW6csB3u+ihszUq5xFdEd1qhZU7I5n3y957kA4wwzWhDW6b/AyjYyfoJmJ
YPyEULWXBMdhkUhiUlM3nEiA5CIZouy7yttxloojKtPwMAW3zn8DnqGY+20xExY2
eJZBpny3Wru5Ch5toTB6HopQiJnKakwwBt5NDIHPOgRNUgjRMixG6Q8b7cmxGGmI
FFKVlz0e3nZL6MvsAjsEY1uM+PuV6uwRqD9+ttwaa1+7gHW/sBTBMBK7OrwyKHAd
wOqEtUmMcKJRlNGs3KYXl0lXovxOgPW+oiO+vg90snCgZkrlvbuWW+2QybrjKkYa
VT4huh+J/6/xypqsv5I+PSI7nFm3tuOCH8wpbioMe1OIS1Wf405H7k1x1GyhqAp2
cXXvBekdAxcFdqHFVsCVEclOk6rFiMn8/9ZxSN3ja53mUIxeXA1dL9P/yokI1l8X
IFDKqrjOVH9pXWuXJ026S+Q1MsBQDocHaZJVFDpsFcxeC21Jf5BRbtKcBWjC34Um
/Tse7k9jvEDMeGQB7QZad+FWIN0gZfsQym8daiF7MPsdxO2Wit0NGZKkC3CqlJ3v
nc4mnxyiOF4EOTdMFv2Oo//DOJ1FG5yhzgeDdqgpahl9AmsNgoWOL/whx3n7lJcF
Oroj/rxRpHtvKodxqu7D2IV5zInjPFGpVnSPSMMRA/BRjZj5lLJrJcXcNm54/PoV
jtaWkMkjCaoqFs+ROsSQ3n3smDPmLSToHFRETyXACvdPHbHdvV0aekf+ztezYv6X
itjPsCy6WbLCsgBt7lvPHuI2CoONQPIuOjfEk+BtWgRchXkqoAk1v91JdrLo8G/x
2y07zS2bkL3QONuGFtOfdxmB2hv29Zd+LzfXc/0X23/OgEEnWaa9UM1eTaP+7/Zy
K4cZjYxdInJz3FDIHuPIAlZTHd7E86ByH4Sr/V3TPls/ReRymf76n/2gQ35vbwvo
zTufRfCTwfTNfI0oUM1hJSoXBCJX2mgBc014Fkzv484Y5QP2UMPMNhNVJ64dU2nv
Wzi5YooBKK045+xQuFmMeSP+tveOy6q2JzBuuMgXALiwd9mEr8nMo/f2mH5TtfXK
VBND+Fs1irGlQpZRNtDI0vZao1RLLXE/Ny/FI7R1sHf4VWk0ngeChM4gnm1Q3d4E
XgUov3Df9Ox/kKCMatLmmliyrTaIJDsSdFCL4s1r4PKGA7btDHALdyHyYiV1cnBX
mXVBKIjpxyegLFmzX00xDsHpkW4Jdm25X9jFBj9x5udLmcU3tl58ofMWHAcDu3bh
1iqHCXouiKAzHDE3QhvKyx71hNfffY8pmRWnuqcJO0Lx/KnICZk9oRVKOJW4y1yl
2SSZGW9MCnzI5E1swzJU/Ct81IJXa+Mmd4KODMZ2unLFtRYAgwJqT/lheOadIB5x
3R1BNcPiwSKyQoSsybyhVlJwlj+ZBb55+lIAaMmkY5uSFGVT/tLGYEpdegG3ELt6
2WocYeiXQtSAmOhgzYjpYC6WuSZgt/MXdt53Qz31Ia42qA3Z05Rpj5SA24PDmLTU
BuetB+haxucKeYGBnvs/50Xp9Zok4CHbOu7kmTxjzyX/IWijeG6R3ArTRpamWwoC
aGBGbI8kZOZuTbjBagUwQekboTkFLovmtXMQAPD8haHBiJbc232iv8QlrLfQ3Ab1
QBiE1B3PuMHAqqNIS1kvEDqVvTBqMdgmXdTXKTFxcv+Q4K1za5Ruxw2mU4OSl+im
2G66rHp/tEcM8BrNV7Ikid3g+xTRBkSVZTPonu6og+LS76LCth1hHmcNtaMT5VdM
cUGsHZHeFmCfAPCF+CfApMDrtdSmbRQCZ3aW2VKOKvTN5VTi5MaVNT92Ke0av+VG
GFD1rzWBeoVrk39+cdExrm9aP4afGXbzM1PKMxqVROqZ00wkYVFrvrs+KAr6s8Xh
LXS/DRLSFQrrqjXuo1KUEm7xIEFpfAqVOF0EVJY8PMzPz0vszHkTMbrL5tjI+Oe6
M4UutV+FhWXRBFcFUFB3bnCaTqQjNzJMxXxqkf3psgfAFXVUnGNOs/FmQ950XsFd
aWMUf+sKXiArnh46CgVZuZ7vNQQ6fTy+Dr5i7dQasV4AbBWMebSQYDE3ngt5vEPO
n9taZdFhEH8DhN+LEFGmZjRLpjKXmdh5Gl75+Yi3pMBuzfVCkqgv1gK+TTfT+IyN
OJFuUPCEHspleUBTvQLs7CnXYhwum76xrN9ckz1ocOE6Poq3W6QJcGXl8Mo5RRYZ
0hiDTx5SMpfuGP+kGfvsVmnkVTtGPPBXiv6aIdmgrCVub1I6btu6PzowTfgLIBF6
maC89QVoB6IloL4kN2kw6v/e/Klra8asibW+80rQ2VpAiRLLqcVo5nPws99jBnz3
kQM04OSHPTr5dHCl/KHgkc35t+FlTkiWqJ9v0PUeJsxD+AL2iVKlYsw9cpRZcmWi
ATbSBcBoklekHX+r5k/UvR9v0sevBmsN4GWxXv/6agWtFL/6ss5FtL/n2pWqGFoh
fR+OIEvL+yhz2PYZazS/FfLYSUSnWA6fwKT31UJlL7WB1sR6y1fXEujB8K4TU/f/
o1jML83CwcXt67jpj25Iiwz3D2V4ZRo+gXuFOAIlyl5EExBvbN7tlRKTEx5FnYpq
r4cp+EewoK7lCuL1MrWRMZqUBZpQaX8iCBZ40bcpd3BfzcR9pLLS6QI1hpBMMY+r
1ty8leHrpGSfCEd7+9C4Yvre48wjOmO6JUggz0OuBQFBzfG6gvLef6CJpeXQLENh
YTJNHgxqUzv+sK1fNzAxWv5SiiNWhK/2IRk9kyPpmBEBIzc1g3LkC04KwLptW8Wr
IGJhG0oN0P15Uqmg1lv2DAht+QL91YZUdsnRwkNvh8QhrudHtKq32XVb6DXN5Egp
kBtmBEDL4TqUft8T2Wf7oPz8NXH4cOZ++0hhnq6K4af1o8P4O1agSSPvFQaewU1y
0yoTeGYgUWmCEtJIAhyKLCCYYqgbLFKzNrTimmiLsdY8Eg6ZBz1RjqqY8X+uhZgm
PGgStCzG8guE7ASAh+NPxKa/DxT8q03e346y6ETmAa1VAiw1pD3i2f/8SWx4Oq2G
ctANgSqH5vbdWMv6ypjDTrQS85VMwtbUrpdaBO0T6B2Dmg/CYn7sXNti+RCO9VZW
8XLecaBhvDBO1fRTgGuzv9AEzDMJS6vSExQttg0ukiSNd3n+EcYjL6srFPhqNc1X
v12seYAApORdWwUJsxOQSR3jHOPQK58RstpNOM9VYAYTZA+36aevm4mbAVQ3V7WW
JknZWQ1s1ov1jieX8GiwArxkTy99iVwOY7ly6kF/Oa069MLp/e9+BBrzILojcOxO
0W5+8BdmuZBZmzY/ywXk6cT/GD0U4IRr6EgZlW32ARUcKaB6/X6i7WodigIWYAUx
Du4OqFdB689MXlIUBKP3KlgGttUM6HA9+GRc5kAUzjlPX3j2AYmeUPkNCpjS74TX
vDDCyaXqV0v4Sev9+LHtsg5HlnbhsbtU4yRXCtBBrb7orukVcpZACcXhwxdr2caB
tojqhPfN7WAEYrLP8jDmLwlkK7gDSW4v10tjCbZct1cEVRM/IZBbuYZfE8Jx+328
oERicBgBDb36vd2EIpjp3mfPHgvtGwgy3j0uYlRVfClrpLin6p4+MBi+f8cVby/F
t+k9mtvUXpPu6/uIvaxpIhOypYQXAIVUC43Yj6lP78NLoJ/UArHZmNolWWMGeL62
oDaETqZXiSNYeCqceFDW1j8LXtBj0/OTWi+3YysUrn4UDmo7ar9tsR4SUoasNcic
490ksXcypN9KZTh3Y9x9BtVgjK8lkXDq5i8Mars89P7JXkNB73ikIc3sLOm6wNg6
48gmnJ9ms+NjFyX6Js58Vm94FgOlbg9m6YM9+fbnHOaYYByVrm+wH5JejgpiSmSG
ZYRxOC5VoXS0px5dB9HMU5aIMQmjy/wiiS1gUZhiEr9l725m4ViFJRF44OnVSo3h
nk2dvX/01/k4WiZ/yYvI0fvqOgs7NlQ2MTxSFyhyLj1ea+2BIhCbSAe9wwcUENRi
4dVAU/JumhKn1mEPg8eQsoVFm65WG6jtf+2xehcDxTLZMrIatVcKI+p/PpKVo6qo
2J/xMXI0eSxS/mVYy3XqJPyIX7eNtrk4rNXdtBsE/LAKEY7du6xeowDOHQgpwvR3
MWFuadsBE2iINsJ9m66N4kR6gdN0fcpPk1sIih5xhiFjuNTL/or7c4Uvejd2S9Ob
1nSJYDKbvMWFDpIsnvBP3AMEGxx6NGNIgROnbfBGGKUqHb7eV5QMpaK/msASzy28
rX21aoxfa/TNJyXDXSLg2JH4Hs8twRENny4zxUKQmE3WDiUgX0Y/Rdi3GKEhBtET
KnB8+mb7vW24PQOtXpt3KbOgDIu+pzN1VCtuANJbPpJj/y8HijEl+wJxxaejxQom
jH4lA68Bun03WTBkltnUF3tQbkM0S3jsuk+nzAmd77GC1FxzslF47WFPM5gaXXI8
ntKIcH2n3ZTRlabjbHbyTQ8K5uBMlkHRW5sqAbWcxefi2hfLS53z3bD+Jd+9UYh4
YbPP781wDS3dtbe9BBfGY+TvgTmnlsiHw6vnrxaYa6tCu/13WHB7jd5O53NFt67f
/qULmOxbpqyhVlUknmDE9r7Di0a4eb7rY/M0eUSe0q/ECkc3hFaU/61M2WSO7WgJ
7EZN+uvBhsdb7KGjRLOJcnr3gnVWVStyDYdySIhOs1+PFLR64e7av4CnT+WQ2Pzl
SerRtA47NkImMCo0YTJwInXJjRmkCRZsIvp+gQx2qUL2WC/VYEBPlAq2abHGoAwp
rM2LF5EwYwPWtoEureYUQyYPVZNnH78JJryewPrhR1BVP732e6GKywdMMgvteKDC
U9gBbKBTCgBXA/Y+tgb8YqIGx4G9qa19iO7pYNWpeHOfwVqqBe7lnKnubl/K/uxU
TBRHr1G+vPMvJkJdF/UOa5FPc1V+kPR1QZJ1X76VA9P22gp5QwR5iKh7sacW8bO/
ySGHgLKjDBoWiqubol7UiclqbE56JDnFrvR1TN0Tml/YpgQQnT0eqVAl+/rV1r5x
rYmiraUJsWaaPT5hgcSRbp9ZQqL7N6GmPeDTJxhaPF8zYlqVpQHHtqz4elumkCWc
a1dwV5F/axmz3M0wy+CQUEKvcabnNzJj7QPYNNvlEttZD0It5WaWUflThSOSvOBu
jhg+Ak8EIGxWvTZ80AWtCR6QgVBbrMGgI+GXtRiZPjkQ3/jIyH/oeHR1j/gOMs2z
cLCum2TAfxFnjQ6m5CeAjq8x6gf0NuPBJ6DN0p6pU3BkarKMkCq0kIISipvNrCJs
e/UZlYib2tOdwKG2EQEJCcFdQfOp7VsEw4P59+GVMbREwvLkeaXjBlikuy+sAU01
5KXFkyd6mdalcQQJX0F44//SHFCltXqSdUC5uGDHvkvmTEQ2YPcJVFuyEn7c+BEn
zYQ6TQhUJQH/bjR6kmhqJJ5Nh+yk88RkPkt5PljGpA7TFEYAkwzbRD7eEd8kiSJZ
DvuXq8QqaTPYXu/K++bGkTOJCALB4BYLVl+RPBcu9B+8MYQgGfyB3H94diSp0xne
8fPFFdAbNTtHtDtcXSFlW1Pd42j2UQl8WrY+OTfb2KgeipvB9068Rr+1LQfd5TYa
yT42Z8ry97ziay9SWOjlYYcuMhSdFcKHj4p6ZJvs7cs5OgE15gXkQsG0cxWXNuT7
RtfCx9EgL6fp5gcnnfZd9tLfvM1S/t/qlUdD2W9ZT9Mnzbre8WJS03CQzrmjen4f
H2FRZLLDShZdNHH3M6sHBu60YdRtCIt4JNyQWdS+5arMXoq5Fepp1SLAfd8kyPFa
oMAe5L+9Vyst4lqkzvEaWSvMnA2FvebuP+Qkk/0XWprGDfmGSdFPbBYeCEUG8dNa
WGT0CYt1jLNTWJmyQqmWeOPrn6NWXs+qMEh0CaGFGVllQ6Q7ijrcplWAQYJim/hv
2duNkY+6LCgwYIszGCrBVZalgps8ngsi+bx8mjDqVppmb1pl9LO7wb0heG5jEF1Y
UTxxtIy6JDMWgHR42Us+jdEtMGvOHO48uKMgtCvtOHW0i1R8HhGDG5V5bmZ8ngYx
DH+ovtxQTkIjdcQcEcabNgQ2xlIPgHrmS6XdG8/8WbdMV8wAMNZQTmOAN78ym9o4
H4brGkGZE/aFlo52MboyEvX4wCt4eV8Djo7zcDBkh7wzlJ2YFQ0IiNdJpczURZvX
QcGHcvlfzcwrM+6Up06Q7V3QO7owhngzhFGQgaxD0V7RknQPlbRhaaMPakgk9R01
qx90fqqvvON7dNrDa/rSeJi+Ew5CgHdIO0nem/JBzGLvsUfOlEgrbNoTXUa6OpM8
z+HO9g6zqviXQzo8rtsdgdJy8kAk8h8ubqCd+5JYppWN2m3BMDO/2WAr1U+zBW5i
2DainMG2yIG9K/Nxg/34xFI7IGMpXNpk8OTf2bzgZwlTkBw+QYPn3ccQIfxwBwTZ
HGBuzA2cyzzWJfz4WRnO+q/DNq/OSJJIeGUSmpFv8qmidODxUU9eUuMYj5ibzQaa
Wx9d0xPwQqDINpDFWGhI6lhsxeJWigas0AQP3QMJcdLvz5+ENL3l7sL5LHNtXWNU
ITG2dQVPr29xWuemYDYVnZ2lQJZlglK1DcUJqrs/szoX30/oa7Yf56qSoWPf3n5b
rUr58RpRbuRFz21MVzt0cpZV80clfu+Wks+d3iPFhQ0rkNY/8XWMRBHg4BON7hng
leQlKgt2k/xRjfe0DK9NYER9P6poH36N/NdUu4sZf6AvcrLGpoZJOqsBEeJa4esb
0lvRRktQ4YJtselikV3l3Po5r/0Ie4zYlvi9loLmgzu5ey9KCpJwaY/BUhG2xyFm
haFBar0qKKcNFi5SMhkXPkvyO2/qvhsg8zm5dys0m1M0cWqmzP99md21Q/xM+AHA
gcRb3n/fhFFKsRX5xowwTHCtuFcl5EaOPESqZvQnBs+u5pzaU2bpYZK1NQ7GAwjP
IfqlzwwwbTBbBjFYJ2PkdZkoVXH61RLVbUBRYqLdyIWzP5f+KxU1tFc+eLRnKGXN
3HwhOO4XVCJP475VceOMSzwveWK1YabeHrFJsQ8bz72HYSBfZ7seMhLt9amx8noF
Kps2UCs/fW965vwZsU2IaQTfCc3YAAjG0Gm4Vd5dcib7gHIs2myWJ7GpwJk0OA3/
fefzp5FniByKrodGkYkaLMw2RnT/aRAZyvc/jZx2jgmVqRLsVPOhGyC3b6sbg/OH
w1YQAttxfsR/JhH6GhCtwBtBmcQBI5sdZCTjHgehma/FqGXa2Gwi+zq8BsyW1gpD
h/fjRaIQaZFXOFzz/iZP3M5SmACKwYZW4CHlJh1t5olCiajqliG9GxjmGmU4gW3O
saijFjoYjRLy1EqaGEnkQpMl5eZDUIhY+Hvz+iQ0j5cP1P2yOgiJGBktD+vafx7j
Zn9hwMlquy4xLEzbque5iDFGjjtDOif2ySwgld1w7lxERV+1g7oc8oUCd5a3iSkl
Pt3nQIRs5EH92G9FchWVJwkrRmHGskD0NkXyVFT5pBNyDULuJHs/phOAKxPzH8NV
LuU792fsBMxlWCPP1rYAkcvUXkxE7Gj3GwtgZbdrOGvhnCN+Z6GzeA6p+PdZP5FD
YCWmOwyP1El06xqiR/xvNmF+0lq9nm5y2FBtcB7rQPzxLAsMCm6wCU2Tjy8p57lZ
q/et9zEth0X3S3DuhmMVnvT00EeWrasnC7NXmjXGFd2eL5T1kQuFiqW4hHhTBPEn
rDOxBqHvpImIZmsO7FqENiDkzv8dzMJA4rWh/ZyLmXKiSn8aX/R7NULgN9b62dI4
Z0RT8NLL4TnIv8OwRyG3v8cWXotLmkeQLDNhJ0ctSTJBbQZwCLPNRDiDxSmcHHyQ
K/4RlxoOTGPtJv2RtrhZtdCk+76vksZeptnP5PafGeIPtr1wpafcRhXLF2ZXGfgV
fhK9FTS1PDmeKSWc1RfcmXYEGwyrxUO4puODNKJjTdAk7kTgb7UpySugZE3feHnn
l0dUvWG0bR0BjFm46qYJDPjE9ZauqEPSsoVEztSZefy5bKA9cZ/iG6nrJUcJ8Kcg
bIMet6nu5wbKxmi6VS9KBHDq1Uk8fC34kHjmdHhsMpeTNGtLai1YHM2/TrA5342V
JlCa9FMWrq+ApFSc98mg/xotlnrxy5Le9qopgxQWBpaIP8wcRu4sWt7NOXX+DmyM
7xSBVplSc2F96+HQwvuTOk5BotcjxMDSqKj7EI+e8KC3PsH1tE4ixylfIe7gouaZ
ZoTYReUToQmKKHJmasqaPLM2W/o9quR98kv9gyIQE4QSgIC6SYhd4A+YNwC7mYFo
nMj6HjlcZbWZGkNazUkg5Yif9ahmGzUyxPDge5ES5YG02rC4VpsFUIn3vGPWXgRY
`protect END_PROTECTED
