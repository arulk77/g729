`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
1tUxEaOYoBsPKnQ3pQ4TRJxpgxwvi1DLa1+QXT6ymj6br2KUy3mjXLNQ81Z1Z/lI
qXE7Tdi+AxUpmqVkKYP/WPEbyelK39H3kh8n+Uc9ZkXdbIy2jN1Atktuz327m9fC
SGzaEQF8OeRG5Yf/GFYwLglQnnKe6Y1sn6XqWWegPWW5cw6VJFhcS0NiAFQIgDeU
1SglXyGkXutvuzOK6+NOOistdZeF8I7I7bBfdNNTwmVvTOhPyfkGGbnXTBowUaZ5
3dWuIzMhU2durkNFEBoPdI71UwW/owTJ/WdxRHyw9g9flPBq0oaily5lx1Vl+139
pzQHvPt0qePENhITd0D4YTcf5LRWM4EOwDOAdCamqSyx4oRiws/5rGanvXHBHcgS
VDjaX+LV8TJ4ZyLiItzg+0pDZlfO1JwPRMSpF/2khg0Xyi2vln8+AdQqYXB5r1Ec
brGfqc2sFR0rETMgRTruYqumdcg09F9cqCLV7g4iJl9tA+cbzYgC+k55SphsTyAS
qfpdy3QLqt9EAM8tCCd8fnKsAB+ti0IFZQLsEZ62F6xgQ8SO4Mev8xlkAKsi39Xw
q76/HvamC1qrTNTfRhw+N0rFyZCpuHL82ItsNIAZwDvxrz/vtiQkzjUe0971esvU
4oSHoYhNROwNBuaY+gwgSuQ5SZQX0E7Dm1YTPWxbJMFLrMEXNaP6a0r6Qtnd9aNj
Hln5+EhrU1rAJxge9vQ2ECdkB6kqQ07aCVLrmIbRQITMwpJfOmNADDkl15ToE/t/
J0ogD++18sUS9PkBm/EZfOG+teus45S3GplcQe1lZusZNYcfx48Ca0F6UGzimIVd
`protect END_PROTECTED
