`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
TnEungXPrmQecSOmy2JWw2mGMULvNMDUdgLVjGzWSuWPG+Y+huY5us5gXHdbaaUm
Ka12l1ZpMEYbuLJYTYfpy2tL+vsyAHNc/huWBxJ4i4qiFFjdmQgjWlU3AYsh2vmN
ubjNgVist3BFFlvNjaAi+w15iLvGBlWAKCbIDLSUvgj9WDm4frtlIbpDsIGXefD8
VVmcwAu7G8MLypG2QZ2IhnsyKXU0J3wZqO5HuYwzCpTsL+33mJK+gE+QlrXsPUaM
4eGg/IM8MnKa6Lg26rGxH8t8PjKlwnV9KEr8PrNOMiPbiC2ItjzNQ+X3PgRPw8hW
s1gaaIcRdcdnqtARFgtPUz04Bn9MitGXSlR3YNfb72Rdeyx1A9LWwSskoWHj0az4
iqoBOK8ZRBMZ8KU4nNrVAQ==
`protect END_PROTECTED
