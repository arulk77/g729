`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2RtTiaLwZbJSuPbraFO4do1HumV01pLYjPcNJNVOSTElmqvqniLuqSUx2hThJFpx
tWeD5WrCEpVh4GIzQE/tGUf1/hM7yzqPTB34ld2UFnFAMCjN+ue04BvC6lLIQ3X+
S5dXiqX/MfDJDtL+9BFKNnFWX2A0HBWMdRjrwuv3S+wCoaHEQY55wn6i6qncMyFE
`protect END_PROTECTED
