`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C03a8BLS4JkxP9BCBvoUJMu+gnuX0meWLwAWYlVOIco8
kyWPVCi8m6vM80nqbSkO9pcUSDwUroWbdWqjTKzf9KVb5vIkkiRB+MN5ccfd/IDq
EMVDYXozxCe1BxJVDjYt0aQpB9gXAAyy1O+I7tcf+n60F99zGXNCqxs714C54Sjd
Lt3g01rVDZahzh5E3Ed0Ato5j/08ASjvquaP6Hy4dE8tSHjUl+EhOmpbseKrpVnC
ojt/bJH/tMBiVqJzzcLZQVjyxdyEDzqcbO7ZOvHjhZFwn3Sn8gCUpep2kKpU1bxq
H13dtxIM59eLQ87lhbPG4ROAQbErBs8tNeaCcNNO6ZrKGXNWkqWkzYwKxpFlRzDs
8g4PyLpGvsgl+LKnaxHJhSZJ3+WJuSPyXhL7yPjjyLQi882QQ5F2C8fjKIw8EKpm
QCeKYb9oT22ARC8tjdAOJwN+X3I+ko45uQQJeqntelN8F4QLjfR4qt8i+ZuXQ2rA
XlQ0QoZ4JW0u0pZABEpndzH7kvwpRmgT4aC8VtAyFt/6qUnh8628VVecfmghAX+m
72rs8PyqAc9VPJfzsbZ0BgZqXW1BTREdZP0c3vyjPl+GpIcEO7FDG/JSPsM6hkNR
cVLO+7yZyuEsY+RpHTmal/A6cpEp19tsVp+x36A0X4uBTnZJpQiGr36X6j603KSc
w42o77vA/se0s0RruTxTbAYhNUzkd/GmVry+SIC4JSRFL2cXEdTvA+Ka5woS71TC
kW8Tvr+0D0S6vhtBNxkSWuTiUFno0cAEVLmRklmW8m5UuzODCGwL93e+AYJrDDfE
PBlOa/MI9f/Pf4bQTxrngi7kG34sHSYLcTmDTSqKQokPjqvYs+aiiTelGzFSyBKq
PWyF8Vyqw1o1FWo8tWPLmfl8QyWW3PFFx8rJvilK1QG1xq6LTa26Z9qVBxeAwWec
P1tWCaABjJIbsWIO6tSrOqKsQRA6mhFBzijXX/PfpH+5sJfcLHKW+Z0C77dzzmtF
Fml5ToLGnx7BKOgFh4wGG7WyCLwy9LXqvpS/n2m96mh68Zq2C22o6y/bdQZev/82
2msyQPvHA7EFURzxtanrBUBHacUpZKPcRbTcqF9Rmb9tt+ihhwR1ch7+oouKQDok
k31kwMThQW5lMIlFyuWycdCkLBCmgP5om42RTTSYRNe8gYUoo/zXZAtNCU1RD0AQ
dbVNOIeP2+6wKdHZJ4sy0epj8LcOrJ2ievEN/4nPco8LUwigJOFwj7oaZRF4mFkE
kpjIluQu98o+s2sXlMClHbl3TF/UuwsOh4A4Ey4NJoU15HUGr66W9TLbRe0f8yqy
xs63TkW9SGfAkpYHGwcbTQc1or/scXO6ubPHb/Yag2z+4lvViLRnji+lUeJOORPI
mD1TIjYTO0nc99KQNpJIns/Os22A0iK9KBMISHhEcZy4UT5Ss3HNC6YDHXn8pcKV
q5RAL5qb8oOb8WNwrEQKC8SzOgaEIBbHUW7+pBgpKyb3pueOA1VydWNTDHhAWEFq
Cmf/ySYtlejiNVjaDIqJEQnOGnvgBELoSAfHGaKV/NpSvhY6fflDOJQ0CKZpf3CG
0AxsH9Sqf3Jwz3OI7shgHuXBz4G1PkgqvTzvBhUPXbbAb/2pwKBqrpgSruEGN0LU
/FqSOgUXtHLqJ9avaolR/+SQ1NJeAAz2IoKKOr6H1MkoYKZr3aSfVkJrP2hCRLp/
L8gSVTukXUA1XxBz9BpB0yMTXoQBbDTtWw735NjvmBP2XdiXtmIFgXKlMHCeB3nE
j0cWD2VoqmwvmZ7QmcHqnQRx9TjahkevWY8cLZunJ6FcrGh+dttHSaPEQrwSFiZn
EBDYl5pn/Ra2IBxD3PvzoMFeKUaJGMw2hr3qjKuy6Wz3e8Bqrq1KJevIFn7YruCj
l2sFzi3s/AucuebeuiKAyOD2JLQ22sXkZJcCfyNV5OyN1byTrXl2LoJDO+A8CT7m
f0twUeyqZmE4J/hXpOVlGoNOBI4ysCs1np4DZe5hzUpFXeifEDOrdz6YSiT/ZxLF
jzUNl+FojK6VrxMwHI4lKSpQ5nXCCt+Hrgt9/zsb8tmRyaR+7jfrcya+E5+Q3ND8
SyAyeNkyWl4vJQXQ6e/hL7vYEWEo3ZIeFvFeKKI+ZTnu1LGjqrew3m5CIxaiN2pG
16I1GqXy76IT6tqXnsdy1DSlmPD8TSasH2ERFuLLw8bvSaDGmLYGPywy9g9sKrZA
ddh+KV8KbwKEHk9hWOyR6McAPGFLDN+ghCYFrKGadSuLlrqgmcs55AwEuY/TdnzV
9YEkTOq2TSCAU9xA2xCo429GIWP2oc28RF0mvGExVSF74sXKwG6KZUJHMUtHnB0x
8n7lckUXwIm75wyVuTesGFp4dS1mRQRgXUxLTrnj1PUzTUOSAzh/1xMsUaX6KnCP
V630uCcOmBa2sDubQ3eh1joR+jWWS/7X7WHcbEIc+124WjPUq0w0gkse51yoJHdf
Zjk81gxAqXqhqnF39D29BQ==
`protect END_PROTECTED
