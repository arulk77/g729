`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD33gSwB1mt7sb3nvFAG9SNW14RCGH5dz/ewo3kOPfOP
44Q2bUxqebwMTP74a8i4qZAEav9aYLy2O/yuKiwi0b8CLNah4MiajKRNMy0nqrma
9+Fe8jEbRxmvA+ZeUglFw/lHZrzpcJI/tvvZUmzhvdpo3UjzHuG0GU90hfcNxKwy
1KeAdcg4N0klY/WWxN8Nc5f8VBYxoyxDqlvN4z6xBLI3vcpI3Vl5GQUJwdR+pU4m
`protect END_PROTECTED
