`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JS6Ee/OUguv3S0KjECptSAlt7ujjzjC+yYTmGGInI3CzH+GlNOTLyr9yC2wLTGz+
DZ5VbtOJgzom2b3T3uwHGkz9NZHLkw61iPKGwbx2TiQ97ohbeFEc6xWsa7bN0A7h
dY5AJcrHayb9iKp/lcNZo7irxXtaLvkV73xxw/GLPx9uTvc9MaygldrMIqlBxlod
XA4wH7JYiPyke7Dj0t0oJeSmr7aj6jOS3DsGZrUBgQtDv46rzB/qgShpLIcZjmCI
qMhKlHiSj/HTQM3St2eU24dUW95vdYYw9MpF2hiMxxjQ4TqQE+NJg7zUYdijS5ID
`protect END_PROTECTED
