`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aXGf1FSPRC9yx1w44MglIL9e3DMWzclxS5S10x6KO3jG
C/+EW/2U0N0OadvJ6kpE1c/tQ9hL/X6RSn4CH3qAQHg9F/h+xtafuqPAPz1yLFwG
1daV1+GbiTb1YK9ha+SYy7BwEcQYLUU3HRk5z4F1+hhvzMwzWXDrakdSzmKMZtcU
/t+Airrhf9s2Pu2oSeW6quq1TSUA6WsjKnPU5T/YqgY5GW2XfoY8WeWsPopA1H2D
Awb0ZrLPViF5eFvvHzkwFRdnPtMx62BvH+/PlWrMtqUM5rAW9WTm1yTr6dBx42uq
Khk0tqxmKc5bWlNV04BVxBVqxGclnIgFS00OfkMm3VWxHrVeg80zzM331vAO3fEn
iXITKJmG/zpb6edw6PxSTfmjfMPX2sYq+UnfnSZ1RTBWk/dqlYtu5x8jGiwMBo71
HCMysdSflx1FGbz/COuxnK11g0nmvy9jwSpTUHgncd/WdiZUPZ/mSgC6oN75KYb1
tTMzov3uGBLt2rFZUk43VT1QorDCS2IXclStxArstP5TiVwgpOODqaBYKZaBMWHW
K56HTflMSnwDkus6rgMzulHkqPkAEnyPvsnxref9eX66W0q3LEaq9oauVPcRFYje
Zi2X5h7cPWHJyEGPYB/aldqATedfS787UmVj8Ve7h8o=
`protect END_PROTECTED
