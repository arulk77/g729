`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
RC4bKCQFPX/jRuTsZp6QkSIk+kQD5lIYDYujJ6T8uvzID18lvexpVBH0yBeTBTWB
EcaNkLzk1CH6FoFq60DoxcoBhUDZ6/kbU2u3PcFSN5Ukdjvv1Bp27M3gXS4cRxR2
YQQnWC0jiTWoAvOPkQ47Ujojk3JHb0SdOHqyZeS7vFHcJkTU6p6Nh0NqfsVS5iaN
`protect END_PROTECTED
