`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
76sFkWaWtW2g4TUTKwVVqiwgecb7cOmKzGaZpSFLOn/oI/GPH7mo6l0CpDimaEIu
klS3a/497yJ1LRPkxoeIX2Aum7EjqtYfCFAHLX76DIi4j2wsQ7u4bdvf3LoFhf8P
n7YpiuKTee3VA+asvM4HU30t3Ag1NSqd/F8lCeg55j7K0o6IYOaAVUmbBjSIEehJ
7T1mC4QhKKyDNDmHX1A9In/Z5s8QwpyRV9RIt+jvC1hlSVb+FUpTBc+sByt0wpGf
502iJdmkgEERha2C5AwFVaVXe0mzMRJDvb1Hwulr9iNTgVoRpLVzbmt3x1l3VL4I
WID9Ui8HzBUeI8jGAnEOZ7CCYztP1nKRY2Up3On0YyAHY27z7gu/iJ70YimlEV0g
tfjQFg8E9iAl72DFc2atT2yIhE1+S7NTN868zyHzvISnhoFdAPcT8wCpeyM+TAbt
oVyKF3v/+OiI/IVTK2IcyQe5hazjakQFX7crjnYwyy0=
`protect END_PROTECTED
