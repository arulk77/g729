`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBdFDE1IJd/c3n5WrRodN5U3V4CSuHrTrIQmn//gLbyl
7Q54z4jcHDFTIw6+koRtEqo6gVb7nG11oInQch/dX4SGYRDAS53A8XQ34Ai66BTz
Dzvm5WA2Ikd6YoHMJSbQY2Z2rFKcCCjy3aCx8NKj4vWOuqosxu+8Pvud7Bb8UxFo
jSm6gfPIU6WXWPBjiygOe5NYSqSBRTiIbk57GVFr2sUbnQgLar9haTD/yg4pKsAl
hJeC3m4ogwsO9D2l9235EUaLedOyLsAbmRvpNqi63GG8wx3yj3qtL3ITQaPcbuoi
53CgARCZ97W+d6GrUNK1nfDqZnu955RVoBiKHsMEsgQ=
`protect END_PROTECTED
