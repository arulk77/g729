`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGom8Fqxb1NJYLnLyhcJGIdiOOQbmnfoWDVdqS1DKjhp
VYQau6stUQtTvBtr4mPOew7il8C7Guee+fCoc1dXKxTSQzqKv/6dQs5DRceEnJkh
D+Eyy3g/Gbj+IKjEGebC+p+6vr/CCIf0x9QXgg0crctIcvaVGM16Btqo6rkt3Vh9
yTDunC2N2/8n/aZangK7Nq567YThywMLSOMQUvZPMHSs167uWXs9IGfKQHeyuSbx
`protect END_PROTECTED
