`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ2e2zO3j8D6I4JSYc+Aes9+pBmX5uBUs7fk2bB4gQ+7
yb3uCdg9O5zb2vDjNKi1ndOdFtAjWgyBLj01P5J5X9MYIXAWGctYMr5Wqo0b+/X/
vSKP3cN/ydMI4akj92aTAfCtlAL2YR5MzUJcF1GRz6UwlkoQcBJ8KMg4QtzuE6z0
8BNSEM5IVQ5yOujn/SI9iQ==
`protect END_PROTECTED
