`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFlYNQJoTS5Tn4WXvWSOe5KWNMn34r2K9UCnSaVXRbnO
4rI16XlKm0XVHUXHC5vF+OcAzJpXx33zDXBqpiHEcMhK8B3Su3/0EMvik4h8mbwd
Qrf18qpKDhkyTo1H3RveiiC1Vyip2KNDwRzDW+kzUl33d3t2pi+OO0SnmJPNhSzB
yY+/uG3ONuHXEpCb9AUTMgZrv9eFw0L/WfdWSgZgHwiA/0bodNDn+2SfWE3XFImC
9MeMArFXdmF1FBoNMotYH8Mgpcg4UJa02kSywMarFYg=
`protect END_PROTECTED
