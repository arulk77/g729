`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JS6Ee/OUguv3S0KjECptSLVHKXoZnyw18B0mZvxk/WLDCkEXISKWXw2xwup7cKbg
CCt4U1+hYkf6KdtEJZJ87Zbo+NJwx0DlJdIQqeATn3lUoyBuHo2636UJAZ0F31T9
qj7LYBxNkeNDPBaJUuJe2142z0FY76GjdvuPfSvJcbhF6TnMFj62oDJ+/liG0d+9
y6WY3b9RDnltQ99Wvaxx5IxnO7D1eHa+xkPX7fF5o1oE0I1BZhPUuLyxfplzXz92
uz55wRV04kS9wAjUVinZc8kfJihcVALTLWbBx1BbPIZYP+2t7+NGJDgKo+EltZob
nGlrp0Q4F66j6tBcNXqTorgmXlDgzcZOWlXAadIhPwfSz5trzOW6XDW3CsbOmqUY
0YqOZpJGcLjbPV+yYROP7R76RgTi2PZO82Nx6egE8vk=
`protect END_PROTECTED
