`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44bQAw6LGpi9yfsVuXHgkanGBek1yrMDlY8tWcY9TAPo
0yjp2xQ9VMCOPq9wOSCaXcZsn2XE2MAPeV2srokAluWyFYaSoOMtMdC301VseiwB
YiJqExf1qXGz/08LGkt8/+qJW/ZCzJJgkMqPhT0n3Sr/wLX3vZCgehPkN13VFNJi
n5DlGDzviEpiM/YdJ60Uujnd4cCpw6YKEmwQ3ko2GX5zylKBfnN5nkDnpkpwVJr5
Di8V4KmvzXkUI2rYMmydeQd3yC+/8NjuZScwao4S19lFZUdlw8g3RC5B9UXKjApD
dUBSH3tNId2d+7DIpI0mhXMQV92Hmg+Y0IDShiV9QsSXIgoCHrohNP2rUbvgUCdM
1WNVTiUeoiHJXYsKBGhZWLkYpmP2BVkU2IER6stO4mjaDQgkw3sFrpQFw+XJL3P8
lCSHl01Y47XilYaga2uZp4aOXlKIUeUe+LPxDE/dRKLksIZbm1/rkKGAQMP4jjEF
`protect END_PROTECTED
