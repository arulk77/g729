`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aSRsG4xUxoPG0zES9e6VmOzhjimkfjlLJKf3MPFXG7mgvIbCT3m0j2OTQzjrW1zt
nTpehstoDdd1dBc5nex/qg+C/pO+XqEW1b843HEViMnwGtGYsorYZDbOP+BT6M3f
s1jB2Zjl1jsK6RwqR0hl2ErLjkz8FSIxgjGIGcEaoDa4D8Oy/nqmoGFO9pqxHCQL
1gtizTaPHkOlqrUSSid4+60rolFt+2I5R5YDUqHk7v3Un4u1y5GVdTLXidpXepMq
1wfwm5lfYsfaB+nW4NnRKKrB0q1Nww6RqPqGxtfWdvsrjU+eD5afCaIPljzOpD1J
EyoCSrQWlrJOlN9skOkEZqPObeH/U9Hbh9N9835yh2/HmAt6ivaqBhJyx1YG+kMN
9wWKdeLpMQGVdMluGD13ypoLVcVbn9jk4z6uetDjgZqqG+8TdTPml/TNbscW7tlz
4NgCfTiBO3AyJYsjDWISuLkgBN3pEG2Z0yF4olWFX5Jw+OFhXYy+YP7MsXGDNFIz
oHtsEqDESL4GkLq4eHxfj6kvAE8A6MVyFm8gWqgIdzBJBj21B72Vww3mf4vXLDsg
GdY+1lJ56PkEkiSeoW0XKQ==
`protect END_PROTECTED
