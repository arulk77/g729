`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1afDCb+PoyxSpneMFdiAR2KmyN/N/WHlmGNAwic1AUD/P
MoS0QxUMP4ks8yaU22kgbW+8P3xhzj41G0LMtvwdJln4AstePGb2I/vBi5k+ww56
9pQwLEk90fY/iOyN36/Xc6O581OrY3oWYuyJSR8qMZZmgJreDZy1PakUeWhOX6Rm
4Oj+IHKAHF+a5GxmeI16liggJUI7oguYLak+dR1qEGel+4HsAD5PqX2CX3XI/470
AD1tsR7NVtkJPV3Kg2lHzNwSDW2bykS2Z8ET6BJvCiW15IR31S+/cmenr9lDN1Ts
`protect END_PROTECTED
