`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFGlC1cSPuk4Y+MnugUW4jC6ewlJJKOyRUdYWVYdM98c
P1qz7sUNc7bDYcXpatw+JCdeG3drRV+CBLeknL2SmsojUuNe04rrlGr5EC8NDMVA
/JC0rCGkb5l/XuWdN0mnUsj/CO7TI/bqJFDSm7sYFD1g6yefOi6V+icTHwo8SNs4
KAngcDvKBT/T1sOC5R+p4RaYonkqVPAdC5Y4i8tYRw3M/lbXxwvxo7tR1ZOhL5oX
sD6KzWviJx/xIyxXPznO5g==
`protect END_PROTECTED
