`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHkIuNCahF7mIhQtQuU+64znHgdBLdFah6kfky7M+y7D
lZldIA5+hBGTFmm2AY2VJMRve9XyWjZ00tciaowq3j+XNjW2YHzQG8PTAkLNJvbM
fAKQBIBR91Z2q3aI8GtPg1shYx7xeEpLxVhE7cIVE8FzvOzjeaZFvYn7CQOa4Bwi
+rQykRiHbT8sfYxsEhduV4Skz2O7AuQlBbQedy1Z9CVTEde/4+Z0r051kFViH4SR
Ap77+G26rE65B+ET0shAhVWpijw7iMdWX+524ho/bfEvMNMwiVYieGGCzFGJpbF2
Mvg2yJ1Tp4cbWvTAdNm/bQ==
`protect END_PROTECTED
