`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JS6Ee/OUguv3S0KjECptSCylAVskuC4DbC6kEC33wWcgesPBmejDGAigIIRj5d2G
gT2tpxKVWxhotNsmVYaIxRZLuxTXgpVOvVu3Fee668YZ4C/jZdQcOHdUXClCrvYn
N6JAlvClrV+g+QY1vR5Y/QbvlXgpFT8gGvybYQgXIkDSy40H7cMW2Bj4sCTUlfyc
5xuoQsIYec8Qoh8wdrDXt3OPAeQLB9M37xbFbkVWycAd0dMsz7/LC3uB8M+OQI+p
jFtyR4dqKdda+KWLuxGgCzbOgBatzN1vp1mbcJRKZtttwAYNEIjqQVbh4E2wNR1F
`protect END_PROTECTED
