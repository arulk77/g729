`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
f7cgJaUcr5TaYOd0PKe5tIQ1XxXZfs1osgx8Dt32Yx5npsXigSefOgWK7xHJDQTG
hseEP0p8ctJ3Xkugdcpfe9EgLQJ0/mV1OYVmhMYb4mxTxGgKh65Dw2kkvp7h19hV
6m/rBamYS17Fc6FH2lXgmtHqj5zFDahtDSAln8im27ZMILXFMp0Zbp92pXj15REg
`protect END_PROTECTED
