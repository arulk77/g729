`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJIJkLwwmHeyVDA6wREo4y7Wbx1gAnyyw6JBl5XlFKj3
XS5blQ7l5fgqiBEeo2zcuXwYFJy3vzRiqmEvg9Gu6C+JQ1WSoJWkt7sgVedZI5HW
EXYorRTsoeKP7wqH9eR1tCNSu1a8dDxVcOKRuIvbqX7XC7FiygDeFcfAN7ByRG3W
lkyYs1QJm8ELKkFUpvJSdmd5DB22CP0Tkbl4fZjrKMN3rFGbD47MQa6ffpKwZKHH
vhtxBRwQKeW4VEmJnkSky5AhkLVpzfo9DOSFtCoOldOWOtGiWO0pberop2H90CKa
dTpZPJg9MnNW86ogwOOsQdy3/Le/geqfiIph+Ohx/N+Y2Uzksvc/oO+9raKBJ85u
bmhUWBYXMnCkOZLX/nBLe7zivBMLkNWK9Q+G6GrUk7lLtRGgmOQheO/sTbuOwYPh
QVMyGwCxu6bbWf/atcjceXUR1pnucNeJ2RaqgNNrMyLNr0dLB11tXMJcP8POhPNG
HIHIDkWS9fny/uc0O5055hP7shRpkpPd9IPBNCQxXXyTTRiKv8DrDXLuw0UZKLZZ
`protect END_PROTECTED
