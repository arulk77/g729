`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SSdwjc0s1o1oWYPuQdeA5Erei3Xf/xIhWvx+eYVeNYvO
VXDf41r4k0AC+2ToS6VoQZcZQrpnDaMJ8nH0/zmuoYdYFtbFPAH3BzQnvV3Mo6X3
P5aLbq9Eu+IIwy/A8+vI8dmS2OeKc4vaZ8CfDIOXh6VE9i0qUHIJ2flte2O8EvEE
2aymuvfF4oUdAb1JVDWbyVP3dSs+szBcCIlq1Mx/TZyWs0ze0GIfPFJcZ5N1zGxq
PMYaxhhJ4ls4x4GLwMiOOwpRf0E6ib9HHsz44NE4X6857jMBmhUQS7aBKPdvO87U
Cs3EUSV6oRfk15liUqk9o+NQy+tAcHSt8q0+gig0Wu9CJqX9ULkCeivbTVPghfUu
x3GbiBPIOTT/Kg6lONer/u4VgK8WpgUr50RVm+SEjTPx/rHbhJBRg644Nm9u92wz
Zw73AMNddhqnqM+sp4Q9UfZRHwKhSuhmlxhgoz6Oup5EAPFznCFr1BKHhYviND/6
0NafEipoEpEpdJ4g1yaYt4KEAFc5MxJmSe1Eo84dXA0cSkv11YMLPB4Wgot4ySQE
liYdzprRXY/ZDgv19wUgyqna1vkkyOhiZ32R141tZrScUm2R4q8hM0k95DGpX30o
UTl9CEerMrXuz0/Gt8+0xKWvOL1kQghGQGKbxAF8UN+iUNR0gEC/aJvRvWbQk/Q5
nEHzU0JBwV+VkMBNPS7/DPO0umBChLqy+eNiPoZzH+xB1OB6j9mFrwknmDF1kfWb
XCk63br1B8PztnP06Vck0ssfUaLAhiJi/jecyRa+LcljwquWvNoA8BHBu2xLGNO8
5xtKckV1cGhOP9b4R0dRsxFen1ozu4ZGaZ3ZkSmfEMTcG2+HdNCeRhiGdOrLBaqB
Em5CtEbwJREPMi4Oe+x8kdj0Z9H3p1v62jiTO+0P8XjAiEmurtuOvIXybfo1Qjwz
dfYmOSwCbERGA5AR8IpRSlgDHhWhWgF7LDN9CBaz/JSAyutJQN6dm/ctgjhfSKTL
eWbt1smEmyLIGRzeONGMq6e7dNw6AqeNBvC/tMcSzZ6o9EnRjzdJ5wstdnxyqNli
LViJst6zGQv/4ACVSX5W0DlNjWDmDm99TkHExWfthHMxqOwo+cVC3Ok4rTKHAS68
ShAuK/iRiOnqwIdzg0Cfsa17FFY4WyZ2rLUOgi8cOnG7ZoPsrFMfT+A1nWimJiR7
Drai9A4EjwswVUCQW2YZ2xJeMvscN/Km49uSnSViFJ9NWIw72Xbe1Mz4uXNDO79o
zuOaCISZgyVEC5UZdQHhW4Z995h/aaGjSjYgxVAJSj0KEPVN1250CeHs/IDQ9Y7u
qbkxuN+xvuyjQPAy80J3yiCBSF3WB5vT+4blVGiGAe9NlnouyMyDJPzJAvzqIpdy
4p+KZOJUe6Sp7TuOdC/zVSAaK0QAqPMoEiAkvNZi1EUXvasyI6vDQJ/twf7keRKN
Rwn7QqEc5FVbADxdVFYeAaFeoAN6zpRTd+Jx9+1jtnbcBnD/QAFbaexHN7Bsgand
NSM1mtZjC2BOg3/gR0vZ3uD1GsI4U8fx8oDa2lw6xndRFUZ84TT8tPT2Y0JvCaSg
uBI4NDK4hFzppWTR7Th2t9DE0E2U1PefWdBrhOKDo2fXng7mJ01EXXBseEr9rX7g
LaeNEH4CmJQClELfzItCK7j/iRgnlXCPbi1h4ydBaF08eybZybRcaXq3m4N528Ek
ncaUND5xpmBHWQMnLz9JriF3OpJQEboBZ5I/55dQ9UsVhldd3XSbHtYpBnBA/k07
1+bw5QcbiH97ond6p6SmEDVa3K3g3XdgFKaW0bd8bVblfTNUsoLxjjZmnpoF6prb
8uyxmuuWybIgScLHkAv4CkOhmXC23/nEP/KiTMvD5yHMsrIQC/EwJNGyuk9jlfyv
VgWYwHGyb4rq93e47mjb5zeBwmITldB5Kt08bBL26wzgc8OLgCerzJwiErvQkzcr
qxl7ZNL1KRahXCcz6WA99HhAsKSE9aaHN3QHpO4/Hg4SNpmF9x+iz9UBPyoK4WAC
6mYvOOjOU2TtRBH0jJMkvjyUF9xQUEIXzGuq9rOc/jAOB0wvIdsX0ZILHlC4h2H4
xo0Dh0qy3YwUboQhLpJFuI/367lmJ9moP0YJAb+VHiW8jfDgyRbeBBSpiH8O9hlA
EUWNklppPBhLR3m3rRAXBIOF9MCuyPkIOg1E16EMFflql2MQjfuQDL5FXpTn3j/X
Wu1UjsvOG4aQ07Kq8va2Aia+g+a0QJ8lQk39ZWDqDtuyA8+rq/OvS3uOzMrMRhKv
frNjIRHOMuw2I6kZ7QEmimHKWHrcAra9+7VgVntbKebhQ7K39ZXLvkakDgseG0H+
BlT5SJndq3Sr3kb1JZUR2IF0lOnxys+l+blljQQIQwTQO6+j9fpZZZP8T/uGjfiH
5t0YpiEkbYfy6svEWpzIQAGW1N6/Px2U24WigDWQHLSyhn3+nfY5E5ADu0KPuKqp
sTy5YFBK9G3UBR1oBZ0HLzXVqceaVRqfP+cxRRm6TaM0xeuk1QZQ/FfmrIYMeN+C
3yk97/lhFa0tSAHP5ISDVcMRXSRHVHY4q3OPEYF+86/FtXFnt+lk/D76Qtr0G2tb
48WZhuKCiz4hgVypXCqbJWJzdZc/PaRQON/rdNK1NnZWK1LRgmMSymw85KqsYxeG
tZwik+a9EaycxoLIesdT75fP1EagXRR+pGvfT6K+x3gwh148lDfkdnauIBFHwVqu
Qe7MWOG3PnK0gekkKnHDIQEEaE2Su8np/nDzluw4o4Mql3YDgfHlTKu1zw2ly1/2
KoKfPPxpTPhxfTlI9Phqj3/hTw7zhc58AxeGxmPEuZo6GiQIi8IsxSxNtexHnsbi
tRCGMkna6bYMXe7rVruJBhTCzys/lmw7mjcVWWuB0CRMYujwg7QzevLZNq9nGJOc
E01PYwPnoAFHnWbAbOpw6V3+a2Sie8AbdgK1U0LCfYp2y7HUB/BlZUWfcWC2yjST
djt4ARSrtP9YXchV6cNa9AIptLFGmlRrxKszPBS85zuQGiCcUKNE93M2IkvKpNdQ
M6HeZHZtO4CfgzbAUF+hcY3nrUwlSeTlbBdLKAocOMmxTIZEs8nH6rAYuMeNMOG4
G/6E2mro6sQcDKpzEWQ6PM9aqqeYfgt3sZyz3y9rVjYw8xqEV+nN9l5cb+w+EEXk
xBgHfbIGBsH1vGjDGcjfnOdApU0JbU2jT5+DGis/Ip9QA6LK8Ld3WWkE+DohMu8e
N6lIKXdXefbDSS8AyfJBzW/Ra4oegGPSzTtSgJyjbUaXsn9C353oV/nfee5/wdeY
7DFhdiF1Wh6v2ZkHBPJqbMeUINwlfsuML6r3Cjy7wi3Q/EmqBaaTBm59AHaVjRRJ
HFogpCgXDL7HMhO7YgPjAh/RjYL5bvEi711pdx1UY1RMjBX7wIpSYOnVn2BeOXd6
1sFu7yMHClqET6/RQIeJxHrkBYd23rCGBZoJ9c7uWx5dFOMMkDMsjrBmn9o6ZGAS
EEZoh2rKO8GRLc3UURyUnvR4NqOZWL+eAzy3YJPWpfpcwQrIJWp/yNLtxn8kPl+J
C0fFehPGiNmnqfAlZk01OKNqA/mjdVzzuuywKiUifdrVmzXFhM/CYRQyoVItD+iH
+LpBDTV95vYEWIJBOK/8uGuWN7k1jn43qNyKC9lOD/AtVObUF8iLvVdrF42rxR0Q
Wr8NaH6+PDQRZaerG2Y2Bg3ICL3hE4cgMee29OGMI46i5qCGbp2B6PWy3DvpUpQq
9EBWWFn8gPKJ4rRGZStG+GeOyhVfJRjmj7WDq1I4SLRS1CNY2mz2Yx3ZwlL1hxR/
wOQrdpAk7DEZzU77NBi/mIPSG0TA0wNTgymq7hAyOp5udnkXH5SGhKkXD9oxDv31
XzbJFb8hK2H4aXAL7cdcEimzk3NlEEuEwMY9UUL+FPaM5YCMIdFko1Rbz86Endff
nkOaY0Sw/EJvtiufcAMRpjuTT+8aqoNHa9re8CTprWbbMJTmZnAjSyV6eRoTYOVb
62GNy1WDokSq1DOXExnYNWPjurS2mbAtmkgeNWcvJnnXomVqbMtf04EH5nza/NS/
BjckQwH3SCvYWkg0+067g5Z0VIVxKfE5xxSGodOICXUVONJOqFbgKvho0WMjHcUC
oVqm+7VEVOLdqyuR6mhk2KiZAWNFfrch0+7mxu180XSsddL4sKchU03PEtkFkyVq
O2W4DM4A4Ceu/LiFZH/cn7XNkSTrQQ1gr0CEuKk07DoCE6w2ogveMdFipIx7hndF
sAY9Drk9ofPpg5bQYnXLY775/lyAepe9Ezm51R29uQ0+Cz8CAIQFDqZpFxDMwPLA
E+DUFbAjuedXEaFL1VrKLpHPih05ascZ9k8lG+pPMVTG7o4y6xaJNnJ9S5Cd5R2R
5gbNAC6dkuP0QXoBlgIKyZV2jkvfmwP/jOtK9gzyvQgLoyKHOeV8swRkRzYKiUc2
iVAjzauc3jQPl/4nZ+N0Hd1jT2/juU4FKYteVuN5FGVEWoPIIJ8C90PxmprHF+/z
ej9YVyyMQ1wb9alRZ+8xp/rIsi+VOKSczFJzMsauFsQGIRqlxip8Wbxm1Vjd4CUu
oD7z72revizWNPFGDiaMDFCGPtQSNu9i6JPNbOCMVYfVdAwcb5r2cxJwOVgIayf/
prMc1NgVvqkszJSlsahAuPqPdY2mxIbITqA9EI+PAwozJO4tcWpeDTRCCtaxko4H
Dx+BefAwm2q+ve/aV1kw8l1hyPGZp1twXlaBMxOu8u2Kl6gKrSNHnjZ+boXoXjBC
zAPWgQjzF8Z5k91Th3UriOvxjGxvk8MtFL9gMO5wMGVMpV9/VazjydTCndeJVOpP
fU1I93SVf4Jzht0nNqziuZNs4s7CMBrHmHUpmm2Rpk6a8qH1FSNpr9TqR9f4G/vG
jzlNk+1zykj9+oXri33G3WvoP7WjGd1JGvIzlaj5svOfNqmTH9w+REfd7j+IU+y7
g68qZT96KAoQq6m4FJQO5I1QzmecECddPojwLaj8rVbdRcr1T5uDfr0ru53klVSj
baeeAVhD2+iKu5eqWndWfxp7ebKJX5gVfCp2tlOCrw8FEnkEA2ZDunnNTW4HyhZJ
UvPHSZkKv4/suwDUqguGr70hPtmEqiN5T3I9/RxF5gwbBoensgXyR4MQQpMRCrcy
wQVl5oA7lcTv0HvgxZgAFiZ6dU9yn4JgsxbffGzNdjtmgyKvQ3qU84OqLIsCK7nF
CQns3UtFMGZBG6myZhBHcz99yCqUjqSfwSUfAhSYY5VG6r1giB2CQahH2gn1HiMt
inoHboOykzOADk0fzJQQIUT9oaTQXM23LUTO6JbO8p8wJ77q62onGZ/u565unhaI
wKjNLIngZDDXpFrLK5yGRcEGJJjhZ09xE1WqMsHNQlAaiiV3XW1jtu8JXWx3PNAt
E53uLZOjCIkT0xc+R/dwPzNXr5Mw8G380O5OyEJRSHkWTS0UlqoLqu+vULID6Z4H
1sFaAbHLIkI0JfWn7+k6/4mz3lgPbDaoJ7I5BlWT6RJ70EIO1tveWqvSlQH79396
Pc11Oh2MF716uLb68neyesYeG+xcxx6C7EVkYWv1XIqdRAAIZbJz2d9t2QYUtGL7
v3mmN8uI8SDT1uFaC9EeHZlOqzr3+CDfrLbQ6fKdkX2D8AhAgQwcP6UM45sSsfEo
EYQc0S9SZO5pYCh8r7PtwOveYRIjDmmRHp868TiecR70LUCHfzVusFeKMz2HdExE
xBOoXYfpULA2GQCb7+fP2oTUdqM4Qx+yrluBGCweD2j3A6vugxjb9O3MGvSbtiIq
Z51fOhMMvPZuemfO4Wp+E+6Y8mR4cJtd6niDmw85V/r7ggkpciOTxBoQwxp1/KJe
Hr0fidYCKePX0V7qu7ysnW0VtEz0T5Vuwqkn1r4q/CQv7ASYa8S/tZ2xUt+QQfnP
ojO+hKPafMCxvCaQrebCCVztORUfRcSvbS/F2zBdv53bLPwfpmElUboYhUlmUL4d
TxjQ4pTlowIRha0aVckSDdT0AfVnirrtPz9wQ6agypTpPT/422nu6/zlhNjVLf+q
1SwSh9p66NFIs6I6Qqx0f8YhYvqlUydBeK1vlw9PxszWesQie31NEC6YGFNkucsT
76vzCZUv0lcQrfE4WtkRh3Z2tOBY4Z2ARhS80KRXp/blkMqbCgxeR6svYFF1rXs9
Lvc1Ji0I40TOBl9tPfIhkYH+6Y69GamPtUjWfVY3AqR0ktjo59mrVPmj4vSIbDp0
mW2zJ6sQXSSnS5msczidp4Sf1j0SMhgNGgw7pLIANqQCeD4geEMvUiC8Z6rLG/8f
MaR+WaZgEYbB+pfWXDuXDLyxdhg9YCJovvqQsh02lvPAOrOd2x4BzAVMw0oSk/8y
H1IZ0Zvxc8AzrqhFfODrA1uQbT3KYRWhhtfaXxcfSOmQXtw0YKKd408oRqHyL5Am
44jFBZ9IHQzqTmxSMbpUgZLhKlyyZoVMix4Gt9dgpS6ofiYzxWK9souXZ4QKa968
YbCyx6uDkw9IliEY8au+OrERttVzQd15lWsNMYkPtcmN1d08BZyPTPmoGnOI7xL5
yNv6kawuSUcvk6G3oELhEX3T94HokcMSYTbLFlO6oh+RC4EFYk5c9JhjAm/a1H6a
ztl05zmOiAPKLrQTR6zZI4yD5sQfX/SLihFvMN7z0mEHVyCUjs9kjgihy8mo7xss
9rNUBUPrdFkr2WkHvTllfkgOTAl1roehli/34JsRsRavkQedjwmJcMUyHk6dUkTx
B3DRwDQ1wvY7pSEbZ8K+9YuZIH3lVuDmxei42FyU7vIgAVE8Vfg/7kO4AxQ4Wh+G
YTHxuGc37s5UawWB4ThnZRxKyQcI53sBP+ZwrHkh7FEBtevAVEOZeTGqpg9Z3EOv
tiG5DP56xxvtyXrHORgRpMg45wDOKpvqo51vuKc4hXbVxvELfBlcv2xbfAuGB5oZ
UUY+juq/aAt75mvjZmE14oTJZ+IZG4NKn7WuVvRCBVPeJdCoz8jkK9cYXG/lwN4/
cEgUmXGs0QUTAS8Pj4rf4JyJeik5NRa1gFOalxI0CrC5pDby3Y02KRnhZBPUZgCS
jtAgnA7Dm+O5NzEy4+h8WK6J+ylHW5OMhK0AQckeeQNOL6N5nbEFl3yjKqNxCRXV
hu04tDJOmpQ5E71FNVZjvHGN1AKYVu/ZBJLwz/ayVFpWKAYV/Dclqaiq1MkdnHxr
/SPnwflPbny7uKLGartYSIW5PQlLiPGGACSw2lLTc7NgN2JAKCshW3LlbFMXugc+
ZEMPemrSgK7MUHeMeQd925sGdcQUULfTCnik5N9yCJuCChb0emO1J/eUhEtnCR3B
9zMJnNkB8HHNSPKAtsE7JKXgyO91RUDRVx3YX8ywhxt+Uuw7mm3GiBR73By7wOAz
GMgUzz2kdc+XuZYU9HP7EGkRcoz7b6czF+H3c17C1effAJp7ZkLrdbTVGE7LyLKU
u/1oX/uUax/xNBNq5660ciWXpes7v0WzlXEgDDKBqIPWUct4mN4QHCZXeOXZYyph
1mM65zWR3VN0gO/SxXC21+YwQiQUlhAxzcuQE2nBfn+YkdwOPbv2M9InUnRgFQJq
Vz8aPeEsmorqjBTpVpA0ctxtJaa7lfqDjfvmgYUNUaq2eA3aXG/IVbmCDYVO3iwH
L5cACTH/zFPoejSAwqySInCdUj4X7GjmGhKPgz5xjdGcVL35dgIj/4l5W6U3ANld
fCQJtUdacY4OOTZ/RRE/tr75sfhY60eFW/m13m+GUvQQdSvliprfBfz8unoLELQm
ssWDq3ZrfwIy8ayzDlCHRqKUFJ6rTyA6VDo37a5wbg3MSOwEGfVNZA9zw8Ls4p6F
0dlF/j0SJSbpXD2duYLLnwzN1JiBqXG2UGF43Slh45t76zqgt25CDZFQoIP91Nji
LfZhhiKtEA1dOHgTfg/5/0Y1YGzS+QyOsDPr3TuhHdGW4A4dkzkhZmMDMg5IJ5Jm
dg0IjMxqtIdREP9oTNgfGdB3eTlN/sZkfaGd1ka4512LrzgPkctooGoR7JUmoffR
mHfclHmngxygDtz8LurvNISGdQLGZsHgWC2x3HqizA6s8ETsk+PE7KnhWuJ8sb+w
c11mTzmv9xN4lH2C7NPO7kpVFk2OhIcUFl7iIZDiHIzHTJcZX7qK/CzL1VvW8P/M
e0q9u3QnOXbfaPkjSLkGuMaXiD+ldUSCD1ujy3NhdApXVlER0VJ5PNy92VjBtJjw
XV4TmuFzV3e6UtaMAO4n99A7yXdx+iylZwrVwyt/8vaIcnwD9Wys3fwwGwoZgN1s
abMr4bpReEzNNG2faULx5ke2CTa04XnGf8oUe43AcoVwqJaICEreJMfkXJnzJv5U
bH001CsOq0KjOM5sbasjd9+M8KKYZmXOIMNptA//+9Z+e205uB+hOJ1ANmYp0qSr
s+/QYXnVZJjfg1QDf9jrReRtviJD0S4PzD3LLvfOKhMN6Lywuq3sZqokMRIeOQNT
2eXsuJAQaARP4hMw5lgv8CeSA1GLYD15PK64RPQIxW2h9hGmKsoPYt4q3Xz5FQxN
v7HSDxi9kseAG7tg0zUKRxFY8o1myp/D+Gc041RzO3W5EyxQdrQ0OslpdXajD7i3
guj0MwfKdyY0oi2Qq+vg/A+oN2xSk15m6g9w9q0v6zsP7MwFVp99DUcllMn9n+oL
bF1GgMXAUVJLvZvVBzJcf2uyxebCtmr9m1cqTho5mRuygQmcNbG1MVi5MhXcuQas
5Po/7jvLmnhYZqBN+4nRlbXYRCpox0b0yyE1icuoizOlMFiOM00Pg4+aYwhcRdQB
5JuPgDbrD+Lu8nmLCsiskmVZakbJCxCULYxhqArsLhMTsmiQqFiFGHeX3qCabGP/
5Tp7OigB8r6r43+FOZaPG/u0eFtYniuI52J2bi5114srwzOZJS+71cZ9OEelmD/i
RgSUQXfkoC5JCKc/rya6NApnP4l4XLU8mk6j2+EJz/TzNGOZB9lWRkgoiBukMBMA
RGFXegNc5fShSmW/20y+KXz87qpuGn/WBB6WsLAXWm864eRTINUOZTls5GzuUEDD
764q6q3ncsn4Tg+DWPP/UXn/I/2sTzfYUqd70v2APCHrtqEyygtynS+b8pyAJO37
jsMFFNyeSPRsaPQbxwG30Oe55UasaoNRN4Sp+1m0P5zi4xJBQmSrNtBtvswMLvT6
RK1W6NuEv2Qr5yULJoF8Iaal0YtqnCkMPlSOasCKcUmdpozw4QteQra5KvhZsiSp
eV2mpXalBFYLDzkE0e+RuKRoA7mvFfhd3MwR/Nr84uKf2D4S0sWmn7+wp4zkEEl8
gp6ODg76lyMGRWBiwmLWE3GkK1t6EsQVn8M+GG0sXBTVVasJY1+4Wo4i17IcJaX7
MXa+8X0Tdg5voMY2Vmh5IJhxSn52jLY+WYcUnyg4mPmMECKbkZcHLr2EE2ZaC60s
g0CtN4kJ5GNN5u0uDc8iVEVoADG2dcyc48V+tuu8mxAMyOkoWo/QgRF5mFMv8ZgU
0YewUSVmwRGykUGPppcdU1SoCDk3idT7K9ztWBFLTS7J4anYmqE4KkuZPuDLFC0q
xi6Ht0/jVlcORlAkoLkrhmX6kQ+YbVJHhaLKw/Xko3pzv3elluvK2DuRSXrle0qa
nZF1GtsHHzzTxIaQE8tQRdf0L/gcGKGpADBoPtGqnXzpm5dGGxwStNc79DapgauB
nMvq3OkajT7THZaavY52iE1vub9fcf7iKOkcgBNv6garVXp5ebjg9ruVvaFhq7JK
Tm3jWM0Z1zOgqY0kQW3KSwqIDFtoUIFeLdUkC3Pzg/yq7pULVTNHirW8iSXOxUCK
K864BQXJNeOSAlpAktIS1uxkxAcMosEC+PB2KPyDuW++3LmdeL0qEXBwwJoO4H0g
aL4lqHWVxFk/Jrs9EtcefvECxTIfc+5WsQJdCOgXuzCN+/saEXE5unBInSl0QYbR
Q4OJgeBlMtMPD/rwTmkJYmiNaUHot3dvQsBl90Lxmm/O9ecwENBonQu1tdQ9pfpp
OxOEl3r6czXCBIxAEQjgmOUXgChy9OoPSmukc7k2LX3c1oXaJJszxbgQHPdw50ce
qdXV5ZBHeg+nEhCgN49/aJ3uGKtygNQJ07WJHUWuowNvEHkUZMnlyhgwrxiH8Z+c
A6Oa0aP04+E8S4rpLCj4ijD8jC01C5ZFaqJjgJins6iBUNsDtl9fFRHgLkhfgjZD
2yI0Zgks+A3PH5Pn7o/FVf0jQCyvKnw5Pow/uy2itef2Whvs59q1pCX5TQKaYVbu
7p4T6d23EWilJrDgMEG2N1SiWz4vS5zzrJ5LitGYbJv9W5/H6rKZWd2981uJxlDL
Nc8QztlC7+4VyI9cSlQdHq0VElpv741UsQ+PR/UER0jfAVEj0VVcTCzsfAlcS2uL
w9ICCeaiBvrcmSv8v1EwQ1svAHG1+IcoyXSz7drbcfAq5h3D7APL1Tov0oaFCuZj
b5N58NxU6TGIo2zhZKtr0YK654HaC7ZEXrHktGKRAJSL801CJuzAV+je0xy/jNcM
04AoLOX/xvHhXjmFhRor40JDFqKmrfaSWhNe0nCKsKLD1Qw0S9BY9WkvNaYrVhHV
EndA8Ist6pmy4czOxVErGWvKSke1u3wPfqZ3lhNUD9wLyxv5M1eNRy8SRUPAmxo0
LHUrTOdOZe12BP4DeH8ww9BHU8t/cmBRaLUK+aGroWJM88QD1lo+MqPtK+yI5At3
1IHrGWx94qyOTKCec3T35faSMiSkpglEai7VNiF37CjCkGbFoMcSEKrIR/0AoeJL
yKrHgc3kzpTEu2nWBXiAcBIDypFLNzkC3p0CRvZHD2iCdoJMumU3Fn+rA3/p+cgb
EjJtQWTbM/8Az+EkLWbKlQat8ZUmg+5J7qRfg27ZViIkzUm5q96hNjgoUMbY0esf
XrP9rzQRC5nIT3eFhCjHr/dwVDpSv+0S77wBwWK6NIKWrdPAuNQDfUS/m8l240kT
erCjeDgSHO3B99f4zFkVpXULby89bPFF5/G8M2zZUzYZ/BW3DesiFlkmM84pGqw3
NixiIPrb6ItNmWHVLKHJllOMov4Bh820a8YVT7kpjPh0pQZrdMbBTcfljnQkoDFm
gdAkhBRKpqGllm29Sku/AonN9r4pjdK1jRJ6ItBGzmJPcnMf+XQ7j32rT0CugM3F
uw4s9xGsrS9suLX23BROElWzcbsOz2psPMffNwtyzPvgFGZzB0sqVIHfXqiWNQ0n
b0wJM1+3jhTwL9P40Qh+SYcJpFtSt0HQ/jqgn5JaNOOyAahVGJoS7z4K+nE9ekN2
ggmXnu1Y1XQ75wfipF8nJEzBCOSiVTS8L7h/qMyOZna/W3OJhP8DyrbEoEUoV4Uj
Y1nzDrFte5xjRdGJOpHKB51BFRTC4Fz4g5vq92I+jb7LK7uczXMkJlq24/fkBTZm
Bhghc9Gll3LnLX+lbl209RgTdOxECgqNdul3JqxjiazSPqiFqzFCMyU+KLQBg7bz
Sz2PAAbDcVwzupJg1TD7lhkJlTteAjKk68FiiOeGoEboCD6e/f+hhr2ngReBHthZ
hufv8dl6nJduGkD7w0TuzvoKDrvXUJ6okVUAQer0YOxXmK0AgIMXTun0Kw06c2ZD
+W8g1WmRmqdGgHE+l4Lk6CWY4qo2zlMB4KOhq46kWWhff3y9TueKUvNeg7Dq/qJZ
OQfgwF32EIVp83n9lSGIz0tft7YRd/gHIaznuKWovNUeDVfO75ci/WSLexldAlpT
0NJ3V/3cSHdX29CX29TySoWrLB5TnH2ikrDLbexZ52zcfae7/2RbY+uDRujqRVNw
9pvhPyTRbpwNYc5xogu4XOOv6W3UDGi0nFBv7KSLO9qL3QZFSTQMga7rZYqFt40Z
OAU56qqoIbpgFUCZFBSbSi5wkFHfuXwtQ+ZPWV7mbv+bc3krEx8h394UzvpaCPup
nxLuaAH5D0agzXta5E0HdQ8/drsjC0RO5Zuj6dRv7DhYf7ZpIvd+Y8ITxPkmsWcA
gFS/SEVYzYnGSXKAy+k9naAImpCOTfiSw0AuoprNNrd4Gol+MxI8tf4AToDNbPph
qdnSADerbGaQaV2fS3aUFyL9cYIK5SmxdVt9Vffoccu6kgJUTBWMkAUrwyDsrF/W
e3yInPbKt35RWLPNksIAfl81EFxBrvrnmp5JUWXwPhm6N05igWJWVJW8uJdph2gj
6GocIKu5Q90sk/z28SgRi3rdVN1vYbe2TG2IsBCvD2+ijQZ2uivi3V/EvPM0iex3
evBBQ20KrS/M6NvxMe/ZAjuPLQm5nEup7ruJNt33ZkJAHq/U/OPjqHzonlj58w6O
uCNX5r+kIhpKERNPMQby2I1jqEA0b8iQmZXN1Gtr0UM2iJRQ9SUvAMh8WJNum5yf
w6iM8cxLZZP5a0Q+1Be8ozSz7vw4HkHYeg8+pFlFMjieAW10lBz+eo7xQaOlRr4T
7jXfAGtMlac12wrCGkWdD3tCPWDPGqQkQ37+Nbo+NR18XiFaXMOova/WjqvlQCNB
/uoLh7f8ALe56VOfudO2m52u+1mOK7QoY6KsCeZRqONaGTHr+ivbGr2ol6I6EXxX
9t+JN1QScN975JQFvPEaTH9LzwmYzJMWbwMJ7zGYCUn6FsxcpFYSPfBe8addP298
PnPdcwoFe9gGL/mUkiSDuT4zRomu3yHoNOSM14miNp1ZAeF4nkzmbRc1HDQMqZkU
hoqHxCjQCyG3SwldCaScJG4ZwZGj5GyAn+1rExEPiq/6nPQMDd1bhd9LzpbmQcAy
D9vYIismsxo4rMQq5JItXDh0htHKrEntDpMgoSAKMDQPCKQHxjNafxfm3XDEiILo
E4plo2FnkvwJgv4O25kgLAjsbuRz3/rKOGj8RkGnh2rG2LZRMCoJxq4isEmItXG1
7NiCfadLvM3YVsC3RvYJiMQwI8rv8EfFOUCXyLQfXio+q/JXXMwHqNIQj8Ms4t8B
t6jgKDH1hfyDxLvzLVnQfYPegEmETZ/5Q5Jq+rwspCgdm6EwB/NsIzFKc/5l0Tia
c8o1usevSIfWmvu/dejoI0kT8QMeGF5h81nONL/XoUzqVXOo+ShpurjceRPgWDcB
aw4n6P4oyL2SjGEHOlMDlTBFN3DC2DfW+UAtbXAYua4JWlsgQcPKoOqx63VC/O6X
v4+BfFer5KweUddpaUjrkYTcKcEdfD4uwI4VAu5ekVjGp42Doj1QXuJ+GpPjcuzQ
D/3lXORlaQEqLOhOq6iqs3cnD75loGgzJlqh8QH0iyToABRZC6rgVFtT1Bn56/u0
UM1djb2bdIb6bX35sd0csI5zAKiRJUVBilFsoeBJYvka55x0i+OM9fCjSwwM62ME
iOnkm2qL9WFS2MvZv2DBt4HNBkRrqedyFtjV8M8a5ZoXYRWoMfng/00cjQd5X6Mh
odD9EZ4/eDuABNWOH0p43N4EUaGQC++FlEwUs+DBid1XYrpxqIJk4/EwewzmZbSF
FfNuUA1mdUuLKD1xEH+XVZQtTb+Zyofbu2GP2Z+Ucdsm9oA13wOlIqAxwAoJusHc
1ebyKyHp4EJH8uGaWkhPsCr4zWXLo6/C+EIQiEKEw2P2dbzJTSmSND1FMEmfsQus
pNDDh/a+gpUTgATQmNtlXb/1EhY3FWS7X5ejl8zLkJgASnNJbCCuhh7a1YKiAFBO
PMdf7ywFWan8of3Nj628chzSssk64SCEl8bVcyFxHGglCrmLp+WVtdgyyKHT4Kak
DoKCaczdzu09kkRYmbcJB84Y+TyEn6d6g13K98VgN/GEQ80GS4FB0CiDEu64Bk/0
ddoeCi/N2y2126TuejPGwJCTb4iFePsWxS49z9yRrH8/OfwjES3n/uIXquEZrDJm
RImqn3LCcZaWO935HAVSjHB0wB7DQdagX93WcBjEOXb+knXcXZksFuWP6QRTS3UZ
yz2vW4xRVQK9K5AKHm9UjIh1oUc0B+OCpn4oDAGL3L23U7WlpyUcZEykzJo60exk
Ue7PFdAhYFAygT/KD3tlyyGs7HWjIS4ojQ+ZsllVz2DnoFTwWwNPS2tDeAxXsZc6
iba7olozf3lgVgwxSNknI4JdmdJMjA3vCT92zfEuTJdXzx9cv1pCesML/Rm3KGi7
3n4DFbC4n1WiZUlfZVkQ/+2Fsc3z4fWrt6l6/cc0qEI7TVnqsMeFt7Iys98uHjJq
S9dCAzJTy8odB2dmwlt9MmcKbkomlpg7kyIm1PAA01B3qL0rCqyEcW0MUGNSKDE+
aAYXSGlYcjOkn0Lpp12DdVyGS2OmZpZ6m7sfXHJZb6/lc+LD4kE9ayKvuhLAIcFZ
ku8RyM4yqsQxiY594zONNayQaoUTpQUkXR5FECHUxnN4IZvVyC/K58Bvx0OK0L1W
XT0+Wwkzmz2+XzQdJQRuFyPryhtSRmZ8juaUmtvKAieeq/I1jnuDBZWett1oh8E4
Zweo6jzEOpB11qSo856buRKY8Vavanxdz2FoOxEGRvv1J1aJz5IUkDKaD1gYrXYw
UsEhqjhKJ1S6zfE6grwE/6YEPFEPWIcN+a61rUEHsVkdXgb35Rp4hesvztqHC6XI
nDAc9QmY18ozmH/whbUZbw2x7k7FNA6ZVxAt0VzOf4RcCnB5jJ/NmGBJgEicVOlY
h3uAY53ih7G3fTxzqAc2gH2QEHLEWrLDPEIgYiPJbybS1H8evCtCksmseywdsOtK
nh+88k940AM9VSJVBHtiNg2UHYeLwGvTBSizDQCpp+qLrZImf0dH3KBfyyB9ZsLP
lKMTiUoJ4P27lHNTvShwanZwAXu1vQrJq2QwwHDdtKq+Dgz7BILc4gp5tQT5OtQq
iI75qXvMBc8aMrVifeYSWW4jEiuMtNqr8FCs+3yR7YwFoz/qs9bIqnIiSxHxDyQv
4jMdGpMcdVTT1qi2FqknGnmggv7jXJ9exHI9s2M+9xOVr97KdQCF0pXBXpx5HKq/
KCXQG6Yn3BLO90SNu+VO5r7TlqgB8RFfTBX+VO3B59kCp7hyLbJUjEE8TpiP+YiA
7Q82a6Vk0pIe4hY6nl6LSTADGHzg7JhxScyemMI2EmoMFTjVMltTXJchCxTEWHY3
Su+Ln4TD0mXqJJHktIkX/Mj0GVVvizncRf3grHOif05sidnX7V4qrHUmqe/pFqoG
fXQhk6m75e32QehF879TBHghMTy6+U1B0Uf++Rl6q51v0pu+k+IEj1JVDdq+F8pG
AYBkvkhtBk2y1fT718qEpdNr7iyyeCj4OywySP5ixFfVNeP5uuJx7NT07uD/lHtS
qQYesIqyhsXtg4j2jBj0ymguCMODD+Ho6DhIM+A/B0FfIQPwWvzdO9VrBXsaRQbi
8rjckkHB+jTHknBkCpnq3AUV3uICIM/Dfe1vHhga0k30/BSfnZE+1246gBYoFQGf
IKGDJz7k3hTv3MjpEx+DEkJ5ZCBCsxRDL+H4fY/dCPCsYPmOHVDUsKOBo90kSfSD
08994cXNxKfQjxGEQmCjC9cTEg0KPhC2ZoNc50LCKLnPT0XR9/MZZ2z0U259lysS
Mmmomsd1syWqBpzDJLyLXvVMdfiJAyEW3MawaKp5RIIMyABv1GCSwAIHtWZx3f4Z
Ht6nIzBU4aaAZjxtFdNRYmDFX5NxFH9WPIz3lrUeLY3HhxpmA3g5CMIvv0IeyA66
KTYKrnCLrng3Jrkj9HugjtRWl9HIeIwke4u93m8bQuUqC9a/9/TNDjUF+4DryCyD
IvWJaryFSHN1t71miA49dLBdUlDe6L+h8Ts+WQYaiUgU9ddzSGI6ALzZh9NF7HC2
JYsVDAZyQAgTOU+sf4xcTkxBs6fv/JoYJjNOh83e4Auwrox3fEYwmH8+chYdSvpB
0+LHZVRY51YQXGwE1hfdauslXDnFByQWgeln8oLANYHwdRbiWYHsPdeQmGpYuSxp
g4GyV8QUhYwDLb3Tsf+eVSf0OLtsuhOIn+4++ROrl+p5i/n9/hnjUDO84AqUR8OU
nWKbeSk30KWbFBGkiFPB02oxeSA1dRan7b5yVXWl0uAPcrfgkxgfHPNClmoJwhAo
lUKLCbj1qQw3+GG++L983TsLXY/+zVqPZPvx4hfDI3iyWvPQ0yCf20NEMAydlAHe
mG5NyitWpKdULBXDi9YWIggUSKH9IX5AQGJy2MN6PGrEfWZ3wl3k5b+xptyE9W86
4vQvzTnDZIl6c6AHcUk1XtjdUOBJpJz9wEk9vclGUYUAP9cY+05eVuYOvsN5caw+
3FmrR/gh3m8Y8X4TcjXd6XAJHVFySBIJpevijCQ5l2j8fwcUTd3yYdjAOWVOcPS3
J03PplZmrAQIAmjtST7GDwEj+RfdCmSKVQl+ijOdL1vtZjmE7KXdYZSADsF75DMc
uNM9R211nyHLYL0OKV2lzBtEqE16OcJJj+baU0eR3HtMM8TuPD/PJirGS46qdLdL
5sgCtbB4VSsnSEYK05y3kxDtNaPoL2NEyfcEFOfNFMWp0V1f3HCPYjUlbT17OdWx
Fyq19UUdGBkvRYsiz1KVrqDR7dpRPTeFozehT0I/I/JKx7V7/4+aNg8BPfj5cdMb
hIlH0/QtKUOPa/3eL+vIXv5Zaj1h3FA20a4qn7MXK8IK/OKtpuuhMAboH5zImUc3
faZPNcVQaPIMKz5fTzrQgu5iR0BrpanRvr1w852UE7vm0b6XxaMkX5rhTIA/81ZE
AFfokYSmK/D2r6EYvhhkN2ATzdfa9X19dlZE8FvrQtpmYmRKgOQWX5XfAoPgOSNx
9uXRb1aKZbEeb9qzDJLDgaQf3K2pcQb+a+/TAlyixm3xFvafGB+HM6tsdT09Bkqq
NO8uVU/umG2rcmbrkaAYEg==
`protect END_PROTECTED
