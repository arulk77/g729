`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pnyY3jxGyCgnwWklYcFi/bU60ySGZRwqjfQALtbh4peRKQPQr5mMFcnnbYUzSY2H
Qz4aVdzq/lCtGFQ2d2NCF2ESag4mGvLw2dXIPmLhhIuVMAg2FuPG5/oZd1QCfJxn
f44W/fhCsQ09bTs1+gcopU3s3RS7xoIZAgaDFXCmRhZgzK76fPbENapuyjyx0pgM
QfbSMy2racYsTkO/moj+kOy6c8o4I5UFj0ohR/e0XfuyVxSd5+MVKBNdjdhUTgLh
g5Q6TsnzBN7D1oBWyWNhfLBbn6vKjHMvRn/hv2zlQi3B08W9Nrnl5qqk9lCchbWP
`protect END_PROTECTED
