`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C8g/1NaGBkCCG0BGv6j6WwUOklHLQEQSlxJXLSlR/5iR
yn6qfWY0Urj+gxZId7ct71fpElrKUzjZkyLPy9xsQH7AKhpCwtyHdUHJ9DVgu7hW
PEFsVKWAqLWEA2wr2ZMogV+Itveg+xxgyWw8APvH7z+jHxjyu41emdf+yhz1rxsR
HFyJW5xQCHPji5vz6r6j2IoMANPgmAOSP9Ofrhx+MI991Cl6KiDg4LvMoCE2xZnl
j4gPz3bKjdFQiOw3ej2cb9w22jpAsGxJKv2mSd5YmKYFqvvF2L1n6zyEuzLKSPyl
0kutbsHAjNK+LqMujtsBJxrUI4//5pYDgmDrlCswzWJleksoTJ5CGGY5clOUM6hR
kYB557klfcw5U3Cv6O53YxoJ9TjdWWE30wBmMk+CIuUH6K5ImAvrQGiDZ7++BB3p
qnCy2TvsjaLfK1P0+IBkKnfnv6ky1LKJSZZU0brdDnVsxpHnCmBVxbMbHVJx87ED
0bNmyZ21YVxlWxbi6ncg8Zqm4j1oo10dju5YwSNAZorKs7aBx2sOvFITyxq0SxkD
J6YRMsDJYXNeeIEUxrLKCb5Stgce+lvQJCbx0qMSRCMSWINDJHEwPXNeMBN2hLwR
tYp8cPTe/vjhLBwv/Q7xF2dJqpy4pBSmNLn+shApkIE2GlV+tagZcFNdC9ose7qy
qmN293d4BQmsvYlqiqstrp+q+mm/mbE+XkNxAihLMfAlGEF9gsJdrLX4FL71FsP9
O9JJ3m+immPaixrPB02FISkh2rkAlIda2wR9e2+iqAkmcSnNvzEHDRAuofpRROGM
A2T65A/BoCyhHrQOPKY8pRZJ08nuVYDzY/8JOStJLwh3hFAbOaC7oYsRF/GX06on
Ke2RU1xW+6QNvFrlBE9AAWQeMMY36EyiBL3tsY/QyHVZ1DchacV3Q19eTkwdeXqv
NiMEnhVyB/BHf0zIMUh9Q+u3wUjful94y6PNgptMXZYvBRrJzKSVR/lueZ2GqTnD
kK7X+1jBaTueRrq665YuoMt5EvJIw+VXhjsO4LLSDDGKw0OlSF+w2YJhKmWnPu0b
trRQdk77stq/LMVaQS0nrYKTojUYreniivVKvez4xK2Vr0Dp0DZ7Au4BtYxp514G
WxO6WMrTwfltUZ08d0spjfuE+xRilkp7iJxtXpJTcaf447GLRIvIdrE2n0FFi0Og
asgkRT9/JGKX9KKtY32ojtxuws30znT9Ud4QGiU+fYhB2SYUnrk6yZuFAOIkZ2UF
oNo7sQB9OpUdqB5FwUWFXfve9/6NHor7VzvJpwWLWUjY4+sAyuTCbGxsJ5YMxvKt
`protect END_PROTECTED
