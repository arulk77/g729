`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJNChMCivPON1fMDrlY9UlWv0g6GA+9uCOW5/WOWs55q
LN1nHKTHqfDqwT1Lxd/NfTygylv9nbwx3FHTGDnyr8bnFBFLxumErQQHmD7zsFUv
ni8M1tuye/0fZgOwRh3SlIgicoyF9RSYdFx7SOoU7I3QVS2xbkMBoh11dOOgfbxI
WC38z1C6wl1mQG9mKl13Ndue8Fk8ly7eEjIlDx4h1Hhwsgyhre8v+5ZEwDJEc8bk
C/Hckd/x69dF9/2JSBo1y5OOR7q5vJ7oHgBsCgXMdnbOS0ZMpEX8uWTAushpUS2F
5RBVR0EHpjhmDEYjRidtP/y6o/wsW4vrIm36vuMceBzxSpZWlJLf7+LE8C28qsnF
`protect END_PROTECTED
