`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJPECNeYzxAa8mlkzhj0OqrUOs4afOmYGvpmGkv/f23h
H8LqNeOdebIh5dSat8iWMY+QUWQScEAdfCTH6r6xzAw8cTbN6qYiJi60EluWDbIR
cWvbse0LwKbwopUc625KHkYUFsiLi/kvxI1UIgUwsEojCq0/PsZpanxZNRoeMqwv
YVSgXAluzCLaZKoCm70LiP1qX8OxuK3SMusX1u4q+HAoSP5c5x1u98vdhleTye4v
iH2PrN5BOZimuvcozqhK8v0XzR1RI8O0vxRFKkI/bJkQT9tk9uHfbN6Ixkq23C2a
+PHyNGW4NLTO5++fdgqluDwv4KnPyOg2JHpxdXSQtjTKtApbPhQX05ZwnTl9oVjq
4s7q06Q8V3Z2Wr3dbGnZPhRJDhx8lAVclFs/Yj6m+9+bYlYBrGELUSpXN1ibJxjR
UtFm5NVvGEpQ6GD+11L/gmztngDv8C4OFy5RujSSt5CvOcTNvcmIB4XPM046R8Qn
YViXt4snabUEfnKEbmupA7OfgxEGRsDDgAwlUfGKWWM1asvMw/2N9REAEgv8D3vd
C7fZljy6MEA4XwyyWfOn6tTaNTa+Wlv71Y8gU7EnLV1hrbd4LHh1mIscGdsNQbXM
kutTBYZk5gVbMv8QyLrVj824/IVwrFp1bI3T41nHp5gJrgZBmMnUt+VlDGfA7wFl
`protect END_PROTECTED
