`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
lpqYIUjoSN94CDZMjMxssIFwDGR4qyeeSfLXi5T10rVnY6H0vyoHN2eVzmEMtzZF
KuiOPl2UCgPSBhTDUQiz6esZQdvv+n+HtDO5ti9SpC3pAuJ7SKv8NRCR52exRZfe
w0B8clqFNY6qfEmVwXw199r9q0Sk5lO6CqQoqdkZhxz8i/BOhsFI8rlbiV3s1MwH
frpPvh698BglD3t850ZrNfMmjF3o0SFrFkt3Lfj/fNjOdzhTtmYO/wahNN38DJBo
yPznMlJJRBpMsEZ06hQ284RpyjECmR+UimrTvldhShxETze/oAVHoO0RROiXRBsZ
`protect END_PROTECTED
