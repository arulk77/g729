`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCdrotuCEtori1Nhcs+YKJVcFBhVpjSTVlH6+zBF3Jjj
3iiAYaURx0aIyqtFno4z7+Wgbvwxi+m05BglVxShXgGC/j9cSOHCeB3I6mIqQyOQ
iojq3tjcAkPCavmEM8zQmWSVJwSiKMNKuysRLpImJluhmPNc8lDH9wInJhlWO/Jy
32wl6b8CeHAfL6yNqknRabdirmNv4qbsx7mOpyI8IaUk9OeCklZpIeZm/ImiaZgy
bmHCUiTjmJ0EGAmvyWCw4r7EqKTpKhQfdZI5ySaFrx2Huni1bYsmGuu+PsPcEKeh
NiIl2ZReFWJ8EMO2Rxq9UP52y5Nq6mVUHSbbn5vn6A3mVAUu2EIXRhUXCRNAyPqJ
`protect END_PROTECTED
