`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIvavP6zYu/wsJUTVCrFo8jwD0at/S/5pJW1G/nPmWzC
lFYhe3Cmd95ugCAR+y6Ek1wAoFPSYesbuWUu0PgZMik7mfRIL1yZy37PLzJiNNiY
L1o48ZlwbAooiX5FtG4kJN+4lz5oXzdG6sqXN/+8wIMLhIuFAkg4rpoySfliuh7Q
rHDmJSvaedsi4O3SgUZp1A==
`protect END_PROTECTED
