`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKgPPS5vUcYsUuLEMcxnHxa6u/Gp2QkG7a8fJB7HIUOx
pEU9RlttVJffXZx6q/1Qm1u23kayebzYtsdGWcqvDGaVH0PPnoefEElvT9i77A4t
NtnoMAZJzSHYYsSl4IlSLuOv/kQrffyebrQ9Gg6+e26eAlxp5jdoW68iEOJ88COq
BjbRHnDtPPnL2SCjz0iim2qZabrR+lX0lFF1WjrjGWG0pYs2ByleNC3f1vCYtRFm
`protect END_PROTECTED
