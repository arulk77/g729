`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1achBXgXuCaO2SzKQbjjF1iO4ZJQEdpDtb2GW+Dyk8XF0
O4TJ7+4uKedi7aN1juOOlBrN1zaAMoihjEb2VwBTnlchZbySLFI1o/3cOm4i2m6j
/e0bm4Dz1sK5eCnQK2s9eCDMyvAmnPlTT0HFNfq9/TG6RWicDduJtyjPWBUyaX2p
opbVmgDZr4IjDax6AvkYVm+4g8jCXjhaCTJNnV8Tta6sRfg/KjPk5DAAuVYmt9iU
TOl3actBqdiZ5omURhomIx1EoZARG1fXNEqo5VfcByMUotRakdqWRCGxzhwfMILR
+NEfD4Ai+BVWgCe8qR4OhQ==
`protect END_PROTECTED
