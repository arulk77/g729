`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAKrY/v3Fcuxs2erZcMXf+BVJO5lq1PljqPioRyZO/qC
wbB4tM5FQq1+775F1ds+BSKCf9EegrHs2r90RWWq3Iffc1oF7WzdduvzUkM3OWwD
ntd3fQyfF9lzoPXTbfS0P9YOmtpjmt/QmbznxASXE6jX0WQ+59lZsx+vqCQTPsFJ
S/WOF8PSxR6znXipJ57ypScPvjLJtOIUVgfiJ1kctHguBoREgeGrKF3Z3VSFAQ/k
yc3P724CqkpO+BkihSsqrI7vM0DUz4pHIKk5ckue5gX7cRJ9WYKX9NqCH0Hgvbjz
zy6rOSVSLBShQRd/VFWBwy+esaGCzGCPKSHSUPV5UXGqb3tulKhvKBu0fJXBnSFs
S21ZkKkKKtj2UgTlK/zz3hQ9Csq3yskKpzIcRTtTmn3OcI+d3kqVNqg6FqXXWxLH
KvFSwucdeJwEOUURCUU3m8cyFaOqYeCyX2RNU1Lfrcox2IWCmMPabGXjXZiIomnZ
meCYJUGqLG7WgpUfNJ/9LwTn+hGBGtqFvhsQZTGW3e3eU93I15UxKtav3m9734qv
HJLPwHyHPEOi2ippjstrNk7Ewjr5iwLTKFJFaMJenk0k1mzwfYHX2RWi2bX8U/T7
mJt2eA3gdwY8ZHDRrPW3LtJj0ceIc9wruWl1TNye3Jk4+V/IN0xx4VQasIe2NMCj
1dIZo0Ez7hhtbFLm+KiPKT0nU0rXp9DmjVQSB6JYRcVShonPKdf6Wg7q/GPGYu/A
yTeNbxfAAv/xF82oPpwPv9JIbg9OMt1gjeu8m9D+oiHgYmPSdzZ/HCtOWKZetH6W
qFPjAvec133si6szniS0hg==
`protect END_PROTECTED
