`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDNDm7hteWBpIJwJ9maQfUpZYOcQFxcFVRG2Mem5vmIi
78fozgs3Jb7z1PlwoX2gC35PmbD3Q/ddZEKcyBR/IuOys2aySFS5payzqWHJcmB6
kE4a8F6t1Rf7bwyEnFbnB10QoTcHnfON7DvTznROG32X/WFhRTyHFMMjDwEcbxcq
FNlTc3Q0uV90rFR7o9v2hiWb4UKJ/RkZDqVIZ+5izli1MQ3HyV/3Mzbw6xp3bUFC
ZrsUCpsYc0FJHN+BIqh4694ZnMWrpKMQRQvOPbz5u95qZvxpsiaVIfuB+DvArjOB
HVhNWHgjUiBa449uCR5n4PFiuD2/IOVt/+DKMkT/qOJVJym2nbiaVTvN8C1gxZe+
yfUqb5lPLbHazzHO2b3YSuB6/bM3pDf/nIr3kn2P/XJrHBjCvxT2YqsJte9Wp51b
zJgB86Z3l4Da9Scd/dhZpg==
`protect END_PROTECTED
