`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
9HEWNC/XJ41aK1wDaGms4Ktu935eztIc/kTZ1xm0ArA+OfiOvgKcB4gdahWTpZnq
ye0fk/K+AsW5oE7jEeu8EG0+BQrw8LnLJw7oNFasSWFOF4LduFI4ODWkKzGeDvCG
VoxeY3iR67HXfwINb4KOOCbXbMNNFjClLJjyYG4hsqFxBjlKuxacSTP4RLss8nd/
22TqygM79M6wSfYZ0OkXWaE3Z1ETFbM5YnTuCVRiVZc4at1SenUS19qaviw9z1on
qVkkJwiun0PEfQPqE7jCFukLwU961WljUMoGazlTwPK3zh4PM6MUUNMedRkK0id2
uCRs5S6Wb9wjvzXuhqqP9alT9EmFImlFwQRNftX83QWH0/ZlXMaU/SWPuLiX5fcy
v9iAuhdDfsj96eJaT8gwRUJQNmIjCQjXezXwtqQPHa6GVVu4TIPNArqUHrKeJWZK
gK2LVSSV97CuMITlj8qcMrY14IAlEp2CE4FDuXHjmhQiW9t9R79UMPJCgRw4KxWN
6mUBRZB61PscwJ0+O3w3VApzMo0OJ8busBEBE9EV9dZFe1L5z7JSXZadywZEooab
Ef13NqAxrBOCqGFy5HuYmx0m+drulCjnPJa4c+C+oTUciouGkyAbb74Ch2QiOg/y
J0Ah1ke4LebQgBE0NpwjkvSMTzlhKm1ixjhE41A2fEGl4Bg2iDtIm9UU8RY1I/yW
IzKBtpGu7J46GhCWcVZ7DRdD6uoAr51Y6SrvozZ4f/PHgt35yFcM9+n6fiuVggOZ
rnLanlBurf/34eVJWs0nOJ42/g2fcQD7OZUn8H6WjsSdVx2wDXMhK0XBrpm8noIF
TwfZxgTBuWlPTqoTCmvEQoYjPpNAtOvdB0FKN554mjRGoSZliJcAFH0Lh1V6ZGoE
0npwDP1WUI387jZnUx77AEtLiZ5bGezncW02P9+cKERj25wD538SbXRiJoToPKc6
E4eruqqLcWRkYg0i1bVxFGaarxUQ3U6+UqadXBoUuKo5uW5ji0onBfKbyzIT8y16
SFemreE3aUhhI9ROE9+zVBa0Dc1O+dGwZzRsSjma+dE9p0dOe5D10ULwyKZboD5G
jFCs7vdr6BpJucCMBcMV6yubCLI7TOhtERpIuAycvSuerHpLv58VJbdIp591wFtv
FMYFAcqR4BO25dUh1tQxWhQaoVvY9BOhAhMQXIdjVUda+JwrbLzG9+ymz56ulx5u
Y3lUForoApvITfc3N6++nY5hlUVTkiAsiGkEBg6Z+1PE4DuaAzxRh8Tu4K8JXtM/
yERIkBRk/ovJsjRRtzX6FrGSS596FOy4khLvKxQryPLX69zvfkE+TAdubunjpyw8
Bd4dlOsTNql6071VL9VIPyAIe2YF0B6WVKzxUEH7PmUS71qnSU4iY0OaZRNd2PE1
ld5Gdp5yf6CCX/nn+zxWJyIJwgjpCWf6jAf/OaOCTSPl6usoBfJ5JykcOSQQ8A8+
5c79C6vHzxiHL48NxwqF7NqyP0NfJevTXbW64KkXGAH70JzKdw+98euDQ2VuWgU+
HpnFR3CHCDZDdMI4L0EtL+2ufJRXO7w211wh6L9PfLfwGarKAC7sSMeXyA03ME+l
lFgy76lFM9g0CHki1tB5fqduUV7wNPn/WOZfO4ZtMbd+vd+auN1Xp6WgqPYHk/SC
Rfpil5v8XVeVovN5NDyG9AjBJhF2pdZnl5CfIKPMHdh6DZK1i7dRA1S0YwYE0FS8
DphhSfM/8tWc1KpDZBkn9Cfpn/KqKvVzusY3OHHOgX3zLPO+f47WgezkdqGQ7dgt
gLCDQBSKMiObClHh5h+eNJdamND3JovGEuW2BJPbvITco4olb4UjjjTUxCGvCEk5
s1LP343urzQqbwuIA0m3kYGBqroi7GWKOPGYPYBmd6TJS1crO/niHU86HzBSobOa
snXhkowbbrTqLNZQEStlBuzC6qKYCQVdPLVcMlFZiEyJdJ98Fyu7Z1Nadvep7cjN
E9qmvmlaOhVTpceESJ6PNmpg4i0QahA/JNb/e3nw6vXOqToib8HGtOmrW1ish9ue
CmpAc6qV5ysTMnPjgUq3+GWSYGJ2PWA6P9P2CHz/r+cjVmsf6AgVrWZVLFiLiFJC
WJTUeS8243sayvS2Nw79clTuk7itHXdcp92iNYVFT0ISur1tSV5AgqDiklKWzIP9
hl1z+u2OlLEUB1dcP9j/3aqUwyPkDpTtsAJwdmVf6DL++tab7hjTbSUVpp9Oc4fn
6u1uHiDOqNJhxhJr162c8OvwKnEwmEvywvAS3OttIeB99trKkf2/2uIV9Q/Mrpvn
T1QUjS8N0YYRdfESAA4ljwDJ+dysWNOwzK0+avzauxEFled6wGh0Ruw7NvyIUK6e
uP54yx2t40dkeGjxLptx1pgUbvptkwR/pFGPPCXSSrEXBscK+N/CAbBfrfg0cmWz
Gz3zNmZXdmYbGMKpH1M3nBwDtRC3K+N8bOwFKUOzIJt/f2Rb+1t9IpXUz6F48B4y
tUCS9KbhRa3JFkIZcpZiCakSZ7v5KWQtglcDNsx1S2miv+eiM1YP2GGrl01l8vNP
hj3OGPTqReQRS09u2GflbiwA6N8skq3oSzDorGkvhyn7xOOyhWb7O0AwT24zLatw
h1Jp+/MStatUWDIczdpDP8iQxlnZao+x3URAScN2+MQxEi2ud9SIGO4fJMupy/F8
PgNCkErdE4d1R4zVLjOU9tpnCK1FeLav8Uo0o9LhP5nq/j43kvC8kTU0rjk6OP3x
EFFn9v+BSlgRKFT1rLGynoYphzWIUsONmdGRjHppMgcHlBOztCOwfS71ztV2zxqa
K8NxtrVme/0serLI2zSzRu9wRokWfmQYObr2RdD98kHjmVPbKJr/f1R6SPmDlLPL
nOmEpa0jmxgU/uNMEG8zlwn+vHxtvEkgmcGyxN06hmEG18j7zvXVfWX8p3lKLGOt
oLhZLcm16SW2D2gxZL9s+u4f1PCLiKVKYW8ONTPNyqYHwd3M9M/XCg13xmE9jja2
lxmJFDHYjXhTuykCcd34xpJkBU9i1xc7vwTKx2YxzCjEjcWJO5FQW7tNGRt1tBpK
kbGDEwuAFBPw7aY1BdAYZxilZRvtlFA5gKx2srsqlH62sm5SbqTHAd6BJcUKEDnK
ECR7MK/dBfAt1665YjZwLLez+sv2+wVaSpRCN/o1de2ur3Ea7sV0n/DB1BF0i4m3
NcyLw64C0nsCezyWZbzuNIlrqom/BPNjWi8mFEoip43tBa6D6EZRCZA1Khyy421d
rO0XVxciDKdN8/y7gNjAkN6yF2jz9qURLpAGZGnyBE1mDhDi8FkiJ0euOUItfogS
kJtSAruNQUWtnOtM7LfpMI0au8rhYohPXmcwfmlaOMmjsYJmh3DiSOy8660EjhO+
1g5tjpF8SkaW8WGhnYwVwxu43FHhgJ0t9ap5X4Oiq3r4gCihfAKWPLn4XI8LejkG
IK9ET5tRHVgaM5ldjnowivXpsxtAYDQEyavzS2+Ipt0Uutr2f6TEkTSprC0qAVbw
4z+Vrs2deQhlC7LwnN7i9IBMvkBxfeYpmpT2acsJWg/n1zwtgJf9jHBANp12pnfc
8Udx/FVjZG0eRJCxr0AT3lvjFMk+oHuh2ZOTKcrkYhE1ST+jMgyCupA0jkKtUser
0ipaXpi1xgWf1qkYvXx6eqtwo29gORJrPVE8YH93nRnsZ4Rd/Wc0zlLQIH9einhl
bQ6KHPGbwu251Hq8sQnuh0+WKXW6FiuQCa1ngxER/YZGYoFLl6N3IXmYbIcEBohr
GF3KsWE30WeITlCoZFKse8w5mcCe5eL63mqbwORJIZQFoZs2KEQLWjjy3xrSh0b6
UmeTlgE6+MtDTUpC5BEwBbg9Y+qQEQWMDFp9eV8ScDCij+awc+MLZSKyNW4B+M7R
Qqn7Bl45xDdTgIElkYCWt5f/1FhRjQfE2fEeOI8i5zo+XEt8vto+K3UNc7uRCOxb
QVkBHortad3wWw4Bm1Xzg9SYP+ilBKWAU1T873LEwil074dwtwPHzPnxLTIRGOjH
o+lxP8n/3+T2R9Uge1/LZJuSKfXpZgCmF1Hn9ZmM0zRFSkLwxzPlgN/8Vu1sFjZZ
OpuO6mUHlTejrWZUbUrETzd25Yuhbiz4WYUUEv+K6S5Sd/J8H+VuRUwrlTej+/3P
zy7IAPpZ2S3mfCH7VEXcffTsOJ6DbN9opvmiPuXIJ7nbjA+4Vm3OsXAKAsTin/pP
xiLzkup4ioYXXM42qGpExYBSim5YOOcW9pzLlFOQG/yGpK+hxqHY9lsjA52FRXIr
zkgNyz+ddzqgNmZd0AD0jKngQQBw893WarAQ8bk7pgWHDBtqrE1HjggYenmc+2a7
H6ELToPd3P6iidjuhs4GiEtBp1FP/4S+Cc1Fn2+iRdnDmajenmFxczOcGMFNzOjx
2uvk9NGsbtQuZoCoF6PoiShTSh0bLc+rmNDCxyjvrLpkToFXO3iXkWJZtkIhT3pJ
XVfjyf34mvivJNDAzmLPdloK5uhhDxR+fV+wIcxRMY9wKdunPVzlM6/aV32n+TX0
otGdYMx/2ZyxLLG7lzV1Fw1PXsFQwJhrrxU7H21pRp8ybZFtctgnKdvFoyPklRZk
9J7IsjckrDn2UscOJ+LSakWudOcyXusiZ5rYyJPVVh/uao3bB2CRZguI05rY9cDY
pxHBP3gx3QWjQGRfdOVJi088EHEMlcMJAxAaO6xjv+fr4yF0U/jUE14bWVXm8+/Y
FK8vb9eV1Y+lywXXSx+fLzeipBH/ox+BJWk51NfuBqC39y3D3H/ucwKboFZ6499Z
3PqUUfYUHpXbnJuemOVrURp1EMNo3lpMji+DEvvw8DrS7sew7jAJAL27OewAeW/O
MHdp2OCcy6xYrczBdntlJe9VOIsupZmeXUVhw5vu/JAoy2dEYwCmKsyF/Qef5zB0
9BWBp9u4WW81MrUv6Bp00rluXJV572vcV7PUA2n8dFKTX9h5236F4y35cHW2nIW2
X7T1ElcYuHiBXGMhOR2nljhrB/7Z1erZJQ4IT5x4eSSVF/togPHK9w4ANudHy9+T
E8cSw0FQiX+4hR2Lw0oJgb4p4Vyh7jasGNQ+fYx7Jj5nQe4iGOgW4UnVl8hvN8FJ
NV4iQ+mgkN7mDq4mTxvf7elsWLZ1EhDetJFJjuLn4itIrBce5QxOdnuvuHI44/FZ
2OnxP2aRsyFMT2VeQcH+v9b1exSULMVWou/WHAtbri6xLFHyjidCTxeTPr5xYGMK
9+D9uJM8AWW/JcYJy7CmkRDvUfFcWHppgWfKF15AKNCUJFU/iDAxhIj1tiHJJZRl
7GHx6xd9H4Na5pG+LbudDLTdfeAnZNJwkU+dOZQbTgCuicg9/4bpOyhc7kglbgeB
V8+RN8y91AZTUPbhM8YGXkwccPdZI/1Eq8kdsC1qioKB8OamXu+AVU4F8H4z62cl
vUMrDjqt0zt0r2Cw7ZabzHj3FuwTbAsBHq1woMbhCWr8mMiKZIii8yzqtKx1XBVb
m3Xg/U7HvCkSKkmkru66xWq2K2gBv3WXf8EBiwSeki5ijMF5Ms0MdBpNs/PcSgpR
Y6v6Xw6mGhyLprWI2OZlBpVmWJrZbh5YIFz6YRiG6Ewmqa7cBVeAiqKnwwjwKpfR
qo8vNDMt15a9CJRE7VEZIMom/L6RnQlGH5V2GacbpY5BWjnMUDdG+Zp5nWT4uhDg
QgEEW+1Wat8uGEdTOx3HTplB0uJK3tSjWFxTp3xtlf8BoaAfsm1uHFi/j+I75bNd
8ybmEUz9axRtZuP9F+xsUdJDE3XiokDWtdy61qOVG31WyeMHVZbPNqFTPsnr48+G
3ni8g2Sje9oPMUcO6WejvoZ3su+1g2GwB7FYTmFCeD7P2DlZuiQY/8ltKK8ogmfM
pHoJvMFGlmoXFt0TP+PWkartldWAv83OLR6YtXSCHxusMcoYWN+xuw/AGmx6Bmyu
VYsu9lhOJvKuWBBcp1HsxpKnhJ0s7+WwT0aYB2icD7klOzJflDsj90wTHApet3cb
C3ZZhLo8oLxPXQp0nTFqWu8QAxfrcFSvpZmpCaVG0n2EIuW1iWpUGUkvzH0vX83w
NCOzoFfpirF9uOMFTCorHMCE+UmAvDXfPFH6wd6A4Df+U2f05kisx9uhZpBygSCA
lKOctHM5Z6G4Ys1D0fMkmfv7Zs3Qs+Fx4Ux/g23HrpTzWH4SH6HDJKknS7+Zv4Mj
GOp0v9tIRf2Z7tnninHWFi0lHGmmDjeRYmwGV675eYd9wx/mAcoRfSKFZ/jvedbc
SNXkQX60N0OgFu7Q6Hk8eFAVpbW4X3hOFvRg/08yYyH3q69EJP3M7jwBsNwcTiPr
ZCQfQdMF9WS6puQHc5VC/qWpdJ6cTYCHfoLBe4XIWyYYu+kQPEe+slFL213RjNnT
WOlr0DnigKAIxygm7QXPuRmcFvKgQTOetSTzoaCt8WveI2NDw7jfk0RttxYUHIqK
rSsuyqKqioqEOFhM5mzRoTMzHGJZ1sBwN00LpuiNtbk45eMadkkigH3M7sTRb/Va
QD4OO5Fg0Mmerb5Nt2iy5FOBFTYrbxRQu6lg1HxkBKDk0SWatndV74Cvbfeeri63
GtWTECX+9QAtC4mTPE9KDbuIzua6lvxoGbb6hQFaW4SBMcUObvSOsx7gnp2pkwyE
siItiTtp64aq2JIwPG9En2T2Pm76Y0mUr7P1GEQl1NyWnDXP3wx/5c343edVNdp8
GCkSItBfodnwF6pOUYkalCdAdyJoZ81if5F0ez0b6FmHeM4YUMS2EBjnzvk3g/V6
hT0NjYYvyRbmywFvHDqJ64X5/3RPqz9O9ar2Y9sho//83dEBLqwTUNeUfUlBPKpi
KpkoqX4pJrR//9FdnQViHYEyEEFINp7Jh7Es6R/ibF2czMuPBtDhz6M9uMUTLxp+
YOorCu8MhZpnb6rntHYEjvVsy9wbTT6tFZ8ZsSTe5I1bRxawIaGPkbLOSm1VHrWu
yBP94Ox5TyBX/ZiuAR0AxlUOwfe0aIKWh5vhIPy8jkMQ4lAPvlcWafM4YUlUSWzB
vNJfHLW4PZOEJRD2nFG/3q0+IjbrRPI/CLFFa5u5Xm9b9qA1TNUDZ2LfKy9ytOJz
LRFxuJn/AZraYZrP9mZsYq9tgw+lLHpWdUWe0+pJBib4AH1wO1A41Il2qJCBK8gc
iUi5I1+2Icz4BG++Mi8RkAqJVK2IYQg9jRW8otJR4N1DYDf3bcNBGQOoAMsrsWoD
IuC7GPi0wur7KcaRvBPD7XweM2zhHm6eyKD8mZZ2rXNHps5pAyB6dG60uqnXsMC1
zpcOEI68OhxZXRNP7oAGjBS4za9cK2V164uHgB6gdh1zQd9AIl1yPK76YYQ6y4uh
kEsxA7n6dHzKhGRDjaBtFwUr4mgqQk9aJJkVGTz5CTU/zO0JL6ksEyw5KFgYUsoH
7mxmtYx5YtF1P/tW6DF9Z89BZByywE9PsvSW4zZodtezc+99+maAMYEQWMR1WJMJ
TQlak7P4DHaV1mFh2Cv8Ifz76Ndfs7QdZ4CSwRkSczWUY2imOnHQ2dnObjNP+qcf
ZCmDrk9IasXmmz4vPa6RkOiMyxVUVKns4GpULnU63X+lNhFvnz20nwBmFK/wMNHa
Yr1X19fPnbkrgnzPoy2+GH8K25StxTPA9eQ59jcpRFUSYLD3xtR6G68et5bFpi/G
kbJjPg3KO8OLGQGysy+l//eYl7d5IKP6wmTZjxvM6EtYeZcQYxend/cgo3xAVT1s
GVwZPrCh/8AXQn6xYCfWWKlFgwkg1/LSl6ZeS9SAsGCOHXfEH0VYVVqpE9psYptv
iVrcqMvpvWK7vGxSWDAuckj3mcWYg1pjNXYX1pgex18JUHmye5+dOy9hC035t1Wk
9qpVQO5PJrKvluybGclOYSJpIEFz6rZ3/OgB1CjLl1K19npcqhD+oXfodrA/fwjf
iIv3dn/eo5iOmAjBx2mVhK0MycXZ2bKFCewN4SET4CDfhpTzck7ezTY77mrHn44/
EnG3v+dT81UnPNdB5w6RPvlj1gVUnydGpJ6oW4UqETjkGkwZLOiB5+tJplBJy+aA
oJ5y1fNMZ/JqhJ+DkPRDd0upLhcHxpFEVSXMvro6cWdQ4H4M8vHRp2lLRrbVq6js
Nx7lelAhwZWS1Vx5pgedXCHUEhs167Kk/+tCG+wjIxzz8EljQWd7pDf3yQUc3Fkl
SUR3Ik/GJZYS/Pamljo6gpDRqrDF1UKwZKMRH/sX6DjZ9PrmwzRbgDGILWHrU4rh
GdNDXqniBPLCeSOg8MPFRiAczY65/K57uwpTSB6vkAPngWa0gw6n9sPxpdqUvKZv
kRMuyc7MpNUZMYZSk5PySDo6SAfVqkSUmcNl5EhcPEVVKa8C5cmhUN1ij+4iTtBY
yJDw/fUnTzkpIXfb8L2548KGAmpWibi8Qjco93WEt5EH943fKEr9ffqflDN388hb
ZBUB4KHvMPzul9VDz9sYfUSFI4+hvWyNBtgNcv2EmDOW+X8Q3sdSgHwsXwFv8CIv
TObkP/H8m+gNKuNEXdmfqZMPjK/8CCTkt6dw7SFMuk+Bbt86EJHzjfosIGZse1JI
FhTSi4ysE2rjsEfFmK3mdmWH4Fa1X3uw7cNekGwRZ2vJPJwo5ALnzb5oYGLx9U3v
1mRPnudXkF0XR/u5hWqChWKR135igJcMyPNA8u5SaQsmRbQLAuw+vSaEpFErN/5E
g1qEbfBVu4DWtNRFXViSv9DLvrR0yPOxzx1fyLIQYnhy3RnIdBE6K8N2GNvr0eY4
vL8NNZp1YRkXvuQKdGFxpz4vxVja2qs8lJWS0Th1AUFHSBxpE/3M/uJcuPya2mqU
Ro/5InF7KsEAFF0cAvLnn/I2OLjQ6JtO22X6SQ6us/B4AL17U4x/BKrbicOl34l2
KLAD9W4b1ev/c3wwH5HEcxlwj1v7geloMIzpwWOA/e3hoAKM92Rx/K/5hQAAHCqy
zvFB/I+aFaRX/UP35q5HO1Ny/gO/W6WPuAYV6u6eKa4xg0xtq0M7F7UnUAD7TMJ6
xxlNlaKH8zTfUtPgOcq1AqF+Y/HMACGOuOIKcnx4zJaJI8iSnR1lArGMeRJd793M
02oOxGTRmWtjVYApVFu+XGgvr/fuzVZNl4+HBLYuPKgdIXW9oO/QujL8p8wd4tJp
N2TZxc2zgyIPUERXrHWYpdVbFcUr1PQ6FyPUX8DSFmrAFpmTg67SQZ4zVrvRc66K
rR2sDuKypNSh3/XwSaygNrWhXvBgoT5dN162hAi/H+SAFl5xFMPlqg6koaTp/84q
dSzOW5D7az2+oXkJ1neZMZfD0ooW7mVUGMrn8KT+jpC+vmYWi55+qUAMskf3f8MW
u3EI4+qpDO72drbIody9e+AyXAk3BSraH+64+00PIkcxgUXWxFqG+OBKXUhRnoJq
M+Cr3QYesRErjmIOtni9vYQVcDrAy5dj9djGTxqU6RXP1KwfCWdFV9MMeH1xZloi
hDgBA1DXzekEnDwRnXyure3SJW3diYlpWj0h4V58KLLEkBkBJgEJk6yDAfJ99VrK
T3HeIcArjW6bTPhZfqee4Eh+XkkoX8AJDzFajdqgtvrGQeL7eDXUnZPxWhc76fUc
naGtiF8XRx1g0iegnHNbMRcWFhV5sUH8CSPw8E9Vw8NwGFYpBz9ndy4QHGMYQ5rH
tshsSvZ/dp+9WNZAvWxohLK6bBIlS9UYckHHRkLMbKuflqTV1lDC40DLNKatVxGU
F8nWoMDdkO4o+b0t659PxCE+XvS+bn3T8Hzk4EpbC9XwYBvS6CHjhquXoQIQRLNu
SprnpNHU1LhOR6JtfnekKo8DGcGJ9hY3eoxmtJZzVifM3cLt5LF7bdkshrrZDHXN
CFB+9ERpmemzRPZU2WVlwqQ2hSD0szyxCvfAn2dEc6/bh4glbUNiaDiQG/SG9T6g
7Ig86tBZed5yCE7DXo5jXlQPqrKfv8SDrOtciQHgYvncc+WtZ7qW2Bh4saF/jx+K
KyqJ3eA2wbuI+Cg9qFicAbhRvCG71qj6cNV5Jo1WLsZfoVnuh8D6/ynLnTblMios
6CNk/heB1MVR+BW7HUnlg0qk3fzScxXSy2F7T6ncqx23cWRLTtSxXneDuXpg3Fn9
b9vimBF/5MRVzY6I9YGCG7ULRuGG4j+WOtzX3eEq36iurK4cf5/pQtfv4v/nS1Wh
7eithHbjNfGFJZbUtvLk9dbDCsMcpxI+DUu00By3lnIsy8OG7ytOiR4jJ44GkRvT
aEh2IgtdEJNpGtAA20Wpb/RR/stsZc9vQv0KSGgO9DSkGJ1PrA+jRdXtHW2gz3r5
03kYSFmJJvuRZdf3MGIfgHlMljZEmDoDcSmst22GoDQgF6uZssIzBJFFIMqTixqI
S3No/5O8c5CkjU55KH2oLlwftcpV2huwnoXe3fDnuNEsV2OGlPKQCU9c398JUIWz
Fa4YkPremayA44gIwA2aG+5PPJog8RQ+n2KkIP9qWArl2tgIWjnbpYQN5D3Srfsv
YZ32Z1c5DJdTB26GV4ELpvHdzIannT68fXSlvbkzbW5rZZyn0EaeWM/PB0yOSKdD
g0IJz9DBJsNfh/3pkzLe37dEFQ0vsvmx2ZetCLq/jHZ/bIX8b3wt6KJrfLPZkel1
YIF3piTsfvPxSbBT1WZS3nESklh2Wh7Fy8YF1dgSahv0WViq9MlxQOu9CENpHO3i
z41bWGQEjWhQTim3OU9e8eEf2xAx5xQtWaLnjvStBchK9YEOA9BElYyLwW4YelFk
SaY2ezupn0ZjLjL9uNGKaM3D5+xR4f4NxcIock9sQyy6gJ4aCLOkGAfuwe+fyyTm
B+nm5okKtbjCxESBTJoq3rnJUmMAa72+CkXPsYqRq8O6/WLUqHPt0wiPOVeraeyR
qfaVhU/DIwi48uErBNWeNyj45j+JoYlr2FUSrBbk2s7/FYMNqXn3Xtolovlkv7pH
0sjZYiVz1AzffrQBpfp8WboKBETvCiprkxL3XdwYBmEHFc7VYNh+Oxu+/Fflp1Js
ENhuRUB7JEMXX/wZY4N6yuzP+IptEe6SrJV0JagfrQ6kT9OBdDI/EjdHO2mdoRxL
q3DpExkH+WDFwhGR0IlqzAc8YZx3L1/0rVEq1Sc5C+awHznF8GuTzqLDb0S+Pj+v
l06CWLJ4+DvngfUgnPixnYs+ssIveBIYFC+Ymq9ZvolAmbhvukgUisTJhW+W7/XZ
cwo3wxja0tILuWv01hrWmWcGEnFHqXmzJKaRGNymYXTIjctRu3ltDMWCNiCHq6wr
xURwgDMKdNkqqpwKgFPPH3EVkfcB9BO6Uv+a2JTKwhZJ9tq5Sy4S95K1Ee2fR497
HakvH3qFfi1HajVhdkV8dRc2XwDfhOa34v1Kwd+Axqdj5LvGkkbHIMEr/OfooUPv
ip8+/2QBgjgo1AvnuhyJRZdKxQBIHEeskktR/6vmSbgjggSrzvNLLWH/dHebvjdV
K8ByAUCkDw2FQyIX5PoqCIVStYsg7KwvYV0TcCxLH5c/Ox1mPppHhy1lXwYhQJKR
MT3KfXtGzzFaDCpfFu+qbWg2lrmOvGAR10QMOJ72ii1F+quiJIyFyn7NIkZwIQ2b
hvmkebfaO7e5R/tjAmkQJgKld6K/PPcakg94p4PsL3KOrKKN+f4eGSnG0OsBksRj
B0GZV9MJfBUV/DfLNICykWwvEPqnskEQKL+qQP4WBXo5CKEyeqlbsat6zxJMvGcH
OnpRjm/MxLpj0nPnjLXz5EjGsir13mjEhrnQRkPQ7zoRQlK9bTsxuiNRaMESyx87
vvfaYE2wSiaZmHR71JB9YtT4muH5yxOgGqWfiBYHQeCKxunpDGTIdWjgpRLiQ9VA
nlwhtvRMknNDXq8XTTER/ahV9K2Dw1a5fYHGuKMQeS4mflNnj+QR1EsDevQNpK51
e+RFKNDX/NiQZXNw/EmLBDMoVQXSqPVKkaebkxuen6Qz15wLm7nI7tUvwV7RU3lH
oxpt03AXFSO52p/YDaZlKvdRjlySLQxyENjykdD5sf2OszZV+mBMl3cWd26hF3Pe
I2iNzb8YEK5QVQJN1F/+avUcQk6e6ymda6uIhditr/GH6ZdG/ygVazDQqs9S3rX5
Qnw7Lx9Z/4QjkJeamDANZQ+XJgs9PXHVezkykdZNT1kgORnMTmMdeIsnLeEXXYem
jC6Kremxx6E3IK6RlNl5XCZ108Rl93nsKhoJ+GhMG4AwBC6PAP18bfvnMCeGQqN7
gL4PEIxihCWNEUrCJXq7tzy7AT5AH2FD8dSgJswsgiuFRwrNesunRHiVMRncjhv+
Zw4WF0XGE+uUT6YvBx4S9hOUSQURK5G18YiH3e9Qo0l1xkpWlTx/rn9L8Um5lFqg
o+G31CjUi+SHgJ9FqSosDzt//BWHBs4UEv/qaF/OKLcrZeNTRxycqYyMJtumQ87E
iz2UEgReT8b9RDgoc/eHAKl94CQcz4Sda7CEUKIqTJOiPhnuS5ZzQvVf/0kJ2K+L
H0kGU/m3YH9vLhOnld+eIFu9pj9e88EGQFX2fOO5qJU4/+ucwMeLkw6DoXXnynIf
KFfZ1gfbC+oZjG9O2fSUCmggdpGnhIoF/JpwvuUiv7oWZTirqDIrewHp76z3heRG
3OAx3UQf04LuuxdOx0rt5bYP3UEXjXdgz9xLrINYo177Y2pdDtKbfoQvTBX2/TFk
ZP1AnARBxxyZ2YfGpdqC5DWu6hs5jcLxKOpqF6CDmNbCUHNMtCnOF0uxMM7HLH9h
HHM0zkubVaSU8JzrIJvrfztX00WJ80R9Xd46XOzuCjxBeze5X/FnT0OD8uh1SC+I
lsvnHOv6auMKq3IkrWpERe2nksCRJyXiDbYbRDuu7RNyz2MIwKsXySjAYl6jeaSy
e2wiNe+BBBOjS7Dsw+IdW5HWef4GGrDdqjRPZ6k9nNfer8VwUmZxVbOL30lSiv55
XRVEcKwDciv9g9B9dkQa6rYGQWBRYSXE6ys7BrfqiaGGm2KpPysU2wey3QU1qQ4I
S9LpuHiaAP7flP7bgRdxZO85oB6CeXDVbXCyhY1XDXkTYhuRF0qT6SixdiQEb32I
9xRbvPthOMcN4lji5rfrzkpy7q3U/BaM/UbGhTICvuoM3NNqLaV/f2Y3dzbwU7hk
cU5E+Aa7eBb2VClH8hpqlyGqF8XitIwlV6Cg+MDbw9hsuqioYGV9teOIsfGxLmoc
t/tlFjzBFXqBb5POOPXNI5cWQBkYrWCA8dp39kr9x+AzcRy7HklVhmGG1eqH1qqv
xeLYqnk9dlHkpMPBoexUyODb4BEZFWCEkeyYf1kGZ6y2u0tpiW4oEGOvWNdLYZ44
aBiFG3NwQSGb4wbtiLJS+bXaBwaYayyEA8e0SCHp+d1DZXrdhvQII83M7tVGZfjK
RBxScnlajHEvPaVHRnqbK/a3PF6H8heZuY7QR4g1IaHCaiqn6vdu3eldYUSt6Oy7
q19cI1ZNHMW1fAeRg3FviPRB/SZPjMEwR/o6Jn7281uksZh7y9kMLzx96XRysNyW
dhltNMgEIBOcREibbC/Qv7SjKJUu5OkJCYwsROmQ1I0igQ8ehea1+h6zQwyDVISi
/eIFB+6gdwthMeHokmnNbbTwS7VXpPUsKNv1XUKFxEeYgdwo0/GwEi9CIMltubxw
Sag0jRgdmM10C15ZPUuy6LX+npWaCrcqmBaoWz/kGXo4/G/1STd2Ej01KOGYPa86
86VAZvT7I+Cc8JWRD/9rjzncWsjOmuRokNXM3JjG1tbYzoLqjAQ3KbBQVvoeBWTm
Gt8Vg3+DjeJMAWHt9R9/AnqboiZwkA2k/CvpJpB8OM7iBGCxh6JKnns6+gzsy2ML
q48dlQYMJOA2G/teYgvp5d8SCOesazSZ0y3PHs2e/4VC1gvSc50tf3I+D+Qjlopj
wAyT/NUEEL8BSFd0HQUzns056aBA5B8sHAmftiDQwkV/3RVuKoWFGke+2uZTxiWs
o7ReFXl34WWuPI0Lqob2JXCoHnBn3FbSy3h8aGDC2eSjMMNSyBAMJPMfqITDCvGZ
LSn4gnsHNep5QCi0k8sSOqL7Hrtjkc0iEVZhdmtLcR86hgzOD7dnNfhPiaO9CCQJ
HHifLtXVr3QkOnFJYoGM9wuhn3v2RgXfnyKNa4cFtA+Jjstkj+vt7ySMAI8nLNs3
IWAzuZ/eYbLI3KMwdzcvVPBrJmqjifRlulQqdx+4oDTgphDZI7CHTZjI3+rkUMhs
UkL4P26kUgReb9zCYnAbizUjVYBLoyyeO96bPMxsg9faDp/ghRrbAjPWQFam5v31
LQvJiHgwVhZuRKe088KKKDe/JX0Jnx6oQPGnb/hfWmFp03J4kmSfFwmb0MSYc7nc
6iPy0OOXL6oS58e5i/0AXZ63IteTuGxw99ZQin3mnCywljLBQsUD9Cn7N+abBvth
xelHuNUiSYZwjyLyWyLegyRHu3dqUA4E7eirQoSqMo6U5k2Oee5qOVTfD/LA9U2Y
F7Zr7YF2a+F9hxTw1gxH/cAc6nSLeQOmiOCcIicIvFkskBxECY8kp2uqtlJO2Ekx
RAe5xwEKrqbEfYWeVmCcI1lPXu3jtGpmGGB3/YnvEhzQm0skg1hLSNgpdiZjBHtL
favTqzPgTo06xVwBMOcW4/LMXFCvlp3uOrkKTyqIQlYw/l/G5wcizefMUe03YK4A
Eh3+g9t9jIs1Ob7hSCktrmn15Kof4cJXed9TH4/LhXA0s77oyqBWIWyhRV1lp+If
eCO3FY+0bNNtAzrAKrMCi6L5krwhm37GIA47rKFCua5yp6Fj20natWmFBXpkn745
QBn5OZTkOnmzp67RIQDjl23UoR5Gx7qbjag4st6D7YkEuzv3frhy2W7WKWpximwU
JkocTtCS+5g7vTxIk+sS4xBygalpdUu9ZpVjvMyxBpyEXpoEdUjw79eJeKox4yML
/KDRj4UTbF2Wwhq9QpBFoDVHnBGEqLkjJTJexJKy+qUbVWujJybGe/XVT+WGXUkL
JOt0NqMF8WabumzrtWhsC6+30ItWZihMXjNlYVCU/9aoTJUN+nvihGCOtyqD37dp
xFY3DUJrEJw1m1crU6YRKKbfZBXGH6D5ZPGke9HHUGc75CcwSrm26+f90DwWbkbw
SbVCAElupowQaHTGYSJN0Bi7GFk+m4rLZsxbioNzQcVJ+/Okx9V2VMdnmKgdtlaB
A4opnnUC4toArKaFaPayU0wmo3s5JkEYzz6rkDRFFcYvBTj93N9V2ZO1TRVW3Bed
NeuT93l4M++MUVNw7LlIUc20eZePvsJ2GB46ygOvN+WmoktqMWC1IGaPzo58WUtE
cJlWfQnXOuq6tZhCNybNRt3cFAE7dFMB0NonqS0+5ul1EbgcSkgHt1DfLSb7Fgy7
pTf3O9yYVevaymzrYHV7KW3fKoTaelWvtw4ujo6p2U2vdaN8eBow1FZbkFGLZkNO
ihl7bNml4N1HImsa8j4lUXG42bXkyIoKXDD6587BKW/hRTcfnucX0iC10YqR8bI9
TjEVte/HM/InHstXGqMrH7hAN8P96CPySMEOgSK64bPwO2to5my4I10lZSOnFEbI
PBeJ6iWSHNja6gLSvBH2nkZWHQ7UW/IwPHEmFgQvhk7YdmlNQ5phevsRJLT7P+VJ
CjBPZXHpvvzbKt4Wj/epgWX+v1587Kp+k/JDarllSxoN5L91ccT7gLPay9aK+Qrl
i/xSDgxqBRcQy9K4m+hPEWwJufsi769ouKQ8JDTSxTRN4O/qAW3FbqV9xYQ4NQcF
o5Geu2z+liZrguwtfDy5MhiOfcFBzmHv/y2OuCQ4CXhvaVUKJKxaOhhB5ycKEqRy
O3N/UT5USKtYxTzudclEj8dOmGtM9PGkvjvmSFsXqBc0qEeWRx5j0FFuaxzmYAoW
Lla5VJciM1su0D4n+vBYkLT3gGwCgLyUql5QfRvE8BVk4aS8DENkTUnKG+pOHBQe
Nt1ob3dQzmEYQ2dA8LjqcOBTML3YVqyYDxI5loBk0EuVBkeWIJr+tyzBQ8tkzYAI
b6bbX0ooGCWHgPc8hI/oeJGpPnvIunZUeJQUDazo4K3vTfRcKy8dovWBrN6jWGpG
SrCHwH4AKDvGe8gwvLzCKQiAdc9hnYvX9dAc2kfBmYx/DG69L9BXqABBY8n+ZsEF
2YUk1revP0QQmIcd8tmT7QfqBIKxT3zRBHZ1NTGL2BWqlezJdqPAXU2NwK0ZcGCx
bh0bW1w/TSOGvrU/1Nj/WnQLNsX4ft9MZLO0vgE2CYbcGMGehLAUBw5oretGbeLq
fVoghn6GPZTAVmJqIfxQ2WZKkUDPnqNL1dKluRF2QmsD41F7jeQn085ErM5kKjz9
TktDb2yDykXXDGnhEsEIBbmK0Dy4QdGb/M+8+COw9QzTRH6Fv8W0urUkqUYbwfGf
GU4nClVwTTZABbFhTsn8FNOBVE9HAAF7AVGgzRv/HIX8uVSNOwD4VjFOaIVIazR7
H2EiF5/Vxnap4FD2/kMakXMWDea7npX0hdOYVsia0rSPrsbiN0LgBts7449v+QdG
LWY+AJxkc9OKO/N2BpkGITr3lYa+Q0b7DcYz1+8rEsdIXPD4ngw8B8EGjD+qLW6c
X3icsGObVY7J6NgAB7RTfPa+WKb621H6/NAFXnXPMVWq7XSMg/UbZmhWP3Pufd4W
7XZGfnp71zo3OZW98HJerTe2XsOVxrufZgJQcVJHnY3FUXado7RKKDlz0WVWINTD
kUfx+KpFlq3nlvx37Ukbe+Aa1vhydgMqdBJtfk4VBf1nitYJir16eNDWvIstUKvp
7ac7G+Wxz3LebGliIFuY7ifOKVYOFVJUFay1VORXDWtcwes192DVOP3GHjQOfhG7
CfjK5jjOkJcAuuPBqTRRBG2IrxCSgr53O9+zE0f+K5bnNAfg9gfGrY/oHJL8RmfT
nZ1FO57XWJQiARRymROCsU68CCyhhc6VInGd0l6/XwXeUZPh4NDacLSG5yINCKJQ
4lpuHeohFtOU466WwuKetYquWsl2uxIZgbbR8zuG3lz7rERXLZPOpNSQ9MIi2tG5
IUOtMxwFkzxn/1BkeAuOuE4Ae9t4vocoR0ks9qFIbG6HKy7vZY4xFzp16pzSE8t2
2AbiG+V+TzPfW4l828xfpQwndpMtMQ8kGLd3uJKLezRvaD+CskYoaW/Iwcss+LsU
EqFcEwlYtsjliM7JDNMXX4Trk0TTCb0+4jN/USY3uAPCgMVjp5Arilx+PUmQ+k/+
YoMGd59cT6Fzz4+WDXwsV4Abm64u/kxLoHj34We8m77Y0xrOaRqdCMgQLbEGdfVR
oF/JqbGk9iuXltYWxZQGWnPC04muT0PxwlSpeGVvvyAAvzW1qaBPwAFtUVVw/PLc
SXVa1rB0KSsN6IMVtYslgsbMG/yiWRFzQrdk4t0OzCtsFwNETLRPqbBlUjnwb0XD
/8ptVPexJBhDP+kgdpoVu36P5I/icRpW2gboM1dOYTW45RiI3bI4FQmfPNNtTWEN
wb7+tpSQHfGb0kYIK9B7ZBZQk01w2dO69UWqdR4Ae4fWvGPrweitcm2lYkOaDJ+p
q18jKhEoIhCEsJhhfHEmyu5EaFS7R5fiXaw6wjebrIQ67SmZxBxWTCEato21mAmC
3dOw9gsWVPCb+wYfP84o42J9OM90jcAkG+4lt7fRHe+yK/deiw1NwgFeMuPmPyGI
kY2ayYcS6FT6hyl2u5gPbpCLf9A8UCf6zjxqqI7cJMCKFuEVxM0JuS5ZZ0KiZQyy
bCi2Bw9NM+QAj2/lEjn5NUNXStZlGcgTnD/BvsARdQzfD5TDl5D3t0toZCE0LZ34
J82i5Ph3Rq04gjrLzVfi2OlSww08xCZnGOmD4lIkSqFQfnsWpX7AiQy1C6ozAQpu
/kRbayhe6yw/GJmdR26EzrnHTtJM+3hbHazf7rCk4ZJtJlyM/uFA1BSoy6C/EPTS
0lhwC/3isJqTDKBHiGPZdMtWN+eodRqkFHp8kMfMHzje0pdQC34Sbe0f2PODxIt5
b6VuCk3Utq6E0i/xU7BhV/oTKOLDUjPX61f7cX2ZSOM/I1itC7R4iiQ9VMyQn/JV
Gohr22J/tu1adGeegxUnYvqGT1HbpllkqprxSvh5vp7ZYDOAsft04HcPBjceC2qZ
i0Ye5AJ5nUD0Gy06mbOykOeRFLXI1oweB4zYVLWYx9OWtZvA9d+ysZUDHBkfuOZF
0HClXq0L3CdL9LNgEkkATPbIu9n2NitBlloymo8GNHXdfG1F65peL2m6P0KS39mR
KFFCeRdeVW1Z/kuXwP+5/aPa4f6vsWaupXGS45LQ93lsiZDKubMtnqWbw4EfdFvE
icckyjnYBze5EKYLImyR+QFRxNkjf/JFfuG0NE1ZoD4jRfG8jSYk8tGG1NjEhQWA
a/vmUjmi53JchA/pQjVR8gcdYgUzzl1tqY/G0SAEG0O57L7eaOmFxtc8LbqMctBf
XR+rUwPAn7+fSKT/1PlKCa7UJwqiCptP7fQ6yXwjuuN/LM57dwtndIQupjiPEsSl
Kb9tsT3AnKMRJZc5K0473V5wx2NpLEcfhOCME2Ad+xOIVRpd06c790W5toQLbe9J
KpAQuLu3TyW92Xvay6lhQ+29tT/FhuV7cVv3QRAaYJ42VOitmcQ3xmoAGmvocqLW
vbVpjeUIn3jRgk2tuPytauyKleVULIiIjBa+Gb78g+tXjllm5Y4RTzSIogzC98x3
CfcmMc17pt99m8PuKATHKADtWqdgj8dVtIi96KhXXZG8DezzCtk/IxM73ZgCFq3h
SH8j0jjUutfwuu90ycJAvDvemsS5jWaWdjsRbF86kihj/YIVl4etS/q3wjOHfkuG
2GquKhJ6VNMi0NFTRnMjI7zEngyeNIJTIA8EdJCvtDjz8+IuvSRH9wAiNOKn+VTL
Lthf/PNKoKDsblFG43YsR+QwfNO1Apt1BWzKXoUmFNH5ihQYys9hIdLSVbJZssnl
Cn0cmCxDj7HZoY2zUA08pDrJA1sLgjyMCcAgsVxdKLiKP/YFD03ot5lO/LpnYFYw
E67JtOCFOA8dF1Iu7YJXb02mRxXhE4rzfb6EreNFAde6bYrh4F5BojzsSLll7qPf
KOMsjxnc++q2BrZi0dxf0vdf+SFtMPR8dB8sTI4nnMKWe3LFnsC3P9/Pv3/vLBSB
s9WVY3a0ijv45KdNRjk88ij4VCmPB9vRBeq/Ru6KBXIzkys+X3E2pz4TQIDuxSHn
Wn65aYxrsgQFdM69UKO9MVc3LvKwp+eSkea4A91bRJNshSH7ltayPLJfOYuqcU/n
+5jNNAyyYYgwxvTeNnvR6+UPUuUkvXQ9xXUv+UdQiukrhkvy/L7dse0FiPuEigmb
oHmKH8/7TP2sGFQFVsqjD/p9z4vyngFtrF1ihvpy5/VRku1eqB5Y8Q02eReA0+J7
dQpDeMIGGnpzOwn7VwMZyiNSDL1qWo4+afaxL/7Oy6y5uXaQOchxfPrZt69VcxCW
ZoFAdbR2KbbUDcQMvEZoAzFjIiT1vmyR8dH2UDIj+KnybGGuNr4hDXy/ZznuVLMz
1zPvBCoSNorE11NkLE2V0L+6xZJoKXaGM2k6LVmt0YfulODNYcWWKZSfKK61JuVJ
mdjN0wiN/hFsyshVwUjamO2c6mefRGe/5JP5rMa9wufFhBJcSULm/b+D0W55+q3F
emTIl2vRzwVHbmigct0cY10kGSPr60QwTaN8VHmAhthDxNaHfRAl0nqCk4itJ9TQ
8VtvDX+qwwWsSgO+YIr84q9mWhqjSIyhfoRd9MoptTVGToDLTI2dI61V/32KrE9R
JbEMZhbCt/K9T4V231V7hhom44IYzV3jWrjNwtJJEcd/H4ONqekd4IYK0Lt4+oyg
IJxdskKxL5q2xVzcGu3TwhLXo96NwnqRdn5CZgX/329RZLMXlKVNhMQUmMqTQmbR
LtsUOYDi65NLmi82jR6IIK0mXEblzEfXrPWim9ncQiivUJhaUUPE1TjG9u2BXvc1
avVwIHCEKIt3Ufa+X+b1KVsUQZUYVtwEKHLE9GTvqHl7bMXAFLuxT/sIQd3JCuau
8NVVPESuFw8Qgkx6eUiw4vhymKBrpnH024e28OodQK1bEZshdgUWasJJsbPQ6t/v
TCbgv46uoj/q1FfADENOdVemiiJCI2rnfGD5Bv9Fu1YocOEEUBEcXkPc9pi9OaUo
NqxaKtlitxsN7fe+GKJ+lj6mVZk9nvb1/HHlbFvBeZPJX9s61uzZ708XSmENZvVB
ZEUBS2xv/08lS3lgoomAsKMYKCT99rALhSKEKNji6K9HKiJ0FjITrbc17id/AQXB
JInxRL/TTwBuuwHX2nLkOfHSpnSMb2T98yeAvJGvFMgohIPQFN2U2e8kUcbqRXZt
3RWcfTIgIt2admTKbpC9V2k+EB/4MDsoLfA3c1C8NK6maHnLuadNOYn5VBKwKyxK
6vekx8ekTvCDjJ0BNC9MiHwQej6nWSFadxIB6HBs74DfWx0VWq0M6UJqCaK2/LWL
OQb/GRTiMMkRWRAz4eKL5PUu9+Xieu73BFIxnRiFwTmsrMzvPzja+U+ospQQXhta
/eZPbQegkUiwvrVPiSRc6v93RD/h63ci+3nH3LyeYVRHtkmGeUPr3VmKstLj32Vr
MV9AJYQySUWYd+KwfsuVpoV7psFi9cTP+ewLIk7VarcLEztaFqld75Rxxj+iSK8t
AOTGRlNiFvy0xmcEwP1ehONqNr7hNG0gB2xK/49Zh7XjhrRcZyLJ0/jwSumDYDkA
9NVKYY1cWIQxSkkykl3nYFzqzN1RolAupEvsNwXjQ0SRN7qbIyyQH3BG4tV+LsDZ
eFItu2O/cF8+DuaF1YgYxPU9oK5X582TPUHH6oln/rzbw4YogMIm5p+u2xaSN8gV
DyrYjgbDsf7NFGqUzKijLGGpDbvY3uY9zpKEi1gMzMt5bdmQLbpqCI0eHE7Z1/Am
cFrLMLoCgWudCTlQZK+wYlRNPDSm4he1F6Jhgw0e2L5NbJXq1tUJBAEfi7LzWoDZ
NcPJEJRSm34xnYQKmSoPN126O8fGCFg55QU4ENBGbwaqSfLoJc7cTgiNxVSTujTJ
RQXreOCGPo9wWIBQdqIYazucg9M2UibFOdP/I97xchZUDhk9S5Y54Wt+6jTlpphJ
c0CqoWdbiGSPt/RMD/WplZ3K/oeN2QzaiwCo/9WgjJiYpGqQVvK7eqhlFyAtgXBv
/j26715LDpcclgGerB2ATTIpL7bg432XjuUeJicI6An2CuQMk7SEOnogK3OBHIbx
V6h4F2uIdWqtCv9xfiBNsuKJZptBwsWiB9lJRtq9sSqxlgAKzB1npWU9kaeUjlan
2LcB1MYJPCFjrmTUxajpvDN+qJuKQQ9NfLeDASiBpvB2nGXm1Fgre8X+kuulIwPh
EehHu9E6XS2VP6R5HTYjukESa2qQDDyJ+7sDZigwcgHafrrMonY07jpYmKkpDHKC
rLmPByiqEeHO5lHvJNWNLYh3tyOKnyd6rQnxNZVFHk6nzZrEYLw6J1z5nnWTb6b1
x3+JcNBwy1srHUK6tNey466hPEyGYa6+zYMTowhmnt51SMwOohjp++wOApRd0s9U
KjHuxxnO1Yo9V4JjjLhP5UXtvc2ffmcGp8prgc12MebQ5taqnQW3DTWJkUiSX3+6
+ScGgcBUPsdweNxW9sLmxUt0t8B3PChx0EcdXIl7oj47IykYT2VQCA97LrCm2PLD
sp1KUZh6IsrfFcGA/xdD95n4ORMBxEFQM6Ma76KbhArMaWXRkXV56ouyeOtH08bi
zznbpUuhXhKiGEtjfOtEZ9J7clHYK3IClZN4iJKl94ZuPydnZMQvhaz22Ynk8eje
m833hG2X38r5s2FQXN7eM+kGfCnDZTIR8EZEq26ryi1mPI2jvR4CalkYJn/s/BYj
46VbhKkWEMGsJwqnczl3b5vEWVUE3+JR2vxJwHZbH3YiRMFZ6SnLmzRWOEEimvCt
63CEGoJW/vVKqhSW1ldAPqdwmu3VwBHFrRvRUFKemLt7V2pea8k3v6JWYHYC70Cm
TerqwGRFUYJGaC8au8cLg/gHFf0an3OBZynk0syH5C3Qed3KnTwulyuV4piKfBDn
U+lRDO6kkmZv4QRoP8FjfKoWy/jIVi61IsZ1cOxvh0VLLoim+/z4WYlgqIxBFY32
sC+NcTXicvejXJ74m8tBOIEoRFsrqbxOwyRp3goa6KiN4JyX11FlVcYaB61YzJZq
BGebDDWpx/IN5R+5YVE/IunH+iFcIszY/7b4Y/hmWXrqesaFeiEoUp/Qag1bjp48
NWuK61Iv1FOjFT+otAj9GHwlFOM5txXJgvRRHv27NwUHWr/8QxxSNh5OpnagU0v4
icbXJQFsQgwpdG8zLTwo721UjzjssniRjjfdrA+9fjq3baEjaTg07KewgdtEGMs8
/vu/SHHYwaGklo8MjEeSqv58V9HwvgVK/RjaCIjS+/Ap74GFLer0f3YCoHbUcjFq
w2YSVsLaYk94geWQ13xM2yrIrlapcXLZeNCkQSSfcuwv8qrb0KaR3h4rhPpmH7G5
C6qBmBHdqKamcSp6kLmK5hzt6fmWo501a654fhTQnmAYBaQma3Fvhcv//KKuX6SD
8v8+0IGw5KnCJGwR51K/S01pIPhBi0CPYOauRicAXTSclxb6qX3QI7hkv2Sp7lwf
jwz5vjXT3B2JIUOPN2HdoAkw0nvez1CBgSia4pUQ3HQdBQrgYFRvrYytbBmoy/jl
EzOYZ+YThMgDwKtI7zk0r3eQV8QLhHIxAi4ZnxiJAsDo1sr8T6vn4AVE+/iN54B9
Iw0oyV1I8+4/mSyyZwG8KKVbytON0ttPN6xJqA0IBVPWeSMBz76fX5173JMaQAB1
uEU19rzPLGRYINjrBWUpvjVJ+RnLxg2Nq7TjVPRx9lzeRET8sha9G3/o7sM/MV+K
UwY9UYKxj/Ni1/O6eSuK5Yc7H8HB9w937FRlIxbU+zQKqSgytc/ths2odu7i/mnB
1/Rai4DmwndjyX576g+ngWhac41/WN1pNrLJqj2ToIHsoAnvdjkzmjhtfDVspO4A
9HU1jTtogopDIjr98OQed9qEPyDhUOrdsf8Bny4M7vEvZv9/PNyUzx1VrkscAFeX
jcatA39Fwfq0cWFeOVB/eHwUawQ6pV66zlQP5j8l0oOc1jAgc90V6MOJ83YOJFA5
rW0Y9iQryEQv9sORKPtIlEeN/Er00aWZBLUyfeplnpnbUJs0ElhhWaTxKws6Vfl5
R13RBaE2CcXOTZW1dY4or9e4ig8BhaHnfn+TBhvERYP2ZwR/Cpra9bfLnyVr0v5j
IN4v3IvZJ2KR6kb81hGctcrnqqrHI8/K2v8oG6TsEGpjICf5JmKKmqx7QT/VImUo
IgRU9VIio1slm9LHuy9+XqzOPUnoopC/xOaZ3zDCDmmdgKBNAV9LdMUZGhcIl1Sr
dCs283xTjVfjZUqFuUspuCueNJfI5RIeoloE2KrEwfI05mxXagV62JLgYX/Ra2jn
8B+PUEMuJVV0pTc7jMrhBLP0NF6I/veFytDubputb3ptFOlgL2Wf35Sso5yEYZsE
GD2Im6l35jWRzdz6YhFgBVp/1yQt/vBJ2L/uKJXClYfr3s2168WOHOjbk9Jv6zo2
6Tr+dqTCPDf+Mt70wyhFgb6IE9JafWqNjs6D0kpSE7AdlisiapVDU8VHtGI+j0ee
9y/+82zHBzCjtlbr3Ih1FXrGWgPJ/uGFTjMPiajZ2J1+W14jtyrcOP9h7jceQneD
ZLiyng3xsuY32QKHKKEigEHaxwdK/TzIgjDIPMLWtq/a9PMH+r8wM7YirWY7W2Uy
EeDs3RIyGmrqz6p+O804N/tM+FbTgc55q25Cj4/3yencYYF/J3J+D2HdsXEuil57
JT+9SjyujEWDpVWAKRcW76PrQOBUuDj0bmeXasmjBy30Rb6V3rPpl3VBVZ8jmWcK
5dEPyxXfFu0rMvqwQUpupwkA69NoFP2pLQ2pqK7SeWcFfi4KKgPzJNfAbgk/3Jrm
7hSbSuB5lgHSske58ji5XlKJYRGaDwLXs/U73mjswMoreFkgUz5Ej75Un4mKIA+h
qm65kLaVTbO8mPM3vI85ACCWaaANWr3TFTOVSDeY7jJtgAn4f0EvJCEFGR/vsQD+
Pw2Fde+ungNBf64EZchMQgHlfMlFtFY8B6vFdPbkb4pHuepevQ68XFTOPZV/HJtI
M7QF9/cKBJYgW8PwtEab+u8wO1GoKv9PANnsyTiQRia4M2tRVmA0DRDBCNTwnyT8
KfvaoL88QHrdU/wwCphFQ0sQ4lbP2yhdLXAfyGrHNj9kULv3Acgk+qx62tpLwr6B
YSDtwqV3pEBSHy/fjHaB09hwPkSh2bn/hGeERamyn4umSAZLwYw9p/KFNhcKC/LX
pKUK0/ezxVI+ctlz4bHaHSr8oL3NDnztVqAYGLothDRKF1IBA/QIwMjB8n4IlSza
yDP0wYWn3WX4PQrEpVR3gbr01ZTu5NTLr9U5Lnu85TSgi0uwDiLBdLXkV2LqbJ6e
iaMjcvpMN4OclqoIAGe/cpbXXfTHGEvzYcYZir191UtNJvmIlCtAh+rKO5p/9Xyn
+I0vow6AXINu7c/JhaRq94rfeEy8eR2K1NOTpnLKHVf9HU0RL1rmzRW8C5itp3yT
6J3iPIYTEXbcS3FZynKCWrzWUxZniJV70G1o5+HJvIZTntltuMdrmlhGvhW9Jv6n
6x3WKfCaQuXVc6W8GYtR3WoQNytE4JyqdLdswAsVmGrHPLlEBvDsdXrpJ36sEmp/
4JyuA1gATXqt2f2+JAN8camvkZEOWp5TBv8aRa9sIWvjjAr1UuKgwiLRxJ02EjW3
CZhHFVToaLstd2SJxDg4pBiFCGSwmUG7F9tvbCO3WXWsaTgp4CnkbtMZRM6co0QS
CDgJM2YU89dLnNbpixA7GTd0ve5bdLlEpYWHXEE9RX0q25w5tP3d/yz6/+LISg4w
RAk6QLWSG4pQGwf2qGaw9j4gJXX44cOCXU/naEy977QU+Wh7mCjAby7OAJ6Vltym
GlqvSx5y61ey1o1euRSiqEIxGVjQQAZP+TSemRqJ9hpCsSG3d5hO/rngoeDd+twU
ntIRU0qL4X3mAs1ioMxpNorHYkvarupvRdlK656Xd5klkySGUoTotsMGlb+Dcfgs
r4rxHK4RX5XvkHefxFEN4FWRiv1jVJ+C4BNUyg40DqMnBzXlvc9iscBg3eM2U6Gl
lawY3yqsRIbVTnu+VQv08Aac7l9O/1Qr8RvWgBg4oaDW3DDP92wVo7qDXw45iTMq
/zKatBYydDSjYaRv/9diKIbSCRR5R/xhe92dKqmrePNRO1LDPU6KpsrZt6/ndT5k
Qlu7BL+rNJDuPIoDoTmaQDXq4gdN2hg63TTczl0D3pwOyUO9lALPL0AwwRVZEJHr
nzLxdsObWrt/OtVgsGIsfkZE063650uMnZ0pEdhOZu8Zr+v2u+E72Xrs7y+yFHQy
5bapBkAlFVCsbdeNlcpeA7HyXuxd0ohIc6kzxtuLcUMtNuLe+RWE7K6O13pkyhLK
mZSP2EamLt+14KnnjkO7CmsaSwWcKjqbE+vMe++CYTfHuZno87qoprBqWCmKlQEX
TYYEgBbZeHJzDc+1hksb1uGiHPvknH/qPGFMkxNOPU/Qdt6CWyC4Zg/2vhWJ3ufz
zLq1v05JeY85nMLfLE4/oP6nFSjVrq18wHmuBrE603WMf7MUllKtFVjuV0oyyshk
YS3Vvk+iRv2aaDu4A7LHQtC/Dlq8o4Kpe9ZQHNl2YP7wHmRhOGSJE9wnBJuPMzIO
LCCUQ9gFxczU7u0CsGjKL0uguF0ZjWPIIspu25FFli1O7EXHQKTokD/Bcc7GpOXc
gdXniKWS6ASGt9Os04K4NLlghD+37yfZnxjfZnDM/FDVqUafNzTwCkd8EnGzF3vT
WSw0W/MO72utCLZoT3EgIS/aWqB79nzsyrhWof3SRmvTh5C9AzQ+eQ2zAflX6AW8
F+5I+Z/F0wqtCHrpUsaDH6OSHYKKJb+o8sfF2+bwHvqrwEGCxhZ+wiQjtXAA9oyC
HA6VLV7zBXUFlGaEVUsgePKqrWBjVrCZckeg/hcSNDYOOUrlWdPg6+GPfnYyu864
1V//D82ZjnD5CR8F4bKRSCHxx37uk1PF5bE1ouFgzWKagvExGVj8OzNRY5ND8G9j
dZsZkf1YAskpzEXr5ds7kW42mLrxng/5r4P1X4dOulBoOyzgelQlmnG1RmCLm301
kFbjVsn0a0slpcxwKAlbj/ZeIqAAVQEpJe2LBtn0hwA=
`protect END_PROTECTED
