`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAfRUd+HgalWFgOGXqg1qhPm9kU8fATJv6/yGt1x/4VE
oX3zlA6ftGn0wKoB3cWno7kck7p8oRU4h/FrnvnR1yrKMiAeRsgFwKYmoJyF7adG
1CwsOO2Vm5YNBMaxX+WZHpcLj/5qa11o4yX//+U5Ngc7A9lLh0zDilR7ZLxzvCm2
k9OmmH79UdCCno3sZQ4U2z6ASpan/X7fYPvRofRqrMiQjb9XUcJA9QyO1jcqAdTs
uc6VBiHMEuJoGaKbmWMIjQ==
`protect END_PROTECTED
