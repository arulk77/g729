`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJziM3rFT1Uui9rstb88XzRBDcCKPiU888ZV/7UupoIh
BEvb2knwxZ7WPFXH+wyAkOjySRgZFvqUKQqvbOHQPFQ3yIGEuyct0WgFBZNE/aEh
oDA1s7qoFJcjfpcYZ5U8zVNY67NHxuJhAPn2+zTnORgrK3bYloaeWtlXJ89i7hxx
QgZp+48WoeY/gQEtwYIFR8Mo/eokIAQr//hsQFOnuRQreALGa+j9OuLKI0iDbYol
gKxqtH6obAC7i18vt5toxnJWNmMxErz39pS2HthF+Pzb2JpfgZiP/xiPCsJdUaL6
m5ZbC8/n/jTqbr25iXioTgTg7CXAZG04oHPMhtGVvvz3/FR7HXgC0p8IkcnN80Kg
nOq3uTM2fzoVPXqAyqJTsYyfg3tJg4zzgBWx59fV/d+81sffNpyvmP/GmaM2Re8z
usHS0p6XmkWsH5KoML4eB31ji8Un5iJ600yeuvzwvFx/4vuJqryl+0laO7ByCAHm
VPfD9PZuBdgxWq8qjyirf3iUqGuUu0b95p5EM4dY6Syhqn163uXXPq3iTWTJcdQu
A+48QLq65pSbWMvMG0ptfwYp8sES0WhjyMeRU886LfOzWOecwpzAhYlbjdo0tdV3
YitJZwuzrlA/F7cTAiBpY3zKhhuASjZphd2QQXcXmZnx2+DX2PnrAbpxFSnQqWS4
Uh6fsmqF8cuQHpbk/axErWOUpmqIWaHtewYuJJsq2Y/T98+D9aTg11k7ratnwKXp
pAOUhd6aF9LzKEVNStR/4eIzSS5Wp/qJnpr4J6AYQhbyt+H4AcJCAXzUhOM+uWkM
sD6fWfJXCDNbuUr5ioWlSOT+J2f3ckR0xWayp4Gy4gY=
`protect END_PROTECTED
