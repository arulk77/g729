`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHzBNbk/BZDictepjHRr2UGrkhLV8wg4e4C7IhFMtmXP
cWBtWVael1xPx5fKwBylMiHsEy0ZG4o8EOA0DTWHdO1cC9vjVAMwOyShAT+ZQWBu
sD2QXcaww7Yq9nnTvem9EK4mawIUuVCZ9o8E3IFBmPwYBBM5fkw81QzXoZJFdVrv
nokO6m6udrC5bF3dzgMQsMoHzliT/vSIcl/T9DUrFBf8dIuPhBl2rTQ7rPygnkMc
ITW/KErKLsPir4y+Q/5ORHzrPT71BIZAKfwG/XriXstuxIxHkx8B5YfPmYBi1sDY
spsKSRU8efXctbpIM/qJep6u6Kt3m6tbpufjbVBerusvh3mK+6XdBeX4H1hoN4xR
ItBi9g2pzleLcQILKMcK9Q==
`protect END_PROTECTED
