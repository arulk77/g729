`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
NIA4ECqsxOGKHi7R+TPmMgHPq+afvlrGHEiVJeUmLRNy1HVvQVeyLwGhYbHs8/ZD
eFhcuaF7B9JRCGa2b0Qnua45kU46ncRlTU+DWddPOS5sG/2qj5Ub6bLNLC4AFrZ8
TB+gPttt5EBcIfi9Ww4YeTIqkdP5/p653I6NjWp0HY/k3VuBr11ocUpwv5nHCKpt
zo7TqdKr12VK0JWJJTfiC9GHa3vJlvrtZXk1taERrmX+9bZWADUAYBEDvsOFaAi2
lmG1Ck9kL7wpJZ3lHV7R/lYfQveTnHbBpqLf5W6MT+MQD6CkErs2frTXuxf+IY2/
g8Wew9nZbfZU/UVXvc1lBpvuF6ClVMnrN0L61V7cUnyARNehz10ybJbAxa+/M0lh
XbvDWsb1r63QGmmkGgRwAa5Dek4KsS9Qlgncc8FdCI8kpvLJK04g5EqQLczAfeMR
fuA7PqzfBmu3vur+EBNs8vajVGKiC3DynfdDbOl/c/tRwtod8UcaaKzTlAK52DF7
7CXQNRp1towyDVKkP0CngM8PlkPag+Ax22cyEhHkZifvWOrLw0hk8AR2/as328m7
GOX20uMnJQrKqp5eISGtl3+KuoC3wZ23MSgmbqOXQVc=
`protect END_PROTECTED
