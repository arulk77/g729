`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD6DMq0Vw3/Urfu7/0ynSNSSL6OxzP7SYJ0TO8ncrqsG
S6XZPsA2RjezR065vkvMSpRxt51l1krPApLB0kaP38UpAeBeRHe6c427R2f81slz
0Xllbj2KAsuTx8ZgV051VJOgYjjN35J9vuxpOC3Vl7JkU/CG+FivvQ15gdVJr0MY
n+a9+5fAkEbYUdSd1nggLx6dWwNvxGMDr3IzJ2UfiVW/LvQ793RLUb2Avfn7sZ71
7DwjYtQUxVH3KbSuApL1da3ECxdZaFkPdx4ZX31n5MxJrYwPgqFeFlHB46d01VEP
UacfDVz3DVoL6QF2B1yCiKWw1Yxtw4HV2Cg2n2+iGJBsAsRUHhBXR9n4jrR7o7sP
`protect END_PROTECTED
