`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41+IJum+IYqwnPRq7qY3V6xH9sv6vIgHEZwi9f2AyujG
UrnKNQLN9kssvWRgi3i3w8ziIfv4eeSBPFQ6falUN6kjCWWP3Af1Tu2C6n5Lcvww
guvCp2eaiSmsSLCtsNYm+q4uIQizBqfwMpEepJ4I0SlP8cAjtxPdizVTHFndk+cZ
mpqFB90uCWjOhLuQFVVt/vl+OEOYgZfITZs6okDAcaMd7H4iZQTdKq8cQzCzavMw
7kmTVyi/g3SQ8ZTBP4o46JvRosRLUOqibyhJ735y2axwMv5gK9sXiQVZHaUsStg/
j1ycue5TiubOpkkhpnALYjozlmkIQPbe+ql5k4m7J/NZ/uIezJkhKak5iUDYeUzw
FzIN0n5uqjSHt9atmzoGKQ==
`protect END_PROTECTED
