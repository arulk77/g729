`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aQzz0UXd4+vrEscJVE491MQUJE/dXItYTbsnknTpAxKg
r0DBUwaAbRKTr3Fss3iQrgvcihvBYt5wm31ZbWM/U62HnYr+Oq5pMVDG7LhObulf
ARThhslMuGDJZ8gdD/f/POFS8CRUYItZWNvKYoZreVXPwqZEW2hel3ivbrSKux90
Wf3I5/udMCJ1NVEU7x21G4LN66WbhqWnohrNQCNfM9Hvk/CgZFEWiBiRP34rPh+b
ikS0v2nIa/OmS0biqcax+nssEJ2r0uAK06uj38F+LAq/lOo4Upx34IlDt7nEIAQz
xsCjpoHVyyxIxCYv+VS8AcLWroIxzOYCZzsctordAg62SkKUe8z7O7M6navVaRvc
KnonafZqGRaPrG0rfyHJNOBQgAL9CanrN2N4hRyFeK0iIwR2GMeDK97YzHzOdXu2
8wXMzPpVBRug/d0TRqZ3QUHOsuh0QKKE++X6henrTAEOl52pz9kg+fHEE4UkFYqd
6Eh4XZlEe2frLawvTdJUuXIB1FrDcrgd5R70BymlDy7DciQTvB017WwJ8pSNtTKG
SGLeEAzFu8cmRh+qkZPQbMhViF8N48tln4Q60dWGKVeDBwVTc16qtO8h4yD/gYPt
OSigMa9vtGxBiWElkfao6K9IOD5DmRqE6Cbh3aKvfYpzhMIMDsuI6VugUWNzgaSg
dVX3GxdLxRIq8Xkf3omun9ZM0GKOEHwsFaGG5j82idSHKq5af4sxb+IQkVhbtznk
l/5On+AqTRoZJYwFe2hBqcZvNwn8/SDRvCkGtnTJftEzGIYYrGXYeNoAE920TUX8
Lo5ymqaB9ZbX2fe7ofVq0uFFH/cEL7DZJL+w2/m7kwZdTSO22Hy86978Ny+NEJ8N
XNGBYDxlDSWTVBRuTTP4EV/iWV9JiMI2JcIzRmJEWqLxvPniE+DJcM7Sh9de6r/h
T8UgsNJ79CdBW8od45RnMhglpaIrk9hwhr2KZ0a9BA1/W2+XgpVfA3BBMWKMjk+9
41k2DEA8lW8PoYgFWUL0lGBe2+h3Qj2Hjo5bXojWhd0MAWiQGqSTrWh9WQawbcP5
57yNXt8Qj8GMkL5RpaUaGH97bx8jm0RE8Jq6J+nUavOWUTB5JUb+P7QofY9MASo5
kftLdwTGdW9wQSuastlHY10cINfpLqQUGybszD2DKCRzXxDIUcVYG85Jc3RHpYWZ
2dBKvOcP9JSsVKKdexVEgCxbvR7MQzj79ALfaOJuP4gMxXqxnfL/Ks4Zi7TBYVIF
POPAlPW0gooyDTptk4RzvITaVoNIlqhNWwPMzegqr3/IxVYbx/PpkA9NRuvnXQiK
k+cWKMvjrRtMdkQvsBklNqBPqWEJzBG8H0K0SKS6zHd/v3jPKbRSxdIHr6t7pZ0f
CrI+uvIAb46cBW3AgMKdnDrN0DpqQOi/ffHjeI1yRmB5gqZ84EW8gxDaov3PPJ0T
OC87PzQwCfmkCzEQXLXo00cQPXmgBGqDpswgLeq4ghynxafAKXeFnbo/nAReI2z3
8tsTXVl4Y6CKTrMF+kvKC9Fn2vIpxQvmyVW9ZRCg1N5jiLydLmnZIecs8Kv1xeoZ
4SBc0DNnevTODklRmB5PF4C76MBOJWRtxSLb1nq43gimmEpO0FbR5ElBr2ki5BCe
aSKYUgFTc31aSOYskPVX9iDHxligrAk7TmFIL5YnFZMIpbHPJgVb/eG8hJn3S8k7
FTeofhNcVBlmDq6MAfn/kCRpuk/P5ylQSyBkEE5Pmu6bpwyC4STTvTcExrYkuGXG
dzjUNsbZ9uRoh0jdFp895YSy/YGHKAbuRC9Jq94F96Tg6CEo3qSisfymAQjHwKoa
WzM8JmtEPQNJ5ALve5DswLLsgVLiw3W/edsggKz4HcY2x4bjZt7zpwmhkbFr8ESb
UtAKyyqmCqJK6tLYXbcdfAdtjvw/QyaJHvXGYNXaXCNZVy+lEqdZVJ/CkD0WeUkK
4qj2yZPxe+8/1F9TDiwzrRVEZ8efmYIBk81kRUvMYBpgq2U/Sy85UQcEPdS9ica4
yi36KkrEep8HG9xAmhcW4pOiljhg6YraWrjzEjWHxYlZg8Yx5XtQgTqVamOsD5g5
OUURzSYsF1TkL47P46z8DNlCBrS0csCFklzGUKYDSadRf4unlThspQ/bXp8511ch
SnI6pzCcvHqWfhuQFHS/9M3fxFx+gP3inGL4HSEj8M3ldlBXEFI9mCMm4JAV7BgF
LwmgTcTSTi3/A0cznPy7666+rXhQSvCPzHeoQbkH8L+wRJd8Djnhnwg+mw7qCFEB
vyCtC6HQDx5DhYMltw6/JA1X74GuWLAV0mmLNe5jOjA=
`protect END_PROTECTED
