`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGV811bll/Z92EmfTIBRbZfJVlV9+NWiZyz7uSHFzpjF
yltK4Va9jAVeZa6CdgbyPQQseg5DdPJAyV5IRwbFYZAeJOdq57WKgln6eIY2Mfe2
LMsjArzJVMW9ZPstHGSNu9jgSFuw501s/7Mi6gFt6Dj6oCP7u6Ec+/r5ZzjDtvuE
Lk/urT+jBOfuRgjqWVPn4wV5J0zowcyfoqT5l1QUW9G9aAJVTCfRnuk+ppVhEfeB
uC4Q09LkRduwExIkqE9gsj6CqXjAliTgECiEEltatPdgk3Fc5q7+WHIKxno7QsU9
d9RmML4PcjKfUznWxo5eIgNib1SlnlFv+9UT18cbRVZuVKU4AJc90dnf+KjX/LU+
`protect END_PROTECTED
