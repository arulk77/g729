`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAsh1P7xL0EtcYlyvopEawgMAOeW2k3/pjbNPHxjYGwM
lLzeFQW8O2LLySzVQeZP35Ikxaj4lC0Gy+zzrUjjGqUh/YGFSgJT2EpWl8JTsMVt
ptXwHBm+WjdyLZ1Ne+l75iHflWjBs4Q5jis++hGW2bRdmTtspfokMvQV5+W9Gjtx
P743/qC3dHo9LaHBdg5aE/eEbSc2Ibs0Imo+ngVEX5zH48qLhdcIFun1bPMKItaf
LWnrSjbvypJ6r0Bh5yJqR+KEmyehjSOaeaoZy9m5FO7tYY/amL3R6kOYLXsjTl7A
P+OJ/K8BTit8kx/J/PnEjXn0296DHpGjqDCC6tXbWbraWP8VVo5fJ8C1J+5/Esl8
lsKJt3Tz2fXFheHI90XSp13OzYLoDXx04Wagpxif0kl8RoWtX3SPPEqFdVXOTePp
ONmvTCRBa0ZsAT/2UfzYEAk9gMprtCv0rgQXgLJ/sg8teT+KxZUJ0RRmVvqi/E5e
HL7NBz0oYn6a+OMZ0X2j/MK7vRnE6l5DWhQSjoqyaYThwxUuaR+F10sNDub+e8Lt
`protect END_PROTECTED
