`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zO9Z4bBvCoEFGiSUl6l1MRlGahs7FY23jrAhc55eUee
gXdtghmHVy4tqaqweQiUKQi43f8gFQJth/eCH8rPrmko48dErUhlQUcALnAggMok
9pdo2HxoFk9JzqIlqjRq1E+lXMl2LfRDuqzTvLt2K8/4g7jdOK68/DpwPatNGGgV
U02lwst28MOVwWb5x2loUdp90lJ1tLaEYZkca0pXlLAezQvkwG6efGmLr+FG3lyH
wRoQnSIYF1tRyopWbI/fMUGHH1frg6Di+A3wYUVLL4nlGMWkWJs3Q+hEP20n4v4Q
kuuyloZYH2MeF9Ueb3wnUA==
`protect END_PROTECTED
