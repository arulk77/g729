`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEFF5cYpwspIkPWmJeD1WDwyPNQVdFN3sGMGBFdBFN82
NSdbNpXovqiszSj9csK/tWp1dDT5TsigYC+6Yjkvccdbk2MDWx8Y0cWXJ5KNpbhJ
8gii74L3GHAjspF+FBEwsiYCbsZhtMOeErgMwXNOLwxfexXMOfB2IS7WS09Gjei0
z5/ri0pNZbUePCMtS10x6tbVARy4TbVvfvnFbMDEx/ju4Nmxy0s4XGttTDYf9Ucf
L7Z+fhmWuaxAiHOm1Y0P1hxmJOSKIFBiZT59V/gHpNeEEeD3XPqE4af/VjnrP7BF
7BP8EuIHVAPRJk1EO2lOWNsINNQ0b0prPkb1cUMRs7uMqaPvJWqceBHS4tNILEV/
T0WmQz4ugsaKFZ+yvpT8AzSaERym65thpstFj+RDAhZok7zQ9yJ8KTVAXcry6BT4
g4hzXMgw2VoD+UMHK6jEvJcye4QMI8Qb0RrXH0hShcYAJgA4rnWyKxOd3FAHIxb6
0VMSDG3uKPhgguFiPpM1Fkakh5SephF23jnh20Xa/P2vwGFjS2HUFP63RvdcDmrs
RGOj+n+RQOanxIaflgW3AAC6uNK7j2+Ds7XfP/ikVuYdT8szfldnRuLWXO5PkvLM
U6v+hPUUwN2rHAdME8dP+Qe1Yin6/ASLzCsICn5Q8+OOzfQM0ys32zxKdlhk2QVe
Buudm4WSNPyP328z4JyFsDPvh8AuqLzVniOAmA+9Upu8/UUg+3MXCek974ecdEaF
usM7OtPbBJDAq0DS4OUnit0Lg4ZAFI/AeeYhpN/8HoVIU0WQTecGBNAjfScN02PQ
JnrYebk3S9fC4tSnc9JTMWzB6lRb3cqzSOj++jdUriSEWjpmtZkrskRfTGxFxvql
heU8EZMcWeUx0RPqoGGOHT3Ir9imbOmlgKB3e4vOR93+hywQ3u9eg9niNwLWPsQ1
7IMQqL9bfbAuREpd+seT+1L9bizWC4yyt4d3M8BdIqaX7PyZd5f9UgsxeqZihva0
y6g70aJINN8NeC14xxcU22BxMzxvCiZSZkbeIMHYyzRFKH3FO5LVHcVsIDd/YKmK
PZQBsrmX6cZ2WJTK1bWBKMoHxpKSFCnlDTn4Wax7xIp2r8WxE0vzMyHA3QDtXkgw
NIo0ngEUQOZOdRvRnb2+xXKFKvPjAQzYoX9rPFeSpAtsyg1Xs1PL7qnGBk81/NT2
htP8UGmWfD6vOa+WP2YX8VjsSzauuPPfj35WRsQWu9o=
`protect END_PROTECTED
