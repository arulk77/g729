`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
CXDo269tkFVLssJhCUcbkePpmo4+0RZxNB7uld9TcMJhkcoX6JpH/W4c9apvvnAv
hB+fdhYxP6QHk3OGcWxKjnByIqkBjExnkPhCk1iwtetL7U72jS0w2RyyJCTlUC7j
lFIkvxqeV9r7aY6C4fgk93lHQKKyj7vUVgRyPveamdjoK007PFYtcuCmvm3xmANc
`protect END_PROTECTED
