`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOj0vKZzgf2pEkO+P+mh2rEzu+Fcfm7VpfmWBHuGSKWa
4egVff+BuspveHD/QkcVunqYDa+zrO9zoJ7gDlGbzhoX6fBzVKSipU80GOyR4LcU
GEbm67OtPNDMiRKyQdxWJqcgWBaeNDinGoGnkSvVxQc14+uQLNrthALn2icnaEQD
IWNvSf77z23vIjlU6xf/8RZX7e3pH6B7P5CE0GA2teR7JxLm5X0ZyCSeoJKmPmVP
AlCQH28t15RnYCVkKsSqTw==
`protect END_PROTECTED
