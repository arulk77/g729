`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHTVIB1VFsYz/+W1MJVVgHpsjOQ8DFfXAEH3YhscLbef
MxyY7BGUdQpO/qJFjTT16bQwgHU/Ka9H83VMAVRWigRES10arBI5GHZ90yqzpNuF
PY/TVG+dgC59kmBnrbT/P31GjoVHKEXR2MKGlQvhY2o+0zHwsZh7Tg95Pr6kPCgK
JQyuDzm4D8Bf5UyxSk9nNd6ndTbgDbZZzkHa0qrawMkhKD3LdsbraZV+/3s9kocH
nfo6CMj37PvhTbVC9iLF0LzCC85H15rYh00OkV0lv5uCZvdxBpB2YyRTk5H0Ok3i
6JOADEgDqo3Ly79z80oLk9g6fLf+s62RZ1RqyV8uu7T2Lv3cnfpmYrvmOhlMLUr+
c0zgqNClELIZmcfC4/DkSLyZYKeUKTiy6RiEDFSigRnTrh53ReS6IuXBJBJCFTlS
loMl8Co1OB/CKe+H6OWcOzLsqRRcWMVNRKvlf1BNe3acV7xvN/xhSo8G0qJLUC9r
u+LSNPHftaldJXZ4G2QaybKuzwfJBW5LXO79EFYPl14DxTQFq07EnyJ0zv27C9nH
`protect END_PROTECTED
