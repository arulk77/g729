`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
02g5fxq6bxKkJROm4+SzQdbkFQTIjMR6l2XBObusOAeqTA9OOJvVjMYLS2Ol0sW2
+CJSQUxmuydcLO3BK0LnNAkTiwrteoQmXZrVgMb7cDDeJIJLegyrXmKf21JR0Vwf
VVdxBEoY0PuMX5UogvGFik/HfKpC0LMycMhsrIQpKEPi/xtC7u5Z327KEvkK6G6r
VMs2mWq9ZdDYWYwbiApjFC8ucn/2b81ZIL4h8jDJsfPfyG9OCvcySW4R0aiK7gtE
Dzm7lJGPI4Yi2RhX7b4xW29IYa/ZEE4HuplsV3Bqd6IXN+yQw5mo2XM2lo3/5+Jo
vR3pKYnsfE8riAjZ9R435Ka/J/8SuX2HD95iWGjvkU345qCJ26shnNPpElUvsDun
Wj1WMdeX6e7NiGm42erVSSOc8HKPRLqqgxuvI5ui8jR8aI5yFq1pkPP463q9VkvR
bnMq5pW5OieGCHW3GTmjC0qNNteGymax2rXCdcCHGARrsneW1WQXpjkqds/8n3pC
7WyA/D613ETa+ICsj5MhWM7UhXdTiUusnkZ9YindfCb0BfxdTosWgH7ZG6WpwEU0
RMbWqbLKoa7iaVSi/12AUp8DmeEYoe8Pgv/GaESthT1Z61h/JaJ9f9h/wzFxcWEL
dt6Rf/gk0jwdFVeQB4vKUWOfsHs6LIWHotPndi9ts3IsWFNnMFJXrWux2QeguoO5
r+mWaI1k7kWtJBLPG5Om7LqSWLVcyIy05XQzhWPV/GfPV0DDsAkXJIjSklPgUCKu
USZRyn0cZcukUPZY2CN+ZTMX2l/Y4g4Rv12X7CcRgyIuPdT6YNfGkkoIuQa0+CRw
c1OVWrpHU9nEQPVfRzb/8QWIeALwxa0CzZcuc3xDRxSI4zSC9iGfZiwdATZKB6be
pknqMEggWxXjfckpAuvAGgzrqzfSYtkOmMYEiOEINTN6ykqc+RCJjckNWeqyGumf
1cVVMcQ4zOHgFEQqbV7OPmqZ/9rm4rzaxjskvlgMRTaOidaScrStev6qQOlju8ub
DEPH0AYtzAPVukam2sQ2s97JJkaAaKg6hqR9B804ytS+tp2BzjvHZWoRJdS6QGXK
hXwsMxZL2X04l1DINWZRZIB6wUXPC2gThmuFpc0EdcYPrm3O1xZTC6u2nhMQKrsR
HfRuM3al6+Ve+jLdYpDa+K5ogcSB6Rj4KhnhqlPWe2neSCXvHBXXKtYZjeQwQhhU
+YgRXsEuNfD5DkhdXa/UlRJacsbnyZFAYt+UZEYw2KAkAx5IHhVuziQ23w1G6H0O
Seol1uPx0aX49QqKEupONkWxUipwGo+L/4HKdD/BUXNL8Oibsay8nrM6Rzi6pOW8
gYWL2XXUXh8dZhsyLgus/6q0S1rwe204jLbBKfNEUTkhReIgsTf5rj6iD65xbUXa
`protect END_PROTECTED
