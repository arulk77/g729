`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFhwgv1nWutDyhc/1zyGN/YeF4LS8M1cshdh6P8MofRk
CLwTYIyIczJif7pOPwiibWM6tUxRBPl9LsRh6371OcZ/JxF85Bx/vBro6YAiBJnm
x7dZq2oeNyZz2iB13I5NKPFkoEuqntEZtpXPyicG+RTWKd2dBkDCcXKn2XshnQtC
MhuIeHvf8KfJV6euukSFIeeweiX7mD5cbQPa1FeIYi/7FlSDXPrqJUn5S47ML/I6
gkECfkYQKiU5cQ60eYtYMaVBnBVG3nKdfQqb7wOZiUg3RZH6bKMp8C++dnc57wKa
aE1tKZPKZH+3oEwong/tyU3l2JeBRLW7e9iDioqPnQrUTZlCI2qXknqDm3195g7u
GfO+CHljLqMjvLDXo28JlfHeDfOOd411PPKAdsySFZk/AGbI+A4PwcW3mzuntgzj
Y7+fP/vsGMv7An8ewllNjkyorh0N55EK0nWToymuiT1yX7IFnAm7WZgyTTRX5M2F
WHulO4O1woHkhD43Z3ayrC1pSKlVOl1+MO/PVj1CBA9MlhV6g89zwtSEmSxhnGoD
ud3Ez7X9iditxKJoOLPqbhC3bj+qSMeWMdi7PpoF+yt2kVAburzaFITYkvcMDWLn
`protect END_PROTECTED
