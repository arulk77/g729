`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAXMRQmNiypx/aGUctHR76Kq/CgJK8GY/6uchO2gKDFL8
ToIiksJrtZg2H8GtHmSEbHcY2u0QT7ZATQ0ACkj5FrDR7L/EP/J7hOlM6LOXT4Lg
AEoViABmZ76RPUKeEJoKFCbWzdC+iepzjtZvgUTzAb5u9nbTo110ugrXEMQvov8p
i7aeV4rjwa5F47GQ0Dy+lH5QkfIG/YoSReC5gymwOkLm1sb71lg2baFDzyqaOs3B
wdjstVUbzLLzPIoRkDVgHFyWIu9NTXK5HvsEtouVmpysmdTSegrwDpCHug3wR2jE
jdTPeiEHgacGg4L5FKDv74W5baDrtDrEz7LL+V0sPfGbuhnXoKrA65q7KHxl6PSB
EuNzbarqLhQd8+QJ5vWglGNPtg7FUrfps4ZG0TQiJFyc0F0ZBj0yKal4jNUthvmi
Z7PxM1hjMd0Oroo26QYRnjJsBbZIOSKMNH0mUXQfK5xESV/DsR8KIoiORD+xUnu9
wiTVHWDoYMdpWggeKPwpO0LjIHaYTe7ghY8/ulSzEFwfixihAQYnzkGRBfPh0qRI
IyevHyU9o3iqx9PE4RLTdMOIMZhTDfuLQJQNWs6msG7plMXn/JD0iuQfndjQaqni
K8eq+tFTnm8GfMwVu4n+XPz1dWdS0ctfRtz94zbj8g9MJWAq7eBCC+sht37/nchX
FAVNFXxjGj0Mu0w6NjKXHBQuI/aqLcvkyfkFVGDFQDE/4yaxo6JlHHsC+faVjm0q
HisCt9iY/QB3qxTQ88AhMBA/Of/+K+A0gKa+xHeCyivOCLWhuVe4f0oc4gDKxhoa
GHJ7sRVdAm2DG3ozU03SPCWS7bU1CAn7NEf3SWUxK2NzAQa53gkOingOlaMYc3qq
aj6OM4wGri5Y7IQgKZ5hwQISE979Syl/SzhKiEHiqCs=
`protect END_PROTECTED
