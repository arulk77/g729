`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAWowuAvuHkRzE9w0c0EJBk+wDemzrJMIRcWBSSwYinDP
hgtbpqu68kWqzidOu1KXBYKT5aAfSSuDtu8wY5H1uPHFE6p7GLxwRU7Z443Oc1lG
c/L3zo1oSJGJLFYmUj8m/iJU4TKbznm9sLRBLWcPgA6SUMAOAGpAlYJMDOAwzBPh
qzr1NNW3kseBx36M2b+4uoMXfbe+p7bOXqFlJ+f4krcNjrqXjDEz6omyhjGOjNWW
Q1T1DQtY5la15hvfhY6Ccau7MUKZ48rbi/Jj1Y/hWXCMuXxtfyBIEjGl6JRjTOuN
5o4NkkF6rgQ8wIUvyYrKAvJMwiGmBc1y0G/Upc/84I8ePhtwn6pSeoFmzIepuPvV
UDyKESzsIW0k7XWKDJyAfQKoxgUUcwJTy7jcbAD6tx3TuENc4vlyer8vKTnlrqrG
gnkC7immW1Ml1jgjdTzkD6m5Dn4JZTvk7nLc7WufHO+q0AQFQJDJfiMPczef8N/m
iBmVo61ehnMI3nYTW63CG7PW4OPsglcknescHByXfkVqiuHkC+5BiqQd2mJWFL3d
KLbuN76Fpt9lXTQh18NBzumER5N4Gs8BYPV+9C2tIkLglxAGKDj7jJAqGLvS/Upf
jYC1XwtaAQkjnvw0cppV4AL0zEoAZYy4/NgemFmFjH9BfyBz655sVsKTbG6M8wXu
+NG0IjmE5xweqpCUAXfL0hSEhRmf/mF54mIeRYjyemVZL/hLHTD7d0DnA++Y5pAI
kKWTtD5gsGvg0Lqtr6fRCsGUf3zUuJ8xqi5/BOnW/kq/2IUUnAlJPYBHL4TzCe7s
A8+yZ1ZYEQSnJt48xPpfuT+pwd9SnYnrVUTIChRl0yT2Cx41i87n3DT84rh9ZO+K
1R2kBJTmHfQGqrgOSgwktwuzux18K2EWLpyTI7YWAiprbrK4EMQu5zS9R/To5wV/
AHf2kHBPQMw4XdskGII/xMa+6/HTWuucYIPjRWCW4UsQCCKyHwf4cGPT7WRZMrP+
lIYnhzUwdO+3/wetNaPEJ17EDzjLf12+2Mouk3A2Wo6C9ciO57MD6LDPnWEyUfv7
TR/qUhQJxmO0Rohhuyp5cireGetiEu8uLuvpxZTQ18gUpw02aXJfh/7eyPdlJFdq
jmB3a1Y366GtmGYAUaZyOxcbHUxFH0lkTllRTpanEonRl1GMXtBppkACGv7EFiv3
1/nG3kf3iRSf8scEgjdsiT5gmZSVKidvgO5FdPYkBzMG+etHJIBX8yXN6sAEGmTi
ujuwglXzYTvIvIO5rrN7UVEc6/NCC4H9+J+iiDJvXcv/UWxis5/o56VJZxILSZxh
wKJPHhVskKzH0T2V6kTftVWg2XxxXMh5vuhkBOl9hk8jKjq/gC3DJuYOO42Wvlqk
6eroxsfqWb1jl2LQWj/B90FwvLkvyNfm02v08T3OWIDD9YXeDAwV/I8NkJ/qjRfq
YMK4sSYUlUCGXu+YD+GSxYgUXMtiZkXu5h5vVROtSOBRSQAnuGG/nMKdkVhHMKIN
cmVec/Z3JEccouKshqz9AZBXNQGp1ujVNqF+EnvUDuGWfNINiWt+Vco/GLMgZqwF
`protect END_PROTECTED
