`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2RtTiaLwZbJSuPbraFO4dv35fsxCibvvj/uPnDo7sDEzL1OaEl63A9UsfmC0b3se
bd4W+/UeJFqLAIbTl5ouOrsCwSjXCdjkpfKDKHmrxHGCszcFhZTB2lcLGh9CbxI2
tXRJvjrfAwoddMV4YMHiq24YXqow2sNOGLN32xumO9jOVsHnns6bypPmTX7qLdXd
`protect END_PROTECTED
