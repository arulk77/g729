`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44jXCk+m3yxu8BVLg9V40A51Apxkvc1uhT1ynp5KVQ17
fscSm6b37bkAFn2ULD1sRBb6vRUY4qQEroC81c1IedJO++cw+MHcU01UcSt9msb9
J7+tkKhijOKBoZdDX5VpWSd2gwvyutbRKP4PwKUOeGbSi57g++csPRyEnVlMR/Sk
KRubGrgDaEOn606pVvyM/r/Pdt+8mE6e0V8/3rXljEbPb8diFOaT1EBBl7yB1UJL
iThmYY33OpYJyPa/VzUPHE8lqU63uB3ZQwFw+Ivbxc679aoPZtz1G/ZA8fu9grx4
zYEbWKXdelu5266q1aPrahgXpBmaLdxj6LaXtIZPHA+qEnlKEmBTuOIHw5GLpfM8
GeBlGjzjWQ7BMotXcTccyQ==
`protect END_PROTECTED
