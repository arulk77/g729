`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOUnsBq8TsfQVWXZz87Rn1TfxCvs73QbfiCcVHXFFtid
YQYPZv4mK1HE8TLCqwDSZTiYCS+i8n960ZpgJzinmMq0FObPMJJNHXS+eQGSbcoU
K51ah8+PTAixzJA5sapzgb8cuYA5c+7RN3VG6m/EBW8ACvWe1+U+ZQmmkOgT+H9T
YxLq91fclZ2OVrOKv1ipnCsNGuHvt4VzGOjDTtYKCwu5UUssnqqxCoSXscqG4V9u
1xoWwSqnRpd2+H41genPLMxjg0Q05JBpZI6Ml/N55InB8Md0nEJePWjBxT9PRKn7
kv2tVjuiwhuwEiiA00aaFDPj6sAAtrXx/15JKfjLDpHBPtWaDjE0zGMZVhR2rQx6
swd+nyR+1Ih+SrkMHfaO6UDFv2/TFUIauFwXm4BhWQXX/xyd+nGbJ6AnJLCKA2mH
/2uGxLCuZT08aeUyIFg0FUmWYCA2spegj1TyeYjDs9M3Ja2unSRV0FYRl6W18QoA
`protect END_PROTECTED
