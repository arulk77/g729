`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHh2zvVFoi6hXp1Li2tviaaMvIn+XGJbML/HWJzOjgr/
xFHKuleIqr0U2CS+xLk8vJk1Du0fsI91EdbbmfFQZA6MC9GWuu91tEuhQ5oJu7Xd
BHYQ6CA2PrWFncomgRCPmWHwoPkw95xvPphdsL8acof3JGngeaR7NiLeQsth1FR4
`protect END_PROTECTED
