`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ/Ezo1EfGIqnQPjqiyBYtBf44gn8roYnZ9p4KU0luEC
0Wm7MVtyUGqiKVZXxMJTI2DMDWPw6DRk4KFn9y/w1VVEbfmVdF1/Om3tgLoDylQW
Z1mq21M9XNH7uiVCFMRQE+cZAMwu/PoqwWjYwJ5fMABq+nKYoyJDLDzKqdnVeI1F
sYhoInbkX3BbQR0nRLjNmctpSofcKHd+fiVoKfxYmV+0sPRlpgRw1nmNu1MY2c9b
`protect END_PROTECTED
