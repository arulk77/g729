`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMt5gdBdti9Wbd0ADTGIBUCoqlwqqfEteojDEh3Fb8RB
C6SkwNIZARZj07FDZxXKi1+CxKWsNxcActT2clejvUvleuttZceI9PgNrlK59KHB
u8LzDWpQJxcSulmBwpXYssdOrISiMVeVjkqlTpZ0ZugVYmEprkNlo4tFc3JpNVlk
bE2LmhuQLFAtbSx4Lq61xXy92XhSmekEGzoJQBdpQWwWIzIwrkK3eQK4ZhP/olph
UEi+r0/D2nF7e+k7ryrtv9di+1VpsSjDkqQwskTu5RNCgZ0Hxm2MJMd6Y9Vs+d8N
XfKGHwVNei2kqFcLJsiVC7C/+WL/snJJT8iBPX9/kDvvX/fzfHT0SgWLc0b4nWEJ
UWxJVEJoEZs5o1DgFj7DG/EcanNVU8CsKDCpknZxUhgKxvxdpLCRa7BewJBTW2Ee
EtyQhAMIkDx+QSaiH1QPdA==
`protect END_PROTECTED
