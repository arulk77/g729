`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4680VGYnsp3/FHPz5TIQEGXQUvaDbYEmssCHtGhuHXWN
22XuvFGdS1meyKDSDy76GFEAgsUhL2f80Kj/blMDcqPVQQgpsE7yhu5VpFZo7A0C
vKuftBhdHRpwneDcE4LGvRYRlYgtE3EHHCRFEBDQLR8XWmWzpq+/X2cYcxk/J54n
VxQGK4lMuJhFcJ1YusfTbp/JaeUqk9sLY7gGeWRmNFB95Nxy9ZwinMqqGo9c7uIa
gtsI0Yeyq43rcGWO52Lu+jZATOLC52QI5MOwbzA/B6ysRIsjHAjbc0YfLVHj3PcF
q2XeSRCZht2r+2JzSpJ6HgfJJgurQ2TpWj65Xnam9ZKhBGZ1WNJj0PG3xgVf9vAg
vZ0CTJSmLn2lLWSQR5lb2YPLLBXrrEaGEDYTwnsSDE+eGEpm1LwBGqnkKhsQGrPo
YgcETGXfNzTdf5V8nkDMcVBfIAr42urCaXJCLcd+E0w61eoYps3ACc5taGixWHLD
GKl0rYUdIrynsQPJS1be7ioFLyQgygY2kJsxMVWtuQccDPUc3JnSKIxXlSOmLKJz
g91F12+u9pch04580VIo9Y1rj/UEKF+uiEp0+j/aWNXqT5QwE/TI3XMChTdNzTYM
B0bhRVMR1tVLSbPlLWiHfd4MDAWWu1PJdfsD7hZOBjT23DLpR3j5Hfji143mL66k
uzQeba2nIAHP7XmSj9ZF3eSwwvtoFE3ESBlw9yrOPqtWEzOpp5Hpl51qC7hFV7wi
rhB2cM6mys2/laboQ+i9Qy+AxMoAeddOH1XthGjbnmXcmeVNZBee5HPmeHl+tsWv
zh1ZuKEQ88jBx2BdPkNIpkxEDUiLjGkpF9CEYfk9o5C72CeUcGek4ZpayIPZ3kVy
6ShDJw2PP+1a/NwZKuEmjsMLHhlHEYIYWGSZDj8haq/8Rr975fXYk7ZuEa3FDCw9
rf4rzDlKwyHrY7rhconyVZXkMsc8te2th542smRVD+GQhCrGiefoCYHIvaU+/vmS
ZA3y1OhVfekfT52eAOMwhi7qJEl0+ilAcaps/IgiLzB2Orc/PQ6C2+5o077FUmv0
I8j8yahUG87X2lpFrGqFhHj9XALxeFDfJfrrCAYEzvWPUhvtHvNK80lsf3kPUa/E
c1qU/uwmQiqhwcWuzyCLvCu7Mu3EVu4l2P19i+dWnbRR0iJ9Y8FjqJFgULEQN8jg
iE9lx2Ixc2psUd5BPPrdvzb8PTSqRXZcaXjtwv0HTY7OdryXkj24IZIX/5sR87Wd
TsSd5+zvfkFL/ZHEjoKSB9ohy3uJmYPWIWJWH4NeC/QkEAyol7Hbp9ylof0h5sKF
x9tV+8ys0cpWg4Alc46vuxFTT8pGU1gpMq+pCfHtl49kjQILAipHQMDGvWF7O2pG
JWXIsmUBhbefQm6A9CdPW/ilMevcWpbBlpOaqin7C6omqxKZdefHWBzwlB1Y3kwM
byFqKSxgiGGxDRLljD5fvrF7YirYNdb2kxRa5IaiDze3nWqmibXBqlkhh3WC4if1
a9FQ7VPEZ4er9xqYvCLmRM3Hc9M6oPPLYigYNyjngkckpQ90rwJiMeqpda3SrWXe
k/GGawVJl5BSG07ie9wLrOgR3hR6GgGaFG3U3a9G+3dDtK4RMwJTa9aNXX06t+Ej
K/13PwVXhlWyZxVn9xrXxejUJ2pGxG29QfPC52fv7vhUSu0St9wBbvzb6WBIOi1h
oPRfOZ7aBsy3yNcEMFqsR9pPY97lbMI9G0roSZ0dTTKMufhhsTQZPcQ3qJ0b7uSE
x1le/dBBQ8ZXwMks+pnW/WRXzuZXZ8xV+IO2FUY1dyn0dpjex6IVW+Ut2Cj8XfY5
UP5XrxGvCzzT3fdyl6WN+CQ2KjnKzEHxNAIOlJ4M05PmPw11zYA9rC+tEfLFI4Lk
ROazC/HLOMNBh7UeXTNrYrNNQ324vbOSZsD/6ZkjS6Zm5fNH6R36Akt/FMBws9nw
6rz9DivLWilq1lwG9nbKU0AEjvrgQkw+Kmbt6O9ouW+zpF7ThGGoiZelPKgzyUTD
8sGvGdd/wD3MLR1vgOlBNlVaQoqm+6wTOCDaCI6NzvoPSwl8sVgBNM7YXU8Doe3b
kdnvC1Jtrl8bPFjqr3sa6G+8U+gC5ZWLqs4XL0XcLFhyXP8RcHqFy627YD+EA+JA
fwfFLV3UrRjmyexbnPHb1xRg3a/e8m5KKYjnXmXZ2PI8Kbgl87fWvGhiJ9O5KPV5
WOLjr01MEc48oxQlx8qDsVao++WU7jR5vk0KWMHgyl7Ata/OHBKTDCmMkd1PfoHt
UwZHnb9pMDRUUojGsiS4kFwtRXpHmM9h/zBPY9X9h4SrC7kddvEmkLTfzOnK5kiT
O2XO+zkSpFyViJcS8G/U0b0Jw3axax+z1Y8UWzVkdgn1xgqi4Un07e0zf7Hw+SgV
f26etxfjuPZPiHDOlpvEY6ZLHhJxJTJzUg2ik1S/TdBOHSbiReWZN2MkwpUa1rx0
Se6Cv9p6Njc/2CyelkCN8ne8GNrBItPvcsEob8Ihq+MqDoQFArzkn+FKMeXYUdwy
3LBhULwaXpbIysJwBI3iIZtHVEffD5vps29ky5L1i1JtiLMS6NjNyuA+3gUPpE74
JGRg3YZ7GIaY4nDLSrEJJWxgvUuQjck9x1+4a78G95U6eQciTaGh+0ykp6ChuuiV
F+4AJd85ZId6Ilp0cCuBlJ4KEnpcN1WgUCjfXoOwm7NNI18xry+Xv+8KJ29BSJvr
1H6JZd8fVJX8iSXhUACuHuOEli5xDKkqkMNm+jZyj1C8JL9zMZWQBJ1TT7mOVfsY
e96cYL5VnQUw9N6gAasvcNz5tjtSUYL56KZpcatEEpubmsXZNoFQtQXqYdihPuEp
Hu751eB7Xk+MVRo7MHnCzEuQD7CxAzKlXptOdprnFXi1OYLIgSnpYI9jd5OOiuXI
5RUxI/nGaaaVcxCjM7LHOeaeAw5Oo0C5vW8n9TQ2b0b+yjRKHhISbY1FTijzTqW9
aAJJ+uWgkvWJRaMTL/NcxjC7TskErjHBrnRC9UY4RuU0ICIPZD45NvP7uqNNu9lu
OqktviAcgGe80BN7E9A/m0ElKaS9b3jSV4iVH3S0DXoOc3V9kcoDTVAJehQdfM+7
RpD5La8uC1fMzIsR/ZciQE3E+gUuvi4E17wTOydMkogsYd7SXEUPG7WSdn1+E3Up
NU/7X+QPtEtfRPRVdz0DBK5sOegH/IIhlfRMjOA1dxiwMRBuS1DQKfINFb19yHPD
Hjo8Hs1n8pkEfIiTGWFJB7xDePRCRCQiqduEr5a2Xa+XOYMu7Dwu0divavNoewjJ
1npozntRnhkIVBbqMiDRn3ob6TE9VLuqoeP1MKk1c8+GI9MraeeNg2TpS7/Z6URG
q4RAlXWFtJveCA5nZofQ94D92i9jdE2+K+cUPYQcRmBQVGsYO/Jlr4kXdbTOx8hO
IEZthoe18PcQaGp25uicm8O38wbxrFmySk/+/u+VOauNNTIuaMg8QkFKs408YL2W
9qbLUK8JSOw2kXxRxQissLptUomibuOQJvetZY6MPb3CT2hX/6OcWTsFq5VQDTWq
ieh6awI1vtrpooIbCw+uZ6KJ8H4kJtJAVkzohPf4/mwCTYnsIYPQZMbnZV/mEoF5
9wc/zyt3HcTwWZ29Q67BuV6HTts6Mdb8IaMyxwIvR9pSaYQ87SjJU6+sKHQvQhXX
Uu4mCgLRtDyoa0kWL3selpZkQ+Mkxj6kryguBERngHzROyaN9reVOjaUbKv+t/2n
n7C/eZR5SJni8SOa4GLZxz9NtkDdQM51my+bDxEfabmvsw3OrVl21HWsD8X6jEsG
h/JvvgUNmeUVEGC/qvItgAFZc3GujuWkEmVAG+cHKiqIY8Ex4wKeFrCGoUwFmBq6
yHSbkA9W9sQ3lxzt7OEYzKOAuRY2FgcZYbVBxlFRzzBcytwDkm+pUrfY9+Fwpqkl
rATaZ//jhT8U573KF523gGPS0u5/Ah8B/J/Z11jPvyKnbcoOuxiZo416vYM0wXuW
OQotp6fAY5y4+jKMNeLzbkPLtQuoHzbLjjBhkZrX8ZZI+9CGn9J/0Ykj4iFZXQ5q
So8JxkkgqS5v9H7q7BZRj2g1zVnpYL7VwllAp92UGo4f823NYiC0J009IDuM+L1k
30AHcvQRd0DtY/GBNYCz4a9cSUrvntQh+zTq7aUi9S2NZ3VZLkVkaPc+Ed1Y3dvk
DfAyG7wR5Sn4tql+6l2++aHcaCs+Cv76uZeuoPetR+KehjEO4qbKPtHaDsxH/mkE
7QfhE8EpPj/jdVXHGdAkByvdB1jay/MhpUGU4ICDnDfK61lwDurUQXDQ2MxB/Bcn
TSd7iDHXrKwSDEObp1AuJZOfNEuI8aTKQJpEzibu91YLK8H4nbALLUnR4prpDVZL
CuQmwBOSyNbP+PjcojAExYjy+eydE5/gQ8rKpgVB5uuEg8KeuolSZMtYoE+MhWa/
DLsPnaoSy4N2dxVO+Gv1ukyIFjSBL8neAiJog56xM84QfQwBOYk6Wb7ZK3PZxV0X
/W1kMCYh9sdQAWh/p553vYhmfVYpVflu+ZK/XtOBejDulL6+G5+waBTOXZuHIZTT
URB32kJ6oopZpeei6bVkxZA5SX76GfaHlLMGH6PJ7BWDK/+bEMA8Eb2CZsUnjdMO
tHvQhm3gSypop/Wddb2cn+qeJBl9twPnklLKQC4dCCeKTVz/Npp1gcDge1hqoFFM
Bd67eFSB/p+UqyQw0IFL79l26jxtLHvEb0IInBdEzYSDlZ4uryGJXr+r0wFGrj4V
Bvsg3qag0h2L+Vz5q94dRqyfOBjJ0UcNWIX/OwNPvgI3ufatTl/80vkrUiJOIPUq
2scSv7U8nyJtljWzlQO0g9le+BfC7gsejfWfR9sd2FN73Rl/CazTyoj+H2+VO/p0
FU0qSG9kZ9YjkCLedi+NxFu9j7p9I1/qsL7hCfBd329oBi8QHGs/qwiZZQFoYHPu
JuSN3Tvvm9QzlayJIMBB6PoVdXrLNcHGFjygHoVGDY6yKuQ8eHP23z/V8vJJnRfk
b9pa+FZO2KWs8qgtzZVkvrcwkUjkS3HPpgsUvk6Oym96/thJ6usGG39oXssegX++
oz3azbeZE/D4t+ucplOg1Qs6Ireou6ErzZR+RBGPKivEGFPSou1wyDoXp8S4MxLI
IAhSawTL7hYIL4Pki08ZEjhzdm13DgKMA/wwQra/z6ImsevUieyMC7hKCwoZn5+5
uoRtLfgDiV7yPe43m5dfBiDfyl4S3VytCNZVJWNtiC1PnKw2soVOcm9vdG6VUPe7
gArcxepVWUYKpkyp0BHoLGlNoDnmBvKhwVrK5PeM8nESB6ULMG2Lh/QRKuMHUTWz
EHKd3tCLOuLFCOSYX3ClcNVJdE4WICiaE56UEoh9IYblbhxpsiwmmUAZdkO6pZnK
OK3238FBOoZsa9zC2Mw7vnLb7RYWJ1GPwpcyLiCBHwF3Wkr48eQzaXerbvJL9w5I
tpgNA0Dbf6RTol7CP/aoB2Pxspv84f81Ra5ReiS26CrGggAvUIfNi5xRGJbeqXZZ
2BJ7AmaRfitDSM22YHOrMOc/VWC3WKx8iJmFiwxFk7UrCSyk8xq55M3e7HAnwaqr
8e7GxuwZfgEmZePeXqEpq5+SJCaiZh6Q/YJnfEDtvsfv8amxJBzS6N7yj3jn+bpU
rC6gznLTnf10OkNp+sdHG7o7kOFWg/ZYHCFSjMgT3vppq5UhmAVw7UGvO94i7dWA
grblNGMGCdmXb2e3SebU7lRAYIcotPG67+uWJYlDOR/Ij1LqpPEjI9mjsBamSWL0
yOAqDuzB/D7JXFNNq3WQRyBdYpd4KNvfVlY5bMs0smjswaImQdeJch4ssg14qrL4
9hcRqCcUGvXXvbwjjaNPaH56VS0fvcj2to8OnUy5ncr6CUqjC259LzYqxqReFqkQ
9lU8G0vwD6JEhLHwkxYlec4R2rJNn1PgDwhWh5Url7E5QZJii7OMcrJ0x3awrhCj
3zJLz7lu0vLOsmHhlUE/K+ZNGrvIVvynYizU9LnXWRAgqWdLZVSu/KmYR/Q5ALKO
FVKRmi/mdQNIK4nscIcwVnJZ81G9EGYgopLGAkhp7d/wJLBAAjsVay3BQXK7PyhU
xZzWvWdIa8wI6rjnCZkh3yWnVfdMtsMhqfAs7l7mutuTQLqBNbLA3H61tnxl0pnK
GYnnS8u033SxYH0PAf9yTGAgt20nKvZ4f9q4BbT7rb8WQlGLQu5Qp16ncdDdb1R4
pxh4BKvC1Omu4BWoTSNLEEUjBaHiml9AjA3ChINI+g77fGdAE/NPQyE1yjItBBc9
aawRWr2wgzSNQhRYLDQ9w9NgHQ8ZO/QvxzkuKT9CtCqOyueMPsbV7Vg736YYM3yg
Pry+SXuQCZahi72L/Rq5YMzDc9dUvqf2oPnl/7BkxY705+RxT2F7lW+xX3a8SMRz
kRDf498d3gW16GVN9BBb//vrfk7t28Y8vpSWAqTHe4JQnkurW660wQK1jKUa+fNb
Q6jM/OiPBwNqs/JQEci6pVjXzjzbrZ/aN/D1rQht5J0zOftxyZDvpi6OTpbO0E10
riqJIc6T+eljvRnHJ1GcTfFRR31FgbTCOF1E78x6xjojQII2FDAxQ/39+XnQE2ER
w0UAVSILhy1tIOSvidWKnsXJuQ4M7/BHEIOxLUFurG4OMDA14BRwQHEgUWzxlaSq
yF4nRtEXXIYAa6lelQzqbuI2PAME4NGr4EJaa7WIjsGw3GTn82xSQJ/avh89iCNm
QLb94SAJB0+jPPkeTBinId7r9SaO8Mv7SO8hZ7lefSFxL9/4Vbs4ReVGyMWW0nqx
zLmOKCEVeAJMKVTYOcxQaidPtfXGyIK0Rm7wWn9QPck/fNgpaQXD0dNfLANLxjvt
HCC4Wv0oAb9F7QPR3qN5of9/ev52EBjgjkd3p4Z/nhJBPbo0Z1HTsnruOar5Cxuo
879GgaNDhZSdZrzGGfh9T4Nri8SMd+K4jEpV2DonRJV68WAV9ko2cojnDd856ZdB
o50PydlKuHXGpHZ/1BHJTwdFPJITZdsGkrOSb64euiw1zwqQSr4KjNvede5YHahj
/Ea7pnPdBLL5jc1XWVwcfKKS1adEsEgANFX/6t0fQjHUD5wkLTqCNJ2gXmA81wQS
4DC9zridhCMM693BN9OuFpqc+9a0FE5cnY575idMthWdWw7M6yrsgoKewAC91j6n
ejFQZe4CvgOeWvXrOyNxaar6wN4jxA+/gzkbfnKkCMYJG8CKIEyiwKFzgsk57vOx
0uYid4yC2T4BwZjcxYhGO/3MQvvvauIj7oCCBUiSO9+Rovd5YRRMzs6VW67FI6LI
A0QtOBKijQE50hM1o5jW78vZHyVXsAHbJDReNkaM6iI31f94emd7712c5N9RhSGQ
HwxfijpvyLJOurBqxBD7mJOFa4cLzoIjHvueJzhGF+j1Bl6mz3+mL4nWmNJm0NlB
UIe8/GPBRsSh+UkX9q4loRlHF03Ro6wIxuyU8Af4BCV9EmJ54qtRYi8YYvf5NFyz
4iVov431Ci1QkDiV+w1Sm1vrRur65kkQQ553z53HcY+/v6pgUd+crkq/ckpPc9u7
lup2E+WsC1L2L862kYiFcuh2QW9G6jan9lqv7cylgZNyboKO5wxjPj+dMpWVXsXn
xPUwlDnndEbfSii1Pj4YwhWoOuEbCxJV8bZ2vYRYoFMhvLYvYKSHaIAI1cRbyHRF
+rPp7Ya1bfbDbN3zZwa6BQ8WwxQr6BlmMIn00WoXlipomb11A5p8mU0stjsH3jsy
Qy+jA6T1oM01DZBK7m906SSh61eifWGOa1AgWKZ9/UzRq23TPQiNcncz1Shhi+q+
zStO15ny1m5U4BQpfbpGvtoQqLrx8TuAC2nOMGCkgEA80S2OSpaIgfLnKK8u4QSM
eid0eGEQgLhZJxUHUW7KWplbnRDLRTXw+XCgErOmp1dVlMSUQuGjnJ1uSAulQS/B
GZQPxLr8r7Z+X8QY4kJnIerHuLA9n1Zy4d4z8Io+41BZSIGsAc4CTvII/lNN/Wtz
o4fKpmoH0PPBG7fDaWSWz/U89a7BU7iw41sGclnGDqbrfGRUcBtsfIh1Eoaiv057
iP4VHj1Fn9iImvRRSQUzdzQftW6tCzoYfLWGrNXqhyIZ0c2RsXMHMX3tLc7SdmWi
oYGHrmtcuFWNG6bnniGZHU8PRnxBmlWVceUwuVLpDibOfQIUExTZU02psYBnwNrK
VU+0wNG88wHKdiUijOKzUrvStg/PLT74ig2gG7i0GEjvmyBGlQUlVtprIaU3Qo/E
sB/j1GFaTAQ9zzX0UQQkVNeXN/8gN1xArYySrZjGhIiNJXeo7Z26wRmq4XE36qh0
930v3oZ1pawiS9J3zquJR5oo2F6IA9ELsDP7kGUfx5p5urvEOdz8xSBzr2ZiKlQ8
/eSy2FsN1jHIqThMOaKiW6u9Zxd8ZqkMnp5xoJdPYG/AqYWaIC3w76MqLl8u6RS8
yertynRaqgvacEq+D6w8z8HI2Wm+6YM+piNT79FCd32xVhqONFDkOT9t3sYovUZS
WceKErax1b13rvzt4+WDttho2oTkTtuEeN+puIzM/b7t4cmARw815DdE2Vv5Ky40
4h8SLNDJK3pDsLXQ1PShoHQ8zwIGOwz180AhISezV3ENb8CWSSE4Al6BCYqckEuE
8iUNwFV7X0Xrs4D+XjzBjufkQAXdTJpgd0GS+FXQA2CSBnuoxTjGEjpuzB0C0UhJ
rqKtfEoKCweQss9qsqPxRnx9LnQKmpcHW2Kqni78Us89JE1jOxKHxePnYvry02Sy
4t0g3M4lnRhptXYfe5OV0FWJa/Z6b/5ahOEGqGF2/rtyrw8BsntjX/Jna/k8r9Cn
S/clPDIzjp9Ic2pSiTqaB8AruiSw3Zw7Ty9lVcQ4kC3JMHG077XxzIRnA+L18UG5
BjLaSzwXUQtXqCV+3+ErA61Nk15WFMasvm73q4qgYkKFl4wUq+iQkKYIx47b9lYC
2h9PcCMJSKQrqv3qhhGhkV1sqTNRdq1MpD9XuYuXDPoYlTyny7JGPDsWYXI4Yfxl
gZbDvO4HPo52mUEte5S19ohsOVvdVih0orIHvAG0cwjIj+rdlCoGTeLBIN4raB5u
kLbeZnFY5TF4U1JTkTH+JKD70z9eqNXmtVDXNMSlNlOTnYXFaPAf3FUQpNqs8kq2
fsTeQXBaECVusCw86BzDwLan0BJkMw0l8QKXVOx2+oDnw7vxKyvCA47HI4FFj/8S
rsdXab8pUJfbWIRVkRCHZUh5i7WUW48Gj2fE/x/1Jv/fsl+WtE4F/P5WayFj4n1X
pJO+IQ9JHjWtcCjVwbNudAY2cOfRK5YdRutBiKI8obb1+nEIyToKgI21sOO4C9SH
4+rfHkZyZBwDNaCZ9PyFGGgYMetOaAKTpFf+riIFDz+PIMs5C9Y/azppculdoOQL
uLQ5aSs0hrGzle52CvskwwmBib6CsW8Tzw4DjkEAcz9CKKZa6Aue1vqWKPSbfXWU
7crqMfXECaWifkGRdgT/5pn26b98tZfTI0fqVyY8HZ2gtvXVR5jY6Hi3EOvo4Gw0
FOjpraw0B3fznDGzYnSQ3HznQXY8VvlPHz9xdOCIlGHqW+JuhqtW1KdwhbBO7UCA
xqwNkCwTCpqD83YXeR03dNj6OKkrVAAjM6cqxOmKNMs/G53iDZvAYRMYu1gvKMNf
J6fqd4wT30sW9dqZdABPFTkje4LZUNIu2DC31ZyjfbB5OCcVvdoinpJZn0YLyvSp
C12Nx2xodzIqlBWg8l9RWOynExaVdvBKe9awR8TbFBdProOZCoeg4v2dM9srEaBQ
B5KqYB7IS7WG97BdxKQWlcUObC2D6AUB28Qf2VlxeYUxt/brt6Ag1ZqCMhvqXC6t
gMB7QxfP4p0qY5kx4uScAIEgXj73+mxUaN+U7Whet6T5wYkORRg1RhMytc/7CCXb
pGTy8XKptdHxQNRurcOOrVszZLmxA4s9nFnYZXqwx8MxdA+Ggl5fCUEpEoKuckpF
CEOBRqkC0dH4gwnPCyyrJ+Jqp5mwaVEZU7MrpakFaxQLiRH+K5BEXyO5Oq2/yDXj
N+uhziV/ym/hlOXDPo8L4bMvnw2DxwLefDJmX0+iAV43dqxG/eKXpvoLwE/rSV9U
cFjrMradd3hhHnP1y2GtvemRE7RT0bwebWjyl9Wtsp20po1kCUOVVx2YAplE/4O1
3qm1KVk+0R6nCYgaL5kmGVJzj2jNBVbUhVOsZ/CGtWw2yfRrQBksP0HJfxOy0kPw
n3Q4fFMoKuqpmR7gRjSJWgVVZOl7iFPgffECLdIMVI/4YHnakqqlGNb8Dmmlx/sn
cU2MlIinLcLEo7pcGwwRU00ez+LCgBiTWtUpZ4XTQ8NRzpWDJHrLUBED77udcrqe
Q/OzxOcQPj+Q/5I6kiMR/7HAJJcSoYUn0qJXNy40fkiwQbFqn+L8tMxCvU8fiRTI
O9j0wi/psWuyiTiNaJmnQtsY+xSRgib5pfDVJoTM+gYkfJrp5BuBYuLxjeMlUwWG
o9V2GT84MFAnrq+kfgXZWfHL7Ph/gOZkJk+JDVqTTrLyuR5H1cn0Ck1vBzkJ05H1
vuTyjNvaeTpF4pmCsJWbv1nzHiEbLAfp16zZiktUJkqDeJaoSoP8QrKJleTv0kvi
XvC/A5/76JFc80GkdSDDyJULonmjHbKQeMXob2g0sevV6yIEnUMx6FB2xZnbnOPf
sdeQY7+67YV0/Eq6191BsBy2E2NBQvkhNVcB0CSB+4YdmdtYTQdNNThdTO+BjdAE
3sxdttA3K4uQBd/j119hneYUdUH6MiWxfIccVMpPc6ebKRXvnZ9PcCwvZx1UCSHp
15XycjAetORleGObMVZyKfv88hhgMn5T9XF9mRQAJFKEWPcUHG1MoTa0a6L386Cg
Dl2tIlFHTa0P+wJULyjTfpNa35XLdlHZEO+OVW0CMiztsRu7CqKbo8hSfdIFxW/t
XzPMe2kXZvrNRx61nKU6DtWbL07MapjqnnpYpZlLcFri+4/UJOBVFB2xuLLXTEY2
aNkAejk/d4RuT5RSuI8fDqWzz42xbh7NqhgxfgBXY3gAwoUuCdPoqfGPJ7QIRk9M
MztW9zTEw1qnxYLh4yBTsfsrc7zDgbwSNLkYqhTIRyMbmCtR8NXdBFXq8ZFMxuqC
h45metXf4+uh6zNVjCT1vkq+n+m07DfvHDwBlcZDFymNZlp+kSb+YjJ1LJbd4HPS
DDVISfkEG6+n4H24wqQF11qRZKgyYxm3IM5ZVb79ay7o6/c1joWn6enfq4Xl0C9P
LXgLszDY12Xd4bK48i/35hrXN3xTWTT5ur+ZWMFP1zDdURHis110f3vRpmQglSoe
024z9yDEnnTsA+C8p4ung9Pj8kko2DGIQCDbDsgUcyHlois2RQjHAxAdXNugS40W
nsWX90t1kOVQDP/9Ubra5lbZkm54AgdpvBWMVD811vhM+19nYos41KeHlmE/eAnf
ZD+/FN/1jscOamquz9yFDF5wkOoQDwRJAAZb/HAphKaEtd2Lspcp+O29kQz90POk
LMGBv9o2wgno9DA+POTKKCP38flvtsZ/wQ/wfpdG3ib8iYGE+KG7FQsPSpyPDHne
cvY3Q/PLZaDzdEQwzY8ZOCZw/D68JcZU0UFcJa2b5dFUWFteYPzzRc5X++9v9v/z
y1nGrVgp5aHaUG4sbUT2VzTwUXcRzRqNV+NJT8/W+l0K8ywaGIvAKRrYG351okuT
ypEkvVga3VV4DlT8e6uChUm2yGKSVJxGkXQqGmbDK71UTSIHVnlpt3K26Oy+uZWe
wCF8e7qbA3zd+Jo5D/27f6ZW73evxwzvRoGfG9m00o7ugEKwEF+/3YwCGCslr/ca
2q7uyubLGDK7xjkSLlmCtM0u+LIMQQ0CgwmGGd6QjpIgTEv69gb39fIdy87l41lz
yssyWuaM1JOsh6x6NDXHtv/3dNrDfR0RBey85lSUW3gpAmrFbUmodTBukhK6nC65
CI23rKPtEd68rJ4pFNrAL+i4mqZJWoy5jErr4pDlumY+vadx+CPV6xTXcLBhRasI
CtYiw+OdV6LgALJsLqsoXaD/QYP23dg6Ugdsb1R+xbjmG2SzNxSwY5mgM0URc+Tk
Vm15iJw08ArwgMdPP+MgkKYsA7U3XJsYcPlb/gNnVBrbvCsm4Q02K4VTn7zCLXTC
L6aOG/rXa6fdfHWWTlUskhQu+uKpPNmFPD80fkNPrtAHyElTsj3gW5XilmwzDkU3
QZAofHhJgWENca2bh9aIm5Z9PSaZyJeY9Qt/kbZ9ZzGkNXm5ap2jVKBKv7Uiyf60
VlsRqVi9wEvr4wlujhL8NnKkUnmyMg7bsQbLFADaJLgtarWrlQtkFYZBnmdRe05J
S0ereeVWQHTBasgKA5nBkWz8rX6lTKvFOfkrzvd7Dk+dPry65pPxiR9OJoruVCgh
VfG0c8PSwNEKFb41AlrjUUcIxlXj13T+poGcTHGG5tOu54SIsWfwbv64kxL/xgod
KYLIgsNTFhYCyDrM0PMZbNefH6Ri0ibxa8oJAbbAXVRbK0jQqnyrG4q8WMDIickN
DbHH+WcvbttpLUENxp7LkUSXvYUL9RzCk0ikf6e+t624pQMhRVCG4XMSjYFajHoB
Srumyj//vic2tGsgmDACMypO+IEUfasbMZsoJ+8lCy8OEp74lOptdy7OY3Knzsyh
7K4KaLv9CkJOJuoWGQTmBlrVkoHl/ksPlde/PROUEPXtsbGw9WUnS6htF72uouCF
pSVMleQ0slKT3s+w3nVVx7jTgaU58A2gruhY3lLpr3I2feNjgAAKSehdxVI/l77m
tgq9mDiFm0Pt69ZEhOSfuAuwjxatVG68o6qKqpfxJcx673O4Nw0XgCRCkEtmJxKD
ycp4luDb6JjUW/q6qa3xtILIMz1G77hDnU3OPs8EC/vEdGeWcj5irWOpbcLeopgd
Co1YF+6Ya0ORRQp2M5yKQGtqUCkjuRV0Tdn5r/gKW6lIk4gMKUWVUfeFAlaqtoLO
KLbgojqjchFfUh8yG8jTRY9KbZQF2iokHzXycjjYViNiYpjW+BQjHZPfpfxMDHbh
0QyrIGSfU39KJwUT3/uo3h3KzCw5Sle0Ud0m3NTRk2df8ygcP/K4KZkTAMkMgDMa
Efd4xlonU6+vMry9hwyyzesust6vSHcuRccM0gw8i2DDarL3+mj2YIF20joqCQhU
KeioL4URtotLh8Z7bkgMnVne3tCRJYhLwOTD1GEfIDd1gnLn7INKuMBlpDx9Kjd8
cIwM7Aroj0La55BEFpBkxzrD+WqdPLP8ihX/Gzc/TIGMwqyjcnqSju3jyb1xnBWm
HguQkmvpK3iILeTi+k2r81CeNKY8jwVe9k/vvaFno9NwdXhe04z8QonhZyQ3AbSr
0QF3/lJjBk4BK3Xe3DPrgbkaiQHcgm8+ih/SzhXaLpPvnsEmeqTqR1TWAYalegWN
t1+Si9APEmsKv4ZC+gzyg5vKDs+B7CTnHw5LI/qvr88jNIDiV7/cEL0Njw4cr0r/
n31565OIDbJYd51nqU2PtW/jniz2ZcQjjKZVviHiOSOqxPwzGa4MK86S7ysv8bn2
PeIJnkDW3SAxJYMbh9zPlD58rwjsl90riSNM2NyP7UTSDvOyxcbFWm8R+5QAy2Pu
N1xYn1rgZJlCYcHjSK2MVW0JmnlGc4KFTdiUzUT2wKy5DeD63bfRGiauQeNhpR0s
OQ0DkWr0MEZuX75MQJqA17vXbnsnH0tIEcMdUeikFzPD2tlHTgDwtTxNpTzQNRbX
iHHEw9djIf16J825qyqbokDY45hJ6yBXfhNCr+Z1XxPZ8QRfmLHB+KvnjlO7ZsBv
v9ZfuDsxdrVuCsHW94ICz7MdsWqyqFxZymy6Q2hSS6yUTny3gnpdLtlkdosCqzRV
KcxYyWct/FBIAyd73n3C2ge0cNcUs0IwwWoxL57b59L9CAHlJjau7eTtUjC2uh3h
LTnHyJl8NRnFqorhz3+opejUxyl85JEHHkT+/URHOYHdlrkwyUKE2utxI6/ybtUi
UYx8egTbcOYYOo2gJ7AmEr8LDr1lAzQoOlPVh25A19I2EZAIIV3lZE80jQkFulgI
bIdjjxlxDSHEXyHImExR/ctYllNXAKKR4//H6ViMH8RvUHAHkJJbLeaLXBarhRFP
i6Nk1ijCF/wNhgd69404J5OHuJncR2KlrDZvngO4xnShaLNN5mAtMnTNFfoIwS+4
ZvFK8oQ3MRrC4jzCMpoaIilS5ve74xbaiExumU2RkjYF1bvunu1qIXHzUDj+FfwX
UMg3L3UduPDoNTz/Sxnt6Hf5EoQcUUWjr97DWFrbW0QFig/EU8xDykUPVUf5Fo6w
PMyYjyq8AGZOloaG9OgMJ72n5XJOH9qSuVS2nnZMQ/M8Fzb3FTV5b+5jw1RnwKQy
UaVxU/NuPKoTyBuD/wKxWP0UZPhd0w12+Myj286du3XT3s19Ej3RVCoceXTrZBxP
bxRuLuWepqKsFmVTdbFxXkzStzP++z4TONdMEuT2icTVqu6+TgvQOmFuz0Rj2vcI
E/68bEE5Ff1xGzGhx2Xg7XuAcR6lC2ge8U02Y2gbYxspwBKS7wAoOWP06vGHmwr6
Z/beFEEd4guw4bTcd2+ZWaHBBlcqJe2YS88wmPHwJ25GVvR+Se4MhmaK3ooiGPjg
YVQIvQmIaHplvd5Zw6A8HSgcCx2yCPSJ7+kn6bLxGzHbJud73ksCL9QFGZs80zqB
4lgezeHwJ22DBpnsNcGCuCwCccB35Xb4ahlzpXuFiXTxojI6XkdGarU3TytAQdu2
VMGH3DtCiVZ+o+vCtyWFVuLVAls9qPyvqgzZ+K//zny7l5VRZTL7933JOAnZo9w/
Qg2w4cGtfQ7fr18bRQk883045CguMiHmsBfMH86Q4W3hubvj+5KaUCSwxXp1rN1q
8rMZL977i+7A8QCWrCD5tt6VjQHshSY2bHKc8WqpQ7MOXCxTh9xfZaAhgy/8mlsh
7WeEPtQPkydJtt2dMFd6hvffHX93l2as5I2HDTv1snevIOli8fCrtU2YM+EZ15Ss
Bso2R+wEyX2cHxv1/mcp7oBJ1JzYxXp9jBomuCQ0DKGYFOW41gw0ApxcCf9MXqoy
qZwj7DikHR+A99MU2I0ERzgJjcCsWSAq4Zclnd9KM6CC03OFxAE+32ohVID/ze2a
+zsd3WIywy490jQGM6knAg+0DrXqMF1uSlORHJssdlYb+jO9Ivi+4s4S0Say3aEB
WPdsXA1z6f060+sH3s7ZrYhz8j/cSotsDZNDLVfB9uXU5nVyKgkl7VC9MxLNLfLe
Pjfte+5NpJ8P9wWmcUQz1vU5WiUL2h8cv4TmiR87PhdfKNNpmVGq2OjsZcmDkJHt
b/qzLK0jQ5uTWEDjHLa8MMeVT9TSB0pOXKeFbgQHCi6g7CMVwSl0jVMfO34Fg19a
cwF5A7BhJSMkj9IBOHzbjmtFXOQisCBEEVterZooTCEGDbE0eXjeANhamgPBXoGd
2OqJ7AuUy94Al2BSy0ZnDPIWGgoTqodsoTKfAMKltiK/FX21VGLfo4RqU2Jhflin
KuCQhhaRcHEE6AvR8ZacXrxMPOJ4NI2WMblc1zRUvo6hwU7xPudOZOFoQpemTrbb
GKweYS/3n4SJYQYnhWkqpWeFm7Ca1VLiQHucZHoVD3Rs+NgUM8XBOPEmyABgmqyv
af2lxl7fLNuc2ks7fKb5s1ki6n2jfDb3NYXE49xJluLTyqAN9GiSEykBbvHzmIRY
oALNtULbsvoz84Mq0nlLkla0XZEZWgRTUo57Of1baLyLxamhuQpk+qMvnfUGG8Nr
ona5VNtr/l2CBEZwDxSbVlTGxAHEqmxoH1bO/YXDKZeNc6dvJr2z/idhklAXlzYb
NLWN0JbI63uzRsgxGpDGDrrLDzmlnY1cLQ8JSaTrv88WN6zzkaIL49PfzWTSuVmE
LKwZ8yFVk0OWgbYc/TdExnozE88HgvCe/oztmXNt6MCu+dna030rjEwfFMcqnHaP
apOmmNSSn7uSLXwK41wArXzcwVtZ8pYnpkTOPBfL5Skp9PnyOoR2qZS8UzROyv5D
bqdyDjyJeEPIJ+C9JK8moqUIdKZ5tmKhGBk2S9HaLg0moL2AqcilE12bkeayjrNn
GgQdXnOYupK1iVHGnkYcm0wNLBkEH2EQ87egoNdOryFK01xN3E864Ve/qeluA6TB
wf75DpXB7if5iVKptWYPF34B+N8xLxAVR38R9crfRHePfMkGvr00/a9Ri5XO8PV7
uoT0rV91+AdX/0h4dxnuMIj4vqAudnYTetZdsq4zoCHC2bH4TZfAmUJOhWhrxU/X
/kV1OU7cCXFIHrB0lUiA0KhmtyNg8fg3yHq60WqGMCStm4inO5apxsnL41rA6Ohh
+6JyU7CO5MScNKp3gLcleIje0tgahFhnpaBPLj/yhyANUHrRDo94k9XFCq3XiUd4
OjRq8hBz2L+fy936cZYKqqfZsoTHU6en0f3XX8qrv8cpLh7YbXogp6bxMTyR/3AO
orC7wsKxmq8C9xP/Cyis3ki1Tn/3M8NUx7UK9kVmZr8j1JW6rRis17fZb1NRF2fK
RlhQLoa6/HcyJ25nTDd4/b9n5a9bLiC7ci/Nbu+ks5j4kYsCwEno/Ua8QYaefCt/
xHvgkAdmPvXMDO1s0neAXmj0NUw8NARAFuRtFUcEkC7JB9yeRzaRZ/cdnXWk5KKJ
jXxibT5G00FvYW++F4ughxVkvw2y19cTPO8sDvRP+M5CrVVvRU4Ogo/UeYSvKfZP
LFoNTS0vrKtguezVwXNgz5dOeovTVBgaspQwITzXn2j/Tr+wLWO+qlVNXdufDNE1
Coi09ICgARHbYHPUa8sF/n52xCIH7vTtZz7hH6IvXEVC0QG3J1b78zy4edwughiY
TQNqzBRlZEq+pyivglTJYomu7Uxl7c3GxZrzO4xgYjv5/nyytHZ5hdtoMzUtbsja
+fU4HsGwLatBTWpHr4MI7LIQOs8ko6SQeSS+EpsLdtRi1YnxQ8kvwuaWTqrkdHat
Ad8njILR+f7Zj2NvhCLEfzouaHbfvoKIdsosCs+aT/OgPuw7X496vbVvULGpagSz
FLKQOIl/Ol2PlXWsy1QC69eKd+qjG9ZDHHT90FbX10Z8S4ovXVoN0hfYY2TXE7V6
e2ELjsqynagIiM02ipJqBF5q2/0FP/K9leCAZkXLTBAdlVl58XJTW2H5NsBS8Xlc
dKq2zerbQwNp2EQdpNeBuKk4qu7nixKX60hmoT5spLU2m06HmSbygcpW+hu/zlcl
r2/hUL0wnM0rAEeJTfZ5oI6+IBlDQuqRaY92mSS9xOBf3uvDq06d6XzH0LpZrF3S
IgjIytGCpmaLrB0Ro/tTHEKV7r1WIqiFXjqbe9iqRqlWDChi3evuyTyQYZsgJAwF
S42VZHysBiYyytAhS0IeNoLvuQAXxWLL3jDYcbYT5coktIyVREP5Dq1lv4MG9JmK
X1Sb5TOT3ul6oiSgV22RGCt9AsR5e9n+6QtXv3OwuHCP5eWJHdKNfeyc6VfaneG4
blawpwpBH9xJzfOHVZDMA3pq8/WoUoMuFKEhIELY5GXa3EzUTRKGb9tpSAELDLJC
kZ0X+5pw69Omx4IkhtRlvGC8aTaUFZfVngiQRAo/loeEdr7vPUzf18PCW7HO49Am
/I5Dyodq/uL2d2PHHasJdKHW2ETtTYFwX2jisliaN/LbkxYDkdE34ChI06D0tS7r
2FHzSJvDxVLiw0qYYMyhXtN6IOgDxP1t1TIqDlGm9P2QpVSC+JowkHtsUxMp0mJ2
ypebq160jLkiKuKtkoPFYsVWTnif8E1lxl9WnR5IWMHCgDR4WTItFFkgVylE5PFA
pvtrSh/Mg4gACG2DgtYu1gAsxwLECk8N9sqGQ/5nNIJ9U5cF1c6QPibwRdUa50fG
IzERKzWIHgCrP25aUyr4pBElfPA39R5wVeJUDxP83qmMfblue+CjmMVaqW2X70ls
5pglD/nXdec8h7Vu99cvWj2HVdRHwzFTbV7++oC28X+Mnm2zxEcEWC3pzonBp5eq
HtZOugnis1ll3y2TRNdnTQRYoAKqPl1nZMVHOUKKtdl9zPTtH45XosS2IMFYKst5
tVeYG9lucelflXm0Dzsa/x9eFLwypyQzSZcO6e+iaORbrFRLwS34FDZngj3Wd6pR
OwN+z/pq3BKHYKw3GKMs9MgQUowTVYnRZYhydNqgbC7MkYqoGeuWs7IVhzhp8Tar
E8F/sJ7C0TyiiwGHb89ikzsIWzZeLFrHBFUXQiVTyMvZDFz16z04S5QujABNjFCb
lwDsJCJPmCPV08hZ2q3t81YurMCxanNpP5vJ1PZDWNINWxBV4qSjU3cr1IOVSADA
hVqMJruiz4TH7vrXzCBIbNTN/mhxalYE0n6P1Ya5eifZ5hohqkHLW9tnyiNqdkYT
nt0T4TNhw6NlebH9RgWMHzGS2tbsdxV5oCH743zm3gBafTHBgrVj1WdFe7B8B8sL
xpNPVY4ArZQ/uiF0BKLE/8zLREXla2XHlZbgIpZgrR2gj/GCoVSkM/V2RHWaM/vc
F6TQ7qQk4bZLfCPCKOh6WXNOiIdVeKeHbR58wcBz6Ii2rKTjo+WX+yY3QoZYQn2x
CTl6iv4mjLocDG9fvypHofatfwDX7RYF9TaJW8Y424DXHeGG/0e9kH2LQcjcuSm1
d6kjSWC545E6EcMJIQHgMqHEtLwnrSSkPlCEWnPfBVUFhIDXkGqPa2415TfKxjkd
k0vWA29mAodu3VC0d6dW0nl03HGK5DuWsAUb5EyIeqBUBqrQvoGnb8JcPQrNR2ml
l1YgLE6hRazgfiF6ttChWVBZMZa9EnA3nXIdtqnswye0LE3aVzB9oTy+fC8wJGO9
TLAq/kHfJXvPHEIwAsC9axV0D2M9OSWamTG9Dkada91riU98GtzAyFpesUDLIBWq
U14GgvwNOf905+JhgTKqBpxUfuzcEtaUvFLAHc2iYp/qgWE1fUhG92ICX5HSkE/5
9j+3UsBhCbAT9RGLVjs9zbA36sjEv4oYRjKY9BLWYo4F2vVn30dP5CRLNBrf8zA/
JIkQegHWjYvDxxkzI4xIs6sHCWZFWWoqA12okR1mN8AN5+bUXsMSDaXwbIZmgB0Y
qAm5ePDk2y3Ra00xNo/JBGNiDGdOvO1M5QlUlGuVoj4wj+VX5VgcjiYFOJlEOS+W
74a1BPBUjZJq47eTZDfFkHKHYwI17ZFjVdst/7/qgTOmuFcWGN3SZBcXqCBKSmhZ
fcBuC2i4CRy/wwDAJ8qeyCZSGXgr+PXCmHYTp0ZuxXlgQl298SXvIhzDikNazU79
TXjuRjtOhuRu8wnjmZAqxCeff6yzW5YkpnPW3XPnXUCSRvVk0n3UX0ZLmhXTQFbc
3RLgPuZMXc71x7G9s4bhZATsU0P499Pa40kPtBEuJsSThnXtXql6TBRWxxPwwHKZ
FRSlAXv+Yy4oi+x/jhQN38brZ4onahMnWfUEMSR2EF6I/pEJCD/t0DYsYfxe9J6v
tUK2ZQ75PiWZDYV/X/oW1P40YLhJ9kVJWTZjz1uYhCXymQYyih2XZx9WYcBF2c9Q
h/BwpzCBxtrlBzVlPPZ6NGGLJqJeqaj1nDwESD/vxb9FlM/jb5rbzSL3naD8dw/+
RM9VMY3aNYOXh5tYSlQR9Qx/WzpdeHgWN/dLdmfu+SiSg40ITpqb20QP18jO0/7v
IaiXoA9k5aghkBMLDHyuBh8PAI/ylAfOa5hW9YBopQuZtV2M4W2EHvGc5gbxkvXY
e8DXojhHrZRNQvekNCDZhwG5vQRHJ1DW1llD7EiQH3LwhHU0rylTzlNBRqVZEb6H
a+p9rOWJbS8xnVY8zv4+hs5TYoaQyzg/BNMPeAU1XmfiDZ01UOBI+1kXVemtJ6kF
D2dJsTvHwJSQtfNfBqqim0JNlO7+w3Ys8xNB1+oSMc8xKwRw83wxsjhkN6IuuNMn
v4FMl6N2IlFqMGPNxf2eu1cwj598wygIFj1+7sdlFzwkuJN2geAOAV3c7MnhQkgM
GoEtb7loW+vgfN/xpWAIeAT9KIDTdW2SYlSaSYNP1PZo7NNH4/drQ2bjSLYW0+NE
p+myGyUIIHrZh3ZIlNCuayCN8En/jMx/ECPcfS2aleNA1BHpgBIMOUYOpWqQUGd+
vVCBiOEhZAX6bWAyyT9g22hOhQnpAsdRJmHVqaJktYjdux7AjjpjSRyF0gX8KJB1
U6uOXrdwIrbn4IkW3Q/5e3G23ZVYV6zRt2s1wAo5nYs35aOAtslkfIKV6I7ycVwR
r6igKPICVNvSivOa8B9hgeU0f4KUl8lKJhQn7F6X52B2XcBV/lIyLcpSSwXJj84I
usDg+ic54FvUDeROXKPUzxUd9Hl0xyRjqYOkxFNbuLKoDuzqywG/DwrXzpkE3cyy
NzVarG4Zi9R0tSDlV5JbpQRYZFyld8tfjGiJQDMXWbSO1o06o0FnelwI7adY8Pem
qdrAGKf5/gq2s4UzIaSFg0dcO/ODK6gzoYV0qdnBjpgMbrSVvK4jki/xDbVmRNYh
WPO5Fpy/vieq2G73i2pQpBgTHAytXUXrBrCjP1VIahnWoh7K/AYkl/rGSSgwK6T/
Q707DR8BRrwhjYKf8aGWAjNK5h7SGg72mpNWBYdc8G2AYu6qVBvg19HJW2lrkdNo
3jl1r40VdJs5254v7FdT0fk1UHs42yc/Bo6kOkS+I2BGA9HNEHrLbrTVoy3oEnCd
XUBRqXJ6UnoX0PIRXNU8NnChTuEz1kFsuuvcZMNAWw4W1AtR9HlwJ3GxKh/QBrh2
MRLLwbamtPPFiJBv2m9V8cg7RY54ZmB3blowFVh101+CYGeur6m0mWwwm1JSKn0A
jS62E6xRlkBJWnjOVRqx2TwsraCGQsERBs4Snp9p6llIZG9OXWHAgHiMEX5zoafO
BKtWv+o0kxeZiLV1JyzDKDj4MpPymP69e+QvYuXhYiUFs3KQpEw1QN9tkWKKj3qB
5frp1B1FKeESKei+4cfI/jEr4fhxLNeYYChuAARuNQSMCWYtgkKLv9UWEja4S3dT
PI0zrya8XPrwWcj3gdpPt1hy5eLMGYWyCSYnFN5W8OCcm3QeTU6UAmRErM5HhZQ6
334wUXfpVzlZZ8SoOOe4B2B/5vP8lojM/f2CF8vl+qVCxJhmpVoZkZygprWzWFMW
L7fIVEXEFbU4/IjazDfb4eEldx5Ye2o3hFPqO+6F4lHVlrisbInaYTQvb8Vcgpkm
rfUMdCw81C9ZsnMRC9+VXVT+XKrA4Mn4Bx2KXiJfqM/jg9yTOHhtwIM7jpMj7l2q
4c+n8WGDemQwjPuRUcZlCvfJYjGCgN5+osOb/xTPJlXtmnrO6NSZTRRgPEhOQiZQ
kazHmMNrQcbRhuQNgdtIT+RKrT+XdDvUDXRceSaToE1aLcqeOoLmRV+LzMUVXHti
QI0huVta3F8Yh2fi+te0NEiPp6Q4Iann9/9VpfDN0AYKTkmHPGBb91N/V1oLKdlJ
JxhWKyDoefQljK6nptcDcBfl5tpIYc0hwYQP/DszWsnyJ10/em4wszamE9RanPYz
4nEk5lyToRWLQ6jFmA1/rlR9Ry9t1T/+4yJYw+DbYHTFD3o0mbNOoCwgPu5ZaIZR
Utglr0tXckUaPeqnpAqMQ8QHJ4T2hPE9A2zfkBg1JrrsPT4hGzA/i3JVZ/9dcdPR
h5NrlFEYoqx+5LJoRDWENRtIKlhac0+U6OOxdgMdA16tImq0RUnuA8+wPfeYl1rn
U0Jgiwx2g7TN2bvSW1GqmnoIdYKme/G4xQ2IftGPBNXVCgcFDGkteApRzelPwueD
Y0TDhU/vh0v5+q9g53jPbyqJrhxDfqf2glP3vC3Pw5owZXmK+i2/1iBhCul2RajL
+z9XjVQK9SUpp05GjzDcac0MmBmSDZd53f0R8VZWf37Te+LiKKO9+8ApomFEiSny
7NvVuloNWHdmUnjHzmVOmQnRPI8HXNK5u6jS11FQLj3A5F2J9xHbRh80mOe9Y+2F
hbyuEcHv/mik8nxTyMg1kqGEs5NaaoQfQ9lACoAQnhyY0xKIXGz5eztiAtK2XyXf
d2qMT4JVZC4G0cs5ggRO1MGZa2atI2zzXkBvRFurBvP/1AM2L3ttEJRqCIL6cc2c
jIrWREbZujl3yd9RQRAKaqcAJseULl5CPJcUwQ4Ovlen62dDgLImwJuXKJ65BcTQ
vg8fyXfoENDMzCJ46HfxygSexPslkCqrsU7j7bh+KmCwFekiRDmXhPeCk+Jp9Wn4
xaiuBG7XEWvERHW9T7h5G9dIUimZBlThU9KuEE1xbEzKUzqXCLo3O8zMtphyz8FY
f5fagWJRJftRDIFqPN4/NEIorg3x/pyIbMYaSqHcs3WuBbR8u9vvkJwvK5b0SiuN
+vQzyDFH1pFUHRja51Kie9WJDTpbyTgkDcBuBYIn3NAQW4Q6U7TwgzYONUSgUbDB
fT/hmmZMh5tLtSLeeorRU6utX5d2MQbx4OY8CpKySKKGBji2DvTg3yFrHJJJS1n4
czboqrWwrQaL4ccr+lcZORJkRrnNdAZYBCaW8augjwpHhFeeTNuL0HmSn68J8/a1
QyEfDhkIGuuEazm/6cFdxWW4z5mOYZZnW/+c9iyFeFhFChwa4lqoohuOGr8C5ktt
uC49vek5LFPOg2ZqeDcVccqjV7AQUnWet8npSJKcn1CPgkWJgG8yK3UPEU8ehsb4
n7owwKQFNoAZkTV1sQnPb3SG11o9R16zF2JtR2BmwWBBVW96KwENuETIAQH8on8r
0GG0EjUeUsZfDl9DTWZvLkdIeq2Bwq01FQx19m2GgcXMxHLSLJZ5XJGPUVlwy6GD
s5qCVBNwkT1MsvRI2fcg7OyLoRqzN+do9YtrLQ8oKl8TmN4qGm8kir2GWryAVq5v
cWxrj56HHONTMlhs/5ToCydbA6UvUlg31505QpHNbAFg7BUkvVgdyDcxkjWV90VO
eT6L+LKyiU3CtO2mSVMW6uOYnEY0zobUQ+U4dxsVp+cIn3mU+I1H03dJkH89iidF
xQseNCxQ+XnEQ9IBE0y8tlCs9mdqqxKyat8qE11pssgZ07PSc46P6iVdIuDWKkyI
IeAheRlfB4eXVSQfPAnim+zojaRTBrmQDscrOIsjDXvhdRbANyAyh6XMuwbQMoL4
4JZy3BfqLtGZcS+ZWcsfi8QRkyp6mE8qpIKKYF9Ogsl0Gm7/B38eYF/EX4dwd3HJ
+D1bu1kUUq5j1PduKHBhCKvfi5tHtMzoXkAiR4QZX3oN33avmzVCPAOxcQWyHVLi
/HGRfuWeRfq9iuBVmZcq43x499DQFDqEoTt1Gg1cdyX3rXhrzvmRU6YSUF+lNYaP
4nVZxcgIQCdqQbSqhjgkWe1GPJSpmLPLsWounNS1j2jZImR6AexkOSsxXlZP/L79
WdgQ9NV9a/5g3B84MrvQOoru+aLZ9Z41MoxQWh6s7R18Onqhf35dPnD1vhHeVldK
9Zs6tScoNV34tECs4TbT0ulxvvNPQa+dB9hMf5mpwN2BBy/9RaabrWEi1Efdu2IM
0Z8wRWgurRae1q4DNak8ahwcGJTiPZ+ge8fjxpnqjybSvtOgC7EadA1H60CGTyAT
LIas1RUcTWUeYEwHO5doaRDv8lSGvsV4EXzHR2HntyYA0gLgCbFeqKfv/SokqDDy
QJXDsjH+9hOvGcU1tNmabje9EN8fkFQo0DIkboSkOYbM2DHl7//iMiV8TpJK4Aeu
hBCC+igHa1a10f5Y7ugC4I6uZpUVWnfQ+f7UPBrblQRGEugnylkFJ4+EVxzy4B5x
jXnIOImIVbHJxrbh462fMF6eOIrHIoCZCp/H+KWnow63vMrL7oQfOSs7iUJmPxpV
I/Pnb5q6Mue8vPHTxznuTMefqTxF57k9/H/QdvT0gooaOh3X8UElbzPJLJM0C0Jx
e8ziQFYgtLdEQcsbaW7aQwz9uu8aITux++nyWOUeXwFMP1UjdR3KOfXlHI/SJQc1
KpnVLIP7iANE/i5TE/hfyqXOOewlB3XCEDIOTYjML+AeYvL4OKV/H4pBAd80NHNC
VRcQ24jMdVDXvaFso3kAvkLGMyVPU6nt8VVhxId72T4CxlU8J42buN9D574XItyN
xYFzJIhjfgRRxrtRM+pIC4awceqD7nF93QGRX4jb74lLLsWFtZmExEsRY9zyAKT+
mCJ9QJKobhHRBcBX67R8C3QfFyNiN/vmjl6Fe/9VR1VE6VuL6IPF7qZrrVHW3tgC
NFpRp4xfvmyjRmMWJu3DBD226OFiBfTRcxNGJJ2W18Z0BBgkJXS4Ky6ijDS4PY3G
BBGphCIC9ewRYX0TnPkT0lAUrC6bgDivBqhJPq4PMq9uNvIYXzL2yLtW/YgXY8Cu
GV96FQkl0EolmvfGdm7+10WN6NaGKAQ34oqYimTtzzEZ9TOeZyOsLm4soR0HeBqg
SsKhUsJ19EvJ4sZbvBF5okvtOHFDDB9Gz8MRwCJkOQ+cFfi49gCWKVn+9eA2i75T
d8cV9AOWhxjiJmV0ttoSJmsGYMdiAl+3AK9PvRO5K5i0IX5CMsQeYp139ovEqRYK
Q9/s6VXPQ3tRejq9+cyUmbjmVcVKF89Wam7+W08lb9SjUgmUOkpbhC1UA4qjVMKH
5bbWfchFk5XobTf1R2EP7X7RyTbsBkT5Ft6Cbr5P7F7VnA1ITXs6/76VlKMFz1Cl
QjJaSw5MgA7kq3SFJxMNLDII+RIdWtpdcFvynQhYXwJ5NbUhgJPhuMQNuSQb3wrt
a8mYWy5/6/aFW0ztonuKNv84cFRWIy1724m4CGyBUNw4CgkPrZFwerta93IbykSD
SJ8Z81Ft0qKx+UBi+KNP64SZX9w9/rpbTosbzWqgKMprmOWY6yVz5JsY5nfWSk1+
jlRdyt2gqfgJ8F3hoUqxTtvGZCslnWIl+SgOML8iiHDV5onBoDCjVdI7/ZCPuxie
kiw3cdDEtvFWYOB5720w3VZ+iT7ez5K/EOwprmWSKJMj9gCZHIL4kJDHAjLtFrBi
bDQmZuL6t442z2MhZ3jsHp3oamJbOVYLLZSzamEuaGCnaOzBN6g4RPUYnXDdetn0
Ua38YLnJLeKOAnZlwrGDt2axzo9gtdb3ASDqT44K8s3ybdNoKW6nA1WoeqGgDISa
MGtjC0/EDvHp/L7xMBEEAyGvRhGIWSBnGBlUOcOwggmoUURGTUX3smTmG9MEsHH2
/C5ufNNfUNH8BH/2/3V+u+HK9BsfBembjHywl+tVqWOREWUKEm3GGXmOmFse1/x+
h+xm747ZVmiOSSD+hzBsNGoQ4hgq4Q1FvzpNNr4xYzL/9Ggzk3RSxBQHWd0xoAp9
rei8dgqS/Dx2D5xPqmsFICx2QUThoXQwk55tNnGWoF7/m9siNwDWTpDMBKwNlCY8
zhHTkWfBD1if7U490oCF5JRIi4CXb5fcWXcUn+Sk+PhWDTe7ypovdsMTl6vLe8sp
uCtrl87VtSde03aUuandTLBeSLJU/powFCK8T7FJswnZbDEOaqUtCmBTIT4jpe5E
9emQTSye7Gcd7O3rb5dH2Kn59sA2xzZp0QdE1Ejp7dGpL24a8Ks+/EEa5xhBAvLO
CP9yosXzTOr6qY7d2tLgHfHxm1vH7MYgR5LiMW4/WyItY3ppXo2rU+eOhUEsTSP/
e1RnTIR1bdUmyqNsbhqU/nOH6AzrqgNOisaFPEcUjeeJljov97tOZ4ZXTwQq/Kcp
BOxRs4jnVDtDbCdk8EEwkbdZwhDx32zfEw2DkAdBwCS02d8z3h5f9U4j9pvVMywM
avsb3EBhLU6Zy9av95NT2KQHpyPFjOkGU45GhCNw/FfrteUrv/vfXax9d4Av3uNI
ktnNnLpquLIc2MMODX8pKvQhLgEE389QTFJcIQcxeiTMwON/tksHYnYXHnFcRDt8
1PtCi/Opt2OOlJhZfzDhgSQkZLk+qgzlAPN4Rea3asKoYZ5dlfX3Bgyp3ZfP2PIW
RRChD9gajHUS0o1e4/CehmN1W9oVEqgntRfAkJo0U5l9vYxeihDz7SnstukExxYw
H2DvzTYCbuYz7MKEnsXKi64SmWu2ybWJSQmARpcoLbeJ+Tp4O1MSp6tN2IKCNP2+
I45Qt+s0mWRseE3D7PWdHFQlEF0zfiSRYOzC/NAY8nQatCZ9O0Dt4a05dTKjzwm5
XUFlleSoBFNkoe35Dt5YeReY9ztcBzVbhLa4BIbNrH+lwHa//qfeQUXCGI1XIHgM
+dFY/lDq5CSd3umZLKg/gyn5MWc5f+vDt5s5i2SvoSLVEOD2X0CddGb6m5pUfOzr
CocNgmuk2QP8He6S8AkaE7a+NsVxoswSHE/0YNK+G0Py10SMcBg0nBxaZjA0T35M
sxAwj9yrfSjC+0GyKT0zMedB0UqwrjP/slXRmNvPXvCfIib1tiThwhUKy3je2Q8d
kB/7HoyjZzYWz7hfiblCy6Agk3djdrIQdmkYi1H7NfbBM7NNvQTLGJRPtkDe5JGW
yVunYQMdwXl37I/8G4sSVFa7q3ga2p5KJhmO0N8If3t2t2XY+ZvKyV2De+EwvRhz
zImPo+9l/RktG1gFYGSvLSio2YCwjVcnc5q0sWgBs0AjqfU/bnfsOAG5FKWMJU61
zDg0fur7SLHaphf3KxZOaFcaAvEWNM0Tj9oSONbBb2XYVtslkYZwlJaupJ27Y/2o
+eiLuCSs2wh+wvJwdM3IiYNm8HBLEM0wJX/TIXN/uO2/4OhYFjfn7Nlqi+gqKIek
jvHAGdW+EiqVsigE3ptyTHy4qEElp1XpXa6hUQ8pFUJuMMsGtD6yeD0/HOdN4aLN
dLfsNaQ6npGBJLuTvw9xuiashE970c/VsGIWf5TvpFCVBF9uCL2fOFAgL4D6dva1
ZrY30BQirlRDoNQ+nex+g+0ogrLDGMPJSXCsOZIlIzDHJFn5P52NYxTOgfbzuwxY
ysQe/wRMsTLSozT+duAZB6Id7vbBFeVdJ+zD4ZLb7Vvh/OkyUm7bmD86eRZv8r+8
tPb+cPFDLGDtJaC98FzVuy+Sei49LNj1cEA5o7a9RlmF20U1vGTT4O2bfT+eFS0Q
bLl1BGZkjHM7MznLuvVr6fDIF1tUre9xAQIdlzTTBjVpwKE2xamHNgfJe6EyCPdk
E/RCCOstBEObYcrkm98ZWN+aReDLWhwrWHkSEXpO8fRNpvg5D/n01JNR+VlFipWD
MPesnhrNRHn6GHwy6pYTBAMHwl4vmXfrF45rQjfHsSPmHv5ddt9/5dEsTrdoYTsP
OoOmtUnPGYG3TonozNiiN+04KRYlAU3qMQfyOo8PCBVNnwtKBkL+IfrUTaHzWHxO
D9bsR43GTqArJF1xgH+OonbFuxX6T2TVD+A8EGfTm0gFX/0rDcVkdeMlw65gFYK4
SfKLazIFnzO6o5JpOVOBuBdup7raSH7NSfT25UScDHYl+uDjvUv8pceRtlzCyI2P
G/gfDk6h7NjJcmwSdYcFShGhkS6qShNvOHul0YxYVkc3U5ep1XRKxNNGUM+F92UG
HdD46nweCrwzcJpsm0EhF1chfymOyKTbz6YGJV2LObJZ7vkpxM2pqvfKOUyfobbC
8mcYvGVsVBWWQlKzR71Eqco2j49I/XYYVquWOKkb46UXTzfI6YEMODTT0cSsYxMy
lSwNJpgwGyO3kOrIpY8czKZA956fJrAvLJV/6YTHvkV3wI8xG3phN+Nw2SDEXJd2
cTXQ/bSugC9nN8esvLym8UTHfCZzmcUVzasck0lPeSFsha4aWEBrzxXNw7IJmDRa
eZvI+XRw84/SC+U1QXJHDMNzNmmTz1I+9iDfvCK6cIwy2RcNbKpT7P3gQNDXDdsn
DZj0oIsMOupVsgL67oL3FFk/5K6tpsLHuTOgrXsHQB0/NRDD3/PvlJ6vI0tRada3
4CabSaOszgRZ+0fL6mrPHswt7t0D4zcWIT/fWQMiZNfU/5yELw2HxwK0AB7FGtEs
uhaibZcVwu/qqLi4wl4OxPO74/synmmkL179juU+iqpt61xftcSVE3Q3FSHwZZa7
x/4+0jajy3+dOAFXCZK9Voxa/b6ByoiZxT+jmtb74wwJomkHPTZ/hRLUDe2SvTUD
72HjyaodInyZtBxxqV6oRcZhGi1txtkI3ByveR4xCdMz0uMEZM4eU1Q8eZQbPC3T
iCcJQKrPbQ6t+pIk3zZ/EWwc+0wewW9hRYxlWU4Ng+JeBlF4WpE+V0gX2BIItPCd
VE0pXDP0ibu/HJJzkBjx5Bz7SPcDbJKvRomX6+McKPyCNDzXjee9IZx0AvtufA/X
PhXiFg74UHv/wW/5AKhJie4qeHuB0aOJnYYwZKezJW91VKt3Kg70PpyjCi/w63lJ
U/f6/ByVClhlzsXcnpSzVewgiOF5ToUtzc/PIjkRQmnMwrinH3JQJg/XiOS7ZP9N
sKA6lYjEr2r2PYRJI959vwAVYSzw5TBC4qn06NhUKJ329jmQrtmHqG4fsuxIwQDS
sXoplJa4zmx9R9j0Ujx4LThEdybszhYtRIvgLLATLeMlvQQsR0BUompmWB4obykW
tGDs+MUbX9kupwydro1NC7mrcWjcYRreRbSTfji0lXf8l8/cvD2u+PNt0UedW1NH
+E1a5IYBKvTmKmeFYqALgsuAoWpSkFBmRYNc8TfzLehfIm4Lbv3SGTduIoSC3hrX
FlefGoKIcelFPRZeRlUAhgPjOCMKGt4AKldGgWZMQJg8nhaTNzL0xu0jB+63rdAO
D6C8Mox6qRurCTtc8FTe+zYWxkM7UenbvVJZ/B4/lQt6WXpm9oOpQCZfHtCdwGSF
YWwXSKY/55SRw8neqkYqRkDBAg46MfPzMok7BhfEnCrJeQFxrJqPOkeP2yE9I4r2
M4rcSLa+5+1XCTYuJWd9NccBsUmwejYat+t22mUkGuyY+9BRjCV8xYJRLKxqo5ao
dF4wgivEQc40lKIZru+xnaIx8G9LCvb9sY2SBdRmuw2QlC51WnTbT89eQJTGutZb
40dM5LkJGxgLlf3rFUnk9INu0lQN1du/S/3DzVEhT1G/5VNb9HimiPuuBbuwfysJ
iFA/4L/ywfW3efXEOBXV9Q8mwxhmc7WN980d2K1AYfjemtzuPOqyBYOoMLeLd4Gz
bbDFv/87vU8N/jofiwQxaoJ6DM8YhhxJ2TZLeFUQf8zh8i8OE9Zrlz+BQxN+XLWm
TdoA9Sld9DtMrTxPmwue6C9ObK5/PfJu4+enMNLlX8lC6e0iCpydQN11XSlch/hQ
UeqLnLtDW0GwDjeICP5dfEAKTxexmauCrY1h9pjwUjPPOCpP4yfLKmouqAbhGLcS
Dos27jPcIaNO7qLff7yamhVm6GpnFvgLsxkKbRDhVtxMBIeXtUb0FNvG9ctOKicD
OpaqimQweGuf32CnXyTzTYQ4KCJEQJ2PTBj8ANT6+4CoCcOoeNa5qRJRoDc/SE8F
iKNHmF3Th18ySkxHO3zpkElCWd8abWfU2Sssp7qzJ57rShce0EUcHm96fgQjeDJh
7G0lq1oVDQ1Qk7v0vYAYp06csbtBHAHKkgoLW4f+A5p1QzgBSQJcP9OKgCMIDG5N
tXMpKc2Mu9NMcxsO17t8XoEQP4bAyf2WGQSrRngrV/QTHOue2ZAeSBWtj9hMYqIC
eZ3Ed+6k6vX36YfW3D2iLkvj25ZIocNzxhEh0CmgeaSKJBu5ZPbBScKUH9XnUsaA
aAVel8Xh3Yi2BXZeC6Q8Ctz9CqnnaLlzKC9iFpvr3I/1RBlD3+UHGU61L6DYP94w
R9QbgVxehnpEebrIKMkJIKi4vwVBYxjZaCseO9Ktr8ufrHgkgZUqSQ4Ze6ImJipe
Aw8B8Mb+YsXMt8b+MsYUJflTc0nAjszEp2ZfjjHrlkpA80/pG0uNf0zAc38RNo3H
Wfhi2kQlOrhyNfLYSC+3qWF+cWdTTbZHqo16ynb59G7b8qZpBPUpciF1M1ffFL90
rBIhZey/Y2L5LaBTlgXDWd4+M/MDzKwp8P+x+xIS9KcbkWQpK+JA7AoASdSjWvi2
Modmpll6FTU/Mu/zuvXUi4lW29hOuhxi9iNoCiqOym3N8bC8SviQfjpFUTUa2Skz
E6WbvbBSOoZxFCOoHk+Ae+Yoru8D00WnGcDUrBRXMqobc0x9W9dxG4Q53BkIGV7+
DOSyveiECCGSpPaUo9Jrp4+xlIdWQI/B57bG3EgwxwQ87GhOQQLJjsIw+v5uOBXQ
HE8IzYHmnrRBywqB4cQ0KFM19wOvi9d8VAB/BX0ShHeBxJ9zUhzM1FFO4ty8XnNV
2ZPK1aSw+5kWQqOcwbJP5ImDKWHnjYEbtO3vxWmc37wYUV17Jk13yCD4KTHSgPt+
ioM+M2Vky7TQNx5nZJiTJWGab2t822YTOHG/gCIxzZrPJSiZBfCo0ZZd6wbx5PFw
oWOzj9Q11ldAWWKyItFjgSvS/Hqn0dRi29NX25Kz0/u8aDOk+kXclC0GsxY7nWws
bD1vJZYKEJJ8G1rzHHoNNgSS3P8ExERj8OqIRZFOe/42tGN01swONSFN907bsT+b
8e666GZovNPiDABs99GWSyjZY8Kyn+v6LpjyeashmfYRc3NYQBRTCJZA1AQkLUfm
s0QwV0nqqcpLR67Ukf1P3Ar1f+P3gvcsQNu6TUvbetNkuKVUgRXlqFIJ1fa//SpT
K6AKqgIvlH+rFMCvYg0J6U2K1y44hOWiuXzHq21CuU8etxAzwNE2XQWxucuL60Cr
ngQp0zaXIzg1MwL4TGlLcZX9GID39+Ean+dFynImTEZgtiBWALtvfNsMn8pk3dLj
E6zU3rJiIX5kWz9OydodE9aHDzBwtGpPOSeF2j3/Ah3luEtu/mz3RUwb5OtXcnLO
TMGxcgQ7Dio539pmbEDNZsWThrbojtluLLcVmQ6LM4jwaiKZ5LcQJGow28TSStbN
F55NlPVKU+c0FsDAgDhk5Py6jr+QNO5o869WBuwN4T935n92vMkzBCY1JUIr+lWW
kQ2VwAfo7qZe9Fh0nbg2hF8iZduK6GYw75Oc+cDlENucSGM4/sNsRbHQS9HVy0YL
yWKntm0VlMfnmUOWa3a6ONZ6XhZTQC+UCVc0wFwC5G1NzXoof9ypV0CXpz9bdLd2
QLEa+o+KBZWfJvPgMEHyEAXtBk5UlaZVpTwWNqF7Y22OnqUKRiJdzYtduJjACeW1
KWzvgOijauPQCZm4M8Zy9Ai3I7gOjyMr6B1QA24oGSqtoPDrvRI/1UU84p/M4J+F
idQxIwebL37xGqqMGrpH30prwvYp2h1+tt4aCN+s1AIUnaD09NarPnc6w42hxNVl
K2krHle1CmhVaxTHu3Jty95InV0spHxjH3Jp9oRNO5gZiFegr1mMtmSCku+HRPEP
fCQ8gXr7dODCQlRh3GPpNSyH4zM3ivY/H1nwZBSQs4LoCutRKgKlMJLF3JaqGtXd
hG2+pUjAf2M8/0QH+tm2r4LnKcOWEorV/HGFN8Tec4skxFr960zR5xkZwgAqCyZ4
tbiQ6p1IFnV2Fqt2pSSg/fnp0DADfeGrbCltpl698iQFGm7z7z+lUSwoUSWlSKIw
tGIOhRU23GOz/AUqNsbVxNt9lFaJCDoqhWam/Gok002ATXXfoPqxcJiWvxL65auc
te/oNIDC+OnniZfyigSn1z7WT4jPCRNnKLKIr/JvtbUjhdSlz83piAORaJ3atGjR
lWEhwDfyknKuUocTLfcNIPKykgB7vZX7Mmewxx9AXgup3vhWkHImUHFASqLszSFR
6qhTKM1DM0nIL44Mqg6wQVo/nGlY4B3XLF1MDG1S0edS/mUpiWxIX3wqkNQ4zxd7
GNnXF/FtewQifObn8kf3B2K8wbD0KF8C1QBWK8T2I3QhZ1uwSPzHl463ayDh9ZQE
QNKkWsmarpxoA2ubl+VPle9quD2B0QJf8nBKVdVGlZ2mwS/d2clIE4MeEf5AKWXn
w4BhfaTLHrPlcCdvPEaqBF+gxEvdgPRtu5YcFPvX736+qluPwFw3Vh2n2exE2ks3
/iDtaLjVc5PELeEHply8TpQsYbkPP6sEDCCC90WtDGLVsSdzlpsSpERhDSyVFtxa
DP8cNjN7cVla+VxdaE2dFstaqlRbJ1khf55fHmQuAZYPwnF4kyc6cuIQ8CmewHvd
b7fbhqiA27ORdd+J8zCPNFbFgsA6pNx5uFglTY+e7ywx3onwr7Yj69nfP4apZwxa
bXrcLzaKE3OPhKkqQ6GzTGD50HTxES9r0l2Bmztb/MRsmFgwuORLsJ+OXlQnCFcq
cQJK+Fz3QXl8AfpNptXG5eUc0WCJ2vJ+cFMhvTDamPCGAwvLCdQTtRZmRantyLNX
FJ4BzQY8ZRNjAHBAOWTBfEXl8VWR97vVkw7JQkGV/WRKG8Oujanx/EiH3FL+4p37
S+0L+h6XXgmaoLuspb9wmrD5UOAaidwqgkemRR8rzOZnzTFG2oJUd+HiURjf29WW
4An69AehvdbafnPuB4TdWJc1/IdgMh66/HrAFa2MCwdzT0LwLmOeV1bu74mntD+o
ANJF9cB42n5l/Bfz1Y18e8lH/yoD6KrpMOyGmcDxv1PpyJgtIsHZtGN3z2yHTqpF
kHWPBSQNu6HbV0I1zU38a6L9P4KaKDSsH4L9ioLGvxGMXzxc31pV+twpVYI97JfH
PweykWqxUzu/+8sCo+XcIg==
`protect END_PROTECTED
