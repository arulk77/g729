`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkZZCKabl+GRgVvFnio3P6ktorljcQloErYryGDytdn1X
K51M4hSEYn2GtEnD5UfYOu7uj/nwv/v2HfRdRW1mO0NhfXSYHRKPygSuNsj5qQ2e
KhBplyfFVLoDcM1N1F5XUa3HSo2iEJWkfhwsNC71pAnKvowASVvdQ08qUfeOb0/5
2hHHXsNGBTPk0NTkxb1pomLNPZUS1IJBYM+uu1FWPrW3BIDNaphHcQJQAbTexpBH
eP8Ly5iBUWHFCHiaigqOvbOLnUpz6EgbIKrgCgEMB0Tr8gZ0SbMyY8kDYSbMgS6l
J/fbeK4gZTVn718buyG9m1TjiBlR6m4IEVHEBZ+iK2Q=
`protect END_PROTECTED
