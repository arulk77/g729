`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
6r7jZbNh5gqKsHgrZIPBqzlt02U93tggAsODocQdsyTci+ykl0LADbK8a6mGoKQs
qk98CVCl3gSapaKnNvFN/3jQfD2fZCaubY5fIIoeVLjtDjCcUcpqomJO4lisTAhA
ebNgHv9SILXLxXWZqY0ptJzNIZySea+Wlxc53nG6EctzZrzN4h8fmxbBL0bINzRw
/mP5PtHWnLvFCWs8U5L2EvR+raH+To1MSdjtFTi2+Mc=
`protect END_PROTECTED
