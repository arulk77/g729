`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
WzkPnEolwQM4IIVczoNyp+SuwOATPtJ3tH5n4oE/ejQ0Le8mwKh1ERE+5tmsCfjK
e6mVMNR3cGh3deTVVAPWBUnPXlO00f3idf+E9BDzBeWPA3FA/ZRiR1N4Z13Q8qyg
uluQhJb5lS5VMZr3byRSfugFaMQh2JhYcZOC222+HRaqaOPOw+t7tyN3A/FH/VkZ
QZXD8LztfDjBFDieHWxl/mVLw1RKtWo06vsL5adZvN3wRwUld4zbTxtsfRl2wsjX
6dSg9fE4x2YNc9WKYLMlP4A/zGSbpa0BZ1gbg6bqMaE=
`protect END_PROTECTED
