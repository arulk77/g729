`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/1EZ7aDk8xLLjp3Rw7zztzOON+os8bLV3y1sG1cXtVx
kQb31WR/pmLDtYb6PgyrVAEiKHvXSa+rIRdoqo93fRgnZHnU0/xUdzyUvdp5YAJk
RmZdlEKAWRZ994nfh7MAo6LSvBYxO6IW0fWYboP8+3JuwYzq4XubeIQBzei06b/t
sl+EMkndn0ent7w+CRqmsCvJEcHYJxarZr+UoOFsntgfxTKNSyJmPDemELI18YGA
m4YE8Qe4mSWnvZqnWl87loF8hVVebj6GraYFTF6W7Sqa7xZonTdr639J84Is53pt
gOyLukMGdzY2Kl2NXKTUKdMI/jynmaizMrtXLn2Ey+AwLt6VZ52bCASHPVHUTcgw
/LSv+6KXY+KE97dmMPNItQ==
`protect END_PROTECTED
