`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFuXURB91KlKSfkLBOlmDZawP+StMpHLgO7XBy8KFQ72
HKU/H4FthoygB3+oB6uKe6EiPDxkDHFEsUmrnonQ4+wkXXCz5/ujaV96buIbFgB0
OBXH3oOX/vT9mnFh9SEGY+YGAVW+u+CWhsAs/arBcEN4YLezGHgMNXWSK75VQlSm
by1PZaPGEDXo0z0W0XCeKAtNfJG0r+hdMXaY6x1t1WoN0iqflD5AGfSsCqWuAq3I
FG+NtKpP7OR5R8fTl5SGw4LSivT4zzL1DN5ctg5X5bM0zk2lvuZbFeXQZB+NDc4P
UmUBfYx9vNqJeAGV/6gh/zJLvhJ+aN7x97HfEJ/Juoc1YibnCbeYU6tgi+VFqGMX
pyDJuXLErSTpYzFSRyZP7vf7cYPEVCbIA5R1R8JIZftzu0t7Wi5FAPuB704Ul6It
ORwef0AgJ2QqDEd3FEqD4MqSXlTv/0tA47yqbzCmvOlMGz3VoYs31pWY7M9vvM0p
DQYivAlpIfoxgTLf8h65kqoW/8nQ+rLWS1BiZr/Aevd1ZPeYThy8eWRDuuH+sbSh
RVdW49ZAVYHIL3Rkz1bvx+IOTn14cFV6eeVD+LwzM3WnAtGnFUAlB/FtpmJhqZIr
yr289rtnpahIhISJIkQztrLnegWxc4F7CAVk9mRRpIk9b5TbedEykBoKM9H10EBy
`protect END_PROTECTED
