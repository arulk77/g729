`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3ON6twM0bRyFDJLDX3Tyeq0h06A5euAW6JnA79geTVhciyrN41scfb2y/BKfB7eu
5IwRII2xweJZ3RPQDbKdLsnwrBOHZwBaFQ9HoRyqWH27KrCU+WWOhICUoH8nok8i
K0GFCGHfJ1qIB7zfkxfyjnoX0CZ1AP+PdTrP6+lfvwK5drFnjKWkuiKtBkdtIB0B
g1w6tds5/wDbcc1whS9aCVHcYAdZC3F86hM9rXdsjvJpKvr/ac+TOCn0HXmhdJhT
26JKcOdKxaQK2z5ituluCnMiMIYJRg4M2fnVmUFy/a3VamuVbXIp7RvIZxr+OdZT
aCxQ8CAwjqGF7ufrmccLzvk+2EEghAwVBcnEgyb4kZEs53i+iRDLyFSVRE/12nQC
D5oU6E2TMzFvF3uDkz6SerBfIvcyWAOpZ3rhYZIyKzyv8/RzMKs2Ldlj1Kz9cSFi
0Y1h4mapW0UhQpWHnp0kRnrrNA/aGuicydbHjho8XDkK3XGfTswoCT096C3fi3+I
R1p3zS1DifKvwDguYbR2gZ5D+hywBXlLLjfXOFINVXF66Q7P3utgVBXinF7xHb/4
RGpu4DrMKPvUpg39h8+68dkLSCUlN2MfFzZSMKkCrufeAh3pMZvIT+Z0aTlE8DPU
b+pofS8gSx1e96Gw8iiKmvv7WIdCRmHp5b6ivIWw9LODHGvA2MRdGeNbMuEn2nfW
oGY5awu5gf254K6MJTfgUF3pSqzfbhh+SI4h+QwXh/DUYrZnYfJmIMhYsGyk+y4X
ZN+hKvo7ksq5YeapGu2Q5HDKvwqRPMupdrz/4UQWlc5+SB7wxxZ2FmzY6IfGLLbL
rUfhY8kQhIAFz8GSF8Pe6BSsofsp4wt8hsYUh8Ub+eViki0kglnMb3cZy876BqxC
WUfLDLfBqQDSQ74xaBbwSXyDTsi/VIHEAJbWJyB7/8jiqt1VZOIew465j02/5TqK
n1ZDo+15KJpOs/ftxCjei02zT6X3emIDS1PyqzDnWllgtKavtc/LdVklcGe5/7ho
/wS/lmaZhxPQsEJ0fP+Z+R1sGdjQ1HHlbSkCQr3zWSvPFU10L9VJ8KfI36ppT1U1
GfaTJz+fDlCO5xpv4UV7JFKYPPG3GWhRq1Ar3D+4316NVcrDj9qVFjssNwR/30zh
cX6jiRLLZCxdq+7WVA+VbGlPfM9yetQ1W2c2sclq7ByKSOVk8fOSu4AYWWvGJ5Zq
4u7X6ZWyQN7Z67Snxb4FH/zDCeKmXb4w7sAO1ISycnLmiXwQxEFG9LetZgcDtQiu
g9eYss6/lN/ne+6bdZihNFFkvdL7cm9d7HIwaQhJPqV1Q46+SgKlL5m0ZfWeJO9r
JYDvRUGvewIdGrPVCzhJd71NMxLnzaxEBob7LF3eDclHK2ey9sW++I1r32pJ0F2k
jtArw8luaqsdIp4gGYNo8F+0vI1xRCvlxdu4rkSDVJ6c5sI+2vSc3J+vWlTzdECA
jG4tr3XCJAXVSFJrO3nrD8aclKKYBikZbFEA1GehwG2x84iCDaGIYsDsjfPz1BF6
IYyi556hoyv9hYlH8ypW8Cc9GhwsdJNwHGWckfavbm1Jolj6XcTl914g9xnQpX0+
sFbA2C+Elpdq/nEstrfzKzz7KrEknsKH7EOlgxM9ehRF+nzgGzkDaCnkXUKd9Tdx
yIMNp3DwbIJI0z7eAZktb/GE0ACr4sR8HocwKMu7/0XbzqSqO0iiIlxSWowL9a5l
3by82X6Y/eG6QTdERGnaiVIPObcIK1CeiNcDssO0FYHiFL/1peJ/RvRpktytYdK3
Bp0Esz/ep2Biqe0+gluO+M4KrI518vel1BhqJcNB7X+mcny1efElWW9vq9x1iTVi
NkMfKGJfptvy5vxLtNY5uLl5dOQgXa+ZBPefHezpwPz3KBR3uBtFplnIGG3V1nWy
zAXnY4teyprKl07dT2aX5GyTxIhC9bMNPsNjMdY5VsweMJfLBo/83PK3roU8JYKw
i2HfnA/qt5lpP/188pfSZgCnWRXuF+8Uop9x9yAW/jzy59ZzdGPVRQt4UhWKZkY3
6rJnadBlNz3EQxD9VVkgEM6qVcxVwDYjrym6pOBVxy2dwGjcLboP8hNBl47rhFZH
YEopZIACDIK1vLwninMmN+vEetlFB1DK0fsWxa8aXynvLSEKs90PJiKmZWkhEBFv
OH91fwniwk9uw+6BJ74ICFvDVx7/5O20takjea5w6nM5TuxI0qXRyU+dVChy2usQ
nnX7rCpR4tFRtINwNFI7WurvwaS4zOjNmsD3p0PDaGjwCLQ5I1BahXkTWXGakpP5
VH2mU2C35F3/PMkXtpBT84RoYS/PJpsVeNPjIJNVu8kgbO1PlqFQLtZSvHARRLGo
J+JtyZarOa0KKKVry9zvX0b7KqEOeJC2sKdBf1jDaPk/oThtjCTnaXCNBig2V3sd
5AYcqOKtyUhPSwuCga7KGicx6hVkgvRSNih8CQLaeqOMLSjQDaw7iiP4u/8pywU6
dpg7oXzBZAUz0En6dlzZxB/RlH/n0LmuYSKRvnWtvgeA81joroz8A7yWuJvMnsur
rleOdzPCTErEx8oB/eFVVYNf3mpx1nBboZaDqm9TVp1s+JoKFUIujrg+xdn+pq0F
ZFq9WtwWM7OBSPP8ASfRzDUnD7H2Wft9aHSDslmj3JEd/IYZRSyKwIJTzHBZmnIY
+YvbuZwHVnPXP4wkRvrNOmlFj4EaaZkNG67XotyPJDulX7ukfU1U7RRf2cbSiVlu
MslkzW+CVn43FxiIIiF6oAm7c0KLCqtyXky59yfuxIyJbqRX/0uy+bcWBGl+CkD6
adJFfveH/y/Vma5lf8H8paRxuLfzHxpJsXK+kU0pCPLQZhO/N8kqw3JftLci1eOF
hVnZGgw4qfV0YWpFCw6j5xsTkm9DqILIuEDMdbUCka3wRdaZ3MXEC6wCnATFpJeO
vI54tz/Q5Ub8LWq9GusKXhCGSLNfOEv85pJ44Lfm42uFd3vDQyu6VLmvazdXuN6V
SsQ/DnAcs1aMS924vXKvV/0a3Z4/MYWYAoYTYCskUovB32ivsmLam3UQFhVjpz/v
MVQfAMsB7B08fCjZU4ARDBGdp7kEJ9+OUICAbQN4imyjbgxL7i+bCDCgP6AoS9Dz
GbV++npAClwOEwi4JIEJL/otkt18RMINxbGMNuLzMHBOXfXg/Aw1jOOQ2zaXmkpi
/fZSKua8FEMJZo8GD/mWbBZSC23Oor1YcDC5EimxLP5g9dp3+HAbzUye08sePgu8
l5Op4hT6DPL4THnsBr6mDfQzsUtiUEZWXoqwEf+WCm82CbQ82Pz3SHP586bO3Jy3
Fqbc3L4GG6KqoaP9VI+CissMnguVDUyufw4J4DcCuj6pm3Lh6E5UzZxk4nHDB8xo
tOd82lewOH+ZuY6d5JhOKTaydRT2QzttNMFUJuC3xXG1wVhOkgX2w4aU0tsocPFu
T/wTSd+z3zLoi9yqZs3m7ErL4hJ+9C4Q0j8He8XHdM+EV8UnY0HHB4P7B9+bJhN+
R9aRBo9vK/s+RExXB2/WuSbg63jhrW9ZZOPXsHWSLgNbyO3/Se23jy5/BfAphw9b
nfjEkAxVEaXPcLK/+s6DtqHRQtvsCmq67nlbj2hippII4Iyn7hTBCbd+Hwdw8eLj
Mnie2/YLfjf16svEs5l+XJaaqxNMZm0PDKXOT9wrBZdsH0hvqp0zgOM/A2S7s2uW
Q+P2ExnbWr5tnbu3Cn/nlw29Ou7B1DdS71jgjXoxSrBtZk0YAJWea6QQxiX599rU
9bu8yc4OegN4Z8AcmOJ4WdVxOfdC2ccKNIn9YMRzSmaLR3h0ww0ThFvak2+vKLiL
HgUgcz7K3pSbIa2D5zXiqS21z7AynB7Q8fLAzYeDUg5Iu99AWm8v+vQL78vNLjT5
+ZK/Xdo/BjjEhSBcetbcO3ZDCSWBsOm9htis3zPrDzzJwn/tqNytbJQ6J8PCnb2K
nj52eq1zyX/aSlx7vCCGSDergDXBkxJE+gaw2pZWAfVoY/ApyXF34tRbjzZ57m1a
Z+Krg7TzMDweMLDSI/k16pphQAvPVHFpw86qlXxYrzFkusgFKMaZp1uHoYE8123G
MI66iqos766NANdCFEVm+/vv2yskqNTBC8CYj6NkeiASx5XM6wsbujCjKAaqtnkV
lAibMUSUwQ8UkwqcOi18j7oTjFk+23OTALDc5aLZ/c8Pduo0r0LWH1IQR6UDzxZW
YO6tSnFNqt54tqIG9CaAUBKmKOAqxmG9ezN6orIJfE2APhboh5ZtcSY5olLVSUq3
Vau0bj1hvyKwujAAZMI7NYZj258ROilnJv47S5T3k4c/zW43OWdchAezgJQmVqS3
ngtMRBGWImeIOjUtlqnPQFFK+ZQPcLD6ZN141a/6MJVAkQVxLWMjg+XBhzVW2/8B
O5YadsDDADnLMSLHl3OaOWIcRsfhQtbK27QJufaq15gQBvD5YlVRYzkAPXYCq3s+
0kjwS1CKJBh1PTr2EvKYIJ+aCqAmgQdQZJ5u1ciq8YtFKIleWqh6G8G2J9V9zDhF
S+NEVJJ8lkE1Xowr5kzxV1tpaPN5sTPJO8Gfs/AFY5+zoun2Ckx5BcJ+KDwwQ/fS
tdqo4e1SppALicjR9oqqL8Qu+6uLZ8uXFprnNA5iti5qb3gi3/0iQlK0Ztl4F+fb
GWYy4Seo1lw+qCuPCVIORWdct3ktB2+K0OplqCryoxr2SeDlRVDBZ1Oh20VSC6YA
crv4UTZhKj3R0zP/fj61KGDkZkq99jrFoQG4AQ2fUGs7EIl6jWzJ5zWjTxky5/8A
JLSOXNy8hO+K2YEKOW+vaVwVdWXtZoTt6CJI82jpDpExcoLVVqzD8FYGkbM35DV8
pZt7DkybgID4tunTx6h0KcJA2doHJ5hvLqQRkZ+AcqM4SDzEPLfcKnFPMHBDqQFV
oME6nmO/3W+f6R35wzP2soaubRsIQf23kOxwd8Z6MZDHgszpwcmnMRvzCJPzBR39
AlnmniD7ulfX5c5RnEZE20xoQ++9jutlCuU/zR+9tocChibJnXQk282JvxJMetjs
uSWcpEvu51d9El+rmZylIXjGaN+WEazqpCogLXsbdZJIchu7hFtukKeowxD86HjD
bI/NurmE0ZibETU+emir8c8kfCpFlMkW0oSZjG/xwstg/kpzO02/vStjDP7Cjq5N
o63ecbOs9YhCydbV+JnVO1MZugiiTPfnQKc8NzXgEI5rpA7oUkuu5G4T+yu4eCPu
CcN97Z3q4et4GW89aH1Tjr4GJ6yhffm92aOIfq98BFySdrKJL494lLLPcD8GFaHy
D82QoEP+GRGwECu+hwA4bGdpDqDaFT5cOpRTJnxB+AJI6rX8MW/0b09KX+ih/sQW
CS3qh8aEL1ZUZloALgMzaWVNN5JlmtMxtAJh7lqJ1npkpwdSWSFXpYeiBoe5Cnzo
rPc3cEMqcsNmQuEqrblK7b4fVXQPFxjtEh29uYTCgfSGyJYlEtP7Jpv7tielxY7N
rNEU08L5cd4RYQXF7UyNTr1ebg2/yOGUXH5KoGy/KEFTzdbQ72A4WWrT57STnvQw
qs9dXx22nBYnrB5/KIcG35t/LCgN8sKxMk6HDT2H9MJd9fCsHWg3fu/s/Tjl8shJ
UIfhLNxLaQBgXWyzI/RmoCTEOtNxf/nPKPgbUZdaUs92rglz2Gp8YgKgR7SG8BXs
m4kEgO+iS5DmOJ9rKUG5/05lsQroqMOUxYEIEjpWu7pyA9xdr1TCtAeRqnuWGCr6
zxrCIP7blgczOZLB25pxCBMNuLIWGMr2KWJ7XkyAFswcHrcb8/5T+pI84gKXN4Rd
y+faS23pmtzJVN0Ek175XKx18NQeI7GJnO8nrHPpiUX9ST5zom0BbbLpKhoGhIEN
ibCcgSRGiS6zITkg4SeU2clLspI3q2vqK1P7Jp6OX8DwKMIU8ZAX9oQYyACkZlBT
B1MeNsU0slcDOxM2vOnk5KhnTc50hZZ9Pad0gscOwLBooB/kO0jH3JZXXCLCI5vf
ht5VTtCazhodulBoY+fJfokDaN9OxKyiZXIThTBfnlTZdV0IbXRZV/+LMwmH1H+H
FZXT3gtoh9R8JAoSENOMyiR2U3GEyLLA/OwhSALGr5on1nIac0JNhIESo4yKR+BA
OzayCKe8sxLGlu3JHquaX8x91bw2Mpkk7uaRRA+gSB59HbfI1Lwa80F558q/EXHO
Bhv2+TpiF4Jd4eO+IAGaRe5B/RGsXWewKvp3L4XUXxug5mK2ieLAichiXWzaKels
AkxbaqrjEp3QW11qu/VpLTTD2Wf/h775l+gScUhdlqk=
`protect END_PROTECTED
