`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNwR5kSSJvzBIvFJ3WCUcgLzVjcjUuTnlVFqKsC7kqwt8
J5qYO7Mf+aD6aOTGHWkbsHERFPBPS6/Z+4Fca+JBlM4I45g5B6CYei74spVkFBd9
4G4zjVjaPR47emtvxJFkBLQKkdEgtm1mO4B2c1yyd2Hvb7iNNHDHsCJmoRrfYuFb
z+RVhwU6H9WAzuWVUTOcxuEb5MdzLM9ZrMT1YB7hwf4XYH4JvTapNhY17Oq99jY9
BbyyWTVbvOz06Ixxd1uUk8YukKdfHXEIlMoHMMPic1fG2E/Kb3/NLDQed1WDcFIS
X0dFJocxQODm3CPM+P02ZgvYCOQLAm9t07IlRONzUw8PKAacJib1KEw1XDxYAAEq
q9SGMnsrSnmyfAev1YrbY+lHEnlVUuhmuiwW5QSmugwnhEByFCNvtUBFqLr74clt
YwOzZoat8g1HCdeBxR8vuqEF0M8AN0hKmHqw8AYhyJ9mBcIRaiqnlgywhuV3VNiG
RRJzJvEU7Nb7BFzj6EfZpc/1favuFj0MIj5nc9dCLvQxbIL9gOiCj+qK3yyCCFe1
AYSoT3eOCLG/FrTyYvCm6xC4k1pgH/G7ELIeIHiANyh+PUonK52+C2Jg+/SnGMUE
czhPwz0lc+AlXUndugJRuHXFxSEYBl5gFXuae2M1+jRssvGOaJAyVl0gtWqar+fV
5k/ITCD42UeqO+f12uWwMu4MkHt9BkFcus+t0i5t3ve8TB2Q1+5mpn1p3xtIrZUN
85H2sxr2qQ5zhjdDSpz5RCpXefQvCZIxTFGZiYd6aD787T0L4WSCiRmtd1MgUvSH
uYGA/5tPIxzFcP8TTvBSybrGLZF3EUmMYROrE5r1gX3nSi1HVkGm6scQdQ6TbMYE
7WqB+E3VlTXYuSpOMH7cpB1pUhnWs0lf31S3oKDmZTy/O1iDvs0F3ZE+YGUYc3b1
UT7V0f9z/c0CpJcI18vrSB+zqvWPSJjhlHty7+bQhhwz/xKM1MTZ0dxYsBZqdntU
QFZ8GBYSujuxlBqYxl+1tugG/hzazU+qXL+g9lm6lpYnl4m59MBKu9qRRRFRRli8
RHRBk3/ZIRNAsiT1Xk779bsVu9rqwbKBC4fywxFt+wz8qNCbPXKDljh1tFXPkRsV
g9427P8ToDeLUqwpO009sI5WQSe9Bw/L/u94/GSDqyVqaxX4dN85YJbFYfEmIh4G
o/1LtVbd1GtfbXSfaW1lfX1S1nDSPJksnsnJxsFxTR7Y/197uX7sqMRZCiVgca0x
AXj6BtUbIpzzrCeobBvaPG/TVAQu6eUTq0li8e2V59IxNbXEBVbTL/Tfx58xsxKE
5CYw5daivmyXorMY4NtVlQGENZGjnCc387XbfJX1vA/0UGlFuHNJTsGwQgfVnJom
PPEb1pupdeT3fjnAt9CqWwTVQhDU4vsRQYUGjg3wxYsHYKKtfrbH+CLNOZxOiGM1
ej4avJDdbSLeOdWe72uuZkwoUGdqwLO9cuVhZ0bDbDbtOIISNoG1c0jptO47ZNsb
kBDf9aPx6pgxLz7rZxxeYBbylQcPR0GdpKouOVlvm/IA4xYWsCuXUFKieJekPhhO
EeWL9WCfrnwkeQptu+y6FhC0H4GASoyMrMwoAh0u3CodLzLmMB0Dd7r0gHRbf+Rg
cwEWHrADZPCWSv9b1N+o3x5rLA7YNQtIeR8QR5F22H3+uguq8PqG/2ygCmaibeSs
0dA7TKu/i4AvecFERwk5ucsth8YZlMiWKyJx+Iw749UHFMlnNCk4nzBnO+cDuNOZ
H+9NsHLwbSaR70sKAOxnXfcpNAO8CYYjuCQa8Wth/S6RGEINcadX2IcYc3yAwM4m
kET0OixeAatHctjS7bkx91uM2UlG0zAf1QS1T8x+YdmtO9nXjTHxENXUwzQFwdML
QAbsTC/KkvBxvsW+oGB37bpekoTdnH7PqtnuQ7u8mTHkGhryPo6QFkmQ1pjj/tYY
smA7L1I7ofI+PKnFSzwP4OP6Nsk+lR6FLQTjVaP5neOiHzl2270YGvL7KZhbOOJA
t2l/QLlRbpNoqOjL2hK0CalYV+gY7Vi+tzd6Y8FbaF7HKmGj7ZhvcwFgbIJ9iVeg
B1WEDEyS6ikrkji3z9qS6eDoaK3JiqkZHvWmC1b8FhE=
`protect END_PROTECTED
