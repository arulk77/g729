`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
zkr4X83T5QFlDr8eI/AdIAiP1vvY6fqaeAQVPCRFjBWsrJ2XWiFfrOLY86FfEX7x
hyhk38osG5A0jdy0C36pIFOYNj0P4lNOU1BWotnCBbah7flkbIdTGszLCzy571JA
+S7jzvOEtXqIaZ+ienJX9gJjMjHMbTwiJm9f/PW1IjHGVt8v9bRXl/C69ano9tfv
RJNkDiw0n8YB1d0MON88EX/usyqxLPl27fTbSR+Ya4ygmVHCSQB9RQlv9/xzfnFF
lQc/0n1k6DhS+14Ya7mTYC7dCOXax7Ug0X1FogTssPJucRI0kcfSOFiqj2X55l4i
vZ1VRoo3GR1j+x/VTuqt54Kgjy56oTwLE4pl4vcs22+B/1hZQH7sGAhWONLhTmrm
XmlyXejJMbvtSkDJR+wT2IflyynCL8Cy1Dm2PGFT+h/7PKpjfR4T1IZGGg1f4hL/
t/CaPVcIheqhnn4U+ytdBUPmdjrJqsQYmmY8O5gJ3Yb+MMLHJY1d9KTHIFVpkSbN
YjGWmiEo+TgCXOdt91Z0Iwd5HHgSEphPORfUkBJ1uMDo5RHtoRtUT6+KwGQSeixq
UVcgqAbn4KPnpZendtZGemyQj6c0GO9CIfs2FTBFSGcnBCkYpmK7dgYZGQ6tGQjx
jZEOcOIOF+g0lgfGXukqZpLMDhrt3DY4W5IEsFT5BZoxPW27BLCYaqzbY6dmU2W6
LhS4tyi30h/reGqXWZTrDA4yeNnQdtDiFRmpU9e3Mo0bNk29mYT6o48Y7R/4c2QY
6ajaG4Ex9KU61P2OWaJRMjTmTUjifZPUfpHnZeKFaCvV8t6eNLATWfn1pt4hgvRA
q4DSZN5KcZEg+D7xWZqpumd6uwu88s24iyURYhUGj4Hlp6xlk8/xu7J7Lx4S8d8T
izYZTZaWePn7MR9D2Y22WabmEUlMekfDJJqtgSN+MGNDSAhZWZri3E8CgNuuSN5K
ShGMqa+AON+ojIsiP9ouSTYbPIhrNhPMhkfPp5dD3Eme3F9ltJLpSTdF0soiO88i
1iF4L2a5W/XbwV6e1amelp7GYVxJFYj5mlTFzbNSUWixVUchwpJEIBGWvm+V/35P
XTBMlBqOKESFLUguHwWs502Ixcl0CMn+63PYiIsGKaMZbgg1+sQggwx4xjctKbZq
x8c7/QjTMOHHIatD/WxAN6mryLM8Sg0CVXVvKCTT1R7WXb3R81CMcRpIhAgO2EUG
sFG85lzQ8V+Vy4PUts1Hlexl52rSDl2nxnQ0kANeaJYH3F8RSXxAdSq+6AsaAWGE
GRdxPuOMjeuJhSREAnBFEGoWqrjxEhG0HdjYHyT8eixxEKvCCTNFj80HOuz0vqSU
6xSqkxJ8EWutifbA1+wxSaLAAopvJ6KA1O5uZPyDUmk9yVTbbEqUuBKp7ewPzuR6
VRVdKwZNUDA2dhBOJlXirE4Kj4rKcYT51Aqhuug7z6q/bvmb66PfJ8kWvmG/2I2v
uJLy65Nb3Vvn8wnyGZEEfgKcws6oThsYkuvvzZ7HsK+2/5kMn8t9+g1A9KNuArQ0
0ADN5+A6zsuRU7DPXNns0ZAXQC7L9tkv+61kAFjMdaPA26+jFDF5oN4R5S884xuI
x6mN2wIOjNdMy8wgjPq9EVsOal9vr5aIqYXEB47x+mkRF1ykxq9VCynEr+kcqPG+
ygAbluGHfdPWhPBUBJO5JfYA/rmaYnJt4ArNgpjSx/dpOStpRIS0fgujEK7eSC/g
15wvdcxmS72TCze1OvmP5k20cp1Pq9DU2aGj78cCQYjBOo/2pQFIfWBEROeN/RSQ
gHxNkFQ7lX7dzQ0c7Y/YJoNWJdcxw93ptQt4GGjRJoooYI9JQ4dKfwT+X4p67mGQ
Hn9Y4AETBbw2X0dAV6z3VZ02QnoZr6adhATwarE3AmkZJBEBwctVt0i08apSJ0j4
+KrYjdcKwu+Wdgaw7NRtoy/2ONxtrtFdpW7xMHx5q+cuU0K4/5iPm2BGqnJtPCrp
Y/JjgDNkbwpIvY4gkojWAg8CF6fDNDllqbcKvUNTKdUcVaUf4UnweTueVMTYy3tH
i7F2NlgmKFz5zf0ZdxO0x6GKky8Pztc0qIF5SHhsFXAT01eUAYGNeHYh7kiwfPBv
Up+y2qIc3/2Gfxi5m8QJkL4V+vKvmAzjLed2auJ4nYuDSwkIZAT5NivPeuJ9Ohbg
6c6f+mQxGrTbSPIzW04gFmB9sh5HMbgUudr9JNi7cpSIn3B/8xMx1qNfnahfIl3S
XF1pZykAd2Nu5embJrz+INxohHqNkdVAJAXD2z8pMnKyxZTxrSnt/x1VBE5K/bYr
7+DoEGR0S6sW1m0uwle02FZnAhz8qFGNv6OPNIR9xPhbc1Ngan/FMY73waNfqZMR
SSoihKwCAmnehAq0d8akg3rTbLve7EmjySSNVxh3vfjfdQl+22fonkHrWIUHWHPN
cMvPePWz+ZWR+ZLdLx8yhTB756L3a4kS7NYVZGq8BmvtvobAOFutaKbriMr9HwFu
W6QFX58AhAmLGX4Wy15rT+C809+ekY8c+wqazDNl6z5X0iGfKUqBFZOHQjJj5MLE
pyGPR/mHv8LZiB4THVRdYb+ZnWjAzM2SSbmhug0FoQ1ackYp54w1Aj2ayOdgEiBT
Ul/lW9rQrQKtgmO0qQZk8j3njo6UdCLn11T+4PZCXYuczgzrU9o0l0yBI+rPZQE+
cH3kvOUdx2oY30y9W8DdT3ePSwyS1o+xdfoJCbz46QarnAg8jnPYzA0j0424wlC0
j51Sc7bRXAnXPFNsDU8cYHPjcxaTUwg6SShil6WFHgLj0ZOMlc9eAaXRm7+YJ2l2
s13hVJnUwVfk9LhRyRv0ejogJUsnnETKp32YBwPR8XtdBQpARavD8WeuWK9fCqCA
mr0g0N+kzZf27BecJvPztTmyjylyQjHS88IQf7TqCvm4K5wdJPMDIpPq4xpizl71
cgS/g5ZadM1GuJ1j07iAQ3AHbqdfG7XxbRHdf5zSIuZg2HcfhNZx5apCeuP5Pzc4
gTHdfJC/IVex+NAGDe9728cEmvIyLIPbfImOC+YKlayj+k8R/2ZUHBWPiss9Tc++
14gjRI1Muulx5U+Z8pJdde4UFIzM3JkFQJJnXAq7byJogXQU7sDdCJlwQdDRZKZY
5gPYWwtc41DpGZxvPQAhP82nSVmrgOLVFbBub9tuqnMJwg3sGk8pRDlqX20oblvy
vZd0dE2L1fLSrOIOZjNlv3wvZyww0K8PfHlRgPKTY09yKSCq61xfsmwbZshZ8DrW
O55IKWt5+XTyxjX74hv93EwlIJlsb2X79/QuZEXjuZqXY6u8vtebavyvOMaLeS3I
j3XRZfKr/djcTgJW8UmHkZE6vZzP3tN6l+2Ay3VD7lhENR+O3ZqGdyFMaqgMT7cA
PWVQCUb4ieqC1QwObY9QCQ7vo4tKbH2hJPjyBlytg2oGyXgB6fNcBOfz2istEFwY
/FuXsGFp367kXrrEgpi+QSlFZCiqU9dgZKE/vaaQi74Fl/pGcVs94sGl8aLc5ajM
NaU3NOjbGVXQIbbCgNV8jXxaHQWx4WQyDH6/RNV1l+H1tHu0Yz70Iu2UXa1A59y+
WdwGw3skkgOErJ0rkpk3RGqYzHtiZ+uRhh1hmTIwQ+g/Pm9HpKYA3ogx4jGmIqzt
OXG5YQJ6X5kudGoZmYWphTCcbRJuP6sZA0t7ZjfvhNzuqJUum62CBVfS/3GhB38F
E4opSuPdlBUvDOPpP1InoYrNeassTqD8L7zT8jFMAMrEvRtyTWlILtf1qcJYisB0
xlm7Hm9FbT4heptHdcJZsmWEFnpwzelOVoF+jfI43awu3sJifz5YG6qEMAYAUCYg
xX3YN80mtNEfcm4aV9nU6R5GyYXEHArkkAdNYfHQ18v6eMp7WUKffXTPmjDo8uUY
qlCrZajitjK8a+TVqAtHQZHyCG5EgD5WRbAQgTjoom/8bXeHGtHf8SO+pbzmRsJI
ENCXC+GNIjpCI+SYrX0AjZttKiVDpep9EVOZ+w5w82Cl/FTJb2RUvWBTQmGgUTDC
I5JtBJ0thjalIdgIItJ6ry0asjdfZMbg6Wfzon5E8YQplHcuTyRg6/Tfk8xYdViG
yDGoo4cqsthcVnPGBbGcFv74c04TfSJ59Ed0faqfnpc6ikBSoAcObAAEDAVfz9uo
v+LdFiNN1aEKDwoUYZJLh2jNwniWQbdIUcsy0C1418rAl0X8E1MJxX6SGkrCDUz7
w/y8ilDmpEzfHFhP34G5p+k3x4lVOf+PBAYtaw0yzNq2nrBH1WEWSeisDTLythJg
14xJHZmzu4pTODF9joERa0zvAL4zSo6wtJ5rCMPVwUkRDckroR6SNJGOlX888dEk
3bzOHXX/JptOAYvPlq6OQgxz3d1stEJ4A3HkgHNthyv3g0XfTEqpAQlKg73iZxTB
kVz/MQe8C+ZihAfxWqFMe4Cu4kb9TdTS7d8640kux5suBdXOaYEk1ag+LcxUuepH
o+c1TTzsJ1SL4GaLteTYNSmV5ptwlM+DyQOUedc6Ne0imoHMBj5egVVXHgHnuFOK
dYxHS40go9HKY72smQwN0+HpWl+Jh9xbtZXAs3fV/2Idzqj6XyHOJqw3fV0M7qqr
goi0SAqUiV8iwznR2LczesJnrr7tYfxbTg49Yh/qssPG/UL1SqHVfPZ6d0a8+FDR
GKeOrnJuGJdGW7Sp0hqtvJ7OWXktf+AWWW/Y2z7xaYLEGVk3/41doOWA6CEEH+Td
QVOrqFTJN1sUy/fY8jXgDCPVc9hyQeAjLP99h8eA1BO+bRenCI/ELGfSlgUF94rC
fuKFrc3tQUu2drGptKJ0HRbobKk6viWuMa5pgYqON41LCdYtSEu6s95XU7aywgwn
NsxRKPoeyZX+CG1MIxTHPbJhjB8P4sVPvQJ9YpG7F1CkEwpEqj7g2cKYON7+DIRl
0FeAEDBjmyS4GXpGPMyxKMRXq/GA4Mf8egB5/dFZWgRrd/cngeM74Bl9l8KwXW9y
TBtBQOFau4Cpiwb/dRqVB5S74SSB3Bi0SgvjeRVYXD//coQj4YROFGLTSdZwOVuA
ljAYzh+8WXwaD+SFfJdNmEygaVZ43Y8q5DgYEl9y7eY89nqYfu/YlUWSjfmXhWjG
pnvufHTV8/axAVFQftJ1240ZQOgXgoVzonKKolYh4XBZ+20SVPeTeK/rxw7jxYCE
r4rKwVGhysuOTKogHBY8RRkxege8+3Fv5+RsxTAVWmJsRj815AgVJFtLHFdFET91
Je25Wyyu3JSOxIadZKXeYtxDtdAkysoatklXGDBS81HQN7+rcuUkQv21BzyYeokT
kn+0uhr9aFjIRiZqf4zqUUJ+mQF0iP76YZgTvfpnpZs7knkdxpZVdbqYdfAGeCEv
8oCPlzTYJ38QHrrf4aXWUcBU2DOmuwXHzURVW8JRUiMgDBqthnU17DZF5fSiAEVh
ToCqjC3ao1SMoQGCQrVfaq6viCLyOXMhQzQZuHIRa3gzpesFpvNttNVkvz76RSZn
v8QspWi90FUVUk8Z6XZFrMKOvKd1gHqo8qkqF4zE7ja/VFE4c+oPBGoeU+Huggv/
L14HmRejxbAYr1c1pP/iOswwlfbmg7IKjsU69PTDY9GoyLGUSIERLOO5xUDWJZ6B
zIGsHdVr5hmegTc3IWRzcskRoSXbsG7m/U0TigAk+arGw87RhcV/qhh7kncdzn5l
iWkfiqMsHkaG+eIWyob6lLB98hTXo9aCzwgPZNqbFvDYW4UQC7wHhxA/vlggEj2P
4fRKTiyvy3VbaqFf+kJ7P7zaWYNPxnpkRXNmCMeMa+g+U64OAXq5lD8ZmN7kXxma
1DX53xr20INQ57bJZGpGqZunUvbVqNpVO5tUj8p3l2VZtYViF0QkLnCmGQMqMzly
B5+KqzIxnlo0Z8LQrmhlHo6bS5Gua96I2he8xcbbWkpllwvfr2LXLfQ1PSZehctc
Kh+L/IW+EjOCrlxnzzZQfXgjYX5ipoFrMvy+StGUWijO57ycbrKKUGIV5xJCmEOH
EAk9BGQiYWy2bIjtbf4vfBMKFCbFQ0FVwdrPFZnvdCxGrPImhY+UjHHMUp7kmAbD
HJzo0JfrKWuAIj1xDLIWptSbje9ZF4TbKA7fIQobZbIy9xm3jAN9T8CToiK3WLmZ
b5mT4sdiwMLgzpRTtdFygbpXHzmEGm74SLB06JvEsingq133AempXwDy5DucQRu4
EWRHf8hGc1z9/131F3f0Tg3ex8fLWX8iu4N5MhP+b/ntX8i45cEhfyV8QnBZENwF
YOvpAgdXmDor/ar0Uz4BN9FYgqV6JBp29q/bVzVQ/qUlv24EVOnbZy6fqBPPECf/
cTFtpkGtkP/m9BHxSlpAhaQBmoTyW+ipYBubGiqnmy6OnLf6f3QzLJCIN35Bcmpp
VAD2/Wa4+m7KOGLmQcoZM+SqJfR96ZsfdfNE5/sLJoJ9yk3b+vYu1UHRwyKgZInr
4xK5v1ihyRYrecJpzuanRkMCmvI1dTNfHv5P3XIT+WQXujrAEH2N4aIkKMlCoMoD
V1H/Zzo0C2sRpk7wfKpXVIRr94qH3kOsCd75QSK9KaZKe3PJPk1G/hng4kAarxgb
HWfBs84AgD2jMgFHlvJaLw+3H5vqNmNzuedogYJqldh4XGtXES8QUfUQKT3xWE4e
EpshyWyV02q8Gli1xtqK3eA6cufpjzNHikKjc04hH/ZLCHpIX7pDdpVuHMDQq3ir
stEYRUzA+Qs8dS/s69P76HTsZVaWXZTChrVE94R+Pv9PFwNnvfL+j+RKMBHBY/0M
7eMRK38Y9M+ZHq71xxwP03sHM26esEZELCQ/Uyd+OUzMVzjuiZHd6Xl/FCw6hs8N
o3h8ynSndy06r6Is1raZEK2e+VjKmvddGSwfO3+z2jlDavNcsjj43HbTlIBBtn9y
sRFbzDHMf5mWACOT9/ixmLpGFIJ1hvCQI1NIRzSziXk7YvWAY5WtspZWB8zjnUDN
Ryj4fxmBJM72tNcsGUAwKOiWDdo/l7xg14iEUR2jyypuCHuWL/8Nge0yPkIwIrCv
cJUnIEVYIAwyFdPlbTM26fOnc/U9qaLkfj3AmGIAzp6ulIbJJ91OVTM3Ku+GV335
rX3BC4Vd4etf3tJKtIJvxU8mkkoJ/p/2vMwEV88B2YbCeqGLbUMsqyZOjGjQaEN4
cYbMAWPbLMiV9SIhsyctv5iv34GvHzCkXgk4zxPQPACnbweueLh/wwy2m/j0FaP2
sJxKD5nK7llJ4N5bQa4DpRYse1I7cFO/e9C88rvYEhWjR+emnovYiTkomP+RytdL
X7ySFVaX6B8nFrhgaoAwNuL7GwP7OcukLNxO0D1rj9C4UC1Ers2qQ2/G0m0Y33V3
7PqgXc1s9aR8KXrTRlA7GpMhl9SfkttCgYxjb8L2XGkhRI+0jiGAFJic6IEu11Kl
UMz+/ZWqvSS8wJN6UpL7E9D7ryIsetLKxVLLBg3uOJKMRxMqDtGV8WO9SNp2gKtL
sNSETv09elqy5QjnJ/iGkogaMwIpVBW9GcvfydORZzVQ1nqSfy9/6sQB0Oh+tC72
YSyBYU0UttUBu7y8HnPZNU9pL/5IAQas+s6DmZ4aYRARfzGykp3XYhiqv+2QY3dR
xmAQ2B0XzeZJoB4CK7lklHjupRX6D6uQYRESgGS0m2w4syU30wCP2tNK0YlKLwis
tDuPsRdu8SKQfbj5P8s4J+p9/oSrfNeR/i5bxSbDsyZ6JoyEHyv4HYQzYu81uDKf
k88LDZXL6McpTTFnuR9O6+3wPQew2euNhmI5u2mFLMJBN4A8HPopnrzXVG3dBfBs
JZamh7juiqteHxJyDOk1hzTBCNhaQMAlw8dREpyIeZJATO81llHj9eglvjFVjmse
ZcTPfK57JYLzB9WjZaBQZdJAxVYO59tn6rHxYZPm7h5efKXlqWhqhGO0bzY70yrn
B8TwThaNhMcMm5oAEYwIHEVEOfpTkfQeXU28aZUwDZGOxcHI+MTdLrtOShflLxXU
IiTDJJveSy5F4xA+pX7AmRCdsC4Tiy2bzgWoqIeobGbIN7pWKYDoC5ArcaSb4jf+
u3ZCB93oywRgPtf2fVsjbRoKWOMSiCi3j+oDiENx2va4p7dTuBrlekkB3HONB32t
S1Ole1/UnwKHBCqIDdWrs9PGGnxXXnJWlAUAgFZ1eMoHlZ/JRYUU4YiYIPu4h4wS
I7KbPRVmzFz86p7ax5ldRxkeG3A1h+dsIqA5F3s15n0vwW9dNaVWvUWBva+TpbCF
CIqHIpYFt4i6V5oUcx1NzyMUaB5/PwijbqSBYDouW3Q5p7Y1UlOTAY11yVatSnOe
XtvE7JV/TJx2q4blXeLe8KIsiJL612BFqo3B7f+RLW1pJw4P79dC0fu69PkbLW7T
Mkd6k3xse5P3NIF3w+8u4GLQMJCPat4N9IQ3q69mMENqKdo0zWk965ILqnaaWv8k
7/14rsAGgQG+cVcfqUlEtQ09f3+UTJP+5cVDc8ddoYwjYcwT4IVEH8LomVJS+Su/
fF1ozQYrZxivEY7Vp3JZCDd0V5wFmbfR24l8Gv0wBSANMi5fRMJA4kaILg83MUP5
9/hctz/8YPy7OtlDCrJ6RxAimxhgg6QrcctIz0ZQyBpuHuL1NyThsL9QFRkvhJ3z
bW//E0hwiO7KU9nkdso8DrKlIx7b75yOwi6bhOmUcqhQ17ToJwFB8VL6CuTUDlc1
lxSoKAjqkYaY/0er3yaA4YicYzOuN1zEO4dR0MQCw2IDjj1To2ClUgbF88FzDNLR
z/1TQNOOspvkhWjY5gttYjQZXLWTCNLF+xU4KUDBWstoVANXYalrc2PCRKQWHThX
nFq5/8cNVXFcOsgQEofGxo+31wD0NQYFW70/EV0mTbzm1VsPyDrnl4Nlm6leHbOp
9JLkhrP+Wbt9zkjZ40eV8eQNTLqVgwUzzK4Tm6vT7micE5CjIYKGg8yNOPDwfhQN
eJaNVtow8P3tS89A1rYhwXK0tskKhE5lPBf6DVO6fvX3kNAJ0ocJQJgGXgAXiz/2
fXqkeKCfG5yp1xN3If0cUw==
`protect END_PROTECTED
