`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
36A/U5tO69wVl401zVMLLURiZ6USZNUcQtYoN84wLin3sv/rEqt7pQXWnj8/34US
Fb90nZ/Q1Jy6G7ZfB6lg7F4m1RyA9hqXDtpsBBQFia+0VzY6ul43bCmZo71LPgV7
c65SH8Rd86bTE6WQ/C/SUFAgX3DrS+GwSqkLpwMQdklRl3TDOFagSsqoPx30P/TB
94PYjbB6Oz658HPbxkZym0VupoiCTOKSB58uvajNVMUGj5gRmzrK+sliutqzChyZ
`protect END_PROTECTED
