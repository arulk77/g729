`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBcRx1sHYAouH57/iKFO02CoXiad/ICaQcAgHzR5Uw+L
BUpVq9X/6mYn8lKIxGRM87VikcS+LrBJe9ap4qyerapmCRS8eQLji9uy/hGCGefg
vpIt62wbnF1E2ZungxpNPQmKFqnGRvruAZTCGPMObPlDfpqbyRRPXc8oifisxsna
I37yBbAQrZJVLTjdHnI9/5b66GgCb42H18VCc+kgPa8BYZTlYErP2KwZAslgSaxp
lgx5Ry4Iev466hgHlMTsdrtORtqR1w0uQCStulQg3oEUrBW3f0H9pU5MSJYdJCVv
4UN2Xaud8aL1UF+HEzlqhOIPbyB81aoJR+vyIvQPFqo/f2gXXvp+QfqOiIm8b4ae
WdMo4/rhoDIKRpmRErqgRA==
`protect END_PROTECTED
