`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43br0BL1iO4w4IkIT3WEf4QKd7apdC+Xb4qKGV2Un1Fn
laY3O2uEM/cVCS8aNw6qOaJVd1n1uDwxz9SpO8NB447vJUn3QSJkuJ0+3jfCN3v+
tL2+r0IjyI3Wz7XtQk6833CcYishjaCeE70+aWN35rcBza0UCkZXFuHZaqYyKRZj
7NAykF7h+QfTxfwVmzF8RPf6igs6PCG2c3jnXmOTTjGcZzd7huQY4PszwhSDXEZA
Gn5WSw5GoWJMlpfeSlIdvEG86u8+FeHU5eiBHSCCL63gta23DoYXc3LzhRzd7qfi
/Z22ap47IocBIuvWiHwQVhf7ww+984geR85l5BqCWXNJ423zVmbkFwNFqmSO1lie
ptgbPqB15F5mTPMFumz7yw==
`protect END_PROTECTED
