`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG7msVRH/PXfD+MGA7zjPl4wfFFBHJLxWWFITuo/lXsY
EeDdgfu6mQmaZ1Z/o50Nbsbg0VuUTwe988hrIJNoRBeOj9C9FUHGYzYb953Y0zyF
A7gFGqSAtlW4yWYMvIv6UvhYih0Q/MZ8HFAjObae6+jaJV7JHx5M163xgYzwcqqm
VA+o/N81gu32Q9N0qkzRVwZ99FlYXbdSPJbso9fDris4MuquA8Zdqt6IzPwMBLMR
`protect END_PROTECTED
