`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aYVAdwc213Uo5YYEBCsIdHGZLyPOjAjxqqLhH8ybpnan
kQqeMQvq6Gv+j1bnXXYF7I2HVwU5ffqdiue50gE2Hf64vM3X2fDhWw5S3q2SCz4T
CXaWk6wXlyqapla40clLPRyuZ8nOZaqBnbeE0jq94pYlXEbWB0n36lXAK7eRcxIS
FXf13VULPHvf5oBOq6yZvLn+/MpkKwE0KRbSH9afr1Djx/27AnRb0vaTL3uAhl9d
mY8kZe8wGUfWMVHRrYhjQ2CYp/3rqHmZ4jgbVmysHaSb2iAbJk/tFtXKdRzy20Tt
vqCXGaTVsAPRm8eAARL6trpLsDjoMe9ezBEGugKAXxs=
`protect END_PROTECTED
