`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGCrZ+MHhG8Q0AKdAW7w+M8MqskwVUVEmLhNLQl6Q8rz
yrz6/ZZh44ntfZFHxEsh4YEbQm3LVbKEUKFBLAkH3r22QXPJYbjV9AvubF5XVep6
DwIZ+8/n4hJQtLQDqr0LePV2hJJLVOfUllIg/BmGG09gJlfPMvW6nwfBv/LXjbUp
`protect END_PROTECTED
