`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
lfFi2O6GByRC0As0HBySRj+UJPhzs4rHIki9zSraQrWEZBuZBMcOs2InLogR7Cuc
x1r2cVrqJ5Q2KJAE3CsL4krNR01k1qdv3KfwVI+tgBKCv4jzNADuY9WOjgGh1och
IQ1e6P8LJUoihGxseZqWtdUyZjk4aiZX+wOyGBS8RqZIqHhBjNB7MyShd1h17yAX
FfKpZ4hWRa4MK4bqbq7uu81grDaT6WyJaKsAcWQiqADF2R10Ac+Y+Dmy1HH8QmxA
zxGURk+XFYgUpjQaek5YuYHj+MKr6lHSMNVj79JOacx7T06be/C7jpmkj63Yp54V
`protect END_PROTECTED
