`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
YxJXscI6clPpnhkvA4Ptt4IDSXp13yvScs8so5Y//BPrUa2vvZeUe0d4niQXngxw
EHZgiAm2JtSpNxW0YM26J7sXFaEgKFmq1UK05QwFsPRB91r4Du97LnGKvjyOljjm
kyGU5LCIZqv6TQjkgAxUFov7ww8FMj5pHGSbU4IN7zWVCtdiDPSyIL8YgOsmmop2
aZ2RjyJ2JetJP18uMO2slkeB26t3HJ8KMd1iJ2FZBZ4=
`protect END_PROTECTED
