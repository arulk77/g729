`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEqqREtS4XcrdNWW0uodHw2GfC5fhpWri6UfH8zfYy4B
KTou2EvblyW/LlwLtuFZp8b2WfTy8BKwKN54nB1g7WO2nWAyRRZUKT1vn7Gxcj9J
El8mrcpX2kryAS/inxvTlG2+a6zc/x/Ag05J7juYuA6eh7poo+Iaesvjt/TdnHz8
rSRqTGNKLSIkm+VtehEvDFfgQDQdE7EOZWGpOhcaqFPWJIROO5F4LZalkNxdC9UU
dEG4Mnddf12DeJUEzVr8CrhIzpp7L4vXs32rnNYaTbjo3TH/Hs6SwKyFGHBGgKrb
NjekIi89x80gGCgjjwyJHX74vOnxsG07GnLSyJcQYa/c06y8Db5qXsV6qpTBIcQO
BtGE0ezLNW4aL9vnD4qrAr4Ba0SAJJwRZZtZfKCkFISmJYSAjU7kUWL3iW/htevN
HTfmPBO0HIjndSmRd9xKRpNaQOzHt384qoNBBcnwTT+SMuFuXzkD905/94PVw+D9
J6CQDMoqiyONg0fKG11eMuXAt9rkHGGthYDYtufUlp5ad6/KKSP2zBTosYXJUHvc
tZTXc6DielSbOOyDq/rOlmLGxrVAGCj4qdOfsKPzubAqXVGZUoQYokIfaZdN17Pw
vV0loZf58YWrP7RLzAumqSGaRO3+pxJnzgso29pxYTBFK/NTvuhJnYL1BmZQQHHc
`protect END_PROTECTED
