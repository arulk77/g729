`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK/v08HCWUxy1aTrL1KHMvyP7BXCe5IT6m9mKhINBqbL
RUtO3i+vYNhtGCLFdpnigH9O4HMyw5q4Ft7YtkEGOkCfXvraBvqyxStwwNYFc166
ZZh0j1FIjQubFvI/dmlMkxwoYjF9fef+rBKf5CdOhBV0+fE9CuwpfSVMa3uYLUId
IX3yZpBudOb0TkivzZetVodBlr9bMIPjN9WGfM9E9N8qdcbZNa9fCELAleI0DTJy
`protect END_PROTECTED
