`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIBSIxjVJhZOvvmpsoqvIuoV3XFvdaOmqwZ3RnAMLqrq
CmNIQpq9bOGJzxWmu0VSwPfbowGY6VNVekd4xQU+vS0FFhwMWqHXoLqyfCg4y2mf
qscsxObyBRRkiktZDZB9L0Y0MnzqTIgItdRmA1NdDbaQJn5McHoRtyVKdpcgs9kb
TtHZAAduTUKfs0EGOI9EnszZOlWSr11BQtOgs2OOGS3Xwl2+w+ZTUI0aLWLLk4wb
923fwwfeg2DYF1AXc58LOzAukgPeo3C1GyD0nkr/6atmfyHFyB72MYPKpFRnBx1J
usvHfPTNmILhIF5gabu3NtvEXymfprJHApMr3Cqfb/msOzeoujqzan+2WWlL4qXF
lB3IDPDBEnCftU0lrzwAPNfzoQZ8gZL2pWd+ZQoqNfleEk/RL+52qxRAcShLM68r
Msp1rnhYG69R//NoHaMXhugnTNdJzMDJKHTWYJsjyIsHTvXVpjN7unI6kio/ln86
v7fYETv21hWzNiv2TICVVzdhuxDmlKAbAXkbxZ4BtgutPNaSzuSdoMGSF0W1jOiU
rVslmucKCpRStcj+42DCFhIf4iMO+B+ITDM5EC+HZCJEN5IoWSoV86grzHcf2izk
`protect END_PROTECTED
