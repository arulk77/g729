`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOhUNLrM4fMs2XuXzAvsmzVdFbp8PkXhY1SEEPRUVuIQ
wfcVIffYQA9kTcLCb+VAI5XLNKTbYHLg9F9z+Vu3yEtsix+hULpIcMLACiZf5HAN
XVUL7W5IBYLet3iGido2BwXMdhguHYcJRe1nn7BWv22A7rU9MIdh6qO4KmnFrZSL
lVdcwqKbz2KgGegt5ttYXmMsXa8nxEt4hdToLG9dBeFkrJiFOYVTdzpbHtPAken0
eG/Tg7XB8973YcjV4mGETqvZsgWhZl0BTsuGFO5DlO5rKV6cYs2RjdrjzQEc5vxX
QGYbZGjpNTE7sU6hO2tdbc2xo1yNOX5J51FaGORBbGyyuqoWX70SaKPq5vp2dY6y
bZActZjNHmhMjC+hjR7UIcQFgxg3fESkUjcWLYV/EWw2yFsVwDIemmCSeAc+238+
bPjzv5kNcfsiZPFb1WHNv8RNs1lJ0pONE5YjjMiufe/thYveaZMXD+CeR3r8LUAL
/i/dVXLo9j1k0gj+KdgPoG9stDxqMqkq3mXKBMxOx432/Vfs3TZ9qJGgOHoG3YzM
`protect END_PROTECTED
