`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
tMI4c9zJ/hxE/lxA8CcP3hHlyFI5j2pw2miRZjy1+JrGcI74+QcKjraBgatGN+A2
nlktCEy0016Ay8bxfevUjMcg+IBtX6KRFVsxiiPlvSVJV3SDSbHEWQSCOErO564a
z39L1njH/OX+MGowtoGwjRLQamP260fJsL7mndKf0+41T9md/bM3ookI870TZJ0i
`protect END_PROTECTED
