`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
V87GIKFlNyr5WzNUfeqnLxq5WIMKqvIhjJvXM/Eo4bdiKagT5c4B5IBB8siNKdVi
s/MJ6//9aAWMfgVgov8rIy03mHLJeYUtryrz1eLVebbqqY7RvsP1/Xp9kskFLVAw
zGOOJLeZc7C77Hvy7U4ZqYaesloEFizKRzD29/hMfPPFiJiDQce0LhqWJBK0B3R7
ey0bBa7+ItReTC6gPK3Y0CyA083sgJhjUSvv3csWpEiG5yIGOmrxQxk/IPK7mk1E
tHcmoKUcXYhDsCNIMXA5iKFTbsEAJULku69ytcrqpmFZ9Ywjw/ryKoVaFRn7SCqf
xH2zXvPKDOT9nHYxEzhyOwLedrAq4tJybplpvk26nc+VZFfGIS5yENTw2YhJC7gI
3ESkbc6C98tqoyw0N+7iePUsEdPPeCuAOjp+lrFRUdb/HUkPc4Kv6i3nhWeLiXNZ
A5jxtY59SeGHKA5oITuv4hyvIZ+hreh7elDaVewzE7wiOsG7bIUVWL2PsBckWIU8
ncS9F+2BO0xxOAjb6YIjz+oKFfV1qpx5FlV6mLtrP1k5KLi5trEyH9j6hn7Kyu9T
4dCelUBkvEol9xcvSkU569f9NAM0gW0iGbj78/Cshhow9RLYr8H2A4gLKvEgUjrI
Yb40P1UiwC5N/aiB1+TXC7UjfTXWGEUe3N4T1y5HyPGFTdKeAZi7U5z8Au/KjUm2
Ydfkz/QJaFaBtKF9YM8LjQ0dEQHMhdRZeWuD+Wn//RzK7YXAu1/fKxluRSn08Rj6
ojlApQ/ukgxgwbsAhuPvwxF0+4aArxtWBfFfAQ2BZWxomp07ewY9C0iCkFMeGEh2
KcKZPOWIdaGQGIuuqcxR7oJIRoPzctXMKqFS6aEOCwS19k+7NT8IIW5+rTYcrPJ0
WOkuAugYkiMw3ierKYp78slmWu74s1yW5IxyegnOc64=
`protect END_PROTECTED
