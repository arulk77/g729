`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu490U4de8pQAEq5t91Cfg9fmE34EH/c1pD6iF8tSCFwSe
aCtK0Ic9/dXj3Rc8lSuwq3cZi9d1k370Os5URo2segk+4HObjXjyrbpoajgaQEGc
CLtgGjgxK2Kw0VLdkMnFjYTELw/brBg00APAXwk2Hnui0Sqywfc4eaEgKdSqPsrO
oZYyY0wl1zgnkKE/GSDmjdrQCJcDK3XKHKa+RsE8Hn4=
`protect END_PROTECTED
