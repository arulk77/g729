`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJmtrPd/q9HD/Jk/kTgckocgkE2aQQ/9xO1TclaKk2RE
IFY+pio5gA2GRF1k44/x7jl4BXAwE9E68QotmTftwaKsMuDE725MbpoRUWtpkA9W
f/WcwcHda3HavqhmkLHJu92gGkBTGb9x4weuidU4OlSbyTW232wIlnHo5ero29W8
xiCYLfHTJTKp7OyNaMxu6g==
`protect END_PROTECTED
