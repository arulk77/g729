`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bwhVnw0s7h7dYMvvIEPR/PbWU49QAYG1QVhTS+mK8Mzb6LLp4zlXT8t8mil9WIMl
z4znJfyPgfOc7M2S5CvJGUhz9JQdKhto8KrK95aO+eGdI25lEbUV31RqodVBguKP
OAkREJLEBRra6tKuOZsOEcP+O4iSeCGZxh+nzqDZOxCGYKt0pDbJx70c9QX/ZN8s
hCoUWdj4Qc5ZX1zjbFCFqdV+Ll4sZkJF868PvPv0ovj91iRKAErExolxN0Gm/CGH
tVHuxf2PWEARQlUhdQIzmlVmCu23o0FO6mDpD3fPmBHUl4jIUsZODvC6AiaPIrL8
r0tgRDKN2xRzTX/1ZY0JNbMOJePnlN/+RkRVVPW6tdE=
`protect END_PROTECTED
