`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu433TPLwcckiWKPUVe7Xx7mzE9GDwE8Lr7mlXZb3ALHef
ZKFZy1tTv3rOmHYUr8t+2wlO3aF05CllEotoxK3m8ZnlAqCM9aO7YlhM013Hw1+f
csk+YpWM20UAYgQxMRTyJlGMwc9+97pk9nbqOG0T9VyXTLIMPuwWxU/1p4Bn87wg
4OkJOEzN/wTzh1V9jb/6bTewcalU/5C9b2rY+bJKwU+LgFoR7ZXyT8X7kIt/yfdt
4vNSDPMYbvFnK0FeadDQqrht89g5d3fkzI+t6uCza+VMn9A4oQF8AOaCkbha8W3c
LLq7G4N5B0t5XXiCMdCRIKrtOsiGEDg9Yqgt9PgyYkAP9VUxfRXzVNIOhhasGWZ+
sHloMHv3HKf61Z4hXD4mvA==
`protect END_PROTECTED
