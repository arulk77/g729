`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
L8RHw65oaY/QicePztbfAPG3X3Lrmw+17BNXm3YuQxesL6WhJ7ZFNGzCF368Uz/p
KPbl6oIdsbSlsbKRbbO/PVgCCR18pDgNCnJwF0rSgm77M19mmAqfCvpv+f2xjIsr
`protect END_PROTECTED
