`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Prgb+lMGK4ankHVaNnLDq+grlOufyX0Ipf3Bd0ERECRMvOuaROpi9J+0505oWJsb
8GA+OlMHUz71WWQlVopQPPi/HR4JicDj93/o4QKhKM0CWWY7PYdJEJdJN4fwyDNI
OogE9GaM97qhYYU1g1s4N/QRUFwVAOr3s9SE47xNfVnNpFuQHTo/a3osuEY1A39M
silGodhQ86ZYqXdc7u6B2o1jfU+vx13nTAhHWBL/w4crX5ncgUBXmMaSBA7Pl3FF
QHakPq2zRFovjDuhYvHVhyncYI2PObfRJOdT4qzjm4DwEeIQSQSGMbQXcumcKrs1
`protect END_PROTECTED
