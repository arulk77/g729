`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN+1nzOkZ3hgDZGaEP2Nl9g1eoCkf8Xzbkk6crkGmIW/b
ggjfSzJZRTx5YPcqfEVcnoDW+VthNN/g+msLru0Md6oqalRp8LrRykk9Ax5Qj9LY
FByHdv9mbYN0oxQ7uEkwLzGC2ukXhxNr4VJWz2wsiIjyo4xejKTk/X0GJrrqT2CM
Ln4iB7udYIoH4vbTsxy9V86Raa6IEaPd4nMyL80WW4KuF6/z0prN3mzCkr0yBSVm
wLndHOpqwTy02IpzYAcl3gfCxk4A/hjOLX7aKBQVVjf3WaeCz+xgEXmjIIw+FCA1
1DHCOfQ7sU5FtqNKwgWYcWRkfjJb6b8SVMadjgvSda8U4G2THiCorciVT22kPNCK
MfQAXLU9FeHvT1D9Uel6qg9PG8qlZsT2fNsuIuSK0JvPEfhv5KeWkACSwfTrAcUd
Can6Pk0ZBIV7p9i5oUPu61gJQ5ZjVUEOHGVSObCESA2BCj0xtHhs6Lkb1O+CkcKL
2l7nCQ6UocSirGDkcSXfhIml5FRYYozuI5SDXQA7zszcyaSwFiq4pSm9zi3O1YIG
CfzxQXETmu/4TmxZF19DevOzxOFFi9TS86jR2J2TKY9YV9Cu9ZJcokWhw5ciE0T7
MdzolsdB+V8nixzxy9AutIxspHveYfPBH70Nt+GDwvfC5MEqdGo52eaWQvVJp499
pARZSnecuRw111YZJyWVlQER74+bKJNIDMBLMtutySEBKzCdwCNFVHLTAWimxNyR
q5zYqiq1XEwf/d43sVq4DBZb4P2p3hQBZIGot4IO01C5LcXfvgnbEXafwAo4ljEx
n3Fvo0XAGnKYYo1CC4uxebhb5pnnTXkjhlRImfKNmEwva6h42iHBa9RtbZltF5nH
EoGCVCVVDpKVE116uQxjTa+V82QUrNxBPwE0PCTBNQzjUE2zl6CpueU4p1XXnRdy
xs6qlUymYpI8Qdxdinm6H+8rcdR3cGnOZFp1uKpZVBocVBxterq4dfvzNSWDFnJ4
qA2QCPK83Izz6YA+H55C1JK/Hi7g8bxrhum/C0EOf8i5WOysaCGcijbtxFREsHtZ
`protect END_PROTECTED
