`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM8ttAtarLIdABHudZ1KgE9uAlWecTLrE1cGm+843ONd
S0kCfFugDW13K9zY3gmgTlri07xJt1x+P6+jzUODKt4RDqbatl/a9khz1II4k0KG
8yWs5tP8pHrl3bAys0Tfe3E0G61bWGXIMOsha9klgeYI0jSzbekw1Zv6NO8BFmrf
jblgSABH17YHpYyq0m+Xqw==
`protect END_PROTECTED
