`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
FTGV/DDFbeID2XtQrXEgEWpKQjMB4VRYpoyMKZEkRZshXerjtz4wPmf7Yqxuyey1
5PIyX3XsbOwtitqwM8UgEVVdxSrTVb58YzhdTU+6wjVnVLGviH79D4E8CgQ5hjkI
lRkiUWbjFxVXDSWEXZR+06PLVgLugyhg+LtcVb8ylBhVgpvjn5eNihKehP35yESz
VGkNNCy8Xz1LFlnn1eQ6qzwe9ad0mLoFy3Pyihj153hWBaGSocD2AoM6ZRAyuZdk
bV/yvw55IvGQl+aFcH2tAEgCOr8aE+Y9KBixRmO7gVugLtAJIappF0EyXGY9Ovvg
GuGiFXTkc8Z1WIxNeh1rjWzMYF9r/Dz8Uxe45DpvTag=
`protect END_PROTECTED
