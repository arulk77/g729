`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePqHSsJts15f14OOibp+v4AU7KIyUDL07E6Vs4HeZ24n
tJOaa/ffoBi+MbPHodgZhbPqJgL2M7b8Vb3t+zpE4fK/wXQGEG4IgoE+ZlXDGKfe
VN7uhAZr6tID1AHN8yls3TVfGsKB+JQQtgaUOkI6h0zBpFWmFGE3sFsEZzqDWkfk
IpYjoVcoQW6u1/IQHdAId4QDfZHA4CH6Mj9C6T6fibiGtC8HvgZJVF/CugFWzmsx
R4zCaiSYey7gnY9gUvpdqCmCp0//EtqczdGoBUCaho5SqkecP9m6d8haaOBMjlzM
Ia7mLHzP15ma44MVddR6GakLSUrKcVw4HiuL1/9ESyf0P+qJCOZmjW8X2zjgnTib
SR4OqY5oxPpIVzjg9jM33FYKdCS2/BrCX8/2DlGdCk5nX3hdmpJ85h1TdMnD7Buj
b6FW/dAIRvnKcPCsLsvN1s6pBVgzxcRQUK2xI9P00GYXzA8Vx36Jx9PhfMXEKFy7
zNGlvHJFfItrQf13QG604LLRGHwEHtXZrlbVzk5ZVtyMcJqsN24H66Bww2aTlR8I
`protect END_PROTECTED
