`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47tk1vmiURxeLt1oi1VqizRZiSGjMp+DxM6t9r9OZqti
W5yPCdPNROaKH9+meGn1aNV23iBIc3zqlJipkhkOXLT/aGsHqsX5V1laPmXRBl4k
6GYXSn5yxhYqw/1xlTs6Sud5lzxkmCAahqr1v9ltEs7SwdMeZkeshhpAoGqZvzT+
u8GqUKZM7e4gucjmxX0jJnyvvh1rBi3kOPO+0TKom7EF/jR9aZcz40AtHWjTOT4v
sC70ygjBwMrjyCXCB2EhgGtOvPLJ5VRwgLC1PtaIvUOO1HKjghIaOPftsV+BAAMe
hD3mosWVlNx5afCcHZjeBWRCi3EjHz0SYX0U6j5aSMJIUdZXmC43gk1qcGnjEfCb
GSEhemN4y0N7DRIOkVXXpSeLvP0BkyuQ1tzbeYJ9giPXI1oCunWt5tkrYxPxUqdl
BSZdxVqL6ZwSRGEGj1rB6GEyV7yK1zzuEvhy0D7XE1lX+XUMkyokh35HWnIZtBrJ
i1v5Mla0fxs31OY2wFU3bon5HwpBei4XKvgLfNbijcf1aRqhN0367skSWUtsrRR3
QROwBGB1NVG4thEctIBiLY/zT8zRiCms/xie1NrLrKztjWz4ut6astDesxKED4we
1/4En1biHkMQMCNMnZvqhtWc6DFsbeCBJX1vw4gyui46JcyvChUalNKCu2e2+1GI
aatZ2AKVhyDnPZbMSuEAxg5PosAJCIyxNZyHGYJbw9WD48Y7/wpck40Fena7G38Y
noOT9Hm5Xcn1qZ9qELSUkIXhcbFXjw+8dYvyZn8zKCB6dJJdJ/WZFlNB42AimcH2
QdXTxyO9EZC87c+fsnEm7qg0TElYvzntLBFu/kDGWEs=
`protect END_PROTECTED
