`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ1V+CLQ2kDKdUyjWLp/EQHACjNe+WYPtymmrOKIVm5f
o8VnB9tixXXPz66Nt+T+sQxRueJfzsvaC72xJmvnTPDuZaVXuVTdE34hst3ahD9T
fUF15f2XJ/f9A8c+qHN9Md6UEs0GrSpwWtaJMpcc5DHKBT7bKnyJQxu0xfj1nnIV
BWmJ1+1iSIU5r+SLxC2Gx/17/jIvt8BBvd3JAASeSe/UCxFN1CfQp2nBzWJc2DgU
b094T7+k6oMRsxUatHdHN7AaHdAayOKulNh1snSF0AvBNdDkZUBD0lVQZ6s+FqZC
G4wF2DudHyOMMcK6agdB4w==
`protect END_PROTECTED
