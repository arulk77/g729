`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JCxgTPGqJbgkDIJrkHLd++v2pPRTs2Dc+g1tLeR3diLKu/FMi2kCc1e8YFVb3Xzg
JAcCjDDawzjcRs4t3i0MKhzyvw+Alsyd3E5IcMdb554EFQbV5Xu7YXtlScIqXjV1
mQV1TIe/sDh4wyJsRQk1qwRJDbYXhTtN8oHJnNmY0qhasmbC7meQrXLlNycuhlJk
`protect END_PROTECTED
