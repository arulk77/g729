`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8Sa4QaLaTxGpLUwgm6jSLGC5WyTKiVf85P12BfzlH8LU3
yv1kBiyOlYy0a13KxnX+vJGLPZQmHCcH62te7k7vppNsyaUt2p8koMa0gWS4gfqu
hqq1eEvnCUeiK/J+UCOsqOTcI/I+nY/LYMuRFTGwRZRZrlhqGhzU4Mqfqd6ktEdk
oGnI3QU3JQFImUbjAA6Alw==
`protect END_PROTECTED
