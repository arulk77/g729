`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41rDnznS51rjxVAEB9i4sGATLq3ZH4qpapptN3fVuZxh
4XlbArqbnH36Em4Siec3JoawRY6Q2hv2zyRocDO3gMSW24yC1AAQE3IHA23Xm5CV
/hOVg05OPK19sFT2dIOqM4ouS2U/wpxIs6VN5Q+BtDejerXTVBEqkP1Hrxo9iDup
CHikjBradwL1NfG+vBvXD6WiXO/9H/CXkgMG2xkla24XO3Kh0RGI55cg6lg5TfbC
xplwWzN0L5V5puRUUigRRA7zEQ/wlBH01r+PrZQlq9BU80OulDrbPLuN3p9uK1kf
VG+d/5s9QF0vKe2Q2hlBRg==
`protect END_PROTECTED
