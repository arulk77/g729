`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePo1kpvT8LSV8CVXpeqN5EySUpghdmWwBYAD2asAsfmh
uY5S8X5BBugzzK+1Izeu9w7AX6oGEjNu4t3Md1utv1EgnjUydRLSE9v9SfQsVPNW
asR5GKsP8lNs25nh44AZTFOX0SPR1XENzH+QseLtB1bP8K9Bfraz6j9CmPWgrUNe
tP/lGTxJXEvyiyXjTRFw5h/PVASf1LpiiabqEI26fXCmrWq4SYMUQh7wptDKkwSe
+5uEBYQI5zxEZ7SZTPaEmKCOr/c+oUU8hkHzcoOfqq/O3Ksrc07EMvZjXfwZQwlp
oUA++8/+87Gq7vE84RguOvxqY1nGxnA8saqs208L4rmCGaYUaWimI1qNA/8pnVor
xUAyWxYa0XYod/bxJcdmst5UHuZCj92PSB04BY9NsSR5+6yDpxaW2EaFJ8GXs9Ew
7lqZSoC0AIMAEuFAs8CuUXc95xqYwA0Qa+zq3mpnRkdACR3w9/avtjUn5Bwt5hD/
dpIudFYpBPur9gu5My0F9e0WJgG4Fbyd7YS3lwY7JNERXgL3YMXYnTcArqtH1Wav
`protect END_PROTECTED
