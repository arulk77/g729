`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCxKuIpHCQTPFRvwkJsxYiwz61Z/BG0x2adbOTpAHXxd
E/PeYY3HY1DINb4FitHc0paljTW7cd0D7Ez8yU3h2DFlnU2UG4Do1s0RG0H/shjh
XBt3SrAMf7tolF6MhhbI4lme7WvUP5lu5pBqs4uOBIGzVaT5HtajOnjrVdTMrzdX
4/N89t7Uy+ELeMxHnju/9pknTB1r8yhhYizhmjebPIuxwTVEVzPF+8XVLb6Cgvo2
J08qjtOmLeob9MGlE0q/rbyQ55RHksVTxSe0NokW3O3rlFxHz85W+7EWDQsw9M2z
0jLuRGiKqO/HmRMuF1zbykmKkTiL2T8chWCla6FlyGvb6eLmnLzF00lfBTq9wDnZ
3uT8sjlTzJ5sjZtz1YILUaVqFoL1Y+ApEb8zfMa2tY+SUFc8mQmmor5MKnZSF/AJ
Q9XnXqm1eNOpAaUE95mL7azSrtUdf6KNh12jlNo41YS4EplBvbiwNYeEMrA/nBmf
aP159k3rm3VzrIWsWDubniYDjHOoSwhl0slaSNXw3+VETt36iBfMI6Rvr+SOhQr8
`protect END_PROTECTED
