`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
773LT3a7WO07feyQV7fNaWArXSFSZCP/XOY90JNE13cWyp205+71kuSU49iYxeDL
VRhJTMXAULE2IPCueenAqwWvC3pHCizCRV+rgOQW36w3xAjE5Yc1iHyZL/T81KNH
bLJGoN/EJT1JWUZINu9vKiZkGuO9vqcXpDBZyj4iUU2kdUrzdsd9b+AEqBnFbToZ
`protect END_PROTECTED
