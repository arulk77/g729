`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveH5yFFafyJwOSxO6WHvqRH8PcVvLeBR0d7NffL9FJN4i
GbJxeZKPRo0aPzbZgFYjT1FRsRSCIdU+49Yr5WKZ8gKdW7C2GS9r0UR5eMRpmytZ
O56mKWIJrbXjixLZ3y7It9Gb9FEIlZEoUB6Spk3Lov5EXIF1Zki4/haQSL3QAlpD
oOYY7BSJerB8qTNyI86OeUnpL+HYBq89qiQ0y1YFfr5iaspTVvu9BEz0Rre7GqWP
b6/dD+0NNBn1GNk05fswFHdlYn+ytYddv/LJldwyow7EPDKh9BaV2iDP4+uWoct7
7YhbSG9vKBXIMNaktNhm6BKY9L9WK4uojc8fh/yCGZXkzhjzNaSe3z8jG6XxsybI
HNH0SSWf8sMMvuZKoSOCh4nVJgmoZkhg8cDqBOSuK0bpomDmT2rgX7YOrQMqLAAl
kPzM7muc5NpHlcDzo7OJdw==
`protect END_PROTECTED
