`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zp6EyZyLa3u/8rC2t2eJqwjQzEKjqQeLAI/4pZL3jFB
g5N5HUefbb7+cEeU9zyvAvvU7tTEUXwNVQCsZv3yRs8HD0P1yBakTv3wnl7bhMYT
QmxCkLVQr8Q7hZ/SwCZNM3JWKVGr3/glph49SUUB/61J1Czze7hhxBjzE3I3Ha72
Jrim46dtqqAjln+TcfXg2B69tWGIWoumNXpWYfaWHTg=
`protect END_PROTECTED
