`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+5GjgdOYA/AcKVctQSbYVUrDFlWV6/kdavpkcYZgQip
sug/9uxWgNtKVuFYGV0CVY0lz42hhGnZ4K6W+leu8RfK4fRoOJ1fbPdwPr7FcCyt
NWvtHaimqSdRrVEsAEF/RsGh0t8tbu0CDwf9cd3HD6OsZj0SHNZMO2YBFStwou47
JpCMffFyTuBi+E2f+9XbrErk9lpOlBWRcFhCwF/oihlfmd3kcmNQtLqkdRW8O45I
WsDiUoFiUn3AggNYiwutHGm6w0ZWXTwXZJ92W3hbI4DUqBcMdL65jRhBgf1Qy4rC
WmTT7Od1UAWOVQSMAncClA==
`protect END_PROTECTED
