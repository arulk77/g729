`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJLcLvzj/MP6rwIkkqjMB3JwIE0V/XTfJ/QepbZirM56
Cw8NhGP5oUiGMnIxaBc6RD3eJabm5kky//JFP/jCZ/1NK4dkkxZbkEcaGt6cSdRr
mik1L9eo+D/6FoDKDcUfEhn0sN1EoBZqJv0Ia38nZWAqaMij59PpO2MsCv7C2zgY
T/y1hqzdwFb0FHJPcWL3ZNXXQghD0iXKSKXlLNbkk98m3ftpJ8as2X/f/X35qMnT
BD0vaZb6zN9cqj9hwPqdsw==
`protect END_PROTECTED
