`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePpnwQ7yzIWUq2HJdy+NTJzh3RHfqqz8NlNa0/yIgIMP
KQJnM8ldjSx8y78UMGSkC+9lwIvsq4RCot7zUdf+XY5G47jvsJ3jucuYcnGy6ILs
TJXNS46SfCTgZJnT7mON13VIM1YWFRrwPS2+oKfl9FG7KsRN69cMbvJjy9JQ2nF/
DEkw2HraCKXh04RbgrSrvbXGwnOMHXt0xIBtibMj0JEg8+Bk5OzBszGfILnwv99b
J1Kxj9LAsJj9rii8NiGwVkvh7HlRxN/6NK0+9ydOpPrvNdbaQZEmcG3epuz1ecb1
koxHT0T0alXh6WKjZUXijxS4AxwtKbrhVycueuwENKhO6K2T/j5T0S7s7DhyeJ+R
/tuPGEpYwOwHUSdMh6QAWnOrxyhklq4aI65woDuEJataWMtz2WcrU9thgZx8Wa3+
ECp/jOJlh8Rq1O7LbkDE4KsceVZXkn7RWUHebgCAVLqFplaLhmRxmFaZIOEQ+9Km
jEZiwx1+eqaZVU3sL3xlyhCedAIKkXbJmOCe3HC2KzJyyn6tA3rBr9Ku3dpk1yXE
bzlLOxl1ay00GkRl9ShHo9n9TMO8IfiXXwjuof4PEuvtj5S3yXdjpOL1xWC2Yszn
PtxesTNezIdtK0AkNQ0Oi0c0ECWkHr8fUI5s9V+A/tapZ8VVhEonZBjPUpSwxpqO
ptz7DfmOsCiWOqf4X9LCl9xZYmqbf8NTo11TBi5ABag125bYohODzcn4Md9fOx5E
6P5KXKe8pBV4XbArQBYm690raePzGd7gXyToTuKvepZAlWNwQ+VwtpeOiauPASmr
xS7a1VfqWbf/74rTTh4iOTmWDsP5NIDtq1JARXFcmig=
`protect END_PROTECTED
