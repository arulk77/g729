`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJIfZD7giK/PdKZN8667zDIrwnm+lmIsJLcQkrqpKbBD
UsVh16t7p5nPj61jexWzIDPQWXgF6EnCsx0Mghoep8Sh6DqAuh1+HNdahRX17Kb4
hfddxhv67GlOTWxBsIcmSJmVprEqbHLZTyKPkGu+qTq6kDXd/Whnv6Fuuwv7xAsq
EtwptH4iwHQDi6eHf3jfkthwP4x/t/hXdqjnVuRWs0zwu2psue5NBzd4phEqze3S
gsnGfIEu6z0dPLU1CQ6DDLOYldpXP79npQstDSrXEPnBhfn3FYtVeZSSixDN7llo
A1qOHTiPxhbptOAxlsfvOeJxU8YHt+HLP9XlfJBVe4YcQITtaMHPbiKXfX7xcU2z
VWnh9u6cHZgSL7RUYHCm2LNQcQuj9gME+2Ms5PBSc39CvXUkpf1kIzGd/zZZ7MXa
gzK94d95XCrLDzcII8H2wVbZZY/mYDzIjKg+JOdklRU5zS5y5lXeaCnOYHHHIuth
`protect END_PROTECTED
