`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAKODJduhCPkfbMhzfrQlwJeaIAmzeLiGqAQzcXQgcG4
zcmPLD12Nch5f1hhx91GPUOj7tSt81hsMmR4vvYUrYUuwXkzWlyns306gzpO94VB
yD5nLkGxVrEbHrEoOimkmjPuyg987uXI5AO6dvmaqk0hC90+Xz+FnjL85RHttMHU
plhDr0fh2hxuDwkbn8cVmg==
`protect END_PROTECTED
