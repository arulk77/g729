`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
0MFlj4yjh9IKSOmhGQccM8kLKY+Sj6rWN1+LuHOJgbOF7/4jN3aPh1ef6+ABJSSo
fUeQYr1NHTe3zooPBcZhUY/S1K9fp5azs+e1H0ik7GjTDm/wDFMAmNaExwyx0T0V
IfqHgxqkTLTxVYUUHPJs+nnF8AUJ29KL0jHQYdTfEPGSVc4bvIW417n4q9A7+KME
lGyxfBuUuLodi01BJIkt7pIi0jsyjJCtrSZyCDmktW23cee92T3SRprKFbh6j1gd
+phPwS5MMXtWkn2BBJoz6p5zXLscCQRFOKSnd1EX5WqQvizTTwPKshrSF8qKhEjf
DCgGOAX8dQZzmNeHD9BpyPTlq8oHI380BdOvGUc7ElHPjRmugsNT2OWsCSgqXAMk
SMTqpfMNBh/L8Z0TUUfDObEpaKoEYvZll8WIB1D0L/Lhc7XR1MSLLF46/PdTEe9i
lgfwyJ+Fu/yrx7fLaIZMz+qd+06iUZYZ1J1l+xo+HK9EVbyb5FoYyn0I1EWygOa1
V9xhj5CogujnPVIjGmmzwGMMMR9qqkuKhcEm0Wtkv4bGB+z95UePZXp3QlzHpErW
+Zw0Y6ctunjZ63RypXJ5UYFwW52f+0umJP82En/FwcBdWC9I1xPi4dOwdkiP7OO6
idDqWpmZWp0inYAOtaO97piIlHt/UDqx7rL5tDpJsx7xIXHiLXjXDFGxdvY4g86x
M97GqfwrxxfAGorKfxoLWlmp40jBtUc83dKvi2doyFoVQLiuVyULqDiicoSIhWmm
GQDY5aPHdajxp53xWo1AN0mggxGENZPS3G8X0N5A+mbUoAWl/S6ZbyM96QOBL5Cp
wWmyzoPZjilKUFkAwsf/4eXZoaO+PzyrzLZIew/lsGKW3o5hhBmoHb/aFvCp5zrF
4O9D5HZXdIxQYdP0CJqcmBa99OWUxF9Omq0MCqj/CINWeDi+0qvhKjbPleX+KeIZ
7N2f9PSrFFgID8j796no9ONknt/8dkTVzKtjxTtVjixX5I2yrJdKXrF/rXnaEhQe
UcOsXg0jz08hGqbIPSjSB6rnJyV8VixyjYXcmdiKy8M1vx/Ftx0ORAQ45N+x1Bmr
9YkipjL4JAztWmNwGTztYtAdvQbuUcwUcTzB+6JFltD0XH3/lisB/EEE6TiuXYZI
nDImniIGNOae+tXuHAZwJPDXFPCWpsdTDexFAFpznSye+x3a5V40LpeVNtBTznis
m+HwffJYXdvC6kehlQBxLUPoiB1zCYBVNKUE5YUldyNbaqHGeTIRz5AJ8VxobB8k
zDwyEYH/ZEY3lV1+04svuJg17H6TmemivfyjBnivKucTM/zIX2FO9zNyhHS99shr
yb9YqKchbnJjyVQOKSS2AbyeHjPDYT2k1OvTfdt/j+0fMaIns9canQqeFl9I5cEt
1qmOoe94AApHjVWZw3qaQZVRdoTMd7Eyf+n3qGEzZ+xzQ3/nGpNn5QZSFc+ZiO2E
AmTs6nOWPLlbP/tSuj82GiR/LIly7P6vyvhU4VkwhJKlMZwcezFzB/uxm2nIvJSv
MDomRU/qrV6pLrE/qs11NNbQhPVWHofCJFohqh68gFC3WJ+Jc4qDnDsnvKvi+ofX
X9QtlEC7/Dqwt7eZ/rof0J8LuQegwF2W9I0py22D/gX2doE74yH++y/QpDq7eZHd
20078S1YGJbudwgDEkMlEnerwvTPFmR+Pssfs0iCr9l6kjH5Ahp9j36oaO8s39Vv
EcyevoiDNB5x/+HE8tQU4rX4RU2V3D5kEbyOZUpnZ/zsmoI602D3zAGGO+auhV8j
/EcodDc+QvXCKcpoRsn+OmKSvVcOASdxOmdLnH4eONKp5X1UZDeLB5432KN1cD81
YgSbLZab9IDyP0Z2b8NUn+mVDSgzLjPESAF0mEOX0bC+68+Fvch8KtwZLdgcT9rL
B1DYH01JB4sHkcErCG4JBnv6Repz+m50tnTxvjejPuY8HQhi2v0XvSJ8xS6lmHnv
xyHIgbXgZZYBP+yGBSPMhWddloJNomjQkMerxuYWHJRXdGh0zcsT912auarqSiH0
9G8BOP8REegL7Ns+udi/4thSJWCaKHAquvNxt4YWK1LbLUCx7f2LtBR+VC6YCVY4
LkXi0025+oewUcTQ/aEBx6j26BjFMbJGqRKPpkjwpVtcmzovgjXC0GHmTUGtorp7
ERwWIj/PfypBrRygCCVGB0CMsVSqCfmgqlD5h5VPlgX56+vrQ243iI8FYK1/ov0v
GaaSdxHM3GwP+xWNNKoJvnvjwBEmtK59Ek+rRBSjRdisYHbnwjQMTZ/gcmW1gP5t
mq6Uln8gZityw2oBdb0zxUonBcj9Oya176oIppyZbSHzQ4aY0PVQZ24JAPBzjzXM
yOJvJ4QHsQHq7ONmsnMQWtFCPFqvsKNYnum+29igrwfwLhPNZ/nPA/H4b3Hi4UVp
mGi1c/nk6PCWLf2b5h8A4E1CDaQO0LLulzj0WBmIc6YFwmmsMVYsdJw1fgHJWMdt
CapBrly0H/qnf1bvv+bbS+FsG7mEk+rUDeHJ0+Djk1RQX1ZknYB/UXGwKEEABfTF
IN9geBm+tXoQaYdbjlCuV5PQBS8wEJ3u9yzvzLM7Kb7cxueJuHHCC2oYMSjrQvXK
hvIGry3AoDKjPu2bgBEqHDzfos+MB2qqYk5HBACOCi/RwuRVkSnr+XPVax9pO00O
Tytd+sQ+ZJKBh6A04oExOEu1JbM+d3EwOpjyUmAw8MJoAHzSuYiWEswuLslqcAyk
EcQ1GU2zXS7I4ZupLfigVSBR6x1Rbf9NVQ4w1K5baqqYcp8Jfd+vr8ljfl/PPxDI
0x66BxVG8u/e5VqVGgGjbPm118piN8wHx8LdWp1Xv/KM7eRpFbAbHSiuHsXw9kAx
xeCBR/tM2F2PR9lTTX7qd//Qwdb3A7hSD9fVHPoRFDbpofkRDP6era86T2ToPxvB
loJP6oHDfqI1Q/IXJces3/R/x684oJ4AJjeOZHjgzUQxiYyrsSBYdg06qKTUYK6s
9Y57BLRTTnMupoNCmdyLz7zeMH5EawN9keXA+Bl4fpXpqg3EgKm2mJXmH0K1wmk8
6J3Ebq5dXWdeGT0ZrSB5D38TTTBdFhwFSVZmkyY7irHqhsI1Urdc6UeCvcrEjFVE
RZ8KVx54xd9LoQ+Dt9y7LJheEh9NU+dixdEcjl8jR3nXJ82MehoBqLYQ27D/B3GY
oRrrU1PE3azkFtgeqBBtSIQK2/y5j3bUVyFccw7mNF1ZeMGriARWybmO0gVRKVjA
xkBWav6hmHT5uRZ8VWnRKz1Cpi4PqAFGeMqN4oafpRW1mUZlPBQwBzm8dKPRXr1Y
QZ/2uJMdYIMlj+prjKntiQ==
`protect END_PROTECTED
