`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGXLz3gLw1ynt4CBzPsHfJxUcuSdslf2wgqcdUBPMbeo
Avp73opUUgii6B0qb4TOfKVKASJBK5b3i0mNQguWYAasyUj+jtwY3jxb89yPFrLG
SYmyoDbXFc8vUGozfhDVixeKn80wTxrs8ZmFz3LLwIgQ+vD9EMCAkMmmzCvRa0C3
i3Ba16jTHkLq+AC4TqoM+4KxJhYG4NErGvCoGmCfpc1qqkRsjfOTHPX7G0AqCbR4
8eR2MOtk3KFtgaKspzVQ8rDEO2UtxumxWLxbN8Jkzjgc804Mkf9zYCvJbBLXfFEF
cSRuI54elA/Z34CTP1nqGc/bUexdlxo92uZFEOcJDqucIUcuL9FmqLac7P1y+Rts
SqN7RQVJPnWvelnyDf2m2v4jspJIUyXFUnetpf0Xv+BcOX0ars3zKMSQQhxMHB8E
djwEzjp5coYoaCP2V4pAGyOe1eLshgVYmR6Kdktajosa6biNzsLWyUoaGSLUro8k
`protect END_PROTECTED
