`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zOulOc3zVNsg/f/9RN0zqRDLptJGRUxzs9tTNJm4MLv
eFgYvrD9Z/uI6LjiZZRmG0Jhkt39RGh1/DRnNTmoR8oUaIxXGgJPspWJSVVAyfwN
K2hda6pBXs0iznu47KhhW6ukMF+Fq/sP0k4zMwR9P5+B11jgG28iOLyGeuK5E4iE
J3ICLckrNx/yNGSYzz+Bf002CbcOI5C7Fdi1XgmxyEMRmaHYLekaBL98DmRaokcC
c2Z0KzlBKQBc/D/VH9F+M+27LO43vZslJMtubUEJwwhjBLunHoo0D1UYJgQfluVd
zRlNxVt5EftG2O78E3KJrA==
`protect END_PROTECTED
