`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41mnpgA3Yc/bV+9AMD1FqPN118XkdrRMHiP0k1bBKAfK
58bnKMmJi3mQcT70Z4kX+CYN+4f/06UyuHr9bnshScwUrAwMEdUs0etIHqnhSI7E
EEmoKVEzwx3CD4jz4DBpnqsBqeGj00KIG4eRRiJEwaMPyixT06fePZ/+inRPynAS
VSW/8mKiFpjRJYq7+Gkr0uydMr+9n7PGKn18/u823t0=
`protect END_PROTECTED
