`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
hU7iXShQLVFcvSQzrfwlg29o0BjAuDfaHIr1gKGU4xGyPDSO1vq1O86GcIIWKLzk
O8TuGndThMuHK0kIQgzjulmAg16J30b/U87M2jtNT9PtCj2NPzdAFoXFv9Xs6Oae
mnYkUVxSkSmM3eUCE7Pj91PJcc2+H0oQ3cGi03F/qLQmA0Kxb5TcknkBoCXEqSfw
D7bdBExsYS8QOuJV4jdYsmWomEQj5Jxa2Pl9T1YM97D3Pn0LV4tEpIQEdJ/cyhXd
Q2itO7uaYAFBQGM98369tmsBK+Nji/A35Oq0sy7cv3M=
`protect END_PROTECTED
