`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHjy2jXU2Lc/DRAJPV8fwB4J1Ug1sAPC5JhxMip6dnA5
mW03Tq/AR0ODOwzkHzZ86OvBY4kuIrw+3yNtzpDwi9YuqDos9FhxZUA+c+4CERQQ
wTzU/zZYW4wuQLhhAVV/CY3IRoZ5HkQJanpS8fgabJJi6AcoHTnvad593G+Yd64+
ag+j1IdM9Uj3meSvq7ripp4Wyr2tZpy8jTECYtVKf+buSmNeUGyvyHyBPqyRkU5t
XSAUeXPs0U7Nl0kiUV7Jdw==
`protect END_PROTECTED
