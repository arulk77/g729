`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBbeHIzmnSBM5RnEvMmpHcW9s+NA8vpFeiF/P6tUTEs0
IEO8r6jEVGq0uPo6NTpiWSJNkPMue3PsnzaXRlK6bwHlH6MuZ3qldpxC4WS2FaqM
WkFiLfKTQukrFeOuRlF6n35lOKwlmtm53xLv2ntBa1pYXiTwBWxot5am+ifoGV9G
8DUaTdSzqOOA8Yr1bgJ/zA==
`protect END_PROTECTED
