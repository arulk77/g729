`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFfTE537FkBpaAzdjqBKJEQCOFA2UlseEBGpMtzLKQGb
gc0B/7anxyBTloVMIRthDf/oqoFYPJ92GkT2vsbhEyBJvuferPTywswd+0gcAGig
Vadmz90FpqwkXjVe+so9DMt1dJ29ZnkCksvQB10izT6CVvhSWmJ9llnhuxayPHKs
aX34zE39gerhcLKHkosr1umZtwXlfU3jXpcZ2nT1OSpR5e8hLlGBVig4Y2MKAUjf
ahS/BX/7n/txQ3wVCj0Pl8OxamlSg6u64KYCFCtVr/omsPj/x2/G8ulxUhb3Vvoi
e7YrvdDhAxSfA9xSNOe5Mp9/Izb2vbW2pMuznpbg0y/ifOcvSUS3HCSS+8bKAhp2
Uvjm6uXsRbQzJZacAs2iwbUxlO7BtVGD5ya+SfqpcOTEzIOKCUaGat0cqr4LeIpO
Y3irgupeuKTCPHw3HNgoibCOYzHYuyWbnO9s4UTEOZjnAuMo3miIm5qE8N1HcI46
`protect END_PROTECTED
