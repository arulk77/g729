`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNWCTkTMA8ob6/OGnwOKU9QOLA+Hls6a5pAPotrcfINW
ScDyCERmcyJeX6bDwwBZ/nAcZJIToCKmIZSP9hvxdl9Os5+n1M4KUIgrfB2vkc3S
Ag+tQfLlt1m3d4DYlbfcYRbinySKGfwcuITEHbNqGSthWKIOAKxti6NDIin1dDaA
w9mDkVnalyRUPvuqmmHhfcQ8LdMJlGRV9ti8Y2lZdng+lNd6wzQz55Uets2IBgn/
Sve/WSZz7r5FUmTf0zhkRL718r6svidNM6jXG7RF765Bsk/zhtWVeBLoJOU0KZGr
rzZMO4l3bHNfKflGAGlmMA==
`protect END_PROTECTED
