`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wdkLGP0Md2sd/ui6YyK0K0YKI/z0+Thx4RQ+BK8vnkI
mFvwbEDUtQn36zb4beJjBb6pLQEsCf8F3apDzACnT1wUSqh43QHmPCluzLkANHhx
vAFSL+lQxpn7kNiLvc/Sm8SgFKeLyCTjnyuWdUKz+ujhVweI2Nxww9JjKiDM5eo4
7aLJkO0yx1AgnGNWaLYABGr6rpBjXFBfW9o94cmd0C66y1J4jLdhWlwkDrqva/jZ
oSa12A4IPQLtHApCyNEUOdbW8yG9DubrLebz9uPUtgs=
`protect END_PROTECTED
