`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJxh08JRLEzoySFOyQJJgdes3NMlrLPKh6O7wmxcq4In
GowGVjpW0GbM+QciA6CI6F5YKkPtRAJP/Nh0Pe8l96cSQoecK/8GkrfzCTAzH6Pf
7V6OiSl4K6v5dh/9Ab7kuZOlQ4IbrbOOuGjYy+UyebjKP09Zs+LMaFhkE0h+VzO1
uEi7FzIllePirxR9CYt5XzkBwylfPBWCvLKqMCLM2uz6am7kprtPj/e5Z+xh6971
AHpa5d21tSxPMrCGYPxZEEi8zg5VjJS8S6t/WyvYtSSsvqRLl+ZhNbgo+xTSAh3i
0X3sgld/R3EgQUD92oJm2WPwvGDNcoV6T8k0NIvp7JM+GK7ALmFXyz4oRQP1onrz
9gZMEnI8rKRPBin1SYBY9kr/WJBhUFrzdjfM/955D2u0Zslleq1q6iOHCctazuQO
a5AL413AF8Cc/3xkTQpN2SL2QJLRRvLJZoG9eB+TDjLz2gtk0PjlWOXDLP6WLDd6
AP6jwwXxGTOnQeOT+5zRjv0SvJanha5lLP4oOKRKMsfYD6ONZBQxXDXCBYlKboqA
d/SEPj+TmNw5ArylQORxow==
`protect END_PROTECTED
