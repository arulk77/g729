`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
WB6TfcMUp3UtzbnwftWfTvI89czRqQdmBh01MvamIw0l8O9wA8DA1fixrhuUX6O4
2TKSTwKprxfUzALOIru8gXtaAylagknAqFIAA+AszVh+RnA6BFDRxUtpMkGiqaDB
DGfOTbUWP7G4vnfpIRtOqfmRhfysZfEkvQ0nQJrow7WNzQ2j7TLWD9t7+T+jJU5e
JbtlGmuTVl6GGH3CU6kZgWgDDx7xswo/tRAo1CBCNhGNLniRfD0RFYvUU5RndKLL
kIOyxN9PSEGPdkn2yA/PLQFD+Z/IkZzuEWXvHIR4+ODRBchQAOR2KqD4Z6LUGxYB
QgnNsKzedYmoYsxkTMXgLrsmNmVnKBzXZp+R+S5SHfDFcD+2OY1OPNWErCfEHn04
9sEaCLMPFG4Ljfc6/KwSXnamQFl1zeoqWsxan1A8omPxuiLs/YSHk4O2rzTEdU2k
eZ02Vi5HeOSWfotKqGUxz9eiRZ7/oHdUmaDWM12mYU2NRNylRi8HU92px9i2bJaa
tFCWw5atm17lmPHzW2PAY4p5ug/0ibc4IJyvQAeEZRIu1f9oCAUkLzaGzw6ylAXC
SYhV7dPQD++PitNdOihInN3CbXCrsXGPj7ZeuVf9NjDFCrrjDNAHkCLsvzhJthTc
hracQd4QLb5TpxS6bJSrYmm0/IKrmQGl3ihgUf/rBqxxpVArheHyJ/FK14emfU6y
y/bObmXN+R/oj6GilT3pPuW9QLBDLPgSTBM/2Dt+6VGIyJ8lZgedeuwz6804U6fA
`protect END_PROTECTED
