`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHy7TjFz8AxuKTlb6LA/DTGWzON2R3oD7EjjFOXRLUF/
Pa+4XEIzGOuKOCRuSxlf5WgjWK2IMZ4h+dfaPyz0XDFh/eDNhOnWlhLadvOEn+QJ
/3DRkDo0eRjJzXawO8OD8N54z3NGsuGEScy3uQfBcFZa4PUswzODNNLgNwJbKL0R
wjwLirllny+32n4ZnxoltEjexhYs7UMdFtMolxfnxnzdRAa+bYyHOuDrChgK+C2a
7CLwAMgh2Wx6oW4/JJjp9Z+M/8egl9NQ3MaQWzEMSnHFTA0kxml7jC+cnjApUc3b
xS+klEySgZC6o7K4HRbes3fBmyXkEMraL5yaNs/70eePv7QrRPhYZqaHb730t2Od
`protect END_PROTECTED
