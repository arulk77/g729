`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMHId6E/dRhOrB6HKfRLhxcxXFtHFAwveYDy9pNK+pLj
Fmu8dhNdgEtn8yTw4QU2zsMRdrXqpxmjJUlUdvIfjs6eX7t3/+r6CHX0hfwP66+R
kEuFPt2hWEkjFVmZgNeF5CQEYKkODYE4HmYETugjZ4gbAI/rtFrf34JdrGrc1Tqs
+rBKhKgQM93BjcWpfcX7Iw==
`protect END_PROTECTED
