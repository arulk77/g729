`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C8/ReCf/IaKkpSjQXIWIdJnLCoP2NAMi/yIje7OatUon
+8LVXnRzyYd170zy86vnq22zo0ZKjiXgyiQDcwtzA+bpPCvtV4PCxL8DKxGyHrpE
6ugM/RBrjPmsoPyuyn6XTt9wL8bTKsWXUG+wuYIX8QARZJianj25NjGUHmUgKFT7
7ta+KPpg/zMdkECvi3J9AAyCtEhcoAjk/QC03a/8tcadhDRnFXkmrtgNPgc2yraE
VHI7378r3HFNp5yG5ny3fqoQJ+ZmNLQa5aMd6/BpL8FDclpRj4yIZQM/kj7wLIrf
GyXrc2AslnwbaoW6wGR0hc6zi5B3L1omh7tQhWQJ22TWmer5n5hAeNmMA8QEOCo6
mltUlM5DzlwnldQq6KXMGi7eGFeHkgBiyvT9GuKHXdKuupO7zedFOu6Fu/cEHoeK
7/G9Q9oKB3p7HeZ7nNSjF6vsNPYV4z5CoYIAm7NoEKMeDxAtQYLoMLNofZDnkA1L
mo+F/q0BNefvbR+Iz+Ujhd5jGO04eqoHXc2tSvH0JKTJTONNfAz2Y1DroC9RCWuX
X1qaDJ2PjPeolLl5eqKzN23Xt20LDPMo3jPnHp3bs1TYvd9TXtnfmmafVB2OiZXW
jwcV1Po/ePFb/tWq43REwqquC4JzXBqO3pgV2So195z3Zwy9yrKJwCdI0uWMpahg
YuBZ71bTdjW35cb1l/+SLxN9QQEY3RZDi/qDphIHDAteV/ydt41LobOMFaWtJjuW
6dpsZbGqGjJcSTttUOI4WBM+hsiLpZjyT/857B+3PipEt/a1eryqkxpfTScjASKQ
XKAuqvNeAS0ZR1YG5c2T9pQ7ZRbO5gvnJc0QrrAP8Qd8QYlwi7HlyPXyU7K5cKq6
9s1MN0D2x+/LLxyTbCsGEgdVsy2TFCoX+LVCAiQUvE6MMMqnxVreULDeZlUMorVU
aldnw5BcB8cvOEBWK+X/Y6UqXSb69LW76ZEbfcRX4sKB5VwkJsnBhcxuyu4FysaY
IOElAzNUG4P6o3Se7mqjXay4Bpt2u8326w8LWy+VfAK9t7Z3eR/pRUmy0AcVn6Xz
ANaLkX9W/UWwyStGwdHr5R9BkTZ6caIoUe0nkMhhsPeflIKPXkDKLEYofepgHJ1u
EUpFxiNDvhcXnfpe3cYbrjRIAW8PkBJcFCLzmx247z1ukmPs/422P49kR/znwxwh
eJx/69tGlV4goy4o39i11LQeb6b9OYUNN43SsUPb2bZB5cjFDEAk5htHbboAeH3V
M9QSgO8QC47mgjnkuEnyDNO/aKN640VRVyi8k/rNtN+s2YE7c/xg7DDCpixjXgOY
IUwBsDPQBHTLp8CmY5Mm8a6qx+0Q5O0qaVG0iWzcTk3p5DSvV2oDeKTKqiBifHP5
UnVcH/rc2cgT0T6+vsVqle3PgLXib4562q2OH5I91jHFUJR0hq5SGmkQJ/CyAEhL
T/3qSg0QOeOIlVgqd7UHo1jHoTsvKI1QrMmV0jef/nxZhm7VB1GzIFqLvjiYkJgS
u6JF0ouv7y3lj+4EZDVJPhXZy+i8622KGJvQuNlvP41X3w/VMXN2ysaIDb5ijPhg
3VijkqhTinRnBv6w/iXwRCnzbTHMi77e5Y/L9iuSOdFsYgfqvWobOeSVBFIbZByJ
yNpZ7g4kFYKpRdja0WBYZMxLIZ9/0YbL8mY7ehvUfqn/cr6n54bZBV/8FWh92MVL
sgYsjHO/9TDv/loHeiJ9vLWjn6lu1wu37NJLReJXZ+kRuIAnFXjSBrwcfKFsTTVy
1BPrJ+3V6YSLGfm8sUSIqdDioJ7rUgUWpi9EVlgb+ArZVCDyixM4tB9nuDFeyDC3
eVHffpcXnrYEXPK/qfv2SOfE4OmRj0HN3mC7dAHC9lFhUegUBcIepIp0axkCEYkX
REiMJVRtPIWZCQjmRcjxypVm9v3HOMqdMefTMRRtPfrssxwY/KBYuD6YY8NM6DFJ
0wnYhbMM4IKis2uV0ubAPYbXZcJWx22Xb2nUhD1aGrn5OQS9QiqJpYCj9Kntlbvw
UgZAyYUKexOhO5BYhcLLUFeEjqzOAufRpqh4tSkTsK88tDawdQ0E1NdBwZqf29Ce
+FSpOHDyfuQPkFW3Np5HIFJptcN9Xmut0zIF60TgECHF9JgbzZ0mShecTCcjz4Q7
0shANoTZYjQvsDXASVvMMU3O+4GfXfIrp2mlJYI1B9tUllJWbWy+IqjAb7eP/lE0
ae3fepuA+LAx/O8toXW0rFRJQJysxaeuTCOvSZHa+x33X3enoMUtuK+buaLoU5Oj
bG3ZpIFKWY8SWUH43YEbsC9pk3sBziMfgg2h6dYTQZWBtibNyofFaU2HKx3KIPqJ
MI5BRT+0Rd7mzblWUuUAikJgZYpkUcETc2riGg8a8unZhtjkPnjsyd/Gh3Y/bGZU
hP86gIurVTRRdfr5f9yg0wKgLzPBWqd1C7QQ8wzEDn7iiAHjeg9zxxhGvVK7uJE5
zqA4srchblZeFZdstw6RwRVIt6e+kpUN5fwoP16B2VmLufRI7IPHAO8d87gfBuTl
76nBX+j8IpIFXyzT3VQv4D0m/ESXMvHDAa29SVfBbXXPUFFatNW8zDbhHCY7yiNs
R7DDFbbcCO3kxFbWafILn+VYztC1CRxsqqA9h5Zi1ywrgiXUQIoulPMNlEViAOiB
B9wLkyMZwvyyqDkyB12bsGEawO4IQ0FjwbqhVeSezTMUgKiqDxF0KJL26ywmDTRB
3rOEO+sIPVFwsEdte/G6yOzh/gGyi1QyIQV9rGDyoETo3bzm5Fd8MhWDoNWEBRTB
xjl6qYG6zfRdGJL+0FPAFNF0S3ak+8cqKoXbUr1yfqRP7oSs+hEY8xj32jW+7Iid
g+eKRznMypDoCk7usB0htC2mzv/s03dkV3JM8JXKRrOZC4g5TaZbK5uI4YgARqYo
dsBRO1s2aLukW9KDh24u0GD4wpTlu2nQx+UUiDq30sUDduA7Aua4E6l8aLK6c17a
AYsiXl0dy2JsNat7sFW4LHJwswyjrQHaOpnHybiyx+gBlFgSUXJkBLcr8NeYPZXm
0+EbQZzEpO3QRrbigcDiEYD9/693HVoYWD6x4Hn8x5s0jdmM5cOnwQ7WwZAhCMao
bbafq/LzZpVfkCQfvt322A==
`protect END_PROTECTED
