`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveA+s/BaojiB3IifO/tJfXtpNeFShpOLX7BHo8vf1x/F6
l6E2FegepaKUhMxxMo44Io/z+3LiHksqFS55GezwU3SRoc+HUiVgLwaR63TWFtTw
X9Je6mUg7/nVQQCSLgC3RPEMLxlgKRUlUob5/fgieIGCh5bR6J5yQ3vkuPRIur6l
4gTtssO6wvnZK5XMpM+fcw9S+r65e/r5ZDUB3f4Q61Q5srsPjl2gMxc9kRdzkh4q
RocZd4X6/p63STwC3Y/lcW0DZIl4sIPfXKHIW7qceF28T/ENWL/CZHraKD5fUhBi
S/CGuq5G1yqMN+HPjaHS7Poky4LXpsuVSG0Oul03+vNuueHm5SO9rxGpAzCWkjlH
SX+WxKbskH2PyO6r9FRN3r6Tk6IGCFDmUUP/u0/T+Rgt52vqdJgkCbQ8ag1p++rQ
kdI9PDPuGTh+xYq0mytLwxvS/XzMsxLjELrkZqjXnc3lcezMMzj1jjDVfwPE3TON
pL2eiNIbx8sFy4E6BFgaZZGlYisRug41DECbnU7WAgzxf+G60kbXd9Ije+h6Y1NU
`protect END_PROTECTED
