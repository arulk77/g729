`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
LMSrLwmaE42X7Ko2szxXFzHy6i5oPLBU81DnF+cqpe6Lv36Op8ruZVLrVQ4ckf1K
WVygQXO1SUorYpH5jHmELaOzo9sE73rF0OwiAiu59KicmtQ9js51kO7CEx9ypJ/6
uOwa6us6AteLy2PCKfgtkNkiM8QOT9s8trLsKfXd5/G2eR9Rt1C4QwlQsQ70sqOd
1lCg+tKF6Yggf0XmbimT3GKOu+BRC+uM1MWyQ62YZyHt2xgTSlT0NfioyiIKOVV9
6iOUrFNcPm3X7QKOq5qB6GeIo6bFy9bdCIZsl1SyMSbsRbbHMoDrTkZZk8HTZu9M
2SKSfxZpoG6xx9c27xI81+a4JU/vujy1zBif7q6omoCCP4sG9RsA7Mr5tNYlLP2o
2ZAC6iJqQac5Fm39CW81aXfZTO2eRAhSogd2FuO4OC00Fg8tfk3/z2ZenZ5aHtNr
kT0wRKAQ9l9kycLRKk9bMw==
`protect END_PROTECTED
