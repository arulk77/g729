`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKPv8p3ZB+fUqbzpuGKd9d/K5SE9verzFmgfcQ9OmAst
lmqpfsOi/ni/5gVc14WtH0HF2msMgc9kbXvXepgHtDgWOC/XY7CEJA4/CljWecLH
ZkTkxu2KC/BrU2sFiEO0Da/4EgNlafzb0B2buq0y6BIn9Hlh6rTHlALDXZzvN6Hz
GGJbKOxcesGRQlIAMMr997ChfTCHIMUA8k/PKOgHJBKNvhvlgi4jXdRrSeYaImbz
cxW+xUB21+zAuMa/kZI9spuvGscLULhVdvNXN2KwoAuvomqE1C3yniXU9MBk156a
m3ID8faPdb9F/udpwYIrkg==
`protect END_PROTECTED
