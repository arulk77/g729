`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
otPgsHEjyWyaUZ9wpgC+VE2F3wJLrhra6fmlAWcWk2kFKymd1vTO7s0laoki36jS
ZIQoUtCAzsOt8iFJgC2T61LOe67msKrx54I+Y/nrEWQX2POcfLW3IlrfohDDztkP
GDfxc97WG7hIvJjTIxxdLoYr28+FrKvTQwhMcEbuJNRx3rXG9zx92ws7s7hrAv8l
XHjoZMP+HsYgHbrxpB4Y7BYQmIXZCNIYY7a7YkaWqtlhpXsUd2+fjquLzWZGEwxa
K11QJei0JHKP5gq5PSyHxgvu+Oq+10JrEofHHjhI8WRXel4wANn9NFkdEA4BnnEi
yitjy/y1vtrKqW8Z+EJ5y+Dd/47drNFrLOQgvLQEpw7u3qTcZlDTVsce5AOVtogh
Iv5PEVfv/YO12MLBBTeI4L7Stp7vufq4W86ndy2sWWalDqBO1uSRUZyFqbGc7ZRa
sOm6Uuz1kIhWeE+dErn+mMyUVejpsrRYxe8fmtfs3CreKNUv06/tMaRJMqHtSc49
Q13+f+jkciza8owmDFGCmbWgnt4nTR4S2Ax7U3gGzKb3JlB2RsnRoTO9OS6Wad70
Bsz09zDxD8v6TJLKXs8mP6YNpwDjYQRxjLFX3fFLTK8rOZ9NlHcM1E+z6vE+vrXB
aTj8pOklEEgNJbnbJ+DgoBKuv1brfkSx7NWJS6WCDIMvgq19aLg4E7GEv9VnMKo9
I8W+MEK8e8WV99u9ee0JLiCTpTd6bv09xbQmNv1KLmYpc555F/r6V+ZmDG+UTc+p
`protect END_PROTECTED
