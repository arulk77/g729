`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveA/C/OkCN+Eq99Z5u+UabY2Cbb6HrmXocaydHcagTITi
1mENG8V9KjpyHInM+6gbCQj+QVTRVDCGGnj3Grzxv23N21kFvYaFY3Tbbv+NU6ib
FDmDR6DOj5Rlr8WgUopiIWwtLEQFQ6r3NydQGEEU6PdgXLyewKg48gALVJGpLU+z
LQxhuvhE2HH7Sk9LuyV4KA==
`protect END_PROTECTED
