`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+seDB+EcWTVFEQKQ/hVIE1/Xb0YHOw3HCRwj3vYjN20
7W/eoIpNqBuvYsU+1Nfk8j+T5F20hbJTML+RBWaKiPaZMWwbB8SE1RXW2Ys6Ai3v
aXT1AlJMChCegqx4OdSOMjWcmyRYxGv7vRaKIUlRXessFAdFwiYD4Z/h9Io4DPvt
VB3m7pDJAViFXldEy6vSl8nFJxDhn1pxOfvtZVTSimGw62DvxPz5LBZrLbbW8K/b
5RzwT/6csy/rOlbWPNW1jlW/Ry7yXQgx1KLB+13idyY=
`protect END_PROTECTED
