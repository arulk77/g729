`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDzBjSudmvFc2zQpuODxXQ4BtXoJOIk6wih5tZN5dXm4
NeZtEW3GapC8XNzWuOT8pHCvx8Zqb/1pOlHir2Ja2iSTAh36Sbr6NmbBdoghiKlj
FvXC2CRylO9XnabgdrOQS74dK4JVvVOxK4Vvw+9h3pz3r6jIrtqHRU6l3ImExvzb
ZK7z8gkG49zss7MQBq3eDa+egQv6vzro+7MdfKUMKJaHOQxBbTd2SmnXugk784wV
FfRbGugFTpfWBT+60vLNAc7ue0PLNUq2amcyWWb4BJIDFCVy/IZ01v96/8HjArWG
BQFCoWwAt8gT0TLggef9QQ==
`protect END_PROTECTED
