`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEq2kIDnyIU8EaKSUNcuU5/Dj89EmFcBlXJ8n61jD7QB
rgcOV/UgMiZcqMH3Dva9wKvgYLeMx8I+BL9MAjbJRnKTEO9rKCPEqjs/jMWGtxyJ
s0GrN+1cEyBVrSOiH0n/rKF9xwLBTR1BJ2NViEnKtRvubVsfDdkzEd+Qh3Hrf42I
Ccy+Lp1xoMTAUjy5Gv7nLQdNzHg/8XuCPwhPS14fLNtvDSQqkbCcww/pJCDOa/5E
Oy1mfuJ57SDdvpS71PANlz4YoGY9ieJZSmQOmA4MsUTsezScJkite8vvw0ZmOuUb
cHCm0EMrmX7JghHtlNpIv6d8d2/0SKiqJWvnrS2sk2XaGbzcfKoCElWX2LLCoOq7
WFC9h9AtaYNOdJnLjJYg5gPD0pBHjt8uukvOWcKjv/BFYlwJXCJGit2ukbK/QZKE
oMQakr+7ifY4Yi6HF0lwihRB19lVIIiVRRaL9acKHNrlONOmVjdgoC40L93g8jWW
`protect END_PROTECTED
