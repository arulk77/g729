`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFzGTGdsxC3gxJvkY+4dPe6pONxO4cnzBmqnafNI5DxD
D9p1aOxeKUfEd22kmCe7k8qEiG3OxY+i7w+XFC0pnA7pJT3QCPZkZpfIH9S15ez/
jGfhLKmGj15aMwTRTya+k5n44jen5SjIiKVTU1vLBSf1AUeWr4mLjxXvGyN7dbdv
Oo9uH6hzPzYYdJESDnw4w6kOai1QRtUDhgirZZjeo+jRhcBzTqyHgHZ0T83DFXwB
2KB09QxbeAwNU9K5/ZGAZkYfM8tjVKh0gAWoJ+JvKcvx4WCWHQL5rS2QI9UNmOyK
aeKhDRgPCVq1hsiWz9mqQ/a5EGYsn3rMe9GdiTE5pN/rZQU9q8GCBIZM4nNYBPPE
OTrC0s106mgvegBLWRAx9t2AZNFnUwV1/o7o51CrlVXykE03L/XzTRHAXlccNEk8
50DfXyMYCHV1H84+pnBE7POrdrmzqoCOC0gqSNiwx2/hoTIYirJ1++tMN6pt+UcR
M4EX+LNeh4A3/Iaeqj2nZdGVYniVFeiQ5Lt47RDajxcmGY9NCAP6zQnsZUMk1CjC
G6H+pOQaFL3fYKiEIIa7wg==
`protect END_PROTECTED
