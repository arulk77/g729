`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHAiLoona79fivs127ZNx0FoOSX1kybm+7vXlGxzrXMR
QYPQ8yp+hgvQQYC5x20C99c2P+X9grm8068hf+QuL3qpK5vOPHj3mJzzsli5LIXH
70RHjyXLN5OTHpxLUDJoet+oUSTmxhmVNscG8fPLOd+dwrJs7DEhBVWJlQCkCY5t
7OUIMAEOvcXzvOe2l5ojMUOD7YT+kqbdT5RqwwdFo6jMeoFsaW1w78mbqzUC851d
b3cA9VxnkNmvErn1RChD7PIUz7KFuCWgVhK9ZVjAspWycYBUAn8qBMEUJsttqDvW
HBx9wBDaow5LkFcND2PNworN9aEag/2p41UYwFjjMh4NBZ1KFX4wLgouOZej6JCm
8+yraLr3nArdGUlXmJnJbXXMdiiCH9FKZJmFgnbnmVk8fl4DOl8ZT2/hXwT2YoIF
8Y1S99znJyzLfJ1ZOYFc6PdQOTIw7FN0IektPn/Ib4ljc2rfq6tGu0uddAzwqOIo
c8Bra9GD021trv1J7LyNGHnATH6d+pej5dRkuCDjtHhpmKgo0zplbr3OZpXyAXg/
`protect END_PROTECTED
