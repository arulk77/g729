`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
WqburvlC15y9F9C8aBkk9ub6JfS8/SMUFzt+Ti6bZx+OgfZS4nRE0WM3JWR3fSsg
Rs5eh7/+W238kT34S8SrUHeeQzjN6faMf0wcBYXyI/33z/chFx1JgyDf9DiJtMJP
fZT41NJ2hi0c9FZt3GSvJH0VB++5SzIXmwiZ9tGg5iS8K6rfBCrxFDLeXxjR7ChJ
`protect END_PROTECTED
