`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIMHW4bSH99frsNzwBASSpkRQqMKDnTr4tYukXXmWu1u
87/y9tKvm0AEWdpis5UIlRkEd7TnSJ2CXDWK61a2TThwFNqZNVGfVBUHyKIIQ+GG
u+kvwfu/kEkVw/WDDiaBOs+4OzRn8RUtWQmxawC+Wc0c7rrmCik020Bhmnr+TF4l
yCgIRD1azkTKsdFTAH9USnEt1QCn4tChlzgJJyEsWvi+jQ8iMcLaQMhx6wCxIqyY
M57LvFU7bGnBYH+s4OE3iRcZb/Tov3rSuJAB2lSclAuNlImvSZtHgyTdJK61lVRv
`protect END_PROTECTED
