`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAfSreRtWcuFVZ4/20qHPTcTVCsCw2XxVUIrZ694bkHAY
zCp7W8MC4UD8ejeWoXdPxL7evr044/OXk7LuYcVPlVWX4/5u0HL/rntnOxlk/xiY
QPSPrAwBTdZNYxNTMKg+/Z3WGUzZ1ddLo/XHkNnFc9ahISooAuaMgQ7lv670ZQg8
FDOMWUhH1Ly+Bf34xD1OrP6cJzCkcKxQ5aWh5LO3j58m/ArvGCIjiMEPO1ijjh+T
5ILQo1YPLK9jeUr+9Fx67F4ENJwegEp3/cbZ0q6qfQX3sGdl4iSLG/Mn6XCaWEJY
Y+fxgBI8fblc+ASKF8zv2Nobg6jAOYQS+rlELW4/7CjKokY4Lr1q6ZQuz/1rPnO7
EPQ2pvl998VTOILjQWTA6AGB2PXXcdhpYSBg3n/s/pb2W9SJdLXkPL7cNGiYQdOR
20bSNn/jwsXSFOXbniV4x67csnIWlDIHd1UWDDBawrLocYJv1TFYa8UpcjLzPMUU
JAYHCY8mcYTEuCLKP5DL/jLR/0VIE20TfKuxqs+A31elKZ/fz+NRJdh5kHuHhDMq
ZwqI/2yDD1sAbFevDYcZ66xVBndLfu1H3FWxj4GTooSoQW4UDv5ueAbYJB6m27sX
j7EmiNo+dFSbRvQpEXtYkuXtBNKNDVEcU75aOIZx0cQZvMK78yS3JVveLrhNHkBN
EuVQ/lEieFPMf2niHmlAzys2cRfYdC4+KzqQ6xlMJlJsI+ggP3bgXRt4nyUjXCYg
24VQd/GV4++8zAK7/MJ7YVqZeHuNaRER60noeGX8MlHzrdTRnRmxGV5WZUoRpnMY
94U2ytJrWXRfrXumx89TQAa/dW4lkhicxuQQOFb6CMTBlW6+ND3zslTTnY1b7MoU
tWJR5+ZEewcPXA3p8XhbijceJHz+2IQGmv206i+KwQV2zE8+1tfZEyxCm86WXxSg
7tR8vI7jXNARbE9vbQVgx+GHeePfgEAgFmajYPaC4VWOm2CA7p1A5flBim3pvpTk
KQIN9Kbt+5u6NfXHrBH03byt5tk/nQTANgMdXxJqiv2yMmct5XJy2dOvNP100PTO
AA/2XjdUjNVWbjJ8eYxNjYSjrUUFXZDh9RWC/GIvdAqQwWZpcf7SlM+aP3p6vw8H
5kN3VwMoRryvtD7FeeZHiGQ5PPK56mKDhVmMAagrkWgUtll8td3d+rIUq9p3bdWf
OEELhBAs614QqC0ubutSYrMD3P4eW/nN/tLngSKRpyeccd6tb6D9+dY6TeUuvOFm
VFs5sOHrz8LM5qpxyxe9KqvFdkTaLRXKbqpa+cMxSflyqrRybk34+w1ktygdFQbd
H4D6V+twqAVMqV2uciEtc/mQa62SGIu3bvYudaQT8TgkZOnr+dSSADJ5F0ueGrEy
L1UivofL9kMUyCYoH3lael7nWeuJ+fwId4maF0dx9JsMcgdCv7qinm9FeIlBMrqS
YAoYSMlQpem4HR71MkcXlq5FoV3Ovoy9MQtwk/p/mAowSS1dGXiGVcpAL/Mz1O7B
jyWL457hVkFscLT7rV2fIRpeMP0El6MqumsYZ0dAeNVxAuNPKvy84zASs5NooE6h
0ZOqZpMIIeU0Lxawxkot7YLsKfWOC9sLkITzNGJuHeK64SFpzCU5/MmHJE7HNQn9
kx7KZ666WM4J1kJK3r4dBfUNV2PijHCXfxhSFOu206OPY6WwPdVndtq/pGOcTx2j
yexwMtq3pVGBFt3Tjfz7jF7gf7K51C439j3zpct4bt3fpOyO6xzh+jJYlaW70lJj
fh41eJ/5g6jSwifgtb0TCpm7eS0GeAFAFrUWboCHkMXXkvcPUq9sKRhSvvwhNNYH
Mg4kMPCVuMuzXBGXjcfWkwdExZ3CG8OxcGp2OEnmv+m1fObN9aJ6gzmjTBLHIX6D
rB1WQSHBHoUtH+VkKtcxD2urrTOo+2VIHm73MfjaBcjq5IFn/KMiG2LaXrx5qwe7
2DhHgB7jcdy0exVM0PvRO/GyNU8+vBssU0W5bYtN2h8t2vnnXU0Yk0zNqxw7iblG
uieYbcPqsSdRrd+dbJSrLS4JIVwUIFRH5TH5Bx7ceix7xrKl207KXualuoWdg4+s
tPWllEN4GjIZIx0szn/S6zqrWYY8y4WKao+q2l2gsmioIsRVgoofgXNK8DtHoVSc
xxAUZGM5SXyYHUj8QLQ5Wx1wUuQjHSItNJPu2zi9csPa1AA+xsUTbzmYeaOJ+1bg
MswRPtgLf3l3uHlMrjgd8CJnb07OxrDamBc9rBQn++aJqXouyQUHn3Nh16uaabnr
Js8z47HVZyQWU3978Y0sEs2xM3RyxYcB+G3dE5RWv9hYd1aa0zBMOu+XLsSd9eoy
TpxAEjfL7wHzWUtHumTeXeGXgahojmSMwFXDOHdF68fXxBkORyVPOb3Y6CRZzPmm
wPUXgf+AgALD/Jj/Hf7zCGClKZQeam/TpGMKSyJyU3qsvPhDfoQqtj3uBmHxV0io
LqBNmdoExLi8HOdUjnhYdOeBU68Fia5+W0ih/82UYEQ/IcDdLcwk1lrDmCIJrnb/
L0hi2O3+6t9cWKjnUNEvWEsnUDArNuvB8b+BwPmlRTGgK6/YMM2wbs435XFwHpWU
opGxSBcOmOHLci+TrObjq3mafc3JeX77OydmKUHYjIRX0c3NaMaVQJJUYdUy5kKE
VQY1cv0M2zh7znHJTDrb5C/q7bcnTvHUqbdp00x5NKMB9Drb/4kmrnqB3SrNdN9z
y98cXMnqmnVDZTXXAUkqG3imST4uA1zlWr9oOL+ri4k05IOYFpDb8jW6SzMLAE4y
0/AYYvKtswB7808gzrJEPg+rX+SwtuqoYuKWGXkAQ9rfYVhiZq6l+aaqDzGBcVnj
Y+HXGqA46k8RA/Mx3HSM85GlduIGSUYAYMqjPjQehKezqBQGWHvO37HEeiaA7ZGh
OtJeWNhVE3049Lmrgmou4o+ABk1MZbXTal7rq4DPdhF0+QGAr1uPXU/mR/OA0Fpo
I1ROagKf+JR6qkbcaSppltiiWjyLtMXWI64XwL9SGfhrSJvj5npDjvKSuHeyIslq
lN6JmbxSVXWEVeH3PQMYqHHw4s5DnL9ZKEaAe481BfsP6MIB2DPCEB+WQsJ51zVx
g2FO9PfBawN0R+uTCODZoIWs4IHKGus+UI3FGefoECP5Secl2C2El3lhar5VUdLb
Znc4OUKan9SV5wNGd5oFYiBBuOpddEnWb+g8W6co+yBTCC+IgM+tKa8aVmxLH4DU
ajfJKoAXHSDgiHl3yD072kAaBJGyCseulseOyl/2rVQ4bxlw7WopolIAAmUv2wRd
BTypTMLUMeYUihupDPgAn2fNr50miQs6ZR8r01A9szA6mkuTR2eIkOcSOirCTl+B
Iatb6BvSHkUgLUD71zlJyh/0osEePZ4Bz54PvrkMICNCoCbFVINTKqRTaGg2AXJn
1+QpnZ/gVMgjfc+JIHMSuqUhkOE4OLmU14SO6OlvzCfEfzxy9MFJkbwYcCArcGpL
mvrkC2lBwpDbd+fVQwY6mFDBcUxH+/+ne2V5uhxpjYfOwMl6Jpwslua/xRxpjvsr
fddgHmM/DofFvz+rxHI29FvgLjUZ9raoypMNWGZjYNhm/xReysRmi9gE6/Y9/MNW
ux6s/M2EMQvLEYJtRAJz+B9NMdlH7rmvb9wfwW11AQpMZppXUkzJlsPDvrFOaMTZ
XY6Gho4NBeYa6YhDgGV+NVNSiHXr4E1LYBbVQiJtfaLpISvv/SGKRWQsF4NK8X6u
/cpWvLVkskv1brDKljma8FRTWllSXPqyQNBxoVJmduJVIicnb9bURpsxoS/lkObs
lzqE6GB1rrCK0ed1P+SOjjSc+8q2xIkaMkm7Fz2R3lgEyiSDO1l8cyk3qd0KdvKR
5qS1I32egShXp1wyjbwk7r1OqLomVs58Xbwp5Ojz1GaHa73z9EZQt/WaT4QGuKp9
ajfoysxTFsVStigTmOUXwSAjCNVzZJjsUnHs0buPecmfYyNSOZhYVe2VmimTb1SO
d/oNkcMwUJgeWVjdfz5WBlN/DM1wAZ7rvs4GJODMnNGYlN+u9yo3qBN1WWPZyW92
kFElO8HD5ym4oc9BX0urLhICj7z2j8pAkOU/DkCRp+y4kVUlKjf7yrAwrjWdpcuk
PGtSHuobjWEtF6apz85z+Krs8Lz5VF3uV9o8TkZ7W++bw1c3uxoZnt0+pFqGlAlU
XQeI21zoNSxyD83ZSUvJ05Io8TrdD0pdu+42y3mhBZcNG54oMYQIFIuC33IuHoSG
1RG+eQCTdI+ZijnqYiXAqdB4WDLqQC8gMlvxOMzM8AmY4/J2RzRmDfDQd4qxHux3
FB266xdrYzP9ynQJ2J5ngsogp63daYGPl7H93O8gRYK9OHk6mcwl2FZGiWG2GbpA
etMuJhofWBf6+WO/LxbEoHTiCFndcu3Eb35kYzf9PY13AcggGxbcnRJimeNOLJ1t
ju7/KusAclP3GyR53ry5axA3Rz+M99ODZmSGPEzofCMDdXjlvD1cAnuahYl3c9DJ
IBNcfitB0GDhjMhWZoy7VwlIGkgHF6CVr2z5pIV3JtfUCEBa7m5SCO4cY0EdOysp
ZfbCYBEFW+uhJtdAIIsU8vLQ77VWF02SeI13QEt6rnw9/6FLMRoEYIYhmP0pOUBV
/vrP37KhXQG+kxQhxEOYh/RVp8y5JmLHp0QwwUp/x4foQtZDH5VW9quo9AzduxsM
9Z0M1cZYYHaD4CyRvzP9pivsynMPQaSbBRhR99WFRNo=
`protect END_PROTECTED
