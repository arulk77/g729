`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xnOyFVGTErl0WrIZfv9PYvPsJIS7+naNpiScchE3AS+
0IaFAXqWR4cliwUqYe1yvfzyhlFHB1detfbBulPfH+Bj/oVaPjilXEU2ZePlZhsf
xGca3LiKk6Qoc1UoCjMi1PCAzJM7I/EAjpdI35ClTfNcIsDtToIQRABfIiLOId/d
xGSI6NSrDuUiTalnIAlKA/gYzZ/G5IxovgzOJYXAToVid6LAVuoOBAQ3bX6nkN18
59MSK/oYu5Z3x0cijvGRtVsodNIUvQne/NhSWAQda7ojBq3MSm4560O8/mt2NA+I
V2d6QMensklTBHED1ujMZw==
`protect END_PROTECTED
