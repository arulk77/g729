`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
iTfj0tllTHaRz/DP/vN7deXsjDDD5+UvwuNRtQowbGUw3vN7muJCRJb3dIky55po
oTz3YMjCl+A6JB4Y4k/+26BcCyoPVDGMYyRgHzpdmwDDymWzxpLBQXX89/123fVM
XW81I8tfizt0VSM6GiEnevff9CaAf85sS65Ltcyjc8f6VCytqx+RR7PSMprQTzPV
`protect END_PROTECTED
