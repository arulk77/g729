`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xrDjMgjEGEauup5I3iXrlU+U2/+790E+tqaJIXYcjpE
Rri7wzXbtAWSxtmRSTbZg6C011cGXQO/jOAd9Qu0b9Pgpb1m6o6Es0D/YIWFFD/S
c9b3uxtRJpwiUsedz2QuRhwX6wVrDFlW3HYMxYRX6bm7CP0o9N9tAqLX54BPrUh8
uRWwkGsGfYSF1s1q5X4JK6XaKH+KMZr6kEtFA7N48jeCE4/UYCS5nlEQXhuOrQtY
o2w/oB5kl2S7QuLrSp4hL+rP4rzVGkuZx33LIoUNdlE=
`protect END_PROTECTED
