`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42uXaiRaQB5CSzfUKhePamQ8ean/PI0u0K1u7IBeaHPJ
PzD6CdMNPXmP1U20GhIdV0uGTq/ocv/qbinnSBkF7jrESj+YVaVuKV2xmcJfkKJG
T/oJ9qpqcPeG58sCtHvLd1HyQALUHYl72pxScjhPRZ03MftvQnedJ091HoB+Sljb
oRVJoB3nBZIUCL1h2IOgybShKJCoX5rryVfVyh5i0kaavBDgkxC1i5723fY9mQIi
m6wzA12BD6w2H4qW/xS17pxQbkfpOaEPyhwxOCJhYxW0NCRRZUAIw7jPEVSBOPci
w+ek2HCsZj4La9YmVIGsPQ==
`protect END_PROTECTED
