`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bmw/HK7/myi/iSiani7k3kW25EBAreWm6xsLNrcWnBVJdydlQAc2C9Omeo9i7qnf
qktPQbOh5omzUmEE3cAtvhRXP4wFAjtF/GGQqp7w8lWzgPJwzR+2YDkVcUUvZ9dH
YBzVOZhW4RUEQlRL6H4SJlVMtApD4D9aFlz5aslNGRIayOel/NjTDGRclY5pvoiw
lZUykahsWa+wDyzSWR13RLN1QD17edurcjHOU/ocrCI88yn2k1PkiDXTppoou8h2
8euEqNTcc5dj7I4hky41B15qgXpUsPXvNRB9lCYG6pHxCxaBmEcJ54BLc9YSOlgk
Jwe9XJRMZdgxpQ8K6/4sHB/B7BRNus8bhWjw/nceWnI=
`protect END_PROTECTED
