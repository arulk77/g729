`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDATGKgaxRen3pNfc/6t8AdKcEv9gMesTDMZLSthKlUzvA
O2qaZyFOYie/dkW6dt00mm0fvuh1mcLftv3dOT6NT/V/01TsxExo4LGPssExALc3
XgcBMUfzwkv59hVn1iL5v7oK/2tZQHFxoN3QkfhslFqU/C4O9afupCbiJinbdmbf
nK3sabw3NaZtGwAsBvwvDWlI4yzaOTQxc9Qq2oGIMX53cZPPij5kq1mX1LDQQVx6
PRRE4LYdiVMClxr3sY51BR58arPo8dSEVHjXymHidRH8PLMcGkHiEWPr9VwFgQ7V
YQsxOS3ztBSSm1CjQHiQ5em/Q3YX6n5PnyQuEcnq6OVSOwKCjVNvSkqASTwR4Bq4
npyCuaYZDBci63lKUG/nCz/o+w63zAdE5yvZNdjXM82Hw4LAaqEcwFJWelpbgWJv
9tJSkI9jZDY6BGsq27hcAdy+zlBYADhnzVVxXqT/75fyn8eTYk3zWV1S3d3wHwUB
oL1cbqS6sKAl7WJq13sPd2X3A1dBQ8oQ/OaNuw64+4YlJ0P+mzB51os0OpurKsfb
W1uYTcSwaNsN+zhBqgyjUCieb002xVg4djiV0k5M6SmXGC8V+WneuSt2HDx1T5Il
KGdUx3vr77fr0eEPK1db2NfL5rZQgeJnUgR7Hwo73BhvMxYs7MN2gs0djvqB4BfK
3dKOCUkQkJhuE8p7IYNWsg9up9Q2tOpu0XlvLiO+Qdoq6o3b/IkqZhUQobGUoNS3
+TZsuoHWH4K82GzzML9bcjF8Zz5diFPJOxDVR2a6DN9w0M3179vKNxQ3iHAEucvf
J15rCDeViPorGzea4foYoGkcSrUsdQs+Sl49s64OeWr9MxdDwMXeFEmQpWDj620W
ggRkjaerYwYEw09hOeLCIfNB9CmIJ0J+SCbs2c/yOPdpsWyDy70CD48Q7dZ6yWcD
CvySOAuHAzqTPiZcTKtcVTBPQeKvUnDq+8rIzsCEsDMzUr1b/gM3AeJDkcRvn+f7
v65W7TKgrhs/RlRy3fvp5elX2wTUE5CblGLYmhR2FXtFNF4nGLCDj/DYoKUyCO42
X17MKyXsr5ag7pyWYAr0i/IRrygJKFQNOkoyzesmFdt7QG+sQHclZk4Nj/Z9i4RK
US1dHVZM9R/m0VQeboqbxF2QyKx4KmS2+uVZZdGtexy8VOekUZUzqcN9MRn00ykx
ZxpdlSjHBz9asXIiVj+lIZMa85prC812kzI64vtpSf5UpmAddjiIyTEXwEQGuqqJ
bkDGzAnI43oo7SgeHqynYP63m66JsSJlN0pG6yYfLWIWHpkz6VAu2zUHF+bhwH7o
f2fyanrs1z0SGGg2axzPgzojbD+GHeZuQT7B3bqNbZAQRF5n4ryF/ALIcZIuxJ6C
7Ag+eF+hr6BH+XYRMapTWX1MhvPXeqmGxPhxJEsIyWHvonvYJqJQsUdRE0ZN50JQ
pAiFJqycV93LDy+pHbwIFw5dBm/AkifcNK1w+qYNDvcdm1wIfiqgDPhOxZjGl7eP
pf5G0x7NDl6SWDEKKeblpZ/MXH4bR+e2SYO+R4xOb/f6P2dtXn5UEC3h8omfpmM1
Q9p3RQLJF3sk+Hj5XOk4oLxwjNI1MZTODT7+z5WO5ke+ezD7CqHu3n7ttLSB+Red
5Bj3kjJdROk+iOdZft2atYTbHYoYT7htr1g86WINN/iywx8Fz5JMgsw+NKW9uHPw
BxiUaWV7O2Ik/TloF5dS7sUR/+mTeqwkoJ/z/q+YSgjNuse63sODWxNjW999Rp8G
metaxid99DsnOqZe9HW+OBvWmCAWGkaiKxNvx5h8ZjHZFr811sJ8U8i+Y59QkSpt
RR/TnA3BWt86yaanAAYHD8/jPs9EVIqAqIck8DMESJkIDfzoqgjJpshfrvm9Jjka
3dKKftOPdVLcVIfSGbOcTG2ELgg45W3rghfs6aIQkXniUmTC2lo0WBL0Ge1FDkUe
ge7HHEeKtWd9q4CXFTSJhwXNBIdnq/ORGNA2mbXs9FsB1Oy73xW5I3lejIKWVIxK
Ts/dCiXZcBesVPmXxJhXmfv1odpnp8NLWgcWIEVIUqBbFSMDbOl9SIZE8+ihyBkS
aDxV0CL/SwUOXNF4Sd4iMwzoW2jkSku1qdfflcK1WG033EukiNnKIHEnHd55RwU0
E/7kRxHb8wUxlAex2383PiO1KiLLvy8/htcjGzTxlyWIA4ShVC7U0SgJm4jMQ5Ht
hngchWsRD0NDgOAal1+BsLGektB+mgYb1EBPhfpJLzyqKrUyJi46kdWTi8yq51sO
Ou955HksPEl4+zp88tT8szPIJFckefjXPe/xz3ESIXLVtMjuE18G9h74D8JGYWsH
dsg3c1AlnmlKn5ET7bSIVVKbkCKOR0qwxhw/0QhkNsOVGykw9EMFEgkFcx7h5NDU
Adx+XcXtsHE3ZIWkDb7tXvtlr3O/Ftsn7M128XimNh0OGnKP5wyr450VhTHdC7uF
/MdspSJuJb2IdQoyrIAflAEbR1A7MSNS9BKlBfsI9jksM7zNgzwkH/uml75Rmscb
8Unc5KOoA4b1+QwPvAGzEWXmI5VS98BmCIEaYEBFY6qtQ/KPmoFOtGMI48LdnoqP
5UqcMPQuvfmhMaNCdgcen6utMib8HGvdATx6QLTHRfZ4SB1j94DzLKjsNcgvyYaD
jnniBw6MQXPzt84GKNf+Ggmg4y+Y0z1RRrveFZ1ombltiMpxG0b43UMe5egXduE4
hkzdKLaElRVdSjU+bKuVMT6YTOYkQ8PyWcttGD5S8CGIsYNCuaFxmvZJzKBoVUbd
OrsXgaCENSLG9tHPl8/eluGNY59Iq9soiQPhuW5nKqWcMC4cABBouBOVXIxfeWgy
ImA4UxjkwxPHeR1jlhSD1ZfO0mD5fa6x3PHcIkT1Vev6ht+vGSTKzhmq2/8HU76V
XBP4+mdZWiPuuXBYV7SrkI/mJ/dD9p3D2iMxOb7VTutfZPED5XKN2rwHvh6W05nn
IjSEvCUjesSpbt8F1y21zA/iAf80pR7HR1Z+n7wya9BqgRah7xgn3Uy7AQbFQ83F
Tazrs3xAS6ErgjNBGTHjsEKLSixKXnTzYoeT4H4VBd09x5dKQLxuoHuKufIIQ6cD
nQAA+u8A6xpC/0L8DJyBdD6mJKzEcx0IR2uT3DAWJU5G+TiavVMKPWppuTHiCPM9
oy2J/VvuLfI/G+AvoMPkcgVdrEKQOMMAuf1b3qRgu017oDvaXn/L86P0MaeO7hyQ
adr/424d+SjXtfLY0Rh1GYm30FKfDeYFJIQJJsGdZsY9/Tvass6DsTFPshCwtBJm
qwgreSGlaKSO5CdN4xGXfHc82GF9ElbG/GsuhYYE3UxLeJjT/I9mU6YNazPenpJc
Kp5wzgR2+kp+sSOUOqRCsxfwdzugju/pLBQLGSkdcW8kJQSSRWvKZyhEuH5bx4ru
WDl1RRuJCdcMjpuPa2MYJuCCnPJsoYf7Fpl7DJAjEqppu7YFy4sj/9F9mEcf1vWg
wJPv+pWvPRziQxQO2fB+rc98jLhHMue7ssibqLh5TGpMibzHfWkumhVY9yFqt9KZ
ExDGNpaTBHvVdroScvAXuuCQPA/HYLIkYM5M9mrmX1eYfuh9OE3wB6/psio4DeR7
druJM/ZKTWUaPelPnaYOj0Mkb/E2DCq37zhF9fPR3VgklWsOIoVxeCtvJAKAWJea
vMTtK+cKUvUg4hzqn4go/ihbpAjpArXAPBtJNI8/I6iBDIg4sqH2KwIsbS1kTXr/
JDVVqSEjBBF5d3pmM24Xrd4jhagHPbUs90RUgxZ14Wk=
`protect END_PROTECTED
