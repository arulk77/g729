`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAfVqPF7QM6I7/gq1F4Fh4m7OdPkX0UteaXYVEBfLialb
gWKRStydSQDFN43gmocg2dCk3/DDjtBnCPzAK71N2bUWVJa0AaeXSMngUgBnBhPA
rd6mxBwxvHxP8KCAVY9xmEp98IRSwGxmZ7eMwEo+pZLDSq8Mmauklt5Unr8ZTKg1
xZLV2wVq4ADaQ4OcfTXA1ZMYn2iNg39+Vp9zrmO3dqgfoyVLnJleKbys1Ek1m6+B
5/pacAdggf9N3u7p3LyFk/7FWy8S1wWeyo+rXgZXfxkVl0TtoIPEyTvQqaAs2qaX
ZTf/qoWEYfyb2LaN7YDVbZPcF+Pdh+MwOB0QXfYraGZz8P/NOU9M5TOkNgyFEvAv
aQ6OoTRb4xbFdysa47jXa3gtpHOilxaEetZhpxYZljTEy6tP8ewWnmQokzgYjCjf
6cn8dWXI/OZfsm9b6hx2Pc5+o51c5zHIdlUfTMwXt60+eSnAdpcMnWbU77RtcLXT
8ovFdqNgLZajZbtDFvGcZ+4Y4yjwADf2L9bLeYvjgXZ9VsGFo3NvNE079Gaoa6HH
+tNncPJieISo31O75f3j6huFxTf1If9fOe8cUl2oiIhAoHDAiEcZdG3jM6FwhUqK
+F8d8wy2EW4yxhhV3TwIIlEdETUuJx6lH0WM2eNGTzUtWeARvmwjK/76d55NLcbV
vzAZShqUtAel5JKUoiPp0hn32op/40WiYvZW/DtNzekxvxrY2J1vXW+uVbJ2DlZG
Ij8SV9HPbmVvhRRRXttjMMqNBQpJVo05LGuQ5gC6IYkv6oFf/VaV03YBck7ytcTJ
SURmNkgh/Ola0JosmyUXit5KvZY5eSJGkEwODj38IJbqsUjkjEm/67tPYIdcGfrR
WjsxJTqIVXAcIkp0br1o5O5ag0zZ9sMW3JEckadCIrqTarGGvTrlf2gR9ehrKJZO
OYVB8Y/KZFY5uzvdNnVE//hpj/3NBy6wDQyJKMT0Gv9moXeS1ioB3ci3Som6mtHs
r/KSX9t/MPWl0WKcm7JHvFJX/Ewvo5LpU0NPFp38ME03rtvTMD3Qan1G4Z0v2tGy
UHjmqrTkLysPRZOMFBCqcDlyQfXS67GlOnfzCZ5/Remk5xGrMBls7CTb6FYInkxs
Iskl4zzpevOk/xq9P5NKdIG56bSn4eaUYqVrm8nq04ojRr4tDJtWVkoRjOlLI8Bh
3sL+vCSYPLaw1ITKLhxN4VhEPC7B8qBs0ZtAcvQQgmk6jQ0ZbR8Q1ikG338Qf/pX
C4ZyS8JRWjQZ6Wji60ciMRoXNQZUGnsFNSpsCKUQh6MyswOZjclrS6I3ZKhUQ24q
SwuwLalXuV9uhsT/bhaEjfaBCt0g9nnJNw/tntzQYUtRR56G+rxPZafO2QKeFTyV
ZWwmmI8Pd7rltaD1/PBKuLRYcLboW5aW6B10BL0EyvYFig9+ck6IiN9CpXmt8eve
zxsm1S2TqvLpIBrP9Dx3BnbKhmL2cFrFgzJyr0Q4UbqVypWei6r/GGiz97aCFBNr
9Uuvc7Gu1eKYIFzTufQ5TbjDRT5R6qB0GuXIx9uzIIxFHUNHh4AU87CFMBbd3yf4
OpI1iJ+TaN3JtUrNAJ/Xscg4fFM8Oby4oTCXm0yX+fXoVmsFU6fJ5anJkNrdrBj1
qTSW3kpnaMj9jpmC1/IHy2kxXEeTIBHSuqPC+LaH7jexrm1qh1Cg25O/ps3bzT9b
29dD3jW7Zj3Tm07w2BvbR1HhyxcFfEB/FQ9G3haQHeuTjSL+v83rKF6ZHKXnIzYY
INz7EImjEg3YlH11mR7UnlHrhX5u2S2FUf+MPlVg5vrPkVB8/fwTH8k0Ke2vWl4X
rPRjXjcB44VD7S3v9ykx/HV6mpEs8njF3reahyQIkyRDfZp+GUhN7nIWBShRXu/T
2Y8zOWAxkURorl6cpJZipzJFOZ+M9AhzJk76Ljra35IcKjSsOoQ2da7a6wnXqsy2
Zd8LEPzQf4cS20PYLerWZbvcx/5OUJVwMjkD9Ywvdxm+sj+h5Bl7wXspMSlFX+E9
+D7HBf6fgO3qBRfx/vSr9uw8yi8gQUQjJlxRc1JjY9IRQd0uKxa5CflgPmnebYjN
DYoPl/qRXvRC5nvrkqT8YL6gChJBZLj7qQYOgydXRHrCXalZPG8UujafQv2eDmEK
fVNTSstQC6TSSpTUbDRU5drdvMSQQdTq807iWamz/TUg6WGsM/VIC90QFQd053x1
6qkC/zpps4vNd93qkjOsg8Cakw8I5eqqJG7x6MRGftmKvAi9HH3rckYynG1K7NKA
N38hgOWxjoBZtopwji4HvqCa9lBTGxCDuV7rTmcD1/D4GaRFxJ2AepK9F7vboIvI
3Os6DhKZeWc5f1UItBxCZz89sqIZ3QCAY7Ub+0P25Zt/bKVqlJgrw7cffcn9Pxki
Hs57A9UPq/wZelJ7mdVT5HJ2SNgDOTvR2rzRKEeOWMp7Sg9lsNc3P8pR/N3wYnQs
j0X5RRsQmi+Nfaeinu10P5UwxW+9Vn3CSVxkjSPmLEPfh0Dtcbp6jHOIHgE/6HIX
HbywWFIj3S1+ymD1miU7K0SnjTIFKStwiNn9o2IXMMcNeuA9lF8129PN18qa/Hyx
g7sDoUKmq6sKgfGMHQRp/3M3X6JKfWkJ7YHqYFNhXl/pRMZXxGp7k54KzoZ0cPP6
mCLUpMze+NXCItJJzwESmDIkXekKPGzwtBKzvpqphVeg6p+QIxW/4m9ZCdx2zdda
DTgc1GbUaRl2rL0oyhtskyU7D57XSpWxgb4KnK6ITj7zzA/0hbTFATkCzZ7VX/cO
t1OWFuA+j0cI7qxCTc/cgki1UTgjbT/6glPP6x3sZ1ijYzzzcLGZe8bQRPlaq8wu
+ZEAX9yP1omndFp3LqLRUbBYipuBwJUwrdIp0w1Yq5h6OoS2U7SPVSsZmbWBRnKD
9GnlKznculSmhrMQ1jDUxRTOjLUz+zJk3ivAEl79ksg5P19m6MMmYR4KKIOrBnzB
xbLYGRbDHQkMvWVg/3qOyqtSJSCyvwp8BzRO6YAMpUl5R1TqI3KPHTRLq/YoVKh1
bEoeptHvqKGbfn9IEmABq43mNxgrukIT5geVwG9YTuCtxUaAEyRkP+DU5Ol4+Xcd
hISJvCC/rwHXh93fPiT5PjJ8B6VotbU0o3MFFyGzMyo=
`protect END_PROTECTED
