`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4976YijzeplrG1JgF6SuKSvJTqIaKihyrsoUMLXJvqpR
0Ab97Mn12k4LgBqfzHDnTnEIGgyuaUujAnkXLbifq69QfyIrzl7c4iP52QhuvE3U
jtmGb3STDWzqzhviuLTBY5PwMuVOyJdrO2yGakustKy1pqCv98+IAoFKdfv3CuW9
poMAVrP0XXyJ85esZVoxFgJVcFoEUCNCEYiMTs9qgwQ=
`protect END_PROTECTED
