`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
iHHao+oqNy2mWM12RDxAG9+XGu7+Z7OEUUemESfIwGl2D/H9THg6M6ipZLDSyh+w
DeWQkLRkFAfem1kLVnbztcdh65pojDMabgZqiOrqHXAeZRb6ohupA8CtMLYvPM4D
dntkSqAmScdms2+6zjU52uJO4xhKYbeor1AkWg7/WBozboK47xwGaK1nGeIbodVG
F9ulZdaJNxKu+U0nq5omiwvIn4Xe3hyWDB/ilzs4kdqkEPhC0XFJW7GbmILA9pEk
8UDgVgmenl7rTgBVtlQCjbgtMJHvRFXexetEm9j1psiQfeLAGDj0P/RvP/aJjXRr
SZxzJzHiDdmkr7OguKvpak9loe00MaspTWz7FguqVFlZChz/CrbtvUirT0Yfy8DY
OUco85hEsesqjMHOL7AauhBXtR+YTFw21QR6gvlpSaO35n5I5avRIh1fINpOFIB5
Si1kLSSxy0NT3qR8NQIC2r2VNPIuLr33zbMlBH6S6udY8WpgFaGuSb7yFX+gPNJm
oMHUeZvTFYCLZ3wV94naKUhsIXwzCHX+ITYd2kOZdROlSfwg56LSqM9P9GbR42xI
hGDw86dPX/+U+CPQkKG5USTUX2l8Y3i4WwQePCxpDET0fEbg1KfGAeRECQqs3gms
7CuRsqxuJlowuwvYXFHvOl5/FXd4XCXnVQwNKE1Vqot6NQCeYU2nIaBuO7l3xHeT
f8uKbZSLXtnsU23Sjl3xX1LlA3SQQOScC7gQyWCyt9Q=
`protect END_PROTECTED
