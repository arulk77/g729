`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
fwMWyer3i6QJ10swv2+Sb6aavKh5c7hMCbQmlNGAli/n9PAnt2HGBAc9hijeVDBk
0ITJi/5GK7b3rsUUntK+uzxcLGHaYObgYo4rlKvViauRh0xb3AucB3lvco+2EiJl
ZyaP2i8AcOVgrwQ14nLJ3wMeNpUY6uRLsCc90TcNpheprlXYQZnJGC51LaTZYVS+
1X5932+wbc+hd8fxZ9opvNWWX3xfjrfrPhCj59nqz6+Zkb6BKei86QGVPMI1VNHn
yuvKHhRlrhb7al/bhwJZqheHp9q1l8G+foKmmHri2aKikgWkellwXSA7Fl7BBnS0
sL3afa4d7+IRuXMT4PCAseaA+z4WNCkwL8iTOaQe+vef+OkDbwruDK4jbJVVq4Lx
0hSWwX6vWUaa2fmYoW+nNA==
`protect END_PROTECTED
