`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
f9hoN5aXPTJcXZFa+HDOYCDqGmdXVBs/9z+ve/WChRKJKzx2X/JqAHSNA8kAxrR3
vJ27vK3cHe/QdhbwLDaGDexMaw3b+IH8FPFGZBgMQsbeKmTw6PtPaIbjLR7ArLvx
UhrOMs0IcAGJzKi+v3fVF/GoY60rbOfZjTHDa6FvOTLLGuDw4b8hdXlS9OMoJeH+
UdHuVtV0bSvwwUcUHb6EqHXJeqDnGoxB0iHhEqb2YZNP8HfSq3jrReZuUa7cq6nY
QUbrotGoeR3XdhHwc/9rHEF/9AL8MeGHQ4pCXXeHSlcOGQkIx3ewuTHxDhOozyqr
i67bG7IL36+hGeeQ9BIkdl3faDSyN267Jxx1hRzRNi4SsdLVGCi+hVXlyYRAoGWC
KOAvPkl5ThIwkYv4HJIAAChjQb0PwG31WEGN3Z5Z5td67hUM57qd7bUYPZrkqYSn
QCp41V+mNFQurekZ7jApQIEhHeDXA+gO3QxduBoKg8ksGwaFART+c2KBZwhyy2w+
HI5L+mapkFT+b1WtISyywKl0gX20rlAMF/E7poWuQB1qBfUIB9B/fkCaAauKwcUD
0WtW/egfuKlcMx3WOAUlWrmI0fkcfiiduJ3/0sHL84oVUxZ4X4B+K537U1IupI6E
78l27AdZx0DAtbzbuJcCpRqHJ6vITU5HZlLEmK+0H33iWvLi2MK+csfb90n/eDJS
m6o162vi+Tp8tp9SA7ApCAxbRNBMasiPEwnJGfAZIbMFm4IcxCAW8sbBSESXpKXv
ttxjLOLVeDefSFnZKZ4kK0M8ONJZio5dYb+WKUujhRK3cxeJyfWRgzjGxC6TSdSe
IxW12WtaeQ5LOFf5wbm52PyLx+SdkupP7DwME6fb9HOq5BLz8IKoyCUOF+9PrFFp
Ki2IfPtwRaaTRlAVtvW1T8VtITbCMsmWxZkCtTvOewjZeUFLaBdor3ei2Vv5AogH
61a9WQr4SobKDUaq46tjuOUSQp9l6O8VJ1SNt0O7Wpn3ToW8bqol4vm8p/Gcqn/c
`protect END_PROTECTED
