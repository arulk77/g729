`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKMam8jO3dn2LQmE+8CKu0tvbfnT0vVG0MyNNfytV8sx
D3aB1Fdl1LrJNiBS85tRTcpU01BMMsGHywPQVgLuhjOsSRpJQbx8SzupF/U6HI9C
HLeDI2PJfMUtm7lKWwRgKxa9hUI72Xd0255nNosQuorQ7CtzZuswyxISxhSWVkYr
nsJJHXi2WXwPLEEK2UkaKe591W3zlftmcczi187Wv2xu1yUVL3KDvc37+B37XNm/
WK9fRww7axZq9d1dLiFWg+wY0P/3ckGtcUK36bwYWm5SE6yJ3HJG+yWi5rz8toPq
Vjm59AJ4pUcQGIZD4dVIAvzRIDea2DA3asEC8fmHy8KneteXML4Z9zFLHhCMPeDi
blB1JM5RlLY3rtNKbTtGbJW2TIUPIdhaF7zzAzUfcFBwvfxd+IshprHNbSbF8Zqo
`protect END_PROTECTED
