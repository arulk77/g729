`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveERAEzdAu1AGJeNvOhrNyJ7bxq9HVHwpCnBsvyC2rHgO
O12dgEmu68vyg9VjW3Zk5iGmvTUYX+dwL024UjSCjWBBQ3PkEoKA5SHFgc52bYsS
bNsERQXwNCnrsTf3spI3Y22BD38Pnk+9SAyE4pZyk/QUnHaZ3OF/gkgyqln5KVRb
2D4s+gKhQZrFy35a/2ONtY/KhLirbk0UtmXB+9s5OJ9visNqRYgZ4SBypBLrQxjm
tciMiZNKNyYeTt0svwXkgrHJ9j7qENelobKzWBvpgQaZEe4Ywl92DAAstycit45j
/sXfyAwd7CrnkSlk+tB1TA==
`protect END_PROTECTED
