`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
72DKe5MEZSH9IT4s+0rFcFee5YB0HhWIITrbQuATsLHB+k5YUFwqXccTEp8sQB3X
YeZkQHH3qPjcxt2812uh/gU93oAlH2BkY/UVryD9EJLptqr8xxUREMeyHsh2k7eN
HNnnGT7Ub1fZFtEWDocvkQHmPGWjh3Jc+PiEfmdQDKCZmuuyhLJAa2RzhUmhYL6p
R0U/hA8SitS2r0o6lkJqfcGmDxvsrueeCe1oT7YxbXPDl1rNVZJOdlw0IFQrM7SH
06OeBNsYepmsFc7zv1GfxG1xw2z+8sX0KAKCJ2dkiMAtExIgao13J+5VvpB6Y3ue
`protect END_PROTECTED
