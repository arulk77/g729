`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
CB3A4srEmGXY9Ppj7DRSTNEbfUAEqG2LDqR3l+fRWSdTX4alkPG4tmKHoo2rN2sh
+bgJWR80BMn0ocMLobvglMl2UkaXaIW7zJzZjuixWRvdCDsJLf1uQ6tfmaaDdJ/x
WgZsdCuf94AAg12dDHXMrZQx1Hs3OddLbkCdfacrTTXl6/eoJMHiEm7cIy3n80rS
nZMUdgK1Hv07C78ac/GDcO77AqTqVHEPGE7nzhk+SBmIxbnCmd5+LNNJfibJ/Ja6
KXXPsXda37Uk8zgBvKiuWJT2ngo4OTZjCFL1l/x5Cmg=
`protect END_PROTECTED
