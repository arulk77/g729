`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aVxZwYhzmnxsIjvatSa2HZfGUBtMVzjsfHvrnbWxH77i
06lOriCbqKVlV+lTJTIg+6/3xRdVXHljuRoW605mwyc7BooKRomeBcPsFQi5ZI7h
xMIt5UjGNdPsX29XQrsMbcwq+GNslma2gN6nbfAG/eKXBpZNdNbHwl1bcJBbYL6f
XgS0mGQ6i09qQjVRPqnVqXJf0MBhIn2D10HHegXgyv5ARBjnXU9DDBujG1ivHOYH
44mh75uKwMxkG+V+09jGtMGNacRPyp61Zf2n1SpTqIN7eaEt+wHHW3m07ReeKA/O
ipKh3XLJ1fb7CwtaMOT35LUXXxGUvrxHOa7eX3Tw8U5rU3bB4qh6siJURR8+qJAO
fu+r7jyoCrBJP2udKmQfxgS/GGYOZBjyqQ7yFw26z8M5EICFpZcxR+uezl//4RbZ
JZlvjlr/sob1rK4XdZK6zh3T4d8E8aGRopRI3q+FYZLD6yc9IZe9WJDxc+CqXxEI
yKujrD04QFKushbAOySw6klvhkTKD+PxXWNE2hTfIrd5oxKzLkvCVWONv+Ruxh7r
JtoF72/y9ismEoTKtplRXO3On2BthOW7uR3bMbsMa2ZdeCXmZ5Z8BhuvBrbvUyz2
AUJu2gSntyxC55o/LqMtqbz/h/3MkEXSpNtlamxIcBFgwozK0cm0OdwAF3P1Sq2k
SBOYNw48Gy/orLoqoIZPOaWVeCbC9fx3nHGM0rK4IwioC2V8g3CWsV9vplRgrOpO
AayieEh3VxUJSGrOarG6Rsx1oadonrE046yLAJhukkPocjbqfoi3PjhnP6Ah/jsa
wykKRtO1vHuV/8O/7d9DuUOdH7jfMAU2hPVl/O/75s57GM5A+910FGGJf4GAXtpI
lq1cpG5IpEB9WNrxEBFKG5SAdzKwkYJlBo5WVmqfSWlfl4zKz1FkKdfhhyKEOiwS
2b7ML9hrYbAd3eGRa1D+LeoajPBwP15B+FL+11F+a2s5eatJSA0KWGPG/QxGrAA9
a2RBwK2UEyff5nQw/QgCF8n8kh1owGMFmJE5e4fjXP5M8sOtX6OOk55QJULx3XHu
EBXwW9bxwn7qh7dXtDipMg==
`protect END_PROTECTED
