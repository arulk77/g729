`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
W42gJPalbz2Q2N/rbLtGCrFJuZBl+RX/8Y6uRvbs6/0KZY5Y6vKH/7ABu07YNO3b
QslNbNmCpgIljkDW2phkaxfQS0zP70PNpdRSqR/Fxkmi8wm1+LmOcDd4iJD94RRy
BQwrJosQcsotnS5BkRQajOXozRAEF8E7ASaAP4sAYDYnh5ztyP83dn5/wlFE4N7i
8QpIJH5HTQpquo/19ESALTB020jmHvFtDfYoV58JhSQ=
`protect END_PROTECTED
