`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDq8BLoFEburJ+JttnLjagC/RwCMfwxxoMxGCetgTDnN
4oaqNhPSzfNwGlOEB6MapmQGttWTvhFftDj7hhAiAxRu8tg+4cnP5CFJ7bQBVqjV
KMIeDBJUN1noP6cdRp4NtqhWg/SJxIe2hjP6XoVjDxJODKXAGK+651j5uEsMznHD
6kJQeg+kI1dkVXgeDu2ygJU3pU+qh6bWBTH422BbUe4xgRxUL8nS85UeLqTQkgNp
`protect END_PROTECTED
