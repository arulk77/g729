`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP0TSKeR/e5OOXEFJRjDx7pIIx1GkJyKeXfeBWhsbTyP
Se8i7osvBeo8rLjfQ02gAgFpRzz2c38PfKbe2K9KMj9LVCM8n6ibSUxgrcHcPf3r
aOSY4973QRRkzeepS2MCqiy2vahE3E2KorEhYgPYU90kr5gYysFXpr6M5kFMHL7E
BOGKTPfJsM8PtPvBf8qWAy2HOsoqY2MbAPT7GwEyrY3WLcQse13OKx5xqoTkvYaQ
bP6OlzhjfZbv/fv4ErJw3HD7xmP0NPEUhJpKEJPuL8e5XOYPVFLSDcBKA0rXmCm5
xs+/QzPhJqjLIdweKO2EHQ==
`protect END_PROTECTED
