`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCLdtTg/QHoYQP4dMpnAXM53DKPEuViqUVVK1jJVxpj1
2z/DWWhi8LOP9TOc77A5GUfIc1UWJDl6Lbu5+OHXwaY3w2uhGCCjXIgLCS6zM+mH
SfxTYSwIMCumRlDRqmC9J3FKnu6ZuYKG3Mv+0wUKN96oWHBnLw8NFnlw70VVsJJY
L5N/rTc86vWI0pLr6Ldf6LQsZIUt/k54xlrFOq2uIfxu5/NhTvNAl5A5NhJIaJMd
ph9pmmDRphfiA4z74MSw3O4/WHtDOw2eiFFhRcdgbOjxkNYlz9slGD9wkmfCFBk0
9UfcsSj6CpjPfihJct+yIDcrsNCjgF40rdn7k7nOTEpv3J9uRuCL7SsfCO5FFgS0
7MTMeEFkXeiBT2REzbTU+A==
`protect END_PROTECTED
