`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44vrPORFQjQQa8O0EAfrE9+1Ch+TTp41GaIv6mhywcZv
xXs9WTqAutONgIdyB4yuz0txWARe6nxSsHE1xV0YS2Vs7O9mHdMEJnVFnPfVaMEA
E26tfpkVDa5xZ1r6ImC0oFmcSzoMsqh5xaY4E5xCx2q0TJQ8kEyofpYFS12Qby+b
EBdNLRRcz+TybGf6zyHl3joYhX+KFedGl9Z8dWfunO3odo2r6MeTLFC7AkLjREXV
BGNcpCrlgeuYm1iMY5L5Q3A6E67coU2/ITC9l+DJSz/rISUHJR+qVZErrZOAcpcK
9/LJQDrn1QW9p3zALJjn5z4GrcnHrSeDYc1ZJn6j+52A26gCfo+OkiUC1aMDwpS8
nOufMw4XoAekG7kS/bkDtw==
`protect END_PROTECTED
