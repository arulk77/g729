`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIgeUD+XGTIM7Rs34xW2dv7UStvRZIl33mCnYCc5qs0O
eBKYPDZjZgMmeJUi06eamNRcLT+xYubCDxaBFmoxHPDvXsOHj/oDsIfd1UdAewR/
XcKE4o/22ut6eFwS7lqxvQ3Rwtyaq5VMYn2cZaPRWAhSG8yISi2T+djrV6mxWwKS
udu9oY+EJacaPgJbYECZrM2yqI8/w7nufPGvPFh8Ph+dKPGibXW7XBh5EyPGvaku
sr2ft82RFbxnokUWYvp0kxIkFrOB9YjiTRzpE2KTk3JpOyfEXG+y9yt4bJOtzwr+
ztZrnFptoA6D+egLKiF3EA==
`protect END_PROTECTED
