`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1acSMhP3J0+VUsjOASvYSaa6T2yf+lguJn9mOcDQDQOZC
JbaHqgCXfD7uX9MIsK1TuwmRubyUoOtbR+T8bbXIxVhf5w+DyRhXnI6az+OxlVcN
Fu0GmUoHfKWcsZATdBjnRuhUIC+4yvg+1UDUVTEv9v7PUk4LpoSIpc9YGG6XWY3c
oqNzJ8QEo9va/OPprvxcQVEKBrdCxJKKcZOOwaHRqvbKhfuOZh4mNt32yi9ShsJt
xf24CViWiIOH7VkZohLuQH9Amimc2Gs0igm4kGmCl6JKCt2L8jEovcLeYvL3FT/c
fl2+qkJFLpQClaosNUKTM1UWfS5oI0GkbPWhoiez7qckRno+br7rYh6LAmYXoSFT
3dwrLGg155rhJzK+0W0wyy0jW8dUyUHP7PXBF1/hEqJTPS+kudTDje817V3PJl86
CHvF7EWS2o+iHDgOkrenGpqPpi/T56QKMv2orU+rsqgp65TGqhviUU21pfZBBp2c
22tH91PgcrK4rXlFVheQEbPiACXdr47pSTsAPf+6U8R7/y3t79HrvsDgIp32D9mn
zQKU9W9eO3Bvw/Wob2qBw+hV+IqMXjmFYYsHl0js8xBgKmlKVQL25AbUY6w6aiRa
kXVEBzWTDjI+tlbIetB/1RtqfWbO7dmSDemb/nstLu/w2iuLEkpn0nah40WWcKf1
7Ltpd4QOddDFvcOX6hWkq+NPpA8l3HK0UGTv7+2Dxp0bUsiV14NjTLiXlm1iNABV
PzQOliTtzgtvNjxf0hWZVpeOob4knpNXX2nq9btaGzZaGuLYZ2tAalLSrNiLzicw
R9Sb9fMR+jfnN0yW9odQJD50nrPAongVsbMZXoaMq78R4Ui2/Wsr+yCFY5oHQ3OQ
dBbXkCyDJtrPkDKBc1laVoM1fatX3HfkedV8z1lj5Y+cmMyLGu/tJCoig2unZvrJ
9oNOK6arkcfxr9bRCakRClmDrxlzoKcceLcYpKwlV0wSphTwYAJVGM55wkJlDjvC
F8+bG3tl6WAWQMbcPfTm1dfaQAL2nuUNkBS5LFchl40QWpMqlJfOaVNd8dr3uqVx
v8E4/byfNCm5GpWZ1k2eNElYPFhbV47KqQolhtyX3m5JRdziwnR/mG/GZJavmKgW
mBZ+DXm79RHRoqa5wsT4dIyGOLhRX1kphbHp3VI3cj/UOaL13xdnZ8bWvE0aQUy3
oODNDgIUbjGrz8CFnOdUV2Dr4JIO7qNtEavvomQzls259TQdNxJGTGdLDcorsUmT
PwaMqlDSUojmcC4J69e2fIBb68CD9bm9tJKgoHhmwVObLTjvP6qIWLa6gXYOLGVG
xbmz8z+JpK73vFb4xqq9m0qHNk7bGPa/TDgTFKxCazAYNf/r0aULO9iy3VSN5YGN
KdthXiF2AwFaZdL/7P4v7rw+BTD1292Y4RgVTpx5UPMAdhUMqAzRjJp8Q6w7orKD
ozxQfgAIwu7GMVoeJlcu+B1EBjDneCQwvG3lFkW2NUTJgNSWW2yUxx8qrtEJ5wOS
ZTpiowAqUwWSwbRrOb5cLT0bpNjnnbXMsfqEGW9HcgRWZME4lIaMadQyymPdn0bS
+qbyFK5l1Ynva27X7XzCNCqVfovNCdxmfpMypRzVfz6axR20RcLu1zSSYXAaCvNH
oCwnUePD162MiXInYKtxje9vMz/SrgOjvA25HYmeR3iN94U6A2b1uUtEOwV3MKgv
zWbzuW0ukdWRoG+iQal8H+QulF0SwK6vT4cWYqV/uRrz20f4ci+CCZbHDrFt+PV2
suQVXrpwvE/yURgadIXmw8yMVE0zlAxAuCLpsbrp+s5UScVkHB75bXx1iMu/30YH
0Ccs6ZODve6JHsS5sek20w==
`protect END_PROTECTED
