`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aa+RyurEPpXoFhHq9eM4nGB7dLmCt90g6O4WNnD6XVeb
mg9uWzr8ZBRBYH6fbOiZ/8+QmUjupXf05dSW8aA450gQRCv00A7yvpZvIMsh9W2d
oOf1ERngdsZmm+r4h+Dun7/iyzW40Wg5YUxF9155f6w+Qw8HRQ99SMpLGopEl43G
k8fKd2IsNHLen7VOFPDjFgeLpZlwZmCzqCYXV0vGBOymQk3AVmHZuAeGIKB4w1J1
NLAgxuOZgM65zqp561TWzyRu7VXRHeyzmLkePPnW8ZuFjIC1Xu51sZgdCn7SQ0ne
6wNLW3RcD0FST/xCVjy3EP6VS8PEftsUju5fWu7C47eM3yRjZY9GjYpkbZXNK3P2
0P77Aq1z0658N2vq87hKzX48SVEcs5kB0HVmlqR5CarKejLUsugplZVLCmrQCX9W
ZRwTwlNOb+bW1rQ72GMex6VVF7pQiMAVHdTn2TNsTeSzSh/rsXbYW1ZN6LGWT1St
BboMVt9dxf7bLAyIZn+J3u0/RteHoBvuz6KQf/0G+cOCrOx/42oegxsuYFA++f7Z
0zOMOPqE/dnGU/G3R9kNL4eS3twgrqYFYCfFZts21lY39eJUfRDLuSDAR14ap8MA
ZeYGnE3rl+m/Tc8KQQVpQ20bxJOcQLmtfjqlcy5TXs6xa6LLB/G9WEvLFdOkFg+9
VcfPe0IIF3nLv/z64PyT3P9/3gThMjHjdN8UMgDMYvmgEsV+st8+nhPGxPjbZj7o
zESe21D0UFJhfmNp0AiE+bsfTd3ABfOezWaTO1nmxlEEcuxbpbrOlQRQqvHZ1/hr
3j+nAuGiR26Ga9IrUoa5fZEJjRuF2RfFodpzQw5ipOCW+BjxdpGmQ7/JQrz+2AH7
fodcEvw4lmTwVwQH3JPlS9aUsXTabLhLGvJt6HlXtSYnq8VQeEeIOU3VKnXTkwRS
iro1nvroRtqvCOAHZJS7IXCBVFR5P21utiDM+TX/IRVXRL0KiJFH00ODJYyeAcW6
O9ce5eJQpKrxS5UpVKp4b1pvriSsUiuAU+9TnbErnsuv8jiBDdOHp51PQjurOEZW
ljO030B7M54XRzMckA/+kX40exmgGMF648hlF7uzeqgVcMdv7ATdhv1awG08NCUh
Szf3LQ/U0hZPOXWc8aPoW4yToTgXjv/iurWpVgI3Nwy6IWCGp4FnPjcMoVv5zkHH
YlFtRX8lGBn1WN5idHzheqg8ziGUXD63hOE8lF4XlmrtbBEVCcDysGlsqZLKCmcg
FdE27R9x0t/CgbBXiBikPW1Z1yeADxWB2d5OeeOYHKXvH2n494TGIGRSFsf5js7P
sle5K731+BpNaWlukexlfEMZ52LHLRc+m8N5KrnRZEhf2+URsVm/D3z8QvQTw5dc
JvpWdC9Jk+vm2p6+f16sh7CEj1pyan8FuYJFX5/jddZwaQLprGoxkBj6eZFb2w1c
skhS3CEJF5pu9jn24Cp54v5ia2xsXTtT1g/Yh+gKFCMV+8j6EID4P1wKi+z3GjsL
2Wg1y3HbNPUKoaojho+66TWZHq5MEKePhhbkaK6rw/6cE1goE7ps0BTsml9+IDyy
UJZSoEfQe0/b4BnwwqPTnNJMvLw+L3aHdjB8riYBxbyVYTllE4g2jtBU2WwWTE9x
+tXHxj3tSGymWLh6CmwNvmEGqg5Tk2w5YhaPyO7+7MkxWbibvVABVvhu8CVRaqfk
IwFzt7akgZk5vDKOcn9ZVEP4KhmsuaMtJMN3xdAtf174df1cfrsknMjeAhuwzQML
gretZd8E+cet1Dgme2mIUic29dLZb4bxVCxklpvnI9jBPg4M3m6UmKwnbVPBv81h
5BcZr/i2vBATwBJT4w5japBa+rTmi76Qg3xo0C6zQ4eYz7VCmxhfa6bs5MZl1PkR
aZuUDQAYtBNQ1MffR6Fu4OQpg9+SwDbMxEp4F7wcA4pmdN8GCjgV4ooQ75TE5yRL
02Arw1smo/ssofIgVGxNqQUSpfVzulBpxDhVmSHnRWP2hjP5goqoozvYCgMI2SGr
JV5rkMx6DverW2S9+53IGVzJjDN6+Tg4CASeiT7hgyqonu4FgoZhWivrKNuNR1JV
n/gCJfyBJU7S1aEBtW9YyIr0k3Dym46RaxBQ0EnyPc6FQOcjO4nYhkVXs7+OdMbf
+kz7GTdR2z1cNxPE3GPao4lYJgN70jCIawpeAirkretGOJPgCxZa64X/99DbHz1p
OVnQ+Vf/GZT05zUn3BX2wrZZNyqgwiSHEg3BJiVzcUGByUw8Dy6t0PAMIokuu4IZ
cfogA0ruxPePHc8TFXibeZEcvjfeLNzewYiMuTm/TPhz4OI+s4rUE9YVhAlB6amp
srTSeNGYuLjTdtIikS+BMTNEtE7Hno2iE0+KM+ER7KByTkIYcszaLZ0WexM00pdq
taiqKbbKv8jZnuS/8no9RM7C5TYUGN2mJI3nl7ORJI1Gn9MWCt+1DZ+DR5oWRX8j
QY/oiP344lWeHwV1qWwRNic5OPGv28Vma0W2+NncRGxSxlBTY3854FBmH5idbPhj
KeDOjNiQZwJEhBUQZP/dRe8hwc+avgiirWdwqee/GA1t5ibLAzohZL1A3iP5kgu1
R3xLl3OVjge/bN0VTRWBpiunxh8ugRvCLOZhup/67dyGMCsT5tnrLRpZovqOgnzg
QLBoEavl9kFvuJPLyP30ltgBPL+3mx0TVyaIejg5T8fGr+zpdH1FP/vObsTHBXtt
zH4WjXIyUpZnZ8q7R7GKo4T7pwvbyY0vUxzY7E3l3VIEnTJdaiBjDsZWl4dcdWwN
7QrdX7vnxm5AzbhqhbDnpRPNTAwU+7zbOjJbOGGm2mnsiz6ciUqVYbaSrLdiSTjo
irtqIOSO1SmcDzLNe9zIuxhT6+yt1B6arFof5uS5WUVGduLa1TqPESIUF/Go+Las
Ini5EZnqCJC6gUja6grPoKCuYCsmJA/KJFL01NaCKc5KiWu4rUxEJVvMmeXKwMlh
hX+SE10pqhYBcCE31HJJvXFGBpW0vz3vZWh2hmTCq82rvQobXWMgNGkQ0dIynoWr
BgfuW8DZnvQJey2qOBWgffTK9euybnphByZMCAGABmE0EFFnUlhsCY4L4X6lGfCy
57ZdPYlhZRS8OBQWUV3jfJTKfLkJJvcZLn1LYdhrwGBJqz/PmAwZRzn2sx6XZxw6
Cr1F9f4+BUMIolIv4/9aJHjmuDvpeohA9yO3dpCqdtvehVuULLZd3Z4Xezl22+17
VIUWS4ekFzSb/r/dEuT16XMY3tXdsUSiKewhs7CMw1UDf04WQ6DXSkMpV8RAyyO7
eYE+kVEJQrkVZeRIKlhguF6HlgTsbNkCYmKl67FHBjpT/SUefEyV9/VMxx8gGJ/h
TYeGBRjtvRi/i6YEYttZHZbjBnySBhcm1v1It9IIYXmodjVNg2BLFVRaED1+W0Uv
pXw/hkE16OZNc6MuY42P2u+MYt4VJI4KamIeZGA+Gh0RjcMOzDUMIi+qt0ZKYWgW
M5SKN4ZLKE8X2FHfbmfBtK92ne//M17mLa+xtS80DY/Peb0UrO60fhfMPzalQaIB
Sdy1fIRuLRGyRI6QTfJ1csiscXS8Y10wfmjlUivlUl/u8bAgNLX7UEhBGiVKK7aQ
e2DunnzKPFiEuAfQsE9BJ501UVlKaOa+v7ZlnlnoYC3Gol8OcmHgE4YrQoc/VKae
qavSTZ3qZGTVlHVmELaYpclFmsz5eAvaONG1XPhiXajQ+nDh+vnXaGN2lucKhtfi
RkBZ8lCSmtOt0fcc9WvcpzgjA5vytSGlXbMxDTsK7u4Qsgq8mg7SXFp4BqIJO06a
PQo2muFIKsCaPzJl+YSVdmzHQUh16VUlj1Acb/WWpaK4HLYz9Mn4eQ633BDiYII5
1Vw8DcyfsA1S6xJE07RwIMpXZoj0Hq1peqWyWHh8WFLtdMjeTcK60REDMpa5GRCJ
0SloxpRdzX0EuqjsbuM6xAUMq0zEEJGrT1oZ2wV7XE6XIlABLzF7ZYY6e8Xe05oA
4qMPK4fXv+wDSs1POaBH0REuVYbHtkkkERWY85XLhWDTbwIlcRkFWJ0xRsu2h+AO
+QNPCprK3P0bBwSzLCHlzj3QEuUWQaFipWW+vUVIe0WepSc19mIZg3b7gAojtAHN
97miGh5KI2v4IsWV9Nyim0nodFKNoP2H2BFIo5GQFkCmIFVYDeswWyGQOEnprgZg
0B74Ez9X03gRPv3h7IucSkdl8YJW5tRXnwed/7w2se1pTGcKfz4/9RGiwB9QTIQY
Es897B9sQbpZfOrYMzAMuVW7+fmlUPl1qmjNEoXNfF+2usrb9upOtxXEO4jw167B
ttTG1QCdH7w1RXcJCzUg+fLBMREsiRO+Iq4L6LzI4QqT12YZGZ5mNJHMeLx4uK0X
YSyOxuuD5Ip6mrErd1nUl6z07oymLeGh8hffAbXCX67FziIgQTx/N4lbYS/6FIUR
tmwY282s3+48bCY+KNNX82mfU1eE0IUZtSz8l3pJuk5b5+LZQ1yWEdQ6eFOKaf4I
kuNM+LvS3tG8b/g3CVKDNtznesm0h5Z+T1bU9YYzcxBVCzc9YwW6QzZ1LUdkqWJX
rkSamFlm4YmEYe/gOKF46sV2WRpUlW6Sz5RMn+R1TfvnvHjMIGPM++fLsPxwqUt3
lJafaEuqEKXCAJqZQUZOoOmW90/r4Xf9iaOd82lADEFlQJqBkZjpe0A1Lntl2wjF
IbOJcw9apWkbNXd0251Ff9iwj0WkHJdVZjemxu6bB//eLhXzkuC/7ggDPtAwsuH6
soqW2OOWqlyRG22Ci/cKaV5M90JwuwsiTPCRYx+SloBmPkez2PK9etDlR44jsHrn
l7pjtcEX19/lR8ZRuLBuS38AgM2obmmKpsVZt5OvKbZvtFnUAgM/kCin2a86Wf5d
fBa2qRn9NSO87aGRGKeji3gQXktOwRc1iRxdq/XN34WZch5hkwkOD3CNwLd1av3h
k1oEJEhDMD01onlSMW6jyNFuhGLuEr+B/eyoRkpH2xLc5a7TgjSR7YWp8rl+nXCa
9s1KG3F5PtmFKXAvm6qxMGc0V/CSEGC0N75J7XdMneQq/zimK54Yi7kj7bLI3A3T
a/M7Bf0iKGXrYy9t7du4e+zy4Fepidhlt0LUzyDBhFZBtm1nbbtIzgXi+7czF6bB
5E0GgrY5ziP1DpTbNvLM4QT7FMCRhCMjESjBTwFdVK2S3NkdZTysgKWQZj0WUivh
k6Ne7IqoBYPIZCvZrjp33XtXcsL3D6WLkG1f97XYHtTshlFSddGbCLrfpynyDAOt
bk+ms8aUkUm9qQh9tmwRap/9rVl7T4uoRUUJntXU8GLZk1OOHXMWbNrxGqwplF4X
8qYlWReEiLGx5ocS+C4mY1r/eCbwh/AropnWeHoJKLl2dqXfVfkt0Qeih5++cBOY
eoWJRNLv7vdwhURXvrRQSC+yGygAxFnLkB57QV5nZzAOTT7+aEKCHt6MiyIBQSGC
WSOKDoZysEHjAAY8eMSr7xsIGM4bBqrTy41kUGczu+2kUvNYbWcKSZG1TFblN8Ma
d/r0AOjUE0spu/YiQ8sefFra60DCzC5K0w6wkNN9F4l46qQvlR6qCW6on9UgwqhX
ZSQoPVphhVxgZRlno6xkpKlQe+ZiM5zHZ0bBKkoU254qgUxVnI5Dyb3gSt22Bdn2
Uv51Avuhbf1ptI+oJjfqJqo4DCpLrCN95MpNDlFhswkXpOgDdzgejNP/I+4GSkw2
NRUaX0y5/fzEXSI23J5YaH6KdmkNk1xK+1QJWv8ifu9bA4eabXpOtjzlL5SGwNdn
q5wk0BJTyDeL47T+R2jQLvfUUrxx6cSC03YgYa1g5qOzG7cVWlndBRdXbFt9d49m
z96ehCqHdIa1+hHzRC4yRR1b1iXB/7d82ZnT95dWgieLMmTXsAds92sDDpuefbaH
htU2WHUDfoqXE+qy13xrzXy9JC5WoaKzWaNTd4Yn+chLdHRHuPBV0H6UDaSzUgJF
QRhP0ZNQ8a9VgpWMJCKzoquL2BIYEAxPr6heQSdF9owMMIa9W0hFjDxnv+cMYnTD
e3NS12tvzws1h4gUaYk9NKgtxiUx5eN91kiD3UrOuzC9nR0qXKuZ1qdt0dY00B/0
cc0a/zc/mXbgAus//5DYOTjqqAkTgFbCosYJByD2BhxmjPHn1iO5cly7EvlB3M5t
2E6VE5K4UGPLUI++Lx8p5Xv/PeW110/3YRfTTW+hbzC7hO6UgDgEXjNuPLaGPTil
MJL3oHmM53msbVCPLyq7YB4jL0VwEdJdoBa7OwAWf1Z81GqDllR/rnYCU8TWMisT
W/Aj0/6Yiqh55BbozMY3uhUBipGhsNpEIIk07dJwGybw2JQZ3O3kZLRJNAWkpxD3
JjzmqN2MPGM/uPXyb9Jr3byvfkulibiPAkigvtCDC1zqiifwAlwCYXAtX0htVu9U
qPs/+L09v8IyjB4yAKmW3emP8+4ErrrzzfU3WusooWdxaH6TE4rDTizxN0/EcPSD
y6xR6KumM4sdxeX+RbIBc/5VMVjdESGbDVQFD5UK0u7XSeuKyjRillZiVzmvI1lz
dXZYgZrQxnMVqrdC0hcPmfhi+/qeEl+Kv2PUUlQPfHqNN3UsNMpd9RDhksXjf2C5
JIl6+NbC2jYJeQtg+aisM7QUukAEmz2xSUYCi8wmslm0KU646jm9J7front5aHDT
rvL8uI64BVUT7I7VagC36H6Cw8Sj6tddGiTFRB4cpiJAzpi4NdNyYpIDEqnbmMH5
Vbcg1Ji3PzEac4H763QknkuvLM+KATpfMYeCeuHAVXF41HWKfHLtbZ8rziexy+HW
2V2YynfFpqzFS6iB4/EjWjuJ4NPLH9PToEm4RU6/j2EsIOyHs9FeVSGXS1Xl1Fdr
R7HLCzp17RbE+OutqVFnXGPcQklM9uWYnj9b/EUys50EUhjXDLZBR/+X6vhQ1uPu
Jm8aP7l9d5K9MX8a8Ua1k/i4XRTu3TlbyZrRgFBTZMhK3Y7wfu71qhmz7/T1AbdU
uP0iNGpPkLjfW+t05V8b9YppwQ43aEi+gX2grQ+vwH0dQUMeOjEgDYHM22fo3h+1
Y50mJKPCBdhHfPFvQzRmz1k0SOIHWVnYZjwZJrhSsEQJL3l/W/H44cEjKnr2IEuK
xhHUprzxBoNbvNqaEetJAEEjDeh/zVHKt63KsmUIKu05hOTKHbBGABSV0M0EzXOW
igMLHgc9sSxRQ6O1s+q6Szv5xYYHuWdMA0W3YxTgzLDAacPMJCF0ecEd1yQmmU3C
e4gCAY6xC39NC32+wX9uWTxyuk/6Wluw0ZDTAenGqR0LLLsi6w1P0wH2StH5zAVI
ouzvmaauM0gwfDeL2HLO1toxbiqCANguHJz4N5r9orsMiPrz7JpPeRsgtzFB3MwV
q2wxY541Rzih3clFkUN+Bf1Whi8/xVghWkurd3AQXl2Pnrz44sUvGYqpdhqCC5Lo
76wJdJQnV9YjCCKXyfMUJtJs/q2FkszKTn7FJz9ZWdxAVkdv+UPSr2oDHxWHYvg1
Xr3rwLUk+l9k6FC6cx8HaUe18YlzvhpKcsuUtezvyL61ymn07Cyp2OKgAcDkVpW3
ME9HVBsrMDbcfNsEGomtHFVfhBNy/IC6vLYA1WghxxtAg4/6mSuCkvz3MKH960DB
qgVaLZ09NpQh8GM2Hq284INL/ZVrn4r3oerbb3sImu9ptCSsxxbuES6k3+C6wfaT
iPPKXO2uZsJ8LIjfOUbQWsmN26AiN+u9KPS9g5FykhP45PC5lbeTMxkMSBYPvtGj
+tUWC7Nck4cAnBx5htzXTwJ+bZkMT6UhXoTLoyVP1A8B5VIyFHtB5ZYqrv+AzMC+
Ds0w02V5jV/06q8ztchC+QomMkmSNI5bdF9QArBmzt0SYcdQwtpxwrST3X4GD+Cx
wYsGBoAdn6bzdAxB6aCTCPpSA3b8ar5CyUQulgtsv0uL7zJZ9hINCggExmXWnZUf
18Xy6tgezw9DtdkRo46hdy6Mf1tA4DnBlXe3ZvlcWGTz0PnkEQC154dcPrIOfZ2j
sQulIe3fC26rvekNuYbHKTRtebB5PU61Vb+7zoUwMEXqJiBFC4wvN1CYKfRD2XYB
Pz4FuMM/2XVyx/EFb3WwOrKF/Rm5yz+9MUAnABk77jxJCQmk73M6cO4oZ4444YOs
bFunKwGLbZs/lttzz993/JYDUsh3J7o8r70ieY+hRMCOg/OpOsHE1QXs2gxELL2k
+e0LTivFJtjhdvl/78gd0V2zuyNQUxEm5LW90oyXa+zT2ASSdA1sfs1OMiR5vnqW
4JtZ1VTZvu4jo74EqqDFZ1W7TrXmrgxiSvtSY7VSowZxblCrqnG1oy4gugf6EAae
KGuyX/DgImiVuaubcvSpdrYiMlRiRofgQisPDAOAzQlmuStifT4LNPZmRUsoAEsU
NFr61l8tpc2fiRYHzPPZZ/95qOoyfWiFV7TNq+7Dsd6OnAvWIfD1cZsz7iERO0FE
J8UkvTCXB9FmuoXOMwH52QvWMNp739y12Y1qdiyT9G97VgvJRSNGPVScRrg19L7G
Ukjn2brvgEzuKxMW6HuuLzosAnselSWW3H7Ck3aro60bvJRkEvixH+qCXwDU6nAe
bxHqygUOUqG2Dhmes49b3H7dMho6LNnzgN4teMbfiRKL4Ai9vtUsZi9TY3hw0Lxm
kTwwWD4+mivmqfWjxXYx8HZBvklX4+RmvXFkRxW/VUf6WYcJBEPNXu8LlZqoCzC7
QlHr5g5PYg3ZbHVHyJ4SVW9FZ32zLSI0xR+w4HRSsAulYk4gruSudKEHyiOtfqxv
Zk1iyTXWG/3hLEC+d31FvrvM8rvFL1UzhyXz/CicrbQnPQRWoyJ0E8qepY2n4WYq
wQ+SStSzdoZI+I/tv4B+jMnxIiV6IFdzDYsgK030mjMwt9Redal2fYuhgA6MdmL5
jV6vHoBtY4hXwv4mF3fQfFYPBnW+F1So4F6wNE1OVrteFbAvVqT1h+PNSk9pLvMi
dd0ICAMbJv1UBSMsZN2r2kXPQ3URdxbzq3A75ovLwG2XWPtJdNRKlpnObxYhlJVO
4+b3tmF9blFxKh1FQ2qDS3zlbRZPPkxdbP/492DXA0u5LPthc9q3Cx0YP2kp65ho
3izEeDTSYvPs9EtHZsGFM0wjUzFv2ihrXozv4/sxzDR9MvOf+kE1ovxTW0HGEEZy
tCRCpClZ/DsHjN/FF8us9JvuGAbDHzHvdosB8Z4IDLd0jNLCqHNxXdgVB3Vom7FK
XAkSwzYz2IbRCrt2RWg81m1EsNYbeoAxIA8nnY8xvj21ENonOX6uwUEiyoH6sSGd
+lpesNQ2qBkF2ivgxCcxaAN3P6Nbi1Yr9tsyquzDPGnuaZ8WR2o9VPwPH4k5CpiF
izoWH7CDGvv8BRq5cvoE+hSBdAww1CABEqllDUW8hyn7pGslQkO90IdycNWooV1e
6z8RHPHiAq/k0ysS9eVYCpiFalHGEBefMqYf4UXNBfTSYgrEhbHCC8RxM9rAbvMD
Eq4W3O8HTNQXzu6Bw1thSSeKWbnRIJyNgwXrmkUBPGQDjt6ZdzNL7x2U2EMCqEbH
Vzi/hIkVHEawcXWcOzm5XI6vr6o7HaoFokWbAQrRhKOM/whqaDEDqbx/7duqXySg
J1Nx0ScjLCnAfO/M9+0eyjPqUIfQTmR/tCuYAbxU/mXDWUr6A0Eexq0bxUhDiuVg
eqxNTak7Pxu7aCV0loKiWCdAVqLvxTd/XQcMHcxBGsKUAKX5bEYpcxOIMfCpgFj5
od08CmQ4CqGPmaQLhzW8BKWB2qaCAhrfzhAV8TkcT3J+aSyMYrMNt0LooGwpT25W
TbYF+r+eSGxjOPGFau8tEOKNzXt1r/jLdZ95p2SmqGFhlUpK9mbrxw85sLGtZHZT
btQesJWybb+2rR1lTgE88SdXxwHkx4qWtw+H4XfkIQASJl8C9ESHVVkdhqwFjKNa
auumcZ0B+wND58kXRyzUyahhqsEcY2FCnTQ/qH4lmB2XjdoiV21C+PNJPlW/FYpL
hsEKNe4kiIT+Hc8B3txd638iTcoyON/NEjStDYjs+M7kKwxH02Wob/B4y64xEbBT
FZQec7mLgM1b6EegiDQ3DQzyanz4vv3bWp+hbJBuH+Rtp+OntrOzTdUbVu8zIDaq
azaukbKzbT8E6p1MuXaO30/fdj8k+EuU213ci9WWdat9snapqGf2ol/OUtX/zK3/
r8U3h5P/CTQWJqYZamrGVV5GRdwBqBpoc46PNtkvg2HfKilRJC/21vunjBvMtC4W
eOYpNiGhccgSxEDEHV8ujY4waD90AUibGJOv9uRAvWBP8k3jMYxT8b2vbxhWeqsS
/Ql1qxnJu/vB04Egeu2tRYc5/yMCo2EhUFgMjScZjNmhDRYFoEriCpnqLb5WLI/5
l1ekPi+EiBKtb7qBP/wNZzJQorUG8jRwA862aCIG61Rq0Vh3kRu8zJLQ/DCoA8yf
19eTiavrltnUgfIidmgvVckai0MegXOJANbx9FUcVs0ICrOkmHR38En+yK2Hr9Ze
mqhYBO2xVRL9KmLsImCw1DPmb3YfyAJd7t1L7vg5zixrSJ+pYZrjfgT8ft0KJHwJ
ETCHkseL+m++OrhjlV3Z/H/kEyii7ML05VrUmLQwlnPUSGn6r57wp54GvCmOMNxl
YD4+0pDh98n8PZC2bT6pRb8thdkC7cl4m2l60S5UFJj+EqzSxyaqMs6rnvky7oKK
MKqYcMpXsfxCszQiRAgrQDEubDgI7XIKV9vqQP/4bx2xARGsqlHezqWdyvGNJjR5
YXTOeYSuFYCrmki0b3SXAh6CPTumuMbpUOylz8TbtgB3hKnL64wqPtr/5q6okZkx
wkH0rBHOVw2IB+rM82Ys52BDkQsKN928jpXb8Tfd3DNhWumbaSdIeL1mP/uAfgO0
nePs/OP9QjF1qgSc9HZVZ+IwdR3Inp3Onk8/PH6+rNbF/GCsl0sexgw4pl50O6y9
O5+cqNIisinoqYzS3TDPO8Tbe1vdZqkoCLu6Ijl0eClpl2F5TiPEon3CtfkycO95
lThEYY6zE9ajfsphEugEo85BWHeWVztUKVrttiLg2JnkJEOj5pvG6ruGmhrdPwH1
smnuSesgJn0Zr28/AQ7YOUr6BqHvq1BqWzEDmNCqsLmEI2myw58M176b9tE9JuAS
o3TSzuOAG0Ara830j2QhKxTeXFWshfD5bhkUnOco6o5AclfT6GvBdaDNmBy0sHEm
diskvUK1cmCLAX/6uNVTIBCN9mxtCxAo4YMT5IHBsfyYaUObwoBG+wbFi1UQDSHz
B6XiE4FGnOkD7r44lU5f0ZCG/+79dhGc4/17txeMx284fFcNUQpdImpXZ0ddzWkc
8QVu1T6nCQWAn2quIcrrUCsdelWGKbz+wK22jqHGKfhBha1YA5sfHJm0/dnzmTOH
+tsME90BBcqCi+y+v3HjcHJw5Tgiy2C2cgrUqTQtMYH+1YuLFWeGOtqGw1bWGIaP
DmWwogWoMj4SYAyZYdaVhdKcpFMwajy8SG83xjgQ19M6YaCl/z+hYDjMSxgsVmbb
PS/4yqyLfvD3uIx4eyK9XwiHFJVbhWsHVtxPK/bWUEuN2RGUuUeBxRbj+kXDrTj3
d1lZaITulIXpwxk45Q/kjnDD/EMqeJArK3PZpyEoZKYOGKPnBQJjSzVjRewQO3z2
IWT8zJhBC+bxLt+7Rr+VmR2X6JBgYBPkDs+m9HhuOkeKrM2PqKeL0x16Bt7NFqnh
OAxoiLH4rUyQ41dUUaF6mIAvRpDW1uf015qvNul2MpsfWZ+o2QX4BgTGAS+K82sN
B2D3dEDponnYoBlUfk0XZjUNfa0ed01ci0db8x6BIVPM9NvgKiKQYV+Q5I9Fiqbg
Oa7J5j0SVLdENwsxEe33szKU7tVVPnOyrKPl35RfTTeoSBpJSnB4kjwC6ACsTJAM
Cwa+9mWdeF7yx2E8YTj4gihdSX7PkiCjYbgkE3h2H6aeoGDv0Wo2CVfxToE7YfP+
LYRvYJR4tRiz8i02v7HTf7a88bm83WyD5DpzZEwmF9NZBbVQyEH7H2ynb3g00Idb
A9kpWxm+rfjRJ0qjMZJhKRcrnTCzdT6FOMe+UvXJkr96FGi6ai7Ij509OnJGBhQM
a0XehsiqwBbYlDykvlhdewMgBoFVINI8LMbLqEhqQ8hXT8jmWstTThmIrcyaPjYi
H8ov9Hr2Q7Um+/6Xneq30qA9cIZGsO5vGrRlUWf2oNDGBnDV1hgO95s0VKTyMna9
QWT6sjVWjVGRh9iVMxLf6DCwY68VjVNdo+Tyk4+9GLakg/qxjD9sAkXvLGQxLSce
55QlgkM5ljJ6VUE3K/30GgFy1hEGTxmZWjiyXtifJ/zIX36WRch5mvf9asewyZdw
V/qIMIZAzVdcqNjny2AS/PeIQOEyJv92Xn2DdCEQjxodEiuZ5PzPXig9rGgYmrR+
5mactTXByqNHUcusYkJv56Zg1QqPlH+IM62BAZAH33o+lvv1eyqptNApR+wWYtpX
xJBGQE8LasmWWSAJXYNHHzp90PZqG9ecaxXp+FhPifG27ef50JXO38rrGm6zuP/s
SvJjRnYhpFJ5BXAN5XOqsIwgmDQZTSkSab2lFqUXVucfw6SnhPUWNWi4677ig/LD
WeMM6kkZQo1MvcJ6+TrjA6oW5FzsaUb6NyuGVjiHsqJ/UzNeimnHxjgAvQHvjNQs
3795DD6FOFyPxZAzzdw0P0YXgeZegwJpoPb8wvbnb742Dski1NtV79LY+H9ZW3+a
5UgqehCqcWpuPTYvj43z6KIAnkw4Cppn4G1c8elrtYpj0X+QvMeBoQB+rzH+rNQJ
qTqljXq5SYrY5DEHqoynbtSF43hDQ4JaJKu+4C8w5gqLPXYG2NYzbtLoFYk2yRWT
TsR3z70zg7ZAXVRGHBCxcmHTQN4i40sNDL1Xhuuowx+PKLycBdaFJlQxBng9DHPR
Dyq2UwGg6OUt3DlylGV6KGfemXMVqQAxm3BE4Qw8kS09Ml9EBYWLICHHfrLtm03e
AxK80hBuSgiwWf2QgEOrCA0VeuCR1zrQTxzM3GlJxftmkSYOhFTKJqYogfWcI25m
kzR4RJKlMccw5qCkHLvtY+iHIVcDS0XuDgyz6XcrXI1Ty23Pple3TPs+h8ivNPTi
6NnY8L89xuDBcKNLKhrtqzgoN2lRBug+cO/4F6BwOnF4z6129Bgv4pyEORRub36E
n7LoLVukB+qxAaui4cpX8KKJQt1Qi5wP9i46EkZ6nh6eNbx4NUzaUaCIcTQgOgxA
rXlbGQWHNL3/KC/DIvFgkFm7hnlqEmvMn+WXOG80+CfyT8nSqvxjGvafVOxquqcu
X91/M7nen8KvWlBFky2UcMIjVVRk+AVZJ+GOBeevbXuqflRnecMszoZrQ5In0OU1
tw3LK3U8ZLMHC1WzJhu2KhgPj0D1ERs5munMTzj1ROQNLDIo5w6KTG/M5YdhVmlb
kKVyBtYQRE52mc5UXwnugRtP5rR9/7K83ZTmtNm1wMH6cuAMctoORVluFsypjxoa
/YIOkM1nBqFUnC0ezYu0JvSbp0cdG+E2UJds6Cah5jDgMJvu11+1LcC4VW7SSSEV
nEFf82coO5vQ8Gnc8g5EirBlhugmtNlZUqkD59EbOCbKFEzZ4jhtNQ0BD0cbhT7d
X/9/gIVFo3ZN/6+IMD23VM7hqpPwbuuT2NkatIulZwvTTFdIgRG87/7gj5N452uV
2fj0dBK7QVOVf4E5Az3kAxqKWNQm2RLZXwldtJ+txP4nfw8EHGHZpiM6xE5XQy/B
UmJY1CqZfBi5/U8aQDsRR2LieEKeUg2kfXAY7SIe7tsUiSPTHQGWB8HSeRKjdOrk
0uCb9jqFcJqlznnz3ir//5iAybowjn+qSV+U7sPpAwVQRZ74I34gxqR8vRpl1sNH
NQCUpxxWDtBtDfWfOQkQ1oP9UOI5087aRydjJRHy216UbtQ8t87Pq0ozVZ6jgpi+
ubn8jcDnlY9h+d8akEJ/1uqBFq8uexnzhj00ztj7hZkIZUIjO4sRvDCGfhxplNGH
4m/xFFXrkb1Y8r+OvdAHUSR9HkH2aP97XZBpdXMhiCQXgVpoiyVaK7KhSrhsOBFs
9Ut26lulqC6BV2lGZpZVtQNfe5n36C/yMiJY2nD709WVDs7AfwaV8yFMFgiBhk80
mpMrTmT++r22tG35Pjvyo1C95VwLVNaw9fvAU+PiAJil5ZooPk4+yQ9sYgI1bACB
ctcK4fHKLoLxnCI8zXsbbKbS3a/cTT85VV4DPpU20HLPP9RmorX1EDVZWmwfKHRB
uErf2PbD7DBTtHzpGZ2FDl3Mxy27NwNAmBR67gFilJE8PUUslG3nNJpkNICzhHlV
pxCDmlp5SA//5k99Z9J72SNboK26CsNwdPI0wLammAdExUEKcGehTnw525aouUBh
kcbogI42qMS3Eg8qphthXd6OcFdTwzpZVcXR9gCeU9LyBRyi6sjHb0GBAsohO73o
o0aInIvImFYSJVT8aVnVQJ3JHwfZMQeYRZ4bMHjkis/GAENmYazTB7zxvCUYh8F4
gS2Cho8JPaDcX7GCMj9v8NZafi4JiZjwufULdhrjUmnBYx+BriQKmPLz40sy3ByB
qCVCxubyrITp+r4WKVyWfyNv5rSyD5FCQLQOd97MffQMzlS3hrdGEGre1Txl5riQ
/4jxolDhQ5D+fo+K6M1vhV8PN4UHk2QCa1u/9WXfIzm+QQcDIN/8XZHESEHhXzky
AkZVT8zINv7RXvk5didEMjbwkEg7zIh5oPhsDwXHa+zpXweHixOaR63RAk4C3dGj
JnPGvODV/X7jItUnEr+Xx7TRheTAJ0FHMcvAYKFBv5v8q/7ybee5soOIQTL8X2R3
z1Ex0GUts9YU4MfLQnE+8QW5OLyz7l8+vK6fTlfEsLpVmINQteQm5ategyCmv2sY
a+qZ/Z4OomFHDFVeJfn6d0S8cMhJfacGU1lEUbKeWi59AsmbgE5k460PpYdzv3XA
IbFnrAOcix9Yxexkg7tMEW01MiKF5dOY5XbODp1VqTfsb2nbQcdOLMbGIOcDZ49X
jdcOyLNKJ9l/R+R3XmIxUNmv5q7QteQN5S1F0Pv3vNkyJGYmy6gh1fqlaZ9k/7Jr
R7+2TVKEVkfOgC7pbTGm7KJ6HU73fhgJgMsEXoQ6D0v+vgpBheQLAqqnL7maNflX
m48b8td+DX9bVSGPTN4fWaQuvEyuO5Jyw6xvZBSpthi08kNpva396gyEUisf5NnK
AeOVoYotw1dga2UEenfqUu2GcEuZvSJFYimpip6ZztynDGJNZDb+nhyYtnbOMEnE
Q+bQ6jeioDoN27yuqON9UvuF6/FxN3EVvNcIZsuVfloOTixN2B5zy3En4rWPKiPG
hZ3F6RlJcY+i5JzNbAWi/mhLLLgbF3H0KiAyPGs0RHBBGuNeG8pM78/DMkDhpCEF
qJYlstB6UTa0BQIgb+UGgifdWzkCTdeLmpsgdoBEDwUusRGoUlnzrZ+ENe6AWyQb
AWBSUVrOXbIiNB3iSwbB8uHDP+ovkSqhns5sjxLkDBsEdfRHlQIw3ItWVDuDHQN4
r/Bzzg6y26SvkzR9h5DZuPyOvOiOumHJPi4XnX0CVGw2qwN5XU+I1owRaH77fjbz
Ptz3CQSLIq0KYgREraTXQma20fvcAkGxqS4avsnTNuaKY6rDY84OuMzqUrko5Wow
3Xq+fh2pGpC+8b0DW0gjj+2ZesXyWrMDvp1MxDgwekxpZhsIffOW7ILf+7YzvAWa
ImRd3/UkKdtFTLgvmOaOiG3+hIEoKB6w8G8rZ0YcZGzACuI60mLxcpbeehf2fGJq
6CZh9daLK81fRrE8ZT3eRd+eeh5XEyI21WIS8UcHyEMNVrODSp8qOmetyh91Kxj8
BBgQ+7bKBddpAPJMjpAprEWOHODCmpwPRegQTg6zwM5hC+kC19qDr9UmAeZ+/SrZ
HIxi3rl7pK8eLT3an3IphDRRBrSGT5kCLq/QmLFBUf8h0tET0ZyX19qugNjlcoQ1
br9JADaim+l0KHQaBh8VO7s6KI6sLvFtEp+a7OfcXe9EvGP+D/Q+WHgMgyEa9cT+
1yf4xSb0HzuL+/SAPyeE2iwOQmacCsEuFKzx4kG5zHZ+wjwtf3uLpzT1U1GbDBb2
5q/nEOkCgxMlvItvWv08uPzAFCQA3FnCx2AxlcoioHAnaMQm3JzGt04ySlW+u/Su
9VNFYNxwjrlVm9rN6F2dDkT6nD4C9xiO2W0l+HAchFtlBow7tO+XKsTc+NH0xIS+
UVRI/l+1jcthZuuMQDlpoZx+Mlon13usKjZTz9EB3QQDl2G6fBzQ74nOdWag/sx7
xaHdAgIHuegqm+tKzLVIQvDeEE8RJE9X4UcJ5ylpTGVtMfctwKjQbRjDTbkkVOra
eucTL8P6v4n8HxfGH01SNMlaHXW0QN+NadRv0h4H/r7OZneBUztA/jBs48CrwM0m
wZ7vq0colRtpvmxPh6dMhzNDicLtn+TVj9VH1SY8b1Y9Eb7qdLLBG7ZObiZTbNUF
2wqjSbzS1SdCZHTCwS3VLB+zZw95w22ZNyMNdYRbm6zV3jc3JwLclN78O5QEpNKe
l34umLAqQXFokPxdkQ2xUxYb5TcePSqqKcmlhK9CYTOqQSVpccvLVAdk5unCnxpL
EStwddQIJRdDJTk/VBKrVMltpMUHgP95VN+ovXbRumIySnYouPMo5K/Hfu4v4P2O
BA8wlbt5co/+mzXWN32eufj63Oq+ystHURA+zYrluo9YAh8S80y/MA/g5JtvjOc7
XbLFj+ixPl8wjaglpq6pI+5BV8ICv7Tl5PGptFOCeLsFYVyoOOepDznA0GAxnADs
dsWG1AtYTRZUOvIwZwaAwg7QMF+9P+71qtdOG5DsAoCa69LiJGO2GMrx4aUFSKnr
7OX4iw6AfIEhayYzM3qshb93nVIyksup5NXfS0XiIxEda3ZwLvgoIGUR3Awz88dO
ox9RJczZB4ySOtoVXasA6riQYc6i/kRpMQegnIuoSrAEzETefB2kLQVlGjROFgvr
uUtYajaffet/alG8cBJI6vl9DElH40ULroUkxKrh0fwMqc5pgkRCQ4UfJZtcrJsK
qqhBCb0hAoIvIkE9XL12BAmGmtRD8w36JPXMSYjJbcAEjtZMaEvjmcqW/4oG7oWU
3jDUnuRXTzMbBYRfBX6BTualfxVaZfDCBKQeCflre7W5M/dFnh1Qyy61Tm7Rq/vY
wZzH7HqtXanLFODdWrCP3cV1zm9OL20REz71Tt50Zhb84vsMYcQJYH/ETTCELSig
K0G2L9/qg9SDQ6MyMJlWMkCHuExjYJjd9vNExd1IYS0DPgQQ+2QW2Chgt3cgHd1e
JSmWzhBNhjQqBrEEBOEoWB07kwGW7GZkSobJzh1WA02iRxrNeQ3XQW6sIStHVt2z
kKYO5nj5ozHKm8BeXBHMGmoGqZNHNJTwvghUkHlbmrbCfg8JFpZscjc+QB4H/5Kv
RvVkemKHfAPgJa3Bg7nSlb85KeLB6+ta15mOtCYG6MMSNoXzI7k1eSDZJ1DrR8tR
5zl1G2rUwaWxzRMWvBmC4heka8t2pPXgxQPLudwzs1ipx9rsPbAzugqLVqS1ugDM
NwjQRZw/r8Fh/kOx7eujLuKI7T01VwR4tyuFi6G8xTQgigjXLvtTPeVSFjRCpSKN
LVQUzlksufRAkxlYlO/DtVMx4qqUZC+J6LbTGJjnAUDjNYXibdeTKcXzYz02/zkD
BbpINxly1qW7W8UHCFyrZuDBKT/tNKHgXH9Ugitq08wv6klcaQNQeIQaaaVeKVjS
I8IQqYdD8xSQNvnaiCEV2g1b47jIMtq8qWZ9LJaSAqOAl+1i4HYB5TiOV/yLYjP3
9RXlws1WnLmswoNdeb8SDZTF107GDGzQYs8TpiuOj6NzVd/BCIvGQHw5P3IOrTLq
2zngsaMnSHaGmp1PQHTV+pwQN3WyQWDylVEYQ+EAr108yF7SdRs/fm5UdsOz0P5g
vvi/O2eIRtPmQPH07t44nQO5xF2sv7jaVT/adG8v4JKpi78RJ5TJ3K6swNEMFrn6
AfYV4uQnz/ZHERePvVgXBze0RHeoVVPQ9aL6ZjDmMsY/1xRH6UORq8WFNf2nn7Gg
Np4hn/x6qzoscu4V2T8z+z7OibAaUsfvh/8Sc7piHUai4SlyQq/wTC92FI6bniwa
wYiyfkhVz1uMKpZd2xvd0qpP2o19nigBsT4B12ve+k4eALk358/oxCgAQeD/cOMU
bflF65nv1/9vRYz+6co3CO9FuqrxhS+jdBt3qTJ90+C7PseS91d2rrlK099NCWmv
lifHHqf9Tof04ioZVdFVh3vgZWvt3TCRlmkF2PPBNn/dHkvv0+7Qj3bLEA6ZXyuy
04ar1Dlrk4GmbCVnPv2dtXwjN9DZbe2TKCHnEVL5u+anAuqHNheUIlCYvcCyKMHL
hdNOzQzFmmi5MmU47CeYfnuuFvQf3XbKfguEfwg2jdDbmrXBniKoRH3N2G/4i6MG
ARabXjtMcp3FMLAhz+ad6VjCkaOsOWGCQtAozz/l6HBzpWMwLW9tmR4dykx2ruCS
VhTEBsLNd4aXb4hsCS+ooVO54f9cpr9EGMi1AZkDsy5pbXXB/BaJ7OUBgfKGz644
dvphCrSDvigGI2+rSJsX/c3ENna3BNk+yGM5sB+mDKWFUIlAmeA+mmm1k6p6qwlh
3cx/xZpcU39nc2ScSe4D4r8LkBdnj0b3kJ/8g/6WrZKhkTDhFFfLQr6qcreSdbRT
a8+9cAiSDb2gw6bMkLE1jFRtvEZCql6eAUVC5AjLdHkYQoVuRYIPQgkRxXfTE+VZ
hrfTUtnypF7SyrRYLtxtrRpPu0wL7T/8Dzd6w2/klfcuWLCZswq/bmSRgiRoQN/Y
D5OxBeZQb94CedFHUlHfj6R5c0DzL5L47jWj8Q288FTfyR7ysZ5NOa/LBMz+gc4+
KHEylgv/QnodftXNof96aANGC6YyURiW4tWylTEezeTSKAQtO+g1JJdxTSg/9UyO
YbcsZzaQNrPN3MeRX1Q5YJI4OuSMvDZR7ifd9+ChFw50QwXAItqBru7zoMkY4JlT
w4HXeq5dx/NcPElN7WdUVg/rH5AfSPaTSBXnGBKM/Kp3O22RSyImSEROt94paCTP
gcg4crx9rarrxEH4HnnDEqpIP2xzucmPti+SmiLyLNU5a9jTYPjcAO8vlEuOY0ND
6bU1sdPDa9pXtbUrAJj5+8tmMQZZ3beLhdJpN8hSrDSClz4faSb7zOYoudkInpT7
7qgvJhoDRTNrEf9mEXv3+GXCjgTOvVRYYu4aeW8Sa5+0/7eM/e3I/y5ZofS3iOJY
Dwe338jgQiWoFgpDpXL4wAAEdWFrJ5keTGUl/RKooMoSGNczkRwexIEXbz1aQfzk
RulCiZbGkDuyd6Vi2eRqHELRn2JnftCQfoWLXWG4kYr0p9LiSHqTwukmmhz+LZRO
IWMgoNq7s2cBH0zx11fG+qQoUIZA02uZqeWWgs/QiWEJHo4ClMaWdnhVVvoND4wC
AkTUvjXjxCgRlq6zv10yTqo1V2ureC6Zd2n2SGIoWBhI1xpVKJ1hKfq4M6dXSLZV
tbrac/+TUR7IUpCw0RSCfGXyRvqhe7K/JdqLHGJA5y4hppZ+FmOLH3iblClmmZpc
ueGsXoKHgNhchXyQfFJIA+I4XQbjWBHBuqzFwiGXBHgt9OLQr02mP6sbBJlpA4Tf
NEHj8F0fBaAO8v4ein2vQLecGN54FnFShKqyXpEJpJcKuuVg4TFUuk0JtoTUhj/T
bJNz0c8/08idWc6+/DFXAR7kBIeitEO4ABwnF5TkZ7BtKFrrOi7mZkH9KBN8JYOz
7j13iX8DqB6dIcQaLVKcL+OAylmSqKR2aZr51VffTcIayhadd8E+ysdDpsmIUWCF
JzBnN7u0eMLteWctiGmP2kXv1hJZGLojy7zJCvodqsUhgms/Cizs/y+do048Moe9
QwItYCLu0iXMq4t8x55dfzJ/MQrN1J2ZMjzyLNd1V6FmuDpkNM3PAFIA6yxC/+HR
Cr/DyFT/Lw23ehlp9K6YOrcP+v4WcNO7sFcwpox7frxhhfq88qJZYYjV02RWiitd
nJS/5QxfGVk6xcduN3HJHqQbFEjc2E/qlH78sbZVolD1N8sET/qgbccNZOtqYaxP
gP5QLijrZnWU9XOKSmDTupj9XWJWioyVlWGRl129EkduMjSn+oCYcxTFDZ/KIB+B
CgXG42oowKoW6HzCShLcqRuOeWhFvBhWoWYzzXV3QM3iGD57Y+my8qkFAZzKlyAA
M0/4rl4TgQgkh0GManuIV0mcvmlRvJQwwBCLTBnY56EH+dJ5i6GZwsesW0zZQON1
yKD/7otQ5EpHGcoE16O72W/3wDRJ1F578TEGB5fyJq/TfCk6f3vUC3h8+LE/vsvH
Qh0Rn5hS0NbgXraSlq1cdpfWGqEQYGjq/7a2T3vY3i68Y6oeqlhUZ2zJwAG5lI5L
CI9JYpkZdBuDmk+lTGr1bjyMuEVqzzU8ClXrf/G5b27UUtzrLXRbkiDhgyNg+vWx
UxBF5kZrGkULmMYWZKTMjhckTGlqxwFpdMCxQCSHaJg/IbP4lrw5I69kIYaI1uYm
uY9oGamsInNx3LBh2hbJ8aHQkfHmV3uw/U64ZwiqJl7GLMMLfuQS6VTLg5jfPhWC
kojIRq2lV2SsmfKie8/UnOIHlzN0aLCXxuGHg44AIDHQ9qFQEqy+wLfhWAPqBeVG
DTwBgp4WtMzq3pE8vcDS5NvMKxfUN1Iw8+JgeGLdkUJtd5ta0N+xcwocYYpwsscZ
n1Cr+RWSfHyBMguuZgH1yDTRGNGWGKKvT/cXe1Coe6IwMaXIFCF26oyZ9oslQOm/
Wz8L2/gYHAC3TWA85qDM7fLurR0jcz6h+pR8zOiG4h1l8MU9NGIQj7Eti4qAf40a
nlm5BXQIKQGb0tBNxIU/CdFZvmesc9EsLIkmAF+VrXvw0sUl8SKDypmxcDVZyDGB
mlDiViT+lYMsxPIPwipjn7jZSA6Ogzqxsw8FaYlpAeMh2QAnLMTA4f3EBIPji2Kw
4Hv36UyIrIZICAX0uTxRLid7YfIVpo9m4LRb+OzQjn9JkGWfr9K4ZX4C0lbkeXhm
B6IkIusKBE83xFGLGjuuHW6cD68k4iI92JvpPpOUELNlcLoKQglu20dZ+0KoGNd6
2LAhpne1YKnU4oOGhbIvOygHl9ieAJts7/E7YH5aZgg15XAIC+Oi69Hl/zH+3+li
LjjvEKlbfBrjVo/rDcH48vaqQajQPgIXZYNW9qUmwVNAhbdkBk2bT9m96aPSEP41
E0cBY2nMpsi7JLaBmcJ6bXyaxJVTLHjbGu23TKmfyzDxnBkLvc0etesx1Wmm6W7I
mYqw4zO1OkExiIj4xqnGz8y0e2Y/s7PrhRJiaNaLtxUQWe2JOQTPoKtnZVbwSFT4
nkXYb8pUmqYeTN77uJ5Tfn9wZVTIBciD0iqyR+eCzpIaYbqFnFM2EtInMxfKO/H3
Y3EHP85nYpnJFmCgKFbbFUA1hviNTkRFfnzXp3bUWgVNGBUNd9WG+jrZoUbj2jqi
EHYQv8eN7XQzNz6EQcU+4zDYI2XRCG4/NrYm75B/4wTzStfxhydJQb3tVkWKNNpZ
KzH/ocfEI0ak2YxCeGoxeYeRpuKdsjP64rSm4PTnLYgSeM+noAsRZGQ6iEL9KW9M
gWE6ZbWFbBrGIG0Q4yda24fZt2dNTEU9X5wyZLbPWmCPHAcVIhz4myskeZ6otDkS
PQ4nF1/nOqS6vRFkkUwbAGgsSFzv+lmhoF0VJp4mgSbhxpbjTVYHff0vyb1qu9Rk
nWZYmLtzHG+wfrrBhDCbS7Ei9v2PZBwltWd3ETU9vvNX7nnsCLn4T19wK9/Y8cpp
wosfPoyAEdySOB16pbYKHynT2R2Vdkax/zG+Js2ig8Hqc1FZqRZoF0eFobDbMEp2
BzJLJDRbx/kjVR6qCA3cHB+OOoIhg+rwbNHYY/hglHAjeoqc7PV8w87+b5oJFkNV
swk/O3ppsU2Ma/klRcTXao9t4Zin/6cpZlHF8V2XE2swyVT0qBhJm5eODNBDQKv/
M0q0ArTXVdJbjJRRdMOJIOhXVfzfHle9Lth7mqOM6iAeEBU4/a+ZHwaDVp12K+Zf
oFFqyrjuSzWPjMq79zcvs5MHf4rNN52zFNHgjP0/ezX/pAZoctNfUL1tdksah7SW
X2JzP8/udm8cZ8gMPak1O+H6NVN7LF3TOgZmJ6anBF2flJQtFULyJAaqee3I8fIP
Q+XQYHJvSI90e5V9S60VVjBJlC0dOS6bV/S9zT30E7DRiB0a3NHNtUTzhzQ0hpws
byX/871pKOA0V9btoXpAYZ5jFV10+VKXor+MiAVyUYjGxrrz+OAHw4zoDhHGIHvL
B5Fi1FD8V9qI5fktcdYYtx/wbEfxJq+K8o+2xYbOQwsc+SupbXxjhcLubdDDizv7
yzgkrlsuYBD96QvlzIdyYNzq3SqTD4gbVBJbYs10oxTLi5H4ASsY1/T/J2KsKNYs
OY91n3qwrT6eqNZaPSMuXmk+T17+3+Z26wS5OLnLQgNRDkYFJdahmva3eYq0zv37
m5feMGOQp5ZyogPEq1dWyphY4tX0FhFhTR4F6NxLjDttW8Xy7sRwLUKw5rvjVjE8
r3Y7cHlbrl8DtcTMEN3YBwNJI3Fla+oOAQsRNsMCHrtJvKvIg1u7/9zv6ZF2C17f
OMY5oulb2uwHg8mxPmzu5O5t894FbI9DuIAlx/iKFaLfx0FAjefXQMMEsOY8NJ83
+IfprKl4CJW8jM9j5sbN6UIPyhFr8AwBg0Ce/4/IXx1JphjSSoJKkxmWVLhTkbU0
HMvUH3eQNIfzTcqdkkSi1tUNYSjcPd1uU6iNKydIvHh38MQ4JC8ISBjb+uxAQtQa
gMgEcBvz+DVI7SouyCkrwec8DUv/Vb++BtmWjBqRs2PFFHsLgPjZVZzmuEYmzXse
o3NBMv4IBJYTp1raQ1GQiKelR7nYGGQzcXYV5dLtmLuoN252UutVbwWYT4lIHjbn
wu6YIJk7dXd3aHnuptkJgw51h2rx2mpgHP7ZJ79z6SGQ2H9M6K9/VtRHDVU3XfgN
YYwhZ9n3oA8sf8lUNeL58Y9sltvAv2K4Ieo5vV3ZCu+ILGN/fJIsmoUtPihYJYcg
jbdNihSEv8n7ctyBDF7R+C1ejuz3jILssC9hSp0Do9Pav6DHHBk45/x/MUMMqDwO
s0oVY67ykxAZpBZubNqh5h/PJK/IOYVmsJpjSddbNT0e+qQNdmdEZ39U7RrqQOef
ZPm780ggkxNFcGXXG/7DbLEm/xaRdJvqceT1kUxpnzjvnuPXB8GJiYEErw6Ticbo
xn5kM2v5Cp7pdYTqhkut6ggpD/JIhaXM30/or+IhPqK5B5gZJxBdlMj7fxd/JBKb
3vDLtye4m2Xns+kUGVsWM40abZnbauGcYnH/3itRqkspDNVr/9tPNk6LpVbAgEsK
qcl8lL3PupgOX1pDfyqYa3QfuXfxh3tE6MvrF9LMEaSjQLkJjBT16F8rkAiM+dQ+
9Py+xbl4gBQ+/Pilxa0TKwnKvfvK0VkfZmuEh7MCQ25+uwWpARs0EJ+jjCb/LKq4
nqDbA+GjONe9YJyx5+XH81/mSgGvtOJAknAwCDck5yBtN4028+7b/pBXCr8ceDub
ZGH02iR33GOe4iHplHDUMG2cRO08tj1HFeutVnXUjLISzODciU9+iOnm74MsEKdC
OZb0DfdCB3UuZW1Lau42QYMmDENjajeivLK+KwK7gSKH9Ix1/xmGp6rbinrWliHN
QLL5pQ63Lsg970l3OaJ4agVt099mS/rSKLci30yFENgGE33x4JyX4cfO+7yl95O6
FptIYKsWNIHGpCb77LOW0v4bAffow+v0GjWkSUAcP9Tk/dMD19PiIn22VrypH84L
buvCVIC8OpzCiL0Q1voYrt4QPzIYwiKmuFOdLepazwhJvjjNwLS/wsQZZgC30NPh
7ia0jwB7/6LB1QsQ6xkfcs3TH6pWAvfsfjG0N9SMUqmo82CVKOW7iZOyvh9fZoaf
yXkOjFl0zFS7C1t5hI9cdb0ON2avXYF15ZU1Dp2ovfiHS8FRJVVS7mb0gi14IR1u
CPlLUGQTs1w6feCk0hdCvZbDpQKzoGKWYL8LjHJpSk7RJGoTZzk9R1B4nlTwDd1W
RZvbpBb8bc35jamhvJ85Ys17uVdM6qtTCMhTgmHqayJhkeJd7xl/9Cn+AYybbIMB
0f6Fr5vjys+9OIs84ghMBears3bXEumXKyecUQUQPzF4FnQC3Z4NXvvO2nwofpm+
Epm+HoRGhtcYqSJ4mXOQIyPiA3D9V8vei7/RQn8MVHUZf7Dp712taGyAnX2i1WW3
5frgpzznfZ4TBYQbrCvsMIWUqxfDhEpADv7l1ADf6oHKBSotl02sHuEKeFzghMpa
JSSyJZVtnUp908zxJwHC/bZm9O8ru5BfQgTolkUDBYZ6fcpPqAh1qrNrUJKpOmHJ
m7oxwX3xM8OWuzcUz7jCHvaX2QdSjrJldqXvEpKG3Q2VjxpKgJ/QbGDrUA8Jn7IQ
l3APgHnQMqRGDihFih3HIO0LeJATXr5ZfY/IcoYLEX6818UpBoMNvrRQ/YSenEV7
49WKp+4Net8uZLg9ZvucXvQtl+rFxJuImuwz+YSvqr14cylZhMklwYqbWz7jd3Xb
T6oCFOAstLz9s7MHgRoYsBsrpVjtk6G+5bbHcBE+LnYLwwXvn70OE3Y+V9HdZNhh
O4rwjjNy4DooUtePhsUZdimt92lGp/Qob5MusaLnLo5wc60zxoqmcVdVuyqA75J5
SnuDwvQIheBOo0+WxVfmyHPaMiLI343p2jpKJxwnUaLQptR4bR7o2b7LX9YdMalN
Ul4GF2D2LwqOTAvcyWjb+C7P2hBlms8djClDUpBIaz6fUJBbiYDeRSCLlo+Zon34
6vPLXGk1VIb8UK+URGGR+BIDhaOy7/Pze00VahGDb/7lRqtmKuQhfWAZ630CIy8X
pvF34L9pc5fIwOrujFB1iWmOeefT5dqt4kZQuQfwYQtmUVp/cj/VfJPgEqdbgGRu
eB/0t+jQc8uOGXoIoMTdfEou3SS0+hj8IidmxGpaSYKR5m6Z98cZkXmnpgD9ZFlX
9lxCrXf3n5c8LUx8b4rQOtbaIq0puNudZ3AbKJtw/GBi0D7yKaofu3g2I878GySf
qtPT2tr1VAlW2XgcrLr7RcPR8+b4luxOZ3/xTQGs0bor4SGKKvFXh4+q/38W+dmI
nP8OghMT1VHEpz3iUaWU3XZRzOt8t18TDaEN3u3IEQlZcPxQS0zIDKtMBc+XDvEC
xZNkOd7Lm8+YgQbGGmps6pY6AFlY10z2stf+YxTNR1w2XoU9He/8MNpO1ohRa3Em
Z8NWhcEDZif5u1IrPttPwtd0Lo0WFYqRrL/y8KX2x7+KiUceBSYCb0GZEZ56uCuA
av7V7BlcknWlNGDTASUai4eXu4fTo5DkZ0++JXfDaO+Efg6IS5wDq1BU9Lmz6tKT
A4dQGlE1Ut+XIiuTDrw1N7CzFDJ/x7xSuwOH0Geyw1j7ANeGbPPz+1wMrRDihbC2
QOHIiyQ2ENP30ax4NICh28TF9RfQvYUfhJeH7Mj9Y+1zCov+fPU/iTztX6QVVoM3
mOLz8Kd/k2bM4/Agd8AbQKriAi288hOROsm1b/gRx8CHvJwiBdG7EBn/BjLJo8cy
HGlVxnSCIv+2QSexNr97arcpDsGhBFmLly31jem/tzJG4GYAFQRbfKAELLLHEJg3
3egx4Zo0sdZAJ4H3Ym+07Jl06PDXlDEsn22LxlRIf1NnlK2eChenZ8q0XUcOAqxi
wDHkR6y5V9lO+vRc5qrOhahA+j17khr31GXpVHjfCcrftBaYurSxlNXfzKk8i3ir
q282UCVXVttRwCKO/BlSuZI09sCvK4txMahrb5ejGAEyJtcb0RDxbO849rAXI3Xq
aNpDT5gdeiQmAd/7GyZ/pBbYtQEpjai3qWRmBeVc/7jsAsHFDvngTZxghgd2g2tY
vTUP7GS6vbCnHEyzbmKaI7rWJFfSjEm9FVuvrHHc4tYJxY/M1OZG0yYLQ2zfwJOl
fiAP13cK11ESQYKGFVzQqwcHO3qVfMvVPajUYnxliV3t7qT9jqbjDWbBFqJrXvJT
vKxNSVLWHO0V3O6tcl6Hne5QsYY2hF9oUTYb8GO/u5SIvxwjgtQhO58YOU6Pl0Ta
HA9Q0IWCz7MEeHJ894s4zAa3I9OHZxIfzap9D4gYx2fNiJ+cLTLMRIpo2Pgq1IEb
dRVQlSEUrvtDQt/+lJC2YHFKkK6vLvE/rHM2SOALkA3EUCU3RHLVfk8fqo3M9h+N
S4eD3vNs6f3vOTJu1PtcR1nAzBTxbfgvJ8QvyPNN7qW/BpQD+CedvHXw0MALHeK9
3noZ+JtDoM1W/sbUDq9OR1xJUiVz7tJhFJzZJsqwYq4jMg8o10b03t3YSdzf+GqE
j9YjfOx2dSZDM8dGD3w/rli8qE0bpDXCeYs72x7WPhf2KtgnH9XDhfgan6jph7pK
bV8U7RfRTRyJNMKyHJB/3aCj/iL/UO7N0SnFxAR2ko1j6DDyP/tDxjg+FuWreVw5
LM8mTi1RWxYHEHvlxQTRhtCa0IjzTi+fL9EnnPAhJoziW61K+cizL8qk31ZLV5Dr
SsdHYeJ+usenxiDndA3WzZGvLwmtj1zqO2cjBBl2y1m3sgVBCpRs0wqa61AvG/u3
JRN/ND9X3RkAidNm/1Nhp9MTBBf9jdnFIEesKLoox4VsrpC4M+rMgpTNoEbKE59e
cjPEL5qF5emNvQdHRc9pMlBOg+7swcIojlfQRZgJ33r3agTidlWNHnm6auvWFeQe
PU804KudxAhI+tZYp6YAPRVgfjJ1crgYEQq5gPIm6p/j6NKDH1gC5af6UFukUDWc
jgQCHATsNLq3+qdAMHN/JrPF5b+ZjwH96wlHxaCDHcgm1ObovPF3TOX/ubNviA/v
SLcFcCl9NbpYcLPQUwmrrXSF77DLeNaIbibCsSqdhPqAiQwi1+KrA2klqob2eXA0
0a5x+KpxI5ONLmTVYF/k67Achd8bKPatsZEhWVT+cU/UcPyZvqnmpiJTKdr9tjH6
YQduY1xQ34ak6A88+bmu5av2mbq95bo3ZmHtjYWepYPFlsN/VV9CeLPqsD0u5C7u
i4hDml3mD49Glz0kRrBo4RLtpNUnP60eCThc/GJWvcjQ55hc8EgGAVol4ggcU7BD
SurvHuQ+/hQO6EdYhtHo9wO63HRXVHrwry1steLdB1ay0qykp66/bSmQDgCssmaU
J/45+cCrfL6xXOefxXgw5Zsz5NLfPgVyJXbaG+bHSiJp7agDDRZswu3t8EpPXKiF
pwaM1lNjmLHtCWDgj0oZc4+3wWlIK4Ca8SqOm6F/ctEJ2Jf8WR1cwtxduMKk4HpU
+cM3vbO/ljsSXGZFjiORd+XMhA7lRQnCQkdYlmsKYhg6wDiQ4LacVwix00eTwpny
f0K+8lekb6PMGqa5i9rWzbDp16q6LUsIp0LP+fPaR7TXFY6YfUKCX0U/QfTyqo1o
mluiFB6El7f8uEMDv8JYbOAnwyq97JBubzWt1DdbHrhOrWXP7vkS83JYH6LxUoLq
rgTW2mJqF/MYRyKMHQFwJlpEed6+Jr5FQv0x/pcRnDc4VUkWVx5BFiC9Uo/YA1Ka
mH5mzXkmrDGHreIRoWj/HQJiWa4u+4bdBBVaP6O0gd4Ey2XhZyaOlgy/Ht+8XAR9
lxU1Y2kyWihKOHpMjVT9NsEO9s6dHEAx8U+XePpLbcsR0M/FmzV+535sKPTcARpM
uz1nNhr+dcJpysrIFsVq9LwIeWd66VV1bHadz/Q0liIgoFSxAqbxxbjsHEvv2LHD
4PEUVSg4DEAfvj8pR1TsO5/OfutWnkLvrNNydKZEEnu7ltmYOx/5TSVA9vf8Ngto
IwO7i/zKR7QfMYfEvGZJKlp2UtOtBRm5zUqeraaA8a1YavVLOGS8mIytvwVZQO9b
xo594alR6Fsl/AcnfkeWR/ktBnKIpqNWs37Anslg58BloaizC7Fdxc1HE66EmF0P
J02oJsO+6uUoZZKliUBECePhRAybzVPtHJXXtdTdovh4m1shbiU8NsDANkTbiaQS
aUhCXZMQgWYVqUoyjK1bFJc4GRrZKOOYUIbqmRf+LDHJFTJrDErjHKs0v12IPc7b
VEXyYAJkMXXH+KV0Gos6pnAUxB1K6I5K09zhIKxGM2FRne1tbeq8FJ731TKB57Ve
qADNmjRHhXVizY1YafAG0t4zy4lTyGKP0hsv0xMtfFeblnm+ue3ufQLCb2ZiX+cz
CxsiNfgNZIBF0j7t+I9yr1yPUVGAY+Lh8SjbAKIxN07K3WfAPduMrbBWZwF3o/1Q
Kkmn2QZBYXtSb9o3qyQQZpy9YLpTKrR6AXhedXJsVJfgfCj7mY7eXD8zirl+ffIx
kWFVufHAzbeKG5o5hNrvXoNyratrZR6Hq3B82WxWCccBNHOmWSVND/Pt60UPaPcU
Ch1qSrR2npm1ugz/mI1KYb4h4GPP8y9OIFkDjcEIUSP2o4sglWD5688PfUGfdDqX
mKlDOOBCWcjbMq/t1+utgiyjO1Sk7uZ73ZM528zVy1kO2WHB7W0Heil380fj8V39
sROVcbTVs4ekobW3vfgpTpaxPMC8guHXXxd+kLPlLSjJe6uV5vjlYvZoKAu/NqOm
J6dm2pe9tnlzk78xL+GoZxYela3+6G8yZ25ffgk7iPMy1Tz5HwGw7uZ+jSfalNRE
x1pMIY4YotHrIIsnD8s/5iJj6ff1glR496gt4c9XD5vVZlfc5t9XU6o5GKXRPlIK
Jc5e3uUJQT0s/6HBFWP6KR68qGJsMf9wgB6ZzuSxijhe04Cpty1v+jtpDia38t6t
fk3kcr2FIqo88zLdEr5EU1atGR0zhI59yQhyCjH52jEW2UBOvHCmGx6KrSL1GEx3
dPeTihQRdNaAW286x6M95HyTN7juLI8PBFcIs2SCJwO07uf9oeDSgto8AaOQYcwh
mAg7StC04XyrsMV03lWmatX7dLCRSlU2ajlqJULVXTzKXWUTvKu60+jaxAGbB24z
XCQT3/+8PEVi8rrgnEzVy6O5VWtI1OhXEuUKcFCpTrQxx/a1EiQbZOzV0gf4w8Wg
FO8N5uh7+R5IEaKrvvDbSTwYL/xVOdhbOVYkhrf8VnplHyb6l8si70ZhDA2jmRhh
qbLvJyLF9RBvbewt9u7NCLUa195hGto1Bbvg5kZMggqLTx6V43pFHumQV3Uhdq9J
4EvIiVrUrRLhHnMujI0+CKJEliWbSUyHixfSiwKdn03u/5LVamNnylU5TJVhVde4
/vJryZ5jgLLK1ofv7Dd5vV9bOY1nXRsVeNBtEQrGSDBMyuR49eypVZOkaT3OB4Iv
CiiYqWnloRgusKVi89v58EvaenTrRiSclbOu33yoLJXX2v/ehuYTNrw8GfClkTY3
bvYKlgc905idDMepFYKji1fBi63FniEElufYXPc4ckhTyx5s6js2WMRC94CLx87H
zuyK6jIkeU3jF28CLdvJLetTiwBRpsbZmf+50X14gFHKRoWAXcZ88j2LhfkGoVRj
mKfqM+yb8yb4OQL92OfHBQHSN7mJb5ZbjJUBCX8YSPfhPwJZrEE7kAvgcf/TKj3x
U1WHbbRYpWk3olntegXYxDVBVENZOYAAHrNogcf4XuPlT0qt0WaltZlrj56xJFFO
VzmI8bzByiwmyrGG4dq9DZZijmGi8Pu+VpJFgOPHZP8CxNS7RgH/iFaVWMxwozKr
2sclUr/mlPKg0oIcFajxFVb7gbOyJzuxOUaN8GK6McwiXOS6bEyxTnfIzgwc1LwW
R5gYhCacSpkJ8gudrNkuvGlBFVfUI8AUhg5vK5/0z/R7Iu8k/MlHiqifNlji4fOf
4HJbkbk4EiCqLbYukFrw+pR48O6/mXQJXqSLclRzFl1WCgYf+XeWWinkQfdXVm3l
S4w5h/br1c9JuE79T2X0yoZ/MtEYkcy8Oxa48HwzWa2itMlDNyDU3p+/pKhNWhb1
MTdnvkMEzlu0KWam20tUVvgaV5lkSjHD6qbFFC5CvY8uV7nOugOR4ZOqEzcOvfZg
dcdpBYpe/r96cNfLQP69tXIqSw8X4Rxo2xOiB9kEcTMlPOtrenBJ84xAQZk2iFYS
OYfahv6fMh/RMfLQ65/zNVu0XeizVOlAhVNZHCeh4hhrjxwlDTKbwamri+AXxRzG
VJIZVecylCmqnRGJj348PjRX5JmNKt12CcD3/VQ2P2HLeAyKt6MPVnmG6miPWANx
zHtzcZFzfHcChpK7pK3UX8kZlYCS7E0YnF2nQHsWGyZBtVUo8UNU8fYr4zttps6R
PDebU3fDmuRQjrElVBZmQeOj1myv0vckHQwU5nqFQA9LjdojeU4y/uKhnP5edV/P
DpEdbeuInerJinW+/etMj8cUX+4oqSVuVrRgFETGVp0bcGLZW3n2aaVjxchZOCVh
GuUzCh4ilA5jw95raHc9q7W2TgAHHB1LghtgrcSvQ07uKVJ9spkYIm/gvNb7z2eY
OcZuQL8/lGGe+xjEa0Wh5U/xH3y0dt5OY33qZa4s+eatqek7WgmhoXbtbQX1uvvp
FhJ2i5oXqP9/WOZKxP1VIVExnT2Cq+JxfTNTH+lT1y5+50wjFg719/TuaAeXN5Xw
DljMhFo31pIfJw5+pF0SmnASZq4r8vfEncKsvnLkILbV0ruhW46NViaOsiIluWPx
iGbMjsgTU/Tj5zbC95BzFfZTymIXwD2Z+CiZeHz/gk/WhipevhAhjijRMQFBT8rN
vuA2bHF2olvGNyHAlsNOTYswybkYe7RLoKXFwdwpYFEji6GUykAnMIjyHUMWKcCq
H3G4WDls1XNw8rsWaXgjfbF2/+DV2tVAUaffY4uab287Rff81m7+/26awjplm8Hc
/LMs1C7jpG56ln9d1endhs0nggd4lHlUvR8I6v1qeLWAI5KGGaw1Q7Xa9ky+vvvY
yJiA8Et9VolamE9RUDMBghtYd0aaDbD7LayV7UZrW104VOPxOrFVyCRd8Bfpz3Sl
xyDJLDxAmtXhW+vvGU5B5/6N4yo+WNhcAKxssyoi6X/O5GXq9hg2oRWWS6aqgDcV
iU0xbChNdxOZsbNsincNy3vBVg2UrkvUHK/r6wQsrc+NfbeiCnTR1xsB9ZMw1Zu5
mRDRvOd2zC6qiJXu7ai3qU/u0WbRXsjIxbk1YJUy5fYmQjJZ3PF8kS2pF0BNSgCR
l4blqnbW2Tzz5vJbdRLyfHDjakj6H145XxI1J1Rj/TaDn7mEZTrd81XLBNLObf9u
O6jB4EZazA2WcnJDrr05k9xkjRFNIEnHL8AdzLEiEEj2J3MGZovs0ju+tQJbllOa
7HxqQa2d9HVAPZjCCAQuo54LGwPahrdVsS6itkS6/3wwfEMkVMoWTB1eNtPS5FRD
KMcWipNHbT/tqXxfJChvKNY2WO5VkensS//RWNq9tZLcdHl2gki01rbS4WkIeaks
fLWLa3Wmy8EDoFQs8npgoM7em3H2zDo2BaY4KMUyXkSqcuvGaY7pVMVgqnAT6VW+
fob9mK0XHsU5+iLrhFdXoQJonoDu4XJL25hm1DE3i3izahvoU68f2N6SeM3NADK4
rqIVxviqI59OfGJrF0ZnObndM/w1yno6k1+YcTKFs+WcSdQcMGDt1yy7rUX79O94
i+dW7uMBx6rZJvePHz9O7MHSd5/h3t/AsrMPekhN5JPnnMyzG1HLDT2PAJFLiDJq
XBpoIX/rSSsL4tjQlacchJJSdUtHh0FlOqX+ZgrsedEKdvQl5oTznpyILdx6oTR9
GbetVuUuthirdHO4uHH1+0mij7lxQ98WSjftQ26H3aU/gFFmQl8bwCTndifbFUHM
IDf4SU4o+SrrZydex0Ade13nB3S6S42RAxtU8GxQ4eghExTMKBYtXII5+MDpMqtH
xEZd0jxkBVCy2LkXfMSa4vBynNcLAP95FK99DnMnuqLg6iDapzhlTEu6locKMAvJ
zEcB6ZQD/vn6iU1dtCShsuSuuyR7nE7b6/fmD8+mOb3JGgans8zJWQBcmfr0gmy0
bI4gjIROaNQbnK/3XVOVCJsJxhHwQImYTNlhylQrUnQY8BaF8joJXd3FJGr8bNVi
KSdpb2DKHD+YX0UcIqaFhDxi1IpghCtAN5b9IaPriXbdpaVkptBD0HVczPYxaWiN
2vSqenQLvuygymGe9ztHF9Kl6oMGjVrLtXC4abBlvtLjs05SFGvGk55kxFXjlfEw
BpOnquCKx9Odes1ZIrwLQ2uyphCTavnWyvMZNexVr/ntP/0ffsmH5h2YUiORZk70
kRzxYggDgUJBsrUMoWH5gEGz3tmVQsN0Ung1PI3knIBL/F2kS857IQDk6dlp1SgB
cWe1wmDq98iFYcH5aTsFvKdicPKaJZcZE3Ogy+2LWelmqbIS9LfGig9dMLhCSQTS
+nMdIGAuaUKYMw/Zn41L79qUG8Wj1MaptYbt7tedY1SRkBAgN5h9n+1WMrEz2DYY
4Wjr1AVQioFU6SEP3/NMvclFTzXZdSfZ+PMmW7V8cmo/gT3hG7KIpUqsNsqK887j
FMeINndal2CraRzPZERoLfGlNEWm0xtrzyFazDkLvjodPe16xvZZUC5zdyb1hG3P
h4mzs2E5nYkmxbgsiW6pFR0dnZNs9/VnJsuL/f75mH52KowZFtLON/II+v+tHV4f
mb2lrp/Yw1Hu/NRAQLyc1F1tSYe/HqwZdvuOMK90DKIim7rrsEi1SBR4wQ2NWwZ8
uHmo0PQLVwz4lQe+lnzth9DrYkUQKG9oXj+VZctdCuI9oAF62MVEAQfHn4Sc0X3T
90Peo8VWLnHwlfb2opOBXbqOXsLIYkk/9+t39BvZRd9mve+fFYT2xPr07FuMcmjt
OU+q6T1fBU+Ih6by/4B0dzSP8X5+/2LMKiCuiGMydvW80rfAzfsGsChmVVlS64oY
AnGUh7VJnzQN4fUq0cHllWgFjrIzyls+uDev+44MIXQ6OrJ0NxrlHlLIkl8HXz+1
8q8U0wfsWdM4VDyjIyDCtCMJIQ83DKw4ZdqH0d+1jTSgK+BDEDl14AHTNOKMlemJ
D/ZSRmTVnGwUqs+Bxin6GThbcwF4D2c8/9Cmp+Ri6Vi/46+wngQg8M1SMxLLDQt2
xk3hcrFgdBhXK6wxHb+WEHmonH5hHC/gkCLCQ9aIFcIzzOTonWCuPffQQuPUv9nF
YViWMLt3nZas6IsgzyT7tBUc1gbZPjju7jtzfTWWV81n42g2cSawcqY0VVImKNyQ
bYCwfFYBgKDx/bleJGkyhDqlb4u+MYqFfKwJ7qOmfzMLpZEoRKW/ZI8ouMcKEa+3
/+sINSXHMxHvyNyjhVQ5b1oietvABLv7k378bLohm9wwK/rz+vWdwsO/9V9I9q2E
tixjo60GaLMLKzqEkBKFcDX5+Keya4eux6bJ3BufRXEXHTVkWseL+MYeQySyLFds
y71MXH8Itd/mF1rOklMV5/AaScgewZ3+PgUvwSHeBsNJJuXXEwrFfW1MxyKu5gcU
NjXFP7K2qOXyl5nq10XDKcyQFHAUb+VfwUFm2Hnf6ru/tE3ZqbbpNrMOO60GEDdY
EyEKwAkgRzWMrqDDE2HnihNEiWYyCc+y6n4wd2qdlxOCINElzKSBdSMeMAw8NyNp
4uLrkKG1uljoq8I3x4W8SMLidkp3JyXiqDYmkOjtnkCzCTGPkpN46bPijLgFb0mR
0i0/yk5EwbDd1AUau2CAbBGXUsu1fQujdF7BgC9MBB+D0pzp92s2LAjHWJn1D+BR
qfJ3OETrpAL1yr6WrOhYComTG99ZzL4qWqw2tHgSsy005tLXjamJk2xmG0F6jP4P
R22kIg/Z2rE6xsIDWRX5JnMDJFjv2hvKTvzbggXhkKmTIm8t65bZXK5O9BQ/HxYh
MjvQ8L19r/Byhlh/7sJW231gFALkUW/Y17nXVqZz6lHkRetHKC8rdVN8HI/CkBNM
jf8QxM9jvItPKKY7OYQ0hiS1G4LgdQE9ZFhHI1i29V6MHcENkYppnBdce0ENElDg
ka6jzLEShqoDnRPcfbRs/RUYEHk6zCt43p5W2mf3Sjbv0ILvcCjVVtHZloG7AjFO
Q/7QmLaP6H6aeToU96cy7qOO7GLwysSgug90FzMLZWZLepNKaG19hQsjRFl08PkT
O2JrUV/PZCXdz8p2fVDDcLyzfR7LozwB/IvgOGJVBpRpKIEbPH49q9t45cdnvhW4
ke71MZ7NL6FuVeR14OhmzEi4gw2HQUcnAWyk5LZdD3p9xaf0J1plydBmkT6HBKR9
SXcko5uj2P0lauhyMuT1alEwOz/Rg1u8ZIyWRlOiodK8N4cJ1ESkBIl03NN4w3G3
RRP1fkdTwgX1VfAM58zu6uEgWEXsj8HOU5RH2G1NbItjL3tp6NtNjd7fjW/FmRL0
oN2jXIgnL0AI/fWMhoav2fuqQZnyZsv2OuNSJ/RdXwhXk6xUMxlqICOCBr1NaKwB
rL86ngAH4RkaBDs1tEy46OQoicK3xcXyrH0euzA+o41OZgtd9uoYdC0Nnxy42pQr
c/6zz+cUyqgd8Nmvs17HaW4ggIbmFuqtMDzaihPhBqBu9/2eMCv2fW67+IgwlgVU
+4t4FSHecpPhwXdoU+c7ILRnmzDPvGxxoZZorVOqqxd82V5tZpVDj1xZQmqsdzLm
mbxSdbCAgNkKRodls9u9Kfp+26iaXPK5zRV+Of/PJ7nLPut8EVzBOWQb1hAIV5WY
UBo4unGSllQgHBr7aefQkwdJ2LyuEc8Kd1g+E1q+gnKGSiOSvWDNQqUoCsUirfMB
kOWFI0RLbl4oz758mz1yxaaBS0DDKRCjDGZrzBTepgy1NM4rSrVkxyQ5ZK/BOI0D
PaU/kq+zeL/qfDk96vrvCEghFXqbTLHbHmeTjuEJHc/7SgpQ/ivztYmAflqPS7nc
hvjrUCDH6h7pwWVAUOx1VFMGQ9V+W2yueSEl+ZsX8wGwq6/13mX2lyTNcJwoKC+M
oEZRKK+O1a54ZyQT7zAz1c/3D5oOubSG7HRR0cpcyVaC7ML4Z0kiYA/LE8Fg02cA
xvagXmtTj+DY6Vqdx2fIJae+wURJ9g7U0NIsON7mjr7LcB5OevWOMtl3rfxRuEg3
5exr8lLXPmSZVojjvMiewjJbx7POfHGDRqEXIP8yBkz7F+NWwXVx9nuBmoe5Yvw1
sTNop2V+5zJga3h73Y9Cp4fiOoM1uQeNQaWh+Dx8LNCqXgBTPoZROdd9fbaLPJm+
p7aEl0nUlMaaIOhXKYrVugtYmRXyis+IM/iCMhLJjwSdYuwWGqmN50WciV5mQSx7
s+7Q0BBJGvVkS/w4zL0DOqEof543nxWc/GAKkizO7nhWNfKX0P3qQNY6D4H2o9vH
gCCjJGkxRWUpzVQs+0pXOR2mgj3wRHtYUL7OfRXYfhBhWTVMaM699HC3lnbj/ioC
GAuJqWdjQqN9IZMi1phN/ZPIckcCxa+/3K/guLGP6Enxjgusfgxa1aqendJxJMBK
zmQYsM5/p4Niij6X0y/ecCBAecgJn4p/kw3LtNL5LvM4HqXDuegfRLdqshogeET9
xYZSo1Ve0+PmF87JoQhcVnPknl1ZxcD7ohXCQd88rfocvgqV4KjSSvBTtTQQO4Mw
sVCZ0UXXG8oLyl83RmI+vBbdIwS6m3Lne37SFQS1CYsF7R3pXXAtBFwbjrFQbnZI
/zLPuBNy6m98jtBJWuvDljuW6q6FwQjJJg1UpvZ96AaR2XuucLkQq/m0sGVqKMXL
MZWuMXkXFbhu9gW8IYfugepjWQcgnrVtejfByMDhr3LpGHD29P1Hdk949DvfDmz3
JOtvHqxtO1SbB4AERYyOfYG5rBt8/NYK6cuSP4zwY5DPtXgmVEkuxFSYr2PsFFCn
ZIhlH/IHQ8HUSqEg6G6OL45Go9eY7IkK2clQzpaqprWW7BdQnj30kENxNhzk/ye2
+zuJK0/Z0UoyEzlBOtAY19olPwEnvI2JykasOKFDak9FB0ywE5K2122xqVhaVYqj
9qB6sbxyjGPeJx7dq8ql6+foprRUWHBKOgwP4z1m6DZFXEZv/fx5bbdyOgxZ+ssI
YFtBHGOymjTSQI/dwlzQrFOiucdj08DvAhG0AAtNJYD4PshQTMLF8XvpWiYALXW3
m+NsdhmyFEBUnjBn3uBzC3Zg6TLHZdkj/UujRfKGYJXx82JtF/E17i8CiyFwRwlD
tKZeEwE/yTGga/8B2fl661yO9nquoZ2ILCoWK9Tou3ppeUa//T85IeAJjEiRu1Za
M9o1deB/5bzR+dfDKyF+EJHD0O7T+j55Skm6L+nkAAyEoXjWQC5mfDwsNAvrtjLj
7MbwDdj+HEjhukx8qHoWbNpOSWtAbB3nXtJAcW//2gK106gt4U1RvTmEDW29Dc9y
IRes0EX6jmNeYo+DkCHWlsLkuTuKqYsY4zjJLnj8HYPZSUNutT9tCKCTEVd99DXx
SI+ng9f6ivSRLkXuSMtNfq9khGZ40nnHpS8SXGIP/WKPIu6O8/Mi2djfSscY0ZdR
AjtbgZLszlJEcGo1622KJygO7GGDZe6psWojGNDPyrqZIZH1IjkVDlzExiOAU1aK
61yBQGPVw/JwqEepgYK1Tf91UfsqOvrvsCmikHdIwr7CpJIz1hC2fIdMB76MhPc2
iKn73L1vGwFJFD3rYHiTbwHm4F8koUIwU5YElmnRcxlL9mtIoYNaizP5nDyQq7ww
oC0Pox850ogPKDUUrTvTenIRtQu3FCxfYGRUMWCS/5H6UlFc6ljfm0NxT6yYs/LU
vKCc3FOb+/rh++G2Lx5fnaNFYylt3rOmBijGAesC+YLyO4Htn9VDzu5x9KRvUxDp
qFT3GljUTsCry+QcpMV0ZaLUXpWucjr7Gw79OZdgTDwdnaDb2DRGt/Shq9WFsoJM
6zhTX3VOp0D+CgWRgW/c+kX0ZcEcEviPt3NVLux7qMOimh92XBt7zzuYtmy664hc
GkBs3Am11rajSsKrUrOHx0N1wT6ZFGGLhTUSlzF2BrBapSe47CowkJk+0yfPaZYI
FMzBna6WXL0O1LHZvVwApZKiHpB53FsaQPZdMPPNBfOE2EQJQ1z2E0Vf08i1pa7M
NKxTgEG/Vi/y9/XF2ArV64HCABs5EaPjgOq7BJC1ClPdJsVCRiWHoi5TJtBYVKLt
m6d4BzToz27i+ghtoeruJ9Qy4/DBAPxm5XvJKqQtzIaD1sec3l3+JkqH17IqjDwR
HOWdCPJArPiIj47cq1Tv84ie4GgAQV1Cz6HgQumYDYyS9W/p2UQu9W5ULwNOVuDh
DtnWKOTN2Xap16x4X4cwIjZscJ7jLccvckO7eQ4n9rBJeloG5hgC8i/HFio27nGg
npvE80SAaiIEsWfjSSkI36fVp4Wdwi+DJoecKdT7duzE4p0Nj4qT2conEe8jUmno
0hmsHOpxHZeLaKKfRwsIlzgAZ/eUk2MNk+chkylfIFitxJdMuHg1Z42wmuYt+Vz/
866EweRSF188Eg6Ys7Lw9pmBWxZQ9ArfFXHYqYHbCdISvIV/s4wVVLCK3Em7pDw4
n+LRc99WL1UTOBoyeWtW0wL26uLgEAabdNOh8kCxvEVE5rd6DmeEtYJWwYWyOlIu
eo6DGOXj3auxE0ZecLiPQLMqvXiapq+kDmQrEwL7ogYbHE1iQ2UFiIgOFrulEVCf
wHaECxdSRWDhcySrtPv7JWYpIiunWFCcPgQTArUXN7478hhqKR8z1in1tO1gO48I
oYn49fo0wy846fKWooODbd5i+TgLAw6mvQSytvScU5ZUho/ZVnXDj0sbDaQKDiSJ
W/zkaAsO4MqwZtlR1n02Uo6n3H8Ik4vMFEaLKtCA8PoIEZbcxPUaFQTVwYDTGwu1
yGuY6aJbDBJHu0DPR1i4jqcllUgealA5LqGNfKC8vNwPsOW+2WyqIpL4k/nMIrxp
kEu6PFnrwtWO2LnQy2j4Xy0UhRqPSD48dXM7eNZ32L4WJcslNzXcNKMkO7yCLvZG
QMvD7r1KuXHvVegqC187tu7HwGzWW6nBFTXgRlfD1H/Kxd2+Rpfe8FQ/CJEQGsib
YnLK71OUnQXBNv+tyW0QrED9k9J0HM/zRVXCzoz8FsXaI6ln3oJkwd3V7bqF5HB6
Z6rdBoF7tgCpXOn2k4iIzOhNw98PIyucWpTXpY+Fq2OKx5BdezhSrfmIWPkbVvkl
eLy1VM9o3YkZ7VeJ/5s8YYthZjlFrJBKMhigOHKrweswN3p/n4U/LdThQEGBM9EN
NvpXScoZUNXH4VmowfJZSPhaLvLXZnWkdXM6SuWWyUUVOWipt+eKVeySc9Iq0geW
I90P3EzJDjc21flXJl7vVPQh5480OwlbQuLFEFN9MQG7/ZKBUpPOghOs9Tgt0Ozf
C7xcHkiLfl4jHSwDOJPJ1BCExy1DHnllPsOTxMwFZHgxTa0zFhyuP+t/1/+iOE+o
pjbD45SALZA72dJZ5l/HIc8BRlB+wnj3cUQHU+0VwvGlBxjNIyb1f2atdpgP7pup
e9cD8Aki7mR40LVb+F+sgROrzJsZm0jAuAfT8ZuEma/BvGrAIJUM8/GMw2dN+rR2
Y6ehF9rQKOtbEvpjcoaO2UErQZsr52ETHJGfEoa+gD34QQHOilC9sr63vYdVa1fj
SWy09RocgWcw/dEAyaWJwq7Mx6Bs8Res7gr8xWuHQvp6ONCGv/bS6zkMB+z9kjRj
IppCW0vUBChKKUEmMfmf52I0bvft0esfjc7JerhBthdhlbAV8g/V4iLgrXBnU5Zo
1Y2WbC0OJsrTgeLfH1Qx0jJVVgCBLc+vnzMhBXg116vOl8bhza/QKF2+yFifNqTb
4RTAqUrkY0kje4wItsRUobRxLWZqnPL5cbKtXoA64UH7GsI/VTXXP1d8ycC/0s9f
5kuv34wiGKkNGU41ueCFoHlSg7GRGBG77tUYHDgMXlTMB6kX7gp1akRMORDE3cd2
mw/+fnRL8Wp28IY+zJgB2XmaD6jWcQLUO2W05FSYb4pgDOahu+HNt7zp1mf/ttfP
1+73VGwotbCrwPoRjrmQGAvcbMc98QugVNpOzFiUErxw6yuXHg7qSCoOLIKuqcZb
menV66EqLuX+sAuJMwMm2ZdaTRlIxoXhdzY0qjVFPoF9Y3P75hSQdsdrLCXypwBx
LtLBHe6SeRoKcU8PxWVr6ZfQG2LpA9hrp6j3eLRNJIyKKNNPKKt3EqOWFd9VJ1Tq
9ABSziL1LZDSohHeCKC7ua7Xynwe8AS+wYQBtAQJCC/tTpJoLkt5piVog0nJJ99O
ocqcnpYk8E6cmY4YraG4xAcbq9rfZYrvHCxU+r2KlwJfXjcpq8UBjSNL5pFtgzUT
1z3ipL7y/4yMVc8ptlhRBPkaELAtgBhoillGgBRHFwpe9E+B+S9RjPOPQpEyT+CN
5iSFMNuNIvXsfcJz8KgzAvESR4s32S+0XR8YXaFXFmlejPre+yA/gCKawMYDnPwl
KloV2EgConS1EGJMXe4uH7H2mLOpNEGkttvAz4CJGg6ytFcJzOFSROz1JeLkPiHe
2XVr/eqqvyCsK5xGyz7sO/YkpnyOwvDSWw45KC/forBEtkVeu0I/Pj8GAJyqkG4I
9pon/D7GGB1KEvJSI3uUJbWGWf7bop3yT7+2YaDqAuF3UbKocCqi0e66glEPIL2H
H4UXQoZht70t33RYfRvPq31kqj2W6KRTcCX+sXQR2diXsT0emSgC2k8wgfGhzyam
YAg2TuQlZS/XD56xWmjZAXIRjYaNTiPZJC1cD9L02LjO6dGhswfnJ3t1isum/wdp
TEzLzDCa4nF1vlH0qDBeEaTiumi84SfaeHrSJ+GnvLQ69FjMr7iQIkGhFEVYej0P
NO/CIaEkatFMQ43DH8tOcdAZBBakaXEax89pt4m2KZWWxtV2nOHiqo/OytTtXbzu
L7eZ6secMhPY5lSK67Dale9yPKe39oZ6hpabEv8Ab7tnxDsa6hrrOPEcLtjmyrFP
FMbxXNgeHbQ4U7q1XNmUo7SxNjQV3jDGbxvzKgSfZaZcGb9wvpzPpc2qS1Wnhqnp
122iS87kNVEX2Jl4iYhZI7AmqGcPdxvjc20oR9SiZ8YFfFi9WeEiHHPA8VxsGcVT
izN/Ry3IqEAy4rIQvinPigwDbTi7Wy0wSku4BAbGQ27RmD2weALpK/4DCg8jhuxP
w6VDTIIJjj8bDT02jvnWFyRQU9DX/KMsL36GeIq7BL6i8+rOxQUi/oMbJWMwbtNH
AsFCwbQ8OHuuUt6QzFBfbVum1AnN0dk/LAyWFuOxWMEEhnVJSfrcneEazbvjExs9
BFJaAd27WyBBXqM+COZ9Z3Xcwj+z0GdUKsM8P1Fwfk0Xw8Jy+llHkv6BkICKemPF
K7mAH5EOZRyKGqle6EKnjJiJyBZjEJztybV4LtKONULmlthHhHHLYWC+OKbp8fKn
V6aUG/rClbyY4K/FvXnRwMibg8oK8qt5z7zyt3AoJe9Lokqs01nxO8FrS4W3BX/2
xIKNolcal3tATNeWo4w14LNiKk0ifZlBOeK+Bl70ZnKx9rvpGaFF/C11HZcxnqMC
mctkVLZWXFgN5H3eYam8ge+/XiU+xNILU6pj3Q9tg+bbgOBHhTLdWRGqwjCM3ayU
G4OqBxgrHHJwQc7vvAQfSkzOe8f7npfuy4yydpspSoAbZ+ZIPB+XH+pk5XFAUIAZ
g11McGbT5C+VrtGLF4buISIVq4H6a5FPRBOjyhYdHxPvGqfA2+KRkdcSzhtxGyaw
yr3VvBcQx+Aj4QMBdJNSdYtukbpSjtNlqgday6AEHwfbA2hnGv2wY5QDNZ3a00DN
OKIH4YdEbrufmSBp3b5AJDGtXUrn2RW/Mbl6ecbMUIO7hL+jukMsQ9miUYw0YHGD
lOOW2vxc4TYosNBXHln5/+zkwiDqd2Ewr2CfIKS6u+7i0TZzva80IzdUhYkuRVEf
6nOWX2RutEUyJyxMGonQkXSHTY2RTcun47IhqialM0Pa+9+OP3wtAGUAYS93e9nn
53Zy70l4krDhXRYDXVyXjLrGx+pc9whMbZYsjl1ZY+zZVQZEzFtGPlk6ARY2We7e
jyij7qoflZtS/UnChPowyAuKOtCKcejY2eh9T9H1KEO4iFLS5QWJAOauY1jvtLKI
pusHalok5npbKSvSmCz3ROMuHCzPTaluJUuBNA/FQL6e7wUrkm6etPCPHt0cYImA
ON4o0AulL6o9hHWZa4mxnYwrvwFaTDfezyYPRANv7HEnZbB4GvOpXonA92+AnpkG
rY78eAucI6yMsG7+78vUfzlQVXHyTwIajDooTnAPdT8bCR9hAtnsFludIsQ805oJ
g0//8DhzpTYl9oQEgYeU93bDsYYcdFrmW7eX0wLV+wa2XSZvRDcD9UDOGJ5xTCmT
1zdVP5V1vYmZw4JYF4y05T62xKdDP7JH/XdKLnfjeUjxeLYa1ZlluQ3TWgoQbcTI
9W2LO9M8J/gjme6JYVeTl/GKpHOwaSafpfezW63BUWp/gMHAwrx3viy5damqJ+eH
7JrDiiW0PKeklFowoUnLYkhNrqlurbIxGfxLUiWS+5PPIk9oD6b/V/IKeVTUwuVi
OJxyFeJVUJXS1B3y82x3aGGv6lccmBwucg/cVTjPB/EfIzsqgC/W6zj1uIDuRS9D
9tvO5AloY7eIGUXHFgO5FGN2/JajvVbhdT744KfM2VH+IDm5E1rvr8AGOHwRWNx6
jsq5L+VpJevRi4h3sYrgwsq1ZZG9mJBFm2a7LdPh28qyE2dXtaes4Bu83BbmH4/s
yXo32SPtWNkmRTorhqkatY+dlgHDNjHH/DyLgZLYlbvS1oMNPDDWIQqjhV8nnjtH
Ov9slSz/HDNmCNm4dCZDvZzpK58j4IF7qwlyvj+WUI64QErsYZClGo2azX7KXS8z
1WVJK19X8LFvecizVqDCU9vCYF8GZ/vJJqrx7IAd5r1Qoq6f83XDAwS1H57vkzea
3nJrukZ8558kbGg6oaaUy1GbTvhaKG+Sds0AUZxgdUNUAPnafJyZK+B4DTXrkp3d
0M+kf3DIsotc6E8OtUqey/N/cjL7bc3SOu2OSHa0UXNKrhFU0nd5xkLRaTamL5VJ
hg/b27BkRXjo3ifEMTZNxFbXH4bXe5dLs2wG0Yh2PeZzX6hc8gdgtVp6m7rF2l1a
E2fQdkt9tl+rPTLo7Q6B6iX4u3z9aQBpWJVvPxTGGNDuxOVleJ6gWQjj/Gc945WD
wiiw/ZAYjelC2f8T3mB1OzxXzTnr1NEZYnu/+2AMTUDUn4KP22KXzJFJ+JgfexUL
lWHglGDuv58m9SaxtsJn4Tml51lYqlmI/NOlii8dOGmKDW42lDEA7WZZAIQ6yn2x
GZmaZ1HJ6VB5OyEKY4eUuWoyXv1G9tjzAwRH3ty8AHpeIGsmieek5h0vL+aapwaF
jzCf17i9z/WKj04Il63ZBwQ2IRZFHnfrAOPUpPhSahlX2GHMdzu2aD/YZUrlpRF2
qn1bkC1vZTbUMFZ8rUjhj4EC3E0428myah2EqLEvrSgG1v2RVA6UHywC4lpjMbwx
xyJpnMwSooWBGTctk7ck7HqOrqdS4ipyMldIpi/MtsTZBZX9o/t8mocHvGed5DR6
ylFAH1yhoNR3AKyav48G+9OhlBxqNGKa7sHLVxQ0fnyK/slTCsk1qLGBU0Kju0UF
WPwWpyqPvhwkTs5PRmW11Cp3xyr6RmrdtUwoQMH4pYiYfUbqTXwM1XbzuIPH/Uio
305g+ZY+AZFreKi5kNDHMTC6g+iNYMoUAaNxXoEReMPQZuPQ4iF3GWuDPTV7+bHj
fyB7JAYGJXTRs2otyUtA/B/xyvim7MQv1/IgxpMlsp62c4Iq0d4MyTMUsqbiZ1i+
WNCKl+/lAyEmeyJMqW9pHs+wyTa2ikUVkwN3sfEdVr8lzPlRowu6gqy7rWeGX5cK
W99DtMRvhILTodusiI9hYWq5lo4oUnduNHeAJZImap4uZOoMX73pFDkL8i4insfE
aZH4eh6LfnrJwAvGAbD6hJRCMfOQ7CY4RqXVp79u9Rg5UIMF+FFBdYRHhGuPCCfQ
SErA/6Pu1cBVEE3Jl4vYyvEeof2jgwZGvgHi8htJrXn2v8Hd2FnkcxEyrOq6vDcO
uJ1Squ3scsz2whEhw893CFyijPTxgG0QVXMMGCHl2OsoNqyyFUunDVo0IdY6fDad
EIt8AiU6sWSk1oAwANhkW1SPzJ1+y93j5Z3RFJHFqCzvIM1gq2Xci6UE+5I51/Xl
4h1LSLpDovSgMErjHEmI5B7pX9jTA3EAh23C8IbJdH1thQRUt152aUWeLymUmGhW
3tsy42ZyKxct0AM10EZJLkWR4pnCT+FYV5xfxNV/c0kK99/+39j8DChgCPwwZuOW
nXgw7fD535o1Pyp4iVZwX+GO1TbSCALgd1lF959kjv0V+guBwzMrT1YyxtwjF2vf
XcbctenLUESi60zMK2U1FSbcqeVToYqVthSr8FOs+pfFMWy6He9sXwf/4yAN9FTl
IraSwbUq4P55OB/kSH8+YTpbLHKgtX/87JVOjyraESkTmizylMP/N+ZPhll87PIc
y6uvhfj6hVhfOfCyZaIU4WfLwctYMztMMDNbiF3mAe8agil2f2Jrt/yM0lXkdCQm
HlXloRzQyFXxiVf1WhBrZeUnyvvvWLjj8oVCskcrQxS6/j18a972BS9WwyDlkc0Z
gl60EMbu2Iq5TfxZVHfsPQ+NFSwCROB0Thl2t7RRNXRTVgPPHF82wKtGtawW6JHc
XLh/45OceSRgj84A7EW3lB+gUKpmbHEqCfgChYcS6cArn7AW1yXdAcByE6lYIOH4
3S/6mAtdu4c6+ZY19Gcmf3u8Bdyg5ZY7P75GuRLiTzRAxH4eRHcPFiJpyWH4SQBW
7alahdggb3JdUpAGu921hQMn8TXKf1wXF502YVv7I2nDV9ZUxvxDnljcv9h6Rxm8
p/zYo6FeY4w16/s7tlRolYZoZv61gdKLkzZ0hktFXv29Kxc313sN7M+yiZzNLxd3
zyll3u6zvMyxO58kyWaSSmLgjYDPmkUKB1nvW6y1wZE+Rk9Fo6lPjJqfmPOOtgre
xgN0BLQDLH7LzR3cEYAcjsfuA+NdO5qKJOrOlXeQfzXe2O/NsSJLlX6fbiBksPrg
hFI5wQw239uV17XnjPtvYZt7Qla6WmtRG5PcG5tYlSNoDq3PsSqxvALmthsKsSwh
X2QluqWyZbNg4gVyn9wzKB14jBMiKQMG9jBMH+NXPdxLbVuVR/dpYgJV0FqZjCf1
0O/We0z4TjG+Pa5u5UIZ/4srqUfpQO4Ehc5AY/xF+lOxVuz5I3ZMiFEmNSY+rkni
jnjlGuDDRYOeZzvdWawQSuFx8ZkKJJzL6b/xVmrQ7Qyug+0gJ+BeEe7C4hreMq6M
FD8k8+SxUqV0oT5kZE7WVyg5tgHpg4NEdDpxApasOlF2x8FkpaQQYlfaceBhVnpA
KkIda4wr+m/6mlcH1Nz+KlTxO2RgkHncKLF8cZyL4Vw1Eb11f/OgRV/jLz+QMJ0i
rFo2sLMNyHAPzyhrc5lwR89GhSYMrIZeILyHWQuirPAunBrEjQ/5O/x+nylUy/T/
k1h1vQMS8RrhoGcleuyuB00p/O0P2zHNVvgocscHNQwLNnp8r8iMn7aL/lHbVZ23
dxD+dLqT4iuDkUuWVLXpWZ1A3bO+OZPb5uq8du8mUrmFMbDqe5WXcHZWinyGzGpS
csCGNfEPkEKGSgeTonfsVnKnGCBk/mwhBaNbnyQS8adOQIeQoRrJi0tNB/vRgAwe
X/SkBaoK6IsrxerEYOHDIIRmw45VQBLZsL9cxaPn8PgE+VwpW7SnYbAsKkbts4GB
RvXrjopOb4ptE6Qt95DZJ1H8cAneHprrW5RSI48YbCnT+V4l5+N8kyT/zohi4yjd
cjqwrYfJjLHG3oy7xPDqnxcOKUW2P2V86Yfo5FjkJRLJ6sq4pA8TEePAn0D0tWcD
boCuS0ft1szaBuItgTzlZfNAEw2GBD9YbzPcx8OgqSCJVTB71DbxPP+YFvgKp91g
t2yY7ySXJK/N7YtfI7NwO1njGDmlciaXU5NdkP/HFTjY19PJqPPR1JFxYnAyjzNz
lLOd+AXYXbVm89D966S3bgKUcoInEAIN5jjcXfts8ctJ13yxlUWThTon8i5OXC8W
Xa3z1zKix0Vperatuh79mR0c7kcl7SzSbtpCfKZiQwTXkfD7tkZzf3IBSCVxDNWt
ry92S4vSvSbzKQMeyKvWkXpnbCzN+K/AZE6wyXUwl8Q/9MCINvYmR03UtYDAC7D2
ulqF9N11VVm8qkcaQ90wEqgLRh+uZ1XjZgefiYolUHhcy4ybHlDGNL4Oaw2bIrSw
T2dvnpRWr1RIyXPXgF7Pb5CVnHReaIxdis2RDGSG74AW0uomO7OZqOzmnBP+Pibd
0PxaU5EoVk+ssfc/fnalnOEA1BV2Y7Evnis57WcsaibGis/Oa8+FqdV4GNHC1+TK
KrzQxfgcz2VSe0Og+NRKwZGCNrvw3NE3YQfS9RRCFBBY2cTaIgGqIk5Dh0SGRPAb
GgmruPJj+JHVDK3I0qOk40qoibtzVDA0SB9xT27qnmRTeWjfJwSE9Lt/fMDvtMnn
1/3DKi6xIl3MIZNsWPUNKJh8DCbCQNqfLrjMJmqbmiNoWg9HvPGJaA+ZurZHglhi
+xH1yitEqdtdvAXPvvqPtRkOoK9xguVdq7zBjzD3X7yBV1e/qbyO1mFuj/Rjjmju
JYHgLEllG8rTF/XzZgMoTWwThEBr8lRMl4ykyHfkLH7SoZQ/H9Ss/oSQaxf0Vd/f
eLAgu97w4qPjG+UXRR7a8f46bU4xW8jQDhfC//uVtK3bykgIzTtw96nasHerj2pV
0Jx5bNi9tSEQZp6htQ9X5rV+ZuACgrhoFhQYFhkhRqc79qh+89k2V6EdZQc0z7oe
D1mQlV2xDI9UMUBsMPYRLXmYKoqF2YjSX4o8nTflbkkJ3mg9cCYKuuVzmTFOy06R
t6babjCEqVZfVXB5lw6fnWiX/BU2SSgYy5puFO/yBo2EbE/NUganK9uIQzVYH/1f
suxNxvr+A3QIYNW3dSMghxNuIM2eRdgvYgaZ3aYAQYo/O2lFVDKfbfRcpKEkaai3
47yEO0nhOr5vxuOsBVY36b1B6cQeovNX01JhSsLlouQVdmctMz57WeGN5l1cHB31
M+8jAR5CVzhdugRb3OLTC2sskFAhBzKEMRzkS0zhq3vPSFWX19oL1B5axqmUoFTc
YfweNzuwP5vWwwaESqFayZs12WfSTAKpeBozQU91uTW/hDqD7IWtfvgrwpy3YyuJ
aVo6sYLIqMyjx2MObztNACsI7mCvlZCEXfBB5ovRWiiOa/6hmrr+njIxfJGYDSKJ
NlroZFgyGYQtMQ3vNF4zH3chiVzJfo0YiZo5HOvwHp326VVoWgfv7AXSoBohhHRp
aLPAcSo+NBMlGjZ8+3a3GPVw8d1TsXJpTKyWDcbIw2FjU7QDdnsDYAR261XJo4lV
lErIvWjlkkJ7pizsWTBCDT9rt74qODBmguSLnD4cALlmYVw/zJA1+y4QhyP4Pe0s
W77MBoU7rBKaOl+IuDbXqmKli/CL4OFWyT3oSvcFuVP9PrTUopXGi5su3qq4AMzP
ia6eVs86GCKUqKiHplrB+Vamv6tB/98zbCDdPsWpDdkaPwmhMWXKiJiXv225SCAh
6s3flvXhN3kvmV9364rjkRetIcMmg744apvMwmHtKVCdaCKOyN0wTH+A1IxZN61d
oq3fdZrkPyw4zSKc4EknC1SnwrEe2G+JTCYk3qgRsGL0jdqZ/phSPzlBjCPGnv+a
vPBCw0UBXvCks44bmAOsG02k51gdQcrcrWpJU7SwZRhhKn1TKGAGxDo/NDNEIZ0L
HFaDjSpEwQrETaqBTwIlTGAoOzbBIxnPPlUmIcMRZ2512viSAkZgXMkwHE8BvZx2
6NAKdlHeZFvBVUa2ISmTiwH7/1VuFmteiEq93cALXDGDEakUXWcMqoOmy88A6SVT
t0/FhNIxcJt5CgWJwjPrGrJ96CbtdO+caXiTz53G4A32k/up/W3zSUxV7WvENrEc
Excwf7jz3JhSeuF8K4he9VrrAVWY13aTNF2qV7NGV5SxfV/F/DDKigOA64OrjWx/
OH6BgFH0BCKiTMRziGtzwB8pOkC6A57rNeHX+zy7Dxi+e438Nk6Fc2+7hetUiCqC
4P1LQpLxODk5WNRdpAhQeipWMTegcNgHeO9MbUV34Rzu45o8gqLWmI0gQ1qneoNs
gbOhkcw37VHiC8keiNVi6M3cuX5F6xGFtSxOPc/sk9+5b1VRGFKff3IrWUO9AbXJ
iBxv6c3N2sVnG4BkCg0wRv5OYlDDlOokmfTsRDx//jDlauqDY14GHdSMH68xBMjR
uvVYJ11kBg2IthD7Yvd7pSlsCjE+rRV8pYN+gKTQgmOhguNHZSTkeiepX2b5TOQB
C0E4SI1yXfmebNcRRbwYPCRCOm9LJSUozawcVWpSEp/4wkZNgDRJLHyxQuFJe4lh
Uz3FDlljrrx+TDGyW9EqAqkLQz4ozlSS8TTt+hAgbm0F3p9j6GJKGH6nSxiKR8Ss
L+M1IAjr5t6XAYPKY3NugsX7zMSAA3rpkoxG5YZUXEkukeDzgufCVzbjR06lJwN1
4jRPVqe8f2m91aHRoEqocLpqSpvnT3cMvcsAX/gujFkvIEmggXJSFGCPRO50eojd
M9mHZQ7tHvQ+jVxRWM5yTQhQVPTLgFaCH2MYWVQLRQGy3iu5/4E2yXDTmoLgpmZQ
EAKaf8nqL/02IakhWkKk4qYsZdhMIxbC8UHoyHuhqApKKUOaBp/FcJGSaGC/N3+V
TQzq4/oe9apFCvHFVvLJSG64DRmdbg24cqCgpPFRNpMIa//DvL/tMDowRVljimtN
qPEMDDsgKzG3+r28QzGRFLQnkDt9Ga5nP6t4dQZaWVNrOS6RIgh0X4/sAsZ9RMRd
FmY5XKx9Z1lw0Nm4WNe9joGKdcNV2gjvT6gmMdDMVanpyeLZO8BdNgoE+PO9mqUN
6MsN3XfP+zX0gexqLbflaV4nt3d3cIWV6n05erxQsF2vOmOhezz+d3uj4/We8Vry
`protect END_PROTECTED
