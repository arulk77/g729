`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIXvlQU04bpvugfhIGgj1DDnt3N8pCmsASMavnkXHT6t
uGy1IRLmPpFu1eOT/BE/a5UvvRCPbuzz/H7xCUMC6CguOJ5d0n0rXfRSHnx1iw4B
4QNCRY6TB/lW6DN50SuQddryV+1wGfSocw9pgGT4UtZ3ODgMqv/X6gX8LQUccmcs
wJ8Kuq26G+/Vircn9XbfmahCXjQztLSNZlnvqJJ5QTFdBU+CL15tuE/cZbrjWo5D
CKdjU03Lr5NE98rfbnJT7g7Qy8eFt/6KKwvxnrISu2Ineb7aKDuzW9vDB+zdq7eB
Sq//X8rXkBcnHNz277fwkw==
`protect END_PROTECTED
