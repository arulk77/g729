`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCPks2jIwjNNMG6c7I1vOWjw3TFpKDa8sfkhfxiObqCA
3sq6ZhsbsKk6NIiiGsBczXU5X/H2InfoMxiUgJzVLKPuhPOt9ro5MRpBNbbDAoU2
9AzBk9kwZYPeF3G/QgQaFlYV+uf6+Eoz0hL126tSOFK54Niar63tvZ6xWt8m+j6P
5YpREuE+IvYAEjmJkBbTiTD9BhkTfAkVnya7ehTgzFzsPTme5USgUEHwUJqwsA8d
IQqy9eVhFb5JlT3fypbwmQqxJTncall0nT5Oicg8mcez5p2TrZfG+Npd6DfT4RT4
KEbzw5D7iCRG8o67lZytuFskJ9dkQ+MoSYCBGJvb+x/w1xhnasXiYNf/lbkOm27n
DoBSVoZzRB6ZAtfXngap4lBgiw+8UAwyT3Hd1F+Q2+SjV8DkEbRoMBQRVjv29cF+
WkP1Lkc61gI0reyWG6UC8+6x0N6xb5JnxO9KraqQUPDZWIZzcbZD3FLTK/RE0qqM
OoXiAkdHXOnsD+Jg3uiItB42lfAe1JjzqCska74As+NfFmmH9MJPPLlhUytrOQfd
LXoByb4rVkBvLEP34r1Di5Z9UR5vneh9z+UP8o5tYa8R1UFtfdgPD7PoI8YMa3KF
eooQ7xMBddBhRTUuEkY7RMaL3W5VlNDg2A1pJmMH6+Nca0ZhN3Ua3OLJnwn4zMSl
dnuvv4K1eJyNsKTIDAYRZeqqPlZxXwxl9z12KjtCYudFrBNvOVwNmGB0mo73RaPZ
QDOzgFa4oRDUoYcszAO/I2f9L//8w5d0orwigkmWmk3h6vEGZu/Oq7FqXblPQPRG
`protect END_PROTECTED
