`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAnmE2oYN//ZSosq09SmrmUZcA7mamnLnc132w4h/HPH
wmyMpHeLTJHV50p9kX/SuWSHGCw1YTLlbhaGnxXrghT/dHWh3OnY+YP5uqQadJUw
KJRXhFkgo/zkBI+BpfbrHbI4qkpIHjs6rIcSBoqA9/rtCHfyI+XMsDU86uzIM5vq
`protect END_PROTECTED
