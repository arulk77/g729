`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
s9CfFsT/EoWPhMDJO3NixQCBHvjx4Wff7gozMrtJfEvt17X1sdpsfompXuI8paEv
uwUu9qE/W+YyCHpRBlHYu7PJiYci77NPCWqkmXpEjfIrweWo+zUXxWe0Yuofz09H
PRRG8MwoSBm9NfntrtmkjtIThzgCCRR/oPEnEMemo/d98ATY1fHUwZ7KcxNTm4TK
Jp5ukfl3a8ixANDfeuikNv5Mdqkfhbd/3LQLcCcSHhs7HP74Kp7CnSfiVqPRbf+p
uPb6PvTrdMigWS1gRp8yDxsnr9nMCbBTsL8mJqtTb0dbS0aUHJMJX6VGA/JUQZME
/1VRJsI9MUFjqdbwCOG6Uahgs76V/t5I80yxJoea5dP49g0RvpkEAdKG+UOJ8F/L
odNH2GL6QAuZ8K0ncdVvPAgWeRntNO4INS4DGEbg+TY/CUDWi9rcHm8xluW7qxxz
9VYIhRxCQqAQrSolLD50DXpqiddxK1Y/jkeeJ4zfLrBs4F8FE/VHYNLgFjLLv5kn
SQPLI91ghB1eqgNBOgBYeJHqqDBVZnO1XuVP8MSSVIrDw5wGFQ3p0fIDhWgyrF+t
Ed6hpgXyZ9vIurPxSLVpwKBAGChgQMLo/q8Fz0f00fFsZQa7zZmOy264DGD2FOzn
iEWcJMjMXxZ12U6q/mLnsqkXW2cbz/0uUolDUsroGclfAcnBRfqW8Kl8KuctG7SA
wWikWzjcfvw1M6NtZknqWrhmbX2TWnBM/cl/lGfBwAd2O2YKtNNSgIYUbFCgU12I
TvZW8QyjzuMs3ycLyD+nwS47s+wSEPV4Y8cfPcOe0OpU1NK7L1XBfT74Oo+hpY0r
ONuE7UUlHS3OKfl1ULltS+cjMk13lVb20Z5AKRxL2QsTqn/IidXjaSuiZTWI0gk0
TsqTs64+d22sFtuKMzwLwOMEZ0IqBQj/Yc2SlXQe5enPX5q0iQwzAj6kXRxbRv1V
NRsl3b7jrMamXas/RKbwmOK8i04r7T8RiCs1jQSNKKKJ+Lf4FKTd3dXueibjLInF
2piZdeoS7DWJxO5p9zwv9qyrSpqG7zqmjV+DtLcslF+cXg0VsQGFSc+xODG4EqY5
f7GXHtvQM6aIW+v+IfavKjLVZu11Ggw1OX8p45EOr9m3soKxce54IVwzZFhhIolw
EGKRvMSzeH8qIuR7aAReL0oaNPwJ47B8b6FLCcTeHmOKFvCJvZLwmuggJsP0ilun
U+028IUT9Ta1dpGUe8kSmnQ2R0whaH1CXOMsWxl8FSBOACA1mSTZaQmRPVLAQKO6
/WicUE037XGMOLixr2V76UIVW+EEwLS6VINae6VScuP203+mPbdDu+cNziEhgy9U
HmxfJQYJrD771sGSxoWQzDtvqC/f6o54yRO+r1DuYmFT6XRI6nIqoWfQhHk8xHvV
RV5PyE7pp+58Hvi95B096RrbPaJYXGoRllfk+AuiD+vTqESu/Twpl68Z8RxPLvvM
RsBP01SLao9B+3dZgwxscZFg73KDyo1tjesksqO4TLRd7zjaV2p1dlDIkAx8HLaY
4qeCJXHq7atbfOzoLG/mPutF5xUoo7gshpeAdG2KzqByn74NqVm1d2vco6T227Tf
hB9aeHhWXyc02mB9VXWgx71iTXRPk7o9vArh5nL5D4LXLmQEqbUENC4QkIX97rTS
7UUNmdvVeUvIit3IHNfj8NkVJWWDGkt+3qlXMx6Ragmj2wUPF6oNmm6U9+DaKAUZ
LwmNupTn1aJV8MZhhMEJoNKvDZF08LWUUKKqEHohqa9UZPjG4Gsu1EKwytJaxmCe
WWnMZ1Y1w26bMp3xltbMLoTK4+k1aiuaX7lpgs5Jb3ovpfJHcdpGP8eOtmPSL+rY
Ke/MA3jvLgSa1+i5ik/5HUpzJ9W5No7zXp5bUOeLt/0wumCFa+wYJ3kg4zEickgH
nN8YwrO3kKS6Yfms2K4yZAUnXakO9vJhJjl4Q5+X2ypidszZlxyGzfCwoh41YFDl
g+FldmmIm3UW2P5nwn28k2cl9MCrCSySiOUS2QcBd/YCTaVrqAIV6a46/iBU2SrD
OYqejmYRlUuT3M0oj2C18b1u/aHoTWClWjZcgqvuSlC7ZiBDSiZkld+GjtJNWgUQ
VRlAhqzx6tEPugdUYSgFJRGMyE3iuUjZcP2AYec344LXThJLZrBVPrWC2qyxF/Lq
gP12PVb8X0pvmfZ191looEF40+zUeAVLj7GEaz+U3g+E3KFDOq3DYHBxz/ITrg68
3zp0szYR69CzKEqFBfXIwop0rOBBy22K7iTyfscpItYw3XRM9wTbA5m4rJGYEvPZ
ImUsC+8bYaWvxKoYD9VBCgexxlCIVtYgx8piJjFHXEFjgEsPoUF8n+3ZzWflfOvX
ZYlfK+qVpEHzJ96qpbqxgVENtScB/JvjuRuYUEyUr5IsnQvxiE+sryjzbrmlrcGs
/LxoYJJNT/beiQbSTgFyinAuME/vFl1ev4fw/Hro2JXrFTgDdMmvGHI/PRvxw/Ud
oHsTg79QRgaisqGJl+Ar5YRHfenoT1515jIXa+0Ak7hShQDJkaa5KIkoY1oyWoXq
SHEFmwTYiWTrF6W4QDYm/j3EFbzcZ315O3zqmYzdomNUQjCX5/HqKdW1hRW04npQ
a+qNTF5tibYaNxi2R5BcBYBGjNoszgZQpxJKlD1wIhw/3yAIunQigj5GasmoPPOS
5z1lp/3aM1Wcl7lWyxb3fzkN/pUpATk3ar0BmHng2WsoVqVi8dgGQogXdJGyJFjR
ZOCwP1qr7kJ3sy457Zj4qCRk4HVabAQKQ2e7rPTl7zkCX5RXQ5AP3qWv7VFfwDMa
BcDma5X0ljk2QWr49lUxJ0ssw5ME5vkgdcbkvUXORGrLa7VxM9RkayhsFtdLxuDk
JR04XAFFmJoI1XfWCudQiRqcS+Q5YB5XEI892KpeDRSKg0nmVaeQZhDju4rLvkMQ
7NJw7LiXElF00i6DWmCJIGMamgaGKTrjEO/4Ugnld3IviGI9mRv5Ay5GQI/O0uea
RmgUOmTZL6GTa5neMaPtY5QNaRk5eof+wgYvORtVS4jnwU/csckaxxAekemTxudG
qtw3utTgsdN/KzbxJxHXA5A4h2M/EdrRg6D7CncCi79G4BAeBsY9UTv3SdYlhJhQ
+UNyKVpTQUc+0j43mbnojFzjVdASOE9kA3Vqh1gzNb+/DY0jNCeP1od9nUxIhhxx
iy+G/wr0CynsL1rbjC1b1DvEhnTBpDcgsxchCNGsLqey6BZ3TCwWOCU/swIr7HdL
GtsBVo8Em436UE0YfWSovigk4UK3lynRxurlufFtpybfpsReCGXA2P2HXBaeIBN1
uPO9ZKLTGzm2CUGjBas6uEeyGtxVo0JXDIc+oY1h0dDoSGxdHsjmvpdOKCEz0DSV
vDtXwrMVoWeJUDCrmDnSNBgMNwyCXOBLvNReD/yiYu6vOdra0g98KusEk3ygga2Q
dhcAtBfq8aUV4hTSQSbmyE7hpoxg8Hq0Xx1+jF30jj/1MLrt6PA/dwb/WuW9csG1
ZiW6Xebq/GiOtotHVUPMXcEoj26FSLrY1VWYVbWqm1BQxtDKCPLxAwnmFrozP9nN
cly23htTE6GFwZgm3Qjs71zwu4PhCIwka9GUhmpAd401GQygTbP7NnqE3Qmasqx4
k/E2LRNAQtR3fCelYjY2C01QQ13ZbOw3NlUu2uikYz02f+TlcuG8rryEGlmjkZna
ORSsIpXXjZ/aKlip5w5me4pe9NbD9VLGCedcptlzSUdVh43M0BMXlucmfJGBwFE+
z3q7IjgK2z1+MqPoHeIKkvgUCyTHHNFgSaQUJ0USaVvEvB3WL4V8m9uNHC/ZlLWv
+34ADo4bBZpTkmCqR37SWMzb9cB5rYMrCuGtR/0YRWaEkE2xYrxHS2GAObl/lZvP
wMA2Z61ID+6eQfu8clDuufbbk8nXL/2zMBPlPch5PlqcIK2WDa5Qp8uQzv0Dvxd6
ROUdjJ5va6n8+cU+eVE6mVUmzGOg1R9Pa9j1FpZfphfy1cM1IzDGkGODLGOckBsy
BKykGk1e+h4e1h6wkOC8M9i+RW/4Kks0iNz0Y8FydFazWA3m/yzWMUVf3QMlI6+t
gOUOITlSqatzrMJFln66j5QCobK/XKUmALhMU17m5MhFK6Ecfh19/5OJ6mRpf13U
ZFe3OSE93mUjj7o6SQ7IIKJ+5YUChexcPaD6jKms+uiIVBWZttl1DzwS5UtKXSjw
2QXuzgsFejQeF+LXafyTygALpt7N9RE5IqNTJr8SpbwrCPfhDCH8J5PMLHatdlDT
lpb4t2oarcdW2HCVpW2fn3eaJ+F3fL3liLj3dbmgTsgPleXaAdWpJnyU6xytriR6
tHe8tncvzKzv+vD45mnRBOrxewjqBzlmBn4i1Fqtw5XrR+2Qaoo35Qae8RqLWrWH
KzITTR5nkxNS0UUQ3fQuMY2UAeKsReEk7j26WqNDgtSeW//t52MV+I7kk3+vCTnx
giKg8I/F35kCa5nV/yy21xGtjYh9rK31k6dRCr0XrkTOIbzvGVMrlXGzrZi35n1B
Jvy5stopTEBH0TtXCE8vackGVcjarXj0ub55ioINvrmrWvx8Vd/XrJq6d2NQ+HAo
mdtn/KJB0x8SzuUfLm5dQFrKT+9cq3OFDI14vrZlExxV7ChfP5T0IEIeaHLWMWne
MEMavnRGsawQvgoj0n/tauFGMuS3umG2rcL0fw9GmeKBZgBGzMcbhmPSoLjaMT2r
uxydIegAqUeSYgkjvnfFo/ChMK/bdGeGIopEPLoL2uqvS+r/wnvkL2UYZPuRca03
RUHEqULQutz5hu0gUc8FsF/LK8LwLpuv4jmjbNbHGHNiVPMao29PKRBICuWJ4rdT
V+hnbE5KWv1nOTnjdlweVgy3Hp89kzn5HM0PWF6Pc8QH36VOlEYavaxPm+HY/FuR
oKUHbVrCrTVQ1FtJqxsradIc2AbWrWmDwJLWS5XEdSOC3xNQ2O8OdYfe+BlgIG5N
CmHRSLCXLscCibEVS0qkPc2d7eVMSXguPypoChyNpqFwavGvVCPZjF/IyY3qTvg1
SdWWx4QNKHBLSvePxvAK1oB7W8IfbNPXzYhYTvTSp41wWDMdQXl/FIdpFXcvkI87
fbDqQiSoh2Wiht2ezOhbbrbLKeRhZYb98+LD4kTCCGe+cdypGU4vOhG0im9HnxI+
JTg3SBxajVGd7pDblOrB4mfHU2VTzZ38dHor4LPAo9skN4WzlJhgqj2Immm/cflV
GMs6PuMoNwtKFSlhwSk8o3sHcXqaDWlNWUNriP5yf8kxDBxe+q3Z+vLSXzwHFlZ6
4KjZEID6V5RdV4S/ww9bO35f7U0yyRx693rcu1iSqHGhW61cDBPPImr+aG6vWBai
+X61bfQKFQ/ksaEwOTChNyNi0AhSVpznzASGPrktWOvVLauMyGwcemBOymvnDOOt
7Gc78sLVOV9rFET5S3ibPxdG3PQi8SWX20iBAxW9yz45ShE5XpVdPfvTl1el+23J
H8iAPv16B6DcmOdKWOfGQ3Dnlkb/Ys94UE2oLd2SzFROP7UBW5dLtJ5kzSt+alCN
tPN38hdABx6sMYHjmYKLmDkCojDerF7HiY+WOT/bgixbYXrD2LUuh8ZFuVWy03vB
jGmAIJbF4apqRW+CbVrPJdQVbj2THDUbwc4jJXEU7ZAZ9b6vL9kPMtHTs2d/M8Cb
Bllp0V27/AsS/CB2dSvaHj13Hzp99jAEp8CS0vBdwssLNrbStVhSJi3YMlHzJcTp
NAUFVxZybO+RmBoLtIVPEjVGYi2163b1YN/j0jrztp3yqJ7w84NayRLHPcWQq/Jb
TiTLCgWUscUm85PnOV9IKOQkVBlR4efqPsTFKXuEHrym66pcy6ez6Cyitz9q6PtZ
188pHKa6hYHSnYJf/qWBLVsLMLP6tqu9gnloq/yDd2CX9xNFFoPc08vEu50uUbq9
AwjxRAskI+97UT9ROm4LE+247x5sFtzIurg/aFlnbrcW7i/rttTEWJ9Pt4zWi36Y
U6pKEMApF3/tgxX7t4qaJpHOCWkvPeZ+DfDgL/NuUEf/EkcPisLWM9aZ763GuYxF
5jkBJjQNc3gdhdSmhg39ZoyWZR85ucnGCW7WPX/6rdZi22LqWIJNmX7WEploWN+F
UiKG39kHcJoTyMvaIa24Qra680bA8chTnLoG3fgzDR7IFEYGYr0alrLAgbsBx7Xg
PW0sOE1ZycbFgjBIgX7+A9q6qqC2Xrfd1ZV1ceYCceNMVTeIxAGDwDyXd28hiriD
2cQuiCI7ZRdBk8QQje0nX3q7Z+lIKeDcB91UaiYtc3XCHSPJ5BFtBSrDyJN7owFJ
reHAeEfO6sqhbIfHjVYc+Dh51cuiYGhfY4TNCqhQf74xjad4B4LfxQ4exkF6exKr
K09eutfLjTdQPftZ8aPftP+0HcDoCxb+5nuCRdhm60/ID22f/n6XIZ8j/dtgzEOn
0LCu7S0ksPoLfIO2ygGwCqAjCUku9qi2+uBkS6GR50urFksfNevcruv9D7jLuxwS
ssoP9EbTKnYINOZVindFkRqaRvE/sHJpqQN0QBRtKfJ/nb9XU2hwSuH10DHQJpWS
cv3pv+d/nMu3ot4q8k4KpoDpQ4FT/ij4HUQ30woiuYpDGH5FqC8tJYbLnkOZsFV2
cChzl8ADLWtWRrK7I18JpBRxZzLoX5mrOEiGYd86XKZaeGeHuAuYQjMLwvtxwGae
5K6m+IeWNLh/6vyir3QUeo33Lu7z9R/goBsd3WU8jatUfFae8uQR+0GgWOeuv6Uo
XtixSjUg9aflqMCl1WUDCX92FgdAetGJByfbS/ldMSb5nAbapf942TtAPJ5fBBj7
n++1xAb3Anj5KESzbjz/xOlie72gZk77zD/y8Q7Oz27uyYnI078OWGU8BAj0k4Bg
W0yv4Mzw72GlsB/YNyJWjh+xEH1TmUWir+jVpsQVvhmshksTBqjXYaPEFCgr/bWL
ytgrzPOm8vt0v2mhvjERikLE13YsjQ4ilESuPI0CK7FH443YCzo/8jcRBhAizuVh
5ovZw4bgCphX2KW6EhMB8XXt+E5G6qCPE9CNMw/CJEvpE6WWzUr7HCogbVobpzso
bHkPoAI3NUX1FXvZ4eguJVl25MCYrExRIYMQapyj1wEbWjIbbhUFrx9jxgi95NG+
FwqGiyEWSaDus91E/Nj+Fo2aZ6z7o4RGIbWuM4kWh4/oL/qUBFlkfItf+PSONeSq
/DZxfcgldc5T4P/ZE5BiNQUh5CKwLz6LpvVtQJxlbCLb7Q8WwkleR1GITskDexs+
TA5712TCD73OtiWFPuzVLmAOxT5g5sHYjlptEK9yReyetVGTbDHdaGdFiHnyeyCZ
DsTO1Rp0uRSuX/xszChil9F7wL1lz/fWRisquqS77v6bB6X9q1DkSm2rF6V54f/y
EwtWxyCoSCJYlIVD8s2SrtAd0DjqxYkmwKYH7H/A5/SVO2eqrPQOg1XpWE4hwK4G
y2+Fztd2NJpGei4T9cPCNzSIEecJW/yuosN+6RYyTVij16x/IMHr+U5rufbXYAHF
J1F0K6L5cgXVqiApBSABvcOB+Z1OCYqbF11ZxBE4QDfdtzHSjjSeCP0q/PnCO2An
Cf0KB/MPGyDKWzKznUs99uDODxYk3ufT95bD23VSumrxccbbgyN8fOPAAR9jdvC4
RfN0M7eaX9hWt3DM0R5mrmGvMXQJMfBI10B6oaiGOruRlDHai9Gceqxdi3x6N81q
fur5KYyZEXrFBPidc4EP4YViMc2XpcUBwC3gmJ1Fw2m5nEGNwSxmZIBJ8RFwnx6y
brwv4WD8FonoNbArMTAB7ORqR+bcGrULwejAqWePps3ySIj1CJ9o/mI3x7qGAS2X
9hGL+gUgnmEsvwCKK366bjZ3RphZIe/9sGkynOeGGrqkbLgO6bsWXkCg4ikwCCpv
sEISRnEVvQJFheE5m/iq7xGODMffpmkr0s7KxzATHEwvC+0bSB9axfcYAEWQEaDt
wm/Q9yAb2KbR/PTomvg2FYU2D5Of/p2CVn+3LuVcyENmuXkfygEOfFQRosSGyP11
BkLOFZ0iGjK7ROAxtRiF4BW1bxqF6cFqmzEmMRaiMyITU7KL0laBmoU2Z6ibu7C3
ThXLGz2aPvN7n8GI35uFnjtwfRGRGLNqqZfLYZk3V+AbCgpuuGqmUKxptnpaBk5k
9/eRmp4m2+/93/WMPz50DFSBY//NkS7IsFH5vubYAM43cbkHgdSK4t1rmZrk1VLo
sWi576ys4IIWZUpBsG9/BU6ey08YqwogXHfW3U/gDIvTvBTweZ+/W1U2/CWMzKt/
cJvlEiJlsua1iIVC8Qb+qkBpRE4g2wPP2FjnFQuX3sZ8v5+OwFtBqsAQ93SWtL1X
XI4Ew62Ks72q9z1Sg+hzoybSM4iAUf0xR/DztNKIUjSmGd4PsxpPoXUeF65QXPIl
fvCNs8V41zTkJC7DRNnW/TvLG2eqFTrRcuwVAMPJd9fpb3Ko0JuyB3T6ASdAFRVS
p4y0/c9LTJq8db8eeLVA7fgumd/UUGq2s6soAXUfNqo7XyBqVkSYOKzMztKCmE0Z
GeTDaUCXlCiLMefFhXJFkaqn/Rm4bYBypPS0b0pg/j60LHdqV0x7Ot/wrM9TSwqu
PcGVBtSfFtqoNVL4Bz4dXHYVnwUgEikYPpL8DLzdLNTT0JMFaPunub7HBkGHkyfz
MpSP0IJkIG5fkQcccq6F7lVUn91S/jfmlIF48dBtJPUxXM2LpUaF2qu38FuzLQun
1eltpkuyAZqY6cDcf4hh20MoiadFbfTLPuM2M0c9YgWLQg7rWu1/hs/hTxJCbys2
2liohmxMsIHxFKBuRLpZcXgGjoQ1eHObHJQ0mILOsK8LOJjRysygFeB6D/ugnKuf
cwU47Y1X80MabfIACeXQ44IljCI9dA/N1Y6wtxEbeLSaNSMQUG9F5/YjHFEiDqNl
JRSAI82vzkI0/5TkKjEmQZLGITNolYRriqH5eavdYmIsbfRsLN4259GSBN1DU1D0
oHsVhRl6xVpIsiQiyVsa5jX1l/fSN0yDhE6Ul4n7icnI6qREqu3gqBC9o2XiTFGE
vXhSH2/o06+y7nFwg23lI6L60e1CX3iVJie2PjGDQvhmM9ElWPmrEpmwK44gT70C
RrsjPi+an+Gm7EZ9t78ObXew5oLg3AxNwcLFpc+gQp3wpDtdur4lDh8rUOFa36Tw
gR7OZHDp8RzfpeNqqpXTVjz8vXn4Vmy1Jp7qXAmcB8Q4kVRbpTSxveU7p/exMIaE
XxRIzKNhpqXpqCc2wnFRYjRiP/nR+g84bO+xZjp1IP9hMQ1kYIjA/VbsMRDKi/dw
LjaSJ1AQbI8hriF7G1ZEUmkjcwEEU1ep+qS7YS/D00QnMHf3oZHxUpXgzuUPE9hG
/p9y1jJa5bnIinqTjfxtNrefZI+lYsprN262NfQ8AZv2WrfzdYlXSVlpEV0ECKKW
jwhtynd55CArbvjWzReCGql+9EWBlJJKJBMGeAauhOKKx0YqPteGMuEHW9MIEzJO
oUsCTwPudHodWzZUPnMDnbJemvi7Ko7Lkgv1/hsE38gBeEQhQzgv+ifTvYpRmDqe
lkVMi2GN0UGo8oo2JUY0Ks9gtP53KAOqk/2b7jrJH4xDDhW2HVj8BNvUFrUGwdpr
BMzXzvThY2x9VEiNN6/g3MJRKiMfXhNfzNjdHnjS3aqPHlxPrP1v/p3xwF98o9gl
aYD/SLftssqEIpJ4aXXDIukaEMhfFoXIORsAVvkb9LYAqg7Lx8NstMCObfBuATFE
lKM3qHyIcNMVrarepPYUb1BXhRBQhUIK24CJvz193N/msvzf6hhG0K78Qn3iMfye
+4UpymcKHSmF4UEk9c3PsT73WIPVn+uihgdaAGHrQenZYSD9p+ec7ChyQRRk/PwF
sem/UjwNbCrrDfxpfDeAOelDDwX/+xlwTAgxjusKRHjgC4zLKuzOhwooGESHtpnO
NmLl72o8hmGZ1fxAIroj+qADxAm22K5TJ5NaOKiBhhgg7TbKmp11Xtpf+SWsB6AF
wRc4KvFoxaCClR7w25o5i/cW6n+yi3Uegtq1Y7pus2KoAn7Vl3wdlLWWl3+iR7+4
iugnAcJWtLo7p4C/ag00qMDO++erH+H2TQUwxrlUZ0MFEZ1yngd9dy6UgLor5+Le
aNe/BUFtYvKFG0NXp5EWo4z1Ce+Ze8Er+NkS8JEOch0sw8+MGIBek/mDfI0rAuXG
IVDbpAkTc6BsrNoqcD/cVwSaatTVSrbIunbSgq+tAB4SKMeybuJJByA5sNZsg81p
R9Sf0Q2P15548K7ouJutH+MpAI1mi3E4rLFFc6YvOUOn1yfHJ0PPwKrmygfwtnJ9
mQ08x6hiAHqB1aDUyWSkjOI7ZZB8UYzH6qTxFgq+H89WrKZ245sIqZ6ScoxdnJ2o
gad7N69yDkOmfKiLTin5Wj87wM8oa42SLwi3umoFM/AIdRvWsw1KoAMNfEcNc9mo
LjlFrWHxdSZ57A4bgqXHJ+EYdDOnCUUpRztU4IeB3ccjVaUP0loKxVka4Y+9TsHH
NopI4fhkLSNPYGYOkTPx8HsHNyBvy0d9p3Ep6s8ItUnKk0LAxrQ5oXn5bDq4IZ4W
9zN2l+qlTKsrNIhh+SFu48GL+YTYffujrxBQE+diNtD+EPlR6Dl0NO41zLW+6VZB
r46HlC2QXMBHpBrxDg2xXf/FLeZfZ9qdEm6WA61isIdkwl6Qc0kKMstWgt3l5BCO
LXDQb6ARWDOypMOcmhucnWEXZyKHywhLQYjxCqYEgZ+SES5MVWhf7xAlvsKbzZ2A
CjjPW8sgfktNWbwlUt8R7TvjJpzdz5w1IOht22MVE3A82n5oR/m/n7gF2ebqykoY
GpM9OYVLy9JRNR9n/ShDTYsByrKRf26r1frQStPFgitC7qv7qItmOrLr8xlRILH1
qdGzjNFkmCfmtiUgog+/Igw6FfcU61o6F7fLds4vrWvQY4fG0UB3dgf2Eq68yI0c
pH8uJEkXfHtSAJVotUTuyH+jI3u35zpaPIk4b7Ht0zhfwdVi2EGmXaNIWsxmv64D
CovPJEzgzLgdvFpYIRHCrJEYmh4UyUXOrSbQtBYqGvgaCzpaLiw1Ph3f19xlO0ne
d1pcDPkUL4/T232Gs24pU+GCawYL0hPXv8iWHdufeT3N24+IeZPTnMXSUgB3nrDe
JXzYeEqSe/2QkjgKsvgoOGi98VyuIPEPt7eFs7TZeO8l+m/bzCZ3lKnowe6wKG4x
4spyyEZCFjYgawesSkF7ISuGGeQ8lZfjx4eTWyQytYz0slzT6ak+kMavURU5XgXD
1/xs/KKClEJqOfbQMTqinRaeF6CueD+S48ktRwk1nbVmQDjv9ujZj0a9jX1Zpfrv
5glYDFtau+cronrzWae+oxmF4p8rwJ+e75xrNBzH0laTQr/bP9WT9NX7Eaywz7P/
lwkx2WYSUfuy4JHuM8iLZ6Uz1fmtOEh86IMlLXntmGIZp/O8zrruYU2UeY3lg70G
neLvJb65XdAz0jr2iJSBReduYy/BaxB1BXHpv4NQm9fF++K5JH9bL5tLK01lokyR
26i/LQuzVrrCQsQj8aoLZ0m1/Y6cODijrEsYFiiqUa88zZE6mqLRJLmPYhtp6yUb
935UgGi2X4nOxaiXhZJsEWq5ndCNTEtw16WZv9qz0NoFaKLC8uKB78pyxRN94msW
D8LQE+YwFoW90A9EkugtajYsamA7XtH6ij9pBwcnRRBHPd/BEv/VTV71+Ge6xFtX
RMi3xxNwt/NK3PrdrHhnN2oL5UINrSm3rAb9+faPo1v486Oa5TiXvz/uFOK8X9lf
Lr1Eg9JOw3ni6ItvWJNQY5+x9ZX25PuohTDmky31CeMSJcCPcPdUN/eViaUx2i7w
/jfkYwrpR5yYjk0w2o8UoO2UcAZC2JkoyyhK+O2Sjo5D8JX/N2InXv/gSUv+fkdP
Z4Kxi2mxjSYAO/euApL2gzKec5l+ufM3Yzso+ybrvxXFUTjrFxQrMn+JjQoHDLQB
4mJTBc0TwB64+cSuAAWS1yGCj0OhgqoL0PCA5xPm7jScAXD3suzqvlDAoftHCVdk
B0fewBz7v6NJSYrbuRjnFflO0SZr8HfZ5X3DpjgayJyc+/bL68/diUe+elJY8xJM
dBQ5itftCoGfw+xaZX4Ab9a0dXW9zvJNw0TLWy5vsCjuTKPjguxri9S5n3B349wR
aqOeNsdatSG/D/jJjx/KOmjO2GyE4/gWBAkyvG1B6dNI+V9ZjQ5oE54Awavwwgq/
IwWqddFspt3NIUT+NuLw2J70KifmcF159LWfbOsE0qKzWOsgG6ZtDXs6BOyUjpZn
smOv9PJ0/npUDBlSmSTbtyePS6tag0aGFilkXQS43bJUDabHBSsDe6C+0iPhvULi
MyaI1lWEp0Pozi9qKysPF5L1ij+aBh5iBM2TyfXd77KCUQYez7tzmW0lXGj4AFPa
4FdQuaY5zSHFT0gweHjTxyRfdjaPGthcswj+ES9r5UtMzjK3VfdQm4tujQyxXjcO
QNTP6v521CuE3s+tpXBTO899CaATfqYLhTMtld60IXAjXztn48dnnoxA/J6CYvPM
AKopse/Iw6YxtEMc8kl96HENOVjhAtPljZ04F9H93APMcI68nZ6qRWDsnE8P8LiE
tt5o+bUAuVMKATvOPyTs5WKz4JhNa2k28v682lGb9m4fR2pQVJ6Ff4Fo9LJ0ipPa
86ZxavVQLl63kehNH6WeOLpnAE63xHPIfCw/rSJEqGutpa4Dv09cRqyylpF6qDf3
keM4tRog40M/1M9D0oL9LwoZJJiqM1+LOhOLORBAa7FxyiBGNVt3TUYFoMnczpaT
sf1MLMCOQL6vEcVJ2+tykqeD/rkAfeUvaqVpPCPwFBgX+5Dihey7k8Jye4UKRLSc
2eXTrmm3X5B0wjxtdPnCLxa8aHmk6mS2jbSIgcx/mZd69X4tFQ16ev1iI52ysUQD
uxg82Y/NwVtOGzrE+o3xXvqbspi9ynkBrp67VXUYEiky2XJNaASCul/eB/wVXEun
9iffzBJmr7wEZzFPAmp5nMa/s+TLzJfJHpWy/JbQFeJZYib1g68gIxJh7t8ZiuFw
CHcAQekhjIRDeoT1MOgctSL9YUbr7UavyFJJnLiS8/pw8FD71b7w9lw5WXFrdI7C
/M3RQVbTgqS5EB4Z7qnR8bZ4DpwSab9yNl+3GZ8InTuQD4vNO8LvUoBSrgL7d0HM
X92i9Mz9lFQql9CU/cpaJZWGVdcvnYVtBGIrSEsypgzjvAkvWcpMBqywFivS/cm/
SzAS4A1Th+K33+CcU1g2Tp15HS5GX9b+l6U/MW92X651htOtvn8TUpt6VlSUanU8
uUfAqCltzAUWxlpQPHB2ItokNu+2iErAKy/bkiF36ENu2xvwVSE3DFEBOhzOrFLb
J9DnnYJS2UwZ/mYwtIj3pEmgHUa5rNOaEvddec8ou0BfOlXDhGMKx7xBqUCt3X2w
a8N9V7Jd28NtErLnb70OX06nzlEX/23R/TEMwS36fmNlMak7cOl8bQArwhOemKkE
2SWR6nNj/fFOt27Ld8DRyO3XssO+E17Aooy6fyRn/u/J7zwi3WtKrqcnNoY3sgQw
BF+R0P//SFlHU5XDd4yJqLn/h9No7bzMfRmhEkOJNLFcrCw8EwCpDBaT/6hiXUbZ
ef2AX4Go+2Vz5eojyBrU0gpcyEzrrOC88Kah0wSH7iw99Jh9aXLgEv0lvuP8EWS2
vBkJWqNIZrmlBxy0f5IxhEV5o8ioF1q3E3Ll6NLeSH2OiL3GAfaB3yrYIdJS8Vil
chv2YMKRra4zSw3+1PLT81u50DczHKesbeqWG+HpbV9ANddPlsCImxPJ0C7K51hF
P6iMoJLrhZHYds9Z9CP6gHLziolZ22HAPofEKQzQnlhdP0UucrmBckZAWiBkCczT
HaOURXQlvB0eyXYxSj/SCG+ScQmX/oG4dWpkKrt2dGEdX7w4pNMC6OMs91jCGH/A
cDNsBxmQ413L++nAlm0hA/eseRNrIQUmSVdL7cTwGE1ZZ+SDrLE0nzRDbckGo8KK
kF2VhBYlQK66+dPw37jFv9zy7xO0K0/6yeXO5Yp+t+FmPv+m1wystKMGili/wPXA
zFsU+rDYG8hgG80T8TrQOsdihGRH7wXiVswF3bRDOnaaQWuLwd7VS1WNfmjQ0Cay
X+QI98TI1vXMEQvktqfjYGzyXt/z4RIRaNcx9c15zNje3HToKgLLsdr+92zKRIg2
ZLoRoAAwuDfOk4iFkcBX/YKLIvOtHDFRy56roM1TkbkPhn+QfLOeY8adgBjV3B6O
HGK7yC3fWLrecmunJy2frHjrdTbXjoq1ifXeyqrmgRwuQ9zzZByLQ27i5oM3buuL
vQ7xbI73kQViqVN7q2BpcTjB6d3ax8OX38f4SvwmQQbt7X7YySmZZfenzcvhRhP2
DwmHbrrxFeOcnuyg4L2E19X/JbgszEPQka0YdGZL7qBprloenK0DVHmYGFxNAS9e
ZD/pWZ2mTX0ui0UhVeIJYC5aOpyyT9PmbFwXdThjM3qkoGYgK8iD89wsju1po4wQ
xuZy3y4TfZL4Mr0g+bu78bC+yTHb1DEJ+zELpQfLVZqOwTQCdpMxmfJJgmHQVhyL
UaGI0uuDUqFNLaEZYHRGKvGA6RMglSWPbOj+i7AjwPkMjQrHF0Yox0CtGiP5bgYN
LTy56g86f4q9z6OWO7OEdc5rfnPsmt/FEfXBA8Lv5aMVZ6Djm+fCGz9u4XK6lg30
TMAJdJsTgalvPNyXPwPCtyWiavDoWSQFe7M/V/vUBTdieYj6cvZp7spA+ZKLHRoi
RGBnJ05P5wVXAwRauhpzsaHDWaVvRsHeueQksa/B5k287iw7B3r4tGcv10OZObIu
VVg6uwW1GK2l1wuNjcDUWnP7q2RK6SlOgGRX16dm4ldU1Gi5ccBwCGsKUd4fO/ei
HJCAzKwygeRynhUsfjN4Xc44OvN0qxCcPkfed9/4iEcs6Oh49BpF/oMMkx4kVFPX
Jb45UuL1ZLWfIQcwsD+LhWZ4aaHvHoRtmgm2JrirquWJsHHw+mWrbnhZjL3HGEQk
r9MngHkc8wooDgSG2tuLUXAp4MWz52plfJEQ60Cg6IayjP74ar3ewWJA/Cd1wNSn
GZePAsNoowD95OPAXZpTqzn984fBUElBa/nXIwYKMJKeI1mFxPAn93aBPoXM7OnU
D2JJldbpgj9D2Et1NAIt0LbIpj9tPuRoioRONjbT7ZqgVQDct4M4lP3+Keyt5Xjw
SxRzJi2GaGB3UpWBPOgocQsjNqT41MyJRbpiruf99cQlT1pTLKBLcRdE8+++k7gY
JyZzFJm/H5EiXeZTZzqAoaNymVBzCUxcQA9gQ1JkC3bs2ZcGW5gGpMsuYcaiXZs7
ELk9bD5knrAb99ixljMuk5p/QJvd8VF22DKG5a0fQBhv5ByEhNE5d55rgPb3YlKw
mx+Pn/XbumuzjAngpqG7CLQQJpseClrKIiJQkuZ4CGk6APCkpLNCd4sL5LPEpEBm
rG+NWLcxyFcu1QQnfeDBiJm9N5Ok2aPhQrRHIdbP/Zq+rHxJVNU34HCO3zT+p5Y0
mV+2UhR3WJUVuOmk4VwfOZm790jIZW3kGmSmUr9Ljjv3NiNHZHoGZUvT9RL5AgDq
aUrDpoDTyiHCUbYPjf126vy17tPU5jyxsAiOnHfuXrXuOvQK0fjuQhlXpsdjmN4v
t5uyOFoJI/TBhlUGwB1hf3ExKK3Py1pb7LcmcNxxZITNjbv498F2JGWzntHChVXl
EGIkl8eIs7fQtZg9NFdo66rkHPXh9x8u1m1hAidiGOzChKEAQDVwJMV9zaSx6T0R
OURDNsYakNEa0rbKnb4dvXI73Te5oMSzusHmgLPZFC/NFQER9Kmp10496aXWea5x
7ABcl3PUPv5jWL5e/odvFTctakbohZUhp0XpdkqMLdOzbhOTtwpy48M8UUG532Wp
O1OuIQ4rKPmbWhIsOz1Ao8+Jr/qsdNAn6qnmJ/PHqR2zOsHlo6OyPcsO5DUyXywh
4NzoPZwQ6sSCX2rvjoYl3+Z6G18r5et/fhVnYBoD3KatXCpjfWKh5NP8rCkL7YPS
STfrLNpjtRcG2HvX/XZRfX+3O9t6sUf3iqe6cbIz6NXp2kE6MKQfLg5lhlBub6I2
aKSPOxf1co/WOzWKUgMqiENT6VcflZzlHOHJFO3mb00ABgtHSEeW7k/ilAi/VZUH
KTyhXY5IzjKy8/3Z9FT3ywKiu0ZuCvrvuwIIIz1QI0SOFmJ9e+LGUEfWUEiH0Ayh
ZQkrdDjmwXcUhgCSFjICCNH3i1XIj7Otze4Liu7RKDDsGsKi/AJTtK6XOeI8F/6W
7s8mg8UbhmKTzsKarshYwIw8UcxnbsXmSWO48TgAoeNUMeS0Zok86FW1RkJWdd92
6cUk0FCZXyjQqXhkGXuxzWBciSqw2wKvU8ad6QV2ehG9zp3QlWZIYeAYGqyovEy4
zrZEOiUnRmvKF7bH5FLGJ5O4dfnQh6zWyyqVByR3DiFhW0DRwuj2C4C8ZC3ul/cs
EPuYwmhn9I/9R8hibf1UIDSj5MdJxJWuVgEn8L89zzowpnTjqEOqGH6AHuPbJH8j
0Yh8ixyLoiilFeZtfY3Zc6WSAv5+Tn0T7OFh501fKog00eiBtBnz5W280HBXCKeh
LyFv2vqvFjWNrWxhkFw6prLUpmbA3DHic+vV51Fy4CCRP9ZGnzko/Ke2V3pkmJKp
oC44hHwej5THyCp7DbrbZkrgqbZCnV+s3sAXlTlaAcgbhZCj/YlomlxMtK+3ylqq
WyO5/dINzbym6ZneivovImPZIHt3Rs5UEANa1eLGC+wn7y8pgAcg8WJTml34sIwB
iu5SHer2fHte2YBVch+1QmlaUM82/LU+sUiubBICLe7raT4kMwaRkEwlB+lKKFn/
lSWcjR38T7lYpHbxwTrywJ9foa7lGHCmeCFkxUKq7mokRMpncqUhrZyF4HVZqAzo
q3b8PPkI77/KPG190kGYspX2PERiKjwP0n59jd744ouv3o3xmg2/8uidYTI50zv2
putq6FYQTkGpPi/sOoFO9dnNRscuYz3QWA384QeSVQrRjWI6jcUleLgnh74KbUf4
qZNgagK1RWKNo1lA2sI7xLf2NSrN03jho//VV0aVcOxo1OiDGrht9jRHQs2SdoFB
xuNWY7zo6tpf882TFQzNsW0sLfE9nufhvFJuAIBf5Xks6ix5c4z+fldLUFqRrDzm
JleObW5M4uLoqjo/D28xYwouaXoVJkV15aHOjzj/5A7xs14R3Xf22nTyfz5GGLrC
T6GHIyvwJXJkHQQMfqhPBOsPzcZXwijnuzUz8echJ/RtFTtyTNARYDRECYJspJ8T
9HjuXDxXTCuwdx4BtiYrYHmShMcpIvuZtykHR0fcJ6NQZ0lemqF+/dZRzn+NkzTj
sV6OcMPmtiaN1cV7p1+AMkytPvLiwVr82GZJTUT87ROhk7MQpM3sCqhaPS3EqQja
jgTAUqLJz2mA3PcPk2qDgV78+1WEVMbG8FBhYbeor7hhjSsf86lkbESWO27EiQrk
2IHGMIVc3E8+6MUy5b88iT93S2qIPRzTDSh1w4G3QFcFRXoxpcWMUkNtIpsLs7IZ
iFfh+bVgR5rQYb9HPFMq/xVMdRHlMZ1seIbKaWZf7Z9NuEZ2m8BnNOvLl5BnGzpG
HQBQ5eE0tjGFtMvNfnSo8gw5E716Rz9xRKsckep4YJXVTWGgDcz+arJTUemOKg/v
EaCYK1INtwAu+J0nsn8TP3IUeMYSDounj4COgdLfgLe/JcSHd3ECl5mCeKG1ylS/
7aBtaEbdEJfTZaEYJArnrSXxjiSizrxXWevs9yesDUNtpfP3xHdOjDdT3zBg5NiN
ac1XPdij+H6eob+G+SbkJMb+JVwt+y5UqnhfdKnaSrfqZMx7rXrfcvoCuX5vyUmP
`protect END_PROTECTED
