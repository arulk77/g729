`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGCqAWcU4H3H6qDCDAKm+OPFugaC/mJXa8gKGEfemq/A
MaKiOFqXntbY3e5MkTeQwzwh2+HGqqRPAwkKUYZb8De3BfYqLAdAv2aWwThUjCrq
Xq2sFUWs0y+1yYf0B7RB+67KPanWdKKec9QmYq9mUnZ8D/S2BS5LNyPgihkwe6px
yvSWk33BggGSEOAcNtu3TBzi1VtmscF56b5vgP2MDP2kvlwLkVNSmdPLbhNK4P+o
`protect END_PROTECTED
