`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
X1lR9L1ZhTrqXb86Lo1AYZ0dFAJmYOTBZ6vsXcsQpL7wyGfT6Z3IIc/LK4nrYZNJ
ugE6C42v5Z2q6K72WdwlYJ3qZfQpSSYiChsGVQr1BZK4mOY6QXX2Qhi2Azvu46d/
vxd0f66kNNVWM4jLc/85KKYGIOphMf5HxofsyZbRvefec3PsgASt2IVl8Ub7ptrm
t2gH6c1Zju24kDbkWoteLg4XU/JSCMcFIe3aa5lScqMXIo2Ihdo6Kq0sXWHUK1rp
TxsfNmfn9LQY9/Mz8XqWrrR0CnkRUXxkL3STtT/6zGM=
`protect END_PROTECTED
