`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAR0OjfZmQGtpl9isCNjUBZs4hkB2I8Tchos76Dpvo3Ae
Sc2ks2sfMal5tvU1Nys44HvXb5iJib+Cog1osR1yjBxN7JXpOKok831TY+1LgZ6+
TZxiqjuNX7gn1356vYn6L/9Cp7wZkF1LB6TdWVWW6Wg19SXRP0tmRIk3k3t25aah
5nb+EzRSm+may1nQDOezuQO1tphN7q+cA9DWVFXy/BDRIEvJxsZVxXRav3IBQqIW
KYr64KquOvLfYFWN1tIFUjV4cZNVYgRDMeC5hIGw5AJYhGkNheeiuRIrQq4wtITW
pLacxF+o/bD3//3FHnt/w8H22dSlnI5Tpkm/qOQNLt5vrum6C8YTJQjvVYPE+Udo
nRt3zVE8YzURMSWMqpLd1wo4EHaeBORNjgKnF7K7hpqpupAX5V8Tul+NPLESN7iP
FVAGUH7egOordWIduNu8FWdCCw1AS939IkcY/HsUP2pxSO5vIsd4i622whdigtbO
Kh/yEwDN65S54oaPHLMfayXpvIVUsMqP4tlwGJo88LvfNjmcptiUqNE2hsxXPo62
3w+Pn0QsYxkJU3IzDDfnGnEiplIafUMxjTJnq6Sk6Y04T4xb6aCwF6C1rk4tT/Sf
4nXrAuqMy22ImMF4Rs0LNwdvOvepJfgJNd2iazJiJ8FvPkTRtbjjQN/ES81dBDPx
i/M5c/74I5n2I5akR+meT2l7IS9uAhwCyM3GynluzFOj2gPma2acLA8VA7Ztmvpj
UuFqKczI8GFPgi91dgSSiNfpuj56iK4qPcMnwzmAbWX+Zvg9OcWTJmGHLUw4OzVq
hzaSpt/Y3C3FoybO6U+cM8HYH6Xjk+OXoyjocjQMgYCTbuQS54WhAhK8+4sGT/vS
BuSJEtJa621KXSqzXQNgDm4z/g18XCdjlydkf9AEx+OyoENXWbCEGBCpXCS+j8+v
Psf4ZEcCIkMJzzYVWfOfper4lPpWpdTjlTLdhtY48Y6cImqJRNOz+JuOOcieUeHM
GHz7ZmDatQ/QtnkuUno3x4O9sb4VEzvcHUHKvHGnat3dOfd4klxsIfNV6lh/8v/E
93BwB64EWsKiNGg8QMonMSAvl3vm7RAi10TwXX32qrYuAk/gaRC4w0Fn1UwKM4lf
AYYf33PpNyq4+bu0cZB8Oqg4GNTw9m+CYqsbr8FqHPXH5Cm6Fa44GxCc+IaWvzNG
nplR+TFZLZdPOAWDgKCElfaWMISjdfYbN517231HgPugDOPbSNTU198KDsYfmrTl
41+fRhw2h+Xcvn4MmGj+pMPLg3+m1TQHOxNjBfW9yEfZg4pmA7x2dmcasKgy5TeA
DNrQ4v+gnZTF+hI88tjCurtnSE0TO6XHe9s9UuqGst+suInAlhqUN2gpdgWlSbQe
WITRGuy56qRmOVQyoIFPBF4sOaF0bqbukg7VnYXlZL3vLy4hgI6QKguOQQPTBOw8
dl7zdw8ZqKQAJ249ZaGlpjCM57H+CGw/QHMbogkHLXWwQciHpMS3puw3yQUWPtns
D83P7S6toK0ce+8NiWePv7BQBzep4N9v7wz70rzDbzby9ogimBD+wq47VRYNzrSS
/xop5zQL3hG9mJGKIQmMGxIxrM1pg3Btc7rIoNUXnum1aeCPok5ZNTsaf5lpPkpl
EjbuU95vqV6f0hRmXBQCzUH93STt05lT0KbWvSKsqTmOV71BJwLcfFKxl0OyY+Jr
R9zzQjY8SsvmaN8wY6M59/q45WStz2yWmCKFQouJ0JLxzXjBlKMhtvSeAc2UH83V
6ASfrt2Ab0YUbywpomWR3b5nvsLOSqgsdKQQb0INpYWM3j7Ll2yEXR2agbbvDIDS
IG+8g+4YiOrnIaAPBPNAWEDHItzr/d/gVAzqXkQnVKsr4ccg312w3mwajer3vZ4m
ywtdIjW8NfGv8//Sn8kDKn/xd3pnbK4jcAC6R43mJcNE1+lI5xYyoK5MUVsKszI4
7otSzY74MxF9vh1bown54/ZzCaI0rF9Bbxsc14eZaPQGLqTOuwNfZNnm/lZWvBu3
0G7sT2Qp/4yPtaJHrkNK95FXVtZH92FYOMF5UFpzUQpxzHu2/jt36GqNbr1Bwyvf
iiESsfeWTZXMVI/uzXfSrAH5t+pOa7Dr1fVhoxbkCw1HiAGvhjBodZ32MTJiiiIL
TDTX2n+Jr/OFOInarT4uq9STC6xwFuh/hMoQpHe8/VH+E+HAiO2aAn1XRY3FlTDs
IDWXlALaFrVqijLUuQt2vqAAM6/ewfyBEl2NhpXfDxO6UP3L2Gnuix1l4zWi57jr
Xi+vaQr3eBEp6Dw6hOWXiXIx6pjg/P64hjK+wvdNNLKd/T4xF59VTiyO5RfJ3YVj
h5tb7zOecX6L/axebibkSxAySR7usXjycDzNqlrSwOO7u+e+IIbN/ThoRp/lLqo5
/z3DOf+gqQQiMAobDT3Y1epKUoV03np7ex2OpyOtI9eTUTW4lXslch0w3Asq1e8V
FGdvNM1UUAQQLequDxMTfJ92kd9AaKtGvLdHsfr4PZTxrbnkZXTvgWVDaIhTuUjR
n8tLpWcVzP/uwBPZPxi4GGTTQmuDng40PMoS+lWoLXabj+F+rAHCPa6eoLm1R3vX
gnxJq2ckI+i4eD4ZwwLEUju4AllzKorMHvgZIvl0VMS8Oek8vtLbE/LkQWEbGtQn
ah5FE7zmSyigdFGlMoOxn+v0zDousZkAggjlOwmv8BNaqJu2cJPqgRF8eBn6oIlU
2bvS9QzV0n0kF7hI8d/0IMn0utw+Mx/Sx4BlZ8dyxQw4cCN/62S+kzfdnjHzrEo5
nqkITdyD8rAbvCZo0w7V44hs5AEXrjfbo5+2gLBr7wVZrSG98bWHAJ1Y95GAnyDk
YR3Zp9Ze0FW8dDBZuHtV9K1zGWZKNG62xOA0mR3mq7AeuwE9FiRD8RlRwXCHrowO
Ofj3+FIxqI89f/t/Shqmn5YMOdeg2kzqSFXXBPC2E7rDE5VhGMhkzO5joY3gyOTu
wXKXClFxCDZhetPVldCVBLWpKio4HG+xEXOgk9esPmHAJR4vsbkltG8ov010ROEJ
wgFmNUXwIxvRKOM0bWCl4i+U2h6bnB1OxY10GRj9B++UXJwAG0jm6eFkjQdORisy
W2/lE3usw9406D/dB9uw0ftHTuo9sOPjCCLeogRXZCFrKtTFj7MbV2QVO3Rg59Oy
gBQ28doRdT5nUX7K/IxAZmLSZWEKADOnAr/kFdnFKeqg7fxEyvZw6s0ppDqgI0Lm
6ELPhdD3h/sgOb+M0KxWSjAcpyrdFlenN8tIWb/5rqqyVe9/GUtgPh66cUK7gMPq
Uka2XOhaHpoN09w5qsWMNOooH3Rms8HqniCaBOq8LsDr4mPZQfag3C8kbW+3S1oD
Q+mG8WkklhgsFQl3c/X+vEuQknU7ihdy78ZMRvGSYJgWBk2gJCk+H/fnRvx/jNt7
NG+4ci3uNqZlu3tkX10vv4m0kq97O/sKuQLLfF+hIfkvK5cKdDluAVIyEMWPzBd8
OQGLuS1fVV1T52TGdOxBPQPUH3P1z+cvnybqmJzJcBl2+l3X7B2db0rQaV5gegPO
gsVi8KXbzd1QBuWq5jtKB0Sr21mwo8qtj3Ozkn1EzDnnYe4aoKz1PsCw9v/Z69cJ
qGhyfbQyA20FiqOP+U7PXLmiC/IPuNRxDnrkHlXDDRYSa9j8WjlpdVQhNTXrP/GA
vOrGsYezlVeY0vL+YHjTXIdCMG9+Bb1ktVN7El1+0Af0UdHvwec7X5aTav8iBKQB
ybdmMnin5R20fGDg7081b2r6jloEG1RK9C+yBzwhOlQdU/TBDiAojfV2/lTpDzVG
S1hZTccWfNx5LSlQjVcl26X4SmOFDOtmrPos9P5vOAl5sura18XCozns6/DCN/uJ
leUeBSTU0le4+JB1eRAgEa/MiQMfnkfD63PzsqLPORNEsx5uTvwBNc5vZ6FaSYMr
T3iQDopdtrZ4O37vYkuIopQxpmt4jF0y/2zFSoRqjya81qHckA5Q9rLG3EiJd3Fe
lcgsc9rqTYHM9AfuNPuwk98qrqk5/CWVVSn70klosAbWS+BUJExbrPs9UymdFreZ
9qXDlxvDvrRiC6LCGsPDttW+Wp+CkZaJTrp+C7H4zdt/tTDnYGgOKZ3I5i2bq4Vx
PfzF4cjTcSzOSlArZAcu2pH1fZwAwVhO2ER8lxDUEuA=
`protect END_PROTECTED
