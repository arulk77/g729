`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMOrGTCV5HBC6lM54YcQGb4YEId+c/wnlndwK+Hx6QRU
l5oHClzuK/1BUXSlY/EiPxyZe4iGa0XkWlEOO/ez4uH3ajejGh9npKhKniVLq1/I
zjOz34etGLrcF8tDnanatvYe7eG61Um0gUg45h5gKzYbrqKuOfcmQEF96xzqyYJB
foqpE7GPto6D7yr06OXRPw==
`protect END_PROTECTED
