`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKmRUlw5BftWlbW5zLyuZcEJ+EINfiMKjpE+vnjajFDX
Bi9RxXar9OndskSW83iqHrkLRKr6gLkNU/PPKh+0X5NXB8WioVPQ9tiGrUFsf1X/
fokDf5IXSmuUT/qd0RYFsS4ujuEqUehLm9bc2JVP8CtJOcaB8y0W3TDa2H9vOeUu
QKdin410BZ+43ZdYgHcXERSlbu5DmM5i0mG703jPgxnO/dh9wHKWClcnr5etkWvs
HVFOT644f3IMJXDaJZpRtwA9hx3xBkLgrfNlUcEwIeGdX/wR0P0wueCdlvRiY8Bt
Qr/eq/BvBC7lUHSde/bXPPaFfyzJysZDM2gmjOLcIbFl6MVInzq0IJ6VnHvMZXXY
ek+ymoHRZGpdfAFaNrbtD1TGHyXI2z66qr1YDDnQG2Eqzrrd+/wRJDlzhcAXfeF/
vD1XFUCE4IzfP9dth0V7Its3Ft4b4vZ0kC9m+SnFFN/vg0RaPJj1eYFipuL2OOmi
2afE809Yu5Hy+0hZYcdRLP/XOLc0LE6zovjt+Mq/JhUk6EI4e6XmQObK8fi7ZhaK
`protect END_PROTECTED
