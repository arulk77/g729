`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveA2JI0xZAXgxoBfomdWgCOVIeuP0H6+xKrZcIx8GocoK
4MuxGuyoW5YOifUtdickrsZAGtvMQTUojm/cql9dqvDG3rY0yaPD7xlHErnybitk
VJK7Nc/kVLuGq5IOw3gqXrV8duIdbXPW7foqAECFGDuuYpVaWCJB32FyS8upW7JH
02p4Yi2/KQJhivqmMIcAZjX3uqEopHzDEnBWizbuSmdtb0T5ct50BCbRKEY+mRNb
`protect END_PROTECTED
