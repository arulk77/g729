`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zAFLohyUR7oHwH2BB/GsJqVDjNeZgbEP9TNwoMhgToj
uf2YM3tWAExM05UoTXwmw4KHAJiOl7XbKuaFx+kpe69PqysHwyTSUt3uiqnISpAL
5dVcxhBmYtGkBFNI3+GfaCheRuYviDGFQcewhSP7vdG4Z8MJpcQzccmA2H+N44kk
2gEwyE6sDr9ZQfWqHle6RXCsQ2xnCxgHZq3f61RnV2VCiFyQ4kniq5zXi105b9kZ
TJnpaKB7o6pFP218py4f2eQwTThIo70ygAsxM6xO2UebdQ2hpbqdWlkyt0dV83VN
VzndHzOGPs0B2gYm/v4A5dmlnOGxynY7giEErYlOV+76t3aUN1BNPgXW5i7y+IFl
cm+Bp9qjKFRkQm4DsLWdrQ==
`protect END_PROTECTED
