`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDARGtWtHadMHVTZ9JKufFygGGgG2+PyWsKPGtpzNmH2Mn
vBzpRBWxfsjdqylJnDLSKTGAC6p1H+XLLqwF6jlWB4qJM2Xd/FdzMZn2w/UJFvkM
XVoNznhbCLYo4GqLAwhRDdSg9JVGixPFNe0u184j+pV7B6iS3yeZE2m0V57moh6h
7nDnPK3tLpi6rTx04CCBY8trC/bH+2asIIXqygqVLW+7vQ7ZygAQe4wC27CVMwTz
RzHUifcazWrN28LqUIvjXbHyZTWWXrgZzi+uLaQmsEY2/owGCMOK+3y17+6MaFUS
DLcOf66IUXE3QzAKg81B1Rrcophr6O3K/qTBETLgxwtX3gAfY/MaPn0rN1TwoTH6
6szy7avGZIqmPrX9xyoD2UmWoBtzkL7boLPjTTohbIsmLChLF60PZkA1HEvEZuCZ
k/CKULVIItVaidzHfm1ujXS5WGzaA+qzktvVdECbyOSuieEwSnzBboRGAu0pHocm
zHqxxqoehOafjNlv5JqiUyWt6VAeT23TZZ5ZzchHlqZweJ6ecw2eKJ8/OUU/G2zZ
HClZNxQQ4qYfVEXtLupTNBWGbixFkJtiiL5d0JsKu0vx+AmiZtytqdtMklIx6QZ8
TgpisBj2UDd7JLoThuE6U6wZCUlCz+AkFJ10xIyuNpFiWZSRShTzec1d71GoFl8c
1prj5MJDHVykewJ3vFpXY5ZRijib0SpfW3b6oNp3N2qoi0thKug6f6eLW8AnzqHi
v6rGCdqIC3RfSKNTgurUwMHYQA/CXKe4j4VX+ZWOqjQfCBmfnLcKdzPAWFvT1wbZ
B15efQajJvEGANkeNsBJc7qY/2FsykL82tPbVVBkUbrTZlFH/iGEeft9fcP/gRES
53r8RUaaKRuhQkiPf1tt3s1+gMOZ12U0Fdawfo98My/njyP3C0dkA19kiP93XvV4
3+m+PUtfGhiBxnn9fihHK0jfr7GZll1GYJlft1sHWIj9gAgLKpRmYaMIkM6++4lQ
ML+2uVqWSdOfk8ifvv9Hch3Be1nZULslbvUtbY+l0odqJeT7iJjJ9+xH6l/zlloD
XLJEV+ZwHonH99g5Ht+HM+3tcH2fQIwpFImgyKJ/SLxB5Gakh4Xwvh6ckirIqa++
aPpwrELqoUDOLfUWnTjuExiBNmnqbgX9k3egYFrmFWOwA/+fzae72PgHb0eBePAm
mHZIkB+8iK9je1H1Dt4i1SYsw6ltyrZ/mWILKfjVqw25QQuWTFeqHPuZ+c+0gLUu
iXd9+hSF74kFXVtRCKPOhq4b7S5bvVco2JXtaTKJxrueg3kPYDjSW03BTk1s20lW
N4wRV5hPq1k2cwhdi1X/fF16A4vWvzPR/G7jwQb6cMg4K2bCv0FZOkdoDKqNJhcU
HzExJRvBu8MWsJizfa2x+yIX/cGopxu2Cy5Wh97J6TDfy2WF3B6TCS0ehpQr5kcC
wih8pIsomwBkOMGE7zhe9W89vIDbboxief38M6DGcq+NfpcAfISDukNDTve+/N37
RP4nNEisO8TjmkfRusRqIahrldWWaVMmeJh92EQV3bhD+7P40Xg/GyCVSOusjsa9
QGSjJw5qbKKdrMMRnGTsN9dfMvFII23nj1kV7uUGhsDg7zmgzSosjCHXDKWqt/s6
84Y+YSoDz+ElL0GKDnsxqLsZGODKK3Tsu6pyi0/u4TsJGXdf/zgB6SA9in/zcB8S
ITGb69SGIWRbA96PzKMV7rNYqYH7IIwYSJo3osB6SgGlZnUomIL5oyUjgkSE9LdT
q6He2ykFREubjjGFFTbdulw2YcJJIye8Kw+Xq3z2b6QQsv6gMCs598KlQJnfwFCl
`protect END_PROTECTED
