`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAQ+kMRSAX6tz3gd0RBiU7LARhIkvl84ZuoVpYB+oZPc4
1VcwWrkT0TZDOKAK9+zMMX0FGTFc2vuM5WDMfNc/sYkzD1tyGGi36xASEDmidQJi
sCNcwhQB6W8hTC/fxv9Y+thQCmAvIZMGpu/v79qBXZDlpJ8khXTI8ZfU8fkMzsI9
qydstZOG8CISnIT00DqEP6u0dHikYUhnsFO8da9XiWUyfXd+E+8Thx/PrHyuYhHk
Gcnp26iZiPttZPcJ2lB1MNGfo1hWbTTvkPKcNX7qPppjtsdQSM6Zm1zA/ahhRMiG
9tiawC1urbeEJHGxtruIclgwO4inFHwEkpCR3UiVfzsQ82iUasVFxuEclOGYHIcg
FOZV4ZHB2V7Y6a2u1MvN8IrEoLpq1YwWlz7f3Sn6Jy0PBgF2tgxNQnM6FgbH8hgv
wCu7NDTIO97bEVI5+5IgNNJPfMIqXAU6RuQhetovb2M4cwzziWuRsjHohTzl7jud
JmvYh5qnGwm49WNgSXfw+2krKlR74YNF5mat5JYU6yfRTqHu6nyYSb6hzTrC+BCO
K5IBbvjnn7/HCLgig38JniJG4ElluVTjPq5TtYcbAfY5+XEgRjCV1FfXT6XQ9FCY
DArdAbgJqCVb+ID455+kXsVg8iOWsajCrbJIXyOnBoTxXkDmyD8qjXIfoNFRDvSY
kAWft0dMe3EyEcmsRuCKP6BulIVinFniOOFOphotF08BT7n4EPOVE3xBlq5b21Ec
Q+d0XoieezNRWoloXhynhW3J5ksYBFLgdkFYPo+YpUdTpRx7kz/HWZBDYkFeqeVM
9XEW2Gf2zK8eBx09FQYzNpPAwwZCRDEiFtPNuDHrdkg7WQc38Afg6+ehHDB6J/UH
KIGIwuTa/suZoSJwNnsCsnXn2jZll8sGnb/QFnI3I/pC4zhzW1CJTW0HhF5SCvIY
COH/Qk7l6plydLYVas7dmhAShf63YxHbh66+HpJVwY5C7hj1nf9XRl8pgmRyzdN2
OPRGN770+hkpS+GyIlMi9fAXOT2vEWhB3JhvO/Mqh8OqkCYBrW6H+IdBOJ/5zSB3
WyXTs/dyjuSPttXvYeSnvuo+w+SAKa38zou/EOOjiofl3Ofh2NiYXWiAim2lkeHH
lI31lnNUa4rUm/Nk4ydphvoLWL4RDtqGZKtkEuLx3T21T+5RayEZt4PFNj3xO2Qz
5yJUfrO3DF9ZvAT3mo9BFZyVGcfxCvNTo+LrbywaxqxkhDlrE6jL/VYnMV4vtcdM
9tfdLqgDAKCA5iLNe6BSmqTmgipwMO7f0o9VZQtFbVR1df/KZu4vsWqRSzwxiQmn
Mxu4yhq5lNdz+d7IuLtOd32QvCa0eBzfTTEjtcxW0ahLFlzt+jjtBVM1oM8WUCwb
lyxljOi5dOrXKgyzymJxKZJ52nZlS8RyyqqQlowNlawW7HwQV0L0wKlrHoS597WP
zSzBq0cbWAm82ju7fGM3Hr7WEXj5IB0N4XnWa51GTrWlcoX8hpX1StOv1YE0w4Du
vT7BfS8cgjdb0YmN7RHCDmevc+e8nKp/zsAkoltiN1b+/hOt+nqpL6kadyWosubU
117NX1Rk+qfqdGGZBg4jp4C7cPX5Z4gvFRNnQ8P9Aenz0bSJcLYEpa3DssSXzAaa
+82vGbuzvrdo6dG4cHDDoXxvCPqDp1AKV9zCaUMnFVWsjfjmWhFvZYAtX0V2Zr4h
bYxThAXSjh77kyGUkuQEMulWEVzr1qRc28w8y2Fpd8qqAMgTgq5KVK1tN/zqd1Un
`protect END_PROTECTED
