`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ZdZVIdCW3a5d/sak29KqYb4Bow82aJ1NXyceUWQoCxfIqWbhWmK6/NfJi/MxSqaI
28Lxjzgwob9wmqiXOe9ShhiRuy6DiR6c9/ghWk+J6GXTRq85YL+VIynR3291HPqg
6tfbIem7dLH9Yoax9vdHQdrkxOGs/4Xc/pjkriyWjg2/XF13KuWHTn45AGP0Ixc5
LB0Q0BptMh7T4rQxJ17TgF1mx5RBzDLEpt1JQDvJdCgmtRPS0ZYh3uHrfqFBA2kr
sf/b/3dObmma99Z7HyATAXwTSZeM9vXOui1Yt7roegYaq0vQPcDWp1KwZN4eTlbI
pOgyFlmwnFiH+OU1gvDPJ4MMKkBfCMK5XVu0nU1nyco=
`protect END_PROTECTED
