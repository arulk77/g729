`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD7jZeW02EYgXkZ5ICC3Y+KhPaIpRRW5z5sy8IwLm9Pq
PG0IzmbE0ll7AnnWCpjxeZzecCmtkCSvq5rioSyNEhXEc35/QdCKmGyU7Rk7D9M8
aYX5x2PB4ptI8brPXqixtgAfnbzZ06S9ZUOydaALyaN6ZQ13D4IXRQanHKLnGMZe
ZblEIi+e3EtlHbPoBjT6plt2eCGvCJM28DFpdVrixDFm4l/M98k5RmAOwVsr88zs
C1e+0SEjsvWavBLewAOB6NEHeuoI/0x3lJjLHhol5mL/1m2IvAtGdDJVFhzK/MXm
Azqq2fB0jSAzvLbvoMEXJGH4iT5RxipRNZCuinzxxU2FU0An6GTXk3qfCL+dmqcO
qFO3jSblLAzoUXrUXxUp2RDNi02abs13oIsOEQUIFPH3tl3SjY/84vAat0Dm4JPn
c7AAunhpfcHdZ1OvnWZZMX8/KgYlXsjQk4P3HvWbeRFoN47ZhxjE/hKu8aJKWbPn
3whM62NXlMsixjeDfJ7W3FO01SkyqscDioHMie5lZl14Za4RW7J0uAASNP3osa8k
AEbUjPOtkcEtC33ca2r9eV1duSSna4vQYsJkFTWFnoDtnmh5r2z0jZYYEQnPfzdy
`protect END_PROTECTED
