`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePwdk0YlaRkygySr7q/647sT/HlUTvTuapxK8Uk1abp+
QT0wiZ5PvcD2rAvzOSzNbkHIiRajtoYq8+12/+VT4Aye5Pj529RxAkt+7irNF24k
Xz+efc1hmDjKHbs8H4XXQ9ERmWzPTprCzbeOCbJKYhGWv3vvUqc4crei7+pz0NVi
YeN3zrnPTAYgUqUBItFvIp8AfCZDtin2dWfKFB7XlT89IbRvqPxVGIvY7zi2FfTF
6SLmrGPYJUvW2nQUl+ukItMEuVqeUKfQL3bM2gkM3NIabCYTP1jEJ9nprW52x0af
pZe2Ei9gJx/9jhaG8Cxju/ZjAvnBbbzzbI/E7YCib3oTyyuZTOsHpVHaUA6WX989
I0adubAZtUbWpbSAimcffYh/wVbM/aFp9m+IcbFYHPMdGWL6txwprmDvJoea9XBz
0O9+cxoHDt4QRkNr0OoF7MiI6+Ncr9Eb9MBqZpTkwUf9H5vMG5JI8MyRZTwonKbI
`protect END_PROTECTED
