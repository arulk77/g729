`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41b9I6f5GT8iCwmaCgybjLZES0jl/OTNQOAABVYPFp9o
WgqKBBKZEC9Bfa4kAJ2dvRSr6NyhP6ppnjQkDaj8gFrKvrX5uWGb3vO0uoIw/o/y
yUj2xCC01gCsUH8IqVc45K7pS3s9zHm54Gw4uhcxvZ95/VjtWsIAFBOe1R58e2OV
RcEtpppOnVEKfOCeannvLqihUrNZV+Q3WeZKihnz7jVyg1Q2W94JU4Fv0YvzJDx+
hPGg6Obsc+rvx1h0xkiOBw==
`protect END_PROTECTED
