`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAdo2AUiFFjOUTsoLpY2aloOkfb5clmibquCgKLAPWxv7
d2mmcUS64JP6tAJC3Nfjj+Mel+/vXjqgpNfdjd6SX4Uq0N4+hWkJW+A2mKvGQrIJ
XRqbWQ4RpPpu7pZ62u3C++8wxhMFb/ohhYJWtuVGAw4MR6eKulumXacxLLS92rZD
XO4NbNQApVYAUYhxjqJY7kZzZcUeFSwDAzGdQAPoGZdwrGVgXwEFcqeu4vCvEf5U
9DEfvKdGuVHOWmRO5yFFqBMjz8c0w+oM6sWusBNqpk2C3TkprJwv0l31BG4pE4qt
ViH7cA8QNrFzPgJl7NKMLT/aM5BZ8CLU2+ZbqrmfYtJbAS60CgZ87s3K2qx+gO+p
wNEKxn7GSvIVBSgwcFckRWp74SMs5MsT+m17aqAMga7h1uG3g36WUIfJ+e3AtO2p
089ZcyAUAlvLkSJqcmK7B7dvZbl46n7qhRdAch/axpPU7l+1m5NO/gUrZGGRxPiR
fmgvbN6GK1Hrs1HhGUvyVVOxRV13NiCCKzFp5VAmcYsDVVXFxiPPTtYcUrdVPyAG
jO73k846XPEfLKkW4Kr83k4jOcq8MttT0uaFBy9fIjCp36EyZgKlfrRbi2UXSObo
DoCUkBQXYMsrlRrqRW+RbAi3bCBlP+YPN5/NiVeS3lduNuyZxVFAAt9RTEmGdwTa
MWWenV8HawkMoQDg2/+UNuBnEcteDCzzXIWz/pQ66J2aosLfnkfIGqqx1rvfopWt
A+WYNSZsXymDvLAXCPWHswXd5U4cClIyEWzuLt98q796DQyfp1M1WFR0ZfRNtwgL
XCgitVWCJJ8C8bNOr6l73BKbajeAXhJuz/vQK8evk+k6dU+KwraTpt1g8d6wVE+T
cUo1uMu/k62+01mqYGFP93oUEClyDPlT0HQKi8tUUB2hhsU+941j4NYb6VET/4cv
EHnbVgiyRQPBsC4i0EeXuRJKspLljbF8nAAD1tRJjnNrupYriq1+GBbF54zq42ap
/Xk8J/Vo8HFshjpgEQsuew750EDCPR5w30fusTDpXZsHbyOncc/LStq1uIuYz1Ah
+F4h4mFgNLMN8GuQGTJNOfm6ODdBcpR6J7um8G1xbRHRAtfVPHIqvpImvsXuhYo7
e1tq9cI3CuS2sEiQaOHzi0W2MEdr1Gher6/xcOQ6vhTUOvLyJDl5Mjz5ybF+wZcg
5R29Zr20Nfp7GgfUGJ+wiKyIR3tg8MskNU1EBlIuYuWEAcuURJ3q8ccb3x+/OOOD
Cmw9CBDkWgI5GvkoK82Wks1HIOqgLmegVedVk1Sl7QT5Rzxz3f/1sLqEU3dyt5Ze
Nj4PF1IZ5eTzXui1WX36ynfoFFkco+B3IkIzKhLk12gTl/RXj7rwEfkrYo6X0YUJ
EkPk3XhgkfPdS9hdZbazDYAtFQKi95ZZd+dRnS2dlbmWuu5DxIIOwqhRbhd+W7kr
koVR1sK2XCwjA/WGEYjMpIQQV5S3zv6rOCQTqIoNH4NjyLV925ZTVqEssZ8a2xmT
oNKq9ALmAtLFvJ3PZGTfwH+JrTX5ngkOEt2FI89f5tToj6VlZ8/k2A1u7iq5buKg
8a+0B+xhSboGCaFNJ5PbSAwgohvYU65llJ1cGhd7BOXbAVAawmxrTxlVFF51SN8T
ChubJdO3iuNfP2E18P71VPMZK74nag/XSWe0FvYvbNHAaI4x7JRYoamQTptu0Yke
qD2fKj5Awprw6XvN0zvX6XkPIrmTZpSazCVIwzr7DEVlsSwp0M5V1XStsAp+oE/L
u4l1i2tLxW9+eCQwf6eSUwag71x0Mdf/fg/NEyGvkSW5JrSb7zHdFPCT84REOqr0
HWX0vVLGPNI13Ciq+O7LK4aNMeTVcB7anZv5KgAJftVaJLf+TKOi4LEAkBZSIUR7
mxc7jiYFn3c3/ItH6HdPIhBCEvxHp6V2FoCNfANVBWBXM31jvGnX7srEJjYY9pcX
PR0Z5WrC3joJDqSrvEAKmggh9DUNIkFDKH6A7DYL58iuwOCdG2Jr2ci5TGgK8rd0
woVXsWp1VGvSO7KL8yyLpOKCWvff8aL/WrF9HzCOfN+I1OJOr/1AWL+wn4wHXC3T
iobt84NtWIiUXgYtLSa/1BTPuWRlnhaXoV4bLMyqDNh5QsnG1nF0NFXF4SBa0Q+U
vJSjYnp9gQbpJf4zr+dAWEzGinIvI/e3oMjrvBQMUBgc/FtFgdMedPNcz4M6bs6B
MvWtJonMd32vBpkrHvHsilRJWn4YJ9RBX7e1kt4RxV/A5s4UTJSN/Qn8Hja1CnCq
2uIMjk0hP68R2qXlcm4nYm300Ipo8pMJhkkG5VCkzKrom7PLEZbjnpTIjAY0CCJL
DqsoukjO4ngUI6LkrkCP8dGxoHp2AGG99EbniwvlUSdWvfAuX/ZQxU+q85l3rAZa
T2Uy4XC+Qt2WdHVQ7g7hRyTaHeWrm+8Uay5ohRNixO8WuuxqVlMCC9jmwFIuD3dH
ImOZcRjaBOiFm+3hmLpqzyrWfEMRrmaoYU3CqYrDyDQfy1tNW2nSLzqppCztLRZl
ALPikLvsWfyOZa1sl4pbK01O1yV0ifNGHaynbsFcsvSpGyOLNNmY2M9Vl10J05q9
In0LYBoMgKE8QKX+LyiU/U9zFwg3v4SryaU8nFb7hYCV+rrWODBzfMkuoHUwJTHb
36zxscdK6Od0tMqnOXKXIyJdfRdq12lqPxVs12x1/mAPMIGE1br3NZB1DV0WAlPd
fhDcIIhFkrnN8qFQVfIJKoA7gvFSqcIWMjp5VUG9jirvUVPD+kGOcilq2jrzNnEG
9Ypc8Tdb2JYeCdOiZ/UKeG+MbPLpIUNftluZlsJwNs7OvYq5vCX9+BUhMxnsjmKC
CsUsAVArOgFopOsuLgP+TANnlIA4rnCUl4z3GAZjDpVE3LOkZTQApkYCOHwmaRVX
ndYAyWkNrCmUa5/Otl6ZMceblk/lIGcSe2q0UquV5pWMRnG0p/OaGpXAvEYAwIEP
Zu7MpShsIs1d9pxtIuRmCNXypR9PcbBWi4qhkI+zpp1kaFlu1EdgGFwUfaEUR6ub
wP2T2ciHVxxTe4LlonJjoKEmKHhvKhi16jqYW20+BL/sRUaQSsxOhB8tA4wDnsWA
DahiUjLUgb+CqQak8O6vPZPsKl477rk8v0ss3pY8t6vUkhA+DOsaAO3mqNKJhoYz
Z+D0qrW0PYl64zlSPo3mnf0KMUI+q3NcaN3vARFiWUGrhWL0350++3caxVIyP4h1
pEAwL6ynnMjaoOteZPxE+v+ty1z1j6dLkP2XAViDQEdX0ethhb7Z/pluNxyZ066q
5f0UvXuYFO4pULV62/6zTFvm6eAS55LsmtDR+7AJQreZ7XJ1j0LNdMegfHg0RaGw
tdeDFLqFyqHxqPYt2ORA+pRy4Hec2Ot2shVckLZL+1WMlo1Ou7lMsJki2POLZQHg
P2EVPa6saLcsMwJ9Yj+ir9pymuDrDEbzqUy1ee4Uui0sPoeGZFi3A6XKG7e+A5aX
dMj0SLXzgwzyK5FXhSiLvQ+mvzUwwGvD2T1tkwpZhpxgvBHyfknUP62SqdlSikZ6
h62wqd6CTkKi3QXncIyMct8o4N64k4cuj6bcLrvLVfbHeFXTyXf0EAoLZCG5mZcQ
tUhSm35rE96PqLkhEiZOv+9TLJu0RDlQEU0XkXVECDWZ1WRbLQWtCW7j0m+mgUui
B3MfrgxEB7d3ZwDUeYr9+OwsWwzXjBMZ6OxFtuEPVLhZ1ROiVJScfSddppxqWKdT
QbjlZ/C7mufJo6BtI+Q1hWdb36RLjuTFQj8FhmLXDX5jkZT++MNNfP6CUiacMDnH
lfqEliq6HCEs5pWcsuWITtcps2q1lgjHi+hnlE1/xF8NpZjcGwec0HodqY3yVDS7
MAIItjUX95EHcZbUxuZggVtayCWJbvhtqLACGePQhxiDGZm4iMMQ80O/GUxs7+OM
aTMg5Y0OtWaN8N1IfKgd7Ax4Ak/G8XoXBMn4cDqc818ixyUs9CAiBE8jp7rCesiY
jnxiJEIwPmXlHGGBikhVdZZxtzdMLfzv/Api3qqCxc8kFPS2wEDExCgExMAfW+86
pCaqWEgT+URB1MMg/HUgVxEpnYCij6I1i9h2RAIlMuHFCST3ps8L+63oTZQwFwDN
L5wauxMC+ARg6tJp8lW2AVsph3JE5Vf4MJvL/sGG9bWT4LstNdq1wYxvPbTZSUce
6CD4khoaA4dVuZP/P+HbKmHxq9GFotuxCdbug5FXSIAdjRnJItaYbrC7oVldSRui
jx/2+G7w80dQr9gj/DjH9MW3ilkGtd2vol8xxivxPCduch/JqI1H+AbiCSnwTmau
wACbPbYviRs/jtJ9TCrjUn4yqh6+8c71BPEMD1J/HHv44nsdJxmhYACYqc4T/nJG
QOFb1FwMcQV5HjRheLmK9x9ZW9Lv3l3YBdcaI0nfjQcvYMjRAkyEnoOrKkfPdDW/
G9BbZ8xPXfVqmWHDbEMWmK+8koiNgl4pt97jsIHx3sQtd5FXDdlA/L1mEQRBZ58+
A4m8/N6aqno7dQa7NQ3W7bg6JWz+aNozkNjzP1KXQnWpBoOezPoGsHWon2eEDDob
DEUTgCniA9EEsaKwEEt/cFVF61ZEcHn7UMCc/uhvmBdiOniVFKJYz9KCB0KTYqPd
coJjRZ2oVO7kE+QX7XpIGeoNAMGjTcVVbaPp+aZHij+dI7lEWZdPeKEk6NrwaeH8
n+G+IlsW5GEWpzKJh6VBV6fM89nk5g3XbbO8mZQJBgER9yjKKgE4LUmkpezFjIKK
oQsGSL5AO/ovtdFFEsaUDJ8ScIMnHwGRBqMOw8OHUzCGiRVKSO4Y1CfJ4EH+Y5st
Yo0SaWCwhBJCGOkj8SmT589iRsUyIiB/MnbwpuaMjTcfDhwFphOmFsEbDIpZnaO6
k3odsUxoQnzDyhH0+BiGeYJ12FlDpe2r5cuvlfhc+Gu4yuBT3j624dT1AwtOsZSn
VjxQ0S902AjWTcoUw6Ub0y7XgomDtJDNotzxZSVGHeFvOpABR8OM6Zy2pbxW4Ptm
ueI98NHSKZbtDVppFJUzfWKJKztC3/otm6WJSdjEvJaS3DC3F0cvVaGvNHJkPsHa
FCEP4ZPnEbNe7QqNhvMINv0tIK3Y6SAsaYynyczxtIq9aeseNwdjYect6tkJsDOw
INARdyK00fsQPb11MQTmejSBSKYOPqHs47CNK+CBvLkb6dSLs9oodXsgEAUwRwMj
pQkikaNdG1WK3XeO1xkspE/zLoI68s3uPsOlfpLYt8LTEL+vs6Xm+/H8l19mWjW2
Qz5Uvc8fMhvJ4sxoGbKOLoS7GuQhElGx5eEIMDMuFvk5KDaFRgmFXWNnoTXOXeT8
l/ivDA/lpndfZ95KmS/16DPgFhXM7zmOBwLVtHGf5sZfbT6Tn/k5MYWvevOSit/Z
6bo0jc1ln8B3dP/xr2W468kR3bUO7ShDIQCrib5hS2AxCKrKGBnD2UfUhB3bLO/7
UgvybESORwtykbYva3j3qLHP2PcDewV9IdFNquNIOT9WMrXgc+RyyIPv3DJkPZMH
vGS4PG31+5yGIQ2dYmCvVXjKbO7+CfdK8INHVCF0leEZw/G2ER+zaGgmiI+t7ajg
Ba7vyyoNTUXXT+FkYoF3pY+8K+vYk6dVBYJlRrgDZZJ3q26QXS8Q3XrZ/zV7ucQ/
26AWdldsUMuL1Zc51IZcEpTp09+RNAzxv+2RrEetEZmJtw7qHtsdqwsJn+gh2AMu
1qism9U6m5A3dGcXNIG2FobTvmrRQ9le9h6fYgJhmheEZTzv7IrQS6khQbbOFJg9
M3xeMKWuQs/zsRlpoWSR9V+YeqS96X1e1lCZIdEpJzEaYdt8KZyQOWROMOZp4zpt
i/TUeQGBqY5fjQsxgJ6RLST+Tlcr3kwWNxdZOFaxCGAMqMeVmgyNcwdjm+4gFXCl
G4Qb5pMkRCSlZsac6pQscHJlb4LnHuf4u2FkkipsroDBQ2ar9CLwxO+vI+3N7sHG
B7Wb+dmoRLlrs7U7Mc6ibOd6PAfPCgErF5NKkEYaBQEcyDezYGpDW19UvKmaYbJU
e/OD06Ky0LJKmosG4XFMFFh+J54mtlvG43naTajR+vuAY2QhjT+X7F7cswZpEF7e
/GHHembKfBCslkKr/KBzgpkm3XRS+bdn4QExoCLXTWDXZT6KYGdLhu+eVLmmenbT
Cxr/pyf2bbrxWTJXwAlwF1HvlPzPEVefPgVG9VXcwHaQSy13EQ3gDlZDYnz6fVly
mgv4+4DtfNfwOSED52FOpJS4OfAALkBhcDqKgfSTe6jpdAcE8qyTE8eMF7oZ8IN9
Or/l1hfkkWRVRoYUZl7NKHpmOKJG8nxGIT2ZDgAacQqF1E6GwmHETiHZchUA3Y27
tJ9aJivMoDvWSWa1dAnnL0hZCw/8xZRsFWkZLcULPvASTWXrtAwdbpz96U7hvBuY
rlKO9sJ9zwjXNFr1J4ET8SQIikou3tkYRword7X0t8iR/pOjFSogmQA84SWWu/pl
vu0QYjfHKBTXs3TrnNewZHUvKo5CGMVWSngiFyqdGiHGMwdFUqZHkP4/Oy1Uloth
/TenUpV5NuX1wgOrm+xyJh66FljRiwj0jdUnr3vx4QIlUKwBII+kfhmWKSg4qEL7
+R/apbkT/8zQDJrZ3Dcbb1tu4+NwEuZe2HlIsf28st739AVERr5GqNQZQO9eZ1sN
cveuWY/fPiFAatxb+CwNPgTIzg3l824HQtHVODCyFa3CQXC/+hlxFkSxAcjsc3Ni
lb0E6bes1sdSlt/CM5wgwWnJCv8d+4IbbvNnD8CFIg76K2C4yGJxoeIWgCcbaloj
sSlERDtog1+EV0w+wiQxOEhabnhKyybwk8H76BQ1mX/+3iewHks5GE+Nd6f3TK7d
Gf96xbOILJIWnkqcqBBtNSVqhhMDM45wbGwZ0MVyvtYUl272W+aCSJ+PYW7Ufqge
KcbPglm6PDFXnFXKq0sbLkpT3xnxsO7uIvB+leCiGgiNWe/jT/Nif3XX8KF+JUIH
jIkju0QYSjw4x2UqbUQKXMkzbPvgtwe+7p1ul/Vd/vlWh5uA0GwDEMkkGsuhQV5U
8wNgrPgdRkwUe8XDSznoAJpXbpO3qcnFnnfjBFA0X5ZVkbrc/cXlht97BqZPP3DH
M27GNbswe12z5VmkEI3Y1f7e0nsA4/3ogR5BWWtW+d+AQRwjtJE5zb2wWWVPzTsd
yLLyRbEhRRYGu5ffgb1Vmz54R/YELeuHadunq1mj9bKe+DMi+7406k4LqL0OfXGE
NaYgufMKtkeN13d/cjcpnaU03ZJDj1pffIw3L1g6RffZntitJqB9Z48hsfoOu6Ct
C12DvzxjF57akJZiRHdYg2kLjkIax3PPHwKdbML1nU9kl/GJgYQeK+13GT/vyum8
b2WNL5bx7m/838z22XTl4mNqgyydDIXLvo1qGRG3umBmx7ALhvEf942usHJ5LrwG
0jxfnBbI3tF9eeZ3o5XBgBhxjymQXD9/6Sy0ldUjqCLlQBQUGogZIarLixqv6ThC
4R5T51mDPhyF72BQpBWcJGZojg1K3BTcrIuWdJ7rf07IjwtxNca4pcp0OUUzZTik
0ij7yKKNSA/AytMhNBbvg0G4/ilnK03UAe7y3zXRs5CiezCJ/fFaVddDmA8PCk4U
SFFA41qvVx4BYvI8syg9iJn2I9wMCBMjc2TXZLO5TrfTw2gzy/eSnnLkrzTbVpu1
sSBj88zEajibp2GtHi0h968pVMAwX0C+tMvUMXDBQn/JOeopFJaEsX4hLdxXqFP7
Se/Q6gkA1QKEd3uGCbq9PnNuKe4rWLeFCbOhxlJwHIUs+ZNjZPigG2IbBPPkFTrF
Y4Ce5zAscHb1Ph7Rn+Ml+fKM+LA6hSBfTwhriXkc6v/bPNg1I/4ZZtZ1fkoRp76N
GrH3fBjNgDODbAo7MVf+goRTCqoGQXnmK+GfACGVR8Eq3UB2sWpR3FR0R65bHmsN
58G8iDi/9jUkNSS+Q0FmlgF/RVihlug7CZ2nNCl/1fmcuztWIMUAh32J0A0SD2X0
tjPg10N1jKiP/yInK4CEe3tQIopCPOcauRgGUT1cuIRYRon83eXK+aWd+tbRS60d
qUDtdNzIFjWBnC6L13v48bXLQJmudorNwQv6T+YMtJW0iCJe2zqF8CwMDr55BDc+
6DiZY6lBgSm0dE2HcslDNaYFik/jgvqu7oEtg0GB4BTvRH0x7HNIvbwDlpBw2vxV
4vxGlQmRs1b2EwcJIaw8BajOybPObF7kzXHBqZSM8HKd0pgBtJarr7tP1HThs0YE
rQo4wIXxonjYpmmvv+/DJeHO58mJcwyTwdvayKfyER4iI/gcGBQGjT4T59rScrcj
AfpL3U0KZkGq+xecHxuuvlDUxWwYpla7TbIPur1CeZuq9Oz64KqfMpBgPSFqRSeo
9kLFRGGhgBiH+nnqTVe2ASzbPSz1sTaKxWnlGpisyMx+ytF27isFXJ0vh/6vc6qq
a3fRXlX31+QD+FOpsL1izEn6VDj9zoaPwDKdlufwQg45GP7djmNNwzpsauXFL7gW
8F1fUUM7fq8Dy6ErPJrg1u2sITOnWFPp2aUKtFbolhLVAt51+QCoAIAglLPqfgx3
xV8IowUGBy5hlS+EtET8e4ddeT2+ZlQBAhmCRtWPdDJfYgBWP/TWrwysxELBnWe0
so4AyuAf8mMloDTqtlELK0LH63g5GwSLUmK3nFBXQUMFffjZEjNQrt6HVTgcqaYj
eNH4pbzSQjFpYMKg7ayEYKMmMkhpfR9RnyG22jBWJ2ebhjeKwRUyHVEZRVoi8e2t
kxF5cWIgPRJHc+nDvPl4oIOQF4zrnfqO8q8Jylt1XYmG7miRrTNAtaBSYILWl0Zh
Zm6Jq+rbB1Ak/ZjXf5CbuRpKxoYcjmH37OWcY1L604GZjdMf8TGza9PwOEbMqQMZ
LZQjXy4NvgCoA2p2u+Trit9AhaZf8URzrex4bXBo288MXSLlAH8S8BdDm5CFThNM
ybg3f/Zd7CmMit3I1BrEQ0PPePDK0b68IzpRQ/Pa8PLWX5i+JwWeOq5+c3YIccw3
O+m5sKgBJ/omEBqTU475JJ7aCPxcmhj/BU1WHOkQgZZbk6rbFEmfC4MRKS9reH4m
HzSm7QKdtLT8+tER5sagzLnd2Qa/pr2xC63gEhKLZPnyvck0yxBebNBLbV8mMJND
6qBF4SqPpRgqhehmOA5DLt/rEWv95AmC7jPsQq0SYNx2GTtoJ0pYEK8URSsZRQaW
XrCkyznMYhNf1KenqFPO6s0TLNgUAgOfxis1D61YUu6ld3rQuLot9fY+LMb80csy
Oi0/pp9qx55oljM9XsTJ4MwdtSGX2ukaecmdSMRu7Ta+evJ6pVcsZkI/iIAg/wO1
BxNRFhRiD1YNntwqZW6cGNmuqyKVS7BcRuxdRsm5Np8ySdeM/bydM4FCNOf3NrZW
UE8Ws/BUpG/Mg+mcCdEvcET5DqKxSJ+bL6AfYqHU5zuAAlBLvONJkoMWs63m+JrU
CGFU+zgo5YLrsRcI04TCVnJHTqpVLbSc0znLmShdVLqJf4itbe/SUkFAmDQ6hRZ6
nmAYWgaU9959glmoajtj07gTkmiNERWz7BaDkiYo8Oetw7I5z/bJV9a8jMpk2aG5
WUws01reQXl7LFDedprv3NNWyOnTdNeHlWbbT0N6gPgo1D596GvDQE1AdUaR6iS4
KY+4Gpr1p1PMKEvlwn4Gfzl2eMdoSydMsTJS0n1n+/fSGoQDggHlGDI4KRCjBFTk
FQSB9vOm4yhaKLXLhRY4EE29w7sIjd2b/dXGVz2Cw0HqIpfxQMZ957gFSBhrFwf2
XB5tWfGX0nuD2nTymxHVrtl4JjGqLKmCVlj+RZOwpg8sihx5fmHX0gHJun30D3Ms
8k7G92RiSNWSdmTyvVE+lak/FsCFbikNM4FNKBUSEThlLmeHWxHk9K0xuFbaeY0S
wd69iVMcpwLtoM/+RmSnESxj3tTLbvLe1zhOrK4r0E+dbGzRaG7oaH+BJ5MYMbsZ
o/AwB1f1510PyMXom9y/AG+/oq/pkRkFtARXNGW1wAuhSSy68xQ305Sw4D03vFDA
PIeyTfnxrvomgGhMwgRn+lgCKJ8XbsoHrbpJk2te70uRpEmTPrGe5D791XF3/G/0
flbbTGUC1r2rPq/7RNJnsdp8rOz7nkR4ty4Ow1for+MAR9aDBjhEDGv6fKmTniMj
RdJwgATM/j+M7ObulLC7yOSxgz7uhHzocd5HUSN/jec5F6km7R8luMt2WygQGzKR
8ZHCj/MVAg9qwLVsCrycwsxwcpGLjR7ysH+bOS7SOmZQvK80yu33nrM5nyb+jLmp
c+vUWJRVGNTJfnxmEvQj4PStxG29tMDNxESCm+8s/X9esksm5HsQAGKssU2a0H1G
iULgbONgdDY++TT3yNSQAtfwKIs7X4B+OhFDBSiCTDwbAeE0FTUNzLQbjx5JQpFi
ou9lWN+AGHOVOd0ryMaSkMSve41frLjOVqq8vk+p+JIcxgsxR069dUE4dZ22+tJC
a6EINtQVPexaghp2s5/6uXZKNfSakI2pvXpze1sxtfLajXmwbW+s65LHbu/r5Gs/
ofmpdWuhA2yGQCtmBC+sy1bCCDz617JtGF0LqIQiJUrVfnEn5+cKtW9Y7C6+N1HA
qegEAiB5u9kR8VDx0TtxyqQi3H6Zs9dnl6rXMvIO9CkHcjeAebV34KzfDVyYeGSe
TgmhpagRzb24ThG9fad4b7ffhRopghS6BkTG1ErIZ+NhStFnpVs4TwoO9AI1oSc+
n3JFRwcxztIYJsEsWDB3J9s8TndnTjRsvqo9LHJGCTDrtTQiJmEnynxXqjudCNpb
8hkSVxMHY/b6V7WFp77n1yDBs4AcKU18ja4Ko3qA1RthYQNO8Py75sU08v8ELcbN
E8ys2Strtn4wA1CIoPCkZP/Kd4iL8NFv1TOQv32jPairSNsZWjLLsZzXxM+YhWkO
hiEa6+/YNgN5mnvkWrTt2YAKnWYWnwnD3KngS2td8LCjA69XlYJ1g4mV+dIwlqiQ
XDx1olw18++7nwTYY/nfLCDkj03Kgs/5+KYSSptjdfUsToVd+P9WQgfg2AOMFvJQ
ILkG/SUnGRZQHffLR4FyXik8b6RrA63j/oKMPLbOQQfozawLpvqZTGGLgftzIGmq
WvpY0JCS9VPwrnPLzTRZwQ5sxxG3zpgGNKHPvs/YoccjaA2GmVNCQ0tHK3bOTdF4
Ut37ZxWbEzWqeMZNbQNPYSCO2iKoRzg5RXXGYTkMZVQanvYxf3/KwxcEMLUasoJR
1xTsd80sVCaNF5NJDXvQA0hTEO0YSZyiHzbfM4QhG10NwhSCX3Jlyh+Cn8lgn97x
yZ3Vw0Oy9mawonocepoYgV6r1EmLvt/8pIpvL/nq5EnNzjUGEnnzv1lvNnN8tdp7
TbgyqGi/UhP+LUyozW5jH7fAZZmrVVFYC6Y9ov4d03PiWPlgMwiZ2dt/4kGwo+dY
j5I5gmx/OWtaRpnsFcfakU6kUhDv4huxTYkrSfdE5V/RzoTjl5q4s3KU0uucD+w7
02F9rx/b/DZfxhQUH9c7C08Y70VbNM/3xAbN2OYY3XYEFGCcPqWH8rbboutDG/VO
5/YDz+GuO+Mq32uL2vjVjMgmvVctsoOufKDZvD8bGSXUmEgAAlzR6x2llHh+fj4A
jUU6A0viXiItLyYf32OUfxRnqRQtS7QIgZx4hvseXGfsjjxvLygqy6UQqNSi7jwJ
XNeGU/bWNkQdTAKd9s7vTB92DkLlIErUHv3MtB4/DQsV+C6oA1DwHgs+WAbRm6tV
nA1TE3bPVDu0tM8500c5JbYfTHNd8ou2FwkYE7q7/giUKBYc6AAflO70wG4zNQ6s
YAxOW9/+UM4TOmCrEx0G1aCOSr0d724Uamyc27vHihOLk1KckK9k4c2PElxgmRJQ
ouCsZuOKFdTiBnHVTQPx3GySXYkCK5rCiEKeZdLd+JILnBm0KJ4Y5akd+5vr0j6n
la0zsse1FJUihgMMGh5x+1Uv9RmU1APCRRIsubra29JTRwaV5EXFR3kXWjowamYn
o9W0JU6ghOAU5HXzTxHvYiknRqvIHfOgPgfmGReiq4HZMQuEHIQ+ItIYlSGkdPmS
duzqBb9AoWn0jkSehIAAjpYy3EFypV2NPXu0Ajky1lzvggbSrWfaYgEOUiDKVgCe
tkwnBlli0g/PKUP+EliAKOkxYQuKid4Y/59sSRpCnyX/u/gFsxusanXWoeGalOmU
S6yxq1hnVWbBOS8B7PD3v8puHIFuSLOWC4TTkHZkJKCFmiAyVHyvLAHK0HiG99E4
oglw1Y9ks9+Uwe7sOTveVfBQ48XvfxuDXKrbZN2y3LenRp/nS8sQ+HekZxbINRhq
hFJU7Jsqa0xwHo8Q9tUw4lUSe4aFYMn6Ad3NuyYypUnZsGxSrnaMd0qjXPkcjezF
SbCbCGK4lN/Kzch8d3rn8GO5Sv18rT+CRGqoTWw3zqtavUudhyQwPpsVnrQU2tRB
7ztxbqgDeqrrffoS1gGf9I41f0z8TyV2Fje80Bnrw6Y8SRe26n9tYV6CG2DhGyjI
SBVWqGT5Cqk39198ADSpapEhp37u03W1G/Dk0HRmX7/JSoL3irfXwekgrYAwj8PY
bJr3dvu/EF3joXHOXEtbYo4SclkTyIlFMx5ScFFXkE5vnqd1emVmygvgibs8GPOg
ZdGGuROdR9lTZfGEXRRe1iXBmQDryJ761REbgTUlzWmO5aoPh6RNJtKUNc/vvg6i
7ikH1/87q8mgbO7cDye3USkC/poVka3LVxvc8yVN6N5IkfhAKwhlPpk3TmI649Cm
48NALLZ6bBQPJE/vQ05CHATWg/BJKAHO13VtflWl1zLhhAWbdGBQmqENRYhK9xuh
fR6Ns6QFr3ngLIOu8rIGklsotdNTIpBDclc5baPokrQ0bSIh9XfgwLR74XPuw5wT
VWbYVw3JUmsMkXvAKeizN6txMwlcKSW4t6BVO67r/yKDu/zmNzj0gsvRC/VjJ7+P
Duoyuc6TYjaMuYO4yK/wiGkC5TlrS1U0GFrBHJlJ3toV9UGltB7ydOwaSo0pEobV
uke4UZy7F8oCY8DjiLG/ff977v441fXvnmCJ8P0QVsBfcZ9D9ethZSho4P2ciqdp
I62rI94J2Oapm0ru2oThORRMTHwBiBtC1T2huwaDzSbq1ShRAQcJ/AFd9GeVZW1H
TPDXXjVyOpgeetOyeRfOGLXDqBgkjN8wwxomVX40DRGmndh1uJn12ftCOhYQDP2A
xl4lXua8J+5sQSuB+GBYjuNHn/+qt/iy073dtxng0DJ3V4chsnDwMFXt6iq1i338
++TPnX+7zxwm+iFOU01GNwRmVByLNSi5YryrD5RnlAVrk70ahycpCqm7zlVb3EaG
KI1Ap+63cPVKesHGIRz0MaydfYWWKf8Lq+44CHeP0n146SQNhCETZpWSyVtN8Rmb
bQ80HpDoMK2Iu9/aHmzPxjLKRlJtrDdCv5UoFjBEo4U9fhlcFZ9F1OCMMf1aEIt2
zjoiurc73AJx5rVL3B4uSk2HnhlLrdsimFmNCcyaWO5LqBaZDGNOa97Wl7gpFlGc
mLMhOM8k/DTTCEq9cAe+3HaV3Fqq4Tgqznpn8bVrIYuPycOS29eTbGADpTa0Xq1k
/yGv1etYL9uLnvqMeuJs/PdVxfhm29+SgxSyArgZG2Hy2uxchtfswS/u/HOjqDpa
kpQOjlAyfskY/JHLOxNBbC2xQHq5O8fXreKq/ly7+P1b0zb1LSRBOH8/zPDP7TPa
9UZqP9GUoqoxyfuG5XBDBI94HqqO9+/iAyBp6Io1hIL33kIUwwIbGKtuJtP5q4nR
MtkOk1ECArhRSL1aXb5a+n9gVLbTTbtkk5Ksoc5WEA/91F7AmdkXAIWY55wZXZKM
gIaubgRe02aR6ipStZYQyEk5bLdgoQ4YPHpA33JB43JSezYOC2YyHJTDkEU/s8ov
cd6bhPURKD1sARYeS8VxwMLWKtnw1O6lq4xatp0D4kiusk1pv4NvkzJ8aJZESxwr
c2H97kJYFLSokST2PfnGsHOTy2MJWcsspFxDallvni1ys2NdV/knuRKcfrRnDv9k
rE5b2VMIMKBheT469BnWLv0YvQ3PJwmH8j2U45U1UAbl5cPupNo6J170Z6Zzhcmz
VXpmS7aMkvvYJfNB5T4aVossM2OBUZuS/F1KysZl9cfKAsCGsCZDyyXFS1MbPbw/
wmoYurYa5FDpcUv1MmsSvZ7DkNw5Ll3UWJIvfdc4mdw4T7cwF4vlU4H6RHksI6YB
1Amb0Ldv84MqbGEIwf4j5JuvLZbsAfCYolHfwBgkylvLUGLk9F9kb1t7hV8+HCfR
4/1CNMUX+4OQxw74vEZQIpVSsXVtoi/jOpq4bPIJzlR+LKEsi0OiieiDRa9XBvr8
SNMFcdDU5hXus/YlczHlhN5s+PEX/XL/aE+DIRMmggnBX+9lloHYVyTgNPd4T316
UO5Nc/l7mBXVrabkBdvYbEWFZFv1ZdqYcDg8UIX47is0nMqgvPQT3gK8nMiCcv5x
pa5tQT3gySDJcRYvG/MLRh/T+bqcuaiLQTbqdvdDkElIC1AirQYqntFiU/WWLyu9
UKqglE2vyres7aEV213qnjfkLcXx3Cw6rfqqggqLc69utDqTPzfktfF7UFQfrMzv
f9Bb8Bgtw8mJn5Qh7YzNgm9B8nX2UMpujQL0Qvcai09aT5NZrcnBKjuDKNWlAoU3
c79o1LfNVeKNgueZxnOgJaRmg+aLGdG8tdKYT4gmJt1a/WWoyTedWD0ZC26nEpzj
RCBIToTGD46VRVEGAL3zv1QEk5jxMz1XevuMeRO/p6QjfUFV1DRxpdEWdbTpiIg6
00z6XPg2gab4v3wcmymz3Ck4wPLgQjycROAVWHSDQ+ofCG4j2leVFxc2EeoTYMZy
FvCIJPh8cGB3GEnGsCIoV+xvQsQK9Fx0PYHb/ETk/nN3OmWM/sTvf+Ia2mUEoYuG
K++52St8T78Qzt0GfhsqGgySPwPybsOlTRHddMF3iGL5iflIdBVqiw1hiWo6azUK
WSgapkGgzTT2rg0ahP0vU/33B4z6pbQG5GVUPbQIVx6EP4p1ugptvvc9lLuV5fv/
8p4hNThJHkdh69ZCLu20kAOq/VJ+VI5vq3O/nKBuoi5MGgviRoSDriXjzzez/oQP
kEK9ygwtL9rW+KrCgh85BBtLtVZKL08K7aqfE1QiVex8wh5MUmvxoUybAN7430eY
iv1Ve6pyAyy1vtrr0JoE8fV4St3O6quYNfYDlm8vg0jr6HbM7hXE01UP6Gog+cjA
38rD+g58D6JvFTIT0s/MounzZ0hsHfilxqnwV2wx+m0qMzso0xBFpwuRNZFdOT9L
kF71vCLUZcrilcDvQ77D0xF+F8oBwOcIZw9ScoBkbHlqzQ4xOUXoEnjEKX1Vq09Y
mhAKrFTuMop7QE3y/EF+1YBBf45uPlWCKDuEOw/f900sadCQpFwRfysbD42Nc86K
kNWSSijz2I2XcA9KlTQdWHN2k6bA7/DAqDyoBHKKv3p3csM8dlpUIwGxzFhVleIH
FKmctTzemkJPp0HMgjDtkdCj04VNNkmP1HPy/r7YsJsd/oCv6jZ8CFx9M9XU6zyv
HUGR5EBq9T23oz3NSLA2ygSF5ChuuM19MuzDBnG6F0QUcuolBxMeDZvMleBqrP3d
vqqOMlcz9tg7bvbcMZd53ZFvi+JSZP7qZTn/i3M86zeesjAltYg66g2XjpUoEV18
`protect END_PROTECTED
