`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD0gHB3ffnA9XzSk4Z9Jxqu7FaJJexOpATcdulOtSeLs
Rdrdky0zgH3zY1gUPsp8o+XD0Q4OHHIPs9LM7q63QLtbNCSCo3JuytDlr7ID4qbS
JuF9Rgq5TtEj4SwlSXeUvQchfUqNM8aiNMKUA212TkRwU70slf8pOjR4ByjzvuV3
bvRr8ZA2pAatkB/yukI8iRX/4cxN4Yeia54EOCP+i1s0r2v01+tBAR/C8slkIPkN
BVeufGK57L9JkFccsS+5AkQmZVO3IMrU88CaiaOEd5ASlc+EgMczjVFn9NSq+h9R
wF5idNyUr9le6AH+Omd70zGDV3MmUS1u9L5jprsAOIOwn6VYQjfNj8dLjOEDy/aI
gt5XM6QfQUGPeG6BU0a2QnUVfy7meXN4iUGDUNFv3NXjBS/yo0BEOxjBO2JXd4mr
7HmfWRp/BQzMjTEAJIt8nXWLDryDU9xd/+RLL/awb+H53oEpga+NPPc5KqAoDe52
v0CGMa+O9NnFGbWMwO685w==
`protect END_PROTECTED
