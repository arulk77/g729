`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHgK7O1TbubXlAvo5yd55qv9dtVq14LzjAJ+olVNJzfz
YKVqZSHhb5+OxRgNx8RznQRivhDKU6wY5uKSZPr++juHADBvspDIlz9bs61xUR94
iHJBcQ2EnkZkQxZ9Xhn1VQDThnpy6CPKxeuLSLVzumiF7dBJYH0rs3PpH1Z1pnhg
NmbK2DnEmOHOUZqdxNBQBQQBzfGm7qLD7tFAWR5+WXj934pCMfvj5fz6/PnOj8y9
gx9Jby6GMhVOEveA4CRMFnqm6VgWn8lBWgX6KyHIIJ37pbsrQ+VF0Am8st1CqMsO
ZsIK7sH/B/FzV3TW9Te1uT1MKg4WbzJeeTL3QW+rWUmakYLQH5P2k4sOAU+5B0JT
GO8gH5Sy7aDoGv6LU4jiizgqV4VHB/R/Ajt0ZpBuSrY=
`protect END_PROTECTED
