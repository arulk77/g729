`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
5fonVpkuKyGiDvk4kbZ788DyHLun4BpGFU6xOJu5bp2pWPpQSxCHMy5qJ/P7ZVHo
O0P0v+sH+yK+kJXK/aIMniVl7ZfU4EmOXk5bjltKQkimgx3fbpU/iH5RVdrWsZaQ
z2O/nP7QqREdVsSoAd00C56EAaiC73CoHLLqg+Yh13k0m91aLopwLxG0piikvu9K
/W2FQTjB6LHVDSrcLkKlkASJ4BlnhJ+VS4HBb/6l/a9kFw/WfKiih1VU2k9Nrp6H
V+MgSzwZySNsrZuwJwOoWc3Er/7jdBPzf0KxHbp6qI7fJ+J5n9pV2UuZXTZ//SlZ
sUiI90T9XczD1JlHegiZhQ==
`protect END_PROTECTED
