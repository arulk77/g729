`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44a++foykZfzUBTEaXfA2Nf6H5bArzJw17oOAasWLMEf
cyRTp0f9vMBjAgV1c+O5LmJzu+iR4mtl1MYq2GE/z8JCwyNYvlV+1MVvMpNZiIvO
keQ6nzIL566EN8N691nfZwSWpMxnBdnNmtomY4UxgIQ0d9LWfAiL7C79JJKNZHSW
j6UYsvwCABizji8Vu74RlVO8Fl1z0e1TNAFyNre7KgLKOBstxSS6Rq9Tc6CdjZWS
HA9dym4ye4e1ZgvJWN9dtlQexbd69mQUjvZ7UtjIB+5qWyxv/o+DTTi9jvbnnrRn
pN1vEZWaYs/FN975HEFeYw==
`protect END_PROTECTED
