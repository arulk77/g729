`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEsuya5UAfPEfFcNkOo3h/ZROMPiYnw2472ZwEbY+XUk
tD2op51nSTHdcOPIwzp8vMPggdbeKRO3Fo9oPc3QFjjICA7OUY0e1zXdEBkZ7Tu/
jFOTTNpMg6lal/EW0SQ5X0INlbtE20LPVEa6jMTTMly9STOv1LBKJ00/1wkEDF9u
MCWuln7DtfOpUgakPNHsQfiu0j+eHCLdJplcxz6nahA4fY6Uoz33url88AopOq7f
`protect END_PROTECTED
