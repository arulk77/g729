`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wSA/JKLV518GviT1UATLt9pb4Q7KBKyKRetTSuoan7X
QaG8n8b5WoV/PbvN9xQ3KsxEa0hFsOgIRDNXW0j3CyT6/IO2eIyqpiZx9kN+FJU+
1ZGT2J/1YDqLQv+gL5FAPckEWlGuDGJs9MxfvUkS3osDDbidqibRHFeVjSInom0W
6vtkYr6s/QrBI6u8HPtN+F2IWE7zHwl1qCXUaeVHmbMIZ5TnHSR0hEMkvMx49ulu
gPhP/TEeRz7xGKVKC7lLKcCUo8S7R9RsFzEmQexmx4a6RFlvRY2U53uMVj+gBfO5
RDpyR7i7pFv5ZRmHlmXmig==
`protect END_PROTECTED
