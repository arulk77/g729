`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
6rDxg+F+hO9hDKPVvgTTA/RstnBX6m92Vws+ecoL1ygJWCNOpNaaFhHQBadTvn+T
QVGpSZMamdYp0JYbqWMnTeDDXAqSLMnFd3H11JYCDHZCPNqE90vq87l6vx3Cx5qz
AjR3Byll7zoBPzVCew92PaYx8hpgctVRpSYI3wklwjRYc/WZJn0feJ6y4NmeJe6K
W2wOBL067h8zcsVSzyVxWUsPwhVu9g2QR6mRsol0zYKOf+0yp8i0QCyEmnBetUa1
Ym9RzUCSTO8zKnpIG9D1yQFnsKrAlygDUygaZWNjkeM=
`protect END_PROTECTED
