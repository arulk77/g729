`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47Jcl25flI8hC1kLNhuMuY9KWWG4/B0bhnIkVffo7mV0
qZkYC9fBhr+egW2yr4KQ+x/quuVPZkg6/xSwgoOD25eR3YPxikvAT+2cjIhlDIY3
Jco/g20Im9G92PoUp7zw5GvE3ZbASB4BeTHmXY6wU1bZxS4gR2fbp+bmw8gCOF8n
FsDkRJyttHKo1PpnT1kFM9ObtTD18RX2KTYqUIC2/4S/Fde8HY0BUbNgmYitCRov
dAlxIJKWpf9GHNBQQM17irJAgUkPIe/SZ2GduQcLFa/manNVum4XBdJIOv3TN/yX
x9+B9v+7gYmgVBtCZWMevKMT+Ks2XC01Hin1p2EiEIprEs/B5/HxIKjHGpbfDGoA
Ax9dgiVijIWLoFdCD9uzBtRl6UszLVpXX+TdSHkCUNwD4yJUu73qy//+6/YiwDlh
081uvVIGjb3EBS2WYqhMqWSjJcYaen6vup4p+tm/eQiZsnmLDCRuKBfLo+Dd/0x0
`protect END_PROTECTED
