`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
9JEMag0WrNXyUwUhDdJvoLH+Ftu10W85rCIXlP+0/uVdiqJKjLwK5iFv2Y0HlNhj
3Z9dDHiqStX+miSkJ4v899dRLdi9rlF3Y5rBsVb7+ZkbJ8FX10HWnG5e3TzfmOuu
kstZ1716M77OaQjtzl40vNkP+Rf/935EKJ3OLBVS3MqeAL8SkCqiVER8kp6y+BMr
60lCkSkRr4+9QQgb39xJYXUKCqBbJrf5n260epg0ATppxuW0F6H4F+7ObuOztT1b
uPnGoGHCWadTvmM3nvmSUh5FAh2mStzDiUmQ4dFSaFk=
`protect END_PROTECTED
