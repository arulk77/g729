`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAbmr2J9Zdvk0Rtee8jPVOWfdSfr2MZC/x4GfySebeVd
6J2RMj//zeVIDSMvR4jVfFXpXjvu5GOyXd28H0N9auf1izNLDHqvF5maL0dW980V
nU34xn8KYnvTq8oJf0upI59XwFCIZ6VmEK395qzrkWQWd1p4lTio3exfNoFu5dHZ
UdHp8usQ2JNawRSXqQ1L8w==
`protect END_PROTECTED
