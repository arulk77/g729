`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAUB9mMd6OqAxtbcrZdRWt46IftpJ6cQIB1ouMycmQz4m
wFZNEs976zmkS5kyS0S7QoqRMFw59qCfuO1a+x/XJxsmT0F2BFpmk6QVrAOCNq/I
gHqLTNvVmEXt+4qWcCMY0D1VEbV4Jm3u+dEsyenjuED87MI8XXVA3wK9vssQGGwM
9u9OFn2tXaHVX8M9DK0pSbrMYzKRa8zsIXxs3pazTy7qNurXUhzJsXJTacuojrxD
bahT+pO970T3bImDMaPO8Qe2ePtYy0UbeKrod0mkiKZWJwCaU6dDv1AG+NowCcit
HRxLFjBL5WSeOdwfT20MarEhtrArIbKkh/kSEj6Vau///T7vCXjoKEDW7PF3QqUT
LswIDIvMtJWbsbSHKr/YaMZcbf/REPNSNJrsCxRy2sTfmI/kwjXbqRXPk0b5Lm61
c8WEHYpqrns2X/J1HyGFudpqH5NLCuwyW6+ZbFpTR9INcaKW82YmreuyWIw8V4bX
gZT0eTNl7HG7PAJ+QKsm7WXqbfnaKuRXsZ6mfqte77qCd2JkA2dL0cjT6YDaAeNP
7bTX/bMSfTaqAZFyQlsON53yG2k8PLaUjv70YaHKtLGuJlWwnRmHbgYzRhYmS8e6
n+7Vb1DxSvNUCT6IfacPuhCLMU1DceaTGG2W5kT7k4DEYyb+w4W3M1yetUW95Qe4
RxCpajeVHG2ov1EXUi2fj6UqTTsTMzbLt9+ww8dXgWdee1vH+8uJgOPOYXh/ZZsq
ZaOS7Wct7DMemkfgzRDG+MKQRI1p2CCBPgXb+dmabaDH6Z4AzB2kM+FLYxTcmq7o
HREkLj0nlLXmelbQ092Gz2JNbmrdt97xgJOE0CsV+lBmbXIq+ev/zbxTFPWm0ieE
gEl4aEk/h0Nb0wWP4ogt9ya3P3Ul1usPRnwJ3Gu/oZ39QAjEK1K8g8Wy5Ec+Bhyg
JH2YSLnZ3JsBOL5VSy+XFfLca+PIdzkwU5eOT7Hvte60yDs8RP/ET963EhouRgVI
arqDwK7sP7BGioZMiq916qlhLNQv+LEqFCtxeUFo0p4avKUv3UcEF4M/8WzxAZ5W
HYvEwHuUDqOei2h2R+jnjZhCp6q+HAO29/7Oc+X4VjB+xaqGAK5vYXtsZNEZDr7I
araP/HBTugpLGG+r2t09hDSSCCoUt1XcpOkSEXAsX98CyRZ+YidRT/6nsMH2TMee
b/wmT2Sgwn8/eeQNjHUqAoZhrM6du9dfVsJkuBgO/SY=
`protect END_PROTECTED
