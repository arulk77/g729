`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePPc9PfB4CqzfS/wJY9l0CzxVKL4VDHTB67Bb8myayRn
AVv50tO4ocH+3XHjaky6NJvUEjEdYf+1hbnLOALgVot5wgfJb+V4r8d/GV4fB0ka
6Z0GbeKlYlxDKH02PURhfhJsjWP34e++HEU8/tZtIJwUCpa0deHnPeftlBIzkW9R
MVPYzaSTmbAdWsr/0vtEKKeaoETG/qDcUFo3mzHiiiSI6ODNtjlRYsd4m4XGteMX
WjX7dqTHgT8Lto60vHeRALr/+qA/7kt/B4W6HlET8AXSILQRM3qbXTvMc6Vk1sf6
/o0AA7bw2M2088DX1jLGOYGRDNaYETjYmH7ItrY4mEKIQ+EzPcFs5OYqAMXzotG+
rzbTvZpS+ebMvQGxdqr5WqhZXSvSQPBE3xIMKr7hJGymkvwlUvfC1CRCtWJBIhK5
NroSbAd4GkYDCEiQun5ADc7XULFa0caBq5l6vLBzLwMwrbnePXMyaMVzliW9CJvG
NH2nQjL8lFZspmI9B9n5NXu1wnwiPQ5zhZsqofSKmPg6jP9+zONwpwYQAOkYhzC1
555KbbYmXjEw27qlbDlUXfFehZINzyRSFMn2rFRdc7nJbHGTBImh63ZqoeaHkVZ5
1ZIDgsZjE6+8/tJQQ41lY4UKuToEFBb40pZa1nHsOI3PMzLJ6uniZ6pfkB5BZWjH
SuCpCG6NQroLrbX5KGfXv5Q7vWMJov7mEuWXVYovnE5aHiR/a/66Vh+58IJmTG3T
3u6JQxNM5RNo0NHPSfd0ed7GVoDWP4yTArw+b7zdZJHlQQ36a2a+RnXzJsM5vf/S
dMDoysnlx0EcQ9g65uXok5o2dmyPaSU1LMlLOVYEKT52HmsiCZAF7xOLa4Fhi7Ni
6WcF80UR379+Nb8FtQoRXCE0GW+zTu3OULKipufj+79s+7H8eZRr883gwTKnZsSg
0oTUu86/JamaN0QWwbYOc4kNPhqMpEzRDrgTpDWQ4tacGlN4LMdu44EE8cMHqEap
q8dRFexsyQRZmIaiwvgvEVbmnTA50ZbJwyB5HNDrcFEG1dh4/RIzd/ALufFA+7J3
K+ID6Z2EKwnUUWAffbyGMvXiTMTNDIwATLxrkasnHucbfQm6bN6RILzzezFVfXjV
EyL3blRYhf5bTtuh3vsPqrim/I9hiius+Wpv5HPrQw9v0Mak/wQn0dgHtu2VnCyx
VsWbsnPwqx+njvvbWaQlE4EA9zzF+MVRuCzD6h1Jtq9kGFn1FThMVZSGf+yCS0Eg
w6+/AfbPQ9t1PQX4Sbkr6DHpXwF97vZF0j1gqQkIJcqJLKY6cedikJyijt05yMTy
`protect END_PROTECTED
