`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNk4JjbDHL9faVeViu/DGm+aPsbcCngK5eoxXZLCFsDD
uPH0bNiU+JvLJbXKO4RtoD0bIioeltWoBqseXEHhXu7PnPjZh7UyxW34YIOXRRxg
OyEn6MduXDxRLdo0pYubE6PbWI9SwOYl7JYKd2nsmJa8hDO/wwKtfPjNohr/W1Zc
eBfVMmQ6jbjJvJ90uHu9NMhE8q3pT9VSSzGTndsKW24XiDaeLL45wiNNX2NSZFuC
60dwL+Ut0sh/4HI5MfbmBDUur9Jh30ODI9nOf3Wgq6rtIiqqON2vC24/Z3Kv4Eku
Ln/2LfQLKsWpINsEbt40NiM6zF+8BT4BSk/sgSYog/Ssn+NYgzeS9NgGjViiquyx
LF13Gbk9luLFXCtAlRLRuioAtcCFdaT7ApHVqU1hMstbIH7uBjrP/jkokqDTauLq
7ByOR7wM/L3Fph+gbICI1e+XMlSwlsg01oRdPy8JFIVQcibBB3Rw17n+SMnj7uk5
D73jdJ3w8eX2+HQyEhlm3St1QjxnjP6hugwPn+o2LBzDYVx2IwX1kjQuETgA+J0q
`protect END_PROTECTED
