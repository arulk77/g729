`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ufZv73vEiMcAQ2Sr8o+uqJ4lKnDPMDjNeydNxzKZtexj8iQ+cDCgwzA8fz8g7KWk
W3A9eJU6KzM45LekjsXsFRhiXa2pZgIPGdd2rzRrczdVj1ccKdVUlMSfya56E3UI
6x4TMmLFj8/jN92LObKFVyGvaA/1IZEBaQxZbPBaXxksoqiIHnFsxn8X7ump1ftK
ib6kiwAqnJYN7orfBdXC5mxP6d9sngTqzcLgx8uh5E0=
`protect END_PROTECTED
