`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2On0KevbSzgQ43BUv6W6JJE77loMXshYx5togdrjV0l3UfcgkwNtZIjZkZhax+dQ
+FWv7ja7ImNuWx6Yq8oX/jjN9vLGGxAzFAnEu13Jg2i0cyt37cwpmH5Z5n4zHPBn
kJQoRVYz7t7r1Cy0wha/k1uM0stHnBg8yNQnGoQi7tufOWlWaE1NZvDgPcdgnLb/
5xORCqdhpo7KCTvz+KbFLMXT5RPYJTNESIRiaRA3c1s=
`protect END_PROTECTED
