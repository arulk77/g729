`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
7mR/631+9IKpzWh8qvmSfoX1mL9rs4sIuMkrfkxmUIzH8Ho81H74KKnIvqTVUBQy
qd/3U7CCt8UxCl85GDJgKB54m2thWS9iWAGMnRVftVNQbFxPF9v3drr04iJoMD9t
KHcoz5n6sQyZF3TLad9igL9Fwz+OiGiCq7hCinKsdj3YXdepr4nKeDkU4eV89w9R
`protect END_PROTECTED
