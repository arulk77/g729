`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42dC5hXdHaMGM60t2l6+vFaOox6YebE/fegAZGSyjM9a
C6yRtZCRapjPNg+C673TyonOK02nmuOoBllpbAFqNaC1rg0sPBp2aH0ErUhFsAhk
EX5QqCPHC/D7WGK7Vfjj7W9Q5TLnEbY0dxhSmMcR63kwndNyFjrCdeVMCpbkiyAD
PRZY7Jl0HcBoMOKUrpXm9XAHNL/u3CQZLOxOhh5b8/pZgZaXmAOrdluassb0tXxP
huXVkoQ9NZewWZpTWEukSgfnbuqiCJ/OlwjaOTT1Y2vlrcSUrLvJlzUym+iWJRuA
xyfJtpk8p+wkseDxuW5Dt0LMZdhVrovLJVQHEdJZH60DwANLdPbBwVdgFmIsHYjX
hmz9jYcXm7TgIY2Z+WR/pQ==
`protect END_PROTECTED
