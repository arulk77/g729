`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMlzlWRpdgNRuE4P9qZFxJaXDELVDi4CoOvPIQoxVuHj
rviHsjE5GW/ELAFa47iS5dmm/5g+eMEcrBsvkKhKlEGO89RRV8bgb9zq2QwwZ0/n
1s0XIkeJOwAScloMQsvOQ4LQtKPCzESd1doqrnlfgYmkjvljaKjMykpEMw210quy
rk2hN9nATvjHXHShIinWuAz6QxZV2cKyuqDXcnvQ0zBuh2LeQDNOJxf8PcE6am7W
uqpYrv2ZweWT7JZ4c0Dr8hCUOO8Plie6vly5fbVZB7jG4hRYRRhtSqMorNzcZjKh
`protect END_PROTECTED
