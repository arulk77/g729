`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveE88B7qdI+kVuB1gJZgVnMAyJ3PGbJtpNzbpnAkgIChx
gKF2TMpzKNXQfawMWTlt7lo2xhdUdKHjLM3FQRU5wWj9k6dXpT05QpFAVK5XLQwY
L1NJNGaa3aD2J/ZSKLtVtau8xZYiwVNqCwbQdsfpBvrd/DiB3mQjxDpMUOqxQbD2
FLbt1yYEdm8vjZTw396f+g==
`protect END_PROTECTED
