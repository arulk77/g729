`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SY9DBh1QLoYWqlWnIcKCA2etEEdUQXAlJERFeP2CCvUO
Osv1iWYyL9fAgMkgGebF7YzYAh2VatW+Gis5aDXwYIqTA27CD3SsC9cn8N9F9+cl
2Rr8chDQxf4xEpS9JDxIlsTEG6cure1MDqaI0f7zRPyf/7ZAp4+LD9as1KKcMKUt
Jb6mcg8bOu8hcD5F+V6TzInrapzDEHfLdqUHCqxUUqqxOtITkhvR7S/oj2/nmMWN
DYjQPVFXjYgHy+ITS2ucMCtv9KrZlG29eJbLXtJJGynDCauIjCT7uCJAcrVHbIIu
XwVYSvUd5EIAVdjF9WvDm9hNHjm/RVxl3wGLZopGeXoUvFsQZGabd8p0GkSLDZVb
qJhW0/0TgWihQXBjKocptOtIWqb4cuJA6kNpyobGTnnVfAqLhqulwi516kaixKJl
F+Ms5Hk7PLHC2B5pwrf6kruveLPY1kk8+urUz7Z0jXPWQFUNWxly+BsgUofqN72D
`protect END_PROTECTED
