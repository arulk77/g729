`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAW9BoLwhUzrqoObh5TeVtd3chwhfXpscfv7NwXaGEmh0
n2xRK8LihmTRUBIFUm8hSm9ZlXdVaTkBAS/+g181gOv0ONk2pi1DoTQ+KwWDe9r/
KmDUXvQyxKA5EUdhF/4LYcsGnhRRcQHWaIUgdGFYyeG0oxfRLqZ0yjsMmrvykgOT
6YGpq5ApcLDzq2SNi7QYVIPxA06IKLF1ElmcDekgYqUZ/XoZ4wPvUkB3bidzXMGb
W98jjpHT+LcUfCW7lBMhQxUhgjcDyWV8b1rwxIRSzTi5dkoEV25v8Lo5CkUhBvuO
QmcNDUWA9RJVYrml6GeaVCCNusbtla/hzjc+V67JsOfp571FVeGQTcSt7fWQkGmx
vxEdMheApgBwq218XJPVbZ0h65wssZmuQcQgBqxJu4LeXyyTda/mZImPeGzThiEQ
OEwGudfNbqj6CLF/Cx5FBdtLQ6QZyU2im8V8NRToHGSUEflTNyt4hFeVH0y7dq6l
vliJKLNITYLSAzLYiDifOmE4amm3UWgLq84O8LHqNKAniGiKeX40lHdu03fnYtHo
3Tud30mq1rdNTnYGObMSB6KE4nDuuWGj7Khk0shAp5wKPgwRwicSPASDSZEF/cM9
bChZdC6VI33VdZw/GYEwZtiXEHHnI+wOiH6ARano3G+LOIoHx7cDaUAWRRl09E+j
nmhBkRO2SFCdv6u1iAKsgLLpbQ5g53Eh+BAugvTgHhbV1laX5uTTeg0/wjzsFC8C
7+ocAHdW9lvZQ7yr++JMnaDNUzVAbqQ5sVD3BPmGk1geHoXchGqU998k3Y4UHPDc
1l0+8/GJfXH6OLq94MuR0KFnh5yKTwgl3hKgwzohgegTsMa8NQ8Xz0yvLRs0gSFd
hxLZTrdZPnb+EFhAckP/3TRpRPwSHp3fBKWAgwOpo9FDFkgXq6KywTUlE5DC6Vx5
W1BHRodhuribSGORGymbMXAhjXX0xtfixGhrhvQIuwjWJoeYbkHJP2aQpkqVNjek
CbMlUSAnMjgbU8kHN8UQ6oon36TdSvTMeYpR5EKDQ4kkOSAFwN/7cacYIBYIemeJ
MFPEXuEf2FgCmmkTamI/fJwjmxPpc1fF3bCU7xK4Mq/cGKWv8u0W2H6gEPWk7jjH
sG9yMlR5EcDCqDFOAlwgQRQyci+09ekdJgfUaBHxa3Fn01Km2L0dDHYEENX7hlAW
0ILD5ECq0FujBzZBgrIW2RJGwvmci9Z21kypw1Mi2kv5Bhwt81KeQ658/5bGQcl3
NInvdF0LzDSevn1B3zUzYYFp0MLHz51jZwy19ILey98NwH/uZ30cWYTJmtXfpwoL
MRi6h/elQHdmv4EZPmQqEMz0y5DskEmY45+V0upD1HOeufXNC6W/uheK/Bv9mlCR
sWP66DgrT5a0qaCmP+NYtwuTHnL0NondzZEIOoOo+6JVY5YaW8tD0YZccLt1VCNP
duUQ/Zw6SVAvwjJpnlWICKbzIqX92aEqMaoqqdhsjJ6gVUysoOj/xHMyhso8mfEG
QNa95xNMNsEpaIirRY0xgb5kZJD37NMSDwKtTiL43w7D3WIWE55U0brjk2XrXOh2
VnAeOWtNftcQLrL9cZvjKkmTrwJMi3/G/CvoO1ns+sDa5qhWeyVxHJWOpm3PE3ke
jaUpd59m7Kunk8iU453YBSnqKGhTF3oAB2GlqeVWvNCIaYGRUX2PbMf+d6LwhnBK
tSGWcRYafr6nJDcS7y1qddk3qogQ9XjVNItDKDAdXbcn9HwqhdrefbNauz230zvX
+DWYWjgXfAwpMzFQzqsNNLWDb7xdboIdjIFswH0Z8A2E5pyUH86Zr8Eq2nw908dy
HVJJSiCdWR2wGDTx1jzaX8VgNzkH15vBeX3dKG2FnGQNa2hOExMZwkzmZWt9iYe5
PFfKBy3oyii/DA1PLWSSHTuEihe0Fkhpm1xaO0Vp+VeYh0dLWpZfOm9F6iUngZYM
cIR+W84QKLvbgCED14y47g9/ciKPFR9ImUZQBfloMJqu4Tc0lZ2nEqXtlnGW6td8
J95b5HrRNkAh876hWlWRUprYdp5WOEVIkIp0q0f0chdL7t12YcWVAdJDFDPix8xF
EdMxLXPwZ3B+uCz0mcGsL7ZyInHqyGOxbexvvZFbjjj9vNmgqZQ1zm6PTclgnk01
34XJsj1uxduvhj/8EAXYLinc7AlgXi0vwsyVe893qsSnbAyvpy5vbfHVjjrp3Ipm
95TsLEdKKwBdy3Da2wiOBLQy0/u3t6TW82dfkzwZBnYciczW2GIMaLKSUqtsf1Bm
TL4zxhfJ5JyprnNaI4Hl8Bwrl0Y3S+b6oRJ1OOXxD/UJccFtCTmtV5l//a6Mj7jo
ZEhFpO8FOAY3/jTB9RFTZa5Kie66Palje22sKguxGa3qdZDsE45tjyBLi25YnO6/
EvoMVgJMoEV9PlCQZl9xRMrOS9aZingq9GcPcVXKhcc4XOuC2rn1m+QKewViiVQb
1M65QEEOYzhqUr80mRm2Y9KNMMbAE7dJo0ElYK3RSJTXyqg+6O2MpIlKB4qhrN0P
orpkXZrGm1z9V19Zguoz+JWQg5bOo1JWYPL/Wo6nmM91ov4vAbY22Q5ZuAx0oMJv
yxCJ3PSakzbWbskpjbsOpqIVAY9FLW//F1c4DZQ8MIRdd6vr2Bj/6w4KVaVuADWz
0rIuKV76W7j0FnJcMSdMS38y4K7cLVaJyFHFqH8vxQV3tEr/9kCHqTfc1VSu5gdn
sC8GQqb75LZqBfr63J3QROYsP8GW4OStQg0lXTYNuQOnqKE+xSQ9Ft0p4jf1f+hc
2fTPaRtZHXIY81SJTb85CJHpmVUf7AI+ok6g0ngjhnQqd+YwW5QOCT903z1k25jq
eaprH4RK0RAovSioWshl97ZVYS5M58rsgjYZCFLQPPUvKhhCFgL+kDzz05quPQ3L
ycmjWf94YMnqMtJt+TqVFEIjZp4zYL847quQGKCqUTV7NghiijV2mgviL2op5HkH
7hnAMhw/q36jMDgTDA6AivWd/GWrBhn/Cy6S0O1mW5bNwYp7rJ038TKfvTjWt6+8
GsCTFfBXExfFRLzAjmpPutF0E5ci+jIROqHzdBr1ACpDmQe8PEScOZLKcywPGS8d
KFCmXyMa8NMIfNsfjxY7Yu69lwmquV+rStK3KmXRMFv6BHxQPl6NQtjA+gQtavPF
6I/EisvGHCxf3rwAPUMH9Dcs3CYrJTUL8mjhaHXco8vYmB4jAcWtZejmiyYWGm+9
I/8uNFaBwusXzUV3N18oeQ57Qt6Zi3s6fZgQz/72JStYJcCoYMISv2/XczG37dC0
vGpG33FLevDJ6UJfLWDXhNuL+p9EXSuUkpapULduVt6BeUi8cHnpsQcCWRGdg+Sf
tmV8YfBtr3gp69LYHCGxKcl5flCBxXIp+1tGw5/N1zMCS7XhseXCtBiQD6Gc2wzv
hoAb8pEByQlo8Qdx4SkrurJ5blht5glzJk8WyyyfC5iNcvB71a3yamDHHLOwEweR
F8UVnue/l6ubACjPjdNqyRMQnTCaKnFEDGh8qK8CWuWdUZutN/bDH/g8EYpUkW6C
AzMI0SB0BwdDbl+pdalSiHYhi6NUHfSrYkliDcmJOQAOwCZyuPoGS8h0Y3gPpwKy
OY3Lte/K1XA7hKbyzpgIEH5ZOK7X0YmvBOQ28+ltMp2n9cdM/0n4mcePZx5g+2fW
APpuk5HDhZhbG0PlGILkp502kgcAfMJjpf0528ZddbNxwUJoBZZIcrRIKFmORttH
VG8jtpznL8CPTyo3Nf14fN4wzPX0Xs0c5n0afKTzqhbtTRxgzDnfUX/0XbyE4OQu
BRQ4FP/RMR3V4tJGUU97vt40ZnohAvGcDBs4A1NPS2lm9U9wzvT9DypZopGq6fiK
yM/1gDOts7gHHndBLkV4G8/rlGSGWyfyyAN0MkFOsJv8PDGSymbc52s8WpZLHumu
UqZpjV6/omDoYxsXrYXyeisCSdNzlGfDqWBa7f5P12GXZfYmWElBn0qauKg06bXZ
Jm9U0BCZ++g2nDIMp4VUcSuOj7+ZQdx6IR2R+PZH9t5JItrXnGV0gEkZnq7xywbG
`protect END_PROTECTED
