`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIj2oTAoPu22hWTnQzQz+LIMzkEGCK0mdwIWXKhr/Oe7
EkEgPidxhCF3xEsuzW2I5hcbe6woZ5tapYW4NQO7vWWiL5w67s7UaHL+wuKlBbA7
s0VfWmrH/ODs15eaECKamU0MRp7ic6fFhwa13TRaucPeqQREpTaQCHEZVBtklqev
658ZnZcZi2UERI0gboqh60kBISasV/nk+6U/doEZfFT5M3qNyb3Ry5D9o3AXlZ7V
ut2htZv5q3mABj+uBYKNHbt5ZpFhwA5dgRokJ/QO9zMjc/Ucwhzg8WHNQ5tVr0Rk
SXoPo0RkEcdM4W/ZjRdgAFg4JNSfaP1FFq53NctQCD2mJ2ME0Xp1sbIm62mGaolA
QrmyonMjRyZuHo86zQ6hHcVBPTfIMy1f8Kjz+Vpc3qOEj5A3jXN3YZwGGz5f33mt
N//L2/tgLaDfZoas8NeUosHFn7zHRYa6CWNtfRpnidm+L9pF/jjD5qWOmZ1Cxmdb
usJNP43069pOxvUjVnvmqArWIn3CUtLeeWmT+pyaE07jSgop6Z8oga7j9Q4jJ1Fh
LZeNZhJR0Cz/LneES9CzRtnQ6i+Us61pe6W15z8Mgs7EdFQ7I2Q3O2FPl2ODvPkH
o45U0N08fvIUmt0BwawPCaTw/B9NGcJFLLwmWs5AFFLvBDloDUPmUJ/QvPI37KIl
w4suZVWhVPLk3EGmiUW7Br49qXhr2HNAdk3LLZB6Fzes04WIjTsuBWVQ41BtGhY1
ei3hXbBstI3hZMNI7avVmbJqGm24ilsU8N/5gSSwHaJyw/HSA3HIjwAPN7cAPjcA
jqwGtchhkY5Y914wgwcgkBW2F42Ivz5pM2KQ+hb46+zcBcXUvoN/5xPlv5/o6NzR
CpmsVU+7rUORqlFKpBYR/HUNL+d+swIAbczByZRDjJIRnj9vtkrFK2NX1tMsubKE
DJnQ1lsdoKtkMP8p0U+8dkV5JxagivMdT2MC5z9FGGL1l46A13MiRKRUANiLO/vr
I9rkn9cvw6AjiOta721KU0Cl1Jv22Jmi9lifg6YiDCi7XeDbpoeOc/AiRjJiG9j9
7ippZf/lfmu+Dmia5+QePMYt6UJPJ5K2sIoiA90O3qc1HOGXL8Hz+H4CZJZ5g76f
3Hwk3ceigBcb13qtOxPKrYgG+IeLWDDGWBeKKWH50SFNOpQ/k1frba4LvfahTisJ
j5Q9fD94w64Z6BwvoM8GnxR1rNzJ7UHAT43AZ+6TBbSpgcAN5+Z4VbmoAkPUr+v5
ca4OQytyOFZPdxhoL5XHkSuB69CKNrNnzEKD17CsHzmAVV6bqSEFxt2yZvx2PQRQ
YxOdziV51lozkG/Q85y9VaStrP/D3Miu/ReLI7vXdk8plZYIaZi+7iA733lHQMUb
RJyiInTvHYpxaMwqflq7JRtSDphzhEcACxoaiUNl+9v9KFij6ZL7QXOZttXLhMh2
LMVa9IjoiYUvqejbl124uzJPdVg83aisJBLvVUZYVSx8SbBkd8F8tYU0LpDEuDbx
nX5WWBEjb5r43CA0Y4TGD/Zmd1CCPFILn1XQBGqAQQ8IytQupqG8CpyzgodbZsta
/bRe5kT6wlrh5HgyyGj8zorIWnR2bul4imbwwNJvFo8L9i8za26Hre5vcH/EcNn/
ZBUdP0LSmTkztoF1imZp4zBnaLHKJUdD7DdX/WcxSqIRa4FA1dTEkxBoW7MkW4nA
2s6qTD7VtDtJI2sB4+yB3IhMjQ5nHqfLz8UVQ9aYce30cbtYxFLmuSm36T3BSJ6m
ljfD0VnTgRFIv94xMSnu7vjPAvnRXsuKUAxPoHQvLnnTJf6Rz+ezrsHde7MYo1CF
41vV/nzKXF0BrtU2mvSC8fR2UB81b1fPlAWwJQCZ30AGXxPEIbYVBkOcduwViBEX
49epmJN54w2dyRv5iugQHeWCaosRhwUDjjrM5OFGnSfEoxTfz4nkJ+/Ao3bWy6bu
1ZYIJnPaD0UsIYBM9v7HA/UfHQ6rVzriXBz3s+/KAaOaxd1kWJ2bQLng4g2fiONR
bwgkETw83VuaS2MoqonsALiqFlce/g4aaATomN5xsOcqKsYGlkzZefv3HnXMsCWf
CqfPo9EcMYRZONhGfHCew9nblf0vB5OyzsrLZz1dOjYalXwOFMA6nSsFXlMof7vv
7f1WAi9Kc6UZqM/CsWASDRGftzxrtERs9PFxQOl+NYhe7OSDNopiCH324yS1If0f
y+lPd8vc+udknUtZydL9pIDn87mXPXqnQ41GFIHJp8GgUUZEZzLJVW3E9qHw+Noh
j45TpxbLICZFBsBL3rArg66X0rcMTOnf/IR7sKxy9fiWSgxFcZ+yOaEawM/q+nrJ
+GYvG9EubCfuN/uHj7foVgDF7OIUYTyeXoBBAGOZoXzh8RYuIOq4K2+1B2kA51Kn
rUqWRimVCW3Wor796WbBCUB9079eGG3j2WcwnjV2le7n9RavUwclW5nrnZP7pUkI
HN5vLN0g2N0SI1ar0g0czPislnnifteVSEwOjb9uo73Tf5muIqa1d39LvnMAGGEO
ZWCm0et8UkOgTk9K0qgZKGf7p2Dyt+ND7fWHcsy8bn7oObAyDHAl2Wr83qzLsOUo
EZvEieo7NDeyAxzXUO1m/r8Avk8sptVk0aaH5k6sBNhEaFO4CnsBVapDH8Nf3pxp
Tqk3+jLFsQSJfPrGLiWrWTo1Ya5gt2JViJGrw2ffTINDvzFR0nuJZG2msRBLWSDr
Y53Ay5VNIyeHRNEWCZi2GTBzydrCc9X2eXUlj+haHySb6iXs3EkLYA1ENgUzmHNr
ZmybSLFNB946qNkMkuTIfnzCGFKw08SUWtVB1H3w1UK1+lXHNkUirw3NDRmOFvie
DPt1HEUrWATJUCa56afHIigLtWkMYG6v39vcVUJUM/d0K3NSRRfpycKllzPZEI+b
+oasZTYdu9da8VjTVbCKnGVhfTAJpsWDNqHZywa5njnBrvqfrwTXK3Pu43kjuneY
bXqBKdE+Z7e+prixzKgAXV6Tzz+BDrgLihFnW3Dsge0hibPEQVB8j+QvXTWsbiYx
S20e9BlUopd2nKH1MdwNZCsQLUyo/WFIUp3emrr7cgE0816tWTUlzuFf7aa9mA3o
UaMHP4M5ZXb1VDJTymSCu2lEA+r36cD0gMTUL9/g25aPclvi/3heyFy+reL4ygdi
GlL5J1H7MSptjKCYNzS6T0n8UA/i8hft0IfONg3z7AMqiXVcLoZrLjvp96E6U/TY
LH4dzyXRaDbtrHhbNrovS9jKiw9snZ/EZII69nC4tmhdVN0w1e0Xj4KniEDR+dmG
x+a37Hicaknw0wJJvxZVylVZUf0hgEYZPWhVREH+fckBxCHvHSd1ha7ktz5IdnX2
zU41ZLKzxg9ZuwxM5KT6NlZac0q9+ZHOdy9Dmrr8p+qQPowjX6+GsL/lW20iqGLR
fg1kXQen3vVjhjn/DbNxvR0uBFOV/pe5+iyqqNlmsSd94PETQhOXznPJpcGpYh/v
sGGWMF9UWAwHFa8CYaHe3KD4jn7PRbQmJIEuHdFX3LEODq8jelLPCynLiE6zJ3Bc
bljekLN5Ub44h2V0raRbYs7hsZ12hwHXQJ7C1/UGghmddwc14sFhSb6QCIhB6HM5
69lvFuCWggY9cUrKb8jt/S+JY2lZ3oYFR+WF4zBWOaCm9XbQwlABLxyiekHBJrqT
89N7pa5GkD5k8mJ3IzHLndKiYb4m5yBdkMVWShoIvX8U4uS6cKh+xUV+lT5iG4Jg
BUhOnOtS0NCDYV2TJKCK7z6vGeB/2TUcf1qWztL9efBjyJnjItNMJs3H2EaYp3Vy
upiFUSRe28H55c/nD3piO3ssUgcDZiiBk1fMnSCN1WPprQJYsrARNZY6GfBTqUw5
ezvhQu/N8oIPmRjMQBdpNmkMzLFWNDQBmh8LySarpRiB/3l6K49COSTHejcLuyJ8
n+Jvjcv/WAcR2qmx3cShxjYxytw81eZe/UCu1B90TyuxWObU5KBpzpz4WHZdn1aO
DrxWDJZkodPmZV7zEJlMigELNDNe+SRJXJ458iQYu7ZZ7iLtkeHxwkGc22dCliZq
2SmaWWNP21/c/H9aUh2hJHNvbwcTwbDTJ+c9dP/Uz2oGW4cnoVY2HFu7BLdd1u21
hMlOKOQvzrE/veBO5gixx3+A8MPLfN63Qp5O+aA/f0pG9Pd3hlggWkPr1p2CJMav
VZmp28Cfv76AwpkDhavWCwYRP+kTZkDC5iMPYsuTSi+D7ZOr0VPevd91mR0dhgxn
bjBogTZybNsqOfu/+ChCO9vfh1O12xuxlWedaiVfEmJuMoweDrE9fC0DcX6N2jQ6
XBEDLkb5YjOey2QAOE4+OUOR1femmYuGIOIpbuCCD9jY+L0Z0mxmtGo7/6C1DNE9
37SX4sbhmEm0JFOcw+QJJkA+CPTuihqzcjgqMYUeQm/FEB0hfC59pDJyCwdxo8qS
NNzO49jIbagD7P7BCZQpNg6Ckd3IdW+R2Y4Uvumsod5aUok4bDnHyPE8pnzAl7VX
pwzuhJVSHg/ORjPJd2XiQ8nq9FoUpw1vB/+5EpJRPCCenbzx72efe5o6Oq0XPbFA
sV8sZl26PYfWxTxsSuzXyNz3lIkRZ/Hus/E+DCMoVxiTR5KyQlejSOBfbc6uACUO
2yBplQE4OYfXBHFcsxQV9sqG4oIOYgTRwZsaizKYhfYYSN7mvslsrJEFZjLGVHUM
9qo4oJlvpfDCDZ5YFWHLTZieC+tkKzapOqYHLu/WXQCWTOSPMPSeXRUHj7tljQ/9
wHD+i6CC8nHa+CrZStlPCpIzcWZsFFBRBlencX3JGXkY9MBWXN2Pc8HPA2VvbP1A
IlTnFhegbHQoma3/KiEc3PK39auBrluxTAtv2XB+WbpO1u2aaIq2HB+ByZy1r4en
MSZJ0UQmpNxYFpD0eW6N41EhX/joqHjr8Se0QFbwKLvYpqc9ftbzOSsd/d4p7+Er
kbufjjb7ZMNSvRABqUs1pAA9+7ZqSgbCxTZ9M8gGBnbVp7pi7Vpk6Ppic36RkqWd
fP9VmEjASfgiYnh6XxvT3rmeschRLNXkDnmFm29qPphKUOnJhEwROgiwmOySY2Ne
7XqxEEdxQZ3y9u2RqyBbkwl5miCiVFjjpmPenT++1u/AAJOG/rPOlozW2RXD0UEM
rxjjg47/vmOnFfwk5a72AP+/CzGIucuI1L6GPa9nUsNqoHAG4iwwTP0QTmYfSo7X
dkvF64W71hB7DDMI7suvcUPecfZJsvbVJvuj3gXZ8XWsuAYiy2773ww0rbkdGIEn
VLMZezShtwEZrOPkRjqQR8kARuhZ8Jh6brhvs5hg6whMgFGWwomzHOV9mMbeHffQ
HB/6LTHPwozmcWm0w/KYErtjLtjxMRDuSj/TPNwufST1hg39ytmcU1dPsbFBsu31
8xLWT/qAKdjAMvGozyLsgt2QbVdZSiH+W5jlO+xLmuOjuQEVo1k12qAnYFwRdJHH
5pWovT3+V3tBjbu6jTgv1d3qPk1iB5TLfsN0aYVA+LLBldVn6/oa+0hyY+e9c/QA
xJJ+CCYhE9zfxsm7gA/MQVXYyuFM8npT6jus5tK9itl6ezKL0xPUnHwHVcUPjZex
xDFzPvI4wc0xkqFE1eTXzVlSs8WFYYFDp9U3zqV9nsEUxWLntw+Rvzh/0Ga/IXla
AN13ALTyxYqUHPBn9+zNWmyiWGpmSzRHlRCcMGOd8ct+gkafT3qpjsBTys7NeVqS
9UmpXrb8DMUxBeIlvwaFaKIff5vJMjTNtvzPE4sd3nDpvZh52SD3wT7nybinDR2x
bLjjAU2OUq0RJK/UVoA3WgdhlD8G0jIP9/bOz5mOP98hCJd92DkG/KQbz+pxLxZ/
sRCrpgsjOm7nHDh8nAmVm5QPONiIKdnCw+8prwXcsASvAhFQDjvnQ3gL6fzI9afR
DjUKsedeJs3KjB64vsb4bi/mmE4v1iDnggt1rIbIF7cuvCkrAcrQiMvduJuxof2v
Hb7gMN18u+NQWrdZkgEWhzM//Mox+zgG/3PzubjsJ0OkdrLijDqCPySK5LCqrl3l
n4YPtW0G5nqekzQWk7Z0iqKSlywczRQDpQlFCm39hfvgeDNeCV66JZni+qu4vSMW
1az3OsAY2TssNNmKoRM5C7sPeCrOYEKrFdQgdfj5hIjjWotKV+nQTU6/J9Aw0eUo
vsxnXI2suXsXu0QK4H2zHJq2FRgj8n/D2rvXZZdMoAtRstbnOyHH0eRPjGgfKCJO
oSCk/iWoI922BYozianKx3utpF/k91gr4uj/fPym1dKbeyNyt2yXOZshuOuS3mMv
2wOp/ZX/EWIV239C/wd4OiXGkeIdXFWd+V0HBKWSJ4FeOxh00kxaO1drSMHJ5eVP
14u7Sm9vSONlqA1OpUbSH/Grf+PPmdnhiRWhbqgCwLa6LNRwTGFHX1fSlFi8GtiJ
gOq/yK9H8Lzsb//7lxEW6nhYwfrF2LAz1RXK2cl9wU3oxlRfuj5nub72fU/8FNE3
3wImi0XQ/kB8r5ZQc5BmayzbDWX9RMhF1YubhzDOceqO8HPyxoPFPg6eDw3klp/c
li2+0Stz5S5pcl5wuiQH4LjgYvy4dXWSky/OVAL3i2KpAm+SMGHDcCLNMxin7m3h
PkyfTL80b72Mv/XOubIZWnHjQdJPu9vkwcgj5OuVAffTBGKRNUz4hlcRIawu8X2p
t+1VlqZLDGke4Etn55C0E0UM2hdldP5mofPWuLdSh+uysY43OigOzgBVwVbm/o1f
eKOYNUhZuHbOi0tCru3v3DFvuNN+qBqoZpmkG44pTVAyuj35NVrKe1cJpFEOmiC+
s8lKr7fUMPmS2nPdDMaZRwrE6xIM1gkdrY/0sOj04xB1Y3zSF9uemdsSvwJromH5
HU+uooiXyuOflgNLislQPcdiD44x0vVOBrSzq4SHKHyG4EBbFZwOJzALPFi0ep68
5HUbcGaWI18+DgU0BNDpvOHiXHubnn3SlzLv2ztenfonhFwcb5v5I7DUW4FuRIgz
Xah44MhZm/grX7p14zhRPjZ5UsybMbYq/Y2M3xKcVar1NoJREpnUGhmlrkdxeURy
CMoHRczQGf5ve5xZAaEB+k7dL9oY8rnisNyDFslRbm5GrW6KeT+WZdSXkLcFMI0+
onj7aqyDg2MrnHfvdMs2XE4eWEe1AR2DPI3EsTN6qvreK20KtRCx+b8Uz0WFmUIO
yjG84zI8ms1JuHD2ClUtyyH4I0sH3KxGwpBqBGv8blAfybkL/fkBZKH4rSMcE3Ym
uh4TExPBTiy+vxysFEqrDMpvpVgEKmLvC5TkJyYAdEx19/uYLd0YLMdIv5ExWr1L
kCP9aC+LUyv93/IqTEkUCWq8mPvPGA+lquI1f1uHqm6S0XpaHYkNREX1jA9Q0K9S
Ivh5KLxPa0CJaY+1RtPhl0fwXSEBCj3N2etxbBQAwlYdlM+x18dTxT74XkqC9dwX
boKCDrjyZabruge2niS2aKI8tOxQ4ekE2bXlbf0OjYhE52WMUBSIvBl8964jzfWn
K7VxTydTOSr7utihxfaYP7Wvhbw3kOGaqlJw/SAUr2QCJgNhGwX6Diz4AmCXQmYS
zYQ3ju+p5dR224O8wPpGPlKzR335fT8lFJKjuBspOUFSp4w7mzKrUsgdRMn56uAJ
3vRmDAVjF1XhCmAHEWBbCA+JEoRsZuhqL4PGnOCNFlh3ArF9E5HnQC4ljdhkSty1
304eauZbOd6GBZzWnMhX/2NbOfLdKwvg0IIDKJMC0h2MEc/nOGq7g5mx4lDxpAQI
iNjmo1WjsD5hmtL+rfJt+eo2Gf4MH0evMWWpFFT0iDXGWWtkhe/WD234kZibMCrN
ktdxZlGdSZ1o2eljJznahqvh5FVKu/7jfjGcIfNJIjVTecw8wktXFPlrqv7VEswm
e6G1mGQ+pWsDupZlfydO6U67f0YofCNVGVadxGDfvQTBui/9bXR/XTnFEauYlzIx
gxdg7mrdSLGKF2ofa5rfIkjcQBveNCOwxWzMubnFgq8FB8ztCZMoOUUQ2m6XU9PQ
rTN2iQss492X3JXHBXfIkpOKkKAYQHJ7asd1O26CrMSjJANXNLJxxsSu6hOm7iBI
xjR69r+HhdwVflItU939uyWMc+kVhYcRXQdHeBQSfng8XH6kPo5tCuipfegk3G6j
chf7BHCZ9NGHYyRtnmhY1r1X8mGU0bx2RufR8A9rkpQPlSlBi5ztPBi038c2sMxa
fWZLVznDcbZPKL6Kv9oJH4M2ANviEkQfmJ8Ytku5YU0qnXFQZyZu6Z/KEVdIhfE1
8lOSc9tsXizQ60U+5lZ1nJ0NSJl8zVpopg2E3MmNPlp5EsLb1TewLglVnDl4Z1/Y
x75tWSEujHVVRpSS0LXKb8/+ZiOcGuNBxaT5CIjW9TSfJbwrSkf5S3WS2L6T+IEX
OC1q21PomXsA4cLd7GGO1xjPrk442f7O6B+lGHa1nBGI6C2Y6ZRZoN7+vBAB44B+
kuE/Y1R2s812YhFrEuJQS5TU+7dsD4nvk0AEy0ISCTiU3+2UiRDIIgAp/N3tqqpZ
0RSq1jOyLnNE+wVKApIgJ54/kDa/SDyCP3/1HBvZNU03UG8INpMgKN6vgDHmMi80
cGP3dPKy/ZYb+vIbRSqd2s5adEn+hIA8pikghVuMzGG9971SI50GvuyV71ezYnIU
jKrEX0Ree39SN23RXOL+wQm2GuyX+596SzY94M6xQFFNNm2FNfxby1PJpTTYnNdN
42nL/PfDFaJIKAwIJ0g4UMdy/HXhs65VQ1E/wKWJyGYjGIfI17z/mUBMMLLcyGu+
a/VRvpveCAScmU9UZEgdt7q1psbLpzt6zXbhk9p9ZXXwviL6YRAg5GqIzmw+oMfJ
QIoRyHAF4bebwBIJxXk6uOIUCmemNPvUq1PNiRY8mXbA9R6UEoy+QQtIF0ocNMUZ
FuQXKsHNOtpYDiHozFfnhsTD2ucePxid2+SXoxgzL5R0lapVtJ/yL5uBzmlpwNUc
xlqjCVMNknvc4XgI7joeGBXfQT+nit4gJjs8ZAVJBa+q/UOsxpOnXDSKPhuGeOh5
uG20sxA4mRDVCA33FaY7KiI7w8f8EVNn+JKll7q8gRo3H9y4YNBGjXvAgdRZFRYU
g36A0EyRgzzqMpwc2MihHMEDqXYhQYJbccWfuyqVJyVPVKMSz9wUzLHNsPUFqvRt
SG9q1thmjRuz9CHq4S8WIXRF5UrCVGNCXf29pX61BnMdZaSeP+PNdxTuTaUPDpE6
kMoIfdau4z4I4hG+BOQLidyHZlgCbswgYFw+4iRrCCAIvkvmMEwg4f0ydioyd+Fq
0JY3PyxJ+mDZczpMMVNAdK145DweeeojPCH7P17qB4Stbbdod5slzchsBJpia+f0
wU2lvUtWywgJvKCnKx2QPOTQ0xr+mzLlWs/L2EsunKt1f6iQftiP/49bF/dfrC3o
iH1xi1FcifcqnTq5PCH5Lr6exmTqRf9p7F2Dh+HLZZcU4Zde460R39U+BJb8vxVC
UCV8VqYPGhjPUqggxE+jlY5zrqVFum3m8uEhd52AOxyJ10oJQ93Pa5jyhMys7Ft/
eS3F9dJ8yAGYePnNUjPw6wURZluLWbCRlFQs0XGytb5B+vZZIARWX0SU1WE3SqEY
6lSM4fY5kyRcm9GtDqSjTkDZsYyST0IZPk9PxrsZzgY0tR/UGpFMkUi81M27RpXP
/qnp4LXGsEMmw6FIJHuP5/M4vpVdqNARUB+2UQP69daZ1wJ2WvRHwuln4tsWcTfl
ARWnnTJMaH+asKQo8OMLULJz4o7Qc7gDnsoEF+4GpPIIH3PFjZ5AbOv2ggcBZR+a
TKSfXfL7AbQTByRF+KOVoUiTE4VNCN3P3fJ4aW6a57aOpquBOBSvhYps7cOIM/NK
Gm2OAUTKbICuJGAKg1TgJLbBbJakV8v0u/zRqOIN/hB2TUqEfxoJYNy6nDZkLSjX
wDIs0UZCa+WiSbpd7e4WklWDsayCDIRA/J3WlPGSz7Zxi542rZcNJeh7qW2KDnYo
NFz5wEYLObp6yymRpSBtJVLlYTK877b9w2r5UWZ841QaE0L4KNEmdyg444u1Hn5u
y9Dw5vZHZb4ICWTkgAPZnBpQoedH1adr5VXly4z0hA6F8MI9+fwIJA68krWgB2rB
yD2ltB1ofRhORx2p6rXA4nOQDh8+NwgGMlv0WqQqiBnDc7o5W4Q12/YAhYZRePji
49oWhtSUcWtwNWx3b8xXLxyZCOhQRrUgfwh9WO1cokZ+35MjhszYRthu7V1BUMN2
1LS47XBjZu+qgyiuI2MvJsIh0NxZ4FpxYDAl9t5oj/59ppxmIT9x367rWgYeGkNM
T9cVnP9QSFt0zmEAQRjw9g5xMXutygXJIgKK65tVpuo7QFNtFetSiAvyyK1xBbTn
Hf2aakrATeC7hWPqYhL4AWNWa8eUqyuaO60A+NfpALPra5w2vPOKAfpJo3NxVLyh
r+9JhTEHv1dlAHC3vlOmoAzTks+Z9M8LoUucPRHrDhf7B7joOXtb4NTSMy+Rd+Ae
50O/1cZH3NLD0eJdhrDW9AcPxkRz3tzbP1tt1LRcXbIng5fVKgetEdWC/A6KLe2b
wvUTHZ98HHiHFQn10BZezpmq+xNE8ww4WqIoNdmEt4/oOoiI2WJkSRKMKYft3D6W
/9ad9yZWr8wl8o0uKoTeGS1LzeAvRJNscGhs+ivqsp7J7UdixpZskDXzeA1/ky54
xNUndnhVVw9CElTvUmr71EHEUDMDMxChs7hgNd71/I9EXf0UhcJqRAiAmXCa5v9w
JleAQtEe10rk0f/KANv3QnX7wnlmPkvHFKBQ8CpTbJIYJqDF04lNq7HThuqeZEWb
ZDgDLMgRDk8R18haOEdSb25v8V2938AI0q6drC5T1lSvQDkpm6RxaPe88U3Sx5kX
WUqO3WLEGkxmFXoJ+KVnUlqFyYRHUPcLq12N+OS7E2J6uoankjOpQnDw0zB/VLRF
CyeLZPtTfVc4Ju+nCTmi9SuxktudhdtTmRVOc90YIDns9uqHk06qEhOC3i+82rff
Ewjr8eqavp81ywHglc/DaJd3Vq5CEbnoRHfZbuN4J0jcESw+caYKWUEAFHCC4vnr
oOKUgH9wNBqpb4jeJHVB6R8lmYandWgT3s+RPCC54mKZzu/QWD8Dv6Mf4aGowPJ0
8nB+2BqUxR9hUaU5l3/VTUjx1Vh6Etf2MLVbQpy91LoYJvu8AZ8bHU8WaZAJOP16
QaDTLoXR2+omi71T7oJkPutsx/sx8VI3ZUsfZ6WZmeihPcqw3IbXwsEZcca2rz4T
W6o/pr9RmVGuyvTgFB6lwrNWFf5BjLjTG0oEtaEYx4BYK9LRgZV+bjyXv7cgIuYp
hW4jg2ABpzS9r0dxj1oGeRfYBk1nzbeh2sdUZ2Cja0Ls9Jgxc4vpf6+cYtB34Mu8
Iqa1JREz8nYEZj1MRQ/hslu41f5ZEoOWmRmfzThr6r7Lv+oh4DfeEcLoLjA0FIfI
Ls30OX1XyAF3pJIiBQyypFY5/ejFaje2xkNZbtb39JcsbOOg8G3yXekZuEVts2n3
BGZ+jw9iwTaEq+puzez4w0NxP0XJUHgd8q+bAvT/04CZ9HZNnk46dqYJyJq+a6UG
yCKbT8+tKBWgP8TB8xNBm5lMdBXgMdRE3ItgstLkTjxjJmjLnKqxc2VwId/7ICLs
qVf0ulf2XUnHhpUnJXiKLbgxk26Iz0Zx7u+Bh7cHn6ZEh+nVDl2H4/ZNR1qAuAWe
cDnoFxvqLkjPEhUuqUubgMBTNPT95x/insIVTbu8azZ8YyoBeGtvrdC+wc3DFZox
z11qxop8pMvjv2hT3C1cq/rJ4pYXxl2qsbLVa8H3jbyQhNK+t67VEx5NaCk0lQd7
xF6Uv4+0YH+bPTE5o/SWVkMKMrDDSqGJ/evw8giZsK1fzF56/szbyKMEYM9MaDRh
QiBj/cZK56csmUifaUZ0agIowDRJFifPezLSD2/kn+4b3megD/t9RiQHDen0Tqam
vwLwi6lib0e8JGOeFmQOuJKYXmf2jMKh/blsbQBastlqGdBKlAoMPme2t1PGCmal
bsoCA06zrFpXRRXEHpN1PFtPK2Y7Jutrf7osfdCOpJwjyqorsgZS1KfJk73j1fCy
r+CUpMKPp2yf3erh+KezbVezaPEbM0xcUrFTqgvM7O3Q65HdBK1hTn+FP2y9uBuy
AK1gsELEPvjJJvt/qL07isEyACLKTBcpOEbmrvbjeF2nd/slPhDSW7QWXO54f5sb
rbglEHWcaInDNKExIB0CIZm9y6vCVDPIG418hZ9yD5Ppt76H7RJthxjSKKDLsGNZ
TnKEErTbX6gODB/VTDLrf3lDgYsteP2f5KXqqKgTygZF5w3QbYn8qEzbo7VRO7wW
jzJnKlcfUg+XHSKseO/7VCh+De7hXRZH6P+cQoou2gjDYmqow0LCo/lay/2VG+eX
USADpzVMq2ZICadUVIczqRe4M4yJsnUibY5ZUmL6edwExWZVYJ1Q5/Y1rBzh9TA0
qOgSU/NpnEJSuo3cj34eRHRq0F6VzbTDqvRrr+lhWSfajU9uvo4cszcnmK2fxgWn
3kl73/XmulB8ALpVEAll0VAfNm6Y4kNm1xfTzN2bGYsjmTVsBNCguK5gXNdRxchh
kbTUsoQBUokfxgdFyOUZu5JNeh6lCHs3fW7mjfY2D3OWjnHTIePZKWFz07Hr7No6
EFw71rt5wY2KkiP35nY+qc79dx9E2AvdqNDPp1JDHmAozG9KxDPYQIcu3XPDJMoO
E/vVKqCSWDgssQuNkzirC6rA0U+dUUzZukAD1Sv6JQbnDfWpFColZXylUQZW18yg
p0wHn7sJGyv3F1ofToKy/6Vn5CqNUXHGv9KTJfpjda0kGRWwGoKF/A1+6ToSlZzd
EkF7Yv36ghtiRvEBKyG+JzwuoY7Zgvq+KSn29DteZM98isqz9pV4JMp/dKTrW9q1
n6qxibOnHeFWzvlX0VG8YGXtG+Kug/jkuZBtsMkSNdmtLuq5DRduVZncvUWeJ5IB
YBgsaZQZ+6/xzMz6lSjl01K5MS2IB9MBpexikinzTl6WmXMmULrY0zxSO3nnHMse
ja+5H5nTCcbLx5bw0he2JuICZRDtsGJL/xDXscBwhRG6XdVcApNe57qACewtw/Vy
j2tjmoJTkaYp+RHDVry2c/xIMQ9aJfvpBbHTX6gi7aRy/XDThNNNW+L/9xb0TS0X
8R7qkVRJGdehyjP/O1FCIiB+QHtF9gYkkDAzOjrYQzkKoyojyGw8Z80ORwMVnw+2
6d67Jk9ir18YXClOI+B3CZBg6n/SL1b/6vU8TkwJrGA7a3rMO0L05QEJJeKxmaV0
mAt0p0Y2QUDSop9nPnyQGY/2Gx2PqiUGLSoF1W1qbtQQoOoyaUOLPcm+bhzpOVIU
hwYq/kAear19aN5v0fryq+P6mRxhM5J9tAFsvan6sNHP7pLsFLiiAVkDPLn1riBE
`protect END_PROTECTED
