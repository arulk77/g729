`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
jHS5iSa3oDAltTeCVxFEa/Z0P24gxZq7280m7DcWd8A7Ff5CqmwSAlGQgqLXRA47
TXB5kOeWsZ8Eu3UVthgxfvoxCDiAGSP7lezvawGkY/iX9cYG2R9zz6y0IbPWMZmd
lxsc0OOkNiptKWsQ2/NIw+gH7sUmD2c5xl8cQR47xsNbgFoIXLEf4UNuKyO7uRIz
UDHw/M0YgLofgcVSKI+3Wx9xQ5snbS1pZ1XvrUKKXvQP8VzN8K6tF1hly/6/u9md
bJsmaw9nDF/glRGwc1eetIvbnVARWV8zM6OcEbJzRU+tVIePOioNBn702TPxd9A7
S2Qs07eGKdXFM6YPy8ootXOkLft2+Y9EAEX9uPpmQirFp+V4Ia18zR97CqN/gMpy
E4CsVbqAq43Wmo4hTQXTnFsR94CMaGiMJXbEkUMA/Q/VNqA9u/hC50Bvnvma5EFM
IuDE5SsOuar/X946/tQ0YQ==
`protect END_PROTECTED
