`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42//vjJamQ8HlxdzIPYyiAgVuUtJZ/Qx1J7jPtKTzRwY
YreGMoTsboqsu8/jOGKk121IndyDFdYHfe94N0TcaMWkIwrZnzYE/qrxj/2sPLFf
gtWz8AlKZ3FHhqqyrLKtPogQrKiExbnu7J5NVt71K3U957hrtFrbIgAQsRhWX1Y8
T7+AwyfVZxzcmBXX+t8u7FBP0p1wsqqScQiyQ7mX2i76wfE+RzyLv8ssMT3sDWHt
kRQClRduJYoZwr79k4DEIDF6degloU6I0K4asQDo/6dUV/v2+eXBQK7CQUIwsNEs
lNLB7Zg+yIhse3kifYbSFQ==
`protect END_PROTECTED
