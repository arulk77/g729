`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
CVynBvPxv/jyZdzGma6sPhltq2pMjVtb6CoOFIgQOMRxnnOX4GiRTi5wuaUQaE4W
Ew2bDMJUpeUKWdPp49TO27Dx66hUVcv4avF5ppL0QRvVLV+3pHGHi7BuGnMg5p/s
+dPfFh0C/AW9xOVWzs7LGV3neXv3zv6tzZMPwvXGEKfjZwUUgWw0NIpvnNhJndAv
V++C1jLRXXUe/5Ag3y1ATuiIjnVxFP/EZDXxhngvjojfYrAAIpycJw5MsEx1eN++
HBHr0z7hQEy/hlFDZ0IlGl0MhPpy/HtWj4pHjRObiwa2DzHhF/WWnSOiKERa052z
jvBqawfUO9F3A+CTQoWrX2LpjJM58yYqa9A6h+VrURJvcmAAsolalZFoeVpAMXz3
rBMkolaSTrGkgfYGSyTd8hsyjMK0GqYujM405r3oh4n+bsj/52DW+p4pwGmV9h0k
h8qqv5mpPfuDVs9U24Ymzh2lqaFQ1qTRXGbpWxMnAyfnq7pVL5aoI5UVa+eYCIve
B4Ef6egukjloUSYavlhjtBf4TPl+jyIWB09+KMdL3Wqop33S3krkUsl/GQMW3npk
yt+t+DnaHZShIJ0iD3f+3QlnLPIR24uwaj401H9BcZ2YcrLYJ/IPSuoKnb0qz7FN
sRLpIMt/IGGV4N1KG47/eqKcT5+9rYDoe3COfybPzcUdF2ILFdoIwZkb8Tihlhyr
4/1YCxOtCFenxLGJXJDihBfF4tpfqWwY/ruzTDhNwNYBwIh3NyOdgEbwLSpJF7H7
rs52uFzcwKObybsEAi6Z7Vh33IQL6nw/uoHWHHImYMJR8jBAST8/p2SPstGpHobU
QmhYS/E/Ctbc2QlcT0G1rmdCyFx+3JF+JUr4seWNzdRtJQ4+OWLH3UgucuY2T3lh
GISl5O+0blwZbuNMzvSKc1qH3i4qPycHeA5sTwgxGFkUiWiiJOrqnz+FaeWrwHHf
jG1zHtgMOa/jCtaT4Ke2YvjiVuMqkkDDSsecNP71pKgWsZZtrkqywnqtH3Qsfwia
byKunSJMwhcibBj37KPsD3xzrbS6bSBc8wGt+7ayguhOAjs2hzPd8QLXFL+IpU3/
I2Hq8XGzlx3y6tmjDfGYvfYpVYV0e2L8QfAndeRDTCxuBw1lFs7Aw5Toyb9YBWEX
yASCJdDoE6n2Zw5Av4u7ReqwDTQUqbhJfp4gvai0SOaRKB8l55opkpaAb77LDcZi
55hrbsJYzRtST9Tu9gkbnKCazXFcENExgRTuV3yTTmw2ns8VA9+R1KnzHOIBCr3E
SiGfKK3e8qaB86Rk9mie5zF9G8GWKf4ySoGJ8eDSkRQ=
`protect END_PROTECTED
