`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47mSMWeVaTjfyEYNtSX/tHBBF2HvP6feyLLE9tR3Mgw+
SIRy66PYeM5AAksPWRY6ZmnoGKLRG0MOPXxCSevEqQKuc92lwZrL+ksWas2eDtmH
OFs7zY4qr2ZY1/kWHJAvm3ynSb/Ip7K8qy3p19wRzJR6PlaGOjP1aJSsaIYqIEa1
kYCSepA2oakww3ilUjZYP2XQqPXe3fsJt9CRA/h26yc=
`protect END_PROTECTED
