`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGs6tOsG0P2u75Yco5VyVqAFC8p6fZvgGdbRhz2yJgqH
L8p2Z3Jn5py5CoEU3kKDUsQQYZcZfW7j89SRy+k8Y4YOC8zhyGZTTepBeTehGek4
vI6+YRyww2xUlG64V0shAuRapRa5mG4uK7ehxuCvGCRZLTxwAHwt6bYmRSpWiiz2
kOq1gbzZOdFUI9fbf+utVIKZdSxqJDeQee2ErMAx1dRXaIjykOH+6p6p9FIXSxF2
`protect END_PROTECTED
