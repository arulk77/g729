`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
PnvCQPATRmTaQoAJ7tdm/jT6oRf0XntShCLzUtVJ412QYJ8yPHxTq74/KMrtoXJF
TZ+iGfFfBHlJZXe9ugzUO9lgGg3jXHX2Kn7C0qs38hwPYwjAJ0wpqPDROH/tB8oe
m+rOpieGwtdqyUCPe7havBbPLbC04nRLoV1oFRloQ+DSWY0vRcNmcX+27pT8lM2p
`protect END_PROTECTED
