`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMAk48PoAWKAk5tVV6l2cqa+AQSS6TbYrwb0fP2d35DW
v96oKiWKhhQb+JCV2HuNTVk/CYxtEULhehhgi2C4CMYqYBgOVp2jA76dNHq8rCHk
ruqsDxWj82i4UmA3dTox6YNSCukbiictY85jnXix3y/b3dRmFVq70UgJ/BFdAR2D
/igMcBGiSate+CwLEn3g2+RHh4OdZdrQKgUD6NAyGCqSpO4ieAJbgq9ICj5sGycP
y/pd8R9xuQvqUwveUU5+F9LP5LQm4UE7qHs6H7lxXYEolmriIGue7Z5Em1Hz1AtO
ob9o3tUQq94CYFny2408zgaURQE0wnRwDaq/+/KP+eTgRCpIrOwT30bGT8E22HBO
zTRziT0fHMK7PcDQnPiuGR+ZFc7Dk1DqSjkfExqLPjIL0fEVQnUsc+ExnrHogY4x
RKyQMY1tjjK32Hu783+B+DILaivS/tNtopH/LBuIqQJ4pHn/VCLyJ2F7pthzRguY
8ma1rUtTtuQjsw2HL05ZT4X/rFAhC4ecYociJuz0oqOR3VSTbvh7LkDvKd35h500
`protect END_PROTECTED
