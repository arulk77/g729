`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKgNmSId6K3MHkYqcQsLEtB6bfEBWESnr+7frMkTt22T
BygVRWs85YZF1Mh0oEU5EP0diW0cMJG0keoi9M1cZkrrLAyeifqZn1tpGqyoMHKs
yZ8JILRiGWRubyJLZKBO0XPR+uFF4nF5Ree8zlzrVDkNQqkYMo7TT2LMKwRuXACw
usyaOietUSshmV67HfbfolT9YutFMY4Z7oKkjNFuxVeClcYbidvLBW6c9LgsH0W8
`protect END_PROTECTED
