`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCD4aauIq+zXy+fcjs3Cw2sJAbgfMYyEZ90YB+AOevJB
ZJ9/+sfdSGxGUwrRDdoJhGbEWsinBVzGjwtE706hiZBHWjj0LI9oKZUdnFZk9GKo
q3Jde++nR0qk78IKrQqle4EX0RmpY2DtynHthkILxSwFvXEj0bO78C2Amv2eseWx
AZUqHz+9H4ID5ehggXmUxA2Ed+h72612ymNN+plcE17j6UdFTj7r37gXrCEx0W9o
8P5DXfQoCZIoVxzn9YTD0M5OPVP4KWMdRa7b6STbhVivDFqC8bgiPRYeQMiWFkRE
dNyS57DzNdSkP1H/9VKXSQ==
`protect END_PROTECTED
