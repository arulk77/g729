`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
8N9okeFYIogwG3lIe+pvlPmUOV41IS3pmP3kMgU6mN2oVtgyvFi6tcbsRZyZ9IjI
ky8N2xv3JZHmUkbQfcvhTX7tdlKcM4zFtqw3vmYs5to2ui8JNBIeRxk1hxi2llj3
SIxIAYMqlK/e9mkkBIu+abA+9U44A04gnq18nvlDe1VQmzBxFSPiS3S9gOExgTzs
cd3CSX4vo1Idm68XVWWS/cDAp3y+bKSxglO/oVBNu2W0D+PqSYi635jUTegiiqWA
W9/5W/PDORQCzcklg5ESzobpvpdW06z+kNgYLnBfyMmTU0p+56O7WR3U/dLtaMEZ
zjDtxSfKI8N4EVES6ajK+Xw2HDobPiTFZHRit+ro4a0=
`protect END_PROTECTED
