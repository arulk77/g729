`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
wDSceBKhzaNnzC+VZH3qDAB1yu93oX+y/ORhvrChElaxtdgsO28QDKktup3MHyWi
9D8QiukuR/V3cbtjDMfjVyXDIgRgYlMqegLIKl3LZqYukEmGx2yOGUnhyW6mhnJz
alN3ngScEbDkCuObGdLZr/XDufQWDhJUHaBa1N70mnul3XyWLjwvVXCdVo7pCBrI
mewK3qIfeBErLq1hT42852eXtVlSO8/E9i0b788N1G1Nv+O1OizXQRX3Pc8l852/
IMTG46IVoD2y4KzmfSc2YmOBW6dReyYfpRzlzim7DmRdXEgJvZM88vxnybdz7waa
COUYgjkUHj/7WCWR1ELT3T5HtI//0aY4waz42x/I+2DkdRT3Y7Xz2b/WJTmFFtgE
cGyZREQEcT0QI1LfoFDOO1pHnWfdrJzhOBuAE3EcyOga1eQW0WvbKV+BE7iFbUmh
Z1qtMULZUiGX8ubjodsjcW2YIkismELvDIkPNkyZ3dWSFHu/0VbusvbOUkMtxDSA
pTDDxDVz+l1OOpj9/S3nPQ==
`protect END_PROTECTED
