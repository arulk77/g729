`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wkvlIEDoaStOrMe/QW7iWiYN5DC3SINJLSvjq4JpNSA
UPmKboVtMmNAtLjZIJG76DfL9MtBiPtKhgXmRcR8PZX1b/fBQmr9LDVAMr3+/jsW
Z2MbNrIAKqIPoTzooHFCfaTV0JIiDUe7oM5pJeQPZdX6PThPSt4VbFqU5LZntsf3
RaCfa+cDJd0844D88saYZgV/kCOHQh8xuYnCG4Bq3oioLyjibYcKF6AHBzc7sxqS
XfR0bumfO62pUsQyYQALENlpRQ1AlRz/O55Y12RSkpi+rDKKsbiiTK7Hl4wZo3qd
kUf3XnkKWPZ57XjLNyuL2dCANHTltoJDzgtxoylafWz6hqvXK6MYQopbHXrySVzg
kRmadjw6K7sAnPopfrRIYTBwcXLIv37KAk1MXMIuPAiLjcb7viQ2fiYCqsdV4nZZ
caOk6V2S3jKsocW8goLavEAPIpmQse4h1sZgM39uIG08ZmeUWRJrVqvXKJ0NpPvf
`protect END_PROTECTED
