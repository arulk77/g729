`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNobg/3DK2qfS0NJ0XgOM3eNaqNmAdwDDdOKBFlRJ/Sz
GPkeSRIf8mSSgvFk3tndPz9XGGbX09oZfgbRhQBl6xnDoKxSbYBaOL4Vd/kbhE0O
qRQYO4IxL0sj2vTmUQQUbpFpUGjvqxT5sggrPE4PbRgmIENFeyUhn98jSCV0VL8A
yO/0SXqQO6xXYEDhWqdYm4ZrfkcShZXt/yMxyTbZhNZyCgu4nl/v9w+LigSeWn3f
SsYr2FoEyR/2MrrpKbi+bQ==
`protect END_PROTECTED
