`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
llAYEjQJaIWeSVV8rEd++4Gj51pr+y2osVJdORI2G74DLNU9uZsHZrdgaqGlQ5vd
N0Z70ppNj9ZcjCSIJk8Vy8S4a8DoBtVwemv3LIAU2JI+zyYXeRY+2ZbvQldkrUsO
N/zgxRjqFYz6A8J5bXcaRV/oQnTYzL982KaI9hMWiO6tLxy59tzODzoHdxP4LvDj
XjjwsDzMk8pTdrM7lUEkoFzNyxNZ6eq1womnVnWcG4aFNNv9GCarlJW+LE+014hw
f8uLxUoDC7+AjjVBn+Kz1RQ2cu0Po8B3Z3FGod5veOat3HyNkEWcm3O1tFQWLJQw
fVp60prn+ujq7U+MVXR092kkEnaQACa5Cfj/zO2eJUYb4TC52CMT6pc8E11xzFj7
if7NUhIm7onPcBBfTBXW/1TnNZ+AzmNfbqi6Os3Bme4XjH9NUQeMHhBSAihmGDcv
ke9nEqnAaR3vb3dap+bjL0uFrUppIgRmWpmACYvGB/BrOMwtF2Cw2WylaZT8pOFB
x7SWjZ3WkAeWNL42LSkl3oi4fm6JJBoBdIGoDa8lfF7sK9pKyf8rRBlv0XV5J52e
jOfzmsSixxfQ/0G7fOUGpOCRj6C025r2VJtkxJ69p+4Enri4aR9fi+iagqvoQ/8w
f2MVVjyTlhM5H4Qlly6JcrQvAqWehfNwQ6JFwqyn4tD1mmM1/qnz9BKQwnTmToLw
jLrxzA/aLOInXsZsV7omb4DZ/75FY3naJXR5VYyTdzUziqvGiNyj1IpAkLqoWIjc
PaK1me6ziQGCpmqd9PhXdZzEU26cwz5sYCH7YkJ+cmFvYBh3FP6euy55C7ugphvn
bXBTrwLiN/IdbM3Ddivh67d9fLYYyBKFqTuFtbYYMZ7bFx2RBFUIZozpcoQKgC/r
FDKK+1+JGvamyCL7tJXYd5xNO5JvJ6r2OHMXiEX/VX+a/OcbRlYivdA3QV4hOsze
WRfYaYgY8Ptx9/dsW3P+O+OAVgdiEXJxp05xWa4e080av9ezB0H041NZQsQJlH+s
YE0vhLZgtjQT7UoTr/eefRDypiTzg3I2BUhojdoGVKk2WrY++dYj4jYKRMnK3XUx
UNNEWrxATOTzXqk3Y421fuDQWOIOVFN053+XUwLNqTLlSzrxodjiXKtMPbV24QhT
cr3ypraje5iV+UV0fhHaMn+9IlpACh2IRPnJicnoEeY8mqPqUvo6/2NHcYMhCNQg
tNPRx9O8ITjbZiXYAj/PWmS3cY73XEI92vUUHSf6iY9IidvC8PMhkyBve+KmJNdp
SApEog8i86dLHlQ/mJWyTxPO4h0Mn1vheCVprYaTFFJjGzfk20XeWkDDFpOeVcFr
fM2c0ORI/DjfB+e6hVdYg73BoQotJGuL2R72kT3Dg4jRssAR9BIYMASxwuirGgag
jFXzAXk9RJujvjeKPrSoJrRC3i/7/bm7UmqGEF5GhQUiH76cIFY7hDxUEWVTfuW9
89PJB4aRKtjEX7A2rEE/GZ6WNvDtlx1c+95X9fCKxuXs0GNnzSqzOJ55qhyTufoS
gOsLL/Gos77eOddqJgb3UTIaP1uUsZVHdCvi4MTOjPKv3JWFr+R0rs7yDJ8TVIu1
mk86ObGTIqiihabmKL50sd0ezPJIUN9jK6fXmiPuefkTVPwnJUzMUl5hFh0Eyr4+
nXW9iC+hdbz9rglDHWOcVUJ8xIHu7xF3IgrS0uSivTC052/YSd7dx6NRQi7E2OW+
gfjGMtaWWFPOxOx23ibbi/88ECJjmAX9aeJ/9KjnT1Sl0ld8A+2MB/Bm66FJprgU
bXO64GzCpaS9WMPUu0jj+VslVTcVeuPezvoU2TOliRKdQc68q2CeHLlarg35tzv9
DxcslO+HV01Ruw09jP8yc8EpOVzHqofctanImhfUL4neHSXVdFEL/3knoNFuRDEr
K/WjfGE5y+NEFylMj/ZNPb+LwFqAQqPTO7vMVU6jtZmxGaB2Pm5xX8+fcfJ41mGo
ZGXQY+YT1qBSqJW8jvdQcknddwFdIBrmArOCAvtLa2dXemmdPFngOsrsOGdYMBnX
bDwjKGucRlO5FjyNU98BbEGgmvAFlRY+7w06adbOFasyPrkfqpcK5a1sIqpoUQnV
8Bl3qWxEeAm2qXJkVQ2NZxfYwyBnAPz91OWhW9guF70oBw4yovmjth20ftqB4fQl
7KeJsaHqsYtYFzaeevKoDjzqezFrer55h1PYn3CMqAIWmhEQ8bAV8VqWOr+JCW5Y
kYGJiNaeAATwkQ+pjtzQbLbY+etpma1EbTk+zqDBkl9DIxyzDKCzvpe55czPJ6FO
JHOTLeHD9LE6meyyWIKDjVSto3WoqnurXw8dDrZiXrFgKPebrfFzCUqY3lRkXsRh
HEh26mtk/0FytxerezbodRsP3XXOLLpOsX+5embdZR+cmAuQ6C11ACa6eMvitJDs
1oGNuJwRdDzeWAYw9FIJRa3ay/qz/zYATaKb+TWvxIG/rW3oi+eyCnMfsR19Y1mg
4clxb1uSB3nVElOJ18/kCUwL8CcEOFqobgxnIts3VwnYECMTze+9WFpm6dRKcwip
PSGG/WupoC5/7ZPimHQGesJuYmPdRs0SFhprQ3sOPs8C0T6qLjIFKlTNue29fkIO
aqyFxKJW8PQGMRaoXlE2r4IgoUxVVbCAfoRmLwzo0P8HtnA50yFmm+D4Zumrlyho
XKVuVB7qWtETIJeyA1zJNQthm9ZGLpfA/txy4x7F2XeTm4RpHUvcA/xOHsxVQzBA
YxZnisGZH1O4VsGwEBCXFWMsNOhtda4QdbGYG3ZuA6DtV4GLhwEEIyGZWA1vpcxt
5yLItJ62Hx55OSRsysFDH+NRxoQE2g1rqCKad/fQu8nNN2m+0puL+vBPPH4zQMw0
/ME+g0Cditdx2crWBPdW9M5LLTH1Rm8v8zgpIYtrkWpyMcc2sudi/cGgMvTuTwot
HX8uGYY8Fh02S+V3bc392QqQxiTWxJc2iJ/dV9MN8ZLkzumeDuurHbwLUYiI6p5W
Biw6M6fNuVH0tcuJDq7sN9k6FDvvl7wR6RB6oJlrewYzQtHV3KDZpgNUzkHxVD2X
H1Mpqyde+wHixaVDF/f7+Qyl+xpvI6+XQ9nZNarw4rVJHs+CbXsfl83GmQzR/zei
AoaDfVBcKFOLDOOEzUieOol8j9dXCZgGuxVac2O0P322II3Us4+VEhm0rZEevLtT
Lktl4yHN+rnkQiJfeKvjtZ2XYWUo8nG2TVNOA5e7Y5p0V3n7pCabY0XEMDJcMiIK
3jhlv1tyS/oZdYyKXe/wp08gGbxM1jccMpxk+S07CCbgpObdg+3bboCb1fQZMN9u
Yx8zjrDCUzmewVLJPjivBzyrwLiDAnYsTSM1wlb1QD8fzXHLMo0u8VUU9KSf11Jk
rPhPmw1sx3hq5YLHm/lfrEAyUaeXXB6AlBzIxBpEePzomio1dfwH+1Q4tGfhFqM3
kgSNBYAbgoU8WimNFmpERAgHnYpmAOPNsPotzVSJA+AQCikWjy3/q6WYl54qy3eA
fchTB+lN4PKBKPtdZu+kEorOZsGID19bqVto6KYatoIhxmyZcS0YSg3z9uo3HAlU
CGqZ03UGYTFNcuMgQiiucq1A3mqAcHKsAdt7IBhV0TwjKbOSxZEEoIuIE8CvRbRu
Py3rekVIqBDN+jkXIr+Zt0txqt9KkwkYrZ5BrXqlU10c5KFuSgg++Gf7fRG8YDoI
+hSttERfyHRWrptyJAqbryh4HV9VioytO3Gee5dZUjaKPzfm6VqA4ngyD9Y+a+qk
+WQS8QHUz0+E/ATaBnTUkGTzJJuFlGJOR8pWFSOCXicqkihXFYnYWYSSXYB0eXxx
mjqBS2CZfTZdahXuaNQgkN+PYal1a5Tu3vVj7nBNLiPlUKiCpTCTurSXe9HN8Z7N
cE4wFFzvINAp4+RvEHTsJRtk+2lRpubmAvvF4iBFCkhl510cDzF+DdSmlLhN1VEi
Qv6VCqHKJSyFpav7goKMyTe00W7pPEfCLTYj3m4jptYaQOOAjamqyeZFeHeDg/wF
i8jQwViXL4wIUYrA6O+TVu4Ew/sO4qU1YZKsVVCUVaOUBCBkTMdMDYMWwRT7Mw71
YJxfLmCZE30Yrwhs2F2nMC36sUUSJadM4CCtqQigq1oDcTvURoqjPza6gszV37oi
jxC1P6k17vWISAJj6Gdk6/t3cbZcz6rsDIGiicjx4Xr6Y0rLft/01cKzTZXE8J19
K/bS8kWGTr9TUMztkYkfSiDYadPZjBwIMm3LkwzQ4EGL/+5GkI+U6U4HRXltbtLK
jmQ5L2TqdVP4rWCo6kP+jkz5XgaqEVzM/HNe6iVHS9TfQMinKLckmIE0S+8hHoSB
bGyKnpnfjfkaRFCnF3XFucGNkmiRt7jU99nK1yIvuRMXf6Ops7tVtarqc/qRl1qe
6sLlQNBLbGCv9aaQAAPkfPjzFLofZyfKCesL87CBnYi3z9Qosnmk3v2lp4z0K2iT
5SDKnUkQYSFUGKIRBllhe5yiHgT8HI/09rSayHu0IGFpfHCkLjn/KkAkqWIpsbDz
Ekf2+HlqUN3K9ET8L9r6W7WYZA7LXbXOFaHQOFAy+q4IhxIi38/ZG57rF7jS5GAZ
qDtA5ca+OV+k3XiN+xZK1MKqJR0zVfzS6cnXzzebOpomjHg2pgCm2Ie6noUjX5m8
b5qxDtcbnx7yRbSZSLSe9ENVQDxmxSd5el7dSoIx1d84uw8Kcx7K3D/xMRhHa0Jd
z58MOwCYol306fagRbDQxyrFeIi+F/NR2PYxXNPbB/lZT5wt/OmBLiZOCBYeY5HZ
vuByI0B9LhC52nRI38yWjGSFs9fcBB0g6XLEP2la0eKYPQudz89XDzbPwe/41dPL
07PJdYs1fK2gqFamCAyKf20jSyTr3hUvPfZoMEW/JVHJeOuTpE7WaVPdWz83XBK+
+KZAsA6ZZXsOwE+fAIcZ/OUM6iojISXSqIimz412aFO1amyNtXjBl4ETvIiJJYGH
tkvzreDMqheZg88E10MxmiQJAH7gSvGzWyFSFTbx1MKqeyoxOoZQUB5hUQUR3e5+
fDJ6xfzMJ6u16+b4BrQTVqzlqKDaFNijlkfmLx/1skVftxBCVFoV+QmxPdpGiFjN
S3x1dAqFDyDGy9rC4iSVZX3e4sTndDHolQI49kF2HE0l9aEyNdcI0sstKddOEpKd
dSBKclFGGQ1QOF5zCpuL9So2fF3zoFzU0iw1GW7aiPmEc6XqyroKnzWitzkhe9H8
5XJy3WBtMu1MmgO/u12gbmYApdM4gBaW6NqwmiqSSWMb9pMRCkkw0vBUMZTc8l/a
7QnKWELOyeOhEWoeuGQSICz2ZrgVHusnS7p0PKR3VkIesRCm2fI9WkF1NT0py5i6
I1Xh6Ajr9yMlgppdPBgfxe5DHXN6xH8JfE5gqHrtkUphwMGO0YTPkdv6vBBOTZqn
9z1v3GikGz/6G4KVVg5u5sfT3KHfp1h/vuDZCF1Ig9jjPLMaYDeTPyaGX9astcrN
4ChO+bZXXfHF80dbnup5PNtMv0OkU+fWAzieB3s3NycF5QL2dwDAqoPaWZzw5ryv
sSS5mdw3PlmHanm7O4ShN1JSoeX3Z8sEJYBB67irQYywXDSI4yN3WgRkmZ0WbBUs
k2uRTL4Uf1+hECaDN7gkpSwX5yJNAgzff3TjhdwpuaLV7NX/oQzxVmnwGe2Ig+7H
ESl8sp0PzbHhfyggsdgth2bdhM7PYQf1kLu4wBEf0imK3M4IRqIiuT5f78q/Z0tl
U43MD1CJzxU43yvV6TkwbEkjMsUa6G9xIKQqP5R2P2krUzp22mqeoEyiJvf8O8QC
2ZsUbTv6lXGjQ6CXFFvCZZ2bpKJf1cJ5goOPyXfXC2xwzTWpapNOaYqdYTaFKWOW
z9DWOmaCccBzn45FIYl2Qa9qbTnFhk1mBzK47FXMRFQxBxfEOvEi30+ZUKxgCYZd
aNrti3JdPR5CYPZfcEBwymyIMEPEPv64xN3yWDool5Ey7Uwr+8lGYkEQUQEzQJkS
deJKUvfFV7wV/XgiM9iBhvRYHwbiCU2H6Ea6hqhsQ/4FYFcVNnRtpRjrj7P8wY/z
4Ki1GX+0mIO61QOT6/zlp9ci3bZblZHQ+5I5Kxj4S2sb0IhIVI+4nePHy3tllGHC
5twkFCg8fNnsoJAlILzaE/IMP1Ru50hdJ54i5Aj2k3C3VAviPj5iE5Dqers0pfQT
unUbYp1iD8a7xwOQ7wJWzRdvYmt/ISEsPEP/EQ9Zi5HNIgj//0kVSgb51urgcNDv
wZG/Xz5RO5HktemqzWQlNAV8XntFqtuTNw/h5q93X7y+EUMAXCXyCwVrF60oFf5i
A6xpvi/heTdC0Tm5YciahW6UfVsQlq0Id7NHi0jg9FlEY13niKTe3ppsUVkKaphE
YJTIFK+WidYwOUXC/0QLi6QmQdBwecaB2msKOtBnxihQ8zDIgqwEb0gq8KnKyB5V
xKLTJxBmKSSSF5lD3Eh7+w44DWyVbun49MiOA5UQ+QfE0rGa/u28T09v2ob81USL
dTugXN1HUYnesq+e4INBiP2mXOxrriWMr0V54mWV540OkgPKuvg7QofB/jzmL4x1
J4C136+5qwtoyPwDCO2lzQpTFJmA1cLiO1L7/SaHJakhqaWWE0zuXYtjutNaThar
M7vkqxgxsjL+WlE2Y7ke9Jg/gMU3NtKzuFixhFDkqq6sIlKr2Gyxn6YBmRBk+CZ7
i9ezb+ZOzt51rMTil6s4oifP+YrBfMNmi/c/0U2HFoMrsKrDRnM3oL4pWx1aa9tJ
T/0XptpqJ67Ueliq4+V4RfDhcUdq4sD46L7QrrWYzKCOBuENM2ye4xUK7jBo0VHY
VXDdiHjSaw+Wsx7qb26+V/34RXXsVlQ0i63sclSjwp3xHOWoXovBvl2Jwb7DTDeJ
jh38qEzGtkGy4wOvAe/duUBr+0iEi6Wvo7jljkve3uPzOhIMg4VCP7lYCenJzmTD
hEXAarnkG9aGTtJbeAtuhPctYTCf7+viR2JryPNmfTbczAkf3kHDhaOeLEXr4i5R
QY2tXeNot5t32jftqEsT+iI9iaLTAE5UHg9gQO7fiUT3GbqOHfdtxpXles+N2ag3
ynuvXjtOOOsM6AiZCqwpbh5kKr2YqUD93TEumNLNIw22j/8yNlb0HpcT2V0/BfXd
+6ughHPgF9b3lthXsxDmlrSDq4Z6MHLxceYxLMICGqYgNmIOIIjS0j9O6XFeBhQa
AbpzKOu9SW3X99RvQR7h8V2QM385+HpDJh0OarTNpIoSXLB39C8XFrJc/3Kd5ixf
VqQ82ndvfsaHMQu8Mdl1kc7r/Gof3mNtW/+kAA3mZp8xlvGQzMlqHUlN7vTTAeHf
IqEQEqEsAYo5MZgKzPFLMBSTd5l9uVHeMnrZxLaBnoT01SUxP/t33yinGRuVcyU8
c4xWW9rrlrCwsoA0mAzDc81t54zYQGKCkCEqI5/UzKAzml0D8xCDJ1ieK7pX2Q0C
1ZPn8UbOBnEaRaZNpSyB5N3SIjtdkZFhOfSOAWVvja0MZ95Upf6hXfgfRJqLN5qo
J0JUyPe2CfC55Hdft4NgGr3rlbtbY1/WQP59mEinRrgSXHK54GbZ4bmEq2u+4GUl
rygjYY2ZYP5TjRii7tmX4m6giuf+NZnqugp4n4In5rPOCfQYgex2Jas2jUKofYB/
esiBcSnlb4ik8a5N64/n4Wsh+PgqNMqCS/ZGWBkWyZ3hmGwqcnyyblsMdLN776Pr
QpLMhSH22RLi0E4m9Dx1KjuWPdfyGTeiSghaMMXZB6ufvWktEhHqadfe28xGFx0P
ZOliJDZRrNdcTfcCE1jcOm68K8pcoU3jkSBge27e9MKxxcxKwYeJSwFbA2XcllGd
WsSzOqENEGA8iNGqNQiq1mpfeaBsWqmjDFl19WDAyxXGFy4DS9IP63VzfZvzUGBK
dGMM8W7f5DGRdp32iweL0KIWVS4Cu5pJ7wT2cSjKGX4GNy//nXcS0HEzrkxuK41u
S3obC/fW74Gk1FRmahjB0zR9L4d6crBZUVceneTpmIEgAwX+gLcb99EdxeTO9Lmo
EqjpCUo5s9GgvCXtglktNWlWyQp1x+zAQYhLEyxssKYHJbzrNHrG4soVrKgGF/0j
kIA85hJdJOdew+oQXYmJCbucidU3tfzUt5BMaAFcZyROysgRkgEnKVsnrAiitBVP
G/GTyQN8aSSVfDgA3h6yM2MsPdUGcbI0fa1tWL0qDzqg4IeqYboH9eRHWZ04nvnL
nHAaRyQq9F+rUyuq+zA8mn4yUFqwO4uxz9bQReyN87knAy3caaFMHXebdRobFu+n
5vjHg+iT8DzYuqR9M5FtATCPMFpCYPFbbqCBqwozYrnouvuRD6dQSrxVofyNJRYQ
iiWcwyoxkDvO3Km2muSDzmSUrqaSTHkL6YSqGbSP9ifsbBu5+xFBcH23i0YJxmsl
TCshcQ+8QqzB+UM1iutnCrt1eSCRdUaqF650vuAeD3RdpbO+pqdTlDh6Vs9xcxKX
PcIxQuJkeRmdgB9gCm8mFXqepsFCwx3phDH/f1W8R3BV8vo7RSRmwYhQH6j4i3Pv
9KhHt93hzzzO5z9hwPQbQSK4VKBRfgA+mxsbm0Set7eSWPu92cFJqB1WWhQPaTmo
lGrcIknPMtuYsClLt2wkTQPXfBrdcY4CxjHAnHciJIsh4zS21vt7+ICJAT7uvDP9
sVrsTQU27RkM9vlJqBcgvdJDra/F1opig65mVVoq2O/4LCdpBTo7Z3Qgovf3ryEb
kqod/8faFikNSdMbg7+hvqhg8CILMnEJgxIW0vWh8+7F0ZRdk75bdRUUR315prPe
wE2RigEbk8CIPZbT0Z9B2nOBdBytGP92V/ImqRxgds6fLFO/ZwQeFhvY7umUv4Zj
c/hX9/fauNk/5YrPyajTO8qbWkheqLm3PC5m46aWo8s3aaL31vkfKS8zZdwcK0zS
NGy2VLMQo2rNVEtRJdLQmZ0oZl3enBx4+gjG4GqFKzw0EjRfpSn2a7YFWfmDeIlE
CMI53c9y+slWSlqOVqwgGkAnYY9Z0z1r7pCbstqmmpNYiVfi9SCKg48s6CWDBJBJ
MPBQSBm14Z1Nyu2H7lSfxLyBidWzwZ7JXQBHSWEdp+z9cNZjF7o+CANipNBeUAze
6eWXZpqCH6dye5Wz216ihP516k0ms/sgpoERh5UmOHzv+2gbefCuk86ZaiWmMsYJ
ZMLjIgfzkAOpgDiwGIDXXIZF9E2Sr2fzJBE71wdVCRLPciWayTzk7uyWOPQYylna
M3c6y3cYPgs29WENld14bj9B4/8KySz74ArAU5CVeOwFECVOfXq+mEATeFg1ZIc3
4VG6f50/HZze9fcG+BhuriQP46egTEL7RnJBDl67DjylTnQUk37k4jJEDYyopTgf
AyBJo6wqXcc4T5aY6/hSEADg4toMn2S2p7VZb0E/rDbxvOkBVQjEP8gPXJFO1b7b
j5LPl9W88odaUYXfHAXfT/Zb23gvA8zYneOki7Q7xmJTIBxPBMM0wxrl5IWMj8sI
uH9KtGGq9Qa09v+jRrGP3ZxAuu21I7V5l1LJFmsLW9+FmrliknbWDrsYm1Stmr0R
V+uHc32E9LRZR8nC06yUoAQMlkAtAGlx5I+SfxqGHXUcBF8aWOPrQyqIaeQtPB5A
k8qhJ7ID643RCrci9vGNXsljxJKjELfMKPm5eAnazJG+Z0iaWkHkf2vhworO0yiq
nzywAEXonRGSDdoPNmHK4BUBqgYcEygYwA7OPr+augHykz5Mapy7quZCcHa/vbIQ
Kjs2VxiSzZykAgwegoYMj0BSsH/iUeIiXUDq6zQ154or667gHzVRwrz2vY3xnYi4
t0rS39Fo9t+wP8QkHRZWaDcYuS2CbfxbkZzyCtfvucBJb7GtQmyxaKMb+ql76lOA
+VV/RxuyScTtdQALAHiQWAA5LLFrzLfPk1jlHUgogjJWDubGSG3K0D9qmlxnH2Vj
a+R4KizivorG0dhoHmY2yJwOnqq5PCCYZBN8HAgKuHJZSux68bmDOMStI/tGdNLD
gfA0kkismLC0HnFOH8hzvLxAiO/NMmPfEjqIV9dGbBEivhk2K2GErYsh0aehILPm
vwt5JPJcaiRt4/E0+T/nSWS1SqIld+cw5wG7cYH9aYhA1fiihOKSwHo7km70A+0a
dFmzICEnIKPq/KsJwaQc4bAnY5d9crt5hCW+4dQnxzNNZVrGsGwU/9pC0sKnSke/
gcRtHfn8QwDr343k1My0Y/pDGTiRdWoLMH6VzjW+ZMvGNg6s2l91+UJwDEvZ8BWx
oPv8y5nD7mHJNvZxIIdPm/IYLYC5K4FXDL0t0IGotZDvliYqU3CcnOTugcC8Hjnz
jh2eqfg2Aj3xOjpUvSD9ejYB1uG/decWlYeRvfIYNm82PM8de/LqoI0fjvyIwegt
KlUVEOfBeiPnrtIDSOrLxpTDmoWwDx8DVvmSFM1uxPe1PU7A8aQ7/RFuWiUDtwqq
JaDJmjSajZCyivJ8S4wl89SpNHUj/kMnY4oUw1UZgHOr4lrkzR12qT2fTXHRMogF
+RHF4stQ/1j21mz7YyhNaszLe2uSfExqsjcm9t37ZXdbquir+oAiJ0PuoiicnWaV
1/sw8/h4Z5h2sM44YV+pXt1MOdkJkmyy3bVMW6ZGku0PluqqKZfPSzJfHFdo++Tr
PnLNxuQatbba/QiRetOrR33h42AFnpn+LieR0RC8vaAriVrOj3pyC19xkpsIINNz
sQF8OYNmXrj+zkQ82Z6JWX+H9bFcb/V4VDExaHW659Clut501QaIefx4DxWB7Xkm
Tqe73OfG5pEWee2bomipWG8hMPgy8cXfhmcTWrq0lsbdz76Ib1o52X6pJvTstYfq
mls1CvtdLfPo8j/5EvlZRlvMHwO5YB6VT39f+S/gCNbGsBSFDpNiZR35vVxMxM41
PmwFiQoUvofguWhNCXO1j69UbB18V0wt7u7k88fxGMQ3XSEbUTSFHuK1coC0OnIq
PO1vDxIwIF0TJ7I5wXYSlFZrDVWpNrSBGpOmErEf3pG9qhTH/mjzSQpoAGRvOcT3
SgsMY49XrCnpe304GD/hlPMK+pKB/h7izjbkO7vceRDVQ1x6EoYXLE4qobWi5nrt
kbRo3aWnsMERKavmGuovNMEF8d+a7TTsIk0PRY6XTtHu1pl/NQR32mlkrcjrd6eF
Bc81iSraObbcTR8/huy3w3fWcR2JvuF7GPaua2Biqmqr+mSD7GVOoStHuM7QliNi
4i6fRwMvNyjw6IBtXK5n4jSqXnnseVeZqX1W30bnDtDAhBpNdFVsyEblwKqjWAMw
w6pq3hknMUbpxMhPQKE7cJsYdcu6b+6r2mTXW3u/tOon4ODI0um5+EfGbkxn4d27
E6KBPYm0Ei0uwD6M9Fbh+tuNq9wJYZuJlwuIkFkqUAlJiI4qEqldVhbr4Xx4F1Sh
h6t3dRF8iUEzbD3+pCWVXZGF9JVj3qyGzbdvyCs5NB5aVEy9KCDrQaE6ue4KWafC
RkOKe6dXTpKL8HxJIWudQ2Li0s5IgHyNjVDu/Ho9CqTSxW9E7wi08yLKgAO6sybR
kCIZ1N7lMveBMaydk75/pnvjKW6NJpWpPFGx46YnGtBXZMQauzHH6nMKmLEPRgqI
dYKDGJ9tQcqlzFoGD8mQNDvtLNANn0gp4CU2mV3YMl7ymWhuF0pViPGJXchI2ZTu
7hBnfJHxH6d5zyB+OLHu0MoNULmt5HTR+t6WOUYBwmKwKbU/xu6M9C/oNP9rQjMI
+VB+vFaMvEIRezk6ofyZQUl8IBh7o4r42uyEJJ/+9i4O2uEOAbTv7lH8AoDSZ+/3
XFUgtyUlgqgNanE0R/5HibKwceoJsvJUSnDuU6CqaRS8vu6Lj4nFdJTejEAqeSlh
4Javs71c2QIG2lrf1r+Pl+K59H1XWjMatiZ1zO/b/dnxR7IzWY0GhmF0AKc2XWKR
9BZx2JhWTQFzsMFdHb/nRL8/KNrfwHBkDvSHD+t8cPZeeGCIgBY6kKpwDcNFDrgT
AMB538LjK81BpGLkPiEJHbMS/qmZUcF2NhkeJpgrgkcc9/2QR1sNNSHy2AgifV29
YEX+iJNA42FVt6z6F5dIlS9K9b+tSe7zmyxsmfHWCCcJtcvJr96TfGcH8ZKiNtA+
nr3VcJA+zWZgOTsmZu0m01mJCsLGyo7aGqz2IIM41PBuK2f7cdbo7/ZgExhtUASJ
7RLpPJWiPGHcd08tE0531fEeaZ+JVK4oiD1tlYGejz0ttdicKtCOFhBy7/5uhwDa
H/MNrQZpA6UGCZwg3RT1Zfnmg4Bh348vt+U4fz7xs1JS+7tfVNe7LcOOtzN5DSWQ
jmE82JUbWV3baIhmO9DJ0Jb7gNGqbexCL7vAYqu2maVmCIIzh7Se7TWxjTWgHpRN
xS5viATFXzOeVLhS8++bQHCu8dlvWFRYspkYCLczFxrPq3lFzXEOFuhQy5YkkbaZ
agAcgdkZJ/R39J5Q9nV7XzBCjsMmjRbcIKJIANsukSg=
`protect END_PROTECTED
