`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41szd8dtCqWo0sJwzZKdM/pnOhUSRrV8Gunoc+5eeoU4
tAfMimvoYbejXzL3gsWyHwsWN+EYJFq2JUgaj5/HpwlWSm+7N7t/p2DuVZNF2R7q
dnkvrr6Cj48WQEfxmWL3XIxEm5M5boix57eFo3/fucPjC94+qKLO5eec75KKTmxn
O18A5CSDk2RbD7O2zY3B9ek2fVJJ5ngKzR1kPEgx+XCKr5kKuL4q21yPiijzxSY+
9R5AnDMzXZMCG7z7lV3k+MaqQQlCOUS1qpqbjTcd/Tg=
`protect END_PROTECTED
