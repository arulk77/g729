`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
zYVqJUZxw01bZ6x9Nfon8Ge84I3KkeUovALNAzE/feTmi7S8DL4HJLY0GeuhLyzD
fPSK7t/w221jr7sd72b25W+p/eU2X7cEv7ldK/j9B4SLw6RR5bC7gaf6DqlwD1gs
ia1qp7P08WLDJlr18X5r56nLEKDHXAQ/jJYIOnYYeT9IN0vuXhNEVhHwBlF+UiDV
BpGvvVwLpN4bWMowrhgMWbmRs4G+pX25EC1+2FyR/9xOKAF9eDtW6c0Br9uy0UzU
Rm8PPrMAei1gXJdNKqx1/rkdhqgV4ayUXWMkZ9uSh5esc/WVXLxMap3utgmDYVX6
U4SULDLmbqvz7tEH3WRSMbhp1Rc2RLZo86v1JDCHK2g1tPiiKo6nd35NnL4cQiq8
m7j3PabA3FmdKuwHvTfIieIuCC00N6feXyMC9TSHgFA=
`protect END_PROTECTED
