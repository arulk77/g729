`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
0RlSXB6g0aAk9+UA8L9XgbwO4ZtZRu69nyQ6mKzbp/73+mgENCqTq4QIi4gSt7c4
VSqdc2GP+uunGzGVzoh/3jiSqxjRzfKw/vS5CmVxvSlLmAKBBxNSGhPXlEb0X9Z6
Es0cohbb+1k2VWI99HlpWlM6g/VrQwcXFxZGXVy5tv6/ISBqtV41XhR9Ka9efXcA
U2+R0AV2QVG2pViqKLBKLO/Tiphc/0UtJksYdzMzD6ZolstI3bVhFVLuFNvt0dK8
8HhTcMp7BobKiDzYIiGGICp88iAmtzc+ZJc6O3AufSOwStwgS4OHa3a7Z99X0Hli
ipnT2zKiTE9HvqekkrMJk4FzVUsWjETX0OSgN7Y5AEg=
`protect END_PROTECTED
