`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAOx5cMeHRLvym6KzQ82UWq9nSWgFN8/set+btTKv1hY
YVIDDZuVhIBV9Lj0RYR3U4wccP8AIVUi4ZnL9E0KD6yHRdyRH2/p7otYqb63Vwj6
Jk5YsBkwh8V/x1dvjRcvViF6Th7joOiBRFfLJHRsuKN5SpOFVaqVEtiECyz76FJl
NwPmmpFhSNs8k65RzeCBOzSM3yWRHtAMiQXw9/OAhzsT+AqvhEN68EEIvsQUkKf4
`protect END_PROTECTED
