`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP1r46JhCFsog0Qaubuf+8uzYGH6krPDtpXKBSLfK344
XeYzwY+nIIc2KFENzxinFLrhy2ouywa1kX3dASMsxMIlCe4fBChwsgt1w4qXelHb
hY+dro7/9gF8+hQnrCmL2S65PIlm0wfWcqJYe2PGRim5wMgZSDmnTMeSQb/wktrk
af6aUptStP5ouvg8P7d5sw==
`protect END_PROTECTED
