`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIJFbpvi6G2W8WqUQ8a0NUdsUcgd0uipbWRjjlsO7IpM
ghti+ZV8UcKfkksLnlL9GAHVhFBmhWcLXrwhhOeQYRWQrbCV4mqU44F/b2dTP1tq
vHu32hBLvH5JYjUwIBPQ3PmKtuvubdsl/KjwdYMKc/tQ9qV7HDcEVeBHeBWd3FSa
h7v7RqjLmN92/o0WnaKOgw==
`protect END_PROTECTED
