`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
K7qH2Na1Dldjz712pwOPyziM2R1bBJt7Q2AocuVhfNeIOE7WSqEzG1xnQTlPLsf8
QyWWFLtQD/DzJQDa8UrM55zrnn7H18sIXctt7mdBgV8jwbFslNGbN+qmMMdhHvUw
`protect END_PROTECTED
