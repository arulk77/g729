`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePzpMTDIrwf8Jnnt8GTj6hj26514P8AilO3VRIqIcDzw
ZSplfAqOjuKuqpBikcfQCRdl+vmb8dt6wCLcZN4WG4aALwRtLFnX13ucxKmT1Dx/
ZsxY+3oTXDN3VofCq4wO61VP7G4cs61G7EQk10sCKBh6tIoLV9qWCT71oVZyaFVb
zz1aaIcE2QKBOX5Or8L9Mg==
`protect END_PROTECTED
