`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
OoqbmtICGEVzswyCA1x1jweZgNnpqGC8g3KUbYF/XjgDF03ODM/GjUtGuSDrZH/j
P8IcEt0S0sbvLCrcyZKYtYXsqh9+ZVbBXW+3Jr5JlJDyNB7PBVdt1SjOVumlUilS
J3gN24MqaSPYmtNOV902dOioDcDrUuQoa8d4CMatU+U2+5Nuhwf3RYQDpzHKnno2
PJvKkhpBkk09Z3aWpR7tsOatNcwNfuLbUZoRybCLaY7arJ302rpqG4uCs9ECZMMb
`protect END_PROTECTED
