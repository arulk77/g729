`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePErcgI5AVj0eI4fPBMJ1SKyUzECjuld5UbtjOV1OXi5
X5MfrLm5tbrufJ7V7o1LrZU5MXAXUrRxnF3lFYnWeXRmKszENsk6CZw9LGqxVfVb
N1OX51qKco7MMBQPZ3+5xQNAWftyo6BsfnUCeiSXQKUzDIUy+CfR9VN+vb7kKU1L
ku7QpzrugoUHeKdZTVXryM2ZR1zRx2puUcPHy2AhfXLH5/SbGBopnfypJM8AXuvq
32m2EncD1Ago1zkNOf/sk6kQBV5dUOejadX3fuDm/P4EZ7RFnKp+QFroj6/eBjg/
fjoixZbcRAvB6JWxGuIbg1rwc+n16NoY6NQdV86KFy3ZMxH9fvlXj/2KfYXTGDUL
iGmgh+b5FH6d6YiwNQRoGD1BDAshx9fvt3CixgjkmNg/HWdAgudQQRovShBX2iZ8
eah4q25/nC7BPxPlfSaZo3P6F67Fi3AlxEu3qigcP4KwrM77JBnKPOCZu9M5AGDG
fgrb7SxBhXiauS/o7TXxR0FGeQDtZsUP+VWySMGg2cMgisyz1GjfqggZh2dBMBsc
3iF3WAlRl1b2FWkWj5U2mlOVhIBg4rGf1WQZLn/Il1OdVdsJANrKMYmOhlwC1y2J
3amSTnFCmD4f+NC6hyX70QY/1RAl4BYDDhZTMkK+7IdDK6tJWAbmumTPAPdUoG1l
oplryUlwqti1BTHE0lqqQ29bDBzxIMJmPbJ2as+MaswAcQODh3GW2neiDUU/ERLO
yBZXICNG21sCKbDF0pqatZ1ykzcMS3H2iDQWC4nr3FJNiwd04IVKBgZUKTjIs0Uq
PdROtHQz7HsrRcSw2UfkgvrfjVlaxDAQZAnJRR3qRMShAE25mIpXpT/5X4dyibVx
3m++JsAFddHsFlrV3FjDNUNxqxQC7V7hYwsKJTPEM4Lc14ATEjvfFD0aT6+8PA91
JFK8EVOAYX/LwRBECPM5bWJXBvrkpyoGQ4CFYWH0bvU=
`protect END_PROTECTED
