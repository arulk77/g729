`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOoXNOpuidwMj9rpRKjaVunEiNUqydzOXNMRvTmIvf73
JQv7aVcaYIi1RHjUMV5JY8+DKiDAtkC1e8olS/xoQyU46eqxLFfAi9HyjaOKv5y/
Vi+0kz70PKHhuci1G2GKjSAtVtiJf23J22jzqICnV9Kbkxkdj32B2zHsMr6VDbo+
V1+5MRXz4WwKsq+VpNFWc9Zh/yFzKDltBZDpVj5+HJRswVKpYvGIXFsJuyzeqmeE
`protect END_PROTECTED
