`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SVRnVBQ/QX9jVcnXPvMIkbXvXifsczn7cFBO+P2MYWYh
ckeL6HT9WX8Z18XknO1rlAZk394Ui1obEn+TuC0yXtao58aSuLUIScnppybDefpr
KKKe9GoEJ0IUxq/k2gazI1bJKMxI0RMX/M7DmyKELEM8yrh1DXX3u8I3TrCycRje
khROAu3wcZZ9sxs2rdQGFpB2SGa6Bp5Fg4fW/WRh4L2ZPACBUFImUnSwaYsRbhHZ
VxrEhDLmF2ZXi+WbsF5pO3j1JQIdc8kC21u6QBWaedvuOwlojIu/8GRphwRF98FE
BsMbEGWhfNX3lJTb+KwwUmN68oLrae7HbcFPE8GX7SuFRoZRAvkX3ztt/zPT0tCy
9jjUfGS1XXAF/OLsZ2U7grhnUg8DoZQQRw4xUcUsAO6WVux9nAGYpS0mCzXC2ljb
72imkNt+Yv0oybh4svEP1fmEDHc0RdmyXR4h47Z8k+4wiT9y6xWDbj3mV3yxIBXI
J3gRXDhDj0zOcDjz1/NjhHxEbWDNAlA+SychT4CwFjzyECoaZ9AZiYbFFjAHAA0s
IRNROPR6zbJtL/17sHaUJ03suWUUkSGTRGbzi6jprGe1W7voEMrSSGEdasmfMkDS
+SnknXxT/T0HpOth6tx9iqsc4xgq8fHoqpG1F27+8b1FHXDzGioXXjImfHMyerca
LLLiiilgr+VcUe5t3Z5huQsZvRFCUJh0Ss8ScNGI1OanDSUqlxpk8TdbUbZcQQ+G
Rqj09zDzQ+n2whPtmOt6e4vQ104lGN57TllsbJ2iDD+tPGfaEcYzS3VxDzl9BQ8U
fs/rArNrpSiERvk+l64NB+qmWqgcgE6hWpSP6xZtP4WW+PYfRARqIdvhFcIJW65O
W+XFJimeRKn1USghcgXRjbIuoDBxynNa2VAgJuholPNJFcH6FmloknAMASgtMn5z
mv5csoxtgILYrtPlZopWSjW0ONIr1unpBMf2t6RUYff3FQIpKzkbqL6IcRo0Y51v
L1hcR/q2slHErFWIN5AbT1wrDYQpshae1TT+zkjLkXMZXWbI3PA061kGFUhyS41C
FEW9M1XTb2Lbt3hChVvMQ3RxldBzUoBIyjQwkbDHTwfw6Qmk6Zopr6sv6qxNSt1I
huijTTG39NZ1HVXU4Zzrwr8S67O1fKrTxAzxJGrXlcrP7Vit2AcMZoOAGkcLNjGg
P1XfTFNv7ttyF6XmzSObw4xkVvG9xAmFFIWwXmwBtpbNmwEtAFbkNSb7Uz+W6Pqv
3LVK0uG8pUb2Q8eyTfEwveoG6IdeiO2pqI3UiRTjH1P1MuQgjhh4gILAAtWnbWwF
1gZ0yJTTH2IuslYcEtFLmzCP6Ky7drsV2LZ6c3tESI1ZduNWYPlYKKkg035FWSp2
OafX2W6N6F8HJUNf98ntUo0kFDzbu5elvE6tEFyf7J90IMzStr7K9AoK3m1K3fjB
jneNQYByeByG7LFoIzsgBMLzJtd/jyeB/tAFL9rGITDyWcLLGde7OxZZu84ZcP7x
yK3gISlhKSXhslGO8T9dHWg8wTz/qUImY94TNLurRMVGBRkJgY5uatYRJAbe/Kg1
DFvKer9zEZnlf8ihxwdvVFbTdq9NOmrtej+m0K7PmsssA3cLGAAC85w1a12WDbCL
jC9gVvoUjnhKNIdFQwvQMAQhDklNOcp5B5iVIt+GE/DsQ+NecqOLUkWnFam+X5Cr
5nz6kerJnNBM8xsTE5uc6AbnYjOKCRanSrfHABgHHZtw+B/HfpXUtZdbNB7OPItT
LQtouAHMWoMX4MXT/BZ7h+SXTYjxsFrHbIxIYWW4IQj11zD7nmCVoEPqogwj6eXQ
rlFoOpDW2631F6EGm9Tmh8/3kRFgpOLhZF4IzFQo5e2zqTmnB2zE6mmlOFAZOT5q
JUpQzQx3TtJM2k+10CfA9sBf+JHdK8KFCfO6c6CH4X2TqFMJfeWXeqRrTpslzTv8
gUVunQs/VyQrzDnOMpff6XX8dJT5Bzcie2H55G1lZngAvhRyAEFLotm8y+ATB9ge
7ydlYsh/bNsAPNzb7nSSnlEN51b3sjcphTQMFxJ7auPQo1qZu/YMvnJ0kyLPO6hu
kxIPzpkzpnum5cB6oGvjz460lSu0Azhvky+hQz3bm+nvRwDvXXrOpRfYUD7FXo8Z
vLsxSVj7Ov/0WKmgyxNq7GzTY9AF2kf2BfBJuOHLjm241POLcGqDRUo7XoupkEW+
B7F2JTMMILnWrQErnUXNFbD0S71sZruA6s/UzyjMNMPaqzShBvCbmDh84WLoppAM
Pd4UAdAEoZToyS14KxZqFUppQTMyQyAiBSLV3nDNyfg8fN3yH6EWAv3/QPnY2HQf
97TJ9ulCKlW9CHKr22QrZR2kh3F1rTkIAnoFJ3lRv7zwuwXjzrubDb6sWgk0QWRL
L11QlTnif3yb4nAYfYw9ZfEJ29jxIv2lYUYbmA+ecJ2ckSczgYEqcic8xvFV1x+e
NNhe29meQvEou6RPtxVkRijo9+VuMXUizheXrcvqTq4ZsDnEULraW0ixKWSSY4PV
nQ3QrPcoFId/kGdVOsT7OKYs8iOJBeiusyl7lXTnvnY6IJvz6zfPSg+DYienIxkO
Qr4kdEbaTCiXDOWEudqiFzUXhlGghISYqgM7F+j5AzXmvNg1loQZkkQJV94QYj+1
xT5HNDL5miWY7+Etk8gczt5Mlxycy+3LPdFVF3YYozOG0DzcIiZvm6jBofMFymRg
izzi3Km9CNMoOweDMk6vV0ndYek9PD8Ap/SAf+MBTiU//MkkWlmsIsttp3LRyAeQ
zxdfTDZdsmQQwQgPHiABeaf9Qd3bizRKm+8ytP41lWJhUmqTR2KVR32p4QlpcOcH
HICEAkPCOjzk8tLhG5EfALz2IBaeEWjQBJ6C9Y0/io0+MFaPODGegjB5pm1KVSaH
gTpdLSk+tQimiYFKJ1rzHbsNXKM9dbNdw5BxIfmAjXWTbHmfia8Vsd+Kqjm+sRXc
lVH/upeCMdh+AmBq985EoxN7dUwWtaA+n2oHaALLdKO67x/6TaWurPBjcJgeAUoH
caT7TkFGe0cFjFvhxvxrVIKfwxHOxJqtleWbqbgG0WROmBqUXSx9ZT9mYr0NDmFw
T4FNgdgLmHLd+P/XNvBecvNhH+8WsQU7EecRJhLvepwOHRbvErkFCbf7p4jJApYQ
MjtKKRqj9hOrf8OxxRDqupsufkkyeLENFGRpDlYMsgJpmHzw4RngN+iyMJlWY7xc
LX0JVHcqqF5G5iwtaZbqHZRflllJPYlBil/ynBLpbdbId3LHv3Ib9hObd/wNt7QY
KrTMqGrL/t82W3n1XQr3gddm281N/tWJnD4EkN3yarTMYrCcmt0jCbr6OGdXwAm1
Ul7tDwAuyULbbhWToSOFQfAQfDB2+VKiGgih29ImFZFrl8N3zGNsBI8WqUqFHvJV
6oD0S7Zwvt1aV4ayxtJVM2M4V5fxuVka6uiCENisSOWsQGWCusxHeSYJ7uczfgAJ
BDKzSk5pyv1ZiMZYoleWr1HRtgxQEwp9dnnNGpqUxyt+PB5wNbD4HoYum+bcAEMh
vZ8mdRVUnfgx2PYg+huqxyeEhEqw9azDIyoS9wg4Jbk=
`protect END_PROTECTED
