`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJZnHDwGQVWkrqImhRDLfMjE/ClZ1QHt7Opy+wfyfUjo
AKlRuztfrS/9eLBXy/Nxqc/jM3iSEclVDt7w5a9oihTaRGMEK8ovJYA+zpcCIihj
UVQMyiLnxrcgCnHfRAjaYaApB59JXsuU201AhxJlCXBuouizLu3mPCt7bXaZ/NHX
NvkiT3VZFD4gXoXjDEmiLaJ+FIefD+ium79SP7lI1kXU2NnbagBmIJMAAeA9Hk1f
`protect END_PROTECTED
