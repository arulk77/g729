`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
hxNm9gMD2520udDdF9g8RLrs0APB7kNVZNuuhuivu3ZoENZ3bGlfBqLSOE49hjQR
HzE8f6sN/Dzm50M/hQdiYp5vz+FndM2jQ3Wo4++u1w55W5gbXBp96K0oFEMzDarM
OZGLFW1+t8rri/0RL9z5YuhVyXeRT9jC2PNRvNFpsAUo2LjR07b4bMIXO3AzxVsR
7PvavOpjOuAmPG9XQxMu3a+khrXKviHjMFbzMnf9srZsSrpIkADvj6HeYD0tib8T
RR0uGX2eM4c78hGeYkxkh+RBnfu5C5ZwtELDWROoJn0dItJPgYh9puzu1qeW2Qj9
98nYiRn8tAh6iSFc2HvC150HWGQrDnUmHxAoSoUyP2c=
`protect END_PROTECTED
