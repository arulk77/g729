`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JCCsCOhOaaovR91eUaqdA06SHn8Fb9Kkgo0IIdSeywSUpYYdUR1o8STQ1qOA1gCS
8g4v8z3h0RqpzhJi4h4EKZ6rC8iqDuqdbOtoCgBYDFlYJKYkeyfoLvjl9dDUIw2P
ZtpKksIjbY40Y8uPt0WEWMyQ7/klxZ/zBRjWxjeNvkc=
`protect END_PROTECTED
