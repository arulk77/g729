`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zm7N7FTJcyXIYpXS5MworFKZTlDPeY8hhUciuPbhj9m
UhgfIt+TgB+L31wOKfS+oganzFgB09Id6WYTU+zwGv1iQydPRm4bCq2QPm8xh0Zh
DgKuev2QZjgSA+Hs4Qpnn6lVeLxAMt3X0wQ+qE5Dg9fDxRD1azjSX4Y8ClMDFxnd
6tmwFoZOAW7pFDlt8sOWvqfQ0F4fbd+t+Qzwf3JS4pOI3Tp0GBk6THfG3ctMETaz
GcUxpcA10OZHRYidu18b6P5zFXSfISpcarGJFnFGKz8bVwqOzLZzWFIAVodfpHKb
eZYupiCctNpFGIw1iQdNeQ==
`protect END_PROTECTED
