`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aUSSvbESxMRFo62RAdKTZEbPARRWrc990sizCrU5mFCx
LsxTKda6ybJJkopI48mhWJbaLDMwXK3LsWp/qb9LKvD4JzzRxOlSXfJRklhvW+Dn
qLV1pFjI2dYBWKp1rhPA9LktX0HlYmzWGSSnzdIMAB3uvLgKlyy341cbXDzABojX
jX/I03jedD9BVUFkk7Au1DWW3hJ5u892ymenFnqkRrwpVIShmvjRT25fZk1rbenv
Z4FK1AzBicqo8Ylfl8Wnp69TFZK9wkfRuYOW07WOJEEE8a0H4yR8KwLnhnTbJYjU
xvJyjuUwcgB908kCrSv0xZJEe3cEsXHSXIHbjHqEK8YvYFgr3uALjzDRaxUxNfhI
yKo/Zvb1d7PZR6Wh9tmfjpvUE2pkqDOqrdyGAyEIYokZfWxQKUGpvBuikIC8T1YV
817t7S8wlS1k2+YlSvwwrB0hAi4Fvz5xkAHqsCTgtV6AdeuoPOGjJrmSXD9uJkxV
IGHGj3kTcaY7XH/OYpmy4tn3mwy+dnLb64toW3ptFXs9B9afN8YuVXdXb1xrDkU0
6DHR0eRscE4lfWeT3OQOlpWJWX2sbapIpt6uH+uRrFcWeKTG+aleUSGZm07Ue7fY
UCVWnXRYBmY3Ax5sQ72vl4p/rUrxyuiHMyBuZjjS9meb1jXTBIJ+bQ2kC9YQVE/8
gDfZh2XaIC6xj1Fwm3An+BnFafwr6x1sA9C3d8yHY+g5akPaedXL2i00/782oCeu
olX0TOYHZ8Bu6uaSDBeK6Mam0w3SkL0iPb2Wn5uKUXMsjwBeNYKS9yeaY/nvMbtF
wZUD1bRPLR0lxIEpecTNM7VaCx8OWyvqXEXiFLwjcmtEwD9z7IEk0ytkI7tJfZzt
AIbkZxfY57CJ0sCTvnB7/8s4JBggNEz7QSXZhlHYeZUjVRmVG58mwK9dAKcx2x8B
jSaX4c2kRFOOR6YQD2WwMeWrhMz+G3f6o4P/4vne+YFHAC6j5nUZ+cjIz942mpEI
EBNiV+BSl1pvFiMlpr264WNBLyz4Rdw1so3NDSYAiG0xOeeEPEh/esfuBdN9WINQ
jYV4VWHS4uTWdbWloEHxMRc+/utLbuwbYs3LfTf76fFxJwV+49EGstyAI0rHvJx8
CrqprTROS6qAYiP/BOk3VwHnidDQV8xE7EwyEuZ0M/fV+iaPvkTqR+Sy1wGihim1
6hdNZMQxfvMbpcI9Oi/5dx3j7mtkbIBkZ0tChXnPzLRlRBglcbrAk5lCaCcN180S
mtoOZlE9HusgHso+4kZ2oEiVbCuML+BKjxRLbUe0iaYAKxg2fDtrngMh79qf2/xm
iLd2ATMMrW7P3unToP7FReB3MJJte6Ru9a/hW4lA6GqWEIpqyKyXuvotWxkeMNUl
MScsHioDO7XjbNVjpLpQDEGssbxCKSb4WyBJ+S5gFxAPDRlzcMBR/rXb7DTNJka+
ok0xJJDAvXDEVMbxW2cJX21D1IJ84DWJmZnMzuy+xERARZStLYqJWZ+7miGis6s7
VSE8zAIT0ihrQmUUFrIhrUBa+RveMDoA9v2grSRmAhDQgzWmKzW1PzUPl2CrHFCy
ogm3FyuVK36hpx9ztc8zrqapFeRrjCXsSrUYNxfdOV2ke5oXxTljfIadPgIvHiWE
`protect END_PROTECTED
