`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SY129Sys52vlPNWCpBv3hfyYaco4TcrsoT9zReAtSCq8
Zwu4DKQoDPPOjEoJuMdT8v2IYQCl7XFX9qNoDmNnr71FyOxbo7k9LX6ayD5HOzVF
p2506Y4T+x4frRivk8zLnKiaLJBjZ6SvIb8vwKg1nVtO9Qb+bb17Pr/Un+/S+1Jl
q3w1h1v7le+QvyYqV9HcLA3/Ym/zIMExPW/cOGqAwTLvO3zAwRSTSbG9oEiP11GG
Gb8BCWsO2d09daFpVXPDtqJeXYZqyHPXwV8OkWX8B/k+hJDbqoci9/vE2MlrTwG5
H1uQaNJjoMJDWoB8xCCHX9I7bTgdZ1twAi9FJtSQ2ptzHqsXnpEsyz4jUTU92LOD
TVTzi32zE+m5pGR3DJzZpHyfF4+IErHLhutRhwWD55BFAX5OvLrKv/IPoSL9ecRY
cCyS2R45aSH7uMTIAxI9gQXkWa6DGha50Nco63Oo9rvsf25mdxe1i9ez4gWo+07K
DWH/BGSgKdElKw7rPAWm2VcSKYcAPwuOI+ehNZfCrNJ45HAv3rDZpB1wQsjjxhV7
TgE0uCciOtdxg4kU7nsu26VbFRTbEZtRAxoaL3EmZQ7AU2+sQsME3Az7W8z3F/jn
uIhsN9mXclhacQ0f7E77kgStQI9SFIOji7zikhA+ZcpzvfuNWMO4OT0SW/m4A3b3
SjfZ0IPT/e2BBvmUOAKf6WNfLxnSNgZU6haTm1J3ptCaZKS4cT/yweTuIK/f88WD
DBlDFde2K1tLqZs6cod/4RdxomiwOpKAT0scn5aYZREHPhrolbcSxpupL666+9M4
1c2NyGuDKEK8lOg/g8enyjfUDo7Pp3lthonDkYWb0qfRiguUADZmGVd18Q3cDinD
IHZOMkK5bhMCEl28O3zuE6vR2vkqWI1miZe/eEFZJncu1vEHO3e2L4jtykbgUZ5b
YbEDXlFhxXZZ3qiWWf0cJn9QCpEOyLQwLoH3Wyzh9FJosTlVHlJ5s342ATq3LHv6
/orATqoPJiFTWyXk0GSRkIGcmbn7ZdQ1LU6lJghRjQHbihQv4+PSfNuPMXZkAj2n
Pc9eEWG4kG+bE46KG6Xc4vXaXyW0kVmkmyLi0DXPzBC+XPCSsgI6hmo7FMJvHdVl
o5KpbBdKt1qJs2gJb21CkpSkZsaY13ryoFUDwTTtJuAs9wxyb2eS04zf3hF78py3
gGScnGPZ9FU2qhUpOOS8HPbrOBA0GcPrYdgS8ik9cMs4JO1oXu15Ql3NEBGpfWCB
GOY19gt+4wgDoX/qpxF/YAJ5QQXO9mezZzVB1A22sIxT759MK2PC2302w9/a9niv
Rg4yj7RNpOwtsYoH5o+7sqgLjfAuNeF35fuK5XqD+tWe7Br/iPyUmcLekz6ckaoK
9VrE0hkagOeH4uJrx1XGKi0eqBKH3aMB9VNWjNYNDSgAv35LduRPBdO3MqYGrKit
z6H9fSRlVZTdH/s/UZCWBBUWdXz/jDb4XAI1BMZY/RrqiRxsUyLuk+fcVHm0NGma
oP2f/OmdmPKEyzboq6YRbtFfZca7Eht5AObsl8nR6oLtYs9sBdk+5RmQoG76Og3o
QQ4qTjA7W4d0y4yw5h1dyRJiomCQMoVxtGv7aSN6+YPqTKF4j+clhxfJN/Ua37FX
TFlteTqTOyGRReolDDYkdV44/cqhsrgUktn17pIaxV2GtrBzVBOnd/LoNevebhDx
ceVAkrb9n0cVSnG+aADV9rN+brD+iYfl+ftF+jytkhUpJWAEavdSmWYi7Miro91R
Ye/cEd10bHehOJkdD/iLW5PBGTdbxwZJwaAs2Krl1KudsnbbNinGu0J2E2gfv4Nr
nFEfmvIiJY1+wFI/i3AYYVqwZGYgXKt/J3m5NR5B5Ri/OrEs0G+d4UsktcGvnhMd
T71aT+TDwN+bRqqwBbEgCae595qktkD3zmKGrdTpedlPrfPF6tX4l0TjM4dzozuz
AjaHOgpDoSkaPFThaAFzzcwuC/VIanGiKIj4sE1om3fv9xDyNzLLFjEsqm/LyoLn
IDrskOkS5VtCbH4i9axwQ6pdxTWqsmoQN7kV83UWxoMESckjtZAEB9QNokCQA0J1
bEEfwQlaDUN7TPippZN2aukna+zKylRw30rJdaP/RqXmmUa+5TwvL+68b/b2kMhw
2Dd//NiTwaCe2e812tAGpl3At5c5sXWwIxBLWPTrle22LpH6g5CJSDFIspszCBa2
Mmnl0TqHoQYLa55Ka3nvoYcTnUPwxwFMF8DXXrHBqfE7YVFcVa2AEQ0HKgKTMtSp
/0Jk+6x9W9ultJedhipafK4DNEa3wLlCiDsI7o8LvN32g+reH/iQRLoIH2Ibjjo2
65u15qQ1NaYz7xhg6JU/VxiXmgqsygG7a2LzSClpWlXc80KmOrHF/UWXGU55gmtz
XloTMSJQw2uFv46kMPjqcXLZSkpiF8MvVcUqpq2uWchpzbkfkvQpEAEcL58atwvc
3gEsKU/0+FvYakVYwYAP7Muuna7kv3do9VjmHfGVhja3egCTjjVKx3jqopT+Sj4t
A9sWli1p4tVEt4NgD+O5isbISqOs4+Tcdcube5su6xTWf1Q0xIGhpyHDoEpkrj35
r2zAOkrupHOPUJkN7wzcQrJQdZSol4Q23qn4KunL9WpGoyNC7CAENXkdsRrY1/lJ
d4V5X4zyZuTkNMvbpFmxJD2e4J/aJ+EJNuD4vuOOBWs3fUHU4I9tUBtAXKKv8H/n
LTTT38uwmgCtGVcZGlYeas4wG3esszDJXVngjeOOk7ZRTU3PkHzvVoXFDH3TWPzF
zooHPyVslwDCFwdZLPmQjp6EdcDpuR6gkbAtB6c5nB7AUn2/Dlmegjn2VgX+gmor
OQEjzkwBVPE/murbayldQCmPBHJOsGOlCB1ks0qoktwvkO6Q8qWaZVpfyggvm4xe
JGSt6k0fR26P0CAEu7bNZlDexLytUINrPMb+YmaL/OKQE9yfoRv8QNjb049h7IIW
VLcotbkAqnfwWN2ImDlP6Swlvydh6T633/fBI4AgoC+jor/vSXtl1qjD7MiPBwm8
twSox/RfegHZPxdB3lyIisHhobvRqCcpIeNGn/bP5IjMenOoyT2ckx/v0KEQFPUc
VsPkpvclBLn1ZZ7gX3qyNj0FxPNOPFv5CwqEu80OlhIhRs11xk3/d+AAC991cIvo
6YKTjrzCSz40xWecS6xTRAJbiafRznjGsLBzV/NP4m2hm5Pf0wsX3sxGprsKP79/
B5r6RmN92mGYAPXuux/zIh1wH5EqGNF+8CmZV01kzyRYXwaVsiV8rav7k9bN7vBy
eyZEKNdzNYHVAzUB80cFE7xNimMiMDQtXRdJMHJQH5gNP9KTC59pJsY15LsEoZ1C
TCyTa4DbNgYlcEXZGFVKlnjqRt18oY8VSiYbeI9SGJaBKxEN9LuGYJq69Pl9e6Fb
tJnNCB63VgYpK+9PFJM88c4PSBY7U7JjmK+gijgD9MSvIy3j4QClxwBreCkWo3Es
PUpRNEB6qU3QO6B8HTa9uHAtrTCEsmkm24rkvdgloaZe0NcLWwbFDjujtFh4ZTjl
mSiBRQeZdNWnSgpqm+7EWmLkCBnZHhrwfV3cMtRXpT0nldoZ15r6GrtJavJ7Ghlr
bzOxGLrdsXa1HOHs73ED3uOSjf34Mthp8dv6L12WaF8V/a1w20JH2KWsXfswjTKK
2anWCDBxwTYU7OopDQNBZah05qpK99e/2lJpCCnGzZqfsqLkmasFoZzusTveabjT
JMs3XizEaJJ4ee7tSDPHZtRoaUdWTR73TYe9vlCAeziQtRhZk2I558EO1LznZHqF
uRFokenchsZfPrCApDcxfISzn3QOwStBefdC4cHYiSPtjtceauhExDbo703UnVTu
do9XviWNYIwAqN3L4Cp6UdzUlCJF6tyqBcd2W693A1/48VfmP3cC6lnj2umyxrsx
yPPL7sjikW3oqA/6gDLAL0jSB/C7vKk6+pM2YfiXvbtWbzfC2lS0SnOos/ME39PC
ybkMiLdL5XYtRRCe3Y7FpT3wGAsLe0ZQovOwgkEhuc/LFNNkrJcgLv24kxnR9rkI
+7bPfS5J6Pj6ULXvOTW/XDxNdOtxwC2QqiMqB5vAuPZIFNlhMy9hyaGwX6Vpt4Wb
xSVPT2plqlRQQRYrPQjdDw==
`protect END_PROTECTED
