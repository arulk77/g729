`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFAmjyx1Hq4nGJ3kz8SE5jlxK1f/3IRBbmxwkxs+v3ZO
tIVL6uGUbERDlvNV7kIbuCwLyu/lfUMR+KSPQ/D/SAjvP/Z//RVS6iI07IoRZWgx
1/nn11nH2XwliBfcnYotqYIsL6zAGRRUNuoXw6LbseG3te4rIeyfDFN6jRIeLCUx
ORuNNaXSgrb/Qm8yYaJkUNI+Ru7XzKcJ3YC8khb0drF8iMSjAnVTjFhhw22EGYa2
SPvzdwKfmUxDkzdjWpl9GyzceQtISBIzvfVkQ8jVyY1cG2GyYPI+DPkBAiNhkkPo
aeqG5rJJesCUrNZ92p3nWICjx1E4cLtLrqW8+7JM5yisEpaugqO57O6HvGGePwJS
PtfMNjnx72MzOaFma5F7t/Rl/KGl4/5fKlwxpAD/XVMNPdOcsdSSe6OMun70d7xP
zyDO4KCD7faKZ80c+2SY4qO5X6dudpRgQcsAIBGdx+hBxfq+xAKKig/DWyIdnZet
98Fo80Fzb1FLgTOhkFwx57X3KwJ8FT5LGbVD4e39qGXKdp2MJMbBlmP8VUEvACrW
zPeHtu2ITNOcJlcwVG5n/AcXEjrqLgAoBWLKq+gn/lNSR51o3Am7jIcz4Xh8myy1
`protect END_PROTECTED
