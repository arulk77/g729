`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLysTbEpl2W9nKQ8orDKqokHWVBeTRZsPkgyFBgaQrMI
hOjsXR6N4hhLYzw/5kvKl2ejjMKteXoUOcX8dH4Lr4N0lUr9o9MFVut7Rk3ZD7Da
f/vJPWwePlMN2Ic5ifnqydE0MK62o4PpUzIg8hQG9DfYuYKU0W65RYL5RB1iaIAG
ZCUx8Kvd4KOyCS8l/SsHvw5mNV5a3Z4M4LRE4vMNPNLE141O+s4OiEx67nrGs4zR
T2BUK7vlC8tSK6PTX588Xkwp5OITunNMEDqWEI4licbr3vqB0rNuw4ST5pn4GO/o
DtXcAoPiE8XCT1EoobsoATh6Uuh4whId2hTXQ3fhWJIJ7/RHBJhOdaVNMGDipkKE
0G+xkX/1TUVKA3nelRm5IWNamB5uWCZS8JZ74m1Li9iCODmFydfJWmmAyXlFVRA4
uLvqpDFEicCP35d41Ov1exOKw7GtCXkbPHpnZajdgySCH0Avs0azPkv/R88Gzqxn
8IYLCLUJgHmVJ6tGAWJjOW5Wj/Pd1uMgqJvGNtHF2t8=
`protect END_PROTECTED
