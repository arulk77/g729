`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
TdZ8XC+THt3hY5VSCX4t0RT/NcpBtuISIPULRn9Pt5uBsOCeCNpfY9acoldqvKjQ
fG2iMcVDW6pFmz7f7T9/GY+LJxdX0cXmbZZZIdfFze2gSP5NrR9G8SmbPiV00fnU
wBJaq/jM7xkF7GkWpMzXJUpA2YxIBI4xMgc2CsjRIR+aw8iOWYhA6djm+xlfgJPX
Xy7iWCHFtQmFOgO5HRNMsmgkld94TOdIdBoYYTLDts6E1CE/4fPClqz3/kxcV2Zl
LnrrNl4grhQlix7RTBGUWDVC6c1V7ExCVJdq0FUgj5nwCqLoGs04Qc2JtRZ57ouX
O8jv9OkOp5Ul8fonCfgnLMvocyBFCMWvFtxCsLyfM0E=
`protect END_PROTECTED
