`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePszB7S5yWIq3IHJCCUcVGxXu4vVM9Eeeb+sRC8h4phV
t4XmopwkkDmTwKGqNPTIST+EduW73pvELR2/eWjK3BDwqqflgS2rv68ET1ov8pF4
4WMRFZWhRrOm0cF5V9iZUoDsiI/pWqFMAqMj4szvKBRN0l5eal4fLctTJS0EZIa+
WHcgn1MCdqpdgQTNDwNHUTNqLo3MzSiuEnkGIZzakCtH5dxoRhupA9nKAVgFljND
`protect END_PROTECTED
