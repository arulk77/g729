`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
0Q3O9BeOpeA/ZkuwWdrpHFfjZs1et5kZL7BHW68FpOomj4skwJuC6zRAwexdSXAs
KsBPzM7zR1cufj3UTnJX4I7xLjp0AZ7Do6UXtB1X7tt1syGvvIYCpsGjKUCUAb3x
JJABKt0DViPJPpMXdMFihfA59JfFeS0CDeJINXj7eZKlbVx8wJJzPvJ9QtAyy+q3
ioITX3eeWHw7vSwcJEoxCKgxzDj/bXLxjWtctE98m+6U859/Cis0XffciiF9JSPv
fQyA8uPDSsy8GgvmDWTDJp/U7so1Zx2o8WRK2Y55lrmVzryaebcC71TkzSvfMNsQ
`protect END_PROTECTED
