`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
LXCy+q4wRxlUrLksQFCyAWwPuPEYAGciSfy9O8COOl0j8M7bKoNnEJCzlwz8OW3b
NF0j/y9+wiM1PwSn98nwXbVyUlJVot2Y8SgGrLBL8iKKOkSsYGiWOWwHkr7t06J5
vnTOGvBjIsUKKTlV06mfq0F/28/cEkZMopJlxGnNNfS0F62FxMA11y1UXcQGxZ05
G/di30Rvxy0Bz6I00tG8j5Ctwi/tXiaRQP/5K4AosIa5RpzR9hNhV9UZM+VZqlJ1
zK0PAhRXpL4jDScFv1+3iSHVy6uJjqWcsIkaljYx9bN54c/XS6yC3XyavZZ7oeg5
frTy8mX8iWHNsFf6/z7MhQ9L4hRSaQdM46dpcqu/Rom4fiAf8s0a/fftjnNrrmKv
QF+Cc9lZ7nAR1S0WgR1clK3Uyvo5xOdBMtfwF0LLWgKsNedhXNvQe002Eh6CJaP6
y64ekMI9TIon+SyraCpapxSylmKu84AiVw/UM2WGrGgL7xWsvTKFAUUXSZne9g00
I2lO/4yk1wRZUDPHbdwSrkqoPljgfRBGEVMlCrXcUcAt2dlF3VpwIN5f4Fp+Z6Vw
y5nna+FkQh7Xcs+rka18femLG9i6rB6hXuaK+uv2HBkvec7HSAGUcrCIxs4YHjfX
GbawayjBqhFTrB/3ELURngIySYEgQC7sZfSSwkGD2PjZ4usWqxw0GAbFUgVv2Ijd
fb3nzSPFYuU1NjG/WUyQ0FVHVq4acDwcWOAejzRSw8M+PnGld341j/Di7ntdopVP
LB0ATOJuo6AAecEWdYOy5pMspZT2IoHjjcOI50BVC9U8NnUtNlGY4HHJRPfgf3tq
eo/4ho+YVf7KnyCHlIt/LWKc1ih/ofOpVumQWQAWlYkWL/ceD5QEnLQ1AzqjzAKO
LvKra88pDS3N7RGHKEuPMjq2FpRzyY1Yyb7KeFSaW6h65nrywoFHP4J9SDI20gtT
QLO1KU9vv0sk7yEgzzKXxId+l4OxQOdhtTGxdZfWJlXLnHI652swQMV1lkbHi0Jb
pXlG9iFkmO+/TY9Iu0jHZ0ls3rOkw4nO/u2MZk+Q3Z7+5K0IUBjanshUyYgGou4B
701+d+MEtLHeLo9Y9GaPyo7ECtmu8Gzyw7bDSa8jpYYa8dLYS3ju0KY+HRzo/gr+
mMKohJAl2aRXnVKjsJKKI2mfFF/GOLHEOPCmwPIl1tJ3HkKbpupcLFdWipvw+dZ6
Byksn0dt4PnxIcat3MYbXMygIwSfY2Erj8acnMQvAH06FtNdZhq0pe4awSv3051p
pRMQZ75dqLEM/oZZF/gzwMfpHv2nbKqMqXHatvdRzbyY+iGGIT74HfAOKnh636Ly
Nozb2DOA6IeAtn8xHezDW+AQXAPvRhetllCpW6u7KARIPYlSJ6Ca9TxPPccjH2H2
CZkO0Eguk+3uTqSyfTt8J/duhjnYjww1yHCTIuWxFdAiEFP8QFP+TcehNULv5xk5
1lvTsqYjZ8LGuookwVjWhb7TZbb3dyHUdXqlVEpvz7GkToxB2uq5FZ5ODzESMo6i
qjlg92ZxGbkk1NksAJ2YMVbNw++kMjD6E37ShahHg26qw3TBb1mkTfDI2KF2fFAz
6qCrX6uJtL03Fa4AGUyF1RbsTLSvNDqu/u9b3IUQw2oRNGM8W7gsEThfkhtOWhoA
+dsXdDWkzAIH3tu2iRXvx72gSUzYrgK/zb+wY5fRBZs6b+IzojRiv0uSfweKdwc3
lCNBeStIwPai80469cK/HtAjBo1IHSJW4EfobYlR4mtlb3B5NJKSk/lQNk3A4PkG
qyGiXWlimvUFgtQajVbA31H0mm/RO3MrRWfukIk4ZOmvkRN2FptzXGFM6NIbFHNs
FJzg8Tyc1E0/pvIquy49ov7F+HI1mq49NEYqUSLLd07tCEH42Aj29gH8PQH3ljqs
2m9HiBArhcSTO11ckTDaxMDV2XDMvquJRvkIg8/EucanHqqwyM6Ha4bLcvC5LKCR
Wv46g30tiOoA8B7JaODlalJawVMfBhU4xGGN4xYwMJv7mdi5C6YJ0ycMPLK7uExa
rJHFxFI7ywseIGX+i2rmZ8kpNBked2tC0ZEDbgjxCPizfVNZfbhrm1jF2lZ+vza2
Rl1Qs7WOCG4o2TT9UYs60ofD5jLbuF2DOB3bt3r6ADe8FMouWrYxjzO9Xutx9AND
ZFsc69Z0RAsfjwcgl/TOGh5LAlK3HveIvQR3Ae6Bhgo=
`protect END_PROTECTED
