`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
76sFkWaWtW2g4TUTKwVVqqaFhY70nDhVe3h+8n9WXU2VMgA4ppw3JdNF/G6iT65q
Oj40QOGpZSQyVe1jpn/FYd9Xh5FFlM+ofgT5+DL2RwZhSt9gkaNl44qLdF8F/xWA
Q03Ie+vabP9OdgVDWUBG76qnYo+qYqMyNMB+0N7Vu5Efu992de9LAMwcg27vLRhq
UCSfDWHlQWqWNr0s56COyZLvgdcxm36C3Tp2uL4qYEf4Zy1PRHeWxOR27gMD/CVG
IRM1ymUsX1eArENuUfTGAbGBesgOpSkuDRehuSmFupUE0SBkDEFB9QqArNmRJodw
GHcNVJGkZW4RgROIUZ1eLlSy6UHf6y8SUUh0QVTgHod3Zg8vrZSxIDkDNtm/FmXk
kOheqRw+U+jIrCk9iyD/zZUoO3cF7qZpXI/s73fX7jujSbuGjEMzMC0KcO39gm+w
xTkNop1a8mLhkHbFQ+Ql4gRfjYreU51/xvd7yVX+IvVd1woL4zj4NsKXfPThHrjb
sPp9GZYycDJ1UYD4Ye11GxecnZJ4hZ53dzswgcXpjhQ=
`protect END_PROTECTED
