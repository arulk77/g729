`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aZYVKa+3Q8Y8JuF6iEchRwhkOpbHLZq6gzGUlObnvHmo
BhG/8Qg3WHx4BKSIFVQzLPz74fINsC06npe8xBHpXPvXwCeiLQ3PaUaV1Ae8L8uL
QG4kBQLYHQT7T7TEJweFQlhyb0r6uLuMBsldo/QNWMhgPFBbQM9ERk3dm5GoEzfa
6IDSvwYgO/nkP9rdegh32P7mTh0wLyaJG5VuKIacIifuMqfLD0ZXTyVW4cMK7m+v
5U+MsY2GCpB6i3FbAC89mOISaC9D/qobVqnbHffpvspnTnXM2w//NlpfjY8XVu82
`protect END_PROTECTED
