`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40MBVyUhZ70j6Mc++qblvcFQXa+s8K0PcojxzKJPD+P7
ipdyJPAe4gHwAvi7HiLzN/U51cR+FnqG6EPL4G3SlxV+PmbK1eYpWUVY+aAI5e0n
uznpzBbfNDQaZBeAZlcUPaJ9EujeXeg1SEIXmnS1EVqkOANPMGOJs9G2eoPFRy0K
tghpncaqrHgvKZBT9hy/zfAuPpkoyEJZeIj/QKYA610=
`protect END_PROTECTED
