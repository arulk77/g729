`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43O1coIhYiYjh0Q0YTkqRgDrwwiszf1NCQYf4B4WSXsk
Z26huadmzs/sPZH8Fimk5FFg+M1sznU+zNYEa13h/SyhKwFWCywN28bW67CEUrgl
b31H5LDe1Xd0kenF4tWlSgzN5McRnXPXmpJgS02u7Xrd7H/7B30Bh9SDGHl5qF9d
AjSknIHRF3A2Xmx4l1lQPsgwpw9YK6oYXFeziJiJuw7zDAwjGdinZVmw0TPRrqeb
zHBNsVP6jjOAP+qF0yYkVdAjLFyF87x0iAxXCf7AOE8=
`protect END_PROTECTED
