`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
DrxA8BWgL8N3S3JiqK1xLoyqdq9LOlYBKFp8sEQZBgxR4wpaw/32gxAKCtlYmhhJ
XWR9aEGrFgmVBBiMdRcdMl8acebXQ5/AegeU4Ams0iqZvtu11lYIDihv+6VMl/98
jdRikPVNKmHv3hTDAjsXhCzP7XmJff2/dwGuOrkFKAed5BdNeNA13ftxMzQaV0IR
BzX8I1A0zBk2Gt3RKdAluSogEfVgKm9D2pXKhnlx2ilpR8DQifqKYXHROHDoJBIv
qoSOBcR+niJ1ibtxMPWh+1mjLkvhRBKWmNY8mHr4usXQQHleKuL6oXF6Qo8EZgEz
MfTw3uo3gyRphsXDw1apKWQYW1Xoed/ELGsRjXVHLEkTWGi79Wda2p2mPzfBLb6G
dAs0FChk7vHLT9XYkG3fiV8gaSAhhXgtN2uLQ+MEhQs6Muj3m1womVz9IsL56GDK
BJOlgWuJFg5bjc63szkdsA5sYWY74uKUDHGrHBjrBob9UXmYPR3N/b88cyOXnswn
mdyAiRYDmUHnvNsV8PmEkit9vF5QCBlzIbtK+vRKUZi2V6rFhXLLzeD13Hqlw9Xl
MNaOB+Ee+QIux6enwVc81B8lg2E0N3piwJLQI+vgLn3KcFJF2eRU29Z9bZI547jT
DFNXDd3YmAeZCY0zkJpmWhfVPyGHRSP2Ir2JyNANVhHDahVMMjgD/tPQbDs0SdxH
gK24FS9PGqFBveTcexFHR5UOVAD4OarwnqlUdap3u/dl5C2y3Ct1FlBDFFyZfkru
p8ZoMn2CZs3i7Lh2PIwQh0ve1Urfj+N+HZ2sOtzl0jothkaYQRzCR5dgiBJK5MPg
PZWNQ1xew6phVKJuyOpTOu8uh2vD4r0JcHy6sY6un1lb7aG3IL0PywOWkj2gbEGA
VHfnY5t4dopLTPAzwKTWjpNUU41ieeN5RMSJIrT+h8DvMoK042ODeqIN2mpu9mtK
v6qs4D8mqlbR5Vs4FrDq/2AEvk/KgbbLosI5qadqR0GmYL1XUKA/wtSOxsskJ9aD
aUz7lDzdrZqcXX/glgS23bdWe86yKAQg4udzYeq+/lIuJsyRLoGoWEZrGpIcPGZN
0f9s0tpKpKc6pPf24UBm2/McqKXRARgXgBkIZbg5nmETMfeyjPhD+mqf5aj0jPT2
DCLFuVkcHcPyt3V95c8/xqC4Qa1u32hInSdZ5p6t37Rs2e+afwN+iO3DPlGHCbSh
cbrb4hj6TPvJ2hDAH6nhoENDE7xIkp4q8ljdSVmCSDDUw8S1vl33xAB0OGR8DVEK
2ZXCLKDw0FycG6LKxHPHi7K+4rpwvgaTtnhJcbS07IxLMlOO9DBOdtNQCBoe4it4
bGvFU9QxYtgrf0OTfvePZPM9XsVV47jcx68ZOwd23NP6YWtYViPNGHKbCEhyNkGS
tbeXXzb6cRm1gij987OO6tR/99e3lTBQGI+nFtK9fPBIU9Wa4gWWmgps2w3AZcUB
w6ILMCF5+n5zOQU1C0vs51WF+VDFGnhMK+7lHlMZJx+4mSifMb4SDd1y3EP4WThK
eBVpcm7F0/5nWgBIP2dEm9i7ZYGlXx/CRL2BRgnHC4phyM6KfD2SD791CT5BLBSZ
utWKoj8xKTIbtYUtfLFq8x9d0DI/f72eGjN4il+/C2/BONu/NV/iIvt8J6zYq9hp
uHWVyS5GmdIHcRUeUxO8Al7RsoJpkbA0XEOi3YJp+COvniZv973CWugLRujYqCFJ
FdLnkyboWM6eAnBEmMK/i/uj26nYJO6au9XIxtkuTw0mrndb8o9J7Wm7MAed1xSE
1wzmjAjJOtdUAM3TKabo4IGIs+xU0Xub3cA13GpE6zHPpwTffpNtKVtnHuFhMY6Y
IuUP+YrMHDjNS5jaMsg6WPh15RjBbfbk3vMb8WEsDfXm+xCXk7rEQGmOkGF9krF2
1FgAdtyFidwtyiwkAe4YBayX8IyS3hnH066XkFGB5KygkJZg8P5yKiDSUADQJ/3b
ciys3MOKLuAijgSEFmherYACSU4J+DLskoenFUtRMR8h768Dp2AY6y5cKSvjPEo4
9vsYkW5Qf73JtWO5JjBpMp1ZK/EJ1pL0JUpWMHXD4pGruBMxxzbEHMSrvGMa3BBY
2/8PogE7GKa8GKZzkd3v3oXm+MKaBO1BBM/ZYztCxoyfiSxD8R14RrGCmT+0oSCd
kmdpLHFe6WNzAPrMGpvrewXBViqFymty5VBCkfOm6FiGDFwGMIU61BRGX4OkkFM1
dOiTIUKs65QHeyE5uK3Pub/T4KfdzzUOp77Tv4q0fyH9PE5tejlL3KTMbCObXEDP
xr8dTFwIVnBZMtf/xjUSWzEabJNY7JpmGIi8IembLkAm6usyZCtg9E+9E1yaNeAA
iHUswzBkjn8l2oqaxTzxZv2bNkc9KXFeU91UvTK5giUXcDATyXTWVS8ORGdxzRAI
PXs2RED+1fDJUHTYEs4VsvJ3k1TIFstBK6VIwIp5I2XznT3E/KNnVDQSfFN9QHv+
MsrW/D+LVFNlrtOH9dy4IQjJsSYZyp97Wxg1mDe6Y2NhCeByS1zGZHiLxQLTjKvJ
+aitlys2arX2Mj6dGFmuV2wQsv/sj/8qWYylylNs5OrRxuhMm1W1PrqPENheN/MV
uFZscSoAyS+N5f2sPD6ChLowUMkeQwAkc7fMzkUfo5iWfd0QIhpW4cHbVUwTQnrf
vGUXE/J1KPjWTw8N/VPb+cJPYa7Y7Jl7mGrf1AfLi6ixKezWPKSWBPojsUq2wlGx
58nBaOtm3bzT8W0gMrgObyEK298D/ifSCWIc74onNX8SEmG+X1/Z9w0K8KtFCz2w
678tYmbCxDgabf5/70sPYhJFQNxW3c8p9rX+ctGeHmP+EXklKnpo5QOaOcp2ERLq
1R6jN09eCBsC/dWGRhbAuw==
`protect END_PROTECTED
