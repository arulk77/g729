`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNksRswszdAyyAwAkP/5RpWJHMXsRnQj8ASAr5mTa9bm
J0CKQ8GMmJilJUt8FBNbNkohEB23PYaqhUlzbR9Qvhj885dqT+qFqG54cME87l20
qevGqD61ZgXbE2aMzL8T6b4OSVSbiIXNJk4WlQfuDACr1TfMREiIvcpjBOSoO/Tw
GYT4FdrC3tLv5EWiIbuLSZ+69m/q5U4dFYrSUz5Bt3h02SBeAutvISb/vOjaMA+v
2kNZWGU82FIN6X2gHkk/kY+JhAHyGhfDjV1WNVACcxauysY1NT0ks7dcgtBTQI3K
CHAKZ3m1DGv51x8QwhXNOLedzPxqsVin0GVWa1lHEAvIQIiehtXDas3LChMtgcBF
XQNRmw3YOut8WncU70v5wHF2thwhjbKI2jTjHU9MtoVHZoPPh9tlYmB88bpr/0BH
ry7TDfq7Y1Hiwt32iPeA6+dIcHjnHh+18m6NJuYwQ0x6klnNwY8sSBlQtUyNXEbT
bsD7bNNyxoei/XxF8s77Kw==
`protect END_PROTECTED
