`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu480A9creWaX0rwdhAuMGCMBZ6KEwZautAFTsj7gsYsTa
kZzByfeNHY9r+XUM5t7Cj7KP8wQ5K0DEIH280VbnyHCUkmfPF5oW/FdTmdPZdcnr
x73yZTHepzmlfm0mCZYCJWkCOOBqvDfNGfGJYvtScprMScWC3yqDNSpozomugTuf
dz86Oq47wyoxDAiv7B4rmHZogqUMDntQbGanlrfR5taE3yCGwy6OrBc6ar9V6oKv
DY2kdaCzpnMIsomm03Lesh5vnyvkPdtWbdy8c1kyG+rZggE0GaQjYTRFqF1X+yu/
PyBj3jiyj/DUXlZKZkLUWA==
`protect END_PROTECTED
