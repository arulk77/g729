`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yHCfITaMNOqNULTI/sKHOSKK0bRdlepiV0WXJ2A4VET
2aT1NReCHsdViP93+HjChnKr/IG7TuaZrEiQeQ/lcS/YM6/9gxvjLA+h+Spfp02t
cuODaKSJn74CBMEVaFo3uKPJn+Lkkf1GXbK2W+kymKm+x9D3v6jIa7VtpT2CJA/v
u166DxzeqDY2gGz8DqdnOD7ZRDRxbgKaDDs6St9g8szNmPpg7pfh/hxbnBsEd+xT
UAb/ecj1sf12Pf9jLIkN/byrsUXMaTZNYVdazhMXmM50kWAdCbijY1CpNKAePRDv
AeAqPjJuKtejb7CCAwbdS+40MDd3LppgMrsuKue4VcO+WpNGfbdZqlwt9Hdd1vtg
Mt8GIBod8sXGLtCx4kd7Ew==
`protect END_PROTECTED
