`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKRyZ5RfkjGOXkUVCoeoMNL1NDqcP5TV+On3UzTs3drB
9htJKDi45oCSt6pg9igX0nAwacJjlWZ1PYg3KCnUewNkODaXcsKM/zqSxXXqoabr
3jBPQVbBdJb4yQlHvDhuTnf1iZgGNsPnp3pRJlRKhAeegD6UsMtzA+NJH2D2XoF1
mS27gHgO9OScl8YYyVakYSaJHZTHrKcz/jj6oONpoHwBIZMNDDY6XME+NoSmW/yP
+yqShR7P/ubewjCoQoe5/wEXJu/IqCxl420zRrZPTfXtc2Oe4loG5OFDXvkVbaYP
kusqOqpwYwqzU7OEMXGx0bXZD9ELhKyreWoKN8P82Ri1JLxZHx2NgY0JnajvKqy8
dfZ4p6WsBgVaqoKSRwm+2g==
`protect END_PROTECTED
