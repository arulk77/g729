`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SViVc2L46XrIVaww78TOiTVP/zyAqEXH5BuPSEmKQvKw
zXcs/Sb36F8BU83Jjha4O5pwQYqqd9D+WHDaIisLCU6qZTn3QvYnSGzFYN2GBvUv
vJCMAbzhL/0e5QTrhI6+AnbctFUsrhPPF4+Z5Yswb1XOGUlD5lVKKrVXo0gUm112
2I5FpSzQeSNsJ5zRSdAYZDz1oY5bBJuDetDf6Wn7Lp8OnrwEg3FyLA9kHusFjCB7
4xT1Axbkiy6HHbZvbJ7dtxvnY2qsHh7hlZ7J5SyRqOs0jPUMTFQ0h7qXMT7f/Zz1
0nf1UpHy0tDyn+qKulumDBwczepyNLwOf8f+AIa2RPZs7g9gmdH5+GWZvFw9Bhwd
VNhze2UYw1AxujjsVxx+8FjNG6YzZ2lSgv4ZmLkKW+WY3K3s4x0QgKkFT5QL7OkF
7S6J/yOW3tSlfiUTodXhihWQWtSAv1B8m1kIQjK0F5tJAuYo2YG5ISLve8vPzPxD
XhnZNWOjjsMYCxveh19joHPXlLqTURpKCNOJ53YE8zp3gG3z1ArbVFd3FHKySbD3
8R5U/Gy8YI8D0p+kaMLoN4f3dkRtcTxJ1x7oEQlhKDVgPbr3Qunde2AbFfxM9LC2
UTeXWWfmZhJdWUNquXBGSe7rgoQibhdbv3aDaMpav1bDmjAK0xuPPJqjmMZ0vPtc
AQDLWAOJWJkpK8eCK6njJHFAjZdWiKLNsqi6+5HFyeZpOWuxnDluzPPcBAR+n5il
mP7co2KYVO6w86A9iUvy54IJYd/vla+TVlvMtqdJDWFucl84WshnT25ATIYvFVma
v5PlxRNGSs96fggrkWLRHIbnGW76QDvabaX/7EZjzjlOIYfWClYjWtjiMmP8sOrs
6qVd4DyO9VWUPzTh8dptaiRxqZIJnuFoyP3REfQkOSJ0wiIxUYiE23pqYtEoSHWh
SVdtR8TGBKRgQsQpAKmyrBitOK4hsf6iZSHpNlUzn5IDIJLAmrX52CvxNi1RP7rf
NuvwbFRU5+pRC50imxTQ2oWKrcgaKyjoFqrSXHR5u+Sf5ooxUf8gM8IUa84ij1wz
CZxtR0O0AtmQdJqqfOjFleVsBSBYE4ejUaf1PkGeKTwseFmrOz77F9BD0tvSCiQZ
fepWH89MRGdk73xNGeom1gCM4JmAoSa4nKMrzsb5kcPcU2W2WAnzw8w9Qv5tuQVV
/fV4ktLTrq1PE2TaSMXp3EGIRXV3W8se02BSxkHQ1LH3+PY/EwGwAR6zIuReyYrB
jyG5xCM7TQNREN36tJI32ZWnY0PPLO7YNoHP0PMSG4vIwmLd3SPyKWArSWx8RMLc
0AWOBP/J+iSqeZM4XNTvLZEt9JHMt8ePwKKtXKSwRrMmJ1+KTVO6d/5PGpLliEV9
WwtX78RAmXCwNaj/qUP55p/YlUrAXnf7mMy0HJ/3bppT/Cq8BU+OQ3zO/gsVPVFn
1etI5nx666OJUJVwGcInqv6Dy76ZLuhRWucAsICvTdVoeXLV3DsAyCZnT9K4BbHg
sXYVjdGlg5djTMuL2nt1e5OJO1OpZMC+n4nx60XaIYpMciV4Q/62RbTgSddTVQqI
/GC0i1l5zxXLf+e59XDGNLyL01Uo5T4NcuPAluI/yY9NzE3paVjV0VbSNdpdnWsr
8QF9h4Xy7DrO5/T1TaoyWz/S520ARdV8LeGZz0/rzANvjimv8hLHd5EKNK1swNbc
Tvte5E7KYjSfp77CkcHsEmi/LhThzWJKfa4vPB3mshik1Vg/zUjdq5ChqWdB7WYi
Zpb8d7Va1roeAnN6g4zVYXSAz4Hk2gwaMnp3YyYTDPITSkZrY2fA+mH484llvqNL
ehhliHsjz8xBQbw7Jx5pZCknrh4Ar+QWL2LEab+5tk5B7ziUB1PidrGGt/7C3R0c
iwbiLSkbwLqiQBW99Msp6Beyav8aayv2suTKz9RAv8VY3vZNgTGp+/Zf5nECbJav
uHi3S6BKTERR4YKMuaejrh5TiDGb0TYC9UVMwaD/kkL1o0S/ZpukajT7ot27yc4+
YLF4NSQxa7Gz1JQ5135Ub9go/WWl5TDBKgCV9/COhj6EY5Xb2HhcHlEOpcnGPMd+
fqNWRxvZ/vYispbsG9w0tuI1UKJK8KJP4CxyMtoJR+LjxUX0rY1NU9m95l6xTQqe
qYl8DM2JhB5zQZbbs7yIkI6NYx7ua8whrnfacXh+BfAgHiuE/842IDLXkrkknsHP
kjWbff6RiNYV5EzyjrvkPCXv8s4q/RbbTcImZRp0Txv+spC9xhkKWE9mJmSjEuK/
a3vEvnDHEGWaq92AuQsdCRER59k2Ix9pmag9OFdNRdGacAYtjRJJq6/8nz63k/YR
mIMUF7B5ZvHo43RqZSMaOofkBZdnyG9M3/G6J8JWX282uTKEKltGyh4nEYmxBXRm
qGgMkhzowd7cf69Ly684fneDgPk+6lU0J64qdBsn378=
`protect END_PROTECTED
