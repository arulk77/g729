`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEKTS7gHYDi0GdRjQJtnAXsNrsXKsRpCV73yrcEzNXng
IepW3dJv/Jfie+HCp50vwCB9Da1Uaowx2IPfyA7gCdBTNpxC0//0Hya0aI9VRrPD
4AfwAYeQMw4xKYLyk0+gSbcxAAlAuUSdEbXLjWGvsXQQKkj73vRvWVE69nnC9zkA
725oLy07ytV7sPSt33p9m/XyVaefu3acxZhQ2MvcdMPoi/kQQBcfZNN6boGQxUmK
sRCaiNegDITLHngsqs2SDgLVRr5/UxAlJqjUrtBWK5nugGbg9m1v1ItG5gRtQuCp
GH4v9BoF82vUNkwUfX1CKzprfr8yKf26RlH7CtFmEL6tqtbH+kPnx909Yf5rO8yt
gtHOS+GprMd9ksAiPywQH5E+oUXjQW+ekY1vnj/Q3Xr+/UXy65tx+6YrGCZTmlsq
Dz46u9IvCGCaarDwTHWj3/ubpE1S6MI2KfcEGz7U2681WRH6QZa8N26ReKIABRYR
bAaQHc36y/qvu1jzyo7DuKWQ4xYEnoBZHn6e+JDuJ6G+h5FkabVjLoHwEDaj5dhL
`protect END_PROTECTED
