`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAZPCf99stF4iL60k4Q52/zckQbGYrCkjfjYFjLojJowL
ddd6c5fyR3gs3UE3dIh2ylmE7G4spuAO790Ha7jEqV6fguWJFWIR4gt6nE4wM3F3
OOk6RRzMd36DTQzzNsGzqKiclFkXVcauykDh/xVzb5zwGHjN8R2e+yLso5aaZG9N
CjfWbX5rxdlL83tYmDv9Uom+wiDg2/V3zwq60yrsv6GmjSK3Iv5+3cjMqgGWUxHz
u8+9V/9nWNzqiQgYsDwSZ+AfEMBPA1rFErevq9ORweA3+KfHKL51HZGolMZRjsiE
WJtMc5MvnKwXmyvFHVU779Rf9gK37HqI5VuilFqdsYbl6zYuGEVTkfpA/wk2seuS
2XDkXYIyfEI4hkSyEKedCe3ydvoJqgAA+GMtHMFXW4GRzkvAZ95g3fhKMMpCkL51
J96jGOMP+fO0JsaOEOLTTtEn/FQjG/t4OmNlH2PE3/jGD822W10XwbzT0SmpSebx
Brfg/n1Bj9jaarM68A4pT4nRVtSDcZPcZ/MPizRfslG2U0z3WIjJV4ZFTBHKe2Hi
ovQEsOQkqC67N7fE0hpiNRzu4aeeQ5Njs9Vpg9DM/slCvxPj15KGZGk4sylcxdoJ
+GC7LP2dpzyWyVFTCgDBXyQKMiha404Wbwbi1K9q1/l6wxeuNBjLo3RwkWyOwJZk
7VIcD9EgiSnH5E0mOeFHAzP8byoP8Gw3CQ0zTY4gdNdbDEYhSuJCVJMDAvspSus2
vmPHZ/ObpTrKP2DhYAS4ia6MwrO+A54kXTX0NVpfprYFgfeKKPJ8XX/vVua516TP
pVBJrBTgZz/zB5SEYAA9c6NFeuIaMPEA3ZHc7SuWrXlw7shswZRUm6j1ZI61BB0W
gRqcClh7hejpO2a+5qPWJUffOKSUQu1gx60+CYNmoAypbBQA7E8SV9i3KzqdAeaf
6kGaVyVBwfCD7PV7J0IejOeTNh5o+BfIQtjlLMfEnbmauykHVg8E2k5yqOo1W9Ei
SHeO8qPOh90RNJrMxKnxwmOiNrhCPpbQjpcL5QuR1QlqPOF7JO/P5jMhwT7QSHPY
+97B1PyWt8T6Xs4c1+dQ76Z72JoNxze5a8dwJhEZZ5+0rvoPk+KRFDm3mzwaH7qK
kX0Tap82+lEWM6j/IQl2TuFheFjVZw+JB1AOyv+txyFJ7Ivwi7v8FL4nWJ+uSjrB
8p68IVHflxvoyxWdj5J1BisleEhu7s3E908ht/S54S7HNWzwTWRdHlVuuKV4uwph
Y5v6tvRCuZTlBDtcTgkIRWutXRmwycQlQHaQy4CDTu7Q4wl4ZYgtT27LLS2CJgu5
eW5ZPHTE/2iz6v8DL3vYkKVJHONKnQFddNpYL4Hefxf7GG+H+4tJUQc3HU3XgLzo
duKlwlFKV9nHzWP7D380wJuorr0E1dpRXUxw0MAg1yWok8b5pEcwaQmUfhxcREkd
`protect END_PROTECTED
