`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN4SKSxdS1T/ra90YF9TLpsXw1NdoeV52uYuskbjhhfua
1Uq/FGmClLO7OP/n9gmvSoM7foijJPEXriXd+n+wDaQ96FUmAPnrR6S12LyCfcmp
jk7+VC5fcOHDTrDlH88OX7wgKmDdHLQmwwP3D8luiHBnngJfuU6aUqWCnyRK676o
8G8EwLc+eIaQSyDdbdUMmNYeiWoS13xnogRHGgCtZXg0rVzGcEGEa6RK1xTRTB/S
urMfzCmXZvjq7q2+tLRgq9Dk+c2g/fFrzrP34zPbY34x6uZPdDdqlPrqLDPOkKCn
hE8wr3+LXD287WvSoqYpDu7J9vkucHnW3ZBPQNBwI9T/FFoKKuIvxi+zSINF8cXA
X94fK2f9AQPqqoiwks17ul3Eq0y/+RG/rtFnSAIOARVu+mPOTNlcQsQM8MBfj00p
H208aKS10g66P1NOMRiiuKcmOtEMnRlyNcNeL+XOH6FkpTkpMfK11i5kfzmzRsTs
OeI5V/5pC18DmLY/D78qmKZ12Jv5n7VCgyK24KMS0icmwFojmOBWctyYN9hWkUAN
ePjQrZdWNoyqTGleSUsLDdar1W+k5QQCdaMQzPlRyN4lEgDIIjA4Vts/5AK+E1/V
dJUye6HK/UEguzNUhDqoxSbej0N7mIN3cc8OM8ClSvjZftxkBFrFUgcH2IhgeJEK
DsruyhPIZaVobkjw/A10Fbuz6leIOb0ABFRF9J06uWWN9B5/3DsSO9w1HQrhKGE2
bqNYcUJve6ChQDVJk5Piuu0/1eJLxtuYlyP0doSnBBCcHi4hffSF5Pc0Iz/9/DKd
tbNhUR2HtYa7hq5YZUnTmvwzsakZ/OxRfPk2BYD0Sf7mpa8d6YXwMt/35QZ87YTi
uqLoougAwxlHnu79JBNeoELq2EcuOMNyOfsROsCSiq8DT/yGGKCCLw/A0hQhByyk
FAVjqHn03hYyqgSFLgFGcNBzeDRa/+fECyBEy9Ia7P/fGIyEik5nkSpN7uh0qBxu
3gVDDyaJfWGw/pclfzziedzlZ83ePMneeoTGKPEk5T8cIfQteEKf8n+6ZX10bcLt
BZc61XruKhNQOqOsEvlXGKjBNh3NDe8gH1TbdI8FxyBC6dt8aM4aw2BjTTYP0jQO
5bIZTrVzMuS43g8REGmnCR6tJNB9D5ByYLEfXuPAEzP/xnU3TNeDbWCL9oC34A/0
Lt1ToTZ9KHVaEmc8EXFFu4TKI4Yq5aWRtdyKQhcsMleoMuqkjrz/Ezi1EpI+4Afs
szBrWX/pMHpjhigJtvwHMXOndnIZIY+6qwqKrjrAE6I1HBkrxa7KQWm1e6v1dhOf
kNomg7LE7Gfednb0swz93Dfg4bKHbCEkpC/AN5sENcc7mhe+wh7v8W/eeKoBFMQg
I0UTpaDdlGKqLwvWEAr0iA==
`protect END_PROTECTED
