`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4036cY3ly4tfsHRN9vyt97UjU8MwAE4HC6AYFrMor95c
TOfF31BFNQMWmRoQqyEsKGo7C309r2D6bj6dPuLtGlLtFAnNPgpsf1gAYve8HQvG
ArsIhCZGM1vzABFlfJDPLNtwoQkWTfBxUig3bfyR9u4cqL5ZJipFg+j2HQl3ViC9
NNkxLx9PRrLAcfaLfEcb3g==
`protect END_PROTECTED
