`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGB1vyOMOr+ofeXci3ENWFeki502CEnOOfXtWdR4nweO
vgAptj0x307lwH8jAJ9aJuh9JH6H6fNKRc2DPbjRofKVjdfbB7UIRZK5qwtYSi/+
Hw7KkYz++tiarqKyN+R/Gj6viJ7hwS9OVuzjuSBugoXHSlKn05QFLsVD6hNenvzg
/yyLIMps42HZ+NKKitb74KKVKHzQgGcwkjkKqELR9uNN13v1MV5ks8Qcnp9n+gs5
xYTZhoDzcXL1OdQlq45yhkdZVuD9wJY8cbdhfmTaJxzdjUpAdMyIlx6TJt2rpJij
foLTaVNwSJweOQqxqwAQQu2lR5AO9eBlYWf6vG2Njl6L3ckNt/hMkdN+uAqSCfCW
vqZ0uIcfq6E3WjftCrWmQkIhnLWT24PhUZy0Q6Q196czzoeM3JSSsPydhmd9gms5
lNSS9M3I0a+qOqqY4Pbqwb1HXpsnUCTLrdiZz6ecMLA0BhRb5hepEgI96QDu13Xd
/JJMBnUEbxHNDsIRNPYtYVytDPmMVhzGXDPESGLO/xajX3Ri9z/x1RwcZc61Tu3i
S6Z+ccevCN4zpzydfDewlynTnmG+rZUAmox1DNOQQ+3nOdP0hoCEod3nEcNKymre
jf5wh32SOtoHAXz5N6fqLNFX1SqDWQtU9MRfNgVE5Yc=
`protect END_PROTECTED
