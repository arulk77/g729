`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
lXr1VGTushHRW+2M9YRdpSQHhhyi0S2Hdx+2Q6Mk/UIJnvRxSKPda1KUgSNq1WVU
SEruVhyVtqVKJcY6B1aAYDC0Hw87rTe/GfRhHUeaRiQsWtNiVoSpC+VAO3ww/Rvj
K8jby0yO4qEInKsqu1/yr/2jEsS7ujFr/q2N/yWQ5xdRrRZOX16FCa2fHPg8upm6
+zDV5ehC/Hqm9NxKa5y1Oq6QDmSRZWLsb28t7lDZgfqGuode5DsReVyKVMT69p9T
9Mz4gs/b3PXxGg3Vnah02qSaysXjfTKZE/J/2kRDvus=
`protect END_PROTECTED
