`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCbN82kX7RCQk9KKg168hApPuMyLITynOyd99o3dn5sk
nlefH0YCLl2aGmKKHWqUavwaTxFGMTOaZgtyeGFvfGDQAT3Z1WMH0K2RGi72DTae
Ssyo3R0ZzR85YPUFlxM3yMyl7Clx6zJ3u6TV7RpqegFm32d6kL3ZML6J1g+5gJSk
20meV2oOz0OfIN787+rDFyi1pENzW+fetaLg9ZCZn8XM7y4hRnohLxnXOR8lHBu7
`protect END_PROTECTED
