`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+1ZMHDJYKPswbfZpOIFIFtC7dPVi5Ion3q35KNqDCnn
yNYJa8Y6ihklqQnTsuzLsOMvmqWsWkkxa3Zn5fxOcOUxD88rpYkjVJ6h/DRRH8vS
8jywm8fRVdgS7jP5W4ug9Dg9aObjuOtC+XD78iFzL9+dGZs5jEg63eFl+DW3BmUq
gVQZLVl1VhLeRSAwFxCGZqMCWvpGaf9VmvnxazHvr+Mzh2Pgb9gtMiuETh6tBJSK
9fSBuun3kScdMEkNicU+bhlgifgDrcUG48oNPkOsjI7RRwN0HbuavUtle4iFf6/B
YXtAtEh3B6OVyN0awUSUvXKuGMUnacaaGT/oxB9kmgn9RbtV5vsAFYfGQ0kX9puW
pByfxX9jRs8xdOa3NqCpUQ==
`protect END_PROTECTED
