`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41nAxzyWoGh6RlGty6FAPtGBdFx+eIOV6jM40P2TkrrN
i4MWx1XWpA0SG5ZPug78cyV2yCv0dDdM8pLpA4dCDZxQAARZsg/p0znZHltt2/yp
fWzCJydkcD2K4/dRvYhnn2B3G3M81lhZ8p3gfiODaJYLI+D5VTMPcf0j94X1L7GB
BKyvqoK3IZnvysn40loWlaaYAdOhxY/PLmasHKSCjoJSfgaiRdtmSzFdEW5NrBF4
XqE8i9D8Lkq9Yrv3Y697PfZ3Y5nO8CDBbgzUAJwFU1j18iZcwlwmc2OTbMoFnzRc
wrIeOdgIg3/z+TgTVbSrxfU/qiOISL696l0+45h+LXUpJUAGev2MdDGrxLd3023C
AWcLcLr2Hv5ZAHpfEpYBnf7aizbqedYf2XKIdOj0BV32btZa2Vz3Fp9h0pB9eHOc
ZrSAavBEmRKeT3J0X4rJNxH4zyNiBJsmHATrFRmw15iL5uuhEQ6aWVwEvoyI9gQx
`protect END_PROTECTED
