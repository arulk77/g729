`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN5AY3F1lmuHotlkE84QoCj+FXzC2HzvVzLOnGlCJ5Ty
xy/xQ4YIFyf9zGS9BUnb6l4nNNh9vvRYsv1D5cPOnRT77VuJq4VOP+/ziO/30zxa
AymE2K1S6QZtFk0yGcexILcwyMOJP8EP2OoTPDSdJzMdG31SZ8487he2cWlqPLeV
JGseulp5jLWGoTvI3Muv8gUEFJcv0AZSZ2GgiYdFyjg8KKVH6vBoHdOk1N+q+A7k
95DbCvkAeu/EfoOudVIeuYgMywn31pSnWaH7WCxAUU6QTL6hRGeIw+7QraTJGWl+
0c1sG9Ux5buFrU7EX57m1Klt+Cl9tnpe54gS7v+Puzmv7f3whmTe/QEZPqMOjl1j
V12IGgOqIPHFht+ueevSupIxt1rjFV8c97DrO6Vw8g2ZaHZSOXKMz/E/n+NoaoRb
rj6ACSWe94HOU5HH1XHJ1rDa02zaJrbaFbJz1XGZz4nivqM03lDilRN41GSuJzSI
LKdew0LhWpES783nmPzHrIMDmVQ+ptF1RiyWYW1/8y/RHbR+OjyUfDAtGCQprL9x
`protect END_PROTECTED
