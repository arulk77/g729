`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41f1zvgjzQFlww/EveYKCQiU2KUYYT4DSWfaLQxk9dO6
nL5ZEq1r90KfQBkc1P975vFwDVBsIgtVVXdK487Lrp3j2cIwPOqLB0tKtZQGsg39
O/B2deNN3rucH10bhrLz15lMFg8WEflx/yXXAXQmIdaO3KUW9aXBAOw9v+MeV1fM
bYGRk6ukmwrjYtrPl9gLxXJ4y5xn40Hh2vRMD5MEsYMG+w/oGqQTuNBDNaOEIQD/
ZTKtZamIccnsGyBwxlcf8e31oB23p1Iao5EQEt0/BTpvAa5qDWYnYsrzPP/JY54o
Zrc5SIMdIiCHaJKlW4TrTg==
`protect END_PROTECTED
