`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
6UMhGKYoe6P1QhXGP1BB5zy6BPrfq7GhMugGtVd9TxIFNaD10TjWAQpa/mayA+Gd
Y7Xo2CawG8RKz5HjwRJTitp6N3VgaWnER4OELcu660Uw2xmT6hnXKOiaV+E4NFkg
DWzQPHtdRzux4X40rQKiBzhGrTNSEsH6rIszDYYxuihBJREXWWqjxPyBdpatLvEq
2UTSMsIFU/McABjj7aDaYGgQe0DxPYUpABTsQpLgCVIFMrICpv7CopA9Ttvibgqk
J5e9WkvNOpeQeTedEJj1p1LGy/PIU3lR8iRVuLwwHhtDVdHl8cN+hOltRzmD4BDm
+4IKbte3PBklw1DxflnsVX3DNm6qCb850n/5Ey9vzMdSimVREqnnhyu5LoVKb4hB
5TdGGXpVpWJpEiqsx7DagLr6GdkiU3aHKHHIYTummwTrkWKS6JqrZs8KKDRFEzSx
GMOM5I/lkDzff+lOsF99D7pOdPr8QT8dhb3ngzXUxEI=
`protect END_PROTECTED
