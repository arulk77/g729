`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
1IipvJZemL9h5dyVUsiiZco0Na5js4KLzvimQTDXytp8344i6dLapvpfT+EPjHeX
juNyrfUdhaC9O7jImWUCMhGGkqQza0+pU4W4fioXn02bBFTnCdy7hqQ3B/WcMd4f
P3B45MqO+bj8tMx/PaoOXc8V0nhXZQ7WRsYykUTqFQA9RxHoR0cMv0PA7BPgM/Rr
A4spEjQkDaklvPYBG84a/XqWjbb+puj64sB+88nxmWxetFp/nkcS7GdE6SxLjdOE
+rJsEpT9dH53wCz1ntlow4EoMrRpOpBMvYYvHdXvZdi0locxzHCSeuZjLrybQ9ED
CNn/mssBMgfY/el77TjBxoaBVJNorK7F2m5D99yARfKYE9u2PfKZ1Bnz5qos32+h
PvHf/p/tBwehezvN8bXlUln4octNLuy8mt7KGqzSBKBRGGCC5ua/Gx5fGBhBLEJC
Jc7SdLKQ1/JtenEVUXgrwto7MKu92zPms35swoKDgRX3Nxc2go2LO6Qr1HiODOSK
Svuf7kMR0WlRCIVyvIbw2PL364XR0UXP+DT16AgTXXBp+YEGYGJ+xK5dvzrc6/yZ
X+3A50GhT7qmE9zJc1O2HQZI1uJRJBMfcyOykKuD1d4K1kJRYM5q/LFiW2WbGe6J
S+oTJ/1w8eYx/oo1gp0XoA==
`protect END_PROTECTED
