`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNRCJURhzvvbnf6sKPa1LHlXO//TyvOj5K0q3DMdqkEG
bW/NyR6e4J/q25DHqBddapsYW1UevxjLCWkjxnhl2tTvEcIwGtC9PYMAlJM4oyBM
aikCf09umcwGgeYR7GwS7f3x8FaypAtf0J7xOlXL8orGwwAm0VwzHZY6qn2esd3K
U0CfjLaFbqU38dxDonFhMwKuyOZQd/73L9yPQCZ9SCS+gwjb8I1roV+wsBASWO54
BMjPMXQJxO0f0/Us+0dMOoJw37jFqD3MUAV0guPqujerDDb4kR0Pzp0CqJiMk5In
/QH/8kM9shdWYoW/0l1IEddB8rYP0mmfNFRbEVWP9OyJXbHfiXDJU1AB5GlvDXLY
Nq5VpUxtIeQpRKehcw9CSA==
`protect END_PROTECTED
