`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOJbME1rCCfTxtD0a1nUHPf2Ioqg/DgrsmGkI/WpIwPo
KlIvR9eA3c1zyC/fJGNcGLO4WIx2fjjW8u59zS7U2aT8M9JLd44QiQz5xlPJPQzf
6KR07DmQ3thH9sU9pjvkqt8EVTH49P3frWTKtk9Tfw36aiOM3MF9Tdv/BHtinq3o
F12pPLMNY9ngQ7fJbzRK1NVpgsCLm2ox7GC0ooObE+oz/DsUjpffS2Zg9Mf/UH+x
`protect END_PROTECTED
