`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGaRCt9JFNmWEn0kUVOrMWNn/lg8qn35iyBsaxIs3q/Y
2EXv2QfFDF/NSi7VqKNuvK7AJboIPWTE/aI925YpSsXAIJymGnE0G0X1lmwakFGE
okLIlcss0IbXxp+Dm8IEm5JFYs1gwIHx8Qsa2vShNhV7hq9Kh2g4Xd48glD4JcEH
K3DR4kwi2HjWF2TCldz9ue8lVTZwrSG2x1wLDloipmEUNyR4+KkCRkcCM2XvxDua
FvvlcLfZLK88AatwCQq3oZlQrqamRrWKQxGEcxoJrjcnEu4r1Hl/zvXWYW6s8WfY
v1Yqr4kZcRP7rhie8butcdgwa9/tPBfoY4TCvwS3R4+gg9Rss2JPs2yXaQWy8gMW
F4hgKxDaxwOnBLKSoc6xxw==
`protect END_PROTECTED
