`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
UMuz+0anZnA2cR3EnLnISRgbh9BCe3KC5SisR60YXIl91uWsjtUWXSMeUTchh1y+
TeI2kN8mIRGKUGkRdTtY5AD/sisp51jb4ye6LKJt32H8hAzwCGILr1W10bZbwAJB
JeaLA5G6pow7KfnLuKpuhPD+biqzCt/whL+TC+yZnHZkm8oF8xdnA5Oy6L5lbSuZ
+l96FWsyv0gQgepRLu7eyVL9018O/oRXslWwZYDD/l2cNcuonmYWuju1U3gI0PM0
hfGENHlT8uWCeyYGdZwvHaGMXjFpXgl3+DLGpTABD4kpJi2mN0HzPhLk8IVx1zot
YOLT3VQ+jJIhnQaBWNY6jkqb1/lMiGGrJm7Hl7fOy4w=
`protect END_PROTECTED
