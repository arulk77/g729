`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveByrfls8nhCILoOyG+mXm3iL1r0rBLcTSwd3hf9eS9fB
gG4M7+NmLiYWqfIzaaceDjJ9gzKeoeXyUmfdZ21QGsw65pnGPN8sVxH3seljolC0
7c6mkjCV6mN4b5s+MxQs3ZzLEYzYdahEOrxV/7jTrhB3AzUOtzTtTE2rLEcpKGni
z+V75opToe5H1gv1O3LkjsjiAxkNK+KfC3iUhMOlr7Z1QWmXwVFLIzmiHhHd6lAs
H2aFiOLrJD2QqMy5xh+0NC6WYOcEPw08ugKM+FXX8EpOJVb1Q2uI0nEohp9p0nyd
NvmPVuy0Kaut4pr/zLGMTJorJCi6gXv4u/evwZb5TyzLCweeOCQtRVHINx/RZ6KZ
kRAHNiT3ykxl4Y6rS96Km7JNruZIjIf1iyx/H5eOqywrBGH1nYdxe8tx3cel5eS1
RVgkGVQNnn8tjJnNnlO1/LDZhO4WlhEsPJEHmD0tHmTSoZ16HRp81h3os8cUKeWa
gwO0xP1mlnDibF1dCgfrwC2/DVYiZESBG1RjM+OAxZ6iu6HGItRa1xf34O4pfN8D
S2tUFmmYlApDpB03KFT8Uff8/walNG/ddtyKJxc+CUtyaNqvDFU1f568YyH/zPOY
W4d3NBcCf/xw72rWtg3X2X+RAWcNeVqqlkXJ2YlCdQRRAWvp2Embpmj8HZdVENjC
gBLLt+vCLhG4+9gi40M/MzhuxurAzM4tqJisKUuwsX+nhCq7qXwVf9FHPrjo1FSx
IuAEC+8CuGCzQCVw+lLHn/swjrsNN/6p3FiPh1HXg5Qk69mBfFVJqTrkEpwHNW/f
usEmdTy+C5C0uBksF7sCrtXLm9U4BN88+L6CpFR1yE4QQKuWITjxQk9ynvhEMtSR
XepqUxNcM6rcEC2TjHEZQMHLZlrBVKiI2NP+gB3FAGtsDnfOAmVxKfZtcQkg4zpR
0ir08ZYYe5JjWwDAe+Lp7rPE751aw2thYiVMrUz0UdvdMmDCpu61si4kcw5zX/0W
LU2WRlo4sSkRBuZxaea4QGxneeernH2tOWe0bVRRzuH7NNtlADoNkAiaZZHpGop/
gCKqzZwgQJr7q5khJ36UV4MPFO2MyVlpp+E+BnhqBG9q61cgoxiP4qOlIgNzneCe
EVHn8Df1sI3aJQKOhj2P5AeANYyhnOiuZIuoubhYPWeQUCi+lD+/DhT+FJ73NvH9
MhoGnbw6zFPysl8RBhwzjkpwGi0qvtmlXlm6QSFu+39xp0Z9eln9+JNcwluz3zT+
/xXcXgA0HQeJ+p8CebAM5XuvMNEpUURPbdZ8KbbYyN/HJQ/YMTU/lVXubxkzUpTk
NvUkzlNEDZaPsluaGdDW0mgPc0caCAntFrR5FPoup6RIDSFO3rF7P/awEoS4dZ0I
/cTk7GCWrOWdtEB+JWMkdDyzcpoR3m3ubuBT+WFl7vZ8UlJR+xiPCAHIGsnCmm9L
0JPFN4noBIxG9xW9KQAMv6371H7M5c2vnX9mf+Iv0UXUTN9FYo7iQxkNzwpUn/wJ
eJmr0w5joLfuGgGNsQ8XZ3ucYBjcawZQnBjITSHHLy2AE1/VOXTc8SiRQzIZgjHv
bkG4BUSctPhbnZHnK7okWXzIfrIYqbJweI4BDTC86vlP+pQWo8NQEoo99iV8KD4A
QAatdJPYdM/nzuMM5FlU10RfNdbnjc1SY5zFHrdlz4SZ/W889GBhLenzuLhmB4Zl
AwYL2nbSxyAbPYJPHBVmoSPrTf1GUdkp47YyNWhCazoJU0oAUymjrVhAnmiJUNGX
`protect END_PROTECTED
