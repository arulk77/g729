`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu476nqoFsgg6iBMEmxA9YsExFH116ko0Ig2l/10kzRpJx
5okvfiEh6FyN8X1lVM0AXZ7Z4jFpn2ImAVpzpfbYPpxFLS6rmquY3YzmNerKNifR
HT+j3JnVDYV513MiM/4O61UDj19DQSu6zCbxZTBndZakk3mbzdvZ0mxKkUsypboo
w04Qc+ZHFJj3tmjgEC/N5YVe1EU/Rgjf+Hb9Q7mPAZfgUEAsxlxPnWTKhfqtQA7b
xv7R0nd2UMLFkjhUuVF94n6wlsXG1Dx7xTImFBDvZXTCRRVoIUjqMt6GPNMMB2Uf
HlMHDbvQnQ4CTbDYa2vIfw==
`protect END_PROTECTED
