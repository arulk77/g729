`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBBI/pcccxtHeWJzAG9oWWvvhKcXFJRDGW7lX/GpNshA
j9YxgYRhYwqM2Dti2FYvo9s0WrJN1PVsVyxEvCkCpL0U9Sunmfd2U4y9xCvDMkgS
Q+f9RDFymda36Ns+BIXs089Njc+2xiA9X3jr/z2X7UBNtmuYlwwqbgUruXg9xcHK
caQ/fPV4ktZd5x2jPyHoF1MENtsRzQd0wQ8Oc7tjzG6moGzXWOoV1gHh9SY4jrxj
PTw/zoQ2qrwhz9MK1zcQB/7yrUiet+xztgTKZ+VfzySRdJbWZIUSi+Hgidosi4T6
RbU5+FE2BRYB/naUbNJFHuwNRo1wMbon8sFQTKKiYbtQANyFwg+hHPQZS1Rti/hI
EySGdUoTL4pVTFljHbdGxZwicUvURA0bwR421clRb11CUHYMf5gb9D4SAwdxavRJ
TeNOXtIx8OFpgFriMh2PySQnR2N7pqdVfIzS5XqvOhUxhd0XCcCqBir/cEK+ykCc
tQonWM4lSsfRhAPDs2qVK+mf6QvGMDrejJYAMvFDlGAPXrrMvdakBRo6XaPLZTFI
A8CQ33buuVy6SCpNx5oCYw==
`protect END_PROTECTED
