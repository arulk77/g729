`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJmiDGVyt8Ax+u740CZ5skABSnhUmezW+3kYn1WsPxw3
VnZWKlL9YrKcypKX5hT1nyohTLnSe4s0zCaBYe3ZS78YJJt/NmJhDNYSdlIEHi+4
9cvzn7CoHyU6ArtEwOnkHoDQZWSrDHSu1rp4TKE/vk6GyoQzO81NdkoLrq59Y+8f
SHvD9NpREqsjbbei+0bwx+y0avJra1UlmESv3fvYJCRZ75GEilPP7M94Q11MO148
RAOI0TQFWecyujpebqYxKnp9YPxICTKZP9SZxz9e6E8wVwsfJvC3uB8fq3W6JDEc
5KRolE4+QpNmxWUXwgSwU7jJ4cpKgzUBq5epQIhlGkPIqVWv8zj4+p5HqhOVqow+
BTnQhnYcSM58RT/AxkhlQkGeYdQLBMZeI8voRIf7c1AUNT/AIRH1Tlr7NTDmFVj3
ujpk6sr/9e90UM7G5A+jf/dmeR90WrQ0dLnvsksyCT6ncH4tNqqR5Imes8xynUaV
XmZ1NmTNP73K6rJ5GHpWDFk+DfsHKjJ3p7H2Omy/8P2ontzjAw1iCiwUk9mEtqHw
bGLmESNe5amVaCoWH+yQNOyj+n9VNLUl8puDDQFXzkw2tLikT9kBFLaOk/qrtEMK
CqWj48zVrXuWr+v19Ae+OLDVPNp8edQjbXzsGuhHt7pqTjAC6G/OqjpPuuRVqfjW
Ht0GKxzeLY3PeGNz0qhAzJ6K3HBHjM6sDKrjQMJA0Yx0OS5ixEW8xq9njsi1MZ5D
NXAJ/3vxgs1eUjgsbAilo51F4IAeR52/6ME3s83mF0ieRVpidAESoPE8aTTU5PZz
jQX1GIun7mo8agtnxz60/2GOQRLvw7wl0imFzPdyYu4=
`protect END_PROTECTED
