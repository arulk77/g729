`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yugXFVUgV30bR77HEHc4n/S2wGyT9wFAkWPqk6RUsAE
cIo4r4BwCP6d8Uh5dTtaCh19ZZNDIbGpq7s9xV08W5qq8+U/8sCaHsvrhP35zfdH
TqaQxnb7OT3t1nqBeVtLBXvcoij78p4kCGjzmrkAPWnpweE+Dif0xYAmvDSD3v9A
7gUZHINm0Wz2f/fsgEOKpNqkbbzTLQzhY33gEXBKzsycgiPOuiaT5KIgkwpujQUL
Rg2ZuF+KhCFH7OD4ywF00l7odBP32okZlr9M5RbmuSOtVaWYyTPdPlA4OBGLkLvO
GY6A37iODIHzPgQcgLJpNpg7gRpnqwFG6OoSmprJoSvGAYER8c2npnMdhZRgmZei
eBhf5IIlav1b3vGP4i7klMWn/2VYAUie9GGOXFStu8315FsayrbVj/lVUyYr07k1
fP3atpFKAvolcPnvKzdOSw==
`protect END_PROTECTED
