`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SbraQvBzm5XwvHjLSGSCV8HuWTAZAu4reMuankTVVRsM
RloFfKTuqqacrdog/hDGmc4xhoVF5AnTY8WZX3iGQJKiWKpPySw53Y/EEhZLC0TN
TV4eF8bv2H5EYreG770f9qRW1EyCPSXKl5AYuVcAh8NpVXsw+Amg/5HXWLiO7qot
+RV01oEgzsk0Vg9Nq33YUFJdPJ6JbHhvCRoeKMmNKnW8D3nG6AGyLp1/uCTE++IB
KjHdfoS59IlkNqiXVBIJHI2PjhJ3yEsb+P4Nzj3ddQrNnzmULIDx0J5BumH81cjD
XkySbitnnf0uWF1inwacHKyjyPMJdpBrOm1T+ueNB+txzs8eK5et3KZfTZLOTAnu
geHnxei51SGjqhbDQGMFPmB72UAKPBGaxqKBd/gyJnmGZoYzPt8BRJU+kAeIYAl0
z22sic/+xF2HIvOIYhfzrYHjEo2cvn8Vl+C6IJhXgKeMvdg1bApfZ1/7HAHJefO/
8iM11odCnOyVq/ZcNVIm0y8xLji6+GWx1eTZ7GwYjGM+AnCBB7KU2qnYHGStXGvr
nimL94XsZPNguKjAbjcwP28HIqnOeGrf2dOP5mnn7NXY0Bw5o5rEwnxGh1sbx9z/
fp72BxpYVkwr5cUqI1z9DlC/GettBQzwozkKKK4bEQOPRHpHEKVtPxIReZRS+WsD
25MZoAm7Fb/mXyHihA8cf4jFzySr0pa2OaudyNpONdyphx6PNxRFYG1vnuAMlREX
vYSGrpaAeEk0MWrRM/avT0u3n/SBWaqlFmZzFKIGiPtQQZNoWNs7bGyRsPb0lR9J
vQr8iCrhXRB7WmIY2SKZxZZanBx5mTvylTfctFK6GGIrcvKe2bUrEGiYvrph7QFy
WSYOLsQt2q5uHrvbWG7MCxsnc61JlX0UeXnVdD7bF9FqkAVbazBH6USH8+VHvkXF
pX3xfG38dKWbS2e5tBN/1GwosIT2m6qhlnFdIWsghbmzCPI4ZRoHTWEZxHWkxz6E
IizlfU/xItYw8OzvA3LkB1nL2rPu685o+GvU7zwcCl5Gu4j5JjO31bifO804t6Mg
7UdvWINhA/W6bvlm4ETbwV4zJZXmabdxqP6H9tV1xAR/XheRtKdsViockb2M5xE9
PPCMurIk55bvNYNjxhpaghbHEX0azqOV6VNntnCvFr+r8rTwzHYZNt3hRsXp6h8N
4ChrwK96IUsNpSRGJxBkWMHPJ8QQQ3i8ODVPao8Oxkkg+3NRawfN8STIiibT9dws
rOeeOOLP0hwoc0oUVzs/MGjgMo1gAFBOhpKcTgQvCav2uQdffG79yhJYsqZx0L9U
J5gcYnqYj03/BPYWaDTsujyIQeohcecviNBvdmNU9mb03C3iuygo1h14ZANRcpUX
CMDeBSbnodwwJ3nhF9tXqyfnQxt0am+QrNljJMt4CbhwE5u4B3jnG58vPn2VR5Xc
SkMZBRa6cW5hR1W4g56NYzKtsapoEz+5ShzktPJQEbi+mVawyMDQ+zzwkINO6W4G
IYSO5qZDN27FCSwCyLSwFODcBalUHYknfXp8VfRUGpy7Ofgtiw4k8hMyzrpFQ2Cu
w6ojncjdz/0BmatvPJOI57rLUjpCeKukIZw272Xz40V6XHXsDDYRIS29lFX9p8jI
zs9iBozfA6XoN6vFzJBiuOkXwv8mvlLlj74DIXYOpQidhXRxw+ga5VN9fQ6q73Q1
1cGHGxGkZ2xNMqSCi7XJpfy/btwVNEoyuHCnuH22JTmd7duX0LjR3yKRZp9r/Q6+
FXy5S+88akNE2sFA551N729vrVt8gNQAOA2vv1/fQOGlJ0Hd3GKlw4vql+mI1oGc
iaz+6NmnrcbDcwQWXis+8FVLQuok4qa9c76uFQZsQK14Jrdv7M0JbXAIK1H87kZD
Y1AbysjaGvVCYZfxGOZ8QwvEVHzFJvwZ9o1DjRrU+I8MLZBoiwrazoFCcYLidax4
8Dzg23NYnGT+tdlnV1/Ww6WkUmZHks23JZRiZFX8OfwlgqmV6BzM/XrRU1MmP2Nc
UtY8nSssEFtj2YWcKUQLPJQJ03GC9j5wjzOT9lsyav8=
`protect END_PROTECTED
