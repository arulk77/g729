`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLJ3mAu5vMKiLE3yKHJRsa/v6hc4Gm1ZrP2TvPgWcqoP
f8W63Y7rqqgyoGtJvziqAPZdPrl1XN5Gm+3CsfwMJKflIYESM4aA6/pgyC5JOqJS
z8EZCHvFeUCOkI0OuybkMWipVic24GB/tfLkLn54HTMYLoVI4uM3l11b2cN3I9VO
Ht0BMlMLl5hMPQCxrzukt+AZ/Cz4qswaOTtf9+fG6zHZjOBVymj6uqizuld1JH6P
FOgPue8uyfI1NnPlZKhsVy71G3x3V5V9Bjy2OK9y9PCJYMMqHWv9NmaN2DDs0dUK
`protect END_PROTECTED
