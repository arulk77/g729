`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
N3fgdnGqXi5j/ITGYxUXZNm6ICbU4P0nFYjp6gCJabaG7UkeDD+yHn7MeHuMCBvr
GY/sgveG4MF5cBPArth04SW5JQ5nsAnLrc+KVeRvg2Gp0K9HoAzVcj3K1LY1vph0
tcxuXq3DdG/gJgChWfdpcB/io8Jd1GLvu6dbSSXYiylLvem4nfxDjSBSYH/fKi5J
eOQiaVNZO36HGDGeLyD9cOhh2EJ/u/GJSx1gFZIgm0FpfrY5yGdvw0fgxuAJhf/L
I3IdctywhfXurO/wyxcMVJxRLhlb/fFRPLCCChGpB/iuG/z7NSBw0qOF5nLgYmxu
msGSA8+JLIiM9+JuLlcuQaSg7XKh/Oj1UngqIO33as0=
`protect END_PROTECTED
