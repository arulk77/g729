`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDn4u/f/XCE0YIb3GYkj+3pDt8icrrp0nv+30+jxHF/V
HfFar7Xj+c6wd9RkJEEg4UYPUOYpa2X1agigsCl1/cA05zmw896jOZtE+vlvmdez
evENOJ7toQfQyxCKYztFCDb+aZhIpe2bzqrDzH+CjjFxGksK04WXM5sQlwnALeyo
Q6AliUMyZ7O48yA7JNfsOysjH8ffDdc3DNgrNioL8yLZND+cDR69ONKHnwTb+D6M
dPKK5rb3FmPdYyUOVCygzrsJvy8f9HdS9ikAkqGvqXr8afEUdyCmJTlAurkneepY
ItBr1YY3ULEHDe+bPX7sNp8FefXY660MWAGkW/DXht46L+jaEJnIVBPp3jhcfMZ9
tZfKaIOzEJzOpNQ4fRhXpouhddSqd/2+Sgn4TElLxkq2EtRGpspDHlp+NdynBZUM
aDS345kkqm2lmef+DILUXT8vpu1MMY/Vp9Fj53iTlOCIGYX4+TYIMN83RqCJNGBf
atwZ5mqbeS2czm+v5vS6zVfRTgny1OJiTm1/L1u4D6IbbTc+k3xnfXyVhGj8Y53L
EXWf9QBqpZfXQszcgKvjp5aD/5NVua2dwwCcXN3TheFM3h0ZnbdBaKtnAIuztBUq
nO4piPPOJm41Q96Or9BWvAB0t2k+TcymxFaYnmEhDnoWjW+oqQHjKuGmqPjGhfOr
2zm5tTewK90lRN5a7IvBk5Kz2eDPFBeHkabcWoiZrC7BAb3sUwXHKQBpR4ZQ11B5
TFU8Z50DfeCZRqFrc/R35AwyTKUO3uCzuEaa1kvSoUE=
`protect END_PROTECTED
