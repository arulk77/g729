`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
AP4/dTkJcFWs/FCSEYml5BaTrt63EdT351OBVATysooS/4TJuzZIUk4WxRGYz0EE
Cly32mcEFLnEuBU8S+a89ybhBly/FVCcGV3Tfl6+N1iwN/2ih7fknisknoIoCZ4a
Bqs97VcL0V3Ml7enFRawTKio21vuBH1ioFZPcwegNg2gQtQdIfN3nlMmLx+dfyO0
PGj877JQCyI21WTvYh+n2/cCasJ+zjLfDLbmqLwtAr925IYpyFTFJN90nQTHOnzh
DLaIzBDOWvK3X3FQmvF6LFj/uSBPsLkizNnaojjB2/n/G9CHKDpg41ulqcLWvGAX
QQRHPV0gr1UVNnbxn/9Sxhii8iSB8pP+pedqCO1kdKg=
`protect END_PROTECTED
