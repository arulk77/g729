`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNTTEDLeeRuk2EVfKiq4KIJHhpVIEt0JSB84cUFXRhfg
ngwUIOIICdsXbcXEMheYQAD4oYixLjDMoPxJVB6VwjTAZHnff/cSlx0KC7Lcoczf
PAkeQvRt68pYFs2pISAXy/iICVjcd++ZSrOvR6IaU/uMVCAlNQgwORADcK8k7UT9
zDvFCzYM+kXbFpUY2PdPEw==
`protect END_PROTECTED
