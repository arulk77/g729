`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIeFI4jYJMiIjPJURFlfbbYFC4rpzs7a12v+iKTXv8hJ
viTrHwmC3XZB8bIMvpURZtIButcvhQ+LpV2aG2ISqYjfz9Rzcqg1ElxBgVoQL+1w
25vcKLLN39Ha9GY9igbEmg/D110HNwQeKDEX1lXlXNDAYImqnqvr1Y3nOZrVWTCR
koeBp8dJrflr2m/20w6/SegHb4Q4aBv0a4Vn+t/keI3Q7GO47b9AZYePrJckeCKF
zcblrT4bKVnt7oDwc7bufWpVHJ68PlV9M8cxpinCd/OLb4ltQihizYSgGewxXqiu
v5k3z3NqMw2/Zo8n4owAnn7t7IQna9anaN2yxM6PAHbfUNblUT8sg5o5t9S5RLiT
4xrpFrnBGsEgnXlbjuNBOGspj6LbAUAwtvcpfMypUDA8PBoWuY7ARNyjfMQL0lPo
u1w6BfF+aKYw08lyzWEA+1Oxf3UhRjtetgfeH+I9ZTNar1cWbWcXMjRqW+57WSU8
hnlO2AtXMBtu34KDEkKi/Fxz2/Fm1eukl/pHQuDMTZGjcN56ijLDox91OTWRz/oT
`protect END_PROTECTED
