`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/il5BEg1EQNDUi4TtFkdZizQkX09t8rbkSrCYczW8b9
YLblvnui0X0zzw1AFYFIuAq0LnXCTnl+vWYmCm/DhMTdtb8Y24V5wTpFf5w2Bx7/
1blSHEfqs+4eqlmJVjTwHmmg/sGfJzIaG00k22Dg/kl41vxSXcU7UerMe7rF2H62
KBDq9VIkjWi6m/Vw3lwXu56/ihJWF6nOOApuCWbeLbUcHakXDYrGINxoDHxTHsQD
H8DKCq2YdP9gDE0VUybs6Wn6dUFxf6AqTU4L4+D8KT7q3/mzNzJ+CnTV2U68cDIE
2/52JnbqNBhBiI+Y1Et+mQ==
`protect END_PROTECTED
