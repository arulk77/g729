`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4gBThrY/vXWVM2XJo+KtgOFZxiRe1geSD8QYMMD4NqTli5sV/o2tYNDLnAyUZRjb
KDeEhUqFtR09cQ7E9jAt6Rg0D2A9HnfS2S2RhOHJugxjVKiQnL2ciwAUnWMBr1Rz
pRHUn0bkPRyrAeOa8/+ASuH/HerbsEy3FpMphUHHCStJnZy24VHPAUTMM78nxePc
NmFoMXsHeHDKzYhLL1dKeU654Jsqio8tqerDStHHrusKI7c53D+qxa6P3JpU47gq
jTjxutPepKeTPGuEPQW3mzn5yqtrs1Y+/zQ15T3iSL4+XFVyjrXpQDkUW5G+5fFK
SiQ6zJFF2dana0UoNlxDT0tFqAKoh0Ux0wuvOg8KJzmub0JAZbHXl5amEXIlDRa5
THJNWbUN8YQ+Fn2lyy882fsLmPqcUaVZ1alAiw3CoMAGZXdwYLbbkIak7bGZjNhr
gWZKI/+pXIPERD7VINDQuW8GGprxHMPJV0wThHGBaK1ap+uAnLUaHSCppNMlPSq+
+PtLVF0r7BTplkkeK7Rsc80hMGmJiYlfUhbwd37Nu7PQhOBPA1yqgrK/kkXudlEn
UDn1BAFIb1Z2Y1FamXEt/fh7+2t5Qr8HKkZpO8mSENg3GwwHaT84vOC1Bby833G1
vlb5gynoJbjvyZAUsoFIziyt+P8A0CcEmNQ3wd0yQ3IZhfFWZ0XDCDkQwHe/EjKW
rln/HhIe9b2IOwpak6nyzolcZoYeYGjXbG7naYy9+IPNo1I6VWfkdzqJ9DaA/F5f
FjSxy5LDil5makaw2sQtF5MjsrULk2YA5hUfw+nuC5M0dmjUY8XDp4dd0rNjy9+f
LKqlLooUL75Bg7tItTdgC4XvDv3GtFByWy5wQbJriUy+xWwwbR/sC5v2HwDHfQg3
un4dOh8s3DABfCDtJIJYzurYlIN5lTFsI3SS2mBt++NVh8+EBNu0v2gmvjAtGBlG
itBAqq5sRkSvGfQs1T1zQfQii7WrXkbqJ4sC2KYxDhGbgqfseViF8V8FG9Sq/tYt
Z1h/CjaDsVq3Fj45Me6rlLvr3m6/rpmtGJJADnAVurUkCh9gtuXhWQwLQ0BlpwUo
tj8FHm/9YK6zB2eGoXMSi9J8AE1iD7MZLFAADXdO2PjtBRbBL/uniXp0DhUbCQlW
hH8Ld7F8hm+6CzfSaCB1ciHkiMTEJF9Rdv8sE/I5XvIkzXmCSD1xXCiOthY9szsV
Xhv6uXNj1Rtsr6Xb+/2seRnqM4Dbe+FAndDzuZoOXUpH8/tC9bBtAYgWRogl37Yy
WOm4m12CSiSYA1VNMUT7LaeY7i8XUUUbis+iJSmlje+oFAxtHcWXpWJ/FHCSV3Ca
WKi0xyoOs67RZQuexbU5BHnDcci1Bb/7nR1qZN2+hQ+WPTr/ija7U07rQIt9UDGv
vb5zPa5wUojWnx+wy4v1FJqzFwNOgv4mwfoDpIfkbqaphebSIHnkg71XjL5RpBwl
Y3gccK8H4eY3saY2wUImF4ZzeVtg0xDrXyh+CyTNl4JRgRX7z4yix4NLjbdvlEyk
zXDfxQ5ExQcQMiBmdrx8d+q5v3k1ifDwiJ7Ed60hXba52Fylj/lLJlVSAP0//5hX
uQzeWp8+taySkkXuWuYmqash1UBvNwH1UFfJlAXO0KgDMJVHmYKNZV3/1oBwPubT
1S73RNQFe/PXOlHDi3Y17KeRBrTozhWYHsp430w8plwEqIIu1gFLvmpz9xHA+dXj
VI9l5ugQ8O//g8HnEO5gGPwd0IxrRtfwaPMZcN0iRhMJijAv2bL9K9y1NFS3x1N3
oBwAShmdVRt1X5nSdkMarTySbZ7ftBRHWdD+VmIIie18A3uILc9D8mBjQ/++24XD
/Jft0qozTr9oVJUYbXjQyLSsDOOOla5wtoB4Zt3UnhZKCkpuD1yO2swvzYEuPDv4
kwxWHTCeGpt9lr46lpmV1Ecioxx5PEfx+QQjT9J9nogaBOZ2Xyw24pdqq9EKhl3t
oa3mAtHi6OPrbYq95pVP/rpZQt4jvyndhKxHCZzEFht7FX+RGZ62Q/8v13GetUou
e6wCXBkt0M1vaZtGl1GKJ40OtLrJwf0ELezqoQtN2huroGXMgTmcP8brW8ahAeEo
XUpdQH7mjx7qDb/P1zSdxL8tsDKIoOSz23indKiOMAQPK00YTiMzpfisuXoDJtLV
CFkyuml3B9u6nsxj+KjX+aMr9RSGctZT68zrd3JOHUEdj0RFBpRO/ZFeGxMr3v1v
CPMo4HrXhQBUR0pWJUrC4xEgehOKZ5k8l1aQHCcLtAjlH3JB6zBnyjIeS0JwtI3s
QTiptrwURNwbNciYYF2Zi12pKFNDDN5q4E5WgKl3IyZccHEYpox/3pCuNMkvqjXY
lbVvpoOdXvV8ZYIbZtQUYsGzwDDBoNdyWSJKhqldMdeVkEPirKG/7l3BnREr+ucx
g7bWFX5W/1J/2EapI8OrrkMfdZ4cdhMzMRWmBQcfuNj04po2BAuOFNdDdAWMp3ab
gYFt4hoZUJH3OMXaq+lDcoE3qS8vZBS4SAxo2dm0yBCBj//YdLAouv13gOwnhuqd
JOHW6OZtNQq0F5laXJVR7I6IhBLwE0FNLsvOE7oId1O2FGgSIcxvk9/V5JT/7jZe
PVvmiCDkMyryM+uH6/AY2KyryHlU4HmH/HIXaw4hJDHnAO9k5GhwDr0RztRNQqa+
+ZbD2jpsxlNPWSwsb9F1x8XCWyv8LOpWmwW7o/7O3kzZYrR/x616zvZmV+nFe4be
A9/xAJ3DbmIa5Z1ip1lJpmjj2oj+V5di1g856UyoB5zED4CvaEAAZMCYxMu2jN+f
HDSz3jcXLAXmfnZhKZhtiXha8sHCNjMx/m5drNu3StBVKXmKQl1azZ5XwryMlTro
3/5xEH6dVLIENvJySLp62Ujlt8zLp0h9Vdi5wsBln+/V7qIzYUXySlJTV8npCyng
BzxAFxlXDSZMgZLmriKXdSoOiKw9Xd3hPo27FWRSpVj/ZOB4hzs7ca1qfrpvaTw3
q5raSUwCToii/rXD2GnfRvRu3iYzzmXTEI6y9CAxvSr6QUUQx9tUjpM8bGpYX9aL
FOm4upWiLIUgwCNV7G4xNDjvP4Mi9lH3451oAgGIEFjTdxktFH1sg4/yRlIvXrhF
YDtD/v2cGxrpThBbgRRYPr/+/oxfjpLxyVs+0GTlL+PGJxp87/PidrTSxK7Kmatn
vNldBrYRlLdsIIimcKw+Lj7/XNs189gDy+1g4TgTAdMRtUkBL/0kODm4fnr0c2Do
Gog2RzBN26iXvcYZpf8Tg202GENtLMoc4hpFQugI3YbCsY9X1L2kxrTP8gDHoq4r
fVj4tUk3LejqAa74aofhaLehY05jEQGhGkBjzTqGhXbrln7kA4/TwftoOs+pWze2
d/pfFsJUfU9JfAMVZMNfDYHZSymzjRglf0mtrQvYZHfoxfaPNrIURGmM+rZEaxhC
lTIgq4EURdoPzVDxD0CiYW82nFDFQNmh2ZO04u8iKNvKADf4vashufD9j3YRWTW2
/jHlW2VgiXo98rzpbrSG3FAWjm/7Vxspb/K59KdDU+3PJwiWKe/oGL2DC/DiVjbJ
Xr3WOt41k4vDIutFyCGtHovp0sA9yckf/+/4UVOcZJdI1MarS40lhG7oS41YHTqk
OIFsw25jHGe1IwKLgjbBsaYhW3PnTFqV8nMddhhT0avTO/ZiAIUGgxbJtOVkgmzv
AbKEVj0XKp+VneXl77T85aqXRnvCppJob7qMas3UwHWoQtpnlaeR7JVsNYEgGd9G
eWD1PHVKQTIP0lM4NAljZVWTbU2j/cVnRmK2fgZvtybvhtjyTPZ0o59v8fbfFXXg
Ao7KFnjGHywOV8wLO724Xesjjf8iehFyr/Ks6NCo+CnktZjWBFRTM1VQBd+gyZWx
s9PZIFQ6bv5GFnG3DHjDnLj1qSuM1LG0YAPHmVwExk03YROzhIk3u+stKULrvwtG
e6s+tK6OiCrw+9H2S3o7hkL26KTN4+z4NKad0tSPnOZL2BXbBPAq4xMmq79BlEFZ
XdYKmcCbiMzSI4j7uM6g32NE2ZbnwFGVb3x5TcyiGlS/q6WEG0y+qULlhkVF321j
90AN8BGwf7lZqb6uIDQ5XhHOpFO7N6Y4ZxPkYHMA1A2tu1pUwVVM95hxP2cQtnTh
SWk8EWDCMsop9oer+zYtGxOQ8Ux2votkzyg4XiMAtFSZ+VGnoOVkOLYTGjJR3wA3
1trmzqsmNTpaTEhSnLF1GUL9uYQxDh4dK4lLvC4CIwvPj3Lkp8jvIXHZkKJRbDyB
lBHtnq2Waa0nDSpnw4izho+uINwebg8+49ldt+GCGCgLLn5vIzzbO+8jKhiWNu+w
EMsX+wp/vlymuRqvUgW6P9o1EwfQ+0ANYpOkvm5JM5W6S4ptU9z9sX3R4ly40ha6
/t/CV1v+4ktqQnSKXmf88G63Z9pC1O3JJHjvJ6qPXOb9GaiQc08eYojhf+pZ+A+Y
7qPKX2O8q3Q31aI6vRJHyVcYYJL3J2+EUyPdH3FlzYe1/qCExuDpSgeilO52bMvq
YXoKF9x9/w28kumXK6qz9CWJCmTrZ89Hc4IppF/imUtUQ5bV6nsuc5+hPyP3TvGO
Do/RjDx4L4ucmnbXl2wknyN+Ief9VngVVjUuJmSpWuCexXy3CcoaiNYpwEa3WhkW
65EuCv6pAOSlEmEiRIe7Y7Vvw9IbNUrxEe9vsvmyj4CvBxVP2sr3JZqN+jnculKQ
KoAyN7S1TdkQpyqG36wU8OIKdeqMG+FcwU2z1SbgeIZrd/ioKgZnouWbu4MPijiJ
OAo7cDQ+ns4gsdc0wZd5Fku2OX/JDIHx56h6ujUijhg1K82s8d9UEv8edlwkBShO
Qd/iGuFRGlxCWUfs0lw/0Af8ScUV+gWxGlzN/RyZUyebGnCV+zlfa1x5VkXZuJU7
oRu8xsPWhQza/6Gt84FUTd1E8NzMFeWrBpw1MmHkVpal/79l11Fj3pSzIK0AqouW
A5BybCAYdSYu7HhXUGWDypq9lyHV2k0GhVbuMez2n1S2jyEdR5AE7c/TujDD0+Ye
ZK9p9Gn9Ug1r4UMfPUSC+QbB8iqJ0dKRsX/CwS+4LeiCxjuhmzLM+CASmpDU0fyc
tFlBrsyX6x1Wc58p3ADS8lhfuJv5nZE/PmLVzwNlNq9McsVnw6GX0x8k+ByCHAoJ
mEgGBkM8urUFE/bMfF4vRrhJz7cV1MiKNI1cc17aLT+nDqNpqYFfB9w9qsnw1T07
Msk/4sznEQbSvjrnwBC/hyEkG4ILzpIeV5Ub1ocqeTZUuRJenVo6KBVb/9RB7siL
miZCEUKVUVKQ2Vg7ewtnoCphxsyroUupQlOsqfFYJJRJSTxDQic7o4gWHgqX9XxB
D7pxLmGTFJoolDVqeo782n2nWuYbkVxwQc1eROSJcjodWgvs3Y3vtypO54Mr121H
x3ytCh01Y8DfYE5tSWBQCTwg9K7mYiGOfMhlKL2lK+Yxl68+Q0s09lwWjCB7OlD5
IbZWKSk2GBLyozpKtiaEWUJXM1dOS9/e6RN8n5FotVoqoHLU3427KysKCiAwHgNu
gikNSv/SCs/lbT9RqDWOQvsEa+kgw8VxT8Sm2GtOSrqykD5SvTOw8plPAwXvs4lh
nC5vmVLJ5SfAiCIN6E7FhlQ3IPMn+00d1IN8UosF1y5y7onQ7bqEkxX26chYr9d3
N0TRqjdbtAq+nb07WaacRfRpSq4ABsl5N6ljBxcvKgz0oxwPP1S8M4VqY8c0Os1/
AB5SvDN6retiI0gvhA4ZnFS4rR/sq2E0go6VSRcXz/6yDx2iqxk7lnsgmAb6oHfB
N+UsQFUHMdhIxkmwy7IOUBiO9ucyUDvrcVA6uyUViggh4OFwpyfHfN2KAIRw2Zkt
7xZAzjTIHKJGCxskcGecWsqEtPxy00Cm8TLOGh/PlJ5LceCiAePm8sr1R4jJT5sN
iXlYb6Jepf16z3ilVaCCvf24s/FgmojaBtGgnhS1UqNE3rohvZmGYBhG182aVOHb
FkY+dzDTAe98SBR7yr+EZUf7rPXkgTpnQX6xwtSrF/+0YftXQoGxwe22gWRvKNPA
yRuEwtXT/EDqKMJzQmk11bcJ0OnkLm5ZccKr1B3Wqrqf9st8kHBA26LR0d5q93LB
pc643LBH+dvnkTDQEtRgm1N2G8+pyXxxCaL3Q4pm4DWX9PTJmdyju9m+W8dRPsWS
WIz1PLdPU1aMWrjJ7f2ZV0btCsLNUt3/5mBgBjRd7rxVbGPrBhlaO9JUjWuU4XjJ
er06FynsNLzeu2kJfdfT2cgo5bBPo8GQbwLm/EXnlTY19rASQMCksngwNS3HXGBr
NUt6X+qIataLPvsFAhumrBrRtcWXkT1Hc3ZMSZ0lNhnnebQrKa6gXo0jINMd+nQn
A6jOdhCHU4D9euOj8uj225XF7AkSwaMOsXmPCIln6Vw/+NcWaXLGjrKz8rTD+TOj
Coko5KeW4b0dVfAcEutcS66vhnfoJ8Y6VNomB4pw5ivrXb5yghXdGSoVXBwB5XK/
mb6pE7+SNG29oyBoleCGBjlnxmWUoHKFF9OrufHbPNMLZckhSDE2dI6t6PxMBzqB
PoYiWIIZdMRQDAwd+yJVJWG3H00JtTFgRrn60Mh29NDr3awJXcm8frl//fUDHbdO
UlX+ew0hX0lricWTmgxIFqJ0uP4IVbLU7c1aEQDPqszaMhaCSP79tQo/Q2r++OmM
A2aKHJD7pPfaik6LHSSOzN9XrMhRWBQaoB9IDmxXaPpkPHbITKsHdPsgNm3ffEm/
TLlX7M9JEy4seJ1/4+cNGvn9lf+tw77dJ8XQhzPkCJMaDbQhy3IW4JDqPXmDBv3M
ohQjnH9ZC1/t2eSUDNDlMcIRc8UGpZiHkxwL2WGapVMWKsrYnhrUjGftwUl3FcCQ
+Q3BDHlvQnzxjxfrtNmREk9ItgQW8d0USARjNoPKk5qhsnqPgv2tOxEFGHhOr9R/
jpQEFUAlNqO4Uoz05VVLNpJkYapW4rAt5eQBlCyl5LPHGOfiBNmhhyVrFG2tB/qs
0a/0uIdwQAKq0AkFVPsAul4zsfcxDXfgkA0i73GKaI3muwtcX31Y5roZ8RtDT/q8
Iudxy7xpEKbYOi9xOdXixLIwNizTYuzV14q73afjhy5QIAIVbYIgkZyc3YeCe11D
q2s5VYZ5uNeAjtJ0JAfBuaFJRV6UqDZZ8TIgeaOt7GbrJIRJu3Y8cPfV2NDenRs7
V1iHxHcDuFb3ANXQu3mSMs5+iYM6bHH8fjxguRuWkezXkpn69tO7x1xyq1EfCRFm
vAgtBs6FOg3XFNlEJqv23QeedX79+TurlEunh5Ok8z2WNPURvnSteFxifnyGs99E
NpYePErNxctW9Y564f8SDcoUAvZoOx22rDC97wN85d6rgAI0Ji+9z8E2dZFStgJk
WI6lNjlxMv8I7IKh4k3LhkThGYe+BJCiADWuayMbrjWthweEfdViDsA+15Q9HOA9
/ATxCk634e01MzJGU35ex8mZ2ZWvQUWohT8Sxelb/tlKdn5X/niCLRcKqg0N1+3t
4lGozc1rxEvGwiLf6Szu8zE/alUdwO/GuzMfuM7fy68M02DIOBfHRDBZ9aAuQJhK
kYI57jeQoQubHOCoDhhwNthPxtEI9BHUgFbCEudBGJGbFqLkRslYk/WqtAsak6SF
Yz8UTuzrRLSfA7jVIayA5KUDYewLJmpJmOcA+Wvormx6Mt55gHiG1eSzv9nsRZbp
9Iu1HJgsYnn1FrCJYb31+3WZzJk3oPcJPPTkIsCnjsCjNOXmuz2+RUUJlYqO8Aza
qali2DYwh2pT2jfNkEq4pGfc4jRUhV6o99Veh4PgNnmTwhhHYdNVqNbmrK52SKAe
3+icxDlXgVb+VdetCiJ6OlCD6rGGERC0A3quqfXcCe0r7dsBB6lFB5qDc8qs+JdC
bgM1HzdylKdCvHCVrEoujsLSdrpnkALU7jSMCUFq3bg6/JAdIfPSCIbH7iR1uaXZ
p3jChoRxGefeNhnepEUb8WeKcxI7thF2k9KymwNxJyCiKFpRqpuiLO/NPc959Jw2
ofRrhaAeg1IYE456yQYMySlgjFI9S4GrXTthYv5y75ccFyX+mPoKxLtf6VymQOAr
47c1T6nuo8Q/BNS3EaCNa3C1Ji/vJKKO5/qCTEt0PcO6W3ttdwjP95LsmBRO/jhZ
rPZ4iTjEX/GNy8MVl2smdOGBpBPACGRZEylEAJR1JKPCoTDbhF+oi2yyM3IwepKt
yiLfnvcicqA16v1LmKukBmxyJKHHGr9+HmUWvXiu25sGmmcn/c0QaypGdpgSNXLV
tIOGqEcz/wM6yruckHTMKhpSZ+0WnMZ8qfcG8eMn9BeCo859TlxOlGzZi4lHZF/m
Et+Hq7BzTGZRVRJwlG9GKlaGd/eMf3w1PkjLdPwiSTWWso/C1ixiPkyDgTshNLZJ
7ztU3+rCUtC/CvyvKRcEjEB4e15ctPylmHP9ZGNhzi1Jryu/iIAppKEdTVoJDD25
1ELLFvHayDn4+3Ih6Ms9NQOjoSZDjCd3b+sxM5gNNLraFIrEAG+LlEzGRQwBjh6y
PP7EHT+/CpdwEEw3FZP3uuWdUDEy0O4/28FpH75mVIaSFxQt84W7/HAHWrKv8Y50
zV3VrE9bwjGaDo6wY6qzPplUycb475I3U8Hzo45boTc8ffl2pVtFSaJrZcOjA47M
NrlGsDu0EiDMFBT8HK5A9wTcO1ic5UpxAIXn2UMokEY+iAoDCLV26QuTXEO+nZ5z
vCdBOrptyxSIbTisKa6onqkYAX0iP6RAx2X4ZvZBpKa3Vhpbe2oILU6Jjm3Mrzqs
x0wpq9vpe8BdhZ14HOmmWEY83N0KdnJL9sQfeQLwDSjsGiqc17mhRB+/xPaPPKpz
T4AM6Otw4x3IzwDlfcO6RwullEW9++Jd8pD82gPX/ekc92uSrD+uLwbK4YkI5xMJ
ENQ3imOVDc98TpbHdT87nIj/SHfIu6Nj2l9o9MhilNARax1VsMyPnd/d8Gk+Jv5M
3LkW2VCoIwd8Yp6UNqYBFE+ypuSQz4LFzjOEZ3aWzMffpVpOcUMzPUu3qfRfnom8
5tNlmWxTzAvNRNjb6upGElT4H5l5SiYok2N0XABQWEpHVGakJ9loUPZkZVPWQ7aJ
+DORYOw3mj1gKrBBuZrRAtDwHcD+6MltxZzhcSZ7Nbc/dexbaMF5LYFmrOKf8Dpd
ccgjXNsDi2BFUJJKOiXL07d+3QiOAm5GRnr2WM9bRoAO2QjnKFM+BZnGm7LykJnN
q2fQTb1FXttZDQHXlYi3TtGI35DU9N7PuRRQDw/B4Ep4Z9GcZJceidhDtkNRILk7
fdQh6ZDODD4WFtU+WmlK5f+o7L7c/xXxvwJArXrkJE95WjYyWPT9vOVNTbObGrV/
n3WI91E29aXXHGzHdURnpe885/t+UPnv2UzuwJfVGFgVTxq35uNMfQg8pRw8hbY5
W/wDkwJFj0QNOEwuLhpINcF1T2kADrKT5Gk4mhCysTrTsgg8amOwMDZrugsszmKu
TreJQX5yd1G8MAJeXjHgJvMS+QQVdaaQTjnYyJtTeHPhUGJ0AB4can8qalZWjmWh
fXOmP6rtv/TPeFEcKcTGHVWh88DY8p3MCW//WHL0OtBjVSIPlvXmYWrCjsFXjibk
XZTbDa+zJLqyWVNZ6s3rABoPDZBbch6whnS6Mt1udIdVPyLZjS6v+mtgjb0mhNAW
q9o4UThJeXEtrY0r10s0ZHMnWq7cLdahvpcV0hOr/tQXzUL+bqzGeriTiMeY5UhW
m5oIREJp4DlKjCgHM5CMcKS6qdKlL/nLxHXLolaOZm1cowoiwDcCd1WjbJBvb7xw
kVyr8ZNDZnjOXpuKZLZXdMqmVOivKG2Jb7U2CbXbIKk4CLmL8PAZvELY+FF8r3iq
GKb26qzYIvAFK4rgZha2KW9rxO78/7DG2t0U138vUGhq/sMHfsdLDZM/WkX3EATS
o4ic3g8KoNu/s+42r7pr7u/GgKXxJuKg7Uv3quAMYnMJWAlwvXF3QkpVpMYPY9pz
/8ejZAFrkRqbbG38e6SnXkB+kyLhtqIZMMgMCZLnChbyBOzWraF0di+Sjh/2XfuZ
MwKZ7/ygmk8NCdeNkXDbTeLrHBSJFd9F31OgfWQ3MUj4xcbvfU81/VIE0K/yyfL3
fzM5w/YzmtD7EjwKYDj+Oibt0Rxb7mjIcVU/5znJh5tquQQypm3tJU9ubXTTuLdR
F4HkW6zkepQ/v+YOI2WwgBwe1Cyy8CrlWZFSibqLg+FKwGi9z/xQHUhcf049Di+5
4mJt+bWZxQtdjLTap3l3rHV1xS0d2UpRbDadpoK8DnsgEbA6dvAZtpPtKwgeEfBh
m6zju8X5CwKV491aSotEE2UKK7uW7q8BunLPdyrQEHr2ya+loCzqTof4hUg/UutW
SZxyHrLeAI27uKBRHKKfTcfMClCOBG285zFexhROggqpy/8TIoR+HCvLfciQAVI5
0RiZ2oMKfh74Hjm/Vn0XIsX408z2btiCSs7Sj9Q9qxOzGm+wSHfk9zpmoAuh7xiE
Mv6EelOTvCJ1nur501C51tRSPXsWISSH/mV8Scehi7YBeP134rkvC7vtzlY2wgFV
wDxCm7rpg4h3J02B1DcQCYwTJI+UoDY8+0EEMv7dE3+cKFsPGoeGUZxK2yxvv4GP
sSF1s5zsSKcQ+oYJ2vPJwlaDAaQLOSpyqNoSQ+9VlG9mvNyObYm0dKPtaqBILJzD
ZcQtljeG6OeJF05UC611pquLI7y26c+QX77Cp/4PE6ocXXDiRw98bzLSn2VJzYfR
94a8oW6mVyzoRy9zzPnRNKwoxbgECDjZP1g0SEUBgA9ADVQ8OxD+CGf6MOZvwa9a
NyykSf3edYAVPk6Ko3QSumoAGKoMSN+jvxCqvJKjodFhMBL3X/WVhaxnkv3+MjUX
EZVwSu91GhJ2TF/TjQFxEhLNCg2FqsQres4/ahsKFiaMprZMa+UEfUU+sVxcW5B9
brCRmq/dEAL1ZmNEu9qdiPw5PdxLmQZprmjRguqbrKKsdiX0XYv8TRNSbvZU0/bj
sTKAbqN5N+B5wT8R1GHypBjsVn8e4r6CAm3PC9iC7YlapNezpWEJ5dMucV8Lkd7y
XyXc66lo/60Ry3bIAR8lZmiShFoYPaBLEYaGxI/rMLL3joAil3wnb+xrI++iXcwx
9gOWe4DDFcOaS/T7MlSjBi+MEXpQCxhkkftwg+tIpGOBFcExs87deYmjSEDKLdB0
z6Upd1OIojrGaSZ9EaVACcuYPAig/vt4fgWvhlOLbtkOudcn12QqsYP4nOOvWbjC
Z/wq8Iss6x9GwUKY/4FZCt10kvmp3kkbwdf8nNS5lw3xVhQmCwYWIZx32Ofx4G4S
oY1z3cyLVCXoBW+1zmTG8Sek98Iaf9eIKkRQlly0M5gArJUwJcwN4d2L5EB7olXS
y0Rx9IIQUFcFO65BNvF9URH9PKrGfEStzINKwONHwR0ZFjSgSTWYyHyhk2joGsTO
huEhxC5miMZpZ/svrgIOTx263anr20YG5Pgx/Fi3/5wI/uzYMkXHNIuaH4dI6+Fl
wc8rP5ASUzdVq64zVbj4s/ltmBj/Mvs0ip5GaeZw1PMNNHWCinKiQUSNjSE4wylZ
VbyYUcgf3zbfAQfef7n0/NEml37RgaF9cdmbvVmA7jSf+etWffknalrQasWeJItq
uwh5uPBdwDR+dIfxkWTMFLUY1OHRMpHiRWfHtM1mXVHZ5ectoR0eFAlA/xPZmzmF
CIN90O95LUHNULKT7ndu865TA4ceC8AUbeSI6XcUbwMfyUCcXcOy9lEPVjk9LVgq
AE6MmYcfIkm8rP4Jm1Gqbk9AUuM47BLt/9BqhjkPyZvzIIrnZ2pqcXEETIDPnYre
HKZOEruktIx6qOMzN/6rw2LFl/CYhSZVF7lnCKZuBnnAy1BnEeEKthnQ4US8CnuH
GXNwr0j8yr8vQGE0gH1SSHapvJcHTHJCGZe+FPueWNxUNPumiyaJibzTsv2yMSCl
xSsNwQNJgn96tJTIjNNqBPTmP8QYPxJsJBQD1tx2T82E2iBXvFWcAEK5Er54Qq20
WxYA2vmgxuRcRJ9uYVXDfSMYJ1Y+PJiXSBqqtDFvkFMdcAWAzNCUyuk8DkzbPwoR
F+tZKR6ydl6AoyaXReqV1trSAi6WOf4EWYkFkaW2RvgEqUc0/9qGg0Galf3HxZh8
2N5gNVUZ4C1vV7251uASWV62miR1QS3TGicpo/5amZ7X6ee/nT0niA4J2EGu46bL
4iv3pC/3oauPdzpdn97b0xicdUnefVBzPyYwGOJkKDMQDIlmejBvG05L8OYJ3T6b
/Gu3WQLadn9ydVPoR83el0yjM9kv4pv76qH4T0BS5lbflYTEEiLPMvuHoC5MH0Zw
SvJMlK377hBkZ0i1redkbPNEci7CrhpzfyjeRL/7/vxSz6p5dOu4dVzDQb2PRJw7
9Bnr9V4oOGT9MhBSOuN2ldg2KbEvhuoEzBJ8xkciiWNuMbwkzqVaz5ga8sVBDXYe
9WJC6PRS394jeq8VoOFXD2mOrDSPJAWNrzbvwblbLnoTu8QrZgZ8iWmIbboyihSm
Cv1efts+qXv4IUsXzW+zepMe0TC0mU/GCbimntxldO3SRuilt9B7VFMwp/HqQemc
eWnG5ix7BDiwapn1Cuykyi10Rlgdg/Hbk2dnLUHCieBAjqjpiQE0T97JfFqG4DCS
o/q8AG+9/uE7mFha4+H8vBBiFdotFEC8EQYLdZGcK3rmV9dm7H13v2TtkcshJrQB
ZucvhEjKVOt3Ls/otuXrMzwUMJRbdRSpMBR+PIvkS9G5vso2UmH5CZQfuy9swYXS
rTByBfkRCDGy5c3Q0I3Mj3UvxLX6LL3Lk41nzyC6HzQQXvad9M53uhKcRZFuOBVo
+GCV7LZ/a+43CWIPCVAgLT2XIm0hRpiHZ1VPf5ZHRyxl79IbhVlzQdvRp39798Ep
50D3mopSqRyKm/ZbxNK3uZ6Pc4xVAkWvBbE3wEdHfF0y/WMVsKkJ3clpmvLS2m6b
rj1JKVx5nuY6jLhsaJkQZkExYF7q/fvx8ghhPiCVUSGP0fzsubwwWLWicql6rVVi
Tp6IFCDFxspq8j8LuuRu6Yf5eRZmqQajvi/BrRQFnepVVSu+GOPJUS3fR8Tzf/X+
2kwGvHLAFR0MQuKVfx1XAaWlMN8zXecrXJft7FE0Bx6w1vITz65mXnBzsfKB/hTq
zi6k2JnRKlVQu3hzQ4LgXcE8gaip9cVrYd3XQDuAS1hLAtDHUwgQoSmb56GhPOjx
gxAl8d6bEaO1oSqC1mnQjGSfqO4u/DDuScDqu9q/Fz6N99mRGBgmOULizdvEn/Xd
ioyIGXky39iVOpkwHcvW/YsY2hJZWCw3M4lsLxufxMWi5ajv96h9wKpaff1s0h49
gT9Axj/cXz1w3zVVsfCNu6ohFMliZxl/8aCZs1qmBQv27GxR0o4XlGH3CFqF05EA
5NKU/AEwgqN0p7USPtzqga5IqC4U9l7CLr/5W3kQ8Rn8fkVYHtOaSvSoVIpQOgMQ
nIwbZSHbdqHv7aMFCvGiiDtf2d3gZGnRjKmCTaTbNygb8vsJUbBqRInGqc/7vbXp
ICuOT4VWGwrn+Znmxnt22SIJM7t7D0r3m2E4Okava8OUHbDCMvAWwytFzs860eRH
Wi+J9QysYN96b3oUMM59GX/Zn/BHJOTSqtY5GuX7ReOIrcd1xggLgcl/L8t8l+o5
g3xAwlG8Zp2U4IaqjRWot4erlazzB4pqhPNBBR28kBN/xP1XmyP9VTzCqlkcusKJ
enVSG/ij8YqjIw6Qz8TTVjiQgkPj4UTQodIOCamBmEBWTzoseZivG+fAWOkVHhEI
s9HM1U2qCGZvchRBSKzDQ6eUvpQMgvXytyqspiGRtiRFVlXkLvKOY0E9CF265OTr
8ngHZQo6aLDTuQsobIWjngIV4lFbDgQY68AaRfpZX/xvZyAa+7XMpsqDKhfubtRI
lSJbWlwAiocKLugFvKD10WDIDMmA876R4Pq3jrHOfzj2M0y8kOr0DM82djzQym9T
RvqLxo7RWfHxinZpY6IaF6WQTgeSlUZQSQTWRzOMit7PQqOvzpaTr2AVEbCFG960
PQpLPt7o6BGu/fKACIF50Xt/ZWA7EY1EP887rVfrouuFozwUjQKzDNqbA+M8jMKt
s7vEpud1qV+nf8b/jBFz06U2D+2GgrgGSz/IvggWZQCikx7T7PSWsVus52hEiArY
+X0snEat22Q5Jnwh6OFtVLFlwQ5WznPq54rOTvk4KHJjLSQDGCR0aezDrhK+vtZp
963BkarJdBrTFPTQy2OpryR0CrezwLqT2qMgyt/go15rAfIH/ssBWlLIHxobbwQv
XBqtucq64WN43e4Puc6V4ZkqvPdH2+XoFzwjCYYvkDuG0L/i45X2lzSxr34Oq4B2
RDS7mOZjA6VXh4fn4Kxk7q3LnTRZIZ+iBib4b00acZa/P7skb08y+d0NH8tekK7I
ydACuGtVT28+aor5o4bs8TZaobLcxVhtaEbnvjO4MVgKacs/AUvL2cxEJ3VH0+eK
cn5rN+eRHWXWox54dZYbvV4PWtnsmAJljm5EATRM4h1Vqi09Yq8w3HOPTkMohzGT
3K5+ptEPkUVulUxAZX3zqC+ZuEamefOF9OH+/ADjEe761N5YgsIORJE+un2dvby7
XEffxkdJ9vwL86GJXM2Cl9ej1Mii3g5G+XBNQl73tvtuuHw+/3nmJGqHeEfPOVL4
B2k18XMOTFjvPp+g54JjmMGsVjHs5JmkCZqYO3LmCtarCrPZQ9ZSIYPiyQVYJJ54
34uVFHkP+p1CcLuSWDVi0GrYNtzHVEfbg5fAMG2cM3pmhPjWmXfoarWr2VkVidU8
T6nHSke21hQHk8TxZ/fTKCaKLiELfZM+e7T+m7Ptb/sxo5JLH18EmFwGTJUKxkD6
ZIPyV+mqxBSxj9CRhDUj9h7/JpWwEhgwtPwovGDcm07cEMjo3Ebsh1DBP5Hks1ea
7VPkmsfA0raGbncT10dhq4R7heBbYkuP0ym5aab637Do8hJ7j3oCj2Gtv6sVhfjo
6fOxqGlW8z263ZHsiq8maIPwhqhkFu7V2sNPl5oPWgLpqdjdZ2Vj60YELNzF0cmu
rgTwxp+efQww8aQMumjlZbV59HVDEfxoHDnh9Im00WuyEDymzNcnv+Je72FXTYna
xTVHm0ZLLM9eVzqmPIDEIcPHcnEu6LW86wnRl1vE7PN0QDcMX5QtzEyO6qPkXSIg
Ne1U9m58Cm3rKeqsGc97cIPqonEUVepUvF0qIhczFh5BMFCJK5TbAbaBM4tIHKrJ
VxkRSAJ9y3u1V2QtZEXmygb5Ulq3HuYcfGuswLpIaO0D+CoxVNxz9DjRfDTwLBqY
Tc88/B+xeIPpvG+OJk8/2HCpsPqZIM5RqjiuAcgaaf30DUGgomTy1SNx36ixvJhJ
kFW0WO0OUoerWd/eFbcw4UaQgF1aUY35wulDxKTR7ri1NFkROKiVT82IElHy+qZk
o9p5QYG+BnYMU/b/4S5GRdNL5QJniAJK34XLcCpAH/N1P1GQhXaVcF5y3Jd5fhQN
NjCI+xjy/X3fTKFAR23j7NZdtz69MY2TDEKFBFfNvwha7HvuDYAMmsaKGJJrCnaL
SE8As6vUGQgOTRvL/1VTeF0uAXxyImPU5PKrHpkx0pj8M8XnHT1hNsUqd3hilgPM
IQ8uSGhfyQpR3MvQgYgSjpEnp3yAJe16RHdKiUJ51rC20JmsTAgmmvuxVn5ykhfg
2EUzxHtuunnB/LLqVFIqYEkcsU9EKX/RJe5xWfkZeV0j+U4n1YyKIbswry318D1O
9xHrdNBMlNnObvlDD74AYLOYNuCkazoKBIDOiSNyP3o7Nx+cg365kWm+MiZcA6xU
iIcUx7PK7NTNPO+jP7kYufP2+tyGJsTqiMNdFqHprkMenOBAN8Zkp6hafOTl1yB1
1JZ8PaRAqve6dvFYfCDOtYfaaEk7OM0dOSsy0d3iM7d/TcxhPyLjyi113k8yObSN
HrGiaPgidtnG6xgC5aUAji7+IfyQK0BVPcH6mWdmvdUjpM4Uk8a5onNo6yv3Gumq
krwLo8mjb+WwXQZVKGvR7JoflIcT6IFMjd1vmo94GptHcqI7291SmXEwrz8glYVD
RCvm9UJpHhWqh41LJ014FMw4ssRRj0N9VZrDs7rh3dIGJZB3hn72Gi1cHMMQE7hB
4P8AZwOrSvEJZySBHHzm6jw2BUOMLiPkb9wSp5O1IswF8+CLus035w+u33p4l6UP
EGFx34LPaHkSz25jD2rP2xJxyG6100p0Ss4+6KYW1ZaSiSraOqb2DNMTfhXfszay
dKJgHDSBuXKSy9dhhJvcaxp65X/O7sugq5PvvWc4aPNdLLAFSf8F8uga+ztQwjeO
PaK4bUcX6O9A3DGmgW6KPLTl2SDIICYylw0GEE4CB74EBLpT5RPKazHPHGyshm+Q
0FAPbJHIpdwGsm+7U2CB1zOJrDob6YEcnVEKBscinzvIEGVZJBY1WDVS+bgVJEyR
J3FYVvtiJjIEMKo5Oe0YV3HN5f/6moRTFe1JASs0X/3ILPTVkS5gIgtgCdrFqkjJ
IDVob2PEI+U+Iec8dGwxVDZOSZiN/Nt92Tr923GSIkQPKswIgDvv+mlMVhVbToaV
C+XWR8Md0hLxCXLBTpoVDxPxNnQpoMZSHADG30L7PFatQmZM/Iw1l4wCLt+qUGUY
YMkizFGgksyqPddw7t/zy6W+S3A7YKlwUtYqEeoMAroT4htBXeGM6OVk5mhbxQYP
oFwcr+xk5o6jYLlBBxzGQcnF/QxxyS+YIoQ54kDU1dCsoFBytzoXGvtLQ7TSXL82
CNIB5KcqVu2G85rMmk0QRnm3p/CxF2OJ4eQAqq4Mq74JSFQg9mwioP8xZJyT+TWU
/KbAoB1R1oQq/addkgcPetp7wxlgUtPx0LUElNSIh3iopT/LzEqKc7Kct/13Kay7
vTP174ciRdreuynjZFVlc5llQeD/mkHnWxxpzuQPo4KfWIG8Ol1+GZ+xpklG4zaa
uVSlNF1kOVvrmfjANpHqkiX7ERnN/FtOzEWHw3CyAzkD10puevr0WhIiKdP8tQY8
bMB9Y7Ck8GHgawCb/KDpQVOIt++/aElmgOPykfyX98BsEHfCppw6ykFl02Us6aba
/GLIhh4qwm42dZQsdTCiw5DXof4zfPBe6rDtkuHoRBk8brWzpmLFbDMXoXTJsC59
8bVTVcD14JuPqfoXY6TwTUaasmDYJ/VlaSzJRWBfANGtwePPzkIY2Ai78vU/sRPk
gjn3y0ixH4b5IQeqiQ9xASJxlpHcfUT++qYEMO9swCHMvP6OaAhJ4CAdxluoH928
+F0CH7+g6GEFAobPvYops++dOBnHOuYvs8NS3wMjxanvgMK/wVWmgyX7+cmcK+FA
GgALEG0jBZaHlBn+A1YaS097O2nQTp5QJ4SlPc7R7TsIqYlLmhdQHnDzcCpxYXWj
m3ikKrUEresxVmJaduGkjIppHYXnfl8gQCGLRPsaLtNALXorTlfPpI9UWGgy+Z+d
BvIlRJh4rahO13KFHOvfeqZZc6aecViGqqdXKhL1KoDCh/oxqmfXMwxeDNRaiNII
mIzObg6hcupNUBIMjkIhc5Io7EhSxvZzoa9VArFAWHtcRhgIKyZGcoc+7KticDcH
utEyMO+EGz+gjgBFuob07AAr8ikkPaZxhsBb057bWUrmEPLlbRnj53t5d5XrgWYV
1BhETrj4Y+83XSVoldL29//FfxPTCNiZdKcxaRoEoxVlk8q6aHolGSk6KU8VPlJy
K5CMGx5u7PMsc6X18zsih3xZbs7GFC5rNzjMQ6K7rHuwvT14ZyDu4e1+eLplCG/3
CnGsoCy35gIitgvk4fwfChGuDN1F8j7AhHD4G5RozayNlWrynPd87+nnIC/GTvnf
JZgFw6jOp65Oo496QZm/eC/LQhLb0FeyACD5Kor0r7OLwoO6iosCe2CCpdHN9H4t
k70DGXQdhSgGvRlA42/PrwEIKJIPYrPC2kzR8yEZ/Lt1VuYG62qvMBgo1SVVMiW2
Q2ERjvF3h23/biDNjHaQAt3CnfbO5DTNJ33XIVbLKLiiXQ4Xpt5VmGea35gbCKWq
haPyVT6lwFndWqJHidMe29WKmLzDKLxLbo9KJo2nRXE1adauMthU0zUT/TID7rqS
+v88kz1RhYU9GpT4vQdafnIwsIGFBJky4JjuvbEcqDrgOofu/0zxvLDlX9NL5nrk
LrQnpx48eedFrE7Rv5Jr174csze+ejK3xOyfdN9yHfln4Jpe86dU1VXBkcYS4lJZ
Injk5NsruUxnUPa6iXWxgn7B9uFg+EpYQRhj+aZWFMPEDj30Z3jbJrYlBdx5l8XY
Zd5EaH58o8HJxpy4G4icEgzXOWHDczI48S6wT93eCDplzjJkVkHiEzIDGwsLux6K
dTs1raZvSTj+UhFBwZXCih0dtBDQwkevqIpbgSnVJcouGQ/QGVWfiJiQ2jFZmG8g
50UPquoo7GjeCmrRKuw1hk1nxl2Qx5/L7CL3k3iSQ0Lm0Sd/GXP5nszhATJrYjAO
X3D3CW6pz9ZzJLQQts6o9X0D/KPF/iXKzi+eocWY0//qIJeun1WVF9Pa/pwpDZDK
bKbch4ASkzCSEE8d5xY8i4+o1jYq2khtdrZLftj7LsVDKOHh0AI/aMYyI0Bwx9Pl
/vshN/r4BW+X+9Tvrb4hAlTXV4YPTgNLiwndxVagPuX/Xhg70k6IasvMEVPmWmom
9la/9I7ge4HRCZ01jpPpM7INKpGQUaQtj4ophEoRA1TkCaKrNTqf5e3ZWYI9NhR5
Q5hE9JG1DveAiFTOh7XJu0Imh3QIxJsCKQTXQ+JYJwOeityBhinqSkyutqR4c5Kw
Hgg+mrnSEC9wdr+ZTg2/sSIVkx0mX9f3U1CFAYj9tYbSwwViNV6JwzWvgHFttkW9
Rkt0oqhCU9itQEzzla3OZAv025WlvqRBlkWIq0U6bf+YIBPIwp1M8pqL8rsWJ16W
ai/R+HQSmhIcotSX3z4X/9G7FmVE2bQlq+0KPgTQSsuHOG6W5HKiXmlOmgY+jT/f
NlIZRNCzCIGPJoRJpbZV/CCqPNpbN6saOBUhOzP2eTnmXhV/dCbkBwsH5bR6QBTB
s9/1T9T7RvB8WtIKz7HYIgTkcCBAb7u0H6S3PrD1STgbFfgUjMX75tFVqZzhIbst
zmQLKGgWqaB+MhVxfBt60nD8EpSGF0uVRcnE6A85BDIs5ljy7vSgJPyLjSfOUaN4
GVt3r1NsZYBiu0grzVd5f2cNvsA6e0GbkqaPF6LrXwBo67+p/ynMQxLX5laABNKw
TVRLRs80uAOU30zNuPdB1As2fLpk61SwdqrKZv2kSrBKKU7hYyUJnjPxc77JjGuK
3fx+cLqU3KB8eUdUkQ074n6M0syA+zj21zyCTdELib/Ro7xxaEe6A0dJGuK6AIg+
vmDDkKtX9UHxUlXrSycQeuC3c4mOrtkeC3rKhTlrWAA0CMXHlsxs4EbcLkBs8xU3
g3rrm2D6Y76WCN5PKkLiOrIfkq04gL3XkApN1wjSUaRqH2WRcbJe7avjl7jPdns7
RsUpYnA6n+k+/efHMosguUf4kA+k/D9rmBHfomuyMIrLeTFaoy6laUH0ndS4/c39
EVAmRONtxvuCbswV0lL23sUXdxWGkldi31NN5dZj6CZF+BVbra7O7389mEgbbQZR
d9gDid6ABKfGNH8vCpINS41GnH9uISITecvn7Q4+2tvPCf1N8XSL1eijjMir78B8
CyscbgIfOSCcaA2x3ByriHvegsniZP/FEQsrJOiy8PC6NDIunySemOjAiubv2U8o
HSs8K2aZGmUPVMSCmfQYTncfo30S88rMbKbwigJ6G0z6KuhWst/C8XdWlAe+e/WY
8nwQm94QMvaOe9v29tGJbYtNcXPv4zq8kl5qGkXGCsNcV7H3f3UaqEvKJwIuKZhf
eLRkAg3GVad03spidEv0h2x/1tLu3TUkaDok0nkdSzH8v8fByFXTDys5zPI+lkog
bl/occKhcfp3MIwd6KVrxFd99KCpGc4ipk4qnad9/pYYvf/tD+2Px7AfSb6Kf2OO
jWOsiTDpXB3e/8fPL2iQIaHzRX4D5RVR+0sdmlYRZ/sDGTvzr46jqgyaATLFHcZq
uCpTceUOFYoSg28rFqjGPXwnKc53HbPqO6KWwTHRz0fDQS6qPlXBlJC5nZRYzUd4
c7iSAmGx83RF/71nzpv8ZrCpGnnPQeZO+/dcckk7FnjhD8QnSh2M1vqGKMhwzzc2
vkrx+20fXKKSkoo3EIHMYIPVyWfFsNL2dJ15hs9l5iAyWdCYx4fzyrxcfcNdxUaQ
30bjpioWYFWGB63B++ewtb/PvvqS2AXKcaMiazJZR2PzrU2FdetxbSKKdTFBBpL5
AA66Svby8KAiO/0QCmmQeOjNBoxP2fEjkQPI3zy7S97/SlKdPBsv7W3ah/IR78Yl
MXsiTwjLjthAgtyESuADIUFuA7e1/ziRclUxOxTA5RJARYBjUbZidjU+1YkQJE8t
abdyxJlwY8QgG5/KT1LSp9NVOpYvLUEECbTfWBAmObkaXD2mzYSfQ/JBK/ooLz1l
NvXWYb49filENzBNIMwWTJXUg85bhf2Ee0t4/wE6GMggTAb8jIVoVhUl6JZKGWp5
XPHMjBFbaXG/+FWZkA6oLno0u0ar09iPT2hIImnY0idra4HQUKe8l/fB8fXWkgmO
i/MmfZhGacMRL59QljK5W0rioETk915saDSkhXEJa1T1F/qRfVE48yNtc9HtNYQd
8n9OJJ3EFlbLr8hoDIpQz4BA0cJbTCGmgFiuDFxQ7bGRxPiNPrR/ksXA/3h5H2up
iLKoq5sd7OtqkWUkFsTkYrdLB4LuCvMhzeqxsw6TRu2m/AwNjSRPFnXDQZJKCVue
habfo+eooj6j19PZuqFS3DRuRDT4QDsbSwCgIt2srOvrtweH+B5CXMrqukMtKYet
SJilCKSqe9NXN24R+6e5LTVv1puaotGXHtL9bHUwGwS6pYZtkDZlukN/54aLHB8u
kYwIjYw++Rxzh2ZzRdiMhbUyoi6Idiiyfyz0M57uPmKmB1ffb6jiDJ9pwKCO9S0n
Cip/yrLLNtBdkyuzX9SaTIWQqihgBvsQGTvKg2kLptrIgHFMkfW+O7bwRZHwGfmL
f0UJNk1f4/EmKpSSdk+onvoFSHmyZ4yn+7fQxdmfv6EBSt+mmIjnBpVw0EV9nMnj
7eTsVf1C9ryNm2xeeDBOt3y02OBWQlkwl2b1d/CM/NDEIaRtGOFRKgWnswb7KEuK
6j6jCy5kJYOcyzmaN71ADXo/TCk+SrZJBf/ysp1TdxGLDQFOyecFk5JjvK02S/yw
G3rm+JzNYM7xYvbb8iXtYfzBreEgP9Br6FEm+ji1cV0p7Hiz2Eviu+llkGkg9zbk
98BEWV/elWiZAphw1KhNkS5/n2BbuazMLxAtJDRj/OYGsC/eQzOi9xt42hu2quAJ
pa7zvKq0XrIDpg091l4mvpBbFORfwTEf9j53RR2GiIIDCAO59Vli4y//CZz9K5WW
3ejdgB7R+mlGptpRbFAsqEcwy973SMjP5Ua6WcJLiT2+KTrnJ24a04CnsYjqGjLt
Ibqku1xW6hwTQcFvYfNxDpu3umCraUN0FCh2f9WnzqaMkOssT3hapi5npxkr/a6+
mXQcMjNYxdRBAdJU1fjQvzztj0vbgHZ09A086sQKHp2VIIp0QPLaVpWu1AkiijV8
O5LR/jZCiGqa062p4L2OUaTUz/fWrRkQZH2mpyrBT4rC/HIe9PMs8vYSy5gcjIfy
tpk6m1SSUJfNj5sBGu6LRdCbWQKWAePI2RDxmzLm+JKWWJJy04AnFdM/TeGkxjF3
vjX8eIfB4b+A09RgZAsX8zB1QNu195giMJIKRbhJQFqUSTnRqzSp6v0Iy2b3Lrlc
/xmLOGu9npCLrn7Nw0ZXZJWFKrJxEV2u5tGcWLpB+IKh9+h2zWgANrwmoOq2fCEE
rB+j9QWyctdizvPmAsjGh618P6E3Lv2yxYFv/HwPE3BCnqM89YTEoHMMAI2h3gcJ
K+rsBUTk0hd0Ww7XFtPYNLRMHFHA2/QKFjouX4UJIckVfQ1hOQtXZqg2baJjOaAI
ilvIU6OlC/F+eip/urw9+oylzPJahRpSfsVWnj+fhOjtH4E5f07h8NhGeb/l/HqA
7DpzbsipkBS0w4o6AmEXzxWgiXbnZZOLQ1f34/V0WrZzYBSH7g3m8aCqsGDWRbid
u9M5rHGsZ2GaWDhbb3UGhr6gkVVo2lVEmRItlf9coPiDuOk6CHHV3Lswjmk+ERHK
L9sB0Gw/nU0xwZ6d5N8a2tboJqVQjktdlXho3KQPXPRGIxuCCc8ZXWXLWYBJGSFI
1qh2GJA5vxHwfmN5Nsuoqv1OlkmM1QZRK//QWkfr6lviwZdVIhSveIeQbl5vreyC
GoqXu0wadnxXCZHXBbvNfQwzqCbi6X1ack1hvbEy6ICKgpPeNNb/bdT2scVi0NQG
rQ+698DwlVKZnKyvtbxmjLYTQsEDNAh2Xmm8ZI8RYhZaYeeN7mmbZHoTpMasA3sT
p8evJp3px8jd/CyM2+R362JTaAostD7zR2aVoYm/PQ5pQFS6sbjW7BaSfzRBl/p7
admi4uNHNmcfl18nSaWAYuYibbn4APFsILE+lfVpkuNx1vzfuylQJzYvV2rV481D
jL6YrlCbC6/pTssufrZefJ9xFAGeKifxcxAjzhanSzq7/ZVmBJBHmG8+GiKOEH1Y
AWGcnH005/JqopKjoT+2lG1s095wNV0Ef+wBTf+BC1wgvmoFbAPGqFGIgfNg6XaU
78ynppoeRTWCpgZv+A5zoQv4iJEgF02MebJgXkNrtRqRSYbVayvZn6Q536mko2ja
B0FJLCoMoNmfmwX7jLf2uxu5gn2cQwa9Ekn0Ry5zB9w2XTJXT7YKNAZbdmYqx1Mi
Ah9KMTnOW8IYt/WINuqqFUG97I4QBCgjNLYwkps0NlLdfkw3kTwOQHJEpi4ktbV0
/o8ZJQZci8sJqXlinnF4Af/G5YB878aXY+ZP0GgvA/SmVI16tJXDhVDtAafWclvL
8oU6DC9rdkjf0PG/T0AiWzduljsOqczvWwbyMsaS7kzL8pzCeVZw2TrjMc7GykvP
92psNsph9s6kCjVmGYfE/fgjzd3Jqu5AvSb7ekrVX9drY9FHQzkZfFZE02EVQ4Id
hnIDjht6LNomRXJufKzObQRffitxP/LFE20nU7SEf4XEPB6fB48zmJ/xgctS3xbF
aNnnG9VVqkrtGUDbpOI1pDUSGLm7zEod4v8YJbno7qlMFW72lL9p0WAjlo2npp0U
jsVfD4ImQ4X7QZZVeGQ4txKza8w0hg4bvGzZ6JKeN65RaKKKwBHVh0yqRNVxiWtP
FjIDHQvrxRO976CJSS/q4Qj8hYfkKQ83ELKW/zrAeyDzkZS1mK3vqJF9ylq9cS+i
lLYVqPsVVb8K7Q6z57inC+yprm9TPVN/jaZc6ErY2vmI/s9yJPj/jU3N1kBmU+JZ
WD5nqeRZbuH89UkxIHlzK/5NBhbUa9HJz5z03gaVJUgBzc6XL7wA31xhacWYQFUK
u/1cJa737BeGDU6DMxmT4Rd5fR/udQtAiHj5NYqZSgzp0cbpDot0f8KY89QS3deh
qfX9xRTSI+ohfTucKQanfukjYEiFpG1I3nmuTp8a0SAhVX85hJ0uVEq9C/ZwGMdK
iBzQlSfQJqL3wBZNZVjMeIJj+AgAoZgPZWyw/5c/dA6t7bcevWSjExqkEsbOqWnE
o9rQJpGY+totRwvHPcE8n2QiwM4/RN8u+8EtUS0Jhhvg8tfAABT4BZ1FZRDBAt4c
kWy93NGSQZpQ7Wd7gFsYPwdoRzNciINiM+x1IerYvLZwfu5TNpw5fcCfeziFehBq
9H5eJTu/wRo6MvO0C1OZ60Odny3+xrwnwbfUkTgYtw1O6ulUmdCUFZ5EPdfwRJX5
32VjAqjL41XvpzmnLZIThBHBtk6iBzi59vQ/3iP4GVs7ZOB0q8ahNU7C7f/C7haD
TWMh5A30F0aqLdlGKZBqa3aNCMpTyChZ4TyKHBMh9PNX8sEg2wlmDsOWc/AfIFLD
wbpBix7ZttGcthxP+HEvjLKdsbBrrtUa0IA2tDvT/VDvgOhkY8xuOgiCKw6jBT3c
tufLY4QI/djFIxUmCLwAVyZoHEHLa96p6OOcH7xRbIXrYF7mcWEV91JcMmGlaCzc
ZFAmr6nKLBqqt77xL0Ef0CfFQC3UhMy/J57N4vohWjH1dVWGNa5yn/ZUaG/ATjjb
bDsZ8BgaKUO7PlcNyjCBTDfzZhcM4zKCGhkcmD3NCGfV2ob8jl8dcLYwbw1qSTld
eFKEAKCbB4Vrv9WQVhM9I59tMeU7SExPLvHmttkYUQpgBmlLW/pTmQI5HKJmgeXU
M0GdXH+fLg9nFESmwk2XXQQ+1FjQiDVf+wbbmfuNvkaGJetLjO8kE0vTdKzi4hD3
hW6EJjA7h3pmj0UGwky748rX5ofRylus4IS+BBSWNEiW2CQqel+8Nx9R41OrbUdU
EJn2+VoPlg9jWhPsw0/PIAhm7WI0r/YszUxc9Tqmxb/ROHTTk7RF2xqLynNQpU9p
S9Oc4hR3s4EDirC696V9+uySSCboQ5d8x0u++Kt9aj8RVR3cmo2H39I80pTFXLUr
J+b5OdmVfivLMpMfb8Wobcfa4nxJq8MXbGPhh17ZBUoiy55ls03RIQa92SCDEbPE
yfGIhh46y6gPi4FAvrjLCaVr3bXeLoyKUIUPj2UYZ7fTRuBtR5Sh42DK0P4rzQU9
p/vzX+f0ARcuecJrxanbeXf/rJUg/s4Az3juetXVbUyPKHqfiH2quOqg8rmIBjoG
gVjiyOm+elkaizVZIC0Hwpb9hz3bXsOjWOucKg07OmmLveIIRWq6nZs+idcpAUux
u+0EAO/9rtRIfclB5hqnkmh/a2AHoo10ZVOF8FyaqiwhzK5kk1TcAmxU/rkc7dRg
glHmSQOIkovVjAFaJlhB1GHqyHlmjDfW/Lzds8Zcx3YUPsCYcMsJ4p5clC9yzdp1
ZfKVaoMEYY3h8PTOfpcbJnrC8UIk1+2KPo0WQBmiNXo2cyiAmGMZb6XC0DbowVVF
EJ+o92x5bNB/q19fcQFWUKZJnc1jKMNQlb41VFpwmBph14SXkNNFwjF5Un10nA0E
BYIWrenUo13NUnSNOhOGcTRwdp6RrqPe/k3dGmeRiZQ9751uEJiEMzxyuejyECli
2q0ZTujxMg0uS0BNdoe9/wopVbm3n3oRvjVvhzSRLHNq+zfLnzWmRchh+l4g/3oY
tfYlXmrLs77PX/+ycZ3tM8wHC24ZzJjnbVeRAhqO1mtW0qiGldPRNaB+JdC44jSQ
B54rTcedsqSxSbQteTDsNtjYNiifFknjKb3gHxmPR8H6GZ4a5KYQ7iX2vNYoipND
1+NKQx++zgTF087QNcrniZqhwUq/+7qSS7N00fOK02l3oXjZIchx3H5P3xdeP27u
I5nR0U4DY30ryg24KthxM/Io/U8Lt9c9bjBeN8LUwQTWeEhOGchqLUo+UaEXcWaG
ud3j6Sf2CoKLmMtm0pb5EjqKzDuZBGbXDsvWWBav3r0pNGj0k9yhE9jcEEFq/rXd
z3wCKqGnvNDeyIpJMvowu2Tx5zGzoANdwTE+GS3Ry64hWzZi5gMCz7AdVLlGPi1h
KJlJM6cftXYFh9FS1jxgzuvPTygjBzbGzT2/0AXSAwcvKPFhUYcr/s6eptrYyFEj
XrKHjJ+4R3YAOlr27OGCnPHxJd6vj7J/MMvCS++uy10o859GiA9ob14p0OJ6kR2j
FF2mAVaFu+t8V3N4YR+3Mn2AS2qmatzjLukw4q7TVFoP85IRtpjzy99U6RxSAkAo
rT8+EhSEc9iXACK+vali3bJXh3Y5epVGxMtO0yfe75t9daNnYf5/gr/qsJat/E/w
Q2DsTZFMvEh3P3syGDxD+xg0ostYuGr71jzMxZl1eetFZY3KgUbrpZCgWxG/8XNb
zA54oPaXREze7pzV9jAvVYHNigJkAcPQ7tNDM9NItM6ThuJit0GPZpEW+NzR3W/K
VdOCNXGTdsEtVL7Wdx7vBwMxceuStMql3p46oPA/ST4XKSoCTRm55MiCbJ9JHoCj
x3UEKEw83ffa569A3FmRd9Yxpb920L4gxVvyzaze5uw07YEjczUxXE+zd0YMfLZ+
cfrPX6nuzBKapRluiKzq2VisTn8tRcut3IhWqM9tL5kzXBAT3yoNF+cZ3h6nihRd
XL088r2PNFDwePziROcapAh2fr48RCIt3QsxC3elUhcTlUEZi7ggnPqyvnGe0R02
05rdWHvng8ISRzu7rlmR5/IJooqeeznLuBEqNV+jUV8CjzT4/5GfZ9xjBS1A24II
3oZzWAZcZHKVEWKu7zAU8pc/TfECpVTyqL83gWzuKHKio6S0KDlBgIoUVpfODWJZ
1X5ln1qPJ6vThAtTznCRgdLi8agh1p57VNJXOBJzp4TtOey8NZHiXEqQ93uk0AlZ
iHWNAyLG6Erw5h2vWTPcZGCKHSzIKaNSAtAzyxMndKwVt+VzAyUkRIrk8I2chEt8
RaIDsWTkm4fn5cXHkUGKdp+SiDbQ7g8nIBbCnHmWKVLNEdyon85K+VGRnPnhOBvw
CXyYVDcnz8utJuBVibF8GlBOrNQnW9UxhS04PhQxjZJdXv+g4Xh5Gt1HfRpX3Tno
ZORK+1uXWkPJMyE/oU/WVp7GzB4oNP9OfscEFXCwKWIwilEPbuqTIBcrdZWisl2M
HjgScjaV/pVxOiyszKaVUhGmufTu6KXYRpR0SblcW2riw0inaDoHTQqAL50m9DsT
OI6Uc5GsBtbG1VBwoKI4YJU0QAO0O5JWw62TfvuYAV//4fPnOH7XT/AbI6pIlnKr
ddi5ymOeZrIM7QviXuF+qlyazjQr71kAw7aM6Uz9bBdW3kkBNuGx8Zy4fLgANsCv
VCmmCEEdxRq0tsiZxtJIGEvks/xA+SnPLcDOG4cgihSkeQLN4YaK/8ZKhigyrWV+
4VFjIWNQ4FEfnywUHNUc+Ur8pM0L0pvgcIaMlojp0y2Oas2d9NQhVjT1SLd0JaFR
F1xzEB81HzCoiRHrsxqcuAS6erI5PZfRO70SoNHiMaJiMKzhIP3GM8og9IKY6oXj
c7m7IvBcnKGExJ1Qf0cS91qbScMfjveoSLeJTudKMJgEkJl7YmOvrwMJtMTKlJsz
4jCnt2pyqatKdBgrWoNX5zvnkSLr3HsAZV4oYg7YyjUAQ81HH2X/MeeGdo9L9FvE
lwbhrdnH3elnZ77YRUXUwRZY9xXmZyt1tVDvbCM/Km4W4a1W+1y3RTu4F43CNZTH
Cr8ieXIzsRDdeBvhBdpOozyyQnfK2G6Zum8Fw/YbCMEPIikSPf7e5+4g6L9tJWg6
/zi7pKmudp9tCWAiNDLJFoP29QZJEyHr8Vx2+M40y/lukgOc+bXpeQrlNZci7TN6
zgZqCjnc41expRSTYg6TdJG+xYn1E9YfzjiDjIyrP9fBC2qhP0Y6jM6NLhuFjHEC
sAP43kTR52lJwAVLHHUuf6scjkwLjllalCV5KOZifQSsORdF0AkVVUMlYmbAYAtU
GOiy51hEAvkF4gbSWW8KB6PL4of4rCVTeRVivXlDFddcUY8++xgqa+bmc1CBwHp6
y5iLewOp8K51Vstktqk6OmvjO3VvqRiuw9mYPLHD1MlEZf7Wq2GtwO1k3djh7Nq+
Rnbx1SrXyLgC60cBIYCBinqvuZL0zRXHJRQyCpEWJa5sVRZ6955QaeVF2CTyA7lX
tGXttMZpvbpnoqiymyDtDmOAuQcS6CqcXTWdfzaWtT5ixChqGmmodAVdUqLMmhIl
QXHzox/73iZVW2r3QznH9c4RL0FH1XtTd7iDfGa5I+fj00JfKWFxzSr4TrSB/ipv
Ld9X7QUHQYMktyrgOmhsoTJYPaM3a6SeKYAawFWhMWkmQdg/ln2D6fX3AM7XRZPV
jTzjjNEekyxdVOzNprM5BSZp5n2U7a+C8Lix/JAAAZHmO4FbcSTbh/izL7094twa
v6GZFOONIdtSwO6fygF88SOsEXv03y9iAW4ZWvSeenSUScr2HI3EUkrKN8GnneZ1
QkYyaHbiu4JpXz8CGl+LpypIO5sDVmb9xv+z9WMybDGfeae7dsncBFJ2D3tdhuD+
WhwpLwKjKRUBFwtuUFZQ13HCvnbxuks4kJOfm6+a2Vf7L3kZWXQqQ2aMkglMy56C
N0WEfIRnJ5GJNq+Znp303vV39ta9nBIgY0NzhY9RdIJftI8HXCf+pJX7CU0AOz8r
zzkE56u/K4JAJWYm2mf//qtAIJenyfXI31//8zVbNuh0G3c7iLCoC+FzPWZMi2mv
7EN0JBy6RNmGvdHonbWaeDXO7ZBwNYzM4o6cQPpIQ9lXiTTsHd+bvlPqW7ftyzbN
2kVGEDbzDTFbsay58laMPlAWRqFMxGbiLsGaDtFS+8LIBLvOZaTAnQ5fF85/FvwN
Chr/AAlrZVUbFFlYCDuuTj8RPj5aOFpW6U3+4pmkxIpf6Uv/9TDM3pA3NPnSVehL
JM2mYKSsDH2SRo4E0XSiEhpmoAQRpDFsgEEGv9VaEKeI5FOi7V1kAFUCBoQME14s
0SJQJe3grQHj+iMR1+rR0eKP6zt+tP3/iE57tbpfhF6dgDZCIFMuAR33KRjhNL8j
doxnCaGUxaGvfGxiNUGvXmBr+NCKsg3bh1Sk4xkK/pTJ7DTKdeWkd06zZIaFINQM
DP456qAb8/5va0UH8fEsytfi6zmdvrh4kiVfbu6QCSpSTE2D5xSJK88DsWge6mQg
QyMS5sx1cE/95DcPvOKHsDb0YaVrEFLofL4BWN9ISLQrMgUD1YGeyKUehbBsVOIA
TY1YFwZr3ex/R8UTgDXH0+ZdcIqJcLfbKyHnenDE+wKAGEFoXjr9FVknZ4hgfIAz
eT/QKkHIHipMA4RaFowHhtIhB7T9PkZ/+boJKRUGHyQhm6giOrguQH9lVOBnlc72
exZrinY8jq6aGXIVlm6W1V8uo7WTdEVLgHWQ4rzu/hqn0IWgHIiat0V3Buk9wOPB
WoB3rexQFk0gi1yHZOmlglz3rrkJSOfbDCLT/CA8/jkPqAfmE6hZyD4c1KyLFvFf
jii8uMvVwhYLqPVmFajhE6XdCNXj2WrKxveiJg5rRPjE352O80ZzkHwCg/9yO1wx
EmfwQno0pKKShlQGtGBtuOZVi+mvBqdGys0l7QSPHbQQlQpYznuwb9CONWZ6IMB/
aRi/dUpw/8OjwDfkroQAO7USp0l9hbXLtZ1+2UR8PmXx8k7K7YVAd1SjhSsuXPJ7
zc6w2lXnNpJgo7nZbW4iRLH5NUgSQTriQPFhbWi5VYp5WBupCTA+6fanVx2pF/Xs
GqnbofeFSVBSKBKDPh0iV2MVHaGFjFFMJky91Ap4SES4YC975hODPwZm5DZtVDQj
XY8npE4cMPaj8WE7QVCLanUSsRF+AJ7BR7O/kTvp1OQo+tOhDTWKiU4kvpgJGKel
+Ft/YM75GJtraM/59oj8Nf83YIypO7/+R2bTUICcBGyl3B3HA8j9XF1/YmV1tEYN
cKBGaA2pz7c9S6MEFFPHTIvOarfuxBN4SiBXp7XElJXVq3f0r2B0vwGNCR1I8v13
6U3NGUOGJMxH9fp57W6H63EQgRJIXgW0O+F2KJpSNdQYm7tftgKpY+oweqgW1b9L
sZnpfbUR2G5eAGMCptaV/YPGjl+JJbjejsXF+tERL9U4lXJQeLuqh7XfUr/s4DN4
EhxowJBxkAXYxxwqyptl+AkeoFEd6b9TTs+3hvEyDuIsxSCSEMaa4G0/s+TgonK3
9p/5CaHnakwp4wX4Hk3+tJ1XsrEniBrwklWd4l2I7oCYgSsLnjZcZYvFoFF4qNVf
eoqHnlO/jvbUpxqetR0TNx7Q/QznUPDWoGbO2EAT5+hK0pYVw6/FQ/07ntRoQLsw
P8GzmyC+7NnfDHDxGbm6ftSjVa8Qv8EL2mlDRji3q1EshOX1JGywn86Mkv3pcgns
fsPOrNv/KxYfuMaFTxSrVA06vw6bpR3XUNpNhb5AsOjSgIdRcqgsn1+jtKhP7f69
aMepo4OvLYdbh41uepvHMuhrJuixX6mdlh6Yyz9tA86QaMiElXDuID4wy+3RABko
/QDfR42iqb5ylG2IsOBLAz6WAbY0LHwAMf1PNrzZB5Ff76+nUaow+LG4dqA8erjF
8BdU40E7ZY5cEQClm2HsjPa6GZQKNfmvjxWQ/T/0ZO3GUPeKR7FeToiqJ9Cqj1rt
a+ONPBGWnWWaZhuwAU2i+rFahsQGwM4Zyc/rKpF5txtMthjTNJGJ+302WyRAfO7C
TfLCj7qfxiUtNlLE1n7XaLuOwV36eGoqm3Ae/+t4DAnn+3OQd6tw0OWcjhMCtodB
GNXuWyVBz0y0rVenajGw5yz5svCjl/qN/ZM7eZ5TWBQza5d8X8E3nxdc8d1g9XZo
qbTq92jNztshjt8Rp5Hkeu4qs+CZCO8fOHliJNMyN51WY+e2PCkV34CST2HG4oMN
AMXl5y1EURUNIFc07ZXlva7dgZS7gRJoIrmKo2YigsC9qbCx2y3NM021UyKvD6Wv
LSib3uiPL0mlz+06k0T2EeuQqHFA+AKbq2E204ep1iyaWlZDgpT4Ue7QKUwZqADw
N5Um9CjgE9jTiudbrJ63E0ydoKZOmNGisfxL5a9bB1CdGxCL7v1NzjIvGhFgaJt4
shETnR8SUJMmtAtKIAsShx/S7tfhHQb6nc6L9wMdgXpeHeG0kGSAxqGLoHYN1N0p
0A6VhviDuaozYVCaoPU67aHuEmB8KTICzdbiniOdjfcFuscFTVoQuGSwF+tw8pLM
vxeAVUJAutgyLAHdQ5mETCJo0DpA48Rlp4iCwm7bFn4t/K5FJxyZiVQJkcrvdlWm
N6UmhVZ58RKoPZxiWB5/ka8r1+qpc9DCuQm/kivCiLjnZSTeQijACwIVzY4vJAwv
5twROThijp6GN5i2pag+LIHkaA72qSp2kQYdY5k3dEaQQHPacTTdOdSHmuM/cgfY
UAmqy6urVDTsS82nI3PiqMJoOeM/XB0tgWKrjkfKQeTJ2YK1Q8wldAi1QhWjh/Ua
npok6EHAVwkiedloXz3US20MwGE9FKTZigxx4xNkpT77aGB/IfYhTkS7G99vF3a0
nSYvkzu83rUxiHh16UGCHAfKegX/MnbIQPrvC//Em0oF9pBhRONLcJ1jrtLqa2g6
24X0ZKX9+/FnfnmE5Yd2BAazfcVP/umTrAbV/3sJ4jzjkrwfkS9XX6iTEGLpWc81
H+Bjqte2NmonG36l/VuvaNZ/ansWcZ7JXDeaeD0SniYub3LzRC3uJLypf75/bXeO
yfhj3aD4B2P2KjE/KrWRYLk8Q+wtuxHm8PSCSjoWcodSJZ1nJec9ly39QVdhK7uw
8UHq44XhhP9lpBMt2f5AkJMPvChCa9SLacYgUIS276YftUVsIf0P+HTaln8NqHG2
wd8GkLfA6avos3K7L1c25NoQit8aEQiBaXCEQRDgKvAWPedVHpX7qfRIIR/JfVMX
NTiUYGCzPCdQlFg0ADa7rTeiDCt0moBP4HjyvmwcF7PH/hFPwj6Njuorm1bvdZ9o
9erDuw21zRRNFK6Q1dvQTnvnnq/Yk/GJwthmcQmz7W81d9Jdy9XS+wjsAzaZm8Br
HVUK3lWswSt4qgjctOkThRH5zr30aAbOqICUFlNVzaqYqYCX2M8M2W++wnQWauOs
SSm0oL1tHBLsHm/IhzMvcK0h5eTc4qhpArNA8PN7s3AmA6cBuKzJ0aB9n89vqDzl
LmwhZCd/4KShO5WX/68F2CmfCybZKym7KhT/LQeeZlG9G6nVfMEK5dXYmNLzR0fW
IJ0Ya9wIwMThFjk930//+XxSQxOgw9J100Vy0QnNF38OJTJ/s8lY/oEdvA6enwnT
cNyGJ72LNHCLNR6A6l9bsMXHFKrsj1AeRG9FIJzjA+2ypnqX5+j2y04h8TCCSXHI
RAPpES/y5DZdblVQACXJCR9Umw+pCpMYMB0jZV01xk+o9m54ovwZA9m5OnpHukWl
YGZWyuRQg2Tn9lnpcG61uYg6AGE+JicIDEi7GufoYx4bl0Sk0tDXwNh8I/D0FA3V
cZqRaAqiWRrheG8cw6deJnT0ig61WIGKE7HVrI6hTxszl3AIDx7don6JXaym8qtr
a/bfUt67QB0I+S3cz9YN7CzngJ3jDHT/gbPDWDiaiTTdclmS9EfoO2EPbKxYEsuQ
lvYVOOVWbeb8f0ya+HtfJ7qV03p2MqriEdjefWfJDqhNPLsclR9rWtG1JDqxagKy
ZrL4wZBB8vepgLPkUS3dX7zcuIAmiRc4kcNKzKcxR/Bcl7kj6dca0jf2+aeVR5gZ
y8qJWcEYnypajkgeJ2NMJnBPZlnVOOszzwacFWhdJnFsh1N8Pnqe6xF64XewR5uv
R38fEynY3WbMF+q8ZcN7/RNp93F8E1tJ7pmArEyjCSh74i6l62j2xAWnMl7/c+2Q
Zkr6IHsDGzs16pfGZblXz4PjJ2dScdG0wQ4uanWNFqylKBqpxghj1qwwOeY3i0Io
cskKxESpDgTOTRMSA7aALTmryjZd6Ny26wlQKOVCos8oUqMRhYYeefqtdqOdJ0qf
RvkVhcsCdTRpJX7CcvJn1WuODLCHp+04HLxhIozX0AWNi4nQo2FOHzz7197ZnUmo
HO/XPHkQT1VGKPS+JhEt+ckhj6qCYOr912yTZThbzn0lRykMTRKssqnkdOocrqtE
fLhwUwCHfqsuqMoNNYh+TR1vPfXOSjwrb6i4qW7E/x0f+TCaOGLAiRu6/M4drVHc
MgADW3M93cgKhRHEiTmuY9b70FQQ8JyiLt0ZN1TR0LglsTMBXg2SA9gxP7tDyAAC
0ctMsKnOGqtk/mrnY80Zlbekd7coWT6kjumuuMB66Xh1KzcLA9Gy+2WiDrgtPmCE
bMkunzfuRfOaLsRxlrOYHG5Ea3m/LkSX+Tq/ZwCG3/IPecaLW9qflOkvC1UmYjGF
sjg4fbaTcBsrNdgI2SYhcths1lGCKH4HVwiYP3hjnuzc2pEg6MnfI0fdfiEPwEiI
bjnth9vxnuANCYbjjCwCQH8APOF47S041uHHn+s291/woaguEP1Q/oWi6G/m8Zxj
3eplu/a2iG1vtOAGxnps3wTPKMUxzVq9cq7DhNvh2iBVPxKUpToaxM+dWpR6WK76
sWTjtjSEvp+HcUuELWSWAmLkjkpRyMx8sXyXyauNlDsZdXncb+A+UOD6m8karBlP
p7zzmcvKO7H07zgGSPggperAE0eaiV6K5ncwij1oDfm6hwQKIw/92qNcXxnZBnvz
XDW/aYwF6NHjqmbi7yEbkGJ0j1T4Z/oNG9O0tFFZFPKsDQVwXinV8BZjG0l7yuRj
SCtww3/9dI42FQp6MxR09o6j6uQrbpJ4LGmZVdvBItnLPM7cEUk5uQwSgtjInLNo
QK6YZ+WiEnig9uapXa5hNSjxuXaM3lyoAxi6rf5ZuxspSzAG/ItvNdAsrXng8AXT
1L9wUIT3wqtXRrpO+0x0/cdAYAszwocfBknufZEhIT1yDgFGgNfjx8nvPmU9z8Pc
QdCRe//Q/TZT80x+TLrbz9I8R1wHDBoMHCf48q3qdwrX5HwzqCSm9hstZudYjFnQ
a1ZRZae5yHDz6Yg8F2OEkNpRJ7sLSlL+eZxYelvc0iKXk/MAh5bCAZjOAdhrKv8s
EIHk4BvBrVEd1KQxThrLVRuBWvXUU2jpQg4vUck784fXZBtSn7eAYkgnr/G4SHi+
v7SYDCecEPMHwMpE6QKUeJcqEg+WryrEAEE2ZtUDqdrQCtKdrnR2wlNZwShhyLw1
Ud9oDX/9m60eliz//U3ohmYs0SoaU1FzlZ4bviPaMAuBNymhw0O08Cl676m7uSd8
sCi0Gbhpk8Zhfymc+zb3ti7JAtsUH7eZZQtFmG6yu6EnQTICNnFJPmaNZTgVTqrU
BDwjwqL04bajDd+SeBtaB9kp7LmPNT0LYKbH3rkOeV4LAJegL4+X65gouyB9KQnj
Hw+SN78hVq5aLOSJDr1LOwTR8RKIMecL2h90F5JVvYnWzivZwdJ9KNstFCt4GEVI
cNm5SSbrHC3MDUMwmjqhaH3p4oEHTrLUt2/xMmmPuG/LzUcKh2lBUzI6UiAsw13b
X032oePNQM8osSemDYHGSK1f96Besrsc8Ln2OrDXOHSgtB3VMHwIJDusn7ZeBrl6
CwNT9BmcCgcsKUTSnxMGZrdRb1lcpuT1N7Z7oC3QPVSw0HT/7Llif8SrrwuBC7Fx
ai1KdrfrhFvfyLcsJMuvLqOosALWxI11So8KHpZcpv/6rkE98jD6E+n1q9JeZQfL
Rmt0Smm4AqspFmiwaoSVo+ekgSKKVv3/JSKYyWGmk/7d4Us+h3Izcyl0mJKFYm0G
tkRsqYWaJdjWCrkL1ey5QRhegr0jTnwITiAoIYavdHROSoNcX7hNOP/lp30d25fr
tUr33JQUybazRMWw6QDhhh5GVA9jATdZliqn1tlyUGHGrA3NzoFdID3n5dnBiAC/
cID1D+qe5FfwLyjTdixLvbg3sw+It7WdQ8Ymm2e0+98xEO3ngxu8/VhgECxvJ342
vX5538b+U+lUPZdhcIODxuZLzoWS66IJSGabuY+bH1eoj+7RFO45mFj69sBDMbUj
BRY7o3KM+6kkoxV9L0P55TudMjLLdb/N9epmRLhvpedehTROor+hFNWuCpbHFp1k
D03Kao8y6WBfzrH/f0CKrN3CRi/k2eLoB0Cbp00FIzlzZBUgcuR3Xuh+Bl6PxH/f
h34m4RYe5Waf0VETawoPlaK3MglUUCxASzAA7FfcfKAlPO3Fz8GwZkXnGLMsRTK5
92AP+0lwiTeET3zdMh6GLFi3hCuyy4wA5bDNHyaWRLg+9uDn22BC9MOGgNxAmusE
7Bow7iR67XqXV2q+aZcXsNy1A7RU5zgoywO7m13cb1P1xhemjXwYpEEo8ZakPZhh
eExv8jAbhglsRayMsnM2l2Q+DSwvEx0hZlV/NHhG6tlpCTXYzBdSrHnFLorjyUlm
LQZ1oTX1MHztAxUlakzcvk+JToOKejjsA5r1CQw2P9eUe9by+E37eZEqbrVgH6pQ
Ieu93cash9mYS3A+FB2Ie5hf0tlv9rMVqGTWqEIvR6mQIfh8UBhOFBOMDPgtrIR4
XSgDq+E7pBw5u5GcVDjQWUdqef3O0+4G5ha33ogBtfEtdbd7nOxjwTUW4rmI7VJQ
/BSGCm+JQmoyFy8TzzYZYbTGXDOc2do6Ln8FwYSdef8GA2I4XycdCExTnexcf7J+
V4HYh+SUAtWv1QnZ9BEtgUVXzxceJ70LVIniq7JKvNXgglVZbQUgzQgk3wWO3DmI
W9DE7g9+UnzSYIhCvZMA+RtaHWMTr3r+XVpMgz+m3+SB1FvFJtGfYu2HuK6RKYBZ
V7iwe6IwQeZNoao4nsf8U6G/9zSfa83g2YdPViPS3dagvaGFZYSru+vfCeqILCi3
g0//QOekok7gs3zuiABayV/TRI9RgnXvumtfFCvpVBtjAoEJVgm1FP/Bd8PmaP5R
SnYXow8hvZWTPXrGW0+qeFRTs3QHRd7ir+/iQWTEDSPvkenr+V+biXOa0m3sH+Sc
HWzt31ygQxzfS6hXgzE4Xd2rybT422xA2UTnHiXg91d4Mhxn0huSzvUnNWDB++UM
O8OvfqXSuXeqRSzEMoxge9jHcR0zZCt+qU5rAdk+ChXbRedhqLQGsrXhu2Vuk6Bp
W1iTXqQybiThpBUFwYcIk2PQYhCovcQPcKVKqRmcWLr4GD+D7CyRgyMjf/NUVCvR
aCkfZe/aaHRSu8PO4MAnFTwzj2+1XSgAV6vE9/33dOfe1M2QwNhHteEhBhpJFibl
ZtdBzS+qjCWOP4cWBEIXn0rHC3z0trOJyR55gQTcXqfop7T7kL0EXiMnHPhc8tHX
SgLO6gFmbV26Kct7EH4N6A5cxsvbsgp9nKxL+W4n2VAnyart8akjJsBYa2cOoTg+
TZ28Cv+3LhvdVry1f1vEYGDb4b13uS6uFFWvx6zquSZlwmW21aJzxQK5Ps+4zH39
PiaBxjgadQ4NvtdKL8RB2Czu+qDW+QFnQWqh28RIExzjIEkvMGvBtCWDJQ/pgDCv
/lUicpZxhSjP+qkiJj1bbmRX+QlYw0QjqptY7oiy/4GW7AObg5pc7mforhWvcEnt
xxFN+61o7/azhR4kiuSF0b9thgp/hpmef27vOBYbJQ8c1x5tPT9PbTrlnGFFPI4/
1h3U/JibL1/oOFgAzpvqdVGruqpV2f8qn+KJ2mHjDnW0nnfwii0nYaWf1ngs5WER
micvAcINNLT/afmYcjSxUSY6MCp2FA5hQfMviFYoXwi9bR6Rxftovxj0GbDPsD0e
rIQPwBz4omppEbjxKT+4KC3A5l/50zT2HE6QCBFxGAQAsICyx8MJyuhtoxm9j94P
NBhuXYJfoISZzcGXvPCR/lopXzO5/koUrX16W7S5EIbDaZwyQ1+hHdmYCl9WqpK/
xMOajHR2smRm/fkm5Fi/XGxYGddqiDYSBYr58JHi0bClMuji//uOla2Jo875Y0fB
F8Nc2BlvMKEsaMH/e5CF7FAGcQE/RyusayKwKGOB+BMpwClLGVyIzk3CVlQQh3VJ
vrU1SiMkXVK6H8zJlH0tuV06K6igkBuItz713YGWbUGwCZYNfchiFwUoAMXysyXg
ptAYCByBIjUwXk0Tcd5yVJHqcTdIPxvXE1GF6XGVvM5iWpL1w/d2Wg48nSI+zBQE
JLJmeqU1gYXPvYlZ8xZxGNON8qITPGcXDpBqd3lSu167/0w1s3ejYzlb9woNe1j+
j2EF0NX3S4O3t+FWxNma/IH+0nzUghCP0XWlOn9BAK5vNmA09SgpXiDmHPRzsq1z
K1fsmmX/9MWvdtB7bPpn9w+KZT71HHnMraKNhFMn+MCNKmXGfCoJuYpJ0AzGUVyB
w9f/XflqmLhZIbz2hlkXOeaFwoEJSpgx6Q7OXQXn+jo1gy34tNG+ZbYGS4RZ8JzJ
SaQrWQki4lbwdGDO1qgHu5NnhsSKQdlVt8PhJi/RPYZzLaGXdmSCQ0kIcv9s63WD
aCk2LzTMxkpex5hm8A5VX2iRk0b7lei86JSMhlxsGMNtIR8cnRAU5HHxzoqfyoWD
R5EtKKgkkY8+lWjvmSWSNwTupfsfhFvTDRgtAkCHinkOZDgNmtdnyYwRsLjD7Sum
YjsIZhrZNwN3cUxaf4ev0q+TI89bQWqki06hJ5qdaVwhmAQsm5Oz2eKi809ezWsO
v9oSGcW0/YXRyoJGON2yBgHUjrx0vkYv+mQ/0JqZ4/994h25kJFtsYHmbkLJ+0dp
7Eq58gemQoYNn6AqQRT+FGeeYlXpeax2j5FG8fZCQFDpUcHPTGz2unKL616VGWrf
Fu3KP7r8qJtg7d63Va4wehmSUTJ+Xv3MZj1qZULSABuDHhlajEifUytMWzGrGFxq
2WBDbnjeaBBerpzp8n/uEQI3X+/3muJpVCje7lEoriiukNXSzMg1tOZ7VTYAaW+S
WzAAuVpmMJgc+9JgpLPMryQdTiHCmctJ4Nclvb5sztTQaJmjwr//FBjjGLDYNKsh
DN9Y04oKyFcrmiWd6jnQqrdsLULAqg6ExYIcCyCWGklq1F+noXwiaFq6MJ5XLpE6
kHc61IQMMxyU9U6I9IDQTgSCGSqoE17UqxYXrUFMQZpvgimJwdc7Sq5CiFcWAM+N
vWVPDty6th6CAEFug9Cklv6nOUcPIMdjro+GCfSKyYJ5yWkkf0XRpyOEw3uQYdW9
GYgIBFm74tuUCbZ4pEBjk6dr5X0ufTYmsF5ncRHvRjNTiyBVAgavYJRnXWsnGiLc
H2apgLq7T7Ec9lmcpZl6QHgFDlnQkuVJ1rST3y4eC4C7QJ7u8jL2QmpmVo/3eLlt
BrNRW7kg3dZODmH0/JrkqcSbsYGhU6AH5BLtclmnBMpdnt5CRcxBs51FzTSVsD17
8g3Fg7K81Ujr8uoFwHRGtfLNfUdyVVIEqkJ/4or9GlgQ8TkOWfIaO8mKIkX1JqPG
y1ZIWrkIGnqoZQ01PhA0HRm7+VCXrmqWkikbl9gxrERWjonCeYBPakQE1B/aoYWt
asx9KezHM2kkTCncyHIuRb2grethomRUkMNmDnBfggXH1im+tjM/tyfCCd61MXno
Fw3CAnCleHu0n1mV/LQj3QxppaX4901eHcCfX5UJEtrGkNnjq7XKfEoeOItBF7Yu
F1SmE+ay9i3WzflpvzG3dFxONdTnr7k3x7lkBLRORm9dZCP7lidZyKX7pR7WA5Vh
oUsDKmeMhO44HbWuHMbjLWkKMrR6AHGuzC8uhaA1AZd9OVYMWLAdhg2Hdr3VMeMy
Me/9eGYVyT23jNru2rsJAzMKg4ZQgbkAvJPE79X6Ytw0MPZPFf2Tk1jBOAaBGxwV
/63zengvhWsQ/nM9Lmo8+0yZoLxSfGIdc07hapiukluBbWxKGHlasipFuWN4Uvgu
L5tSnaCQ//8bPTlKK3n9r9ImQ/4ghm9nGN2YxHcme3kBl1UoHboUYbE8UN/0BbFB
ww1rjJJrG37dXxwWHvRsIxMp4i1VaVcnO++AfdM+zT/FglRSt/wWMHLg5yYhWVVm
coEBb01fWHjsP1rphyJKIqVVBv5dpQGMfuwjavTV/qHemoG6WNkjHEDaB8V0aaoa
k+ijpxcdQvBMrjwFLZ4b/PoSzdd2g71zaUljewJ/VVZdurcMQDZWr/chRoj3qaPY
FloDojPreBRKF5zKH/9ODx+wQkDBmq3hX2aEFAN+Urtirgdfa5edHyfzaY/jb5mi
VMdQWkuKyDMEJrnESxIUZ+Blr1iXOlF6PYKKk/g+tfW0ywWHC6aZdHcz4PeFlbW8
p6rblN8fTGlfJkyoH5bZgfHAMyoJI/zgUn0cryoEF+LPQcZEChDdc6/bqHuPxwGc
8F5ScRVtuIzX8zwVEYl3ShdpY7nP6SXW5rlacczo061g4V8Alt0OrRNfhJ7eS99T
30lUeHm6gOJjYB1ElafIaYJDtMpu2N+efDB++dt85WOJc+bCTNvexwwn3jXIbNUf
A9BFNN+XOta6A4zCOrJPZQLqnrwh/uMvXH5wfmd2hrH4ShJw4lrpqtPr34RQj8I1
HQtJZihhBSCjwa3ICxGMyCx3wyW7EEGG26uAwaCYFE7IRGuGQOQYC09WUfFIM9xp
omJ5lCDZiDiTDU6IXc0UXjLtBTzodveRXWNB5mI6KaCar/D6ICy5k3owDh9qOD+W
tt4Zd5SbPdC5VMr1u2/R8s4YogYDJruwlsIEYHd19DBZdJxfi35BOPeNYDuR6tO2
NZcSyOxtiiFbBKPxpvFXn87TIHJToJznz/CByHO8Qg6G1smD8+gV8FCEJJ/HxsOQ
hGfMNz/unx/7amXohR4GphZ802Y/ZG6x2VQnLAjkeWmUdOykXyKk0R75nuYduxOB
srwBlrsxL0IqWUDCM4sGQIAw3TKZus6N7cI2RUuQP245t3HhgEsFmr3wJaTaquE2
j1A7HJJZ1QuTeqasZl6hblNQDfq5LW57bFAe7s0N1wFyEXPjzxuy0llcupPSBZ+E
UwKfY3yhVLmlq5U3jHRJ/bjvz9Wp9ofmG/duKT13SqBmso3JZIQUCgnDXzZwmvLS
ALkN+EC3Jm+ouaaWXvfCWuP4KmziKYkwCGJSeCM4SAK3FpSWBCHqCOIjz5NHA2Ha
Ft17DhyBjDMjUsbXjsE1KKwLK/vbujUliX4EQ1UxfrrlGwkq1VE4GzpUuX6CXkik
VVd4ZoOgrDZ7play7F7b9zVfEuacNArdDMP9e6vehFT2OwxuBc/Q+O4RyEyUY75s
mrKKr61/VNN0LpjZwUekBUWNztKmOdIahFFJJYdbJXN5eRCi5n4/6/3u9AS4c09V
E3faByz+CWsXvs8AnQeQGAyHEjCK6XH+DOu/bQG94O1fWiUIFPVF6e9D03MrEeez
cI/Jva4HEcUot/32lai1W8Yb1Utbhap3awqHp0ess1YLGXxYbMzYNF+4ZuJfXpQl
e8N+VNWkqadBcpIBgG3l4KJx/0bIm48IKGJ7+B2FNd95ruT6s5APkGgbNPNkiF9G
KYMn5xdf7g0HZXVqWtvtKyhD6NYLZkxbeGBjd7HKzmWWMHTA5QDxXBFlGs2A1tJl
QBO9PT7w33uM3kO63tMylG5KTWdGo8e9dXwnWEJEmjW1F2RYQeafyLlrOjarvMbP
JUXUwU/B7atInVhSp1dPqiThU+P+gTYzG9D+mS4dpNACY9ppfVOTK13QFvSxkT/F
YPp1L24sLYeUwWSM6HihY9a7xCcXgPFjTI+biidsVTnJ7NDcBQnKBZYkJCrjVbXJ
TnG9IzIjsuzzv7mprPnGoIojfPZl65xXwvq9lv2V61WXzes01SC/zNr0VjnfaQl5
X3kli848EzfSkGt6CNKboV24FbjRAYWQRaChtR8b5kskbArRVw9Yd2BjDa7tFb+s
rY6J2hHruqvlpUgqbJ8wooSCQUEtcz6Cn1F6s/ZoYKg6lCh1h7YyIQgTb/Q8V5sO
mevQTVxGsUnofhy/QCagM5r8g8R51b4658QOBlD5vPsq1NIObHOGfyFgnLN7ieZo
oKo8DS6UJK5F/otUwKAmC7sXBqY68WruzLPzCwRF521K848HJObCPVUIcnpVtwx3
idITpY7z9wNgUpB7xJF/NNCSTZK0eMADwwJGc1TXaYJ9vmF7QbdmbxSe83M6dsM9
BGutOn+q2NSlDrOpYeRB6P00IpAOEYJs8AjDhcxx7zeIideOImw7JFosc4aVvWGQ
HYK5hpSGyb6OReN9p3+hyobZP5M0UMnlEHXsdbFp5Z2j6braW2ZpkPxGQVwj7u0v
SsRloV9VitElFAcWgQ+Gu6DwmUlhkk4/qVyePgUPZL3DvRqf3Rk6ISCxRQKcabg9
c8EY58TSgR2Psm/1Qe1B/Tt+g9TOrchul4QgDIJwhTUxDLvQYWIPZ5F/KBEWn9Nr
3dLfAR7wpe8bwfQDa9hVRl5AE40epqU144I3gRJs+QhON1ce+u2QzhoP38kEBvOO
f61EoEFkzvhyqo8qLnelZ0XCmceVyy0J6glmnJ7bKXOAKtjxqR6jUWlD2OgG6QPA
bpsX01cWsxqm+VsVx+tXa9VNki7stJViEfsCOaYh0/Fpp+BzLPX4KuUgf7Xov/wW
LeOb/zbFVe0n5h2YWo84W1bXH8uyoYI6wkIf1ENPut7UrF6IKu7vaGjqbb2wAEe4
mTLjvHG74x2TdjT7SErAFpKzry0GM6rSiEtDKZr/+VJaG522YQtrw+cNZ5ss+bL+
HsFOmRqI0udMbc/lKtqvPEj2i5pe/XLFZ8SZoyNOp32++yNY14X9eBHyp5vWGDiQ
cuoF7n1xzwedGu5pv1++LIZUx23NyU1GYYls5F7+HF/PhGtPtZYfU192XuTD3msi
E1Kfxb+qwJF8ycS7B3SlY7d4R4dmlZ7F0Hy8OgZC9BtIynIOtRwoEOL3c5kUAIJR
oZ42wY7e8MP3jrgIQUlgw7woUBdsyUt2LYCisUN67e+k0AuShuWB4SrTPkWv/odC
Ntj3pnKpnDtY9mdd0n53oD9z9E7uBeIdcKfgfaBjM315D2km4O77palBWyo3AVeP
hwvOK0YBjgUZFVJC2lYB8nePZDk5htsP8oe5aPD61ZDfLAlxXDGfZoDSUaJzR0Ah
6IPcstuMzE9EgTmHK9SXxc6B4jjUDhp66aDusETSq0yYXWleKmW2E8et/LdVLsug
gEjXqKs8stJUmYIjQTgoOQevAwMYtYQVog/DGlkO5beF2GgjruvP/Se9a8wK+Ykc
W32R0k5e+pvvkOJO83v22fJ0yRQXfQSeu37CLKjiuSxmJD3ilMyqv/qgnnDbHHqj
u8Cl8gFGmansLBXWceiLqAkbpSsiTYR6CUWvCXsDSFVE+1cdqOyvTsb0/BlDGcQ+
b68t5YNMzFHmf8qyzZlcc6tCXBWPgF07nRjvSQ/4u2xvnUfqEk/YgmjGgm1r1++S
IhFbtsszXmGz1Dbl+sVvKr+zRy6zFqJOdsxEArbWEkLzI3OdHPlTgeo7fi7KVX7b
nknB+nVdzp7Vq8orUNslXmIjcmde14PJxrTchOTrh2ooPaexomvDgJN2dkoOHIKf
RaxXmPaRUgskQWpjnE1l5ofZJz4uUnHAl7r+ir34U6I/hYJMngLqvdz1WPUBRvp4
TLkqBHWkb5niVw/rAHQLtqyFJ32iM5pY6RVc33drxKR6WRjWUbDjLHI6xaIyPwkv
2w/9wtWn6ABtLEFImIQVlfSm2uKDrGYagOKb9ZvAZ5mm5Yw4rGYsxvslg7RQ55pC
VbttQ7cPWEKAbuZK7MyzoL5FiVppjbbAvMJnPJPmSZly8Whmq42jDwKMywFa7MYt
wAqhPxeN1OT73wELJmlEGmtPDPQqkEOCD3UrF+9OXXdm3OEJqYz+9VnF4OL99HXQ
KL+NfWO42sOeHSTDwYlHyPvagWPqvIRoyVut6xG+ntO2E25kZkaf9iv240lbvKC4
gUFLojEu4KMFCa8WZW1jGXrvaIrXQ+daucMpcb3kY/e0cJQUX43jDCvgxEesXSQO
oulVNhEHmnmL2ebt/dgiFRgqLUTy/H0Qt/dTsX8ujK/mWzlbfE1xprhmWofuB8mm
68AbHfqLnYzRMGT+KIzSzU+4ephFsngymiqbUEKEj3n3uX+9vEC2QIQCFi4rA4fY
mrkVxQrTGC/+BKGvVKETmEud4wW0KLKuR6h47kP5N9XXkp9OgoMUGIMlvkN96V4J
sEXqd1ulXzoyjoH4IYctIsY+0mNC79UAD5MVtW4EntcfaTmJnX20Ls4eR1D9Grw+
QJHVwi7pfxmYP7n6D7eQkToaDUa+OIPIAc1oIrJbLZzjyai26H7K2TzQx0QaWKAc
uSgfZu8c+gaFPpKyCv01GR5cNoT8wvE8Puz1XBn8CtH8lSoefME9j6zthzCw8ZKG
y+jdDecN+yA9E5h009NEyamlXbwQeGJsFog1MgVxCb+eaklZCvQyXUrflO7t/pSU
wsKMYwHqZvL0JV6ThhGvOT5Vl2+/bDwJX1MPK6yHwN6sLaqTNiALBJXeMIYnThIO
aGSIlwlYEL23vsBAdJ/evB2BQ+1qBOunbvf1hvgp0YNQr4IcwLu4hpPpqAyMVH+6
26DfpdG1tIPYUyetViMhfLd0QJ5rFoKFAOlfF5p9iqQGwbybYZARUsQ1mCYgL7tb
aFmfMy+1r2i6bdZDpLDESn3urq4DIuQEkH5cglZkqSq0PqC62D7pMxoe3/e532dq
Qeci+9Obe8DVfzS4eAa5ka6l55wbXksO70p53IhuQ94m4sXWH+jrZe7Ck7CJ3TI0
kNvoUcrBqMWCWWrKVycy7i/MNQ3twW/41VLZWXBIsMkinfrX9sTq7spkO3ACWM8S
SqYryOJ2InH+FcYnaa06xA8HBuGoC/Du5wfhg2OjdpvGQAOY9ysQ51eLUwYHp9MY
k8j18tRXG0KV7s0Eg1aKhWEMZIcTONezwDm8/F0jhmqBg/v9VMIn4WUf91J7iPkI
EYz10nHCMTeg8DlG1PtDKopRl5aPtVDNeTo8BLIr2+KlEk4Jge8PM2LadG1VHAes
e8PRGn4WyQDKBy3LqUCJ+xxfm00UnYKqor6pDJKOL44g45IBtFgNHPZoKXMT3vgg
xoZAh9Ns9MAEFXK5fB4f8wW6GxJFylR0LKiWjixeSdEEdiP64fs4KNG1O4imjkYm
0c9mJQwjXZL58q8aO1UhTsRlvcJsCfDrf9kW5sgqBxwJyTtqLYpiypTBeVc/drUu
k7UwbZ2rqm8VcgdZ9p3uZA9UYGB5wD3QYmpU+hrtzGjdReMWaMvyAaBaz4ZYRwIs
ow1svHuV9J65SZvQdEPSwF6lTXL13uz3a9aIJG5cnj1uB6SgB8ypjGBWe7Etpjb3
lEqrCatsaY+7AjbmxjiSCv0V5vYbT127xPT6uOdo7LjONkHGxuZqZaKX0moep+hi
aEe8kaqhRtEUOTvwqh3tPPgzr5Vs9dqzJWOD3KyJl/Wki4efS83tknGsnH2CUfmn
E1PqBRqzSkcO8pRlFUIrwh5g6tnXw3g9uO1C/8fdY6/ID/JogQw15rq7GxC/z8hs
M0D/CR0b0ICoFJyV8j0El2PjPnnrQ2rZIxAOHEJ1jULuELF5EF7eJ8Y9FhMvaCTR
hUZe8Ih6HUnkd/UxsZo7hwtlt3q1UKaiF5V0XX/j7umZckj9Fb0NsM/FwK0FI5tM
X1aIgkhPnMpKCYm5ZHcEp59xZNz/E/bwxarMCKFuy7IyuxAEBLCnsocD4yMqeIJ+
i+mAwlg9dgCdLeBxlIGSj+p9itgZ06Tqx4cuYMIgQL8nwLPt6rNomD5bE+DwWT6d
zyPKZUtJxdUwyU5ZQnA7RwxeOBi0lhRbHAMdXjmnC9w4AwgV70F8e7/GFbK7ZeJF
AMN6e72nlFkx+vVXkALCN4Fw3+l4B66ozl3tez4SiuxQWxdVlCDqEYzRqMeJzvsN
LcWrE+hREiltrucXc7ibDtmLEXitjWnVfpjtM6anyeqV2MpZFih9CAhgMUv7C+nh
tO9/hoqqYCb62jXEkBen9DERHHxZQUPBN5ZY6p354ZBSSnKdeUKA3g1igF/mtwX/
RqbSsmfblIoEh9++nfyRfh+vObLwNzLcvzzl+Hd/ENsDzkvaL65lmh2RMl+4ztWW
/Aqh9lL+VgIm6zsvbQK2qiFzWnPLExAo837aB+z3pT6J2zMfwV4mLOf6wnjeYyma
CSQRD6zGUXO+G+Jp/NL4TdvR/cNneQyxzlyEbTW27rbZ1qrEqaRzQ6xtzle2BRpQ
WmYOXEms8DMmigWLJpqheDYi/1gxRPN0kjC0Ypn7r6/I2eqo6f/R+ziKUJs8UUc+
PPcSzVCAzss313Bu6Rn/s/4QJvJQ9rbTT3Ytv/iy9f5TSpnfFGlV3IQX+UF2SRrg
1rdnI+EZ53Lzy2pSSvPtxw==
`protect END_PROTECTED
