`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C1ZhEOaXC+BA+UzucvEJusJcKr6/CdBAddFfzG7Dj98P
zrZs4xOcPh144xE4VQ0OV5Wj9gUuMU47AFSW43i6MXYkCKpzjWCWlWwEYRywH4Mm
evbgGo7Ixqm3hVHFUBje6DuH2HEWTEVBreUfPloUiXgBZE9yHwtI0JabO6Y50iKC
Jne/ka7skJdeN2jYK+Qj8f9MjiBhIV7MeGEXOSgvki/pWQFIHODowoQM4GiDVrSF
C5iBsF9plp2y6Rt7Ap/BIxwv6DVTqOOetmNnukqkmfZDwbMvlTFuzMdhMC9TuxEj
XllISa1WvaMLR2rxJhZoRk7YJmZMJKHisAnoywQ1E42J3h4LGOIREH24rcZVtYv3
Q7pAuLuKh3a7f3IXgX+Q68OfzTRBwD3Yw3o+G7FCaTgjmL2EvTSPBYz3WAtAdiBA
B2Mdv4lZn5HZZNMQDl6qI1DpmdJJ8iuykpIJl2U+4z9tO8+m9kNzILZsY0eDtIoD
J/Q9zL5dcFc3YekRV/7zsm+LjStGR4NnHNKFdhPqxl1GAWKSNG8S5gR7QV6Ohh+I
eZ0X/NsAI+UF6mKTbEiwREMnC+xRSYe6wROwzYRaa4iPVONCcq81VOMa13vjEjoj
9fK3uFXcKQL/tSLZXAL2b7S6wM9hDSCfJ+LkqTx1i/8F4EFCJFVfWckZINP2hHz6
`protect END_PROTECTED
