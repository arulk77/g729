`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
y1d4abfL0XrPTolgTKzgbljDiwVZyACd+S1X/NOQNXggd1X2pMyaRNxzjnXfOdjQ
Qw0Dui9CMKGlyV3KTymIsjuiD1yxDG4/OLLuBJHvBOgGXvHarPdf/i3rM7EdLP1N
hJqvA3EsNCUA4mD/oaOKcZ0G3LPzqW96Kkzex54+XAYcD3RcbedNLScffHF1E8gU
OTCR8WswQLWMkWdY7O91HtjudITmmvvfB/bT15dig+H2woNa1WPLscfu1RrHp8kB
L2bpu29er/DLgHSM7kcWc0pxTInmdk56cmtBJo4hRP9eiaIKvVNSgszeGoSZH8T0
fgqdu19LLtRHsyCxCKjExqbTZlrI2q3K7+0fiEWBZxTwjI2DLCdO9TpWpm1goSpU
zhKuWXBNMuWvBBWUwWLYNeJqMn2aBh0ILoqi1VBZsnX9FjqGL6ZG3qXcKjTziiRN
2W2L4xRoJSORahVs+d+J3ZGbOdwXBmxeaRLWp6XDlUPIat1+zMUoDGEuGz1qoDL4
rpFl9TUpf1Num3re5i9RMQ/elBoQYGiwxto0ZyhhCdBcEHDFsYqB/Y2FO2Y3ZFcK
mAaV4zvZpxum/MadHD6Q8yXCFFqIlZCZmKXKXa/PhilrwyYWkjYDuNpcXVMRRPcF
gAeLygJejVA3kTCE0KkjhLgEaB1w+NtdKZLE8c2bacb+ge70RZ50w8dmo4OrqPGq
qotmKbb3s6cnI/22Y7AX+g==
`protect END_PROTECTED
