`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGCkTAUoHgc0AYhVCyXDm7ySB/hWQcftYhLVX1LmxfSB
DCu+CmWVH5N7PbrF8czmPD4pZIeYWvP2KhUqiCmfUGjjTUONM80xxV3o5Ih1IDtO
p7VHbIbncgEAArpHmk832Khs7Ysg/HrxGBNgPSVzX1n6h8CKlDogQdlCT/3GA8ku
PNkXrcY/V04gDv6BGUJQlhCcOSLxjas2KFUzmF/pRycwYBNdZ0rLHXGMRq1uznI5
KSVIpVWvD+6sYWlAlj6O838ZMAzmENzbL9Lp7LzRPvssslA47nmEyH6Px6LXJxoX
QP9eKEq0dhfQQyJ4/fTJ029BVvt9OtlLRaJGkzHgUPyb5di7CwK5+XjfWCHXjUq4
RMOdNQLQCO9BteeUMGOKfuNKr2W2m+6pnTPkzXwXlv7xL7yVWom4wx6Oe3BnlRdg
o1W0risBsI9pCLeW08zwFnFMQuCcCV3DFk9JE4mjxNLwWuZ0S4U8b4GQhhBvm0/g
3vHoCFyxBXmnEXNl0QTLG+w+IwIfMXSdWordezQnsApwVYYz6j0khvGRqsl/Fwf6
1aEYzMw2XemrmSYnpbeGZAvKu9kLzhIHa6cE9X3pPAOSuwFeFnHLX8EIuCHFteN+
M6go4pTlezN3xv2bhf9yRIyyTLhBzPtonCltMIlnnPpMmRywi9nx4Yixyb0maSp0
laXnGoEd3G1NBMdDSFW4Omn+xX3FfLIimotz/jUpZpKjKaYuKRRc0GY59oisTgcz
HuLibc10SueaSbot6dEvCiLNtbI5DMfkFoI84gw//Hg=
`protect END_PROTECTED
