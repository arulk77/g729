`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHZ4iAk+EPZXC5YHRGXIJL9ImLSCrCzzMgICc2WEApqi
c+28dII0dLihRt+rB4IzRP9YSKxkSxaWBBH1ttK70LYvGyLdZxLPbSWZ+0qi1Mxd
r5H4BmN/CN0Tzv1ODC7jGPL3MAMkaEj7JsR8625G/2OaqiVG1Qx7vKrqB14WNhNf
YOldtZ83T2zyzl451NABuZhYl84S/e/8AxyvaJ5C2p+u0bmuk/JzzGseFSeM6gwZ
r33eiBvgN7FgxRJn6Zzog7H4VgWM7qWjHyBSSVGVwngFAU11iUWqtMWidU7SLlaf
5XqsOO1qbiOtJnA64fe2hY/1oPbcMTIyL4A+zJdqEgt7BLh3qp1ETwHFLLdMwjkI
GXAFTnXjj/1x4dSWwfHC7jNDaTFWuZ4g6DzlH3lv0aPaoVb6dpCHYR5cs2oY41vU
njrBCXbYVQHtnz8ucAUdco4fTLYilW6SdCB8TLOhKdoponVrsfNY3OZyhC4DqgAu
KWUYB7erGZF6VKowrHIhBXHoUGTe3A7SunHQfNf3Aw05yv/8cbru0m8FHJCfPyok
myC58OKh+733AHj7QWaa4OGxqBO74/BLJaWzN0QO/TxEccAsfU769acSKWfZHLV2
PAGLtOaaKUdjznaYlF14ErPz6VaTZp6gBg61ph4Idbc9DrsMP7ymInQm17Nh25Li
`protect END_PROTECTED
