`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLztSNUybFEF8GROXzsHq4GBViaijnJYMnQxfVH92Mbj
Q8xFnDWRWZDiw9ZC/ivqbOBw548R2Uq5CHRRK16SltJLevAQ4vWp7EPeSYhYL9y+
sGIImmIyZ+9JDfwVPMdIeYqoWAAcQ0kvv9KZ6O2LNpoVwhEiCFEKdfQce/Ggxyys
`protect END_PROTECTED
