`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
5Ve3PeZ6UdMVjZB7s6azwmFg6onQbinxrJ0yP2E/VQNFjs6v5YAuxCAh1khVNl1O
AQanBaVH9cy7taeg4YoRvaAvfOZB4fZCl3onKYDt2d9+xl5CQikjnNs/YjZkYDVw
ufFLnR1YayfNJWIYbbVJQr7qoNXrarh17YtYTIDl9FMPK2W/6QTOpzsEYMOKq83j
2D0YTPdKGOpRoCCurWYaEPKCFHbcAVQRgXLhKxlcSec8O+ElX1gg4ih/KHzYtIeI
yxNFB9ygkz5JuNkl/uD12Qr6rabJUjXJmE2jN7frZthLj59U2ZQ2aLTNMYexYMhX
5BKuSfsLPBqr6HAENOhWQBEvMYlCVyDDNRT9bzc/vOQaWAGp4DGUHJ/lmL1z9SfZ
kpMMEwB1/T9nLeuEuW9pmZKNy7Q2gWWkmRmKjvxslJA=
`protect END_PROTECTED
