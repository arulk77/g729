`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41bY3oXy7VVeQGXojz/aHjzZXZNr3yCOsEv5JBIXHoTh
e9pk3YO2123dQ8eZbLUduS2J29aU2H35oNJaF772WNT1iT4OnJAQymp1thvjZR8L
jo5k66Cw5xzixFTymvVCjJqyB8V4MvzlPyxQmgjK+RJgOIQGnfXZOnCTGb9wWHd9
GyK58iGsoG0qvTDTLIGitzL4arxI/wgKq1YC91F0qwh0CTKW0prLSW4+UJKZkG36
HikR6/ruPDU3ZtJuHKUst9AjCOQkfa3Ht947h9eMkTRGr4TZJCeKm0Bn4ajIMIaW
HA9teA94E2TAC0SUJnDdlc7RAiQBoHLvbrUhd+xjac3HZJoRv2JoMC0UdwoI7iFw
9AlzLHoxY2k2J7qHn5pO3AtFjtR9gDzxnuCwDMlwIKi138PhghtAelXnS3Mzd18c
m3y6Jfm//UvIjCss9JpkVQ==
`protect END_PROTECTED
