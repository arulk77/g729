`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDVd1Hcg+cx0aQjp1rMGx+dDaRCjkNxXQmSpZkATFiUm
jciWjBvKFc0aKnjHG98PvWMHgdZqmY1pyjQXLqkXbho4y0BBYYEqiCAo5N9/PBxz
SFmuBMvUA5UsluTlDU1TV2TI/Esw8zBrkvGX4GlN2PWAGN/TgVQ1vMWwQBm41ra1
UO1tA1pejf0W5ydLtOpdpV0v+CXmaVlYxDzoZFfrGTx6Tbf1E9M4n3RC+uEkMrCP
z7m78siRNhLnqWYYHJ0+/AjtjPGwbHp+j98CrgIYoDU53R1D9d5PabEUNFceLuhA
xcSILvpxKp06sL8bPftIYXpsqjf4OrZEeMmf6/OsOx9RvNuznVUCRiQQlNpT/DGV
eB1ln/h1fQ86uHTv4CeqnuyKl0wKI45kJKQtNLQNbHYhBp1//oFEA64Wf4mxSp/S
QumizTFwnuzbmpjeVUcJg7VLh3b6RW78ZhujDUNtwn1tDPK5NwlTA0aXmOZpXNyI
+V1oiVXgbMWekGd2+mRNQA==
`protect END_PROTECTED
