`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM4Dro9GKEX8/lxbZH6ATZil0fsHkJPZ/oKV+7qgDIfj
Qno+02XGmaT2PQekU8TnW6xLtEIIFExyEZWlhTLyEDH8oyPFXu+NKIcJlAmsiq2p
YAXtY8sexrmcXRDUZpaxm5KzVGsuN0ZOQC8WSU7GFF+ZsDtymHo9SNCWV2m5GCB0
BMezS1cCl4iCuqECV5hTPriQAl2zBecc8ioSrt6fJg0QTmmDN3rCoattlXu1tJjU
YWW1BBAEpnilZ0eD6iC7Calr+sh3AOUMprwbZ9dhwf9Lw6CIUcHDwe6NT7K/stoE
V6MIzWLSGqWdwOyIyKeMsXpE/mDyoCPDPXXzcAuidERiIuqECiNqYJXOs5OcLFwl
vZoUw72skUvA9chEijQsCjUBEBGGITLuCqBOBM1OsVWmzz5pDUqavNKdvSAKFBGl
U8OJX+15TPA7Sb4SfN5/EBalZwpa2hxwIhOGqyrMbiaA3yzun9FaO9MJqr9B3Zjt
sedcGbf5MjYZ3wipkd1synO/iMQCCt+YYtVT+mJecXJZ8LgwRjulm5J6yEINIw7K
P4utj36d7OcX3mhqmxrS5XBEgsT9ApNVNqeimUNtqYMuoq2fgt77q7WOV+N2bH8v
6AT749zpjFRlxDaUNOIBw623wruHNd0GQ4L/1qTlBNXfQM4mBdRwoWUSp/lHjUbO
`protect END_PROTECTED
