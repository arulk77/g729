`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zP4WGPgrY3Pig2X73My4ylvC2c1GKGz5SMqM8XXRtxb
4xnHRmrp1w69jEQQ0BnlREkEFcBrcnn0lev5jDsUkKlisHtApUwe+uklLjnrocPH
89g1opoRfFYgMquP5t3slN2L6UzXCS1cUVKESU4nEJOApL8sP54w02j4mi2v7G+5
V9wnN8cVM5ePr544wc1z4ETxM2mZHXH12yo+0ryssCPEy0hcp0OEPUWhnOFdRIAR
dyM9CB8uC+7zppYEQMLAfa4i0BeY3zSzNbfpGo8bPJF9CZ8VJ/kjQxr716YjmPDH
xWzf0RDWwPGFQXTSRpTqjA==
`protect END_PROTECTED
