`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47MKYjewgcsnNsa9gwCnj9c9zTuZheieV71EswwNc0i7
aJ67ZgUrFKvMv5YBliYHWqqHPKXnPHV2c9kHpGYM9uZe7BIslNwCQCnhbDl0L1Nu
v3MMG/2VHmLB1U2qYrN8btky+QaFcuE59dSRF9ViF/JiR4UEKaOnKotg6nuWff/e
sKNi4qXX3fQ1m6by9pIwOI6JMFMKWnywF6/7ZUw16TY=
`protect END_PROTECTED
