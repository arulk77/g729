`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAl2EdSsVyxD/g1MVgbvMQvyckqRhOsEJ4d37G3gSus3
nusSwskxlpr2/E8ma2+naiL1JpRuXQKbHM1HbHpMiXkuX3ZX6jrx/QzmCofHaZSQ
sQx+SSEL0oL86KE62HEBMuCwLkwD3SnhBuuNHkS+QeY1vMtBWirjLeOVyohE01vw
bFXt1Zlh6wcznCCbNK6vllxzXkq1cM2ItNUntAj9JqAlG+HPacJ7ouh+m+tGlfNa
/d3mbYkbpU6s1dTfSw3BQ9awlFE9g/6UZLfSydxTrRywfi04idB/MU/0p+8Idrym
A1rz6Bb2jNGwpcD5Cbddo5UGCXbASAV1ONhazhYGD9/E0fomx2tCIKrJpz8qA3MF
aOx7u5G65m+jIKdRxebuJV+jWusApYfRn3UdHNUcjfUgK31wQcGJ1cURORXfa3ie
1rH7Mv/uGC4thE84BqMB5BUNvLwKS0QjrqJlOOA082kYHVMm4KqfwWG9eq7/gdQv
`protect END_PROTECTED
