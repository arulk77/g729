`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFL/1UobLBUmWkfCBODM4Cr3n22IUxgPnZaezjBfl5y7
Zdu4chbSeF+MvZB8+J0KXQq32EFQ5lY8VsJ0ShcZxcFP40SHG+ub+D4ax3Kktcgo
dswdGD15dfDPe9jBIclgpTi4eyJT87sfhaQiHBwq5wtoSPsZln9opkPe5PH35AGa
NFPUsKOv0YhaPgV5kqd20fAIaapwgpz1Qx6w3otMWXuNIPwOza7+7N/Pt7Cek496
XmFueAJE2DbzHF0CfZZ1N8ABvW39hLYBc/x4ZtFVFMN9xxRqjqPpMhjEHikoxkQU
X4wv8Gs7BAuV0cGypPr0pQ==
`protect END_PROTECTED
