`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKptuRERAaOvk1gKJp/GeNZFigcRAl6Mw5Lk36v7NRl9
4tAy/yTHl/4zy8NG9M479z0W4KI1+AC3t3qG7lQqZT9aDv8//8ZhrCKrA7qadak8
SSzpuY4T7j1HO3ndb6xXwqze9COoSXtpoHIHiH+2rse2C43riJMjozn4La3Nq1ta
gLD9L6D0zt7m5YIh80dXkMrwMzEx1b3WwelXFnyaK8ED8SVdA5LXiPTcmbw7PEpz
`protect END_PROTECTED
