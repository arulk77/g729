`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKrIBq6WtzfceHDmXZIFunIMQg7G0CXjwXyVvYcQJn4Z
Dze9dfVfUDUCqTtsPm09ENJ3OU2Zdq4283LXYTjjvvbH8mUbVbWzUGg8IM5MtomP
N/aaODjGHWezeKJYiBV+K1WFM3pnUmeNySOcL1ZB9WAvMhWUH4QhlRIr7j4zXl7n
SD3hAqNhP3xCv2R2NEI7bw==
`protect END_PROTECTED
