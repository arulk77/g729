`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFsUkVbyfWwRpqazO0573GnW9gJYL5D1ze0aQuz+7VFj
svPHotpmRC8eT3yozRm1yvuo2OzAk5X9rXaFfxdfw6hQsgukmRLr2bG5r691gN1j
HR7kY56cSnZY2tUYpSLK+XID00C76rc2FEO+HASpXoad1Ui2yYSzlU2p3cCxU4+8
tJGj+tldGcx7lFw7vhpEMGfzmLYEB2g+o3rNjDHRtH8PSLhsLDx8LZ8DWrzhltO/
yYlSNcbWLlwhlWlNTX+9y25LlPCrNZIfq2tA0z9RsJ1OXsIj7PpuTxiuo0DgH9qb
Y1bXgCibI0a0S/+Y5uSRNiJHQAkiBjyBjaFKS+b27Jy+dOAwDXfKUVC805bKB/LA
YmmtNQj8l031Sd8dBEKSsl1npTWl7PY0qrB0a+v4gh1PL3TubD/SSC4TR/Lu0SUU
`protect END_PROTECTED
