`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFMKsBW+AGJ3v9cqK5uYoRRDQgj03okaLcGg2Xa3X8oD
pk1epYAbsL5oArLreqjl6V95/Gort5zEypqgolN++GFarnI5kMY0vYQdWYxLnrPg
O9qfjNVgU1g8osAWhaTgxMz2E9ChKRo+BYSjujnZFQWQFdJB0PzKkZyFrZ0/8Rr/
DH6YeTdI9KI5cZTuZd8/HD3tKqCDq1S2u+ikxBEfj/Z8dhJCxqBb23BU2jCNfCOS
ecw+5MQv+YL8XDgAYFyncdZEzPED+kdTzS16jxi30tg+a7QliMIzlDokpYMUJDoY
VFzHZHe6i+Afjw3NLuo0Fl3AD35DkSa5QfXuGICVKy/+BFwdvd2L35Id2EACHcmY
6Yl37WjppvOFCCXxKgkJxbAzQJaJx2EUz8LFsVNgilLFBIwgalCoXNGnJkZfOVPl
WZHpYobZa827aE40vByyOpHxUpJvnL6WXw0wbA8tF7AO0EmXw2e2ctKnCwgJTK0F
cXd5OwcBe0TCmDxBPUXVoed9l54DNHn22r6Tc3GtU1wmmgC5pC5SbZ2GLpNwBOzq
`protect END_PROTECTED
