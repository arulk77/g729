`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
laXZPAbodayOq1/doDth3UBLrVQvxC3wAey1jaYIz4HcsQPQqmJ89mhYnW/Lx04k
bTQy8gYszSOJ3zXXzZcUfPMcYb/Asj9k+15FA5XEaoYbJyRsDzrcfv7CyWc0v5pD
c3XZshImHJj8SjOcfMCk2jM3lhdzkosBVj0ZGclFdIs8CIsxloixr1dtgsRr+tXl
DdIJdJnY3HFIc+0JMqoNACDhLIklxh+CLVycAnCBvLk=
`protect END_PROTECTED
