`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
f11uP3tAS38J+2XEq2c6cJ9DO8EC2dg3+2ZuuyUhSDwlxNIptF0QhUpYFdJCytCX
/FgaUbPR1WdMszTaDyW5b9gOmGUOcO5akqg+qoOErA79xL8u9PJ+iyw2k0aR4JxQ
ZztZKcV98oorDvoRjde0NuLQdCufWRsp0PvJJRErwAOyg4yr4TNM0aqXwLb4SLci
`protect END_PROTECTED
