`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAb2FNGHExkITsaESrD64FLMPu2vrQ88A6xdVca+XCxR
FEiLrGLycOqvYn90CBWLc91NwP/imuNw59b4ENpr5V7jcADT+QUsja5tLhspP680
8J5KLpuuWeBcPBtdylBBff1HoYlcLjQw6hLtwEwdnr3hOXNk36031Q/4WNyt6C0s
w3ArkRUoTfiPzlc5v+ZEjg==
`protect END_PROTECTED
