`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44RhMRV2BlLalMF6CIPbrasvFLeZropTVYTIwB89Hd/a
FJ22Uj3IIXq3YYBA4a7JkIWygrx/fXwVuhe3Wx/trVVBe8h2k1m8xY+L39BWD+gy
a28AGe7qQoSrS53Y0SpHzJd+ZRnGJZfZsuQo7NBJo67aoeoxw8Sackv3iimC5YXl
ftESoObe+bnKXJ0ybnE6uKdNT2us/9sAimJ/t9Zx8I2G+cyBu034k8Y65hdxjREs
uRaDJG4sjVNXyVvHRoRVy0DvUaI7vUc1jn95alApR1WYamId6JJUORzWbsCETf0X
cqLDePIjd7LcCEvu/uZhgw==
`protect END_PROTECTED
