`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFWjsnysCHBmgMKf4/vIYbyi3gsn+PO93fmyVK3ZjY5K
9AaoizzS6VJPvh+H8cfIy17eKZVqXaXuVBs5H6eqnWrb0hkFR0bVg4u/y+w2Wf02
iKJWQrqkt38rnM10UeerENLHyumDN1KWv89+Ju5hPwCRv+HQymQtm/2LltcmZ7Hc
CTY6WK9xhF/kWYFd4uExTFfSmhCJ7NiWadVnv8zuLnlbuncHnFJ87GOk6IMGtkr7
`protect END_PROTECTED
