`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/5LXBdnk60Dq7uSvaM4ninTwU4ODsnYMhv93aWShBgy
gvNKIFLvGQQkiSjMSJEFFIzyvX8QRBSkJWdje1EJjmUHxCHMu+eEzvAYfI3Dt68B
3APSvIbpuu4gmubNaT4EyjOvr42gURC06aKtHh5qerwHQTRt4vbjrIX/4w11OgW8
NdUbi4UI3adp9v5oYXTMI/BloA2w4H+Io1DxTE6l+pHkD7l0naSXBdmqLXWS2Yn+
J4bJguMCz+iWbn8LhAE4PJQuc/fx+IgAVMF+JbCOOpptdbWw0DxkfC5cokr//Os3
jYK/aPt2JJqSyv0uVD3UuvU8UYFi1mNGZBA+Jx09etsadlh/lNsxbY5E91lB0+Iv
Q+KCQzujwrFkpXAtZsJT/QNtdecGZs7m5JJTmGCqJ9j5xO1GuCzQ8Q6+EMPD+8DP
WTofWtJCLJMgN0W5Fb7KnAQj0dBp7QcdL1BP42fLBe36VajHRBGpRH010zuRTC2J
LxPGGkxLXts4/fNFiSOCJ3jpC1y9ahN9jQr3inkXtiwfcNSzdY9nBUpsShO4WrDI
vEEMU/SHv47CEFCVzmhzTm9qzeahWKTsAJwUDpjhGIJKpmaKQKxOWyPJJnJIN9Hn
`protect END_PROTECTED
