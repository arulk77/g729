`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
COEjt4J6JtbQ9Ym4tbYeeOggwivaD/1OPvjlwyWLXQXRIBaXZ4Kjpi8JWimnGA4a
HMvY/XHkkexN2QxuAxNVRPYnEl43oNtQnwcDC8sSsse8RuMb4dlZQ+rGBVZ6ffb1
1oX2Q68gGX8fIc6Xz7w7G0d/dYV1e/ZZ05WjtsUrOm/8yVBAGf/WyEsAFzjiSGgn
MNc1Y6B9yRs3vRp/5UlI8aFqzm+GXZsKPxegCA1k8P9vR7qLJAkHvwtGgvnyBYOG
bPaNiEsGjIzQCSki8U5NlGjULR/JqBohLIRK3x9wKbVpsbV9dnbCMC+IO+HAjf2J
3I4XvNDf3IUIGzRdxAReC2o3djv2YwA1ohVDnb+P9a2eylSxEQEt+G7oQsJHab0Z
11NNxRTKjytzK7dKnwNMVUOJXNbNX2qkW/2Qksh5ThPreDos36bUXPofoGfpze2I
xlfKRQavJ1PE5JsJW2iA1V3ZvoLfJ4mIetUDck/JegGsNqPZEebwpbKZo9RkVqHE
ftyjMDo4nGsPAdNb3sXY1zE5lZZ0jxf2ZJdIUH/f7tsi9jQCu+pHWeg0gPcelRco
EOtO86Y3qnr3AuysNFBfKznMMGVSm89dRPWjZ+9OhyZEtoVTR4uoCgg4mclzpQ0M
zN44H715nrx6y0dgps36nmoWRIare+vaZVb3vmul59hECUWfj6U2exgPXdUdruuk
xP3dyeZ+O2yJBUE2qN7v8jPMQ3yEa8hEANLx3QmlCgxFtvQMPAcJheN9tM878KpE
ol6LUnL51nIFYmCImpcEIVmjmSho542bIS8K1Upv+7Q3aC2zY5USu/byY3HcXVyG
ZsOgBHE6m5LWr5KPTjhY9h8xPBXt8aAnNgQ8db6dMeZyVi/ZMv0SgXu0RppeT0J6
rhga9kpIBpYBuTBGblH4cPhQmtUn4PUEuYUJ4jfTwjLqn0zzbKwyVQCmV49Jd2Eh
M0FxnTzEyN0k14HtpYO62pkR2zBNwdUcNWWQA3eHJrZ6cDyQtqEIRGSxcqFDRk6W
JMGfmlcaXCUca9vDqw9Frb+p4zVv9TJQjXKIJaMtLhKKjBYNPeWkGwwenabUlZd1
zglEUZBLjStBcocDR1CAAALck3fjOUnA4ZOqp7cdQrBSg7hoqLFznd4a8sWXMlcB
pBjhPQNGm92PPuKKJpAUnDl2yLrYIhdmogxM7plmaDIMPHRUaQhYQWxj3oZqMHfe
jvqDq0+0xh+Oudm/qk8oc30wbobB4WhXJiMHOZGrPjUpukOlDQjLA4vKS8xkdMNf
OhtfCrwItlTOGxUHFvt5gKpudwuuIEduoP521UVRZV4fm4d0vICmY19X1XTvOg+V
Gy1U1KkWyNoQydNxOG6G1M5xrKrku+E4YW3i2rMO2YEwU4RikquApr8RncY3Fjwd
+5decB1tN3/UhOu4MW4LCUP9SddFRWRBMVcK+7/1WOkpDn9mw0vFoDdyr55pprVb
X3gMXczCwM4c8T4BnS11J/N2Fxun0PRjWdCMaI7pba5C5u5gvNBrTmW4fEBkcPTy
Wy6kXfqPjybweO/XPz8aCWNdzWCXjjYEUbfBcJChOblnvlJJCeQrERuiJYulFybD
vp+HOP36Gx64k21HqP4ebqm7nE0a2lOKAjrSsPRlUezs9KFHu/Z4ebUxmmM7NHGJ
INeZoF18iZl8SVts8e+srTdj6fytauI0lvNcuMVImygIbqaBg95b5b1Iqu14aYxl
HGnVp9bqJI8/A9u/kJjfgee3Ckz+Tl4F81N+Fmxobx9DiGQnBvph+NRqVyxNRjwX
nRilnNEyxe55cq8uDS2AEV52TiePaePPd1ktuAUyYUKGKHPjBh9HXQZiYnQbwUcM
nO/Wnx2VN2Ms9jjRZ8Qi3uLXCC1KkxwljBDLQPvx6rAz9hFgvfpPPLBMf5sI1mKn
roG/BEnUKmGIG+CLNWGLJLlzeVTFEoRKyucxqGK7AiCIEsutoP3DYDbMq0Ub1vvZ
fdfz/xySaNOEmLXVNYZW7oJ4oB+HWX6oV4wNPgnDU/UcEv1fAkwOwfRqJa426mPp
9M0HeRIvkkOYUXueVDWcqKzs+eXtUoQZOCEqMv9IIg1YV1qDTUAIRMgvibC8qiDF
SBuFlInNIO2ia2EA4x56uDfRsCrXx3ocuAzSjz1cRsbOtQ4vLFD/tDPdLmRjszcY
7Ey/9CDsLsYZTTvzCbFmWYsOSPbgostnJBBY83pJSaLKsFXIiaggthpkyT1H0x4w
iPa5Ic9baK6rYgx43IVEiKl2lKt0J3jAJgtoCyvDPiAoblgysAR1hS1eOrB6Pkho
TNe2LDjaaxpfJ03D9PXa5LMUUFfEUWMcUCk1vFGGzNrHw7a5rH+FGbC7e9gNy217
Bpn3UdVQhE9LOwvzJezaKRi4/p2FvgE5Oti5gcibAyYYqK6ZVC0Jd3xbHIUTHbZD
7DshkuTSp7vXWMjXtEdEgOp3f0xzU2I5T/f6evonBswsDyThWo18gyyXHnxrcgFo
5dKM9HSkj4sOFlxfCBjlpFrRpAhwtA5UitpYH/nuBjwLorn3OQ2gIp/8nQgTbjt9
PyXFJC5mh36lZ1pHlxxzfr/OKDEbt56W92zEMnS0CvOnRXS78RDQCxp77TyIkInb
Bo9XkeEHKTTD0VukNzuyCCJ6+t2pQOMcXiKe5eCcOLG/EGdoIkV1UtWaU949KKAk
MsYu4NayVRow1uxviEV79c0vZGrKl7/0rygbpLYL6DMpDlcNP4IGO5ITomOE3ipe
0dItC1JQxa0X1zUDLi86/AGS0P1b+eyoOwHzmrEK/SUbsYawJHBma9yC48igd+AY
sYv8tQG6TbzpTeeXZ7Y5evCY/HHpmgYD1fVyccnm5ZzQR17jce2p9ibd64jsmckV
/aPVRFW3PF2GJzj1QgtRsQz0wNof9pVcZMZkQWXJxNG1mPmRK33GLMODGShjFZCE
wbGwwTj3AY7l3REGCAtPFWg/MVzqreFQZ3dqvt0hlFt5ZBVTAUtwXlumlYkw0j0w
63TW5Bl87yJ78Zcqk8ISCpw9MchcyqnbA5WCCyyqjc+tZaOUbiHe3ujENESevRw/
L22ShVd4aezQP0AEi47oxImGVidYIUCVP6XWguRnqiyDl14JTO8zhfemCDYYzM0o
iyJTNDixmIIfbZKsCu2V+Wf3TpH2o4rB8GEsCyApMmJOS0cyufQ1Haqnck1PqGtd
Sfk6kSxQKD/FKOeRZuP2leUAOYqSh8u182n69LOnLWfH5veiZlbuG2ISureqMM+1
c3uU6GKmKb7eJ84jy9qrQKJhXBtjZtRarAxy1li/kL5hFyJgFLdoYt8NZ8HuvyeR
qhUCXY091KmR8f1zfhXjDFwFEch537/vH8uascDTMRkUstnEZlfDtb2mWhKofqdp
m+UUf1Ak7VjlIPk64GfdrUCMWTI/8Mzcnzd6A+Cfbzi7wui7UHmBeWjDeiztygld
cYQ9jbc4SgOZTXkf5ytVKNxm9XsozvMYg2nBwp8CgRaIf/3fKYKLA4cMFWDdWAno
ARrWjqRTfqXd/rgEKzS5hfCD0CEB2lgrgjmm4EcBxCUEvaS09J/mjywadnNTaEnL
jCRn6glGnhdafNymSvRs3Gch/SZYGmq1rFr2haKkgkJrj9xNV/IZMr1ljsM0Ai1A
y4s/vB8xLpkXdgcaFsCO2z3mkghPaJYZsqn1lzF6h2bEqD+82buVnifcdNsYUS2Z
jl0WVWErUG1jN7v+GLLi5+rTq5I23xNI+e94n+IlYmbho53vTGgS4+HrQ7kekpBn
hprto6Pz1ylq52UIioaD95n3D082xcPibJ4v0snLm4LNTkAlbEj8UBUF2zTHJtSc
hAPz0fWxJ6ZosgKoceI5issodPEPUGliIuJ/b0Tj6BbWtBwZ0iEBiVKQLtT/uubQ
e3p6ppFpuvsr6QGuspfLWSRspzdENStA7IRFeXipxs+OVjrTHd1LnGXPK5CJLhGs
hJSusfyBMZLLH3NRzODPErd+wAFiKk9CMz20YaEhaMUCj0lYK5tjrCG4dwMqaVVl
r4ylh2sNFeGPUacdqNyStYfMH8X+A+wQmW21jHhacU9IACdyzV9puXrRKcg2KqoC
Oais13rmWjallqEvi7BF3yCZL99vhiYfMrgQSurjgpgmSqu6y7ZeahSW5lPWub+g
NeLEaddLoU1B1bYpoqss1R/WQcUd4uAm1F8n6h/czixq6thVS4lpogQkLRB1wrxu
pmYB8VoO//WS+Yd3GkGpRDi1VYv0MOye6YbQJhhDuOmJVKRSy20hY05VEgnMaOTa
uXt2zT5USn4fS5yD7/dOPmaINTDy++YiwV6iMn/0osJ3033TBwAl1+XmGlvXDjv6
TWdlcNhGk/FzYFGfhPH/x3wAe0qZUtJOw04bgIflTlQ8G1qmOvycoxzNAL/Pg7Mc
9vlwDeqV3p3pbIX/x8SP9PND2arQH+THIvYaeSE8Y1H579Q6eao1M6FVafS1mfMb
/A4NORvrYQmXfsYBsIfO1hhc4wJcVQfbF8H00iVVyzHXAE3d/v4CAFUF+2G+6KK8
sgbZonarZnV6MVgMH8n3fiE9xAbaxGxqsGKBYRwrxj4zcoKOOAtG1PoEupP0Xeh2
OYIocZY8mUbdlHeSeCY8RPBP6IXWhWHKwbnQmn9Mh9nZwbH2GsmKgBogmG0IU6Vq
FJEOaJROY6WeEurdgaFHL+ZJUKeHT9/YOffgyJEAB+pTvVjonaeLGzkAKxbmtN9r
b4xDm0lwQKBUV/R5TNdkCSSLUl5sfGkj3xpo6215+Ob4WmknU1IUVw+3xjZphZNj
Ar8RFMohQWo8R6sY1hJp5Rl1nNKFGdcFA7d5puO/Olkkc2PEgD868uPbSJuaF2gd
PQIJNkgG2LvwRAQaafG21yjhmCnsTnB5TT0hTz6GCPA98sBhf/yEx/bbFCdx4rIe
t4HMSWwawhEXLmbwHWz55VlBEHignZjcTRRFYhB64UfBAdkOTJc6nSYAlPYZKs7N
XqTxbl+i+u6ZDHxl0Xp+UWfacm2EJLw4ByLK4LNR5+XWVqLDGaEHEXp1UIQmmGno
en2pIrxEk6DyIQey0repl0LXIMZjyJhDVrdI6BZ7X4cRz7S1NQCPQcCTl6HIq+DS
0vm8a7eJgpqX3DhC7arG4ybBqDqMh7gR3wRIF8MKp32ZtKq6RGqzb6aGx82Btbqr
WHr4q0lJg7jKJ0gszrTAfYApkif0lGpEC4XIZmZqhXDgQxruJICK4QPmvQb6/Oxo
NlJH0QjGkbT5avNK9Y8qwiN7NN4rEY2pmcmYP9tcVhgs7R0HxBmHSjcsvCElgqqp
xNLzLDMntbJT6xeIoeiu9LTtR/NC7Ae7GaQwRs3YxZ9SUWQrIprSDFrI6yhJjBCL
59DQwVA4S4hrzG+qnMCTnvU1PsdsEhiXbXJiv6qHXxYBGhGI/zw45M1W8uMEOHtb
tppE1TCI+n2rX96R88IUh6eyOTEGS91nRUEQBrXFZNxH+HAc8jnl91dDu8lynCXo
6o9+CCz0TORpJjKPGvFEwb4ghPzvz7TSFiJd8QIxMylZDrUntY63Him1FP1KQr37
fDM82O7s498CNTGR4WU6+kefGntm76uruYoK1/JxDnHZ4HflYXyy8wUR0QLgNfg8
iFL8FX+KelK8BCNPXFgPHYokvdcmzN2XDs5+UIn+s37xeq0ZcWzYnV6gKjnWWJGu
kM0z2H6el2alxWg1gSCsw28E8keKdfPgEJSGOiLAI4fxifndz0NWIDTKGo4b8FYu
1L3El+B1BzGaMoj8wUmc6tr+DdxEihFuYFUXlSMGUBDLB6v444lg6oNcMu2HzpiJ
5uCOHLpYkcXY/zfHegOpWywrCQznsKpiFlDr5a/YnwyJs0uJj0h7uQn58sLc8hZk
3gQk6KNqUXxj9fgEuBFDT83xZ5AGFe6FLTXHs4hiL69NDtFW29MDk1NAGeDeSYgK
DGcLr75uF2HWnV3qQ+u/EHLoRzRuLHTr+BndmLarwSEkFyIwL01WBT3XOTQKz/Fe
X0W8M7wP7jUUlV0DHUA6a5AJKSO3z9eRzZoLq5VO2AZmaJEt2fkYC5grP5uSfYGy
Kxzorntdsc5hC4eXs38zkDK9MFcBlWcT/e78R+JOyaSbynXATPjGUqUNLkNVphYM
PfKm/Tyj5ZvcGl0zMBks+De3yyAknxRv7br5zXhUTJGrzJ3Lra6gNs6bfEJwgnfA
MA+T6epy7kOjVMIxmvIyYYRkKOdZJZqDI6zmOEjgqFohPu/OkXm/hsOcR3mW0HyA
nqeNvCgbtnwCUKTXWOdJqHrW5Xo92jdbSdO1mo3dzULDhyDcWFrLgV1FNz2pLWMw
X04s47rAkA2GqTBXyQb8DhCCjYO+yev3iNM3VT1FD8iX5jnFIzG146CyK5Jekqfo
OARJkNmCeVjjAu3EypFpG5K/acQBQvC2WQqBBIMiitvtTNUXKxNLiNhUg9WLSr5y
WUBVegqPJeyN1iZxQAdt3pxXjPo4Negm5Y1Fplv9i8AC+/zvp1xCF+rUnfSdIKS3
HijHdaa6gajaM9OGRO7CY9CraWl2LCv4tOozwyxAIgTM3qJc7OD0bsdoJWWloUwV
DOvMW/vSKi+c2Ew+We+4G7a9zFANPd/SWG8jEdEAqYpEE4XKDQXLU3Qmwcj0bvrl
ekXnu/caKU03Z2NF85NF6gMpU4EgDzJ+VOfpKJyAJHzzom6C4XmvQ+KOxtbD9/MH
bPpe2Kyl+/rb6ZRsSoaetQ0gVE2pVmGoAlOru71v47TmRcCkFcpmElc16SMNAnve
4SVMquKzk6c8VwVl2XIllVWJI7XsEovRdwh0jj+Prs1dhnd6nMG8AvdxEguT0yyc
HkRULL/yp5z6W3s/QkikMS5iomAJGtj2mhwMsEHkhOetwtSbZ7PfxWqtnPEl0Sqx
D5v37c1CV7XlWeJPceZuFi+at3RfDqVcTQN8pq8on7RVYzERns9zbEqnWN9yGFU1
SNMen7Rl/EsLM/YIsp2hLIE3N7/KRpgrVuAWorXcuWssanjRzL5gs6/XgeDkei49
6Uul3rLzyWaiflzEfUEwkgrWl87cJnR67bpWkSA+hVvEqX+AhjTk2q3rRV/YohBM
yozGqjA+c3cox0rN+jmWk5gNDp9F1WdxL+0rcueNiFpDfFcJuVOR49M3Q3Cfmema
6wbmeIiGri7V/Hrm/mW4aoYLmrJG8Jp5iOaIvbA6cNSiZLLrT1XLa/BZCjody4x4
UukCs4BFVRs+LVk3BCaIQN+NPfUNG4aHBfPmxYgiBV1ycNvXXE71+KkAWWX54mWa
eY90YMH9QDWso+t97I3aifwX95vDtLfvX9gsWV7d9aTGKQEffK+EtWBjqfXDz8Qe
UsFzVtFb4fxbUVNca1sSatCsUyM7/ZNKwHTalnMjL5cHwOJRXB+B6t8VwO+0Sbcm
26dBMwZKIwpLunX0yqungXyAEsr7Cb/un0MHYgq8nkZ53gqs1+JiYngWD8Sn0MRs
YxxsWmidbgw4qRmPtzwNozKlC4Qc9g/Z+0nO28qZTialsBWrQWQrzI+znExK8Yff
h08zFXLdP95S98yF8srAVofZSpiLPOlrgf0cqAWOs6OmqiJKHIyMMoMxiEKr4vu8
ZE9xHbhRgwh0hXXSAwxlsY0jSl/ArcAJvcppb/nJ0ZqPujT3wIla0uGLO5/0EJck
OeToo1rca7xuMU0rF0ja4Wybp/8TApvXbxLYa/pwzX+/6CmEiSgrp9pv+ZAc65Bn
SZ6cb/qYCSStwegKH2/DZhDaZJxHzvZCizewMNMaBZhrNAEA0JEgsMWeGgpfyKpY
F69RoKP2Y/UBfz6xNz74Vl/zxpEoyudUWAJNZfapIDTChBE6g2jI9LFGzZf1S+bc
WqQY0supDC2XQNm4qMSDNC8hKiSHZFlgvkxXVG8sAmONuoFnm1ipJi4VZTEHEbXR
pQEWl6rzUZsUmF2/35sGWdYfV924c4EOTS1/nimXOmfZyhiX24abW/65czTRyfnY
knnqk3LfQ4o2HE79YqJ6SaY7v2Fk5ZRnCXZwbF0vxGrsnss7Q1fLt94nP/SFLPml
KnvS9O9FAlwfUZOteRiOy+mw254+q48W9MRRl0RW/izI5d/zJp8ynCaHnKJdHAiN
buIfUOjwibNE06qOFvBEE9jayYH19tkpS55HRgD7pQjP2lyTJcoSZuITNVrqp7Mf
TU/PNOQovn3F8HF9YR3jZTgf8v/p4RwdJtZS8k+Z+BPXcZhO8u+WaWqIdCXW/NXD
gUAu8VtXdr3qMoCKkXCZywREsvlKx+hovdguTtdRGFDnuwD4oTRLlKDkXJqs97OP
zp/j3B370ZJr+lsTF4HsN26uAgMOM5U1mCvaxAF4oezIDlunF0Gc9KY2MWJgzF1Q
70xuJU2fs4AKnhclm+5S/my4vtrLEFenh3EA5kMe/CW43CXotQ6fJgnKIpyn8E4m
/evWjBM9IXbsHClFAjkxV5Z+00odxBVezU8vR97mREggMIQrjh/j9F8OYn2EMA/0
bvtUcgA88poF0H+lOMOZ3vHinfAnucYg2RzMUqY9vsF3GOeKo6676HrXbsyBo2wl
xDifssnNID9yXFTkb+r5BJlC9+syirwVmaq2PYJLbXLjy3J+vOtktTKTk2+OHlDr
E8qb7HCO/0fSWSahLoGjRnFOglMbdcSWMvzWUhvDpgPYjIVFhnypYZh2XmQ5dHlw
rVh4e/IwSynGCj8CizSxNQLpgptgr6z4eytsi9pHKsVZoN8AP0yxTMkzmOCj9xpU
1yoEIJlashO6oA+aYtUlI0xpXoavxXzDre4DA4UM6sm78vqrQQp5WNUsOtJg8/EB
Wt6CBNoxlU4TJ5XhqM+iAAEHsrr5MYHIlth+fAb8/3V8X/PkDEG6u2ET9nBeIutq
vx61gNsQ+KpCAfj2EIzcp3v9asn/jTAA9KawKBB2lGX7o/0HOsjTI+C6fk2STFjh
7kEYW3zrxGzmV9OPLhollMdVkX1p7CbuQ2JV8nfTqUin6nekGN1rusE2x0Dp1k8Z
epc0ZjMxqTofHwt3mdkKykaHqvqZiORubzHGGa1veHsxYCL7tCwk3gYy2glYRb/s
nx2xwqSXOTd/09dX6Z0BZLqwVD99GUmulYnMi7LKpVmiK4oQPetLemWM8Vml6Rps
h/IUbZWkWXtmhIDyr7xJcWyvLlwHoC5tu8NBhzJCh/DzVFKRFy+5SxQGnBF03RtL
dGj7FRLX1MRLFIDFbDBZSSzLbOAFol4difY37toc3gThCfbE3/Bl19NyZ1REtpiE
toVR5lFaN5WjqRLvUfcBi/15pityop9pG9jqcEI97QEiXG5kYkYUyK6fjkaHBuQ/
LvlIgk/HUNhYcRLSWbaYKD2r2GiOCarAvbvy4MKt5vAglEWG9fE3fiNJ/1OqToZU
JZEbwGE1MEm0+y5TmscoeYDVPOg7e1yXMFdf38A9EZqYx2andd5AleaD5P4i7lH1
re78tbSiOa9yPaIX6bT3YUY7iDJu7BDCWJPtHGPubYnfD/HEpUOqf9EoRfnYVEk0
yKEDa3w067VJFpAQyPVq481TsL/Q0a9Mqw+ZELnJ70w0OFUtkZ/uH2rmsJyK7tEv
opDmjOnXNLYycQfOSHwpHaa6pI/Qj/KvkTvzq8Uzc8Kja92ls57+GsQ5jdjEzAfi
YxzIkcy981+tRg6is47x1L3JW7xlBo3vGpA+UKau0v4qi7qGwSlSi39qR4zzT+mP
ykbOiM6NamgBEauvJMsB4WRQDIfPS0fEi2dhhmXd1gHu6JllhAMhYXGNBH6EYWAi
/NrirwTc7qVJ/ejOdZ91G9YpaencYjprlut9nlZtA8XGsyRSzC9YUDhPjv5f0Ygc
LmmqSpwNTHOc16pushJ2jNrUPBSc8BNeoj41KZ08r1eqQ9xS9a5bHuZTx3YvobS8
GgmTQbE07L9JtHggtT+3wxq0Io+zI1bccgIq7k3tBqNG/xAxUk3OmNVTlJ8f4ZOJ
e7oeYeWDk7pfjVQzVj0KiCz2ibjgHgCNLne71ArdRpeN3nK+ZjD+829ki+4zLsO3
ZmywFNuIkGr8OMYG9q0wm3vgoJ9qR9EoQ4jf9e8lCZ4rDzQiasP+Uxe4SAjoFtAW
+rmWUAzHFX/yooJYge6Gkq63SYffmjViQeywdFDdBRQloBoshMOWCQ3EeY6VrgmQ
F0DsOCwjP8miypaxu7tO1tXwX09AoVMPrvIcHPg0I5h+P9C3yGNq/ecJrUjPhHFK
Z0tDtmaoOvJG08W9+gGy3Ea3MkyEIjGZ6UYKX2px9Z8JeAajhzWLnY0D29kvyAw7
/TH198m/SjOdT5K59Ghbm4BYLHJszMWnCX+VKTfPrlKIwa2q2YxCUmvq9puUqBT/
2u+MFKPdQl1ul5lbfW67m5S1NoHsu0NpaH2pZ8+pVhT8MpnKzsvc5JoiXF6uxtav
RoXJ2sgXuDP5yuMV3nz1FbyBm2OsitbvJIGuB0gLWj7uBrXwCuKY6f1BhTlkhKEJ
QEe75YbdlfZXAGRKEFf2OzswXBNzSK/8S5JPTdkA9WBmgjghNqIpPX+80LTPsG8x
LbotiorFsUI5pM3BIHZj35cD8t+IzRtF4FnuzdXp245a8wMIpR7lzhAM5yzTiq9Y
ICHSBlt6E7u9Sz3uzKy93XbpVzkX1NLlrdxqL4clwe8u1GsB8b7BEiLZzbG6nY3R
2PDPSlM4X3io6C4yTegkf/W+g+1tuF+yHaEOsjQIXM+kCgKr3WQj/KiNgo6WKN5O
eyW/I6e0QY93R4kB/4VlaSTKBWcLlYb5Mm03SeSwj5uQPyJ6rV2k474OC9H4tCQH
ACh85nMf/RJCITGHbaN82FRvnZicIJdpXHjbivzt2ji1Mw7U3508cxvL6MXN3ptY
WG3/TBkTVMzfeuD+6SIBsb+GHD4SOvqSTdyvY/vJRm1VQUOhs2AvwBhmwFTFQbKI
U4DYh6i2BpyHOospF1wpDZ1Y5HAGDybFhIi1IJVcT9OHRCKvpIiE09n0Gbu9UX6i
rzV7T0SyTiqEutuxkU/SZkkmSlAZAIFQnFCvo0RIivkC7d23Yg6ZCHuHqkLSXqym
pFctMRM21zsijDzoCPMHb15tUdb+vD/Ivfhqi/rCJvFcCk2FOkY+VEFGpa6wN+M/
Yzzi6WKhM76IL05Pz3YXUH3y9OejyxrhVUDrrD0zdedi/PrBHhA/nZn85MAtEWux
UNA0XeNhvCr+11a0FX7RPW+e6sUVnmeco0GyyLI/LJ+Qv0x+cditRK7oWK/VqFCM
mAUy1Ex758tTEnjb2dNoWaQifPh4MeKiEHM4cAdLLs3Agi+xIOpzy4HoryS/M0lv
4bZ7bsu6Oq53ECrdDRrpm32TG27pm6FSWeCH7G3KBtC0AcmEZBiyM+Np8kI0YRfc
eXIDO7d09j0owlYB577x4GxKrbCEir+uagGHNrArHENl8v+vx0p0GekwnPOXWhg/
Gi29uqSyvQrd+tMC2wMCkl/wJu8mhEM3ynHNjdwgGKAtVkPN+RIMxqEL8sakNQ3w
X39h0GJtABXL72WBQMj849HwqP5xsHRiie/DMnNxU2x7Y/OI0GZjOaScMZQUtPxE
lEgcyFtfHt/Acc2dby+sG8ITbBGd0yRXiFc7wpdj3724N0GjDC/87efyW3ObTzM0
`protect END_PROTECTED
