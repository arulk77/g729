`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDTs4brU11Zqx6RwP7Z0hc8X00YexHJO0/G50vU8F53A
CHqQYq+yrlmvsuEvbgoJaWTkl0lCb1RiRpiImQbJAwyQzXRJSVkSdhSUJ71UXBYn
aGJf+lTsPQ4/H46xhOXywI45eQvsbcXLXZzGEuWn6yrGciWu51pqw/wyBciD84/Q
Fqkm3OfeEUheT9NXTgk/gYb5c0NskGEm37UhteFoczqScgnjWlaAZTeAncWMhDX6
`protect END_PROTECTED
