`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKqZiyitniBQekf+a+zS5EduoqGVknhawxSvYrlQz7IR
4bh0GziuFCW8XB/ibQv5zIfGTg6XaiaqMA511aNSKWEZuuVw0UTlNxGsZ78YEH2I
FNATEmGHc2jjL6shT3ermR8eeOQdA2r4nGHG4dO5/DrKVdz+lPgWxXAh6c5r6wLi
Yyn7caesuMjSFUo1HIOBAaj27ULZ0HXRc39uA1KWOj0EI3oiQomFH60jRPH9+DKB
NXYeJTvtizQKiGCucRIK+/jsPLKfFEVyZV87FBhTb8CcS3/PK8h1U0EAi3M2qgZf
0vnL2zDQPTuOrkIlXk5yPeEEBJn2EvgiIOBQSgIe6J1iWPiLcoE4bVVT7sLES6pS
7psrgC/B9E7JjKU89aFY5M/+EIOTqgCFmGjNdS9gIgj8THu4eQPm7peZ4kndaJKn
FLsLkYOam57bV2R5Ph+ZDZqQ7Kn6iwGUQN0PwX+zWh4QYA7ytFLmCGxt3z7F96ij
yFhGRipL9KBAvCxM3fQZyQGurkBYnazwKhBbp9no87ADrCGSR/+J1pubh3BY3R+3
dZMJyZzcM6aU37hS6outFUpMCoFf/N3b9+0++DthbEqEEm1QL8wSTlj/U0sYsdc7
`protect END_PROTECTED
