`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIQJcY0rOdZPmmxeMcB1tAW6jgaztlvuT9WcaG2B0dJE
x73VmFKrfYgYf6HpzZBdhubEECOCQ+a+/bP21fY7cNr/NZPC6F+c5X4Xb3P8Jm12
DLFczW1CkWHi3ah4tdZ4a4hQDtT4k6Rm5Q2Q2Mva7tJjtt6P94558GYQeqAqSfPS
OseVMZxytnJapcOM+m17Q7qtSBWSrb4919IgRqP+D/qtaL0+BQCZzDmi3rPsrHiB
8l6dhiPCh65Dg1lrNRwaLS9aUgQYYNkNRnCRmWIwO2lw9Fhi8Qpck0H44rSV5X0W
BbWplUpe0EI/+pAt2diwfqUp/H9uNUoz/iOjLHQiT+QnagdSSinVphsypAJyxeul
`protect END_PROTECTED
