`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45qyd60MJtrBb4exetwTZEabLWSf9+yb75QRcV0mDrfd
lMHYkX9ttKUPw83MXwKq41O/R/w5Zve4qEar2TwrsatPgSOn8bn7JSnRBL4IrrFA
v71xjgp6i6skT1pkxEjT9OYNQvtYQzJZW9grs9LAN/29ms+Ds8hLz23LS+O+rJIU
FJKmyXu923N8njn8nIwX07atEUXJhnCegg1VgzZnw/ltO+F0Z9lI1oyx3K4dVsgG
7/Lxn6mzVhKr2sCVHM/pbP7lvfUChdqZ0o9QAw6iTCY4cjuxfpJFziSM4u7EUM1G
9LLXAs+9HEcbY052i4ca18Fs9xDKnR/V0Nrahp2j2MQaLtuTJRkcLcTnJpbCz5Xu
mDBj8Klkwc4srBcY3j4ZCg==
`protect END_PROTECTED
