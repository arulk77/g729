`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu444tHTWPXvBZRzn8eAwQ3KDhNRDGrAxA1ovfUfZK0uAt
sDYb+R90QibuUAUDHsu45Rb7GVsfCe8pqWGWOPwGrDaMrT7l05eircXMhEPjgUPE
gs2FNwciClNbsQknsd2pXZp8FGXMVqLBKW3q2aendCUFjX7HYBzDNjJxfaoMHaHg
uLJIEMMsS4XAGBJ5OfnkefkM679m+MOAcvy8FI3spOjOKz+EXmtAAP1INBtr+KBP
FwPP5ZMnYR84YKAqksTMFbqQf0aU/Tx3DgD5ZhP0CR/k1/GvqwPMVfXWQLm7ihQY
/SBM/H4hM5dvxCAYLV3EI6b/nlAlmlYmMCh7wlCL602wUCjBCEz1ITJmXAdgWA/U
wmzY44GlmmoHBxSzuZTBbA==
`protect END_PROTECTED
