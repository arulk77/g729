`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
BpcQZjPbz7GrN4Df/7wuTrzhHrgu79v0Bz5IGj8pzmRShSEJMwqavWs4FIsm2P1C
uOJd02PmI4Mh9UqQdqJozhgYYqBbwCcrTN3KfbGHOB3JqxngImbCynpjp8hG6P98
O9wXeUEA0PNhSALdXIOfkUOhJ1cTG/RG9OqQ9izWW5ERd0J73ETfDCfF1dSfQBF2
3avH/VNogR1Y33crNyFUct7weYf9B66i8avUySaT1cFI3bzXCB14qHT5d4Z7YhFa
37vAkgu6bjWd3B9TOptnojjRKbyJ2hbh1E/0uOBCfptNkReb3wjjlxR/fuGBS0Mb
odWZvFNkyInWthtgYLO5mQblE9XOVN0FowXJs/CKkWWiRET/GPKaKSVw4Vf1AEmu
2DBwE/tEZJCzK1ewtPd+IZxfMZQKcRJzAbZ8OWrsHVQ=
`protect END_PROTECTED
