`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePla6NOnO/kbb1oFDwwSxPCvwVt6vABGVeGLdR53Oa4V
E0WnezC+Dcwde7sUlos+4mZ6Vu8+ayL2Qd7oOtAI/9Sb0/ls8cEmNDvYTdv4a7Mc
QmYcvoPOtRB9Es9QN2/SJTk01kLdzv0nyulvaXSuVdd+SXJuPncgVXQVdpPfu7n7
kLYIuZLKQ782bNKhfPuG4QcXm8O9zG9B+fFaeD5d3zBdYEtbcm+PLS2JLgxH2GP1
XVcDu8c/MkvMBhpKdzYHtFfcdE7sFtItoMZd7S0sKjkG1yvDNxKmrceQv8LfJDlc
fQ/aRfWSvXoJC1IVLhrKA/tT8/ScmdbPpwePdjgk5Dd/D1IPh4LWuevhwKtVy+DE
Wwn3walATHVpkk8rZ6VBj6LbMWhExCQCmggQ/4EBG9vk8zOLTue1ZpNmiA2hN57i
7/d7fPs9uEtyJmlJ/+JewvehlKE4EETBSNYlVIzKAk1cm8skdfibLW6eTl3asbbj
2fLa1cJyLhH82Cy+hcwKzQYuqM7pgpHwFtTml92qJAFUnPQkEVJ/gkArvhKVC7SW
`protect END_PROTECTED
