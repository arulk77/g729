`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFOXJSvEbS8LAWK0mkPMrW/DKVwU+kfTAvv1g4X+buQa
y6brzM+4KqzAQz4lzDCzh0LK59ayrJP7ChXQzcNObJ3qRTazCbr10K4+Zx05lUCA
A1G8xAdKqpJS6io7uRIt+T4il6qpq187Z5tUejQj3u5DfZ4FWhBpAUQzlrlYsg4S
L697+82vFV+qP2mMFwETzrM1yLg1XYpYEWonMn6r+JG6GjI3G+7rxFSwhZakw6x8
EiOykQITqaDIMBNZ5DEkUA92rASdCK1ULz71JfDOKAb2Za6Z8yvhSQASCmSmuFFa
ocDvFpxVZne86wXefRMFMUtEdctgi62FaM3In8mfVviWIl/NlqZVYPbB3iqNnOEL
Zx/RkTvCfxGikcKG0tEE1BVYQs+pJJ5kfusDgqqdQLS6W9VT6mlTJqtVd9b9Iv3a
BcpZpDqo97B3JTbfXKj5G+fRjMOrOBbX1OwCGFGYPqQFHZ4ozNcvyg2wOFxJDI7c
Kx0sHzgtgFPfmgv1x9IesV5/lZEEvkkFL7IWhc1uT2I5Qdko+ghdoozvRKfFoHm9
XC0Ou1sZOpGADxcAA66YoYv6muNiVU+TX9xOcSSOQT8Q44y3/b2txkOM5t6A1FEt
GFkKam6gLaytTaE+Rv3yg/05lhB/CKQzrnQEY6xq4nm2x3UrIQRud5zukUOwdpX7
`protect END_PROTECTED
