`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4z5F3I5iPPw0oFQYpIFc6gJqqa24HefJHA07M1GQPmpG
Ew9AUSkgQl6AV4nRXOyyN8fbWhcGLf+pT2dEFkBFJjV2djyrHQsBOm/3Sn+jvKWZ
C2xggeMWl2DUagTGrdYAaG8FlWZbtjaVNQL9Q84wfteMFxXAa0h5suEfezmUW/fQ
HfQrsLUnW8G2VLxlUCxvVCe0DnyfhlwTvclZG8aPAVrHt8yS8hSV5VK7f6bSZTLH
2ezAPR1Xj59YBD24RSKp5JgCefKIn4/Rq80joGEdPfWKwY6mzp7NH+/NVBJTcsGi
W1Flfo41ZCbVJqtqa/WeVIiqjFyazzuKEAD2mW4xafNwprCnnJsblI41FPZMExpZ
9XDozSFZmINa73+7GXa+pll/g3f6vERD3BLIBVf1PAkjSSRWd+my7br7fIB4A/TJ
s+zdAslbIM+NsGTL6xt71Q==
`protect END_PROTECTED
