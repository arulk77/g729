`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP/66y/WWuc8J5NmE+cYi1bnKlaPDFe8HctoFzsy9rDz
HSaZWzLRJrB0E8MvQeFP/gCnwKQTFRHERXlHf9ribMwI1BgdXBvNyqBKiI5Afy79
BKUy4raYY0WsLGZs0RNcPtbIy9cpI+ZVFhCXGA8OovaZXu0RcCfNP5lC82Nnqyoa
dR5oJRy4xvgeWPbR2IdiZQ==
`protect END_PROTECTED
