`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCwumoNBMh5z9fqbyve6aaHuVOyvNKUprZOcFLZ8h2Qc
UCASR3M6X9NDHQz8AlUxQ9zwYn235whUMKJwWy3DXyrQSLbzqcB4DYReJE79qcs4
K+INa2C8V8OozSfiCljukoORlvv6blDLbKO1XGhTvNgIK6I0SqweC8epymDmr/qg
3SQGuMz2/1GbOrh/uNVKyZkpMXV4aDPbdILc4T0OM+ZHooRLwLpIJdvnTPVE3zYK
JNbNIeS051Ypc0TaIc9L0OCNMUC9FpUJDlEwNGlEhu8Vd/mSwLDsfygqo9N4EAFY
KVb6jWmS6I/8SViKPeg59w6vf+MUje2uE2LyNg9UOq1/T6Ke+4bjHWDrdhsCPT7L
2RxCbXZUvP8qFKzfU1tgfwcoFjKfK2EnRW4po1Mx6EoEKeKTdDk5ZHZupSmxYTdB
mEpGLyQkSPAZWgumc8D2yG/eNTKg4hdQ5+1MLzkFAK92Hf96/9u1jV7pEgFDmAiI
CBFRu+OaQsC26q+NgGeSR08v+mRxymol/mIVsfXPKIvFBgWLXhm3Jpchm8pgXWit
`protect END_PROTECTED
