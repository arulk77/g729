`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
wX+z6W6KU+6ZnDmzndevQHKPIwbR09nci/2CWC4Vg6EUdcaua8KagTZEvWIs6eNn
pnAEiF1mTqB4XA//O5XTbwZhArOxQg32bz4277cRFq3s/hvuaUCllE5NtiBCxj76
ldE2dROD8Q3+hKsi41cE+GnXELS8htGwBXwRZb/aRgZJgnWPs17kp7eGuYE4ZXTZ
nWHLTq9uKabtHtellBvAo8RIbPaTlFh1Iu6tZus1vXgzrd0lpyMOc9xt26Jlnbh7
ohM+xyqaru6J1sDIsgDbeuUhv/MbVG1xbgtHIGmUO88KmmGg2H8MsRKl1hq5TOLu
LceHwn3LRrYF0CaFeX26PookhOYfVRbKHu9Fv3YEcaZC88+ipJTpUygSSqExEhbc
OCIKdkrPJ9kNiyO51fpzAX0QQZrHa5/Oj+pjdQbrNHT1wZRW3288CUTOxZZ7UN1P
cS/noX1cjuWHfZVbnrViD8WI7H7iDB0k1Obfgiz6hRdONYA3qEpN9JLKSxAwCaQz
soyt+7rwkrYY3uMsBTH7QEKulLIi1kcfN6gAWt+U0m8k4tQdOIfsnVimRvZyD1bM
XyLvynKjwRdLjpZsKHD3aNj8LwqIIu+5WuxG1xry+pQQYm6uKJP+ZYsSjHH2lbSo
mMVil3NAdH44XEJAOkOJeTZhPVCpNvLUcFQVIUB3Cl0X7rWjoXt48OsBupJFptz7
WcpZZcsO2pMrwEa+IhaAHHXeDTX2eOWTQ9n9HY4+QIDGQsmucUD/zkaW2l7LgVbp
9Ief3yhmFtGevl/OFK3Gx2EJuNuDreerg0pC01U4ijsChKv5kBPeRcfY51uq5UMj
PMdDoIZMUlK/xX0fpWcygU/KB0ydpSMTa3R3JGr1n+OSdPdLAbRKgq0JwbKM4hJ8
/3JCOc3OaVfNB943PrvJuF84TLzZWwQ/eA4vNvagq+aMqgYUN72d9Y5nOLayJZHe
dFr44bP05/GIsmS6kBMwJ0YVPSCF6QgUqtzUzTECNLSdj4cDZ8aDn4nHNlc5JxgU
ZvAG34m6YEWyS93tnELS8zPjzIbH/QZhJZeSXWIK5G/tRc6dSTgLNtxr3hGJ06Zm
MRPb5yfjK2FMstAmEo+gzIK/pE7ooXoZp3NEX+ypH3e1HGdhG9YL5RlqgznkCt1v
E2I6wDfHI9JnjrzTR40L/pRWGL7RYPmaRgxYgAXiuIWvnmJFKsiZXYSx+7utMeBD
9xjSmYt4baqAkeNP2jmAzTyI2zGoeYkE1YU8rbuC1qpAdvhH0FS2kXcWp8Kfdx+9
dd2C5DsQzU54lYoSCmRAxsIL1HvYZAEQvMbMFh8Ruz5n1Zc8p58h2jjr1NqiHsqw
pSY+tWy65M13Bo3bc5Omlss9+kg0XQgNXmbodhL2w/Hde8+Ynuomhay3z3OPzRL/
tzXdiULLBIa/208JsqAij+j+WzLd1lfhyWflcDHDBguV0WJK6+OuQ8o57I5jDOqK
Yr/NTs2KMQC025WIZf8EZBe9e0bQsP0Pxjep1kFgaWa4tJ7IX4DTxVl4GVdVEnhL
FGiKTdna8VqxN04gwByle9cnTUdfxvqWv/t/YTnjUYd0Bv670vutabsFwhSViE3T
UPI3PpBlog+fsbqz5dTk8yCfzWy+eZBWNCKUISPzNDfb8RLX2oXRrdR5WBbsQDEo
6tsFPXMN7JxS//QGmuNfbt3jI4G4qVCA70N4NC5lIkGDPGykdazcvNkE6u+tY0vh
QPyLr91PQT9kl2IpluqmGK4AHchKIDJig3KdW5VHkc3D73DH0abxjzv5wnmfqkSo
usAchydErq0CCk0goCkxss4wMeRALH88MF4g491yaYtWDHdFDPGVvgRD30D9JKnc
YWkmRXID0d3jgQUWQAGzU7BxEqyEIE0orvYzeX89/APiXODqrsESec8XIHu6/SYR
4iJMc4jYwmvRuqJ0n3wIEG1G4YF5L+o7nL1Gy+nNiZ3utyqGD5vzkoU6wW6wVgYy
T9+GStf5hMoCGtF8Gqj8TvR8CuXigY7Ao0HA7Hx1GI+r79zxA+czoDMx27rOAjA9
VTxc7f8htYH5Ly23WHX0p3G2X8nZM4lngB80CO6OmFhSNww6Sp2eIMxTHL7H1+b1
LpGMcZm8KaBjLEkMCXKAelZNI/HtvdNQHL7BiXljSl9tMWI1LlHb4BNcT1GYFaf3
Dbk4BwPo1vHgHFFYGJRK2VDgSB3D16Jf5rUbt3N/4G0odeul1gmjMbX8xD5LSp22
+Qzd/jlh0iIoHPqQhelfqIo2SyrKxqD/jZXC58pIbTsvAHmfJHqEElSgydZAwavC
9xx6JhOabukMOvuN9ooGw2i57Tzu2SgDrRPKDNeAuFV//SmWY1dMcQzmV22YOORE
VHkvGhq7KymrofWcdFdoEvkfvxCxyKdIIto6/9lSYsVkX4FtqWvsov5X5/vYbNeU
49u3zDbuTLQ7+4LWnvhBIcGna1xbXamT07f3lO8txB5qA4NhFoaduGTsHRPcAqRm
5285wOnnm7dFWZBVdcX/sBtLEksX4XBOZ+qzenQ8RUApx5mJiLuREBnKmgeHxiZ1
WdvbHd0m1FoDu0pUEg7FDSWTt3U6tOtVQ+jhm1iKfLEb1SWq0FBW7o8kHRcEHlgM
IGd8Ky9k3IAFgxO16JZqQaViApEE4cTOYuNw+1M+4PNtaJCo8nbNWNQun3VqjTiJ
Q14pI7PMkncSCHtezKeOkhSGPRDN2nomBa7GYIJ01BSSHGyMlhCjGsuXJqZ2yUT4
mpiVQjTBDC9uUh7lt49sRZoB3wxfQC+Vb01Y81glFQ+Hg7hQPe3I+c442An28XC7
LahUXN70+Y8d9nKApwcQuGEtD9qRd2kIK+gAQDgWNnMkE0YO2+vlj5j3dQontM4v
EzFFBtUYugxnx4PvbdCDfEn1MEM/ejp0oELL48lGLdnih9SOoL7p0yvgf4GF5LVy
+oDhWcsJtYozOw8Kst7nwn2/DbYOgQhvfe7TrGiENEcKGt4U9I5tYk55tDEn+fbq
B5OuSbEl7UbVPcFSgP4IGMinpMtJj6EKjoukcMxIJlHQW2abNWwTDDkBKkDx+xZK
qB3XCsq3tF4gVGQTBaeON7iog3THC3sL8Vx9yrJWw2PhyBIXgIX+BO2jF09LMyo6
tVtvuCccQ1r1VOdCXXYVTiX7RIgXsuvaNvWhlinftWSW1EYD7uqtrGXeI6NC6Lhx
JJQqxI1em4jr09j2MZKWyaoMxXwi/bngisbIwz6qF4xXcZ5ici3XdSv6ZBcDiEA8
TlyBgr4TFkt5OumtintembJ4hLKY/2DE9JKgO8tNvwdA29WOFxxnFANlzqlPrera
dNPmj7xBCdhhlqKy0XyLBkdFjTsPqW4AehpEYbX5FG/7ku0wVSv/093ufod6mHMm
/WXoUI4Iwv4EmwLhY1szuPrCY8cO76XoVacec+vrMmqkTBMYAOwlJfZsqsoxIKmy
swaLM0P57kxq6m01GsPKtNc3PgQCHB+ut6l6jIJtxR3LNoLhU4JQdgXLbcGFgexL
RaIDRCN+7N7k8zZZ54brsm3UYzp9ksnh4IzLarwaOJP9dIFNztM6kztZJOxhrSt4
KES3Gg+xJESIaAZPx6ZOJcyKgAjsW7dwmFmaHYcic1VclGHav1n0oJ0iBg4XfiAP
cyOrEVwjE0t+R43rfQk0UG9CzKqbBVq9WTd8NpRAdfDdTqFDhp1tbj86GRhMxl+H
rnyxtrsUT0GhTM83Yb4RsAbKkz8gb4th+uj4owfoEH46K0UubQyXH4QfFLIae4nc
GHVUDuBiG4NG8FZ8eOn+WVSxq+77kGDhE5KK+QCQtiCRdSPDfdH9QiUlcec0WsZb
COwvoMpQxNAnKYV+KTY4egdBndzRXO+zd7rwx7bZFeboF+hBYZlzlvZO2DrVJVVn
vuCfxF8RACjrKk0QHM8nG05yVvznElfd9+6BfmsHgwGABy15/V64t6ZTwOLcNXVA
1G3oG4VE963QVkS3GtykK0ElfMvImkwTsaMAThNyRf4NKOqQGMYNnDqAz2BKBvMM
pgisouoPpES027JVoYPK3FxcZUdZBgeAYVmh1BPF6dvWD2anUj1d7OTdiKAn3n94
8RQ3uTsO42AtLJY4lIgXJWIRyO1/7JxBeUV8mVeVom73MRr5jMhDUccCbVTyMqTL
2QSVy6lniRJzNIFsD+WR3KGtziWjE1NzgXHN5zZmR9ZtoIRIsdwvPLwy91NmpkKN
/ubSSMkYNU6hMWZlN4QNxjt1vIYgGqwdGUfMTljthjF24PvGP7DpuRrmcci2+k47
ESCfQzJ8B/HnnzJu4jZFkUybDGOxt/j0sBkZRF3bSJToUIAOoq+rRyTVdMZPEEGu
VumN3DeqWijnh6mM/qzu5acL142mLONvPlJ8hmKTkY2/f+JLwxLPiImindtdMMvg
Z0lwn6TrPnpB/33T6SVRa4pZWpZ1+Sn53AXorRgWcbxiyxCLkwpCuXfMMiEuuQja
N2JHukJ8kbSOkdn9lNduTg2kUbNdo0pT3ETzFOJOTzLI/nWnmRf7Bp4RM1Sv7KHz
HeZeFs9jM6SaTokrd3LXrdlc1pn+OiU5LRihM6cWRznCyEb9KDlYW8ia8oqVqS5s
agnfYSwQgmMwjZGHntffjTBaSE4ioTo6WjR+mdV4ooZYw7RldprIQVoAzgyjXJNb
CcM8OGeAT/BqzFAE2DEThM2qzlvQxkc61ftQEbqLur2XulNsNEor5VtfKYHQgnjs
CyNRJtrI2XQPawBLCKzFZdJvFQWoTw80Yffy/Lu+Tuh88zmeVAqEXpffPr7v9cfC
E01sqWI4GP4VItGS0xlf9JferIkG01HMxFvY4OQiTOi7BuchGwfyEgilvsZ2krmb
00QDSQZurPwCDsl2vpKOcwJWAOHWIh7drnnltVb1vY1lTm5KhUynJo6qZ8fHYSMW
myHDNN2jz1Pm0fxeDXmgo+57VuqEw+S8y5KRRH13UA/OJEciNLTtJ8RKYm2WeMQ3
pSvO3Q0xNY4h5isqm1ax+fUFZolJpi5mlPfMweO8sfBWaF1io2vOesiGSI3xkMDR
VIWlbu1dMjZzodzi+DEYLjS2nJWJI3bqvbBqUSuY5KhI1snCHqEiilpuXp0VfAs3
YvOpIVJYB6OX4lSnN0Bob56ZlGC2UXBQCa8+dm78FrunoHEwcDnDY7SscPu+EY1b
Z+5Gvrqyg+hs7f8/jopO/Mz/OFZTMxBQSWLr0vDJhOEgDritxSjSa2P463UOvbnj
VC/G60R9sh7hijf4bmpiX/pu0TZ8yl8GLZ7T8zukZYCEg3lgeIlZRi6SRyHYBvrc
sieXK6Dsjasor5jjj5VRCm5K5QrNWLQrEGfu/bpUEK8v8/623jY1OYY+ST8xrK2z
gL5Iojgdq80veXvC+ZcaJe/T2rJqDlRjUIyXcdhAQf+O7upOL0FiqCSWiuVQ9p9O
TpbCgXOINpYj+WeVy/Jg+fBxwDxtu21VGam1psO7+FkVr9PDYq7v9PVxy1wefSRf
1v501C72BhMVtCK596sC1xnTYbvmv2FGdmpvxLTewxzRLvlY0oRHv2xLYwb54zqL
jYSLb+16qstNfZ7cLNGdX5vBbSuDpy2nb9GvBzgXIoO+DpL7jfDHHCOsKMqFq6Bg
+zG1ZEDi+YkDgCnoWp4sxadZ+RHveoSg6lt/Lssv6Mpypd89/bZK5v7UUdbDVHFj
CU6rMDfIXshm2FJAQo9pRmozctE4fF9UCYgf/r5mEXaDkmzgD0yrYN6c7wJC4O0h
ZQR3q6ujjwXkUDCKYLz8R6eYU1SX/p2iJ1WAP0m/XlGM3xHEP7olJwhJsBdvDZBd
pUAaqvVy9l+wdlU+ri8Jh4eip/c74P40Q9W7uIONKB4cH4q7O4ahCqo3PXO3n2xS
ztegnzrQD87x3dVe5DXUj2P3XqgJsHh05NJ6/xwpmkxMA0Q9PP7f4mGvaR8dQJwX
0zBKM/e0nOSlWNwiHTwC7H6SsbWyF3ttLxT6bhsFohnFcVNhLIMtppWjucqcCE4b
wOgmskDuxJTQV1TYmozPKLfR76eoJ4sS4oaXjIdEunpEaX/YNUsEgYwr8ewjQT3T
FoN7QG3RrqcPAkRAPK7rhKPLg9qnV0hSx3I/AQnXkT5saz7kFz5v+dxFICih2jss
L5yaQafyizwnx/Nj6ieaG3Pg+lu84nqUtpm+L/cnzPA09hpQ7g6wqfp9Y40sIXqa
Y8S7WqZCpazftdJoogQFE7kOiFkTPpTxk9MZGk2t6AAMuclB/Z+f3XAjMRFAmiAp
O4Vuc08s0tsesNNmXVrZq8ff8rwvzzS78Ud70h6IpxEqsg5SB72/vqAnojdZDj3w
aHDXVqZNCaEPXJdtQ9a7nu/RYqtbUVl+gu0eC3U5uD6Je71UCbO1svjTxK2AO5Dx
jlLcirauOs77vngXg7AAvk5Q7fidxk4So7gJNRheKlgbKGf0TfJnXDs0M1KE55Qe
h+Qe5D1ycPl4sYrJp59iUIeZ4GHamWic3weF3vNDkLALzTD7DELs3f/+0o5b8ysp
t1N/OtgeuNyc+TVx2ut1thWortCnvUSskvoLHb8mYSmonD2BZ2uNkImvAoQpEoDP
N5tZ0/cMx+CBj7nR9Oytsv6D5DtjGikmiKs+maxt32yG+mOehi5wm2nSC8iri/Mb
KssYz7tEyA/6HP2J4s7weqeMNDj5/4SlOP2tvah7e1Ll7qQoY+oIPrnkcwOIYrox
rRAJU8i+B3Cyn6ZBmln2KFjOTJdaZO0gZSGCrzzfQslFyYFNS3URSHP9PRqqR6OT
SinLpLtRCDCLRVOqdBHpYcumBY1nYVk4GY1yVLAwrVqiayQ/PXWjHCRDP801lif6
fJb2t066EmfA31sW2LQoEdOGHNy99PsHSLsExTbgJBpzKGtwQJrWVjFm6UGhMezW
YutjIX8LHKaAGYc9Wy0o7Bqyf3F5Qr0mewDRLjo+UKDzV8nEgX/A2ZMmdMDgvOHW
U4KTEdxHuV6gD25fmGJgstHfV73+kL9S1vO4GUX6zI2p9TTAJYL4WMoH+STS+uIg
PoIhbdv/vW/gaYlJa9Bja5WE+tbLewL0fPaA5GWiXsqs6c1yOIs4TXR2QleVFLEF
Qc6Esz8sVSbxWumGELmHi05749pPaIh3pV5/Ex+rZh5l5+HXsyIQu+cxNKfv86LF
Z867fGSjkjMSdeaB3oCL8poYYfovpiv43Z0GO5Yfcoq8g5NrqbIdUW491RiV5g1I
b3bpmXO7DbWNA8WaFg3XJLsljijCIx6ANLvIa2V09g5wQ+AxEgcnUdPNpxm/A3Tn
TXjD7OEOv2r22RrU0Ywr3cWsKTWKvFAu3NvHHm91R7BF6dBIVJvmZcj7UkQgIyk9
cNEOm4+qbSA9B2qZ0vcqJAkHb/MHYEh7ASvTPr12C1rU0gtbWNgkX7U9FpqGs5d8
EfEV/eYwu6uqe5o5eKsgeehFR/EpI/0E5rVNy0/MkTevVlP1hjr3zMP0W/KyE2bj
c6W4P09VayR7epuQHGBzqgyqu3wNemlf7Y7K3PHFP++cU/9ZoYQBN9q/+PSszCai
uG6npDgvCRQMh26hMy9lLTtSr2uxul5sRdcgk0ZLebSyYnFR9lrgGnK+Wc6EJw7q
i1oODvmOOCY9DnS4wFPjhErGjmJ8ZDxM0HXwzmPDt60a1UTGfkCmgszivUMM/oUN
4in+O1OS2eSxiAQOMzD0JcO4HaElEenQ8zK/oHIt5UpDq2VNyHdDdteqeJrF2hiv
74aO2oeIAi60NBVXiZcb8IqJt4z6IJGlZ73Bxz9enpzJjYTcq9qdBTuh1hH3pzj8
FSnXWcirQe7h+cJIwkfPhsQADeCp1311UEpnSF5oKgxcj15VMnF05Z/J2D7MS4gx
Oxvx4HbF4PgETun8L0yZFCCP70RHtfWs3sO7izSsJAF/bPll0rXhQELSCL12mN4P
Ii9jJUevtBvLNUzcwscBK8JBcGVsUP13ezFDpxPYiAcIuH4WObv/EHlljPsGUv2D
pHMwwSJcWVOpXeCEilcHGF1sySCj57hl9QWQoy48XNn+vR2TSkb4+GF2qHRTOZMe
zPr26CO1239tCdZ9RbCHT1aM7DcbdDQFtYNNosddFKRVSsM30v8WVYPAp2L/ttEH
h+y+GEa5GEhDroAi/GirwAb/1wxVGaci8FqYIsNTYpd76WAt7Qu9vbY8XIjRCNJj
2OrFPpxdWscgYToUKosBZPLVGShUuJYKwgB6xqzZJmiI1qRrg+GNXccblO0rCwzL
CjgAdzHF1vB3+yuxdSCDK2bocYK0QVopIIP31DJZuwVpanyLYe/6rEga6NAgDTmx
acrkec9YtVyztQiU0oBSuj80yK6Wdr2AMuzGVg+ya5b8Am0mR1hnc7pKgiKytUkT
`protect END_PROTECTED
