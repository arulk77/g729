`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aZd8AsW6YMve8d/Fo0zk0ILA2g2wWXgc0NXRvQDL5uJY
k7YwUmw8MJrjbMkz0iyO8Pwv7cLN2U3qmjEmwlXytyN3ccnTUhPUmYPE8uZh2Qa3
txGtdSXNHHmW9RPHn//CLrZMdO6kSQG1JyhoQe4hO4c5MCRK1FeaIz4l4eS9w5r6
RbX2YcWQZE0iFalnI8iiUGJDfLpeovvJc5JP2PJmqQgNMbdxwJM1lKlYzJUZl3Q5
vPLF7zuh+xpcWMiAyU9U0DbhyI4aLk8FhJgX3wgHDug8VqDqV3Lgl922rB5xb8NH
JaeSYxNSfdp7MWsnSRHutthcFfmp534Ik03wHTh7gxOs3Q+WOpAGjMxyTCd4o5xs
AKWYRDN0EDhGp+Ff44NH4xzi0LPzuzafoQU76dTcvHOTEhaWVgR65QT+5uQFs+7j
xjZqHFyUJNOs2oQIuXbn1awP6OpGFLaY/kTLKiX3sgzRvm+T9FCWXpqZs0Kxww9k
jVh23ft+023RJNe/E23fIV+1ds31lqRn24yeSYhAGmC+aRNq9IDUw6rcJ0jGKiso
0qYXmdNnErOFgSOxMc4NpGHiZ4GbQXZ1QJZr/aTrvh/bbB+yX5PFxpB7K8Qwhgra
1HjCAeI8BeR8SZDMG8E7Lzn1GK3zGIOpBxJZnG5G1K2oHS1fWNV0OdFFT8vje/Pi
oFvXSaiscpkt0JpvKpZRe/i+VmkL6k6idjQAtgNYGSle/cR8vF4e9WCPydoDWn3o
XfYieEWVFxaZd9upbho7moWuhPhtSvtnCKPbX0PHz8BdX4JZPZh1Ndy+ZeSWR5nT
+ZABJ0ZlsXeU5X6/jzdiTSZ2BDNtAXoYhaq4J9pZw4QdfwGmCHDt6fpqJEOHvKi2
`protect END_PROTECTED
