`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL2UfY3naBHWt7SaTNrWgil0dnXGVCQAUXA0HlMhRrDI
rM+DMDVt9V8D7vx3t6sVEYbJAvgK0VvcxlrVkz2U3SaNS74PGzjtb7j6++fdvWSt
eeSRCzFWrpinqaUc3y6JLMLZ8qxddH3Bbi+DkUSWw+COBaUzCx6Qf6hHNpNEpVPm
Yq/6oBH3njrvf0rnlghCvvFY5y56UnBFU1wDyRMRJqUk0h2tLcsNBSJ8vfc1ZZSV
qXqniI/b82+w9qXtQRHsrXRGWqi5TEMhqFwF8+zb+VVkE4tvI26TVbMzXlWq27Wh
tx1VEcLTaVDCnP+amGTB1La8kyZoiOjt8d2XjbvsBRv3Ii/0qCxtvtMoS3ahIAEO
Ik50X76LHprKhM805cTGKdgbB6k5EXdBNyAhzNUFpKI0YUv8DKWiAs72RlL5QYBA
oW9xkRqC2mlDb9kM1oFOx1ZZJxzG4BAVg7Rfb92Jf4a6SNbvvwmwpcrPDZIoyVNn
N25459eIIgn8BN/gH3zfmfyshcVmTD6bKUaaYGbNAVi3O4W9Y38e3DWm9oxJKD9w
`protect END_PROTECTED
