`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4jUYkdt5VjR8oFbu7ZiLktDBETznpTCrkCGu7b9E07XodzsaMb3ZVz4j+azpjcPy
wY44F4eWHDho0NHQ2fEHIU7QaEPiC0p4RXQst0+uTwvzUpbF7AabbyCIE/HtzOIR
AbaGsmoDRQILrGE4Q2itiWT9F1Oz20CUoq2y0RWom605jzJoTxr94ygnBtCztKbv
wiwKqoxtuYvvKrCUFCTixnOW249maBqcU9h1DRlY5HSWYFxzJAg3PwLY+wxB1k1r
vFD0GM6FdGoIBIzbAGhkXxU4pu5AIam6Sygz3GVSZ5/IhUZapImHxtDeNaowB/yY
GC3Y8cnJ8u5I3SIy1ZjRxyVSsMQWCimpZC/nMdMfuJU+jPXw5K+HpsgvoJ9kpvqk
gZPpGpuD4I8ntwuL93hHoNMTS+oPeuNLo4ZuM6Cc91P0T3WjLtzUhkdpqFgQcseo
Pu43ShYLKapwiXQ8j+u9oyec2LULXkWoeUjN7pazR2l68LEEw53RSimcOvcdth2u
iccsEQF9gpZJuxKixCSvgL98Jdg3k1tBIojJ+r6FR1bZkAaSqCbS2xMKvQw52ChJ
U5nF4idXSypOvTQxVqz0gqlTxqAeXdvVY8p+5GnslPYax/Y/ja/2RSS61vC659s4
UT/n6W18J9qsfaRFujCMnNfD9+jzUZA/hgakTwHNYoY8BW6wPxVIOLMS007PoHVM
V9+cEp57lyZM9GKGDiBrnI0f1bkZZnKsKrRmQ3ngTDLBYT4ANABL7lqc1Y4eyDZt
rm2T3kRLf2ZG2Pv7GOqYMitK8ENwhTsfpSs+zT90v50gkQToLkFAz4uevaJtssev
jGqwfx0F3xNmBFHE6avAAKOZCljf+Lesr+tJhEbK3CZpaedUkolPt3hAZcSGOecD
UJ8DpeLT8joy9UtR5UTjEivoF4cCH60e/WSykrbFT7jgG1Wx/DJ+B46qN3lgCeSn
CBzDZznBYb4qi5X+FOd+6cSI/FpenBRgFLWsAgp3A5sPtJj+ADBQiICbeRRXHM+m
uaTdHzQMcR3+hHz3GpDCVN+LC/SJllXwZb3IaxKHLmjbYOQghgUFPxVGntrNbdwi
C1EEUChoKWHntUsHpKZCzK+KFqPRuNELJVy8wi/+lfcAOCpKJFGNh0s8eAroCAHu
Rd5Adxm1Sq/2hq+tS8a3o7wka/zlPiS2HkJaISEUHaOCqH8IRrYLlTHhdqFUgOt9
idF1Y7ATAlE3jhtegvG8LfFvi1zXb1H6VvCQpN+Y8MvSuJ7V9esafvMali7tse6e
IV7MW5/RNnSj3m57krw/GQkL2ltU74jZ6E26TfeRyBvJzWgbr8MFxsABFNUXKJFC
F0gHTumXsD6JtuI1CNt+gmDTYZ7zyeQHlkJAJljJcw4mJhaMDkEtGFUCQNT0IX9c
M7EsKSb5NEUNRDTq82HjTuC9dk3EwwH0jlObtX8Zgvq+yOAOPimN30Jyi2mb/9ti
oxBQn+3OJR/DhQTN2qIoq3ceRHgH5b7SnoWkZLrcyaoexP5gp6AS49p0RFIzhulw
5Ug+/LbOuQ1yVqGZp8d8+zuW7pmV3B9Z8CfnLy7rbdyAu2fIGbzvvV4RZu9OQcfU
noAPQYyx0hL6sj0XY474IiRFN6qqZRcIDNuyAisqnUX31ZIfbab0AQs9U1ApBRRV
F/CNQ++M0UJKxyYACAqhINo6jA65VQINcpT0LePJ3/cHhn5ou/QW8cEFQUFIzCHN
GZ44mmaqMtweH1zTjYxK3gEFM24SIJvFpdtPw+yjpyNjPLHmVlsQlOwwOgbx4tZt
O5ykVI7jONWkXlanbXlclTCqP5h38/Zu/sntd373tL1JtA7TkNNcZFkq0OlvYRnv
YiQ9+8yEAvW/fZihkQobMXXZAHkKYKl9lSKVbOo0OLrTUXOxSaIzhkjr7mP8afFR
cAhyTJIKcdomUI1R8KfYtNP2bJ8lTIzDFWGKis+h49zr+9O4NpOahg+KJzdC1VXa
63WTOm/FA6PcEiqqaAb1I8VjorWN9PI4+u3KjqwIKo89eUyN3c6CuzebXPX1AKG2
7r6YOLKWB5mi8xHiSUQjSnu5NWyXDpHL7ONd0cU69CO0U6j90K1EST6ssGLHP6Ef
mw6H4wfGx674I02Fa9NF9vbW6b9UgWsFcRYl4vJTl0y3e/OqOLKpKV8kizj6Qamv
ZGp3ZBBnWlZHi6dJduNUA+K9oBwhkgbhUvZ0r/iuslozClOzJ9/ak90bTcirLyYs
NamaboKknD96OgwFP446MdP8wV/nTTWYjQNVeGud0sOriZyqPmBvd1+CVKIEQOIE
17u1fKau2k4P2518dWxiM9PFiFY0VlwnqJ+T89ympcCXJflEXxA759/IVgNwIIEm
lRs9NyyjjD18rPec18CojoPXLysJkHUJjNGxxeoEfRB+Uc8egYVGWr4XIoUbcsl4
zOAWSXniT62TnHIF7Dmwbg2HkokW355NMGZe3pdh6srZeEbrg53I8WzSZWtz7FR8
7Zujinvatnvd4lV9bYUjupq1RleKi+Y5qvzQ/YEzD8kyHyM5S4dKkI9hSHxiSavz
n1H1FidRR8ixEIcXixVyqJ2RkTVf4KPVbVtwwzZRhs26aP9XW4e8StyhfJkW3SiK
5QRMBDKVSZ8xpy/hQPf6PkNsKyb6q2LX4yKNU/6s/RPxXMp5QwFaXz94CXPb9VfO
ch7FLECPX3Q8yYXTtqp763D062AOyyHk2b7rY1CBkHW2HM2HEyTqSRqBsedCI9jo
TxTXroawqMxwut1AWHz/iS8H8Lih47YZ9Xgx5XGq271T922weKRJ4yoh3knn9ynd
H9COk+ESOve8q96lOjS0a7/bHVBmRgnAFdRKR3h5HN60rB05uDGCu2EvBSsyrAH2
mvQ8WWAYWuoOk1Cf0Db6CsUfMqH4tnT8kvRDL88TSrVxSclxGGHxRiy0UARsTyfG
gSR0fl7u27TwsU2hhF0wGRH62MjKyA8oHHVIr2FUbGbxZePtwN9iIpL2kqZsUUvw
xM6s/SSzbq0mS/9SCcw6hNg/QgHmW1BAk5eQ02hr+PjTMwfaHHvHny3p0hC7jCIi
nkJgpA4xTHq2xnJAQ6Gb/ZDSts1Zt7/1JibESPRlfpxZQXtQ1bYRMWK2jQ+Tu82j
99FCTNqENaeuud72MH+wuOZJRlw7RT1jw4HfKa9v52fdVmbVQh7+9SmNoL+LW0Pa
o8cLCjVOj8Vhj9DFAeZMNyZSU7eCaznBoevaNPOCk4/AXCwG0Wr4QIlq+EOfVEfa
UhlI57fPEz8V570D1E6cuRpGClDC0s5jbvAKVuuGF4Ck+Piag7Cwg7/T9eb8bohk
hJwBnscEanHlYHlaI0x4AEeDoZ0GP21DnjXDdDnqL4oAHmZiCXq2FbnO6DwTDz8U
`protect END_PROTECTED
