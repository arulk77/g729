`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNokLKV/alS786hu/OcE+8dFJllbJGNY9bK2aDt1RNKj
5x+BCA0d60MJ87bBzKoTL4GXRgAsGUJXmej0HUUSEVcrmeqxoSaslpIbR4IpKLgH
0GGTROknvlZv1To05tHtnscHXYdMAtnS3EcPy73e1DnFPPjNM/OjFn9w15diWiCR
bR2sBSCA0vNEweTz9qn1hR5yDCBgiD4DMzMFoeBtpoYmvpcUDXznq8GBYXb2XsPd
C5BHzhI2/JF0FRajPMXhKQx//U98eGMkkWIxSGj3a3WTR3FDH2HrI5sQex6siEOd
yJmk+QJlgR3DfVOGwztEVMWui951sf4Vvd0jqDI3KWEJkeAMXugtqXJCKBusvVUV
7zbJd4Sq4Ta7774KztMJA+/+zs8YcugxPA+LdThW2/D041NBirJzYgxsJj7EW778
UCG9D2NHyv6bOSsR6uV3p2YN9t7AZrN83PYA8VNCi1pBcrs7ZWNYnFF+h5kqvLv1
mGaFoNrd8uIY/Tb2YN1sexK4FN48GnVf/hgEZLJ12sq9p+TBf86DgwMrHSirFmN7
8/KZmrOmCONLTb1Aotyzfk8WIWdiSNHKGhlv1Sf1cYOC96g11AJRbQVW32YiKiF+
ALzmpM0+u5257W2makDcL8t6YTtNOJERRG+PpjbhHNbUSF1bTd042tqNQiPOJ914
7OPzxNNjSCh9EZb3MQdxIeGrto/kbZZ0TcwaQiYxxm4aIwCaDiPfsd7lckhzrHc3
MDEcSWv0ueMLdR4mT8R5RerIQrLhdMBpuJPtDwIIDxzMY0ds3OCfb20WYZ/m+8Pc
pEbC2g761DEc8WbTqDzRi99QkxqFOEovNI88MdUZze+8HRrMtcIraIBdLELzEBjq
BRW3fA56ks7RU5mZVrj+M4b52qCAoCy2AnZlM4haaPJoqGekUfD3vA2XcMDhEoc4
oIsaY/+7KSVQfOqlQ2+OnTjXyXP8/pLxg0+MFirCTpB1kb1ZzPkY4dVV2eKIi/E9
KPoT5tmJoKnGQsC5K74oV4dmvHh/4qL8JGfV1UV0UQNfv9kpoTVjSQEkKVqOVY6i
vksVNUjPYyW6KeLaPKqATv6yJuSBg0Eimctl0dItDPZ0vRLV518RnYbqleryiV7f
dovJcLWayjhwozlsTzABNJmINpx4vPA5M1wQryPFB8AJsS6xFIqq+hEfOAuU9oG5
mRgL6R6zSeJLs60pciYcKg34005APGlo9lM7qe+OJTpGkjv4BzXTaKa6YGVxfb6+
fwatSBBxE0+Vy5/QsM6pYjkbBMHOh/plJVsRgqIkkuUyapxSStHdVwrvwDGDOIwi
n4MYJFx7ikFEc3lZgGTs16vnzsS9Gv9Gm1ZMRv4+VYoiWR0USDnjnY9O/pxZ2WL7
KCWbHkon8o73wEgPQJurj8XkpVhgwbTsvV6jMLNg3eZioA25Dwoc1/zv38RZ0pkS
bJjne6nKdhdtU2O6rXlTEE0hup866N08iqzRwaWSN/dnFTsMx8UeOtC7X/7wqPqP
bXmpiy0/lgffNMkYTgk90N+6YrEW98BCKvri3vtH84J8k4UmzPXMzuLqfrDMBdGe
pTS2uUZ0C/JaauNa4eZPG6dd+SzgUaUrGDi7Q18otc6Pzjdyuw3CKpJoM4f/uiRU
n4mfl5hdZiiIwfyhpIbjmh+mJtlIWw75XTAILxcKio/HrdA/3TImMZ5649YxH+07
S66HtxFKe2RFCh+8t1VzRBqhYPv8MXqJTM6ma8zjXfpV1Ppy/6ZxJ65yTZ9dzfkJ
JQDsGIP6IJrTMQn8iDJ+GDPISkWkQfsOVsTv0qJOXgDGgAhzAlc2ful0L/4expaG
tGNz/rmHZAgwLBH8mhVOw+BpyvLV+FCaFl6FUY7cdfsfubHnZr2zv8romZWyZpfk
smoYLDbIZv17iJx6yH4T/8xGe8Utcit9yBAit3J94FGstN+VwocSbGoajgJUsNhi
295OoJ4gjJPzLRenR9mKXBpwPtBFkOBD15c/O++pNCdJVWUlXBVdhktAo4mNqKwQ
242ivWUOZVcJftPyc2W5C6WbkCZ00M0OyZOKbOWAk8ZpIeP1cNqjUuR942WXd4Fc
/aGQJgnKMmQ0VdfEFRLExKec+UGlVRSWhb8WgLIXE0JUDwpxa0AYzlqih+kG7XUI
EX/ZWq0rGnK89J7nYeEozWIYKzUL4Dz9pjvVKGEGy7wiLw/EliSrbL0UdeP3Ht4V
ZnkqqpX/JvyRU33ew1+SumgjzRD08MEniyAVXPBbgK4VE7VzUYGTuR1vPQszPhkm
s9WCmvYPe7raQ2QHWBy6vMxOhVmJoAgbjY0jtwm822DpWcNxwrnPZXbyB2EnYVDK
aCYEZ2bw2UxFBgFWEW3Sk2zxU31KMaREIGx+pG2I94hr2DzteeHK/a66nfhGGgYX
lKUgGU126zLKQbn8e5ADscbJLGb3qkjCqE8B9+E0pKz452TbOYGEQBGPdH6PwThU
VnlIp01yHaXkJ/APaOh6yTfRLPSAHO6vvmOCWGq6TDGKBTjmH045nnub0uZnXv1k
unhPDw9pjC86WXPHEJQiyu8/s63p9jqZoRQJnOpsZ2wYsFKRn3NSLKattEB+yMpg
B/MkAj84TqFO2Nzl/ZNEB+2ItpIsi4p9wBZl60aR2Y0/tw9yZCMZ6AnobcH0bHhB
x8q/JpPPx13zJzwthQgoHK1HnLjPzbnjj1ALTtgIHaB8JJmweGJoxWm6sZfb9PVR
Ug9JSQfnZlrQC2GjdC7iOEZxoY0cb0e+JssEvwk2D84g2xjhLWPFmpcy9HObYtRM
Rg4hi8V4k0X1fk1HN1fY5JrH1mllak4Nh3FaEXH02t+vLzjQYXd5hOxiT3PjzdGp
AmGzBRCm57vhZgeCQGpJBe3sOgA6rtdBh1bDyZLHjxCXncuVkEwM3GccqK9YrePO
SiYkdFm36pIQ6yy78BxAS9RR6tUGPSm/efOC6nN1weV2ABmqj3Rej4TWCHMnYyII
R6UO/Op+oAD51HrZ1etwaFvXFECSngZ+0vo5a+0q8V8LvT0PFaYLKl32ghBgei7L
a57FoGB15cqhrBZ1apktqEqAQSKumlqaAZke3Vm+nv5cgk4ML+Vjn5YRJ0TVw3bG
bQxOidVjvfOXQ54m+4YrOHUyBxmtoLTizYGWrYRr5byM+7/P0kDEUtSWO3Yd3Na+
/3h33dKnI5JFuA/YB652qH/jsLIiAKf/zsbGzlZS2TB5HAXEkeaSYuHoDccVRiWd
w1d8mhP1h6YaPFWEAF3nIa+XR420nyELMKFmcXOTuLRyHA9BFWzox9Xh0co3ELos
o3m4BVpuz0EYxqNed8s73ilrh1lQwf3ctn59VSbBMSwGkXddAApm4pTxrz51YfRh
E1qRpzYEVnTX4W21QbJaBdIXnXtiaa6hdn084HwHHSP1Yzb+w4VN8EpzZkbA0VaT
/V9Mn7UufhyQOkCiDjepWf8qp0m3LwIqcS3m3Wl3uiPw1AmeQ/870iqts7nDmuws
vy1JTmacv4E7OUEvtqA6VI06zjyW8M4gFjcf9Jl5nT3PkjRzHBLZEcl6Lt5m73Ya
Fvl87YD/8mIx7BaUENAffoyvFWHddbe3duPzyBjCw5Ox7YQlXAdI0l3/BMNCs+Y2
0Ohxf03K+tHyoIg7Wze5Jo9J0RbW6lxAAiCyDOcw+pKq5U+TU/UQNAytFR8SMCWO
X+odxZvlGM6id8Gb5TdLhClSZ/nWCuXVuPeeyJGr1Pt2FVdlSAVbUdRGjh2319bx
7hATCErJ6Gz9rVF9iSnjrbwQgQTsK8UGIkcq88zsHOIjEgkuEOQ3DQNY3GZJ29E6
K+wvDO0LTpiSoqOxIOAu8O9ur1DIZZlaCuYQiAxr5Qx2LXb8tqPkLb0jqw9TLE0t
3V7C/ZLYNk+hUQyCLf2OCjv432ZVIhL6nfYbT9QqvXm/qo214Uc6pMtC+Dws73DF
NTHedmBwyYLvXLdqo8L5ySqNsKwFUs4UAmvSprEW18r0bPf9JyvCDPDqisUS3BWY
ieoUc5KPq4ez6VSlVC8Oif7RKxLtKZ51JcJI/nh9JcRlvnCVZlkxgQ5z+4lxI8qs
wFbbY8c8iT76EK4IUPmWqolQZGRCm0sh8ZTq0muVuce18dgXlW5nJ5owUZxO1gQ9
qUQFunT1qeHH/clf6uf5yez9B6vM0Al2vcripD3tzRPR0FukS0EbaKkbifUAzICh
hVup9htTr+Ktmpk0VLZ2U6cDdp82DeOX3BxZRi4J73RYSR5N8wkEi8dgcWH77f4b
Hwx+aBW/x8a1FDgppBlhjgIfTT3mboFmSoTnwUXmirGWPYQUSXkZ8Pi89wSMrXgr
u89mn36rTQgAZxv6M3VgG1VUCcFaDGskvM2KiJdOQ7etBDeUHnqT3yjvqhnKvCkp
c7RPdgmTL11/mCH6Axhmpk9QjsHFb+YzlaqFu9uvFu6wqUSeLDZi7WeiK0EGHWZK
YSDQqs/8rNWHobMjNmcfdy9C0dhPTgLl+qdy2Ua6nsYwHH/oUxMn+iUyb5ansTGT
c+7KX925rBN0gYTIK9ajaDcsUCMrUlHY+qgh7/OEPaYvljkw1hXBvT7FItT1EG0E
YQD1wUQOpG44t4tn5BvSdCQgatir6oJXVMhKxxg5m+n2R94LQNTQRB6X3PG+pBg6
9xTxoS+rH3wRulmkNUqRKkz+dy/RoDXkxKw8HYGkqTc4kZ3wyE6t75YKCqS2yB6J
qfAdyJ3Cj9jd3lQKLlU71112nK8NUNHACUfY5XtOfT/OOSE+q4Qfe6+Ry5FEMR5q
SHPHJYWEt+VB/Mdb9OSLYobYd8xC7KOrJysKcUXiN+gmVvPFRGxqFVH6RZ28EO++
Z2Wq6tYWtAflYXX0TnJJUzzOCuipr8sgFc/f7Z0JYZV3aI7PKOsGKT9ZeMKHSkwE
aHpSCwpPRNkchofkaQuD78mbCVeaTNlyncrtzgo+oO8uHaGRUzPk7KyLn63+ftMI
qwBO7LXMJZFl4xT/NN6kK4asNGR/xUVFS3hNsan7Frhu7CuoNxCZKQJ+OqZ8Y79f
JLasOMwoluI2Xr+FeDRhYib1/MqLlkK3ihiYij+hBjmrwQuGu9ZX4SHkI+cQiL4r
GdKq/v1Q46HS+g5fwOiyJemfapJiuAgawg28UVzKIO5cLSZHThl6+FyKf83zr0J4
7kChAHciXlC8VClHsif4XxubsY3yF+cCh6RH33QTVcqmD4UY/rOwHLFZcj+FQyCn
1a7/sYO763IHGBG0jrWMZzIBDRilezIVRUzAS2ZAkyKOvgrry+VtqUlp1aslBIq4
9aEP6weOLuGna+up5ISGRwZVnvCKxmhiUBh/dZt/XqR73YzTSchJ8iqbuZUcVN5i
vUhWBC6s5i8BYi5bnP4Qhg7Dzfc+Yj+MDYO6dcLBDXHlpWx1BMRCsGymEU7hM65M
fBmhoeTN+KdFPtbbk06ljtqgGFM7Hnaip2019dqEGF6/C7H3c5vDFgKHcIQFxHBT
SIMx7GyBTSXzDRmQGVrzG9MYrOIGKKeC/KW+uxP0oSKefjov7gBj6FvP5yz/vW4B
vqXDjSmiFUsNcea9XotVRithYplXZgY2DEGNmiZeHubahtudl3fveSRf9efGljPc
PAtFe1B5VtF9815cSNQzy4R/Ey+ziRLosX6oZ4+2Ap9iCxL8fNCnofEIqhlybfpv
aszWKlG3PooeKd1QgMQTl+0iKA7TuU1ZzeQj2PUvubW4wcKqN0uBps1vkulpGoiW
fYuAmMAEq98E0SGNFHhcsXVMim6QnGhSFUltt9E+XDpDLclElXHFbgL7DMVklMRU
n5hQpX4M1dYwAUvUqNVq1aCVDDgL53AYcx3w0wUxEZbt7/1QMjF3yf0rTr1e/q8S
+EGyF9wpAli++UG0j50nRA22JlvlIeVYoPK5BU6tLjzN37yFr23fM4KeXF1NwqwQ
BIZ0P4xk1lfqBP9CnUZhbbtyIYctwCsAYlWrAV3afeP4f6lud4a6T77+El2PC1qi
c/d4YY+jzYBspuU1bAVo9KrZ2OaBCJkWDZ1pA15Jdzr3ibzrrgQ92nxOvY9eHfcf
5gzBJ5KaofsYjHCW7FqoAVcUnn6BS1LSM58773+SE0Gzp6WxtdQlYwKrjl6ka32d
XTArJ8ZIJt6y2H3eoXAbDW5XmollysFB5GRvY16vsXDPrwuYAAEGYTKMHD+bgIEJ
j7LockYdIgo6Pu6Lp/8cNx5VQE94opC8IN2f9ft5GCQjFhu0N5yifPy76rBcch+O
i+TKIDCA7ujK/8d33+JBfT5+JGCk/xfhfwSOFI2WJa09q69BfJDCvenPhAtJljw9
BioienmFyUJ/Z6sfDePhR9ljchp9nIFMzPQ6URxTKHyZ57K9QzSowNw74KbW7+Im
5i9UZddXP3ea50pm/y5iuJs4AhgsFQjO0gakPsd3IkyZo5mP5HVOxugcBjKUSGfX
0F86O7GPjvhxF3A8GPE7c8OZ89Sx5KzsHSTxT+xAKUF+JT71W2Up/k0SQLN4xGR3
ptpkf7LUxyR1fjwjE7CDbUDPvckqxqgwbiMnWepM5gFySJf1ByY58d0ZkHIcxbOT
FNcFhwc+NJx2YFTjTFxIpsXneVNDR2YcxBAlL4I2hWRqyU1wFf8S1Z/PIgoxOA4U
iE4snQcJJmBPB8RuhF8Fx17gIaWSevxHfjr2Mo5LeYynQ8X6kmRYEl+wwyGcN6ih
sPUD8fHhxhr1Yk2Fdt/vpgG4yayI5lJvD9sNx/H1PdaF7q25YiokB9V7eMl4bYgy
3IqghhvkhUJL9ISnnL1Jd5tVL9WzZu8pOF3anKI9fOl4uaVZw+dq+e0k2kEX915Z
Lw8o4+vgTLMN7IFAwwrtX7F7mHjq44i1kJVwBXbmXPkxlohJ9Wg/0Lr0dHTZxBhA
rEko7FokEp6bbKl6ozu3idMsvt4x0cH2id271ftBSuePP18XB8SNLjAu3JRzWkLd
engCLGBx9WPuwLKF9IYDbllTqPX01EBoUAsMZTtVVvdYnqycyvbbbnquU7XzrXnD
DjKIQskGPs6/TXhSFFuitkSzyf+8tBt+IHeFrw70moXl+gf2ltxEsmSCfSrSDeE5
2GUsiwscjCW3AUJKTeC86zbktgISYublqXc6eO+pcQqvVXHJx6B4pY3mbPDt1Xuw
4ETh5taTVObpwzvGzmlq1k2By2kO6NFbADuYBNQ3jHEb0bw8Xe84gK+uvvvha2++
MXoF0Mrs2T+J7CEj535IPw==
`protect END_PROTECTED
