`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN4Z0L4yddOgou275gX+J8xLP+mXhv20POK4QGumSql7o
i6aRNTY0IIfWTdy+hJeFhWf9csIxBFA2Uc8sjlZXlC7nHWQnURe8k/BKHGqz4njw
bwmr+ttKyL/sCL79DguUUJHrkMXRGMR5LjLS8NTcLm30XLvqtlHiRRcL76RH3jTn
VUjxU2qIb51o8c8A7uNgT+W6L2kbpycjGIqzr57AhdJb5QaV/96NRxT7XIxHScJ1
g/dspo8NfiyqKO1lmXLqaaAI0HZ8NPgWnwgOFFBEbilDoiewaIPbvtFlUrcrHZyj
z2Hgaap+ZBXruQoPJmJTSpj2Zu+JTGq7LCNJPoMfjdK3GpvTVVWTJwykVQWwCibp
HnZl+KQLjVk31K2Su1gGeKPTv95FtW1HH1oJoJv2t75booZApA3uXBYSkNMQjsGa
Zuv4318hzaHS7Tq7kaOlLPLRY5uflJ58Nvc9J4jVbkhguA/8Hvqjy5RkBvlFN2fb
HowA72TSDOuY06lzeOiEy9mxo9TBDeR8XQhqDKDESP99PPCmGQYGb9XWPAAeNbMq
Um0j19ReRY/dpNmK1GdDHSWu17mLRpGIM2NhSlfWJx3IU/BV/6y3vV1wOnL8EU1r
9+1SE9QHF+EXic1E0wzNdu1oRejaPu+X6/xYcfSV5GDWJAlkViMRc78hvEijM0Ur
ZYmh7Sb90PJD4Z2or2Bdeo2r3pbsSpnJMwkbnXDYAqnqmDWO+yTE/BcxhyNz4mwG
cluGSc1r0GdY9djAq2th6w2RAY2+xEG9LRFLIDFllBv24tP+TIHJzBtgm1Nq1cLQ
W4UeTJzbeAb8usKJdc2qNMFavSYG8mT1Tn33051qVb5BljmKPGGP3V0tfsupr+Oa
FfRVEMTGzKfXB315lUfIeTz8hOnqFjoMHYQgtl5p7TRHoeGUOgyYD7hFiNYGkAQi
8stcNGJEhMqfOapYY8himtd1ou0Lgx7qwSYUzh2oyOI7AN4uzh3XjxZw60fAzJOO
IdDe5YKjb1gbnhNdBgFRJuyyQ04gJAMWGch2sOX5Rnw67HSsUimf7V/FFh9A8v85
g0Cq6UGnOgtJC/B8RxbR5a/cuAeciicvY+xF3UxHrIX/eefBKFzSetOv5I/0uCRt
dQ/p6LaJV41+xuUUICMN6YS40we2bmlFP3oelm0fgbYVG42ko9rdZ96Joo0mvxVV
CoxiGjz5IYAQ40QyTo/QVTxccLp6YpXsKzXusPbwv/Qsrp0wPPStyD79PlVskGgy
IPBnujiCVMUCj6AfsXH/OtXxX2esoQ8+gLPLS0ZXOm6LWrFsiwuZkLqKlls1USOY
1RzcIaddsbYC6PWtQ6eE6A==
`protect END_PROTECTED
