`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEOr6Mb+tVHhedoPZkJdYKnq+Lu7OAar4NfSeYvxqXYy
ZyCfFLQ26HsMrMd1D392gd9SChU0/YDvLvG1M9QWyJqsnCBsSYPRYp5+k165TSC6
hRDJ2K4SUna09/ZqRp4gS9fOCANzRWBleEC0RyU3ucCyF65h8On78+2UlpnwjTnz
+06PMq2LvUpYvxsi4eBOQDM7vcMR2KwHrvWbAYn1GrVykJGFEN0GvUXYcZryENZ1
`protect END_PROTECTED
