`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49bRhPQVKXn6CjmROA5NJShQoSZL86nfQZQ4wNu6aJE0
Lh381xgNvR2NhVGHePbt4EPYvwWKvwV8RhEujjnSbqFDzDsV6M2UN0ACwjTwEiQ2
VK5EBIRinWryPnGOnuQRvxLO4BD8MlVBS8BcBhZB0Lw21s/QvUmVmT5sCxCTMA+y
gY2TkYq9rRA1VqVFqvuEBTPPFTtLDr2LTiu1U6UypzIh9dinunxlCWn1vWII+TbC
6HxtFLfiB2CauJ8c/HeIOZbtsWdn2Lej0crJwo55e7Gof945MhTuNRTDaYabG7uC
TEv6yl/Ql1ga0ZBbH5gASo+j4wpFsYnjlmiMQ8C8ae+soTupFlVrBFDTkgZ5kVeW
UJl5fCc6fq4JGjtIeOJoaA==
`protect END_PROTECTED
