`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCeC0qNjsVZGfYpv6ZxurHmukoVYHIezuKHmRNZcYqW+
IFq1PHVzLGQkKxCtNvd6NXa+pgSW8rSJJ88cG9QXL+rjWZgqm7SIXPQODc2x3yom
reKfejhoSWdVwxWTQ8Q7kxLY+ZyMC+lKzTWq1jRBz8iQMEXUJxPkmcMcsQKHtwYg
k3hGng/vU7RQZaQCG1PCDNZu7rC5JW45zHtqebNyH3dOo1nGk3ZlEKQqTuIEYfu3
pf4+5OWG/K+HABOEgQjJoHCIuwVmhu77c+t6p2xr4NFydcviXNbF4kllrQnSZNLM
a8GDikhEnOwY0p1buBG9Fg==
`protect END_PROTECTED
