`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGriS0O606R37YXu+xje0r+t5q2vQDOVtMC8okpF+zZK
UD4yJpQvmrNW+97tjq4UpC+rBhT5W6VBZRcJzlYr1nvFZtFRxJD78DFs7Fp1gRT/
y05lPQeWL9sbDTXdK21kpCEjrLVqeY9JSPECy1JIz+ImvHPzuotlNQOvUzqKq7VV
Hb/y6HYMZ3B3WDo0ipaEB936enWcEjjjrz0ao6IEXbxaVA8l2y/b9fDkK5L9eZEZ
`protect END_PROTECTED
