`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu454ow8RvlxyUZoji0I9VlcUscdEJjTc+umuUu+jAKK4D
uqGdEFC8+akWLDDz8Cz0Y4ix5WdSUvDBCmaCnmqDFuZaZ4XlZ5B1i/5dQJhO2cLZ
s03gU/HLN9qLG7tJA1X2n1MJo44TE9jdxgJdxcY8tddWHW0uhemr2zY5ZqCS7q2j
ID44CVLbXT9QPMndtg0ZgXlzmEP2lKiy2i8luWzpQy4+kn6JVwUODP4W2TW2UtCs
8WEMGfoI1hnwiK235ZXkSTwovh2BcCJGkNC5sKDvFMU1+Zej93uvr8SmhWyuraNn
VXcyYicjzMFr0zDiyJUflQ==
`protect END_PROTECTED
