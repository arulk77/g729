`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
lN4nr/xCpvZPj/ok3CADEtJtKnRw1Pc6RvQ4Z0SFx0fwBkhxLtP1ZztHSvIAN3hH
7fHq5mOPI1CKzeGBfySH5zLy3FCdBMuROYEctwtFccKnF2mfTokYQOUPi+1Ud4H/
yyccyhojrmpbavSZInutOqF7IJfJFBSyczhnLqOYQ5yhePDBAaMUrx6Mt58FGouv
hE1yNXfXhtuQ1FAwuQicVO5cTCHpsdG4CeD5YyQznYh9S3PBL9nfVEgnBZRMeekI
V0Uzd531PrF2dJUKZ33lBRsR1qblo99tVAGATzRSBL1zBvo2azFP+n5q20BFXEl8
FCDXiOM7QLRYFb+xGLPadH8uX0JiHc2CENNyhhB+sSOPctVOraT+bHn9wFhIe2+S
E8W4IhHBQu+viZYtcH17o8a2HB+SYOH9FOdHKMdLVn18BUu3SX3wcE71yzC9Kh8/
EbIxlCr/TEd65CMoCAkZFNwyJuaufHNrttBVyIAEJ1k=
`protect END_PROTECTED
