`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aDZEVmmeUSXIlN4WQQ8o0WaLsU76TiZ2JgTiDMuTgY/p/+Wwb16cUrRUKgGnABUH
nrg3dCqGuJIxHs86NoyKtrkGhyPFUdzmyCl3/Eolt2uIdhdi0cqSKcrI6Ml1iRqa
4B4YRVYe164o8rDpRf8STkwx61Jaw5Rmm/w9YMMcGIOrwE2BNqH7J9xumPxX71HS
`protect END_PROTECTED
