`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCtm7jA/MXmj6pVHO4+rdJccan3u8KJLZ35UHztSmVrX
y9vz219FeLlLPEVb5JYqQbH/E1EGJ8QB8+UTGzaZEAicKIIynvbkvTVyGLho2+FS
UO3RTFOKOuxhLhKNXhKhEYrvgcliIyKOKWvF+VwSFBSlh8962s3soFDTOsKV8+jJ
hiHYi50IYK4YL0wmX2SOsg==
`protect END_PROTECTED
