`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAJmKR/c3b8ex3mxkT2UbPpGBucRqhLwnty2cj/ly8Md
DP7xGqqmUoryKR6RRFDZr+zG6+7rD5x43A23aO//ycnrW3LOR6aW6usGsM7src6M
SWzAYF40902hwsC6uIZoMMzXKHI0FVdOHhi6MvtKs7BKb+KSPi+ZKKrNOnNO3rl0
KMwKfvmCCoh7hNEEgSFNug==
`protect END_PROTECTED
