`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
W52by5FksJUdhgHLv4Ym9A4G6smMA1Yg3crfUao4pbrJC6Z7KCgzU5ph4Te2MkTo
qzRZu2XdSJdGacCl8zY1uywz4HPhVe/Cl1jpklYWchx3T0s8mfkezF+pxVTnKoeB
NH7NlTlxUKc/GsV8Ugt0jyf7EeeedEIQ1iGPt+C7vugQcpDyeVTke66cebdafq20
TM8kSeCwV4zxhf6aM/GM3sVj2ZKHtnS7GTLlVFbVtloeVfdJB5Jooa2XR+U3GuZq
ipqG4qpg5AR8GzVwoqXpUHchxLQ9n4I1kdq8DILTfB659610z2t4ucilixO3A6tp
`protect END_PROTECTED
