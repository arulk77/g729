`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aVt2nubnIFPJEkb+9WAelkHeIarluJVNa5e02kSuftIl
ezuvCLsLwZ7Id9rreALhjW+x08/iq0W+t40MgSbI9uuMyUMkU2pG6yQH69f4FrLZ
6very9IdqVHCpWQJIaggpQde58ABwUQsKKZdlCT2LOqC98O7o+12uHwM5Vj8lpMR
xvzMW/bKVCfmel0k4OL9tgQsBrDqbWYw3F0Whbce9MeYYHxqjKf/sPGFdRPI0b+I
I18vJX34V6g76kuYL7DOF82KwQm/CSswd3Fw30zZ4h7MRaHEPE25Ba/5nRePScIt
C0yapzauOLnA3OIii0kktn849BuZiV0AQ0vCLfZ1BNTwygrgKJ1ab3Hlf/NFQCiG
FTGoX9cjLK6vwp8OzyDkEP39V9wdTqa4/IEgUYNEg3Q=
`protect END_PROTECTED
