`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG6Fp7/FzxbxvRzkd6Ic48TpJzh2aGoOnTcfmYcLV556
o8/cgWTccISH2lAMWA9jUj13SVJQJsTXLukM9t4/xydNvFet6hGOImCeJINBZAJ4
CoW/igQMu++nH8q5WxxWDU7PFrhmA/ldMCUrGnui+VyFPtsjZvWip6ok0obmp6CS
ztdgJ7pvyOm0B1fGdEyxEg==
`protect END_PROTECTED
