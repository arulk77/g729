`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNzdW15j3feu9U0XFCEInyDh9lFotUoxdE63x+QFEslX
7BhnNSUzurvGeNl5VhoXXgBrTmA+cjGFXPdidhSNTR8A2iQAcsyh6bxlPwlYUg/X
1Ea3KaOXCPwFU4eIvFLqpvHKAabKgCR2Vg+tLJ/1ktbj7UQZ88DqnUNFK14wVqip
Qcpjx3UKc3z+dPRBnq1OiGCwh/nBZLvZpRK4wg9JadXR+kJXnaMYwxUu06bj7dH3
O4mveb82Tu6T1aLV+B4VTg==
`protect END_PROTECTED
