`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHCGuO3jq7W0opveZE7WL8rxBcNAsFd00rNp7ZaZl6SO
Z2Sd9LD8jeUSI83Yz+x1t3LefyDXOFHeDYF3Bh4x60GBgCWVQa8dE7A9D83ImNlQ
7BwX5WWfk4H2Vv2dXKbvpJZBxdYe4xmT/Ji2SHXm+91k7PofLbN7/MibNpFBp6Bf
hk4JDwlcIcxOoShATDqOXsnEeJUTQjN4LTJk1ERoi62CPx0j48lhM3K3RIKH6Ksv
WxUEs/Wz8WZ9pr8YYhfpWUt29DrZ4GAd271ek1dokSe7BCAlwUXdMkY1ayTfTDhc
uknqVA4lz8qOBTAWuPb38695m5LfGzbFGffFmGXD2PghcAUFggLmJZSLSWJbxXcK
snPqyvmrGViEA11ANBtjPV4R/feayLBHcV6YZvmwc6xQbSo7HcrjIpkZI9zok+zc
qhrRWxCqlNY2dKY/jyGVHurRHgmf3JVdQjt0przTQmOTr+l/egtq/JYAIs7Vmalo
3Oo6+nfsJE6DdI8NKgUdM5HxnUz1i5orRcuRpaW0LMOUl+fjuCEIvTipm9x9l6P/
mVByKKsZ2IcR0F8gRhOFHPa/kS5Aotk30I7Ud828ydHyZAZvcyo5DnRnaJVdOBDL
1/SqJDUvHXqul4ob65cTDGd3c9mz6vva7rECTbly1TmEricRJuSD/SAGNEyKazlp
7Yvmj5q53J8dBFIlz0hP9r1TYACwENCK+51K8s5e+nZSLN4Ojlp9jHeHakOlT1nS
a/n9if9Wo92hxpkzTlsfds3tOr8Qr5CisTYwTq1h8+NGtZSHQDJxe4o4k1gOxowW
8Ur35CznWJufXKuJRQztMF4PW1t+C1/QyzHrulbYDW30Eczqicg0rOYl0NiylZMz
sV4I9P7AHiHL3nZVA8vvu5OsP3Vt9loNfzN3R2PNARmvQJVXwwnxbA2OazFXM+bL
52PsSdAMRSKhSG7gOCNen9pqyYlbD38ZI6j7EPxXAptapKQt9acsgIdrXLCFPYay
VAWRQruumB1SLRgHK0gziatrHyl+39i5G8qNfsWMLDNfG5dykir6bUaOCqdoWoFH
rpZ+PH9+y7mYdKEp4Hegali+dSBgFazfcza/k7JAucA=
`protect END_PROTECTED
