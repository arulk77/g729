`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
AbbudKXJ3ZVdktf1WfU48iL7xcBZES0T06XD2qLXXtzR+6vPp1cFnlTj6gEp/9Os
xSHXw+PgBl7MSO+HqfApmIIobT1sEoYZciGSca6dQFCHzmSl47/enEIyDsqi0dNV
PG3dCugnJkxOEF6E9hkGrDkLFZk/IZRXuBYFE5kPpkFU75HxE3fRJtbAFr7TBimN
`protect END_PROTECTED
