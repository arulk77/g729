`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIOVagOKIYAoA0N2+X0H7bm2RwnTpQYpsUMSyWGmsmOp
/V/Ui1f96R6hV6DROhxxGlp+uLeIpfqQxfy/I0QnsJRs8lHQyPLHgTgzCmnXCgBb
vV/WoDZo/jz+PTtvDaaH4em8Bs6n3GtwBcLsRyTKSHeoRTYtE5QS1hipxXgr0fuM
OFwbnDrnVLb3DgGFZhPtos/42nZjS6OgQRvlUvm4nBZRbxT0xyHcVaw5DzTdWiJg
oKJAiX9UoIRO95EgxVK51ufnsQhEB7MQsCjQvtO2+AHT/ODBLhkcy8qGhmvAYtj6
8oSF2qpfuRHduWiabtqL5JwFR29kCq6kHbqYbIF3Be5a2fSegOqzHH4QIyN2kBj9
QXdsNqq1XZBWoQbm6ZaCghZgvOYi6x80wDFDfatIK4eVOE5RfwqT488Rhh3MQQyY
GA9DOz3GXaL4e54XWJzSTUVr4ges66rTsQRw6rohaqs+dw4T+hfg75V3I/Khjk/5
InBZbbkvsTg6xezkPSppuYWqojG2rGQeK3OoTSLhQj4+l4iHVuiOcE9FjKIkmqGL
8Pigngp4g2p2NfjXukL04jzdjWi+q3id9VSwRIAt98jH9IT2ZvXbdgBTcD1857sD
WUkWevLkxfD2pLdynCanSnOgqaSPk2KEyRliTzqOZTxtickxDYGkyQVTSuGEO3G/
X/at4qUl56hkadWWqE4iTD5/sLtBuYu0UvvwGL8r4bFeCGq/3AZREM+YPBczUyA1
g2ycpIubZcZX2x0xvFA6vw1hUdPI7WeQFxpY9nZzGNLP9ZJfWa4GrIZo+r+ruz+l
UZrwPmI+BWog6sOWxnw/spPeHpzULfCV5lw/zhxRqQZsWDwjmq9XB+J5o1xPed5s
G8RNQKChQFprLUM6iD/UVRazKrVqP0WSY9hGTvX690DwNAERJlVLw5swMn3C+jAL
yszVHoWL3JlrXrugL8OjFnyNJO+hbkHp32Dwg/VGa9hGFUBUhCxsMQ+WcW4p+kPv
ZwWPrzFnrb7FKokNMGbOTDhMH9qAAb5gBj+s078WXFa2k6ZuDBunwSczVQ0cBJRc
K3d3bYQs2H//kub/4Mkc+b04A3k+/Cx3rqU+siRG96QG63fcq3uBAn4bpmdh4EXg
WHV4CtxB7Kzre5WbP477V8+dO4kFcdV7D5AHbI5po2XlBQxPUl7zdbMN13F23zLw
MZu35VJaz/yc+tXyGZnEPd6WqbVVCh7S0HYgrd0pb1loNcjfPJBgGRto/UAn1i/D
++D5afpiqZA0KgtgwXQRawNWvjUKLjVeNKSWSnxB1kH4OeTGqdG36lMid5p+x/lZ
m5PnwHwaIq+NC7QVxVlO9r8fEhuwFpWI4H/aUQGkY0BeqZeFmxPO3j7FVu1B3EX9
Rzks0sLygHdTiFV5XIjEaLCrvQ7EINoInKNo6kFqRCrh83Pl3rf3fDdHzk0r6MF/
zdsnYc7iI6VOomw+V9bjTGucAXxq1KT7wDRp/2bNjjtf1Rj8VN1z7jcliqPtwkm6
gLHfrwo9Pi9DYAT/SzDXtApvq4QHqGJUh9g53dddkF60ujDtiRSdx3wkOlb1Cp1I
N+xn8BMYLG+tbinoP6tLxN4U5RWW/nR7xePSx6yfbcKZK7lt7BE60INGsPa/qLQZ
/jOHK4SQ0bGNh2OwtnYWHmgLA4WQuZ3tdGBHvLVlZ9mRmmnlzMz4mHkfW9hMNliP
NpRbrY4n04SNJ5SJp50Cq2t5tNG1B4NxdbGNNIkFMiF1qWBFOkizbj9GhhfVQMpz
a0Pfgl+s4Zse4H0J0kggO4Mr5MiNZauo/zDHb2NYV+oNt7aFo8bGkvJDAIea53CX
fbduNVV+OIIr/7hGyqzWL3ARgqb2GjDDgF0eRHVv70Q/TR0eE+RYHoRSjMVn9n47
SjQZyS0mX27zfGX34JUjt9RGa2cZXCvdxzuN1b2qesu8iXtU2mcSuwUCK4sbUx0Z
gWPOnfu4ByFv2ehuEqVh5bDkHKA7n5G2Z76nYZX6RTsWhx3uIU14JjnvdB1MXeMD
p7MmN2MX4mZVq7Tzkuy5WuLzspUSA0Y+r4GiCebQ5Hgry6s6wJm18NWy9CWgBuWd
/RIiCT5yzsNfCBt1TXCr55Gm70A1QCcbMMDKcGIPoyJZjMTnBIAD1syLeh2jOoJ9
MAKgNVLA0D9XHOX0lT0T+H7kWipKOU/bzdXp2tFxBNSElzQ9Z8o0KYL0rDkFP9Ja
zCenAjq5Tbb1wxTRHRQpxYcY/SrUY3bu+2W0JM+XDTe8KONfCoLx0i1x8OOaxlKA
XJBpVNhFRGWbndLhl0tyLuKmqkuPbV+If8Fab8IDJurMS5qlTKibMd2km0NoiWAB
ijCOJNO2mQPqpB5cRVdtFvTvjQCe/36fp+3yBBCMd6WYRs6hFGeT3Y2lg+egasb0
QTT9aw2I7e10i5o6TzGQcOTvrpq5QxybwiJvn1TUJXGyl+q7wZJTRlazx6It5sjM
ZMd1AP0mwErDEXdDDJib0PuocHJgg8cOtKgbQq5I/YP33cO4Orx/HgECRigP47ks
pebWwI1H4TrVGBQ600tQ/HlLjgPR/wVPu6UcgQWCJz5dfauWcOEEKF5JXZ0ShSuE
r8eSjYPMOnEPDXIZBKBR2VgCbncWK7iy+6mB5zp6yHgFZ/bJ5dFaowcV6NhpZrXV
my/bkmSsnuEnsL93nTzjxTm1ibZtYdoGw/jl0atBoZ1GWh8D6uoOsbKjNw6ZKmS2
wygMTcsleF/SsigsX+4y7hhq1ZhZrK7SSeOcg+IPxhzl1SPUgK82ixh95sp9alig
nCCznQxsIEwo7AhOYi36ZQpu39t6t0/kCPA7k/KGhzbsjXHqP6wov9lMikWZIQo7
d0IBrtbF1W/6EpD2aRTGM4Wf1g5xB/SXP1jO65Tg/cAE3P6VbWK5TEdXI/e9Nual
cgzxHj5YDeqnxU44C9J3uuLwi+iIZ+EKKoRkX3+VWT0RKzqv1VZlWy+AlWE1y+LO
xY1fTT8CZ1MBDPB1BzPx4D7v+W2irXyhIC1hmDA4w3NwQdOiKcm2GTZZP5wxuMad
wCx4mfZsrbaWXl4LuRmvyYG6ENzMaDw+wMZKiSsHBBzlZ7wUDGyRwUQVyqHNQEXl
tm1cXzrFswzLB21z5d3MJDbwNS9EU2rVbanc6YYAaq0umfX9R5W20c7JxelDhMFq
OvUT3a8OZLyhLNGGvMcD8VfEG6tuabmL8NyouCEWUVPnuBo5QeVpQ2rUTTYtY0Tu
X5C2qydXCRHSrcdgBnA5YYdM/gvbUy9Ppr27rGuw97+Z38POyjMnvkrDOoRCC4lW
HFwl3CYSBosGMOtLGHLLg3LAd82G58UrCWdU2PuyTnD5b3aA4qc/kUD0AYgUiRoy
lf6ukdHtx9sAxVg/+DAcOmU4WXoJYCzwhSiuKe+K1GEIcdPf+eyModbTPjxvWmFt
aGXgZvrDN1jojxU+08o1D+bzvwcZYRfTKKOEfR/llZqHWbl5PRen9x9M13Xs2/9m
1cKMkj/BBM4p+0WbWEhhqigTnw1cotWGw+6T1ZxjsAxeSGf0vzboYak5LJ04lodw
TZUOR7/MqxxKrr2RYinZp+OueqQ5GdxwdZtGhdT0MoTHXqKAgrnyz3hoQUzmTG1n
xofsVkKuNXMXwYZosb8LyVXvTkWFatTT7wBBEuCJYKR9CWGVgZqKoBQoX0zcW0gA
tYjw2o3CkvuUDk82F7cs5AD3frq+dcC/MElDI1IU+XhhmWc7xla/bGrrhnwJReCf
h/BEB309PLVryZ+XrowAOE6gplx1lDophaytQ0viQQEsZPBfTEkInsGTEsfb2FBU
//qVJIMqrFYLfb4KsmXq4R8g5O7BfHJ3V/S00vTroQ6mLR2ACcWnISNOuvgPX9ys
iNkkjsF33K4JUyAq+bD254uNfz13xnMzZHXyTTTbRuSkDXWaF8Nju9abVL3gEjDy
iAtnDiBCtQu3V4qL3qliqLcdsAas+nrNDHpQKiKyDIzds25rJRjPb9dWo3O07oiU
EjtxCns4RsFc7ud0oo1DaqAwiBc8Aony/k56GgNyl29WCL9nzJoMmWIyY553j9Oz
qnfWt2+2Gv1Lr2ucXvtN1cOrJRdBB1R1SvlochB+QZ6XKkOAB+OuKHXeJmThD6ae
a7t2xCfi5Eba20W4Qie66wMjFLTskFhcVIhFri/ig54VQbzXwE5bADHvJ4GbZxYP
XDky16cefdeEJHXpyiQvgO+nnwisj+C0HWW3CveRYld4patlrImzK8uVz9HRmur6
xuFsM1JFVJ0Q0GYDlck/3cM9b02NZ4nYkb7mPFVa5XwZZS9kI1Dx0ovx6DSBzGaC
X8SPyS3AkkOPmaPgglQQ18hXUwARvikeQeXoDiR93METGBkx/wM81ifV80mBDCwO
Qwd1QhRJIv8PNMaL21vyXM31FEIsXpWnLgjE76CIOkFtNicU7IRtuJ7N9jMk9lze
lBQRKdvY0sljhuS0nr8/d9GThdz5Tf7sebhFXCZteaIo9K0RPDYVVZh4a7WMRAEg
j4fhFL2Rg6ljbQoOBi/yiMgIyoz1ZikLnVceS4gA006Cm/11HcI1MAFFWT9PdZUa
NRy4oKfGgYa/jBSIWGt3PMFt/XOMx6sImmJsdwuROPMBj2IQTb5Bt2qOto5osDoO
vGpvWIRZp8/02cQXCEK2hd1933kp6IPGhrsiBNkFUueD7G2IiyAZdKb7smYII6h2
yT+Om4U4p2FKfFVY8IZOiaSmeMWjF4R4znOCFRxzVz7SFUvkTzfAIMxvBPwnI1/4
ToCevExgt461fB4hXj1yURMmvg+AA1u4yLTJPWxxqGRV6xl2ALprC3UGcJ5g7Mwl
7IcunkvvVshHhSvGoKKZ/iXOPrwtjkD9FkqkVasM0zLEa8bLXD2YBgr2U7vELkDq
S9rIFs8j354HOzNCatSdcSU1ayALxj+gqI6AnjL1O+B8HmNLc+7goSLZ4ovN1Jlr
E6346DBqpVjvqBWbXkdHvKHwnHQY6sNk/1n1zzhRxRA7mgOjxcX6KoWv0ZbGrSYV
5eGEE5WwwardracUWdi6MoxPRhmEXBA75308dtYhXijEt3mZbDNk0jyw/B9r9mhx
Cy/Isnw6fstIYDVLyycKucnSNWEUk2KKCONgn2sHfrbid4+r3cz32f0kIReLq8v7
tmWBgky/B5Qng2lB9c3Rb8ubsn5QouHqVKtpP7W5K6xeqx8VAteyp0gyzK+pde2M
ZMD1MuGixonIOmUSofyTOWoF7ShN3vu+Tb1oUXGZ4d7Dsxc5+TWK4JGWmu+VOVp/
u99GltbM8KTiMSTQKTNdAjYvIlP40wXPOcp31YLmlhTpc+2GPF4Dg2CWCT+p6okE
KMkm3lKGrIp9O9pv2N+2AXJPdpPclGANzFnWD6l9BAQMudzmtmrIdEZ7QmC4garM
Oqyi7FGLcivNaFNG14lmQZSc6oUwMAUNPkYMA1bMAaGsv5Q1sPuS5r/E09wwu9e3
rfYHxqCAwbdS0Ev4PzjQwLDMRNU06AdwccKiipi4avvNc04lSDYYsR+5lyfD6x0P
PRkqUzFknic2TqLlIoBkSJJuwkRopge2wmJK+Fd/2gmP+yH6wHK8xRqHmV+lV5K9
RUXVmO2Pu0v+er5EcU7ubTMZxRtklqzK3XG7ONsl8H6LjGDjSZDHB65l8FcOwWRv
K1BNDyfYEFRRdBgsgOSAzlEhvOpaqU8wKwsXZsEapjjCm2rpxGZ9jWlJIrzDCBQX
em4wBt9yoyhUpHoBXp5eEfUEckeNGV279//BudQjD3FEOmfq552Vr3+CXF2axtan
4AtKcX1+/razQb1/pS8N7qrhUB7AqMKAQmVusLcP62HCEg0EjBcg9DwWkdvxOI6k
Uxq9P0/ROcB863Ytzprj4ETwNY3uwgOpRcaHysfpUt9Iv4CQtFgo4N4mQUMqV0QY
83J5RBZQ6BQ1z3QMI7PB4eC0O+ak0r9pjvRF5a8sn34x2sfa1qJV/jFB3bAIxdlm
ayl7kUyET6sAEhX/7FSYyAMqUZfLtz+nr0okKdZObtgkutr3weAJAzko4dAuU/VI
GQ4EkLqhDNCoqnjbY+k3ALQu7b9Dl0zvCO3IOeED1yHK5KZlTH2Uo0lQw2VdodiZ
3mx3vVElYABvPWM3fZ/F8WIw0NOy96SGs+KwKwnKRsLhhatlt+2ZHKJCUfd536NE
g8Ik425fPnih/FvIX1kjNt8vKOoodU26n0PodZiCAArTqy/xz9Mt8EU0fXhafXNA
s4G1ghwOguS+ulAMpsBGXmg7GI3WpoWo2jGfk4g7dCJb+uxhMJwXKh5puWNoeAv5
XFXQA1E/oKa/pA92DqVltVDeyko3pf/k/K5mxsn7kqSRUbFWRtSZLR0bIcns/Jef
UjVbeBZj//yPztFzcmTRA/vCCYvPflKWfTAXtkh0amtreR2diJArS1OHmVD0qs1/
WmTyk5gHWwOjY/U/EcXUMehGm9mkZZi77/SUgeA71znzxL4JgBOeBNNX957SYK4v
6LAs9UyQ8DzeDuCCrLeTBEQsMi5brWsQ3EI74KdfSIm3w8NFsh4X3THCu6l64hhq
SsnyBqp37lul9DJ8ZjCWUvt2HGF4x1u1aKavKLoGFIH4KulOS2Tdz9dh0QOoq6v4
61kHUFSXy2ey/nftZ9cST2NxN1MXjcBzh7h5YP4joct1v1G5s496LTs2AZpthQS4
Oqk3Lr6E9cOPIwo7Jk4uarz+4Ar0r0g0KmBaTolOVgURrg57Hu0wCIUiae2Xq+kr
jxA9lbwh4tWGhFXNnT7KzG4cjL2xGMXtT2LD8i+38fdSqZPpwdmq7LjlbmTI3b7A
iDxUIeUYv9kvgm5jB00QZueBlhu8T2GIMmgTvY188SoL06EzuYwoDnkXb43LfLnh
mlrcG7t3j+7NbIkajhPUL7sJLguYU4fp9iwWzfnMpSBbRGmAjSK6G3lWxCYiwdem
Sba6R/l4tywa+ZInaxHtQOnAKldQNGLdZae+RyswTWglZtnBnCuibOm65a4c1TqY
fQrj+GTkrj7Y3h9mjh6BmUPR+9RfetEf3WeugeEd1QzFOwVRwf44qDbXek59kvnp
fPGDu6nBLX12AaLkZZOkr+9NOKpIFZ78wNdFXen+/TMFkK7TKUqupx83BarrT42g
vr0hoYAlLu4KxSnK/mIas90hfa5rOpFEKI2hfGv3ZFZrNANjxgcJa386LMxP66yx
vi2hOop5dAoBLaFvmGvCWYg5JPXjr7jEsMLNwDVGOhrckaU+ogm6dd9oO2Mal5/Q
s/FGKtTjrwinacencMWpRMi+SkKw+X19vbtKi4EuBUlV/odpz+flMZ8LtkkTcO04
XjMowq7tpY6zKRlXfdhMKuiKkNEU75pMcYqBwyEgo1PpOL0opfHtIm7w3W7ZNXua
9gol7PzMUKFEYoswk6NKOTxV93zBk2IX3lECbv9C3ljbMxJSo2mEaFUpwtmLArVh
wU5LECYmu1cyC7I84nSmGeqpyzWfRIn9V3vafiqFlzGX3VGBa6f5xbZnZmbNWSgG
CXi0ZeZoGxFkbRmllJ2JLknQPU8AzxC0JPneZbZ9GyyuASv09vjqXwDNUW+4ie3p
XRWQ/itIvwJhbO3uUvEZDf1w3zTHvUCOItOkXUAzyr2yHaPZwkU59IC33R5VSvgp
fd1QqqWCcS0lxb5iTJS4kGY4we0A2j2sNo6MQRw/v6akZQBKuBREy+jkK8RsD2Qs
kEDPmgJ16bWnCeqaLrAmOn3yiQnYaUXpwuCEmCipqQRal1cZOX3vx6dMRXHIheo3
y9DIuMzYbQtlWrltRkFHr24vTJ5loY/SvCDdgA/wMFA8dk4tR2kodcJoBrZ/r6oC
o8D253rBvVbGNrLusHisbgcJn+xLs0EWkCcoZqSvgyjFrS+xQgbbyeCO404wUua/
K9zpCaL+K50juuD+RADrGmfoxTjwEcw9a1SohbUp5RAMKU376jnUdUE6q8Gu1l7Y
ZeuBgeGUIrATb+BQ+rV6ahOfS7wv5ldqp5+dVWnJum11woVXai+OCl7XEFYkRTgh
CkDesJsD78XOBDZlrLrwD+8ZMSQxK2LfWjCeXV7n3hhjGxJsfgDZ6BseuMxSkYBr
0cxyWFO+loMifIRAHwtrjrEZpsW58rRtms2kyM7jN9vz0qXKslQyP5SIix3k7FcW
3Zq610IeogQR10J8kit0xunhFQWuJgQkazeM1zYCxfThj8wF1JAuQ6ZFnGQA+/lm
kd1Y2qyZZ2MQhTG7JSh34NmQYoJ7EBj2Q46h6KV0/ra3ElAE+Z6OAxCLe+TTvL4k
SgmQKcK0vljWnR2QX3H/npwbrT0w2SaERwHHdRnD1IMg5JOedvXkWdtzIi2upxUY
KWptmvuDprKs5Oo8xpSn73wFVM13bCwq1Sq/Kkmx+5Y=
`protect END_PROTECTED
