`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDiP6jA7G8lFHPBFX9OtlCcAEbchQbg8oTK/k2Kdxfat
p3+79989svglFWvF0djQWS/ZmXdhWGp6dwJSsggrq6WIS+may3cBGp1+6uOHw5HP
OEESUiA7lLN/lR0tAjtsAUj2CiQW6xycKQPkgrXfc8vci2nVbRSrkzYXXtunQSMk
9nDTh4eWN17UmSo+HPN0xPkabSHMMcl4No83zUsGEgroWmg8Fd9ce/wqXm72p2cK
yhpbsmXcRVUcb+zDgQ8iLqJFwjv3XVE/inr73bFvqxCbuocW4egWbUQ5JU54ENhc
d6+qGzNf/XUHsbJkbtIYGXVPTZXzUVoQ8X6b/QrNMWLb7LDKLshhyfQQ5HCEJ1/F
l03ZSzJGE+7dZaeOEDvqh6dxrwOGPNHtQooGS9VWbaSrS5i4OgkQD6XycMcVM/76
MT+BoD/xeqGBbJ2KbuCBujFZr5wYyUCpK2uScd4ScbPCETzInjEKtU81LLf8a9Vk
BOv/SpeteqVSI6mV7L2dt+QoJO90yTtsCixWkqADJEqudUijjGV5CXNxrWo+504C
b+4Ftl7CTyJsRRzlI/YAYco54dRwYmo6iDk2Bz5mBFLr/t178lzjsPgFkd/Gr9zr
wAIBs3qpDpV2gcA0+vx9H0p7t7g1bEOvsMDYgLxoD4SVonY5+/gTnC8bYUVbdlmo
PmVisygQYf7nQDktd3CWhHpLR0WJpppHkyutgoDD0n+PkNriiEfXpktTIxhGXfhy
mNkK0cqoDF3ziEnxn18tM8Jrzp+clElSRvPxvAw4BtmbUcBx5B4i8gosnZW+E5u/
LYgQQ4RgrixXfMHOPxLh1wKg3Sz2v0cAe09QQYV8uIg=
`protect END_PROTECTED
