`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42W4HL7DXC5haKjjdm4Z1PpJ0przEXJ3J8D9jfCDep0U
T18xixbg9LB+x64FnQk5dZ+utBCyy8gGkKL1r1YJ++AByMpPylsB/bFhaoJ41SIs
p43lFChzBGompJovJkRBfa0VN20hgdriyh4DAWRYuR85+MQffjjGHmpBWLvYc4VO
WJ0P7MCcMS7rtUb37a2izRDXZ0DsmwWXeBxq6KofT0kILJz3kOWCjI2JAudJtzBe
G2mcQZ6LPBd55hIjV6cVJAFAyn47x0JNTyiU66ed+jNWN0BpwtGducIa1ukrajM1
6MlAczlCite6wMmngvJFRA==
`protect END_PROTECTED
