`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
E6E1iIhcb3E80aTtq92MsNp7zJpaCp5flGZcLERn9SXInW3WRfsYkSzoTA0hymno
+BZjnFYfYCraD0+S2dbCuJDver7HJ2mpF8m9YrdO1IGWiEIRdClFBgLsPWmYSgbB
XvqQZWvyeuATmC2za939nbKOhIc1WMZZm4R8URyLqKtVHauVo3xjegw8ECpLu0bs
k7HOwHaQUJhSWTuiX2DDJsLR8GcMEYEQYqoNife/gz8=
`protect END_PROTECTED
