`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bY5En+hAb4o0+9RgxYkBc/lS/GBWg3jG6lbbA1nREGkCvmzbHp8yFjhk4ZMO3Iae
34UxgkJ8dBKdxUgb33stt04KjjHAvS5JB33EDHN6DXKAx170JYD3sUAa9cFlFPMx
fEE2XSzkLNchPHyqANwNssFYLNiwOxirwGM2HiyDzMM+Yiu+d4kck48qQke4izl+
dWmXYgiUmdzhqy3y/NcgsaK+GMBEc2t9gx7eqvSm1ULwn2G7/dlnqNDkZVgI3nUB
32PQDiqPNLBYlNljAbdm9tgxe8PFPt+HTrYDf0z8Ck+4YBqi1y1sJ/NintAMP2xH
5YQmSlW6GuEMIwriua9OQFvFptjMhqP9BpBxeSz1D5o=
`protect END_PROTECTED
