`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOc8qigpl8tEe54zBvvbvfWPCzLtWtzKP3IosvrfrLL/
IyFAjFZVqMpzD8J612oqQ/fNlIVqcPc1Z03nKUbQwaKckbAURe4K9NODhS5QP4/J
ESHH8Udp5QRf4rty+QkKxqa4pODaRbHqK4iIUJZT3SxURd2tOsEgLUlKVrs3P2Tc
T9OgBprAluDu/TCcUponTYiT27+eCLc+mc0F8HjTMB9uwlDuMvS06CvDFTTZOsAx
URy/PqCUcYqbWceBt1BJmG8QV1Obzs5HLNf2sXIMILlZvrwbsLXfWJF8GopXxg/5
9ACXaEO6e2vidoM+Bg3SQjWk4lfBaISZithrBxul+oTPkwMSX2FQTdrZPfEEai9e
pVamzYLsGjNopqjj48Otiju/ZltVLsFau99vcr5gyafbUks+oMZcPw435QHRB4yB
nB2GrIBKQFpfcTLDVT89/bxsmzT9eVWk6yF6xIz16RAquMKWH13ao0mS6/ndIz+j
JC2ycOoyZx3Cg8COjYQ3GCnVw1tGh0XDbv/cR4F0sz2uddf70Un57gm38gmtzT4t
zUzw8E9DljiFzQsbRsLdcA==
`protect END_PROTECTED
