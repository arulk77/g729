`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFra+XZfZuscL67H9okrA3mTUS6t7pnRrcWYCYiNaZbZ
SP/fDG/cwmQVrbchjHeK7aoMJeX8QEJbh+ki6z+K4eW86c8Qqu+dUQx9eBaSBlhx
Un2R7GYBXOG5X98xhRPZSC3ePvS4BU9gFlM4U36z9X+PnXUxq5hQ78RQluxk8ZJ+
YePQJu68deBUx5BuCAE5IJ+0kIkV+9MxtroEb/fkp4arlEsRBcR4ACFcMhq/Hp5A
U6M1ecw2icPtaVzo+QsDoVkvNAN7dvt+oKUnH3j/7KPrt3SXvy5WrFHt/FJf1GwD
O5RqOM2zQQLAVnnuLY1R5g==
`protect END_PROTECTED
