`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBZMHhDbU5rR1qzLcIGRReIaMm8Ftu/0AOqyY442r8ca
zrYZEa0oUTp5Ltrr0Xd2VyhWNHrEm/ytQhFgxZT/tWqyi4LeMvvg3BYV09mBDvVi
2xekQLyDBPGkWbmkZTKIx0NrZo3xjNk3MqIc8JbqJsnS5OjcJSJ45mNW/q71fYsA
DkDK4WJNBlDnwPGtdwmJTw==
`protect END_PROTECTED
