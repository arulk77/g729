`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLMNu/EqeTDYS0XVPSC2Ujm4GUGLEGdYli1+LjhMySea
Qi3iWGsx7lkNXj0kRnya5uvu0qmLJghPM1/R4hvDsv0Ag7uV5/sApAjNiqT/5OXT
C/BsmgBmLyaR4bGiUlvkn8qS7X83Zxa0iA1lMKpBtazgHDdDo1Zo8tOhG0z6MFFd
N07jt5kUFcHHED4lQGKtT7XOs5aOqXMexqi6MG4+HsMSHzarzPMFfqIB1tLRxRi4
i5rGQz80oYu4vtnwDnZo3QMsqPwVPpFMbVNxmR9dJTrgN8kvgRxPZc2Aprj/FOQi
eb9sxlnmmT2vXIs5OrGDgDok6eGCo0w6/LhnXVerdcI6mYwszYVOPFB/XiHmaTDn
Zl/GLfYk5jKxngs4b0Prmw==
`protect END_PROTECTED
