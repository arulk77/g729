`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xS+mB2blxWJqvuV3Da8PYxok3NlRs0O293h+CTRGp1n
i8z90GxfdgLskDf4keJgZz3eYyI9T55IZ+mUkk/MqKz2rTDcy1i6GMKWRkf2zS++
suTGW4E/yEnZPoUEZxgh8UTYbVW6PlmAAag7HX3t6cxNTdEmno0tHgRbTupN9fPJ
/Mn/ZHAm9j+0GGT3lAE2kPGkpHGD4erFbxbbCpfPVXTSXteO4pCnS8vbV5vt8tYf
IEdcfFmSCQMHfa3s2uXImspUBoxCqUT6UWX6ZB4e21Y=
`protect END_PROTECTED
