`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
5+fw2ufX/PDi8aZmV4KbEdZZLNmiPmIHUQm4nrODn3fYA63EIYBR1qw46FeoRfXn
4s+IqaphUAwi5yoUCG+d9JYQwE5jmXfTlBPMJeMVZhGbd2fsYlnb7mgzGHvKhhKN
iYsxPTegH+Vb8RWeD4C7dqX19yUXI1rT5uc6H7IRMqyuDoHowlEof4jJxALWaq8p
FRcXcTfQm9Lb6k2Lk8pGUFmv4JtvRD66X8aV6IU/djmOdYey1aVVM12q/esD34UF
cgmVNvbpa6NUqs6SBVgr8tnn5vt0+pmTi6veBr2rUEPF2FERf6oTUOBXYqlfK2Ti
rSrgShtGICVlJzMQbCCDT2byP5hadVKkQqrWne74p/5gnCzNYInRDgaqUp/YlMZC
ltAHN0zu0AVmjeatjvfCApZiA2yqz4l8Xnr7h2oTgBq/5u9OUGFzXPX/cOVJ+Va/
OakLzrGLHaQ91BBjei3rZKxAyqARNJJcly67un4Y0iaRC+/TcoMQs6AGia8S8mj+
Aml1Qb5lecer7dtLB2OSPOcNeQp0mwtuZwTXr9wP6u0=
`protect END_PROTECTED
