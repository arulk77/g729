`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
if7OW3neLerq5QTb0GME93TVVYdTk/nR3kkMz2CrTmUdOavJWLu5iZAw98fii6nB
8pnsKNhtnW+8vAW+QBWvKnh6S8wuW/PCkXyUDgqDkuP7oqo4ZnZznkY5hP0sQ9Ov
mkh2jLoCNNrkBWJjwhjwS4Ei8SceEM309SwMWQaxjhkmIACqd1XqTBBigxafW4ke
oLfFS8Pbgt5I114fvV2KPdg1X2dlsLjOqKFcS4/qJGPXkuONYbLrGXzzEM3sJ7e+
`protect END_PROTECTED
