`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEklOXSqxxD4JSG3oLfILHo7x46oPCkHqDuy55PcrAEb
TN65/K7GRMpG44N+Lxmq7+jI8lapgW3al0VtdVfm+BzLfuj8Em1nqgfnYyNHWlQT
4zJRJ1o4XjiJDTp1TXmS3lZIXSL0cOc5wHttN86OrTgtciw2Q+yGXjtDgiyWNWEI
Ry0LUWygUPMUPrdviSwYwGQzCkY651Eh5VLbrBnnsTXo4W+e0ROJtDlLvzzaFY2w
BzWwafpKqZwAGqIFHqMNx/J/CTAOf6cxlXdouZxDI6H5EIXbkn7ifXmK5deFSvRJ
`protect END_PROTECTED
