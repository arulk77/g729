`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAy+8EqZbz7auDHkJ/eCVHLbGeLaHnhsilwJXUxH9UDx
BwC8ur5zhL3WPOXjLitM/ch66BczbKwQJw8Nv4dXOnGxJ/6tUdAFC5ivsUTCP1Zj
WNlt+3AEs/N/MIJKMVSiDe5dbONSPmF/RlQNDXkgCPFBDgsJT8lKpBE7s0BnW1Cy
vPijb8cbhsr8W0QJOQvMaD6BT26t+DOr4emwCRyYIwJGjfOGF68eWMAGzmgvfI+9
`protect END_PROTECTED
