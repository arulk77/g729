`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44BphSFs/+JJVxUHG/Wxoynifvj4oVns+ortf/jvRhb9
Hmfmo8soJf6KB74IArvE1JDleqCGL3xp92SkMI7cwDUbAP4YybqhRUO/FLZRvu8S
4vReBImkdyrC4wLHJfJA/7/KIboiu8Yd/14oBwCF0O5W3Aj9BvSvpKgtr3YNGDrX
cGaqF4inaAq6wPMPfx94aQ==
`protect END_PROTECTED
