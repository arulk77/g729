`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJRDY+W+L5STAhQtzc/bluoAGC5KKlY9gywnpHlmERqN
u9jnNa9zgMasbIM/CbKTZTs3l8HSgMakTJHUCcfgZUcGv0YlSnv4pIHUV3vLTfRJ
ziFIBybB0C3BpQiJor04g4KojisgYfQub5RWRspyS37NwUs07xw4jOAZW3FmY+GE
kgCX69NIr4Zu0TVd6eXdjsstTmpO2PEq5mjrL5k8kuko53BtMn+kmoKqvu9h7MbB
0/JI/bh2DQ5x2WXz1fldnYuTNgZ1QdCk8YOQzlGnLVJ9G3STJ2T2F+AUFYakRa0f
rEunbp0GjiYLcSIzbQxnHv+ZL9lr7zMA8RwMrCtO9NDjrwkl4nnKYAvJ23twdBZn
`protect END_PROTECTED
