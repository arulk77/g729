`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C710svjsiC/cyMPC9/xXb+EuTZZbNf9lHondu9X+YEGX
IhMkULOxyU66GhA6W+51n43sxN7pdKN+Q+goIiUafdL9BkoAeBVCGWNi1AbeIJ08
rAhOtFVx3VgbnWQ5URMCAvvA+K4TiQgX/J21Q5yPdjPf45w+bHdGXyop3b/CnSTZ
4VEwxAVLakBQJUcOGvrsC0OzwIRUFhVZUw7MP2dZbpOASpgeOgIYn7JRWvQXuqmh
4KEMN2tN+lJSqefowDQJwr3JGWEv/YSszhSKXcDPzNRytKlUNcHdIrnU3Y31XbNb
ZUNaH/RLOlETwFjBTcsgWQwGcP+3JwdE/l/gXXqyKm9PrieVGHJklFyepHj9Cwgr
yYfPfOZdZeakr6z9F6/TJTDBt/jPKtt/HmFQdf9n8eNc+LwzR0XxqCtCN9pwshRd
H4KvfIaLnWUaeG9JtrZJxzyCAJ6r3+mOaKVmwNkMNK0n2I6LCfXgFLm1aEbrMOOK
rjRuO3kgOK3jJiOpnKU25HFcIW0gF4jNSQHPI7MLBfCQkfqUKH8bRwvKy0FltdpG
TQdMhmk38GTewyozerxeK+Cq2JgR7Y6wwJhZfddSvwJa6xKuq8dmldvFvJhrp8fB
LSUHMKEeU6azaJch5use923sIcpKWxnBFTwb3RWZgcXwcW07A7lXHOfDWHDWpST9
5mW1fyx5F7geFzse9J6T5g==
`protect END_PROTECTED
