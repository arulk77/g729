`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
WdYtQaMEMviVfvde8jxk8Eybbkx/IEek8d5iXxPByOy+QKoSuGviXGocw7R78ZXp
oQDjxcri4yeLPvjFDes/rc1Ua8hJixlDm76ceGB4JKk1sWxn3c0FVoixfhbtMhsb
WuYCdNMNHamZbVOcyZi5pG6Wbtd3znsm5KEABBXYBk12OGJ50YDkj2wej0JjSwF7
ozCIGzBrZSux0SLWkyiRLMX1zvZ+m/6vl+dRU6qiKH5kBoyK9/FBnZKud84IW/ll
mFHGj880v03ztgRxDzewpGq7JFEAq9SLbplnpkcQlKi7Vw2izyrXfTRlvypubQBv
CuQkG6mUM9FMeIhIBDt2etUp40kbAwiIWTC6xSB8Wpw=
`protect END_PROTECTED
