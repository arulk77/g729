`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF0yh3zbhPySj4KxgSrezfxYLW3kjQxRTEmgYaQTz3j8
jKLRQujBw8uQwbA09bouONigftw5JNGb6voIQwumdf/RfGCpRs5gbw2/h77EMety
9LSOZfkrTQV7Y/EzsptI56FTrxxazkK+3aX8Jm0hyIXJcCH5IOYYzBvZABrL5OL9
E7QAR/NRHySk9zhljzy9+xhaqJkceJZo13b2fNsLj4sg98+yq6CyXVXRHv+BUc3q
blTeQPe0QXhAOk+JfxEB7oqQ/EbS2KLQI/fY24Bknqipvv5YohzNId5VNJwI0RAy
0g0gKp7AsW6E0hnrPO0+L89h/pUM0btrtvj8SMuhXJ/+VKmi7XluYlnG3IbiBY68
uOI4k4xVJM+2aqWaZDVwlqXjosBMNFmf0ZYWCKrNV5RsAtgMXHMQwH1otf7+UQpK
tH7Jx/y0VmS1S4b82KMqApBc4mI61nLno9ZUsVY2LQlloZ/ihsmP0RbeM+7Ms6vp
KLcXy2RZs6rMag3OcADZ/lK+qRaKeHtQiW+n5kfK50sXTUTUqF/UmPdvcpoLfFQQ
PaL2yOIyQnu3MmRb6RlFnDk7QoEnYwq9ZCBH0gwK23zLfHfnXiTct4/5qbgzs2xX
fTFbXUlXFTnzopPuSBixjYvDVp9Aj5ddqhogZrmo22ftmiA/TfL/VjGVFq4kVgXh
lwMjtPKq5mL3IXa33FRTRxzEEp/OeKdysYfT0ZVekSE31dwPj1JLoTsm7SrGF47M
MhqrWNxULKolcq08dBnfTrJjckpIvScw0sjq/LbYRoQ=
`protect END_PROTECTED
