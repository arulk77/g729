`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN8utsj+AWXAwbfyrtLgcc0gjnrWiHjZ8c93RHJ2Wr1f
osxwEoInMU+TYPWTmx2ETNr9fZf0ELXI4F20oSXgN7EpWx2JjMJwh2QuocIPtug3
DmucpZVQiDxJJrjhbpPTsPTTh50o49NO7wOUBH/P3rS9IlwdyhE+nMt4YD3QVOtD
`protect END_PROTECTED
