`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
niIVou0AAt0vRfZnOa98IsMdccCcYBlHcdPnrd6TwVeB6XLIqrambYittgW/YQZj
/eVABYzPiEAGCwk5RK/gPXQVzCNL/ICornYYQhhhqljWu7Cxxago+O0/qmP/F464
OOVZ4QnG28dvQ372u8UYOrWhB4hCa1yKR2GrnamIp796pSgZoXEJJ+7TYJ24gYRE
mTHtglIucO2nRm4HpM5rp/loZakTB1nPLC6PWO//0oeu9WYWvdBj1uUJcsrXrg4Y
VfWCtqVOTRQ2EULSDFsaIn/IRUJyh5EKgaR0pdNAG40=
`protect END_PROTECTED
