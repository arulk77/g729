`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAaE2uCWbAy5NGfc3pIoj5LFIOGaZ712pPdCM3SWb5Qc
RT7OdSAGHiX0OcvzsmUfL9/GluFj6Rboew7bDHWJ7Vp4Q2d49bY/hJPYvRpbw95n
vY81hS6mvjnBjM81NyTLRA0E8cWW5ZxL8GcX8AHWjTdnkKMkKODdhTlzPed/pyQM
Za6CfCx0Hi0fEEYMHixuJ3dpFfmK3O8h1Agi8TUT04J0e0JvO2Ngu0jREHkdg0Dc
fh1gzBYbQKFrWv7tfvhpHA1l0W0TMAX8SUx8tWwKgGS+TovlZyPhs14b8PrNOB7S
FSMdx4Cl5vwb3PKK58phx+15Ij1YaHopjzOoFSTuAA9xT0s8r3LkFHT5FZo2v7Vg
t9RJ89Z2AIffzlP/y8U6qBG+02m17t6CEDLlHBUH4JP88Nj+IZqGWK29df6JmVZW
fJGWY0R+Kg958C8RCdjxdT/HzWHzPXH/5cmHMHNAHZDhPm6mChxSEjSajUoIC7dz
Giu62gcaY7iX/qcDEA2uLN9B+X49psZcq9s0iANOVQYXo29KtzAmSFx72wBBBaTG
vRipAHCp9TRnf999aDsqAaKL/izHMqIgJCTaJKFzPcCTfxe2S+K1h/ZzDY7jfvzh
TtCPjFr2SlXzV8T7tcstsPuHCkiwKhKLsUeZV/CEpeJUbmqfYARSjnakRvLJkQ2J
QNwUJgafH7uJyiEXBqwJd742OSiyIalt3qsxGKEjowEM1W2lvS6wbN+eQkk08IAa
4192exxfbr8u+yhcJH3Bae0gl7K7F7pPSLz/PGY0r4Cm0O+BJ/pNA3t0e1NjWOYU
o0eWWPqrkGT6KveaL+hUE9ekl2sbg/nIo/SJHEEHMD1fN7C4pZvUuBhtdnu+77zA
EN6b1Tx8ZQRB1lUMMnmD06mNgp3oYqQ016BpkO+dCmUYKs0CgFGLhHX1RKmvS+TU
wUJSqHk6XKW7FjG5ZkxUcy+mB1i7HHbuVCGISVJwzVmUqjDeRkxZ3CutTbgmll80
`protect END_PROTECTED
