`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMjGnkW21yuSYRiK37Z2KG1n+Z1q65diaPzcgDp3bCle
axXW0v3Jjz57QUiuKCNXzfsnA2lT9ejqZkoGpbSmpQpPm7hRGAb5zWc6YZjFEkeu
IC1QudcOOozR4FR+PBPwuQzVLuN63PgkOyNWXrCNK8hZs9TwdzbtIqc5S3YYB1K+
3SjQzkQHAFDTdEUi2LEyLnnGJKFmPw8a1ENC4X2GgM1mXxBr9hnoF/GbH6Ai3ift
okF99BMjuXRYF98MXbJZK831fJeYt4tJW5jP/ZNT1F9XvlIQYFr4Z3vhoQ1QrmRO
0AFLFMaqE1zhVwcVVpPYrCVU+3yrcMW1eUb8w2hdsBiAe4BRCHsyunzUSwyrt1nj
Ogx1pmLy6gIOCRWUj2OZ5zgnmcHYiv85JHyGSp7s1uhmFdnrRbMa/XNyHjADXFr1
rk0OCLeGNQBBxqLws6U5Ru4Mlg5TAXotdn4A+51w9+tmV2PORCrBZw8uc7gTnM6D
g0HW9hXkESmyJdVEc2pnQbrGwjcQOuhuFtDzZg1m0QMS++bPxjrf13hJH5sKw5cN
R+o5svKh2ZpKD2PsPijFxUAq1ORF+KV6/obkiRLRi2fBK0cLFloN4ZhZ3wVu4A/E
5OB2yv0Ncx8Ozcdmayz2wIfGg6uhgEjNNGP6aGPcN5QCsuIXVTuWRXtVprmhb+de
`protect END_PROTECTED
