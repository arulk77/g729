`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDARWpjELK6yxXLRNdZdYX70jykqn2n2MAF+/JicYUgIcB
nAl93ohmyycP+cYTqSPlqOoSt2AfojN5VjdO97NLqzgW11VDf0xHd0zVXPflPkhK
sBwiUmdxcUZfbO/3KmC+QKMyQEDixNVZmBB+G2YJLX2SGF25OwtPvMLgZZrx5B/L
xo4H1PZDpsmu6w78KsrfA4oKDeSqtmJ4qtydcVXdIMGb3IFRaaNekaCHsKlgLkhH
yBIxl+qykFkVISkpCFiO+501/gGngyE6AwTjy7mh2nANGTiMb05pfjDidNkUaL+M
GX1KycRZZ94A+rxTof1JZ1U+R52gDH5WXmjK4B7yZB/kDuSK+/BJL3KwNRtMW7uz
jBjhHOvoe5mEdiUohmmEMrjwF080d8EcDq2q7AamwqeYzWYIHTsxf/WJHUKsM35R
w2dMPpQ/SPgBsSQ6jENjHs3WRpBYO5qro1nd1VO1TGJH+NJ+oTQXlXXLn6Co9aRW
RoRN09XzvLdnYKZA9o9wzQOSrlRtl/u/pXpi3IapsLkE3D39Bie4rN6JpnkqavjI
sBrmIbje92XSbXGoLnYUZLK/2vAc2bs1jzPkv0faOsVVbbC8utet2WsnL3PRnzGq
7uKiYrnu5AjjC6PLdZB7zcAPm/WKYn2FzDHrXYoFWmVu9i+8D+98oGLwL3q9kuRk
OBvLhI6rm1voXMwSPyrxviS7CLVLgNdcOweVq9OosJvf+jtvwmA9y/nuiPz8ZDyM
bIOb6tQUhDPmvqfGMiIfQUC45538QD9DQhsGzxLQfTmOeRDP2Im90S/RzkENPE5p
JB2oft86VQ1YkwKNFoJtFwFQBg5gWdlIR1GWRzqEYtM3pdwJiSOg4ZrWlC7qIJBh
+iwsbGZuGErIa/UyhqJQQHJuL6k3wjtsXtQYCPsk1LHYweK7uCw+nJOBn6bYuLkf
hgA8BzBCwly+4cZrBlion6gigSfD7TFoCs3h2glHWhqeDjHazksBaQzsYzUBrn5r
iMxNix4tEgo/4r6z1ztWG/5AkUCIHl8VdP25G6QOAiiebnLMu7t8hKoGOW+Mfkjy
+6l83fLgtrP0ZXaDzLrR70ZzdRAnD/FB1K5wK/re4csEVDF+yDgu+8YHOAPi0NEW
LVZrd5xRTqr3VUpKgdCnM/WAFHWgcpLy8sEI1uBethMZSomAm59qWQ6twMzqMDGE
`protect END_PROTECTED
