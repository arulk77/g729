`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHT/yukZomR91UCnSczOJAKgJjYgzxNOQQ6IGHjM+ZqO
+cUDe220H26OBBEgB2y+JHEyJK2rXkyaF+armfoJqPVjT5B2/BCA4pJMO/fIIdKP
+hYjXRrrv+ktrn9CmcSaCZmHC7K1WaxqPft26Qy+aV1kpyhj2QQSE8itVj4i2MSL
Oe1uYYL1fKX0ck49c1ScAhhhS5EPSeY/K5jWGgm8lXckdss3l962CQOaWE/zxnvE
PHBUVPQXAkWzJ5iJrnj1NJqRlN0cfcnDWgEAxZ1fyNhQMdFPMQOzOZsI5WjNkCF5
p5wNXFdrQ4xgIIweV/yQM5l9Be+iwNypOFSZ6dFr5nrbbK6wQ3lx8mCP3J/akfUs
hD0RK7Y5zQqR8N5VsqY/YKeGwOp7YteVOkXlOxlIaAbI/eMOQRdUZuUUes8akk5u
1w6mKPcIHV+62HIcRVi4NfS6rGuZy8BSJDT/+Q0F6DdDiTykUAayhd3U2G9UhgJW
QYmue7CNgHMjHEq2Dk+yCG3WCRbrH6CakstlKlGeGmNqPGWnBP0yZCY5xpeubwsm
`protect END_PROTECTED
