`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
R4XVF3TkhtcHz4A2h54rdljtZ7not6+EbjFlPm3zYIXOcY/5B75b0s9gaN1TZgro
BQGx08oD8x7pmYAaRUi4ddfDWyxgYQU1eAld9z9JiU6JIdFao/vktjkvgYRWXNNz
yxJOLxL0vbLaF8aN+t5uPB9vYh/RARLALKKsONqZ7tQXYGJksSf8pvH1o/BmPlMI
WfYbktQ/2JPrR2Nn9QViFwUfi1a2LlCi2SooceRBuLI=
`protect END_PROTECTED
