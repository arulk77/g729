`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIqLH0tC215bVS9GOnphHQsy8LHF2aFneHnwdpfkBNtj
/m/VuGgGtQlbkzaUONjiSfibq4GJN1QsV0AmG1MfE8QryYeF0Z3cy9iIadwH+WKy
ybyDxaH2L7x0q/mc6Yt2D8rRWimanaEvBryTYJmViqg5j5d4irXgCdw4BosF8XiE
CoEG+gINPV5t5geh1MY/pw==
`protect END_PROTECTED
