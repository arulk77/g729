`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB0fK6JUfXC14ll/lvX2rLswzNsZgUXfSnGlE6eu7QRG
CpJ5OlYf1KcTTBVI6OIs7RlqfuYZWG6o3A+6DPuKx3R1quUDgoe4xPImA7XvfBjG
NRDmg/UZlfLIJ6lnb2OtTsOj7CklhalJN7A4DRPSg4JBa6YYzCjTcsLFXpevu1pG
DGEnArud1OyE0SP6bS63J8sTn+vdKxCRgUtRtFUEyjYTLauewCosIf7by9oY4z7I
xjl7EdgSUFCIao65jGiYU5h40rwUTRxJ1cY2b0MPZ6/o8qm4Q22e++yXES1pMf20
G+Po/TERl5/n2R36f1aQXcUALmFDWiy66WlP9btE4ciRPG4mjlzOtEylgP3Ac/R8
P2YKztn9AYwI4zthmYGbUfj3w2fsv8DCTaAIejrUDIBuQtwn5YTDR+ynyiLvxcEJ
`protect END_PROTECTED
