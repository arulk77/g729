`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIGDrEI0H7L3pGZkxxho8kx5A0c3w9H0mm5kUoAgcsb6
JFFSet0QxR2a/yM8KIu59zykDOuJC14JhqHw4BtDxoppYcfjqgHsdjlT1GoqNCVB
LHR0sChsVIAIxQqqICjguAJhRdry4n0GI8tLkAg8DPscqIPj6m5eP2+QfTXRiRll
ycGi/N+QAoGmY+g5TjSGbAfUOdrnGe9emXZv64xLu8vVG8WDe7I4eHSqXoEekWMO
DS8xDk4oEOFmS54J7sdTnLe2j+JpxC28Gg5gQXhwLFrM+JIbZs2dLuPSZzsEXvRv
otzg7WiUkN8OXvwyoG80DAxqgShTW4tqwQ7XAC7+mdsdot1BbHfLm4qco0tHMmaf
`protect END_PROTECTED
