`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Ulcm6poJPW7dyMU/oxOw9yDIG5q4MvaiRKj4WK5J1Gz7EcqA0YsG46Sehu2+Rg9I
QS3+I493X3GrFw4PcDYe/c8nYsAn2Bwl61sotuApaXnrLSu+ijjo0wFP02iofMaA
39wdvVWy3vmr0KUV7s28cVdpB3SSHPQyxa1/s+nChOzy9idDxA/fJD0Og8Pi7cUp
8fzcPOJ6pJcOGoEFYjdbyTR68qn8jtSz1ffokIjBctUeZiEz8W5Xr1F2Zc+Fbpeh
LGLr2G37A6vMFt9iy+4vpOZ6zOIbQyfRkx5utuuN9c4msNbH+L8Rwmf+RfXnqUj4
7he1Te9fPx5q69A7wNtEpPGcHz1/CpIt4r/KCX3GMga/oCd//UDB/CAfgS/Uph7y
oJVUv4iXTKZzNaZOKS8x+nkcFZoMn5gKgEex3ByvzTL5hBtWg+7Fu6ewtd+mO3ct
Frw23rM5x87FH18tZIGKGBOd7/ltv9dd7BrNFMlOnucP0syFJuRYm9m8uOvhMCBp
OolWgCGyucPBa+Dw+cCp//a3YAAtL9PrMAtT0gcUYo0L0NrUTG0SEcR8osfQyHSQ
q37ivaJLJcnxdJEZwkD0M1IWvukC3ocxdUFr3gLMqz4FKXuXDE1s9nlFAkpF45sk
zGXR/ww1VZlXrBc0SrXlSzaTyelaF19S13y8nkyeVcB3RGeolXvMn2nevCh5oA77
nNU435ORDlMl6Bn3p3ekQJNRVARZwY4MNiBQ0vATMTa0YWk4ZBeszYAiER5WpPX9
zBd16K1X1C5SO2kfHxkXonva1rZ7dJnm7M/7Zvb/ceqcrQTo2gR0eO41r1GIpSi/
Y31d6sp/CZ8bZyp/euSNBclojVRY9O/SUzr7gxo35DUEBgQAM79+WPhmpbgOaaa2
dS8I30iAnPg+nBQXOFL/sJdQfcu/EZS+uqoLgUccdyx4BgurY4ai/UQSbZqCp3Lv
AoxNqIc48949UnW3WuEB8t+2B8pZRQGfCHleLiYICUBa7UsDf3XwSDFkssgPQBm0
OwO+QFTHql6pRUDenkjVsGgtF79h2BodWetVGhCPdKDwt43/6+Hs1al5vqFPEzAd
mDR/9xjw7q22Z6/pvWFoRuBtKo3v3Mc4cMzny0B4vC2SNHeDlDEJ4j6fVv3HWT8M
`protect END_PROTECTED
