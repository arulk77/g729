`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yM+0dM83lZujxfX35+MakZpk8d0HiLUmzGfcdMWmn8O
r3E+/Pjnd2qijce5T3p9QK0Su3/HZWnGKzXITFkOm6wP+zThSIdeziFAvmi+TRrO
n9UySofQ7S00pOhBS3ea15BCHRK1bYPX1mrzqYWzyNU8tstj7jYBZ1kmPckiphPv
ryr80Ol5HmCzJFfCfqo9HJR0ZB6eYUAkMz2i4GSm9tI6B7FgU7ePfwt+Ajy3QQ+v
HIwS62cTBJ578bc/xXG/mUxVoeUxQfhdfmevugQOBvA9ZviEXjQozhXvig+Djp7n
ZQG1r9/wqekAMuUiYL5zHw==
`protect END_PROTECTED
