`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+zh/sXlLcYC9nuQb7fBMPo7E83nhpQR3TfFdZA+Bwxq
g3oGWORCAElW2Ro9tFA4mzHzYvmZqvfas27lFxYQdumnGXCyh9dR6rieVUw5yWBf
zbgQrlxRA3zmqsZWJWC9UtIw34f0EsVwPVjEqCuMjV0PPJWlZdInHC6fE87jlRRk
FpQ8Yq1jwPysNVfCwXGgcFJKOvTHC/8FGuJKiG1qGp/oAMJ2wnG85xCo2jmPG7TW
rvfCO5jZX3/kuEdAD79M3SGXnFZWpU7nggqn32LMLggLhRs9flJ2Q3JpDl1NEj8S
sVFq026PovBeOXO0xzkkfA==
`protect END_PROTECTED
