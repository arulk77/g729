`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ErcVd8iE7AzCLfsiYqiVxPRPgJAMbln7/9M6zt42AITUEXOuf+lGdvaLfTUchcXN
rgXyBIsQrbQqMvcJJYXI2zKGFof+y8hQlLNWZb++alogUjLVtotm0LYLt9y1XEYk
jXJgDuH28xPwkGDYI305KCfvw5wWs2vJEoGjSUvuAJL0MoVHvDaJ9zKwZvZ89+Vj
`protect END_PROTECTED
