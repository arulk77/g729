`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveClVFsTfqsTjD44qjU+0ZBzSPQcng/WZAQTcj2qC8XYg
tV4aQxRo35G5LFBB1YyO3xLTD13VArXRxyoC3fpVfwmydZed5WCJugJV1w0r82oH
FD/sY+UZA64zazI7xdCWYBlF2ISVMQO0hkXDtcBjV9LbdnuShbvL8pHGIBSYiD5p
gXjW6ixRcDprcvdtxFB9KYAB/YCWieypIvQKZckeOoWvOla3u9UjfgVxdHrPdouW
1wh7vftv/EA2RSPgeDvUG9a1dycEbWvncBMd54eLZIBtGQuRfUCq/QXjS1GzIL41
BVWOQZw+lEtJa29uxJ2enpEmmGPafD7vEBYKeBn9e5c3BgUx+cjCNKNKAtKdhHQH
sVi5pDvcR2MguGh/LiMA3NOAy8ouRFoEKAepJWMjR/TBGQeqCyn1FL2eS+tLvoNE
WqIJJHhxCaJ04rw18/YG4q4OFuWCMk9ru67A66/MNcsQlRSBrHVj4z1U8cav6sgQ
OfP/CbK0XsRwOpAFeTxrRmsIl3ze65nwhgdQbig/jfWw7dnzsrpwKnifwjQd/eAi
frXWaiiOpuewxNQWtbMhbmr3PfRqGsQ50h3YeI+lWh+xRyFes1Kkd6ci56Oohail
Pz6Hs3eYgqcuoVeidtI/oP+zxi+N1pqctzGZi43sQLF0g03K0/DSQhMZ5rgl2RGq
DNt9jxCct/R+9xKrUTooqEVo+SkRRmi/bqK5KkQrSSOLbTRmmLzd8KUSKagGTLov
xmLH09AraBpxunLcvHMK3vWWaA03WsiXUU2VAWE2b3YWsEvDhgVVaD7oE+FrV7vp
UgMqjTM2jCO1uMwIkIFonvfq3CGec4+RMHofZA7hdrboKJ7dfsi8hGqhrvjC2vf4
PA2D1yF2Z7Mm2NJ/HA35qfYQ85yCa0qSUw4XmVCmKETIrMK2QC8YmdOC28/mc62D
Ch3LZMCTasiA2xrcs6+XyfcYpsIjxgMK9q1c+8IthNPRxZXA++jl2eUrugxRRiuV
mNjyDb2o8nNJz5NI7rQkH9vO2ngUUpacUQPl1Gyi1DZ4xqv0gUQy/r1ZdzYeAXS2
iwXXww1GeVRnE7DYMA5xdV3Ef5V+l5tddz22s+sHGh46ArW25T3TzYYBl0iGwOIT
rZVwWoIAd8RRzcVCpRoSnLCI9D3oaGUCZc68LYjoAue7bEExSkG+tiPhnxmu4/t6
s5qb2myza3SKVbHPXZ6X0K3Tn5ESLUWNcfLkDMri0lvxpBLb+qo2XwFNdSemOd37
7WUoudkoQ9kG19x+ftsTTSMfdxNgtONv74CMhDldGNJGTNamb6/2JmCoOT36NJic
eW2wNdN0urfMo+x5Eu+u5X0570fb+5qzwXiY9zmA1KwN3Xe/pPxG9NVRYlf4BQ6K
ouuBwDyxWnOU6Zb/eWuPpdTF3PZVnxX7z2pXgmYEdfThbV9/y4voFodhiHv15MW4
KPTQNmBTWvyeUgY6hodlvmo3tqrBdHWQ/z2nNktTw95/eh4DujeTu3W9iXU3aVnt
UX9zXtuGpEK2lT8rbz9HXXwxyR+o64L5VTNWEYUq2hXFn1UFqJfh7MjN5x2UqeMT
gWlx1fcCf5ReFBX2Na7o50hjWxKBCAM3/VfB+L4jbj61jPMBgrEScMQdF1P5UQ3Y
nMshG5wYMCilooShvI9A3jt93ALp3f9A+iGFciToLVx1E2E3e0ltrY3Dk4c45D/S
`protect END_PROTECTED
