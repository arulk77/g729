`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBN0WKxUmLrXs+ORCIHVbVGelcfDlhBbhLzcKZ02Q8t5
RxmoE/s/no3u+MG4N8+Mcgn5Q7naRVltbZBD8l7aV4CiBhsD6CpdwacHS4bWzeAh
xjLHIINS96xRC0cdWigOTmFmBt2Sp2+FcZBzcidnRhA4Bhk2VD/dryeuHczNW/lD
GjG2jOoXiSMvF17vdzHz7IjqolZ8oSDDmn6iMYKTUMFt9KPl9kuGC5JoB22wKw58
CU+5i1SFGGN8DlcgSm/D/w==
`protect END_PROTECTED
