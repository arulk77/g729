`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40N6YFGheAmuQSzf4ZSngDEohUI9Cv8NIocTBLbIo/CJ
kXTsAfmkcV9E65F/1Da1EViaf6d+DgHjX13VQK6gn1pCJaKdKp4E7uj137r5SxFS
VJXZpDu4XsgpTPjidFzOguCHGEXHPiK7oBFMxEENzwfFh+NDVeUhXvzNhhguGOlx
rk5bm4aJ19Fh/bMTaRZVQhjblF8TGnNfFpDYvTDTxWDe5eD4ID9DveD1pFZSF7LA
kKLrTSx81X0uhJvymxE2y+GDHhSkNlWP5R9B9UlDm6lK4rcOn0eA454+UwIs8RT5
8/eHdT5CzkhPPHCeVd+i7vbBFAz+Px3KzDsuyiog1KgLqzwfTaFyXZaJoMsMDDp1
4GFr0CfhmFtCN9iE34oI9w==
`protect END_PROTECTED
