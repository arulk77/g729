`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
VN3cZiJB9f6xREOOK65F2r3xrK0/QkVytXdQqH97UuyDVIU+/sCCGckJgNmtG9vp
i/OWmum2RsGfQS/45qGtTNxZnQcdnqSZMgCF2Ss7MK8JhKT+A+Xaw6HOlsCxRAt4
+67ww8simTW9zuSyHsKXHI6D0rw0cholIDNQbe/uFH4WyJwNEMFl0XexTFBXnqno
rCmHODc/jOF223wJmbC+//ljR5Dxmi5jbAbolnfmUl8k8agbRN1xkfQJNWhHKQ3d
uMbIMoTxlpTnkWhdO7GEdf1qi5EfV/g48p6Ub6MizIfvKyFBm/dp3V0t2hD47txX
BAxUDtd1pcA389CARLS2q9cgZ3c1ceCiOV9awZvFUy3CuojAAj/NUVBEnRVTp8jS
CfN9jzCKd9jdQvAqOtk9F/XEWtA0NEXzbNhkUlUvWa7IoFCXN+xMYnwv4pdARxhJ
700OotPbzrXZ8mJoid/xoJCbToptFUBiAdVsQBYHtSdRQ25QuasjmzXhoCLujwZv
CS1c/8R2D07GsU0QCU8+nicEciqM77Iot6KK1JHYlOvxqb+Vn/aZUv3arggXQq/q
45Wvt5zrr1y1wLK7w6iZDsa9VLSOe6z08hMTr3iaDAVL0A+stkIr1rCWadlxR2ph
6dCurrxwCbcqjIAAZ3k7ieaJKrLjgyknCXYZ+59HZgL81xM4hVYxhMVz6ARFlfjh
jXW3yJLwz6GqoFY5fuJdOrV8myol5QbCsaPqzo/dU7JFtpFoNpZBesy/hc8EUKlT
NK80SL5YyWZpaNypdobORZo35nDV70JlNlbkN48v4FTSXOedeZA2oQd425Syz/M6
T+P3PjL30UHGkQKOza6rJW1DWoDbECbaYK5A7HKKQFXPDvaWJ3DhYAPf85d/Hg2p
sHC2yBHB6pgXosom1W4M5/0t49bwCI2dojcgm4ldqdN/iwb3HKUjktb1LmVvLVt4
nVkh4N1/vZn0/pEt69rWsTUR4LQZ89eFjMXkTmowmgw=
`protect END_PROTECTED
