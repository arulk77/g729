`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
V1m5O3Gm4c8wXl8T8mQk6jke8NPlrHMzFxzD9+6NRuAiFYjjcc1pgFUkgD/AhS1+
JI8/Xhdu277Y43X6wHM7dUaCNANvLW5oTcq+g7zd5G1a+orLfx3NntDlwrgqJyYA
m/yNCUGNEKGHY1zaM8/Gbeb5A8XhQCySKEpnDlOhuWkTsU+njdmh5R9s7oM1O2uK
tuBi1z0H8wUPpi2v73THdaEvXPeVlnBNqynBLSxuJsrk5Jtj9Cct9X59xyX407mX
QwN/8G5GK0MHajAIGQli4itAd7fPJM0RFfKTFNvflIA6ss0J5Oetw3m26P0Bo6z5
h0r+lPUvYaQ4+hxq4dQcjj1aYxCc2cbG+Kw0D/WPB8s=
`protect END_PROTECTED
