`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
EKU0KeoEu4S7LQG4xgfMseuwueTIFl/aZjZ/gFhnqirCHW+Psy5p/9RGY3/oWagB
p61Eb+EDErcc1dAtQ9RNtaeznm8kB66l6K3BP393ihpe3SHSBRqEGzgbeWKambeY
tkfZyedHxVvvAAZpN4Ju+7edX+W2+Gj8dnIDVEzSrh5ZcR5BntHfJtpqH6H6lxZ/
0NKzkScziqfvUL25AIUoKXFxImGIxrszhtoQsSnmzpIYtmjV8+iXzedh7hPMMBok
gzmmxiDEMuqnGKTCnJyGQbQnPX2PYL6fwp2qZVPL/4SkRd8Ig2Ndn7m0iNHjuth5
nL1QZoa8dkh3t46UwxukQv5Ez7DPHG951o6VV4DWeZc/mv110Zbir45jmiYJ9TfI
s8q8Uj5bGhZaT4hHguQzN8jWm7sQL2uwcansQCCLmgc=
`protect END_PROTECTED
