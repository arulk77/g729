`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47QFeX0Ww5p7Ux0yLQBJ4bdvrEMPFfHo+n5w+ywna7Ly
DrP3OSvae3dkuWeZ8D+6vVCyJKjgKsaC4/IR3QCySp5gcPIira9xuI0KQpqjidd/
6UvX/RP9l3upVvVAzNPrhS0sBxC6vWO16KFYCwhPC/8QyoG9HxfAKGVwdm7+ZSOm
WAGSoXRB8JpUVB/p1pvgh/JlI/vVByPXRv9rAP5g7Zk=
`protect END_PROTECTED
