`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xdlvtITYyoFFOIveD33PICfwBWBCgpTm6pS0tS3KL2y
UB4ZL1kln+Aa54n0QtY50Bx9Li6DDejxpAcUHViYGt9brYyodHJ2ApEPekwYjfJn
b/FnggKmryRVmbIcaneDgLtm6lfO3QANht/A/CoQO47XZwaAwKwuZpA+xIsbr11c
4qYf+mCtkG9s7ipA2SqmgoFYWz8wP7kWMiDqxiO2n3o+/r87bVhr3on1jui5+u0t
R/oXOCBe3yqKZuO+b9qHwAFWGMS4zR9tVF6o/C0kp179vyeDzd4dr/2S20a5BsjT
EhQxm9+ashIg1jX0XsUKRJ/RUFGbePI5+GbjEHhDPp+i5bQJUROUQJqwsXDeAlt+
FCsubStlvzu7CRW81zv97Q==
`protect END_PROTECTED
