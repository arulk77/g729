`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aSv6JxF8Y/OUI84srszgBHSJxBNBXEUiQaeYVV7GrKxn
uofyRE6CQRX6cqGpHe9NmL9DZXOW+N5V+BInAzOyeOfGBU9VplGhSUUQuLYn/oPM
vFxu/7Hi15YBANlRiwRtAIU3ouJjIMZyV0CWJUAdZcYV6UjHHEWo+F63cCv1Va3v
51k1Y4AfgcWcMelkWxcURDdg1VgRHYzDPRsrI51t1d+wSEXluwDhakecr+gMEiaE
u5ygAcNFshd0Ze6dvwnFWnbswdARoIj4E2Cq2grPmqI8k6quNX0+jnR1rgCJKPg7
DsXv8Q8juWhjq9TfBvG+An3jeBCIXv1sH+g6MXJkiYZBE0p3yZuGsaoj8IhxMnkg
JSprIbA5xeOwnQ5NCm1/JsJyv0NSZ2lomJizUK6X27mixU34QvFJIKpWwqeH0CeL
z1GgpNGHHpF+tmFJ6KajF2Btdx/tgGUhHmdQGiBGb3uU0GA6jwUKbJHsN1Hq/kq3
vPWvEY+WN48fogZSnOcyvxKat1fxcvecMjIjv4FTu9IZ84dAzMnuZP3TVzRFdtZ4
mbhkyzUG3zOkZ42xP5TE5akQnAGKpKItnwyi2tFDR4a2ZLHte2rsCgVrSDs46oxl
c8IFr4Bbifu/K9flbU4ilWshRuGF4ivhPwDU8tSjpsID4wAWCN1ahXWyZiTbS8ZQ
E3nW3MjqGvlKvQ1l6RdQmpXpJJ/rV8+xiDxFR5oC2OxzaNPUxjNDO3GNHfNVx6A2
AsfdupeLkNkbJIFCT3bXBGm73fXZyPka2Cb+6nWvm0qBp1SENu639Zb9r2CTOqtW
M5I92DbZLaD47WbBaV4ics8iAovlp/cubO9Dp2+IPZrBS/Oy6BktF5+riooEPDew
BSVhzch79f69Iuw3BCY6FnMmzqAlGoog6jJPpDLDtseCclSFHw2Gw9ZWQUFMeB8V
W3a0qF02WzTK8cqddkyaLU5K7b1kZ8TmKmcQOBoqTn4iqM2+pFXpbp7KkG/DPqLq
N6f/KyntNBKK5gxw1iHt/Xqc2RzvkCC7YjNT9s8dgeaf8Ag5+CNbN/18ARlAIxv0
UOocfj4oTBJHljdQ6odIz5RVyp2xkEa1SXLTeEGc10Z6DEAVypJS9DtL/Ohcd9Sq
CVg1Nz+ZQTaxZR4viJRCVLowWeBS53zuUWmpRPaCzeZxVn7Mxcpz6CzmUo4uG0SR
3dxQf/2VxPqxGSMBcBF2WnJi23MInmTzeqZzx+VF/HrN0IMC8hlVbz/X08wMFJoL
/mDeOsDDN849as3U3MmxxMuidlAHePeno1/ZYSqTfuy/qLtEDV1NhejvHmOzm/W8
U2lnK8/vsoeZ52l+2XzzjKgNDquOQIKuqSRNteWGxaPBtwaRaFZ0bFLQtRzxVjgl
XdGCPmhiSSLE7RlgJtkxQNTRGQcN7WVy20taYpq/U2USnIFSXkKoPj3npPkfH09S
L8UyYVSy5/qXzYHMox1Ryte+VaEjcMhqBpDYKp7ZuAdtijMYx8U4ILTTi4KRXj6S
eP/lmRMuDAM/lhPYQvW9urpSXhY1D1XLVvJsMzaKRPX0JUj6W72NF+PMJTqY4MxT
CQZnFOxyN8YtyGgdgmJn8xrp1ssV8n+0G06gmQ6RLVmJhTf0J9824frlCNaKJX7w
pc+LcMkiXeTlW5DBvZgXVwi9GEKgC7C5e/i02IdKkEXnH/mypOUlThCIbCcmRreh
/kOfUjVBXUVbdGrmYXQktGy+/c988nNmeT8XdeWyRIHXU2pgBk8MtrMk/siCAwJe
fix6dNQL65uvoRMvGqBldlZqZiypzkyNGEqG0CTQcGmx6TDsEB7Zn1FSFxtV5V0Q
Vzq3elaeIzOyI6zRPLuDBSKiN9lG9vuKLtlp/SpD5pQe4HlMqVoSeyBf7LdgUylG
q1VAXIMwOZEX6ra4IJNTyk0majTUAh5sDyO7YHgR/WcOp3eLyqa5PuHKzEg1YyJ7
V9YP8phV5nBWVa+kuKJTmUxnJWmjUCkKHCP5Gl6NcJ6Y2eXYmpCSkdARRJ/MpzQS
fdevfm2FNIsOgRR4led8bOu4Zdg7+xC+7w84lFsH6Xn2aVK9zcXA1UrsONmt6cYh
3Kb3kFSMB7Ezij+jieCxGeCyUSngmtnmo72KPVW2DuFbp2wtY/aG4DjZLcThwUUf
BZtZBX/aQa4CEop1TtQAeNajpwCj2dFTsINpA48P9o/ZiOaEVnxyuGjZibw5G/VL
B6RldbQp9JGa2t+KKmmE6Am5iP5EBgDyHURs5B296ZigzC3VmwZk3LIzAGwT677V
Kt2xt8UiA1DkUIEdyFand6pLQ9GmFQ/79IfIshqBRXI6Ykx2/xGx9NDSZVHm0Bln
goe1jV5KlKmN1o3Y3efXyv2U78QUAV29WyMNbDxB4kqf7BewILBOOd5PwU0eMXVi
0t8WqjWbe7LlNVeomXd53HeL5JfpiSWQaPyv9D+OYifNIrxHrFIWVYeORd+foSiB
i6HLKpwydNr2TUh/Mv/Qf7tXJMyES39JL9WD8ulMjbU+55FKCr32F22GoX2vIy1j
XCtUk3ndBZltRDx1dUZVBZxTHrdWtR36fRgQ+1d1EtO6A3a8P4SRZFeVtwl79s+o
SCSDIscuVewRng8MAxqRR1p5CYNcl/lNg/iig+locP5xsIO1GhIBjgJxXvraHAt9
QuVW9feo/ANrA+g2/pycbi9gA0cPz5vpKjRxGt5u1/DKQqi0pybvWid8lQEwDBNX
S2L2RfT9VGq7uN2qdn9W8yt3BzrvDmfv6llKqyGVSHhT1ICO77wwleclzSmIRR4z
ld7c4g/Tx7YgMZbtJQqEG/DN6teOyhL5nJptAM19Eh0CwfP9Rdjc+EysULCIgcJj
HxygFr+rtipJbBmakxUyDPhfNVskiv99nV4MGRnvgkoz2YzZqEcfosoDQB+Dtk/S
u0VJWSn0NJZK/1OMjfA9RU8NjF/BIwjOIRAxaDhaMkEISYNrbKFpcGtWXq5Fwm2O
aqTDEqOBfHX+giSvtxHNRShO3iHgRdaSfEtFFxKfO86YRVoF6PpOM7q36zI8yDK7
W1NLlHH7jODXswSy7f0H2qXcppvmzSHBMd5VUIMfuUr9eGkenACIMf7sKOJaXdQA
IDVz7GC57eGfMgivhAUsH0RrGokNtMMiHPau65t5CDYr5BLbaFOOCMGSWtdKoS8j
1OTscZSUwmFvuQ185Eme6kd2crGOQ9KlasDU5rI5F8RvkiEkl+tUlMLi8vVr72lq
8AjqSSDhlLfhNIF/0aZPFq7WoYrZ/Ikxa+mkv2BWEwrkpoEfGVdo9opyfiT0fCoN
z7RaCWwanW9hMoydqvspIehlCG7G03nJcMkjzNGhITirfAP0BwAxagCNv04kRZ77
wb5yFGJ90u2jT9qL9yI8Cbe+Isa8v/wUwe88mXvEQONjI7552SrmdaTplliywbRy
1EssZp0wpTTcgE9N4hphRbM3uU7bF8p8MGj5HnJl0wHjrocPq5d1SI9Au75wd9aj
xU1ZJINoCya+EWIn1n/KKGn19crW963tukdLrSReVL4RxgG2mcsK5QRCMqJMD3zb
/qatiQ+ViSwVq30js8jDvkB6ZcKYWRIt6Cw4U156OvvoMUzcZ2V/6edZcsj1Ahao
sQBZ0tsn2vj5EjOhvqA7XD4Mblww5sPBCh14VVUXEdyk6kd2EoOCaBuKv4KAGWGu
hQzltVrINKU3iHRJcR/PmN7MeThsKJal34188fyvNawKJbITIjDBura/tufIB+w1
pQr30vEBTfKTolxXnU3N5mVt3xahhsMJ84ZVwl4Q59pG+XdGpWCTv2eqO87wlSKK
gamo22whYWFvWjAwVoIlUzT3JypwKYjRj29ZUuzsUdp8mzJ1C6r1TluBKSOEt5dm
RCT3pztjZJwqsJyPRgsx5nnW4V3e8rTisNiDskjrYnY8eQItp8DiIcubq1QXllG0
TwDmTIL/A6slvUo69+mc8wcWoizvANNBNgYffWtJl9YXRMWGJlNJuFvYaygcH/q7
QcazVWDYLTUkN4LKEMBf3NhUkMN+uT9gh7DE2wEFixd2A0FZBxrPuD+ynrUHAFyQ
Yyu42XTzwqVCAQ0PGGsv63TPSL0x3b29bUTQOgTASZb1ScB4VVYtvUDDl30hBoXC
WweRf1sYZg6LSTbzmnUT4xsmVOyK2r4sMDnXFBgpvWsHHPIDxrFoc8Sl8k7SxqUQ
Nu6jIlAqwRCMIa+7L4c2rZ1ppc6H9gfitnTviiY6LMiQIfp5QvqgsVTNd38tZcEF
+/kYxrsx9kg1in/oouf7hbvDVPPolHlrD935z+QRir4EkUcUqhJ49PaA+EVHILEp
CPO6UiztbWOi+JpzU+fZf83EJqB0+RddZ1f6yD518mtd+wD1TU/TOPBN76pzcY10
s+lG7HSrGn2yc4jIAFEY7pOt7AFRG8hRhc718KE8aD7u5yicrJXX6yYhCR1NTKnQ
bUtOmZSMdkJm0MMHg3BtzFNgJ/f4y2gIWUeGNmliu2Yl0a91/cBDESYzFZ9Rkf4i
XD7Kv20Yc7p8jbBvP0rHniDRlZIflyO589kNW0x9mOq/nFNTMz5VeAOvFh4bV4n7
zvyB+UDc2fhnbuOj+7jdwpjeBv4cwUooUnawF/n7YdfE8CtObPFvBw9PFXaBrYTE
lhFxyfC2Fw0rmP7OMiFCYWZYwqS/oq+cmEcMX0XxW7t0OX9hoq2DiGp+ZYJFIWOn
fqHIMa7dOFIhqiTBX6ocFjYP1SYhaME0cqLrilYkEvX4KMPagDmn5fq5GRfTCJI4
WJGvvoP7Nvx6hX4uK/os6wMXhyNA49905G1oEl08sipUDTItUYAcIY0DnYYVJEwM
qGvxt9V2h/he/X7YNsQkTHKaSU3NVM/QCoQhGDKgYAKD7KW2MhcBMyB8ao7lo3AZ
L1rP0uFMECJ4ruf7S2ZJ8XzrIEyQbBcbgHR2UvNFMVsr1rjEmcrTCbiHcOOh9Xl/
Oda8H3u6obyzzC4wgXQF8+cRoR50GU274Xr6xOQXlrQN9h7dzYOJaIIn2ZoQrEJ1
euYmm+UV3yt44vy/vpvNhIdu0sBLZX/qBrqliPYU7YLOvVSBgXwolK+/a2+7I/6r
s7WQ/HSxJ2lgh7bbmXurLEucjOd2KHFqGNn5JDRcg4912z+58ZQ0oacU9KORngMp
eQ+0/KXFcLuZ1L2TGIhii1Sj8r0vuO07a2+fBcUoXvVzrvEIHx/hOfqa6nl/sgUH
+R+Uojqun0yt3IaqxESYL/qqdnEs4R6vP053pneWlIXqcm8cLxVF1EtkcmeCRxkR
SnWe/xSWY4dUkMAuTEhEc5JnWJavjf5ZRAiv0Mw9rYpzCNutiph1fcNGi5yq1icE
XV2CDbdNQfhFZaABJ7bl1H2QkxTDgIZF8hd7vomk8G6CQVwatsidoYlSxoQAlclr
xJoJSYpByHbRTl0iSRCM6ajm8BzPtkNrgXe4IkVvKLDMYIQtdJmamkrlCZUPYT4t
ZMts4MEhuRkAIaZu3QG3sYRXNRWndOKmPme8HdAyKqHxhyCMDrsWjU0mJZX1V84t
y6RtrDmKLPxReAI2e7icPVylHHoVdPiEfY3ozLH0u9PvDTd4O95Nilq4+BMTZ5z5
zv+9bF1L2QTzXMgXfjQ5OKZY81haaw/0rvuCvUaK1tAOvlk2/257EyPRzT+okj6a
Vro7/foRLyE9byX+snMZ39TFGmVyha2DWdxODLQyeGtEvjaRaHsqcXcMyefQV4S2
oek+pGmL5um/0AXfb8unQuovvASQ407X1skQcljbotQHCelMZzXvzEDAt6YEOThD
HazxX6U9tbQ9m01p+Fb4X8E21iylKaR2pay0k54Kew4a5bpJHqQgKnHDEPA+weQA
78vPOou+mwdAztls9GrE43YF9zQV2nZy8FBcaEpGodFctB5U/OT7T5xpXSd9UMNb
WTVNVsAvMyI51VyleEy4ZFmLO1KyVQ1v9ySQ6vHdMY8xB4MHNzOrvw788iFqDcU8
bXQgeMOFrOXD3YzfvGyIw6PGZAp5qISBxhwJoZAV96rNHLFRmE2EVs+urM4Ei8cd
1zKQVpdDgciH1R+g4ol4YWl/S402/cHzu8ZSmIP7VNQUXY1ZWpPnnWMjXM/soY+s
CQcDhJJZolCHKRsKBChVFOsChWYNrtKzphqi2OnPFaa0HPD/kzz028SniS7ozRDC
OxqDVW/Cp/xSeADAUk8w1bMfSkEETlxDFTGADUs0/8K0f+59nNWCQt9vL+9LmLDv
o077W9PBIo98GBGfyc+1LBUCJuo/pnX5pM2QjS/JQ4DGOeHLPLsxhklc0Oeik44W
UjwoSYkJzo+Hjlox4C/Xeki3e46+yfVUU7PEc9z50F5GBBOGqKWgzjM5VBmRRQN8
pZ3ZtzqXcm8XKmnEwUSxCbdoR9jBotqy+UgDBLq04FtoIyCwx+vsgc7TQu9vx/um
Gcnf7KPH3UkPKkNMvr4/K9Y0UqS1Ht42oFz2KQ2ZdfCyQhKcFh0+Sf98TBxk2Y/u
W0u06BrkaeiSr2dHRAmyr6Wcbso7sklH+3cJOfxL1fYfPmaadDO1BT4WMUs9+X2E
4+EvD/hMIiOCRpDCo2U4+33NpWS3bdFJqeeA9QHe9DVz77Rsp7dOE1p97eNDcWp/
MHGIYE4IS1JTJmVKIzpLXOO3jZQmZ0lw7W6pmcffGEaDpX0gbmpowLSaHn3HxgJd
NuVJIWnAd5yK+E8fbacOTUKQFFRdCFhC/1UiQHjLDiLaLTRFjSXzSYrmaecNUqck
zKKaT1nnD34eWRIDtNjjm/BVxVmlhmHtOT/D8xGsKfG2IkukAVUpZmfw92pOeSPy
ywYSYA/TlxfPkd4IBPNT8qT6HbAAJE+RK5Dm3RGUUIyDiT+BqpI9W5m7bUsrYkZU
kDp1BGbHXqcP/RQI3gujzB5qdCC9YZpDexeHyuGRT7wj8vmYfwSBKtGFau3D4d57
zVBvbATL1RpsOzoReiIQkrSQyed479LUckeWdBal4eoEaPQxEYwWrTxkFJu8dZZA
4QTEQ1yKXyXh8+0703nXEUoxePqiLMucvoh8iBSTqZ5lydcFMxnMxy2XUmcqTH07
yx3LCNz3yXdl2d68KEoxNzWpRUVRIq/QMBGKF79ybSnYaJlekhBR91VE8W09rZVn
Lc88ULCf+mad2KJ3Z0zs9NLMDivuoxfpO/YgFxr3jrVUBAWArA8X6+OxgjcXDZDd
jKV1OqqEnmXg8uo5wxfCCd7ANua+aG7uEEfsK/0eYoJf/YPcjlVPDFtl2ISBTJBd
vNLsVsew7otHEa8N89GFlqkzycMfT4eNRQUTyVKDxIYtRgNDa/kUP2QKYTtN6yKu
DUkJCE2Mc/qDiHxgEZi/lDaFUhSeg94TUA+dLAuJ93nTY9BkAQ4C9RTcm63uKW/F
bVm71CYHMzscAqp3G/0O0U9JFGSsdtDH4UCDsTY1tZ1gM5JjQH1MYpbwzNgQrSxa
C9eIdH0Z9/4QamsboIQJN3+6pIAaIylwV9SWnuTl2BskS6C6vP/QB0P3TBqbe4ZH
yNNtz8I+Iav3Mz+y8soDTu/FJb/vFHm1xZ3GChQ+6MpbazZBBOh70gOxhejr8Ikr
8lWLacv/fTh2gf3nM4RBhZUy9mYnrHJE57Fp/bFeeVmnlOPzMiwT5f9AwYkJp/dL
KWR/GJ90Evi3FAhrXzGFYGFxyFgnoffHjdNt+MrxkuvZndzk7X/vBZIL4jnc+vj9
nRl5D2qQ13afkqvls+C0eTum9qqUxmHcqCGajjt9GoABDgZ0FaU+6xDGm1ursK9C
j6Wa8Ks4DEv9Ietd4vOD7ERAgZ9uM+rJa2F2paLcYH7hEfa74dV69uSxqnN184gk
fIgjSR9jxsM5iMybajg4RlMfOco+Au3pZ5WfUSe7iUfpgmwDn7KfTLOSJP/ZFRyA
5NV5XVX/cNyr0LYQF5dXtXn6RcQwAVDuL+xfB22buwsb4nqOmYcrWUOhbf3Enojq
jxCzq61++NOHNRSARrqHFmwaauD8UO7OD21bhfoLthYzCAbMLj4ykSPz7xVZACf4
Pamzk1sfaF+JiRu7/cTnndZ4CQPBYVCUJP24DBi0B+aFzf7evnR+IxLfNAOxouhF
0yx4I9nQ8zLrysNrTBDY5cjh5lb0aDMcUIv1aac3RW29g4PZ0Ukc4CDG/62aCEwZ
tMuBkwLVsybbW4yo6sjGwr5wzZp9XOPER6eCCcLa9iJvostw7flRwDm2cDG5aNkw
XHsf2ofnoSr20NfphSnQk51CGvOSvvD6YjVPoTzS6MD76HbX9tSEBQm451pDH14c
MJHpKx3lHJXaBuksTX6y5XPA8OFNi3/ZYOda42y93E9kLnkHGN6dQ/xZzU13UsPi
oSZrF3jiMDAYHu1DmUZtgKZBqS97KuX3/H0vVEwC7bOOGRyjKKfCAuHCY6+pLF7R
RkdLCcHnpeoydvDlknJdUT7Gbtt6kAoBqnUKDxYlbLla81X/OR7+cPAzDQqemYwl
GUZdofXtSncmF3GMpWcU0df2XmCDljbLrb9r0IR6zS+jlJDKIPsihkd7WU7BIdPA
up12N605T5Caw/8ZLEOrAdxoIIgYm3DUWJKQjTv24gUPW9aoB1n54vr16tu3T98o
N93J1pKbD+07vmdC+V4wUaCAtj8hPg5UzpGVk/qhGiO3LF+u4OjCX9hrNmaGwSaf
PsZ1KxxxUrXDrCdYE3rvhj3XhkT29ohQ43CVDRyeZmNZSoeOQFwIB6dYQ9pJ0zHC
5JTV21wYIlPl5mGIwIbIzpH4khP2wd87yCTtS+ihrAP3vYWTFIlSe39H685nA54M
X1CohSHmxBua6qQUZFNnkpYAikBJt5KeaVpZyHdz8vV7dvK+ZhOhew1pOHWDDOq/
EJdGnANK9vm75urRgrYflqqihCG9U5eWi/6I0jyFOaOJPc3hDSGo954a5OZO3WuC
xPt/azHTcxu4GyrqLNjCo7jVeJcA4sMhK/s6pcpr4a/NCiYYdVjzzwx6v3JIjJaK
EVMYYSjYctOBIpBouZLZ1rtYYrkzkW5BHMc3mwebgcubskINmUUCkV6Korw+WvnK
1Xm3myrDPkhoQLD7u3Wh+Sl6GXwJIqIGr6oRSI32VisXTyd2kXr1pqkUJVtvUMtc
X0Ki+i2EscgZI51F+QSfy63H1xAfUxsdcMn2gIIWGX+13HzNPlCqNYS5Mdb2CjRf
ob15cSMd/uwnPzgmb/ZpQgNgT9LHnnBat47s4wAEO8uKB99VVgHf8r7uxkRxECgL
IcWTMH2p4j6rr5Iysv3ZhVEAgtCpF8zDUcOfb9Mn5eiVip/BKqUdQos7xBpnndx5
TYx3+r/amh7hcMHZCc1V/B5K7pQ9mH0cBT9mxHRHvp35n5uX8wQrMhooW+KWvaLP
lUcyETwOZ1KPssvXENKAWSQcwQP2ZVj5k3Agx6T/PEKx+crm/7Jgw1T8+LND6dJp
7MCe9eVMBn7xxXwJL3HBA5xALbsJmcclvY1p7dvfq/QsbCFMTBm6WI1BzJZTWbXM
4qdDrfXIksFeNhMnqhqGXE18YFMYlfMmKX7fv5xQjVJ/9RR/YYOrmjl8+GjLSL5F
Px3BKXfp5Tdd/aB+wkAYWNPVMAw6tAX2SoTjt44FicmTlYimqO5WCUBCrZio3zEP
5SwBiLdNcmyDmRo8Mwu9ons/QyFx45FF7B/mCwzs5uYbnncN7Qn74iTF90TJOAWc
mIXqlAhB040OWMdWJowVU/Jv0kBIVaWcyIKh9R9dHdif2HH9uxxgkibeoEPjrbQM
GOwudcJ4PX6DcOxi4DfEV5qBhg4DIx4/omUAGOFaBk4dkshHamB7BJGP4n82oBUE
fMPColT5Xj12Pa64y9YM+JyjEfQASLtJtA/XKUetlsdtcTd1m3rcRSAOwGhdHwwp
arG848z7hgwgDGw1UReJgfhQhj8bAnwjomVS4ZN4iTOnJF3x5HdS8W/7EVQB2Dy+
Ix6Wu44TnKizeMVY/lZ46vnh+QTH4GHny3z1KxtmEgBwlqv0lekTxzPgryMpI+Ji
jBX7YhzAVZJaXZY4xyJsaLXoMli7Ik9CdDgXuGrjDiNtjjaTEGqGUGBzqec3kOQI
hXERwyd9XbAcUXi4bHISOAZ6UM+82UfjpKZEjNmCJ2i9vZQ2Jm8cAx/eX//kFp0J
bIyxpKFFpM7YVK1PBMKNuaKl9Sz2iIL7q7H46YYYPjb0T7GVSsDs/6e5gBMl2x7o
zjtEGKHVIuHb/RvfG2xElSFO82fVoSIieTIA8lgPfT8hSAqTKv6n5mU60KMvfbTd
lDtY9uF9ilz6JsChb/N8DQmHcHJ5Nc6iVffgdm04KhY/xAgG9XDLrFPeW1xQo9Hl
dHGXBbY6/AUlDMrdSSOsww2ZA/kklhE13ZrNQM72zQcu0YZiXOyk60Tz3b269RXD
RzQnbZ7gXu3eEvRuVvwMLxiPkg6uDlPceVT3J0tZmvz7oeZTYJ6lhGV6ZwGaBBcP
TVXllnYfT3ZWNF2H6I4edJQbpszHQcRDhNb3S+e+JqjBQPl4ipGM19dGrtDJ81ow
0U9LpCoKpRWuQFYrgDzAqtunYuIDVjeAso/yZ298e39WzPI944wWMkgY35CAmX5b
IOaBFxoFqaJ1tqLnzDNtMgc3HKO+GZ19QyChrJHKAntL6iVZjaFZmvOJFUw9IacQ
QmfaPnNmkeE5ssCRJRQYgxF5PBRIiJ+NPls35fe44fSzLaza8I8oM/SX4GUA4SEk
OhdYKercMYPxMHPISq92CCX0mWaDfgg8zBmeG5IA+5dlrfUZz/gKTGVan/sYryax
XZehYbcQ+Q4Eb7prZCULe+5TMRaJcKk9519FOu7Wo8m41NuiBNuSFaBDT/ZCvUJ9
1QjZoHlD6W62mZ+BkbD4ODPwXh8Ij3dMj9bb/b8/3gfJ2/merSTDFN6EZ3X8jRF9
ic6vUwg5lj9aGdEQYJot4Jvd86EGTa+6ba5VXSjoLbUykekR2F9sLV0Nl18IOfZT
Npjjpf6ex3au5ZFjJjIdHPAFzHhoQ9Ned2AX3+yHaG0mloADF2VnFQbLhJu8EZCg
pgvFychv3YAQibGoJpKZDGawftxacltWgAyEe5fPBL/BgLtXnbh3Xnfa6coPQdxS
5r9ycl359DeHune0pak1jfoV5S/KZeAm3iNX61nZXEQGVd0LeHZbd5LTaEGjqluO
fU1SHtycX+WnrmE2Kdb9tj5R9aQhcOu8EUih1GMxqL4LPlFhfif9N4W7m2LZGLdI
i4UjFWPc3mJ9Yrf1BKCie1scJxcYLhg3iVNR3r16QEaK/p5nSb1DX2CDDKDWtVhu
KS0R5zqSOD2MNz/Mmvgln7lOWvVQi4zRobDvxQuc0sN6rsns7/pJNPUtL/PT5KRl
xoZXUWt4g/ssPxSGIchoRoO2z43HIam5zteSXtYTbB0/KyuQEhSPe1yvFdkp5JeC
z1kYzKBLQbiWr935ahmkrbvN3H8yqAX1iGjZFwbtBwGS6lGdJhMO13d8as4cdbUN
CzGegpZTar1vp5NFMwcPFElZ6fa2HOR21vwdPMH+jvk7zcoZVAX2p3NnQvS87dtA
zn2WVl68BVsJXOp4F7xtEYS2GPr7LBPHtJ5PATBESrAurAqmLRiS5kmbmoAfG5pf
Tba9WKHCFNrjITI06aSO7iEgUEqu15/Dd1nwAhKjpVncbKOb0PBprpLyk383Ji5j
OY6sV7VaBhWHr2Jquotlkb4Qlar7Zscz65P37fkAC3C+jqSJ9LLSP9Ks4N3miUAd
wbxj/Lp/NUR7enq8Q9GH6DQL1V3G4gP5+othss37nNt/WyuFsVg1E0dqvBzH89PB
hhD+nx3uaUtkT2nA7LKENlCXX1nMI14PgNIMj4dR1FlRa5B0VP9LNhwFX3Du9rbh
lledD938fTei6QPQux3XVOJ3xYuDQSqPevmrP5C4LZYo9gifJTuRTC2EsLWrfDBE
k4QuQQbIAX/Z9+LgkHC6MQlSvT95Mhfsc4SpIvVtnqKISqK8dgbbZ+ZjixxoJ0kH
ttxvsjNqlHQgvmK6lO+1vtZoWIYAVknl8FXlWf9pmffQ2mOzdVzqZt/ay3bnQVzw
HijKlxkVpTv+HVwD5I9xNSF+pO6ZOkHC/teLUICZ7P0Z9hHyjChF4kfgyw/WHi3+
3lQU1dwm0GsYze28+C8s2d2Kdya0MwOOizOtWhamo3+YFnUzY4Qq9GjPvbujQKoV
SEcThjugLeK2f31wbyIrwTkU71I4h0ln7OzbwXIuHo8QGlDX4dGFFLH1eYh7eutM
+89Vxw8QEA4GcUzS/hK8s2Wt0brNXRMUi0+xjj1Lm01c0i365kvUsLqamOQr+l5v
JcYR/TTEqqRZkPVNkXUro8dAgEBqN14yVkMaoabdB9gVbJQx0vE4L9nnu/CsNUFe
xB0C+a3ulyu0qc88kwKCUjn8YTkxDnZ1Liw8LjNai0tmRnf4KZ1ykEM2ud4UeyeR
74Mgs8i9IgacpB7o/VfANw1h4ori6EyZD9M30r9cumMj2qxCbEb1tFKypmzMjuN4
x29OBrVMA16akqXZjGClH8kPM2Zm6wNyFaO6s2kwA0BPY+lJ00fgR+U6v9d2bFVe
GI5QLEAYCRe0m9gWS76V4jQAeUyVhWOIp6Kn0Rrr+CnnCVRspdWZECrTMNiCT36O
S4LToxdBJiyAgUPpZrdo9uqnmvn3sUkdB1dLOSeJovZ0YLFlTEm3EuGDZ6bUDVIX
D/6l92MAABehza35V/FL6O3gkjsoXa23yXKSKC2I3J2GVPUuohIRG6ePMGelu4n4
X1Dli9sPmDwDqV3YsvekWkH782ux5qQiyccexx3MB9CzoVZ9QZBVNy27Yr/h6dtN
K7c5TImIolbpAKB/IwmfPQkMkr9UxUCa25eRuFMp3rzTqPZTR5/axA9J957iwYPf
GijWykqOZj9lj4s+me0ZId5mT1K/QkRDOkppcdIJ/vz0h6fc6+WgSzS4wR5lBBL0
T/HwoilwKY+SXpac1ktF36Gb3mgtmO4EF5nHwo2SBfUA4YSecv/JhmelLejpzDat
YbPspl8s7iZMV0L9TBeFiGLzmE6xs3MjsvWEBiDT/hVxNXhTi98zTlvjfpet+c1x
30DOWrv/GxI7PLjB8CM0IBnwPjKF/VpAiuBMUMY2+H16tBkAA0EIukARmAzhWZEE
7nX2JJ1XcKAqi+nKdKtxXBTioGIs2kYFw73r1SrD10SKHHF+3A8+PPkO3zDrvVm6
Vnbzi6ct5HLtFJN7YIz8fRr835ZxhgcbqU5g5nhkvXz0t5pj0zzjwsoPpg0xJ778
OdUTXvFfXlqMegLKVHQjEZBdYD6T5OJnYGEl4fZSuwUNZdtkhmB3HA68pESga2OI
PofDhZdhmzDS0lklYnEjRbUBSn9MPRfWtPSzn88FvOGUH2Dohc6NKzTqowott0GO
xu5JT9G0gjd4FczJMKBP67mg7Z0xm/jM1XGGfpGaLXq1p+W/f2PNZdBmuIdOK+Xu
E1s20jPBuNosX1AGAoTD/eU4VSs+2wO7cF2i/4l0Dw7Je6HKhwYaeQcQykTkcfe1
tzutAeP42ryIoKgs4+Htm4jfPk3aVwGMNXei85mX6p7QiHW+jNkxTqRj2Xj9bo/K
j4tQgVGYRTlkC/OTFUrkR+i7rJjhdTEWfjFU5UfAz6/UiFX9A/p4kqfLanA49lR0
S/M7Qx0e3izqbcovZ2sVzTsq6Md/6hKJ9tTLo5ChtDZrNpT1PjuwTA0NgSSevnbo
x0rfTQb5Dzva0dwQPvwORD/IIUNUCIFsKDSGcgE7mAWqUUxWZTLvIMikE+ZqjU8f
0APROSjz/8aqDGOqibrwnGLJqyIYWOHzKTcieGoQ55giNs4E+/jR/M/uEeuY/nOB
YGBVC8loVep89YxoIwgJzbbiejRYoGPBL9mREhnBGmZYBf1mgQUqrAKetouU+Ano
B2P8HofrsL31KRYRNe/6fXKaEhQlawshGsdCHrozz1ltOwXB2vDo0FwlBGaNfw0x
MY+5o+PPEDT6p0M8PoMbGedJaCdndhXgGSxtvvJ1npG1oGCzhONZNseSGlMMq1Uv
cUHIcG6YafAsJzC1VHaIW4fnCCJeCjudee7ERL4EZp83BzYFr10nWOZSzCACMdft
83a8/uv10VQh0wkFnuo3F4anWnlOHEkxdU0v6iQ4dOseoeWH+ad0v6va5Pfk46hK
tFjUuWDt69LFTZgGJ3EysUzmuzZkotcHeWHR7fb0nOtaruKhoqCj225D42gzeAr2
Ta8zPjaiXWis1yFE+d9qdN51Ltjj6iYDYj3s/dnX63S6jtCMg6ZLjBpJCRD+Bo7O
q7xCy6AOo/MVnoK/mXIgOFS4S7UVC601hTLuq0Dtx8zhg9bxlDNMuqXZ+Eoj0NIy
2ygFj9dle2cKXKwADvJCj6CmT3SiXpHhBm6OsQI/C/unYvP1cgVyWv8q2FMoryLL
B6zzQe14X+0Sp02bf1aSwGSSwYj428DshdMGmIJ0v/LqMm4KCn8YLPYmNIlzYnOu
z0iVcc6S9DJItv3HEl9ng3IyJnk6vmR7iLrEiO4rrpJWNn15qWUiMuhMZrxeI264
V/LdU6DXciEE8wY6bA0qjKgVbmu0MvgURoPGefPDbVYfiiVD5+szZGt3B05VOPi8
KcrcDAL5cVfmjyVegG4g2sG5A4I+F7/vVNEjxzD5wBACEhL2vhxyQC3Mw1R05x7f
ClCoqSaIUm2wHny704g+BC7cCYdlmDSj6D7d3FYZIITC+wjBvlNP7SIDCjHhsW+t
L70w28hQuO7/zlgP0jlnW9fAv8qCKBLLCygZMAf0gwsy02Vr8LXdwE8Pbwc+5ikK
W2uKBwJv2wVbARP7N8aX9+JL3TYqQ+PLKeLtm0GsMCaAOwoDdYARCjKM+hkQJlrt
zt2QPEhs9SsQxfjDzXesVZ3QeHARsBTWs+nHa7J0mDV5v9MOf3gCFmGc/A0to4XN
zR+YHA6701/p5a9MbqJyhFbQ/Y0i+FLi51jXvpXzhOzn9iAnmx3g0pkyDx9GLbxd
BvnG7PNVJYJ/nRfcBmAK4LJCa55tVQegxSgEScDok41if1nlvRFBE8kJ0/bwFYIs
EgG4T441eBUbJfEWGbToEf061fwWrKpKEhZ0rerMB0qTl8vk6+bwPFHJxVGXIQY5
0k/6aPNhUB1D6nvL8jGGiA+1Vdz120CNVNq3frVOLkTTbJxQ1u/4s51c1cqyP82m
8k2p6xysM6J8kMIlhUuT6/adGgayyzclVqE573lm99mTk0YGFnVgO+Tm08YWsrUb
WnupJv8cF63iGjsrhrTPmy+LwvY3jnNIsS5HwULFRihtWnFO5wwGUQEABB3Ecqge
Zi76EFNmj6Uh/PbPF3jcOcjLhQPEGAV4iF+eO6v9mQDv4Fxm/FdHvS9Umz+vJZ/g
CvXgzax+wqGII3jHmKSjVptbPqsiP2amKvyS6kCXLhvHcp0uQwFk1zidlS6w/u8e
k7hqZm6NK2Fui6VK9G2nTrDRHRZmOYjSgw6hX6dcEzSJMqvF/EswUsiPFbiKPwsr
nU7aqLeOxxAekAGGt/Mu4BNDL/wKmxTGzjIo/2Thmvhf5QZ0YBBpX30MfxdaSgK8
i6sjmLr6CTyTVgnuH11r3Hl0T+bNc7umoSSofhRKKakwXHrBH3VkWfusXO1ZUcrg
Kb08Lg6xagxE/jNuZa3G7Ks1jtDLCa33/puzxoMwID8xpLYCt9cCnsbboMB4J5Z6
I/6MJ1gcjpaMCeGnt6wk1KvvX7hXpfUvE9uLApmAAeBc5GB73+CwqdRdmrL9hAv3
GDTCy7KRK2CVDeF5NLhkFV7alMhCgXGBxZo9fG2uvfpVZ2pXIe8CPb9N0ElQIUrf
VEp/oq+GkKd1ZCWK1cbmRaaT2ppz2Awy9Sa+UYZrHxipJD3OgkdMHSN+ypguSVGg
lWqarwnMHT2J88TviaPrcSyROzpDDGWNUEMvkQJAwRW2NhvsBj0xXPCl1JXdx1Rg
AY4/7nkFN8eROb7xevFPdrQ2SFtoAvXDSXBkXVNSSOygxCObrLORUr2Jj2v3HTPX
5B3bqS7RQkWRvdfFKVY2kBKCU54i89vJ/4BAtaT4AGBYhnuuAQvLjHjrzfMCSoO7
f9JYx60KazXRnMwgZla3tByXr1u7mkpQRbEJ6wMtMuYWWC6et2phB+MCkW/UBSc2
wkJbcZ3eNkTYwdTgt5N3NRk2MNndHsOKuDVushAavMP0UPsPXWwKmiiF154IdVyt
8FjHOqgwf8AOQvSF9qljIT7olh+N4jmtazolldRId/4GSq8Uo2YYK1SFXA7ZSwXN
jfo5h5761zaK66QLH63MYjU0gPngj9AUkjLauWJ9BW9+FSfzPeC72xRLjIOMLZbZ
bhvNbcnqroqP63hA0uoQcZMSzryg+oqjtTUCHsjGkWZqu6Ul/sqkLnI/t4adOLIC
djNKSDCf/clTFtvo+yAB7LLz4tI/ii2pacG81AwiChQmjCRCv2Dwqlv3tFRHLt3J
vs2flZK3KIKVPdCnhxXullBozPrrLGnf056Zv5i4FzBbkE+MV8ZPobdDhJJs93my
mWVZL4D/7r23hTP399p5dzW033jXMQTHCmkd4wOnYdhF1DmMHu313P1g8IR8yHuW
XqlOR8XTyZarIE0NYl0YjvWWmdG64Igj4au82aHhzKURK/DkGBP0qSR0MpXPH26W
bXKHW1G52d4zL2/tI7601E7xM83P1mqUWjQnVHc/26KkaaarxDfBq/ujDviaYyUX
r0VAZ2M903l2IX/337VHJklWEnNdRRCBSwGqSx7jGu4=
`protect END_PROTECTED
