`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG+BpycMjsMlaSswuBxDyG2wMAGRjbRswZONjIVdSEW7
2bwT8ZfZk0FxoyopWOIZ1UsFffyzsnJkNsu8UoehQk0Qe+KzXe0tn6huExZusaR2
7qFeSUSkSwbIFbIgpZ7DLyWznOyOhyBCm2PGe3TwGw9+kuoU8U3drDpewrYLiLoV
a0Wu4ZjbcEyMovZPWe6+T/gjc4l7oqMSPaKQQDfotRjjLMvJlfYPtpvokwhApiou
ZObgCAaOK2IuG6vVUIhZuEjVok/kMz+xGJTxEALBy4onERA9pzhzSjIUZ9IxbwzF
kJ4Ype/bI52vBskVEqkGh88hsWf7nF3SbBRI+DyjlMPQWsa/9qJO1qn28sGb67qL
mq2EJJva/y86WCPFAPUCTw==
`protect END_PROTECTED
