`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pLYeKKoP5v2ViFUwYgl5O8IqHvbLL8hNRwtp0nE9Uj7rDtd67ZzuCUP2zSS2VYfv
q8G+HMp0tPycbTVhaCJRAfa61YCWScU6+AvgzPU0rHBOsteTtqZugYbu+eTgkFny
m8mQQ00IWaytdjn/pSuIGLkIXgScxx1v3ejPjHDLWhgv3IqhzLenWsselz02ZllQ
fUQckjLZnJmM1N86TaLv7EOd051UoJ21zRyWMLW0kVqXwN+AdyxQoAHXYGUkb6WR
xfVq3OImr7eIPBrHwHjzzULTZmC7BxNCDRLIwwug8HWt5LoAASxod0my0l7v227s
`protect END_PROTECTED
