`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aac/t9SOIgudUB80UtKfxL0MwzAdlkGO73Z5NmozYRrH
9PPlDYF8NjhDla1yABs71urHna1TPqPXrwSvcoXsmobL9wCGYR14Cxs0NV2pYVe1
Kr/H5qVtexPM2L+D/uQcFXO1NzeeLJhEyteB+3tPLGc4H0juPHJqY2jhYvsFTnxI
xEtSJnw2eUdJtH3a4jODG8i2us2rhGWVxE9XygWB2jktr8684RXqKKd7n7xDWRMy
ed3ImQ0mDInyqjKekWAp0yQh92MhPFx1Cea9IPrWJy8hYMOeY16UCdIBGLL1NNtA
411Qu1Mt8etK0pqqjGwPpk7iFudTvY3k2R3nlhcrC4/1wTtMIrKNZ0+22JISl9MC
CKSQAFHiWZ+LnJD/rIoVWukY8M9rXW2CyAmIvbu2UAv4DKiOZZw6m2q1V66/u832
u2LNqI2Hnu+gT1Z2+rkz8BHZt9Xm7Mk0OXLrlhsMlE5Yr71L+9XKSVbhOK8SsdoI
N77XClUDLYbi3Ss7qAx+/qkus0X3+/p6pKQoXyBbQbAucieqfL7rt2myVmsdTKwB
8TXeBGE2Cm5J/nXobOGvpTaymcG1rnWRCrCjvc4w8sQfmCcQHergOkMSrE8xUzJX
LN7gTDraFiQrzOrUk2cHRnFHN6tC9xbetq0eV5Pc0/QfFnxyLMcYimVqp9oEqYI0
+8PMJmBnh4w31MWhOFFHcjys7+mHZHnwdDWi00I8QP4O9X/qdHKftM1+94Bbzwnx
vaSFzmKtZHG3EZYafHDxBd85cO4VA5bif8O292DR6FHzGBwZC65w9hn56HnKCLhx
PuvRIl874NtdSQMK3KLdhZlTrYT0O6IViCHGodFsQA1bQPhb4tNgaaeyQf0EQ9qg
4Jx1OeJQK77KCHoFLARv6BwnoK5fOlwA/h4sAxhdbn0UXit1sv0cEhjbfVmbB0k1
xdrsvA4JxoShvnEnKlIPhQlXXpwOnHF7DBhBOv08IXZYDVbNGqewTPYuaGwTgXDg
0qCXqCtncpHOZ0bXH9JIqeamMy7l6JYZ5UUqDeZ+gEKGQcC+8bK5atSkS5PIzoLJ
oCfT9BC+KSFRmOg4uzhCqQPnW1Gtt++VSiEBz9YpUSpX+Wxn95X6xOetvVhgYaWR
vrbbFYKt6Lps4r6fb7vAQQM4tATneGKEYexWU6L1S5b0h22AjNJR8ieaBEGY8k0D
Pjiz7HzSLXamsDzBOS4u9m126GqfH8E7r3tWviakalbp16k3NBLsoYYdHuI/elXq
TBmbO/5vt0Jk3eDVHAdVNqW2guVXpiwGUxhcLgwg3z+IYa7Txu8kblZ94jvS0p2d
ZmNVZznbmCLgsU9uowVusuqsCkmEugxU0gts41+u9SwY2Dovc3WbSPm4d1Ts7n5x
kG447ydXP3WirKmnF3fHqCP1+Td27x0yjRSX9ytHcAK5PGfftQrAAxSCIWs7aq2b
LMTasEp1XRwqSZjTgauHyys4AeCHAkco8NWI6XyWlWf/upeA/+rJP8xUeYp/67br
5lC27Q0TuEBIEkFUvuoQVQ/o5/OhOGVcVyIODC21X0Lt4DceM7xgVYMo/CyGF8Jh
X/dI4dHduN+D7O3svzDr5d6zsivYcL9rZUKL6BIeriUE8at6n3Tj7Q/Rj2VqrbjS
8wBuKzseSmrHj9Zam5zttrsUpBYHmwKJLBFmVWcrYccA+nIV1bUIVTDR/7uFp7HM
4gkygcKs9VdXyriiLd5fEQDaAiqrqQsD1RVs5Uy1Kz1nml0TF/Fq+nBEQF20lD4C
GP2ufq0FwV53cmGl7iGW1vP8zbqFe0qJQaRtxIQlBIH7j+wQrSpK62evZ52eYSVU
kAdjoHQmgPC4nJq6iX/WfeKSjZehzvszhF6BiSSSlDP6D4Sgjw75MQwMLjsJLGvw
c8iLzkjq0rwQyOoALXOSOCClVxCLEOhP0ds063sSQhojUjB4CwwHtekuARLqarU1
gXfaj4hPBZ+e90wWweOu/rzbAyJW77XBV8IA5sa3a0+KCxgD1TcVSeWH3MGJJbZC
iLb5IJ3xJoBQjy4ORGWDPpTephnfca53xrZ211YSKL3YosbsB46ZGoyks3yvrZxj
g6/BBfgj3LaqMzhirBEZOSeF0978F9pUjmoRBmN+FQbcQtZKmhBbm66AB/HN6P2f
8f3bwE/GNycgsygQQB0YJ3cP3vPrHC5B7jNoVGjmcWuYqWMyEW/+VBW/F31S5iJF
w/mcCK25Pe+o7S/PvZlDBP8QZ7a+JxjFwHj/3bCuMrsp5JUhRQK7h3RYnasBwM2K
yvQ9cB06uawHmCjfs8xEkL1O1/48tplBTg0YvZzhz8GbZvtj638XVkxWxZ8v8hoy
SFNcT21JirIIEb8We3YwByCgyI1Ft0PsapxVinlnXoLe0bRy0Hu16V85Pg2uHdKt
pj2rX4xUpS7/UYgwPjVLXUVUe8o9ND2CraZAcbTQfpOMuJUSL/Irt2Ulyw14H/1Q
vol170FuNtaV5tf6qhc2+m2mYdTyetEBZ333GVq9DVuoUJV4cRq8ubGpqeLZde5M
9Afx6nhIDA5d0LMyOURMFRKKorXbM4cQ3STyLVdS0yPw+2Wnet/jBTZFJhVrFC5d
Poc3zvIeXAVEvTycJf0+s+7MOPc7AzswPCHbfdzUJgfgH5qBfUyVeo+G8IZjKtt1
2FehhEuMGBmfD3T/Dhc75X5XNOs5jvH784imcrI5820vMzigh3f1LxoeaPTpewPR
foGe12nlqnmWd9kB8E2UX0dFImhr8M091L+RmUhzXkhd1K9rQ4zI+qCv71ZLISI8
ZDlJQ71C22h0xEErFyfeHOeNZjT3qNoGkmwJh5KcJ90D2u7l2e8aUVB1SN+Cuu02
k1ViG330LKx8ncxLSO8nwGrmyp4pH2NBQHaBh5LOxJaIj8c1zWNEesgZ9JmfUJ6+
va/7eGWyVtbCzElxruodsizVTWAF5WkltmQ33HmXKvVFIpflCmwGMiUEYw3N0jrF
UqDMu6XKn9CRFMddyGYbIsWafR9HTXz+ZtgKoNLk6t2zWn1XXuWA/Qaw0bcCYxeN
XjeFAMi0/FF3bJ+Svm066fzN0gu4tAyapZlKcPbRKsPDA0ZEpUWYvlAQRPina8qf
5HidjoXN2/L8M1gKBdZZwUD3GTAQhRrx8cmCkTmh3Y4m9kFB5ZwA0ek2dy50FzcI
s2mAsjx/vT8p+Xr/OG+m8/+9AboZKIfYvCmXy0ZwBJ2D0brhMn2fsLhUMcMJm26w
YM+yrd7LfibakaPJXmr1xHDp4UtkX+tBXDcgLOOBji3IIKM+2D1stsubeHzbBcm2
mPRfZiWwws4lPfGzc/+/m6CY/ryR1gXXfJ+wyUn2UZU2zshMn3mZKKAXJ8wqC4b1
HVtMcOFO1u07J7SdN00flhvVvfM2qEY+4GZEOdD+atVb3lk8RFOHH95yCcO1oQId
oFAhUxcx0XtrvXrsr5JFAijlp7EgE57iJvhLH6Kg+k/VFTgUjxnJ8hqooM64gcpt
vteCld0X0hRXvMU3+Ocwv7HDTSM7V118c5bZXTouGjoBUDdRR2XXO0bGUkpOTAjx
SkWw3dWENOSg01HZ/OAbNuYUg4WhfJSKAmdal0GCnZj/M3Dxq8yZ8T+lpFxuVoAX
GaVL46cakILmJACizJF94Ig3y1a6G4WyP7/fj0Re1OPVQU2M8xQMShXskwTxgeXM
AKYAyZhYIlmB/vV/WExVeGk3r4kqy43MoI/c4OyqmWHwt/tvJDMAD43V7ty14R8i
Mq8VFYh0c+cf1jythNXiJX9RwjA17rjh74esFkRGhxSILWpB01bQmJMgP95iI5IT
4p3vdWfnOZg7bXz7KPtvYBccipcdQzptJjiFNNfShc5mEe0vEfy9jRZEBHuMs2s5
NCuSwPGK8GYmKDxBNuhm8Y+VRutzIlYWNS6ZkHma3rI2Ynqq3ZvPwTSWzliFtec6
j8325RrrV+sXCGYWHiHf+99lw5E/RpJ8z+vRhCZbM2Y9oD6cx8h/gYM3v+OPq0tr
JpujuKMLCSIOWBy7irm0ej17UIdEfbz8lJ4rIVyVhsHti7Stq2zlIIvzilMe72jB
V2VZfvYYXfM0hlESrfJACQokFDM2WkPcijO4Vo9/EoFvsZaNrwFiQdlHLrHJ9kJi
vtFjKxDcvSx/zgnDPAx3wmShOBejODwFc7XYEfvYe9OSEiO3mTKCQwZ8YFPqBl1K
tQXR03xWuGjEjEhB0Z/nfTGfRJY6kLr38Nb26NtIVGg5CK11wo6iMx7cuGm08jGR
2qmVzfmTMFTDmija/LrPF2Wh//8EJANJLKRpzMj5CGYuFu7iLTu9s1Kf9dCNrmlT
qm5ARLot3Pt5oZKPI5ynEphuQvnf+uUBTjQQKhJfY3UBwjXxKm0QsK1GsJWKAvIF
yC67m45KM6Ru0K8uOKONeJptWxipfdOviQVpc2E90y4=
`protect END_PROTECTED
