`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
hM0uWiMykzCsTVvW4ivy1CgLaoxn9AtdLQx6X5/0yy8FqOnOpuYs31j0ZmwFAOi3
m+eCZ5B95YvAP2DF9ym2omxNFWe8zlw4wWA28fF/cUEbLDyL9jGmbIdvwGzQqa8V
r3Oz0gbgV0zWMCGodIWO1JfBmKC2WZoCo+j0b7Loc71DkemE2DE3Elh94kO5X6lp
7hKRF15nHW6hXABQI+/53BpzY3+YKYj7EeMvxOocBGzvEQSQzw19t9mtA8cg0aSj
0FzamdWN2Ij6+tx1r+Akp5mIa/krkNHVKoz0q4NXhQPyZxKI/9H/1BlX3SrkTnPY
sJMqNboyhPlrBWvR/iN2zlY7gcVdAhik+TjN/eGbfvU=
`protect END_PROTECTED
