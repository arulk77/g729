`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMbX/Hf3EgW0y2K68cfobP5uTieV8E15M5eNdhoaMDSJ
GhnChBjJ2xTpXiFE87Mvq7ytDrW3I0c4qA+uG797nWCq6GUPfQ4l6lK6M62x3qh0
Cve5J/yKXcgXf9360cJLrMLocUY2iy1PaWrTLn2maOo0NiTByODaVK9fAgW6FcnN
/Rr36umLdvSXQaYGePhRh2NBURl/9eQQJmU7wm6B6sCP2s3uRstwe2hHpswx/MNv
WF1irPwG1QYyjzLImP2u+6KdXC5jUqeZI0VwBuuuCSxIYxQDleEu14bzvGT7px1B
`protect END_PROTECTED
