`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44lYa84Kc37S5EPH8e/pnGVodC/lzlDPeZxAFuHq8ibV
AmS3awDvo8fFS4OTIZGdU2Fd/Jf5vLdb1nQPXcITGrNRO0vgiSD14RsRNdn1QCc3
hyW0diFhJxIV5J3iMe6Xu8zX7pSKtrLHwX0PavvAXG1cSOR+48v1tvkrCS9v43Kv
9mylxeivcJz/9aXSOX/eeYQRcQiUM61Etg1We0DaATax3xex6JqhsLSjWQGiF+Uz
hDohIjiQdEQX+i+QxjZKy/asQctjOw6xo58g7EWzhNUD3TH43ge6wnBP/hcd3eHI
MdaUVovPPS+n9D1XnrI9Qw==
`protect END_PROTECTED
