`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveE+bGDDSe/sfjIp5QypQMbHYXCEffUNr9BzE8zkh5tD2
yK543+WL/JcV40t1JyoJ3WSD7aa+MByMluyqtnJSje5Y3Vwhe8t2915iqMGjN1Us
ao/za07KGtwQPtuW8RKaNlMsiZyD8vUBsYGl5LzSzg3hDirpaeuKxMHFuGWVgS5G
disgSHYDqflfdLJtdqJl0OEAy5KCpjUarzuNNUPe2F/a5Ei2px1HgjtrqZXAvE8U
x5YbTOotrohqdm93g69mP05U1f4+4Y69px3XdeY+1z87+8RKZMNHOpkz06QQLb9a
AMxw/PyL5eUcm2VbrWRkS0gGU0wM3QakhuWJLUrc7Vt0YHZkYh013nHiTPPV+hFR
JUrx79hF9+ftdjZUHaPQVA==
`protect END_PROTECTED
