`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu474zy22keXiAWa4CPJLqL+ZSiE6xSy0NYjVbrqjB4ryD
j4E30O7Pl17tKB0RQVTxMiz3/pu5turcDnKEfX2IaZmIcOdxihwiKdo8k753PIZ2
Z8y5MjQvO0hrs3Eu7ycRibGQThBVfaQgEGJyJE6OCrSZqefPRR8DYWRZ2CqucQgV
HzE70jlk4XI3HnfRFAWeteZCuvLN23Ca+Qh9sfAxw9W21JJsSvPeGNjWbBXPsumW
QNcWa6oeXfXNsjcjHSH0EwUoyqa4W6fm90uONYASolPiaV+Y87DFHVCfjRlhXkSo
Q4CclPKwauSVLb2ZbcDwtw==
`protect END_PROTECTED
