`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIfXd83EuByKrJOEgzQJUVrPcow1adcqxk1QqjerRSYk
8mf+HkEVmaGip7WLF4zo/QwB0SyFhI0XqDYeRizE0ofVvABKsx+vKR8Y9TRNcLfv
DyTxfMJbZd7oKT3571yvsNAQVyB4mnuj6DQyC5NgZViTdqodqTdWnRiydvzVji1u
PHPMAOvfMz8cceZam+gHJiLr4DWsrEeqezsqIeu6khyugljClguO5soLSlw9KihH
Ocb8Q9oew520FCKlcqwK1w==
`protect END_PROTECTED
