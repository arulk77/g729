`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGIH8MW49t/9qebG3jNBOZPgGxjtVsSMrsN8Wf1FpVij
1x2r9Fm49oK4NF909etpb8eDquUvipaRGXosqOIGekArhT92W/8s6B0PyG26ganL
DlRpXxfhQiiwvdwTTHrW2xu0dZRGm9oqE5RxUEz+4x97bcj7fUOWS/JbnJsUcb/z
Af76lTv8snb8UaY/6+TMNDd2xIhC1l++OH7A/hDGHZ+p4vAsl079/TpIWCOAjUmO
wX/8uytbR0ituE9JBqPRYPnw3lMf+VOBGK6sxiKl2Hh+nm6jA/5mMd4cgC1FAYnJ
2B8hUH+jbu775YQkJknqfw==
`protect END_PROTECTED
