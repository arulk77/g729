`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN50k8OgEko9HcOWNofTd2F/g9oLgZmeqLcnhJYUgtPHa
ha0DgdcxfLIMdrIfMNNvTpc31OtTh3GcdwnRUojqp4Ra4ic0n/byPN1j2KHZ6YU1
ddd/0EYLg5K+z3/x19uAagx/Qgi0S5bW5Ez49wTnYmfp4XIoh9hp0zCN7hiWnUN8
tkNnNYU+dqpphY1aElitHzhHiMp/KuxXIV/17rdlBuUUabtATXo7RO3c+AoNnmih
IwMTXJ6S10MuK7+T0CbSwrlEWPBasUCrlWanjry7dg6NEQdBk3QwXuFafWYmbh3C
S8pWIGMj3c8DK97hPIWDEQB7xLFJYC32FIgbbL57l4Gjr6/KM4hLJYSyV8xR16Rv
yzjMt/UPMkV3XJjmsoqWGBJJ03ZO21g+/flmk78PaCbJ+v0qwyaGNqV1JawoQtsW
JkXFNFN1PTAjHXq5O9djrrv8oA1+uezmSjajT67XWOuuOAxTDrJgnJrWifbB2waE
PqEICBH44d/D3ON04SKYDtvNN2QmdSl0Prav7HDXnVEaJD8AOIzVEXCNUD+PZppc
vMVELUInlTQtj8icPCcHb84pSWBgxBhNsywtfGywgq1LWUG2/k5ly1KwHolJU2K0
AvgUjai6YHancUqJQjkKEVXDL+Pq4+YX887ACgXzKMDLvTHuKz0md7LCO2gvQ8XR
ZNTxuZ1ZTY1DrIU5i99fbiIK1+B5b4E4lzll+zHmplq7gQBpolqjEV2Uv0tAD5Sq
4X7kizcZGWunFv0d+1E89rrYoeZkF7Hd9xSXJoJP/asKWim875Q/FsKntUwZDPm3
EFL+G9K1WhObj+WT49nKkmbbWhFgUsMeAkxh6FFgBNUXNy4d/Dl+RR9HhsmVVf9l
aODBEVBuLeMls1vKyGXXHMtQB832AMdUoj2ZwVJ9e7Gz8mEyQn9ozaVjClla9WpG
ryWh1a7URsePuY2t2KWzl07UGze076x5DZxVnpITVy/3Cuu2tjzq2DYOQByRwQMm
A/7i9T5Q+//yWIkl26YIvSXGD7v8EcL4tmXWazJY6RtsvhcZjHgZnnJdgUekhv4h
shjG4OUdYcRKCLikrt/uRB55XslD2fyiyHDxASPbsfXWpagfwZmgN0XwTBrM7Hw1
0g+Hacd1ZTjAZs/1VyukZOUfrNl1vJhpWAUg/1EGNPsiHOv0hkWFHulsh3de5sVW
DQWKuJQIV97eLC5js4jl/BZpoBJdSWJNPRGlPyQ344C297nEuT/c1Lwa4Z3mfy/a
KDUzvOiUEFU2tnJXT6kb/vuArY30p8PFg68t4QJQMUhqOUprkucFjv/IrK5oMeSA
txidEsVATTfWQKyNHmOrRHXkB71M0gcG800/I4IzldxzgByv2DdSQ/af7LsqCocj
kYT1ZtaPF9ZcoUGDAkNi69PvhhAjN7Y8qgzn2xSscjjQa3HICe5ygabUvq82ZYru
m1FhKpeLIMfrhIUoZmtxpQt+4/6a/ik33J7EKkJ9/DDXVAKLeohD76iBehIckWzi
DQfmws/XHGSxaMq7yn+xycFo7iEGIu3DRX0+xwV7CM/Zsv+pD7s7nXNn4fAQWYMr
Cn703iNUKBR8knhTUX1m4/K6bAESvxZgXsWULZp0+mdkSIhHxbwm/NW14ROh9FbQ
EwWupA6wdXipbOSKORx9/+kBthHwRgltP1xY1hX1utwG6XjwkI5X5pyfac+2hTHH
BN+fRVL4OKs9cEfZRTkMDZV676w/39GtkO+XONp0yCkpzdwr0Nzm7fQqc+W4lj9A
LgMJ/uiNxppEIDnD3pwcgQYHUeXPo6aJC43dq+pZAqRKg3gzBYBD0i1VHHP82u5n
eEDt361UUryLfKRKu0EWs9xnKgALkdrLewrBmaQn2F+GgkGCyVokdyUaj5kz1Ck1
ygod1Wmj9niGD/vqq8+rfowenA7Pw2/vTjBA3lf2OtNf3kpopZ3GcxSF/k68azEp
wyxRbyzIy3AgyFvBTeETxHK+iZK9NK8RJ6v4imdgDScB76d3CIAM1L8+BB8gT8cd
MkMtK0ebkzjJuy16uethAA87Pujax/IkeRwk8p7b+IiMeKgZzsTv4Pb5GgKXqwwi
pBNeq/cNDykCYdQOh4PvG+N6I7yuQOpTFIZPkbj/tlsgQSFeLbro5TS+OGIvExwK
gKPYT+FJwAhwxuwWt8+71pn72lHubHBQulue4AaZXVNdB/A65r4jiXk5jFYmI6q9
bIIc8mwFi8gU77Q8lJTpnR0STNoFEh1K6+bdVXRznWn3V6CuurwZE/4RO0YpMo7l
MCRrd+frikKhmYdyp19jr7cUizw/76e9ce0CXJcRUZVd/TLYXnPVP05TkFQ5E6l8
FipGFFOt8ccEwpVC3DwqqZwLWUjrUtc1nAhSaADvqRIW1BobPcJw9NKeUGaRDTHa
S+Z2yVXQCAUkaqCxk9/VSalmLrW8UpCTxOTK3VY5Qr7oE8SaoRFgRMPuw9lWfu0R
MqwlXDZDPk/T5J/gl8rGGcoVN+Muq9/94LW1mFW1BZgSTzJfhvbrA6Cf+/1GkgmW
BCf+1Ra7Otssa5t/620PqSFIrSrEA1lJ3VY6oSUiV4wCMKJwU8EJ7DrfsnmWkx37
F73hr3AWzQvMDNhdOt4qHYcTySvrG1bbQ4m6ih3BZsLcTgVYWr1GbZHi5vAWOvrc
jVg//q6FYg/5kcNMSLd8L3YG0RhqqEKS5XoeDYgU/tnvEsLgYm2Pl/bFv7rWGO97
glj0m83emWYkH5Axi/bnKH8txe57iH1f5PnvuHbx0ez7GpIBJuQhQWSgZJE21o/R
3CHx6/9IKors80Nkzn1AEHmBoPywMkQ3hB8hSFKjrXNl1vbK0vUehe9XLc0PHCxf
LwAbq02WhGMZNN2vtNKYnEC09kyB3pbtah4EQuMghVUJSM5M2pveu5Cj67PSlQoA
rQKtBAG9oQBlZ7Exjlc+7povO9KTqBXkKKJfxc43deIL/k2tjH36sE61AJL9cVQT
b4YUnW8/KfSPbqunVx+WngDJe/gfaSSiS8FiPj/wBnvEG/XJ3jsuaT4mhj5EtXzk
9ACWiBPUsbQrvai/v3NPRAvG4vHcr6V3SEZZuSXVzxNrh2/uzhhML88MXM0+ZX+Z
LWuk5hB4NkMhNTLqHRoMFKBbvWD3tYpbPpzhwXVKQ+R7zZhSGoVqy/vRhsEMdv0T
xJ37pbpCBgU4STfwqMwfSBs8SS3IIHLVKcItXenGEeBohvjI8AD+rRBzzlp2EAsS
3OhI0cX7/qzHlPglgIygxb59pie5Qrxh+VJU4aAdJcELgLjsBru0DWh7e88vHLbm
+urlH8vgWi+ZOhz1xKfzRAkqHw0IWP4Yi1vZlSbHW3Q=
`protect END_PROTECTED
