`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu423CXaWKz6ddhTmX1gvHHIkdO1CQIj4DftH1jshgi+uY
qbZjHx1uHFN9POiAl5012mjWeDCOGzlWBIaOZwz+/t8qRBSy0cNuQqprShw33+ez
+XA71vJ7Mzf+5xA0uqxKPjPanmi2RZwYmByn6ocOoc+7JjHWhzdwuDtDIJq0RuLO
FIy2U41sdiY98hQTtLOS5mCMBjEvvC8/mjI9tq/qfV5ubM3rrZAZqHXabMJSuK9X
WLH5z10jyCHXu748QQJ+WUtwohZ2UZphQY7uQMreim8=
`protect END_PROTECTED
