`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu400hNs9Cr2JxN4Sw5SjtJ/0Eg7zsbZ3/+kUvXWjhjdx5
ixgldM9DZNX21dFBz0qkb61LH2bzjOWWsPhVIFY3jolvpgsEBvax6giMKAAvlSMJ
amvWuH9ZV4lVAx2IZrt+LuV+S6+aO+pvq1q8s7oDaXJDIpV1Fb4QclDDoPDiEAb6
/NWnHOpii5LK155cfMf3rCK3T9i1DR4lvEjBqL0o/7s=
`protect END_PROTECTED
