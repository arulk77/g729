`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73Cw7wR+s1vMDD7gzrrwdnFq5aYJYRFEiZsl5DFa9n9LUM
s6KmUukZnVUJqn0f5qGlyVpBREkZopnc+gVFJJx/ceibXvr+sZIECA9oPYh0eh9N
LCCb3cBT7Z69GWfK+Oc/ygRS9fw+44zFb0GEfexc4W0m80neozk75l7OrSyDm9cW
ANLjcKqzMcGrSM03oR3zPYn5yTuBwe6NecK48381iLJpZb0ru/mo+af/3qWde6jU
QUQKPYU5T6nPYl/VSwVqKCeeGo4LHv5JC8HVXW1lYfoBLaatsGacKBiEk14dscm3
HbUZQETr0f7rCGQcPqU2S0H/ryV17ibxP435rXPtO8I7RogK0NXNaQJqq5o2kt3s
lZU5bfAqUlNweMg7nkE/QJu3XrrMHG0Yu1/FNM2fPJ93cfNo9xfM15k8VBEfaYfz
W7VspdPkJi9HeaFHgDweD6KOKuJ5yXG7R2O4z/T77R3txDBysEyPdFZwvmRGcogF
oZUGNQH219SKAMIiGNQuZgLWYjwjOqnAmDC/WoMAIE2NTiZT5ZgcEsNIkll5SU5O
AEJDZfyz0uDUDPsiAYB8HYe3H5ie5vNdOlv+nUUcue3aPlyRmoTlbgN9roK0+ITb
HE/CBTwjZnM+UkgUQUy9DnaeG3vDtBwjPHr17afS3SXHQXO71uIfi8BJQp4OLiNB
uSDTgL8YAmNljJJ2e14OaRl8+rUv08UNAhA9NKb4d1evuUVCTNO9Gu2rGRnm9h06
xZ3LPZJ+LBgb73ovktNPGPQ4jrX6XvdtGiIuBdoJ4+458RVcnpxoiIIIV4TPUpZZ
IrCSfMPp4K8KpdIa1+W/VKNDlSH89r0QI9h66NoCKTAfxKcgJ2jy+WAKK5m1z9rp
G3XJ55i64bSkLs4z9R7s5KXObsXwSi3XY+09KzfWKuZ8vGBlEvcjoOCIGC/BTijC
RT8peYK1m8RXizqVWrLwI+z9AbOfYV1x3nmt+ks7pnKH8+0Dg9uz8BHVIzdGL9P6
eZCCI1eoRH8HQDdnQNacqXfQpe4V5RUifnyahN+yF7mTs05F3QWGa2EwsaJMhHV2
GKv/5iazR/FyJUFv/7C4OZjxN1vklqb0ajlg0YtDIzFBpsE810Qp8KHxw4hSFQP2
E8H66SmqQEdH9flJAxNlazXxY4PpY5+KA7/cm31lOEWKqKwRmAT05DG59bMc+2X8
Gy+TJbill3sBw9ZjAYCDvFl0UNWxludHePgVCnbbnT4J2R8J1ZwE/O1Do/CsN1ll
wH1KYItgIqRCrYi/CZnsMaS0ufE62CuEUb4xwP53L1IAmGWJybjgRREAOUFy6cpF
5VFwrJJiQAhGGB4TDans+DTByi3pnqfr1/9BQ6LH1IHgHhDEESAZqyvUVkCKHPWc
T1OsPgKizTZD5fQd4UIWQPkOtPxaH59C2hTTAEikBNkrT9xHOXRZMe6cZjKQM6Zs
N5qR5YIP8cjcB571OePDugmN2ZwT2vXoetIHJvLOL8ljDaP5oDAfDzzMKrakU04v
2QQ1Fpq4vcEiWgplMoPNPUXeC42SCuZymYy5rsqGIyOK5zfs5yapi0oYVzBxPC2M
c811dMBpQToX7vFXZxGR59iq30jcoGLWsL6aqm6CyCX2p8IHlU/XMVjeWtovNBpB
auTn8SwI9CGZFmK1dpAEh/lzYRVNT0+oV3LSBjqiN7cOP0Dkl6Af72RvqO0CUc9D
b1BCAWlDfX0R2bRwJrsOA3Tze5L2FYbMe1r+77xe5CN17wRQ/dlpTXbvCbnT0Qxz
ypasAxeXQF8kyjJAW2/Q6mNRt0ACLmZjt+qVoL2vpt2Q5lu0G+ZJQIEDhXm4kUV0
QVlW4bc/nPQIx/iiI4GK1omLxibmn+fRsClyLwroU4JOfvET9OMbuQtFwak9S1Gn
agl7F/6jsqJFJ6p4kKSwIf6f7D+Jmui+f3wRkbZlyOCrAK2lUwbAGXW/ioW7RDKW
Tu2cA/vT3TuobeqcJ3e4HSi0Rr7QDx9LkUHnOKLzDfe85/DsmsDv6DVsbYQnC7XF
bgcU62HocAFWQrcoi1n6fp226Q7v3zqY5Ml59+MtBzVRJjLRs7NYQ8vqSi61KVo7
RcWSai3YCELQWsjtyT0998O31l2V6bbBLc3jrXxxZNe4FZu/WLm05vff4jHeiKrK
m7XTqnrR5CeVApDwd9CXr8mQlOjG42HfJ2G2kMAQdrpxumNlw3d6DgLnpHoki3HF
wRNwU7F9hZ04RI69sw8FL28wJOxC6QMrYLe2gMJNQ0YDV8FG3lUWP1jM/Ombpw2C
cV3Qt1xdOid6MNv6HckAJOOzKrMOja6cIxQuZ7rnibXDdDCqMscGVExuwGnrxe62
rIAJ0x7FMYXJmbCYRgDqXv3WV01FHgG5M7MvIf+Amx/QxiBQlNLyuXzQ7vVjDl/i
yZCN+z3WS+bJ+epUZpE/3QALR6CGh3hv7dzm5u8I3Ctv0Y985+jj9rJ4YOJ/Fp3e
5dTm3LcTFlu1sXdoGs1CjGSBtKFJ/AeQISGU3NCYf2Bb2YWXokJ1iizVKvhUrI8S
Uf+jv+6hEgMc19y82wC29+RVKkreW8y2yVqVVmO1BJBq9YZQznnLCVy9g8n+5ux/
KwmQKqEyknl9Iowt28W/3/JOastTkl/k4atNZ9HafSDRGtkoniXfcoP1wz7uZzqg
CMjAxiEPhleyvs7QRuifPEa4jxEh4smqSOc91zi2zYse/xOf791qC4QfUxlbHJ3j
ITvpmhD3O3hXsSVyK6sZkR4Zus3CVZVZTZMEILjyzYdbl2HG0PRR1StjHI4OL+ow
FVssmtXRpMxOypLeYhTe/h0OaAujrXTo2r5+OuKYuILxBfCq9Vls0KgQ/CFNIOOX
f5/9vBu0n1o+hrf7se48lb64km0xXgRfGbfmYRt5SgWLTk97PI9PaDz1LimRsD+e
IX70eREdhRVkfPYtOG44Lx9+AL1XW0IHHVXkXDjhdL/69u/CBfEt0B/m/XD723Nx
60PZuF3nroFsvBFnV2MD3VZFmj63OOfxDGPf8B8v696jRanDwZFK+Krhhv3La76F
ikPvAcJZGTEMkQCwuHFbut9FWZbVNxTlwGecVWzq34XP8O0qRnjtqSCcUscnDB4b
ZrLLm7y8IBzjLlHztFbNl2cIUQO1hNfOvLp0JU6/MViflnIfPkGFL8esdiaAI/gI
bA7dxrJ1dH+uuD5UuFq1OWKAFkM+M3g0uLt9piZor39FheZk0AlNg042jKR2qMJY
Ji51OEr/HPDVuRECLl4090WLuBZVCKwu0yJ79MnL+9nIAmotnSXsiWL/tWduGmoW
kKz0hgw56T6IbxRwJtKWfQZkApa8WKcmXxZumn/JcOFb9vlcECg2c9xe0Z0Q0Z9E
yQO58vYDqwgzsYTaTUy0/C10cxb0c2evb5jNzIPLUtPZNEuC0ZBGErPeMVkUDbOX
IOVHEOevJv5JvyACJViNj5xD/MkhiyR8M5/rLZRRaKCTo7/tao6O7SHsI77qT6n6
6y3QZ9F1QU54csnI57PXigJRR3FVNbRN885x/j+gLVG4paXHI3uGRM0drwtob6Cx
xG+rWoRqnZhLoqF7VKfnQtcihu4rEA0JiUuh9V4mkumhAA1tVaMUFKb+f7y35GXP
H+uWE4RMhOh1/vS4e028EhN7THEicFZEzIJE4Gdcdcpo/AGB5ya5XuUsWyQKrgTZ
AeOsK8hKRqV1v4Z7rWVqNntrU6/QOjmk/8QamsmIMl38FTmA9ZFK1U3zUXpfJPvp
+D1SPQYRjT4rvma/UvRXn9u+AW6Vos7m10dbZPsMq3/ZLHKUhFDLXo/Hn0A0jeM5
YwdidHCGSljlCBJ6dCKv301EARS2ewpMTWrY27dWynFvdL1GY7NxFw0C10NV0Fwk
KF6DCaUu5SLBw+XJhGqKHB1BLdCbqmP0nCd/zaZHUxbGYHeu1lo9iocuJdREuwN1
3hF8rROL2NKvoHIphwS/dUMAonznvHiVY+xrm7M4gqC7ssekfwYZ/wCZoyKA5t7q
9Nr3rpSflV936ugMsF5wkVTAI+KXk30d0JE41knhWNeBhSUzZd8pxE0cr2j/nuXt
zJh5/CtY7SGEHaKp8kVGseNwE9OSS+hapw/rEPcc6Yrt0JpHkTOshuOmo4plJqcF
qY61OavtIJK01lbp6SkmmSyUEh1Ndf7ZntZSbNlpCLRU6EAf/bcC8TqYGm5kCEVA
gROzM9uAYWtHsfeAFlQVo1wPh61FFiqwlvy01hLRryrrBPHQdF6Q3WYRo60dGroQ
uT3sNYJCKz0R/+EfNkNXBsmrx8zET40lKFqhcE1Yfj/Z2h3gU3i4d+yXHx42iFkY
lC/0rOcBEgh6i5R/q29S16VGwTtD/z0hyK2GyJEmEUSY6u5vphRRd+M8ycM4UCLw
UNGLTlNniwz9tJU65VrPU2VygRHVSAnTN1dbpSsZ/iXq5+XoOMlWWNS6YtDRoL+7
k3zYTPmnlnHTBGhOMNylVDbK1LLdJcyW+dWE2Sbb8sfyEYW0X8+jv5hKR6aVizdf
wZF9/kgklcu2E/c4Aogzwn28ceH7p4FBUFzbwEZSp5YBV3lcZu1hldTP6VHmsUWB
kB0vkZLihoNaUEbFOCb7OPz/2h4dOCVCe1QrhyPYIEIzYgcnZ1hv5wbdrtx8wE59
S/zBIgc+HLb1r4f3KsIcF+kOc72iF5UC8eGqz4EqczlrVyHibzbp3n0oS91BPTVM
uGriMZ1tKcLjx9iSaDxCuHn9kPLvzlmterEUuvYTyVwXed5PxciIDyl6lh/eb19I
KbRpyBKi4urI7BbAiQnvZ+oDCQRLgZrYVEoNawNbnwMASTKYpVNYMANcvGJkz5xV
F37UJbi2zUcRearZaysjIbXy7g5Wke5ZyOWFzBNb4O8cdW4cJO6BNB6weT7OoZvV
9nO7AvF5BcXdR/TXW4mJEXB7cKKZ06gIuAe1pZe2LOK75A/5pTLH6v+RL7ZeMqSn
BlSaVd9PH/DGdSIfdIoRNa9nmhDBNlqGoby3xp53ffPf5wmdkEgTedNIDOHHbsan
O8nZiPiJQLp/sPZCwSuOhpWeb8J1BjvPN9LiuZGHQKqK7YO+os6m0zHYfA6ooD2H
gZzX+hzvlBOoDJh8I+vkgEMkvuNGbJjhJ3dEhN6Sa9gkvVjikh2XboUGyVpLdvke
y03AvINh0/HwY8K4neoXH7UaNT8PAD+OGzP38YWfxgaY02fxQ6+rornngVUoU7tl
DZh4JD6j8VqaaVeyZUA4IRrwWmqFaPr+xd1n28t48hmvTJSSd0BX3prUP2TrpaIb
sZ3lU1UrU5DCTq71CNaxoeQYJUDeHLpAfeVkRx57QTZeowq3QQtBnAKoMJlqAARk
EZIuh3sbso7BUmNxY8j9MTEqeXa/ZbZ8P4cGWynv7CKI/TctL+QUNw95Nn03uoLo
0q+OaZmfJnK5/0xBXdWbadIVrB2S7u+yvoaQXST2q2sn83hq1KwGGHYB9L1JFJ1c
Oni1MUZn5vt4dG9NFh8BP9cGsRMjWNb5I5qmrFBWFx6NTqdd/TulEw+eMp92Tmdi
7NtHuULAal1hQ83ybOtsCDZxk9Cxp1GAOr97++j5Bba92x5It4Fs5xWlZ90NngOW
+VjpBHRcXZJt/SDuv9DRvZ8fJCt44+deZkbtN4LdByTqVZ2WGF1vHE9aW1IiCVyR
dWQvF9IMgrF69AUhyGyrg/adWlNFaAHQMbkz3+s2Wx4kzl6qWc6j4W4BuZYCydtu
ecVvoTBoj4XMsi8Y9vOoGlst3G1SND4SGJE4hRfjKul068dmrN8tz3CtXO9gbsPm
3Q2J+zwHmCv4wlcYYMIDExQUxHtSGqKla4kZcUN3LL8JiPz70sCaRWfX9vjGOn96
BWP1YRwsGm+E7FLB2cL0DFhhYk4hEvHVm9BWufQeDZaw8aFdcpuCPAhbLAEqbhdr
ZMPo2qE4Q6kFTnusrWUl7wu2hVDWvCHKfmp6ET9C73ETYmR7njmwOUY+sA7zD/sX
svGBcEFoOEUly9BHBiLrXRadbgUrTQUfgzDiYq/843krOSW9Jk0GYZGI/N2nfgFp
URztQdZcAN4XQjwXWiyO6LS9MYfErfJbAMOYgKEfiDRySco3SWBUNT2W2a47KkNF
WHnC+c+eIo1No1Ruq4YMp0yd3xg3wG/npn5STW+2zILVJrGzjwZxGVTqmSk44Mhc
Qgb+cKMjov6tMLwJbKi/xVfDlXwuDa2x1VD5FcWS6YvNyf9Ur7GylrTB2Inf+QBl
my1z+1htttw5nZVjIi+nT+uO0b13LbpXBL0oTQU5sI48qLCLh6/e01LRRdYrEe7T
niP5TZveSMw8uwYVyiT/Te+Othy9QvZNkkB8RMAg5JKdS2f0bzlwbih7ZE4uEZt3
S970OjticSlgSAD/ER92VZmx98MTkGML8L4sFM3n7SjLAHEvMEGmqZTzxJt3n0Ba
mP7xPpfj6dTsCN2fWCegB+zxIpTEpoE6nUz301LiKwJyqJJqE85rVp/TRq8YliTP
FeVOG8KEHjnqzY+OAWwpnWKlKmqAymUZ9Bvs6vdUfdIAbdt87NkJgQ1AJGrJoV51
qsLQzYudrbGELogeGY+vRbslxeXU59S0/D2a0dvFcI8wA3lAJVjy7CJ6M26CRmd8
iyJSRC1UsjYebf/1eS9hfThzEX4abiNGJJzCRln/lcr+AO6Va+K/OhhtIk/MsUjC
DOPoby5X92TeLjsf/KqUGtBF9N6zvSUIxkpnMB49HUgdDGXv5XsIoIIfqp9rcH6h
kaw0+1ET0HkUlouhe5YIW/tUtfqHaQdZtPcAoAXsjSt3CsCL7KNEPNYnRSKXCyTZ
gxTNdvBvigw27yNHeu1DWTC/SurijsMBDONe0JEOqrLpFVIhwUwgxYsKlPwRkFrG
ZbBa2ASRETkOefRzlbjYK0yyhNqOHVvxkKWj6mrq6vuyLwE17z8fAm5caoSO1IGv
fAldhZcNVnZcMQzdlCHVVDlcFj4UiAWtpSOl98KDP2/hFaX3mLg2edK5PfpqIQP7
Gmbjq6lZv8+FNJbq0g09w+DvkBFI242KZLVV+lJEeDrwkD16OD0Wg5dS9eJ09h5U
AiLJxYL5R7Wg4kdAVUOhfImu80U4Hx4AgbcUTECxUXz9AZhZQFLhN6XrC4auBIvV
ikFBHL6WtKdTD9cXc6+W5+F1UlLr8CmYQDyx6IFzP1hLYu/Dd2ZppkFwHU7I6CzF
eV/SybGhcwDprWtL+7Yo87C0jyElrONWhOsi+g6RoWAgidnL9iyTBzYZBISvhVfx
UcNmrZ8PqUl9fyIEZGxh7W1QrJcDfz83famLWcTqwQpc/AfMzsw+dx2nosL0qcRQ
yzzXS/MXfxAvqjnGKirQzFzbGch4OUdfDFAiSd+Q/si4s3j7k8gWGBzAQ7Dd7wq6
ru+7GwGt7T9mGssGMRAFuzwrLVgmUvFYVyvKwYXRHSbij3+IiOSaxx6/mxZSnL+q
wvJxTnNg74HEvlE69MHMTUOiNQM22w+58VIrthfijn04ENTDSvv8+rgKcx0w2N6V
S+vPIpIcWxSzQjyYUxxyOBhETnmEmZKxKQScw5EBQ00Z7Uk6ShUW21jSnhpWPsin
tFeVBfqjpMFvr9qEMgcjz/f23QcBbD8bWjH6rrz3Rs2+FXByEwaaM0IZHhc/g/5w
4pTGZFace7nVroBEOwmfjowTW3wfgFx2dT1okJLs+44fI2sndHjXBnLul0ELd0LL
lt8YJ0jc3rnMviQ95l7aQPhveoZi7mCx6AtX2QOvaqOlVAb39baNHDaelEsR527/
v3bMtdsN00lOCeuC3AlM2Qwm+jQghZprehuVjFZ/gZUnENtxrRxU2N2KMX6GcEF+
hP1EY2FDfl8dyWeNhlzFoChIVx0cDgQ5KxpvxPeZvQuP9Y4XE4sjy0b7UDv3XGPU
u8Omzuua+jjoNLhCqUaqFYisdg9STjDng6/6D5u1rkXH5cy67YrSe8B09/9ANkht
S1yIchoupZ85cu4OPa58by581shekRIoiXQVpMSIGBUkDH/8GsvIdQHLDhqXY5Lf
43CU6WteLtmhA1NV+a/Vl3OBp6V0AN3cHRGdlx1DKQsi1MSYno9I6cXXYqPYTRYb
9UODFw2Qy+3cNhG1O8ncZ8Kj6XsxpYmIzQh/yQhv1pMifTKzI36MH4yVJTUBEaio
chFej9XN8+rxqq8HR8ruTqKtG9sAFPfc0EKA1ZSeJ88tCvMlijCq1NJUdZClwEps
q200EhphTuNKlWD28C1wRDhsKthh5W6lSKDgJVjNNrUSfFmdyG0tPx0nFyGfoBZi
1/+onnIUsgdxjCe+6k/eLBLiQRC8PwJIZ2F46hJbTVmzuTtjDKtxUI2hK8vM/U83
hcB/2YYn+u5fdLX2fYgrklJpP/T1fXupgj675kz0yGSxc+7jw+pM9xLLUPIJzmst
qbwChz1gSy2sVAmLIrz+0YXtz46UH+Nc9x8FS8qMRVzM2D6E3FjYntx5JbQNHsAe
q0ah211SMdpLCrKF/+GtpTdaFB3clkM3V8cHvGj1Be7Gg+SIZUJvwM7yj8quQ6HS
DsRNlbMBHSWzeEVoiYgwkMTghNMDQOifoSMeiRcGi4gzqawAHwkMVJU5CxEwJ29p
2dLiyc/MMaiOWXHLKiabxCl4ska/0bVCSmdT6/VmNkWHWhh4RmntOCWruB4fovD/
zI1KzLqfgAwWixvH5h4uB3SzBd+VExjGkpLfVg1+Zcu0LEuNOyvLnIY4EiN+0O/p
4caSwZXiM92x8+ZCkVDWATPycLXKLtCEVhWI9NUP66vJCIow4OyA0pLVlZztM4L6
R84LoIoqYqpa50+EkZYpT7cfcOrxe4iOSM2ouALClcXpOwMufyuIggYrO61Okk+s
zCx81AG4eK5OX6juHlfVkS8noV52rD9BbV9C/bs26nAJvTHJo98tLYIJl7wG8xvh
6EMJoD/M+CBNDvpcymb8DV5SLbfKJJ45neQUlSdRhIB2OSE6tXoh5LKnyIf9XO14
WAu604ua2yepPY6DpujdE6EL91lALd25AQa6M3fxgnCZa+9sHwRRLaftJipmF/Px
P2+1L+K/K/+qN0U+D6CN636/zOOaWQkr8gB8MM5OM4nixAaMKFCKf1A6RWIIa6Y7
Wm2kCd5sHchU4Au6OdT3XIGvhO+2HTZGMIE9gPa4EqGGJiKLCDolIO+cTyCvfuCN
0fCM1Fg877ixEnj5HMhADHmuVCIz/VN/CFVWJe54nnJpG8xFunFVnkCWxWBZNiak
KueL23NZydAtVQLoM9E6rg==
`protect END_PROTECTED
