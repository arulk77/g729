`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
xLp2NpiN/jV1McKCx0Y633Be94pIUfq6OTd+cfLWXwdflUnNMAAHWCsb8upZorHm
UdWlQHs5/YTuk3F8VwewPkkYX9Ylk+KKa3+Pc/Jb11fONERBBxLwgm3vEjgWid9m
HuDdkrFSNcmUhz0l+JMxU/ePg7/VUty/d/MHOmFt8EmSqCcqngR5zpMKi5PvikqB
`protect END_PROTECTED
