`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAU37LFgeFoZovHqLBwAXE5Bllc8AV2l9t85wy3maJpxn
gLL1dWi0KVGtrg3cgur4R49kH7Mp450fJ3hSttvmLFWcUUcGcT/IeJq9fMkGaP1l
hXiQSfwX+5vS39f5batC/bSR3yTknYvfFhvH0Tdtp8tdCQJxP4nv2mpF3y5ZUaUl
Bdxp2rGzSM/2SzrSPzmnsFdutfMKA/PN3BJ9POZNZE1veuYlXiDixSOa6RSd5iN4
SOujJpW2cSUVOa9LXBBMhnBIauWWKW7sZqe4gYlOer0hX5mi0Ua7tG9knLyDA8nt
jnMH7Zr1JHC0ldvzUdZyfH/ksKjQGvMK+/6vwNj/4Q0MdikBrR+2Et4bUt+aI5y3
KAE4i1X4tPCfW9NSEpl5h2/+ayhob4+v9sGc6V/CyoPiwjrEHeB/ZNf3eiRoQjeC
rc2nogh9C0vOVVBsXZmkc0Ppgmcps2L+EHdN3wx2DG9Aed99npbymkB0TIqb+60r
pOXPra97yXd0YQvY6SIufVrdhPOW/CD+ZOr5BH0o7mZpkDzuEubFSyudlaJ+H1Ew
JzxfdfiyD2paS8xOiI37mkI7FO1QPW6zJDyvukHJud4bayouHDjo0yAPDudMNnXL
4+0kvYdUM4nHWhj8ZptF0EYxeCtaJyJi/j7J+3bNzImqIy7vMZE/UgT1SQUWznDa
e0vL6cgyLdJGQu4+Qi3xTU0xz1V434OZ4CA8fAh44rfueU1U2LAMKfRGsbcUHByj
jrXSkqD2/d2HzvoCnVOTKCkFCII95Va4DQ5HW+TpftmsT4FwmxquluBwnpsKz4Hc
Z8kvBT14gbnCX05EpHzBEAO4C6Yh5oiMFUcLX/jO4xlfT6M3gacH1rZNZvgYTTMJ
49cnMpI2LmwZ6Vtch+IY2PRpunBUkQf9BsW6tzLhUTdMpcIjIALih5wrUEMMXNbb
x9yPrkm4Ase6/hrbt5lodjwF7Z1ylQYf43OOWLQXnk/Ey8I12TLwD11VipezANJh
2h6ib23r+dYZaudm+yvWlJE9DuqwihE3H20+d670ofYTe9Nr9eXMzlkYRPtMUEZC
N4GByE0W6MxwU1HArrfoyHrSMhLUAS6FtP5kNGwMg+E8bnOi9PUCOJHayVipNf/y
D1kUBVKTLhnG4vx8fpfsHn0BVNUDKgxZE3mDWvuu9tzdp0B5KrE0FchAWFSjHMuD
9kEn8UFqryOMoSxRVCXEAmPNK4UHhX8Iqfa5gC+1v7GLsaKn3y4ppcI0vQ4TKixb
gV+4jTVmy35hc5vGMyC+Kex3c/8hWwmixswhaneVeWf1aHdaB7rEZT7I+oOPsMA/
9ZcEf6PWjEiLtiNjpkp5Y5Gck5UD+FstB0RQPrifGRzSeTFAONBrG6vXX7pE1kuN
nJbP9eZBdoEf+gsS10hxCWUc/4x7rufEyhV4xOPOZeUnJASnQbb5md56EBgQct8u
HfwXjgT6nFmvyC+X39xXO0dQqKh74SndyZs+deAoyW5tWz1CmL4U5eWnePSYEW64
sCunRvUyQiRX9BA2hfBYxmfZMMmneiOq6wsA+iuX5NjPR/EXZrqk9qydkmJ0+DF0
c8v+ZZ5iM/mpknhTG/DPWznbLwWIfT4MRQFv1UPYLUI2pvxE/0XR/sjO5zvPwcmh
LelYVVVtHrq5trACwwxxTIzJj4PMsHj6Xd5/JozgvCHfwGA788gOIXk2XJVYp0g9
UPQU3GNTAECf2cga2xO/PB4q7RPUD2lLAmjJxVCJfPi4o+joj07DezA3lbJ+o+5b
FxOxQO9AlWYN0fGFaT5ZLXODHKjvPhWBDmrgELyHvBH59zdEthdCu9ys/5tcID4+
M2a3JGJUCYeF+e1Z3u6a3OHsRDgDwLOvq/FQ6/PgPRNHXnHTYyQ1iSK5TUvdEtaT
pDxNJgliTIAa9/vOoLet+E+ORhyuIm40F3yafM853iEDDYQGcRAt4dNuJGkiIIm+
z07FB70x8o2dedHM6ld55Tpif1VgprhQIRx4hAOFCqf9V3DYJIhRp0PuAtjYK9hE
KpdTfWyfHee68tjq4h2XuNfzZtq6W9PRPyXVPYF9/IT3xTNUedX4n02bd9vrfr0w
zkrNAanmVUIWeVkPtO800cVeGcx3rbvU/Z7ErdVvj8dxnXZhUf1GrdgBdSnAQZCW
EGjyYHIpPdX+KDuUY2hAYUd527NgFR+mKHs8g1n49qnu5DuWAQgdwUizRt/p84Z9
5CtCuziisOHjKhlOxilKCUkt812I1kCACTZ95p9AXVA9C3d4QbZ7Nvt6T7UK4hx9
MK/5xuI+V0mQ63Ja6KT9chGM9398cMZH0bhTnZ7FTeNJGArcM1Q++J7G+2T11i91
0Rgug2QWF2giEYQVE1OGrgh+vaRT13t7DZw+qUdUzHPGHp5CKQXVtWJrFBfb2HFR
TbZTiMwsdE10TzOTgz1S250ShNNYrcKOHE8CrUZ7W2k+AY0/XrD1t3wJX8qe8a7/
SAep9GYjSgXEYoRNTrxuUllMWp/bBtBQ8Igp8SWnZ4C2iWb48aPO0SbelystAoLi
aNec+CMsJq/2bqGoTM67WwyQEQeBzmovkXJqVknrzMoslyCWC3bcpQSsLpDRGM9N
f3ulJG0PO/Gj789XBlW5s1yze73haPecjW2OHKJ3zjIiapg0sL3PPPshRNLVnaWU
8mBs8y9Qk1AOhDiEvOeB8P9Wf/SpoaKhGBGEnBOkype84K14ocvHl7wZQpES4IDb
SIGENbFpCiNY8KLcGaqJvnTxBBnQ67xv/654pA59Eu3QlUb8/GZnXKkLry/4Dv3n
vkXztzT5fCEGu0SLFw+B9SGGPgJ8smsxp2uZ8/mb1HvLoqZ8Tvh80J/MU+fMISJh
9sc/4bAmgXLB/uLhdt/jMR0O5jPezbnT1uI868JSPRI0NWiwFXurn8FL5KNJlGU2
FrEP9MHBx0B3ux4flcvjmOk0ENtvDFkyq3KKoxmxQpIJ0UaxJJ2IAAVuEJgj25e1
gpwFNCwELckEMaDEb+K90sUf5iReIPd3JZjCerYofQnORnQvcGNK6OxdMINJCMVq
IbptSSLgjAxBW4Ohwb69H2OEjVdC/E5K39sAV0Us4AuqVkYmH7Y4Jb+8eVeCcTF5
M8usp2IT0GhzvDhvVU8EBIiSbrgvbegslrfoytmgksxHhrkSi459VJk0LamTB1h+
Ha9kdeaORucHdH1ymKLZwHkvO1UiO0WUQo2uKXsAApxl/AzMy1jZcYXln0Xc42iT
oP6paqAJ1u9T5r4t5sPsC3omSk1pmX+++914nvgRbviCyYSvJZadcjeTyX+SKOKV
/UBW+WyOJRcLRwlt3aPvihOGPR+yW1eHIQfjrmeYy+8r5FcPqSZwt9sfxBrc2Ob4
3jQHLDTv9HfYqk1fqe5NqxsnSWZJHR5bqBPCPgKZ89xmXr2/JjyGpnN/bEZLUJHQ
MWI9X5neiTdg03VQc18yOPDWtzFvIM9KOs9oB19nXZ4N2JT9Oj7yfzLkY+/b0gX1
5pFb0w9fvtDZLGjPx3ZIdYaDFM0Od693HLN1whHOfgg5Zxdm565MfDz5o6MNE4zC
1eQsH35pPuD2KxKNOeNWqHKoIfECa0qJCD3jmcydigTv/FtMY2r0Obgz/zYYZGp6
gs9vQaHT59hYfYGVnq6Zon5F9PB1AdGzKDJlx0aehSgKBJwumh7TdcF9hac1wEGj
tFxAwMppt0ZYtJvWovBFGyyoUyfGL+32l5HBcfdY2mmcb5rUyFULNqsHSm856/Ir
EYfqKN7M4CYqGw4lVfN8KZZzH/qdj+bNUwvl9GcgskDP4eH+NzFxo7t1Um616CI5
H97rm2RBdBFwKXavzgJrAbXslPFTBqyzbf09p+uAHzkHuA7VZ1nCdXBriO8dJTqg
M8ncyJ+rWjW5/p9fvQ8RqVEsSyphEthsIq/AIrPZj7t6VYDTD11rVcDcvXUv7EXB
8zTMfRA2iO/u4ST0/983sThrzwnfANeHXEOlAy8VqeMBvE74oivZz2KGYi28bWP1
wXcD1ntq54wi6XbIe/3qUkVPjojB+TCTJpCc2z+/aHf0eg/LXewOg9FB7GObKrau
4AMstUMe6fAKSUgasuGO+8NjtELINgycoLlusnMGRNbkliJno2/shK5Q/tOBr6eX
yu4puagcGjzoL8dVCwxan4jdGj0lKsWQOAqIzzXdJorqUXNRla6vIzho0diySDeo
R+JNThoAWzhkK8nhQnGjyQWj0n8xA97zXrZMhyUHgn5RwNOPtC/RtAzNaPtTpkoQ
F9Q4ndkO/VaK8WGFK1ERBfZe9/yyEvMf2+a/jNGtFJdI0kPoNerKHz/8yiAM8263
gdrzJ3tXFGTVA3Zh7DldV/5SFE7RLvTDq+T1lOcXSufj31fpgyPRMXifqFuFHRYY
YN1sh4q/dux5wePWSShodVfztbi0ILFWCdPUscP2V4oqyHid2XpXTVVVkkTMB7UL
fOGwPbcT3rX2YlTcevUQr7M0E61DtFBCLtcC49wqNNvXvtBHDdUxfdl+8VTx4CFZ
V77B2yp/emGdJ2Zgyy8fY1m+rZvRS80AYbypig2uy5h36+MROF24OHWgccipGQtc
3/A4FlaBBcJxpwrXsVShRjDqFuwc8WJIHMLMGpRvQRUzyQWQBEPUTZOV9OZs4sul
cU3RKkB0S4MxTXkNrfdW8pXJTl91LR9SdqmJzCo70gbsWsO5r2OqbzQklC3kKDZH
vbuJIuA1k5tIoGa1g6O3dVlFErWpygp7ouWrLpc9PH0f4ZgfizfHoIJB/98PE2Ak
pBR3ZaFtLSUn5Z3Wk0AH9hD6mymEJNCeX/O8Coiilz0iIeSGGXsJPukHH6ac6dK6
t8AUcGM8D7KWsG/Pz+lF3Mk70kXLD3XNLr0tLovF39MMwXN4R1Tk9YnyF/7DIbjt
bRgNwtb4tVMEQSNDgDIo3mpAAdQQ7+Ce+6ism0kJcF1dGp7u9XbqJsUKKV/1mj09
dCz44dNvIPmb6OCCa1KyK68+k5sSOeYfyiaaF6tNdV4d2s+ldPP2vUzQxBkPNNbg
v1y8EYqqViCZgDVd4FGu6jyyB1Pxvc5tRmUv0sekst8Qn8N53tiYlrT9qn/8VmB3
uXdkSGV1oKyJORgsnajNGsE9sPvIrn1wJVB8upIcK2tNZshritOIszxMSDoJqRAx
DRIiKCCm8vxY51hZ8Xekq3aWXAQPTubjXf+3H9SIX0URUdd7BFibsD1lDSmKmSGC
NnEJBtWUKPM6XlCmXagYzyp/XBaU+dWPZV99zNxoJnNMJdiIyj+L6pCnWQzZWMfp
104jB02yUDRGDotEe+qasp6ZXU3MnGo42pHoeKLTN4l8NqdLlH4DXi86PZB9pG2F
CvIvyUgTYcPkA3NkywGfYXGD64T6jyBNdYoq0Vk+VL9JGgOYraexwzOI/yXvgjwP
n62BSZVXYdip91Dpmt7wFOw4ZP72r15Z/HKpGpsJSxSM7QGE34G2MWK3pafqlV4P
XrzYbVq+vO2cbhcaItYxkHF3PDbllfnLiBZid2ga/5hvL+dir4g7ND6Ylf+UOHu2
zl8A2OLvifCEHnoSznSzDEImhiVPtYRiRl9ur79kJu5c0PeqKIgVqsoUCuAlBlrz
GunujmFK3gI0JbynKHZ9LA==
`protect END_PROTECTED
