`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mkWIkUzW+CxA7V+X5F8J8pnDEEKmLDrwHSrWIr2lc6yr1NZwp3eMe3+SC7Wb68XP
xKZ/XCLWIy4jnvra5QulYwExOOFPkrUeFw8+gCqR/jVMHDytVDE0uku3WbXlRf47
znbny/AhmKalGP7ZUI/u+8b+r7WQkSsK5jOIPD4NDQGpwVyMWxqoBMOg0RrS/ptE
KDlxt47nY7WGGkUbCM8peBErXD32vPexWvrXGdcxOdxoKZSIpqb47y0dpB0bpmaz
ptZSuyh/4Rd7Tu9B+voP4m10IEdV4sCL3nMgjH2Whi/mIfaQHS03R4gQoGqM05Fl
QOR9UY1sLsQm36r+CQsbyUVD3fPc3pTcWV42c3vUvss=
`protect END_PROTECTED
