`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
z3RLqhUAdbi5v/dq8FrVjxqkTzwh34oL3Yncpl6JQ530LiTxProLMliYXIj5zCy6
LWJz3mOB7SIcvtfEPo5f4C4GXETJTFq6yr3llEA5J3z5hc0hg1xiAqZvDfCQOubb
ziBzVLoqF7dOL8SFJ8yak43iXHQt1emzeeQ8JuVvFE51xAy2w/UkLQWrVObMHjfH
98yoGicXIMdkn58x3MVU5Ev65cgaqqEZSmPDDJIMU+u+ZDcdF1cFBOCX7gWhg7ma
`protect END_PROTECTED
