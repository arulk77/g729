`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SXf5Q3HSNjEyuq6+V9h6p4AepCKeg6lIlmakF9U557s6
rXY/b8BUB/+KLlJX0h9dYvEekl9h8CrCUqd+8j8qJfs+ovXV8ZChM+iAt3vJjacd
1ZOxDee3QqmwoYnZZhkgMtqbrKFII9uFcYPJq7g4CkUjjFc5G6CEoyJeoftP8I7F
baadBFpOtfOuTjyFNtyPTqyJFBbOByxQMi7mlPVRG0yDQKvw6SO+8jhFrA8dC5on
bQmTA9ZO/ouhcywHp5GnLaziE15l1XNtYEyEBZfQdyp0VALSwXh19yAM5H47+lFr
efSwBNND5xeBr7nD7ib8AdUYFKAvlxcx+cia8pkZg1vaS2AVlKys9Pl1nOveOa5B
WKzPOXA9Gci3O25SghqIBltOMpdPjVaTKJhxY70J1ctjOauM9BzaG/IjPrNMlw8S
iOgfn9XIWohh6dqKPRjY6Jek+FBZpQwv1uPxrsrZw+mUK7n1IdTbvGusxR++m8dm
0nxhgcQUOel6XheoPTXqIV9HOCGcy7ZKzIue542yFLy0gbDkeMlQKpMqBgeA8ixb
Rjcz/3tjJNKI9Em2OeFrbNA/IMUvjG6kmnEi+nMVhqiAcsk0TOUiWBAbttyxicoe
eQfABqnIhJmiuul3aCp4cyHfPE8nHAp5DPuHNzKlqC/IACBJljhyWrkwLoApFYYT
RxMyPMuqv9cXulXMfc0bQlFs7XkTAkRjwi7cLyYB0bfZXRd/TxFNbfnpiUt6eWT/
0ZAv8L2aAYDEYUx7jTT7ohAu0dfwrR2X/VQQFZ6u9W5WP1gkolsVeDBdeIJPSeMK
FtMLSVAvWTbgQd/xdfGIOzenks+cTVCEENyJtqDeWJYkWUXlPO7/3OzuaCHutC+D
p/xwjUiELB5c+wLRsMSDBbeXByHzhh6oCjimo5TPJKArJZGKFT5FdLpEytaskjOh
a0K7IJhJJVpz/u9dMkmODQH9/NE3BgRsc2j04bGXBZdpXEWkLIXHe1ghQkQyAdb8
VaplI8smgwhkGqPeuk4/B6Kdib/VF8f9mCly7+adpFozUAdduNwNNNBLzVASVUeq
u64QpyxAe/W2Yi11UioDuEMIqSvIi1YTfMYhPl/izIRYUD3gDDLBefG4LlZotG8n
Lp7yKPPLDMJ4k3XZqnc7XiGVq6JsvyFv6Lv6aqYpqFSmKO0Qf09fE5qLkm9pn+rN
WzC8CzKeCaMllanXR2JUNu54M0JYInev2gU66uuDGvhKXcUFKsftRwYCwjz72ay9
wmv1kNmprbQkvlrVdB4NS74mEaXcL96YSQ6clrj/NVMEeccidk3yXggC+kkuWE/q
pBaHvXLPg8lxJQHT/yFxZMs5Nwhq3uyrkRXjuHmO4XBhgiS2mOy0POuLIqNxBZI6
1WknfzfBegnrvh+Ec39Kd/I6xiVkh1z1xk/63hPIeftX8QxbBaVFyalfmm1KTiYp
Wytcq6GETAc8QYpwl0C9NgIAnhRTyEFJBTJD+HBeslsWf5jUE2PctOLXxxJWZNxz
IP5sYYtfJB2cugUARklnIsW6z+jpbcPCPmjMX+emGQgV3UzvoZoGRRarqSfMdzW7
j0N524iATrs+DA/mK1arUUIE1w32EwsKgPGwVEjyjZVBVgXnnjxgogwGkPyhH+q6
79FiavMGxqi7qFUTyi7ctdwhQ939Eov96+RzTVS/s4KS6Pmf9AFVLm+LptWkHOyq
GZcD0D+6PjMgWy+12XIGLx+f8Wq2Gy4eHGYeni8tXQNNYKHXfowP/B63IprxwKxw
y0IQJQ0YMoyErTl9aM+7qwsdwVkCbO00VURWeGEG6yL3mO/KC6gCzMAFbGoi1XGe
2UcBn+DMHNzcb+MkqD1W32kTcHPDDO3upuedpM2N0JT6Axn2+7Upd6zJR5mXZ0OV
oKtwDkEBUBuJUXy0M4U8hVP+FMnIfkv95/QBCxc2x1dhRX/yFSudFcqMwubx0cZR
QpqDeOBRtRSHxc9zUgUF2OE+sWiIa6k9ofYTtT2L/NvFJenxQMX2YeZykA0YDJMh
PAi7Ch8NHcYZ9sZS2SHYLoDbNV0DCr5gSaeubY7igIcuQhnV8Hawt8YQmHhlq4ts
iV4q0cfrCoSO7sl9tpXLn7tes9x3KaQQcTuGxMoGWA2mqSwxI/WseNcv32dwryNn
cfeFWplLx8l4Ju1gdLiVWgyW+vU4In4vCUcOcnEJYydfFAY7ti4XUYVJAiTRGiPv
+0X+eEBljJQTyt3+PyuuWDJgkOE02y3/arBBN+Uv0wXWp/TwRskdQkmX8bu8JY3M
TDx8YSTKmtUY6yOYDNHym15WblYl7vHR6Yyk1AnW8iLVHUlihzgKK3CHEWOQdiMK
vxMujvPU70Q7xqvRQChiT4VLAkNeKbyiMiDc/d+WHHwUBlw/Zu49k0oiVpYViR4O
LTvt5BV8cE+Fz6RlSEHWI2dRDhM7YO9OuDqUujkYsPHULuXWhm3HMjMdiiahv31E
lyFgksIs9tGl12058O51vwIMorQaCjIixdsYTONPakHvreTW642dVSQ0xWDV+fJT
tTih4i8MCku1FZBYn8TbHdJnJ7SQMbBjBZXdm4BMllqEalyPMy3ljKDHUIABdVEn
PjQNvAEGClvlWsPwVyVlMWZ1aYE6jo8i7Q66hs/KuMCnkpvrtdFepTEWpwsMoi3L
JYq0urDuFhJZ0qRGgdvcJbavt6E4OyMQI6EmSlNDu8UOVSSmr4pRb5kGIMlNCDor
0otwcQsR1dcIbYgmdDkMozFuGcv+d9xd1xSu+RwA6Mzi3adkKenfnVRfuktsgz0o
DiaquFKH+jM3TLxtluen4wyIm+yXDlb20n0GPbhqq/Z5M/Rlei+j0M4PrMA7bKcM
6+5AKGEqo+EiyHIBRSoQwrYIwQXRDhvsra2ckDM9LjL+/ulXuw1/tWGkVv7pAecW
Dj6FwCoSUlaeqtR/2cUdfU/BL8iFWajYJPcldUqDniYWKHY9Rk9/S1cJ995WfjjA
GzbHuULhTY3mAgyfoxGEkmbe5+/ExbikieIScssJBP/mpMV6+WeLJCIpEESjb8BC
+tr9g2x8gEdMjVIax9VBFNtEEDLVdNcNefRWiVaXDB0G0FF+5dxDOA2FwXg9cLLc
O7OqY6hwYg9eyqRrcd99Wav6QoTTV6p3sWFUTzk3TocRiIDGQlKRh2J+xQwZZwvC
K2hptKGe7UIy13imq3abF9wt3MauzoeoZekC3XpwrMqZ+Ui7DC2hkoyBMo1UxNdx
gpG5kHafxA/WHafCfwu/MmcuF1GSOdUs2uSNFgfkwhQk9PMCKJzQr8JFH1y7DM2s
j8yeWr3iaUghMyFG+6Qqjz8glz57iGbzT/+6Kc1os0wq7DQ3kLsxSLj0Z0wemJCe
YYVtqI3Om2nTP1MZ5THKUb6bTRe0UKH8NyF2WFhwg80hQMqweExnZc0QKFUOgyjL
AIVoleokI2C2AfjHu5lE4UuxFHvde8eq0WtqecU3hqMH4vaq61f4MVZcVSmaGNws
SGsfHpGyg+MG3bBOvua5PPPqzLuVF/8Md0eJNdM87Vnp9a9sJJeQ7KrEHHf9zZys
05bsaDjjenKgcODLXIRkSum2w7V+JqMELLQxi2RitlGKKjSIeQGt/cU9qBuNuMfV
qZkTM3eSZime/Gv+rlpgsYtHB+bkDt4vV5/eJboFFZ+DY0n/8frP2VAynLreVnqV
hzIJxwGU8SBrBbTTG6FM+4AwQ+PPizgrdqs3jobxuAibHuq0vxbj6c0YvuoOdzMK
o6D/jMKsez3pIg54I12DGq1NOhkVfEgvtXYPS2Qy7lagy8rzGe6cgu5ywCtJbDpY
H0EiaLd7zbkAt20hUwpEsShQK896TQQAUEuXsi09IGwtcmZ82R5gtpvxM0vDipdZ
2BxDp+5g02nAEP3t/RVVR75dTz7USb3SgXB+oM3HFz516t/tx2ckpaC9ceMo1stx
OlermhNlaUsKz1TI8c+OYobefTsSdDuONrlzonNLiwNbSrOL/WqOvpppNfQ9Z1bp
JEWm1Cd05NAghLMZChpzUwzSmaA8zIezFym55noKn6CrUI53REBP6remxyVrAq8N
vqAKIGNbOmAJ/NEOMvUXTdRvOgX8XIpmHYF6WLgstSqWnJRy6kNgjwdcLWy0nVs1
flQcWOlMKHBw1OmR6Lyx9T1jhHXZyMPU4jD4kwXpKa1cZsQWoMTbjcs+nNGSOmyx
ENdfzi6L/vIlZMMTyE5P5UOjSRu9WuFAtNaEIQje+bnqb+ldL5bdP94EssoXSn8m
PJ7D34XGTgfn6fVjoNfK7Z8zHJofsIfLMd7kt6PYog+I5Bx1BI4LaIM+Q1K3K8+x
jeEnDTEHr/tWORImNFeqnS7B/d/vCWueSm2djr0Kj7gtKjBQpr3omHo2mKPTb58s
Vwv6G8uQHSLU78/j+kZghfMrlHKjvhs2dN6PDYU5V7q4yqsB+gUQfRYUDmmkmjBH
lG+g2mY7ZzRqmYc8yr/e4DJk5spuJ0KxeGpmdhaj/oLxT7YrgVWLtCdO26u5tQQ4
owShEmGDIizYBxn6oGHmBgpyJZDleje5WU4cqOvvk5+9xfe1dxMKJPTN3fNHo7CB
85xXY7qM03qdtlGQJqqFlBO51t9wNFYxO0AMsswtDJmyGZI10lkhJippu3Ze3Qqu
X2bd+HBNquzt/9lIt0OdM5VIdS142XkKjvlKDJrq2uNJ6uavTRbO5y1OKQW7XUWI
GGJCqZ9oIHvCweTkAWE6FBF1XfRKARZJeOzheidGVI+xzF2Snsc54CML6k6uGN+9
5g8Mkkbxa2w5GTxCKke6KwXHtAyu+zxfXp8wsTbo9acksE7tuQRJTnOJJ0qi4fmT
8rjY7u/fM/gcGbaXBPKk5icTCemZyGMXxMwXM+8WmfFGp8u6/Oq0tK/bRTitqqkS
W+K/mJ1F3ex1j41vyCeG8DIGJ9TEiHXnFX5A2iPi4sIu4e6942s2VlxEyYFIFsrl
jNYz3cU3MG2GrVkGdu41Bott8OrnX6B1zzEBzQ8qguJbRWRAoOLryg3QvSn6W5Wm
KxWWJ1ZKk94NREp+wgDMf6aVoG9MfOWJeBY+oC/n4Pkop4EYnInu1X2k1kowomGD
DImCtYmKm8H9tiipoWQOh2shvTW0DnCogqETJ54Vl5bGFXALUaUQ+aaAsE0+nryK
WYen0cHrXG6bD6Wz40C+UbQr6aUdWH71y1Gfnu8GRGAiqBETQ2eyrX74bP5OHWfh
unyv0jFx0YYhc8RSAjQOwyTh8QvBFgDlNgYLxuSJDijNqoTaS254A0MN330KSJRM
m/aTVOcnKbqDPte7JMXWrWECeoRcMpz3TCx1pYCLAGPubRs2evwSgRTayGeF3nEg
k8OsCCLNpwiHdU0bK9W7LB+VjIMVFZALmdlV0+WShvngAMq9uBxImYGZsAghWOns
uYHzE+xtXbp8kvXfwnj4qkc8Nso1PS+ITEk4FQ1F/vmK3agttUrrxLafpvRA8M9x
n+QW5I7e3Z9f4jmj8CgF5JgFSxOTlkUDSetVNuMK/fQW8ej1Pf9ycz+fEFU4A8SP
4UxHz5JDLZxtn754arGYcHFQvJ1eLPpKs2YodxOO6sgnPd4MoWb0Ht3T8MUyMjJk
07i2HU+H6V6YzU/JwKtcM9GIL6WYN/oCRLs7RU77SqUQyQgJzanJCOB6yzjiYIgV
4OqJkzPT675aUKFlOtWH2ebEy/t6617R6dgJO+QNahnfd9Ox1hGsEnY/ircjiyCB
rXG7gFyC4Qfepo/ZnZcO6f7FqB/xm754gI9kONSaCfd/j6jzbitW+stRMPpIvlor
S978okbYceKca3+eF/N4pwUj0xau+GpCZXERlqgrsVzaTQvj7jpBwiZIbw8us++m
LpkZGv5HysCo7KWGi0io+SuepKkdfAjet3/0TiBxuGa5q7lTKKnSR9W1EaSjlges
WB2V6FwHg4O0xoFNwOWqnC1LtygBJOMp7bn+V3unTV87WYLAw+v4hbPd8T2cA++0
3X6SE7FCL1cJh87KVk/6tjkPoY0vFoWkTe/VNvKM4RGlvkYOXADJC4RNm0QlSVZW
+WXvg1wZWkr6BOQivIoCqPoP9lefV3zbdj8HDVYZLB63WTSyRt0y8VWuJ1+RIiQW
4D13WD3cy/B2Sw8m9z97ByFHy4MDCMCwCa6Hd05gZ6WhPZQrzyQWmQ7zMOH+LaAC
jfgR8h7kQYzl5sERILG7PvTI4dPsId9qFqsu9A/QSoA6x/kHOqi5afHpTaU219U3
mR6v6Tp/z1Ww5qYiyvSg736k0Wzvmnibdj0VT1AkPtfQwERbXjL1qJjtS/959M1y
aOaC8JBJJ3NOhi6M4v3BWaMm86BUrEzqSYiPQFF6iwaauHyk3mKacOY6IWB8Iox3
v2p/kJIFl6la39tDfogUPchmh/FCO/pBa63c5EfUbiaxNs8dUqMhh1RkfLee+uxM
XBzVGjCoQ+UM23Lx5N29QaRNsXSeczs2A9jb1yLbQWmaPY+I0aLawv7XqPcr+GUi
5vW/aklSFWrgXJDlKLV2LqVLeBO6b/TuIj/ttNexxyMorG5yf4/9tdrNHG3b+hYR
BYR5EgCup/p89Ml0FBjyHvr2rCM35cG1kT8S/27BFGQ95I8kIGRXbqp1pvorOlvf
T3TYMT4v7iVTMJgC81z2UQm1tF3e+llEMy/kpgc8dp1e2ng2t4umCJDpNFu26lvT
a8Y6G1yrpmBzlhgYjcp98/i3bZNl/JzddIT6YPpvOd/uM9wlioqdUswJJYNySovD
tN/n4PWgvnz9TCLEITcIvOFcES8NDxmcUuqchvtcURE6UugcanEoS1CaXZx9didg
3pUf3Hr66p5uC6H3CkahLUsCRjkCZp/cSV1eAnmpe0u78OB6u9TG2Du63DtwHG29
0UQPhT1hFPfaNN429iqeR/iOA7A3/0nQwohOmFFB8K3dkz122/hR7WJdP2mkBUo3
cZU4PJdERvN4auHHLTlfvvvrQzxXnHQHUyI8dAGQ4QYCH2TdxCR8BXjRmEXqamX0
ywxZqELc+fu95Akq16vjwcJZQfGUUaIwhNsZ3yoZS0oZJ6uV7ReUMRqaihtjBdv8
ejE8SVXvoylZz07dxYNtsZcjiCcqZdwdFMyvK8HcaikBHvcpN5PI5u2KEOlHL9VF
ig7RdYbp+wPPfh9nC9fiTmxJ+/j4hXR5KOjKv1soWpcxmcHavAg5otXQ7KR+Ab7v
PnFw20y6pr4wAPS8d1iPjmv3XHvPyaFu3tFKIkA9ZXY6Pew8ZVT/wdXPg75wU7JN
upwxyhQnZPsClUqtx2takl+0tV1kzs6pDJ8ysPCYTXo8R2SIDHMDcjWZPxLJYbRd
q7HfoYkpVuCd+GzUXJqDBLLa8j/HEJWk6TQAuZ1TzJMTsTGthSpBklQ1MxJi8mZg
ARPfL9fuLODziEeCGBEB/M5vdsHSa6cVoSmrtv/DmjSGaivI6KNjOZER3xULlGKq
10nJdrB/M9wJ22qo796FWpxOTC4KMtt1QeppwnGzO68Nlb3jGxUuTzd6EXVL/CSk
QlPMfYd+ZBxUwUy7Wby4Gn1kr+JK8d79dglOERB8gP0xK5rtsY8a/32g92PWx0kI
yhSkJNRzhve/tSQ2IcMhObFekGs0T2vslQr1BarV+YB/2MYBkFyFFIJmmEjKPrbg
D5hnQ5Kp9g5kGlstD6T2g5g0Gi35GZ18SpZJ5/8ph05yrnjyTiKazPZoYxmRynIi
bL2TVXXADWARy++I+xFmOETvc6A1s3eriB1UrhRHunn8UUTp51zD/O0toAq1Wfpw
7PKOeS1enbg8Chz/u6NVhEYlHChQEf3Y+/REqKNU2XwENMaTK+ecZSkt1s8HMNsi
SqVyJD1Fw1gjYx2F+F5RZxG9NQLF6XGc6pEN79UVpuknTxfVt1YfL+8GkdUyReJV
DOVyRkov915A4l6QuwMbM+nUz78aqXQ4NGSDs7OOXE15q8zWMeCdAHR9NFPTloN+
3YH3XVCfF9GkkMAAN5Ni/hCF1xidhYmratGJ/mHAEJVLUS2VkxNB/8R80hhIscta
rLk6jDf1Nf8IBj7uz/Ty5pTEahDVpynNzEmcTuEquJCaB1QKy9BSVmbI5VKi+ADI
5ADgcHyNi08vfFf3nN4qQ4vZiJblj5yfMS2gH2anka7ZXOrcHZGxILAHh/We7Kq0
FBxpwO4rBkemGqNo0iVKpVebDGgeWhr70+/ZzTz6r6VKnL+QeeHeafWA//2RVZqu
z9sMUnNTu177dhAHZC3vdSuhw9hSDcq7ekt0IMbPc0G8D5+XyHwy6P11zPUDOWpc
leoTPcsAieGtduhN+pAHM+e4inU0eXCjWcUCCpclId2zKmJjzv63lOWxoYB5ZNeU
bw7e+QjwrtYmOBms7kNtkZcvoRBujrYuwJs2dUArPjYiKSgoDKfrRAIRP5nyb4JU
lIbocb/FhOeD0uUTxHsJXa/9KWCmlKjcPpaeZJD+DcfeCdM+U+tqOhqMAM+uUeR6
rE6IUtmNDP2koVQBvKQht6p0+TRuz8s0bVWfmiSzoen+qjb9iiJRW+zIaaFy+IIK
KFhq+DxOFpG3CO9ymA5pPPOdPMFX8abyvafVU6yw9Bb5ChDAaj3a85PyMRhEkdDN
HvCsMFUwRM66z5YoWR3PwZ0z/2I1s2eaS2cUTW6WSYgu7mz4bOkRV7Pepz7a1kZK
Xv4+eWes34niobnSKduuZkaPtizpkjBWj+/fG3p/DWyjF4T+uXwm2yRJfi3M1b1g
zke2tPXbhWQv8DRKARLtXL3B8roeEZcIkfUvqVC10D18p/b2DMFO1jk/8uYW94tn
hHJCgdwpeqlIbjP7BCaINHhaPHmBcPxHJOESFNcUSXiSoo6YHMObBvQ3lcoZQrny
hLF3dJefJfvsgPuqV2DvRl5zEkwtAvzUmaoATmMpZo9cpliFzTJ9iZ4VqW3dXaFv
PAv+sNVymafaPoEBjL/CHSw4er6bO9jrR2UydsLM+w8FFg/5JFhsFa/8xsWG6i7B
7QOZS2PM5KRztiafcjvgwbCUb2Vre/FL5AB1N5egPTj2/g7DrRUscMmuxc7Flgn7
Tu5ITdzXtRb+tW/Pe0i9SJI1E4sanxy33bobv45Oq4WLsZFYDZOnakrjvpS7ZKl1
VkPzi6E2p/bycafZA3P86y1TMkXd8Mzx/VaurfYP3yjC5FqcEq+nj1941PgrH2YM
1JcCBJeTTfu5nzP6bgWqha3DzGA2quOjyXK7io+9kJAMHajHRM676TPXxMfB1pJP
8Ez/yrAvQBdaPPpJjpIVfxsxEtfmb2D9CBVglKihfLWF9YDAcG6cfmpN8WrMB3Sm
pe0pD4xVxV2aORTtSuI0+ywFn/AJhfMC7Se/CFrZkFNYAkKqQKER0gf9YsIj/H1G
Kpl2P6GPCaDfFr/m1xdVVUfhN/ZQy8Q7Oazwn93d0xF9pHrr1yqTERGzY5yq66zr
gvKPWp9gX75La/CSJ5fsod8rPPjaMgqoG2+BP3Gp8vd/WGW9/PnXkOPt+/EQhBJd
IqlU1qs+d1XJx9IQ/JGyHjHy00yArVfnoCezJcF3sAi7GlO8GeUfH/rZQtfe2ihs
7rdZxYwuZuNIchKeaP1mm2zP3PzQWwkz4z4WPqgcQF+b5um6pgjU5UQuiOLnzr7A
Nws5QxnZ0j5WNdyqh696dg7px3LGWEL7jPTAbP2wXaoVjYnqEHvnHqkJGHAaN6a+
ysA274nfBxMMF9oKr7ZWDXPqKomcp6VZZJpHe01tYYiY94Kicv0/dKqLLt4SrS2I
+kChyu14z9e6XyTOcF1kiBh/vQssdaaewJvmzhNc+SYRrnrTmDIjM3jOc5baIN9P
RKG0CFO5eLw6JnmT5fdy/so7DzZwpiwNFhfR7e35ITFoPLkKBclQY6u4I2OsMQ8L
Nv5zIC+Pc5nyJxc5GRJ89P5tfWE+5NELYfgMxYLAskR8/65O6LMF1h75bFvWzlFC
iWU/w/BlY4nSY43TuCLP+OBhuHiHK3B1BU+DW0iKkOTdH3OcVnlJk4OQH/MuqRZ9
Yk6jSVlxtxktIYQHcE/AjMz3sjQ1g7a1S8G6FLIYIUcmwXmH1UdNNYvg/SRJIgFA
VpVxKbxFRIlZmNYcnKkN+eg+his+ME18Qngcsy8kKXGB1P/zNmfxcvyfr3aJ/LRj
NtmVsDj40q3DvYFPqxEctZWYQ9FLAOVLDArfaYZKbC5AKSSYoP6skKVHulgqCvtT
OBB3A5Ayf8Z0b/wwYB4tuwQYJjR8EpX9GLqZi7W3hlpIr03pMDk9tkCGA4njU0tw
18Es7F+A1ThRplWiDOX1CsDOGYvbjY+AA16yWdK7Fd9D3DU30bQ60sLYdoohdOHh
q1sHF/zXRmSAMxBWEcg3GGt9yoDNelDMriajdmeadksWs3BdFZNbT10H3+kuzh5u
b2NrHCkOsMtHJqoQeyzG70TAGjn++KY5LU3chHgvtqxb7S+MLAMUfFR0QoMmPmJT
Do4pi6Pp1UR9V0EkLFImqqh/k2AYOLKAigtGho/LviNQQcGRfLAjHn+B/NKCpeqX
sO6z8TPTuU1eMZgwa0yeleYuG+OEewlNT2WBqIS0PNPMndOSOmo0lAuJN1kXltkf
xmdktMbfOh4RrwwLw9hkQvmjCo2Zh0ecxr/9H2JWPy9ZAkgFpMSzVRiKn6kZRORd
dRjxCFwmCzgVud6EBBQRRKt+xu8Nnem53dgX1OwydpDixUjOyShh72Kmyoia4EKH
hCzNvDc8DaU2HuAhCE3ziwioWh4ZxbM94L4jLhWkaxxClDPaSVHxGN1YLRZ3Akg5
QugRPq4Np/UztJ2SDmRbcHxhem9ilZjBXFCm0rIDB/C8RJc5vAo70pRGsL359raJ
71vddCiQnK6oqgfmf7jc7g5dOFV/anbiSA99bwqWUfNPgLCpoNKp7pK3PZp6jKEF
9r2O2zeW4w2cJzfcvkVaUeR/x7xo2yZat5XTu18HATsZdlXSHATjl/tOFVhD8Irh
E2vGxQHOFwrOLm9ujliVuoX/dwgjHazOEa9UPikWBbsdLEpcFJKK0v1sK3JbzkaM
jO5XkfkANCzOBF05fC7L9ZLhth0+iDhjT05L36CgHg1Fy8LXtb08kcwoSXold4kA
dJMOQJIkaOvGzl+RZc38iXc7zBm81JA9IN2TdZq1KXYtT18anuSVNvi78UmGRE7c
kLYhlSYzRGY6buzM4UugC2bJL+j4BRWnOwhEY/vJJj2Q23XB2dk141A3KcT6F4Db
VY+zobZmTcqljIZFCCPino2UIpVKXX+8tQ3lEG0WAwvu2SdE39rbYaNl2rhGn4ug
170++ewmk0mu4rZP4C41lsnHvK5aAJAsmqbPUgbpe5FD2GY90QKkiZzAceNverA3
fBGncV5xE3QaNmpA7OZHC4MYdd2bmwCZNf2Og7LIGjG7kIlvEKISxRTnIbt4vQrf
geki2WlGi6klLoABuCDjHDcRVmZ6KaTlnjbVRLQcpO2ieBdidlG62mp0yginM0Sr
I3ans//RRLoLlTFUk3tlWOzPupR6Ylq3cTJSec7qk+DCqju0MGrEL48JOyoBfi5R
Hnzv2wHXVyz9GZwno8E1HPBst7LbxSqYN7myage3/qy2v+ThI4nidhvhKxHn+g2B
CcLABrRsVz0krFyr9n/lOksIDpysSGuNOeF9w+JLPTawA+LLs49fEZv1JVZoglIp
nPePvXhuSx+CPbBboZ4VayvnRH6Yht4ILDSYaTybkCaQ1vP6yiOuuyTPi3rmd5LO
kLR3eUKex+7Ig0iQZHsZbO+BoL2lsPAw2oOhCbTZvEe6N7lk6xNxXAyMcmDcoAMN
yF9magZaSpcIsEwkAbxytH4OP/DV1GwkSQyzuAtOMUlrqs+lCRltDqN8JyYO4b2d
paYutKfmMJRzK+t1Z9grE0pnyNE4OlNlj1wkxHIkCN/p4JkIt0uGSwR94p7KIyte
uQib+nHYxJPKGzSR9pBPf33gjVzw7pKcwL4N0xLiNUwn2/js8hUrPnwxqhQ3GzhU
5nOzFF7cQ/hVjjhEy8pRm9OhV3Ahuvfm5B9GrrsAqOebiphH/eJnmoHEnwxW+1mk
C2CCKrQnAWw66J2F+1ikcOw/EpaxbtFM+ZKHSXK8xvm5sjrcCG6Geeacl43I13Nz
FuzCQxrNVk+D7UsKI9nIuKCUX1X0VyEeXH/VZa5G+Yv1eE+0TqA04H501zLl8zr9
la5q2NPY5UC0kdpDIc1zJElvZwZ2HBIw74u+Bc1m9Hf/v+DksrvgJ3u8yvsc7IWu
wOk4/OyUY+0gOO1RHqVMPO27xlTmJrbNKgGUsMkMeX5XH2ehJ7wfA5kxkTUO1zi3
N35vKTTiXWWJwc45o+R171Pie/CYZHMJR5QZ2dFjyzk99iQjl4HWMV64c0nwEng7
NPZgyIVhJrZp4R3nHCFt6kiNTmRT33w1GA1M4hky0ITl9np2uwYo+jO83lJt8dTA
q03bztdH9J6o61ICuFXvngOBeT65ND9KSD5CJCz5OUqsJlb6PRksftJnW6cQuKSs
TY2tVxYFE7Ni0nvrV+1pBOUM97Mcp/8EnvKKNZopjCxjy98XqS6JMC2oAeuOqvkj
Al+1mL3VExbt8A5RPwIl6t3zguYk420ujsyzuWI56e5kMNDQi79FR/saol9GWrFk
9magEByF9ZVh+/lM9G3lI1e28V4Ft7vLXqocTEFdNCIX+QId9+Yctt80Azk9dxvf
vIyg1M+JmJpjCA5gWRpmdAtvZPtKI24cN5r4D8rbnQdEPr8xZ0RLATNiVe8c23y9
/rVzQDUg1Z8h41WTT8iwj1lNWOMa7S1m6XmCPqQhsfMHjRH0uPiJ6RJf4yPIYP5H
eoNbnguN8/5D4x2K7m0cJG0lakSHN20eGsF0fWhImXMaZ7taaEMCBhTTqny0OJy8
WHVDedjhbU/W4ZdMLr0ZnIYHDX1au7sgHOsL32t895zHfe/pnqlIZPlpMzF9GfLN
YlEA3tNXpHGx8YoRiACuJcc6/iSGDPLxb6eZoLyy6c+pLKftXw/tjlNHe6ed8ROF
/skNUAvt+ZV5vc3luSU3AHuD63KswBfZb/bY8LZLm+tzfKVY/mo4dnR8i6wQvTZU
0K65Kt7ovMlEeO0vnvcWqZI8cak1pjA6p+tM5+u7tdpZsKl92bI5g3v6xdpnDWw1
FonwfzR2r1o+bEQEQQbPUQS9Vkh1sttsbywwhXnzHDidc/7at43QlKGjXu7W4iZf
yUrlKk/7JLxvEor9JNfx4PZrbo9V7nZcRNpbMG5NALEaJOD4CtSJw/0l/G4THo3E
7T9Ayb1AaIBtOVi7ivHktWy64KCRSsVRf4emJW+QR8+SipSnsmKZhDjoG0gFY/4X
sw7ohar0nFEBQ4bLLTjUjCeLpaEJHSUWWZtH/Imb4D98rZzPzqL0QFI//WgkmyWq
zOqaBma3JSOdPpg0IM+AKA==
`protect END_PROTECTED
