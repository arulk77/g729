`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42l97wk2XYwDj43Zz/yWiL7bd2DwVnej6nOlap0kHfWU
1tQplsMUtnOc5s9clECfT6AutmGqba4f0L7YP/kwlj586o7vj8Hnc7cqsrYuUV5l
UJG6WcrvBm0fTTSZNWD9jdX+EKwgxTXnHmIV3r0bSW8y+DJD84aNt+jl28qrwK9t
XdypWjJAFaOpq0nWTdhNH1PjSkMLBjfnwxiblAyjw3XPKaa4PK3EEVv87Z+EhsaJ
QtU/9ZwzfZuNIAZ/JwfnFU5jG/JYNvAL/KXMMLDe5ZL7Imd44TzMFKOUcnakq2l1
xH+NfYnUoY+ObihDmXcJToRh3V4aMIQ8sx0EStBHeqsgQ6PyHBKDQiNlYd5u4Ii+
3lFBDqWljD3ZWHd5Nad/WNTem7GwDNxEx8tUEGy9XushEktR0d4hGft5CnMm6o42
0KIlMCtblUFJi0N2BmAjzaOadHtkQdcWBubAi3OafX0eqUm7ZnddtRn1b3381KUD
`protect END_PROTECTED
