`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
iqfUR79qpq0vtxjmrGoHJf7dgU13r30g3qebSD57RLcXIQI2TLk6AsAsDW5OCCCa
d57WiVcVv5t9xpOwuKZhkExbSRA6YV/kAODnBD6ZJtrAoc1lMQ6OqpPjRuImZ/l/
rdEGFa1iMRL7j07RU/b48m7dc4Yjb80rNRHej2jlE5LaljDyP0ziVuTMgjjhT9UU
jgAJBdEhYCH9fbOYinPCxkIsqcFYOtQYAyTX0mwxvWDi1BCmtUa7I3wXQKZKzEHb
UMsN2rarpdF+vSyWfWYiwe5VOQdYl8u7DRiQXN/iyic=
`protect END_PROTECTED
