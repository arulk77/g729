`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAY6iJtdXMo86CQLMtxAicQJ7RvXXhOnEy76onazDGpqX
lNbYPeg12PE1wrlW6u8CpmcR48Rj/p7tRQknKaRBr5bbcikBGDAMGS60ZXdqLAxY
dhTJhlXMLrCaMCKt2GoZQ1+OuPzc8YBM0/boMl8mOT50eG6J1MDhSFOgupWHxvCB
rgnhrZaHXNnSCEZEUtyhieOIw0/++feiRXvsYaDyM/j2OjVdieEUH3b3R+Xd3TQh
/xzLJGX3EZwGfeVLRnlCRkIvZCb0Vvq+3IKTtBihS+m2RJN3w0hshHhoiAPjIgbg
PrZPYQG8qXg7slthiWn5z5F89+5wDtuKvSNtERHnLRZVU8uYxSpqxy1J8tyi2O5h
9ukraMtShgRaGRp+GCx5PW0LpN+3plHSnYOrzIQ9xoUsFmRXYUsDAYK4tY3X9Gq9
j12jknq3Re4oZUFXZhrQR2ONA3H3phLGsqwvEV51nF+d3pMTAniPMfMUehDC055c
oz8eceaVMZcGfxWnCQ/CkAXOfwSEeZM1oTeS56VCqx0lTRzwxYnyGOLNs1bfn1ft
3/XpkMUi7V7wEh3ESldsMdrGOcsXsvQAIY/RWKCCPw6YG9OxmYT3BvztV6i/3+PP
QTiUjrJey2MIbaz3/DPvao7XQG7Uywfn/XXWrL6jKtMTTSh1UiNg6lV6lHFKNOfk
s+aoYq26e8JkQrJTGo83rQk89FoK6OQD+lo4GdJtLVZTHipDbz0W6LXrwdErSil4
z/kIxHBYakje8hA37Xa/emXzAB4JhI1prjrz5DBUcoMhFioyISiNtgDHqvAaO+2c
GznJpLV6z3PRfyhQOVc8jBk/GZ0c7JYlw/8D5/9EuiKvquVrNsraXuVIyq5yHhKO
tQyKMm/LnvTNSB3s01E0AlPwzW3HUFYWDb3RqZCki7Ydl1CVqEkAWOdxyTrQPRJZ
eElWW+pPx9+10wK8w9U7gRK4+tni1kUl6HwGNd7j2bfkYlzensAC+PnPIBQ8+15j
QioOJaWRiRWM6s3iZDnvYOzyE5SUK858VsBrGlLPI+TJFhMx0W5GsRu3y/rnQqKT
TdY0eMGpRYq81oRrh+scbgFmt8LhQ8/HXN5zf7IAk3LYGRYCbTDIC4WEjS9Z+yoH
gxFQFnaDdYASOtNOjDRihgsHX81GjH4np/rEv/QiM7DAelDKJoFFPtAZQm8VxTq4
FkrV3Q5c5XMZBs3ckTbTnCJBo7RRzB1k+9h817/Qc16Jw/9ijLHlBOIsnqdvz4Ch
pYYpk9chNUia+/w/HH/aF9MOc1TLM/CS2PCGPt1y1sXF1Iiu2iOCwgczpNjwmlxS
dOGHSJFsGNyZPXSNW4ZcqEYmOJLXKRZISSJlt4t0LeIdSaFsvZJljhwxb67oxSsQ
XMbVSEQStYl7W65J5UqcTVDOW7a6YGvzQBEh8L/aqRg/uBxPtk8UyoRxZFQGgAA/
yH5R8oT7cM35UDBiLU+AhVpFCG/9JM/K1jA5f8k+1+8YcQzIPbpP0DJX+woJTqMQ
5S+QKEwI4F43FDwmUBwiuxScw3ljXC3pn7qFdhYG63qkscft7IucZ9BNu5+tMvK7
8T3jXL43DQx14BKj011jsftj9O9VCTLQdfrTo9xNzyi8sa+N1y376kQmRsOkiKNQ
3oIx0puOKAQABrt0vD8Ynqiu/F6qyImaYk9V6GDEWPnKHo1uLZj/Boph5OksWrHw
shnx7UiomeyXbfTFtSoQkd+CoVbLh/HxWgUdO7Yka2ZnugGGxcA10KEc5yY5hhtB
oQFDThjP2Aa5rg0AUSeh6LzM0TL4iapZshY95NLUFp3vXOMNlbNYhm03f7owkHEo
7gAtWY/FvREX0apE58QNnUVuP28EDVyz4GxwB60hAamIOfOHpH170k+/tWz/RpYr
Qd74t1cbcyC2/UVkgvl13WNFew++CNTrSMzJKr3GhiTmpEDr9/t7ABqBFaI5RzGn
XB2R6UkgxAF/a5VktsFBrXaT2puSnhpgYS4XTC+7pZB6lfhUePVJiTPqd+OKNSXO
CUXwmpFotKJgp+/M1bKwQM07hyjN9Rx6X6Yf0MgR91zXPJlDYrr5ZV6pYBUP/Kh7
AVshRdy/9FQSIcsbKdpb7DnUhst52Bq4xRujWUyTg7rmUXOeFgi2abs2jmi59vNe
3BlVE2CuvBamFDgwPAZiuo7myXM9d+FpRqKQ2aIK/C+3bkBUSN0uUvrpo4co+nkM
AUZVfgXpaeuuK7KEa6ICrCy/Urk1/4tEnfDM0vuvZCmEw70+7R4NFMgBRfMVgcwY
vcnLcpDfTv0IeTqEc9UKPyOqj4q6cn6AwXAZyCbh5Vgrp7bV1JK8rjYpD5NPxHsj
U2f0/nQT1jCAVfFj0cG3WJ7dSuiXDBsMc4wqXi81EYH1NrRbw4rGK837UUt2ZiPv
WU2dMJ0y9akkLkLGIRwdMwNdv18eb7cRVfiqcU6o7U0A04ma/dpFMP7UabvHb26i
1/AFj8HdqZGxuZnTvrBNkwtXbzBX74qm/dewzNbzD/+7asBiYgWL8+ybtWDqonhI
4PK0qZ59KBlL7Kc193VbAlNq33Bh6dmHTZf9hqp3wOCaTzQGnu4kxqPD8Rz9Hm54
37nPyR1Koia0SYNyWkSSeGtoMcAlnq+rjt7dUt1QrpOM9dTSDriMZNZ5UaObX3re
UUz6bWHPz5P8YNpjACms71N2wZ9hMBdv9aDEH04pAUdfC3AxYHLle+DnlBwpeNNj
oN8rOYiZtPmCcLcRkmnB0axvO5RmLsXXmSUWVU3nJFAtAfkyP+cChnmt9B904bRJ
wFRj02N/QiSufPg7XoQ1WCD5ecGKe9zZjUPAN+iOJMiApXlqp0GkUbj7WV9iz+bg
Quv/+Ya5Xq1w6Dk8ccRof/yugBAgMnTG3VjkzWDw0W+qg+YQebg/o1AAsZ41uhu4
aQVlpJpgRx2eyCc4/J1LNl5M5ryCwhfnBVj4HaP7qZf4Vpj1+lGwbYbJpp+8ITCx
UYfmXnyMid1QoS4poNotG8C9yeQtbbD8VX9QNKvemxO4gJIYY9RM+ONc4+0IB6z9
IaEwOaxMQD7VMEarrieh6ltuEHxhj0YqDMK+3p3bHsRnkA0l9B//A1KX12pIpM6S
roQ2Rqdp8dY0jP6SVko95wiTpcyE165dt+MbNnAsMo+jFQ4lGoRqkGyA+JYoefNv
lXPmydMR17BqUONwjSUqyDYRmyO4/WYtuonik5lYocKAw9KxclSfOM0x9bkJ7YNk
80shCeQi/BAb6wzmr+xypjE38BdBGPnnAzl+ycuLhBitmD1LO1/hMHcREkL+GQTu
rLfDEMm1igp79vqKxgxJoHJCZ7K8pngBRZpcRva+q0u3CJEho0SA9pkCRbZH2412
bii0IwHbOWrqGtkr3FxbUwDbkMT5vpVznPZIVUhRYAKBKs+va6C8OaH8R2rfWbo8
lSa0TFRikM1JglVEhoHwXBRY0SDxMBIIBzj+TAUwNYCAz1b4dKpCYdjH1BBiTAPH
IjhMCQF3OPnTeb0uolFjqmvh16G6KmRwAmAuF4cWXgtACZidVsVssNC9++QhaIYU
HLtLTl8fVgdY6ip97FwjsmDX48fGnsl0+FrHW8gkMbKOxD0EhX6BqgAZFS3vy748
8KgvspRXlZs4x6z41FlZKfkSSLxQhZETw1jv4M0DYarEDLPGOnSieeCHJR8xz8k3
SiWPAvqOtkpo35sEA7PEsu6YSr2sn5drlg/x3StEC9zN0tn0YFZNDc1Za+Ek40+8
ubsQCdn8mQmBsX9CtxKr987MoTvJgt8I/2aNmeOVyO6gvNhDJP75yv2A1klh6l30
c4otmdVYwvsXfnPs9Mg+Rw0OPGBIllRMLzx/4qmm/WYm5qo7IuOH67EV5vIT2e3i
UQA5lKMMLyLB0Z7uUL8maYR5nLUWKDznu1arnnlnI24oL9VPYCzL4rYTQYCL8qmi
wEPdf3iLpiAzU+0dmIhMNotTO0IX036BtipTOxejjtZzFT5VZBx72Gp/pcVp7iGk
8DGHcsBi8OQIAvvRC5FvrZ70ZSQgjw8wqQt0/4epZ9Ib61Km+4Jsr2DucA6WDuIy
GJP2juCCkSTI+4ldDoQlzXkZjOGT+Bi4RDj3pSYnj2DfZevDhPAiGffQHBolt8KC
zi8LW+b0bZlfqHR5qUmvwUGXHIce0XlBY3g725390XvndHC3vzMc3yCN1/J6cr8H
xrIQsRAX2rUJukuNzGgq73MyJeN58NhJg/ZIBAlCygu331Ux6CX6U8VpT5TAwW8E
L3PdZKxzLCv1LxTCHOtWuXI397673I3WGJ3iNVrykD6GlBovDdsskZ1DsL9Z2wbC
JV/sQPzlQjD4uM5Rqdv8EiK5q22qjbN+1z2oiUIyJn2TgEJcjSeRg9oYFsVkdA4k
hs9m5ZqNsRj37QlhrzZAHV0vVsb2WSIEIRP4arCKEJJUTiSGRdJRSHK/j5M+JCYF
x5vvMzuQ+8vrooMIPoaKhXtujzNF0GYhQRGv3HnjwOqDyo8pBzHpr4iwtyFiwHIT
kuGXRupbiXAvLVJ51lEbvDQSyUi4AG1E7LTioauNWGbhyHHVEe7D3KYu0APiIogr
lPlXYsDk0Ux9KnxQKij7hvmeqnCAAlHJuFl6UtKWPHFiZXKQUyfSe+oa4c9VTa8Q
aoEevDmDkNacgT+sihubQWOTNxACDtgNZpGYXEyJYGQ0n3z/jT/ZDrxS45p+zBs5
uPJ3/KM3XgtCr42D9USltvFuaoQluHbpUO6Ezy6qHljPmjidYu26U6LYy5X80dtx
mzspHBE1ZlnjskDBMWDQLXpt8+ooqZQmWztWM1Ilhzfot9Y8Rl8IpBebAIf8Ce4k
E8reQreR72qC3EXicleJhbwC+CiAHl1XRYhUI1jHffL0fhQ1j5WyZlKs7cHysYSF
cAOiJzediwbOpzPIe+NkJ04rAH+wJM1GQM38Jfh9WFXWIuUPUFg4EZ2BBF8rJPUP
Vpyr/Zs+eMus6PHBTXsQlEC7nEOlsKuY4CCeHcw/EnOFJSAKrpUtgkzJghBU8c2i
RUaCsz8KZfBe5+rCgF17aDbfPkJOajpP248J2hjE8t02I196AjzzEHq05w3Hpk7I
QQMwxFN4y0J6OuMka2lpjZ5G7vEXoyI18sTf/s/0C/SGKI1hH53qibl1jerC3qIw
/WUF37MuBizrU722s1MEqWMZhwDYAc8/vFLVrK15BRmecVwwVkwkNzNjlFJrRrCH
jkGL0NHFieTSd3ujDEtKFvzulBq9qmnwu0X1EHMihcBNInv7NtB79EiOn3TX0dYm
BxmdFi+vsgBKAoLZ/EhWwXyQ+Q7WXUkZ64yL0+dXQXZQItWy5p6gihKR/pqVFF+0
gN8gBHLuOjmm8nx0927g4LuhPXa7k41DW+9D+BPsNUvTUA0KOLSQENsAteJQUbR1
bq0xMLjt586dlKqgjmXz7CJRL1tYy68GB3gGRC2HdLl4S8Y9Dy+xGk5myR/4OXmO
7rm31CiY0rKKgGtNpAy+5udKYlBzdiqk+iTcJJ1+nCsk4Dr+frQspW5UL1kA5gJj
UVW0nFz2X8OZIwTt1Ww7IEPV8VfdXgSlOPNK6ndZELH+Bgdjo4rJa3bME8itfyeZ
51Rl+UgEFkh8JjxIwCAFp+saAndUFfSc+qwb+lfly8NF7YEJ5g2cseCDHDL9TShB
vG2EpfdqGOLmPKox7ZbEZ/9jdEnOOJZYcIEtSdQRXMMAZ7xybb9sIip4YWhbTQwD
zNENf24qcglNcXZlmw4jDQl/XwON6Up/bnbfampPght8ZIjFXqrwdpIJbspbBlmH
FSFlP+miVb1nskmgvUkGiQ6F8L/BqxWr//0n1ShnEjSaZWydiPMeWaHoBHwYppRy
oX9BTcKERSOgP+FhyTLw1ld2fty+j9k4t/04Ieu6HkOHUctavj9Wa8W5PZXsa+G0
1MOHIYWHa8mVHa1PzVBhz0BNBTTtI6iurhR+L3RxhXjzKdkmmwGYxudDZz04qDK4
CvTZpLrKOkyzfmr0GCiAR/HGdkiMtyzXEIzbW5ViDn6zWWNxffIauKAQ75/zw+FS
luXWGOVwyfUT0livvUMwi6IaFaJM2VnWQx9fHqNqbY42D9NiWEcs1zrFx5WKf+Te
Gz8eTUfyCAe3p4sXmq7M5vaDYKKe8iQMRoELLAY4crUIU0XyHMoi4u5Amt9IuyzD
dyFRFyfn1rpeETZ4Wq08IrGddrjmMCX1q9U2RjasmO/LvCCRLni/IAiPqpz1fggY
Pr0IV4TOBXmPqVZJzT2WLfgnSoquLfZfGodSeYo2KHRlSkQ04MCLXsc/EMZg42d1
IwGFlUUfzam/1YSFE316Ib+ivqg+Pmpedtipt52rI7XO81ZNcXSfM1QrUN/izkQO
f9MgTJ3BwpAWWVB/iWKuYNIS6Ygu7RnIyUkj3SK6CYVbOAInqOkfPH6PU/sBQ4p8
+YPR3zVILQKkile7sJ1PspvSfoFLI3nBOjYSAieU28XzqtpyXeif+dJT6UEcW7lh
YEwSJE8EINfjnmRhtWmQBVGWbVPCVGT05YNEGO5Qmvh8hXc/E8f7xJkGdY2rcEkn
UcNMWTOuEMBFUAMAqMJPeCzcw8AZn4j3NCkzqor4F91pH9XbqPrzn0SycODgwhns
V5tu5QGhXzC3vekwmoYTXUhnG8sJnnBA1YyQoCr/xRvKovWNx49qDfa29pAp25VK
uWQI8mY4XjW03/vs5oK4jT+971H1IjhqK2g5wpdEO/zNcC7VeER/8/peDDeDWAD7
2AamnBGKgmhaLm4ayKpwpm5c9c6V+DxiXP1ZK9oFXhO1AUIaTBIrtMJIGE2ZFxZD
jXtMgWRi5e1eMV9Ma7RPs8z5ttzZesoWYSlXF4HwrISU3Z538nlWqXqgEiVsxFVT
7TX1HE16yFOrzXdvIHYpRlbT1BvucxqhHxuEhNjpWaG1DJqgCFL9YSUbQpGCyPnf
upyOnmyBrnqo4JNdo755naznHtQ0O/qMckwj6ov3POPH+eqiLx21tiVs2MCi+xEm
eHnhof4kRyG4xPdUvVNLQfwOyd8s9iXvxvW+QYSDWUsYKHbp1Kz2Dq1UK3XCXnsq
4Iqat01RrJAA5ZKAf1eEqJitO9+0+YY96cOU4G86AOQvSS6Dz1za8Km1cVdTiIvI
10boXRWNeGxVNPl+M/6RlDEv4DG3JhodDKyvu6zdY1hYLw7j7q4a7d90aKi21Y+J
oH5E/WU1JPgSm6P7icBtNByGHrHfJl49Ib+ojAZzndl2Cb4SdVMbkynw8G/3W7BJ
0tpC7Xz3znTPw6fqqJsGyZrNX6J9rMSmgjnR8jLTSXlkys0SYNBzcNRB8S7R6Rkp
Np995mquL0lFCTn1RwDObfP3Xrn5tT8QSq1xXn2jVRCzf+jJd9etY4qBmzHJChM7
hXdAZ7U5XKKNH2nD7bqfN76PRS9sBTyudbzBQowBLSZkGikeESNb8POpJIzjt10I
mXz/BX0DroOtfi1QyUyIdVGkQypw0Xt1olR4wWgyg7R2arAQPaC+UNA1Anr1MkLz
NDjEDeKX9OdD4lYnojx9QNNS0WjyVxEnLxxZzEe2G3KrEQAkxY7qZYPE9lqckdaA
m5ytN5dBHOeqxAeJT4eWY07T7ZLkz4XcMJQ0HRseAyylDAphhsvx4DSlQmSJKXji
jas4YLPdMBNmErNNPhwMmxrKXzb+b5SYHx8KuEfnTEzroGVuqZwDkgo2E2Bj5nIQ
Mva1uGwWMICq5cXZ/iWFl5mLEYhCX7Ald+HSLKyF2Dq30R9s4iPn+Jz5aZgC/oe5
PBb9Jl5gS32yyQkE6uvo7fmrpo1HuOaIgrR9Hwq4Vz+C42MibosghLPuxsoIHp53
2/q+ju/mDLP44IBlxLUE66pOL68+OteFfrY7DiB4mV44Y74v4z6CwBfT5VWehBs5
ZkNpoJYIGXJ7g/ON5ZnkCgjBRy4aywIjWsYhe4/Dm8wlvtbnnLof65nQWM3olzwY
Rk0/73bxJ0tfbjPneEE0gmyEWBDnNLBBcfixtvD1q02JJ4OjSOxqkZKv2E0bxtRV
4hU9XNjQE/U1dEC4TA1wWbs+zzqGcIHF4YAnhqiShI5F635rHj9T3IoiYPO1BWYb
SWDtBqWozsLnyIc20uKY5edmnKnbaGvE3W4L3l/8H8cI5foU+616H++Jv3xkJ5ZU
HdPfBbgyHc2sh/hAU5p2g5HAfot8FPhxJbbZZghVc7LjcA2k0tcWEM0ORbHAJZXp
nGugydhXJrRUP6KeXzK3ODMy0yp3dqzBOXC2n0G5VHXf8/NCdXX/jAwRVFn0Srpt
IwX+zNm5F4X6kx8yCUzp71W11z9LwczpFavHqvkrhFfQdg92mVSV7sfrh5Fd6JDj
tvdML5UaQsQQGUsOegc7wWlONkuD432YmVR8cJQqXQtMALvwoGoMAFJrpBcgMaiC
NurdtP6p07lw0XDqyQdOWC86Ygn2VNoncj1t1beDHurlyzzaz/OlAv46ijDjS7+c
ApgyQyic3MdJmHLqm+tGHp93BS4z+qnRqLufU7au0GcUrZ0CjV9W9MZTgwb8+SLd
Q/5u20PRjAMq/6y95gwNIXOjvyNdKZ9JBFiTvJ7aDgRh8WLsvRTMzwEElbobpHmZ
kF9lP/MbHwQ0uXvG4KmpHyMfFIuziNOHpbulMh96woGHi8oIrWP4Pa13qfekIGDL
dMGeLJT+xO2nP0H9pxwCWBgcp1sfmbnf9yeKj6qRTZ/jfLRZB5Am2gh2h6vVwOQg
kNg8HkS2YtJH2NE8VZRaXmwKUiU9Ax3vJoyjIENlLZPiMcCkaRD+CXAv5bIez0fN
OQfe4yL1XdSquKRVsgavwvvA4y0Vasmi4tyM0tJg7XHf0Z4KU4XTIEPCtTPH/UAV
IIfUHH3G4xncjIT92eD/s7ITeP2mezlbS7hwbOFDUMg6cdl1M0b5aXJzTmkXidil
xeX0kwH8ntm+1qnR1zFsR40MjivbAlmgp5s9vhK26TUzHws2o7DX+LP71BwvOowr
51YVuA0AWgwiqRtrncyhQZAQIqZIXciuHmca2s9H4TY+aHr8vDRSu041qjnlLtCq
uJVtG/XUVw1UgIsCX3j0yAHIM96pDaqjaRQgEx+cHVtFjkMpXdUScdo+nWHzgh3l
k4a1fk9W4NTDrbdPcttIFxqt5W/U339fxfcX/AZ67KHLwml3MSTl3GW+FKOD76E2
e2gWOrOZid5lmvDejDxDcvDBbjUPhzUOa9xaaDSUapswq+1dhE9vJ1H44UOrIKe3
GF58TnLj9KkdAL8T0JFU/mC18ynoc28egEabyJBqxvgRtJS2pkavHLdzn7soUn0N
OIFpliggSXECnkbWr3+UYE7UYwovlwr07vCdZ72/Lutd1vkenRZil1ZUsWrUjYWE
d8X/d5beicGglR7qh1GYH8as7QanEGpo94LKPpNpFcpeOHPXoQuFUDj3/HbTUAgn
PwWqdnKNqG4E0Vay2LMtz9wn08EcvubaWCl+xyiNM0KbJsDOgPExHtxI3yEZZLcc
kaMKWbJ2GnlgUCGohHhHmxmQbDh8KCNd0Fylxd3ff0flC33nlKJNRXAUqG+8aa0v
eKwgHnX6Ook5o+RfBsxs4L+Z50t6s5kOYp0NGxUYSrEt/UCklbLZgOTuDQodhU+j
8+6AYc6pARf8JAgdQtAV2g8cP7dgv6LM5PUrvfAS+xZ59aZMr/GgS3QmxdF01keZ
bhfMPucfGN4BnffHUYOIAcJ3etqE8VU4hfDhFTpt9rQ+l4SWfm9fpag79GhmLPgI
hxgL6llcF85IX444S3BvG4qbWPLU7SJL3Q7xTgOrUefD/w3PvFaywx/oxj9ESken
CDmG/qSBiXZVxC5RMvApjf/gRaECYc01FovYFc2BjwWOmVtLsYAcQRh8dBcVkJSM
aPoYihkys5kjT/i78Szh/rOGP1u59dKWLIdp4URk3IFN0bvn8vK+vxkjNZ7apNsp
C/39r+v1AlU2itZ0vsvLeI2du86usA5bO8ipdSMv942IJQJFqf/PDs42XDHiUlOI
3sQtN2NTFz6yKrVXucLpzpkNP9fs+jU4AB4As1KdekQwgNbX/W3F1X5AfYTd2pWA
TClZy2m8vICY6+KNR8t8Fmbu7/qCUnl8g/sh1i3Jx37qIOqAXFDaNPQ6pBpu11pX
d8UQFDfuMYNhYuAizogIM03yfh6jehPGt64ciUMCYX6C3uKm+MqqLptrF0f7ROFc
KBgwubPVGlOwDEjAxfGxNalsqCPV+Qh2gEkJasLRi2yy+XaZBUE3sLIDPu08ooTw
lrpDjpix4kDabAPSYBXM6+7lDT1GE7L/pn7ThxuU6QycMmUak17mM1V/fXMgCsgZ
SaNpoyrm457R2pKZ4FI51jmHuPtV/U0DPDbI+UneJG5dveuedSTXfNlO6y4A2RIC
PMMK3wx9kJQiuFmMCN6KqFUPh2P5/iD7TXvHnaJge2PYs7WCVfapv82JVkAp07RI
Vvl2wsmJh3LDUMS6RiCeiNKbKG8cM1qwAk9cCiMXGB0HKW+oTQu7bOEKEY4vciCX
E2iCtBl+uFsv2c05G2QFPqvTFOyr9HARhv512+Imx497rAEpnpuxVJTRYjX/vQFE
rfGJtAFGalEUDAikmxkCCSH3fKzofBC3ra3vUz3/KjV1rj0rtqoc/mhVYfKaH3/0
nti3d32WMQvZLG4cbOTadpR9GAvUYS0VjPRgIOO5Z3e8Vk4L4JiTcANQEZb072z3
Lo5NCVyfqmwTK8J1oeWtYhURmxZKpshiO/UNas/83+8QHZzzIdSnsYW/YPOiT7wl
NstNkCmsOjC5+StoKxLFUB8VtYGMrN5zngLiH/PDYAlXVQLPQtagRxpqChIzRkr4
17zdglz1h+ku0JMVp6rL6wQ6fuiZnZijfXmd5HZ3Ipk5WU2M756k1y43H245VLQg
rEEd8wFR59pD+g1NuVZ95iV7YkZmWhDuqmff9vnT81VOffUfnLHtkZJYwXFncHJV
XR9FPNX8D9i9Qefew/qfdNwv5DYqj58iS0/eDPQmPuarhVibYPE2dtYdBbZ/qHlx
N+yCCJss4loAJJilXanunOKyKRfcahfSsVtWXrXJ/HM+6WJWRQR0pyCV7KxIJ9Az
/RKyM1EysFZ4RobnK8eKVAneA8wzdELKSZQZPiFXGoXS/n88Wf26clOR1Z51aKXA
Mr6BpVwWyiMsA7VPBwbdvgo2GhsoBuGe5HRH6zx5HTh4FItmyx6DTvHMBLKl3nw6
Ln5EnD2oFmdauk3Y7RfjiYr6jmwAScNtDXmZlm2NO6cFD0OUaUDxueq5Bsr9Tw2P
xeWWFCKLa32CTiYB0ytY8o+rX26LnzH5E00TSkt8YuV5Rw7KT8VcmQrGlntnsHj0
ao8fabEYp9gdHY3tbKDfNo2+8bQWOTm/2G5mvd8gAKxau53OhD3UdtDwLs+Fsu5R
90ef0l4O9aTkjPD6yjqzAT7hSGnFCKTCvRWD9UzzRT60KOTRbLH8SgAftMrn1IPZ
nK16+begZyfvCgVq3sJ3gZT9cUo6Ctmd36pZuXeM1Lm1ck/+rlID+1sNHcQsxAOf
K15bD1G61bni7wwYmoXk/oMokf+hZuLsUs2fjWUltSltbX1sw6BS+CPUE7UEwiZ1
1a6sostn1/OMH4G9CWEOQhaSQopZssYGUaO/1+IZ9B9gqaibG5cKX6tOnOp1RPLe
m/egp6/Pmdii/olGlu+vICs8dHDUYkAfh351/4Gzr/MV2/N1vR/V/IYBs6czUbUa
TFEUsm+pvgM5YrAmTz+mc6Eyq0qjNDxfGW2uCbyiWgRKNJ1a+BiFUjcA9lEjoi4f
NKbwxix/vn9NB30Gv5YqXzUfCbIeQRqsZyutu8WVwv0z8yjGLsp1k5f6S64lJbLn
0g9pMZRhRcXFOhEOTzGzThXyePSP2s+5+qSyQ32KxBqCxKQv6Lwen3Hy95l9WRzC
V5oFmGXstCEni607xo+IlROOZ7dGD/yZAuMuA6SDBIxoR8RNBePXpsQhHurnysMB
ewTK60Sw5Xp9EDXWQsGuMsajarjZx9WQ1SeDiEex8ntOfex3mSzh1h9dv4+GWSD1
SeUu0vge3CjlWF0gkxGIrWRgSAdoC25iSbx0bWSWfvrFMTWucIWXIaYUsUN5unSp
lV+pNkyMjIUuhzFa5jk8NGYgHh3RaGvTFXRZxYD6VdXdRTUJuopDWDNv7mliDR1x
vDCXaajwLX6bDQI/JNHqJAP0vuVa92HHFUypTudLg8CGQCJ3DF31WzIua8M2y1Qb
Uf4rEpteFOLx6LRuvBPwUEB5BrtfyH78MRxbrT9SObzrtF+Y5trUOBJMhMxBRRzh
LJVXSuwt8MNXb1U7HFrCIcugwUYs4jGfLkNDO9QVO/nT30a3KvelSeEfTEuCtZq3
Mu0Tq9cvgJIwysnt4uWssMVl0xEJAjEWzldaRzdQn7cDhBsCFlIG8AQS/zMouYcb
6M+wsIPyez/SLMcG4yU8xA0B0B8/FUNcrX9byk1mEWhXPtfZhmMx0e6DhtxuvlOj
VHQlnHuN/nS+6b67acilv97BPZPeQrU9hRxF9Znz45M5QWQNBQ9q4mLyU1BJ7uMg
/XAr4tH7qwmZJ1MxpirzWyCbu2Sa1R+Sv7aWf6IyaNnCLPDzZyU2f71BikZ9F+yH
eLx7tl6tCEeBqsUrV7thtqsDM/uWa1cEXPk6qrRj+78L/IUffDzkilwrR+IqKan7
CU3XVa5Miw/JwOu41ePugC3uKxWcXW0wp58g/g8Fxt3cTjVcKvtXHLaKQovQvjhE
WZDo0tkrqWCiuqv9MBkUVXkwJulEKxuQtnOgxcZb29fgC2QPfoBLRoQqN/k3s21A
fV3tXO7Z1VvH+lDUTXtFXRJgK+oeSK2oXER1FdNEBTRhQMtBepD9IumWC19ReFd8
Suzef1MJNpdcvExr1kUR16QUpdxR+jPa3SqBDRvpViMjYozWdtuhEdaUpXGNN/bn
M7iw7/G406s6HjI75zL/Ic4ZBr1kjxI2X2vqsCkHxVh+QCYJ8QRLUwsyEAo3SOKl
HIdP3K67rQnusDx9nBtI74yGiXxALTG1DTyrlyoO8N7g1+2jBe0RcOHn1gdW4yU1
QuNOZ0DRE6yv1lsUFj0RnDCNK9QnJ4isoba1R+bWLPvUaB3VPm5OAV5kEvmDmcUj
B49g157mvEXyuvAadsIXT9DpcSZK1qpjVeK75r7PUqUS6gdT0vYDZskk0urBKc2z
l8bwnu/7t4aZvkSdQmBftotaMt29Tk80aNfWtBcOxvl6yVUEzfWhgoTjeYZ4puk4
hv6zoWyNiA5/1X7zHphSZvwgA/8ZNmTgU3HEIAi7BEXVEQ/WnzCFO/+4QLPVycl9
31OInZZm/11J8cb0VUs5NffmV9PecTDEO0nvVydFQ2bjIEAWlVn8Mtv+KPxd8px4
mo8Mv7MHBgjAqhI0ZXotb9gv6AurR/+1na3QkO9X2Zbo2ppSofESviQuJy8+D22M
sn6aSqiYDec4hteNExT0aAHPjC8kymd6OWquqZEiEJDCa2ivgmwAZpVHt9C/pS/A
TSZFpEfLkUU6A7VhLg+F4vdOcxWUkUhj/kYjoAPwTGWK08kpyoVVS56wSKyVNp5G
sHoXfAL3HaOeU8khSpJe8rFOkLIr7S8qEtI893Nf3WJupkcHhHTLR1WcGXot7bnb
cTeuEIe8NuWmPBw05eNRbxk+eMLW4N7G36PJifH0l6vESoD1hSPZfBHaxBGQzlIA
gElQsBYX5zzZwglbQ/XfnWjpFt3u8bUlp191PA/3Ue77XgdQC5jlqZlrZHtPoWxI
PtM+dZ1kawoWqNyOf3R4BGEvKZH5YrVc2yrlGj6al9ywtqm3Vkk3pBSXWPKX1+mG
wEcbkK86j8jFMcHo3aDX6OtY1E9b/ohZ2LWNL1E+wcP7e4U29+w2dh/9AUSnZYif
l0R11GKuzWSofOmK5URGnRufZ7pH4KFILh6PfvueoAf3QakQPYRmO9mkbaVv+fTj
bZWwxfFcpZh4CnRR+ihdvVpwaiixlErZXxY68A9MrtquissFidAE0wIt/AkTw0JY
yFZGAE15u/KpVhTGLwi3PhvSFWc75GAwtmCRhkeY1apqgTNal6G+fvjJeZyFAra8
jAdUnvnUFp2mit8ljd2iasPiJovFB0LdHc9lNDbOs1jIGn9K5tWwJsayQ62wgMgI
qvPYoG2DSYo48jqeQaUQP0/I6NIrGUJDqzuV62U7Fl80cvF8KfgtNfRIBp7pbOGP
1fBZv/+1Sy900JP9xKdfsYKfoUSs7Pcw7bWxxb+dWHF9hsyKeQgtCeuRLwV14rdq
jnNfWsJjmnBEF5jDXJaj8zKsUzWdpRzoY5LIQLRTHZIdjzdH5cFJfg7AQur75QfR
lU169Ch3PNskx/FOzWU9ozwja18OCgdHkYEFNy+p0uIeCZcXthClQoQuiOVLOiwd
BDHlvAgZ/dYQprEy2XM/BLZb4imYRn/KvX4hOOyZkWUg97OYvl4kxHFGyqhd/J3C
xLH63UZVxsUih5sIx++3ejtSVnrf5si9FiNX/qU7tYguqdODeg5HdYJVhPAUee/1
pJRrB/ZfirwId/+Ayvnnh+r1ZWZLgrCAt8kQ9EWzFzCpgXF6I2aOvJYeNqWyIUbB
PhoIdlekeAWH+0VusXyaGt58xw3mCk6ebu7HFs21hBGvTSPgTek+4WiHQvg2DpZM
gInRlhE+hUiPPakpIol2EGtzpYhItCgIOuPNOpKxj9LwlhNJB+wwWN46Ajik38Y2
fWkdG2VqURKJFdIloAh+YioH5md7fReMemrYpYBU8QMoyKUPBn7gaWW/ooMvNpgF
8CUfk8ir5vZTAS5dAjuDbKIma1dJtl9NN+luRpLx3nPHFlL4FmE1WsZC/BG1Qbhc
0hG/LlBQeA3GgCylfLe2Gdg+0uSED1kzwkhRXe6S5klHC4IH3nm4oHpNPPxRv+sF
qZe/auWa0tn3uz0rYKaI8KilXCF/YRimaQzLgpXZA/01E0PHS35oGyCVl7vnSkom
6APbDg1aVxEAkRysnga+pxoP5G/KOPV+SmA3EoDU4XLrgmIqZo7B1OK8DlBfzVZY
gPxi0uZPjooLjtjarMhGu++z6elhMvrxWgPVzKQID81thrcOL0ohzQRF6IfAaUkM
BdsvFi6USuj2zmvVydHeaWQJHv0Pc8kg4SHcqyd0lhKjxwdKCIJ1sZoZSo8gQDx5
DaUgF49xJhNZEcOuW1vXPdGnxeWNsiVUJwXblgobayV0le1OQ/pqXMZkD2Mo6od7
w1iHjIZ0q1N/wuhREfYIsOLfvKkEyPbKM1dzArtSe3SJNLuyTVs81uVJa2UldiG+
afe2pzh+g3y6apLpT0IJatgzHw3sZv1JTGAQ/fFP4CIfLA1ayzg/9OvYiY9yHN6L
Pxzr0ExDDcXvmCI7F99PRt2fkb/F73UBwFhguRs1CN6UP8BDCJCW2iNitb6Acnms
yA3vl5oZ630bEqrFf97DAlZG+WYkwkDi2f5y3zg/pmDRgpizE3UYBU2FJYzG+IX5
WTGLOcC1DEPZaFBuCPFhh34r62E58djMpRfHM0C7Nak6OQH6iSCM5iVf4+HA4nab
2pY4/3jgFjMHRWN8d2Ihp+CQ7c5/cTDKL7rFHdmrgQlmII/xAYHFgZp0VKnMJ/L3
l7yQ1irHUVjSpTXWfJeYkXaKhWYn8AcYZrHfCkmdNaWx/Aym42ULz7tsghzJlY1V
0VaJ/VFY0v9zFoBscVC6c3P6MPLUisTEsoc4MiAg9lx384cugckFzPYbNeBonLkT
RBX2vzuu0dnoLd3aZaLGvrwDlPV20QzEYcF2sROYD/l2rQssqd1m78dMLA1BwfWR
+AfPabMsYEssX2tMsb2/16Eq5KsB1jhW8uIe9kDmTAN7h+vfqOLpGUoYMGVoHEPA
RZpkJKTIr5XwKdYYbk5Mvl9CKxgMoUuEELvObs+vEiQR3Mcz/UKz6lzPGuC8zm9N
bujs5t5Vn3DhANn8AzHa2ctW1iqde1ZgP4edFBlc/T4sswy2UjpbJfpWOMUplGYd
BvB+ccLJnxxwePQwv9GOFOvCJzlyVybGtyD9p24YvpgcSG38/KnFZXiEfSXx1RW4
okWR9KnlMWLixCSFVFFXSAkkzYZE1ljT6Urshp8IS2exvN3rAWchlYjbVjESPmZG
TqjpqdnrsamIQPh1kQLPpykSZfxYfKDTLiGUyToWQ0uWZ3mbqit7h1iNlhZotxzf
toPxhKlPu+3c6Nik7ZXb3fp9lA1/KeKDJMPMeqFx/yCgv+4RlwWTxez2WUAV4WTH
Thrkr8fSM9wnWrUUVRfMT3exgT/YgCzOeaiM6akgpERVsvoAE1OpdwafCdwGGhfU
cr6mPfFj7SDupg7yX5/eQgVzOEXhXqNtNuXs+JkPHtfmYNAJAWUbcWoeVBP0jzge
MceBLxSHjuQz+fCi3Zfh3WZZkeJERWaSAuKn0inlqraex3uOGlGRiUY6B7s9MGb1
+Kls3GVswOHZN92kz9OnGTVXDqlezPX9YyROPKK7iAehVKlYPaqMMUWBMZBlrPpU
2G5KFB4B12TKr8QDuonfJ36yrERMaLzAL8Py9WvWo+bR4JY/PLOThDMjW6hllUgg
Msgsz9Cwzjj2WH3TM3bN+XGFvrJRy7Vabs/nPq/QNAsMKvWRZqZWZI739wplyoqP
zSx2/GjxtILoAPt1KTkqZJQ7Rd+M4Dtus02ZAccn65s6OTpPQeYZqRK5RLBch4aA
PTuX7UFDHBx2e0r1XpiYHzKQdP1TNF1MDFH/Dsp+OfFMiyRsFWHF+7hup75ZHFYf
l6nZ5NRd7imsls01rb4wi0z9lg/b9SNoKCz2WDcyuc3OKSaz/ERHSZCZZNqlvqf6
x/gr2RIkYBM8Jxu3frTw7EifcrCUF7PcN9GbzJEUkMRFQoik08RS0up/7sy5kmsF
e3vAnDWunzrdSrpThENNmSRv8rAzRj5/uEF/ffDJtfhT+EENmTh0vU0WPXKejrsl
Xd7Mqc/OYl3vFmeljsKad/6hjctRAZ5Ai3/HzZ2VyKHgEweaoq1xeBSELuRRoP2i
0jQ6BDS6G619T6hU9Uf0KS0ilzcg6Rk8NKHbRcjRMql/5MD0gKmbP9xcE1Vgy43b
fQji/j5GGZBcrt5s/xWzaOnIq/VBwmxIa0UvDJ2mjzyrbGjup8ykNIf9wC0HmZyG
hRH4R67Jre3N3K0sZ73p1pcVeRJ8KgrsjvruLDd4OVWtCFDhal8VSemSf9dTL5kV
ZpXV+sR4plhbSQs4LWKjADPmleEyQ87a+IHQakkmNg9/wzTmL8oLLBoaTEi80eGH
QTkYslrXL50ijUfyflYBB1a9eHyKH0ycs5gxkoLOlBE9jYCP0RS198d/WYmgMPIm
pX2+kSZEoWXn7gi4/yMY50kWlam7hI92552ZIEvnO6ZPRMYwmwqYOKokbS/yglac
qMp6aYEPHj2sOVbvBROzuwIAigvwAwUQYgTJDWDYYyrTOybft408USa0WKiCgcMv
aknchzEPhnzgIsY84L5lXGzX65FmIGMYCvnLt78UsMO69UiWpJ4OAc5lQ77DioJM
Gm3dl+JMmecTzg0wvykRb5vk7IukP53/yUtKn7tEXypo5olALfcpoQ6voX0wGHQ+
kx5XIocBnEWXM0qx7rr40WBDZEotclTlNK0woQsXnNIwCijg+VoqLInCWtQQ0iKu
7wqw63YMPxQMB0BhDISB/mCmqZN2N/vnGp9+V1h7KvYYTMam1dMhTKrvLglmh27X
K4wVUZR5HxW/dfBj5I1hSfAfC8lYKKrxPMd4N+5DHZtq5+RF9D2JeoYixYxW2QW/
NqNN4++w6Wjymu67Jb5aDozfsbcGzKy8yr2F1j5bNp06K7PFLuQiiMs9xSX7DICR
izsrXetcryuzBYrHYjILYHBEic2Mi9AJ7qRcjF/Nir/ft49MXYdDdqrs+I3twWW0
498tIzon2d2vNPXD6LDfNL8LIu2DaQUuI3mjVMn5Ess+MUbbO0h4BzSwt6aV8hC0
J/zTWRB139EjKVpN1R87oQgC6ecYDAfjT0ruMrpGpROQfPP7DX07ReccERe5kBlj
0GRz1Upo3OouBJxIKGzaFKedMBYUQq+mbagKCg4282GzfH+c6vy2vZgxxlya4s68
7PABG0XPFdOjX+Q9qwqXkVyQpU30q4GPVeisL0faiVOOte1PeOUnv/xYX6ZIbj7j
aDsjvgVac3lVLn+ZVuONwz58IIZmbwrvOVW/rrWkSJQT8n0o9MNst1etJBFhxoKc
s8xWSIX/X4S6lWaFf9++hdOtpVz6vjMTMNTSeu+0i9rGunJ3LIHzrBdxcMtdGz5J
7IrLfH+Vi02kpNt2p5lxm6cF2qHY7tAPjqRbmHwxkSiefdxzyS2rtd1SN7NOe3HL
2wzVPiup2ezl1LFg1OY1osLXEaXUTAz6RBhS//UBp9JXUBUflhHf8wVVfAqtEMmd
rwHKFynXqvu4ZncXz2573Z4ed1V6BKvrkIxDX4lWY6xcafImD16RuNXnDE71/8QP
6dwlce719c5c1/C/IIPUN9R5P6f5NzNLxjbu87zEdcKl2t4rAx9i57LLGqPFEhCI
OPoIiFPLgQFMeTVlVqgsT3HPpkVnBoiqA2MhquePZJb5PDDwlfCoE8TeWoRfqVke
tMY9i/XH6EKf5g9mbTFs9mbX1PjRlgwHVzGNeFUC7yausQMFUS7OuR5b+xrhO5+w
cJrQzTJ86izBHe93Sb/DZtyd1iQjA0v6qKr+v7Dzp2/AI0aRwDKfTrseEYWGdp8X
AA1ypgrLeuyD/tdBOnqOb5R5RxTAT1EnKTBd4AqIvjvEH7lF7eW0Km+ShT/DC3ul
sVR3zA+DK4jpw7LZP+rwTkx6w00G/0u7C9oU33De8sEgsWoZ4LAmzCKsnz50csae
36/mYMtXddnag1owouy8oiq/ixteK/Do+II7AehZZLRpYbec57g8PM5FLyqzipNe
zRTyOfC9l3OwC+TD6zzBwwTEiSWbpM2BlZH50iJPdjLZrWsSRBemXHZpUJqbLiTi
wMo8cAzKqjjBy09o2eilK0rcZKbyWQmrLZRHeSkwwv9Nfv9bG9NaFEPz4yLW9VO1
RnpxNl5i1mT50Zuq46BMYodxLJ0raGY+jSlacS8+FiqeAvOGnTDdHyOIg694iW8x
cZyWO9LsI8Q0pX2VB4bJlsnLRIMH/e504vnUnchx2/xlTmsxTUnWvn7X7CYXZnQd
M4IkYze7R8i0E6LFp/0GG+8lyIZCsNFvn4OoVtB1+VjxmNj/shhZdMgnOMbIYytX
iUpvp6cpvPxL8XiziL3lilcV6SADV2nYAGSKI4zZDepDS7ZrfEqTVt3ET3Ygco/k
qQmHGQm06RwxZ6RxEjBKtA/qBCAEI/PhOBt/BkULkIV0wiBP05o72OwoZkHVbBE8
TYNavo35toDemF96YURsfFqFaRPZhkx9IDWV2yml/WMKEoYYfndo6k2RkJR5zi0/
xGMeQEe54PeVSjHZcIX7o54nNMgb4F428BZEd6S40LgPFt6rux/HSlnSlXh1YNsq
MHAzVYR7PsCsr5QjxsEwMOd8YQSLENyNmWQxGAQVqWlnwWzoSGwrqu70VrpiY83V
6Daotp5UflcLTEC0eSjrfl8yNKQ11FjxwK3aT5+pI5ldvDhzjVuUQLhPfDxSozA6
L69Nre00sDPZ8hufsM5A0MXSLMZPXwOOsnWEw1qiQdJC9J+PlaQiZ+cOsobZBpgB
zNJ4deYGgr1P+t7uAjnsbniJwyo2qoZY3ZfwYLQutXrFuhYjmmE3HXr/f8uPpyGG
CrdNBKUTq9PgTQwIBKSOFOmcXO05kFla6dTBIpEU0AfFKUpoOfRinYlwauqrshfQ
L/lFm1kcniHR1hAkBM5zHqlgCKQgjyfC2/MgMg2q/9lPfkDrZ+Cq7I++nVnAyd6w
XoC87/zRBXSHqM12UC4ADucmxRZhMYIpi3X4jjr10rPoaVEGRI5z5MHi/MW4Nrl4
LZem7Q2cHNepUYDYbRQIpma1D1Mk5ZNK3C4R4AxGBVSmcTQMG1h9SQBzZJrswzKN
MALtiw7yQmg4xVdWjyC0IDKekgTXlvOjhCcw1iTFZo0dxF4HHcWOhrNxV043PN4t
/RLSbw1Oeh37OlZLh5a20Z23L0zGycGG0fEqcdUVd0JNzrI2UMJk0r6dMiOj9DX/
EuvCSsmK2BcbV1ME3u87iWbFQCQuARNXmC6p1eolPNc9sXM9HU6LdtX48RBZsl62
GG6C6Vu1J78PEhmpFuidbb04IhGI6CRhfjdq1ggZd1ZtKp1AyB/Uhhc7XZKMfNEr
VLVOdB+hdltr9lRsxVjJ2JZ9PvuAvh9MgspzWMCRThhHtNcRKXdhJklzwi7W5PO7
3Amtq+fnj/Q7fLDJd979q6S8FpXOJFPci/xYrzMj9IEM2u4BJIOMQqdblnz7okM1
bvLq6zV4wezdwpTSzC0pqzJbplC4hAYvYi3ihlKHoLm1MEiDa/xFtRqjPUm54QtJ
DpP1gmieLZqBCB5/G4k5Kvn6ABDsgmKWSMy1+/mq6KMEJivzyNtx3Jmd9IpNBt+s
fXgEerjiysfnr+JjyTBJdc+5qDbg/prOTQzDz1djZcRBFZ8Y0Op07WkFBz6bjoI2
dW/qyK2syPZZc5Oq/v9VhvOKOkJ9ZCV3rDmA0pAuZ6HWGCr2/eXz+Iq0xLeMNdbJ
P3fYzPuXdxQlJ2oLaa1f683I8+mnHQD/1DZpZPZ5MjHMrnS1UrBlqB/bKOd2BfcY
14XRiFmBhAu8PkuxEpY1EfTrpa/KX3VDoBxt/s3u3qZshVilzbCfaO8aSzWGv3u1
cyluqNHBpaMLUPLuGOoXVFf6URwRULzd2NyD7KcXeyAexcVVsKK+WrrO/Lp63aE8
XQ/wlPBowODtNNMJAfRf3Jp9Q//p7Wdmy+SQOLJIkOxhdyg6Ne2aASn2SPkFAs7O
cwmX2hUjOAwxX8t9tuwK9Xuof2YDR84151TpUSin7LmL1QxwTxKfScPQ1ATQx+Rh
I9u7ciu+CWxBLuzoJlizW847R6POpQEgnyUkYeqJpqK/uKD7wYrz/k/DzLbqZXo9
y1L7RTxt6hBZ2YMeQ+Bi7Km77PsH93UPzPk3mtkvvv9FYSkRcXD+jiVnL3iE3dry
R3FIBickZEVAVlmPLWuUxSyevXI1r4J7JxOmbV3g2pC7PJolM3gKtHu+hgriCFW8
ehUaLG63uEVFqIasrtXjwleSDEYMS5YufQfhW8ZekASASlLJs6IF/dUDTLxltJ1j
EkkoJXqagfB/eF12XX/epJZfaNTkM9OZeF4x+Ky3sgb0tgOt5ueccg4Jxl3F/YcQ
n4AkemZASTUN67dni56GUX6X/86QH6FNh7KHv5XJV4BOPjhg8rCwZVSwAe0jJ2ms
EauL1bWoBTat2IS/V8ppf9LTW0D849R6TjJjKUHZ18HNO9gGkZ0lcv/A+eQtyEju
Bw5qqhBzGZPqd7yJkrxp6s7TuAu6DZLXLYgehT8mjzl1q9c6bFYGl5E15qxVETsI
egne8gnt5rHsmNKyS89rNgRO67wTm4cqc7lNgrXXVLNYGwd4AjvjvJ4H/K4Nx4BF
eZXsZFOif6yDoaDnK5/zVRyrzKGpI1hDFvPiJN3vaoOFHyZNyFNywgTodq+h0OhF
J4dTtIyaZqWeVbFHAACNFNTfF51qpDVZVoblw5kOnDpMLk9R9le5ETKKCTQqXgdp
gYLcNC9vlgIygjhGF8R+EgRiLu0koOt+VOLfQXHfs2QqKXRBYdzhm0oTwVf8qzq0
CmyMSkjtu9ICT/t7uK+jYNY1B9suuynqfRyi+7IKNdZFdb/q3nNusW2YV/SD0ARj
nw2stg1ew6sjm9HMo3dHSehMHjjIKnRaSpHrE/qdWD42CLcfsU4yEExVTHM0XqE1
y4z1Lk/93ruoIXUjoPnuxs+HHsv0oMDPF8WXT9rz+1Bd5DGNNYfY9X//7dRA14mk
Ybx7pWY5/46aiIiOSLxsPeXkNvtSK6WBEFhivnrIE07r2Lw4F9Pa41+ZfPXw+O1c
vTbLXdHe61lG7YcH6LaGE4qQ/+WSWAcVaSXle+fOz50Y5YhsHpt1YsxRdP290l02
RY0Ckq4fmre5CQfkzkDFg1SxBTfkZd8ytVgqSfzdLq5yIOUESfY7gstrKXSg/vEP
ND20ySDVa3uxi9orc3b9YdGrYJnpScygMos+VdvThDTOysE0HBcRl1VXlT0gNxDh
4vXO9w7o2xxjSa6dQvfp0ZnT+H2EwQBTneLD2UGMZEMFpwQD+Q7+0dz4LEdbZrUI
kGWGgwsUa4X1h9VQW2VaROdKisB/7c0O2h9z9733RdrnN5yeF3doIdPYTa5ZdP80
jFoyWCquYnF9WSEj5HA/3foIQnc0B2a93QtAjGeKvjqRIT6Uz9Rm5rRqddVEvlsw
ciVhaUvVydMhQIpnlnEp+sG3e/nH+PaKab7yqjT0sIE1XRax20iQ67CG03tTJKUH
A+LLzjRU/TONHIig6kKLih1COBBLoXHaVh/fmJLg9JMwrflb2kYLGP1lE26RZFlD
lyqxreBYyPGRU4fCzRh++5YqBNLre+7VSYMMx2cNRiV10O4wkQskytkZrwAzsGKq
cb7ll5UMLM9ijEiGKqnYXfZ/qGAJ1RRdrz+pkiE1h8pMv/PqwcnntpZJSaqt13xN
pQSN7t76KjH3GcsprB/QcTiKkHQ4IscUmLI5ib+apZYgthkd8eqAX4/iTFn3qkCz
ojWvI6asnItf1ew4xhtFsX4pPg9d+M1wdagDMTUXRlGerv6nnGgpIYDPUgV9FDrX
JQkZSuhQ/Qp63vE07TspfoSUE+bm1G0iB96U0L0Nhxx8L3FUKiE01a03BKeiWhRz
FDQJjhUeXYxBDaLBCxF1tTBXnbs1N19613ZOufX35YxNF6Jb7QrHz+ux4butZZvf
WeAEsp8QkPL+mNa31XeYRHfObGZaa+iZcvLAJSIm6v73gDT8naiIZ7pCU07ZoZ/I
tRM3YbP4xUSBUjVQ+jM6+TrAcMrUO6Q3JqoPTsv5o3W2Fv9+xzZ1JZD3gopl6KiV
FbMxh+LXIvUy0uZiu+0rg+wnQ/Gv0s9n8VFQkCBY4StHbBlxGMxL5Pot0EC7H/gi
5Kocx2OlefvePOm13LEAsLJn0iMBXRzhIdMFTAHFGpXADNBjAaAfBVLM58WIqt8n
XtsV0k/y1rS38ih/qEr3JEpmnr5i0dRx/UozCSrkaeD1k+WqL2HVJGxV1iXk2HOy
d4VpZ/WDQ2DAzP4LyYj8gbYuPyzkYgSr/g6aGWPjpXEBZM3r7aaDGxUwqUtBmm/A
ke8RXgBG7dw3jt/0ulmBCqEFUCKqrna7J8+xedb658+wfX59eRG+LYXchNZKvh3V
JnkwnwGQtqbY87UMOxUMx727V89ZvinbVKNpmN6n9FbO/sEij8SU0YisWk6zvlQS
TLvShxV2nmvCmFdNFAWyQRvvwGLAIK3TQMOR5N/1z6L4AcToRc55uvBkurCr3bzx
zD9NWI7qzqqpvhHS7p+ddkErQ44nD3R2K9svTD2XfQXsOIyh5T7zswtCXc6Ebaio
fzIaD4YtduWtSLS/fNr99ZEW5Ukn/CqhiLJwxE+fmyfFRY4C4pUNDBKAGTQIK7bA
N0UdNbcBmNGlrRcEqLBsbIfc9HhwM9JUDCRA4qR+YZhli1KZRxP775sr53ckcy6b
ZhnmnaPH+qyFy8wGxHyvM24qMmd2JcIBTMQPU8tKyqFGL0EZ25vreecY9bWcK5PS
n4VRcK4msaz0kdlQ4TtQeXdB0yJczOgZDt5SCaZ9gofcYR1qUZQSNPVQzjpqz2zU
+x/PZVWsVqEdHTNof0W+KDNgxJLxC3YHBqRlLwwbM3kv5LOPZljOQvjWFcveRA3K
8lIPl0KY8xNtG3W6IFDy2YUi2jUCkX2aK9LMQNwXZFY0uitUwMncFhqIAe2tL0Jw
qfvrEO/D9y+VUpSatgjBIrnxYb3kcYIC0qCJ91iAnwGxIwFF7MLQyvlhT75bQzJ7
KnqKYVF2RngDrb46mWVwNE+8+9oFN4Xu7kS2c14DHXizkLxlAOdTPOF9RGS4/HO0
9gXREu3fnc8LiLLXC8aVQ+zXv9KrGdz1vRjQzKiwq8gXehKORgcIj/ooZ3slgSsg
UffDGAeUb2DJB6oTKh46Ered3XJKdZmkIEQ2AOoTx3r8nG+vuKwVo1z4XV6sGw24
BADeKxDZ4nnBxarhegOy9LwFWSf5gF9IfdyOq+eYo/jniu5kB+fleUaPQylw2od8
DzoxXAVYxPfDHYCHBbUWACf3g+PX3VSObPkzdNRi3+Kc0Jm22t+/0WL4hzebuL1C
7MSnuxVGyP2OR4yn0AttDM7tzsShP2u3OqXQLuHmoYJnnLWtYAkMjpWA5XHy41uz
9zKubcLa5WWXDJsDiqjwgst5Xo5qBP2m3gH5rOXg/Be3LcVHmAuMOPl1FioDjGJX
f7BgNMm/D7cQ2DHZCFp6G4VguCSqmWJQrheYrKssC7LfZ27AmJ6mXa12Gmv7dArf
1M8Kz8iog3uo2rPAANa5VseuPrtqHFGEDMVy5KmDUmmGQ2q+kmRKk7UuS8sS4TUx
J8493NPneHEMN6vUGefXKf0M4PY//RoymmNVHT6+hTQtu1r6D8qptf/Mly+E1elc
mqX+oUHCENOqTmY79y0BHWWpPvLnrdyrvNSD17ANr+zLMrev/v1vbohb+Pa1DVJM
LscNoyl/M3/st08usiNabMHevFDBaxvLNsmoQp+tIi+/spvvtKDgAUhDEdx415EA
uMgDCLBmnZPIFFnF/jqV8yXCESVzGzQkAnaY5mgE2DEwPfu7nQmHWi7FocEEjKSV
KOh7PR7G669IcrfsApHAklk92qDP//Bb8cu5J9so+boj07SzF+Me1Rc5eBmLxi8t
2+thJexqF7HLkP+XynYVQtnIhYwkzaB1rSJX2AM3rb2Bx+CjX9dh4LAjct6wTx4c
nNjrS+N3i0RshbD4z564PThjEu3h36xVy6xrSb+XL94e9aXXnlQs7L/6H8wV/Ezp
CsQw4TchSzodXmbY1LrJ4E18LoVTe75vxvq97u6b5EyvMkXs83MjSH1tfbY/oqbd
m2GFx/3q6ZF+Nh63EwcDWCe1tSlc5rLd9hNSYv7X8QkIo09LDcCkbh1f10Fq4NmW
3QfZwd/PV/0Q1ZDneshLf3gVg5UcJh0HzyB37CZgQ6BzWgUn32p/c4KEvGVFN/fK
kJGZ7tclQs8DC4jleKwo022oYvNi29ItFsO0dKP+8ylgztMdqaep998rOc79HpZm
PMjpEAi8B1py4xwD5NZyveUzKhkUnemsIbItxjFyi7khlCsXAtDH9gzugs/rkO6d
aPsT2X2FCtCheDF4O1OQImtw9Mty6dA9smEHj9D5RiBuw9nULZR4uaz9NZcOFpYM
TZXw6Q+SsihogM2AXTfn2CY1VTT1KBlmDzvH9Eq2OUyKLYOuQorWge3C0Bj1s9UI
0Bpbm3pJAUijCADIJM5ux+BVb33Fz0OOulR41WDXDK86oZYfd+SfXx+b1poUeWFO
N4AFdjKzLB2yyFzUiSjn6GLgK38UChUDDI7JgLpf0siH11J/O8tIC6wKgdNcfMw4
et42gUtPTYcHUPrVndD2tqsPiZDKzgaPSy7Yj6B6KWzV3nfNlE+QCiRNrzyapZ4A
PCOCB/cz+XD0Bt34h4ltdRD4Mcz1l4A748mGcjn2tVqtQpaO9YRUJ7P631RI5kCa
FBoRiwJtGG/whB7YTnDHVoZY0QdvQnLase0zFcbEiUiZSFpnB7Skwz1W7Gk+50lo
Bwc5L9ApRg1EjBsEWgid20GRiIbHsJXsh8IrddNTQpp2sR3KsxMQSodsLWS6rFul
MKLb5neiT4p4iz3aGcnR8VAPJwOveaizNbAMezwqofEz4cgPvGeigL3LcD3JVD3p
IYpolgsOt2qdUPvPDIOSnziqMHg50LxR0XOzT29mHFmzLDGYs2DJVQJky89phQHQ
8XavlrjYiSEsP5eTrJ0YqzvzP/BiIlZsiE8tjYRiRVxCrQnPkh2GK/B5qxYAqPej
BJHsW9dKAr+F1Y1lTlSYrfd0Lfidcqu7ax4IC8ZrTUJ6UaF1eXZF0bp9bBScHYAa
g43lQVykRwLXGVZ3sBeFo9FCM8B1VLF+4rGzXczR0wD3G1PIXrknM1ss3yvETpcb
V0VebTmQSueXB2CJy8mn+32O5bHQoO3KEAsbdoUp5ZwcHXVq0W95N63QYkadlAi5
vhc/0Q0BUaOpUmK7FPzbDDFPThqBpWVGfqREwGCwRzMJCAeJUSGBNmxD/8mpnGuy
pfSVSTjF11vMcRdjBHMFX2wXwi1S+vjQbIIONtE7ku7XXF5611gMXmpwWtsJITBf
DCrj7anT5TXLBbAbmsVR6S4DKC6bA+ILKovRPIjo5BzmSGLeSV8fseN503aXk4j+
P/iDxIDycDkIBSIef/C8jkmlXxE+S3MCneKWsX/2Iwf80QLhVct98++kUYUbuCGJ
rQZNV/CkwpA23uI8vMElRlvwBvYkqC260zoQvTUX6DK2/0AFRT0PO3p66437SRCW
bAga9tIm76mbsru8VSGH6wqldfwAJE1aloZSzRwLdVtbCrDIfe+ujBLB53M7A6g7
UfsQWY71Wq628Z8fw8gBagalP1LxHOeFmncTXt2KK5XVqPlAmioJvtA7O+87bEqL
dooe7xWKYhgq45Iw/NWYoHW91CLdQjY4WR6nI5u+BFcW/oUIBy40RJEadKJxzQHh
DiwLv7vfO47gqKZJZVKFwdn0jXxsRsbngdtJS0bDHxntWTM6Q+XMUY/IFQBrKBfy
lNZjsAS2gDd3ha9G8xRctmYlul841kt4QnX3TdPPnto8D/V9qxs8uWUphmnaiDo8
+93rxrSJ4r1ba7GRELhFJQwlvEFZylL5uqXNsFbz5yyR0YTx725pUZOj7LO36Aex
We/zTTtu4pTZbC4k9VHJlsuVcLj/YZxZqu5jnw63Xw0zTN2lcL4b+IS/D7AJYsh1
zOQBY4q6a7NTlsjoqBNPkppezYNNaBMhvC1RH2WlyC86WpEExWcxvLIwYOHzvxKJ
SvjUfyxnb4Eu2/wtc0G8z92Ghr58QP55kqo1OboSg5NA5OO2m77TABamMgUxdU1W
UOHtz20fclfwd9Y9Li55R/QkDQxNcHLlfGVawsjSxdnLKfTzb5wZwOEBqP8Z82I3
UaUoYMKNFG+pFfZ52Tz3+0vcdKphGRNgFE5giKM5Pfjlcj78I59HqZWYhkIwqVvo
AtpRgKe1R4CGs+oFx5ZRcaVTCXIQPmSYFqeVMm6YpoWoveBpnHt8E0NLAZtZIHBB
/QKGiIo5vMBgQ6ofJQKQc5/iv+hotFYIZMhikLDxWDZS8ZjENqe6ZswqAzWyt7et
QMCQaIe7N1wfCZFPujf3fAFSCsWVA+voyeAEL1Rc2MD+MuezA339QWdB1qsX5dU6
7FPZJoT5Jq3FL6kwzb7E/5ss2WJNSI3UdxYDpFmM0g+VMUWgA8h1Q4lLOC7IxCd6
t8n1/FGBTPS/A1HzgBifIdYq+NKfp2bfbAv8fKj3UyyOcmRYxn0iEmyKzE6kMa4X
oGnoebInLsPUNkJVeWQUuVd6POA83Y3WwHCfrFTI/hSdM4SZzfQ4sIXgepjHn7/F
q6bink1RmP/WLw812v4PGB2rYV2L6CYCuDapsNQGVPB+X7NSx+l5W5Ai+XoZFzyq
k+48/iOiPKYozzDnGNL2LWJTNvEz4RuIoVirnxec8Pa4UMvokKResGfXHjwTVnN2
K+aRdxahMBrfz9SN2H0J31lsrdPBVC8GacgBsWaD7zhrBmEiJ2SosvF6Ot1bnSqH
StjKILdGUFogyYT91hwnpj2Y00OJkj596U0QZqtJVKzWuEe/A/8ya8KyQzFm9Z8h
nE4/3Gtx/UVIIx16Xfz33vWwEBlyFgdTCthc3zGWiQfMdom2KZ2zJXSaUuKE/dVC
HOtx248XQK2TO+Yhn1cLcm+WdTVpWQA3rWXxFYC6xGSuit5c3rrtcGTI3rYCEMkg
9SkrhmYgqDS3RxqLjt4NGm/Szek1O/XNaQMBqA9b5qy5LiwCQtxpzQAf5hG0pH1d
kkA8rD7XAwkOCgLpfAjsXuuvnuBURRtjWHJiNq+u3ajwDRUuknclZHBzpvFi6VnH
0pvlBM2kupit3kXEseE0t4/ZsVa3e/5q0qUQNmRFM9rJ910O2H9QU8D0UAnk6L7T
NfRg7dAvK10wO6QkScWHAG3iT4J/AMwfEEqynjaa/RuE7SgstDsCSuqBMJl0Yd6D
HPPDxd2Rri7Odq89fPyGZCh2e/juzCEfr2+cVcok5g/0vGZO3mRakwsAd4MU/JTl
op/2x011YOoqaR+u7UK3epTHgljZlFDlUeUDv1ufTCjvggpfW8ti6rFDgHhGwkxU
geUtaAYMiNmvDGyX4aQaI6RImAgxJyzZF/YkrMTz1Ao49pH/JvrN6izHwD/fy7Q2
6tplre1gT858bcRQtXeWxak8bGE7IMBdpE5rpL0yKUOL5WZQePMbFqauq/w/JHGM
wzNaSfTVCiMoPagU8k18ZKzDHjgw9SZHCNHeUpssRHydgnW7UiFLMfJUAOGasWuY
VCnZs9irSRBja02B8Fmh2TU1CE3yULZLzlqjYZfEfd0QRAheomj9EJcPAtHPjue3
paV1o7DODDdPern57BGt8iWFxsPMTIICqciS6wKrNGC9AHOtzdLT/dOPLnwJ34TL
8oQl1JqyD4tPIOd+ssNEW5Vs5uW7ys+nHhdTg4pnKz1bh1igtDCf1KMtXR2fwyYU
V5qrhR4pmuj7OD2fqjvrV8X8wVIGhBOXkecENowPoJWlPW261SN1UwTjqYd/qRfw
HsFcLXuzDqdYgr5Ubed3A/gZ7yg9Kg8C0ANuq9FS9kLWTZ5y9b4+55sNQOl14z6e
SdiU6pv59VwUN4V4Kj0CwgWiqfazYJrAo02BLgS3jIK6m0oDjuzMTrCvxHbQhANf
QT+E5EmNxnoNN7dJTQgWRwPYkxJ1XECrv0GAgmMnui+Ej0n45N5jtPftMgUZLlf8
vdLFcs7Ia4vyl0MI2PnTj8fQfn7sp7MQhpC1q12kVpX6/wHewCRD2QZb7h0lLn3t
iFgZZfgvQHukeIHOXoFtvelfEdw8UhrX8RxfRiPiqU833mtP2oK9zWF9c6YvU/rl
Rlh8doiB+odzmtPxh9G6AuFRTTp9s4lAeaFRk/WNPWRTgdOJ0ULfSy+T8oL+A7Lx
5/LpfixSYXENhU5miFjxZjkFsvtLSCSkUa6whr6XHobyp8LJ5vbr3fOl38pnCKV7
5/YPXNTpNuwniFztV/cENxO6XfNYXPlS9nqC92fTxd0974YprFtUWddP+D5Gz78x
22Hjz2ggstYHMIks0ax0PIpHcMa4+l+2glgyfej4hFcCtkMsnw/qm/WXI+no6HNp
PrmvOfBk3sC17NMp7mhH+t8riEOB+2ABYoWG1/Xt3NlvPjNTePxbGCW1/sBdD34p
ECi14vbpy9LaXV6NSO7WEFk5rQxvfVIJ3Etrig9Lz/vsGD6tDcnRbo1Fy2PIlTKV
WPDsELHDfTjgZoejNTAHPKvEen2Ui/dMHZFUWCcHgJOVA7iHCjTvP9CVlg7PT2x1
tIX09PIw9l0GK+qswFHFJuZXwJQpjYBQlXkcbZNbryRYjJVIzkA4JPbUSKqZS50O
HGT4Iyn6DSWY6EIoct8+fW+WAOt5S/AjRXn/Ns/7IV0Gr2g2Mu7xDvGx4W/ZbAvv
YEDEW5yNXAPXWLcrPu/I5uyIDUzHhZQikwgJ6Yv/0IfWUduHJ4Kx6fUe6yfm/+Oo
8wnnwPqGXgpyzyeEJQu7kXzHCshsJA/1xyXnpK82uDd37zSVlI1gwR348INzUX9J
1lDSYJc9HZ52/7z4l9HkBnedBvb/D+IHYFHjAkSGSmFul8UAnUicBu2sfpdD7GVB
s/xXWCmICuTWvpcY3oV6I2jI2iGpCtUQLsWDnhb7Bcmzc6Fu3k7tJxH9F1WttUjA
cNcVdloix2n/9CE0dcioZTy4/CS22gYxbsbcbdNutJe82cm1VJBMe101RouIAcX3
QQJT6RmHGI/t7aA4GEfL8pBIO2niSaW53GqGvj4Ivzx56owtShbIY2rRlZszJbdr
sZDwXJyBLeZHIONXerstNNFGUbVlBN4EV5I2M8UDPHXwRDzZFmjpXux1ycu59wwV
AaJlMHfHuEgrK684RMApWRlWvHXgDqrKoYYyD7Ilgk7KHga1FJXq4yzXSIyQS61R
BCHHIaJGK6AoLK7PSzASSqbCiLOCJj22yiHshyEUU5Rj8fz2D21/j/J0SX5BXgPs
r/B1k5iRVT+my7A/HmLC9x1ifqfXqlQP0JAT6br6CmyxwrkT+4PJEKmYq3N6A+pb
Bg5l5A7RcuGn2Hn26gt5atKDHgNoh4PVv3GsQfzw9k+CzpPgeIRfyTD9TsY+nsup
L7cbZFvrwxsiEVav/SDKAyape+Z+Zv/UbtWRo9AmgmTGSt6xWQcE2KL72KZ9jdXF
aTI8N+ioW2ZBhkNTlQU5GfVw8M10vSDQ5jskXhMbslurl2RUT4L5hBTFgE/sn27z
29CU1nlfu983JrkpRMyFQkeJ/vsP11r1tL5VQaGS8l83MRjRxscD+5+35SLp1pBf
5bgE1D4VqgbdnB7nUK9rprbTowDPo6tmUCd/6piIN+RhRdN3glyIu+mPNS1OWijr
KVe78wF/1XCn94mR7M0ubBwxxry/7q672Z2sh4LGOQXyVCAWo+V7lMUblA0xmz0G
DrwfhbbBIvhjV4DI6eKgURCpEiwwAw6mQCB8T2ppweZusoizOnIxX5Xp3oO+C+Ni
Tb6F8J8UXPycTmbT5Y3/jy2jL0ARgPNKOlLqMNhefO08Q/tU8uWT+M7vwrvqfj6x
1KrAMBENMMwglYKr0+y1k2IB9aoCEX0+cUHCem2FmgsVjs8PVjPfXZ/0XsKYy1TL
xlxfcyJZ3TEja0MbiW5ICEI2vKIjIRrMN9z4TLSJkdXzgM+AakVBqTaQ2+YhTrd6
FKYrWp4BSOEUAUSexgJlKQ37SbPF5l+b1GvoLAiHpxFnErzy8WQGQHklb06PDz6E
tg3Y7bzxQY7F3l+2dQ5BM9knT3YIs/gcx+Dx16GQ0PFiyKtTDpJRA+vtFXDRSvzp
73Jue5mj80EVLN6eOkHROhz5h2Rt47X5+BoLWWtEEY8iOnXMYEH+CFNtqR/8Dyp0
8/kO1mfM2hUquDxE2tKj1OkJxT1q1BnmAqud7+nwdcaQYLbq+x8jRBnCVjqRA0vx
4Dpz4g5OgiZHrk8HRTuwgblEgwX+BdgD9P/Wqn5OK0RgzOnEdxcs53QSkqA2CY0S
ESSmOvr8jmxpLL+aFlSr5kQORelZMlkTV2EtchCC4vqLNNos2g4O2wdGfdrcjB8J
GGaHhaidaLzgSeBhd2e/GNwjaBgI6W9siMhYOJ+Ljo3sH8fLZnYw9PwBuAB+eqWR
MGr0/fi7eB1ODdye0dE1Nj5TgHHMKVygTW9yvYwvAfmv22xxrZ8om9KVyltbV3wC
447Q6TLjQfoq6w8erS/DKroWZ9K025sV0AfgAq7uicTYhq1vLnL4IJOdXdef70h3
e5l7coL6Q7Tc3FXfzFxxSNiCWyQD6Sxf5qpE45vqXBuNknOgXKoNrL2jYWnxNTev
q6YrC3YN29YdxvwrRU8t5EIZdoq/tRT4n1zWgdPSFDmAtbcJ3/77hMnknvs1NKz0
bBJCvq2CuOPGrDX0DSwJ2wj5+3VwZct35Aea8RSXcZ5zXQepQ7OQd+8PNQ0ZyUws
Q9dYZIXsnfrtjjZmIwIbVDxJW94tu23bI7PN4afDveg9AJ1NHr4NDg1h78h75PRc
rMjgjJPRnRqK3w3o83Nql+xp47mtdeht1iSZ4AXLyPFou3fY0Md1h9CwzIq7b3X7
VOiBu65pHvVrJxg43JQdTLXFxAdy6hGyN3v1Qlnt5WInk7AQeqatAnvRq5/pH55D
1lZmG0HAIrdJaVaLG6NnYWyj2IDEaGDVBZdbXc82SsAvhFAYU7nV4yAkb3rc2edu
PfH0rxJ/ECCiSfJ/dLaZLrOpmG+sY0ehv1K7NATl2nEpqx2vyUeQzhhPQjt+w1xe
1bBPP+4VEWwVd5vkHAmFt4JsldjV2gy6SBWmym/KUXAL7EJ4UJrBPeU5Yck/4Oqj
w/VsQgl2qkGoNd4qu8mQfIk9QaDSE+yzEpY6qDQlbJTlEY4H1UDIupMkfvAjNMY7
5NvcsnJYu9EI5n+LrP1WgbxYOIKcUsx68vdmV7HnHRoqOHag1V2XCA8YrwKdJh7X
vjPTUosRAREdIzuUe0qMqRwMhlZ8FC1KaMyyI0zitx5yb/aAVQWnBDNrwJLUX8qQ
AZezSA+1TkEOhZSRyAm3Fn1OYyNJGLytO9Ypx+ngM2mfKiHqIY+L4aGmKpW6TQVZ
28ikW/EbLpe4PI3/BF2xY2pmOkQqmmBlKyMuO5D1ebdFFPLgRRwj6NnT285dEq/Y
jYWBjVqiO0zLQz3mXUXr03Am/JLyEZjYDwUO2X3V5pWGtLLPPcFL/BhowD71EuzL
rUdwrJwwZYsEwgLjB0O8jVTrVTlNJYlUbqkLVcxXKeZmnUpEb1/c3s5NVhOh+927
JNg9ev5D2Rz0VSQqT7BVzCSmHZUcUNT98kp4TpGQAX36drc9MQ1iuWFv0VQWQtL5
LmhDUomVD7lO0Qb5z5xJ9UWVV8XByFGVk9tpJ13pRAgqE4TPGkgdb3Ua+SbQeWTa
l+vBotAZAp+L1TKWNw4PMreEi5IuuThrobLURR8zmkIXYsBDiGN9z1jIprmn2wzb
VS2dEb7ehJj01HC3W4cgejZJj9TDlPGGTCh5YIF08C4huTAwri4pEKEjcYkmCxgE
iQYIOe7V3/DyNxEmax9WQ0TyTbAhMO5kxHppt10wOi5VSZA2MAc7RSWmSZAiEhlv
hN3AlGTAgKqxJk34Fm+akbAVIcA8EqhXTxeXSANEZQvxikWuFs5jCsG9UZJAHYGj
k1FnhPNfhE1bsDfjycUcTBm4Lmg0fsh9Cj1A5RqKqSHgWj24egexxUw0BKl+NF0e
3yw+t5iIGqRawk9HY1t5Q0br7VATNG2KVPUBGYlxm6YjTFNPNAD83O85B8EySS4+
P/5bcKJcvLVuMfMtAx3ZdNpcx0ITMytBsr+pj0F1n7+eh/HH2D9nYDZkQ3XiIduF
2g9HL63tuNZki15KloZq58PtWDBS96ykJQnD7di1+CAoRzx+2nzmI+ejK/4HH/Ni
FPOPDXajDlUwiuiV/0dpvjRcKu9pvZGv6Yjc9NpoMd/OPu0IjyKVUcGtE2j+STOO
iG+zTlxIG0QVf/NVQB7iVytQTWWF2kmG/OeqMkucG6sXxw+g1T7Dkzqyr8vuoYaM
YXc2QM5zbjhzJm6zv0j86rqQeAktd1NGFYau5Zwo3UHDK/4NZz7SKrDe6Xd7ZWej
n61Tl0zTkWShx5kowfKhbLMwGF/4isfTUk7H71PGKcU0TAcY2Ye2Qqc4alEC77ZX
iUDw4t6IS6VncoJzDQXA6KvofacOeNBtyM8hx3G5JlT+JbgkYXVKAfJ/s+JEK2Zk
pg8nNLzhupQTKpriO6c5O+9QZx+CLrzOs1PccVA7gRQuuK9QLg7HhzykutARIEiX
bK4BbtxaETxdSJt5caRb2k8jtF9Ax3tYcGjLdJyuiUaDueergTlQAa4ndw/Gb5PO
oVmRfDBH4+AzZHETwjxVDIOWXUNGynkAW5eV8eYW96Vt2WLJFW8dvCk4FH4DRWSU
rLKP7Rvu2CgL8Ca1REwiQO/QH7E2LLh0NeTUon91A7G+tDYRlt2l/v7SIjOThJ0O
vKjEnqaoDMhCaCXSoIFdrPZZhVHOpOVPWYlX88C5KciEBQVxB87efC6xqs9rZDkG
Ag4Hpbn6dkVxGc+57+GZI5icbsm097itW2ZAhLWbMi7jMTHrYrvi0CS8rQVXzZ0+
RyY0jqriuInQ2tBGXgnIC5AlETw7F+jbbxn6HRUydh+AQ4O4B49FE0NvCepPJY+j
hzEhFLIU9auIQ5oSEpdx6gZqjnQf3+2nwsFBs36lvzbK5+9KvG2zlWTEoAmwCY+A
9K0FpJwU0nNn9cyh9lNGF0+mSPFP0fpB0CmpG0lRYT2FzATS0W/mdkhwj00BSSBD
9D5a4omzfdGaMKXs7L0y8TthAN93yS8GX9bIsNiGyL7lPwjyoFZRzzJjGmxsiWhf
ksbc4Uu5jx2MtzlqqSf3RGIweuDlFLFhTB2tK1dXFkdxTRepsB1d0/w11AgF7+tL
/8sN0e0Zzf2I5l/S8hxn94imW7i1huvZTkshdKOmQIH2kANbvhImAX8ZRdIk5DGR
dDeR366Gsfs13ztq0/Cvb7T06TbkTnn5Eed7OGPZ3uDYXWjD+lgJwIds5Ftmaqc/
ItFtmp2E2VIywzmXnMnCB1ylV93x4m7iANrXnWELlfyzp88qq6IdS3E9CNrkIbax
CM1/SUATlGyhH0JtTxMXgxmS+vsfere3NNlaOqrRtN+m/5p1LmomIoG9eCfR9Ay2
aGb7omlG28UWUrk/4+J8f7VPUexFK8bQLuraYzbcoP8TqOGvg15TvoiytgUr7YH8
0w0ra7ts0NctvdhlVvic/8RjkBCJYRU2ivhzlxp9doMIpep8jXEmz+kqDMm/i6/h
D/bYMygok38eBEeldGFurzMB2oNZHFVJ1cjjT6Vo5rWsydu3YScCiJ7c+DvvGmUn
IGwymg9fWnpf5rSb8tDNS8O3ZJ/jup3GofdiN3RbypGTaV5Fjhpb+3+Z2aNOvct5
DjFC8ghICm82wodfMMzERAZumVPJjS0gCm3WOTnJueqzpZfbTMwTfwrN6Bz9W5Mv
m2+DMCXqTJ79dlJBz8yzgt1ZKT93JKEzF1245/hiYpB4Rv4F+Ci2WLrmplCPr4zW
j4zhfiJ4RKU4TUy4852psQS4lT8I3xNdNxrAsuZWvIu4eIvEfBlijoIXunlXlXzO
4lpU3TDD17mS4Tu0h3g7UShX2I4Zn49PHwJH98CKQl6mmPGQ3e7oxVTzDnGoikqH
ECy6/d47xvP8EqyBIQD9ETYyEXLXePrV9XHVUc3NexD+xxwUG+hiFTusCuNo4ZPO
lSjs0p3PsM4xttjlAnqYbrho7JufpkSP8C9LSNzdyPLxdUmtN2+/IA+WfRWhm5WW
l+8wS+JOwtyxERs1lFR8CZkKA76DkHOSoous8LLQ5d6PmZ44aJUQgpbQCRsgpGBQ
Sutl7MUTI8vuuUFLkJOCnkmsoER/cwxY5TO/ReFwW3mrSv+CnX3HYqGu0aJJ4yl4
XjLrP7XcjLWpBo5RWerr9nQXEztuwV0kEnSrWAfaRrWu3J0Hf2jC5x9lzLvSJW6G
+yOv6rMF/4VomXARvX6jcOAakux1wJ+Os61rPS0aDorLVdjC0JN1n/MYsY8Kj8I5
OFVOSQ9TlkY4iHEFDBRyeiY79SLbre2g3nYkzJgrHVQ+oY5f7VGgU6+HCDmScE/E
aMGuMLUTT3tIGjEf9YwmcSUzOGHYrpJvcQQqclNqXmcMTgx3IfYTyacxT/ENAjpI
Zt06Usdd88VJlfCEnX1NHpwMr65AXQ2SMAYmTQOh71wPa7fY3ALx9U59ZXc0Z4SH
p1dX+9lGLEjXLBuRSg65YSJwxUBf+eXVd5HmpQeIXsuliPhLgWfBJXQ2f8HkZmcr
ITANhKX8W2KvbORNPw4y0tgIjM0h9MYBqMntlxaBxNr4c6/Z8oSZ6VpNdUMBQ56w
rUhWfHEnOMTLzExIiR+3NLP824elTIzbCv8kF7ugONvMu1cNtTnCeK7Id6uZ0n51
2RtGdBLFtfpDGzVL+3DtPMIOff7WJJs95XJe1WidNoDXquBZ3yH8qAX3vC1DaAal
s022S+9tWwAxrKDTJgtSehxK+EGcmXMySzbCs8EW8XSYh0RDnapVCmxXxLl6UCcw
nZiGXwqW2lMPIrLy5QssgeeEKllvF7aA8DL1yf2dQKGpWxbDpYQ/hQrRNFId5qxD
Ymkve1969rD+KghuzHioqcwSFxsuNSY5JmOHCi8U52Hj7ron4Y96UZfOG61FQJvc
6TClWnxpmlCeR0jDNhae9cZQsBHfjrRvmDCz0p8qN/uGrCyoREKQJsvok/EMnbff
ajmHFML9yJMfHI2+9QsuCgGFA/N2mA+2a2HRFUHVuKHPpB8CIjNFcaF7Q6RJhXgG
rxA+A5gPlf/VXQ0mOyFNDdTo+4Aublj0yT6rWbHSm6IBnOBbLawdBYWEpZWvrxHl
omtu/Xfl2osvCX1uTeTIkjSjpXJaBWIPKUd/xieBy0g65mQhUz7zRc499I/v+Ue4
DEKFdZOvhH/RPEJfyIdFUCpCVZm8nD0B9Ew3KUVrHI2eQsSIR4X8j413sOMvKULH
QxuJxKLfEogmVjYT0j3/2d98E9vwFRh40x7t0YMoZSYo4Gy2XFC8k/jIlpm5EYyn
3079Z10n39S+EWuvDfpSK/zHLrG2KGRBHkJR3CQt+6V6utOTy06KBjrsSH3IToJB
hadGhnL88PaU/rL/QsvpJoocd323rEFOko8r3CTicB7ZqyujP+y0mFKGAP8SWuNR
cRLmNmNeg6/tx00gyVs8f8GJmlvVbYfV4DFJTMGvjvRtnbyfgKzhLh9Xss8/tQ8/
j1/w/F2x7V5jwaRBmZyeOscBCy8qdhtVvopexf2ZcZqWhzJtp3SjNZfO0y6BZrV1
MIFIhOk8FHd80I88EH85+0VOKfg2mMtQVy5Dq+aH4SYYYPNjKTP3O23+ezHbYHGE
o9u0U1oogThJNLxp8Tpgv26ACUT2TDVpzYMia3o6JCEVGFgJP6sww940IxF4NfAZ
PhDE3I6W9U9VZ0SeReZhtXnUqeE1dkvw3TSnGK15TkrcSis+/tFUJKptpuRbMoXQ
KMMhOAhRD8aNcOq3YXIYYjKdhsfuVdmpTH+OjhUcmlobQ8pfeZ5jLSq8xUX6+k3G
fFuOy+477+k3YfDgK6C3QPVInQr+rF0OEJX8hzxqZLn2OWLL7oJqDfFl9oT2JHgR
fjqcPuy8LYa9/HwOTJzKGUwGWVwe8/6kjfTczDLdsF4fazlHDAu7JVD67T97ayuz
XCd/b0zbN/ScbgCXO+aWzflUtbTn1KrHUdOt55rrEyUz2U6dgIWyMWVdZLKmYgPu
VtbUg9l23/WZVK20Mx5oIi/GFLOjzGK1b8EID3WqPr1ZO7VblOnX2iDxbLRcL00B
9K20V1j6S+mUE9NBJINBjH0pz8pu9XnPRRE9TzxEaAF5U4gPmxtbmJsZn2vAqLWw
njVdDqUKypw7a82kF66HhMkFKAnEuL3c334ZYFbt8/XTYp5IjI45BWozUU8/0NAk
uI2HZ3sVWJtRstrDrmBm7Isa2Rtzj0MWyWxOu75XdKR6q5vVn1oQogV4bJQAXg5c
PMoppzvmL9kaPDj7fypQ9v76N6tuH5YmpDw95i/9Y8JlpBOBrVwEy6faKx/3DOoV
UFCTS0WIDfWf+0NVXn6BzJs/54Utr8FSKHleOx5cLZY0JW7z7fTA2oIV/Pxcxv0K
/Q0aW3sQsDCkO5lGY/SYwuPQLLpli0ftWEeMQCDPXWO6MMmRRStIOBi4EboowKJq
PW1XkG1GcX1D080imf9tO/3Yrkzl0g5MSTIp9pmlkwOUGVjsp50vsLBL6RRZER5Z
AFlWZE6ft96COubMeuyIFy6TXAaD7U6j9kT0S9Mipq6fVCiJdnVe6T4vJ6sQ22wV
MLu/yMZvnmgHw9oIR6ueH65t7VLIn48SILNQqg0csLucTzYaogHW0WF5Gz8L5wzS
9xzanctKDdfWLz4ekSJ6j8t+5v8Z9eSlL1aJ9/vQFoSvDszOLFdRq7LxfXdPpgUq
rJ63d8Ldt4lo8ZmVnbiJnGrdoygyS/77qWx8v6syz1j489vfM4CMghWn3tpm1saQ
KQZM5jtY19MqbkvIFkdN4dTekDK9X0no4uzILm5UEpYEOYmykZyGm+C5YPHXVlNJ
5IIv+5mVeLaR6YCaNLCB0iuXSbw7ICHUB1P6vnxKDLtymv2zAEr4T1Y5zlWTK+Ti
/sfIqHIMkxSi+eq6HMTCPe89AdEzc/Wyr/Or12IXcgESsbzO7a4Bz5TcyHL1UuZq
Cy8Fn/g51UEyrVvzB10ry11430ziHHjv8b53JeE4lqHJGlQm8S7+wp3dvSXkzrlt
ErR5jFlwWftPID7v6CSTIPR7qsZRJpC92LxTX5WywrxKvkDAU6gDvLBDG3wFHjpf
sC31bhK3UqupRb9lp2BtOsb9Gfx63x9pTUxW61V7h9tBNOmM0N/rDKE7ou3E7Ucr
vis4B+qS1APFVAntb7bhU3hMhmextyjyr7gXZ0Kclhc3/QGKViPCsAJgthDaQ+km
m4eCtuTLuejuP/loBtzEyAbgei7SnUEfqvWovlmcdsJi9ya4EkxET0/JHVvwuZvu
zklvneJ033djPS3BASc3KCHeDzbiZBXF83PgAHSjwwp3KYaG9RAmMs+oNC+2l958
JxiytuUa0jOrIrqFokeMuv4yvqhoAk+EpVH/9/qzpDyE6It3chTTXFSmEN/n78ZH
yVbmMJSWge96EM8ZTtgzWYSZmxluh4ZvhUB3J2r3xwFyVg0p87cEPwsnyXxwKxAX
N6CwoSnBnnabNTCqvJUzai+Jj0OebWcevXoQjrY9uFn1fRj8dQ+NRFIkIqMmWQlI
oucv61zMsvEOkB3Q4gT5rDQYGXTGT1cb/l3jJEoKSBjoOYLovHz+SyOZkVH21e5q
837k/29Uk10oKpoZ6yRC3Gg1qEgfkY5/zAv8CI6XI5GswuUgeYIHvi71q1qkK4mT
xBIVxSDjduzanNSw2VRepGp09//4r9kI1sjFaSCjMLlyUbVcPFN2aTHSDtS7Duf0
1i8PlXQCR+u821wacQAlFz6Fyupm+ObacTVqR9oDcgRQXL9uGT+ouHresv72ISZC
43fP7I4Utt2kFwyOocpWvxpRo0wAplUSYEvHlEfknhDNwIlrEjA+NT1ESxrsJnzC
OS18MXFm5pZnARiMOXBeLYLgb3Qar7vzsapJ7J0yT+v/N8agpZ+fK/F0yAou2Lal
uEhbAza372t6jbkLYllJ7Q4zTVRGOoTwrBO2Fh3XZO8oWmw84S1oMWjByY1kd7Hw
a36P7vni7o375nK9i+FJZ37FrlKBPHRxoOxSlxbC6xgAwGWKApwPHLZlYtLTUPq2
fJfXgC8XRLUpEvjdxmJLRU3vGgvkP0U/uQYHKC9BcS+4K4fg3m0SxPSjOC/G/lUz
LG4TLD6O27iRIBZOJbJZRU5Y0S21daP+ZHnt9vKqrHPYUYPdHQy/McMeKP+pEKxS
+N8MZurEQokxJgBD8D+ifMT2g84NenrlmfZE9m+rwQPFp/CiO/0n4hGo+Kvxxll1
OutfWGax62vI3iXHg5LnSRr/aYji0D5OEiIuFf7/ol0Oo+nD+PS9Qkno520cacq4
5WMU1oHuqzZUn42+OG2cuWgNTJRCkzR1N3e93zJDA4wYlwZiYgCKxzNqjENtnGEa
MuMjEfrgjKV0c7tNUZabrMyOtms1EMRW1NSniqOLqGHpdwt1h1cYNUY48op0dEb+
STYn9gLxBmXUYEPfxO/tX0aack/WHUnVQVz9n1sD+Wu1ez4HxJqLueRm1bI6owtF
uoPdPENwlpWTBloFbNqc/UkcIshLps8qZMoA2s6gLpp/4Rm3NWp6p1NEKMZfPmep
UDiGBcGVbsf/V84FXsZWXtHmmTeyn4xPVYT65q4Wc3Zz45naU6O/BJkbklvey/KH
SCfZ62yhQJhEuj9JYPQxS1m511+cV1xQwb9I0gCj6s6eaqVdEeayQ90gUAheMqIm
TAqWDCOa1uilxb0osoYs9kv87I1CKXQqOu5erbt7jbmz/Q6i7cesPqrbzwEl8LzK
xrclLCLinHUKdfoW2zOnIZsFcGlwFytv0VWiG6doB6FWCabZtgNZsASvKW+cxhVA
uek/BaeaO7QNRyXpLrqneU7GInbNtKXYKGevDtV1/vmSVaWxB9qCO2HtSoccsT6F
sr/XyOhiZ1VJgWVYDjRZMBxPJreXK/vB9zg6w0d+n1e2qqI0f1wOlnbndJMrKcOw
aapKcCbypV9eM2yvxUAmUEAtyzvdU8Nk46wxJqBxfgh83HYuWtxetONrBdevWsUi
kTR8cu6/zyksiRE4IRbnpCFVdNLCrESy/WCVrIAj0t2wvom4tXsYacR6qNb5/JJE
YS25hrniAf3qukYZjsELEyjhJGDnvY4Uo8mXPwN9kTYdsh9qG9NtrellyMluFRwd
lwzh7WWEc09/Hmb/TqAGaUIdH8oGZpLMCTZ5SiHV2IHWhTOtDHJXiXXzjPW28tDu
OUaHxnplvQeE+JjTwNIqA91aZJFheDkg1xPe5TOG1e/ZvH8sQ5D0xus94wBGK03f
EjQ7launehU53xRegLryO8JksU5i421kxDE6VZ4gQA2p3lRb7KGIfcK/OY9/jyT/
Weo5oVxCRfsvogaXCYbGeGZj91R4WjkmwUjjpdsHhexKyXVCb7zw/GgOlD7fvME4
AKxmuJyWl0zAYnqogVRRUP9ky7kpoWJqXXjDX66NINbTrRwFeg6IP3ibmHxIFsX1
jEjPXr57QtFPgbrTqN+J6NCojaUg+T9zce0hDce6f+BEHHc8rd8rVSMocW2p+EoB
VrCgQ8XzPg6uOZ7CDDN4jxQbjHJTFYLUq7zS3MQG4nzw2XbScD9hU5WtsejQkOqQ
HhnkuJuWoV6TYPuwGbVa1jeVx8Tu2AFeo4w5/EiMuoHxTIleI4IA2OW0c2toKHPD
70xjuHttmp7uV+LHCw0Wqe84SueDOlz9pTanCOlT2AGgqxFaq2Sa3Rin+MtLJvK0
W/FzuvDaDfySu0e0CAXjPmyhoakOgkuwNzwc3yLLdKVXUdwm5EYDuLBj4IarcsZm
KCBnU2UoZhVijYwFkE6G78ObTeVwH7yK6KK0JEG4ZUWJzqTGNG64r+4YkKIzz21I
8YvFrfGNaQ+YsTgTtGjQbNURA3T9eHa3ivlrIK5gX7eUVtuXPewVxT0hqoJ+OCie
lsttYqZU+WOg6Ug4zzwXzMMm8pYNcaY+aht+3J7h2/lgYNhwESMjK0akU3Xl5ECz
Xn1OMiSj1ajvzPQWkNRgPCqeBsCjTbwJO42oN9UUt/TrGWkfvjNMX7JPP+gsNWOW
AkI3dA04YqFJ/kQBNL/RJltBYgS7zFIMXflGhfOYdqg12tpUm/VDpPIHJeoDxBBJ
CWrduYvL/wURPZ5AdtMNpb+5RgHsFVtDGngqS8aSrbYDk8bwzrD92BAEMrnidsZa
pdTf5O4x3/KbUDlVw/7AglCqJgwNJeM85B+41QZ9leZZ2a/LawoOOVjfMt1vZzJ/
HrUxoFRVrF8MvWvPO8l10YkLyrRjijE8CUl26s7N/GFrxLjDTnih+CVU2FxekrsG
exqmF58m/2V0loLuzmL6B+CBTplaMzC0oaBeFyueEmmQ1TZNQtKazlyN3sVtKzuc
9ZgGpjSvnqn/+il99ZsM2sAP/Gd4rdITW5jjgLC0uAyDKFLHWdelY8Ubr57DP1hD
qp5binY+qxI2TOPU9UJx0X31xCpGWR0KZL/ELXWp/gJ82rR9Q3u0lJmaXOuct/v8
bY7cZXu86CoOeZ3+DqclQu1XQOrh0PX8MYRrbgQ0am6uRn4ub83S7d5hkmrbCBUH
xAkxfYpVLw+d8aBJxRggjJfdvWL9yQ0UIyWWWZSvO+nTOX8jhVVQsm18NFInUfIe
R6sERoBzgUXwV8rw0L2x9TbVJAs9BmQhX+UYqDHL6pllWo/jM2HuYXAmc6Y+27GI
lhFmZk9lnWhpcQRmIShH9IOS0bFFU5FvR8N3gdiB9wbINKzBMhLljISl5RWakkC0
ePYL5NDeisev4f9aUD1fvys/5Y4YPHTcAOJ9h7G/bNx/iiV8GYesm/XxDfghTTZJ
VJUO/gIbzQbNWLeEydX1GJjPPHQMIpCi14K6XFZCJZsQBGbJWM7XtFIlD2ktmYOT
0ojho2OxsGNQkmcQUDMYV3fHr1EQzTZIoqBNG3je0y2oXV1cDyQktHp6cpcvrcaZ
+gAK1KxHRj9TZ5zdE/v9+FTzKKWbnM6Lh0dZEvXUFFCLZM4dri6N4P5Hs3RrD13o
lq0RJnHaKQQ5vyqmsTWVd05+tC6OSEzWY8VwAnvHQWt/JpA7/hTndB/ASy5Uj3rI
aJSSxz3Pre9IfOu77UXYDUgcjcF1BfDNilbxArZ5OMP5DacB9R6w5hDTLw+MG+dB
b1um37E0O5Fu9H88AkkAH77WljegE7gK6+xYW6Kr4HkCva3FzVaBo1Sj62FhsSuj
G6RObEZ/nbFcZ9p6bj+wVHgEWy4HaRM3iobbkGVQF9DkIGm6RPZrqVQiN2DX63uv
axn+4X7pv1ZrQQU1b2KkTStQTy/F+8Iet8c5thPwJg+j9zD6dU7XUR/QIHtXk8IK
eOxWiSgFtszGMXBnt4KAuLFPWMZVR3rv6TnN0BjdC6dSFy9+kPrPCvqkskS706TH
ZR1h6aurgQNUK4JauMduMBVrOIIJGJ+TAFqY5SJs6CN6+L3jK8ieAeO2gDkYEZyo
OWRE3ao14UAWUOH7T4y5bYCF7oqXFWMK/xQbgfHz1p5MideWEeuy/SEzpPg46B4I
So7pW7Bvz/FdAp1LBwDVS1zc09jxdtVM2w8z3suri6abw64e8JylpYZYlnuPcXj3
KaUddKMsK5RI/UrQcVjJs+UvOk+1ELbNYcB7ApZclQouHEbDbYLKBq1UqM5S2oN1
JbLrikUpjIWNMpd/ePQ5/il1HHg4bJ2PYxvlWdk/lyaK+igrTValMBOXFx/7CXSS
N5t/2jsBEnLGjTwFNGN509PORQzBMuheIZ/Vg/XkzhRCyILWfBgxP5ZnBQXvSq0y
tKPNHaegY3UBipVp9LJK7I791/+bAAZqLi6hkfzcQK3pA5IuLiDoqMi7frl4YjQ2
zF1dwhJfHhkNnFdcs+C6YyQGTZz41ytcBf3hHQaxBzQBTw/S+9h3WwZUevIkP+Ua
8/TmFPitFYpAAtUU/MqzKaaUlCLGEeIQrz5nDvgh53rBdZ7rktNzmwzhq6DO3F/M
DZ13HudxXWeqUd6HNZa0/L8g3MDEpto410wI/Gzu7uiW7iqMIoYaUxSY3c+IfzxA
PSSCUq+Dy6sfYDFOMR1cVOpZ8GK/2192S0Esjp2BEQfptGrMxMCuHpCmh24UN8UM
BPuzyG+qnYiyLGYLQHgoa10oEXCw0V/M4XA5LTbg15t3PApHXEPazMqwjXAWjAyI
WrUnK35tUC9P6vHwwBBBzSaMq8mg73BrTeYJ5HTrl8ETgib3Dynwzm9TmFw4hx3P
P0bXNGtnNGdiXzWOnGLnQXczWKHVUwDKPffO0nx09RrEI5u60RZj69VobKx68r81
GFB4LiqyLl1UOYJIPxtAFZbaEXlqj2bryePTmBknKtD5MS2/VaqDXInXFwNwyb1S
tWa/pV+/BE/JLNEzG9QSRMWYazzqUFzqmHwUbmBKmUjo55RgAYVrU5UoBg8IQ0kw
kOyshDOVEty97dYl5XITUeAWjbCp8m5lFpDiVy0jRRqZ+ZYNhHE5Db7YsY1el/bY
XSvvUFQegmNKeXL0djlST6Ebjh1VQc6VDqKdlAwC+shIQTv9y2MDzzaLGe1Yhi4p
17+aaNT5t01uxIRiMYHJh2/zgPSNoo4JoOYu8uEV4dIYanDd/JTG26Ia6SfuXNJX
kRKL4iSniVAn+lSY01UFXOLPtEwCKw4gaj29JIklMab/aaDcTuqoHHcqIfxUQTdz
+165Imj3iZuG5XP6TlsI48jhg/FfrF9Ebl6Ac0w561QKksUaNpBXogsQTIURUhJh
l7iVvkvskIoTTvfyJw+VUf9N0pOEsKuhr/AUz7hNNQIxD7S6ooBN7uLuSplblh1B
0ZWYaWSPEfB82S8spWO7BewW1SnLMC11cDYGmBQ3e6IFAgWo8ISyW2xEo8HoR7Rz
MUMQFrzUa8zLB+6ushwIlHAv6VG2axZ/C4cbPvysHdQCJiFg87d0MLhocJeP8pHF
eZFvk/BWHt+z+IWGgyQKzj7t1Z0hILm+ucXpOinQG67GrjekuD24dqDu2rdDKfG9
8dsPYeEO4OuHLouW51rCw9sgLL2R0OecYTYGv8vvXRSngrMxA+ChRgRzIlw5LcT5
Wv7xcuwQAC2qKk4DsvGLjaskm9qiz1Oz0LfIfPBqA/QEGqwsS145HLMB2Wj+2vpe
f9vfITWKp8wDeClivjTb+bX2xunsDrVXacih8o1MEeEon7rUdngt5PXrwxZ1G1yj
zmwzcIpURnqWSzO/3C9tZj1CchDekThNlNLTOsk418jKzIAn5o0dZX5hWd/gkPR/
5ABBfpVbo7uY9uEw0jUMB7trD5L8iyKBMN1OqYF/BLrt0IwUBtDYxLJanjIOX1it
e0UeVDzGY0YKkSw0O0Ro7ckUw6Wpf2gZobEe/5PguQLKkIomo6zhxu14YHllMW1w
Qdd6WKz2pQHChEobW9SnvyqZW2HdjZySk7t3anN54zSKPR5NMJoUK8ohvbM1No4f
u+LX+D796no9VbIdKIlySCl1QbeMFxiFvQxZKCEPKlLiuaSEmmpofJs9I7XFaqg4
PDw2Z6qqrMm9uwrfBkBEbLaTD9iCdtCu6e42RkftojUg2ESgvhcqDEruMKzaR/fr
g1Lwk8O6LoPOVMKxE4S36X7+xTjNdNqH8mjVY1H+rTnziqWMuEh9U3Q7ytyTk5Xq
IoYNm5XvxDLEYgZCNuoDzRl0uuALnrla38q7gvY6YwN/LujAdEfZtXLUpE3E0sjH
ZR94Kjj3LXDfeIYibtNT/xw67llFXeMMli+0M2hnGg9ZzckREP5LfiHaZifSii/s
Gg4VTZwvGb7H+mPEunOFNEXDntz/yehBmxgN3btI3LiL6NcgesB4d/Ey/pf1n9H9
bcdv7txRTh0VjqiggKfaCY8KnPLmR2bDdTKuSO1IiQsEuMfcx2+891w/Z7s2i69s
bGpdLoxBxNdzdgr3q5LDdSrORg5TCO3GvmK/Pjq/adsJETTWfWVmV1TYeeeE+9hr
MGAz4XlNTTRPmfwCvU7hVrJfTP5erX97DSyFrrCg9xHBmiLcVrJ/O1q+nWQCfBjq
6BBJ7uAK24qvYLxlpi0HdcVG7ttmw9fURENoQIS9Bynr0JYdY92Ft/+B7/GD7hUQ
OHwkSh6JKd/9kcuu30YJwNvihNwbsUzLZrCXgoPT8J+PsJT1xb5/hZmoZTb7egCs
Gllb6YjfXyZ7ulwJ+0T5YuxtrNITtmiMZ4OE5iyP1te1PH4y2AJh9+0kpDDZkfxA
9oeKzUW2q4KoR5eWIHSkgvKCtBFNYTK6d3H8RLKkIdSuZEXjBZGPQa30G1ii12LJ
Ima5Aj6VSx6RmhqGoIz6C/A0TitT6DRy9Mt5tPVj9hm215khy6XTeR4vRf5yukuG
L42Sw/F38liPAMe9KK1f1OsOn86mTVe3GQzEUYz14b55k7blxWBDMYiLtXvRjcxi
jj4fzTKtYIRCdmeU9M/pMrTfyhqOJEmuiSYjFlPD2W3/fELXVy68SgDMZICqegvz
dvITwRrCurRfQf4xOyQLWp+LIoYkLt7Q2+ffLI8lXjefIhTzqdEHM7U+RS6TzcjK
nNsl560TZG9WTJujdmVGiYy1dxU18ZEigMEWbgrjHPNN48SpLbWT5LmxCmtAeyOW
ZsHisRyuJn3Jb4Fjw52cO11hmHH2NOGRce1rxfYHwT7OiG5mjreAwzy/CyUR42b8
GIDqUI0otxwJsFa0DUzsJvlepaJyWebBZcc3GLr2Qq4715xK4hgE+036xSfHVXa6
y9P2w2nV7VYRp0hqJ730GhnbI2eMnHJT4tDgOJTHKD9vOjyEAY7wnyjUmFChbP6d
re4ho+BVnUxaUEoLkONOXA2LNQRAQ08+Q34KiMpi80DdJfgRNkDZtgHFMb8zZ5SX
H/AlylBHQA9HvbpJKR1Z+oU1V1+vrJlEwWdUR01t8ZHmTHhFvRkYcA2GWgBVz0Fe
xGJc6+6yaCWr3iu7eeNZviDCPv18E8gT3y8PcjXr0LB8QdoLkjEZ6QK8OZYHTzTs
ly3gUIHZBH5k9+m7+TfA5cSy9JRp3+gWau1acKpqcnm4l8v0lKO9dUPbvtSwcinf
0cBq+rN6FAShtKJ6YpTDF09MoFmxyo2rGv7UH15nj1bDbTm25NcwmMJtBaH4k77i
O4UE/TRoW8Dv/73/sXVywzzKJxCoh3GXsrfcyaZZ9UTsPkhC2CNLti0E1LwxIVQT
W/7XNhrN7hNhvyqoTpo3YJTEaiuvLvxSZ75Lmau9TNLz0sVawQsyGsJ4EuAkCVCH
OnN0oz/8RgV1MD40LLDTB5ygvzkBbPXOekBg/v5IqOXqYn+laxffE93bwcsY8Y9k
bwpntu2Yahe3EMYJlT4Qvb8slgcSmeA2Z/eaubCg4UgnzwCiuyuXACLuUe9Q3yde
YHi8ZA+Mc/w3nT0mxVYSfq7nGUndlnUvIQiyncMLq7lWWmm1AVljSMGPoT6x9PQR
CSXkyzn6Y43BP2POtgqyROltGxfIWiBfwO/Xv5ZGVgFhsPTHlB3g0vyx5AU28aZt
9Qlybd68S1Lz6sxGdJZKM2HORrupANaSKmdy/M0Mo2w1RicxQiZp8GRSqBV5lXoz
TjgHpjLNnT4mevexWZfk6NUUNrxp259jyin8Gua1bS2TtEV1QpqbBUg1tNKQ6SnN
jdZr9rM+XExTLojiK1ug49ogzwgsmGgnEl60lfMiTvKNPT75O+1P7VICz+niiZ28
wG6LNgB3Dz+R2qWTlJxU9AEM1kDFkmgTTZyJNvUqO8Tvdid21Fqr69cWS3fCs6xZ
xpe/LUz8nkUTwjyE/Mnu85dCuY0ilfBSm6mYJtMtUroNfTO83gDHpZyNE6YVwXqF
hNv0THRX8ec4j4/VBAlv0tNdPHoOQ9yRT0ahJFtsJkSLiLlmaK3exHbqsyv8cw6S
ARo87a3or/CdRFlzElwqDAn4OJF1HjQm1XmJ39Ilq+hmb0ee4pV1xyJ+scbOBEXt
uwRO2b1wopjeTIKp8vexVRLH1Vs93Vh4t2SssEvPi6nXCfb3Abt4c2Ro7zmCqyOG
lpq1uE5sgvEqgSTvmbU+BGQ0eGdhLSIz9d2aUOO42paV1TiAg7lxK6HodewGRS8d
T9O7TdVW4ELHEfMEjt620QVs4O/ZSAWeWhfKDn6c4o8hDJWn3wLGaNVB6rt7u8om
rjx8Qi5SymVHjVjLp2Dw+7tXPkgiad+OYeKG39B2ZS5XlegQ7dGY+jRHdhra6deL
YFP1l8dYw2qtsUv1j4avz4J6wMZcqUqDMAisG/bpPVF1Ex2CMwpG4GKyCDFQkgCJ
EKEcmO2zw+tO1q2B83Yjpov8rxUc5ypDj1sYDz3UUASI8+wOVY+id/2a68ZD38FG
l3pTm8yacqLaU0mnh6BIETeoflaL/nOBhxTwDwxZ6vBfj1+Z1QskawFwGfOU4BCi
HPq6p3e8DsUs+44qBV+PwbDq4WUhKhZL6bKoSwCnbadzh7/WtcfV0P8VwseVy3Za
kwTuf5jUooaEuBtyUUQJVIfx1/DDizA93CC8T+3qWcn7pgwG/exHKjzwiTEISaBR
DgNxOViRyag8hUY9AmY9Y8mvIg/YUNsbMZUnMjp4XEOVWislnQhCJK2tWr/hsCDG
0M1QIdXMep+cIZ8I/3yiblEWb8wje5tZOTEN13Io3B/ShIKsoZJaNmeX3ZLVBFDD
KpcgqO8zgWNi9BqrLjRXsYP6p+LULfZ2mKDoQzrxXQoIU4D29RaMj23baa3fAqPX
KVHXOMKYFd2TGaxRztSa7W6zqtaFpVgyllrHk6+Dc6AA6FLO7Z3hi7now/m3y8Mx
d0mZZytFgGUDIK1Op+QJJvKfqubenhQlijJwNs3haDoraeu8dLSpL2Qul+UBSSrj
kw9U/iazxK4dKB6hGgEzbQrPCpaXeSlDjdojp5AcAGq4KSAO3AzOkHEPMGhLdr+f
osD629aua0k1TE2qEtwTBJ0SpQd1bJ3mNH2ZHigg0h+Q53QNQg+0+HrSCa/Ey2gk
NR5yyDQK3X4EmpsxHfxv3jm4OFehb9zEzdYL2aHyYe4jtGxwivuv4oNSlRgW96Z7
RTTEn8/TbxJMsjczowWqadxYfWrWDHQ9rvn9EAvBPJMBP64NEBL5KvyONlsSyB3E
PoweVB2X+5/RI3kclbX5SXS+MqlSWT1EyFwbDreZSM0s/jBLpdtWsfQNznqx5enK
yAUCNHC+p8BFcuD/Ct1wCHuyH607zChq0glOQmcKOdHLAnbdMHHZ6aoD6YonIfHg
7/b/IV1dWsF+bZ/PRjxGxY2lb6A0KJmfwuqfMbFynpFeq6VrLefa7CxBkQrRQQJi
uZ36+ZC1IyR+myjfODDCWamA92/g6wwzmAYMkUz7p2O8Fo6s6Epgw4ILD8+qmfFT
uO6ZtMWXZ67r/ccAjvCPtl7X5iwd7f/VkkpThETOHHlTjBZhgH0BO8YHgYMoDTUF
o6UHqPctVeCIViKm1Q3+Ynnsvhxu18jzOIX8qTKxBv7vdQ180LejLTIJXMWM3gO5
0WBz6hHn/Gy4al0m8xExOm1diw3nTx6b6vi815levryfAYTftnJBe3vKPnlAUbrU
dcV9Cnvqo1q8F8Xj8w5s9gZXOEJM0kNv61MwaX2JMhom3jeQd4mA5tPx+hjE6NY7
Rigsl3XYNpE7MYNYN4E1Yp+F9ZaQLSTlL5pP6FJL9EZoG1Bv4BV5Pgzru9emCij9
xi+4QRfpa2VFbLC4cSKfWlZTJzQsTBIDUzxyyOHeYXId7C2ZOcAIx9KY4wjNNoy4
zgm7sFACjp/ICJUXtLZ1xR3d1o0Dy3p7myU5maKwKdzr1J/LDdOo6msjshjl7wc2
iktO8/qNW2S26ldYc1XaV/MWI0hNL9lg1BjbqaXUKN4jG1QCAzMO1PzHV0+bOzEm
vSUCm0n4ff9q1Ei0LLJC4k78qqYEyR+fWWSMlE+jiN4MI9uhuMpMm8TIvWrnggm7
nlQrY/ALtYElhRjU+eLJUU5Mk7NiqTBuL86c5bqTVDzVzJcyziFGoBZTVhXYG7cN
XyQm9C+NxTBOFBLm2lWexc+t2oagvliMj3HqG23DEgnjPs0pY9p1YILvlPavVNW5
ssN8o2MR+ux4U/DVGK3QUfGjHjHm4TjwSbDMaqfUBWiZwTxdav4WcRiaDOBs+ILo
pv+oie39q6PTxmeHTyTZ149oi7mptLt+H0UwwqByrj/NlaiQ+DlGuFC5Nizl2oxE
Yf4zjWJwHnLO0UbLMf3PG6nzkczFf9HCK5ov9JEHxJ1wDQO+lKfmklSZvyE/bnD/
afiAn8TsPCWY3rTglhnhINLkVt0bFnA1YNuaPQUN6JroxtYxT/gLoo15KH1QjXbW
3d3K6V0mCaW1TVakeURzkOTIEs8ISmPFuyZtncQsjyy+V/dAO2fRt1aWWs62Mno4
MaIK1fUsUu3ZWkV3Ho8Vfh7HeyFNRn0VoKPmHxfvvVLg+F/t226neqx7qnrpgzQ5
b/73/R44d2JGVqqa3gSk5hGYPUvl3ovNAzMiETQKoyPBoqbMA1xGzm6pGHlBtbB9
Mb1Btfgg+Nsu2McUl9uIWAaBN/TsLgKrGMi6cqB6mvrpfCIYlV7jesPDFufy9m5e
oj64oZ7/22jr1yTDM+b22IZiezeGdjo+llw9kjL8ZHwuYV6DAmgD1LJ/30OWodhs
4xw3nC5LQPcHZ59Opld4YbptlJ4/UIluaVT13XzstCvXdgeRwh9jHZL09ldO4k77
mSQ0Q05E1DqoX020egOfBdPEJniCJJghJBeTlzqXhP3x/WYc0fQQroAyRSBJ6dXh
qSBr04oNnUtANhx/IYcoQq/f9XHGdva60u1oUh3XTzjaty335GChqKLlczZ1PbAT
90F/CNbT4acSEmEuLKTrbeLgKtJWrvtYYTnSHSoWCwrQT8S3FzzQc+/zEkZC/lRs
cgh6VrCXkVBwhUG0LJPLlAxp+32p4zxoffySJUlhJZOSp1qF/ftfngYQNiY5+y9n
qF2bakEz2WkDt6miqFVB0csbOr/09skXoeq5zG/Vpimmh3ZdvTKyRlnZlH1k3ag3
RHUSD7CN96lpeTZygvUVdhgdM1S9vmbodsy8UzLY2gjf2bQdmn7u57KWM7/4AHNc
47x0R9RmuExc/ZI5GA78X1wlCsC0rOd6DhHll4smeF9/kdBp9xqti5mkccChdki9
U5IFOQvcQH0DzQGf62gb6mqv8nbeQL+vpFdFpn+CkyRMPK8RifOEn+hhsgm5zdoL
nsD3l5rLJL90/fQi7rP2YJcumLuBM90PGOiqMfQcqt/62XrmBqmhYL+ErF7zEFFn
3GETulMGncfDjWxxQTZuUa3itn3ATTZ9CKLWJeO9t5esVphJCY+jTB8koRjbivz1
Yc4JCORwnp45RJ458FLb9h3IgPY3dj3oygxq501hjrOHqGNswiIsFBtGoLBqnJFg
zEEWYJIOihzHwztH8OGjkFCsZCzYdKqxO+6l/eJcLoaKGqc1fNq7exZGoamBmPKr
SEFnn2nTsFP7r+IVYlgnXvR4kTY8jla9ubTlK8YdpAG6NyYuMEhycIGmEZzyakr1
RZAjOpgQhTxkhN9mlIbsYZpYAeoaj6DM8r6A+k0vAQbQE8MVinycsKp85sRGnsKH
6kbt3OUshg6KrXDL+app5X+k9/clm2N6evwb0gZOR20ujKn9GWD3Ch+1HPyzorCt
/q/F+MdvZHRNkuaP36+0uyXetjt6FLf91oXduhnTPxzcdB0fjX3sjil7OkknrHJ9
zyCvwTDocHxrKY6BIGshpb9d9z0M2QbR+0k3ES1KmgTEamtjIpyaP7iQPaNP7AQD
SrfPKyQNWsLXAJhZD5SMZbECr25tgsyzm9lLh2Feim2oJJICbAm5TkK5n59GFgxf
7Zmbs4mg1PhhUwxyDI6TkZmhf7F1zWVsuDVd2QGwLgPOiVmLzcuvgft2WH4F7az4
c7WPBfrxvvXf9gWrldP9SLAmj4dm10uXHCMx+3JJhhH/UUtK9IHdjyyQS8VBmnj2
efH+qVdXzgMhcKwwZJjPb3srS3DtWm0S54i6Ec6xaz4w3ZQb8qBKOQGSbRr32oZK
vUfMdDQs6M3PFBEgerLsO2uRcxgy66UtmCauhbUsPNcKNFWewaFg54GBcdBYOOZA
aXYLiWO3LkeCmjHGKb+YpwqUYfgD3Yq6cLJSu5LpnfTddhc2IN38xGSDQWSwwe1+
aPt1nuQ9vUK1GRBAJnV9DNYF48PzOHGmBqhaFpa15+YfWG1NRGyphBjsG+jkDxRx
MxGB/71JzYSDAHKkfhImBy7Z4tt5aAITivkvvrL6/127L5zh+R83nzWSGacuOoaH
fjdltLqN3vh75HzpFuDtOQgIqmZvsa+n1JX1rpqSOYUQutjPtBIXY+nsYMfdKk9b
qYfWccnUOHD+lsID94E0VGGR8lL55fe9a0IJpJV4K1/Hat/SLWMg0s9ALeC/40ZV
zh/pVy1Ykt8GcZSk6TxaOlLFSzRysbx4SYBdnJs/jYIGbvk0qzG5OXnK+MbBJp5X
OUe671obmOFGar8DhGNNYwGCGMKhxTyiV2rS5pQYIuPPB/BfDWmM0BUf8VdbVumr
9eJwdjxsG1OziDPHpklEjzbK7CQT5wx8l6Xkw9kk5m9L8R/28XVZvG92sUPni6ye
hKLFgPUd6csMU84ZeWKAMbnsUSEicCxL0NsIUAk6yY9N/JWTzPwFmZKAFxHZiDDM
dRfvZjaekaRGqUBm59IxfNbDJEkV6xrguBMCpvvwdJIY99Ps12UOegOuopyFXnvc
h64KzCoIkZ6CLtBp5MvnMuH84nGSv1Hx78Ly6B1x3dSTp5w/shBQvN9VVTZon3vc
RZ8pYGWgvJPtZKdVUGbwJH59AumwFb0+WThjHj2PY/v2FVGuTGRI17SugqJiRxYy
DK8A+nMYV9vayIyiLXuclAAUZQgtsvwmjPDlW8JFKDDnUSkM5HtkhJPaoZAehusJ
7O1WYBDDuLR0iqdakKFEd9Fo8B/mpbzQUyLhVzqREEi8PoUApX0TV7DgQGPzFTrv
hvYWxoJrEDC4SnV3G1i89ruYKjqXAjSg/b+fnznOmfWERLVQN1x5IgGH0KOPJQma
LICPPfrC9ZlMTs/judf7vhEeDa7oXivqoM3+i856CEq2wylLq7zrryz1/zkua9PD
L0d1+/uiUugZZr9e6ze9vg405Ujz7M5GetwpWoIDveSFH5j72ykLkdDSmsxShSNz
My4JrFx71RHYp63C/rBRhWG7DUcGosCaDZsugB1k/wFOcaSkDsVZ1I9Cxpc1FnEP
Rm6+NSGoL8B5Z+33iHnhNv2DZprw+aAPTF3wOKmAG+xbTrFV32jS6k60LGHNzZqv
RMpjx6YX/YBGx78OL0OprB+5BW5IpzB+T4QxvT6uDdvMpxGHL+nowjuVmMnct3V0
XPSnmUpQwqAr9IupBFqH+0NsIR6H0NN4cn1QoN52Jh3OQb0kTpuqtN5bhe69Gjhb
4uPD1JheNqeBjdDknqMN0jHOKVV7/2BLF7xg/72gFjJWXgrW6kIjpDx3/eAobZ7j
WaTJG9KrSn+VoV2n4tNMBUSYWlRssc4hrmIRrrhL7YVi1rZlZWywaOp0r5NIM4n2
m9qM1jeJNRP39pI9K0PpE7SwzQGX1MrIWRU7IvbaibpSciUnlqnpbuxinIR7GHAB
f/N+49vzPNWLtDzDU/sXFwTf2FCe4VdWuNgg7HhYDAZz2Ix28Spj2uQFA4gi5Me/
vQaEcI2KOHH7K5AwhrqVs3hGLqG4Tijz30EOef6vIrQ8bRsxX04lHXwJEau2Uwhr
CpxkbrhUvhuA/0c/XmoZqlvXC/6DLqtDRCI8wXr1BlH9IA7BVlMu3vSKTKYbBivT
eI/9oVfd3OarQKHWmObrEdvB9aYbMfhXB6hWjZEGID+LL9FlExBNRIp5CYTT5wwO
esthR6hB+dG/W86iqxfAqLhByUFnZ5VGDvWItCgEkgYY8dpcfGv5PEqTsBCJozWk
Jn2sEoXwt1JD6sqPS4Tdd/a5PKorT6RXve/IHZy7nIU0bJMJ8TMrmnxKEyWZCuO7
P4aGBaFynWZZIRFdMgUmonXgPRTHibH3ebPCbpzDd5KpdlTFdEqFYZn5CrHtygT7
yFrAnjya1JfoXBanjWcdGKLcgVAlvCI+nJPnxw7IK11BDN8engvFGZbKs8otgKju
WwUUp3iolrcCDn/Xs7J96IaEwrnFO1Bd3jX7UaDSlzqOxjQOAyppcAw3t3ih5SEo
2/muE8/+GEKOGuUKhkQq4/f/74DOC0cyQ3J2Zbe/+nOLb4OwnGtcopdT8RNJjTbJ
/2CqcOlm17Yxd+wQyfUICciQquyRlrEv0qAdkdzHXXBnOHtZMsETEqiTi0odtnnm
jk34f4QGH0bizC/c64B8ZE+GVQSkoNTxYHk6l4MxzjfM7V3KYbPaLp2sVpvFg7HN
q/4ivkaQztKhXq1/YUi5YcupkkSR8dMP/zHLgCREzKI/e+Xa0Xzy6Q6ZakGxQ4F7
HWIm6XaJQkDSRG20mwYCfOLRR3frEJ2a0GDwmWuf61KaftGX0Q/V5UUGQGoJ37Cj
DOl5X5HakPo0JiFOAtd1fA6y0xEEYANEPRIem3F+ZonitqgljEiBVtvdH90drUzh
JA20nIKHN7Ti4TpDaTT0tWHJgG4eObpHwKgOgXvURZnmXxAcSniSX8G4I9D/kwXu
iAHAmh+KaZoS/Jty4LohkmP6yay4ZDLFbpZD5NyOBvRoDXpwnRmuovUJm0CyfbNK
LssBjWAjPmSosFJ4cKKuO/rl8Dv0KWMDvJmdY1wHBtu7VYNTyfCN6v1zUgqkzD7Q
5eFM2mBjR476fNEVp9Yb8m0KhSoeGLE6m48/6A4OmP3dJWiRq3y++0TIWCBMeuii
Bdhjb/qgWIechqN8nIWSa7xec7wZ5rM3B0smLZA3OyN2Hbg+dOKGOHsYKq76h8cM
+2TKlDp+XaTVAqkDzMBvdOz/6WEm8Uw7UiJe8oDTZ9p80YexVdVb2ShvTKq30iBE
QWhG4aBjF0OgWOBAVfNB9n9eFcVsAxi3IEMu1I4qao9engAAWIS3BYzseB5D42s1
vBHnVAZHjvWIs/sexxyBMryJQ1Zuh52847rmNHgeV7la/XLW855VwzQlJY7xFS1Z
+y2i/8DWkdzS93fS5uYyLIoelzlduVlGeDGqHW6jLikwrlLlIJ34LPXLVXf98lOy
YQGA1T/uH4SS/uOG+ttrCuIbDS/Imvg821Xbz6NIHhg0Zu0je2oPWidt2IvGiks0
thGNvQ0g2d8ot1ZUS+VFgdh+F/F9QP2HzsDkbRPK/+fkb2b3sVTEAyjsd4aBbxWi
rUXOaMDdr4F0ZdUeFV3A8VztW+UQjy8uxxOfhex4OJMP01pBX/xTzcnm3MPwJNjQ
eNirnqexlDJdSsLt3Jxz3itwF+Z0ffR3YMm1L/UzE3AWEz2muH4kmQ/gekPFr19S
YzQkji0nOUPxhvZyfhIdz1DVmXn8HPyr0ps1WNOkOhjNwmgOS0fKfiDBz10ReLhl
nf0lVQ+uH/l4qhgORSWiNp1+u1IskBs3zdTMZcqIYArcfWq/Wj1U22fKcRsoCi+1
jL8mJiAW/QEZR1FA1f1a4V/jo4oHtPCpGdtQLmAnH9eGubJaDEJSON4YMo+xnaP1
3fASwRWqzPjhVUYNxt27dBb9APEEI+nHlyzjZJ4U4MP3UGQo92hcHFx1aJWF7At0
W9Wjc9WTerbNqjmizzhb4QG5X7O6iDYxy2OIFy0R4XY1NpdA+8abNL0D/dZkO+WR
MDhVkDL20hsG+03WmYMIP/KrodtY0Zqtc2Y3i/Zk0pz1fzjIOlPfXNnZb8NIMIfw
+WXf3t7VpGtUikwAjDIWxriHM99TlupFqHUJVv5w7OOwPVsvF+ajHHcU8tsILVYA
hQrlejmh+AvU0Kp3jOSBpAoFK9ktVdU0FDoOCiEvwzM1h2vbmYHZZSl6/ErG4ilB
zIjpKjkpcjQJe+8mReoMNfK0QtdTp4sbBkVdJfyEvl+0rA063J+HVxBE+feTmih5
AAz15psKRYx89+8XhNdEc8BACx8llWXoG8iqZa5c5Wrx+44qmOI/JSnsIi7jdeya
csMiLFO+IBpR290USLvw5yHBManjQE4+yotoIdiS+fltnbiykpPM9xacEzwJcPia
++a8BX/O5/cZI6i3iDwaV3vJFP2JV0MRH/J6w9G5RAT8rBqNB1W051+ttdm2UkTn
3BEHx1+tcpiORAxouh6W2ruuX/qUgk+6zMwcsPu/5c+OEmJyLZky9lmOJa8wrPdH
zpkmh41KBGh3X5MQVxIae75sg6pKnsQDWMEZeEZjdmlOrZZ9gNCHqvM5F+W242Zq
dehuWyWmEJRTY2zFWDd/SdXKEiLemGOyNudX7I+dyy8pRwWYfPdsWKKJmz4vFyHY
i2CmlbXofeZ2s2v75N4ri2bwaMpBf6YbXAswXKrK0fJ578BHebsjHXgEYWrMJKVO
I4xG0NYM6s5q1VSE0CFLkXz/aekSBur7Eg71iSTQg7jGKN737oIRsYDTkR3Noi5s
TkgNaxQAQwKQ7bWx1AFqXLTNAMWKlCoeP72OJvR8PyweYVw1/fhMm20PpnimSfdT
Wkh4RBKDht54Nk+yfAXQswJe6T/k1a8REGZZXEXY9/XrO5j1JQkjg5sASWnLXCOC
/1mfcnDZ1zqgT0hd7ZM3uNcM4cY0I39oBL2YnPybCmK4lWqLUCL57pZ+/+N2P8Zc
iCtZoauntzQFtpYThvB7IIObUQqO2kN3wBvQn9j26/FT7UWWKc43Lt7mHffcXyyc
sQ4aQsS2GAwDfqM7mh0Y4S2CKvfJVTVmSnMPAdJhbwB9MVmXWzqj9/4sLJS3UT5S
HZPBpv2zJ+Rwicm+2gueSDpZLy7h7J35BOciSJHB1qMKDVqNIpzU2D7O+1In2L4q
oa4J9LNSsa8He0Mo3kwTPIr7j3xvSwBOY6/pGKJ4v8BdVBoGi+h/UEyvVQRsIMNi
d9oF/PC3m16S+z6H4Ce9Zp4POjgmK6nRFOq0YM+fbG0sBczY2L75fD4UrFxT4Nsu
dJFBr/CQS9v6baj3iA/4SGIoik3InY/Ubeu9xg/MxLvA1lRMgsCJ3TFA8PmJsXW1
RSci187+Cx8TEvFRXCLozrCFeWs81SYFrehd8kMBzfTviw5HBE6GBW49wLb6Gwhz
USeri6N2rzdPpEGGA1PirwfrhvuuKCjL8+dFLo0LiNUHgGOIgt1GAlfR9Zp/sZr6
oXGBJkoSaFEmX4eZ3f4JcS6qOV1UvCeVgjzXCNLG4+tSbY2crWiqJOJrF+i037ms
drnc0+oJmZQBrfWVhB5FnyvES8PtWDSG0uLW+A62JqLaU+PxEhpGfKGbS7e7KjZ0
yBQJTrZyIqJzpL6m8SgpR7VVOHVk6J+1iTD8/mw7/whgErrFSTWVa57Ro36wj3oQ
Wv/i4tfRbvwypsscpF0/XC0AGZFb27UPKhuGs70pkxDN+V4jJC8YP9urPDsi5TW2
ruMBXFLsGJXrbgq20+Taotd4vox/wvPJNYrFj8H6w4WyeRrpsVe7A1W5DJqBCUP3
7alFHc76LmskhcM2B0bGolKHGWD3mnEMWHbh4e8ZhiqCBNqJ4K/k2A6cL3mQd50a
5w8LOV16PH8ymVUUhXoGQZUkWo30Q5oZWyRmJr0ARqML5fOD19w9WdkWAMfDuPzc
OIxmmk2ORRpL/2yikGTw+HrjG0Ht+dO7KM2UURgOPB2f/KC7k6qOCxRpgc5L6Xsp
HdwU/pa/Q3XVuMYDnirliGHcfKNN+hZH/lueUT02X9jlqbLWAtRN8sOUay0X9bRe
SUOFjGu5kIuhdMh4sx3PCd70334jv1OK+tH10UNwaRqBCoHzfhHi4FfX/yYvTw8+
zBQjkUqfrBsvwRu223m5AbAjE+dstmTBKGlFYreDpWsVYkIz5382+ShNxDx+apKv
MOGrvABteI+w7OzJ2C1jO/UiUSVuGR2xEZwmtz3yVEO9MB4MM8b/gtO4a9+6nzr1
A8fzveFK4V9TAy4hhzv6/iOvYbiKjC1JnYHjj+1SzIgJ9QI+V3q2wYiaPzwsB25l
CF/JhancoKm/2eUFhD21ybayewT7+WLZfRlaRwvj8VvkBswrfXrAUcgAuwan82Rn
aPCUa5CN2wgPfuEc/6Nlx7hxPPRtJIO4MZnCWkaH5iWYSL2R5Sn1baG8avIbtBNA
uE8Wqwtihe0wMv7dDxhSMKwwEaEQpIob+2qwTfOh5wppzqgMvbdkq4uQHWp9BMiG
IJDHW7fJVXfjGf/ZS1jwswN7nZzPZ6HZReB3YuS6wIzSZUfYBWNVSF4LWGf2FLGb
M1uqOUv3MmrvUOJW6L3DbGU4EjGe+p5rvSBD79gIKXxcJXx72+MIKoyaoppoRvO0
HfBatjvaIOFCJDcgNE7oDmm1W6sU2NA6HPmHxyn9sDfrQdWH59E64ilklWgqLJCj
MlhJA7Z4lj0W4IQPJ4SMTlmsUwWXZeNbpLbrzbPUdJwSJDIEenHcHyJYftFpmdUp
F7gXA9GWMNGNFnjY0Y4GKjGLLwXsjwBEqyqhxMOga3dkU6BiW2iitJgEtHa3nJcv
0iyB8csacYAVFEEbI5W69QI0fKiZrQ1T/llVS4CjHlhMr7myl/aOxLbgLm7vgrKQ
E0GUhMLgnHpXusfEYLBryUDV0lNmkfefWPup8nntwO80QW7CdvumTulq3M1Wkn3C
0n6X8xTsMJMdZpcAQACwfgzLQcdfhtLAFbm0ZC/arPp3I5Txjs44XrvZYCT6yMyi
6DFhFZSlFdBaZ+gnukVkgS+jIg1eIylVuNNH4qoCoWdZZ+6t8oOMNZny+gVmK4iU
BG5HKm2wffwHk3WMzk9TRm53CF6zkOhVD4UzAN5HlmN+0177ilTWEHVGKKg4ZCI8
1nKwuNHiV/VGFRl6mJUVDra9RNsuQSwPtrtki3wr+JgClKvK5JDFkjTaSlRuQgfI
lnqYSsIoKdvEXsz7o0NMRu2b0tEGgCBGG8PNX5eni4+8bfdqXhvE98Azbb70p5lj
Gq8tu39OvBX8YfxFaEYwgiYarQrVnAIfdQgBMWJuBCiqVFXQlBjjNfu1CLGgA2vM
Y7f8WBcQ2XhxnSrzopBb5baF5GWGLqSOoOlTZgrQOSE9vaKNJ3L3yuuvuNovtfOB
bLhjI9YDr16s1blFgggnFs6q2Y2eAUAgEp8xFq3/iPNGfi912pnT9dCHbyEocFXe
+1VaSyZYkiDkl0zlDrI0C3lyVkSs2meho4lUZVQX/P2QMy/BbGPMxvJicZt1g/q2
lQhH0hEKbYnu0pqb9RwwjKZsQXOhvoM9pGp9KpLTKlPMPD4j8838khF/536UtkU7
/bjc5OhYEZhrzxQ/H5czdkVI/UrZkUC0Ji3znAvmmNCXtkTV8xAeW8hMYyw20UUS
7BrAAIXpSG3C2Veukccb5O6uSaj0oeieD+N/zGHV/5E+ZNCSz86KHywyZ6hunSNb
kGpNoM2RzvPdZq/ACB6T63P5R6pt02/jLHZPc+xxigozXXQ6mqrXBUQvCMfq8//Z
WSh4BZtG2nWVkRmUpbZ9g/qWpII3nqpi5pkpBX1Izmp57292JABHi9E/KoP0PlnH
76ss81bnL3/nqIgHOPbacuebAdWn/vpgVapcH1YsD0fSQOLUOec+72bpALjJGx7z
phwbl7s6GPTOqEcsPngyn/JX7M4TkjocyIwMHv6t+skNw5nrB36zZXXCWoCdTPRU
pFhkMCDkClMbhySgGlClsB6qnhrWjDPKTBfdvqiOehu2sahhFN3vfV218A68b5e6
gEs+IL0yQNFWl+JFnUEPZwVAJ/kE/QO+EQxK++KHcNjbkzGldkZtceGbdj7awvij
ZDntb9QZNqUL/HwL5AU+UlYVLv9v1Z9aBP+hTgnTer0GNMdG2sQXruYA8Sce7U4Y
5oJe+lwSm1C0pKeBC8yk5feos6KpRH33xYggGndiKwHp3/UKr1uXRjGub2PgxTi+
/GsNUB0z4/H8/rXYQLEaREnQDgtZIxu7HmP20y7xM1xg5vA1PBKEIq8y6thq8m2L
g4uGzynlFj9JJjofYLy/nLE9Yo+2tFekgMuTW072QoHn+dj3W7NjBkivC+QnjuMx
SxQe0Rqfr5++iDCJKbIn6JVqRtQLWGGYZYByLjyLN62vY4vSAFirh6CKvz79JE3f
2ritMgAnM4rn07pMxyNX/A7TvnITD+I1lkN/N6/X5MoQJA2l0//0+LgYwB41Gg8i
cGyRIEpoY+uburPbY2eseNS/2GHCW93YjGTXsyxOFdYgG/DvRILce6SxGui6YzwJ
Yxy1XJPLZUkFT1oteuOhFL8bBFVWQTwz+8no9wf0F7oOq3YQxDcRL6Hc8A7VC0n5
6kwgvoXb2fGkuf8u0VBxU0UqxmIf03t6l1r64yQsmi3YTTSpMfMDup28VTVYBGSG
OP8oU1qHMO5yvYBckapA7LMBXsTHx+kwf6+lPe72+BaDxv/pvbzw91kFGKDMVX44
6PyhyG7xrUzwHvVliHSiQBnxidPnJ/mjCGxTjt0VRl8jxoPzJnhgPDf1FrHqfAUy
M43lv/OJBKcUFuzrdvioJIaGRZzZN27GscA3cNsrpG1aA14SUy0pcAItPruYKYRI
5HuVRoVYgk9Z/PKNCEoJ60cHfV4+sffZWzvID3zCb43VgNLsvD+a4jFdnSkY/du1
2KQsg+uNOosFCAsdGQVQ/8KppQSkX44hOooQrAI1t7TwQn+HVVlPqf0GsjjBMn7+
YoT3TucasEYR9Wy+97IgL3CdfOwfQunO/RUPw3CQHLo7IcMhL1kRZTfTWDblQUMP
yu6gZ3vAFS/mzMD3vSyZ4AWUfafXv1Z9lNXdkuEiAbGm1rVd77dwcqiqpm0S5clu
K792OC+U6GzL5suqssBmLIwXaKc4XxMDKc0O8UxIrG+i6psEKNPLWnDmzkVIpcPF
nvlxBpQx5GRO/djF/h/BgX0DE3G1SK13Y9k0QXGO58KKNd9GskTL8w6KTeRaVADm
5QM+s6SHX0xEC34by1dDLkibl0q8dXv2kWPOqjtHfOLlJSRQx89KOLsQJ+sd7NPX
k55uJMIeL0CC99n3wSKLb85xatXVvP8KWu17RQ+6CueG9pp58I58IoTnp80pMDDH
1TTwEJBGnAu6II1AOKRoEpwkrH/lGdNdY5/PBWFHhHS1X985m+t+Lwh7AzSQcIRK
iC6BvZ/6TllrU8MO20E38JFmnfAL+YArhvCS2IJwtIeyTG4KVy3I5tJ8wUXgu4p6
gpAHrXA/eJa9j/dGGNeqQoYPX1k0hZd/n/3h2+x6wvngkZUK5bVixcUOZ2cAddVh
tfBzKJsrRA4Zv/cpZz4O8wLsCsvRiZ/rLX4cwZY4i7YttyoLQYbXptLlUKtvCnfE
yNS8IgC/msB980SSGEE2CxYbMEv2pbmVSVhvAUELs5Yhpb5B+KvTrqpFl5/0z3HR
rBudQHRCBpIQxdCvYBMMpFlALvYcum+pTiWfh2cdPg/snSRcRjz9fOHcXfrWo3oi
6r3XkyD4299+CxKhmrta6QOQUCQnkXHHpy+IFp3OWK5gpCRMfIL4esLdjPlA/kx/
jIMpg/68GVgSewLG0VE3DuCZaSLFtO0GF0Anu7m9YpPgJkh282QPaHXcm0cHN2jz
pgsomrd5iR73icv6ZqjiwlWqAPnHtxC/2Rc/xkVTJoV6oe363gw/5qKhSI65ufzZ
a3uBNT8+nInAaq8lo6a8rOibyMMKxMWjLPfQFhpatyP90ELf2gp8T/EY8UYqyYNU
RlluBqa2R4wea61pp27+bwRvsOizYoeCBKvb9HerAUJHGzqowFIc9QNRB55X07Rt
k71PyfqrjQzN5owwVt4shmD+RyJ3tFL+KfWiEyAM10q3+UNbFO5kBPp40CESBRsw
muepfvscmC2QkZ2FbpWdwGZdDVdp4sXaKHVkBpOhPy6epTpAqDUpe38xa/X5iBMh
J7b983VvaOk5AI5mVWETRiHza1w4S6MDIdFd6vFJjcKTbQaK87mkaYyW1Zut5Gn2
+YF1uIUUbqaJNrgHlNFyg9SOVqd9oscq0YI5x62hc/T0MhaQAB1efUyenJC/JyuF
bINbjL7xKVL7+OTTjw7HsWjo3o6DuTq16z1dWCKs5U/MQYZxqz4H+68pVHqHPu9l
8fJ4kOhFjBipuVj/XsIPXwpHm4B23vPpVn0DXJuMLL6pFpO9XSgprYZ42Q1C30N8
+9K27DSqZ44qV5s3XLvVTIfDf9P5VH2OSQe8SLmpT8tLRbjKUDtvVzCl4xMIK5eF
a5isThUEhokwuARLzBqdXApAaIOn04l39psWryqjL3iB0P7/fjM1yABIQKZFXiWN
jXClUo+Lgds0JXZd77DadTxa5l+c81aU1kJUecjgk8fQKItGuwmUU3moqzNkIBRe
ysU+YbNWQWfxXAQDnT5yOt+DwqnMsogu9w69UYUaYkkBnZblLvkM+JbNGQty2eY+
n9hlF2p/4doW+ud6sc/3BDwnppKT2od9zfR1Rr5QGrXMUSMVBm01zz8YLxlfIzXL
gwWREDVQ3WZTr0O6kWbnzSHLKZkOxj4mvtUOrgCDPB7X4u3G8uq/wpmPANKs3PBX
Ewgp1K6CPqPY+uaOnkug+sq3WmGy7d6Ioce4ufeeHfynUCtsVdUOiqk1xRkPLzD+
SGWz4yOLM6iG6gf0Vp7ITHrXKgBMaJzVKvRRUM5FFoqwP8wcpD0KrTv/5tJwWjGy
selq5gJe4EWdZ7fbgKrJjlkPTzzBGSW0oTL6CeVorIlv1hPmDcAyWi1HBJR74ZuV
obcybfLvgoJTypfiUWYJcEB5ibFfLSlQ5niaunCa7i1pni96XYXVOP4AhS43qKFQ
kB3qHVtikO/NiO8IySGU3VFFwL8tYBb80PnjlFcnCDHPI2Cl96d2itukoYAx0Ozm
/strb5iEnKhttGhvJM4gpvNaD3YeImU6ZMkiJ50qQZmhLv2YymWTxd8leetsca5Y
MVFOndEo8CI7AWztAYoWyiVZjdJsARRBy2/wSVK5vc5nXtdJU39jdBux0r3CMZDk
Eh3PM3/Er/rKM1/eT+m7GJicEYdS5yxfyddxPLU7roxIBHqs3b9enz0u5XWCMY4X
rvinfA6ZjwFQQ5ysETDbjJa728z1KNWCGMfcDijuVlJ9g0Hq4kHuEOp5f0VzpcCq
BK42NIsbBNMdkld5H+WTEbGRVTHyTZ71zhsJPv+9hfKXYLKcvdfqmxpx6uepx9FH
aT9NePMtny9j7K7V6foIiXBajeNqTeuNacD05vJVB0sJTErgjKvfwPo0ti/dAUMu
24svRCcAE4vFo7f5+KUSsxDL8+6+Yio8oRFr3ZFJ4IrDx01Ygv5JyN02czuLFbIK
YDOqMozZitEkXIQD0eNVissWYZHqg9Oyjwof4yrlCEgbckVXp9QGAtMTXzYWroDP
TuKrk7bF9vNetN3ovS+RTvRQj89uKfcgCmk844en/yuP0vkc0MAmS5dGxIgKCpqe
2XO2dUjD6SSFt6HOHPypXyR7NhgTvN7RWNbztK1Lar90ChorHFQ5pF3p4ab03qLM
DIJlIDGyhGzVW0t28JNbWJQFKTW2wf2oi2QTg1RHMixQhqPwlzr/ODbuW5JLrlc6
wZ+KyLtvr8VBzMqpOi97S/UQNB80AxDTJLnVon2hTteuDSn4l1TfER4MedtJXrMx
yJgkTJXEIC6ziMmGyIRB9vwoP2lP2b0SYO3DSwSAoewpIrvHe7wAqTZP6WXoEP4B
RG0F66vJXC8WTP/SGW8caBJsWutDwjIPbmBOYwsUzHyaZhwxKmt06MiWVngkPJTP
wW+JN5JK+obF3K5teonLBOdo+prYULNUGMT7iTFoUN0npDEJ9KTrJYW0EvdgalI8
BTvGoVXiyox8ZAMXzueVbRhT6gh0IHA8nCVKcWbOmf+dDsMSMQ56Oo2A7cSov8WQ
INCtTzfeRlvd44xrbJFGeZgsqqkwNtdvhE6fNybxlhqV8/qbwpFKulPOKUiYtRmz
NNXsjcm3APzVTkMRaUwN1YZooua+JlgKLRDuHH2n3r9t8FXGk9qIfJfHDPG3UUvO
P85EjxZhnqHymLg2z+wWEkrgdbGG77Nu2OWrq0jB44pd1b2Hb6Zr+fpJ71P2SQxi
GQVMLG4viE9Gyp5X3BK+oF1f4NFyRLAgSLlbTbCMdCKZfAPbczuR/Wle5Y9JBX43
V/JiSsSLxoBUgcn77Wu7njF4lB7LFOzSPQ3ThTeAFrc00OpoSvO5SMeQzx4g3Hd1
A7/NyjQCqUhpQBmC3EDO99yxMuVeS0JALtf8lrDoUSOM+FI4xSfcLo7vX5XwlkA6
uDU2JooyHKRkczK9HsPDNr0AXWpF0tlUwpeYb45SrDnHGH7fe0hiXFybRZup+tWv
RiaPOgvqq2pf6vv3s477Jzep25uGXjFkHHrGDkBDJJoVt1T0f2RKUZPYv7KtCa0V
WzkRuRpIkoUHj8WD6CmwlC8BZTiJGNFSjppnDgwhxrMOnc98qKxwUUlo0/jGW0DP
ElP8j8NpSU+62NOBvnxfdUsp97S6PnZmVmPA+mApwJ4LgNqLikliCvB0gOXGOiHY
SnShbkiG884aYSkYrN5xBOgjIB+5l+OAMOTyHBh9+VdBekGX7mkYxC4jE3OM6yzy
rrpv/EUxLG8qpJ4feV0Dg4m26m2Kl7XpBOoUSLnUKHLGljh4zLLj/b6851oSLPkk
K12TpmAmRROUuTJXTC7BTynvsy3OUeQmaSfLYPP3BRJo76VrZFemF2lBKCWlhzgC
nuvHqv/+lNRw8zq+6lIumKxd5c7gBTmOXVQMn5J1qXQ25mv3HrbvDiU9T99bUt2O
LYDNUP4+nGkWhr1EA4FgEUJctwayGraCX1QmaxqSgPcCYiWB3ku6KhC3CFZCdYIf
q69MOdNdoO9pRl1NDFjgq2rVc3bvAQP0vp6rMJNdZuDCc80m7D/snQtpMpNeEbZh
nkdfRGsNp7e6Csrm1WQl9dWjIR54iaBlu6bvhKlAWRIJnxN3DkG/kZ/6wtBef1rv
jYPGNv98HxNILoAVyFwpdy4NwSsPil5i27cChLA/Xb1mQHjXn0BmxupfY7VjBDpu
IKCndkJj6Qfxf06RnJAr6IC0JqdGR8c623mMV17HxXsY4txKcgglt7pb1gON/Cpz
LzvkXWY2ZHX9z9za5Yh0zJamtF7WwUUWVoFeJ1KogWY7paRRaqhJa7rvd1DqP0gL
uFEtNIsxiWRoS+/pRUWfsNNTQ/bqwG30zq9Q904vNtRgg1WLv7vXaV6k0QeJre+K
mRYX80p+wGWueLG+8obJhCwFMZAvPdFhDQ5b/fRCJs87WjNUDqB65gqKx0j47s2C
G1488MN06QUKRJVofXXo8KxNeEGtOcJ1FZiZk4J5LI9A1cBS2pVmYXLuuYMd/TpE
A4Te+zbeFCyKAWcE45ZP9Iy0Tri285t+u4Q7YeuHlTWymdJi2o8DGVzqP6scmzfM
uXTqbnhuceElg5FJP8uCQXyTKDO6uh/TK2k+K9dBrbxAe5T9QFLg5d+4yv7k9ZlJ
ReBUbWUwIBChKs8pSQCn58RHnpTZFYcm318cMxUAEOExPT64uASglNH7xGa69yq1
eddOvabRJWRcggE/c1ol/h/ZEYWivpty5oIqx4xu54M+Cy/LRF2n3rwDhrPmSjHb
jNUacgRLZVGS5P4BI4hXpUiTkM9bAw+S7b00e7dft9xZuaOSm05yvf5vj8poyoLJ
cpswaC5AgYPbAFtGOvS4gdyBuhkAqVC5TH9RkBChtUodKIs0F6SgdEIAEy90IRaj
N3S56qKvaUnGbN/zKXGcZ989WG4VWF6rcsRhxQoxBKdgtLBBmh9mgJBTjjFoyFpn
bvJF68ZzZoX6rFY9fxWJVcp203VRiMaeRcRt7Pjhu7Zk89dMOjfjmbrvGAggAfZQ
aANNmifutDFqJNPYxBQ9WgAdmH6pcP/J0JjaQt1KmkBWgbye4Qg2+f2Fp3BWW4dn
COe6epN4HYLy1hdqgJB5md3mDNsCznTjmRqAwV/YJYpRi/4WXIAVdrBvcpu4UPXg
t+uQ38+16JDN2GKnqdXeccgh+yjLB1E/QM69BY0zWmNXVppvOBo8/m28IBf7yEMK
5Dc8WZLsVwqynnoDx3X51wPMFJtX47h90v5yJhtsP2+Wl/9P+3Iux6e+dyITHT7Z
6A7VxTZCZGtR2twkAwjLGepEvb7dAaJeQk1M9/yUBSWg3nqZqRYemFzAkH6xKW0G
V6B4G2zIIJXmNS7lHqFDe16E/ptsuuCTkb1DOfQ64AXZL668tEdZbjn2oTZjL17E
ye8IEgzfn8SJyelTr/a/kgt35CGLnQ203c6y/fI506gwW5qgx32gvaEmF/ngq4fw
cU8wZzocLW2JQPuOB58rkdaYbvGdWQfJO9rHL5xsJTL439o6G6mt2YGb0TkLDS34
ITO7a4Ig1yWtf/samDTLKcENdzNGpahyreJvAE0bw2FcMdIyx1Hql+0YUWOJg977
mnP1+aUnTp7NLOyKvXdSCVaL0zPFv1jG3NmOZ4ihM/f52QfqJtR6pc1ESMBROnvq
89FcT/rtIDpjlno5IRDQCQ8Vf5mu6DkJzWD/0KmmL6nvFfr9uPsjKypJXWAiTap6
B7yBWbFKpMduBfQjgpgkAmshN424LU5f5O0hCtb974LiBazWKdn61Uz2oKDkg0tx
rSiXBMPo2TdM1NhWwzqTAwAld/JBu2GchfYpEfvmsP1NM6ol54oA+MT8DYPHX28s
QByS5tevwtcd5xjyCesUrRjjCT+OUthuBy6cSWTC1lb2q4cToxscduA/VdR0dXad
zj/zdjNFLOzPe6XImvXMc26O8Ngg2XTtG6niCi2ZEC8v4YH10N5nX6hmJ0zzH/si
XDEFrnpHEP+CUZY239cvXWNsh9Z2Covp6T4WL6v4BsF86PijLkMe8G5lhlP79f+t
wWSCD/QaxqYMaYfXqakvWcBERJNsPO6BAwyywzWwJUMRnAo0NPXnQNEwxBOiE3MT
WNZOmXccGT7yeg/OK9N09HaTTI3I63Gwedn9Nub7fPbe8lSYXwauetgEByEvD8gm
HlPheJq8jxR53NvYw4LIpR/EUbjrWeZPFBQ0j5gMlsbFX79cv1JJGb0GDXqsYbX2
L+Si4oopZTlESNaIcCBLBWdJQSn04p4YyOw3QJrcla5vRtEedi+ZEpQT0kHdNQB1
AcBtcPboxM4aXIwhEsWEl7kUr54l9DEM9zC3xoNbCmpM5wz/HFJVvzhks5GAYDzl
Y2jJi4ab6ZsGUumyFzxEShWteO/S3tOI/yp031QrYjgnqoO/bwaTCaS3HXUDVEW+
c/M2JsFmgU7DQifYAXplJFBPL/21ceI6DTu226YuI9D+Q58SC7tNH7ISMMnukdW3
HvwRw2bUp38thYW0l97uQhZweG+wxyZ7PqsOGEQ6hk8KmTIfgE7tV/J9JJMj9e1T
s9ruClDHwfwuGircnVX/Q6j0avRtQ8t9g98eHdV+WkYJEd8iX8MGcqpkrIir4abh
/HR/Q/M2et5p3PhSzecoxOovqnYjXkkMmpu7La22S3B2DYLvWrBTZEWrmVQ8h9Up
YFbJayQrayNVF/jQ0m0hCmDwf7LKetXuchcK8LGOKHhRWKA9Uyr8SDe2vIdrqg5h
9V9P+5tjrEVUL6EF1gQatCYEelOQQ2Xjq+YBaYpWTzR2P2ZusW28h4wGJboQXWBF
7EF/F4wpLwvxRPyjeuVyy/ggYn8RO6Sldp+mNroJhAJH+fAuVB5zoT8HmjPkGGSt
mDgZX/GPB6qIcDyxqf6biB2MMkb0Y5Dqd5kR3mtZrqvQZZxI0B04kCXGPAvIeUBw
xjeAvs/T1PFcwQ9E9z+tCos9fBoU62rQBHXSYPqqAr4jvW7dNnCp1T64D0MUHfnI
2iLY+WOFrkh515dP3ePInXFza6GPPzauH5F3cDfSfzSiWr2rVbfi2X0Ev5bnh9AU
69HCuHSiMa93OuVbFVuQv/3LW/4ySu/EUL6YTph7NZf0M9i6SCycRgeKwekIFSkZ
Uccn+5hOTvFfJl9CNukeafv8a9OGUG2zMtPhlD7zCeOtcbkx22QbcV1DqSOU8IZS
6XkgA2K92+V6S5ZQucuP58O8F1wx6P13xQSJyeLUz3/drkcsPVY2CneCXq4FFIeW
tFy3el8CCXX/QgnM4QCpzLNJfdabw5+RhJcnra/TSz7KlC5f0uJL3674gCQl26sh
3l03H77TD2dSGT1Qtavhxk90eeKr5cU1C+3dszV5mJZlyywG1iVfjIwVdFTVvuVt
7fQ3ezqslXQtP54O5OV54RkxBsLolO2XKkuv1yFoM1VQanLJ4R/yr5mwN2/VAjPC
E5aavna6Px8Axo15D35lz1Ro+ndlxlo1M1tT1/8o7xYWhMOSDP9NT16vk1RLITmO
1gbNuTmHGBhJZHuQl8IaFC9mTASz639JqiqlYGsdP8Y9W3eZ61MnPbIXCq3XW8mE
Iz6AeQIEMRjWYlfaI9xyHwtvkFHgibXYABgl38spxdchmZ4TRw1Z0YFjcgk0xKKp
zj3fOOnWOk2QahHUjpgztCLNqzECYzJs7BOl4HTl93pyhHf152b+wkTce978xdld
3aq18DxJeogeao8QjMyVfTvuZGSIAkQN7AGRu/H3X8vvoPkMBWYkldU8EQ2UhNre
H0aw6DI8qYNU6jqxXT+mQX6wHTHjDJ+hbUbNIfqqq25/s+q4xWbaWSsVa+YikBYn
mhHUsi9F1/zp055UuRff+H1mP5mjNymSiMDGxgLlylu6VeHFaVQnAVgExyoCRA+/
QFbY/65JF5TcNU9b6Mkd+2JgpAjddOSxb6T8ApUxHcZgYwXhbLAS1nCIqzsJTlvw
SQVr20NOvRilFtc04SUn4Td0nLtL/SWwrQH0aJd5PVeHIUyPRfha40d9aQR+ui6H
MqrcE0piFs/7CIZVGTWSS3+6svyqhXxAr/PPb6nm9J18ArhSldvjeiTI4VCOdB/W
scgQQYPx3232VCAwdNOyr7t1HCCbiGqf3PFtPFNr/XCD+FqmaF96FPYidshs1f44
D9/r926ql/SoViRSEfmNVCYGiR6cii2T/7/pIUiRMp+q4+0OFs5Aip9neItGF7sr
OZTlEbeKRhtvI3VxZVhBkCjLZsqhV9QV8ybm3Q4m+b5V0wNV+YVTfs51sMDLcvwd
Z6N4yYBAW7UuihCiCVxkWn/BI0CDWSPXpIvvBDgeoSQCP5t0uk/FxDKfnI5JRJfI
wnu8XyCpvLpTE4ow51cTE7yTBRIABSExN74Lc8o0iDzuMZLgKnldckzwt4cavmZL
nxSmccFINZnqkeJHBxm4+uvt7+dVWE0DIM9WF87Te1rgAYEBX5pnzK2/y8p58ioW
DwhMJhT6yVJRMdcnRzXw9hu3CcTp57HsVrCAqP5BdaZ2noOjZVsm83bjVf6D0O9n
wDIW+7KT6E7azWMA/Q3tx2D1KHktEeFDsZcl9UWWXQ5cgo4KsYRv4xtE7EwuxrT2
IUvi36H4c4u2X85W5N5tCApscPZPHIpa+wuh1UuAPcJ/d/241b2ravcF8qbhdJYl
67FOw3ig1b7HG5NreKqVCCHTE3ECWHRdGcEfwBlCj5LSL3UqY3cN06x/Pso3KibR
wo14+b9vu0zCqXjBDVclwXYbejiboIN8E7AvKWCx/kYn5Sph/Qgz2wtk0Pmv+PiI
OzkHJuMg9iiAtTd+kaiBCEMUgfBiMHDObmEe1IRIysXXVGWuPBo1GBaUhzfb+8Tr
0QkNARbMFsiXQq511amvNCOoNA/6WXCc8RbsprTyC5H535QzUzqJAzuXbV+h3Bqs
02EWt8mlJt6tjZSTyvSyv74hXLCGixCOuEunMlp0SGNxeVeKQK/WuZr4zFnAxN7C
TviK/uithzbpb4YnPYvXI3Y2fWleAnCsgzeTO57GI1iJ9fSMyHacSiSoFZFUF660
dLqgxeqEoVyUDP4LWg2o6tGusFoV2Jwk3ZguFOgcBOa+dgD0u4gW17rbv57Bscy3
Vv7SKc1fbXhajmkTTyt3HO+5edVn2ANKPK5LnuFDYpB6i3kxHn41/ASxtuiyxeAM
2ooEXsYFD1sTvh5QGDe38laX2nN+PSi5yVFjRGzU3a1B4vU52RPbl+W2MX4ENnQ1
ncx6AAh+OVG6YS8u9SGkQgdMO8KOTWhUvRqwILKOknqeVRvrOOg2EU/3ITLHNtgT
Df5MiNMZcrk5n9OYwu3cbQdB+ppUfda/knK+HI0HJ98y0aVKTLf4frWfPQab6KGv
Ow1wQHEDvHqgoBrChXkyeI1PuNrh+nrr2aTrAB9WLOdEkui1qDoyZe8TEVe245ro
+pR1L1v4qhJudgsr04JZfPGm8tlhy12ika3qPB3yVGZbUPZjMbs6vn2G+qETXYMt
MaQ7H5kaFMZebITWvux9yTU2/e2UI/mqLtGvhPg2Va6mrmAXXTPOncjE7DhImaFu
PECsFT3DXfLRzWsO+PpQaOAcuh3mI2tYml7G/qfZT/VxhOb0Nl29oxJb2JBmMnUo
3lPnHjmPkBHcpYCaADUt3AwmVlKcognldS/ylJo5QTizsh6fDeKBr3A/Hdel/TL8
8GnVZJgfm238/MYMWP4V/QedNFlHN17a/b49706N+aVyTfzPR/Lc5ojy+SPhmAIO
l9aV/3w8/nhUTOYNdiwlbiMmib1XYtLaAzuvrqAK6AU8rEfiNsWjv7KTWpfjID9E
gatodk8m+R9OFlWXDMqKeIOpuPFx6P6UQxbYPvlEpRojdQY+COF8tqF9btjVPmAO
lN7WO8XmCuSPXfAqfYfAkcNsZEGkysbj703T4TuTu6erlTOmbdiS1S4nSkd6VFCO
CEyJwlPL9ToMkl8vAp7o5FqQnoRX7WWa1onZr2bGdVPUqeKmaOJjvalVN+8Odddc
S2+2g8dmON3cFlrCLU+H2dIqztkgPLlFvARVsnL2GzTTbfxbuGVsIaNIfs76h1Qp
/4bR1yZMbjFPHvAz6wpb0YOKgRjoNTqb3Qr3iNFzMakJdqGARARR2VbjITUHgXZ+
YCTiVF5jv9jZQD7cewGnN2Bk4N9bXeD6Re1f+Hb5fYLIsY6aIG9B9U3UAWrQ1eCe
6IBLCFsta/l4EGWaPcWtzgJoTiz66zlV6yxb98MOk4ZzuELMiYUXp7qsZLQDq0P3
vPbQra2gTI6YwOThftXurLqh51/bC1XhTpwhQbaT4ExINQLE+ieADU+af0tqmOVE
TZFQEQlL4aHFLyNMcvtdoSkTw0hYOWxZjdApNwiDpL6WdvLQGWK2Jt9vze82Vbux
G5CFo9PUyiLLcPAessNNRieeKk4qr7Dmpn5HaIxi62Y/iuzUcFW0nOQ1v5DeIYoY
MuZ3bMSo1kkSnTvhjV3fMaOBQArVxYeZ4XwtZA2DYF1v+bB2SgiM9BatcjWrWLl3
zTACjyuEv8Qm0Dhw+XVg74qWp2DzveyDnq5a+HNouKbKQcDAptfm8qDIWuAFKY9l
TXVtPeNoMUMhMkfPvSnPxuEp4VzfHM5Pyi/TOCIIJCcnqKQl0B0ay4gwGRpvmDlE
ubWmAXkjDEOY4lxHgziNt49kkK7V3JxjI2c1XpzTq/mYZN99PwnXvxk2HC68Sn7D
V+DPy7pJFeqvMYw4S7Y9PhMrkYSR2P7NFZMWsPw/QyitYqX7CEtik8ktEmXl4E4R
dhvsTj57vxrUstan7aQNKBvn92kLJ7U7/+omoGWrGyxlrxvpRYudMZtws8OjJ7tz
n2upcxi38v6rKHdUS921QranaPnbN17V5oZOxIDopwJbpiXbjZ4CR9UDDnynBxzF
FOILQkPcCOfHKYYi1SUnOe0K9A2TvzX4CrCjLbO/GpUSmVcFjqd0ISXQ7wRJM82t
eqFYuTt5cTcn12X+B63l8+bTiZkPeSUkp03ndHtH+6UMb8aEyCJoCP3+QVMWMLhw
pWm3TbqNH+X6OHgk5aVgBsw0I5Y8TzCbg3vc6IxumJju/g+w/mwurr0jtlt5+ZaN
xyHNY3FRoYvFBxu1XejArC6nFPa20UbZAjpy3Wma5zMWMufeSHKK38H8lkB6mrIE
GRyHl4YK3ulWQQss+ssnRhby1VisTRRGLEodJXWON+mz05+AR6eHlVOWFmc1OKUF
rk+Mx0WXGvbCqrZxfqr9neFtGZm/tx3BfqsJohGt//l+EgYcqLdXvgOBXFSA9gEh
hwgwRGx1iYuRYBhA9jqiOwV5M1ebJ2o1bBCs+ZLvBOadHSqxQzrDXQeyll+1Wq81
edrd1FwkJA0eZPagBp0XqYNkReHzXzjaXRcMYDwfeVQIXyW8IxpeYRJ1Icd4GyR6
e0Y21Pg3ozlwVOG0gDOOAJYU64vspJqaGHXSmG09YUFLpqM/EQ2Pr73pBn9lSr1b
n+wdNb+6qjtD57YD8Xu/p6BTkjatxpCGNVrdM5FAwAUdqbVapYacntT62yqeeQUf
9F0uVRXhO6mpJ3p0WJUoKv731RG859RocXSm/zXn9gSXJaD/7rQk86+eqwMguyqQ
umpMZjXNOQ9Tb3UfkpCfP8qLVEitLHWiL0Zt9sKVwLkB1WjxC/rq7lmwRuEvR4hd
LxKEged4ZYbnQFbs2NwN8QVKgCBsGZWZAXilBFmppFhkwa5NVRLDCwr1oivcRcUp
L0HA8Gt0roB8LSVM/aL55XZx73Da8F+BmiElp0O071igPDZ82E6gfwhHTI82O3TC
jqjhW/DcnHodcKjjRU0yYeUmSJnzgZi0WaLJnMFNPQ8BSKaWuuuAhmwU5a3bYfgP
u0F0/7O0sBhbreMg6PeTw7O1TS2Pord7s+43pxq4hT+bc65Cliax4+e0nxfojsvI
rgjyi82ooagrUvHjdRWlSXsShO400MuEDyyAjRgaRIZbA4Yv2taJHmnlSktoooW8
pNEjlZTBxKp7QE0DGdGUY2JIgizqS2PJ8pQdcPhocKSg7013UPdVxk9wRkzV/vaM
r7n8ZonuBWU5IBro8kAEDw7fDTggVBiU83GgOFXxpIAYh3c3xOQqQea1jYI1GLQA
13+Tcs1fAI5DYe7J1IHNCjsnRjkungdxqVx+2R2wVhsTYaombCqLS8ElueI4RO3g
Y+vhfpi6KLbqR6wljOtWhK0WBkcK0rD16j2+jNuuXcPt+dNRRqjl/ohYVPkq1Qoo
ZdXE8pcWyL3LXRKN6DMAxCBFAzpKMLbTNd/UNe65+rULDJ7dKmeOO6FnvAgbD49F
J4QHu/Pwuqsb9jYEORvyNPO2gB2O0/9nXwFHW6eE/6vAk2mylHQQcAFJXETrbBhZ
bvDcLcNP6VhfGzyaHRJhFk0nKSp2rM44gTG7+evsMSxkLZm3nirlm8a8vtrq7wxz
7zxo9AGRL0TRPvmZs2Zpm1m2PlzYcZd2+kePTkMEvj2HgPItcN3Ox8vCajNkeWXr
GSiIYsZtqjv6cTdZcW1yDsJopz9JNGlXse9jwjugIeobkURObwNvxtI42qfFBiRi
ZKZCLFPayBJqW2nbtIVlU9H47ePrMn4YCwEThI7PaQQnXVYdnulQyCIYDYLGrF+q
lanWjPf6Jss2uadi0tFCOdpmEinAC4wlkgIzvaOgK68Jcc2U1Fj5dfuwKyFq+vMn
9LTRmdzvX13plBo/kabsxqrx+XBZ16MjYCZAbnmcwKQCUgeSGIDDKLtRJyVIaU4I
Bn6om85nt/HU/60ogbzQphJC5UcCR9eOTUijcrbGjya6Xkon41ZqeML46Oex7JkG
B2FPgb+YQoqEFAEaHNa0iRyQ994y0UEEsiU09mFKS8GuhlUxB8fl4Xp/VjpLNOWD
Fd2msl1X5dwmn4zjh9tLYrpFgBe7ohhjGS1PzHYewqFojPakaOJfkJrNqCI+ar4U
ZQb71oCt35yfC/epPpEEhgfP/dBm1ohAp2vD+ctGH3xPG40Q2WYmC/tz3DyupM69
AM2q5j2QAuVGEWx67Ex4f2L77/vFJlHffD0pm+N1xGzaIbxEUY88ZtZ1sQn9WSvX
aUk7DGMn9C9l/P3QggwDTRfieIyGwB8VBYU/n8XeHJ+C6y4NTy2l8U2agTamAe9s
rtgxcD5CqOCNneCWmwqQmBk0wwOO30VDqkZE6C72aG1TWrG1PuULZ/MfsaLmEVdM
XIyTcNX8Ft0pDJqubizwjXJ/gEFxKqPLR2O77rWK2Lvz4wKDxvnRTrEg2HQDThFj
O5LC3jhUJUepH/W+RW3Oyvao3sqwgA3PMeHMeUczM4kkXqM35yT0N8hDZbKP+Ocj
KWl5kIiehfT6wHicxUloHv9jusHCeMjj9LmH1C0suF63xjbLguTHtpIVp8k1rJ1J
Lg5ltWEeoRr/WMStbADpPqF50KBF1yKVNlSsIpD/+TJoRkkthtPnNkvOJFdAXMR5
U8VG39vNal86iZ+3gasR9Vw6nWQ3nl26R8anR3k/ohLOTT02NfDXqF6Y/u8eXAqW
9AKvz41baRKmBfuUl+DLwZ5xq0BDGyGiy869Fde8BMRh+++nUo09UFAGoMRoJP+1
l4iNJdDlWQnU3YqDjiDnsApXOUjN4Pe84OGPUuhHyu73GOVbqXGJQccJqdPr1WRT
hQhcC6qeJLE9X8i4UraSzH2m8UPXM+t0D83JRFo7i482HL7om72+h/FviCN9/hwt
v1NNSsBzl6WzKoHOkTsbgRgXgtWGFg7KmiOE8FFt0WrQNC7p7/gCY9nKsnd2PAVz
xHftkDIhIbOAsLVxt30Hr+4bY2wHk7F1XL4UNeuxMa24m2h7lMhoLLTpaboGx9Ao
O2FqAiisBMPhjfVSBY0IlTLI89B0QIrb9BDOJwl6hQWPB0q+49pljB5oR7i9Q5TA
HxLZ5UQQLrV2X+NGbQWHiqpMviIIjmZNC/vHhpLWvy2iYTo+mRhWlqmWzOzhFPU/
hNqr3qxeKGW+cuivxsWG64L37rDKwBMBneiFqe6v+TJM23re84r1VF8T9nSdh08F
r5AZiokt5e9XgitPOk939LIt1FyDqRuuxewJArxOiN/4kT3xfg4ZaJh49XKAEKF8
a60qXDPR0OzpJTY9IXo9hua7Un8uwS+Eq13xvDly1SuBuhm2EIQJXLP2LdgNOwYP
prtLFxhlNPY7kx9rJBhrnT3z4fj/+/FROZwwFc96l1nbyd8EHLBYfNBrF93K1G9o
AXB7pLq1OXmK8/5j4nEonW2HjnSbHcP6J4MaJCmZW4lVhlrXRdqEAeTZBteq5V0h
U/rNzKXj0LNQBlc5fxC75Kh9LoqfqAdhgtUfzOazoNMcxGvMu1JoLoZSl6+VA43j
Ecb8a1TisNddycqjh2h1CPMkYhIPXGsnwC1Zask919J9sRWMB6wN//IWcOAP0Jor
n47CGLVE2lppq1Oy2SM8KgJVCFyL8NUpIyc1FjfbtxLS3gOa+qk/iBWv9WQwOTv3
rjQdDxmRK22Jciy79fOcJGWKgVcM1WR11TZfUwZk92qFUP7JdfRsozRcA1Mjt3hh
ro1rlCMLHKdZXmRMvOipiSujY3vkfU2fMa7wRA/nI2hY2dNnGoxf4g0CPVykviyl
vCWnj13Y+dk6guPo9XsbbCg8DZEj7KTmaD49V/UyVDI5af8q3MItu330he5J3JLK
+Ns7/ErypnbPiupAnzjsXK9yo6/bH/7p62D6wNUYIVMzAQAtlOdz4ChLvSGh2rRS
mWnHYBwzuO/VhrasJaFdD7kXdl5hPzyMCWYfPtDgHhUP43srcTnFhBYf5o5wFQSm
Isvk04Vh+woRibX4XFpew8uwVuBOAEYvMC2tCorukJNnbyi0ZSg7nVlKKpacblRy
0PpKRmGjbaKoV7r+gye7BhQh9ZcSl91ODg2rLpeWV1zoGVJ6zLZoq+0P8MQO0J2W
X+1cGxfTRFjsqI7NUusMm9hvFVa5PAp693z3vdQfPjlJI515oF6gEPAyEbH106mr
UL44YGhxqEjNF5FBkJ25nhMDtAXugoePcQdxnXjg4XvfYoAiYaWfmK7jTSrEp38Q
NNIN92Yq5sNH1dd8gJfRZYw05ndn7E1Kg74l0Omt61B/qVsVoYQVkYCQ4p7Sbbty
H09Gy87Yz0pneJhIFgNpeLT2muDmYYlx+sNiG+KzJ6D2b51By34eImRE4+cUUD8D
7EvTJVVfx/H2vx5XZtlp5ON7ptL9NAcXnUhfhSA0T20Wu73b+cCv5KoHCWwnilyu
Mg6/NEyzFa1f2nKhiv9cYXu1ZeNV8eYcPY+y5sF1apK2/HrTMlvrXQDFE0cacgdk
LAkO7H2EPwifvqd5PrSIcKt6Dgfhpo1vFUZ4WoJb7DASeI+sImCYkPkZWgYtrvsS
7j77hXDvynRxlBu1iwiqaeprxNxIVsZwuB80fuWXeNCMeVRvSTIy/EG3ye+v47eg
RuxDAA0J4onqsRUVfes/5E1FYKpAcoyyzIjnmTyih4sj2hJ9mwLSldM/D4DBt5qd
7jPg3dEh3+nGAJ5QxrBAM5s0QMyEEub/haaceYFAsNh6jIQhdi6ooLmcvEpgagU8
C/jg+6NTBE2Aa6XGu2HbnacPNFG/GQFg/dg1H13OVchv7DkAwDIMVygZftgpd8fe
enosjSduYdFY0JPIbQR6WRwCGJHrZGKUPeM9eyIyoohq40950Deudp5ewoC8JUpt
aIBwsP4i2qVJoLNb4OVpbuRCxgzYKFI5gzUe88jLmXyhQ3u5j0yjhz6MKyDQFkE0
wbZZThdF+eZfpraZIh3n20S7unIETVLdz3iwLt4B+STlfeX+yTNYccAW3xR83jdw
F10+xmp2nFbWi4TxWPNaatNttiaYxpwjnGBh12v6Ka3ymHI1dFlWXkUIc+RIum8p
AWiSA8fvwcKgd3yffpAKzxA0QNGtQ63b4myEjJNImSmWKEl/a8N0JzVtX0SImPYA
AujyFRQxaUxGYcvqVVKq0/mU+Q7M+TZc+0mY8ZQ+fURLMhtDXyQb1ztyrhKplHyN
/04v0YwkezXTd2QkocwI5Zid+1MjFSlYU2DrGUdtKensAWsRCDeXfyengg8jixCH
eSC0VbcnfGPN+QStCmBQ0wSEJxJIZWuKqGVYA3YzfehfVGjJ136CXshAweQqGvkr
ymEcWsjhzt7muxqE4ie4UXtn/4nd63bC3gaJ5PtZRAPpg7zF1cJc8ogEGUtJHpVa
LJC9RtuLDAISIvoWNpBRq0L6lc1Jwlr9pAYq8Q6RRedea5YGrZd1jRc9GagGaSaA
L3Y2gruzMbyDtpj6gqOFRiW3V074FRFMa97/Bznn9Dta05Ml3995GSaHWKucG8RM
pSyiTsGlSF/W8mWNTwoTsQ446sD1N2RpukkdVZFHCL4c+mxZeIgIHv6DBUHT5mQN
8IOQJowbdURZROOlMDGL68VYSYOqTH4qH3BYLjph8GikO6uNKV/zTtraGIx13kXU
jSjUrlh56Vriakkpap5JhWKhDKqhcb9HdFmqa87u2dF/wSVo/2uSL5cIU42dt6UX
VRAKUkbSkiJbqbeEZ0GiTEwijV5zCUqHfu9RISCmS4aplCHIBwne4b//2sOLlByw
tm9WUfoD0Z42hwUPCxu5iSSWiU/f2CAyKa+/sHaaRNXFwLwZkz0SbrdCHgOv/JiL
OMUHHQtZg7X8XygYgWS7zmxhWyY20rUI9Ez9VzmvrMPbFs4lb2zM/v0+VEazKn0e
dfuJAftXuJou27fgUwuA/ibLTtaDwoSn9EO9z4rHcR4jQrgBiVTiXVDtMuGXCwYI
pI8+mKj9PjHMClII0aZEyK79cDas7R5UZmHP6leKULU65ccFIAJNEsF0QuqdFuPE
uHOKlUJYi9Q/Tx85yZNQUEXvGhqJ/Z3YXNKggZYS7t4mmGyCFdW0oewA7rG+0GHc
yJGTGI4LQuiXFL5vnLBD+6/sBgyuGvFoqTOsPPJIANlrm7UXPzmC6wg8Yth6t07J
itsrwggX1l5tXdsnRxF0RPoBkkC4KODVSQJyKPoveA6aJf5SfI87ARhMguaCdsB+
n4Lwot/cHaDICtQX3Vl2vHJfoWC8A3JouojmH15V7fR5zPrMgyyKO6OQdCqHd7bQ
SwRkr9jjkPU5m6yHnYPa+urGmNEAUg7PLlBShg1nxJq8JSY0ZjOuth3QAWypnPKB
PaZaL39Zsak/vHgH3MlZin5WhaMGZB1ssa/T3W5Zse7Ksa9qWIGDgjGVegunW4xI
p1NiwUYihzt9rFf43OoD5k+4tlwmXwNI6vtzJ+SA1eaVaoxLVzsh6Y8R4EmtJdOh
ZYfPbCMNHV6MZseSmDGqNakKajM43sSW52Rsrmjz8KEKzftc7zfcBMr6xbYUFSkg
UeLIeHsfVbAG5wOFF8b37qHC56j3wCK+kRO0bLM2yhVDPwZbq/TTdmveoU4S8yZw
xQlIHemIcRAH63QcP16bi+uenVlMBKK3pgNk4UJ6KwJK5axGmcweAHjMAscJz/5g
cmEkq5+d93ZqLIPYl+Pg4xxh5dQqKhGM2iX9zMzOtNmePouFXeh69di/1cY61BwD
gciEVN3j0sR0WfpBVTbg0dHiWd0wQM19++DyIEAxsD3UzRXloaBmDvphvLFaXpt+
WTBTBc5sEhpg3+m0DZxTHh0yqNIY+rB/DjR5CLXLYaJDOlK12sY+NdDkRX6JynAw
qLuDq2kU1FhiuVoEsUMQpRtmNs5KBjHnHGhbK95AmKGOaWCyDKhqodlCPLgQTl03
JZAnUTl6yPMGeG9dSgE+Dhnot0VIwaQQ9IWBm8K7XHiyKvEU8bYZqEUSgc6pRGfN
hSBaaqcjgkNWNfcBOS5shN3AjUyiW7Xth6S0JAEaM+Lk7JzhvpwNRJBC1TyvYEbi
dH1ohzhChwct7FVaJaNn0t+bGj72nUJdi0jexgOnLk9ysbQbGF1IX2zupnM82pPs
3vtgjPb0tAJTvbKH+v+KJu6qzj1xGGEHhhs1ga1DtJsPSsIB6IDLruEZOiFxqAIJ
FidEuhxnVhb21xPFCKiAcY7mPaKfPDBPNfiM8i+fo69GYHsq7sasJzT4iYynm1ik
dHVWjN36Ym1Ym4T7VkzfZeNN+3BKk7DxGx/Oa10f46qFfLuMp1HZV7vmlKoi6LWa
nGRSI/ZVlzddEYI5HCSIpVHic6oI7GUYryb4f66ts7VdcluaosIhwTfbOrhEC2mv
OaQKtx2LbDwpKC/mzF+mfsYe3CqLB8xXdXyIYXuaK0tts4kBGifx6zpRc51fGH5m
7+VonL438T2ndctLbQ08oJYXvimQOjjTXj8gO/JwxpINazuTRQmNvUgSGFTOffqr
p/HfOxyiUEklL3/Uj/8hGQ/5/GCE67hoclKHs8ii6l8e0sDQg6cUHDPPQunVCDqt
qoFE6FwyXOApnjrCTBWziKWD45urmXHG6zmxfvR5+XdcUJN9r5BV99r8x6XLRc3q
KS3vc33M6zewAZz1dF/g/M+xDDfCFEbZZDdq0gpMUjM0mjcxaJ1yiVxUrPQGhR00
yibTRMI0pNYainxQ88rsWW+RLifjScDsofZWiWsT/ibCigybuxAORkuuYqvG24te
ibzZwqWNxPmxgRghDRCE3oeDbFpEd0FIAzkj0vD1CkXUWUwPcUgMhNOKa51xHUX4
W5o21crExIGIy3bRTSX3Smc1D5wENZXXXBA+3SWepO3hzsAs78ljXAC67B8Zcmh9
MoEtnZ054TxDBss0xW4d4sWDdxpLpGOZ/D1FwqrrL5MHmtSOg9Bb/A9xhOdctHPM
X1V8Qzs37H2TzetjrsY0fGDZ4OE/vWHeSRrN1JcuiDdJ2DZag2ZookSlaJ3pOKJx
t0ctGJaqPXPwu0zPG26nenrXG9oCG5+pixc6mXeXRdNteMCaafk2xWecNDXy0Oj2
CKgrE1mBX0VDuDPLElOVfo1y4uI4s0qp9FpZ6yGFHO7OBssuDnhfn3Fqo+QxB+U2
kl7qlhCpCbhPBNmtEcEpI8QxK4f2WhR7elmEpdSIWpYNxgPgLSZJQnCJHpHZLx9n
kBInMPVRRQCPJqlHlaAtXHWB9qMu96odE4eNwynaBRzDKwgTQxto3vs2/Lske05q
ZOpG6PPsPPFP86ON3xxZVlIMH2lirpQQM4WTf3XWAdRyLYptc4cRT0bK8OYfIW3r
8g+uZpREuyI6FA24g14ydvX70foYiAq6ciIf+2NBJQKd0aOLLNB4RE3Pd4Hgcotn
PwlIryu4HhHyA7yGi/qgMWuJZT5LePgUuIh2Ky9mc1ZiSBI7G8xlfygz/8JH/AYb
pU74mCmJVTHARnsXivJjVi+42wWnrIXOVwzDQFHbj4SkIDwLJdT/JMkIcBUBbUqS
Vr8tfAxGMhyC+IxmNASji4VyFH7oI5OI9M+3Tpxcc3jUZ+zFe1zndHpH3y9WdJih
p3yaWidzWZa0CxQ1aT9OX/ipj0FV76rXW9uaqx8QclMvC9qsjIoCoFxHh2RI6vkv
mqMyAVXZoKzWd+uyVb8JdqcyEDmdYqFAm/j/O469lAx4Pc/xmLiLwOxDE9nk/vLJ
EpffDkaTZx7urPBzQMZbwIzRS338ATP8kZEYvMiL3aJK/gZ6CAijQSfGfqTNnHF0
l958QEXQoNgypo8NMl+97bVj5QcCLQBQj1PbnB0zKoOCloXSEpWGHMQpKmj44tPr
t+vOg/ebEtfy1TnCB0O0DX9/MH5D/tPfn5PnkJy9yhwG0Lhla0RMdFGK01p4lvlX
BBB4JY2DQRY58BE3iXZh4f7xSNbrxO/4UijiHj5ZGVWLhXEMZVB/Kw/rAZzB8VuB
EcR6I9yoCjuXoVs1d8XWou4TsjPSUbQeeeDVJPa4CYVMYUvHEQi0afX2NzAVX4JK
ODUfQNc+ugucH4O4ByQDiHG3P1yYRATgN3zk2o47oIbT6w3KKqMWEc6IBgyRcDik
TatmxXfEAVLLLecnnFjglO8305uc/esPbspff8PqCX3ffZKeVZcBwYgS2xQ5vJuV
a1h2Rf+URDHT9tL5EWgSUED4Nv0cxXtWT3ORYyjl4UL5rqu/yyeePsSN9KXSvgc1
w/2utuAf/56CcouPnYBpX4BXubjUQ2Rxak5TT1H02cUTdNDBvQhVoTkCyzWxhFD6
SCoxSCFuFFnqbuegbTSBtcDnEjjyf8FWlKxhEqfJojF5G3XcBzM99XJO/JQirSTr
giizLzfCmolG6qsxJf2zLGL1gEhinR4kCGj/sOY/FB32rz5h8hQNV4rskQycX2yj
bsQiCkMTjpolDRLNZkgnJDiULCU1/ccqhJcZ/jyUNP/kvj8KXfj+8uKLguz5NFIG
nI6Q6fdGej+5uiR120Dubuy4dlR+TL7NSnyS5zsddN3nBi+hjCW3ZVIEd+JsHkyo
PEjOisaBBMny4/N9GnxWA+0WR9oNorHt42u2/+P4kteF6Fzo2GJ2Dbd8OxxmyHyd
ietn823+6T7Gez6k4RbNfdpwX3VopmqnpvxWZ15HGIEO+ri4PI7aPhuF6L6JF3jp
cJdUXcXOw81dmqrB25nuOnhV8sSopCz003mA2MVF0GiYdp5wNE56Mfi8hFIx7ryl
Y5sKkmPErfvzzz6JcoDQc60t8Sth+JbzktpvK9XxuJiArsHdoXSuTti3upORXC6j
nDF+vZsJyILD8zgtNO/lEQ9hMy+mVwGClMMoWhlw4wSUxUhIimBb8YJi5IUFhxUc
MTGlNpriPSAWAH1irQhUgBNT27GQ98ibwslzsA5JNXIaC75lL6FWptXy5trsA5KR
OCMPPg7pBi3imszjzTWKymWCimzZW/dPjqguZTrbdpwX125F82L4iix+WBJcK3h/
DBk6OJrswAC8psnj7kMs7qDb+oveln5CPsOJhxuM+YztQR3Me7B+1ru0uzIQzRlb
f1PJSZk1bnk2d51z1kmCmoNwiXw6SbIGH1dZDT3E3TOWLDoTMT+AHIePhrh3nYzP
nTuJYnUpU6wKJ4S1ZCdQ2LEtXWPsmWn+Ot800ljK4Use74WJTWGr5CRaLWscoHnA
ifd4Y8IOj2RlVzjdqT7yCbsdi2UgYND5gfEL7J/2Zy9szpDm3XHC/mCATcvqXqWP
UfNfa2NnFQcqp4VzWYKV15bABfXhVCExcXU1vH27X1NdyVq8b5psFOiJsAiVRU5C
HLt/Uxt+mUprBVUn9Kn+D/E5arAiXcsgoyftJQjyfsbWVM2imsPgXRMYD0Dr/HEZ
2+SeSUVcqfgcfm4HB0KuhzX0o/+OSsXoNkLQUK0hGXFQTFcfIFQidXrO5B2C3yq0
hOhxNPQirei/LpPM2AYYhceXAj6MKoUjM5LpexCv7eh2zNSvU1tfet04COhLgTk2
bUx0l0wytlp8MyXZfi0w0YbXBJSK//9MPLOINl5pVrEqkO9PWF1Qu4egqpFXhFwc
LBPGglXQFpexwN7WnKDvOEQ7x4jNG+q5OIUo2/yKUcRGVoDzIpMNIminR47GC49F
jjdnPIyXNm0bpEis/o+2mFkqIr+iBltRBR6PhxVNWUizAvFhhn4KbPne9Gv85Ycm
9Wit1vKFmO1sg97CuD9vjriAa6HmyhK+CCwSEIIJ+85kYt523uT+cgSfDAEec6CT
WSYxhoMAkzu+G2u4tyBdWrCjqn3zp6sDUhQ8s32/X9KiUrc2q1oSddcHpWC5agPD
h8oRdwX9HyLIt2gCa3qNCsnKS0BzYq1uWuwoJ7Zbf7EsxAn7UNQ4QBWLVaOO3OG3
191JSQ+7EKz7tScX95Fuo8dC2N9ZSimUVUluGG9xbBkmme6xlVO5JYcfV9TtKW1s
ym4QaUQSDs9GYIXYajnsrcWIGjQCo33lzRTHj6qc8+kR1r5/hm3DKEC3xHWb/xzp
Le9ei2PGxsaoq3OpeHZks+4+7hha4wsDtDY2Yy5iLuSPS/nFfsBiNhRBrjjxxcod
uUUBAiMUdnRTWQQMVCuW61RZlNz20YQpIPr/hyrT9nRITcPgLuLsZ1Ds6uzNNqZL
a7ZXARjgp3+324SBYV+dmTyJ1DCcbeTQRHpY1GGbzc8tVteH8L9pjS45DqiWrSTw
dYrmN5963xzWTcoq0Vqw223fCO2ftq8jQbSr6TaAYdFpYCuUP0xAg1ZwIi6HzcE6
VdisuYSUcOFqEl+BvEU5WqzEIiOw9umYsBX+kqafM5SPLGHhtQSnzUKQMAnt9BsC
FyH6OxpzMs62DpjqpaFYnP7jMnzrPGitdr+kRW3JT3yI0otn8DQQ6XzY1FslS+Q5
Xl1Hs3KGLiP3/0254ym3rfF52jmxwI3yGvlDtbXAe78uOx+JvyaFDZmgJTGKUeMY
ENpX+vS/r/yGQ98DCZVHCAXGaq+2h8DmoWQNYriXUuaIaXZiOB4t/KRT//4uB9OB
J6SnvXeq2Jh3URo9raKnHAY6UyqxucF4q49Pq+B87Uzs8pPTHn5J9tXldgAnM1VF
tImU0W9L3Vzwi+dvcJTzGWuSVDhENyQZktNyneANmaXeYh2tXZt0Ol32ZTAynRaT
fGBz1O61+fYVXpgoa0ofQT2vhByK6CuI1Bfnqv20bJKBCEFLvHbi7sqpkJeIa5CH
pzqQpXQOvs1dqCce4mkqRDdkdNEmH7/ixXwK/tQsjrBif4Zd0pKBoLwLrpg2uNKM
hQh5JBqLKAhZEMXspdEFY/kxMlNT6MDGBphSFDlRhWn1XYucwCciCvMfcGDfL2Yk
RQHZ6VkII4Gg8gDggJ2At7DOVhOtLyKWQlmSfGV0kC7Hyt/PLFPGRdzSxvUGqoly
0oXxng7Vca5ShE0CWiWc2J1VlKLbx/Hq4KLiATJQE1OKNgjKqcGb2UfNnnid/BuA
G+fvq167mkH33NAGGTQL/qb++Sy+jlpnFxkqhrfUIUXljp7qGHVD6w+ws1vd0xgL
la+dkDTncy0DrJrAwduHdUFyGuWBZKB6iXFeOKwknXCIY7cZBUwmlj3s4UKilChc
G4il9T6HUDniU594utXKebL/+OQ26FEor0JA+VrP1E8SCLmSX2l3wOoUe5CqMFoh
tLjiyTj+SSJ17C0FywR/yuBv1t22eeXroZgDP0scSGoD7wqoJGMEoZBvNK+7RMoe
CNRR82z64v/b5hedTnTJQsVDCi4cz4hChXRrpZJyekICN0W820jVO7VA/a8C5he7
zTf4cVQQ98w1NM8hxHicYSETyojIflbHrTY5VsCtlQugmawi+irboFu5V1wfAFmA
qHq9+HqdguleB62ugX5krvhUkcf65ZId0i2c9etMM2wC6xylWuQC/FAKq1NgMI29
ncdsMJo8VZHyegB4w8YAnMHoSWouu36rgaDG1ywusQPLpP4StXRzJZUPiIEAh9/A
q2nOIJD7yPsls0Ld/B6OXg5WSI6yiwd30m7/Yxf4uCjXkMq7R1A6Wvs5exJj/sHJ
SFBBOKWA5eeEEKnOrwvTsXoHqEjSfA3z8tFrbfHDa+HR92ODJ3TlG7vPVAWXVXVv
VmVr4suOY6kraWu38KPnb4yJe/nHzXTVmQ6gYKPoegtgbVfZNb0qfPz9vSbxWZut
68VvIzbc7xz8v3gYPQPzw0qGumIUjYL4jgut097j5nAeiATleDjciAlpAZ8lwXWE
cn4LFk4VD2pfUDLJcPuo41zPNavd0MiGt6JNmp2P9M58mhAayBkEWI8a8fMnt2Kl
rzj249fUBFQ1qlE2i+En8zAObuIRAmwcUnl8GJ9JNd2rmrN+F3rZFrXlfN/9bx9O
fF2DoInEgEviHid5vLf6n073ogaXAq/mPuJjkNbjOzS/mZN8Lf6jvC7EFVXeCt/j
b+w//9NiX1VNFX2wVMBn58D0jLaN2llWcOYv6Tc3Bglij9L4g2wx+/bYaO0pterT
Z3a9oJ21O1QBD5WsIav2qi/VqNzPgg4tsaoWP6Iox+tLM0vO7baH9KjHoABHHUHv
4b2sUj443C9wWvHXRwx0Mzm31xWJs/xOQG57+Lprpv0khZmhqf5ysFcqVxJZqLhr
T+3BjJXw3JpftR9YsEcWBRjT/f+kgO5n1NcKnbpwUcrZpdAbF8VqxVSn6aq0qd3x
oUQf2aXreAn5kxX/KExRZhz5PVNBClLR3bem2n6zoSpZ8V9r7pjBUj7sDoF+Zxux
zt+XaAaCBzrIbrVZMuklsmUUTjgJM//3+F/WJCn9NEFzFXK5c+l6G27DTzFjR3qt
Hr2rdoyZ+j3r4af4IxB7DWvBhzIeNz2r60adgkzXvyi78KL3nZyDPo6eo/NMWEoT
1EtcpX58pArRjGzjt1Mti1nLDRSIJI+WHYbeiE7Opxf2m9fmdFfUlJosj7IwDpbn
QKrAhEFLQHi3a6Yxf/utxE+vvvWms/55QOcelj0okMPGtHWFAwrUEGRQNPBCeYgP
q6WKzQSy/2MaRclj8CxqQv9zi+Mz0asxnOTWUU3+9cA6VbWooBfiXA0ldFDsarW2
Nkz0oyHmSX4BX94XF/JKZM/ZS5oxK98j1R1zsVPPTSzkpKpScR4tHOOS5F8YxCN6
RzzOCI7x5OxPkbkLXq7NyKCJkXhhY8OKp17QsJCaRsoflV6ujJooHQSxJqsiwMKK
iUbGX//nQT7WR3YiZyJ7o9Z6y94ECqI53ZdMD13QthiHpIZESnAGAUgyByRJ8ez9
0zxCWEpExzZo9+1TgE2/dls5CKW0fsr0FHawbY2XAp1DNvEfpg1LC6sVzSUDV+kv
5ClwBxWkCFrPI+ezNY6fyIIuKIDwvBZRvS3mZfQauTWTgv+SXeDFv04XUsq9ElbA
YexyusOsfRbAA9iabLylxVN1VwoOioUkm0n0GLBRfnTnm7ZAVq0nCa+xJOOGJlCi
A1H3pjaU1NvTkQQD17A8wE5+A7zL2yY+/lScMnkQStVHdpweMeflKhCDO6XTLoU4
Zys2Mkf8rZ7OQVTB5KU2hEM4XNgqyGjk6OciMd2fXF4UDUuov/UojvCNvq2LfRq5
+E6rK/sRbOia357IZlUGUqc2HRxw1W0ewwdMZIeNrCs+WklKAcdXeYKYsVLAJDcu
1w7PVmmaEnQX7uqHgeOAm4BzyzIUy9aAtFwxbl3ZY6JtHFzlL2aL5q0m0lM959pM
lmzactSYvL+AviZYqhcxjDEKGa7kLCyKeV7MY3D0lsCGgXsZO4fPJTF2tPKxFVSZ
SCyijuniEBqrAroIN2G5Sgn94vjBtbZuk/UaQJYw0o7nihjWeVZHgHLclOXDvKmg
vm0U+R8N5lgAzAfjhpQ9IzW0fCAksADq7tc9RPAb5wfZIphT3EZ90ThiJCBNswXm
GCyedtvRfZCQZD63cQX9m2cvLRHsu4ooDszZ4D5pVZKwO3NZKQ3ggd54jp7N3RXv
UAZIKVZnLaILeK9BP3nYrnWDPOWx2ABS3hpqwwOlgWnP7mUANSib5v6E7WQRTS04
LDWyUIEoOrQVHGZPL1C9eC61hQs9cG4dxfeM5nUKiiVlIlULfeWXdrh3Afbw5Y/M
D2mBS0/Jkzy0MJ5G5EN6hrZ8uVLXUdiusC79N9gEDbKEBor9wXPCQS1NWAd5Jv+x
vuooyaFqCDuQhFjHLcM22LD8j2sfZa+Xg/450z+TLBANbSFwQ6qt51F6msrU3MFZ
gTz3q2xTqvLYxKEOE4tpUjaEhDP1KgdRSiqfV66SK6l2TdjneTBRkb3uXBcVXwMK
OXlGjsAfRDx0DG8O6W4OkOTzDkEqjxZ/EfW5GAS86vaN03m/HAh9CTyDRJr2GR8P
h1mRmxrjREyabgka7a7j9jbx9IDKOt1RLUX8fQI6eX+OI2bvE7VtG17VlzSaFD6+
D6t3s0lmmzFqaW64XYwDdUsMgI4qQOCBaFRunZjgZmgUVFnRbDgU1Icut53SkEHG
lkNenaMGyPa6QXLAW+D45gD0ERKzcCCni1uWDWyltGCInWWxxsX/G7gJbQ//ARf0
9vp/1bdOm9xyv2MqdcASdyRamFS0xYV32+0D0u3wAvGOsOUHt8zbf/guJsKGajnH
i3oQy02YDeGoH4z/SocDvy5/VZ/8R+5vjVlyuitElRBBQ6FkltZUahWDh0QlMhdk
qQDTXehorOx23qx4rVkGJmJ9LBcCUEZiY4ODZ72gNrNaNRhYdtGenyhKRdVfWAj4
nWy+1ekvUihMaYpvd98h2bm0+iouBPLUbH7BaUWF5AoLQIUC1wv9vxWc+Z0OJENf
xOjap4Tul5qgpgLzggNukXD2JOunQ0I0kzejDVMynDv6pHlI/Ekqioq5fie2VoyW
LOAk2aqFIkRXKsGSowpmOMcwSmIPQDM/IWDHtrRFmSP9wlO8vf2s1QWqtq7D8ten
27ODrUW1OcmrKv09M30fLhcVWZUsCIoo5Ooc57M+VwhSFiLbU5trRjTpp9N3daWX
2j7THdQ7Z2UUixV9oyBTAKdAww+qozVE1Md7BkvMtdZFuc92aUo7kzYIk3hfIdkZ
LZnpZVaxTgsLUeNx5qY1UlZ+rjq7Jzcr45PxoyU97r5tJwWnmIvMhYB7n+XbrYfe
WjLatvTvJgXmrMyqpRK3sTYbpUsHtLaGu1WOaMlMFKnzUsmCQ0xpF3HO9WklFXnV
+fVNrsxAu1+cG/26kIrfQPmNsBWJeYK1wX25fABRnV4SzoJHR0o1OSHcsJm3addh
3pJs2B5HrYyA9gBZiuf169Ior4oogN4cYTM0sNrFdElYjp3lK2u9NEuI0df7Qiux
rwYUegeVStMUCQLDD+CGlhJokgSCqFkDrx9dqLRwOVNyAwlDCEAimrTbrp2TzBQw
WBcSVGJJTTpIUjeJM2di7CKwpLtuLQLR4QzvC6fw6JXzaXtPeWSdz7LwGWTHHhRZ
oqcw9xAAEu3k3aKDdui3HW6iGm7nF4W/KgzT2TVaKA5aGk481NQDj40M+WJ9fdSO
K+sr5vDulkB0KEN2QMbihyB2AyI7mO8PeSkfHLqcvqjAEPoxiatxSgfzWXgKDhlD
eT8oc/xQfIP8kK9XWmt/5Omh5fjY0P9OoFlrHvsciF/+ZBRIbSvdD1VJuypYzaWw
RcEvi/zvmaFctE+1tIhFrU206MAs8hLFhclPTajDahsgeU1/QZEX3fAnkEfNd4sT
xTQkw0S3ESLcJTZtUwmJiSfy+MI8DJblidTtBj1I0yWjSfRUvEnldJ2jcLT5XLIM
WO8XfNqPRxbAlHiIVn4NH/b6raLpWb8eLmxlvnxZL95cBygpKxbTvjuP5KaiH6NH
B7AHqkF09KlhJtaQ7dxXqVWlnHLIL1B6oYxp6Vr5thn9TCOM8khr3r6+BQwb/8SH
J/8NpYTh3Y6bSp1MLOOEjcggqQDL4SqzUo5eUw2smlje23cnUUHWTYAX9SUlgqBn
fHSyeD4nqaD3zB1+ROz3qPer4wtVCPsvMLSFiuCvem5B1SJnhHANHIkaheSkmSo/
Afjkjpq9hJ4Q2S4NLkH1m/zlQZRZdYTVCx4OwQc5l/88ggbL1I1Cj6huqAOq9NKM
4zv5W9A6Q7+JH7ODl2VWf5w3Yf7UiKo3kNVxnlBwS/p86PaBu0GlB36YVI+G94ff
mp5DNtkB1Qqprn1VsNoXxyT+Gm2vK1O03GELiXHIhNbxkTymjzUjoVh55W9ZTBDs
gtU2JjdwVISW9zVmKcglkv3xJeMJ1Z6MFU+cSRzXcKmD5ExZgJxQiV6FTAfuYAME
KJb0VlVYPkNB/Q5LAY1ySCl4L5N4RQeVz90e42ZZDBhbaHyJIvtkxPbkvNiILmYA
bMxz1LpPeuLXAxPtTEujlvkf+rkA3RrXBXpbAbj8eL4jM6V1NAVPW/dFMt2YQfPz
8CRzDa46zPhg387a2QJ21DvE8UiFGuexKw0GZvsUXDILyQxUokHkZCsOzrLpvapq
Ufv/gWzIXsSncHY6l8qw5mBh3JiMZ5a4agnV0791T7AscNv06JMZltjX5kQflimz
lsihfvRLi5VWM6JMpL5B5GMDXfMvMfeF5RdHd3IumoHEB1U5q9rv+Z6t5/xdPpBo
tyPDh3gOOeG+61BY+TLRb1SxK84XFywAtBWKF53FDs9qR1Qq6f0HK696a5/4TSJi
sdGH9nVBS0nyoFlCC/Mp6ZAvUG4kC+VRlViKmzmBp/FiJ/NW54Pm5T2dIcs8ocG+
b+K1WXJLucmTUUpjXuQgoWmeYKPbyHJSJAL35lBxZsE4hqzGzYNJ6LRnbHu9Fqra
6YAoIX7q/0lhZOTviX0sTl+1vgta1sJfOVecTgw521kzOx8Ma2wBPz6tnygNiiHZ
IqJ/ZfoNnSPwrp2XBmj7vPi5fjuoPdMoYsOgxLfjkTqcS79Elp9sbqJICKjha/LU
IzDIxdrfgcAoZMB2lf11B0kfCOdvmyAk3TVv+3LGDLvcYqup664sJ4ZLFoc/5/qZ
ctf4BlNtBcyw2czFPjf1JV7uCdFodJA6eHsxVTGOXP58+bPB8e4SQyv6BmhwWX3B
eXwj56/r1e+xOWZIx3b5Thz6zA/8Qdi8LasSr1HMuArRXyjGOzb1zcapX+o+blAU
NX9r3Dxb3ZQ4GmPk5KLtBbm/TzTY2UUZM2rZDcih0UuEXpGnFpd/sfQlekA8elba
G5JS1yBHLxfCYoFe2PxXoCVneMcieABvw7QxnkeceGWOk00Q9n9Tfunjnun5mTMY
ly6f6KOJoX2hXvlUcijz3DcBz1kCI30KI4FuXghdzosXFqbEyUiYZBe8ybe2XqBl
DFUSkYBkrFiMGxawOamNvNjNjjdmSGuqpV+vWHhnyUZWc5P+m9FuupPIBtAeUVKh
xJWk7/zzSZOwjc3lJutzAwgcr45Bcxjo5IF+5S4WT0i2Y5uRpQbZpTtdhaTScP4F
Ip0raeFe5rXtt4wGcmuSQ3aDqp7R/9cFCE0QlJJiWWXDZ3F6te6DyjvHWt/Tmj5b
SS1iWz+CRJqKPczKrrP1JbiDbLamw3Vi5oOgXlECiwe3KKw1IqhYznWBUal19DIf
OXP9Loct3P3/FmUc0oRHo/I615MCmJlTxsqoZ02cPimUbgJQp47geYt4e10z9c6J
QUm+owG0YnUf6Lp07b0XH8NvQEI00GKYVVMXANfPVisp6zd7jwsmZNa5XzzW9Xyf
0ZtqWmyTIrnVgheIv/DJfxOd+8TGgUDUy+4MZrHMEQ84xGD29WAcMq+cpinZqwOk
682/Z1R0FZkpSe02jNm+cRff1QgJdHnbipxkVdRkFD7fV067M5pjWrKNJfehrAbB
XaqgCgDlkaI2KadFemnxLyeig1zbr/X21SnGs/s1g40yzD4uaGE15Ok4lskhMh+c
ZAVpf4YCkKS1qXrg5AOogOjcdxtItf3L6RYgLp4NYQhFSG0F8E32NP8izzreaO51
qhBjYuz4Vi1lbq8ZXgNAKx/scYaXCggbml0rEHRaqjRnxzaFBHKJ6hrpnfLquuLp
AjRChm1uNTmN7T8cTLMJ5kObn+3youkLujgN4Dvt+vYVJ364VD0moCykl8URtTdR
I1k7fvxf/B9YylW7qD63RDLhdvQHdvTshMkDx3A3raWWmVa31+S49sMVW0F9QtMO
spnq6Qi8cDrOGpw75fyt9Asjhl1Lxrtp4kh4nDCdHEBiespcfK6O5k6OM5156skM
9hQAmgoZRB5haSRFxXtvu0yOjr2+exxkHwL4AImRJyC+HbC4MGN/iJIrOfR0VaaI
lGa9ydaUMwg8l6D2TA2sLr56ik+9BFFI9yG+mt/wbCrEo+RYDNVt+a2RfFM6wxQo
78H9qsoAMT/Nytr4TkeiSVBi6EhVQREzM3NHPstaiaOmqhVR8j4GFCXobUbTpcZq
lecJkzKKEiLG/NPXkhKaxk+mraLnpVLM2bhw07fkdiT7XlSBz3aeKNfowfkWMJxK
7Blnpq3smF5q1cdiEMk//67L61DDcalpJlwKlbNf66VGvQKyBLLX9EGOId7c6faE
a/cZ3E7Bhjsts1AAZONQSxdsjLECEKiMOsmL3dMoEmlycY2+alyC93a5pcag40NH
3pDOCS8pyowkPAvvWHR6FVanFMLmpp2sVoXki+UEHq4GJKNBWYjRo36MbuZZrDYe
WJoxBddMYuBqrHUQnlV89ohaL4EgFvRIwsnYjLWCUmm4ac7WBgmBQjNhBBRlOD1E
smhFy5D3vh9Zj5EOyrLuW1BuSWP9bRLMpPrAhTHNwiLFGLxFbIWjJqNmhB/JHsTe
qsMlLRG32jqMYgiiF8lNTcUoK6QEZETQaYAFv5XSgYlf55uZbVI5Z/L0krbBLqWh
4V3679bmUwkbf5ct1dtRL/1+p/CfOoFiC9ntSJm74WMpUw6AUV/zaihvs5PcNEQm
JjeCVOrW1kFvMizxLtwUTR9ffm6mW8IimzWTLHbjMJ3UQbWoTMSpysRIgPehWzCN
xuXn6F9IWbuA1NuebgJODN/GO+9+Cwt6sjM+46ciMi83RAzLc39s5U/dWAgx7X3a
etO++b0Wpnv5yfAtkBSk5GijFGaY8NJ2CCxeQ6uHHLplgVbWlgbbnZu3mSQAiG28
edimUn0fEjmij93yk+cB9LBY5zk/NEJpa/GYmN3YS3v4Zejr43WRBgMzG2BuhiD0
tR729gOTu7tPmYHDfwLaQ5M+zhozkR2YmhUjq41Tg2AklKAYuBUzG7oGuubZbtbN
8up4Du1YExwapYYioRjVlsUE6TYEaZPt2LyedU5E2C4cQxGOISQVKB/97KxUTP6K
d80dPMwQbg7/AIjb+WsBm1YMKJPcpHNhwLSh+Jzk4xkGpR06Flsfj7TfzwUkAhSS
Ejx+7Hs5QiK8G0+p3LAWEKbkz8yZLhBYEf1bPvtwKbuyRwWtGFtUsHuPwi/tTnNJ
kuOqCp4fzSvF6MUCMBLaYgLzAlt2Ji/Jg9caNSugL4Um1Cq5IQ2ibkhLusggBc9g
El8DdSHbkyz9MafvXhgLHXh5t0Cc+Y6WyuY4yK8ZHofvZvufRP322hp5q0qx3dB4
ekBdvhhFIDOVH3ObnmOXGezwk9TEUxhWNqAEv4I2JwNmnOaXGhmCBFbXo0azRoo6
FqIOhTOdsXwgKq12lM6ymZpJ+SeglbEBvZeMrp85Ag6QB/aOIKzEw532dgqP/Tb3
HA96ENTlD8rPWqMS9BAtuRfY8cQpbnE6AjnOAmu6yUQGc8fJ4vi1zydyWO748p9b
ls+PsJYlP+U8IoVOG8a3/bxFWCQgwk8rtOEiaFtRwl2DX3ZQGVM8dZr8FhwiyDd3
Xg2t/+bUgE9CmFvNEsqPjpIYIMq8DLEYBGveNfNYV3nEroIEOb1LpCYvbNamQeTU
cmszaei1gT+nGiwGYjXWInD3Erb4qkhSYiM/uS2xJ8Apm1OVxmIyey2utSBOb0lT
IQvL+znw5tSA5sfFUNS3N3RRaGxq+mXRDm+R6rVjl68W0KJNMyBuObQMMn0Zfsx+
6ZlrQbDmmisuj27QChO933eu1vqubF6Nk8RQhdrpp0eBmZu3dTQ5e7rrANFlaxWc
Y7F61AUgQMBV5jkyOO4d7uO1nFGZqdKs41/9dzSuRld/oPk6hzzi+EMJvKmcuhJz
16DM1ziunP2BQlxAQk7HNSJXNGzs8mkgsJjNvFjM3mse8ohkXSNy5DPoDRpvwHjn
4gxATcMahSonyW+2IWFR7EFiHuppOUA65uDPflfiGh3o0WO9fHxf3whPXKUwHibe
c2mTC/MOMB2YEI6P2qF4C55ruXLZq+tGGj2NbhmzJ41hnfXkXD4jsbxIJh1kQdhf
DQyafqudfPp+2MCGnFp0G/s2ssvQrVTpdQX8+f7P10k/Y6CApXnCRcx2/kXHqcBE
YYrR0Fk7A8I39+9AZY8bD6BjcTXm9iBZZ19pKVMc4u9u6sh8ubQfXqL3nbYXTroh
wpxk4R7i1RHglfUBOHRmv1IHsyk0X6m+nEGuCAJUoo4USA1XiQpJb7tpfU2pvxiI
N/cnTOclmRIgWkIrgZbSQGFu0HkpqsKLa+S25MAghsOZdiWnf/gk9hBQzj7212TX
QNzTRt7ln/I47Upu+6JkmPpwh7Mk4QoeNRiJbbdsBr0CH0ggnLL3+LJFIrEZ7bgw
XT0gUXvL4zEy2+33G7mPNdN7Paxah96W0GS31OZT58Ex7dhOY54fY5s6O2lfHyBk
3jLy7aTbCb1W/Y2W3BehIDdUz2OOORphKVy0qM/d0XzALCNgWURk55uGJ7hzFlB6
KXlYb4msid3dKnw+/Hzg6aV15WSmt8q7OWFrsSeiTh3QJDcHG6G/Vsl8z+zVsUxs
LGiu/PMebovBOpgRtMPRJsvcA3qUpNieSbXRuQPg/QyD69oSbsVBH+07LKpjIgF9
p71B/+fnWdxAFoHWezKRb3yJIZHjchH7wmdwl99Joz8PsPS8IfezzWvaRAM2Bbvn
kXymRHnTV5A65aemEdjxlB2INiwM+9q/m5qyV4VRu16q6XT3xBi3ZAWRRGLiMf8a
vlQvLR/xEEc93y97dLGXh5Lmf6Pac7TAymP9D7GxeL8F9lwP7LGQjljySQlJwAF3
7XmHCTmDjhnBbVqlO6+oSiaDqOT/aKuQQQq62JK9S/vhA3vc5uczdMsAeeMhLVX4
oZ9L75Xn1oCTE9ZQOAm0w8jo+QJo/p9X97SzKIlRc0ljuUsR6sE/JpbhZsfcOYd2
cxxarNsHM+ou1tvIl2U/khNZKPbQaUTKi5ZqeLK+TzEjj9LsUI8gNSvvrwCQ8zGd
mD4jZQmYeQ+ou+LumuOqSjyVEeNe5boJ6J8jNB+Hz2uOCrCWaCTubosML4KtEY8F
Om+OqwuPNdCBVC6DZ5taxko8HZIo5Wsstf0vft09bmA5USN7DGXKEVlSUYhzJSLT
dLr8c37JU/NmScOceM7R/PBB9k4njFza+RwkvyTesw7AQnC0RGgBGaRf8xiIYAfO
DXw845FbgpEA8Ny+fdGosvbe//RTymwgRGcDCIJ3mLZIDHqimauF8Yftf1HWEoOw
z19QAzI4P1iQ0dBuKEpITEZEs2vBlRuXIdjVln8EBMojXviNQGZ18a4g11O44lu8
bEwcIhXghbzVDPACnz88pmUl2P8DPQOfrOs4lvsQAeK/AU2w9hd9A9pflVckVAbA
0MU2hysHOlSsfvH2Fr2bJ80q82EJa7OFdzgnEgR+4gt3jSJSmlaq2DHhqFovdUmI
ldRaa9Ralf6zTRaAvgvdVvhrXRm72QmQj3Wz8PwX33PZYty3fkbm/1SRRwIxHR75
FySHtpsGW5UDC2aLh/KoVrVQm/Uv/at2xMRJoKuYQ1r/+86G7guMF6jPIbreU0XE
d5VMFViv0UQKGfhCXQFoqHJYLUVVaS+1BunGtAp0SBoNB5PS0xSOtByewXrh/0ZT
bgyMj5LXTxpOIIEcB93SKDwbmPj/xf/jXn35iR1s5w22aEUSWdrA7aUrc5ysdkVi
o0737P7Xges5gpwvf86HOfG8NJfgLj//h3e9oFHu1yre/fHUT65c+CHT6C+ao+AL
IH+f7RdWFe7jffhzkxf8XxwBU170eVWwRjvhxE4HlMewjJJ+CgvxYn1fuZbbHyes
lg3iCTpppxmM9Mse2CJHZQp2cuo0IQBT/jn6w9WOOHyHNvj9BgB8e7NTJ97njjaL
pPV7M3o1AGbIz5iozko9VR1atuObVDRu4m/ozarH3L5BAjb00vgOiHVrqXbyUfnK
8JFDiCcZ83PUWdmMxrLovQrH9UMrh09zN+IDZBndGEHLUzVCTBG2+Djx6mvRSHrM
wewPgbkQy5A2FX97rqoZc4of6fS1b+C+rIsfOUOvDIOn0lX22tKwt/s6N0zzsNBk
183BquE6tn58iv0Zc9toV/MO1fZT14H6gg++SB9ii85xPdYSeEQOqIktgikrSGXT
06DT+haUp7XYlXxnR3dYnuA9HDjr+Cfy2AFXd6SIAxtA8013qnxy34SUsRBVE/0r
bGKQ3bnt+TWCCImus8Ao4hS6tZr5qdPM31d9NNPqncL9ODFguabWU8yEET7BEMjA
vkVyMFs7lcVbKsIjdzl7qdvH07mGMr/HvvlNXYQfuqTOZ8lMfvz2DiDzLEx+U13w
Aw/OP/dgQzobLSZfj18j4UjgdZ/4+JI0Ye6VsZCCOEY5y0eax8OHUty1quMJRjmR
/gWZTUqfVTHIAw15hbwlgQOADJ+VlaYv+ei//Omr5pmcSXFefpcnqsjl9BUfglyN
OQbrL7j3LGSsf3TuCarEtfieRW5vh90qQlf2LE98ZLo+bqHocFlOXCwUPG/U0Pmc
hXDFMDFpMmL8MP6fVytsO4+j+MrzroPCaTPYP84EQ4DTrHjyK9pGkFgrOHw2sjln
/J6VQfWJq348SYwqBgf1oMTs8Ybs3espZmMXBsBF3QbOesmZlyGrao6OzlhhHrZm
tMkEOx6ga1KMFNNp0IhB2+Ifis6yuE9Mt7vo9DeA8nG4l/uciUutaAUuxIS1inAe
OwS4Dx1WRMXG1dq9Ooy7MoEMWwB6AeP6lYIv6cu85ehkC8o3N+ZT5sd1zx1Rmvug
pQeDkviD3ZYWIAk9CEDNV8NeNbK++2rBwqRyte9p0MqwSBHX1x4Og1550m5cqYHs
/L3NbBEkhEdzNVT7tugapZDCoOKDo1zRpoqdY+AJJFv/jcgRXLquFURt77L75+k6
o8E/2eP0O6QoRDjn4q2qkp1nkl5KJ7oM+/Mk3+AMg/Ip3ZxjeOSZVZUz8Ka+Bssn
7vIjD4+6sbz6yfXXe/DJ2fr5TUhEbTteVb+1A0mbo64PVRcUKkKCIZLfYw0XehzV
heIzYdF4PreS17jaPK7CTi4wW2ESNoYnhWbeifDz7pPlhysdXB1l2Xn7dlaNw9wF
Il2Wv+C+dUZ/Dmf1oqQIngrfBsgwrsdqMCdR6pVZEbCqBoTqksicwa2kN26TL8mf
6dj34hARCK9Gryzyfqu6EAk/hyGJa9N11nwa1yqLMzvIUhWks5dQpqpmLtXqmc/U
BfdQS0DVNv8EgU5KnmvvVcAuHMKQz7OmmkP8ucfzNFLE5qwV8J5XouBBmah09Tdz
jOKOHRQ66b4uCEPeMMPo7w5SfHSLrE2a+RTXl5GA9cQIaO7XNjYH6Cgt+KasAK+V
fBnhpPh20rsxEjZ/3DqetEXMsd6qFUQ9gBsp/4dR84tck4x2U7TbFIH9SxRsSJKg
l3n0eu5lAoaDK4lGVaEmBJK67m4dFg5dkPnzSY9O3NPcrd3kW5nUtTZzb2bshiTV
SrtuRs0iaBSXxTNJ9XbfD/LBDQdxwcEQf9aqR+vzf4z79DuilSMolv0/zauDU5xs
hDnrITz5zJ12uaSFUG1EP0VgpjEj6MwuqypvlNDSYkdR+MmiDzaatdSw2arp8FRq
/pV+c01cWAVsF15d6XryuR3D26XfeO4CieaWjHutoyMTNmuI7kn18IWiSnZ/RzCz
C+8vcz+Oq20Bm81xvTFSlk1PiTXs54eZx5p/M01+dpR/JkS/zWB/CxSAn0xHqxTA
B0jAcNJXTWeeXgdZWrwTqlk5daxz8+H1XjhmCc9WCEdWyUXN4US+b8pFKZFI9i6X
gpfhm289848P6Yt+opRg3Ye5JRQDlWTzdty3MVnqOTNNqrdvZprNdSTQYYoSBad5
DG3/rFdnOWZO5VowaGloalhIdHsbSEEEBHDZXauABW+M+k7epjJWysYqTgHMWDGH
9bUxIJgkX2NbfonN6YxKOKHeBOLQx1tW3uFPOwbfsBztat2om9GwPplRcMg2hw6i
wLTb3chkzcnUk6GIeDnkuQ7hEG8IO1yE0CWGyaEEP+42gFwMtcIuTq4252OeTlYy
GyZS9MVZW55VJ/hPqoS1vAOhtWRqZxVUcPka4UPw4mxBIM6NQ2/HnyYINdnusC9j
V+3MmjvUbBR7V+Ty3+3LW8e+vaBE8jlvuDhcTnBO27CL/uzNVKpR6yKLageLXIZm
6dl1gZWYGy+lTvWG4x/jpokOhjsIiVSFvZmKDjTtoDV03TJ9SDi8v0Ow2NjlDRP2
KEpW2z5Erd+wUT9Td4sz/QCyYCiqgK6oJ7LmFiBrOP5oImDmXjsAwTS2lqJ6r48/
oW9noNt+J8pKx3pPyAq9EyGRvnpmxuyyjQ2MIYuVpl65J81hw9WyymakkDg6xzzo
o/OvAqJOTxMuIvKs7z1Q0/KCOhgHyYDxpNqkBzvsZwgMk6vo3yG5LC/o51sumOJc
utsh8xwqJlWV3AOsbM1pgOdcGZ7gWqhPAxMW1L9LKoXRbqDDs1PJj/5wNvbqRax8
6EZ7+7E2oAe+dTHWdb+ishKGhkemHq3cJK+z4xPoDyVKjqJ4XAw2mQrTuveSIxC7
lQhwDd+ZCfYQ7Fu99vxEf9C2BiPAzUGB3p/1ySvb3VOIDCiwa0vQ0emzV+tp0zxL
cAfjTPiuGHHmQiwu68TuoVIA66sCBdLMosNgt65LbTJ8wkU6+2V3Y4TUjW24+e5P
uN9014k4IgexE5d5rH7T/pKkOdDm7exFQOl6VOueSK8veECz4c/4fCGjY5O1out7
MoPf3HLcTI9x2YOZwNQR8tr/zUxTeHV30WQbg7oXfA+2rT2YExtA4BP13JyZxqYS
shLBcQDcSQmOVQLHIMT/nnPyDjV/ZYitzG2P1FZ49Lu8GRKdg4NZuQvssIKNgmYR
pGlmsh/9RvyZnBNAHjCJ8KOIjhU2bcYIkJYgLKSKkYkF5BWCI9yJwSDC9UnadBud
PyvYtKgX52ThBIS+L5R1wcweHndnwQxqt68DY/8ZAFejMcM5ctzk+NmSoh+Ek+aJ
5GsfIkdmX8gIiTZOgIquz4sjmUpQYPhNiBkfVdW2aV6FJZ+vU44QokvYZhmPL/GN
l0GD5fFg1aeIYDWJckrllYc5jZW0dI72VYaI7q9RKtPymgdi2H4W5EKwxjPG58w3
3g7vPyw/tH8O33hsZTF9tn24rifJO3kZ5PdFRbPOeECDcAz480QQovLzoSMsbojU
vwVpIYoTS5rB2iLiGXoX41oRw4DBuyByNlCBFdkGlELfaDivYggb+huNzaZMOr79
8yOyo8HVTS29Ea4IUBTtE4IyroliutxfALzSbFfBFLfdXxcsirkn1L+NcAQc07dp
47oQps4sQwLVRFYw1i9hoOjN8UuQuoZUhB9pCV/Xd9ytvLk/2zbOJ0SNkuey/Hln
jeF9NRgAQlUavylTfuLKxQGUN2jqX8cUbrid1tVGs2A29cqVLi5OViRW6bWTKRxo
JQtr+OnkTc62/3yOqQHmjXiZC88MrbjnE/bxJDfIeuppnaRmzStnCudlIqgrhpbJ
3DhWA85NWIhXtcYPFdQiHekR8x1RycC86qnbPZdxTemhSE3RpGEuf99pZaFJuKdt
wMSkh+petm6glg9l24RPsYQSDBtrFcfWo+ODIcTXShrYoCA/Kw6DdabrsjdP1O2T
0Ot7XxMlgsLqyCaRhi91vjfwUnh2SCX/tAEUGbSMax0p1AGNUM4dxladdpJ57I9A
QBqL8AdYnFFTR0yJ41vh9tu01/QFSE4hZZVKA2ktuDaHX3CBY48aLnFLoDCbCCMP
gghT3xg6k/6GlKuF66ErVPMwMnt4V22vMCERR+J6JYd5ZMiE56HRLt+0CxM5C433
stJknXZnA3LrKFpCHfyT2Ou6jQ+J820LzP+KIiZR9jab508MqpbcUtyGS2u9ObfD
NkvIuh0unMYIZ9ER5W2FOm+yWw36Hx+964gmnwZV18Q5a3sVSPx09X79eUo3fJ1q
pC04UZTZIDJbyc9GPlqN6PPDrG3IUpdfZSIUUSGkUgZld2WGBjgrMUHWNJnxqBDL
QLedx60Ae6vKNKPOj/BfGeg/xlAuERuygd4akkL6ZGfrNi2xfmtV8xJGlgeH74Bv
mBvN+jdcLPAvD5HYREgG+EVEV4luJScv5p5imizCvgcSc5PvayZ2kF6PcNvghLvZ
XSjjtYnKBNlA+Q+zGqNl1hJ/BnKjjnwG6hyJuAe+ZN+KhGMOeE/bNMMed8avomhW
5gShTKP3wFMW1QGtZlHB9/kcYUMK9WWrMqLdKPJfqGcSvrWSr/bAkX6KC3uTcoTw
3Hb3i1YxyQ+pd+q494f6QfDT7tSQhBtIxebltM+g8yEaME9R0qEKDOBj28nfyfgJ
7073eDq2yH1m1Jk1KgYjtQeEEBpYQ7QQg+ZCGgj7xOIsLkd1273JO/nhvCq7c3Oa
joNNU4bSPw2nx+VCQgj97wiwewo2zJnmTWXoDVUp5GSRbh9xaxBZ95PhvI6qMNVM
2JPg/Ns/9scohri2+GdRBGBs96GP//OOBL2wQoKXv5NcOENLYvIq+lvHapTFKjV6
8tsdj4EbnsyVjGl65h1hly04ZCSVYxY5tH2xdYxPIwezYKvl1DMGqU2EgpjNMSGE
sq2s8yaqLM2z/XoDsuo4M74ZZjXqPBWANWEgMVx+8YFkJc74OsjJ/xBNisLMtP/7
qXC+wWWw/k8e9ia3tYy6mlTzxhWXHcQtKWFM4+sOwJ1+/nFeO7xnegzIuEB5EXK5
gO1PIpwIvjJwB30fwr49rb3hoNNdli2UYsLWUxf62QAUsG/tZhvmL2t23mUffwth
VWmsxW+3gKVsLGqIdj7O/tRBJdnOj4uwy/Thd3Q2NGj+oAz0CDzKRuJHOh2rR3Ve
rspeDGcLRTy/Vybd4mXWjQME7bhPcOK7VX0TIShbeElF6ZZNn05ReNblwZBB1i7+
ZQZ7Dg2nkzH9McpBDC+sq9ykO5SyxI2KfOVT8yZPq8B4FbfSRVOFKh/zln1fchU5
9BcsVP8E8CCh/Or0Wuu1jULhF5nbT2puRgVpyIyTl1AphuoQWSCEuHoxDjtWKHUo
YHq/a4dr/5I7uwxpx3RttFnT8HdIVOMk5SeohiwvuMFkqLa9Znkar8ef601bcKcJ
SOOQo/XHUUNgLeKWO+Y11NGV1iHSYE3WejwxJFbNGfzCnDtuzYhbn94hvYfKLPZ8
OJ68/1JQcppWi7TRrVJFfeDc+iGXILcrjrlsW18trxJ+1VJeNTyrzke0YsvGcRv8
WZqMKeCpoi8Lb2QAZu5dEyeRdwRmuvWb0D9VxdJHnjWuOAMQNyIWGy92HNeypg9Q
CMXFrSnWwpV1orWle0fAXaRQouvhLh22B+uJLR2I/bQ6Oe1jXLeMRhvu3ITnXE6O
iwY/KsQJlCfviDqLYyS2e1VYXiDQMgwIyDfu4Q2wEXWDsd0fkN8B4Sbgnib5A3l1
wFLhvUNfGstuSPTP0PQ6tCxbkSih3vHcqMNWG/bRNOu124We5vf7pH5pVo+wBgzU
enlotJNWChBwFPa21i/jQY20pPb/ksOQRZfpTfZzRDPnXonVBtwZkCHcL6mJs1ck
xyIxf0hh7BRHH4g4X5xC0VQH3DWPiDfXedFz9UJ8kxPcRKeb0FCdqZhjbhWifE85
jdJRqDCaF6Dnh8USd1eW6c4lE808uN5Q03OGEdTer9CsG4U9Ub/Yj4Z7UrWrtZoI
zqdzcOxlMD5qwG/r8z2vC6HQZkZTC0/H6A23LhhuLzhToP1c9NUZepaJu7omPB6f
0lqLwsgIHuK8g+9hjzViyqgMSYPXrFUcxeXwzLGe+autRc5rzPdYgoEBRnPYCOxF
N1Y3BhUGNJ6RV75R9SNeFltSrxIN4rPjNF5bV/6v96898VaoOlhmc+BVgROEyMxL
ADYB76bjJGwSsL4RVOnwgOwX4mw2aFlAz9gv0jfzCj3L3SIscRwg7nubWw9R/9mW
OsgOl/M4QfR0aXvnV4f4LgfAO1scBFert0f7Ls66z/9QVsyczC6GMPssfPO8sswf
lkyPXUM/xa10+mu3DQ5Uqg8HLwOU6saU41L7jGQAAwSoiCIGVsgTbcCmyYmKOHGR
D/UMjBHxryVPapPdtQOjFkpMsAI7iNcmKDW8TKEnC+fESmML/0AxiS9qpVDeLPkI
pTIhOq160AIfoD/ddE5+dGq0l7dRL0dbW/g9dbEnr7z7wCwEn/Pc9qRMPixW3R/O
y8l5ntrlRkbrSTlh93/jD4PdYuJWkjA0JPyJ/kI6y4osri96OPJzokOCed8cxRpA
b9HdkinCZTB/fD1I8fFNWSj0HVGhFmaRLeyLX6ZpbQLPphUn2AUzUN6AJTp/8bAX
GFcCK2MwAIfEZCyRoKrAHcbP9Fy97QSJveUDi3HtlQzM4oj0aqy5OuHH/HZEcXrQ
CvX88wGM60S5L2vfC4baP2fm5/N/A4bdcVApOm8Hq/2iISUzSyvaUfZDk6Cw1IQz
LKbWgwBXvaG883g8mJDLveH3z8vXHUr856aPNWqzpmEywnSNGGf2ZxdgE1yBD98T
2SGxykJ8Xk5ue89C+QqP93DhvihWckd/nOB5V+ZdPdaHzkBRV1jyHnpVTiwdbxIL
yCmdEs2S3IxRhVz2MHW8XSXJ8sjNNX/DV08Q6i7KxHfORQSGIK63HsAp0Sm3yZ7L
UZ3D9Uep/iftMhNqjizSN3q8pMLHPV6rrPWRWhykHaU4ztn/MwTNGkcjx55AvneF
lA5DQ/rcfTqkEKJFKQdXWqxJ9SWmkmf4MgY2g4R/gu1AbHQDc0N3caxFf8sMp0GC
k3g0BuQrXZda68DKO8PxumavCbn0Ya343yHnMMq+7LRBpqykLtx8g4sNd47fB6KX
rQ8B/WpYlFV0hLLa2zBqlMNZEd1H2x+I88TF1f/FvrSpSm5LnLkNn9wKFOeQ4kNN
Nxu8cp9EcRtHqbiViUvxsUxEMjeaM6+Rsn3GYuO8ckzVn5xf0VqDSMi1zX/93rvB
GUdxvLJ4cEOV7AUFFtPGK8i6sWMZLZgWXPIC6raXexKL1cp/UBR1C53tvMB8EFTq
+rd2NjOAEVAXhyZFbZzaJ4bZJ78R784cQ8ddW+FlUarNhcXZSxzqwRWAdyoNgbFh
F6lXCF7BvOp6OLD6KawICXmoK/ovTOeuABA/27M7xmU4Nh0GsIj138Z7NKvGjZNT
rAMwP8qME2e/TtOYaOKVWg9o1JKppg8vxgwaNaORCzPuCg5bfJWjMWgbEutRx0AM
mFPuaHy7rGmSeLM/qHPfkkc476uScDHM7D8YcZOqBGgKB+K+IDx5YyJpjmx2MkcN
0sdVw09TdaCZsm+3PzxaqrJWvsbjvSBCYn5hUiMfTV+D3kjJKYQlV9ozDMValPou
6tG9cIg0smd+D109K6di9suaykerCMiZRe5sGbGmLSRmDlXIt55TRfl1TFCCJPW9
uKmrx/RLMx/zge0zKO4IpbXTducCf/JRc2Q4u+EGdO78aMH8QKdbt1r7E6dMGkQT
9i0O7tb8Dlv09tbIQy4mXUdZQsau6yU4dNWfFaKDFmW1MV9tstcCyq5BVtje4dI7
iGs2/zckdzTbPJt+U/yXE045uelL8WtnaW89T3Vw340P9zWP3fxQNsPgzrtQM0CY
VDlOnv6je6aE1+iyPjf8QrHxLv8eseI+enCjjOkK4Nlwp/Ksbt5iZPoeupKqks4w
CYwttprcaSEKyL1HlqQfkXO7PTsZJ82D4Xe+9CZ5ztcrYpD5f3pP0q108x6sRihq
USXf+qvw/eDcNThAbB5IJs6iujqIZHMpHyFKckPWO8cO+Vna74/BvwEOwzrJxXwD
gGuHaHO12vkoH0Pck3df489rtSke5pYRJ4m6T3l5s2Pwj6sMgOrZ08wPrrZV2QKB
QDJvcbIJAQHKRf7or11KnRfeR1aXtygWS20UHcSF0qrUHqHiErqGn4BPlXwhneV8
4g67Hb0b+UI1pgIKcjqlhjBHZVD14peLUZZ5irLl1DdtltmfRCbbbeRAJw4VYhBx
07gAjUR6uYYYPU2QAxdvpfiZ00a5NNdTqUJdvF+HZ+VzLU9PrtMX4+Qp47PaYpIj
hw+OeHutRP+oh3QYBq+JQKMHVptjRGuZxZMjXgK+dO1emKo0FzGGf7Hn23R8ivGt
gMcV3dAf1FlSF17vlZNtVjI8MsOx6baYurdbDx0Vvet3/79nOVwIJsW1nF+lRaqQ
/x0YPggDvXFKP2TIDJWBTPI1c2WzcCWk7VbqWmyyaB7hKCGxha/A6TTntsSlq+LM
vWZ7LsBScgMhyrz4HtVpadBTlxJYl8z72lBf1+IW6WUxJKU3X/MT/PKR2e5ZWwCn
zpz8cjF3rLSxXzGacuDAdcUCJbRTwQ0I3KGPeSMApegQxxdbKqZtRGSQzmJWhgDQ
RVq/yx9D6bcJ4PeBCyqOpYEGeBbcxg3iPB8Dp1w9y6Z3/uDRde3iOtgmG3vNLHwY
+NL9eidbR+zsb1FpQsyoY6iS58rURh6oPaawlpQCitOjBXI1MMEhzg25PFnzh8td
xc0yzf83Yaz0PoYQf85OZjUHfnJMIV1scsR0GgrshfwZPdt0p3S9Ec54lM7+Ar49
WMDGeZcPW9le8VmhmqV1uFUmZjeaxAUnFwHdb/f5OD9Mc6aJxbs/H8KbEfGWvINF
WbAIt4DM7a7hpA6JBfwXUnr0spINeMhFisVmBvrUB7slV4s59iUFnsg31SWJQuFG
wDqp7dfJ2LNUqSNS8UCzC9H9RPBVf4kjMCg05rJlJ1fHa5xoXI28qQ5gJSm4/njp
NqbP6GJoWoWL5v8n2aMDmComuWtr3VCIx5DBHtz9DxaXCuTMRcUfOPM3lQb4S3zc
5CYBR8MCA0yVBIvaXmokn0QPboPmw9A0w3brfnJ6ap8NyUkcPUguIw2FHGGEx+1F
oh48ShnGKaNZjONb/baUEC/I/+87dCrbEZG9ghRXcmfG/PINxDA/5o90X7ji9rmD
sDgeMymOLea42T9CWu5oBPJJmdK4roFLT7sjbW2DG5CkzZ7jsuuzmLECi71q+pkJ
7Ym6q7d9NNySkxdU9H/OEDER7j7iQBxkhrge0in/zQcGTFMANYMOO75yX7rmkd1A
n3YKHI73wCYINChzgYfNBF5PLYCGhspquY2Cb62QepBinTePL3edxBBuRdb3HHFP
VfL8+jyloGgvtyuy5HfNvu72KTzUpAZ8K4/D3Y+4WLFkL4z86h8BhHzoazJeIEEx
4zp8KocPj0JEOcYfu89+sucISC4tjQYVQxiV7AfCdIMITWz04V8woy6QsAOZG3LM
nanuiz87kKtftneYicvPPChjG1LIs85j4BFTWSo8BxmtlNTwzkhVIasvVBm+5zkt
3qden02Wra/48VKQYFQAfYf9L+uW7ZGQ0OO0cZsvnsVWjebZdMO8HFYsqc0gk11K
aDLPeK/MKFSHurYtVOWvEHw5fGhnVFSD37t27qsq/D8vs4paY7fYAm7fL2/IMIGB
GwJjNOUHbD8tRA/nlsL0GceTlY9g7Q0m4PqucI1NQRewjbM5cW/FBblnOvpk87fl
vKGWI+ya3yMFjaB77VObBqD9eiOOK3cyb2NGB5YJmfEvw1wxji+T2gyBtfsWjEzu
N/sE8tu+KznJ5rx3Emx+Uzh4sjYj2odUZbc05ViMlWSsbBKK2nyWKut7gzIKaAFi
XyayXD4jpJcolpnlbGTuSG5KofjCEleOst6SNVYyOKVxQv9yipzEK2h5POpBxhFr
B10s/WEni1vlUWQDyN8gXnTFhfR905PVbmbfBL02FCr1nqx1hkbBULO99EcRHKGN
q9TLD95XFM6E0lMoU2EeyRS/tDHja109Wapw/lZRidXRjwhT0+2KWEZKlo75ZoMp
C5VXL+lFbB9Q5hQQaWsrHWzpO01Cnb0TgiHzVa54OU2xcZGYGRRyErFoDLrmQrfW
bb7Uq20UpShfjR+8sY5sXkXBDenfCGr8+e+c7LT086a1+8zLC4clexENFfohnRLp
RCQ0BL2b2YBVrjjlvPi962LIUM2YvAlRSxQjyjq7otKk5alJmn0nAExUzl8B6VlQ
3IiZD95G0T976ffRO5QW+aCZekUxyu+sPPY7rLCSJjdQt/2VGGDzLKgdR1NR95HM
F7TnE7ojWL5lKLHvelOCPqo9QaajQplUFRUzMwXJCOCXzdEZLJ8CDP2ZlBqcbl1o
pIxgjQnom2i8gY/LIOITz63QFcOeu4ZAdWw/XU3GnCR+KGAmNI9jK/H8+WmOxUtS
tTcaFOc0ihmXXWuO+5OIbbxpSOIIfTEY6LC3+2Hpu+YVF++jzXNS9VoW52x/wbPX
TNs+BFmTWSnY4MxeEz4nCqJoTZp3Y13ZVWqAznWIHFP1KjnkN8GXrFtwWgxND/l3
HB7f+PpoQq/P/7XVcCgHcTB4uxF7y8tmxYFP+DSQwvzGvPDA8Tfn9sQCihO/FnGH
u6C1YPhRZC+VTG1mP/+80WCSs3Xl0LkV4X2tapUDPekrHFVnuR0aLC2R04P7/yV5
Rd0ufQc4ov4ISKldWjD5XgBtYmP/bShXCGovibX56c4dyjXAqC0EpqXQQkyKv5C7
1PJ5DX0e5QuKPqoJQGZoPhDs/0erJ4cUa1+pYZ743bD9l889723Ra3aVf1HMT6Ef
x3bYpbDtC2svkCPnIbdffCAOddnA8EcGRsQeZi8eYgIoHrrzqKDywgpuEYOJAIm5
aKRnXTRCN1NHOJzrZ2uueZXp2pHvE2TX35qaIo/XoCgA0NYfCf6CvGTy2I5Qy3SE
kWTNrt1MX6qBPk4UYsnxfWOgnmmwwzD1Pc54G0OqvnLE8Wa3SXJF5tNvVfd2tLwC
XfufQz84za62MDEMOFBMWhX24hxclsS3bEOTHySuzo0mg+uHYw48g+2xPtig8phy
dVs5rrPibn7eaAq/qORvMaknlLAxdWmzEL7kHoFRep8VBknH6NDAeE4kA3graEMt
28T1XtPbQfgnDYLExZgfsrcGlYIdxcmus3ajOFfj6XdShwe6Il4VWvzNQMnNQJRv
/ZVcEHlDEjhLwYs3s8Fm6spdy4rJhoYoVscuijLbeqahUP8SAGkTBHzZ3G4joZD0
Cf/LIQiHF1jhoLBy8kmAgX/GFdXBuZXRWWzLrRhgoKO89pUFx0QLuMPQY0J0at6l
lkjEZhkmxOcw4wSWjRjjAzHpzrGiadawmDWPgIfcbcsrcRc5KCGvgmp3erln2kz7
7+lNDNmJ4N0Su/iSjMohOLPVJskJLsg5+Nki+AWCm1XXvNF6eaQHoFv2vNICBQm2
xgoXypu08jinGXAY3x6iRQZi4QvIJeWII7Bcl7LbNcC7JW4sa35DsggC+C/Hy9Jd
1HPSjpjXvwnOcClV2cngBNIG2rN4Bhcc2yx55apO5s4IDiDhsmoFC5lRC3gPe6K+
fgZk89mm7ThAW2L1WQeKwbkPx0/nVtdaBmSzBD055h9ZrZWrV1tX5N/LiiAF6/aw
ME6JrtU9VeDrzutuE+F1iit3bZEqK5NreplqL3qvoiJgFWT2B0rXomChEkQMnTxL
csgTcei9a+riyj4kKMkSmaqpbgT9UpEnurtVS/MniSGO50B1IRZZAQvCxz2k3+p/
qE0n4I5UD7ve3a0LIWBFIYSacl3AhHTD6YyxpGcxkEBReIn7FwfV7yllguNT87NG
0TMbhnlq3V1sw7H6MwUsIwFV07dC2b7YJ1/8A0ha24+pENvrv4dGG+HH1EpzIlkx
6UU+a2EbdrnWSF1JIEWsMlo3qjDTJkNMsxBOmVcbSpZztnhMsoxaMHqkqdGQQ3bS
yBAc1o1i0OWEHsvXJY1vl1k/wJwNImx8pUIqcnOjPcMfc2Ebjz5EW7pU2nOZAu8U
GIpEVULzI7jDAe8TfiJzela2rvD1LpxxhggqNeEgC5eIk1xrMe9fewUx/is57ETU
mNpCOAm8SDvFRAPvuVpKT0yt0KmayjmZejzZt80shYbDnL/ysQFd2FphL6Y0JzEe
RWTEicG17/Uw2b9rxCFu42iOxUCRHKANLqgymTuUhxHm+uv9MAR6dqIMeac4KcFO
BB0im09XiVl589M8d+d+QEGXIbOaay3ltnH9PbHSldWqw++4LzmRO7iFKgwPcdKW
hiqFnx5goZtfQG+JqymneOQX4TDy7Hk9PLSR2xN+F4vbsr6Gaou9PlefTS6+rfcp
PvRu0c5sLs2ADvsxT1G3FzmNeX1+GdTlj/Sv4GtQSCvSPQ2Qk2tFF/a4RYfV8uPf
KYTA2i3uq8sS+9y0HtL+DcAANUiDYRCKc5q55HkFAnuXVOKYXgdtj6FnbE7ysq61
RVBWg6js6rSE7wuzXfThlU3CrpEzSW0KE29+obF8ETKPumxnNtNFksxRso+pKEUM
9M/945srWTKGvOe68XvevGsJmtuepRyXiiLL87LNZTkwuzgS0Id2Iii6bz15+Tdy
S+g3I9RvrSEE1NyEwnHeXKESNn9uioswN0D4H7gVUUe3gtBpZ1arS4YPnd+vLmRH
66I9pKu8J8m8IGBJPi+30nWY7CfAKwzLIkguzMSAct3d3yOF7IZfdt5J0Q70Dm5N
Np5Jwa0Iudxa8DSfR1XovV6KQXQa33HEcJftUWTjIRHIQOZSeMKP9iyJJbpWFWVG
OIOZYbmaFlD8QsumEVmKepfP9JcpbZDLkHmRl9lJQNAsSAiXiYo6IGleinwVmvKc
VMM16xtxILV/bixs3v2fDsODHFwxQVpsMJKABdGOtnkO/wZ//PokT4TuZqJZDBPT
XnA7oLE2Bm/BFxgkWHnBKp4z9KhTVA48MXGkRa8g97wiVXFVjcf/IXH4EEvwC2+f
mNgF1nLuEpq+brd/6lTzjrd9K9e/Fbb0XnVU8ZqTkL0CyGsXOcaEud+VzaCRPuO8
lL1R7w7YDWPoLyWCr+Dk0ShfwRtgcch5JPrGyTSfT4TGccTC0OZSUrtezC4y7dLM
lEP6shZbJi8MVkTvnDcJ8Z97Qp4WNViDoeby8IIJ0r9ZKCX27W4/yBDu39l3lB3Z
jQya+xWLyj+i/BM9ER6eP1lb/gY4JXyHOwfCwqSD/auKAuC+oDpBAXVG9s12cOb8
AqnaluI5OxSfEkeCsu/N9E2vIg0Jq8j0sXHWh0seSjqDAZYZjKkstHbOU1UV+B7P
JZaFLz8juQpxxgQqBbwI01l5fUwuGo6b8Cnq2VwXjh5UbioEpzUUeornpt2mPngF
YTeRyXdbS53FeqzPlOInXjv1ZeSkBIF7fhyXb4UDjb13wnXQmw1BU+p6cWpZnE4z
QzmDQ8d8blO2A4H4mn1Vj+CBm6JJj3wH5kuPb6LJBq7jlAr38sweSLmbeIxk5cC+
X0rPSPN7cl0Dl9u8cCLOv3k11VdkZoSN3OOLKzkLFf4QPzixVpxuendURp4HGj2P
wpSyGVrWXsjPPdugMtMTHGOGgZxXNbyqxERmpUTciEZBETg2YWpZhbcyDrLeuBOl
CtThZdAs4ry4aQVMffLLAOsPv1xnIbRWV+trFF7JJwi0iy03C7lDKp+dkoUhdpMp
DuJtV2gqEK26Sn0TlXMgcAeNErCvzdpbTP4IsRQnAMN6HBXBDtBYWipDKKKvUxd9
EhToSrLEb8S2bZPfS/0RdfV+sGArMModtd+Alat9c9kJdcKZeO3ByEaD2WYKH+UD
nTRc7yrjM/PMapX2Bw8iqhpKfjLEFTF7y11sDUuc3AHpuSwMw0dymrqNE7j1FEcs
S9SC2ndI7rtaXL3PRaSdx0J9v58cfz8GTVEBbKF23fIQxmYhumlx+cZrs96IIaU7
DiqaguQn5CmrL/0G7IFxKlNhp+PydhxCqAMpJKBPQYWHF28EKoeJGQFRHO0cyKMK
fFzovVARV22ex4posQSwnSrdp4zOiCgnPKdWrxrhIu+T378PPS1Fo9/Vlo56X1YB
+ctnvBg9TI7hAdjNac1YPO8/fSjUiNSthG+S0ehQ32bBlz4gsYzEBodeyEDkCg/0
VR7XINTaP0YkE26Yxed5uKMtRRFrrxVHl0VXoPctZ4ZIY6YtOJqf1omyfGKlmUce
fbWYM2Hoy7EZnxfcEFHwIJ+xEMs3FoMhZl2Oln0gy+74T/FQPdXbwTyl1zslixPV
FKCAbx86DytliqeOZck99GK0KaLpgCG3vnyH7TFHbND+o0S6O41/66QdhFzK4og+
qVYaWPd3OuYxkxTeRJ0sbrYAiBEtYr+wQNzf8X33krNlIBhBe1m2B1USs100rGIn
Wy2mC+nv5nRUG+JM0slqrbcK7LMuGPnet6DzhI6w0/1CUesi+FYbjlcztTji7DdO
qM/SnhI0pj8B1/jsfDDQhFLbcSiQehqxd9grqK4IqB3mTlfQf98YTWs+GQ09EwVS
YTLRCaGQ8MJCvMHBsP/T4PpJg0qk5bPdGpYyj3VqJZkI5Ycyvg5RJbZMwT31Is6f
S8olhRvy6BKmgWa5FBw0Tm+9vWyETJJoU8Yt0pV4AHYaQILzsvg3srb3NRoS923R
YNkLbuXgZcg9fBazoINe1XUkzkGZi7LvSI27oX/OoD+6x3D977sjkn1FmSv3lbOZ
XzgEX36YmyQrxui+ssaXQdA3avRtie1ApvHaMssrHfbpRf/v54Y8eyEPoK+2eHLQ
gJt4u07RX0SChMHoH2/7O8ozlm4xHiF3qd8HSlDKxPF276augu/YCrERV50G7afp
+EmlZVp+dxHboIiKmC5lcWmJ2UFJ0C3X/XzTGA3PwZTz3hNTOfRIHXTM33PooAyu
0Y+1BwdYmCEEWGAxpsLlwrysVxTSFVZ8xFvCCuyjcUv4QCNqmj7YIbqKPwn3BUqE
DoMcvNwTVobpBscfjfjVj/9O+i2pCI+CUdd5zbcqaSxwwnh/2UlVExzTbvIcB6EK
nxdLU4p822UcXwJGSf7q0g1ImcEuZX47ionH8c14NqPWJuS91MmoW4KMKBSZIujr
ttbZY9M7HiJRF4p1bC28+cxjSHsp/OePZD2HkvtT2Rejskss+D6UTSkvtcksskmR
eAV8d1SvjPNoWU2ZZJC2PPElu3nXkFximFXHlN/PnkgeTsI30n/+soyz2qaC6qsj
L4l9vgLEtFGvyHYyphvIZM5muXhOnfcPZIS7aGJvR47eRDk8zQlb9AqWYBtGPVhm
hwVnvXkln2h9wDMVNvJMtotpaXnQ5W7FSstHgBBKz5bR2j2TBgF0TRucsASXB7VB
J6U5GcvI8POdXYpwwxJxrFUlrSxb7G+IP2blTp1jtDjB6NuL/1dTdnwO3sdkkI/T
yS3rEt7vWyF19TxL4yOl94WQX3195kkzAbUgxU1MMrEmnvCttfHkcDEUGkD1PgSD
A0Ea7twbSUekHwlKiKg08w2cmOXDoEpv6omKuMvyCoXe1rZUtQdKcHF0N2YoiqQX
gUbx8UE9W8jkC7NIYkj7PzCW1IHzd4mqjJJ3t+M+MkOvBdtOv6tn1scOs96syRAa
APZwcZQ5FWd7X/nqV1LfoaeiTj1dAXa8oCt3UeN/gpzr4NkUipqtN5axdCx6Cgl1
SfgIEkXRV/AXi1d8mpSmVPEacXpjZMdG4l076qjyEGqQh/ny5A4PwXe3t5eMTfZ2
pnjDIUOFCC06/Br0RVrBaJ7sdCwYJ9Y2UQKwwr3fxOpc8IdP+x7A0e03msXalZ7L
T1GCjBCMkGmr2NBSkOYV3CIbS6VF/LlyvbXdnFjP9AeMyUWDzxuf7CFOCtYfGCLR
BXpdJe8NM4ghsRTAtjDjZXtM4NKEN3OxrxSMlPe8JTuNruD1A2lZIHWETlus8/hn
W2ggrmYOr749pPa2yw/q31j+j3qszYF5l6ecfu6OvmdEVD8CWDd69j9GKdcsnM3Y
LkgPvsDYkNKBTXtBrM7fr8dbXJwtM3WQeHJ4p+jFcQfPUXk3jr38XAeTvIyDaAIp
fXoQedDAV0zBbqcEKGpSrLGN38gK2gORa170M2DWFXX4yRuH3NvX9NmwP4keSy0+
zzrODr+1BRV0BPJyk8zKOWaXryt52tKY1pr36j8MOH21EDNONYXDXdDjcdcq9IFX
E5CG4azhxFasBnjENcTssmrnPX2v9ks2Wz8HuYXxFufIqzYmOOH70+9pP3ZoTZoW
2dLuGcetiGUq4iqxX5pOsXN/+06yQvRQ+Qo0C3+UHHWsElyn9RJ5WA/ztDxwVhL3
+XR8BIsjwousrUQxkkvqyUN9eccLI+5jn+tbDNoSgITXi4MY81lNwIIKHIAyXySc
c4U4tve/KAOo7OP9qkgUKvpFLr7UZkg/ZYtGiGC1jw4lHXWdv0IRuvMFiS1Xte07
2VYcAkPWI4CH2hoefjkSBFZ72lH9JNck9BPrCFEb9CkaRkb/DfP9JhrGWg6rVsxT
s5r9zh9r3VWUBS4Dvke32Eq2sAyDTVWdW2S0C9xcET2A+wfL/aDHLhmeo8FO0XqK
ULdbBnl5vYtm/xwqnz2jxQJdqiiLKPeUiP58qYkPtMTLP5z3dclO/pSc3N834zAb
zv/lOVTku0v513c60nTLSTcWpDG7aTGAv+wPaNWWWS0anvFmu3/hYPbiIsvqkHcf
80UTca5zYfLwWqw1EbZyndoZQaXg7Id3c5qyAmTS4m5VK1C+QWn0oBs4R5u8GVP1
nEhi1wtM3KSG+IS3FFJaPNl6wRDPAd6zOP4YbgHwvkzpiNcEQYOHt9oQJZkk1GPN
HQUZQJ4g7sYxeaT7o5D3IoVA4gy46+Ok3a1w0hKvEnk1rbgaBGz/Pll7Pz6xqVhA
xy2Ajxnjx4TDnK6sBNKAqanK46f6es+zxgmJMx+Pr+EcP5DzfuEiz775IXdi/EvC
GB/IGmGMlhuwSA3bUILUQYCGO91TJGRPIhKAH1uYHOQHerplEYxa0wnIZ8uOcDSP
8ryU36sW5vIHTD2dBYY2v5sh+ckllUsfrhgKtx3FLfDbXSgnb5XoeSa1Tweb0b3c
/OyMT1N6ligaEpU4dsQaPQ7be/QWDykUmKeVcYDJIB9M48a+QVEB7yMtSmcYkISO
R5QfRQk3jEyCsz4ulZHL3rS6xXHFUZBxQIwyKXW6VZrREYkU54z8/XpEEyMeCl5d
LaGX9L73yfZ2O8qms0EA8yOY0zhehZSt+H/nramSbf1/Nm+3WNuDZJHvkVqcnusc
qnoyd/+SAQ8bGvc3mJViX0VLbhVVlrQzlkSlNCxIW4nwO2ueYaWVpTnasHUlhSif
Bwc9rN+Ud2JikstCoiV32dmU9rrMGJOR7qDNpGfq4wMCpVWXPKm7vkDlddxKE1uV
CiPhuz+Stlk+8IgrdMO/Mb/Zv4qWDph0+UpSg+QTBKLMYYLfCWsaX0UUDqcIIFV+
+b4QH6TunvIN/eoal69iHosNdU2IE/RV25xE17CJJ6SKgUSlOPy0tN4aInXj61vi
f66pa8VZm5LOyq+mD4kmON82jhB76UJvNWNxNHQZap4Kq6MvhGRxfJabHIwfDMf8
zM+g2kl5aTXJcoNNiyWm3K4kLNu0X5frM/tNSI4Z5RM1BDIbBwlQ1qcxrbWNt8nK
u86yx701xG9OPjgP87d0gmVHxOQ3opGnkLrZxkD/9WxT+5oCiIs7hbS6nLh4XRR6
hOIJWvYJfey6q/3vg+bDXOlrYHrb6RnOZJNFNbG5fTd26n0caAaZSpg64WH4iP5E
Dy6u5PGcLYoA7mKD70kZ18zLePC26tOEo8Z7XDVN5IXnBnv3/NJQhMD6FSQbgFQD
8O3bBTskprUrPtjuR53967+vjPuNwh8a4ymMKEpDR4w0DwcXtEd8dcJawckTePxR
K+L+FX0PjvC98Rk4/pmZj19RaX/Hyr1/cZd4+EuXegtPnlBAS699qG0EA/plvewE
GitCthD1uyyvPjIw6tQFA877G80tmOxoasr2qmkjaFDk0EtBLnxeMeoiwFKYc+wi
PWFEJEhpdJASyhiEnTAWAIM+N1tZZxUsArtD648L/cUyE1nyo/ihMZVuohckr/5Q
ZFbDS8zsheJeVcMXdPBd/pHxH8KxI98UBdO5Saq8GYSit694GxEn+PyAHmBmFi86
BiChPg6Z48LqJgHLYdtm2leB2L765OI1DrkosFFBC8Vt1SgTzxqPDqAsvfM7wqep
qw5uzaR5okztF7RDRCb5bNBbTvE6f5y2FN5UKHSzskPxowu+fxxx8qGDp1Dg4zQW
9sqNB0ZvuuW8P8U0RciXuGW3ArjQWtYNLRTs3DvtDQhFnj9mTZuS+Fk9E7PJ2yT3
Et5FedwpMXKE0BKeg+KzpGz24dICYEe3pH0voohoiHjyzb/x+mMeHdfUhyasX4MZ
1gUk9OyULfiUBs94xIWSgscBxf/g3k1X0RVc7VJQfGrJMgDZyRxDO1uh33fSsppL
BjASWlL9oy8obX6wByAvPypQOVwzwu4wJJd3OqexIH8L1/5HtK2419GiRw6IjS/U
M++Ux2lukdUPD3B3xnmg6R/Ni9mdwOyj/2N0Qou6N3DJKyFx6JW8/EghZXaejOql
1qAZmVpyusaefZiWxxQPvdPcSEKbdtbLsTEmMpqTnMiFLERJS04pgXShPOaPsP3W
9uy6D2UHp447HFDgz5lEw4ibwfvXilocobey8QacU7ah91GgIC9zcxzCgJ0nWybi
CV9Fgg4+5fqLYbEUELIkYx0UtJ+RdCNOFoshhPVZrTcax5q+S/mpZrtscJ2UY9Ia
cy/n7Zo0owTL5fcvSDo9hgD1eX6GPYDaWjzOQetQwZfrh6gCWhwPDdAO0kz/qHl4
UVMaw3bIKA6tEtflEQvWGGLIDiTG1pdO6NJM9+Tr+Uz94EE4JjiS9wBEHH5I2dU0
7HEFUaIJYBNzEWn++ieEnHFB0h0k7N+fCL9tS+XtkGXKdsGCVk34qqckql/h8J2h
+oivxr0CE/bBDiDs4RjNYDs3osdGgWOYP2lFNHHY0n2I756jU2aNs5Upl8VAewNb
omstlYIlKlaitsNUN6uBKNQqSe/1oFhEw3nZD7LMmWf/4N3/zFJCXrVzrVq0FN6C
s0ehhmGCLOr2TGTL3uIiWLHC02s/tfZe2Kvdju9ss2Jso4WzEXydA54rX5DOoZWH
b79osjmqFE/aaDzNWlJwWVGE9x1j6qwgBHtb4XyKHbh9t+caFqCqI0XgbvqUHiSf
T5XdgTDfHPuJ+dzWHbFPpx0mKYxKMywlDoMPKCAHM2vMdjrxOaY9RYgzZwKiDGgx
0rU65SEYAZR9GHDc9CrQxq+lVx6hBYiUgdYXwwHFD+GC8o53bB2WAzqDO3iYrMoL
dBW73476/by4Qk/kb0unaaB8yxMetnewchH7yO7P6fMrorilpANH55XWDSm3f5+T
XzsDdTMcIXcqUpoywPYO/IbqaC6Www3lVocYDvrOx72aPRVwQI4ABKPal0yQ8l2F
A1kjWwI5Xxi/7NNt0eZGSKhU7ThD0ZCKZBBNFxTWPBMMCGu1Hfd3MKKbyPTFn0wB
MP2P9dW3rR81JvqnQ7l8YECuNS5hV5LGuFnjul8MMkQlC97l5U073c6rAXjKKrNC
4tbnxIQ/BtPkOyo0MoV6497q/NVTvdsxwL7rYSxlbI9kYzdcLzUnZa0MNEMYTVOx
VTtOav0z5V04Wvri+18O9Tw7NKpi6C7peVh0VQ37yYGwjdxSoIXy/zcwYrctdjpB
kzpfa7PElve++VEkniHZTwO95HI1Q+kTyjCF4BsnineD9+2tQbaqECTkAldZ/Zgr
2avLRw7CqpJnuXk3mfr9ydNysHafp9Ib1I4/Ga4/PGgiq3MC4x/T59VW3f33tMDu
rAKAR5xDw2tjvlHrl7YGSQ+Zvdmr5/FUrY+pIBpfbYJgftlpHMcQ1RYEqu/i/LQk
j89kJKH7nCZqxLFAreMf4INJf8rWb+YnZxav0QprZU7vwSIBlHPxwWUwiSO+6t81
r8m3qpMIZn0bvRi5WFPS/qi2vYZYZtNMa4avYCgGcQPEuaxdKhSjNoiwlxuMd0gl
hPEo1evnSa3Uh9ZqGVO6LP+Ak0GsVHGQ8l1dlJVD++0vSVXzdZOpGvnuI9Gnp5yA
XA7mosUVHKrW4RAiww0QGNmtSpJbA6b6+dazl9BvYWb52LZFpyxTXHZ/OWYHQatQ
mmt2Y+pDHmMCajvrIoCGlpVmHlQ5dDRruBwHL68gSudGq35fifglVYuAe/DXCBvZ
Lx1P8CAwsjik0FapsB4HinD1eWWmtzfE9SR4gplvLmYgZDxNGTWrUryMANpabSg4
IS5FoGVwk/FOy3R5GaqLovYH78TWh3oO/7lJ+oNEeA1EHU5BbzIGpTidnQAj3T0M
wjz/95OEwZM4/wKiqKbmk/DhIy2l7evIHtdqSW44AjreK20ZubhXB5i90fm65Ern
jLhF/e7qvgnKIzq82OcoYUDi5qDBgSLlphcPf+dzOufL2WOegxwh4Hbypz9JZ7dx
Ku22rAcrpoTodkYpafWd9tBMmykHEKwLD2K5/57OR9Sz1cNc2B9XCs/1uGSNb3qZ
YIrWteBjRt1hFGCAS7CtHVXrrq1GVL0PdW8s9z4aMiDtY+yZQjmb8GGoLoHA6YsQ
AZftcYS5dNk6NcEDiBYxMH6jqwxfO1K/3Ihf7ksFlA7Tl/SQBD6lzPwzCx4fq2OP
6iHmjJYFypmXa5fLchoq95zvPC1oojHtGhCLloMMUtD+OFj4iJO3aJF5USldZvRY
4IYtXOEaoEX2EkWLH6QpDcMtyBtmaQX87jM8DIWhY8id73423Qg8OEXPAfqPvSmQ
IQsVeq0yVuqYENjkdrqCK3zRP9KrGS+8a+bSS4RfBx81pY3Kes2t1//HZ3t3lOYs
QfWyrLFTMw1XUXegRLkZ9yvbIFqHmwnP99t8ai/nrOYH44qq2C9aBtCAJHDq0Rsb
PyOLIq7nndX3tKv6my32pJlqOMVxeiOfDhRvqxAP0rx66vGlfn4/7xR3TN1pC9x2
cE4H5Rnl3dBeJtC4GTUAS/fbDWVX5mIX74smeA5Iy6N7ESFhaeRWG9pg9fOQAXMR
sNzydaK5wg0yUVzYCB15/aUNe6bZiwkvdGZJJnjB3HxmEP5KRITeF0CnXGByFASx
jVmfTU2XpUP0ZKGnagsBSoeLFoAXwtWU2/NssMzqGwuz6eYxgQTQXfS2ORWGzt34
7oKh3IaSiqQ52BhOIGU//o7t0H+XbBYc2naiM6cXzXPr5dwUtPsMhwY1NN/mSogl
i2wRpP8jUngvI3AdUP4HOxMfRfZl/mghPNkpXbUphsZz8aIXoxVPB5ncOspgjytm
6XAoSizpBAXWzo/r18L7lT2Mjtvb5kGGAwJyxUoNWzAJGZeNZH37jUIYizN/gMpv
nAsodADJ2a4OeOUbjCFtZf2wD1PVVWF+7jI8OXpLwcJhhr/JBMTSK/cKAWd03WZf
Pk+1LBhFugsCLW9HgjpHo+M86u28t27jkf3EYBYpNgxOlSiAXuNJclZjHt6kFn5p
5/t82bIeYQY3WKjvMd9YIi9KThWT/F2gqw7AjpAC9FLRTFcIHUzqYcdI+v/5CwXh
ZyGWmFYcwY2He2FabW838sPkJ/s29rd+N/8c3Zn9RvnG6kHBnVwvPuy8mXJpzGqz
hqQqALg3wknf8z/V+tR5gNi7BRuZ+zfk7nZkn6+kWX5M79cC8nsU4DTrK1/y8xwS
AX0hYT2a5xrXTGdctfjgRUm2nRXwI5kJ+tpFLTM6FqyCRXgAo2NQ6YWiQOW/bYL6
ed34GaQUDr+JnaJlmCZ30milrEDEMhKDwfEqZxduTOcYe/pahtZ37AtcoOClDnvM
cyUIFL+kxRiQQjaxMzWL3r+BaVSaByeeuDWiris8Jj0zxYJB24ZHkkVd2cKlwf8B
az4ifCijfUu/hxViKXLK5+C5Oi8KJhN6GXxwOQZoCQvyGL5q5DOC12pUJY2vxSWn
dj00IJfjcU84XIAAIyqJJrPyMm7d8y+Qjy/EKf+zvh/2uG0q6cxL4RU1L2OcoTGm
GrV6d8D0rNLNuWB96xOSQeo6cfmVgJbjm10I66wEyc8yHWd+HK5GzMo37yPYgmyZ
4UKw4lPJNnzt/UCzK/u9UJAcuAx2v7Eb0/nT2zWQnHtf1qks6Cnzj8dpUMgbYaOz
okAGqlc4hC7PB5k4JlUS1tDuQocor5RX2sSqkAV3PaSEUi3lPk7UCtPhsWVBqlNb
gz38+ynzLVw+XKCFGVQozfeuAUVH2Owda/KoM9Snb6CP15Y8/3UyHCYN4AZ/2qDz
SdaHPhKzrALAf9K7elEXuQQ+htZwAmqMcc8cae03a1gq4Yu6vyZMjy5tR3YTQgeK
Kel0ByzGTciBILCauXdmU+ZYZeXEk75GIHLpJ6YHFn9sG1kRT6cQ0Dj5m0RvTViK
wY0bzODFvSwkE2B6EXJPlqh40KnVQ1HtUsIxi+5aELs6vRdUVblAfjmWgqbhVuvu
4cXlow/PPqk8Lco6aGRB22RKCPHS1acaDwe7+0S+4j1CF+Px0fHJBWV4EFmYqac1
lMLyq/GtH58e8U3A5q3idLxD8CHfymqTSj/gXV61nRNIALVCCO+kEFFKgkbb/m36
u8nbREkBR4Ace7cd1Ci82dIHKs2XIk9oC8+CwC2bMhiTwq4RIpPMyKESuwegGpQA
bWTditTVRu5TUTyaCCHdSI9g3FQcyORo2F1tQmreYTYCkKYtUHs4MsgRe8nZk1xF
Y0p4QqvBEx82qm9t8ijnANUNOH/cGQb4+q0NrGWQIovAGkFBzG2ZbvgjHOoieT4p
7wxlOsKeu9azVsWh3sD9pij73cr5TXSI7/goVq0ecVQjlH0URttBts+LhYsdIP1k
9oSwG5ZkAUMZnAyxa4PGjp2Idte8s0fy7BtK4rMLMOC+sdAm1hdwE3wmyl/NVB5r
/2XeQHOV+ianyvEM6jVvtXn3gEefsqRKDrt4WkLAXfM51jM4vlO4HsF5FLZSeFfT
fga2oF9FnAjsNRaPc3YoyKU9RjM8xYuHOLDk7TliJp0atPi1GRqdTD6UALcHDte+
Jtmag5Y6mK9YIxk9NFDVwDh6ylPiw3g2pOAqX6AHolCosj9g0vhE0WuSQ0ykkc63
VHZ8/10dxo1yVIfz/p0/XPIV0K5sytCVX6QOwAxvV05y4qyk+3dYdDhU3AeJHEnq
zHQXnakW8h823XUqpKqzGmJGUAK6UOhdKz1LwZZexR12U/W9B0LuGA6W//fFcRd+
retTn/BPbuwmZexPnyit0Ta8Kwo2QHZn2jLv+alMWa9dZ7NEY80OIH0YtS2qQDAG
QT1tEN7FnT4ZcDXn1z0W+bLhJlX3TLEk3JPuCezTqEM83dAAi0mso14GY1EflIWv
FEjjxF2zxpDqbKRTKwzNfT8n5pKVW2HwD4K/KNr1pmUAQOJD0EbNm8di44MnMb6K
AET7dUuBQM4BCMXecF6GnMKSHD+LB6R7WvsjnzV1N1n1X+JHkWNYao0sCxZd7EQW
H5KhkMQ6biIe6QzZXKLs66THStQ40Eh72r+G2O5rpDy5aijsp9rz69kkP61AFkm1
oG8zqaMICySecHxiOhetvJ2+4fVrDG1R7QFkR4qzkdFdKbJUlaawgxaShrqiS03l
oRmQxjGlsyffHSA3MeuWvK6GAyEBtw2Jo2RzgUHV5J6hR50088gaaGjZDoNrd1j6
/oIg2DUpX+5vmMxBeQ/QjoD3uTvJWFaTpTWV/NLEHrQpFYUfruphJyQPSggy+spg
KZ213lmim6UbgGMZqEv4c2yu8NJ6qUZ7pX6xfjVoOf5ZhrdvC+qo/SKNX8rpzhsR
fGUBrY5QgoC8BnAFbsmLHMCRmgElOpE+LYPQMcW/ywQEJDI5q7CAdovPcWfYRAlp
a6RuB7J42xoB01hSJSzNF1nwfzuRewvWVccsAlqX8HvPuq/Cnz7V+4hC2jbk164v
jVzCEcyd5mgkhKg/Bm9VEvM9hSdzy/kItEh6C+6hhG8Cp/K7kiw/LpG6iZjXEhAd
fb0GkveDpkgWOZOSthZj1m0hGDYjD4/6ct70GnJYogBXNpPM1E0681uXehTLfTy0
o8WbfMAJyJESdx47t/CWwP6U0rQJSuYx7W+QCwGLrByXcWn3cryIsnolWcEjuxtV
BsypqKrtkUSI0Vxkqd7dJlAwFM7pKcOl+7j0Na/z3G6bRE49aie52nDxNsbsWUvg
8DkoXH8Wif2XndevMSmfwIP0Ac1LQcOCkHNAxrYKev6GqEOtZD5edOQqB/Ki2UZX
YMbtnoK6orVhesDUunKA+1GwcvpDibwVowkchzJhIGrqy8lnq/Pd1djpUgiybjn2
2TkjEvowtZD63ytEg17r+GBcPQGbT8AIujfjUlv1fSc=
`protect END_PROTECTED
