`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAdAdQWYmaPnZOOZYw0QVauJZKqX76cVq6RsTysRP/4P4
5Z0d92wuU0tV+79ZzdlXG3vZmOw0S/EYf9w+vXwv0JAqYLbZ17iLBCTQMq1qcJq2
LhEAdswBGSIhw3n5UMz7EJ+jv7nJFsbCMgaq1QpoxkPv6lNK59H27IlHQiSDM5QO
RV0cSVjzDJYjt2s5c6ygGYZUVAqjob1FFhURP9hETb6InnvfW3PJPfrOH6hCJX4D
HEwqZHf8e6OISPbWxGoB0agQlkvZlmqRFumUzhykGSlkpvKmAfQZ8qeVLzPcG1g/
DXUb3ClH+y6dkDlxQq8LCVZ3uKg4JSKeS16gJcobvrw1zRy/EyKGpYcvLzKWixNO
Ncxvf8KjFgH5bJb+Vj+EKnePfYRy1e52uiVNiopFxBSC2xkeEt/XmbPhwGL+IKro
F0zylyCUvZG6hBG/HXpjoGR+PjegXUQOM3zk3WuI0HhRtAf7deldt33Y3e/9Vvfc
NlVqeYlrmtwxUQcGxJJDCdzL7wOO4sYftYJgpAuA+pPItd0bxGDPYLWx0SiDG7Cp
XmilU+79WHpPsQUoipEVYKeuplQFlIPsc2+ywDKUhI4jBIYRZC94WjPjxe/hnuXn
6JU/LzY2PcjkpLCW1wPSTDu981YRCkt2J/YAFJBzBrAhlZ1ZwBdcwd6xCt0qsOIE
qwXZf1p1Nw1KY1mwcU3WqW97ztQHUwYSWzpvtGpz9Ct0yS+DZw3b9pE/6ALn12E0
TNa9wz89f3Hc6om26oqp3Q==
`protect END_PROTECTED
