`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN8CFJCPCLtr1azo6zvRgPhu/p6ghNqKsUoU1dIOjhKBc
er9mX3hFFCx/7TVfQ2OvoECWwA7KpP35t8og+qWBLeopEPw59uSamR0fdsQ1Jkmk
prmRhNmwcmW4UVT47eh/g6EkTHtyHJ+Q9WGclwCdWq6Zl3RV6ADpOWLhwT+rISt7
s1JdEFwkS3cYWg9HGxL8HwjX/z39sV/kwGaMlyJQDjrdfP1TjjGvXlu0382t88JC
IJr7IhcD11p4mul2d+Gsx8xQwvcIPneATY9k0f+X/O5wgNghRwULixKJaEmMyDuv
utsQC9bVBqwE7kBqq1QqDYWxoxZ/bBGiRnVQESGw2CThJuHwMIOSIui4Dbp+lEhY
B0rGEixbyJsva9SSVdKVMXXFBST3BrlrMS5qrF3yK1/UMy+62WPLR+fbQZVyyWRX
TBSSW2rk5HZDYFqSZ4xgqnjPt4hmTmu7a0GeB8wFJk0w9AKnYvRtC1CP/3+HnMiQ
3RTZsU9IDVoCFH4SPp68eTJAI3gVZ+BuOPVkfEyYNX8aHKnj0aQIXH0b4PZ+e/k+
8n62kdvNAuB57+MAaSLRy/sPBz4oCd3UoTJpEqdIppziSsocXPk3JSHFia+uHsXs
ox7knOYgQSFhuypfT+yuWIkVLhbbAjsuTn3DnLrtneOj0p3R72OudL6mPIyG/rov
HluGp06Bd3B3GNoinlmd1t2GlcWfm4J4HGe9XYlVAVaKakU5nhfNucitSq1pm5T7
rqeBRXO6yNH1mocOpigIPBbbpVyMqGlvleLL+1HWoeZGxNRxDvOzZraQLhwWnmqX
DTJj6bMFBUeISXI06yq/5VIs3HVn0ss57WnuN2cWvEN7jFnitSEmyB2XyCgudt2J
WQW2wam5QZMxpog08fyg8a3iSjb9fwJhlgD0PEBBXIKLaNL++dCxKx8LWt0ZzVX1
C4UNuEKK8H+uVA4vvJ1VcUhKkXuruZMKxb5QnprisFIn5JdzkhLq6UTMkEK6RjLa
E2Uws0X70a8H0f2d6vkwXYBVp0xtK3jbRm21yzacw8OjZaXPtp3B28c5OMXcEEMp
7coIW97QvzGBLj3LEcqznwiX9ZimlNFPxGzCHFVRgLTarjsD2yenCaDTuowug937
zIZBDBwC6dJ9b8tYeDRBbwpboax/NcCIEmDpwgY+PMX4k6UGSnaySfio+tL3IEMJ
V1MWZ20DUrFOFfEtPhykEnxUnpIljues2szSwC4ucT4PfbT52wyHZnd9zPXZtoSh
2q3jdeE4V2YSLhOMoiKg0u5wDz0uVwRImjLbXSUZi3t0IAHzQZDA5wrWQcM1dIWK
BTIM8irtMs78OyZtX04PZpluFHYOYcskytDvevNGS3+XIfEFKq/q3muTJtSRxs6q
4d+9rQc6FAItVudJnOhASOo5oJPPfr1ZH6EZm/nee3fcxln/Wkp4DLubbYCUK913
FjsR7cngQVNv+BMF1khnWpPgG2Q1BoVZYfZbsRYyL287hPWhOoukist45tHIYNOr
rMkCSkGvSUz4RyifxLQVQ7Hfw1C3gEz3Ek6kzUAETdLA9VEOkgajSrQtamRX0mhc
ekqGcQFAAWX/7geHX0o2yzrrKQT/3uCkQsmJo8EkhN3ZAOQZljQzZSym+MlG2V5p
fmAlyhB60RWcDchg7pFMPC72PqaK5G0XT8Fhk5KpK0YWzKx7bxocfw1EmIhH/CRY
BHzuQW42OfQveNIICICrV4v9d6y4XSOJkkJnXZHmBsQ7YkudBzChwX0mYCN0TMMl
/Kh/sXM7EAq0usqI0ITnGEDnoN6GJfIbFIetPfXZ6n0RGdZH1JQCapIdijeFeJVk
VCZB0q+cK8cfGdpmX3akk8UdMkpYhrUMRKkPfqGIzkb462sbZVZrW712vw/Ubl7w
L2qpZGyd+rTbxoX5/RaWqjvSTJq7eP4Z0XCYBx4Ey8rVcqFbZEwww1IusqRR45nC
6xSDxkX+z/Cm2QPGdNyCLtC+7YWKddax8sL1jcoyRyfiPSpM9uY7e8hvKYT2QB0t
Jb4DxFhD3pOh9Ws9DO4Xvdt0lkaBYcsurbKEZDoi5AC5vYBJ73KsVgH1xxE1KZ6X
Q7jmxiDzSxn4oC8TEN1+yy9zKu2dgenYWc+Q0LpcILadY4lPj7IqlSUVOLksoAjF
ZCZXOY4srsOdJs/z+JAW+w/K5ox5sqkb8qirl288nekLH+LUkqMqJ92ww5icb4ms
m0uhRQqoHQG1HzS78Ce9IfFHXhGl2zyumoeCOOx1B/lNnlM2uittPg1ljZGaui7r
CBCT7LMzG7gPqpmhIsqXjHU/guZw0nKt6ePBWDFrRW5RhOEX9Gg4ObY+EZF+3L3E
d7zhbLsdFQxBGuPG8QA0kq/0IZh7thXeJUlZF3vNENP1OR1MzFffhihB2YmXSNKS
E82DCUYpoEKcEhqkPKgFsmso/WuH8L5qzwBDaIizsoeGlEX006NupdwWz5svaSmO
DKYPS1xLkbXCmPdb9CAHs+T/PNL7uyKaIbaagdirfict3QSpTQvVNJitYZj2C4Qm
fTYtg3mxnry1GrgiYkuHBITO/XNbNq21bLDSPIySaKqVmG3ZT1BXaPkqyXsdlMZM
0bkW3d2YRbsj1CMjlhbPI/DxkRAl9obYMdjH0FUx8BgqfScEJFTkc3/rwlZEXUfl
tw01cjPc74KyceuwWZSt8ve6KkOMGkNZq4NCx2nJN8O/3h7nMAiZqD2pgYpRdhNW
ZovjiY/tHY+d0IWi1/AZ4dzY6lYQK51cECPvvwB9eRcSZ0jb66YJDUhJ4ieFEW+x
hsNPXFjxBKv5xankP33u0Ec+zGTpjy7MyiL3f6gj2+jQAjKQJtgQUsk5fLq43gZ0
U0cTrdyTl46QBSVP6q4a8ZUKrol7sPQ3qle2POlmn0cqLtFAi+mTmWcWeslmkj0G
BA6wGA04a++4iIhsDsSa7gm7cuHBYCrCmk/JQs+mh0M+bp6ahLoAvPsLYMfv6cK/
0ueCzQSViRlkLjQy8Nn8Q2DrzMeW4f+ljYEtIDzRI+XmeHl23BHoSXw5UgM3cGPn
oXQ2zIpUTdz8LKTwi3AbyzEFagT7wodRRhWaSNMt8XEm/vcEVxkwN4T+jILQa2MH
gceKV7vpi8p8Lb1Y9LocKqrZX+PN9CIUce/eALN9mSW/AhTn3MOQaCFW3hYYsnMW
QyjaDt6K7I5oaFKvC9Zv5WuUW/EpulMJlRfOe1IEMkLwT/UImBZAObA6ueDbv3cb
V+28flKI3hQ3Wax+SyU8AdjCQfny+a6nHpi8n3wwhgpWBDRpvbsoANGfRZdKNj5g
X4NT3ZYciwXS72lPrcXz156EaGuE/aqcqFrWCabHkxzuzsPYIsrPhzZd5Jap1NyR
NvEKfm+d5Zod/Qd1tbKzl3z1t6VpNNXJQ5FKDhrg8dzd2Zs/KWYWAJQcnkRCMZ2L
oWRRBZLpBri+bmzM4JfVIXFy0Lm5rdziJUdi/XtdR7NO5xteWgpZ5IupsL6Fd/O3
q4BIgrst1xKTi69b4azDGa0KbGXgNdF7Sy7ZfKfh8FkTwT8uoFVRtGdMyui2zutt
Oj7sgzUnJ9C5tIoQFJaCsYGe3iHZeCcPaDjWhN3W5Tlas1PYI4NrOhcdl4NKSd6V
NiNeI4R+SMmwHRSYkQMNhHOz5SiiQekC/0TLOt+hJYQWMjZEY0tn13ofz2n9c/wy
pMlFuNLHNR87sMU/WCdLI4UYf+pUDvrSBBtrup90OT7/U+OKe8/NHCmXvNOVpw3b
TJw9rQhHt6PzxzK5n9tTFcks+ZWlKcZIXc4XZeYQUbNLlr3t+pNQ+jfJAXj8/LO3
hvGIO2PRutUG4OFXmA2S72Yw7johlXN0oIf2NZQt0O8Fl37uAKYp1VGf1Tm4Tzwo
8Gh0/lyjUJEm40cjpTHCapHi0bWucd0PesGrGJdRe0tdI3B2e/TlMknR2HIlzo98
RR3tFo4UQEEYk/hjPbReOFknxK1j9lI2Gm50i9Ubqy/8OAARm7hFmeGgE5tNZYDd
9XRh6QmmND43c4VoF3YQo2X5atEgaC+4KEyN1UVfBmqPvyI8QJC16KKvApWY08tW
CrP0xnvtyoPnGnFOjjAzLVyVe/6lmtKWfqb/erkun3tE6NQnVf+Fh/GGPTG+eiR4
Q9XD7cx/KOZzYDudXKkohqrHK2cDzTp4qIapUY5giMj9tpd/S+/xZSFWFMA0zSJU
F20i3Js1OPJQRrWzHl0wMs1mq27AJtbKj2Tfyz3qenixIPHTmiXUt7Pd2dyhe2zZ
fJrRbh+Rznh9p4kx9uJwMMDgoac39FvxqlQjly/ovH5HpniMwEwnnCdABK6K52Rn
Rc5O6WkslioEfibxFyGdwiZHDWgmzElkHTFn3A5vnDnZ69fvWqLxwR8VBsMOINuQ
+3yfOCge+Ew7csR3spUdWyYl598ZTaLhJ0mG5RdT1xWacUIc7xoXz5+wDdpPk21u
p2SxnJNSQCjxCrZb6NpKAGQkDF1xD0xJ3/gTK5HxOjd+7kQ5I7IUeNrLPnwTIo8m
i2HfM//CAET3g6f7vk6zmH0c4+FejAcVbtcTsvWaGOr3CrYTPJxdDzvOmlEs7/u2
9ctsXt6BPzUFhXg2aGZNHf05wRgb2wWKccOV3cZ+c26MZY8joEX/P7ssgkSig6mW
uJFMGo7cFX/DT0yOMEbuJqTh3EyM1GGtYU7/WFDge3gVNKJuF1j7cyZEG8ig0/e/
aNL0V+Qq6/EHSzOyROP1a74VODjbivksN/99MUYA9cizaQZmboQn/Wcaoe3HgrXu
bDkhBZBGgp2QMnuNwxz+wdHPUXo7mjZYG03aFa5+lTz1eQzGnsUcX+5uo4i+rfdW
HT0c+e5rL17yztMKRWtXauJJ7Ja1LyTpC6AZSRDZVa0aFY7jP0MaoAxk2Q+Wjt/N
6379/MqPjCSBxjr/+23vnxudv4HajPRYao5ol7j78BGbbX6u+Af+AOHM+2H+3KS/
GhtwHaC0uNjta9nagdy06UIH+78jO+pMtmSe3Aghw9iqtlbW3zTgbWBFc5Es1jmt
SmgtqzTyVKV8wofcqWWM+yYzueOEYg6W1aR7bxOKKNCOD6ThB9TcZOA6VNNN+u3u
XlDjImwcRPCX/9EU+6i+KUFxbmL8gK19z36tK7pYpYop7rybcgMWH39rnUHy36Pv
E9ZMSqXP/Kt/hgFjl4W1GhuFi6YzmYW5MIm6N6cQIXd+NbvNohHONjdhBeH1Nxta
fmZx+BhAS5ToFvzY6S5QLcm3KRuI3iEuO4g6cIUDkkMj2mmruAmRLH44sXFzipQ2
pDkjHuuUlP5/izMGVg/KcujvaMUm0Ce8pkC/zFg3bB9COynyHpgNl/2Y9iPaB2Qo
cOAxOkB5cAT/5iPBHo8ueFJs3l6WH/pv8rgyNikdbrPhIzIxPSJENxAQzr3Sc43m
HFfLQqY1PwWKILNgXA9QK+3HVMmBtyZp7h1Vch+bgg6VU23Qnf/F3MBVod/PRo+9
uchX2dZQdUgFcSFoQ+LRZvyEu3tKBNwybnGxIsYJyVeuUQ1QGJF1WcSQZIi9RGLS
AqZ9pW2G3AEIAmmuFj0d3s9a1cOg7sKzCoW6GuJC6xM+wB3SdS3AMSYAQsxUeCpN
v4zflf7w6HTNTJXrgBbjdkf2TiKl5ha3Cp+eshviPi1Qgle0nMdNyawF3Hh2kXSZ
/AHTGJicyL2X2O7Vo5FR+CJqbp3tkNli9K8GzVzE7lFp+YtOHWsTXoenitt+YkPa
SBwdlgqcyXuUgTS8bsA08uxsRDKpxBS1Vn0xPxog0QAWVFqvfGRGqdfseB0s3h0w
76l24g8RYbpAVqjCuIHvHtDj99yzy+1/Z3J4aaDOJYr0JpjuFlEwr/axiMpL6YqB
cNlAGBT0EMp6JM/j59DfjsCIt4IRjGLzg/hagnnD1e/0Z675E6TJHO0nX+k/ywPl
/guY0KgN32PotKBO4r/oaUP31BKnQz0EaYy+0pKybzAG/0hlSESMp9ZV2GuE4cXE
Q4mFu9UAkJ4lprYdijB7MRZ3/gOiIx2eAk36Nylwrcr1SaqsmWZwzF+/gUTvH8Ou
dF/RTALzAs4x7GpCRBws+08n6IOcMxFe6buQRHvhCWASZ9WkBL9fZEHAY2cit7QL
kx0EqS5cUq9konpseevG4R4lNRGFi75v7NaKleL8ZnY6tOgsCRkCHJP1Fvz7banM
ynX99f+0au7zGD4tRVMEw1VOH/1rJim1ExloseTTg7xVuHBh80QTr3qzkRDLuG6r
yMlmaGOE/W6ANfpIfJm0C8fYNwL35QaBwgCGiAX62RofIAdIEWqq5PDoHj4y5+O8
JQ2Hrr0o84h5XB6J5UIZdPx1ZkwbZOZBymopG4jrjcHCOoGNJY1BtkpxW4QIc3OZ
jM6yyPtnawFbv8hLO8r3JOLdL+XeVSqF7HPKLJbF3WG9tg9W8N8JjWM3gEEJjeA6
fOsBQcI8cMPS+yZg50xMktXfL94dcLbx5qThr8W2kVo/eqXdgTSZCrxyw86Lq9xn
1zei130BCsWVEcxvc79BNYx2QG+5mD1KHkpyKKK1x452UhMWzh93jnjtpWC++KBB
ZxDX0DEk+49c/fxgFHlCaZr6/8qQ73tN7c6zhik0DLnU4poF5UsceV0pLlJSdjKZ
7vWvEQanSpRnjSQyeV2cEgDjNwKX297gNnqFemB7Os+bhVMRQen4cXz5AysbIxBW
rQypsn/K20dQA7+3JpTZaYvs6LJu7HQH8gy5G2pfLdv+Vn9E7RoEm7FxlWDRFjmJ
uBPOxkm+Wzc4dBBmz1cKsRMn3UOYWRReUjVUFgwcfcgmCxTgECk0eWyZ9QZUAoto
+Jpa+hcq3z5TEjJsMLDFLoZMAk54ScHdGs8DgGS2gUy/rKjf2qMD8AUPGyxaKKu5
Bp24rEH4vBRz60LepCfwoOe2G3DM/OKWTc2CO3fPw93MoLpx+IEj173bCMDOEFfk
IhCE5jPSqYlrwIfIIDPjD66sCGt1B9KK4b1cfvps7No6xFKnVyZVe46LquBLIna3
S9ljTFVQpwpwji3HLcjIxBOB4DRE7IeMuuJYw+XGX3jupzvkfd2LAU4CLmoY0HxX
fD7aCkzy4RO8QgxzBsM4Q0BS2DrsWkk9oEXpRUx2JwOlQ5nGJwgUd+3XP93WFHV0
8lxJOiwf9s+WPXgI4ufvdT9UDoX8MzxLh84vQu/6wiZFJbxbCnc7FQjuO4HiZmy8
N6CWLH8qH3XbJma9Mc/011Ps5rItOO8qbXQXLcz3vnlnlp6pCtPD5nwHa30gLwfb
hHUCb+2tN45YlWsRt0N6FSSQWb4WDfKrYH08BAV9kcRCiyeEsSH0RDeSvO5x9cgW
0CM3hK9wWn1dVIMxIDnbr5NMuC0CDFjFfQkOGhqO83DzQYaZM/cntYX0u2f/KN3B
4IOElf3FwV6mlhKNJOvv5mFzth5NiXno+jQB6j36yKpqFw/LfaOSlGQ50hb2bW+A
5Q5ucwPQ6gTjEHX+7GetWZPG0dz6giWV2aF62JCwLi0qIHYdOyDPoQ9gW1sex1oY
C4RuBaHmUFSf2Azzz/V9tZZ3UZSQgurl5KM9HY1BeBtKaXjCoeC+YpxWS4LY623J
D+79Qw942GSdMm2onfHsdHwRWSuKQxAE5MUEqJ/OrLfNwGNiVRtRCNkL+OAQ8qiZ
yp2CW2h5s5XiN9ozMQ+qOe/K8+ZGD384U0RjQln0dV2bP9AIOZlLZvQDGSFXMJcN
aJGx/V8yro/If7Fy9l+vY51HoEIy6m1H+N3eNNrbWOjGTEAV3+KP4pfKOZ5P6xuZ
IWkLwYe5akA9A/Xm5RRXmNO59fliKCMSBxHjBEBxLpnjQJj7W9nEUsDZwG/Rd4dV
6+SYQjAZ8+/VNDdnadeJwx9aPc/lvDyp2JEpHe3qeGdK3Uc27xsXKAOd5gUbT1LO
a89EZ1lG2jU2+/d0GqZTteNQlUg7Sxryh+yaJr/chVlcZphGnG31jv1JA++0NGc+
Sd7J2Vw6aRzgCa/G7XLt0cLRpeK6fGc7ofAnoyfCo/5UeazQgIMcarufI3CKcVBv
rMlPE0pP2W3xi+gXwY701c6xyQe8+k6NsIZ8bOoa+dAu5srdAjqjMLHcrxGXYiuO
+T6336yeCmZF7lt35ZSjpCSVHiUj2aN+YnHlBqEKDHbuDUE4HhbcG23PbNKBv46v
bFkM3Q1h51vCB0chKJP+bgoRP0kmAXpnP3myVd6F5iWrftiqDprGjcU5IQJqRe+P
qOan7i7R9RlVT9P73vtlB6TnggbqEF4c+EwR0yPTpjwoE9CYLIPpQJ7Ame+Oyi8M
DDtM0iuqnytCeZ2h0m0R2EYODDljopVMU4B/QwEfJeB4E2KilDATUzmGgNakePPI
1rfLkleRkckNBTw0cMVTLhx5OJL4L6zRD0r5SizcyBQcWu5WKogbO55x5gU26t4G
/9YjdkfL+dF1WjsDULbavi5Usj6DK9CXwOxJp/uoJm7bRWO6AgPnGtw4BxmMSIZL
Ob03EdxVx6dPtm8Bdd57x3Q+2549Z/tBgAWOyjr8yHsRNAmWs+u9nObmgyQPltgS
MZ2HPyHUN9M9luiGibNAPO0bDtlMiTYyI9H53WgLflSLMHEEhe7/WqqpahK7AMXg
1isQIjLMbmoCEfcEiWKo6JExiBDBF3AbvxHYRsiWw0gzeqAuleOCIOMW4y/mycGT
+1hol/0QZ9WDCym/57l4tOcEMvYp7btO0d9rOK45qjkg96OQiwxhDL7cZIGx0nYN
+Op+VZwcagDJBEhVaRRG6s7TCuN14hcBNlBnnp4gjfaW//CpLswXKrBmBv5r7t7b
ZLssb02nnjr+eZpZMTVGfLR+o89PaHIOJVwCNYbCawEmb9qwgHeke9mnn/moJqqk
kIFbf03mrbUwCxw9QiQnFbmaPr+3VbihL7K9fMJOh5tZWzmbe0aJCDYfDim9+ZNN
wQNSMKJwSxa/vKkOLJggn/C7xCFgynMH9Tv9xLTQHVxRILGIbRuXKx78yChWJoOM
rxCzSBUPxcDHzniWDos6RAAGENuPdWdGg6WUtzvaUuZ9MQ5K/7/g6sT8cH+NiopK
COpIzrRMbUKY/qPq0ZPhaSw1QuxrDw+b6frowHlJ4bPLybvkm1MGkD4AFokc0jUj
reGNSKSLVLzr02ucMYWSKG8c6AkmBwShXjM7IOpbhE9pkBwNxs9T0z2kss9PHq9v
XjjvlJp/uat5A7O7joLZAn6AT0f0X+x+JwvAiXQXGOWGffoN8g2v5hKEG51yhb4F
h3Nu7xKDFcaOkfDh8jm5Vt4Uc0j6xQixsxqqAElaQXRumHPaOVRoCNlgWv5ZM7Fj
WMrMg3UNdQpK7BsMrmhMTTng4oVou74InDviV9cQhbSV9bTA/LWwjGd9AIJsExqm
CCEN4QVchAfglUKcW5K3MqL7cuhG2reiponIVEOx1eNh8BJb+ODcrUo+49FrIQ0x
7bS8LCziN+w8q0ZC3mWTUY8ipP2XkrdaYkem4PDUiZxh4lCJqxlAoP6kAtqLGp5m
8h7+wBCJZXmh1FCtXNtpC6cqORNh/bCMjdgofjBRFXWjMsK6jz+W0dT50O6c/iJe
D63snFOVpPjUyDUYLzp+UR6yxKgxXkwAMWWNmyZOBTsVFvHqUt5295aSwFDteaUR
zbIr0K0YNsT4a/h1XUfD8/gnhW/o3Co3eL3j/I7LhcRBL1Fp7ldQYKmlxs79Bt6I
P3czOlvsJExoKK1msajz2rJKW2oYt48/YacPWjP5OHK1c1d3yb/+le4IEgGPwXEC
9eDEb1TeORGZe67E/kDo82GznhecNgg4vkp/QliuD2N68V9FybeUTQkOdbdYiXru
pcGJ45JtQdDapt2i3NJoZYA3jpPmS5LtCog1C4hQWfq3o0zM53JkSt2x1miKq55M
19RsYEIGJvYQHjb0oyF8MpDJPB0TA1uU8PSHA2zTF4S4g9KIFSPI3Lae2LED0Z3C
WspWTmcacPtYDsXJo7XxQjYgiIsMxwTDwwlmUjqBlqpb0FYe7kCpXkhmd+4yvIn4
v5O2kq5rAHjtb7cM4KRnuHkfZuGtU4qpLKfti77YFkClE2Fve1y1kev22SerhVNQ
dbEq/AdNy/hQDYujgKpKngbOiWf0xLwwGvuooblaFZ0t8keUMVls2AV9/Vdt4t72
kHZIpBPV1RYydgMHzv5bT5DaD9yOgDL85tpg1BaCt47sqrHptEcOuKzRjk4cZqOZ
lqqy+esx2QF7Msiw/S7BfgMHIqK+Gh6cReoB8OKnoOoP46Q/SFfLczBSQNh9ZKzW
jt0O1WsX0N3McxFpPCVJhv76gOk21Ll1sCOM23B4TYw1UnugEoNZaM05scPuARG1
3ks3/NygfvfBSE7EMu4Se9skbsOCxtHFCaGo3JB1DrhHFdxw4M9FkdIc36zdKQzP
Uy7/dbtvJE8UnHgI7yfNy3svFYHCE9Ut6pS1TK0pmQSWMu5CQrPsV02JwJYXECTv
XveEoJ0fp3Z0/LgTqgnGHS2SnaphM/y309FScmbh6a4ifCueNDzJPWwxv8Bj9cY6
aiHLTqpICnUahQdDTLDk6c4mmCsofAuIhhvt6/ZycMZ0gUQ3lbpCLTCLGbzrPvru
MVhhPaD7/gwBvHWkI5K++PJQbFEV7C866j5xbEUp5ZYZUAL/IZbdn4G5c9ouPXTZ
t2ANQ0opofVjc/zQ+sKiWI0/7WyQtDssCpwLn75GKhh0GGLa3OQ2mMg0Ecqjl2Hf
bhQ+2otCzIOLm4hhJe49r3akJDyKNI9/QvSpalhKC+pSfI3qgHUiHf2nrARTgUqa
6pv4kvsOVYQ3HiaseoQEezByweEdnmxuME+lVCB5POg83nf+QEFzuqgJV8FAMsOn
x+L6PoAjEsCJ29qf5kz4JK71Wk+D0mSmqxORekkZfP/qz6q3t29sp7tZCR1WegCe
fbjpefChFq7sRmhIKS/OM0xhs6wZ0XkbqLZ80flLktUIFBuaZZ68E3qCQqyUWWwS
XagJOlSVZD4gNqQwPrHeqUTsu31ReoIGI+vz2FF92wcXg/qzk8X8rWw/dx7tPqUI
UY8U3Bxtfux8h7HZkdKeZEzw+zu391Y64iRFMEyJoyZPS6Nf7V9nm6dRp2MgbN6b
oRxbRXJE67kQJ3P2jaz0gUGZHatI+ncnWOz0iaSWNroBesjF7nD59D+Z9FWtsrA2
boTqFfw1zER2HFkIx9+W1MsDQFr3CWBiK+opo2nilCMsf9HTwiXG4ZPC5DVkDbOp
63Wd2t55InTnUxOzLmswCxWoL8+izoe47cacYfl2aFxFREYnnOT+yWDTHRdAOQg2
J5YWoQgJkGZgRPaMHGT3g1cC6P3CQ4wFGKBkZ/zQdVlc+Mgu/Byk2DbNRANHWKDz
QaohAcJvrpkPAVChG+WN6Cj2DmLkejpncUtw7NVPDwW4i04Scf4HUe3puDsyIld6
F0WRm4V1k1jJS2imfQNQM2mX5AGYy/nkNWXhOyjmWz+bIrTkKzbjOopX0YDDuWsv
ppKG6gCAzG/K7Xj7rhoWPHyZz/dwG72Rii3RQE3JwUMbznXmSPEly/1aGWWw/qwS
MR20iK3n3+BsaPXyQTAoRlB1yrCotptPI0jPry4MmIkJU61cD2AWOg+Cl559gnFY
mtlbdJoAaTZ0uJQLeqpi4eU0vj4FxzkiJcNmjQhFI6UbIv56J9P3SM4W6ch0gFxp
K7o3LPkVfLyHeDquyN0O+NSDlLT30wO2ppleFLHVERrGgRVGqUSzAEOFpIpv7L1B
m9lAT21r6zbvHkPwyfMpLlTmR9479RtgyFuaqc9YL2kVSS7gXKDVRYnu/mXxONCL
0Z9d8qn/r+8KeiBTM6fJwrKG8meo63xOl7M2ILRiTK6WfUyiEK8FHl7R2SfIPix1
Zl3ypOJiu3dIEoEq8itTg/0jqLaC7ZKHITy32uChL73mgK18rahEKpuUzKIbiamg
vMbjaq+R49v5wWJrZUb0DHimeSp92QXtw4os1y7zeafgQ0bEwg/PAKrYdpDYp+yI
OAeSemIE5w53YC4xhJoNCOXeVv/NSp+3FsqEGl1gf1t4Sg5UKVb3EfrzdtFHjRVq
0d/DkybCOqHXFxrmd2nzNzccU9pV5ReNiQLA1svlNotsmRPj4DRaUmWWsb1gMNU2
ryAzup6PeJQXE2qrb/65iC3ePfcge4zh0QcbuawELjP7+MH79et+PGJocpTnrsE/
BUdiww72CpxDS2RcnlmR5X+8WwlA17Xu+Dq40UejwUroZKED5yePHDGkb6LA7XeF
uEXMMUsoGJyZ/2rDVHKKXJMXwBwwpYlKNM48IHgwjvFkurV/ccuHgSKFT0XE5n9j
PgmhoCQLNtt/881i/7s2/pnCiJvYnsNhKk5oF+HBiDgV1S3QDFKrXuMDorq58tgs
m9bzKTu6zQgI87VsM/MoLmpvvA2LoPEahnXD9pBACRW8HxqiFprZXyCXTa8Hti4Q
l0tcYTx8PezRDIcvU2owF+pfIDqHf9Pf5w3RSPdJoTyOBTuQ8wMwQPULJFPZ01gk
i2DT8QV/85uQyIWHm720NGzKsAiYdnC8A1aQ5HUjW6WbvqEz13XuWNZg+dj0rygf
S8EF7kaAtGKfnAFJXpE7u8HhpOPs43SGd5scgKzUu+aZLMS/gHU35kzJQ7QGVCjK
c4v8N+WYSIATqiSY66K4llGuzdRNSYDu+yLaWcxXCtxfHvN0olkKtZOLPzRiTcqV
saq9sAczrZkDdPiw9nyhetqpVURYz2hgpfb/YGyY4LYDPuOQMIkOu//K9DVpkyn6
q7PN8PAUqz16HLRmB712cP7F8hW9egvPiFAII8m4C8YTYt8zS6Dany1kQpGrBOLo
YLGtnczYzRWD7wfgH7eGjpW34jzA5iRX/qorR4NYLspcwTHbvDFRqe6n+dSUXBkH
nIJzNh6vm6rnPvG7C+wbB2f3TlPmN0QDeS2JxJ496uTQlUMuIDvvmmQIKyFSgyHp
ZyfRL6ZcfLFTr1ric3AyyVO1UmGDuNQczqVHEZu5fiqsqMvjLOs219UxQdOnSOEy
96a45fpkgu/pQaswqJfQyZIyuwMKAZZbC769SjV7bCJJU5Puw+OhlbijqRlSO5ma
LquW95ZXL6Vwb9tEkmO0AqKaGyC+HnynkkKAGER71pbwRzRfZx4kZ5bk9QtTMfOW
X7RuXfrRKlBqrybYTPAcO+9beAbsgZVqcPdbD3FfB9kXq0YsTAG81AztFqjNCNO7
JkwWIM6ZYXUemYoqCqkpuNgFAa2mM32y5SgGeQoULoqGUuI6ecpV10DmlSWl6W2b
v2j/8Kx7tBkxEFJfCk8K4iNig4zeaU+OJjvRzfdyiKPnuZUTO0ReVe8hCC1PjOBW
7qPz2Tasb9pHaqWKIZ1wDhXbM17YLQlZ1F3B8/syqFFI3L6oLmrC5boJmcgQVcOk
DVmELcRNP0/Kxkkr1JIRNzQTaCHskEj6xFpqqR9vnzQCc1IWiNrnANtcYWAMHleG
BenVmbXx9Ylmb1ZY/HFl9K17gxqV/KFSr9jlCVl40f8XHVjfCweq0M2LOYcUHKnA
/5HsuWAlINRXQDlBE4LSNeHph0m/QgGt1z/fdNLStbUz/nPb8KFPkIxFHygWJKEJ
w0k7YWIg1M75CH2BofXgSotmq3EmtX8xL3QsogPXuqX3Cif7SgyL0barcWQ9z62+
IQtAAHyTxqQuRPPJgiw5cA3zCexxzhrXh8ib/KtfHL3p9LTc4UZXp96er+226AMH
I2ns80JWeKNeSPUaaJfhhnTKwsZhttXyocX0+GefTNWfkNB+a05RAKBT4RS3zhEL
UGlu72h2H0fHCu25rYHCHe6YYKUPDh/SSmAJvYVA7trC9sOPRoplA9zxhV9odSiR
Rm625BCb2yP7Vlq/zFI7oLoOX744gNG6kbDyal1GKwlvYow9cCbNV5IuzSdx4We5
avNv2BIaUVQ2jtyDClCY3LSMA4b9z7hyXwFnOUM6F2P9cbkyVtgz9bhghNnHqnMq
IwmJ+qAomgpuQB31+qtn71x41Wdv1IJOaG+AKkjtZbnBe0prf/C9LBqgYlKDkr0e
mSg4zjcoHUgpUS5QqQ6oYab9K/K+gKAzSogChlYY0c3SNOWXJgx+60SB8YckCJmC
M4xG94gdWlYQyaBUuU5bMQuZAGmEVGkc/efPwZgpqLnsD99D6HHlQ0vKVU0m3KrH
LqRfn5PYj+qb0zVGkHkhLAGr5aB5AjYJwOZfFl+ZicGkw7l9xoTJZTa4RBm2bygc
39q2GMtRv/C0G9BVjRcPEWrj6tWLMbiyNsp7X+hhOo7Q2bYAFiPqH7UpaMSVBVMX
0TZe3ItZo1pM6XYCof812OpX73atZv5RIme1d4sdg/bvxvP2tOf25CO2iv3/e3HQ
ypGeOVOcPXmdvVf88W0tsdEPTi+eeYiej6XLzH5yDbiA0pjmB2s0394l/K+J8esW
jeYmjmZvUOCFnENv/XVigRwPBK+1bSWkJnOTozYyV9X92ODHMYU97FDtfJ9lqBVR
hMfzNIIVd1u2E3uP0ljQOAboSJ5lJVS4wq43HQDo3nmnkmWwcpoLMmDPoQOky+dm
IU1XcjpxoISSsjcdASQATgoJAstX6vwtzPsyue4pSt2m6IKzkz0zP63Nvx23S+iC
fPBImOTJ+jI60w8opYmbQl4IlqRZ6LE4g91ZMPuXanzSS6Ec8cECwXLYOk6VWSTr
2lkLgcxf/t/pDCkORTakM5fnzGarUcke7XkbizFuXiRNj5/6tpMhOGRD0iYtLsKN
0GhrL9s122cwhU+mbbJpZ5e4PGRfumVUDfooQd6FUAVYijv//70L93tvXkVRLrcD
q2ZPVo33WBZ5h2ST79I8YWXClJ5u4HftlZNo314Eaeoak4G9h3vwiS/fX+VEnIGZ
hD+7VAwOj+09uRU2YkqQZHOLqJTmtOBQf0injM8OQWfbZSmvzWt6ulhO+qj6sTMj
7IQykVzHJT5Eu5+/lxZ/z6Q/wlfjdZQEyCn8ugrch8cNbi9jnvXshl5qdomX2mDH
56LTCe39m6Xcn1QMsWPpY1uHpXnMT4b6cqXxspyOWthctFnn5n0Dt32CLggWzmTp
6QryqYU9MYqyrsfhVm97nD3aqz4iOoBSrlkwscXo872bfcLBINXZxDbeTjO70Igb
qRyaxyKBD2o9xp70Xx62Iggg00QG2znXWIgSauyzafSEXL/O/UP5fbhGqd5pxKXn
O/4yLeW54RMTihqj8SeTH0VywzLuJDiM0r6rU3Obv0V/A0xjshl9f2Ve1tEkJyQD
Ol9jS3zPM0CNjXjUNpBvcZtTiBAjl56QSYm9x4s46hp4RyQdgrTi5Fwm95OnVZKh
w6RC8VlNAMRC+s/eTlXey35unQWAWkR3csgml9niYmiGBlmXuo8gfcfr80quIW7+
yjOfDgCovRo9jBjuWYWhtZGW+vnpTMldUh9L7XxYq9yUEq24mgjEAx5SLJDTZbMW
MB/6+mW4eiRWaY8ecZGwtNcZPEMAm2aArBvKveq/CHPzr9tsZtf9ZevOUUeHBSDS
esIK2Er7tsaJ/OETXwysz7FSNCjgxUGpeXHhTPLhK3HoJBV6MBCUQuccZ0eTmkBv
qYIFOw1sk9YVNdBztvYKCREo/m3EBe/qGI0yKL4ep3fan5YYqqY2S8nRr7XOFWo6
tzB6Dg7ZX7QATgcIulUoMzlenIQAg3moMtE2aEkgg00HxR2P8zJLAZM1THTNL19O
cIepbhBvu1Pe88ZL0a5fU4WfCd3MXTNcmOiBhZtAAoBaKESXHB3d2VvagX2R9N0h
EnsQTtcQrSSii+VStgsif22rl+R94miEOH8FyGt31Tjtq/VfCM2SKcsa2XNx46Ak
WOXc9pjLLmOPu3X2IZfPwWg0a4GHnbyupNXHm3lA1uYn/qJJ76cuoLmhyx/LF/Hw
IO8aAnixoZgFb+rjh++o4MJ0M7VrXcOIGn/SDy+eddh8U89dzMTkOuCA/nRrCWvZ
Mv0YJXIg5/XAzmMjGIn7NWF5lFwGnfLblVYSFLBYRnuXdjeI2vIGWjf4YudV1z83
+MniM/TmsfNqPGgzvPjfkhdVC204fW8U/Y8685Ojzsio4rK/5s6KqRzGBf7B0UUW
E/lK8NKX9t711ILwqakTyXJJ9I8zJoNOVVhMM3UyVoxJGuPRot5bKi454X1QfUzw
0PZF54bmLPE3VnNMToCb3uIi9Huns94Lc0VC1edybhQpKMkxhynguPDN6dyk5hje
XIqoFBDe+uomInFMdIK29uw2t4b5N0GaPcKjXLCaIbQhU7zktF1XuELc0CthFW7l
LZsOESIkmQa670Ax64wh20hUMPRnpb8DYOVpbH0B+iV89jObDrM+SgmBCcpZbZ+h
ACUzc/SOX0T7ZsOj1zMALdEp1LmwVChM+qB4ubPidfj2CPRqD2echHGFEX2h2s10
YVSiY7qrtfMGYSnj65mtnbtowCquIZDq0MQg1b+WOBKs7dEFt/ZtB7hfQUM1zQ5u
s5dbDmy1TRZYrqRWdS/fTmTrlrELmYlfHkro/V8DB7XMQVEjuPxEdh5661VXCjX0
MWbC2gpOFvI7LX742KtGlU98+Od0FMF3otlklrNXo3GthZQGWnBgizXQwOrUVO1K
t4OsD8cZnQNsjBPdIkTGTl0nDJW3j0nIXARj0bekEy7nTddIkUYWD97ntroa4oOI
jI/Zzkho8FofeNjXkRSdg182ay0FYkHSPPSJLywkUTdSf3LgffuGKyS9CjHBoX6O
Yywq4vt8Q5N/j5efKfuUbLuCSuPcenuPSzw+L3wDxQBM8EeNM/iFM0rbdF3bHDcL
U9EUVJFsPVilVYdM6Qzq6S8ywt/a2kSQ41Xz1yxPpDk26lZSmnxEWP/X/Otn8M3X
AWWimQHFvEIyKwmDiAVRWO33Ijszo2wRNPY92cjYGBaJ0BVrWsWS9O4LAD3fc8jm
YcYR+XbewrL3IOjedIYzFC9XBkfifbXwLOlU/x3G0plgsC8vF2A23NVks/tg/cvd
d+n6omyTiQLcxME2sM37vNJgZl4hTB+mtT3yisblicakCMtrZsLNsmJa3PvJJyad
42XA1LB/JMW6mKNc0Ad0oTCcrvtuDWZ9JGgWfNEMqHbQoLGL4Tw9nNcCYsl7J/Vr
IxVFWOD2gj0cfIt2jMuc+RbLxIdrhwFbFCkTsmtTlcT/Q59YZy4AINDmoEAFQm1F
9WXkPFdbzONL/xCfSLCGIunB/X042Lu6JNI9YMUe7SrwiX7WihM6fZtsqIHSV+rr
iOjGlgS/tUrCladysEuTpu1DnzPI8W0sWL4Qtrm6/U2K7v3s7fKT7uB5BgpC9iqL
Vy9+17JPKiFZKdJvV2Ux99McUVE9v/9abVzCiU7YG6M34uGZCX6TBq2TuRrlrB83
UxARLNVfpJhXEspE0PbR0UolDokmwL8Fq5YLD/8RPUbf1OL9u1by9X2upwuwNYKc
WuGx7Gkl9Qnne/1q4K9uHtDufNDDx+csztP7+Xe+Vv2v3hu/cZGNW8Nsb8RA9xRe
tfWvy3C/7jHhQSoDCZmtsrPI3VN4vmwFJGX8JI2tsAjZXG8gCbjqaBCg9TfZiv2C
n9npK/d7NB7awdWj1qNtn1eL/F4UgpHnpRyIx+hHawVM7lSa4PzZq7etBaBOAiAx
dx9/zSsWsCSPgUnzVgcqDD5K5nyy568BqBqWXBNbX6TpCjEGPUQUrY2LEJcSWfd0
BioLMygqQIh/nk8n2ot4+6NBE58d2hIlpgSh7yUjnj/wCYNjlneb81gdlZmWAGu0
whuwNktc87fI1SIzkMpaZQq3gJmW9CYC7FMo4W2Qien+btMEBbAfx2GZqVL/Eu55
VcQrKWlOn2lwGy9Pk8o/srR8fXcCh5oQdT5NJEHTjWX5BonRNupYt/kG/k9frEW7
yCJnYJmpa2lXMxmfg/KknWzKARObM6fAX6UXyaZH+MWYdthZ83MPbNkO2qYOZFOR
6uu2ML3qXOksv2NUmy1B9RnG6qLAjBZ7rrX7io0/gE/lKhBpBw+y8uL8B2EfHuWH
YJno8TOCwO8vkOaZiFgLYm0cM5Yew//17zjeY6DIWwjYV/27KgN6NoxRQJxoiBH+
EeenzJ+hyaYvFSdJUP/VwTlzByMiALTOSeukUiHv3J5r0Sc9eXa6DcIG3EJDxT7+
KaVMwK5/o7UyPgy+QTJYBekPKsokv8Ba5Ohri1oZ/295gmuFddyGyW7pQH0ZJKIu
iKsOERQENPnU6npjBV2MywHd8S9dq/pVsEU0DHwIRG4UhCTV5e720QzS7TlXCZ+8
7Wk3JZVGuwIQNtNFvgnnls8U790NhLMMZc+nIMUJUJQwS6FmK1ZRvENzfZSA18Xr
I0Cv1NnAlgSCOQSR3fKG6M9BwAUParKtRwtDfIBRFqSGwgVF60XN+7ef154Aw4kU
AH/OtX0X6T9ZplZ89kpeA0JimrtMjSw8ssbctsi+L98zzW+RpfsF9mlLwReH3dbG
hCem5G4ybai/+Kx2RLlbEIbDJ7o+bFTFxjJGmAOKwr2DjuOrcwaFYN4KeqhP/D/+
5TzwlTCLQfyj6Fzvti0JgAm9QXqaRtGckdLGJ+2hk5Bej9oMTNm1dWJCWQh0I1dP
mU+yCF0sHTvpt5ewwaE0TFZgOyRR7QMpTBMDpF7Scfg6Kzwfa2StTVWYHZdzNpRJ
WHj35ulUayDsoBqCB7ZY2LRID9wHr9BQS17FwJ1aOZaoGMN8B364ARFWugYsf4lj
bhXT3cf+tSqnI1Cm/UL0ksrrjeCZYIa9ouyYO/xfedyC8D/DGVMP4Eyb/IcHglfF
3w+rSowKNF7LJS7wEiRqBn5SLMXOu0ij3uhS3dG1DmtfZ7eWDVawpJMqz884pOA8
kqh5xeS0ND/ETPyBUz6kutkBQnRBO5hW+Qn4qmUzhlCVbML/+oBx8LwEyLr1zB1I
rZj2z3MEBSFIJwt8JSct0ZzEwXjQjiqtciach1wvlmtM4GIxAhML/yz8T92xd5vs
0Li8BM34LffFIZpI4mJ/7Ny8yu1/QItxeP4qex4DvkljeeP094CydBQooFNtCuhe
XmA97gjRwv3ovzrfFm8GMRyTBNnRNd17gTnDDwWPrj2vPD3dY1pm0zIjgBukM5ku
aT8EDpziS+yeimNxTsatZD+aIAsSpMmOtkdI5qdEpO6i1/SWmvCggOsAW2gaV05z
flllA0IaK4p0h5s1WOa3zBHWCBc0cdn4nHv93TbBUZ3EnX89RyDY0MgVBO2QQQme
Emj4ksQjtZcVlEd2TmA24TzjvYHO+mPVIbuLT2uAdbBTVAPx2bKb8nACx+fXukkW
pfc4AGWrdJwWXSZE5fhACJYRY+3OLA7PKwOkJ0KliVl8yQF3K4St6NWRDda+/ewH
E9AcQI9EEmomRgOIloq/4mc8QhEzP423KyxOthI2gi3Mdtd9b+YEHzyxuzHfh/KD
fM4LDOazVNG74FqRlwfdzbIe7J5A9rUR3avrlKGqqFvmYhCF/zRgJge5Fc0+WHLa
239RW/QCpR21x5g00fhd+9NjxxWg4vLozPyiIGODVq/5PGrjTN6cDKK5/224VBoe
WlPfs17SLin1zu2PoI5WfPZW7/GyPXtm8LU8kx39z5wKNVhMBDzlDqPqwBUvjB1z
8YSVtt+/3kQDu3N1Fe7RMhi7E5vJxMCq4Rc4nOEFKiNrAWlOU4ihVXBKzFbm7OLY
t1v520HdrU/iO4JR7iSbpxcrNPdoRRiKf6YQUA3+wz+r3Wb5R61wu2EKtt2OY7lm
BzSvmDKOuzXNjIOpgooDkLm36vuJa2lBJUzEdq01WZN/8SW12svfG8Ui3bPMbiqC
eoSunKGk0ApI8c+KIxX+hgY4tB1wu5kFxK+w4w0+SntewKUcV8aYgxx5FrlrWmdV
2jK4ScILclZJJEoLuV47Q/POzNEBC/fUkbvc61tXfN0+BDYvOqijBgLxfr8yN3CA
oELkEV0J3shjImKIAkwaw1+KJ9HHN1dTXc80F8SSYecC54AalWYHZEdzoNFCSKcu
3VIMcihQZtsJNmb5+HuQ9RDatATComwiiCHA9qtUuMeWYjZ4bJ/sDq/VVHAD6TH7
QBmxfn92Tm9YlezGyMLYONw9nZnV5CtSPT3yYOb5Lqjev4czUK5KgTdzHUBuJ1Y9
X4L+dW+ikNmPHVLwmhNC6wJJOF5RTOSwoCwmO+tNNhq+bJT78Ed16962IQErCDle
rzEX26Qdn0/82Q5M81CqeLGTuHcbzcnqmSkbBYtW0BfMdHl89u5XO9G8bSVgJXEW
ftoBSunvXXNlacUFSwEh58QlaU1ev+fBhHBNqaqQplg2yY3mAcOV5ud7seVGKIBL
vP/xkDLNNnrgjjjIvLj5YPsrQI/ebLpWxSClP25OZuuUVmmfCJibko+e/k4sFAk0
kjwMsFzD2Yw7lepCgQWHmHFnCDrwYEhcydECMZIRWhk46wfuHypf/KsGYR9osp/9
mXADoGCsQNoMmvEREPFH0zemur8epfM5gZ5P+jU04u4T844gwaZzcIybjaFTacEj
5UL2gxjUbLRXr4LtoIDBiIcpUQ+V/A5Cl/c08foJe4Y2ct/loMPBMK4KH8X7dhqd
M+giN/4hF3VGgCTUX11q76xFXsjEaTwvxcf4yaCumgWXA8LZmJ+NU6ZdVYlecpIU
sNVg7yxTTl6hETFayu8wzKkz3b7XB9yTwYQua8rnSQgIa8ey2QWm7F+rt3o9zmOj
/Hqd5Rk17+El97Nd2v2bTUiOlYmFzdKzpopJIagATi1LxJYt1OX+2tipVg1LO/vN
bG0o7mP4T5dZZ5Yed5vDfjyf5TV8iOvWJCl69w8voZSQBl25fpG+hNr6RUstVfSz
w7aDKW8fGVaK8wpAi/iEqy7Ew9H04nGffZv8MphBsGAcfB8rXWr3WQQg/ipCwX6T
N0ZsyWk2TuP0UVzBLmSqY/hDm+f9bekaBwUJZV58fTTjmngar0VyYN6RGVmD3ldM
4jcrbJfOJkf07emlo7mK49wr6VM1mYtqSvahhi+8wPp75mkhJCsfgKNcCcEiedl5
zUj51WcwRWypv6dTzCJFTwRQ+DkXn17Axq6laBwrjdynr7yRtVxDN7CC0Sa32lfi
s6NiiJ4YTkZeoBczNr+/pxqKKCI/wT7SecEqZrXrZyR/qLeqywpDnp3jBd/JTYi+
PVHlXZTKxVcaosBftvu2Z6zbPXTzd9Qa3q07miPLzDt3YsEiG89o5c101ynPWhYD
1pv3si6KqOZjhITLGA8QuyXWvRtYUHsYSMPg37ItYQvhgdMb5YdO8cx/sveb0BCJ
IX8XPY9HCC8hdoLW9vHzsZ6WbjdMmwTu+N++3IyVJQIh7KhxXZr7Z+cmzNuId/2c
90G/FEP1yd1lVIB9FZwjU3BPgjOhj/X2I3XfLaNh9ea18PoGeZmtJudy6MmMJBvP
Srqc2Blr9sCUXdOHcj8nReQbvuAN/o+Mdluf7YROMmrXtChf/PuGiqRIC40kxlGG
Cy2OhA//BCjDM2gr7S+kifjMisWa4WA6Fh7sh3yRLIpLboEpBjpCb1iA0wOw+122
JZCZmBtxZYW7LM+Ujn7pcUh4UKJVbjmdDps10DdYN2YV6XLtFpII2cO6LNCcZb4/
fXrz6fXfTZZXjNQUUkUvdCEmFCZO+JAuIUbPd2WoehQmfbgejNcaOfGpI1eYRcWH
M2TaJ6O2w9WNLaBlUaSaxcsByRAjLq/crLB/y5Y868r6mRuMQzkxwukPiErmrnI6
NZRbO1cIbS2wn/OyPpqq8bc7MQGUmtDi/eanP6cNZxLmZkzIdJgIcov/DDqMV5s+
kIexCEw0GHc3zgIVgel5KDF/lMcRmLDyX1cB9feRNZ+nqwxDE4Y4m7H0aouDnQfz
9zFBYO4zflJescDK5IQDFeZ0SU6OJG2hadzjLrNpBy42GR8l9UAF+55NZzEDSYLF
srGoFX1Wy5bN7C5C9FREcXKHq2sXkV4VqL3jlXa3UF8l7H0uOCPnvQTkYBjder0y
6+DVe/wCdAe8i3H8lrhn3As1uYv+RhfrOVAlDz3+HAtEvu10xtjIy48Z9AywjV4n
AYhDpsM3HkLUwY1mYJpBGDbvve5+QNcCn0aMV40zNebjXbb/W3X1sHaY0QK/xjzk
6zk3Uu/czQnt0BqKf5vsCns0hjMqjSbrkZWQh+ac/Og+38yUydSAF2hcaWcDUAzf
MaEpn9O+4E8qwqTM4BwWq6xC1xy6LnExAcOwEuLMvzmLxvZqAovAmwTdzBOae1te
1Mwsl6+CaczmjDuJivtI0EbKw0Dvx57MellZieLimPuIJFc712THBR7OprTp5PGT
DUngwF/v2UnG6b5HoAaYcs/QBs5GW0Adpr/4seoR2cxPhJ7ziM+X2SeBBWged3a2
cPlEkDhNC3I4tBWDkOc4wz0CleW/swyqwgY/nvIpuBKOdp14cf0BfgI3OO7xJMj2
In7MvDQNc6hmYGoLIuCrqTidzYSTYuJeZEBpV/S1j4X3xZ8CjXX6/I4WhnZKSp9s
P1iFXljOU3wc6v5w3/4J0+RRMILBl/Uaeozr1fHk2yF5WkxSrqRPpTIKoKTCfZXW
FRguqhe3BefmxTpi2dZG1EZyfpT0TI7864LQB1LNelNrGu2AVpKLVhN4x3/4rl5N
ORw8j7HS8iq4TIraWH7K/xzmJK4VGhMV9aItd8KVZTZcOYzPSNBWpCYfnH5nKQ5B
HeXcd1ROvWE/eOfyEx6KW7tErh1+vpx380RnrFYbJjjm81EaVQv7nmRx+54QjRP7
qNhiiOsUMU5fK84Si76FjkKwVWHgwpHXzk9bMZI40esYYGlEajREY25GNOi83cKb
HtMUOhEjOvHwmg5kKIXgOfRi00qbZlR33j+0WI7XI9dwgzxvZx1NjNwZwwTR55G5
JeaHKt8EWaHmnXiX2PrVOtr47GNDSX6Cw/hkgN8AUxLmOTrxB4QgvgKbTq+M4zZU
iVommG3HPNIr3t1dGVB1tQpWmctGv8hN1FUhBJjiPBMvokaWQtB0DaVMW36WVwEx
5R75mdHC8yCzT8+5PMLcyJ3ujrl/873rTT+dLj8oevL9kEyRVnrwRW5WWRvUbjGu
BYRYOBQhvyoYXMla/ztBU88IyTXMQogMqBD0tb1wP1ZeWbx21st40/PrZreo+o0K
I0GUg+TGCMpuAqL2CvQ6hwVwchJhGcLY1OHFk6Je8S7triLkxVEfnhcsHpzvfaiB
tsAsUc1horF/KLxV+dAfWJj0WNObMeS3hjkn7hHufUDPSwloYKl5RHEoAVwLCbCl
h5ZUcYHRlxAM98/kRjMNUJo60YEcYU4YNYGXvH8GU55Ewq+JolaJljW+JnzMQClW
6TiftptF2BOVgsw/6uHwacve7HiSnNJTafAVXCxoYZfOgwviyta9y8xshJwb/fq9
G7vdsQB3CR3DHIZSsSLzvdexZtv3SPCnOBb92MedrET9kNszI3SHcFpkLnzNyW9/
DjuGXHbj1/Txal7l/YG1+I6z1BqCAeL3Wrham0Bk5i2EdCjeOfHYWycZxSiI7zzw
zvBFOr2SYVOZD2Gbu8Ht6qwuYw8WAW/GEX4NL0C2yDsQX1Oy9bxrt6fgyy7sdIs/
XAsiQ7ttzdbgSoK6rhjISRLw33Te7b0R1OF7MFwEBTYgI+sBN9cWtn4iZESJkkVP
p6CHA76jaCe7AZiFN3S90p/tqzCCbsO1zUATZyavSY7bNxOtzJ//mheu2QovDJJm
Lw51wPXgFYSyngB9rbQzJmai2EshqQX6EMlv+g05eVLkp1T9IEePhYQWtgUjOwRB
zKaTxsdMeo7YcDBc/aVJtZKMFM1VnAyAjkiYyge0aa5+i8K3n47gSIPkRvzKdt4q
a22RLgSBdGpRYOuIWxehhbvf0LrQVuWvho04kolVAEj0RXpTKSTk7ie3m1pt3O9x
8JcdrIpKUHHoZomBqGui8nHuLp92TOaDDw8EFGKm4dDFzybr0GKFaFeDdjb/yT6l
isabTKf2R8T1MBE6894hKRb/qVqMhSRMz0vIeO41KDd/7hB62Swl9uPESfFk2kx6
2ED/U0qlNnxzyStqsGjpfP1UNjFyNJvz1ambFKaMlJys/JlX2ImVXIzUStI4Tqf1
ywPACPg2n03bKx11zwgOiHfoI8bm+y1Pv8gt/HT1O4KLKkhArQe5WmKITeIsgeWa
epbIntlK3XPsO/ALytDkpTEzCd6FpPgaEU0pdIuJOylIIHOVy19AOsEIIpdA1BJL
xZg1TRnooJAUyVAjmIaGRxHXnjdHfeaalIUeOeObD67JEVv8CCupEVKyQXnm1Gjx
Qa9jMjz/86Wn+lTnPkn0zdrqrfk0YMAxkBFIipBAeaPdwK6iq9IUp8O9q03f+Brt
CYufGblEly5+nhKPDM1NyfZ00qBXDjBhcR3YRAy0LOBJfEM7tD/veVoEIRTzVusE
DEqB4uJPUVuGBGY0x2iCG7F3okNS04SlZTkv0NSPWAihUHEOaFg57+2NBzOUBVuF
WQ2707eRFFDOTsl+zpmx9hKqqhPRoJvq1fE+VwsmmSVbJtsHG0h9h76zprvRf5zg
e3DJXQZ0Lw761Dz3YCAeWHtzsI9LpwiWTfE8GTKUAv9UOr+P+UJHxjFQIIkh0YP/
MfwC2LgQ/I96vzlmH18y1iGM2nS7bpTeGR6nVGdceVOoEwEmh3i9VdZxMvWna4BC
CQPbAW2jlb3aWRbZc1SYC2DU+QXro2mv6csnkDodoaecmdqlFE40CJ5IE+6/9mwD
GoxOrwGZkPcvbDcMu7xHsc7WlhrD+LK482MINjjdClJzUNVBIS7EYt7AUfoxawjR
JPnXhVt+Ski8ii4Y5sfVihdAQHmIC9Dfgoe189wuCLxV4ZEXJs6u83KJWkNrLzUl
v4tB0b2kqjTXFXXoLdzGEPCc9X4IjdLkRqDEEjaLCsHWcoG45roTyhzCc19Uz+BP
JTNVTylG/m8Q4PecdvW6vXP8lMrfTeQVu4v3EhlIBa2t6MrbADgrkgo33vogB/6z
1FZE/NkLGrjrS0mvuVgX4sKZgH4MUpqEplK2Z+AtEehESO8aUiCH2PqjbV58ommK
9JZLOIrLHZvc7QpTFuEjAjgrovlXFt86Mu0rvBHZiAC4Ok8hJbrtkaqPGGZctCOl
PAPun5wH3UPp9x0oTCtYaA86zeBuBuVpXY+OFggxb8FqV4gbQddvEYmLPRCinIgP
cO6n3gLbhVCgHzgmCXP9uCdj+NW+41Uaun0uqc5CvV0T5/BAqM4G9gxYSaEqs0U/
v/Qu9qf+eeBuD60fvs2BQx4Y87HDjidFH1N/5KphHFO+8MBzJV+PHS94YD2LEOTX
zSDqI0/Ddfr2XWP6qBI4g2W0sK6i7rn5DRRvI46YqvPcZqdEUoVIAHrtjXiBvaEz
daknqNq9HLA0NvVq3jQ5z4MdlNFQ3Lhtn0bvt92ZNBjoOWP0hz6T1vsA5WcJH2lL
gp+b4J4dIb53vXeV5MLVaXgKKGx4iz2KBTHDxbtEbBdADyU4u28Yl++Zvl9cjcqJ
G1+wsmsAQmzqEBBvB7TKNTU/A5nJvFsnf9H9cx18wU6IOdrNp4RbD/xmjnllhP7K
TbEfxaC1OYpJlngdLMSes+c93/43UcXqEJbj6AsNStTKtoSplOG82aqsx8c04dXF
JOBHWCS0Jff7IuBvv+zhjnWIcJ44cenIu41TLqpbR2CXXFk3dT1gEYIDAvqHcx2v
EH4TZUIQxnFz1hCuuImv1y8Yv//StqptCiUCFw4ut8GdZdgNaUqvyvbQ0mhESJlf
b1eWc8lV0B9ZptmILltMjylWpEihHQHOruFADcMDJxjgAfR91D4ZYG9tpYAiyxuc
vJmhVcRqu7+T5OFXtzLTbuiiYZsYOk4yPbssYLn/5YEIjYHrwWfyTs/IgNwdT8Xb
dgUn+MRkEyBqPaaGc4yzrIbxfCePN8YYlpTHh9Q1GLmY2j+plEqqhWi/lOXgiWQO
hbn0W1lYnjPfjRhswCjFse3QaQWAK9PkXsDwL/zmi3C+ebmXzqjab1QsRtLK/1H/
bWQujOeHqEbTm+SsY95NK2f/ygt21rPMFBT1AC9UYAtYDRbHG/nLXUJ0au8HYnhQ
+7UF+n6zQTRuFCVD6OyCRlsQ58F7+/+yaSbS/DoyhcKTtmmjjUxY34wBInVQZIxA
XmV5mupdRWCXEyfll+J5firaGHuMSv5Se1gBWydlQB53i7teFyU+cPl/1+xbLkRx
x8Ex/GEx9zF92i15+uJTd4wXdNIPRFICgwsJ2MYdIRiwhzYUmH0K5yvjEyOYYGFS
sQJ3EFgCpie0fe01XsdfQ9UjW9D0tmlx1cKc84ptV6D/L8TClYJ6MkjkE3R6xh/i
QEK95V+uC6Dxx1Ys8hkd3quQk7tI6TydMzGKJ/Gg19V86EW1pehIThBBNwRs6/PM
n3AA3Mtk1yPjq8v5FcoVlTkKFfa8zLlCTZuSVArA9NYpcv+g3DeR8yEDg9+MPXlw
HePmYPWldS9yVboYFYywGJJv/JIpUnRqQHiv6l8FxuqhAGegrJ4t2ihvEF9b88Qa
2H0PbIxeJTxwh5c9YnnWbi3UnYYmiUmbPNhNkrH5g2rAtOpwrSt7Pp9BEZMkdSK9
C6MkXXnIBsx0lHZ/oF+xbtfU4s6ysYPGtS6iBHizTGkywpiQZIItJm4TrwrqV5BO
G6y1qcqRp8MfpgIPJIdwcWWlFAomCJzYVA6JAWoxHl4ZAl+XmS9wRUJ+v7f+J4cX
MKfiC90qyMGMDktDfqitb84wY7bckLxTIZSEWRWUiTyFSIndO0ThhEMM3tNirWAa
sP9l9jOodHbKLHYhSzTqAYpk6b5yofmbZ7n2KMZoo+QOBDsSBx6P/rHalDBpu8T3
h1Qdw6BVLaMKeW+R7L5z0eqn7M6lFoWjA2fXdOVWBJJT3ORdkVLoRO2n5g0W6mSZ
V4nYSiEGQx/COrlxo7ZPI88ZqWV3Ms7ffIc/wdDZJBcyq5a9YTeuCTJqlN9fpzkC
C7k60r4HTgFE26eYrsik6oudhsjXu5SJ36QGwuMhJ1R2335JnzD5uglZUQN4RXVS
yCLTzcupvwKGorRDwAoL0IibnFxTr0tYjy5eDRbQq/f+9QJuslV6KAqY2DfxpkAZ
bVuBAeYMnXvemJrLgU/eMNTfF32pTGwr3AWQ3JJXV+p/UobxlzlWInKtapiaEzxx
w51mMX5xF1unYemqSKMMuV3C5EOo9FXgE/rbYB2I3bhVrfklOxNF7PbW55vdnuI9
zarKkH4fFXNJtUpCvbRx+xahab2aAkOwGowtoJtMIIZJHOrF9ra/OnseYCKAkn6p
KGglgJWTo+PtKm0jaIYDwtNif/8YVuxzv3gWrNmfIzftYl0t2TOTfz7ohXQIacbS
KLEUM+1V/F2NpMuTUW0W0OpM5k13nbESTgGuPXxl3h91KCcjd3GXoJzVgyJLJmiz
hj+JkFBpx/i5cY5bfeVftVGKGx+ugVycQS5C1Q7JTlyNXRx8wW3LxpL5z4+RsN02
JzC8i73pEzi6YE/2XpOW59S1kdq3UDz9cp80rL47t/i+E4xWGYYYdkGOijptWBEb
+o1kSgcq4JE6JuQlNDYFinDXhMkCg5hag8yWmjceyZo7hyUUu2lq6UYbU4b8yayj
ykaD0iLUgpBUcqHGuTylTQIHrZxwExPfM2qG7VuceY1i10hmnI3PV5LKjf+Um0Mw
Y1LEb/3gzsFHOR/2Anw7nwGKWjH2h6dFbmTEQx5EvpJzvUUMYgsa8/JCq0aiyjgQ
axl3ZPra3otvuIwRZwzRT+TJLCdAoaGpAZzMXxDyzrPB7sIXXzIfHZRseg75OK+R
1WTkEPuqTp3C8L0NmcrP7U3F7bAbuFYZZn7V8/sCXkt99qw3a+XF2IaawTmiFMTk
fYXF51DoLegxnT8BFqT0F7hyjJJiFG8ITFikXdZtum66UrBKOnDnG9Rco0Amlsug
1ITuhTqRI9z+/XL9lJfQV8VK27nbdoQ02AvEzIYFlqp2MOuft27EPk4jmmtXqlex
FAD7AzOKn5snfuzFIL39vULhUUFY4wEZVcN+w9SIdDmt1Whdvv1CFQPtswSomUOh
xBOGESJ3WoJ5cxthqU/LOeKqlqiA6sXbET7asvN7388m+H6FbtSP/yvlIzpJNKfB
YRvHyekgQ0WIMm+kg60XZM5GspQq97JNFdDvOAP9fDe7oMM34rjF5KHCvrkc9K2b
wwnBNXZEdq6KBNKj3aazXZZmr4c0EMYJmLpSq+xmSx7m/cDT9SHslF2l6MKaCPjy
IXGV3LpzKVatlZouQAZysKastC3LIPWJZ0e+AMwuXGmg12LLl1e7DR87k/iyJWVl
BMaSBo2Us3AeHN2symcaU35S22p3Od80QvQzQgTaWwRjFkjE5NxzE9ulz3/BJXEz
zh5stOVJpu9KkC1JKTIc5Etos95K2y44LS7V5ay5qtFM1T23kHr0PZ9VilUxNAw7
f+Et33w5rAgpriH3nGGAGP3Yfzpe0W8BPVK5UrLj4Xf6yEmI/SxflZkYmwlGrGSi
T+9lk5vRn0OqtTa3Hw2FaUpSVb1ebHV65i4P87gpx7fw4DeDIcmUAElf+KRWw1OO
kYkSX8Yk5fqrEqKYoTzZifRXQrgDFw0r9ShlA/x2uXCdqW79V8e11wRpTc29//dM
bksckkrKeFtOBZg1iWAKsgFdT3jZro0vav26AzropkaW+XAZSv8qh0BmE2yskmeZ
eLFXsakI4wKk6BgQMScrd+XvtSqDWNvG4EfNIAeAWc4sTpKM8MFcopCoPJGh8Zwx
kYqjbOhZnH3V5zYYtN1en19AJHdBaUg+HB8z3zcpw0WRpYHgCWvfeH5AFfX/Tyr4
yyD87oQAy0qvmdPAz9U04JtjFx6Dnm0GUVPHS3wq+ViJcW+UjH0fU9i0DyfI+/ZF
y1Lt3/an7pDs6QwUcf3BYk60QIAARxPNfhm9laXkY3GdK6nHD3z7D+Wvh4QDMDbU
PUwJvF1mjPK+5BgJkmnXTlxKSmnPh013G4PQGG/KuYEjRFiJW+FiqC+SOflzlBPv
KRStw7v5Ysk6j22blfUyRcAvcBxVapqr8huchUD7TR21JE+Yt4Saubbs4iByQiWe
Yc6NQv72aDkmGaArJP+NOGw9qAY4tgLiFFVj1lhHP0l2r+OfNGGCIdKx3rd5Ivjj
t7bUQ9pJWvY3VyCF50yJyKn8JWX6X48ObpQrXDisdzvS8iksKT13ws3a7T4TO8Te
50tlV80E3JhNSj8X8CmQR8pdjmXe2Ca7qqmHf6203+DmPoqVgEL5n66OyQj96doI
dW5c2/E0gobsxX8kNzkjldAdhi1tb7hl36PnDSavrLmCbSd7XcODOmxLclS9Lxg6
D04eTQVs1MrpuOUPivm7gWuTT12JZWCc859lMyyZQu4vdXVtxhcSvhdS/y6qXYfs
e3afeJKp62k6CSqc5RwBrI0JN8TjscboT7ufFSWorkRu4eQpH5TzavItUGAAUnou
yZ0RVG0OavBu7x4JTNeHwRCrvNqCK8tmmDtYotb+7fyscTCpI8m7weS5UEAKCOIF
6GlDLoQ1mRjkg9xwmjeydmwREBuxGbkaIcJFJiOJz1ZS1P7vDCf7Ftvi29zT2aDK
L0a6XuNGqhFxAXJkaLVLv1fntqw2HyBt3bRZbOJOQvcoVYrv/IsilAVqZZYn0sRc
I/MrWDIzY5eZUb+T9ztnR1sT4ErLNWs1pJ24owqaYFBAWUpd6bUBsGrrF7eD0Pzt
ZAz70j9jDB/oyrID1z3wxH/8L1vBxysC8XsFNmGZBYs9a9sUynMOrOiL6mPJfjnc
WVk4JjTYUgn9Tpwa7eioEKpGuRc7XJuzBeiX6wz7HlIxFuXrPKhwIkVszmvmxm3Y
/ypjmmCupcywJ4dW9lf4KrCeAJjj31/fshIVnRSRx/LUVEYOyfqC/6fJp3SNKlO8
bkAxoHPmi6mozemhykJiVoc3n0cKbkR0uwd6titSuZQP8CGhO0nlu7lnij7KOfl+
CD4OudSN25qX5jP+W2WZZb8xyTeUx03GXE7jByS9Hg7HsrcMJkHySG/moLqmFaCG
lWaR/hVjOpZmu51rivpH7fiZTtaVLWprZjTAMalXxR8f+BdqMo2fXqzz2j0Jk+/7
p/cQKZsA9EP0Pxz6hN3dWxjG4aJpttooM0XqHeCWCQcF8LWL8+ndl9Il+zmtx0/A
QAmI0U/qoQvR6xXyLd+NxHYB7dJBw06r69RdVz4b/+HWVgFsTeb6THhIESVXClCa
WszIgQ8yY4Y7ZFoBOuNwsbXVxmSCzmzPq4I+sz0a/vgMZKKd3w0UiU++u/HZ4Adf
mla6juSxYDi8Q2XqqNqHbBnI0UYnT7ZDT12FN3aCyQu4NOMgrV/jxWC8b2KKu7oP
HCzBkB8yRvDl/jRM/kTV42BN5vEwSVocjdLpnZrkBgqyCISf0+pFJtMCerPMNDto
XXBP6+rGtPQ5s+5S8P9PeqWeVXKe4XOYsi9jzbFX5OS+mf9TyPAKkUjTy8/gXXMU
au38A+ANYq/wn7Ki13LUOqdwsvnE/2OUC8RRc41JOjGrXX3wfelMmCx8qnAMHl2w
x71/HOZsoEqJs28VB8nuKdMSlIVB71oSXIxF/EivmkrR2Fpn8W3Vud/7WeHCUs/X
BMcqgdpXD7vieYZx71J7uxDJUGp7GNouExMB8aTr3gJmJNaLwqkCBRBBCthC+JEV
9mxFOy7Mc8UD23UMMb6098QlIXp+EVHCGYlIiLfN9IQjY3zGUaoPu2EdNh1h1Gdt
7cpIagA1BTx++tMqFMQoNYMht+iGDtqtQ6VhoQEHtFUja6t31SRafguKJ9D9P3wZ
h6Zjm1xfKFgxE/nkdqCs5ORk3aTtfFDMGRP1OOByaw05pEzogfVak/GkXAq3AYo7
xb6hY4sH0g4xrp60zuhUg5nIkTYlNYq0haoVbfGqC+4YMWLU7ymPygKZ2kXpMTBU
DUbwjlPLp1pHxaMsj7N74yaurK7BNMnWe/VjNovTvkH3JN8AXL8VNZxXTOBj6CHQ
8+ivlvW4BDWA9LPT4025u6+f4UA2/vVDCFBavfpb2W1GbogYJBKUYg5iv5Z0XYLI
Qo5s87n/n203v/XWJ4GwWyTkp2eUaQeV8i6+H1wd7FXV9YpJCkFz5aswX/AUZJkL
bE4bAxDDYU6WtR5xiHgg9Kfayy5gBOMjCFjhBI1RWGSQrTXn8PVCHZ+VlHlQU//2
chyBGn1GLJaAakoJ2eFOSglmF5uK19FL4ezFrWCx34o4RugnKgWt+2IOqucKXjBp
wrq9u7cQgFFMCksWKC7hJTFd2a9pd8wXO9dMWvHa43orCCMfdCFVgBop7d0mCmPa
2TYMYQKhMFEMWoF5tJSRC9JY3hYsrRmtrDNf5uCjIPZ4egx3Rl9xzCAtGKvtXEgG
bs0V/+NZU6Xx6/SasC7N9H/iEbmMV8n63abDiawog/LNweDq0JeKpJWMFsiesWsB
75+ZKG7Y+wXv4+XvJweerRxymdGNMvTTFMk3nGkUAR1x49P1CGtNeqK2OF4vkA6u
FWZYjIb46jPi2krE9ui7W8w6bUygQARgG/5T4SXgmgdSHNTOWGkqCLZCFWWAAHqd
10Ttb+EqTaEXU0wNjLXcHugkFSWe2wp5vJNnvAtJRx3MaFRfuXj3Ikc9ciU+/NA9
RZlPseAVEpK2hFScqPj5QCU+ZPAKVpaAtOcJoa+6Hh/pjcRp8pRA63x77sOPkuX/
sQPo2jT+dhXR7EW+kqpca2EkcWq0tnKNxqGLTgoVdEgcVOtbgZ2regoAxB75cBR3
gzDMRLfGkTUnPCzItsus9vABzkzIXDIEaod50/G8M8OU56QATD6dCWaIYdaJv6bN
36PY01AZjUmdPV/HX5c+geXZHw3juDXfuoWufESJXkdauBmo5Pnq/v7yffnUgQia
NMfTSUbf4pPBld9drVIi2SMocncy8knkucgXkXyskdYkCvNjjDSz8rba0LlN/WfJ
h7h88Zrv8Ze69EkakzutY41mYs6Jxi0N9TZIZZKfyskcM98HE7NX6g812YYuFSEN
LHkS7XaJScuG22QunyhBMs5gqzNgAOprEVhsi9pqdq67hRZHJmW4jkINJF5jXlTa
eRWUmUCiZlLEIxYuPCJRV6VNxjGkFCr//D9rn0143oz1S24OcMwCb9cIbp6KTZhV
jLSLVtbJ0aa/Tmn+FLWOto3QrmuCIpND+8/ntDQAKDPbl2d9MXoZQt5v/o9Magn8
wMneEqEIN23BfFyHJIsRhGqfdrR+NUygw7tuNeRvM4IfDLlf537D+enISwnJEfpB
l5J31hjW0v+ue8NzzlqKG/YKtViQxSd2QR5AZP5GQTXtdZ6I89+p/SbaZuWUYijD
g3jkR5bjWQq7m1cNtz2PZGKz7TKrx29cobiymtu1PZnZdhBmozLwiqqO9KwUVb2d
qaqPpjpJ6KL4aTdVkzeuOUshFoicLlOYUsGKeFayeNrwBue6IN4WUPfHH7bMAjvt
3OaSjYBjaI3ZLvLzrSg+cBlx19nWWFjkT5YX2SK6Vr3xoFGgjd2UkKjS0zP+lXr1
YQLNRMEgn92VRO4Mgs/wkZKxD6iOuizJ0pIRXR9h/wFCE/fbXsmuQQJCCiBcqXb2
iWPb72D4R8jtYR6IhwfXdcJWTsOCg/zi1Ri+6z6dxnOpLVVC3eociSEkvpsKZukw
F15luM395IlTeaQNW1uoZlavufme2uGzd9oto6anb+g3puNfBYwcCkRuq/zGYMCe
h8bIQ3st4WuuQsyFFlsexQ5wEiRilIjeLKDlFF1eAEdOWYAXfMt68FyQzT22r1oL
02uqthtn/bMT0O60oi9yloXp4ojg0kRqACvHqifg54vD1sUOFmj6PBqulV715ZKE
objWpEwgPd+5rcfvf5+ljTQSI2WDjVc8iVzXbGCKWWhHg5VQcyajaEwis1IeLQjk
DfHciPLDbmPWvFj35caZQQTvUZ+g5PGMZ8Gd4js3S5FUAHTqlGp/4lF3NQwKwTm2
M12SGPisyxijuOnIPSVJGma2CqbxS06+N369GFV+fvPiRX+RMSBgymhOHbqJruOz
kkWABbz1HRFl1gNcGxMDlUFzYDsA0hInNFJw/+U5iIzcXbldvpcC0pW7BkW2+0a9
+TeonURxLVOyD6Hjn0b5aIH7CY81h9EPuFkh5YR7CqDivCs2rWXa92f9I9m6Xxuq
KLpokHQRNQET1B5qz8J3/Pma6LrUDlmzxQ//CCQNeZRONGkhUCJDHe5cHva2BMJv
W3Ub0EPW+RLpW4xvQI0UKSLN/BLVyNMiWeDiokPeAfYM8XEYDjzpmT2mvdK0Vim5
r+sk8y03WUdnCakyZlEoeREx/Q60FEWQXjCvMNdmC7YfDYchp0cPaU5AbWfk8pjc
v+WkYWnGL6p41DZaNwlHSgt6eMafrlwY/5WiBKxwG5RvUlPnpY8Fg6gouvXpLf1+
/YhwsM3cOpLaOY1dF+NJyvbj37g8gyDiED+Mr7bgAQYb+VxVC1ECFKTL1GiawuY2
ZT2/Stt2TA616o6V+dPzuWzGqm4yv48gvTN8LWBocoPXsW6ew4nCnBf4wa8EU9DU
sFK7yXuT4AbrIUvsiSbiBrseUUwyx/q3qgAoAbppgQCj0J+1ebcsgN4aPnwy15WG
c8MnNdH7NFLfRO3rRKqfTPQsGJG5ZrgW04JBxP3uPa39ZHgbUnk5ypiuSxoMqzVH
LirhBbMTdNNCpo9pOiPuBQoex+tk/4zKDSvQwo/cxgsRe5Ljusf/X07fMxOCcSQm
K6aL1M7rIN8RQwAFmVMjhl0lWvX+sagiQKObTgl/RcKza7WMzOKPFzbcIZQZtwuI
tD/XrReiHq7XiPb88yXhmDmv4TtI40GdEIc8GLf3k0V7CeTy+776hxLKoujEu3Fb
L7MhGKR1SAthaPLxqtJPxBfZNcfBT4nuZuFWnJ2lLE9E30xgJovnHgGIX9Cy4TlE
Pye2EdBmoqhXzpJLZao+BiYO4Qa7HTw61UVYOLr1JL5cIJbaZrOWFSewF+ft1nho
ognRm4oOZxb9G5rUZepXF8GXzgkBGEb0uE8u7mrBAf3JKVAgwBQf6Ns5XBzOumJM
3ScwXE4h0faDQMGWoCPPxogsVKrH/9eBesMh7uU3YDiH1lVZrZmm772zp5gdfFmN
34rbTx+rpSzXfZqsOIvny7rwKyv0fNqws3qAQbuc+VlvtszxPuwrtOgSb0OIVQ1v
CsU1M7oKiKzhBlQqJ43wMtLdjeJqT9HbI12vLx3hq7xcwcPMVwZ+TX/aoZxqegYg
jRhaBTMCgnW0aAP1dyPc/bqjqk0qaeGFZ4MoMvmem3KKLbYYVGm33onu0gvdPbO3
5DzeDKnh0OI4C/kyoeFKgl62thXIlDqjAdRBpRb+mguHSp5TuSIXdpS1PjUHVlLK
nwZFfvL/rq8dfEYvEBw0oNZOY1wYTD7Y7cDC2LuKFpeShvzXymt6UOid0CXEYGC4
HRsIVI3yAI80jaal30n5t+2foTk+CM4PghA7bh6sQZ5jIZf75miw/JE3A492dEZu
TFLPv1SP6bV2KwCIPVCCXvoMPUvHV2FWPYXM38pd4lSJHhn+p6aMQrx5sgLYOUr8
vc8RBofUcNW6APmXc8NuoUXr9CkAZ+eL5o0Zo9yCUb6/0PInVqfntZasCBBuBpRZ
F2P1Gc7YurETaAe5PKpIZhJeg7lYROXnynkuUp6o7Z1C1vCeJ48PWYnxJU0KC4K5
zbtKV6UxtYc2dzPIa4Sxp6yWVBhEpyJvxoa9p9YdV0bkzi/DSjfl5IXani6Et2EL
CvvYkDX7LmGhWMRYKTEL5V7LzNHY0NsopBA9Zmc5Euk/7JPM2tgtqA2JQ3rgGY4O
KG0JCpO5lZE1dwDwosr7wIwalKiu76+AFJ0ogkgK+6HNuwiK0ido9AnKQHTyQIJq
vNDj55y2H8Fl23YxDC+6CakZoThNXn3/+9YnfPvg+arPiDy2PjL78zCxEsUFz486
jSotBlLH2ZFQbgWRKbNgOPqOKMmt7EBIqGrBaeqaMdsfPoz/SdqfnoYobSLEUmSK
lASmj2auCBQAWlW1niYgd7QyWBr/jNBW2pkOcpD1dJbpqZeyTwfyi71uzfrct9dw
DHxroQO1tlb5M8z5bNZaUSnxiQCCDftUCCUIxpIppFUJQsE7z50AVxWV5T8saFEz
OpA71XGPebQ8NmCgaAVBs+fLwEoAt1GQCym3zv3T4MMJ50wllN/6ZtTKRvrSikRM
defmnYbVM07atYDDPHo0QUshce7fsN/1HstxZSb15xXmt5YOrI19aSUJ3faJ41CM
JALcU1y0rK6qOvTiXr5qhoWSYNAHCjVhVTnENYaZLfba8k7iIwLC1koedHiXLwLT
usg0jlkr3qVKrRP0hifjZvJQcvq4R92Rh+8E6ys+nHCpvwRySil+jkyvDUNnfla/
V6rLlJ70TgoW0ngBys/vX9KA63P/3cirtALl0d46yfmcBVxzjfUaayqQ4oT3DbWu
UMQe+qDfrCEZLYWW2jRs4iVmBbbTDZ2y1iDbIwlmnxVcXyEznrJthoNkfau7++Oc
FFItKrvjnEgQ5PUUX0TT4uI8iaQ91vGvWOVcf5DccnS03k1vdX9fExHdFb3T/m8N
06GsxeBpunOP66CFN5rihVG2c9Jl4hQoWjBM0TRHZOe5+0mBYHsJFBfRYz8mw+jc
RTSMJx91yqTPHwv6mZ6eWNHnjpM0kxz4QnMaKOQa9VOpmLQ0V2FGsp1a/WIkV2YM
MfhrsdiH4Hyve7k8V9r0aSTBh+IaT/iHmBki5f+jblHAu60o3KlWdJlyQWJo1kdk
qBgHU2CG5zCHd/UxoCqwIRqcrVdh0BRZmx/7lejPl++sCL23bz43+zNu+BLvWAxI
KSWD9p0DgmEqUCbjvQOFjCAoPk1Z1+nxTtkgndyfFGWLBtvqulQwNIjYQ9v+nY+N
xM21oo6iKtzaYv+DSvtCBlBExcqzJrzgjFJE0HzCUTXfEihOD3aeVEp1XnMx29B2
hNsiknQeRiuOBHe9bhFTSUBPa3jbKbY34UFU+xHn7FVecufdm8JgTw6z+L49vEbR
8W97SNFBmMWf66xQAOK/NbnwdZeQSkA6f1FJZSqmMI3Oyf38I1JJg1bDEg10uFu8
otlg6lC9t3jOAI5sBbSLkZw0o8MtvEAj/EI6xPoY2Lo2f9IkYQlAr6OhzRJST/dz
7OeHHcHhhHv0GEhcXPQMIReXM6IIpkUmQkGSLtGI9qkgDPK9Vs24G7JdLLtOCPKc
6rfaF+epGkTN460cnBCU9KTadyiFjtEiRe3eiFBxYfIxmo1E4Ys6126T2oUgKDaz
1Ak9rsl/neZkV7o+AR7lXQ3/8CD/TlyRey3jlS2dhoL7fjeZt6OsIxrUVFmFB+yL
sZEYt20yGbgOBWGrd+gQmWtHgUTuIoPg6/J0BPt3MSYeaZ/aEFzds27aGhELonbP
9AVnw+5+HvVNw0EO8W4Uu1bLpBnaaoRCZaIAvYhVUYllhq/eCXi80CnPs1FG80xm
MlWyXGRnZqLTL7zt74aRklbDdgJHbiRFNVvLgIXcm0bBzbZm/OdTYxYwsNvUh/0Q
Tq3ZYIjy+ZAa2GfGmpjZmSMH0wYj8slkZT41dVioiZrcKkbr5fcqQFFU45njhl3V
YXiR0IpQI0vfjGb9Gqd6zYV2twiPK48Gp6fBE+rRIamhhPRYJfnBw33ji9P24/UK
KWF5oF7ElBrZyYLV6btnMrhkoQWUzXk6YOH9zP96dxb5265Z6QOuFMaX/Ozk1kqO
Z/QJmT+OqYztazMPnFVApui2yJb+NpBzR+ScptdgC9mz5EDpOBhquQT7MX8YRCi6
GXHxwFxHlwWbtvfgy5fL6Djx7whAKWsjc6LryUAXFxL5nXfnJGqgVRBWHJXAviJK
u+ZppYRCjYBEPemrbM/FEFe2F0/bZwm13H/TW5kcara12HjyKxNI+w+Utta3E53s
3067T+FhsAygtGNNxRLWcY8zzIgTnvg2Qn2VFtGQNjQ11XDGhVKYBXd6FXj60gJl
rBMDfo9J0Eh6XDcUZN/IoJROy5g2Yduwb6hO+Byk5IsBOxcl1czf5ru6mGxtgp78
zOk568XDyvlViu/JS5+uQczUkSLcVo1akDBeIvHiHfbOEIWEcwyo0ItR89Mn7bjb
KC9L0dYbSZjiy9eLSlzS0qo8Ly9WbKs1y2D/KksYIG9zrR4klzO4syDGZ4TEMKz/
8OZ6D3rRkUoq3QwiZ6+CEN4YDhDMWtnBqTG2bikXYd8GeJU4ZI5km8FDyP7llnz4
iZmjUzNMY3JHxm1SwkMLLzelUC7XubRBxe1Tvqs0f8/F+tNKTIUNrvIfJNRdlagB
J2s1y+CNgTaUs0TV1OXsonh/pQhan9liX4ymW0BO4BB+z9xGPbIaKSkgxfZYvLv8
IcK4PZDRgK29bfoAk0V5xTxGD5fuuCFH8dfPCbFjhfe1Nr6ReH+sMxGn85DIP28k
2GRBywZTOYXEYqonPf6PALqGiJBzfjv0kzf3rrmxOjCV7tcB0ywnUFDw2Mvhd4nm
acCNzLyG4JFiSkynpnMj5fOFNGb9iW3R8yyu4+PgxOjlGk1gW7fuF41fu/zo/dwo
R9l0RODnvkT/U//2NfDJ8ehGEhj8+EQl9eOJHJVuimm4kozDR+DIBQT5/momIYy0
dVIyG3YGmA8XuPUB0r9yBU5Xv9blXlOMLThjjR2tqzRstzqiSgII+hq0VEyJoLnR
95NtimPKTUUFSAqF3ttuWxVcTCyA+AgBMUZ2SxXkHiRK1scvVruhOj5a16avJpfg
huS/J/mxUv3QxvRXGqQCTYtPzEZZ1KLZOkTUf6uhOgNdWw6TiJfBspP9BXx3qjbA
CPHhUFmje34Da22yOOFVDVTBhwI4ZNa/t/rlGaUYZ+btP0h8CMwrArMTN/FsOgas
4IMtzi96MuCLD01BhAtDtu/T2fcEEM5eQjl1jwXHO9bhTzv8WRgIZynEafkNscsK
wswLc5gMZHmQBL6i6ISb797whYDOJX/72Mg17vXfi7GVeeKhkj/s5ne0z1NcaApl
1d353CaP1tDY/4nVX63fwWF1V5kQX7MQ+TOtg6psWsYatl8TqBtGTXYZSyVQYTDa
mh5C4IyI7qGTTZ1EAqWf0nweN3pt6+sGxSodydt3Dt7yXMo4LJ3HILwsTGj3VLl/
Th5SwYjG8OOOpuXS/GdLNArr7Pr2hjx1OqU4qoWDAW41SMtvqtLxqIbwR5HwSRSx
rF2Nt4wnUlkKvYWJLWMegXiWV7jgm6aGa74xBpXDxKVRmKYTPrVnsumMP7VdfiSW
+TK8y56Yxx8ZI+XZwcSQJ1lDmgtZmt+fNExyUuZ4WiNLX6csSaPrirgFmzt8YFzf
K5gy8uCcMnMZh2Vqj8Wkp+UQcWg0dzqDs06HYoFEXaad3bg1afTOxhY2784XHH9x
3KM35mydtUHmF1p6lTBK3wss7FvNpgigjoVIO/XWxf0zewZYkppbEylz118RiMQ+
liRePlaHBgI3L02zz4z/EWvx/FfK4qv6RUE8lLeVt7U9ruFpDk5kYRKmseCk0NYq
B/kTh+ZR1gE/F2xxE3qb/a9PllcvzpFnWyYjVAyPKk9kH1gPG/cuiUvbruGZeJ7i
Lb87A872hbBBafMBjM5RhIYGrCDCcCT/zw0BN6RMuStsB5dHQjpPno7B1rn8lXic
6z2af++jKEf3Wv4iFIP9fN6B/wF9DrQYkVBTgqDQ1mKk+1X63eTGBTmcjBK5DGlY
mjtdiQBufHg9uUd2zx5JqU1yrFI80nKUpwl9VFJr9oTTyWYyEdVL1NU6AdbozR+g
LkVva4w20xuUXqn6qFKOMM0I+Ml9Gmo97BQVVlpVIZiF6cwvo8f+WC1X7OC6sLOK
ZwocJ56RIJMIm0ds3ZLEPETL/hahbEWU/EMSaylll6Ttz+pejmXn/OcyLqKvOjJD
BJelp0vyP7o5VEgrD30FV9PcEUDXNK+L4I28Q/u+i+09ZWuN5cEBms5Gp0e5i5KR
SHKzhVClOJF3jpZpU6Ly0kfaN0wWQEmUuQUdS0/6aA7rzDPUW2y/01EARb2QT9R5
0uwHC3r10VO+ZjM+kfDlHLX8JAO0RfjYSrBfF2sqAl5O2OL2OPhzyKTotIPArk+a
MbNxhHcfZxHrFSY/a+eyMJ1WlLldvwrdUZpSv6rBuIMbSLNXz6nDcoTlH2AdOAxh
TtZ0totQOx5HNcYKTL1yiivQDutTO5MvVNy8H4TzpuuVVxr/v71JI1Z6Lu6MeMwG
Ik6wXzEdYKe6BHr6KJiPnOVGwKEOjn/j5UQ0SdYlUnSGMSGWqNVmswu9Q7AQlA14
bXCTw2e8keEyhIkrDuyLgg7eIQ+ENl3S1Wmr6wDthySNqmu+lJX4ND7hn6h7LkjK
Weel9DucsA0W8xbMoLIRXejRpWAxnDImqsfTyqGZubQHiJXnPUkgK0wf1yJ7Z9Ya
mGWdGAgzcA/G1JhJCluWu8E/minQmqpTR+FflLi6OZIFURq/a1lNvxJ7YO//Uhli
ZD1lMNQUtbRPg3hkWy+R6kibw/GLhOoYJw4JErSBzyVP7vQeTNDVU6wL+gju7TYn
8GuPk7mSRWKUCIrQZhLIr8ktmF6pjX6vc4obeGnZpAKEhhe6vfvvh5A9FA6FagFY
fck3d+uBhGoyn2ojkyHcSHna6Mjj2jKmzW4b8mEFzyTTz0sIwQjXMQOoiW4JTzyi
JvO2Ep58UWN8Hn/PaoJbhnLf58Nj7wjAbNwK0GNCiu/ywpMIkU2/jdCmoqH5ZaQ1
mcLzgf3nNuVpg/y0vMfGm/RCYPPwVvIwlnEYdFs3HDpXBCAps70FedKJon4xufXC
xN/zGz0Iyb+1kDLcUwQKHJ/LszUFKJHTQ64BRFPq8/I=
`protect END_PROTECTED
