`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
y5nAakIkEoOUdNBYULfkB8KwGm3qQgVtn/7Hqag6Isb+52Naf/6nfuCfiAXXntV9
ibrdT3bR6GK8f+RuxCju6ipady6HiLVtnl6dA2AGuExDgA+8TeTkTQe9SZjschIr
qQi/hkXDxI6BEfcTG/iIROGdUJSscsYgTFw8Ng9+wOHJzaiT2uftGQB6x3y90bMh
eX9QLle7g3o6vkMJJizjSU6XD9AKxNP5h2NJeiTyHcVth0tMMzHga4oen6maILxI
nvoxPqmYxOYbJpazA5n+2YKVR2AcX/ZccFHgkyIg2G9Zjm+3Y2klIGHx6f1l5voQ
sgkKlTN/JCoEIryVq3AJkHP4vhnaVL6CFCy7zG1z1aw8KEu76fy92U4Psz4b7Fui
vB03so8HqbY1al3jP91L45E6+gUORCfGl9w83tAZ61pJnmfek7MrcmXFf8WYeaw6
Y85n0zNpMMZSzAYmVKGyOxvqSdHVU3jhF0mBfJ1G9ccTfpbJb/LSi2YrOk0lOdMs
q5H2XIaj1emkpADXWDIiI4XOXIyofsGy7zjp8icRmw1Pywy2JtHuRywoHHUhJjtQ
Av30iiFd6flqUAOTW05OeLiAipel9XRjdVYW9f9KSUr/sD12pz0+H+wgNpdjh2Y6
ipELXq2C/i8rJ20+aw1soqeDd1bbW3rwxYnyY63xPMn+Kn0kA3Bya71X2/Zs6YoV
369wNexfHmoRYZLMu5uLNwdA/KtchVeBJ9i03QyrVxWkJQZlcqG/VNRRY1YFPvuu
fWaU07LjWg2Wf6cCjIX6gU0HDmZoWI7Zw9QwcwMM0e8S6Oarc33t+ZRH4K+o2bYr
2sD409xqfu/UukztozznXPIpqeDC6E/Zg5tDQ+wZEbmpE3ZprcMNi13DnWZceDwU
XmpTusMS7msUBeTPaj58We3DFOgYO2tCHpZll9SWGHkU40M3urqnIt66JLHZ2btG
bX7CtkK7LgyfvKSfOyqa4cZSaHLbTrTCnDMUQhAqD3ffR6W1DbGbBYfHKT6mHwrH
qEwCFbvBuWbjSc1nz76UR9ZK8iwP+sbjLNBfCbWlWE5JWLari3pG9fYzuFHHeEo2
j+Bh68sfFsc85a79JkHpbo3/naRwWxenKdygjB75r/vAdoP2dkfBnOcZ/q8hSgTK
T6gEIyCbjmtfvoKq3mwz0hJLY2QwaXQkNykGKrEuRvRwoKTQCmNojP6WL2h7Xq7g
anClOdEH+HP6FHXguCiSGP6+WJxhmHH7HCbTbU6NydV04WR31CCIyCXQw6x1AYF+
zQmVf5zsNIxciiA1fx6mW3ZQ0oi2F27yRv1KJwjer+IObeEZiopc8JEva2HyLhA0
IXWI7wCjVJ5PSki1PgLWo3hNsDy/EocPq2RCgjvkyagJvHGbxCXHvwATAHu6F9iD
ALXKNSehkelydwypZNifxFSl67F0EO/CJ/xJYoGc7ZOdsJgNIqLjYLXctk3rA3KF
/A0y10W1TWCTWeQ6eAIw4BA6pdscj15mlhVdrCzecAiPt2awLYJ8RHajqwDPmesB
nkvtePTylD9ur/GCqP7DWxK6JJ5m1Q+AAVpBeTpRbxNERCqEGOPSUuF4l1c0E2rv
ik8OYjwqOrkK+qFclrdfObmCd3oJXeAKi6HFM+rkWEbidwJvOP7wz+yZxhC3K9BN
uiYDTn7jt8VK4bx0MPSZiJixJ63McOA5nqrQAT5jFdAa10YFrvRTAn+aX9G56TZ5
soSJElS7eLJ+MehL0rNTOhz0dQMGK4PzSubVTbmqnm45mEHxai0CEKXBQPQdCSWd
jlQv3KMxQ0210be+e99OwED6A9fVrsjwl1Gbn224Jx6fiO02YSRhJ0Q+cZkQuibd
7rhzZiSEwl/YFIPRfl4Oz1e+oJcHJGRdYHcGUYkIHGEvvjNdzJm6BjJYWQO+TVZD
7iST3pZnI02zI+R5AvxVZziCL28Qkm2I5K2Q9ZfWHfIDjTbIcHWAEeWqMBPoFBMO
kzfw44qerWI2dAJVCoQoqsTg4UIFNjTaPztJtGCQjeA9bAAvd6moRsUdX2fheOfQ
/5mxl6PWO1kNebmjeF6pBQcQVIgLngsyOQcNJwkSQ7YTGT65vG4peyWeNBMr2HU5
z7g21TnzailIyk88jx8zI1xYStbFxaCTqcNAFIau+4YdwHsD6SxAnSVqCcf+cq2y
Tc6kLzGIwodPO0HCm4xoRkrbMHnuuVV1yrh75H9CQRK9Jm6/6gy2dKipd4wVH+M8
rEaDEf8Ds4a4y52vjzZtXx8Wx6FZhBL9UUl7YRIZP3yqelS+U7qBOqzt3OP+AOTK
7UFJccFeTkI/2VPFCQhgiUSa4gQ+pztpedOZO6yk03yAiswuUB2rUY0MHLsy2Ep9
rV0Xh+tXY8oMdVQXNGznu3dUvtTTkzZBUC6oFurHoN90Lp/nrhRWOmzKhwdX+HWV
OzyTC1WFcXDu0OBYMGafL0qEZN82x74Cv/hqVBIViu5r4GufFXMz4SDIp+0wdwrP
C24UPIluqB4gWw8cVPYa5NVlTT9+wTuVwF+/tX7bM+/YKm4BagsPoyB1mHJx0RTa
uTRX2K14YfOUm5vRkGTA6PPYI7YtHCRfb1M2Hpe2mv3WTnHoYcjte6enbvW/+PM+
q2vVyfcy00QOt1B5+MIA5R2TEhw/dDAtc6YzD4QvkIOn13/kP96mIOm8j2DeB+OR
LmO8Z04NABztUMJVxp9JcHo31NjoRv1CGrtvKJ9cpHR2hBzoWWMBxT2IFsYnnnr0
uiIjzsV9Mf507r+nUh91yysVTkTrfkUzD/EfkhKksM0=
`protect END_PROTECTED
