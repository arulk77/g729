`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47GiR2qIzPN8YpL4dyaEMdRGWnrm6GM/BkK8OYcQeRaT
/OF44hAp4Vdt+La9Hx746JlWnzjzoc51pA/A/nc6ur3BBPskGA0LjSN/TwMAeJJa
dJBkt2r9/Y/QUwnyHhpj33uB+DFLZwrO7gALKX4OmioMZFX2u6WspBB3V54+BCvg
hlxW9Q9ZUh1+FxrRGThykVL33LKtEoSzNMon9fjKAEADlt2ODTshuyUqV8UQuxFH
cx3o5aZgTBXoRNwGIFvgr5GCjzsclBY2Y5MDw5RBT3accBYNF7rZNzxr5PUCpLLz
wTwZcm2VazGnd8AADJXp8GSU6oN7fxIXA+8RX13kZEgIlioGisre+f6Y8/3aiRPx
dOk71FXhBsuwrgT/CmiqJKLY1ZNSuPZiWw+Uj45+sr5Dd8RBAlWUUKcXSaPYuWUm
pU5VFVvmzVZ0gxgCLd3t46saAFAMf+coq9L5wC7Gytywq7gQplm3mXbkCTQmcRNu
C/pQ9lm8tevR9vAHMCpzNYhECLgE8l1kMSbmp+JwHsLKvI99yw/omUQfAUMja+ax
ncVygrcfnMzVb86JfTMBAZ6jtjUiWbmRsjrJVwe9mNDMhRGCWCenDhAHh2+dH+k8
hz7oZdSc9nOgX3XoC7FF3sIWnpGOWGRUoHqbfNI8uun3QRht32P5vnkBtB3BZygr
Rb6C7lH9f54Yn5mWuyx4Ow5/zdMN5TiyNXXm/Bx8a5LGNO7IPHZOxCRdFk9/wGyz
AG7ifxsNSfQ0NKaDFW6vRAJCUcYXSX4IQF3j6t3IqKSLq94PxO9xUfAGQPh5RPLa
gHsLZ9Y227U5e2vr2onnOHcGx5O+OBp+wE8oFpUL3u9xrB/U0SN2ugrme9jYVrhs
BmSo4bWmQBIePFquUm0i3w0d41kLZ8iZOgfvnl1lDpP6E/1DlMwXM2zYtP3Vr1Ls
iPKDHslly6w7EhgKYl2PpIRNIHDKPYeGAzxjl+9VFE8xJRs6ZQ7MnvMcs77HV9JB
qgNZHTAhkAs7XPM68Fkvq3vxE4LrgRVev17tCbzCRHTGfAbnclJ6s8Wwi1eQ7lL5
cxy5gFZsbXjUEpMGFAbUfdMWSeYNt1ni8xVokKij0xlqqkoUpUAJ+TbX7QnhKSll
/HmcD4FLk+qljvXSyZ6bwYtQkRQdTkpfoktwyujk+PaS0aOSz4ToRaa/LmATQfvY
avDYoeU98Ld8s3IsGWwEEqF9QdFqV2lDELrWMPcb+jPBc+AGww4mJS9tk8LTtao5
pbhkZj0iEqB1GR5KFFUSyDl4Rrj0YCbKOV+8n6AZSJcdVLnvV9oqoDgib634KET+
8r2Y6XfQq15nQ45ZAIgEhDhTzlADHOab9aDM5BpqPXuOkxxqFulGqUdJnrEWQIrq
5xp8Oao5fYITlMW9r6brp4o5vK5zWOVRp2gLYJ+/enQLpQTHFVxcjMUurrcfat1i
UpOwm8AN8paa12Z1H/BLvXBzK+Wkg8CuCnfoLmluKgGk8w9srF7FQd2RosvJnZLK
iBbq455GZjSkHsiZBlVDCTqY4GMe9+JoGRSP+gF8g5gCeQpkN3kUxCIO7QSktXg2
2HfPVW6/bHp5TxA4YY/zGTXEtzR0cbrz6eD0JkgUCa1fAhtBlCf7odhjXVtaRR8v
Sr53Fn32lKZklJSjDg65oYOg/pbmyrVI0t8HA/uF93q5FceqNUW9RqNmzuwRBEhZ
Qe/5B+o7aeHg/0xwTh+9/smP1XizER7RgLkbv4GSwD/tcWFbhswlNaa/EpC9QGIS
auuZQhH1/8+lAI/Ne44jfqtvqokmfDw1fxOhDTSSIgdMP7/9eF05TE8GhH1NNbca
EjJKynPU/S5hkhPOwE4Yr2dGOQdv6ZVzFxYj9+I61Jrb52hUN4kG/IJOiZj0IK5k
vYoMEbJIFPqc9ev4qDNygPFsperr9Nm3wMUhYLeqkxwJpP+3WA6kNox+ZEWm3wbQ
LggTx7lUUDiO+pDmtAa8y4lqgGnqS3iAeWanagMAagUPJI5cSgNYmFc06xeQcvIA
g/RKq+bbD4HNxSq5nYzAnbCPmudUjPWxq/OMsWUvhEx8/jf/2RwFZHuy6tpzCG/P
RROdw6wkak6XDVT4HW9KHEVhQXDzlKlq4zMwaaCnyxnE33E517bC6FzH38rxNIW2
cnyD6S6aJLLNHQlEomKZkVBn7zLg8NvtBTA7EhEoSmSHAjunyuRhyo8In3jmm2BA
DsCGDIwMYV4hbCIU7kAtFyC4qhMZPZrGGyTEujvXAM2ahKDqZJtgPDJvmBk1Pf+r
v/PsNfCQu7a8GZ1UghUe72iNqDPDkXshs594YjTu5XU7m4X8nTrgIM0I4m+vUJGx
DUyCoDuFF3CkhCal4Cv4ybmTgZbzlcldNxHL2SfkycKNcpkjCqjfGEWNI7DrAjT7
yo6VSsWfBkMND9rGZYiahTGgjVm0d59DXL9LEnfsLBakcwFcyYJ5wAp218JotcGw
x3gbQQAC6k4XSjztU97hAVtAg0o8gUl/wLpuUdGcWcmZiHBCnWpz5V2T+U7+Txfd
Bx3fp/sHat+1ZidlMgt5pqdcLneSOY2th0xhPk2Qr1Pcz51XmERXcVP4L5Q/DU12
TNtFOLvzoDT85djLqUqFjCdM8KxzVge0mk4l3XK7qQEDlh2TGRuicLEPz0vyHp6Z
N55KlOtI8V68Q+0zhDh7m6s5Ff4W6vl/lbtSM0JuGw8DpkeXH+bsgF5xWbb6Nl9f
b9E8sdZUdHVXS+/fuuJie9v3bZU9atG2hDlFFClAorAbXtjpGRc7oeJoSsUZLmUm
Xhl0rTtTXU55/2Ypcu5dsA==
`protect END_PROTECTED
