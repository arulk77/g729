`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP7Jy9M/WiMqEDs13kZsqE7Sz0gqhr/+Yvv8yqJjXayZ
qy1CozVwC9uRXWTj9Typ0qdfSs4hXyx5ccLx8BO8HQ9txMgFMPmKXHxs9HRpwPIM
abY/zlSS8fOQQWF0ZiVAoU28AWdo/25EY9dtJGowi+yPrio/+wuY4buZiiPxFrkb
ufpDOfokkK36fIpV+hfJiEMoZ6GjExN576ZwzePv4L1B/JtBCjVJjhvdtpxGbM5t
FX5lf063AX0QWJu8MC5FRI/bNQUtxfZFwPhUb/OHuJv/3trmCyAXRUnHEGRnZXK0
3YdnoxIYPM69HzIV2811zw==
`protect END_PROTECTED
