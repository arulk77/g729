`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHq1Wyrolg1H1ovSky9LnKaxQboLDocHddTKKJE56j37
IYeBDcs+vGI5mVIslE9WiY+QvFXmlJ/XHFoaRO3YXP4S94gHzRsYrnovDayk2lIw
44BIOZCMKE277VUW4HRqcErd+dQvC8eE2bMIjisZEfIm80e65I2Xe3l8iiMWA4Ub
`protect END_PROTECTED
