`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveECcthAeuo6AMCaNLWbjOQcrZ4Y1tR41nV9TcfAA1FKG
M167x9HQV8KCdeKyOmLjHKrjvmLOicqNI700qTxvV9p977G+5lrHrHkQSpFoyceG
dUy9NYv0Q5sriXQ1wPiOdS1FnCzh555bcipGE7TEYQm6kV7oMiV+IaJkQe8tBsZo
XRJ9c+eBWytVrJtAdCMI6w==
`protect END_PROTECTED
