`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
xXLmoGGSVurXvsofX0aY1sR8hhiGr4pFI16e1F3tqbc4GeHCE+TH/kiEDq+RunFW
BniwGA/8xRUe+lmfDwgtot9rnOw0zO9CGwvB5zaSQwFsDRTl7xTvFLrQvklPLnQ/
8MO1XN8d7jtHak3YJkVA2/y790MXwq0jGSjAEy/9PQMzAxM/p35DPMY+qaBwPx2d
ltQ5WhKwR+X30ROVHQRlTyj1QbRfJqnRBwahG/5zc6A=
`protect END_PROTECTED
