`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8Sdkc/lph7Kcv5ukSvsNl0W+uQN7DjXGn/7CUp3UtoY7u
aGkLeaJraxOBJoe4/jJBE+lN9vrIs7TMO7JpqS6QSLFdQ1svJegcjWcx66AtJCNB
8hzH6uoQkFAqtpS1caHvsrkInGtpo+ipoTjFAnry/Pb5DAvKdD/76l4K7F+9rT8s
NfzPvau4fD36CibvuPTVbhtt4Kdh7TWMhKef48j4NWQhy57U5/G+aifMRanG00wl
LzCe1d9HjMx6d8/44yTxXa1mf/jDuKBsDaEmKQOFE8MaHx+gFbmvOwDiG11NPqNi
fuaq2TRjZfUVHFz3PFy0UKmjF1NYDq9WgIMkk6HQi/ZsGhy908j0sbsl+DexAn6W
nybOm7OChOaPi2sg7Y2qRC5PsXKpee0URM3SJs9xUccgMiLTOcfgPqE1bGA7aOyA
rkbm3OyjyR0nCf6sAB/MQPYcntWWxKEDeZjHGDCL57OTUniuB0XLa3/SCRMlPVHk
5sIdLyC3YgformswGCf8d7YAfJH4Xnf/P0ET1J4AC6AIjfZYrTDrQxkzW5RtjxHV
eOAdB2zfQCoR4xO+7wEC8WR5P1Tdq45dvUmVXC9pruSPXivZtVJf+nTYzT8VSGWk
OMvJQ5rZ9PS/t+xysq/THP8rTBWALl98ibJ90Z9BdOxWdHjUee1M09r27hOap9Nt
jsAPj7c0xiZqQSwsVX3MYdcqZ58a4K0Q4/3JmK7z/DI2rBDPLl79D4sbLGdWBFjb
n9ZGGRiKe96cHls4bm/sSzLa1YTUeOSQIW4h33eD5Q00C93D+5LDWiP7nqerJ2Ir
0ofchWt7RxBRZIp4nQu/9E5H13gdrmC3wCpgHijGQy7NY7kfxAxy3UZbNRhDAjEk
6+S4Q5tE+YNlBTKf4WGw4SbNTylhQGeupPouLFbxRAFOEGclxoBpcLtWXpZ8NHni
GVc0OkBj59KTjsOiZsSsZUqFXMezZOEnDCfVMGyl+j22+bIBzo0ZWvohpaC4bGJw
WBRZwajREZkbhGfYL6EkS8Ng4PMHFhCeCORiwahO0ZxQiUgmRwno7BaO4eQAkiuA
tE7Q3w1y82MCyVMO1j+cf/iV6T/+LitqbsZl2BkRERiZ4ggmbbaKt3nkOgyDZun5
Ett0G9H1C7HtpXlBTbSvIlm4AYo1jkXL9GvIrm3knLA79JCxwg0g0H1etHI/JC2H
aEXPVEND0wk45uOy18iCUZ/jxLQ4i0Roypj4LgAzlc61tFACXlYFRaIx0xjFUloy
IFDvSXhI7aVcqWDHJog7XXOZtTt3K2xNTX7VAxO63k8BGA/hclt9e/Ys4BZaIzft
X2r7CZWeC3gsll9TwlPZiyF3Rhdal3lRJUCbem/Bmx/XJ9Fe5FnMAhwov87VOh3v
aOmiIfycMcATOkq4Z85AYYhC2keHVT0oXoHqkVwXFwdgxfHf6npMAHaC05AGm3I3
q3hB5k1aw/pRAsVj/0eIZxaiBbNDbam7sDlVCZ0HArq8mWB6B4jtUtWDomxCSq3S
eA51J4oo+Ai+GStLKJV8wYi/v5mryxaZ88U8rEaSWeH5r0JX/eDiTOhz9ds4I9lE
nHc54AWV4qib/MJ9qVuOXQB2LcjsL+Oq6Tt1T2jpfTI9h048Qe21KbV0lRhtEwmR
wWv5ZjrFumpKtBxMijL+zwpua0C3DgWj2GLPDcV7e2mEt/3brWLkgJ93MsS4/h/Q
4GX2kiQCHcQ68Y+uM1e0a9LNsigLaGDxKRbvx3ldHuBY35zR09+F1Mo5PD0+Hhmz
3V0iNDoL0DdHvL6RlCK7n1VAL2A/oio7kLBStZIQZKa9Ra7BmU/YlyRa5l/NVIso
dz2R3jpz0d7seE3OrHZk8Zj3IZR42BQbgh8TVpmS5qAHE91eRWQbTNxkNWjGfRbL
+XbFQyAdB1Bp8aUep2yEebwHwCTV4c0lDolAH492R1qfK3abEzDcLUspU1F7AG0y
nSMY+hI6ErsCyoz0qjtRea74xJTLpSZjciBHgmMDR/zxTkg4VBg3MhLTl/yP/V7S
YnCm64EGaQq26R8FtmNqMy5B8GbWzAX4uA+6FTj9qxziaic39EaODFNlsUZEEEcR
i/aXGCE6BzSM1HI1wuu3B5my2MB2lXZaeSWJyl/RPJ11niZG73uLaUsFs6dBvvNH
5TaIaaVP0ksXv9pupOJ+upjn2bKxKw/hBnGIDGxcA62Tf8Deepggyw8NLiARS4VQ
ko+s/DHX7Y2u7BQRcit30Tkl/zVbqCOXT5Iyannb7x3/AWcOFI7E7EkvN29PnCr3
6eeXBgpU3t6hFye8Z8HB8GvU7Oxna+Yrvkn5iEqCuiFFkmyJVHdlaHQWnGIGfZFy
W9to4bTQKzgpJ/6Q5e4xzBhRfLLZvKRT0tbqmGW47gWE5R5n1w8nyMX3SaHw4ltZ
D8Zw4JtWmDVySu9PAmZZEaS8Y9v/MGf6iXOt/+9Q3f6HcOGnO/wGfFSBUYwBGohr
stsaXHVo5d0bv0aDQlzTBfSpfVbRmtLe+SyzQi6tYg78WnUJBN9bNtamhY8GRkKm
6qheZVvMHi3BLpsFuhcBTCn1p+B37n1GP0bz8NnSg70vX4satELBkKWAMHZbfECk
q5++4t19X1N7nkRqun4cxk+bQrOwb/Wp5Z5Qscb52JiUlBg7o6M1xDR50l1QnG3C
8/pZ7HVWBXKcRaJgVoMP0Qisq8L6Ow+8REveG1WrXxPnnCNgCkEQdmdySdaYfiet
gEU/7PhwEo7cUblpFb5oIJef/AEGo9vB/W8x4Uwhm4LaWoxsI7TK6GxGDdaCadXn
L/2fzEqsOrzr82ZBT5bT9kDsYTEDzF+/bBYzm3yuzwBVYf5xCH6ZIC1k4RQoA1Ll
n6WfK3Sa/lnK7pA+UR8aMj7kKekmurrLHI1ybC1cMf+KnnWnrVxq1056u7So+cjw
MXLQzBCrzTn1efsys/wn0SRZSJlW3MvntOhxD3zplOhbbZP5AVDgJP3+DZaMOgmm
yxnmR/DFYDPdoNRIxd4C0sBnK7iq7nyBGbnkDeSOdxt27QyaQy1+SnacNX/t870Q
756LhlPorBvdAjn8xEQudAoTMEYlsQuV2WF5jNwkw1yLpHr/qHbJVFjRC6Z+jdWr
dsx/G4K7inV8NLA8ZUAh2L/+Ur+yY/a1YIQTUpGOA09anUP/F7GsA8jYQMXTzFip
An4cQIGWM0D5mEVglzAjuTu/aWOx6HForY4PMboR2rueEO3Ukws7Ct0K0GF8A0Vw
3jpQx0SmA1dGDMtfj19RD1tMaUnxYl/Vwk6S3TIwpVj7jYITZNK13LCMyvAHkXcI
V8XV9t41noB+8Wgi3E+pDhCnulCZgQJTyOV4BzUU5SRSUf3PaVFzX4Y8s9NZwRRl
8YJm4wNeioiI6UAl8Gx+TyiYeQHyuH3amf3hnTK5vXfOE8KV0NSlKzbxNKUoU65+
2eV64e5pXwF/KKjk6C1Y+yf3O0EQCuY0IN7gjgMwNaX2qQwMJArESv+c30Eq2CDL
XF6P6ibeP9cF1ud9x7SNxi2MkzcvZgWwwYqHvfC0HwvN2LQKK+PmpCmfuZ519Dar
PiGkggUqq3Y1p1dP6h5ody1d8aBvln1gcpU1+WfBlGy/8Tak37NCwvJA8hu3wyAh
LKBxzh6sR7mkjPFgkq2dwkc6qFN3UBUBMGYVqfXbiCD/dlgPEgUV9eH7S78o5Szz
sGR4QMfTQD7FtO3CLIQRQbBB/g/OXStPWtmr+SiTcGtC/ydSiSzD5oxdfXXQpzMu
fjix6x+HrnQ4GKfhs740QuVj0DJMjAlXwbs9kKuzCe+SP1R6BWUynbZ+7kN3+cO5
wdHJgM/l8BdV/DC9c2/tUudgQKQdWutJqLDIOb8LqxfkubXfPPwMVy3UwOn1g886
W3pqMOw/qV3atr7xm56STdW942ncMCIFRuDXGZL6tbFdzvXbRZ41W8YsGprbcFVP
gcNizvzIyORDHwb1jm1V0fT/h443sl9Wr6Jke2n3latFbOUViFegsn1ghz6LHAJ7
CRYYszZfSauTOJPpr4gcF45KAHfOkps1H86jaDzAkenQ5zTydl4pF/LRS66BpdNo
mnlwWdyhdJakP7fobNFC72cSDe9+XVDMi0jj83rxoWp6xGlMtciZfaY73tQdm6AY
/+6Wa+8Nr+ob32JApKQplHe1GH7E9epDozZWuG6Qbpy65JszUy0QdbUV4FyrlXRQ
yvR9Qf1//imZXo0t7XuYMtj4PWgjUwEW/Gf7y2z53Nx9dQLt+7GVxIVcIGPUyOa+
ts9hFgNplfhPNmMU3Wt+1tx0+W2B45zhsOfjXe+Flf6ULVJDv8MFPQJY+nCnqsDg
CJFa67xbX+jGOw5KJVGVvhbQVFHhF70/uYtFDxOH8k5om2rm3cZ6UMJgzjLtrnSy
cPkm6w93dpIatJKggDDAh2BGhsa2xeO1jHDc4kI3IOJEC0j5bBnpNnzdtS+OQxyv
PMUJxTiMdcdvEp3s2ERop20Dss6QGzw3na2rLWzWQelrFAuwhwHpT3sm+oYWE3lw
OqWGEyphEHAm4AwoRGYYb9Jy85iI34mrnnHElS0HbTA04T3vuDwyr/hqGTdlkz49
sc4zKwxx4rmergDNJS5J+37N+oiG1fIbMHLV3OTAIWY070nyyZnUtj1mKnWEFn31
AcoYOX516fyz4wPONlxwqN/zz4RVJYEEB8rmPsINwV6tRfMpXm8v60ROZfvv9UmK
Otz4kiSew2W79sxYLaN8Us+hCX18XIbaFcoKRzDbY7IHDE3gHvBSNnO9576BwIsT
D+1sOae6xOGOZeXnBx3ChFrj9FQ5WpmC/bhEKEa6iWskCldkhUWtoSOz8QvN8vPX
3TQF2cC9gse7HVgBBpvgepSAb21WcI/R5sRb0Cvxe0KGScZiRvv4G6Zm8e5grjSL
/Elc9LRvVu5lDe8FPBtnu/QDQJIHAym3G3XXW0Qpi0zwxp3KXNX7rmOYu65qHLx5
Fa38btXyyeaDccWEUtjQ+oGiFWBgzMBkeOA5gBF95RtAVYDm+ubITSWQXyFHLvQ5
jpEMP7eoV7rqZkEnXDqvwUGp+7Cgx+Q1kLhVFJJ879SgzSCcXGsDnc2usPzY4NiB
D9jJgfWOqIfWrj76O1IBhGu48DIe1bvVYKcSs22bZgmt1iP75EBSZJgo+xLrnXwK
wvqFw8DTy/XHmX5lJOwHdvxVXXYDWwKDUo/SsOKBqvvXMCAxJYGr59D+d/D+UUL9
ZXF4oP+ztX7bRlXLNA06glX75wIwolTZ71QWqDwxO3FJClXrKZJzY2sLFvFUBA8l
wpBx7g34USu3uekBW+jRDS8tHD5qxdW2H2wJfoW5CEWpRyQoklrU1uF2xmC/OUKT
40vtxzPlppP9Fxc+trEi003UYqWHTPutIMg1jz6O1Eyp2xTXBnhB0L0+zRbImiMS
S+OzXeH3RQkKEbnVzgdJnken5ldobqDX1x3F0sq7YyDN+h1Z1DYGNBOzvjJEu2R9
Jas2+N6avYqgVUUr+RT4xAOHd8b8SjpLvNkgg+YkV8Cjr8H0qETmjgx+cOh5FC5N
PehNkwO3n4bw8Xo6Eg5eLsbjK1GmXciJTrOx6A+3/PLs8CnPbMM/bpYhRzhPc9vd
bUy5GriRd3WIApxmuZ6kueqfnpaz8cJjDyhIcOa7zPBddO2hJ6sQh/N/wTsP+lmz
cXQgmD+51PyQDHcLmIHO0a1FqMQS+Z1s/W8fSBF6LED0++aTWu6jGZeO/YfgfPiQ
iqGD+R8uQHQ36lRBIDPhLfg1ltjwsiE9sy0XedCuS/dIq+0BdaQofdqMz5l9BnJr
k4ij7BnhQ5LyIVg8U9641OzT1WUWQcOuYZL9xtF2sPEAoyuPuwgNcRDIZ3iauSzI
IBF02jxwMftWoR+5VDlz6xehKIYiooLP3itE9y0RJ7Zm+HFh1NShgyYeDjVbf23I
PJkSId/48erjYCaunnA8jSD/a+2Z89ldLBLVvLjRcKFyZNC4pqTct5o4T+Zizh9J
6MQdufIzvkZ9ES6hbLGzt4g+3AzY/Q2mvigk6px2wqWHfkA6/5U4gj18dT8gHpPU
IPRU9i7WxQPipfm9MHaRVJkgQDYf9c6gmQloIqN5vPNI1YYxzrQeN6RXHj63Q1Ek
GKRb5oLcyu9jcJZnd1oemHed0wtcUYZWNK7BuNsgDSl+aTCpY51FN3cNnDcCBOi1
KvsuUNV+ylCfNkpWuN3ot6/BDoKnkKEyveI49qN77qccf9m2P0nN/Mz/LGuVVYd5
wRGnr+IQTi6i21fJDlD/N9wOuoIsrGsktsW83SPx5KV9CVofrK3mvihq0Xly6phJ
r6t1NYK575QxYp1ewGRRXZ8CyRBrFmJUT5xDOo6PP5N/LpSZPYUdX77PKdWFLJuo
1oD50Qlygs/WnFspkW37H1MohzSRXWAvpeu+MTLECgnAQLu/KvBkgMb7kQ8uhtK8
YOyo6OMXBwHWhcjCdGB2yzkP+b8q6XdlEUvAzBvzsS0YXa+0ouNADvKR9R8JcD/J
D1RU338suNlrmVGtdqcPjBnjUKx28Ipyn2P9ibsNSpZeJKckTCqqZE0MjXxayMmP
Z3zdQSNkPiyiQixANuJKyUcdPCJdFzuly3e8VDgvulDxwsK1V4A7kwnp7hkqwMdZ
xHr44XblpY8ZVARcsmEweXW7T8MANW2J8/rDMFqGmkBZ7vSG750bk/JC0DOx0u6D
CYNg30nMgy1hk6VnXZ+3d+dWg1QraAQ4r8fxxaWXiO/7//jr7nC3cXMlHvrafcmV
orvXvD3kGnMixfzaBYmD9mh8bUK4ldSmRyo1FNjAMvmO5R3blQJv9b3tZYdc7k0M
oH7BxtammS3JfTibMTXTQLe7s2GHNMWmDvB/R2wnwoIyJGAaT3GXZXd17EsFHzPt
oZ4mJmm8FAVJ4UQ0G2EksogiJ9qj9YWcvAJC68+PCVi+RunkFxRH+xijbboDKCzy
LzsG0/+qgk//TyiN7XAr0SdBVdywNafmhHAmwEQ9HWEQhLXWutD0E1XpVIVE1Gpy
ArE9aCZY3Qpf5gtx5kDqeMkiXN1BG5c2b0U5BDe/rGcT30e0ZWIgKRiP1rXJ8ZqD
6NQQvRmTvBLwV1qj0TYXOvWzWYJBL1ATnYiKVKAnI7vVbikFifjpXhm2Z36lHyjJ
MOkFZFSgVkK1TR7rTV5M6g0+gVG6RQEMyJ37gNOhGrQlPZkmGdawymBjZ5IoFoYx
U62ILgH6IMQtquHmOjwlnpP2prnr0yVTl5qf9QVKxUkGCOYoxzaZdiGuJdenrBvC
e+zIsiuSRZSMD29Vo5OLiazWO3E/ko3r/ck0/eKBdYopX0o2VISh1DOIFmpWuUIp
cA1JrB1pMF73P20SBRnu2qtAdK7k7KPb5wAKh8knHBu8IuZ+3ToLsaqXhYAbasfN
ZE5qgN7OWfEn6odJSnKuvSe7oNeMYZXijQZC4l5c80wvMiCctQJ/E3TKEPsNp32f
yQSqel0D/347holZEaUELO7K3rlRzviY0kLjUkuu1b5Hu+h3kuJPcQF9ZgeIVX6e
H40O1WojWKXYbaOinlThUcKA99CDB84FgsnLsYJgjnLa+FEYrN6f9hfiBJ7+v5SI
I7KE11GWyfcQX14CVf66jXjMfl6pt17ctOJtTEMSZ9XJfK6sE7TxBAbFeFxNWJFw
MZCYK/DGLEe4B/RhNqcbZa0LpSzh5hvGsf8R7CKQJ+y4oZ4PVJBwtYWu8xDQA/6S
xCf5UkdNk+adeIFXA3S/EN4EFEzatm+vIkgsPJUf1gCFhc/hn70qbjpT0LpU0pYi
zFA+ivFeJM+CtoeyfHdWS+JzIN7XuxqShcCOPEVqzadJtZV3dhT6yEjrMZ2lM++m
ZkQIhvJBydb+RvJ4Mufx1OX2v+e2fgqoOERaa1ZCP39hP/ZOKapbELFdgt46OWte
xCwDCx6KcQmiLOruMqd2IGdxYvNfykllDqvfmQfD1ysmvAGSt3Rf8/eJnAHvaBvU
XUJreCZ6dI/1amxpYIXhxfaS04xMTNSMzD+7vyM0ZrzXOz5Qeh4y7y8USd94fKSe
FNkJLQtYVqfdYbMw61emMMtOHioB9Egw3uRRwOhOXIXTmOt5wM/7pil6XpHNWzHh
1NtRsNbkkk3d+WFIB60776yYyfMhXaqVoSy/XQxT3v2z/a/+wWXX6eRgC61uFdEA
/BBG3hoiLCl1GIlRKtVTdKojz0mdw4DpmClvm4woqmD5lO8rfX/BbEBx/vCuLv9G
dDAiwrGR8T3C3Z1d9IWbPYYGtlfGj5CO0P17jw1xIr+1WDRHXPVD29+aIaq4+Ypf
/2j535ep1JjFlF9WZm5+hwdGcyZ5IYVF+TjVbcdwG0gC0bjvvXA+703UBL9xQbwP
puAdCxt50laa9OJxYmQOSkUCqy+/K4pcsCElwBihxYEY8WN32B/Zho2KmrtMhjMQ
aeiJUQT1oTYgQA5d8ioeB3v4qOUA/BhgvOjBbfxcMA06I/e3uak4CXPMsbh3Ao+D
NHHL/95IiXFeG6M7WbLq4Otu4uTSIWuzorvzMNO0te/JKOPZvv/ItdMQa/4q+fEP
JJvDWejK42gdXQSAiiaFNaR0MzPVTUioI5lS0OxSn1w8clgvZV/XLzwkDj9P6QI2
gws8rBhPwALRdDxKODDY89PpGd5vS5QFb7k55SzpE4qNluBXH393vfkGZqV+71nC
Bn8ChtdPQ2QNp5D1foU7Kg60fEnBa0Sgl+jqIxqKepdX8YGnVOqD6uP2V9B3r4s7
OEbu1uIEjbOjN31iOjMc/51doBWb2MWZk4/6u5sDU8wjgBibChzOW0iD7ZTx8+Fp
G6b8F1mCXeF7C0CpNA6Gx3x8il/ZCJimYY98SB2XhjVhNV/rH/3qeXPpRvVqMq4Y
FzuZBJ2E2gp+Hs20DaRG0ZWCikbbv5oTw8DGUxAO8rzJ51bznbAF5YfSqju3fxA8
OEd8vaaytfO1OuCVGI6pkQ+350vctzVvUJYjPPVZgokuiGxGGVip2OC0X/ia3uSL
woWPJO40yH/yZR1zwo52iy4uxQNMxEEV1HoNo5Kzjv9a65p0PHbB7Ge34luX+eOJ
ZoKsWKc7HJBJl8pbEtByU+cHW2XitM1sJyyefd1tpvn+zy53Vt1OIvCIy6riCRYd
j7/Yff1/5OkQ+IEW8syhnbWteU0qA2SYcinW7J+KyX5Uyld9NJsKmxZNi3Cnp7KH
mODXt1IneM9mxsdgb++6eutHgt7wUEG4x7XZVMIkGRMIG8ZtbCgVc47sQEhYYkwI
0oJR0oPEbM5SQinRzWwvfOvWhEp3MVl+mAuvS89eWmKpcuwSvISoSCFncduZixFg
rFZzJ9PSnQToTLigoIQwDH8UmK+OETZ1RUAwKlpjoyW9B/e51b9DhMFLMPq+Tk25
bpTrQDFOWpyuDs1EBOybfjlmVAteDiORQ8o25FznUiQvS4I4+uaZmcGpkbV8GHcM
bGa5mW69VJB+A/DMcCqqqPc8a/HmU105xHFg4hd5pmKu5oDdAQKrbhnMy3W1dGHJ
bzJ1R5wHpyJeP9Q/6ToSqDBCDJUge0HTeEKeGBTOA8A28/ToxUGj1lSy6yjXgb0w
lrU/zb1kS88V/aARfWj0yGecmtK04sf6bM+x4eI6CD6KRc+dlRT77Ky2ZKMjg6Md
S5zLmA+5Gzw4dTT009vNOzssnRTq5m6VbCzki5bc0G/DdZR9RU96+Z2jowyv4uCW
B1ircVYs5Raim9DfA95/Jsm9NWzma73nHOkD0yStZ6wcYwVMb0+BcJ3qbXAvJAMh
cJNjzaTPwIk/7XKDawUF2Dj/SAoOfj7bX16JLrRuo3nFZZp2UvYo8YoIA4LOyr7I
IXlvB7MjCA2gg8nTJiJHsWtyyGKwjacg9Rk4VVBRljLHBSlm11y82phXPLw3KiwU
cP+inGqULqIMkjMf+e0oPkoHrTm+AcshoHMrElnsomRieO9hmD7KYvKQtinfc0Iv
gd4jRolBePQ5nrrqDp5A80b9HV1DST4DioOgD9RHxX0N6OzcWdXs7ISIvJXnSaZI
TLOu5VzHoZJA7JeFK31IN1DCE1bBQGvAdMUuere9tUp4AjQb5MNlYvqMP2YQcVx2
UBdELlXTcG9G9+20Finaq/QSLM86Qjzkaay/sw3T/lfSikg2thcoIboAJPizcHNz
ryQ2K5gPZlpuGO/n4v+bJVe9S+fXwtU3QiQHUaiLvSr5ZYzilxrGCzH3rnxt2K26
0I0P6pRw6r9dJy9tfay+zijvo3HDhssS+fznqnFctK72aedWk8/kemmRffmTJhbN
a1fEIo8WtGHI0u/d8kef1WW+Qjw+BDwln85OMASiS2AFUm+gn8GYLMiux9gGQ8as
GZ5bNxqjZOWsn+5uC2FJsX9ik5iC/t8j0cX5KaaHzfndSgQADBktAd+cg8KgJAaI
UuzDdmEbfaTlKe2vL1gmfeBREZKLy0qTRyEsJdVfni2HdDEhvcIycCQesx2FgZyg
qawPjcuJmqYURe658x4D71XTkavZj552PKqRJG+TERrM3rFZy86kZXv8qiRwJPev
8gr0MN50zoqgaCxI7igwVNA/iau0KJrQ6EfoTNcpk46NH3fbhqz/zzVz3tr8twxK
aZlxuX6qFfZ7kBQYNahZrA0qgNJdAZ2j7iYlmMRLcO5NoyojC0NLAJckeqTmJa9T
wRzyqnLWBXpqDZy/z4wQjfexpfGfGh24UNNWZRebbtFLdsxTZWByxF/29MzrVC4M
4cALdAyvz1icvzVvdmJ+YUHu4ueYMrdqqIJ4sZ5SRdfDkQAuU7sl7Wk3GPjjps39
K+GH8RBRr32Ac6ycRpajKltLYO6iG/SWFMfYu+T1Cloh2UQeU931zk14l++IndvG
0mpxCynfqXygkk8hcebxpQgjGQaL1jWZZtmIPpnxu/MtLmrR5SOUGBjEQI2ODID2
XQhl82L8rRArV1eMU/tyAfQLvncmkM1eBpNN7eYf+tS9Bbu3/uRp/NaDtBGmxKZm
QnjGp0cJKybfWM84YKj+9nAuTvqQnIhzgwERgOUAqsWUgTLxAPsU7wDqin/hxnXL
QEKLNBmA5tk81plWaSqj5CpI+CFkGcMq2GiK2TQZhWQN+EVZDzZHvYUdpaernUXm
zeISlaGp9LphFUkvmrsAX2/RNteqAutIbkSm3UGl7MKGKsFekvJSrKPABbc6eUc0
UnG5uSTu678oVeKGC+DPFHx2ImWcx/2x9xhwnUiKOZ3BrwfGnNAr1kZJXsnmq7jg
NGyKDCmixDKby0Ko9EOpOBeOQHeOVMzZyOlt6VPwF+wz8OKWkSprp2P1lV9jIA0L
jtsr87O7dakNPYZOOecf4ZQKp3ix3TJfpC3ZUkUeqDGdNOnJAwz5N+PVQyVoBUZh
lgDC10dsOoHaKQ+GK6n+xT3b4BzA2ifVgXnnOV7ajxar6AUeN8hYRfL1nw+x+39A
i0YX2DNMlkekaZsrjWRbQT2Y0BEpPju1I8mxRM7tCzUe+z2Y7TaniP8nGWNbbl3q
iUbOUZvNbasafPhd8vvaHihsWU2FKTIZDADm8qdVlwRr1/843sRd6Y3WG0GC0IBM
RZXjo9vlUdhpVWc/7fsdUZDoA6gh7g8L4CkpIiJ9X8iADQlBUXNSAoBok4vY6E9z
tA+nJ9xVD+/kfPot9FHLkPdxZLAemHXA2LHy2S6uo7uTeYf5tSDZm0LGdQQ32RsT
XrQqxcWAogSBMk5yjVirMTVWbkXLAUm6zj5h5xn8llFYMOcOxL/TMgymIQPTM0pX
JdO7LhPXQR0zodAJHpclNvM6jqGFajbfy0yqEEmo96u1XbexfS5OuzBNcYnMPfKF
QG8qU+7YVbwHhQhsE/9bVeAEdrTCnS3iXpOp+mIvMHDTb+wGxGdxWk5n5Q7Zh2aZ
j4YCrepedmCs5HMMvGScLfY5LL9lgmOBaushh8Vb5f5iWoFrD3HcBXwgfn/6T6WM
dg700yqsR3KeMfIhyMOIL/y9fDTQlzqhVB/SsBZUaa9lSW0QQ902q4CfVH0D/pGY
/jjZIn6mafs5LOHuC3wnyvvvbxPvQDCdlhSkuveeY+8=
`protect END_PROTECTED
