`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAVsAamanEUjb7AXzpGvcnSQ2KgMtZ6fWKjIWvEvdpKr
QQou1ZLUs3V8dZUyih3uj6Bfk5CueZFmoVeWV0Zc7TAAz4gV8UMEMbCPJaMocFTk
G0XMRiNt0re6HyezaYG54gIz7/fZmDIp1r/SD0xn+7nBjvdTwekUNhgPPzxpXJCQ
uTqFYDuKtRNQOThA+OtUC04LPZh43u+5l6o+/9W5H5GHAshzIF5dUDBIY/7myVYZ
6hYe7pFHI/h3ptf9C+04DG2HyxCmZ7jKF0TbedYxZhoiNPaTBpOAowZYcWAGCvTj
1xUemo1xQ4ydEYbOPxPmOLU3Gwj4Uq7bbO80wZXNwH6KQ19J02I0JkjhpguHSnpp
HTZjEpGDJgLB3X7f8UDBOi+XwwzbRCOrvBkgBWSKUC/zty7K1oDPSLvVL619bj+k
Nz2JyEDduWqjAZgBW3U2NXuvCJQvITWp/w9u+GOi11DaP4CJf9a+AOzBoEM+uBMV
fYmqymWWS9ctlEVVeU5df13fIoFv4uE7sT7E9MhkLT7+iwJoPgt4AXTnw71KSAQY
QJ9lxt5Z53h/St+6epGE9nFMF1lY2/GNIXIra8O71o4XL/nLxr2wnxfimnzHoBRW
`protect END_PROTECTED
