`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJvmwD6kERvnV/wIGNH9rJFnnlBM0Af3/f0mXzKKYYsV
9gA/dPyiLC2Ir08ZpnVH8k17YLKAT91yRVwFeKSg1Vbg0VO/GLFHFnnTW1JWYVJ/
RxZWLlrXNPr52b2YYiYZNfg5O6vAQbGz4OlSRBpNyA0Hm0zgKIXnse6uiAt9Znkl
sMSwwHsEkwfJeufA6kf78VzVghHY+pKQAyIsChFOZwfMA/WwlZot7P0kxlc1yvm/
N5Q8LM3HxNqr9R5lZfVMnEgSKFdRb1m7JRpAvQ2mGVn6Pk+5ZdZTPJ8/8Yn0a1Pc
TtZy718Pif4cszbeLO5jY9v2mNwu8YSKRKASH7r9CpLrD4iJyYOe5HSMNRZxjqgh
kSZJeVQxHsY2s2vqnCbjFbfMWPsipVjuuIVniyHqStZiaRozOA5jfyjbTDerQPKn
MQHeXATfoGWDz3bjt5XoqQ==
`protect END_PROTECTED
