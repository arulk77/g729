`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
rJ2uhDo0HKhNfUi2z7yXQBUfeBqr65MW7SVTo/WQLwGEUW6KjJdGOUK3Qjh/zRJv
MHL/iwrMHc/AERrVqffZKWJps+FUqf7AgdotzQjbzs60NVTYP4FcnIhF369UyKW0
5mNFgFqseuq7gxWkNafAgla8B1ELdLnp/vKaUYEdKlKZvhYLn5Dt9X91P1CoN4H7
BDTVYZGcbsz2MUtFlLHcBpBZ7q+qwNIw3CeHRdSI7mub+AZukpJYFpaiOw0RfenF
4S1UqtjWD/j5XVsQk35fPBqTS/TGS8Xs1vhGWEHDdGRfDOty/0wjBcHazYhK/Hus
AvsSqbQ+CA9rL6HyIns1rqKJ2vG5GW1P1nLIgHlBDpWwKm4bCBrLYA1iwiAG7VbT
l1I/pCgc5o3U+0tafvhQN+w3OMzUAcN3v7PfuK6aY7g=
`protect END_PROTECTED
