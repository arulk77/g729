`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C7TTHlLHswIYDan5Ph1XyBd+w4WC/Fz8xKiXgPojFR8b
PiwQz+4gUctuDGM2fj1sFyvai2XEXu21hYJPXijTiTaMr82nfMT4ydoDCVd7HXSw
+VUT4zY+N2QkDzfBYGM+pgTNEYRBDMjjg7anZspadRBq7XtXhrodwBpPPM6xyeJa
60JpIcrFrf+111E8v8dINiBQGp/Nz38NNS8dTP2TSnJ9CCYTfb0TY+VOps+6zoCj
QLityEL7U6FywKE04LhMrw==
`protect END_PROTECTED
