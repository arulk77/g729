`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1abD76e4NseFV+KvW9QS65kmRJ1U2EoPILYML9jMpcwDC
OWuYdCGCYO0mvzGixkxdmxm+MIlHjXAYoc0w2LZns1ff3GwOs7WYc596jgzsYBYv
NHJj4TOiNUgsl9tyyDj+Go7GshH4LLgR4sshkVsXCMqY9/z++N2fzck52BbsN6oj
AsrvddvcU8dGnhIS2ATuJlWd2ZangnqUIgJaHwhSj6O/NusS735TWjOeXn0+zA5Y
sdGvOftegiG5p++g1gaq3T+JxytitwnYRJVOraUqeDc2uPoYHvCYKalhQEoVYZRT
9W8tM69XbWKlRnPXpT4nPiOfbX/IJ/lH+tu/NZTTT7iJpJLpdiH89N4zSqZEO3eV
ACXOhw1nwZCIGBgmaQG2JS+mchAj9ALLVDEvDGuu23EH8aITNhdoVf2LsLJa1Mg/
UpshE+HyEqE8eMj4NFIBmsvQXpcscT22F4ACwjh6Gys=
`protect END_PROTECTED
