`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SeKIdscyBvBb+cOch1RaVYoe6Ix/+Y9D+Z7O0NFfAwR7
5MnNIZC4Kv5t3y3MhyF9YnPGc3m3vIrZKKu3ARCE7FqwTAfIgdOT8xfMx8Fnmdrd
yDA+At35yMQYcuJqBdqknDWax5QnUHoktWvmd6PdzALR4gMP0/lqEC2kJ6jNoIEc
joXv5pmV5o5AQ86NOvwS7Jug/mQrw+zIlsNWDooxiZ6PhMqx0EsWCmOH2EzPHFao
Qf+widYFq2NUfD6u9wSVTfomkI1Dk2KumLo1TNDbQJ+KbUCfErHjdXDoR320QeZC
/ddK8FZx6EAIA2knzxg1WQdVV4QEIkuvXOyqz1QxhWmFOz5yCEeH9mejZwXbedK6
4/sru4OTzcrFbyDaGGvgy+/LB0IBTPpI92q8SiHCjA4oZ+6p4agpfVxOcZ15T3K5
eWHrGUcp7nmR0LQOlftykUEW7EayefcqpdnYESOlSeHDmtl/h3iotgXIdJJl/fv7
um7nuGjvObF45l0kojRSDFZZDkDxmO/bG4VwTEbCrh+J6qH+YoDKPMm1qOgVUWY3
iJRT3saRpNto00IPZTCPTGzdq/sP4LWb1nUKxmaBygJT4wEpLlxuFO4wBCE3Q32+
sAfppiHupSTDZTuw64d/Jop7vq6jTE5VTaKhId4eiP7OQoHxVsUR4gtoesiKg7wV
5O2cJpsISug00hjnRqQdTf8yixoEjo0OSf1iqd9l2NFH3CwndpIZWgIp6do76DlP
O21dkKDy4xT/wtvu2MPZd0xjY7UhtGIVvM+u5bbn1ZfLyuKmaLMpfyOHAPFtrgfG
TBdv9NFiuVGzkdwIDWaW88gMiMiMEj+6wBuSJeSgLBw7G5LM19/xl0CVuhSS6uDX
NDCoyW9e/2uKVei5c4tfFDZM8bH/ptKQMsTqeSHq5JEEQSbibBZhMiB+VcngF51E
cf2YUSQxTadkMbbWz7+IiTdhESqKYAaN3HgV+TlO1a8xgqCOS8xhTDHCRySYdcAr
pQXNeIDns71aJ/Ad1MPkzYv/VYUX46liD7zTgOcebL1PJvYokOC/KvMVWKwO6jnr
sF+Mqyzn5P47q1BXgkaBOQml2j3LhxhiD9xTUcNNwlNyS2uzMKOWGAuLBBI8F4L3
eR6Q/O9S+mPKGnq+jm5hChaGKVqTa9vbkqDGWVi5+SQgtjjj+jZyLiZ5p5k4yDcH
9hQEtvqggXCYN/9zmVD9TUlEhDGnLllM9C0kKOEy+omVLwZGpghQzcR6oL7+nGDF
czGD3TP2xsln0+8QgDFhdontVIGejRLXTSYHy54aXVX2TD9CIWhuwCi6X96kgH5s
locySDz4eq3YRD5+JXbMOvVQry5R1HllEGDTfrM/GhjhiHL29dG0QDAP3Q50FKw/
ySQNYNAw2ZiW738Rm0EQuja9asE5yEFDhXQ72AGv29cqALbOGMTGIgXolfYWtTFh
vGuyXPgVRSTjsMz5myhpAkRkQTYLUXVWSyyNz5vbWFjfHyz2Z+4vNBVMI1UkRnAM
CjVeLHWzBe0XP+y9MjLs9XGdPbwySn0qLOlSlzXoF8rQSwMcI1sRgvzxltY4ZuqR
yBnS2cnWJB4r6umy5w9X0aK2fcKapKmEUKzB2MP2yxmaD4MFcnh5Kkf5iYuz2LMS
09K1ExuJrXCGfLzDMyMxemguKLKwkjAudWo76fv+a7FVxkbSNGFgGAkoE8bqma3T
XPh1nS/nQ39DaXVuYkR6bNZIxI2EYACqaoqly7C7/6BnBDhIt3p2itCykEGee7Lw
XLRCI3TlkwOPNJj+zlnHBREFn4/gES5NsqfP5CMakJjps2Ve2/7MNwbk5uKhbM3w
H7KJjvawd3s9tfwqKhoc1Q8aMCNgYb/gCWjO7URJxSMhycG09lMjK5SE1JJTknBx
vdDt5g8WlhsB18T0jIS2MJc3VfROQLA9mlH6M2I6dbo=
`protect END_PROTECTED
