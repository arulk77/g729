`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44guqqI4DK02QTSsNwLmveFkab3F0/uUdks1X/U8xnVh
iTYVMcfYP6xJBSe41tqcn9V68jC1aHafl9fKzr7HwCogvlv2yuhUhYawulzW63WT
LAAA1X8o/OnrWHT+vty7KcRLJ+U8BKTG6402KNbMa9s+PofnJllCEzMJsHhf/TKv
rdDVXmPKFqWV3VWxcU7eTt+yVkbsnB3rI6DKaGb+lUE5wM+WXCjSrWYqanQofpVB
edtf+Zui6koEDg+6ddI60T6700wD/ee4FgUH76LuibCuFSUB+BioiZovD2FAiToo
99a5Us358VOTkqLbnxOMaA0RkRnr7RfFWDmpCVRJCm74nBt9EAWVciZ1yCjmsOz2
DgpRguElf0CZC2hYtr8Mp+2hLt4SQdNMpnmv1LnjfCHLN7qnh6vjGotRHr1xO99U
xuNfWSDlj/SBKmAWOl9gQ6wurTInJvYDf6AhdV9bMwqO8WLVntJoGtllqGPtpgdE
zj6DGV8N/4TBtFE5DiFX43Zbs4t/+ZDnJv3BtguHIAjxhWU9xusiGz6G22v9mzk4
pVe5XOdj+cPJJSq/AUDz7HcFFg3DFdCNYyKZUsSPVlzW0B1jwTDELl5r1XgTw6Ml
`protect END_PROTECTED
