`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QNw40IqJrFvY2E8HYWz+j3MJewolNyNQqVyin0JuZqGRQ3uNJUpbd5ua+snlpV5/
YzUjDWayVBQjYmEBStg9qqoJznQEZfzYl8dNfs9K58lkf7+Cl3yUUG5CD6BiMX06
kYd/0X3bNYf6I9uxCyZKBUTnaw3ohu5/ak90FmyzlHj/eqyj6KpGhvhez5TYvPcN
`protect END_PROTECTED
