`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2EBoZu9tBf8wFLCnm6xiM9vAnzloldyh/0cABezxEDiCVTZ7bmDWLch9cTrxwTuc
lLrgbnqMzhd+R2yBtXsdg88d9g8zwJPLTECkBHXkrcw/FOb4FcJIFDGyTh1i7qIh
mO3RHAWyfP2vu8+Dg4U0lvl1Q1bYLGEXbTAdAwN6R20rsPnn+Rk0RueYCbReLUHg
ELLqEDgh/qVPbj7BDzuOaw==
`protect END_PROTECTED
