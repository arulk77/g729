`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
OcpW7aqzNBmSyx0ifJQBYFrxJpPCXm2afhyrisqh5TJZIOvp0nE0bFVRdV3rklLV
9xZsFh/HfWF3gQLH7Xqiv+FFIs438G20f3bHQpLHFm8CaiIQ1z/HWKcr5oMsR1nB
dQwFherTowdR6tu0sxDJJFQ+h63cL1kPRLitWJBNBNBtBQRMSPmHktkovYbydb24
cDgbcejyH7GwHZVjcGuFZKPCAPu8rCcldnn5WCx+s8kqw5qd0j+ihkGKgtYRP/Bo
wSz2Pe9qIqN5MRSHTQKWntGnW4JDrOu1kL/EhBcIEzKy9HGIdsNjfrCzEU2GxrDG
E4SqJLgiqYZglZp7SjlBYW/DrD+sP55UqZW5/Rr/hn/tY71G+yIow0xlCT4+eRXm
2iGBQkAAgYwhcaCHCLYfkQdfGF04ZTfsH3GOMKvSAfQ=
`protect END_PROTECTED
