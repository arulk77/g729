`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBMAWReuD364D50EpBQJSMx6mwNFGGTEBpt5son7xb8s
uuRvr68QN6tsKtdwC/0D+7KIOxXHcJd6gE7TrwmhIUpJx3yAsK9HKvuhalsK5INX
vbgp57JRrX0ZYlX8LJXDs0CiPPez121vJM1no8NPaACaIjSDvywMS+Z7EfpDqQo6
v9qzKk2m4U/xEkMWZorh2Q==
`protect END_PROTECTED
