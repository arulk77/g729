`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Prgb+lMGK4ankHVaNnLDqzQwUH70aPheR+jaCKJJ3ycojufdGUDacmrlWSOWf2HS
TW5/BBnFwN7tOw3lz3KmYz6dgyym9EN1Yt9hVCR+dIokVfm3c02oZhaAds8Fd5HW
P3Gfek1tg+xlPXOsFJCrin43/X0oVQwK+9dNprineyQupHLBEPmJ7kIfiRZD7rsw
PvhOtJlthXRcd/tXGlmJkvekLX3/cWL5Buuq+E8ooeI1YD6zpQy69uVZr56BZoV6
lsjpz7eTX8M+m6bCHDKrvh4uG0Cj6zaj4Xu8FIlUPZO0DHlsQXg4QlIJ6RVVb7ky
VowNXq3MoRcSDAwxwWE/oQxNB/pnlcj8sxADNziIq81EBa78IFaU4eUULJhKfYpY
`protect END_PROTECTED
