`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL805ECx/QdBMKUCH99fs4+eofNGLqJ7DVKu0ru84RPlCe
zOwDTBiHLSPFfImvhAX/V0c9ugFVkHtSxAbrkRKj86xci7SvA4zNW815bnvAwSk4
CWWQPx76BuT+Zpky+trc4TlwqNUMnZTcwmz2OAU3EXPZ4/aLyr8M06WReJd0rNtV
GeqRySwSAwsYfZGz1AqFkOquDwdJUrzl++FhARcs1uTrWnFzPAhgjcdpM25Wo9KI
RRTgHr2yD2kpmjMLexveopOLXFVqBjYKKkrm6+WqmAz8cnDCQX3A+wkiSnFytouA
NutmnVhP2LoZNUV3lmcyJ4mZN8FvCuO+364m+LQMP2+iRJlxjHSggzEEVagL1LHh
O/Np1p0WoxvPT54rHlDsQWWFiM2c8DpS6PEBKE+sxbUDEi7HE6BB0SCvqXLWJD1t
GP0SIE6xWECUDF1uEQ6S51egzyyEhq6YcBwhIRpSHew7qZ2E+KBoGNeuRakMRDjY
4CNOr+Mmgr0gqzzr6GPrQJf7c7mifV5H7zG8a6VXTT+zuLUvXSbTQErEygb0bbTS
lSea+As2I2sIEcQZW4ptzjhWKOlj6H3RA1dQdmDxaN1Pw8XDAs7hKvsQe0/uBQ2Z
u5bFDADJWei4oTEyUCMyLmb0wUi4H/8SevhuoFQRSQymLadW4UlCEKfHfi5gIGkj
n0zeo7q06CDo3wIv39iOyhVpSd6Lwv9jrZ2M3DCwrvu1Vs3qSdJzoOjvOxEIAIxB
qm+5fOiIHiQY+B6qeXrHyktVWebf/k3y0HVwz+jwhL0WnJdQCvsZZVgozpjPD2+H
dRNl/T/LEn/CnjTMu6QuSnJsschflb1IzI97AoD74b6WmvczOHcv5vdgR/25paw+
zRl4XocXUoJVI8SS6G1i/LeTsuHZHVB/azPoZ95qx3MkZpy1Dq+S7wsxfLhG0y2g
YBAHJl648m10VDzG/pTt3dDYegxvo2fO9f6qvuNRWrEVs3XWw28i5Nng8RszQBEG
2UtjZNFq7khVtw9DpLpUZyHTVjvoSLYcKPpFxWXqZbDo7mo44v3AzlfkoLP8meMw
VNrG2TzCUi6XBNmncG5p0lcavBADxoYxUyOH0N98/5FOZEWuT0YcDXHQU6kJvHN9
fuEKTkNReRrZnXZ6cO9X4CZ2U0awvleIsvMnQtY9mey6pIvcniHI5EvmlVNiTMc1
EXnBQ73mX+/yczd+nWbeccCQrY75WVQwpeA9Ovy/tOGWqeJVor4FsDzPx3GnTwp0
9cOm8qe/A3WFY8DI67iU58OoyDZLfylZEU0tVsSSzInGklRVV2/kc9M6iAWDaijt
Fb6xjAL/VM2fn3gi+g+b5Q97iNscvcwxI6E+tljUPGWjvKu1rPy0/QDGKPIkQlPN
Edy8FK9rpFCX8thH8mcXRDn66Bow3OGcYD4b8PUhjTSdyfBUcHr4LEDbWstsYl/l
5pvqEh8tUNo8MvT1zZFegb7bTJOXOV+UfoP0xJ1KgQtNeE4vCAnQfkluOX8uND4L
hPy8W0YsPMpEdEZEOy5D1WbiHnu4TWxkGkZVlMWabC9FfE7mdMeLjSiKPBuNnpmF
Y4UVqqPKBEMqDAhi6H70Xx7lHUaUxHDCUCebei84gNqEGO81RHf53OWigp8Y8Rzy
lSuoohe3wbRWB5Qag0JfsAtq+tP0m+jNsLjxlyV66neWUA99ByUlDq0jU6CkT/Vj
fHevJtgthKX/OtXiUXOFrpvYjgoPZ4u3FPjy0y5v3ZdDJHS7pPEFqGtNn3fJ+Zvk
lmDE64XaviFbkCednoffCdaxNF1x6xRyykRYuxT+SWmUFtzV5sEnZif/GsWLd+rR
GOQUiagDx9g+aS8FsZBa7ITKHtfGUj8zeiFc4RNtOMbzcFDgouFsnwGj2O9Ci0Jg
iVPj8bbdJ1imfPJPTxFdWiXgP7R8YTsh8foJ/tAyf1K7tX+G1J2wAJohJTvmcPQl
reUVAd1CpeA5KMwb84hTxhvvY9+RmfcPAvYMJJSxhl4FdwwrJwmQhTqz1b+N9QVA
0/nip/ZczkY/cW1+AmjKDqFcgTJBnJQ0Fh5XtPGabugWWFTPkqfidlGlSDDjxQs0
tNsJWjHIsMVsV+APZgsPcL9t8plR59XzG7xcmWAJpzj4H9Bo8WG0zeEPKpVFIVTW
LOUD2yaiwz7XRMAyfM7Vd1oUJpCgG/0mfSe3eq+7sHQ2DW82YIICxahgUMA578il
Aybz+BWb0u3vsWRgXS7SBGKKw1nnKpAyqYGTmJNOehYNm354PuNAnbwKMDw3qj+w
2Z3eldXayYG5TD8y/kf7ofN6uPU6pYfo0nHq8jKHi0jY1XdAYYVdllfXFGgP9gP3
qNyOVH/rKlseFqfTnMxW3Y8iPewipn6LhhicVwsRhiKghabWLZ2Ew7PNKXZl8o81
Gj07pwSJ7w53fbzQKSbobnUojD7l3gB4zdn2ReLhzu6zXoVJqoFCt9Erj1Rzs7nf
qbN8HSVVIJqzJpnOgLXv69TmLgKUzf/CXkzuKv4cz/tlU4yj4oIJPZT068mDESmy
RMwSgtbBPZRRb2XNcErSRZSQ7dPfbAbDbrlC2mCS8AC0uq8PVIayHC8yT19UkQpg
Dj77lsSrNfjn9zPsmZjNuuWENGFF5HVyz/r2x9xpi3mSbNo08XEiIbOp7OOj1sUU
acNLuSL4fLtZo9NK1pYxARxISaTEtmmEoUBI1xZLF1u8OkI6TOql19evhZdEqBDP
QQb3sbHzECQw923IK9esObyYyowojbjZIXoika82fw0gpwaurMZ6f3UzQs0dMJH9
6Pp1rwwit+o4EpRYmTIiI1G7h0U2vMGw/HZX4emuNVtQoKOBkd0+PbrKgM4GXZ0q
8XdBu3YWXfNi4Q99Tz5DTRhefCWEJYsU7PGXa8RqbagX3hpqN0kpWpAqdBd4qRqi
TGCiGo+0spgPLGPPCc5uz7NR9OVtZ2789T5iNhlnXxULiwa3R1OFLB3ov8W53QEY
7SHWXDc7X8y242kCzZgWaBWrAvd1dDHDMdegweJNxJ4G1dRRiohk5gm9OaA8KazP
hwjUchXlGQHJTIXBHKIiIsxXfhFqQ2880/HdMbZhHBmoHgip7D5SF51jqwb+qdKs
dM3RmsHLsGV/J2/WQIGR77oM507brtm9knFsqIhuuYuiWhBFn5sf0iGO/H37mTON
Kj7meOUAr9aq2oPTVcz+BYOWyRDAKzNwkJx5kOpqaEG6EPAJ2DEIXVxumPGEWJhY
UCO+P3yfKFrhQDFGtcSGPw1Poibee4NoVaGK7oRm/4T+ZnHee2gCWM4S/dwowREv
wb3ot7Vmp3+XrgRPOaT75xf4+Pidft8o/EkjyuWYol9rp10lpXZz3bzuI+eItGoV
sdTp+HFB6Lz+FNvjf+yqkOGJB92T06wWDKO6q/RBq2zlC5xM3Wbi4DoJDY/XxRhn
kZ2xiQx9LHbKpt7vI3+l2QuPptn4PQm1uW5xUnZYdQzeMEv3aCqiDFxeRXzRPmPk
R+op+8fb97l9X+TM7sY4NHiTWGYzecUaWMI80kfajK7uix5hNbEjEduZSlWPZDiz
86XGZS2rOtWVjNWEjr2k5vaa82c08Iyn1gNis62wnrODQ7/QHCXMoZPSTrS7bsTR
MC4ifPOBhbqydLT92/hbQpOqCFHDNoxe90ySzC6IZT8OeNek31W0FBQezEtOejp7
Wgch1CEiNwmRJnyuwAUFxqGNUzN+ST0dSbYoSp22DQA0jjH0/ABZiC2q/rzJNVu4
BdTYATQU0XzADuXiVMKBZBLQqNO5nQ3vL1ifOWZ/gtrlljeZc0ris7eBWhXTVwxD
Wfd9yYUN/yX6VLmhhsD1E72fd6dKzhi8r+Ull14ldgvr0utLgOaNgOyBNTLwLVv8
4AeaK4G4G+Ob3eRVDJ7Y+5yd3xkwKLP2uB5qsfowYkjoGCKU93PoedXrVmIdd2ZM
btajFZ/dohQxgMD1Jp+vFTmq8yWVhiXgnGM9FxJh7HIST48De2xPMAB69jxa7tNP
8OJher/bGOi14POgOQZX26g5bUqz+G7XAAomuWodl++JYDIDBZAllB1lYbcRbfO9
d4qT9xw2oQp15uuKOKPX9qRJmZ7r2SS3Xs/yXEqYvNo225oA+u5Ki5qiXE5mEjL/
xR296/d+sKZtBGLExDrVp2jQeUneM2TVB4P+IsiC+EXXaUMEK0mpv0yQaE8LQ48m
el/AXrw+s+BYoKu4s2iQNpFrUweeI3aWyfqBSEM5VeXm+4W5Y7FRW0h9x6xX51RB
1lFzOq20Y3KDAu09LjekmmBFxKXsswQQMj3S5ZrUysABHMNcH5kP3qTzSwZKULbp
6R9jsE/yaW9MgSDnP/fuk98VRCsLCTYQY2lfrksIhwofOIJVZoIfyoxfef3Y03TR
gQj1HwMi9c/KCP/kPFFzdaVQ/aa4Qx13dzhECc+aSrAbirexS2+zJVwo3TOuWssg
cm++kAtOkZHtBT14uNsCbqjNFPk7HdcTl4r7eu/V8ivzLZjyqL5dwC1jSVOuFjKF
I4q5fTrtIqdO0pH8JqcAxuPj/0MBypOT9R3OXjYaQC2edPmTZKrk5CX316pmLW5D
99rlQDp4XgN8b6FcyzKkaxQsGpi/5AdB0oinufV2SitTQ63MRMtx8r10pLF33bor
1x+hHHXIqskiVi13nM3s4TvLl+uN0fqz6VGcKdxfu1qMQfrCJkeyjFc8O72WYyWy
JQDLjzlLLb+4113kPgQ5JfaZnjPn8GdZaSZM6Va/boy36sb5RM+IjwOigpSkt2p2
qWAUWo572P7AJNvIF5J7irXHFOZZYd18mCU8r/Et/dtcEJ4LDPNRgX3hw4kMslGk
SHaMX87E+2KNjZAUuHWdm94uhJT/QgKyj0gzFDawdRFk8I61EizB/TPOU5/+hfC0
qd6cgu1hYSbXQICuTNyZuSN85hmkxR5ZIzj5/AIoE5o6/n/ZGVpu/m+wvub/akuH
Na5K4gOAqTgfYrJ9QBJtMatTHhCV64vwMGjO31Tm+hLK0KnzLlZ4tXRtyFSR9DOA
IUQw0LVhvlnEj2gNLnlTW/2Ivo0c1XpbDpHr4AbsN2x2DCSPzapphWK8jrbpWMSa
qAgrqwXJJrp5KXfPOeIKWzYOUzK27fthC+MhI/vwIZ/o80SkJwSucA7mhLgoqRZ0
z+JYWr/ohWq/Q7csfBH2pdhR+RhQugIpkHclZCRh+b2lW2jI394PLPl9y4aijWpp
jCE1kgRQ+34nHmFZtKMzql1LR1LmShN5aRPpTHSabascGbj6gf2tBXSgSOtLW2vF
h6f1XZbDLtulAYpW2+22xDvqE1xn7ftapguTj6I8lHgVxxExReX/wbejzK+JFgn1
pfcruoZ4KEgyn3o/l1hw1or+sro/83U9PbG5eYQO0AF46UhJ93g9cKfDnYa0usSR
XbVj6eNqPWJpolfRRAm5mDfJg0gBb/alb5VibyV1mR1dOoA+OuW1S9emFV/lwnK9
NpDJ+nME4l2J8X1Z1iLcp7RpFjM61pYVPe6kGKJlL4RIVhXWOFFz4xcBVzHEp10d
Dx+khTtjm9YLCYNGiSotRALAuGKmAVCBJTX8yjyLyfr9ZQ3ceIpQ/OX2Kj57/Kxc
A2CkVOn+UkqL1+XDkErroR6MpBhk1vKanTqDLD35xwy76vs74iCJ8R3/xlTmf0tD
BEcUfj9S2PqtG+J6PiktAsC/62jlW+0HMTdxWbR7jfvayFyuU02/8VUtKigKucay
0wIHZ0hGje+OZVZTWInsa5i+SeKHk3DDMUWzRp3V+MAsFkg/8vhI4K5+E3xSGdy3
kWskb6eSJM7ilA+wn0E1lMp17ug7KlBysKVvI4dgBvQYwgjl4EiETtpyp6zVeeNx
4qLJfF+xZUXlXPWLmhMNWMibGD8o+k2Qe510KS8eb08Yv2rPrNiYX3dmur94WFBS
YnM2hB0hlAs9NUI1YCt39W1c7bW/ysLCJ9XOylTyHA2tgkp/oYEtj9Tob5bTU0eT
7A/Ho/GybxIetvq/XhPHi//ZTpvRdzAF9MeObZVMou/1SqoJmBnYacVtObHn5toh
kxhMKJSfb1uTxMC7OnPcjTv6cM/wdjvMCeZduVBH6l3DOEpKRnubHpG4IThB1fuI
PCw5wsN2iVEQ6s2ooHndzBOVbM4fPDZu9/684P/NpsYM5sJQEZD9gzAoj1vo7349
jjEvyg5UauW0gYb1ZW0Q3bDdYk9xdAsghBH4VPaHXgphpXqvFol5aIVFqe1TuHaj
BZLF2AAj8V/HW8wejgqQWhLreoghowrr4mnB5TM5VpLq+OZZkzHQ66B4pr1G5y17
6Mfe5CFm24ywg33O2cdh18uZq9Wl4aBdnscIqoobM/ynCJnfo0UPRqpm7ygpAp7o
Ao0XzG0jGrs9Uq92vaxRGO1UCKfP/bdiO7YijiDoiHcxYvpVitwJmBKxr0Bpz7Uw
HKw8b4S/6GUfrGQO6GcMY1cuLHKbI51LQysuV3+JyokaK4glx8eJ1ySbW3tAvAG3
2GLpcrfXNLHoH8OKrZzzxTZ+y62ZjaCuZvsS6jRcsEzQSB44HVa1qozxbHduPQ41
SBdw1ROCrYvUdAU6roZc8W7ZXl/GRykDzp9jSFMit1ARdeTBNDmTvzDKQ8t4XUEL
ye8gcDL17fCoK8rynQ4c/6iOc+4+xWm72Jw35nqJ6NCly+gHvGQncOcS9EyVymJs
JeOwZA0zNSbWkuyj1jdC/w2t0TfSjVtKuUGr93fL52UPRPs2gnfKTq1TcCRyDMU1
uerdBW8hsrfRzb5jgQ5gyOPOxo6qjUzr1HZAAm087i+JTpecqKZArv3sijjaVsX4
GLB5gj+Pf6M+4fzoJxaayLgWapSIE5/zEr5c7TYhPa5+TCga3sJx3dOx00i5mowT
SNPhmbd2aXUcy5gbdPboIYKEZIBHFOpRmwqnVtZ0Yn2TFyNIENz/Sj3NCMMVgI4v
CcniLC/JyUxOzdfTYIWHwwW29OSXA6kLkhfnEdj82FsLuia2kp9Htc194mEyfuAY
PKYleucgvKAqkFkNO7rlHKmlvb0Vpw06xUdGMcxoxrY9yKbhIQH0U+nZJPX6iIft
PFtiABwGlawRRqchDjB5G04ePcRyyvF54h/QvV6ydcDCbgIZDhJI1NrwaW7wKgxL
+yD88oKeH9nO7X3yw6tJexeIP5uBl9WpWlMg0v1U3h75mxrmkcYxsBosC8goqZEq
pCkr+SrGyJi+H4N074R+pvqVhG2Sg3fZdRa2pNO/syjr04vdxYG0UJjlMB4OxjLk
3ICZ8fjyab8MG6e2fBcqnGhnPuBgazYgU3/P1QhiW0zz556Gv8Y6NLuTQfYhto3l
bL77m0g/x1Xf9Qfj4OeWjMWGHc0gWs+h+UKbWNLV68vktU9YrnRvSUsI/LdQFOTo
nOF6Vd6e5IjW4FQqpWArSN0D47t0yOeL/yh5zXhuXJ+OxjwSSSGjb4/s0bVJmqfN
6dHZ2jHv+QRxRBGL25snCHQJWcTgLXTkAp1JyNKfJPn3CdWcp63qZJPgRH8DNTTO
gYJ8EkWEl6j1FLvssptNrY8smStN4aSsBgoDDrUUXnnVTaTeT6gz0JYjg6yPhp+c
QXNHqawtxCRZ3StvBtUrFa02Ua4cAWPHTkCDjng4TAXp+0NKGLlJ3nCh/dlrWOH5
ysMFN1E1sbAy8wRv7G+pNJgfBH6xI8e6Dlj/Iridz13xDd3MZgxjjZlS9PrE5dmn
g0qlJCOfFYHQl6pQ2DI4PFijxHIm3iHdwKgjboHmaPuyByL9gw1/lWkgqmR98/Aa
uDM2Wi+LnxjpikNYWgLRxxieBJpp1X9lAugABSXlwhp1Es2EzruijjgmkC4stlBy
oPRPmgXRNMaShpow0K+q4jjFu7HUcME9Dh11WB06y8mFb+2PzQskBrnyjMdNapxk
O+KkEOnZ9ID61zC8cxqePC/HQTJougo1GZy3sGnyrMXUxILORBs4VVSlp5vQ+CRk
JJE4GSJhX2zMwaLhodlIAihE6wYR1LHspUD95Y0nmeDunVqZxFyuNCxy9WNZteCK
flHQati8bgmtt7JB7WgBdhZE9KPgZqSIzl00EQJn45LcKwcFHMzee/VhSX04wLom
gX9q9nnu6+wEEYC5lUQ+wzfrf/oDuz7sf6HQqaZ+e4zzVoQtqrEdPJdn9XKNkBE/
H40Tn6w8rbdtluxn5Qsmy4V6n57Mfp0xv/skK7cUxQNsfuZf2rW6AQfH4e4KjLej
7FimMFop+orc/aar3cXG2nEo2vXUeFlo3mCKBZTmoDg=
`protect END_PROTECTED
