`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
8v53/UA7yagnqWuIJvyp7keEpADxHSYPlWd2+Mk4TA3zwLB83DTNsWz0gdjtq5AH
PPNKNEiW44G8rSy/lEgGRqPiq0kQOabvoXFueSRrwRSvUnZ4JEXy9jJBRczoRYw1
jl8O/h7/36iggHzrHfE07Rcsfvk5AvSkGEeW54+EYLcAARq6Yu3yD+NOAz9jcvnW
jIhumj5bOzLRqYtoJpjjihnlnM7jzIC1CygyqaXLzaADMBC1rTDzd3UI0lQpdQFV
Cg3Fq36C/YmBjzQJ1E+egU0ldU2b5gy7z4FtjXll9Xk=
`protect END_PROTECTED
