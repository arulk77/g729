`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOUrCv+e+frIydDIGdLd2xhQ3DZuwH4L+cjFzVBzR2tB
hW+lwAE8eCGx41NNQXSbdb3fmzp/qB4WBy4ZzGqH35rFVZPOiNr0F5yTT+vWVKlW
UoKHKR0dGDE+bUdcN0veIdN5L/7lie6ikQ7c7SGM8X0ehvZ6W+Cy096xeP+cH5oW
+wBDAPnTKPItdnEZ4D4iNZlF3so20WYAUOvWs/y26IMqSCTYhKs5UxHJh4zRqTLT
6PWV1gU8cLrqOMaZ+I3t5Sc8THhAByF/rnqf+q7koRKdSaUdd7c1vz+vEdu+2e1E
kJQjg8FwsOfSCtw5Vu6uPScU7V3j7GZCHiQwZl25JgchvG+0Ze4udssXMj3j5GcP
m6sLXrXGmlhzc2IE2LlgpWxJzz4SI3Xu9hErPEexWsp1jGHTGyyPLD0eRpUBdboW
dv0WV0m7SwykpS9Eo1lDLOWYsiSyPYVrc9iH0TsknCLcKN7AS88R8BWsZ8D/27U1
`protect END_PROTECTED
