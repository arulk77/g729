`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKWomLwnM+OYEVfduOJkEcprrmtQZmXsczMrokLDpVmg
MIp38lGEk8eAXD2e3rJAHjeV1bWVaFpdkIzWDpGO4Fkj8oKNbDNnJGshuNu33hRW
UiittLNRLkajQfhHPa9HUrYbTZnNj0xkJYgHBWamgl/2nBFB83uY/J4uQhm1iO1A
7HZwcR256SqMVf2oJmKR83nB3zBuTQT/JcEyPHeyMEu+j6cT18exBxVNKxsPnylt
osY/4Uc6JKMPueJZIjoZH/Ub8vC1NRxpnnvvjM+wWDtpGxhfg99kbT7CeV3fouek
vT3b9RV/rDFoBiWp8gijd3Hldinkwxz6Rn6YHGmH81GzFo3OA+zru7qnJ8L9BnJT
lc0nPKkYLeM3yb256ufyxg==
`protect END_PROTECTED
