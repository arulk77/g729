`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFxMsZKBZ4FMkgv4RPq1vCG6SMyGdCTLc6/x4f7zukoj
6nBfwInuS/SmruwysjVz8XU4rAzs/K5IS0f634R/uZ/JGr7zYybs4plMl6Wv8KoR
IEPXAr2p3RCjl4baSXvRt0wyCfHeeiHuiwHRM3FXVkCYKW+poH8iZyrJHPiaHVsX
BqukL9jgwS/SkSn+3GiZSMomh+YhENuhn8NXhLIcONjBtNDaHzd1tKq9Otw74MWb
`protect END_PROTECTED
