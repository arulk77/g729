`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SX8Ra3rE0zpchDldYqLqCIA7BuH1+j+hgDISdL2PkDvE
gHkIW/wI5yyvXL5V8ir7dbrLmpt5NSpugKYx5WC1mvDLN0JC7nj+Cl6Fip9I/wYt
Ft2dkYUJrNmCIeqXA4hi8RkBposWx5IvbSL5vQ0yhw78lZzv/i1pF4inhq054CDH
FUw/tfuhTWycMVbkUYZRbg+AoKzOv0GdW2qLjHCBo5xFnEcvrsAMFa2onTmv5gAW
WIunsiYfLQns1+Bq6DmcFFBLrOzNgL++EkkN2l/zEa6ny2ZVV/QdSrJrdqsGGcNB
V3QxQORpkdED/7xxZfQ+FFBrod3U8hzdZwY44z/RM/SkcdmV+R+aVVeuPLpUFTiC
`protect END_PROTECTED
