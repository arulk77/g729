`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+Z78/NtQ7XU+GkkWrqYCxOjsqontXrPLK75xeRfv1yO
rg3YSK8/VSjUaupxECKkZ39zvc/CQdRSWKBtkZxTxRhvrVaDq0/ruKXkQrcUggD3
9bvJzC9y+TCafHaREqzqrxPXhXTPdq/gBpG7/BkB4avJan2vloPoGe3tSOqoCP88
WEL68G+Ctk1xYnkzHLYaztdF1tMj1kek53lPeS+iC7xKJX3hVft5CHp167xjST1N
1Esv4DDZfK7OzzxBtZlmVyL/IJmo45m2jEUzjBzlbVb7e168LWAbvzjeTEQLAcx7
dRwCtv/40aLA6WLONa/w93tUhacZwK175WE900XoCUpVZzkXTkJZThELIZ1u9HvT
zrixyXjT/MG6Ey6wegRDNg==
`protect END_PROTECTED
