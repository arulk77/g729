`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
N16Ktw6phCJGhyCi1me/Z/MNC1u1Ku83Fxdknu+I2OFCslU/pTlGfFme9GwLqoHu
iddJ5vtKh29LNgNaZLQCG5sZnZZlzExebSY1v0slVGS48V5sWO6jB+IaZU2jQj5g
ZLA1nSoIMTdRwDzE8N0b0iIwwxYf8DauIx7ZqbTPzKU7naw8mGUAxmTHDaJGmQt/
wzNegoFee0R5US+AXKZri4kn6Xbgcux++gRa3tpP4YLVJJA8LAhDtjIYXwfQ9Qr9
qaZLwXaww6LAL44pof7bVwYKoIamn9E6fmoj6sDr0Py/J6Ny2IFqKRapBudBRQBr
jtNLqA/ObuVAuWGdgGXVuAVMQx1jf7nVNBqygoMiqvb29ypClpLt9N21mx/BpIR7
Y5Sp3Lc57Zb/lETWPg4rfp0lHH9L+/FLqMKOPA15xxkPRrpAZv8fpZEGAvHpnWzs
t29pr41oFpcQxrsk5qp8hJoLLYJH68sbnDnueIARTKGCfPtyXqf1fYrMUt2+Vgko
k5fkMyT+UYatxTJFX3xTc6hqyqw7n2oKEBbhq7m7N/dzk95/89jtnNg6G4Wc39HC
nxenMI5jFR1ndguU54EZ0sZSmL9qJwqT4qotoEf/tho=
`protect END_PROTECTED
