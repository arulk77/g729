`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1afFafNLynlQMpubqZYNqnblN9xrAUvk/fDzrmG1OVdXJ
Uc2awsicKAhue9KzBclHEmbnxoT33wL8aJEImvY5bWzIH8vhbQ/um6hfJfRGepA8
ZlRG5UuIoD9+4PMs0h1AfnYTVvxafh/8+WaecgeVtkC7BniD9u2muyy5EgVkNyak
Ixgy+ZCoxkv+KarxYFxOMsTr82u19aUVV6NKVBw9nWx5gVgEau3B87ErB2vG57WH
KgaognZWpvM9ZWJDz0rYSxrJeXILx8p6gjHJrAAWAJFABx7mbNNMo+eIPPVqaA85
Lfuj0vJfg3V+fhAiHZ7mIeN7mw46k9V//L9r2MxNCt6gFZzIpZ/JpdYt+Ds2+ONp
lXEYk6OHXdWGl1x96AgaBrOSw3X3M7F4tRrOucVB9LYLvqshwpQch+6mkRAnS1rf
2UHfYCqQNrZsUvCheJo/NP8zzbB+OYppBHk2zQZEAMd6zL6Ms4fkdv81tXCbDn/0
3bw9+TO1LdocArw+S8PVCJft046OkkQfzrXva4jc88THG2RHWQncQhugkNmBaUlq
6yC0NCBk1pgnzRJxKUaxaP1/Pc4F6Sgz/KE42LFGE7WxC0E6jaj1IEBbv69dOyTY
CbHmAFwA1j5Mn75BvvRMeu6hAhMVwltWeh+7If7daIRk2/xjhaxIs7ubup98HLx7
ATW2k9mq4PemPIJVle9qDynQ7m3hrSWAt8SI8qCdOVs5IMf1jFi3leVTPgTHlmmc
E6MHw3p5C6By6jNgQFBxiZZwVRXbMS1zGV2LQVML2vAtaLfjOF+aAbcor4Tclo2q
IsBstNrU7VDBh0UboG3J1wppg14QFPWqsYUrCOhacnE=
`protect END_PROTECTED
