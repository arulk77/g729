`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4jUYkdt5VjR8oFbu7ZiLknE165ZkMl0bpqFZeIqCJ1d6U7SzwyeyF5smR0jnhyB2
XWLmhefMNn3hiusEhmrej/WO3i5TMlcpEdLigl48387T6nuQNWQKZ9xpOYDxpsGn
zSFGDkRITw72EsYwm4L7msp/B3uMXr+695Tom+s1VtxB2YmGjIqTNPAVHbLHrqp0
UcGx1kcO8CBOTwiCTWYfS38IU6ADeoTi7jbxIQSj/wT9m1yov8Ami+vSi+fkqOlI
IRTZGcdr27H9lNsEyJMKG3Grdw3wJYd3E5T2qeP+fJ79wFjgI15FyhTjvVglMfwT
`protect END_PROTECTED
