`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
b13W6hvBWWwb3mHPEaWtCnmBcen04ggNsUOqio2Mls4vf7up4z1x/bpRN+yiHo42
/181x+v6kjnEJ/mirwdytzt3PyU2wEo7yA187qbN6lfoggGThP8Lpl1TCpli3kW/
7YJ0ebpAfblFm+y4JUJHxah1fNC0Ewb76lOuvDm/Jrqw8ke1sSAAsyGxrwN0kafh
hNocUdVbBMJmupww3Aw4AgaWEzZoMXEaRdsPrwh+7ZIxWXlzm7mwwxKnlz+3pEY6
JWSrZL5qyXhVnQoLNs2hcvYGVoKuMLpYSewfe4NOXXFXn28QljsBof/EhJyTtORD
yD6EKElakfISoZmsbGOHNkQlFl83W5g1oCx7PdhzjpLALYAn+WXhjQORcNB2RGQw
rLoXKtiYTwsJ4R7tErmm03FyMf+x+FximkCkwHFH+YXN32DYWOvTo2IRPmiL6WlM
fq2zfBUNQU5T46WV041yMyy/0i4MALAP7M65OT9L7jNTPGr/OCI3umqtdIJ9fryg
3uh0Vro0ThltasM5/w3nHMn3gn+386YVQM7D01404X2MOn/jGP/9a5D9MXNDF6qz
l+eyMXptT30Qo5JZFkOhexcCHiP3TDTbg/yoyZqSP0VAUZPwM/S3v7RZo1gaiDhV
KS9wlctSn3EL1zdcHksQZXFwSx7jZvCRofDWcF5EP/X8VG4Zn6oq7QrIYt0kaMaz
qdT56vwqxtzTv7xBURqF1143UQEDfNACn+nqAseXvc6yckqCn8FUb30ftqMAoeV5
5Y4L4rZYHMSvMCKQMjxpdvhrehofgotzTu+VRY1Cb7P9Qs8R0eEX+W/5U5V9p5r7
rlGdZKoyqzeB2WG2GLNHrxlq7pGfEbkVqOgVPXljWx4KTWvy6O2Qhq1cCyplVJPn
y99lq1rlajLB/ACTZmQF5v0QSxRwY9/irT3h6B2FzPFbsWcqhzrumMpd8AT1jCqs
dbPUyca7lM6eYiz68UFzfsquur/eGbWzV1hA3F6qduBVX5pYveBCbFGw+oXzrYCR
oYto6uTbK0abjYjNtvxcxAzsWvD37DpWk03WCLqAhzg=
`protect END_PROTECTED
