`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOx/otv46fOIHvKragnn3tmmOwHB8OE+4Qii5WA+l9Ha
iY7vL7tmufcSVjGXfP8cmNcTbjTptoEk8EUzQbu8350514K+gfl83hbffM1pr42C
DMqjwVBkWUm2TY+C9wVEvVf4nvO2TOJ+dDPDv/XTVIbSJNKQ9ox+TxqAlibG9GbR
IoDdBQRrR3+OpO9u8ohcgWYo8voic6jOrl0t7xIpLt6v63RvYpU9DQ9cmpcDkRgN
sSgZe+AX4iniww/XDWMS4MaOBPRzTDOVFzydgu0XUfgLJEpZaeGW1/X6uU7enPzq
Oqd2wSmepzlqLwquUMtg/Q==
`protect END_PROTECTED
