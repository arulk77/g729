`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLv6iZ4a2kmkrAzMzaEypxEwoEiXxNMo7/8Q2uEoeKpP
zUDf5IYXJ9KWycqCv8M6N/B4OLkC3WzT7Y5HP0TKimsx9X7GBXZrRSPuVucnpmJJ
Y+mx9uwMAV01OojpzORTG4lUO4GrxH5PRhK8PpqWfVRQApBR+fFANFramf/artBQ
`protect END_PROTECTED
