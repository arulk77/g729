`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN2almsg6V2Odv3IoepGIKqXic/+S14ctSE5mQTL2Ig9
z+LwAkGjKCjlPezOCJY2WcJcY3VqwVM6s0dTPT+qJ4yV5VCR65/063Sav4YnrMz3
tRiXsaozCWAqpGg3akAUJsPmCSWAhgKW4pMbRuQ5/b5lZEPCumfEqLhJ7r4c6asQ
uM6nNx8/Y9rJfl5PciME9v/w2Ncn3Lht+pYrJkJyA4U6GehnL+I+3ioQdBO5BUpq
uwwB8zxQyENyh1wH+ryG2w==
`protect END_PROTECTED
