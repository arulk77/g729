`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
9l396gn4v0WMqeUS3TXhTJi50IaWiHAkXRvtkxLKHR6kA1wExGfVngRAKcz+2N/H
Jx4zb2nrTnKQMmC0ZojXYcnaHsSC0bwV2/beiJ81203eC72sBIOC6GwT0ypY4dT0
HCMypSONkVa/iRxciACtVArIjC76e+TYf+skT81EdfNFhajlJrSSlKzaXxS0Xref
Fc4Ali8VSwmj7u3lX6Ay+mq5wgHhMNWJBonjPu/1qVKfl/7uCRqCvKqAi7b2Sr9E
ebWmIlVy6/ICEVw5dqNkJs2ylcBwHVINV/kGfZ7bcZs=
`protect END_PROTECTED
