`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF8d7W+YFhp+mn/SQrX+hhNZwQxCIsnjA34ez29qu9kH
yXx/5PIaE+2ixzTt2FsUse8R1Ej5i8h/qHe/j7VTWPvRZV6Bgaol1uMQBiUDNV4B
TP3eWSRU+XtRYr3FCvFvTRdZrbtcfXEEy4zC6TuSxhvN+jVWJphOby/5idxSO4cI
BlbyffGqF5e3CoqkxzDLWmZa71sPLwzu98/V7+Ppx5AjzSjNCrrX+qcuzojFRjbp
`protect END_PROTECTED
