`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wNdUjwV6i1ua3a9Ac3J1DBJQdS4Brn97pquxr24Sjpc
TpsFvfelmO62mNtTW9uizVLxnQS3doFkFkjNmSg9+FnlU2LNoEK8STwW0CKpo6ye
PbNO0Xz8OaSP9kH6qew+G0gIfIjXK0b7WTqKzEOjvEhCWCzMflMJI0nwSHpeTOP4
RswyO9jB+Jo3d9IPwjW1nGLLWjnmmBtCQBpB9YwcfsqLNto9P8zuMCflwAXZ0yTb
Eiy1+yiMNx5N7ayxhiQLBUWcaG0aRP26lrytHZMt2tlT7vGR9Wt61xj/puTDyCIJ
F5sYsLUGzxBh3lWOSVLRN0n2HyypZsH/rvQft2wSOSqh9nwxKTlrL43u0IqA+9zk
B12lhi7JNZJHfM6tThv9G9u9seEqdZfmWZZ6crT6jpjkFtHbdl3/xsUHuHkvG1Sd
2r+f6C6rIYrgUhdb5s9xIqwRJKm186oMT70nR2fWoa7HCga0c3i07L2+RIWMTrZb
`protect END_PROTECTED
