`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJv7m1N0Eim+B8grj1Ar0v+CEueVI5oDw97mOsMqP6eD
VDM2XZj7deDd/c4hFZiwy72wam/o7BXmP31DN/JmIn+kAxDkPdZp0AgVJajOuRDa
DIA6FsOyAl5B+8tMB7ONcfI/xLltC5/bZGcYVuJzq4VYpMat5rGak7sPPxALWiGe
t+2UUnhsqGEZdyqC87fdyMPgr207Kp/4dpcpvDpG4FJH7rn1COk3lOlCVjutrWul
SiApS9zS/wATShyBdYv/ZMSznGYb7gOso3sYlPO2jqfSDGtsbZ7IpT9QLC6CfYq+
ThIrrYiptnNz3QKDwmqyXKmKW3ma3RnMD08icmldFeFG5QFfgo80g7BcA2Lh4vnE
QTb4Uqn7JVOJ7z7V4NvQ5d6/qQJil2M5nLm0bx9UqDmhZc3QfT5rAnyxh7JH5dUx
a5/BiaYfeQLOUwbt4HgkxYma0fQRDBz0/9Ux41cuMDqid8Gad2wEWO/ydF0Z/Rly
GKiyzdO6QTk5dTOe9ss5NQclgIbaBk7YhVKoG+eWEhhm/jXKXdjsTXl/UjNPEnYd
`protect END_PROTECTED
