`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40vz7FZVzSw7x6zD2NP8Cl5m0Zx4ILzIjSWzfy5ZeuFl
lLekfthj0sMQxNwI+Y+DeIMrwLHI2R8oilO3ae6dKv71+qa6g4kwp5rlYAsDhu8H
p5wqWeLs+vg6Z2nkvTWoQDWgqmSRf7WTysh9p3HhekMLK++Ecn52Hcj3By7x+xW9
CwJBYJqAPh/Xx0T1rLI7TybyJ7BK5Z/g6AfEShuSQm2xpGo2L+eM4a9XyTGqPaDr
+mXAM/pZ2H/nhUuqpPY/nrGGQDtTG5XAOZH7q9MsQ8mZNl1FtkszW6tkemynk278
jzyu+IIF1bf3SsgZG0t7PaRy4OzTdz/ptYzzgrfoIHzvKm8EUQlZWIrmz3Uq7Y/V
VUNEJshdiKp5Gue+VdyPFh4li4i0uyJlrSWLJObDJOmhWHeFfN9VkzBlq2va1/dN
sjM26tiacL7ISV+R6P6jPg==
`protect END_PROTECTED
