`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
0bu5FScASrJloErt5HifvFYtWwo5BZw/UUgqCApUVPFjQMyO8l2lEvUfm4clT8xG
jtk39DOPhIJLKbdwhybi449brXDeqF/D/GHFBVjCfauSg8rJ5pX+fj1wyUE+7LcL
EAOvS9T+CQoJVWV3kXdbHWqIk3iDzjdAYNlAELFIbQCEjfekgJeK52auyT41nvUG
B92imzRUm5OjFuLGH6uLtS0XkbqRpWL1uDY0EdAYzh1KHO0OpV2c82aMfxqHlQ9j
T4AAjzWyBMUjelF6NHjkDak0sT04ydIVl3m6tBftnxYFh/PlQ9Oc7gmOXVE1WL4a
wMepGC694NZ+PR5JpeUUECyhgDWq7ScJC6yn+y3HoRkvw3uNhE29KyaFR9XwBycH
dAVL4fGUUpgJ6h47wwKRzrjqmPC10bNEZ66yqNH9xCI=
`protect END_PROTECTED
