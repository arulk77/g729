`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
hqQ9c1Fory5Mn3+VggGYywsMl+75evxbeMhoYuAFCElGPk/ZebUAHj5yeDC7VZeZ
HJpdaGPUNMLTg0PuykrNoKnj19ftiT6UbEehJi4IVP/GWy87W3Q01UkWrd9cK8Tf
5mALdjKsB0GKFoIMv+9ZuRafuLW2kRlP8tmaEqh1I0a/w3O0RS0xljyiWgQx4S4T
Qa258ro+dQ3/KLQUH4ibTetjGmBnBNHvNrDSW19Y8nxzTC92KXFTfuW4lVpLiqVu
RnrKr7GkU8QQWSWAX0ro6E7fn/Q6TlA21qX8mobPGV9SUkqAb9I2hAw6UqQg2s6Z
6JWfMzsGiXQ04EGQ//PocE02XtgeGGWz9HmrjvmLxS9Ic7C7wUdpzy9D6uMjVdCq
nk8eDPRPC3MxJ+M/c1pA9PwYPat99b4a9std9IFWqtqq9qPA6K4eiVzkHNQs+/va
YQvgbiyPb3yv/xlFcSYePCxfo4KqZQLUTaG1B9zifcIDVV5ICNxJpjIkPObyptDX
`protect END_PROTECTED
