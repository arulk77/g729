`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHP8UNJxT+MXSCDbt4+ANXxvIBEwvHgre4iEoTQN3qCd
pUDlZ0E9NbA8FFALLpNbXuwLNX9e/zWqFZ4F/zvtKe/DZPf2PTpmou3hNOnR3jC6
dd1H60H96s+qVOR9BHXD2qwVXcVtJ8IF2XO5JyJ0fXEYzwOMUBsBzpOY9l/wT3AM
Ijnxo2lyiyMZOyOfb/JTxeF3QFh9bTfNdPngvwKtzZqNcRbgUNvDDnzCWHACaMVI
`protect END_PROTECTED
