`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43+335v3/hOdzpszcXKnBn8I8C1BTnSFXEtrN8FDB764
o2vJXIAns4dgCJW3zNAXsg5UtvxiZUTkwf+i38MCw9YENLIy10j+xMO80b2dRcwn
R9trlqEOaLNGz56F8ZLCYpZ0+EIUW4b90a+k4U4pKKpfcTI22JYVZCJOwV4GbwRT
LrJGasLGv57iHFFrU1N0px4DFZNG3KeCcgeHO2GCpA7oJUxixsVcSqg5Qltlcxu5
jGwwP0+WnKs7wb6LjEu7vSv/nRqFNVUAgEG732ivrDI=
`protect END_PROTECTED
