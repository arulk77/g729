`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIMAryh38jzV8DXcARTfr4ZwqWgVv6ihPYMYh41GSjiZ
fSyKQDUdZau+8BcTDjdfHzGi2irYkDZv9UHVPlINu1JVvAVpnlMLJ6AaWd0wlYaM
k1zaUMSJfD4jMRMene2FW03ohcoqapOo2MtQHnJ5m4xUKCnXSnaay3cR4DCzkVT3
O8lEB5fsf5jxa4DiUmMo2bW8+hu++p+CWcdSm+LCLSh4LYKKleRgm2yZ7h1Bs2Jq
knXhFBYUWBor1wK0hoGDruwSW5SnsuP4tjlXEThM9sI/5YO8xm2bymldEB5emmbU
DJ8OudkbRd7KwxIwG4/Uak6IKJdtIXnA+Rye4ArfrdEFUiIE1Vs00FFQKnYG4FV0
fZ+Ryak5Sl7mNRFvGH6FPWeMc0OCacbaT4b+Dtk2TlT/iStQQUdtnqSWKmSmnczO
Y4SNmMRijYFFllfWX0E10OtjqVoAxKUM9v5uHkSg2hmdJm2fWYKuC0PnJ5ukoVKE
ukDvcWtNwhLcPbBx1Nl89TCbmsswSueApm4Y2Sp8j/C1L+I2E7L0b5rYGB7X5vd9
d51lGOi5Fm3KgrbdN+VMrw==
`protect END_PROTECTED
