`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDM7SO6AmlFP2HJcZcc4C+xWIFrvRAw1YgexLvTSQVtx
v6H7aO4yYrKSH40SskVR9XJkUOx440yMXml/JOyAN94Vr6m14QPy/qTCAPu0I/wY
sWkfxXc++JpCS6K4y83HButw4IdsSACcOMIYStyS1S/NT4pl94BZFQ0o/CCJZzew
pqFVTnnLlT49aqJNyURyqHeIR05/Ju1X72m0qkLYxQqN2rbhk51fixsB1khcXMlw
hCI58YhLM/xSlc7zoNzOgHorcAkfNtkkMFN6JO6QOZYC+9GQaelV08vKERqvWDEk
XvL/lg2YgNWQ5nyNoKd2lmiTCD7NqTeQ5Ovg3wZdfr9amwdRER6MJz7lMBI41J4n
ji2Yan/7uqcgxdeLYE74jJcCz9XI8hXNM+HVQTMdO2xSxByyZlhrzzrHxT6y+8aW
Y3NmRRzhnCew8d0ljUo/o0sSFIaD01pFt7c/jHXYc535NMyhJZjNFUC1CHvIt13a
aCeu9fwy6/lDvsa6XS6Q9jCKJ7PnkN7uS+LDs1g3oJyMN0S/kOyMdguSlhCA887B
FtPBkwtU/x1MyF0VlLgXdw==
`protect END_PROTECTED
