`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKLucIzmVo4thnjyJ2bfn1qwXIqBPV94Vn1UpOi+3cQT
KPaHAp/vTnO2q6TngcvCYok1CWoQB8SC61vonxmUeCDX5EoJK5iAeFPYaUDh1N57
9x/JdAhrrjgBvwpSrINig4Ozz6Bg1Wx9lpcCXnhxT3K/zEDeCF77xF5bfDSw0PAy
NCMIh6pFdpa8ceOle5OZAs8cw9dQhAO110AbR2KIYy/gwjK2ow/VFAiWQR/qb5VI
99FvnpDoMIqU3mCA7Vz5mEZBn8UI2Q5DYYGJdkzP1xbk8qf4aUvguJtDFApcIy/J
cVlxzXM16qUm4V/jnkjhsRymPGL9AwmxB66vCAxqe5Zdu9r6iEytXuULZ3G+ScE0
S/Odv2V60js9FvMUmdnmOi9YsFl4hSpupJ+/C2W3g1TKutgMcURQvOGeY9mYDncu
zNCNBZkXsYU8uFFlCSg5XfqwP4ggGohFXMlAY1Lj8XKgjeTNncGFmw2jG2mfOApl
wSYUIvuWBQqkp0cc9rKf8XajFLGbFh/0kM7nkO8kwqZUx+Op7l2RsvQE5JmOS9TH
VbNC45JHIcWxhFz6bbXqSmo9LkeBQla3V43KXOUyD934+sIZv0c/dqlmDno/WzCY
`protect END_PROTECTED
