`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
edp8+9mz5fVrbvFgF/ad+15IFJY3SjZJ13ZrBe/ICmDbDbu/P9sfTTGmFh8j2ppV
/nwXAL0XBIKTG4+D8GbwfSLoKYF6S6U+jI8bfU/CpRWi2u2wbvXRa1dZ2ov+n7ae
lUM1HCDQr6J92FzLkS4gpvxop78neJ2b/Goo90y9jEUjGWLtcPmGl3czE7uZW87C
qMSVgqInOMTuzQmXDd9r17+9VVyXdkrvkgbHOf4ziAorXAnx9HiyOI1Kjl1TXyLj
taSypEPboU/JTTDnnMtb0oCqqZoflTOxOnDoTG1sPg0wRyrSRXlDzm7ZmaRCgU9y
e70OjFKB6Ko/XUz6Sij8tBw/2Y55RDqcjq/a5beGSG8=
`protect END_PROTECTED
