`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40tGbMSlyM63Pev77GvV47dmnRiQsA0gtmq4dQvT4K9H
xTEQMPZS6sUtog1YDs68G23J+UN7TUAQOK8DXGgBiN8DWtCSBfW8w+h0hdImDxLN
Nb3/16y2+NFhAmEA3dM7eQ+SmK0MHj782NlLgjVfYywn8Nj+ENNPvO5gEnhKExa9
lzWd+v5G7952gdeFo+2Uke9IcznFtaVENcmad+ClsduT/7mpDd3CUFFDQIpFM4X5
8tuBy1+Otn6O6hSa6D3Hha/FHP5j1LF/k256qvbi7TNLJnXd16Zcxduc9DfXo1Uk
zDEzenTYhtj/vPkyd9G4iTaHtnIFhPBEklhPaTfBMak4y7H00Astru1dhG8JOpak
TTBf6qLbgXs1gOnBMgMI1O97cO1ALeEfWeKxDvO2y/BEwOko5HETgfNLqcE9tnPv
BPAe/gkKhUU+WBwhCz0iblt7UuHSj6GtUDFLbSLLiRymg9EX+CiQYIe346FZwJxB
`protect END_PROTECTED
