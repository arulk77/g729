`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
O6tX8V5i8XwMokRWGsAhFOlFuFg2mrV5YbqQ+5NIVzXZiZ1Ohh5ogNvsbEbPLnQI
Q08Yt5HKXHn+1X8NAzNlHbEO9zGuuy30kPr8t7PSpr0ZKS8MtPAl0fmsfyIRS/Bq
7sJURJJM3r7R5wfwA5QgddxQQ8MBrw1UMmpLZAQf5YI9Pu5x39FpEOQOVpAUUNlY
SokSMyFfVPYFQjVKZskA7uqfo8VVVAov+143U5Qxjri5NbTFrSdurBHWsK1KVHDA
gm2MtXdB+t9U2Z2jenmHMZlNyqSEHoPSpr7I0wRuYiwFWHSgvbiKIQMgQcEN5fV/
JtynUdq/lYeYEQ+hGNw1vDHnq2bSEU7dCrywu09AswZQA4245sop9s/f3R+4WnKq
itNQ6xr4yIj2lhV3UmNnSPPVLPV57jhBm2rStHeyVYz7+NKHLRU3HLxhSfU7gXho
NbHxhIXLijVNIx+U1QuUYl1SAheIJpqyDLE3XcGqyDKXtHEIVJg9AJtIjrB7vXBm
Z74pBepCOcEFGhzEPl+gDwLXiTQjvpfT+gbCE/o9jWkjM91+/dAD98AJgNc7IyJ9
HFLaAT5mzbJHbdGIWUafibkj/lgkfHp414l2TIGf4fuXkgWgGVb6es1EtUNtdekD
K+E3GSGY14xowgXw2aheoCqLuu5SHvmQg8ASmq0qvfSUkVnpoVDYCfMRMsEyBfdA
`protect END_PROTECTED
