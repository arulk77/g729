`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yIxS1dtYD3kXN36og0HpuPxZI5WogQio3emwa6owAjk
2RNRWWFRYpsFjTA+H8Rz94N6LNGvLcXcfYxoSYOOpNXvZOLbDNyNxGnTZSE4FGK9
CNWWtLcmhJnf7bH5IRGOSg0iplYe2On29m2XHi56PatzJt3SdAfA2pRKp0MdeuXh
ILl2anaA+Nw8buS1iZaKQEkStPK8DvXU+prNNOn7zAE=
`protect END_PROTECTED
