`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45MIAx1X2IZ/Y50a6Oh6aszrPQL13WxzKU7wsFMuQMRU
zouJokhozJaKeZOQu04Q8DsU//vZIAs2sJpT+QQQyiHFIq8/Mu/5xqqE4fQW36dU
ibj035iwfzDpMvcudSzZT1RF6RSL4W1BZBC8554FIX0iFhHuzQ2paIPMlFvpw7LS
Sov84Kd0a8YQB1C11P8toQ==
`protect END_PROTECTED
