`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73Cx7S6fIYlIp3wbExnUmwb+j8329PzxK3kl2tGAIZMOf8
zfd2LlD1455n8hRCZjIqpXu6G4z4fn4Lb79po1S06HUppvF4n03BLEwg1n7fjxPn
Ct92sSiatw1wuIy18Hoh7hRcPCKcbBvvUrYJDrW12zPtr17S5VmIHZaYMU5keGsf
NS96cJU5H+vb5AOEPz0kNq4d+XrM8zkwceP2yCBka2SCHR+guftF3Ec1S7jLaJXK
Fe0J5O17yyeoxThU4LCIALLVAkvBU4PKP9meXphIlLzFbBpHmdKejy8LFFpM8cHt
GKCkrfqgQ5afY0rnueN49hGS4nWuMrnsQemjFtYDL9oBLLnMV2z0VG46ZLx1qbF6
yuzWFKZtPay12xIH8m2qJ4/HLyc+x8bLWklhFjUouDzfwwGiQba3FHacyJRixMwk
ZyJuBkonzPthBOoPdi9MUXV3c+aLYN+4u2oCCyC13ZpHYN+Kt0UOjoovt0wB82ne
JSa+MjBhjVRj4Z+o/n7Tyn7llmJeYy9WlFRAapZUXhLyFZyyrCTZwSLVh2qZaHE1
2/yPLIEeOdAdWynT4ll3Llg4JgeJT7ASM1zrJgTiXu0=
`protect END_PROTECTED
