`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCjKUoGT7dHURt3tYKoDxh+mU20Na2wd65E4ZEiEF3SE
MYwI8zk/dQpYDvEkbG7qCL+lFuwkbwTO4sJbh8yLcAomKQGy8i/hQvEiSYAAcu4x
YW1wLnAGbQ8d8YWxYZdSHJkFUuAyzB3fc6r2heSZO7WuVkt+138MFAKrBSQXqDQk
uHN0lRAMAPsVLfP2e3lpgCDKMz9/JUYhtzNT64HhWpbFBNdYn6+28i7zOEoJ095u
+nUSxu+T8QFtDtClZfy4Q741aNywsA0iq7g3v5vqh2mS3nRZY+sz3NQxgx4RcEtg
YuYtcutgGI32yGh+J0QiSLf6v6FNgtTRAwoumbw5OspKiDCJsVqCHD8kei36W6nQ
bytL6Mj0f9aF4KcYmmtRixwHNsu+3SBbRZJ+PbNRv4yI5psYWqCNJGVwjGxRI3Ra
4OeqVs0CflOab933CgxrS9sGok6rdX9xdRF+jjZkxyC3tyiCl2CMKUPv45Bg6jrF
UkA8jKGX4Xr4faI/dBlKl6JdOEBG0hI6ZivJTJQFm41pzeVNy1hiUy23O1xCVudF
6w3Xt35oAUv2zlRZoKJgcAbLOuwpb4aapSzCMHGtDbg=
`protect END_PROTECTED
