`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IJkKReClnivQ7hyAdiXpo6VEI/+en4DmNWTj6f0wVlBHtbTKCddSnuVuYi2qetJY
pVYH74KYFr7zhFNLJuPCi8ITjtjowm9cu/XECTgi+RU6OIBiXuXjF4bgH+JseJZd
Z6mNFHCVPt7AErWWVmgKl1nN6uMo47VSmBT8YwiXEUY=
`protect END_PROTECTED
