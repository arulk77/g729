`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOoyoq8xH49T15Ep7NYJ4xYRzdjvKfJL27r8lVnuf5g4
NP/O9wPZttausRPDBMfH5dCMV9suYJkak0eC1+Hb+f3NprO17BiAO9ag84ojrKWX
6ibgX32QCgOGrYlBFYjZ/BKjB42Ov2VcS0/s3sQSqpdh8fEkR56kh20EnqqD9xOk
+52ZpGkPGCwBHdi5vcLIbeFgpA1IHxDgdOulH5pXtQY8QQfCZ0sIqEc9Hvbxcfvd
X4vrlfGrEoiocze3L8u8w+GRGcm+cJKIHaAECJNKNpxW3jey5ZkI47NLth9V9ZRj
JQHOBZaXaK5lttorAsUgJ1qG58nFABgd0wtAsZFYZ0f6EN4GXUnJPNAsdVwTNI+7
IWyrDt8psuzOIEX5HLR0WqBb+lNX8Tu3Hv8MtsXjDf2IBlViD3LbWYnRhvyznto0
N+nUc7+UuF+lV4T3MxAri+hVcD/DidUtgSoDxsI1v+lrLHXkMJt6rh/8hTPQc107
7vJSJmLZKyhuZQtgsTxP37tlAoOz7EZA/5emLYDzNo4D1zUlYmaBpwVwzNgli4ku
onM0wJQ0snSRo50vEvh0Fhi8ZoshZW/VfQxPhk/d1m59AilvuDb8DvM0PFaLilqO
H5iWNGiOS+zPsGwX8hDXLmpYKCw9gmSo0wW8IirKyRb/5nJyUfLWlJnkNu5iDgob
zcXdzDt0ziuE8MJwBuDhKsBciLw2sMky/yJ/FuD6B19RXeQ6168IQEG8b6OlM6aL
`protect END_PROTECTED
