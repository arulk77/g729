`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C2vEUoBidMdJ+8nmWBQseNhEfM454oAsjpmrwhBP6VP7
1VSpPQFf6dNhSj7bzmaCs2gMXLUV22999Pjwt0dRfz0Ug70Ra8LFT7YEou6hqda0
LheqdeSxqFdQM05sMZW8c/P2YRZ106bVdShKXbAnRM3teWfbE6qSYHNsS/SSxNEp
t/T9WIfsV2Mk7anRH0HJAiNBueXmAzuyOTdf5k9LHgRov82n2im9YEwwCKDyOTwT
kpkownzp7FqFA22DHyQxtur0ezM1rvPoudpwLr8qJMUbDqtRVNBu9g3b3htedI2I
7gQP93XZFZJqrnE/4oEnImbHyIGo+YL0uRpK+XgQvFb9exuQKhfSk2/Gt9ANscZf
ThDXMsRGahTz4uhU60T9fwZQazoqUbjkMPHI+3Dtq4EXGRrxLaLzp+cRWdHecZII
`protect END_PROTECTED
