`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIUjuqFCV347uzpKAcueGXkbQyF3rBPsP37frYSKgwKF
DD6UOqqpaM5IvM69w8cdAY2hZTgdzSyLnVlP9KzUU2gF0/oLm5/BuICt6R+HYhXG
w7OozDmA5Ow96agJDVy8CR50AmRVedxcMnobFis1T0sG6wdcaVawVmz14SbzYXoZ
iP+Vo95zJdgo85LkPgje85Dn5S0e9cwgcv8wxJUacY0Ntu7dW0YO7iu047dSBNbV
QXNhr2WRrISvgl+KfA32xaDXKKLcHOkt0ZRgEIsO8NIvXKJs/CFDvJb/X75EziXC
01z5zMjPOP9ChHukJ/PteXbBOtQTKdJEJtCmEoyi4RHAaetiJEKBX9LY+Zxo7oWP
`protect END_PROTECTED
