`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SdlPG3PedBW8WMByA1mQfWAm+WbfrYEpXGuy+BUGBY/d
F6pTYJzFqkQm+BAkMf60ZC/pW66w72ibn4zmgxMDUU3S+PJBqU815GRPPPV0jVRB
nl9XpFX6mS29wucb+kXrh5qIFo9U5A4cVmqMrSqH5Dcr1G9dmMAoi9I7WRcTqhLP
oN8ZJLJntW2AfuMJOC3ub+JzhzOJ4tLriIFf4WAQoONLDd/L0162eTDM45Y1xXgJ
oXgBQFnF/ZuUq49Avy2+hdAOiPnyTsABR3cwoCnEG9CuVVjloAexuVUU2GTyj76H
8nCcMCIamks9CKtgJdQbpm0kAj8xZeXCt600Z57bzdaYVzERuf6LhZOyxjkH7KQz
SRl0K4r7jzV1RBMxo6Dl+dFagg/m6aTxyrPk29u09VXrBv0IbbhfhZTvBXG2ZFnG
jsEuUqaSkKUmGiQfCGLiCYc/tZqJPwOBFdoLNz1p5C7OHvLX+hSlKrnUAMkE/6j4
XULDLZ3KkFZpn3QFfYCdAbD3uLlJWB53hQiV3bn+EjogKO+gsBOMJFCVAHcLewov
01AkJlfNO2VX3eUS9PJv8vNIFjirju5IdnfcyGdR52Gbf5u6u4rXTZ8zvpO6Yape
Q8yuUs8Lq/6d+UY4USCs6pnWI283lF7zF9MHahX6i7xxd0/KajwdFQYoyWNsRlk6
FGFE1EjJiBtaJjPCyXW1b9jgwbinsKuXhqAjCPa5qd00p+eakqj9rDNBLvnufKa4
6CwQLnpZUQUqlqPYwMGWJSw3EiWAR1fBi9VuVIFaKKCirbkW2D/RK1FNFL+OFUuC
bwNzSu69QsC804JP/8JtHeKzaNwMbfybm0Ut1qTbnLqno8Sd610eoncZu4nLBV43
sNJAa6tg4heigHXrtd9Np2bp/OuINpE19jJC4wmKZiE/mrkgWv2Sfiz6fKmEcFum
nKHszC93CHzCD7brQEGwlOe7l5OlmnoLHyj3a0XlwfEjReeXdwqF/oTwz4okF/1/
JCE++jHGBb1ZCA6ZgGlyBahaY/GKlkPBtWQ5lCFqiEbjrX/QafcjQ5F3eFpGCBe2
cqTH8+TyR8wPOlXWUPGfttBWOdu5hT7UlX7YcdRKGGN3/vhJF4mTZWlQMkScmioo
ALiIcBWrkcgYittHyeL+SBvUgkw1M31T9VHSbvNZCi7roaG2j56w9XbfXjKBZBz+
EvbSVXAU+gbeZ4tIp7lgNRl8Ez2JuYfzXzd6MEun0fRqAi+uSvjxjubJfIT2owlK
n9yPwMx1lrWFArYPKErZeE7ZYpxLDqOqrEjuEoYz49ifgwBnfITkJYoaIbho6z2Q
93XNYsoxn5F1fk4zFoQo8w==
`protect END_PROTECTED
