`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C4nbHx00p7qQmvDRuIrSaKKrfXWuytDeMdf9fyRClSfo
Oe3KLSFJkhZlXMNtDUx2rc66Tle73f3pxbhTyXzZGVowWfsCoXjkNjoXEm2ATB3f
zlIAcJtBC/7+4LEE3O9YZWEYdqMVxh7XPeVawbktO3kJSBZ9vQprkCjtijtgnMlU
0LSDQw/W950LurhesspZOvH6bPAXzcB9UDkATWZds4Bm/TpGdJpwe+7sbaEENBDM
PvROKTxrm2P04Lu3VKKbgeOOj73UwQ9tP78We13fjHBBKFiupxB3pvkD82lyHrBd
LjwVh8eeMjEy66rsatYE7BhVyaDSO9zPxnnNHrfd0rmLgD7WBzpwvYtyYRi1HrPg
XnPRKBjVk1t2+fkM+WGp7ruCZxCFxRGeRBIinm9/DWxGZaK4ATXj9Sixj+mYvqxV
6w7Zptd9euFQikgL/YOqafzBOES4vAzomEKj+/vFhWkyGFvqpMLgWuTGEozWhdLj
LY0ZF+uzPoCclEFKDi2fjm7DELmP/RRyNHkjOCydap7mfpcalk4daVeFii9rBlJ9
TL51jrQaob24f4hgmkwqmXpGO7R2uY/I+YYNfGQolH8=
`protect END_PROTECTED
