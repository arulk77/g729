`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yeGg+WPk9j64IV+6DVg/5JBlFvXMnvK9+Wl6nxJwthO
HBVnRxfPflE1T1Ju9joSKwCkqa67ukZaT/kFgUflS6axWHY+NCUDuo5eI9JuGd4Q
yKgyDFfa/DIgkSPsYqZRedv+juUWsZvTVAn1gTwm205nSJK55ZjxGyiGxMy2omKQ
kuP4/PhYalfljgwlLSa22qpUkLHS+mJPd74NkhTPc30gsuO6RBUpsyW59+93MxEe
q6g+I50wKYkiiZgGQnvvKf6zqhBs5F0B+G9134zdvRVRCrup9xFMeaeYkZTdHxrm
F3RePJOPZOsVozFW8Sn40g==
`protect END_PROTECTED
