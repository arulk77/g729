`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN0Q1GweRA/TODb+/3GF0FTKiMK1QBpS4L74r7+IxLsYq
nYg7BBVXjXHeyfzCXNv0ak0WXMTuPJpmtzyctBzrZOdBeVX80GS9II6f81+9Xglf
jL3QVYJywOSD0To8JdNqZ8fjJdQDf5cLowjdHXXXauMkRWq9hagkp5ubFErZfEUo
oyMU2aGwVfjarOF5zKechj3e6q4EJdZfQ9mumqrJOzeAnBV1x0IjqLUTZiTXkCrd
m4andTdHHR62I3g+YyEWpcU/IgK1ChFsVee8I7u8nSFYjJbjiS6fQZ9+1P2ECKg2
qtOp4DZGpmLiyoKidKSXz8+D6Avv8iX/+jOgNHvziXUz0SAjYsF6S7XNn2sjlxYv
aOhsiShOV/Iw2rGPDy2HsiOFy8XJv97vTDYeKkr93BhykcaWsmczSzEExAZcUdja
i8TGE/ftXtG25H0pzb5UCv+R0cjGvun26mpn8gcLuN/w5zw8qdLryR/mZT1qNYKN
nbnB66uajD4zmOnp22cGOjLSCBAuZoW3AJ3wO3CXUlTgsyDCM3sDq582kJnpnIlA
c3hzt+RAdmxfT8WR8ZxkLCfLwmgDHchgeYkKne1kqvC1PXkPO9+Le95Ig9y+Jdnj
z+eH327bj6PhegGYb3hURDyBuVpC0Byj6RT94HG4mk/F5BqQCyoErVQz9DZV4b+i
nd1w/85QL3aN9k4BtgicD2/NS2edWO5W5HmflgiHEY8bzQpzmwH9hY4BMUOt4+q8
1qZgrTbk/YLnZhXj5lhrfirRLH5KDkvD92RpiZ8L/uMtvhBNUSNJ1ImtFsUyZtsy
DlFCMHU3CIh8anxfikvugdKXZ6pDVuiMbW8KZmP7pQ7y7d1I6kGONCVpT7bklRj/
cHvF9YYHxdNEepfMOLrj6mJnLkqZES+CAqj+2dcwmFgf8+VpH0t+3in9dVDLXnNm
zwLr3a4zJ5Yswd+ex18BO9x+8G7SuxAnu8b652U64qwaYbPwReDvo5ieXfkPjZOj
3yQtvhs3agh44rVkNtBH/HvT8WQPA8Ok1r+Zq4+YoIpqlhV2QE7ZOTm9gQJdVqdF
tgaY8w8OP54uEnfm9wXe4ArCLhN9OvYFzHCsDHD82G2oI34K+XseQmwG9Z/7PAD0
JY9JEGoTOcwMVFWJgqJLxSZxzTGsAO7i/ekz0lvjoFpepk1k5HNRTMCj0sDHEUq2
1Z3o1SB9Dh2MMUp78S287CPEKV3kt/+adkrthTDO4/drMQQpauzwcSFKxU9c0o/l
TN6k9+roiCcln8uaht24tVBpvfUZ2m8ZOM1xog95TCq5+jLOj0PTLzM6qG9GlnpK
UjKBKlEqyv1yi+PMw3ZfZSzZGOTGvP+ebAaWesfHFMYJL1IAPsaCyeigwaARwTot
bQ+ehea40OFz9isKy+mmO/zFwNRSGvO9SAG88mjZL15bTu5sL26pdo1gyVA+fPQ/
orMUbvi/PDCtyEXaORtdpHi5BlvXUIOViQOFuqKJ+aa8LRCdY0yb4nPxvP5orDz5
fnS2i9ly4gUO09YV96J/mHiIfsD9f28xWu4xmMSIfJbLbYZZ238se1jN+kDWoAb+
5FRz5lbtNyLhjSAXxdPzO7OpiDflLe+CW3Swz0x4ADBbolW4bLKt4ND191BxXNns
uO6M+jyG9WAqkdFF2tEDnvg5MqYrdTZTQt7nd+Vhl/f6EQe1cO2YSHry/FGSbuv+
FmUCuJYkTBsvyoouw4r1a5g31obJApPVl0ezUAwAhRxEQJOovwA6TfuZMiLgQpYF
NcVgL9uXLEwIbBFpyrRhAmA/8Q5X1FZP6NVMl0+VsnWrrkTXf1Olk8LnL7AoK6vH
zfjY6H3mSBEeSqGr4abb3A4eRNbN0GwfsyKqXzkPxZFPj3iyOik/n1F50ZVX8tzJ
brmmuVHplvruZI9dqigSUdRpfyvgHq7n4TB0YsHQqmnYxJlfqjnC5gO95woJ9YNo
/V/f6Vor+gYDQ/3JnyOZC4K2vhXghNOR62nL92ui7ivzRskd4obPiu5g6dzGbn66
qGzkiTdxDP90y59WEX/AzWW66h9xEB1Etf4p69ydJTJvEmIYe4PCDND6qIDG/tWh
Tbvxm658xfQi6sffsOfLslTCeD6TPcN6CcWwJBklwjUxvbaGmDD1YSz4nH9Qg6ST
sLZv39yt3OdclbDGo1ZfHRZ4ZG8exIITg7EuCButu8X39F+lKVHpcNlRgrm8hmWi
fVSGeFtcoIG7pouxk6WmARIjivmC0I6p5BHwCPaS1iI0TmbUoR5YUXyCn+g15QU1
YurccfyYRS2ew1O4CUk9A90rqcT8gz9+zTcy6SoOzXDSy5Tsw7N92kzI9lefesN0
Cjrg2ZaZnXz+A5H7KzH7SaRVjxhQK7vWW0gfb+Fbhphrp71wvyn9f/vmS+Y7AUFm
OVQyOcSlMr7ozA1A1ZNlqkfJr63m5Z5/HOKoZf6kLD47cTuXiM+XtjU90lLNGT4r
ILgVIkgwX8/Rb3fNksC0c+QBYPwTZBfJYfCI6bGME7NdlqPs0TfGfhTd0M05c8es
np26bZi5IHuSf+R4tlRG/yypKOiQJ+khDQmkLAqEP/T3Tsj4b2hgs4naT7cr+de+
O+zgB+UAEdJIhPMTHNFecr7VMJQ7NXdTa3IGX2dWMQXYtj0lfMf73bi3y7oubQrl
2mlWMfOgTdTbXs07VTZwtfjQOUDDyChxzMS+1/kIBVowMPYtRZvlhnM3GUgQxxvF
XyReROD3L8z8ltbnMcMaxxxsxd6aFSHyl3l4EDi1+W+uJCutJrM2kFPfBfuOFJrY
dZDF3MZpTJu7gQ82JaK0mRKpWrIyXWjsC4TvV/kM/EPBzJNcTit15UA1XkXZUfBR
esz9Qv0mxYDF2hhZLG2S925ApgmS9gAPZ7kBpZsavsK2rHpibQKHH+3pSrNocmKw
9kdFstRuJKhjw0aiSU05mF0cWjCkbtRKaaVOq0jPyNnQb3kDfa+8V0qPo56RGV0g
yx3PjkGfy/LnRjPoBuaCcA5nRYL0mmXiD0jmI8JC09AtQUhkUyZkBiw/GoHMqaMG
iDiyOGtR2mBFVdxu86ChYkH29XkmqCorQpsM0RgYS7Uf23cZINIo4en8nPSP7BwA
FQGbiA8XzxeBUx2q7kn4FxzlKNpeZUYpCcjhnLMK/iS7p3enuDFM6pckDF2I6ZHf
3H9AZ/k5fex6YJDJT4lhQx51S9XKI5AGnIdebpI1djwuFvT8D4Nl33eScttq4mHU
NqPXsy3UYF1fb7zis/vBBIhn87vPAk2XlON6/SdBqSCqmTTKPqf8kdGaPVuiLyr5
hql3u+k2J7XE+VGC1//7bhRXZD8P27nxtYDMskg1+i2RdWdI+Xj11yJOMCa63jwH
GL61hXdyMMG42egq3EWVNA==
`protect END_PROTECTED
