`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKgQOnn1j9A6NvWHQ3Ln1SNktT3Lo2lFFe37UXgobwQP
U1JHwi8UYkbwwBH1RVfk3zE0WpPezlYtth+zYPP/aRgt2Cny2fdm3pggEntaSlYX
h40X+FGfuifJzzYzR0mSNPYOc2NJwC4Dmt09O6u+dtjbTuVlGbZHpdvMdOJMiJRz
ePMZj0iGqIXzu5XpXMPYBE+M/LAlZSeUpXDWl5kVFM0OQXzMhNQdhlyDqT+Tzm0l
1lD9XoOcguCbNYny2n4SNdbt7JFNLILK++r56lq3WpDJzJI8UWBD60neon6Vve05
hUKRK3llQp2GH3VhbA5awvq0e9l7RtGCS5M8jZkIheD2arWuZ5zHD5yDOXFRFWPv
K3NOooGVUnT++69jdkTZEvuDL45qqf/uIVCbXTNtMorUpm2EPZyXYlm2pdCa1Ena
M101qxVoGymsBW3JxEAIyB118N21C5akjv6K/0Qf4vZvo7UCIDa7BMDQKONvemuL
vJ0/Rip19aW6JLTwmAqJHrgnlmcO9hK3gwqfPN6AdS9ISfzw1aPslQ5TN7OTz2H8
m1HGiV8Z+51dGw/WXo6KGSk45jjBQorWXSMk4pQw6DR+O0Hyfl9sPzjyHGULVxJt
DtoZE71T6BpB6pnSlJApkUcutIMK2Dx2oB1tyVxhlMSFdeWVq7S/CPIrDgStyuJN
yAUMMHzLxWxtrq6P+ZdXeekUWjCTHmG5vEASXAq+/J6l9apgfBfWdcL0bL94kPez
pKtyWmPb3dALfF8dRg7g91hvqrGVXJ6ovTz/KuubeVskvcz54Dy5UkTDhAV/3Wrx
erqrV5P39vBUTZU8wVHSlaimTW3wHi7rfYRw8Fwa24sPbkNs1w6UzZOBneltsDqY
7xgVIOboOCegvh+X72/BD5+kpJSOmRBhLectOm1otsHPT4eR7kmaUGZyI8btu079
NrtyHsXFVAKCbAD93c+IjhTQ7G90fO6St76HzMPGiDbdFWbnDIlZ7UlQWhL1N8Tb
rLASt8P4IxCT9StPnQS6FvaA/cFb8OewVb+C892TafEuheUyN8fmpUXgbfls0rrI
0rEN5yDXS52nfwbMbnlQOD9p7DqbD/UgU0SyDsLaLtixN5ITxL170+rnjlrXhHd/
RzVhaf36c9Q/5D4b6hLPrc3kuaZN681HHGMLeTYqVy2LUZGjR5VFCqwZxRVoz175
B/DCZ1dYYW5BMi4Ubyd/wi4lHsf7MeysXKTfqzSNlK/CzUIasyy0e6fDtilvH7Sd
QE6kj+6pDBZpmp7wvqJr7iw815EzPDl3uoIR8ReT7TOh3xF1Fjkx8RWSpQUPW5yp
9WKAWTHtGc2wI4hXq73Ha3HMyj9ZfjkeR+BWW4RX2W8XAYBKA5QVAY75VytwrHCS
PrD0yqBW1OZsVR/dEWbccg1U7LpHYf6pXzoAIgGDCB7OTrgzrKAEav3tUWCxpUod
GV5ZPpacZ3HMuOBAmvLPcos3BH4423LbHvBNxMLV+ljKJJFnwYqT4H0PVVf+jd20
E0Vpnw05dsTA6QBSfz8bVRAVXk7dRgIuw26qVGJZkmodh6GqaQz9ONu7e0O6/y45
Ozv/yhH2idpHK8PgogMuqNU3BFWhahXjVGwORKNAFghpNazrHGH0YMqaQAuD6vfY
cNBokPKhs5fxji+WFE8fRrZy9ubnOefwtgYU+RF/nzfE8rxsu6zLQciEjM53KT9Y
exUm9LSK/88JIgVb0lCAB5CgQ2iCnAaBW06MA/0P+qJbTzgzNIQ9njrpZ4oyxWK7
YUkhIhUeX5XaVOWLLN51p60EPMDSYuYYDH//O9VI5YKsRG6yirr+oHv7FGB54ZYb
koBr/ZJWVLgF9c6KUJ1r3+M4UFWXzMNeNADo1Nv277IhMiEjhqZabLd7342rzfFi
IlxsqwfopTopZtulwAk2FhUMyLb5480isHfatK55gC29vn/JMplDLB2GtEsIuSsQ
MGMOfuc6hOKfrNvVy4NNb/jFAbzm5WXIG8XjwSE1dMlliFGqrNWYsJYa4Hi5nR0q
P5zwiror3DzRcRlkrMN4arobf4EuX1k7lgqAZWkWQ3PdjYTwAyTprAhfZBSfWQ82
lXnXAGHFwWHMvNVepwKuBNkc08iKDNBs5IJ/2FjJUM/xTrG7T8lL5VdfQAHAoBTr
7N4jFaBzqfwSRCDRUPnITOel7PVDNU1Jjj/mj+ka9vxWTFupB62tTnqhd4zC2duU
UKZDOPKyqCzCeJspXfdgY+YOU+M7PijmePnXiLy7fjy8GfLx0EKuyO7lp7/qFe7A
0IlGMFE68+O5yKUhMbjhY3J8+cFvPdvQz2YgyI7u/r79oPxb6mLgPLhdEXvOPMjl
lBOjfBIdzwtx4s0vM665cvX1DgOeAk5KJ0uu6GWAWeLj023POgOu0uW+tkixvE6U
IITzw82eDsbSzwJ4bSdiiaJSc4BYDstDJINKoHPeO5UhkN2pPJqoGD42kvOgWIAS
8zRR0SSEVkUjofq3jb1kRUBy4+SaXzqUnTtOrz85CsABINm5HpR5h0XdTkOWn9l3
46QkaCGhW4MBNOliO/OGT2x9tdW0/WPodDhvUtAv4BwvvSsqft+/vkITb5eKjsr1
rSVyxBvqR6c92p9GdUZljWLgAUhRWYMLpsxo846vsFd1hRlYUc7GhWVlyiUZVzyo
fxXJZzC7PG/NAtMtZ4UccnlOjA+jYwu+kD+JvfKgGOLjs3t7X8sWnuUpItnBeknc
TeOWnLYo8Mhu9zuxBojUXVifT5o1h+uohhYbf/0zTjBmrBatFFbmgGnVv0dV6/8y
JfMTekhsqxb05JEz2MNj+3d2FiOdMiCIEFjiFurA/Dt77oANNlV5blG7GVukzuL+
gZsB/dyoftIEeReK5Ul+HYpS9yYD1T0yqH88qeaFEYgPK1n7/+r8DEK9yMcO4Kig
kjKiUifEQweFfONkN1qokZN7F8py3jONcon643BxDwBDXV4IuQx3oHGCLDWW6G+x
5DoACx+AxQ/QqfKAtLQSYGWiK8w6OJ2D38cWINWLUqE18bpPC7gmBU7MoFe/h4pN
pWoozcvT7tGqG3t6G/bsa8Vf+qRFZBmocLswJZ8oPVGNUooryNeOt7XkB5HC0y6I
dN25rFpGVtPpYvC24+K11Zx8HW2mquLmkAq97m1GB+TTQdGYMi8nNCLpRjsvNXt1
c0TZlEqTUUvSHuegPrpTeiY97GKEW9i52uYMJe9bNilUGu65KIWj5oGjmGxo9C/w
bxUk00HPG1wllkLXF8pjGCVTiDYXRgIfX0goyczDchdquEWku4edsNLXMwSgIZ01
lpmR73WWXeRYhdPh+aVENjBz0h6MAutoAZAfi5PdfYuKcS5XvKNnQLB+BEb4zDJy
awXL8IgkPsmcegrq+wD+2kYehVKgDbtqi9a1ZcuDO89mnAeokiwXqogS0oAbBWvq
6nt9fd0uEuZDRL/ygDB1Uz8gn+OnUXxBBmO84LyUsov+lntRSGRnJzursjPFyHJT
RuM4hp5LU21psN9WRfniAPozseSWTaVkzlyy6Om6vkQqmNib5N8k8ZYbBqjw+L6O
ERpVXKzi2ra49x6kZl9rtx6OOHw94Z0+78nT1sA14iKCERLlZTnQoNMZz4ajsqmg
GUjhD6hK6QLlxMZLzOUMf7FAOgU2++WhljvB8jhyaPQWAx7yLPKcaIxpZdzcdBsJ
6lPW6ZQ2Vapow1EPKVtwGmhqY3/QfmihAdJpDbJuAS2y2qrnwHqYWCNuoET1ZBh6
kcWv+Gags4LSAHKqCeDjPZi8v1tgl7VsMvEZwIuasakxMxXIBcZTH4u1YFPoqjgQ
mVnmp2Ci/ArKw/2iOLpEyqLi9EnJCVa6iq9BsT3u04cAwANiPNwKVekf0H9H4iws
SoGhgeT/hI4gRxJSDmv0qHatE7dRCAFapF0+AgF9xEnlvPqLbmYwQvsP0xr2b4gh
hYp3uIzWSTpZzdEUFWVyJlbJKl7h4374dbt9M66UBydyeP8cr3hUGsrCarAjGk7i
As2+uwisuvBjqk6wVHx3FHjUlxXh4fbEB8rH6Rs9xXl8fzTVpUU2zXxARnQ+cxqR
wOkMDPCGrKZt1tRJl1D4WFve47CgBFqFG3HQBV8bIkaVhpWhbXS8OFr+Uf2uclxE
ZJKYX3OhAkrBC2hOpS0CZtf9COHb9wMzBUCg1ftzzZzbBi3IjnQ1f/h3m7rwKihq
yv/1etnTAUQ/v7MIadEPLLbO7EeQzlDIp+4FF9TLntuGEtwHwbDJuq30pcdTGzdQ
m5Llgoau9lqDQdJsK0yCeBoix2FqS9H1aDjYRdbpoloJE/GHGM9J4gScctZBrdQn
Pwda6FpfnX7+jDB7/JRU0OXkdq4lf6/6zfEILQXd5/snPyfipuKyXZUI53N5A/Bk
Kum8Inb1/bV7ezo55yi1MDMCYPWib766CgNaD2XeQpTVdSxCArYViScRAThie9/y
8JFBQF+gN4SGuZZUEx1hePNEpOXZdtHEzQXeaI/zbiSyWFyfiaq1YwLn38Ip+OOk
SITSf0BG231oOcnpVvaDxCxvgReVsIFM+Nj+YSCLiixbIC9dJ3SdI2MA3/8+FO//
xa89t1xDRmS9SSBWgy7XYB8L7UOZjvxPgz2oA3AzuOIil2v22MAMLoigNeQjMMeW
aSS+yLHh9ayjPNF3Mcr5S3P81Mo3tXMp0kzy2KkQ+XwiXq+Clv1YeDJXIBaDHBCQ
RHN/MLAmXtZT+TgYbgW2Kxfoh3VBdxfG07yLZofbJcJYY01cfNeGs3CQFm6RomkP
9P4NBHrSo7R13eAHDjVM27YGPW2WYct0fAn3jEGKc6OSOBoaIgOuZAbLOdDuCd+k
KYfZ0qGzMzES/6jBusmaaSyE4B08oY1XCvohmjANlaT/MMuo0FGPdynnOIVPEKfo
XKd8ZzQ6/aMJw/OW0EimHTEg30ZakhVb8PWTaEzljctZnMDTaLgP7v1xylGsXmXJ
MwMukoyhvZeOtS437DyIGcTDpaLaVJZPe7PNTRzpZkAPr7JaIv7I9KaFZoCwSwNE
P47bgaj+mEJ/ONQYd6UmrvCSVO4+MnxN14pp7B0/dx78RBWSCAQ3V3YCoRbYGS//
f7zuOmsxtUcOF8+pcTmMwYdAgqIEeNvONvbgmRwWMw3frRx8V3+hxPxmosYmPgY5
lcH2iqEVDxKb2lIDydwieI9+r5oxM+TZ74LnjTAo9YP0wsFyJrnElu6LO+oy+sz2
iTksOSvaBooQ1An/yy3umRwCl2OUBMFt4DrFMM9PLMIt983a+Ej8FL8yJbpp7sq+
aelUk6BpW9Vjt8NEqsIqTb6WbHljgM6PYyxLueoK31+UcMdOt8+J16VhgEMVgfKQ
rSCEpq/143ckTAHxHSlAssmyB8Nl4LXyt1Zq7v7sPRMIDVc9Z4EPkm3qQxbH7LMi
qMSrb/mNneamedFhVNmbYphVcroOb/vJzqVvlefTTqGLkxKuUOnsKYFJCL2MDBCP
rAYn0aV8TMI6QH27imqjpvaIbYxwjDuJ9gqBYiKVAOIIEHpC09Hp2JGcsO5b0Mpr
h8gke2yJcLXzTdSYLCkR9TBHtrv1pSA9hV9kymKwD41xm5EG0VL8STfc1p0QuLjV
fOWNREhP+nVw1ifohIC/EwN5NSr/MjK3dJkCEVJPS6sjm+v7/ySw9y445FnlYXex
AqlHlmnm+WnviKGzY2nbi0kimttrbcExCCr5zbdOyPA2fmZW8wZbwQOHippXx3CY
hq3BiJlAYoHz+wfZ3ovFZlqh44dOgHf9AVNH21d9ucVnNaHKSHElRx150JU6gJ4X
OAlREphN2GrX+RqopCWTugFX6REdoz02qTRHu/jsnHzGnlpqyjPwAd3e3uq9Qpri
tclAt03LZcD1OICS3NGaeYbJyHutzGMOSkZ+XObjSfRpQupgM119nTa3vMwh9Qlo
QcQyPFnzDw+wR5JcCGCYs5qlGajrEH9A0uzOSG3M0YqoWV18iuuItnSSs61Z9hWi
i+Z6HHt8QjxkAFHaSVC5YemPyNJpc/ZBH0mjqJFxCD7ZmXxFA+TSFUWhEqXRGV/a
oYgZw56VmFxuxejs48vB9oq5H7I2vr4CMxPPUOpbnFjqZd7vzVdTl6iIJMzq+s4X
nKuktL8jfK5yiCkG7xRYO2SBy7WFHHU3OJW5alRLxvwVqe8cQvMSZcu0bTLKv1G2
QXaSJSbrtSBqzSfk2zWzWWoSZ4rGkx0vHhbs4HpH2xG5peOBkIyTJDpELEeA11Gz
6yADp7+1jifWurD7buEqhr0ZfxvaYiBZQzbytB76Ff6BfVqCJKTXTrpgrPIGn2mB
TfzpwAAYZXHjLy2tJ29q8N53Rc10hsWUP3McDRL7U7PfDCL7vLRc9x9luPUBYIaP
rlfqOzwR1ZkYbqaCgU45VHrbfL9EmQMk07wKzt4L8nIjnZ8CFbIAstVYGDeRW+1c
UZB0LRTkD34y9ilC8o8FG/+/kWr6zocZIo2Bz4wmQrx8OQIisgk7XrxoK3DgEuPT
gD52q42CcLLFKxDjGyYjeRjk+e1wLhY21qXBmbroPm7flwqZC4khRdrPGasPdyy0
pzDPzvZAKn8ZEnjjiVQ+QDZeKMvXiM1HRwPWZCMBTrBKHFdmZXj9oBxrwXkYokm9
kziwBjrVYpojoyZnxgYqldjTtGoIy8ZekdewtgL/JlTwnNtIxZ4iWPfp91FaXQen
TLpJ4IGwK46y/t7mblSlBTFUMKiubEo8UFk12Kp0W7gv5ssBFExR+ZaA/Rc0NDGk
7DbBpS2EVi/76GKHRwzhM4fAn77zQ2dQuWw5VKk1GxdUhG1Ve+xXsOrqvoaYyzuI
ZpsC3VxJRUAlVrpu+YzcudTBt9MGMktDx5qrWqAjXPVMFcfxQmQfidsGojHoAt9J
HxqbmF0dWx6U4uHuYp0uS778ZeKemtCCLraA7jV0uVN355SXQE3SQpkLVtam4rQu
FrtOrI69u7mf1tTpIL1wJ9/5fK/snUtbbJKQjLABxKusxgVq4NvGY+ZSGk286Vzh
qAcjet4CbOCO0ilATQRTEzSsjn4NYMY8ydENphK/o5KUW2rO9hg0OvDoEiR2MsM8
bLHgeGpRbQSBAvVTRn6BlV2c0Jn86P2e7zG+djJfsBpDIEfN6x6etGWb7IqQ4yD3
cy7p1Uj1y4wyCcdyScicBpSnRfaBAEFLx4D6cWLz4+lo8m8m+bxg4PFjpwJhID+L
bwiLo3TRdvWcd6PLZOYUOu83uYCBIWr5E0mbJLTbFFfPuKAAc78gLJpcTSKx+Ezm
6OYLM9VbVtG4kAxCAhzvwmAtCriEJ3/AR5dys2UvdJ+ubUZF+0UZtI1mydoG2M5P
Z5hybHuQDuRl1eXFjEH/Er5MPQbdPMzihqRJjruyufa8k5o3tyiAlN7AosISHwiJ
B/63oPRpuly5ciRAPEI248wy+2EY/ZDAvaUIoNfIjCnTKCuJb6RD4hsGyARleUrr
IbZKWvDygYkkBTZFuEq7+aZ4NjCsspOg5VErgq0j/ps1xKZsZKBqpxbS31rIXvCU
zvfePHI5NzeTaKvZQeP649Ed7aLHMlWxb95zrsyQWEAMEk8XQT2Sd4rTxnpDZ6rp
uB8PzUTP2Tn4lGAgJGQCcg2I5ARfumSs1jwBLqSM+5jQ1dVfzSXErjw+pBnRcWAV
iPjftIc36nAGKw1FYk5wobRyU/r7uxDxfezyP55jHay2SXUNBJC4UZ6QudGvFA/J
0CwFINwKlAkwVhYdMIpzCLWT4mLC1XDOQCfZIDkx1UPyvR5cpApfhpkVQZRTNMdz
soFVEMBLyQxeYFZVSV2mOsG8LoGVxHcaKMd7e9lZM0DaGJHd7y5P+0QzpgH9/zGS
y6Lb7W4SjqCh6dJHGLzOK5PvqvsaCaGnarFREkGQz/t4h8ppNZJ5SnUVtP/moqD6
hIZYxmgqEyUjxOkcXkCx30bjBmOQmoPMJwZM8wLi127LGYGMU+19y8/0yl+8IvRe
xHTt0rM+KltL3MDLAXfMI9Aa2+UZhf+cFQvVCrssF3hTreUVt34Sb8CUXAUx+LLJ
3sc1vwZ/jmaHPixdCcLy76EO5jChJq44XWcoXnJ8muaU0cxi/NLSDRZ3mUkEh2q+
ZnVDM5cWAFZW1F2k8mNPrsgJ28iIaZ1GQDYOvnT4j6pBqcdX/sm/UpM6rE5QcMX7
I7DQCz1o6/TnYoEtcDnK6KL2sIAkZNyC8UKu7U9szJpmg1b8Hjalbda0JjGrBTW0
fTZ2/+oWM6AV2aEUIdumZ/jnRfcQefa594FjN+EUfbde+LqxThPvsbKBBgGu+pMG
eb5NKNHdDD0XLUDHjB2IyK+xjETirD7S5wUgAEzbSt3sZ32Jb/CdUlp0PSzjjaPh
essoXE7yDiyhkx4UYOebePMwfvuS8CsA2oXskwObtzCvSGohfbmkU7QI/2PGaXy2
BFpB/jOoa8nOgOGQv87mYpqh1f3bGxKpPXDI+UbRYi10nOizo5tG3Dr9jUOeikGS
WzEDFvcov6wbffWTbld/gZN11FlR3nz/iKEt6HLv8tpnQ20SprTML2cg+mWplNZc
zdiP+KRoK0DDRqn3/cS1oTWNDPwsd5bys9vRJ7GopW/6KvWxZtL45EBkZeKtN08j
DB6jep/LYC2Uf1VFs2uu5485hdFylUXOUyrRmZ1LnVhUu8J9p0dHLq13vUZ4OsmU
2WeLs+lM/Xfv3UAXtU6gmhaOFP1mYDM+ZJey3q0JUdi0tCWONmOgRqGSfbdKA10m
vmpjEbfUw7r3IFL4Dvle+SZGqXv0tfK8pS00NwQ2XJuQ1jp/SoW7+u8f/RfnsH0M
lKRxNvYyotULv+8NZ8xdxRyzLI29a1TKRokw+dQsxIsfMiLu9Km5KYL2mI+0kv8p
70IEnH+3avoGmUyGKIJEW982/6nb6sObiPgQmyHVcOdCEcQ+WhHNwwB45p1wojuj
X7yK5tCIwi7882a9jMAlBAtLB4mxtZLrfxeusKlgEbMn06O1J0nglbeOV5AgpOEc
peruZb7wor7Ka/Lhdhnx5BN09oVQslTWnnXRod92JzW5h9zpjfLBf9AbK6lYLaVc
KfBlQpyocFFIXWb2P5CmHZTAKtg1VuyALtKSZZzGO+nRhSfXCd2HQNU91l4FDaB3
uaYLfurmNRBpBMOtK5QqzbR1O7LX1tMadZ33FApFgv/w0B9rCIbSZvG48OiWfDLl
JPFCfK34zSJq9as9N1fYR0Pkz6Wkeck+fecljZRXPt3ZZ+wZxRdKQdsa0mE7AzP/
y0+Xvf5s05zxY0pX1vitMtAU4LVM5BqqVaD0gzzOSyC7urHGNQK5vBRo4QBzXIT5
Q1DFXBWecX/3yduOiAv13VHx5vhE08EoqNbFBqYwOReCMnTmCkIxV7YeDLTN2g5r
/EadASH7a1T92q5ClV4k+LxsKybOplv+47hVXhomGwV6bo8wp5ljXP8PRgq1eOXo
f/vV5L7tSpe/8fdLsrldkuvHOI0Fb7JMTJfx7My9O+IuOcsR1lHXGqGxukF/7VSh
CWWJ+uMeWOcZPxBI4mh5AZRYvO/iz80KVaeYh8WNQb6/O4rTe3h9PK5I5tLGNaMs
l7wYEvx1adDR9VLQ2H6OERR2ieRImhAj3KSwpr+2g03cdcuLhj0dL6TktmOZ0hrX
gXzvmSBmsyiXdK95sfsloSHp1tRsC0uB5H/0wqxh1PhekI1RcxF2QNidI9fCznD6
E93jVH7kJb/KfPcZk9jOYlM8TkvUUCm5myhHbTMdeca9wCkKkF4QfCa3Nnk6S6qY
4GQIQI+LRUApTyL50IaLuPIK/VxDFPE0kV8CqMen2bmA4p+Wqp54rmR0Ss5roNnl
YFyHyPXyrJEk7MAXwLo4SwBk9b9U6nI9/MD5cBgpCcwgoFfuAkquFE0jTHBtr7iz
veotq60fJsNAlmCpFqKhUENQboR+xSEM/1YkB+fbCmUTodR29g1FVX989T+G37SG
VfzFHc6TamjnP1seKI6o3enAuLsHRACKKillkfrA5GKfnwNC9vKPeBDc27/yBrw6
SZqkIpB/pEpyj0eD6dLJ96JbIsbpPG7wxv1nn8nIExcIjQF5lTjQViI5tJSefo/5
9iqOBPqD5z3UxY4ipJqOLdRIyjcKpIOy4TObebiIkCEkXbaW0R81mHS7aBTDvzcB
Zzetp8MXj4renobPsZ9rUEgdIq1wttmt9kyLGphDRKmCMofiy+tcXn/VW9lkJd2Z
HdAfXSV07oR53wl+Z2iCqExnY/6kPywTJRTuO2hKDhpNgiRRPuU9P7H+Jt4GWk75
sPT/zJQaw/VFFqAOBL+BTeSNZQt+BmYnZQqcTSrN4kNvcd2meItRFGmdbgpMo1YE
UhK9gz+p0VxIr2yPc74QnKmJjUQEX1z8W/EuILScAUACWfsomXb12LNq5xnvsTlJ
r30uMiKou6SjSFJhum/pw6gPkJSlb/jbeCBZI1LXb3XAxsEQtLqd3uUNWNrX0a3U
urRN652NyDUuwQDPlUEebnEniYHxbIRzVW1i8cW4WwDb1eJOKeY50Y6JDkXl4/al
tlauZcO1Z77cLWbU2P6+12LMAL6LWdIi0/bwJIWKE93HxDcpaBPtFYtXbNhFXMsh
4lwFfZYMErj9KXIcDVIituCyVFRTtmlH9NtdjW78mf2N/x4LyGoCTiyAJeLUuJWp
5SDXtNVK8x6fSsZBTlIAU/ZIMGz4tCntDN/lbyJw7pFF/QWsDSMSXNWSUijVSbnj
0GV/dd4LPwC5pM4A2xBV6iEJnK6o6ZR/Qo41LMt+lcrwpHUy2tjMAXoknOMIw0Uy
1ohqmRvaN1NT9pRrQofUkmJqY+vf9JPjJdxTqrji61YTCIgzp46lFLh5FpsIoL74
mm5r0BDsb2W0cWpj07+gHAxs5fT3fp+1Ami4nZqbsouoZiNc/jh6ZmlwOZILdX66
kKmFcozE9PPR/ZXYfdWWbLxeaImX3lVBZq1ncUeCA9utZmJpL/cUNoC4C6/Gtxv2
Tu7kB96HUWZJgPkLBBSvi96vuMjfW5ULxgXZA9JKWtgks1hftpPETcuUCOMwf2jq
TVjeMeGzkUPaGLvzwITouhV3sslizCptal7dzrWu2ALiWGmR9oFXMCR9IGD355xy
SfuH7RDC7gpUwTUfI1wxKhp9QOazTTd8eGK3Wr6mh+b+WbjybUnDQ730ftLA3hlA
5FcFhNU6dRefWCzzd+qM0TuxEn5wa45j8gmNRtchkbkDkAwrdFXc5YbBbtkr5vgJ
bazOALR7rb8Nmgxt2gzYHjGqNT9/HipUTQ3LUGJGY4Rq9WRvatjzZXbcN4TLpHJu
qZK8o6XiOrGLBgnJB8NRQYtUkFF3PuMTimTVEkShDF43FL65PF9wWMHJkgBDBptu
wwKt+8g07GF5aOrS3sVt5M67kWDfkTUL4JCkFej+BjiCuGmYEwZWdP8tNmG7TmmN
Yvj8Jp/4eIHCcITPpQPrw+xtGYc8qZ7p9csO9q1ZamNvfQHs2iqiMbaTW/PcAfEB
u7UZK5QjzWUx8XjhrI1L5F7XoXO95o4sRskm9TvgmdZNN080hNvDZsMQ4y94OlWS
6ukF0XrHImiJpwSLCI65AV+hxViug18vgjLXyr5FHWrlj2NDIMB2fuA68Hqjtjid
/9YealHez9YO0yFuZsesJnBN9kumbKgEaHQILTwfHoV94dsavsMMZ9w9th8tOAJN
xMpoGIabDo1K+Pt+vWW4v8qd/XESKYlpcMdnAXKy8ifakBgAzuMtFeybvD9Bbd8y
XH4w3D6SffaeIZMcOSaiQDt1KF5yHJ+goODcoITnn5g3/KsDK+r1GVZkufkk/iXa
wQC6kKKQkdctl3ezHoBIF3ojZGIo/itT1yvMfNW1a8LOQz/bzqhhzBvN5mqeeXB9
vyo9o5f8VxlL2YVjTrHbVBfNTjAY6yAJWuLyB0vMXFX+vca7WiJW2X9qrAejgb2P
sGXjbhBsJTOduhZ+AdkviOVI+QKhz3x2nETxUHvJyzjDPMGsmarsJZpMEkLX/N4r
61oorSQVeHQ2gKrp+BXtt4ecmjZqp2IlB1jL0gRDOp16eWvcWDmkiX4Jmy45jBOn
l70A/yydmRkvVi5+gJUsvKVgQJnFCHznUrSTsBHKKEZvoTaOnpW6gYg0YRsUH/Il
7i9JyIX+rxqD11neJt90t3AXsXd2h36vjRllhjXqVF2G1+RBXmI1xs18awv+/x2C
pwC5sky8Uvvf37X5+DdXvlxxh12v8vq225uIro88U0kfHb58c/I9MuAVUMmgIng9
+7bh4gPuNfWaJ9qZGys1Q6bUpJnysxjZfJRcTvhlb1OdvPSn7unoUBW7dfo9CsJG
upK8wuzMoYIM/e22G4ftLolzSdbNFop+dANdoiRXBVTQy8jdfXs6gP4wbYbqHoXd
Fpu6IcZU/Cpy++MX8Bia95kDwJjukB6fZQjad7WG7FAJaBcP29XfjvFtFrO+64Qm
regBd4i/i5yb2z00YEnohYnD6VaESwwATOBJwXSM0tCqqNbv2nqRGc2G9iiS9a+v
J8t7HTL3t1WIsO6vQP0eIlMRz1PDnP91LGYO1pouCN+ZPBIEtBZdAsyZr4KAbcdV
7DIUkfqzNNpXOTnXQ8vv9CSu/Fbw3F+DyGNKn3p4zf+d5+Z+tqv1VyBQfvwghAZ4
gSSd9j40FJPnTfX6GqDvj0j7OW9LY1KjJNZ9Bu7VAHQPL/IODtOkZsM73ho6R6TG
sRWm8FjO+92PNWCpNBcxH7EOE2biVSXAkcKbZibVmjfraftr9Ku3LjmCwPJY1+LX
sl+vA1vMKOb37AArbS8h/A9bdASAOQ3q/ayRifv6C7IDL/ink87nG/ZQtHyZfpGS
wcI/Fwrn4Ja+eDcTYtBy2W03ZdYRMq7F025MEyeeHiJ9ws4Hm2oPyKhMgdcAHkms
gN135H58ki5/6+tUxHd+QYD6iSemL/l+8DKwlIeC2DEMxIWgweSUPhevEafvjnzR
LY6qdm+F8aN1H48mnUf7FBIAfJIo4eYbaFF2DIkaE5GNsDBQboug3FPyItKaFKJQ
BXO11B7PmJR1ZytIR5WGgmGZ+s3bKyH2zzmyDwonIBCLXUPasF7YqXRSGnxUj5QS
t3c5g6zia+uIczVyhebo+RVw+0DM7vZCMfistuzQ9iszA8c6Wo0zuSJSeSfvxCa0
SxcvRJyPce3KHEe5LrEN7Mz7EwJXXMbRyUFLrn63hUBpnkQWE0z9Bv7NQWTnObde
f3vbSwa2QbOal/As5PAO12Z8VPsrkpmeDsDc2GwbN1VtSWCPkGTP2rtpvtlaMRx3
76evmhufnKyELYXGfDgBVh712sL0iJ+QxwdZoyItGlD1rOKUXMNbSHD0b2Fi9NcQ
As8CWk8Xij4CDnE2PLW1qaPlbLXXUW2cgyJrhDv0nlQQUn1xMLq2LDfgNa4A5qU6
ZcM2p2EDccWtbMNtAcACE1p/8dwRTXsk5dtIiRVD667dvLXi5e5jLYBwC7WLn73e
YtPPwrmlApV7CEVMqNgr0XjLEDfrs6B1BJIywtRJMY1ZpIPKbHQZCReKelGLpBgH
Kira6OjjTtKd+icb+wqUT4+0aZZIme+1mc1nG4dvnbj4X7chmkfLty54gOuYJdEh
5z4Rsf+aXhM01VqibI+hqYkfJzrEKTQ8xgvux97tbJesayymONG7vW/AWPd0jSIz
OVRr/dx6K0XOk5v9O+xocCFdU4lLq/Ivr5m5UvJ95iNePuowy9GeTMTEFUPdV2UU
AzR+WSO4IAr5o6akmDuwz5ZW1T7jdji8cSj1Uzok4tcfa0q+M9eFhlxGnhri/bBC
MQgdUQy5iAbXmzm9A/TATMj6JzJCLE8y68oghN3rRjivKY8UKKw1L+4GEp5jrzxf
XLLkaNRYvZrC9SjsCZD60F9McnRDa9ohOWkwSns+W65r16pGygT8gsGsgb23IrXR
5S72Q9urR5+zONi8fDMriK049do+sXSAvXLwNl7T1xqhmdQzHFYDkKSzZT17NQJI
On8YKSfR6NQdRXjcnDIBqB7LJmjx3OEZEnaQmHvKTuFr0ruipDglHRv4QQgI9nWh
8wHP428E0mFzdN/8sWN3zlvXvX9nOWjqbXK3DhVwn2mm6Jvobwti+MgUjeympjEU
sNOKYuvPx0HOo/fk1rP6EdEOFFLqdtOA+n9qMLssebMuU28TcM9wVHpDpAQIN2l/
AYBpyG4TDZlhayhJJMiog7iOSL7zdLGPNjnK7J7/D7oju4NiOV7972l2c6IiQzvF
eJTKpq5LVcdEma3niPVpeX6+srN4kf1Al8m9bFlt6YlWzQIWo5WEAbis5fwS/0PV
WpspFmom1mfZzrepCJejZArgiPFjc5HDgu7a8hCRdmGwNTRIw3JWhup6Qf0nzi16
pKrf/FPvGeAx0zvfkYQcat1DxU4I9sksTHKvYaVkzljCoXkvQzksh9Q2tWIrDpX9
YHfj6g3U8cXyglvrbi/JhHawTon6L6DbWt5zcOzyKIz/m+XAzsFzhoOOI2JbP4T6
NwbhpHoa8qd1qov2A6Acr1FDfG/Hlf0jjpywViYk0NufvMEh1T0d/cVDovNsQaTW
9B1XQxb7VAN/4glaHAf4YKCfh6keN0E8vYx4cGkIw57MmREywFUbvIZ3QlNEzMEs
0TpuGoHB5MIavq8NAaIx84l8B7Z+lppRTrzns/vgzkps1BemT9qwPgxuRwYfSwy6
IQL6CD55LHP+P8zF3nDdURzA2mUM2vYYKHstnjaomf63deyp4wmV5+v683LWS9Q9
3JyoznOcu2rvkoqpx3DSS/l6KuEe+D2cSmgTyvBdiwP7WOtskh0SzrJJsB0YMhsm
3w32dYhP+AMoULqEfxTmR6iinFrgdz7fYDBfzXTXV53d/rFftC44mARuiW65RV0y
SLKG3OTVQOa6pvY3M+qnXq6HUMLNZPUzLo0VbYOWSj3WiPXpKT0JLynSNeJzdftF
sIMnk2aRYBlkS7b2H4KUdsVL4s0toa0LnU4kqsRxGkkoXqAFTvTk4A3+ICcQay8i
jcyOYhybXSc9rbmbc5NKeSX19czPV1flOzTh85HWWM5FfjdhdlQCGAHLSPm3U2+y
2Yj9iMcC8GIaTSc6IyyWHWqXHkdNSGQWuUZIi05XNtryHXxNKx1P3bflz1b00ACn
EfXD5A4nASDBGmg+dMh1ASEjWQLKQsHLX5VpOJ1ojAODmpQv5VEHmI1HsWc28je/
aun5VuSqTZzwVxU5gi5mBNaggCVhi5WfzrplO9dprOxeOL+8HJXGZjTvSwmy66UM
U5/adMR0aaKdH1q4m/CSOg8weovF9uTAZyTdzD6nJQV3tqJE1CwM21E+pm+JIexu
UWKPNqJfcfpPLyWauE7fcFqOx19Lv4JelP4540/OYA3aMcmgEh1p1/fj7TDII+lq
Nj8+HJGPtAFo2vLMm3bwbNzkjYdxUNvikxZkWrwx5lkNpm8g0VbX1LJ0NAua1oa3
VN8SF435fHTeBsGy+HzgBRhFaYZF+LN2dy0RIkMaD34FbXXn6xr38qMKnCDFKWrB
QXxwjdroYx8ZUT/gQc4CZaplSEfW5atkLk0Ob8fTo6ZNIlvjr2WumGsnKSaevyCP
Im8rql5X3Rh3JvRl2nKXQe1olviagc8k0GZ0HkYNZAGJIy37wLH88StFR+yoJDOk
8HAxa7AgZKsW9w7fJcLYYllA8URjjym21WnLpEg7H0ZC7pMEL6lqqcviQe7OPlIU
wdSxi6T2ozS92ZpxmhZpzKhDNoPex2WdH+wiV/2d2alwdN5IUkazsJEtjsWCyd+E
bb/PxEsALwKZdvN3VP0WOlVLb34uShkwH80UX2G+qT42sGH6Q+6PxBjIJE3eHalo
3QpVLLLcxAtgKBDfluR/sU80hfjH/eeNutOC4fziUs6MOc6cE7O6fpCA9GmQeTyH
OWic1Zo6KXuaezObxK3jrZ67N9qnTB0A1P85skVjLAB3tc3mCpw+uo2TYp39rX3j
FhIAfR03yY0hZFESc0DATDyonzDLpTn9UcxOJRkbgHuJ7pu7NnmA0KY4WGhYdiaM
6MMsxIUaO3qjyjOgPPjL2evfdHv+FkEN46lRBVLjh4OxZ+7MRFvTMCzsLKRwH6Yw
Sst5PXq+OrsD2WKyZ6k+VPJe4XaYI3DnMSGH+M8VSDz7CMHyeloZ6zmPJ0ahljv5
xURWlqwXrswDdxUH2VqSbtm4Ni7mAlNleMIBrR/wvL+mmbKHq2jh67ln82DfCk9M
zYjvcPahzDMWsu8acDzQ4ect1mih5SAzjONobTeYgARmRAs3c7fWjuBruYKpaIgG
D+lOhDLUO5383hbn+ekB+scMNE31glgp0WAFCWcDrSuSzUOEdjoFqKMFJB0vUq/N
ZxgW2w8I3EW1cz+LVhRtkZXraapoXQyPwXUQcqspNh1ZJ1yKtIW7EU055995udXP
8uPn/OcVewhNS8Zacc0zJRqQ4ZWi5fdRjbAYEuPQxWhBNPuhgsPmqc+1DG72PtRL
AF3Rjyv3wEm+t07qDfwqiCVEyXHijz5M9v0IuGiCYVAi3bAhqDVyKtFAFHRTZIUT
1vEDaKyPfhEnFDg0SnEdw6vja7sAoufNE9XPKr+cR5QqmNXIwtVDOJaVhN5AT3rm
6OJYa0BsD+V/90WcPqdG0On8lAYxFSxNdld29vubOUsBDwWlTTbHhPKa5F3ZQ9lt
vsAHeDQ/Db/nKKgT8SADuJKIv4IGzMuBdKY7aKecKj8S4YT2C0FapDQc7P0jWroI
8vnBZMc86r56NTyyAdNUPnm051YPNjLpQl0rlfUSTkmqQ0bJ6b2Tkev64KN98nZ4
9Z7kbS0kr2oAsU29XySwhL8GCwiJhZKKGTD+qKgw08M++fTdUwsaY9r4lGdTqTRI
pR4ytGOEa+5P3WckwvU4E6Yb1T2F6InlRkvwT7lCVr8Ntjguoz1pXwrolD0CnX6c
qDISZuKvRd1Yi2JKkyIQj5fFXhNQhOLbbZyj70SOfCsBy1IHQO1w3dHMPdOUld8z
V1V8pypSY3Nx7TA9R8KXVEdzYC2D+28v6PyGUoIs5ra1C7rllCDAnUXDytvWGkBw
do9WUXlOLN7Yqy9BJZe9Yj+p/MYhYQlHjMsBSAf15n/8/CByx1+w1WdaJD8vrWpU
hA9nOqbwbf0Dgn/MyVVgw3SHaSP2+ZLY5deboifseOdqzQOdFfFj5iHG1f6q1HlJ
TlSU3xRtgQnF9MRpO3iF42hN+avQX2xdT0QFOu8Gy6zIXxH47w+MVDqWobgAnr4X
rINrNujZxj5Saw2vjneFakNNczCo18HLLxUYM+IYR9nTznF36zsNrzZwYCImIVH3
ku+mMBPP5mmIJEeKY12qW6AloRvOuuOClm86Gqlcar2yi3MCnx3qmH/fVybgddrL
qMQKOiiccjEZkKnQ4Dhr9o71FLgE6TrzrBkxA5zHzTKMiRI5Mxuxmi9XKNnTh3aM
rblP2CEVoX6rC7fElFfQ00OaIykZ3ExvoSN+WOfW4qIHHl+cxZhNqf9px/us6xAK
+hLEBXEKdUtiaxUqtHdj+kZQ9+cHFfG+hp0Ir03SI+F6rURBsgg43A6IOoCMHZZx
dpVxjDsTwmuNKq6dHXkbLP0l2rcTjOu3gnQvj1OV6JAJNl1cSf+t9f7scn2O/RXZ
EZDT3Gigb97CThHbykeV61maJlb+RdIuWuEDmMHqzoFfZobdj9+UtiB2u2cT2d0L
aguX75JRM/X/weel0oQzYKoxP9p4DbxBB6q9Nn2gaM6R2Qi6F6iHkglhr2QZNhwC
Qc34NcoADRwE5kYYM+nqkd0naU0wWkYLg41lep+7u0zzueCdR7OjkfI56JcBMMam
nROUl+kpElI5DhPmV2KSUbZcNjByhIE9tvBEzqQ2m0Mcg8QX3/Ui5sWRGFSiu/Py
oLf7IXRvSsV66WOUGsWtao+gXITttXx6CgvRFjmZqItoiw5bKCFyK/wV4C5+nw70
vqMoliYGVim5UNQgiiewc5TQkUj+80goyE+AVx14Cxi2bGX4V3IKynf0Kef4Ywu0
BQyHFRUs+/76UXhNlHjeX9iJx/1+1xz6+BH64QnoMYooQZRu+9QP/BhotAoRxRp1
tpIdvw52ARThOKQdoqzGiNP8oWQN2XM6kDBgP9BnS1nhLvMcXeNlSEL86JWMiRZT
c8AXONSln+C2hcSicEITqbogrNKIDvLuRWg/AYK6kwxt/tRwKEzhPmLs6uhMwayE
eTZp6Qqd6n40W97RuUkHDRWmsJOnU9iQp2KVkACI85Ngd8yGexNL+SwMmxRO9daN
a/LUUalRxaqG71lhksA/GfRlacQB9ga+ImaC97lPdE+UJi+9u5BIcujMSjc66mT4
SWiQFzWeaW8NGIiuodiHZqikeeFLrUjTTHY2FaJEAChMOqyafxx4gbZfIh3y9lZP
xmGHw2QvUbrjESfbYzaVuuDqvkoS48IMVEvfI0RzWZcivDkztLPHQ4QvOxQwIRNF
gD4fDbZSSmwpbKOlmg7gGd8QTEQwOngyy+tWVxdeaC6Z3MX/snI4UNU3WlIsNUxs
LP2DiEaGymDC7Ay1rKlOoY8rMZDUzvb+0H1L86mfp793hVKATHUBDGL09xmMrLhQ
NyPJ/ZHKTeXokojzOdT9R6cF2qeSeB7TxZpzMrSwMOeTDmpyUHYckvstkoHF333g
gbdC+WCwVW8IcJNFNPcFrD+gafM6smHTIRw1IBLXcB/o4UVgCuMQJWbvhRPkljlq
1f6FxKK2nYGTD5/+146yLaBo5uTKNEAyAb30MYbpHouSsLoRAiNzAw37OyRQZZfv
mp3jqa2lkWfbyuWBGLDlEb12VsMOULMR2dJTpxCdSuR1ZTb3o8TRQMWw/whz3IdO
NGF0EIdVz45Z6pW2sYjf0TLtA9NbxcBTLhgOe41FtKcGs6Pheqv08Jx9T6sWdIuy
2ggXKzfr8VlavtGKFFzGvRCnssqhx1nTC2djX/jHyJ6Buo57QbRoY7wz4VNo2HfZ
autuJ6k1YOIfxqOK5tdXYQU2eKZiVnL8YRCIWl8OPcso2RrYQZH6apLeZmk4bzSO
sni8FNg2rwsUuj1qvrIKNW/6OjecvNpNTJNRy3RiD4FUog0i1lK9vLRxJm1rl3LJ
LMV9sTNUrUphBuqnoZOmNw05k/d9yLaQW7Tegk7wWxMaIV8yEt2jPUzEXQ6RWhxD
oC7p56E4O6otA94+jp8RXXhw0F2NLBPdzKCRzPqNsUMPCuYEzDrlKeC5HScMRcz+
/EXGVUJxMZmm3BsnA1uHMXUUUKnrKCHW2NBkNFI7wKZNWDDrI+d8ecmpTu52rudV
FsprVhLQCG+Yj9nRGz1aoDsbf7Wp4TUBkdny8/ONAQLTq9Z0whueXikrlJ8aN+IL
4SCUo1vv826QzuWoYcvzLptEOPeubuW2/iVKQUNIL2X155BZKCBjx2hVw3XIAnxA
85/lvv0Y7jFwAWJx7ZhuS4BoH16nDE3MJ9hvQE25uwCW4C4nB84FBQ+GcxIWDwBA
lY7k5+UbKTYg8L68wXkyW6MUozGNxQLVQiLLYfiETcFXf7qDSIJ8MH7b2lKtcQhD
`protect END_PROTECTED
