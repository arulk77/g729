`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
7lGEhjLAsNjjFc/QLdH1Cogw+5MP9n8kkGjkRT9PZV5ygsB1ikugauiIC9cDecc3
OeDrukuqnJEMDSpSkmdBPwmcJxujsZeESTlTDA72rHl1uATdjmKUuUnlSKBnnWJ0
qmBxRe9UG9ZNck+H3QBjBL3CtSZtFHvYZrFiYFcRwfMh4fFbO7Q53vixF/G7lKRt
`protect END_PROTECTED
