`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wKm9+9PAFunYx31WcS7sQj0l7ns++NwHm29S5qdlYtM
ZB3rq92q33qmR8+b0pvjVCgLS7C19LP66adwFECpY8mz/EfgCcVLDLMNk/hh4UpH
MmY914JHFImKp4IdyBpmRB8mU/H6qE84raMuz7QuDbuV/QWVAJnSgSc8ylkA07z7
AcWaE4aS9IZMLBSq1GLpOfGJYYs3YljxDJdyMQTBBmAqMbOMSgpEkM08kU2PpsAv
o7kKceBnxjIcVcxLWTPaoLfYowsDhygl5cUfSg+vkwKVnTWLcn4+q0nP1dxCanoG
Z/cUjXLLbmOS+RH9YKoNCmj4XvOCL8hhK65D0MzbHh1mpFT85VHayPjuzDGUQwUO
xK2FEGW6EExczwhQUOYCi25I0v1pHRHJ8+EcMTIzqubGgk88Oc9kZxM7sBQOv56V
pqqEPWLGQkNsYO/9Rf2u3dSbu/yrO6WzY1yor7qKnw9jQzB9Zxyaw2K0OVQ1JX47
`protect END_PROTECTED
