`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNa3gmiQGMurtxWZd56Z/irfNX7Z/U4m2bgVqsfOWZL0
kFcVrj8h8/vP1gHdlJTpPSJwU/RqX1NvWQvAvBwJGnHOhm2zpEYHA4XdBMBKxC1h
smkbgrBM9wD6//prSDKIs5enIJewHlHf+dgI7L+aGOQ14EFCAYBV0WTOcqQ5N6Gh
/EbeKsH0MLkCFZmUm3tuvHmgdVk3MLPTsnoyvCTzY5tiIhHL3X0LICrw+P4WgRfa
d3i/S/5T99PfpUghaAvOCI6sb7zh1BTralGuB49ZQ3N5oO2zBmZ447Db0nVCzTnM
rgWjWd6ap5OI7+dXV237/Q==
`protect END_PROTECTED
