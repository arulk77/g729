`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
WiuRYEYfH9iWb5h4iAI1sDUelwm1xFQZ2NwdbYGkayfqrjztwKa4rXqQXN6yOaXl
/rUHCFl/pnICUe6aB0tTSxAbXYmqhM6e6Ntrl58qDGPhXHbAjNjGlgQOZ7N29VrK
cMiRV4/JyPQCFrlwfEeC4VVYsapQ2qNbnZkEBdaz8NWEWrX2FcE6ocT9KutGoNdv
DofH4wGY96VGDKZ/TjXWdGwDr2qDQG5eF/805chdLeqxy4E/J/Q+lDxi7lAszSBb
8LnETSpzQhslPmiSu/f3xQ18GUx8HJx6X4e8r7UCQVCdwo47v44YWf0LSKlCGBwy
kueJjTFHzx4tbhU2StjCus14mz9moTcCatLRV8zYbvhHskgRX9FFgicZU7LQ8Tcs
6QUNciQa8kszNOWf+HiCNVgAmUiqb7VuSdZd+5nEmG4SNyn3eq3uToyiYWmCm2hs
CjBsH559JZiXYfXaueZAaJIs+xehpNMRHifKlzWqyEQ68JGOqGCQvfKblLVE2zU+
dBGx9EhEgFqD/1chq2VESb+zvsAbc7dzkQTQQ+MiQLDwy4GDhNvFAlbd9mdv9hOI
AJMkmdqkFheCPl2r7ELzdAq4+6mWXsd8gV2Z2Y+j3sKV0uqp7BPxS3Chr6Zsolhb
Hs80/rDCKRbPatqMon5igw==
`protect END_PROTECTED
