`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
37RQhHNi4JDXEBrfcfibbIIFKXJsoK41gkFdneU0vaBe1J+OZBJgewnbAVcmnUO1
sE3zAx8M2NV3APP9eSnQPtYPG7WxBO63fVAYeZ4wJyBpU7po6Xys96UFTDmy35+l
1WtokBicvgRFjXnA7rB7C449+HcOU47fU8TrpPJ1xQA0diq76u/iKN3te2bAGznf
E6VLq08cGNAUefJzBiwTklDPj9i7hgCQP1Od0QTwFDuwR/GnM6/89LGXg194wUmN
eT5NtCvdysNxYyJweoa3NNM/G40SxGyIECQlEy+nrvt/3eF09KYr+mxb48Y4VdBt
vd8OE1taF+A1QDc2RByYRDWO8l86Q8uN70I2e93DBeABJu1dgZZfcrjsLzK7ysYC
tMbh8r5s481y8pzofYNOw6a31SqI7KUcZFy3Nzg2qDHDjHt6clWEgqziJ7y7qYRb
k+/ftxqI1OZGSHaJvOi1JoeQJIEKyfozzxLWZeZ8Stdy1PFmFpmpizx4D4bbc/aw
R1xHhE9oGbGLajAZEqVihzgNLMxMwd2KAjrzNwkAU5wiQB7tSg1NJUx9o1Hy7QHJ
iZ9qWx/tvCAqFhzwrHZFJw==
`protect END_PROTECTED
