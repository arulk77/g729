`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
NBI+FEyqb2xGNT+rpfQNUhBszhX0dw6ErwCYaZYvHeq8cw858njXEJidpvB4bb1N
R2jOWALR+LHRtR5HcSP9E9iVb/13b+1u26xgAld39rJey5Z/P7zQC3lp5KEOM2Ha
h4VF8i7HkR2HvWPXPlAtzxnBK3aPyz5IHwi+fZ6NoHsqy0GFcuZmHwMcRPtmRU2O
taj2xSRzh14asyvkdUCqYoF0GPH6gEKlHvHpbElfQirjTZAq1eFMEuiwI0ZqD7S1
p2sTUpJyOjSk7q0S2zWKWptvkuNDdKwxs1IHaIL2i1aEsFgoM9JofyLs31XYQ3rU
m01eYxP/PfGz8nNllO+nj6NsuOJsGBZThsnVlr+yOLsLS50h40sg4fJoO6IqNV/e
+IQc/sp6TMMwWHWRtplPgzHt1DPm2eLnlwwfEuNv0M4n+jhzw6ZGZXnHkRGm2SZg
yf6PUu/+DXcdSqWO5zvPFw==
`protect END_PROTECTED
