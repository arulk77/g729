`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePB0PkEbH7wyjUH1VUvwroiLYPOCDimuwpDeSKRPdsN1
Inbxfj8Ttt86jfX8MKJPYDDiL4es0BWeWdfbO/UzLgof6yBYlhhoRqhtlq0FEuaf
F05IaAKaeXso3s9zBSHBe0S+mMJOtH5TZjz+yWGRXstc+t+rRWcQUkfId6sPIVp8
QnBOwKNDGs0VRayHbObOyS6yElIk1ZYsp3c151lgN/2z6d6/zFwCz9W405IX/ete
`protect END_PROTECTED
