`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
AvAh5vKZHQ5geOwcJmbRCupZw4iAnJgtb8Ps1AVLKaHGQvYd6I6V7zTqwAC4MC4t
KYh3avnQNEr5ycbjknfOfx5M5MjtKuVSL0QGG6Lv+f2Mx9blXUmJijj1IrrgBSUr
rxRxn2cERP49wItioJLIjggr6gjCFsrhF6iOnayGbykl7G9fd2j8E9xN9R8fghkY
6KksVk5e7wuIlNoWWFfB8ZQXAQR5sc54IBgi9aXKAcJo53y/uZfBasbYozzSCBnY
61gHxou2nABZCTr9aQ4exxfa9PHqIo2T4Ctk1rIhiRXF0CFTsMYxjBMuS4/skGgq
52HrNJs8BXdM46755AxvPSINoSNNWYTFqBVwPjYf5Ifs6hCYkkNgAYwNXwDwWO0i
nKQv6K+2utkR5jGnRBKQe4mp2GyRoaQPjfLwEpG11rC6JrJXob2ZVLQIrmci0jpm
lnYgdxxK66evSNU9Z0N9zw==
`protect END_PROTECTED
