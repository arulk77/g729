`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePrSx7aWZWflLKGmEjEiyki4hwVEgv4hJdPYul8GZwz9
nX/Da8CRfvIuJzQnTkfdbqUFucECUENaUrv5rqEn1RaYJhb9lRVuaVtjuhQw1XVg
E4HUuv8rqwFRgK/+atEQIPI+AddKJ48cScr0gGamfCtot5wGEpnN+FHArIf2RI41
`protect END_PROTECTED
