`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNwvqtLYvwLNkro3KSzLOqETdF/wCIkfpJI0T+O9dLIx
uvNCaFLwarlB60ianljMkLzw/75XoG72TpKhWqNXFjCZINoXR8ENeq3/jP1O5/Ju
WhCVzrNqVdJX87BUgriEnsLKGou0hwXeXBx/Slo/HBGt0B2WbdUxK4XWEowCUOqK
t6X9PCrrk0+nY8qiQQRhEw==
`protect END_PROTECTED
