`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SWsnmnYhpmjsBqqLIYmA3MsqGaV9K2qfm78uuXaWqB3B
o8Sg83WReN8CA7ZQfbHh/kaSujIjlVs80E05WEVpGOy0E7SZ0PyPAp1hKoL/zxcd
ZIk8CS7MQDyyTdqwhUlWE932TWpek6NxWCL0YsigLIr7pq/HVudoAQfiLIyRfmfJ
oSOxYAvc0iCLwmdbLcpET8o0wC07ATNn+t4pMLh/+AaWBm9NSOIlOsVXqnITYuEt
dQh69hbmD1OAmjnrsnzsGKWMsOOrqam9FliIGsKnbtUXgBn+L+RZ8174yTARByoT
TBxNzD599JJVNpSePJXkaMYvp7Dp50zjG+I6ped3R9ucDCo6/GbHKTM2+KhvVUV4
rBVhaq0nVI0Mn3X5GDMHU87BKH72B1Xs3AlAspmbLfG2c+ayVYG8syxIcAsHu95F
tqEUzwbWukpxcSCdhqYIxY/AAOYJvPVW/oj4CcBobvLfcV4fTjUYNTNrLmdfvDTQ
jBtQzvwoBqlYlcXPAwl3HVyd/+SzWknAlFR3oR0aZ/Zw6mIJxVUYlRfS0Pi+rNyt
VaW6SHfs8FGsEAnzbFTNuPwuaJolsgtgDdpDEm9UDB9hQQ+NS/dRQyHimSLjEPCu
0srZ4iEVrafJxGVhiZyG2Qg9eikRWMXzW7Zhg9FEweUB8X8DC9aJsTE8ThSlVy46
FNoQa/SdQfUL2SH6j6JmozNlseIOjqfX4Ry32+cX8OargT8B015MQqzpTOLbyqyF
NTkHDXUePMKsOzzr2h24nmY+bPgH9fUsGZoxSLiyFHspiLBZ1PE10lfeZQrJDghY
IASeTrO94P3EokMYllBarE61UwLNzONbSG/F8D4UthVGKFGEiDKqivUZiE5KLKPf
6Rx2Y4N/hNXHNiQEsOsxM4vW2sNTuSfYLsYKWCXMLMs2abqNa7CzQvUIn5LtzwYE
OTRgKlmmfbOUvhJ9MHQcCKM8fqmVAy7GC9o6yCpmz0EpBu2m9SuPp7O+7wEZhI8i
o2dxMjBU02u2HXCDU0V0WoL2i+8ZG14p/i8G8CAru/Sqym2g4jp3yMy4QYOqkU3c
byVWKLEQiyqAQ/ZnvD0DQyvUUY+Nk9fOY+/GrNgrZtuDgF26G4C3UEORE4Za2KeG
kkvrOE+5UCxjsuJTxi9eisjVIuyonymiQWO9yELczviHaGsNNM60ppX1t62QRK/n
LMA7lDRZevG6baNFwRg/P6MQGKeQbgQ0tCmZ3JXzprFpZc+l6RRo4eKO6tQ6N9cs
9Z9vV93UMSQPiUQdVgWkJ+m0X46LsvcbkVVGCadcAgqglwowwfViNWPBD3LDecjN
RjU5FvEpsCMabeCcW7mcpHA913yx4nEdiFU9pPlmsO5x5ZwekIQYJBxoOmP2DNR2
kieHQnmG1+SpwSYjq4ocNojsX0zM4Prcde0pHpz7VIR7mB5JTmIXY5dxAHZVTjJm
FE9mXCDzpMU5R78WDyIkhKbRpcRACRwOa5AyCZU/SdLuwHDPL5LnfzmWkEwj0Mt8
CPoTMoTfUHFwBYvnnm1FEnZxFGXl09qfGh2tX+K0lKabpmruuAe30iCcf17fuTaK
RPQjIXRI3XWGEtRVp5Bz0ZwdXqboqBbPc26tYnLRamrgWsvwkv/Kclvy/gc5TzL/
gSLi3lhqAXPgT1SfxQX43LnmBQigIwlpcvYfuyIWO1pzrFFdAu5tOFbr5CjbEa1/
ZJU3AOm4HcVLydyL+dXorDvF1mfsubHZpIcAg3aJkvXA5GuEXvy1gEGf0mVJh469
c8BFYv9E78EdkHIMTbqfBbwu5pIIoN/8hOSLqFexGk1LN41tGtm141jr1FTJysGE
p/BwfpijxHxBZgs88b89H43P7n3wWubTZGX3Zf88A4S8velvUzwHIJr26kkx1+y/
S/K+pd6GBF9FtAou09nVrNsBCiqMhVSjjRWI2WnduLCipF012JQsIkR9AP0JdW4n
bRYcSSXycnQyLSciptuJSiHVBmmodSibAbJ1OydcK0WfFl2M7jh74Lizsm8lmSlx
q7aquTPOiHQs53TeIjeQrOxte+6+PARSGRb/kW14/W/08bN2ty4TFT602wIo3flr
LLY3qzydccAIMJ798Ads4OUn0MUQpuPSBbiPDtEiEfkD8IzcVW9IchDzmo4akQHY
+30HwCnTJSNWumj1CtESLtqnWHwTc0BRQHN1vLSLRH75rMTYLi5vesdjI/CaRlJ6
wRrvls7d0DqPL4y1EJj43n4Vg8YDNBDGaIsASzscjn+B6zI6LoF3AwY3s+DXTI0R
FaZK6xxqKiyTreMj0TXgsImN88m+p4s26xe6gUB+Ybk9oQfYbasJUQNW72FOVLeq
jyvLKSo92Xrf+u9EEwcGcJ9Hirhmm46uCkBgTCbDcAlMD9ty2+5hbZ0zJuj8MWjJ
Yi//QqOYnfVBQH+bLI5IP2Gzo6pt+ziScCVCkzJ56LOIXe6w8zTt0Voza2LRvUpX
ItbGM6ZNSKdzzF166M/EhjWX0KDr7mvK0HAFSCKpUBno5kgZ6FQwX2fV1pPA1v9m
YpSY8bEXYYNrcud92aLlZDXJWWONs7RKyzo/V6WDRgs78+VO+5xVEJiLQfjVK5ub
294hm8lYUO5C+fIvoReSuOTZc40s7OxcvYMsfstkCHkbw79wznyiyath0OjGs+ws
oVMOH+Au3k8gx7QzoKvpHkFUypK5t459CZUegcD0Xgj24z0eI1aoUWxuzuqMZErX
SkciB8/YkaRz+NR+oOFIIggymtljCyBYicN5J6e1w4QFITRO/hpQsGMZL09x3lEv
EAJoslmcuQdNpo71Vl5b2JX/UuiZa/LEJ+h/j3lr7b8xwKATc2frtrhKWpGP+115
1Ie2DsTjBxS9ezQ1jQsnNhv4xtTJooPAqnFfclFP6n2vF0zW+vrQZJRJrX+dmrfB
RK0hZH+ehl5zdgeC+amuEbwroyoUH2+TISwdhvPEjD2yx+BeEv0KnpC73Xmw/O/R
Gm4n4deoAThDg9YcxiR32/IIjUPV09XNFGhcmyUBTizE9+V4v+5AXU6o2Vu5OEEe
HVFPreevSU+0/ELYLh1Xsk+vuAU889OFUcaLT5Ch4ticBXhMxN6A6ncv8VzOf4YT
hPRoWCe7vWP6LjXktxwRyybBfLQO2lsv6SsIjnIEeoCV2WI7zQJybTwAtoBs2fpt
WxcSm/Ytt6ccZD6Mr0rmN3M2PApciesc45db8luVRge0J6PXp+h5dU3xC+wsnKce
JV9gur//VCukVHlXZfQefL8FKimjrYWndhX5tfeYYYiwo9dmh7r6awFxnAZbFWwA
8INuDTJBmrWCU0rxqURafwFW8UPRZOPiMhy/Yv91TN+dva4NO/NQNF6dHAyyNodJ
X83EXL5l+56zpPuf/f8MX/M5uF83siMzzsmbhqNPrPvdxI9kgNdtoLbygX0fBfLE
PIfv5mjYhVzYDkhUFbUYm442GhHi4O2R97XX+OUxclZuzA03ytjr/hwGjVzE1+rw
/A5GPI17TGHhzv6wlsSdmM3+iwiiluZtH9npFOQFUDEK9BJv9pL/EWq4rmFyiQ6i
aWXEQQzVJNAIzy4Tc+IxJSYnqmbV4V/EXo0vkkb12E3AxPONlBo/7BFSb7tS1rlG
VPu9hb8cWGAJ9XYrcCqhB9wMi42sILcWOvLW6nG+OQGzmtujV6eiSvtvQyvyNTSq
yLN0Z9t4HYhbJl5uUiNVRe2JnBhGXMSjOdjDlBY2mepfDEsg1ZQhmjG2SjWXbcFY
OpSrrmoPQbU8mZiRMigOJwTdH3vf4r5lhyYbaM7VIbb9jF5qudkIi/WaM50gs39D
ZmlKWqOk7j28QMwxeBEGXC+QUbfGgM3t9JwxfwBh68oRkoEoG9K9KTKhv6sI/SsR
njiHSaPWBodEIeo1c+CoVKQXq7IyiK0JMHRBVnHoiO6doFR+520ZbJiv7+R02ECZ
oOS2aV6bryT4bLC0TuWcypDEIbuATu8FpWZ2jloYU5VoktFiX0LTwr88V6uA62EZ
PPzOJHujhxy8XSLB3lz3sblnxzWvcKYsu3VeaVR4FI4Q7szYCuawH5X30/l78IHQ
krUD75FT9Wokstu4TTAKn+o3u25dhKdfw3kMeYthREprgEpxMB7YMDzK3bZnDI/A
/I0ADB2CptHs0c8PZwrbVsWZeyWCTJUGGdCdYuSUBlimoIkPuz8RhhTc50DK7PpK
jDeadOBBYmy5U3FeMZSsheE/67OSZdZegiAFOLU9q8kCy8gIe56hRUokxNNcMZhV
BZ8OSwdO5OISboD3vvpPOqPoSTvxnHLOjGXndQ0doPR3PFH/7WbHDGRAyg2tSDT0
K/bRs3o87eHQ01ARp/QHSIwyKFfPGXdUPPhmCRM/D/qT8Qp7ovhIaPqqfgXKivSp
J0ZoxkUDgkE33qxTTJHo3Nn3HJqnyijz0wmgomPxfD9CGUcGefTnLN/EV43IyeX0
xmQxFCwOIdtG9nB/FcLyvNUZTNZCXECPW9srTm7kE4X33ceQo4OVgUfK1n1QMCtk
AY9f7U3i3M1Q+TKtRuqIKTUiYyKIii8OFrMfpb35G8q5dAwlJKRcsKv8g+T3Xhig
KzRyGr96cKKsIiU/N+dF18OVsgK6WQ5rTDujBE8GgMiaG4dR42+s5lvTY/DMt2XE
sYYZ3JNursIm/jYOHZ72h57L1eD2DISqCdYwciD7LdcVewYC4UzgQubePHx7wzMP
VrFzQ+xyTk7oz/6RPtDbUmRomDi43rMo/mHJt62RXIgLDe+AZeKWpCONtC3Nnzv/
0SGHTcqBF6B0BxLislZQzK34QOiS7i0R9tc4tlbuwlhwndUfCc7MqKMzE2H77PQi
uY78frWbtl1fBtk3IkNla6DKk4SdR3u0tEcEC0+nRnXuTNGKlOl44pmcV9J5LXl1
ChdiAAl2l1X1pTg9YjFzpAe5QJK1mAFz62wBVnO0ngCcHxMPvkmflAMmNVF93pWd
TB5P8EY3cdr3l2iNQ/2hjGoCxnYxZJPW2qkw0mLQq3+4SZadPeGD+2jHmvszaaou
sLqd5YF++AVk0a8DMUQIW1QWmOlEvXQpOICLBaFnoWUJ5JW57znCnyTTHGlLLIik
Bz2l8ge1c8dxE++8ND0B0knugvEY3mdeAbdpgmH9kyTCV2nYyZ7bTuPeZn9f/bIw
48iDcbONHknvkSqewl0ZY3Shjp0CdAPj02VvUUBZT9ws9Ao09rQWygRwI3X9t6qt
LKMVoG2q58Bi7hZU6FWnGIsJT62wUgyrftxm1Jgqh6QlgLY7oFOohaXCuPbg2peG
aOSdJzjbgTPFqP7UcHRyAe6+Bbf48eTrzeylBv45nLBad+k1BbMScgHcfrHmzS92
`protect END_PROTECTED
