`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOpmX0N5i0kH78i3PsokOA242qkVZ0AE7BunOb1zgSEg
MeOe1ELhoyLwwzoU6R30Nxmp6Jp3GOvtM//hwuRneR7pPpcl0wpicnZ8071srdui
IWnVJGFSYTMDpM9qSya8gFTmcyP1UT2j8su2V29VkQYINSUvD1YcXICE6kwbdpGI
/V6rAMH6iASAABiAYH6h+9SiHxSAn9L9jS++wlu6RE9IqPm465KAufmWy+4XPLWG
`protect END_PROTECTED
