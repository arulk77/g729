`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNX94aJGqTStUI8vA5QD1eEPAnR75r7bouRm58ob5T60
sCsGoSou+GKintxXaiw1CAuHBH4FopbTuDyU2CSzMsqSj2QoaWsCkBwuTQ9ZcAfe
khKcvsoMJVnHDbzmmx/2tPxiPPJ4KKPFwoNmaFz8/GK3YCmwVpcqpyDBrVoRuzW5
XecAsqRD6yawWdter241NF4y4byk3+ZPHbjhvp8s6xeAm6CVr7mvbqbKGmtbV8O9
`protect END_PROTECTED
