`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveInpWsC+DRXt2uRa5slDDUm0m81RtIvIdi2zMGyjX8yN
RRa4UnGGS1oSU6IsPS+D+Q5Wl9l4eNMDjfoCMfhIn94uRE7Ufd6OX7fooXejon9i
hUgsZD6JQMHApy/y8/3X17OoC3funEChd+GtQNFiSHQUly81y9+PGN3iwDw3Ab85
u7jl8lHY4UNxrlFV/QqUpc6onlLrC/rDGmRP9C0MUPTvoENKboTDJBQhX/bsZ/cs
S2w3zxvEmSPGDLv457kPN/eOSYs9+vidU0xmETwNOvVOKjAnzj6QY80oLRC36Y6Y
BH//Jcg+3WynOXxHFaAqpQ==
`protect END_PROTECTED
