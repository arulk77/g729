`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8Se49Z//iDF+hgI88+oy1lUzSn2hwr74zrDcHRMATFiY8
FYfv2JcLXgPCBKXUfvmcan501Mn/vxNsyp+YIMCOh+JK4NwKJUikkd0J75JDHm5p
sI5Tc2BulPgj+iO+67EJy7JObRNk2spujWlSkrMbgfzMjYeY4PmiEqhLpuc1TB0t
76gVcKOgaqkssNAyE6fswRm11BniI+/FmE2OqQAtOhj9uL92fWNoRe3XIa5W6fb4
LwbyHucZjvo+qDS60/CYDJ1QP1hfYAcaTmG2Twqr6L3tbKY9sjxDZJsF/Kd4RNye
1hBa5utkMzuVsubquOUMS6ICVOVw8vkKutKUsznv5xs1TCcS9f4CXQUA2LoEqxXM
a5QU3poNgtDKxp3XyQqqUoGnd51L+jNFLExoPFv9IPsYnOGtBqyowubbfHq0yCj8
0Hs/ts7rrjp+Jh8TZ48wIceIV3WgqTnNYsUIWsQkY3Ls7y5B02UsLE+0TKmIity9
zHA/AjLpCtPNR3UuHPupoQPzbjQxtLmK3ZjBPUrt3S5eo3BgD6M6AU84N+azXHe6
lkj1N2cDSJH6aq4zmQs6SbTfaeJ+SQOyg2P068/J7IL4QVey2rcYLAvzM3/Dgr69
hrb6XpFcprGYgd8ztrD9w8Pkx69X6aNnc0epqaSID3DIx1iLRYvJnhdQbmlotERw
LhSfSug88TJBdo9oDALVWIz7XamsqjMzriVPruragahKrCo7VymQHAUSvZCIDb9n
ieZppF0CBi4Hj05nvALTQLa4y0NoDwwp9BdT3cRBoz6w9ATCxxgs/oOsa/Ts31Va
cu2ZiRAbspnrWI8p9Neawt3BTUIqvPrjIGxA7GKN4THS2Jaj7NiolmR79jfVXlxc
qoLqeimhIyF2ZUthdfm9evbQxj39AzX7KRdyQpwYsNRRNqimGF0emltruGx0bmBf
nJITvqjJje9TN+ofBddra2JyVyZqS2G9kzCCCugH/cV1cfJvLAEpYNczXwPKtQlM
QisjsiFV9k/oUZPtHR4slU6KIv8XHQaRIHbVTbMG7JyaCdvrqd1sTTwlqdWnSAdr
o4A8bGCt5ya5WYBIYWmACcp4rFKhHkdymrIq+XgsT6JsRz3L+WlfZzTL+am6y8n+
1nG0VLM5YPud6P2UPRH9X+v6188duReD/xqisI7P3BLy+9ugxhcqwijO3ypH5Bej
gLBr1QzN9jUoJUsXyr+Fy0irCrNluA0Ya99lzf18DII3o455p8qJT1czWqtu2Otd
7OfWwr/h3NOjavTjCp3RAo0ffl1pBrtd9KGcJJhnC1JyeeVvOibwLkwcOHUfFULq
uU2FD7vGwsM4NHUH/U8UHNbUQpjlJHSAp1eEvKPrdm1DyU+BfeHJ4/Um5mEPIYBC
5QTUopU621J6LyDobEAYpau9fQ3O1fltLXWKSNm9Ca4D+CL9v2T87MjW/ByKsQR3
JhaiAuJQET09HiD0lcvq84Z/+9FShoIoApdPChf75WCDAbnKRyV4Jt6EwnWhd24Z
1b2rZ+JnUEiBAhANmG5rNeSjeaygm50ifXP2NLskPgwoy5hWuHltoE/WVkms0tRw
p/uPLzLPpegRegkvt7jAXBTF3ZOaHllGhAaeLtYa1BY5ycVy9x230JDtnagbrw8O
LF3my+FvxUJKXSN6sIQ5hDX/LnZB2tMon6o0kgUjXs607qOZNQUxnkHEkB8BccLt
x2rGOMaUOFjN8IquxQMN/G8WW+q69MUqH4y9zA+R/mFHyMFJPhXvtUm1xpn/8X/K
3Zu88YwKX8ula4MSDaCwSetvdTLNHodeE2JsG36ngTZ1sGQ4h8WQ/A0bETmHfjcv
2JouHPo789eJ9c6YOAHVJExP58qmZ0HZ8yXTUQz+mKCRp1ej+Mj/NYpizCiXw7JZ
uOgoBGUs8rAySIJmxF/qpEIfPipRVeqvwlim6o3qRAtBht4CqLE0hpOkWDhz3wyi
HdsLbS0Vj+NKJOBU1L/MIB3FK/IMsDWLIwuwWXHee1SzKU8NPDy8Q6g/J/3mIZzL
kz0rJN1iSUuKkEnWhTx3o+oSiUj7zI+RbVQqJrG108iZotAy1hKCIast2dR7bxuv
Anv48iRk2O0N2Iz99UhyG9E1rPN6nZlejiSdvHW0SG3K4SAZPOhm+4IvuzHYbcqD
+wuqj8+7urz9m/3IN6grzza66c2QiakxzyViNDX9Ljt02lLG+TKN8fcRIo9twBX6
O/n0deA9CJDnQfbAH23I/xCHGHLKdU+mfjOzBA6yC35jsFrGd+N/7jbynNvF3DAw
B28YI2QdNY+LDABXLXKn2XkVo1LcHelMXKhugqIfOXWBZAvJlgpabSvBhHzFOy+Z
EzYNdqesglZ05YTVoRjKJ/YhRpCEw1/mbACWdSEIUUk=
`protect END_PROTECTED
