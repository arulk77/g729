`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C2iZxZjH+wksX7iIO5kbaQ5AZDABxdfg8gEteZlq0Iku
gQiLCjheu120VgmWYZoFq73X47ycf/grLqDm9voG6+O+NOnsb44r9hiv4HOgwhVW
5n6TtB+GvFYwkbLfna0AGfBTf+9+t3CfKq3CbhY7iE9yztz6YVnnvPg7AZN8xaiq
Krz0e5j8Ad8qaCCcnRKt/gPUGY+ojciMeaCWV3HxMV1AkJZM8M01Wm6Ur27Kwp04
+p+lj49PM8uMQOBah3d80Z3QPS35avRG4jHgQ3Gp56P/bWYv68+czLh0ZHBz/DzA
Jj3AJ/qb3lyARDd97mQrnz+MXC/wJzNZSTQ0w21Pwaaqam2ArC8UINC07NvwPSV6
dFaekj5uvN5sv4nbsk5vJUzAYGHVzvFCI4HDXrFSRJOB2AyPDBO49fxh4/X79yXH
XHaClnPR5Yrizp7M/DE2Set7Il3e4/dHv++/qbuMFwnrDgO4XPwtDbbXqhpViaDP
HuE+pP6JVJelfYbJN5dRN1ScSqb5feqysnVDosJh01eK7GBBqMhB2/mpzu3Rwc1S
xM0E8+zmv0tT+L0Y8PvS6MJ/BaQ9PmEuDHg81qcz/BlFXQipwMCgCaJaS1qqldS4
r4AvfKiE7EFSZR5heobbGg+DzppXt/D1elkckVSYG1VC/2zL27UnYx1vGgJTerZa
KG/vEHyBJFTOH5nIxHuu8ZQJJvan5xYGR2aAysOtlh42MraeZk64XCqbRsD/r6dl
i4yCIrqye5r53IXoNLAzVU664QtuzPfc+4fO1qdViMXKI9BtJAHYRXf4Q09B48Kt
D3UJJR2oq0TLJcT70NBr+sRyPFs4LTDdwlf9IU5S9WqIg+vvaSXNfUQhhByHUZAP
hHTrs59w1YhCj+D/7AgJYxodgs+hVXneN9tLns+RRK7tw2T78Y0OX7sERyUVMoP3
qZkkkNkTBTd7wfDXKoq6iez1cQVPyTiIpR2ko0jFplRHuiqgGKRt3O6fc04NKtly
n/XXuYAcQF5RCOeDIeR7EdfhntRh1onds14rcUp/CKw8OqGl7UyNKS/K7CMmdwY1
EWCReftjPrD5WkNeBprsHHJ9YDENxNvBYn785AppPxtF6J46qbqucIkep2oK84KY
5HDvQitvttqzEap4M/asVJI70wHbqgdoEXq/1EiU1d41phEGJN6CVrLeOGQsmaIX
oNZ4UWp9jLsnqcGXGpfoiduKJaqFZA2Ttr9AKjsrkITW7KyBD/rM43+g/ljn2d5W
TKZhF6Nqf1cBeOW2WuXdiQ74f6bimr04yZPDm6PJ+HQiyMJc/2sTwbHQnIiY4Z+D
lb+nFTITVhHlJOWQ9/avoWuAd1UwM7wEgO+yjHJCF2vi0LIkHtPCdV5AYB5OPnob
wHY1QBF3wrPcvIf+ZAnE46HaPgKO7ZKA0Lq6S+junZhcZpXWvHFCt+qkx0OnYwlB
CmjHU+7h37ZDrCeH+3rKtjCWHi6WO5/inx4eYc/W3QEWnLaVEk3QsUKpryk/vomG
/7DRC96L8Gs2G7cVrroZgVxBb84IU2N3uQGLhVTWBUwCbdw6zHAo+NEoygtYomHv
gPFQNIr3gL/P10k9Yn4JKJpB1YnuGXGf1zeyqgybviOKmVgmyNY/d3f7b/z7DrdG
syGuv3TsrZp7tT7S1gDZEE1YjOVv/pIzs6vPnUtIEjWlWVYYfkQ99ITGNNc1PcSc
fFuusImZ/BjsFADw5fwFfCctYkiFcMqSt9hjf7UhpyqK+oNu2uMr11OPBEON+/fq
FuCUrphhZBgD/obC05t6rIZSlDKcmNTxVcC+1FmtyyE=
`protect END_PROTECTED
