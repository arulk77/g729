`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
LlxB5YqF/qI2GenX9CNpgsvuCiwu7ome8U4oYtaVqhQfLi8eIL5wljgXcjVzIcJb
iRWKGyOfAZ2ps6SQWvIi5DCHo4/03/kGJy/XY3YMh6M83hFI6YRg9nSIJfNIACru
IpA//2jQzGfvFHJKKPmHk9wOexEr9BNSocHlU0mFMdZBAJvCV0Volgn/WoKIo3SK
2gDrovhUyxQjSWaMqgelwUq09n08r1HIq8/refbIcqhTzXp9Oi/Cb+Mv/FAKKfWP
NDR8CW0trXr70OKTYw+dLIGfv/BR5pyjE24VsnIDuxf2LkPIhVNjnA+/haY3MHPD
mLFlTJ65L9d+ihJGJEJueLmF/wD5kCbZEmfFl4CnbJI=
`protect END_PROTECTED
