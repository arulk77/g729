`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aJ/0Z2p58rwGIy25OY1AHDhYpi5z1uc6UopGdzb3S8QMZa1jYx4mITAs33IEDIgf
JthSXCxmnikost6EiHFwRb/Ct2h8O7/6cWX561OB6Zob1ItMxFEaiRvbkdQLSbUV
JoBaO7TlqFF17sP5Xxe+TvMkhaJHLKUJH1dHRggYCni5V/Ogv3NtjZTw6MfJO3Zl
XhGaRQsBtdDxxlKPtHl0gj3s1TnuhGG8Z6wXoBgbpJHLqSEzhqQ5pfpGs2oEgWzG
7+S1hywHSn8dd2FmT9ytfuGdOl6Ow82RpQ8xmCpiUU6IlJ5YaGhf4q/gjSMasntW
ZhX+O6x1dJWDCBti3xwCR5bgRC6P+SQV9qzfJyW0MYpePC5HOxqjH94Xe2FGH5Ek
JUzNf34KtawSMgyM4h+OdGBMKGNKJvItFrgKQs+fX0qJPfuJa5Z9K2bkjnkE4jbB
gdjqA7vNbHW4EYABv+a1l02yOEBsnYgeWyTXqiTh1RXp3LowMkiNzrQ+hwg28Hkg
wZdlIYkSYLH73MIQp2dC/tSr330UsGyZDh9pcH5I9AYbpdJHHQuGOLdpn2ed3wbs
KF17Jqv+zuXXwdTrAkjb6bx+kdxEMCS0HYyChVi0YvyJNazEvmlcvrz2RhDNugis
EBpBpqjWf6pQfgbIlzc1D9cSgiMkrMChCYQnawVCMF2xmmnFQbMD36zL9xzFtKW1
9DOuVcthzjZuZzu1yLTHNIMa2oaiCXLUrKOEzKrBhWgb2BnVSxZYHm1pJnVXelzA
j5CzXjUGEFW2Xmp6VPNudTSwX7WZ61lyt8qT9+AWUcem6GzDEg2+iMyVwvB4ECB9
/oAcwanrmB3+MLkk3eiKAAW9tWzD/J6DGL11AuqNXjum/IBZ15Ufoxug80mWwFuc
qvMxgkxC2y30rRpblzkvaPcS0JaXp84L7RDLFt1ij+67AfkwuFly+xmtwg/PAihR
UfWxuYRkb/xNkETMRdQOdXokg78eUt8Xhy2Qj/TtroSO6SCbtLDl5I9IHu/BfAPU
63ed+R1CB6SlvTDd9compA==
`protect END_PROTECTED
