`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN6a0D4ImYzNbYPd8yVSJhS3cuLVvyepi7jjd1ZcuC+8b
dkbyRZbchmFf3xfCJon1vuGPGOWqQDwkjsXTMVO50Ls1zDz1ZKyEzOxCGEgGhNqN
TR59Z89bHturi0muGK3E334EaY2tGMPDwdBopM0DcuDwe+OuKsMzRrWxSVDfrsfI
iELrzeTZH70ZlUX/7/yVhS/fSen4fPDp5AT5afmFX5m81svJmfVcrKKFVa1oqgEE
VBOJizIdpcJf9XdMp+WlNqteUdPak01nBhUGB7JDeMuu/Ddhu1rWkSDs+L+Slj+5
tMUXgynabcZDWn0pZT0/fqWt/MnwhOu8St54HSsfvh4U4A1hV12Hwyi5MphBK5ul
8BA4v1t4oJOsrSs6fPYSs8ER5WL/LM3lfDsDhHD2m4R2kGn0Hf67evAeWqoReEfE
kVdCgRQE42Un1MG4fq4idLSTdNQrJTdtjrwjVHLPIHc7UVGdPKJPv3tTSfpKq6M8
oScPf8tKYbNRoLGzLj3pr8yr2RYTcCqCMNOYJt5lRpzWTERQ+9UGSaCZ0Xn4gDCB
caIJ1Y/ddCO4DlTBX2ChtPn0r8fMjBJbrkzuWW6EtxA+A2n94OrRbPIh6fiEkFwG
v5Vap7YDgB/OFP29KrLg/mMtCwU9UNk03ZuOLk+IE2iMqLwqELpdu8eZPnnKDMJw
IeRA6Tq/+elgD7qCn0AnmSFaajMl1buP9SpOGCtJYQpYBe0O4jJHoRdPPImV65Hx
SdZmIdIZI1of0IgXpojTP3w2jZo1+/Ogztc7rKSVAwFQc7aElS58JyCiwFz17nZb
6rrFUvEhxsz0UBCS+/5F8qzMEcu9qMJQRfy3kfB+FvwYfw2OGFo++xQeVIUhmqFO
0NL1fcCG98HIKLnrb1iG7fCO89qdwqHJDm7R/MbJYULRAxHQ5YkZBtVNFl5AtxDN
3fOm+k41KxSWbRKRBfPejgVLwJQqS/n9eLMPZ4Y71u04u38RM985PATPLioi5EjI
D9DBgMyoZ8G5n69xsaMGLdRw6GAixsgM+9aBHudqBMS/h1zIF0M6s1j845wbVaSg
RbeMFk6t/i2rrep2MpAsVsIzg+wmvEovWyleIuqzKojBDiwYtaWG1vxSUW13V5Mt
euXf/d2K+3oGOkrs4OjsF3IGbiIq7YobzcXZ3v0NIbJ6qYu93orJkY+2sXzRTL1G
mGuuJ4w0Fr1bUDODe4R3aRVRgDHIVC+Y4wA/ZJtI4pU2jO7oCUy9GmMwp7cDoui7
DPRDWxwAd1Q1J47GcGONDqaPnUxTM/JewXlLK0+1IdxN4TON4DNHwr77sx8SWycA
SlimVTixJoqRMhE0R6e+/e8dRmSvaqq/DdE/qt4FFBOzlnd2t2PV6JYdICTonjqU
CZnU/2Acv9XdRcJgajHMWWLF2CFMpVyRViVHd8dOQpAnuunbPQpD5uTIRYVA1zp7
9UrMeDporcwR4K+A/wZaIMy5xV3XYtIx4pmuLXdKMHCs0x0LTSID+rp0MVMJhQtk
wecYmvi8URz29EwiskQ+zLrt3vrqqziz8FyyXWhu2oE4RNcWBCC3SjTNrb4oV+VD
`protect END_PROTECTED
