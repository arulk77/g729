`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHK9zqsvS0S5bkTIUJhVlyN7S/7xlPQcqXvgEAIfdwGZ
8HCIQj+61hkHDZMyBl0e49dm+6T31n07HLHnSS4IWjJ3lsIJ6Q+5m83RafblgLYQ
jIzHcNBiLxdF0iPyNEIV7vAsJGfZs+6vw/FZwv733AFmPMU91A4f3H1YMz+P+/Tx
4Vm9clgls1l6DrRZB8nFDuLPcQf5OX9eKWPN4G5GEHy6l8CYzvcyYlLzWc5usxD4
dXi3LGSIPBe3zhXdL2nfyQzn0MDvAM8LW5Ts8OTq94yM/G5IVdsE8ktD3GTMnt1A
MiWsDxC8XbVN+MW3UYk4pnjb1d8CsZr+R1zXix8zJqUazW1eqyKSbLkjv2ruDscT
dbthYX5NebPtkwmpgKLdt6H1gYKW2ZUTbmIm/iFOBH92FNxRPoXxCD3t1ouZrF2U
IqUpGJYeQwR5wZeZ8axrrsUU34r62FHmNcZDMAAjjUsVL1ZJ8bi3gv7a211HcTc5
fdqorf9h9nGWxVHCKPw78kOrZzi0lj/z6X2JHdRvDO4Y8p1caz6uLjefV1C6dq+r
pkLCz7kRhSHbnFQjwwsDQdFO+y8z0JFJNk3DIRzKnQwOVd2nYtGeKZwyppKJyOzY
9dlIjfbQick3HH97ciUcU9JYy1ckOCbOwYzvUbbF2X25Rmv7pGF+SZSp9Yzihlgk
`protect END_PROTECTED
