`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
f11uP3tAS38J+2XEq2c6cKXT/yGjZKW/iZ5YOvE0j1O/RcwqiQaaP44y9LPLErGk
0T4Cr+w3gMTd+JQpmi16aCaalAH0kK9BMSr3ZBvj6x29kgJVJ2aMGz5fzaZQjZhj
EU7zMZeJst8x3kuHocG8bQe8xPii7gm4FMbAwG8DYhiohI2nQ1IwkWwg6D1mSvoW
`protect END_PROTECTED
