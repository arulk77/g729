`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJdYZZDk3tJU46VBCXAXIKhtkhsdGdWLiwhxHErwqTyi
qpeQfZzygVJZqxjjfPEzKSub1cHoxkDVu2A4f517eV23Eu3/q+ydJcN7hP+P+1+/
QkKTeJ+47Ms7ws4DKwFtXQEZVbvvYGqn5u/KGCNg7aRnOyn+56F38Y0Uv2xJfy6g
9iD/iu4yetBbQhfoS3HAQBJq6DW4RgFhxYDRVrAh7kbk+nrzXl2T0OZT2rLneJMS
ZrqNYlJnXDcuftbRKSeSDob8CgiiLkWUZfheiB5AzRkEZs2nwmZh7SNV2sQujLM8
N7MXWwWiSDoYfL/36PtW7gkHi4UxqGHgn0AgImtGvBUJnnYiOSjqbByL0CzjbW0Y
t3Rq5l3MiuoExdXhoV6NCbLiD27OVDeC0cExmNey15Yxc4RwnuuxdCoF6tHiqAfF
ENj88RrkEmjeSTUqDj9egJVZz7t8i8S5JOnir+0rM7M6Gn0vgqoEPS0nK3Lh228+
YtnDS8eB/mzPd7fZ7iohhg==
`protect END_PROTECTED
