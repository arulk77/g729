`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveH/HGwjn3YxicjNqUiFQlp7qxAkSJn4YIWAx5RUQLlX1
JWHN2kA03TgmGydqGWCurpUjHd0h/67T4TPnOHgel9dK2/F+r13xipMvQS4n9pSR
yLfrGJzdTv3qEYhwjlGYNcHTtuOHllwuBXOoltiQumc60UC3rn5PDFFQEb4B5UjM
DKM2rGDQPZF/zeUUQCXe0pabj3BjIOiRoU3tW2snmoHBsHehWC4LfeNhoarEcyOG
4HvRsGXia7rOIraBN6WfJ4q0IfwLN0TmlyPZrvwSEkclriQt5cw2LqJl49/3uI5+
mQEorzsSHqpAIF76w1qgUd0eMSL4dCEsDBEATCKiXQhbGPcXqctnB3gcfZC9nS9R
4ZajJR8VXfPYJmeMAqSJ4uu3x0ogR84wHlKjqSJ7/hr1mSR++Dv+LHUB6gJZYvuU
+qfWz4uCRisM4GIZwCi/GV4YlYusaO8xX4B8iAHs9vrPx1j9klQIifEMu/S4b21s
hi7BNmfjKKchtL/+l6iCHL4MWRaVnq3gawUglQ6ZE8/Bt7IZ2w00qzgKi8QBbDTw
mbkBbBj08ka/1WGn3HVfcvhe7kDiH22eCLQ60e+HRmUzOPw2To+EANmPyU1L17xB
`protect END_PROTECTED
