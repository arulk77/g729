`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ2m1kEEfQJ7ykHjDyCMwRh/3N1LSGK8hcLWQU1RQ2s/
zmy3Vl+Pin/WxQFn5jQ7k7yGBMLsTJgigJhqSrtufTnKYezodpQo3AnqgkWnH8fb
kD3PNX+9P5R3g+qyxBn45DLzYNHYPEqxvdzbjcha+qghdTk2wULD1H7U4JxWYbtW
+dMvR0fLttzvuM/86Y3lcY1Bve56Of1PpPA9TMSBieEcFF5UVohFNBbkrKrTPabZ
`protect END_PROTECTED
