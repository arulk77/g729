`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCBdTl4oEEWumAwJ5X/fXbn8b70EL4rkb3ddoXN+EAp/
apdRmkEYMqTC9CIdBnDTsxzrrOkPP11NurXhTZN7tuM8hDKJuwiM6Cze1icAE/gT
zYeabPPr8AoLklqrROsEm43VBsp3PAuH+otmjqjzItmUN/zyJcQEojFJexr8unC6
udl8IFejIXm7WnZLHGZN2V+vO6c22tkCG7FVVHA5YGgP/DkTO8egW2bo/NVtQ0+p
YEb06a6qaNW2onNJwEMC7w+MNlH2Nm2A8El5FXSEgEYhbibrJu+7wMIuzX+TaVQV
T+B6i8qdv4miXje2ZRbKB19BWcFvtaDcRvd37IqLNMUYebL+6ceA2eo+OO0ju0Vj
gvjFjTQjDSRnjepba5sEcJVTtUefb6TE1nE0AxhyzFUphw52vV77I2mfPwMmH0u6
MjCtjYKjCZ4YDHxs9O7Ap1KSLL4QWapXHMVky6gxz/5WtzKE8qBa+u6JcALMSBB5
LOO7wQXYkgkyCT5LkWub0g9DJl9Uwm/WJnwudYYeWIRl/TWmcBYNVhVXHcO+sq3E
0TylmOlcvysqaAN9V5Qgvx5RmYRc+2FiQeMPM6NeHPjH0XCK8sAgSdynnshlOgbI
hrSIybjWnBFxNI9s4dDs1CG/XrQdc7SwAQdpfrBkwroryPzSZqhgYv+Cu2eNqiKY
ZZJ077lazNfxoRrH+W7MK2Z+wizzheHIFRc90zXq9Qw3LNrV5sqXuxJgTm2VdLWq
TVKv08OfdTO8jrd5Tw0qGNG36X7HUb6psnY4AZm4F6wu6RKwSrwPF9Hv85IYhC46
XIzEKdAuvqUBiZTDfMb7Y7+FEZ37/ch0xVxyqmm6fq/uIFR7xckqj9pKB7VaSsI/
lhETM/XZi81gfo9PasEqQVlbefA1dVq8yLG9WqyPxzqt8Jz/EnkatDpu6XTvt0IN
FEuKL6J7iCg9CFI9Zjrewv0CV0l1yzT18lV5QiovoZSScWVq37bJz6fJVM00rcYl
2628v0po7qsMyo9jCNtfZhoB7mdjnuwHxtQXDoHXIP4oGbw8JVnVRpcwL6LOrQSD
qLx6VXqZH1pkQCLbT0b//EqpL9islM9vHAzUiHln6hppM/Cq6RcOQoG0XKs7xLBe
B9VkFUs0oqb/TGgrDraHTGXQDc44Fkf0K9XGoPGQljVWN9qCFSjhwpUEjoDti0dM
F6n5Okma/2U4T2BXlvH5oorLVYT6QI49/DLPOCVpZ7/75cwnMMr8BHdH4WXmupCw
aTGXOEKzo+tcO5Uem9DXn3k+76uNTEETE0uEErxOz/n0/FOTckLrA7oPaRB8PbfJ
QbRqayru8G2kB0zwkSnDwbHnuQv9Sz71TndEAT1s+ntVKoTnCS2SVwENhiyvvVTm
2ZJ3qzhecTviCcji41nL2+062zlg0iOe0023RKYxXWDMWwmByL4YkfeR0L6CR6pW
DwuSka9KS3nYUj4WSpnJEk3tlVpKXVY5BA4JsuM+6nVept61a+SlnjbEEFi23qOS
O84+mWVY7x6fixzUv1+JO8Sj8qCgQxOE6t6ik+ZbYBjp+F9Csy4jznlKwFobb45/
yfGCPasiH1YWTAp8QF5Fs4F7mksc+48/srvFcE3lKF1XUUcx1O8iCfVyBDli6e2b
WwlMCqbr/CmqKjdYJHoN9isdLwA5ErRfy+m2BCPA5ZjDmk3sF32YelYkoTV6CRwL
QU+u/rEM6v+BoxpkjQlXjLjuIlwrrqYmqlukGudXDOxpQe//iYshijudBCM/2Gqj
fnDBW28Iu43c2tMJMpt6fHPD4wjSjV/O2oy67BNwF+9DKaX8rSo+EsWWWT9awW8l
GSv2DUyd+39HWlpbpDtLhqXO1ND7Piw+E/RZ1g1SGMjkxDkQfK84UJXW3NY7TFar
shWkg/9p+vcnWRUQQHpF0TKoCY+tB1AGQkdCUCNOcNi4glb6bXnyhO7zy5mAOu+o
8MxmfIVmu6Rpe6lBI/YMfwvzlM/xAnblPnZl5YcgS+eYOPLiASv4QVtg6ptwmZ7V
8Yyo9A84UPvyiqeLAMkl5yc2MrJMENWpsHJu3uTethUFK59eO8QfXYES26pJyAvs
JvQ+7u1NPimH1TLFDvsbM3TI08mldvZkrME+MPAIQe7QmChV3dRCGnqIHX9pTmmE
RtwpU5X7QNiaGmP/w7dizYkd8PnUpqMb7L6dvbitfV+Ep1Y2rf6zXnxfne2XjwzO
N4M2+5+0SiDZnk4XGBOSTIPO/plsP29Ambp1v40TIIG+XYC0zrQmsxTm04TeNRX1
qhmrSayA9SK0JDnypeof/HwGirqLw4wSozRhb/knc+7Ad7lyA8y5fLB/E6ZUSMs3
hk+cvLrdf7xGovL2m4s2SRTG9jPGxm4cnPQjkl5p6nuwxgeFW9Yjk+F54/8GIj/U
yJSab+jfvE/E1qcKUlsot046n83AwVo/GAA95tdZUsVNFD0J/AnB252z201Yuhqn
W7FDmjS4rwDqvf0NO8kgWYwajTrfUpVW3QPns6oKTCw7D0VlsOvWmX4j7FZoUqGC
viov7rvjUcB6LF/w9YHm6HBcAP/YInR8QZPLbLybt+FYTlX7uoz22CvIWLG5Gmle
9BNmQXOAfYRygBPDBcs7nJAbvfc58G5Fzrsvxl2TK8aXd7D6J7sb7x8T0WjRNhp+
sbI/9K+jHvTfCw31OS2NDl/ZM62tqj7GHf8Hkqrq5G5hk78AME9pOHeyQdh9bj5c
HYGPGcsWm/s+2S4Dj5uPvoWb3C97+/EMMsgyn4N7AvKL0rGbEpUEqnFemPCn28GD
KX0VpEguoDZ3hK7U1ttH08LpkDcLFbO8Ue6PDW9CnjxB9w/0bYrY9zp4QRSkUdzE
ebF9XaH4mdeQImP9z7HhBkLT9mp4x2J8LYe8vMzZ9jodWF1LLVJXCNKICzGcqg+c
d/IcImrBltMSXGLIEi65XpWTwH4eTEbLJUA23DszOta/DFNROY1ntC/pVuoFL+IB
QZrw3wONkZOROASBKREB+YOonaQybG3uOofPJnzhhq6mY/YIHyRa4SC1AHJUkzna
WQU3C2Si8YCMf6Traa4OS0QLZnwhQpeTQbAr+JD/DFH8mzIw+t1oDILOU/5xi8sh
oie/DduXJn5iycCZu8YdolQw6x0UYLyqAr4lKhxqQJ2BIZouwvKLfQDyMCYwMBSW
x6sbtjfaO2cPQXaL5nLvKp+dWu43VCQEueoqeGYYJC10jrvY9I+oa7QtrZmK9i/n
fU3LVy7Os3a+9HSIuwmYW05LkpKxYVbZrIx1BQEsGssSusIy3n+zOlXi9gk8NIRk
ttogmDRacBvKWBL++Fnrv3qHDJRpa6wrw+g6+NZC8rXoP3uMLx8hz7p++CCnTmKY
7yD5yq3ndbvfi1FIdzhY4my3IFhUTrSM1pV8RnAPRZforkj1VSJ5NIs1smOJYsSM
V422NulU4i9ptYuUhmFVV3QWWTbrnO0Rs7Z+DB3GmhlhjiHzoiE4Hvo4F65JFgFI
5INY9ey9xQXcUGayO31CFaD100tAuNlRswxkWrdF91fuyYFrtWWd9WjRBQdY30I1
3nRaavTCfXjZHRPxHd8wDnq7HMgab21MKJcPdfXTjvwMHDOjOmjIAFefDBSRkaX4
zQ18glNgRahDWDH/H7SfzPRZVD11GC+bBIXoQymOYEfo1Gpo1P+gi9Z9CF0AGMN0
ktdnEQH+QU3L2LLkACt07PfCEsgnBVKbmPtsMZwt8EwVmxMlDL/F77X4v1Dz9Aeo
xYwy7dvs9UXHPZBUpsUBBYDYj8/3ZWyrA75LP3bt8wNhzQzAv+NiRQdi/cR+lUcV
XKThXwVn9PCeMJvchIgRI/8YIls+fx2wS2SQVDgjZJ5wHGOv+ljb1PmLHJ7gpk9i
yHnae5Dpul9x0qKxmk3wn712mUo6jbsxvQUPX+FhRbiX8TuRMW3+5VXLpj8WXUDL
nrxFWjWKIeY+ozTYQj+FWnMrjzICWsFIfMatM/QDgLJBXWsUrnKfKzL39Rk1AorH
OJ6bzcAIfo1ZyJSmtc+0RCPL8BV2/13rqJcgFOjO36olN8T+Tw6fgU9b0qNin5BM
ZzJVT53B8YiOMXhLaARCDLnZRhZN95SIakK+O75xBAoKhQfDMJhfSMikJTS8cap6
40XvOVR96+s18JbSpCBAOLNLlOEaeKGlklqa6wiilvHFKWOa2sMFw5+sEQ3a7cFa
bIgW604XT1JQZiJJ6KFhVPFOsjxMryag2aZXtJNVzle9MQb2sSXCboY1rLKYKNhL
MZdCabD9dEy7xLsHivrfjv3EoW5BLwrf7KAZC8j641Xyqwn54RvfzEFPPPE9vn9p
yFeCWx8JROAn2mfCOoSVwszQ0Oi5oTAmqq3wzqFthQrWYo6i51sokayfzBzcJriQ
icb8zaATghyla9Ma93G+oLy5uSwu1M7J2PjewpkwAMupjKx2xU544JJWi/WesNda
UE9AfHsb7sKsWdR541gHhFfSMHAgx+beYTr/erJ3lk8Y9CSqsF/9THn5fIUV3zXA
+9S4BJAtnO4kC2wnqzGD0ExRIvD6F/0pNtFGSNuxJtuipva+evGKkupnw+NhRQs3
a8feAveun73obYtcsJC6o/DIN2HdgABvZZF6G/yC3i3eFEO95prDal60wTI1KKlg
I8/ynVQtLLSIEthUXw740DMwOzMSKJdEwAknPisKVQ5Eg1XbhexTNBBaFtn+BvAx
YWvDLGa3+ZEsBMuR0NwgbgfYT2CBDccSs5oGfinsbvByqmW8a9o9EyxdH/V9ovGy
wLKlHxi09oogH/wCPMXP8moqSTtnUnRUxwfmV2/Pxs12+hkhgFzi2NbKHq5T7U/X
d7PKBQZahHoxDtgWFAex06ivtlaZglIqllMENnwhu3IlPz0H70gy5O2wyiB9x08h
M3E6KxQXGKxPThE4UVID7WNcXhy4pwgcZnC2rLN+zT4I5/tKCfVvGS5j2vbEKIj6
IyJi8nJQhOWRy2GWcNhMtZeWpx2NzXxB5BCv345/iGNVygpc1kFOuDQ7lRsZVIWH
/9mG4Ng35keiucJ1bJ7WFg9SyGriuW7RrYMc6kLPkst3RccyObr5z7GXeMN0J9L1
S880qS7UBmi3QXqohvB1I4JCjGcxheRK2qDS9Pvx3pmk4D8aXO4RWfOK/dzUjprA
bdMk1dLMCYGDj8IcVQLT9ScRgh3DThhMNmLXoi02oqOcnw/Mq5j29KDQYECuZkiW
cBsrOaPhTe1hJVrRcQkN7PYUVLgQcGU8keyfABesx/QVuOTK7xoPL4VGX1gNIcVp
CT3py0LbVJO+H4QWUCpjRD4hLzs9Xi/IwpmOMqzd002juo8m6x4BvmVlpffiEYyP
m0qZRsggWmYCJVMhLPqUO/xNXKbMKXWG1WhKFqBJwGalAne2INoi+1Kij4ZeLc3a
LYjW2Ff8C4yIc2shryf0HHwqZUba9I21egJ9BBkTnGFQvlep8E7RIowbDrFCrQCk
rTPENps+UEpaj5cfnLhFojofQDJCx0oKQwcugAo1/DFejC2PMMMov8BsaP4uzzvT
Brp6Q4GDaBdeikNlx0ueOx99S2UJrPfmJpbJamwMPiwgcRi3FK1YgRiyNMO5zjmK
CB324SxaJ7YoyfK0WUQ+a5GnMYjgjHg8TS6DbZGwvIBaHprhfq3tAqhLKGQXiwaD
YDIECHY/a9VHrSkVRnEzhfrRL1iqTtvlYzXpk/UBK3is+kiskt/PU+qTy8X7NElA
ySGXtdDOdITUKaIKnziplpcyaEGK5Cjo6Z8Shi/gsX8H7HJK5wyneXVc/jJDbyQL
J68ZG2h1/KAxIiWHK20RGaJeXGwkxfo/znvUs7kvlaQUyJWCefkpVUOgkXJ4fZsm
TWlFaCHSybe81nPm48S2I3IzBcj3dl2lnAirqBer+3gtztLS+TDdPkeQTjkMQ4DH
HXOa40d9aDBTte0VF0ZgBYWQfXDK5QjnX2QG77ovSBI+NDeGld/vkozQNZ9OT5KL
CFhHHmyDPTrOcs1KIoz2Q8JofeAApPwiDPTKjHwKsKrCOXNfCjHuU5nbIlTt/VGG
cTRfqhKmdf2rSq5wLqpl1PQCIn6UNJgvLo9GocF1L7kswu21o2WRQG+yvgGXQriD
RiGsMC0o0rgwTYZ8sWGmd298RGgG7A+Wf23KPk77MvRw84ZTfYnX7AcWAlUBlUna
1pb6i7uPx2sDFlJgxHr4spbEd4zVvMrLAtqn2aW6W902LDblBhdv7Ld8lvN49vbO
eSY3ukQyG7yqRS6bin3pkar/DyFvr3DHB5N8Cy54KjZAS/H11eMsxjBGaXK3f5Za
iBJUKNLlTo8K+JCIoiuk6wq3ZY0M0FzDRkED3PdgWC+i3A8z8eghx38NMLNb84Vn
7qxllqfc1NcUEy3RS4OEC6LmJqRfpW7N+GWwsADytbdZDRT3o9uardskkTrY+DOA
lfF/ZfqBra1NF+zOl/pyFLZXutaF5jX7cXg8kyiZnxcrghKt8R1EhxkPXjB18Erq
+ENZv+qevuNaDCpZHo+z6WhRNqK56UvrfckdhiBSpvubT/mfsR59nPtAQqTiwO7r
acRIMgKw1rc2ckPw+OZbIB7EiJXGaoLDz1k/2EBwxqiENMDslR4VBx90ppDGJ+Hn
tXB6nVQM0LkxW/j8d/rntNAIHgi6Nx7sowysutpQgc2Jwvue/CXRs+GmsGcNOZKi
j/v532JDV1rZhRaOPp/wvKcTUFlBJBruQ02iAWxmW+5/62Ini7LCUJoj7C54zD3d
PxcvXxtc3ZjCN2qcm92gOxck2wfgAm9zZTWK6yWpyccJDMArYP8/yp+FQVku0fRy
TuxpnWpXDLWX9ohDqeHEsoCl0bdL5S+j75YKPYXwYOcLNY4dxVapDNo2YswU6LIQ
dz/Pme5ygwkk/jUgpSOMeXChKTJyL5YFHSZZNKhLg3dW1cdlsGKb71oF/VSOuG0F
J1MXAKyelB9cNMrOq1v+m47eQakuqNPraePAOnYFKAb6L8qPrXgCmz25VjW38E7i
aFuFD3bvgcwixI4ncpmrJc6NgNIX2cs+1QjSyFq3VWrE88wWe/l69nnXtyo7c9UN
OoezNjAQ344fz9mg1/PgFLD3vwu9QLj+MO836pW2L6HIv9cytnJX243o2WlEDFij
RVQcV9OFEp5jKtV2Gh6n+NWLMWeMs4+oxGemylBnerOw0Y8pSj82hLnZrhXNrECF
KSMaMLCM4POTtzEQzAvBM42pbd5ii9B0rxaf890BAzxP2Or8ZmnX9hnE6tIi52ES
h20vgnc1qSD2Xp58IuRBmJMYKVseOj/Fac5U8NLQMfrbI8ilJt3e4tg3pZ96U7G8
bpqGnLcSBc1kxaMJAFO88Mz/jnETmH1NoMVOyCyyp/v5r/quZh1eIUykMKFMBZjT
9FeYYxz6aE1AV67SUVrnCE4BT4MigYKxKHr0Et8Ej/PQ+nYtm4YQ+R9GFEnCp7FK
MkPVgQWa0fPrIRb0GelfFjlUF3BqryX5hbN8aHXERAW9qJKiOpywckMSfPl+MvL+
GdvOLOqEAxCtWNEmkwOmKmFKnbdTLIBu3+iY8UtfXMVs2jE+WJVoK2xNM2YWVQvq
9B7uiW6i9e9+dlt0WtknkdNGQi3UysMoj8cVRESXppnzDTmZm+iqQkQu8HzouvBK
Woldl/mKTrvS59Py/S4j9PJiTqP01+JHU6sV382Muwzus0JPVR89Q9bDCdm8o4D0
cQOFCYgMl9sX9xWxj6x6/sGlU2bGSfEA4k06idjp3ekvdYghI4wo7laePACF7Xvh
s2sJMRkdpIqnO1EY9AdzgsFOgBPR6I3YA0M+zwqxSdeIvclGwwWgr7IJoBJFGoJk
69Z+kNkOsfWDjLemdf3Izu5BTgP14QUycRVBq5+se+eRoH+1+8s/DU5/mj4H4Yx9
jApjFqFcilqjPJqGKGEdPPBHaijsw8RS7MBXAqJ/tYp/iggpdslGqREgW1damfX0
mtWTcD7/XXzcreP5GqJfIgUvd/l+nRnk/2gYcMZHKsMiqc3bGpHTC7PwHFOa2KbP
dFY/9cCbLJHg2WEI/zCOGQc3Dl0hGp2xjpndL1Bcmg/1ZmZU9+yfDYOpw70CB8Io
5NgBZVfuJy0GRUg6Sk1kJHlgn2Aelep+2+sp+mI+DYT1sSYJaap0RS9X8wE5mQsv
WuecwlrmXa6Rcs3XM1GVYnq7THrW194dtemK4+fO9jI5p68T/ex64h5T45nChbMJ
aKXgu5ln3lz9F666vVC/C9KsekiCv6nXPpoaQbgO1XIaGfvjgwF37dTHg/n8DBQM
hCpusRMUVqkMMBjEO1v8Ka5ao/kyWSCIfvzrqyunY0keDNbnil30hWpwDtsIFuDT
gd0spY5A85q4bW+1ISvi8nu1pjnmQFTuJhJJ6coaUy7lP09Q+GHJ0BmzZmtugPi4
bjdHZA2jDpaf+2lZ3IqLDTm/sBEq5Rbq5qwRoq+w4b2feougE94ssit5Hp7llAyy
aZaenwPf8CBJS0f4HzzLe/BbW33dNNxmI8C409XqWs73Whac0js5+3j0wGTrggZD
uC4ZCMebJycdObriOkHPaDkoAEZDJ0l3kH+YBn/QmlkXTHnblNTWQORS7pX/Gizz
Nr6vW/BP8JSPt3Mvsqz0hqVnPZbMTRavPs5s3h3mjM8hrUbXbUpFEwWntTmjPIJg
oNiI1S3V+HKAROkHrGPRDWYTLAguonSMGOMC33nBw3KbnbGtbDtSEyx+TLk2izEK
J3mJWl3KwfVEboeVJPy6YHGt7l/ZAk/vTZO4AzOu5B/XX2W91Y6Icz3d7wix8OFJ
RAAFTix2vlUlYc6m42TTdLVNL5ueJSboRnbPocUgCt2xdzdgKd9rUj2eB1a+1MpT
KYPDhMOe6BaLgPwP85q/A28Jf/Vcyjz2WtNyXB7EaVCs7N7B/iMaKgObFZdHTjAm
LtbcD4YsF9nspAhq/+kdAkJyqtR1e2AsRXotQmG9Dvb3QrzAL3dngkx7FY3xlxkK
49v+Dg7MlKg/iJkSVVKvHwjNeP9sZooeHnanYwf+qLPK2HypJMg/gdXyr2aAPdAQ
URK8y0Lmkt6MqOCepP+SaQrP/i/HN7VvJBjQPdIxPq5U9eWT5kIdthl10l7H8zjv
wcn11qdmQyIn6QKH1j8N2tmjB64Mz/4sZU4fRU1iGt0m0tYT5wdStOiSxvmmkszc
8OH5cD4ozrFHDDoxumoDnPQSEzAZ3OU6gUsB6hDs+5xLnJ2ktWA1z5JqCjImtf7D
A/WSrVSc1utHeBuCNaCtsYBfQeY7UL3rElCgNLynVF0q1ffVmNKHbZT3BnX600eU
mbMZt9hLdtpqkTyoW8h48ffpvTU6pim5SvT+b+w4uNkNlVKhPGYcsi5fqN63FgcT
j7gSOCZ+4fExjxprSniXGijVLBEwoax48cLyhj669JXDR276PFScXmWfHjJ0auRz
Q4Du8ElBkbbjs4Aw1wicn5BUGxuqFD1feARt4zSLD31PgeENJuuU7ESrwb1cAG+Q
tqIF1hEGRnTtl/BAmsj0YNOfW1tmrHRwrCu1wvqjmH7Yg45c2mcjkAC3HYw12T75
PDJredpv+vwoEj/HXMEFFIDjxhwzR4dx4vTq3uOvywTlRhNFyIZX8Ki5mr5YVcqj
iVKZD2DBmzTjaHiGxuNAfW5zNlTnNWF09wAJEHDeM/rbYq4RWPvXFIML+QMlhem4
aTf3bmvFEO8pEQ7YfKkM0rqeuOu4OQAd4vOlRKPtR8uM0OYhHvnqwRp8VhR67J1M
3eIhRHB+cUe8HOcx6rsg46nC4mItQWbWeR7B7qoowicA/DCJcIyTZvQEJcYabgY/
c6xHztinygLjGyq18L8nEmjCmmsToBmiq4vChqSppYHJ8xf0FYnWbi0dTqO7nnMb
LSNu3EmH9J4fm9ko4WVuEstybAMP+kIRFXcbu388FuRaWtpIKOjFyd1kUQUCdLvq
c+bLmg4DI6mzVYTFjFRsAbnbsiqOML3McGdeZjQWhciIdiHmc6LfiQzzfbF1Fdwe
ULU1a1gLmtzukp0BLcM+OQIYwdhljQRvQD3nYGLjbZtZ8WAFywk3K6edkZR4aNOa
96IvAFWd4BbGYugO/fQ57mpc3HVZDr1GzTcIKRNYP61LAdaCK+dQWy75j7osEv12
NhL2gXesQNXfQ/FwrK/c2fsb81X+qQJDBgaN9VBOaPhf+M5A4YhzETVa9pVyVRL2
AhYEjRZmBZ70EJUFB17/pv2V9N8Js2zobmdvtFSB4a74Fz9tqnfS5XLMyrOnp6Ji
oazPUKsos+Vbc7NkluhH1xhym/VhJZvthypxyx979ZshV7cBfHSR1sSj7j+yIuT8
s1ZoXAprnSG5+oGLCPiLNgk4chymlaeuPtfTNKBqHzDa9bnjIoZbp87gvGWybQsd
nNZCBvp+rV8FDzeghADImz8EEahtbVjGiWwqV9WGFad2Q1Yj9ar+VVgT7B93UFyI
+r54r43egbZ5I+gjC7iB0slDBhmENHiPUMHGpnQjE5P/UJ8S/AuISVSuLrf5Eohj
wYMHQkHnugX+KVC/YpOAR+ftQdmzHmbYsJ+fpBz3Xa/9lz9j3iqaNFyOyaD7Em0l
qFX/LBM+JGsgN8S0HtwhJ3+zjgzuF2FvI6wZIXXLgrLF4s4trEe5P5xldJZQfmQe
69c/L11xi2hmk5Wv7tgq4DiJauk928UDVwJw9SsOZp6HOduAu8gpUhfn8FqquCIh
BgnkXxgtNv0VnjXbIISDul38pY2e/avJsiqTo6/d4RXOebX5xAzGcq/wtzY7DO5t
IQ0k9eTTAgLjWKBZ9IgkPXpmprGh9CgOfycWM4cs5Uiqv7ybra+fN9gYhB1p7LxR
kttDCR8eYN5cY/A26ZYmsdu8e9ozM47e339X3AXLkuuqD5K7K50EcG44qmmat45/
vE7Md06vHa7ctFeBrZhFencrF9JPdnWg1t0DMq7XHCkSl9prV2lWhc5TpLAhRQtP
PFuUDLzaEuNQVLMp2nhRMHHDSXTrOGT0nTVhc766Z75XDbqbP2ueHITAc2hqecVl
SMpUMipOXyIWeFhdX/SKrab23ihZiiW17j2MocipcDoKeFRraT7AcdbIlNH0hldm
qG2XZKv5ZyoIfJmQbFV7gb4oJ7PiWaJRB4cHImixtUj21N5heagEafyhO0cyVtHm
6qH7iQysOFoauSmmKqAfhg6fSjLfJqQS58ASMTnkydg6RMTR9Tb4yXb8KY7e0O0F
S8HIOQcvDbUG+XJCU1ZCkwiNXBc3Dl+u+oS5WzvXjS8DZOYPKG0c2PmuwZT4JZFl
O1BrlQDfFh2oBloGepNTwTc5kPy2ovUtAV9OHWBQ0/Em+IbCuWlOUWpzj8DWl81X
ZvHPS8ajIE17Bs5KKJ9c6i3yg6bI+TDTAIdpLhTgZf0dlFMr8KhC8+WAVrsrGSra
HKmQiFF/2NTh3F5iArHnzpy+kjHuo7Z2e1tFNUAPFBnizSEUpZjpiZgsQOv4HVoj
MgyJJTU3pMb1tSRaxPP+KhupeC4BqKe3XatocHlYPdfmCJ9XitsJLNDg4XbMo38z
pO6xHTXhlyTQa9WIpm3f7ezIkhj3V3qDoxjOeYjG4N9Qw55ca8cG0RXiQ5LH7pxQ
nROzWW71PqUhNA23QsTPxUFp5ea85D9f4PLnTW8Rq1725+CJMrpCH0VgYfq4Ydc/
Mak78Ad2jWR+s76Ga4F/QKvhqOpsgp0kQefTxMZ7HfiAaYaUrG4rnpsOHkB1dcWq
VMW7+97GcMV4fTm2QBXSd0A6DIGh48ZERS/ux2rw9awnPpHcmos66Uy1EniB7Qif
FnORVV2K6mk4T5AxmdScNGmRwVk/cR6sZrcFDhVn+hp8cK6B9FiSkHR0V15DotWx
q4sxof92blH0Z1FCfDTI1BuXN7k+OvCpsgllzhXcPat5V6gMj+OjUR2Z1GHWUC+x
92DT074m3Yk+7ldqyT20+WpVEYDIFwMu9oBrqlt8f1WWqC3Nq0HcyworO9aLP9lJ
+rtq8XZHkLa/JfwRKoQK+4ikb24STyzgtwp7RLLpgJX96YIKE8x742U6P/HYrwNP
HumCKoWYf8X9lQ8ifUPEIn6h9LewGKZok1hAG6JdmsVE3ziCMepWlYSLWFtJ2xZI
+J/UERe8XebEYUsKYvE4PedXFRejB3RTsGqCPIVDfRkEMHXl1uPx2eXHfTNqQ+qn
X3+wwV1AGmPpxwuBn34jY4TJeV8cIN1PB9VtpXBWQGemeE7OHd/vqfafWDyKfVuT
UyioftF0oknyXDG5Rvs4N1cDvPhOLUnwA0l2UUtnV7jGjT4pwjbdoGVui/OuBCsg
ewbVkFh9z4BoJOWYyJUjiTOzJk/jiw3PhXoW7nqZn4GH0ZIkX2UeGW8TOGUZtk4A
Th+w6NhdoSparlm747n0Fg7RVMwNq+VM2iMflWsEB5WYARQrUTQOegCRLvnOY5pJ
Ka+H420BclocQBn0WsD+Qcm2auOUltPtFTHGMLf6UKZGBQMyBm31eFWhq3lXVb1u
x9WQLoLikalS1s77HmRlkISzoa8mSdp4PFYcarx4YWD6v9VxljI1DupMxnfTugyy
09wWnEGDHgF8bbVzBs+vODp3rGKfYuf0IttvDm+MCXe/kdBytaehxOiJNBQCDvIC
Ya3MKObUxtLl54kJlDjtjflCJ+RHqOKa7NEZ2amhUjherXV9HSI9lAaohk68Hl8x
9TlT8IL4TL2O5Y6GeRxGmiVG28LZLxFDv9dQ26tctNlcZlQ5NJGGMoEs9ZoDSgnv
R4ApHFuh+IWIoFGReMIi7wuQSmU+8TV2NeJXjHkXBTc78+aGq1YbjQQD6hin+QZ1
+mq+Mr2PRGgkP+IKc7KvatHX/ykc6wRuWhN7XzenDbyRQmpyiEFGZgtt6HknJ3Pz
hjbTGeXIOWmLH+j+l2q9WMYN593pZfnq5jYpGX6m6jfvYEs5HqIx3gz7ynOqBu6L
anjW3tJuJ4cR3gjMvnAm8s49bJhRWa6OwbL2Dv+x02ZGFRRn3Bqr/ZwXUjMn0Ywc
6/YzOh0c0TNEMhjAs1tWfhYpS2Y6H9jYZwqEpG4dSGRrib9UZ8tEGhVurmXDPcK4
CjnYORiUToOHItKnVIQPv980PXQAU8YJClgRkpYBAQ7rfZXdt9y6jD/9/JS1zV6c
wW1fx23YRG3AgWj2+50UMN1eKFGy2ttK/2NwKdEMjZ+U33HRECLFzl0FBYRjGmAq
YFiOAg43w7eSSVfr+DTrdusgTGLtSBNtlFYEeN0DyI6SZgr4zclTXkNZ+DiS4HC8
UdpwDToePrPGdbNflOQOihILirAlKovwz22R6NY+SXSKPFkhUgTNt4Cssg+QxRaX
RaRd0as/4/7Z4+9tEetdhl11p96oN24eKtyolLE8iHMd1DnVP43Ue9/OrslNjh/w
Ha430OzTEfUaZUcaFervg7W2QBwOoz8Ig9QgQrojeQWdJKGGaOHdXiKiMS0uwKjl
MisNz51qhSKEuFEBg1tUTevifTc3sQSsUbSBxwocrlyQT8XoUFZZxlNsrLT87DMO
yjWd0w3rhFLgzrykBOvMfQDF1n7C4QyQJtpnaUpOvBFOw2QURtgtwWawRpzqOk8H
dDdLnTgPzJ68VEQtg0AmUn1Z4S8O8footyzNT65E0LI11CiPp2I2Xmo7xX29naZf
McbM+1o27qRws+9Uj+AkDZVHduBFYVNuW62w7Jf3HEJXVYzhtl+zQyH+qAeQjQYz
8InZzG1IuIW59Y6CBqTd2Iks9DWDWKONfXXqeTERAsJMDAxmYujLoPVJEN7Xa8Zw
cE3KhBZiQ/kdlrK9fWGWZjmSzHBa1ch29ggFP8FzyxvkWh/qjoEAT4cFMXVrQAzG
U4Ctpoe4h2XWHK2NmTo7bGnkHE4f8XuWa4FX69jZ38/vSY5gdzHLKxLCgnaKr6S6
3PeMhJa6oSokvo3W+FiRkbRxYX1xsX46ZP/eOaq+cL6Tmw+7wwyTg7TbySl8hClT
mtsI1w8t7/75LcRohuRCrwQ1K4q+6yr9D30OscbXfGqsU5HHVzWnj4aOm7a/P+zn
PlAVOv75a5GRsw0vEjq6e3Lk0D3tjtjwzjyEFb2ZOWzOEvA3NYppXkyFYER1Swpl
7HL30scpl2CFV8cH5Pca01QknjkGi8c2wPCqhCXG5OCkLcq4ZIcS9GaPzeE8uVHm
oLCXIRy9ctbLuLAMsl9sdbvmcPUo9d9IzuWkGasreKANa5241obgVlzfUr6TSCpU
OKDFUVj5FAP0nxH7cRUegot3zhCbSJrEWbMEYI4KI1NkE4z/GpPPg3HcEmLCQVGz
dcXWjpMIOomrq/SrwktFgBfqMrwRrjzMP4qoTvkyw9p9XajbtXig/vDywjdCa489
OemrDOaGlVvEop56hlkiZ+1ksII+hNY1A15Z2n6Fdak8u8vncmSNAeU0qEkPegeu
s2NqBAVqHlZ6W8ryuz1aVITRRYkWayM9SgSK9YxC0UTCKHRRjolqr2wJO49tWqNb
ppZX7P2Hz3f5IG4O0qj6OMdsAlpQC0FiNSBXYCLehcCL0QjYy9FxT228lE3V9hg6
A+tdBi4BxAZ795TxIS1C0Brkqz3MkSjr0geU6cBjY02uc1R90QCfDqD7wlCToWMC
u7j2lV4qBsL2egi4Wy4MGMzisE/uf2V50i8n5XkA+8FzW/nvL5EeFm9SesZfls7z
ds+bV4P9Tit9LnWhbr2MKPkcJnRiVhRnJ7xiiysCOEm9Vy0ftMWXYdMBGMamLy65
LHm/XSmpEo24trqbwXzuhQNkjiaBBSQhbgLjTenXH28DEBfmoaAcdx1OsiuB0gwW
Pumrz9JqtiKRik1BVKNIR8HEGq0gteWMhES0cv0Kurk4NxRSWbh5Akey9WUtRLCg
pMQBsSWr/Wbjdw7ueogtX9xTMqCNkUzDE3rEIInI4Rg1+tGAYEksMfDY8B2RD5Wd
MruVZ2Gu5i/3giOroZ3bTP9CeEzbkGko66/W1QYz9LJShrjiDHLxPsk4IMB/9ged
vNTUuvjYiQS5K3j1424U7gmwEfDVepJ+0D+fRaLKAmIz7ttOxO13DZhYZdRVqvyc
IHNYrH4vFlg/G0VhoQMkhtTHaKX4A3rLupu7ZkiJRav0lczO9RWK9cZWo8Si81RF
ihlYzRr50YbsGvcwvSILjp3xqeBQGY1PQxC8cj5TZ+tMReCROhjSD5DdezjxAo9c
/rON4XX5QfdrIAcD9YsXiTx4+Z5DHJbJHZxBb1dvX2SwGBKdMqGMyNLijMmHXgyW
qGnlHO+mdE1SuM9PO8uuDmQruIjKxW6GcHXL41cxAizqXwxzwhdDxvLsPQtr66RD
/+2MXu+oj+oBWJvOkJhrEZYdZ99mVho6jLa30gWGB3nDOAgxGEd4LJNaTZw9iV5c
UOcVaRiQfMemyrDpU5LMM4fxylvyNQsZjqhPBAi/ntViU3YYu4vxZpQVGL+Qv8ll
5goO4TGoypDeBwSJ+Se8P6EKNniMgbJcR3/wAzGVcYkVhFCOsHGgpHAg0uJSviEH
lbx9TmRhHjjkFJfsD4cZN0wQsWVqDI+8cWRITOpEYcImuefCVuYMLXOocI3+6Xoh
SIU8ZWb8AQJVU6OIfhs3VJJQY2aUnZ+jEHmDn+4lZZ+OE1GxXmcGZuausL6Hq8+F
wrs1T//bvVODPRgFolIRp+E5gX093wmbSp1GHkCCJOl+bWhhO+oo0iHeUswdkrSK
mD2TpJZRN0/n7dqLjfmvSHT+hQtQXgLmEKQeN09v7w1gAc0ijFZpMyQx826DmqPZ
bc4csCUXoaLCdHF/u/Ut5YFARVkoqGzFXHd4TKM44QH7pGqrfR7GmlAj8dfVYYnn
BDP2d8RYQ+1jwv4irTcR5rzBn1KNJ44r25JqKVulzdrZ6c+wggRjI21/C3vwzXK/
KXQATNY+QpgJ0Uq1BdDYKhl0xk3J0VOwZrqUSPQquRuQCIDUB6rCXCkfH0f1nDzm
YuANmqPCttxPj2NoYF4tLq00Bq+b+Az8PbkxyBpnP5iLIEEgnsJlrqql4ffxsGDy
DjZAjdvJc+LnFORStEPQpYXj2pG5VQLqcJbJEcN/6iC9Eewvsl7NTTmrdHgTF2Va
ucb5/U3MvSMBwu9ZSgPawjuboyppfUbIXoNC/pjNjgwtmbnFBD73QwAsB3fEYykI
5xTJJij7FpWhlkUzZCc9k0xWi4gGUzd4a0bU8d06k6YVk3OukIPpw1a+FtjCFTYv
v1/gcXGoqxPvcgIAEseu+w5HTgdhA+9Vw8VkI9X61DQXqgbQDPQGQ7+ohfQ1Jx6+
lauM7J33/AFpfwrOTL4ahT1FZ3fFUNuuqoKYVmAAznQVbLTBG2utXfTlDl+/hacP
M21GkJ24UAQeIAi2um5YNg69CITg6EkRivHB0JEctxjwqbZYP4LCpGGoQj/m9zaS
lWkvmMIAuMjCHCi44VAxCER+s3OUf+3s00Aatn6tcKpaMpRQuDAxvAvWw44ZlHyB
ER/tc0Zi+RvIhBdDoj7S2gSgVg/3SCLcowS1XMuXH6xH46f2Q5kQ1myAF+ZoQ7Vx
u/rSGfBP4o4Kz7QRyTDq0UvifqjPeUmPpPNCo7CiyFzlyXM2tzRaX9UMkER3Yoov
JhP2D17SVJW3L5kQHW5jk7ASEjf6wzYgoauSxA0cqwBmwQKp7JmQMdoyhSOXVWp7
pd25k/QVfnKxAyhX1F8Fzct3M3Y3XVgMQ4GwOa/8VUgvZNGSQ0kC1Tl5bv1SoUcD
z+sbvk40FdFhWvyeKXfShsinwoysyL7+8Dvt/Axkd69qwSYiA8U5cHRJviD71Jo+
MOIolvnrFXoY68M0THa+TGe4w39BkUZ21LWJxG1BbiqionVrMTFuYImZ3U7B21BA
PfhB0dbOPVEG96ywcNZ7MP/p6Ufn6PQI/ntdKAAdSuKPP+1qdnSksRCNXwJfAIvS
CeRsmXVOmBUPc58tcdfreAf6E3ncMarePcChli8Y7f4AXS7l2LrsE5rbs069X14/
zBoaX1gDtCP3/4iwEcUe9w4C9nQdSrXMLLRNbNjiYclzYeYn/RmYoIi0gNetSmlx
6mSt8oyaNbv3d3PoG9Ka5gJaeuGZRZXK8G4tmC3tMclVc5YW24vCKCxHN4SRjS+c
JfCb+gup+Y1CGeG/+oUC82Tzt/fbhndi/wDotuFn/uGpkeklUo5UmzNvNUFMV7K/
r7lmnilgbcePkDw5/rBcKa5WMT+74yi22QSpOMZaKcwb14QH/EN3ij8EFWyw9Wrd
btzLatr6hWOdXwT6tBfDMURh8V3/ntzuSRz/cNXBMfKMYjOUI3WnQWiCWatLQd9J
akOss5c+9advWfjMx3jC9Qbi9/7uZYi77aQ0NlLgS6dB/vV+r83aQs3+kGUqlppr
JzZoeesHW6QkP/ezOjI+iP2taYRsJDMSRLJWN6t3KyIYmTneU6APtoBPo+d2RSK7
u8MNQvmnSF5DTJghXKrprVWdJloMRgN2Ntknj4zNI0tNjAik/6zhls+QrwmKUfG1
Y/zjHk+8DeZWh7jjHgFDjryVeHawhEGkV1XN3pRp6rJEc+kBw5xeaXWfCdGr4O95
RQvnycsdfQZsPumPGNge7CMQKf+qtUHgHjzZwo+OYcX8lvciofaVW0Bx8LrNIGAi
kW5P7g/dY73Grj8ALF88GvHvLL/JkiMh2euNrC3WK9uTA0ZJ7i6pvj3rv/lnqQuc
+qJFQj47LSKdGgakOBqroGrMPIWuormNVVQ4LHwnrevp9eEFb4tjzmNlE6qNwf00
p/8XQQArKXBRxSFi+t9yZHb5/BRmqO5OIkkvIV/Hh6oyocO7DoOG2OjB2AnAOCdF
KMxTUSEngDvul9CgMiNu1T9aBMn/MKYq7Q7zSuNg/uqkP6nPXMs1jVtJqS72EtOp
sjO5VuzTYIYs1dYcCLtsIpKK+gBSnXbePgcb/hc2VZEOS38/ARhTE7PKZpQSrkj3
AfeYrD61yYkAEle6d1GAlE7kAPhjM+zJbDBRYbjUle8r88Q5Oo5OtS77pc1QMy3K
yo6kmrHz2LDUzdLA5lw2Z3GUewUjDeoTgZqDhdt9e9l2z4AgRJsFRt88vU6jZoRO
5qMPiS7CU/Z58tNhd6y/pMR/kUckoaCv2ZIkqgTMG7UUp/fttuGBwNEKQYEUc6FZ
zB1HQtlxL+qKnzR+qnaoySQPpv3ifrel/WiK6cjFuk73MutB0rtjtbq2WRRqtP0o
In5O3VY7Izdd8CF/AFnSEafk0eHLw2HGGot9C+SYpVDCD0NduzBP5uXejFn7Xvt2
NYpqGmOOWSgyeAXDJi/3EvLhKYfQD54Q+BGpsPanjVV7LGArOQ80s2MRrqGdUdOd
t7JmQ7VWD5gGkXES7XDt2X2J4lN1yRQtVNr2yh7vdF2mMqb8c4PiBpdnL1E2qjZL
1m2N9Mj+EUJR67lW61iVmElay5gUunG4TyoXFRyHDs6Z0mnM/2msA+5n0xclPLZS
vC7MItXGAEBAu54PSADo50INE1vOOm02BX6lm6P5UrfmC7Ipvpxq8s89HCox+mag
I0ljs/b36dNJI7yVeJdJNWTrlme3Kt/c+njxx8ipP9t7RzXcrMN+TKzkfbskDMVc
LPXBxf84iv2w9mEFmkcYkU85imFwatbbUFcAcQDuK0+ypwfRssCa5WmqdaR+jEfS
myPtwGcxm+u3dJ3WZMQk6Ae0jKR8BKp2beLkRU3MzsJihimZOUPnJMKJANFYI+kQ
7aGZdwTW6B4yw5LjQrWAN2LMyR8SVGuG7g38294lzVNHeeYJtHXOwzXzFLCz8x+n
OxP+lyCCBtS+1QRccmTbaR17jtG29YYSXQNdyPoaUmdxT1pWDVH7MO5CdEjj2aJ6
vkVLeJ6JF2w3s4xzu0mPlErRbeEOvays4zvlOXdhVgWR+l8xR89lofqKnNWRSfsR
8W6z+uLC7BInm8aT3p1lnxwtn29bW5zqqVNI5uGInMzFskDCMVuoe8NL0wor4x+l
L8VbgJ9srq4I/3bK01ddz9dikJCGC5JA6Rs8P9jMyiX5BitETTb65DNxsWTmZPHD
BZdSqjThVseyEwLmsLUXEpcaXaa9b8vTg0Vdxu5WAOuZZqTuOi+LM6bzqJx/Hlqs
uO5gNbWZaG+SHRgIn7UxeTdXwrHtvUjzgV2OIRHEN2c1YSZWEqO6y1yP09UaTzla
9pmY23uAAqbE9HQT+7F8V6+Bvjd90wmV9+T8EUfrSOaL5RXIwyfsUPlT9Ayh0ckM
Y+BP+xAcHnbz9abG5Gw05kiVnxukwzDlA4y3uhNxOXkIDGcZTlP2cyYYYwdMaypo
krRltrr8uI+kokT7X1oZzFe/fvlxVIoSwqwixLoesamLOaYkdu3lR9K7SMXpaWOY
rNgc0Vy1z6UDulp1qy2rtHr1DcuhSGXU5GsNJD82MGlt4o0wYNILceXKVqQhe99F
tB/uFHe7J9OS5gAzMLcU4HKQXIYfyO5w38wmoq6amlOpZntyNw3KW3B4OdwPwgXQ
Z6YIBXlIJGnqT3BT22FwwdPEZszPWMe847TVcuOk9Dl0CKNpAJ/UaAiAWj9uSpBh
DLf2fjHQ9ElMYyDYxOBZQAfQFK+UMCBBOECkn1r7EMjzqsNO02VoPbD1EFtkx83j
4h7DNL2WqF9/kpu33uV6oaUnnQcnoInQQEkJBn3GvtgFPTaiNEjd4HfUVt02lizm
knv2yWSFXZh27vJaHYhrP5Ad1x8hJRCCK88ELcB/WO7m1f7pIOabqrDjdPfTdj0e
RK6yXHMaQMhHyvdOWV4REn1qLGMz/L4N29+h4FAQNh7fDIIREvu3nCWzszP8TYRI
CXzUe12wtLUPWTCqrJsJBrxwMOjVyD1BDGxg8j4hYvBAE3uE+v5YYiwykYJLKQYf
cxPqUqkDTh5bUVvrpXw1Ffq400IKb/mEQav0LQ0/WbqP0FrIHSMZL7fdglt8zFcV
JRhyx6Ir/N6i6Sxso7EaVNwxDRqTUIsboOlnfzJncxn9YjKmC3Rmw+XDCDc0FBKJ
WF8dPk6Lc5Gs/wXkUHTqq+m33fgS6wKqZjQk6ahfgQPi40T+pkMIZ2L2PITs03d+
eRRf04uaLt9U+QnnrSzuVbX0csjhoz7kp1nFXU3/2awOtBQg57j4lbUDmdzD2j7m
S0c0/3APbsK0tWo1Xskh8SaaP+62QxgPL5tMCn0hFTTC7PqbWHOxeQcdT4uLvXaS
gP4yY0hEOOC1Bhxa5cFXQI3lhPV+cmWHYFsYVxHGub8bY4PX+kDlXZwCgOsR6O8k
I3/XKb4lyDVyKyVY5E949FsRem7IUVxluy+qpuwiqXXuIKkHBVYbcIWqe2GEgnV0
IceCQETNfF7nPX7uCr2Hi9QIC57T/7GT0Xa2ZSN8nv9nV2v3O4TNDIKVNVYxq7KM
Axzl3qrjK3a3K9cSaIB4jKd9llaBqBl1aeOTS02Zkr9ARaRqrSz1raTSlZqVu9gd
xPvP9CItUpGcGXRf79UwKBVdkrz/1dS+X5bgJNFcqtq+YhmvOvAOt654IMi8JAag
yIYMkQAIaQyaej8HV0PTBu3IbolurM66cKbSY2iSeLV/urmvGsqvaTt7bgEqABQJ
mjZVIsaEa2L+xcjFEFfzoapZk0FL2YTXqX6ABwe3W/dPmlaGX6S3R7/yzkW2V2C3
5RQrNIk76sbM2RJ6sKB1d2iAkcHDN6KSewXApvbjzAfn/fJJ/JgPYvunIRxOAVo8
8a3iAtnHmm3feOJC6WXoT2diR5oZx/yedYZq5BY7imiGJ3UOKQscxGyvmbmG6zSl
Tba6qRvI1B2k8I1cMVn+xBPSibPtcKAY0JMY+G5HTNJae3Pn97RgR2bG4AQ43k9D
Nc3rb7Or7q+ElvO0H6T0DmKdQ1g0publlYE6ymJ8Mhy3kKT3iIVhRavgeSL6p8ld
P8EX3+JvRaYjkK8mtjKhbBHHF4cofRCtfFfai8D+YGVWiTu56LF7h4DoSryB+GQw
mRS6mk8LK8PiYRRA9rztJvWknferTxYND7eBMwLuDL7pO8pfSSsUBxhx9KxpsUQk
dQ7dhkkiy5MYcifcbiVjL6BPznQRpPuu0wHKXsalKvPmMN+alLvt32BPCIuZenPA
UknCnE5Gf05sHh0KqO6gh/fzqSuF2hKwBQ1fwV1n76KGlvJw0WjI5N+hzfnlnT9U
SvlhlhPddLvIQoISVLn0HmLDIs0EnJSvoGAujHarR/t7vPiYtzccHk7HUCHJ57I8
7Qcrn9CTHHXJzFLo/RMkzZyY2Hybwued6mh9dBsC1EOQj6cQP4TYS6BYIA7oUXXq
U9xIJpdFYO215Fgx0SXFrIbXplNSLxuNPqs12FxPCWMXprRWM0O7IsYPg3YLhVgq
YDZFtDwbLL38qwbXIm23u/cTLevJniI1+U3uCrT/vBiiTBBWnzVPRP92D0AP2KJo
Nx3B2bpVoD6C+/vdExfSJ2y5vBUzBVuqq5jio5Gnbt3kRjszTbdsyZJM02co01Pm
B3eoJzGYGCZ1UT2OHaj15aiOVXAhhhlBGd8T0saev/kGtpVw+xsHhfkel68fFDN2
bupHBxt8Qrmbqrjmy2sIjALs/wwobOOCzjcF08JQOnhM4iTf42lxVer/6+I+Pxmc
ci/ERVRVuNfRQRoIDNFt+N8aAQYAzLmR/KV2ateb/JgudJHFWrn0rr1Do5ROCkvD
ZVBOCifhIgZs0rCgIUXbv9fR9/n9hZmTpVA3G4HxfhBi1bPfYMd1kX72dJuth5Cz
94ItxXwtm2YFEJ63MoTX7Asgn52twuwcJpJd3/xptS8t0THXOB2JpjCQ6pRHUHl/
cYLjZsV7E7XEBrDk/S6QIx3cEQQ4I3CwGca6aEU5TJIdi/T04tGivbaR9Dvlvvka
aGr9lp1Dh878s5qxoF7ZWF3+skWmyUxSlwxwwD5e+Yz4ohwFxL4b2T34em5qsLPE
LeOEHZ4u/EI0/Q0QrJXoIIEY8wYDiJ4AB+/GUrR4UKvryzER6+76NoKW9N/AMjFD
PjAcPAQmk31C7zIyQzzkbb5/thjV+rgNcoDxbdfwbzyqgGhuZm5tbHKodVZEIPPV
JO3sJAK99v0ZEheyVgZgFFXpBcIcg/8F3aKlf4pqiK2aKHb6VY/O5+4B8sxE8F3R
H4Zn48sLzqFG+NmjJ/zJWQGfVaJpt1pc72VNM9ZF7LH7oo9c3vqAo8RAWaxlhf5M
pglWSybwE1466MaVv7uKt/LdLb9ZILw6+XDC8EeT2pLY/CEeKF5s1FJS5UvotJd4
nFboL7b+W9psUMErpk2gUwkGXNWlrG/QkgTLy1mIhx+wop5vGiFvFCUXW8gFNBEL
6F5EUOXmex2rHt667xLxrusxlZMeDk25K+aHCLIaInBf2uSRxWZM9pFVfOmjS/Da
jwYXuf/KZ6FNILAFquWIAU1kg65Lf4K93V90ggtqS3BtowgPhyAL/aNu3lRLpQ2g
BoirMkIRmqPf4blJz1hrJzOYD5MEggejYLWCjwhNF52h1eJ1tLVqEC/vuNaGHY+P
J6tn6gVDARaLUX/U70fi9xlZyd6choNHepfdlHXZwj3Nk0e74hRuo+mBhVH6P7P3
sVfYS0+73QxHX+XzdlX4KnZVVjf9Lzszb/VB833DwRfmQTibBNHHQmWIYZ7mtSVL
yh3jUsOHkF//AWkJgFzi5/myqftGPIMjkGA0aHFpcgt6ASRtyXEbJW4k1M/0EQ3D
Ad5MVoMUUX1QQl/sVdqJVmdU7Yi0q893Lx37buixH0VW7qhD//xeR8PbhvOH4x2W
l2EodeXxPA0B5uKuOrZ/5QtSs00s90o50icOjbHs4ZD04zCtjWzcZb7A+6kB/qH2
ZHTLXTBo/t7BcUsJcO+zmgeUwVLbHicbzBov25QDtxSMTxvvldAZjwjG6YkALnfm
jFnUnr5+I33pimtfNpvqVPHZEQaFq4S10ExlzT99wqlKSNEDuMbdzdHIJvIrTzm4
ixHZ6GYnWR5W5v2aWMN9frQjmEJP3iWxD8wiq/y3njo77O+IKu+/xbhONbRvHXX4
JZVZW/jpfRG+QSgA+SmoMWg+qhzJR2sDu03AAh8HBoojBbhB/jzT39Zum4IWtPse
MmSzrBzCvuYcCOWIuZ6jGb+OiVPM1DKEi5qulz8TYrElQVRU8JTrCq8uk06TrvE+
tAiw5cHHANtwZqITleYYqWOGUxwdESdio5zP+Ykw8FKapcbeA3ah63EsxUqdrA9H
1wsReZvdyadTivp7PYSQSMVU0xYPjK9QG6zuJC2O11aJnZjmcco1kHpkDAybvEx0
+7ewiemZXLd8Oj4emsCQXrs9vcOkPr4iFd29Du1nih5mhuvTx5V6E+bY/DhSHBXZ
khEKTzAdZ34odCwt+IGZq3eDK4VfJJ14vryEx661E2VZn0EX0ZDdsYWiz3fx6gyu
fFl2s5Q/yFS68V1n4Yt9likxzPf3SXC/z/HTOGkknLWXcKoCD2XRLYtWD21IHAtc
DTOWQA/+Kjxfe4awogtVK8RJ7GCAEWQfHWG3mOpBIpcy5iklIt1FUkp1bzL4zJ9t
fLDg6kMH7xze/RMomWsZ7sdqo7A0SLXXfKh4Em89k0kOgd+Git3XR69VyPcXpfEg
1fR7Aqr7oyU/4/qRfnziWrbB6atC3Zw0FQIpsS/G5J2bpmDk+w04ROIdkuGCUZoQ
+89TAmnawk4+XItVdka6ue5VMgpWPzc2YUTQk1oKHbla0TjLAp1NW9ThvnU3uW/x
/r9csEYLMyi+Ha2XeYZZ8V5Aijlafs+J3jImEk61LqWl4yAYJj7ljX1MMRcthlWy
GXU4jL6yD6smNw2nY6j7mJg5lKpdJMikohZmGlBBjU8VFGpZXUJKP3b7SKT5oKAy
8amquu7lDUhhWFbgRETs8ZllaBRTlJ6ECdBMjjNgRTNKO6NinAUGWhWsaK5XIvab
lhTPdfOH0R+pmij670NKDEDbevKv+ZWNUJ17tiMQ4wM4lRp9OsqMcEfwr5dAoSsN
fUxpxtmhJrA/jQuHbOzjOpEiDvpPjgc5hXxBFz/222QtS0KueRKT6cIFFnqB7rFd
JmhmbPzf2iQkYdiEBqf2PlSmSSs8iD109KT9Ik6E52NpwBaas9TM/NiUXFm9JUxg
288HzfM9on4oa+pNjRsoLAKBIq5Rq/yrjjrMg+slY2cfqQ+vm7yFNbf60HbKLUZH
JYMG4LDr8ZMWxvdDnQ4ruwSW0tBfRElzCoengb7lI8tBWpBlxw3PYEcz0ZAaLTIj
vVwqLC+GRDwdEyx/3g61Cvp1D0PoR1v37PQrmc8B/Lq8ceWJ5Pp34xon3EloZjB6
B6Or8NfjOuBuNe8b4hiW3vrXSWFRxfVxYs8E8gd9zqENCKJUm+6/N46o+XKNUqVr
DZ6SjgEY9C5O3Ba5BsgvgwHaRl8Vlr7D9q41en8nGL6rHzMnDTuuJE9p3aEyqvuW
5y8ahFOFe8u3S7FA6cT0dacITMCeOblS/NadcQgJ/gL1caD59S7+/bUeGx0F6v+t
Kfm7IBV7EipLRebAHpyNge7MaJL2ovnjF1kLetjlF2FGcwhAGL7A09Cl34TJaBGi
2ipz3AGClG9ljPWJz6O2lEofxZTpWWXoWOjsVWA+ciWzbc6Zlf7DKB/3P6+uHlJu
ROZNNfe40dmpbR93lvLXQ3S/rWgdFg+mt+lgshk0b4pYs+lQmUYN6tYkeWwj0F0a
19w7seUlI3CXoTAAvSw9cNuAV3ZwEupnnP/NS6YBqlq79M5dOo0qhXbGJAKa3SRC
7kD6tgAuDQTUAjrI6ai7pI2mQuAGDRJrNiPeLkAAnQLEmKsJ1VlZv6PhI84PHKE+
1HQr6QPThD6dTJ3BygjqVzOxfJ7D1/XURyc8jZhxWqX7hakpFRZOgCq3Z2WIxsDt
n+0klw8Ss9xYoXp0xQpHESBVm0Zj9ks6vVyRGnrHMoZw+DscJ15nYr0oj5opdnsL
0QyeF6K4Gs9svKfY5xWJJ7PM8MxXQBNjrWDH88CLrmLHQLqmdaEQ9yYOCDnSJsd7
AuPGMm6Ff1JbyXzyFzkDYBQjK6Dt9tFXBginrKQTGSNY0qXtvUVgZB0nHYtCSQIx
dysM1ZUjypr3ZzmhnlSaxCucUNlTkbNigEnVEHAQAkfs+4RY1nnwk0/Yu//bQga2
JRiHLcrYoe2IgUzqNpOZjneD8qL/hc18iVb7rxVnXX33XJdxtUUga79d+Vhl1L0M
LTuI0f3gQmL2JZKdvjYCnrauzqKMKX8Wyw8rZEXtWcvFcHHAUZt4gvUpHmAixH3i
SrdNmvyBRBXkBxHfVJWgRKjZZ93QL4msWHCGHptY1fULBlapYQopFgmzdkf0Yopk
WqZhywBSESt777SNrSqGzOvjKoKYaC/TomVEfp1Eqj9X/xs8Iu+uPYUWh/CQulbe
YHOWIYiGJIdtd7h97YDMtEzvwq0ljdGAPH7RFteUgC1u/lh9LkC/6JTWRR0dwLkx
I+wnFAqK32n01Mg8PwbbXPbj37teUlILMP3kr6SZ0ChRbaHaf9W69fBTRkqCIwqm
WqBPVXGzQ9YgfhkD61O07MuQu0PVYu7FZRMzhzhIroRjG+WxMzrwFRkh4lJERPip
e1YGAHKk3JrinOFBcyYUDLu7GltBwo1T9dgm+cNZYkNhBMsjJ5HqCJD4Cn96QjIq
/BF8p7yR9e8WxHNL1IuxdWkecownlPKsOKQ+EH2xOCJx1i7tAN3c14PveGD4rAvR
y8bXm1HJcb6Wu0kYMyiKgm7IaDESesks9yOE8ifexTEq57cbZAm3tNW09l/x1gnN
GaLpVUjFynNxReCA9LajdPePb5aANgSFe23FXJo4UC3MlNINxD1QB+CQpZ938pBs
a/3DfICixxgEvsVl9nnQaj1DJJs5wfLaw+5LKVYhpfQRXCc/ki1YzIneMm2O5Qrk
PNlkk3fc0E7wOAxi6VN80un+0dTDClta0jpwrCRRX+pXvJXYU0wJtoK2s8ykuPMZ
KH4g74haf6NVh9iAp8swYFCIPUKvaD6j4Pkz+FQLNXN01ExxnoxDQ02qjx5vow3S
644MbfARfywhte+UzPLLBjNOTJFCOZwwFLXZcV9bgH3GfLbnyeYveqaEvPGrplP7
Kay363HSqR05z+DAe5pxsr0YPcTV1tWtCopNkJMKkoXbMYyRrv9ES2U29o8n5A7A
LK6lK+BUBBKVh3mUmcMktdpFWC8mc/cwFmwZaeIRGINjgNztuRRMaYM8qjbpYC28
qCULWYQKer4v3eifFdY6QvHHL5VwFlmbCph/3chLZehPCiRgf//L2hwTwBfTCoQ7
CZVW7U4+w09gFpEHU5+Njvoca4/SeyxYEo3kXpZ4jb1fSs78eDyoVRXm8yq13ka5
iwDXrP23szCBMmvhXE9n5EDXpAvNPorPmnYxle+6dxoaU8GBt68bq314+XcmLSu6
26XMGKk35agyllI3xZa8Pau8uvBThFmZe1g1KgJzzVEGG2ANQy+TKlJGicbGOCGy
U0MkxQGJzZUEETYtahlxoKR87S9IPA8oroHL0XnRmnsOpSSmD3CKMIWgwwxvX38Y
RysaTax4fb7MOp1SNgGTCvkkZBYcZF6tOG7E22d3f3hkVOAaB/y6mPnr+4XDDlVk
40IAHK56a7+Actc3Y85Ed/MfVBykL1AzowFPkQqzXfjSwLSzk6UI/cLeFpzsTev/
APB1iJdHtNxFUk2uhFrNxAmV2U7EGY+2uhXXc8deLC12aikn4yZqQgJ8SsogG01w
oS9NqO4Dk6Y6L7GsYgim9CWn17ylizuq+56ZhrxGMwY+KD7ZylxufzCAEWg7kDGT
Rbub8zPLmOCbyPSkyg67zQ7Tkln59FTUTI+y5pOrzXQOn9RUDPrtCr6zaSdUxlFl
odO3ZJMiD7TrYadpzzIQQ+jgwSJHUUE7YVpD337JXSYeKsEYd6jGel6sy9tUWmM+
C/1wVkQiNmbFiwD26IWBCt2leGTCoKB9DDsNgyy7fvIOxZK5pAwPPG/uivA51oon
73YUVn9A3zLN782b0M6qcLgJMKtMRRlP+XzQpKj6f0FhGOfsGGYA1zoRBNdoQdIR
Tjp1fcdR0USdhxckW7joOGyibA3igiBX0zGq3JUoBOayIo2fSSgpmpLqCDj6sDhu
Wdd3HaHntV00QZW0xgkOUZHoA9fs53mnY2Xq2wtM2pHcUfijBo5YtLRsQmeYTo+I
ksWAhO+0nquc7ou4uYCw/RzuYkvoAZgPnLn/qEnumW7Na3xc2/EmThDSY+JIw0IP
m7iSeRQtZzoqBRKxXYQp+xVo+B9VIEkPskCUfEVLCpb+Vj/k7pQ1YNAX+y5rD0Gw
QlAChp3GcfbK/M6d6df1AltKipvTfD6TPkoZoCg4XBd2imXSbKxGzwNuFcHoc9zG
Jz6YB3PLLxklvCVYv16kPzUBvbKQgelC+MEmEPUuPzprSLs9NPnD1xUeGTy+in5a
BjEOwHtYQM0eJ5tpKml7hCwRQgSf3oyHHEgIZA2f5YoC9B2QWP5j4ySHCjHWmEwW
mcnXpwRJ6iH/nWWJpegH4Fm9Yabh8FDz+Yz20zRBI310xKoZX4EZSRxxeT2jhc9G
ZbkuJbrCqZNqPQfEwzKUcejn8uk737Wqqrgf4l6AuIkuIRaNN8BS1LWUhtQpF10G
9WHFqT1wGMpLWM2geOQZgWOO6fICauRaJKvNSAlqNVLSahsCikF/STZ+ElnTGBzV
8WHNXtYHgplHeZb7wATcC9yncwX1gQhTAC0WOeCXgz9VeDdAU5NPg0SeIQ4dG4ks
1ZzU/e8f/BdvdlsF7F3KyZnLo06CLGNAhEXBOZPE+FVzrwCiKxeX2kDiTcnXn+DV
kygVj32qBVga/v+lEI2XH5vaJm+1KC9239O9NjlrniA/ndwajbvi5YRfSkDBjIe4
nbhuZVg/CT/1zZpMssHdXxthU2wR9amjfPgKoEQxYBKnALhmo9YwbZwQiQw8HMCx
hHvrPNGPuZkKdH258rUL5iuP5J5CvPeNkaFjKWvefVwyUU8sDGheDeYWsIeWAJbm
474V5mW1jMLjXvSPjN14gtDlzkCzEootlm041lCmuiygnuuBX+P2nmIT2TpqqYbT
JAPI3vhwb07GOKb6dQz2YZlwFmYQpBX3aFz4mtBwXE5Qah0yjf/a8K78cHy06KaE
0pF0HUfZsiJtADJF8eM9PvPI0hWq4tbEvAX9+2sHPd+CuYm2LgmHhsO449bXQhvR
e9dnCGwM0erolB8SI3tMFBEV3TliZVUF3bMUtiAUk+kY7rcTwwbHTk59Jje1BRce
U+sNl4K+GL4EHxN91ANuqQjNvdM3E46bQXuiQT/iBZvceVgaotwWrzNK+3S0QJfL
QnlyMQqvo5/8a6YVxalDOxzLXPPNDbx5MAicFO7qEAibTmL5X/lHtNPWaBWjQ6G8
w7s4PW2009emZx+HZ+1F5xxKriIF6ThS0iaRWbXXygOwY2Jz0zcFn4tAH4OcIFMp
cSOVOkmeGu5FjS0xzQTE19hMKbE1Luz5uzE4i+kS+5YeHadpQbP6MqRCkOEvQ35Z
Izx0z9YjwMr9aWiCuTh6WyM+MstPGJh4CbRUlY7RUqy04pjU9l+D1kmNLzLU97bs
Ey1g0YBiFEE9ls0bFKwZUFsyz8z9LHrPiT9y4EqfFltpbrsSO9WxFeJOnCU1/5w4
kOoaj/dYzpA4IxadC3vB+m2nR/70gRl5+2DlmsMfGzSiSHq4a/fnodG/D6Z/dkkS
eulqjiPAOHoyH/AHiQKg7W+njqg8aOoA7ZLnooyCnG460h29juuPuHv0PVHSl3gB
eT235UX6t2Vp1KBEmtwBQXSaKQy/yAnlUAiyPITcQGicp4zmQPjZocSnyMpHan9l
8pp5fhc2QfBDbP9lNJiOY+nSnflye+2mYz//iIIr1YhgFRnYmRSp9uvDPvO5y/pB
W91h3SAj4zBcOuSthqqNXrwfAV1yCHZInNSUSAiFUyh28XzJZ/pnG05sMRkjgIh2
v/X2Lk/hM08VNEhZdXeVby9bKS2KjT+zEu4Mr2bUhiaKEy5d/6Phoog5TLMJpHkr
fUnQvwynaMAAvO2P8yrhEhSrW8I77/JOWen7FQ12s9SqW3Qlc/rx9nr+dks7266C
AtOwtF/V8+IVuHSO+sk7l9H+R3Ajy7P7qQWG/KlAMNtWuV3PECs3FKbdXaNT8y13
WqizG9mnhRDruPk4pNIkUmbiQ29r3elfkV+EAmf0bXV+44MgXsNavpyokNyxaatW
PAjY0KNuhp2X3ibs9hRHEkE3bDfU37MlZEvldjoDz0uHf0kpE3qJldE+Bw3Ixq+O
RQpI40DI9hLwZafPU7tLQgDQsbmrw5zaU1uFiS9PBtawYUI/RTiQT8fnq+QveAm8
z8NpUDSSDehBvwb8e42fYcwe5xajdbCXJoqXdiY82XONMLQHu43udOWhFvrE7j/b
Qe+bqxtTxggsd+zklcUrw071jatItoxK122lYwbYCf2/fDSfocORy3abzQ/uo8Ml
9r6sFe2qr9nulyv3KlavS850gfspO64OcpPHWE8Gin+6pU/X/39LBppzYyGzYvZ3
cMCTviEMcbbUAuEQRXB+PifmnwJzg9JUIoHtDQWQrIZT4Melgm0aJRlVFXQ8HO7q
lliDxFUiO4pOtB48kugbeWnOhyCxTmw+zRp/Wwx1Pxokuy8qEynPO+Qspf+EDruW
6a8CVRF4e3L3WVl0gsX73wh4GNj3cekAOQNVJajFywthy8p+G/s5inCZS+x9lkQx
+Ir8WwcN6Klcy+fIEMtAYpIPdktyw5CsIPC+/4r0HkNYqVyvNhqh5lKYQDsSJ/ou
0G3th9E4bEX/glV284lzItPtGYGe9CX8bBYKEX2q0r2ln7LMwVzH6vfTI6D0fMtj
aK9d6UQOlZ/gfwTf/QntGqTk2Sd5iPiOu/RWNwZlvUhKTVRFzQ/xpzXj4cTm2cJv
xnKfkt9x6XOaXQf7LR3ywNEY/TcTR18LviVHL7UK2nrEr1QzNLmKFkG3E1owzmag
YwZ1ZG9fGF10eaDcXP8f44G6wyRwBQHz6wU/90dgUX2KNtzKV9FUmzatVllJbTK0
tAGGcDKAGHNAJ173ZsXEfIcC+306XxEX5475Hn1MPr6b8ZGyo6vbF7nhaWj6br2Y
Uik6Pqv8hQsIH1BOXUtqoht5JEpgiFNWPkG/LfuLFKexTfETcqliiLUBg4GVygIh
APUzZw5qV1AGYyjoKVwPP6KAyLA7wM00joUVRSz94tgiPGk9YV91Nolni1ITKuG5
CgjIYqDlq2zLqDhMsBGlIAMUCQJAut8J5KVGG3sUDKbzHfdGWjmMW6UYo6quUXmR
Xe4xVTEzq6IpbwZoG0W6DK8SUVh5vtTLCRvGHOx6DmaLQdkk6Ul0uI1lHz9rIgvS
n10xnvZqPtt3CCLu3AhEaQ==
`protect END_PROTECTED
