`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLLNp+qMXfNkQ69O1qye37pNxjkoMQOgYFfsXd6b606s
LUJO7Vx0Qe6LlEl2BEzsScnYVJ/fUb4JKyOk8qzGfYpqQhNbib5ka+WKJgP+nSHc
+7TgiPqpqlpi65nnk6++98Dn3rBhHToyLrZgruCeUu8grKMmLwv9gsBFQui6pPWZ
BTvt5O0wj4aJ+hmfWHf8bQ==
`protect END_PROTECTED
