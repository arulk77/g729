`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46LIDVuQUZ/eTvdw8rPCs5GSzi5JUt39uummyth7r0R+
DWzUp3dgR3ORatAoDThSW/HlecmIVUzv/R2XZwwLn80vefaBgBlErDick8A6Q0YW
1c8YbPrBnU5ueUT7pQkfe/44vxP8Z/eIAbrsXXwt5gTWHs29C8uC2nNg9HBLa7xP
mwMgdUJ6muX/1LhKz/5+zbzJgzHZcFjVbXiunYfJRRoLh37tmJyitcxw7jJslLVv
j7t2zMHo1FJvDxiJDjWFqDj0Y9l+yn9ASS24/JhCa+IYobt5aqzXNRCe4zPZfczT
+/TDNC7KrbPnJYTdaF9N6WKUxkOWw5Y9YpCW3arvfG4j2NsO8EB8scGGIdrtsnH7
t7Qez9+idvtdJCy1v+uTFg==
`protect END_PROTECTED
