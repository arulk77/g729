`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48ZDUsxUU8SEfyT9wFvfXaK7vS2mvRjMnoF8Mx5KihoC
zKoNROLQrmcgyRAfACxI+deDm3JDZ2dVqB9+be8wyqKBbfXO4ridRqWjFdGD9lVb
vFnBYZTXhfM4NmFgIR3SQicQHBCm/pXI/bB2jNRmb0HuZwohAQHQ/EnR5/G5L7Ui
AXJwn4d1XbKxOHmLlRUJP2Sq9Q8IUOPRpdDGVz5DF1Xd7PLYikGGl1togQUOD3tD
ZTqaA65Iz98F8TPJfzdYZMH/0hueRTjMdL+u+4TARzUtZpQ01ygpB4Yqbs8nslUo
omNyoU2gUh5+sflRcF5y7rfSK4D5U+tG7zMUn0qXpN5ARM+1QCy9w9IAF+LO6Wsj
MkDj4Sf6Z90aiuniQOE3KMXbit01R4xJjJ98mA5squDJ8fVQehSLCjYNxGcQb9Gq
q8Htob/A/SjH8tdX9Hn+ChkBWc8l5awKAWVJtoq2uZZvjNLHeC+zRjB0tNYtJrWd
n8J3UlKWQKaTkaBMFZYBQF0DT2AgYN6TtVDTPC7JS8JnxR+N/68XzB+sgME4Jz+j
gJ1+qnoHlAyFWpZhtjOqhi142uD68aQLYmyhm5SFqRzEH3Q2WvbfxN2bnty/tLFP
6zjpy3EpvxG+AeDKuBx0tzcKT2OYDHQ06hJk+YrSiRKD9c1B5I2zKjOlYf3ZGJk7
tuXV5q6pZ41RxNQ2iFXKP2GB6LnWdqKosd6RmO2T1alvmfSvGq+m2nr91XcwONgv
15bDw1IFzKGXp+LlEpRnJoWC9CX0Th8hIxERIsKZjgOWcr+kVT4G0Erq0Q6fexwe
n6wWfd9O4iKdOuIBTEuLWQPIUwTxY672oz4kJ2aobeIWEMQ/OnbE/OkLFZOgLnNu
It4ueyaHx+jpPiOl0oZC/Dweao3j8vOvcTsUTfDu+ezotRrmmSav6DDJEbG/u2yW
egjup4zdLtv3FGRDf3zS0h0xkeTRAP+HWh24nPLYw9PX8SIXaS0vzhISTHvRhCYD
+M3MJ6DEwPTHdcTjrQUbenV7b4MN7L3pf45VpMgBeBL+H+EPcA/qZD8j0/pq0qlS
ZryNV0s99ZDSjZmisT1TE+HTi28Bj0+c6qo8NviB6wOOqhkGSgaJihwCIpb9g3bF
RZs00lgIRPwk3UI9tUD5z+QmVSOxYjXBs3DidW0UOo/0HkSTiu1J3riQZBq6eBsS
YgXbZsjD078TtKAKz0gXgMDOafpVLxQz6v+1V2mIf3mQQCS6Jqpz4C/LcH6JfVLU
8mymxqRzoQnMts64w2lLmbOqpjxjVtW8SWbpcEoqA9uskNmEj+6aoBQ89hYPnq7R
JcfpvQD0M8EDVtLkV560hSPjRBu3PnzfJb14bYUDAtvKuaYlAOktUhfED8JmGWht
qWonq6mtH8DWKzc7WijvT/d8eYJ22DEv19nbinUbUWgDw+LAVVWPN7xtuxn+BamC
Eoc+tpVz3a9+OnylFlfA59aXZHqoMoavNFCfeYHP8zKT9d0krtJ29do1xHbAX/93
R5K3eRXkvwNrCmPggUUM0HdHGSTFFRKVFgodWnEEidhJPiGhdoUbh/t69fkBZiUF
Nz8g+SpNs74I4gcFqSeG3vFKOCGPg3ojvqOQGeGHhAKUL2f3KU1k+0umGagoJEg2
8/L8tiQiyfeYXmRJUsLFsbjyuxY+0qxpAonckS0vrBW6S5qsZoJaanqykIQ8MfHK
zBI3Dy0KJfFm4P301Ea97e1b01UUB3QCbOVXfCn8cXDd0mZjPh3sjQmJZhsSU/xh
iekrVw9ZeZjVWuXIhSYfnbavaO8ppbB5W+DnbbPpjjFloQlBs2RvjFlLb3V5pqyg
shg3L9NoeQl0TEucCgtrBDlQB0W6fSDp4XrzmdwVPzL5SUeJDAopQVCl5qLW92ZM
BaUN877tv40aHtjz2YE6IZ7HkTu31t2tihxBg7ArB0lZQ5Vct9A4XYvrd07CaRIF
SnXTYlv11oSvahbxEBNBd1Y+5kzTR5mmkymXvI5PKERVXD/Bl/SeDfrcxYCkDydf
9cDL6VAkXLxVH8YYRHpovz9fWQ32jkf/vtEl1pRmCpGYM6BHk0ICBFyhaZdm1Ttu
yMBAX72NWlFIFzGetuO1FFY0C61wyU87qrWTPm/ns6IoLzd7g7BgeGWlCPK+jKf5
JE2/uTJ7ZF3PtoknSuqdMqR5A1L/2NgmEBVzL7EyV4Xb7rX3Pwim6cyePko1JENJ
fvBNPxlVbBfZnU0v7Cnzwsbwjop/URfnbLGV5PMVl4tCP8EDWa7vHGRTkuGglHAI
kxg/c5JqLvIvUbAQzEnSIizW+ympl3c7NgoAVrwamlmvnPvXwCCD3YSe5zhcYaMO
R+gE5YQGXHqO91GMsCZbTJsbmXa6n9yvnYuvqDzi04czX4gah3oM9XFAHQvwxu+y
DTo6X4e5tgmsLpnGJUHu8P/LQzlr8osGQ9Zt37/uVzhgTFHu44UDOILgxpdzRivr
CbijBVxHT8jvcRSSSdtqC3GC+U24T6355ms9NQSd7bC5D8oLecXwsvFabpGcIZKo
116eM3orQUCrkXA/pOyVuuErOejcI3jEK2FB9PSKPBC0/z3tADfmLdqMnPm/J6dP
Gzb28Zaf5egS+TlaUhws5TgSMjnOPVGy/SPXDyKtHjg=
`protect END_PROTECTED
