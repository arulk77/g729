`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIK6dF3o5S8xB+THW1JAgebDDGhx+HKx2yxTYOp4tIwd
EDLt7iaB6k977nNijoI6nsIDXC+bEhlwOR+Hm4b97ELQDXs3a2kAY+18rbfNff6e
JyaRjg18XcTupatfmSbljGdpf5p505ZofJQ/X6qEnBzET1GY/2dCCUf+rPuJFyy+
8cf3v64HiV7v4cDhSCZuvw==
`protect END_PROTECTED
