`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFZYhZP1MNeJ/qYN0GI8qvEtPvM4wNL3xPIC2Jf5iOUg
wOL6yf8nibVuBiTyMnPXVfdiASrGFJLdDrrY5rcON+ntXqLTR+z0WZieJ+s7nZOL
OMt866RmVmH9Zj/eS//udShPlYkY9vA9Yq52MqIGelFAskSveI39mTMoeAu0h8KY
QEFiI7wLFtbicTtXz9HRWZ9gWQibNOS1q0BwobKPi9iXlJiyXdFSstkb4Aoz2yBV
bYkxafYil5yX+PaC4YboUmioruonVGe1pkcCUyXRCs+vC50JMqINWmgXxt9JojtT
pQkRoxwAZniep8AZCrGbCg==
`protect END_PROTECTED
