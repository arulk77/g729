`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD1Ssa0no1A+DVGtPXtKpcHSy2AoAqHHiMRUnDjb/NXC
abFLuHyVazhAracd9COdoZHacuA5AwCN1RxVIuLFW9VEl9/l/aAotLU/GxZVGF6M
hw5DsPZcqmgVVWSQGdYc0PDf+vXi9qZ/qg1fDp2Gs4tSIZlSUf0UpSeZNoe/zb1h
piSajtioALIFVhT3gOfQP0nfz3KViBb+n8akxV3+YxK3qkdje0frFX8utYCoclBU
`protect END_PROTECTED
