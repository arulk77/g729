`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCPmw44Ct5+iQQrVSgQKhZ46Gi57PdBBN0Kw9N4tZAPj
lD4KYN2LKobMcmo6Dd+eigYHKz8BoVChIXMANdT56hidozWRNcNMWZzinFk/oJ2B
juVyXuB3GzruJp5VWO6VkWNYGB5W4HuxIWSx8XEnmEmk/CIrRzK+Fl/cTQRTi9cR
lmiBGL82UwDa/+lmgFRgbH7w7pLiJcUoUQFA8/XPd2C4vdzq7x3iSB8xlJueCF4O
1876JQmEgmvbLT/rpBdoWtYMhzISL62NVmiEz5PSf5cM9kpM0gY10ake1thd+Cuq
tH5/d3B7MXxckRU1RbvKBw2gDcWYgpgCA7ItL3v81jf3DOkp0waDuh2Cyy3GBi4r
RV5v/kqSW0qCU7ckWIFc1nsQukIXebSmLCNN+1rGMAtWYMgyzHaFbxdUkXRCBb6r
OwJC4iQMSyoWz3e5wf0TrGgtg5vN7kc1Po4Qys2jc7JNva8wuUlUfR4hGNkoJ99S
uRD4JnGajYULeJOVbu8y2ebXmYrx13g20WZlOPXw5bJqNwd+7oreBviDcNFYeC/V
qr/uMfAQDzNfUqMkUUcf1q968sME2Faq4soPFXkSIPbkCclgYP6hqYQpCMSTrXLr
UNQ7ui2JIIa+3yv2rDuuFL/JUnz53WoNWAGAJxH27qHE5JfPnlEwF1Jf8EDZND7M
/m0al4t45AH+qBe/2NO7kSDx++Pb5j1qs4b+oAb7hAysTL4Vejcj+P/4N/V2shub
OPrJsKVl6eyy/XP+SUWkeBuPfOjcQG/yLCEElnZnjwmdT4zcQagD5qIRUgbsoXi9
Mz/sAWYz4cP3SkirHUgLRq0q4x1WUXEapD1Wdsa0jQI=
`protect END_PROTECTED
