`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMUSHNuYyiJAUMD6O2be11nARpClRWJN1S+ox9+aEgMA
thsbrDxrWZt2s8Ci0RUTLfRq6+Y5qRtIIwWX6micCiZ5Onm1PmJ0SJJJ4J11PdO4
v4+qkB9L+y3xyLiRoTs2O18Jii/BXOsMoVMUXKaRhelcFLBMLNvf7+BJgI0VP5Dx
j6PWiiGa/mXYekBY79+P5kn4QC3QRWK23Vjfyjx8fRXo4oOaHY8l/X+aBP/X4O/B
CZmQnykQib2hZBySYeq9Jr4ECWSmX3hfeHSB7s8ECQ3LcCShtB8RR9pLUix8pvi6
Mol6vABjIs2pjgfW6yfG4VsETaFvWtrUXeyaJaw74dFwfb3JW65Sp+TGaDlw9f/5
LPGvkS1A93Rdl536A95XnF0ggKKA9HZaNdBM0uLadOi143535RFARADCw+cNbs/b
VOw7Ri9JYXIGdjWYcBAq8GTigoVB+rh94ove8rrzvsnOFPDeFi7k9VmTM5t/IpuK
cDKcYHBxHwyFg/BPPbjWrC+10QljWjAuWQhiV/kaOssgHqqd1c3BEigzNpymUqIV
KUH9GcDokwt7bHWkaL2C29rl9hFLVdw7LsjBM7Ra6hVfee0Qy46AYPeUpFfIsq64
pAnHRzxD4yE0jIIDFS2Y7nNP98e04PuBQfZvoYa3GdxvcreuY9aiAecnC3xs4qNM
Nl92iXGwkJ38lB4gVagTKO9qusb9uSaee3vi5BXCj7QeSHNPd7W+am/JAaBoc9sG
uR+gpQUYt3t7O5F92/gXYJmFRFBzcG7TCWDr4dDgJMaT1MwX7QsHN0IxWAhCBhQz
sMh/9kbmu0ieWFxem0iMqUK6jK/s0W910C8WilFqgLM=
`protect END_PROTECTED
