`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB+Hl10heg5hAB35WGdW58s+UoA6r0MIlkeQzjJub86l
4kkz+OxrDThvmqnaEgrlirQzx2WCiFQzEMt+yITRNlh0iZ2EiTDT3lsl3YSX7pIz
chMI05L+sx1qwrjK4eoBOBBiCIB3GdUaj4gyYGWpK7NRZiwWlTASx8I0tITjU+fX
NJmapxFjI0wfP2+XSH4+jrBhZS8EZuys0g+g0YVNd8NYbhvWinh7buQcaVd2BN4F
TjkfIa4ibs5eXiB21OtZk38KfFTkbbTvkJvVYJwsixfRYAkPGR54S4JkOd3TeNUZ
M6/znydwEW7J9KYaJGrMLg==
`protect END_PROTECTED
