`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMm3CJzdyajfmxEqkMdZD7KHLPL3FdUgSnSBmxzijZCL
ADO/7f+LUSfjza/pH2JfKAwZvr463GRirBhfaGbB29Aj251QnIixhBkgi5nj2NVV
NyCw85ikdAXKTyreRWilv3V7dIliU6HTFbAU/jgybsQRPmQCRbyMkGhV/cOuNh3+
uDCFm54VcDxxk4vkJWqDvA==
`protect END_PROTECTED
