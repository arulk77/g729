`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zkK7/vEeIFsekLoSDYfZ3fZSw8hsOzuLR8odzsc8l15
FJwbY+0R53rTHCbE0PUiTtRP4/aUlm2PH6uE4SRwGfog3B/w66zqEPHHf/4/sDqZ
oc190u7eEDj7HxTJi3pnCEhECpXTqy8ZPwJ2vmmrH0LaUiiqF9P8TT4ZuMvChtXT
VmLNHzuKZqtb+a+qMKFSSS+oDFmZSRQdyIT3767r9cKTgbAq0BMBiREvyFnUdu0Y
xAeOMk1ej3XKwyyanRY18KLdbv94wxi+eG5lDzIzoaI=
`protect END_PROTECTED
