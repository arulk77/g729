`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveO+tIeAhxyVy2EyE+yVioN0aGf5AUOdGMiHzOL9iG9NT
z/lsds0jlVo87kJVK8s5whvRXf5nntkkqpt+0IwjnrkCpAyUGu9WvuZcJYLEuJJ4
c0wOfmu4osNDVE2Ub4jKfPVKhYmcy6ATD7u83uwNqUCfYNWUs3Vq+SpMvF2+NuMp
vHxt0ta1rkwfHXO+6zTaBAjkA2+98ESaY84WttOQ3znLdQ+i4fDnVh79qesL6VSi
F5m/Vy4QyBgd5h072I37r0mXAcFsNu53Z7VyDBjR0AbhFSrHnZ4AtbL+Rf69Nws5
tijJXmOGFa8f+I4NN1h7u8Bhk3X/mmAlTgBJN8nf3pKhoU5A7cnqMNo3le6D32OI
g4WSbHePvxo9Oxe8J/vB9VfZ+dZjUNNlVlesMqOsdRvFNALVInZ6qBJCk8V3YU3L
3eeULaKx41DtrEBUMNdqSS6IYotv1ZguLthFDF7Z00wWpSis6vgvy7/+11CA/DgV
zclmwUke6ZXTneMIxeKSXvGnLVQE1X7VT436g4yEUBHLgisOKELJPkft6LXpi6Cq
s+UVXtteqcT9XbBkFYyc0IaS38OaPU/aw24s6iunz66qQVQQm7Bu33O5drAb2cD4
3O7ydhKJi+HctwPh88doAv9LWEPBAcdo0x6p1RSf2lAEY5tqtO+ulRQsDlGAh+8M
NlHTsm2k8+H5Qc5g0p871eSonVA+EAgBryJW5mATyAZhf4VGlPCbUjP8or1JXWHd
iJ+fB0fH0iCeKaCJszDtGf8znu77aFu2T/23lvZQRTE=
`protect END_PROTECTED
