`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4z7tKyeVYYu/WtuqJz7spgRT9ZgjJKDS+dpo1+G49Wky
LL4puzMYA8UTzFFD1OVQZPoiYuPliZr1IdKtYKMjSu/mAHddAg8X/4M0tnd4cMHc
r5LV2umQKL7GLnMY/2gIu+kbVYJcQilc/oZlTR78qFHg+B2wUt7Z2csO/BDLh1IE
moY0bRxCJwkcUEUFafLhCGKNpKzwz+O13DCXE2ih1hgYnP/Y8Pd/uRfuWD98N0l5
MSuw/fMYpnCDPO7Qar/ilLdbcssKY0G4wF0PAWSVMfHyVNPoQhiRPSt0MQQUlhdw
IisA6ng1y3YAXHKXxvWUykPRPeAnOXrZNTLrXcC348wpeqqZd0OuUVjYsq8cSuU6
rHQKhDTGmMJLAGum2MK0YQ==
`protect END_PROTECTED
