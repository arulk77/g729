`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOTxoaEP+/C+f8vklr2tIDLc0atvvBDX2RugKXYIrK0Z
OvV0dKIxCYfmOJWyBg5ZSRBK9NwfSsuufpr0kRmF46J0FjZZvnZArM7ulymbHwaO
gm2CarNpcYPPLyu6oGM2fKOd5wnMDVcyemdr5JXwN6gfI3Z7OUy1ppZurPJH+vtG
Pm+3qP6kgia/7OVarv21QwWxsRtz4KkQO7Alk/yRBUa3zKInCC22bd9JHxDIhOEw
`protect END_PROTECTED
