`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMxWfp/cSJguywilA/HQNldf38EfONfeRM2ZstcYcwuK
YHNMB8BSOjXwO+zwvOxMPjdLpd2cwSN+vDEAomKsDtkXyAIZdmLzAZH9P6aCEsB4
5eF7qxeg/5B3lfYZMpbD6jAl83n8wwQwCtXXvuf8N1IDxHSp6l7cpjTBMH/IQ4WM
5MOBMoTor042JmJXcdhEKJH4r/1O/yhw9J2O2+t+Cs+T0FU3GKuklIeNAsWRcvgb
+SCVxyiSfDuokBWJn2rY6XRmoL6X/qVWql99rn03MxpnXFwId05i9bQpONaOPIRl
3X7a8Z37ZKYhV16Br6EtGFT2nxAVYMCT5CiaKoj6EOwkYKzdDg3Redh6LhkgabMr
nUSKbIBPVvEruNlpX9OI9A==
`protect END_PROTECTED
