`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK57ehCYzCwPW7BT6KGR6d0E9qIFQQGzlITiNZeK1ct1
LfRsWCaR1Kg8wRucB0OoimLC2xOENxM8tUT1WUteCCKNjwvt1yqvvjuh+zRGs0ux
I+SBT0wBGOXaKlQxXnaD9Rrx/98OMITTvKmW4iDqal27Ecc73W7La1Q+D+cEYqOU
ytw3n97K6uff/hLSU4Bzt6e38RpN40XKaLruRxDlTTUcIeYvF6sW5oV+piAMdei2
22CEpuRJUoJ3KRt0aNoy1QZNOHTTNpiC8KvuF5dI/Xxf0DyWTJKrEmXGXSNnIq+L
gRnLiZ8oM9xd37zFHhtWGcZ5hejlOt5dKIT4HvQMiKdESjZjlge+ah9FYawG52Vh
H7dNGc1dawdeDZJuyQ8uEPtsMxxIoVrKYMQY/ff9qMNgsEpkgKiHeEEmAJBPuKSY
ujmBKem0K4kjBhiyUYrTXZkmBsuaMBS5eSTNxL7jrUFEQKomZb59kBEYCWRbEwzw
`protect END_PROTECTED
