`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43N+bCXKWQButyrGdL42li0z2rWCBbG06foIsw4jwuhB
p5FUTPzeAsqGKIUbJi5peuUGJog0E+Tio1CKDTLcEhi8bSqH5GcgzUzFlLeyqy+g
Cfcc/3qW58pIH5N0BBhUPJg1RrCLLLE+pPrWy+EjwryTE/GWrIl2hTH7v/0Z7mmh
yuIBXmM1O+pYyN4ZpHfsgodyc1plhdmloPNSsG1etGxM5SR1mAShTJB5bMzgcHqy
ox6MHgeKZ9XahUhzy++6tL4RIdAZOsNeG/0AwG3wDXo=
`protect END_PROTECTED
