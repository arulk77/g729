`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xGagIvjabk8z39JGUbmlO9/wj4UfIoLo/YXw3a31N7U
LQZK83hZz3HKDjQwPz2R8FTZ80P40TmjREWh3pxA8RyMdxWQqbeRRg7aCUNpWzyY
Voh6fH/hDN1rvYuE5871rGlJoywvL7ENtd7bnJ4Jvt0STprGi9W+p50QyWUD+OoJ
QH1XCE2zMdrSgBl0220jaex2JH9pFW4PVs3o3/er11LXWHsPMAG8kQsuSrukMrR5
aBWbcxABhs/kFa5zzvuDpNsHMlrDcnHAo5euW8uEP5rRPXyP+y3NGAoKgl4V6zb4
nmk7mOQZ1Bro2HER9jGCkw==
`protect END_PROTECTED
