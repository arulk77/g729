`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
K9dt447uqsIDu0rwzISswHyMCo0jIu7wKnb2AZeziA8CLbSK0MMzW2M9MTP9qdza
HyVqncEZcTl2UJdptWX5PNh07caaKuDa8/tn+egakMMzU+5H53+/EQCVYtkKocM8
X01WrtVOxRBEvDNKFDhwQA/GI+DYT9aoF9Jtfn+DCtkygpJ82oikCZexbG8u1z3J
`protect END_PROTECTED
