`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMXgDWI1yYbuIpEm2VInSNKFyJs2f3SntgRNIMb3ukbu
MrPi6qjWC+rvVN0XUTxCs77a+xMhfilgu00M3JagS4k1P7j4/SILqHnvAEjyu4Um
2aDvT9Q2gE9qEpJaeXfvwkZHUZhdMjkyunnqXmW3GODG0w3xx1XfkiQlla3xE6+D
HDdfNnb6bz7/YG3cxq7udDmrrGYuF0zoPWJL9zTNtakD88LzMRveu4c6peH7cZwp
+1XDhf8N/FR+dkNi1wlBo/REIhfbYH5xhTF+IopP3hIhQWTGClM1+QrTbKsxEskH
nnZXbA72D4VVmTpee1V6ng==
`protect END_PROTECTED
