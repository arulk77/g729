`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG8uvhytn3tOHnwJnixz4hvsOflI1nmIluFzerRfpy/F
zcFCFo8WULzthiyF2r1ZT77H8EgUsgyFKJkTsbeQdaoJ7A/lROM/F461QxXAYyvX
jopvJQI9iKp60UjALrJzad5Qb3cKI7ywOjjAMFchLn7B3SJ5+L1Jx6A8sZoNsnJ3
vl1ext8dDhQDtWf+aIk3L1ySHLf1ZTu179JqU3x0qTBdPNx0n4h39D3434/FZ6cM
g9zr+UBvDKiYmZzAuhbL7OLr0Y3LaOj5DWp0MNaVn95jw2NaV5HWlUfaVWqx3ixH
e2wG5oMzIZBUV1o3rnD5EqrZDUDvs7dzYCUz6DgViFho846T+6xnftHUXzHO2X4q
yw6J0SS69TkhBxkakSu+AZYSU4k5oeQAqvyYjSL6Glj0lyzBD0kzHCAes1YLfBxn
8lvjVMg2v7HjDy0CKcxVOxVSnRCj8a5Y4k73ou5H1xnPQ+qqEWuULEPwymDH4FAR
cRThw4J1TqlebDN/CoAEFa+3jgwMe4Y7rqOyGFPE3Dl2IFYJx+tPFt8B/TnTtFCb
+JiF+HgrQguqjRR5bDoybo9+TMtJgjoxVyqo3PMDYl5qFtE8dUqE1wXpIfVezar7
sJY57Tp/VNkQYo5Z/94m4zlJuLu3dj7O3xFrMaoPZT740HiRqlbUEXuihahbWEyy
`protect END_PROTECTED
