`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1ab91WZOK6GBEzmZgt1rHXSiWK/vkdf0JBpTAKayg0eg8
LcxL697N1SE8r5aGP1gTLV23+uO6ChTKvMI1hGRImX80C6pQi9Kd8SWgSL/tvnBM
T4TMeXSqBhSMaz5FkbVV7INjqHdzwy4mW9DoLKH+iVg2c7Q6z2nb4mVM1ej8QW08
0JBMKs+soUFj34isS9X7jztvGtoPRIFtniBuJQNJhsN9fF7QnPV6yRlH2WZKc7ek
RDitLbRE6SYwX+oCk/KkPIMGmjOrJMpR9mofxhndx1A8n5pDlxBf97kjfY+CbaHa
vQD9G3PYSkyaHChJa5ffWe5ovsXXbj6GRU9v3MJpZmnN/41KL36UQpzcKDcR3pNX
sXw54v9gDb04YuEKqcs+JQMzdwgAT00/77WFADJIFeQUEDqZpFFiIw1eDlyRvMhr
HMIb9pHzUdsmjrYTg+gpqoNhepmG2LWPRAiutSjqdu4=
`protect END_PROTECTED
