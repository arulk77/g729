`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
SOghyPlkbcsGMkiPIgwlJSuLkymkI2xwsTcu0y1DTG6zLQhlqiRB8lDSYDFbBN/0
W3MIwt+2sNyhj8ImX0rWcwvJ5vfTC35Qn9omZ1bBJlb4+Ski2yPtX+uhFJpW2pwO
kvrH1oLOu9y/1e5/B4p6ikVhFh7IG5PMb+kU4h2YYFqSpj+FhEBMOppmRP6zOWPt
AWT6XzXwgZla6ZXF4RS6qRkQSbuyg6PJF6vicgm8rnzxGYY9T812k/+j9RvGOTYX
urpM0kkGskmAonLyUplhQLZdTxlOyPGupb3guTPgwYftI6JpG1H+uaKaMFj5A/5d
`protect END_PROTECTED
