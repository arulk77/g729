`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
VaOyk62LqGf2zAUQqX+P2mImgm3h5otsBkvG68ySHukm0wQBZ9dwHBdL5HjkQl0f
+aI7K5aPowdGBvp8gn73LEpNNoeQFpKMVpquSGSvtwzw2rDrD+iHmPFAqi80yvnl
h2/QyzeU/uYBBxQCJ1ICG4+hGXdbeXRUZ/QPZAXFROW5zPuHIgH8Nq1gKUoYABmn
`protect END_PROTECTED
