`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveE4+wQL3NDCfbDwv96zhGjCg9mi2KV7ejQXK08rfAChE
nQS9PUQNnqBX+qgqIFbNfduw+8mWiGbtteeA5W7wnMyUiS+SZ35jPgz/xD1BheMs
OmrEjNm7eIapVd6O34IT02xDISOHm+DzVXO9XxLMmb4U02FD2IdSduJ+6QcdkIsM
kh60iT5So0EObIrsFOO6BzKQSEi9pP82Vne9fKl6ispoFxdUO3tdEx3xpD7bzCTa
BfqkoHeRgirs+7AOy7s6n6pMp0FYQKNe+GbkofmoGE7MBoI/k4KwPJoUCVA/HDh8
I+zVkrDYKTuum5Z4xw2uJmyYRZ7mieKKs3L9p9ocVsfvX0MJz1QH0BtJ2rbUEl/7
d93hR+K/KuoBv2NhSctMRvmIsg3Ceq6rVzfDpXPtpKYwvKW9rcEPT9q2lYyPATDK
zC/5M/lbZu1Qs1+ukCEj6Hg5/bEYT4zsrceqtKlsyHA=
`protect END_PROTECTED
