`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+PWJsb4fbJinHq2NRc/yR6DOAxMF5a37C6ZddPeAbQ8
hgsNT1xMrw6CtxbofNXfVPgruYsRlKyZbd6THYU52bwXRF/XIeYYK+yV3xWYWKRk
KsjcbUzuNrm+RzOQTqbppif7QyqMsmYa0DHnmZB733SQNsNUXDnWV782gkPnIlFl
f4t45TBWke1cEyU59DLfyaU6cTeB8/jJ7OU4MwJyr97a+tiv+vRIuDsrxjVA1O/b
HtmyUkDtRTuyMhGLuHRchRCbZwylCf8bla+4yBtG5hI=
`protect END_PROTECTED
