`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+I0xjoFMQoqo7U1btgQoKaJf6Y0laM3s3fn17ix74dbmh+uNjLJZVDd0My20Q2vc
baWg9aUsUS1HHx4bxWH6+saOcCZEQgdrftC+RZYKEQtGlpAj+2m2B+Zyx7plOtTN
BmqGiFuvCOHIY3qI8BNuTxCXXCm3OV0ib7sw19kDJP2quwSe3WSAlijIk7k5TwuF
V027R0AElbAJyoRV4bxFO3jvWl7pRfLiIq2uQ1qcj71Mj8CLiqyyWeqGTR5NkrPV
DJ5r7QhQK3QusnF26MHhYjFN/zPqlbtZENZBawiGvWI=
`protect END_PROTECTED
