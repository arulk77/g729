`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveH86m0dkMXBl3ks6oVZhzdvuGMefE0rNWREb8+ogH12x
G+6L5TmchdLyreYOtkA2ft0VAOkHJUqLql9CC+qPoPZEIiwxODm7p2hdP2YixnZZ
3D/YkvrLxIHEZoGqoz0WvWx3gTdii3oYMs1JZOPizZ30Y2SekCjXoY1fuzfr3too
vNJuFNeglK68LzZL4Q69mcytrnlc53LAZvhd2+ISEQLmDSdbH6uFx/V4AyuGn3J1
5DqwM8OTr2d6e+m4OCxMhmy0U/XRJ9gqKYKMszozdVCoa/8FY/SUSUKc/oEHpdf+
J/EF153lxrQc78aRZhjpmqZWJ5mMPYtCZUdKmWCcS+XuHch6BWzZmB10TovfhA/w
F0RGyB3mgaaGJ8BoXcCReueQSEyJGuouZObiZATePS7tZxenfEF3wPT9CGGt9XCH
mVWiJNfvKE98jA8S0AJUAkA3RXQ04IPplndx8e3tgbVLzkgsuA7hOVsL2RNggMLk
G/6UVWVMrlC5kWHcXgdpqaOeK15xe4zrU8UPrJoqKFbBfr7VCIccbFNEs13SzigX
l9BGA2qSiR2YQPoDfTibxA==
`protect END_PROTECTED
