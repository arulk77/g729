`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB15Xl6Jxl2I4yp+ws+3BGMQsNFDavM2dXSV7woXZWw+
2DZDK+RtHMpeNdUWGeeD/UphErRr/MJUQCd/mWevvKc6dPI36d8hlFOPcuUrAQab
xbTDib/L5XNP86LeeIWGH5xE+YLmPS3RD+QYM7AeGp38EwCz+em3RcbdzYgvTSy5
vGgZGvN+bG8GXVs/+LNlBcP3VdNFrJsM1FLgZ0dp6p5u73OkEv3rVIJ2Qmfy+1el
thD/MQU+LYdKQVdLaKltfdHwYXqdDBN/KNpzIKkc4tYXitEMZW9uU1O9GVvlH7v9
Yta4hfxI3sMN+Gy/flMBObFNTVl4tRJS7U3a2zDf+ojUNjdVhcOGQ92I+s734Fl6
S3YHrpu2O9alWh8RNnkMPtyf3881WYHaznedlYc6t7q5w1HmLkORz8wigjtQe+UA
1Ryi4Ivj2n31B1jA/yzel5b5PQmrK2a3SKeXBquKqJKkTsWUK9NtFULCS4Zqp871
Kphd3znfOX6J8DG/AS9a8DDxqFmI+WvcJdgGPX9c0cP7RiafiYteYfT61sPxYWP5
w/D1KCp67yrO1DDaMmrgrNTrSgMTpWLVluznzeKD9yDOsDHeWDl+tMs2rxGr6Fyh
z83/Ns/6bvbUiJ4WhJ0Z5ijtoJoSOkbsuFDCRhIb1SmYTM2FXdaRtsfNWazV9btK
ENDEkDG72SBEWwSZAqyVReX7isXDOf4lKPX6c6HSGJ36OPYiGhP4hABdQvEnIfpE
QCruNeB3ffstu47PavCDyYyBUCpCicKsAYOpytDJZ7ouXbLMYfMZMCMyhh2X3Onu
`protect END_PROTECTED
