`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAUd2mH5ol71BkTrQao8i92bys70e4lN2iQd0/lADpjta
RW2ZmG/WyaSamBySjATF7lSmMFPHKLKe9QP1omQLIj4ZplSTGzZwGMz4S2ViNyNE
PhnECFNBJ/YtnpL1m4DaBy8CRYGj0ioVyw4O45kROtbpQG/pLHheim4iUXeMevHw
5RA6X7FZxX6xbVMcjnnOdQOCCEaGxEv0CdN66zMGU5Q6n1MkjUT5RXqAahmSdlkZ
4D/dR+d7b3wqBIDmnQDWJTeDG54nwpVloSRRcnT2nIeuVVM9P+RwgdsVxdrOdFOg
jM+IVRUG1wQvpn+pIDAau5a57a2RX+i5Hl38z3q3rpyKfFJOFnEekRmx1HaXjCs0
mtyc4r1goNmvjjryBaF9PCfHObXVW3jSL/YVDhnk6+9aNmw3fF36FBmPB/dt9Ccn
eYDrLbnXtomsqrH1/f65RddbeNXhU3veLFNOrouYpLIOMCSK9VLoLScIBtmuy49E
29w8j0LSO52WMoZ0BGWRYbm0wCidzcsEsht+lEFGgQjYnznvsvO1WAKdetp3Cgb+
5RznHbgjWfuiuc7/1kA5tuCYyYQb7KppClDydfkuWlQvLjtnnkuDsd9qk3GKuVYB
Tz0oN57CtRgneKSkOmBDhIi0i2EHwYzu2mZHxJiEJYWaCoX3YfnTfZJEkfs0iRdL
ziIfJzlPyLmzqbH9MwNy/Te0ms9hnu0c19IYWchpT47NZ2NMfaWmvPRa95VRaq/x
J06Fd4bzOu4ouhGrmWMnc/EuMWMplq30DXWwF/KJLvrOgGSAdeThCfJ2sBppFozr
9hfpFwrYwEufLEd6dNH9IlZLncCoeSFlv6APPuR/wGexYBrESGxfsLT4dTxs58H8
ZRV/de1tESKvYgsAW4ryPn/OBYgeaV8ijxwQCu/zk5u0yrzz9uJ2xHnC4FpA7dsw
6jvQwT2dC+LeYW4Wtbkif9v06omdpyB1w7zv4V9iG4ugmQDquOjwObmh5muDeevm
Jk7e+07h9dFZ77Rc1oM70JwKRp2YRFmbDHg1oRaqb7o3yzoW+shAycQyQuVxL90A
IlDoCz03rOZLftD1x1SbZrZU0ze40XzW7viXqjyW8PzviudjrSUGbWeHIUEnBLoC
7e1J4pYQimhGAN7lrzBIpgId628YHtuHmHSRqbtWoAqv78oUxckef7zdBoHOylm0
zqj+b117/1v6Xy53EHxMII1yaJ2CGzhb9/Wpbh64v3CduqNYc7eli8wBwMcfiA1r
PJBaaYZLLeOIJkFrggNJedxCT1nlkHt370derdoMcofy0OSyQy3O9lHWO95Eo+Pk
dJBTAp90w7doM/nMN/OE9xfU6TNxugA9BHXfWYkmD6ToPBOR9ZAEVHdP6cOJy+y4
l2/RjP9hEMvNT994OMM3IxjRqpg5a0OFjnSKy8wvXUhGvICqo7xA4ODU/JDN5+jx
xIORmoP9fcooMAVn5Cl/iZ5TtiNNK/R5SRDr7kRAwdMaY8yrPHzpPtczHhxNOl2/
ay+XZiRMXDNgoWvt0ugJSWf2SHvnB6PaPE7tLHG1fYRW9TBS7eGLjKDeg9dnPMzG
AASwPDL82Q+IGc8KPU6Af5lCx1pSjDrci+VTooG/r8OZXfW7uZOZzVqVCokBECZ4
f2Oa302ERSAvdWg5nTKHlsf1WFawlJ6lWpINfFuh38u65IqOaxkOp7qYBFg4Hc8t
GZyy4zdGNvkdxsB1sG4t0FrpA4LIFy0eUC85Jvjb4rAwmKH0q582fgZcFqZyJUCW
jBVIrDEFmSY0EC/65cF8LtZhZ1T2ZjcjqZNZ2bcxC7vOuCSpplwWYsQl8tg79Kic
XnhsKWXbm9+B9v/6PzXtbIsTnk7PeT/89rEIraunqVLFHaWmDAI3wEMVsc9R3MHI
FIkUt1ToOgRmLsU5+SrzzSyTNKUIBhzecb9QCAtogtZEpiuPIbgFMNMfgJx7sypu
V979K+m1QkMJAO0hgMa7NWT4P182Ezx0DJzqIq/3QQRazFeBqIkdnduGQ0j0T+8S
4ISxk/swcltMeIO382bgJCNMnefUzF9h5NK9yo7yQXlRrY6bLsLr3rdktH8WIYrX
nvRYgrH5hziakgbwPJa1pGdI0gJmZIRVnJN8Z3fU3f32lQLqGOmNqe45ErdOrI0n
LFvpbV60VEa42WZUNcxuyBOj92VNHo/rLDFZt41N6YxfV5cG/5wZA4qA9qIGgKTG
6GxU2KiugguM25kphS7nPoDrSePZobxvGv9zAt44EH1PouZqk0xgiQmXXhYb9SFq
iTYBftFhhGZwhsNHz1lRfoKRZaTpM4mocTM1i2VhRjafd0GL9YZWIATpetO48v+B
Fs3RTU6/WPEsAJ48Cu0EXfQiWdpJ77rpAT9p2YAUDE/6cPYJuz0KXJs4ucpjpJG3
estZruw6r5dzQP+jnkADGMNQfjZ0hgWRLmRFlJpKWbJ7zl/dvzdsfHbDpsnBC1Qz
qFHgjYdOJd5Pvfn/4GLc9uAyRixpFGPlprWnqLNSd2IpxvQMPM56xTHakBmfIkjI
7srLWCZ/PW7dYDnAyfuvn+kaObuF1cwe+DDRnobjUtxhMr90HwKDGeqtA9IXnOJr
NCK+9rgHuCph52jSbWKEFshDsJIl7RqNQO1RGno46xojTIuyVtuc61xzMA8TNclZ
T6gQt/s7hPgwztkiKXJb8JPoxbror3APGopTtuw+OSGrSDDFv8ouTORHCERGA5yx
YCn7O25PywB6UhIKmud4UHAFQP5Wnm0JTgH1UPxeSSxDHkeHzm/YEDyC+dL4JWWI
iod9hBm24jiqg52OtT4jxTXGAfvrb74O0Fq2DAjLLNDVThU6fUwd5B1CZMKUk7x+
nLK5+R/2RN745fOwpZnDd2uIb+9De2KxM60j8QKuhxBeVu4zGL9Y7hhaO8QqLMHY
`protect END_PROTECTED
