`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49QnAd9Gitz8qtu4Ns/tRadlqwT+b2UJ1m7BzwCsAqX/
zxx0TQcQ/brwa1CHAgteYLfY/SSvENvBB8iCHz6xtbB9xM2RmQyliMxWPLz7tgi1
ehw0funET5vm5pNK2BFw2FgO2ehgkyXUjSCuG/Vzah3GaO66MfssUGzj2O6u8yJX
g8HKUG+JQ8xkmEBMPTyvkCChduOX2I3P7dmqTAJBG4Vh9YTN6zLSrh97hrbEFWXb
eVN1tMmxttQtk7ZaC4493fh+/wlAemH8zKq+lTE1fYCRNiSH2Wa6t+RGomFRu8pC
VUDCn9TBYa2Kk/iD52yhBKP8yWYVmJXqhSTu51DWRuFDcQS+COBVXyks8Y6ehGFM
iNq+Pe4XxhiHczMgQGZ3Lg==
`protect END_PROTECTED
