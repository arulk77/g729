`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
FTtl/A7/jSjCriV2QVQR5uHJRzDrpAvkHzrKpR1arbK3wkeWEIz1hnJ3d/ooPE72
+DQNxPQrubsxmi6+0zcIan3+tM4IQWe1yYF0cwNGEEzmIMAzNkP0VYEMokGfmfa+
POTz3jcf5VIg3hJxqvwkeOyyBJx4lvSMLzjrvlmlO+0mq2WRJxMVWmpLs7nWIPXh
qHxzNbkZdwghRbzW7JH82ZpuyqbYHSODm9mAcdyRjnTWp19oZLuyF6DXdXvSgty6
nT+ZgqAVdi9n7Q0aDo9XWrrdFVZF4qx9ZrSNQSxIJAicd0dY9kGhI2rRpIXHzhz1
jUaYmYQgkjH+oHvvrDJYaSHI735W8MKZianktG06uGrskI6SJadeQt91xPVQGKM5
wYVx9wZEhBvaG23ZbXcNFJ/9ybp3dOI+TanvU/EAgCiiuS6VNDpniqLo0eIgu0Ir
nr9NEPbBMGGfp/r2eDKisG6YeRMqNjQbTTn2cXvvx090s9N8gbR/d8h+odJK/E6H
h9SMrQAwMdFuXX2jG5bv56NB6Gr0TB+AK2W/yzR+r/JxOmvIOn778bKGnmvb9Zvg
1RFoYfWT2Xd+h9spvHIX1RbMZHdvBORRXlThB+fToyzKpG/XOIcWptLp/3i2t8uN
lXnadqiqJVIMmb/JWbriMyeovIgUlk6vy9rA3mw1Xat8mrnfVboEkujj68fb9Ptc
ED5G28jO/0bluSmoF+7QrdezbmsBsfRIqdIRuLphgjHMfh1nPx21sJyOZTRa5bqh
R1hpc0vLMxgQyPdWbFfCHg==
`protect END_PROTECTED
