`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
dLnPMJHCTxqoSTbPpI1/1DdkXdJnoQEduAbawXCD9lutjTOmdbMUdXvadAz2HuR/
/rL8B8wHHRSpJ03sndqOGGjTImcY1igM7DhzYLgDPtHdkHujz357bM7eTjK9VNgd
Xf6jTndFxxs46qrz4GYNNOeJ0vXHubtfIl+xFnkKbiG2dT2kMkXOQTSN+evsQEo0
xkla/dgB+AH7jTCbQLv2/Qi5uHXTgV8IQO8VLyTzW89Z3jzks1MXou4K+3Kg5355
UVRrULcknzHWM9oOp+WBURc60mqzWDqr8SNNsZ5WhlcPGBkxpQQ8UI45bI7Ethz3
MkIv/2Ue6FaLsX6XdguDInkoilUaVpH8yy9ilQ2psIjH+MHNoCFQpvDUCHTAyKjb
2Fb4c2AWu6OlqBTddQFr/1gr3qUa6tDqbJDcDHoCxIJBqDZQXN7F/m/ir028Kh11
SF502KZ12HzDsUGVOXtnzg==
`protect END_PROTECTED
