`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDSo+2Yyhppqlpwd4fbPyiSrYOC5JBvWHDoSwgUHqU54
LtOs1k92RlJlcnvtA1lQe7SDRmxQWhIYI4MVzDRtjBP0HNzuPSirr3ywOEmcF2gE
UXfp7wsV0aZ4dTxvrEnockefjSfrYayz2zVx3G+AOzcQOL5yLlQiWcxt1B80s5d0
gVV0a7AV2wEVgjYqIUoF06LIGS1n6TyRD6UPnisWhgOEcvnbLDW6y0+W/mlj2aHQ
`protect END_PROTECTED
