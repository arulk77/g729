`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
OHsFqDPLhGtkHHMIDlXAwFfKalWI+g61HzEHAN7Et0IPofp1PQQnaePbS5ljtGb9
bbRqKloLdx/onbcyjEG0TVHr8vwVYdaz+8ZUKUTYVWKKACo+ERLaRcaBC/e1hM8v
Dok2M/g4FpEW/FBdQS8s56dQzaIBk3CmmurYootomiOi1WpVPRhQTuKJT+PwarjN
`protect END_PROTECTED
