`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
tLmzDNF6zJumdyd0+b9FjE4tEuJsb2IzYUlZlplIUNCPnB3UfVC6HvHLOIdDKEan
PP/xBcC4kSnMp3CPQPEWo/Wu5t1bgO03e5fG2HYOeuapIqYDVx2Q+1BvH8qVu+Tk
p6xCLiAntVGi4rdmsF90xMes2+IstqTIiMQZ7pKihhwzFiSzBDTIX4LnG3sXsBOW
Cb5/Lml9tKo8JkV+q2LwMVOZ6HQo9daNl032EbCmzw9lhOLN/P3l/bZfFYPMoVio
qduqX7vZTDk/8087k9RJ1K0p1NXZV2fuFFYQat8fa4AM0/dbueYJXPJB3hcsyPjU
whEzgHQ8XnJnnL5W/Smb9RI3hAg+K8+CJZdvo+RzpKv7DbkraPmzqAdBznqNvgsS
jqOdA47ow9eh/NUfpAOO0LViu3kuAAPqn+1RMmTBa1YTtk/kdD+AVbScBLQM/ByZ
o5eTTaqyHbps+k0dNvZ+mns8jfoEFV5dF5VAkkNU4BFHzJDnkPgpxEVq4aK4MMpI
VLApF2U4LPfnotgaaiWjDyM2M2TPgqKkLvA+CQcNokR92CUpHhsc1+IFCTbFKSec
T+7HznaTEA7GgBGzMmHyxcsO/MRxqFcEW6UlXHiVlLdN2xquHGOKCcsPpaDX66p3
6o0o1ekAI/BNVTUn85g0/tSAPFmsaX0CPs/JKviEnoMt06RSq6seuUAGFAzKgTY9
1Jvc5lOkbezNm8vMrZTM26BAQ9ikFx3/isjF7BrPd8v1iIblW9H/6wZfuhegwPnV
Q1HTYTknjoHjABPjYF2PSaIhDfODE9ztzWKmwkVdRPlxV6FJWyYSHHjD6OzKMFZR
IW+obVK+NhsKAffahX4CSRFXsMZX9o2t2aY2RntNmnnVy4qNBqizthBnJm736K3b
HWerE43Fh//En0vzykEu5J/wvo3NE/6ujRhdG0czew4cur4cGae1OHSxsGwKkspm
PbvGAG+S2LF8idiljMAhC6kDRbvmThDMDlNIi5nkqQBcm5EdHTg46ThFZ7azKsNI
NVZGE+7sM6vy593JLv8SC0mvHTfKvGYRizjLU/xrGcR5Tp5Y87lrRJgKzqP50i02
kO2fzqCsIYz2ZFWQZcqy4E/RiqLLfgjNcl5xc27ZlnfLnlUHm2rpXuDYKdozbr3A
CG1DBZY6CtZyV1zZdUa7pFeFskWzWsp9hZpBAeBvmkpXz2QngTRQ+Rcr3S1GNptF
QSUlBFptRxb5sXmVqvU4PtRldaNvSyr2DreD0PoO1u6VdOXpD1uZZl9jt6g+StwI
6+ioOmwJATwNDhFSl+0F1fUzk7kDEmZlYlj6JoMAhjSUSzA6fbDjAhal7cmRWmzJ
wdJnWFtRK9fEmY16LdOd8EIik5EzLSXv7rfzjkTO4POkC86ZtMimRxgSuJkiodNk
0KlqlgqmUISc+akYagT2kOO9YXFUzA2e9R8t9e56znUNE/Pa6OQeGXm9NWBFTeil
Yql3PQD5DVWfUzcsywk7sNeZZbqMhoRyHJodrOFs7e2zL9VvCF6pZOSYX5vjYOx3
5leQ/hnyBuO4g+mcGRwny+iWxSUjuBCz7040KTwUh994zbuikGQCOfqKMuj+3FeF
kyZoKdXd2TqRnmRmWiYbPKtRrXGEZSBu8ReUWeAz2roHQVYCmPnVc7cDLva/+3mR
1OKpiwp0k4c1CQaQGiqP3q31nTNM70EkHLP92h8S4mYI0+vyTF0lfiVvqe8Laoc4
PrEFU4uNcsuJIsXS4G7v9/jiJ+YCYHtGfz+USMiN46NHJiDdtqXpGyIPRpG00P2D
eMh/Upf69H/FP+QDU5O+xeodE4MCizkjAcND1ZioYbm7lAzH02rR4FAld7SiNkkB
pE7UYL5n7BXP0hLXaUHBcwYALExLmjn5BOHE6Z6122Rm0QDO2RU32rUkFtB4LCuz
PaXEpbW5Pzly1hDw+2FZvirL1UX1EbbItS2SgcJmmFNfKB3lTsJ2SEPl9xEIoVt7
vxcUEhWloXIjPYvrP31yiv5Rj84U/VH76N7guLVoIATzV4aP6dpNGlUPTzn6hO9G
K5LrPLcBozPF3+SUnw0bUJA4fyHpWq9fCFozZ7mA+Qf/Py4/7rfJ+bIKRReybmCB
TDLSHEdITX2/x7bRNYfZE0gzCGuKk0d+w7i8oPBHL61moRp43CquzgbDyGAF1hAg
2yfTsFSddrv0VKwMC2pHgMF1kYjzJ6CwymmBN65dDQ5T9RTwS3PuGVqI2X5Ad71v
n8I75pD7IZNYCm2cioEmJYLQG3Y4sZcPvDfsRr1swBfSm3Lmz7BRCtQ9chgFPf5V
oiHZqf1yT/FFu/RTeL55Dt8Ze0y2gMKVFIblDoDymBl5KYzOMWByakLtd7iO+Xl9
H+0SUL/BvReu1fBXNkX4VlDgGPd4pvSxQ8jp4rmGeIsr3O1YimWaYMqVFqEphhR6
Pl93cgPv2kHbIg4yGoZvGawc4kfqWp3sutSP+6tQWbeQyrL1MuGbIWa34OPzI0at
DoOXsXrMCG9sTjIna3O7nXn11fWgFvrYYbv75Zci1UWWfSht2j/9NX1vQh+VqTxe
T9uT3XyM6dKS887Z4O100CC2WyzTXjMkVTRZ7+rS91OXch+pzoTFyqyA+stnonmh
Bvb1MQsfqmrpoe17eAW72lQ8oJo+7ccAZYLlWj/8BeI29Hfpm5U1ppFFq4AJo8zR
BwC2U9NO1hcKyUcWwO5HMlOp6mVr5wGZCQP7mzDcga4ZX/Fu2C9f9ykGYF+/62lb
vaQmuT7ANZ4ZqN6jpdv+YSYU8+w3QbuVdKFJUSOKZeh6rxC4oSkG5HUcOsVbvrJN
Es/CG8OqfnWPRmBlg5ZNs18+beCsYSxVQ9gC1B8njjsVFtDQKDYIN9H5wCQtEupN
ljRn4sV1wnm1l4opEVnxn8/7nDVz9k0SpFuw9sfMg5FHCzHqj5WBZH7EyVRxmX/7
sQPfzKWgWZ6yvVqW84JqJ0jlSU4hGrVk9V7ASoMQMiN62ojUOw3niBA24J+6RcM3
KGapku6cg+iSW4BOf0X7qwXchx3Fwj9+MuKQENF9Rr/IrEt/EkpxP9GRL9S/5wh2
rR3yP3C9VbiOtpXg+RfcX0hDZ72QF7IqChcJnz3CfEBIVzrCNuVjv1hCI7tdWWlZ
99u1c1kd3VRUQMajEbS7w38IMLsYUNaBS6lHayofrLWkNCGGKmJL90VTJD78O3Qh
WkfXu+X69Z+zgZjOOcTaRL+0p3WvG1AVSYDw15potGdQCu4mK4m4l0uCU7LjIItC
ue8x5kUSVkhOfjgmNjQhSIeIgpbuqU6M3uHgiAl1K8TMd5YsRm9hBk9zfiKA8/EO
7c6OIwed/uHiKctfPLHpHwlGuUB/CWBgQ9ssfJWYZdw+W533Maa7IHhfFrvZa0MV
1uIwAd1Hcg3xskDFTCcalfXN/BCu+flQ4GTAyPdB8LNQEAxp40t8O9pFm72ehxwj
jsyXhk/pkCV4cpQDD0OjN0gf4kW/LWNlUfJvwerX6UPEM+xcpnoZoUr1Mxw9EJpx
urmDqcRaUIj2ARDjdguu/X8Lzp5mu9GFs/8lJGbmYdcnO3BDfdJJgokIoCNrT5f4
dy29SZ8CmpfaJrSL5to/+36xNK2MeLDTNfRq2PpwIDIl7RS9zU7F+EWR8ZKk7+n0
LfBqVCVjYeHlGfSgBT1OePQUPrOdI/iwwXMshY0+4aXZ8pKI1FummHYpzAVchMJ5
RBQ2TBD6SQr09AHUDEcRQDIdelkpSKX4M7lVcsdXFKfydh+DVEIPNCLxKeWK9Nws
d1rc9fmXsgBC95PiSwr10zrNhC7PpROJgmGzHrilQzJ0hgg9uqDeOykZWR7AiRT3
bTG5Ao7WPB71oJUqubnhAkQbCyaUmAoLWIixm18WYyhH7UeBi0VEbGKK7NA84Pek
WDwHFNNXWGuvqg3h/pbZbctiug6NzylviNnFohKHhof5X42A8u8HnbGB1piXKbya
izunoW0EkweWZA0IMnvcGJ7Wch5ejlv5c99r114jkIDuvYJV5PG48Bya7klvk/CQ
2123/BuLABq5fzOBLHSCt4ZqHs2QjiMuYmEt9TA0OQcyngdCabYMIWB4rIOJnmWf
PcilKIzOQ4fXGIxgK/aEUG8ntAKdnDIpY6TI/xbrh8nClld/sdCVTHaF5hQKYJgk
Kl9LhPgVi0YZrRRgX8sJEtOZrxq5ZCL98DOBubmM5Akmnp9YJX29VtnNCmvuiubS
YXh2sIcm0Pb29T+Fy+6pn1TAGOAYFUEDw5WnimIK9mwaaIn72QTXDiuXY05quO6x
YghIzkB6pYVDFVbKSN+DDvzHsiHAoeQI8zK7cYypbxubxCSFmepr8QPk9ZY0kq0O
zVEvLMLBvtF5azq0SIcnF/h4M0yxcvONmHXKm+tSN1Rkh77GOlQJr6DqaJXk0jOK
kvsfS6mN4TNmlaaTmBBglEazEuUH/27LrQRIqeqJZ3h2O58P/E25IsP0RdLBOBzV
87l4ZihRrAIdKR70DJT+BQmsPVGmjpdoYa2JTml4GYl46fZKt4S30l4IPsAhQMiD
mnzjqZ/SjQ7kAs9vau/nKgNUvBjGiwKnN9qYdxRNks9TEC2BvkAA37ON7LwT9Fko
M3XwVaKmEVCyI+FEgZDLHRfnzVAnkLZQJHVU5w09ewNMzka3ut7Q8vCWmD+O/zaf
pAKKcxpaIxQjb0nd0RjA3OLDBltCOQ+HbeASH2X7JgVajyM5ehWfgQapk7I3qp5D
r4b8tcLAFhRPJpTmHa/k19KB7d5yD8c5GEio9jul0JWrJIIsrtOnjcrL7eF8o4uD
TKQOy0mK9d+MK9NIfNfgr11+0RFPsdrhQyxr1O8bfvmUIQRWltKsFz99os6XQtrl
aeGxF1IqOLWnHn44ZTXLRBaUEOnpHiafCsT082SPz5RMjgTXJjhb4bdLX8povN1T
J8em870QzU9hoV5ED3bFY8an0sy2IuQHoXHJoEv/jIlFCF7ZRLn6/U8hyhwzv4TX
mrj6jOceShBOa6gQRsfa8wOqt8nG4s5QaZIpzPvGBqx+DBKUVt5RCMl1CNq4yHYu
kRRljmXaunQ7CHJp+AIwLDbGEtcIgsaK6fC8Iw/qxEplPfJg/VANgAxpCdG6/gVj
3Izg9M2zAhoO7gCXICi9XK3gTGXZEZoJ/vpNCEl8OBPbao5O4IDtS5n93zD1caA0
B5zreUBJPP4wYVYKQRBmK9XNbyieYytNt9airK8TjaeLzFMXWMaxqFQ1Ra5tovkX
ayoh5sr5+CHgz5kCf9tlXkwIKVf3D+1l/lGiTXBHTMBn4o12wU1+S2d++lQZ9ibc
iAdVOexdfhPWbNBq6NdQCDxpUSXTBhFG8g+2YW7EAjoaCikRhrqpX43r4ZxC7cSD
x4NS0a7x9fMsio++pt8NLCVn3c69XtrzQsi9Tfka9+pB8GudXdss+WwHvaIsRGNc
iFMKyXsdO4OPsPDUMhAPFODW3ZoKpTblhBIbcWYdkpVdhRRif4O8HRpTjhENkt+5
d6Pvn2WiKjFs9dE7VCNN47oZr6l8ivDkQ+QnjT5gXdXyCDIXFvotzX5hDJTsuR0S
JHr9wgO7XtcwwLRBZEdPvanV2sI3OSmLV2jRFmbBzg1OTqzU70gztpb5oLS8GV9m
H5/N8uiVJlTX8rby/H4fIDrv/0AY/ErLF3xIiXW8VyU39RwZtm7yb31wh+u/YBUL
xIivKRLyszjVZlTaUyycTB8ukFy481MC2qJDC9CzA/NLsnsXbfonCQ4K2PdilwWz
DlI6kWTq+6qe9I2qHDSKVM6qXE2yfBpCAqutORUZfh5CSB4HNf3L+qrpxysemh7Z
unAoggYu+xbAyd8/escxt3DK+oNRXe7yM45GLWeghIHjFAq+Wv6CEHZFJ6BPTpb7
EpudXozUfDUGj9Vkci17JYgkB72ml0RHP/634pP3GfJcCFEWfEmSexkn7rj473xH
xal28XE+9wd5yWQUwjVf8ToqvL6NNxu2Q0qH5ztmgM/xwc7nuaD2JYlLCfdStoMj
DrVMDG4ghOdLAXSHOiFofs4j50uZomebSQFYFmJEgJ1gp0yVMzeWML01uGQ3g+lF
4SZAZIBknS/HbJSbjPuejAKmIbxTlelNGEHFNaMykScQmNk9TA/HMDT/MvRzRJMv
GSRxNsK7RXp3SGIuLYIVL4/7JXhGOcHS8/w+q4LD/6CoIqMwm28Rimz+M5uzufch
o/uNt7nVckzk05QSXohNsg==
`protect END_PROTECTED
