`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wiXRV7vWFgyUPzpU+Ee/pbNU2rhkLinFK63j3NFxO7J
GFXDIlnF1yiHmh4d0QROIRM9emT0jHAZd1+O+btVCYRuHdssLcJ46YI0r5uxJE/w
yYvA42anVw2RAetLc+8pBLzqzvcaN19uPu7GJCgVIpsKbjJk9ieu36aF6/mFSsYu
YY10Su4afX+Zage1q7KeGbC3aCqN9IMwg+HErIqDzo4mRGclpcOemrrKI3QJ78Bf
/LxutKKYLmHVzPx2gSENsHzs1wkr7U2M7B0pwJOTXIFmIItSSq3MsPJbdJvDhjZm
2FIgC8q7O4rbkDRxHmFFgutVm0vK6ieCU5EoNHoS70RE+dJckccpScHKpZhhnoZu
IgcxlH80JQNnpZQDkEsjnmBSJ4aGnMQa50moDwgk5WEax80v42cTd2A5434mbbFG
OCz5FIMiDu23GZHGT9O4qFLwMjQ1RzMg9zeQYo+bXEIqEcRFEz7LR81krK//EEBP
UfskZEF5FG+6iZyG5IVTF1VZSgzlpNLJ622/yrYPJMd9kTz925B5HjjkEPeFyDXj
nYfPOmIRkivo0plV0+UyRERnP3h24QCmW53YyPTMq4nG8y7yJ8Gq1XI+ukVlcSLG
nhBDvd2gZymyrFpJ8wmaSw==
`protect END_PROTECTED
