`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG4rTPOnHdFSDII2+8eTTrYyzdkWzfQFpbN8R5RzgOuj
2FGgzu2qqqayHt/3q+Wpd8O6JJrfLk1nkLzEklCp/w9fPRPpPSIJlcvOtLsuobfq
IeO850PRzI1CV2fHLAccOc6lhbFnYkdT1g3Qp3tPRSRlkD2OkdnMrjd6SzRKxyeB
BEKMq16bUkYnUJifI4CncWzSdO3Qz2gSaqFa42l29Z2GWS9uV3tuEpUffWpQTh+s
3ZVQLHZc8CXW6IcIdmOZTysvXnyWxKO69eFCTzahNDMJ65YvFLQ8n8c9lbHQWa8Q
SGiYrAAhuIHYAZqufQa73h2x2VxgjbZ3a5VeoTCfepeS+j8uXujYxv0m6oa4W217
OvTn/fKscNYoSVQQv/Vk1BanN9WPDN9335GOXg1FjuE8yccu0YPP8KmCMWscI3Vy
oklFd8ZeUt3AjsKkcmNANQtV1zOo/jakl6g+cnNVYjgHdLkILnOWLeq1rgOMTEdu
EGD22/Y7atFq98nXOIJ7TIgw1VXe6B/Jg5PuFmmFEJtmngmEBfwehpog52CLtz/P
u0C2Pgf7Q5+kpP+Yn1IRSKspUq5IvIJeyRRQwYlOaMZsys3meCu1eHRVp13xI2FB
WQbfbc8Vp5XlsycNXGr9wY+0kOxZUgS/hf2tZWQRQso=
`protect END_PROTECTED
