`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFngQuYDAogzHUV/buWeLXPO5eYsP5XFXO0vlN3sxie3
2HcTXk0EpAwJ6rRkp48u4VlZD5u89HhdkvLIPq6fyOEnu6EkuHNBl2uB+oK50DnI
5K64xb9Fvn9UEBE3szn3j9Ggii1sOgO5ZBeg0F9uYAmvwK4pxx4tRAyipuWG9lEv
POk5wtMoC5VKBKzKALsXfVsD9w8Jexgh5I17IGeVW2IroFtkVzzu3JmsnnzFc+N7
xO1qHdl2JwVunz94kTVv62LlShoAWOqUh2ArAZrazvHy7J7vunp/Kcm1rLDbXQUL
3eA5h7iKsm+INkVFvtp7Q2OupNfoTQdRs7EEkXOAgnGwRDVHI1clk9jMfkCloWNj
CoT+5PPSr4sRy8V0edt0WIRiS3Beiu0Sbolw5dDS0fmtHtT4Z1tbybYkX7J15Fib
X7289IR0bdjjmZ07iNYplK1k3EcUMohCMHlY56m2t8ajcz0Z3dy8WBjEkQNj+KSe
N3W9yJA2J0InOFysQOlCUQ==
`protect END_PROTECTED
