`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJYAzivdVafqNdvatZKNt/oriSLSUQxTtKDt3eloEgr1
U/dZVmpp67SNxrDo8D73RNs1Rg4EHzS2+OIYy7p3Jj9Od1rYdJStmsNrHB43PT/m
uc+V1DExDa2JA4dYOT97ABPtjUNPQZsAbiqlKmsCaI+IqKUssTv2K2kfK92f3LMm
2KwaeG5W5DyYooy2dNdIshp0BO6jZdEeWmsAxGh3VKVYI8zC6TMIwP+dx8UFWLaw
IzmCCYXmMJPS/uFE0gwnrKUp9IerBgFG+qw2ohI8Ry1ImhXNwJLL+kApLFhasmdO
dXoLnriXSxNWgykNvuoSxBIinhm2axJ5KMNEMCnSqZUqB6xINe8WnW4leW2cKXBq
`protect END_PROTECTED
