`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1acgfq8IkPt8dvgOdaF5TzCEuDKeeyiDKzU2le3HfLsZQ
40wjdDiUQb+u+HDMLbloeEqPrHAXDS/P7ljWEZYeSCim/3HaNB+irAfz/41TNYD7
9LkRNYkAktAdaoPoVRpJ4F3DrvX/yc1Gw+suxJ6h2TPkijZ0lChpoBdc/o/0vzdx
9NQPjkyzy/azMapl+jj+YVBCAdzikvOu5lnPLU5MVxQJdu2VjffqJlxsQCjHRbJj
`protect END_PROTECTED
