`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEp98zZzGiyrkoZFB6OIp+naWTg5TbYyfiV/y+nVT08D
ltZ7mNnCX+W3MYY0gmgA0Na87lNgPTULnTNPI+0Twhp1x83W5F33Qz2EM7VpZQVQ
++PecJNFFSQn0YB/HlrXDWd2leEWD41JCSygPCVLiyMxn/JMfEHsCI0Fq6EMMH+P
SyvCeYfsmlxu9mjYWhfIFaSjkGCwc9m1SQVEQKzNm7eTi+DdCcLCXjQ+G6Sfw9tM
ttqLmtkk9M7CvHEcmtRI+5FTmgkBdCr1fu9VCMhkzmu8ccEet4QYs9LMpYL+KZWI
NFwFjMwzknJ2+p5AHsE6oQ9etmR6UijEuQ5RTO4FYTpJH55quC0+Smx/5zWwBV1M
ydwJkZH027V6Oo0y/r7NRgU61/p/OK5n6TOdxCuZrCf2v31oTs693G4QHQWUAUdN
pXjQI3TZJbT0E8KxD7NIaW2zCybKzMe2ONUfHpBcGYhINU6WFj7t4u9fd2lGD2m5
/jyHOQ2cVeu90S2/2kTyQ7OvxgyoeyXQSB9chjWg/jOiLNKbj53I2b8eSAG+hFun
Jf4LQlRWBk5SzJqq+slRSLdJXjopy67ToxcyVLY9JFU=
`protect END_PROTECTED
