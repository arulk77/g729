`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
zmGG0SL6BskVn9A9Qw7AwrwgeIEwLBKtv2kABrzrHC68FY59ExK21c6AK+DToCH7
RKQE8St3C14pUo+aYU8P4M19BFmH9TlzhSNcRDvCz4rr/CoVdOq3hlsM2K93RAyy
5L8GYcPIjKZb2+7aM44+/Ql4RxQ2fFABKY6D2NmQ6rjgcdHp3nD8/nv/YuC6ihXj
+wtDDbAGRbj40kpjHP3jfGra2u5m5EA/asSv7nv+SqZDDXLXQOspqIN9Kzty1to4
+J+xhTAtstNWw6j1OUG9AeyuH4DQaeX8/1B+0IUWBvkvwGy69rCG/7ZB5iCXy3UN
Z28i9tMkusYNwbpOtTK47sqcyvlDn8NWVBrGOCuvHAYbJ3/XMfOOGlxC4q2RJ9TC
EaiDlI/F7SWdNXbZTk01/VxGIERbPJVTPYapBQeH/dL51kSlwumKP3KbhRajs/Jv
zu4XDl4DymBC6lwidqJycYpKVe5p0ZuRAfM93dp7pWnGq7+pBgqhiBcnv0cLwGSz
BWj4pwY68OICmJiaJlKtesLt5d0rqFqFuw3Qbku1yvHerLSTrwPzsHeJrs0Mre7r
iVJTktS4rBS9MTLEjja7XY4mLebrjqLcfg2+GvPQs5+42XMa7AcWxiQLL0E9Eubt
aifHZnnbipCWT79zyf8WUJotvHQaddwvzpGvm2+kJlI/Ath9/hvA3TPnFCASdS6r
0R3eKdzLXrv/S82WPP2TRHID+VtpjATyZCn42HvcH1B1HuFzaKsYCsW9/Q6SQugA
WSmWc8l0yLY6a6FsinajYsHSrQC+8uwJmtDI5JcFvExrS9zAvP9YeylC16s7LtjA
qUYbJGCOISUQUifG/McHUPAWOJEOeNWCmAMtxhLonKCUvlu+KUVBkk49cNayGetc
IUMumochYlzyVGvwxQDU2Z4tMdMG+nTB14bbEIV78Sct0X2EsAW2s7gKcQdX6ioT
dLAIpFVxscdx+GF1FESmLko9Kijnt4pdjywG/svG6UQP1H4qXrkZApGa6lskRM42
YHb6iMhKvdODbDWdC9g1cFG7UkEt9UGvfjQDvrDonp2WHLEvM8koTCS86y5+yRWd
8UB5GxHqAYiR6jg/FkudpHZYoRNKhrxOQXYvrWKjFpLstwhn9Nh33T/ZZvsO2UyG
Mz04qPgJq/LPLeT7iId/QxHWym0KmZg7ww34Om+TYZreO/BJyH60LCKWJLPqPqdx
Ym4dSsmJUx01eZDk/Pbf6fIvoS7ki/7LKjAMuMjQ9QGL8MgkUsCLcJbPcl8PJPRW
b+3R7+KBaoqoQRH5+DHGL1Nfn2xP6AM9WvuYQi5ORNuAvAcM94LQLMydjj9eLTJg
89BFT9Ywi8DMK9JxYLxA69vjYVm0oPM/Clsk8B6L0kdNRyg6gRPbKfs0byQa6ZJK
FQlv7U74JyGigS5Gd8uLhdmRfURi5SCLPO3O3Mpzx/AsU9cvGFSZTCn/cLoFAKkC
HBENRrBHpjm0Vz3ClNFrT906vIVRtgiEk/ENM/OsxRlgGEhlK6pkPvJpYW7dA98C
sx4u4wHomEAV0clVw0GzpWSwimyTwF0SrNXCkBx0XxINa7rg7YShnGMJSOfaI6jT
1TQb+WITmRmf1KKsWz4BiozijnusD1JNzhlh16bYITau0ArZ9YkAVY1ROGwTG1Fx
NYr6dIioLERw+TwjpPXFOJJgh6eoYLqo8hxmD5RwIZ+REJJyybI+QVfI9ZCD55uY
GhuuF04hTKB4DM1KWimvsFaDQDRAJUYmskAhglyKKHrdVfKoHOmUF0xgRZcd95Bu
OovEAquxaau46pye8EiQ9vxbqy0F7lcH4naIP4vbsrOlmUiHPJp1lyF6ftiqqSjB
2gMWivzKrqsfykzAZbGGU3HXs/v5EVK3VYSxKle9siD7w9p4HABhNY04Ms8GuBy9
lzSjFMGY9qr18tOiAA++yZ2AJbwoNP8uCwkuCaWy9CCPKd9hHFsqw9GTxlwTjvWA
ab25lbAfS4VI+9BAihOrUEHRtD8h5vZ+u6/pXj28PzgtZh7iMXr7+cNYY2g9Egph
SNpYJ+W5YVYzdwGan1Gr/Q5PXVzZB8Qb6z1Tv/Br6y3EKTHLSwt5UkSn3VHDioSh
zmsJIi5J8XlR4/ZbG96vM7g9i9rObyFu71faMdJM7zqLKU8HU8cVxO4lz5VIK/o+
x54VWX1J8QfjcVUwD40I57HMd9yQwm0tC8+fJLvxicnws5MpelLpaauCBoGUtQnx
0jmqLdLHGLz5M3zOug/CEtp2hJJaNsXTqOAiukuEIWREmvGXVMKIHHI4aZ4GBzOn
l67EIP/qxwexFOd2JE0mlMSGhU10FQxgjqUlJTRqZMe5XVYh+O80hOtBgTZeQbCa
GAArZPudWT2v6RbbP9eoQvtKKd+6iGe7q65N7vS3DWeDVMLkEsLZISz5qR6SONEV
E1xIt3F0c/DBp1/SkY9g1OofONPOQAbkOoO536ce+tlLS8ybQ+FGTo1yEf/J+XL0
NSS8Nj67oV30dga1I0W/WT9OfWz7YEAhtHAdRfZiO4ahGr/gCqeaA0+9Jeg3fJzz
ZVK/Cb3+BAlVwDrR5xqDE2fpFDFPDdAkWq/CQ5R/Nqj9RTjwvF+n/fToiA00U5yL
6BDJKOx7GLMVhZjbAmE3qe7ivamJwIAj6eeG498PYIeU1ccbbf5gzibzdZdKPpVA
ajT7rqLnASltV/LBGcZ/d+yeG5nWdxgf2p4WnUtOoTiFjyu3RnabO/cHt/ZDamr+
haz/CusQr7DVPjY8WNe6zpDq4Pz0YA+L2nHjC6pB/avYEu9il8PARAhDhQet2RQ5
iTWhl9Xz90ScUzFfXP/G1PNpJX1CunzQi3BeFvtPrY/YA7gYGsoEWFXrPEUKYOrp
15iL8MR1jqy/tBa4VrsW1kQ0kArSkSbwqUf839br3QqUPqJODC6Sb1364acBtW8m
mxMaBOeKJKJE7eTiePplmYmf0M0fpo4qlWl+T0ecYTohi5To2VJFor2EUZ7r13Em
AZr3Nw1MJFbWR9REqYbUxq4fgDHkhMZYYw87VMfb9YLcu8PMTdUtRHqDWk8ssuFF
hPnUFijOnHNc0gciZnf3duqP4NPQGvsiIUc9jRUVRI/DDmNt4OdfTqw6QN+bMEdn
MHNJZf8iSI5Oqt2q+OfewKsn3UuxCMO5ZO29VjeOnzn8BZjR2SSsgFbcWQdGRhii
wMTnGgXXpveIRFMh73zC2FR8tFFd5cGIcj4Zz1/QiGuUFFoSp/JU1s30H9ZrIRfP
uaRf833mwoxnrmbHIS8vdd7hH0SNmhOAPTYEM9XUM9478n57fgfDpF3WGi+R/1tw
fp2zYPfK4ZQyS/6DM6fJwVj4sWD2E8fybTvZyVpd7DuORKo6jUfqp5RCoEg8Psn+
jeCiybJPkjmzLRk03ea8Bpz6JfyvPRgwtouiIbmdSRM6jhvyET3G0A41l6nYU4d0
Ax5IszfRie+1u5KjysEPpbv0+p4VCXknm5DQiXcWxzL6uq8RYcRaPY5iUH06oxTz
7Sy4B8pqxFvijC3XZNc3TLKkuutS8uOuoJSBO0vlCDkIKW+51ijH7ECbp3PqiH1V
49kpHgNNeO4ppsiTH68NAhlInP/tjgJMTNUDmfqAQ+ernKMygqreT6KgRYVKUfs9
RXqa2rWg9YRjmNDLbUjaUeRBoAZylGqsBEA3kb1N4N6sbZ0lwe3yaYhfbXi2kcGJ
J0P7IWiQ6A3lH1PJ6xEJ+ZML4EOldxPFmTQNWhGO1USVHmqjva1nGr8ySOAyUip3
JC2NPTmk/yIh/zaeHmaia/kZiNEQaAAeUOsaWKQLmxE2X9v2CjoS9U6WDU+ld4Ct
WZVYwO+MPJ4igmLIADz8DSpr/rJLEr/L46GhXc/4eWB3AP3+ZLaU1BYbRpYiyOqZ
kuND5sIW8WN3HB2TOeY/Dv1ahKkFy5FRSznqI/ZJcj2Vqiy6Ey5Ez12pfmaaqXHQ
ojFrGjWa4uU/zlqe7hpcpWoqDYvInzrbHCuUxpfgog0YupEfKOaxrCEQmRQieuMG
nhdGc/xKxgcf85FE84Aay3uxrVQ9xPOKLZiPY3cB6JEG4XBo7IJjDVeE6Hu9bF97
`protect END_PROTECTED
