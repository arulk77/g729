`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
SH6z4RN6pqLkMO+0eZaunXbqaiHJheW557haWK73WARtsVrBbrMIHUye36Waom95
IaCNRbx10BnEv7nnFzc2njEyt7x0iGHDdy9KY3yTFolkkJAIvxsDbfvX5avy4yNo
Oeq0DtxQWVXZNKKpoEgMBmXG8CmumgurytADAoIcXovGAIMpw9BOKouslKhSlkTM
2feP9FwhjaxnwlcG0BIZQclfSrVhG6zhw+5gRspTYmZdkj2YsnrrGHD+/l9EYzVN
7Ov23lEuBiKgMNYwmHI8ez1A2rbi4Eh6BwFRbbGe3PZcLVTAcI5i4X8QDifaM2Uy
Bj8Itz7f9b3RXRN/qZZn5xXObLP1fzV4U+rSt3QfBKUCAEHVltfB2IT8FbBjS43f
1ZoxeLJ47VoMMv91BgA6M9I24Kp87aeLjyS10nPojza9P9meECbQarJWMsKANIhy
L8EWrnkRSyMqTDhz7esJTOQLLsSwYY/rpU5qJnWr4m0XqSQ24SYXGIRbIzFSBS7i
2V8B+dVjO28Dtvp1cJgTkjU3OqMWhtJ1aqF5Oe+hMtwmh6//z908YUymXl/36/0j
1IXbUqet9Bp5T5Bb5bJqdwDf5tbmZffnqepzLI0t8GTMQ7NUUDpT4NUYo0QDflb5
FVg4xIGdt52m+5ptZeUm2m5O02RQg00PsjAdAGKnRC8G6F13kDOm7vQeM8lnZCu6
Ddlg3jT7z5I6TjIa1HhOX8Q5zxO4ZKYYJvafa0tKaFjsBSgFQCkpva2grGso+zhd
iAV+a8e/lrT0qQcV9+PVLD5SSRVAYnnKI+dH38A8f1gYlfWJzZskaJkWmlc/8XIo
3pW+RGRe8zAUzceX2ZdtVw145x12EgI6Pq11cgjpdglsKO86MH6rRGXQ0Bu7mQ1M
DrOh628oIy03hRA5fbNZE2TuwLiNf1UFj0ze63FXhEuvXlyN61RCSgJuYM+sVcfN
Ghv/I7w5f4VUGPF+O/3lpUyEuLZ4PyC3KmhW6a2G8b1sptDYTl8azLnThiQERPg3
z+yrkXRaTxnkmRmXShWjLVPbXivD97QZr1gXOsWdKb0k7q6/yi6b/mXJgn8eelg1
Ge5vH/+eyTk0jrPfPAH+OWI5I5xA6I3tcfartIRVm/ylRbbxX9iWzPzsptJLoRWa
whRWayKO+tBx6JznwcyIvAtydLzh7jY6W5r2AbtK72eEuJG3mR7d5hU9YG9M2Akn
pbShBnCMG4iUqzkSyYF39kyrd3ytmawaMv9Ezs5tO5L2enysYoaV4rKmGL6xDAwZ
i5glUGwcG5l5om8upBbtCzXHDr0OK2NLZp9SMWhn0s8LfTjv/72U/c3FMZMNlPVW
SlkFPOWMoi28/ips7iew6xD/C5LW4GkLlihCYJ6zBLU9RnK9218KwAeks9lf8w+c
6SSs1n/PWzgkfPYxu9kqmkQp5SywLgHpytZfxsJl7zU68W99Yj3KKy3is0RvBRSq
wTqSYMrhH1F6vtbQYSal1VaqD+aFOA5Sjov/hR+FmP1QRIOW0QT0mUlESVjGjnv+
fGOHzVuknFh+N1hAy5jzaaJpv+Xrc2FowNIdOsxUg99sgqZ1dIBzqEgRM9IwtJIe
emOzq7qFcIa7isRrGhfE6cEm4Gpi3Yy2n0s/LojJpMrWxP7IJ5gpt3G9Xb663Jmi
XcFCzr1YNnmbDt+yQX2HLwmQbON0pzMsnQjuB0qPauGfdEB7uSUEPrbrm2K2xCij
r8GaYDy+827OnPh0CQl3pA==
`protect END_PROTECTED
