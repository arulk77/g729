`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48+63tYJz+4hQjd+Icf+YETmLRg9jak/F9+6s29fDuFc
FKSasLJbeJWsmLteBbAtwRpCR5kM85LTDcxkVJvxbGmXo3eN3MDo9AgHHrPnJBIm
F5kWDO312nLJ/n4A2NLsPAfXbSFdr8xja6IG+Qbd2xCdDylUQsxu/DARE1iZC2pZ
BVly8fko/ib0ANA0lC3/1/GCrtcz28yXmKOZbkCFXl+EH6a8IU6kEbkvdr1QfyRr
+4lbO3sNgwrNT3Z88cSM7pZ5gQUBJN7zPj+IgC1eeFgLK0uPlEORMvPneouBftBY
pR7KecPbdcuVkFiO3NDLfQ==
`protect END_PROTECTED
