`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
eSW9UCz6UWHfjkdZqQwjQaKrtfjVX3wgieIMZb4/qubT5JluLTd1r3M7zvZ9JuEe
Geer9MENm17xJA80Cw8lASlCNBilSLLSy4tnV5Cuy81SjfkIrY/1HKmm3yqby7fv
FgnoHXqFyphOtcBACZ/cOvOMXvD2RoDBAgm+Wyly5p7+4qF0ATLuNP0EKtxAnMKj
+VNKBaj16mKroEEKmxgp/tE4xi5Vdr6dE4uKX9SGOTfLa762Lo9neyaptjYKt+7v
/+fB1WGJcrvLOKBJaqcs5g6z8lsRnbbGoJhju0G7R7HJKm9qyKBIM7/dYuFxqCP/
qmtiwuJQyWxELczIxIHQwHUDyQquM99Z7wRxCFhMOwg=
`protect END_PROTECTED
