`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAU0c2b+kuonQSYj0j8EiDLTQKDGkTzpPyJbsJZj7zZv
RUmH4CqsY6GEPQTegBgLCztCHA/EwgvRfdhgIh3au/bD6w+KcYeM/u4f/O5Yf2QU
9a7wp3q+npCe937pt4AK/aA/reSUTtlRhg8SCwRm6o04g1H6BHmvdljr3qXRD+6e
2fWBRGfWYdGF50JbTUxRPFheqmnk0TD8PnlOWRJI8qBp8XWF7GAN8VEVdFz0yo3P
6Y4FDe1TBE1ZBf70smGr3wa9g1wSpJNVlupIOmqxpTLUQRvrbAsEaDKPzgcjwN69
ekxujkWffrXAxctJe8DUkn1bEMCSYCsEe3ULqiUukNkDrXvjo+AZj4NsBPOzb9K5
Mraa2oJhyP0oRiuvS40HOMRWc+fI6GT89aMDNgv3X6FmJHNvcYDbctLgTqyhj+mx
ZtuChHOBj5LXSz+LK36vpghhJqhLAeDmM1vZm+XUsLoGWeUSH6Wqksq6GUSJF9Qu
IOvzpSo279nquYpGXwUewM/GuHQKXKfpfbjwKZSLRGjho+hmO+Yk8j2bA9SBCPUO
`protect END_PROTECTED
