`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
AXf8jFGAkzY5pwJv88Vkbsz6e4kKEWpuErkZakzK195+ppUtW+EfhKOomsYGPj7s
8u01bX97SMxv9SRU/lfgRz1OVuTEzmxGP0suoYY4NqnauZKr2xVHyhZzEBVeBLcY
R8A6hSKMo+T7t77rRZqu6u/NFRHuivPsrnfKE3CYAo/k9gZ4Sq4s9LaSmhWd7tsI
eJl+DMetcSEqmL+N5Zkb9C9hmsbawjRt3xB3T/PFepCPBywXIIPB/s7M0G3kVxv1
+KH7ocCV7PqsiVVgMMrQFoFcUwm0FOVOCK2PT6kX5gA=
`protect END_PROTECTED
