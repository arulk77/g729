`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40qiD0Iz4rvttWrzQflv+4MBCWWDvvQ+vbZW6xBL/WN2
38qRX2XIu3a8v0mtw6QyAKCF3S5hfugfmWQ2kF8MQCn/95E6Ru0MSjHjWecmgjlW
121xopp9MStAYIQt+GFRkGfftKODiVYbyv/ENv5FMpO//3lYfm6JV6ZqKrvEbL5E
hIAXx3qP5FUrfha4hQ/KQ8CrL2g5+qgeHQjf4OHbb9eVbzKq1hXSKCWTe1JMnrni
buAzzx6hIA9MuEi0tNhnk7CGnIzhZsml81zsYHWS97a5Hd/y/M7eoyJqyEkIVpod
FcoufTMH1cgFR9J2HotqqcQvp+BTROnfhIO336loTaS5O8PVi88+0DMKkYew6Vhs
4snjiNyu4P+P+NVSMKiz/jjMLkiljFXo9pctDhFUQO6X1++PTgc4xNMtNWNpML4n
qsTcYx7eWwFCjwpVt8Wvkp8hWa3VKMFeR7WXduY7li3+FjSCMOdvtra6edIUwwgB
spjlHlSpUiC5OXfUf2RrKAbwK+7zsxhad2+nl+x37zfq7bAV/rXbf9HPsaAESmtu
lm3QjB7pEW8nGoxlpL8jlJ5bWfRjWGcitIIqYSQrHaYcmHFaafLs8tCmFcbGxRFH
`protect END_PROTECTED
