`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44h97pWwZDPl5H3xC0vt3J3IhP7pUBhRNravDIE+3Kkn
etUcU6uMTMtLjQyfB8E3xTIwBndsLiACtklJLsDm6WIkz/g3xmf60nGy4vI34Zgp
mf+CSESnbLxBhkSubMvrp+1SPoSaPRtGXOxZd2CmsFeFXJ8DLlpfB6qkJitNBsNF
V+kfvZkDvzfksV9Mf6kxug==
`protect END_PROTECTED
