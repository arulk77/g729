`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBIG5IVqpWqllScnPKiEGZYP6V203b27nWDfIbXvR7gM
8IWg0VCHKMydQJjLqAhIIaHipLpxtqQKEaMHA7TLzBZ2Cvyq1NefT2+LFn1NW3V8
etUOl/WTzqasnFdlnYbQoLf32NP38cStPI/5lO0wxMrRkpV0HJpjQ0WH47V1tbEw
MYUn8qh5g7zaYGwckslIg8YtVbTYflmMCYbJIGo5ZqUeQVkK9pUexgr4pFc1U4Qj
0wwLloQcVrsYu1saeXnI5po839BLShWtFEYfRw7rQppL/drS9fq/RAOmlsCHQ7D0
8ieyPujRrci+tFaciaSj5Kf66R8tuJ6EZiqo7XgZwkomEjTP89HaP2YKCsTYou4z
fyJ7VzpdI4WaPcofVtioHg==
`protect END_PROTECTED
