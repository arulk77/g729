`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SbAIs47ECn7iHKuT4/trKoQ6Ch/x1EBBjWTSbYBUlH1a
ZaaYM0JqAXIaOW4TWKApVt32+s/pcaBzsu4iQ8izU/+KF9A7lSJxaPnIlwT2vDkt
A0JRbXSZ2qtOcNi1CXdJDucLIlm9LVqwkAKNgyddcaxkxgHU5+WTSnOZulgyj7Ni
KbJsWdnOgZMRt14kAO1YdKdkV9wL5nJcQJ68cn8A5yVtwaMzWsH7gLOdmd0PeBWP
Qf8pwSJrTm6Al0Z30RcXOZqvvvLd0pBckGussA3B6a4z+U660QjB28TsDQiKH7U4
W+fQ+hPga9PYUPQZonYc+iV15/ddbS7XptzkwYIvQDCkBTi/k68iz+U0NuD8EQwG
qWkOwMTKPMWh6kkL7W4tk0i85Eubi25goSeIUUiqYzb7qK7An+J5TRpk//cjzJkt
jioKjR7ipVtcI2hP+cNQ8HaL56j/UFY1aYRyE28A/Scwr3EiSui3Cn9IJivW3fJ1
oy7SsBmhXH6wfPkOK8Rn+aiumq2L6LeC3pnkfwXGgsJwIZsLr1anq/ndfhyOizJl
VxnrBum+jI9SeGPwzUDGLyDyhBpTUQso36crei9o3Mn122IkRfTCe9lQL45A4Ec+
q2UbCiffqQBNRLIWSt5Umj3a/TH6R94p5s4fmM2QZRULFPE+KVbieLwpo285XkOq
G2LdyqOI+5baXB01SUClee4XEd4VIdDrdk/YbHGGJ2TS65o2aPYKIO8XPUCPQdcy
MP0bgD/f16WCa1l3f1JUbUTkCPIB4KK4PAv6WgC80i1WRtFB9b+yWBla0bkYWGM+
KPEh2G2q+f0Ho9O9LUXrxfapLKNz/wr/ubFMuyzv/LUfIqoPekgBVCRjhtKYwKkv
OnD3gNS6alR1FSIGFhd1LQcChzb3/j2IC3EugmBGIs1EzpZENC4Aj0iprYJnzV7C
64mrkDSr07ssSCW7efge5GdOaSp+dHTAud08WU/+1FzLFV6SxS2GtEomK0JwTb5J
KVvFDc/7QnSr/a/j11BDyT+vOaMYJah2eAfkHPi8yJiVBwHnEgr//z6D93gDprxv
tB0zRY6W8xsnhQ2yteW5vZp0K/XcZcAaQ3vfywrDN7Toe3sJxTrDmQIH/7UJQvkx
q0vmmyyzyO6oWg59ua8PS0Eqj1Eb2XHOB9IWODT0iY1stQQfkuV3mf5cz0pdLAt9
1k9HqXT80oStvCnTuNXRm8B5k9twvklQ7yEB3gN3B+FLpzPAgOvRjXt4H4ClwLf7
T3SLcOguA9jniRumOr3yaJi7+u13cJ9Sa/wdj4RV/f45aIkG33c70mzgoWS/1p4l
NbZC/Aaaz7vjWr2RqE1wnFv/oTCzTI5AFjt82+xlb/kVt6xQ9I4N+BDpt3GKou2Z
/hQR2PWfcQxjBw9ioSMGyeSgG8S3z5URddSU95DwqgM2Xs4Rl5WRxtR9dp1KaYKd
yMnfEajIR7lkwjm/PbN7ytcpHNWAjeKQPQANCbj3CxEJmn3VhL5Gbum8je+n+o35
oFeE821hFd2H24Lw9C2tdIUOCRYm9oLYP1AKj/c7EAnXel6Xw+cuVqsUReJRUq6Y
kMDpgmFkPEssjnQWr3rMp20hOejrZ6Slrj2sA8hcs1fUzNRMnK940qTlmICa8Yvu
5LQg6UL/HFCh1fihsB1jo6EhyIej7qYbTqKxerRLd9c+stuv9+aY5YMIHwuM47zF
mcO5NpdFZTozQ23zlWE/hzbMTJz7v2e2LXix9ZG480Oc89O4pmAegV++ARL+Cy7N
EFypevsPFM7ksxIgy+5x3CIIqoFDnasXiXWeJHm9g4Z+Oz/cc47ZVTCpkpXXm1BH
KfvtQ+6UyUDxhU9h1t2giDZQJeXKT8aAhpmBWYl2sdhm/ICMZmc8JGZ8GuKeXFCX
r1xnEzpFRFwajB9eKhRt/MG1dQXJbRL+qFZKRywiZFHcrZLctLwanvdYNi3U9WvE
xyQCtAunilAWpHVWjTQzFuyFewhQKCwpEJCsJcgtCqkdKh4/GrR9UWdHm0/Jbfcg
gVJXtpgwgoGe8Wt1KGNr1JxvDO0EHEBt/1cUZEOVw2fHdoCUFypH2rsuv0W8UCK+
5GtS2fOfArMPK1EYTeUZuNZx6ay4YOoIZkrw/jeCRPb2Nt9C6Y8M4XrRjBcjYgpN
21CuEBZPzvbLGRRuB4EPNhaYSds9X2L3373Ycar8BoRKrOtOR/EsMfhhOWTsSHj+
1afLRZojtndTp/l4UOw81kmPTKXeTy94fGiC+XGr0HpqJV2CsRSXO9iY6+ffTueG
PD+ISNDysmX0TLTKkCsimkWcfTORA0vVfwNVYebRbF8etkGjKhN5WulRmMQkmae5
hU3q/U1WrNtCcsZppUnpH+fOfR3N3W6gEO7s3HTQW6w5KMimddZS+2Mw+QODD0jr
guTlwYNoP6sk7U9iBeMZnHjGPsbe+cI8LiOF+F2fFgBH9GV5CcUi3+WWYfxxMcLn
Pnd19qvZhug3u3FikCAbvJKCHW9ZyVmE8DDTFMjodARvEsN6JW/zPDfl/0D2N/Jz
TGl78oVfP0PpejQCkl5bS0AZnTd/lCzWKv0hK7ZO++m5x6D+tktMPUMXSzfRZLrL
ZPwnLgS5qV5UJnCK8Q4Bhxah5WupZIMGa5uKqlp9HvXNA9khpIkEZZBm8Msh5dM/
VtxeD4AIPzJdOwbmdDyubrh9m6PO/L7qWawn6nZltvOPBVhY/B3w9EKjlXLW7gp8
ZP8/KyWezg7igYCw6DGYbOMf4OxoSAhvPKyDbHESXFYkxHk6Zw/IpkCp5fv/PYuW
yqPAL9D3af6i/L8mIqiyTgCfMPZ5tE+MznBwkNeRPqwVmxE5bSzIlwbWuEE9sMWW
Cf2ERchrq+vMhTV99u3ZVq35tCjgw+q3hpzKvyXkbEXtv+/F9HSMoXmZAOJwAxXT
`protect END_PROTECTED
