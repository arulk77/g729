`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveORtkbGOyPSfa50Ru+LufH0637XcidhAcf4X88aoWyJv
PfrjlO+owjFHVt2HCp34hz2YCzK5mGXEHr+a7nF9B/v5Y7ym81u/mttbD/nrBk7m
G5hBSEh04OLB1ZijsAfDr4CE8pBhsh8wkHBp+RWnpNpsUfaBhlE1HhYqEjQyTxwx
gJJQsAkKPsYb1QAHqigNvLP+OulN83QRqtUrnp2wkMqJuaC76bJ7qnnnfS/6nF9I
io/NuGNS2JVgEDBj2Ut/YfnzAdRQtSRWpZETdAzQN1+00ht4/nJTvS4cFQDEprr1
irPqNbV6vNkRb78LhPpQoaqVZyUscN5qjXTMEF2JhIsQgwQO1D5neAm1EE8+rUDk
5ze7iJg56SGrl0JyCaUyWjj1KQzzMLbT36m+VB+GhthGBF0iLaBgYEw+d96R0QsB
fj9uRuqm8/pkiBfWHaJEplUxh3twm7CnjYEh1iLXkC6xOlVBITd9UWcNonWR3ZFW
CiZoXakJX3Z8pGxkVFe1HlS44rwx0HWWXrwLUxuuUMxoOdMiX4ayAqlBRDEErHgy
hryRFuw8mdjbZhEKkCxMbYbB6NckoKsaslHWuz3iOjD/2C97yE5YHDu8jedccdrc
`protect END_PROTECTED
