`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCdHwJVqI6izZAGZAZ9mPVJ9ZUsm0GPvnWbn3ib0A+2D
kY0kGG81UFBeTwscFgK+HUQC4UdK7nsvRpEmkzdH3FoBIfayitIOKoyF7jlO3CKq
fHrhFORDeJKkhrd7df22n3F7uMhDVSMhNanyo1NWk7PmmXeTPiEiZG1s1Ujed3YY
etQI4CnVuiSwvVLSRjLFR0KxbUhXREc8hkPULJbhn/kffXAAd/DsJ8vsMpp9Q3q3
LMNjK185Kv7evyS9ilOizw==
`protect END_PROTECTED
