`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDjJ1wmWpVdRAEITyurrQSQd9QXXnmPwDt4xkXImFabE
gAHe46CTEqhP9WbN1m2MsyoeSHNzaJvkbK9ywFYz0pqFHDLRFYu48fI7VLOGmbyU
a290zqIx76uG8Onb52s3nyief4wLzDQGiVK9QczHepUy3M7SNoNhwxZvpog3WFUl
osDedkXnp3SJcn9Ku++XkcX1hVu/SE3fLYRClNZc0VpobWBz1gwWOVV+yQRoqPuP
PU9+b+O2CCY+7xokiGksTL1c9If7gqO5enfTmk7fOegS3Ziaj8uIURkpd1AxHcHm
LZN8hOu6w7cVv5MytV7ZjOj5Pr/TvKUqTQWGl3XWJPnka/dlOithMDXIBIWCrnIi
pk/OYtNOM1ikutjer/ib7bD21sLxMb6tiXlO+eW2cYiptA/wcBPY2Rdf4cNST+Jl
BDssWFMyLSddwfz+5T0AW+PSOC9G6iLZj72cfn3luWNpxsaN2XnYLsYZGhk8wh+s
`protect END_PROTECTED
