`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pnyY3jxGyCgnwWklYcFi/U8jBw5uz5nXmHa3RXFz8rBaQ2veFKysULvpWHnaoiGe
b5qC556kjY4Nqok1sViLMFNOPQSrGOaruqnGYMquxqHhNU3A5WCrQC28JVpztM5T
gy1fjuI8xZQ0Bx3d3oef1FN2sp3OmcKO5f3/k2Yd838h6BAs0SIKI90ucoqGbN0i
RpKg21io7pI+k/apvdnqBhxim/iYju2rjhWAtXt6JXPEhlxdl38WHNjeJFlqcnr1
SMk65YXlBQBhfVxGXFIzzQPE0dq5I4xpaGk4M45RFYpZyZ6TzLwxrwEGmZeheSCc
hJ3esI/kJIO9TtFQ6Cz55PuagpH1oejr0ZTU2CHsdzYF3m0XIuGujN4TaicovlBa
aQjD/bFKYTgP93bll6Q7ORVngJ+r8cd9LgRf627iukbtyfn3AfTi2VIL0iVK6hNI
q21njjStYCGi/MfSSjG/cDPyyJ/fcW4tTR+4waqpC/M=
`protect END_PROTECTED
