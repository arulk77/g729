`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN3UgzCCrridg7vRorzqX22gh22r38LSJes6aVSTpCOwg
8xshWI2hxeYlhEkssR1DTFH5aEvkGeSpuqMZzcvjYJ514Wqf+s335AHwelD5eEtb
7MdStriWkp11He/pCGG4yDOERJZZRCY/sCCE7Dra7ytnsNxkt5bPCkBrdErrXe/q
9aaRFcR0PD4ac7wfKFDbUlLNxmz6eRD+BfYTGMpoB28TQ5V/PvGNztWKHJFBCIIz
IfMedWhsNqOd9J4AXyZZGarF3zRv1bkAvzJGckgeQwgQNuIlyv3c8VztuSMh/xVs
UfVmByrgZ5I+90NC0ar1yQWE+sLffQUOlDjlhvWCZPZGiaiDRZ/K47V2a5kXcHBe
DcmEKjfaeZAdMhgEXNAKjYkMyhBRAMM+m5J//W+qfUWa8jtodLHBbm6J4kiKNZiG
Bp7nY4xv2eSaG3Nlq/fDQsQuLGGJOUZEc5ge6DJNJrFrxwKxQjAuwX4N1rLzk4Lm
LTm4AcEzpk5nQT3N5QiiQ9wiF0ucE8Wd3x1t2VC2kWmvPEUs+bGAAfiynOqQP21c
Oy82xr1XmFtngidBt1XxG89LWBhnrCJdsnrIW/g3E/hhtxiUBjuLGccZD+R+LPLD
jyJUfajYj73KEBaIwwxMH9viVCaN9T8dX5Jzjgw/AvqmGGBwe5yGoZciefT34mmj
i9uq+Oh7jxRioOkW92pQ0Mpy6WOi7xNNc3EbyZ6QKSbkUtT+73zeFX0VKw76i9/c
Nde+pZTO0K2VFwROonRejXTNhEmt/xmBcf/WcEX3Uy5w+6Hqml82aPK1nDAPpLWc
gXVV9k3ItjIFPHifKGOuctiL9CMAABU1yRBivd9lKASeqr3PyInX0jp2lRsPxqg5
XkUGJtUsRJnje4H7EQhiAhm7oh2yLFfSm3Ko53coLI1ogzTbgJukFZ6d4EUR61u6
nTy4O2fkDHOf/+b8OtWanKjj/9DOaX7eJdXZU2tXg0eEWqVLw235S/5x4Hzhdt6c
6ZDbfRpAIobaj/2u0+nKGprqGFLbfM/H1aHF5A993d/VxmrUgSYpLl4fZutPDcDN
mqvJ+64yzTMDR/pQX0w+oD4Iv0/KKM4fYRhLfkBnDy6lZRBkW3vv/bzK3jqApA57
4zbLHEF/VFmkLPdU5Se617HH5kCwxYFgyPosR7J2pOkvqRvHAj/SsxUct+2Twkc5
KyrW+7nT377AO+7C+xtKbhtfZJSibRmy3guRWd6K2/RlwfL3SozkTxkHQrPLfu2r
KtOffCcg6htRfCpOY6qJTei5N4c+HbYTLZ3xmw4akjcpWvm+9XzZihLg96LsuKxY
r8pJjy4OZ9vEI8Fv5/U0FwRYg/7+p6wmCZz9D5zr9F9Qq8E2lYKRjrmLzpodae9N
UQjYvsaxpV0Z6B/FIx9/TASsDLYdGZiQwh3jToAcCZFAVfukgnUEIRY+kA9gtGFX
3JryXV1iGiaBxdvsTo4AirDLyHbW/JCNMvzFXC17YQBo+pt0+MxVD4jWdDx/uiVJ
VlstKTvDCgv88StKoQ7cV+CV3T2a0QxxNuuE3QkECK3NIrL6b5Ec1UmTCX6+s9fU
f3z1VC6BXjE0bXxbU+Y2xbpLfd1Yu2oM4TNgyqOAEiKwtPh1Zql+krDAir0G8gMq
0oKL3gVQyzG3HgVJQLKeNt4HxPs9vXULaixQFgg2qV5idRWeY/JYJws7kPla7/o/
RMli1cDIeL5mHlPxR1gZa+V7Uhl2OqqTk0v+PZMTWVIjC2hU3Egct36TRMZGKNyq
iHjgGJ5CDnBS2/g2JXFgyA==
`protect END_PROTECTED
