`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SaLDcVt8EXnKNLrpF5sbgElB6b7xzVa38fLuFEygM4D3
NVKsEJCHw2Ei0yUUW+h7Zx3oMnx6aSGbbTk08lVOJXKvD1UM6tCrJKwoFR5+imzr
gmKWu1AIuiGrxPK1OLRANcJ0U1FY5bY9JxvjxKxvNVOmX5vr8yIbBr64NtZVNqWY
Dcz9yQji1uj+j7XbMIeiKnDwHLibxUXl/mXgyqutvon7gSxcRMJhw5L5hhWjhwk9
4tZk+xWTggM+aZN/MUNryQI0xL7PJetrrlxJ9o7WOZGZIaa0fn6F9SD/Dw9TysB6
YUOaC2e9wvIh1AupLlAv2Et//7YYy3HZYKur7qda8KN8lKg4oulOWrTFl7HCI9WM
FSn1hsyYEDCgKfbunysTvpES4JFEteaMnO3sG9p13uv0GhSUwCSfYhMfOBr3znG5
NC3xRXO6fL04HxUYvJUd4OzZWa5rFCF4SYszFZGD1m+FvKIHqPprWvQzQAhEx+0i
gEMne1+LCiDDOLt3uAY0F3gQEbccvRKuh5cbb1qxrdDucSIRrFm7BBu0+7dFQ3E5
VzUv4Hz9fH+i5le4GpNjaBOekmUwKSxvVUWVHiqcAzb2jJIMcPMERVqhk80/FfYW
KYGcV3NFwvCnGailB9pCjqNV51FoGkppJtjiUGQUmOmm226Ka7D/4Tuu1iDsADQy
53QfySrHxOwnPkVW86ZstvR62LCY4j8eqiMbeExSpZlooM8rMnqQjBuFk16Dnkug
CEmmUp+HhBLlYMBz2sNNvlRsvj65n9HT8wD7CRLdeIR0Piw+lhnHuFak/doQW4Wi
Ovg+8A+9hlKoC+6WC/IVheBbViiWI5+xFBrPp9VxulT78GM9OwzHscGYQZZVIXkW
ZZ3TTIu5JbfCaop0WNZGkirXQ0eXmH2f5tbgu2MNY3cNC4zaiy3qYuYJFPCUe+Vs
HI/SrUlWLecQv6vy82tKT7uotqXCfDbqPE0QwsIDCpoHApjRMu3nyr3XZXxYtuYq
tFjmpi+SrDNysWjWh6HUtBWo4rrG4/lPASOfTP7acJ6w7M7j/FwJfoJ3WwZY1GuK
opUxdPlLdvBgxnYzFFCNAt38Ve2DoaffcTCDhZ4/Wb08pPC5x0HvRWZJgwNH12ic
RGTda4exWr/i7j/2Bq4m1EGdG5OaTgibXu8A7HpPi+lKnRBsexXZJD+rviL9xRC8
Sq5L2dXvpTE7gFOiuilfKjo6ObPBAloAq5+IcSczZlB3uNShlnRGfC545BxdFzsj
01+e761AHnhZ0x4Jlt1Nfi//F16W8q00WjywXrzdylahOjIP26JZYt7HQhL//8aY
XshRmHE94I97MkTW4oQQVby6iu5FjfQ2aqHJVKNuo35o2ZNzZ+fUHfouvYv0Dy+z
kb3bEUCWQJVpB8p3CwISjADQQAl2KAaHu4wVyu4ycXCuPfE4sL3d/EDY/P9v8GqV
yLI2dtAZHEflrwh4d76Zo2lGtiP6mlSWC7gDuyFy3jQlpYnfQL9V4T4oDct8DgSr
sDfWtQtWn9CZL6w6+oOZOkppAS3EDGa63AOCFUckhI8slyCCYl+Rd7a5NJ5axKI1
YuQ2aJMGAHg2mVIy1z6haqKMnmM5XXpNIlBJY7+lEyU109ySxeou6aMIiAHNTGtT
BmAncJdCjYpxnZcqBzbtGlqPGNtiq5qxHtZr7h5xt4b53WA2W1aHtgaLm8jwisRy
7eUErRLgv7mkmGHEdlzxHVcuzLJXEYTkPEFQFRazFIj1Scj231k5pjUpE+U8S2kK
oW0dRhfE9Ow1cxLy2/we7CuRpm5OG7M/fIfBC1/uKlz5LJvTtuUpOGZcPCd43CrV
6CVqofAxLU4AA4XPnMQNaGu72g7Z2ec+/dGyDWt8sLPIovQunjJnUfahRmzyKww2
+AAzzWOmo4zaiCQNzSsrWCFO3SxU1ruf8tGPIPYKPC41+dN5AQRiJe2B4qrZeVvs
xZiT9RVnxbp2x6IAdwym2L4uYxxx12oi6ZjZCB1sxAoRg+KHwnMU8SF/sP4Vvv7t
WctHL1RQtetL4DPdOkiveV3Ls8/qMrP8fsFnoTDeonaNS3vORvpMeXAI7iWC0j7i
vLzZRRt/c8tOmzC0lNEBMTPDNL54XcltUZ2BqC9VCR9tVVCRANIju4vPxN5BZ+Qn
bUKpq0bh4gBZ6SXDqm0X/C4LvS9As4tGC9PzYAY+TrgljOWOj5ug19PmJ1BkLaue
hnR5pvVaCir2K9If8V9RC6yGYcvnAbEhEWjtulfzJoOJjKgxbZ7+y3tmTUKwQt/E
S1Jf7Gj0T51yLJJLcCILYW9LoyWXN6J7CzoytD5DLSjAV4bXruV2xvPPCGaRHU+Y
RPwwNQGXqY1+tbg40G7vgZugyt8z8HG1DoaofBMhHBBteliqkwOMIOZR2WyO6N9D
YOANGtDj128N78M5t15ZDFTudUMHRWBJLw616DEqRZ+VS9M8u8tpNIPJvPtSb9fQ
lpKgL6qlmjWCS3Ea7ziPm+o5dCac2P11wYfLSCrzZYzJ7nO8NL3wlh0McrXMbwDU
MUWCnRFYud4n9v1awIJ5uRYmzcJKds9TR51KoNo7p88nR2vE+egvlit3tPgGbOiB
EcyLWMyxb/qj0+w+skh2KtKR5HaAOnYI/SzM7JY/djHBPhqXm/aoC/X+BjHHMZXR
dFDiQFy3+a1qWYMlY4aXJ2RuBLJVZEbKwwYki83ZMZdKxX4HlVrvR7ITzC+G1Gsa
q8QlnebnaGRCRIwLmPv45Pv7o0jpgkBFZBtion3bD6Uvi1u9Q2iWD3TKVToFxcbx
eOoHx9byNU5Iht5ekOazK9w3Zio7JnvFHvvGawkyPFe5S1GP7iRPiKG+VYjnI0qx
pcvvSJpanivWdq2UwNwqFgAtHAVRpDXIvi1NJ5xXLb+w/z0nkOppEWx3d++IN84j
1p0rZPZ3wVw0yL0fP05nWL+oaBw9ChepR6qLidgmQCy7nLInjqNOj2RQ3f8FBiDl
/ymW+Bf1dwcPdaGeWmssRoEBMWWmU7R3a33HxcIFwCMi/zF1ZJLNsZdqUI4r5jjr
fg8+j65SrLSnKx0J2ob5Ar+4My24tIPbAGg0KOC0NRnQULYUHbvB+cPH0nV1no/E
Ln1v8WMZ9F0jZBDHsGxOIKWlfWvso3AMt2e/Pc/WfXcEmFDmksI0vz7Nb3h1dmS0
WVYN/m2VW8OPEDFkRaARQJ3hwGgbeNfey/7xpuZHi3VvM8+zJ9uoRSeNPOwSiNaJ
/NU+iSi7ntaT4bD/v9A0/GpP6He81CtDSAuPZ5wj7cNswMXm6fZZgIBNmBgUJTtk
zUXubPy7zOsX/J8248EhkSq5WxOZriWXqvOlzkOpwpql22+Z1lfzDNPldJ0p55M7
8ogEkAsARmoLpNcPR1gnaadn8uqyL5RzKfqXCaUdpqKLt0M+DpTQDoBwwUTCSN0P
RlC7FRbswh6d5qHO9nXKvoP4TzgNCWnqlO2BPBa7DEnFlWyMSt8twhRFEmDDWGfn
eHcNOxmol/+r4RfQmjhAHDSyh17vYkUQq6J3/sptZyPVvXZg+x7lYC0pnt/v6bnS
Md4bvg9ddiZm8/5SzXDjtxLadJceFolTu7Ft9qvi/p1t7IWJu0LiF1d1h3Az/pDv
+Xz/d/MRid2lKvPoD2ujC4BktiPuVbvLLWFOkLlsuzl1Eql6iGRHAg977NTAjxTJ
uFzOaw3eyUMsaTGf8luqgFtDx2op29Lny8L8lBy87dBmRmEdyN+3XNYStLc3UMm3
9DGM9QHphwwgQG2yZRLywA0LZOuoW2O0iEFn3Bn86ZlurLKsDnbVRCpnlGeAisSE
z8C+kHvxKgvCLu944Af5C4o1ydQXaD7xZocq3PM0VI4vM76oziVNNR2hatwe6RsL
M0twh8C918urxEaDgog8KtlP7ed/v3OUnenhcVl71VBK8QR2yqEpnSHJ9qg9j+GY
qKuY6j87Jqh05Ex9mTwXyAeleuPuhwqd0uIWbYzq6ORrby/cst8nWqs/6SBp6pna
aMc5WKdmn8eFOO5JvLusDf6F2Uu6hnQCaR11Xl933qZHr8UyIE5Z1gQraO8XYmvE
f7+ojtlcb7hT/le9mgx2AOArfBGacAA12RG43AuqdMiyQapWIJgZ0AAUXf8RMG+l
Wf6kWyuZ0h3fH1dbsgg/H0KvVRh0zIVcSgfpmVUmOeuy/iXV5LKX52v9ZHDmNz38
WihxZQaRK0viuwTm87XH1GSE53LKotfFNLo630Ogstxst67b1T5nqMlNxr/t2pGK
VGK2BP2Pz+xZRURpKDh8k0l3zkATLEPkJ9UzhupLt+qi99H48AjfRlSt9lGYuXPR
vsd20ge59STWfP3LGlpWFrS9yc71HCkCdYWC505dPdxAQdHqLc55Up7/GwFuTdt0
2uaM9r2RRAmQDn1bsp4sfcTVbtJDaZUzEVUJtmnYrQzjYZTXDh3tosBd2M7c09Kx
gyimnHfnrkiHK1VyfPo5usly3LuqvPry+TPvdbT++AAA8h6+W5169hFeN0bnJr9y
XItpLBlErBnk2L33Xz8eal+m3N987ytSKQ0Diiyw3/LGXuje0xCHYaqf2Bs0G9Bg
0JdUQpNNSgJbaki8WezfbY5e7wPWNp3OCHFwX47gSGwFN0Qdi652DsDVkzZ8f35c
yEpxrnb/OapH94ia4DbosBa+1/uuKnptZ32JYqt219RNzwMwCthkv+XaS9SPmDKe
BjmapLbs3hT8WCLCKTMpN5SxFRz2n7lyIxCNYEsQ1+jNdEgCrYoxrbL1aeU+WZqb
Vfdo4mLxeyShEgrVfTYn4iEh+S/JDFwjSGm8YhynhNFO528Ny2+IKRK1BpjAu3NT
DoVbk+ErfPL25K3vbRuZs2UTd1xN8Yf+10eeFPyA4ePChSReTyG+3z4jbC7ACYX5
3fOsUZvvy3hGLxL3o+IimRax+0DHE23MMjXftLYYJm8Pf6wxIVvTsvmNrdq17vi2
A9yi0KdU8llnH8C+vaXGda7or8ZrKz+QRhg+JXxSKzW/t79XsBAJl2Wi7Hx088r9
ob6l5ImpHVARELqmWMSmygYePudfygiqltgD5BWps3O1dsKoLam5otuHNzwlvD+x
ZsgoOXk28vrd0SGPKlqNpjBzfVJPMNQL0JDQU2ysGCijgsnphz599BV/0NiJkKnz
eS9iqqatHJ+BeOEQkxPvX628p8aSlooqMd+d1nHqR3brLGRs19OPzyyqg5ZNyZd3
GZPEqCLAqb2/Y1FESlndY7NlQP0uVqOjPIPFr3PWefDkmgE3PQI9r/z8jFOvQXPb
KihvdJl5twkoeIrVNNHbiNf2cT62q60ofqA3iCyWe/jEcr0Rxv4zIARoc/K/jLz6
tWxb4ChFyo34MKrEVHqt+JlIOtdlFUciZEm50vY4wBNpmYN1x1abE4VYxZtYv8cg
JFwn+62+vtZhg7GWcGMtZ/ODFTTf6fkcUdwZo9nHiVqrWtPcjdGQe5EVOiVByr8N
nSCIbcR7ENHlRfU1kkpy77cQTEKahsL9jZogh+YTqO34DRveTlxJTYO3pTVW65cJ
lJBeaH4nONv5BYRWw97ckY6kOAnRGPT8qfNaT690nin+SQY/NKqLjwW6ubI6BP9N
pqdT0eK/Vp4h68WivimILnO9KlAYZlqamcBQgHakiUhNwCdVfUsBQM9j8LnUYGdc
VInSeDspFbhW7izJvUWMd+Bcx2e7OrGu/yoobRDQItUfWbEs/YfOERx9Ux3EDULD
RAApoB8L7SSdJtnvOoFtMII9DhJvjNfnltapJo3edAck+X34ExffmIF2OwPoPcEO
phq5Yp3e5C5/q35LWslUOGK+OuNY49pGIIhYTuxcxw5HeGrYb2DYl0/3NctlqDbU
2ZOtAQW09Km8qM3ACGoOIOKEWMI5sDdz46szpIClUR9PA5viqmfifzJm1U9NTokH
Dtngem4hgSc5QgXrkiaWLP1sqT5Ol95KehFbtLrAUnejZ/gmGO7nqIkhy6Jsxaws
xSqDmGqDgc0+2DF3F/05Ou0xCLvuBTN8UQejItRcZq3jFyEExd+gUjx+cMO7HRos
U9y63LEO0STJXvYbghHaVOYSnJh9/w4KJwoHitpeJoK4sUb4aLk8+8QP88E/8R7M
d72A1v6r/Z3SOrIBIPjfHmaCTZn8x5TLjJbaQ8nx/IGOgRTXu+fmAHj3yH/Bsezi
utEqh8aw7b8+qLU7RpVhH39ghj8CrDfh2NLgUDpwwDp1uzoWX3g1fpE/XLVS4otm
knjc8IOvhvYPbubv4Hbmzkndr/Vc+HAFI0hSSTK8xbcMCTx+nsd3rK9k36jvvP9P
C+h1Z1uzMJn1BnTCkBaPvubVl4ov3rSEs3KD/R9VOpGchy1pR8XJ4+NCKsfTXWjr
yXe+sp0Pika6voIcmdT0im6xhPG/RiFW689DOyu8roBBDuGGqrBTgtiB+2UvfpNW
Cd4QeOgfYlYVmHAIvTuxswQmIvz1qARCmL+DcSmP9dSL/jEG9wTQYCCvA2bCmoJT
L1XDjHttKDP2CuvWxpSkeE3EKF0MyM4ZtNrpPSFrVI2XoBDsMeUwXkv/Xywj1Z45
WvEXzlz7j+soYO+eQ3VtZDDh3m0QbMY9H8Zk8mGBSQtef6C6xH4nozlxt/FuP4hz
iq8kxD1GmoJKNspy3nk+a3476QnmbT2OhWOVTAaa/dvGiLv8i8JpTyMyM7kIL1Ku
ja64gvUrY64p/Ia6PJr3M+fpoN80v9xoP8kWb2zAteKWVg70VMgrKJpNCEv2oZCW
pqf7VtjhKld60Fd4fnFKItN6ZbqFc8KuCUklJe0TNxoH7UNiQV+VPNbdeUgKQ4Ir
uNLSyc4LqoaGnmfH2Ahldxkr0R+HK5yvSKs4jPaXnfsVZ0Z5C4DfaZB0wzdfX08a
rhaO7dbwRWIBI1vPAbp22EhxIXP1GkA2XT1Ch2awe2LakvI/K1177LWG0Su/9AIA
kbT936LnQTryjyOYNqmihGpIQoX4o5rpWDep1XEaHfjCM/XQIlmZtVD+IYarkMqa
ud0HL5SxhJAFloSHWgeId/WnbKpyR+KXt0Bnll0T+2/EN/awS26m/POe0URoFMMD
/0aCnp8FLgJLyzGK8rsTRDSkhjDxuijKI7jwWjSqySRzp8DSZ8SliaEXwM+393iY
rYlvcHNWsWMiJtbN/sYvSqIhbo4+zKBp2+wZcrtqDNp1wnW16K67Z30guAEoXzmz
lb19DiHG9SV94FfHrljnq8NZs/J50j8ta3ZDI0jYR/H+T2b81MAE7ZFwurWjusU6
UJFSTIQ603XsswfBEbePMSIjVxNwUx5XJmc0LeEOMuAsYGllOMRofQvpiZIYjHb1
uA40KVRZcdRHDsKgZY/ZtgeBaToRBaDOPFTtHmcood6J2FDNjnj0raRpuQiQwNzb
QRKsOBtJiY9kstebn8PR6dAa6yDxk+Tyjp9s8my+BZsIwv7G0g7sD9CEWtcsWxD4
HODKhh8EMfsGLHVT4tdXMjd8RRlYDsIU5hC4Cc7pMsXA7CzB7JJU0Q1Fj6mmFsGk
Hy+/IShubcmdVx/6oI130TTIi3azcoABYHE6N4EhYkzUUZ3KveFF9JrXAR97Wws1
FnUbgAObjGJOHE6qHaW00fQ1CCe96Y5LgtaJzz7tgcbpdHu7Tv946gnD3n2y9V0/
2qTpWawC8Q+xYxy2HtKXtOH/iLLH5GeEv8nE7y8UOOtPE8tm2f+oDDcJODUuAhkF
s1/zk31Hg5adPTSURdjd5Wcv9oXYh0VUozAsk6I/+D1eBEYk49+dMLrYGFutGXHr
fZSUidwc3eZO3p67YBZZ3KoLPuHjLD+fje1hs1O+5QfhO/fv0mjcJt/LJT20PfxZ
zk2bkDvGeTZ90cL+nPq2NBnQpt9SjQRuqS9cYquxoXZW1BTufVKyYWrPMjp/Y1EH
XD6iwtL9mLWxNB0LthLRel8j8/DejnSiAivft4hRpjwciSTjmCXBZJ5kI7k2dFQz
nH8ptzPmtvvu7n+0TJ5XTUEgjXb/lX1ksfm9DGRH7fodMg/9ftsmi/RKP5zRfsGb
HVTJTY+kyTjpWVI4fhfkD/GQ8+squwNUWM6LUTtMn23iCArt0z0d7VPYCqEzLgnV
KDoD+qYH3rX8o14tfnGH3cyVswHkyrzIK2GDu2hOY+oUXK9J0r0Yx1aLnboH3GkJ
Kw7AqGt95uwNmAp2o8cbQSR07AUOwXgUzWeeqq6z2B3XAHmg4BoTYTQ5+l38DkPh
//KQoCNRIsPMAe2DtxwYypC3T7D+//Npfx+AEIiVOnHM5PIbThFkbBQx5DDK6TyM
a9NKFrSYtFtsk/Cnj1U+qZ0Q0RVVtlUXk9U3H0/1EuORwXvtNftJriO6IErsm2Bb
p3KjqmyY7SCUCYiR6QqgH5H7MazYgBXNrCPS7DZgezoQ2rfxGUPa9Gr/CJjJzOiy
KQzjreq3Y1l93oyutzUiNPQ5ngLtu1Hf5qR4/Z8hYdl1zZbJ/T5oZo7jiuTAVZfj
vJMEVfYcnfHUGkLudN9oTe9tu5qJC1bY1szA454hFLCYZZSLXyr1XE6f/6GoRMyV
ymoUFE9TKUezKPQuK4VbZtp0PwqrqbLVNXcIuijNMgdJxAY0j6V8T700VRaRL5Vk
97cPyY/t1x14MUDPvdAEvQ==
`protect END_PROTECTED
