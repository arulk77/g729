`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLDIzUJviymGnnueOb8XQuKdx4+yIczJcNEJDdz++z8p
lMh+9FuKhLJovrAAXnDq5tXmVLwiXnpk+FUYQ5i6XvddCl/T/jdGAbtkdSS8JwxL
HituU3tQxSzgjIT2t+D6DplJAnfZNZ/h3Eou9+HRsIm8/kTAXgHCrjaF78tuvyqp
KHfWXgPdAQtC6XHzoFDofcMjKxfhwa+gMPCbFxpTqRYBoifX9MxOrzs1NohXBL6k
+KcKTYoNicpm4GEJhvK4Qb7dX+3doPZf3SqpcKTAYngudK8Nw7tPvvphzni+2faH
gYYf7YEpMOvKzSvfJb17uw+yRru3OO0+DuwX5TTwK1IDeF7XeawDjq4NlGY9iVis
84kGiVaAV4Bj2X/mEVTr+OJop5AUyFyg9I2rqmLm83qRSLhy/uTdM1MgKbHtNXC1
29cXi2/XJ9BAl8SldP3SbMDiqg3FuCdeCF/NipbcAZqZTRHqCPCBb9aq6jXrWmeZ
lkkFFL0Scg/MZJ5eoatvLN5EBPIPoZsZFj2aOvksxddhXatzJD9Rh3HrNOIfP/kn
bhHgdUwHEiv2M7KQ60nyyVz0P6a3TjdgIC0+eBCeIlF5EqigW83i+JrfygTUvMcR
`protect END_PROTECTED
