`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Q064xpZucn7/1GOSQ7+zmhvRCW8UN55r+4+v0l7fBGiHCXKksX3u2i29COcXEOqG
59FANnN00Ha2U/hXSxN+WkG8XGdP6wedwtYBYdSA8Q0qcgQh2QxIFjeobmAFiWJ6
CJVoJqs0tzTdOCBDVxHNkJAWSTMLzouoy1LV6kh2pzHJKTKlvuimzyYjJVD5nPoV
yKjCM2uba2B/SIG/hXFYnxKrYJALofhaUBKzn4AeXqo4AWBbI3SEN0rIcytQGuEW
qHJxtYf2/l47//AOp4CwqMuf0nnWrS/XsS80enrDZyuFHqg7sEBHia+lXLYMQhNd
XgxhZ/QFvykvgGIdQ1oeQGF6MqjwZZ4EbPskZZhLWGmUQOtvklAQDNSQsedo0IOZ
Zw2JaniSEAzVhxd1VUR9CiS8R77GgZ7iYiGLiKAqkSywi+IH5Ets+NYJ29oeu5Xk
9Pus0Vpb4VMyK38sK9vhyDCob1GpWVLg2PqqDplmIFM=
`protect END_PROTECTED
