`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8ScpNhBxd337yrg5iueZ7O8yH/8S70PH19kNw6dw4p8T4
NjtQrtIeXo4GNap0DJUfBbbauZAVec9KboUKXirkOhPKEzEZQL3AbeZYQ0vmVq4z
tU5TESo7SSzHcxYxMzgTxbgVbBEuQQYWCEjq5S3hlatvJZNycqoPcFW/sa6EQk4t
Ytb7R3R+nd4x5tIgtqInSZoWQyTX0X82yCxuPr+ghTRL5ek8LeEItdtrcww2wmaT
hVgmVjshgRrMBJX7v33DAOcvQV9mMshotmaRzTRI8Gz0JCr2TNdA76OZG6Ojm795
mnuKa9NcKMnwWxoKVayyN2CCzKFLXJZZsCWGX/vn7vaS8Rh3v2PVN457cYDDfz1d
xt/a8pA8x9P1bDhZLxaH2Z7YXA0k5s4nBym2bQmllDzgdivipX7THiNfnCdrwvBJ
NcmlzrDtHmMRA0NoAJY7bP+FdlD3oNKWFttdS9GF8ri20ziZfV/XeipWhg755Jpz
+4oYSsd2QFaknZiMZSKClYaX9XzjGla16CiEspHlw2JloT4QIqcD8zO8BHarWbk4
lsVm0x/qvY4qhynZ1iITQ131ZbZB01mpKPgPPpD9qd0pkqi3m8MDJRzfLrXvyawx
uOx5Ox9wJTF8d7X9z3ao9zpxYZtyGRPesCeb9smRPzJYSAKa8K7kLYtHCFSwkXHS
l4cbrvqTEb4ZlcdR1Xwut/wm0g+S3rxxGTCIUqztUoWwAHAX346AvU0tTvt8shcA
6+o0mgIM2I1CxweeydZRpAXgVC/ncLjskKPH9seM/soDoy81IhWk4kfvo74hRw1I
eTyxJd3zqbZqchzI7AJ2+PIR4/yfY/mmWkn6KjZt8y3/Y5UqGrgBHZuOuvSiWYqT
5099bo/6QVTK6aPBPCoeEhBPL50FLFIWU2M5gkl2ITU7DnCr+hSKqVpjEE64Tj4V
zCheSo7kxQIoBarBePEV8WJyWexClSTEn6zl4vb9D03oOWLkFOMYX7x7lMW89Q4d
IiUo0GDYzd53VlmY6iWluwfwsFKbzslYAJu13qhF9p9ZB9XvNIyonJM1f7dI7rp9
9t3anLaY9yuXLCkdREEhiRLzmSWS7f4rlS+Pdr67Sk2O/7xLJ7eAVAsmN79zC3Kq
E4AFAMMgXDmHA6bDOKN5yYA4zayKBZM7IloxyLIdp4xLPFbbGeJnvN36h+90bh/y
2YOLcrdvh/blJ4AMwAWbsBYBqOCs5fvnqp476iGfodiWjUYhJm/3lGahBjq8tYYB
GuJltr/oX8Gh5ul2nfJDNg==
`protect END_PROTECTED
