`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/t7IxVfK97stk/yojokaI3lyz+Wm4KgSTiZ2uRahEyw
gMyxEoJl8uenazTqUUFDFTtqVuPQ2nmYeEEKegtrgbkBEWYEq8ekffNTFntsiufe
bQ6DYFRnN3xpvFfKdaOJg8qKtCCQplW0m8U7C4Sh3jLMU7qTq5GKf7gCfGzd7YS8
FjLvvfz24X5GhZL67uuGYqV0Ahgx969M+HZTC8lFYj57RD6auu2nrHGTc162b14G
wq7lHnlc/vfcqGvzChaClG3HuFRCuhU2qaDv3LnLP+KK0yk+/HPiSEni2GSO30xa
e9DzlTyM/RQ4bHD/yihF1xjzTDScuxRvsRj0chuTbUDvPjL08lmhDZc2hwtwauYC
B/JDRTWDaWE0uB4kMLZ8uA==
`protect END_PROTECTED
