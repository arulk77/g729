`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN3jF14HdD4nL13s1WxRd7+TFD2AYUCnexCSJ1/pa2J6a
OUA3Z+FSj71W12OuTgdRfvYEHUS8F2ywOtjWm85jd5eEO0Z/+zjkoGo3KmP2A08l
eHQmMjDqktSycZMSam9kJPJbx05Ghbf8JwDxFWHudM7zgxTZ0Fgghfw3Fq/n74rU
Wbtsc9i0gzN9bK3Rf5uRAYgHE26FZbx6bNI6DTNgyzAV3MxwaVtihsGj9HekdMoE
hdaHDCf9G/OdTujdKk5ucQI/jpw1cbBFxicfQysBms/l8iyrjbKFrlXV+p2zvfAB
1IxjUunT8YcgLQj38EnFT2a4OSp2tA5iCHnWNgFonHP8JQNJMFPshpTWRn/zotu0
gI/hxu7fg6OaEyvkfyU0CUgFlmI7GdY0yELFrwffPkpvbMQf8sdKpP5ynEa1XFlv
lvxFj0Q4RLqw0N2MC1nw5HJ37Jbxi+h0kmHpC9QYwdHOosr2UDX45MfPfsH4ZMpQ
43SH0czq25pg2ENqjkOOQwHXdBH2FG3jQvB8jB8nioG3rc+CRmZes+5mAzQz9oC0
Iv8D8WaP6EVzb60SRWvuGyVWo/ySUoC+3UhC3gI7fCDWwp6JlWmUwIix3ol0rqgr
GfhNJMpM2JrclrcBkaHRrC7PvX01l+Mxoz3RSYHoQUNb8Z2Vv/5WVopxKeRMr4ml
blD/i6YVflEhNH04YY+74BIK6bt8hX1izbuUVhOPjVqC9chKS6dC5InXmoT1Av5t
YDNKk6NS+Jc1qQtLNznbYh0Y4XCI0ECILmHTq7A0veXg7jxT/D0obe4D+zZE2/1d
Hu99teZUnENIrbMz0cQ3JMcLzThggw81WiEZ23c9LPAdxrBlQBrcX5ONfknPae/J
w315+uU3wJYFkQCW6W5Z8TRV1ue2bV4QiZ/0D7w/HF26NnXYIc3+atCxXLoaWxrU
dp+gCoy93BF5SNd8u1ni6dRKiSno4iA5iriE44/Scv6VzFO5+lKxQfBqF3jEc1rV
zEjoZzi720AwGoRKEteYmga/35C0wrKjXrHiO5LYSt1EmEp+GXercWiAnF4JQTEz
LLlwuombVy252gAF4UOrT28QS8Erb8+feuYf32tFx0Tbts2YeEnadMl0P1pUiI+h
qwjgTJ/mKc0nkIeG/2epkulbgvCtcqUVeilgc/Bn8yCUrvx/OspusqjlMQ5dC9il
x+VMAjZ047IpyxkccPsENNcMGf5LWKuhLu4kzVBiDGsXoV8Stvq+wI6tI3Q0P3U2
XCrWNIxQgAfB3e/xLE6xiNtXT1TT7hNCbBKKjQDm2//nPfu+nZVDhJIvdGDC3Z01
PVTI5sWrCYASQ57Xae9zTwMR0dxh4pM4BxZ04/bt7HokHpCF9uohnq1w6C8PmDEb
SyVgh2xE8Dy7Mwe4A3gh3A==
`protect END_PROTECTED
