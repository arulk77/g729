`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCHdHQDTzBpvWEYXUbIPNgWkV/MtncJcXEfDkMX+8urH
TfAdNov6qnFHPNkiByEFWtlCqgVfmO3UcS6H32KyOg5v7ocbDbgEQDGQRwuKmpum
vtmY6M4qEgBnp3KQqm/wCP8MGROh7aJZHQI/2Kb2Vbgo3PBQK/nsla2huq7H91OU
NzWKRNZ6CsANjztwDv8SW4lHr46mROtbKlFD+KkcZp9u2h9zSMTHy2PGUpzmVoek
h1fFD4hJaVqAPkRJ0JrWX9YutGD5FZGp9EwOwTG0COHDUlHfkGfMJK86EVpGZQq1
bcg004OShuF1TbSGu3d5ZDq7vWehc4Mjl0xunCEZvjsFIwG40AJsfL3xxCIlu4Yk
NXXJpkiYI1vDFIls61EZZjgjYv2unHucwHgPNwQZfCAOZhBwN1ed5MGVhu/04BpS
GzN3Ln4FyZRYK5E5bbRklSWFCx+6rb4KAEhHQYlHX/MM7Mk2Is1ZwiqgNyP38Ngf
zJlRSiDXNXPnOjKDH3C5sUC9ldvwj5ZpGQ+qGPB2dvmDdfJXqDruFN4zYky8Cp7V
khR0NWABxQd71uvpyFxDzywzls7ptt+dhvHS9pdEKBJsd8QNkgBQE5GIE8nW06yx
JkfEMQGmLrUtWXv93/3wTJZ+TWTXldmOFU54miXMoiGF6TaSUFF/CvykBhlbRbYZ
xjtHwpcGrKl/RKzUgzXNVGkvoVRPIeUmTD58XuIMhpsXkjheXmB55dbtVKa1aEM0
1oVNbSsrR7ko+9KiE2N6GgdFrjASKq48vgtVjSykEO+c4bXaotVV80rmVhMb3ufb
va3edKp9Xz3X+rSjCI3ryxJjbJuRztUPILJ/8j7WQnA=
`protect END_PROTECTED
