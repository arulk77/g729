`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOW/0qd+Ptc89naLJVUdI37872AQtrndKdZT2sCBC7Yx
Ca4BKHFaGyPSS7D2OaVD3/DfgGxNuIvIUAOf2osHnPDQZW8/rrwLFaxz1wlyugD3
fVS+3+mL2cpdUTe88BdfnTwT1YeINLeyuXq24m6tYxLECdf0wkQ9J30uJPt78n7w
bNBOmxaGVzF5tWF6ww0v9qoTLud/+eOnA1fUpcy5sSStJZA+QrTy55v2ayNVDPth
FxdwBQgZIXRKgZVUygr2BLw1BuSTWtYtuHhU+QaE3we32Bej0YOZQPLGPcy6KKLy
9WobgUEorUa6kI7U+zOQvg==
`protect END_PROTECTED
