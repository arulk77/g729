`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIhkl4lw2V6MtF11fjmR9OfXdBB81U4hva+YbpnZV6jf
Co7NWiLzqko1yaEvO+1LwVk85CkkqTDIQssJhAyH2NkwoZn/aU0QeY2NYQ1fHgsI
yXovKtIdbrN1JmFMTPwsvSdicd8dCCnGOBKXBCSHJ/CDNvDupmjsIeFZIis6HJLy
2XjJBLQKEAWp8CONdiPoXA==
`protect END_PROTECTED
