`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF/TO0N0d+VzgXzJqxrhGJg8qrLSedyTG8ey2GG3owbJ
sdF5Fj67QPyaT6rAJltMgECjuRajwCqOe0GWvyYnpK/OGV6MME2zAhYu/oGOsVd0
Yag8hbfnEKvQceOeLthyoih1pn2sLl3ClXttQB4pvc/+CVlA3WtCfUDudjFPQ9Bc
WWUTUV0OAOOADj2/pplMbg==
`protect END_PROTECTED
