`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN1ZVyl+ofQ7DKfRdVD/xIRuihM6qSF3ByoDizcI1Ckv
tc74S74NZuLKI9WqVfxAkHiVxJdm1rUQR0Q0/9sjX8sjY+94VqMImcWk84rsU3Of
bJD11TNtcl6MHxScLOq/LMt2CsJGhFIxIfxR1V4/BynIB/pleQMjHgk55iwv6V4S
VkgWEgTasgmLBNTd4zC/Jw==
`protect END_PROTECTED
