`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDMe1neoAEdC87RmttUad39hdHJQ24OBM4WsAQ+Tuw0n
iKMMSTHpRq11wcthcsAAk1OxxREW6VK5HUY1H6HrZ7R/peRJDGpzKUHP3wnzy29o
97MdS9ocUYtU5I2+/KWkogcQxlIAg/JyJNGw2i588ruEcciCIVW0rMljMbJRSj7R
lgIISPcANmfwgQrp/FKduCo+/vWVGQA7eDLfqrW7t1ZNoQp5dfbdN2IBh+qj6hjc
8fzbMOb1NQFtnJ1i3ROkNoJZeCyg+gtuZz4lkpwBXoAigkwRH6/z/Lx4z5pPr4DI
jXW9h2uuwnMO57zJvlru6EH8bNJsiXekXF7FPfAB2p0u/2VNTtsHc8j8MRkaFpPR
Fey9x1iS3OAlaHy9TQeBbQ==
`protect END_PROTECTED
