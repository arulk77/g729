`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAy03H8BrXXc9FNpcJD8tneFhwkGMwBj23boaKYM3z4h
b8fZDJLTrYzDLeNpRJYH5/VTNTtDTdB4E7Itdbo20jNZgQJKdae4RKXC1gG0Hdg4
YpXF5QYkKEfUAeaqVw4+i8F/jf9hSGb1/7/Y7s/9bceDaImH5jhr8k0xF3rOwOlJ
lClAhPht/ihtXGa8qQ7dN610nAVwLMtwox0B+mKBry273+x3zOJHrsqI3R3vXiIZ
eZwtq9v7Dtk2h1LvgS1JYUXOt0HoCcAwJGdUQxGOFSWTjXLEUCiDuVNjYoSd2hvP
7oXm0cf+hldTZxflXoKLrUO92fGWrTgh/dXNDa0vN4WE0WWyZkR1cp5fuVOMJnYg
Ocj8GmialhdmkA7tf8ojyGEavC0D0UvtUp3mEgApQhDYuzrQSOUFDHtIpqgD2836
SSZ3D2KNh+DlZ+Kty4H25UV0fY3Dj1hMexuEWobn5stOA1a12kxSftAEAzV4u8yV
Iru6vmpHOnQlc9CDl5myBfcmZwoq0HIhjeaMJDkbr1lfKY7oPKf9TeMmvl3nirEZ
`protect END_PROTECTED
