`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDrigwZ091T47PSn+SIaNlGLlUapLOwa8HDv5eLbkWG7
PEb8vIU4CM//guo7QfNVH2GLqSZI3LqmIjYR6Q7tLlWR0vlZw2qKWgT1+k/AWJRa
wqPrQrk8nT7X4NlaeYFE4RMA9sYSZe8+Mxz5QnQ8dKoENAlljPUzWTN8EbDLQPYo
8vjByTrgw5HxOXJBkYpim2iGjQygRjsE4xjkuOskA+SQFuKInlpC6StcnVD8dOg+
vzR+D3SALTzTK3qk3uJWhuRPO292ILvyrtD5nS4um5jz67GimAoj+ap1j3mop8um
me8YkDh2RNiksaljsmSdsVbPKi2MasBunV5VF7oBNg6/pvXoGuffpfveC8Nnzdvs
yZpGP0l23b6mW3T2VOus3j4nPY6Ge0Y4ckdTS6t5syrc3VYdr+XYBq9gXpNj3fc4
txSZaoLjffYXzhB/6MNgj9xbzC055TEu1e8jn6E+1WgZJB2dUBdA7lA2oqtAZwLH
k71LzZUvKqDWvPYcey30uOKd1P/GBZSxygPDWLlOjhDv3lCbts5HMwqs2H/ovGZk
B0az5H0Yljl0nOUDEnYQTnfSUuE0vqHyhjZId3Pcwx4Hmprsb9T0KEp+p1K3mHj7
kUs59TDagz3MUTpDwQY4EFpAbGmr39jsNk7A6uLd5Y1kr8Mq0B4jk31LwJ19oGit
jUfsZpKKs5nW7PtnnQa7Ew==
`protect END_PROTECTED
