`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
PpUBwPTObDEXpd6oVhn/bzvpXDrH2A0kbi+OI2OccAdsV17OS3MYrfsDtxTeFK9F
gdg2tOXVO0Mx5q3d42f6WS3ND62csph223s9ktY8Oha2oszTqZZ05vYaTj7W2dXv
i5Go6CgG1/YPsMgxVM1LyPrrJ7i2utz+korSsW+2cAkbZFqkoZbx1haMgfCgtsNu
c5yh0jwtpeymbNUGaI2tLiwDbLmnQ3+jTMbr53BJ5bo1QONh1IjnEgmTn0LOLJ0D
aAxvTLKJ/hQjzlOR247ppWC4yWf6of1uPRIIN4BDEHc=
`protect END_PROTECTED
