`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI8zSHU2v0egibI4D27mevlrIm3iEHzOgJ5PwMMYze0H
dttXTjd0Fng8yrRwyChtQ6c6NPs0FIw0Gew+A9hsr2XKiZEsXWPOrE9pZ6/QUUQv
txfY78sODqUK5a04d77zvnIDfoj3ClEdp/m467mJn4b2Pvlsn4o05+LsrYASVZFW
B1uXjoZpTBW6v2uM/v4Lz8uIrRAhJfVvLMd8DpyYFqNHhbxSSSbC7HXFISUbA6sG
IYdK50wMSwDt/RT91glOqxaM9ry0+YUL6GhwiU2EeaOnDdhbPAOQ+kyiay7JXhGj
UB30oeNiFHWlBEzybdqG89uIqxSUD8tnjKs+lnu011iwkv+OSXr3okreAIkouC0B
Ylj6jBCBgbsXCkEyYdV54emNnl4BSYp+L+z9xxeBKLLx0fNC6ve/R2IM8Un9ECHA
AtmdXarLUAAr48DH/7jXqpc+2/ibADpJPY10jZ6WrqqcgwEVLDnr3JIpJKmwXMaC
zs+Pa8zMgWvQVQluOoM04Zv/k0EhEfZr4TBGGG9gm3yGIXIK06LUZ2rABu8Xaewt
TczWPaBqNoO2K12xMwxs3foYdTQsK+ed8eTlPCsacwpXmR4i2y8duClDL5i32Rj5
zYWy5s+GsmhNeQCW351fXK6VR4/HeOuYJooP+AoRqNvZAWxeb0IqiEU3SrYDjsA9
Hdqz89vCF0GrRvyPqmuqcyR4S16kmSe7G5tX0Rk8+7/XIM4jow+6DWBeXpNxNQhq
`protect END_PROTECTED
