`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48dk6voWlcV/Qlh5OS+FC1biX6daGDX76vjZ6fBuWger
q3MLH6LtUCwDRfrInhLIsnToLIbqKXWxvIwVqVql5xgLgmAoyr5jE6rnmqRAiq7Y
xqaeC+6AGYP31vqtiHE+yqhccts7urIbFRPA02A1bT9XZzXWEhQ4Unm5v0BNroFj
bONsnH6nzA6mYqEuWbQm6i302Lm1I8qvxHG5HyKIrLk/ucXXM67J/QyUXVA0se8U
N6aieYHb2p5HprP73/0rO7Un8dFlXnAoG2QXo4ODanYEaXLQQtwk1giVBDfmGNOF
jU4kwkuA4fUK8Tzhq2JUMyywF/7M5Lr6Ick29uB4Z+DVrxlt3o8fo4cCdtqKycQV
eib/8kYKSPtvHHmWQZ3kIA==
`protect END_PROTECTED
