`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/VwebrcMfJ/thDIv6pjva3Fnw0gnS0wikoRpiX1VO65
x6cXUARaEVL7Tu7NwjiMCGxqgtFnhMVA69sVuRYwOboeZLzeDZyLOBJocwV6bJJ2
EjKWsjXnkDkX5WaVso+kcQvaM+/77PnX581FRB3tu1pEGtkhSbnWkcPNMhVLWi63
2hiXTwuopawJD1q9Vpei+Wf+NPDddHkZiO80bgqcdRHRNjHJXpaoVuR9E3iygbG/
OQaadRyuzK9yf6zAAhIUFxbjUwj5wsQyc/L+t/bHPyY=
`protect END_PROTECTED
