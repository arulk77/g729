`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveA2JSu8xPA6b36A0v7aMVKiB09xGPbImcVS/oAzIfxs4
QOkfdWsRe9qkWQZP23IV7ayYaIwD9UsainciQyRY/mg5jXGaACMDW2TQMd1mckO8
lQ/81XScQ32TYO88WAY0qnljMfIp0zr6bwOlBXtMefri/WNKJ9M6BJxAbwC8oXkD
Ub1BGMcyEMDz+H/tXeo4jwjkqaql8IhT5nSOP3fa1ESeMm5Aie69pP5jtQKE1AxQ
38f+r1+nYGYu+MV1CmsLCGAkzAoNKl8xdCQku+GbssCfPMY9AlJdzNi6t8aRPuk6
ohm1yMmLpi2dF2Ozpvvd7vuMBtH7JiN8Iezk9WDnDzVKYOfEjW5FZKO4SbE7Lxhp
HMPBwdpiE11Fo4/SM97l9eHt8QZcM99r2SffqwYpWqYEUWX3H8A45+mJlipnI+Kw
vqFwRlhzONsoOW2jRuKeIqukhlGTgOQVcJwItxaPVvpPJoall+DIrOHseHnfNs87
eyvRjawIoF/29aGIh1XtiZqclHVQHP3rfo5hGKOTr2Z/xAKPxtki4EyXHYYcTDXz
`protect END_PROTECTED
