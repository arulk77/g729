`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49UQqksgk5pIPbqS2BF7GwErdidc970FsQMuveawSdRb
UvnSsAcaZpwSGbT7Zq8SCUWrgT8apUAzC+NnTanSS+AMJ83RHEE8KSk/3l0ul/Sz
lYrfM5kCm0a/VYbf4rdMSSbpMQDISyPdQdOvei21qWjijtDuE4wnsTkF/0PAYeqN
V9mZkRxC80+N807sUVe+/pIhJ5VyUgZXTDjDZr3eAjcBwbhqmqGudOAU3TZq2eOP
cmVS7Ezy7GPg+ychJRfS7NdvUCUwTMjV5Qmpgpx2+Rs=
`protect END_PROTECTED
