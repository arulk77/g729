`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
VR6ocQpY6dr2GjpOl8KyUb/le/ytvlIshy2qpb9AE++IwUqw2gKDsXHyFS+G44TK
+ntN6vMqlAs754A/utNFtClJHLHvx89Vbh5lSJg6eMGZuTj/We3eHYSZgtiClnoE
BW0HinlomHkMhMttunJZFeA03Aiinf3W83RjYx7OQezuoQTdLWlg6eOyZrSNYaXQ
Dxqrxr3VUlS80XXvGXY+63oe93Pz8ujzjFWzRUoeLag=
`protect END_PROTECTED
