`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM3jbLp5VrYA/7DhGRkOQYfcKCUKpqt7ovOy9exUWFoX
wh0qYtNOn5fuhHC8dLLUa10HsYb2BbfuuHzwexf+5sy32xG7lUdU2DVTsbQ66uBr
1OElzJvMZ3X5yPMt5heVfKoW6IFb7+VaIbcvERLUDg+PJzs2OUfsQ9A9eo08bwil
ZLYYb83tq+2KKyCaY0c+bhyn1Ok8UH2dfYRQoYiIsVQXs1l5XDZ9xvBzTX/7SsKE
yKyd4IBfbjB/Gy/wQvPQOmIbMAeNnWCKUvQN+BvnywbKMS1Y2W6rjfmkS8OCbiXQ
DBbWHsM7minxLt5icTBxvLxuNfK4i5vCCXFFlz1YFlPpXNppkx3TG0AjGmejEDJ4
M/Amc6zKXWokaKdDn8pVGg==
`protect END_PROTECTED
