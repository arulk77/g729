`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SfiKHKe+dYjSwh9b9sEujV040YwF6+kuiNOYFuYppeya
UxTowb4Bm94YOcnTwohzQ9PT+4nDu4E40GN+64aMONZsc9ntVxid1Nv85MfiA2sF
AuRwJkyVN3rziLx24Ej46/uMRtLl54EIQIS1t8uQ5IjRv7AV0YF64kBFuxdkwmko
Ej2aGw54ZOGG5Zof9OoUI7WA6AKgVLnnuCh2210r/r/VDIKMk9G/W4HBUASfMyyQ
`protect END_PROTECTED
