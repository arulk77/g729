`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEjtsy6VThjxHh7s98WYElze7IwnZc8NkHVIfttCofwS
P2NDJgDGoGIV33kGPhOL4BbCX40BTZiGrjFGpMsIz77e0Mx48CQjjR71xDSMw8pp
3wfca1fpEFNuFI4hrXIFhHOKDP6ACA9dQMtLW/IqGBLVhf7hgXqOR9wcfYqxrKOi
bdXH8ZQ8YMJfeS1JVnxJ+jon98+mX15p81cu1GQE7BXbbWgU64TfC4oF7qRdfvH8
0Slp8gvt59pod2rPE4coovfkSDhyn59YnFBOeHFHxOKXFGFLvRFxoe6pBr/Xpqqf
+mIs52z6gdRRlMh7rAWbK+g6bb/YfncHUEIZ8VXUkrIGQiK9DC0d9aHo4BBwwThp
Fb1YWn0BhU9EsgRch63ALIpdEj6XYPwEB2KT/7ndKhwr7AUoRtlkf6Wx41gWd7I2
x0TOHp1XvFAOiZLlMJbw2Hj3/dJXLzcYvMh9lsd9lPNJ7BO9vTig3F1va4kNNDiV
mB/DLsdZZ81lWENsKX1mRyAeie+xMxXSQBx/qLCYZlUocYX+xohY2MtE91GqRt38
TASVlYEdOq5MGglRRhLedCYB8bYFdpCRY1Af7nZsVU4=
`protect END_PROTECTED
