`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDCQD6EYdrPEXg88XEjJ/Ko0bmsI/mw6eC64dAn0LwoL
WvVGsu+kTHUtIMQJDaiOZaG8p+9AmmAXWSy5uHxLQ+xDFbmT1PjZ8+jP6B7tswKC
gtt89nTuMSwg0qMruUB6WO2qKMuHldG3BWDNfysjt9qv3qXkijfDbGI5N5pQWQ5Z
pODJ7nGJ5SwT7FEAEC3WXBXzGfTKMwDytVMroATA1ga6SyT75MZ92T9FOJjqvP56
`protect END_PROTECTED
