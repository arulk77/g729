`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu423hYURvF3hfCU4F1gvTJwTmYo/kOGuTDrI0X7Td88Bj
OEiVPPKDFP4505jCwXP9oOpTzrMTAP1tL2ivLpxVVWnO1Krq6lLB+eVRttlK1oQf
i4JwKwyscvyNPDg5r48E1O5QokyZqk+aXNQF0Tic/MeETB4v3fSvFzoya/7fFUO3
AIfL86t0/yEKd9im/63BEhaX/lvo2Gv/kgc3nCNkR/k=
`protect END_PROTECTED
