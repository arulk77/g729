`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJLySdhSUjfzz2hHfkZvHkpDtS+BY4iGfTGfNiN2AxRZ
RYUsSTKMS90kAIgX1TjiMlk8LZHb+VE1bey9CA5t2F+twomHSJmZ33jrPWwwJmUq
hoZyqlcGeJQt3eh9h+0UEzG8HfXx6fr2r/JixJ8zPeECiYYx/rC9Hryzk8FaTBAJ
cabB9LF97x8wNOxrGDwOZiNEkvlrD5ix99f3+dok1S+0PnS1YNbmDA1+zxU4YSEz
A+LdN8UkiI02tQL7+Bqkw7/a1MOS1HCecOlCknjbNFAUD1fR9M+ZwiT5aXEFUrA9
JwEp+/yqwqhjLvCZC77y0dSah4QaISk9jMURjkOXb2hPmZub5VGu03JcEPYIn2GA
lxNAf2cc2RDssgh72XvIbL3/8Dxr9dNVVoOwy/jJ6M+JaUBseHPgVIAgBuPNhzd0
ftRmBTpoE9+UwH+ilDwYE2SA7mXK/F/61mFBL8oZUn4g897Geez5XIBzOowo1ZuF
wSOjx1vJmc8g3vx9vnxt78qZ2pa4HLSpk6hKsEbcr41HQRBHI1l8UdOARnQqs5xq
G0r912XPAyn5KBy20ge4/A==
`protect END_PROTECTED
