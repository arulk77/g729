`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4ykVTguZrWGBFL/iYsgTRrVp/H5J3fmluCXRIZoCXkwx
HWilUShl/iZXGZ35p4MCpQ/v4usDuo7Fqm5VdPbtJtP6VB0iEpwjXVnqSwGNZqFL
GXbuclwhQxU39ZUI2dnMcBnEmSquDKaxg/I1Q0c0sR9TWYFM5uk0+27d1j6EObsO
IMETof2CUQla6p4qHG/3LloQaGIInye3E9a3N/opoMvjcxFAEPCeJqnmESYrUTwc
uSAToTe2y8gFBuN5mbWta+LfltVqS9I8IsHgYY1xfYRO5VW6AEwnccR8znW9JEB4
6bdEo1BVjdgf68+tcYNTc5XRsA+JzgXOZvLcNcCaIZkRj+RkOXgiIjoXEWIOmTt7
bcuNixQJ74PIS71XiaKrShetUehbMfUxh5vHnLcCwQyyReg/aAX+OsY5KjsZZ2f3
AeNRWQg7KNpPry3NAt6lf1rkAXGU0VjnpRqn3s2Tqm/wdtsfnNiBedUdVhfxxEup
kFQW91smSwlLLN3+rL7MDl/pr7TzXmURYahasMK8THJzpjgHxXFzI0CLBOKHMTCi
8k4w6RQF5tvscHelJI8wV0ts6+Lz7aQmiSBvStUHpq6Mv+7ivkBYMwe9YjNEf5I4
CMgmW+Z2MpolHvWpPPPVVfosdB6mc4GeMojPlauUX5XXDeXTiLCts8euCMCopKQk
+kvUsFRfJrev59k5a3Rz+YbxLeGmzT0APdB1R6KCIpQd890LUgfzMdgUVCjx/tuC
ese9S9s9YWuzSclvpeWookPlM/2Y9qEYaoio9bgET31osSWuPeH/TS48vcGfjctc
X/8/ch0/X1Ssz2ZO7eDfEa4wTnhvfvRKKrLOO1ag+329oJVjDGXljFLnrPKxmu09
6HlmTxIKQCXtk6oVSeSVdkFQMqEqv12xVkzyZa9xHOstMj+IwCD8NSJxrRud5WpA
ktFeceYanwToTfpGkjEV8wGsXu4ljTh96RlnPeCf2BX1QxMCY5QWEX+a+M2mJbp+
hWT2NMv9dMXIkItbMMtddC3G4xeM9XCuNeRTGOu7IbjIRRotMHbjEdVbawoWNfcx
cP84hOnTovT9eop3TF6m9XZvDG55fRcLuYsMkL4OcwttjCCh8/xnt0K6cNSsxpDq
wL0T4LZkXvxl36HILYMBn7PdxfG/CsLIcoVOO+dl6qF1rUxcQUMzGm5tdNw4p3cw
xgY33rDQoZrRFY5ATn64qNvxWqES7X1BRLbQFZd9bLBKnJNkSZf+6rO0g4y5+Wzq
6Ob8v0g99MPVox4bLmHng0gvwz7cUwSDZr27y87PGDhZw0gM9Qpr8NuyUxtZKDn0
4kNrZjDF7UVUGJ4xrzck8iCCCpQvvAoYUsc79aGHzqSI+GGo2HAz7QxkQQQevbd1
M8aqmOAWY/EZUzmaIKJ/giGiBSPwkjj9HipGCOGtk1P5eIgZBu1PkFdth6aYLuNm
2HmbhVIkFx2hLe3MWS2s3CF7DyXP/vT5oALLVzaKCSvBXWDqUUXoXbMZiWOsJkCM
n7OSo+rCWiAMwExM8XADXFuNga1SwHpOc+YFbLVRXKyiyF6R8oxeizJGEgT/tF4b
2LCltHHquShv0H5EWtOxVfFnrxpwB95EBev2qurwsZjVZcQU1kGeeBTK+0UuU584
HBJ+w/HEPchMfXplxpW9iXSDT42a+s0NvO4/E+JH1x15ofMH0sUG+UsxnUn7By69
sfn2MkCpUsn3qpWPt4QVIxxfVXRij1SOPAM31dQRcWC7Z66oPsU0EHIC9+/J9Di2
tnHWbU4bOH43YQOc0CsTtUaANNLndo6Yy1DkYVso0suz2OMzZtbKUcCw6PnAsSRE
U6OlsRUAF/LFX4Qh4SNm+nk8Fms1Trondn2e1p3Nh+qJh0h3UjTmAfECXcE+Atd+
HotMRLuGij6Id3LPIZu9mY3SBYhFN8m1KVmUffVM5vQKvA5fEUju0bMZmHJWWD8n
BRzfUQ7kJvcIGPDgyqdKvyo3EmC5rw6G6JheFQboJ69hdskdozY3iQA1Y9Yvf3fi
3af3SeYQOSoDKPSXevNRI4kPMOPMg/4ULhz9CylrW+42Xk6Kj1k9zz+gzDl7y9Cb
joq9KfOUuGE7YtFFBakeD2iART9vdFRrDBueFbANdqQ29FiS5HPgwxc1P4stwW4o
2va9u0UPzPZuPVQ+xmSB37Wi2UoLRNULBRCS/q8NruyHi+5lZ6fSDxo7AsyygClY
zTk7Vx2LfHU2rf+R4Josn9u2Oy5aAAkYmlr2patro7EbWsZ/rvihXPLhZB4kepjG
nCLNa2LfjAtFggCj1GcvmNmNbqF6TE5U7dnhg3wPhNuBja4fzC/UctuOzG8kUV0D
ZElDLxqTInr4FifuQ6NTOVQ+k1ngDI57NE9UzmUK5wdB8fDH2SQKbwhSihYXzfTy
ZcFkGBeTReM1PL7rJS09eu/xdjV0hVuJL1NnYaSu8SkTBd08YwwuaULP8xPIkNgr
G3c1LbRwWXu4wbHZGLGE/3gDFB1oiFl1ub0YiEILzGifMxf5h576h9exyglPQ6ss
6UZ4JZwOUCinAMEavDBCBBoz3+STu5xYQg+Fo+4awq65am6VbDG8cLuHKLz0EgiN
p/DEve9M3ny3W02ofqGFMMnckiyuBRv6DJpFRxLqGagglhlEeC9pDEEOpIH4dYI0
bbABgn7Eq5fe6NQZYuxOVq807Lau66bIVjUpIOVCt5BA9GG2KTxsvnJygOVcjvpn
KsDvSW3nkWUuLzVF/Updu7n7Io7tpj64+svyqhA9A58Oy8oXVKYnDIWEhGBeRjeC
O4LJLwg7iefH5NvzBY8Rhz+3zFwW660T/4c0JYc+6tOnIOW0BZTLBYkOPNS1B8IV
GkCKLg5ZeCVXyxyr+As1h9dzBC6XycRXtgRJrhSGqWgVxenK2XlF9MVfvZZhSULE
F5EugXv0ljEswTQc+ukhJgq/Vbco3YzAGGvjKxS13etvd/s2xgdunEQzJJBOoq1r
heqP8NZXgqp7MFKsJ/SbkjYUVzQCjcFFPfpenviO+qDo/L8PxV+ObEPwA0WnkpPs
rbn61WasJfV6jAkifltfWvNC6LKvfkCHG9G3PLH5K/kDiDstGoYHq4Bzcea9ws9J
iShyZ0DTDHSbNUM99J+Pp96NKLH1HohQzPDSw2zSmVrnU+zmcWXJDqSB2CeKfKBP
p4F6Ua+AhE4ST24eQtUNEq4mcySkuBR/OZrosKmfn2GDB5xSbqr6RHNsRG68H9cn
h+ymbRsV2VdLHBA+f+n3R0JJjsp/xkJhSpJSRQ0oljQ5yRvStcRD2AL4HjHvm7/a
IzGjVoFm3g6bxdZFDdl1vRREwHCwTLlGCzVT/gJATS3yEl481tnSpEur2ERgULnm
L3vegbyST90cxLhJcoCFhEaYZXBqW7VffA/moZMag9DLFnHORXm6zTrT5dl181QJ
Cl1RZQBFkGGlKy6bvZ4luCbN90Q3eZLupq+CgrAvAYG+aH4pe5arX5oWXgGJGkFf
qc6CGRGFdYBn5SHBPwE6nSSJNUky5mKt6unS4yiiYCoTXZQYDmILJEjIjSjLcRES
MgQQWLUd+LaAuKDGDWPt0i9ilnjwMISf+aeL5qIg4Y3fhOjFPfqozCtBtg/9HQo/
VR5Xw4pwJY+dnrv3Cl6PuLXeT811WN73Bf2Fa5vJ+LmSBYaU6DtCwVaDlwCZ8AHc
876sCMQ4SfTRg/tXLgzYh6imZVVAyfUT8WHDzpo/4jJX1TVCxMblvIfamrc12CQa
Agc0bgbv0eJX+B6kbN/SFJKX1pqM2Kvzcf8PZkq1Z3aR7pAcqlQUU+2ItLzbc+EG
xfLQy85PIPlyfCOo5VGvnF/XvpONDWNWS/IAeyWFILUj+iFUNE6DewMW0qxhiE9c
fffx35S6ZzdNu+oFffG8h8sA5R1wz+roYzp0qOz6j+zprDwCmPb484N85gGX4545
VY/MWGF47OAPmOVSjk3rQWOdh9O3MdEzaZtclXMZQ2peN8mYn2Nr1+2WdqyBChkJ
PzF0Xhl+uICeS7Ru2QZKW6U6krNR5fiCNGWuM5boprl1in2HDDryNHDOPO1/Kn2M
FCcd3jVHM2fLLvnZJJRf4JzdI+bjXc3KcibYTAJjMGzuywqVs9UJO3ZSaiJtkZGR
5dU1+HNg+hyAElqzPvmv2N7JcMWXnen8hYAIxjMf6vbNLpZ3bgTIP9I0t7cbn3Cy
YnFof/tQMkvHrIKHHq1krx+MacLKeaNIgP8mLE7SQiHtE8TAlgor5derloYgziQ/
yc+Wz4gE/Y/1+PvG8NZ2ZloU8LlHkos+SHWxXY3+dbltZ9hs07tJ2w+W5/wWLNg5
uoWA7BlaooYPl3Cu7wdECGu8NoeYxtb1VbcvSTznfarJacNQ11y3SLC/3bnQcwVz
NDnOeXdKKTpCaut4X2ow2S6K3ZgCjliLfvqjlw2vdrptswjmrRkFv0onleSqwqCC
lz7C88zwXTbW0M44hXkJV0QxB1CDfcUA0mFoq50bNVkyzqRLLm6Z7OK3E9+XvyV0
O950TS9uCVFSFbnjcf1wDYpcGpR9MX1/sztMqba7clsGYxAxG5vxTh034Ke3aZy/
lLCYUg9M4YLa7y+axbU8Na98Dk78rC7XV3zlVzFqOn+YWabEaFy+3upQwOkYxTGz
F/TqgBDarYwNr22wv1fx7bRwrNaGQYTwMRqgIogKJ8OsNtr5lmqP45W2p4zyXzP/
RGnSMBm9wUJuQcf1qgrNpSyLM0j5xlhV9+JFBdmevfjkRWzemzBfUrV+wQbtgYaG
JNA5RVsGd8aL2pyxFs3RhJjKpezuKYUqFK4h7gvdmihNZxlQubnTf2d1g81aiJOU
6f7JhL04XsJDquDQwOCDUISmj+cWyano7oQS1+UvVHuZcrRO9Fp5PGNk1yUNdooV
iXu3KCIV5pPpEg8OWfXEtUl1ZXmdWJF8FPap/anC+fRLVlARbYIw1WHzsgOI2Yww
sQTk0KnkAVMiCm/ECBLWrA1p72zTQOMwJlQp/wJLLCreERMhHEpa2fW3uJc34gmu
qlIB2dcIH60fpcl/HqLbcm3tU/kzm0IvqEnwT8yzmRXHaQ/05wi1Vzgqf8/BFuyD
0tPDprnpeVHEMBur1aOP5ETx5WoxB9PVbviSOIHtf9hCR0sLGCWhDwLQasxTBLye
qObgIB91imLGQckC2gy49nqrxG/vpvP6m+P4VgDZRyVpJTGge7DQTk+Id4n1iu+e
J+lXFIX5Sr/HPZJSuJEKt7OwhIW12LBoOBlbhqDGj5O1sHtVHC7uIeylLUZC2eyi
INBWnPEdjCZFffurhDi9pwZl9RkKnZcs8LL4StOszwx6igK+VtapLMAYvzSX86v+
SwIptL6TrsCmODFg+A9bnnPKEbnLoQJ9wYdmkH8OfL053O5089fRqrBUTTBdAsZd
ubRCo+S5MEXMneQOMAFSWynVO737d05stEFgCBALgVEoUSXG6PPLKeooAFtNKuTc
YeKllakeatYEVZjz1m6Ma+mJnRsxhdwOSPvSKdx7L7sdKqL6Kj8qZjlPNIPrZQ+x
omkZCfSupDCMNioKlBFWJUq/TsFDyVNe2++U0YgfDxpV8zJAS+PZM7U+tUZoy3Mu
ai3G+8/y3dw4x7sxXZghhprAqLp689RN0VWelkaVMlC5/J7FKBxRfboJLORbeRli
ZoVuzA1xLquWMSDvDxguzolnQNCKtDZNnsef2GZtyxlER6P9pcLAyD1aMmMuBr54
j0bBwQe6qN3/XGG7Uz2xBw2FwIGxsvd26a00rzDGWRJU//jxWegde12EzpTOQKnK
45M1m51rx5VzYnWGtYCy1Wrxn1gNwlteRe6Dd4Bebyow7eIh7eYJWDU4K/Ii0nea
2z0mh1zLDzY6P/nh3PT2y/281KDoZDdMKE7WVB3SLB/ffUnDLApO69j2hCbCGxKB
GUEj17Bzptjv6TEFBnsOFj6moIfYdt8e9y32zR04Fi41m47HxmTTOV0yLHSDZMao
8MORJemLTL4du7P29gtemtz2zxQBFgKIr/ZwLpBX29rnR3G5kTAVqB1EV74gvPLq
3+YfKBfXAtDHj5WIxuK0rYCiZoLPIz5Os6qjtg4tLQRY+uRF+q0UD7/Kv+0EMnNW
FGhW3DYNkrD3hMyZN9jPU8hYtVs9ZXRrNIZTjcLhySErmPJmdcoNmJ2ogykq8QlT
ebFyQlsgRhDPW1CcXchKUAm6qhAR1XVz0f33r7kPHHBpcqzdGNQKhj/yj3HlQ4CU
vWGzrUkYvVH1KZ28W3Ro6uvMmDxqhBMcTg9Jb4fqcZJhIAdkr9eIVRxr4RqCfbuM
Rc89FWbx2BWoA6Yz5GoPJr90sz7LCwtKovSnW++lYg0WVCbDW0o6av83czRxrQx3
ErjDV+stxkYS/84Ironw56ezfX4bAjXHdhGFLsHd49jzZOt7s3BSoxihRen/kbdB
ET0FfRLoHaicbdTkUljk9RBjxje665ZcCbbntLOGOgRnFWqFaNsUtXD40yeWFCkX
qX1PAEsPn4QLG8/fRVRq+TArz7H+OxMaHVT4Qs5hW+OleAaC964HaQrzjP41KVVD
MotB3yVigZ5kIFzwWdNBwx6qvSGovkoxbi209QM4hnp1S/xKIB+GmXIp394cFOsw
nEyI3UIN04JMRsBDxl3vJQafsT3lXWjLFR9v9y0K2WhPu4ZuF6V9kcUTAqrOWcjo
A/vuK2bul4xdFFpLvR1hOCDzMs+f2G2SvwsX7AgYwIFWhM58/o/a3RVDYR3BAYDC
gbHdn9rp0tt+VaRLfIvGvpgYyAYRyIvedn3DcZvOStl7VrWTerEkXJljgA6V75qx
dQbWtIXasqGVwGD966ssM4ndgBYl/gbbUEADKPWXoIYsbYUivyUfHLpWbiBrTAAR
ZCfdp5FppXiJybYeX+Ys6lLeRIpTGqnzNwBNfCAf8ncfbgO/o/dKPiZO9HzmYtt3
HHfo/r8SUVSZI4rHSJnqpPCpG/ceXT38Y1c8FxMC5Cf0kv5cefBLCGue/ZLt33g8
HgKJnJJQcdIzG82Ha2Ib1gI2bRumW9uc4EDWqq22cqItq/X2mnxJlfOEa4kYBkRH
502TNcx+VG/I0NoAxeNpzlXBpjtftulosr9l/iG3az7MbkrC7VPwpuJeRG9z8Bx7
egIidRs/5PrmYprh3Gu0v6gQmk19Kbvz8FI6AIQjILdDTcvxQ+IzW8c1Vz1y9ahK
HoTgF18ugp4hHkMgsOwSwmOOVT1fqPV1HyMq+YmieGP3S/ceA8mxgpPO8F8ygDtk
NxpoMTYU7SfjRoCHwTvrbmNSDBDJC0pvYJEZf8sZpdhtNXRv6K1HXGowkVM/cfTX
p7Uenr2IVGZgNhBcR6o7r/JvYmoYkoJgu8iCeQ4lZmzN0wf8Z8a1k3dmjToPvgdB
Xrnth6PQJKu59z6dQYS8WvwhmLk2Tnm5KTCey77yQiBFNMKDYpT4v/33o2/CZ0Wc
5Ax2+CALC9mLyILp5Qd1l7gLL7tinKP/cDvDP6vW609lIMRwewYXG1/bGC5JvMpN
IcLLwQce/dTm9biyudHinslJ2cOzoqzu26ZHuGOY0GlEz1EEf9aCbTEc32ri4XNA
JWQ1P75ohnq6pHcD3ra3eKR2EDOAlYLoU+NDEoIiZSb6zeOysZEjPCSmZ+Y9fd8R
zoi8SMkvYgBZG4VR4va77QfAkcKABj0tyqmiWiwXpjcA1n7TDTj0sfitnuroUean
Ae8nJqmeb/UYpP1B1xp8HaLi0r7lIJj3rqXIKuQI9hTMRl4+HETQiEF1sTRaWT1v
9tfKUdGjy3yP0HKu1W/dzHYyKzkt+ePwtv/UzUndAcQMTilqAQrTQgea2LwcanEA
f5UFcAr2sotz3TuYrMnnI0ij8lZxrpnsuiNHO8v+CVOqq4ZEwQHyYhh2Q14cT+tg
Vwax5AfPhYGhQLi2ZLglFbtDwqqfmqaCeMIj3pfunFlpsAjt5xfQ8jG8hAZMrVUV
eMcwlj6FdnL97/PsM4m50/E508p+WhKJrbUksgJzhQy+loTglUtL7ulDTXby75Xy
Wd2SQHNyLps9PaTH3PRchAqezLS2hwSB0onwwAGVUQvzCTl6VO1atWje3GnuW8H3
didz/cg9Esof5Bis60GYfSRha9BcyIieBb4FQsazgOnsbGNNTtXSn9X+zTnOvNx4
Lly9qvOAKcXIK3pw246Hit6LnS9qAEz58FQbuRX5JG3cZYD1EuQg36CfP51XTybX
64tpmkr0G5OomsFxLA0rguHoaaViQnWLMMynPMxF6w4eIDc9rCCZ2Vtj6+TQLW3H
oj9+W00dSqWZLrikYAVh8cAezcpm/K52qczlTUaL3X2aEM4o+8BNqazPAc9pof1o
8VpdzoJ/IHmb430FrxWv6r+keOOklQvMcLy+vBmUZpfsjcFybWBefaDOPVCbReoE
4JzNd+lOR/Y485PwRGb3lS5kMD+LCFFxQM7ikodZ3TmA8woQmuRD+/acpqmBoe+a
fIpMTzFGMalRuuBvFgT9+b/zsQMAvgyTUrqp7ogRhy2+x4xoCyKaBa/6A6QU/0ss
MLgbmTM8Sa3lGKDkO2SmOq7DeDN/arQv39Y8KgutMjxaajo+6jGXjt/TMuAqOJpD
TbkR/Ei3m8mgu8gN2qnwwU9NuVBH3SQgaC/84EHBlCfFPUQnI/+/sJzTvXhnn2pp
Gsr/Mh7O9uKoda7biWnYct87bJlBDvpmYaeR+aY8/r1BQWh8DP1P0lxZjvvagB4P
dktTQwStS00qzvyprXUq3UrSccKxDYu275fpFzKZe+mpCQQJoWm1dn1dBF0z8OZ9
o95T0xPTqOrwnZpbk+T5pNKuEVdTJR4esUWqp3E54uMO7a8Veq+QSGS2Qab6dy1a
XRXemcfcowHBUrti0OujlQOzW2rKjl1INDnBFbO2kD7lkgJ8Iez3btJyfSRrdmx8
srT/KPEWpLCOZEmRYlm2d0tm76d57Yi3RdQ7WJzARnAyydPKpVZ6jeB0nWUjG2y1
KbKWuzD65jzc0yfZrJmhn7PfxysRdXm4t5bEIHxqvdp5iIMk464NgCgmjBK/3xsU
RhGLrk8TqE/AYIjcv7LEMDrort2XjxylR0M73SWXrKmewnJ/Hz6XLJxgzP7eXHBQ
Ij7bMCV4mUM6WsV1/uLmgJVRblPxBfpkNU1nGhIf0Ae/4Txhpdc3Yujp1snvo+8C
XBQ0vVx1e82tkRm+8y15m6WTzAwZQLqAohSUbZaGfyEa/TOueOk3mC2jbelr8/SK
UlrXYIqUcG6Azkz2etO5IR7TOmjF6CwwUAEzBHXdRuQArKE6Dg2AFdGdywIKnevQ
YjFntlSxdjFjK9UYkaL/fPwhRaofCW2ZMlIzM2/j1ZUY9Km+QDuSJBmPxB9qpEWw
+izA1rAQDBU4pxHWq+XVxn7ZJhg3w8SE3wBOmdX//7lgq00BZyoh7mLbmNFSUZiy
m0mo91/pJK4Vva0iJENst2DeoA8rhjCHySv+wcu4HgDswYpmGowMBn/jtjvG5m2X
klh0iEcplkyLWz5syC+itIy8jM44MdgwTVHpGIhjnXAaTojxnTQh1h3M2Q20CoVL
a02vyaX3MUYL/upwaxj+qv9tdNzTr4LeQ5NYwlrzIqE5Ui8E4HqKHIkxuleoc/hH
ZO6/pNALkBAylBBYuIwWhd+XsD4o1tpoXfD7P0PFBaU1/4REO3EOkwQiZeQHsK8e
zwcpNqWqBIHfKOs8Shblfs3fgmitihFpEczj/YfajoD7Kx5rB0iqaNTfStQ3I4gR
ODvpevGWCk/2R6SdTlFsjJpP1Tg7zuY+vwcqB0fktpEjEX4rftJ1xJDHC+dYBOcB
q2lGENGOzIeZ4xmlYf7RZ7M/ZrPZkuDdHoaTrpy3xNKh2in/3cV2+LpuNClDOyir
9gjxotx6hJX8xrXtwdiM3pDDO5wQYhgGJwKKSLvIlpVwNf8aBXKgu5uYabualz6s
Oc0QCXy+Y6w1mgYAJGLm72Tev7R0L3ILo2f/piA04oZeF813FOnml9d6PBxAM4GJ
+EzwpOjLQwbYnkF8wgxyE7m+QZfSJGyjaFcRrBxuiDtRqIkcR5sIfOpMczrF46l6
mVsMma1NPdEZmvu29Nd20oaZ9ZXDhvDrlyvt+RSIkGp2DUy/7KqmwKyn6dH9PHf0
jEzYD1Hq/5x4FMqOa3CYd6AZmDVBdVVq/YX/Dz9XBAV27vlH1RWMekfjRjT1064e
OhlpF/Mgk+hamgX754bI5WKdSZqm62W+9Dyz1DRe7lzTBL571WKh+TPA7ltYFTT5
NvRBLiwMI2jlkCFoZE7EB/fzFWdMmKKPtYrO3klN5C8HazlC7CqCEW8ZrjHrUcDM
VIij3D/BW4EVQGZg9svqouMQBRFvooj86x5u54XZP7payBctlaBk5LnkwzTe2b0Q
2QkOZ76WNQAptZV6FnnoSuk0doxTwwACeQSmMZTqFpyHyuc/tqmEzj0UOaxLbReK
htultJunHOJmmd1D83touHUiPmuNSVzTZaeRVYXHmuq43XcN2brdNFooV9mL+sEO
wmAbsaKadXY/otO2LR8RD2VmIt89cVJ/RtEV4B20l2BJRA2G8/GVR3bAIXKJIIZS
aEvFG0G93HHGXb8MrDlC7yHlMo9Zn2cr8bXMqGT70DTUJmHRtLDrEY8Js/E2plJI
PrsW/SAsDaFttcTUYJA5YnQv0yyEkfzS3/+SHhfTntLt4ELQBs8OgEAniI4wNeQR
wLiTeXu7/7ugzFQByYHXG9CIexm6EtvjeoD59jb6rs5HThhAeP4dsjCK3h5PyqCo
d3YWeWwoDibx+/zGazYVuKABl4nZAuOWoIXlPCONqZ2BqzqJ0A2SZR6jxJpAwamg
HWE/qeQuAEMhGEY2wbx+Z1xp18jXrTWEJUrwOSuf8mBll0JwT6hXrkr+X4Qtsn27
cwJft/WIYHJTMsjSeBZ74HMfi1CU+8JMNN4PDaezWVVebOxiois6EPJgNRSjoAl8
8CQ01dUDGgwbZbnisfe40KihlVUgU8sn8UgGlx4C9h0Pb9L0bQZOByNhbwOACbT4
97TqR/lVxOGx3QZkba6VHSJXenpCT6WYkDFM+BjdZH5EUowPdcqWCbpwBSihmVVa
kXBOBfKr5kiKZY4TIPLm6EdABmnidHsLU/Txue5B4feF4gMjr9LltkyVrH1Doxkf
m2JuV1/rkXi+t/k/Nj3oaTkyPV9kjjQnjUu+0s/oFG3L98JEf6uw6QS/FUpq6gqR
fE3+0RqyItSc2zeSeyXoljNYTpPIHQ/TkjYNapXqF+Qpz0x6bnJG3kskrb11jpzN
kQDQkkfDPEbh5m87BgiHp1xg2AiygHWaDM54ak7DfzmD9PQaJjBcNNvvAwAT9EPp
Yp2F30hoFaXQln2dJHKdBOBH96QSnDE2MUc7VT4PIYjprtLGpGwe95mtXLDdBMgs
4iBTa84y1KI22LAdP/yOnGt5se6KULl8qTO/2hIiF/bGk1p6TdRhUtnXrToqTyeb
JTcWlt4bxLB3x1YZcCSFAXuwWav40zWkJmkk01A7ruWeoEswNuxOac04opNj+nx+
Wnh/OyJfht/tDmQcAA6nIJddKRB3a3XuOcYykkaoKIWYQdRDaIn6zQrMYpDUC49y
/TcL/LG/4d5wbtksVeouJNLfJdKmxaVZ1gBfplDTsXnbpqNBAeDw+SjyCrPvqhZn
nrl8mAKm9pH87t0AW5B8bgM3MplB3hWSDoUJo1wRhQPlzrPTdD/0HI396//+KVZ/
EM/5Vafq1cv355Dn3tCPH97pATT08dKdBOkw45LMAV5PoAk2070P1hsNnDu836Ua
VAZ4r1hHQ6CTTjG4niqj7uYAOThADYpVn4HkXRlouxyUXjhUlFe0HJBjcKfNrG5c
ZYCfhlwJmlYls6qQCKTt70WRghee6Th4E2CKr3EWE3mEdHWpEcpto2u7Rxa37N1z
bDbbHayzOvFsY0bVt3hRr87dgReOqa/cdh848uIcSzA16BJCV3xWVzKTQg4eX5BF
P4rjlY2aVOuuNyhxznU+oUJehT6S1/iNSY/bbX13Q7CJmDk48JMXiMBJTQZ5i4Qz
UMqYvu43wHIQsKFVnbj0sdpi3oGiadB5/40JIBJeViBUCJy2Q1qUT+1WDn7CqY0A
yN1CkInuL/DdR+M4/ZVWVB4BldhUYrni9pPmOUtt1Pk0tJv5kZHKX3a7byJc1gKO
hKAe+a8VQtqVEfFoHX9cRSRSnQrZ6PjHB0uK0MZMZBYMqeLSXYmd+eUPp4mWyabw
QRgHxHJ+ZWtrqDlkTSysYdU0WViK29MnRhzM4EcugxWQVQ9rzUeNBHlqlVMgCXtz
BQKQOGVL3CJzrhFFlB+NMmk1NVPH8Uo/HQIcTzZy62pPG/38kSeydkX2mCwGjclQ
UrPiz+6YdACirFJp1SDjdNMo87TifiARPkfzAd7K6DH4ALCojwPIzZyEsJO0Nj6F
OsIx62uUQHMd3UlhiVX28qPUWu4Wkejp1zbSZaicnczqm60yNmbkVKbM/+LBJ9Px
Jg0BDZMYxbELWt+PUy9i2CBt/d0VWFPCOE514Qm8aM/KwldDaw/Lb0MrRSAKKWa7
ZAye1miY3/SDOnsEXmMNmsKtnwSdkWZVXht1tOBZvBeP8o02b04FnGsxkDqUr/F8
C50smGj7byGfehrXljQwVLSHq1M4UfbkLBiD7xzdkpbYm0QELOM1flkHXoqXmR8Z
9cc2BOin25C9DzUiaCCt+5yY6muAPTRwi3fdkRn7l9FF3GEShw9u8pudplJIfDKj
bqYpJ8oySUa2IYUGWUxpQJaLgtsMZ2pv7K50UawdHvZLnsygvCbqDJY3fJvfwB25
nXePJgAwXzFaQdZXj3xVQmhRKAcy2p1EB7XLCFI4dEUyi99mbUtljMa+3h/nVqIK
MHDG0rEH91yNtgtp7O2zktaCdLgY7Wpb4KSXj3qPGivtt49YYbE+RXNrJ/GwLsaa
NXW7QukuROF+XU+RAZOovKfuRYcEfdFLSvINbW0yW0nqA9W/nLjX+/ssCeWHVvn2
VI25q9Y1qiXABwQ2J2RciS6WmP6FV9K66VcETVdzQ+dFatvpXIPt3zI5nYc7anF4
80iiwT5m9WNPNv+wRToAxI4Ppv3bAO70PR4yFZz4jeA02TVcAsB3yPy+TASgG5R3
bt/W2vW8Vos4xr3uN6UdI0vwE/N+YkjTh3qHKoX7B65jDFNYa9sR0tTOE4Uz8bpe
MoOFDqSnCJIEk+1I3RF7GnCvXRE6pDfbXvQ2wJqTjUQvpvoWl29TkAJVRSRwCsW+
l/9gUUkwcmpH2G7zxbC4Dto8UVxA1W2CqSGerBlvVHqZNl5SnPMVKV/y3YZbUhlr
OCQSV9+yusDOZrJ+Uadr6W+6j5+kZ+F77mF8QvMikGt2I2+DF+InFVPTbPyfFh3E
LVxWtiu5ZafWG1UQxMBLYieVDuQ+NRgRz4OEtJt2i6eM6oy7bxR2iJEAd4ygSzBl
2Ncyv4sRzICcNGbrqzh6McXWL36w1P4X3+pY9HomeoQUEEtNxhCi6ModpRLdv+3g
v6ClfiGObi+KjKSPCWTd/lyzEGd9/MQQtUFaHl3RizuX1oWLn27bRsrnhtHMfK2o
abax5bNZtrkOZc+ZV6JGVFehYeC8ADovGowY+c4jedcWSN8x5LMKepO7OzsmUo5r
/NRztwLXdDLR734a/EySZY7IheTPynpYuIemPmeFRFrbYs/rdtE+Vtm8M+QYsB3D
YBf2HDGo9/En5LHed77SIQfJ4oRwWmLPiXA42BmBh6DKbAsHjynwfSndAbcHHnrI
RFxnO09kN0QlXplQTBMGQzEp73QY8wUMQn5GBP08mRffFG5uEC2T/f4CDjby1oyX
6mPRp7FW7JG0RMugwUMVfxvuOXA92sY35YPKxvLFoM/ugrb+B7Xi6LeKFOH/AdGO
aB501QR22HtGKPlSAg9i4nlUvtHGpLUao4B3wxSQJL74MR3yLqd+oK8yy6Bq7o0N
tcF2i6lXRCCG1neKLzjCjc4oQ06PIy1cA1kyeURB6EcnpqY2xTC/zStXwvBOaW5p
LvPev3foZll3fmMJqB3T+yCJRA9kSJxCIS1F7ybgsEnwpRtE+DwgsnfapQr1K+Cg
fb7MJffkKyg6bP0wadS15fLj/MZUn/eQkjOmG2D+33zTGYNTig3uPavT1MLsmtv7
5Z0QzJKgBgiQDL8WZte1qlJyCnkMcIBjvlMxXK7GS04WUfJ33MR/2wpS7lGlDCKX
DY5tdKARvWmMTqjdUC7z931+XtRc+gcIE9Z1toYjthMj5wGGVHEfoWS5GRv7BhlQ
xRvhHljvn8+DesENDaYQ3LlT/WeQ7T4eCkCF+PpbkEx8GB6qBOowfhtPaibxlL/S
3C/9Wze6U4j599ca4hazDC5b2+uupxyuWj/u3mN57yZKP4dxluOyFBTYLc7vXnmZ
W8YZgpEe1V57QRFk491wLR+HDwSRXfQvu0aakToX0v1KEtEoWskG+lGA+ZNLJC7j
6kolkGGDvP1l4E3wVBE0nWFhvGbRBWtw59csBXpw32J44h06tsXFwJIPj5cn1e5p
Z5dWk18r9dftYQyO2irmUNoR55PJZWP2M9SJLuC7/wbdCgoYJEz0mHVHZ4Ga8E9m
YwCy/vZAWqZ4V2hRIEM/cIv1A61piSRMqcCDEfvzRjuWtid5aBW0FalcmnVWIZUe
YXt65pSuTkyS5VgEee1RuaUzI2FZF2E6rl5+gGpc27Xel1SfTvQPcx+JE8wKVKiZ
RazV0WOeP0OC8iKEoS9zrpWdkd9Q8B1/a7MIaDit6dyZgC8fTqs1Upoy9oTcRba0
tnL2ntvSWbUu4BpNRBiHzl+BxuU79fkIrTNNhuYE+gHOiQzRFbeUAASzLP+a5jKc
fejnFEZ/t9wB5/DUE+SK/kcz3/QLkGQI8na10o4a+o96vgP4KF/RAI4m9jjsrSE+
8V/V3mUKUn9kRNnwUZ487/Z4ZgxfdZUIz9WL7dEQ2q6Ict9TvkKyUqxowmIM9eKK
wVx8SR5/wsLhJBXAx7SdQ7oxh8zsCijZA0yen/hiQLmVAhtHMf+O+q5w1NlCh3YU
VvMyY5Xv2XcgODSWJVJXIHsl7sKdlB7u/P0lsu8GlN2Mz0MIC2jDik+rVR9Nfcct
gVzivOuq76bIAEFHuOI3mQQnZT/pQHvJpqK9O16QWXIrf8tPwg/N8hD7l1fhiySC
xNCGNwl0CDsXnsWx1+cygYoIfv5lWg1kD7uWMsSQ9W1DUQCIIZ0A4CFKtE1D8NEx
Dvlz6llbZhWz8ZBuitAgl+7Wkf2ByGsmn76F2/TqCwU7OuHOLwt7Y2vvT9Zm7We/
EgBh+waQrIpr8t9K6Rp7uG71aYUhvuBnC4iexxb/kwoqHQNvNHjy6TOgZshfNSgt
joMgjojzXKXGG5ZKafZ/tHFPn1w4dqHOoMg1DRc2P7zhx0n43UcyWdo2h2Ne50ji
9m+ZjQHOGiWEoTMWhhSwXE18OVm6DpTVsBQUKiS3BYg+ZvYfQdviZcuLQxW/Aiyg
pbNbb2tq3n5g1nhiF911c0sYJAWeO/khr2CqAsyEkLtFhJHdhRzUwmEWJu773yda
hzpS8Vj9gQqASLvPiy6umv2/Q3oRzIKbwXFWB7EXJnwDfnBLmhSdKH6h/F+ctfc2
3KNRKzSZAHECMTr34g1GznTJY6c4WeznNSjn+RipphzCU+e2OVM2zBEpwYJyaSqT
MajtsvMogk0z+3c/qXLuaKMwdlamiQG6GUfgA6YTsv/G7x0pdZ7FwXQpovze7d3C
IIse7aJDAuXtdkFpncNCYXs0g1mhdhIGdWI+rXPbuZaG9Cle+i3IwrSD7G2LUsBs
a3epGAgXHacTczEm1tH/IumZMp8NYgEkEu9xzWgqvv9/tBvT4YYrsRtzvSAGm0ok
hnfoUwy0KoQhwGonwk9HmHvjEBIQ4BzrS17A4oS5LzLEY9AjPJzbGQJI1h2rV91o
srRqwbPr+b79Sbyi08rjsQjdFRn9idZgDJ1dap1zw/dqJjR3rkAcyT9Cstf3tIta
tOD6qySTBrxhtSXpqUD3Vgij0c54LklreR0T5xeG4fqz7mrCt1mXU3Eb6o007THg
gycFSxeQVyCMBrcizhpMJ6J3nawONkKtFBqLrUitEtAaphRE4Zr8OKgrsbQkalqr
w9yVrsS0pOFNtkp4qdqlRrS8MaKY2uR536OoZUKZ45MbIqI3SZGSlJAG7n3BfAuM
xBKQ3YIIXI/cwmDxYjroXEtlL33bPWHi5hBK5air8D2s+DMlzcMJwif/HcKAf28z
eli9TIx65pNXzffQTPYt83CGAkLUiCMOVHbQZt4Qg+z5Cy27cghJLQAXXoU91oLS
qWbOyDRilQZZ89Vt87VKYP6nZJRVu3GQOFMKxFReY0gbFBfGts9WFtTcsVb2thOX
Ub4R/Rx/hPipkEeNpETX8GqG0lzeIoz+FM3qiLoFncwn3IetV8T93ynwlVDDTTMm
tiy0Si9zrPwMQ8yfVQY11hZh6na42XpYb6eJZ8vPrVGGhT2HoVt1nbWVGsKyNP1b
0Kxgl0gpx8KHSyKw65hFAagnhmC7Y1WyGi1Lh75TYyZsyWf25xzhYzo9lDAmFhrU
iEBuie3nf/Zaz6Ip0KOj4WIg/HuIlss4IKxUjWGXaNaDyBU88FT8KgTbOXovHC45
N10MMF/9N+Kz7hyCSEU9zEe8PT72hYuHIVnFyUwpr9NbPPpzAOHIbL6Nq9bufkfl
K1MU8BNLjBExZ5d+IIXusd53XN+hgRDEO990FZVMRwnJxtVK8SkURU2tj2EWNZSH
1lBJHd2g+iYE8+DTkIuCHUNAHd8Qols/LY8YwCUFu78wujIO3ELbIxPpmYhYEH4n
pay2Pp9woxuIbURjN0lW9QdlqRssKsC1sn0WiPnPg8TiycTTXq7SAMEYjBxTuIrp
0SS4HMTNPMWkyduO/Zp+KDM9XeXXv0yJrY4YbyyCAfvuMm1DYkXfGu913xhoHDuJ
nk3/8Xtx5x3mc1jjOOZJkbFFtM73itsljSZQ4g/K4cvWDbYlguBWmHpGy+ZKNZJd
+XlgWjAlaHkDm3N1WXpPXufJeq7ZeCTLFo1730vHkzxL8gKs/cEMRe5x5MWV0QVk
wqNh68vP0JAK5t8NKhtoZqwMw1RpvoihMXN8GNBuCd0JDvHL3RXNcXwB/A494W+R
sRti4047sw2zqmPQXottAjoMFDRKDz3pRC8r8z97XhWzdfLRzCVVBoOzEs/9uUrf
b56aUZrFGFARjewVCdVD3x3bb+EJdEcex0+EKgnA352PWjndPrCUjh1O/8DJXxxZ
csHsugQqNB2MG+MTdu/bCjL5f/eHeVllNyRgHsYGJgqYPuDc27tMaTC7etCJnzRr
wpdqorsCqezKEVwAiOJDrtk26GWkN1Nl4iR65c839LhNdUtJCw3sYpOBVqhamQYs
FdJwyJYFQ2clSzVVNOcawvu74bEZnQj3p4YdQ8AzNQGsYRNhfYIQ9cIUPv9HGqJz
ni2erH5vA8R5bJsdUrgMGD9RaN3aW8Uyw/p/YKE8uvwh7fc/uHi33kFDkGSier8P
4tNFmG8KgADeBuZuP+ztl0dOQY2RTHcRYed+F59ccuzpvi/pE7NgCuFRU36eiCPx
MXgKdZ4PmP24yOrjaBUHNyLlOmOdM15GjjH1paeJgJmDDaEh1L+VB4eFUs//mfWm
3K3TPCXZUi5Y+cyKwdyPf8IhcZ8Obio/7crtKOBKXJQKYca3EZwFV+8L7ZoxR+Cm
rjP/W2nQO7sc6qODHdMz2/sKlnfcrr+cj/Pxyn0E9HuGw525Y3WY0vm2a17c+tgb
4DMycUciJr+urlTzGY8kooFJkxYz9OPN50NWcvFu0Fgr1P5O28DmxH1NO91uFzyg
VmkEeVgpaKymNEqSwZ1ZKEp0EZ5YFDoTNjQW/USyMMM5vYAI07+ra1FkiHLlkuk8
wJVjHiQoHTdrzb6nSQCBjYGNGD/9QyNO+tSftzRa76vwO3ya+x07vkjVVU4xGoeJ
P+fB9J7LQHK9zzPyQj9T8II2tUYSXtn7UIk8xuiQJkSqBpsaKbLScObBei8XeNGh
yebNcN4rmbMezu+NK+G0bLvDJsYHAlIM//4ikzOZ8HBYqneFoF9//F0Z99okvtBo
wv6d7qf53Z6HWLw74pv+cpkaqEQBLGdy59UaMuCr5Bl5BJ53bUc2cyHJ0Mq4ljUz
4/+eCmTxIVnwjBbKL5G+EmW8hZ+sxXa/KAtcLcob1cpTXzaFkPLwpbNMNiupndCy
gKXk683ZlqQscYCyiys+xCtgfMQlEdgv3vMSRsFwheVImZhnftDckJG0U8q/HyO1
tvUsT2tgf8+hto6yTDMUu8D2z254AKcsCAXsLEXVwTD1AmY3wCw3CZNzlrBjp6vU
3GdICeOOUY/qSUb5+mrEtP+Qm4s2ejToogLU5tGnXBxQr67kTBoBTRkqrGRyJoZB
zs0PWgPjJvngM94e3NSuGr3ALqXlKfdZK0HS56J3yw7hjexWBx0fnWTJ2bRgrjh+
y9R7dpasQuMiYWBzEbiOxpneCr+acYENugiNIXztgdHFsxzKNouBYw/qEinPU5fY
nH5Uwc9dPdZRjoakmRklIro42g65azhsDmZMJIUMZbaK6npD+B4MDA6q4p6hggPr
Ri12xkN6UGJHS7CLfttOFclKAMi7N/GXUTKtNztkIv0J3ou8tv71NSTitM7TUtYr
icZcJvhlOYOSwTvbd4uwj3hOijAz6ak3e3ncKggT2khzuJStWhRo/H6eOyEhLrG0
Uq0jZG1GRLDbhp5tqJTwjFyuo7+Dr3VKeTuQ+lZx/Thdu4y/xtdaMpdKf0jrZs/Q
HbS2oBk4QM4IxL2ekuLsw0ZFbqZ4lXntgvZGxv0ia9XfnOtq/O6Lp0ROYkMFBNZj
MllFJmdG/utDleo6eYVjSn5vRn/D/g60xjWhM6x/tDBvfDqRQoiwDUFODHhG107Z
TR/mQ7yZ/zROyRRy8zi9/+httZnYpw1WZ60c184pTQ2mACyLKqm2YnReA5OUVolc
C4gGFlh7Hcy/6EtlL4hgj1SGn5o0AsmpaEsi5cuUK8nEhw/wNLkvA33aT8946v3z
AN5KlDqGTlBkD70EJhketHlR4dnS4lftmuuXxh+iaj+07yipUom6U/+l2AUu4nl1
0ZrU4fxHpdk9vXW2iaCoASUjkXf/h5l4zIflNPnfwams5vSzr5w139nMr0ukaEoD
jLPyXmDeUREgOLM4RqqIgwzsQ82rcW2QABbVXSw7qU101QeDuE713XnWjMMDUuxL
CEg+Qh+53LRbb2i7gIJB6w8h734vBfw9CiJgQQrIiElFNFNmXkSCBkwzBzHQJVuL
pv9VDWfoqDrWLHeVRtcsakwmcFj6veAVgtvfPmoDLEhNolSR/mV6BQ4smz99WknL
H34Bxv0rEfLFG/BowlMJIb9LVJlWOx3tQmm29jd2WFNB4o0rr3SPlMllMKgc0YvM
MkNB699OZWDiAidQT2s1pCrLl+e6HGSDTzOXWzpc9earGRgKHifKCrwCTHEi7ZxR
Tdl922sh/7lZg3oCBISPDzJV5uCHxz4WFPw3+qstjckP0MH/DeLn8esD6jKR2+Pl
PM52SFzwrj9O3I+qIQJmehwEwGtjUuZyPxm8Tegwid4vJd7ZYSkaZjmfRIO/7WIf
YBzf+4T4XNeHmE8AkALRcFF2zaCamNSSMb2QqWFvRnaEONyJHgUJO9SUzwcxWCB9
fYVb3zftnCoCeiTYXoSNXwDf8bgol+V59Gqp8J47IuDp6Ortq0GpgLLU8NrOWwUh
cRyfUj9jAE/IyrMu8nCfQQBoPl3MCLnKosr1aZusXltbHDB3jZ4FVVeEj3OQSG3j
jMy0PPul27ZawgnJK3rJ6PncFERy576Ni2YBb678PnzuXNf/8Bvv+UorYQc+p2af
UJY7QmX9xl/mamDzFkR6WsSUtIiZ5sg7ygRqgElbjq66LH7mOPDnvFVVAdaIxxl5
npwpzG2gmRsp9/JUX0ZE6T5C0aghQZrL8vWURWIdO0Q4zQMfr3skoSDxEDOdwfFq
MwdNDg3HWj6dF+eWSWXC/j8P6/OhVI2yFlEGBtOK2ictvAH8vsL3Xmd9Jtojt8Rl
k02ltW+KlxRgeTNbiOx9vTdT0JokMHcKSpjIv4eXLRWZ3ebAxAWP1c2+0jTH1aKw
buPz2A0MVISRzLgVjqIQFqVKL6Tq1vvBMfbbe7UGDRcSx+fB5BJ6ZnViFAyVn/pS
SEF24HSSfJXj+k+hsQ4eSXXhoxUYkDNAe4aKI8r3/32Bzk07+zPigOqzgRdw8844
5Cp+62e/ev8ZzS17dCGOFktQWmyykJqk5mqgsqlAZ4Y12ZwpSf8qPQUFISLN3Z82
xaMz+l/AwqAOAt0uQq95P5/AZDvjm3E902+ZA4ulun8z1QRJTZ+Z3/ixgHaLYVqu
j3wXXAWzfYgd853ZjfTTVg+SEwDIMKBRiJOKG9h14qy0ivPSpU5l1MIU1NflQ1FR
OMuSQWBeYFBG3//h62FbSpXVkraIf4IaZloNwPLA6cFnnrvqqP/9Q22a39q636rv
mNlUmwuLVQEGN1ng32UMjhlkEbSnq1Mf9RpRv/kDTFViBE0LAIq/kQ1B4ac3p95y
L7wlza5FaAFiLBRfH0FEoDVjFNKbVrJnPmawdDx36YyEaFaumVz8mdnSNqHhamp6
mxTN8bg06n+vzSkmKKnXcIJZYY3VAFMdN7J7qCYKk+fA3DKr2TIjdBsMprHmzrfn
7jUQnjfqwTCfxrTME+VPqTK7oD81wAHM76JsF2WTFkNdka6lJq4bvDy5gEL9ObVM
wT3z905kW7LferL6jv87Ljm1e5ePdDlbuCZK1xuqNV4qSPa7a02NIWcKBwqCuiHm
s3qKNHb7T+SnSeZgqWHyHtPw9Br5gjFIRlQwA5Ss5eDbxzq8TUsnLnY1XBYlhOAq
2niFPipSqFktvvlQ26SFDp59U9IOyWW5JoTneVRri5UABlffS7wIBDdTafeSNUQK
km+3dqp+PZch3uoHe4fxxls2HZ6mQsRRMcenAPWfTSesd90tu804qOFiyij95Qqc
Qdvw3i7oNSec2xkD3KnF4s2BsjhahIg0Yn3vdif53pzPUUB5rCgtuiHtO4yR1M9e
A/tT58IheQQ6RZv25lhpg5g55MHwkhAc8ynKz3LSfspqzGuRlxGqHp8UgbkIIdE8
DKMPmtdwFrgHPu8WUU2Az8HyGGKGI3R6Z1zSezQsd0HbIfp9P4VS0aRNGeZW1ozC
SZJwcsFSSDEImWdzALk3T8AMZAQOloq4IyV2HexO+gj1jYLhdsznoXcBXnYi2ImP
GuUn2DGjzw1Pg3I8TO5JswDoQf1xwwxzBqfZxDY4E7ahlgg/EGYPWenH/HwwD7Wj
0Inww0edf7yA8d0qzHKND08JY2+paiju/ebqd1l0Baz3JxnaIR3zhXBmGxoJ0Ff2
LVPs8ayvoVAj/c1oRoYumdkZfd2+1NleE7QD8aH6O6jffiS9xoIM8+WM74FYuVqG
jCG+4Zi/gxSfz+bRU86IPsUwsepRFjlA4I/MMG37XrjkCCrzwdE6A4ltS5OVWnyB
/foHvY00jwJhypqmtwYeg/gt62dbAOzcdS0pke2DBt473WvxzOPqlAqs1otR5mUD
zxbMrezMLEDWC0ccf/MfGYBU5ovjTj2h61G91kqkC0Sk3GQeKYVpxcPm/+GfpO36
daCFtznPhCvbEJO5McKl/irD+q47RCoVRhF1V1TMrP+bWrda1UFz29TI3jKfsbFS
2O8U/RJ3ro5jIQnxSdhwk6QeEDfewxMZejSQMArkkN6iEcZqw+jyTni5oOgwkWgU
yPYbvEn8N8bgRYGEXd/mq5GmJqjui+b6AwQ1bNQkimVbYN3rxMcvzwPrR4/00LqZ
z36A67fjX70ZvHV2aMgX+OjXBzI04+19aSCZsuQMnvK78fJC4TwlqwNWvvSiVoyE
BQ015c9c1dkj50pNMOAhdeE6ih9EiEZOxDVZwQoVRPy8JEXKEpyEd0+pf/rmigDu
YRUmb6B1QiB4Oy1t8H+n8hAW5rYZkx+4rAV3Dpaw5MNVY/tKo1sW0NZhUo6HwfFD
749owZkCmXTyv9s8SzpV9B0qBDqH/x0g7vbHhZwF97KK6EjfVgckBcexrpWNWo+5
lPNbiZmDTLsIIyLKnj4CR9U8UQcflvL6BrlY4wd6UGabjoHOuE4SefDEsQMYKsK2
SORDd4M6ckwOlA1/aAdj5lf+dmLQ40Zg8K/aNCU1cJEBWUEHZnuot4Q0+y13BfKh
rChUIDBs1cikQv4Vu4IdSTpbNNKz6cjIhhqkF595Xxd1NVNxai+nccEXnWuD37V8
faHX3vmAf9n20pCn8ZoZWe1iR+20uUO1Zg+q8izczcxiQnOmvzcJ9pbe+nFaE5f2
YmP3VA0if6WQN7G4OJccxP7MYcwQ6ldNx4bdKUQ0aeCImG0+oDFYeTKIc0TnuFjH
Chy+v//yQKtz0eBsedrGAYwOwF1McV/lZ7Au0PkGFLyLU4i3SJi6aqtuc3n4CgTv
e9SfsIIl69yeoDIJayCu1+zhEtUffaUUuMwheF4QVClAHrER3CLpyO7Q5c3aF04V
ibT7qqV4dcC7PkXnFt42E5gwTRUBslDWatXAeZ8zcOAyt5LTQzCvpaF7A7I2yv7I
LW9Sp8DGcgy60F0WXNZe1yY+qGyw6MUNMM9V2xOHEDlPC3tczTwCW1XsVpLk0Pjb
b59pInk0uhGNMcVoGVYGlHhkcCpgrcCfCTtrCkOu9NCooIWoHfIPRRDqxtiZMAZ5
CUGe2z0OQVYVdx3GSZYfIiVNJPYWJekLvenUjrDzt4RvA6XXxqxREmHdJqxoHkZs
ZAiAjABSMq47zvsXJqsw1kULzlzvvaOshGrBzUikVT5DKmM9v25JCJzbo9H3Y5a4
R0slGaGIHbx21tOsi9BXUHYsV+h7RfytNpfQ4ZekWWuiprYXT4hWsnwMnbXpbIae
Zr2a2Opm6UOOPzcL4oJR8oePL0h1749IUToce1Ah9lQ1kVE38YCTmQnIN3W5m0na
LKbKstWEg8DNU4L9I/XMKdglW6a+sIR5ZZTjg4Cvz0FkWJRMKbrOj8D4NtXUFoMO
2NpdzxiDQPf/0TA+d+2XKtLp+XMb120n1vwGKNIL+8s70pYshhbH1iuWdlKI+08F
XfzhV3Ku3BAS/5Tju9yWdxLvNAVuMPPw07q2+ZVcs6JKjkC0rGeKv/2sxKx9Lyi+
gjRywsIX0mZ3y0dD7EYcRL7mi/mwJV7GSbdu8ZdwLA1lhff/NogBACLjbuf4ucWn
pyCeyXxu9QG3vz9CdGqOWRY7P7Qd81sXlPnNf2JbFJlN4SEv/R2wOkCFhzrqs7X+
meSDI4tmyi3AkgeFdY1/SogJjoM+kvmgN9LSxV+riNcMqmZTpZhIA2oU6c8Q1NH4
sVtRRPUNQqV1nPEBYNqrpxgcS9SwU+g5r1TQ9orkoSOa24IMywdtLg+ABJwJJKwR
PRIGLdY//Vh7Hk2s46m0kqP830dQz1Pfqyg2hFm8tdTvVwtdu0lOKv26vVg+1Hmk
t6H9Pzhxf2dd1z9F27Rf0YhJfiEHPA2PplBUGMOJbcBRN8LdAJh/73e884bPI2Sd
p14V50VHievFoyTUx/FNnonCoGFIXGB4M7Y5Ef11bnBjzmJdt9BKXXrq5EowbOn2
VYJA/mnniSncotYhiJTmJb27s65TUDTo5vffddvBW9ZG13QBgoUfz/7J47k1FRBI
EWBRMWn/nmFDR2sHez2C7CRbniO8640wSs1z/0x9ZEGVfGyvTfsLvU5k3LGJHfBH
WY2dG/MuJQtnsaFNAY9d1Yz88M2pH00dbmBHmoakPD7zWGsEPJruBNhz1+aSkRNC
xt25Y1yMiXKF93mYWfA1YX6fmBFAfHeoL39GVBmQGahqGVIpn0Z9ACkl8qgxmlnS
kxP/ZtwqtiFtv1RbQs1D4kYgtHqTq9BDpZgHc2yEr6vVZ94iEWyH2BN671TXW/MM
1vByOSurEzwDq8T9gZPFawGOL4+Ega7+YXiujJynmR/H5JG6dFpOv3vQ3wk7t4vA
Dj26l+Dtg2NmncDu6Y4OBClpINEd196dpEDP1ivQ1CSIkouVDV5m0KZ64IzgIhEv
HsixHVr2wKEJ84wjhcQxwalf5AgWgW/QPyWuTyXpXef/WA1B4tc5DfYhBEjs/WNA
z+OpkA7KlefEib66iZLuD1Cxf9Nw6VTXkZ3uAUsnE/Q5mUStq+OaPfH6BCcZb0lr
itaSyTJs/lyIg4Ez+QmLEcLU/yYoodFi3BraZb5qCSHsBekAc85CRNug657LqI4X
BjJ7b1XPKeVhNf/aiL7Dpc9hmYHnjOavwhlq/PTLW/3/I8reJe4k1ZEkxPYQY1lz
jOAkV3hoEf2ziTZuVHyCcoHchWBzF19O2AT0J4cBqEuBpgLWQrhsFXA+bgrphIEm
Rwm5BzcWKqJH4vS3cCX97ay69ATqEHigi13RvkalqXML+w7adBnL916I47ZhNT2P
UZjWjcFEjpqKmZkKsStuODVf3/Aamvevelxd7WaUkKRxovhKTFB0xbt3d87LF3tb
j3wynneK/C0f9G8ca0FZtcqEH0TTlip6JS4tRFAYYLXs0Er+C4k7uonuAiaLu/y8
8Q/MG6xl40KX0xQ2Czqr2mvuYxNNE79S88x4FDZwSOpviDVKUazBZ1cSAobR/i2c
J74D8bJFDP+ZTTbJIZovuMHLJFIPs3etOsczRIEvNFZNmYVvob7FNsLMFJajWPUI
fJv6roUi+Gqm7BrIId4upj7JM59Jk/dRfhOEGXhJej6vtiT3r0inGpwkkTVq/fSp
iUonL81KgzSI+mgOpr/BXNOrpEwESBZ20F0JUttCSJdke0k2NeOUmoMqHw8FStnC
rT6NhezoWisve77wIjdMjMqn4eSRBxorux6FoT+GqOOp2mmxkVqeU4cJb12WB02f
8sw2DXdhfraOBWbfxzxhG7WKC19wpaGTzJLL/HAhFsDdI5WO+KklmHZeEdZ86S1/
vw3n+BBW/ZEtlRpcXq+VR2fy722a+z+jZJ/5zaH1bOvs7Mf7zU0YuOPMuhXDmlRl
5oR+9YsRkUvmbO/w7gvMte4eEr9g818dUnx9Sahp11zgkxwlfXWjHyt+Vn+NuAc+
0vSOCzQuTpmFxnYqk0+FwxB94Lm0w2T/jP4Jcp/3j20wV5hF5CzOuG0bM1Noknkp
o2HcnEIq+mu/cw1OPgP7gqWKgyYr8NyhmWiYnuuJkw9Ln0F4/BPUEtv4VyFzB6aF
T2jVkYaOKMj5B5HjWc84s+O6yEPtudwSBlnHrHjCwTu6n2kDwCE1HC7PRttSzm0A
4hD+JPWyFO6pzFvmtTwKD+pHp3OciNouEWf/t6DgNxmSaLzYK1boBrIWsFV9iMu7
Ml652iulrdo4JXqMOCZl2jTQmM9UMxie4L3y208HIHPNQaY4ufiLYGNHLjWR2yUA
UP2q8jZp7UBODEa6ZbNVkDRoWOykcgKFcmfmNjEuZZYJUL89eEXQ1Fw9xD9QeM3m
ySPAmNiUy4J0JcQExGDC4kZlnr+iqTA2bBew+U5mm+pnF5zUhf1RiFygeT97mWGz
07J9K38qw2XJ/7idW9KkuHqWb0nDKqNJUIKI2jNN652D1Mg42ZcbnZyN5B67fTwa
4hzuy/8UGQyuM1/OsAlK6OGuhEoayFFvNTgR58p/yTDvuHkDnOPEa68WbqKkkISw
HDJM7n24SAOAswA9/cRnWvHTS8x3v3UNJsYyOU8z8jzcyAXdj8KWnvUipbNW4PqZ
gT92LmWbXlz2eOgRddXxf9tvu5FPhC6zyRuUu57TmtdHk9MXIxPPdkdvPMEsnEEu
YQaCpczHnL/Kl8fWvlDkzZEFm4S2AkNr1QiIWnBGzM4R/QA0qms7WLIEGGO4YqxH
dTFMOZUmwyY87HkIcAUnrXWgDpaqMuEHLAxkAjqdXKDSOMw9uJcIQl2jmj9S1b6L
HiFDZM/5VVlo9VFKH7pbqo9zfAThzZp5q4jUQwfmqVXezKIYdxRLsjJH4y7pxJ5v
KS1dpFdzQUoSWWhkt+cIV8hY0dSNX1nPCHNGn31VGLvmTun4EMubcy2cn+2r/MgG
aMmQJVhjj5/DXNQ6BQD6VsbswuiYeMqzEvFGCVn1o925yZGnO6IQiOjLfSQIuee9
g6ua6+v3xF/Sxw6tH2XJSoBZCAs5CUAIMDUGLJJErptad0M7JWyxvl4F5ks8EgLu
Ch2MHnyI1Z9XDNHUso7KH+SkfKKtaIBOjcn6696QjxAcGDSeacPdMyUGmLP7vmzq
ygY8UfjQdTBygjhT9Xw7uyWayjFgbX4MgkYziF/S2GlgJ44ACgvH7CW+LtHR/Rb6
DhRbxxXuJKG6rzpwg9u1iEd1ZePP1eMk7DjKCkq5Hin9z+y1n8gimMy3O/xISE+T
TDkK4jgf9wx+VkB4PFIjmYXytp8dFOA88pDE9d/ujNmiw4aXfi8JQlm1hgSktuIe
Qbc3vraoQ1xtQXlIHs52NpMkGfx7H0KHlLRpK+du0AXi7aSeJr/3id0QfD54ScV+
IB0AEQ8N0ESHVaYkzsak9zlR1557xKfWIkec+1Y6UxjxQHLIxaK0QBJEApfepDvw
fygKKc0KWl8fke9td62L4DjJeFfcbE/SfN6+qCSgd360Q3v0V9aWLKJRLjAP86oa
XjljWzt4DbjRqiTAqn/467fSl5Uvqx8mtxm/ISXbz933MFfCUg58YtUAMJY1tki2
qhFeWH4Hqx7us3rR1g50H652/tHF5FGk1JvluSCBoKBtlxH9UVcbFCNQ6WJAwmYD
vuqKYBGy0k+M8cT/3bJ3hWCT23JgUfq84q2YnKlEWDq9BxRXuphp5MxFq+gTVbwK
AfmsMk+Hf5uXPoZeqjSYURi974MvHRy9fboq95qniEQq3PbZ5OtAddtJIe8Nh6py
Fb8rClQCkt+X43Z7N8CHCPDqImacKzo4zaXp5q6AE881ynkAdJ3CYC2GSI6t8c1n
EYpWTNkfR8mMwAOiwMHufrbqHxuS4C/KBkaFZU2U58u0OCtNGvlK42sXOeXYX2TY
1q9yNf/dk3GebDMXLig/IQEvCqwlTmx/usc1yp44miUgwR4rChenlLwoyHTb1qcA
VIn2OQoNI0z18RSOAGmzsEx7QFD+XUBi5OO7jKNjNiAHPywcb2p0kM4ih1wgWkNh
0Qi34v+pYSz9udoGMhvItOMTQ3Xbf3PEP98hBNWicO//X1OnuTIWozvYny/hLpVX
kfHPmSXcuIJEscFJPVk90QGWjPgCxdLlJQzJQ/3d9uN0edxF/shoSDOgQ0Lqg0OY
pr3amTwV0PMqjfFd6b3uDZDtrwqdIpMAjc7TlY7ha4K4tDi9mMJI4xDGX6EfK+ft
kvSYpW0u9oUkSkJOfFj/jZ6Tamab+qgq7NycWyu1/ieSBLNrDdFn3l/PfjvBnKx+
KuCK2DLTO9f3/GdTZaGhE0yE7/+y6x5b4fWfJg7U2uIa7ZkI5Ifi4CQRQv5EC3k2
P688mzlRIUvUsLZnWG5WYXmlpvuNq6EWeyKHZnJ3s/6QgIv6orvzQUuxw7kLV1AN
wsaqMrLewgPY/yb0rx8n5rBJU9H8J/70fwmbeMGIGKhjCK3B5aa2FCq+6BRkpVcW
cZ5VbjXxXLIFg+CH6JTikpU5YeUdpgUyD1aODaqqu06g+SZoAe0CzdSjUXTQq8sS
bJxIACqmYRRtH3qZXRqeSEuK7oIYJh1O32dFYos+JvrxbPMU1Z0bzLMzjzwixkcQ
OT3AJs3UuWrQ/Hisb0vkO9TRc69ZvwtnMu65q6YM0qesSsbJNkjptJJeGWja3Dno
3x5t4YvvF9C4UYqccpCSJOb/FxWDchR4Ma75QImOSipD1uevZ5YLBA4ibIfBSvAU
GaQK2yMwQvOjQxc8XGkykDHfZ5sCXwADtJXhzBMyZyvHYgBbraHBJlnJ2mtE766c
wvmtrfR53dUVMLJ1A43hSkDD052x7Liwr66FwT4dVCmZFV3ReOQZlN/Psax1T3fs
BsNnWShzgBT2m6yB6s23YPB0G6NYHSSy+mHWB1BIydzmwhQg2DjMx0Lu1NI/0KBL
+Fb+gcp69k31VpLfT+xsGHSDUCLtXHDLCQ6Y7Hi/ctCIMGxFgsRAdJjUVoKhhnu+
MgBApq2z9J+g11liBEpwFaAdbpUuMSklEMiNSZAzj02lVifzk+JkEFyGqOPj0Iok
2NgitwmdddxfwuXthSeGBVpGziCQAWtHcLf0Wqzfc79G+gpZJc9tmx5kYkBTV4PR
PN0S+TrYOvvD/eFodQB1FGo8PuQiU8cNm2NWII5CfUGsxaRjxD2/CPgZp1yZMb9e
GCNOQWyanUpMxYoUsXkJI+mK8kIdlqBKtF7KYBPE1rcNZ+L9JKo4qzbaJMj187Jq
WdsGtYOekrfiLzxINcqoUhXNCtWq34JXV83MHRzqT5HDvxoE+Z4I4KlVA+66e4v2
i4pld9PtxJIKxzOQ3MzS0MI3fOv0Bdha3KaeIttPXM2cIZUPar2+aPhYlmL2OBrk
+ZBwNqkxhJFAYVavqs+dUfIATjIxm8R9BncOATEcL5J5ksEiqTsnNsK9FJzFE8WX
Oysh6nUJV4SQCLNle22WYexpTXuaW4tzsCAwpxL94gUFjdT810magaOh5lSBq3Iu
PGLO0JADmHxt1J9DrgPYlPY4eueg9CYHIdNiZY3XfwnOlvQFugPxpIdpOeL6gw6Z
bBR9hQhAqJT3NGFOnAhOjeQHBenBJsKaJPSO9WJ1HMuj5GSOx30wGKBS5OiKmyVB
FT7MS08c0gF+IVB/cA7K23Ax58qZy9sOxaZRrYijFMYYoqiy0/tFAysoE8PlRrls
afYHK+LGg5X0+wGHmJWGkY/7n/cWNXeurQPnNfdIXSV8aF2JhkLEArm/XpUCIXyA
QLiZEgVBiH4VbrrfZgwvMMqjIa+HaOUeD6csInPCz7QmVqZV94uZkKff0B2lseO4
Mh7KjPSWMkjLvi0V1l8A6/7c8dfGOSo1dQyptnOj9wFnnHMuRTKr5auJtpuGN0uX
cryAM6c9fXFT1aCsaEvaQ6x62aNJ0KQljQ1DdocAWKknLiPjuAiZKJSqV/1OZ5SC
THb8tfOU/jlkD5VcPSW9QowF7/minq1UDupAIDJKkHeAtoAYiJj+M7t1TVcmW9sa
JOuc+aoD3MZIHawcN2O18JUm6wvaF/lEnqVlArfHa7b/WycDhbo27U86iIxLoNSD
WNWRd8IlHy9e9dKsZnbrE+xtsY97E4eaNsDilX5G0nMp4fPwH+VGcUb6/+3Zv4lo
5W5ss7PUZb0HSXCil61ftDOeF6cYCLwn0JAomSnJkomAZMHjW8uxhbdlphvFrsXP
VP8YWrNcjjwrCiurGey93aOP/YvhVw4K5DsUcAyYgbGsL1G06OUXLiTRT5ou2UYe
x15OV6Jt1kxcvJBVl3jRhV+4HzH4yYQJvNQJvAfE9GLv7/EiB+HTxF+jqV/B+xLw
CXhvFHIxaQzVJYChayQLac5oqN3Mz+RSG5k6RmWLiR5yDsyr95rMCGBjThsiAq38
fjgveLyQj9NriUtSN6Qyfj363DA0Nad18lnPXenPNs8kVVkJGyVSmJcWDKkWnBLj
Avw7Mr/XI3oi/08gOkaBPhsIc1OaCOlctWr0juOxRr2PAqynWQsnUJoemeGtGMQa
itBLrBMQK/fu+kOJD2KrQe0d+NBAAUDTgK3GJSOWpLu/bv5SvcZ6VBjgGYegEIRC
eQNEUvfsRIrQde0dLvDuez6c9du3R8od0GwZfgHKPJEBppB8kYsBWEwCjvTe4Lqh
yMizU8RIUNI7PFTnCn9hxqg9/1WMRQI2Lv8dPd6Z+qPSruHpr8hcWpaJ3N8ocbZM
vvO5ZBihBNSYFtG3FWnejXMd5eVOghF3j1+V7r20Jae1OT/l2mjT5WFsgHmMemCq
uBwEvVWVeXJ3PFKiKXnoKcsrR1H1/N4y+MMdN8P/07s1UJ5U/3y6QiDZy/0qzQFQ
1Bzom+RAxws5B6kJosfWzf8lTIu+763bywc3Rrh6cuy88fpzCy4ZhZZ7eBIpRjqw
6MjSGyzpvgbt1x8mstFhE3wK2l3fSstnEG5E6BlasFLiHchh1f1MatTdIKj1kIpQ
TvvgzJxF8kGZE19GZI31xxWwvcVYdFPMXO4ADap+LQm3gvJH8317T3DDRd0sw/N9
/+G2525i5JKIAwxh87PPSv1QhHpg6e/OxYu17uiBLh38ZkAuCB3Iz1GRu0ptz2lu
g19Xb4Glv8kFWbBbN6ab/9pk27Y2C38Hbu4qdmsJN6fO8B3YQDEq9aJEh/Z8Bkg1
FBZDVnT1qFQQHcZlJ9ENEZwrVU/IR8xe08N3aaR7XRRVHXXQodHQ/lFoN2MTXpeY
++9IWDH5bZJZnB1RNWgUJlOsfAVwD4q+bPjlyYfnxEMZS7sGDPozGtnm9t/weH3a
kM3KmUNY3JdHAwgvBL/artEwWuTb5QIYB89kHyjubVHcN7IHKfFV8IcdBJzY2Llj
IdPuU4wO5eWwFSF4bDRRwP1RwaCx97YyK+ccDyULH7sUdLK4BVyflnLwM6E4sgNv
bZaq6sKio/sUETFpb5YBJ50uRkLrXW8//u8v11k3kg0I/8ldEi+aa4DcOYTvd87t
4cIx2H1FI2q3AgQeHjKWiMVkg3SkU2Nzo0tBbhkt8QsVlTBdo9kpBQ5lKa0iMZgV
u0vrnpYjlWveF8+Odh9CjrEazdCJD35ndBdvSwVllWbo8Dv/QUXMchpOupl7NKaT
ARHNJp3mYrpr7TzHtFIJX5MR5yOFPN9VR21PfrnHFuli/4wATVjvF2o86j3Dw2Rs
489LxkmFJnYko4vD9oOEozkSaBwIyrf3S/BHL44BlZF8/LIYMx868ryeJXdHvElI
GyFuuNtmRlhQ/ZVHbsRbpG9nHRD30eRIyfcuZiMnbFiYoOjXGFifehIj+A18DaMW
kv5NYN3LVZ+hTWJE3E/YzmYsW7h2dbWmGx14vJiygI9SFe2ufw1zv3l9ChlhjLgC
CExLxcRpWv39BcvkP43i3hCkum78HwJ6D/ED48Q4fi8xcotd//hzreeE/1wsDfOs
dBhSUOYUf2kOGJ6Odx6Z7AC6JHEFhA8iPqAp5WqqQ9XYsCSWKHoiPNDXCFrVB1Y3
/jc46724/9NP96pvjOEtnPzEtWTpjbB5xc4fYSusapd8eRLMVvKcFUbClWF2Il9K
sFp4X4ZpOYTTuj3I3k9X187LSjpEUKTcctadJZhO/a6Yilw5sbLzMMwjJjH2SS++
S4nnnP9fyscDbq7oq5Lm6g3dsev4APSYuCjPEf3D+Jgbf6iKQl+OSiaxL8NoI8xO
Yiy2absyTADkla2WpPf/mXz/Un2aDnOlTi9pUZ+peOLLl76PzeMOderk9nQxNEYo
eYHdSzoqgcQMII5RIXjXrzByt3UFMDy+wp7+WDIAVeS48N9XROfqmccKFaBvazCz
NXOdlvxVP/O5P0HL5mf8bCQ/e+ZwVkAOMoJOzvMeCcWuytEzqzInpOlrwhlHkBVy
3jI7/r7epIX4lt6DfYHL+IKfConizDJeyfRDt2AG8gbEvMkX4oQbCsw48ST4y3s1
QG/9purt3YRNNpLnM+qPtTtk7+Bl6qzBfkRkW5xFggdB6c1RPzWCVjT60CmbUY2E
4bVo7EYFiL81Jw3/HknDAK4+8PoLhJEnyJx8xwIFrHjvRMb14ZIkH1pPCdFxYW/D
bCS8dRj9DcGltMWZRYHRSOYs5V6JTCZ7Ox3rjmYmK1ctlExWF4EDsCSXKpwOpmxi
2WDed89hK0b9K1ZFmn85dGI5jr6Lo1TQU6Ww40FsuOQ1Gh8ahdAm3RXtV++E3eWo
fXo0xBO1frDg/sI9rjeaVBpcoKG+V/ZlCh8ZDgrLxrr4Bs+UZnWZuZTNAbty4Nyr
fjL7tEmdiX2YvSwdsNtQoj4dyxAsS1J9n2HUAYEitbeRZLQsSKo+zea8WLPlUy4Z
a+x3vh5Ct02Zo+/e1qZchshN2feHn2mspyQfc62uPJ8etnbB4gZ7A1dzw8jg2USK
0ni4yOX2dHElPxubgE4OxD44RHAUbHbqrC3tAKlDRLbCrjceYodD/qzrRUWppvq4
w9M8saf6lihO7Bf97BOyQc3iXyrCkwTug9QTMRSAcLhwMgINdgEn/2vSztIwjuaS
jciPJX1V/Wff+PEkPd7YdbW8iYr+sncSAl0dmtXCcK3btXsP3BHcn2701nHBNY7A
N+OUZzqLszpoAPlRP8byqoZtNv1KgqvWbD7MWL8h5e6Jr5L2TY25WIjwNdB75ugD
VY4ijzFQMt1lLvsbmLp1CRxbX4V4h2esLrbwuNTJwQx07pnBGEbeSq6wv9ezZvQw
a2RX3Wnh6kZhUUvweaYAvySx+ScW80wkDe+DWtTCtrhRF6y86+TUdFYmYit+zLJO
X96GJjukCvpcQLsmw//6fwLrVgZM2nZTMyxrk1LIEUEkb5U3oBDbUukxamtcDrpp
ITh/G/Sua/BVXxIEqiZM9BbHgjYGO+nGHLZS7fqeAbd1qeoBZaERNEU5HlHNBrAq
s418FRgKfu1WkOPE8iLekT3Oiba/kOKxwlnPCdSQHR17wNvbXtViZ3YkuaPm2TQx
NeLU/VqIZMKsC8FuDbmv8w==
`protect END_PROTECTED
