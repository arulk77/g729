`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOvBMLxob/Tq9Z4PZWEoaiztHjXwxTKaeb4fv03fXMnf
dTPfYadbgo3/70csEeLTCvRhWnBcMXR4FD6ilTn7m3dtTNwOdLyEY4ZTJOR6VEx2
AtZnyVffeKPbKqOxRnduYwpM46kg2R9SKOVBiTsQsB7elnx1cS6ZMJjo5bl0VhTG
mJPyDXb/ynkJNwttAqd2NClzPotEEDERdDfbm+5bHoK466DHdF/Ud4PWJKeSjVdZ
bCGo4qWW37EUkl5GWHJg+XXlicvmbwF1CjKHzmkOYPiW1jQGMh38v2FivY4irCap
6P0WN1GQhu9TBj/I+KE7MQ==
`protect END_PROTECTED
