`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48IZ2z/xI8QiYCRYDCJI0hZj5dR5kedxsIm+bVxNTTER
BuP6jqX7/I+8lDNDpoIb2tbQzXD1oJ78rPDFPgn1wu+temoZpr43rIciERDW1bbw
GfYKuiCjJbgprF2Nd92wmnX98qqwn9InJ9tOQUxLek34vG9NaBT1DJpa9ayd6Jke
YVMJ1wzi+aiDvUOnNBphm+PdFquud6cxnYd9+Ry4/68=
`protect END_PROTECTED
