`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aZNRnQoxpSrcnTtnOijVBWhA2g9VIMK7kFHnojaajK48
jZXe6js9bULxyCcnAIqMdbP8eA0DgLgzztmra6mu7IkDKUUByogGjVhOVoP+JxYE
XdxUPFw78rBZRiaAzU7WG1nsFfffzYvour6QOk6BNAsU6sAKIKZ4fY1qjAyGyIPd
CVG3iGj2tW7pKpxEEo4AG/4i6rUvlKUEuDR/IglTAaQloAUqJCVpoPLXI1a/LBUn
DzKEg2INhXCEShuRxaWHWiqVzuqM6kNKM6EsVR1EM4cVrpIWy6911Y13CPUlSkbn
BVAdJBVZVw6ryALkcn26W4goa6ICgc2qW19hxowqZimGKtTZzMMEMbSvSlQ39v6G
ypBL6+GM8Zg99fdjuIjeJeET3hsiogk81QJJfdX3cXuKg1tmzLyc1x3MMfxuV/HU
`protect END_PROTECTED
