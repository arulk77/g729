`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAIwK2yciyQT+8QbT2oAccj7RAcWObEZo8AKfBMnJdQ0
DolobwBHQei01zBObAopVVygk5PfQEsYcsGNpZNgYauhnfCaa3a4Il+N8Q9oADOH
jpFRcKIVsQZqUEycU5KudVB+Qmq+ONfDPlQCW+CR0sv3offb4Llj0kjj/9XaEB0s
59+MdOWZD8x1Xcw4CcSbsDDrdevn7eEE1rg7MDTMAg3OqE4ofpX3nvEQzypjtVJQ
7TLN3nNtjCqP4BftJnOIIg77MnFCGxS9r9P4rgtsbGda2DT7euP3wJBPRYuJhOWE
Fqg6LJS5ZCeORvi6PrspoTBzxxDxJrzreymW8Vuu79Q9Kzu20DqyhQHXu2iQfYrz
u3M5dO0FN0to7L0VdHI4mZkxdxnzfnX6bYbCgFpeeqKCd9wE6rvZ1A1GQKKBe6kw
`protect END_PROTECTED
