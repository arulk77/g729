`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
adbzkDZFya55avLeDhCFU2pTe9sIZKgdHku8eCFjB+SiKs35hGA5Pmu9QkXGLHIU
0xZ5Xa4GjLiiMAi2b7KwVVUFYILvkILDsrVZXSRprUAVgGvJq481cJHmF/1vPk9Z
E1H1qwmxwZ4atCXFw/rSX8wEZzJtROdqJLP63z0ehUGbtQp0Q5WDRgr2hjtDvlxM
`protect END_PROTECTED
