`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SU4ZhEgWY/QoA7WZkf0nxYPaJGcfGuGcl+1aXZBvHoDj
ATtEbqK/+f/sYdF67Tf+sWqcUouRXRWaUpItalhNFjb3E46Il919QQkt8rqWZtHf
wOeh9AL4t/mP7f6B5KXCl2uIWJ6gvjg0Li2ugIlwBryA8ekB4aXOATJ83Y4CXYBh
a/4CMb8UgbQHpQhD8o56vejk2jL6QnHDoTbdBexpaovWryjP4WT4swWIKrVk/eB2
TOAU8oqmJgR+qchT3I/nYxvN6z/HePWDUexsFVPBLOWfm3AauKf9vYztIGlV1eSZ
MoVW3URw7xocoVzcfSh0OshUfmmU84tudng3fKdHGTkLltK+7MTzPDsZk4OGmqBr
72/pZerDjSpH1iVbm61R6VqjFnAdSDsOU1nBEB2LuQ32G7lsHAFjSqTWNMGIzBPY
N21RFl7G4XasMaRhHsvC9eKKWXvhGSy8yC4RK5CRWzQy5PtjL8WRixx9UU7Xp/El
vhOMjazZhuDrbDKtRx+g/YyLEaYfWIwoSergl5aGe99i4uhCUTHEJk5fojxH3Jkd
DuJGM7KT3Ksa8aNIp2/bS/2c/UtxKti8P3L3oeBtIT0A2lmQNbJz9UVE4QLpupZN
JEl7KFgAjuOi7Lligscf5DRDshnaeZvxRZ95U0YXTqS8VDIN3ee1TJc+nr5peJ7c
wZeNsi+vFzcgxe/8sMUfCjPKRaD/CqKeDizKtrz3uGGEP5zKJ/D12mnQqhgiyLsH
/NhHmxn3FRp0vwLhYrm/hwfuwzF4IUBv4L4bHav80jUDpnv4TGoA1dMI6pPJwQVb
HvXPvZlDOTQOn5gd2Rx4TB1+aWRw+tWp8HwNUqX99RrdZw/lEqyu2PuoNLw5Xr5V
sUABiIjpOB8GdiZbhRzmUYY/JsKpHKTTOAF4jMZ0tLTJ5Loff4G7cGf9HDW42yvl
M1EZ5bkJFjIY8jEuQ9o8Q2EXSlbqoIMXQyxD9mpEzuY0+MwbtYeNET5q9YSwLYSE
wO2G8Hj3Xq9H26d3DvP1oDcwMZUePE/UfLK6m1tWoucdFCuop6Z8PhMmAw8K7Fy4
MfuNnHWzL08ksizNjz9hexFejGbbQ9gAa/IOaLhtuaPhW81Ht9RSQUOXj+IlFAJM
cJChKXmSsbUXQ3OhHMCl8d1IgRU03DjxG/NIuv16QgfI94Ux2gb7jF3I8D/iw4Zd
`protect END_PROTECTED
