`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD3toDfK9CAIswk3WRx8JB/gr4rPChtJmesSelTM1MEZ
P0IwFwNX2xPjVdxWoHd3BechmwtOzfJfEZp7ov326Ny7ugXa4HEITtAxlDNvVXHJ
jGCX1arlIHDH3aT6jrioyNWUw8QTbcgrx/5+f6lpv5hKNthVOVD/uEOqszS5UXJH
q1eTPPXRfpTeB320cQ0XKbooVZe7nqIJ7lMhx3O+1th2J1W60lLcUcC1GCVjd8ej
QdH7Ll7JlwG9wf++4kTGQffjulMVTdnj5d2puXLwd0w1s+gRAA0P/vuToOaBbetv
bXiUhgr1RJsnH6ZKfBNipz24O/Dp7NRn4BmE5JsVl27rzlnZL514W0pSXOe02hJ4
OkKc6HUcEHg6YvQg2o03dg==
`protect END_PROTECTED
