`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4hW+SM1ADUh9FO//GIe36ZrkP9PFkOPjAsNomr3a8Nlptw0opUMksbj5sSgqMjtw
HzpDmsduBnRyQ3qJJPILTonGw5GTS5m2969M56CDTmXb9GGCuszXfUtHRxW54E90
d/CNOJ7u2OGHsT7CQT/VHTMDJcHz6bQU0g6kE5CNpW0BJYKJSvkvS4wG7YFbaaoe
mhmodK1WYxjkimxX2Th2AgV7otKNjyfIFzCNJrZTtPIih5Fn6qt9wOxx5rveOB3S
+ZSwK2VXAnn4wBl+lbTJwdbQ0x0hATmtzpihsw0gicFyodJDcN/o1ZaSQTO7zHnS
pd1awji9xnExALSS42oew4GlJ1HfivbIugVry3wMlXyt/NDyrohdngUt0bE5h8ev
KjkrDoP500iJV+2lBVBNn636snH4GhOOLHPcQeUQnqPfhthG3wS82wBj9jZKXXvC
9Blxfgb2yE/iivZ3Z2va/xIT8q1SPGQ7OLeU0Rv2VKGaPvtaezyxpXzqsXBaXUmO
fIORPL90oJOu3uiL9wbVgv6rfyZVdQYmduHefJ3Wbd+4halE1znrBUjkjLvMF9mB
OLakuMrbQvvvj1PkckaSRW90Y7ivFeEB6flqY0/pBhqp4OWIlxxlnGU60lDx+Z3P
MFR5AOKe6Et4dvJzw2RwAO7eMjKRB2tvWrowtFF0ZHzyK19asZQh4F73dU1n8TRu
UBA1W3Zs6Vfw9jhe93W8uDXG7laudxJbrF0AGUmtmj+dYrDwBienTAs9XDr7Ot24
`protect END_PROTECTED
