`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
gelQm+1nPbcmrRl4+p52R2thWO9kDrC90vPFFuylbYYNoJLHbWveFxkql2n5O31N
uMfFKTrIG5y7zvFpd69q/ZeN1SFAMpXyxrJmroeVcZloPtSowvkkI7H9VkYErAsW
KeosYnFdt9PWqJ18TuoGBRY0HHwMrCJmt+dy9cKgtKytW04fC7mV4SMI3jMk5cyy
`protect END_PROTECTED
