`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveObkJq8ygWKYz22EMFyOobnNWzs/LnmocqoKry/kWXyD
Fs11Y6ypotSDWnSyjERtqsrUa1QsPQ6VIcdj6rVdl6lQZvZb+6VKqYV9JoHRiYQl
Sl5G1YXnx3O1/CL+U8qzDhuuzEH0kNCrt6jhN6WZi/45eGqN8+Rd+xUsilhAoXKo
Z9q9qBBRU9osTptH+ZA+DUdhtm2hAuskOLkMN90+6/UZjnCBIIAqDAhaAO6QUi90
NYA2Bmg6oOGob9vUpNHbE24dqg1cOHKKSc8s625pRFDksNIyiuxBXSRge0mDf18j
VDgM15mEVkghXJdozqBHmL7yhSEuPhT/HtJNYCdLlGXnidwwCLsAEFYqI7zy267G
6lYkxexVk9zgI9VkOtR/EeyIsA3hpYk45o3rwXJKvxYu6hcbzqQj/4KKRSa/7ZsC
njS1v+5vopuUFV4v8pFMAJrukYWRPFkfmPLhBKgyEc+f77dQ/Q5A2xAhvQazPHF1
p9u6XktBycrGIb2uf7XsogLNrlVb+zfjyAOmZeqM5nIrRtQIT1FKmgZ6l07WT8ls
`protect END_PROTECTED
