`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
dBLQhQV49S+rSe2ZvL5JUswrH2lt3Y55a6qncqbdSulyXvs/0jDaoAHfeUAVlyf6
N+B1QI1535iBWY9mO83r4KjR5UFgOqjrm6zClyI99Avu4Y909NdYUw5jGgkvsXs0
ZBmKnw3YYkvPqJbmdJWTchD6W8nq8OwMQ5R08f7YcsirISKzrugbaMecM0oLUx0L
UfzWecNM4ncE2apNRFWq4cahLGTgP+H5062xAuWgAGmRiLc4UsQgXzAMORZcfLAQ
XtROUEFoNrrIUZTe58HrpfVjZW3UBKM72Qk1RCbl4A0=
`protect END_PROTECTED
