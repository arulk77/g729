`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42pMXMfplN4rkXrcj+v1ZmEREAWK4w8vzIYFpvxotMLU
9cvnsb/UT0A+FNdtI8KopIrOFGtWx5HFCr+L7ZmTaOP2sjezvY7o1rY496jzqxDh
ELgOgKNWnBTKONAkPq709r9p31ofXE2HMPzicCVuvPStmUBxSTc4BfPImF278ZqZ
KcsEAlrsmDin1FVBcieAbVDTfKdQtll6hbgxLzDJkOtcciZz6sUr2JTmc/Nln0HY
Ot39x+LPwy22GrAJap1CYbBHrPIMmKdYtaHgPhZ12fs=
`protect END_PROTECTED
