`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveE+beW8IYMDaVnbsoSac416vTmTjrWzouYcoMLUePhk3
pothHrKOGZDk8CoNR54B5KUX9EeIwBXPfCKaSPJcigpXyg+rpqdFNby2R5+i6Qn4
wfo0GO6DQylOnfqthuBOsCrw1RmQyJYneTvAFy9LD6jmSX453FiHKZnmQJLEzm8l
1HZf0zJ+FC7b+GhYtN/a80B87P++A8MaMKEnKeUm0VbhoCeJNWynblQjxNcU/h//
GZZ2JTDSAcx7v3UZjeJPB+6rHP8zQgV7VkBbGbLDJ7wEWjDb5OjrbjoFDKi7Outl
ESSktRl4eUDUf03Ftm9+5hPnwFGYXJrcUPHPd69CtvqFO/W83rnlFFau0+1eLhGq
aKkurx+QQSbbX5m77uabkfQPmYyWpB0B23oGX5spSZ6rWUn76MDYjGXEgdb33Ym1
OpKiBtLOg5/IA7ZUyZlAB6RIxDCK9uzGdGtBxugVxT6KFgjdSBl6ASrWlZmT0oBP
WfVMKLrkCGDsmwirGykEZol7FJUOeJWGWJh/POEQA6zwlRlz/defBfAaPMxVw8I8
S4Op+aNs/wnWhC7naDDlxooF25/R2putMIv60xY+7yfupkDNQIol8NmsK4KM/wGz
JgwX0wO/t5EDYUByPkjOGEEQNEihc2Un26kWAq8AweRieL8hBbw9Hk+e0+AqwCyN
NnLCFBvSb5kuVjvQNF1k0td/JYV2oGU5rV40NYIlgDykCf1YOxaI52J3/oIPMvS+
/L7HzX6g4qUI2wfxWtzUnIb8uu1a7ErpTop8T+hF/b91iqH9LCUDxpRJ2B+eS56U
OBXT/rcvwovv9wCReKjmfBAa+p+mEg1ndVyJ71BKqM5VgGou4sjaSWWXtVxxOedL
4admRGJyitKahD1eQwZ/Ivo+q8T6sHJt7yvAruULC6+OW2zFxkk1F1/E3QFFyYPU
EYwTaAOiQIaSb5KLVB7WYO+yuGTUszVBLG4m7iTrbMx3s/0B6fj/su7TdDyEJ+vT
Ca5inatyKohBoqEjTR8ZYAIdcGWQJFUEZL58S/L17ok110wrD33gUJ1QHkzHE5rH
k/HZthb++RJnYUyn99+twgP5Lkq34281aQ5lR3+iyOOG5fTNB8Qj4edF5Naji8Id
dPuEzITef/64ZvmkATmy6100cWtjCiqFaRkzlebLxHgDbp5wU3tO9TdBpWQpzOpF
`protect END_PROTECTED
