`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePDplQ40b/JnteJVC7rox5lRLpLMNkMLdZWPLMGrwY0b
qIt1kAzX8S3nHIXWwlZw2pA/KpoN+yU8cJ8m3LcdBk0u6z4ly2WbaSe+D0oWn58H
3QT0N8lNh3At/3PnSN0QyPU5RE2ZUZGqUSomAjlTbvyfAoh2VlcPv3HzWpmqIwNQ
iCVfsVMnCQeUJjC+e66Kj3DoWe1CyfT3yBfBvFWvlbIemybjADQ7mlidCnFFK8sx
td9Y3vZiNmhdbiMl6JRYMv6CSS61EJhsW4xi71D72yrPej+aWpuNIfbWFW6jR3gU
VLTtK5+LKjC05A1YdxCkOpuc8crYaLK7FxN1zVODo6oDee91jUGPXwZYQpn5ab4R
cLV3Pv7737f9mjTkAm556iksGEg62eoWI2ip0/4CRWKTbrjdSu61yuzNhodcxSS6
XQlk0vnN3emagB7QnI0asimxZLuWkkr1sJP+Pb5WVYS5F7DEVPIN6c0YSpuawhV4
OyXwH+HOe5mxGIlTVh2HQg6YV2oF/5pu6VDho7coopC+gWZ/drYsO8FH6GXP93tq
6o7YBCPrtQcYO8kbRAjTR8Z5HBhdNYtCE5wV/hXzMhYbUDzB7uif062TqKUmXZ3y
EL6DKVgVYAD3J68gmQvm3uMe/XBj2wd4UtUPa9aTRSrIPhG05eTOlHZo9HrLliNc
`protect END_PROTECTED
