`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOyoQ8deWQLsZHq9Ie/nmEXhteI3GM9eH0OhngSsIV4V
NDT6Q9KLvIRBnoiuZEu6xqLNcLp7hYGk9SvHJQa+vrx6F/SDGLOt9/QeRUg9ux1p
VSVErkjPR3t3LXbdUDD9mnfu8u/Al13xvnj79gN4k5Fjxh93WcocC4f1X6AXgQ90
hTNelwkeLaeBIH7QNKrLaVtnnzISwZE5aX0qH0031m73atQD75uaUJUYQrJDvhgA
sHzevPPzKT9En5gbiEvinA==
`protect END_PROTECTED
