`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGE6cojXywzI8gWwQHTnHE04pSB8z/c2nfTAiqu9OaBG
0H9EP1gjptUpO3CUus1GJLsu4a2+lS+U3gXChLpaDFysX/RNXm4sLSONH6fnRU42
siOUvWJyJlPiy8Wmf8mhEWPF5FoVYimAIXI8X5BxRCv9fj9v5wmLLq/nRS1DHeb6
wIYDI/QXhVk7Y3GIEczlE4QsBVgV428a3JZSAQSS+sBPArACbMiN95eHWusjaiVT
EBfBEPJXrvovAUeXx37disABC/+B/4z3cZx4eTW6ZNcBntAh6iH+48gLP4vrT+v7
arC/7DRXz0mjfUMvWY49tP8qTSoRBTk97nwBbuGHK5ZdM8g3AGBj5Dlg89Z8lodr
yIVjx/cBT3TdPfxJss0po5h1EVts8PWI6ckE4L/tYT2Aj5hqEXfEzjEMsFHKp4Kn
8VW6yAg2WvNyEkejrFkstMtCSgz9a0r6BsxAsLNpJTFPPhJ+czca2E60KNALW/VV
Mc0QMEkMhm1A2xMHh2coH7epnv0VYuLFbRPm/LAI6lu0T7FYcsh0r7MxBGnBEfqD
9HqZbRBVsmKkHXO64UoOLg==
`protect END_PROTECTED
