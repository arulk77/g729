`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAaRv4oL6VK9eKyuIZfGdIuBnp9Ul5Nq+Bod0KsmOAddQ
x4+eTHQ+cLcJIb4a/7YP/6PZJNbTW+hdGCbGxeHu4N+lfRbONKnEwofNequD3FFL
atqT2qeQelsI566dT8YfwLNakctZHUNtNEkbJLp+Omg+XEaIEf6kRSbVqhXS6hu3
+c9rViBxxG+Z7YSlurChZX1T9ynqYe6Fb6PiDZJM0c27P/76TbHUxLMKAA+HAe1j
6g/GIvKdOeeBghTM1ui4ICqBnEBGPS95u1+dATH0K0HbUl1D7MHatrA2X9wk58ha
7XKOvV5zOrglqf+Ln7nAIfES7KqfID+KWlqBQ1g7WKkn4WZimUCQAKSkO1Kj3yvv
LVVp9VBh1HlPjtCgK+XnGv3WdpODxEjQrmOfkurSavNpzFRXAKnrwESbaKgGIJLg
Me4xPqr339vOZkXZvw1g8XqhemIf/Ub/zlZkFlkAZIhYCGV1EGZ3qKJ0KbAYQiXB
1dGyw90yFxlYrxFrnfTTM1i3YrT/B5zR0dndLxY5tvKNjwC7FOQWpwbTcrRxAokw
JyKCK4ZVVGzoMl4l+imVIHMAdR9qmvJfX5esdzNKoZjkaG8GKjosxfB1ls2JjMHt
l7hEHkjBacRt+IHPrQOMGZPSv4e4+eXxI0vOO5a98bigSz52YrP6ce8UPBK8HWAH
XqvGZ+OpvRPnDZDbBDX0aW3VFVn86qvAPcqA4xLDjuDtBV2eUgIn4nuJlrEbh71a
WawU+jKXNg9/0mDh9lBC1PArWNtZxp8L5x4Soepa8hqXV110ODWFcAW4Vq3+POIl
j3xPO+3TOpHtkoV3Adx0Vzi4jFCAjvLeIiYyRx2Le59pLsL4q5H3YC5SHEfzsytQ
TQc1XrLpdAv80vFDeKUfarQJiXq2uxeEUlQG4iHLganqo0jucYeXDNznW08jaIlO
FHXXKtfJLnoqLyjKwMUBZHipL5+MYCnDROO5+4QVesO2iibDkSZG2YOu1JiI193C
WdYGo+awcyqS/GWosx9WiEvZsvnH8gHSMIX6VcKKfSnBBA7Vskc/oeBzoC/V4art
x9wBS7J73V31xtWpxWnGPUAOjpC9OgTySCQ5e7cqUCdwX+iziIshkIwQRz4uf0Tm
N+QuIvEhxGZopcnh5nK9QxtD3HFw2GIFWcxSWHYebRxXVXHWgofll1coZd2DkJEW
uSFrbn26G3srYPu6szMXnQFlQk4J0LyL2TCp1XLBv6WC00ackFocmU5r5hFTNCNp
pSE6Nx4AKIcYzvahxTP6cjuBXn1nbUp1k5NTODeutIPXULbDjxYwB5WclpU084CM
43o/rmp1wt5QHLo+GSqiLRuIe0rqfjGN3DMY8M8VARuxogZlZFRLgDxnkx8cgQGx
xRL+wxcNh57bMQVR3xFOFWmPjXnPRLl1PGjZKW9m32yyBas8uFwZihY0RjzjLX0k
3lXS9Y+SxjQSmAhywuEaWlVg99jv1VrzzGNUIgW6iA88X1dSyA/CEhIFRjpbtP+H
wQ1j1mcjNk3U0u7zqURFrpAMfghE71Q/jO9Wf0jCnkfhRGyv/eqFmSr15hwCSZqZ
PAbAK8TJEg1BlN9dcbukZr1k8MhaqphC7Tw8QUEHUnIcmM9gnM4pl45RFpOWuJ6n
eVCAWn5M3fGKEQjPz8O61fJvitSQHVu9WPRrNXE3m6dWj7uj5noRrEhmRvQX0e8+
P6u5689MftDJ8u5w0k8sRNpYrtlXBX62p34zzqTckX/W4HnMV3FdMLkDbivlFjV8
LoEXqtphvQqx6wRQtAE1Ul5Gb9zXqM5w/Da/IERcdVY=
`protect END_PROTECTED
