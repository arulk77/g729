`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFpYd30QEM5IYxoOjNbkPvCMS2s+Ab5xQBKq/9qi4Rzh
qTryZNM+wZbmz13m6J1a/fIQnlewnoQo3NVx1HxgUmIiWsNBtOH+GaTX4uyK43zr
WDuO3MZpmK8RLG03NI1FiKUogCAtlwwIYzGxuLVSUBmXFL9781pzg/BK4kPTKOvc
U6Eu90kpqTceG3QJRstQRZoVPE+Z69u5OBISKPHQj27D8uY7XtZAe4F/4+M22t/d
Jvd/HIChXN9I918oP40rsS/0LqOSTddxXoWlyYLx5XHP7vljKaQT0gl70BQ1kBTk
KApDV5XfXbtYxbYDzo87gDU7dIWCsJfnt9tfEPD6liWi80XQj1yYtPHzUoLiOv8b
4E5H9vBgdPjJWUhxVy6BpzsHmbvsRApvRjidaMT/v1snYFSzOcpN170wFtiFWZQ2
uRrv5mDj1p7XqL/8kvB0mkp2cZdnF2DDS7Yapx5qxyRgePbs0qDggnYnlsx79mmR
CmfLk2IZ7YWC2dWup7+q80ndWnT+kYqsjr4G4GFB0gEg3g8gXDTor+XVGg/A62kw
rsRzPs6QWpRrFftbgoRxEUQXnev2uD/6XKgG4D3WMrbSevXIV82FleZ7zrb8Ikec
x1Bc3er0E9aNrEwZb13zfUBDA4IQ4eVJjpUZAlr5Zxvn1NtQUygl6M8K3Ys9McHZ
XjmzrbHTBs/HrLvoL2uEiTwA1m8vNrx9NFIOdT4TL0OdVTdkcAkZ3Wq0bbOOig+0
PDUcVf5bpi4OqRuW3F8fcZqKygJ8c9XlBSgfOOV0EmbTs1K5hj8cS0ODqWgCRZB8
`protect END_PROTECTED
