`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
7RWERbz/SCu29vx1yp3KRBbD0haMaP6H6gC2idhw1j2a52qcuR/Wd/wT3b4CqPqZ
9zooS6lLNuHvyybP4LWrG3zZNhGWGFcuAlyPf473H52SZJfam9nKJxlLgyHmXg3Z
0RUr2oRZQWebjb7P+3nfwByvmJnp604nG+jriBicx+FrKhmVVPNtooZyktmfGwGf
`protect END_PROTECTED
