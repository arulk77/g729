`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zL1VWgL22qS1t1U59sxgp3A9xIzQTxfIKaT5bhzrQ66
iFaSYINPcew9vYij2kah7w34/dGK7BDvGV9MNmdgGGTUQedQeNeeUTKuCz0MZyb/
yDdEMZvk30YCT4umywBiitwyVEqdwPi171Gqao9HuCJM3lRK9vlCcN9hCWy32KLr
m7BGuoD06FQDIbye3/rFHCfrco1B3HwN5CzE93fCGcU+OGlKSMBce+FDHBolqWbW
VVbeQPQgz6aj3QU7ppE2ZLC6HU++DDbNrhBk6EP8hok=
`protect END_PROTECTED
