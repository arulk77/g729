`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
W0kpc4Yy+X+TYmIF7tJ62+UihkP/J7vsUQ/zeKuek2AVWgwHLN4ESsh8rdQU/iR9
ZPHXpNTPyRZ1VNTt+W33R9JGcEvScBwSHR8TLgmoE2GwnQFx7C3n95L4mzM/62/m
Awv7UBJYhiyGN9JUCKOSmtdtdAIhtcmIjX4y228jDUPMV19WxNwiL8bNKlp+YE5m
9vP2GH0e1FA0MvFkbb0dacZXOg8oO8R4rbxECwPJwb4IjLpAJKJTyt2JhPc4odHL
tiVO3LAMuBwi/8TZ5fc6bCLXjHcrM/dBj65T9h4WPI6DbJeLQ3c3l9ybkm9cgcfC
Z0+bSB0lMMQZ27ptopQqzL0mGpzW5j/lc59q4IbyBxc2SXgXQDfDnujbcqe+9GOt
8LABgPcGOpihztCbLr7IuOUvqLB8ETNpsOwrhPwm0YrBY/T3lBabEKAuFRJPSVkV
yg2M1loeKTnXP6aZvQl6ahDESnIbTZrHlbeI0Qg6K6gIqFka3ROB064A0eZNc8Q4
owGWgYOe1IsX1vaeQ2CpW7YRalno3i21NXIFUB3VhpnZSKFppZpMeJQ+wwHa2Yrt
lvxi5dkKyXOuUoXUo2e2RChlRBJkwZccSVheQnEL0FiDpfJHHZQGKbuRSwCazKTu
83bBwEwYe2xsYwBmECGif5aUkso/6kbTLMM9c53ImAOXbFFgNZ1JDqlbLaA983Je
lKBXDbiHnvpakZlwWTw3yg+Bue+MAyV0OmwmLOB2OCR36r5nhV29ZU81thLWzTgA
49UINFgxAXdHcr39JXjnfqZ3VwYMKsfgnA8c+fbM+t03+vQyTi0WM6Q+kW+18MnM
EQVbYVuAxHy+NcK5IPRls9yksGgT0+LoGrQyKo01MGE1madjoJQF0EOSfBqTKoTr
pMVnZvc9snAxNnbEhcRE5NxMSyBwTVCHScvbbb2XOlTBEjLlZ39r0pl6aIdRGzaP
KyUYuN+ifwV3OdJTBJPXUOApnBE7qf68HtrQXdzfNHwSQIsCXTHyXx2yJSnvAPKD
WGxH17NuOA52dPGoSXMaKANxVviHabmNf7pQpPCC4lbEPvVSBG7DClamWvI2nz2r
Ejya1mPKGt39hKaxF9Qlkr53AZ5PX/OWw/VDUSemTcAE/3X+sFNhIFUrbmGAA3lm
S6RzNmks7lCCswCIka71onDLTlLs4Dj+Mc1PJ8Dtlw3nqkrqQKTU+ukfHErPnDXO
BlJ78Ytm+MTtR5Gq+Z9IrtV137f/EwiOa2cuwK8LG3WDfUh7zfu8aD4DkVmKPEBR
FavkLfJtjM0xZ2mgTul4dh4mBNrXVIv4oo4NnazQhD9s+DfASkXNHKuJrg7a2tFB
S4wRi6AS3OADKsDSaxk5SV2zUMQk+38hoTnCrAsm4WA=
`protect END_PROTECTED
