`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wzQAs/in2TgOcJY+NSR6d9Z850Z1bqyb1rMXRWXMyKM
fyeL9UzXr2afX5vepwVUUf3WerbJafNWD2pjBryZF/p4btF0BFlPtEQln9Vs7qUp
c2jWJM9odtiht/5paSKOzYEn0P6wIadS0uEs18gAMO/ezyjD3kpZXP9K9CbINs2J
7Pgp6ZiJ5Ajx+smz/Ki0ebUt3IupDHcDTSstPlfGt7D4MdT5qWmWWqOrn+OQr0cZ
3t4JdDwSAEbRgqZTGRCyhOTE2y0mpi+BjnwOst1bDAnEX6pGYDSS6rTFZkHHniPf
01K7e4fPIzyOd5FoQmQ8h30z0G1TMwg/assrB5cnwLUTHO6HIheVOiTbSJ89Seuy
H2qIgUjnjlq4jq75iT4NCA==
`protect END_PROTECTED
