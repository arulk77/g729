`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aZFhmBc2F/bSrQkh1U1z049aHzwBectbV1qtfUU3/dbS
4vRsaDbObj9g8J92AciC6/D5fnicjry2NehWUhc8MGuNrssgb/vmG3zQVSuL7J52
BJ1753sLT2HPluCSJ7OGCyd6DJaQYDi92gQgaxLF1Yqj1u9cWYPe7LMvLriqhPQc
S8wS6oZc6FY9sxJOlsmPfw+gUdoXtC0+vzmmbSSnySkWhsCin6bqxjBcEJAzuD/r
n4Ww8vv+YTiYaG1vtcl/w/YdJg3UitJKmYONCT6Pfhf8WYCc9MRSGtkQ2fLQdv7r
cFidDL10E0AjuqQH0ZYL6KPh6j1L0WQxDAbQhC+R7b6mCc8Upk7S+mPv3EffTri0
m96cIHCR5rC7BtKEEHivnqizzSZTYKkeFGGe5DC6aCFHesfsyTDXLnNNB0PWozMb
auQa6dQgWQDYcrRjx73UdBA4rkvpT8xRtu7cXKj3NnvEoJ8uBeubwOX7wrXLGIIK
0Ee/ToxVYWdsZu4RLqzGD4b9pokGmzsT9eWyq9xaUbroTdo5paBAeCJn07ERJTW/
16hB31eIMgIhT/kQjlMIBvwZMG7BXiqifrI88mmOpVvTqw0EAX4WLNIlTuOVezLa
5DSxiukiR35zlG0Cc4ImXrJtZybXAZjmIH3zO5asA+IWCBZ2M4bC+S9fp/ID/tyB
tJknqpdgXg0RErzxJcBcWHqgtJbKMpAGzs3sqq84x6an9w1bUXZaGr/zE4Q9cxqz
DQQ7kkgmgX4/6gDjtWUk04WJxaRtPsUUnpWzLWY9XCpim2LiIrRS/CGqBmYvOc1g
oKJzTXdzbqdhtpGW+h5dLvVYQcl4eyZ3teVVmv1wTXftTvIWG5A7/YYHsbokS7QE
sHkvpBeKejb3KVAP1GpG6vfydczMhuxl1o6zRyVOU9k3na/YdKzv7G5lh7VLTU0k
TIYDy3fyM5AOCKMdA5TQmaHFwuGZeF8CQtjk51O6pURtIGugYUgpjMnE6budperu
ppcHAuAhtHMcRR22sK3Ke5t9jXuo1u2eYAUQ33vKQwyT00iwdCxKq6jEnwY2YQ8A
CbwT57VV4YBun3dlRQ40rUMWWmdNihOh2OjKvsOdXbswhXFvwyq/0Xv+3+RSV+Xn
eFgIL+MD+D3vOqFrUKmJkXiXeWn4s1myfqgNP78vo5+XlwiK1pODz0R2/8IKRChH
vBgKXw9nGo8cYlGVa1rUfwYpQyAi3ResoFHCRBLWK/0vtUM1D701eropcfjrC8Q1
JyM8lvsHHKuEiNnJFCMORXxDKsW1f9tUndScmQB3jW8K3L0P1TWdk1uMrVSGVAp7
oo35na8aVBrsZ6DnQNA/SdiPcnjcGCuzB9aOEBTFEcB+uTPJl9rz/jf6pj5rvEQp
IH025G0heFZLySZ+YX6HVJmS0fXzcrqMsb0NWKjt/hW2HhOVwTJA0YsVIKEy6hpz
uMpZQBYT8g1wGpxF+3Zp7D7VOVPJ7iAnkXZ06Qsy95sK/hnTR/jvrE2oWYY/CMah
0i/ja3MAs4/HKB4ZnIfEuXv4W1M4bXwCggnX8xaeylvEAZWKfScAsaRb7ClaYZ6p
fgbJ6yvi5cFAfLBSaIma8PC45QcVupmtMx6bTPYTT5vA5pZUitTlLIGWKkX7VlSa
t0RymCIcWUfiycu3+cJ8WHlbTvZHJSZ0c0QZAfE3+puLe1qiKehceDT8L6M9zY7F
Iwy0DZUFQ1BcpwbGhL96SwCXynGmlvJOpgSOLSDtatIDjp869mACbGjWeUhF55Vm
hs8fnq7DcavDtDUpWTGRXrFyfkMQrPrI/axF0iYrmaUMnlSdm/HQXxDfRZSUU4dH
SSEGUI7K0UzNaNXLWof94oDxm6HMmmeD/qk8fwLU6KQY9PPNf43ATJf4/arXLDKI
49ADNKpgg07f4tA2CB0rzyw6PwIe9YntxRvdOKi+HZlKSAdF+ZuY8KTonEcJIu2k
oqjWt6dffBS3/POGyySVdXZ+vEhDYOkNZfj6V80tGY65o+gBk3SteGPdcIrAgdSb
31srHeSCfdtiXZw9GumHsTREx5EES2a6pW0GDmbef71KjL2kEp45DU7Fg0F44pCA
MBCDerKD9rWFeGvBqlFpR8V+IHkAE8TxDU20EJD4IZkVQV0Qg03JBP79tTbjhivy
4djcsriAcIwwDHe0UeADewLIC/b40Plz/KEovLwFcN4TCtPGuZ3gt6jKd6jMmlCY
31FC8jOajrIVyctJU9X31d4tRmp/cHVwltIoN3UEPiTdVCEmIq5Yr+97Kj9RBH5M
ZvVDsBPe4CxqMiyE5vlDIOELPX/VBgBxijzK6BA7EuLBNRVnbRD4xRLj5f8qx3og
91iLZkbRXKaHyeF0DIpZWiZwokHO8xa5PX36g2YrGA5g9FqudjHrU1bkR1sKwDlJ
LHRtEdxalgYdKQvhofQ+L5vo20mwYvkpBxvyLgsruTDhaGhtvBUj4ZcxHg9JZ6z7
xvtqRd7hZ37V+AcSlx+FhlhTjKe/hCAJsxgyCC+muG8sJ5KMhnMTqDXqd4osI9qJ
gAbCxecesvX+LzjU7ZFjSmzA7OLEwaAW97V5qeaL7gJ2nmiUeDvPMvmVEq5TlOTp
DQ/VnvWB/hNi2T0gYi2nwqjfz/pKydV/28CW1FQ7p06FPqKsYI6nBYRgka+8MG9O
iDUdSYeD7IIxasy36m0UogqZpKn0L431CqKmc6vP8w2THOWJ7//ZNCxHfwnCtnyg
NxMm55rJ91RkCk9TrFf5ac07Q6eGakadf7E4u9k+ptHJHJ/OF2qjEUGrfwRYHeh8
qiWzw6qMAF/AA5ZHis/36Xscj3C8msMjSriHo0Zy88vW2WVuKvLdgVB9kmteE4+r
TxEKIxiFTFnfZdxoE3KnJXucEfH/+NfNVmD6T8KdeWT6uAkV1wUhc9OQXD3kC1lg
RCzz959DcTOwyV29vlrNYfsL8FiJnajDD3VWWNtOCPiCPGU20KZUSpb+0N6c+EFI
N2VfOb4OY5Mk3pyfnh3EUdgCA5MgsLrnLCqu77gooD2OvXmbe/mCZyHoIRaRLj15
xzRTZdvqcGtT+B8TmJ/iTZY69ZIfet8xziTfXbxbucDSx7i7SDIQI4yO2BQPmM2J
Hyqs8tII+RZ3QHN1f7jrN6ts8PSTYGStu7d1bAaGiuE2pGg4z+H9j8bYE7b9SMFv
3y8tm2TiRmEUThHakXaggcDoCYpH8dTneVNIq4xDlps0Asa8KRtVimeQ8Y2B1yEJ
21fV6P/omf7/NzwtmiYzfOC0eFup/Hc/L7h0MCopkhno5ysQ/Urgq96apOXwnvD4
ZJpIuvLsLbtd7YIpyfJ1STrwiMxcH19x52rCGEdvCyCDnPQpzqDoQJe7aIvr/GKC
9mRHbPIbsmw1VywGmJNncE8XTLyY3VK8sIm9VJQ97Qe50NumLHkPhVPhP0YISiNx
s7WMwsuVUgDZ1FNEZMfjvFUfSzbSu2/U8jgmsajHG8E9A3uWJJQlAbwDQTHBqIiV
Q4VScDpj9qPLbOAov836xvFk9EjyHRtQ4Wz9ENfEuLtYQiTHQHGxyxmGOyPSU6EC
4tzKQNCdw60kNSxeL6sxQXXzS5pLZZbhSObYgX0Vgsh9DEka8UQVA1phw4dKzgnW
2UZWNSwNuA5JGG6Akbvuo2nrztaxPgnRyKN7fLRS2I5MhMqHUVUgMuROLYVv0+V9
nIppyXtvjyhkGkEIxW0upn6fJIT/CTE8aLXh3Hb5b/TkrLYaXd8E+D3rNUTQaIz+
PIbIWr89B445whTUbM27sTlfPaMp7TyirXp6PMPEyOHNivcjdG/1lVDVYx8jByf+
DRGgMq1+Tth7lZk5pIZb2WDpnE5DcFfVY5BOCzxUduEcipnYmsBR62CV+/HTW7Xv
YSMESvOKVlV2poKAjr1BSITpI1QwUtbCKwPT/5Mk+A+SM6+/9MHeQDo4yMw2ZkyH
tjPfXYxSxTL15m00waT5T85isaef9fcz9O1jW5Fz7L6dWtq2Naqg/T4/5kJ4XGdq
MCBlUN8WTxjZTtO0cq21He0cK5v+FUtKbfatLhGxorTTOWPw0P56bf52jQ1TkAVL
2ylz/ZIvSHcUsNd9UHbrMdbcK9fNyiDaAmQDNl/7n+eFYuRpeQ0+1x/yAWccL6zi
J6RmvceO2n2mXXaOlYCDPfCI/gc+aXKibw0VxaobCNZ31tSHItQtwWYUAkVR/rzB
LUIYloZzvFs8odRWTywdm33dtya4eXy5ScF3EoqOukguhyIPryiCwx4xuTRb03eJ
nD4D3JfBij0BnnOPvaJ7S7K5Ilz9VAxwiNkHCwaDRQgBu8y3s5XwToY4P5uCHkHk
oz34ZgPO9Xy5+aS3QIfEZOZqFgniJrJFvSa3006bV29kE06pvY9UM8mHGdERdPS2
Kc9Z8z23/LCuleST7RQeEUWkM9xtYNytauriyD49CT/TfWvKGrYhpihcr3+QOy0N
8yU2JgSpxNrQ66aLs6sGiTDu1tilFpg20iYU1kDnyP3NmXWGYSY4LRM/Ngmj9dZS
tF37F8mWo3l3K+KR50OW98S+QY3yR1O/dztX/cJnRj9o220FYqRYz9WeNYzdpI6R
+aK7kMaDBUVIaWEOfF8DY9iNwKYg60W8AOpflQmMeF9GsUW/JoYdcndtrxkpR+Ya
ypSl3Bx+PUsv3OWKHT963rsd7ZA2CdI9LZ1eQxVq4W/hcuQJtz1MeCf5JQlZC72Q
xYq7Hr+dPBEsUhpYYjd63V6YMzI2+KW4lLMObFZED8AlISZWQs+SWLWhXGikS8sR
WIntZ//TsVRrRfmws6Bh8gOTGteTyDPccR40X1E/oWQhLKahYtn0Ue6VFgTMpxJN
is9kwrolKEsqmxDBGWsODDLigPG3kaC9268t09ikUK3zcg3khVKsSy7U839Lfgpm
9L8hDJBdhpVQmSFadUlNfGxBcgSnFJ3A5UwkAWmvP9BTrwuIPYgfqU0V1nJKdc+U
aHBjlfH1brASw0045/6ysOJ6qUaF2jfTxMKKU590mMq+u0zCAvxuK7C587gXBeSt
ZwGKDmSEXF6cWruCutZM5FVDby06zQp/L6JIWhyjVnrc8E43mWnEa50V+fY6Y5Nz
gadhsarOGwrFMXfQ0UtNpUD2noWUpoAvSnB4qYLALdvdOEcGRK1BdurGwe7oAR+7
+I5wdvCn7Hg9dR4+5e66emtebLKVOflN3qDPU3tU8hcDr8N6cTlUD15Kcqh3Vwu4
IHLOpUecPemolf7LMwgaKJbC5nL3wjP+bhjkWoa9gre1UyE/gcjpTlHhHV3ZLQ7G
2TqIZ4HqsLX2aeQl3elE+kCHdiY+6s8EgFdxsRjCuL4zwmP20mSvjz4dXqtrv8ug
OC9jEgmiZJpMt7c/38I2bKS5X0yqBxdPJp4M3yM3gIXdsmA40mKftjOeESJ4m7jX
L13O9/bv3S0f32D/bMTDFcejfyW8iE3pwJ9SAsZcWqY19cAqTXi4XA0AoDM0NhBk
I+vxRvvC5GNp1xwy7heTXSKyP7OiauJjJljfT3/Jnc+RHNb6GMLREedmccunMSqZ
u5db368Nfg38671m9AWl4CJLwRg9adP9jPx8yLOg8Fvv+oW59xLfUjOPgTajdFI4
vUJXbH6E8Dqe62J4EbQCAUBNPHICQYRu0Fq0zdK4vwLDhPEJBXvIWbtaLVUlgeM+
gQ7qtwFUPZS9rhF+gWg5bs0RTsugqJOFOK7yla1+iHtWUeH2pgmpKC/qnsReVJp+
585iM0FsjxvzWw7p3jbu0OQ5C4YJXy5QbUYk/mFjxTNBRKbhc5pD6GlUWAaeWcjb
lSybeY6fK9KVFlgH9nUzRWmBcdJRNrY9xK5mZDxKH2NpoBUImQ3ElfAt7vv1zYSE
AyOWf1s3tj5h+LIGePFKmrRuKPP9/N9gv/yV3G552lfhz2q+i52AzFC9Azlu24nN
QHSD6ksImbCT5kZzdyZbmFyAVoED5ZRNHV1kw/sgvJBpmtc6hRjWkvBZNNx+1gCg
1b0KrW6/KUOYrnVQy5dDsBFhY6MfM+6YEBqYrzwrHhUsILxxr2L6byrM8oESYH1a
wEeLWGSZ/IWxpF5xRdnLEuP13XW1E0w2C9fMCWNJXQxhNNlrj+RrZAldcyhBOEgT
OVjnm4rkQETDBZwikI8vHcEQY1k8Ez4ZQUhRiN6Ip2+tdySiq/RMZH/Yst2FFJsS
6SKMvO2nCd7xNjB6qPN9wpxga8hifMd5e75po3IbKx9dTX6Fn58JpsnAqQK7KQgC
4U84Ajgkf+un5jc/eeknUIAxyiiEVaoVtVqWs746O0UhGp1DkQiCnYpeqfqjolRQ
TU1ymmE2bo4B8pUMJfs6KATkLazU9A6OvDnsShUjX0CKNUNU+oDbjsIsoBKKh1a+
fTGwcPip/NqJcQWs5pHGcsAyTVlHa15U+5yAyBO92i1GFzenLlfcVWyzlcMXJo1n
6BKM0BneP35ZHQ2eQVcrQsBIevlvnlt+jXUXQYqnOmLagDt7g6GnpE0182nAKpEz
vxqxaH+JWdkx1wGqsXXIqO0Z/xeWPRNcsP9bME7YkCGtfm1H4626Lq1gaRkVmImQ
HsZ/F4wy9v3CHtkTDJJlc1VjOEEiXRcMrFzeVu5SADhjC0is7h8kYDDDgRdJ2xu6
nb8Wx+I0c+sVujGr5wnbSyPkKbAFCEluX0fezIMuHAc5jzXBKH4LAIAgs5a0hzeN
PIk7/OXZlnTiLqcuNdQV++kN0Qy7FldT0VFY53RYI2B4oWkB9vOljunU866OTuM8
jdpigfMk+NdtcCos/SYmRcTJwmM2dAyZtwl0vVjelv56EOTfzeMq2Ox37Ek82cYZ
SdRJ6UchVQDwOrKFfdMeeGG77DOOg0wvcZPLihoYl7JJvcpsktlpd0FIWVlrQmCE
QQoqPt4l6bJjn5IN+783EueyjON08P/ujTfQJBatIQZT1ny9kF22EiSwdsJs823s
Xp3QFdVZPElEsP+dPIpDPEBl1pYQhuvlj7b/s7FzBqXKKA12EHAz9zdFyFjEb38X
5zvcuVQpomcLL7r1975wh/Fk9fTaM6MsN/A6d4yqdKRdojQzc4kbS3FuIDzlBWIx
CWD2pzvpAvlbPD5vknWqV6owCkTjf3GNbBKZ6NC3mh3Teri4qUwaRCBAfFUka62h
RY9gfLjGWRBaCMmHS8abr/kBE02awgMo4WNI0VP2rmMeReBYKKHk+PCxHEir2ixX
aGcgCGb23mIhV2TkiKwUrLD3Kfh/GizC5stY+4JnwBPxQvXTjCsdbCnaiMbNnMHl
xk4N/vjVPH5gxRbZg86hIlIwIzRkwtcLXYgFyd45EPEE8NNXyetLfAq6Nj9McItu
tfm2xyTQ1x13DU4UX86O/6JoYE3IoC9auHwozSZQFumUnDWDjU0xn0M0MPUEJTaL
S7Ip694Iuc6Z2brC9cSD+2aMx04vnaASDBuZ+WYGy7qnvyKi/OAaZ/QB0idL3lfH
uARrpgpbBXZRENQGxL49YjG5nTPyp1WzjNpAiF2UbwBZtzEdB/tiDDKBb2IG/pjr
VZzq2CZzqh4/wIuGlzFNjuQZ8tGrvmtbmvCEDv3tdDPO4m2Wheb6KHqHeY+Tg21N
PbH3KWEvYtI8xoBq4rEqnvKquqCHZpoVdS1jbC9yr/Iu1HofBkC43zddH9lA4Mkm
27adU8F/Rv51t6xkqkkLuUDMtte2hfPGTb0viYNSD9kBw+W1jsSUy1ZGQL8ba797
UCSMEMUbbFKSRbAbZ2qo2yzRJQSZObm0HUPghMwIhBMWKmFwBeBYVAe2FGC1Wojn
ZTNqF/ZdT7fBr7QWBgKBJA==
`protect END_PROTECTED
