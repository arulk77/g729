`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGBP0MktkoTNQJGPcilTSBuYT+LSr+oXroDPxZqYCsc1
+QnbuAUFGbj55t0sC464yMqWSH5iUoHlL77A8+bFK3TWe9X/VAk3dRPOhTrjCBUj
l5ehkJpyATsbJy/LPEIQ8VPklTIlvGmfo/fGwCPV/PyuFRHi0C66ckjwZGfNhJWq
`protect END_PROTECTED
