`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
h/qQTAaMOYyjha08xDqnrymF1/xT8+adVrkuEHZ+1JC3ZG0qk0cUoIOliTPaaaJx
I22QXu6fjiQ9pbH+3ebynMCUyq57iVjos6UTgGJP/9Ka9Ezxhios4WwYFn50VCum
JxYtLnaxJL3LBM1YDNurerMf/zH1+G4uAj5fh1spNLEJ5p3DTSB/Pev59LB9YWDt
pZWPMgtT9Eb4dnlkvdsXLjngkD1Lk1IHpNTHoz4i12QHn5UahmEYeweCJeq6ivPH
cm7PadkR09+Ph/M+ck3tsCSDMluchi20vQpGdt/yzQ0DWw9vzvqNnrnSVJGUzCrD
lqr/hVYLui+q73hjCt6cxmCJ5JJGJY8o/dMIzTuXdH0EgR1rHmL/bylf2GfLuM1L
fcFO5J9r/mSmKiWa9WRTCOCCIqx6P9gBt+YlyVDotp7pm6brn+lFy9ZJr8UtHCgm
mlzwmN9C5XW0C1j9KzMWjURS1LC7snOu1w4ayQbt4om+UiwpiLuR7yUtJI3pFPFJ
mcSuCy7L2nL5tmj7YIlVkgYh4D0NY9QsOUEJX4gOmx0jiAloFhXGrZ4bvxWq/gqK
aQMSoFCf8nH4d7soGz35VfP04W3ptanx116cP+uEevyJfsCnhorg5hn407yppkg3
`protect END_PROTECTED
