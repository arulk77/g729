`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1ab+KgortBga6r1WXzxR9wvU7HShHUV9zE2/eKx4rFzzL
5gy0BM/6WOHkikgCiuGV1Yqhw1IJwdW+Dc7zBHvpOgWSDaE9EETAi9xaYfXVC7Qj
Y9GIyTq85ukH/924WzKSsU2XiOVK2EnnvgbNbz9KzHAMGfdfNOHrgf8++Krn5p65
Xl/LEHmcHM3CA+Imy8EuGWIkRsBUNma4ZYKfdI8vShVUBpg2of2L90E19lMtvhTb
veE/Uk/SHgnHlcMJFTNU3gmod/kuGYeYz8xOEQsncLPSdgCZTnjNaLCxNx3/Z9JW
VdKhb4TEumeKfU94ezk4bJzDQd65OLjA9pxb/TQrPf3LtNK0WptpLgwjnClR13hG
uyBC2dDeVDJNzKnoRRclEoBn+jh7kBy+Egtxgf/THKof7BW6nnlBhAN7lrdp3dct
8BfFT9rUBDnC59VlC3+yjsW9h+ok8LfpCutim3wfKB5WxOl0pBrWs05hVGRHHR/0
7rqKcBB+WqoOvSUB+4BGOwkIuUnY673AawtVICYRoNc+9SUoP6nKCaIFTnPvIHps
ICz0DA7o5UPFqUYFodbgGh83x5xpN5WgZpbytH7fzK52p5tgSh3cE3v2FjnhER0B
JdCXjwIROLBMYc+thiVBUmD8EfDjoupYyxYZbBgysT0rZM39kfy+dzizzw930EK0
Ms9XsmMdhbTqQ7c8d1sgg9tNayVwkImm6FqA8ZlSaM4zTF6mDa9iPrz9pQJvHJf1
sS/tFH6piX3ftaTudenrysblA5Wu20ObIrBqhJZebFIXfKvErWFx/KMcSGJdboR9
h0PMmiQuYCXyD0ypdrtMQ6qmlNcs450qr3BwkEMAn/N5irSsQP0cIxR/rNE++SKw
ksrtCxSE7egiAxsIgBICu1RVfrPX2VJZugZTl3lcLCzitkTeEjGhOdrEFgLxAvgS
sSz1hLlXX44kCISg5rN2T0rAns4GwQ4h1fUIQ97+fgc0kpLGB1i+akwmWSC89lUB
jaJEi3Yrd6Mp6balvT4NmgHdTa2CD7JoAJQPrEyxYCwNooQBrsx6VVjNuxsSKpxC
0k6LAsC6o/KdmxHW1gjPGXYFT8hb5GMskZoRU0gwqJaISui3emal7qAIJ+xMRSO6
lvCLHfLNvu+dheSgRLqIyQfsJQa0rVBXHVRf3goUahwpxrwY+X3AV+CI8LZMAXjL
y2Yc8DesH3+q5rDjqk7Z6cZ+xUn4s5Wj35qmdxew5Q71+eUV/MbuTETYsAaWgApq
x0vNUYzCy3JnK0D2bgn47k4HhueWi49ykB9RXr39cjV3/bFV1XFKM4siE7vqJzXQ
UMKfkuJqOkehMRv5GGXjDf1wjO3z6a9LIWjloZpxEjIs37sWdz73sW2RfRBxHBky
ObQhbaSaIS+EBUAzEQUmhdUJq9EMMu3uA6zApg8ZH+PSS/JLUDU5N+gUE/5m9RCz
PFDwTtE8e80nwjnggPSORcmgL58bTzhGcmvO1kIgmhuaMQAWg45P7weC6ImGlEtq
2pJm39bZGeMw9w5ELv0T+WQTvVYOwVXY1fL6pAWe2JDPdXfghJ7O07hRA0SiXkQr
wWEh5WfwJCESnjKg+701NGjLibsHjEGJL2/Ngo4T3v6RCtn8rTr7u8A+XbTSLf8Z
siRtmUq/9KRvWMKQx54/rdthFhE+Z0Z9mPKAxzNc3BhKic9n2m4LzfDD2IbBT8z3
NjZCZ3j/VcUKRN02e/0N9wPV7XMlKTwYL1JM1zZ5WfPj04oQKSM6R2nEj74kSjaF
mJjmxGIVgRYdCd35rEiPLliBrJxZc0fZ3zjjYgqVeuMEMs/WMtZ9SrdJcxy6CZlu
K8oNjpB0eKt8fKp2LqnyvXhTMFBf/qoUydtZehhuHK8El6sQBHWSWig8NMndW2tx
J7PGHn/NeW9FaUB5X4fQxYRsP19H70agYpaCen416aLG5KELC/ACvT1WPbQzg/yu
2p4ziYhrLh8r9omMepcv/D/tIq3hPpIlwktCge7pHDw9gq8m4nOfK82FeaAjzkAM
wK1AGLCKppjP36OiJcsuaRpjNlL0tMjO8ghgu6DRrM8caGUNdF7MQoq0CET1at/Y
v+kxK890lgxlLGywOoefXqnBQ607u+cWNyvQzVo+4ytld/UQle9GQ1ROghk6P6/y
aOxtOY6o/Dgdj1dO1bdHDWEk5uU+qAIW00wUJ0Ozu1XCenw3bHrlq7JCp02LH4Kv
MLP6k6ufgfHC6Fw8ivyeVmOTzBEFotOnzLRpd+V1l4ZV2pYZjUYVCOtlfTK1B1sz
JWUGuq0VtY/5hqoSEA2/B9N4ZghguKPfVmXUyh395uiknDI9h4ZnymxRS0eNmBk+
S9WaCs6R691FmsghOGXFg326Ne0NgNS8ZievthMShXz7drIay4iuSK/hczeupEBd
x2t/UUyMtAQO0L0SFA0OK1QvH4CrQ0WcSWPH1feCmw8Sdbi9hIzNTdujj2ecvMiN
ICxuWEgbwJTsagByHtdTsCdyP5rJE5zrO6GSCKiXLo75fytDwif6ZY1HD+JzdukT
wZSyAOkSzq5/EWSjrZmJlo7jw0CULsbQL0b+HjBF77vPqzTFJkFSA+2RlBW91DSv
XQ80/fc5f8Zi0FQ+zGoHMPBXnQaY8oSufVO3fNzdxJ20VMt602Xkqx7gS+usOl79
v1dbrNkfArxe0UifX7m5bJoXGH8nnkVpORkIx+ueBqBice5VNVY6CCl33nN78bpR
YLRihg9iST+DKu27dd8QG1SAK/GOgXj+yJrrd04F/TRHjPo9+3eWfleGcqQMLbVO
bLHBib8F1mDbe3d9waLoqO2UMlg3+HzRqf/NnW1wiUzozrRZcb3stzx2ujcSSrr/
IVeEFVosartT2LHhw2DkxLDXNYo6T4t21xeldPhD7ET5XypsKLeeHJ+M4yLLp8ah
nIFgUIQQm6inZ/uU+Yp0pmuM/lNE76N4kgWDMFp4f96dWGPpKCqdvTAYXu5AqCWv
gXX4nX9Kk99JyE7kBytg6HCsfJMMNxlah70p7AjnemQDuxQMk6a11+6TOmryrI7U
5pBYbbw1ADdBr4TG3TAWFYLQpo65n0E3jvdYasYdJMnM4Yk/4g/MapT0ghG5KDv1
dsuPKQxb3AZkMhIYIGbl8Bji3S+y/TfpVEGD7zm+uqlJDC3u2U/UHRz5WExPZkRo
MOyZLzLFgB8PIlNxfJ0o3xHgqn7Zguxi3SPcFpMQTHop4lyhLNnraTCAjZ8hG2Fw
02yAumxW6ytxsyGtUdnMwgxdRl7Cls5Yy3rEZrkXztmkoUyMri8zSpvrJyykKXmB
hz/cFamvZ9i9/5Fn5s1lE9gfgH3SiiT+Sj6qq8A+bNwY02KO/qOCs6wY7QoysvKj
8DeiIgjG4b6QWSIHzKfG944Q5O2bQXSeGIQPgb0/aoEr6/nFg/QxeMQog61Exrbj
qNQnMs8cb1FdhmT6z4K8l05BGq4hyD83GFOttfM1ljtj+9076ImUUxC7DPsJm8nz
l05zbNKSwZ2VRj+OSGmeRRXr3LXMrJMlGYqPI9Ca5L+/CeBZBagCZnwAY1EbpGsI
2ueHLbsKK/T4qqJQ2YG/xWdU5Dao9iZ/bbNe/jh55Bn0HvtmUatXFPLrSCQitqDO
84rkUEdZfslf0o0exB2d3sQI2SBT1rlGgt3ndpksEe+1zyzjDND3gC1SNYe/9TGX
9OqLLs4cOea6SjwEraSeM8EfAiISBq8Bj4fc8hcpFfh293RYg0VxgxcEm1RcN0t+
dAeYxHdWlpUAG5jlUmLO1iRvUz7ICCJGcq0FJ1eeq830AAdXiPvQRQh6DEDIbTvR
QRoMFyiosCiyRperb/wTDyFQuNadiT4p34gAdqZo1qz0o+Ymd+doIHHtYVgF8u7y
TPNtujgp72EDI0SpEUJQE0yRnMM7Vx1ftEXUcPYaVNCMme1HD0BrE1hksJfjjwqE
FkIVU+JhxIqPsxQCk6ZSpBtuaCZuRHxc0KKa2qgMUjNuXiJH4g5hY0KPL7Rmt3lk
oVm6PGJ7RhZ7vFe+9UWgxQRsIfU4kTWSPxcZHBI429QSzO087RkGPJwIcRA7GVle
t30IYLkPwoIoDNNnTgU4xdQRFizCLSRxwxUAXcSlsVXHpahSO28nNPqa6F0Gc4Yk
6HC86hKgFKUUKOhNkiDNj7OFL5UCk1GsnRz3Sig2Ku0iLKA5j1Mc4AJW8ehChtTm
cTnzNIcb9Qk8NcQwHfqgvOw/1j3zQHiQlyuhH9DdsXlxhmXiWjGZhEJZI9gAGfhM
3PQ5CGeGUf810kr2k9me1LKUQBnksnXUetcvSJpDrdJhM22s2mMCQoRUr4tlGCf6
vx0Xcx8DWsgKbZStF9Z04DvAThGV4bKqZSb4/muuAVdiDebtIb63bWNPmJkNoFsR
3lYlkoBcJu54+l0bV6ltgmQ0irdJluXewAsmly4ax35Uvz+MMrfNOIECDyYwH+DK
0kqhdytqI/gGSDCgnQbWBGHJzUaw7SacL6IA2A/30DODJjR1wZAVyrLm5AorB6J7
NixF7NWh7U6zam/9m1F9FtdGyA5PhDN7453/zjteZYYQLjpGeIN0PCFwfUdjtDYA
YuBujRPYxNXxvFy9Ls+bTsKKKz61HDm/ZMedTXjdnjqC+PZdvW+Ghy0fsxghHhpU
k+yevUcFVBvjmgfi6ADi0iGVIHboI66yfMKMsfFEc1+Qu9wJL74JsxB2qgty+hQm
ekifTp9VOn46IMfUdtMB+St4XR80uu/feC1R6HYNYXJGrstKEAN5VRP34yEviFZr
GwUrC+zk+fqRsg3wsymPunR0GY3S1pjbJJ53PRpLFsEiipgwxUwf1fLTASqg9+3z
a4wuPXB/yiD/bk6uVDubLly94sJoKgPHgGJ6u5WjZZGPQl7y+NXyqfgH6BDi/6iP
DldSVSQoZoxR2/IMUeHYN6zP7KCOO9ukFyFft9WSV9TDUNOUhq09fTM2gzpmw7u7
Mqvwc6sKvLb2BAeiMaj4cAZzyh5FkvQiDP0iPiqS90PLb0wQtZRx6MNQLJtz+RsX
zROxAevnpic1NCgS+ymULVnPUfaQ4QAJSqz75eeC7ZVtFZRonZl+8JuYrVQqyOKO
9JRaNsyYbKEoape1l2QEo2Y443JaskH4e60jKX1lMHoorTru5hJhOuVJzdkeQK1p
3oQCEvGCZcrvjqkeJin8q7YWcH/Cpih3PLK23JVMmDHxF8xygQig9+xCWTvq+DSU
IakrI8YrHOwRFJbRF8pYH2f6M4kv5ZO70C+31o9qmgMZcfBomi2KcEGQUm5DSvma
KGF1bWeS4YXguqlhAOPMrMfW+lnrC7CWUpgOpMuKsS2NltvuHlfcmF79oCfl9fk6
yzN5iE/XTb2oXwNmWKMm7jtyT4zPixEchadvgOiaV3zofvUr13yCXpYPU30JbUb4
H2DnDn6SYnM2l3JjIM7kb7BIYsdjGeN1x2Y5xu5YvN7RY9hQ7yyzDRwLgxtQ2S11
jY41+MsgS+hJMkRaHZdDVbtwjnMcQ0pBbaSRIGGUEXmB8oIGQLvocL15Dv45rDhj
/nQQ8SHfpbhAA420poOfJtX/TwBI++DQ7Ac/MeL9u6Vxhk/+SkZV/L21u4aPLETD
HOrEkD3POliSRaovezCDkzyblWVVZjzbQtL8UDDRH99e2gW53v05g/scW0OvCELI
UrTW9kn1zR4JiEICxsXSv04b/HbBnWSzrmgZ4+x3WQ1zlhg94Jy6XmgsMoYY+tGh
MUMrakj9Y2NPmYhe4sVoKL0OTImg0FLIUEtHatR61SbDeS0v3TRJuiWb0Y+BXZML
u78CiQYEQVyvoaKdAqKC4A/JDt1+PGMtuJW5+RP4AvDC1k3kTQB7ZmFwSajyYxwv
BBDFEe9Nv9KIUV6n0bxIDRL8JKW6yj7ZHUEOzlzKHjPmEaiV9bwxFWhHOTYG1cwe
WdSUP4+GV9rAEihAn8w/SrCvPw0YAPQXHIg0SU3leQJ4jdGza6ncpqVJjea9EQjP
TtKLJbvf13Hd/jYWZSdgoafV0rlfPvOTVK3W2UNkkcxzjKcDSqz76x/uhe/KyeD0
eCQ9MThPEsyAvbxliOa5O1wzw6Y8qaHht/UW+oVdsweNVzfbm0pkUESuMEGUYxHH
aIVOT7uTXsvtNMMJQHQI1L+s1Q9GqI76+1QvGv1Hc8rE4LBh1L26axHJjj+CUra1
p9IHrQl/hEJ7K1CokWEch6LCodncj4Q7mbnlJ0fniTCkGmjb7Br551LnC+U4jCV6
4PiRf3b1KmiimL63bzlQQIoEwfXe1s2M7JC1gimHrdWe8gziQvXY/2u1lyx4nmL9
YReFqV0thHNyKDocWf8j86LgePu96NVZD3MJ0sbJPIDvQcwP2ZqsIhmHMzpETenx
AIN/wZtmyKdzXZz78OrB3mCsWVKZKTUmwtvUZBQY4+k8pdPVA6nCIwdL9qJjDHd/
fUljvcOHH2Nmcj6tUD16nfMwDphjJBG07NTSOXl8Z3I2eThWPLO7ORd9bNNwpCn2
WQ3XlGqbEQN1nCugQCbeIXrdGBhvAFlcPd5PfHVmQxZ9aChjtoKPo5WnWLb7e1Yn
JFxFcplEg69Lisdh7C8dBq5r4OKUYs5zvFsUcKi4YuGBQVF6TTdmHS0MckX0ESrR
iTErHBSe0TbDerYGpZXB+54CI381f+IZBG1h/e8CjwrVbt6yUnZ/86xUKzEJUXAF
cndr+mrKRUIFrDUdkgI/va2i8qcqHHXGBwEgJzH44valYcMccNCa29oEb6Dg7ZaS
fsXZZo8aS91gKUp0X+QURG30uqdK4FFIGnTH/10rQaTSRv7P74Ow9NlQivkrC0kj
3MfRusxxT3PVB/z9bi8pQ9n+qp921sRJvexiGJen4ibsRa4l2So0MWqIdNO24ynx
wGD9FmBk3vDv1gvpePkgzLLkjZjAZRwJTkrZYyGaIvd9t+erAbXIu7MUJubvi+51
C7OCo32KXwpZUoZccyKl88vsUO4cDx8m+gWJM0T6TQbgmUSMQkkJhxCWO5cVXeUg
q3+sGlChf8rdq2PmwItvKyH+DxRRW1DNLkj+lMBGGbMv7m+qagTDui7gVi1DnEQY
YqAltwaDdK1+kPG7PJJlBYcDzWoS59uRkMZH/j4FamVHJFRmFmcD2T25ZQgYlPyn
tTTRs4kQluplu3LiZTPtcqSoPPYo+iDBdEq1VYk4yIMf5h3WU2OaqEmk2GPqOzFE
J4ZQk/VJkayBM0zL7+K/V9eTVXm+PvXkVFf6N66xsu37zGe0pQUQvRT9LPoyu6Rm
hdC+QjkyxjlQu1iK4UV8H95ghSP63onYSFH7HXhpiIiXxN73zarVU8eUpS6ChJoO
HAdsfe0RxoNaLNvxd50C0jIpTtjOCpcn3oUAUZ9quny+yuc+xWvfOJRtMGhAGEbz
By7oFh66v6dsRBaow67opn58Bp33Rr7RJyavjlC8tr4U9K3T3+bpxv8sYxBXb1iS
HDT+SzPB/bkpCXSX9B06A6QAD5aojFqq+ZU57Ps6yx+PrCZMvA7jFu6DdL5lL3vN
1lcmiCEpkx/Iebte31aT/Tatk11ZHUMsBP/97rja8HuSAxyLl3Rbk556mruQwEyE
b34s4y2OlumvcP+tFEF+Xq7fS44aHQ0y7Imw7Radr3CKy0OXTf8DDt7WXBNkmx/1
RM2PA86Z3JwUbuimM2YfXiw98R+x3wAcT7wX+6rxDN7epTgSO8IweiNrFdZUQmHP
Ku6drDc+bClliG40LilTr+4tkHQSUgtvtEWjpKsSCT7amBu83aVIUQdxBxsWUk2e
4dPGzgZIgQUGEFY1zNJesehSaYya4aw0spUSHt081ubvjumMmmWI9KCFGr/PhBBR
m3axJLHEyh9QVrpZvVrCke1AaJlP50aPLSYeluYoJiRclRJ/3xUxTcQoRXqWsLpf
tMGfCXbnc7mHgtca5lYJSDCdVMZW2TytA+ct55FqBDs7Nc7TnpfjxKEI02vgD8yJ
xXyFkeCZ/ygWdH1xcPziGVgbCjvIRwkZzhShy38OZTtb2Qrb3LJmSIVjNDbqhMA+
byaGjKK4Pj7pSTN4uXVsjSP4/PZfFPOR+S+j442Xr480LvfGSJaUm95+Lw5DztH8
fFX+QsPqSPnL2ebRDsOYlYUHfiPVuJeeO5iZLjSS8HswdGLN6IuejdrLimgP82lw
IB8GPM+JtGr+SzbL2bjZEX/DUegARYdk8+wJEpZVf9bpbmJDOyM4AKgvB9icBcAK
kzoBev4LXBGKvifUAJ0arO8Cv1/DGpxPAGzX28ug3lY6QbAtTvAAfP07VuWZeAFz
+3FO03jv2gxdnmOGzQrTI1QM9c5zcU0N2T1roXj8WZrEMIc+UGNzZ8Qo1BvAa+lP
y5/D6Dh84UkKhfT44/xK6lE76Xo1Qi7bkgptfYhvItvWDOLmkN5xJpWdIAtzKqM+
CyVNgGi2GQ5jK1GOoGqL40RwkTxcPCP2nsBK2bylJtCPTrrW17pSKx09YYwF0iB1
CQqA3eWRptO5IzNg+Cm9WvOt+hWQ40Vl7u7kEXMxjnB1dcNWOrUtyk3jHokI5zUo
9Z1kzn+EZprV7KQnTzaTeBrVRWE3sFpPpRYmywMEGWh7e9t13+k+775dxj39AHrC
Z6Gteb8ZqJwMdSJ+qwwJUo8mwxcBw5Dp5OAG0V0JhUuBoZ05dSW5Y/h+mrgQlzPo
MlBC1L9maFjVcGwSglThcwyzIL+YRWEhU4uFtiI6ZvU=
`protect END_PROTECTED
