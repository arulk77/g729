`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN7119M0mTaQwRKogiQX89AdplDBe0D26ztiReY5ehWm0
yx+PIus+4s2CVTl0GM/79+ONXoWxBHEdIH2TKP+GdU413M9VBMcNB97nVg1Bd9eE
1mQpQyEvR/4j3j3lLN0Jo0OTHWwW6K+StVUfqxSqruOP9Ucejd/NV6nufp1rCuuN
3EvVYGSSN3oIqfCRAE2b0bMzTgeHbUPuA/fnVVlsll14y+x3LUPeqMOKOTeRja8S
hqgxmF5WfdVYfaMohYyRdnzhplAXHSqP5Bi7Kp7T7HymtfPxLl0XVZeUcxljBhkM
0goToSlJyCCCPM4lNTCqBGCMOdugtXJOAAZPVRPTudBpSSC2Y32PTkzY3DfsCSZS
QkAr66MQ5fm9J/uOm57CID3A50w9VAp4CeuadYkyhd2Dhu88EI5WDF1AtAqHH64c
qA7084jQCLqd0996D/tBsSRcPIpFIBx+qnGrSWc2aqtryWYZ2/Xt14mEUNaqO+6c
Cm62bOCGH8nUW+L4f9zsy27DY/6Fx93KMJWYMlicLZ4AlO0F6RyftqRuQ5kbxYVC
zuNEEfV1iMqmgXn4M6PshzMTVf0G+PrW0MAi+0Y1JP+74tFxJFjknK9JXYpIV5GE
I0WAWbEtfSdZKOS7lVhqTa60eSwTfqu1ARUUAvxk4QggQCXdTQ8+Q+CmPzbCoN21
IbVV9WGD+HHEIiOEtRdKSzFmmg4U3Fuj7d/1Guy3OUOjqe0vsDVeawXV/6zFEENX
2t9Pf17L5nmslk2WuRtFkS5jGok/MF7EW1yA79XAqtuDaRFNety5qq6QbAOHSRSL
PVvW7uSRDAzmABPDvu04QqpqAAk7kArZil2yDyNFprQwIztVYrCdZMYAEZdWq9eN
Ju3sDaEBpvBkdBNHJwUE8lLRnx3nIa9vgyM3g8+JUWmp6qrZGzIaksLe9Ti8SzCd
96tNTKbGd2xYePeSVHAti5VDZ6VdZz08IrnCTgA5A2V3eN1muguGyjPNSJ8dMw/a
C64IQAENE0n2EJN7tQAv/tmwyhG79Z57cDgGSWas4N+tPAfWJ4tOrq1Ym4mXEz7w
Bhi5x6jEpZBQ1V7WqN/gtfs1wKBHTLKECAV8/JIKsS4pHKK2dm6vQypBXJ57vZqo
9EBBK/ph1CZvwwPQmgg54tsp1XhgJ1t5nWnbsDW6yHMPNnbCjaTZB+Nt5l+8Gz+P
R9O01azvmHVQeKpSZ9fhyuQxsVeQQD6OLKL8NQvMOS3YZSt9G5LFaRrRsNIsKQ0+
ukDuo7JiZ6l6sb3Jfu+gyYdXTqG7tdEh2RdckKZkk/JucCe0o4GW9hs06A9wSus3
7qlo4y0mpjIMwzq8rCG60Bgpul0LaIozMFszxBD5dcKBsn4cT/CI7mGY4U+6S5wp
xx2IYLqXYm/4AGbFI1ofeqxD/QlVIfjN78cJbubE/0JmYw15DlyetzM38aV3o7Va
ap3p1nexv6L5DE0/4xDnTve9uCQY5u/OPCJBu8R7dI6tR3JVGCpbBNc480F+r8Xn
+CSkIGFC9NoCaS+JDIr58VoHSdE5D7INCBDX4DDRbrY08mWY6SUiQOXwBxQ6wAP6
R9odg0GxmkVdhfBDzA1NA3nMT+cr/nMDmkT5Y13QmYHhiut8fz9zdTZezVgyQOAi
pQ2/t3WabCNtQY0FTGwGDYB7vB4AUIlsLPpDABwipR9yrCYj1Jz3iHGW+rIk4zDG
HnwLzO4OWx+qtnvPmjTwu1K67viEsqnzkfAYoZwWBJQ/Cosk1nzklLTUajwZEKXJ
T5VVJHjQ6kgUFcvXn9yvPvGBdRjzzUOqFGHfgY1iZfxUsWqak8I3wIGGLMDa9T5Z
ZFc2FsyO8YFICWQhWPHrQgbH75fjNw58Cq34dL1+r6BZJ2x/EuuV2VmDf8/H0oyd
OvRGSwMXlejHqpl6KeK69kCOQacfW6r75ra2LKsUAvQr94VtAUlLZ/8f7KNq+iQc
9Rp+38OyYdd042ZQQP3HiOk5vpfIV+tolHNaQpBWHyvNepnLf//Q1ZqQlpZ1fkd8
cHNrXmFtIslzxBEUaTv8AnolVLEQeQSMuOLMARTO1PCim5So2W2Vnuhb2PvCG+ir
hoIYLstf8bO+8aM1wLvCOnvn4jaHPcy28bkuCe2kwY8A6t7SrwoPak91fVudF/Ji
Se9tf4sr15FG9DsP0t5SjgviugGwarl41I90/shi3sog6uKS2BFfPMGgfmEN/bFu
Iz0g1CxZYbPZOly1/ApkMHr2qoqFP8cEU0Zywl7Z8xrM55UahE/ZUZT+rEXe8j/w
2L7p9UXmPgv2UXK1x4dRv98VIt4aOzRAg2YUPfwvtbSSV/joXXgj2prwIyrxsw8w
/jRabmQu/rMCUJn3zaDGUfZBZ+qp6k1KQ7UaQp+zfDivZKdHUV+A0JCke7a8iiIC
mMsXMCrVkUZmpj3EQyQuUrwjhD0qpfx+SSGlbCgcGv+KcbdmK52jRt1jw/nKlGgg
J1/xvyG/nJRRqqjLswo8ywIRmVZXc6anlT3qmVbqG6VK/CgLW984NtTIWl/V56Cq
F5bqem36iCDBtFfUFQaOhbMrJ5eCAH8wfXefttgfYzxDxDIu3atz50sNFxQe6gKs
B1iqcIe3UIWAneycNx0kTrKKvXWHOHomA92LQN70Wd1GWDFihnLy7F+7p738mNsy
O1RML7DzACfdIygGG9p5F2UCM11VME0a6hGlcGNHz+D+5FyKQlADu885q861ja3F
H5Ay+GU/zhTgxf4tcXjHFA9+uZfKRgQ9yaYzWUiVH7gBIIhiwesaGdF/vPMxr7cN
3u13zz6wuz7TwuXJLuNDR03btutC/S1GtSSkJMHo+X6oh/YaYwkMMb68y2+hNCkz
2VDg1MP2ADWyj9YyxVOKTr9EOS+284pykjBXbfVXwC+A8MlsMd8yutCcQk4Oa634
rnhZK/5FXxC1YyOf3VqNejO3mKNU+AGKFJpfecyaywl4HKkqH0gR1l+FQtR+7ExZ
XDbLV2lIOwWw6CsGTbz99U1gCcxO/5q8h/9n3fFnnaMNCKSGhiivlwZBMha66WUb
JQtNaPT5dKCrBwnWAJ+BIsV8YVtKttMlP8iF1KCrubO085noxIsTVAbCbzGkj70I
lncgFMAns6eYWfBU1pqdl/b3R8GdDPnYQz7UEEysrE82zfiFPG5wqSawvbUJjIsh
Fu2aZC/+/hqL6KSjkxDaXV78WjWrO3K3ncYzOF99kzClMDkN6j5TGtxcS9s1BYzW
hopJJe7O83AJB3vz1wK5RG8vJJKQ/l4nffILyaoCMl4nT0Wc2/DwFQUnbng+bLQv
m71+xctC3BqfpvmjYytEhIU7pVK/JUqoEJpA406vC2tite1Dow9nxv+9NmzH1Ndg
N6SHRbvVV+MJz9skTFtF0+IBevKhkxBq+nnaB3r8xR47I1+4kyRAA+6pPr3CJgpl
0kcy8kbiOq1RLwWuOP+nnYSM0uvGjYjx5FngcukARMdkHquRjNHTmEE+O6QjSqU7
6vEMWsfAGuABvqPxSi61AkbYSolnGcqthh8ImN+vzFr2iwVD2Sw8DHM+CRdf/FHG
sterP7xmCYnJuWV3Bz9CO5iqYJxGkKeFw671GXQA6d+KS5XHrtXxIYxxdcmhg6q1
gLtyJXuMyqhwuHQqoe+R6/ZdryWXVvUG8nJ7B7Hazv1jA6M0a8xtyd7YtiGXfpMl
XkEXzeDMWiGrMmSwcZVP6MuETQcclc4YlRCUuXFIkZAdZI/CePJjyeGVmRKhP/29
pUQyv/PqCAN+qWwgSCcY6wZxUrHcSUUz3DOXd4CsKHShRWDFOBkPAyVDJ42K4Wa8
VyaJwCN2kj8PbvfQmJw36uPtC05w9H+YEMku6tjgf/tWRt5ko7EzkedGS2jfl8U0
5PcG3rattoGhpDXNFSPjYDaB8UlRbKq8ludJ5pZGnPSVJc1Sm/+KT5V9FxoBTh4I
CmcY3OIJos3a8sk2ZnJ9iEGN1J88io2Asij7Ci2EbpGUPCJ+oEYcDa+SLmVD2sT0
zyuQ9LQlTMSVzz64Tl6xv4XQWQNIV3E/g/k6bfcq8xGni5VxHz0VAA7sSYMl3Zd3
XBgF7DbrlWm4H8uPNLABTlLnyRNXajllbtFEaX7GDccP/ScBXAWar8MipzQlAfCE
MWX0RBmtTM3Qg/XiYZWNS/dQ5GdCK9Of5do+44EuZciOquItjqpnM8bqyOBTZy39
QhlpgHrnfdGCmpZ1SNngy2K6MbvfIbvl9wYlICCrq9deR6G62UffO0KFqLW6ZZRp
gbiaEjg0rBqLs373gsuDJVrW8SFjrIBA3dFIWXdgKKnfnPp2bPGVDiGgPisxi7l3
Q78bZkXEcpW5ZXawxM5QD9hAV4CDRBP/hb44FMxWf9QoSjW/SrlkcLuuaCgE1yBl
nrlcLxYblR/SclkJ0lsg2nP0Buz88Cvnir3WcdC8cbX67CCNkQAufMeTNhsFVNDm
E/ra3jhqRMMpkx7YdqkRRD9DUNgNDfdvDrwqXhsGu5O+GatfEsQFuaZQX61S+TQL
CBCoV2ld/ZT3BqqaaSqbgWPkhfUECpL7q8fj0iXdcXmkF3/t+GupUdEe5QtWzZBl
Zl+/8u0CYpbPr1E734n3xFTxOnstI+q8hOxilSnPmhBCHEiRvx/8cOP8B2I0xMod
4wrFQFsxQVFMAW34/28zfCyATzdy0SjTMhq68yaSPk4ZCIfSU73F0q58RuUU6BQD
VUdjpv85P+UyhVVv9NWn8vZlJ4XAtAcrlx3vTS23aCsApne9kbuIRQIHQD0dQJEx
KX7AxtrAQ8sWP4GOx902fQnp/EyVCwhXB94Wd737hJoWbKA+J1TUtDmBkei+vVlP
rr1qskIVffEfijzFIssf5U2T/N2OdOnLGVN8lVmOL+nLcJufC7SMOl1Eyrfxl4yk
oq/k1V9gDLSXzTTNree+XXLDY3bFjnJkVIeQAwU2f4qG+vEYEV96gM00hPw4cPFW
I0KjSytnRsaX8MwouSk0IsIVmoAwiYlwUyPxuUNakYy6odScJUYzvhkToy9+X6u/
bm/73qSdpqWb9swXMNWH8hS4yICJFnawQtBOb/TfowfUQ+f+RadCIdFqZEIVzZnI
6BtyMpl7uuJIQR27k1bYtTyT0SolIstZdTDE1tRlhRmBdlciIt0AoCH2aERXPoad
kD0NmhV+P8tI4IWp1tdfOil0tdG01WhEkk6JZEVTl9rJzDx8mpc8adWbfhZY7Oyd
uoLCeiBv2ZADU64KhxebzP3w/pzloaD+wExzUhbcC441XkxLRwc8+dviAdTJKmBa
em2JunPYbNx+z3M1Ha+Gvl23nXZ3YD28a8Ee/aXEPaT1cdC5iG4muUmoTm9QV6I2
RrWvKwAfIDb/HFDIvIZ8m1BzAfQZw1MvAoOaKzSO2mbZnpeEPL76qMPb3Gcp9UuM
17ASFDmxb3J6QlPwKYx+ECFp0MIJxSaeJeKneMFPfCYU1OlU2E9YpOWyAYsG+4SD
lVk1qdKYXDqhSpe43RP4gqTsgTB4Mk/dqs3+NteVeOdTUlmfIihj73WOt4KBDhlG
dh8UKDoANtyBBWppTuuFCTHSxk7mTLal/kPcJ+jrVfS1apXh/ubvr6iPfJyGasFX
DnZXCyXZ3vgYQgog/C+1N5eoK+w5mhC8FpkRBiksCyLORBgFLJCZFzJCq4kJWxP3
gWXwdsGhUPHEeq/cShYWG5m5eVISeg1c1nbYMX65MwxRUqa5KBb5m8aNqymbDcvd
+uZhE8C0M6R3pHkoC4YpJLC3tbyBZGB8fTG+gquDStZ+H1sDeK6q6pfgIx4MaLGg
jWAfzAUlI4mNY7eonvGyqJr0VDb2ZCTkDCB4IDCpxmBdEFcinUf8Yv7toYjk18qZ
/dwfd96nX9zD+xsIYo3R9m9tr5omC4aQ/LtgU6TNZ+wkkAjxj6+RThAmZLHcZjNe
YVfkZSHihdaKzg9PzJ+HwDmQO3K4bAIQbxNW2JQci3T/0rMVmPgLVTHmSfS6RuBz
pWWfhMwGtDPtLS/ZupB2sj8T0YAj6aBrbSISCFyVVmvJAJVXwe+IdZZggo75+4gA
ZHg8jU3Orep8W1dhQaRkreEzZtll8porK+4bMxxZrkPwAhjx4QwcblCtIY+ZvfGY
RueRxDz140OGYvHKgwb847OkgTowaCvb/66ZlDxYZEicf9cYnHADOveY3mh/k66v
mdIFjae3ha7SgD6L/ZiTYQYmDttkvTxfUzN4D3DeAEv3e//WU5f1k5PjqCAX/gbz
eNAqfPCsWZRy6EM1QZB8d0T/3t+qhrQlg0mpRYQEfxaM/W4bmC0LT/1dS+06DmsL
lmrfWMNlvDd2hjePGQ/RRSgBfwAbi587r9GOOFLCzTG7vOSZNTiOowf4tSLUYhsE
vvsIlx92pPxF0DPvOetK6bmOGrENAXBiHT5nxMs12es7aVx0nIS1QwlBePR4AnvM
q8GloxnsTpjxT2qkQutkBilOUDxhIfffGR03s17LYEq8hj4DUZ2Fal26l8o/Ds1l
IUULTqzmGVHb5/6MB2352smwlHhGbGyv5mHpDj5eyKwWI7SXZ6sbmxNuM/W85QIz
MzhvbFmTLqYfga76XOU+veXYRJTzFiss3KGDSafftAzJgZbQXwqh1JF4QhyMXShl
df55ecLxHBWUeYXQNFDAb7cIOkgRSGlu4YwrVRT7ccT2Y5eWgHTVSMyz6iUdKwMb
8Xq9XPhs1pacBB89M0leZbA2IwwDj0EZDaRgR+wZyS5sX7rUunMsycIJmU16xXtg
UTBjuW29218iEDfiw1UF0u1VFPbYKVlMxEudgZbPA19Zp8qaYB3g6hM2Q/F1FrXK
KMdJpepp4Nqll34ceP3+/VkdLiDcFzDn+b/MaGsh3LcKGB4O5skb11FEZM86AwzI
hQPeu8t0GkKo2zvFRNikg9ggBT0GCLMhBoXlooFTfcN5CBXgHinuUJ24aa/nwJ5a
jmu1k7nwXUlBitk1o4RrK10y9qQuj7U3WYzqr8VubwoF2MBD9l1rgafuMgQYtEKY
NrfafED//H/gGcbgLFtLenUz0Hz4DXvnc7uHLAAuBAgArbY2QEVnrek0WyEDR/bu
qj5F4Ye7yaq8wZe/FEJpkmjH4q5xceiLFeVCXJC8CspqrmkBlevYtoL4QNNXQsIC
jVu0fVifbi43gr9xCzmE73oxK/kA+EQ5//Qy9AO4vBNbu7MqfGnS+OtKbHTbSCdg
js1wQpY3nyTIo9INUNc7UrbuBypr4+21wbBMsOMphsIYWT4ssb1asAxIKRSwuWNX
tirbjxzwB0TJBjrUvDSxrXvVtbDIl4DQ6oeempvJ5ORWqW180uGrQMXWOIoyMrXK
CgNpO/z1Hc4fFs+VsG5USUc0Frrj06crOFqw0Y/j1b6gTWxndP8ROhzKI1/19t+b
RTF94dfuTIbcBbC03CuO79e0wiS0142y8+2H4dtDAZWCvve+1QuVSFKxISL2eX4G
kOBKXvy7Zc2KkF/oSESphZd5caWUI3xFoWGQQuB4aNyhbtifPmMPnlDti6IQyNu9
jy73Z4wOor5WivnUaVjQJHHO4j4qkjXfkf6J6d4gpb0DkjfiGbNnMebPy6WG6XqZ
GCH/LvEolvQusCF+p3Y1tsSeU5sQ7SjS59UE8dKzgVg/SxLQCv/P3PDeDhWlt69o
qCPvWaYj0Sf7QP8mTAC7JJU1SnVYWOPHT3Dfyp4yoOjJ91hUkk4g3D61T4PnUfMC
VVWqG8PJ/Gyf8W/U7L+dqQXofA4Jq85oBjGo3qgyQEM8WZScZSeHzsUAy4QWO0Ht
icKlX5ByFy+y9rZ1c1r2opNJIDEEFGt08uQjgA8g5nVPpvoKcj81kBTSg6IInDFP
L8RelAymvqkeptviksy1TSdS6cdfUd4BE1j7f+OpOg9eZnVqNnWbjKtqOgBBLkZI
HPLRC3Q4I8kZyJPDpXduW50Z1OCZGga5P5qqfRLfPydWFY2bkAtDFZ1N5D+Pa5Ha
myqsqDQ+g0zZT2e6RIS1WALuxq5rQtAhwsRDN9OUqa+zY7nAWRWncP3gxNe7ExrJ
VIgKGpIS6qcmsX42g+Ujd5WNAq1rXUS92MQ1ixTDiyfcHlmKrEUMgAEuWlBjC+8W
qt5PdC/swgyi8ocpRO2bZBSgseApUwxMiTjSRM+x/rMsMJitqq5+ujFWCEIdELpv
AIC1tFFMfyIqwRWXMauw1STkT0657UkWFbj3By+7KD3nq6NTFQ9G0s1duSOO1afU
XIUVd5cb7I70Js+hJd1/UivEH95PTw1PGcLAH5RZR2CXM76wUfbWYEUqGO1lKR/8
tgwB8WM1C+KhiK1qkPHFV3nowZW4rbVcNwMLJt5S/NVz8ne42bl2hzRdZ3eTPhEB
+ZVwfFl2AvyCJl2qBGUqjwAxBP5VwsDJRk6gjJU8detN4FPVrwrFNI9sRtVuAg7r
bgtfayqVSeCOXFQPwV9vecjjrUqopJspYmU67NaQdyxeAlp9DYtZFjBtxEBrPkjm
HUYVH0UHcoNLrefUo5HABaIcFkbr2BkCEU8lEXEcfhxWF7/2BCiWZ4xHrIux5M4O
n5iM2MYjeU/lyhS6ijvpNlwJUElUfGGMD658vV32ERDc5CHw+F5PmE3TsK3adbEX
1mcHlQqsqA/rSlQTdaQBe7FaShC1qrUNoWWtWF5mOjHeV1AShJ2B0j/Ls3OkrUx1
B/pZlDa3QPK2ZkYcL3cyJCeSTm1XhSeEEH60w50NF/yxB4AlJku6hxmw2B84Dhc/
KsMQHYLgnUYKWSfw5lgs2d9ygh+12VAkGomQk4pUGUXPyizGAUMCLpdqss7Vk3QX
GGJGpvI7UaAJQCF9QUcJMOB9AW7mmM4UqcrSbBpwESg8lMvwkZM+safduxwhZRqT
j2NjWhCZ3Xl8wxHXl6Wu81ZoQDlQ8c9TsaxWR9pD2xJZNAglxK6YTDHOQlYhOSc9
BPYtHbfTh5G8mRIvYdgqEoUKUJijPeH5KwL+8NXvdrmTnrEtnmVQnDLJYuAEphaD
OaDD2WMufHKUT8R+SG0MNFWmPS4FOGFkRYrrlu4+01Q9MWW5eus/PCgFqPNC40F7
9RJrkd3qfGXPyVBIzG25rd1lwhfYOaEYiwR3jXX92t2ZicXSjDO+GL0WOcQJOLNl
vxr72l6mFnUsM61Yp9TJF01oBARx66rnLpdumStTUcFYNx+esgNxKifTgi39c0NV
HAWFFwTnqPDc5+jWklW9T4MQTZkwolc4YZxq2ptBY1jPS6Q2BgVhMgxWCt9WkflJ
YtRWlryrrt0lGFhG49maTcE+bi3jJshYhnXTV38yRyMj68cs7n5TBLCwrX0/kl4q
rBxvMm7GSErr6iEJcR9heDWP+xmYYOxJN2ZzSc3hTvFBz8vJpHaEWPc877Se86nd
DWy7eLIYhCNnS5/0GR4VbBDOk4NANMahzw3q7wvc0+h+dsJ+CsYSCJbs8jWujMUR
1pvn+RWdYP63VcS3rsLLP/sqStKIJwjBccTK+RuRMUjrBoESs1bbJaK3qWqse7Z1
yf7S73AIJ1FZCnALEUC/VnQMwNYJDbWENqPip9iWrRBRAyB2r7RYhJ7RPpzUYgTe
VnpEqg4wT6TtIgv2RBFlr6qirTaFTunDm0m56PpMhN/Gl0k3URFVa4CgO8HKZYPG
UBNoIh+McLIZEQmiqptsRc8FDQEmy4zuC5HRqu3e8zaSValTDHqX61jMrXb4Xcbc
k/JsUFC33Ig1eZzwLHakjdpmY1C0HgIANY1ZUcpuYHy0m/egLPDv80Wlfhyf2mOu
T6c29Q3bcUP5HiZpUlsXGjGKE+aFaV/hXGSS3heAKXHIrrB6boEezK9zzMwq6HqO
JGAG/+idOTMKm0RxSItXwn8oQXtGa+ra8WqzfLcRPBeKmZD1osTFq8qlNlbt2nJS
OG1N41NUyQ/A5JBq1Qc4PUdNuZyVR8rAg6b/twECdQasgzym/aRnxNcgnAee+Tki
BEaIePseGSXmJ+F085O7fP4Q+V1PSIEQbnfK3bXNYzE1Hz8ZNb8s4i2VwQ/FIOs9
/aIGCzR61TJdPJ2ae2mlosOtGDVROdItr/iir/rOnh3r+khhqeveGfBj9vr+nmp/
WR1Sss9IFg3RVgAgCWAcpAgYAbLQThQfA7Rx40lwHCD6Pdn0+2wqTruyvTR5igBw
O11sQb0fsDJukJS/lkOBkAZ39T37mtcp3RuTzOcAmmthwIAVnGWF0lR5W2l8lYeN
L6rOflVglpskPxKfhvi/LpnxzGnsQ9cS1ndgvuSN5ub3tfoQqn9jFYQM44qo1Q/T
Zs8VpyUhDAqRZWLeWwt3pUkbBbuCKc811DbGJzaYPUXAjIMDxQFfUNZt0alHUHNz
hc8KkVy2HwpkEAU6PpucLd5Duq69ZaXo4KZjSY9c8zgKLJwfOIKPdfefA2e19imx
4FIThV8UaFc90IAPYUzNE2l1jeTCjqsePDyDd7WNRd8YSpaTPy7IiqFSkMJW2CYT
/RZV+2RdztoG8kDqEZZ0gwZ1PWUeTU1pA00X/aO6l5DGnLV7qcjdDUl60fIaHjyC
cXTSTEj+a7tbEo8VnwyWzVFs8E36csh5orSaRdpXa87JyPbBPCPYHNMfIGvTjZ0f
qRf2soFIles5T8Pw7I6Z+nu64YkjUSTip2sfxD7E5rxRF9l7xu2hP0fodGSs9Y3W
f0FUTwUZzVKxya1R+XsQq0A9L8BfgYv9yM0aZfzDMwvtKC7DF6ECd0mfhiO8SLbw
o+mAXPEAMP7cboQdszZZMllWTpLX7vtzENjPyJ2XNc5GAGAPFZmkNIzwkyvWEN7h
CQfCMEE4k0WhTvexUQ1bKw7mPgJxXt64h7JCogpLOPhpIsL1f16R8UgDN06Zk2zf
TGzHDRgWKEOcLRyie6S81iDuwaHiUF4F/Lwk99sWhVY2BO1uGH9ag3JLqn3raQBK
ftg5hr8UlP4YQVr+3Rc0qFg0bhZqH9k8MAyu6/sTe5FZmj9dA7GxKo9ttQ3sf0WU
g1+DU63yM/9vL3XZmPehSaUp8Jh6fCfdGQHp4xaqxQJxis/Mb0uc2aCpJsFzfXpC
sluzEYEYJAbgLez9CUm/qtK6gIC1GxuOK985dIm9r+7KP+uYvSyo9DiPvJAB4YQ1
GfN8Uf9TNUY8jtai4h2RMdoo7ZVYunbAJ7WQWsDXmEFlW7QxekNYApPHWyRfXODt
4aj2JKiOstyWHnrolR8owb2LvSTAjDprn7kqpYLsDhY7jD7ntr8LdbT/7wsw8BAT
SgSUZp/cqwPNo1BdNJt4rzAvI9Iijjncr2WtYpgl7LiNx5nnG1s+hcIKmRRsBQ/e
5HygKsBTwYvXgRuGnzMh5k6oz5yqa08/HpnIbdC27ke+qmPC1INQRbtRvzORly3l
v9qzfetS+nRtVMcB8lzi7LT9r6e8Rw+/n5cLcWYqRWNsn54J3ibYQ//zwLZBecKz
457x+TGG/IXcn/eseQce7Dz+lkn5ClOLSi4FpIiVv6PcBDMYies/ytXkXU9mxt+w
8lpE767wCg/kSPmZ5thIJugvUI5Y6IpS0WxF9pLKMgBNDntiw8CwOD4LMn71flor
dFRR1gLpGbB4EBDKtPuYez9ijk0RNoqrl+4JoSNJXCNGIWHHPvARzxuxIe4YT19u
vzyJ14m5U1A/pMvLxFJnXEY1eJnzKzJ2qgLtgenk9bZH2sEs0iUouv/T0cWj2kwU
F6qPWF7mW62QV52XZKj08leCYrv9LVeyI+GnKyAUEIPI2lPLaNeAgtjb20pA5a+I
hhJWLxh+FE2G/k3AXweNq7SfJtHiWiMcAEAb9q+G1p+Lq4eaC8DouFPjMfK+v90H
00k7TivYutwa+UU09POYxFcOQnhS/sX72JEgEgyokoNPpaXlnCw4tZterrM3eH+3
2V9oojBSj20SrFGpwtMk1yzC46V0giYPxMUzQ6Vzg7r0VE1iku39oLqZDhb6k7W2
wYSKnuLsORdD6YGTtr8xdd3jUaJwrZwf5M6O+vW6EnukIYEBopFFkr/N4Gi264wC
VMcLUzOL9teBeg4vAsf0Kq6oAT3f0DBm2Qvh6KmK2gv7BsyKOaTwlvuAZ3pMLR9d
dHgBHMCOeCWm3JxQFDiLtUzT0beR12sM46a5i6sbDujThLdN5Kd3+B6/bHBqHQFM
fmhMjwfDy0MWaag/nFQYBVsF/JnPGR7cTpcPbhuRO9SLh4Ipl6wjitMcdOzXZmGo
t2fwVPY9BpdsRVZygwxK68tQb98pLFF4qu2jR/UllsuiU2LzyXhRC8I9yvkVmoZ7
GM+Sh6DeO/NYbuWvlPvJEg9bY6hlDUPa/hinGHzbVd3mK3XW/6zMv5OKE4e1gvwa
ukEIkzSw7N9vb/dcV0JDX6TyugucIFuX1ME9giifcyIEJZ16EFQOjlzogpl3igDr
jqxZehp0jJ5mi26M8AY8LjrKUkLKYC1uMEapApxUioF9il+UK3PXsidGXh6JTgPE
iuVkcvvLbGS0cK4Nx7zvtSY2kj4xq9vY266UdZtg7LzyBn07OadFUe1a0Jh0iVps
WqVyjvC47+NCe7tskDPHroydCe/yrG+7xHT7293FW5mLRUUVT9M7yBm2u4LkjFdr
ISqORkR5W/mH0HvQr/khyyvMAxxEiv5ZoR1q9oOZjdK3BMNT8VOPUs/FwggoYkcL
481+2E3PYtcXlXurHm+TaRF9nV3V0YjC0d5aDcX4NXBCnQnEzJVaehW48Go77PWO
hIJb+rem4F0ad0wukke6ccQl8s+SGX9zKG1E5FP71h3sevralXPKY061JmMUqTjM
+u59WLtBaw93B4LZGhNcJbLNuyrkesUAP86Sr+GjlqZVLwmWvYkQTu9lv+CNZfVx
soUGFeRjCHtMNr8DVj8CPGyXjBP1rehaujsLj2WrgJ6VfyV1Tau+Qlly+dP0L/5T
soCYbGTUdis5PRebg3Su1ikARpTTaBI0MxvMlTUFAKXuxZJrrTRFg5cUtTJS0vhT
LceQhrCtckbKU6JAGVJkmvw/gHjtaQyqwua4ke3X4QocWURyjGr7wbcm7/5LIMLB
WWjOJc5fWSLlnGr7axQwOvonXKjaN9bRp++37zXTcdh512E0WRFdgudcWtt92rKJ
krlIWZPfSKXlHsl73WrNSIDRXRVXSH4DSofSvHlypilqsZnf3n1OZz9lz9yIl4is
syNmVpWYjvUuKsbFBVHGcnZYSJ5AnfKryD1lqZuADHhWqgBw31vrmPHd7JbCh+hH
bz2qxvp6ukSJcKn1fFSonnIRslyvv6iNX54DCojDz8zlzII599dZfd7PqW0lPjSa
wQ8RFJ+mCsTvYZUZSEKl5FaVL67LpmPIbMLJOC7g5e+GJQLnSi/me9OacE6Zgm6O
bds/gTP3A2pXRfdkw/k0+7iVwMY0WkgaC2PSdoWxTsZsRFzlmW7d7Ys5DIVaEU9+
swSbvW6Sii5pei9/tlSaibBVXUMXek1OC292zp1ZV/KD/Zj8hjofKJh0Dn7L26Q2
i+3psVy+foTARHbAea1JTvhuqFpMtFKqKFuz8Pa6u4+3+0opKKzDo7jiT2wBHwVS
wmXvxgBEoekT3A12EagMKqBhuxHgGNsFSQ4k33Q5PozBRyJeOzySWosFf0LIzK3u
8yGhm9OwiUUEIwszewt+YrKLnKay0iC7yyDE/wVlHMV604lcXXMjlcmqac9yuYcD
bEaDJeSZXq9DkvFcFE95EJ6D9wxCTgZNoiIFP1ymW7Fq9fyy7oxna5Zu1JvpDDC/
X7EL2bUUXE5TrtUoGzgJD5onHwgRHtlGjtaOZM8goUWYnZTvrtLaiLk9Y8iVUH4u
mCi1Uvand6Q2J2u62znL7TFElzlxcg2+YjRs7qe7+3phlOSSjhLqxXbUlEXi0ZV8
SwzBqetrmT9Jz5VuyV5U8QHSAkNDg8N/HYz9Hqv60UGAKJzyrm+qujm6pEtR0ahj
goDw6DEVBCLYwT+7jcfDIBuWVVneqLbxfI2Iw9cfi0oNKCDAo07C5ddLC0/ljm09
gr3N0zgeSqD3oZkk6yT6zQ6PWfA6eky/bsUFbE4UK/4cUfc9/A2KCzwMQnAXnozs
oCoWfpbTcNR5Ep55PkbOh0UYQSF2aCsEwukCJnfbmo3ZgzbQNQ7zGu6NldiXAk0w
HoewWcfqH8kCowvYNfoPostfO438HEx5mnV35QztTcIuaNMd9sf2CJli1x7/3Mo1
JA4JdcRbilVofnexs0dsMZz5aOMgj9Vu96beM6GmybVbc9fwXmpUP2U6fyaM0DJz
KApW+GxRgz/1mNJVj8zfYtDLOiXv3MOycj23A1lqd3ff4E1l0neiqE3G+gkJyrzG
4YgTboMnHEZDkPbp8kIfpwyL3Q63ZplYm0fUcystSRskTevzNj5rX4NFUrLrNrkh
cvSPx0r+fi3AeOKmmy6eaDler5Tb+c5W/UZUF8NTInqvjSKQ5jXnSIoMn/Nu2Oia
dUSVP3QOwKjyUkx05lMUXSuneRn/X7phmiRoy8cEeJsXfzSEPn8WtLN1haRtQTC+
qeNTw37+vOnhey4sBJrfgyuQa2j1fOTd51vu1kpfXY5CZh1kowxQTrVC6z5V31rG
JuW3njc9orkXqw/laMJ9CScmaNT4L3vJeJfx+AZoNJK9241Uvv57Qf47lJ76084V
V65NIwqfHXJlWOmvxVSow4CLDK7E3EOs8wIl+ZNs0eRqLqPQyg23i7AXnSvXVl61
Z0QorMb+NUAstWmDfhUA/S2VkJqYbZL19BQDaZL2BUGW9+nHxJGQcsWK5/cXPkq1
JH2jynUm8cSRgqngGF3PcFgVbcM0AU1Rvb4ph2ygRml05dHqCCgHLVVtiMrK4Di4
hxyUqtdgLwbw7ELe162caD1AY/43XlGqDGVJq395Eaix10a3B1IE2aU5c86qdgeO
wiQGQK37jkxCKx6Ey+qaES3jIMawixqVTuaCCBp1r47PD//MkuJksryUmo0SqseF
Kil3oDBT6r2svhWdAmsiPsaug+Isda5QFA3UYaUA8Ne5IVjb0LS75+hK/4EjaKiP
VP9TBOPpeRuhUXaCgo6WSFnXIhSAeXCyHMuv886zjHk5V0bN9Kmk/RrJQQPf54Fb
uwUayNbYijAEqQA08x7JyIkmg5c2N0IRoKonyQkYhBVehgaHytw8a8skA6VjcIpx
xXbZaaggRHMDre0czjOJfThbSzVlUlwPwo2K4n/hoEF7Dn2WND9xN/3ew1QxNtas
7KJTIoJz2rQfIO4pGNOqrCpqS/2U1AwkXxep8FnAnAN0VXIObcSlJheg8nhh45gk
mWHSSDX5RZbiinOFrFJtmkDqSrl9M81Gi75Uo+WZsEyclU2YjHwd269p+ZWXYBJB
LO1IoxQFduWjFFVaNHt4AwaeXbqT7Ha4AHQcyySBJtlgCVIYFk3b1OPM1hDf+Pwe
Cr/JB+oe73Le8pwxvMChDyn4giDqMTATSPemDCFjku198/SwLdaae+IMLhX5Ub16
rB6DfXimxRkWGgBylGPor4zxdw2sdWafPh9HhcM+6Q2cWOEXCGQ8GN2LQON242Q+
nlg3lm+4RGkQy8jOOo1UItvS5wCgKcHXYdz/6ALMrVgJhr+bLRDb25gilCtiIUTj
ilnjiFHFPRqjvys1mbJYBeYCjOGVIP0l5RWvCGG3dFd8IcK2qpCVtvbfFjq5V87r
hh2IomdHwCzfECbomWC5L8Rx9bTXMKwzgqgvO/nQI7R/AIzI4cXEYOLpmvgh3Zge
1lYZTIiw7HIAHkY01Z27HLFiHtSbGJBR/QZo36Yv9vU2E9d89rASMCOiGOhYDpG+
cMk1vEYzmpbmXzHMrM35pbuTEMF2K/G60FwRIya13XwIpcsSfIHLEjNfX1ZVf2bg
GkzD/HLCOENoA2fATFe1KzK82R1os5gykiRQYP0klnEQBtQt+xl+x3+DfEByXk20
TJO4FatA1eeL/lBxavjSUxccV5DQVqMqZ/h0A8Ui3YjbGXVfvzAtJdiB4JocEA31
ce/+5tUnXUs56F6f2Md1+osKTc7qTRSP/Hzd818XIpYQNCXDZ4tdslcOAeyzZ7zU
r1xLvwOIbmoFIo9fC72R+cpPaEIV2FCRt7opgtgJe8mBtQ8GQ7kwxVuHUIFeYumV
YmmrgSoM9lwDHrOU8QNF7rp3aT+s0LWWIAsWINGJsEwInlAcgN2ubIpQ09xBlccL
UUeU5HCHXJCpCjb72haSa6HjYPX7zyGnqNBo2cCKFGcjTgbPhflDaJd9extilyaO
XQ4XhZX6DqzIxdf8vbNt6STW+czc47JU4I5dG8xn4MzjqusPvAjZaJQxq8oVj+hb
tp9KrHvQ2X17QDuXHaahb1zqmYVcvjGAcpygE9XOHDObIe9Xri/J0RrOBxf41TCt
SbA0h9fls1brxmPILC5v+wJ3cFtCn0rwt/WSiRAgRM/byX6dfWpZSXC7kSEblAVv
H7G2VjMHKfLQbkl4QzfdE7jJEM7OJ+WEU5fp3lWZsq9M0Zfohf2lBn41zPl2naDc
WVEd2uEdcRWOi3NNaTMIY34CCMYRNTlE2yowjekHAIGtxuVWx7MFGnCzg9Tm7QFV
8FWDtMgsYyhGGL9kxYZdHAqgxtaEwFr4sGNjkg8MtgDQfd8UyQ987jAXC7tMgMGY
Dcr83FCe4IAWFrABnB8sh5ILoDjehghM5tOnb/hghJ34+QuFI56UqsjO63iRXtdC
DAzsrxUZdD+8NZpoc7nL1c6oDrRfuy/0fKrhXc/n20AmwUoC8fV98qade10X1GUf
wtIHWEtb3i9L9LCSsj7LcAmXGM3hv/7m2os5ssFw4WY7+2ZDi7I6FA171eW0RP54
rRWki9Bdig88uXQ7qTnH4+Nh75wEBxPWofpD9VHyJRZU1u9WLWqDlHo11/faF0dU
aHyHkLNOFqRw5YJXfoIyGzC9MxoBNuTUa8QZ3UKqzGiNfb3Nyb90Z2S85YwEhVOE
g8YnQ37wG1augEck2ZChXkCoDhW+VSrnPphIsZ+0rkrSgZXNpvFPNE0L7s1ZYKO+
k7Z37I9TxZOqlu081aj6zPpDun+QmvDKJ4tTP57YUVAuBY/EiNulsrG6SDibz7Ta
jczTMFpRG5eE0jgyUS/jxLAoo6Hbcd/PIJBO+L9tjeDtWUEEupIDq739fCfvn5Rs
S7lg4itBUCVQkzmxm1KVdyDiOVsO/AqTC5/pc+iFT/znxiE8FqJ7tsBAWBgbdGIW
tjJMXMZPh359esatKbwalYut+ofQdka+CpBvAbKa+fr7JyfujUkPT9qyr6uYYgwc
HTRZESY2Km96/Ufw6xITBpfR/mhr9ZZp/6Z1M5D74SlJpfS9U4N91CmedFB5wEFk
j8sTNGj1cTQ7ekGBOhlhN6mN7g+KYtwJs6HCqt3JvU8vwZWuYITPOnoHmeGg4whV
vnyVKzc5LkTahkAQsaPu5N5QoCWRyly1uh6VNXjnoL8vCfJatybZeGd09ZmRDwRs
CRwq6Gl+oKr3LiHh94UMFwzmUJFJz9qF+DrBjNGoC38zTZ547sHSm2pWcckUMbCE
lsBVcgHZrin+Q/Swk+tzMK57Bvkp2YbndWtDRBDhTy3VgDHVmLfiporeQqxRdlmq
V1Qod6JAUplEaKgKKUxAGYraGrub+LOTlUV8RT39rSMYPfaFt9S8X9x+Fw/xnMwi
BMYHwbP30KeIXjMtK0ST+zhgJ0XOJ2TOqLqUL+VXZEptUXkmqsLspUmKIa7MvGSC
PASdvFBdJORSPGm+RmqwewIj5sMlCjIgO+0aa4L4pnkufGE7XIMEsSl9z7vkyVOo
QekaOZS7fDCACKckOz+ACXwawzF43C7gtVRY4xjRfwas3ejjE7X1jmMLh0L0MAGu
oSs/tZk2twhH8y+ZEcETWD2525URVgM+E/5F3aUxaq8RfFae8LZi9VP+jUcEJv2U
vffkhxwPyvslRbiykE6y8+msGe17ysoK/7Lz9WiNC6CXHP32J2W1SHYdBv5H06aL
088UJCUjf+9ZtrexcnO2SLcMBrknFdxpg6sYso8mspQdntKVs60C9oKj2KRcsNNV
DT3fugAGS6v8aQbzdBG2n6FtN1aw6FJshzSK21fwWYQULkbD72lPAb32sJCKKj2X
KXXHXxPN8THaH8lgFcEUF1qR5znZ3zKHdc5fhXcdgQ5hrVL5exd12xIOE9uxzQmJ
xpMBGXYvxTdcwP+3zZWXCHTm5ENuJxwCS5eoz9PFcz2ZkMcKiWS3JjGi4GY0Zxdb
ddWPaGx5CPNYSu2cmih1ZXXBgVeBQq2FIETkJ34RGkhg9EAWU4tAgsBJXYiTw1X3
YzbBQqmxsyezW/bnW6KHWAkAQphI9n1D/Xug72JVMZlz82P/8a0MK7NxGcvRsZON
AYkBN3D93Mol9Pey0jwbSyaILmGEnxB7bBWOHE2JBKwNPf0rcat/55MAQvognxdl
+Q3cCIL9FS0gYm5G5j5ULs99GNkUtVAWI/aYyJRYfhjgTi0VVwcC6JpsQ+mpW+lx
g870ngAI922wbN55/QpuPFpFYB+DBYFKjJvexqKJsgiAJZThXGDoWPtdrmLJnx6p
PsRz9Glj6oYn62yq5t+FhDXftKYQenoC9ksWzYiaU9X0uHVLINkSb04yKMeMHUc1
64yrakLJuLjcNkXY99f4YwEz4V9ssUpJ1Gq+SjwXzsfv38/dy1LyZ4r48Mrs23qY
Ldv78XVFa/AwMZUs9zI6ciYfxAcmaLmwbTewsA2q317/5tYrQGensSPfZkgGLdTk
DbqjuGMFEV2lTr9bxWKZwJhoEvyqqClMQku+cCAFQ1PNXMUqt6NlwWazdl14Nl+P
XwI5W1Ble7eIvydw9DfNSUVxMh+V9q9sK8j8iFOn4wO36ZUN5xLpuwMXVGIlToVR
Dcr2CzEKFnrud63IJ5zUNNFAqmZvfCgoeAuDAnnnEDoj2PsePq6f7U2zT2eGR70C
E0odV7vdlDtnUkx3qbfiL19TzLNMlQGJH8oUH2zSvqLPoe3NKBCeG0ANeA7aLa1r
lBef0iVgxm5qrWd+NgRBLTNPcZGVZ08+ZnXu30Owi2bfbsxINQEEjj+n9NG6V7wf
U4jULu6FTjB1k8K15rBw3L/HkND9inS3NVJJu1z5UgV/5+HiuKg2GF4Z6nGqF37f
KWvZTOOYp8giFYyzbZZ9CtZsLW8i3V7XeRCbFG4+6zENUC1cB4vsKlcb3T2tP7ud
DVyBJMkMnzwj5mjvBLLpxuCxYjQLNIHzvsBw76718xKAjpmVLn3gGHnxdkQfoWjm
8EZ82McTYX1NxUQLcJ1jcQPDSiJjvYD3aukmzxA0fVRRhQm8msipOsfRxC3TRK3S
SsoFVHegBUJQkhXJ3efGD9s+sVe+lp3fkgJ7DQWV+SQXBe02AYDCMHC/mahNdjH9
6NM8I2HbrM2cziccoi+fmicHTm8sNIgDZP3habIl/jc5as/orx+Gg1crZ8ySoM2V
53xOJlYZg9raHSyltkw/9b5Ah2TiD6vD4M0vH+2/LoykTW8DGnqe3MHypwJ4vHc+
XXegZJyDXPnl41BY5yXzYIpj8RdXGpY7ocxS+fmjdA6A7yXymZzxU4GtJrT8Hi3m
n1I4sW2xtAnGATvLSIfUZU4o9ecbqV7aVweL5oHkjzysdU29u1RsSIlX6WXiaoUT
iQ3klS8zWJYN5YWi8vGsXEbMi0I10jsMYZdQfgS5OPd09cJpKjIZ4e1wqefqYALN
mJnJvv7kZy4TCQmvEv4VAT9xgDziTwdIe6QDMVyuDH2OSjEdXVTrkLaI/FZcomPl
yD1E1/4NfQ+7OUiX7tF0khYL7eBL+DRQbSV1BTF7hy+Ej4ezHOTElJeiGrqzt884
MV8Gt/Xf9yo7co9We9yDmhBcm9lhVNFSRZN5CIwQZ090CoCoJq8qP/zAzY51kt2g
iCFyAhgQo4aoRVmVQ/nIUQCkrla1dFyG1Rg3n2BnxrXpgOC6eflMQ2vY7qzqC25a
8GB2on78TjCy1fjCez6e5BS+so406ZwHVOB/giB4K6/joA+TIA4zuj1kG0reVIa7
4thjpKpaOPxvBtb7YXCCJiPetOFs4TTPzvqdsYp7aIYTuNxkZBmJUMl6WYcMjK1U
HH0/jaKy7wI/ycv00GyQsq7VuJupFSldPGzfVnrTFRW2C2FS87rC7FgZhn8kU+mj
T0/HkPmeclfE87iuak2rfrKaVr7wABFNMZdXyMFgH+86dbhjLA2YuD+k1Mvp6dTd
XtgTg/5+eVhLGzzl9ZWIEjxNfF/HVSnpVrTQglSQSs7ICGEQNTL8b2Pc9bxjRZDw
jm69IQBsibjInGkevrICxNFSH8sA44U0+/mSgqwLjGzEUN3CzWets6YdOMuoi9vw
7dEupoWukXODs3+5JKftj7aNYgsp5DoolSVjSoLSQMICDoXzmA+TNSa33np2hbSw
/djWS1QeuFYyqjrjgs6cdNBhfji8u+crhg6BDSM3wFpjp02dCiNklux4Rz+oM73C
bLZqfEOIiVHNwSM0uTjZgqhAjjh00WoM1iBmsJ0SXNTmUnz9kVVWqxX3snSGSesF
ynyGx1B1gs+bU0bq5uWcf4f8aHWW+auqKouiRp6Hd7IOm0mZB2FEV8caD200plMr
hfBQuCJ++L6JPxLafgLk/qPLITO87rRaJ7CtUtGoFOMJRpuTXjvQ/jPi+3N2QXbJ
S3WxrHemN2ign0HiwU8leGtk3ELjxVWwA9dN0jI5g30+K5f0UNtnvw2jV3elt1l6
IOso/6hxRcl4kPXsW4WtLisl8dHCH3m0fYUn9BbaIDflub75+DNbhRkDyyncwqiU
vq3OoqQJUTC66P+winz9E7FiTsKveiw+gLDz0x3v951dFfj1JEN9JE4sDQRI8woD
6rSSyC1Q/nx1U2E3NvlJoumUzvaPIesh2MXY6b6Gd4Pxatlhk8lA4RiUBtG9zasw
koz0XD5x+6VXPxpQQSXcvvpkW2b6pPPm/f2+wyA11aBxQC67UGNstT4ZVsIYxqHG
l6A0MoCrdAswYcAu5SvQcA8JdKQDt1GqwK2HQFtqYbIHkNTJOvraxd6H/2HZK3j7
kV8v611iTdhxBqq4A3708QM8eAJgAT/gk5Jws65b7r3CKXU2cKIeQlG7tf9CqFnY
N72jvDqdCbcigAeKgKvViozFTfX51+j2fdjbhShtRwNLLI9yIc+eWaD/2qjrMIkh
TBN2RrVmkANMW+VrM2btQP4ESHf/ZyiqVnetK0dNB4bTSZ00cw9FQ1+yTFVPdwD0
57stboIlUhLpB82syrHKg1mhdcaI8r5r1sRjrFy720S/sLR05gcdD3sqOSFnM5I1
sh4oWYr/C/sEsuLs5asQPlhVt8HHu83lXkK46uGo7TPjrxmhxPtvRusVg6CHUNl1
UgdcQewIXo3Y0WCtPUjeoFk4vhQU1lBq9p1NBMuBRNS1LFXRJswPDKK343Skk3eo
ToS2wIYy7EqqZ+9ex1CWYe0677Mx5MqacJgcIDk1Rzpk/DuDUe37slozu4g7IvLH
HBhrF9AmPfI5riEfAZgPlMo6+GZQ+EUFrRgwE8ps9WxTzb2kHOWhqUoLbCtEjxZi
n3VwERxbtkCJJ8lWXG9iFYd9sYJU1usejTWBMKadJ9VX94hGWDQ/fda646sIe+o0
8Nq+IgT/SGCdW19d+tDQCHDw/53ujLptBaJbnn13YST63iLmSJkha2Ecmxdb0M8N
isSZQ2DsiLZo2/Bb98wz7VrjArkoGVSD8OFaHFmJsVOf1zwwPBPE7R3VmCAOkhoa
rWaJSiTLjrVB2FIp24JK+GAjdkWWQoJgK4SgJQCmDhoAFUhPaPfLUY6foxi1s6rk
fd/zumPHAw9NeweTu9nkXwAbI2SGmkp+Y9FE8bnf6mS9S00gQ3gfYubrsc1ar/TK
LVoBEMCyktTDhQAIMFb1FVHZP1jCrtDwJu9oQDR/VTx3vObVkGDcI7GE/Bje8Nge
xM0qRXRhskLcE6vbOPLGrBg0BPLGg4xvHjEEhtEPM5GPDo257Qs8lfDyXdmAhe0u
Dz7qpNBb0qhXN+CqSPL1pV98keFYNtIWLxgdwzE2TPEAUAShgqpIOlSP1ln9leJX
tWQqyweVdnFQPSBCleuGPcZ228QsjyeuRDam8QCTRyw1tj5f5ssAFYyvFjDVOyJ/
yfMk+jvjsaUwueKlg5foLpMyQ2ngIFt6nlIP36YOkF2CqX/hDQ+umgQ1jQxAO1g9
vcdAIoLAkFYkDkuMI0fgiMdeH1W3fQKDSPA8EYDeN7IjXEYD38RfZPKbjAuoOFzz
Ijryqg8hTa9riDIF9l421DMT5k4gtEi4ec3SwfYeLHcjU1Njqo4lpDM2dgUmWS/5
+fb6wOLZgGWULpaAGmYYhVd6gnWghp/60w7FCY8fO7tkqqp9a0zTrVc4hRVHhoXe
jXeEk4M4hkFVHxOsHhHASm7hNCJQmvcex1WYZNVP0N3ithCgc65xOs1ePdvew22c
PZdTmWkIXKWbgdMcLl9XnQWhT9+4gg5jyUXKyYiXpD7spieHyJQYLb0NViBRhqQ/
ADaFdpMdOZQVr0NUlL3slEWF0Wb8J36pE9I13yY7YpkELgI1qkSJCX5WIH6Q1guH
Rao7SrSyLpFk6lLmHdjyEsmSA0MTGxbIaY847p69wPeZF4zg5WVRO8/2eGnr2ESL
LWcW2ThYaOt4/qALfNat/JoDHQ0RafxlCGIsVx64Ves/e5OGiNfspeeJBPtN5Y1A
054gH2QtN7D+5bNatXNCe7JmSWbeRZBQ9sngn8gNapTrFVhvfpf8ld6090UJhqjB
fa1NcezvPda3nhl92HA95As5yGABxEjMtfdXBUyg/6+lLO3l9JnzOvi87vuVktxp
wO6Gv2m75IUiT1q1ACLG5YGMAWcNb9JKJ16WkCdswPmN75OVRpDXOCQEns90z0/V
2yJPEHrCf2eR6UN6BcR6vM0r5r8H+jQDWv3xJK7IymE4v8RnUQQmbheSRn2TUdyW
SiBkbKYA6MUn/dlJXWGyJ/UicEjzNLny9JfuUJiWleV9otn6dmQs3ViRThQC75vA
4/V7gVuv8hmiybOLyIpGLenWJMO+jSMKEa6dmvuVLs8YdDI+7i2/3JuBQ+8IYYq1
gzdVAJvWw4H1nNhMysD2SPDXYpH45SPJoGlzoGojFjDliMGBNpk2i2/Cy5avdEDu
uVcO7ULIh0pWWqm7jXD5RrsJiasUL/JLih3yrOxaPGa8TWl0gWBhpXjKSSRMpm92
3T2/W3I7i+h8RJ0qu22Dm80AWrZxjHPpQWvunYStwz6ITIkqtJvudhuun2cQdkVM
fJiKCvQwVS21Nam3QFjdeKlDd7bm9/j64n33tRKcu5vulZ4QHgnhCCGM6UwTfjfA
alv2FnFC0Kieu3UfXGoiooSzg+VrmCy4gfxJoQWhUR/jktq+f2YamGeslupaNEsJ
KD061855T6Pussk9AYZzHZXwNa31bbn3Y1FFxyR1OGyLLiU39kY/OwV9kSjkpxC4
bvqYTvIGqPG1awTpxPrxBUCJCu2Et59y3ivjDqs0ogRDTid/MM35t9UXuOzzT4fE
5ORjI8tQSSW/qsxbr4b47grdLqfSP6FPISJ7ExscdwQ9dk8lq7JwJkknQjojkxc1
DrY6HfW34FEgyIxKyoSq+Ahp/ZzI3qxom3UGcMpoYeahHSk4jfYY1TK2ShGcH8XX
AHGm1tzyQp14sb8K9hchm5abURXLaAEYEnzQxWHH5Rdy2ecs5hhdtzYmiFkjhWkZ
4oJADLIguVGHZQmYSnXqk9y4DNiy7JjRtWlZ4Vq9HOFS4bpNRvIdsx1xCpq4xiDK
6awrL6bN1uiCyF4DFb4otDuMZZceKgIyDpx1zAOkqyjCdM+V6GNR+KVDQGz3PV0h
pp8IzQdNZJDo2ZQVOFALfuFRqhcL8EnjirzkzDoBZDm/fjCqlbNgGpINiOSbb26V
FhUw1ziAu6vDUsquPl88Eb5kGn9tJ62AQPtr35T+NIvfWf1d1NSP83EZyZINf6kF
m9EqlTPooE9SdlJCfE1VkWvxjeefydvgu6fu7ayVamWwfhpA+8I4jbygED04/c8t
Xc3SS+woCR0JYlkUHugLNR6mZ7U1vVYTatFzppQRXqJ7OoNxu3JFaEps4bANt0//
ZAKKLqLqRCpH9wGWYExnfZE2Tib8Joy0e7vwPxYZ04IslrgHqjzoFD4uJq+ZLAEP
fDqFtZwA3RHX1ot1QxltvUEGibR8pA3qqvbyOJ3TsPWP94RTttO/ROiZFuQjdZKd
62NrCpwQFi0NTkVe1tfUakiQqhUsiTVCTxZKHf+CSrX3Bs6mirAYhppwiF4U0HV+
pWfEv960r9Cjdfzfhv3rJwGjm87lVy5LK+zrx/cYHQxO2M0dPlsJLDZiIGqlHZPk
dBh/D/vY+Rx7LspY5uz7jGvE0F6drWdR1c0gKIuFGD83BzTpxSgpuZC7bLe6ti4e
XGyjH9hthNRn6C/tYOSz+cBvf+J0C7tJBOmV78OzQNvFPoooW+9ebH+2h42pW1ho
dBgvDBKrzk7gbHN9Rg6bePSUu0CGQqlyIxB5fMSG0O2U7yP37H73pXWc8e6JP1YN
RryIDhj01K68543z3EqrHPuuX0dqB2p3ye75t7+g5RklWi369QxeXkDjlN4YpXlk
IU3QDYj9dxqf9V0b1U8zfJ8OoKDqwS6yLCcD0QYOODx/Ow5XnyNatkEacvdcqC7f
HMxScLJk4QfRITc711EwKUkJPl7q5z5GhMxBPHjwpKzDGidNq13zCG4AUXKLjN9r
0YDOw0NiUM/97KaW6fwg4q6gFaXUbWDZuslTHjLBOLLl7h2cqkJzjHDnggJ2qHve
81d5D8qDfIPrNiXdivBqeJrlpA5Scyo19QiHn2HzNU/CIBm8GdbUQmuqCffAde6G
2hNc0l/pkdllaJCmHgl+C1UGu4q9PlzzWaQ/IUey6SFijOzGdJVXuUdSmakIvu/Y
acKZrRjovietj714T3N/0d5lIoKuD/6qj1SuI+BAfSrYNwNEqCf0l3ligGyUYNME
QLI6VVZPVlJ78UV9/B7GxNFtn/S1+jeU3cEkP2Rc1G6EN+gOQ8FRrasdJZtPLd6B
S+iwtQWkfoyfJyCMLN+DSS9LO+JBLyzJ+v77stY5UBIlTry5jBE4LKxBMP7qZAoT
XUDKz33Du6YFh7AbkMEnGTyKaSzLMQciGnPYh62Ft+lXYCHGhsGWiCd/pBD8oFnJ
+Z10uFIQcCdruIpvfozgXetNTzP9gCQgIq4HXgm3QBN4uzm9hd1hdNbPLi4m84gX
00ipq22onRGAaHxe0nATQ5lq19IEk1qF7vAmbNfk2hsiFfP/H+9MzDYFM3j/EQ9E
99DS8n2+CttO4CNtJWr8J1zK4VLX3GW2IP4mkpjpm6mhMyDtSDuxgUwtHVJPzi1a
g82GNmIk9F6U12J5FuGHonLtpohHCrpwsYcRg9INa7rH9QsxIw74JxmPc89ygaPP
dATjMvuvsU92bwy0ezuirAByBn+F4iZ+D3vEkdbi/V95T1ruidrlkKjZ7eV8nsf4
rlmF65rIGiN+7UYJ5f5RqhrrMuD/kMmfct1ATLOQuh0TYvOZMIBAHvJ1a1xr41V4
Zf26UCimk1Y4BSZi9zCE1eqPQNyc0N9meCxLJJe0zGgLj5ZgVR+UiUzj4Z+dXrg+
xl/+7yDLDybUP/bWvYzNPl9dGqxcajTo/nTJkZM39+3OKpbQWYpo2ZKcSPvCynMC
+KevEaypOmsQLydngwgG7x76bmUPJzp8h1rbUL7ONBOlNkdOucdeDQNnKNPoBnlz
joDt38y0IC/dvlxFKkcu7KC+0tTVaz5iIKtxewO2e54AQh9SeUV+mclOGBnTo0/5
m/EywxeLVSxgg0UxRivFW7XfB//1e9hUhwbeTboG8ohSiTvNm4K1EFhcSX2HgxBE
k6ZBuNxCDoeeEJ3ekZtHM21c2rF3SCDlEFmZ77TrbcIPm1Wf3PwuziIy2oWrPW7z
MLgisesrwc/7zvZDj/fcINzw7Wp9LtJ/8o4vlyZZB72jA/9aShqWy6QF7GfYMs2j
eUdTMbwaIauj1E+1f5FTvPZI6vw+yMQQ47tLxZHgPb299SWyhl87wZv+WRFdgsnX
rAL599ebGMKNlO+k6bzYz754wRZfrUa07zj65uPxdlBiys4CUPhaRt5m+5iVisDY
cVC6N198k2sVqSbE39h01uq/Ss0H0SwSgHvTddZSOQ7n8PNWwTZB5QPHJejQ5Uis
Zpyro618dXzS/SyWb9XYcxlg4orGyxQxzJsf9x+cOZANnr1B59X8R/tFPhagIEt2
ceinXgmV6jmpRRIHa0vlnmG2UxflRzjRGKu8FspEgBPly2oHxzxQdUHREM94QizG
oVMRUbC7mMfLXjkMkjFkthL9zJOL8G/L7xibkFdwvIe2I9hxTPQFhHYrp2FtYgFX
d7a1+xBIE84YzyIN6km24AyB6Ycm40KxnVPgI/p5Js9gmWfC49MVGbj5rlCapWDr
X+3OKqLveUpnjPceBtPceWf4G2rWfErJDBVJb8D+pHjKZlI+apbwOxCm0DFhRDAY
5Y+mjWGr/QO/l9528+xY1SH3cDmoaEIYQoFfL++qZ3B10aa7P7gxAiY9/73uSFik
QNBLdwA3uufgjPBz8sIrcbDS4+KV3Z9rgoTv/7skeKLhYSwA+WuJ37UqyiN0EXX1
0VFJ6YWKS6LsHRrlCfXXOCUj9u//6cyhZqqG3QiN3RrnZr4XKyPjXRhyXN/Ln4pF
iWae1MhcFNx+gUGjwocwb0Z88saShSExC0dlyeINWq3dp0DPEaEBQCqT8NdiPY3P
uR7WlHB2WQ7aDizZCdNKw6segM/TsDCzC8K9B/E8FzOOwNPv6Y1GpLGel7qMJbb1
5MCQrP0kD6weI+k//ULPVh8jMHWcnCjvCMv9laAMj6YJouL+2pNTqxJChizL2V5A
K+5siU+Bn3Bdd+fz4ra4NNjNDhkUndNBT26q7D32av4cZnKkrcSU6Emu4H7Fhn5x
AHkCEutHGK84NZtuy40twlPZgqM7ffl9mNgzuWosyd0CK+qVcCUSz+bFNZzCmni9
gm+lvj3o9yWNFyowHnXXRBcmx+raFcfEzYEJMsegomoAAqTgixngr9OGK+TAVdbI
/j5GMmeuPd+1xBvnCHTbWirMj4e94pcMCvSwUbCM3KedGFBZjYxNqwv5Jgex++Dx
rPm3wYwfGZtCwDVdYXBoUHKNhSqoodZv7IpaeAPoMG/6QVQsspDnrZsqPvqQDMH3
nIN0OBZRl1PVQU+M0CwmVP4/jm2N09aNsrVg9l1DN3IawxY9rUfDGUCdXG9XZKbn
fgbwClskKJfp8XAOQAnZ2Lr75bPaFyzCK7QiFP/DFkGdmrO5uteqyJf6HRmIWtzO
vjuHh5Tw7EBTus0E54JhKPyZ6sPC67xeK9DgkF9Jmk0P4kpgyOm4R/jUeDZs0crT
wbErGtN6MJIU96g3p5MdAgQkDjvUhQt/fNYUrZ1Sq9yzbomrkGhctfZGDXggzcqi
PVvKmAtBXZjBJxagIccWZQPAk1K2P4DHq00nTEWDY6y9LTGTJ2QkSaks7QJIRvL3
BP0YFgYriLb4Nf3m/gDuMcyYJYMClxjJXfUlbRnWztjsaXIg2KCMjfjAVA2nqzQ3
TowGA2Krkds8OujYXK8ZphV80AC8kPgBq9D4kXQ3NVUe2aniVFaE/3Iert5tHXV4
ZP8kEPIuc+VoWi9edwbeKXNszDQqoJtIRHMKlmHiWVKuB/ZTGCGZ20uTHPQUEkzl
XfEiCUaMl31guEUV6pq+xnZkO/J7ykXbOAGgzXW/a/Q6ucNrA+vdimTpdPRKRnmO
NNHntM4rw7lBewgxYXKFEqu/ZnHMn8qzA44Q+QWN82mCvyJX2HxVj8/ROsMgYodG
NsvOv/RmZaiKECyYy22AyAFpi1bmYhD3lI4adsrWwJVFP5J2yBZ3mFqlTRegzmuG
FtkqTGqxW5dPfGDtmmw1EvltSYVehH1idoXVkwUSFYYUd41ORngL1ZgEKtFoP4Ll
Ss2xvLXPHpTVt74LJ1rP16FPH3lx9BC2NpzIS4Kgg5W+TYJAPdsD3dhmqQMXJzha
k7q8hiifjPZeowPGJoITs5ItxCwKooxpqr4b3X980QeoBm/+DltlA0f79y7LYUzI
5OfYNkusAqMqDd9Xp1aqUbyQEyX5pW74JsXNfHBaYkZ0bVJ7mGEgFIjpmbaTaFzF
2om66eaAusvHZEr5VtZkRFJvq4zsrykoQ9S1lJiT7UQIcHaSlU6AE9cciIwjcHMu
Fon2/GBZuJg1RlgG0+o/zg8piTBWa/+PXxFc6njJHj8ag3AzwhY6DMef6pUvE8H3
R5estmLfbAdAjyEv8ntV6FjYYFHeN+ffSOmy9rZpTPCbIb4LcFXuf5u840tcVvnT
oMSlp5pJu/+H48oWjZ0SCiajyaYE1XmmWhBQNC3ARSh4BuzAxjFrRvIhncAt71rs
XCNlnZrkk02K1iLJt5BrC/y9L/BEJN8dU+whZiKGN6+ANExQ45ElX5TEZKLGHAdr
Ocj+thV3WRKwukv6/SL2vtkh2wmr4lPCkEIUcLTTrTRgUFlHwCLO+EBisBdYan1V
OM6BLjSjjPH/gEn1Q1sw4E6YYfhJTRywjkMRKuuZXAMWeomP2mGVZntS6hldRK2h
EfkwBIgiTxMkEN1l8LoLP2Ou4MnWfFqLiCR6DDIwGNafiT4hdJHLakZEIB/Gc7SQ
VPvONqVq4TIng8NhxBL7phOZ8XACdRls4nsIUMo32X13gmRIH0lMYQXpZKxNqjOw
8oJyMmg7rydMU6yQE7R/HWqu2IqB/TA8JTbDP6oaxqRohzFhkQo+U6dOVN+qpV2q
X+Y6ZxloiP5EUVVJpd1U6b5bQ86/saZXDO0H+JbIt+trtQ/nrU9DYhiThIE+eI/A
gPQrULuwUEIlT/27IVld4EdlcPxu0skJUUUm2rP/+oZqXkt33/9Hph+wN87xgkt1
8v4cph3m8icHh9ce/ilZbWsEIRloLIsJlt5gj8va1TBYOPujcvhZum2ZG7lgxHqI
7DlP8Z4Gq699mFrdOyRXhH7jdjF0ziBp4meFqlqLk6RUn8iVlkJHFXBDPPRlvJSi
zyDcilfovkElafWe+sdwq+ce8vUI4V2FakSfAZnQGSGW/dEJOUb5SukDL2uqvKV8
S/wz4kxWhipUyhs+QWZeLy2LwgUbaTJjWI0Hh0JlOHZrv650VvklGDz+r722iiYr
t1Elno851yc1WAHJ2SswJDCfITQSV/lNUcyDdsoPZo3MSqabZ6slQ+7y9X/IyC8w
7SOPBziNCyS4gjtk+WZ2O4uOzR4hIiEKJaNAgia+Kx2wgUNb7fmlq3+YJqvq8+qz
7uYupME0SfU0zizeQ+FtlaMFTwO9X5XdIeYHSy1IGKT9tGi99sbuSn2e62AM1J0K
X88OL5PCIjodil5fs0no6qnNwPC2Pq4yn+SbgtiHcz0VWL06HIbAnH7nwnnFOR8G
D/EVbnKBTto/F1oKPYwrXXw5YS9O1d3j4cR8RGVcP+KMO6Pe1mltM3X3BCgWPntH
j8ceuAC5KEz/ft4yglsVOIJozNFWWhE6mCoEz7uIJqnxU2FQ7k2mzrK8I+0ta6NZ
efD/jJ6gyUQARsoLf/UtPJDTIJEjce6t0o+gP8qSJdjMIOD1k4chHx4K6c8BJ8zf
B+c5h/8ZHhrlpx5M3ZdsNpTgPPvpD8LI/BPdTAuMr4F25vf8kMRg9Y2s/Cp+Akzi
I418i+4g8b1IDV0ef5+wP8FH/HG6q4Iu6ppEKcl9ONbKxZPtgtW8M892yMuxcEhm
EXiiNw8ITXXUIDwTb+h2p2Sp5S8/T9QIvioQXJ8NHvI1Fq6XBcv0VzeBKyvBgOQb
gOypbxUazIX6T5xrfc+sLDhLtdlkHB0kJdiOPd3rvd3yIAGd+O2XRBuVzY3kaN2k
7kLhGaqFyTYRaNo4tbRK3dXH7ncywerBtdHZoKnkgOMW3YWLuad3ZxTX507bMdPs
ACxlzy5OxdDUPCGOKVE5zFpAbbaBvHPDG4Y4CvkM7H3aVNd4CWsh7Ld3xhj0QWCg
khRguDBBH1mCtk+ew2K+sIor9UcC59nJ32dnDgOMXqpjgttUlOx+aZTapu6nT4+w
zCtKTpUaZ0ZMoeOiblFy4dJvZtcNHGsbRVat/qZs2j9O8dHsf2GzOZpehn0d9fz/
uFxJcB/MWeqmjEUMlXmKiR8hF71QceJVyJv+QFR04eihXKqSBKsnbZ0D9zv76sXM
a5+TTSFtg0PUSOFFg+N2FvhNz/KvMj751HTtMKjhMxTe3Gz0T6qVJflOJS1kQd19
LLT5WYKXkDOV7BVFK3Ga1jRdDUmliHRa5B7E9+PxP25/jB7bamYZxyyONRqsTi44
9u8Iy+OI6zIfvkXKV1c6ot/vqlHEeK9FpLyjcwNzpTNQpMSSysKm3WQltxYABddT
OtPQBxi5rog7mbVW6Vqv67HYmYkqX1TNDn0VPT0rkBAsqAMclxZ/TSx2cvqwhLrr
KQw3XYrmGIf216ji05Aw7lEbRxGoyaV8DqB1jjv6RKljW+2jqsMjCyO12tqg7k7x
mCoE3NLdaRlLZ0kri9DO/iEAKAZa9Y6DdOq7AhmeWGs2f770WHywFxtxirMEg6Cq
KAZer407OjyQJefPsRJBAJHWDPp8igVNl8PzQQCvaiUjyedSpfGqhfcZmSM+Dvhb
9AclKEhXQYjglZPseZLCKaxat0iexF4/Gtf7/JezIlzAkFTBUNwZ7Vtzbt8Wxdl5
0wXwPCK5WsW5E6uZAqYpeN5BoncdSsoa1xxlupEeUEPr2nArVRmbrtLJ1fKWXFY8
81EY/9lXXb8AtWSkPEKOCY5gy03dNfnbRazd1CsLO5AjTrKm8MA0g3NcKmEEh3xh
u3ImK9PORd9834LaOpSGHYakK6y3lhiLWjov0T7eSmD9H8iS2knInlaDVbOaR3MR
Y+6IkPHl1e31RdXrYCBQvoc1xAL5iwewbadDqafcQnCf1W36cmxj+OVjajfi9Vz7
Ita/1uakyqIQnkNbeXfyUUaRqRdtVI7YzxYr501TVA3ml/7eSExX0LoOjMnBTYwx
4gvfZoqchOAtY7xOOU0yzgY7JmtzL84aBD4d+OoVd5UT+qbjb8NbUDZLXNJvjDV8
0WSJtMFNTnWBWlFPnAS2LEdq9UlZoZaONrqIMHwfxp8JQezGr/IbeXH1AhtcUUF7
q5fJ4bSGHxEdkpE2zvcpcxPlTsMHQMuA1EjBDluo0W2sfVc0C4peTi5tzAKd28XV
d6woup1098WO/M1DhQSNgyltUjHrhfkIcwtqDuq6nYPNxa5PLxbao5n2YBd+naQu
zJFx5eOzCtKTctz3LuSXKeA7HEdnhDeczavKTYT1+ayI6tFqVR95yqzM7XbZwwJh
obyNJB5FXyNTcH0SU4Ok32DymglrVeBkBJWaHTkqSnY7/2VaFARnumfyi3vcnQwh
2tZfUl7HtFWKPXjEHYy+C6WrK5DFzO85VQFpsM/DXTF8nXa33VoDRBUSefyBuMaD
KEJtapf4GBRfZrsPWAMpwm5+4boPW/vP6OqIJbNt2SMHGN5xznJJq9/3cK8p9tAy
ymBT/PWurd2/7CQUDNTpMLhVREx4eCMQfEG+Y3HyNvQTMBpsDrQDnOHgztK4yHEa
96NmIqGjqqQtkezYeOh+XOOAW6qmiNJjuf4XKZUr6AZoG2aX7D6J7jUjMxcQF0Z7
0ScPc3kE0WKNIwfu1AYlNRY+QMHVwRDUQJBbQUWTKqss326RpExg1EGsFX0TYls1
lMaGvkKSodFotVqUrZN3P61DTWZlGa7LcIJpQ7394AMR9xn5P3+dTu3cJZtEZm4P
9WSWq8NZHCaALdz1QC+rNyArVL+BzfF7UajS30ujj3hklAPtC5OkfVtwMj28yk96
YyBWPnBCzej5+ZrMV1r0tXkA+6eAtwLbxYC92w075ZdDjuB0AkOE6HQYPkysb9o0
cDWmiT3ILl/39KEYlAsUeOa3F5wp0oyCpITDIjhS306MjT1Oy85M24SPxQ3Ncrzx
gQYwqYPCF5dqo4hEcp3R6xz3oe4DcRXOKre9UgXPryfB3iHd/5ONqnPeG6kdiKrq
+szRjOqfLfvLOl51+HSSQRY3jCQ4cZvyKbSmp9bEqe7a1K5xFBo4FmBqhoXhegoK
d6fXY7gYRSPsrTg54vBWu6/44005o9ws6U3QZApc+7SG87cenGwhqHgp/M6wE8Md
b1Lz00w2SJN+5qeR10MAbmN2NHw4b4NbH/Vx4NP/xu/GfE6pEg6DP1HjE3BW43l9
UaKZlXlC2tlXRraL34graqXEHR+hMRqjj0maFpEdCX2URWUYkkafHhOqnpQK3sPB
K+CXQ5GTahkBQLp+/Da4QwOX2CJtIbPA4IneVWtjUoPbJcKpmyJikVLrS9BAyTOK
3+yIOrBxb6iW31w6flqC+IugHztZgPj5X0eYKRIhCeCEN/2K3OiwA9sNqOkrKaic
bh7ExjhhJYYi6IA+41w940m3mEz7TBxp3JomqfjDiMxdc7tXkJ7DPGKoz27s//TR
pM1bAWcLfzZET8GQjp06m5dikgb2yeOwQ6tbXtIew4XQ1QuNzVvFsF4shcV7tYUV
G8VFFLyr3+VvyVCGlSmZRQdsyifcOScxVFeJ0Pe067Jgq1/2s1R8m+HNv4NhvP5g
hRcIdL69+UUMIUBSlem/qccXyHjQftfFkg60yLYpwVqsnJrZ5UgbSdmn4qdM1rff
I7PPdiBshZLHhNqmFMPvpGLoKa/7GBYTRjaCSKNr2BBwl7CBslWhf7amZuSk0g1a
zjA54jxpYpAbX31F1HAg3ASKzhs/dH9Qs58vmfdO64gakjzl606zG3i0DYtY06jT
82LPrrOW/bL1bgE0ULyPxHcWHvh1NNa4yCfUonMjDQp6R+kIyR9gEQmKTySCiQPB
ofqTDFmAn+qwpTH5trR5YOSgDwdUBMDoptaIdMhgD9eWCVhAS2s4623Atx6pPWa/
ox3PidxG40tlamhmwFu/8hxd7PoSBT9Jx0a2lZzIKHoyfXrMoWQf4skHuovW9C3e
HWFsdY2OuSImwdGzBewfbYqNoljLL3KVpIEtdcJ+UopEL+V7gLPe6UuSNow43+KS
qXlI1jM5k4l3THPd/v2ETsGeEB36AHaGpHGBWMAGWf9KSE0kGQytKA77qJ0EbwXG
5MBWHChUAsJr78CqbN2UM8J8IU2vY2XOSoniGoTQlb7xm+mNthoipOj0nJpxOjEA
40gZlIGZzkuyQbAzqhlKc4M73OkqlzBQsvbFjn0UNUoJ+kfblhvODjCBS48nAWKe
/qV1TsAT4YyhbRsq8KZM1MMVhlsWoeFv/T9jc6FR8myPzSvUDiEffC1toUumjttm
IEYbzKHj0Nw49aT6DH9gHLPVVLrd1Q2N0Yfvqsl016TQa+x0qpXi9foP+Vz7a7/O
eqaR9jd60XFbeWKg6XMiVR2CDsi0PiSXIpsjeBZpCGgpZ813kjRNKl57uK3LiPOi
OQ+x5gBv7lEsKNfSRp8GdwGzyJfgpNtQnyFOOvWnakIstyigpXzU2bKH22U0jfj/
8jBtd+Kjd/5onk+KTrpVBBRvLec0p6ZKHakk/DcmbMtflOiiZPHJJZvrNK0H6Ax1
hA4ko0nV78TC/8uUPUDxz8ncVF+eF3GxHUlkE/PA/7eVJIXWb8lRxevEQuIAxtNW
5wF1AkVihPFc4iOlrv2E3cgzIMMDkh//jWLkmLqvc8fCA+h74aXRba1XTm84vr1Y
J+p64I+ecyGpgMP+6yHBPwPGYIDusvahZYJlfRWFqIbJTk9W86K5x8vW5rbKhyhl
q+g0FQHoAzwS7tF5L6nC7UwSMVdA61Odc6M6yr1/1qYmanKFk2CbtuDmwpqgYtiP
SaSePaRU3jOvNnj8u/y0VojshX2pG3E+SWCDAk2sJAw/EANcaBkGZLYKfVqA/U+m
41t5/YZ0N4WE0S9ChL/CN+Meh4A/cltraCar8xrew2B2eey3H+5hkPOYZ65RLsUj
eMxQHs2R0HxW5Uo7zEdvQKmYd5CMRrOIyyHsEvhB87aQvO+2yVyndtrqXSyQdNGk
XRX9pq5Fp8rFJxj3IP1+eglL2QNXI9BEBU4SYplGu1vZp7rXWluvczgkv9tle4Zt
zK4b1xvmmqJhhvftIP41yxDPhnjIuCj9gLu1mzoFZUdxHbEH/By6jp0gghq8FnM1
pwLtC4WZOVbNuBduGdRPrK8lVtiK8a47o9vmGE+yUtQeM5nrBj8a6qQW4Ke0bU0r
BsASa5wGY+MdHlvfrqQoz2VmntBxqQ0qvIpNNOcZYE7E9gjJwfGqaYHY3IIIpwR6
B5yzpXFNrvPX7DBt3TGWRMfUDni7f20d6eSn7+10IUeDAyIczw0JyXyZANvKp8yH
VvSrquzrzXC5mIP/V4IgQ5U+GRIw9X78x2g7rLyPvxU57xUrlkfXrSaSbkwB91Kj
7hwBpRbm0GKLMhqIchNsnjC8QfOmnULfcGGnASJEKN8pYfQ7r9dyX6oQirS9nSbI
LrYQIMp/d7ASdj/DPTvHzbYkXkdciLXCy4O2nzvpaQtCbnmzYxKsGLkcFZ/Ea604
vTU3xaBupKBgaPZPGdAinB9l90PSu0PSq79C/BAydxd6NiUeIli2oFiUu5hYv/gj
0IwvhrvqJLgkC+YlJAmcReGqJZHkeNFdRRwhOBEh2tMyd39vm/LHfqpvDp48V057
I/+9rRtyMKnwslS/6DC7sPRgQUJBRSTD6t03vsCVFjfWNOUCOPy7L+gU1whpJqxC
YJxiYeQGx7O2MgqeJlAYgdEz/03S8iUfC4iHrIwb3Utga33+UsB80d83QNrDkM6p
KNONiBasgA3kGg+911bjSyCJ4ozXxXkYkU2f9+UZAg/ikUyXAAht7X0ViHIYr00H
VbxVNq+JF0yAMurkGAel+wwlQW2AvURTT6iIecS5AepNRrd7kVIufWCN9sDyN+mH
QNmk92s3xtmpZJucXNu2E4M7EThAeQzBxQkNqY3miFA/YVrHyeLh+zuzcJ6BdsiZ
zQjAaqZBfMhn28++j3EaslxqA1kj+NcVU0g3U8J7CeX98pS37dNx13LN5/HZtdHN
8WsiAFrnRe7n4iUnzn8JdHRMKyENn4Bq5JcWEIWFJWGjOb22Ehko7xhfbN/vSVlP
2JzqRAeum1ZXsQj1evGJjEQPmNoZpqw7m4GbGt6xubMZMmr75flblhHMI0j3OAqP
EXdODXzECKgj/8ZO6lKntG0KVuygbjRVJ89uzgDRk87YZrc0hbQlgf6VAb2J1fZn
o+BLvrWFUaC3FsSnNmZCpZYtWRpPwL3kEoVVSQV2zwsiD95DkROG20/GJQDxd+5h
kC+HMU4NBgP7hwNz72QfDSlA444fod/Xj+v1weUDQ2PSQhS8DztHUxIC+kpWMbj0
jsmGPQba36YQAG5MlQZGEH2nvcrU961j5dioWm1GaGE4ugwuul6ef0uzv516Qf4r
6/2eut4q7kBm0f31rW9LDYcOYoKRBGAHeGUP34lukfe64MlHi2K3luaFQW5I46cK
r3DcmLk+ggC8q9Bci34J+ud+FG3BbfpQZ5Iv8SjNmP5mKrEz3+nrp3N15uCnhHjX
dkHe9M9kj1LjCAnW8Avsbxq0pN7z4qhc8vo9X+SdLzrocQCn8QG5MubHhYuiTQ9G
IEW7hqq4pwgqnMM2UzMxtYJGJCZtqFiTFxPKfEFh4sfR5hq1exBe/XXMODSPHaWQ
o8LN+wfSkwtL/Zvx0O2PWSd+VQezwIRzZo65kL4KdC9gFDg+xllD+E8NwsXq79tH
q3ZA9k0z+56hFacpSExNfDgodTLXY/kb67bssr3CsPon42UZ7MKbaadjyWsI/Xte
lcrCerQ0tXJksFXChOOnA6au1qeT0HkLoElFcGQrF8GhXbL2iVxdXIB0yrx9q8Li
VIvmK3wHBDM1ZXR3O5I6slqAiMlEJjsIfer6BbYMHGLxks5xD8aTaR5qfCTHZkKu
ldNXTlRjCNIJn+5C/ZP7H+qr1ZenJKYvSQBgMjGIFk0Xka7GT78HsqV5r4YkoREr
aaX5juRsTa9hEFqpEn49acitC9e1uzvtM660X9uBuqPkZokBxfLKjlLcPSpK45hq
zZBx/ajWs+gpS3u7P8mkamlmRYkt3UL/+9ouqzeUYl6L6ShzdFmv5Ciy8wDCyQBo
upqqyzDrQQRAkvpUCiuJ+WyF0Q2nGt8SF0jVBDbPjr2go9TD3b2JvdMVaYWNEJKz
Ney3RKgDjqOJ31LcJUDx2kTaWJYGS1O15IYA6UtEi8dtAgiDS19UQ828dl16Z5DW
+bmtcGKfP031yNB1QkJJmwmEbqtAdosjSY73t1LixampvbjqgqXbTfNWW+3bjgM4
F4mZvf9aaBPxQ9kf45/SIi3IffGU3pAC3lYJ3ycMim5VuTJrhdnizeDFRm9lTJ+z
8KYVwga2eRQJTCCsAfWBanEsDCn1rIT8+QHg0l1/1g7PkrWDAtdV7ama9n/1f/vz
h/9KHVe1pSXGtPlVOhGqrVSgAKOGwo3VA32VZ0Dpqyjn5t49/iwGvmx0tSAhnTND
h0+gkYN6j4UJlfqR/URIPd57U0CdxurRXbpQP62hGjeQRS78GjejfQdOVGWftwAo
DIqhKbiWj0hbVzeNzAJCvpk6g0EHk+KgLAqyylPK9QGf09+WQZX+9TI5JZSRJx1L
gZHUVCs2x6nsDRSOv+5oByRiTHV8Ml2TN37T5uo7phvKlGd4nBi6RkKHB2LdKZim
HZ2W68eyrVElnCpLXQCAlzkX1jTo4jZFY/m89sPSrMp8xDllTrPVKkGO6wgj7ibB
KB0xoEs39dS9CAUuPq8oSvGy9sDCOmm/lTFI1W6JgJSTTSqRJsAO0wXU4/aeFv3+
aYDwCMAbWp6gMTFJnbLrY8Jf8dNd2bbiBbEaGJ/RK4eraaS8jye8zp3kg/yOLrwm
XlQt7HDYiPyZJTE36ppjYwZGF70BvLR67kECWquDvkPF4WHV0BGVDKQ7Nus1B1o6
elauOexYK27y3OYu/hUYF0pMthm5pWC3Fx26iku1yI1AJor6eHc4vWUeo5t6StZc
GTZLfwapUvs0MwThB6hbu44XwdzBg4TqbLD61mvlAhLTKplFRkuVr3wwVfl5FqUB
eImDk1/encd54NttA6nPizccZ3Cj+GkC0VAXUBFjNFQWdMo0xhUcBytricl8sz7k
+v39McS+HKP1FTKZugJMTQusCL+kb7sNiIWgAfVt+VCZTriQIgip90MpBHW57pad
vJlBHjbwuOAdT71D65G66pw0LX+Lbqcfeg6jd2+217CPOqYcTcjbH2A9TNDvIjzU
mD01a7ZoSkHE4GURY9Qy10FsNyU3DXwkro6sOSujPC8Q/ik4w3zybImadYz2GUqA
1plyBmyHZFSPQsyprSVWnADEFzO2n7/mYKF1xaaLJZdRBpjzHJ/SjA1ECvlw4p14
qcE2HRmWKnQxlY4EsW1+HvWRwnqV+JjQPlQw4gD+acGbJ4k3PAzInA+fVx+JF0Pc
DQ6G3nZC1uZ4Mkz+b6Ii5rWMZQmxbcEhdXLBeKXFWCe99oa8A20aSvMIQtw2Gq64
aKzluFQRBxx5sriHajgo1U2VJf+ySpVpyzJ0OSU3h6KZSr9Ha72xG8tTCn9hRUOY
6vYhAtQhJ8m3q5SyLRmFHhPGFFvI7yElbRMeAiu9ZMgYvy4r/8S0LsyWov2IkYB1
JCeImgXuzYCqMAnOHNRC78nc0+AdMSASUSR0LQLPNmUmvwkJIbmjOElGbSSI07m/
9ArB2kV25o75t38XWEuJBvZZtw3c/+YOXzQUlOKC+ffgKnkzhADnF9skEgOvkUr0
mUiKzOw+6Gi4trjb91Y+Hk7XaDZS9dHzPLVaL9reLbBwWf3rGICuJdS48A0sVQig
Y4ZL8FMt117YYd2aO184Lmni/NFthwxVr2+1EyxlRQs41uqtchqJ35xSb9nKBhJL
ONnBfJXJiZmLXdzcgwFJRBkg/k3Euun+RAfEqOUJp5L+2t08H1KwxJkFL6oBHj/r
lrOxIm1UkrK1CddfCxTr+Nij1AFeov5mh7RTCbKzC+oE7tbRrFkK9C3hhmEB7Ud/
nt2i2BfyUXYsAax04DKhKLAYOV97UsJK12Wszi/lPzgtvk0+QUmxPjqY64th7zsL
Yo2k1zMe6ikj+kLwME0x7GCbhAJRO6Fac5kfGAvskspXS6NVtTOx+ggh78KB1oPf
wyUsCiOOp5kUV9jLRkVgvZGw1A+EziWY/BgwF+ZoXMYbHye7p1ZGMSNwFZt37Axf
NklSlyNczMgnswvIyS3J5pWkEVQQBXNUVbb6eNP8ILpgF2Z3yOLi9Vm+9trPV4HF
Wp/9fRnqBqiJ+ytvlbEO+azoV0ySLX1/kkLCYnPf+lBVPAtXXVCbI/TjaSbFMNF4
+f/mAsZpOFZcGRa/zX2qny4Dcww5HveZ5BtfxGE9jooFxbztaBRkquvLnMaRQ4KY
2ccBlIeqXyxWhaSkIccGMQdjLEUzuQ1iy3GZM3L+mOxOacooTtYzfis+uzV4EViO
/ssZxFWkWlw9D2KnvtLNnQ27K8kEhK3kZHnocLCGxgEKVWdoGs+C/xOWaxZUv/4/
zimDHPwAcr2okOg6VECbwlAAkTcHFXxuVf/cJDcGn9LWyXElYGc2z4tvtL38xE6Q
JiHwckgReydyGmucM9YGINJegNNs9u5fWTLd8zK8oNySruyaTZIUYegeUdyYe/Cp
9DM0vLPJgw5riwWRo8L0Pbm2ddbOQ04+fAHzs2gDxN2bBL5LFqwogS5YCuf2ZEhc
INUtgp4UmAXqYRgvcjfeZyBuVau1dQPbcHBArzkJgqW5yJ5NyV6cLYriJS/13667
OXEw+Vi+mGg5nl39x7tmdsRrJmcrt5QDw/IE/uLT0YYrpfyiDGZ4B15I+95u2TkM
CHHJo3T3lEY5h+M3lnvkUv6mcWH4F8GhoRz3kYC4HEw+GRrYZXSkvejS+PpBBNnw
+uWlxZ+xw6qvDy2UqEHmct1KoZtwWpgx9XTEzPEPbQdvhi0OYlFVYGv83aUwr6sW
24zPRngatot1vr0T8yHav0SWfSQO5hrAGfXPEZiyYhWe32OyXEF0uHM5D6zitPq/
BTRn0g97hxCx/uMgw1SF6kGVC7StS2mgB9I2qxPCAv5SXYBslCTtdMVALvo/hir4
hCUynghR1qGJu3XJgMDlXYJBftcS6RI3gSKYSxkI/znBg0iLmL2D+VFHOskNZETE
iRoARDbTDur4cjcCxeVSMdM6pd9Ig87zcSM3fBD+MXeBomQk29rGxOucipOHVZRC
/x4clgrLEWNjZwtR8/kpy6E3nqfbuQLgx0tAhvAQiR4bTr3PHy0ZTh7tg6ZFOtDm
ChXZVpoyNOaa20HoLOMu6rKQjnYZ50rnkftVYfCVTA33i2XhfDtwveOvZVj+aG7c
xzRhMVlM3z3nH78ZUL7HCccRkVg8D7BkMuyuyNRq1vmgeyzC5vDino2g/kJAvjj0
DRml71XF0XsQ1mY5XQBiJZ9djWpD8Ey85cmh2rYc7QL0pRE3Qyz3toTU8o9eptAG
XAilXSmn5Lb+fTBQC/78hgpyYX1pPTGnSaeWnuhIfpdau+M0nLY3iJDBXX4beDOL
08VtR3foSkgfocVSUs0jdda2JC0UEHTOGJackK2nFlOHc02mG1ZENazzLi5MuGOz
lvNe94z6YtXz2QuXoedRcT8Ep9ICOjRBYQDG4ThQNovilL35ZmalEFYyzoRdxUaU
8Ul82qRvlYAEoMO2B0SJM1neJVOgPtHOfjeWQKcVhSK8sPdAC8EQoIkfwOhcoLyf
tT2VhIndHHhY7cbi2GNUwHhdiKClgAnVZUUQlyPmGTNYxZjGjgqWQtS1yVM2n4sY
NTR37fNtCPGkTnLZ4Msv+mPElo31PA7wbSPNmk9ogTHZ8jECGR/yIMBQh+ft1uqh
cZduGJZ7ARAvEmLO3tUjcBgw/IoKZJ1DWJpUt4eI4rKILARAYIawPqLp/ZVFgJJf
EApEbYJzqA2vCsXeWml+whISlSgkKquLNkQbX4gRNiXCgY5TUoX/MyIbkFz1+VD7
Ry8XrIfPDkokWqqqkWt0kA5Xx19aFH5Ja9UIM5vK6DfycLTHsD/aNqPng1/qWEqI
k0wgUhUC7Xw3aoXAKLKHvjJ7+N9eUiRPtg83WrALOpWegQwrsG2fI8vEM6RiHYN2
DhQTkEjblY+K2iChY6aPVhAy2w4PVMG6LPErOUTe3liZ78CEjDCBX4zu+Ao6xByq
SXUJHtB+14AZIh60v4Shx3/UgUzcl61/kRKCIDl4rP1pC0QW7VMDULvQ3v75e4z1
TSiZhYamqKo8yIMtLGo469tA/sd3JwVG4J65BApKWHTyiHP9Du5CSDCgEUO9/v4t
NboPkwbJLB2mhHBLcL5wZ78Ejp5732bVi8dvLxV8is1AOOcBI9bWgXTf2xsM+ZGs
JqJq5vUVcTVGz+bwvC9UDfMny7yMvh5E2xBOUNKzQb/eCz4Bc0NZesWdkO8mYAiT
Kj/A651WjYxgOBxxcZL//zj9J2Cic/KDITjvER5dLWO3Uxs3cKEC6/yc6niIfLr4
yAh4MsBQePRKmmedUPKIeD3YSg4q6rkAVkARqJkkQeCG/Zj+vDZWCXrsl6B3LaUn
rYvIVp3yvuFsky2DLSeRydnxXkUzugSgdmozAxs+Dvhzg/RvvYrkS+gBugW846Yg
6ciJDTbfaC6pmwAwYtodCsluXzhjscs9yGEBE9Yh7KkJR3isAcIOednSOYnPwShn
UniXD8G28F6FkOhWaqbAJ1GN0cz/hdPxB/R+aSo0OabdaWzXrJ9fvMmHMocCkoe6
RBOU9H1nFhrmb+D57Au7d0evHbXfARN7IbanM0aN9BBuLNRM6RjriCfcJ6KCCctL
+i7IPm2GVusjllyc9opGa4btMX9Ti9DkbIn1IDNWGXpYgwHhDR3C4KUYR0ghtgMO
A830po6kdvWOCqnKbJ7oU8JP3oCodHsGE0+dAWJXvRbvFZqGs0MbYcm61WFoJzON
vIq8qlF9MZQDXDCtxPVDO/8sxFGEx1ECQLo3fYDBc2ATkwRoCyOJRJIHaJWksQju
EpFiS2sj1enlf2j0s1vvjaOlmnSpvS7qNa+Aa6Hh+wJ0DPevUspdbemOy+Er2M8x
+C4ScsIZu3s4qi4GfLs+8nrB+6Ik+k47PPOPVumjFfac+JYOagsJoyDf1tZb7n57
O2SwKkhDO8aX3uvuqbpc6HF0xHWbTaZgRqKxqrI4bNDaJKa/AhG0sJKDLZC5qdZu
qC/xlCs8NUfs90IiiNXURQcdTYY1HRZ8ftPoCdN5Mv44UmmHSo0vCvWQyLIMotQE
PM3XFCR41KwKFZY0ERZZbx5SLZkgOyjpraAQH/3+2Y+k7dhw7Evp0pbTu6wrhcEO
x5YGyZ24ql9TTPyPLTB3GDjZo0LYuCGkXBB/ZExldrbkyaRTeqlgQBe6mJ/gByLe
hSEB9+RDmNbWTllzT+TbGlULyGVgdvonXPsTa3AGf+G5Ui4vSjEr4ODXs/2O5HTM
KLqPz7Ns2aynG21PI8MJkqnynOGB4zjTpYaitEIi8dAAQU2idbiONnyyQGKwBQso
doPV6Mx1nWq70Z+pRbwNuGmiL1GNnH8x3BrpnX66f2RFX6LY7fWpd5hyrs4xg1Gg
A2rofLWpuYC06CDrr2m8QWViEh61ykfdlcYwuh9+J0nzbibDh1JnLyc/qrAuDWOl
UNke55V1JGHVu9uM26GYsntx2hthL37tRTSrFbKIokLGLJGYVoF9YsNOzFt08o5S
GIIwGK+FpUXcAo4B4jwt1YujxM7v0UCLqnNJPgj+hQ0Y3Bjb+5HVJFD1/rl+fu4Y
MCVy7fiTe/g+MyvJgmT9hFnIDs/eYRE2MbpBthJ/8gWj4DJvh+sjIEFSiWDNTuMP
1bUOF0O5YrASjF3Ok5ocmMIyq/HLTdSReAANQP8oZkNInc5BhgMQ/Ul9n6eomG4N
70YfvoO4rYPGcUAqlhMrXGhiZ3fn2Nmo36J+SPgyY87n/CfLs/QLsh/LLnwQNJJd
zKNpJ5kc14zno570JVh4GSaoXSqUf95DlQASp96goQkhncSqbbDZ8nUPloZbSnr9
jfiglgzTlSPxvhEuDL0znzWI6zsC8jYEREeYmz0sJqmGyN4/AWM97PtF783zaCD5
fApsylPzBjER/diEqgFxbu6QLeQPCqsFYT6QW1B7lvLNIr+wrUSLAYB4f7rVJS+t
p9YNdWPCW7oX3G6qUQjkLRoMdDNy6CEuSXgaM8ZPJL+Qg360wspRnA2Eg0g0991E
p2t7ggf7byr1ej+qxhs1BLouBAr6+7Lvfc0OOLBzujfrIcU8bf4ATDLcbpEKrUPL
hDJqnf7kD70QwxfZU9jShW0fh5eCaCs77M5QFvHRpubdhbgT7AuZtQmL+8nw1eGv
yz6tSNy/FSGW2il+3fOIPTvakBSSnTkKAkrOJX3dpe6RoguXPM2QS0PEffGw/oL5
njMbt4sYXHAZSiMUUUp87BZwJMq9cRTystUJx0vJuEcyropLUYFmczOQ16CMrnhs
KygkFta699fhKzUZ+D8LsYSDu3FsIk6R1Z6LPCDmDO5r/p2YLba4+D5FJVYGrZbW
OcPx23fhJNMRTNHwqCndQjEhpsiFm7qvNnP3HxBBKQ4HkLdJbKAR2IHHJv12RlJN
U0uIzYrJybcWeEkErb8yxf45eip6oE4LnV5NIptUc+kIVTfSTJbq7d2qerES2VXj
v8EtOXleo7hWWeQ28B/ppw==
`protect END_PROTECTED
