`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOJKx5WWY7Pnym+sysr94WYr/HhvVnbyD+ozmqb41wYn
GQS66+rv5ZUHo7Nk1D49F5ciSeYT/AbcmU4Ep7iPOqTk/VehPfgWNNT6PQ7R4H2x
yx7VQGD1m8ar5tl2zMldQvyKVgkWY7ubVOgSRn+zWArqbYDdK6YSPSyA9BRY0bUg
TxQDDsajd8QrRB676bFXbOHjq8qFyyXTx8kaSqyAukF+AQPpVX2fum6FXWpCZXy9
HRMYR1zJ4rtFBONMJlGqUlLWrx1m5JSKtpoWHBxl9dKmxh2Rxa3dgefTuWG/z5+y
cBdgsDXCFMvddhuVSVqSej86UbYFGl5kFbaVJZwa+xDW9iRaH48/v5mqWCPExk9j
`protect END_PROTECTED
