`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMCOZI0GvMqy/hUABqSLIJfd7o00BFpb/qc7lQnTWvzQ
8fS//0kJVaaMu09nYe7DdM4nlesb2y98ICdIAPwY4Rx+S8czc7ROu84Y8rVkjqgM
1Jsg0ZFrJVkIeTisxuBXpxYNdE2S+8O1+arf49di9wI0LGBVsUuy2NOF7L2oC0Cj
kCj6yTuTnBlCWFZ3IE5IQQ==
`protect END_PROTECTED
