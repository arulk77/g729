`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41lmq+zstvvtk63CZV4oDOWUZsMY/fwNYaDP4YXr2kG9
MOPpS95CMYuVU7p8Yi/w87tlV/xlTXdVFamKAQB+WJ/S7kXYLl9gmmYiR/0SNGgB
of46gcGzXBDPO8+BHQyIa5/WGNpMnh6kRRDsjX9bAkJHOc7TpvN2F6JLxaUCquf6
sWRh6P8kMPu5XRryEGOghQvcBeCTtCGFw9xl9nS0WAhkpSNXD2YVC/DCIIr/SVoo
vzu0xSSdCZ1+7tX+S8NbAuZ0qIi49EANwUopEViorRgvX+45GHV7yRFeI15bPjOU
6aKjutycLK7XnNshQMTp6CCU2iovOQ9iYRcQRFPHvcNuj6lQe6UJf6uStUno3D/+
uyLD876iidrohpvh+/zSx3m0NfYq8fqTbQSIjikfMrfogguIgmMQhcK6PRWP5q8d
JlATQPisoZuH6/OskHi5OA==
`protect END_PROTECTED
