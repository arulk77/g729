`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGlsGU19gyylcVDDerr6pv97T1CL1482qxAng8gFq1kX
Q9C3NOWSKgu6rBiNbU+/u+iajqqFq7LNmz/p3uLrGEu8MJCGh0ye9GBlHpM16gOw
r3T057SwT+9O4WBFgbcrSJal8LXOUXwLsFAX3PccurraJSdyvf3IcW3PShePB5+x
y8aaeER2oyE8A+bKshnrZQ==
`protect END_PROTECTED
