`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHICjC0P/IV5fvhHZS4AJyZOUo3fmUEUgx+/vWT37CUg
3xlqoFZWfP8ZmAyFvvxSiHngjopOdB+rP5ljGo/0eBvk8wPnNog+uFF/bBGbOhrD
/U6BLw+3X5XUgn6buloPlrxAxPd274cmB/RwOzzjvPxLz7paT2EvMA4DNrYMMCqB
szM1sP69xTfDjMdHKzJ+Kot+t0r20KNqlFGD6ZX4IplThF9kDBUfDJigtzjsEfth
`protect END_PROTECTED
