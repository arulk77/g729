`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL86PnUjo8/XckcM9oDd2UQolBZrsfFgN6Iu9PufaewlJK
PgQLAVlk5UcFhIqv2NTnOsmr9fnCE2FolIWmJLfifkpaY1VOQ2FH82j+hvyms9g2
bkJFisRr1+PJ1kQclYMFptfSKPVYry+Rh/9eJFarS3peBzeAmPBFQ5sypaSZhltC
OyVd1bumppFGPKuN/kJvToNYkJu4z7CJr/vM/7RGjCMp+s1Cukwj7R2qZNcTz+nY
1050NgSpku2kMDkMrK1eNiGu2TyLw+1Pn5TJLAL1eszLNOHWqVJRHkwXwqOgMaIW
Dl5+9AYY/pU0VfX9RzKNp9hQI+GyjEeQqB3XI9TkUE5nJa1aTgJ/gUYbiZVrx06/
U1Igv1fNHI5tpdqR0GR3TlgAIIJeUrlwxHkHLKQFgfO8WjNTf2oEeLYMnFZ/02WS
c2dW1bii0Qdb+M0H74SqvDgHntNU+7vZ4OxeGZZfvi8fqG4WPu9izf5WtZ669juT
Yskk1Btsk+lCV0vedGtjb71OqswEHnaI9UPtjZZ6IqhE9VppWA8lVtD3dith1oKq
2n0sdYQImg5n3Em+Srl/Za9a9FoCFyWUYkBvGknLGtVprHGDkubF9PqXYyjF5m/6
JNE8TLu9LWTRxcVxYK4acAZBpRJOkxQG5JgV2xynSWo+LlUVfNtu1Wkg/I6OuK0D
JZyffrONgpWuEP+Jt0F5o/MX4uWFvQCGdDnZHvYN4sAROLqkbRgYji39Pu6Qb8a6
2Gr1UgeAvfajTEL6k1XLItB1Nlqud7xZhXXsjFQhSrlLd0v76UQseQhk6Q7K4KaB
AM33MPRoCKPu5t9MzJEIIw==
`protect END_PROTECTED
