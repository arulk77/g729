`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wEb5x3ZFs2lL9SLSvM5L45sbTUQCSd3Vz0g7msHgW3G
ERGVF+lLHgML38yHJgK3KMIVPQUEwKg1SGy7enieWRMZyY1yNyZsBvjK+Uh8VAFa
41TVFMIfsJNEdsW9FvuZBkfANoHVZ+333dztLrKzvg8c4Z9bvwsNUB0bexcaCg6p
aTMawlC/frtosbmrYpEXbI4zDouPp3SqgXPu6yLAU0d/WokcVRGg/SeytksxeYEB
PFQSmo9/zzx6ZEYNruqKY/4SF0c1/gVd2Jt/4mkRG6eneBGm04Rfbt871m3PkQTP
KyZgdbDk3j8cGPyNJDM4GbRN48yP6fb5FOFYgtfOcE3an50j2wl5M7tsUrW+suAU
Jzt4WbPGja1Og0+wAj52vg==
`protect END_PROTECTED
