`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOGqzYrpEDHvapwcv+9webHadqy1gynyx04havr2NhDR
Cw0pZTx9Wi1H4fX9HreVpTCm+B3pc2MJsH5CrucHcumPMzvDSo70oYdYTGLLUq8M
46iHSDD7gd4dh338AnKV0Mhy+G4AigiOlaHrQ1Voukf3cMKXqhhgZ8sfRiUadl7v
eu/ldlrXlkskcuiv+qHPymmqvYbh0rsq02iy33WSkp/0z/MQElf0BL2F5b6zPtwP
QQWAkKNIBPs/ndiOlxJUl3zogimbeIT/w7eg2AicLNgAfQVBCZkk5VLi/dE3e4C7
pwvjcGW81XurgFV4hwVLRmtUBlL2xhXL+X9UrBbbBX/ysQj0xayCJi0ESjp+uXzG
LYpquxqDx5o035YZeNSnw4SO0eYmBfGm8wl/Lzr4pPcUkkzreCWdXZQidNBG/azZ
RjTaEp+yF9TBwUVBypS2o0aCdoAZlAe4ClYuIkQHo+IQDJFtXAKIQb+CFqzu6jQ1
pYeQMokbI+TH1KsqICtveuepTqsRU3cwP1dsb5b73EStBNX1A+vUGaz6W0+zCfto
1v3cdZ/AsVsjws0P4iav6/Xg1+9+Wv/gSsoZLs8Tjp/JaBeDp15g/hcPLus07F1u
9gczERz7zQZU+iRl8Rq7YXRJZCtl42KRBS34ZJK5e8GYp8bFVYerrYr5T4SBkcnn
`protect END_PROTECTED
