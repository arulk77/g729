`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDClgg7mzi5cmjTMOa61jh+mTu/a2CBc0gY2bHCAaqsV
PcGQ/f+dfffvwKxvNCYbBIdnsESOYjNHMUc8sGAsfbI2bT1tgQLW7sslbjX1STT3
yLigt8jlcYpWJWg1P5i8qcEnnNd3jpEJzqK5l/UIRAiQR7dCtlna47o1DviGUB0E
SYmx325mjH4lPVuiyGkfhd676KLZYRJp6bBHIXeUjnFk7tdvwG3g6v5yrdo29L1t
`protect END_PROTECTED
