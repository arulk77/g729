`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEPDEcIfsk4o5YkyqUfwLtpT4lDAnzdwb8ouW7gCMwr0
/1cmpOusThQQzhy+tq5n9NDzjwrwY7hYF7Bfq/vcbrHpm0yKlXz4OAjDaUhrSh89
3+Wl/5thtlF5rxaaerhWNEub/s6RXxStuWXbgsYtsSwSHuiv4BZZahSbfCWLMixM
2XcDT8YMjsYAkhuw+aIKSPMl4xl0njDK1J9TL3hPCP7McnI7KWjkgZ20q6ffbLfT
9rF/C8GOaShQ7a4AoRqRcw==
`protect END_PROTECTED
