`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDASfd6muvCZBmZ83YUiuYstWXfU3E6ZQSfEECM15fzoic
QnxM60QwJT35BBejgPvIRMswt0Br9ibVF2nYmXoQ/Ifd2/svSxvbpLwDgSdrCxhn
wUKHTVz2pSsERJ92r/Gr/t3k5Y6X1J4vYFT6+ufOfVXKePtgArdgraGgwtm+Oj4m
xwt3IKREJT+ICmR0bsXC8HP141ToVCLuDIQZUMM+FyyaOEtE8cfAknw/TVjdQtcX
2UPDigmHxwOeP92c1IRMVXAuynw8RlTLNeQlOJzcFjI8Gm47UvfagFdFccM2kx1O
QMZxGEl29/lQMob3xzXZ7iZ8prshYV17yWV+UFgMUFtO32aWtPg3YETgJV6Si6eH
6NB3Vxn6WpEgqbxZEahLsupgYFLJ952RMTsv6uM1ET46RB+94CIfml4Q6BGLfATj
e9nVt5zjKi9fsozr1kGjN7KH8bbiZpraGbK9UKZDd6tfPSoI8ChzAkZhhkYluYOG
Z86XUVsgDSIrh6N/39X/H3rQ2oFA+hLl/2mKk4ZXCOQZYeEC+oAb4Ow+xXiwEP8u
r9tJCR5PVV6dLVQMLQ1buiLMtTPzL5LiIkaKVudvzxkiwjCdqP+Gx6bxddUm5D4s
xZhPvO46SXpzKduMTSQ9CiCxKD0L6f5L24xpUF7mYRU4ym+bYu4X56/UrpvfLkQP
AFbvEP4jbTd9iCSTt/H3+G+t7uU+aUCbnQJsjDjIN0WysBtwU4tlLfiPG0+k3D5p
Qr7grYLFhvMZsx/05ak85QCq4F7JngsKvU2iLx9rCk1e699G39wgbmOT9sLPy9cI
iBuHtnzVRVra/r0SU6krLIpJ+l809DEb8BtSX8COsLP23SxvRVacQ5sLziNX7WAz
8VbYWCqazQNzmuPYPdV8LQ==
`protect END_PROTECTED
