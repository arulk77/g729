`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ab3t38y2wf5+qsH/48ktMKrytsIe4bC0ISqCoGY5JZ8UEwT26TaG66+oYNSbAF4t
36CbZU/FBmFAhat6ojU5yVhEVSNzrNvz0RgBN4WPSGaA5Odd1nLcBlUxV5RoY52Y
iqkX06IAwFojqJjiA7OY9wpT68Y2rmaewHaWAbdDdTLIJxIFuI3LiYngp5YptNRo
eMfhFYp2tOwXtAQxKwlY2SdxN9lILjTGO+6fFOGPUxpTNagjQfFg3/9aoKLQa3Ig
0qe8eClyoxUGBwVu4gMUbTj1y6LKrg21syKG6a7qEdjeCi8WBr08KpjJ+dUPf/Qq
hNjDCrGnmX1krxiV5rD3mBWPswjp1/eZXJascPlNFI+sgeqf3HFjv784tj0eAMP3
u9yWpcwkyh5sMwlmEfnRKW8WBDo6lybROLBuSyHkS4I=
`protect END_PROTECTED
