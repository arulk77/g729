`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOrMcm4rNraZWQQOVwInh/EDYWSFiRj1RFKcv1ti3zov
AgiM7jiXGRJXY+msoJOxgXa2dHRlRDN70UqG8cbiovOuOX4ZlPajO/+Wo/e148B7
pd7oe9DkAJE/myBhJWuDc4rhUnDCCScGtpMO8WtBw2FpDg7JBGxD2yABZ40MvpBp
iDCMXlYDhEyscJnqaWZpVtCszCQa1RxhxlTQ2aN+cGO/dxKXN9ryrIFEXuJ55LN7
o41Dty7yA2kUPnAc7kh2iQ==
`protect END_PROTECTED
