`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SW7nHk88U12dDE48Rw9mF4kBCeesxm/Mo0K57eRTR/6W
2ZJ2oSEGrGdduJsxNCrrNSqFsdhq4x59RDfNy17WRMVkUzJIkoN3RF3NKUyIYh2s
Cl0mh4FiJmTpCy7zAZGn3jUXmkUOKWSGGTMt44oK4mzD+NCw962ILgnubFZOgoJl
`protect END_PROTECTED
