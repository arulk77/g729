`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49MOhmsSoBqZZqTyx+lnD/WKbmdyXbbbGVUXaC4iTYKj
bYI72pDl3aPACGq5WDrnz1XUXl1cFYwZ4cuk+6VPkJdUMXZVOqZm0roIkVztbih4
fH/L7e0dlkc5dtT+f+83Jd8l3UwR/vsMO22tgozNbs8=
`protect END_PROTECTED
