`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/lx99wpZgE5utV+z5BhtDvqcnAoghXW5WGhqc+6qvnm
n6aIWYouinUG0VTwkyxjMkzcNcH6daSyV/+ojR6oznq9pSusqogtxU5PLKugl7f1
+FPeMLzvKRjg+yM4HSlpyGpDyJIioIDmDybAA+BLK+gery5JZJcdtl97nz1SQiuN
ROGC0aDUk8mH1hzcwQW8MVzECuP38g6sNcoUkf3ron4+vKEYEK8eukFwkCfsXV4a
ff9yvrz/ecYZyqVJTQQLBVabH+L+UAuwMEqbzoadr9cv5Hb4miN62EaeFh8mKPcK
sg9OCj+WwZxqsUvsNcKsGuFgnxGKzfLEOZvY4HIQXPvszA9vpQqJACbFvxrBhmei
QaAbtFNwmFE+1k8uQyytZfUGKcv6UuSIakTDEq6D3Ng20hEJlrBYa8/kAxysA47O
usiP5D2YU+Cw3A/Bs34h7I9WBU6ol5vd38g4ZgNL7aZgCGOwcGLelA9IUwWsjvut
`protect END_PROTECTED
