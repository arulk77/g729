`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73CyPqi24IbCfbD/n+VM0+bk41MJsI/nUgRKWsK+TY0gnn
bKz/uCoLqJdUAX5WXeqTfXunp+H5uYRCC914VrS8u/ke3jbMjvQKKc3y56vSJH8U
7N7Vowveg2RmLUXdA/YCOiUPVrPfTB+iUyEru4lNxP4Y6tMKjNR07xejluLlGg3a
Jsyw8b+kBK2xSqBQAFvWjfWMPZjM5aptxVCZVtqvpWxw88LXZqvWPIBmJNjsDSJc
e1UezA6dhKqnsmG0sFsWkVbyi4GHC2FX6Aea85cw6B3/b2QiIzpXEFS/1RxrRN2R
iABW6fMtDX3ecv1txevqjw==
`protect END_PROTECTED
