`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46adUxbWn3vOCcltc9MWsG6LAX9I3ysxcgRYEATubVoj
9Xcs0sfXucwOsMtvV/nkzHc43AVVNMGW2pzgAom5q+p08eNmq67KpqqSEaV2hT/n
km7R7LBZmJyc1caU0PkhhsBgkLRL4gtQF5j9jv7lRP5YkuFV7Qj87E2EJLK91tO7
iuHnjDr45muWgGaGbTiKwtFgM2FMlHhPSVsk584l3M80ukgcf7tgf1JUUB91ZEpf
um5ui0Lrt+bDkjsisTCcfOmO9PefQWPIRudDG6BX5ZM=
`protect END_PROTECTED
