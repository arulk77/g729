`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
72DKe5MEZSH9IT4s+0rFcE7NjYK5fCdis9nahs3McC0nW4087j3kx2Kc8JC7giUa
PVdEnSJmaAOSKKnQReWFPyKEn5thOg77LRknxPhOS/I6W7YDhqkIHe9OtN0NFDfo
XrPICsRxCfhvtGXy6hLicSfWoVTm0Yos6/yqZKlkm+y8lzEmJaZjN9DzDBoUlC7q
6DOSqO907zD/+lSW/7euVfMFooC/s2/R75Fk5Aq7j2iRsga279wIsvBFg0ZaguXn
m/yUAnjyTGCYmQkjwP7rBPKCxSn+lc7XO+o+OwqQ7J1skc1rXVolbMd2oKDtJqtn
`protect END_PROTECTED
