`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40YZ7QtRm/or0jwgAuS1NzlKgcY9V9ry/ULRiI46TfR0
HkmDViUsCUSW7hDfk54Q3n86I5lUEg5qNbGAijmfLKqp38dpft/8EEGu3hxw0jk0
n/GsCHDjtY/JpSHKShoWo+PgqSuMx11pOnyFljGfhSIl50yBvCl6YkCuhR8iE4la
asj24YZjjnJj9CP4mb7CnR4qw+aW5W9WOsI+ddBdYMXvcQL04/I/6Xpf6CoNgErc
zdjoaZiW47YD8h3oz9oTUGNK3L8+0J8ZhnqDpz3XrBFiDCEoOYV/JoXgSln5bS/A
8qCYCVkevpMuf5T2fEgtAA==
`protect END_PROTECTED
