`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
zbNaVR9vcQVAIvjS0Qt3GUqjpUbB28LCcbjSu6f9kL6K7bVR587hf4oIuB8WhgpN
jZUG6L4NfxVku+QPnpePZYGNMxg7OBZ4uboIKpAwXbnvQ6uRX3DIDtWe6nl8v0AI
SIlFai/2cF+cIbhciPRcMgV+62wlOPo0LTIayA9OzjVbgOagJLOd1OUsxrYlvsd6
3B8XyPJRY6Y/baIAFG99YIPQRzft22Lgq9TdCd3RJMDiRuQbRgMuZhbZlQl/bmSQ
E3f4D2H/fyXqh0wT2uE75JKWYXU5z2JvMLPt0bb5RQ80F0G5ppysYVHj3sV5QbzK
i86oxjUfv4uJLyoCu8TNskMGawVC1hqkH3NtjI6jQItpSBfaJg6erGy5VuX7Hgey
al7tT191J1q+VCtXBxYEc2bARCWK55ZI9iLcYRogvj6IU8A2ixogEc67e0FjA0KS
WP1QkPjHKJlmgrq2PV8T9Q==
`protect END_PROTECTED
