`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
l5eymvnnLdY9K5G2Pcs5AP+aic/HDZsHOYMaSWlvTJfs1YiZlkWJB9/fIDiez02Q
ooJLpmdHK73A+z25UBezTj+uoPOeblhPMK3Jyr0MXPXy+i5q6/QMrRvrnAOe7S1B
64u3DSPteb5fCfWlvH/RyFjPbY/3O1EWrf8BxlV/GxwO590s2Vv2ViYuVHWUolMm
+zKgJD1ctsK3DwmGOOBzOmQ4VSNoJuRgDBAgKfilf5ts6Ak7JGgeq7GeS0ZaZMSh
iOFVACGQdzzT+t5Jdfl8vsGNtMt16PaP23Ud6pb9klRhZscwDYcqu+VByDZ28I05
S0kybjivRVdQ/vWdxXwFW+oB2SscOzmv2hJU1oznqtMsHNdQBLA/HmU8XlaGZouH
um/kiREu+IMlz1rwQcEo+/Nd339qYpBHjnBw82g3K8YFLC+OYm/4vwZSizfT2NJC
OdTCzGYvkc3rfgcnVn5pvMpURAiynNGG6SBR8jXrNtmNYGQIpPZ4cQTLOfbp6YjX
i3aTq1z8bqzFPcmFSgwLKWJe0DMAbwQRszBu9gSLD99WKRX6u0A2pXWc7f4F4StK
GJEd/j5L73IOiHVI4kvNDArG6AcAKxsXOM8YWcj4IgudQTgGylixBzFDyx5+wWQT
pNY/4ZFWakrBlYZSOaedDQBF+GO1wwJZhTp2udk8l2pcj+q7Mr+33moaT4HXPsX9
g34s2ZqAG67hdYEkgqoHIPwh5rbkktDKVCSm/LoCWpE=
`protect END_PROTECTED
