`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFl8sZ36zr5sAyaj9WJNTa4qb/1lnuT4OUW4Ck5o+9Lh
rM4UL31s9g7epYw+LGX+d74KJ0FN1rz85ELqhmj5tjnWoODOwzFBDzd+qeGPhhgi
m77N8QsOdccoFh9WUSzE5Azr9ws+71+AU4c0WYC3Xzx30NN3RuCUATflsklwiFMA
VqGnMJMgilT7BfjFigCJuJGodBoFAh7ZCy3nEhmkBAB6tGKa1jlK8eC51Uwz2Vdm
epGCMsZJrdlIEdYrQL+K7A==
`protect END_PROTECTED
