`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMJrQw/z1b1/C+bAFXw5NofEUU4c6TiqMvpijAolI3Nq
dZl8R0tdfMfXTm9Rbne6t7t0mQRIbAYm43eBgjDXg1C37tDi942c/0MXSJNjvx6c
ebdy6Y7owQtVCN6Bv1O6TsPai09A3GTllI6GWTmkhzovwzCEaBbvc9hpDjsx0JVz
BAPjWRfCg5T80Q0vI/pMpJaj+NQw7it71W5juiC2bhBrEqq2XoSwEjyNDckYfaLh
rw9XBEzWYRzHdVYkyib6cVq7B3liy6Du1WR3/FoMXAorTrDvhV5PXb9zI3arcLLI
T6l70Faq1zkYlLT4j8+S8Q==
`protect END_PROTECTED
