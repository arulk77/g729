`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveH8GiwGA3paK7mK6RFR7TNuRBNmwYEY0mEVLT4uxPe6z
AiLpWDU/5r3bwNf7cyz+kp7LXqLZJhjoFyG6NI0ZcdGneiBFB6XD7ODf1K2LQC5j
0nzxC2bhHWGAUUUYxUX3CoQWJc8MYbzx78ubUj0bCsYD+P0yMbi6Y+IDXSUTNlmd
tq463+EtB1MWACylnneSDXdMtRXPTUhynCCAvy3OVAmA4+AtbZzvIGeSjtMxn/2K
HCrMGC9eZIOVvR1XdQo6UcMCm5h6quoZ4YSdsCRTxSuatGAqluTPaS4vfK6a4prc
dMRFYsZdMMU1M+/pomHAOW/kPRZz4QOEn6QRjeiCsyQbOZtpMLGdNbHj25cazznU
yPVo6Ld0+pdXKSseT0uu1MHvagLz30+KtWelchlzBEqj+ZPtqxGJy864zK3639b6
ULSrbtpzWKkVNbibxbzc1TNZEKzLLvFYRVTgtvzibAQnWVqoDhGcFvDPV/NXki95
ZmX2izlcGjoV/TmbQZ7UUwNDHkM6bRZKk4akcZYfPz67qfsxKjvfta6V9QQkNteV
`protect END_PROTECTED
