`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
K0HxfhmGSPSX2e3D5Ay55iSyJLeP0DcIgomOgAvHFnuYIUnOS2BXHJKPbLo1sWfF
fFUI8FxHE4RP+/2pfailWsMDBnELR77p+AJR/LBOCypz4v4sH4MIBRWIr6XPg4dm
MJY1efSO17qyKjdcKUPAlhJGpdnMwg9V9fHnDv/+3S/P4zl2NaubO1Qzx7slydi1
aOw7FL6QeZY3GU5wT6lHd9Oju3EYURErZOebQMjfvxVL+26MOfZyqJO1N2K23iQA
pUUpnjJWMjJz3m4WrFy3JAqNVkZwDVAYSCvfg4SpxwUr79ISNWSbPsOF+C6KUz2j
agppePpOCu4gn65Z2grU+UzTh6XM/sD0SyTWme8/xwf05Ym+35OyQF+WBcBeL38J
L87qbJerCEJVuqIYsbN3RjI1pwo85ng6OFrSLHUo0tfc0DuU23UHJofS/MsfC9vE
MfT+u5D3A5BaJxRta28e7DJdthAn3XbxrOPuTN9Yao+KrvnwrlIrgcSTfKokA5FH
GPm6CJqvHGSn7qW5C3vatVFswxwwJVCmtjMdwUslsX0=
`protect END_PROTECTED
