`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGATEhDP7vEEVTqeM0u0ZTFwMkm91vYxxmvRoV/WLdBs
hJuLXmx8N52q6I2wWvU5+ETmkHgf0uutLyEB5pJ2xjFe/YzNEftKEBiT17nowH0L
gWNtHtc9qUvU26UGdcnVKaTezgmJZ+29OwDGuhQT/AIyJjbP34GXglPWprhsYNH5
nl5Wj239SkT9qBdUEv1Kpb96UFEDbjFqdZ5ENlPvscAoq0upyMv094+BlYcDPG5K
/La0goYzdSR7NB8R18Mpds02vkN0Vbq9/8uYcpVBSvhPhCvuowmyLT7InmpUl6pW
9ndvZJHt+8bc5mRRDTFPdA==
`protect END_PROTECTED
