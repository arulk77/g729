`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN59OFlWsGSLWJfNJ3mNZ5kEP6Hd0H9CaP/8jHiLbZlJ2
gXJiHkryfwpK3puQt11rQYGpmJb6i9ge5lEWbMldhErP6oVMgqxJA3a3gJgK1Ks8
1mQHCrQc82AOMsdTSN4XGfKabk02VjupcrTzn2ZXdGT4YeB1qJCWJcgU7DsOiBVa
zTXS++6PYIZO9AzJ1vMu9C9KQ1455e5SJd5VKfBTnJpI6WY9N++pZ+DSq0ZJX0rx
+6UrKXoiMel5bAAdOYIK+YxxKia1B0EGJmB2KLzMeQqd/y524SUEDL/FlJ/sVIft
fCrM8ngWxhoygGoC4uCCm4CYQ3LJ8xe/IChIF3+iH7UrawOJR+P39TMl5NqGJoRX
jOrQ8GQSx3Of0Cs75FavsTse22VEvq7Sxf+/XhqS6uY/8Xy+grm7+yLl8dalmL/l
OF2Sy2WoF6u/GDmqisqo8F2ieSIKAh/NQj+AgXCpIPbNTRE0cCXCgDmHcF2Bqyg0
idBsI1Nm/6ty+wa0wiGVWOGEwKyUvrV8i7aV5w3lrmwwxWJaIpobzVOxFqgNXeDP
c56tA4bjfMGR2M4BOERThWPJxrtmYvM968KY+m1rUV55L+mxbg81efUMdc0t05RJ
zDi8rrRDNB5AOM48Kb5C8Yu+xxsVer1Ca/eLo3NPZ4t9FfZ8e7xJ1JTFJzZDce/s
igDevCys7ihoeFQL/XyLT3OWFrL3vpqA8I2M3kTj0Nfc46gAK9pANF4Hh6LF0629
JsykJW+GtTcjNw0tDzwClATp4c3SweRwYS1xr49Pz+9et/tJ9Tof/sgA/bkGoc5L
8S0TV8TBLb2u9jHyjkyYvfUG3BF/RgaeYFaL+BjQVRHklPuklGYwM46QL3pJ2yhG
gdoFup2E3eqObtOtTlQb/FLZe6aSfwCGHmXgAPi+8vc4wt8PXEPlM5XYnkZVTEo2
idw4MF4X+UxVVqFJ6zPuUH95FVpx411QGWbRrgKttstrvDPV7Uh5Tguv4NBLwYD5
Q+0kIMVK9F9/5PqL7pQTphGhYBLkyc+nsWPaF6ttb+P5BWJMIG+Xf69i6OIwgudi
r5yuZ8tUHASkOfsvoX40RZEtbgQHbFZNRA6rNHBLIQuzZkFb3qI89PIq6BJ+5XVm
IXRPwYn2g/1zez3WMK5suGiBnm8dXXoFcO7W+cM25EOghxRvGDrADZ3ZFBFfn3ry
227z9suK9GQ3uxU+6L9EhYnRaNMvRDq59XhsB8fvqS3saM1YG96KsJc+kHJ9G+7j
QyacNBqqick6pjfsEVEpW3STZfvCQYNecpMfGdW7r1fcZbeZDXc0IOwIl8e67UBm
O+m/9HFAS0kqBvny0TRyhBcbNGsBtnmeo+j9okHS89NhxXi/XC22YwVgUd0jbczH
wHZuh+ulP10CNEtKSMxycRZHhh9aSXZV83qh6/EH8L8gELG+BrBaT4B7+uIxQlLF
2q81MLpBplCTWu8hwfqpZ8e2pcw3m4Z06G/p27RsGjvOg8adHnDHPxANbc8aHZgr
VmFvwOGngrcDWjafNboLKCenO2XCvcvaqJI21BiT5OhgtGDNOjnN2ueHXb6KZ9EJ
m87Kq3+wAflfsTMent6zApqIWrkoIH3dA3ZphmDpPjfvZzQdRXoVQKIcpOl+3yKc
Uf6T3gE/iOatZ73KBWGCPT//1L7QuUIE6TiihMRjExsQhC64Ifn84GZq+O4wHU5T
5I1la7DqnLDKpnmhzJUf6g==
`protect END_PROTECTED
