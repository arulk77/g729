`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Uzo3mA/mwHt5TnYI8qcNLIItoY8/YjcP2srOFf1t5Ibqv38xhGz+XyfcSlm15MAE
SQqzTvSfvFwyYR0xRjO99eBOqS1Fy2fUZwW2SfE5+o2xpQCTdY9e0aOQjcNIzqwL
+OwnV56zqglR0BznZv14CO5+mYLVO3clELy1X+sMSRP1fB2gzew5qBDdr2SssaLz
VzSS/lLj9/IBsG1LzGGh/jMuvesVltEUqDUjB8hE+CS4rrOT/WIbAudZL2Z+HYcU
0GWSho4Hlo7+TMNLINarCmDHyb3xinlZ/KfIHJM6ahvI7wm7MMt5UFDowhSEW9kk
bF/TZXCBfxVexHfDmkSx+mvq2e9Tt1oUAfbF5w2I9n82Ydz4EPbBXYueZju5Lxta
d4NcI4QvLU8crLOa3FJ90nufk4RzRxRc839v68mpXhtLedTtV8f6dlenyF4tLjno
3LORknqh9dzhNVNo+V5Aj7EQge5LTQNZ3xmNUNukHU90ib1S7jzdKFmHXlQTi/Km
u+ygjOj3eytbF4rQa6ffqdPBLOUBadKC/LNRvbmX2eC2LnrUeoh0W1QpE4dW+pS1
e+eTifyLqffH1zVXgIEILAZ/zrNXnl4vrpLNoFsD3XgNsn9F05zMIH+aHg5hE49y
MJmXWbFDgVSSHoGiDgJskac9Hc0UaM61sW7O5JPqg5375mxR0YS/FgcYJsqwPbAZ
+811qQ0hl1JDcrW+49zOuA5T+oUnroEL4IMUp4JylLbXdfWN9GVtYlsnQl7TvzD8
GCo9wys5EV5Ty/sZyinKPsMVZGLBmb/7Wuhvxtlc1HxdqOe1YSfnP3gTFrDUFY0z
0hE0+xHbty1YX7VCUzxMqXuDslmm95q6jR80Er0WQqKA2SY+wiNX68T0I3raXbEG
lR4R4/Jcx6JEQXKN+EIytqJYoe3oskNyVeQk4T9dLVvkrMmy/rGTGTYsmaQ0FxP9
VON2fxdFoBXUAKR3SMmUho8S8QN/rw/AfwQM1x3KIU8p6Bq346tIuJw0RTPjJa+y
xgZ6hK/D6vJLgIn3GO+otJ73pehlz8r18w3bxlMXcaUdzUFc+yWanCrMIQc6OTvR
2/Thrg/900/fwESznPxGCR6u572qKhG4H+8y6RLfboFWF3zQY39Kr4tmMA0Wo/nv
YrOA8WdkiYXWqHm0vKk2HSIW7Zp4HYrRccsTsis8pIS6NLvcs266KFz19DpjxLni
bLFvEm8hZ6BS1qa0PtQ7tv52vwmVRJvHj0/NVIrN3KJZmFmXeZTvF9WZ0tVjMK/V
EuAbxHRpEkSb3N5OYJI8wJDR+kjlsBsl9qzfj7/bXG6zrv7kxL+21Xc1TswA76PI
X4572/jxuNhPCF4+6X0t2oNmIoAPCSPiQUz5gK5e+Lg=
`protect END_PROTECTED
