`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ev6Ax10uWO40yuyR0lcYM2VGlLXOUQEiNU1EoEiQ6CGoGQ5lO3Uq1ab4uzUyAs3x
p9HonOGclTG1g2A+XTS2wN+qn0DKntNcbBC251GEh8FmAedlf0kM/mphV+FWEP3i
BAsaNBpXeyPW5O/bsZG8Fv8ZmFv7jQ5ESMrB9T97RH1fBzIaM/Fgath1GlNNRmUV
IvC34Zs3eJniF3MeYzndNjM13Q350P6atjnq4oKpNp0MRJ1fKnVsBpbKIQ0p48fx
bl+6BlTVj6q/uUaewz1ePNpUBpbxpkBT2v/oR/T6ceo=
`protect END_PROTECTED
