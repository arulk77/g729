`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJsFk/aYqzLiLjUoOs0rENzQ1hP6y8FR56y7ylWtxi88
sOkfVVOG1pnODrq6CrhbsjXaF2U1pBuOSi1Tp578KL6nig+0Ff398u3q9Lo639Dm
O12gQBCP6lgwvzklBe89A+B+gzmXnI3gWXfTnrwB70TORLJKZQK7xIJYKiR0W06y
FXmUVxXabR3m7DVCRIW3aH3d4TipUaVZVD4Z3zIt/n3TpiyeCFFEHTuLcqutZBd1
cpx/Da+NZXa3QKDCK8QiOw==
`protect END_PROTECTED
