`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aZzzFBPHyuyY2HHDUtUyDABo3WAtFGWurWf59NNSxLtG
+NNyciVjJg6wR3lH91r+V6uhqNItfI+grJEbHyCiqkpK+DYA1AWM6jXALr0G7xKY
STlWmqvsgoof4nn+j83Hf1dWMUyJ5Ery9eX7phYvhnIHZ4M57a4cel/YWfv6lKm9
xdKcDa65aFLlxfcw74tcoRDzAWYGU7ylIWmHM8C+GpLHge/SFsdzNoqgPjdopJ92
o+kfF5FsnZenrfVjlOJNx9mldjI1F2GSZqURR/nVmSqZiN08f7N5poZyUL4ZWZy3
TcxlS2sUd6aRyiO3ogijR4Vj17PHOQaZKESnDKFOnq+TyjnSqJwcae5NgQI7QBFt
LfUEpyosCBxYtc5IcEHXW8oR3M4G8INFSu5KVbmb6Zhwy5FOXNFMig7EeMyJGLip
gZLE7+sKU9bQDStWLEnyh8yIiwJ4sVcwlTGN2hLZN1nH97/cW1Z77pKXe+VMMGE8
hSYUGtKW+FOgZGMB2BwfjzyvLhNkLFzXCI378fvssEkSWBTBc9B5bN22InGKEvtr
Kx4i43yaizznVnhZFBSyxdEMK5V+BLf6XrbIh+qlnhd/pduvUh67xkJ3m1PByExY
Ii5Rzt5cKgAvicDHVxJVUYV3JXrgTmCWdY1G0Z+q0vUeY9QVfsngBS5gnAsqRXfn
Em4A8ml4JAI2dMTm1JV3QAC7sZ4tRjEvZO8b69qF2vNilloquhJdDMlsuIKg8oP8
I4ZPMdGZ6Lw9odz7Cw4ecwgnklizuU0q92ralANpW1gob57uYKlasAkwc1KS8eCO
Nl99/3G/QKbTsy3Ch07IovsBt2d6tD03bkxBXcN7JoIxwQ2UMg2OXROUt5y95hvf
H++hbryALxmhBv0VQwCFrMUlh3wWY1vsONxI+wTTahWZ7CgPWegIMLt3zA5Aey4v
L/jH7SDBv3wM807AP9yy5xerlLzQSQ19co200+wBSwNJC+Bun9WSPgJpRQdeR3rl
cglrN9W7pQWVQwPjnFrnqm2UXdbXXcW3f4tF540n/iKFVSukQKQCFHTj5E1uIIAf
rv1mn/Eky3igPAOjL38NfjLy8Y1v3z+EPJbkgPc2BB7wTuCZuDqTniw5AHz0oJpY
oQVgcLgE5nEKaqwCpRULo3qmCCyddhOv7WSi1zkmB1Qz89Rb1XRA8s2Q4+tpSi7Q
EF+YU3XtN9V/Rd4FcnUhTW+1v3yiq/6+PthDB1Rh9c5c5MEwPEW2WztLNgqLV/2R
1FZ869kSqFzLxyaP1E39leLNlGes1Vn2CiwuL03RSuvjh6K9jKPXp3pdkxj1b9ly
HwjGDB3DexOfHLQfAwmIzLWgnU6vGm9QfwnQaw3XOyC9+o4C5bECdP1oCCwASrXX
nFkOdVIeRL2f6PDQatjyYlJeIxjQPTeB7l6pbSjVWz31WXBm3EnSCPYiwEx/Osyy
XDCF4g23ev6Wefaay1LgkXAdEOPPz6b2cLU8mCmjshnA7ajzx5PK8KVvq7J5MLpp
i6E0FLSWt0LgAD5NQ1Omsb7MYA0U203VsjrPc8xnTWMHZ8p4CIm5rmp72R/5omG8
J+tQYobbpl7TlINupRCQPnQt+8UEkFPP6DXXF0TsREssSOq4q1m/1BNE/3F16wgM
l3dH0xzvE4K5dzMsO6uu3mzzvBK3SnQXihJKIhbWi3R6BY45SZxQDan/De98ezlF
RftgqKi9jB5CMh6wwjLwpvlbxfiWSIuDbM6ieIIzfkpQ7V0GOElhs3ZgYiK4rnZv
ZBu9uHJxtqSiXOCh0ixtXKe0SgrPcqAXsYGAQweC5lJfXBMRa3XANZ48RFeX/YKA
i0Rx/F3BKMzJalKJiZKxemG1GYk6mtgZkH3eYK69UYCb12Z6OvWyj1FKsmH9hjpO
87iE0RZNE1eFemmugwG9mbuNq+7PJSqLLtLs99kWMeMjoVIb/AV0J3jwj3X+sMHm
09NLsOgMPNe0I6utEEaNRWco/NdeWBCpPiCAx0CKdw2maV0XbTpDIcPjFifcKd1u
TRrpTB1YtnUOPxFaPgh4ivCEZLjXcKi8HtB+LXlFvPhgnyMFUH6F7A2uSEl0FWMx
u6zs+IKdOvb8MF9BQhxaJ1Tg4sx3sfTpZYJche1KomklXMEDZvSMHvTgBqZr4lqp
k40Eq/StCVnVjipPXRqK5pXd/tvmU7vtcyHCG2iOk5gHabepkW5Hl5yzEGV2/B3k
on3gKrBhQoW13wRFElyDHF/TNsenHm4tqRQvJkpIjEN5ZFTXaX1jUAy/cPT6FzEf
fcWYd30Jz8feCENp6QpgoJxm16kj8HC6GVDEnTaz1LjeoFdZ5GDKq45qPP5J4IaG
GZKtYz80dUUK9S41UbQKa9e/Db6KfhARD44pwbcwcIMq2eYmCJAG60k4RMhmQivN
2sI6xLhddoLHWwr/fzMv6vayRrrh7gdn38bZQuOsfBum5uh3c3BX9oFY5aZz2DoB
S5ihQ9NSR+Z/VDFF+3iDGU3APFxgetP8s66vslw/k2q5Bge2hW4vSSau9xXw0e3a
/U6oDhyr0NTABtnhoCvVdcIIsY5H+arLoTr3kKHYN7nrR1UHxEDunmpRAyMj/I0E
3UekUsaSuQhVfyYE5TPxMrogJYi0YbtrbO5oGptuEmALmOjyEOzK6G4D42BZ/dSi
nBnogjHTRWKWPBCnLhV8OFsQa2JRwoyl0g78UKj+eepGJ77+1RqSZoIA2Gl41sST
+yky9MLe8/oOupk6accqSidtwDNRvvixWdmemi6HBGsMV6D0b23g+bOPecgG3ND2
Rc4KcOo2bAizfsrxz/k3b2i1ImeUzDw2DYLtTX6RJ5Hg7MpZz98HBsWCJrF4YRfv
tSxzEvoawBhrSxVuetltLikNHA8RJDcTDBCOmZGfCKHqmciE7MPz5ryGzyMAuhIr
puVZjne5VRS8w4apcwt5nFCtnufyVoKXVrVhXM79y9qI9vnpGVgAekO54twhPRS7
waH/uZko16CBdvSQ3EcwsEeidE+LBJk2IasH2lxzPwpDs5rhcKPD44YPqyivDVxX
uwGwQ9uDtKXgdJj1BcB1tUDK0iBMRcAkzk3scpkNwAsHpOfjhMZgDqdHqGFr1KVW
+hb8RWoGrZDhMZ6lmBQEWDFA/Dcf6K/bi/Su6bidn1UrD3LI8b3F1k4eTbxMrfVx
MSGBmVp10eXcKuA5+n5Qi2aV/xWwIoOF39S9p5ZkvbjU3JK07pr3n50IJPt2LQRQ
Irub/f1wR/U/+YdPhcT8tWezL+LuMgv403sDbqg61sseDLGm256Q/BBUabnY/MNK
vfhIDu8pbzGe6QigUMxBv3aozzZqqAQ9AG3bL7ggsu1lagn6EebJh6Rl1Qe/jRfJ
KFmsWfkSM5R0BjyYKuNOImHIcD/fUnUjZk3d8y4da2MSgeks5XiN62R0nUcWBRLg
67JCYVzLuxcSuxTA3P2wTacFRHqKdusNjQCpSUE8cP/87SZsRjCC8y6PrOOA7gPM
4Q0qu51AX3H34NgVdu2FNWyZvQv9O4Am+0Nrtpfb9vgDhjKQ+pr69uKeP0QzbJz9
bcW7kNAldDuTTA7b3ykl3PgE6iwtWECcGLU6wMZwT9dxRAv6ytmuVt5jfJXuEKzz
vITX0QtK0EaYSUE0w5fHRrlsL3TJLm4blON4dvoTjeVHlU3F2uyxNur81ZQtGZDd
8Z3MiZNoZDOkvFWqA/5f/8QtiSr9F9fLudGcjKmdK6w/wFOelSj4QLXHb9wv2w6S
Dx/lON5FDPxJSynpciAsgsdY37ZGwJnnagIsWa9Us5HUsiBE53WJbMHRM+aotPSS
XotecruNl5LBzhexlqra5SQ0KwaWEuloO7njg5wqg/vQ+wxpLoNhstjyaFHy5GmQ
zJBjqMABjqmZN6mTJou2K4vQDyRcw4f3fi0kQCuJGR0DfImNu+4W76jSK3RvqgXI
kGJNn6Tymt+LI/CYnh7WEdm/s/aHHdZTn71WYmZv1Q7XgbipYXvsBss81rL1IsLG
MDKC2Lv9BYi9PabzKC3bmwZgHsiQ2DnZ8xcztPi+fQYFKmY+1cNiN1Alt1qZPy6m
9uWWyIjxMc8ndF7N+eAdiTupNjuit5kkbldzoVfR8cjO+kcaCobtJCxDcuRj9Abt
q3hKT/ATsAF8q6VcqCryV34i12+jHXHs7L1nrE+SOhFTdoLxYuTjtnW5MDCeLt28
JWlDtK88stL60xWyoUNQLoang6mTYr+kQf6yr2SGBsswLUKvu+23CtfQlmJHpOZg
sKVFRYdtTISv37BwfaYNBIrqxwWzzMyfCjghqihGbf2iYfIv0oBhd6PUS83FzXio
YE1iGqipWFe7Sm3qkRBGOVqCvJylwlmywHi5xHk38nU2apzY87gI/mfDrnECDDWV
VPGLUeZ4JWnVTNDKJXrnYUvGCHVwKapaAY5r4Z0jWkbHUomD20rBotGezOmwtZl5
jG4GuXIWH4cKInbjh9mTIpKPPLi3W9kEH+r61vlhq3kwUOQ36UhCl80ytK7DYeLB
R5tUw06RikzV+9hmqxvZ0HZ3nVUuiuF7ONtlUQODskzWixMcaT+ZrpMPFig7mmZv
mvuUuiQBtJAfip8Rzqqymw5xYPhnqxZExxrOvIZCVBpW+ZTgdyNGFO4jhnnVcSWo
du98L0hLaxZdZ93tukno3Hr6XuPDMr76vPGUNLbMPJMOvm46kExcuE2o3cog/Q/i
oJvFe80N+WLyNV0BQpi0O/Wm5J8PXHK0C8BKP6+7uX1tMLLK4SAHm/6cI4eTGRkR
tMhlFyzx5IO1U/hmR2EfBnrAo2Ua/TZpMo1M4gAdj7mC6f9iSh4+wmVrl/XP5Y5O
ocM7nNfQRTuk/humLw1LJv07i4BtzIKZ1IpeoOLpAi9FRqgRLBwjQUu/pB5Y3qFD
AfhicWKKy3p7iEudDBCBTEm99TrzG5RF7CM9FzEX8G8iJ3HA4Th0eLhCiYRGxczG
p9TJ/+3k1IAVUvTXGZC3qBKW57o5QRi5g00CqUkRKWsg7QKP8i+3mVjRsov9d+6v
HQX5Ddq0SivcNsnAmOdt9NP7qHk+uURiKMyaf9GYKFuAuFH2UdYoUn/RZ87Gh6pI
BnEICC7YOsTdhl54q5c1/omoSNrb+BkGn8SG0IB+FHI8oZYYmUgI7vUWSYMAYDEh
tK5NgETP8Ro9VlPTzHpRABm4L4y2Q9YxH5/SQAdZQoFhjnPlMDRafojU7TD+wvhk
y4HVO3Ua8k2stJcsv7u5Dmu1bpNoyovYjihd/Zk6sXKjeyRAmx9YCIxodQcgVfJH
Hv8KRjOzyqHSXSLWzYUcR/5WxJtOiV+/PZ3xGmWNWGIxUncdKv3ASFsA1j821CYt
QjeakE5PQkT0Y+pp6SHg3ZTajtSdVWo2vkdMNrlteKnB8A1KFT5iwtgoWfxKK/Oq
YlUpP8iD7gbI3z9PAKmOZvkXLdSt3Li5RQ1OCQWK2p/PiSEyE2fFLz2vVtShyv3M
zRsXMuwG7wyeCOC3PT30tlBKkXIgPIueEReR3iad6nxkJgtlfoHEGrwDcDv0Z3wc
Azli/r2e9zpHn3Lb5jdgWLADfkI3FrI/KZ93uiVCLeUIWb9ilSll8nXE9o8oLVTP
IkhJl4NOlaS5wPfi9L3/t/YhU/zv4biykXNxc+K7jUbKH3dzEBh970RfPB4bPq1H
DzWu85Tor5vZVJ/j+N9r1llep84XLyYGQ69xHggLYudBI1yQ0ibks8/hzteEXnD5
TKF1h480IRuzC3UesDNDci3/lBlT3YA9lDUnaFr73sDdSkAIkNhvGVmzlFolg9Pb
f9P9UNnMrm9aDswOHturjzyJoh/IUKnkKvk/vmxwzzEMrJ3pQxCPRQWKruC/uYTQ
xAilEG4b1aIFv9fhv5NiWujTrvQQ16hm6OgIOsZBUcnab7Y+7N/3+gXFyRp5hpqn
HMOMJaHZcsHgVfLXf4/XgaFnHzkkyl2uO8IYgEHH4jNjhsRm0XGWnfur3KzeOBWy
sU//uu1xF9ySs8xRTlrmwfE5RB+G5VOq3hZjO76V/7J7MgpVjq9gReylxS2tbbIU
gktNxItjQfubJ4kBUNpVxZxzEELMpxMadA2fMjCuMO1yc/Ju/FuocT/n/7rE3NSO
9HNdwpJc88Xj4TJvMZdfg9VWOR+t69zcBJEM1na2qDizP9AKeYz28g0w77kMcReS
19qcGp5Ye+R4r2GIeW+BelxdxuShih3roDaciJcB9jdmHxBn0dgjvKfM7bQOzx4p
xuKrwtBkNSHigtfqHuuuyfe0q55oj8MGCe4nDBqsAK/Khf5yj8BgH2Rg9kARP5N7
x4HJANZX5pULjwFl8iLMGbSRGUy9wpz681LAv70IXhil6L0NwXVEDO3qS352tgKS
PVBUBWaLF6/TWYqmQOpknAa3/0rz+v5Gtn7Ymv3YcwLnMGx1vxpLGs1vpAXVop5N
rhiGqiH+0dLWK9QEgz1D1BzvjL16VHHczV3ANEzdmNydKAaExomeGIqwzg/IJYSO
kZl5iTyoZLDbRv9r+TvSXYL2MZsR7yqKhnB83Gll62AjXOarU3R38PwyAmjRPKv+
50MUd5EhQHV6j/U6YrmdKpDRc5p7THsU55Yv5lCuC+WUxmk83n7UobAE3lAZy+Vl
IkidSSReziQ+Hn5fVpC+fQArY2rMmFFBJza1UZRgj3NR5CFjqzgMOiGXN7euaAbm
tX/fdeoWGF6WE37fDNNqeXdVDu8fhJlcdD0Wsg2S42ohUQnFd9scrMDpJgKh5Kuo
xPJpnjTE9+c8uYBZi6iufcUTACf+/jWkkjkhVGNwNuhFO/F8ACJPYBnhCT6YiER6
Z4o10ohoXdcqla3H0JjdHRrnGmTPsWlcqjn4mX9Bz6D8NvYgXRlSWZDGX39Hodqm
aiUlSxJs1TKtdD3MFDbNiAwUkCLv/u+DqNb4LSRqIplhEc+1J2DNMJmdSB4JTpFS
SEXfPOtGaCG4PUrlHZMTlz+K0rbbRSsoez3sokir0L7unaeyInuLvx0WL8bLfbo8
HdvFsiyTh0DmI+QATFLiThYWY4NW3i2k1mGh9MB2qA+06kwN90lwWZnUbbnTL1Kq
qMBScVdP279bMxlSpzfeN7PuAe5470ZII2U38O9RxZ3OJQsasQbGJPkDrULNPSwo
AHLWw1vG9N1OnO9RzQbUrHBtDrp4Uc1exlL0q8n6VARHuGzPFUTSap9rR2YDuyMJ
LtUrKMwQIIScxVyfvLrO0vL6+0/bUpTs5MKYmZyZg/D9klSkYFNJIxLYGACRrS6J
lJK3oQeAMq7J4QlYKcJZgm0pqUCl9pa5b04DNqp1Fm2G3DQvoSdw/FWG+/PtNJAV
toQirEKljs673ZeDebO4igFRJGQH0JTBjHqYnPgkkl0I4eN43XUsFIH1pfrSFnJi
rRfwwpsGFdtPj2fGxMmj0yEEWBllxF3xRjjWDFZzvHvLKUgd4wY9KppMIK+lV3zJ
GaK0si4RfaWg6bTSdWLsRt79j1CZVcKX+5hwrcRIQDYtqUhU54cFqm2ZNKiyaFBt
bWvJe3PmkeROzJzmybQLvj0Qb8NPqbntSh4rj7/XX7xq8Y30X9BPXGKrjwSO5JNw
p45YRBdUjx6dqL6VIKUMkhb1Z/o2MV/ODpEcsoNxLAs2tICaFg1LJ3PtzFvMg4nF
fey+vc1ZllvKYG6lnBnKuo9ci6R3rmjz2r3fwytxV+ea1LFuBrSwwdUiFxVI6QNo
HBwYtwatkn+WoUfpF30CkmJO4Qirh7u0xP/1oW5ZkwkC0tAhCVUBC8SUkMVzgYWs
p+q+UtaNBCF2bZ2GHlq+6RsvA6fk2jLA88K9I1k74mMlfLqiqhI7WeNh1RBmWIiA
ORUMdydboiL0f8anzAkJ1hu6IL74c8exIKvHDXO88aXlyGWdjlwUqZHFG7wX+PGF
Fzdnyu7Z8krEXiUs1jC0/sBmddyxExXpZctNTLhBoy3A7uW8klxDZ45o3+x21OY4
OcbcokobZtUzJXGOqHP37zG+67vS21oCOZtnAb+F0TmZV3ANoooFXHyqX/R5bwZY
cR4zEINUuLCfq559nnTfSGnLqgosXvhKAitWIrgkfYELqcvlcqHhVYVhJgT4pgaJ
z8VyJPxnmR8WsEiAiGkPr9QCm6TOtuVjRoaWrmeYhpVMV90KrbixwZGNNu4ix2ne
6af4W8oiTJGCBPLxwH2rRk87oESh3+6qKvGYieqFAceLWTYvWvIqQvWQhWaelSKO
lMQj9E71JwMlzvDBlQ7cogRlR5DGNXc0vYrG+GRv3oEYvoEvKnS+FJcVQkAeuIz4
gulHwn4RB2nhr8llbfJAC3/UBD97stds50EfOHv08YbhfM17XERIR/OgAmkLiazm
fL7ZgfkPZd6MxlZ4Ecvw2Sh2vwRStmDUuSc7infsnKz+TfD6las4vpACaXUbGdsC
T7qP4GxFnyxN1P42Vb4Y1rm3Wf5O9nZYMPFpccKBLuDeVReP5t4h2b/tBLoRtn1u
5ra8ea7py0sf/pDIgexnW0rbDYy+00Jan6vNs7mvUA4YODgWIMyc+TLsBs+4rniQ
8EtEuyVXPnv0KVi8U9HRh0UJ59M+mMc1nxET6z8GfyvHl4I+G2FDDpb+IjsMIdWa
UwvSirrAHHyPryNAbU4XwYPyvrS15Co1ZYiUbp1NMIQ97GO2rrKZdVTuzE5+4sKi
P/otNU805qJgP5S+mPB53hAietFzjKCzcP8LHccRCmg64hPYvwJDUSz7ragRauDd
NmX/ENNiK0y2ZwV9dPHuM6AYRbrmP0FjCHHD4yTTfXJ+Cr1ttVPAs19Tut8w2ft8
Av6FAoDGxbOiVS6MaRt7spRtOt428Ykt8MRd/d3lk1dCmmLdlK0XSzpG9MAka6ma
9yUouCftM/ZX+Rxi34xnnrRdpbhN2flQoyDKl9CQPqUOV3K/Xfl5cNQ7lia2BWTp
8xkfj8e446KBneuolA/bHPOQ4qTIN9P1PlWZbvc0jiLVbjo42BRrmMx6sCnPEQM7
YVvcCtVm07P8kn3S2aLsfvQ2KawnN9cbYpzEX6XnQHWq0tD1xt9Jaw+w3mmjAewy
b7oPnmRbo4lBufiVdZk0NefRZSjcyHvGbDYcNRbg/F7oCroRaE0WYQYJ2WdW5g+h
Yf+Ug6mCveXQo6lG1kZjXMnPleCxoUTiQLjM5w2KSZxsBEd/AoF/jB83YTFA1SY5
nAo8z3IS10T5GdcWze1x5/TKfhq0TcVv3amWEj6EkrKTVHaMq+K5ISWBYIAqh7m/
j8NgMONAcwvgzHbzEoi1SafqWHu1YsbrWVEmrAnCljRGbnMP2Y+Mnsf5+ibjHG6L
s/7PYFl0kiUXghuuM+34TVK8s1uup1RhyerZpTB9mXw0HyZ+Zl/ELlbQVptpLqa1
En9ZYI08M7POiHvzdjRpzRxy/DbX3hy2dQuZHeaJM/bCYHWfEOtedKLvy+eup6dg
If4xAKPd3kpXTxTBfZ9OJTFs1SxO/t+x0Tq10Mn+kEcBhcG3T3nNfYuRry4BsYiE
ayhp8U2k+r1eBek+3MM02tQTdIi/d7KAt8TAOgEd5krPd5+KUyIxshrLsNXENpMT
TDffj9GTmKPTkRygLX7wJNuHyFKqEuoOYyrKGdKMMyl8evO/Zm521o1EOYPoGiZY
lOTAXWb5q0l46LAGgpa1O/QwveB0+3H7yqTMGPZv0kaoZuD/7ebBUXWZktCjuedp
MLTEAHuFwC7jjd+gSXJ9Zv+dSF3P21eiPlJzm2rrsS61jJexwqd1Pvbb7jkfT+UV
hGq9tW5/zFoUO/2Av5DUz5pezazDWwbtPA7aboqV4de+2ObOJRiefVnOTwBDQp1r
iX2hBD46RnNjK0w7hJi9iGNm8dX0G/E0mQavVJDlkiFIZQC2aGQV8CTYns86T9oF
+VioSjS16AxbAYQmZ4D4cSzbdnFAFOMXY9J8SP6dxXzbX/O+nXFXM8JOQ2guFeko
4ILRBmJ/AJloFxVPeKW4NusFnXo3Y/Y8xlIkKYEiABOS1CafkJZmTZ4OE1vRlGn5
W+JvBC49l+BgY9L1pgamo8Tg6rFnm/GkzLtve66DhWrpKIAyGWNCxs7T2RGyE2/1
WMduX+7HovX80cT4xrZZqkSV6d4T5OUqMpMO350JhXlzuRmUtUjUK6Xb5lzXGNv1
IZrTqMeSurKpB0rUcvlpy2OfjgqYKASLal7H5oIC9tmuGxCkNURB2c58aiz9RYtl
36HPIz+heiRrVaxaHl6OEqAoQWTnjoon3WLUEaUCG+gtwW/lsr2HbrAJ6g4AJCoH
EaaWTu4Ir0Wl78YnCppMVrmPnnL8Ezt9QiPwNje77x5NCWKrunH3iQD018nAmf2k
XOq2euxq92xcCpoYVAEINlx8HGtCb2cOKke0aJ9jUs3I4RtrDbPjB1jeTnZpOZcG
WRPEQdUkLzIb99p5a+nFiOeGRYoulYbLk6qaNk7X2SGDlBVKrTpfM6jfB4GI9HSG
Zy716MM3Snvqcglc6PiXqm5/JGhDkDp5Z8ShgJqncom4+tdrUBacJnN/rMKk7BtE
owOEtkzEEBEpOds46YTurgh8TAyRqNNC+ygy/aBv8KT0XZOnCzfOnLfI2+a/4Jqu
MVd9uez+r6W+tbC1tHGZm/WsEzPP2VkOtLK9ex4s2NBPRcWSuENayOvUtCBiETME
JWaZNhWpvXVsFO/FgB6Ndm4kit4lm1TrrR3zxYibL5OpNAD3p/EsjlUbTiJBuvgS
ask0EDnlPxeuNazvIAY5rSPfYerSEG07/s0o6/WCAzS8eG9G5qvSEq6ZCu2CU8qi
3vr/jLoUDz8GRUTb58KDnb7OH+85CwH2cuFYojfK5amIiCyFB9Sh28z2LYQtcoeT
Hoi3Jmfvo8UXGCgNm6bZGW/gx6NtBe5k2XDV9LgwDZ6pXAoUtxQQkQyFxn8ctMJh
xJL08AWw8UM5oVSvB3Q/0IUWhOWMcXZQyvWrXak5AdD8Nl2y2Fapuag+Vxxt5yCA
+OrYFniuY+cnwe/P66+jpEuf45PfMQMZZZyMCzciv9ifnC3AgFLd+CVlGhplFOkQ
onKKQjdeSiWG/iJRTE8ytdzqCVWuOya2GCYN2KNI6EIrHy9JGV3LrHQiEq+zzqL5
RmDvLlvnn6XeMxPZZlgOEAScp96yKDUkDpTTOL86E1wMwxSfSeR4i3fRd8Qsdj3A
2RaAJdPCpy2/P4e0+QKu71eYeTu0e4i7O9F49L5OXjcydg6Lg/o4sB6ySkTPcTjU
vHTPV3SH/p0xM673iNEGBPTcG+H4/aSRLsHuGb06lTVvurKqRSIFl1GgAc0aCIHM
krhgELT5t6lyfaOtjABG1mY9daexK6KDYkH4C3HFPZs+EC8MxbAw6zTM0adxtr6c
OApdtlZNWfZSTLA5ZxpQztH870GhV7f4ch0x+Ek2xBfnBzLrvhBl3AbZcdSsKByb
cX7y4oBPueeni9C693BEKxZoVLtytWRgUkS5Vbj7pUk1V3dnXTMxQ0MkQIk50vZq
gpsAKiMwhF6+KgfXaGvuEKLYvkhpf21KHN8zDt8ULVi5Dy9uHneLalLwNZmLodpv
Y0rjySbYh+vdTxBgPRuCEtBoTiBsD/SQpRpY3G+5ryYrCXjBJsSNwNjM5GTypXu3
WZVql+AFJq12Qn2Yzd5Iip2/v6ep548q6x9aPi2whOjvy9zZnCMbJx2pOG3y5wL+
7fC2E8osmBTlf1+9Uf4/MGy6jMhLwvVZRWzR20XpcBrNAs5e2oqujtnBR81TIgR7
zM4i3HgqlOg/koH7LzcHb/1dZn+0BzFaxQLBOO4oTW2yFmrJKdJWXKB+m4ily2h4
JGVgnTKrP7/2WMhM1y6FwL8tYz0Jksb9T0lrnUZTixmVxQWUZVd8UFcwjHHWDbWD
8cpclvFhnjhFSXbHsOdGzkLJ5uo7VZ6nelmaqWDn+vCDe5avxSN0ndwfczG3CbW4
uLdbgSdW0fK+D6MaFDa7wKhRwEKnZx2TYWHsb+TqluBxRLqt3IM9v4LbRTDSx6Hj
epTvljALBEowK3LDZG/Z9BpL6hjJpStC0+iLJulvAJfvHDhjdQW4NwdtgQNc+JrI
OxTysdjsiRalUqTX71nXKyssxkix+EP9a3q7zx9Q6xsK2bLSL5woq001VEFL/HiD
Pnd43g6IaIu5xfDqYTTrkWYZ+X5XkHFsYCDHdsyODV7MzXyIBnuseTNC6OP3OFqM
R51pqomzpQ505tpEdKDJwtYpkjaz/21Kz1M/dJWnaQ43d3BdJ6VvRyDyEwDeIQlU
CCPVY7uuTs2I+mtn+RvWGE3LmoG1k454qpCYf2Q7UoKdnKqZONAoJVN7qAUfg54n
ZMZvOm8iAF5pbsCI7XpC+VGOASv0irjzAtPOeCMBZ3x1X5yd+SmSreme0ZyvD5kc
fShoFkDTxMX192F8iJnAHADeh/vKXNUUuIcmK/0TDfgtNHQsVFGFZJ5XisQs+jph
yZuYM89yM6xi/FIz4Vn7YVMIMN3WNMUqoBL8ZGHaKJ1qmP5KbPPycouK2NSJbetV
XDzKNd9mY8etKAdVxfyotLFhiF2+qogjwbCixtJPBszPXB9DXUFnufL5cgCRK5dv
Hv7kbtogcsAF3nCsGMCAlPGdRPmgpBtrmqYAcpefBdJlzH3Hmqy009/MCei2fT1D
r23XPAP7Gi8x1k7hK3whUdunwX3cUchGq8o6xMs9BIb4iPRNWv4puXyPPROGCXuN
uSp8KzqEmixJkxvkSa3WTss3zOBchj27yZRKp1rryQC9DbZlScmIoXD+8nwioZtz
mN0FyEXViWgdAysLpt3Ozr2xb7cvUHozZ1KQ/j5O0wZZQC7TH40uKjK5IRu86s0z
njw/KE06iQV0At670ZwMmhPE1su6CN9icYJQtC8bLY3HVmwKvJrHn8bz14Q3N5/z
eZa2hcxAAg3it1iC0QRdSxL75ivlbfPc/3jUcjuKkI3oluV/JEOoUgPN28ObWlVT
pblK4qCNZH0x5VzPvmIr8Cp6Opw88RSwGcWOGwo+bjzszvexAtWWlBmJ+FfRcD0h
zkTDUvQk0ov0CxjKK39ASIURPbF3jJYdEheBN2ln7g3vA7aQMVWeXpRinDVdN7vZ
s4r1cz4aly3jloAxUJ5b379T2LHIjgAO4XOYdRa4dfdBZu/1gvNUnNC37rYh3Tza
z8Jvxb0G0oc8u6bH4h4QvYkZkGnCNqSZpZKUvwDgxvbzfKwIE33KR5T72sqLDgVs
DmnR58zuAD7LpNOuheBK9y6XulYJZV8ekRknCEObBdaezlAgTwfNrDnTiH3/JQC6
zji8e+NuQSBHOBBwWz5gRvDOpXG1JmFXoGFDrSntayve7KbBksBgbITOn6Ks2GtT
AEffXdZS0S4wH3pr/ZEJF807xAl+u08kexXy0oZddkkIOoTd3Qb+iT3Cc2kpiDSO
OIG0UEa+B8dBt2Bemd5RtKgPFp83lABfF4hO4Iqu36j55SniK+A6dbxoapARABUI
2N2icclDdSEOqncffAYV/drkHq8t/S9eIibLyjsUmW0sqUzti4Nw09hU82JS7K7M
MnwNNYBlhPc04f4Mee80zDYMO2H8CXYYy9DdmYoIC5Ecgxpg6XfJghAEukRYOfYN
vFszEh7EyDEZ/ZRM2rZwNLBlz0xgyZOpKXrcJpuBhC1toJIUtDDszNOrK3DcNPa5
y8OQdTyh0diKFiiCcj3EJRcfjOQQRntzEBzWXLuBXxRnruqKeDnQ8xJnUt9cD9k5
uih7u+pAPTqEKEWadnRtjehRU0uYRGxaER2kcmnIw7snEG+Wx3Ndm4e10r4HCYwK
62GfPdLhuTqXj6mnzEnBiO/QjgezqR9W2R3JP77nHYTUpz4Hq4wk3ZDAbNINJg8R
38TNcV83Ex5DTAn5jJtitamF04NsWFblrFHTE2xuEst4xb90R57ImJoh/m+FshYy
2tw0TSTvBZ6mf8e8e8yfMwGTUUIEQmLl8ICRmI+pvpY/MxzuOIVTg+qL/jZXMwQJ
VQ9oucsPAXGAmgkkziKRTNqTWOgmEe8YgJZFsNS2EIWzIFxgAooesFjLJV7kWWRc
kDgSrPdwkFPFueolqMSNRRjgdPo3FqKhQClO/2CL5OFyafStLpHSlSrNgQP8wYuq
45cJSFZONoIMW0K5tu+ZSaSbu0X6KMG4e3zjrT7pTFx6+OY9yJU9Y1PpenkAindf
xIxrKpct3pMJEqeFHH5wKCxLOI8PAh55PkE1jK6X5t3Pt5y0mSOjRAGwlV0XgZo2
4wE8kfIcCAmMykKOSMvi+fWCSSM/I49XPQjEazYvA4bk98TxhQE40m7PPJlrrqOk
VjZf67ivHGcLjOrA8DUWEoF9lRQ7vKA0TD4Rih1Uwj/XnN0Thuq4NNbTy6V8Tr7v
XP+Y6gObjIqNOoDzR3uvzf/TbhQPzwg0KDuGayrCTTJZloQ8+gr5YI6xZnLrc4I8
FKHzxPwlD66cjtXfw59Z/pJaxJeTqel4+Xw7XRdkI6CliiLlHEps+oWt+073o4jX
qCZqEgl+Em2WS6tTYNeejVAM42+EYnmgLvxte973VF5+Vt5L4JzieHBeD8W2v5TY
B31fEuJFvzCQtAb3JSOjAEUqWch2fxDrZkJh35cUrCn1bHgOPMrQM1oVF4IzcI/2
Qc11qYvdbLfhdeeXgX0jL57UyVKd6idGnWY51lxEn+vNMufj6S03ezyG4Z+O7twV
zzg0fq8dWOxgNKE22t/UjNRE1/awFMBLY+LwMv9Yc5XTMjaWFSmg5E17oZr5om/4
JuMeun73vAJeUhEmQP1012pAENrMX143FPK0q3ptiyyH0Z0QSbVB6hjYkTT8uXxR
qSk5PEk7EXWZ3DOoWzCufcBJ+TEaZTo5hdRU76pU0OcG6ypIYYklKGcc8nyXJbZl
/WsqdxanDLwOhWzeeuLcZ3rrm1YqMgInYBFGzbHMXBs/H5bQZZgudC043AnM7Unj
DJ5E7ZLBuBSCBg7JixVpNcjwuWZ2Kyxlof47M7R+dtawLdkGgLi9bsoCwE0QuT6V
UQ+0M20gY1u3Y9WEg18nFy5EjtSHVhhUTF71zlWfnUMdrRQGfo2hSMex2Z5l/y8q
abZDivzW2yJhkKrJ6Map4P4LV0diG1BlDoL3dcrcjdhsS5dWubn6/CKxI3Ri2rUD
mQ1PwXM00RjEl4+ziWYUu4Zfr7KDEL/s77r4lsW86hAs5lvJQwQC7vgDXjTZqeAN
M5csW7HykQH25/cAk8Q+E+WnNUanXrkttzncPbqM5SiV1bGfyafwstpgJ4tmKzXj
URuRGJG+nVN5uVLmQXnyMfABsESq9g5wsk30hlgIRCKCSOskrBNtba3XwuoLEV4i
DoNXtWvgDqgBlQDRBfvonfSuvHjfE+2DN4H+zyEIlafF9RIkfzkopi4Y3BjeocaH
eKgTnGnT/DagvS4if1sjl/c1iC9og9PBxhRca9iYlQYfdKVT+/YBC4HNrj2EECyq
vb8QuSR9T1KEeTF2D/IupXi2C1RW0RUI/yy803KWBNFysW+NYvlcuiU/08JEtXtM
JJPg+TJvoIyOhQFhcmZFKKH7lrbYY1AqrQiKWbCEKdp/0Fv1eYTmS0wIao3eNzr2
CmbMsqmmofOqliMQ349HYeCsrYnQ2ijSJYmfzEZoT/Z7H/XGqeQdV3DVAWXjQhIY
lwVG9EyN42lMHu4egeCGOmXk/hJ1seEdPRVCrQa8l9KsGeA5U4v0pvKf4zHrWBnv
WC0sjPYeKSbZS8ovNkqzMokLxzEcL5KJY8WqGdnlqHAz5Msvp/lPih4WSQOFnDlz
hiZBb0MWnK5SZ5Ji1S8KpKObqPxza27jFAxI8JbmXCva27i5c2ibbn5FGS+/A2eE
sZNUf0riEeRH+fWgEOFcyBPRWV1YJ0X0gbyHxmAIC2zH2uvot0GfaDHy25HfL9kc
AXwXchUyzP0wiv/I1Bt5XsEEA16XOy1McDYsRH5Gi8NKPwLsHzD1ELApdDlnZjSu
OJPpA3cHG01S0jv8M4UoGflmA7OvI0+j6QqJ7Q+LtDk4Y0xOg6qbUrTd3emQC56B
rD8QX8T8ikJlObbEC027rk+cNQ24HFJV8BFTClV/pyn59AyUVoN+IxEX4QaN6FpL
XLjXHR+q0znCJvLuKgM3mdIn6gmeYGiQqTowkDQYF4HlESzJdnRS+BVoPLrG0DpF
o7lmFVmo13JJX3VHfNZkZ8uxvYtyjt++wwlI4bV5hrO6taHcGvbVUrR4JdG/Q10S
6Pne+Ue7G4TRRIozG5qkuLGSar5/FzVIsMS5qdsXJwbyI6f9vp2KtCLAWd+G92iG
dWi40pawFLFYonq9PNrNiqw6NBG9CTvXyfvGFA/57d57wDx2k4MX9Y0xhlLr1vrj
Zm0VusaTqmVo28QtERvqFIzn3BLoej93ea/QdI6N/h3wKB8LjKGzWEn/WT8+aBPQ
7HTgASPlh7v1wefNXRkB8eLhrxVZqM7URR4eClgh0CPVrZk1lh4bM07UQ7DT4jVy
qcolpy0Z83MBzBniJaST+cnOdpzQZq/Wh6KQZzWlRXZyPfakKkOA9AOZ384ZivJG
Blcx37FMOFS2MLWRewjwq7OTQtmv7OfdNIX07HwZkYVC/yiPb+pq7FLFgQVZ+Mof
tR/42RfV1K52/KVythCUjSBGZMpxZlu+p4thQBDDjlFq6UAplXC5BcXmKaqVnY9v
DbL6lUidIkYvRGiOKQXj7DRHVDqLqYdBt1pBdhbV+DJlJpGqYw9oa/0iIl2A/WGB
jbYZaL7TEVgdVD1Yuh0npeh+tgVapUxrqmF6/1AZ1bF1tvztHeHo+M2COfGwG8P4
m/9GzUMCHIIU2oUKFjH/S5gXXz0iStr++H7nSsoSolAAIN2NOKJfXrun/tn0vaKr
udOUbPcK+lB4C/PQKFtOIIqAHq5gHfkRS/4/FV/lQ7cd3LMdR8SwJVh8NoBheW57
XnW9UC5Y9Ps6dD6rPSYEWrDzJ1oX15jfJYupGLuiIcBn7hldgXeqwR1kMt5ZvyTT
3Kw5iSPY8aZOm8rCrgaKxvue3/FDweheIEZiuTO73KYI6CGKui9EYVs0xhoYpFa0
NNg3PZQki1XqyqUGUXhrBgsu9WeiTZDczwkmZrsUuAQpSNIsa2nWRgpCXSZffqu+
fmikAJx+Xxs1HeawMI94+qOB7De3mXJhSpq2hJeR3Oh7Ob1W/2/xl5jIHFkZBsZL
/07W05oNb5bkmbkpuIZSdpO2fQMtl1ydPRxSyfMGcT8g0CgvIl+7VJTrKBw/20Mw
RmsJyHh1HiOpVUPPf+26UjzI3Tr6mCSZN4fXLksMGPHbxBaP2VT+nahzjGG7Os9N
sN50V6SRU6MvMFBzynybes9q2afI/e4B/8MF5KakSQaOeD9TOAjkps0ijWk3VG6j
VwWDoeQrWqDJjUMC3tcK+ObySxTCEBzmBMDY1aReqsuQKwsm+s65ZWUXZ3gJXSjw
OgkQ5caVOO6Nx6UTD3vW3zIgqbPsaNcz/ig/Rl+F3mLdTuxd9+tn3xzsHOmX8ARW
5L322n2nZlM7a4atDlsxRMVsGtjAqZ4+ntfxGpoOMt6z+dNKs1rHt6pK5NYJvjkP
He1A29iADLxD8oNmDeYyWWiX1ji/QJ2v2HSNMbGhxvzNw6ChKw6OHPWaAHIv4UDh
aXkha6LxiT/ko6yZKoHgLijpnX4MsNTRxnDkbsSgslw93g+zPLCKyRhgcvRuJRN2
PP77kpIHwzU1VHDcng2rX8uZr8nxbWn+Hd25K4SycXDmG8D14uZXJCoLVf3AW8dk
1PYKpwLq6dWGT3JPJvhr99bvlxiG3Xi29HZa2n0nEZ6PyRsr1EMF8Gn9ESjKJvn0
p1aE/sTaQSpsyRr/sV0tUIyGDe7HuvJBUnXBv4G+Rx338hYRS1kAL8hK+Cjl6HAj
eCTdjLYrGMrwpeyjoeFAnHpYxAmOZbHhEMbRpAvkhZ02gLpvF9Ivs9Bo3iksWJEO
nBAYDb/dUP7HlX8RamydyQHLon5UTALEkBh3iLMOYSimyNMnWHB1ylOhZ3WSRKtP
Lj8JUBZI+YrpguY1ZzU6AotdtAYRQ+FKcAMgoG01oMYc3Warex5Vl+F7OQ+oqr01
9ltFE6UR0RKhNNfJUsAko5BK9gaKXYPA/e7+UwKTDN16x75U1XHJ2iF4SNfzts6K
dAlHaqFHdODW+/LE8A3VFNqBrJpghPT1zBHZ8HtBfcR9AtXN2k1xLexAE3Qd6pBX
/0fJY8qlWJuoSc2+j+eQnkIkkGlm13NzJ+KnVlFQUG5PSm2T1C2fZXlNtLUtPWni
v7Cc2hS612lkOx1JKN/a2RyxlKr9LDGcktzE1/BKKbau7y5gxdlGQh0OHtx8Y7tf
UluQ/NHWnIQxPsEAM0SxR9c6AwlZQvRYbRnbMmOhd3e23KlWJbvvQ0v53YYnmoJ0
VYyUqC86s+r7AJcBdnN5NAg8j1g6VuAqMYTCbhUeRu/+i6oO8jC2tN/wCNMzThFb
p8YTTeLFbR+Z/yqVdImihftP+XePzFTTL4RYhJz2WfO+PPMIvMLWISWhWNTyvx36
QT3UIBofkB9mhwIhc0v3zJNl1wkwwWK810MQJZZ43H4eEzMNIZ3k3/fyuf5+Ih4H
n/c7vHrTFVQnkTdNENc1wYqoijHfJDeOcfYwgRPBZ77n3MZG4WqgzMFWx5UgTaSv
5yFoomKX1YWmTxP70m2B/myx28XhFYVqvlztPbLI77r92/iwJ1zaZVAorlFe2rGs
BY0mkzqBV//XQdX9/zacNRx1mNwfPpK+KDdFs4RRhIm/0IzdxBZMf0HFW8Tqt1/Y
cPT0lfQ0W33op5gh3mzVxPRsX/sWEWEKqJdNTIaWwV7NWoNTZKoL669FhqD8cidd
f2KluGDOnrTTqPnaayfSNFHTy/ThvDkKMWVzN+5JZRYbg+M+pgkQW6+2DtrgvT83
K52VI+V+diYQfqBC2H7SFok2m5Ugp/r1ZOCw4PHbYe/W4fQucANIERgmqhpXpR7R
NeOf7RrjZg99UytXivfBkVRIYdZr/ftasSV6GE0JMhKuKvoJe43yMU2iaeTf1Xgo
xSpLCSp4IcV5IE2Z4u0r6nOpljFbHyz33BA88LDTdRVq4S9M9AC8fbRAryeue5pf
r0W8SYKyOi4OW2Zwiavyimdmvf3AJDZoZBFu3pPwmPTywmHhiBzmUJtdPceIUL+l
27mgKQjmh63n29YDuHDN+L2V0lCT/tCaLmqWNxkXU5YiLZWK607tgXST/gvf4jQa
+pXcpJtnkuZYwFE0Dm9futxL5uBBT5TTb8Yrq6Kax++cxtF2HC2ob3hiYCqGG6wD
Opf7d3TvBlD0BvYSSq50+wBiiTzXzMT3tJVzeJb0if99l6RZFwBrI+UsM+lSF+O2
/NhRqpa4VLhaXVQkCPFhYuge9C/ATJE2YpmU3N8lb0pRrx8zp0FXI3FVsh3qPKe6
L45Xv5D6pdGWbht6EWHcM1HDemvbtAStH+Vx/wECrIhpk7c/V4dq1MVhoyqJHuDx
6zyAmOvwLvXq4fGGhesBnqMMj/r3SS66NvYQE+9Hi05MUJwrc6Lx4/a6D9VpceaV
q0TnN8t0gOyrMhdJF1sl8Uf9hdzm5Zw0n9aIRNePwcJqLI9BQmC0LWCN4NHaLHUc
plBR2WsY0kroz3gp3l9r9FyWk6WYR2a/jmY/eR0aoqFFeeO74e28jDedpk0eKNip
/m+AjbKhlDeMgYst4BH/bBgkSkEOBYNjEtcn/I/Ja/PtHG2I0Q0CyZFRoAviBqdE
34M4FP9yb8PGRDthl/V37IfH6XrY0LpVFyhjHY1d0ohJnCqe1q89kxI22tPqV+Lv
8D64igoIVIACQAjyzKOWkbwScqXlpzCljfcLDOMXJ/o9lVCO3Y3fQoDOgcb5EW79
slGwPoU3qldHEAertZPQVlFxPoBEj+quYSvVQI22iivjORb+W36v5wpr4Ieeh3U7
4ZYkGiVRZMVWr8gtyuekS+D8o6V2oxR11FA8bP3F8XTfqK6u3BMVceKnnrvEcDYn
IbS8rPoi7MHet9fJumJZnB90YmSlLEDFDVD/+chaNglPIO+9U+J/gfi7QdoYTJwh
YCp5sQpN8U+vEUgIHbOga2iju5w2wicQduS8KG4hgMk2RSQiV6MxbXH3mzbykIZf
R6FenrmRnbiKV3n240hIfkArwp04QDLtRAhJQg99a19SEjUfxa5j+noi8bIoJ9tW
SHxIqddiDH7i0mdEzPL9MX11cNsGQB/+KnTo6JNc77m3ZM7YAnIwJUaUolmt5nQ/
74Fp9FF/nYxMm0ou+RKF8gb3zOWWXOfXyqHNbzCgnkCLiuZp9R7X8AWYfZa9LeMR
PRIyS8Jqg0WlM5ItqkecOW8qW3v7QUNYX7zvG1RIHmwYbiCg4q73TvhKc6SWbqoz
cNxFcBAivCMjCLn3Tvm/q/S8AjXLwNEOwE7uMDFZqNE9D1sZxcy4hS9H7UmpuZbi
SyGRYECLuTMVQviAzbQqaPR+3VCosCofW0UJVtYqtTANVXfwL3k8o8VDTzNhoUKE
lSyQheV5rYAwVgMFRCPRTuk7dRygo2V450SILq5uAeqenwlw2j+2UgNnkFIfLRHn
lXK1ZRrXFynov8IraHAteLdeevPGR/xm0/XliXlvVrWt6sQ/dKcFlRbjARoRDrAu
GnSW74ZE0rf28l1IW8gQB+Vwf/5Yj/+Cs909fLXaHH+aerZhBhuKJrHlHO+GR5Pq
tncMAyv5eOPka2p4qZTStdH780SB947G2vQR9lNb6D6+LYyzZ+yitpdFzw0Bdpu6
STvFPzn5qpF4LtLrxHj/qFztogDYRU13GMsOMZMDQWBaOUOBTYeBZ5qYypshWuS8
oKwezWctEDkvxhMins6bc+m+65eKU2EWpgMaWuhv5rcb0+7LxiW8MkDntaNG4onI
FhnF02rTyj+0DMqMTWrl8NTUd0cL38dwBZA4vPaotLaFDTZu3vo1jyJabYXGCkck
MyOAG3tIiaAPXdaY008OoqAE4RBprqzFyEIfSW0s5BrX8ZIoFSfRwlrB0NoNug4p
PSGeTfrJPrL06Lycr4f92sVcFn7ttgTnrjI1T2Q7/CJYz4Z3RCvGMXKt3JzP9sPc
OR14Qsb3X75NzHv++Ux7Us9eZ0SD+XOtfAvWwPAvfNpqrDtMhiWl6kd8GA5VbjRN
wpWsgjnUOPG27IdF9VjHIJJW10hIMfd0n3QPNpWUt+v0dy2TEzElWEyeAaT0VMjT
GrOG+oyVYGTL1Stt2Kb+n97ijfcZABh4f6C5lNfrbEosk7Wejy9q+cqt0+raxbLC
92etPm15WM59/LBpcWsUs6Y0TT5g2jlH1dNTlFPEFR+F+sz/XJLW8gUvNOeGELx+
AvNS6Kzf86OB46Kc+UJxJQG0wsZ7ZjpKmp885qlUJoOPP1KnNHi0WNgOrPuaAza0
jBDAI1bHReLxD6yK3q5Iu41LAAym3kWFNNmPl7FMicX+rV9KPWcb8zjMwE1d+GPt
aZ1F9p4eHqkJ+gt9vLdYKhXI1FVfTTJQzogMTh7F9IIB5WU6WdLLOWY7CjU0vD88
x+CPu7azcXo+gHceVbv2KeyYjX3CuszhiBeOC0mPVgQD+3XNXvlWLgfCEyNEcCP1
e9geIUb0Iv/MsU2idY8vz4iRVaAiLKFsnbNS+ejO+Qwaq+mx8QZQH/0ZU8UEKWLB
JvXk1MVVCLq/MlVuqFx6jFws6ZlBswooChLfWPV/mbDczDECicaHzvSCJR6yvFmD
7tu6UR9aFPSOY5Hww+TFBU58iT1UPOUQM/pZNqdfYbbF91yO3/jtXSBHH+TX1TMw
NUr2t1D9JdiVMyWPb5FTLLIqAS8voBrxmPTMzIdh7vHWrDCwIqd1TXnVl82tj0fZ
EutZ4IGxXoWgxvwwXvxjx+04mtJ+ea+MG5odna0x1/kycbY2VUBnF5b1gbGlaTDl
Kl8nLLLQKi5mLuMIeFLB5Dx5q7HIqjHJoBVV9bKmW3CDqcC4sAss6awhSbuwfOBw
RD80cooqak8W0SYnvdAUfP9JWeEq3LY+XJUchfGB0U+35OpL9cBemHIqop/pIjHB
kxVeHqTxDBf1kINCrZAk/8lFWpeN6j90H9WWuUkEphEcPJpss/VAQWGNBfNW9vgS
up6LrK59mhc788keCsoE9wf/b4D1hwy2kzNljgBCxKf+8jr0+zZJBYWfJ9zqXRvS
DDBe10zqu0kJd04A3zoyAbMbRbVicpAdSVeXk7wBw7t5dhh1VodUEHzAp1BmDMRC
Un+XziHK5PFEwUsLNEAHMBdScyiPi7AKeSFRFRstkA0x/mWgHghcf7n1TewlJLsc
OJTJrDXCos4mAKB8S2KNv3rVuwuJ02tBOJrjAgfifnKhvTyn9a1GV2pG8FszRl+k
y8fcIzCQFnwgIwV1sK1bo2Mnw3obG/eHcgKjtpeO+TgGXnvOIISXWHR3iu7SFE6t
vESVCtuWXbdlClWRQwUBQt/eVNayrGDzXkw0UEQCqvAG7viSBAPoAv4PAa9pAO9c
/uFqSVAZRunDUnxwUeNmTu7oDGvVusapNc6IRX/tq2pbzZtVgzAPPRTC6YFftlj/
voSFBQNrYWLPiyT2fA7BOMtsL0wMydnbSh8ti4vcg6WUJNND0AX2P9c8e3DP6aHj
myBVXA5in7ib7R9zyuonD561PN3Bbno02iZXYTaEh5fWYXxgKLPHZLwtNiJWmqI9
omMvxCuDa+kOh89SauHaXZo22Ow5UN9ZidYaTxhj5+zI6Y/+aDL52lqETZTYK9OB
7lwBZsTh7NBQ1dIi62eYN4a0yJPJgnwOK8S8XgLB8pGGW3K8YOzAw9TgIuCF1UzP
cpo5QTQaZtsYhYIlZcQH5VrAzd3Gh2XQ7Q8wveeziphqXR59rP0avQI+U++L2bOu
tsDXZDQ32urdVD8J0wfWeBcJtzryq8H1Lln1ZfzygVNMw1/+1FF9tRSqRnPuHeDe
tdcBXN3whRcD3rfNfQE5uxLM+mFp4MuZorZFUwrvLagwTlfHqPCKwQWI29IvonsW
QDsBpHnttMvhzV+teULRTh706H2o/MIZPRqwscgRWCQTXjBHa7ChqshKWVsSvPMR
Eg3yOTkriymCpmFhlU0TjbLL+y/2L1guB7JbWMsw79i5GYiktdk0YzudlKQaKMAT
kXK1jD0TwhTwonUGN0nP8Ppon/TdgD7IOzvTYI+KkWxMnWvGoXWuPUkyhEjdHM3x
KQUVJP/waoUSexXW4Tlvlj8izPlvBUWcJWHlGWwmQkqdOMBe03z4SiBJt1HVLkVB
Tfp4qtqAZKQtfRcjeu/BQ+gz9UiTyxYOj2X1t6u+UUFnzY2vyafnpSPY/+2eIiJc
WU20dd9PBkgBlpLUFqyXIHEIzkRmxEBso9mNjxzgVjwNC6ky2IKQYwMt1tWjOXgi
OXk5djDlgDcSqs+x5ml5B1tK3j1IFi9JcSB7IUQCBit13FtYHEDPzsgNSH09Fmdb
INsMj4DKmrrCF51nDJ6VuIx01mFkbpyoFqIF6N3kGyDwiMk9KmnjwpxY0xTMBWQ9
8gLugOTyalGDlDfYZJnK9ghoJAGhm93C/P51pq1mFVo/iGVSTsnufplcPvEnhfLQ
/v9xwnm6Qh54G1OSRXZauRv7xzO771FloAhw3Sob0Y+0C4KOVk9ZcBSnkL2MDbxg
1rwJzcHoBemOzW4QpHAC6ZHfYaWubTmZMJnSG/ubdu8C0WtldK1HLyzTJle6lvHh
ni3BJI/x1qGNZaFIjb2eF2DjPZw8dDABz9e5pedAdV1nM8VLhpexd0lgRIqCUDjm
Z7hCay5RBwhxpq8/z+hD+JnJ5BbWcIKx+t4/PQuw7gkzN0pKdVAvSzNCn9peEWgI
aHHlnSmJrPktRlELMCwTEht+SNyFYJTORP9ukSHZGI9aQpmj7hO3yCZBZS7DUQyY
zoRH1aViB8QcBlr1UV3K362vtHq0VCYFNpj78V8GHbsz79iVNW9NbB+8/02odGj7
wgj01wsIZWJRZdGpIp2nMrFigMCxnZdPv6E+8E4Zo8nlzFInHzR0qsOOjgKRzZvV
XWL2iSObd4BYDPt161Telv8WA9AWJQFiD5yO0SVVW7Qc0n25qyomJFj3bEKuuQy/
kWqmQ3HEEq6wNv9spjLq0BSFlcbohfv6zmguaErP/8CnEMi1RjGPlQoWum07Qz8k
vGaWe3JYVtjUMXqp9KvoyoxI4mBVZW/9rPrSsbvgs2LtDypH9ZMwdQiMdfYJARU/
/qg/nhCIHNYv8BTB607id53jAhg8jr2Z6lAkZ2BR1+eNDFcaAw4CcHhCOAwjHbD4
NIRenYeKsIIZkkJIVujj308ebKTtPHtTRKAsqClauqexHRH1PY/Gpj4ztCEQU79k
GWdN/qLJ4YLj72SpvB8pgL5WO19WWbgDfoS1cvBhA2osUt68TTQ3wqZQHmqzhLw1
6hvXVD8b3hWtQ8IPLd2+amnbOFeVCISYj+OkO56eOhsBp1G0O9wG3wfzenlJ9Zq1
Vxb3wwCaFaxS+2bRJeMLmvkktyC5R9Zp84a3cFc32rNJ2nEsiRe5KHR9YQwAcCjE
AmjHtnVUPrHX8fPZtKeJYa91Jc6GMJUgq7cHVZLJS1rxLdeFW5x5UfRPclyuL4/7
3LJBN8Iy+1MaJPVt8f/xkjUoDra1FUWMWi6UlymzeWqrkaBH33R4XwEtEzap5tY2
1R1UA3x19mDbbYTYkq3GS8PmbaEaaQyUridw9zHfaNl3IgpkTuyuaxmp9+5IFdPr
CM1WCk2nOz2A+PGbsUpBsfV8e6LYRaGRPKwnfVrN088WmmeiYAC3YB9K9whgGkxt
Z3hIVIhXIEyCLh5xSM1P0Bw9G1CUEEfZyI2H38PzC/w8oO5KeqHPM+qagBbe4vYZ
j8xTivjxuoEc5uC0OfGE4jh/LNFue8BxAT/6h9IbCwnVxUZBqEi+ZWvaverEPeRQ
/VQKMs2Pe24M3s6v4zPAmHwM291n2sqxXo6dPE3eaNAo4sImIRGGwaFsZL7Z5huo
78PHtsZx8wMPB5+7dTU40BRl/Azb6ObCNJ0RayXBXoDFOcX837QLNHEyl5iaoLAM
z8r2XMmcQwn86HNRXu/JAixlRpuM7b6kNbF3kCuOvbhScn4NFUjh5TPH+pgLM/jg
IlyafHV92UTN0kdsclAxdElOyDIfJsAfvxM6qxYmXr3y8TTN7/Y74WoC3B0vbWll
gZdVMfXd2B6md40qie1i6TFfux4lguaHlEFk89aNassfpC0d5S/7xbMnjuf2jO3m
VQ4K4g1BjJG7fM3bq+LZRuXvevS6MhA9T3IMf6FG31ButL9a9y7nhCo8dYv8Y9cD
yWsQQOuxZ42kzusn2AgSgJIqa0W8DDfofG538FeGL5bzBHa6U+6mCSFjN/TnG5p3
bhwXItQtiYHqcUC69K1EYsmc+X1Ljf1BJ/4SAgvyQzwRAu29jxHbuh1iXNyuyqx3
uI6iXZltk8IB5d/lNOmrwuvQgH073UIScPQbXrpWruM4lU3MfVBgFnk5p3Y3B7mU
2zjOCvlf91D+VjAusGP15iRZpLxW3pmTybMI/2B+ERziWlZUaapdBtAjzGaB3YFe
Gm+4aPv/rbfhSEe3nMIT3ZIbPNbAzo4KiJHWl/OEekGkOlUOrftXQLLtd6R54bqG
LJJnuiOFdyvNrC8t7DQr22Cbqfo43zrOJ9ea/9+8IbQ/zwn+7x6Qpz5a5qv3RRKx
3lu/bJvXQvRFNx5zlT99O436/ogmc7afDQtpChZkOwdpwTxbZgUBeNfQsO7/HaeD
ciIYTRY8jwGULttnYgsl/2uCeSWYdS6wSSr/MAH+9/DKfXgxSKAPtANc+2qBppqZ
VRkoD6VjqjIjgmAwtGoQMclP0Po9zhUz+kTZ3iRcSlLsGZOS25JKF5y8x1Y0Jl7L
SjQjVQUWH6l5TDf8q8FZ9EcRE3Ah2eyPp3tP8Dt5t81+3Ag7M+T5uNFAOF9blwbM
dw6uA2oQ7ftEYTrTnGop4HOhMArGzM2DO2s0qufqgNNoS4cSfsLP/xJczS+ja02A
c0EFJFw4b3j7rO89Pi+qsHFd1W1XY+y6yPrqv4Czl1a3bQagr6tYLU1ZfafFulrC
69+qDos2tHhnY8pB0sRpkBF8s2fRRU5J2kgPK2W+EGTxN3IzXw1sJVL49kuAGWMF
Y5uzp/tdZNlSlCWAqv+sBplMHbDyfXqcmsi1ovJjkfeRZEj+/bZpXOCRwBM5GwBP
GcGspDHpMhWJ6HJUdNf7UzGqMe07DR28uCKGaWSX07PHt5QE4zpcX05r24YXVupX
JwNBQswjvu75kh7zcnFdfRk+x1KKhrKfxAKLGjWozC85FcxkYU11WgW7VfxrCECr
m5CpdZAZ+ODkYbPcZNzyAWsgoXTihKYcfeLMPnKCQ6t3IT5/hjchsbIThP2DcGj8
0DjYNxrAGFIxSyPHqMjweHPgZ7AALM3P5bcqe34QWed0kWzJqQNT4bqhoYRnh8+u
ewpLyOixU8uu6g1+KvIHLubMKqSIWl1zJLl3DCHHmAktceZRwMaudLva+kmYBaBJ
W12IM4ezr9JoHyfMpZ5S75APbaWOPdF6yu/s8i8zBD8A2WAMVGnn4hcORBqxTVkE
R8XqU9zean7NlwW/HIRwPzzyx3PDU7xviaYkpvx94Hm7SoRtM+TKHtTCAicRM5Dd
uARq/Fx7Qkj9k0vesd/BuYbsPmP75d8be8sglaHq9DXVkAthJh6ve6fpsDhdtpxx
ilRT/1nBzHX3upH3vAmliSoIotQlvK+A+KvMa3BW4bVoy9/cCj0/J+niqxZNYD1/
xh6FM446hJ6Xo3BQl96xMnD8Uc7V0OPpnBBNpI0t9kk6Geav/T4Sq4vP961i6Cg1
HXJBMxFukqAxJtK2pMtO7KbsftAi0kIStZmWmWSQqlimX6P3zCaiPNmuRQDhddql
CoOtPHR6PBpRmKsQmUXTrQIg0SmPAUWEgWRHFyGyjYCh3hHbFIB4RwEBxyY2bX2a
ZO34KmPOoy5gttNnYjIj7ZxXWQDFXleonNbxLnCZyBLhDqdc2fY7uS7Y0dr2X6cT
D4sWUw17drYwMWgvNFYwUO08fbCbcWlAfBM0iZj4iIeOLo1Qr6IReTwFMYyNYXwa
j2NLGRRKNTYrlaH/wDW2QA9nZaaURh6SHnonZZ+6KoPTrSeqCO/hhRprhDx4/tHH
e3n9JmGfaZWJPH4wbdBjk258lIKBEQiz2+eb0LSkm5iBoi/eJOL5v+sEHAUil8rz
Eri/LUVKMTxWKuo6u9R6zwKYs9S+PdLz4N2IwZOQcRtj5MrFmgIZXeNTaqrPZAeA
gpFAZQZGEo/3OxEg479XhauBpB1xtXPY9I9ZRFzMIW7tzpFbROFTffZ6t8YyOwOk
BDtfCF446T/UdRkLmtFmwOkQYgdd+22WKTZaXUuwiIZYyIzoR5e0feJzVDb8BgLD
gUNEiMvwDRJ6xp+uzEVkL3ubIvbK7V0efz7Pu1JGZGocZOKNfT5yCdVNJPadc1YI
f3JxPWfnouhHSjjU4CUGyCujo1bnseO+Zz+zNpKYDNacwr8bt1db7WLzm8lb4xkt
jCMIx/uukZcxlqqTB3N+xvWOoXHyXXHCSxtpmNuq+m+9uUTUcaDy/pZnbANlPHi0
P3n2HwYZ+9ZFEKo+FBIrR6UHF6gCoF6eEaf2DE/k5xQO7/VDISSmsuRGclM3na4P
ZQhifKc4Zg6FV6/I6rto6uo2KWTVBFeXo2KRqU9RW1PJpU9+FUmJVL80meZq4Sem
WzsHpbMrw1A2IsoAmKihslAVQTuseAPbcB+iserXI0/WgP6zDkgjFsX9ItsVfM59
Po/Srphi9yrXGP4rDzLjk0ddKyRR2A/kNcTFNaOArBLbShNZFzOv7YW81b4ZFpgY
45ePwv1VD6Et/QJ1wlM2PLFjESsjOhUHdFTgIhoWYtR0/pneh9GdDuG8uwlw0CUV
GtY1wBPqvy8JEPD8inV8L4i/cR7gLkUmh6sIrwWm9MvNmRiKHx58LJ5gChl/RqqS
5KyG0c69vUn4ok/2xipiN4h/ZRuW8QPHdxHUQae3UbCB692Mk6exjdCjnd0L4roQ
DM6WBgO6HeqNr+JY6FEHe9hbFhiXTdWEItC6cNU2iBiQ12aqpoEvSWv2CD0RDqi/
NOrKgwEhJUXUMYspNjrCAvZgMk58ExX2126+wjRSVk0vWgYZ0wQIjlhfohTVT2Wp
KbGLL1+jUqtexxUAqO3kpN0NBIsM0BhrwUtfEiay3xg7USW5+s1ggMs3RjQwdvMh
0EK3+/OZsE8TuL92D2eUrnL6U0OOITy/VnhHML4kNDGJN3SnHb5TyU3rut1n5Oo9
clOtg9efjAGeE1ztk+8LyRrIP9TnL+/GkEeFLwtuXyLPkYrE08XxwUSQCnmRJN4l
BzuBqPZys1bBNsuPO+5HglxcNEm4D2EFeUJAkqMsdG33GGP4FVjjtNr+N/LRUNCM
j8B9wbks49rim2r8Opg50pqDYfOSg+4480iqaQ3TR1p0NSl06Te5t9OSPFC0RlKW
CZc8iPeSFUIKF2pzRhWG5q+3dqA/9NGkRPnDJdEi6Ja0/FvwlVf6gHifRRSdPBno
O9MVlqEPRVI/4ckeF5+1LIbE436ahCjXkHn5TYCuQLjfDMLjzx9wEzOIOmBr6t63
sGIjLqo1fGSWJPtICR9KWYSb/lwA2YShG/Ve189+outiNFHgia9Ythy+uEKe07zU
rBW8udp8oBoDoqY5Y2pWqhveurvti51fVjwgZ7xMLk/jl2bCCv1On1XPTC6WBrNB
Akk34rE+P4V61VFkNgWm/sl6+4TJo8QaKoYE0qwsSQyfhyjV5c7agwgcencYypNg
dFeKZZ/Slv5zzRCi0fRo0bv6/EmYZA3eqHwhB6oyS0jlNsw5vNnYRl0diVHltOg5
QHueFkvQf0qFfJt6IdKI4pAZ4i0gKldZ10JMhv1igI9WSlaHi48lH1AvQe2928Q3
bzAncJUa4pDc0mS1Wg7e4LYGLfOvMnXGJ8Zme2lAfAWaSTNAZM+v24PioILjTa9u
36Q1XxxGcUVRr5EydpwsqO6v3NeBvE8cqYK8O7fGASJwoqMaBWPNmuVOjJZPR8st
KAs5Eb46K4AB0RtujrH1skkWQSRnOH8pXU8PIuRU6RGtTErZQBKCo3JadA2CcmTj
EougCPxfd2LVS5pDQtuVedhhj9JibnFGQQMAczEinQgHCgNb+4wFUF2VWQOGLLH+
mmAD9Dxv7Er8yfy0rWrwMM1iesKeuuFJbOaAQLpJZcpYrbSHO1HYPMHnaBNFL7k+
lUm0HOU+zuLSKyfDeN/5SRzYX9L0Zoe92WHwnPWcmRcLlAjTgUnKSsQX5l4ZDRBq
jYKx+rswXjIbCmNFrrB4466k7rQXZGBem20UYsbIiA8EDjjAYpUXaveDSLMDbdMr
4LjFNibG+S5+Sa7wrY0vuHwrQ+MY++dgd5whfXK1s5fQ3qBuL3IScoeeugpeADEr
KDPCb79UHIEw6qZMKE1wv9n7dq/HCaS+u5us6/PMlM8l6W6brbJPsSpnlihOUsXW
GvZSq+8XULGQBR3z7f/CZw5W8fvVCI8ZcrWwAjI0lgobJ8f9XnSG0qovEbf9IZRl
JP6mZvzST0GeD7LG+ddBJReDMdGNENPfuibBF8EhFNFKe4YQJWnQSgALYExUjGL6
NUKH2Q7rPq0oqbiq/YCIAvJnPRe+UCKNdSp3nzdIGLlYu5rogVCXFS7ii98IokWg
/5lhld2I/4fwvfhWLGiZy3ul+BbUnyvB79Re0E9zBwHJuh8vff+pLwM1aEcLXzzS
OWkvX72Ys/If68RCxxD43nSmigZbcWQEMceJrTa5WHDPHlffFSndNA/Jg9leiKAH
QhA1Y20x0y5DOmk0luoDEjkcHJkelS3OEGaWJy7/tabYS7WjOMJV9Lhg+sdOE5Cs
PpvRJmGK8HIA513o7fn3PzmvceqkHrs4SksGD8xBdfhyfTU97cm54L6iLvyE2S+f
4f/x7Jo78k91Br0MxdwXTmJshPXp9CK3v3qSyyFIeIQN3cOTGjFo9DMJUL1Jr+12
l8NJCaV4j2KkvTBH01HxFqiEKq+7rtCI6ljQd+QdLT++ZRFrIG3UhKwS6smo3ATh
ellXTuzJwY0AY20/4F9MPlCVhwZWyjqBmlNIbZRNWz9r63yIgwu1I3KXI1g1wO/3
berqpu8wLDeRDKNG+pEu0o17HsYZRKLeGo5fn6KfSG2yoG8IHYnQsiOxoh9xa5Dl
iyJJ+5Z/3OwmJMNRAFCmlw43QeS4vYYz1KiWwEJal9GqAAhO9caL2GelUKUw8sgs
/ra3v74ZSLSNtMTceHIfp7/E6IkfPbIoZ62NRVjTR0XnXFoNRxH965LoFqgb7FEY
B00vPBVB/l6xzHVAeqdi6kOX4rbdA9fuK9CopFzG0yN+lveDBlsZjyYmMb7hNzJ+
QoSKRjOmfn/a/yvrKH1FeZoqyFSik+RlXIzQUJdQXv0llMucZe6xCXx9WYQ3iMI4
x2mup8dFL8whbY3smd4QZx02MoxPunhBnj9dMdPFItkyVeiJiQeprLGNRDxvZIzO
Qmts5H2hgVQqBikhi8uoBzT9STEurAH2Rc0pfcDfuyQZzcKj3F2mZzys9h9oNNKl
47BNsNVfYKQ/A8mZr5El+AE5pQ9tlFxadvuAskwt9Yb9uw/lgNzG0gEUvITZet/t
V06rk1qMz4Rnp898fnrM2sxpZt4l15n3cSPFida03U5hKiNXA17+zwPPQlFIC9a7
RBpfS6s+IRekPRnrWPvZwshZ0mxxC7PYj2wjnhVP8W5xVm3720NMtwinNIXapcLp
dHfGhpPwmVrm9TujPOJ08u7V5//V31eJ1LErZxrzWhNr8vXdkXwI3GAs9XnWf/UD
E6wUiplicMfFX3UF1817r8iKuun++qQDrajZvGtFwpnlalqsG+VwDFZD0mVbNNvr
j8QNUChwMjQbOvBx/mHg7BWo+Lkwd9khlUuq54UaWy+mU59jiXEUvnKq3cTF8nzV
7P9R8rMsfsCWPvMfIM5IypZmVsh/MZpyWhbMT3dujxop+4515xGgeRpoiQ3jRRyB
lJV8WbUM6vVhkDLber9MhAoy3ysgiDFSb9fzUeqkTci07tj8jGWbBaSNmgItT05S
P1Txq288xj/ZuIFj1NwEX1tf7TJsIh5QQwnxbcNURaVJwWp61kH1ZFpEthLogxDA
XrIZycqvnKD5sZOSXhAFZMejpiZ6CdibUsNn3ONzNSH8aO3DWo9L1e3QRGOW7cvo
6zgMPQtGo0IyvqLS8ZbHV9wiv7fPIS8JI9nYGNfQtqiN/vRdwO2W9QJp5JUkrEK5
FdG1itZzr3dU+1NlhYH+owATjnUzg+HzbptRKrXok1rNlHrntOLnjlkJzmEFraQe
3vwUyl+JEu1Zj9I8dh9B73mGf4Sm8FJfjl9FcDbihH6VTMbYdtMXS+Ve1H4G/B8a
8yV4B2V+xcuiT9tSmjarFFFBm3zfU6Uuj2/hBqczg7hO7yuSymTd13n6pdNZzJBa
gOtgtSr24IDH19a21TXKJU+u1iK/+fyzJsH+tZNv7EVNStp6rpF+PY+YYdGg3yXy
M3K/klCRyvmv4A/vu1MNg22AWONTT/+lRO206/FK4EJFq4rX9CUgDlCAVGTORlQz
jgAmWLgA30bwzuk5LHivweC0OMdgkmvN+Vg4912IzdZB51JePKeV/lSgpZqeWH6I
ZCkpRIG355tTjauMi+wE/ul9iHD/VMaon6mYJ/rGN4hX84LvLU5+A4fpJD3v3dU2
XCTPhRaSAky916wzcJyGwF+xDz99tPtcOkq7WuQer37AQQPNTie2ELlXeB6yIm9c
vj8P3UiWFPs9GPDXCzygTsfXa/tZJs5psfNZaRHNPzSyK8tlHcVf0rGLn2QeBW+K
Ipoq3QI4vY/pZENprxjuz5kOo94NHEqO8cVd1VBziCqNL7ex7lG6FLI79XMQj+/j
lPouxRH91W0y0OrMrq0E/sQkgRhACSC523Zo9jZjy0C/Y/ErDqME4yo/uUzwNA2n
ct69k6TKTJdnMyUeqecmpSDq0KEAg88Vu4RMOBZQt9OfH39ydAHi4tGFKWMRhx1x
lxrJgbUdCvGb8NqR6pJ1AfvlkuNuQp5gHsLseKY4mlkjTImGfqWDNaiDRawczDZ8
4h6fWJptz4HOJMZPuPLYGW8e3QC84fQADrRdEkP5ValgtoU7Ae0i+nJXN2c1/WsI
T7UtohG+8o4dTMhiPFW5x/ZTmzn9g9Z2hs59pAyAFvHK8j1QwJdgRBJk4jGsQEbW
7BDrpXKAkrf0FBrJgmrCj7+oAmQ7/8nSMyWzZ7ZQFYKYZP+MWFHlwW6vhK/MHLju
PjNCrLlq+cDhrBhEKwWcV00/7Syirz3NxrJJY2Yz5XZWNmtWe029e5lSCVUAoQ/C
CDDmHTaKko3nsU9S4AhroRV4f7mL24uallTZ8O+VY1uTpaFUgVoVBVZffCoUoUHj
pp11bhS96zZ7XbgqniXUQBoIKL1FR05HfToaLlWdzrUgL++RgpfTd1VX2a6/mkKi
MZZKirw03Jx86j3EY2Q7I+r9G2VRyga5Y4saFmMmAo8MnpM6WKX5UNpF7hjwJHa9
qkI3P1hOtDxXnS3KLZu3PDykyZLqNyO0FdALeak9irETReW7wAkeKaVbC/yWeNrw
1qB8gT+pZvfDQ6m08I7KjdibK5Oa1cksj5Yi9Chr5mCDSSJhxCytj9eKCgdvsKSG
mEERXwpqFngu+ymZeefKSJpXk4ed+eNpsNOhEM4fZYGpnXmdlVMH7cyNeKQo1VD6
smjO5x3ULjkw5v4Z2lr4EhEV1CpbHxVoisbV6p09kMqFbP0HRa+XkszyFLj75BjC
ELHUL+v7xPEIWPW92ghdfvLuhM2L9D0PGr2IFOmd8kLzM/S9C2yvcAur3rwEFwOc
W2EzPmoRxODZlDnzci1M46pYJntyc3n7chazKeKMd+/cJWjnjma0ikIUIWVZ24hF
RW+yLLefvR2WWqf/xH99XghsDKZB5eSimmMB2WxfgBKS18T+izssFUVLguOF/Ej5
RHKSpXhhsWydYZItQfy5UlxP1tMlfzH3WMnH9nzMFj0BO+SxKe74Pujnj2GrXFU4
Z38WgpxgWMxoPltORohNYZEoWVh9hKcgPP2lg8L3l5hZ1QYAlBxOJRb9kGBQkK3w
CBIHDMaoecQTVh0CCtQ5l+orQlbAJC4YCQ0BMPWbiesl30FzNQK8MYiGUyBOhFIj
FwTSHgPtdB9zViXY4VEwWx+kOjkTMTSMrXWs80rjV6Y5LJFHb6Figi+q84ybnZco
4l52Gb3D94Cf/ZweNzzlXzDVPM0KbXpQp3Js3Fn9DKomLbgkiJQOebnG4JBIPJ3n
Y6i4qEiBZkaWSlDA14odop+Qs7gqF6ni6FVAS4a7KVlBSVSAhL2HONYxgKYX2YwM
u4OZP60oOIFc1lTK7jBxc5YY1hhJykYdw81hrvXScb+3LuqfYRU2jHIQtkn8LExX
Uy71yA9ONtlszMDF7jSJ1YfMwAsMJv9OLdnSWK64/iFglzqugJcaiZNdoM1ax440
fA0kALYmm3vUIGfK3iVx56zJ1BPRB1XVrc+HRhPBIFZvTzX9ON/m1Nc2QIxxseRc
T3SNHv8P9CEjNeoZ9op1ewEH9eSq+BV2ce6hxSEFhGxOjHPqObyZA2Bzn3vlyUZw
Yvd3LWAN3BfQ4iaDgEH69K0dNQPA9Ko6fVYuXC4do32s3NxMt5yxZP43xbtn9dLk
6g9IIUv/24CFSWx5cVzCQbU78Nh2Wltwy3iMGuTJCfQQIb+brBodP1X5fhW/MM9I
xr39MkS334s0SWA6+O8a7t9crixlGdjqlUaNK/0VRTfbp2BN0QEw8naSPd4saLX7
msSyasQl9RYZK5pTTOuOHnF5XxVVxOfB4DJq2Txs6MgDy8PmDOVqexAJ6tsHApn0
JFzI0XLJ48tcaZuwSeHyP6dbjidJb8miyNF63LzLD2LlVpOAqj7gHMPeKVD7LKvU
M8GvsDjVnHATuKy/KLfBzabXLRCXlpL9/Tw5VLVMhsWMt/0dwXIMVwP8YLMpsxrs
VYwzFOAjKOeJ0tll9Y8Hc8kf099JFYiGvKexe8DIYand5aRZGTSKcV7B18m7w53a
2iBhlI8bB7xqiXJ5klnpKM7cjxSHivZ35ig1ZOfx6ZhXMUf4Sebqt1HEUHxKJOlt
4JMmeTDSXENl7ISRogCxNowuLgedetuFefiqr7DakDVQjh1CuqKG2nQ7TKR6IzGw
L9lyN4ZiTuFNeWrfm8BlPINqUgyduAaQlEpDtZuBxKgwzfU0/zGD2+LlJPdrgolc
ZOcb8N4m1wFddKUeZaemWB5rtFkpejZOngTDjEHPo7kWaraoDq+kZGfoQhDtN4Hd
ERVsZ1Ilb8y36go2Tt6LbirYoOkxNpKU3YYEfjo51nM+c0PIjJHQ+dFFzMlBgU/M
F+tzzDhEokSBLn9fnHXSO0//FcdNu8CZVxmLocTEWL/0hh3YguHdIV6urayAasZg
ely7Rajh34Vbi9rF5kSNhqQb87CesB3rLm4gYq8oSVx/6vkREQi70i2peBCA2fAR
wFh1zhKCmIZIK7wXfhn5tv1K+UXnVSGyks4K9IaBcK9gN5+OzosqcSLP6sy58s4s
yM38QDd5GWhSy57usth2s72jQKeAZkOTdcKmOEleNpuf0ZNf3mBcEz4Dtd6TEMNP
UK3Li67aLDOAJu1Hb6mVx3yZclUiaOWRbuyFx94URRCIVRDbzEle0/cWQ9wLYBBH
9X1XuwB4wxRjSxP0WmIuMpcjYjNrx5uN81GTsv9kEb0fOwVAmFxYmTcRblabrKjz
3MGrHmOgOUMLIK7w8DuyEfjLTbBK1OUYkCZ0mCXtfzdv4sDn3uWHyrCtFz09I66/
5aGw/O9hiUiXXs3nSQ+yORboRw3Lhbdhvo/3/c9oN5RhGmD7SCF0jHU/fjP3mT09
X/Oo+zoShRnGrygeBN/SVqylVeJfHekW72+DYwtRV23UdwQov8vndUysDlLnHqpu
T2mXBPaAHx2dyL73ti8aJYoB1NCDVyRxN7//kHdBPCnDSLwZR8oBwJYHpFjxNS7h
U4wVFTVQ6Gfc77LMEdIP9isOLbAY960OK1OfVJwiQ8rxIZLIqybE4GF2Y3l1RlcC
S1PXgzNoRzYYrP7UVeNhrh04BydtQxeHLYamHS1Y0JZPzAzrt8WKm3WU52Grd2p/
8qIlZDmylXqD6W80gs38e74mB04m6BS3ukVJREB47t9ZMhr4zBP5aQKzi/SwwaCs
8tiz+2kAn1va8DOHMQ9wGx7zrBCszlJDYdPT9SjzDXmioLeYXFjA56ylHZzfW3TI
HlED4a5Wlnkk1MO2d2c6w3NdPgF74eh2NSGlZIv5HWydpfEuvW/XAmPPZzhEHDr1
gR8Lcc8SYsxESowcDBk2aOy0Ey/smeCnAM1Dd70GGUD4QtWZ7uDA7oaW4itEhifl
iZRUlzCDZlEF+LYe+MJwGssWA466dUv36iARmtGYF4CSVeAUobzmXRF2CjGBnpWD
e2YbaN59MtWKGuFQ2H2p0QgIHKxsGUpqa9SjwWQ6kMU+NjFEptvSuzsa/iHiqGyb
mvy1gDOxD+4lmPk1VBvORJe3/xDWnT3ciJHVrf1deIEKEVvKDD+RkiS0PKWS20QI
b39AJQU3XMtYi453FhQ3VtGOrQVB4b+4NIDGsMvmZnd8CY88zgIZMwoRAiRzTjAR
uYkO1fi+A2KBq2WfcwLVIsVpLHLCj3Pc+tiK1Dz4ddiCaVzqQImjwPhMRrrjkUv7
TTlVxu0N4yKOINhsa52ktMfaKJV9pyV+4Ic9yMeXPeTNKoF1a8wbqu98DAYaN5eq
2nMAMkJwlO9hGh/Q9qnf4tGeq1D7IDfBsFSgc65gaoyI9ZaLECur1Qigw/Cz8mwg
AASspmwYtH/Bm1JKfY/BUhTngykgZu52+QZZtesbBtI/p/OSD6DiZ4lg0JbZZr51
P+++piezwUyQOjcUMZo3+ynHRyxzltFqqMC1lwfIa4NSbONYJGvWiQl0S7EudQhM
LwW5FoVUC7NcmUrzi0I7WSNQj53cuxeXNe3nVkAc0g3QgUIiKH8Q6CPX9ZsGHcHU
8daB52wvEoiXeprhDdTdsKBr+OQqMQOqVqrAGXJcIFOXdXLxU8KKlSu9+XbU86Qx
tfOPVO7akMKl002jlkNAhgHOtAF4xKwKOgkUuAcT+n771VqDgb7DYTQ3omGW0nWt
vNSGRjh6VLYxkOY0vc/QNi07Vko5qZH7X0UNKrrMq1kdGj9WObdxntlakeQ/Fhvg
7bKVKmfJ5Rwx9UT29ty0OMtCa747cI/RsNU8sFwehPTU6jUruijsRXZwDzDKNcqV
Ej9Im4NULKbgBTmMqsrLUna2gYrr/VfHtBayT+wZiz1fimf2VRmPhRf/tf/KYgHr
K/hIdotZCakdBZbs3yO1oaBpoR0UTkb04btXq9Onzkqx+SaJJpBgk9xaRU6+MkCD
0XbM88CS2PxPUruCKn0pnE3gGtFA5xpcD9R3cnNS9WLzXvwm1BF5v9Tw2XfofGRE
cdyI0hV1yr0OVG8F+uQACTfjv+lYgRqKD0CMZb87dP1i0S0Hunol2PvdJbOeO5mn
Dno2HpvAshNBdTpiB0RhB1YORvHM8LjSxNPO/MOEQcxGXSVFEm1fJnoWEyzCu606
O97LxmJNSMiDGJHBJ1KielMYdFMIucO4o3iRIr8ZD9dVB9YOjr6YsMnbaTCIboM8
JFOGelTmfI2cualY4fuu/Z7L62XexML0j2wLoY3JuNBzYuofouwvwA/QIAk/u20Q
Vd/g2G2oVQjMClVupmdd6nHXt9iaJc/66K0kg6TTLL10hw9EJxw6sw4TnUkcOvPH
n3HacIY87pPsXebz7YCSTXeLHz7PV/kjA3KdT6RR5+c/tFZHainwHkiUR33trk7b
y+++2sF083ixyX/jTEeSftE3PKSSDqbMIRp3hAi2WBvmp2OzmH3YuAkHYnnlkWnk
/2WZkxePzwfcohg5jnI1iIdTTOz3GHHxyAcYihHrxC1XlttoDCSpVGGZbvkxnMKO
iaHbHfVdJrpJjZH+jYWkhCfsLLMM27eWzC+9MFuD+T+h8TNzQTWenyuUxaYm/8xO
hGRuJCynHydPfKPlooXYpIKSM2oya6Eqmt7qeS6mcRjxeDcdPEQeesrrKkgAM09D
j/rUGikDlFZqU4Cxb0bU0XAGDD3Ue+XuxWxyGQnbC5cDcMzbiBGHWrdN1Z153/8l
8dhVs5Vpl2Sh6KldA2kffqlATGqo0rAVJwYx+LNdtbkM8jP9oVo4IHsBXgML//1u
NLYQvSPb5FFYdgZHz8QfTf7Q2SHCFsBMoT4qlF2bgIu+ZsdvpfbaqvqJg1b2oC85
redNtLHb43X0yhmpIjNnL3UgIa1wsJ+R36IZ+WkLWzKx2T7NcCzAd2Tg4p+imUi0
p+Zgk4+U3+jfWAcU1V9l9/RnhR3GMazA+9L+93YLBVm/SvGlBDziPr//1/Wc7bws
KuOcYqVnE3rR0kP3ywzkhND15pBRWSllx9oOc36WeXpo27N7dqX6O8VnHvkqQONy
snFLg64qGuwrkw90Re0CtCidvyKtTD7comnFnpaMCYqpWnWJgjzMhl5q2Boh4Oco
KutDQZ9vI4j9gcXpObBu0Yfyf4btp2pBM5AmUahr6t3Zwk6fupYSXk2EPLJvqpme
aeDcQl3hVSF4QQhjXbpaRI2JLTLib/sKwVTvyz0bu0Nxa3k/QKddQsPZLyJR0ObT
G3dSRcXY4ZUMXgkS/UtVIl5mq7bOCKHoSiFdOLjR3UUT1R5v/1WKt47uok0c06To
3VLT/Jr+jHH3Dp1Z3JvrveJwLXOJg6ZbFNMbPd1HS3Po4yKmONn9mgyvWonuiz4j
322EfDkoktUe/ZSxGFbao3VQ9ALQkiyqH/BZWT7Kv+ZfU+HUymO2jEYEzUS59j63
YBg9S91fo5yHk5V3zBuTYoMNsoTvwEqSbz8hC/Gy3x5C37gGkqU9B+OvXX4387QW
T43GbW0cuexetzLfEc0FtRTGiM/dSC6tUSWVcLOyrAknuxnZy09CZTjKl+p1KnnM
WBKrsNm8XwiPvwKmCRiuIqnorxY8eMS5AwkBEDFCn9SEBbwtWmY9wfF2JL4d0fN6
oqJXQ0HsY1FVbuzB6uog/w+PNlIleG8jlstsvwIm/a+WsNZhUNTK2kzVUOGKpAUw
3obun6gPVQiflpE8qf1s8fvrig28OBDaJxwW7+3ztD1QxfStetiT2fVRk10SjNn6
bDXh0hq2ROiSydqICWo6gRA4rMj6/zEdub0ryjRmv8GWxfTeRh54eTd0Hh3FqiFB
Q5b0Kxnr60R6augFwlC1Li/iLmw8ROJ6tsAws/c6WwoWrFbMKkcQkPdZkEY6NEz0
OInQi3Jp34VaqUxT+A5DBLmMzX4AD/Oio2cUyYeBlwbQ+xfW318qnCG08IuqXlg2
ASjFpAQaqTs+D5oW4q3onO2vgSa63+4Hi1GNljmdDY4+xAbEYJPJ3xWpStGZZxaS
bDwhoW4aOax3dbG/umt6ZqKiA7VDcix4gQZcr5q6KI6rZvNp/PhhUc2vmBXnGUVF
uDHBBeNWcmjRvFQg6B61gae65B1Xp8B5VN6aAgqPY2m2NEX3ESPD6XynUpm8wcIm
QaylxeYveUPO+HFxYiwerNM+ILp5uau75ArCJdqAxmwIPbIFIuKB5JanQp1yX5s6
gGmGrwERSM7I6P2yqVQZKkkwBxBjsBvd5BKe1PtAbO+0my+4O6NQYZ2u3a7zqytC
FckTSMl8BsdeF1VKtkYNEXc/XsbM39v7eXpUevmVZB91XnmYqlQ2WeHoq5zRIX4O
9764zcr/DcukVyqfvToYjkN53Xf93Z26Fg5L/8H445JoKflOyPjZxFOwvojINfDz
A+vE8LcozLX7xFoxvF0M95oQYpct5znimwct6LOcbPaIdK3yt/fv2shEj/mFSfiD
KH0bzt4fqFEbgi5J2JiuQd9b1jL65dl+pVvoKG6QE9Xbh6agUx9Qz5UCTRvByTPZ
6DhRyM6eGK2gsQ65KpNxDca8c/MbNXsKTAuiOSNlr2dXMv0+ozoOUqKfkxonkj+L
iyKAboX3SyEX80A1iUMq57XyNj9NMIIW06qfHCQ4Nf+cHcjNYm0TLiTCPp1bA5jR
CGEWXzXqMiJq/rWUfCYqloxq8nvdsauZkCEkyZ96PzPKfj8VqOHw9VAH5ZJXh8qz
+pNZv2xXjx50oM3O4CV9FelNdYF0Ju4Da3QJxcG0kNQkJCloBzw52wPTZxHcF4cE
4jeAUfr7AonUF4B849eqhGonKxHR5VudtWdet9CvAThO3vGEO6x98v5T47h/j4OQ
xKMR1A2lMK5/ib4k6XdzDAaWeqGcNEOm3pWZ23gNOJ+7nntHs/D9dN06HxWyvO+s
43aIFmnODxM9aua6LapHQ9gZn6k8HJ9PCtZO0BJTBJMnaFJNH2up5ej4h/wWYf2S
8hpCckhNmhu13B/2H/GuE29qWBs5EzAySKU+0S8dwF9D33P0W8HkNynIgPeB/C/A
9i1PRr4pxl5gkSIS15VFKcQ5beV16w9gSxtIn1uIsXlKn2uYaeO1IxdzhXt0foBr
HvX/CTQLG/Y5hskiPGspRr7Tsvox38A1GBLRsbwy/LaSupjdjmnBJgwFIeaJ3Syo
sYbdcMCtxupovoxZQH5nORtZmRzKnKJeLNRi0ce+YtIVcwR3H/dzuJV4ywSL0iBW
SSOf3lHeUQpSySInR9wbD6DQjZIhbaLSosJH7NqLGBh0CIKaPr8wnoSTmehu55qz
3kmsQjNxd3w9D36ScNABnS5ipfqL+SSnCPksXFtoMY4mtKSzcgMKP/ToliwSBONX
KQBz3Klz/02u6TehMLEaR/9fjsrR7MEILRBR4QyJsgVmqLr4HBBgvfxiKSMhG9Ea
TrhqsAfgTg89RAaYxG/V3t2gFjBn6D0d65TUPUt156q/H/D8A0lU5J8HfHjKk++u
nyli2dRl9S7sBAT4/z7bOaEBAyDH08Z5G1AsDeLxADEh7egYnQ0er9QvDdjp4snw
zZCP7mWpxSAY4zDNOSiUffWcvt4lpYUF/dwEOyn1DOfwlCI7fk037FjOFa1G4mJS
seoa/Ipu8bTLZ6QKZpHmNFT9lnuaF85DJ8MoVbyGY+mE4pfCmf/Wz+y+z5N7McUL
f7sRJ9Kid3dB4Kv+OLH0xkiqEL0tZiRZwOKC/K0YrFlhn1STpV4/XuD3C/DA4FHG
lLDALmj5PWF9wKbvSWoFZEauYcv1u09UHwcSYdmdaLU9VQZRO7e2oKLLeq7fUBd9
x/9RFcqHTiRAwGTod7KROUtaq9wgK50tOY1dQvQZIYKxFt1tvVs2TEsNYDNe7sJ5
9iUvNjLgBoqpE8L1npHqXrK9bBQW1GcWbD4TEsEht6a7LFy8KgUd8GBRf2BtxDyi
xxPB1vMa3Cc4ewKmRmT98YEgXBS27yvYxYMomlDurvEbFqSf8qiIOWhVcgs+EafB
mBmNmVNKw39yW+PP1gRGo5/I07r2MxKsT91SicG1KGOfYiuqE0nejvGR/h1urxLK
iPxe1IMNUu0t/Ohpm6HbkstpsukinapO3sAAYAoLn8mbMkVRWZm3E2fw1F/c7sK0
yP+Jp+lmMCk9EHNW88Nth8K3Rn2uqkRJxpbmI5m8yEExH/s+pomqbHmF43OmTsQa
LEQ6Qg/eOYPjUSoWGBDtEGZ99eBz9hUb5sEJU/L15Wv6upNrHK8u1QbJuj1XI0N7
b6w9Y3fcc7ZWeLd5kEhclxg60dIbis/RNyFc5cotQi11vYlBNqllwZo06B8dg4lt
C+jWDl/Jd/vuEzQ3RN++zESdf/RFTV8dt04oNxSz7qC5hOxj4BVFhWiVZEEd5t/7
Xol5Rf7cLnTbMZMXbuxuQsvgJ2W5D/CdFKX+oKRNg9b/y/rIhBerFblv0rY+MXzv
CS7IBYg2CfnQzGUrzgdKA+16HkvWIqve1M0Hcw+eQPys5oEmw/L5HDgjAOZ+HWGt
Xt/FcPRnbWyeRITvw6+zgilyUXT1kZrBwMIKQXylFNTgk2rh+LNfOu4Iniuv242C
1OC0gGvyGsa9fUxJzpqJHcGBbIW2Knd1gw24tWJ4gMyppLq/6XFoMvyicwbtDgP4
TCjEf0WzjQpLbDLw8ZejZwUzMu58/dTjCOdv02YUUWgFwOpZ6x4dqycAoHjyFZdT
Gq2iFLdY78IpKmCP6ipZu4/nlCySeZjZgWk22KXkyj4yHw/PUOu7xGxc+b8vUzPn
BeTZD3qZSExSDQuZtWSIaXnRqZcG6E7RBcII/1DXTw+J7JmIGMJExCyH1zHHoeeb
BLFjF41v6vyW99PW27R6VD68KSxwQPRUyLVihhnxdWWrdZw2YaYIrOfzl2lD9KR2
8Rbv7doo26L4qYcIR9zbLrz5G3iQtzDmAonHUbrYfEXL+Kz0ylWltnZchbO7PUTl
WdxNTnP1p3q8hggMrF9/iBJ2zxjHhfAyjfClN6wMdFcAtrgGVtmG5lC5aKCsjJ02
VKzIuwYntqX1kpY83f6mETWYk4/oPognCBpeqzC4Q40wkUgRkw2IQTpouPBL0wjd
Nc1vcyaoZPUuAlqzgl+oPtmgV/obnjEjEYqEPF5mqxyz1NWBiiOQOv6yO+jhwsUy
mJGTy/305vTTN1NIzNKQ8djZ7ElgXHmpRa1KffD5Xh0gtF+kUy9D5jxXzDAjo8BS
b/P9y5vgCKu+pO1XguyWWjA0x/AU7tYkaFJmv5di/q0ER8UFUl+pPgMFTBY1DzI8
3Es6K9DWDRLJBiFLejDmg4Ig5H9elYyQg1Ld+0LdjSAe+uL8lHh4bZ4/Mo7+YtmF
cA21r/NrCTQ41tr4QeWjYcQA5f5bc2GR8OnVooPv5xJz27eDZ+Ldht0+C8b+Xvii
nexxTPtONWoDibIBZR4bbgfXySKPz9XFdrDks7f2feAhmP3+8SzO+xk3qJV+w99F
OU9WXKA3yHB80apFOjxuvgQErCc0hzrLpjPy7T0/4gErTfgLgNEki369sFX+BpYj
brO2He63IbZpzbqWXVjAnKY6cwMvREhiKdLrEPEd25mFkU9vTqwJDVtpSfxfTMPU
Qmc4rFKkcVndNjmI9tl+rwdmgsToZ9FlQf9WqemRl+ED24Op54G4ClqvET6jbEKC
IWNT1NNJiQd6x1h2rp54g2BDMOnAZiFSZhCJaKhWXEh9qW/vXs09HEAFuBWew8tT
XZnh4IaWJr5C5ib7bZV5wh+REd1cpl/RrZ4MzT1cEDbI93SsG+fv6ei9v+t1aaPJ
sPVM7kSc0550P5S4IoCxZw97b5gv2Qxj+fHs9b5zSBpwEG6WcdyauMc4LXdttZPL
ePl6QPYasT3nxjQP1qrZC9UQpsljYbevzoiD1Ytmrqb3FL9Nq4VsCrnvEbWMaYJg
/Xhs51ySGUhlaonhK3+rk8w3woF1tqy6JR45gaQfhh2rtx4mprc8ho9mN1QSKswn
g+rsi6CUCpaXE+ynIGUMM3LCqFMOx9btsN8JgOX4XRtuVicwaRIAKqP0iUTTs1hs
xmriKpxOarcVyBUa/nb5N8qvdvEPR0jI5UHqNuPc6SJSsbVatVV1RMYa6Kdl4P9d
Ieub7/fxrcZyVcICdgWLvG2xZAJbIr2qeZi4oD8+kzakA8ZeREtiD9We+MVcBK4T
XHlmU76oQkTcS0WYcX1KLqeFEyRc4yyEA14p2wZ4ZxMaTBcmfadWYQAZfv9hoEZe
`protect END_PROTECTED
