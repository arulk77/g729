`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNxeY9oQpmCXkW4r1atYeUttgpGEI6HZFC8jE06OLeq4w
eKV/8gs1nPUuPLGdUHiqrnYXysmnBofFLlbqVyZxjDqRyB5PJz8wDrFloPHlFFIA
lEVYQJ87EZVXKF5OIISXblT3v25yoPkIZAVbwp4wWbsvuX1LCFQGcy/gc97DGDr/
zC5uZuSy1oWdk037MULFTjc83F56x+oCSGZWAKUJlZfOm43qDedChSn1sOYb6png
1DumcbQFbfJqp7YubIjXFvz61TX6iL5D8RckB5h0kzMtR7u6+w3dJUCuBGILvpcG
+6TJZN6P9Uggb5qR7yKSm5a6H2wuPoaj1AeOVyDA/b+o2B/Xmv505f44k4RWrZaU
GUT7ROyeTsCtDK4kDFsvsAurEDqzNsnSIPIdt4dwNSxO4pDnAE/DE5I0qBAGJa1+
Hx6kY5jI/MAeNbWr1dmlaebdPyPF/5GXQfsfNTOJZjkemaj/8GTGR2R0GZptWeGz
f5OIMN/NKVyAKhe4M9vDBQcSO7lLa4EfVedM2D/HgDL5axCB6Uj92rda47Zmycap
7I80F6JGy75rSCaLaZnZcAQe9bW1UXAMtH40R8t8N94t1LOKRdYo4YcCQc6ADi5l
l7kwLhzybMIm0RkMLz6aAnJpETHRqSh1TEnqGdZr6zhc62N16y7RsTcIVJSY/Vxm
YAiG2Z7K9ZtfNsjm2D/9CNiCzlidC9F00I+/fln7ZFnAB+kmVE9XcE1Rf+T7LIt5
AjTbMJyj/bvf0kVLMSZt2MWmDJtJDsF2reNTswZJDb10rBwuxkn46uKYEJ8ggHFW
DV1JJ1eCt/TUcOYRcnL7H4waUqcn9pBpKvnbFcS3XXNgt2lDHL5BVqE349Zy+o8R
m0z1KqzY3HOwFl9B6ddXfilUwSiIuSSHKddxPFoFB0PE73Iom4qUXGdlHZCbQ4qN
ZIzJii0b+Qib2W5wW0aLmmv1bxdiM4PLrYAlGDtZwmnvE4jeIsQUHiE7ahYKhIls
Xde6B2VgCkAF46lyL6jGBnw1+Hvi88F8S6/vdq5ufSxKKt409oOiall3SAPNgsiD
SFHp/vX7HLACE1nN4t7fjQ6VZOiRLKctfm9byZHmI/T1CoG76tFHReHooIW6Yk7C
tP2pSkVx1/47YCZp17JqDcNbVhmEODSGjmHxfclb7CxFWga6guOtEeSG363Yp1Rz
DLEV/XndhYoMHrNfucNxm1AUG4csWbQEWL0CchZoAqy1vYX4YesvBNPj/NyIfWOp
/gC/X8Qov5VC18EqhEsTdpnER9o/5xyxyk2Tiz9gnW1uGwov8qzPT+nQ+tLIjGWf
olPkn9FYgKXEh8lqE6Vq+zr8OZxEDfukJmFlF+yYBuwF+BuRg3gRUtZBRjGfzqF/
bfjZONQkXPCMoj7fKqKDHUxGpFxhyZfF1DkEFbAH2kVzIYXSqLKYlgLyyG7e0xIk
qUEq9T+TeNjeEWbdOyGLMCGUmr6X7AM1xt8I5gDNNVL6jfj6C8up9ya1IPsVHW/t
oOx4U0ji3ujkhrwhOo/owqd+OFaHySNqmrogWml0VMm5SofMokPpPMqCElFXuDjl
qqozX3R7KPXf4W5NElyDSsn52qpK6GtaWepbe2Y9xIA=
`protect END_PROTECTED
