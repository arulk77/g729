`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
B4uwvAg3LkJ9lZO5eZPoKJE5COCLvlgYteGlHSos2b6EJjnzYNdqLWfbj3co1Qtn
T6Dy87suaac/+pSVxo2BcomvIsStNvErtKfoptAfNpwwWAAyIoYCOvlt7b5F9el+
44bg5ggu+EIjnlSen8Mx9JbUrpE9mFcGQQ+Fqg/onFzffVdHxFdaamBKYt9teVdK
zZoUtLb9FtsqOuMayPbt4zpU/uRD8BZUfSZLj+j/rT/DsQyzdeBayiYWnaqXPWam
V2ibqSqe5scciIzEn/63aU3kfQHjcKjdjjEbyreHuIivHin51+9jG1hrTR5vS+Jy
sdlraHuRzN0hjOTN4B2qTYZw/MeqmStE5qJyvEfyLpYhPqJjG1xSVlDF7uvvg2Qj
hEV+IykgyC9dM5NrP8TdRkCgx1PVZem60LYzp/2j/xGLK7vdOtifdOpHVqKitGmz
9HfuEDv1+AxAlwNRIsLsbIUW6MyB++Ge6KQf3YJre44ynAx62xNtUPZJfBbhJ4sq
kerDCr80/G4/SyIAVk4LXg==
`protect END_PROTECTED
