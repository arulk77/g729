`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aYCqwlcvJ2LozT54cot28F2GHY3ycG507IA+AxFSp2aN
q/IzywAfJW7zq75WnnNR6ZaGzJhWJfjtcrTy0kVg0Gj10hCy0OTdrYzKga4qU2eB
8/s3dHuMeG+bPDYF3Sh6lnl+/h2bVn4KgHs8DFNR0PCoT1S04pP4eR3hhpjkILe/
hTYLLL1vLuySWdWjj4KR5ILKnrBqDoyniYPn10E/QhzyMreuV7GXlbRDlK517LBy
SHGI4f7D/rFwd94cT1//kRvR06u3/SJWMFDHI5im1ebhsKNDMQ+pNZj5qGzUxUE5
f3NZWJLVE6f5lJo3jIpPI9PxYjNECpIzcBc8m/nByhBujLlUqcueXbw5t1qkmlDI
4hdnyDw2hsoPYx8dvjo26EuycBqk7t6JNTDRHQFzFqTeE+81/JvciDr/inPDdF9r
j5RznVmX/24XFPEKQbE5SApOBz/6rplws33QuQnZpkiA3rKdhhhKrTT+7aQFo+9a
E2xCr2J5X463SRkDE9fACCmA4Z5FPWAexSSKll5wne9D6gt5OiTYQaYKP25OXd0q
V/FzrTtbm7wny3cXI57jQUpK3vkcGJhYEArnpPD04cUlLrQZl0QzkyQmzX1rO6pB
jBW+wJLHw0E+Ht8s2kHqE0qSte7Dnf5T3h1nbpAzXOEXG4rkjDwwZbFCdeBrFBW8
lBvV+UdxB8SuncjQl9uSOUegDVqx+AlE1Fd+pBBNGn15nzbVNGabvQvVVX82vWKG
htkGfPBB5m3Hg/YFuvkxC4OwkABX8PdG4Qmswc+pToTurHrVNCg+LFsAfPYc+UW7
WxDdF/Mg8OUD4MlJN4vJ3mGupYgmFeG3HO2v8fOMbK8krYzuUZHV7kwbQEz0IYTI
RXnBMMVS+1zc3J5cfdqWynzh1TpfgntBc8+WUAXctkH1DblRHdwagLXZKA6AE3fG
TMy94Hv7n5kX1XYQ9hCcHI7XI5eA2UvH8IgzxttmUvyucdS5p6eWkNAwQrSjssyQ
7ePLOwB2tMIvOZxkWkqa+iN0TcY8+I1ip/ZbrW4jOHpFEMsYO84w/HJ/supgUzNq
My9tt9WG4sw/gAr+FX5MUC0HoUc5IQELGD60CTz9iDqyHajAOaMWbCJhMnbK2wib
zPoYPJTtSHwg8xff3kDXGMmMdBkoF3zbCRYfmOH9cSuJUqqdfyK30PUHbdJq06eJ
BrrJL1BlojRHzF9yWOpkUuBWol5TRfGY5jxmbz/jz60V7/NPB6ZWZ+YYfkB8xYrz
iKNElMLMb8JreH4Fgl6l2UMORCG3kbl/wGwky7RPbDzgaRwf4YHSVIkS/e480s2H
QqnrBYegY+XMlAox44XEeV7xb5njcShJzIZAUeaDX4md7yGFngiiQn5MM6QLluC4
78L3TIzU/+1DM206v4gPWIl3dlf4KZ/nq/dt7IG/KhprHGJ70nFHfUPnoMulcsvE
doSPHelueLOoAM0TmwavdRgvsHEcwfGRV84jPd7wrtQ47HyOoNJy+13qsMtadTxG
LN6xF5p/Uh0OKEbEKBcuFjGcLl+KzIEGoVY8tNytQTnSWmwhcbNAd5lbsiGwsCxc
ytaBKNOTaJQRIK1frnPr1/88rqIuUwFyQ4TzZhlW9wEJZQdJ5Nh31n2fM3kWZybA
ov5gspZ9yqGk22EQmRZy4NzUY0FLyvHXI98CZVV6seA4dzNXcRJ76OXj4n5ncHlz
cRjLi9w8GNRPE+rwzDT4ic57Go83LvVOTG7iPOntL5uQNBrY7X9XxU1t/1E3TJ33
FIVxsxf3dQYZIF89KrMtu0HbOgqodf4mqVS5AVPsNFAO8SZCXb5WPq6J4zpPXrtM
cpbGiWejOk59KT9fgdgeoiJfCbREh52vtP0nhLW5eyVyAYKI4eNFEfnx/HzRaR3K
TgKRf9zu2yKDnR7ZdIxOTcL0ZprvfFJB8YTS6gB9TA4kPDb92oxZJr4F2tTU6EIs
7Fn+TOHpx9ZbmevREe7DD7wOLC3HY2NbfXzHisijQfNgIjuEefWcapC2VWJBp3rM
t0hOEZ9rYvS40/z3Js80I4NuncK/Rzj0ryH3NblDqRu6C0dWkqAPrYUNvdWBTUol
sbzFAhoG7z+AC87ds6lTdyO7E0zNIZ9GIj86xgO4IXguiYw7aNUZhyNoFlvx9JCt
h9R7CTYiTtWpK6XDl5kAwDAVpQ7s02QQv5GCUkLtBgRANJ3KMUvwLytS7116qUX3
Q3f/zRaceOSZxc9w6H30WY6upfkM9HR5FhyXvnnRBOePNuSwQQ8+YwnahWTMCi1O
fZdYYqPBjoWiMwJvUUo4//W/vE8wzLfVHXZkGKnclzxcb+VNUxWGhowPKI8R5Khx
XiuQki/vv5ORMHSYL+4QF5d1kyQXWbzdIee3I9lgAuJSm77PPyqsO9rm7N3oppQi
kU29KKPnpP9L+ljzP06DluduYx7empvqnxyKr1rpQ4LBGzvo00+j7jBaS0PjcPXA
FZROhJVtdDcq2EH0lKDKOFAgyVpLPaqTAsPabKh6dMbBFouz9ZPmgIZNgpYZbjhc
/75jrh19rQbjwUojJu/3n9OKJwjV3u7cUFiBwkbR12k7nzh9vM/Ug/95BiyWuzxU
SuuK+321jZZ+ay9ZjMxqkUQ9+VkP+vtx9L6pjAB8ifM12CooQK6Si7hUF7a+EhBv
WXm/fwFtCfcfnIOXB536uqHGyG9t2HW/1ifLV5FrNOohbdAVkh0s5tR6ccwuWVA6
OfaxLPz1xLL0g3iEdg8OW+KXgRFbbC75SN5QMerQDSJ2OHSAdjPaiAYN830h1oga
Cc0BeesuKoxlLW0Z+bpktU5SxMGIveVL1lzUb3j1GTTklPLvMZ+QWb7btT9NET+n
d3Ps6AwmV6nCynWuvqVXBhyIYt590cjXrXDW8/gn47xlerxRzdgF968y0snv72Hf
dMkp1Cii0PgZZ2K55kfag5lf9SATifbNRb9AYmofAvtua/lpbhBWoL5Hafefw0Bd
/1/3pJc2uHDPfXcDkbfcxgbQbbYQ0RQcq67YCegfRJE1WdNZ30XntZ/jQ4q5KzN8
40rAjgmlrdkmT8Gj9Oh0Xg/4CFKX2QMZ0+n1Exm0+z57xv9y1NtWnOevRm8nfcvS
KQx6qeSVmIz94Fnfz+SeTPsrWFktfxNAiKrp85qkchjhKH3fSg3NTTOgG7zbfybH
2UesA7bb3RzqlTfG1C8I1AIsRt7knCE99APY49YQcg00A+AI1PlV+UzGT5neVQyI
EHc+1ER7rqbZquSuVXO01/141JdWUNaWyPklQjnSIh9oLnU5vAoWfRsz59f6acDa
/cc1wlwLrp/l2lfWC+su/m/fLq665glOh0P9Bo6SJfnNqPQdVPdEwgv+i50evAkb
MwF00Nqk74uo3JAg1Q1CUXOhnKzezcQsaB19z1PCLLIA7c5n5Ko7t7u5uRv5DTjc
uBAXF7Ck0zah7zA5XZo+sX942CVBKAZBfapLJ45jDVH66coixo0AhGKZmFgX4jQj
N8P26lEZSI5kBE777bA4PuGZ2kPkM5kPFdChRXMMZErdELqaMzvW1jl/R123psty
gaN8+pwsTzcRj8iRDNu+h7aGgGBd+R4UDcVrgoFniv5qnajkrVQ1aQHD/ch9Y7hm
g1W4BjlZmWS9jm6Dypruxy+DS2gIccRk8L09A/YRRaBiJxtaiLSFc5aamiWxYgnx
YPkVnOMU63nz3RW/cGlN+SK3mpBUV5i3EDhIFctz45wHkGzD8u8WOda31BWIr7zh
G6jQ9YY6wAmBuyDKrK3V7Jq2YZ7y7mGpbtVGF/1+aBC7eV0tCUYJc+A3ptNfekm3
8o5YdSIfbv7aJq+In1odknjOsI11GCDfD47dfhc50+3oUrPhjjFUY27HSbTC9luG
2i8TwT/MiFiyqARxj0Fzz/Pn7LdG2k1cYDpMxU/88+jnvt9yBemZagewVxkNkcZl
ulyvOoCtDPNPGIRL5q8b7oAHoNMK/Aj4L/pqljH/fsbRM5QDBJpgPIDh5My5n/FJ
yV7f9i9y/cRwl83HpYYpTzDx2tzAP1pJTEqZHGgAN461Iu+cfXegwXjclUh1qTJY
Wi8vlVrupejcgl/pyBQbnx1uYIfUB9jP3OyUmP3SVuou8Ny6mEiFH8aqq6BsGvT1
+jf3qM1shfnIBv9Rl35W7oCfussYwIQgmigjNRf9wjJMwKNWE9vmYmmzbNQD8lU3
iqWkeoSuz+USEzB7GQRXzDXEeMb+GUF8p+I9uT3x4dat4oZc/0jUQREcHo1K/+DY
tiQFLwB68DF+4oj5Wz72cIyHqnpvLwy4/c6oAGhXTQM4RpzwvekjBQU7Jj5++JsT
wbgw4gJtEMeq5pgEuBQYiXWbzmopk/U76GkO+vIF1zIrU13PpgHALbmtorJ3IazR
bXmSs5RLdhUYQS8rP+GCE0eAdmhP5ve8KLuvKB4D+IcMRvkWHpK13Jd19Jupqm88
bcVjJsPLou/CcTv98uH/yb7IPqIzQFV1a2wFXtkh/3uRyvZ1cfTjMf1myOxW3kzS
0ZBrfS8qDFIA7oQGnGPG5a0/iAuPHZOlMlyNNTMpi9c7/V9/H2rY5ttH8Lr4GMg7
6rACOtsUfwwPmlS1tCnR/MZa8Ceg19HA4LQcpnESo+np5WdIaybkSW0vJ/h3nyNH
nZ6a/dUJvIIOSNsb862D3g/cHFIjMVSh9Laz4KrjyVdZahqO4JTSkEW4QbYIUd4r
bDyTot2FYTwccKXe2bnv0TTAb4/iACL+pCvlnyFn7gH22llACWHERdxWRgXYfUH9
hYsPbW8I55UQ6dtPb7S+sbojv5Fqk3ZUVNgr7P7pErrpA6uoERIxLQvDqyeKdv56
KSUESNNhalJ087TXJZj27z1hbehJwR6Pbhrm2Ie8IPljUlh2bKwj8PBi9ThwnocB
b72MHY/83IUN6BVWT2HCK9kB4GMGsKSotzTwnkaKhWyKhS4Ggj98ZdwYcvDnTkAi
oWHVKEKsBTdfeVI91wGLF/2DUjXb/GdGSlVz9eOk8QP8OjWSFlRfe4C0Im9Sjb2P
+bjutQJno6MjRhMhnU1zF7Dit/hQv2cx3n+uZwQyf47dbw9fa+pgdhkJTKDAsQOI
n1we6EkarjohSsr5JcezRiZlIfA0sQVBw7Uy0ddB+Ak8chqxQHwBKojrF6tC6ONe
rtKyUWYADFXOCqeDLze1HzbAVpmhdsz2xdwoAQd+arNRx+GSDj3EAowNb18uRGCQ
pdp7EWXf3be7e2KHMvouhLY3wsCiaeZUhbfQCYazxq47kmseVa+CHhJAiITkFnuw
nkgt6lOsEk0fwTnstaWiVa9q87+ynugBznkH+q69/vQgY9FTwP0775JEI0YFbAcA
hUGr5nL3OEmdufKwp3ADvP0Ya0U/eNA83LyN97GiXXMmVMQtGi6GvpMD6jGwfcaE
G10Arahwd0ONqADd+waur3XGX4b1+pwE3OST7Vyg5ZVaMCmgLy5enySe5WMTyIol
/qk8dPASmMA/2k9VPtxduVeQmAwkZdLmvRtMJGXwMgN8hI8AOMWqHVCMiepxJhbv
HwkqfL05G/eJU3+GQWy0iO2ks5qhA6K9xVkq4edPIz3RqO0Qn8ux3c0y/PDFIe9A
WgjLApXmWKe99ZngEKCcKTSfQovRx4micmwlB8eLj20Q9xH2wcq4BfjBYTRLOc/1
uj15xmF4ayfWxK6ctq37vJ0/icrD1Z36l0WX2Agp1ovTZQTsMqYUYm2USNgylref
KIC4T2IMCA4XV2gxJWopyHG3cDXbAV8TvXmKFbcw8h9NXtK3nmkQLn6PPhiGyy/L
43hPa/FwSkft6DpLXx3km0bZn/wegklpn6cHYzUWDUx/PoPa+AmgTs27CzbH3CfI
qABJ/nxn1sRl8C5qgkzN0TFCowa4JxHY/l+KxlniP6c9L7v4DCEsoJsgtfwMPRd+
C0pIiO3zoRnbybmbffVni7yIGRQsDiIdhEkToOxuhDMME+hWpUnB/hSlmNQ0dKRB
IkHYlEPVuaAiTHN8u0pq2t9oAJpCgQY2p0pnZdxaZDmH8ELBTlElRLEgcj6Jvr0k
/YfCIayWwg7VbkIy0HvptUsk/72NLpATneHFRwWfwKMQeYj2WaOQJPNOrPlCX1zX
t3OG6YeUMHIIM5j0CvwIrNp2eulSRgvXt4jL4fGn6bEAKz8P+gc0qDRivswcNZuK
YufWz5F43T6KruhbMabOufo3k2BO7UNUrw9VDAyErKedzySy8T7/O31N1nf6evba
5IrYEbAo7VT3H8eOFO+VzFKfijSvs1vWBuoF27de1bSJCg3+wOcX//M4nQRDb+o/
rKSKUAEFlcNyZni5Jp0m0CwbhnF7gdWEe4RcDhmQOQXhOf/GrN9itTpibzo0M4Nf
W8IKt80BVxgAgXXgJUVctnWMGxkPZ5rLa5Jhw25eMrRQTLz85xsFWhu+RpncM00k
vxa4s+J6MKlXDl+Z8rKF2H82Oxm31TB7o11s0ZQnxxhE8dQfwTO8K2Wof74/jM08
8+i2FNVRGO8iRgJVUdqzUUMWqPF2EgYMOe2cOdw9AIUEfFY3L8htI7bNllnnU7kT
aUdS5lSFfqgfafhQC+NpTMYYX9mrJMf6dZ2Tk6uXDVUumxUqXon40lManqBfk0hl
eofzB7tYr2lf7acIFK27LJQwm/f8GA2ncacyowH4Zce9V6/hViYn05MAKyh+mAZE
xSxRgpZ+S8x5liwAtwzDkHmBowyzve6Ynb9h9DAgoZhky+7R5+OPe799LAThmcmj
wPTvg5KMxBXcDdZIg2zsUyMDUhtdhsNeVPPlzV0Vi5lVWOKbJCZ4+zvoptrAClG+
qlIHKmuJwYnXScI7mElpl0j1T7XpuJHGrH/M0bJl4jOlwdG2HHL5wktiqYEysTIM
+zTAjh/73rz3qx9SjzLeyPquRQUXQYf9wLg4aAmgqJ1fItkOOIranY17q3SlAmQB
IxmZ8lOtJCzNTCHcyFgvIbapN7OovHqsWoFreYcTw+h4ap2uTEr51fvJUpTAUbim
bRNGx21SLdFjYKLvdN2tCoztb+gf3spmwy3pnAGjvnKV6TtVgku8VLOAGMHJ9MO6
1qT0ctgj9skt5JvAeKme47SaktsIRmcBcpR2pKJXq3bUGM/D6O/H0w3z5qniaAWP
ZJYT6meQ4rBZL94hnUH8SiVy8b2tV/y2Tf+7ZSfghkJAFaNzeDvHxYtq9K2Z3QAA
aVkTKXFjhyiMC4sR7nqu2PbmNufqhG2iX3QEEsdfie88H3lpUc4KgECAi9TqseaE
s4Wno+6BJ0F681U6KiYfim4jXW15UKM/q1cCIuoa8kroAKXyzX/++8HWtj020y7R
Nik4ZJDrcdi7tAPIEHDqLMy5/5IRNJ19I2XnKAmzq4pQYVnUH+ESx6SBNUcH+ffW
oKJOgTuaf6nayYGM71BPEZtVdA5P4Nlg21d3IxFM4rGvJ0jkz4iEslDvSAHH/csF
4WP6XV7Mh1fxEehus5SPIg6y/FH4sBjt8V0I/dnJOBOZ2u+6Vy+A7Y6haVxND1HI
g+D39OpApSCb/R5YYJL+w1sNXyYzM13KHpePhwSF9d62ZN/cuk1TZVfEXqCuor05
mYmRjzZw1LAuX3x9b5eaiYLJCmQdNHMBbNJd+Wz1vZFFHkDywj/XGA6nZiLRMy5h
Vy2vJo7LiKaFivNbSqOATxGY9LDIctLwJ2uXeadhE5YsSxwG2jmtAXmk98a9c0En
0qbVxzU+9Wm84XdT+AkOBCPM2XK8JasKWJyoHgH1yEB7G1EYZa3F9TA/yBbn0s/e
WBTKUPtErsBqEaA2P1CScPiWnf8iafi9+gyFxvnSKTB848RHors+5XtA2zRCYaxP
cEBcs2OGFEPNDqhcYMXBTHI+jIqbns+3ssqmC8oU7xfMfjbZnUmC4PwqdBctg5Js
1MUrFsjAi9yGUphgwq0mbzRT6HXQhXtR5G/MvlTb23O2/1D6B5hMbqJ63XYxcaG1
xuaGsU0IUdloRoZV7HsYKbdgaUoqDhpNC8Usy/mxQr/MoT5yJpIH01UOobye13Zw
mJIRgGGZ/m18KMZ2o5eHp3kbc5GdPCC52Pg17hYjSFMIV623W+IMwJGxXaySVcf3
+Nm2AVy4/dJW9YHTpKLBP//nsGPmn5HUSyZyrOJE69XQJDBRFDxYSaiXhQ1KJAxa
+ssl+LKrIRdR3AOxE17P+HKG2bgpP7iWJK/2PG+8POTbH0MCzcKeujFoUwsR/ot6
i3basV7EioZ0ZoH8vCqTh+0bmch2nufQV3a0/CMStj+wq5JIZTS8b4R9jf2gJYdF
wEn5LnKBt609u4kxs1XTzzmoVx95q3UkPDD86XhR6YWdeEkmPVe9RDdWk8x8myRd
n7i3et6NdwePRxKE1U66XWM5lWJj8CCmxRs1cnufi74TzhTOuzYTdXcsDPIhAdHP
aR986Jf1zqYy9z/sajdFRM2eYy+8nOcyD59EJS0WWBTA0KnUeCKUVVjFeXn2Q/dI
PowE7PIekNRzJTT/XMrQ7YcviOJ3oxVBYFHNXSz1QT5PlzYbIgPlRHLNh/MG77dU
pz7sQ4LPdQe1iCqDRw8f2o8vB9I/A7/rcN7PZklUAqw4gQgOt6o4666VvPmdn9YT
f8dTjwJs8PJy97e6yaPTrjW6nSv9pMITY2N8ljQRn6WeEe/BBftIvG6dIPt/XUtx
Tq2UJw3lI9xTD2iAlMYdOBfeUc5P0yunfqQX8CRINzf720CS0bc659lFbl3PrWdd
9DX/rWaVr5PzmOzNvO5eKv4qDRare6KrSjarSbNpXXwMrai9/boVWEBi08ss8Wv7
iKGhEAl0F8tl0TUuJSgBQMFOjELpKyL4tBsco0cYWjE+nZyQuBI/85+kuF8HlUkn
5+bGlgR2Uiqgi+WPF6+ICFIJXGlHW7IesEvvQbYO/3yGDbEudiCBQQdR4agfa+yq
CQKPt39jOHJTYCkSo2k+F/bB7HgbNWiwJKK4LR+xEx5F9+20Naffe7xWaZ/Cd+Ps
560+26LNTCOCplZMgD/PJWY28DCtUzevZFgPvMIHdFMUYV9XU8K5frcBbh0IgVM9
C9ngBKdt5nT7xlBB4N8fl793a5zINz2N/7kHdI2Ptg1CNqEyH13A/o162KPIlbqj
JPEJncZGjTVH8txjk2Rom9ugCs1kboDarQyUW3D/4EdozJ1yfykjQwqIk6VP7Sjd
/mMVW3bWlTo9q33U8sDFhrpH/bLkbBAxWdnd0ZEjjmDAfmarqFq24UKG7qQYEsp+
JIA6leH4ykFJCTFimLdT4EPPnJ8aANLOuUQUOFh35uiU+6w8aQ2z2y3N0EdBYwMp
uKrXj9j8yrqa/4e3XG7Y7CC+IFk0+L0IBEYbweYKorGyWG5t4PEVN6oakW1VQeBH
daJ/069EHxQyNOQvQ3f8CfysUt7Q4Id+tPCFrPpNcfiValaGERAq/4+D/We4dFkB
0mxrBtjg7XtI45vtIMsqirm+59wu6IVTWkqNcMrbXyMVTz7RTCuBdNyU4Rso3DYK
MAKxMr5haY6ONDuSyggY7aeO8hlg+Iw73fxyt3VN12pmv8/TaXDYCotzSA/5779H
17kWdpIHJuTjSGqG14t5BlIjeiz2tAxsAmxRFT114oH+Ez4fFEVEUdxSY7KU1EN+
46HQz1T2GF3V8t8f+kNIVkpCBC2byltnYjFEPvhYd8ZQaYcAoileApVQ7VbOcfHK
blCJzJKD26H6k349I9+i9eFnVlmnj19l82VSoPjdbMX5NHY7E6xWuyqKA/qH32nt
fJ+9LxFNnXdawYQHz8EtLg==
`protect END_PROTECTED
