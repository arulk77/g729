`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNaeFglsk/RD0SWJrr854pY49i2jtF1a9uR9qUQ0j5mH
+E4kNaN8NScCLY+7/Oww+0sD8okl/UADorQd3Qm5rEhfQ0XqKl3+G/CcHU0Mh5Lt
ywbOUhPX7CCNwwpWmQ9X92Jy9Y9ZY1Tm8sKpWJvL+6qaJid9/J0lCZ9bN6BWQIRo
iPvTe0A8J7inbk33bKt3XrSx/DARLr9G3Spt3uqIgS/uuupcNyjjeTOa0fligcck
XiOmKsBg6UPp25WIjxJCRw==
`protect END_PROTECTED
