`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SR4nr0nVpKxgeuUQnpNRjbb9a1spos0HtX2R7QQvBlxd
nA3qg7QvyApUb7o6X3H+i/K9BlWeDCwl0G3YZrDZ34AGw1wBlas4hXPdkC2ewmwF
IRiRfJWCMI3hayLmF1ChYy36mK2x5HfXb8uGwMDENKxMeWHcAaHvoD3kPvOEpKEN
GqYe0HJkEi7UC+yckcvME2Ce9ZCZn8Yl3y+zs5cq28JDmOhU0dUKvTDHwHZ2ju2n
95c4EPsw0RT2A9s8OXgcr5ZPqEgdgdP9OiAY+b8vUhZ8Tppnzy++Z6dBXWWVf0AA
FKK0zI9CfEEgo9UZmAQ+twWj8vJLuyG9+owiBP8vZn21PyGfXYb52TKOBAcAcCdt
ZII6eWaI7YrGoZGtiBWDP8YFqM4uBZ8ftnwN11GCUYDOljgO3WcWPOP/f+iQjL2Y
z0qLYwDArrbAlGIMhsVZCszxfyijcM7VbkFfQOjEIN+P/IOA7twT7sLNGk1uCgKH
dlHq8Oof79m3Fyu79uaINLTHdu0P1wmD3ch1dAfrX379BEvfKDrhJxRMGyjmCDTg
nUAjmWQ+b0p9QOHjnMjU2bbbkeg1htwXC6AOwBpqaKxYx2RooH/tTm97iY+7MueV
/TLVTbMJn1Qgs9FxU6r7ltEtkoIym75lfK2mCoNoS+ZOGsX5br4+AJzT3aTXsoeK
Mw+lyyifTUQkbH/Nj94bNTj8PgKSgeftF4rE0Acg8jw2o2OKfzCeqg+PR8+p4sSf
E8v+dsbjkMOxYMah9TDZLF3NvXzcijxsBc0h2Sf64CGkHIDdpVKds/dszvVejDlq
58I+GmizcPJYBUTJQ2hdUMrdctjRHymDnOqbfUp0cPHf6Z+cQJbZ5W3BnqEV+tjw
TSuCYOv6LWZBL0QMLnxsBo/6C+bVuTEvfT83JHSHz5uospeTHiWnwn3bmg5MYjBP
ILDTBITinMdzx3lXIk7E0T+cloQbeMq9amc9kxlsevyPYey/R4eaSz/C4LYTLDBf
PHwKEmQzLV+aHr6dws+qNH1Yjgrjg6DujCPp0RVitAZA8Fv06H6JufSv8QiqA1rI
Io8paALPJ93lXpz/Su0vYE0iZjNL0bfPkS4v5pL05KXOIV/RQnmJUzoQxL/DfsI7
rdBM9YsW+m92a0mXU0FNh39UYBq9MeQIO9AIrw++7qvNVjQe+LgYPyL/ognuf11m
mpKTVA3WFjD9xxdS1rVy0kCt9Nj/MgiDGbKQ76ruu4moaj5vjUGELJ+375aztHFY
T0vkLD3I16l26U95B0Y/k0gajYHj83NdeRTXr+2Tk3ItlDSoq1V59fhvGdkmiTMJ
QHqkv/y5tACelsuEeZ9PWH67wSShlsy2kAq1XlmV0siZ4/A6bSPlJChHZoMSSjr6
U6e/M+HjVCmsq1PDRlogX8JLJ1J7nv6nqSpstmvC4QTA8QOut4uVYp2/5gDdHrZq
UuVGO7d9I/Chqt8fcjDs5gAhMz542ebHeG8+JGcoBfPcAV88fuMBWR24hemWkKLE
v1Rer1tgV43o1eA1Gd5s4041tZNg/PpqjkwXU/5XfxcaVFPntICLVMKt049rlTkJ
`protect END_PROTECTED
