`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOnKgkQGDhna8OQyvAlfZPtu8eOE0vEkLHnD2G2WF3a3
oWVcETped5TIIxVrtRP3cwPjCZegfm7ALYjbPUiKBv6XnYZqI9/cNRje1cVSd5Qh
oSZkD0MeGdAd8D7eg550ksMwtTXmQKI76xVstQ4N4zjwf/Msf+ye4aSg8OWRVU6i
4HpjJYgVPa1w/S/4vr6TxkBidH0hEfqiItGURWcmZlXfPnsxGwgtxjo72s+7EW5b
7PHKqBvR7fBlnenBQhodng==
`protect END_PROTECTED
