`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAPjOyotI8CD97Hr1GQMYNpwzsZgq46J372c7Mf+woBg
ksuzNA/hoQU39XTeowTjb7p54AGAX3BAGO6DqkKo2rr7c+OnYnPmV43PKqwTg6l+
mjlw8Ij3YhTX4+xYfDg9FipYryG2GfF1lGhLRFwOHbaikiSPC6xy8ypq3fw+I0ms
7wUZopDaRTqGgoFDb6dpdmsMM1EFVja13++GAoDdreU5JvOjK2sUYXVzk17iG9/F
Y2TXpGqJLbIxKzjfaM70dUZtXV4RYzGd6yapDKI4W5KM8dz4oh5qSS3Uxa8rCdqR
Md9hcIb8P15QdZrTZ7GxHio3Rv17OLSWxmK60JxkQqrjG3OjoYcuc8iikciXODnz
I7pxaNrj6qmklmAsDjJFuA==
`protect END_PROTECTED
