`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveC4ywCkF6xk1lpdBRkxpCYXbiPf+1S/A7wP3OFDblGI0
d8vNR1DpdN5+MttYrttRImY/FxEXEQX8lB4JUlbaRRsu4QqWcmOYDIXX7eBYa3EF
mWPQKzV5qK8aiu+urIFD3I12TrbVkyDgzApmhJgr5MwCKgrdxdHIdd+0CHWSyANZ
2CyjmxDvwkTS60ztAZCsTsRMmmjKQaue7LeafaE1Fkeu8CyYbLquyqptwBfN+9A7
Uhxf3iBAG2F9/ovcxNkyYcSl6vsA9zl7FTbpxTv4XnRbLtE/292sofT7XwumhpTn
FJB6TotvoT7+7Ohy6/IrdA==
`protect END_PROTECTED
