`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
/eYN3ayVHaBELoSQ2Kh9QnhMXpxo5pCrED6aqJ75MraI/csU06tzrFNYnp2KP0Pf
Iqe6eFRL4kGBo4q5faQ4ytPOFzrO6Ts0Z+Z/O6lhIJhOZH0huBhIQQCm0lj/w3nT
cHyGJz/NzcEK5FfEHu2EJZO/eqE04h/wkhFgK4vBB9Oz9NkatadNczcNqXIOjxQA
4YJsO2V4b6zBW/zN1Mmlm6Eo7BIsFIkOnaX8cfGVi+4kRQPVkr/pn1O4Nz/8WdiF
w5EqSB2UEFQgeutCYSQ9yD01xuQZz6NwKSvgS+NOa0yIu3e2nAB+zk9XO1STUV+r
YUV4jFD3b74Iv4ITxVkt3qWnQNiJh6cT0vc9mSYBuvLqMt0rYy6azR+CGKVHCCCF
mBt8aui58ctFzJQhAiBfH7cX9K3WI8YaAn3n3zBF+MSS7UBjxMTS3aX6v1U1VO05
sWL5F6fRTfso9oe9ZSUzmR4QOXJf7jc2coiLMK3eBzdJwb7tjX8rCu9xaxZcqoAt
dj9YtHmjoru1DMS2FPuAosaYDQZvA07ZRoq/YF/LHSqNkqTB1Q6ub8mYkbYEgj3s
xfnDCzr1Qms8pa+jjvppJ4h4pgQke1hGRXpF8c0BVpsojx25Actsn2+wEJ26Zz8N
l7KEb3xC2CKI57UAY/bmYfXYOnEeepOMtD1ZTgwydZ0gYovS/vTJbxBipx0AJzRG
PWd4k8UpC33UQrCA/S+bLjp3SdQWTYHb1+SoFQ2gHl2BC4vpOjHU1fWGVBDCaJOI
LsDiemcx/Gh5bGHplQMTy9N7ascKkebUsMqHhS64y5nlYhrEyiHNoBLnw/K1FbjZ
g76y2ZrUYPlgRF6JkVbJQ1WcHjRyminFLFt/zE0wvEuhc36iXET3j56CX71IwX5P
dgttSSkC20yNPDLuC9Y1l5hFTkyVXzR+ktsC52gTFiFCmsHfy9P5FxZZaSBVX4gf
XPtgxYV9SrsEEvdXNUHYBFSDLIFUajjJi3Bb1NwhRXLwug1V1d+DQa1k6uoTK881
t7MaJwmVmDHWR2pBCYdor7vwi2rUCo6gQWmB6kEWPqJtyG7R8kKQnuzrrShOUCys
RCAizLeHEcvwVgMcdoqe5StykuSwNJ+aOLeP3KH6mY/YdFaL++w62WCo/d4uhYPw
87U6p8tMptLHQg1iS2Fxu8IwPSu40x/Z6uxj0E4IrKNjDRyrMIW6kiPW4czJiE5b
k9p30EYgkfO6d1Hm2srh8ensnolljsVA3RftvZ87a9BQsKFSXrJnFP+LgRxHd+jX
qZf/iLvv7p+9sU/mbtON+mCbVPjVfCLtucCSxZTIdyieArGGGBvFOrZzQngYpgAe
2u0xUF/ccPbF/T7QQnKCvTgevcx9dkGRaR/IL26WAUYPKZuVvXftfZXyqiWc7bm+
YbCvb638YqRY4ZJ7/jKG9/sTQuQtiHf66NWYOXHaQJprU98wqBJ7EDu1GLkWymbp
LqOuti8Tq+HN55K2k8WVQprRomkiskFNQIYC+N+w4yvm8RVJrY/3Tad8EhCOZVwy
UMB5jpp7am9fgJvPI8MRWxIXdql4EC2zNJt3O2w1zqdAQYZHc1AY20nmta2rRNiF
rJ8+UE09q+JBX3J6riHjsNplKM57uZhEUez4Fpts8FTcrLqcA0EKZPjzbdC6LIsL
2cq00F/+71aP/cLZoYxRDngfruRX1WoWxvi2neeCib9uwJ7Cg/HR0AX0oN5IFRAc
KOfl/usd0WDNAsKBb7M7mAWPbMY4uR/nMalE9gFJyMxk0Ysknew2tjM4GhXZlL+L
wUVhx1geJuwL/a0/fl2TV4jASyuNRi4eccez6CLnYcMAxdX906UnuHTWnMyGDz/v
eYLYjCEJDyThUGGvu3XPdIx8nes+5DPRzqFLmBr6lzjV6JYq3mZ/RJq1gS1W7onW
HNLSBXv0PYUjCKiY8Kc4Ya/iN4Y1sbKJCK3yhZ23lM3BtGj3CE7ElhAcDiPZFRIz
A4rFd2VCwJ7Pai+B43DhmRXkqpAqkmBqSJrKTI8rBF4O4tIlAZ9MJid6KnkiFfES
Pfa6mAQyzS/tyNSO/84AjqrTbZwu1PYzgJ8WDPmQ4tj5liYgJTeVEUjx3E4MhZr8
mQFCNmyf3JPt40iBhVFMEa1fz+onTIRHlEzhAKCguw9H+mWuSbjzb1PR2wlhhwto
lhEJP0VOnW13vrV9m42ujN7OLS/1SHNbMUBozvdxtS3RHfa4ocYkKJjux6nc4R96
f/pLOUEdOkZGNiylcpDlKHB7M0VjnFlVlx9xTgpaUn6lXCEl8DKyL/nvtQgrYr4n
vhKaee9VHjG3Lerolp4qSfcA4VuF6n8I23PvX/yA6lyiBs7eIZVGkNK4gvC1dXsX
E1V/s4lTJSQ3Jt0UxbH7/QrAjPyV7QkTasyPV9ZA+fghI6Jb8P6QrxYGEzn8MLsu
Gm9xnfv/QGLG9bBviz2O0rc+hhfb8CJT0lCrGT9aIIlMyMcdh0BEMZoY5+be3eS0
v5CJwUHSxMXJG7j2iHLU4QAAEFtlbKwtjvkmDtdu88SCg1R72y8r9pLtZULFtikC
n8gJdNe+v5MtV+ggNMPV7gKE6X7hZ0NcwhLUj+/eAfZw2iUM+U1U1kJg4sEPk0XQ
1OF+pAV4I+I2xsMgITEtAbIhBGsRcjAresGxUTVz0czBU2BVaWZFseTIt0+YoWdM
/jVU/fgRLmOjc83l+Q8DbhIPmW3abIeCIzzzcAK2il41DbAxExz84K4JWfOiLjxU
6Jel/H+L5ca4bK7ZzV2XCNE36I6LQeV7P7jaDfQGKXHuJM3f+xY60DbJisjUeGVn
s7mGRwN58g3x4EySWW2Ro0EzoNk9DipHqfQvBtuJWi2A0YcCI2H3Zk8fW1fsgA79
hVHajy3BaFJLi2gGi07aHpxgPjVthMvzebFpOaaHR86Aqsc6mRyZGRtRdzqZq5w0
gYUHzGp99Vwh6Iwkp/NPxXXYVWh7yXY4ISXgudKTtpPBP6tL6A8EGgYbUwXses6R
LcRwOBJDLeLc1gZTxtI6BA==
`protect END_PROTECTED
