`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCC8E4GL+HN/IRlVp9FrXiIHaAjxUis8VPSG4bM745Kw
iHM02fvmHpfRKqdBh7tOzE0OOh7osFwh38pGR8/KqbA/h7/9K/BS15Vg8HiTDvJq
biSiapi+Y48RjAT9wHOE649tTCWY1+TdkUFMxAWgovyKawm5LpQLuSI1ifXOJgVa
sW2HP2eWf0fr67hRcwCmxg==
`protect END_PROTECTED
