`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePdhWDk3Ia818TQtzH4iCJlzkQ3k3+mgPEcELEo6Pxxm
a408jtbEZ+9TheWg6KIF6HwkFBSgneVtpmZB6AzmMFKEHZ3jwWZhbeIzUoqC6s6l
6gPZLqnHAkY3lyj39yemjo9hxQAVqytt8jSABr/kMQeU7EW7FjVQVuQXwJrTuWMh
LyGyrkrwysgmFNE9GN3zsUFm0BNjZy/0cF5U2luNjy5b2PtxpxckWfsuYsHvWCP2
s726OCPic2e8nd/zNVVUF0rVnh4y1fSIIEWeKlnPDz5L+vMDGnN7vM6Se39KLb4W
8GrdOf3gdv89EWkAaBND5ZPMaYu9Nu5TZckHnZa7gttqrpETCvoho+Rhpexl0D6L
IySNH6X+jK7MGcX7ecffefEqzgO4j2iFj8wHf/Yn82S2wF2i27vwq7KHYsbiXc6S
`protect END_PROTECTED
