`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3ON6twM0bRyFDJLDX3Tyer8fsNKdRAeCA82M9Jn7LrsvWPKUeManybWOL8WrjJs5
CrHYuDhQriV3urpGan8VXnU/CFX7eGuh8Gn2DzmSb/iOrSvtIaEqAqDFWHxFZJ0y
M98Q7MAIZEoeM4qB0b+zxXT5ASLiceFOhMT4mrsQ3xEMIZ6doFQJZlev/iXYvMrH
ZkLVnuid85IFWctokDGWkg==
`protect END_PROTECTED
