`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGpcLrj677yAxkbHMiqeq35/s5P7CdLoO6kqK7UEt26u
VPM/O2+0pFwhxWt9/dCEN0GxY/A2ILAIfe3N+3InHxeG3pZiD50EzzXuyjqpcrcY
v5nsGWLb6CP24OlI+gN87hrW6dOKiKnZWxMgEmEuBgso7GDK6K2E9gDXGE6plbso
Kj1F0nVr52Myq9W0RCTjyFUHaM06RVSmVx+hrVPW4gRVA90TJmGIBYz/G7LF9FHp
u5r62LQGL0qtUqkyy6gbyaZEzBhtTpsED6wxk0l6EONuh+iDRSMHzkLgq2TKmxkY
PqSptaWvmC1s0Xsg+VUZWKjcw94mO7J5fzBSHECNTVDzXW/scGTySV6oc54eYRXr
TQdY1uQPZem/quQGIf5b0JcSJhWDBJTe/OiWZeBUMa1eUGFupqr4iP0/Kkqyo4Zt
`protect END_PROTECTED
