`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDATiu6lfJ4iAqVZNsC/G5SmymAu7jL7BEYI7w2KbH+LdH
IrcJLrmgDtqQ6F64cZTEUu5x+gChHhvM61o8h3ucdE+enz/rEOSs9Ua4VPcpi6OF
fgNhT7jx/cVxTwt+P8GOVKgqK3Y6oKj0JeM4Ewbm8rY2RJ/C/rBm9mq1JNEsv6fl
oZsR4qVyhDcdI6DV6wiKgwEqNOwlAkqwMJ0PvBHX6x1BqkxsayBUyUMmXyFHwnhJ
JQ3YYuEsHHOEqVh/vibPkkjnMmVqHI/bEiVFl5y2FxYVkGTTZ3wPnHNNm650Wesv
zsqkD4vPJqvomUgCpF6rIegZ1rBIfRpLiekkTAu25QOdaAiswi8BTlWiqBSy0zv+
E8jXblZv+ZCOWah5wPKv+8n3VfWE8Pufbiuu7wQu0IkyfLDpTV5Jc5hTjUJGYvXj
M3k/VAQyJ/1YL9shQE7w//rmSICV4GTwyKTGKkz7nyEk/ZCYp/eUFRrxYy11bXn7
Wa+41cnndPlOEcyZxsOu9aN1+15hnBQDobh8E2jYjcHYiqqeP8MaCTUr/hthagAW
RFm23a41cQcaXrAkrZUaMTg1KcX1ch/AXcoppmvQh9wMs6cSbst1OuDlmiDOWeta
PW0L6FzgdtfeerXBjBwfR73VEyKXysnWXWmihDvVS+6nxXK4XpoUkxOw84AUYvrf
F7ggsrWn9kcI0O7zBbVktmGuv7p7Oe27PB9Nbn+DMdUcTC4B6odKzssDuTMQd2sN
jdtRQFGtOvKoTyO87XsAut4aEpBDvDCKLN1dMtQCL9PmNebEDsCNrkXxhIxAoWSj
aeQnjrOwip5GcK9xqNccjDX7CORaod73PZ2cAQr0jO20JFQQAonBKiJufS551mv5
`protect END_PROTECTED
