`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
5FEZCWPUqFgG4fF8vxvrvV0mI2WRXGof34q2b3x5EzFYetjJzx+0I6omVdMRYWIi
DoFOYktKIRIDtV9MuIfCfyw9VchDggIjUZSU4SVt0QoB/wLcYJUbgvwmHQpihK6f
n/+2MjbOkVnxjwMyH4Zv3AwmjyuhOtgS10ghvlRVBx7ij5bMWwXnPeejvOVcIXfX
Rgl08tGsB2+Eb/LLpPyw5hoA01yS8ishVvwTWvSvcILGJS0Qw/rUiY6RjwX8zmYs
254y5v5CwtmPQM8WTqpPacU+JCXTfuuJxhzuoO/sRJ6s7CIkvEUWgr52iiIEQFCD
RLy3z5Dt74oVadZgCEc25PrCvXJ9OSTM8WyWTyE9x05+VkXtpZTDrsj1a1NYQtqw
AjEFur14G6yC5gz3YlIAqfNIEvGgCrtIU0Jq/y9YYhQ=
`protect END_PROTECTED
