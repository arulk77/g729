`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
LrymQcokOQf1jAtJ1xL/etuAIvO5I4Ec5vr0chvjb/i1xpGF6+qgBmJR59vB5GBN
wvUMT30GOsO0QQwrNBeE7qjJrIR4+2yQKWHAfWiT6llgJ2Wn8DR71yhQRCcwzC6t
IGSqnhCapuqNP679ChFg+RfjLfMMikckUJ5S5TdS6+XuzICXmnl2gfrYybMGat8M
zHMKjMK0gzIv/5QjOAg1QTOZXVvlZf9Mp2gXZisgg2hkbmvIpf+2TTnjVhwQs/EZ
sjrVuWMq7i13T6vjkJCnBsfX6knSZivW2UlkS5gNUHq5j30WfrzMI63mzxut1w1y
HNLyHing7znTf/H8vvkr6r8MqYx71ILKGG10dAASF24=
`protect END_PROTECTED
