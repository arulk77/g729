`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMMXhiZ8AODhBMwtOwL81RRMhhefQz9E/tTTKjLv06DQ
z3AZ8la9mnG+k1lVQa0zBvATxDcOj8A2nuEaqKsBBvy+3nGyvSRVOvP72/8UHdDH
2xrRx3BE0ymG+O/A70OYzajoCm29/XYVa2YDRDu1FNOoM5bBpkNlkG3iieoWjLNZ
QWBO3DAoc7NgDoqCpVXBB5aPW10MBLdrrlSVKUKZNAvgvkTT13eDwWWHpM2mWAzX
S4HhRSHR6SJYzAO4RBW5dfM0jn6bMxXi1SUlv7X90F5/Ja++5Cj+7COA1v1Z3s17
TGmZa2DEh5qRQ5t8cKgrQM307gXJq/AkY0Hzes/7epVq2eyBbPJ7SUS6yA0GO1nf
6SHsGwgCz6hTNvTH62R4z/wjSN5Eg6cN5dVtlVAkO8sqGmG82CNix5jGub3ZYPN0
8e5ZraGom1i53ONTrH/bx0gMQ4tkAzu7gb/PuXMTrR/I/NaOytFa9A0SQcY8J0iv
bmhjBidXHHtSqwWCohBccQA2enTrhH0ZbR5pHMh7ieWLw9J+3+xdkYsk6QL/Nn8i
qsTEyzcqQNfBNSLBCkkS/A==
`protect END_PROTECTED
