`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aSzaByWvdCbzr8lAEqi28PW06NYBYUyIJXXxhLCQH6lC
V291dihPyRwTmfSz+302YGla8bViVi3HD8PSAuxxbfCnk65G/3qxotX2Ljo3Utck
y90U1hVvrzrL4KSVxE5JDt6eYeO4gYAa2ZsjB2WVjfkMACPtKcYKskY1rXKV/T+8
EApeORdkkSqHNOtFzIStDLusxQKCSwXnT/ldSe4fkHFOlmA1MdAPTQYT2luFmD2v
3kJzK7I/h0bnMOxOJ/7JoG3ZO+5NUMRdrzaIH2MGL51fBw96vVTqdyE/es114ulk
`protect END_PROTECTED
