`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePkb7W9G3bHuWIOWxyvCIQDomGyLX7tDHRBuPk4aKfek
z5UBhq/Dm7oVvvXiYUbqxyK892dw7gNXp/PLJ9QLe9TBAIfETnzTNHlqcjKxm+XF
dY4ywVcXSSHCygneMsj9WWtpBrdCYFQBpcOPMaUXUYzZM6CGy+Qu6U3VP9eawjVC
HYW7ZTg5Kcafw864NS+ll6/awvr1/G4exRNgf63OOxhKTV2tmw4CjwO+2nlgxhIK
Q/x43IN18cJC8rc2SIBj/hnXwSqdCes7Ow9oM57ngQ3KGfDqlP1KfMEgmLDvkxNW
wwfsO8urrgitZ3rd4/X6p4N8X1Fh+/6wjj9n/PRw+f9yEyzUdSIzahzcDx9HRCIc
TXWVpOtFj3qtWyE1BgVdU65hu50gIoB59EzUHlKbd51myvqNFjhZPXjSqw51RGhY
15h786E0oxqlEbbrfNCF8tXP7rr8f++xse1S8JyA+xaOl+qNacSB3yDt/mot0v2u
QNlW9w/wHKDSL43xcjO/gkJfSZuA00xFAOBs/GHahO5wvqXw/d14nJPWeU76roHe
QldFD4lIa+PAf5E6oB3DpodBwKqIpIPxiXHXr3NCFavA5GTonhJtRSPgleAwuX6+
7bNupyMsF+FthnzWsy29FiH0yKvOwwoxVZmJjqDCQT1LgSqhj0r5VAOHSPv7U63e
NfAIoLCL5C4/cQh/Kzt3kB8U4zolc3Z+ufPcFPr31P7wINRotMuj1vTtjhEPyEw6
uNykAtOjGe4NnvIUw+onbSmwsym7L4wxpPdu9VrxrSCB9XyA3k+v5gBdOL+rjJmh
pXRzGpTBiKxu1cQm8yco2bRvHRHAJ2YEq3xhOVvEJjYa+umEgtP/nytzmH8hSIFM
QpTJ6Uy3h5f3rpebQmfo5vIPSBb62pLJHtinYYrlcW1sjnS9X35r6ew20828IAKB
ia9Iione/l7V3/4+Rfk3iWyeYV4r2smiPt506HpVCbonTEDhJMnuMmdxnlo+ktJw
ouKs/AZhubyyLcKZHTCJQ4dczSceQnLS2BhXEyMiBbW//jKUbFdJgshp670V6j4H
5yV46zhgVPpWufqecly6oj8DLwD+3I9fd/hrTaOEVpGjPj+knsS5BCwwBhXnFMmC
qssuU+sudAdPo497hGu8mSAMPETpq6RuQq1UrnMozvd023GhAwgQb7BT5qwmZWq6
E/iG6pBs+/drb+ZwC5lBt2wtT0KCjNUTxqj0cf1u4Z8NEDvqqgUEWtcl+kD8hpYW
eafEUfwyHbkkj76NhpPjBfJRuD/1fYiINiL9n7YTjv/COl/NQhUTbVfYehL+9GDt
x8mrpKA3b9BBS6Xs62eSPjqqZjYYfcZiRz3PXYpcdLB/vDYpssoDUIaQ2Ik6LUf6
i5eOEc/O9gkQHHc15aUDwJuFka+j7e49zID1gYhv+0K4LV3lghEk6jK08NyczjmA
IXq5eWuei+NrUx3o1tQnK3XoeiaNnMF45WSMQ7MSUQZ/gYWvv5EUt3Fc5fIcilzg
dCAWLeBFVUu4+TWaqvBryP6QzBF2dR7vibspEGaZaSWKr4yVABllOk37EfS2EDIg
bp1ee8Kg7v1OLVUxSz+n+ME9K3Pb0Z1dRvyJUUEiwLVgYINqnEq0vMf3d5Bz0KSg
aiMeOLFLqMbk7ntUomJsrkhF5pyWoPGM4fLSo5fxuSzFaKiOHotus1amioE7CntU
p2DRhFiqLv6MWjkakKfXc9r93Q7ODZ26yhDdIKlQjFrugWwp2RUryWxMMx8huMCF
2nducezuAX06oSer3xFARVgBc3uMskQbrfR0x5FurL53PFg8SRM3ClQZqgNxUJ6q
/9nolgK1xpwdsMr0BhILSm7N0D7xMgdnWSFkOovvL8ZXYxDQtW97oaTpmkNh93G+
nwLVngX/T/zCLs+AiBMLv13A327dc/aHYGX0DYkmFiO95DZpX+z52SEeDyfo1bA7
r4OfqJynh2cSJBo1BrqZnaAo1fqSh1f3FT2GMdP/gHsF3jpe4IHDIFH6jdUBKC6Z
QIuYiXJnKalMqd3Vh226PdY3Dw6FzLdOTV/hIn0jxeySdBMW9h7f6BODVE2IHuVu
joTxGyZ8BYm7xOXodz8chBFJVkYFX5P8ydEJ9QHI/bK59Gt9EdJbWv6F8BoHFQjn
zUFGSsqwtfAmZVeYXU2l/JGD1sIp7FN3mi/s6+8U54SOOgVJEbsiKEmy7YbaQaDQ
pVEQzl07HcIYZLQ2dkP1vgkmU3eE3ht3oCba8lKJvp9iKdMzk0VLZT+Mg5CtLTQ+
UUXWodClmTMrS4CTrDxPPklb5vXbfEdyZTwVogZPCOK82BgYW2eU2gci6kQW8LCz
ocTltxS63Uk/w5MfLJmcNHdGNClif1lnX1BjY/PC4hwfaz0A3Du1Ov/nAKX+xTaC
nMfG138pPUlsKYeUy6XrtErtXlK2YmSzlpf1Mfk2KsE3AP7zGisleXiby2MQTyxO
J98RnQ14uK219dzlTO8UrhTht5Ch0jgDXpuqSvG4I4k24pC3UA3wxJ7tw+yBpaHs
6lPfNHL4I77+soyQymFjDzWtYzVlZ0NnS6QxxqGFL6wZ4FSQYjX+pb9hU1i5B6wg
mhC/sZGb68NaifGNumfTDBQOXAUHlR2IlrqYQWv420jWSOg2j50qw7TrwyjLPhXr
2t4ExNSxkG978WzbbgYMnOoXrjJXLzAbkcVz3FWZ8z/mSxm8XzZJ56IHM2ncPhEQ
1QFGY8lS3DMF7I9ADtLzVht3IZHUBSPFgulOO+zSQbpFhxmm8xJvru89/ZsreRVa
4hSrkeJu6ysYr/iG0uu1rkA59vp5/INvoN40+VkNRJobAMJEXwUmPh/vbfKVsdro
C+dPKSKGbTGXmVOpDGoWiOgac91e5+RwjR4nh+td83bbTJlxu4g/wU3JG/WqfuQ2
AqnSU2dPXe3DBsi8WVQeOft3GR7ue4ojN0iMXgMG2WNR8ahbYZqxmJ2k6d18M8bK
Q703qC1a/6B0xO01zFK5mHtGSA9zsODpfMdpCKfc6hc9rDjn7tMZYBXP2aPoZV5u
02PhJ28i4fF4K1e3naqMPeWguWWZpHM+yPzuFfYhHI5QDgdIpVNITg34uZGAabSc
R2P0whPVas5vPIqWwmn8f+IjNmoKWf2aGExYUAXLaIEL82rrFDcCqY+6vIhsscCx
T2LJn34jn03e46lM0h9spQMSZkj81HOUVupFtfXbfQFhknE3D7aUTfkmcuPK/9qr
bgB/YzxtyFtX4QfQvDNUcNS8YsxKFSMQ/WS+QbhM7ucfSFeizUbAWolVSHI0vQTo
OrHU/EEqM3X2xZnTYAQUSJoLAyYTfhZ0HkwhbCRufjQAeaq5AnApQiIVygSsM2WV
H3DPhhx02PEpu3bTOmew3trRsKL25J67MO2ifvxr6VRUZzmn0Bpvm7UcBu4eSTdr
OadRWDe6If9ZUMun7S7aj5YW46OvoIeNSTGXkdFZhHozfroEcuggP4E2k4pqA6Vh
uBtYq26/7qY4BymMS3ywbcjYiWeXsnj+q8wyn9MqgQoSWKB2mp477w7D0BhxHfNr
vGi9pBE272njKbLatlZptBfLxerBEoRq7Vb4RD81BauRS2PUOo494cPqRSzOlpuD
6JrCFJ1urz+0TMyzkkCkBMS3hPjOIa90DNVlwXiBzDRhALUyQ2d+FyqsxudhQi8N
GOuN54QLn+5Bz9dVIxTvkjSFlsoSaqLnDqEoDlXbw1kufPB7zAmeBY9mfG3Q/IqX
p9cO/nP2i9xfn7Qz6Fzs51GYJHllmWEDc9iQHLPG5dySyrrAyHSE4yrkAjgFJnYb
0oYWTZ6594fYZSw0K2m+zrAinm1bQ9O984cOtc9NulUfR3x/5OEj8Ke9dzqip526
mssmbTT2/l/+KlfQACHJll9WpAmcH/Wa8a0KBFeVn4v84RZx7eYBBiyfGYlZlXES
3apmRGeGWy8B7yRCYIwhjVwsee+ze0HBTDo8p+dvgP17cKI0E8eeTciPE+60bXHq
+Jtp5gcG0YxqVC3GgNn8+Ix2qR/593r/r11C2SWJ5BD2gOfM262bhU4Z1fFjTGFB
aXfSe1cJeRr2md/ws1ebTguG7RM2t9aQE7P27AInx9DsfW38wFV/pxM1R4hm1XuE
8s/5INn+YxR0ClPjU4WfMuTuz96WuC5dXxwU60S4mclNjXdADGBtUovXgTb3jbFy
0JBEvN4ABCDUi7K2x7F5Uifh4xohC3N10AOqvusqGs1C4TC5lxROA2bgaxkb6JrG
CpbRfY4hlvZe/HlINg+aPpAfwPbgPby2kJ3HLzCwm3dLT9BiwIc0VTgYxg2ynu87
uGCbvAplKeBeZ3srKxuKgG3QDuSb5z3hI/mco9Go24vymT4kFfnr7YgpyyvQeEYR
S/oT26eyTtLEZTFb5eZuk7tWpIR0QIj4RXhtt+ZRwnKaWXmc5MpMuzk2TWJmQuWz
Aa/MBjsnDJhYy8MxorRP8L7pPzzLx9r1CtAKgLeHItbPw5j1NGvf2fIgxQPs3I4P
ka2NCw2TLpbPHSK1JSwdray6HMmBHed4Qk2NZa3bqyBpaiNSD/VmJj0MjLtIlPZe
FMUFFwwpI3Dzf/UhV32LdsX7VhJeWqd30aVH1JVdYn4q6aSOzvwEKdM0Htc2+Ca0
u4h+3P6bFr1mPbRPCEv5Dzrk7hKGaE+sqF7YhmeAwXBQ/IBz3Ux9PKKlbnV0op08
pSl1OoBJK7VBPWLisZ8IxVyA7MVW42g0XB5qAC3OLHr0TpYv7TWZI5lxm2Srpiu0
NMZrB1RAIUE7YP6knlps7b9rnRtK2vrC4oqoe5K+EiiuUdMp05Y5NiYpO8Ax3+Dj
RG/cdwqaGLm0z+Sfi81ZFQWpePXl0EWjmxYwEwuFpQSrrPqAT6Mg/xbHf7wWKSfY
l4PHoWYGo9XXGxEJVposle9wdYYLWyh3wWO+FyTdw6lt+MXDsL/kYpkRp4JSK151
7fXoNi/BbxHpOAX91iWzOvgtUojVCyXv6ET/97r6O3eZLBv7EpfV6sA2ql4t5st1
RUodzATNpuuX+7gw9N0/wwtCQ2vB1of5rbjh4U+8KeX/xtwoP0u2L8g1ggvlKIh+
cRORLy7lAr2qz45A6uWQw4UOEsiVM/7mNTHEwNJVOz9nui/YmWjds8BSUUNzBB/G
0u0G1LetLilZf0kZX8nMDPl8SZZ8I5DpL83Jc5JH2OL5Ge/VCEtzjiBZ6bvJCzpG
6VLsmLAryqI70GSb/UmeU51+9RbKCimj9yoMIrZdI1Pqv16lQEUBhqiYJG4ZkcD+
KYa3Q1SNV0PiKkRap003hb5kvEXXChv48odG6DQtXBUssorf63AT6NqzbQdIPVfu
pZTm5qwQHchs28KnKJCWBlHNvz2gkbQqUyPz7plBKJe1PeExM6I/7N8naPjBirGo
Zs12VMZxfcC1DmOVVbpqo6TYl6lBF5NlWL3uUnWhJ39K/O86bKC3DbiEcd1LAppJ
W9PqYm+edp86RmErTqsiwBMzkyPXKj0+DL6mI7UCLsfUtf5K7Q+vNx4aiwnuixP5
mo/P2uv//+B9dxGv2fZNrIbatnCWQlOwW8ObRy9+FEfvxlIYqeCzmpo1iQ5tUSgk
aYRPxRn0Q5e3m2388mBO5R9iOH2VrWM5ZUNgAZ2J9/cimTppHK2spSLD5hqwghE6
TVo5U20wucS9WaLr36r6ZVSya1XfhoUyz5CKHte2p6CAJSdi0JKBIHlyXMASS/gp
QjldeYjA4iOkPlQVt6W3/snEX3GTnkqJOZaW2AUnnL+W1MgYzl6sa/T+lMBLGKOF
kK7QD8ufO4RI6iyLgqjvyP59XsgT3pUAOalL+GPvZjODfC4z3+H92VZn9lgZ4z5k
k6jT2hIqbHcIrLaxZm1bLdxFEgiKQuduk1v2KeUnBwZoHNtLC0G3sFgBvpeL7X3D
/E/WLC0QZMmWvbQI4TOSNQuPzKRm1csWolSl/BhrfCHBGM+dJZyOvqhB6OTsRxT7
RVatg6mZ36iRZpgxLMLzhiDiRek0IK9bYzU4cwzPFGE4zu8qlOEOHeWdxfmXF5Sc
Q/yCOqPmnHXaI+eV/GDMy8z0EsQ13FEBJHxYiubTTVlKFXLdd3w99vLamZLOYQ9c
hyfgkIeL0fNJ7Tbz2lS/cjwVuwyFDjIVH0isFKYWfAm2cUdNBE+b7flDBKQ7GZFI
m62eXNhUNu6BQ5afTF89Dnbr4JZ2TkQRkJsk0KfoLDZhbtO3pnoT7TjZl6fxmB3U
CkhasHC4WD5SjGHxBGOuLsSjH+IoL4RkMbuusyxXNFQ8H1wKht0uT7If1mxB9Z52
Pcz3KKWx5DVTTj8AbN6fDJr9tLnQmziCDDn4uMrIYzgsMdzjXOJugsSLjI8k3drL
6+7t96TL8LEoFGRkhk6O6toBkpHdbOV74nLIsTtT+dGxMjsSBoRF+FhYvnX+fKzX
Rb2sCoHWgREmtzjURODeNuOQwfLGndi2bSsIIHWMeYyRzmyt5uRvSYiZMJpklYqC
9JXQoDlEhpGOzQXmf/2GeRO1h7LhBy4hDce2Qob/g704iQCgp+7ldvye3Ab7vT6o
aiU9mPW4rUJD28TS1sGiMGqGRm2zKTHAExHRj877bEL4svOfVjx8d4Qb66edNSMl
dmndhgH059bJN6/CYQIS9uY/CE1KUMuFehA99In4IxIQbUt2A7SJJlgsIk4xvJBu
IaHqz2Fc6dXLrMIBcxPmSR1fbhxTlENKwHdbchpbmNuah8kJ6Falv5Xo0ytov0hv
Bsy0YUOFSv+wayU+R19HbUw/MAsFAjqcdcdf0sx9Buxp1x2lHj69pHLYm13Yh+Ww
XY5fu8mQZsBfO9CpJAszHtLYE1gzgYk+3Eqy2rhn4fE0GHpERZhDlsEWIOxwCDNy
DcsGoHjlz4bJEyP/qdAVpjdA5t5INqf+8tm0RS2uxgRIHBhk1d3MMmHNPr1ANkl8
r2+Ix8XoMPVYZeMX+MSbNRdObd2aDatoM8yuhpN4KBl3Oy8KpQJ5/SUTI6unEtlR
+jAw8Fr24l3V4bz1xzxdqhsvH6O3mO931XBgkRHcui21KoJ1UGz76aRWQB/wLNUj
XiCtwtbHmGpFDvSuOc/1qXngyx5eUrQXN82F+e6St2q7UCz8SeTk7bp/Rj7EkuAz
qrBsgQCdf1rmfhPJf0fwh9/1bxe5mjbVDkwPjnMLYcmoDymW9AkQihD+lgUjHYZ6
c+vgG5WBsEb5k69R9gDXuwC8hWxLZSedmSPFeYFsOfk18SUOn4K48vtnabtnqvu2
jgFaIQn64Xtw9shz0opCv7KBEL6CbOzNi2an22wJhFGcr15bZLqzDXGcvrl0+YUt
2Kj+W9PSEk2UQAHLWn6rgxcbb1tQtbVD5Jp5Y2CBHdbzbuEo0et1gC+BrPM2jWtN
HqykNCKpaquEEXq+ucAm+4omVSOlkIhDJEcfwIm8yob6gDUldtMDz1vHavyJiZ/H
CeLfdeHUyr6O3iai4Uv2jhWcI+yR/NZBEEV/ZrMGb0w+9dYvZtzYkEUq3I2l435T
Js4gSFlwIVEQVHappRxgqS8ACcAzAoBN+YbIl3/qyXoD/OKO4q2kwFvYXkbdjsoE
rGuAj8uRdtje2tsiL7UKxG5UyshQQ1r0l63ZHU/w5ptyxMOgDRQM8O6KuKXaTosF
lR9vQGK7W1qgOBit6V+zdm5xyBP3ILX6T8niTftErC8tBNYfZQiwr5mnPA0jgGtc
sJTlzF2+aTptATzcb36yPIFjYoDh5/o2vMIiVpbv7yD1wPkhfyzLdAd4E0Ih/oie
WkZ4L0X/lN0gX1M2RWZXSFVRJmjEsfr05NQ5/LAtdJ/A9aFPw1ARBu8c2su5kyiK
PC6mV+C9CDQTjZcu8k/TW0yPTGpCERnVy5i4Eu4K9EUUBqJuOIn99jqMDc9RBlLI
ROuzyGkGm1jbOUxfkD62SEaYBdJeRyaeZBRLG0coQgG35PAQOBXFGqabwYu0tY+C
H6apeIMbRe85zXFnYcnLM1ZJSitt2PSmTPk8IYRyGuWBK6GG1UGmtLrhMpzceDjL
lwE6Xu/kx4Jw4FoLEhewsoVmoybrInzTWJOjy9TZ+18sRX03tYqJqBWC785Mp4zN
SZCqIKoZ/SPvphJyfMljpfczHyc+iMLz6JdNOmzS1EoEgwD8TO9N7FJb3gYrhnDO
qiCbXODmqtEoJz+TQWW+9CvyD200XZJGxKyO67WZ+3KtqNYlCijjCGjmw9wozoEY
IOf8RzoTHGYYozbRz5shgrTrXGgMYQevlJwq0XkO5XFcHMZx6eGW8FufudNgq9T3
vSk2qHdV/LR4dIrIMV48rmbEJoNtiGxWLNTC06tQuIpmKlhMRk3Rsj7itKVoZKYM
H6+FlsQVL4kSn9RiqsMWHI6of4K8Uhj7RURlmMCHeG10x8vQfg3oBQZ1xUJWk2Ze
yxAJmKnM1RU2YJ0PdGwKD+gHvqzzuy3+kw0JLNQhC0yYRrg358InOpAZtDwfomlS
YZYmtGKytaWhzG5YB1QBGMp9FfGIQpol7ysEYeAkqMDffsM6PKozdGngFaAl9PgW
HXE4jKMhcNlO6K235bQ69HtTLdvLKq/DmuKoidWfpsBs310ZAGY8K7gtOGhrmpDx
6sMUv8wRBCtqTIPCljKjXimZf8mou83GsPcDpHk0cGBW7oUJ1cA7Um0+5nGvyF9x
+LKEW9ZV9FGkoWdsXULKISamhIU0rOTFsk+loWIA6fnJHfbAIivWhSRSNMrCFmgu
OXCLOOwMZdQpB8D16zkxeI7r8OLKR7jU5RKmJ84+Y3IdvBh8oI2vPtwApwbLBqFA
2fkazoDEZjTokBLIkYKyWfVZGOcTSSVf9b1V1NbNjj5kDQMnp6xNY3NgwoRCn6Wb
Y5A4JP8tRRYW5GckJ9/6AjdZZiMUB/Kf9B3fZKnU2pnCZPKcLCNLvb+jB1CqNXcL
stqSE03DHAru+7pjVKEAhtelHBOGLUraeAsaMMLAC/yRxcMkl4xiudfs9euYoqpT
BUFmdishInbQvrv3xMa77R3/A6G7y7RFn6T1T3PCR/K5E7JsTm5H+s9rQA1T2ty0
rf4bpj+wFd+ws0Ot8NKN8f/+adTpcv/CUmgnV58gjx/Q2wLCu9YJA0GaUPzDeMD9
/7XYDJwf3s6cPq/6f1V8mrO53p4p7mlb4M1697ErLfXXd+dETyTUZokdw9tqzQwf
kkf8ZZsA8F92J0+5nnwzHKnLmZZVcKz543Ju5sNdmlE02rVPJ36d3igOwEIXnKVP
tCp9mRGt/brM0uJtuCsjZRailHcieGYuOP8Fo7fpkjXoPF9V/iBfKGGax9Y9sPt2
2BuuEyfFhqxIzVJONAkB/tdnQBfFlPgNTN7haRLzQiQQbpBi4u+3u+0pCrsri+s2
QCB/wZuGZsWuShKNY18CubUo42fKTs/mWtAILZqwRuf+XYtcLnSOnAFxcXB5n3W4
zCV86QULRtIlHeRFguMZMk1GjxPgX8lHhl4ctQ8cXf2ZBkHY5uGwkCjFOiu/+1T7
8DEFGeXjrGhtyykgmmcOWloEqQ0Rzlr/tWxVtsqOfesy+tVzDP5HGPkM1HCCzbiQ
YWP2qnUdMF00Zwzx7cJZwZdzeg0kXZviLhPZsg18IyUycAjotvvbrkY/mIMYEk53
2scP61rV7EdYR0fhWPmWYzdov821fvZqH16z4gavpz53pObMhdVQSAftvp6Ti7lx
sywI2Z71jFVxxZQpvh3z6LY0qkCHf8f8byMylZAqUqyKmoneZWNajgL2Pyf2KEUm
6N+ZVCWsPwhV/SK9EDh+0glYsyOaihkHW/ugqsvCdXIM9AkmhjngwYP5IhPRnI6t
9Um0xjQCSprGvB+Pzg339l1HPv4Eaxxi6HeaqJE75vpraKDCjBgfClkh+mr5c++9
qIiQEMWJbqCYOKtEGRh7pmn/g7GPvsYiPWxKMkMuRyvxHZhYh4aHi3o2EXVYnklw
Ro5d5P76GhD2tle1JUUyEdRetP4jAeUZ9lx7ujceLFtrESp9AaFfCzlhfjwFmgoc
MfxK1+qtV39havovB0aeljyBQ+wullFfBZEYfu8+y5jcpBLymr3ejKdSlKRGpw+m
wI0xnT5S4Ytb4eNZTYkh4Ut1ZeSFBw8BHYIHBIvvvpGB7+eD4DH1b0FRv2Q4gUBR
BrL1z8l/u7kZge4dJewFLNLX1aseW+1z8hPjSS80ymwFRKJXGjjK5wY28pmjVPqY
eyOIKfbi95GupKpxKIaBs+ZsbcTfl2H9aMB733RarD18PgWTxZMabwKT4sYnVsBY
3Q7xlP+QviMpSQsjqXr5Tld/awWoqpCD4StMzXqW6v17ZOFOA6lGQWwIk3qhOTrO
6o10jkMlO9nTOJwNURIZr6X0jOrKXuJe3s6Y9A5mV0jaIebqna49RLrmYVRU++C1
LcMIM1QZa0/toUiDn0669mHCE0KDKQm5GKJQunocLHOUVrP20ifXqu2YxdYmNmEK
dxzHP6/xjO/RMnhYPcPnoYtuzicMuMC1UQSfAUsQJ+TSLwGonafAEB9N7vSYDz3u
aoTgr1E3KOYwZ5zI6p6D+CnIwi2FE3WOceIGEHbU7AZ8Zcp4TvIs7jE5upVwoYb9
Z/GOAM6ZqmNz5btUfqVs7MkODQNJHErsrwk+kundFTmLno8B52a3T109Dm7LtrGE
ZpP52xFwcN7V0LC/E0Dyuh8FQiyeLmhiKNb7TV+vvcBTHa8C+L4PZYckeROnDxss
q49xQmSsLlGMuxzgBGH3rXclo4USaxBZVlwTY0kVRbMlQfgZ8RWLJGdaMlPkJWbW
MQo5AGL4mLy29ymQdPgea7B6LWum4YOpGHtc3k8N6u6tFc2pWbP1OwDyLjk2Ejgc
lhmMX0HpY3lG/jlU5SW3S0O5P15oLw8XS8YwAavJVkRA3CqSKAvJU7Vz57KgxZLa
/5tEqc9ynFHNWdzweERhs5iVTHws5cnjg1NLKBUwQfy2VHcjjeCuMTZEECS775+6
tPRsRGMuAZirGGIK2dVZGNxNY8E7jEd1DdlzttaEsYsc4fehCQ3rgU0KYM4lJr03
kRAeSEM6hpWkjC3nwojSZpR3IzQKWOBALSkhVFWzAHVBXh7k419AlWSjWfVmC7we
fH6w8podmwsFhibEDOkiQKYVCN9bnUFl5wCvjZdZTQypUULYlYKO2ZoJl5Erkgv5
ZpsmeGWG68JZIV4tHQ22jK3wKV4UgsuNQXUWfNCzOwIuqP/P4wV/pFA7A/kKTBD/
sN9gazDhIccwxPTZdfAsV/KJEI4N8FREsh8riXyk0wyIWTuWktnqZXgwFcJ1oYx8
ceduwH+RkL5QRPe3KiZDah/dbADTRUqyC9+ZlheZzf8lNauPsHy/Gu/Sn58DfyJL
yROG11JA2lCiCu5/wXWsOcV3L0GjldLB0IY2j7GiCn0WOG6VjnTG22n/gi/GJ73l
jLEVql40FmrTsNFTk3Y27XmPDywIBvhu8KOZey4uHSyUqZuUSVbi6/KSvPSGMJ5Q
TI9iiJNs/7oizpokt672Dfzk1VzFdRILoKMIF4YJfSmk5a5BToz5ThT4NyTY36Na
FWpAiLaR560hp/qkd/jtryNE4DzA7s6RvB1/9D1VAGkqrtcnaJKOfu99/IsmDZR+
SoBtftgE/pPrm0Ctf9AO4wL/x5sRO/qihI9HddTl4nzg6/Jt8zfjefskZqwC1Ja7
moCQfm86+xpZkNRyewjhl0X0p3ggKi/tl0u0S7wLvmEnjVOPGnBYsIGglq+GyDEq
GIjDODQWE1SuMaIUsszm3yY2xHLudr9EMWC6aEuUWlNhzvMjhOp4PLj+kky9Mhz1
9b7cOq5yOjUnesx42xPpiltxJKvoQxW1EOLLRTXhq+W3tfwGjp/bbh9bqAVF4MO1
OW9k8HaR/4pKdhSDv8Fn+l0TeFkEt53YL4Ayez/JsciwAipGJJU7FFZxdIuew2+4
EJ5bO3tIT4D58+meDG01mIqsRKZe+FKmuPSKqD3qRCWeik6oHySgirAOOPUvor4/
YMzoEJ3GwqYlzxdr0cHw8U8uhWmlBBU3JTFbxPv+EGwGC2B1rlYO1FvqfkUH2N63
vy+eXw5QgXMfXbGXVgJhTIOYYRpwWCHisxt2/LjxPT1GMrHM6WE3Bo+7UawQx8PY
gLUhSONAV1xq/MCTpqB9Vd8NJyz/JNnkYeuMXQnpxYE5bz/0658s1/hCXFlE4fxs
g+s9e3vF3B12IANjfL85R22XKeNQOtmHQ692WVHaxelE2g8QnFwdGzuwlqf+2S6g
OT0XRW5eZPF0UfjYveapxE3jmj67johbDBpluhyzIzSs8l2hj7hC5uYswZJeBsMj
BS10+06p26Rac+Rtayivy/YIlX23kFW44nJ1xjC8A2ZDhnV6a1Yi8BI7qU89vy+P
GQLst/EiEyAAOQO7kmDHtUsLPGXnJ0Xy8yLC23tNX/JV23NxLZ1BkMYrm4zwChJw
UuSZ+/AaqvPx/5Dh/x7Rlm6eIRQBwMAxe1X7Px5+zgudEKh+w+1Ek80nfYReqGNc
hwPepgyM3buSM0CXmSb1NbEStBipGbFNjiTYDb9oSPK7dDBOialY8F4EWw5CE1Vj
fwWLpf7ziR1kMMHb4FDrdivEf8nAIiugSjU9d+u5K5+Tu92/WXtjBw12ugpox5mQ
whUbivpXsvf9BHT6eVD2ckdvhSc+gjZmDYDH9Qbo84j2A+HcFv94O7sy06BzhiTU
tSnqBkTZL77O0ZGY6PgGWndR/BevPnapUYbNL4X2YUakasudYcMHq+DLa1VW6kiG
LGPNUpqBhz6+Scrz2XbZK1wNSO1qQxCkGF3tLs7R25gYwkQM+y5Wze53U66whxp4
9siVuLnh0L3nfut/Q1xFJqYumRr1XepEdpIl2Xp4qpo7av4fKFlVxQpEnKZrDFL+
LkGgXuz3xJs0OpLSXw6RJrS5/5eYQKYfHNjTcXUgZb5kbQ38QtQqj+oasc6vjCUU
/Fo5yo/tSeLHAQqd5dUV7ey1TqcG8R9F4Ld8ubYEYQCXhNY4+Gbui/5kf0n1EVCP
a3DulJyOVU2niPmnNN4XDR/Meg4RlDnLTtZXq0oqEyAdySNJ6Nx2SfRCMSynZe+E
9z9gVO/S0RBk1cH/X0G6cb79eivgxlMchkoDTsZu47Lotp0vZiTTbPgVatdkju3Y
RDO4/0wUzXxjYlz/3HoZsgkyMrszJUGNa4TxeT7C0Cjz1QU69MKYzQrPVlSyRwJ8
oKcG0iAXPYOQSRZ1fMvJ22YApc/tO5SD5WQeC6tmo1mHjaEwyBsKiP/Q4iis6RHu
s3dT/CXQXY3ILAlWe60EHfTYt4KAXot/YaKeTLkvXWtuAkYdR2281pgXqwnrQnYI
VqUprxvbOqRzZ+xir3rF+u3ozY58tSMm4fpofvXdOz9BU2e3OEk+TAzTmE00vLMx
igm/DEonmU/q1snqDqrov3khswDQHz6XYMtfHLkGpHQqrhH2zr9mlO0Lg9CYXjIg
8IOVEtYKgOKMEJ1pS/XNbWTHJh3QbOBedd5epmU8yLLMigD/ICUZQeBwq1rDGxJO
Q12TZwjASd+p8DhKWxpw2r1HvjUIykUjdd2R9G1Mng1iY3Vbe946TIeQi5d9TUaN
HTeWJP7CkjxrTY+8UQyoiYtXybjPgbDf3tVgAYsica9ESIhPaMr1NJZ+q0/eQHST
8b8T7uZCMmC/ovkxgv+IbTaweVCzb8Zdtb70t7Deg3J1IRhZxRcZaY/OdjPIR09J
1u8ILS8v7cxFwbL+CPnErhklv2kIQyVKknTBzXAvF8kn/iV3tWt+lnRD00NhXDvS
BdahVgmOqUtlPRrdKqassPRmX/yXXR2Qv51y8+dqN2hzNrjx+GReEc+tXsq1Uvii
KVh8Ts4upOWk6Rca4R1diAujc6Ee4QWkLCQ0oKH9BuJunhoB3lwE5WywIEVTFBn4
nTxXgUb+KgDZWjKfmCmwx5d/FAHuifsQjva/RwA2l0W/fXWjqUed2CaSOJQ+xLZb
4FTjso1cgyaGEs1GVyyFlw1SpBjglLk0QcblusjTf1mvOcIQluhBGm/cUHxP8K//
yRUFL2gFa1fh/GF+fUzo+EEJN1EJbrYbfRET3UNgI6gWu7vyeVFfOuLTSsbNiGpG
z0ltZhXKJ6W2Fd/d0ynKC44K9dK6/5eTZDn178P7yXZZEXAdW/FDre2NV/CtfNMt
H+mGGO0uLk0BkBzK/sxJqWEUzI073gzb0t/KBYn7ANgIlDqbR52Q5OM5Ox3p6jNT
CkVZyvbVowHc2vfVEVRfFQiTNuOl3c+VuFdP2VWDkDyriv0gMIhhVOuACDzNUDV1
GOsFdDO1WYcoAbAoE5Xiv2DMwhiZ1lrFPKlfPYMuWAtDLYbcfEPPHUlBR11M6X9K
HK3DSChH/ZOQYO7UoiSF1Y6GMiIrWMzq7k2OCKa/LUeSG75iLFHEzg2xfVqHwybV
vnjt2ceLJZ4eomDUYAhC3nmcFPS9IZkBo/+3h51RlFB9UKiGFgSRV1ZI750IPDxy
qJGIcnA3nDvj8Qd972zTNnfLwiZ7+qTe2wloF1Ce1zZgsSawLdYwPrlajR8bWuGv
apGk/miGPq1vxGfWca2HjFIYXDTfDX4bPpkXfA+uOkJanC29xtLVwTgw8zjV/Xyb
0il1FifVzBMBsmq7VDaVOT69iGi0hfmWs9b9oo9GwqNa0SRwgySrcnLzdt3n51IW
DTGj1rlEgwfYAlvIevX/JLep9IVTiKNDXo/z9dpJlhQhK/+K26ybDRN7m9RuqpDW
fWff/0TWu4js+r5zcJ9SKiNaJqrCgO+YkVFbEKCxHts1fLSjmzAywVfQQyPnRb/d
vi7h0D74sUVZDS9prfYb33ZjM5ak66nXjD9q1j39s9kpNgKw+n1kxLO6pwD3eYbK
u/POnL+TIoORKyy44PTUAT1wlXdIT7iodxHFoMoVOvqOuplbJGtEFgtxdrAHPSNM
fR2a440J6SAdDRgdUb0KWMulbuqU7Z1sUlm+dOsWrA51n2M1vTg4jfsUUENqzgro
2pFcV/B1iVBsFeZuJzhlclVSIHJkRaMAf1rkRcQ5nsWxiHlvAw8C88deCSUsPulm
5okqH6PazCLOkJkk+JuU4D0uCivLSPxz2XOhIDz3jhEmbBSMeZyG0yuD8Q+U4Oz0
xEfs1jK5mag805cpl+qOcnsyr+/e4kpI3kL2ooFGnrvwZ928UnhxYZmq7XwebNOu
E6YpmpqOx3gFkyu6U+xgnnU1gyJkCwFDfZhwI7GLJQ+MwtyOG7BcmMLn8kIm53Yo
g+L/Jt/qsNNCGC5LubooGI3g+U4Lqa1GTg/p0RYzntYAb7kTNaiSR2kpvY+TB0Q+
ihJjbSrGc+/aUanZ2DNH9J5/iEtPnlc9SpdXNd6jATZGfRJ8vbm1ciYk4Ok3htM1
LXmxjDCTiY2CE7naDLL/2OCDlteXRrGZFwvLEb5bV5h52noVAd24UfPgC6NRjL9s
8mAYCSTmGsHZJwiibKMxNuO7ZTIG1WLqPrnFGLYm+B54diqb0/ueTU2vxuBghyxS
PCnAylbxzDH7pY8T4bA5JN+K1Jzi2Z8essQXgW9P7PqHtVYhKsCNq3rHDAOH2SDA
aQ8yZwYcCKuRO6Sd446aZQr6+8ppHe33aWtwUUvc26r/H5kRB5mnwsw/gUGoOvK0
5WIFHueBT2mQgP80CpPZAQjj5y8e1Vb/81kUnMwL3awbdOUM9jpRYup6+wpAYExF
Q2+qZZWG8zsTTXY4QTNDx/bfWK+j9VqFt44YSvQBSFx5YPR6+FIS/C1L/o4+YQ7/
t/WhQVOyyKrVCAEVjHyJoa19AaUYKgwSgK8sgd7n7wFXxkENGVDovxUfI659t91n
qmtaptOxth2E/YMs+1aNtczfsZGLa8g5yW9oLp4IwW1qg6Ca0jFweUeBc9A0Y7Nr
hiITeyTy0lzZfodbym5/JQAlLJ58hioNwz98QaCUp3tQCrpxwe9HlHfiasqFwSDA
VYmUO3Awg9oM746fPPzbXphcyFTMWwA9InZ8HstC+B5rZxo+OvL8OOpXxkTYGYzV
42rVaYo2lH+dDcm6jxA3SHG+T+if7/Y4ERgVljqP6Uy+mvbZUDEaJVxJOZqLM0l4
UyyGSZhQkTlwDxRAuSDl+KUD32Q2Yt5/kghWQLClT+b5FU0C2Dy3xLJ8MxNfrubV
022zJgO56INWAyknvgpU/xRLB+CWR4JALRM8yB+SMmR1WrQMAIJI1+m2mzWBSz/l
5eWO7q+ldMLGsR8pJfgkKVzUUGSNZauEdYs7A1kZm0Zb2OiJHC/ixAGEOBo8yK0O
1+oassxHwc5Dydhj8KKk5ACvNddY8cBPKOjmK0Fm4uOcFkNJRPuAvlxZSWQBW5Pv
Vvf3n8mfDybtUshuAjCei4D9eAW5oIKrxMqI732IytwF3bfySJguQkR5W+rKI6aR
SewHn8q53BFKuuEGCWMSPauAZRoNmkfctp0UDjyFetJaJlIwdKEBCFeCUw+f4W9r
cHSMaQyHoNGA9jisPZ3CJfDvLs/tuEwn/6t9ktS+tMwwLLlNV5Ax3BI5joiQzx+n
8cttTwT3Gx72Nj3BGi2z4vF3r5+IqmCyURBPAoor9fp7dAWUKCy0Gv6PICOATY0a
G1m7rQvbu+CYENxJIQgDIw==
`protect END_PROTECTED
