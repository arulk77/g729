`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL8xdC5TRW/BPyHgukHwxYFBttrHEGXeszfgMcfpEnjGkM
TdFvdSBuifHDJKGu6Gz5pH7Gk03ikTMfpfVBqReE60AtffazPtIiMaI2Hj3sEr5L
G3R+xMC6lYU63uP/kaH/O8YqIQLNf4WBaKcu+D40ksiz5rC/hEmU8kIg0cKRBfgf
40hAfUnLgSatnjPz7uvYLKGGNaJK2ez5mfux3XGbZcdnicwp1uJIeYNng36XMN6i
pbUGzn4JLLWUB+nPHYDZjslIYo//gY3bodp8fOx8RvNmbKoqyoXvMdXfGzkN/SzD
DNVo9S4AeftH1MopB2pEKVshMbQhqhxeH6pGAOI/wbyaqx6eHx0AHUbgY17KFrLZ
9fxlQ7Ezvex0swUtyTjOlJpFl9Gp7snv0MqUde42OjGdj6J4nrxu+bcJ1JJL9mva
RgYt+924u6wv4x7smVbfHNDux1eRyiottj8yXNrqbFAmSgT2aLdQQxnM/Gy/6DvU
finRt7M7weHroCOVols5CrlgKgFRK2AQfpzynD9ZAgij7hC1TEzPRXbMz5/mczVt
7RG1JND6er0SngcywRmRNEKKnpa0KcopvUuYhTiUMr18CX/wRuyvM56/v2YzI0By
4v2myOFg2jQ0hxDOeTcWLOouzIHPrNBUR7DZeNrUYdV20XaYFh9n9TfgqWo0qjP2
YKVvfD/DIBMiFyI7d3XNOz/nGYxKOM71wqDXZXa9ZpJdeq7tGDpMTwEaA4b2y+NS
7abWgE7Kka9dxwb+KUXyRljVb6Kd9JLzV33Oa9yMJg30D/xLlPGGDzwlVicctCiC
qdxa8cFZIlQC8FsNL3bbKNMhP8yeifiimHUepC2DGklNHBrCJSzz3LJ2wiK9eh5r
BwSw2/Sdlm2tzowL0xCAUcCslqg/0yobNBzzSTB5aINFraeEYlYTsdDZF6z+W2xA
FypCzB5cI6byTDyFpHadRExwsZ+7CnxY+FyGG+bMVLBFL6vjswvHCEDSinHXemCE
RnRYkrPBeVPmGpDvEojUVTggXlo2vqkqMZDREpGcgZ0BEVaE2xaG6VMBNrxr7APr
KrVBqR/Bnfmq29kw8Vf8oEY7sl0QSoS7YKn7d80naMUrWs2AItEZnfptqng/YIPq
0W8laeuGZPqTV8qLsrEuCkCRPXbBL7aiZhPHXKo5UX3xgHvH3cqMAN4Ce8+AlgPZ
9X18JbVrcB0wdaOob7MLrFZdi9JEpZZVxmqVSLORQalF9FTLhXTui2Z+5K60AVkP
YetszO2bxIqZzkfAav9TxHdRjh0MQVNBBPJ2S8IBSq0CPUnSZuCsBKLRrjnDuhFc
/EXAWSQkNxk3YuB0dcRLvc5Ggsiez/5hOnKgOHWcUS6pVfQs0T+TheAzsr3bxf2h
BlswSudsUoF7VlMWmFaki+mS1Z3ET9r3doXIQJuq3XyBstdiulbz1RofiHAI5N9d
A2fbgkbVOM3KxIMI9bmVgitxKkYQTE0CMF+Su6IGel3WLNhKZ4wj22eJai6WIJIC
9wJc4R12K5XMP25hLgT119v7evZMDmG9WS47jEf9pekiaooDrre0J9xVkTJaXP3k
SNjtO+waCy/1RTzH08ldhyPenSXgFXQ0lIzpgrEq/wU3RQqVRgr7g7khNz6A+EGF
U+pBH42sbFUWsQc/Y9phkq0qHqDeuG2A4jhUAcRQ7AQ2LWXcKCzpMEbZg4kOcG5V
41uuLxk6KDL8ka1r+kuwsk6GVtD791ybC2uoiLEkEJ/Zz8XDTZC1V27MdpmObIx9
Rawcr0xriJz/zCURNH/NqbfIy1+oVYXUgF3p3GMbmOp5qbtp6LnYRLQ8oLRqL0lL
GNrt20iHdRhz4mAP2i6KuVOLaulxcnj5UxGSKPRAlo1D1ibzYda4ZZM0eMf99BWa
XAKuW8rkWdJyqQEWQt5IXYAZHR+IXXm4BwOys53rn5UiWyIhyn28sq1yhOqu/Qva
AkSryjfFkq0ZzxlStlGP0S6u54BjD9Nec2XkrKAE3LWFmuvwzROk5ezpEtDSEv6P
hYWp0+UxICPSEyNISbx2q4Qj29beIzyM2CyTOdHu50jjDgBHLffQBPBxzmCgVYo6
MKuRSRk0M27ltw0tfdZBAYr6cnbqmRZZC0hkZEejmjckH1rpXzyGoGWdX4qet/Vv
cngI0EVB417C2yZpes5b9JsgjzRsPYKEgdb55nvYAo3LH+YNPPoM98o6JgYVimtf
pHTdmWqDGSMcppd50iwBIQec2Lv+/MWqyp9ixKfZbK71nE8t1k8cWhaYxirQ2ntV
6nUrlWB77UgCazhppp1Q1rvu0U828rkgMGlQsiXG4PK3XauYi5TiZanIFmtZbWBd
gpjZ7Pwj4GmdnU8sqbpWCBAqJmrzfW51U7WW/B/mQcS+cgqxDpkjDSlJXL8qwB0c
x/LFIIJU4D5hom8boJ64npo1/9C18KHchRN6z4Pp/Kxlh0zojPoHSgVaY/dXbGWl
Lp+4GrdlpDjsBrAKN2OwajVlYcDHUltPJLEowLoSooUTnuNk1qOKVYwJKXFGoO+h
5LDVG3ewJhzu1u2zGmclZgSv9+yTI2CsZLCVHlnCtHFyk40MshjcXofUYAUbCAGm
LkQo4Lvi43nICPpGRkc04mcBujAR7PnJ0tIkFqtp4n6hRXVmJlUD1aL3VyVTSQGK
psFgGXxLDo5+Jcxv8mPOvs27Z9Zeu8W6EVfJEHAuMhoIFvS9NRuKI4dZ3QdB70c7
6RqSzyTaBMw7qNn5LRywWBZW7q4wPL6fEVHl/WHHYMucQBi1ysenJnUouihnHDGa
2S0BUjQ+GH8jkloPF0S887/dgTJXcCL8k96vkFrvREz5Uj9MvuZhQPt2PBXd33kr
JtI8by0UrDj+xcFjRX82AVY9k5mAC9UL1LH2VEZSW6GMU+off2flWNDIrjqvz6om
MVLYVCXVcseSaNhErDWhsitnLV241YqObefznwK5BAAnoNDlFroHdjC22Uw4Qy56
qOf8LEX9njU1CXOGL43M/BNhkTVMXorX/UFYBIeT2cfO/ANCxbCAnaVhuq3B/Mb+
izH+o0LHv3jxSNNVsP4NURC/nOR1E5dyM7pHkudf/ruGNWwwivyAGc4I688OhrvN
J4+YrENzF1ztALoaVWNOexDNbO4ppB4SKv9AnbiQRQfAi33DVFgX0qQL0Y513rf7
C1hvZ1N1Pmm0mqy2SRpy8yW5urbaCwobuFiLUIpXqUT5UAjA3LRgTZ702M+qDcO/
VWqhOFFkRXnxCMfd+6w5oI2FujzKU5I7whzAZOg3hUdKS8LCfe142rNtqQeKxaJX
HREIg8bcuJYN2xrli1vVJ6HsfFFyymA6SSHOb3tK2IXE4XmwMZlAUwiyFVDyj9b4
B0ofYLuD7t3k2cDPgg4tIDQZfKJhm3hLRAejjORbCH5wyHKrTDluNsWh7SbKp4TO
FrAKHsBSfXTqem1Ua2Hmie8RF7XRUm8Muo1hcuwrK2oJVlJ6A0/hfAsJlUOtGABJ
RtWrWkgCKB9DCLGPCJAb+pM1SWLXpdbMNr+3m1m1hL81SL98sgW/lUrPuGj8jY4N
UXNQZJqmClsoPbXqG4ov+cpeQi4InJs7BWMaplsyu9Scg0qsRKHo1Nilp3jhe2i4
yuifm8cy7Gs91JxmYZIMZRH91xM14BYG8sRzVKRrpoE=
`protect END_PROTECTED
