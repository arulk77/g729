`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aUPUgQwNZ4mZea+tt6ExX4nl11y6B9XWz7doJ/c+EZDx
Su6CkOMRll89we8DJj2RqXr95oB4xuM15g1pys4TT2r5bClFMg1NM2uyHMXxbXM4
T+IzZ4g+RBZLo0Od783IIJzmvXLRqsNkzV8D2oHwbjlbp2m2nUZb9SAK8x3UR7k4
83IIUwvlljMpAsT/nekM2f55zMmIYhfgb0pKsfeJjm2O42STwm1/M4WClz82G+fo
KBHhjGpKyjxz26iX2Lct+Kt+PjlpsNRH12k6+9fPh2Z92gvwWAgtZLRPJECJyMin
mslfPro3+lxXWPlAF9POVusoBTDxwnibE8nBu8OREQiXE1hUYsbr4k//sA20meiQ
KvVLzIT4Kbid/Fdz3ZoO0C6HJLl38pmt0MbUfdp3x+MsjEzoIXZCWhK4vLeBQYuA
FmlsFJG98JcLnKGzLVpDlJHIiBV5Io1xiCG7WPsOFW3/9nuqWSLD77ETsp/NNvck
Df0aUy2Jy/HX3fb3Tb13A6bN9LeK3fVv5LuYHniH4D2CJRPGD02nuGnDwOe7y605
c+XdprSsnyRy6uHouKv0nH7JZZONolyt7hEB4RI7BSy+pvs+hG9vUC0c2r4m7cAi
BxPCbS39snQeUvWOrc+7P2hAEoQyOAYTcJoznKeJAqveb8SxsFITUxxUXiXxG+Fw
jHtDFuTP/c/RulKatU1wTTiQ5y6WMyYI83pFFdDQyydavD+ts03CPW56Vwi9bKuE
S86Wej9N/vVzuASC/eJj2jV4fJ9SWtozBkDjqPEyj4/R8Ny9WqAlKIO+x76xmrF4
0rTQcVU86aI51uUFqra11oWuMsitU6OgdYWtGAzJbX5IrvLgLZ91/eXJTyG0doOG
EgT/yYDVznjjy7nHx42vW+C5scugUzMXWc8pDeBLTvonybWCh06EAUPhYDa++qGc
AXPiOyGR49lY0Zjv7zt/QKXm961um/yhsxXSgAxOQcaL2mWUMQfm6iL+sj5NdNjB
vQlSKPXTst6Hat4qjkAs7hIOGBK0pUfGsBHQyVXsRO90YXZ0yP0Hw4n4X5tdunBn
6vumzsjmuAEqE+k7VlSGLNOoopEqIyfdN0Ssn85fjwqrqMXb7hvoEpMF+pa7IBrx
+bpPFRFjpgySXVbPdIs1wKWIfLCZIfURqsrR7IAdzHl2mtAuuD6piGfWS3dHKZ+h
Zhq7Hf+MQMOc7dycbFA43ZnAvQQBAC5azmGmppZpoAxaPn+o4044xUQgLjPg5Bki
QfUXZzRFSuWxm633bj029wypvB9V73xjuZOpZiXLuWw+v98AKYdlfuBlp4NGcPAQ
YUHQgkubgsVL+Nm2prAcHBv9XewbGFx9M0lXcQI5YTNg6oSFOgB/zBnb4ODpzy6U
7mJc/bomlycg05u+yzQlWDDuCF2nYJoChGsTFkwBEcqNtbwmaPTYVrtFC7oVg2Hb
JRdQBbl//etIGxgjKByyXtexjOAzyxKGNT5ebZkBe9GpT64mRKKUp345mVEyxTs0
es/JhK/TPyshwxjz52yr43UkA0MuZiI1OuNJaFupGJu2RJuIt8u4nLU+iYzuDyL2
6A2pK7y4hzqIA3tUOJqRHLHW1TxZmPcJrkVZxxYlsIpCBhsedtJiFyHEm5s8WlK1
vxjbSCkSZfQ/sw6JaL/6ddsdMYi4A7osCT5WA7TcQM5x+cP0dUDXPMTjbMdaFTun
A5XwiFYXnT2MGheAsEX4Dfy1RBeO8eiDNy8r9Mv5K2ELm3x3DqFZK0Wj01YmLu8d
pvDmKrBErILgtEN0BNUznJkep8tT2EdU09nbaYLbOTe5ddEH8e1oMF0L82whE1C/
szIXqX1qGpb+oxwxeSZ8q8AfuqnXab7CIjiBaoqnIqGEM07BRlOycJLUVFGZPEsH
TY3Y4LCqHEFXMYB4esJXZx/vXb0tSj6wl9+ML4C4HmVv/So+shyO/Suo0NS+8WlG
GZpEQJrsKjZ9g26BW7GugZKwxoS5ZbITZnh6miyTMksvQrNX6eEo1T93JQvKSTKK
/Z8yo7v1m6Cz7Hs8bp2252ggB4UxQENHxY+XS+KHxXI65QQNU5/zr/NtdGVH+pn/
egvX/B+8CA90M3AkJqfkvNxk0uBZMycHM5jVKybfvd4WpcSp+Cxo3RqEBxpqL49L
1OwYHfIO8l+Fa3UgAuQFgY3ouynrnZfyU7N2KiBPIM1wOyFf+zzeCvutj30+qYrn
+m2I6WGrg/AL10hKGOsnHd0ZtJpr8M7oqRvZSUU6GV5bt91W6RL+my6sD5Ajvycg
xCPhYR8QORlSgA6CNowPRRdUkWa38bnkNikHIu+0aKeixZl4xJQ9NDREkaGsjoZ4
+g1imJH7FpVFWjGyAldKCuiR3f42KGA/4yGAkvf72vzEtIr16fD88FHpGNaBylDA
mwAhA7cnQKoBYQk5EyGwlQfvmqZ3jQ4HRBtYlXTXoULXbCjNdvJEuXGdQiWVLkUz
c5UsrHaIZOWzmMDvDTCIbJGD8EoRkQmRfXxFqPwI5Vo6FHin8Bho82VPl8d3SG0R
Wbd5EwNO5AhiaKo1rVVjOvayWqpK1noC81LY47xZq0sI5k7uRZslGIf+xgdRIJmb
/d3Nro9CAk5RTPw9UuOG8qTReg2guJxrHoWX3JvsFHSS9XtsdWqO675RJOlgoR7L
IXiIYR8tuVAx4hzCoftZyruD4dR728AI1IPvB6fT8aa8CvOaDdyD98TDVuHDbdT6
YRx1Ma1y4+8LBwSQlY0zvW1faP4p8C6uHyTV3rDp7kYWMNhmwVAjH9IWLthw3YGo
gIkHwYY/yKZGqB4W5FOvA+DjpbHfgA0jLLu1A4CjEv5q31IcJ7XKYnRJ/DZ1BNhB
3sppc6XqH+cb6G4FoR3NzoRHQKzebyQocRdNAsPXyPfn54sSSdj95K8UvnwXY1Ix
2gjuIx2RP+WMDz0T6joA3xYpWPAYx8FXb3D7WlmVx/Czf66cBKcDnjEWuFruWi84
GG0VPqGOnzL4FSRgkFncKncK6TItyp9l4LSnrQ8r8Ua5qbRfP+oAZJHUX2ZtILLM
sxxVMOCcNsLZD72z79jg7APF2XuEMTn2hgut9vMxls7t5PzK16Sniaqa3eqp0BPf
Iy83kLe2EF11qycFvKtvHNmoZNmPIx5OiX/z4OajtHZhlhRrWDOjhODidO+7wqQj
RVBHlTdg/a3Zb8Fq/DCB2Z/0IjZ4L4vlu5TsFw9W3B7+5I5WxpdJy/mK7uCxuaXg
h7qwpbESbXhTqosYph6hP5UkOx0iujfWlr9OoP+7zFKEX/js9k6BoB0mPWmo2PLE
gH1a/HN32je8OdM2hzvQ3ztfDekw7MccYHsrtpUKlKB/DVWx5c5lZsTIHQspslfu
RLvyqDQ/uC6as/Iqv7v+1TJwCX1n9ErBfSHZqBCZoSR9BHTqyuLRE0/tIWsdT/BW
I3Ov12C1qY7TiXj1Y9kBTSHinus2pav5VVbR9TWERwUm+xkjZdSLqOwB4w8JSX8k
OcyK+UVSY4fhPaBcDAWmXXJ1xChlSPKlm3YJoFdisNeIkgNQFwhaA62F7qX425hF
U7i7qsCLtDrRprV7tQBQ1pgdWzV4Ry+H/BpEq0qEaoYY9sf5Ho8WGMUcho81zC9i
UDoW/QjixM8hVh4g58s1p44RTNqkrm/d7KyNxjtFqVcn0oFiwrgKNhsFztQC9rSf
clA7DqQKlxd777x47zOgmB2+edBnFVVdZ3mgQhDR9oV11mX+DBHEf3c4XxwqECxI
ocuzAfpkRl0gKeGntoh0XiY63GymX0OtApC7AflgCRz5KJmelwAsaEHOGb2IP8oB
NDh4Cojbdlt9yIf/EGDZabA+thtxCI7GwNBBx6zVYNNE3t3Ga0wzoAoJ5x7MyGG1
usB2Umoh6+LkxPB9OwOxdncJCwYzqKbgjtU/kyNWSWl1HMkk0OxKZazoB1jqrRFw
LYFfTFqL+RHpMQ4oAUtTwT3fx5zfr+3dbv/piyYkzwM9V5GSohkp1At+V/Z+ojIK
RIvYjn1AuKPGTXA1Cmk6YJksWXSuqJvpEsJANOJWtCT5W+2oeAZNtFW5IPsFn80A
bXDLqiBdvYVn8bctcTv57Xa1L5kemavI4U9Qan34tqlYozwYEQMeV/d4PKqmidKu
NNgQ+hBT7rs/mGEW2uQCJMzPYK6YxStoIoJD1t7HwSf0RwoHj0l0GAzNqrbqyJS+
tAxMkun6lasDGLuDgLTdXDPwGRr1vr8CzS+Ohi6IyJ32KiY7dD/Sa+CY8hbWOzMW
JvczzmhOf+a3uMWkxEqmX90kLkFFQ5ZPtMkegMAFyd2qnTt7wSrAKF2Uj1GIe/Yv
VquprPhBSIooqW3nnYALIah0mnH1cuG5CAofzu/KYS4YouH7jM47nB4jEhS98cw6
fLkOTgM20sZFduw8eis2PFgf0iP+/xrDowH0jAsdC8agJamnbaaH8ttX0bTrQyyL
tSTV9BEnKqw+uql4ERCNoXPYKm+XV8M8DvceZhkTixptVSNHt1wEoIEY56A86gcb
Cs2cdwzIcdu0444wNRjz198hxqPnNS3ZET4PjbWNciymXAI3gd1XAPAOKFWNYIWN
bLtjRkdQP6oDIll/O+iS+wkzSWe+H/wgy2yPVADjc55Ng32NQ4fX4Ri/QIKi3r2y
3rfhhGdYNM1pSU6shKu1eTzM3xopLT7f9hb0nm/o4u84Pw+14oN8ZTJneEqFxePN
Uq7HvfRxuLf6To1901+jwoxfpdzt0QykjKe6tfeH4pkgCW3xFLyWfm7sE8wWT+b2
qdvvWFoB/hSMMDTiz3HVQV55MHLeiRdtdbA1DRE5+C6xKpgt4LdXjMXZi0FiwOzz
nsIQI2cTm+NVfpAv4nu1wLFroWStQKdjNVEPddazwW3ZSuVi47BluEuD6Zb6MZ6z
v4KBmOXlb38gurEjUsDQQz0zLxg+L+GQr/95AXTL6n17NCS3Z1zo2ytr1Hdo0v/B
UAsE/CzfrRiTFVg6TCTAIU30gq6b3VMuhmLdmr/1j525VDAAF1PWPCUPe1dfVFTo
gyv+ftxd6RySwLSF30Of0xrFAIBdhGCuQIhGptz0PMh7Szmxb25PSjTOfW/lKkda
2E290QXWXE0e9hcRjuCC7k0YsHaZuaE02gLiYF1NIvVQwdmAWM1lCWFjI44cyFtb
NCgNSJEnPfTPPdrwL1If5UEr4orZH2GMuhZ1z7JwfC6vy1m2E75y2I2Ps+TXnk6Y
SA8tcJspqPubWcIz9hw8EMfo0Ekpo6hz9KjWvLG+TBq5vvPeVyX4WZecDg4jhvcw
EODz8xvLoLZWGw+9k6jzGj/V0NDz4Z3hUKaKrivYURj0NIOxZI83s3I4mWJyFomF
W4WfdKJ+elkB+G6CJqDNciwnpUujFDaaglArNBmZmSJxFEOupbjkOLLUJGJJM+MN
VOZpGLY4NJCjn8XrI8xwEokEiHAfSG8zBASWcoWDfDazE8q5crXEo2MXyiGXCMtb
NvDtmb9kplVyWMJW8dqXv+dc/wel9mzlIXRLM+3txeVhmoRe0PMafEJhecCq2geH
EvWHZhCkiMk8KW5KUShj+3DbG8aO9+tQcG7SR/BPwNfWEphQocgFOJhja6POskMY
tarhijUNFOoO661D+Bj6/w==
`protect END_PROTECTED
