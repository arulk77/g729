`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46N71z+XHT5cw280/2AtymgZSLqGEdTBATBW6Yn9z9we
pP2zeBZmWkpkM8/UhDyrqC6ojwr5LtGRH/2ejKpDxaP/NNUfPtUpNtZoMs3WS6u3
N9lIhK0uRh3+4aT/jD6ew4NudDdU1ZFC8jiTkJ+K9pgNloBCGccI8qrQnyz2VFHJ
3FaCr/kTrpkYw12H8iMy+cHCmluraJfhyT7lISQTiAp0nDQtZoUjYMHMmkUnr9jX
y7y6FNGs/eQ4UAuRizwHLFmaDwTZ4NPokRMpNH7MMrCeiYYT354XwjAn8wK7PiH8
Wg+ih9Y7HbisGQCBzkaQVMEPcPjcCi3vf1KvEKUM9PeWsd27ZMm8/qL7G9T36emt
XIfrWX9hAHKD61zlurShXKQ1ZPmTNndCBwXRFBIkuYwPd+Q37RmTAqW+bwHDkNSP
ByAZsOeUcog6UpNgiUEJMXJ+Rgt678ZQP+OH3MmgRnmRsuCU00+b2XA5QTFvKpgG
EExE+vgxs3lsa7zyHf3JRM+LDDY1ATkb2tPIYxJypq6oa8jtHmQbDgQaMNVMHnwu
v2KRjxL4bgg/6VFZMAgUcaALlnx4Yox0RWYxBz+obTydLKTaIxqWyB4nR020ub8/
uDWc9vWKnfMOePwmbtMJ9aAlny7LlmN4xjSfOOw604gnptPs2StGUCpFe2kYpGnU
aRcBTYdxkmyO4bWaElt/KcIPAhY/yPj7vQTGV8JxEL+hKmi+ntTQO1GcK5mFoE3+
jPO+1wRhSf9x5TFyp8GpsedSjj+6ZjdVN8BG/vCz4dQhr8owCcghaGgoFyPpo2bR
YTNHmHs2gDyJz2QgcBekyuTT5FufEi+7RobOkXCFDOpE1kZOIVKAdKFhtitvmmTF
Xab03e5sY8NzQsr8LjePzxA3oVQi79txzfQqRogfb0/pfojQGhDA4FO4eJv4EO+M
h4XpZmP9mKOPDxVz62s/YUhxl87QSLPYIhsdpP4L+u3ytqT+aYvcU6TvApAVxErM
593uqlPvkrWMLgjjy3iwcmeHi5u8L69vYgkzR7rSaspUXKXmHr3UoLeYWd0K7kDm
LN52WesWTaxGdGs4ODsRHNVO6bobpvMXvyT7KlvRAMNcQcZlyJnvSNNfl2MMeT+k
iYA16DzbpWbG0p3mPpIzlKKqlYNq8A1UKo0fa6EM/BrArA7DWM4DBi9LIm/0pbEE
+HNOMlhZ0b5Qf4CQPjmfUG/OtdS+KKVzrZZ92JZ0AmRjsRMv+F98+Q+w4w/kFJeq
AeosRKAby+HLEnXqhCqKLrSNvdvPnlSQLPlD5U7lvS35ik3xE8UpDkKsjBLyJknt
bywDT2f5ucGbnVk+DIjUXEwSisB35JVGhvotfEmhqkM4rpBx4wxiyRAwzyP7qb0X
BworXRidYyJ/yKAIuuJHqMW0TBxHNTHzd4d2j/oKQLACf/+uVAIqRoZdfqq+I/T+
yfXvbxOVLei4eo1Hn6LHvd9NTK/dgQQNLiQlKntWkcfFgUelXQtha31/3o9vUB8G
1jJD5dA9DxQibvlEe1NTovVzlQmH6nsQuufVso6zktmzQGQZLLgmT6H+iViqAaXJ
YtUvNz/FFvCzwfoBBKV5zvswIIFh6rXK/8jwdShqLBNepcZ4a93psXeUFB6W29nQ
IqeV9Kam44RtvWWV6Vuu2+4bhGU16Qvp4qr73MVefc0FK2Ne9qNcZNGxh/GlpOjz
sVC1pBsx9BiCKCmzkn7qRzmZ/KU1EoZrNbblpnWJTujovPA3nUd2obFQAoOH8QD6
`protect END_PROTECTED
