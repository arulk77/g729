`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
LVa/rSj7hvdtNZCd1KQwburIatSzRdmPjRRTxzsxdjH3As/5I1+xR1eVNqERkfeN
NcFP29fMcD/01L3aHQBFvptN2GLVqe1otoCsCvN/7DDpJNXGtoJqCdWDqWgo4qw9
TnJVe9yzqdA11PxDAH6grlhwImvemeboggnn+bNdgKZ3pAa1aDd+i+5pd/KiZ/QS
Om8RqZVWYS454PNZOGe3gqOdhK9CR7Rudjp0yKalzcDNubf2cDfo0FWKRMtqUZJT
SOMqYfUp4O8JBLwZAjwIu3p0Dupnbcwc6e3mx4jx9O5zQWF4SnuxyZ7p/V1OWq0C
qxFjoG37hFhRIV+j1xoAisQeyZij+RLUyATVoy6RGbaFCtzEF2BFG+NqN7sjqCSe
goL2Tks7kMKHrS0NSW424cH8WJirPe6lGEm7WuJXh1WLwxCwMUywUTveFi3W0cJO
k31AM31NvTGKuNu4T5KrjBG6xDfqmc6TViCC5kKqvOzWCientPfi/aBAPqcjrJMZ
b89AsyYtYjDnd9RCMYbXAQS8nGFNIBC6fCXgOCnBEIWMQ8JQyWWAArCYcFrdfwVm
GElB/p+lJnTCBg2kajVvY0yHSvRtaq5RCGzLAv4SuSgKs3kQgCy81caW3ZRmEWCK
fxHbfvDxG8+uaxxkUn1+ywY4BqCphjHtEX7/T0t13SVCghPG/2wCWJNLzsSwwvcv
WB2BR9gZFBLJm0zk1kbSFWhwA8Dp0CQW2gItpD5/q5eZj6OIxy7XYgsfosYomE19
MoNswACab6snQeV1sVhhpDadKmbV/qeAvT8XnwmB0sizSxh37j7CZeuMQiTvLbe5
dK22d1sSsCDErQCdleMZAXlceh45aVHcx5QAFkQKBPw=
`protect END_PROTECTED
