`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
s2X6u2oN+fx2UEmqIhy52AWjENOwuFFBRuwwcEVwjkz1bhpccI4cNSdm4nhoDusL
S6OI5e7nP1lLHhZbJG45YSfC27b9RoIKYjAPG47ieXB1c+8uZywq5L7dAxgVyd1q
KYGV4HMdCApJBwZHMcSTDjoHdTF2m1TQAwwYcIy2BBimdxAsSLE1s276qTJ5OQNo
+j+vKi3KxQTWSEgdEmaaxDR4ym4efDXRYWcZLtsDZa6hIQIgrnNK82ov8fIYCDb2
nGrjNQl4Y/DskVZnwwqaJjgpQXa2/tMnKbesPUZkhYzeeZBCwlBGKNh6kljMlHaX
waHX0rxlrZfdIztKvms0vLU81zigCwflB+CUr9XfVH3luWb0EKXAcsRGjTShUU+g
sPzxou7Wz2Qf2zyJS9r/hpFO346ISqnkZocYd0C3iG6kYiu7cZj52DCgQwRju1oe
1mfZIAPnQYgVuve0ffjzKK8DtdfCVNpQyBLe+PWAtE7atjl9YTsBuH0fJoNkXDfE
PSBkKNOX0FRHA91X3xMtv0vMO6t+lstzS/yFVM1S5X3gKttIRF86md3hyaVbMOql
qKFE9ta/dnlMZggq7uS+AMx8HeIkpBOZvYn/8E3LUHY+PxrgFP7GpoMUGuYnwrnB
lDp6L8Oyz2eaOPOhRnLgFYzzLjKI1/bjcZKSk2ZjyBawL6z3oDy3VdJxdDAxrXbz
PnkFujG65ngaqXLT9uoGPKei2qRVjcWRaG26I5m0UGjqBQwRUEpoTL12F5rOGWzj
FC3EEkSoQ9LRslmikrHrJ0/BCXj14G/sQ9/X6AEC5VmHlVE3X5FHRe9flbP0HCwD
ikOkpz7YfnslPMRx9+uGLfvlWCmdiNcEPpIuzddL70IXZkm5vcy3r3vnL6U67BMp
lBlDAQAG5tStBmpOQVPvIj63Iy5zpGL2oS9blrhkd1FyOCDtLQif9yGmx56DeIhl
HxxxVw1h+VhzMAItr3uzF11btEygFBD3ekJ4rbmI4TzBIpzHRSMcJhW6p+Pc9SBN
6AbWWAk46NOi4Wi7fe98XmDxmgZD5urRtiKtZGHlnrXSaVOV0QY/N3f7FeKD58O8
vsauWIdnfKmr0ZWx6Sl5mOlaZHVMnj2xTx5fWGp6LaK2RsNnIeyLMDIKu17pEuPi
OizaDTg3GdA4+gw4V1JYcbNQESOxWsuxJ65SwaKw6NHcsifUgopsHFvG8NmIyIL1
P+U/s81IqryOqpWRrE/MWsUvs0K8H7UEL2W/BNNHcgX7Tf85EDHkuc6f53l/h3ik
gurHGIkp6WZVa1u5Gs84aAG6twiQSBnBJDqbHuH3N19kSdMqe4hY2KdQNSa97iEC
QbVBzyan9lulmBWTQlCja4vPlStaKNpnhQzGZ0ECGoI2K411cbJwsTG79ZkXhTej
/VpFiyfn6ZXoYUPBids0479pIixjae3YzfPspGzAL/sFe26vITdK74p+tcoJsF5G
u7qZQIidhe1ec+bIHO3v9HM8ONmkK0FR0ywsnMGMSLNkrgUwTiyBMrc83YAAGbB7
gPWvHokm+NerrHF7vTI5XCVlaSorVj0/IUNJ6V/NUwlO3KAHe73yJE0XwW0hKY0s
V7+R7xUQHgnDZatslN9mWYbmReR7u2VDYSj55pR9NS/1T4N7FCwFeDisPB4pIYXk
bTE2WvNWh0SZ3Ndxinre4YbHeXabClrE+9Uwf/hf9mY1AxWvwajS/w1jj8usZMlr
WqrmA2dnzwI/PqPp0MJC/b/9GPK6MvsdLt/OYegjPzdDO7q/xqyYsQiUeCQSkf3j
wGcAcpvQ7NFzjse//FMdL7Km401Pc4IrxzYLaYir63w0KvrO2kzXlrgBWvXk79QD
szuP0IGe3IYIb+PfyN1XEc5dBnm/wqJT6He9z8L61XlvZqaxXklIzOy4dyAxL5ok
qP4KVu8Hqtd8934oLylIAErnnWTyt4tHrQmfSJD3l932+Om9UfOg4HdR95cw7fVl
TjZVhs5FPpTULxrLxgNo3yk6NKMm9c6Y+mosUm1pvOnVOK7oG7LhNROo6DwUKCOE
dgUv8a3zbcl+aMG7nTi3czWR2LGGmRrSHvyOZ9/9b7uKPAIs5n92+1GwOKAvD1pr
PoQ80Kxl4G1HBPngsWrAld9uaDQ9il1za7H+1Z+VwLrDQPOdnx2VkYUpVkJzzt95
zEeS/ejRuFjsVyK4zaPR4h/YdbVDNwgEN/L7B+mtAOAngF31S7iH2XoOiv2WRC15
eWWucw/DpethYlAm4foeIS01QYNUboDW2Hg5ch5VIrL/RqcAVus4dRj9++nNDaeg
jo8TN2zOHwXpB8xB0cm8uVczPsfmhSg+Ef4Ikyuc1sSKqoObVIu6botAQYjtQkuQ
8uyzyxo8pNEcuDXyi9OtbM0ql9T55YHLLA8K8NxlyyCqU9q8MVPixgfx+ZxIqZET
ay13ZDkXaIfEPcZkOEJGVviYR5uR2zm7xqy9mNz8xGCWBJIWG/loxruYUB5HJP3G
m9DEQ9OI546EO7wE4Z2s9um892AivEwciYOl2PVCUaX6Rzdk6snRgoLtHNpfMZeT
Eth2b4q5YTLEhGJJwYZZVsYbl2MDN+4Uy2/LCKDrp0i4rQEribUJ+W6miQcAB/0A
Xz6BlT2IXbKD88OELwnLUpVL7zJ8breMH7qRPuC34x5Iun3qG8stHMiaOPG2P7iJ
0g85Ttu4BbYWp57Us9ccOqr7/W0lilPat24cq44BSLiYxz/PdSwWULClhcAYvHPq
0zskzy35d5ephjHP4dCEM0OORbiU75JuJr4HuLrpgMO8QlUpZEiUgmZx2j1I8i69
tIYzxX7Zd4N4Gq0hNSTMv5b+BD0KBRSb0HIW7CQ23pAMcFGMH6lzTStNVFoYkG0b
zQmHCeTQwSc/nJHzsQiWShFMtPbPRzzKZX3QQilOblTZBRhUhk3m8vPH4nJ02GVf
wOmW/iyn8MJDRZYD6Wh9ubTS9Js7NtkOhaGbDZVO0CLvbn6WXL25P9nI0j4zZmYA
BGHM/QZCFgUfDxJQvR2D8jUndxokMggr3u0zCEjLPiik9FvyeLUS4Ex96rjWJrXS
2LV9AJ3H27pgLTCK+rMtr8o0mIRyJs3A5NSioHs/jfM0nPvocg1dHl+oGa7raH75
WteO62d9EcgzTY4LXSO12hGxdYjHuQeVhly0j2rKrU2OkTvftUnArqeWAXIPuUQA
ElPVHzGkah2FbiGu9xz/mP2iNMHoJneOvhORuyQnS5A4L1eBKttv/65tYvMzjBMb
CZsU6s4BmQyT7q3W76bOneF+76pE0evu4Os1rdmkmLqBBN/HYdYCODeK2dBc429R
RsOOI75Wdl+LfWI50rrD0A/IUANLdOZf7G1arwMy5qnom+9B/GVy+oKKKHUcSLTB
KeOtb/hjYjrbX+JTZ3LYfVU39E8siQmqS6cNlZBYyhqLOVtiuhu+xUI52xrLOxkv
6Ts//U8h7rS7YdzlLoFM6T1OOAta1qg5ttoNYYGyMJshhPgz0wMOvLW+m1njsL3v
Xe6IyY45Jo91urUup0YU3nHwraPXVYgPt+PiX4sNCNmL8W5RfCy/RPyZcloiudTj
/acjD8hHPcmXR3F6C/DjMEDudjB9C2DfvcJWZ3a2C6vsHR3pceyVPjGDOL+1sacj
+YPaNiU+XBB28QeMDEec9D9L32AT5TrtEGT4M7qQoVKXYfT9Pyq3c6Hqr/2K3GfA
DApeBdgV8fvPBqMaU5IA76yi6TFYoIS262HxmCzDxAXIVA0Mc5sCM+rXSMbbqudM
+C+vu14OhLHFYJBmptQe27w90ewurFfOUzlZwAQTSWhRYiP8nBWaNTs5ZH3qwT50
P5cyhfgeXR7NYjTr/qmQma3yRJY0EC1SjYCilqI2q9V0TiuDXCczOQYzQYfAfB4A
WWbd/7oHE7qrodmBbr1bA6JMh53bYrpzY0TLFjqrIQNH+CgppaoSCQ//JKgn4swt
asQfJZICS4IZXvah+hnH2IxQPlbtF2ATfFaVaYgxJny9zwQi9b2petnqyvX9aCQ4
9dpuAMzHjPM2Clf2Ky34z5K9/Jq5tAetCNjrl/z5JBFv3xnUW1ZlcHpGZ8pzRyfn
+VpqDpberumynLoM8FGUOFxlJJCZPlTcXlzsIgqI6TzqolfJnpUf7wBL4D7qQPv9
AlCE74Iz+n+pzgyxOw8M28ST8Vcs1N7YLPVC6XiRuEyAwwJi9cCdq1cMnL8dwVIS
7AwgPKhq+hL3y78i4CUqw92xZzCKa96Y0HpHpqNf9D6iwHVg4P/eiwIwxFtVbEwU
Cpn91R7cSLemLOjxEKzgL4ye+E2P7JUPeCVaN/wjFNGvD3+X9p6M0OP+wZdduijb
2xT86UnnFjY5NBB9xkZL/E2sLJXSyASVktfK9q8U1UwSIkOa9Posr9U/8nz7iIAj
hFBtrMHTpmtl11rHbChaDJsqkO2B82UYz/fahsGE2+759898TmCBEdfgKEkZQgSP
C3p0BieB3ZhS+nzt1QbOTvO4JVSkAZafP72GoO9uCT64puL7gx9FVgoY6gxP6Yix
cHDh/gFzqEemBHQ+CO07snymWUuub88CZZgBEoy3+yXSan1pyXZ9W21c3xEL34NI
9S5u+nGpbiR1m0fZKCACxyFrcFL3HMxBa7g9cuRnR4RcjL7pxhyQSuM5Ulyegxf2
Pfam/qz6ZhrOz9YUSSKn3z6MHmFoQLY4Y+SrYqK4M6KcIJJ2HeDTN8lCO99FEkm9
`protect END_PROTECTED
