`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNyclb/qx4+O3KWpn3SnnJY10DKYLecCnDnDKxMeiIKec
8tvT61lGcxiE5RNUdvZwAXiWkxFOOf2CcuUNC/FjD+HVp9xZOqIkWXEZJgHO/e36
OECgV4KxGxrVC/myjR00qjBW3fR99X4XcUWb3g2riwkf2SBpokG30sg8cq637v7W
IDE7d10WHo/5UEK5oo/XEJk+UmW/T3fgMO+hLMlBkf2o6+pxrpGEKVgoyrKWgRwm
PzseQ+nUMUcY/37oz9Q7Icw3a1T95WIJ+/GHgjn4J2Q6ykATAXchkZZru3aQXAjk
+jYDcZJWDL8Weew7EDHvvtdeOP+HTG3nsKSNYtQtzv3mjgWYKkgUPQeb4fp6B52B
qWujvZPX0jxdhohswc2ZdwkDmTtUZFiAzsHCe8l2KMo+O42adyyDcG5f1ML/4lJc
OtU2YoHBKVF+HNu5/NtbWGZAJwKop5mD6Wzw7P64O6fmnlAy3X++IGLn3k5FLdnQ
MSRsV3iLValZsevGDG7VMXFmfcRg0r5vcgnKWbNu8RywG8zdZv75s/FlyxJgGrJa
Vi+UApVzgkCE3hSYaxn3m7h9pQIDfKW47gsNDxWg2vhNwJrInTBPruOoVmRnM6hZ
wtJZSkl9QxNu2I5Fh0RhKG9Bm+WYwe//CxC2M9B4h+IfHaADCobwLKTbmJwFVGdR
C7TBzLTV0/5xwmKTF51Iriulpx1a4NmWPKJr4LPw4zC6pjyQh851/eDGMJO/nJ3s
EokEpyoDcjcTSPBF/XHvneC8jIfL9IlNiwoxJKyaMVXasPjTE/Dm/fnSL8ig7PIT
o8NRfm55pGjhchbfQCXm9V/J6efMb6GyJmQF0M55b+c1PlIJJlIvJsgrfJA9ZVgQ
iJ0m7BFqnXAG5epYzgD+84TIaQ7qvwW3BFAhzrkROfXQXPegcUGM/YLns4qbxaq8
MWrWdQNI0dGlPXnLcuO0HBUtKs2e8yg/Zt+LKuXQa4M=
`protect END_PROTECTED
