`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLC/JYm2+2zaKSx4LD+rsfoccuSUVQ/TOWz5Ye1F7Mtt
HZrhAS/uU0E8Aq2iSAs8uuHdAn26T/vPLoKNrpWirId/3HHYyuE8IxthIFYJ4NV6
zo3NvAYXor9WaurTgz6IsHiRZWzkFi0+qQfA1ofRa1aD2aTplqgNtmg/w2xPIiHm
2ZCqs5RtU4jmeEjXL7V06aSd+uXVJsPARZGLfi9AWjVC2+kopQQmEOymawXXqhVR
Vkwca5JA8IFpUE7SKTVo//Znqv9K2NEVUg6Zc4VuAEinvUxkcyJCNQJh1WC+FZsg
Tm02P8XYf0ZJKKlIPA3mzk49FFHxhlB721ckpH5j/IZ1Z58RPd/93Os4zy96LBMh
Z4C9PoHXGaFNCPHtFwrspwJaW8RUtm2GaswRt3/A4pNdMT+P5qDJSEJWyafWuynI
axnZeGnMFIQetdgZ1qCLSb6DGEfnXQjxAE+zUf5C+Z+vL0cvOacEFZk2NkGVhDJ2
7dP9eRPwvuYPBCef789Nl6BJXaUVUDFWgbsPh9ABGeOMyXfCvIgtyoHdGvMBA9cS
iKhYUBirtoNWPtaSFsrg8xlXiE2MNpgZ/vsx4UBFyXiMQOLB1maIelrbRBRLSTwU
bpm9V11iEQIBZWnvMQ6+GWoyNKsEOhDDF6MnEltz24IJQMY2xgAefaqVP3sIZx1e
6S3h54zuiDWh2gsHyE+EfTcWpksKNvaUJmsJfYH+sTilkFV28Pt8jDkJcyzeKdZH
OGNibfgPd5w349IjPuPOZppF1Y8TPkUlh1UE4JNVDBhesTWn9UKNwdErkWrPKtT4
533V+gM7sOYVJjIabeqfqLSYQT+yWKmKCdWWoqczRdI=
`protect END_PROTECTED
