`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4jUYkdt5VjR8oFbu7ZiLkgWFImDkI6iB7DYuMS4ipjvDRFYzpPZ45WZr9XopwCcJ
kdUHQxqViV7AmbusDB6lD/t5JzolI7nDklp4EslnStUUplRTHr27fv4CyUq6iKef
kIO7Ud5PUUXut0GDtozCdze9I6YuRcmf9ylkAL9w6rtjVPuOQc3RsJF6msHnD+kO
1wsOCfsAIwBCf5RYcItbu9kXjfBBFZ7cTjavimaHj1PcnmRgEZVjlVT88+/hx7RI
`protect END_PROTECTED
