`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ZtuA0r9nLUvY74CVfMikKlNwdi/9SHIXtJ6HdUpAendvO7bAurSM6OzmF5r60B3n
gXPYVqpDjlwY+RquZ8b+jXFeTajt+Ivgd+vVqovVxnEVeimpAjKiBfro9Xo006MB
Ddq7gY8DpFwhhMoxfjDmcSTbe4T7GgfEoxFsA+9CiNg97YwiRy2eG84F/BLYLx08
`protect END_PROTECTED
