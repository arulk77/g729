`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHISHUFb5eDLItN5EAaEh+TW+XC3P99NFiViniFSwXBI
/T6x7qHBNmoHpfFNKXvnJ1HsRXB5ffTpQm9wTdkWxM/yJmwK/Hiaah/gfwfmsFs1
idQPhpWQXA5owovThnRyjbq7wSIRp1bOllEIwHNcC+IjJ7o24isJ4r2Vo5oIahAP
4UaC6dMkemBom4m8dpB8qxmG+TqomE0n+VkL41l7qqI2D8ZHAZ/Eo9+7k/4BY4QU
c2Qd7DYeYL+yqhy+HRKpBZVPx1aGFTdRIuxfs+clYYTJdoB5kUWw1l3wfvT9fOB/
`protect END_PROTECTED
