`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
g7ZawmzwoRa3Hw0l4KuUfKL/4dPdt/C2h6G8sf5rEMs25vIKsD4gRsZQj4PyUQyH
b5duZdHyr6rhZ6QTBhAgJHU3aqCpI6wq2y2cAX0YVrUSf/2Tm+IxVBBDtaGID/oQ
aeltEX9ibCBlha6S9IkeAalJgc/mCttQBSD0fXy9WaOt0YXbe8xs5Q6E3Ce2Y6oE
XQBl6RTlpodXLWJkYBWaCcqM2Qm4R4LJjEATlUyx/fRFYLH88j0pajo9rRYOe1hh
sDFsekrvzl1XQVg0l2yrmmXD7c1kjOVA09pYtZwbPNCt6riuL/mCgrm9iRQzxuCE
RC8E3xCQGcju4puXXLghiIYNyETh/SXCPl8EFob3WGj902p+o4YmjeoLGsWm1L5U
1w7caQtsuPPTT56+981RBSigOQSpsHcreHBhs9n+FCRIokXzIiG+w/FvG/uf0gx0
tz8+nAZVIY3f3lNHs0Neyks9MYshtLKbPZSO4ks6aEvhBxdiK1hmvPvV1lMhpMOs
0mx+zCMsVVaM63hwXWMSAqce/yWK/tEcwkAWP9qEKN3iI2dvWjjcjox0MgVDDnnD
xx+dDFVkG1QkT2pelUKLIYRhlNMfwCShSL6dCuL82r29roVF06PhNJA0VqHALmDr
pOZZePz1mWN0tycVgXwSBoo1gBDbrTAlSBX+sL1oDmj1Zgo+O96riC8Wq6Ql89pD
Zg90TlgDO5xJCCwGU+y8y4yUpANVl7obolgH7SAZem9qqeSgb210eHPSXYMIC6TU
6WhUsrHTp2EjXNsfw0zNzDdq6VKc2f1UQC0YArbARZ4oYVb8lI5UQugLBLYjhIq/
XectdaEKad4ujCjKD3sHduND4q87av/nswv5xzRzgssZ6/LBLKUCB4+ChZa9Lkgt
P91XVkT4/HNgO9wAFMGxXNKq3/cVMqdggw302Ijv9rgfnJDbrxcNddg7+QZSQZjw
ZQ37CF6g6XPnYlsI3VwFVd4NN2fxPuOSyCz4tIEnzaGPH1pOFGrZOcQElL1nc6XE
8rZdI9R7bKRkjNwWa6+0eMken08KkP1tFiu7f+zMgwfbpiQ85jC4JZZXg7C8m9GQ
9oLS+6JwNXnzt7zIaydwr4zmPJeUtWDjPQ0SpL3a6W3lS2om56FxOC5Bs7jKB+O/
jSqRcIPgRYtmTsCQrW0sJIHOJMPlD8hmCtgmZgkwiF9tCz6OLrAJyXRA8S9WwHOU
QOxeMle03fvKgJ7khmIIir/jbFUY3WzaoP9pcX2ujaSwRfKwga4joyPndQ9BSCox
nTQqUqaFLhMKTFncC27i7R/GSf+P/kpS0iXTQB35e5NeZVt2S+HN0tYGmDY8DCj6
BvjchNATqUCW/lbwj9AKGjbKLnwAgCNXp1SEKS5v0zvn53uwLhfm+q9Js+qdAZxD
GM0wHN9Vr37bQ/WOTKOukT9llBY/5J8secEuPx0mf7Qdj772H5j3ZX7UVt5BwWq8
SJh7+chdvsLOEZ+yADZdqH1IO4ibG7ZgmrbpWwjrRC+xA1lDGzx4nV58LDrcnMx5
IyLtfSQCT9gNU4B+RvM7jmzSMOG5YlmPS2HfpSFTwxru0p69UxqRJ0MDRQUBUYDq
gDgRXjDgbJXXF1g954dn2FjYB8qhY9QL4LN4DkCatPXUYutCQzkNqnm59iEgdihl
j9akv25R9yatRCPRGIEo5QgNDBEL19+/XEKfESmA7DTunQdtn6jLMsEj6+JWup42
+ivfGX3mneYA9s32CbKC5nWLMDUI9bIuubrNRp2gp2saQQlzg2+KfJH2zxF6E8ms
RFpwVwpj/ArAG3PgXo4e3MGoBrdyn0cBv1FAVgOlbK72nQcQDbTj8EI/IQzgfqkL
gxf1jieZ9BG6ryC7qGSgnWkcxWyqKeyiGpXAM4rpTf5Om/WVtKdW1Qqvkq9UyK5F
fR9MHoDsCFxILqhcQQ5TcOkpQwpDc2DCWcZfX3bfTGyLkI6t8/aNu+xqVnwUDh1q
2RzITRyLXa2yL/CR5OWDFhET+jBURRW70Ax6EIG9TxU293XJKeTJ6/m5dtHLLKtl
FkrFjEZpuZg9qKNTOilQDvNN9nQxC+1HLMyBzRj+gS40EHLjmyaOu4jhvBStzGsN
DM7LKLiya3xc0J0k2xPyn1VQ9xnv0av2PyULv1ahwR6SwCaPxlihJaV3YgbsP63v
ooq/JnWke3bUeSIkfJuq2QpJ+9pEutl2RnOC9WDZi+gWFBT+1ze/JFwChmSYMNWT
+Wb92o2/MXtVwIkVD0mfjzXDT9eQrPW4sfa5HY9atf2KwQTyYHq+SOrVVG0AtqIS
p9Mu+/e/93Eu+37tnT87NlZFjXxs9hBM30EEWzEbgocvml97ISfmj4T56c4PGpEl
rTpfS5GfRGb4OkP/8TdazOM9AXqzF2VI7jVvhkpvjGnIWQZeCZF/b7PHnh83QzhF
RVKKNVJck0FI2byCwIwnSkibkNQS0bpyQ6xazq3QXJUNBfL0K86j43I3VEi8J6Qn
bUkgAhuWlGTOCCsEV9egkTxGGaj3VnZJLylhVC1zWcbtz0I8PygVTJ1/SD2x2drX
UG0oCjKtxYjNp2ayILiw7ygUyJtHlxPWl60UUbeZBLI3y33MS4Hhpe8oHanvZ1UT
RjBSzgm+i+c1uc/OV5H4Kk0fXQ+1w8Pfk5Wr/zvafHH+2rl7zDrL3a5LClAbrcUY
fYnzeCogLQa0JE/bDvTJredRT3yCXXBlbGsmeWX7XzjoXEvONaVNuUENoAArqH2R
jlMVYSMZ/zWa/f0AZOadvXlUgev6N9/Z8Svz/YCKOOTNa5saYWdFExjQNrSOajo6
Oi2uDmrNILp17CT1dkq+lV0bKiTVFhCQF8lvxDZchugvzebAa8o35bmoTSDeG2c+
he6BhZWr/YvBuCN2N15XLxZ/WPc6tPMLki68dpv9Naa6aVE4RWGCNNVL6vZop0oj
609/Q2aVH7LswMvHlZTbk+ZNeeUzMORvgvaqDFY8aW2svVO5cC2098cxHAgPgqqE
/acGPS80z2KDiwYb6/BHGFIxPtUEXfl2GvuQgxi2uQKU1jSxCT8030YIMnWQ+c09
w++/3bzkHQzmYeO0S83Z66gX/Ry6nY/MK49YsWEH1PoFVFDpAd7JSGUNaCo22DY9
Dl8JROz4k47BfZL42LPDwvAUWGBTxxyz/1Eyex4A3WxeAhT2k8XBfpB3aIJ4VBF9
FwVcSr772hnfRuj2AC71nayF34+DG5ogVtCnQrstCroKF/CnrdzcpOh16OmA/tcy
Rt7G35bbt04w69mlPUDxggTqqcaPq6Qx9wfx73DGAgYhoEszPU1zzU8g3TMxqXJL
h95OVbYZPFYSnqBK2PdLuPbqIMbLNfFkKMigWqWZoDVJCgxVqD9MXWdyyWrn288B
2Id5VwiDHngLC/iDK++s4CC0JPWGh6CajOLUzkMwj4NEMAmONJBFHpPa4Gkn8vuX
+upYtIZdAgBa7DescUz40qCDkFT13wlVnVfK7WFmCeZ39/rK5lbMU3Nc5jrdVTzn
7f5rKCoLwwXuLEKcCiIfhqYkNafsKloFp+AABnFAK4F1NXglKWtGo1r5F2iJoo7l
k3AMwYYW893eG7mS/BLZQ3+B/5mOgm8WUmGV4edYDfPfogPwOkhCf6QgoPKIah6l
Z+BsdSppSx5Zd25Zx6spoEinyn59mu4NZpE7S3Ma9zAP9zqP5i3zClfcuqkUU+qw
gfhgEh/OIQbT5qOWi2zzv1aX3xtVoadi2lV/GdnlR0a1TIGnMMA1jlNhqeAwd157
cRzi8gZgK3eKEamPk0larpGpTduPCvGKvwtA0+498Y1HIBZdwwfN4Rh57Xqd0KdO
FtHM310lOUHYlUudfa5GGz5y7Ztymwm4E7VHn+yUcN/qePdktGwuEmK9j6f3vgep
EryxD629OFNGy+IDa4ZFewckq+jgo43xDNl1H1Z4yftWY/J1OHgGRkw0HKxzc2tL
FTh0swzbF2W6R+cCMlVdqugX7emNDyYtpia59Q8V4VlPcqgvSRGAhWCZjF52Pm0y
7ExpzNYCSXnQqenC2k1Jb8Ou9PUlBVz3nxYfmSMIYR/evSq7BwR01eGLgAIdjMkE
tZEMAR8G+gZTpJ6zaWgf0Z8TRqEANRab0mGhsM2dW4UetZabs56R14WzlYyUUo8L
DLdvR59AIJr3bLu2vyElZjcI2a0vossgxe4vFyFukCUhcmhVbLNeog/MUDiRRMzP
mky5GyCMJZxTEVhRaQg3axkf1+J/v50tokmPnB3a3X+rudwuoGgC7HYhop+8vB2s
VXCRR4PL3YOOw0lExEyVV1fiftEXJomeGGpQzVBYKRWMdbcZODLvwqwsY535HSzX
PTbvoPrHCufStkP4M/1Pg7SDBr+Ek07hRBDPIoFg5OdRN/GqrQwNDPlK4WS8Owze
0ojbP1TNMvz5I1pgsZnGn/+rWjvT5V97UZdGDFWBIh2TB3wnuiI1ZCxXJZ+RkK27
tqbwW9lywYkcmufqbDXHI+GEYx2Bk8SVYPiUrT42+AfrVSQLNplyhyptMEGe3bYO
2b+TzxvjBM0c+LXEXNjuFNjT36EGNbscOE0YrEVUOjvYi2/2TWGNF5WR8+A/1t5f
ODPXFMJ5uJn6L6nyEDVi7PaHk8pq+CGKlzGZSeLDr6+187tAsnkMAbowAxZNwUQo
m9WxViX2MQmVMZraIUgh3xO5JbtZOAkRw47dJ7mshdhEiwdQ+S1EWDvsVYzbl9un
AOkwUM7GcIJQBqzQx/CJFZgVGK8uEQZcLV86D2JctUj5R37pwO899B3QkC8gZnDa
6tLsrvwrX4LYusb5MpV11J1BqhOfLpingJeInHis4QoFDMs+Dm5NAciNIr0LMHjI
VIPUFK5rCRGX3Fo2bV3WGx1h/NApOlAXxOYNYRQ5hfrfmgBHljNveDAZ6Er8Mb5x
UGQ2XLYG6ay3aFwE+XLU/Q5pj4vLjZSTR3Ts9sV36ihVX1HLcvMy/B7KEnUcHjNV
kMFl2LF4ZJc9dXERqN3o90LHwcOSG8DZZ0SKeppyITBt3tcSIjDNn2wjxnLaxGnx
0tnDbkDqlm/Y/i5SDRlXX9yYUnQQ5f1lmQKaOfyZKcvfItlT3O5YNB3Ob97frkln
/vBlZyMoA7HDqfk95QBn/hcABG7/2jCdRAXAPTWSXYix0Ut/kyL+yOHXPy6Qdzfu
T42mz5U7q7DxF7OoxMmGYMPGTYfvt9zmdrGnOZaDQg77ltiFSetQ61JBIAvhzlCM
q3WZTPlfqzWv2YgD/O9Ov8ADj9fr5enRv9GkdRN0WItABfmVRPQ3aNROtA/sdMNB
hEd/GuiDvN0mmXTA4RU5WQC4qGo2TM9qqnBlO2/U/sVBnbGfVhkYss0NHfYMiWW5
xG4HE7ox5fsH9koAbcCWvibJQSEoIhp5iaT+p0ZDQluqFF5hdGgNVX+HsGihEY/W
Zy+Ke1d5Z8IvHhibAWsgk9youTo59TKjY7Uby2+U2/9E+TBwdFOM573kGrXXEDHl
yUH2g7kNd6o3F4CeAC+HUzGLDTWddxSSp9rh9ExrN6xmyJoiS9h6yRT03dy7GD/G
KR0eiHovyZ9zu/2Fo9CJEEOUCXr2ZBDCda/qlAsqfimXRY05YzPUzBhEv02I3YrV
Lw1v6DZpKUL9jS1OAwctWh0rsJIPkD4ePzc0EBujpec95ygBJ6XDvvuRIsK+2iFD
Rhsw+S6vVmaVcRnCiKt8T2feboKKjj3UWDaug8BwRvVMuEoa5lcBSnZ/qZPUUa6C
fOj47QoGKByuIluhT+AxsLxkrrEye7UvMsbTdz3Yoft34RvhJMgTqP9esP4gH+v/
SekgAdk9VQ364KvYSLCPmn2EItzsslo0+52WllLLZHKiqLsYJ6pN1NGVop5PVPDZ
6IsC1uegKeE0kX5czhYBwBGOM1uqz8M+ZB2u5qTtcAUt9oG/JPJqhLib/xvYe8LU
BP+rLE08tXaqWEMS2SJ56IvjW2MqYd/Y3AphOYuw9aYKUPHqmhStc7cX+32Ox7rQ
ROwF5GZXM53LKp6P24/kgvq+Fhojc1EpzVp5x8o83tvZvH3SyJgM2LfwxuGazwCo
58FYZK6xcFpH/SqxObpw7qp2uklNhvfF0r0lYKeQQi1Ea0ew3cmwLML45LheAFnF
VZIp2r28GGGwsCKMCcVzWGBC6UayojmIb4ELWZFEES3dJ7G3fP/+g3nSlSDA3mAy
ATZe4V/EG7YNq+2Fx5b1lLqwmDjctgScb2WWO/XRJW5z2v/AG5Ao1fBVSEoWiUac
vtXU0NIXdaGFd/PMNW5IwGg79Lg5o2hGzmMHmX5k0q2Np2YRAzFgg/i251Zbc+ra
CyJFUkcnqkRQ5Objh+z02RhlS2911NEjKm2Ue/kkJAfDvgE9EoOZlP6s5FVmeosf
b0pSRk+I4rvhwdvat04CfnncscwwzUMDmk0c54gjv2K24ZlylWkwluiU2BhqABwN
FJpectoaCAUnFAkKxbD2cQLAabWZZk5WyUinyPS81kirYb4ML5nzHCEH2Kw6u2WH
KHEdK8g9fYAxjNJ51X7jSI3mrP+Ysx8soedBUZVcNGN+Jrf4xKQO6U4U4Ib8YG3d
yrRE9jP4On3ZkQs+qK6b9Ft1GWOu7UBX/rqfdapzq7DGQTWhwYz0DGDoNlHA+v/J
FyQcq0vNmMhJIozBeA3uPgpVYBU5zfKCQeW3AMSmydAxpNbB6qmY/KD5s4k9T+pj
RkPLkVXhkUyoagCwV+kZdqWj2fVJMFtkMxqKHlHrZ7pC3eTcO4EIC7v0zANtlgPX
TCiwiI3LTVDYs8q+qOsxqbtrbQt8uPZ3QVHSk+Aen+V1L9L2lIiwLAZ0QOXef6t+
pfTcCHsioPpuMAsifWZNUDIOl4c9kHgRjOtB3Tlz+2HCAHSVgCZ3eJYJfsPMdIV7
cpYmh8HJQZOcX5bTzud4EgoEMkL1TgPnD2w7qNP1g+ng6vBcwiZBInSdLwt1H/zn
Gicuv2tUutcLBGeZjbvOxHfnHr9uo/1qaLVybxQBbnOm59JjqFJTcC82B8+FIPyH
21qvpHSyxxAh+gEoPasa3uVdb6eHMcZGiFS9rzXH6PFYjJsFsVqw6gF5UZMj2hT3
LWFCnc6xSr/xy2QgJoZr+9aw38uE8N/f5U0CknBhqgP5rJc/oaw+9wNjsM+/but2
Wz+7r98kFDBtW85yjXmzGBb0PvWgRy5W7hLE55+kmXHuZoa4xJudyexYG/UETIyz
dFiAqljwt5HGUv8Ep1PypQssGAiDnWHH8BjpYIuk5F1UKXlntyaAKRIioe5f9szJ
5PHwdUS6/lQv1v8nq4Zy5xi8Fz7eYU8TO2j5ewXRQNH+VbYpIEdHldww1XBTXsKv
UR18J+p4972j9Kl+htM4q4hBd3aQxusjz5YrAH/baT89ZynyBFvnaIxKzKTO3S06
T3n81AQw6PiGbuI3nI/FNjbTLQVC7WSW0YRi7pkNc8Z/Wyub8r4BC2njRFQbNydd
NcJYBtEtzJddQJdDUtKfaH9CkhH4LyQ2N5A9FbDPEM9LAnr5jPuajo5r8aEtHY4O
ZZ1v6g8xOgparCJApa77UResdw3J1iSphjQwyW15JZ4n8iPHsEsrNZY3jkFgm+Iw
5Uq6VJ2BsbUA1tNI4LSrXYRFQcicZdfiCb6jKJEBsXEEOygFwWS2gQbehOIOIdw4
`protect END_PROTECTED
