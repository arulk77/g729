`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mCDnWIcVhICwjHB+c4faLL+Ibr15uW0w30lEcsJDKJZHnI0FNa/1wSnVvpQSuC1m
ifKvpvuhyT7zrc91DxUJOWivyLJ/cUk+2YtoFKOW05aS1BwEt92JrACVYON+cVUu
c1apmj+0r6AvQ+gZCQ4A09vqtbcdG6PAxWNAAfmyr5fGdVHsWcnlY3E4f1ycF2Zo
Tkk8AP2dtIhJbbMv/oKSkVPpbPqW1f22ehz67Ug2VPKcRZBWB49HYhlUaU7JYzIX
i71bfOpje+OONGAdaz94cD2pwCUDHe/bpqzLdmFg3xA0I4FHkHfyLYztdeA3MeNv
3BKV7d9e53iP1jGVMz6rlaIQof8VCw2AiX0ZP4solMM=
`protect END_PROTECTED
