`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveO1ic5FGaLENZKfvAP/Kz2iKo53OQgw3M6E4PIyqaJut
4RbFr+2yS+o1FvgfExaA0ktiReKbis4tZip6pwS9tt+Gk4OdM+aLYmY/FZFxZDxO
LzExB2uN9o2HlkgUmN1sARDR/BMXiT2W/mf2fANMO0T8BrZjc8mZpUfL1R5hpkMD
iehKPJ3hjiQlepe95ZAgyufJbHV8l6Nvm/LfXKI55E9XJdsh7/cIPj4Xc3hBaNW6
`protect END_PROTECTED
