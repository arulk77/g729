`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
adUeznlRy3CxlnF7PqxVEz8O63epPTXptOGo4T88a0CPAXZZVw6wUuBI04GKNUdv
sMf0IXVMFLsmhIWWLlKC36prftZfXUY5GU0OD7yg3zZbTcdwXMokJaOEYxR6Vt7U
yo2D6Wm641nzKttFsDy0Gzez4mukxTlWhnukSf488/LhkUce984cKBoQv9YgYGZM
ycwgWzcNrc06ZL4nhNhKextvgUrDeNUEGFG0TBbtmUXg2QeCjm0mx4iLK9Y6s+VN
uPDgvsjJkpjxcwBT10gw/XkadObSFHxWZoAw06Q/d5P0abbLbFyzbF6ySnH7tb0y
hhnRX/H+BuDKXEuijBTq4tfzuUNkNBcQs+cdAX0vV5M=
`protect END_PROTECTED
