`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHLOq4dz9RmQjQdqMv9HpatbcAc4o234k3fkQZQwwYMk
TWBvo390NZtoN73NVR8lvyaxr/FlkBo67eyi9J+qEiGEB+fPnl82OgROEkirjWaj
q5F3rZd4PMWxmQqUTdCPfLGiHY8S5UgGWQB9/HtlKKbg0CZjOr7pbMGO310ONNTX
p8qJZxaH8IPParJsZ+l1igtVFyiF1NkcTPJ2Xnf4zKWTmqeg0ZWMVbea9fXTQMFD
v4WFMWA71Yat+I0tEFrQ+wR5Wiosb3uWVZFCHdOe4F2G9TxjPyY+8q6VBg23AqOC
14/PMLBCnAQnH1dXKZFUUlRJVEIXYkJW9vOPSK+rhYkscbmkJ2HzGfKSeVBhXI/F
QWQsMNp104/NYrOXhWjLqjJwZRdQlDhTauKF3SWEQlyYx7U0xMlqLgxCq9ycCTaT
z98ctzS+1J3N5kZtRybRs4E0U1pNgfGKEtN8vj0P2yu8u8am9n/JSp0COAXJlU3Y
H8ZIc8hiGKoymt7BFtj/xUdaaVDQ4jy0wGqY522OlfoPdKrAQ5ju2RNqNuXw+x2F
eKFmud5HGsifYyGn7kGMBOGfrLaJ6fl6TUJI0FkS49+oIrH5OcX761GElZAFXRIA
j2iOz1RmaXDxAog4ASnRuolzKWxUrkK6eUoexQ2ZP8gD5mH7o19B9ybHO006g07O
vlWgPPW0DrxlU7JHihmrkjGuqjvmKKgNgdwXilcKSPBeXhiMCCFSAG8KO8sLMUaZ
5aEhFtaB0BcTlMskPA6Ey20+jcF9JUTvr1r6231+vVQLi6kGMPOh+mvvQqMamrlY
BwKk3/tB8gFID3nfohlLIwxZ3quH2EEI7PoGz6G3QD4=
`protect END_PROTECTED
