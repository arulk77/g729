`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePOndvP05hUgkFVaawP+IoZI0EkiUIbDEh/qNt3lTdm+
8MWL7NuG0H6cuF3GSzpEpie3a+3zTdrELAxP1ypcARV90IGBiF/3HJMwh0m+CdTI
txm6K5ldI5BVW9AK/5IYFdQu4uLTrtZZ/lJqHP2lEYBi8OmvjPJLh/1uAcO1zTYK
g/xG1jsqqVG5GW0BwKmnyKrjRZSIxUu4vdrK/xlWEUZAwr7c4UbeRLXZAPfai9Ym
`protect END_PROTECTED
