`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
A1/S5Y9ZsMsv8F6rmZwNLIWlZTnyJec0l/1RboX9DBGypjv9oJgqAYKt8NIexgTU
tC+k3ESbXJBEWw43mzR9OAtHvtLNO0AKE2RAULzwyGuxeI8O+V/mCJRidWmKhEVm
jMH3Wz1Dww3jCJ+cnxJv4T6AJh9Gq+hnmjdjX4ErbGpvkDd5tVrhiDeqkJUip0+h
PMz7i1RJLlQk4N/4gbWrBfuAn9gjfqpvWUaNojlAM7wmEMIJ/u2m5caAsmWSbjCZ
i5HETsDuoXqsv4vQLTwoOalrkiO/SnQP0Y8yP4zDwX/4Gs8J0Vn2qde88aT67XA2
7qUIXUrwg8xOsciUJWuHyNMo0ajU15aSRXhqtVQzfWw5o0R5XNNVreCz3peT77VI
w8413hbpBXZa1XpqJncseDfzwZdLEldGWUJR7N6e3MpPAXgVMT+IcxctyW4kMtKK
n+JGruZBeewmnjpP+PrpEMiKsokb2+kwGab7BzCsdZQN/Q836rP7rqAaVBw/UuBb
2L8dNQcKRR1RpMS898gKJ8MnFai5QlkF2cVBqeiZIthFLlJ9sxgLdFQyNbW1wjFR
sZDB7fTlV94+RLZM371NMFtsCmqudaZDJ1Z3XBdVdOUZnvcF4yQcME+nN/c7SBmx
uuMceTA7jJq+w/hWQvoGm/kF7dlgxw1fAQcRrUyYXXgWO/Sk9uF07O4TM5eDYHp7
G9pwmoJfW6JcOjkfVbvmeA==
`protect END_PROTECTED
