`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C1dfV0tHrnnghlTEtZ8J9cITkrJ/xR5yZ+mafvSAm3mT
KU2m2rkDygbcrt4oBGhnJ0+09wEq6pQNiD0nreafP5sYAJgZ0FRIcDNXw1PUg+TL
ONXpLlf55bDavX5ichggwaMdHCV89CSmsRZyPxJpr9SmibKhLwnk1DFv0YsKL+WV
eV1LgtyL1YGc3h0038rFujixPrZgY1u6qmJEVzUXEx0teknuhSBNJVy2aqieRsmw
z2el+FFvHMVjp3Qy1SuIa9RwPGKvNxi06fwVsAoTxD/WccOi4QhsBnWfUyKisuuQ
U5UEkmTILxclfyQbYCPkrH6Ga8v96EySzw57Pw06U8EXnCf9aorp7pJr0eXIkHLP
/DIRRKcu4a+wBg3n/1pDobL2fVG4dKyJLL9JWG8n6WnzzPUhqmRB5cNwZRa2Fl/i
gyNihJituZwD02XO1U11CGukohfwWajGILARBFTVMp0GXuUIZeGw+cU18hP7kTrm
DK11JxQWwgkU5iBkT1ZfyP78ln9Es0MT/ulk9MdIZWcu4cZZCSZRaCiWb0b6H4IY
Dl5gFMHtWuGtsvCV3TmH8ZT7javmT+LceT0DDIDKXbpjlKnYini1UJyDz5PAEIL2
+nm/XfW9t0e855pKx/rJR4H3VtYXuos7tzWr99xw7qwqS93G7vgGQ5EX5BVRzFcu
vEQ6Id7ytc0wwS6IRa+bSopNnlLDdmYe9FQRf1s5plyVEDsV79QtHsbJqv3HFn7Y
uAgy559SoSRJES+m1jcU918Stv1NCGdYhXMjCdsw+aqyQtPamJbZu7lYfomkHN/k
exGN/TRw/IOF7kG9eBFWOmTOuKUVhiQ1IKXHOKJy57a2QVREEeGr2INI/eG9i6fs
TkjPBQU+pSGfbnZaEuOcpt3iRRyWZgmwagRIHOYINfz9Fz/xlTuaPKZFKMbqv/IC
x5I5OLAQaP4tgAx1/2Yzr6o9/RgU+Orjf+dy1vWbOJg3j3uxilkaL5Ie9gQWN+Ny
zDGgFNfxLDZOA4WVjKNyjeK7OgN05p+vKPofFQPLLJ522GTC46NzAkZiszty+goO
7oUFXvzZqFhiMF/adMG8Wj1ypC/gRcCyJGxTg3sh63jZuzDon74wy2Cuo7T6dA0t
acjhRNdWyuAms4mmDGqgqzWVsGwnbojqUn8cEDXc8uIo0iOXggIjz4LZMToVshKs
yYWh0HcR6AnLomdli8CfJGX7QNe8PC3ntq49ZKLxdZ4nzZ8guFq0raZfLigcLD6y
Bj3+dy1pV4lN1kkkv02/R60+yA1v0AojBG9zW2ABac9TLW2ZYh7HV0t5piiIrtvE
lVj4/bkJxdWF0Zg/rQD0jllrgVqnW4QvNFAaTJN/pOGsURVHai77A50CyDjkZTS3
I/SfKIzssj1xq4zznXnRb4YwoS3hjmxxzNAhWrQyb4g=
`protect END_PROTECTED
