`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xMJQkt68bTRDxHrYfJOwxJw2YyQvOG/rJz6C//noGzE
YnNDod3SpzLBwkUdQXfjmpZ+M+NVz9VuvCaSnz20iEQQQni56Vcu++YPzx53T906
/1O5Wkx6Wz9vC4qYUDVGAhz6/MQ2m3Jhx+0D4V4eQPq7yuIQBwMFzbaSCikoenFq
MKgJTSDmeIcwuE/Q08/pRZ2wLl7W2CY5IRoUA6TLdhlUEFIyN89RMJLWrkQsExzd
OhMxeWfaVqlbG6KlUB/bxbQtJ9JXE1HZHCBAj1DM4mpwdesgVF3LC7rTm3gVSDGi
xR79mQneDduJYxsQh5ixTjXUqdnt0uWHxon/PxCpzmDUYjPvmTfhhxbfVL9bl+09
DvlboTQAbrngN5oLAZygwocZ4KBkhxzj13zThwxp4GQA8QR1BFCn/4OUFtclr4ez
6Or+0Zthv5XHJTIgmZdljfsighrurkftQ3fB8fgChuoDYG13gr/0m1rAxY9S2YSc
fKIFtAPhVOCDHvp+SlTIl4u5+MBUFZkERtMyI4qH+iUXtEZ4C0FGbVvyg8ZMvG//
ccroCewFAjaNnk/sw79idN+MztXYIUc3S6CuHsYnga/RNMX9GzRauxuRxcNjgqgf
21+IODVglM9Az6MwnSiR8xnYmKrLuiYCy+kNLNIqxV6BZd1/ODt45IUuvEzIcE0V
Zu1Fz5Zsrg2mJUMU7mszZqt+LijkJ65cwJX1s7VJcy5esWPoEzxysSvvwit70uJw
C4M1xE7rE2bf+zd0v12wNR8x25lyt6bMWYDOkO8FfyBkavKkP+ZKgLM1KWCh1E9E
M/WSgJcADEpSBeoEerk0i5iFmliO3ZE9RO6XRZPEhaJwRbL8cWx9aU+ndI/mCc+3
x5J2MFM3dTzBjyghEOA7569hhHenNgntd9f6j9AxmrBDsgBWtth5hWhclCl1+dFs
nQRA8cuHQylnUavFROT6fn+qEm0NWxzV4pel30vA6PArAzvdclyT/iUEeDoo4B1Q
cQUoEAfKqSGUkjMoKkrWj7SZsBrlz8Log+fWsRoYkr3TikLrGJFUyoryQh0IUuv3
y18l01EGqrsuFRHzTVFC/p/90w5539Gl2GF5OmEExQohrMc5NrB6JtWF9p6qN30q
KFKWezdoToSFV5vN3K3OmvqdjxEtJOhm5U9xxAos8uDG/tJU6e2v5eryO5fL2Bu1
w2tuS0vZQFZU59go7ij35IFbrX8isnYUjppgIkkFrnZ+PqKK1ZdSQujFluVBT/mG
KKODkSUiCW45O1xZbBmJNVjtOGugTV+3sZEQvCBbtazS1f9iJVuCX6ZeoiOsfjjd
8bwacs3X0RfmWgzCY1J83Rtwcps8XFEt2VFG9hJE5e5wKQmbe4/cG7YgeiKYDdMl
7LTpElh3b9e2VgzHWqTPm72kT085Ww/9yYfvxFSNAqCdaZote55KSOOxV9NdkXCQ
voswInvanSsx2IcEUmUZFTO46FJJ/QEBbdWabRL4ZV8KFF1Csp7Uw/4aCUyvHc3v
rWUDX3Q884LnbxiZSG8gusKQmBz6oPVgz7t6EXBlE6NwWP+q3yAMRAnjw2HZi53E
8Dem7ciYtp3TZFbr3xdmtQ/A4dvWKdzZv8m0UEmmcrmPeVzjl7hc9FLiQIChFaFo
UFgM+r+kBk2qLde2iUgpSBfK5uBLMF3yx55tC5b6Y1a4yFUzA7ec03oJkF04L22N
GHnu1sVcKqUj6LG+mycSjXAMTOwjUfMgYrc8pBBKdocno6RXJ8vusDax77QY7kTc
xplIkxbUZ2NYhmVlMFxIXMe5H17rILb2YICD/fYdO5+E0i5Drl0/z5q7AV8PBWEc
v2e3YGyAw9mSm1+1ojVeL7RgzCQ+fzIBeFBdsbMPNC3zaq7TaAePAq82BIaHlHNJ
wkpVYN7Z6iBsVF0te4nTsNAnCW4op6czyS6LwFUOArBUN85JCkixQVyWCQdppRtk
ocWAUnsnF6fUCeVyuuw/aeVTNrSqJ9fZDrAyg26ltGZL6idq9DnWIpcHUpVJhYey
8PomAmEDHKlUefEYsySzCTONiisrWQbZh1wRoBZZElkDGhmDhA3co+y61v5kF2wX
ZvJMW0z1VWHwdVB61b0/NnCzrOfIKXKo8mQwgCTILcA=
`protect END_PROTECTED
