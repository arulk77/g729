`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
7RWERbz/SCu29vx1yp3KREDbsy+We8lfDOE2Bcpt5dhZ7V+7EnWPv3YUPYz7wE1R
VfNecQbxn2NW+q6xBQs+Ety3CYKH2rkOUjplJTwraHIXMVPmsQRzT1qlmApE8U3T
Su/QmORWkbGzgeM1qKquYj1PCLLB5GmIwtq7KKhj9mWrTsd2qHAb1AkvrUtWXDjd
`protect END_PROTECTED
