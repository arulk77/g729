`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveICBeCDO+RCmCpu3ZFjKG7y/nyKNRdy8LNrc2SnBW8S7
LxepetJJvlU7G+6vKL4qsFRPlTLCBsHzt+5oI/3WywAp4cOb/4SneVoxIHSaJDBT
RCXbojYCa88pBLiNE4BzIytZPOjDt+BnuGo9HyuMetozb/sP5y9O80B70v32ESZE
LerIiP9d8FhfGPy8/PGB+g==
`protect END_PROTECTED
