`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
nm3Xlzn9zUn4PtKhF86EKMT0NOgqrRhSMouGvhD9K2X3W99yhb+vMBpZHUi7K4sO
xNP3tHQv+RdD56YfUZBDH73xwdP/QpPVeWOxZGiEH5f4II7NwvDuepVa7KAVpvoL
HJR3oNZS8fJVcQsRAlbd77hAW2XeEtl9pJSUBn2JCssDtWOczubhaow2uIoDuJy4
EutFNbxwqyY2IJ6pdbvrfWpTNO3Xy7TBTEnUSyDadJs4k1tnQ+Y9MUN0jn7Oc3D7
M2kDhsmROFufRQECcsc409m+oU6V3YqVQb7t29uGAKpBZc78XUmMq7tA8OCKEvNX
ocWdPAOsVZdij0h+XVhSlibU0YceqiK6BnUHLw8MlQSfoOtlJgs3OfIdHMDiNcci
V3osZ5Mxm0D65gPo5l76VumL1FCA9PXw81GfmeRQ2HRmgQh6p60+XkPOXLfwDjP3
qFyp0eDbmJVd8HkTRwFTwgPkJ37r9YSM+kC68RcHUzv7pxKTjLwC5HZFKGsAglGm
WFjdm2i+tp1DANUOGpjxHuCNg4i8uIlPPLxnf+gy76LpkM08+PYXtl6cXfZTjNEO
krZL28u1mf6nGpWujC/etcpKBdZ1Z7ImMNyUq8HqcLmT4SkCt2hYWY5rI/aeVDn0
QnL+HfWao2Xqn2iqV+cyfJfxmXL5wb+VCEOcmm/KFVZOvlb2fOqoi88Dw7nAHU+d
8E7EMZ7ZsTp+V/FDDGOriJuyg4kQ5pIgwv8AGZjuftVLBs2GULh8TC+yeobfiRhf
`protect END_PROTECTED
