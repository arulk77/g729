`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42q3n4YfWB39ytlIUt8m0d2WDmxpBLh/iuyAnYXHUIie
JTRov+hZ+Uo8yDusNZc7mN6oSadTcgarO6fyJvxVDwhRdNwM3b1ywjBjDz+wxXCC
zjmxV2mm+YSoSwf6j/1COZkuVx9G0DB6ebZTtge1Ewz3QAKU1FrEsVGR2edo0BgK
c2GcxatQg8Pprm5PF3bsz/HrJmt5H5lpbur4nMfDLx07YPzQ9cHtnCydonXFYrk0
J79OBK5/JHJ7wgIqnfGqbe58ik0o+DwIYzG13AKkU3YE9j17a5v8sewkozibKNZs
p8DFhMgpo49EL3DlzdJ7HAha4++nqk9TL/TGsK7MEFIur8wk5yHSh7engiYcJgE3
VpQ+UBJjemiGJqCyt3drYg==
`protect END_PROTECTED
