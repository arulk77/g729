`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN2c70kzG5Pcqowoz/cgAIfPfw41qec8s6np6Zhi0eJbn
UWQLFQzaOMxolO2tcQCOxNj6/m1eYLNpnrDX5bajfEvH9nH2fVEd/urq6j3AyK1r
jIJUxgEnibCTYnxRxcTH1W1ayXMJwQsxI8PuZ+Cfbi5PEA5fsxVwb1rhRy58qxpj
A1pu6jJRG+gJn2ROvop/Lr0xIOIet4tXAHW5kuMHQP4lBAAhkrcIW4uA9sG8I1px
if+BK8viUybnOMcK+YHy+r5nknKTwL957fIEHZn8HdYtGY+Y/ZOZV1UJqW5iu6TS
2/ZDslZ+j0Xb9m//JJ5lmb8er+iM3UC5Ms74XNhMUTP3d4TD+n+rgm01YX+Mzr4a
M2ZfEqS+glKFa12G9elI/T8iidpJxHnQ9CrPUlQz5m22qeKS6t92x4WxacTu7yDH
gyJ9yXD2SA2oLSkOZj6K9GPVRiCZ9F97Qcd/MLvvFlBpvUv9YcvPHqaz6zZXwaQx
qRz3PSh3Y2RhGpGRPH6WgxsK7Sf31v686rdkxrDsiMCENU2uPya4J0H7hf9nczQw
c0xTD5+bFALAhzrzrwxt8ICuq6UGCiIpwvHnt7GJgbVDT5Mm3wiz4IUSpimgtAnO
jWMSlSOwB3lj7B7/YQ4HPQMtIV5fQ1qUf7o3Xr4zIsxkTmMnt7rI9D+GO/v5Zg6H
cnoqqfgldwF4oxJcDVvE3lb4jMyIs2ymVvAPedHOegOy2Vd8tLq6qhAl10JzQAn9
gvYMbA5ryD7VfLuHWFAOC/ZTA7leSkl61xDPHKljJn1C+s5Y06umsqxSftMV+WM4
HDUAiBc5EU31QwZbyYPNYAmLm3SQKeAbFyJPf287q0fh96k5oc5/mXCH4+NME2Mi
CRymkQ/tplPtJg/dvW3I320J14mudVcHZsvcaFQVbjo+F+Up3V1IwLsQuwbb14On
xuYtsMXWnbyvOSvLcn8B4WPcl77lRwsmn0LnqwwGBzMI/S5rciGk3CzWKswJug5q
uP0lD8Xrbj0q2wCoC6y7VJqnjLKWkSKV5iCl/bADee5DZ86jLT+w0Cjc6K2ifPnf
3Eu9Qt+yFIaGrQ5XTqvXS6FR2NhG+oEiD0DlBPfUFJByDGZTZpzz183Yp5nLafvf
qZyHpNq32PB6eNVMuK4yP7URS1cvR+hGI+nIrlIHoQFjRoiDJCelv4QyWlKPPFO0
V8DSSqbzCf9n9u5GpLfijstYrpNjCt6a5/bJgWg+fp/jjCTkcZZsyIgRZhqkeQOF
keO5zis/ZJRDIjKWeVlmBkqmwHFsCGWnPez81nqEM6JNPbv1Ch8aU9q7FPppt5gQ
gWix/FJaTESn+8WHeQaJahLDNvUkADYO9naLPIZzMhCiL1WHKwEjDiQKzeIojFwE
CtWGtnRxTS38/Y2KttviDKMIW0lPPogL6ulIpi1PiC/Q7YIPF6ohnVfUCgSFHy7n
LJDsbljoOtTCDqgpjne9b0PhPvv330q8k6/ci0z112gwL5VCvEy5MROcK+VRoEMn
XqbvjjhjG5Ne7k6ncJY6BnvxiPKZeQh9L4RT0y+o4mJrVMLwLdr1jvJQGi3/U/cd
r9rvplsWEaT4rlmnDwD4VQAoyCi7NyCN6fX5/SNINMY+RqOJNA1oqO8q8Yqoj3aR
k1pnWSzm947ZZnvWcaCRQpVFJag9rms391R5A+kccqlgyLC/UN363YCzYyPptkKW
C08Xgj1O3fcClyWuWP2jxtsjqhWIFJrBwiuhp7G4DrWopYNZZ8CKFY70rfbeTgfU
5rV0GRf0XtZej8Z2F71paPBp54x8ZFwLPECv31T6w18z1jPoLGAf6CDoDbSGDxee
hQ7rqMpduVywk39V0xJI1owquDK7qQA3isIW6wzPrvQoQrT4Idz/+LrYRhUxQO8I
VMKFj7wj4+wElb3UgebHw+xLIFOUU4uHv0kA/jm1280hN86Z0ZytE+Xv0K/T5qok
FG04BpV2FfJTKiBlk1KsvbI6CtU/5DTotjzjAdeSDeFx2a3J0UZ9r8l+YiH++WlZ
/suOarinV2gsy4AzHYDUOSuQqAUeBTwxDrrVTU5IgJXFChkS4SjHXzx6NOkPEBE2
h6z7VEzmOKxBSp1DSuSZHxgNxfzlZUoGBvtJenkeBUtzvmbKebotTb1JttCvo+IM
B4XW20a+33fvgzBJMpwPwcb24S1iM0NPs3sExM8jo7s5EKDIfk2R+SJW6HsR5wrw
eyJI+dGaBd/nnHZuaOYhVDbo0lDnPj/SaTIL1AAY4Ly4woPpJK4qbPXNXGrJGD0J
1yhlRsRp/bfCW5Pn+gNy/9CXj4UvOYynjZsoMoWT6WvtRNOe5rGMEhjL2xR1ycgy
/J939glpVx5ToQor2slaF/+U6toJLY/JaZAmPa0RuKgaAklCF/VNx5K+SxZI48g+
QLaDAdnDWySbHgbFSNm+8s9O6ZdCSgE8n0vH5C2nYGlc21UOoe8NY7aQIS7k4aiv
YxAWRgOZdPJLPe5Vzs1JbecwQWI6frBZZB9BhAgN3LOxPqvV2h0AaPxEvGSHyDmx
JkiTLzabhuBZe4LbDlJFjcOyjVOgyjUpFkGfom+oZmGmOtGe1CaMxm1Ky7IFITyc
Ycag3L2fDkCR6hB+yBaia0bo+kNkZXGEepJ4k0n+NrjuQ4eSFuUR72FlRgJrGNdb
o+fGemfPeCezSxBruM78FfAWM0Ierdpvmm7ZWe409MfqrEtncDoJC90iSRvkhQ9W
q6mjb6JfH9YI+vIOzYLfEFWuf+9fZiQIHR5CuqXxLJESPOAPN+o0Cj5MCpTZeIyy
Yfy8srcIR3+Wzti7hSNmbsk9X0ZMCJwhnGACL9LXvVV9gL8RqhL6N6ORjMJEYKTC
nf9oKfTdOCw8+jQg4OQ5lN1y5xupVykvw7LMMUxL/9AciG+ZeCiOHO3WSEkkDOeC
568OqqTKBLhyo8rXQMV2R2H5saldAqW77bBDz578RPuV9GwRWq4RwVW257Trbntq
+6MHXF40hGFn/NPFECeO1MdB+AEQTBgMZ3Yt6YZIbgCUVsZ6bJdl6rbwCGY/E+82
/2B1aqHx6/TWUBBxci4gpcZMLa+/CEa/vDMoFTLxbUok8uT4kiIHvoR3GRhUiUKV
3GrjFCzouMo0x9uV4S6MbbvcdaJYTrU9YDEDONbW6AFuq+DUWfk0QoCvk7N+Pzw3
imF5ZK72XvZc6tzoCVczyMvJCpx0Tdrduhry5EN/fuxP63ABEAh4Ppho0A3IktVf
w5DDYzbPX8uLkoyjvYu61z9uKYOrIp4l3yFuK/zS31RbVr9ixpv6AEduCPLGw/W1
hEz0IrtRnhVpGWsRbr7teJKZx1euRf0dNLlsmu4PLselpBmwfpmLxW2FCdedhBnS
hTjj2srk5UA9j4u8MFRyxcDtr7noQ+En3oZDvYY6x7Y6whhNgKasQP49U/93QQHT
TGudEEzdK5epruUXvIhRhdCsfWRfJM9JVorYs3GGraADJz+vjvXBK79MFgOut6bf
1sPCuizCALTR/0q+gNDFWeSOypzZb/rMWnT7F/KLg7F+0ecRww0SKdexd1pRCfAK
WsVZrfbGI3Ozs8ta6AY3Jf+dyT2bGlQzCSRyGzJCooxRJhJHYYnsAuEks5WLDG1f
qTkHq5B44rzfMeBfDQWE9Bitr29vmxO+a2d9N3uht6/IjM4pd/1P/KsvLbjkIwor
cKr3YLBF9Y0b54KfzKbJEGkfQBrZi6r6PM3C31GNTzsJe8Ohfg8zowBBzfRflGxQ
c2bGnh3UlcOqzIXcrxYZr7mvGO7KArN9VoNqu0teRmyT8yUnHK3MWA7M94t0gv1v
EP5SKLC/OK0w5WvrcC3hWsBDA1WQVJUMVKJxBgVBHuOnfdRQfPoaqY1C+wz939Hp
slTfIYP/cEVEhtILehuqzb843XVp6TJ3PhZvRq3vuh9FfwB4g2Zws/ikIor9lTdB
f3PZYg9umVRNPHNly29F31hed7zoH/MrymfoJp6i1zOTj8GcjnPa7rM4ZYldeDBX
jfJS2I0yrUqSWMEEk1gWNcXxTPMoXoKofn8bzdZURK/05oomDlpGu9flrpsscsnB
OJ9vWMabupXsPCEkVmiHcEVW7lJ1TvWIU/S15AFUTgiWP1Y01KwOyr1G7x8BlgPj
V1j9Xrcj/kpQGciawfP4lrBEoTIqVT0Qn2GSJRFUkIQ2tn9kp/oCGRxohsiLNe2q
yKGmGM7jzm4VQ1v/xKfU98mL5BCBagYtZ/VGKPNcomfGMFvCYeprLqzrsB3TSffb
M1fkYiN/qUl0ifWUK/0Dz6fNd4+y2w6rBcAJ3k6Ufiq8ff6uB7hhD4GjWUkdRLfh
wTOCEuE8qTWuwUxM5+oJUUpr2MIhVNvyLHLY9mXGqBHYhZjqlF8v789lUebw9IQv
u0hZHOfOHwVV7VhfGqv4H1LXMRsfbmL494bokzZP4qXOCz5TJBisBXHAWlHZ8rvM
2oMrH6+FUenVe/1R9LoS/paoUBs8OQzajFmpGy6KlKjqLlCc0tHykUatnZCTnjqZ
chrv+SqZAdeI7iOuHu6PP7dfyJcRCN4LOXnn0KWPwsMYD6I+G9WIg6y/C+4i5gMa
ibE0byWEuhjTBj3NqOAFaiSeAQqX5jmVsCvLi3b8Nmo5QpuQWadu6jibPjoDEMA8
5XOm5SVsH51emRKKiRTbyDSDYE0X9DFkdijIO2YfCO3oW8Aaw4iOBOiju41ZALPh
o9Ivhz2okl1KGuDhbTXWgj9u1goPgySTVSZyFhoAHAaIXjJQCtFaBCBANGSw6TZl
mUxg0gaPkJJveaYtM1NZPyPzaOwGuzUb1P0E64XkoFfd6fDOZ6pF27OxS8eF4Ncx
uuzD0itpwfIST28OjzJ6mSkTBLmp/dKdNvEqxQpnFdZSpHoPUtVBj85Z2z8kb37I
7y8gp0suomDR2TTARYYOaGWzL7ImxmXOVSSY4t7Nyxlqi6LjXS4MBvSCRhsgln9V
B+2bXBk+Aw3LJIwBCS4H6Y5fgZPqfmS148wNWB0JKBFt3/86tFec01lJK5pHKt/F
2dThllW/+9a7qdlKU12VAv6K/aKz6/Qpue0ARbQRUerMh+iKy08SekgvYUeeYTNU
Wl64OXJ5OLWEe47JJy7J8EMymgraGtj5KW1JoJql8BN6Ww6IGJ+ATslfe9N5HJSc
IHZWn5VFSkwpKoRSH6R4FfF1E+0j2h9II1MzTG58Af/LbabfwGksIAOYW2Ax9PQP
6y4w6wbxsLFRLVT+zWMoMAdolNQyiB+i1tqr72vd91+sIeAZjFNPd9d/ZTDOj5e5
s9BmWZHWsWp7hJAXFiNjwDAjp733WlV4mOU3b01FJ7WeSztOVVrk7G9ckxRGGWR2
9Su7jx5Ti9rleAA8tZJgFdfRa5O65oSh35t+wW+PCkv3uSyvFEEmoG30gAzrrAeg
logCZrcoso//dUNyttB9KI6fqsbCyoVkrvjYhnlV6Bv7nvLHrtG2ChwPjS0faM+l
pYAH7QZPS6M6WBoFlgxwhq2FAN2fKbhNXZ0wAFb78b1d89MAE1JPSv6jElEnTQtk
xkuj9fS4f0SaMOsE0ZRXulb+gb/duRGP+QWmLJMvwUOYL/N9k6fMfyST5ArKFtoF
ZVJfynmPE5anF+43UhBd2dTldSmjHhss4wCimZjgyXWKB4/QJOqryyGvtSqdp4Bo
50bdoXsqzNYLqX17YFmcuD9qsfbfoWFQ3sYocpjiKYMlUhti6cP2a9E1H3vBH6ex
w9j5Q/y5sFUdmWuebigMZPU5OEzgzlKR7pCur82zE08oFR+KDqWm42q8q/vxsCne
3RV7vkC4mPNhifU2VtB2QJtay1vB3OM3aVoaN0SW/yQawhsQNvvwUz/tVTWLixIi
iX2MREdXm45RW/LZa2bIu8zRV26Oci2LzI2jTiloTEmIlxaQdgB1Kyvbiv4XpaVd
RUnYXa1u1+k7fx4YxgfNjdmqAiO0yhbu5Gs0lyggiIMqc7hcKGjDBRFRfCfIoT0x
LNKI/5aH9dY3l9nNE0TyunCGerbgf2LdfQyQDEggcXJYnWOMLfQfZJbKIPYk/wPh
WxNLW0dLcUEPofd3YRicSAzCugdI0iJKs6Hw4jdp1jojrRqlb+kQUrasGS51pMxk
8rDh7RQJHtQEPnP5CK2QtOcw+rwBt1kirOirbBhlQTWUNlsLPr1lJGiYINwKwcjM
SLPE6MM1CVcq4GtZpZXIHsn1xAWOrKVOY436VkcaTFvs49xrh5LQvj+YWdOryKQT
DSstC/2LZ75bDvPcQZTDam/Cy6h88Dwin/jXb9YIgiE1pGrJzVVhEIcUhREVRSjj
FLlVpnRBuPLYpaws74ZW4Xwg3ofGjJ7NSIhjmVS/FoSy/WqcPhLWOB/05wKr9bVG
ilprK6Rux9PpQ9O60vlKKrPi5Vyj9KAklxNX53Q2CitJJpanxNHIgGh1xHs/oArS
mJObLaR5tK9EX4nGCfDSCMx1bn+7/+bGizKOEPsr9LuYYVnqZ/Oes4+ABPArFN47
y8a7ZMtFQJ+ANBxp//4z4gOU6G3kJytByJsquqBn6sU4qn9qUHGl1WN8pB5QBORR
+D0TpgMBwTjoAjosTdD/xKNhIr6r9MaLRDPaqsxoKEhrgvGHkOE0nOeFDu9NPDcA
nlt0peVbvCqPTJ4juAR1Pr4K4m9VuUj/LA1AWWVgqfTQJZ9hb1mJo865X1JqUHw8
R9iBesDWd08yVLbWok3t5b9VRIMKZqc7M452jx4+7xfT1nVrl/pEvTtqPN/bK+ol
CNPT/t8lzkN+vf78WpgTkqEQbOqKU4Gx2LNnDYsJNJDGsJRV58jcVOJ5mhVTzbos
/k2lAxjVpQR2Avv2Y4SpEp7JGCOn7k7cQTadoF8jX8pL+txm4JKEYd1JtYuWEBS8
zoblUXro4CRMW7ZRnh/0HOxwfPkjZrQiIdM7fOluFvrAU9DJ3wAfsE4NpCFzKQM4
0se56wVAMMgPluj6CeGJwz9sO+/XY1JI3BaNWwUclni8U95NIQuqG6GAlWW+E2Qa
IM/Spw32NSDG4WAjk4duDpo6GkNlu4QKTHqy14BYWKCDldg9f9oeYhugNhbNAjDU
4Lm0QRhmJ/Wyn4zFCX8Dl1e97vf/ZFr5dONGZwQS0Wz6rcps6jg/LhJP18GF+/Ay
VrWg4uwiE3/tiB3P/L4pRy5PjSIcpunjeX/av8Jdev0Lxm2XDy7Q4MD6Ve55eK68
N3iQ58OceW4H4dQTGKUaSgHcHi3ePsAfElvFxROfmeAce7x2sP9SbJ9d1w6wQQbB
cNXbsHkEwNA01QAwcmla0wW9hVgO6Jt9oiJRYKGSUjR4SSznKNWmP9HiS2yuzVSb
aSW8JpbQtWSxSr7LgYEz40tAC2BJr43LmbDU9JnXuKQmFyT1BRvJcuAo2emrDxrE
B657amiojnkm6OumfF2CMCGh140Ez59UsDFEr2R68VOXPhfFbE9WDx8Uqn8pNiGz
yU3DfC/9lElf9u2Xj5+KAa3Vdj2N1CMEgUegfXMgJkWwHNu8/SJITAEKZAdcuhN9
oo1RwDWxXy3bvHIi5fY9SPS1wVtHSIJN0ZCEHPBhi9SPwWc93w9zHo+tpVRGByC3
aBB+6ltSUhGXtC3uhiG680ItBpsWE+6jytO7gF2DrEkUyg6wsJwGoo27eTaR+Zne
hQcHlXNF2wo8qtkMdFjL+zLKhRS3rUWL4Yn0zY3LgCICX1TGXNOv9Pf/i43LRzhI
z6bW4zpcVjs/hPY4yeglmJamcqKBcQIRn4vTul9RqIVSKmuzu2XfAm5rNX/Y+0oB
RlNZBs+EgfWEPhO5exoHpE6VTOdHzG+B5vNsZXiGNbCyiV0TTpMXwHiBSxeQCTfp
4B2zH2mxk7Uap0Ees2/cGFMK7w9a/z6P43iJ8W7ydvbuZPDHQMB6Me589diL+9Sl
hdD61BnvZ9uG0QomaKjNMLg1a5aB3EdmqqIdgXf32nfpO31CbHzCQT8+ACiVqYi3
bSFsFOu1/Tz/cmRS89vF89BPTxgeFLDNqihs2ecUAyvEyzZ9plRNdRE+0gNmM7Xb
/szwe/WWGTLPDoDf6yUiETpPU2cJCshbxRzMldnKMQIW1zMs/Ro1LJemfe+/hjgx
mBRB37lPY1w+VsUoWt8EhvN9a39Tgxw8QrXWm0hOddUQAZqmwhi2/vdisehpywyl
Rh6Z2gHYCX5Xe7USc9IIqrtWWzqXUyYKarGP8/KECqT7aWmrdEMQFi7XvYo+CD9D
oz2iWov/IQ1y4fXhNNDdMHZC4tLif6XzUPZY6Jp2qU6h2w75lZ9CWuHEDKidRDvs
eh9fmi/csG3+vuxDbfEsbhk8vrDsXB5x/2xsEQnPgfTJPscicmZRccDJ6Q5uguAD
4/8HaLIsafqCTe5t2BfP5XwBrqYWgzcUgyCD6q8+DKVmkPqn94VX5KSVZM8hOvU2
HRh2psC8KuxC4/66EwhJl/tgYpXrt/SaZjZ/ba083Aa8776Bu82rhlc0DulmqLMg
L9d9t5lIHXoP2jcaZ644pDVvDG6vx/2GPeUVwTe/RPUq/CsDmdWM+bKR7wgss9Ra
OIb47YClHO4N/JNYLkzexiCZQClrLrn8jpZLQOAabIRfnatlSVeS7QYChW6Scbw9
orQHz6jOMLaLxf898iznwTfrjXDsme2CwJcq5tMkvKCz8HujieZ4TO2diuMenDPV
bKFkpTR0si811ndnfLpI2VnU1JuByL73jqryA2GDJRY0E/EKenHCY6AC+sJerckL
nUrPTK82v8q6p2wKVIuBW6ZPwg8OKkRRPsuoiylH+RGKZMSsgoFaHwq44KqrfXrB
6WEyuUB/8YMipn5EqhEj7nW8C6o/g4ps9rd5AAvR+NDExnbvOL1EtcEQ9mAMhmnf
7KW/y634lnp65AbpGp4pEdeXEDJ35NW8GOoxH5ROijnpt2233s+CnsICdHdzClhR
g632oW0umtZcpvnJqARnao6Tr8r1RXysZj1v13kJh1mvjOhkGeRVDJgE6cnOVzGK
9NckAKsyBoiYQHmOWcDd+qzmXJx3SwnFLbkH1xn24XJt5uLLDeTHn8Y+M82RjMpE
u4SmlXIzbAHCFH0i6hL+Jbm8nKPaHwKA+eLKiuxMjfGll6V+dS3NHqfXQp0pOH18
1I/GD5rKGGttWCWdo537EGWs02qoOU63yQLOY4N3bqev67ZE+7ZewaGBQB30+4bh
l7qP5EVDgv6fYzfoQmSVeSQqYX4EVYkOBSoluSowcHp3VqtuCZWtw3Hz+H8MS1uv
mKJ6Yyq6VCaJoDXAhkX85Uon4A1/fAh7lVYpteiNViAFvk6Xt/LZl0lUNgQUxDAp
bG2WCQuS6Tmf0H/99iPZv1/IeFSKERwTdEB7zIt6CA90IWza4ZsLHdyjTEEv/cXj
jE/uTe+DvZJ4TBu+qVo3TPp4UUsapw3B7RKiYUv0QWsYOn4rwDl568cwB0hvPOhV
nYIDprM53Sj18c5vlIvbnHt17XsAlEYlMflgBC+PNnZbspo41FOox8W1zqYMocvC
ODNJlKXOM0rSBIXQnmfiQrQK4CAlY1galpBipWNm8GpRUpXaa/N55SnnsXMuOBqu
bsMstGH2Z9BOxWKi5b9yBXrVhjhKwooBsJdA8X47mwtxpZ9i5eTIwYj5Z/CVb4vW
PXNwi96wVkBea8e+U5RrNtC6HQS8H35wrtgmitD2QMlYipoVioTVDjSrQN7y8Bot
57Gtpa761QHzPUpG0qW7KILiwkPkWAtWzGVWuSgBrsC/Rdy9ls1+Sz0ohPVLWNF9
umk2SrMQJZsEThY+TVVDNUn7w9jZlcIJHfiWUbI66VSrRTvt9XmFxs4qGVVeA3pb
atAniyqIUcduT3zQAJ1iBZ/GyhOjzVwRk5EXOLQIEudHWTNhyyhG80HrEWok6tXS
d/XN3h5m75+T8i5e6MN1EmMqQKWdgm9JjLZTbNG97nLQqLqoo3E+WHbxPqDvqsSj
m6DH9KUN+yLy+YrGec44ZM+dNzeUJGfVBcjfU+65qbiRAPY2mgEcODxxz41uDHaV
p1mTx7ZqSUB5aYjJPZ52vRnzXRteS8/WuvRAqoX3k+uxIafkL9heUBT6y3NuoYkS
F3IE2lB3Jtg5Gh07I2hiyBQhYHkAjL/FB3FIQfcAtLGSSkrfymR18rpsL9vaKvba
wz3wCOEUhBSlHb8g9LY3HNTGx/4OsqUkjD/ip2q2WbIP0W232fhLgjePEMwO1pf1
lzL677PCHJ98nq7T4Jq5d/bsTFgURQeCBoRxxfD/fq56KOZw15hO1gPtEYko0n/F
Rico3DG57yWNmRSSx58wpbB5efC6y7OxUTOvyk4ekgmbp3LNfAPAQIx2hBP4T7OC
iQKwzts9I8QBmT9UpoJExZWg6vW/g9VQN3R45qaxcXpJwyeKd5wAQsQ25AYbLZ5r
Mw0IBmufr6s4ScrSY1q+rqUXW6ufELltBFny0FQTsjqXYmNExoJqwrlwACjgw5Tr
8zVgrPUqdTd4zlYoCqJxqlD2/R+ohWxNUY2NNSOB+d6i4Az7AB6RJiSk9hHFPUCl
U46iGJPPqkfbFWKB9qkiQDmpE5uMw3E0Ld9SAw0jl4vvDMpdsoPJoINaHwJPDgEW
dO3CGYgNIWa0bcbhLjThZZ7PfvMFK9nZdzD/ZBbvj4To0btsLrNI3FQv7XlKwRXm
ByHyEym8mw9kSCHrNyrQTErlK56alIVq7upKIhvhFjbfVqLMmXAD+hE9AIWGFxLl
ppDLlqPwU9+TyOnlcIztWTjsO+diLgPHvHIf8W6zbEKyN+1gztViHs3EpaxoYeaM
AuLIvQ3E0j1iGH2xeRLQ1152jBMPaUA8JDBCYMPmy/0FNOXj7pD5tLWYM+Sz9l3W
5L6yUU+8Hm9nKjEA1sEXYb+Bg8/LA2ZxdsaDUlrCZxCSiE7RrJ5jYBXV9OFOPfIW
qL46xeYuDpel3Pz6GtBWO6ms+SzvWCQPol5Of7Q7TR+n/6FVPH5QFINB7erYG9vo
K327K7an+nRGiP1CVUEiWQ/laRdxYYM6HDbz2TcEz63bsecnrZmr0pUetZSt4/B0
IlafoZm7TdtiUtIQ/oDvag1qk280WoYZ9a6a9X0w1BZqVTekTjcDBwJVFrIT3VH5
A2OFpgnGaJsxhrK3PQqjJ687rio8ouOxo/tHBGRw0KUhvtnJOYpDEV7DDmvy3Ldr
pHjjY2mqmMt3UDMWBBpOlNp60SJ3+qUJ05ZXnuZ+xExKj75RohbEOr0bF29/k6uU
dTOqIq7FLjZpphKvL45GT2CWBVdTu5qyv8A9j28vwbrhZBULhxsJksepBrPxfUoh
/bhQKXrrYD/G48kxbJC9qSdXKpiA3huASDHvuFbvfvQspDIpFYXnEATjlQ1Lb/hj
vtAuw/hRJ6bhlU4tXfhBUKnqkmsFHs7qC03tTPDX3GpVGltM+daiU7Y+Vb28Pqch
AyNayuBS7vasz4ydaTSpopTgUZuuwWHPAQcSP4PlD6Up6zfHQyY5JvZxrx2yat66
eO7je795o+YFfWCga+3Zvpj+2CtHeJLaqKUmq8vudj6zX7nuG/m5u+D5fA3Ju+Ic
iRZQ28hbzYreoBUYzIHuVWtkqQ0uhzQNm2qQqpDOJ4e/niGTi/x3p3oCsoYm+9oY
MQQ8BdOr3etBBbvOs28t2rB1/ffy2x8QjbT2lnvn7ShcE4wmZ89YQk8e5S20h3yG
k9rb3gq3ESLgTWHFp+6pwSa5YO6A4b6kHbG5B1+a46EOT+XwcnKuYbCjjFJEUSA6
jLQGWgptSuNaYUIbJM4SadX2gUi/HMHIh87l2r5vZPXGhn4azlRofRy7LaV15p4g
TZGetW5up0vafu27ai1KrqZcFT7OGaOpwMepZHHTH28RInNCnmHHZ3RgF75UX7EK
m3NBJEXjgKMGu4WApE86+bWCZkOfAgnNybB2m3SECjsdn4LCP8WnOZ7Is4ivs9wN
AXLLQil05AkqLKr0g/Ckmoa8fijqRRrE7kL9tiiggRPPaClSRqmL4xzycUiu/B6u
+YwEPe6VtLkv1MDT70YjwRbDHnYGdEQ5BvoGV0LUOVzgf04//3vOxSE/LXb4+q0D
3lknDVkXGRYNW7tSfUJed+bP6Wz3FS+h5TpLxwO5NtB1ZQYo8vzqaIffSeIU3or+
bJB6kdMzPgz9S422+M9kXHo04+5IKxsUocJ1aNKw20wO2wXaIBQgzDegmoBcTwj+
TYOWp04lr+s5kYEoHayNgX1QPD654S2imRrw/ib2k2qmLgEnKsCOL/ybgQucvVYW
pyu5ljVRclP9/nIVShLJ0aASQGlqZMAjm8Rq4XSrEYADQ0HhDcHwJSmkWU91X8Ce
UEVXshkA8DMb59Ih+BLGmg2BEv0jf3pf7PzvtBi+uCSvcViRt7m59cqfY4YY0Wds
GKx/4ZkVYeRy0rnIH1JvtjSEtT5qY1NEF4h76C3kFHktVVZkuGcMH4Mw9FY2KF1T
L0vC7/W6RAAmx2R1uM19i01oHxzv3DUCT3wyWGfI4dU5+FR8/k+pt4V4AlKMCNTl
EfiDgZdWU9ybxSn+7M4IrbvEOzfo3aCMOxaJh1catwrRCQYF2u8sqpBHv4CVjrbn
z9ETM1EyUQgaQ9mQbRCB4/dPoeLD4e9IS67RoIVIm7o5Gboak13zroHOnOrHfuQ4
tW5W//noAvlqJaZuKE6fkbyj2jwOyxk8c9sAdRfYl8CvNbpq8xA2F2ev6bA0URQZ
7WSlDiPQma5xFH+HU7KvZ553Sip1k/oqLwgxuXoLp9wN2PxLigMSq5GC6Q7Id53/
3G0G54kq20wNUEdLmZzZ2QvWz0Gcl1di1robjHPfNKMrtYFsiu+n4nXp+J5n9yB5
c5k9ZsTHUwWiB0kCRFQk/28Fyt9FMZ+HnBU8W9SQU4yldPPRxFRvVen7LFGKBpNJ
bRmcc2INP+N8rl1qk6pEk/++Hs3sHuET8CAVxOJRRnlq6Bsmewfc7bOwCh4c7Zn5
GWfqB3S7hdhL+XX+OxAH9uJxLTJRSBPWbjHk/lyXSmTUAn3aCbzzOeY9czm4cMci
4jWnqvWbgG4J4g5je+AFUDcw4EQBX+wP6f1X4czpVjdnq3rcp6FLuQYQLj9sJyUA
6bFEtOnQgwYpvudGavJZEcWbrkWfaf8VlQ8aKmV7cZYrXV3bZPCHZvtBWB0XYw4E
ynV+7XS6AGt+islerfIt580dTU/4z2dlznDTLfmfvX+uuHDG2TZPN1dIcgrD0+3Q
riX7vnp5SBkzcMjmiuJZb8o2bDKSz/gbm6hFBibsujandheGzNpIZTmlK51CHOnk
1IuqlhwsSgSPKFlacJs+y/rTFH+pfx8+V7JU3s8Re05wxzqpH2rQ4RlDoVa0d3Tt
DQnM0bOKy9/EtwK/OwMK8yx/4fvGjI3/pperxNTg9y+sfWRF09NRdSwIw/Pvs8ey
++A4MtZCG714TNeXaDU7m2ybJuvm+hTA7TFDZWHGoyLBtN2hA/JzfETuPkczJJZ/
QhOkiN4mYuw6Rkx8rALL3udBHhPeYlWdkauvEGWgrAGwfitSLJeE3ZyaL/bgmz5K
06PVqwcV6cc7iVBrrbyq85Zb1WSl3fAZojm6NAHgV/x7Jw5l59RGFBII/quhXCk1
5+6mt8Rhx2rd8mQS5IZiha9F0asExGHuZqZeCkD4K6l9fRAuvJZ03v1LTYUECDFm
ySVPAnr+Hcfv3iGyGt2HTENl8Q9s3veheroaH4MRoqEqA93+Etcf389AYE7TQSZ0
LELvf1roM/yVLQtoTpcwb9VE0Xp1ZWfoNy5bVT4llNB9W4fL/diSPfRAY9qFGNFQ
rUQ/SzBjaxiKHIT+LHYFCQEAcq5nQCoMSurM+Z7bVVDNnRxC43HotgfsG6hYKhEE
igV+Scv/Eb5FOW/fj/5E3p64tCi0DkSxvp93meQpbi97UToIQfdDj+c6AagHKzF8
oPiemgjdQggBI+pmkwBg2lpMP0O9jTrY/VMxJwe2SUWEELmkY1YGB95nIlSQHSyj
9g2B73IqHX5hzUNyQD3bZ8kBgYIw4vdAWMoCQQsWDCe/XuVJABes0I71YtjFloAj
399xIV/KeXLeyXrjRYIzB15//Wsbqng/cfcDAk0JMKo7PVgqWpI335UOyjR/leJM
0SGkmWrFLtJBoBmak9mIvAri+U6+9qplb7lqtj8vVJ9IMA3Bi+6XeSfpvf1YtKKz
IcRSfhSWaTXjq9Y+vbYKx0vL/zKnuGkPkuqVxc6sNGt3o9l6EfKbaBnwfC6T3UQp
zCJXU4t4EKjefJnIPAXgh1SS6XyCRJS9wvuwhFdTIeQP1R6W0EUktuK45WAgjGKa
WMWZcQoBKnNCSt+zDb5Cpwjj40I0gQuNYY8KYSocWl4wx4j4S8se2blVvaU9xO2h
P9DD1n01nzLkaKXN714ustmR+tjJqJ4mPJ95uPeepaZzY97su6NNwXvO15HGfPnO
vRKpzEteALey94HEBJCUAECc4N8AgmdvRNaUmpwfHKmikmp5ljDyDGtSgZE22EPj
y4dKJsM9OfId+t6TU0QMry1pHfHjM3cDyLr2O5t746tyLZeyocSEzezZGHDndtc/
Pq14OjP/iC1xiVEyGz6KvELR3BP76/4nZPj3oxzy5r9K6anRfAK2pXaoL6CaTjV6
OcfgQfTwUCnsGfrEwn34Cqyju10rwvfQwlbzd5f2b8Nh9dkOrCil3uiLe0C4WIup
9nSVwbriGrIqt0a8VFMN0qRU/GDxP7VJGwqUKkmtjqiEGXZQk5V920k5AkdD2J/c
9PePQ1g0TGBoCELn1wMYo28jD7UmRyqFPqPYtwUlF+SYeHVWnAg7fZnCWQyuNEn8
v6Q9mlZTEGOzQYXTB05FAxCMl/18EkckP6XJEyE/Mq22wE5Y5vMql5e/Q+QKKLCj
LSi6h+UQslMLSy3mP1fJv+Gn10fEn7JNbdRzMQAbSygav7ajgJESabBq466IJZ2T
UMig0iQogi056uUSl30UKM4AFlG1UP02/02vCWIkmnj0S8GLtcG9J7xE7/2VESeY
fIjMNDafIWGo2mEhOwFqUzx62AKBISh8J7gnUKu4Inq8PFd/lmHrVTQfZDNT/01x
+FLY5csHqqCdAACZx2BShHHfLXmWq77ZWzWqe6yBbYRN4XBrXSpxydlTcZ0Y22PM
9nC8iv/M8vtKJYJQ2cKSfN0d5Y7Nzv3vqFfwIDP7pXPBx3GvKy9WZP91NCuckAP7
4LxRhmsiCChdnZtKVZQpjS9oFQwnCvH7jRapyWcTvxQTDg9N+qs3+dYR8YaYUCyL
SCS96wYKZLqAUYk/WuISWVEIgYM/zWrNUwiS7VKUO3MMnadyXqwBs1GXTDNgyVoA
O3UVycnv8iZLGjH5bGu38kZt+UusH/7fD0oJ+hmRnXPHJ0Y5Ek+ImBr/dl3EtNM3
3lsdvtOnR4nwOIkqC9b48TpMIhjjAtEz9DsPIvHk0GDuDnLl0RMftjI/Mrti4WiU
SRFoWc3Y3SsGUaVkk7Oe0CoJzM2ys/N9YWKd0I7kZuyVsUSp7l6/IRwnTqs3EaWz
xIayaiwjTlGazX1fyy4jN0cs3ppzfdUpQmJ6mBa6XaGRYi4qoQd+SZpeJIMoxKFB
haNoVGI6X+JLwKiB05ZwE+WSHY4Nc+L2QU3EUl1YJaqXigluUeyNIpB7J3IJvroA
ZFmQsFOPOtt6fpAT3R94ZD9W/pKiHlhWnmNez7pX1vPWXdpDzdBewFAIQGtufWog
JBN8vEQB2bYNIzNyZm7xE6C99bhAG2AmRxTW3PILsOndUgLt+B0PhCGQKlXVx8Wm
9L+nKhHh7dEeKFctpj6b5qVxw4UncmbtnXBbdQuxr0erwFHi4ZwHjvZy/Q829L0d
fgcXJTccie51gYj3Si+Nprl5E2WORKyAtBSyrIyrkwQEc3cULIjZxd+D88ovX1Vi
ZphII6NO5jZrzj2mxvJCgKa/7E5Oo+Rqo3doUI93wcs3soSlMQamkIKUSxkNUhMJ
qs80RY8YwS9H+Lk+m6i+s5Sx6bDLVrCbYw7s2LzKUB3hK58S89vL1CHGLDYDBoDw
/4GwT5HMKft2LRDQAksYknyDfr/KLfw6N6LAi3ibuPE2Ki05A9M1bXnMg4FOG9IZ
gCI5R996o98rNIKzRtCIc7j+QrlBDFiH5DzokD8ALAOIZYgI6gWHWhWtfCwI4M5N
HPqvt6ub2LI6EiZjJB2hP+BAWsjJd7MaDkRMOPgr94PPftLiuZ/urM5j9ZfpM4jP
YFQRUWpGLcYTaDG7PyfpV+bya9MyNpU1iyOjv0jHO6wYMUAHslk3bAKGZzXNYhwx
HEmLrJbES5dsWWxRE6LZ0uveDxnURG8nGhTsXMq61linOuH3pHujhVKGEbyPHlNZ
Ae0NkAsfb4+qj2v1ctP8WKki411WARjQ4w8LZdaoU2yu2Wqf6sVMJi/ivz+BrfUP
Pt19ANixAZmHNNh8oGnF8QS2d5ei0dq+lKLNbKL4ZhWlWml7VqOlyc4rblt1rieZ
pXmPkiagXGYE6E8NBrYGYxkCVDDrA85+HNBz4nmnxLC4y6+jEsVR/1crAnQX3Vov
+1z0UOMMLmH1m3au+edNJMlmJE+EsAUK+pv7Hmqot4d8+xSJz+w6xMFiX6wGhyT3
gkthKtOVAlAeP9y8J9wenqAAtUG5K1TNTUMYEKkSfb0Fog/Ahlap+OTW4aLeZWFt
WsKMLb7HA0+cyUyGWA3uuL+VKcsYQuari52ajhf58Vypf1iDtOKzncYutpRXkKGx
P56TeFPf9HbhQW52iEGFDuzLUw7ALbrzte67hPm7ZuGvTbTVOeY+QnLlz2cxejib
SoFtFApKxjti+/0NpZWf8YwWY2QBDxk80LhOWA7J/gQeFbADplVkHh7Xp3in/xI8
vwq5+LnvHhoP6VCDEGpdBDoEtMZZfzT/CsBeLFRX8KCvEVWjSsCHWQalQnpLYNti
zC717CXVfBKkQ4qjci9dtJVNVRa9KaLSwTKUDWqessNBakqIgtqGrK6/XsEdchBr
awAaLUYJAmyDOzO3YdHoe2jUSi9VP1HDZyMTGzJ+ZLHDWyPTHPK9nOXiS7K9dpSI
tA4vXiVkr3+yb14HtZAr1nQjSXrEtFA2Te5GryMNr7NrrxK5p2Te1k5g9sKjae4J
6cVuYcn/6Icji9oRsYPJOzxIrZyxCnEJ96QYj0O3Iz8PeS5DKiieADrPnTzN4SeE
9yrZJxHkjhGeR0yh2XV6ybN+Oul1ohWwhodVWV28GYqQEXTBJ82lLiS4f4CRVpxg
9ObCiTVdIjeOnOhMlBuRppS5UCErRGdYw6IIv0ImlPIzEfZpmp2VDj/Y0yLltEXD
+HlKD0n58TbaRvG0O/Rx2L0Ic9xiJqpNZEUzNEAUrlJBSQP1DImDIg6ZmPKFZ4vX
OpGmM8kuBBGVgwMua1CmdYTLL1ettEZ/VVqQ5ehu4P2aGM+UGg7Kk47rR6rjROI2
A7o7qEeti7snjL83Ak4CwkJhGhrk+Y1xJjf8bV8LXkB8FweQjnUFPqMcned3WHxL
IkQNQAuKhTJkdkJjX49uykSpIKTKBw3BhR5IaXEcUyD/qQHHmxOP2Hq/Jfmxje/m
RlXiDqPJ4t+NB83s5tQmpkCC4jJohbOglVDIPO9MNdYsK7R3S4qxGoxIc1dfAXUz
Dd8y1Sc/GINijncNMqkCmxMIhd0tR6PbFebr1kMc8eEubyI8BevLE33exeFML2T5
HrD2yWsJ8K3drTDnplsSetDliZPbzQP+gHMQ19UxJW8z6hcQ0qRCLQ61oknVwtUG
fFO0hE7HSDVBC6dlYClU2bAvzanKHp8e/I3LDuzzX/UcLxQZ3i6SDFxG6Vws5zJK
sYOOWiJyGWIGhqMxB1BXwNxDxbkZfVahkwjpZUOCXRIUd9mGOOb9qV8bKvq1YhW3
46K25TyGJSSHVHcN989n7u/faUn2uxXWAkU0Dj+8AmQEquDbcp65XGqQnL901LvJ
dJr6pXTpt//u6t26ve1K++wp33YBjca75fMfmEjGE7vqr3T29bnu9sMfQ+O2pjFa
ppV7MddHWBxHU5bBlJBDQi1wlclK9tANVlg++Vzn4F/iNbdXiv4xus63UyD/vBwS
x+076hwFIWrsCxUK0IQvnbh0BWe6frCMiQNxPBgyovaUw4outcX1iyL6gj7cox+T
TCWahh1kaLjtez9jLQN7pNisq3Hox837nRFsa0nzdWAyr/v0iIzcyPY3zeJ7V075
DnL1ntQI6OyW8uYrakdPeOFmTDX8vPiCeHZ25+jSZn0ZZTacDF7djFFbpm9VDIRr
ZxrflX9ep/gilFFzOb1FORkx4I07Tks8Wvf8mSD8fr5STPuq9NfiXAgtM/Wncktn
OcvsumedJq9PJL5J/pafD+9wdWJuZrIMHlmGeVYkmxDwg88xq0H/4paJh4n6a7sr
h1jYdkrRDyqMqCS+iXOKHXCRr82Pzf4ZXX+oZWyS1wHyeZ2GLeyPtnXAiC2CdkJq
OrRv1BYZcXUE9+Lw52sD2oHtExD20WZPdOPio1vGq+VnFd+zZHzifNGsS0HzLJVO
AVMmgFNEoKy7gSsdKbxKPH2cP0qmxvkgT+WGIYIHxs82V6qD3TGfi8i0NngrjxfE
WJf3RBIGGDgiDaNUMFHzYoGzoj1MrsgfW1xMxIix6k+Xvz1ZMitpBY/sEQtlEIky
vY+H2NKGjvKjL505rJj02jIL/aQzGPqMj0pLgsGiBAn/9Bk/nqmZ6d7QJyKGd/4n
rjwlwJI9zvG8xX8ziX8iCSpW77iC8/BeoUCrctw98BTY/8rRF/DJnfmxjYdzEJKM
zM6zzMdp8bfNwQN53GJaamW01zFqp+zsbPAn2kQOeoVdo+E4a5/DPc3cRQkgXQG5
QJtIUfhG9A7IaAcFqyyqm9A7sssbcN//A8ybpj+pvpLNIhoi55cNchfvJh+gpkjZ
/G9yiatsIraJxvmHKZS9RL0Zyed9u9B6t6tqldqY79RHpIb6EUECU5ZsNnEUSujN
qVRyQLpN/KNuWVtShsohsSejHIKRHPrwlvLh4fTUTnbxxpcl3X6oIy50nDWWv26G
SJK9dcKpMciyCHE2/eCoD7ZtDOQTlrknZgoSsKvmV9Yme8isYGc7LW+DnldSiJYg
6ZxASwJW7EWnixx3w15mY85XujXjBv2GFcb+iR+nsGTZewiV1xaweFuiV7ZTVrSR
d+O8gdIJO7UvLjKYdoDPtp4SjAkQm+28hDUO8fbf4mgtl1nlNQ+T6/jy3vy9lYEH
/hin9q199izZac5GBtKSUJ9NewExhMfb7lyGyOpIzoNToXrQvQLEmgtNXF+luMSu
jZDNz47wDUHVduQejJ8H6ezJNREx/l2HMt4RRdc5MgnvmuNTfyavP3/rQrEXyg2L
1f/rCCp/vlvOz6aJTnGM9YNBgsk89quVXNA8gYvxjKzJzYL6rtxDnCn5uJoiAe8Z
hmNzr0hFBjSoN7Mh0ibfNDrbymzy2NBcMqbkZtrxPqAUYnAq60axL+EZMAQIjaNv
mQ0nsowfgHOwWqe6I7CXbQ9aRC4ToNbzoq94dDlnkmEmpRQ/BVxp4YuQVtj51BmE
CWJj/lhkmhJ44/gtC9dkcLuRrUsvSmYi0dFMk0rhCxIRtl18V0AOHcSgG2vVm2Bp
4OlhEsjO4drzEfGsMthz5QXPMfQVCUShRUAoB/Yfcona3y944107665W0zaOo2kf
9cDjUBT4cjKPQ8xatvA877NFpjxRwOIwjtkE6sasyvTvgUlfH2h1F4IeC3Y2LlgR
MDCeRMKt6GSDHXkxKDkuKI1hNHrcbB01XUSQIiVvhlGc2yboYXWXoVxZE4Q/gvZl
9m3Pu3ZA1tRtsjvlt/15ImCBobCvc19Z5vpD8XjIZwr6ik3uOfbDV8ElhSCK2r7q
paLy+aubsryL7n2SVant4DUoK9va8qrABidllpmDJ5BdtUmJwmQQk3Ti7aRy2aI5
VHT6O4X0p+6OnSus8wkWj++LecUXdxKUWOCa5OH4Dg5GJatHlZWnIp6CLc/IbQEj
Tfm0GDuHji4LCSBsIWwPKDtrGGun3IS3wXGQsS49I8jL5JSwG2J//6Wzay6f7NNr
RkB89vfZg9lQYPOpUVRgjQZmXXZdUa7s+h8JJrTUKyBBul5tqn77V6RiRD5A7X4A
ze27lg2HJMezlS0gnKnrgtiT5GxkO2e6SFW4G/ostE1Qp4CnDlLQi/s6Bx3buq0K
gX6R7mPbi7jk8qShLcXlycveWQmP5VqoE90r2GlwrBjEMt5zyrgmyLbc9KrIxtLz
PZbSOs21/J8/4Xuh+GQBN/58Ciyn6IrbQhg/pFUBH6V5ay0ZrqDT+zp2Ep+V1NUr
7NXLV8m5CNXCHkr4gGS+iO0YuMHObZpvTZGc/pwvznoYvyklTzjhh1Ll8F70vGQM
dJpuN8VEcnEF3nXO1ZX183OmeD0Eh2fLxovI2+FNaVBQTF/D+Oj6Zv5/9TywYePK
QbHMfxzJSJgXm1ZigBL7V2hpGNf8OcC0JSFGBTrhYtkfNbAjIalOtfG9aKGcyVWF
4tPi+CBpOTZZ6Q6g+tpiNre/QGGmyiY3we5R1RJpdXwFecDOn9xP9AsZfulq9mDK
Wyez2mqk0B3H6XHjN7XCBMcQF+bxpc9Qth9DdwO9cye0IAQuT7/6npB7FOEdiIas
k5J4BdTI1xqq9RqfRK2qhqkBlTGkPtTbV8DwHtimD3xE3Z4kgEOXHGSvWJp0RtJq
8IfTnIXEk+Pnw4Lm1myY7rGfvmLf5hErQgdxeaCla58aQmrhKoKZqvecMORYAvo5
7z1ZyWhy6AdeVH11c0MZiu5y4Citnxkq+wZqUKwuE6a8hCdXZMLB1wHPK9HLpGL4
QZopZG+91yri3NqDIpco7wmCVrDnqCBKP1T9M+JQZVif5otJl/CddEpSrzmTAFIo
8WrGWljDFY5c/7+4dn4QlPCwQLXlXlXJyO6FwCbzUSX8AJa/GTkXkKg2v2GZbaI2
PEIsBzo0mhUc4ktqtsvAMojkSKB0IvEUX/H0MrCiOKDzjRhM5DPU0NGLSnZS2bK2
YTk5+IfzJF7MyzkSJF+69CUENaLe3za+NDct4hD8rCk0LmMZtRz3KtBRLMV9ilud
sthV4VS4xnyq/eM662qY3DCDUgjdrwdW6/A4o8P0ZDZPae8Q/Tk8u6X1TU7637EP
ZwQ1++ap7atujpoZn0nDGkQDMXjqlwzfyI7WmrM7X+4lN6XungkBgxmjNJWWG4FV
NMxok1bF74yh8bA3eg0ZHFrshHwqcrkx4WlZVt6U6DsYsWmqKJxyDmSo9cjFlMY/
980CiFN4BUeHfMD6DRqEiqGFRENVdbjGP1jd1eFodjyYWdTGx6hSR/9pVBgwUSgi
ncpI3xPiUXagXNT9kyIwmxumXpmfXSM5v8cZhcH/EzP0qItCT8AV1AveqpGPYgcd
om4iPExTb7u+3dltjwItrhmSqOnRtHxbcGm39nNmcwdKJ+lcaEdL7lqx4OpsByjs
/fE+aKTt86nh+CzznvxNtQxaIt8j1zry1S2bTRtP4T2umQPZ7b3alygJtAKbKzSb
cmUtPj79eZBtdEVGskxV9Jarox/illsBzQfwaS4VTsIKsHPP6Yq3OZUMLyHQCYYJ
qnUa55TkmwzNpkd8CNpETjV7kNNyYkRfsjLpPH66giHeGhGWeDfv+LVfmQ/xiLR8
/jAE2SbtumF9wP12wTEbGS303q5O1hGQYVI/4eThOotQNP+a7QUOqsA4N6ynMKBH
g7xUWe6HjGd90wl6kQfOhc1Z33MYRbo1lPuAqVR8S8jC/KBHoqO/nxCTlhXdUBR1
wB4WsC//3muFfMHubPCE5uLSPf4gTpgauR7XJRGgnk6RwgzpCiuh/cAQpUUiBp1P
+QXvVu7DNCnOoRY5Y+bw0n4lOelFwJuFmkTUCzTbKZfaKgB3pdCi9t4Jwxg9qVkR
1G+2MLiOficz1+vHs/It8gK8qj7JcMRbCwpmGYwFgC9sNVrV2q0JntqzdINyv/nV
uPYYpkRPVGgMKTJYJw5+KzF4pBV4I0Y9MYTIyVcRSqOBOquOccrK3nNfy4I7zDlE
DFBsnb9IXsgVRwkX9aL7H1vz080Oa1zCIDxZFzdO1bpPIoBoVrxugd8X10g8BmNT
umtprlTmaH9sX9yeQYd58BAG7+kH0LzRMuZviEZ8BfyRf/EyJcezvf6jlEV4Ovvz
qkp4J5QJNXQ+OJTsCwxkXmDz08kBXgBvXj54UA+tlfmUhUs6BXDURL1wAqxU5tzH
9luHmLNF4cia31v+atf/rdSXbelftg6iEyH5PpfuV9r2JbcA9hNdD64AVXul2ez2
YH89DOrcvdq4PNUoF+N0wnyNnYyakOAJ16FjB0VSaxYX0o0hhzuEWTC05Zw7Opa2
2ncr8ufS9DrVTIolpF4KHbowD3ObfWe7ulZNgfQv0MjSeH/4hY5f1BXxJ8dsjxL8
FwDwq/Sd82B8Zsdu6YhuC6Fl+C24rqrzV/CNedYwFG0JV1lfalGUtZoJ9KzP94E7
F9UlUngpDH1fv+zONSFgh+u+tcSyga2JvrY8LsBVC10oHDEvJjiRWDoPFjPYxxLh
e7rbKm+Lpxu8FTnbvWceQPdv9O3KhmPSqnEwU50/qquhIPvHUGfAP6CL9yhTkLZe
KdqwwnRVyqp2Vc3SM5yHwnwuwbWCqWq7b73uTzjz45d7F6j7I/TFxhf9XeGWlN2u
NsMFV8/4XXEE2rKCGRgZmqCHItLL9zOCsz/Y5vh6AzQnUKhrrVAPK4Pk4Dgquc2Y
OEfLnXxx4cDcpfYZ4o64u1wDVgPWgTjfI34n93Fp7P29v7//3PJb5Ps1NVR8hP4f
qhAzgSj6zMQSUz5EtYgK816wDrepWytiggcWrqNuqGm0wqvB7chTOCGJE4DmjCwo
bwXzDl80AYKX26rCzFbWo159BZWvm3Lc3io5/v2TV74+EL+ipc9mP9QLciDf2U5O
E61goamT0Dzw6Qp1Zc77iXlCghyHGdMRQEcXAkoYMxtX6Zt56Ng1EiVKvl4qoGNe
7lC6JD+MGDeEP7QxqyAZkxdDZH7+MGoX/JikqafuuniwuZ5qrPngbocHpTHK/CKI
GyaD/nd8EqbPsrNrmEoEHOEkdEg4XKoMYQS8Y5DOOVjH7tVbo4WJTY7V4Hm9vhBq
eBO5QM7XD0ZJnMsr1BEey2KsdNhYx1sW51/ZZ9V0b7C812ThdpXiLFAzYmOo4wFm
b6UAzN9HfILGPrsmNaeTUGgBIrUumldW/bPl1lHr8eiiwx490i0rQaKNgh4nZaM/
fQ/mE7yS1mNa8hiTXRbUqZ+Ecg0cSwjl18ZMcKSIkJ3IQPU72aNO4ygcGmsYjuaP
kUeCJpJ169rYEbZP7L2h1TCinlqFPi4SYefmoNkY7ZqJFl4YcIbOu1LtLTxq+aj8
LbovxrtaK2hX5aQ2MzjUukJlptDlfsq+F4Vzxr3S6a1NgE4GIXO9OtxvlWPF6Iiv
rPf9o0Z84odEi81fs1zHKGUmfMJ6qUqW0iIEqlzF/HM0ucVU7p4VYJj1vmawbfmh
VWh9guVn/lJrUkb0na29RJRIcuhcfCVbXfTO173HLK6U0iapm1W2YQRN3D70tQJm
66I/p8C3TIsGtWttGkXTi08mNzYesTTDQRl1HRrePCDj4TxHo0BKout/Bb1xoncD
tBzYglFPCWOP+feUN5dbkBOCKAic71LMJ1dd8WWvhkdZ5jVy6kFbOzhRnaLznLXo
lrqPKhcrY1aXU+Btm7XFiOFTdU+D4fYvCUhXjG4DUwnrKurEes1t56fDlwFgji5h
gDl4xmze5/Lsru9NM+42T6GtuiqKhz19gHSiNFoZNAov3pJan5UMAVQ1YWt6g2Jk
FVsO8aGNiTaPKPCcPZ89UW5+7+Vozn+5+QRq+4PHvyXkpk8Ii1JeRRJOBUyenv1i
58PBOmM4fZm+ZEx5uMY6rKO1q1WIK2LQXgSRzIW7CfYut8lx6KquQOg7OXNDgXy0
Yl5IDmNqUH/Sw3gO9aJQELvOW0fLoW934CdWsh+HVAbYtaGxhKhMDNWGyPzhyDiO
1vIhCuWEbHUHCvQfADUUrfswMHBTauuNdQ7dpffPhGCLGhTLfJ5xmSO2NcUxqepU
kL1V3KsqHvzD+t7K5ywgLs1zx2jAgSm8dsWg7wc5wTdgPWmjORl4oWzkaO7A6aST
7x2S2FI7RlC6jWCnqocNVPyfWQFuKuV97FodG/tax8A2ZI3yqq/utfSUbOu7a3Wk
hTjH+XG2dp/aQl4jGtsXygfvZmAMZg6PzbPOlNOcM35qkuWLeB6StP/3ZLBgRwPF
dciNQKErJK0zxDA0ZLU20KCzkBA07op6nOk/WTaqUwRZi/iQRgC/4HEBkx9uOP/G
CQJo653goMtVi458cv3u7cd9f8sv/8o3tkFVCT5Sjd4AhYCLLVEW6lHP+E+aR7nT
484M4o0kppc769WQMIud3kaJT2L5PlJB3dUhlPd8fjYks0uT6hUjQeVbRGKAWviH
kpFq4y8baL2ZIi9/bdFWXljcnoJ17olzZFuVU3rdhc3oRs2bb5pHt8SmcU7tPzWc
g8vjQ6CYyhb0LdJOQBmABrQtlLH+KYXIF4D1iJwoO9ZBGSkTxptXmSEtiVD+w5+r
sj3Iysu4KGD8ER8oPwYMCZdKKFb3J8X05EdkRB0rwKMAsjr+GDzsYsAAeQah2Hqz
HDc2az0W/ldJ3o1HRwG+ixb8lFah0Pz1VWOLtcjyP0AY4dvdDGeimJRUCDdXfUzc
oOAnHB5vxwkg0aHzHuc2M/i6rumbMx3Pc30zDlPcoIvHijxNRUJA5khZExTXEB4T
7uypPmcKdISi0EdEid2edgUGiLaoNL5VGEmPg5mhn8rDiNBACssN/m5WA8/FZ9a6
BALP24bOve0DzNR+9i4GZ6b8yGLeVW8aK8F3rbs/M7cqvWEWafJFqhTzjRbxhtRK
0eNUNkKUWDw3J7pGETFV4TqMHKww4/WmQzCRhZMakgHQQ/bPrOTHbXkfVaEldnJS
2ieGisZoHc9dX+UE7HxAdT4VXyXpxUkaN521sY6SpVrSEbAbo/8Z9HL521G3Dc+l
ko4RUbXiBkgQ86HDOR5JoK5BtfkUuMjb+hhulqHZVLq4KYOvox0uC1TxVUTCzr8B
sPHvff7z6Fc1xWOLFFWosmvgsIjuLMLYz50pQVr6IjK8mU/cvo01aeKvUcWx7Q/t
YoY3N0SWB1TsvKlYPDflKf8Q3y5kfMgj4Ci4SRtpCG7F7E4NHNaHD+FDZZW/G9kI
PzfR1XNHr45GsAX9RPOxk3J7/MSW6PgCJP08vfDUQ5JPJVT05X6Jz5aPVz48Pb3g
WddifcazA3rLNfuXMSu3bytK1YwrbZM3BuUS6uGQUfldJWqpbF6GkuSuBPMgKGnZ
QZSxtADk+XIOfqrDeBvoxV6mKd/6otpG9JFZeJaRKTQ3zj381tRZvzuXl0g/cNLN
9SzB2XYVWlID3cuUwOwwZzaz4QCfqj3OlfOTabsm76182ltXiVLCiADW5sIcZD6/
dnIt+FhUJO0Lli9onyvZdgcuSq1JT5Fe5nFGLtwjDIyaU/mShvJ2XKBkH1HhKoPr
rdWfN2thzmKB4dsvEg7Z4mdXCQsJS0m2JFtFajFClSC5k8WkwMmpc4cZVrCxIB0J
g2mTC22PAN2Gn/5qeRlxb2l4fUS4f2l3GWhpVJbS0Her4V+NCcD8hsghFIH6V6qW
ewz6b10hfrqDoOnwyKlxJpsANPWIJPE7iN2O6G01pLpTvDQo/PTa1dlI8nESCnPY
0Q1uq/w9Nqi6U6mWuVz/uLBR7YnBgKgotkJ70mPoOq+r3ONcYy6UIoN7maRXtRvK
ZvMUL6TLUwrgTLIWH5pAa6IRAgt+MpRE2puzBq1iIGsTTqaZjX7aNOOnH3axaMJr
oXr0l4Kw82vshO05ApxdzYk7VpBRTCOPxSciPqHKHsby523BYIxHh/1xJ72qV9G4
YCbdRuHcQnyclHuiXh2afyx31OIUZV5Z/WcF8A128jwI40dQeudWQw159gt2d90h
G4cUYz3gYNm8Ss1uAw2tP6Vx8Zsbxc7WW2tKGSao1yicuJaJH4dar+l9KiOwjZwZ
e+4PJxTq3cjDDEDW672JaACCh0BqnnMBBYgH4VlGRSglwPLtP5uej3PUNLIHaFVc
WBFQ6Bm/nImddgQRa1bDG7hgYZeEnnB32Pu6n3YITYc1eBonjh+9EED+/2Vzs5eO
MaBWr8BJ7wu9qkONl0KM7OPKbfOzF2f6+rQhFzprwczgwvw+vFXjji97SPtOwGhz
hQxPRdxe/srXKh1PJiVwerN0wGnXeLIQgsreFPiSYdLydEGeF/PQFdJv/A7irsbo
h8atMmGIKMmCxOZwwFS2APeFk7dSP6dsNe9Jzy+9yrTNh3FkDOjNBdO6oxK/i7iJ
JNBqLNf/9+losPWNv0TxbyNgneyRwYzO84+0qyyiWRgJ+nzI5/lgcN3Rte4pdSRy
DujSqUAsOidZBoyvFNzYCU6tyCBC44FWasLXbHwpsRfuP2LZUEEl6WxpvKRrCWw1
9QDFMkYykd3CjSA4NowVL8AQHQgoi3NjPDBsUR1Y91YaG/IhVSYg5qaALP0zT7Pk
xqtUGGidbIinXdq+y3DdLCFf2HbkmFKb5EM5FYNw28IF2R/HXZpNmG8KdKrfvC4t
fy2562WNFgXosHwl/Qyb4L7hc+JxZPX/LwqRmbOWn3tg2Pq96dQR2oYJjzZRqJKc
1bfqsMKRJBS+978tZjsxLZXwkCbJvXKuiMl0bNfAfQFgZIZO0Zc/LewQ+XHhKcr6
gYxsByGDJN7c7EH9CK+u+4Phq3/E5g5Jh19SgU/PQdr9N7Kf+qu/aUWW8+llVwmq
oOY3N7Z/UchpEPLPpkqgVDR+bgqkqvZKL/DkfEpKSeFvu8hohe+g+lDTiU20CSH6
AXQh8C15GeNpVjKaBiwDATUZZWNr7RUlhpYlCwBT0Aw3ee1EbV5/Ul1OmW7B6Wip
SHromYcylpjRlwG5zKlXJvywmIcKsMF7J5L5RDO6g0p9eTzYfeMztssniaWW82ZW
sB9ydX7jyDJX3vIaNvGRXkcJ0ipq8M7p0cxn3m9ZkWXkPKOsJ28J4snPCj02TwfA
0vDPoI/JtUSbkt0ljCRJ2sGElWhfDkGFg8jI8Kx6Qr7ubqeuf8mHFcK7I1CNPlaP
MGz7wtG2ha6jQ4O5FejF7YvljycMp+JbmeGti4l4UrKhMujb8E9SSunr05xfgcm4
90csnL0Sc2B0azFn5EgxxC+I7QNWmW6ztTFjTJa92ke1RXmRpT0VVQnedSGqE1jv
qRjF7tnY6Dyq7K6GzedmifR+/roVMagd6Mu6yDinPm8jknRRSpEBEGRpPidHyjm3
DOC3j24VFhQ4lioIZhMa0yTMxnpeoBb1lQrtWTklQxYs+CUcz+p6eoHoPn+7eao4
q+Bo4c0DwBv8G9+2Bm8ySWwiMbaBw4VlMRQr4qrrUVuyE1PWHiFAplpvjmQOdN8m
WwARSww5ZXB2rqdhelz4aS0q1xpLdEauQthJu2TtLdrJYimLrRdYilnu0XpiQapv
x/unBhd+9CJncC6rGY01xLxRP29aSFlpMliANritVH2Citdi/ko5X4UsFMl+T1oZ
bpbx+xeiWw0RrQ7HF8d9zeBrEnBHdmvvPWFmmhh2iFtn1H5zgGgOOTZu1OZDh4vk
ghuUNAzAAsSHWJC9NFfoE9B+Mb1lGWtq2PZlt3VSg0LKh11g1C+1TBD3ndGCdx7N
KYjKPL6x4du79Ur52qdUUqED39wEKe25oC7XZCqPk6Tr8ZXDLF0sBCxptjgzFZKf
QZ9RAyiVtVAXKqgwQlnolgJuULd320xLYSI6u7LPdiYlFIbw8EBFjIuibInJ5SeX
vteayyVLWDzmOUhLgJ2Ev+URfbZyXKQ77/pkyaRjLyNTWtw9NDtL+FVfRgYgEB3D
SqXLpWILhFRRY9Wrs7lEYjAcam73ie5l8aq1jp7PHTujYSxh6qrTRLvpsrm3DQJL
FTNJfzYQ3DlYLki/Aeff4lpV5hG8RrUPWnG0RgfK2QUnbB4RXakU9O+HoDxWQWPZ
8gl09A0sy+jSJleS0vbc9HVR0lOmaQirMbJYL81PyCtbZxKZ6PcGrATdYP0fvceX
ZJ7SYXm8956PkHQPmlMF58qYzPfoc5E7qjLbxIyshv/hwTBqMPRXPkbbWzUfwrRl
NGbQSUgpkB8yAAN1M1/P9ZwnH8FZF3lbt3k7wb4PhSvUXeyCtKUWA3xEp4jUNRt3
9WPqn/jawiJGffHTVmb3KRLdD+k7lujb2AdFtUPHkLZMDEnwxDgOqJMfZz+VtXkc
0FE9GXs0pw9zl9aAEWjVD/EjRMcB25TSCGiHedPbA6Vhmqhp9JX+DcxHmWPcgmOX
sHPEbY4fc/pPSGl7DVu9GuaPdztPGKsXoDUjj1l9C82gnm4VQhG5b554wV+bKQAH
0bPQ8spbQpgjk1A5x2PFss6H6+BJ50ad5VH1WcELE/2zl108bXu87bND/J9nfhFa
pVUOPE8GKZvIZcJ2JxnhMRkWb9busooxwT9elvISbuCyLKCdAVLA5fof71SaInKr
LzPITRDyc9t8MmraAuck5K/GQ/fJe5sTMmfWINeiU7TaculNO7wpI11sxz+ot5LA
DHz/OHPHGODVqDE3+esESLvQJespaKP2guCosePwCT9sSl8e//Y43LYgMW8tlPne
u8cfBokv5Zhtr5/qxbObo56PnYpAWqdt9fJgyjmadwwLyWYAXP0K35XDNtmGdE+e
J9UUi7rgJnoGFSgMEx7jsg1cKquVHZhqsOTSepfkrVtwNETUXBB48/SPw4lEmX0e
T5GMHXFoC1v/kq4/Aw18oSNYl8c4IKA0leMWwV5xn4WVoreHZhHW1mwDNWbGA2cQ
2ya5GCJYxe0q9gwNX4tVYdNjdZQqSMZB6xR2YNnjlOALPCYknIMWwKFS0fpQkanB
68mnEJEYrS+s8MnxjF5FPFE35wu0GaZyNu7t5YvdFwMXwhW517CTXgrVqwFlvith
2I5GR4jLAnQ+Onzy6PrdE3nVr5DiBB7KPhqC1U3lzwKpCgwVvPcWlWVVepVVfqcE
DvGrMJTFL37zY6vhGKzzu9ed1xilcgLdL6jcC+uytR/NopXEx+VRorRrl7Aytqb7
zMa8BzSWvEi6+2jmySgYi5MzGYLNSedm0Akk1/tdsiQCyebkJwN/zrXeBm9qMwmj
J8YTgXMJMM1/e1ogg/J4IFw0yh283wn9EhL6GyOQ5+zgU6VF4QrZ71qBzEud9Bjt
XTn2A39CiA2+PvBD7UOwLj1wdSaHYSLAyA/pqEwPmEYM0eTA4WYUXCTmQ5RbM949
1stMte/PNyZBcXDnz/p3JewiKwRPvaKirBgrefaYkuZqlHdgMCMoA8dZAIGt242s
m/7yjVQJMeji8QgktVmIopPStx4fkLEu70hUEf5RSmu3+4s8zE+0MHcB9Gfkiy2x
99P7TnwxNmZhzB+M+JDFS7sSESs5x/Xl6+WRS/AriuL2DcjPaEcX3RYKl5Xhd2/u
tor48dIsB+LpmKDa0gY/+obBIJR7CGOZYbutWyBiBl4IZnatRTI3JEj5dhrOJDpp
WR06HK9IpXce0tiypYjFb+e7nHY6N4REzS8XBYnzl1AkUu+dXqfdDgZOrnt6XoEy
KF7cQXNPi1e0NJ/Vm/jdEbNiYgY3beRMFs6JUif8yaHAsChcbZjwhPwwQtCIy+TV
SRHxr9eCitYxBOC0z8+/CWdeHPLBUMNjbLNhpLdePSVKFD7O0hjeuE8Palin89BO
gyjrNErg5W5oMdahl5/u2y6p7Zp29IjHzVY5gWCR0ud0/Tb9tR0TYFp6awpvspW1
22qUx1gBemTQif04bnlIunKXp/X7+XOGYexNaAWO55DW/wO0Pl3FtZYEUA+buyKA
w7shkvKb3hLMlJZrl0BLaX+BDUqWcRCrNdJnXpjysfMLIysmrQRzNPCqai9Qh9+7
IKYeLo0HQzXDvAq9szEnzKCbiaeLev2pDTvv+5yPwgqph2lNA5esno8Zfxlig27n
UlpjINOO9n/YoQl0cZe0IUv0xQCJoX0CxfCS0wgSBQK+IES3ymaUfioC6CCn0cJP
ioScnxVkjST9qzjc4n2YZDPIfLioTENgvXFnWmyvUaPku4cQhSTNml2aeovrDtTy
ldFcZAAczPw9eCkpDoMGL69S2ZScOoPg3uQWc9a+YMDMVC1QyzRVtZw/hBmamXw6
ARfIdzNUYNf+BLTIAu6dh9dLQjMHdwic70V4jlW0zUa9SYnzWm+54R3Fjnke+BO9
eb+gm5xg43fWQXGOHD6jP0GiKyfqTAVS0GHSaHoXHD8W7s60eVs3xHtgMmj5ZkrI
XEf1NyQc7M4oDOBNqxwqHxZNHMbxl/580d79tw++34RUocWqhZ3YoWfhRmlDSTPY
VOGPuY6R6U8PaVxKsQxRShSvR6jfiM/aslYeldP28oKHQShha6yYVGDBJOKXMNUr
ltU1zP0HPIEppkgjadXUu2UBL1/QouYoK0Rtp16Q4bu6Ly5Rdo/wByVstuqVcDu/
sIQoKOvXj/cURiby5sO+OBTpwu5Ek/LKuvXh6ALGcgh/sBnctSxEv8uGiyV96bgG
mPaPm+6hf+zC4FPmHuJlFjq/xtqx+/xUHz3YIEXnZsxlOHssbQ793oE2LCkHET3r
7azHrqJh+0QjXbMaX3dZB7FxWakxJwaZgKHySQe6UegNMO3+Qx/9SSSR9CEj7Q/7
Bgu0FPf3Nt9RfAaevch+9Wj7nspcHq8kF2KJIX4l0jAN4A0a3OAQSFbIAH0oxJF3
Lk5t40qVnAHPeGYe/y8ilKbLn7ckQahL8a2JvEwlor5+u9NOl5BKblSxbgjk2/Tw
aDj7yWFx2MuZW4cqmtmdoKDdRHydIIY/8AgNI+UljiQnfRcifaTaQCd87trGsbxB
rcplBSPBcLEb2hxJkg1QxUzdqRnfCRAUN39X0UxYPGHXBUrID6xPXFiBqhYuoIAi
woKi29KG16rao/d3B/OJPt4kOhMnjFKqxOCCM9o8eU2UpJjRqShKSUwQlxWpanNL
5AZRV5Q/+ILHWUDOtetY4XrpcMz6xHT0PG3j46B1Ya7ExA3AP28PEVOzJ7O5CjPs
JtM7lfrpEYMWV68rwjOfZ18NhH2EiWBrCM4Ous6g1QZis1C54YdGXt7Q2g3wj8gY
CcVSjpDPHGp3rEX20KkLtjapO/B2i9IJUUi6IN/9LIPqOF9kn0gcDS1ImyFiKaAJ
ovGwyMQRFo9Zwg6BDmCUc5S/uU3KdRRJy+neTpQE/p07wz1pcsYdGBEONT19RAyy
RvDMI3zl7fzblBbipBdE5h1o8ohesioKqNhqFssfrLbc3V8atMiR0Ey+p2NigzRd
V4hbLv9p13PT6KZQf7cE1ulix3OrM/AX4AN9SyzdiFkXWrql9KsXzC68OFQ0nzSI
2/M/l6N1jdrD53xHRk8kyhOMk4ovwdJb2TDZmW3PZ1XfejrIYs0EIolCZpeQodxT
ewX8LzOq1Eo8e1yQEQO3/fmqH0ihjWQHnRjSVOnTBWnlMkwn/NKcx9pI621Wk3GU
Q2MEpFY8Uj/9n8xL0oikFNcoM3qjz4ijK4kwMXcCR7H0+lt4isMaN9/crFVZEgR8
1AvaPmHaI5y11Y2M963v7QpbViz8YkBZiMVKoS0sUKiPXFMoiVzTJI8m8vJHzE8k
hLiL+8JnqH7Ak4xi1WC3XZPZf1uRIS1iM28jKSf8by3sULCaiJvDlHk5A1xwkWob
JLATr56DzKAjySRhvwTynzVy934p1o030iL5TtfdIWqtLpgp/3qeUgcT9BIThBFn
Ljg5am0Zf2Gr3Q185WwZ3vGkISUEWW3YFq8A79yXqbwPcjHyenzvDeKrA1fTE8SB
tX78dMrMrEBluKrXSVYkMDirngq6sRS2jR6hj57/ozPJR9bvQM9dOKD/UPTBrCN8
AtiZpFUtHBENTUiG2BS7RNOgspR5TBOHYBrYyNxIQ2P+zUiaXbLI6BTKMiPi47RO
MntwDuJoJlY0Q/VxdY1k2zURNI8RpyDe05YAF9dw1hQTl6tmHdWqENtTaYoHf/oi
R/7Ibkj5+hf5BzmXyE7c6CRaDjj7WE4cUwsPEHBSsBPh9eoJbSQ6XBTUE5u0iG8c
BOuj3uupfgNU8HIPIjWb3JUHUHrfSu+yX493Oz46eoOruf74ycDwkg2T4LHS5n6e
xFt6iJc1uXVXYATz4E8Qv2NnddgTrh3m2wodx5eluJUKL78RxKFjXp+Vt630i55G
0o7qMOL1eIhaYNhYXfky/HhoKx9i/bmSkhAA6ncoPzzrn8UKr/aZGP/MXvAwEjbM
z7c9iTrlovYK4lnFrWWbiuPz+rDF8SxWMZzwzPhJafwj54I1stS3CYgKb1dY/Aac
kEEelMN8cM0ovxKWrACg9JPqtA7q7QbK8jrmTz78Q8bjNNES58m2hgu8nwEH6mrv
hdzY0WfBbh2rlqiWAKVZIr9MpS0II+Tc/gHEEJUMdBTbzpYD/XbTETdeUTXfSmEz
YHbl5JJy9PuN6Mq+mZPilWnGGoDkrKHjtqOS0692pbigspxaEz9gco5ILsTgne/D
2nN6+adqZwU4IRhixPI4kuds4FKpDZM01nDIuN46NxDuWndIAhu6Eb9YMdBXiHMH
0T7fcZqY9cS1PgEzQQ347KQYbVc4F7bMroiolTuFIzpRdwNP9HnaZNv+jPOVVWVF
vjl50DksfWcL27xwWnHvdz+P/qaPz64vTrAKpVvTeFyD2Rtw7MwjHq/GspDEM0L1
XO3ir1oSHfpqJH0Eo0dVVrRhU/HqL77ptkKdt4bIBiuE/DGbJeux7lR5vT9MX+nk
QRnb3KTDh6DOFOSjNlYDKnFzzGQmFVJoBCO2YPUN8no7/pYvOSM1D3WZ1DKHdWYy
cMLTNrUSGLelYosKcm+LULz2k34FjunHN0Zx9tMgxMkQlOIQJAyukXmDsTsvo19b
8+jLjy8nVfKAxvHlxCh4n2gH673xrKVhDEKX6XkMjdoQXSAsWmEVCgB+1rQEr9tC
TVaW7kPkccAsPVn+/uW8jg9GdEfsVMJfM5mbed2F2cDdDOTTd5H7RwpgZQPYzRe5
YcZiKA1MW2erfWoRCtf2OQohf5EyObi0RRZSl+icYLdBqFmftniqGmMdhPimyfr7
wi5I6s/tjI1Wk/DfFanbmwvSA9hyvRQS+HIxVPv9dyJgdAiaKLszHhlCTyyOQWDM
yL5qJIobawBOXcJEND+pTUK2iNMUNXrOBTf2fFH4Tp/6DzzV7qx8p1xqCLJ8NY/Y
XEVIPn6VkVrBk+OJfoSUgMEvoE6eifgKtzqrNaQhd1XOjkyPECnKGgf94rDcZN8t
9qtKrZ58eemWxg36YWMi9nPwkYouKyO4Knq1tnVQZEnzUVoIai2GFpDcW0kDncyX
tdD3n2QTBToNmk8VU/tRxSnJYy7EFvAbxFXg8Ql1Xe/EVEKOQKoe2xFnDcERLyT2
7GG2rPk2Fe/nXfPoqh4btdEz4qnYjGfIvCngBjKE9DIQLPHreRjDtjciXD5HBuTV
gAB0/sfASnUcdvH9aCjhTvXlRDSyx5iotN0eWaoaUV1ipM6SF+1FEvSpzYwSPLrG
aU0nZYm77/YPbhpsnugeQyfpvTrG252a1UEuRWV3ly6scDXCmF7mPJiY0oVh2Uuf
NdyDuY0Pr2CCnLSNy73q+5mmfXVUi1N6S6+zHjTGz53WPNJEOvqyCzY6MhBGhrMg
k4otoujT8ssmfQyz7sUDov4aqg8GTHqnpBu6qobiI2VoRxRqd38rXzeBy7I2KuuT
QDZOffze9ehkyGTZlzHBW9UA4jcuVeN+lnSvmWmuRa/jyJuqcJtqX3S4eqNSJzID
kK/9S287LresseEGBHrLCLyKmYlUydj6Aweb7cxgYWgj4kDsCkapTupWDo75+bvm
Zx9XEa0ssK2AiViWbigO3tS7CgZRUEusj/o1Iy2YlRrsKowe/IiZif5xU9xtnySN
7cQaLwLWo6GKMSSfrQAH0GjtviQcXyvAR56NRpbUI8pWNEm9d4Mn9pBRcIuMcwFV
E96v0Ax6uHuZ1R+Tqh79Oy7tWhOVejHdYkWCTZ0SU75xhbC6h0cf+ljs7qcTMnew
PTYP9RI34jTxmVy3Z/eNwSB3ymRNf6Ht9/bMIu1RbigfvDfijCZx/rquX34IKkad
tKUVwhB9bQh3Enkkk75sCZnSsje4NfC6y0aMwrafDUx2olFsuKnpNOYRsBZCpXsm
4o644V2e2sbtr2vmXEQEUPAQ66E7AZhZWLub6RtuQ1/Uh0E4i4YlkS3BC7yQRm30
oJwS2zUJ5yI5mD9k4p0QMVfV6gdgMwR+Ea++x/5ky9y5l6Jy1MHonGunMdnpWuUW
D9ik70wi2tJaWe+3p6SF3CUwji9AVyfG96af/FMlOK9zM0UYtYyS4qaiZq7dWch5
buoILm5rYE44hOczhgzziNfMAXDu1wr/GICf2zUx/HIPSGhE4KlEXq8WHHSbHcWm
8VHCUtBfRK8GBIIdxAcbFlTvaMOXEjH0P2GDIhp1V9YcDEKux6Z2GMOdOYxgXZch
Y5sCoXfNcSWlcNByCawGrXSUG10e3GARlwR9tJi+DooNi8XzpdZ2ZrtEvJo+Z2Qx
HjtKvaZx7pcaSirD2lFW4dA7QORwBx4xoMv9JXZ06mUeADFdRb3EyC45N7FHUt6J
tLJoQcdzCozGdwu2KhYVTQDsLN1WLrnoGuznGE9kltfiaCi+UCUMtff98tF3mkNW
x/ay7Ot5sCvAN9VfJHltmt9OJm9OYg/GvGy9L1JJtKKEVDNu4eFUOQJZgY36r5fx
r1MCupD59erQ/82ByOD38yx9bdRxo17PSIIgW/znaMqLfQinVAfZpu97OFcaviBj
EsdgVXcnOsC9EdverCsJvb08DZgoedNSYKJLYhbDmswNwMxSHMEpBAl2PC+cjFyf
tUmhnV/apbCYcE7RkQ4G9jLYhbCdC5QIWPEsAuLcidOgPI7IaSCOCjJP8Q/eTRY+
JXtgAxMIozqz7Ym2Dj08RWKtZmqyhTuPYAMFIYgW4BeIPhVv1BMFwVGJpk3Lwetf
5nteZxuIFHcLH9PnYtG5IE1+Z0DJAkfep9HVudKaUYJ7uyG5U6EoV+HaTQEvqATO
d+X8L01koVhV2Dmuo5l0wC2lb4LnNP8GD9AdHkhlGo10QZWdXAPWRRE0QQfswHKZ
yG22M7+LhhX/zUnRkEUsKL+cuELxEckb8KPAKgJLe9cvSSWhX6KNBgiZl85vPju8
gddcMs6Bh/5smNuPxcrPTMSzOHpQHYfrfhEbua6OiZHOvcqm4ZC2uwsGaHQrDGS1
K7VlPaIwV1NU+fViXu2s4YmwmRcOKuCQirG9YLrex6opm8hQMO6iZAsdf3Ax8iyf
FstQ/qkbS+sdUZA1sKQAigoSFwfu7CfG4bakm34Ocj+bJC9SPVkr6Qt/Mx0Me1l5
RPAxzMteX+R1KTVzqROILSbhLkT5IqfMU5WwDkxBikXyZcI2QMMoZ4tHXpVXTP60
HTk7scR1uI1eR4NQnk0F+fA6OBkuagDm16dOP4REJqzeCn4z2NtUMHpbJasGYTNn
nIZg4t0CdC5D/K/P31I3B2GC4HbTZLNOzP/27i5svSc29MZMlcV0wToxxZbdcYEQ
Od+C0BdX/5W3Y93Ro5emqbo/GL5u1blsxL5QeHUV+rkjXcrk400r3AB3gp9Nhphw
Tqi7i6gIk97EYhC5Y+/TW3sbEbsoBlLBqLEkbn4fROC57H1/GU0q3bux6EjX1130
u1Ppawl49BgYRzuH09IjhFEdJstRp2eEp4SN6bfE2p30EaVp+e/eDUVTxvEb4Mai
1flk8q8sa+iPiJxENKs5bMCzeuI8ZTkRe3uwev02ilXNy0G0KHOV2C2cQTTiJPKN
LghJ8j01AmiRIQXyrkKGDWcXH+Sx62ky5iKXIKViwj8vPGbQdHAW6Ln8nAFvuQ4R
qquqkRcN8PD1tp8N/CJbbfGz2aPPV9G3CMWfunpTGmrK6+s7++biFQei1POTet1t
eUpRSERCQw+nRg1rLRz6HgvJokJ52nbEmzpy+CVlnIfgOiAlfH0zTMgiOOSklBN+
RD38GxawICjUpF0hAcl3fH0ANwxGtJ5dZzVZR/qP7msH6UHory5uBsaAMcSy8ebV
5X3AjF1SrUuWth+wYEwatAgV8ocGLJ3RzhhxM570dIohAHj9vCmH9ZnBa9cvkfsL
m2SKno0ki2wLlxHA/z/9Uye/wvlE6dC/PJ8JPRBaUIn/ezXY1XDcfT9BPBvsIlmW
OvtpQHEC38D4PMRLYKeWSI+l7P92wGciVIRLxAehJTNFZJ3VszD3XlZcYLSHDquO
YW7Tl4xmuTM3n3JX6tGNvUfxqKN7xY/AWZ3dIV1rNB0ODIaU8GgueiWgo3BsQ0T0
f4sb0BL64eHBza4ciZ7p5ASXrIfrGjTjFJO/FgePTvtZ3zIljGsF6ClxVaAbaAZc
WVbfSpYcJgnm13Uw1lvax7XS+geAPbzZXyhaETXznEIEkntfhNKsUaQgC44ixvj/
rS17BPq/EN6DZNdr5GbNdXdt0s9CcxnoKeXwMe2GMVGp2KQ98v0W9PCjhvJGbqG4
NRmXC+QDUT6zqzrQDnzkNTcJIp1zT+UnwxzAq0ieXBjIgxs4nbVyuoDY/jpYN71S
iej8V8teTHGBBLOTaCSdncT7gfCWvWp7q3wXZQkuTrFkqbkW6AGs1qwLoR2DTEkE
VUhLU2xXdT24vaG4iMMD2PNbpv1GSDyEn1av1W38ei4RBvLGqvWws1IuWDb8qAnP
MBOjnQW6gyI73gmuy6cVL/W9XTMilOzUg1uJXFVSlyTqE0xAEx97FJS8JCJ+42r/
Jf4D//ViBrwDDcKaxpMFjpVcxrCeqxuKCkP7XqaWSzmWtui/FCn4XcdItSIF3D0Y
LU4x6/JS9KwPL1GoLCIn4nM+jGFJaPkq+kWCosGaOjMzU1ls6NDlgBiMyZxsCEcf
0T1jLg+qFC5WoYcWJ7vOaw4sU2eDLNCh7973nanweb9l/IMNDnbRvvqH9o6fWUYY
glS9byuCYkqmWlZOlbrrIH39qfCV+/BEyjTzPwhCsjJOoScPMKNl1p4JQi8Gkv86
l/1WoNqeIjSRDXuV+JQzZcdg+8f9L0nNXnqUT5RPVkyU38z6nUaZwPhKRWeqNvKW
yuomQc+VufMeOn131kYk18HdYePe2mmkSX+HLcZQqgLj7Md9sitgEkr/TjCXk3DZ
pLMHeP+q82NSzLOfwRgoPtZgjvHWzMi+K4EGLkJipXpPrkoVs7kT458P0r/2iV4n
JZiUQoNyODayRB7bFT81Sp0CarkrcDvpn1Dcnlpjng44KVVjMYm1gEo5lxInneUx
X+wovXjhmT9Aj2b4dpYx2FmNvMsJuv/Gdyk6dxeuTFVzRb2+mqDTd3q0gvdgsujY
0j7tHAh9soh+Bb/Gt7KL/NxdX1Z0jCmv72w/BvArMofiB4JpSpZXt+403EHpJR0Z
g0Tpx2Wre1crwXqDBoWkWbqh9LbLl9MuRaz7qc/FY/W2cfzC/08cBubCyhQstF6+
HSZp55x1gukctGPq1piBS3pQ5CCmu2U8tVfH5e/51PeiK9oXtrWXnWmCifkFSVm6
m0DQcQUbEwbxBVmixHTh23tJrK8qPEY8SrsSn61pDAjPdMEQERWF6+3DQ1joCLny
N5QonLSJ1yVYusUJMsiN9IiOin5GNrhFg7pPUUi4xxzYJN6wSBLDrYHiymaBGTd4
t6Pc3EBqSLw7tU8kQ6D8ZJGM3T8v2aQ9wqE+r276fz5mNylkfQaGgLBYNxKbY+xl
58rGaq86P0eKO69ft0GEqfuRaD2BbpeVimiojpJ6iiJUEULYrrOWmDpfPUFY/d/0
UZJbmxObIuwrD+a5yPNpMFlV3eZ6i1/Cv4Sj+IPPxWOFV7evV+yccVj4DDanB9Pq
shPb5MpmCZ//KDg7dAT+hfqYg4BVXiTW0NIP1QFORZ5hW1LgQ6lLIu/FEWrngrHD
0lnAchB6rC9zEhY4ptpuqsC0/hAolIaJIlTqzbrSoCiS9WIpu0dOBxyi1lOkRYJh
JHOe367TlQgfVzaPfzNbxACJv4oUJ94zbaaVGpotf/qGxjsnR/e93KLiaSg6/5LB
cGmApk8Rf52NfakOAhkHiLlODHHD/JGJ1UbZLy7qaHo2SgfL0Wm43LBZSa8xccqG
2pijw1BKq5AqV1NXLYtAvQ43VFdFDMHWwkpBGMDjXeAm574tb0Ii51/jD2s/Qi2V
lA5pcXmZ6YoJ/HmlGtG9vwYPvo4X7/pqiGjlJ9PZwKt0noFN0Ht3omlDaK06z9+6
NFdUNU2ayMp1gYkjEfYIP+hYzC277kPhtyVafZ00O55s+UevLiitDTM32a3nUjGM
4PdAZezyWr3Si3vVQN2DaLTe0P96UViJDnV5ZSnb1sQxC9K7f9S365guV/Df0v8T
gldlIG/gze2VlVHNYt65Vgs9YQFqiIsdmSDyo6cSUjd4K4eWhrAbJPCco9Ebx9kJ
QGvzZyteamAB99Pw9SmHwr80nqrHp7vVQR2/U3h5o5vCEpNYs82O5h809ommuJBD
D79W6PIzxTB4Vx4E8WvcMS/uGn4F5Qk6kXIY30vG2c/4fo7rXlXYZXqKEy9izzW9
F0ztWr18cW6xQoN928e6ufAfIvEKdWcz/sAODxawMmzBN5BYJygD4gjXdTy1ZLX+
1vy/ocq9fUrMljKU62j0RA6qOx1j8IrLS7hujgWkPYw95XJzaP+a7GY38ml/nC+k
2L/BKpBAIj9AqskgoOONRzXPw5gwAKV5u4NIKcEPFhDiEnWSSnDXX0aPKOb1Eg9R
AxAOtHXyurPZME9sUAXOmYOWodras2plzFNrneYzgBEFiF+5TwGFxSLVfrAKKgap
OBKOLbkhoFASfIBKLZIfZl5HICm39/4c2tg4tEyZJzqjrMkvgLyI/CwmvpzePeR1
gGKYZmTfglh1TULDYg1xmEVEjslS44Jy40uFePfYWcNir8OXNs3tvysoH6YHKIz/
08022JWIh6dUGcZ4aQpANz0kZ0hlEwUSBFTEzRJRgPeS4KGBnhPwpwTShvW3x703
xZASMmdemqNczDbiigLeGX1kzESXlw/i1w/di5hdq0QnRiz1xE219bLuOr6a6RtR
mRSHQrerbXVOnPiYpo8N6zpG8+Ncm0b4MDeUROsQBOEpHgvne3MoCPxkv6yHoh0a
66gyjb40K22Qi4dzUIdwlpy/hEPMdm2Xo1kxCu1qsi4FEZGjvOQq86kOBRcdIwKt
PE3BhrHwWoYCT/Om/214M4a4vD3Et8WBUxncvtizKSYE0IUL/Q3kU4TgwswuqHH4
F2IpAc9NVtql2Kt/rWKJwxmSH9Xu+5ivE+RW6a6cY4roaAtWQaB3ecO9P7PaLnKG
m3oDr8Dw1W6ytN5Q4GaILstXnSc0bNWNqJCbaiAgTCn5KFaBa3AdtaHn5OJMb19K
IfR8QKgmx3MM6vAYZ07Y2bI9xAN+wtLGDoTrTB87Il/3vlcbsAnDjkZy3PsQSsdL
ekDEBms9tsNl9s50gYlxGwpMR7+ipfHFC6xITJye1ujNNvGmUH+3HLpoTuNFN3bE
XjrZfD+YyKQti7U88arwuKU94vszhf0cXrKEpyTENeoAm0fzRNiwU1ctHHAvesl4
vzKZqE/RdvMuBotXMOio8gmwJDQTxi8RWOJuSuDPufxSfpsu6BUUOi4pHAL6myEX
QPI+LYLJHNXrIQg0/BtSj40okNQYSHwUOxIHNxpwDqZX9E3rddrQdQ9e5ZT7UejB
lNWTtV5VvVkghOmBDWCSUmwwtTm6QEdeKOQqh2w0cJ7/nzz23tZlGFd8kEHzec/0
3eECu0d6ddsnKJMFvONx5esR6XOqUm66mmNWwVfxloq89c0iqVhnQH4g7BIExMuX
MkJgCgY9b76g6z8jKIubBM5kvK4oC14nfAoVT629qnTxr+bvgzyh3NI4sAWczsIJ
5LVq/vl6Gzl37itA1ql1SfF3aIlsGVlGqMM1H2hl1ieB302TE7GmcEbG0bIhNhwG
qntXUI4Pbt3Zqqpe1hcOmf/uLJP7+0eII4KHopfkiHD9cLGbzW14+6XuteY01gFQ
89rpi5lyup8ffbWBVE5+u6Vj9vvqqgwwaDSr9XJziQmZyOgrsgO5D/uA89EK/SUO
eJZmmj/Ukx3PVKubCPpCV41rEqY0r2PYvj4XGfSrBvbfFgPTF4w4q+Foq+cgDe2e
PR6rxP3xoGQqG7MlXWjVunVbAgoT+ALeD4VjAWPYjLNvINIPj8M4TIbbKQrpRGhB
4K9mAa4vT4jtery35iPRdoozM/zQdgKHB7rMKF0FpNxSFoQipfe9jkvQW2PlIyBw
HYvOjRSpiKarP2Kg9QLUt880qlKd067LEYAPSfgEL+d9nuzbQZInIvsIgP7bkk6+
oLLnavb0uPdd1w4QoRqLc3/WPpEtfRHuYKa3SCXZ0A4W/3kphjr0YYTz6JE2xZds
8KLF3AJQjruRjDbQqE42Xt/H1TiQY9u7NnofmQuOjmljN1ryZHOvY3ao1K962SDG
oIiXFB5Zr3q6xl2jqiNHKxboDPZzha10Talo1ul1hpelwil5ioAzheqvwqKsg3+A
jZZamDd2ZpalUruqsTj56vuRO0bjgUJhwGwAo9M0P15yTk5t5a+wQe1F25fqK1Dm
O7hLObYXNi9gw/PJa9wyE7A4su/s3jSWevbiN81NEftPhe85svyRaMMymbiboajL
DohdtIfC87lLXf9x7nLpWv90sGjSPHbcTPu3IzSb67MFBxYG6UkQaF4BwOHeL3t9
T+J9ptAeS/M/DLxTYknUIxl+7xK+FiCBvZEuE3iKBt6wHmIdI6MdIQYEzMk8EziP
J7qqfrseFPygWjjeO2to0LXPUq/bwImh/i3WUarDRgmJoR0+SITfcwiocWOH1Lv+
q6yOjkBKzhf6PArGXbyZokzMBbLKp3X3HGsGjoSydVoNCmKvvXhtQuwqkm2SVmek
PmKUg3xvnShs9qXSzr+f2hh+keqV8/X8lZIG8eujq76SGrLB5mniSX4fm/qrcQ6y
+Qv9K5pSSL4kPKbeKVO5UMWLWIWlhurzaKqWfwWt3+uL34imdWKARmr/JL7K26WS
yUQOcNESZYlcbdq0UdDupL56yO9EDeJzGrj/6p5JceTjywXp9vCmHLNmmcIyGe1E
D0SUGK3o4maHtRcLGcUjKyX50fssrg2aVHrtHzRnjolVuauhQ8K+Kn8P2jz/jfGE
9oblMT+ZV+SllA9cyX+EauTvUVI2lwRa6W4JryViwrXCB7wXX76kqV1e/ALiEEiN
O5tEsRaQ1Y7NSS6cjYN2OGxNN40ZRr8ok4ktmIDT4HgcJNnkVajXVhyUE28OsLu9
2E+nCwgj0307cJkCwypB+x9moDkGVJArM2RLEAI5hvoZ2rhGh+nvshTKQ6DMlt3q
ZkqkqrJBqEXtikyD2qo1xMBYYY3wNB8zxSc7Bng9jBr39Mai0kmpF5N2BZso5aXZ
bv5V8gahAcVHfUKuBwgDXyHktIUff8l5iCIZ5iXvIRVJSWeZ4y6OrEFq6gCf4Pp7
Q8vmF6YNKT+s5gPVW8h/5mZgbpe95pEVcLoKhxItyao3edNifVxASkVeZui755Le
lCF1ZONEf9+Gu4QtdKW4Bwm99YGtVKHF37KfYxCOkZMWwUrMvbzQwsYCyIuImIGh
JYleF5u/FP6/Vksi19V5GJ8urDyWnYrEdb8UNoH/ZLwmGozOZspKAgCEYRcfAS65
B4pQwODbwjKlSdfRuZbLB9PMtx5txQO00JCcYN1UtNfNWtrc6OrSiBBGAaeG26QF
2702EPC7sDW7C+LAwiPcu7RhE2l8hOMFxBvKX63T2eC7exzvSVv8h+H5PZVOwuiS
5opCYhMtdec0P8H6lO8YER0bcjsfXk0DvSIpXT6tbC3uz9CaHrU5Lq7S94KJgKcu
68AzzNWNk1bw1s7JTE6NOQhTckZ6YPVkyKL6RKxqcy1EJ87dbMEAoWgPVxRDWxh/
Ijj9n3i4lOIL5O7S9AtGRLCThGkPkxwia3P5lErtgugSKevkIStyXILRjkAXrc1M
9845IDYZX1MpmFBuGZRwa8T8MJUuD466/xw30Uzky7pBjQjFUdsOtUToznufi/zT
3FYXcgGIlGxl837YdHyFuEz/3t9GudNWU6jIWbppP0awRYe1iiphZZMkmDwC7CWA
ZsZj2Rl3ssz56UxOo8OQ33qoKwu7VOmMWbvV7rrZ3FijHQRmOqeODkdiUhNoEaBG
SHok8HV7kx6qXS89VMhnslpnPPLMpKQKuQrVkv7mYgQfFQefh/IhJxuGeQ7ONWqQ
rt1CFIQpxekhtbDbC6xkT4+DnitVrEP8km/jg67Zu8zwwUWwSJ4ZdvDkYLsfk167
/FBq+UZyqtij56cDGEhTwRxapDNWtGY2Is/K7StjYwnFXUxIc1fDHZuv+SBou6zh
f0PS/BHpelOLA2fJs1iDVHgFuJDufRoXzjh9hXxlnz+KGm41Ydaj8TcE5bls2vtA
4ORFZLt0ekDrrBfsk1a9/dRYUeUm9iQiu/TEmFr0nI74BM4VQ48LzEkx7vrskOq8
XyrS5gWaIYAngPELC56AJyP2EHaojXh1zcjo2+9eHVmAGXKtbx7JQm0n+9wurnZ1
KDkapbGfAU6f9m+ObBrIVrE2dieRvnL+UVblFpz57DazgAHthK8eGFftsN1Mr8FM
IvzpHFBo9Wqkn8/q6ozhyY6Jw8iKZ5+LqWhbzZLXla4FmuFzBOOm5HVwxnuD/e50
Z/uldi44SUWDSV3etvKgYYeQtIYWZ2tMnRyUybt5k3whW1HIPCXd1Ra/yePB2hyW
qnEnJTT/rBnZHsrz9+CpN0kN99Sh8i2TQkVIeO1vtvOnaOuxJc1PvZt5nlpu1gq8
loNksehTqxEy0fFCv2/KHqSHFGQ/hYCKtSUc1wqJXNWt4d3qa5UeRO7Vbxhop91o
NbDFeBMU2TwSjjUjUkfBdIC5/spp8n09Gza1zRAjn0pPHipNVE+8gZCJkiVzynK7
yfzcQcaCw7+pZtA5inL1DDEISGAXtNTYTtwmdoEDlG2KLslpth02H4Xal+UKVNI0
mXvzJ5Gaq6uHCIvq6Mjq0TZUAj6hbQPTPdztm/pATZouiV1fJQ79heHUBEtmu3fD
C8maTIJY/mqHIle2/U69vvYdToNfZx6C7UPW2P4INAcRLM6UdYV8HaZwSITwErLH
tXgxFk4EMoTeFXJWTtyT+fxRnnQr0VWwFnJWJsgaEE0UvkowjuoeK3aUQrrnBo8y
1rbYIQOHHY7Oegg2AamCEYRWD7iTT4Y4vWXJ6+YxcBkFf7dxAWBB9Z8YM/yC8+ZM
XNMucNrI3DdmgFqjaQGpnA6c4H7VWbMjxi4BXX2oma7UseuCmbq6jb7rAMPQq3LY
dM0EJwUNdqF8SsweobbfrjjznF3wYMf+hd0iggBCjSCKlooBuRpsj2l3fi/yCxa2
mnqHRjw5H8XLLRhBbgrcEqw6bykbjzDf7rHtFSLQ6BgUpUok8Qjwmy2FQNxc/62I
jpWiKkwbEGQXQBSRvi8amlZxQIMitUyfyenNSuMdjCpzuneFtoUlK8PkU90wcs/7
HdD/tpa04T7SxvfgdfcSVhYMXZWoRwDiA6LkX5Y32Mdd+xYFBBUoDvATIrBhPZbn
U6O4pbxJRuw5Yit5WwzVQ1ncnQovdnvb+g3ytuBGzTWv/C1TvzHH5wYw8C7VTbfu
hvuIIEVUiqABJPjHTY0uAMkIbn8FKwSz5m6LPLHKtj2ic7m95D8W+DluzeXfrppa
IYSb0UM5+oRulPpzobFcniCkmmddlige05k8GXBki+czg4iePiy4u818sk8rNR01
semMCxLFAwssM5Lf0jwrDC+YABg/CGHis8iKRHxSDtl2LAN3yV2jgc4vqcDJ7Grf
w7aqHmMUECrrVjH8zmbB888eZTH/CUvMXPf3F5ZLIZr3GUQadZplg4M2dSLBGg5o
sbS8vrrCYkodCrfMdAHPsRZdOdQrLvNPXkpfhTVWEvytAlW2O4b7IizvUv+IIHmV
Nfd4oXhVoYx75Z9fDTHboYdC3m8rBT26HuwY3TWB4ycPFwJIxOiFvh9xWhfc3Fh/
bQeqJwuND2v9QNlndJIWIAzqX1m0xwkjkZpd3haJTTpL6v8/V1X6zvEBx9q1832U
15drhPFZyCdNYEpqvqRihvELh/HkHdftLFgJERj85aU347hCnpzYBF44p6m4iJUw
ZJ0ORQR5wVL2OzN7I1DlzfUcbOaFUk3KDSpmKfJ9d8cWTh8YVHV7c4YQaG5nsC/Z
3ohGDsUMK7FWIv2earQBSbYkRfvcVZAwHL707kHzDQ/w3DodqOYhdLvQFqYqovED
efrzN5RDtZEbU9UOwvOAqjJNjuHXVIBfA1bOqb1q9w9QoGtCcOr6oOvzv9ZmhSEo
xCldc+HxlbZ5Zvo6h2A/W3l0ZGjBSQOaOeBgEZJff92zwG47CUPP6CpnAF7cAXvl
LgIYZJysxVSlKj0Ifx4WmAIXXfV+EHBRL9SFO8y0kfaFyVbbFOHsEc/TiBGr4kvQ
7QKDA8n2RJMM5XsHW6T8b8G8RfiO+GXMxYX9OFqyA+XNnWSlKxGCpnGZaU6zKs9Y
zPL8epUOkdwFV/T5o0Z5tpQ61SNhKAdAqDCYZM/pGV3TSRStyJnp94GxzBzauT74
U83XIZ/Wf7m6mVdyUC0Uis1C4o8W+RjahR//UUB1ka3x5B8+BVwgQ317Na1Jr35u
PZAQLA4V/PrsQSlQTGWLTJryhY6zBt61bGSkgvjPaOo2zF3Jh570MF/BB6Jn+FJD
mA7uPrzR1Dh5eGLWAY0YmRR26yuIwE89BiqdzmAMAr3CQFWgEyX3js+kzN67DnOM
f4WEus6uzc7YyUnToVBcfG3Ctyy5CRXUfb5WMnLhMqs5I/qY8PQFZ1a/MTUKl6cq
qxIRu/9VtUlqc4/2IJi73tg0F+D7ggN/R66hqN09LtTqo1qZWT9r/Ipp4opdI9a7
Sgi/56toPEfi2DMIfF/3Dm8x4sBs9TLfChZfKCNDFFxTsDXk6RaqWQqWyYPmF4n6
lvQxjC1vB0+YuEhbr23efjcCj0Q+sN6gHVCbDCMzW5Wb2KLAtru41mn+sxEy5D24
pDBh3sU0I9iH1BBWFp9PPMvW8WK9KznKJKd0lpbNjD2ZSfh5+bqCrI84qibsVamh
8Jbw+M5gSqX5Wc+EBbmHpb9qPu7KybgPz0GI2IBJWvebnuoUdcL1FUCeq3Ki/161
3hW6a2As6zvFO/vpz5SB9Y2mlGEopL2Abn5ThgvjDPjGoFauwHOHtwhDqG8CXvXR
EXqw4nfGh+el0MLoWkk1RfxLVi6WAE/0iwYxSlbGXj1kfDfNut8vHjdN60k4eq0r
NvJavySVLRgOuX4uBjL3cNBeA3FxDHweXrKOLJx0lv+1B/Sep62YXBxnnTj38GH4
h1tc1WyxXWlnrfGe+x1k37l6asr/0tI8SuPu103RvMilsA3b+HnyL/FArKfkgVmd
T5tK2GYXJFkUuMRMBQvw0I/d9HKtqz8vFuuI/jCji4FdUoaTvNQNS1gJeh7YxojD
7FClH9NhMjTr6XkQEwEyZ/gXUrWQviquttyqiJgU/8T+BYQ2xst1bvxdMQ//LU56
uDifofd4ohj7LEl2YmtfciHHIdVm5u07ba1QG29yERcAhRaaTkviUvjpgy+QgLMI
1jHmIoiclDpe9lR9PJHHaBCU+upTmv/r4xia4SHcjYY1Hhw6yQmiJ3h6ZRYFRuHk
WDvz+y5B8xQ+xAqm1iWVE+dHH0eMN3tH1X9Srxhx0VRfFHzOwYb84ThbLKMLVrA1
2UUN41FAb+ICLH9xPUTSePv+7a9a9RzIRHaOXm49HGDBXJ3FoY1K5DDMs0VyNkoq
q0WJmldJZVEFiY6kE7T+4ZM5FjqHnadUB73fscx7Wh41NmrL34fNfMKuPp078SnV
chNYpYCuMU3Ev8X5O/c2RXuSQypC6NvK6jQTwWaub0j3B9C2Kydjca4r4/OwAQXs
qy2y51mHwospAy7oki2ybMwQNjJH3wyntDkVSsKVwh5UdhO4ks1NfhnhYolYtGda
ieIx2bfUvlqluG9oxzN+nWT6PygSFHz9MO54DoUDEqy0Vz7XAL7RcAuHA2QCYyeG
vnBgsXA527leS3te0PWXQupvQv5HcsXgZEVgFeA7N6g//GArcssL1xxPuihu+C7e
hLeeQP9I7RI5ujVdvgdpQAru/FZkAjffYCzvv3RSbLrs9j01TD3H/XbfBJ1gb6r0
zEIR8uLp3Bp4WzinH8fIzHkOdjWeW9fmYkkqewxCGYgdYoJTzYqejLBv/FAw5t57
9qSuRCCEdpkoTS+iWVPyj+y8bdeUzDLZu4w1oBsduA2oOppeeeSI0s4DMjp/I5t3
19sMnP5iDmOY3llUzuZyf3dINCLVSDkwHn+PecZNCwjnN8J1tnG0dVbbU+3dY6ez
7tcFrvc3xsiKcdAw/zvkDgiQnPZEfwzJHCG7ZgvntKSgV9bxtfPHNxxLugVu7zS3
5DqKSKyiXAsMZ7cb5RNgPwZhQGQZp//rlgyUJ0rYyTlBZ60yBD2ozGI6OImFQKDa
eIKGxlE8lHwDT63Ib+i+EIHcXO2ePBFaK3gCwae7Moe9rVe5phfs9y2agkCFXjfH
ptgr+B6+IkoRZz3ObGpJ4uA/daOcb8l0MAP1ACjcOCsXaev2x7yLQ8L7SYrAk6Oy
tgFo4Y72ik41CvNzm/zOjQAy08aAz1V5AHTc3bMLpvNo+ihM4oIQAulgQhCZBi4M
6t2mhF9sUQKruQqoCMWOIie2TBYgL1/HSF8DLr/C9sLD2mzH6dmXe0fY0EaHGmfY
PiIcoN23K4BM5cNZQFWtKBzcp881AFizbnaqKTrOaPbL/WODtuk2FyvB9cKrJljY
othU/o4o5FJiubtZbzlkxa/u6Ja5rZBxcLJ/loqC9Y3R/d6xk/11/wXgiBB+ktoJ
XfLZ8cgph8ejg1uQFB/l7nmxrBEdhSkEL5zSfiKeJrtP50kiI51aafZMlzSg4ion
BLtSkGCMoopHnjNeJX9uyk1kQru6JHz5+jhY6naBjltKfdz5RT7nTFqRV/wQ/reB
y/AEvYGsTvRNhZWkmnmEQDRC/85tQVOf0LlHhms47c+Zt/Uhclzx/EyRnk/9YNTw
g1jnchSZ+Hlv/0OOMuuU7ZTb4abI6b1O2HdvM/z+m9Ld5A1SPmx5N0Zl7zkirsW7
QF9DjKhYV+h2hCHf1x0e9/ZN9E1qarzAOU1aoeSVpQ8DRlgtWMXIOdNgI6zxXIiN
w0CCZd1HmullC/qAko7RSs5UEmN6s5N32iuov0/BGoaYQyE3x8dhq9VIzWLDtf6S
5a03VOBaOf6Wu3V8zZvSSJpwJaVAVYi7hDvRYo9N6HxqGAoESnYklO2pkGKx7Zy8
sr84QSsyx8Vk8yvWVh4C0snPfGndTgRnKdGioZ86d2t7hqPRCnbVykvCtRfJRd5F
F2aCFrLlSCUzrgCnGQygjst4OSovfAGxCUQzYc6rDf3ZeHfHE79SxqkFfkL2JRmu
IpWxlV4/0EzHFoQqruT/ZgCE0t4jkrvtKxqzP/enyzHQYGOiJdX8lnbVvI8r4XW0
mjNfayg9gu8gnJV8VyO3rov4/KfvF2CM00marqTWseO5fdyhU44N3XlzOm2Bo5Rj
rf2jfZAV2F3IkhrMLWjpnEp1d8YvyjOK7nEc9qw1r9k652O67G0riz6KO842hQnN
EFHHRmPNz/ULH0V89uiEP5UUo5PP8dxUIOvW0AFLg6gJxsj+cmWqCZZWF+X2FDWX
tqJYMQueRHcwurs1pugj2qaNpp+Hk6072hNcSwugb95LUin9k24pGcsW3AYcS55n
ni9Q5MLjE80T3+0bKP9RGNsHHCihySpooq7I4xO4qDWiRTTo5r67062iYJcC8b7s
19oWiznl/5UPsQTIPRCZ88MnAUb3DFz75IEHdsell9P3SOiinjpn/8Eix3A7dWrd
Mbaa5ef+yk0DYolU2q9bboSAkzvPwp6rD4Gb1i1ZLhOfrkDNlsTuEEwEpx7UBdgj
RUyiiH2wZfOh0M5x2Zg5409hYAQJHgZbD+kuaiDGhr34KLwnZlytwO9FWmgFbjUK
uLXfFXkhXoJdfR952DwcFJTmuVKRJYDlxQd2tzAGi6ULb+bKm6zE0Gi5MImS+4lm
FgeoMeMLO2r+v9Emf2HY3573IqkK14/70B40xyXs5lfa7GB5ZhrvK9vp1DONnJrO
p2wEY3mSE7IXzwFbhF7xbIZzs5AHfgdw0GXbTHQf7W20VkhlGrv8E3aMFL/fPpmj
0wPYEMUMngscK4g0Ovtllx5IhsIZc3mEoLgeLgQHEEWm7LkQP7DBq9uue0dgEYDY
rGeY/7u8AKMHYc8AZu5ITA9UoGCCpDg6fFVZyupESjMG/FSsyKZgDcpkQigkE071
ZcGbzITvfGTMFzfzPS92PuPmkmXRMq7A/SDKxE6sZpbueJe4I4+tPBDvA7cPXLQG
NCAObaxKI9BN3rBTdB+0Oezsiq9HjyWSj9/taZ88n7EQPwVPWAF/6B0NDf+zPJhh
213QqW9SOAUfHWnuWuZm8SzpaSzYAWWAORAQm1oTXrcjTb3VOV64G2vY8G8K1tRs
U4mhAJMASxoyez7YsE9FwhuB0iNjPL78Pbexn8A9WgbctP793IapeeQEMqa7cyFf
nkCBwBbvAneKLm4SmASJVsIH/t6B1YxukEe2yiMwctBIb7y3IJN/g7Oqfm30LSS9
sqZ59vhy4zt7f708+M12YhRFqSCDzVE/WkuMoJRpiqzP1k+ufBc0FxyaJKxTn7M9
diVJ1n5EQZwSjN7yUT9Mdbe+yS/NJVCOCUm88tBjf+EDyZzj6efNbZJ6k7Up+qvL
sDUTYU1EkYrNFHEf8gGsd/tJMnZB5z4n56FEjTDbZA7c0iHlBNRPGINAIWiHDRtq
cQFBbFGN2006cYQqNyoFm5A/n6jOkmdFaTKOuZZDFRp/k8Lqh0PVaSE0+KJOBwuR
NDnBxzgok1pHstUSdJeiPepztKCg/HoZioRVmtYWxplMcanRwMbcXtyxD9InMtAZ
EMd5Z6vFUDLS3bHHFbrLVE/VAeN7QWP3wJkHIX8AS/TKkUIwHd0UsTc7irrbBNam
0kGqJPjgrCdWWvhcZr8YeuWl6dc5S1iUhlfK6H8Q1RqlaL3uZ4KnnIeGIcjYGHNu
20JhqTedKcijhsIOcBg49uoFxDs/472z5kg6xCkjD+/2kby2khF83SAxkVNhlw8V
qGr8/3noigsvxZ7sWFiuJ5Ofjo7vv+0+Ac/JcN+xme5d1ijrFv1MSg3wRdCmI44o
MxxZnXYiAFYfHFmgpCuRIMj9XwaBbFjT63x8qiWsYopmeBcv8snBxInMonrRiVTf
5OUZlbdLCk3pUFCKzQC4hNyJjrYjexxnfzi3AnO+yA/8dzwsUa4hqw2qGh+R48xi
q9NlXTVrtnSl4s0HrRD/jS0d1JbszjvHCK+e+Cb+mox+aAKkqxxZds0I/Dh+Y5vS
mKrrOXVUKcgyN7CPapimWiWl+6oqZFIosViGWMJ4hGY/Cd18JTiRNYnQ0dDCuMyU
WPtgOzySlnmAiJUFMXwKbzugLofwUSZ4I+GgkWkjzU1U+fw4BPSzcDVhd1CgYdpd
SKg/RTmxK6Y1mRslk8T+/NXuEsORRZKvUMNMpPwogBRTDf/kFiMKHwjT6tDPGQUv
ZrE+9CK/qd2CgJEeWVVYkl42l+Xkez6Us0efyKiy99+z+sxw3H+djRzaxA3cL7a6
EeiO/ZazoRzHaEdyb+UqJzBVNrp28zGxe0Uh3cVQRlIy+FlUDXuVoUmS/2HVaKY9
vyNfK4ORCbzqENuLMZoTnHarLpOI6nlF5AkrBxlVZ3oGmuq6hvNdRsSoPlkg8EJ6
ZyyEANtnIVkPSntwKnrmAj2Wpu7DQBOzM27EMgrSa0NFBTIRkaDQNZoyX506j9by
AQZxMfhaI9SXa0rj9QuMUNkqlJF0KVF6ItvR80/fKc0OvhfXhrJQdHDOSp9Dm/ZB
3Wzy/RlcrHgs17gjLpEGE0YOILriCXA8Ungnuw3I3YaUDEfR9ytp+HbX5aSzgL1Q
+EX0t94DZbXCVMnxia8BIMKbR3ou+UVXqG6SD/fC0hZkKWVGKdVMYAAf1XyjbkNI
VAUbCeY+cHKv1BoB45msvhL4hBsTEY9pBv0GD3aVFFLorv2J99LSXQ1AZYLOcJin
An27D3RUdqbo0QGGt1jFZevhql1pt9NVfyQqu36C5zx00kDcQRhE9l1LWcC4Uj/W
D6T6GhlCFsjsVbiKBSKhNk+2nGX+/4HQ9cuKlhHRbU+/xi75kQ3zcVXN2Jk26eOb
9J/Se87N2DCy9VN6NhfpP6D4iaJwf3GaJkyF/AbzA/V6PbRM1EHx7TZCtFAB3JK0
kOTHcsMdb+rM9gaDYFL5f62sjdJr8ALugY5KHp3CMpIuBqSEi+gI0fv5Ip3HxbXY
hKHLOlRPuIY7oFD3Vi11kD/AfCMfL7MCD1oy7+4zx1FF8GARawnoRQ7Dhkgi9dQe
KbR361tX3XBKncGscf/uTcu83nZn1kGrQ91EraXho1P8Acj+pSX2GbpGHlNPjH7W
MupS8KX9dk0Jb37wL4F0PYO6dVvxRicPOLHCTp4R9YSVembTbmjoMRKa12foJEr/
dl4HwxbDpEXXa/n05ojyLC1zB/aia7i8KWT47qo0f5Z/vItG9XIDhH3O/C3p8PUE
j6SRqGwQmOazW6BDP9keCKkT0t4FXx5IbAB5Nz0F0qnrXlezgw1EbvR/0iXN2U7H
uw9z8ubd+gdGfIFqo8l3EfsSDQuYUZUfk51S850FK7rQEKU7QokTmOLM71VeZF0+
aKioQaLXTKW1lHOFO8/5pvGI+BDd+4immIJ5yFzQHumvvlNxdOHMgYp8PYII2rzH
lxtFDjml+ENnsQ+gGvlTg1/GRS8mBF1u9slekw+RpxwKJUHGdrlsiyyY8Lfei37i
jgvKKZaz/bNPXz871d9HdOHeErUBgSFFeVYn4yFH+ku/FIxX+9KD82Ur0j9T1mEV
3+i4S+5ujx/gbi6xWRtUTodZb3z/PI7KnMRnAiP9f/z8wprZEMi1FBUOxrNMebWu
2oIgsWrPC21X6bhjEAfkUIaIt/6JX+gGH+CKgk++hJcFyogcbLlsdBtcZ5eXvpTs
QoMUWu3JDS6HEtvwbxLMwLNOeSR0DPY4rXSwfUUKFJ/2fFsu7hUEwCyViOCaeUrX
0RiNrdetrPgVtUeXuFickVq3g21YyP76NToBvoktt8MI+VmyQMJQM4Fh957j5K0G
VjxO5mMVe1nW2WipSYJL2YDB6j3q8LTbUwnfEsBgkkJwYF6ZZcODXZNSxDbmUAmy
ACjNX+DsA4Wn001txVbZ/g5gTZGRJ6USHloAjvqSPvnAdCclQ9vmOV1m53atPKjk
LwI/rRt+pgqDnktUk8D7sjxsXH/OAQp1ZalhvmbeEOzqt81/hJJ2YshIGNQH3asy
4x6OQCIDD3bv6vEQYAY+8Ntyp9J6qOBSG7qoksJbLKzEtTH3IcZGyYWOgFio9ciW
GcNtFnxYkYjRF5OBCj7UIEbXOv2/OZfwLFTO+rLqQ2f9BkGk3PzA2fktSXRu1EJU
Yi+XDl63yCeYqIdEzX/eaIh1F6BOoYB5JyrjuJNaRRkOkY/Kl0kndnlMa/OjkAZN
1Ly3MfPB0bSuL7vGuwvoJPYbu+eWCP4nhxWRO0a6Rb0IsEm0sMli9aS9+EguaSK9
FNFHsTSDt2P504rrwI6ysGwbR9Wdib4IpXYankvZGNTMg3HdDtHIBgsyIEQ06HjJ
K1adRQe0JmUfqZJ0K1S0kuBVNgVB/n8Q+TycihdcdAnvjG/Ealmg/kd+iqyTmAK8
xYdR0dN/oZjhF1F49PxR8RuidcGzNi9u6PDtnh/XMXM+oooNbapDCXzIq4FUYRzh
Bbc5ZEaahdXFI3Jq2GMfwIhQM630I7fBUo0VwSSdV7u84D1iYUGVt6exDWQq1lfr
pXcGq/ymjlRffwLMn1EILTzl9hv23kSPd9kQLG8If+B1Pczjwbh4ljHbNqr9gx/h
PXHyCBEg/8nD4vHDOAtQWN6xaXgAK9I+cNxvgLGzpfueioKw4uo8bqJ7D4KYfb0e
lSXlA0ihu3l6f1lWBwiPSyEZrB4upNNGZvH2Goravc5CPKtBBm3Cic7gIu5knkJH
aClMv9haXQX6nxWy5RBqG1rzL+XW0ggUObPDomjff6KoelEmLtc//scS2DbCqoX3
YeoaBontITz8qB4MvOKTrOBxLGIhCJY6Hl1aD/Q4Dkb++ddWsXuAncMWd8ergdeo
vfwAUv+dYegPM/EXX6Ud9pblNJ4amWt6A9eT4BjJdn0q/k+OLd2GTirozIArG5fJ
JUFVJshBLubVda7wOZm6k3cJhcYSygrrQQIW+ps6RlbzSk2oa1ebiipbRzQB9wuu
EOXvdUK2bx/zVLeYruV8SAzxAJF3Jg+JNlize7Fl4QqKb6m4Tyd+vnYIG1ynLXhl
I3WtVC6Pv9fFNQYqv/GZvb4xO4r2SypLAePj7G79eXYkGzQSjdUWsdWmoGGglAGb
jf4Vz+98POoSl8/PlflcJOXvyB4jgTUM2XysTqnw/gYxClOnwze0kRbEoDcbERCP
XrndZZSMF0zv4+thTR1uZnFCYVFccgDFbTmAXgUGz7wEV/pKIxnaU6X9fY02sDjz
l7r5nkZle2JUgiys8aB+iaX7+NszwxMk8rnDkMJccQTPT4T/q905XOIEh1oebIUQ
Vn3j2MI3hrIfbTtHWquzWW8Nw8Uvxchj/Ka6JAyBjfGTbNUjZvVSW7rRmIsjrdOX
FoEMRv0Rj0ZEJsDyxeFU1+x6EJ4YTcHeJg6l+miV5M/JVs2T8GZSaS4zHrhd2Ugw
DHpraDd6XUQG/Ub9x/QCXErmR6jP97bR0make472HFwnIvlNayQjnzESB9jb+K6j
KdEp+/r331OA94bqXIF3/wRBcPAPV3qBCI2ZLvzKXs4jNuFzLODWTD99/MWC8HbW
pXjx2RLHrvWeX6/HwrPmJnnhyaG510ZOdK1J4aan4FEz6xVT2ul+uEIT9Q/vfD+m
v7Zqr9q6d7Nytp769ce+hz/y9mZNh4mNlMfH9/AxjtL38zoHmqCw4PAWmXCGnzKU
vviNzG/86xaz3B8v5oita32nPzoGrFGTXEeOov9zYhy+7XQ/XNrGotMs+bBuB9mL
ye4Qkjdqsz1KxiCLoiEm4bJFlACpx7hV4SvwPcpnso7hIEmoJK+sR7FXp95rhWE1
zInW4ai4rUP/PJamVe3o1m+UubJzC3pNQM8qOLEBLLoRIbC1k8clXGIgir/Fc/MH
uk1q46VjTLZvWdbsZT8eIpRsfYLlnZH2NjisVTjTFCLuER0II+gDx92y2+GiujC6
7WkbLlcJJT/8YKAQ34e421pi5SUgDExR4A8LDc2XKQYNxrLf17tpaf96A7vpMIph
nmn1RMjz0yTB7irh6aNAfBp4RzkzSvJLyrHNaFdW4ff88LeadDR8HYMztoIXkgs/
eCDMu90TnqF76J2Ak/rdTbzvsZuxbaNXxMK5aJgaeu8Y9+SOe4Rm23BW1C8AYlEu
JbmL5vwMfFSzJ/wk+36R8GLAneDsPp5s/cnVlJ2c/FhaXoQPa/aVTwt2MbPwdzUN
SQ6qkpiArRqwxDR3nf3sakYcv1TxnVHSGadQVpI3BBj5owj59zbLgggfaacJ7SmB
PY6NS7IQ9VHJxAuqQoZrmhbu7yfscNYLOum6T1OQBSry0oWzxlW62j6SU4NjnSYD
9ORbwmBwKSQkY0X4U9cscbjDh6Y06rnzLQpw0GOsU7Yz1h3HLLNmKe3gYLq9QFsj
rcVUn4/O+Kf80fMy9qZUirAXKZSj6vhGohD2K2OarOl8GuupaHhDpTO6R7AFcZM/
DahbQbJf6O3JrmedOX2YCKbNOskgavmMcS4s2427QdLdvQ0PBx2OqPpA5qNjIq24
Z/+7wIzmTYbbnBvjJzOzS9wLlGzJ0RjaPNEQNfxdFyZt/+FAz9Pq+0qFf9z4gJIp
Y7PLoWvmc83qtuUkOs/37YsrS6SGxb8KZORDAVH6EA8URD8YKPUBTbD20k+/NcT3
aPXsL+tsGnvef5yVGbYG8HVWjMvQHZIkbw2KijgLwuT3tgVf+B0DnCvOfUA2CPdp
YkTKhNSMsYTMU/TDMCVYrP1iCa3ZRL3DYGHB/dwr9LyklgyBrWszLqUhGmVspuPx
Lg2DeVXUi2zVRob8OX6vOCsy2lFRRFlUYK95heF+A+ENoRl4wH4ULfym3i9GV9s7
+OedfiPYRMrpuB6pUsIZsDR9xYBmR2SXZR7St23z5X3ud7We5t+tMms1QKXbOUBG
RQtTgOnVb1gr3rmWbG5WC4UuchCLhy2dpyOhOI4Jzudfc41XdhhEA2JtwQ6cmr1s
9wbid35hkDGMTkAMW8UUvJgwYg7/Z8g2Nf0kk220fWYjhLy0UYKah+HcPSKP6mXd
4kW1menebsI9TnCkiZOKUry4EYtZ4JK3wY00fokMJpXWGHM++Gdn+B7LxESVh25x
SNiURASSLD/o6aFwBT2myRHxRC9N27tDLABcajJj3Zw5/GiUlJ8PY1QbE35xZipp
tza/WG2U1YdAaE7nzJ5dT5Gk13Cxkz7R5fArpGqoySUmJ3Wj3aLVu4nND9s/OrnY
gW6E8xQDKSMjQQikFo/WAjSaAoQvZkniYvp/zzU+EEz46e8ZuCWh4N4lVFI9C1ni
yD6x8UU15A6rz5mTLdmIAo8TKqf9HL1LUiNmhEzaJcPZGP6bjdvZeA8yjlUB5UOO
boTugf4XO5Ir1J/VbEImvo3khZ01i9+zjP9h1ioZCnIDPBeXb97IWrg5Iglla2oc
qwxEct28ut51lHEb9oaA54oYZ1MNXPDS/maGUP2kCrbLolzjSR4HTg76TslMr5Ot
kj2U32vLBGlmhVhl2vvWnxbI8IlN7q/zM4Yia0LOIHXhhdBJMN8QYRIi9R/IVRD7
DGXoTp/2TxAYZTykOCOip+viL4Or97Cser3kuyoIDHciDJ399/4fV+0IJdzahkpc
r1TtaldYj4U0UHFSX7ubydZwcR26nQnyM40nf+yn/nOedoy1r+hdcUK5Y51bchz3
GEaWuQjL1dyXxNsZHNCwELzMmc8QC+nEVmyjfHY99yA0yJ61hl1bObGZgoigL6TZ
f9upL1gsZ9mTtGmZstSiFk/p13xpB/pWfEWBO35b3K/c7p3iRH7QmNehcCAQDjz0
neeDVObK9lYmedZmRMY+KlrvfBSeHcKUEEKOI9X1iEznb65XdScsACclvhOgLPah
IQE3ILS5lBxdgLW3LWAmvh3SZX4Rj/wU07Bo2KpOj/OGehVuuBVBcKkBCk39fYhd
luCyXZh94NYECYuG74NaCLrXOk12F/ipxX/dHroUESZ3dYhhO9D0VrJROkYiGRBz
MuE0jlFdHqgG0MgJItzESDUJexV09LXqT2TU1W2Mb3SI0qzNs/2jesv46zN1u+Dk
ML17Eabuvmbim/JE+RISyWiuORha/TsD3c+aeQ9OQVyyW1xnU6Fxbr3PJWNBxTEa
MJWcRCzcKmKTYDSDPB6ZWoOt+cK9k0UY6DD4AqcfE7tWejJGizhlOctC/FyPjma4
l0EHRyuaLNU12yEEGGgqkjkR+jOsDVrNJ3F6L6aX2AhghrB4hWD+cKj1qT9L8Nnx
83lu1hmwFUtYXR/DkE+hxdWZZD97virx2kLcQRIDU24xhraGOFze86TlpQ5jhVAK
rAk6EydaGU6HNmsmzPiQsuOAmQaioc7aEi4W1f3xEj0Q8dZz5YsAtGBj4Ou9EzXm
M6N87Z9A4po95iO/s/1RhLLxY7kZxkeOtkgJ+t50bdqLoBNSNVsCaCFFSIYQFl6+
5g2EBVrnwTxFOKku3KvQeFH1QyHiauzJ/JdVrv+LLk9pcgvulgZSCbODAqLmR+gT
OVsMQc2Paq8BWsUpXnPS6R84SE2I3NTyHSnQ8fI5hBHqfOC806zi4SX/LftKvgjH
vr3oFhOXawoP8hg4AINU1XvKSynC3j8T+8mDVeWwWX/IgjihJWy8qLfbZ6+dwp8u
of9eBWP7wVDRZKHrarQcB8p1vsnLDNOmfCamCk3Ylf4bH9OuIt894xnBNgTPMtOY
IPIK52uox5kyydqKekz6pFblkmjdnliJoN/mZhls5yvEGWuBMwh/BII7B+qtXrUj
yC7pvW6zunTKhmCciAm4zbCqPQNqkPu99ceOHqozvyPe4SSwR3cg0LZrlgI6gn9Z
Z58roPfv2+ESu3HmJg/ehZ8J+nCEG+iMoZc/8LV2Z4BLtr8z8iTJEbHQ6QvZG61T
oemCxMzcupujNv8AyYvW3xiQ1QaQRNVMpSz+VBWCdVl4sNJ3jyabLHa8A8XCKRZJ
cWk1A3ESNxbj1tAnm978+JrnCetOXvgPzeDNZ7uQxgbSo5Gh/RXVOd0hV5ivXURA
lim5q/isCY+5j1ediqm5fSF6XmuFto4m2hGvgpYz8WOOi/C/anQXR4btm79L86r6
kpweeDg8xb6fBHY3w3kWwurF6C1/xoHeahIfvg3+8KA3vuIJuChZLEJfZGE5uRRC
iCVz/2b3Dvtp+jYZ34KFiwF/u6rG//Z2wWkqdBopo3tw4n9RMcth8C7rQXuYSQWQ
QrAfVBWVQQNBfzJrA+yok6m67GAoSaRnGqWdTWf6sB3dUlre8xAGnjBRHYhDSWE6
EYShrz7eyeT444kjxeKxysPOLH4SvcFWXOr/uPXp2njb9Ay35pCHIhlvK+9FWobH
j+LEIozG13Zn5Ksn4wytDoLC/XrUmU21Tqg12MOZwmIKP2lkvHVsrJ2eTRNzUOaj
gDxhVxhfYP0PV/QGr6QJz+l73y+ta3d8d9233iCm5G+L4vsXjdfVBpqqPhGBXuyz
6V8VG6/Bhchz+3xPzMWUuWteIm+JB/DCEjmekF2J9KLdDcuPd806DTd458OL7Zrl
rRQmG6aafAJG83ppe7LzYHxBegADNQDcwihfFPNZ0u1QDE9GNGClJO0s6aq+AAMZ
KmCwKH8hRW2868vU913yVhcjZ0llUF+wnFmYcjmDCrlhsPQ7Ne4F8tdPAnC3JtEt
+WAC6mw22RN18tNFtlnCQNjMwQpN7NmRuSw1D02cuOfL+vk5f2aHfI+Vqv5AW+e/
LGoDd5yu/rLDBZNjY2tXyFte61rBj0eztkxFkzyul8kQ9IMRFy+sohMfVyrI0Tam
I4gES/VmFBZIaROsjjwi9vppUrM5Uin15ecSjI5gj8Zjm9RlD7M2et0343NwHhoz
btufAE7Phsfx/A5gucfTMLZ844SYpGJj0v6drJk67m3lE+hvjI3enjnOPnMjp6IR
NA/sJHZ+HNR3qQaGTWJrqeQ47MExyE+Tbl7KXOovCxE3tsOYds5LszmhBTuBs7Vm
7YrrfrKSJqkR+o8B+FvCJ2jvJY7unWAz8xi/2Ci7ap5jF9koVC7odDt7AB4jLPex
VLJnlZSh332XAjNKlbe8GooMQGEngFNu421doHCI/AcX6gfIzl8V/Y3CMVdJqGEJ
7hMQ1Z1/vCM4QUptBbMhFB88KN0GrEYFYNkVHokWwvjYrALj8OKdgQJIA1xApHdk
DeJ0MFkB0Vfs4cii82+f7hJY+xPtCCWtSm3u8593vvA6lpDYcXm0OPbLwIPLXEQ3
xaC2uOx1+L32AJ1k8qI6RBMKb/9Dw/DvO/XKYkmDGnvZ6cCZOVt8hWxqIpRZ4vff
bIdkcy/8AUZ3Kwj2eaOdcLgLrwB8M0TM/nRLPjDtZF1SFPUNf+FqFF0OzjQmeTNc
FnIy1i2esrdwNDhoIXOfWofFJclJ+SVV0AWTvHG76wGnXcxduwmHzJSf3whW1Uog
WhHR/PQbrqgp6NX44mrWXXUBW5b77A3qpu5t8G9yjDInVWuTMgagQ6jsxLJ8ryfP
4fhWN44QJ4eVPNRTxUiG7rkvmxfoSh99akbHGDSk1zAbk5rvowPY7Kv+jJfuJzOO
GosHdSfepU90aqj+6aqqOWQAC4yIhlF/mq9sMs/NKyEEy0rEVk4gy9dQ+amlTS6M
h3fVNAzPuDRssFSJy2ieRBYjup4cyo0CH94AA8CwNhxSwtQAVU7HPW3N6IXEfE6E
uVf4v40YlHML9w2PLJ7Wq6NlofO9VYG4ufnpOwYBcudon3o0I6XAZSjlN6wsrYcR
p+FEXVMLGRkdGLSzv95f5R6koSazaoYwXE+R5kZqmlz7cYe/08j+30rR5v11W2JY
aMZHv8FS/T9r53F+zs2vGstZSu7LWmaAYE0MiXnbdBpZC5AoCQ5udYOYXdALOqF0
ODqGFRGozBOqEtAeEu8WGTV2wnkKm+tEMWkcCg+2DY/tp8El0whonrQGwIjQYtnT
jgPQ/6EBvaYFhmpKIu6YbyDL9BRt5qbOmFJFOtQDAiR90FYwh6BAxtS5v2+KU9iw
GRjemcT+3mIxKuC0u0360S3buwT3Xlylm/c6za1bS2T6dzoZvKObB/CWL4O7P2fi
nMh06wgAt+DuuGK7eocQAjqgQ4b/AMjrrqlSSENP/+V3IqzprX+LVtWOsR1ZUCii
3bMtlzEW/E/f44ZSjsLJaV9dGUxFa8SNHGW2MLX5ARYSA3q31mD4DjGr7OrJW9tJ
Tu4d0MGJhVDmL+WBWHJ91ZwBQQwq+BicbvVp8E+fx1/EU1sCUBkorlOVR6lIF8O2
rOZC0cYtPA1joI4Ivx7GuAnnVDHcr9r2zL99wfgL7Krwf/RPqA4mHByRnmXam4Xw
gpmkz5eXPc1eMg7+Gcn9phUS45fe4Mh469arTdvVUHTvf6/AMxQPnyd3mrEjhNs5
GAzlf+Ah4nWcThIxLfzJ7/MJyMy024ZZ0/KaxgdeaTBo68gsRYfm3l4EkXszXbpg
s+R9dybJiGurOV3J3GyOriYt8FJ9/nt9k+ShaZ2Cbfz4XLLTT06xI6eqjdDIpOO0
hOMS4CzW6bEIIrJOwOYhDutrzqWZSzKie8X6X/V61277My11Fqq40iZT+6ZP7OUD
+Fi/DpDSFRSYBOxICxhm7ZwH3DHmH8jbMNtUzpZM8htF6CHkjlpUaLxbGrCcbMST
e4X9W+MnNAVcVmhhdIwS8vylIrAig2/iSm5dORrITwX2C4PK5bQhdENzqxuQwGrQ
XGGGoKG1gR2UrIbnUjtRRByVJ2Lkvj1drIIBRb6NrkULLNlEmVh8p65L01yvt94d
wmsVbALjIWGIz8R3pSikRc89EFeRK5hOYDqk+LZSUMTnsch0CmgGcT4IA2d2E19a
PWsRrMLT5WdIq2+fl3TBR6Zz2IFYYzPACwtXVdcZ/ozqJWbAhT56HLVTobdjhXYU
PwaJKkuvQvxfHjABbFsOIlCLKWkKsCxnaQlki4RMknHiiOpLYX/tWBwT4PUY1pgo
WdqH6/WEI9xlwWaTi4KZSRzILQBSpgNcmBPIztPHr2PGpUJ0KhNTZFNZR6tnohcc
Pz5KQFJz5xBidy42xtNZb6o6py7qG5NsxcXqG6iiEWHCWUPzEFb61KRC4R6Uok3Z
4VP79ZqgRMX6l8Ytc+n9J2Pm/JIAlBOm/oHuPremDseR1XN2Wk7h4TFZUyPV55hk
XkHX+VqRP37xPEUDBa7q39WkdA0tRdQxCurDg1Vu9jwC+0zVvMjnVAz0KdlgCORC
h1dJYGR+ueFfJWA1gKTNOqdKSQ43NjyNzbvKw3dqaCvAgUqp+rfMA2V/Xlb/5suc
BNKF6UB6Unag8RhpxsmaIcHh4NfVtZ+0IKS9Xblnzo+/DPU9RKnkoJ+Y1x0wJ+2R
dZqiooq5E+Z4cOIe0ScXCL8uIrV7fr1fWl4GF96F0zn2wL091mkzViD/So3wN9pu
zOYJtDg+eunwwaK1AKyonGSdzdEaz4IvPWmvFdV7E1bvIwpabuhwOcctpUCN15TV
YShNx7P0szUR7YAY85wpL6Nr9hKBNg1A3X30LNcu/wQVToWgAZxheQFJH6+HL+8s
vszwa7w9acJ4EQMhrS4XauVzu0a1/hXQClkYo4QYHcshueOM8IIh+43sEuHbn2IA
X1zb7aeFs1VpfsFKh1isw6xP4YRi+i15fFHfX17sIq+JqyBEWas28u5INFCfaF46
cL70CrZq9Lj+27x+1rld5Cw0TYkxIkVuABKrVrPIhT6ZHTTnzIZYu2j1B0l0pOhP
gS6TTM88mmVDCpzhsuKTie/L1b7Xf410rObE/JQxMI1KwMIzWsVYJ5Dxtoilgi8C
pAm6W8IB2WZLb9WA96l/GKXlMRx6KLXWqJ0FluIHmbyR4KmQpf+/gAgRaxUhde0K
o3BM+QMP56FKtnUYWryqF9UE37aGL+hIUPqhD7+qHNHbjshd9x7NNzt3SeS0O3rS
YpZUy8vygNWgfudokxB5MnDzxl/N6ATUhPWTRxwiq+x6ZCJF3uulwEEfe5ifL42H
lXpQyyy0rhmVgoE97WL9xGQIKiteSBogoNdZjmpfXcei1levm9BHseBXw6C4maLh
l2RrMaXMrnQvrTptiCoTeSyspHruZBynb2lyoHU8JatsLFWQIs2XhM8CWq/qV5K1
i9wrz9lEO6rkrhohY6PJFo1igwime4LESbNgCqO6f3ABN7xUnpPCr9P7jZPEDXY5
pRcodIwP9T7EyAJsXnCFmQuigiUohq25rS7i8Fp1YzDZpspG270Nhfu5uUrKAgrH
oTwpPXWvEsQQIawgE9oARKBG8aBpGbzHO38W5TwhmmZdgqeXDFA5mx3CebkwKng8
Fsb/fpvTrX3Bi6Avt//4Ov6+vKpSM0kd0PmVEXmeu53bj0IwKKuXjwxgclViJret
BtRy/N2/wMgupPMcdbioCA7fOyTnFSSVhWVpJCaF4R0VNANY8ku6dNXay/WDah7Z
BRh5PbEB6m2QTy8xOtxGztit4bI9p9xpM4vrfPk/0OWJVkbNHnlOlMWB5Qup56Ku
lJBqhAT+M7Mfj9eRvoN7LYR/p0M5yiUPOcqVvFFVOmGYAqcpIkF45ihbUf7loh9+
I9cobOWAMZoY0Ufy1Q87fC0WFCS/O6SxFKI23RCfLIEhNHAZP/3ZpQV/KHhblrVe
O9CyRMjY6ALFfdJDuJO2X3BiVzm9co0DxQcAUYo5jCejYY/7lwEscUfGqdiOoNzN
R07YDaptpyN9zIwlyZZRPHcxb2adPryuII3XjITGGUQ0mSZlVCdm/5H9ypkKdLOV
Va3a0KQlYUZwEHz9CNJeLsx5z8Ue1hEHHbGakjuxacpKiWTYcrxyg/EUwzUqw0X7
fPUXfq2rYChfndckSAHg7VJhB7JNwIuSMM4dk+1F2fYznycGtt8pWrfTh6TTX0C5
mICs7xI3Xh+QEgCg0nReYt3xOEHg760kVQ7dVphuxYVHvXwzfJCay4xtoiETNAst
ecneEd3Bffl/ww7KA9Nt648DspktApxwiPYjKNRTzyoX4U+MO2wxzy8wdE+V7P/W
Xt3kPs4R/cDEDnlkqAh05XFjoVCtdzYbD5n9jCHy1JKdJ+97EalxCMQtYbOZ4Ad+
pL/r1D+IZiRdAYTIL/c+D7LwT2x1PIltwL7NS9pOGv4AIf8hQ6Sn9Bl+ydH/GtZd
XCo+w8PzCBs3Dh5FYIwD1wbaLUCyCL2xZR05sZaREGcpZIMcyFkrcsNh8q0srFrZ
cfKDDZ7W75rIXpeq/EWcPRriCrFe1VYIG8dqgj4mWzp2IXcA5pLumaWHP1pj+br1
YJa4UKP7rjBtVj0QBGU5ZB8elPOyASJzjdp208NOJEVAlSlRwKwI9Fd9P8jtsVt5
nccfWY9uxqSjekzY2jEYGm/JNhTp+NPCa4BUATz99RMWPlWsxVFXXKBS1/xR4sQ7
B+OJSHN6CHt9KHQvF6txd1W9WwouxcZPwsPYmizP0gmOgIOhITo+1349AlHfDjz9
v13sYV4rHRlXNSY0g/WR334nZqgVNlEMV13hkvHn1ja1/oc45k6XCqkLVeZMmRI5
0DhF4M8WnVEtxVGfJxQ0ftzfC/tZw9caOSmKDo9yQ/Zcw3n3wcvknpDBFJ62SAAq
ZS9k2U/VMxtLX2Jv+U0/M3iZXpexNxZFXEpuMhsjxkmggzXrdy/GWcQNvPFXV7Xa
ojCFzFbCLkPuFovpmpz3Rr1XKbmd0Yd6Hqjy5fSDq2PIzwsWSY/uu/OxWjLmuMOn
dHm6t0pwbc4iw8jnMTMuaw5JeXVC4RiSu5Ra1Q9d7BzPgWAimmuYxhzRWcsLVB0q
N+BymfcfKOocX/AlyDXj2+oiMH0R/VE3/6h/50SB5e07svsGpmiepwFxNbrro/ek
pEebnabC2MHf38MwwdQrLSFqTw25QckiYGbqr7ZAiSLcwMCW9qsDhx2lhfT5InI2
Rkwf0UQyq4e/HYZBYY08pwverYzMHgT+JCrmP7CC+10Jg6SGvXR9rVo6Wq1qAUmu
igf2P1mZNI+WjfH8eb+P5C2Fh98UycLDWL6Ah5RbaZyveQ7PRz5tsUZNo4GoCsBa
XjDPAcq8D75ak+0EoET5t4WFOkZGjJjGXewgZnqOBMdFaU19asmtDF+BAGtUpy6Z
o0vyofQbSDc4oKe+v1gJLaV3EoeS8Q7eCcA87KKdvAR2RNS5Z3p6AT2ZPYMyXQeU
An2e3q99Bmwi8ALqf1Q9hnQLvMb+EqeCP8S26jjEfrXvGTD5HUoNVEe5lP9DElH/
/0ZosiSY2X5tvHLUL7q/ryJfox8GBOYe/Qdzu6VYWSN+QgKYBw+RICOW1oQ6c32o
Z9E1EVpsvrzN0d5kcS8qZu+5GviE1OH5rm+rkJQ0NGavw/hqHsy47s9CQYjiRRrr
R6PvHQ+nY3i6vqpOWr7sd/hEFyOSTq3+fSrYCFe/7Bwcl94bIBsFm3I1Skes9mwW
3AMRKKI4s//0+hrT1mGUTaMBW76Sr0X6zAmdiFcuC++pXEdxoav+MhBzM0rO+nHD
stgcH/GQj1IZTsIVXrQSXZdJU5rozOFSlRhEN0Q62SCvXk/DPwX+AhM5SJUL8NJv
m60lQFWouL+Myv8JuFSScxr9SDtrnCi832L8JI1Lorkwcgskdc0b9dARoCCYOMd7
6VGv6cW1CcM7ifuSWf2lpNwjKplmcy41ax9pr5Am65L63Mcn2UQQOgbG6a4+3D4t
+bmPNb/ASizbnhWCOwTkK6d7Ixhs1C8l0nk/e56urVX3dMsMh+bhg/gbE+BaZN/6
NMGfl2OlhzpybvviW/pWjNRsIT6cPurQmBHDzeBPfJ3l737Dnw90LWzhSxuf8pgB
+8f4vh5mQYtbNXuVxmPCDBACHKp5AVN4DqUYjIG7rQoZxSJtml+EmWQpRsJcW2n8
vIsQHqvwudsbBX6HFxLHX18saSmIgUEsVKq2/jYReOkibliA3u/GQFN26wKFmcoX
S8PjK6ihckaURCx0hviILvHPoF0KugYm1WwXWN7NYWkguq8TM+ZSXKyCTn0SFbsP
f+gzqJT9DfR8XQDRVWpl2q53PQMWhG9dD4neX8l3uNRaG2bxHfHIqVxBiwrZWLzW
Y57BIun3c+nxzrz3ryytplNCSoEtHXX8+k2ryROcZe9PtiAZEjHUi/wlj5ObGoPy
1P0+2fXyjsYl0ns6Vnez5A89XfGO6x4eoO8jP84VRlE7WZxutixJ7N1wU94uSS+Y
v4bf+37CtbESymS+Ey/g0Muj+WRZ5DIZeUBbtulifCAfhORJEpr1XAQ838BiUWoT
kmblH+envTb2hd+LulWaRtSiGuzX6nfpnmW3nBDRRizsenmAidpwitXlWnX3yqva
u7AXULLv9Wjzpauau8XutDVv4ZNEIx2TRK/Vyu68vS9RpmtfltOri2oYVDEhM9qK
kOz48EySLNwrUcCMybNIDp9rAIJZGoac2mN4Poy/ux6T08nv3iG1LMhLpMzRhR9/
pSGa24BxcwneRqsigfKGaW5R38qxjJo1FCoy03ucYP1y2RcZ3uA04CVE0nJcA4ay
MYG/uI6z9t/N6qy7kpGGwEygK9v5mWKVgLVVu4dkfn5SxJwgCk18FNGJ8pVmM3FN
UqBJHpKH6jM5SWi2KeZUpcstUEDD+OfmRFFuy8lskjSUT3khmU9o4HAcd/k/yU9k
njpECWNX/hZOPZCb6XQ9b9fajfjD3Fjwyfn4qxpGwvak/WMxvTzhgdtRst+vjfJx
boUXf1wX3fpFV+KadxmERh7VwGRz9kIM493whb5lyr9oai4T9wL/Yq7l41RUiCf8
RAuXU5/ayJAV3ZlDDF90tKJ3Q9E4f8LH8XC9qs09O1MN6WGTXbnah3yItWFCN09n
Xw8gGWqZHlGr39L7Y7N1ZUn3wCoqvrMkT23SOJaAU13vrEZP7sEvurxDJAl02pxk
S06NQ/RgPkTXMLc0IIIQoTcUUHrOGiEOEr2X0O7rIqrsBJVqGKJBdz7qjIEf08fI
B6zDulBborGSuU9FuSeQ3SK0268Ho+v3zF63/izwopuOnGXsqPxnWr+eP7arG459
IrsyEUPyNjpd1t9VYarfpAGORNgARwt0nTpBooQaDMtsZTcV3zWYoIBpI7lxiIHg
AC8ZyZk3YJ79WzAbnnBdWevCAem6TlE7fpqUza91wjFO1gYCPbtcrAEzN+4Ni0gy
c2cPqqBKLdcCVvxY6rxZMC67CiC33qheUOvZXfITI65rEMR+VwbO0mRixFihOSIb
8ImyGoiN0/RDvErPHoVAMqRL1Mr+l2HOXaZd617u26FRPIvkYoguI7UV15clDjos
0am/R9AmiQxsK0YXne6bEwzdcGXpE4t/M3zvtgUcQPqSC1iaBa4Yiqdv7gr7aRdT
e/pRznvANe/6oTGPRPSUG88ra81PlCWlv42LOrcSo8I1D/7QdXBzCGm7PReu7ozJ
cdodrgsiebSsZi4+Ancjew5lftQ+xr/HRaAIEQKePDADZpdx4Z6cv9Z5g3S9MHU6
1R/9nIeSbqAJBiVyM7W6PsQE3tFIem/J/qbfDRe6LFbSiopdM9mMIilV+R5iUkBJ
W9TTxFi0qejdaOGn4XzSevoqDtFBJkJcwi173UGeZwYjWxb8oF5e+gxHA19oGpXx
t49HgPI/SBgAH7+DgfVzT5kJItbKOUzM2z0Igl/0xIlZuSlikfs/z8q2yWYHs6Fo
q56Rfi6mZQzGZ4/jmVFprAHCsoYB3Xq9VApZrRm43QRzTqllr8sFYM1Uu6HOa3EJ
YP0LmhiXuMfw+7sFjXfF6ZjfWNojfLFrXmyNy9+/bd1sbRGp3I2k3lPQbugbuDHW
HMqRut1upF3nav+LajlAlteZqsuHDWc0Cx+Xyd5ngnmnJgqy8F6iLsm0bRf+wLCo
cFxhMhR86qFfQA/b0WkZXopPmiRyzF65p7jb4wEg3z0zMxdTlzTUqIYxHlIMz9vf
SVYiDt+MA/W/h4cV0MPxnLap//3zIDPvLx+/by+O5c9xaOqyRxbIhde3SXLw5j5u
Nxv0ku/6iAM2BgpdfXCv6mftp0slq44WM2bHmNrnjYNmeZMZexPDBAMpJ5rB5X30
gXrdFrp6uhEal2/jmnQnWYog3snMAGQStY7hchz4XQxS5ymsbn3AkjF0lXEOD5jw
VFTl8YrI4L1udKgVLj1tjUhU3KJTe7uZBh+RQHTbCvEAw4iTRekVKJxwL2QJwnSP
FWv/M3NCMTxw2JY+3w3xcYC5u8CAKDiEz+R99q30mRnCXZQhxf9GGuy2QxAsv431
uWXVGthVpmkW5LyX2IMWN/5qLYDl8xZSIY2/kigqKT0V7jgaAdHHEhswtkT9kk8R
ToG2+IQP9aAyU0HlPPJilazdW84mzB4IZaoy9HXo8pMP9cn7BDizfwBmuT8WvMd7
iDh22x0pQarWF4DSLnv57gDcK62j/L2YGP2Zmn8UC/lWoo1rCa65re1Nfie+WH3/
2zmfPKRZaZRfhqAKcIf1wkKe8x603kaHz+gKagBKdqSeL0Qz+Ikq6nARmK6yg9TB
0BFO9E5cB3UbY5ooJBfA5YAGhl0SqYpmj7l/yeu+nvy0DgkkCQGjOspHOZ2kfWyY
D0qtIgJcRtYGDkzraTVLyZ+/nEhR8ETwZ3drhsPS9q4gzPOXCketpgPxgLXM+BvS
5CmfhPXCaBQgd3aRx1huRqDcVvvOqL+6Nqi6UIlDYnUsyo9ig9Fkfcd7djc5BbD+
LKVA7EJ0kQ7YYsksr4MXgwM7ogOXfthoULP2DRZjVf0SBQ9NJf2GICjOy5Pu+zky
hz7wFmP3Y4imqofTDN1XFSNGNMm0LAymroIUdopHNJzHvrfKu8jJVnZqS1mB5tSh
dKX/GTwZdWwMyZTwZ8AaJh0fOCHUrUr0L1gx1MmTpfm8yA3CMhjXZvLVp7fdJGWn
kR+ufp4qPgRHzteLw3LNGP7TqX0MLV4imnlmOSERc5BUHnob06d9O59+WKZA6ZGO
VgZvvfewZPSd/Xr04hDW4KDAX7S86fco2AHR79LChTD0m440YS3srC3QjL1zefpZ
33B31Zpxq3O9qvysKZH1wJZIOwbHvawbU8Wuuy8lQ/jMpOdheVX+NsobvMQWce/G
unq3Lo5EvLaABWzfIiFYgov33ItFBgfmyGKAG2DunwrIfcmrt0nFBTbJPBqOkxMQ
clrEqZvR5FQcddCImai9bz8uUYsWXlMsxL8F6tErUGWzVL56tJzL1g3jgBlsuTJI
bbm4WS61Bq8mSka/x3DDCSWWDcsmJ6mZRvPJxAV+0vYTDWr6UhNyulaC10Sh38DE
otk1q9NAp4H9rfNW6Gv94U0yvL4mkn2eGzoKEFDpevK9GuFtYEjijan/A0ueL30R
FkpZgiKtT2m2jxo0V6xc6BYIVifNsVD+Lw/FRG/Sz3Cs+O6Jpk8Cp5//suktN+Zz
WUZrGOniu8B6lwa3d5al9OglUbMTz4MQMOJdN/yr0ELJXhhWkRQoVWBspu9RHTAV
nQ7Uznx2FUTvkLB9yJ0OdGetNMaknM6f6bIQWJDTs2+RQzzrKjMgCjQ/L7d7H7zj
MAQNhFfHMmqbVj8WRZ9rwA7q2yLKCivvjY+GnVtIDCJejH5sMf+rgsv5n+PDpFW8
i4laSkpRza6OLTAwlRFj8koIsxrErr6s8DDrblvDOhrY7IfAnvAUTmdwWJwy2BY5
zDMtuOt1HxL8S79cvEbFVQx6VybH4BV+kQTp3IUL3Zr1ErIgFjVLNBrPk8bmum6d
cw8Ww6s3tT7ohpkSCN47oaKiKS/vBVNk8oW7+8LtHS42Vq0GYGbehs2IsbB4agN+
IzAvOjja1wvEEfup7TKIVKdEPmeDhib/7Wm49hjeoUNb8CBhRmLOaIglWbpB5R3A
wB+K8niB/hBDE2H4Q1V8TMAuKjRNybvIkkspCRb9AgRXaeO6TFwMkCNH23FoBHtw
j1N9da4GM2NGUZIJhrFFjD8/8EbQPy1cSzmzOyeyUMMG3pWispgshhADe+0JtNim
I0USiUUaCBwHEa5ARdj8c7MzZ4VBU7VfJLxE2JXH6tDRKPk97jBWPqohjMjXO0QR
ANegAS+ZOQuHyS7TlbZyDhq3UUQM8reUB6eKUUIcnmERZR7MmAPFkSRuPB597xBs
Wia2LgUqxNUo57x0sJOXsjfnvFkX7dgiSfaOqHYDmVLxpFWG7RfTL3e7FRUR+NP4
JgGkjxHiK47wzDrIXUjL8Pi2Wwz3TE/4JK8Ietgkn9KGMlF6ohLDzZzinnRmrNOw
OiEquQo5w8VnJM668v8zVgvC9NAeLNYpMV3QcVI+ayJkc3rMbtvOkL0cBiQcY1Pc
4QU6aAXh5cKooyM5ugmmfOlIsHPAeKmztMEMkFwQiXKEF6lR83xGuHe0k1GWRkcy
8RJjG81T6FmAdA9gr/3Lwdq1DcltHHIBHoK28B0LXRwnAlnxCaQr0AqAFNdp0xG7
051r/ZnQsguKkVmq0q6TWApYWpDukWJWmJCFoiZMW2tWmAeqFHJFJqjkPzsp7xJ1
sLZBWs8Hzh07mEQX3+g2hYb4RUUyvR6LyCp2kRrlB9mTFZJ4gwGGaeyiqKon8g/1
A4YStILtpCDpI2BOb/BTB7OL+gpQ+nia8jVLB5ZoyKzT0lx0aJ9wzNDYQ0eQPUFG
p2dC+PQIuX3njdJIWVykM+EO5w15NClstsKZd3nA7eafYCP9MGOFichEfVWA2YsV
g3P2u1iFCPLRvUSa4y4LlyevRq7jIGC18p3ZgLbiC2VUax3WEFrm10dl1pAxhFCV
jVu3KmSQXSMBuYyhVuKybHMdO2rN+LSM4NelzQdkomafC3KHcjZJLAD554KIo1fA
NwxfhwyNRtPPIUKdkCEOuA==
`protect END_PROTECTED
