`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Hk5/KZXnABi/slIb0Rw84bi1ZMojFgGHW5svYAKlpRZWdcGQcKGpcYXFNfc9Bneg
dDWUtE07M0TdKOzZJqY5/3uXUPKdghBSWFdfOh/3RycwO7L5X3IudYeo//kMsDKA
1Y+B22FM3ikAminjjz8yGNKZE0AlX6sJFim7gfcymXyGFD8ul0eeRWZXt8E+NswV
alIJRP26hbi0uF9t4KuzXQ9jbdZlKQLWBbf6y8p3KetPgFA+rQ34X6FnAj815IiI
`protect END_PROTECTED
