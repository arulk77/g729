`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHK+5n+kgTcZC4IEoOrK3QfmLyaxOwd0bvEK1mNIKcAw
iQFauwhZcJ1EEeXs7G62eG2t2e3hVqRuTSGgwKAi/goWi+ab0yTbv1oI8CoLbuA9
TgDQmSMutP5Al0f+5IJFQ3/kd2GEW14opOIvIWwIeDlePk4osLqOZ6n/wdF/hw07
/J04o+Ab1wJE6P5oI1d07jMLqottWCTYjFF9ljaLIqk9d7mXZufoUEsnLyBny8z2
ip4eYy17R2sPZ16t2uBek1oNIcuRhI0jKTS1qtVC2ePgHV2G3SpxprbVgWkau056
7gkvo/zQ8FEUhYcVS1XnOfTdKF6mt5eoyO80WYZ8wj11Miv53Ln84Ie7cYFynj/f
ijkP/ZjVhzbM4WU7rLWUqQ==
`protect END_PROTECTED
