`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C8yxELulwIiZGqXVChkN32dsZHq0zo3xgT/EJD6EfAQo
mtxIkahWaTW06khSifMqeLYRJ7J2+HQMWgdL8jKEZZorT35CgYvK72rLk/vFCy54
8dw1JSCYvolEPVqjEIn24sY2QbrFMmXQzPcrxzPP2CKIQNTBJLeLUcfWafQA/5pm
lDON3O8JF9vtvgSjKx3g/NDSP74nu/Y1QwiMH3FkRhnyMbUw8VV99ceTnSZb/zvD
5J/kF2nD0HUXc1oICqKz3wdvTHsWm9KcT9zv6qDgN0EsNaAmxIqsvCURqkZlK7A+
zKW5AglAAVDNQtnBbf7IgcxL773XcXwseHy3nBh+E/QByAIFk5W4KPzrjjbBoYgb
NO/FUhFJhjkmLVhHHHa1SmrTzpOOxqM/+gGfHHqrGsCKwiorQNjF+pU/EjQEpgHj
LSB5N30vJZyRhvpTFQvWhXIiML4YT5qavzsaDQvOBSqCrWmzibiiWgOHyXjq1Swb
Mm2a1O1ICJp/5pbGaG7AUdU/Q5Iolz9JNmLAhLLPwli0PAf9mEqxTGKeHseZW6vK
qZvJs8Xh/FPdnjuGBR1bezF8Op5HilSNLnrlqGE4hnz9ulFxxGi3Fiia/rVPnyQR
AMGgUjY9RsMiRttxeD8QVLqDPu3crERJIuFbGPPxQ9vpP6s4P6HwGNJh2FTQsppE
Vq9CDs8xZI1YmKsmkF1n+xT/MxA00IIa+E9EJVnEjnz2HUaSAYYBrd7+r1PBCWz1
A9HPCnwD1kipZbta3NMKREcnjggBMnH8nRPJfxybdjG7+JSm9DowcGCEPolDcHQ7
aFzmAjaY/ZrCGiGdw1c1ZsY/ydU6WibwwHtPNUMMFhPerral9Yjhk9LDGTzlxz72
zwg+ipqoVyx1sGiju39kV7WqnF9/KJaWpUvZGKyBuQVMNRkl1KPAKNTfyGI0Y5v2
ei+d5KqSc7T2q28SwIIE+EgOnG8u5ZRZS311h36H09hUPI2ZCt5R0cn9kUaeP9AI
Cp/HIi4wWWfv1WOyv8JV5INpgJwFOgB3biAU0b5kUmHqLX4qsVDJEbD2NFwKYBbn
iyc4tX1T2do3Wl+S7sgI0XJVCMNTcVfYUWJKuzE0Wr484Tpud4Lfnav1eswTkcaf
x5Hox9DXbpIVvbHKA3ML+VVAk42txH5/ck6ugRJ94aqeB2yQuYrbr4q7bgNrXY+1
oALEppy+sKM8FgNhgJvk4MKIdWVSBW+xRIJSJIf2wgYp+khE4O3+wE+OMK3tpbQo
vmYhNN0mGdGFTW6+ZsuC/ZLun4rgQMj/z+NYQBMqJtWQ+5MiJP1K1KWPF+fVMgF/
g+yFV2erI+mJhfw8kaJr8G7hSATQZ5mRwKvRG6rz0udrgZTfkNdTtBxoFEnVzzjE
m4t3psT1EeFG+qcZvYZblJPj9JN0LMI7ppQ4EReLNOTCwTl3I0LvShrVhMlLDNil
QZmGd06adDq7IhPpfYauoS0UMUARAqe8Y5za0lqNbB7fwk8tkW1kfx8pT7QO3u/b
pre4suNMlDmr6PpYydFgFaWCc2lcfTK23zGCa0g30vQTrZH4i+jaPA3gQFMyaSl8
L/0GM76u/hTZLgzN7BLHc3HVhnzAwHGp3Aig9ZLx9dw5T0YVEtVDTCjtKFVeE/U6
5QdFzkedNX+dYwoUjMZMOZ3acq8lboiIBNjfX7kJY2TfX+UpgWymmcQHySixF35Z
5QreQDInkdwSbmvGw2udMAlR1nwJ00SgmvBNtNgVpdgXvXz9f9rSsbIO1MdnTnGn
kOH6ftld5h2Y/fIdtXPMcCfrOgT53qvCSFMVRG6sntYmUuY2nJcQ79ewbv/aFaOj
0t/EZnB34giQ3B2sGLJUcDDa0P0OgeLU95XNKbLHfNL6SscWNfcExuC+Cub3VblK
mW+k6OLDH1z+WqKkhs+02cfm8E4tevt0PyKHfFNkAQSMSyH5o/CSwP5CqalaO+1H
07toXAo66Sc+dt7piq7LtKmNKZJwlwMGorFktDOKpmP5+nU0Yh/yuIRky7mvdxdP
z1riPl9qsqLe3e6jtMz8yfmVTMjdjaCydg1TiLr1vzJZ+ICsjCBtum+5gGPu54rr
qfpveg3sk+659new3j+/MVehoTE4Ta1e7l2GFW9n441jrKMdST1f2RvbdtjDHTa1
4gnv1mhcFTBUnn2ABLIeM+et86uwNrYs8J9BRjRnM2q3H4+5CACtVhnaDAOa5qeQ
/tIIuId2/HktBT2uC/PzrjmGkUZ5tv5aNUbYTb5CJ66X13aZmh7ScS1xSMMfpJ1u
7diYeKf8V58Dp1Zg6zDcWgZZFGnN75VHPV7kBdj7S+m/Ff/JIkyJHDfMJPuRnv9j
MtWjf9dtyrUa/P4Zw4Ho3zh7qFuEbgnIKqZifmDns1ozh1BSw2zb5mJCK+JM/LJU
I5eOKzN5iYgOi325/XUeOjeghbj23fjs12CX6IUF31mEXEZrZkvimS1f6G5XJt/V
DLvUGlQ56fHZBcgdJzf9ACXrTKnVNJA/4tuASVarXx9oVdj9JTVsmQRhNiULrddB
lxdwf5Tin7BJ7d2uut3InfKLSjtWH1eeZaWJDxmhMRvcCSrFRr3LcF0EusG+DHE5
s6e259dIk6FIa9hVZBKBmYcY7FqFWVsKqbSEM9qd5bAdFn/1Th9XUR7J0v4wi8x3
AVdJmuW+0xThfDjT13EmnLOtgXBcxYDAYBOxVFt4XORFMijUf6n3PrbGYLIELh8w
w6/4gR8kWMI9mJdhsSDw0Z4sux2qsabR+nBqBTCkbpc5rryQT6tq4p+cdNfZCBOu
GlspC2vtk9FGcfCSZHIXSpFSiOVTUd6vF3Ru05QPOeqvUMFDDpwmPBPbrELFpAyT
PXaBQ2XnLvj7SUGCVpGR9jIvP1Qkc0ttlZvvKAnG8Su9yvql6w5T9kIPBGq5ZvYr
k19cbglWhNwtNp9WjJOdQytun3xKqDZ3XeYnPaqN9spEyi7MpPOEfGnWdLBzKSEF
Im2WlqjB8ahqlhQRGjkvDz/7WAINbTc4uR4/MHj8VZ7SHEyvl+B7F5wVLF1O6Tkx
2RmW6fLYujpEFNldalK+KY7HfW9DYvGuweR06fyBP24fkqaTrFSOeqnVqqIX1r/G
K+uDIIvNpRR04rzwvRM/hbW1eBygY0UcE0NrWTlw00NE/PHrStss4iL0N0MMTS44
YGXc5Q3I9DjVf11O6+ueCqfMBwHOiiXnxefIpnxHq+WK51lUPohIFsi2PlgaZMS2
Y25kO8/swe0BhIp+2awQqC5kbFmleWYFzP2Tfg1jOwytZhs2k1Keor9i107VMOKd
3ZA1KrnPc1TO2rzhLfWxl5xObjxzo+uoFOVLB/aoPySEmgwitPzQp1d6rWAq+m9h
ob073tmkOarlFClg6FYc7YVn3pzUE4nYzvKanD64SwwvL+tP7LpA4t5r7zeR7NGf
EB5B/xCNR5qkshvqj6iU5OBCnfV18tb6ObghMue5g+E+t+Q+y6ODdC0j/RBxl9mA
C1zjQ1ADbZIncSfMbdfxiTV7MBnihq9ojfEMeeEJOcodaMo2v4uXoLnge8mKzJhu
mWYA7UDk75N0m6D9y7PaxiBhIu9rosmF1yce43lHHGQapubVMqP9UavM6N6Y3YBJ
CAb/irEi0m3cpw4+2E1tK8BbPRZXs8JXdE84IjupzryPGJYx2hu5e9/z0RX0a3qU
QGPEUXJ6Kr61Fj02NyIsT33p5vUizf/l6gQVR8XSmRjxqtT283/jZHA31pHmcJ0c
jtT55n+OmtF6xUY7DlYtPpM031Uva9u3TUM2My9ZBpx3cM2yspF3U2yXmCvnx/IF
gNhUAkaGwtl/ksxkaF7kftxtG8SWQvnFgtcwkSmO3InpGp3w3Mt6M0njg73oBVVw
Zni81ykvJUeTcfq68jKDGlGvVx1J75u3RcUZjauHYt+nd5nA7fjFdI0ScugK4xiC
Larq6V5TkzcyQA2AL3B0tsJJktLPYXXUtAVQElEyWTyoDe76CVBnUQhUdJl6Uysc
vjgjgDPj4vGTR637v73ae1lZIgdpSdAFUzp7+yWWgpawDXNa+uL1Mnn+E62ZovEn
5DvTr0u43WovoaJUjGdg9jAOpTyV/k0uvhANeUGb6GMWa9Qvckae9H2yQ5/IHiF1
C3ua58Bq3bJNWkbksHg3iIltnnYB6H0Ffg4i49yiHRhG+E48qgRlytZR+35ZZXQF
8uAIS53AhQP9KGIWQfvncctJ95Ew4aP22+shGIrYalI1JyrWj95UfUZGF9J6jeTN
c4zzvvBj83xklsjJvnEwjVgaNf1mfSXM60QGJJ85JYe17IeyS2zYqDhLWUSJX0dB
UeV4nwRIQHI0sKakrtWFZHP5+QRk50llh4hxOFeL/59DC/IxMfuO2xXKFZGueio9
A641HlCo/pXRiXB5AdyjOHipOqRUB8Gq/ZWZoZsbi4HTj9gc7OUSpiipituHlo+b
Tlfyu+nvadYzZRGIefu3ohOavCqgHD7xSWu86cEHDrs8bWWQ1EUSza7eM2hBDIOQ
QAdCrpQtUOnPGCwNPyS0NKx9I2EeoLBSE8+hWcyBibPQ2PuNeUohZVJ9vZHAgUpN
JX5duzrZ/hkTZ/rpu+q/8MLwhleJYecC/jOTAk6IZJhddiw5UnQzCFlk0wAVXW7V
bB3QycJGTKwvy6L4D6LsgESj1epz36pYz0sVs6HPGCGBifmR/TsICO2H7wkvYer2
Xmhrxi79H+nXaYXjoLn9sQBPvsPY1Tp7JKGppQf50LakKLKgFPw+HUIW0MtYOW85
1jbNG1HoEP22MOkV6C100UdfoyQ3jF65SSWjLjXvAPB2r2cU3PHn8NsW/Fp3Aw2r
3aZTTERm1kH5YLabQlu8tH4bbco0789xeJBTcX4o2649n9eMo+8P3y/S3G0yPntp
d9+dmLuOgGZ3YwWk9fYOx3bg5tobiAokRWhUyCDdgvLYZTcHJpjK43py3WAucZGw
YuDJiz1qb0Fxz0KfmB5cJFIM60LfmPkb98AEHhiPdn50K+Om+ChfHaZ4uFMVWbDs
CDhumBLW88wdvcz3BKvSUy3Cd6JE/3vxuGRUJSriqOWAHNmoHpa1OQ8Upo+oURKB
t1iGtf2J7Ex59h0Edu6u+VhRVvJ+eSWPX60wghiC292kV0dUZZaXggzDGxJgkFkt
ag/TmBFT3amedSjTqRkymhVw/XVEYJVrb2n28J30ml3VUDvhVpjGsB7WLtqNUJP/
8NTervuJimHviaGQs//XZcDgNqFyAw0CKGa3EsbEkl2t0IhK1UE2r7SajM3UtXOp
id+jaNew4L4OnjnoWat1z4jFhqjeyE5IdB61Ze7SYg0M49EFljXeZGo8ukXtDgxc
68vheyoXC+Y1YlSNxLQNPKnDmM1P0ZWhVKO61xGP7yUO/OADIo2CyP/aJhZ7v19E
bEoLXUdVlju4siWKdkkfMAR+wIng7JwWG0aNRJ2v3LlIJc+QWR0C37F89LXoXT2G
7qNypmRTRXf9XYhgfVHOQPlO1J4mRyJn/8e3YBNNvq0XH81JCtBNd9OEJ7IIYnzy
09XDCUtFf1u4S6yHpkNJ2sn7uWh6I9bLm1o7oapFV1k5rmht/Hc6G2le31h1NbrH
ziuc8ft4NzkIaPmxFQWOkD71cRoO5QtsuL4gm89TAp6RtIKOGClKjeoVk0oeb1+R
XMVnxFtpB06TbUYREaPwh8l9FM4Pz4zh3TmHEpz9qwldRqshb3P69w7YFJANlE1r
254/4p4nIteCxDUHmi8YSHPWhtKCRv4SmRYvnVRhEdJPejmYJ2ZPkbds3GggGEiG
QF1blE/3NtYg9HaK6sqrpmYVSLfplhpqA+hAHSs0AGk49JrX0qbYg+zw93Qy/T8t
zVDzc9AqBwi9puVLVcPJAGkacm5JOh1XMA2woDXBy34nfolgwKwBF7nDjnxlMl/h
BRUuUk3M2ObORxjxLG1XPRitCW6sNG4+TCrBcXhWAFtqDWyYZ+58WG9TmuDFKyLm
1QgL5cRpOzM8QMc7+QnccEEd9WtTpCffNvGq7W0k7C6LNiX6rG8vcX3504sqn+oI
bs/TN7YVu+fZ+4C8jhNvlMuszW1mKm/xO/2bpqPqsJEaHtsDyP456hrgtW+EeNdt
1fA4UQ+GYDYWWzsoXipV/9c3ZsnHt74y1v7v2aSmhTcQdksFZJam8JpiTwizK3VO
QT8KozDn0TXQoCOQhTGveLEcf0PzuL/7cQn10T+08OU1FYbX7XOTSxOjb9Ie4HM4
iQHfLnZFR4XtdDcUfzoTju7g4NOQXROWtweMI0UgriPd9zn5gpE1Tvx9LlMz6kk8
XczpYuFfGO0PNUe3EtuQXuDevpJzxatB5ustGcpVZPPGvDNBhrxKByFWGxGG1ktz
1LpkL69XTJpJekVm1LHiQ1mNTweg9b02RXkKX7sjL+Y1pndiYxUZqM5xCj3m24sM
DNd83hb4klKPQAmPW8rnaTO413E0g5lljCvz8kjJa2IFBh4ambHIwx9YInE05wnv
Tyyc0jT25/S3g6LAh0ZTrcffrZJJWW2hOElXCG+12eXOzNkjn01TwtZOxTabVTjo
8a4NjaS1YmMfJ7z+1D/3AnwXL7+mWmINuSeha8P8eRig0y+HeEuKU/g0URl5a0jd
GoOMbI5N/1+bXysEgoscQWCRGNrNkJ6pLG2d2BYQa+XwGfpQNihJRCj4AN8r83+J
N7fNuAXfZbO6MO7y/JVwGzP+9wDWLmvDKPknyEqJczYeM95ePQYJ1Ze6Qf2xeY8Z
ua54ezOwfXINFx+c6bV/vgtXz2NHVkjzQ5EUj4IZHGXjkFBIbk4+dCNHB7mPs+1P
+5J7TPlkUHfiMOvUcWlH2zTXHUZk7gEgLjseHV5ZL3ehxR1BtWSVd9p3Y8Qfyt4R
/p9Uf5C+7YHE8lkRP8UZM0SFTlALmiityB9YclkjqqnvoK5BlBFhV8HUsOQrjZC9
TujCxjyGU2q9ESErLukg7t/85oslQcmFLP6NrN+quS5SihOVf+VowVzfh0o6yKmi
lVqmvd/CfOkHxG7ZY+U2leP7+v9okdD/vyzchR0BwBiXpkYU4Zh0kQ0XHsuubgo+
E3a5KP6PYfOorbbTYL3/UN59w1AlggwauuBQpsvdtt85zA5rH7iDlNuekoO1zBYl
efEdioN/usH6XPBe1enGPVO/1v9HALk0nLHcO2NtfrLD/axv+UiPpbjOCz/U5DEX
VmzA0mVIX3VVUbsY23SrxTRjfL/xYbcEVMZOIYVRyJZh58+y7cugXarDMCSJxU91
H8I7/cS31i1ogrxlqN90ySE5QSuMQJ40Xwea7D4DbWpcSetTabZuMroOE5P+bM18
+BQMr0eiumRlTgHDPy3B2LdnuDb10StRQxzG6H3FgoehycfLRzVE1dgAlShsZUZY
jYzs2cJrsQ9jdvfQbJ+7KzZuSfaI+0mqHDyI5AcoZN/wP8RdrE12EP9L6pS5z42p
IPJDGetbcavONH2Px0X+aKb8zm0/yzSZDGqN3J5/YbNwu9lRPUBRXYnc+TOK2kpO
JQ1JtF4rTxCBi+icO76d5z5LZqY4q3DXBjlyCMNHao42n2A9dXPgfvRBRZdb3kEM
T/2hoMF6NTrAGkZ0JdVuKcU+8CwysKLVRCRQbSP8xYiOgxISGDZZ279levDqlAwC
9yebfAwGxFBRrRIpZUnmRrD2tR5kst2ZKQsY6LjOG5P6QqEmkOMJaIHPqnBEJmBo
p01bdZS5KNkAc4+Y1RhGP3BJ5FEzf4nEg/leTbIGlEBl5CnOHlCWiUgYFO/SGCDv
XT3RJihW9YdYL6fT/Syzdpu2xqR8TksX4g9rB3pCRPvnjyVN4yONXYhFDelopmJS
NrTgA2vIc8HyJUfDtpohiszhSjZj7913GGny8AUbPIROeaQyPwVnIjl41U10Rqkm
NtBsq47qJFbxl7jPv7WGIoW+OMZrjkfUFW0pWMpOuGFa40EH37yzTYl3MiMJvewq
wsy7mVN1r83esjt5FWcX19q0b/Aud3PkJUZlxifLCWU/+yPnsRReW4aaq3okROfU
I5S3FxiK1Ls5CTBFDHLHw2Ixkx4m9gRaXraKHR0xc1PraeeA5181IuPlv9mmsRT+
PDZihuC9Yfy+MJOAfYJnInT41NPoDGH5MnHYzKFy6MFwqvCQijqop+cCgHDYSDkY
J3zRZtfc7jKLqqCeDuha1tw0eIFUev/jL0R8K/zOcMmo7ZLxX77uir0NVnnnPlFG
o06Q2YDogMmO2NqAztfODdS2f5CK1jyFvqKIa8r2YainTClL7IMQM+KM9gsYP5I8
dNCS//gyGZ7yo4cQ+OQgaT++bKZr/pXcClp0YkF2dUz4JjCQNovvKElbusbyUAfu
apyxFvii1J4dfD4QhvtPLsOqpVOPSZpWEi3ShF1pQzEnLE8ioMXgC4BqckdueFW3
bzkkiKbwGWZbHGVyw7aHh9A7S4CUqQgzVAf7a4n08+zu6C+1A9dI5sBjrpB4japw
qIPHevVxqfk5O0w6ssxeKmv9udRWCH5eut6ehMglLnjQt9C8r+do2QiH0q8huzcU
Uf8lNFDeCTWFhdeOXe2ZVHVec4G6pjpXKoVjVC3VlfinOqRwgDJMadXZPtqNDsWC
A8n+eJRNs1E81hk0xuwpl1MYC/I1ULOl3nV4saz0iTUCSucpg6aKVfBKBiP0gvEN
iK63CprVy4E+c8OhPOJhH+W4dI9EZZC0KSP2Un+JSPh5pygtgFBUGPZpR+pfXemp
vqDkjJkST5XlfNg2jycI1G7kePxVb7tMtzuZ8FKCHjuKkMnwIYovRcid5UEWm27X
qfrgqZeeLfTWfL/xIl24Vlb80+/sC/2/J5xO0G8rZU3/GBghBcQY48vKnNA4Ckah
aCDGF1WtkRsj7plzt6D6nJ/eG9/SZZ/rpAYU9OJISDdy3gIQC4Xrh25CjrG6Tlq0
5YEEBCTjkJ9kGWRD9A+BP2nZymiI7YSzduw38SnDBDitMitfMyXT6V0bOI1et7TZ
qOimo4Ykz4+rdf3EDsG9ZagS3p4J8aCr16pCxrIjF9rHqqoiwQol7umVx0mXEpST
zJzYG+Qu55vao3ios9/aWNFHImfJeWLq31nG0BRpmpI7+p42vKP/i03gLMgKPwjJ
rrKCPE9MZqwpE1z76+RvvlTvWHVR63v0wcHk/+sUOBrwznrMr71w7DXafMox6Wml
B3OS5e4qzy4KrbOdvOyVlgScnXtmKyCDIJuH0jK8OFRfdNtW/SOXlWCnHBNd8T5v
MdrPcP91A0dwp8xhBlFdj+Z+23qWIUu7CuTiDCbGGp84P9e3JfhHqtbvFOsTrG3Y
3kBIGZlEJctHaJpbHYR0f1fjIznOkN5vDkDGhInI4VniSkQJYhGj1EMtVgw2yzwT
FCAYrB82Maw7M4x2xm0TbHojB73raWUVnQiFq+wSlVdTfgAJ42NXEV56FWNCqM1U
czAYLPF7sJC2dumFZw870wBVFMaINR/2Ok2Ob2YHJWoueOjtkvh8xwA2cqLGfGfT
v9Y5g52FGvmZEjLRrw2FyV2+K430qJuFUWRGaSnmwoA53MzSxV/4U+/wPTN4wyJ+
Tpiwk9A+DqYJneLwKDspMCE2nJdDz5jFbPIHzuzDZjFrSVhK5J/6nOi14HtLcC/u
cPcEzssKsHL475Y9sfjiLmfaRlfS3X00a1GQfGDC6MUsMq11JJOlBontLggmBHVP
4vppa0cOrgQ8FFM4P7RYSUAPi9DWZOf+v2nrAUJ9Kp8yAzcFVzvyX4wPuJR9doL/
tgxpSHfPyy3oe850MYDPdxsHRu2Bmha90YU5aKTvOUTpx9Qk/k0Sl391BvkBtyq9
C/z5fqG4XTJ2vLsQL5AUJxA5WN5BKYZGJEQvCYosn1aw4eO5sULwTY7m99Z0/vDD
O9OHMmYp1ovmZrMRbKXxQikK8lP/Mo8JPMXrDJqwaNl70KoV2Xs7vmw1YC9U+zOK
I+wZYJD2toRNc6b3WNnDKzXkWZP25hEjy+/gGtp2X9bm8v/1i59gUl48DSAAL8pw
gT6ayKt3tb0vMd29ZqnpVFyLXTV2zZNESTC+Qb7vkF0BrnrXojKlYk9Rl4BEZpT9
cU3pzmxxUjbDhhNuATXUfokdXGEHN3U8clVIh/i/RkGHSkmLniIAXnipAPXOs7TA
v/g83EgRhy89Dgr40lt5LpIZzid9HGy8Dkgx/FAFEO9GhqaS8EkxxLFaQd8le7SG
0AvGqFLy182KLdWIM6fLXJAso6B+Uj4ZRePVAmb11P5ysyw+MIc1vEFnnRVreqfW
wFxK6x8opSEyOXP2Akouv2Jq/HGrPyvgtZ8YkljWkUMeYiTVsBtL/3BEYH3WR9Ic
3ldWlMS/UDE8TXWsiO7jTURlrqycakACPXqN8LltIlUOBLLDuK5edRd7ZRR8WgoD
zDFfOPjrjIB996YakGondBQHcCLzMXCE1THYyKCJalHXk6enXcBpXz6dcqfQ2LOa
0MUSI2jDCbf8koecHfusH++Aa0VgDACPnlbH+Ix43d6s3EzDC46iH/x/8z7HJ2D5
7rnVyMOFIAfCeGFR1rEFDusGVcsoTEvz0qz2zHmo/OshMW5XyzolMGNPp60M1xHx
xbOWuPcFIChntNt7qvlyUEv0jq1EvzRHQLLfS2XTszuH9UMocmYo0OwJTPsAclC9
RoU4AV5M0GzQMUvDeJxeXo4vUxpYT4IDTQzLUDiiZpb880Vc1sL0DWGVpZrtLbKZ
NeXicP+WBMIoDOHLpVVqOc1WW2YAc31D5VcaoznYMETGW2K35cA/UGLlIOgFL6si
2l6d35k7JZSHoEHs899sXXgOp2CfXCoUCtOcDSdpRbhbdAxpiZ3tSLxnMX2+/AHk
d25NTZuTCodetQG3N1LYpp3GqasyBijp6YkBKsDBHawLcKFHr+WKUjnT5G/pPj/B
MG58IWegwZAheHOj9ha+8x8RnhmdjE4R5acsLgU/FKgzWjAASoV2dJYCVy5eg0Sd
cN5D+QdHIhzB/93CWaYl8b3QekNxu+OQu31p1f5atE85K8Vk6tQPTo4Ya/cRBSh8
kE5bU5iRvk3QLEznUMC21x+/BlhYXdZ85G0IA8RlRpI7uwWkbdIFMpL9DZdNbwJA
c+EcAYv71sUJyAeKBHidgNTBJh0ghRYoU1olaQKDxGZsMIl5YzM3f7zAo4tnvioG
TH7mlMZmCNetepY2sSjlXd+0FKOKjRcTA7HmxYVJNLphjArjfoDQpgIbMyYFgWa2
Hy6gTJ8diZDsygPawhF3D5pcU9qYBpMqvxmuMVQj+2NJEfGe5Yg8EH417/eWCODp
bqBxtpY+nuUIvDdhzzJrONJZfDKJ5sx0/yS7kOJ3pJGw4pR5pY0XGQy1ESnZmC6y
3gwjv3j+gqCJ7z76fEA1WdTyLqFYwvTtcGt1Wj/odn/gZ02Qn3Z4HzAm5GpiCzKQ
pQM5y2WB3/x++MysfKG4yiM7qpGt4fS60bBlN+AryCu9etpZYBQmY6ZQ4/x07LCJ
puTlYe9JQ5lN4x9s7HjqeJt9Ga8od9jb/7+svwqhBcQntNC9inK49rb7SiExD45n
t5POp76PIOAf/XA7hR9vkEYWTaqtX8dowtrL8lnKzeCbswlFTxY4nBaOTM1Mt/mI
Ez0tzKnZZkdJuTqK1C3wA8BmYFcNnGfeAGuqdFSRZDj8rCNgVjz0FlkrMzqiOz75
/BS/vVhXvIjT9zUuB13Dt9K1kYMTrmqsxjqc1TVmVHMpKzchDaiT4ZzkE1JSl1jM
FZRPbtsvST+U/Ngel5FmPRcb0Zboi5sxhT8FaOM2e4CyPt15A6kCBHco1S2fwpK/
diFJupmsGkoadIjlxxjZvGyLy5u/FpG1Eb830IolUz1yXT5IWX+aSMLSeagtiFe0
bD5iMpPZc0VLcjCbVYux0n+p1DR+fa1+ex/V1VaugsRq9nkYnFUyrLYfyLqsL0Mm
5FBsO5ze3w0w10uFiq/2DigVT+wun2jRFagCtLscnjB5a4OdkvmnecQcbE99isHS
+69SyaINX/iV/oo4HlC6o1E1n/hcDGCUVX2Hd4VwcgA4/okFnFzkbgwk19cnac4+
H2MAkR0FzFFYNAAybeBMzUq4y44mjiMUjnzAKwIfJ8z0otNDW2ZTI6w8GtA2j63R
R8Dk7S/dJEQUT96nVMW6dKLK22EB/7oBCagxUv3GLeX4eFJvEwbtfDTgiEpmwrWJ
MDPoDVa7qUmzRjUghRukNNg8lpHnndp7igoL4KmlIpRAnjR8fbS0VWw4hRtZCLHK
EStIlpJQ8XbnSbSUoC4g1mKDtLqQL6jV+nqxwc1S66qSejDlFq3Ij+mkG7tdACeU
2OZFG4F8XEXQW5LP4vvgXjOQ1iUVgoqoQIWTUOPmVsNgkZIScVknnFuye0fqeqJr
cK/VeL09PwPjGbxeWzUdSEqmrJnEUZ8Mg1LFMjM8AqJhDYDYqOixgsPV7CMTkkEK
5A6mHIMymyeCJwpa8Ag36y5PHvzxkCjcjhbGpt3VYMoZ+aC3XKiWD/7gyyofp+3L
o1uG2PyxkLX1qMhtp3dd9j/FwwZLo75h7a3gememeWFN35FxbmZVs9BvzV3Wu1s6
2A0/eLbSECcvB65Z/GN+VYiT+sw5ZnN/P70afTykdDBnIoUVfYgphMq3Gu+EtdbG
3JncSZOzmoVsAnDzOX0QyuE2J7l0HygXuk8zIfnBXt+n8qcXPPrYJ6xsDjlkhMWN
dP/krCPlYGJNa6aFlRT1kVqMmCpGtoTAdYs+H9kET6oa4ez1bxLxVdupabZibeN5
7Nez7ewwg37TT1WeTqTSDwft7U6ORTOkKmz1iURitLG0dLTmBhoUaUGKh3DPqXuc
TNtC2zqbSgrLDtgJLVutDQTZfKNMcjyzN+JkUFiEzNFv/ryTeqqFBXAeedpaEawa
Lv1501Ok7BrpCgTcwE8MrXtfkYpPgh9tCRwaslpcrrRIhY5dPMz9iKON9fspMjOU
Ie0KEBpvep8x3hPpa1J0Am2HrWkufZ0GKz7Hc9BSSg3ZsWp1QRpiMRolzP83Cx/2
7wFTtJ/cTL6OYpu6BnZCw8MB1+85x6UXaNkX+UmOpYJgIQYEVhaO/+loIqAtvT9q
Ixze2bkLqFM/TvQV1Hzz+DDH/fGNkI2vCXJIbmq8UC3KeES61WFouDE3OVYw8Clz
dv6EvRpd9HSDnIqtsQEnc9bjjGtgU90uF9+38nx9Btcil2eeTJQUHEuEMc0JJ6tV
9k+7fUeyENS3MIfqFjtS7LZJm6F/8cte8wTd9h9M5M2kIFsKIsXoSrMdOhRFkQxG
hORVdHXonRGhi8ZjnlmornQHV9i+YE+prHdZ7MJn/k8+ZI0FiDia8x7YEVVmlvnG
9XjB3qbYXpvUoKUrM+5CnUgDOJ+1emN+nmNty5CKzcDP5Qss88lfx5xla9tLYAra
I9mP2+4gxr4iC7N8VvWLcVE5WKUzErdFC8PXZPfloM+iC1taJFtZ7akwO/9kafPd
9VNITLudTlMLUCS5ez6FT2D7+1UFsKC/aoduXpo2+8Ij6THZ4MbVKDPhocXnp17O
449Wj2wX8GvOKJRyJKba9iOdFlGQGU+xjyg+xF12euJRmUcPpqqIiJQ5YMzbFq+T
gR6GhanNM9rku7Wt3h7ZTwNJEJJGdEqNI3Aici1NIleIreDrf2kPprcrOYpYxUH3
xog881Z4l22MRelcZaSLGsrGpMxa6suByp4FTFr8BtNpjhotUtJOzRgdq1lRNjp7
SGTm3Gh6D6RoyX99bufRB7Q85Yt5ZJ9ZXkX+d5HXGe/yZQ8WpODZvoQki+86Ne4K
B7yzNZ/at1TeRwtW/mZpnwpv97Q2yhYaCCGHzrHoYTcSGkO7J/qY9DwFl7WPtVP9
6aLuybYrQnHAB+tYCpr74vzuSZGC4DynAsznzg5YhQVllScqrsoiuwgQgUKFWT21
x5ycZK6PG74YyzPJa9mD7FM+bBpcPoMnCKHMVMgh2VHk8v6elmDXEoRNA1etRCUf
vn2+NoH1r1I3VYoRMcDeVKoHduCXZgRU+WfOPYgzC1l2w53oev2vek5bSAq+hs7U
ce82G98rcYHT3VJqFGccbUgy+O7L7nV+AFeabpxAYbGPL7OlsxMMmeO5QPu9QVKE
M3dzuzNnSG6iTUpj2qjoEGbto6DM4Twz+UtfLq3dWHhTZWXraH/BOkZ/VwsEZPbs
ZOY583gX6BqmQd5lYdeSoxtUVX3D8yZsxaToFDjAEq6kf4hL0OKUkYOcQQB99oWe
fGAzAPT98V0qy2e0h+OEsJ44oqCilHzA+Vkzo8DDWInPfIOTUXWHSwXAlY3MelYM
ZAsikXg7WzTp1bufNo9tIYGllJTRMso0vAqQjIpliXrZbvNEv+S6f568kD9OX0Xn
Vq8mLBgPblaO6ZC77hMRUi79bKCV0kGIzhPQBDNfiWd2+AuCn3vQkt/I17FooCqE
PhSTjCNyIczyfgFx9jxVnwIZ6OkH95rpbKnVnI/2O5/4SadAO316HMA03rjhgjVj
Yvv2VkRKZzWFVlIdKDAX7dzif0iXfCD8gl44YdP+iOaUrsPk/j7OfVXF3TW4Hs9t
1iWhPvYTlQ9Y06uXNNOwPufi75j6G2Xnu/QTkMZS05gIJnZ1QUF9cS+vO3gE02en
JP0n/Wcfh5d+WzFExj+Ssgyn3nqobi3Vg/zdv9KWdftaUND6twT1KY43L5/UAp75
pLJllv5k81XZIPg9KlFQZYlZknpZEx4VELKndzEEcmBHaYK3VfVC3JK+MK0VxBvL
tXyYDlk/tegRZ87kTV3w2Eqn9iajulzZNddfSwikQvMOGaqH2W+wfIadd4/dypGo
jETFXB1+/R56HksVKIKZkTw72poCMILZIeKZdsv6LadGNtly7JTeQuvfhU2hCUI5
emyPHvq/YCkx/7UJwQW8mMMSBAFlrk9ZV+TWPmzdqB9Tw8JnAI/YWHUFGN7TcauF
v+6hFQ9HGt88foCANM4z8ubvcV57RnwgxtHFzs7z31C9YDAHdN5O4kahhblXR10b
0gENd/UNcezVPFRLWV/NZJ38MIc2uaZ/qG5bhSqN7Tx36FAg9mhtf30qQ2OkIOi3
BRU4pcBtp+6Ez120PMmgzZC7/5s9KhvLi/i9PyF0/xl5vpIiN/oIvKzuyJAobbEs
CNw/oJUiBKxYqCK618NJtNLAX8V3OR5+gY5rvtXRSEqHVKiQpJqrfK/6mFvgTKC6
gSKpELbMenkZ+8kBEq6bmB/hCS0+Egat70ChawgehtQ4nrjzJkBdrYjJS2ABRFbw
suMvaJ9b+OuLbyOgKJAwWdOidJirHNfIyYA79ImdtRboBCYuiwwafQu2+xh8xwTG
MG5pTm5ykHYzE1hKolWth7EWB6u95RaelZwv4OSWK+CAbOUgGToPzWFKfiS59q2D
IO7b5z/E872dbbJZI/8EzCDorvt52FxbEWm80IrjxZ8xtexdfeGnPZnfkMKDILKG
zVHA0y0ofDug9rgTIWY+5cZo6DgZRu3EMGUwagfJVJw0TfLVMFFGhOCyir1R9gL6
WuztVlGtpCoLoUzaTZ/FPmJEcNTYv+EOE1BtDloLQ+uYkaYAm7uEudzon41UmAdm
KdlwccDVMqRanZUR1yFsGNfkPM60udKrK/XNHVXsotXjZQA2f2C6Cv7DHqZ6iclV
HRaEWEADqjL8p+90pauuN5gFfziR6qqoUvZkDgS1rbDdp1LUw8/ZxuAAXRhmLiuh
XVOJ6A0iHkDLh7tQ6sqp4DS+x6lJYLlBEwfWfWK2X9dT+8EHeMv/NVige3Mla/OX
fm0xZ8ZaebVU9TsEsAWsugrIJwN8PkC42SFrJGhOv48tWMU4PECvQe0OKdPdVsp1
iTSkctEHXNEk7Uk8OiuK+QsrVHvht6OSVoQAYPaIiyt2TaQECPlgcxRrRVD0+Cql
n2y+mqscbj9Dt249UUszao7loKHowVWmq+p4zFqGGHLgpiavaqLLQijptsjEwoAG
Do3qn5aZ5zNnVa5dgUG0aJ1nQ/TqU8tdNWNWL+9+cHJi0If4be4TvV2nSiqQ67ox
BkXD0GsptcaanZ1rAL3JHw4UZJbJqCmOlL4RxVK7rO/D+CJWdqih+CNoVKo7izxT
fqRCmbUTOqAWsf32u4a8zQO/FLUNfSm+Hu2eVQkavvzHcPfd2POEit5F7PszbroR
kpBW63zzOwwSjnrg9S0WMZvytp+jtWZ5Puq2bD0A98QcaCywRyHBezgzU22QBBcX
xJrsDHOfThB3PbNSYSCPirZ7Lw5Obh2ozRNkLVHLxe3+t+XvtM2cl5PnupgIc7M6
egV5vgwuB6ZYm0u4EeZkckYOpoDvTqwpD/403u5za9LWj4Cd5BVMZkpZxVSwkjci
JRhSijZ3x50x2yrlL27ObQ9yJ1YDURLMRWIspU3Df29BpZ36Nrs4yf/pnL/YsBRt
wcc4w5x27yWGHM5biouD+wLax2wrGqR9YQPT+TDeBU70j315Nw19ONaTUXDmHp+O
eg18nxBZ8/CK77Ip7pGH6xYi9MWiUnRtlY404HuAF5O+UcYhkQcyV+ki2OWfctuw
DHrC0W5lsC4wYJfGjV0Lu9VMSTcUCjN7pfY3K7EopzP2nYsKN6iwH4ZW+VdNF/8m
qjoJehu/NpeNLITQfHcizKUM6lOxuGG8M4i5rn63SX16N/mnTuPOTiHu4/BbXFsQ
AWPCkGFBurGHe0LdNaD1JcwyqD0mEHI222bRi4Nd3W+9SlEr7FFFvH0CvL40uYUX
xdwxcjI5nUGLxwBpu19hmS6z5tTk3nna72+vNXuvPMonOoRa/j7/dKsubDGc/mIg
s78pMvtiXc1L1Z4qX4M7vkp1C8ORP3d8NaRoyHA85R26G1/Gi+u2PivPYt4In4xC
h5FRyQfdBjdbvdDidjUQUWQhSejheqORuZftViD8MNsFsQ2jgYDkrsOHMLBPbGSm
s8u4BV54ln1TE0O7ArytEmhGADM05hewWf3Gq+b4UrpiodUL7lNOPF7dg23phkHB
oBXQcZUUGNNG1uk43mxz0J/kEmROumYPRKA81KRqi/MoIWwzyy5WpLWybWdEaRcL
XskEXAwGvEhMD2wCRYTDkhsHtx+KMqdTW208PSuOqu33nAZvABgWHceu53oAYzt/
uBtyJnjKyhzFalSlHo4TEH8DPRF3hKOBOYeZdinKU8WUwP9UWXVwq2Shnf+LFpfk
8Lr/1Aepgss/hmzH2TtX7NhZi14KyNm9tESOFL6xxjxoGBvHA5iCu/IFlvoUxDMf
HwdJmxvoU/aMvTKb0E7n6q/ulYxJcHfwkoyZE7Lnx27pKJUj/psqt7NuKVclEvdB
ZK5CH+JnAS/6Lqag9R7WrgatdplJxFDLx2toRfy9NbrcSmwIROC30xGnhR9XQyB8
7acpjgYK69VxdNCKwrxwrb6uZzlN6cBhT0ohvd+JIcfngI/MGhznML3H/CXpVqQu
KX13iwN1kjGR857+2cKgfExoFnLfs2nuqpxxxo+1AZhLEgogGiX/nlrzUnL0ZdbY
eAZcxjueZwy46jmWi7/NEhvulxOoD6vdTHTsQKk/QLsWlBd7Auqrjmif8Frkqo0I
cwfTf+dhtIEOqyOBde7yYRskCa5MMBVYQnoD7BnSnTf4MWHRPZY9APrha30MX18O
38VVZoN6ypRFb6Z5y/JX6A3dhODYgCljXuRRUZ+Y0ZV75PK5SDFfHjLOsftlRquz
FSPOw+JUNHdyJ/CAkXaJ7bK5LQ36YbJVrhq9GldyQmSJswvig3FlajP0HDDp0qR0
AChxg4WOGDijWp32XorcHcSlAqHjY3p1AiMwVbnYzmB2HXD60iHOhiHXvuhkHnYt
XKBBTmaj0Hdd6fR4B2kZpNcDDhxer/yVQsBZoFubQuBhcjdCTaE7/86dHNVpZw2z
3fFS5v3HVyWpC9ZmPhPM+K7tTlcnG9sSD1Iv3hs7jxtIcHIhMMQQaRHPgi4LkgFj
TDGz5RKTOJylGHuRUXnwfFwVwLANnbyU8zw3wRsX4lBT1uVIy+VCOMDLiProqyaB
+a9XCSt4XlpgzJ0SDVNu+ZM6QAumhlXLNxZUJ0utp9wiIqGi93vIxWz5sA4LiXt6
193zg9wZFgY2AHrhsq5LL5Q3ZHB6z9ESLGtLLGkPl3XRU/6RneSd+UqjmPKqHeT7
UlgtUOZlNm/gcb+MEbeU1T5fMmAw9YA9gQoSFCghO8Kq23AkdZoISJ6B1Z3foslj
cTiqCn/iapHuzdnC0vi1ifpnmLSmhYa97fpxd/lxlcyBDcZ48etqrw7sCeINrM7v
R1bwVLYlbHwrd4CIgyblKjbEXod4cqny22o48Hz4Sf5wYdPfxNEz55upRDVQ+vqw
6jq50WogKrjN8gNRdiHKY2bpceuOuHGzV1akidowbxMayRMqY5/FS55mQ4g8kf9J
Cjcg3KcVGhIKm1ocXQdVWRVwH01FytzYqXCqBaoUF9d0oD57zi3wqE6dyP273nYw
m3WgNQKqSc3ORqyl5qZ2fT1MfYEx2WYbs/e1s1vmxIfJhL2REqC9CWYU03FwrEL3
f+AoVQGr/QQMqPMS5D+XUPvszhXoZgzz1kPl8sE5aMZmzpWeP9IkzMn/wS8DipLp
Ywirx56dObmhckv/LPTbLhmVxvxNlP8tl9J0QLjKrBze4Qa5FMwfhD7evg1835vN
Rm3M1ilzcEEkZ4eF6rXW4o+W5++3O8D6B+AY78LvMmZeKlupKLlV7TiW4uJxzC9Y
cNj0p3rkG76TaH0M7NQmkIJqtRc/xiDNiHxBFPoTt8bOVCaCqSA+DQaWbM6P4x1D
OU6WAK2dPGHDYt3niIXlV+cy9iDeeh8MEKE5qsnOxkJrSWuzjlzkjxXxOTwnpx3G
lAQiGSBbmw1DYuo8O9hb6/ruMng1yJbCXFzRXZhJxWKjnpkKKFtHmyfgu5+AAQsa
FPeTECVwTpQnaI//e1gG/VY8Je4XhRg3NaocE8Ml+L6W3WS+VjBlMDcquO/d5NUK
u6p7yzKBzEDlG300njTPqSGGMs7r+5uBOSq4GUkOW3CNnMTsAXu0edxlQ9+MCze1
JLU14V+qqt3HCdBNT37PT5+dJ5wtPHwHUqHlGkapgZucprFWHCeXZyPZtrYZZHl3
Drt0K6i0b4kps1UoXqwaDABkzmuoXC23YUWET7kZBWsJip0e/xC2MDZeA9TPW+Ay
2+i5d0N18eut9GfGugzIUI48aSmZ4/JBdkhqzOI72IO27r6gPw94V07qyhHyRA3r
Cdy76Dm+cM+7eANlREh1VwIjyRtkfWVJGiE9arZrwSC1CkO+2n1yCZ+HWDjtEOKb
zDMOcz+cMHUjyHdEyHAPPKK2yTCZ+5Ffz6yD2Lw0YjwMRmQn+CdxhpgGioUxPeG+
GjPO/kIHesIhJDP+FY33x4gSi0TwqRioAxG98qaWNddrMUZRhF0VnTzM73vDFcyw
L2IVJKb6kdw+gwhpr+Fnhrm43R47A5bf8rgPB8cSbqwRTFg7ZWZUUc194GBuxP/r
WVRR7QNg8sb+ocUEr90np6onKblCe7+OBEFAl5D8R3Wuzz5uHURHhB5LqWF/b7YJ
qhmF7FkA/NekE4WE9EfUSqoetikegj7wEY6yJ+3pVXPcULgGOTS93ZcxvgKJsfZI
7aVd0tQlCcPytyt8Bef8ciuuYHH5DgWe345xzxORia4QZFpv1D4z7tU7K/XFkGu3
GsTJhFNmr9hpkroCkUbNnACMmBbgHiqs8ZKbIi+LDENO+QHaXoSalEKSwpft9O0F
vdFNW2O7hBhvw/vluVMLmRPAzJX79AraU78fXHP/tNHfHyj65gaG5q4+2u1VpMC2
Kn/hrpockPnufEfmMPeIKheKD67cx/XUlb85H+UTFS/CsyJ85EMVl+G2KL3E4bPQ
7I5roVqr1Wb4kJA5GuJiBqZIRxsDkqJeBREP6EAbCZHCNh6Ob+moCNuivtHInMr2
uysfjrBLBDpiWNRObF2VFz6kQcm4yuxcf09HPAXKWgIhAJjO4mdBU1dIJ4ho60SO
CVFk0Zbdd7/Y4MsbSsT6cMhHjE4nf0zrcCqYONJ/g2L2+GFi4LkYQYmAifO7DwV7
QkzT/nalEHlyJmZZCsj0+wKRV32woTXK/mgzX1ckcI3g7WGZ83fDypCeLj0v/a21
KaM4A1Hwsmftyy6jR/S/Km0pesu0/CT1rRFCwLjElaTcFxYlVVWNajzjq85iVZE5
WtoFnL6W49yojNKEnPSZNkD+JyCZ8uAKEqgciP2b/37Jl2wjEETzt2DiCrCHkRQC
AS4H8cxVhrPM8miGJNBNsUE3f+ra9iKl4Zd3DFS3yZdRMv+I3A6c+kgheKsRNlRT
2mlNgzQp/VncSheQA55gDMG6bf3G9ARI10umDu2599UjhLLnzV4ItUeNKfHcC91l
ToW+8yrgin1FT75JeKR24yO/kLM5OmIR66S28kbc0pKnXLPO3tlSI1IU6f6FyhP2
aYgWYJ0Xp0XI0PXHDAZJ3y8dDMsWfMNoJs55oJW/mLUBNsCfpKS82JoiXelFIXvO
QEGYvD7/vDBA05PAhiloyo9HeU0UVmJjR1gASQxJLZVv1q4mK+wXgUnqVzcFZtcZ
+KW2S/zRQmmJZS95wKwi7ULkUgX48BjUzXziwGI8Lzuh/hA9MfsAJ+Ta0NOlrL7p
Ed96zBp5Hl+A1R8IH8SL3pZxVf8X6YGrkTz5f935lJemXOyhL4UnIEljmmx73H9a
kEf6uHXZubRz4Ys5zKHwD5bKIMGiSgDpDxzYOSf8cPw9qiRtFwOvECUfmwqd+pOW
mKA+JLpbMWG4MEl6ydJFfOp+lgpNh8eFmH2M3U6xurm2ya6LHjIKzA+Hx08S9Ye/
EXsfY4CCunfXjNp6ZkVDcJhffPkEavVmbXMfFW4PX2UUxRvRJamA+edJH15QO21B
NFAadofguuVaShelW8HbPJx3ZIbHUcpV3SLxpITgAunFKzl+uCjjt+Cz0jTnlp0K
0l+Xd4mmsbViouLJ3YcddREmOsZJob8P5p8j7/V7hX+1s9G6QOKJOMkfcJWiDl0l
UOMDOYRovbBN5AaRibtPat13XNTUniXO7ccU0B2l3Hk3K5HA3/coxVMrqzDYNJz/
a/HLaQ8ZaVfPJuNDShAFpac7Ndyo0PrWAuWF90O24JfktNgbt9q02/hbmSej05FZ
wQJMKhyzps2L5KT12t0aRUifGIowK3BqmRP+uT8DuDqEuJB/YOBDM4dAk5Jbs1kN
iNus+5m43EufrH1JqTqGDkzVlL4sneudSExBQLJ5jn9yEN8JuU2WigGT7QUQY2z5
V5SCCLYDNjDu7ylO/6UJ59/JJ/y6PQcTOfHkb+5DVceR+x672SLFj3xZM/Zx6BvX
xOXfkc+w4uXxTFPYEN4eTeHnnt9j7wao4ShMhHa41HEhsH8MCsr06AtxwuiaHOzA
t5PYzOuVW8GTDIuK17wus/s9Psaw0YJL52dMTOsWELDDQ0R3fDe9GtePB8+G5dC2
HA5L9UMNBSFPoaNmK+kSaS9i/YN5T1a5A4beeYeFLRXQ1JF0n8gbtdwrexAmkXx6
8gYuN6Rl4BgaG6+qzvncdh3ph/YbMhguDlT7rgPPWblaYkrnIYN0VZ8KNB1P0Kts
XW3FihjUwANpYFlF3sCpz3xewUgg2f517d7uZUVmGtEWja9td7+ole73osMPrP6r
52b/XbDDCcPv2Nm7j3dmj8N5/gquLLEPVDbqKvzvRblRMnjS1h0YMGrSaLcNFjQw
lCbqxt1da9CzSaPY/CLuBtJFULzliptpWZU+87Z4EqTB/AVKnBz0dAq5LsZdZ9o2
q4FQ0Qx02SWNrA7iSJd6/fpbgitCsA9EBgpJkRAIehYYU0dv1InkFqz+nm5zE7qz
+JR8hcLSSgLHU/UNV5npBKxSExpgZIQR2wQi0GRapyjhZx1rp5N2RuIGWQ5ZRMv6
5KLm5CLova6whagedIsiOECNkyPv5RzxXHOG1ROb8wi6o9LV4cyXCsjEqUAX+Ofg
jTqGnI2JLxkszZoUtmR8qwyi73H5pZEyFjhoOqtLvMl8duYUhGeH8aWI1lNm+CQJ
+8UEnshS4cBpRUGyKwvyBQURu3xrQt1Lc/QkYIHBtmA9e6c1jEj8Ukq+nkQjgWIz
RNLOC0sEOVOIrhfaQk2EQsLfkwjZF7PMOaA8iHhn/G7Ice0FZKcQH6KtE8N+uKlI
XRjz7UuZ7Wm9ubxlOWYlUaqHX+vOTj5gnVkSjCkSVsGy5MeMweR/yqoEzKtaZei4
JaCOXfKZ2jUOGwDaSlDlZ5X2RHRuy4X7mx2oP+2XKep5KJslaPUeOMdb3wKn6EFx
9A30bAmwSUOZ9lo+Fvm8I1BVi/N+8rN7LvtksFMWlijTZqEqsUeC9voyuznzXELt
EIP1df2gQLSi6P59fJtIBwzRNnlycF9f5j2MqEbGyFMI86LzZ5DBG96zXHB4TDI2
vL0gGiWs9QkN3tADb1gU7n6hVDrIRa0XJJIRheDSimbCkOSi0uSPEK9psEfXUrPQ
05XvziaBAOH4OCTQH9z2wmKInbLYiMiyZ4hSDR/WZxlea7J5JnyXWBf1rOl0Sqva
qBYS0qOKHh0QUF+2eQBkWLxwHSyofnob9Yz0BoZiids5MeuAkkhu+Y2tK4XU33ID
feLJKS6tzYJQAjYzXpc7nmL08TtfUumb1Hss6I18BCvwYkOuMG977D/qp3cuc6/p
ZOgLJyGnV/SvwS1o7J2DUhR1IlUfWmCqtTaPtCyVJh2dX3Cni/ICHL2IffvvXhcO
jjX1Iol4Byu8mHir6uzazC79d47rYRyMT3B4LRQrqAuLAYlcHLGJDXpCCaByVCOj
e/HzNZ7eTBHXtzXqZGY0M0GveF52z5TsotlZAblrzH6sSYyE1YajrUct2IW8s6ZV
qsJ1s11+ziUAKDfWn8Zewo4pWLmNK9lVmTI3lojcmI99O+PwwquTFQA+4vezgwcu
EqVEpWUuS/TGC0i9eCYE2fAXOKo2ooCRwp+QYActRzFWikxel+n2XOd7hiukwbzQ
I6TCWroGfbeRp48CGiVCksjJgyvbsWn606OjbkWgbObQLFCvq39OcWMeC6Z6Y3yA
40gWdq6esv2UIQ3Pt+0WnfJjWsP7Gjt4OzwAcCfN/gVKWRe9X1c0VxMM2UKPYGpr
0GG+1BdrSItT3q7f8UTXgcX6k+ITGawShVMNPtvFptRkjDZJBWfQuV3W01dVIDko
9MsS4QhwUZPNkh9vz6ZTZmQzDvw8iNrw5fRPjXoODFD4YcJY1f4cn1EPOmlUDbjL
G5ZSEiKF3Myo152IDsBARHA9UwuY99E47LTfSkYJZoP8RCPqVunWTrBk5zfzLnFE
AEXtmUmnffrSqLUlHdY8Bd3YdKnYgUADbzljRcvsLtBbbFrBYnduqsDsAp6FS1IA
MnUGpHJ2PbSDN9TJ07nOx9u+kbLtKA/Xh8/NHNLPBSWZuBP+PUC5BY02cC8yLyW6
aAlysfzyh7TEdWOwGHl/iace0jcCTsBVRnENom0jz3q4gncSChS/EdXxURVr3928
4eCt+JsXMFuJr98CVpG8FNXKSGtpyvKmmFUNK7TddK07Czld0jfJwz09/PgYVxUm
qktpI7fdbOOKS4HTaXy4JR+jukmqb5L6wRZT/p/YUr/IEWN5IjwRObkruIzRdE/e
+ihfsF0RzyeR+tPkAHyWsVpkPKE6vkERZFmGLIOA3bnHDNbuaNyu0hSY3w3ugu5m
A231ZwFHm2eagYadTxOTBSmWg4iFznEHjRZbFrJQV+ndgyTmCTkGwIXgYmbV+Le3
1UHzJJv7Ksb14iZeJB22GUOUKb7KxD+3HL+8mWYuByNt0YsDhuP1lIjH/PHVDPsi
7mem1YDmtIzb7ghLNKQ7yODdde3+SD681mrlO+/j33DuJVOY7U7wEEqKWfJ3wu4k
JEreKxQJ9B1npTbm5T5rR0Bje33NKLyV2mpYgqDGUtVqwjs0jAY3i4yR/fmvgAJy
EtT7n+2BeP7JvoZi2Ktt2F5idHKM/r1cWs6g5zHyBHmfu63Vhy2UE7D69P+XNEtu
Tk0GB6W3CYbT9ecgudfmduUxi4kRmsyA4DnwkNRdHiICFCsmT4jsKJ/t9SEZqUdO
0uok/4RbwMjdE7C4CaANPtwHpVCIWL++oC3BkOZ9x5cbHPOwiC7zsV6E2iTnQBFV
RNi/zIV74JrwiDZqox+t+f3mJos9y2e5mQCDcFYmZ61oYjKPE81r5F+lbjHygw/r
SO3IF5LDFfoHKij6paUuBKTMIqhXKwErZ38MU+8TWS9O7LAGfGl8U+21d4lD42pQ
XI+KbCyaVsPCLhyndet6wqZTmX3YFOnIXgHuVz1VBHpQo5j9Wzto/u+c9tZjkMPI
budTweTgzIBvrjpRBEmb6IUzQpg4iQ/9dGl6Y/5UDfeSsAy4MtGeqWCFXiAf4aIv
nvFDjo05ad6j/bE7LEMIw36waPx+U2+xJfyCIUOwrllvIpBFHbIMX0a0QZW1i5ny
CrSYwctB+5uCbXrqHXrTKq2YJxU56wq4V3RdyK8GJzmyZ8Gnf5kOAUAOQd9PJ4YU
9OhPefYUu6yOCDFKyikQbeMDQeNaKRsKFsUaXuZ1cwycPYB8qnYyRqeiDkW6XLyE
Yp3OJcCZRprKMxhm/Y9p7K6qGB6dF6hN244DqkypmEyNT0hZIDJIwK8dg+kyi2bn
OV7BQ0Emo5273sx/UatnkG7RByjChxg/8RZT46Qt6wYTPj9pqUpbbMkmVLvZuUVC
Qk8rCIbzqUzD0rlZLpC8T10wySp7mFYQRvO841hv//96w5LFbidCWyQokFRgB+WO
zaW1StOG9SurclSfohTac9jqCPFEcQrqorA7GEwOEbYD9Ifi0xxYi0Tapb1hJyup
Lar0pnP+0CEd3X/7OaVLNMxXXtrkT2/z0Jr89puh7pTD207x9s7UANLxcQnDc0K8
1QxaZlJNx5YAro7L8LvvLzKgrOjjX6qfjSjG0MOvtcbPqX4gnDeDM0IcbZX9r5us
SiFGLT+BIjR352KLZIJwIBloLZAy0x8ShaHgGDb5XKKlrLl+HAKE015Pnc5rOHm9
sEuN5y4FlYjPakfKTmzpHt2aouncrnAKpvO6VubmXM6vVOXkgX4Z11YUL+rQZ/p+
HNwA2dqzQ31EmBMjaYdAIURJ7CraBIxYfgV6geuJSYegdEheLZaSebcL4dYFe/Uy
B/M6Z5wIeAEw5/tdFFb/WXjxRr8JPXPAMhG+p/wUGNsjx2aVaXC2QPAPibVo1o7z
utH+7zJuQBlpSuvjgqWbKjuekE0m103DKKe4chwjQkYNC9O0vsgfjf1shi5Pna1q
W0xXQcKCjN1sx5oQ3JjcZOBdKpOO/lEE99lGDsV3KCMmMGb7dGfGULaKhvNAFSvo
jZaHHYFWUR14EwwIdvBpldBYpIop+oWesStc/xZoNWgwddJw7QHjovH8krlN3R7F
bvKQ0arpBk0xIqrQVu5+G2p4qG5ygW7c6dGBIW6SZJ4UGt+DPQE+gTokS+vlTpF+
Oi/bXar4jio210UJTbliDny/xfz16IYFbV0g2WMg3Es9tZxb+Wm8Bb7E4uksld0x
hID6AB9mukS8bjKaPgSQwxX1EAPKQqhwb4b9qGwUEtAfB854xvtGs9XqTEhD18T/
5+7BU6tH+79oIxfh82HCv/OXK3VkcME9QW2W8MYr+SRPrwyCB8pxP07o6fPEev1x
eAvK876+C3fFANfMR9g1GbDg3kzhghojuRb3mkIrG2GBmLlz7v9v72Nfc3Yi9svQ
KzZKZNzRTBJgX7e18C1cBnmn+P886xEAP0bdTEJDAAFg3YcnvU1jYFk6KEZpuKSb
9smgeG+jHv8nM/JudUgtdDhA58GXTrsy0k2+ZiQ7FKrkpSeyPeVREE//cAJMRA27
Cnbx8dppaFijuSKo+Fvt++4zX7MjNoNVrNEtC4eY1iwfLXSFBrVpR7eFoQxjcsW4
D34xYEd/NCvhmGc6a4UQqHN5mwT8lptMu1XdoCYPLUHdaC8CZOxyvmFmOrbn1OoU
fymYoTN9cxYWQaSazadrBB+bBs72/izYd9zAmqnBxpvfv/tcsbZkbGWSy8Jvk77n
qYSN6xY26WyimlS6QEUoOr4lZl/xY8Y0bfpswy+p7SR/ylWK+qibo+gYvgTsDUFu
7+LppXWbHfWNlts1eKtqaQuuBzMMP9wk8Tsd50BDdkk1nfgueo+B1fIbE5agHsOj
YAnlRF0YzEBw/tRwPM/n5FfZz0JGxV28Sxw5mEPCx2UpSB4D3w8Q9IGwD/GCqLT/
Xpvcjadr455yRGD5E20tKDso24S9oAnYdmOCejAqB9fIemg+aWt1MUCKELYEnAG1
gQcaKOXIto83OQlXsdTHe6LuRfPrdrU1Q7+uxMd/rHRIuU5mMGgj1UADprtw4sMu
BU+kIl+fLtQyrHBgpNOkpRCbwEt0w0qhDiffghj35LVk6dNrkbJ+1gDIJXXLxcKX
awJwns2R6uuMSaMKAsznJDeeiCgV4iHJe0fg3n148tyePN8DXEMf3l8gYAWvWUtL
xK8MJ1ppQIh3ovM5f4LeNxP37ETF3R0BcA/ZL3+y6jwwVpSflkyE+2IPvUJHicfm
fxb72hhWLjAduHdqKWu2sshw9DZiUj8eRxxu7e1SSM8n0vhR8d9a4xORkMD4ebdt
Qx/CQJXcXmnOMAtM9tfalYpBHqEhTcq77CoXzNTpg8L4IZVNmTP0ZRXxrJHadjPl
pApBsIXM5l4S8X6zoxC2B+K/MUZ/4Dlhk9gHuiMLNzoDOjB00V3zPuJLYKeFwj6w
5sLmuZ/qmoQRTL10n7bPtBenJIKnt/9MFbSMDDmrGLdTfCGpY2IL2NDCk3sNFI5b
3lzqoEN4Eww1g685SwUX2cUa9Gp/3qHz3m0ImI1AghkgOjL4MkhGLCCadKmtfEQ8
xKDndu2Ba+iCP1DT5cWKLq9wLDJto43RufJ5BSLZ6OXgE8z9SFWfTZoVtVjTJEGZ
BmBQ7g2WS51t4zvXkGkh/6nNTtQVjRZ9RgS0kMNfIZo8fAKNg/pmup7g/Ca9oPzg
JPStlcILs0UDNbNccq20fi1FKtg6P0gd8Hmkfi/uMRzJJiejT7OrgTq7PCtO2r3o
xW1R1M9p2pBwEGuXG7UlkzXD4dhi/uPQh1OqgbGn/GONC0U3pDXrXatQ2DS963ZV
AmgTSRVrNqJnreikhk4osCUqtg/c1H2LehknOvHc/5sWqRAH6Sbmo1agOb7tH7mg
QrHSRwD7Iuv3c4BSqWtyUQ+gIxTHOsJJhUlpPhrd5wI0a92v0QjyQ9/tBSrIUu4d
KIKKX9tWdx3J3a8Sq+QLXxxGS71EbJO4hDy1HbD6sdsDSFQxRkpm0q/CNfoRME4q
XKQbEaoZKTjS4y7OKLj62HUzjcptF+hffhiJy/EobKJPw1CZ5vgApYFFCvwudEWd
Zc6yCs0DKuqo7aCRJKj+NXklVgPkddZM7cFiZIGmMDo6EerbhZxoha5Ys7/aV6f0
bw+HnNLW80HfUdKDtu+7QpPRwWvIY+A/fkKs+uiJa9FvVNoT4xkmZt7GRmx8GPcw
J2QN/F0dRXrvoq69s4v7wGxomo+iJeDHc7DEn3KC8diasXzeCktIvkje6/rq3v/G
EgZw531LiHxsGhGgC5ZVRl8s3Jl4u5EWjxm0pON397aUeIj7ZwBxqPe43ZqfajoF
TcrWJsSOTcHYU30+ZJmKzj7HW+qko6VfjfiNIdpD+PAyJlC0q58Dj6bHhxmAVzcu
wsiYE9n4uU+O6Qhi7ltgZ899xtrgVNv+CNEDeuW6CZcAjm5KWn9V9Lr13SU1ITYv
qy4FK6fAf8CkzOECiqXjWiL1BD4308AXAEPI8q8eZnLMaRpn1AImjwKfRXVapNYJ
3IpQCa5yPsuWMi4YNyO/82PBdbCt6IeUx5DDxdAm/Sk/57/3fabm717zBv7g/8Hl
EuPDo3uQH7m8qxU6witJncXQoJnrVU7Zoe+93VhMUqn9Y4x5SwGj+0DFFhL5cyph
vGlfXGzbdwBqh73MAksJBnxk9CaCIZnusjwbyTajdq11PqE6CtFVjD7ELzDtTA2K
5bQ6cPTsji7Rw/2iv1ltYKBKB9TSSXxRIsNwQnBQ6mVxDTfoupZ9vw61zMNl+uRS
xbDEJkOBAnmB4QRm14jwGwn8XEpd8pXU1lLLJMX2p/lQIEZhBJeW5GbsMPZIVFhR
AtgtljHnCJU6jLqmipDCAmTMvv52e6v7ScX4yHP+21Yt4Z5I6XHNfXk25jNIbhth
aSYezc4KhahdKhrWIsYRbu5adFvCbwhAKfeBh7c99KoE3nQVq9sC6bKf1+EcFuZn
qrjEoCC+jYXVNCEItePjPxdhxr81iLCRuf9mOUAgszQnfmbMMLXvcc4USR3syvGl
cynKmnv2IYK/p5/wabgoeWNq2yajEdip/+6goHAvyFCzIupgobSlrJlVgcu+MUs9
qDDwsdsyzBdjYHFoawzWSA/X7zJG+DPRW2m4+S8FM+/VLR93/SU4Y3J96W5B44G5
lw9A/8DLWh+6GY5F6hSK+33L8KpWWQRx7wBKAoMik44PMIDyVK2SvtJUy7SmFovd
fUyJar3zeE+QTJseVY26CB/0DI7nT3tHnenqdnSEPZG2Pa+aLDJtVWuFI3ZvE1qT
38g6DgBZgLpSbBUXpqiMgz9eXNovxxn3Er3nr38HgV8sOCN+S3X+iA5a7kbaFLvx
nucmBpYNF8Haq7CJ3RU4FQq7+4nQ4f52qw671nL0SUzXrNn82OzdWGBgnTHBUL4E
pzreNHGP/+N9TXJUWx1BysQIM0o4jBnsftyNLKGeev2a+ukgVfqNnGpEJNankIqJ
Fnz0dS89irdIRuBQ0KMokZXgNaTnmb1qSUm1H7cP1dt1+zGiZQCfgb83GheBEI9C
gr/omXLCLFDv5DwmBhVH5Zmli10lHHKaQmIgntH8nwBg4bECO72DbRTAvFCRgw8z
S2/EAS7qRuDGwxfG2RPRs+1Ye0WfDL7dowjxae0v1zsV7zNTrOIwph6W6+y+EbBW
mKbCjbrQTo+2nlRnhr/c9fXCvKj+eW33AfuWLSYh5qX/v+8+3B4oWhxqCuCFlIvT
tabN28TlNjNJrPpDLsuo3/4RfKheNOd/63y21wcaz9WhaMxv3tnqpARP0BmRKabq
WOeDsHfo5jnti0bt6onMtpjbLRiAod6QQXwR3M4/uELjCADbKGICZ7RJ0oWaKjXI
qNbv9XuI9ubBH72RMuLIUwXlZtH8S6EOl86kpViy0CZNHStjqPH08ezDRbF7eM1o
2tZ1Ne5sttG+NIFoHJ80HN5RtcWkGTPST6cvMzMoh2zwXtTjPPGY/Y/SXN+mcDyA
WBhIMlSqkNFgzNJuDEC0lZvM57PqsTh3EE4GoHdZDdYjmNblbxQO/BPq3vF3vk/p
+lypgU5kP3jKwgkYYukpWlx8+Bf+yc9tzPnqVQqbYfwtgud6HNwzGq7BzFDE/uvv
OjzIkajKynTRN3NStfbfYU4813LzQDs5dhNKLyJ3O/lOTZMXtT11/L7MvLQHDZVm
Jz7x+N4qt8q6B6FxyILwByIl55CJjl7yRQu35FQIPa49Gp6ifk+ffV9Nb+/UFnOA
guHu3DHDCLacYMj6Oxj+tXWm3IrCMVvtwyw8QFgxsuEiHv9yS+ByFTUc0uSb3YLD
DjzZrWQtiD7TACdd5u2uVbY0acf0BkMPmg+ynWMdco1yHEnmouJUsqGSSsg8OPSC
gE2Eva8N3BDZAH+iomj3X2L2bcrmZ985Are17Kzcq/qv9RIXnBJCZMjPPtuJgQqV
mrQNQlX0t9Myt+zF40/u+EKSEnnUccJ14WgNmwQnrz6POmS+WLWUAnCMmIHrQ786
flil9Tt9gcbWreaUGwQ5Jpmv+s+Y2WCoU27HBUckZLb7lNDD+CQrO3FtKUTp6N5H
Te5qDu3pBRjOhiGkV3BCa4Zd9skfPh9bjt5/HB4NIe9ynxJ/RdQJi8sXfDh3BQvZ
IFWrTljRD2XvONsD6eQ7f+yUAGCmlvVkkLTME4s3XsCetjZlqsjPU/vc1W961qPv
v3vd5N1GGyfSlcpCTLQvUk+lOxD0WXKcmxnpuaxOQk++OC5pGxtP2+jktsz4sRSI
0sH6OQVo7Z/MJ7xigAQEbNr9+3cO4Nx4RcnLiRCFJU2Z4BJB8biZJs9nd/wfYO3s
zHCXmdDj9QtjQqX8Yke/HA+jilVG8Y8fGTqUWzmhwPq0TYk/Gg9vl5keCMWCLfpE
MQruobu8CwrXm4PMfnU0vKJljJ/RheubFAq5O86OD3bm6cseYo/32qcAcB4KvmID
6fKwuQDClbtiOwPqrWioEe+PvmBgYQh5iS9QE816b/qMSzQ2X7Fi6IZnqoRG4rr5
OySnPVb7zJtZ5e8i50b1ym5bzPJrNXN8hgODd3zxUUUgSOTu7qaa2wlXlk3p9rA1
FAc4IfavYqT14nZzEDsWIPEuzzx3pOI45X0mlMdXuJ5BnknKy/dbLnI3JviSXfNR
etkcf4fze2nQsTiC78L/X/T0IFPJ10kF0UdQJGF9irNLpo+a9jYBUNDBB++cxq2W
JXcQkNRouKmPcWIgBtFFlQjBT/kUgyZeCMmjQBQvWk+c8cuwS/MB5VjE/MIymoyW
AZ/T7+Sib67aRJnf3wxuThdVDUZdNW303ej13dC0uM7fqkgqwmOuKbjGYRKXpx1P
UHzvYPsQ4DbGLUq5mhnaNPQGdLb3LVdsszTBGCLgCkeo7Xgi7Pf/Kl4u0P7RiiSM
cabsxyWS+HYADXa1AZKIDNjuEIylV7Aa8gDSb7BcKGimEI0KS/0IeDMw84O9yLX5
SNH3FN85bPd6uB1oeV/+IEZGtzty0a7eaRDYaUkkGwxe5qb1xnC8l4fRov4fMXbt
wyDJqBu71cHCcPXXCh8wC35qCFZNp/PjMr4eaQRbw3qYJmxTxc6gcTrJWxk9I9no
hGd0/Ckxzl/pDjVBI7VhmrbMJualaoKrgeSSbcsgBKLwIFc+u2W+LsNrX92nP530
R2UZZtmiawUi0KvSLIi+5tr3oiuLaHdt7vWlL/oquLlTaBDDRzJu8UFtkqz8gkXN
U93xVQi8yyz6hPRn22lnDrLrg13fKYoHDJq41+Br8YMbdv/xHCup4D15FIvRy3qh
ATTguFEaTt0MabXhlKFlwRh+vh/DiekwyipZhDd6VPRJqMZYSwcsQ/nLOzli4csI
QLJ8jy1612pDSskjpOiiyIO6hovCxiCHIoeUukfJAK69sT7WfkdYwO05YfWMfyoJ
dlOXEKywPJob/DDQByp9EMVCRUsFx0E++dXfTeyJBmqxTh1Pe5paZ8uE1OGYs5kV
8kbsHCGiNaiIw+YFZdW3zhJrpUZXAlFk67c9mD26HuK6jQ2C730JTKHKky8nBzNl
ZiFHSi1BBVCBzi+J9OzqoPgKnYpSA3dUWGOmCYx3dbw5iuUydUpBXylxMsHd/SgN
7ZUKhdDuNipxSzBFKDSp2+qmM4IQCW8nos9jn7TIlaGM0E/X5DyE9bmEHoDukTzl
XTtG4KyQ7VneQiYkYzE4mnYyJLFrouUhA/hhyW5e8VbKfK8G6cKUcLzyiVe3c3Gi
HEf3O90RjJitdwExH83kPDhQYVzdV1aNHL4q3yKzMl1pBEjrpE85FMA8moHtdrTa
SzpY5MJP5jdAr3E2HRymy1CBXJBpmbbJMAVxHN/ejeUU2MiE4i7tt0Yq001Y/j9j
Jw2bfIQwmUTpsR2dt9mH96ZGkV0NR50rM74BmTjRqsDfFT97wyMkpfCHkwLmrQPV
kukP/cos6iFgDlQNgR7E+Nn9A33f1oQdtxTSk2914n0ix6a5hLOTC/kjuZRrIF/U
G7RDeMtxy/WhH388a7F21BXoXarMnozqDJQ6nbLEPWYDWXTRmdz8zFU6+tYvA05c
Rg5bITr0/YLA1zFOsQR1NTWyWJ50Mwj2OfUsmfYZsm3pUFs8NlsDIVtOr/nPnnLx
LSK7Kv/F/MqaeY7NDU+/kipJUynz80b64SdQeoiakswoydIGWD/PISkzB8Em3Nga
y0beg0PjE907yz6eKGelBlh2HnAMh43jt+ny9AKtTlqONEsNVcOp3HW4CfcKF3UL
80Vc3gpI2TrfIqtJAl8AptTv3bPbd0ojpQDWinNYNJ0tzEw5hh+aphK1nPvdiQPi
1hCU8RT1LDA8dc8Hh6sWaZFo4cRaR/zGWiYHUTnaYHoYO5zTmQTutlfs0vDzu8fw
5om9ONPSNcWjnsRuuCdPNG1L0op6kDuNNKG1LtDsGzB6FCtmlwQ/y0b7+ny6GY94
AlfjvTO/Z/qkGeVYSFP1s0+tmRSFKNrKxUCZe1AC3oxTJNNlr2BJHNOJwvJ1sQ/K
L0AZ1lxqocjZPMSJ24eg+uY5qUkBjelQvxMvnNKMg8zHcgkqtNKrKhmk4NGKBg20
ZjThi8YB7TVVX48EB/beGx4eZfuaeP4L6OVA10Z6YBSaLMaRjG29+xpz9HZ2ZHTt
b6igukhE/Onu6F04d+7Y7hnhwrk3tAtxybWFM74cKzGfMkyhArSYP9ath28yxEjh
DknCmNZtHoeDqEw0Qf85q7fsOX4u7FcI6z6/yBEdKFR3vvvmI170VmjDKAwgaRUh
RrXk4PFLa4EHUhHYRYVczfv6hmas0nR5SUsY5kNGVDlUhiKtytcG+HNO2nDjgjnb
kl3XLlGwVwttEb/6C+d2mBu8vnfeg/Q+EtTK+euhJCkqbCvlp9o9s7Sc8ATHULAz
orbggSio8QBX55lqQkX5O3Pbgwxd6dlgrOON7OaEuoEGI2IpAU8cbTJgAPRVb293
TpGvMdsamL/Kt+X3aqMfNhTGeNaM0H38CydTaE5CRsfTL72GXaYTBdPRPbltAWtK
sEIr3EFr010ttEBrPGcZELk8TnEdM6jG6Zw8PtmUeLPZapHgcgTeWqJlIMMqlZp9
+5lbi6WbItZf2mgJAdzTu4qL59d4+iWoYvlanVCubDlFsnUPMRVq12eCqgJP3EXL
WNORcN/i2U9ckmKXXqtT3UHhyXo7A26vovylXoArNS17nWZuAmG5Ree0+GgmU2cN
HwWU1N11Kq3l4QmS0HrFpwAtQ0+850+eq738erZYX9JPdH31Io3YiAHqy4wg6PnO
eEKGGJIe4IzIbkdlqFNcwQrKU87ciwESRMF8kV5/sU/nrfdrG8+G+hQ3ftgm9bBa
gSDYwVOewZIjub4gU+1KNyzw5uYSXQQLKrHquHegcew2DxVhAaZUToVk3WgSIZ1x
RchpksYDuIl2ZUM69f0FlmvlfEbGP3SCi8GPBBNzf6M59+UThcP/KKeff1I1WTFn
W+a8SsJr8cuM40ZN88vv70TTGBgkkzhA8EeHLo+GTqCoA9bSoxVC80UJgHHBXXfF
dXpQBRtIHDsfRLj9D0rR5V484NR3c/Q+0YXXRayvOA17yvP46x2jdsYgsNwcwFXf
QJoz2VdyWLuS5duVIWxy1fiWpmr2CLtk2J+78qYU7ZmMg4WEFF22y4GprrbqGUKC
wY0wI8XbKX9Qw1D8BnOVNTY526Z5stfOZfDWGU2nXyWH/jeBh7XmZZv/3m1CbfJB
kejyxuIjlSE94Q7s1+EQYm6HumbznoOmm3vKEwI4RupD9SdA/a4o+q7AyjRmAiNI
P7VDEmU5Aow+kogFRWB9CGiiF/03hA2yy9m+gVAQuLPmndhOq69KHzfn9MbqRXAx
DyhwtaAbDUq3XxJ8wK5w3G+GUpAQAutkMlBcOY+Jw/34PnB3ayGMbKBG82U2Inez
R5LaAjDO1XbnHtAleg8HpL8kwc7k+hlQGNf26EQ0SfkYlqk2T8p5OKscHONpXfM7
kej8AxNMGr+lQ04Fe1FPDIS9HojpiBImbov5ZAnf/lPVgIH97jp492P9hPOT0f/r
5nH058T4Csv8oFhnUcB7VPMSlmlSAaVg2JETsObvE+o66ZKx0yS2kMpKXbMe74gs
ns9utNSkRkG/a2QduXLGeMnNmeoGDrsbnfFhJmT+gNYUz4Z00FJvi0CS38QPeNHo
jt72bc4wfuxQkNAfbi80nB9FsuLZhgZjXheZ0eK2QyPCEgJa7i0YdW7Gyztekwmm
usatKtZEKYWAFVt1tcJ1jL7L6fvmltTwrie8zZS6WTHAjphW0T7/zxdWhgx9MJf6
wSZHN925dEdHCTrqHA2BWlGYP1iV1LIux9pqIbIOpvLFQI2tuN4gSvJhA9KMqKle
kzm9CcPxKv4166aMlH4QCN7lpPflNGrxsLLIYjx6WZKhDlGpSuV+WeUUrNLQK8/L
9PXwC7ioy5F2xzQCY4Amhkv0cgBH4/0afG3RtFiM6nkbo9UkMyr/bp04iUzo6BvY
Z6ka9m6qdh4doNvH/tJDpl9ksXbl005ePiu9X7gAcjf5Z+mv0+jn8AmDAA+qTE4F
8QA/41YxHTN3KbakEg3Eo9tpnCWA458txb+4YdTLGOXRwSkno8yu7vT4BnCpGgMc
ldOQeyuBLxH78H6IuvRt7uSr/ZZVjwTBfcW7uucDSWK5ecBoAE0zF94Vp/YGRNuC
QqxYEJS7zwPJSW2S1DmgjZBHo/eR67bK+V/fT6iRaZFvF4Q41nLl+LDDSuvPc5Cw
P77RhmCTvR5fKhEDaRov0YkBC7r0cgt+8BtkyZCnjb6I3rggNmVE7J3AGefuCFHz
6n9G1rFuxgeapY0x5vY8rydxGP7vsNIcwXd0M1XbfeamRe9YtRUTRlUf3b4/CdyN
infMN8izDLgDkbNmIZiYWoqzBMmj3LvRUyeXm1XlogwvblAmun4LN8mvRTWsBhck
sQRXa/kHP2NcKKld8bRgbBdcvchp86RbsIlyyeCzUppFpMMuv+eWYUGuHvlWTAtH
lE+UqNdKTzHn5Exf5BUKdmSPnjbsUBIIfXdlu8qMflMyDjGFA8B6bn56Cb/qNYi/
f5YBPda7Cm4vZxI+R7gfpb8/NW+0jL2KE3vWsdjb1sGUIDrQ5dTVHnDwr0o0c1IK
TgeiXPnwVV6u+19AYXyyPugnmO4FeMcX9UUV4U6aw29EVXMC4YqgirTXf7xb/iRg
Pny6AZiAx9Oj+PYeJA4fUeRLcuOrRc8cX0v5A5KouaLho8Bmt0XDGtqku4sdH8cB
uiPvPYBvqqBTV8KE4R3AjMnK6YiJb2iYc2esL6EJ21e6Dwa9udZ9ABY2hDTmp4NQ
fPBHwYDkBeucfYMxyP2tXSjjAfCWQ1fYVl54D5l/My3X0/rBzYjLPGgUGJ9P2uYK
DL8nwEY1CtzIpLa7ZuhwIvjWQ3jI4U3xzLlNoSyW+Yy8sdFvBXPbQzSLz+igd9Tf
Aa3U6Hme/5aJ2w2YhyOgTKpyy2W0jxHCW+jxyyUJe7wbzPxJftT64BsbCgh+ZZQx
T4uroUcpkmyeOf7+FvzfYNIPhtWRcKj6V1ReLyhc3aCC7PcmK5TYujn/H8SBJeHx
E+0jCq1ays5UQ7Ppl1b0HsnNjqL2viUQgruqlMjK8J4PTl+xiD2Dc99OQlNUvPEv
ekbLh7CZ6eDmxAqr0bng3j+afDiv/kk/IEJB5zrWGySogH15K5mxOlU1MO8avawy
a2CWWrlHiRud9MiQ6JDpQw3nD6O0GhdaiaA+eSaIVYutsJpIpzhC8tKaEuxKo2Me
gJaQnNw4AOwdE/GN7dMBOaJemicVDkVnwBCvqsxCWbY4hTYbo6xiMvQyDPOQ1epw
IxymcjrYwZqTcAMLIrVFpL+sG+SQMrTOYGfGE0pVBn45HUh4yg+2kmYvExH0qScE
tyoRvfRrnrussq3fKrzExAQlheO/nAscWixnaOOqf3IcMHISRQLfo7OUm6OPcD2b
LSwormUnGsTg7Qh9cxVUIhghowiUb5yp6jGsJ2MavECRaj0BUvs8q3iI2GVoKTGp
e1rnJEs93rr9VRlzfQMny2ni9zMKeAgwk0KlW5iI0XR35/lZQc9zP+PV96Nlq8h4
OCFjWo2p2rQsrS4jH4pbvqQ8SlbTCanCaxffmlMXaFX+1Q7auCE+5lR7B9b07A4l
qepqDFe9HWKK26dQgbyylb93MJ0/QjxahXc7vLcNrkYoq+HslnotGKKgaYEntG6H
7Jc6VjYhg8SZLzF2Hf7YjHbV6rNYsO7gDg8V/sYGTsULHzH+OnRsgaaEeihWyg0e
JsJMJQ6AaLnarzltIyJl0+ddzUcPrx1FAwTJbdqFFtpvzW8Ql/MEIoddi4gOxP1b
Ooa5WU2ctJF5ZiD7GGZ73wKPexrWGDa8cWzXRsrbd4rO6LEWoqwPynkAOnXRRRGp
ei9ysBgqom6GZtUAucEtCQ4gfVWSIowzApiFBYcuETQ5Iw3DZgvboB0n62+kiABa
7UE5BRBKPfJ3UxV1GvmQUP5e56HfWYcMMGwF3Cw2dCj1zneeCn+38Q7Kgh/Yn0W8
xXxMUDqKZOFCS+Zzqb1sSX6662D4Wkrphmldggtdf5cypoE5hWhPFdr+yNNfWPmb
KSZ1URol7SzM6TNcM3QnrxpSSYKleMSk5gEx0wyQVJcPdXqQMXQHzuu3gDkWEo/l
4dHQpqWIi7WgN8zQseKk9bk87nhW3RwvjnYHaMqMBvb5QuzXtr7uDlekDpP9w09G
5k2yRhYBekUollhEYSM9aMyodpqqq4O+yDj6OYog2cbkMnp1XNcDa1YZzXx4LEjz
CnpWkebZWnJoBkinxger0mvOuG8+bZykVSKLyo78O8WzcT3MWGo9ObJXMY7uJC/1
2lJRrucA2thiWSYb//8q1jvLIy/F5Syo/cYODC696byyMTeuB5Zdyxi+pnZ2i1fs
kCL4cWIIe2zQcWYJf2cstvFo3Vtd9GT1fqyxl+6WxQhMOtHCC4sIVqANernplphS
NveFt6k4xDKgxkWWe/3CwFMK7rok5Ss5QZKhNKvNeHM5zpWZHbvENDicXCzz8Pfu
KTbl9BNlStRtVd8qvubRP5ciZ3g03HJYrvH0sYJBim9YhrH32rRPzbdBnW96X0S+
qYkBZ2iDyYj/NXBDg4eA/4bI4KT/KfDylBPu+hMssHDW2kmsyEgKFWR3VLS34j7J
utKs+f7qIA7YlWmQDUwQWzwpNWM7qPJ/XS8aRYreulGkqYgFqwNaOxGlab0xMeyd
ZoATfNqDLxRMML15AJR9cV8v0tprxNaeOevgiornqkOXxfSoCO82/uo88h0FTsWH
EX3OKTuVXoiVe6WFU5EP3sMb8B1WObouw1ILm5W19Uz1taxVRFeINf73lRUkjw6K
4B/pYyP5wPvyKussQeCJOjzpt0I5/WRxsfXzWyXeml+OoY//F0Kwefqv+U36YZNX
04xrJRr1ObLaBnq7HAqKxw4vH2WsT3oJlKl4QqPhk4y6SgD56xLzEsflTvWmABBD
6y+KXs5iP/PW4eoZhzHrg8pxYlmTmwgcDV850vXNg6eoKGAEHL+SRLe5+0GrzMwi
bGSWQvshy5W6hOCPQRQvzyJJa8jvf22CgXRHITKcVM2U1N1v0GcPvMbOQv5F48HI
X0e1WI0wUYUy0G47O8xRADD7WfTq4Cr3YSjvrxHQthgkGGP9F0AIrYS070nbtaN+
qYDYf2cdrKOl8yFRpNa2XRhGFc6dK8WhRaxgMoQAK0HBTZj+40DVra+U42CVuvJA
qtrPn9cElSg9QsinIWL5r0wu5BxcU4K4+gh9A6j57PNGVt2Y5K37ZFvxklpcgu0P
oX5G4Sbtlv53LNZLvHHlJ8eUEKi3//6JTNlx9BIXkcDikRZClMuUZCsBGm0BMm0m
XjkDkBSvNMf8Yje5Gx4Jz4/VCHGszlgNDPRmp+meKA8l8PJ4F0VP05RTYKRodzBZ
0NygNgJrFw6famGykt28IZQ/743dK+CNO5f4nT+Na6p2kQ1HQDZ0uF2qAxjNE5+w
Dxq9LrSzoRfoJrQ7VbC2ttRCF7ZjEGPWX8XeesdA6gSgC4G2XYmwBtQy8p6grmMv
HYVdeUh9aaZBPvscRWxHGeU6HsnmHXZ6ZWoQeJ0jTwXYk9IR3Pphk46X/FDVuKVJ
rwYvHK/fT3PRg483q28XT8bmhRaOHTdwsRPELh9LQEHuycGmfNGl72/0brFqwN3W
nDQzTAzfSDrgNMaj2x2PeBW/mM8MAdg3LJrv8eynZJh+XeeYGQp3vt4CmdcwGie6
D0YEpOitGvtT6LhdyfCNMlDo4Gt2PFngsjM+GiPgEjJsi3tB7ViMzefCDt2yQGjK
eNBPesewp64Lj3VZh1BbeChkINml9Oxshugnl6PpuFGK1KJ0rg17Agj3G13sD4bv
up6ppQMBAc3PYWgUDyu1/dnglnUTIWO/NAhpU1GkaukEDI02Qpk0u3Q7XB1ATt9w
wiYkQSJ5Gh8mmQkOotVMjfsX4shnR6GFxaz5BicUHs5N8D8w8BlIjb34JM9cplDC
z4rFq1llG3XkvxC4FsAzl+/UGlN2iFqSttoxjKAtW2Car6mf4DZIXVih6gxEyYYc
V1UZpy/NDE5WTEJ9/UwgbseQmMu0yF482P9ReCxUjTUDmBH3BPrTxiAXqB8D2SdR
EAfhpScZBuRfAGLBcRPg+z+DRhY8QoHq7xmV3JLei9uK4R5AbmwsD6XyYywkJkty
OpQ1LbdO1ms+iwOH1lII5a6uBnSxgNy76n0PaUmslkRos4O9OydjpvOH/yS5YAIY
vswbNT0Qwj1zb1gI1+S4A9/8QLFAiH/oYVa5jwPxRvF7kfvo2mp3H2HfbmrXd9Vr
AK6bOQMnSgUa+xG4CIyVP/5jkyIMELJDnbjI11YUj5gKWyhIdCLy+MZWt54icV2E
dI+hGmMewDwUl9WDtqK9GvBz0hcQqF5JQwbgnD/gJ8zwQSK5PxKHeBLhnba9Og2A
fB9pzNI4yiQUYZXT+RWxpjOOClHIBoPViRso+Uhur68wgN06tcFJpOaZtmVlYJQC
K9Oasz14A9gstJ8a8z1wFKm6pE/EMgL3ghsw9bg1z9H/VQtQZfVQWeHIcBUk0Ory
Yp/3BosgVq3KM1utN4SnOHyB1kwqlgfdNCPJJ+7CiCkY/+n8qr1VvLbM3viPOczQ
j4xIQKjSQ1fe45649IYz+31Da4IOxc4dHkA8K7T/nx6AESqi0bvIiQJIxI3fO1xG
c3KZEeVTAmXik+rP20+jB5LzxfKU+eJxuc+7GhjnAXGnXEx7zL2duzwXRoeFTZdt
HYJVTjzJSPXMzKzmSnZ5QOtPG9QOQ/yCvmudafBfhFXdXtCVp7ff4X9ktsWQrpRH
4m/kb2JT749DWM70qSKEznSYzMO+e8ogpvslFuTwIyqtIYj3x9Xmo7kPO95DyuI5
VauvsQ6WsGb0myyW0M2ZLyJuLi36tV0P5eVT8s67DBWuQWzi1qhZgcbDGQ5LiS0A
7xutfTAMk/ZbF+72/sfOYIclVehCegpVSPG3ljJB2flZfoRvfY5t7zeeZXt3oyeL
+hIuZB7HeK/Mdq/o2fsNgfJrxkH9YPyblAv5Flc96PuNfrF48Rzx9Ob4hlroMzxb
xzJqLcfHcfjKIDYb6w0avDC7QnrR0BqFglc5aIjYhkWeZLFySvMntTjgevvnLP2+
B1Uk54S4LuX/l+DR6tGjhMgQGe69S65VkhP8uGePgH8CjgUkhQsAFaqxiTVvM488
KNtKPtDxGikLh1ooiItDrbchW7QTiEaPcqZxW1r7KBafoc4VrumGKSaeUnnLru5+
MCgUWCwF5GdOPbKLxsopbB4VbTisgV24DlpHeifv5mFl/ng+pTZaQM47bgrFYJlx
KPqq87N+Qmexp5R7DbIcn822TuXfqeP+d/gqhy5LDmy76LVWf4R+zP4d3+QWgGti
V8qiNRDyIZ4sC6SrZWK7aQQEhMtP6k3NxXNGu6CHaYblTP32Rnw60xcVfTwhDpiE
JZf2trXA83d1508JSgXj9PtemtL7An1+sj/Y0t8gfnsPIjRiv+nDimC/9zkz6Rjb
dNdLGCEZ851C9QkKp12lOxltWzzTi335VwkGTd8rENQe8ZQ3kQXs5qqhPtqlakkE
AXJE0p4EizkQD/ZYV8ZnzO6nlgbGUPvJ/F8UEx39x6B4jEk47L5jbDZXC1UBT79v
tuRSXZsy+M81fvmcjKpq6X1SZWTsmDMDjTnU2anFSyHjoboADPdnJUjSa/JrBXuE
2Kw6hczfBsn45NjXQSD80mldc6Q2iyCyTkkakGBQeXEOPHDQIu3/EkNNX/pSdAYU
/XVLWHk7O/zAyCjmD6xnyDvRxlZvmYC9lq6awFI+63ZWRC4HvcY84vYGyDkzVtO4
gO7MQpbPftiSoNOmrTSjVtJCnpf5Vhl22P4ixXnkQQBbUwM97bUjJ7pTEWcKHn8R
ulkNc0wRw/PO34pgQMLQBapWsRVEXxs5h/Ic7mlLP7SJ9IjWoU0y/k7gwJZZnxJi
3hlDZlPQjlZzpkfeTtvYm/sCT5QJdmaIyUWNmMMvwq7JOwawKjiZya7at7+YgA5W
Qhz9GILlbti2+tVCtTlUOy2hK7TwSqCVyYd4er0hDRhJO+zf/uZjH6C8DDtf7nxt
ZBgBXSYefND9vnDJSfgEYgX5MXHQSKayPcOt25l24BXjm0EhKDNh2GWCzqz3MLWG
cgBNF/ENCiM9003nQ/Yy95wk6yIiWJm+etTpCVxDihP2ibQMaEpU7WbDfZ6/KJCk
ATvjh9Z5+U2U/FVfS27fRQKcwL+4PE21EsZVKFu2SwwT01UGNHM+oGttbFBJO8Ie
nJIPOKkzRn++w+IU9oDSDyWzHrZuoijPhTus+ovGQQV8z8iB2O2X379TMn6DhAvb
XIyBzhJ3HRgUO6VsPyB4GH9QbSEubXBUeziJPslU+QOu6M25jLgxnsBv2ho3+xNH
m/Vp/dzf0NdcW66v50lFM+E0PFmmbqS2NCGwJrmMh+ajV+p+iYd89fS6dBZEuBun
vjzmAxjVkDT9iEiYacxSqmpPOlNh8wAkp2uxbYu0+E2wOm8WPrNe5fVUhnF2LF5k
jaT/kIoI5Z1FQE4/95On8w/FPlh980ZiVMORQA6vmHBtkc6G+7POUocqLaMPPeqM
RgMqUgL/XqcUY6ikIPuolKett3apK6xij15bRI8ZChHAXRzZ03ZD8oaD9+naqIpj
A0/WZcI+HT4k/Yh370kWXasopIhHXNoqIGDuWzn0FFnmM4j/USBJK7O4uZSIQlSB
MdCxI6vxJr52uC1uw3zExMaHWoLoFVNPAOeB4QauSp3bwSwoCnyA01oUWvKiDI3Z
9womZmSp3PdF325Lkek5Sqq5j/l1pAx9x8fhF5c0nSSpoSRZzSGYtt6LkbZnDv0i
mAEzVHZnbK92d7GWNz1NphbxrM/iCgFBSG7fbb/N6MT44VomRWz6mDFLsXbQOqwN
6Y30XuzawkW205GR6+CvWSjV8woRbTHWUc2Jub0pqaSkmDLaC11RkeqvSgcDIj/W
B93LPHdq1+g5YcmH6s1j7Q==
`protect END_PROTECTED
