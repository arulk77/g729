`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42baTleneWOiZ07imBxpi1FbeuUBovBiPtTkttfBvjZx
fxhWvgTu5T8OSpbg33Sg63LDyzaKYKGUImP4vpC/FyR4X+nwhSoRw576Zcjvtbib
vlk+rsxBNqlOg7owFjyk5liR7WhSU2IPxpsIrMNG2FWlFnFgzyEZZlUMIbipki2s
2Ej2BXW0nNB2XDR5lBOqoRDJrspPUfRwQn8ijalTYR8uBAck9aR53Hlw1GtVzbSW
lMuX4vdeD7juZ3OvMiPFbGkTFPMiDwKShW7wvIBqYzivRLLz0aS9LlwHMrQ1vu44
jhjsEvGMZC+BNeLfcAUfxUTSefhHZLQOHwQrnTGqzCFwGF34e7ySei/X40NtTPNc
13jcUWOtisb3KuTf4wsXjQ==
`protect END_PROTECTED
