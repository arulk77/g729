`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47VG9nI4O3E41XwY/C05Kp7bimmjYp02d/41KhYSlQyY
V/HoBuybMDFGuJbeuibnzKls3Hv/SjOeEbsaZP3UM2dW5V3QVL7ys4q0Jo2lN2Lt
hbDhJstbWa6kN0FtdzdrEfG/ASJZFKx3+rERZNOcW25dbjf5mszi8Lfgfqxfu9YN
l121kQUSSCU6VHCwqtKrebuRLEGzZF0OrAh2RoKUerhHkr+Ici1hk3JJP5H3s7ku
IPLaHPkQN32pm8HXoFnQ1oo3maHK7gpidF2Cx+3Gh2sWxLB7/U4Y64cXz+uiT4rG
mh6yLcQIk0yD8rAwNCDFooxYf70A0pNLB/CJXonOoveHvDUArrReS6UKjHhoG0xM
U9OIOB8mQLYr2TzcRNDwodGTl4iMAjevbjNtI17gEvqiiuWGBeMdyCtaUbkoFVss
ZTjkfe/GILBwhzYs9/TdcOIpczjbeyZ5CU+iNAskPf0deLPWyv85JX6XPYd8pIec
`protect END_PROTECTED
