`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNbKMVjEglxeHLok5D1rh6MXt618vx56nj66tPa5FiQB
I94xKFMKvrI3Rj49RPOnlhAJ+ZahEAI7nXT4y9Qxc/BVQa+je1W6pm8nHjIBTOaY
cwC2vRVT4tINqzlIimhdbrVadHbBxFm4An6HYqnUZiSdBynHp9AMRuYZokgGxJre
OS0tcLyNF3xorC9a1J/Ic371ib/aJFwFT9XGPNxRbxCfBXotr6f5y/1KobgBrUP7
cnN2wlKnFxMnaesx03urYOJG9mG8ZUILup3KB5HJBcysDDOaSuE1mOYKBBMZrH2/
lupKJRQ3ry+gGBfaX0Ya47oe+RXeBv7e35diaeQUVzIK0Km00HRJlfg+mJdu8pkN
n9Y+wABtAtuRinFH/L5noSUveYVNGcT3Qs3q02v2oyRbFIqo4YfcTrNoyu7cDHvd
c+ALGcPtFNdRtAV9yr26aNaMimuy2e/qeER40r2g9WYV104O1SoR9rWsz7Ie7wfP
v49rWA0Se79r39+wj0PgvIBDGRj9MflX8GI3jmzDYG4/fE8ooKtF+KPYm1R8SAYy
gOSeEazJixUC3gqatQ0t8S0g+RITBcKK63RQIcRaRpcjN6t5hWaewDZsczp2sSNG
`protect END_PROTECTED
