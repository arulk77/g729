`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKh9OhgzasBJcWZ8Xl6AwgWL2caeZFpPoG8y96Bmefj2
r68t5bjxkmGZ1vE1Gs62X0iglX9LkEil/oSSBIqUBpWjHcaWiVtRa8XmLIxNhFaJ
7SQcgjKMOcLQmXus241tmrpEzc04kWkDt9HO8U6vV+tfloeop0y25kRBU7/uGdpy
`protect END_PROTECTED
