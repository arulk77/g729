`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAe2SF6GGWeAjUVbaflFpsdznGL22u7/XCr2ucJvSDhU
Ut73em7fwcL4OT8WcFb5CbRA8cBs5jr1aMXgEJOxzAS0qWTxjsgdc3CYU2KCrfLX
QJIr6reCxhc9NkG/IScl3a/XT7l71NblGJeyJNQ14uFCxE64KkPmCoKyD9hSwNea
ClJWUsS0uePez2jsrRUq4QuuIn/UUyoRBQxwuDhntLOAih1WkBDgEMsksUayC3cC
RLy7UbNQQrNSSKUgU97hYKsichgJqxN3a7w/KPRuy/lLn5am/HcnYa4jeuWH1S2X
Jy/WECUmZOkyWBrOm/98OKc5CGLtqHxIpSKgeQjwA9uTvsz/jPptXoisS/p2JoG4
lhbgKG4U2yX//G8jMz9i+mJvAOwSUJLnfgbK+maEBrzKmvm/pNlNpHzZJvWRaVgX
uF9e8g4cMMWPfElOHVLjLfX/K22/94xxc9fasQx9HYfakQcpcTsVznNT2LuAUo6t
rGXmo5Nod5qKwfcczOhdWYf+4022l9btqZEQ8dlEDz3MHhkR9rAtJjxrsw646OZV
lC1uaE1EC9Ox7fzm9TbOROmfOHmFE1E8yIw5gnV+0MlIk0YWzNIl6wFPMUL3ujBL
BX1N5YEqBv8HDDgbClfhXH1lGezsfxXVOP7eG+5lgYnCNNrIL0E+wxScpgCo8Sjr
`protect END_PROTECTED
