`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJJohN6R6NenwQ2l8TEnnQWkB/f2ZePP4Yu8Unj8Kjpm
DRyoS5jiB8CSBboI7/pHSKh/iJDkpGmw60YPsV3ABVtY86w9mEvDuymtl7JdSK8G
RQQJuJ43XVCROBo2OtBkTleuLSzScdOzJLtotOVyeetDoQBNM9YGNV8YrMqc7WM6
HhIs9mJadMR6HWH9CHfj3MlVgtRfbaFTpsVwNMgvac6sKz0aaJfhPX7YkvCmRfSQ
Qdt5hJLM+ZkH65dxMEPhDDSe4IHpM0Notgy+XWcQ0O+CkKDT2ukMd8IivUGOW4ui
1K9xHN9IAApGCNslPkI+OYHOHKUT+ZrIUwa1NHU59tQ=
`protect END_PROTECTED
