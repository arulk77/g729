`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCXztt8zAEJKTP25Vw6ZWrgZtCyh78wRnw8riB0ac3re
ZllOg69jgkw9RwFMi7iz5sVayN7l68XJgwBITJZdMcfol/duYcUTTpAfNuUIP9V2
5XxskaN8phCqnU4Tz/kN567mERjdNBfOLoGzbn9F4keGbn97w22RLkEA2WB4+8BV
WJd13Ge+2TxR3ooVKoSP4chWnsfK+s6nYqWIIRds5u6Ktni9x/FE5j301A6r5PhM
q47xdsFfvAdBKs74o5XXrA==
`protect END_PROTECTED
