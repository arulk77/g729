`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNwfMmp09d3q1m6voS4MB8ZknkWGkuy9USyVBjJSCoVV
z6mIAN3GgOwAGQBV10Zst8gyToJUKYM+hi4vQYA6OQZ81l1vMWdGzk9hZwE3fQ3k
NtEJ1NL/6JinD/uyB5wDNZYhhVCcii44XVsFzGbwUUpXWnTLgliLvX4Mj5Qlzxxp
fATtSrB8rAri1PgdyYew+FV63Zu2uubE8wy5DS9wwUo0mGhKfj9jiBKQ/mxHZhDg
3MsHbnaJEpH9oi+y8MYnnPaWtmt4F9N1pOA48AFhOFa7IH/LeoS/+2L+kAfXWJu7
5s4uJSYTO2qIAy1/tRS19DJ7If39RM7ZeWQewfSNNiYYmC9llN80oVvXY2Enm3Az
PuChMEFrTDcaSkoctyLiAGsLabURAb8uYxO4nblNeu7lR41yKYsRQlzNb87wyOd/
AogUXr7g9fLixvVhn2kf+EU+/OxHXU/KRJGnNO5YFZAbi1omDPOPI0Spcr9N6niC
AfjfTRzWUvRwlpRIxnNznuPuDD9w7yCraIT0c+2u1cP0c2wS0UaWYlOm1ZfVVILo
VG2HyOseSzheILumW6/81A==
`protect END_PROTECTED
