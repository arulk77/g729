`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aRfHAkGo7+8VD5pQW91LEpmOjyI8a0jIlULOu1ryNa0N
gISC189hA5oLgdkVDe4/P8qkenshAdNUaJq+egm8iFznpT49Ax1Z9v4E5STfrUpR
X1mBBTej3n/hXz6ArTI5/TOBii9oSx/zuO3AzCgajIJ67gU2Unw8efIC1isQC0bC
WZja59FC5YS80coCnbX+kUxvh/f0pojVK5vrOdP+whF5qYxyMvjZcSJ8MfcY64F6
gP2Txj4tfCQ1RFskiT0A10RcEfyFjqclU83cVR3hMSlCslQ/KnnwbxiHEB8IcpWi
x/SYw10kTFnSO8QkFtKefja/e7ZH6RUJLoCIFovQA/GnvH7FHWoyRocv+d/A1RtW
8BnVLtw4F2dmNjMdM/k9YpgWH7Y/B7nGuBkwkgCDgiyVosRdH+/QAezCFxor05Q1
3DSK1XvwbCn+EkokvtCdjItCz/IC60NlT6Wu9XonNglKSvP7tVhK3dXkije8W2dQ
XXCMETgPHttSF9Q2KLe5c4NvkCGYGCIpIpx0Mi7rWyoGkANzKjSjr1VjMzgpwOiB
TPDonFovFOimQscIYn/tFlqqE8c8egKsZFxMWS035tc8Q1zug+Vh6Ggr8qUfohCH
`protect END_PROTECTED
