`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
BZ/ypQ3j2ajQr9xqu7n0Z0Dy1XmcYicYWLtSUDnaUippV4+6lpmNldn9adw70PAt
D790z4xXXHvSTXq4OQt7KgnYZowGqSuEMj8EJ7icc197IE5oI68t6PX0lfCsmPEu
kqXY101IHx2MpcDiyYZg5pEKFAWT3fRn7c2z2OwPHAJMgAsoglZd8lNb3yryT3+/
pkHnP/x0rQyy7hTr5jSRHsD5EBS7v6ToK4E32UH3ytg=
`protect END_PROTECTED
