`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
nMV2ol/PWO8eqZvX4PHeGqp6068Ycb+FEjAoyOYLgIZF/+d1FPTk2uJhj0cV1feh
h6pllCYN42JHkgYCZfmpEpXSEJAE7ubLJ3+uJlTDeuCswoVc3Ogm0hi+BU4MD6V0
IZFBiBZratUqs1Qw40e9HMYwCGMVKNNRODR+K56tyaz6bLu+SXAvKoamwLoGudrX
fhzdkNOitEIXhvL8F+9o5z+rH/DlXf3SLnCfAyjXgTtRclncP8zg5AY/CfFVufLi
A/z5ae1u24xplYZ5A5u1Ti4nsv8xG7WVrpqT3ONdYMC7Ulh2wdti0AAsbz63wvCk
iMk8exU/70Ie0wlLnO/MqNcXdOMGXFnOVNAQX0NoGTnrZSycolAfQGWUdkiNJ2cx
mgz7SY8hoJNCgyMNkXr68J4NvVDbSRDhW4hyPgfs4WL9o3TrCyPS7BVXS8gOtHTc
247oa9H7RijZVUZenQsXKTIqlm2yN9DtJK0raNy3xIh1y8kdW02ALibQGO27a3Pa
Aafvl04NLH57q/D5QutI7FHmle/MOalCNdz3alkT14JJiY0IdH2KNGr4yeeP4t4r
uaniyjwhcH2Hm/kM13UrZljK3mFZUKQFIkjVuGVC6IksMdbiSw8dr/qsVDWU1XBq
nvonr3jNPNovOXTfRY+iGtfLmMuOKIwO++IZre6UnWTkiQgSADPyVyT2wC8zVkIi
BNF8oPIZoVrLaTZ6UIbki7sG6kZYauAbfuOqeS8RZUv0VN6PJ6vcI6lJ046Ca+6A
UPjFg55A3Ev4A7lyAQuBPLHgMtasqyUDbgIu6rEY+1mhKSSdR5IFFvV03y3LHNrz
apNsCxoZ+yDluAcEhV28fyw+LXhB5ttbOlOnwYEDsgtQpfSfN2xBaeiySXDg4msd
qXB6fo0EGxhfM0gPJAOi70UajJYrmV9fNyOj/DxwmuzpWo1SN2UT1xxZqD0+t9m+
pvkh4DQtK1r4OcmhnvpCMBxGDnOgI3KA2RfgROLv96tUaa8R0c2k+Wh/k4KFvwFH
`protect END_PROTECTED
