`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SaVB79dvnbJ0GWENU0coCSyZsGsy44eBJ7tR0VxhXN4K
Y0N/3MKkVVYhzZJK/JeFCQOKOCvZfQbItG8Q7fe9C20V8r+vFaICokvWZKKlXqae
4W5z5rFRXFPxQtPeRBPTS2UzXd0v37gPnN1HHj6ZH7RY/0rVH/s58cKLN+4Dc5EO
1Vj3ZtbtaD5uQ3JyKabOulXT84EJ9jMZ5bUg1Syy175ep12AY88fS9IFRU0xscPl
bGHRP3+1BQCx4r/2AfgYvwQHht7mhHkH5Y8nrTwpBumdYVNIU74NfQ+W5DryETNn
BUbzkH5KPTp/WjPo7RvXBQJ9ZIZg7ww1OGcCYCGbaye2gVUmoPVhKoINlqI27uA/
gH7rWqliGeB3uwq2oX1nQa50Pb97gkllN/dZrXpSKBKO8fw+bafDT2DeymB0mp//
s29fmiQtKZuLN7Ea59hKKTcw+LScnpXb9QAH0COuJVYvMynh+xgMtAualbrty7cY
Ez73Fto7gp32MtqU8Ndg6A93BjkHn3rAZ03q/M4TDKZh2wXNb/IT5dKYF0BtIakE
xd6q8PfCCINvfTI2cc5JKtHkFZppkmTu2fZ5PhSQnHzWilEPVgkgEGRZG1JJs6zS
e6vGTCjM5AioxxeLyj6NtDzdK8XfALXqD6IjMRLxk4FSuoXV+oWNDfHriZr4UUk1
P8ZAYJkWLeNiDeJcjOZjMJzqnJ87DAhigFn/wD8ucpr2lTYKrU02NNbPmOAwICcO
52KpfQgYRYuCkKS7MSzH934pa1e/gnLgQh4lQdI8yL299+mabkeFEIgA+gt7gcQX
dzu3bhL9qJqwBG5ClXCsG6TO01eRXhrha79t9tdOyvCK4frynuCUoXGurqU2gniN
PXrYLXFtjim8MH5V8EgWBYKi4iLuR5RI+IFzvoc4llONapamY+ZmSKUWiAtqoXSC
y2b6OX365TBJ+IttDoOyyQKJi+CGgFzVgGW7MiPsjTvD6KZDcUmhYqX00aS0M2Vh
/3oyH0RoFz1U5Ep8oqcgiGvh+jDY4Bbe6v9QxDFOhSKduYwEvztjMCF1I+Fxfjcr
Aq1KZt3reTz2zBvCfH4IoLa1yYWreB03UMS2en1W2Ul/7XSmG6tFnS1LqrztzlGn
+9JidD8DFTkJTvReQaKbqZQqg4IkTC6t3l42pEbuDjOousCLlf5p01ywld7kD03b
bnoHxaiYm/sc36nM6wNKPiKnUYLIDlSmDFYnRzoJNv97NKfxxr2uMm/VUQUnlnGE
42uPokCeJz3pa4hB8xxnUcSztcQ10S0FofqROTK1836A1hMYX+tiHpzgLEGROAif
ww28tpxyxRrIWrWZg8Vx7bm9Xwq6aktUqwV80szKrYhqVNxQUK3X8436PGE9iml7
zvMlie7qhkVt951bkyTqVnq24bqiWrJWwt4ayJLQS0pzKs3nMl8xl5O/YZZqZg/d
mZSBCTx17a0B1dhR5BpKcQ==
`protect END_PROTECTED
