`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCOUvfmTnN1PgQhAmfvi8dyPnY71m53UajxDwdOICScV
23dXT3uetZ0pUIG+RXq82A4hUEUOXKvx7JUd1lk5PyynLY+K65gY6fhqwL4unI4g
KQkzWiSDnhOeX7kjGBfM4YTzFa6Bj57oT3Rvb4DFXKH+e0JjNWz/O0Zrd0QND3XR
ktlVAuHNhTWv/cYSvLIGPxcROxusstZFAcgypf8lruCo4EcVmnDzkRDM4lJ/pGO3
EQjEpeZepdOdp0VozADj3Rcziidgjm/5KUig7iq6M+rzKUKNVk5QyK17jkbEUjn6
T/mvew0mqgwH+tytzcTF9ACVl3GzBBUUmnFHV4mQniA3Pe6IKg70CFcCfyWXWaJs
2qDRP5fgFIAqvEDUwamCStJmX1n7zpGpI/eMwfYzRgdEPvemg7v858G4Vm8n8YCS
8XFfLixVYJB6u8znMLTGuKv1uyYeO8SgoM8qL5Y4JAYQsZx6he1YKx9ssqssjWH5
ZUDBoIbCVPkbdqBpczpCcZ4+RWTZ0Lrm+K/sBJgH6d4bP+rzGxI0Bxgsbg/utdJX
`protect END_PROTECTED
