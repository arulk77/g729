`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu433gKUjOaWlpgpQ7WP6Jsz+i7PGN5nskD4LxD5v+jLDq
XyRXFlAHgi1rsbMEaX8tSjVZioIw0kNwxPZ/a7yNl3t+a9NU9XpqfFh9frH/c7Ew
T/2XncNNQ1cQLmFBWHK/gJ2dJLRPFcc7SAsKpBl31hHrMgnbIzCRFwHub75ULnFT
iBrA4RFfh7NeTQZJn9plnamQrziAu7TuOLxVINclGUU=
`protect END_PROTECTED
