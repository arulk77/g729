`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40zRLzeUXAZyC/6RQ/FcsfgC078C1W8Vy91XHQeqqtPy
74SAOBYKgY1HvnHTs18DINFMsUAPs/PvcQfvUjvdQX6NTey6vPE3myK3CFKdRJ2F
p4IkdGaP2X4TgsgypYUi7eVhY+ZCGVCLZAUF6TkGwgDw+q1qxp9tARWq3xJIzrfq
tuR+N7PoovoYqZIi+/AF75Ev1FBVUR6JZcOnYJECQs7+Milk6oQjDhnVUwpO4LcW
VrE0ZqPDJ1nQ6f0av6PHgaKOaTwHhUN1MeR5WNdrMydzQ18MVPOjKhgiasXpiBXb
P0+zG+hPLeCLecnu2KiY+A==
`protect END_PROTECTED
