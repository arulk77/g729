`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3mFUa0YdhA+Sio6uroqSflh/1tVgQJpe5VRTot9H2LUbMBykuZroC8B+IRaGEFAc
a7osGC2ZJZIpaPp6m0HQXMnmaPgDNSLN3qq9NWcGAEr55if9h8987c0ZgvqRod3W
7iVHLE1m+JxQybr+Nww+1xaFhQPuub0DuClgCiefpOlzu353912MgV13cDntjlMS
hpw4XM5dTVi+pyO/5CPtWeMqxBLTx1VCRjK0hJ7a9McBS8hWX6yoOEPr9xkTBhpN
Cw8CZfMlyTKDrDYXlpxlXoQi39dcrOGly5uT6J1z8nKDGl+rb51OE4AwGGlZ3DPX
6NPNPW5m9wyn1C6y9CXOiUfoHMegd/dBvWsF76x/WlfRNrMnQ8bJVr+mdjE9FJDL
tX+D/pVxzm+yk9JvYeDkRmb7Jdkd3N0MPYUxzgaoq0pbzlMaoSXSJ5Pk+R0sSyCr
HO+VW4Dt99iDwP8VnYPNGxKb4OvyL1LlJnKbCn+mV4s+GXybBpPf10+49jRwSZzI
sNxRIzGgAkAqSppkICeNW7nVAaRhS/UiAlcJGa2vdQ84gLQS4oRbrYLflL4kThBr
Tn4sAemvCBA1okhCvFnJ+7bFqa7CI8xWKHAfHiIzU9Nv/e9lw1rz3bnXRDJM9rb2
4itd2z0ehreQPfo0TFTYmnKPZAQDM42mdLLzxAUo7TMXonnpX+v3PVeV68kSdssC
arQTHYboFAOEqc1aVVVvVg==
`protect END_PROTECTED
