`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
CXDo269tkFVLssJhCUcbkYG8O0BsCJolj04ZKMPaLD0S+edh3WwpLcyTX+w9CWqD
UQvnzKDJl1Lv2k7Ix93sDjka07Y9V926T76pQ+9je6oM3+gwq6c0EXmiSgwMQmQN
F/bD6v3+eDpGt5iUMl8JjIo3d6NXN7UmhdPPMkGg2kgwEXyDtcIWSqQNpfvHLgHU
`protect END_PROTECTED
