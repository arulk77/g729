`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL45ClRdBVBBY0sr9A87boACkTLFWvvLLEhpux1C8J9a
B7No+fYN0vr86nogSfoZRX85wUP6nmCY5jCWdObpc5qUZT7Wkr4Yqx3PvMx13xKi
QnGG42C3KAdyWy9epI2JvgNiKzSSB75Vy9sobnUm7pcWPDo4brTYzgO+QPJCBktQ
6HPvIwD3HknTjZwFtfikcOniieH503xW9VspYa4m7cCCRIjRaMiww0e4Z6IPuX+u
h7/81NXlLdiaDASDTfefQeBL0vM9rqBCAII/q6DiH8tmpu3jHCClXRMu0kC/qPvY
G5SwqLceRPEOxfKECFtvn1dCkM0rwHpFSQhSEVt1/E9DmU12oMt4dbrSqjTMQORB
Zc+AXK1ZjL04rYlhoDmX3NdGwORZ57sJsnqMhznZAzJQ08+BaoidYrXGO4KuIRgS
Xt6Zhc1zC2MVG1Hm+a3yf2uoQW2h6e/ocf5Y4bTYucFaVlyKhmX7cW/Ah5TLtIFf
7yyuYgPLW7dO/zgkt7aHPf4zovvPpRyh+XrztaqUE+zlO/aWE2UW5Zje7Vsht/oI
SCddKvmkig7sYkCvZE6Xri2IZs1Qdr50vhbXGAkk+/g=
`protect END_PROTECTED
