`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBqwiFELuCkfoRWUl48w1BApgtr49DAPsxranV8Aj4mD
oR9Kgd4PC6KcQYFVwtxON8bEjNw/x5NQKEPVxsNL9bPizqnHXl1XqRPfBjXcku3I
lBUwbbWPMpf3OBrLy1fGt2sTDDpYWHJXdQY6WTdBkr1fZjJHJwRz/un7NF60v2Yg
1RbhLn+m54JKss2HfhNJjbr14rnxwNGqFSsrbCZCnEd1pfoVLnaaiCK4D7ucjZAw
CM/6qcTqlrm1+Y6ZolZcurZzyxX8m1Sdvt5kWJeDXxSzoT7qe3bIL8s4Na3SG7Gs
O51Jxq/C+wPm5mzWNXKDMARVGAxgA1BgIHPDU9csfYNiUlPdHHSF+eIZVaxesGA1
ObVF2/kykzcBmmqaF6rVOS7dyM6uh4Xig8ZecxTxGtEtgwW5mevjMAKgTq+D+/45
`protect END_PROTECTED
