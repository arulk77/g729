`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveO7P3YmN6ncCgwtDQPOP/fd71V9T74Kz3LSKgjvzBYYp
K1qFZkdaCVJbKpifWsu7YeHT9zj8bd2v35i5RlgVwo3aBkjszyJS1gFe5iQDqwEA
RHPSFhe+ZSfB18uvFRisQOeU7G//pjIGiod1DXfQ3EscZ+ut8TmW9Vl1lFWNsJHv
XT+EdGxEA/F04/Tj5HmWpISq9dXtZ3+u5gYDBEikc73Ts8RWo6+wsJ5DFZcCaMRT
mn5AqUjzvsRpw+xqT1oCatvZdtB7nJr5NCMndRiO4MZQay7XjpAJdXsmDeCZM6rd
aUjXSmiO7c+ykuz/6DHKUQ==
`protect END_PROTECTED
