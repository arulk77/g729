`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
G2lyJLtFYpJoGV+0/I2UmoeN/VLlVPk5RGwt8R0tP55L8pHKKqL5moiM0p1Z3KxD
y8DBTP/L6rjWNNpWyVNzYwYdvc7ETVT16vfTdJo4pR+pG140L60Vj7QrAiZCKmfh
4APhy+LVgYKbNNKvZXB6A3Di9mcBgovYwqJPEODElsUf6q5AMl3zmNiCCz8Qr9MX
`protect END_PROTECTED
