`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
LRVAfdoFKx6URBusEDw9ZR9mi8bqj5Pv9GnLBaz1NsjbutypQ87TKaCADqFmRpCE
/ChmJpEmSGUTRnVaQ7CzZhJHzrm34BydEoqjUp/s3yDOzPJs4q+LbKfijpz43Usg
UHaCjJRijl/Oq3o2WZMQAm52bzTVcxLNrJsYhe12otzVjjy6WVXm8U3QabOzFjGh
BGfJxwYO7x788V+nOeOR8D0bj6+VtgSSD267KC/2JYDSCuyf2LUVLn4Xu+0m7A/w
69Jg/wZWcCC8GQKrj1OTEm7QzhbRo27POru4rv+aOMkDKzXDp+PXik8aecxe4JxM
9t6EfAhwaGynokPEtow/Q9RdTeaJI4XlsDmPfsdlJ33qnOuw5l3Yvx+6B2jyDRLB
DiFlNpa7uWkv63Drmch4w8wpO8xI8IBBTOTLzwCWFWLT/5LrEdEZ+O6mo7lxcpsY
nL1RQlxxo6MRq6DLdNROJ2kOGpxNhsNc/AOxT+ql8nJBVoPf81ZUJnhTG90q+mNK
eb56HQ08tolUBDNUGC/XznnSEde5H83wtLdLDyt8fhabHdIljAWXOBN8d+7uR+2C
ArDNuV5ymKsghWjzMV1B1aPJVUPeEf//s9PsZXd1KVmbfm2u7fuOq2M5n2RFHDFG
TKNe02oH3UM8RkSYk9Xn6EPKKdMpOct1jIrdRuv93Eotc61ONqIrN3bnH3S7qvMF
DiJUSLaR2d6zCHymzsU3u+CoZz5q1p+9oKQbHvPOGg9ZWHOqFi6/4E/Se81kUktv
Ys4vnlDi0u56J5VONd1gdQ2hICIbytxePwVm1661Po3anhRg/s7WDl/74Z7IbNzf
wHFR9JuuOMLGawygItV+L6xkRceiUhN27mCY7CUJyqSEDS0ptvL5FrS1DUbvXaxu
0IYIqw8VrAncbGk7xa3g8WZn4TZyg7h3/i4HL5qqRNDjTZmhZTNbAstUhfRg5YwT
u8G33bUrqi8Je+12aqqGRKkKvXfW9bY/PMKKqCzfgGM/t9MMQt//K1eOx5Fl6kBL
sa012HCGeqowDndkVorlVpHiFi1K7tiMCukI7nBG3pfu8uqWw4UG2sYD6R03E1FG
l53equPnfTnr7ElCMI8dtUAslHcn412llmMANqL0QNmq8c76Juw2DkliFURowmKz
4s8albQySsLaoefJkOBevvAuHYVGDWKSeL1U6rCj0MHy27Hiv+z3TvyTXLDcAJyf
`protect END_PROTECTED
