`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePGicrKUuR9ueMTyteEGJ1LiQPNdC3ocoIf9EcDPKMs2
FwA0VdmN3daPRIGwYq9wX3eKyK/1Mrd0sqUXMEY1H6IvzjhZqN3S1MIFSN3+s9Fz
Vlo+8Pv+GoDAcka0l3zLEoro+XY+GplfzxAp2WomtzacY+jhHfqRbtxbR1XmTAYH
L5djDZoEVLR+Vc/aBDNxi7duhNTSEKWUjIUq4Idvc+eydXlg4YQwIZvA7F0revRr
6C0uSWGM5IQ1hnWGsGXSXg==
`protect END_PROTECTED
