`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP/kN7uuZa+FEnhyTmEUWowTYl6XtZueC4cbFzqmg1jW
kcu94J2eyq1f4tQFmmG1EGWl5RCNzT/IhYjbTDF6FnjsoIC2RcNt7IHktH/Y3prT
sVCsZ2+npewgIaEqSLEmZaoTIJuLgJ8cj2skdJ8Umo1lcEPYa9jhG2U3C/THOQBd
ptKUjYSGlK7kpJuX3sP2PyUz8L0tg8F5E8dX2QE973j6F2l/iBr9mlCiEciYBFYD
aQoDsu0VDhEyr6+CTjRxTwibzUmP8VS1KVqtvKwD2SYYai74vkyXVVdWlYh0qLIK
OevL/8GJFWTUt4xywuC7UAcHWb/CbFoxYliRtSoIAnjj3Ug5CqmvM21xOL1Cqzfw
cRNCd2GxAFXqd5qY68CwpHhOD+kqZECvk0crla7TlYoYwMCPGXUZ2ula7H9+QEBa
AsvJIKuQbt2mqyXHuh0E4/ZMFOjmTLLOksqu1FTifu2+/O5JBvzQGEgwPcxSxvKj
cLqTzmk1Ejha0h+MGw9wcf+zN0/m3qmNEj573s24/eSEr4yGXWSxnfOjurv66JJr
`protect END_PROTECTED
