`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zYQ9Kjn4alIKRi0PNo5ljw69U7gpANLoODtTJMfyzim
dy4r8qNWbvHQepfeDHnBfawRejmULQrgJXsZVA+YZlLe9YhpR/XxqS8QtGa2L71m
wF22NYPheGHDbARJzK0er6FDMiFOJy1jyO8952zq0ZQAi1m6HMj84btek5Das2WR
sFNK0/fw2Lc/z9RcR1ubaf2kuXLeJbqlq/qVBxu2gjw=
`protect END_PROTECTED
