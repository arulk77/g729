`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJZGZ0M4yzD7vxvEhN9JFnR1kguQUPGsMerAdSP/2xmp
q2CMrxYNiBQOTqcFe3frjjN35ZYu3WlJ3SFiK6YIrMP4cKKmvBoDz2xO2OCuJqNN
aiGXeYJcOD3Lkyno/NGQ6XmuYhM0bblRUBfjKNZg48qT8fkQOxxBj4rEhMFw5LWV
XzCElhOctJmZp+HpKUpDLhFchcLpldpqKHsAdX2EqEJ9Ui3IgKRwYzgtTLZ4ZJxc
`protect END_PROTECTED
