`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAzE+aeMLe0WFwjqSZbv386dvvrND2bgqfOxfQ7ZLhr8
u97uBfdGUGbq7sxxK+MgySY8vMdUyn4ilJgajIyeQmx3eOOIC1YncMXPLI5bEgbw
mRk1FmVNSrdms9X4FGh+MgMwaS/AYWrv04rkfOpMnUdaCjj634MhUrGO/ELsAhjO
+ettb48GVKBtNtBriI7CI98vWYIjpxP1PDNKeG27Yyk/mXz4yx36tFfwz+EXR5dz
YUxwMT/aaB8OUW8dMhf6e0tiyqEMUsXG4tI2cprehiHQbQY0yoiwnqmfzhKb78Co
0LO6dE5YWJTjEgq5pOAuKQ==
`protect END_PROTECTED
