`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
HkfpqTCjR3ahsiK64E6opa2h270vPu0KnRZozUxVjIIk6QCE9s6G3UgqqUIBMraj
TEZyhOcvx4pRMKyFviXHX4ucD0PIErYwIDEZPJELAL3EyLqUkiDLOHrD1fbcmZDc
ed/JaJS408M64W+nEvtMNIhdTcnC1iEhWnDTCsot0O8=
`protect END_PROTECTED
