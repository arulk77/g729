`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJMFXIe8uEzOXfAc6L6qHNtKZA+vsCX2Lrv4ECddLKAD
CGt3V1rwndsJXJwYGtUi+AFX0PgEi+Bs7F4lx+yUh+u0EmtyioevjiwpniD61X+D
BYS5bhV6VeS3CiKnTcXrzfgKBsghHYB8RbbygAcrM3Kcb/cgBazAXh8+sZ+P00pF
FAHITlV3YK5urDFXS+12G9ZmDJv+eEAkuqaweah8zKrTILZxweVNhImLsK9fiw5u
`protect END_PROTECTED
