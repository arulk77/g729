`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
7RfCgSSEYuAmMsOKUiuNAWmx8iVTz5mCGy2rAwqMT8plDdG4Pqm/puSMqx4d2ij/
9The7nMqp5WrQYljRh8XCmyUzWE1DJ5tDBT4cCFEthVOOHN46qmJ4qEX9I51go4w
U/G2V7dkK2c/bDfgOzPZjXY6hg426fl9usAMFLT4SxlSxoD7dnpKFF0X6HPlvD+l
iG3eJNOqJDX6od102GhDlwJfK0Ljdx67s4TT5x/iQmAJZ9Ynob2FPCZT9XebgwXn
u0TjiZaO/hij30VqohvNBvfnnIgQuU/B01Jc7jU4YeY=
`protect END_PROTECTED
