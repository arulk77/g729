`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAQb/up9fznfdhYCfQH2AlFG7w2IuIU2IrbNqMUcZlPQ
n0ti8UarA3QF2VLz0xX6+InyQOSK5r4JTXMI6MwD8A43iLYPIIA6Ed77KJbVgZ3Z
DqHc+R6gUKyDNzoIUW1MZkwTr5z1CXUHV2qTLj7PidRm6878v5+lkpstX1nsqcby
1zJ7fj8SEsA0aIq3dxw3rTo/F5ks+TFMVm5kqyY8VKcR85az88fAtt/xkEUgc2y+
P149b5qopOTvFNnpBoTuYy1ZEjwAmuwZP04yTHeOjUPscqaMUB1kaQSaabEaDV/H
dddslf6Um8S8ZwFx9KqPZYQon+lVUSvtmwPKQJ05CzX3hMVXEscrynqJVzwmttfL
hlP3u3+n8gjHWZ8Do9I5YgFcBLl3N7WiXQ953JMTE3I+VpAsqAXsoSwTdr0+5exB
QUvGD//RkJQts6zNDxYEWgUlLlGlgxHBj3IYNxwNWQaqOB77pKWJg9EqUypq8ofh
`protect END_PROTECTED
