`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Y7qB1uVeRlsqTjIbhSm8PzmioY9IB/6SphIAPETXuNO6tbBLJaPcAJFzR3GKti2a
Fclrjh3F25OzXo7qnU7cqDThsntg8MHZMBsB8jEhnF8rNYDPArSEjV3unl6wocer
auX0Qw6JrzKgXzG7ou5W39pMhsQn6PKEotKa8MCf9Pit3xiqrd/zV+or8apLgBa+
62hCJRY9Z+2ogTr8Dp60I0K5acjId0P5Uw/rIXx3qUWVdSUfXtNY64safHpHTF7s
a9A8+rMqylAbo6pWEA6YBzisjuxpPKpEe7YiRIgPN/A=
`protect END_PROTECTED
