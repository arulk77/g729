`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJSAX+6dIUc3Vup9tqfQww3YUEPnlIlST/1nT63lEy2t
dIfDS10bZO8p0a3idoZ6/mphtur7DovMwLdLslNVMlDaqOTCyrJTURmoeC+RmRSw
RjWAkZ/ZLVru1GvcJBlOP08suR0kaeWx8J4RowblMRlNO6oX/OJ1JPtrhd38RvaO
Jf4Iy6ey1Wj+YdKkofBXep0ZJ1M9sgTGGvZ6ESay6G8fM3LcgUN8OnNNRfOPvCjW
SX8C7pJS/LNNDMXUz7cmrq4HabRGsR9FR3zF3F9TRtvVPiDp0BPXk04LyJUjPgha
5THdlJK+39PCKM6Hp4JZ8Hs76EEDpn96WIeQ0yx5inw4IqNSBHML6bDvrbeotWoC
4ia+CLoS4pHqeMNXRRr4BlCN5As/97U3w8wZNZH7Nm3kgXuRVFdhwh4UCU4UCNNH
BJpusqbMG+ii72NjiHFUnKtDNuQJQNfBBQzJBFPl0Fc6j3zzguRRwDMzXL9h7eHG
NJsZwzeknHGwHVZ2ZRyvI7ruRX+DW+cPztmET0SGATt9f4fkZ1XEqg/39ftwI77+
`protect END_PROTECTED
