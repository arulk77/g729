`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42CRYY1k3h1DI5Zx5kk9oerC0hhL/GNSz8Qc9tzCP6R4
xlrMxVrzc9RXaXGFZVZ/jZ5z7iys+2g29jOv/Qn6fpZFf+X8Lj3SnMud3lfIxb2L
lEFBBs3Fuqrnw8hzlKSXr2igqE5ZhC0HzIdxTvvUorbnqTmh9472hgjE7X28ObhN
scH6gES46x1GF0vS2YA+GqvdGjcZnXMI9iV1eM67vbnoSfEi9DZChUpvZTOjqI3U
wF/7x0xfL2Jmtifw2/MPf5ViNFyAW3e7ZbcNHydNYgw=
`protect END_PROTECTED
