`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGAsYINQIsHkBfp/JCHvgeBE+mwB9d0BlDEMUcAM0fGy
9DCzvjDQK17mSNTFVhUJAX8Jhejohstusk+HEgv+O395NonlLMr4Zjb1AGRuIe5h
v/A++lbIhScMfWD8jmtKYeSSHIsTyU95Ilqpk1VM8zEotwcgx28P2mnMzDbpd08K
Z/Ghz35VR8KtffRr8Vjqj8cxSmdReRi5mQONFvu2vsFq8T5sDln52NgMON/g5eP4
`protect END_PROTECTED
