`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aZXLjlLAjubvdr/D86EVWUc3wo7I+jsb8JO7YVsol2Jb
MlSSnuK8qibtH+i3+CWTXfkA9uQoIu5vVfmjnuLKhXu7ng11HVqrMyD+0lWQDdCL
hFyb6sEk6NoVVab+yA799vsCYJnN8dSdZ9mL5ShXuTXju+aX0YNjmnc44bE1kdPn
b7z0GmU8u8xfQqbesJdlhytQa28olLkjIovNqc0tfdfTpRxyQvg9+AF2rK1uvRaD
/mgc9QWZN1e8Cb6ShwLXHNm/ojteqwcBK1Xu/7zimBNfnAMICzF9Hgcr9ZDBQ5Dj
zitSOtfi59Pq2Xqo8SMAyQge68nSCaSD42QeUtLcSsm+w/SCzjxadM6gyP8TUwYw
EVSwvm98F2AfmCTx635Du3NkEc1xCZLG0v0mDK+kNS4Sz17pg++tfjG1nZJVNY9M
bCkkIpxg9MMU3LxWPoFtWSpTl6tyWUtGIYcaKpY4boR9Ha5lrmx2QgmzTRv5Hgix
9640BzwnTgaVsZhpoBP99En3oF+I+RcOmDfOjU1HA8pA6/MhlcxTzaov3fppnYXt
fORAGMX/XAF3U68AOkV8Yag3FTqXEl2w8Db5tAN/W7LRiGVVBw8UdRbEe2yvydxB
8Ci8MOGb5zbLII60Rlrnb4OkwQDVvdy+/sTQxM7zJ7E2RF6Q4XtBh3NRuLKCVk95
TFuLQVv0ZYOAqou2f/lwrB8OH/Q9hiytGRRiOWiYPOqxc3X2u+Ye9dhyQLL/Lgzg
XCJKHTMV9DRHFnnTZ0TB7/6j6E2efVG2QYIzZLEbAGHpdznbEbGnpez5aF1x40sF
cjCXp3AHTovI1WurzaGg+Cdtgn+8uGzhgQWN1gu0RdmD61kVYF+wQhtEJcdgveoT
AXAi9skYty9Nrr0U50s3WJWLOeLykO9+8IeWbU0r1kBGYTUQ8EVo5XWIYT/qY+3L
OtE++F7FRQhYAvKHqy5HGS2GudZKvT25VrU1fjnFMPpm5ZeudLLGoI7GaZjkX0aR
mID/3lgDMF9dthtNTaJClZMEP1GYnjGyCwOhsFJWJXe/2UaekNMTx2ceFa7x9Ja4
DifNsYo0tTy3NW/kDZ7/RDaDFbrn1ueuMGyEYasew8DyIyDwP2I13jz4QYwKxvS8
UJNWHW221QRbqi/9EtAVu9dZ6wcj8DcViSMLs9L8mhI=
`protect END_PROTECTED
