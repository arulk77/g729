`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47889/2GpiGhIv+ELZFyO0SMX3WA7fpsJEZwOdJCuypo
v78FTkQqOo1xgCsQAFJPyfvhh7mJBmTtB2mEqYbxT08f2rlL8eJ2jz2zH641/cdV
stQielXBJwWtdXSid8sCs+LmXuN4jqg4VoUNn9VTirn3Xwfjk9aGnuk03yUEcnou
x2G5YeWb5IZZ5ZokKFGgIeJTYy81NZE3syz6prPht5w=
`protect END_PROTECTED
