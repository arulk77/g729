`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN0YZ5/PjYL48eoIjISzfciZ/Ct3YnH/P1wqjclFCwQGv
dQyXXm5+86R6fag+fhsRfEwd9Y4on/80PAi1IsjvMTvJrczPxUedtKdcFfOb/IMj
gtRUuInUMijvOHMiKeDgSLH6/bWFvq+U4aPm8TaVMgzFT5xQtxtYdA/AlCSvQGnU
m9pH3PgkjK//0MRTb4sAa1tNsiSp5IDWHHzB7n7Ctmd9HGqIPbV3lpCB/Ca9qwIw
jXPxhxt05M76LKJIrWBuAp721DTJAI7d6cPuSf7jSUMZygSlN9bS0j2ddlwbQenF
iY5oIeCti92SPsD3JBjt9fObsDljU3RvQdNC5CKSwt/G2iK4Rh8AkOoQ+bf3dwC9
1ZoXZLfNcULzsICOoo2GpUlcRD4uTShCZBtLR4FFe8R6XV2AxUvO20Bk5M4iZjpu
zCaEE0rT9j8Yf7thWTdUFzBQolTDKfXxtOezBbKQI5gSrH5MLaGIDKICxZqw9+Ge
+kHGWNP5EqfQZuy9wHwB2mJwSb90YKBP579X2UeUq7Qo0zYHlBRi2vEZMpjJqxoO
5hYN5y3u/a4bKj4r14F4vV2EtcsejOoOlc3kUZngbTa/n2yvhAddgze9nEPC9VOy
S43eoRInJE+Pi4qx3oukVnSPzUx/a8/rfG3JfPgjYeBwm5u9oUitYtKflQZsmRv8
1g6ABIrq+8kdZqau30eWytvyLWTM8qpYZ0wJGfn9X79hfJgEV2N2oLlrmFVitun0
y3DNR4gQRiG8Bnsk8BwB0mG/d0Cu5vFn1wx4xCgl+W01A5kmKvL9syTmWiZibO2L
Uyd3MyK6x6H0GNgu6GPMdUfKx6tD2ynnY0Z5v8W8z6UonYhmi3Z7aiSXm09jdbMk
33ImMi2NeJ+0yg/aPyA6boJdl3dhW6qLJL6JtlEF4TV7DQZQgEhElwyl8bvy8xgG
0B8U6Hf1deeaoYpwn55g8TmXVy4FKkzsdFNzbZoeu5MPtYCdmuuMqkkYPCw1hFqU
WrSKDMywgLX7YF+VWf7x8v4hRkIUXyAp22N5t9YL27/t9LNFfpqZulc4SXb2eUE7
4vX7cVlMjeBJo/bP/DVA1K6Zlv3ehHszsLPi8H1rQqkWfCEmDvUJw6f+pGZcJZQk
0TYLSlky7vLvD7sKwknts0vK+ypeq4R2xrNGsNgFrCazYO6D+76dYLmgHmHk8uSI
Rt4ifmIp5jyG7KdM46czJj1ShjMOwBTFvxJI4Po2vaNe497xGmxxVLWTDQSmPpdX
srgh1aZBFHqLkZWKmE4TyOKDxi/q0EblXqcWGq7Q4e8KaUs5IEeGL2N1Tz4U/dZo
E9j64K8oPlfEqIrpy9rzyIkFQBSA4G5+jvMVVWXlAPZn4Wv0yi2FFWnzumdz6rf5
iSE4X5HxGPhZkhDBZZUqenGg3CMVOu5EEl5nsEk0zVvZJ/1oQMp1R/NGVHc63yYr
TT9JZruZ6YDtWl9nayKJ0Is3649pIs/rQAsLDysNmOXajNaU1XolrKmMlU5WmVn/
tS9H6CJwXug3b1t2bVXAQ7Lo1QL0QQx4RS1xq3avds1Dg4FxScNw8geVUniMvXx2
U252dtyXxtmp/L27rgaQtZAIWpsV2ojh+l3Rme+i2qjJCLkNfJL8GX71oyJaSpWT
qanETf/hJWnuH7X2t5DqtfxsrGLXh6qq7AT5f4ewVtx9/uXQpTri3J4WnRfiOtdI
30OzahaHFa4KY4mXne8E2KBrEpApfEdKcELLJE68WDVlp3iPMp7EJSIyxSXu5AdM
1Q5y4GMy2GScSn/cPmIc6AciK0tOFMH4ujvXgvgmEt4/VIeFTAkv9lbUkwAyzuDo
jq2sEU5ZRnGEe9X88pYjw6m6d4vXiKXMLfEsA0miTeHhqIPpjlonYyjQwvbxSbyG
WO8UrShHm/sk2LKUuXWNja1+I4EapeLs71o5zAVDlBlYcjqoptzteQSdMiTKBhNj
tg0eKAbLB142nhtd9u7c0h/2wcGzMiucCzGKIXwuZcPuTcRuRrvcKNq72/lcZOaA
iHVAalnc24uGAq0jIt/A/Jt64tIn4LCuYxUwNKmZ634B2VfQUu4M9LdBqB8rpUj7
aDUiL8w5OoqiaXceYp5/Rs04EJQW/aI1K0JEaZTt7c6v53vySvft/7u6Ws1TDt5N
5oeUJKO8l7K8R/sGmOYm4p6FQ7iKpPnHHQsFnrNGkuzmdOzpUnx/MOw6g98/j/Bn
QFO//AOXbAWdFxzhC1mn33SFzpjLbbkdBAcjxevqiI88cntk02a92UaGmNsyzENW
f+bnI1uYcOvYcPz/nvqr/u4jq/NWYKxDb1nZQ/Hjg7pnjtcxx+pbMBfnQfpgg1Vw
vvYHjbiTBVSy7Wh2ltWR8vt48LITiBFzDtnZAYpv1ZI1ccbJMP5vb+Aw1IYRoRbu
T82rEBWamMS7eWv06Qw2Samsllbpe+dqHtQDG+ZMnKmfCOjzSFjBnfcTj+DfTdLN
EgzWQYr9tflTCnTfG0IT1u87fQ3qls4MdEDYNG4eqo+cfcqZyHCOyvmX51J8Rz35
uZlwbZP8dmyMZOwCfusDaJ0ugi5IIhsppO5Rv9BM0rYUAV/QP/4c1K20iEGLYnTr
8nke6c3Vm8d0oV3teTRqC3XUO6cmpPCGWqXfsFKlhhjq9lYBlXOvHGMFdsRF8QZH
h9smc39F2BB6brIXsqSuTZNZ82GmVoi0y0K1J87O/A0=
`protect END_PROTECTED
