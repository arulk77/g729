`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM+gSCzjgR4NH26GxIGGovH0/xoPmDg0PRDNAbCEAfIP
GJhE+shyNThJA0AP0xSdIj2b9r7uaOH1K9N8Uwk480JD1SS9DhKig33uVtP1KlNv
1P+F8qEt08BDViSpB/raii+Yr6SONi9rVELqGgWVlcF4SpritIiN/DbFQrV/Z5Gb
uLFpWKT5jhRRp2D8TOZZ6fnRPeJBJmmaD1lsJ37huKxPgvI34diu3kGDjUwsTGaF
5jiiXJN0D8ARDarMNR26szWo9l04ro+fY1mGdh2bKiQyz04bCX6I/k3/EPOaIgxz
GfrGuTUqUQ6YymQP9RYGkBUA/RWLsAaYYW7B+REeT1uuYZsZJiGjBHKVydVJzWiF
C67wLcul4g0JkwmYmjICEQbOnQ6hfkLPb1XDa9s3pNrlyruJM4TIQc/CxN48MyOz
ibLz/mWQ3ONEtHmnxAeo1BQrqVUKTbBhujSpkoH8l/8KWJ+Xp5N33G8TCOpgmD+C
`protect END_PROTECTED
