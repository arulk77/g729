`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBhy4t8joRwD5Af7w9oSIPF5QJ0t+rCTNK7tFk8JmiU+
AqLESZKB3h4DT11ArHV0vZb3GFaM+lIi9ZtCwAMEgIPx2eBCcHtPj77+FF5ZN9vK
3UO7A9mwCl15dArCHcy4xMQRry7qHmzb4GLzWKsmvSPq3PQA6xu5hkWgvebhtkjn
o+3zphmA4WVl5Y5gNaWxLUHy4Pf7tw0rC0KzDWqn4xgxSOxe6vYVlu1IwfYxJBMr
mXrKhNtVtFLxq95N+P/LXZWRcUmA0EQu/BaDyqsVprYTYjkiKDA60vzlGmu5scBT
1RzQ7EoaY7/xdsg+Fz+RchCfIDZZilc3ZDZRLPoWUDvtphggfKG2lfSXFapzTvwP
TXl4trRoFICiFFdz2wyElCxaoJ9ubInbixQIHvh5L/GWmFHknm+sdEXpeTE754hl
UBMlVzfaGG15wGcepqs/qJ5BQMCIFPCrUcUNPJxrguOwGeG0hN2QTWfzwcN5aG1B
`protect END_PROTECTED
