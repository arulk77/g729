`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP4BLzoT/pGRTee4F54LRnguiZW61y7lDzMXviPUTDuc
UUEYGIF+TllvyDhbQ1oOpPWLBzUrg9vn27eHz/v0oDh0nqbGHlH+XjfdThI7Il1F
9Fuu0eKIq8nQU7wUF3EVwOkh+qgMO9w/8ESpQkTKay1H59tk1ENBYOO8H7U7JjlG
t07Z6ZPS3uk8gIEUJA5J4Z5Xz4wkOtTNu0FkqKWyoLvj5VWDkAJB93kcA5KuMnOx
GTzYVzecUAuuwMhE1d++vQR7zUy4GiI5TwHpvWDEFTUheYcNAxvweD7DLWchvcpF
Zuvp178F5I6D6+cXXZt8UuW924C3o7kJPOmMDSI7eD3P4Q7fnN2Z8BFaq+C2BI3b
uWcsZYAIkmWm6IeTx+BYf8biiaOT7iBDTF2ORsk1EHiLfKBkkvGEaKM5D5+/+U7T
aemP2n9VRzb/tACs2UQ9ORBZUQOeKy3O3fay+BK88rBoqzPkttCZ0eIjQ5tWy21q
`protect END_PROTECTED
