`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIRO9KZmQibfkbeppo29UGJF4zPa0Kd+exgNwlRSVzHX
ebTzYtIpMoX9lYGyTX941YLHIcCQ0Usm4ML4pwrO8z2fGHRi3MIHdpPjVgmS3bcl
/tgzxKY7gDqr8Bu2hNmls1S7Yflmc82vbFl4EZsqYsed9sVPVzNdxJJWycQC0hZ0
2viyIIgQYEPrI4SewcHlbXR08YHH73u+Ayqtv0acw9CsK3eT+K8f2yUdFv+98+Ow
wCUK4nI0/qT+kScwxXEbXxWrvfuxRQSvsdPBesbPRU1T+o/LRX5C2J52Ul6NX9Ox
uf9VPfepCPL9envy00HXc8hNICHmpXYP439ztYE0st/epNPST3V29xtHKjASswPX
2e4J/St8paotxXnlX+dE3wnD7MT2OlpnSishjthWdtefpmfSVTuvX+SYWf5yK/0p
rJI4FumPEApxCRPFAfRlvOAdDpgruTZrn6gRM1VsT9ukCFPM1fLdjvmmXcS0nD++
`protect END_PROTECTED
