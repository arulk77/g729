`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBJ7BqHUR0YTKgeZHjb1P09HYMSs8agT+CoZ6AHY/mGO
krPTBh+ghyHUbFgGIWjRN2fQCq0TA96hVDKhYhJnBkyC/6IX4EgqyrDtW6QRCI5j
qBvqu5iydvyVy7w/nWMmPwAMinlzkgEoKzBaShAMPk0YVk8OA7s6GbctD6huQWQ8
`protect END_PROTECTED
