`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMHLkvyE/rFUhhbGeCrSUXNsadtjV03eaJt870gqcHFp
cw65YbeSZZyDA/p+isRhH1vZtAPArn6DNXp4VTNYzquOriVtY6b7Tn9w5M3TnnAu
GbvGq4LDdtq+D76YjxVRJYTQSR4hni+u1KiP+sb8nD+LskVkOYSsOsxxqoWcN55i
oIC05BhbvyPAOSE4zLJQzvHS+JHr7AbdBEZb6yhKFHe7awSyMtE+jcLLTazP7FYQ
U8NdK/TXlLxDpqrLrmNJ4uqvxZwPGiOylrTFNNArnQLdHrWrxNtxeakdRZ98cLe6
4dsm19d85/5TM/zc0CokRDsXSPFrZ9grjPMVZYGRgaLiYt+41jHHy0mowjRiPdnk
vXpGgi9xW0rui6l3fFh2G8SdaBzd5AWrbNN5u6Ovcbz2t54JztoEDZFsP43WMfUC
WxL5ojYQFc8C22TyQk/bH/4DTT14o4/ikJlbw+G+WQtxxjvNqA47T/TwrttZ4AGn
zCoW/2EE1RtwpGm02xcmOiGMjHLd4Ii7bwxiqZiAamFqTq38xABnShjNFopuj8UN
2jLae6proVE9W3HjZVlWI/E2DV5EjSgM1h1F5qRDM90nSoD2vWA23s4/9Rm6PuhU
4OeUitcaPLWO6nSb1ELQpaeNd3HmYXF6QrVZfsD8yh0wbybSg7H7B4pyXi1fhiGS
oODMRcHMG7C2zulOVFDcfKQwf9sGXPxpIOnD9pUkwl6CFBfU/wDrIdyP+BA8MyQP
pRtNSecYWzvx5m8AoUbiE1DqOEuXBGh5S9ylu2q2cvo/dDs4iWOxzvsqLhz9CIeG
1cw13c/3rMVJT3JfXl+Ufve87MOuF0SlyFmTpSf7cPfTbd1mgsaV7AbXCRb0zqHY
BtNixTXJN4XOwW13a41AtVUJzDJttTDksgWEODebUBvrNYsUWSskW+/kDDkSYnof
B/jMM/pSQxDgd9MkFiTWrolLTLDcByEx62h1lfY4KBIDH+d48LjTd8s4k2nciCQc
fGrYuH7QG3/jHJkicAE/b3lxJtJrA3K23fggKqWmlFrNgHssSD2lrhI01oNbLgZO
+fCxcrSYGv86RDhNAdhcNAgOqNPQGi1wyXkEwep8wH91Vo7IpcUmpGzGdbfijcap
W75F+OX19kimBnRZDD69e+pbgj/Sr7Q5/XkGm83WcyPPWJzW1dDzuHMQuUcjN/sy
1eWvpjkx/oSYB4IXd42jjIIngoXSZJ+bTUSoR7dsvN5kDNbfcVQkRgXMezbEy9RM
fC/AqsjNwVKqxsQrv21y1puObydzBsPVScoXXYFFsUSHUxzCfjeVhGkhc0uQHu47
WsaN2Pkv2PIiJVBsJNb4HDH9/xLeQow5YBAyFGS2me9B4qGxZy/sHmpbRBxzd0jb
6zDqbDzLlbOoIuX/8D2Nqew9JmhdGy0aieSs0JI2c3W/lJhH7N1ZZ50DdSRJqf9d
+G3dhWS2uThi+pPyl/X+aUHA6CKCzpGW86LzstqBKMFiEgU7dCOPD9JOPYm/9ih2
SqazehB7q6MrZQJBZHT2wAj0oMemn+AlxLl7E58boMPOv9z1MLXGqkIyeIZBF5mF
yPpxH0ZSdRPrXI7s+XqnEk7ug5aaTQ1T1XmSfjPpxDpPmfD3KgKZlKFSTCq54kXX
F959LPD8E9kFVS56AtDVBBZnSu68hfFU2euD9VJdmSbVyOBu0U5iKXj6m/P5vI1I
nDD7/ueZ5o5ReN3o6l7p1AzqtlDNa9pt98Py7lDNnVMsuCwnshZwI8WuOnyg5cJZ
sMwaYErZjq9Za+SDzu16vgQWKj2anZyhH1I0IHH1dRbhD+eNy2LRF/SQGZR3Zbk2
gva+BPilVMFyqluZLhRT5NkFaWx/RooQtHGuyXo7267vvQaPN4YhFJagkahFzlxA
QxBLtsSnBBArTNiaVcX5d61Ot4jGCpNFyTCefsxh3sMz6gS9qeZl+j4gk02GfYM7
Dg3//CmahXgL4vI3o2zIteOoltXTJ33GUVd5NxyVFzSI53CH2rhLcV86O5j/CM88
p4MqsgfzIIl31/XR61i9ezsvxbCXJMkBBhQ5L921PGBcKvCAcUtNAzeLGI9t3YzF
0tDfKrsaM3JHw/EnL9fjbmjQnLXO/uM2qh+3inCJqp7vB5Zk3xVDGhbVjW8JCVLe
mn0rFed9/80X1nb+R5sk+ZsiYd8LdqZhwdzpWIaXotimLIP/OTDWHz4pHEv0Q6HP
gO8A/R1VqH9mBz0Yfzbt9G/BDsHCYU/FufyRka++sr3ptsx0RxpfexzuVw/qZJ0J
Fw1JE8rO/WNcwzqdLc1vtWcfvwwwvFyxnVLYf0UFFm87brs2yKHSSYvSaftPA022
cThFbIESkUZ+/ajNM3v96Z/vWXIrsOcCU4D7/hJmgW0G8CYH1mmQOjTjLRN7QWZ+
oPQalUihrULS+W7TxOT4KGFpjhFELIPBuptSlLAlgB2Vr03TdCbfEj6Hlnk2fP66
1RFtcPt4JPDoFEcSfq0vwcpNc22fyI1EoS7XyzooJkYn794IWWTWoejnOpw03CrT
/WyZUL3YqyzOXpx6HEtBvHpyd5FIKHhIVu7IzrNbhgSfj7PPE2n1a5VkDc9goGcW
GBy8OkiB+pt6z5fbFjvE4cgS98xBXjFRSCvBSSlP31pS4Hdq+biiJoBkRrspwoHj
XeM54ylEkXIlXVmK3mp1ojB+rQeF3/fuhH/UmK8Uo0dHwAO1TGuTaYu0EdD7D+vA
Pv0LFkGziVKnbpwWXgDSNEHZR1AzJQHPkaKc7qvv3NZZn9JIJEB4nZHdsfcj7MoT
CQWNDvC8ig30G93rUv/ObnCEneRHQHLsVd5nzYpm7WCPNnJeOtASWzSFkes7qg9S
gJWZf4ZtN93qGoZ84VSdas7Kk/cUWz5SlDPQNHx8DJU6lgY+vvGqKRrGbhQ/E635
wOuhika3k8OuYz97ksOzMIPN68RJH5qAlCJwKYLShakGt52eUxnbrtE75LHjjCXJ
gbfEwgFkGlDsLbbb+QRDuZqpnbvsQE4S8Mkr1vfp+cOJ4ERxko6/eiD+GJOQv8ta
L0nLdBE9V5ph5xwXhBqPExYFQ13/eMe5i4+O3MOyEjKPbrjz48xgEbPrgVQKeDLL
aUXf1eDV5u78tK8zlsOD4Uvltr0d2o8bu8Wm3AmIYzlN9IBwXPh3G5DN0DldDUhw
wOL/+YK7FFHfSmWC8FjnIPu0ro7HUWiQ4elJoqlucj6uS7POoOa40qlVtvh1fyxQ
OR8bPbSM9yTcAp/0G/84qhLWK08csuFkXidwVZE0HaWdrwU8qjIybD4iyyvyAivm
lJzwGqv7DwaXkwGp4QnX76q9AqMgXsPwAT8DjpxW56BKeL18iudsGr3mwk3I4AXp
m7oko8jAfqU8NXjGGupls9vjNHiK+MY0VqSW69Ac+eD2lOI5ZmjZya2FeyUj1PYB
HN4bl4HrSh5diWqhA8dk2qSpVcMKK3JeqJZKz/cRqtroKxB8e886laWftHAU10cF
RXABJLkOsI/y5zXiSHHtCK/xqFok8hE6zU+w/iitawTclHZ7m1CaJvHYlCm7FH2I
JwOOCCqJ2U7y68zOGR/pPZFL7Bd+8a5G6Q+09zXN8qFzCH1iJRg819VUMgFy96pQ
amesdbL61YICWxBHxXi5o1/7wBqbmhzIjFWGn7hEJ6XYo5cfvht3o29tLCprU+jC
ZMgbxgLJN7FfZ/ScJ8HGUHkA37aHbxEWo4rMOuZuqQqzT6UaaOLaYYWGmFQmrALm
n5diEE+JiXAirDyg9ll8dvuEFrfkHD6NKj3ppfn9QnoPGELpDxL9vn8pjqF9z3si
Wdza2zwPkWGijc+2pCVzuglNkDjHg9vVqTF+NKJb1VjVSUIwATsxHPKZGN9uAQbL
NTaw3dPtf8RKnVXdRE/oUecvNKlBlkrrm4dgXH83oZXKh942e4VtGyDH1KB/0ri1
nWPUVEhW2P9zWLUWcvCyMTYHwcfseKXbn1RtUsAPBHlMEgGgHdrUYW3lcAVviwGK
714ztBAlJPsYaTN3YkUR7JQ4VCf60si8hQeyBaA95+nSlFOsc+xsufmoJIA7UITR
5ZYLoCDGFTJZp5fGz5ivPW4J1BS+QCrBYFDcH2wiH13fR32QhqwQJmzdY7w1HGnC
vetTR4QBzTOV4sHAugsvhGJaDCIpIQGK+CorgHxk/Bumk1y2EK2pHEq0fmgXckxi
YudRYfaSzdCitEn7Sl3wbxJ5h42OjsbCM6/pMYMQJ4TQ5u9zSkg5pRBxMIC/ZgY6
fiq+OVfK/BnymlYF+fvCtw8Ec8uPoCl9gF0wS20t219P6zmc02syoH8bhLscD+cA
2l87yXJhxDjZtNwLThHrTEd5SVIGtT08CkRZR3XsLg5X4wtqk25ULf4L1A0vW9I1
AFaUWMsfytW6mw88CjC7bpqVLftxzXCp8xgnyK60IxEqZcTyAfBqxMNk2cJ4H3ra
6QTCL4Fv/b674CMZYldXxRNO6CHn4PDWBzfL+kH4HfCpV0k5zEYaSMgXMbqFJ8kd
inS9q71iiNJwnMWDLoaJ4RZE55yXmBlv1FkrM1pZgY/ud1QPnd2oVTcrvSKmOKUd
W9MIEyn4wg0e/pyhcqN99bd+wypSRDGrd7n2QlETz8LcFolIEqIkwo0oTCKdvW8x
wxZ8wdlw1ctkKPr/KXnZvwFWiowzZoogQyekUkKrJzHtwxkcK+g8bFScGfyNFoFT
8UveUCoPpd5J9ewWhTdLruvm55d87WypsIMMxHT+gKGuEnjHY+z/2Jw42wegylAN
mpPqt6bWF3/vw5fiQ/xkmF10PcxErkhJkpHSiKq7314an71e0WEq5t2WYlGrtmIs
q7Ch4Gcg1WvpGlZbY0ATgQXUI1R11vmwvrUY7zhYolJuECozGyplkZbWo5k7Aj+a
P7IQ4OMPSx6DRz5MQiJRdo04+WgNXvXnTcOm07IKQY0FHhI8kRwzbuhP+s6raDUX
WWVAx5R6s9l/ucrKadzCMzbCa2as5zds7Xm6DtyIkerEjQqwyyxos8Q0QocvChPS
l0ZQXUO/hf/UEg35adGz5aV6jU6A+L2ytMFtalY7kFWfEe9mnxxPqiDfKhq0RoBA
jNPbQ1t+LuSsrXfKYm5JM0Vgw3FO50Wu63cjG3npU3x3VKoVwiwp9EteuXruRtxg
MtOwlf9DcIPSTy7VuCmkxgpTjVHM6WNsCiRMDcrk+H/5ErDb18qut5lyeecSl3Uk
B6SAQpcGHJGzm7B7wIHUKmSqKddUOsIjJMMidTZYO0Eh9fKQx42dFtiznHfFfOuL
NUZoBEm3smQu+fad7ucBWgGSR3ra8AOtkzF0ZrgqoSR9XGKcVLQgop6FP7cy29dU
ukvRdTKx41+xRSC7yARKN/i4Qack4vBHP41Tkl0I8pnCxDF+l6CuczUS4j/dT0ml
gJdVN8ezx0s965oGl0p02Lxyg6VSgHeYYg89IUJyZ6YGnwGFkwTu4FhicNii+8qW
2X7MtnsXZ8xCgml7ZhMxcmK+LjCv5DNFPHelPW1MnYN7YEFM2jMQNyUGawUgklJ+
mdaMpOKXBBJQTlIwt0iY7I5TlGVJgWmfbmwgTYwAH1Q=
`protect END_PROTECTED
