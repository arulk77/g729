`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePESuM2n28GveFondiXTM6G1PEI4fheGTapagIrDYBqp
YTw1oRToabRl65DgpvOby0H/g6SZqEmabn6KSTVKpbLoZZmp34zvEgINbe2OneQk
po4sStZJJ1AFI30khuQ5stUP6980UnnUuhlsT4biHg2gk43sBt+ZlBX0OVpnwG8Z
ORSSNJzVOsTHKn42pyx+X7L1WmPe2yUcqsClvolcNWQyhb/UWiQ9Q6bqAZ90Gbs3
P7P2ERcFDqydQdHra1kX29YvDZX04KH91qoW+BpSvOPGSmE1f7fvFcOwONtJPRSo
iH4ljF6sV2KZ6Yl/q6G0+A==
`protect END_PROTECTED
