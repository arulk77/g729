`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wLpve5xOvaRBAwWc+e+bQzK6y1DfWLF6kCSVbCX1ZHx
OiMbcwOv56sa8Nz3XBGud7I1V3u4ttD8Hf4yjC1Bc42YhYdZtMcmOMVPA9G7cTer
+BFFlnC1M63UuY2K7aDJpPyyYmfjgVj1WyNhePKWatbv7dGppfdtetDKisuTLD6e
J2nV9Kh4HYi7Q0XqivpS9h8RrXk2f/FSE9Cek4AWi3UFETKutuuy6y5OiHDfrzFy
LgX+NJqwFll+LnN2Mk8stAH9Z35hKJScKqATNvYYaeI=
`protect END_PROTECTED
