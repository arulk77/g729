`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu417HXcUnXXe6VRiDBbGoNEsJHWRROXJNo0LjZwD2hfIo
l0cydhFVNaBFkR2pLJeXD9yc+d3xFKnlpFgHAvAAmLKhv8juMw30WNjRBX3cm98l
EZnyWfg1PH+Q//Zl0zbmSyhMFAMWI5HpHJdoEM3xFENP99wRykS2p8OaP7QRm2Oi
vXVBDP9Tk/fWuYf1r+f4Y1Xwa9glcX/tQN72+iS8lkwnUoJ/z0jT0UGn9b+TUdNL
dhbUunh166NJToQ3sqpv0DKsbirV/iccDiX0ThzJbog=
`protect END_PROTECTED
