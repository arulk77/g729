`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL85J2U6KCgO4On3Y6PKen9SflezalsCaAL1FXtn8OLYdT
Rv0tApqNcb5IgtoNkgbrVMeRMImXQq/WBBYIvLPdIbdF0aagzlLd3UfjdlWeee5/
fgAQfVIDH4m5Ge2Y1yUxR9M+qGiCX1Gv2aFV/I1X0iGfghen04+EcyW5mFtdxKsA
hQlk7jHcjywyfI9qbfqyOIJjzgMjVg21g0exoUllLiwsrSNMNZcAQkrZuBk0gmYL
IH8GocxLSkgpTLA9aCbUnqkaBk47FCxm6epY8vqUTs8+uuiCNnaMv6YCeSU2pny7
/tNZ152+IHWV6mNj6IieQEuoMUFsWzHorYNf0omVwwEmzSAxuPMNbAa+/N1NlpXO
jeh1nHhWkpIwE3kySHXpfxvquoM3ecZFy+EKrfZkrFU=
`protect END_PROTECTED
