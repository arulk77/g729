`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1abZ9+vOBY0r2p/T3mNC59w7G67ITSAcKMl3RGgPdbw29
TniktxuAomoSGoHPOlw7XDMcHX8Q4UZrFXaQVZ/xhgseT/u9vhopHe9P3xixK27V
/+6Vj4xKqS1rXHb5kN05tT6FyaNszjwp3U92NccQZfTfcNI/G9FcZ9Vl272i6tQb
GloeBw5lT4+2X/H811kTirFJRNL7jnmwzPsZ5a0IK0G0sNOrSUgwhqrC5Vc/776e
c04753n8A9THZ3xaN29DbMJFPz7KnJi0z3N773LJOv2Revv5TszodzA38aRxGe1B
sDHVF8oyQczciM9p/pI2psiJXQRR0FCq6hv5Tq1HJnVGKg9Wd7xyWHrLr8EJTRY8
xPrx/6RszxzUyOPK+r8GdJj2l+6r11gSlJZmu5xyCSnYhxw7Q7DzPxjFMD8xZIXU
BVTxsTQdC6GH4ideGaXkwr4czKWu7vhIdF5MIgnrAgogND0HjvKnZOINC7VCdLoP
PubQkZ4F5wo5lY+x6yh2adqeHoR3ARB/yG2oSckKvkQU0lGsNVae/uOwpvxl8lq9
2ICgpgSXZOjHT9wt+gFJ/ufE6YwMDrHlwgtyJ76+uNXMp3z+nSzBwq/cvJkSXbfo
XD0dyxHVJcNNLIWsViq+Oklr2E7ySiECdHphbT+iHVNUxWbUBL/e0ZUvGgI2G55L
aSbSBYoQ/KB5CTslANIZKHI2F6ISv9mi9Fz8GT3ppp6xqKvLTP3+JChRUDdABE0y
WVhdW41d76yk1b1P+QD1tfksYWseb3Rs/rrRTolXnpftzznrR6htV1X4uOg9AJdv
tQ9w9A1VErkABGrEY+emvmROvrIMewl0bRGByC4xDrknQk2/q9IE7C1Un9iFKZpa
Kubm7mhF0uawU9vQi7nq5RcGaHLNVN0E/esCORO9g+ngC9ZaVPKpzHraeTpdaUXI
MFNfW+rKsb5y+i/Gm6L5ulbDxbpxLV+O7b6ZhQhl1GW4voNeilxvOGmOnFoBYVNy
+o8Y7BA/ydAgVhwWjNHCJUd2OC1D6oq4aMojZdJlM9Mpa3JHlg3dG9Z1CEb6RNSK
C4Dn58UTzJi/CnqJmz65RQJuk3eKff2S/4b8p0egbS6+tYAPFxusU4nfB6xlykEV
TRB/8lhRkveHqKYEx79f0f3C3LH0cS+XQpADWfCnR0e/DRjOVb/MnOVtNV9TRS3y
Ark+g7nyA1FoIe1giv1vF64AhjuCAzmxk/oBPycfisQnCe4oB0+dL527bVfCFORY
xMnPGM7+TlkQakj5bSXIrfS3fOsJwYKQaYjZlQzCpvI=
`protect END_PROTECTED
