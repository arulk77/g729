`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1ab//8JSKsrpv81panrErcVJoeGkGtPWlYaJ/JW/YCxUx
IBipntw1yhONJsVV+LjayV3tQTN6sSK2r6dv16YFNClzrjrYQdNlOtn+71cmvGGW
p8uXp4ePVSqZZpzCmftxyiDqOC1srAUeRckGCafb8T4ClQU1xdlTo2nDGSuHrwQp
IAp4cO+v7Bla2PD+u7M4a/6cuWjnDGC8E2ou9mOJHVU4BL/ZmyPcgnrrwxQsmHOk
kS5h1x6tCoGG/7ctLA1P/CYA5yulGxfppcv+8Os/3bsOiRPn4il7IW9onZHfpSCx
8pG74Lno7p7qs7KoKwzh2+BSDdrnqSM+YTzzgTgAHE1fzyutfnbcIcPzmI+i2Ouh
`protect END_PROTECTED
