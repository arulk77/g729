`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOclkM0ROJA3sV2QuzO8nxtCB5a4Vr4KZoNPajraikff
0NHvb6TO9hVBWmmw4Zb69qrEeiRYcR/LCcQ9ndvsjRMTm10k7BJy1PQXJxtkgLgO
CwB2xp3/wr01aDeztK1Jb+k1CReWZKDj3mkguhE8+1g71Tybsyp+SCG7JbSeylpk
UV3abJKqsO9b1rIaX4u2lRTQNhwV9/X64yQCdgaed2qagGIDmoJyb3BLJUsIKiES
VeSxd0OJ9DLn1h7VxMkclw==
`protect END_PROTECTED
