`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDQZS63bDHJKj7XDBlYufwnii6LIocExMafYkMU1uYX3
s9dVO2q+McxrJbQMghRktwhrW2M0dEeOFL36lJPrOP4xqbKSDl6Y91YQbzNK+RtH
BpEFTZAXxkeOjWIIlir9pOcNLc1uBPsjYSIaZQ40U0D3UDSuVr0W67eq2ZBchwsb
Epz0aVjt5fuY7DoQ9AY4e7UTVzNPBBjASsFeNM/83lACOiCIvyV0F6Rmd8hqdhJr
ChSNfPiziHr+zivQxM+22M7noESZCcgUhXPPlcWDoTl/3xy10nSxALQefXpQruTo
ojfwUEM9ZZgzqKYcP1vj80cE85f2YDqT4wZlhGJFbATB8r6c+O/KP3zh5/n6h1FH
vNGVr10zg4K3oVYWBHh0AMTj/xRetHlBhSM0XLdmg2kvsECGmPv+QNF7a1L8bCYA
Yu5rH0qcHDgjk7a4dD66JQ75VhWuyM8vzMF1A5xlYA6S3s+AG/OhvIhCqIpjJTWL
CcyLfG/lybwC43mqHp0m06CX3ZMDlmm/hKX+mPOze8o6NiSM7bkYhKLunlsOHHkx
OekiiJ7Nc+ugbLb+pYqVgqAzlOtHDn3PYBaiPmAKpxKUoVHwWdlYKD97TD6bfmHX
BxTHLeA3LKLUH+S6IX4KQLP6ZXBsOLdveuFHX8vfqMVudIi7Nj8S5HsRqz3vaiL0
36pE9UKvQ9wzIhMqtSoga3KZGksQZMJftkeX4s5XxwW2sten/fvBUFoGeXnP2rn4
rQOobg35QeQSwnpxg4fT/v0ebvwbBlkAcK0C4eBODqrGkF0764B/+EfFpUWBu34t
BBoAs46OtJw7eXqYFZYTmP5ODpZ5fh0Sw+m+KVKrNbE=
`protect END_PROTECTED
