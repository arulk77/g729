`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEpSv7myuR5lg8i57/giq8jauqpsIcwv6H110/nykcZm
4OjyXhjSSf+kELGcDcud7WOQrRt1thdmCKnPhPeaxKu+c9Km/wAJMdW8VoKlrwK3
KPrJEeonM3R4UkyKTu/LxxWvfBGFSSSGTku3sOS27V0GZEu9Gqb5+aVA7Y/f2pal
jPESOm+keIWFUMvwlOTYIrzRDWKHzyOzzSyruU71TWM11dYEgX/ohXTGA5+H0MhH
h7538DxPUbMF/YF1uZGyzo/JYoy+isHXHq5bDLMISRlvcY6KlBYDw2c9s8v2U4fm
mhlxpf9J91Zdo353G8WF4kxNdIpafwpLkWzwpAIzapP9DRUc5nPQmrk6CWFZFH/5
KsxL6YWRSQ2q5FL/oWfZRCzRq+054nx5Ygny+yYMHr8IUNnPLds2SxLwHY0j70x0
UvJQ2+lEPIeQgaUzFxx0ub1ZmOyiRB66hJu1DMkzJBOJhxYCynkxDPF3DZBexcH/
PmwJHVisz5zpVCYMqmhKLyVEapPnRJZ0de59PFbSE7c3p0XMeuhIkyxwCT4CbYMm
`protect END_PROTECTED
