`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMDxktAbl2PV3o6+xvsMZvYQ0QGuwPE9BiIe+wz3SNs/
CmS84KF68N3ifK/HUUj4DmucWBylJRNniytcUVkPGXJBi6HomG9/chK8yo2d0xUB
+9lti9ZAy8S/Xo10WcXeZV1W0Wg4wAKth3Wm+nt2X3LAlFVo641ie/7/TaofSBij
4kTrpgprQ59vOxO/uuaxQs0L1PBZOSLJeXVDHDK9DsjuUyyuqEwwmeaAo719Qi7o
3+6Qc6EMc7pJKJO62ewFD3Gccqe68vMwhDNVr9cwl5dtK5SIbh2E3xhQhSaIZx25
0cqpDyJa40XAd2En6BJUZq1SYiLniFwDx4sg3Uagq4xLHZ8Nz6Djgrf15OnqpiHh
y7TbjlpC50rO4Qi0fDs+i/YZmipygUhYQ3p1HaRJDG+xd5P1nW4U+8u7yUB0ZgjL
IQ3bym3D8X5KzDl34SpDy/u51JsUjAuZxjLukpW02Y/kGhL3ZBFe8pkKjtKHmpAE
DKGsC3XyIjN4Huif2ccDu8NZLAH0mzqHE+JZy2LHao8QR/GO9bu/Q06mMBIAxlss
`protect END_PROTECTED
