`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
d3YsfdZuSKfKDP/BUY/MvbJrCrAgkRkARUNBkx7ohSkkH18xAIdJhpr3ZlWUVAQp
aMWEgE3mFYd0pzwa5wuDWFVoR8QKY/tJCF7pGXiSrQuF6EE0+PtWghcawSqJeHC9
tbojxllnp4OQSuTfDGb+GnEu67N8yAoHW1vErZujre3KJn0YWjkTbDc7xSDYttUm
NyfH5K/5mesG28XJKu9qOniYKCi4UcZmo3qM/nEBSI3euARMIWAVbA5JPuU8xEML
OcHN3osjYGRXZJ3/UM+2Kx7aEDYlYPDXzUeE+okuHTcttsmmCfAjLF2tPx7sWXuC
NJJ7TRJScLd7ZFZeMH8oMv07O8rJJESjWdpkLO1BMRje4sdYlGgijZx1FBiNoleD
W7CiI2v6K5QIbY4OJCCgZ+d+DeOfz6hqmXzbP5/ZlfgBo4XysQLtn5mj1XnagvSA
qnzn/sFJjs4ZVU4NAslG/+mED2FdsGhTRuG5TpJjQ6FiQkyn7zBU0dIEyQ4KLgOX
TnxzFEfaCiFeDq7ANi2y76v3X/cnaSQ9dj/yr113wNP0Mgz+tGfuhP2+S0ROZcvg
g4YxyFu1rJfp6CfC2yOeZoNwp8M6LU5rgoZABZLKXFLrfBIweORZIb/BJDR5Cqkp
lpwdN7bnPQG2T3+7npPdthQteM54bNgy5Ooa0ELlKuNCMJvQdgotY20+Kfl5QcUd
zeRxaTB+vctlOTxwH1WgynH1Lsrbs2tt+Q1XoBPbCulZj52buz6f4vqRE/xVipUA
SVwZnnoJX2Bl/dIoJbwMpB4bgIzH2arE2u+Wg8ckysjz4qTw2U3Gyv1T8b6TEkv6
vodqpYk0vrDrKayW0CmZGIm5NBpUT/kaoiFrgB2y3nYImcA6AzCMHwl41+tVQnFi
J7MVLQCRGbj//63hq6jKkrq5jQaKDn8eJAkbhgUW5IOaBGYgmSy8Wg8ZeA2SNLBp
oyIO2zufj2MNe5HduywdxZ54eY/aNWp/K4dRa3J9RtRUOOiJ1MWhZzXAZX+7wvtF
hs29R056OVylKD5DkDtea+rLJTvVKtfW3WJrwCgaeyR4CzrnKUdrnMvp9l074V5z
lDpkYs5Ja+zRJVv7jXhRGcJmC3AILgj4xafjt4HqJ1VEjP4ABe3F2pKNbWfyY9+a
HCX0AtSiXiHjW/dZEMOkKKVM8Xwsrn9XrNa5O2pFrdejbby5kMEcB012ytGS2N6b
ujKdEF3UTMredw/zPAlzZxfnpBKDqaZc7mXnnmuK8AoIfKNovAsVsp/IG48Oq37m
gNBcjGDv5SxbGmrBtd4HfBqvltEZ2OYN2dLMszy4aWWJ+iY6E49Zc6n2y3KIlB+Z
SuWlFApXnx6KisMgO+2qUtV7aZWaDUdiD1Cr8Vkf0bO18D4lSZ17KQouULuGvrlU
ZX2a9+2wgNnmmCZuuEqGtmnDY8T9R1IjymV1F9vEfXUm+FkeofWLbtrzMxgUfZgS
Tu6Y4CZkVmWfvv6N8HZrox3oRTYIwn38nhrp1PZvvQcMkGdiiYb+b1gXKivsCj2W
PTSbpYO60hGLrrukpJVBkG64FCMXarVWjmw0xvWbx03r1fKdYLMtnO+cE2swa/Ot
/l+sYGYpqhNeS1Hd1kVU10zLpEdcvW8Sg2rpFup+29y0xxhPGgnM646a8pC9FaYj
PK+BHvpLDy0N7nYwAjdBkTORfYV3U2SvkW4VCenDCW7Dnc5D/+FK8ztesY+cKg5f
T6h4ogLPdD6eQe84AlYKco5I8wi5krtgjrntIgRLMqQpyB9dDxkoNO9CT51yg1x6
7RdBS/xjS2gGb1biZT0zYZNA0J77Mm1xhq5H90/u6WH42xspVUbCHXA+oAMz/+QY
S6M5aSbIi/7epc6mey1064XOGpjtKLZVgVQKk322Eyd+1kJzo6rAH/N1jmoeWGzV
FHb33xx7BeLnGOuhhRYckUyxzaFLCkW/42KXXQ5QQuIW+/alt1yJjIrVUTOnN9Uv
08sIUu+6rqK8v4yay0RbjD8C/6LiGrVxBmlG2s6cTmo3zQ9PzzpTCkMZ/xzpJboL
rXPxU740YKZkAZvghOD7DN0QYDi61kSjMbvndkQWrfM2LnXs02ADDmKIAQX+j3SZ
LjRlnDAra6jcRlV0XUMjHmv2R5Bm79GGSq1jDhamp2djd+ZrN6WYo9ksX8aUU+c9
Jk/lrn5CIqkPKJLKhKRBmYFNpF65bkPJpzdfecbvJj9obWbiAkofeLGiG+BO57MR
dDFgcIiNcsbYRFk5fQOVQRC/549zjbWUZL+xKcAGflWa9XBd6nmnrzYOBYypbgs7
Xce0qcV0JJn95JagZPUhAg8l8JhmOocE6A5mqRX1Ih/gr/ZSTrSygFjHrfpy9t1x
wRy68Fbf49lFoqXwbHSlbB1lN2oXaFBLbt5Ai32C5y3vaJ0r7MhGeI8UzpPJHtyY
RJqDxYjt80UnYLUjK8wI3t6dnZUkbkMnn91mPGJZt8mKvgX4iYfmV9fM3RP/C2I8
of/nRjdeQMnptKYpUw45DnOoHBgPQefOryPmYGYTg8YXDb9qMJh6ft1uEJmBeKNc
GS4P5TdlVhTHaCbDESQNgdGHowDfxGD1Td6EYFi/9Koo/BGus3DBOrtL3Ol+jHEs
RTPvYkTTy5LWAT+8eaMS9b81pPPVdIZj2dp/H2MYaO8v3zLjbjPNWNCx5gbbyuzW
6y6aQt8xqcjApSO8BpwK36Cj4l17ujfNT6/rlpHXyaX6gtLrTZSS+v+9vV8nZ9lV
I7UDduuwL1cXmaEIBQ2M6lU/lW2BjEPl6Gf51beW1WEa5chJuKWPWd3JqxpcQrog
GkFQLTq//s1/85YEWHXpaVsPjbTHY8iwvfX3kvecN4CwezmFC5qPE8FoYAg4d5t5
zLpt2oG21VjK/lk0DXXiW+AYzt9aZ4IdUgEj8xuZwcHdkHXV9+5fFqR4j3ksR18S
++8TMU/5+NWfPlg+UqrRB6+5pcuGutFKDN+cDNqFa9U+Yh65cWvqF1UViVT6BO7t
Lx0KL9jY56ex94j6YeXgcclNrrwJkoHT/0ZvyroozjWoPO5dYaj1WvmDeeeo1Blo
kYzEUETwsZXlTWEzZz+i5z5BzQv60B4YmxJoRaGrIEkaMscYl9Rog7DCrv9RoRa+
QsJdbAEfvinKnNdNnCWPBFZTaDSYJS8xfrQr64FmtZQCZYj1WdBaXZBZcNVzsSV2
wlVA5EzYOxOtWxF/KS+UtbZIU0bHH+rbiQrouVo/XCa1Kng0B+NuWdGQ57MTbNt2
1jyE3vR2ApDQCnM4yLsasyUD6dNW82Bby1mckfChaLuXqfh1jQnNuXUC+KNMAIVx
BUELeXYCNnYZXkMcTqhTCCR6VcGi9ZeqsXNtwTG9xZkxSBB1VZcso4dztPVUcRGo
H4IaoM6/cUj7BuHEcYMVXlJWRtLpSyPrwFmGax1GrThLVdyGpwpeT2b1qiuSdmMj
yUdPa6i9hIWOvDnKOeflkE2OJ+K/ZIBuEi8fvLRv0Cl3yGwyMhcsBgBgT3HZt9zl
IehTIrN/JoKNI1icqLCtXxdK+5QmqNsTFuItCiK7j6gNL8i0ZbPLNjD11RWZAa1C
CmlcgL49B2SejBxXgqNFEbHfvQ4Dym+SBd4YwfhQo33mzVz1xJJ+flBIYokSCSJq
EyYwsAGfxHDp1XdZJFSiUtDH6lVDgBmcf+wXBEv8zeY2DFy+Xgq6vw0oH1iAv3lt
A1qGTxfQYieXRW6rsO/EgSS31KKbs8Ectg3rWAL2/xLQK15sictxJo6ZjNXIYZCA
DIqUR3tmb+QV9zdI1SRkslQ6qt2Neu7oVvRLwmkaU2Z0L8sOMkSKNnP8YKRhocuC
x6p0fsOUjJ3+aRy3i26yX3q8AvjqKUB1q6amCXKkqwbxa7RCvyWIN0HDNYpSC2Ez
AkA7TmFfrhQS7oluF2yidkEOP8EQKIcwQsxck+cCzzHZwAOOyeVrmtqG6+MnoLfe
M8YpycxWVQc2ya+hchd+ZMN0Np2BrqmHk3IzPZzg7sYnQTxGSiwqKYmCmQVKNN/0
kEPUZbwrzKBUox3yyeeDNDYFC9RVTUjNaHjXDEcF951VggWKyfCOxTevPcNx0MEa
8nQ0y3YZvJg3UgHPjCimB32QaBLJJtGRh3GAVb0OZmVFZjShi1KIf7GFykf8Now6
XxDYZTIaQC9nZhvLqtMpYViYs7/Y/+j++P2/ynzv/zz4uWDLS48QYPhoGFSngvY5
y3IQ3/kdchHBiS4eVmrRdBhVSpxvrUFh3sTkhWjXYWVpdIjU1hasxUEpEV4ge+jN
u9eF1J1ovzVhwUfqV4UVABM+xOczF5ftald1706NAlq2Iwxx1/x+sKidKgPxat1Z
5hjxcgwkr4PoPqeCrCe4KUJdRQHWNcCCFE5IQI43M89+D0htr7veuVumwYOVpoLQ
UaZ/Fkrhvgj8W6v2vOnUukcJXDj9EKLjiML+JPr2r4Q5Xkylq6e/PBUt9iTuLSh/
Uf6GbKxvfouIXlMBcJLbVytJmOCJa7eQsc5BCmW990j3e73TDGWpz3RxTmcxXnKj
keASTdAgKFq5Bcy9NWrWsxGB6UfYLtVfE6pI6oEHIGetnBcUAcNgcOSIFgmEgGRk
sCql0hV2jxsyC/B2g8DV7h0I43aTHetUO4TxtWZZQ1FAQkjIlaJcwr/Y9IzX2X9t
Gchet3LppaoF2NZw05vy7lh5eS5cc9GH2BF/D9p2kGOQQX2CrcMeLjSOIwZhdLPI
aU2NguZ3VW8btOp0YPDDkN8Yl2qj+UV80J8haNV/CA1WZFx/Oewnf/97moon7chD
Zb9bKzk6v0D5OZHlF7Kn7rYLLG6+wLO3JvDzu+W5QVRA8tItkmpjTSEmeTDL//Z+
Wk+vp0JTci3GsGvVUpivw/qfwDZ4+7kkMZFrdu3jugie4ipHyuw8PRtliGuuWFGk
O58QSMO253uFIBDDyMQSM7aETjAtbepZNMgTHhaFH8OzSWdOdMsSFDYof+1pnvCo
m/GXaHpBEXhKaK59KeYNjM+E9Mi7sH1ZO9mw+d+KSpX06xfn9USKdBSVw6qVtcaJ
o1m5whxIuFMVqFV6JisD3Ul6BvAToVrnsgXy78lT6myVj//6EYldlNlMRgNEOB0T
ehmvoU2SJDfeIcTQuCPWK1p5i7Bw7C6TY7ujSQxcZWSWAHEVS4/9b5E8Sp5HSyTx
uMRnLgQunIHe3D8K3SXtdQfy8FanPK7O20ZnQ5EFM/oGbSOm9PkFv7jgRjGqSJ6I
eJdJvfbD5Gi+msVylTcXHU3Dloh9I2BakSeDAkEt1aqLnoEr4Apw7ER83/SCu2kY
hOn2fosaIjLk+dv+voh5uWmirl0dhbSi1biKe6JmoWZl0T4yEsb3xC1PWeccM9Ii
H/OCgO6LbE5aAZXLNY+0zM7foJT3GnonieyG/beMX4wY4bsqUX6mrrDb7jkjxplc
YdKyMC52nA1eS7aexRXC2fCvLStHUuO1Fd30g4e8oQ4JztdSElA5Nr3sVAV0OOXz
naBFKuaT+croblUZqxu8uv/D84MxF8L3eeTD8thVMKLXcEdusk1SJQGD/pPvkL+e
OwYE+UG7SWQtUu6aK47uHVmjJVZQuQCFJFtziaXqEfRc2Ohw9q668j2em+panzKL
FGIy9u143PgVNfEtt3lh/QtUnEDQChMup0EzLkahpqZw08KaXecQFB94tpBYqBHx
CqCZO+5OTglcyMVepLJAmZkzb+Mrv3xtFlICV09E3zTuKGLTZs0qFm665BU9Kmoc
5hKFPNQ1Tb72mYomjRPX0II9xAXusUNVuynS8rO+mK9tuZ6XOCTZfSvyfhQ6cgya
69iccYGLYrOLzdY7nYFIGtVqWT4P2Ft+0/P8kklUZVjrs+ALdGdyelqZFJ4nGEln
TBy6Bk5MaztXztgLrTxdgiVsN7JePprOdF3OtLTrtzlakxiXAAMKmPV/W6Y1D8Wx
virJcN4NgQtV8qk41MyUj+0mKoBxZsoVcUjbqP9W8qWh7Pe+mSgA7lKaBF3gOIjb
8WxUM3yKhK9FyloEOS6Bx8pbRF5uptBA0puWY9Tx+wa0dHIdTNPxnngr9zxwZfqE
CrbQSnlN/pji4AKbZnkTtPMOeqWpJSM2rVhUjbQYqfIZwwT50GcQohVnl4LP+uG4
TU7ZyNmKbCJCNBNT8iTye0BKMzhvLPQXyRgrZWouOoe9A+P94zTFT8gZVUqQBz4q
odoYmbgNgE1iL6DnTvBfHy49sp+WPNwEY8lqunyhFVrGjXSU+CiHraQIsOt8NpHk
X9Ew2Tqfpt3ErfBg83vupIFJJiMlZshjRCf4wZ/ZJyXtrmYsSMQkeMQgc07X0/Ej
Y0U6d/39sT+buiMZKy8K9gVMBMBQ3UzusZoH+fPASKX8dXmNHx3Am/b61IpkDH4E
5+8irsh0wGHawNiAlglAwyXgmaLoGPSFF8lZyNahcKQcpcbmS40yz1zbXJnDHRvs
6hV8QF5uSS8nqmL63EENni7oNtp00iL93lg6CFBPw8DNT1lqCNYrJ71d0Ca6dC6b
MB+bCoSf0KHg7dHtpZKpHKpjjH57DMOxWAueVqOtyGdIRAe3e2EJoTYuXbRE6grn
suPjQ0wF2TNGCvU13NDuHTygONBgbynpb095Tta1dx8o9Je9wA7T0iZDTcN8coIP
Q6iSczXxgSry3bn5v8UhUWKLCgEp1FRFqUXgFTmjxlH8L+eHjIXg+2jn7EPxolp3
LQu0XfaOeA6w783S8Z0vkVB6dqzDd7jbHeRm+c9lGGd1M0WxRXWqdR493g4OleQK
rk7YtMB4gyBo2unSbKkvE7J1D5UViCCxu7pcPOYOSTQ8ERiQIRg6Tz/e7JsJy40d
CFsyKWjefTzb3pqAMotxheC0Z4WgPF7cRv4qO0AbqV4l39sxcZtz3jQHOe1o2ib/
9v2voq4ZGA1v7vzGKHGQHBXR+rLm23iiupU8gsoixIWQXCJ0OtIbtOEu9wiKdbfa
Jf/cFidQ1H8Uz41PBhiveqjbOqexS4F5Gg9/WbsVCGWanlMq4niJBMMFzg/CPCls
Jdq/KUOTqs9NOUZgbP75rbzCkGLu2l0owP6swtYkmHVsI8nk0ByNir/FwADJjF0Y
xqGLdgBNJ0CuZVEWNP/bMVqXM/G24bjuyXja9Ev8E751jSJOmYgO0+bLA8tVb7/s
kJoNCjz2VpG+lxT8jdKr8Cez7b6ZJcOD1efmpUvQPWD5K5iYt8v/kmTZhA8zJZhO
xntV+gM0W9wNz81nANr260KAkaxl/7cKJco5A84M2N8/+armj0Q4IIlfQzfcHuv+
PizwNow4lsUdihpUwNWveX27HHKbb3afWo6GVLghRdLFTJ4FL8DYyWXltbornE9G
XQOcN0geqDGUOkTGYcXbXq4zqc+zvoNLv38YiBuCi7ZRI6sf1YkcQqs4pryAKwl3
nh+c8GuIDEopWuuTgkFhi1Xzn+yuGIGKJB1j65Kuu+B+bCzfKIyGtNgMy+KCnCI2
5Y+P4Js8HARtWg19ckFhrJK6Pu1WQ5fkRbJcrcNJHvtnsdOj4Sdjzu9P/Wo429Qp
S0lnM9H6ypPVfNSVROQa9L5jEcnxcBf0s8VkZHZ/BtS/+JOMkzufKSIMx3JgD48+
ais7YtkC+wZ6R89HnP1DmwXfXucqvAF+mjFIW90F+Y85QGEcyh2RvN2qhfpAkOgs
60DHNlqV63WpnGIj3gAhtG623fqaXIaINIL3PQiwworC2WMqvs8O/IuIQAU/q/4a
jQSAFgaPM30FKxQKupZZxzrQ+T77e2Ob8OrpDnUAzg1W7x1dpw5zzlV2XwBjrqBB
yFCKogPu0qgwbCvBusd4/yTZmu/Xs0QETG4QKJ7fVHP4kHRUViPSm7nv8G8NvorK
xauAaFygO2q2ygKYCHx2P5u1lZVAGlIvN1fc4dQ9fpdazIc0pJhX/Uby2DcQS7f5
HvheHXE3l3ZD5wICKmfXkfEUxusQs4phzIx5nHkOV9nbPxex4wzNJopFIBrKBmyK
EAuT0Wreg7t5S4UH9P9bgXLLzREQm/ku5EACFZBHRUC0cbV2Tk/gUBdge9t+S0XD
S1m4WeXqW4yia8AkgqChaClVjhmHUlhif72qHoTrXhDpymwPFZWwwSKCO726jRE7
q5K0OCGutZKs0nCIkIfzI535Oi0yQylVvBgOey/TVPQOPieqmHp0VI1unv6ey1XC
wSj2DI5SSeLy4yYxnMpBlAAVqYiMOCY7YaE016KC/LcV0iG+5s+uKTgkDDAEvzhv
hF0x/3VMvY8IypI4RM6k4bNO5wPPg9BzrNBz70BH5uY2ilO2/Du0uFICZ36k21OT
GrhYEY8+x/7AONa6LDSnWTFePZz0tlVVkNUYxBcNzJXf4MpWCvLF5tpdyoNY2vQ2
OYVvxMn7EviVy/6cupOePHJWnFYq3jO11aDLWl4wIkk5E/KzDDx1/jP1pKOAZIc+
qBD3441ogWsGKMFcm5VyUGFwTUK6IlD+NVt/+/TAYEeD0awVd5F3k+NPj9kfe58U
YGD+f1yBq0YdiJHg2h14e2bRxPENyYVLOaFyyT2p0+oMY2av3CAzvo8noUNcVZ1d
YeoFfojjK3EmPsfaDC6a637YBhNe4UtIVA/Ox+A2CzBiCH9tTldQNwUblnlyeS1R
+MR69GX/1Xaf+OxHxGpcgHt5Kp5dAQltyhZL0EuPbeJgVHq4fMUVSwDdrTwkHOKL
eyhH2ZtFYq1g4c8KOf8fzARu8DX8egR9/jrFxNR+/lkFMkCv3JJjExCkQ5Nu+dgW
8felUhQR7zxaBjErxTBfBS+rUZJnohJo2nhXEBl3BqJGNaEde+HFvYZ1R0CxkSIx
VThHEuiLaBlOJUtkoW+052cIdU2ZJzLwH/owHj2PMkzah+EoQmPrIIjeB+fUp6C8
2Kl2+1vbiC1IN2IN68VgUCd43oP9eIPxNNm+2F5FeCJYhH80w9V2B/PBAsI2Eg++
n0SCZ+iZglpjuencNFPHw5y73sT4nTuXn8KvQJH8yixYzk/ulSBtu0MG+dywDmtD
MWF00GByFykEWZZ497qtm6oQvnvycFE0dfzSAOMP+LN62tHCxNWsF5XQj/E53kDm
TcYqLNKfokTW+bYnqEqaFar7eM0lP21hdDTCpIZ41ozjMtAM6sn/ZT+G7pCzKH7y
9OZP72LwDRyP7pYA4ewkio6QaBIA0AijhFm7ob7PCL9ULkabsHDls7RIsd81VM/h
VcH3FmI3D4w/2Uoxdrsj+bG4gHTpHmZyKGfWvnVZQZH19ivuSJ5Mdhr+1bSgDfzj
piLtbSSmyi27cbkXqT+AhKc+zrz9ELNqsLOBY6e1hKRKaIuOIzzB+tKT0ggnvJwp
ybVm+jxTMQ2u2EWLTH3od+fCxpSt232fVDRu5D9I+gTAlkLo/qC5GCWBolzVQ8y/
IR7lHnDm/nfKJkk8cgnS9vKgaUqzEtYO4vIVmaL5RlJgSQ/gYNMszcHolCA376So
HzQ6QsaHC9KWfZuup1QPrEcOcdcBq7IkOQfNWpV+RhTTVln04TGQrN7GPfLpjOEV
/3pAr17x+cXW9FzWP/Rygdtd3rV2d4UBs08E49sdqV6DJJgxwlM4P5eb1nUNCRnD
egHueiR5DUiP1liEtL8tflQ261f6+bhkdVyTxY/ugeiOthOjiU26GasZx5SGF5IT
eISptC+ZrzaTcWA2DwBJe4y+gRjaEB0sMwDRZseox6T/qelqDil9LOA4iA9VmSfG
Tn7Ah0m8QwVm3G9RB63QWV95ACm7ljAMSUPe7zHmQqXWLd1DGPkHu/oLuOC+l46y
tTK+vs7Q98ml0vsxj/YMW3SxcagECjSevPPHfCnJGNkq8WtzOGTDAj+qYyLU3mrs
t4tCs+iPy8BxQNIodQDOOZQFwRYJ62Xz3xwaJ5YetrL06v4Zujkcz746x2VI8x7Q
mxuqeE2JXX8G2RtIzBFt9Af1t3E6PZWbqsOO3gKjuGmQhrEdo40CNvdvOjDzhQOP
7wU+9GMw1VKMkndmFDFPH+H1HJtvcJPdxel8ZAf5j2abk8MwB7jzUyhiw2oViXnQ
DkOhJfXjwvEsoLzUBkPj914tEvvc/EDhjPdj2AnDp8y39rWE+8eYVXxb/iFRr3+k
HItuSlvFuZu9pFYkjw1FZX+RtsqpFqPaBqPs4vRYtg/j+JEk0+Yt+czq0F4QKth3
rmAsYhnqqG3ppwkRq20y13XSCBsV+E3TKsNElZH6+t6CHORhD37cT0eizm1SKmCV
dnCSq8AUK50ssm5OKWj2/tX019Xk3mmB1vzxq3BrzgUj24hNPJahvJrYs1Ijer5Q
CeME1nV/C2AiRePE/ruJsKaPNBnNyf2KeX/LlZL5yOIqxBZ59NCJFfVb6drzjrnr
MwXsWtvE+zG6xmqLbaLepFwPkhCU75bZp4vqCEhvHtCYs0/F4385JTapXL+i1HYh
8bDb9dbJSrxoJG+2+9JDEQ8iKhXeef78cUWhbuzt8qS7brWqxx0FFwDLl7mGet9g
KkN3e2colZ5D0dRkK6SRW4ODiKwjqW3kML5J3cbYLQooMKd9dOEzm4JG9PpigCUC
6j5npAL37VGK0T/faGN9A5y0sEB14E29s0mujxe8sBmv8LdN4ZdyLN8hv2Ze+MQK
BCQTwpOlTaQOcLy7eARDrFfCqnMF3Aifie0YCP/be6JgKZe7dMxbB1Z49ZR4jVBZ
tnQE5b8HjQC6XFA7jzB8JJbSFlXURQWrzWWYu/HtVF8cUKxkmfmtyFTeaw3n0Csu
4A5hDt9CuSzumVf0U/2MDMbsyn7SCeiuJD6p/a6XLwVKLCIoh12WmceiI8XUMQ16
vyv+j/JXS+BNf34RRogSFpxBccn2ugAYr4CN0po33gkCj6SsywXv+gMWvIX7MLVV
tzJD5hBPBLT71L8Je2mW/M4qpGtRGsL88ynhIJq47Z9N0Y7SoR8LSE0akUW9Uwnq
UiimCMIRHF+2R9/oaFVcc7oRb3zh0ySmqIU2JjfilXOWhCACxbchSZdjwIujX1Om
/lSwZ8srQVJUhcArouYm/Q77ey3sxyEve6ms0B27co5sdQPXevKWmH7r79T9jtT3
VGyRc3ZhsPD2EtO2HaPubOBH3Jr64VDcCzHcZhRVvEqD/KDSqT4UAxIaerWnfW/Z
aWpfs0zdaa49X0Di8bXQhOdSmwU1S4UJjXYoXGpvVbmkPPeP4Rn9w6rkKshCa0xU
g1aLZnLR0Jhcm7/YVnNRxhLpTrkTnnpL6yi99k26B39oMnE8A5jy6sMU5+ffL2sG
WEvgqx6pEzyM2sAF63glK68bN8xOLw6Fo/dp3wzxAgsoUj3VtC3hKGQnDo9QqYfW
VnTO8WFrljBvYiWz+khiHdIh43LZHtfEboKls8x3Qqrav2rNky4jN9Wae0K6NMi8
cbJprBIrYjGDSU6k33/uFT3dcwj8b3nlcsUSlrw+fCeA1klQksW4Gu4vD8L2riYd
VB7dvSvEIIk5uAgDcJzpwRdcxct1ASJs2Oiw3PbfnoEIplUbZwnpYIZxq5Rdgxa+
DbB9UzC83sDq9dvDaoRMaCT+eGGMR0PboWSEwrYAxUh/IkUl0y1XGK0dAoFaodaC
lWonrC4XkShhLWEQqP0oUNCO2AFYSUApJ83ruQL72mYRdBAXyDjnyH5w0s+Fkqyc
8eTDNEjQ7HcOfmzhpqHbqlMhEJCF5oReRlf1t3xKZKlFkVoq3eGBDJYKzjAiQ0gQ
aLXzWbCoUnUyxBr2LMEP/qRXeQQWFegamiHWk93QBK7R/Q3zc0HY783P49vXsiML
u4RBhH7W0KpuSj+iwdE+2rH3PTPkJOMXreVRsL8yKuMqML7yOINKM2VP7zb9ieVt
QFJ97JKDPSmRGjTk1nDkIoaK1QASPfJYaFG6IPf9h64Cv8yIhQicoLA6AFhnlKw3
wwZoOeZ1fsDZ4/l7cPNjplzWhJMUHNYXED3UovZGA7XFPgaFVqV+I48cNiN1wQZR
arDK9RhsJfr0iCvNUSthSO/Lia6HuI3jw8xF+ddl2+1tvmuy+SRtdsm7i/f48kIT
B47chcxaCbLrY/D6Y+42pGprn3ZTd1/p/0CnDFB0rDWcpFZldzZSPX1iYFM41ZoM
Smhit6CJNt6UN04YXrxtLfDMEGx9hi0CJTkRFBu28tM6vEhV20uFEqPwDdL5mhFQ
0Xzg0PY+PcbOUgPYWGSoILGdjVpIoPdO3+ojzt+tABrkpTfJbTqNbE2QI8Bro3js
yLElojGgYz1CmKTpX6YRmUjrJkhptEpFdEplm6bUFucPCb+ZNV5D1tO+P4Bt8Qfk
ZLbtw2XBbCU3P7f0lZ6SwtZ1J9+rIWZMEzCbkrteAytTyuRD0ysa67Haqidt5+jj
PqS0kPG7ladpwluebbs6ASwTc3wKLagFdI+re3CWESP3KxD+jcf1hB9wngSwn+/c
wg1qmiYsMHk46yfEQyth7A+et73fTwv27s1jPF7Q6+ao1HB9m0QCkFsI3oNhuUfF
dVq7jyPc/IHdwhOPCwUTCrJfdC2LWdRzaGsM10Hw39E5THmjnBIqC3R2EqQeTrX3
KZKeqEXUgrt4HPa5Tq3jgUBNSo3Yhb3o/fDTUqEuA/PTjGWH6Ps3fi4tTZ2DVYbf
c3Gg+vbrwKh5F6zP2RCg6Gh3W8IjGR2wv8lQPqUKauiL3dSXQ6OSq223o15lC4ek
wmoOGSh3p3bu4+s6bpN/aIEFG+7r1KOm/l+xreqmjh3eDD8Q+2cd1/TMjBfER23U
EWajIvNqj9Gc704xYilJI2ldMMp5upvyzc3U5NssLA4Nvmy1l0Stzlqo+1iIznEw
lWfjEI5Kbd3ihK6rUu3Rs+fFxO5H8T0HmhNWT6rMfTGgbQWPPoILAV4LqHjx3HbQ
emwnCws0wO8I9csVqFYms7SFSnfT4FdrvOwb+OwsargflzS1oeAbPVQ72fVJ+T3U
0no+Zy4NCG4/PRRGo+aOu4zfvz1uXze6hERQSP8q53YVqkQ5n7jLMu2ultvjqLzV
0wqr3wj88806gDysz+lb4oci1/tWow7+bgty7nbXy0z1tG0op8a4HuoqT+E8IAR0
wilc8rd428aSjZMlu3GdJENId5TxU6IQRpGA1waK3Z9YaY5NdHG4ZgnifFtWW9dQ
1flGInxcK5xE00bqvbW9gpxwP49WhWwGWCxpKIciphBeuvh8RcCcKOlsP74YTCoc
HjKfUB32rNsbwGf+WL7vgxMfwbKG///knj3+mmauqYapD7FlbWva7FRL8Z4LKoTY
yaSAUcbhGwEldTthTnl+35HO+0bzecaM+dEvIQmx+66UooaR+E2aKeFRFws064Tt
Kh6z8iMmhG2WpX1xBmamEjWqvq7iRH9z6rja7ynNLSrypdqXQJ4UtkCOmUbZ7sDM
AkbMF8j+vJ1vr6NraZT9UILLVoC1n51AdaAKO3P8xiVdgoUT4FBe+E3/qL+4Epro
+6zQY2gLd50np2TNE+5lCsv8F92XXrKQJ9B5HJEFJHAWRMiFzDuTpnhfWiUc+74R
Uoh1u+Vg8eHPTk+z9vloXnqyMfCHo8U6BMP9Lwn36d8BEi47PnSi5ehZPCGaXqP5
eaDQ2ZmB7XlaC7Mb9bG/i0ZGNTQ1NqEp3Eame93MMwbD7ddqmC9z1AQa6lZvrSIP
DZ4C/w3qBGoDsjhijNiqz/RzQQFDNVp1zlAtvTyn/1miy7JtsYqw0qGHj3kXgiD0
aifNN4jbF1tgrfx41cBg9MdXqHE7X+e5xKMwMqerRVCSSRnt8yLnlg5NfKn6g7t3
p3hmxIjiwFLBPIeG5DA4yA==
`protect END_PROTECTED
