`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePCFEvFySC3iBMuMD9x57euCXF9r1VQostOqwrKv8A++
sZhOGd+xB5/9FnwOAwwOmU1ysUXKBdpi4wEqQHwNQkX18Ea8tLM0r9NH7MCIdo9w
wMZAAZ4vDCpaCX3SDLCrcl7PBl9g/KXZbf2Ca2aP2qJ695YAmra1udWQrhwutDkP
mnPL9x5qWZ0qWez/nqwps3EvaaWdMt4bSET2LeVEptECTYeIy5xVgjl/SqIgf+46
cK7smJdJuzP0eAnRo3X1Ng==
`protect END_PROTECTED
