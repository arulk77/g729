`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
W/2My2ND0aqTrq9yucSJF+nMjus2Z6SodAGH2La/CNIvZvJWubnDbrMZVLO73hLv
7kG0ZdDptz8gTqGi1RKNRop4XdcOia5h5dxnGGiGwO8gVpELV5MZUIUP7oMYCXcY
XbDw2lobWDbIRrMwazOfHhmjzrSYDozeFY6DNLq3w/bRKTewvPUiA3r7YsfISpYl
DUq1KptXn2xssklM/VcbNzRLpSbjCVQzYsAjsnQekKw=
`protect END_PROTECTED
