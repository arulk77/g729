`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
GDj17RJoBojAXqXV7N+zLAJ7AyG4+hjL9Cg/3Bc1eFck6nQ/mwDeKOs/xkDzITgm
fv1yukqSe896LwB9k9dGovQTfTlnX1TUMgmZbfv4ZbUQpdSeHn5dv0QHbU5OKGlP
rj8CP1tyfURlTKAl9+dppynqtbT0ykPRC5UoUo4W0RU4BEnwRgpUG56nP70CX1xK
1Jvgy1M+2qvOLIBQ2tapcwiLgc44vZJ/rtaYYpFBSHKPtDz/OccEX8MfrcvJf7G4
OzRLvhsELEs0u7Cog51IdVMDe/VuPkUoUhEd0GCbi9xCf1CTyfjV+txF9e6ei9dS
lFIC/mpcbUyZUHQN6nr73j/RJtx4wexDJSg0n7SDWnoj950wZOd58dUuWxQ5FkD9
EEaAGKE/visQHdinnet5bNqgOo0Xn+nU9Eid+YLeSOCG73rALYcloRl74T0FxWpK
IQZCmtc271kV0AgE4FAZgSrvyL9hzUEU+nB/d3ICITQ6XAz+eVzBmvnt+QOpOUay
EwJKt1dtQTgmgz6Lz34PRLPwZIrq6kQ0AAsRq8hvcGcP8iDISGHYcmhTmiauBart
qT1HH4O7m8mc1+cmLVVYN0Shyc27N/B/HgStMr47iUO6UBW3MVzmAV5ogkvU3qoQ
s0V0O/cp+cEQGSPjXSUGuVfrQmL0rcY86szjmK3L9xDxOsMo7XHimrKT/AKCrSmw
+AM/E2DyBHhZg5Bxbd0qgXrq5JLvBS10ncfiiEgFK/1P+0+Os0rpkJ6QG0I83x4o
0CHxBxjmy5dhaOuNsLFu52VanvATEgc4JQSb4dK+y4zymgunyZm0t+swaUse25DV
q6zMsy+3gWE/VMrlw+qQMt7OdQ5UI/LSTF1KA06EdK3Hd5rARZjVw7hmPyzZj1UE
PByg3tlFMzYC/Ko/8YhC84SZ+PFCTEDh3vil41V2ADY6C56XxQs0KsxICE10jvnB
liDcqARJ1YuIyMAUz21Rnjh1msWL6ca/sC6gN1ZFcqOj/L/VrXp/q4ywoiufgj/d
/ol0l1YvDhUHp9cHqqTYlx8bOi3ljRfXQSycFOKoXRImZhEAK/9uitE/6SYXqNze
Ub8bCs6jquJOYofcDyj7DQdRg1lIYZ0Abrpv4p9GOCvLfk3in+N66P15WCdBzOgx
ILeWa7tLQhLkt3HafJuGzisdlfHFlcJxtTne41C1X8s=
`protect END_PROTECTED
