`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN3zfFnIiGDwzN8kmZ+7U+HXGlVOVOQ7uS1rBxKJv0Vvm
`protect END_PROTECTED
