`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
dZy+ShJZLseY/kB72Q2suoeg9vtu6R3sdpDGUqbwxFGvVGCV1To0XhstVbaIXzim
nyvZl1zDoJAh/f/VK5FubYTLjwLQhc+c6NTA18E9wN+qXioqrhFOc9IQLTWp6o8q
T0IcWnXRi+tniSmP5Lozsihze8t910smwP9fC95l5ROUF1aLY5xFkAiHGLpPclVp
osVFzOj+JBQsGs0pqy5AmEMrPRt1z2biS8KYDAhdcn8=
`protect END_PROTECTED
