`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SRXHZlIZxMUrcmY1YS9rmbzL9kYUZjaKSVLt55+z5Kih
8/2LSRf/cCf7/njV+Srvpr+GOaNQB1gPJU41lJvPIRrHT4q6ho8lsXI5izCV5uDc
BJJsTVfxKJR5k/WDfnOH1sFKZObOnljb0Ox3y/knZ90Yj/v7WmtnYfPXwMsS6V6e
1uEPX28huSK6XxpZhLubOSJKsKwAyUwfCpcErYVbYETW3+Z8dE+OWnKjwrUQQJvq
ZDA4fmLeVHLaKuoZVIdHgnJobX524XQfWSgk33BQGIEm/uij3jvrdyKnW/NsACdw
qyIbuJwYL9rLRdT8Ez/vL9Lu6hOF+mZRa9Ytt1mHE0dyXHzfYDPdwtoiMthf1SD3
FQNVpsXCihSeSeyrhQv8US7Aj0+b2pL4z82MCkJQKX/PZeIFvBZqu4o6ffh9rfQd
d7sDsqfXFoDEhMS0fnaDpzQWNNX8RX8SwaRQ37aBzI7eTLLG9543hpKtN2e7etUJ
Y1KWvSGXSCy7nStl2U9RSFVa0P9D4KcZQSoZmGLSgtPhpbsMXmN8WtS0VEDp7rkd
1WTwKP++786W/fV99fd5HzBUrD4po4Bb9mF0UP0I0fqJWT/VcSdD6jwy4i3VpX/H
7/KU8ykbEwrvXpZTPtWJ5f6ZvevmnJBsL/P7KKD4cCi4xqJmRlYYeejAj4nxmWB/
ys6ib6wE9H6HifnTHyH1/O7/za28+oxZ0X/ynUb5OwWZr+hwmEtffsv0VnJ11K8+
t5DyTW/Iq59kNYXrTxGQeC7IgS5Qurm2iwMYlD81riSlkUL1AFzvw13VQZLiNrRA
Zu53fXuva3V36XNH73o1dil9hWEEYZdXzfvVCR1ZUkAZx3a5pWejRgocjxKTTG8I
W/ZHr/xUoks2Hlch48GEzbCMmAhnb1HXKfZEJ4SXMb7ndufPUBS0Lq5lVEO0EgUy
AXk9KSK/y5lglZUtv4rzIi8bG9319RN/L7ovnfBwT8Y+6F4grkuOJBdJfOPOIitb
mar7PDtmXVyNNxoDoHDdaiBKANjeVOzzOIwbvOmbY9Ycx/ziNBCnEIi/3W4rQ/b8
uFS1G4vIVUtw71mSekwL7scQhcPVziPmUywjNhyAt/KwWcqjptSV9bYSUJSEXwxX
/9vPZm0vuB3TILn2aXgMnIyHUZn4CRSvjMFTuFILQSYGJE0fKPXVexCbYxHJn4G+
iHQisWviSRnIJaQuKnRBSRIAZeDZ+pz8pinMITLnLStOBKynxmhdi6x0XOgeZOUS
EdRBqGaatATOK/GoETi+d7bjrX2qbeKPIjv5WgrnKBAyAWCIJB38PIhLxswbrjgH
Twhstu9Way73L0E6FOoHL0BWHl8Vt4FcckWvX8i1aj5q0H4m4q9r0wQ2d0e2fMkS
vIL4hshRNhKTjjSUSOM3DQOS6er1h8jhdT8z/Lu9Mt97MjTup2qzh6zTVAvxWwlg
DSj9qfr64GpDevk7nsNjMVXqMbLQNexU5MuW9N6iPhMSJaUTi6BZK55XDXG19MO9
fowJJoH8XPgzSKClRHF61/SzNTOV2Nd13pn1ymeuYij302AtlOlqqcKcGRJnu6FZ
aFUdvGsE634ZuxXTZ/z5K3cj/oKhaiO+je7SXeZ1HVWuLVjz2AG+uwUo1y3CYYD2
C/zJ6QR7o+nhyTVI6IwQAUL7ypcFbE0Don+xGdpPTMgrf9SlKqqHQg8dpoaCCLlN
ugi9mcxZtxZrxJiJibxieKPFXxXEY/xCpK2En3lDli9A8zN1EG7X70dcH8f5HYRZ
0ulsoKUUAu2FpIuZ9SsrGiYYMfbsI+/U31MG3s9spgfxw06jR+n+tdSH2b6GZVgC
eUBRLhN2f2apU9nUEqFVVz2e2SNJCd/o8uyCWkQm8EVFzO8wVWFdJnXHXQk2q+U/
urg+hCQ5nM57ldNAynFyzwrkTrpWy5c42M7HJv5PWjEHtGKJTHoUv/trnJiJzw8b
AMd33q61IqYZ0Zb52Om4xMK1/h03foUn101O9DTS+6CpWumg6fRKRdUyjMh09Y5t
2T6TMsRdF3UT1Y7PTMAqfAIslSljtXQ/HU0XZDZixIJMYRbA0CaCoLWyzqvEODzT
hha4N94VFO9aG4xOlzdoqdg0XDoDkZdzHayqfW6cq1sFFWrExdHDjYh0gu50L+8C
+Wwzsn8hPy60LO8/197sZp8i04QV3w5ZL9EmoicrdhRFfLRdd+16qb5fk11ol7Z5
Eh3fVn0qc1F9+2sN0KxAvR3CnuRltwHhuNINXhXhWcoZNYdrWKMdSnoR1j7ViJ9T
coZD3Hf+8RJqQ7bnjiMGgsfrKSokje00Mrtl8naQFJGF+xcZxfQuYrSCgzUVy89W
tktSsstA5Ux7E9/DvF2iTdhSoJBtHLWnJDtgIsskVBvCoc4emFeNl64PvN355eVA
lQuCf5Q8TEm8ZJOp1WDLyQDiFTjIK102PvudcKbaYQpn02fAgVuuqlCCUXZ6M5Zj
KPE/qHjUsuh/HXQDsprUIzg03kZZQ9BPI2TG8PHrvpkrq/G4Rk6280MSCpYAgMlK
qa18SJH0WUnlKtIwPBAhwVUJxyGFBOQXQSrYjpdsWXJ/rkOlhAPMB22xG44vPMoF
1nQQQ+MXk/Nd0U4NdVAORwSJ9EghC+A12MHQtVqJ5xBc9kzpzevZ/5S7iBA26A0s
vHmEk0cMW8Trs62IrJRmLP9ZYnms7TP6+X8u3FxrpiZg71rJXuilElP8wxj9s17U
RTruQ2MEm5wDLx09ngivnFlFY6sfjjHs+ioGaPIof1EUh20mWutdSWmTKoaD0/tg
Ob7k8I/mriqMV4s5XMxAQ7oVBUq3on1UcnXdENNP29jhL6kbNJ4vV5KhZCfhwVMg
ViEqfFEiS2ve0vbJLZSyLVzyFIdml/kirH6ecVXFROd4kjJ2vjD8uDcekYNcIgRE
`protect END_PROTECTED
