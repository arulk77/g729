`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
EgjeWzNT66dNouyGH0l7cDQRoCYsxUlIBsscedh5QPaGQ+v6q5L6OqZYREbozmL5
E3nC1EmfoC0kiR8ZQTly44etFjM3nGrkMYLVABQbnjbugdD7siVV1heSCWJ7huEo
uXdnt6kytMV6nJ3hVyIHkpGccnyC0HGZQ954IQJwvHyX88+GQCCgTvZyuuPOcUw/
`protect END_PROTECTED
