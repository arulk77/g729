`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
1sEQtvj8m2vMaJfS3BzRom0fcEcc5JDbJhD4dYQJwhWonqUhXCVK59FVSkdiG4gv
6/BVlK/jkvhSB6xz4H7xWaKv9mJV67lPc7x5nHaQsWBOq/kj2qx3jQ4a4OKtE+6a
kiEc0izM47SpG+gDI9v641UmMO28Ine8S1uXClBj/ZHJinW7wxZFwO1kjxUyX1xh
gYyMDytV4Cen9zD2+aql7aZ3To258Ne+9nUPLTx1zdX8P0uuGToYUs/gcaWktb7I
ZJA98lm8ZF4E/IILYN2hKligP00eC0DBnxhdLa5vEk325KfjDbzEnB3P2LXcodfD
7Q8+PjJTRnrQw0V21nzBCreQOjxtcEepyWgxCDcvwpvA6Deee2pxD24nUOyUH52c
i+vC20VcNz2VFOHSQXDvLOTe0i+f//tdOJ1S1HxCycZ5NQmgQnLdE4l+MJiSsaYX
pkKdWOLOxz9bD/EEVuFUdYb7ncvUJTKk9UGS1Nl/ONp1pF2ASuhVJE2lnPYnzzrg
F1wsQGstkzmgx6e5u0oLM5mbnoucQOrzLMknU/uzHX+c7NGSeqmwLGCPi5WPgQOM
N8wwDOBcF+UcA6MSS08ww8wd9rThKi9kwBwiDsYUpfiUBm0o9G2pr3bW/Zt1N9xW
L3xHtn8K18f3Ptab/Y5NATijYMalC5+9GYy0Wh5GnL76XaeVk5LkMf1ybjKV1wSK
zpDUUduwBhvw/Kr0hKqJEUR/BaLsfH1Qi54EHZzEeE9nhK+ZhIfF0xpv0JDveQ2+
Le4imyE67k7rUCJ722/nRiIVmOIBipvsIuTY34FekAXEeFazANqFp6y4rlmqsRMl
DITw5F4BCHkLmfgTMxXvSPWCailHCb+QQ/5//e8IkdBlnkRrsrldR0ZhsmJuylmJ
QYcukV68WUHth/Jl9GEFpk+wj6iUPBsW2OxVbRQN0YkI0Q/BZvtsQZ349hN91iuI
UvZoqiRJ4p32BRGmVG/5mrVTPcwDsKeECA0Dmn2JLvf+TlrY7406GU2ZET8XdDC7
piEgQx+l871t5BunznKx46P7ZbCFBPd6OWR23eehjzxbubDpbVh2qNGFz4CJy0Fz
rWRZi4lBrqiFQRJlhaQO+yew2qs7TdaQtKkDYC6cW3yY7jEjTA0fLX/mmS9YGwl/
Uxr1KGtwwXgFA/nK2RiYLVZ7VmA2WMxPvi/KbiOWfSTwXXQoJgLW/3M+X2P4pjsN
zgUqeBlau3MmSlNHGhXi5L2FrViKLhcncpttxeoRnRCmpBftB8qxBpoMQzRi3tk7
pdYLEHeAe10Hq1mUqzQ2gtF119nAuSVEdRlo+5Mg7jVKr4O+WXDbK2LKPAmd1Jqa
z/Y2b8i2xwG/z62MoXVkyehE/gXFd4MFhqQcMogScDihiLPbff9Ny+JlBDJJq1Ky
u8gVj2sOgFMdwcOOwiNYrY7s1WL/FPg68A/IWEC9oI+4AOoH6ESWn8QunGX+671P
DYPiXO4WM8eFntW2iKMF7Pn/vzypK3JC/AkKjCk6sdyBRiEHhocXHMQGfUaAMsyB
OR61h8KJYP6p2CH+VQMNHhQLvpVU5qK/beWLC8QfMcD9D72IUWDpZKsZkcMXNc02
V9ogRHi3D8YMWoNToTsWO5Yhpi5g6LrsHgBceF7G7FiN1/1V8Z63/1B2ijCfIXr6
Kcfvsm5Nsq2DhT4EBlFZ+Rh+ORhetrzdz4cphOhZUxDmmSygVHDsK43cyAkYd52E
pAstQMrUql/LIXgl+pRwULHqOqNjd4XVvXblPErugqDxvJBlY6JC5RsC8QUF2Weo
rqT7jK3DwVjNXJgbKrA2QhBMBNsiHjkpbfvbVzLKnWdXZyGoHNJ4bkZwEzgLQH0R
yFJ+W0qYzZnefYyWzM9Io0WAEbrJ8xs0AfLv6Gfsen/eTNu8oRgDENZC9iq+O74n
JCNUKCr29ZgK0yZPCJ0DG1YS4ThDECb+bHN/aaOjjwnVCZpjVjd/GQi/rtvbLb6P
SDzDyZ+pzbEGtELBeL/AOPA+bJs9wsGR2ZuFtHjDeevlP8+r8inENcLTaRH1bbfx
YAPrbODODO49AvktWIeyNmcXNJkv24fv5I9/4oGIZ/2FhS08eak++/gd8JGeXthG
OwA+bX9RJk0qK/AROIKSzIeIbE9bJobThKKTBdWnmahLi2j238ncrVIE0Gj6U6PE
zDFdm6d6WPB0Df5Jon8WG4Kaq/XSa2gDQWr6ZDk5rJksSUj2fKFXO8nmw3vlj1w2
6eGS1ZA+gkW0SkOjg3PMD8v3hSBs/GyRoubmpPqyiILZ/J9VAJPHLsO+IYQv+DoZ
3P7MmO8UnwNbDvd822tWKc8B0qgGkf9La6j4UcPV/0qqZYfrwHLXpp7y9nD/uBl2
WnazmMgoLfVu4OZgoPg5VjRfZqsdAGBdC6rofD7z/dKyI/TwhH/fS7KDZFaV7o+J
BVsrGGNe+3IAifnfyQG46wAxJp55TAfIqYL3UNd0dGVcqprG44BTXd9EA53NWzNi
JCwLSzYC3QX+B8hgiu/wF7+/KY1mzgugf9bu7NOip8Dlfu1p0wR6w5szp9FiVXHO
PLhtIQ2VPK76AFrrmyJ4K2H3XJENRO23ktoZBjKn+hrXPo+GBh10HMZfn+3xLkiu
c75IEG/vsxFs+09SH5tn8IrQGtOg8mNJLgP4vf21YD7YHBu7j/TW40rpz4pvZFYj
gAjjEs8ZmJAt26bD1FOgF6CQSMuGyGnerVctnDE2CpzbaxZmerF+N9SWw2xTwMgt
QHN8BNT2kJri2LvkSoVNBfp7FXvA8HOT9mxe0CKXal9Vmd/YqDHx09/GRkr3Qhsn
eFrmPLUG1P0/w4X2Ca/5iXQnP+oBKigcBIy8N3TwzQFMJTCVEx/0fqq/j2NckLvz
YhBxHCTbidOx3ZNUnpYGsHQsTwnDqIvODNLQWxpfNeccUR+oa3BXvT0M5KJ+msf3
xSbSXbcDWRa2vBpbzCoAqbNeHbHEm6MseD7HkYBzISRc5a9VYCWtLyvGBVJlWCHv
pVHnudBopcxOk2ZrAXbHC6LteIEUYxcn34OYzdkxd/ExjhJDzzcEKA5Bz+zAZewf
9tA2dT60lYttmF3f841guw+wKfIM5Tri0JaW5H2RyRy913l3J8zJ7qlwoQwX4xiQ
AfYFd5BJ5nwcGelx0jrsR55hNqwLpS+8YmFN1oziXU/yEMa8ioLPLyzKzgEvH3zB
MdNnL99oNp9ccnq5mCzxXC0jdubTZ2ijDsrbrCw01jsXXYmKnQ0gb2fZ3Mp5pPbG
sdzSsEv5UjLAa+7cEEcKxRKblhHfa3VLO/u32l61R4Mk6qetvmI3Si+RPNQF1pu1
/13hB9D6RRZUPagTxljjsLJmvVWpXC2RFqFphaqFijfDWZ3fzd0rv3dFxU1ne7W9
sLz3mne0VxFKZguvZglM1IJBJvR+jWoZV9RgNTVciNp0ehCluuLY+JiGdWfnYdYx
wbZRQVWafQ9K3mTEP+3hUB6PLnP8UPYeCiKeyPgnfpTJQrMNb9szuMeLLIoXkGEh
K50IfbEWAz7AR7i1oob0jBMkhfBRayCUTIAa9wgl6YY9B/D0/psY2WoMadtvmmdG
a9xk7txVs1+4Oj1gUpZqsBdOIxBJkhnnjw+XWYYAzvYW/tvQDsZsfIKXQNmi2eVC
OPPYD/PPJPXQXae9HKqTpuEVKxPFwZ+7y/BQgFOrBf0z+UNsi7Z9ky7vFTKVu4vv
q82+e/9QjrzAVDb45UqwMV+Jt1ZXdGLGngRTrfsWCSobmmact+mPWsvAYz+WiyjF
ELP+her0lcZ+bq4QVn0wVSgqpnpmuuxGB3cbi6b52sSXTZ8eLVxxkcZTbxIPA68c
/0s30nndAp3JVCHFah8X/CzKvP9stXtBsv+sYAfMz4UWYnQMrq57nwy6fNqc8uIo
aqj70jrgoyNnDVOtncHJ6ZLSU5tnoV9ChE2lbmUX1hXO16sdn7874pKpWxxGdEmA
xAtKgd1Lojh7ncjFETEPDbhqiZYzODr4WD/D7KXp/l6M7lCRc6tlHm/Ab0YPkyUE
JVuJbXcnYa9Kqw9HOUJV1Fg7G2uEJ4iwDgfgoyFXxlE8Of2vvzEbE/XgQ0xKO37h
Wyqz0yMTTANdvDDm/Wa9RZ5QRmzp/TWK+LJSIYEBofgQ3XQMgsS7ECACXdsmz+b9
tQnL2NApyK9acyfHyu0C7g4b+Md/zP9q88Qy3Zk0KRWJrbW2D8/5rBe1Of1sdEmE
q5g7laAC67Ln84dxRFNER34qDfP4G1pzbVVxlFCyL4uS3ig/cwQCFgNhn3/zJF0s
FprG6k+3qpzc1+mU1sAuTe9mDvZMlPFQ3E6h+s/y275/esBdsH4ZxwU2p7Pe6lzj
dy2yu5g+alM4plkB9MtCTdMelUQW5C0TCTXmhbr7KesNskTtKCNFcxr7qhpZqm1q
mRctxvmUngWDNxAXXI4BRiCakzm0SlMLNgN7KIXEOcEmjjP6/QdQJeY/mqJcIe2z
eE8JRh1szq/tjmU1tWr7woMk8xBikAsIevrvRZNyVpllBmUy5OrYueoPWGZoEKiA
UXWscuV/KxXdZPgEkHgOkEYLEFbdzljrmgQgASipwHHSxJBzjXoSvO7HYimJtTPg
AwGLz5WVINg9ivrnEYD+EHDK2Ll5YI4+8Q9VwnYKXG+3EAMM8ANgG5WFchbFnVJf
hF9OnQMSC3VoDhl6INXICDkaWUHACLC861lZ4uKTamm5rT5YH9uhxuXqpyXYW8Ci
ZCfHyXYOqpB0VOopQu7d0Ds3kpmxPn6Ve0GwqIvBz0lD7w30fYSAZSfwEyWOFQsf
wbp6IpP2f38mko40eVfMymd7bg5kUxpfPteKMgl+P5AGgVtigichPuOm4a/B0MBd
QmKE0mWGwfZybDRcOg0pvDokzTZyLAOIxSUPyXYhKF/CUfq0Yb/Onkz5+ftnCOc6
nStwXQAHqj/6TG1WMY3jCjINfaBHjvCXV7uNd4NcVpCRjRTDNiAE+xE8uS9Te8i3
Y0wSqFJhduTq2EtOxaRt7JErzLESQwcSiDfg/DF//W1muPlgkZqVurkW5niz7usE
KN0dsqFsl1LE8GH1j/d2+A==
`protect END_PROTECTED
