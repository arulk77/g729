`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF1K8V9gl+QLDfxWYfXHENpfq6eXf/1PveKP1GpNcDIH
kkS1eNZs5WGIp9X95ONb3bMtGGQyq6TUR2p+Yv/59ORnMdrQQCXVGCbeIYdsPupg
04jRj0xZPBgaCGWPxH2k1F2iF2v1bA9pXopuZbF8ncA1pnj5hng2vczJOeMrD4YK
HzqEBH1/gfXO5No+6P4aG+0yURCgPswnPt7CPVGd1K6IoDE3YuNX5M+Li0H5Mu/A
qw8gasFs9n9DF57J2klK+ew9RIoASxIv/nZHjdCd41hBdeKGtYNW0/+U1wr2q2s6
SYxSocg54U4SIRsRbL9jIyfvUrjj3SMloGa6cNtRvzVFJS1WGxxszzgpdSXnJ97j
kH7cY989v/3hbvnoWxXQoqBuxHem3xpfsTZNY8rlY9SVoYgwtSf9Gf6d3+r3yzGg
s9OzrxTL0FMV7nKaIpClYgAScMWD64CDMOcHBn/7wF2Dmzi7iWQQ1CKZ1gKojC9p
`protect END_PROTECTED
