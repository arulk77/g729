`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveITvwy/a8ODMS4mOAVsA0eAYdYGQyKLeOZ8zRMfbcsau
7ds/om3OWdWpTLAgYOWAK0mWq2z4UTVUqeyZHNfZl3ZFrjd8kUsFJKEnf/HxJKFS
UN127NuveUOovVvIh6VCjypzjLUq5CDdL1extY7qZtwgm0OEDjsEXRvtIOEnzeu6
ODMiyQU7FsdQ8lZkfBjoXw==
`protect END_PROTECTED
