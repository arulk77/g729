`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKeUc39TqcYUZzedDtUEHWG3sWaXCuosOmxkhYfqT36b
u7j1YRIV9QrqlMZxQ1VtZnW3/LekR8+dot5FTH9WrAKKtU18hRBdsyYJWUrajiRB
wq4xxx3zTKSuyVCtaJu9Wc3oDSVvLdHnEqEorstticETFRU11HI3vLrbZb/pFBUE
rqusGKi2nJUkQBHs4Nq5QKVv4Ugh7TeGmvaWjcul209cAXto2FOYOaJRUpec5xwN
oJKdXxVEJkRk0UeafqOBnqVqJo4ujWheAz+8dGu2WHnzPSx+BKNYypdvM8PlR2WA
1Q9wLK2mQEB/aF7KLrTD9MW88e8jq5BbI3yixNbu9/KCPKeCpgfWTj56no9TFIK8
8I88lum/jxf/+twyS89URcgbyLCoFm5xum3FdnarQ8g=
`protect END_PROTECTED
