`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aXvb5QpSnZA5XkXUBQVjPVYZdalSp1hpOA79lAJ8zen8
b3PFAIvHuNbxATrQSKr+dRB/gihFQCqQPg0tJw1ujcj7Ghl6xac8LCva/ttfs9Ss
syfEg5+mTEipS/quvF5NdiNbRQ5T4ozCCLsIwVNBnDKySUldprt4+2eVeiPHf3D0
ErYjbXHVRzUGuOH/kpbvml7RZ9fthA+qAs1RqYV8DpRGq59RFBo4xNl45rvA5/QL
bayK9AgDfasWlPlttzqZn1nI4WJgn8fC7htsD16ZNT74g19YkzxQPIUVYX2g90Wu
8h+Q72YTY3uEzRHE/9hjt7F5QeEau4tX8Jaq8ZESg+Dad+1tzjF9XAhUjxMHurQQ
oVeds4AX4qsFqLkvxsFBbyjQFFNKIyrXKdXJGwG+HC4CfkPug23nX8jWF7x0zaNz
dnIopCq5P1XV341aBZpGJOTMIzgZymoK61kFc3Uov6cuiB6Ncz3XLwSDpdpU7D1p
D+AYd9w9uy7dQvG2cAvXKeutXv30CZMNsU56JwTtoalsbT6Da/gtUy+umPsrUIwA
hO7ikMmEpYhuxpPqHGylznzAgjqLvIgstiQc0Ace9rTlzCEai7/+CUxp4RtRDm5J
ldJ4luPqqerLfKCdEhLSqvSSO9nKJRrU06ByWotZ1JiY6anJkS/UtcKhe7q6tPbO
X37khfk3nbc2DwuBDOHLyzQo7F/mW7WnOMPEdru2BFiCmCn0KIxWzu7D4D/mJrXx
EjGIwtEHVxVsCBs/OljjNnsxT14B5nejvgB7+uwT848VredIyKyrpyyCj7nCxDTg
lAkdLZ485oMgqjJ1XLd4XLOVNBvOU+yl38TYIFu8KoGgalqCwojOCEuE3y67Y6NR
MduY+blPkL7ybbN8ok3CGgBMQzqtPlR9CcLKDVx5bV7L2IXfQPh0k+3n+xPMmue2
7fhOw4FCsJQfeQ3BDVAQnU2bXMeUgekwWJai57heSFPOVh+Dznc+xgeV9qKy7NQm
y1vLsuiDE4a0Sd+S7GcfLNomM0LQLCcn+YvUsZa8pU0KdCoMjjVLvMe8x+fPQd4B
lS8RYSAOphouD98ODm7/ejcjn0gipk6mrsUFd46A2z55yiPlM0XzqUgaZdnUJ7RL
G+PxxTf7LDyvA/ac4m2uSyZ/RJ3gR1pVl0XxQ3cxRh6K2XuxxSi+FYNpwgp0X9nN
d8kq38J0zPL8jBvQuot5hQ2Id4Lfo11Vr+IRuN4EOr5swxnf5KMDGzZMY2K57Vju
fbGDxbQ7llwVrrHvlI9qN7FrfJFhL744bzGDhTlUDWkxHmAdqpOPtC2x/RaQLH+Z
VYL+bWErOnaqZuQy96XNnos9qeHpjP3t6ZhXD7w2fwb5D8+Jmp2JPsVP/OsEruk1
Vp1Z+jBtzrMB9Wok426DApMoeOQesqKZT18WaZO+KSepInG5GZd5HIo2slcLEuBW
3BuHleput05jwJ7TxzUwjVP9o/jv5sFcDvhj4c9uXdfy8QsFfHgJGG/0SfpKzW2i
o2VSvPyv5kfRLgnwjiCfi9onRWKnVI+KP1J5Y4adayetgKE+VoMwel3A47nIgyTr
1yEnd9UXjqlHg4PDmG8D3RKS0qyoOELFYPbqxcI7c4o3a47QDi2d5WkfM8soL26T
E/AOp9izH1g6Dyo30zxthDbKT4eXQgwVx8Eifp9yGT4CZt8nIfmM+kJQRU/hDJBR
9dtY4J2fWQiukIf59mlP/95p8T9quFs/k6sXavDdCs7Xa8khAMLtcNy2llr2qaDE
21LKMZ6E0Wi7UDVp/yzr462tXmSSCv63r+Uy7gX84GUGlibkviUFkJ5y4sP5Jyos
A+reAR+K84m4unE0fAoPeK0NxCEMHW1+c6fA8Tt7lMBe1JcBZByTUDMIhiqLkRJv
2Vm+Gx3g4hEs1sZVpGEVigOnOjRJhMbnDdZYHjyKWHOY4GlU8DdIBN+Ff7huaKA+
HjT5nVRAx7X22ESPcrtq+oy+GSR+EbW6XlmwHfzAEkaVWzbEGmxslv+1rUj/V1U7
r82LkQnjHE5yfiZv1RrfwDvy5yrkRwDu/O35CorrXLS6EcyKCsj8B5NKHhHcGmq3
kaCSJ/OxRyzg/bNW9f5/65rZyq+YBOxm1O7dNj4YXtQGLRuO34z2Pruvb2UsYXXt
kSSDl6xtGo9jIiHo+LweoHCIEv7p7Mklfc4FYF9kCmh89ze2gAuz0PdBGGQavf3B
NuMmexpKD/8yQAPcoYyIW6ns4bzJNUh6brHeh10SjtKAoFixkbE9bhVRy3mN4boz
Xc7EmNdfG8f1fFP28gTlbba+BFQUZoU+AV+1C7ai9NALs/T243LbY4FbREf1+X06
cvj6M6CU9hzA7n6ZFObxxLVTabm+J+ennBSO6wt7w4ojjIM8L6ggRk8xjeeEWmmY
UgegJLKtmRldO3d+Wuhdv6/5j9cXIcs6OK7SIo959f1qaVWwafcNaCF1s52k0Dme
nuy1TbcoHtGe7fkvkRkHdQaJoAwbgNj6GNI/NCpRCtwka2fM1POwFfQNF2LrpcIf
fh02twZWp8xYZ7OC0nSJ0Ikd4g8pQydulI0su5RQIiM2FuIYqR22I1xiTvCRnGFi
CIFBWFysth3Y0gCDAuKOtOyBKHIDaClKwcVIK9UzFFYEzdVYYNIAwh5LxhF7J7+1
0aDbr+s1ZYYeKFVUIbUoqc8HCYbWeDtPJkqHFOBVaGzirMQyIuHfx3hqGzidG9Wv
x9iTPocXSJFQToWmchuMSumXJ+lvVOAfCPGKHNIp1HaFiU9Xim5ni+TIBmw0U1Yl
UDADBUDEV2IZPI7mq7yo0xdNhn/5XrMRMTwaE6fr7k9PlCXOvf/Nvb3ipB24Bdgo
giQw7BWw9Sbg8fwUokcA6YBuaIXb/CcKzwsM8iyH0MxuREIie/zw0ub+YkWcaUzm
J4Lub0gzZownURN8bWnbsiC9Qb6kbFPOi6EZI290Q/l2SaaPbnvCzgBKybWS1+r6
sVvaF7vjQ8g2DYhTKXzh2k4hkKxuuqQERZpLRsrZapzjzOS51Aq4M1VBFnv/cpkb
50VJggmG35/pDT2dsVnRDZWrDRT7xdgVbi7Vl0InCHuPOOlfaVLVYPZ93F3bvrh4
M7XLmLqUgtvCpTIgsgwU1pPSJyU7On+ximOH8s1LYIXsFqm48U9bYryq6FjiiX41
oZvuXzY/m66z3C3r5Z0LrWeZE3bDwK5z/SpEVqQmYh9UY9CIBnGrUvkyMxEC8G/b
0Ne1A2LxEr25FllpkRp9eGfVWoR2vyUyWMcnCfKFAonPgXJ2kMwl8vLPddYR1JIE
4JQE3iitb/ExYr9jbREyrKK5QxzBL23bj0IQvOzOJ0rUubgBupK2PhpXwKPEJsQw
AFgVFk0H8Sylr7Obdn5xCaq/NEkNXey/U4Sqluq133JGy2N9C2/LzM+47DEQv84V
I+EO1r4Y7UeINgbxIkQF9thryvwdzPkuBEdOS1czcU2AeCFxIojoDxKume2hrQj7
52UOf7aQ85dQTBGkHyLM/yopOn5vzx9qDAWXJ+nX+RM6ummsW/E4fHP0LnHIXvDU
17n9Smt+ZO3egFvpoMZUadd8YmmYJ8wr34c36M04cFojPEIt8tGauR7qk3rx/AuP
gC0qQ27LxVnWcz3aw8FkhCcfwqDG5nCay0QjPsk3Gf1y4WobEDGJQCPtUXMF8bxv
RgLnAebI7b/UkXiZBh3pL1riz8RC0Iapd1DbkoBzs66DLhGXMezV2clVw6PB8Qv6
NKC/oHW774F/0QKL3Cxac4zY9WUnD2283J4v50EsVRvNsMIeUTHyVf3JeT8oPsC0
FSuQYTAcFKpuYezU9Qpg0l/363f6CzwmI2ix/MCXyo2TGgg9IY8i8KzTcQuLEjNp
bJVhsOQzI46Gol5t/H9rIXJRyWUobThwsaXX6iV96k+O4dZgHgDZnQZTx4nLXbjX
IoNxLpNqtqCS2XOH9NswHAvwdN7FAMwH8i+165czihvXEFNWWiYko5Vs5xArv5EO
da2GCRDk0rn32pe1MUvjsQYqXo5XhwbMjyKj1oOO1ZDPE3InSXRbA3t0IkEC62/E
iE8h2H1Idj9K2Z3T/0QavN/DxDU/4ZiR4PGMb43t77iu1NveaE828suxaDawOm8Y
b7TY1QwE/68HcjSgBEmKvfyL6da2PQYEdTxy5Q7fweBOp79udCI3xpTALzb/ySKs
Yum8Zfbnm+WufAx6GDOVi0d0tO/2xrX3/bj3iRbAscaMe3Nk9yqUdVRPjYA4xyfr
UJgvAi84djEHAv+rAY6vCZ/mIBGrVS1CMiHpISENJZUQsXpgr8l9VMnb5MMTtKZd
XDI97yh1Oef+W2su7LqLeICmlJ3gSJ/GzObZfQ/h8hpwoSWclEH0zBGWERppM+ga
Co6hmMKyvpLI5y7RNFRT/nyZTEVmC7ZCiHZF3xDuDJZK+WnQXWLv9VsHtNpSXTrC
SlhztuK7tZ5y7ZDuOM8pdZqneXfJskUwGlgbGVwYihomo79uQZSASpGB/i7rcFM6
7moV+jEp2hmk5rcVXoQ0Dt+7W9seWYRtOpvqlThNsH/JpeNRw4cd5AoKbBDDBvzX
/yi4cIwyx5irizB6p17Hp9x59eh/sXkbL0JCP9llq7nKnyf03ugsTJp1RAJGqH0e
i7lm0yKJBK6osJtACOG/EZDvHPGLS66w5ZOrzX/53XQfoWtbnz8EmKX3UFEh9OL/
IbM4QIMLwShzHqaDzoQwXei/4UCR5Gi7fdgOjfytuiiAV6f4XNQSxyn0CWbS2BJS
tWQ5aVJ+jz31FHESaoi0KiAULKlWVQroIlhkT12Sof3dQO0Gmv6Si130SxkSZIg3
kQSn1ANz31W9ZAW63CLPybAxZercxqWkyGJjn3+Jj+uqaD1cu2n1gsdZKia8Rg9C
4QeT24O6SOWqDGFVLjhHWP3S+lUkPB9iS3rI9SoYFyL6n91GdY/GZiYj/xvzC1lA
5kS7cw90N5FS/60Yvb8gYgaImTzpVETQ0IfvNOyfnJqFKMpPIsM1GS6qXwmdvhJy
gJHRdTgyqhOMTcLivx3koc80NhJiCe2qSEQRahJmgqBFmLVrcD2M+fQUnSqnSIRj
szsh/Uow5qT2uL8DtMhJj0TjpqLCTLYdqs8lYCtFHn9/bl+KZkQeeKrjs2x5VThn
I3SmLrxKMZTjH3jZATjz+1+tlgE0olu11y4+uH4b1GdrA1mRQge5ozPOh0aQgozG
X3rljwkLBpQGGNNoeFjrsTJ3tlQPI9AE9O0ZJb+PcPfldoILEIoGrqpBvFM1qSfE
pVIaokWgnM7ZbT2h6g2aie1hL8S6YDDb8FJmMYgffeCF8fjL+2htYItdpBqWPSE6
KX1lSBU8x8tMdAEmae2vWZV5pcvzMwESI0ife8hdooHWljslBSharPw+ZuEF3zH6
gYEEdfEsITamkN5HhCl/AqCfOsD+X7FcnbutTsI4aSvXgJ/rA7vd8ah2TwJsnmvy
o/2ilwGpYDquFvd74rF/PJXG3ka+J5fB4iUkIIEywE/0ZL9Q2UHhQ4/7oV6iWR6V
P1YomFzLn6KtObyKhUDrs1QNGYwLiyTX3Wr6uKYbnyLwQ9OSpEVYBQhyzezQWv4E
QAtXYYOnUSYQFCxRyCQL62kGW/z4YvySA3EaQR/8A5xtlewc+qED7RGaJ3oCbgaj
nV6yPV4cSAYOXSyKu8gSCCOW1fymPt/90O8xLHvBOIhiG1dPOphjpm/clOm/JY8i
cOg6A1zVI1Bt2EMqzYi0F/Qkjb2KoWsl2bwinvBBcEgWKD10SISyZ4tCIz1uh84O
yVscAvOMoh9PnEf+9JPIxfJwXwEcwAP06uszH94vyg9XRY4cPH2vpKBd1+7oClWA
CzkmaBv/n2N2XQbbK61KoPMagdP/BAx4NW2rO0KMjSVaHKiz50fzYASstl6FclW/
2pihWHG+Iz6Qn9iprdam0XKX4tjZe4LFIzS4qRzd+NigOiU2QzaRy7vluakoycHN
zEJqeqbKCeKeQxrfuLICGZDOQlkW6hUMEp6P3GV3XS7+ZUBarhuzaGxfYrrAsEvM
Ahd+Nuoo3oVG17UAwk6t8wBK7ivtLVQMqu0dPXQNcjWuv2+PjH3JfUoOqz04lozP
vHIadZW41G4q+2Jl41nBLMrl8MMmwxs21DcrjlIasIMzSS9Eep0kw+H4k8D+NSBQ
o+n5xq70wkm+c+qhWSrka/2a4ajeCYJgfuUrm8PIpmMYPsexzJO6W0C+2xnpCkld
/gn/fTQU56gcte6sOuZaoL55wcdJxu7zCUQMkpzNNdunPvVV2FXDJlOcRSv13p/N
RlIeIMPQclaxZ2dK5fwI+x0QIJ78SWzs826qOR65rRVw6lHetr+XyT9ldSDPYBAw
B8sBjoc0lUTuSslC/LO1d68N2/5QNwVxoTKHJ1lzG/X9sNHpIr/X/73zk9zZC1ER
VhxSjRh/mq+3BPoOfEapejcP+afiNiCbXaZ95z8byYvi5IRjcvU+E9CHuqroXMoF
g4AV1HEz2kh8uy3KHzw1VEpllqQwwUXwM0RxwW0u0NXn3oFfhpPdAVD3AH7BMiSH
NF/B2xCcvp7WZyUTov6GKn51Dpbvq0drtsOdPo4p7/DMAxry2yD++qKaxhEnAzXU
Dm3PMh4/FmB/fT551dGpDacQKidgagyHUyiPdhbId49BKyJPF1SwzHu04VFbSwAD
won6al7GBFSTLJB951iSXI2BNsejL1nDkFqWFXDZTWbss7GzIOmGxRaqYOGGnvWa
/LyetRzYWr60roeWSc+H4FsBdO9F7qpmdwpAPPOsiaO+5V24B+PxGD95JIEWbZBB
vkDI03Qd2CsgBQMODQ+tBfGOPVkwzRoRqOvB+flLJnpM095NKskVHTRKSp4t6lUD
x0uxgjpsMI37CXVWkXhzUNXJ/meft4KyppDgk76OZJBNYfVq6L4wGQrBmt/VY1F9
g3GbWfIuH3coTPzVl06kT4BNKi9ObugLk9QZv2sFpbt61LZlo+p3JuRUxE5JEJRE
tcGHbUCE2qDBy0FTlsVAkPWZOmfeWORWjy/Pt5ovjXcVKhxkLfg8di2X9z/dKbwa
90weKffCrtHwpGnTaZtnc5DmQ19ffVnv3D9Zj12SujTFWGbrPxaEiOwg2foX/PhH
fV543UBIkvEH7t4w2PWe4Euohb+ctaLisTMuGcHHiNxzK0JWfsZuzefvsvGVQ2BV
Kxx5v7pW2H3JLNVjFcXJW5mCYcSGkoIk2tfDCf4gORFQwnXg8Yy7mBrMfcMl4jYe
2C3l0DJjyR9V9w92fmTH3YNzhJrnrvXO8U4LF6Q0fiajmu3C1WmN4Rlie/Qu++CK
GDyxmdZCFCoWWUuZbDjhJY8TZidH69WMyvjKufh6BdydU+DQ+WZbRMrJI5TVVCZU
8F5gk/Fw16CKXBwVGXLNjEjRJ6yFuXbLBVwaEG66aa6vs213jPW9Wa2/BzQhB7gc
oQZR4KzvHERdnpdZybdhLqHjNCzw7Z+juxtOYTa9uOLt6Ce2F117UDkHIYuxBmJN
0cUpPquzGYPL2shkXmPgokM/MGSCLdG8/yHj2a/gVhpx2prgzg8iMzY9sOoOATkg
yQM5A4edbaXXcSLBNyryHJwkSAcr0L2F/JJ/7hJqYeXNZqvvRJZcjePZJ6X13iDf
A5tssUeXAVysHUp9tCpKJctoPUbJXcY1BWbylKW5XFVRSFJ7wT2gxWriyq4WusW8
eqSkTlwBmQguBtyR8lDmv2mf893E/WSFI265JPKt8CLVr+D02Plo1X7Bw1ExTOpV
JVSwaoZGADoSWViOyLRNxCO6l5oYPC1vMYvVoWz/qXFdqBY6ALlxvH2MLEfhF3TA
czHjCYPbScuhvcg/DPRaB2fK6XZFPfdLWoBbFnqkFCe9zY56rMKA+Sa6Q69VFOQB
FO4hrJfMnu4TtchsOqUBvzU1vw5CKQqcqmzSvD79ovm2U5E7PeaEvR35J17iN2bA
K6kEKuIIr6rMUduOJm/2UCMVOvYj3qsetKO+WZEIFDoh77La3DHymUZVxxfHzDE3
3TOuwPCShBplj0tK1wCyHhFd08bIaONLYAPK6JdspsZuRZvTkhus8/6FgtVrT089
Q2ubL6sAb02ciRKM5hUiwGRKe3t0vTNG+UDMR0bz3w/JYJWJuFcQMHJsxCcQXykI
IMstHlvCafjZMnWnuCtMANJFmPjasgWW3PGx6rgLLSvXVw5qX7ZUe00TjHlhzlUj
TGNKS8fvANXKsUQWKa0l29MJtgeosJFPALRsZTXqB5Rz8+GFGSFFfDtzBYYwpk3m
HfDmUNsrs6azFlnKG0dVGlthSG03IL1Ki5Fgi8C4iwnTUSGHx0JSEbn0ZIGRUF/N
pq26kiingeRLy4P2u83aecmzhqGFzm6o17SFxOkmLaE0oiqFhej7RU4UGTl4p+JD
sCUtWmSdRwVrqfYTKaoNSOnCvr1bgj/dfUNq4D6sxI6gjS+TpG1LSu/+ELGmgxUx
6NvKTJRtJcfLlIoToP7IkbkNPOW45ixBngQJAXNTbim3P+76dYdq3xrPpQ8OIXoz
F6en5wNmthmS8mQ/TRzRkmcf1cJeJofIHbRhX7IoTXK2h82Xw6JnXzX9o2Mh/Std
bBv37THNB9EkWwT+ABPx15+hF8Pgj1AZbibYEOpp7c7QnzcqLdckOyYdKZRDbNLm
ravGWozrEhRVwCPktevdZXqAbUBAdWNC0BsM+mf/NtJ8J0fD3F7h/zWF3yyjUt/f
4Ha+nOSdi437yHh6Dq57IIUE7sL1WM5YO4ntyT76nKYEc2stSShTpjuo2F/90KbH
LC2O4L6j3Zhwx4rKmW8rQxr9KhSil8X40XwKRWuCKy5csCSk0XPq03P/DhF46V4l
DOvuObFw+aP3UTIf0O/Q26O/y52OzULgJUd5RIgVe7vvkNEaUbDuurJUi1oGMGFY
CBWTLfucpOoE/L0GBL9yvoeDk/uY3arH9eFnDeNVSlbBozVTvOB+xNS9XDGW202D
I9yxZW/hOhP8I7dwauNPfeswZrJKnVbFDJpyasE7RPeolySDw4uKlr0RhQAwMKtf
PCca0K+X49hJ/P0lcN9WJgCeM81EVtV1TD8iw+G0UyRSeHD1/iVPUr60uuwHc3Pu
1ygebFgjhhpC+KPOXqkH5FdIzJL3ubhk+DVO1Jo2q2El7anm1e0tLESAD6TK4rvm
CBGz2KitevVEQGN4go6iYjjBXu2AezY4lA+PQU3v/+hS0ECfPBQ7H4+9dywz7JLD
8d1ycpA1eLR+EaUA/y+0qm0F+Z4MAHMNfEUarU8QudVTay996eM4Dgh8Rj+tGFu4
3BwjOPLtVKyGha4BvgZpDJhEg5lU7agXtN83M/apA/D8mfkuZVBSEzBfLdlvZI23
FA1znvuPNOUMg1B1FpR84RE3V4ess+IlB5ThL8PXY6wPgZmoL3aUjEEi2USbi0Xg
ePSNDi/I3TU5G2GjEqjC2vqUP6Z6rAs8kYPynPsN0yGVOsSO5HkxnEPuB2EQUWux
nM8mHknAsu9SeeASu7qc+MKuv/sKHo9f+JDxR7WizYD5/+DrMsYxu6+Liyi7DghT
54Qs+dP1s1Hv1ydz496Qapiy7hSqgt0W5WidQKEbTWAAlnb0AJncNC0JBLK7UThH
aSt1qsRKltKOTRXLGPL1bwZc1KwcGlI0MqS7dSgPk3h0FO/6+IoOeViCGEvbC1AP
SGq2K2OdNlszD+SyKv4bPxAazF51Htw63HIPIdyGQ7L9ka7QlUdiRyZ/x93lBb5a
teJdKxrz4CnoQLlcizt9mGBt9qv6lVtfw3VivAJ6Jz8FI2+FyngRCNLqIaF/b3LZ
8MCM9mV78hQM2hqdHLdRUXvg2Db9OeEhPyBChTxie47duaPD7aNaK0s4ZACX/6vz
/7224QAGoiD+47fUHNpCnS1b7uUbjvnJyOzNJgk9tuxqCzXokSmYQXGY0XQ2xpCp
m73fY9Rc6uuSaOFlzb/nxlyVlhSRJvRayd5MJvhaPVeQlMdNYdWOLXu8XvuUJW6Y
p47RuV1unQ7TYD3kUXlDnvfgqLgOvCR5Q4Gspgjka4LrF3fJyvYsiguU4BZMxwSf
DQg6ZPE6M9NL7CIwkuae9iqLYa8gBAu5U0Zyfbi977sVNv43ZMvoOk5FVpmhTRqg
LI/bFdhhDB4WV9+NJGv3MpVhp/VHxWawdbpkLQ4BGgUTWeqT/GtyGcXX9HVszyGN
gKrk5DHSoS+fkkzCjeLfCl2ATtBgjrGvE2EjIVb2RXeWfxc9e7crLlAaBxHzD6rv
YgvqM6kTVjQ1nP9qeI2QRtxRGvzGlyX8YeKJe72GpaRKLfqku6V2Rc6rJoGY+Yce
VkiefT2r8h9ySmy2lPX2nx8G3B90qsgzAPw6g/V4tPaRh1h06cQspMyOoIijdfbN
SXvczVQQp8gLneRktfOSjSeFMFWBwGndAVw2FWMBl75HtXGLWmhkrEWkb4eCbusm
oKiC8xkA007hcwuhy7pwb+KmLKQVNnuM5Nq9OXT7u0FE3AuEKELxIjki5bRHprgd
nla3eHLxIOV8xDlFLUbtfeRjynQp6ecOVRVEKtF/Z/vXv3j2A71h6NNaToQkgKSw
oxSiO+ha/ZxHCLKauqT+nXkhlUE9V4031TPgva/y6QBd8Vy6nV2Rbz6I5oWArD6G
hfmEattGSqyi/Gi/n6KOtQprczhAnauJ2wF3K2mPa3rAsmfrdK8rVGVhHfGEd+47
/oJ9PRgnMcXy/6wu2NzpUw0w6zh5GU4ldEMx5zPRwZOSgUeexo6ORKfNYiY1XDpm
t/Mt2Y0jGkHJVAlabMaar0yrRoqB1yMMXj7aOtbcNTss4PRX6QtdDqTSj59hqH1f
U6vGuoyEfAYTEOi+/caZATyrSprtgsxM+FFZ0/jr76iqQKhPOyhCqaEeSGpcadiX
3V5WGbrq8TwSRMI2kP7OE/vzI2kFgQHVkxKN+06H9umz0pRtGOhdwcXx0IlzPUsZ
Fx3bEVmPuTBCENGNuk5BW8r24W7vPP/CTeLLPfPpJJ++YQSntxmf/g9w0CgCvzAW
vv/eR671sKzrg7fM3++CHPtQPMLRLa8C75qzr/VWdd2SLFIku0I679Vq8N27xlaB
b04sXRmGwuXjKV9lpa4uikZ/a4yK5707yILMwnMsJnz9D6cWlSwwtmFbu4A/idkg
5E38oGurOer5U9r7kG9AozNu0+CUTU2Dtrxe4wZzmRoc1oRzT17XfTmYcyLKBe/U
T5yapCFEMNTv7YeHOaq5BwmvQ9RIDLhw7Yli64XGlmSK63eceGyu9Lzun8+3KGsl
sN9/n+271rDxfN9wHjFGB0Af6liEBFkpVmuCR0GfZQNt1Q/aBi0rroGXexs4PaZq
LXb1dofCtN+pnLpm6uADI0oAGtoa/SWgnh0VtsCpzVc6I/G4uMn4dxafA5Bf6ppn
Y7EiAKWOhn8wrUY4K7MXP7CxpKlC3NPtFdP+mxbvB7X9jS9MchknvkM9UQ0xHWcM
CGO2aEd6X6u5ZxxvyoY+UGdVSzScWvw+fWhmM8mZWlN7FSBZUn5uzBQur7EtkfOm
nWrxEdNHGT3Kw7lvgEjiHjTwTg+9GKRIOb6P5fq7YADVD04pa/QGQT+YXPYRZSAh
rcgZ/hmz6CDwQmyd2JfBG+r7iwte93NgMMZ75/I3Uy67etfXrPVW94UJ21JoMMOp
DUPaUmCg8pLETK+PZK5YVQB/33mQkpRtggwPFRNwKS1KktTXjbu5HRwzjiTEf2Vm
PhX95cc0ZYpSEmq2it8XJy4JflJVqDTbtNJABf8kJPEfDeQ+0xaoWFWtxwL75g8A
pv7Yi6VqRE5a8qJA7uJ5/zX/oC+TCTno5BowVebGx/Lu5YbXfvl+KH12xYezQfZC
FGzVEwuRoVGnnRfUGNFLa5RPaZ03Bq1web5syabyu7Ma+3pJbv8efH3RbGVz4hcQ
3tM4QouXyp59K5JQ7OJNaE+z3MpQOx2jm17lVY0VfMo63hGR3+rifklO9a+wvZaR
SmGyg00On+kg7UigMSdiylBMuIi21wpuVbM57hNODO15kcR9ynAICNRJP1nD3EdJ
i7Bsp30gawMCELxMz+bdSmbdCuPKkF110uaD01tKJnmE5h6Q/Bj2Ezn+gRWfX+uQ
iy7oJTa2dNXxsq6XtUzrNfDJFGJzysOMIGD7qgn/6BJiWUWhv3sPb2Se+EUU65r3
CaeFiG22Mp1gENRzGKWxTHXdEewGpUgf+AcyZ2KU3/DpPr2pgUcIf8omKwIer77e
RBHfGEziwYN8l77XYkWJd4RONLxg4TlBvkCxLsOuzo6xHajXAtW3bweabfMQUFDJ
/+yqtO1XqdEvB7++BJqd2TI+aM9LElQaHyK4hU2H+SP763DX1gP/xrjPjkKWOBNE
FCzT+y+V7uZxe74BagH0WpRayoOBO6AoJxecMMXobPHczfWucwk9rl/Qk206sg4u
ZmgSSwv+g4FGH4hw73/WW2/E5lpj/lvOHp0Mme90pUjMe7Xc6m2nP2AzEqdR/4CG
xYb/dOtPIlHE8RRbTdedsswobmnIrkBVanZ0hq3qnLJG6oCHkSVoDJ7r1iyi7h9D
iP6Zwd0aM38va7KVcHypiBkRaMPFlrg/NY3oSIneiJBxjaByDgF958KKvGaL3yb9
avSSisRVfqc5B1lg+Vjvf7xrjzhla54xoRGAouWl1JqS9bFLKai1qTBiBp4GLHlm
hI5C/c5/0odIQJUn5OZ+0kVoIqL/wKEPKU63bS1yK16F/0UFB6A0G2l7yGNxYPXv
d5aotzEXBy59/n5vYf0N9HKQa62S1u2kCQ9ufk81s4ddl8jJ9tltw9LUvPfbN/QK
esBkERSWjpa6LQo1+nqzitSLe8WWXwjyRu/bXPHwS3874fTbWQUudwPVykoO1zZ6
KrQKOquDPHQfkYb6EVWhiBSOcQOz6O5l9rmoBLiaanWyKv10vimxz1mRuKAkp6gJ
5vRRis2T2HBZSOrikwsT6Jz8Fkyyc9dzs6n7wMAZgQNXwzTLj++eE5214omc6SPo
fR41K3nmyy5r/MRGYq+Muqe68YFWJ+lNVenh9acPktX0dfN1yg9CzG0Siejz30v0
pw/my4h/h7fz8Z1YR6hd+CVLDfIvXwWEmXB3xxTrh1pvuaY9IWSVrsWoxI5dBCka
5dB/STjQ1YPa3pCiOOPChPEPG5tr0OXf02ZOqoTrtk5y4l/g6Fx/LYphoU3h+DNQ
q6P8HCTHirpr6fNHSw5lpqNzyD39CezCO1o3+Pkm/Ijh9d3kpjFCBGoPPi/LL7I6
zhrx72eOY+3Lw9gY5pT/g9yqjc/iQ08pjenIQKOqZX0fM51+6wZz6t3OZKsqK4QR
oizfJwwbGqsvrFOn/15mF+xOhcUPaBHUs1BNkkiOUBQHapkQcDvElMwq2GbPO3Pf
RwRSJ2KxQZu43kIlGxic8MEQQ7EGJPZ8L+zXp4iGCIQ1+uKpDIYwx71wenDLQ48u
JobKo1zcrGbWnvO2c2s9XW2SDHA0z2xJrIhWPtr+nWQNKNEWOuACrfTX/156mRJ5
HX5STHpqwvncyaeEsyksDiil/wIvDJ/i574NN9DJ0alyYWfbVE1z7LYEBbtN4q2P
1ZrX4yvxkHFW2zpKx9XDzMkiC2qecys8FrYx4z8nSe7ge6wz6HXLpNRIUHn0CyBj
rCNZ1TnAJoJZCLaljVUVng6YgbaL57AADd4Ld96e1x8t/EA8SERDbNTwGH53S2PV
KvukqGTkKsY2TbuUwerB0hWSHel5xHLhibNwzGp2C9KluaCjPNc7XbWt+xhqk12R
KITKdhpc38vgg4HmcVgpukSI4wlmpi31SCz3OwQuF8YVNI0xaDCR9enIrYga/ff4
qlaEI4HDHius7yU5GFw9FfXvJzWWYuocULOnbABFD3+X5zaIUZbJ6dpEhZ8eYeqd
gyD31pAD95KTPR5MdjH8+/9EvbcwPUXDYUkNFi+/vozlHllAIESLT/7dKxUx4ZCD
WTNZepy5yBwoyRVyNXvx2Q75Bcxj9kgTbfzVh+TuDvPr9a4kNVweFHBs4lg/FDGF
GbTAwzozW1XiLde7ADIaF97ElFi7XH3binHuh+6ePdgF2AaijPkOWCZa4Q5POkoY
A2ldoLQYSyVHCSRCm6ujxmJTGSW1wZN1ujhdLi1PIaOdvFY86EqErSvhkpfNXSuJ
jxgyQNA+Q7hRKLyy9uT6W2vWaYoF8PhVQEFk9b6xvKVZmNxn+8xEHGmZSECPegnV
ss6EH+EgREHI0tC3TOcFeUG/8faAHeGfKYm8l+aUvayroSOwkjM8kJsho8E/ioQJ
eP/1khDVBI1i3KGNCKZ0C6uExPkxut81RZ9l5cFJwftXxU72nPvsxffEODZ61gv+
U4qfsnGs28cLu/V2c5iBoRaXBxZZcnWT0yqx0QPRu3mfARPhQiRdYT6v5upQbjZq
6shLE2BgxK2fUFyHuMcEM01ibHYqmmKsfGWt/6TU9GL6wRmyipsQxJ5hlpCBQan+
HLy8gFb9ZYJIoGYub8Lt8LvS5YGrdlZoIEBtXGuRFh6D3DkmGl14BhklPux/ZseH
hKCrKgmSjsGLfTAJUtnBqyVitiYJ2b2cApDAxkiZantVMvneEMGGzJn2G4vUCaxg
1KZ9xqn8q0voTXYEw4AGLm/2DY+MO8CQ7LplW7ndHIGmxZQ+lr7gaKIOuBARlgoy
ciHF0D2WH1QIXoAB47dYkXPQy5/ACatlUa+QiTcucQsa25mDLenX9s7mNBfyn0BC
mI8k7IJBM+vrrNhBf4cfg/LQ65Ugu4I46rgGZD/UOqSzUjA7uTqS2nRTTSiYC4uA
ExgpS4a+54tvZA6UnEqd7r69oH9oi2bQR5fY6YLQLuem6H3LW/TUKQ+eZDGZiY3W
cn2IsSt9fJ+7yfzBoWSAB4I0f2/lLDb3t+5SOXD3V/irwTSzWqTPuVfQ0glMBC3U
GRLyjgRqx9K0mln7anzf0+nQQ3jGWPdsvzsOjN+rUyaWXOUUH6IuTX9Nh1opDmFI
FkEfOUwjQwjW6pdvIEYsH6qzlcfkabgFTRhSkgCkEIs1Kdcetx5fqvmD9xspL/KA
0M7RxMh26E4L+UGEMAV9WdKe6m7uT6+cBEGd+AnirjYkXaZeQ+hhFekTabm1Nx2a
RnjYG4X4u/trq0KehH3yPz1/WcfUCNHoyKZ6D4iRipIoQi7K/FUz9B7Zsfo9NVDh
dA9+eNd3dB1ZVkwM4h918vYN0NAOUyPfpEX+IPaTZ8oeECM6TfIujMiZ7WQz8V4Y
afCYpH6vTrkTQNJ+XjHaKGTd6gMNTUQmLC7maFGfuOEWEmkqLMc3BwBetX+HGhOo
mt0B4UaHkonVID/gv7Va+w7mBR/frmWNIUkwrBba+qUikoKWOQSFlD3wXll/O3mW
vT0jfelKLlRqcqWOGvpWoNDNGH1wF4EP5EsxJJhvzJEONrGodMWKTt2XX/N1b7LK
bs6U1WhFRbLREepAmkHDV8FFdEKMYgGpa5e3l73+abovXJnGEnNRSEzZlau0HO//
7CuVLGwszPxyhyoHryBxf3FplqW1TiSr32TlzbRwu8rs7wtIL/H8sPd0TErAXQnx
NgeefDo3W2e5VrOtY1zS9qFDpNuOkjMV26hskh3NoefHS9kQmQAS6beaekk8AL4H
M/cWzf7lA8zx31Dei1JyG241/w0LU/Yzx/lQkLG5w41i5nsQ1SMeH0OkAyqDKqi8
LJTFiq7NeT6Gdk3ien23QY6Sne+K5ywRiNUpXFdZEFJpvhXylQJv5ClbaNgDtEU5
ERUl/MN8sdnTNHoI6M4RylEyGW/sM+I9CcKMiUfQA5ieRwyNBEXDXCLp2JCwuWUO
iFX7BkLiT8fTYnYsYCkHPQXx7AzXKpyp5ZiSXTygq1OFQJW0OIAS38CVnLDI8JlA
I2RtGX2/5b7eIcEHZMm36Buvy8LdvbemJ7dcsy1PkkqI2rjWTC8Pp2vS48jYhKpL
FvMLr9wohZODmGvpscyG427p/FauonA0lLTPpim6HTmRtTq1eef55ZO6b8769W96
lp/4hbvKaD6cndumaLNwndDLjcMsendd6UOzh73jwcIhQ/6wdzcMX85pw+6mjEup
pNzdDs27soFmpb4umsDCl8SP/4N8vKG/Uz3q+6GznSYhyJOqA+vVJ5SsnIE4ncIy
y20bF8KG3VlGTmN/7IZA4cm8axVfXqVqWQVC253An5cjJFcZPw3Eg1/7vyzucR7V
N/MPgbipTB5psloKVli7VMSwomIjQPGCYiYisDNEL4MkWirv8RvZ8U2pKxtd79fL
2rgC5Lu7bvQlJsHACridHf5Ki+tGuuGGL4bu7vHOsdedd+fpUghfgokGRpfNKzih
DGZLFhWGNMQk4ILIndKg1gaUz4RdRNo5gmHVb7EY04ZI7i2uTeMNxGmhhH8nP0mJ
ApTE2JMqO2eXtyTs/gr82JoemCaBQrm9XiMHsZyRzAuwBmysQ8Yt/VMYXCVyxdWA
kxur8md2WcyJE29gq17TOsMxD53n3VxVS5TLqQZLt/HbN4WfMJ4bZcEBE+aIPeTR
lM8MyeaqJ8NXWRpcbpsARVkgG/d8AHlqZOQYr58NHesgT6EWAieLme/0ZwdzjnNi
Xl5Z4c5UXmUo1OnNrcJE/LefExLYnre7BNvCGOfG2PYu0j18b7tOHLgk8392Bb/p
iflV80NHP5TQed9EWLL2zlA1wObl2XIuB1R0n2zifFn4vshYZgw5vsZxNa+65myt
6GETihRtFYtpjx/4PtiJbjQ4OH/7lFBzsTC3N/0Radf8N4W2LIBP26g8PvW+Plhj
hqKKOA+e7S+VQ0O6o8kesl2bZdXXbXO29CPNd1uRyzA33rwnSZYyy/+pb1kTDc+Q
mOfqTTDB3YMJ9XqE8mgd0ULbGLQPxgHnjkRjxQMi3TSWvuTi7MlLMMEXj1rXKZxD
xoYed0nlGR73/5qq0Avj4phx1EamHg2ialFda27L+saGq9huDRMQ+nmMqNRcQceA
h0XUccdEFwVwlW3Pau8CAdXD8uPMfoNokv+BKGU+ZnKLgrBm7tGcxWEBh66YQERb
T9DOPIK8Y4tf037nS/Lrgmaf9InqeoxMRP0Am001uReUu2qLEmBPVgruzcEgCRht
A5LrTKrNCVGMegUmm+/O0M7aRlfs7lnA6LkUrXflW9fLF2TsYusfKZ+Je7cM0/eG
Co44sq9bZ4tPgERr81v+hw+FkWCjwZ9g68ej76UThaQPKtz0u7jVQBzB+pryEzB1
4TmMSwYwa0yHss1kzRkPwg3PbkpzIu023Gs/ko6UdXEEnTyW7qe0A5J5w7KqbJeU
atgdo9cdp/AtxmNG5BTME0YDGtgWIS0sFuL9xqHh1xAh666QC2cO75ggCcvt2S+a
RFZg0kwpd23FMTY83zCJU5DmRRUO0eBWwKy/CO9CaQWWOuwfokChz8qDF9OOTo95
OTE3HIa7wHps9EPjcEH9EhyZQpVM+n4AoE3czd+Y+cyx6xyVdxjfie1rHxA2xXuy
dOVD2zgNFFvPSJLIqhGnhiAcJWCo7l0SGYEpWSkkXtdsrN42978uk7VQ91YO7+RG
VHMTAMR9veyctMM+LQN6mC2Qw9H6MsMSkZPsjkeukTIG8or1Bc/QNsEcp57U9lWz
VbcwuN9d6wxahvOpCQUaxbveKy0tXvW54E6Lis1zYXXe1mUlbrjeUcUtOAalvnUU
AfClbPHue5duyRwGdF9lTt8UWy01k0W4TpTKFNJUN4SzBhopLuXZBjhbBrKKGVv6
TG3ECWDugh23+6xYIzqyW+DNWT81u5RFv3b+aq9YltlSrvJ3hHoZtebSe0Cc0EKa
mJVQgxS8nscIHc6EL8tdJGkhCyQJXSQUV4yEeE0oNDccWn29tU4sdqA+2h5SupDN
nFY9h5s5XNSEynr2Ox6iJu5MLCwWQeGASlTZ4ft1BT8sQQl3XnKf6jf3jeBxcSr9
5z4nYb7wVw0LumgtAz0k0G0LzqF2gxS4J4CbHiGksl1iv+u9laa55GDWmHoV7fLJ
Byt25DgVIP30cO8gMR0ELXon/OKKX2pzyKv404c8wXfq923b/Gaoq20mmxpJbJ/z
2S6yYoR54jOmNoX8dCEtMBJI3lqf4cZ1A9pEM4qErwgcabyF2S9tj3egrabqkNxB
EOdpJSETNPxoXH3Cx/Nn2+4kXPHvoOAMf2Ttm65o7eoj2eKHKH/eZdpvJLHnxM1E
cKLvm8AKFBRvqfBBB4cbdip/Lmo6ZdMObuJW+ubjnQHGq4ZZWmCfonAHRPhqIPnZ
YlndzGMovnrCYeg068RuTl546qJz/MHwE2kS7Ai8LF4h+9PjubGveB+/5xaIKjcv
RWlFWTQRP4ogcT2g6NMaFk/HcF0fSkqdTlUlPg9OzrUd8J1cr8pCWsByZ3/JAlwT
BFXYaIZr3SmWacVdVWC+m3QNtoMyAtY5h595+ZWvP57Owx5TqO/7Vp1sCIbjl8FF
NokrKcMl2gYEmwL1RQQs4T43TayXGRgR1iAjs00IOoLchuMe2kCQVBufS4+jkkad
V00tJaRpoCTnX+v6MCcY2aGfl1ezJ7fFEiKllc8nCCkEYpEzrZC+MfTZiH6d0vEy
+r+plm24lR6WDZqbVEtXEfq+7y6n1PNipZEGLANc0CBU8IDyYY+Ilx+1lSQ4I0MR
m7h6Bf5bvYltHzrCLdqmeHRQU1IDR4cPp6cpZ5c+qhqmSpTZdmHbqx9bMudHS822
jqWu3kT2wAVpqg54fukwbQ1jCK3vfYCLGWLzb2je/Pi4uDF+wBxVWRJGN8NaaQRv
3ZQzV23L5ijxXkRkMQZdKW1cvqH+DEotZoWGTpLY0heLG0VkE5e1bfFOjvr594uf
3Bjo8s0fK0vR7ejGXA5GSTzXY/pKjfLStM/LdGIzsnVBIxWiINtv+9wjdCk6rvsx
nFrEfWoEQ0TkQhZ0TRkRgwb0S93AhpWdDjAtITPNwkm0OYDzSNooh3/K5sV/VttM
Yz4InWHwjbKEGe/hFPNYqQHdYFanAxrQDbNBeIDvc+Wd7c5gH7CQ7at7xWJ4tS8N
ZrW6HrUWfVkjsjaANHxloDKUP5baf3xF7WGd1QbnhLiaHTAgL1eVimc9v/ychLRQ
zy36tl4dwYcB1OXmGR3m3WNyTVVGVldmNTikJvrJe9qZVkStt3cdDWBfvOXaGJ1w
WS9TfsBCSuxMQwAXfoCO62yN0d7a7tMvup7w7N+tbKeBlytt34qfoPTqyvB2qPM7
Hr47wIReROxr9TWNxAWZEUMj/9E9UniheE7tMeXiHs8eGUGgNCbWVwb9Cei05c/H
uf14tF1w3lwmLXSyK262BAchfqhOs8khNIsK7nKpHL6X917Desi/ofYSOb2Dmzl7
fJODvnqCPNBQ+/1ZZHnlf+adasz+2nCstLmRDUpm3eK0XBHqM1Gj/RluLYJReqzS
IByw7tfqqd54+/Aa1P7ewV7cWgDyH01/2CKIbgBav4LZ7DO8V4YjisFVUsxStYEs
RkHmuFv8/HGvk5rbKND88EXdNC75fSevsIj1T05K0y5Qt2FqqmMo7aUuVNSCxzkO
47sUCmriaLTq4SJwkZzRLARF7YJmmvIHqCPn2gcQdQwxnfQYKQp/VF0VGoRN0hBY
hvj8sTPog+T2YTdgnAYScQyHPkGjd4UMY8CqU+6SG1B8ymFiEDDa5m3np6xpHkhG
CDtfaLH4Q2GJ3PjhL1iVykNT/8SlpL32UWi0fPbNOQQhEHhrma8cKdPRyX7G9Xp+
WEJBNln55umsmgJqPJ76u7urUOn5grRrwnP2HQpd0f8j+04yRwi+2dnhshdQfWO3
hK7dYM9Q3vV4xO3loTiCFBF69Jd9PzyoFdEKMgkJiWzyQI2xt5qe8eFDNyXPxSEG
3VJWzomjYbfmSY5Pf75KaxUqDLlLM7pU+O/1c3/voFt1wNOppQYOE1I9ng/vj1X1
VgD2IX2hKCJAXnqDD9DwProO/xH5VBvKQB5xzWHg/lPopOEbDXADVJeKhLmKnh/d
cXaWBRzakjxmvvlwx4UPoMmM+QM53WwDA57tw9yvsSScsxewS92QTIbxm5dG+Fti
Kp1HPXcKdVKAvp8izbNDTb/XXHQQhxXwuw+fgZ57xoT4o65QFPPMqaPPX6h8cz61
nUQ5PSh0ETt+xJtzWn/tn87GH83UNRYMc1JHCUfYEea8uCiEzG++vCmGxHbif/ef
TLxkoi/AMPN7s5zOR39QYJkCObO13oiSc7/v60PF5yyfXNv5kOKofoY+6q2uKsPY
kjFVvYSYIxhsX29oRIS48cUWUCE889Z0B8H2AwLhN5SibzqfU4im2GwhUzYaFunF
ir0a1mIfOmmCsZDcdeCzYtqdvdzqJJFETfskYdU6KrGZ1Us4E+RAhFWDxuDzppzJ
evMJGhkh8xsOExZ3GW7Oeyq65Yi91x3/HmBDQB8mwxgYmCAAU2DL0WJOQ40dGf82
x+NyltL5zSaYb2kKKZPKryqNt5OxNSgRkKoDHd4XVa5rjqh5ofBPxD7Cq5XHmkM5
WhVNtw28qFuQ492M0b8gJZHujTsydHal7cK+UZieXct6bGyjqthNlyryrHyfBaEH
XUet2mavJvZWSNvMB9J3PN/2l9I17HCP2pZg0iJkjia70Qbdr1991TxJ0Sj8mPWz
3U4Hj1SNLpfOcwufl8Ya2kcxi6XtHg6hDairIrZofdl4OEBZ49OiOA7ZFBufGr1e
NmrlCndiaclBVoNSajRuy8Ls9/lknzc9JqmyG9/mY1bsjBtWePQZHCOaNW20BHEY
RB/OWL/QIxLK9Ego/YGhX8LzNXN7L2Sx+RxFltOriXYx9Y78eO696v1TVpagI2vK
Rb1EbaAUAC6BwAbTZc8SZ9v81wjGcsEFcYCJ0lI8DD9OV3MWa6pW+ffhUPg6iwhf
p/Fl7NFZy6cOKwMnk6B4YWZqXmdgSHosopux56faDV5+UZ31J/+gV54oaIMuIt4p
syhcpcfA3q11x+9VVKrtT3zLPQ9GgbnNmey6oWta0TuGeAejTqtJXE/69h8DuEW/
im0LC25DS6wiIGraJEWkIV4BHcN6Q/k8jK8YylpeuuhaDB1ee/QikHhzOwi8cclN
tKff3qnGHEBXP6t2d1U6EFpusWyHiBNe6qS+MAoLMl2m8OE7YU+o6GV2xzdrgCyT
6QkVnTI8EgWVzSQeMxafRKzPSW+RPLbNsrTeJkUuEFWe87BSAPxmizW9peiQr7Jx
+TWvnqipYG1rbfYUW7IRJBBJ3B3GTncvTrwsVTPXaufhb0dPC3QZShReUjCQVEAc
LB4VElo20hNvMezwJfJnln65HvHHdNwQ6gDkO6OCSVV8lRs4BBDBehAOh8/4A9Iw
OGGBvHNDS1ixIMfJVlVF0ISjl+j1M9usY/bUZL+Bnm5Zu5SRLO/j9p47F2Wum2eu
SHzMrelaNakbTTL++UM2qZAortXRe+AEEHwjxNMS1gYehOSQRh4q0BGxW8oUCLcq
duaFUMaJLFvFaEULxO3aquBWrRlU1eLhj+FsiNv2gqyWZAQ95XdSfi4BE6oXIKe7
H+A46mmAnUmeU7j4V9q42RIHN864VZo1lyhZLXxmWSVqaUnD9bwZOxPrAJ0IepTy
4fxi0crnzSH1vKc3HvPtdLNVBBDmabdvQhVZfp8+F22xhLSyQEyGc/8uXXQBWgc6
MykAggWU6FvrZYSgzFwkYZyieRLqSV9NImRGZoOFqPIfnmjnSgAWP+Myd+fFL1mE
uWvezzz+12Wzkj+xJs1LNmuRyar+l+AbCiZTzqQh3W4gBxWSuL1GVlPUNht+c7pZ
HSfKKYti+BAktToRv0FhqBISfyBblNtlMHywJ6QI11CZjMzS8zhIZ7677D0qrzS3
+7NwougYplmlkijzeDfT8U3LKcUZnEOhNasnqofcla2aK2ZmnPPW+ZslyAbxm2Oh
Uu8X9AWlORhQ+kT8pvUyB8Oy5zxZ6kuXCVImqGvKRk5aPNHpfwt9DbiiWLPovKHt
obpeGmAPTI6RXvyLWRr2XFHWzPWaFiIlaqZZxHGn2TkusAaLB1LGawJ57/jdWP7p
ntarp21EXLmhuasihylOVAmoA3ca2KNKy+FRoYfd5mC4V2QStMun4RS4jXzKIz7z
WEAnvIryvfUuZrpSigasyu71SaOgD7GzgbM8cSzaIacefggLFYrmV5HLwfO5sPV6
W4okGPr+JX+ycY8PX8z/HYGSeoo/ST9qbSfIa7ny/u4MT+mHc8cZFJI9J7hM3LT7
Dma5kGYtcELtov2v/ko6sZPBjteprKXumZ7GQ9dgm/xNyBxfk9eukXvtCOZQzbC+
b5Jt15v68CuoB+ProqB4zE0ACicgBPzdBKaXnDd1p6xCj3iKyWgXGcwIKdRJuGSz
fZSI49M4n8mAmvrlQx0SKiKkSkJL4evu52Bi0Oh0C5wgCzBApuD//hpWGhSqzNC4
iYcuJEPMPr1Ek2QAj8PpTFJQiPPtbZpfgCquR+MNhtmRQ7JKcfNBp8q1HdR32Llj
o0EOmtkzi7PLIJNvfYoLM1mvJPYzHkh2kmRGMPAPkZPtVDntBlJcNNghLGBTO9wS
kERo2g28e1QoB5s3YF8iIHPKPdp1EeATNe2dnhHYW8aZgtAUGP0aG9FLWBhN0y4X
aNT62k6i0/PbVwbfnQ5xrBz8HoCMdSBV7a8KNUPscWGbfrxyOsHanMmGw1mIMM2C
n/sp7Fy8JhehMxJ2z3CYMVP4IGG5qYiKajM236dIKoOgMAU/DHlwKfywT8aat9Et
kt2Qybixiit1mAbeWGy//CY6+o1Dj9HCBeSte8rk+JI5e3q1nH5WdRwFSIImIVcL
mIbSF26ESSQHxD74sY53aSL7KSOwewRyZ264jXRxnHkEOlcF6uy4KHwa/kxkWReZ
YDuMJsErd6mq9nhNKR3/85Ihfc/v4sYJvHbBxUH444rtPb4y5s4VSuoa+oLqib1V
dqIYcuJFMi4FSrQFLI+6x/d9nTuwKkA5ZzpRPNQveJUkaFpq8uGeSvn6YTkcyHLx
LTpVyQ+kUS4u1YI5nMKOREmZOv5Cza63+z+E1Qv6YZZViXVxDO4SI3vB3edT2F9x
Me/EOeDCsNCNmWTFpqdmLAUF0P/wujqNWjQsStbZki74NWnFvRcTdiNj1qLfU5AE
AiZosmBumfiz+HVGAWU5/mN1x0Y62rSne4Xnj+tWW519Mms+E40/uAC1guTBJoj4
D5lRpTxKdjkrxI/gHIxodA95iUtcRj6heViUpaDTGvMLs80hwi9/VqhTkpmufY9b
REbBExts8Y3gF7CMaxd9MDtDQHMHj0cms2Uuw0UjKrHEXzCznLlnvcpMXdSFSNv6
fGVQW9N3cS63kef92WaiFyQTVwuczQM/k0AdE/+WlXMgubMYKO1aGekpSgbeH86W
2hohwQuYL+93rXMBpiV44YPXLoQmJxmX3xGL87Lyl+8N2MPO8p2vg0S8MtE6bRZk
5ejogeTRJHRqceHdI+NZCd76SEd24cnATaHAP1easpRlMoQgUdINp/yoRN/VHuEn
bolnnqxbxiIdOTcC0w5nRDIqypVPDXV1ZGXi1t4TzN2q9yNZctzvurbXmZkvJx32
Q3K4LqaAv/zgoB2tVrg/yzU23dW9llULk+ePQ0UxQ+zRiyYqKB2yS1asinRvexSf
9T8b3l9rt45XmjqWEhEMtd+sPxTP9Vgb9aZnoDb4/EkoGJsic+Gdk+cAoosxE60L
YX51l4VTvYsRGs8Hmey07yf5kJH79ocTUsrvVhfRG5c32B5VSXes6XiJMpTQWA+N
rmzEloGdQxYUzQwYPVexlk4IZwn9G5pW5D8GZInbRmjCuAXpRxiBhZTNv3ALatHK
b41FxpFkLE1kO4wwJrlJVSlqy/ivL2Dk3XWT+1NYS3wNAlqpnSZdcGjvUkBTGgLo
n6BqvEBYlLfJuYishe5qN3XieHvHkwgFYSfsu/hFIPkDMzk3MfSbTgs+9cE+EKw9
AyYogGW5VyQxusjOAHe8CFSbSRPFucJz71A4t98kUYlhIBQhbaHmo7+n/kfQfa9n
CdjfcKaZmUKBWvsOsXXAY9Y3Oc5jnuJRAF81vmMdVmPoIlIZ2HPlWk64+R3spoze
jA++uDszZzGvhCL3KGpIbhAEwOiJ4nfA2cBSYsxZj7A4C+EFtZFkKvsE/zNVBKB6
pErcU982vuGDnQVgqCVBTv3SYnAy9LdMFX181JWWPI0Cz6q7x7jm/EC87kGHc1ec
v92equmKIdHmilWCd0+6PwC/+bPII/ZXQwSAs0L33Fzoz5O2XXzxeDU4fg1YtA1M
Pv+gAXA/HaczHOkg4QlBuT0nZ/pfsokx95FcNUZ3j3+roYRHz8rFoZlhTf3/kMtl
FfF1KjXTpdrqMX8JIZGNar7k8WGFj59ffLfNz5FcX+Krv8agVTlFaz4Tj74NUUPp
bjcQVTwkKtImD+SDVaM45qDqUkwriWx787kvPwSe2Ly911jEwF43nCuLn2fYHRDX
qRoSq9Kod/c/8mhyAEraEm+KFvLMuDeH1dlwomKnV05enm1SPxWtcNZ1OH2Kddq6
GWjccmGZ1rLs8FYtKSq9GaD3oCOCFWlknohmXTmsG9oslcT0bPSqIJSLFKgRbGdW
3wRmQa14/GOR3kFne9qs1URP5TJ5t2O4UJXZS4+/LzCu1sYslJ/E/MInWkSFXoMv
rg4o92Nw9Uk3EeX8GnmIaN7vG3tXyYQUTV79lye5Dk5+PsAXnl8RtaXHSxxmfuxW
uzYB59zS8fU+VOcJxwlnFSzxMJ/yMvZQ9LN8qd3aRsmhmIS1cCc1tlTkOJLDXEn5
S1lqQRQ950HqgwdHgtRUtpauxaIsO2H0U6wGGoi2dZb492xIKaxjZNCnbXZTkyvs
u9Ynus2XS57JTEzu0vXj6RoHCpdYFD6JdYShgqrASqxnt9C5P1OdkwM5bPUPXyVU
pahKZHBcHJTxWXGByDmWXwxlxNWEPapRpejQTjY41kV+d26lEPEMkIByBoVZ7/ak
bB1EmGtR29ntOvtawvrra3kdBKvfz//OJ4yI2oISDXUGneY3+m+8kmsnldK6CrBq
zR58upNB7tv4gzGXLkRG6gDdDeDShBK8T24ia8uS3V5BKbVqGw3YU3Tn2d2H4yqo
r9c3XO6TnRVEMLictaa5GYkvgKMBBWfSgYLddmMYhRwkYodIfvxZkUV9lYadP2OU
Q3jv1HSFKEzWfwximg+p206Iz5B7OwR8ro3cFtKYVkw7HG/5OthYOZI+N+WMYYuY
OSa4F17jci/NourRfHx3dxG0M74bpqeFxEl6UTqhK+RHa5UbQeXIQp/xmZ+bEHF3
WB8/wWXaxzP5qhobOsruypT9nMFj0/ZA6/6ebY6KCOWV2mANJaHzPl7dL6E5IIMB
e41hxrXcJ8hCdjA/ipgqUQx6phmb3U3AYyYvkI1I9MT9J9KC0EoWrHm9HCS8pwOe
BmH2amCXLPgk9bL1yxlc7yExivlsajaulqr4GybpHLqsVe13ddQIVc38piSi4ztX
kfV698lJlBCtuI3Deha39sVh1Q4I8HR1RK+lS9VrO1A+j24+4QSuhju4om3ns1fl
XgHlClwp3vkwTshRQNPWxBQP0AstZ9SaXhP97iZZ2jAPfPTcAI1jv4/bSFpnwu4h
yyKITWdwQfYoer/YRXPG0MZutPdLPoZaJrmKi9L3VGwviQdDb/NsXEyOBkDHyKdl
v7amkBYvbBAgiRqaukB/AP2jifYCsHlHM+0M0zeVnaJ1t7Jh44zgv1fErF9tDzVP
fpvkGBzhDJBkqSK3IgFLCGuJUr8O8OA+Bu4FR7L18L4/HU6BjCXy7kh/eu0OM4IZ
6iJggLj2DzSYiN4vuc0Fl+ZfHJ89da9qR2TLG79iDI3kG+5H8e4dS+UUFFrUUJaF
zWGgYgp/cKlZ4QOXmQ08Tm4JNYhb95LdTfnRvqJsCm5XSvFpuHv85cnIAGkiPU7D
9nj4KBAGJskr/KPRqoojH5E+nWtUBdVGTb880Y+bfNWxWW6LZhKG7R12ONZZpN08
kyKOkaOkyNwv2uEGM7NRUc7MLS4HUIsrSp3IF3NI7VztopEkd2F4KA6GyxwQxiMo
KFFE30UookIpW3+Qg9xrzcVs9tP+WjxJ+I6kFZaMoSy9OUMjH7NTz1RIp1FAKC+O
0JqTHd8g9uRDzGGHChBoQVBypoiEe0cRrEnevnlC7g/ChMBzAEbTxrc/J3agtBXA
VLu0bIYadA1pBbIlBaDRULR348iflUjojFnFx5DGhvlfEmKMfL3FYdB60fvoyzjO
Rywh5NEAtoOsRfNNV1MnEoow9FXmHzYPwBfX3SD3gAPXwS+RT2upPfjaMjOXULIk
TuNgVKfxzyD0LXgDCte2m5HIJoQ0E8PNYptQVqOQX/7qnlS+RK0uaQyVVQDk5BxG
+Iw+EdS2ISIvCU23bWk6ArST/RHQTG5ktSltpv0Pq2zEyri75jMxr9f4pZHO1eZa
yEL+jZmPozVBhhaILWM8ZF1bqnyKJfcnzZIzoawrC/3bRaJSzFcJFm9N5NXmquTb
ZTDj5pxnlkE5mj3jHJTG2+YnSpZ9ksHhd0oUxoGOfAXTB5ofh3TOWqim21P9PS7g
PWsdnjG68/75TgeS9UMYnM9V8rocZA8IrVj7U8gOJdlIB0tQDT8ZEnr5ljfPjocL
MKXF/qqQLtpTFKdLlMRYAexG6fvoSBDfXwH/wj2wX1wrd7AS7xILyLfCEG38EURj
RUniJge70Zik2khKeByPBtEZ8C7dZ/8gZkOgqovZFmG1D0ukSaHaGmoPKQJYFbhk
+Yuex0NgEn3wdgIONoa6rqsbwdjURc1JAv/EEFywVvrSpMb2cqBqzyA3aaOUdaL1
REz9OPJlZLLlsECEebij2x8U+Z0Q3ZM4puQQbbqsfhz/ERxTSSlZnB/IawCo9nQ/
VciBIilUA32ZJsFiN13BG0bBMwXpIk8sM6Ce2U0n4u5wtw52UgPLaIt7SXnQpHop
IBe5X5+KoNlMefyI/rLkR7kO3ImFOTJITcGIUwKyO1K//Owws3+y5ssJXePTbsTf
gPwzXL5/paMZUDfdExkrxEBse+fOFkEV8WBTk5kGAfYZD3++sB60NtUxtSpvLgQk
ccGD43KqPqsXOwEZuAKQAC/Ja8H8q+1BhmcP/Xqm4ToLTCfkyUrdcLDrZbBw6CAt
tFkMj6BjL1vhAExPUJB/rfoYpiHldzB1Y5Z47casJuoqCWQKBBIZmIbB6s+lNG92
8cG9Y12OzbMEoASsL3dpDVeEtdXfXI2hOyWTJVT3Fbk992OfzkO3TbCkxTXJAESw
kHezZl+YhbTm2xD9ZoRqjzCEGPEZQeuozpWG00wHwg49hK41sk+kwFUpztIqLVdD
YsLfYKLzag6NEiQp5qnk7mwCFreIJkilggxAaWJGN2+1Vcqg5VBJBdBAW5s9Ndrq
K2ajXWrVBKT4BwuafOkIjpFWpy6CAABXzjuVIG9XUulCruR59epOZC8iNE7U7gxx
KT5HTvg2pnWAUaekcqOebufR3Y8+TzAjFAK/7vsG53JS2k7tEzv8Jd2RSGV63ogn
w7jv/NwulxjHr+aqH1Zx5GZ6O+3T2iXjcy1ioOAenrbNRvVpkG6mRyd+rGkRi6kH
IeDomJFu/kw7wC0bURqXibEwJTgoxXTBHv0gJuOnIiKrnGxv8/gRVn6yXmczisBm
R0Hw6UhV0edZi7Ff6n8IYGS7gDXID1/1V1gyYCmekg4bmV1MaH3YcOhtVe+gz3TL
mEYV0W5g/KVhVM6OJdI2/OrqQmccSHuReoJu3MvqQ6wIFe8pr5JJSWHAChNHd7PO
9GQu82MaNc9FXB92L8sQ3RlVbjJWgWS5zKxupwhvkrZoXVypMMCe4NJpHxXVzjDf
ZHVAoRDADjlnW1GOiDZ1zHmNACIMzOhWGQ5pQVWs0Ir5c0hTmlSn9jr12XQy8IK8
l6YEHLzYbXPWU0+A3Yz6VjDZWVHvGVnOGU8Rsfe+jwn8y1PCcyo8yb9s7zqMkzIq
RY2JXpxNnuXQI4hpnv/jP+Az+nKNsok/0SclyotpSOyxU9veaF1PHjf3qoKyWE5W
uuxcZ7Xhfb9A77lVBseBSPDaMn4PjhjOq9WUWttY0nkhrmPvt7sYvqTs/ztfsBwN
ROBN704CYr478N0jl7eXHrWVbWBRXtKY+jaJ+BbFOHuO5NgJNKiXFpI/Ykp+2+RN
3EmmGs0j3RUdcGAVoe0LsDQaZQeTYOp/cy5CE4kpVuPlDA+r+hLl4nvZmpRwtd+h
p9d83itGwY+TxRsn/JssN7b6xyaYgwDK3OSoHDkcEDFPZAQ8PlvmvPT9jf6mHcud
PQYvsnTXsEOTV8wL6qUuil4CgLNT/nV+MbLFOGbdne8L1PChdK/hlULe2Ahiysq2
8AIilK/xeTplnICzHmJy/PbSEyf/n5cA07SavTTbopDS3LnbUbFFhwpq/XA2z92T
0C7jIDn61VQeeR42rl0o3Iz84S1LwtnbtfzXxCkamzsswB1N5eXIGp1Kj+mkNl89
f5kovncmX9bSoOEzM1o0Qk/zNj+0WLwDfaXnk++p7oLkatXWycWUbaKzpFqthrZM
cgWKyk/gLpRfeLzRCQ3mX7biUT3j+eCwXHxjU2AGRGFIpqItU7VS3L1Yq9xUBr6A
yD0b8uaqdx2KyZArDloTemStbOhaEyzprBfCkU0AftlvZJ0QjYfGfRr9uBey/CQ/
hWJYjGGAFFQSXeXYAXMwlYVOLsHpUEEJg59AYYVp5eJ0iRYawSrs6Vbx7LoaJXGp
wOrh7G9to4cwvUMjAYsg1Q3OE+ac3y5g7dsSDhKTGLe8v7tIPsU3EZ8TCw4UcuX9
NRrRSRH9gSi8gfHlcuNXMZJnURmYtSX6ZLktIn43MYVtsWdUdjxIViT8MqYfx5Jz
5AuEMoLzUL7cOEo39X+sFxuUenMKD64a7+nuIGe6/fFazahdvBkkuJqRWLEdg474
Nk1uCucQdcsOAQ5kRuo0AZ/wQ9Fi9oXNfkzii0304C40c5uxhv3J99v6Kdx18eA9
Y2GQYH+0HQB1/f2sLkVHFhM2USdI9jRKorKp0+U/EZMQBd7FAJcc1KkppkP+6L1z
X3BSDqXg+5MqRX7+rMEcW+qgaUQhOaDmXE4fTL7CvCllUYz4rXyHX64/MlTiTz7V
OFlPT7Qy39wzFFdObE8iI9D8yOGhZfCeC80YY2lWqF+9KThQEnXuRVFwepNVsd3j
GUN8WQ+tazemyBi3ffylDMBAKqmIzeQTi3z9X9xtxfXOOXzHVm9n7soLJVJ9Q2Wn
4wj53AoAKk6Lrn0w4MjiahukBjl9F8EOT95ZzYpUKZmXxgoSx3lVt1wLM1vDZIA7
ODXEH8Lb9kJGtpl+3pb9Z2Chm3vsTEBXEViJ8NbdXIzeUGOhp3Sner4/uUa3qimv
JL0A8rFQNXsmqMqr43jekl4LhL5tvPGUtntWQgRL9x43ht//uaj6k/MmFQGm8r4G
1MHEk3b7ktVtMqP2aKTJXgiFehS6pXzuWwUd8ch/9iHl4WWjy17/Uq07VJEuckeS
QnNegBR6sIeGrRtF8JWyfB7w9PSteVT0lSdrv8JCI0cVhGDn5+6FyzYssJINoFgK
j+BZb5z9yxX1SnAolMVT0tqVnoLyaWSH52t/kKyLkWQh02rZgHE43idUQ5N2eQhg
X86h8PJQ2M+rmmkImZJNOgW1bEslYBpdDgpvaHew6p+jAJhde6O5W39dGYDMO18P
PRUlOkUcWs08kq/Zhr1nKZKhCwc5qfsQI4bvOTOhwM1T8j1skbyseYaP7e18p81d
tPNFbrHky3KaMbj3dVFeGOY3QAaMKkoeb3k8u1mBf+MOSQMIwzyPg3vP+0m7RxTa
PkfCM5QWtkkZWp4Au4PZaBA4B3BsjhJRk7kaxooz25HesSgifUklEKc+u6ViUM0X
DQW8Z4bu1zSSbvNDzpDeAjnXJIUJIOlUb2udWe05dsWvRRVXl8DhHxFBFqS0L0Z8
knaai0gmJzkl2Ji8ajG9WDVzxNWEp2cnZ3jfxV9dFzJmhwveU9JTx6wecoE65u57
iGvqSMeAwMXE+B2dkM+9pli23q8PtsOC3xYbR4fnvReqE6XHpz6gDU0EisKPrDz5
U1PcZITfLhVOyKWHi5VOkPmvyflVWRRTT1r0z40EZVQqZU0ttRiT3TVXWpR4T3Ed
mtKbNDRWhdp2A6rZhIDY6uPXguj4i3lyyvouYGLsdyCD1krUUl6T19Bfbru0NKvQ
v0hiId939rt2hrswqUgfFMfFMXiAo8Wx3Y9X8+IR97WJigHbeMB/OdBPu0VkH6ZJ
f82clyg+/z3V0Vouh1YnLVpBq2mOvBSDfee8gt9V0iOY10XVNGkKCUR24/Zde98T
XEIEMcIHlN2hbDVrGQqKHwgeX8cXN337NiaKjfn7YAgTrQCX2zJy30ghqjlPaqVD
Ho+iDO69D9dYk8bgrpdqJb8h9lhF8BT9K3xs7Xor0AM1UTW/ap/APRroKnpbsS3c
JN4uxtDcryrg1z+T+B/usDKBU0ldCw2k78nIUB0gW9L5gVL2XjgLZoUssaLoIqZg
z61Pt+vniMRj+MNs8d1lQwNxaMmViVzKfpM9bbocjCMuLiFLyGq9EgkMIraSg3gf
CcdSUm10mss2QBiHqxbiSo8+jEf8i0Yyn2npaP8PFlpxysMtbA9auuJDSGQq7y8S
rCJNGXfUQnAK6acRInHRrurOzC6xx9xELQGItYhh0AK4OYfLY5KQOIFmjsrcuzqn
vn1kunDVdJ0TAkOdF4P6Pz7bC2OeMFs2ymSjR/Tx30WPvzGOcagHcGGSxkL3HEww
K84u8n8fPoVVmNOcvTYi/KXC8uQAbP9lf0bUeiamWQtBAC2Lo8OU9lhN5dXF9Z2j
+EWIV2IZE1gsY/h5GcSi8g7Tqw8bBz+73K91BAJomVPt2IdwysHN5dDAhuifK9GX
syhanLmDEE0bPdvuNHS5CiBsPswiZExi68OlUDVd+OxD2kTE1WjzDAG0rQEWsFKg
4AO2WLRo6cacewv8z/PIfPd6zh5jsEp1gTFzHtETPwN5R3EHPwkp8umpdvL5B5kf
2ATgpbj36YCw2CoKDY8eO+LgLKm+ymPyJHai7F2oJoFHxIQjMBh3pQYlr5tUoig8
yTnBUm6Hcx7tO+7l2Is/seHws2+flADXafiPaS8+Gc3yC2PcV7qM9C4BfgaKbW6Z
dEuQuSFTvIF9aiKk/RqO9GjEs517ygIf35SngARUVDeLjzn1HwiS4hETNoo3rViO
1ZiqCCz14Z4w7LHLCQCjT2AcEWrC3jphvRuWvNEJHiOhcD55n0v7fiVpHVWGOFfB
EFFsbsNuuz4XZAeQFpDecA0S5yySHcVGv+1NK4X8sBkOg6Sm0GexB0To9JOypE00
dtxE/1T3YlVXo+uqKOohxonoBOhijp2mbiIaOxEdGYgGvI9UYcX+wNzxnrC6EQSo
zanIiLpMhsH2owc6gEDxmbAcLvTXHDBbrjoVYm9Ryt7U88Y0iYrvhOJAjsUIO0Ha
pMJkoBP+sCORuLBcvf+mwQ44mAejANT/GaxKp+Eu7Euh2wqq3tVF8DABg2U/WSVn
rlHn7CGuaOV41bBZojyflZqJjLIGcfngk/gljVDhAhnsdnrOHhCHuhMCZQK3BffX
x3NgsnDPboWIWsJjvfSj8ZoFhe+X9/VVCVA2dlmRuJ8KEO8c09qhZGGkN6H4nWRC
ZW7GyjWHoX4tIAu6GHjowATfjfNAPpujw7qUBztslNlU2FlR/cn8T5GKuhdUDdlg
rhxYOKjmDvfVW7wREaHGCr2YpXUkpce1iiJ98NDUKNszOmTBGHNyObQwIdgjM5PB
OxyJNGjrppVsGgoq4VA0tpiGnpL33boJw1rxsMmO1S3kxa47RuA0iWSUFQKqdR7v
INY3l5KEGeYMr+pH1Ejru3+ZF300aK3fQp+mRdwfPHb3obtUBbP61hkrEIcJ9zve
BRcGEPaqSHpk7McauPEMeGnNLogrL/UTwUcIXgL+PrMQ8LGHIVS9yvArBF5VKqoT
r+f99Xsxkr57vZ8GkGtJsqiUZcqgDBdWMZI+fO77PvDjcW3skJjLAKJcWhR1mPVn
H1aXqRrCYlZYTB+PK+eZDqNWnkh7XFwURBZgjxL+NNvwuSTJqRohTB6e+M/oKFer
jZyCFzJD+ZtH2hJZcP/vXgGxzLD7RIqF3yGOjsMgxYdzZ/UdRuH1WtA62iUjUSPg
hBABZV7RGBPkMv3uFrvF3zeQIZFyi4200wxlbNXyscn0QOFVRGRlpaBeS3F/y8PK
SsaXF8E9KAYXTFRiH1kBHabuGIvjN4JXzqlGptOcCpNBmD4WX34vqlnpsjMe+6pd
sg9hFAEputwycLX872PYsHPBeSwiJYoMAm6W5OlBGVg8DGOvkgexYGrfi0gXjV2A
nuyKDHM+dh1/oHm0h2/JK4t2/V2O/lz41zBY3WYvYFfrValCJTE7nfBb0kwSRKY6
24p8syfNyT1Uk9MwIf4rkSfBRJezxsro3doEjO7WTgNQz2kMo7Jrm5IjXlrvMGTs
YWKWwzYXHAY+akec9UtMx0xY+5gAb6Iy2/6jH3W/nctNwejkI+Fq7eo8J17MUvTW
s+S2KNTEQ1/vTvS0Bm+a+/GVgDMD8/w44JwhY0toTerGvjltMoF5EW92LorwYj45
E1GgUqgceK+Qx+tINjZIZ+wlKtHW0FdzjWAJbtnU+TrBBrZLbJ5hNj1yv4TtgQvK
sjGLh2CJnlvpDEnRaMq6UKNO0idlTSJLf/b4dh1+0+ZsitTHkZQaZDJQAa7QQFnl
B0dbc7VdG2v17jFs1JdKx5kOupiIhrw1QUquyAnIhrgtVcwROyym3E/UpipG7FBx
Fzr9+KD3aSk1yooYxlq8qPV405qXDwcHYsOdbQWM6bgzq9uLXeYIQHjz5UEgCdcV
JNVdZQdfhCZFnqlns/gRwHGjqvtCqq4RgAsCtidPWXkHXsa2YdXZA1cnh0gg2V4Y
84gUbSUS6NEwRVvCt8sNHfL2VEQ0ESOws3nTwp72B3rUOLZ/l8MOxj9VKbu3zOZS
T+Fg1iWXbe/4/rU1JjvY+ttDU4H3P5+a2yN+JfpU59352K/prslQgu+aUkNssQn5
q3ov4U9rq7G903NeQ/4LYZCEFE2HzYPbupfcRPhomJO8llQA8NA6sScRD1GzLOKg
0jLbzI20mSRhQ1nDMp9tfasYO6nhu2Q+2DIkjks3g3/H/dUoEa89+yW1L5whDwsa
RV6A88l5Pm084dzn0xxQNy6oj0t5gcDBdJ839FbRkWQM+pWqJGgj1nAtqBMT0GMe
i/A3OH8pD/W6BeR15f3duCW2IIrB8FaKlTOW5zLer8LNSQrZDPdgjoBDGrg9JLFo
d///D5p/lGjizHUM4Riyf1MVrP3ogJ599o+mKxC8CSLJPXeOKGJ09CJWm8ZeDp8f
jUBA8ld3l3QygKp30JhjiBtR4/ByVq4WkFF8zw6u6fr49hYUyRP6B1IfUzVDEqTh
Y/qg3B2y40Av7FHTl6IY2bbH8YTMMT5jq93v4B2u/SFrRIeznEj3lOKbpFX3gqJP
wtszUF2R7UnjYTP5v2YpSBfLhdoR8UzJbmRtpwbl2m0OEBBX2V13FlwZVcgK+huc
sXyNL4SrlkCvcvXU+iy5MVENHi84ngoOAGoEo6m7vhSbG41cqU3J9r0FCOrZxd/t
4WD80QnABdJy1a+ji2D1BXlOxHYW1yfUBtTm5uNR7KxJFSe4QG59MlGptRcOhTmp
Vfah5s0Rgb03pRvjfU5/E/CuchudLPy2PzbgPF+el+mBUFOB5dG5p2iZIkDg1Ky0
qVj0XTWczHdbmUtGy7Nu04UvkZflq1n6gOE+0ajXytB5b347zmDBO3RSLtaYfkPf
XFLp/nLzjitk+LFOr29LDvRe3kCKK4l9dHgDiM667fPZ7pgYD8ofp7AIXLxP3lfe
HrKySiNlCvIFCHmBVDAdjfj0he8d5TCz/v9dkVrpFMTmjxERCWjsq2wbct62+gtD
2cHnDHzEfYdgIW7jimk/GDrQHuKl53gCmXvAlyeoqB/rkKIEaJXsbj7WpYY0utdE
FxdEwj63vVDqiudIzrJum0gGxS2oAlVZHD9vimZfJitWbmAzfcQ0juKvrS3tY/V3
Qq9A6OVbd0CLEssVuaWnr57BGZ6Op3DJW/+oQEw4yu71lHm2hms4bNxQ431riFD+
rc4APD+19P2//jwIaW4kTeyx9xqydd05nLw1uYqY6vn9Tqb/8LbMNKPv82XGQWHU
/gVIDveznrt0KqvycXFassiY1XA1WxK5H3JlC8i2RUXixBxfkLpZue48fp4dFMwG
7poMRtla56kLwbA+4TqLsA5VrOWUpVWhGx7XGiZma3jvMb4RSaUSTLXpe30+8Nmt
So++zgAFIOhiVUN5RFWPfLpncSDvoH7WNMAdDG48zirsh5Y7lBTMWXJ1kVnFHnKE
vPk43ioivrfWpKFK6WT3p5V85yY280lZ6W2yU4eE/id9t5xpDyzd7lr8BDZsgc4t
e10ly3lAYD9i82dvE2Z2/AjTrruTpjMEy4XtOKryYIWV1yM2f4HDttdCc4MQQGDo
itFdv/i324P7xsfnl0PBoTwaMXU74IVrlznbP7zZ7faC7JxhOhB+SSptpu4+kKap
pislE0NJ6fr11wz3WOE3NNYTA1jc1puGeyqSKvtgZD30/5yz7aGFElTDlBnetbRK
TXCSSRetMbwWxU6kDpRkxN3nh6h3gK/G035vTDTxAUv4DGlntRwMZVHiWimSJIF9
jJegvRmrQEAejkT6iP/CGs34imk1R0QHadtfZFd9tNeBkvNFHP4mFhCTPdhplzrc
GWGmHcjMFojLzEETe8IGpNpT0bo6/DNe7yv90ICGqR4mdjYf8c6uj9p0noJCaXto
QuHugom6/Qa8bmQVk7LOBsvihpiYlbp6sZ4dF+Rja6/5holjkJKkMi95gwEPS0df
4GFiuS85wfM087VVEhRVsl7BI0xLPNLtKpljdjafgUpyxQiRWqbaL7fv3os/NhBQ
i9CXdSVMHE/J6RI6RQxvzNGOGQFAKLob4+EIsJ7A8PgH3485PsbthqQY6TOy0JWQ
j0pYpPJinl+bqi4lQ9VydDIMaHV7RKc5ohBPZLVcpa+bLkableVNjhGkbD1WroiG
CigSC9i5GUUwcpA0eGtbusyXM8bPOpwahulFb/g3pPQuxjpgVZmisH3JOuaHbrVZ
kigbrieEZF9gbXhMKsMIYGP3Q3TYJwtKKgLkjEGfJ5devwwyTdIMLT5/PIHzYXM1
d5IOSRTUuddxj9+hG6Swl6++x2CloWNS8s5UCyJBetxaDuISdoU9WbZkztgCjG1t
rLyuF082Lf/UXBa0JK9Z2YW3gFDvBnYQOUchQ40Q8LFiROGDfidHGt8wEbBUd47W
8hLsedMOC7/97XPqf6xZ7y1pkpCCb1avCjA6VldwTS9aO/BG7wOdVpjeZrTY+d3E
94O5LEkoA4FPV6mPko/ywhlALbuS7opQZkOe3eIHIWPH3KNxc4sQlIAyKjpXmN/N
sVZY24UhUJbe6oMH3rmUmqD8QD0nYvUHjA+3rCM56+HxZWSi77zjCTIc0dW1EE2h
MlojHNv82kkqd+CBnokO3fNBD2WP64nwrc6rsiZhvVhnXaVsILW2liLuQ1u7Vpo1
IDJQEXb7j0LLMhWySaCzuhPA0EWfqmWNix0xoaR460XScE4TzmFOrenyuURXbTnb
KdWNeprC0BGy72hxTt1o7rIc0ZWC0uTDlpTKM8VGExXKanhgZ2Tk1KZBd96iub6o
M14pZOWKKn2udemgKVOd5WlpBSmwjLLUjGE3vXnGNXqD/iNFzF+EqDKFddbaOh5E
zaHVzVt4StYnnEoaa46TjqUSo6mzveXsGJtocF7TaTAgdWkDLEyon5Oo1auEP/8Y
n2PpBI1DMQu9xjZBFzwikxEVLag+KoOyXdQUSH2ecBwma9dhzDgoHKidlVl1ncSv
2ByvoUh/rXf2+MUd10fOVCdImW/GDjezGgueE6rkEGcubkMAZrhU86mJp9IcQNvh
B8wstMD1e96Em2cQLPrkc4mkg4yPnOcEp1UT2lmd3RhX+d61lN28Z16a8ARce0+a
mSs0KUJV2Pk404NogPLBRtUUeyyZpq9n3zPxIg5z95FuMl/15O6NtwcUUpZEkUWI
/QyHg90l+d1yMm6Al6PBeC+z2hz7jM57CXzaxZia9i5nMnUDhqyQkdYKf0mtj7rV
b4N6JX/2Jgf28yrpgnYE8gqfV5K4IXzj0/YAOFif2CJmx6mSkahF6GNV6k1DJg+V
A/KMm6z0n36vF0oHckvt+EPX/1ezNN5Lo+RMYKU4T0g0iBA+chygavqoqEd8XI70
D7nV3fvOpeIkPZhdpDaJogdX490jUJL0DRZwfEeeOGK7IFoBudrQVB3NbtJfgYy8
YJs5xUz/VY3Lf2UtBL9LUMNKcCzowKUj1/3zT9AB+g4Jefr9ufv+CzvIC9f12Rm9
3W/OoLiYKo27rBZ3xctpEx1/AHxV0A0YcOv8MPFnBB/DdwoJjaBSK+JvoDG05lu9
G+dyrS+ho2w7kE1qqnNowTlRDNIxmuPMBKjXqlpLyeYLdLkGjSydeeJnPz3O1Kjz
LDwQurf526zRaYnh7C6SDgbQNy1wyMGwm5NxiSSnuI4VRs25jGD/vx3IQDOYkW3V
hGDGcgyfCDmOJHaZRlJexBfEffqYLhSDUfXtvm9X1/9jQovqtrlW7r+CPFxPQKJs
hkIDVNmz7CmRVxGtaiIOAtCVWfu64R/w6CX+eSIiuzOw4jUa4cBsltzqsKpHq1LG
KQZGyu4IR3K7zcn5oWWMVea2VnK0i1wWEArRiUBp/xw91lMk7HiSoO8vpt9vihod
7RuDqUOSUs8swMSjT/4PF59FZ2gCf6g4Mzwq5pKnjiaNj6PzCCyRNhLiSkRZnDgW
/+tz3+3IY0of6WMORlLoabCiol3dzr9AxqnsYWNI5SDg7vhuZaRc+c4NlY0xlEd1
DYC+W1mLzSSgcAMOZRRGNAtOX+CnuVBSJxLr3om9ylti6HFyCdNcz9MBYqQH9ayx
dSMsVgh12I+OON0F6fzHsZASdqCDFXR/itBmArJjX56uEK/iv2GyTbTe9d/m+1Sj
synl7bsW8C45HfnKeKGBlqs01z6OEu5j/+BaSqfUARQTgI/nWzVkEzYmkB1zFoz/
SLgUA5h1MTZ/wzzLZXu5vHKt/GbKHWS94i36VS7VHRgjzJCS//Aw/50VuvMgVurE
N7guM6+8oC9Z5ujZaY5THbT8ZQW9y3DTgPkHuyZ5rVuxeDCXx3583KR+iVTKN+St
+PcOKLhQWLtP8/EHZ/CODSFqkiZ1Ufxxi0k/GyCIoePtBnyH6EnQ057ZihpqRPaC
/XjbX+ydQMU5OQhYj0r+j66i2qEK3XCFQ5oZ+64oH68/G5H9AXxeuNyHrjLVMSHG
jX6fCe0JIv348IPTWMolOYFJ5gawF2ptRRyiL+KLjII7+MaFtaPy0TpI8K0G/0gb
oEIxSrze/kxUsyWRmirOVeCfEjbmPzDfJ5FRo9PO3R34lrHI3hCAmpb25+7xPbto
jWqwLA4Q3YBbrSz1ISOontpD0xPo8Kikc/TsXuvOmXl9m8/vi/3f1IHSbkQ/FWQR
A4uTmmjRs1K56z9/ZXdFd5nolvMcyewE/cWbW1VGiwkvWc4ee5Di7l3uZ3EHa5Jf
ux51bT4tpHQVY4C64vRIJ3mhbKkFcFdmKjc3IZZ2Rq2KhMs2wO0Fn44GAPEquF+l
JsfbKa7BoieyfqnrodMw5pILHI0FZiSJ79XLVT2lNegcHvgnDAPCTdCC8ETl4PMA
x9jvz50cf3KDDyrw8TMFjvP+NjI9wkSAdy8bwEGV8KA2j6AOmpHdm6SMSncp/1Ss
DW5ZnZ5bGHGl9VHtdVGkLPIDAaYzBrN8SHc5TV46a++gVroo5CCqZqTEQ1lZzrRa
lrf2vofBe1m5qMiWbVnxIRtml+7vgSTRaS5TgW9jmB2VYOhsK433Ez/g3szLJ5iV
H24yEDi1NjAEgYRBGCzPJqSpa1ElMPPPsI5XQrHgYmCeGt9Oex8nmjMgtZsNTlWw
wyMrhs9ePSFSdrx5iHqATGUfV19HWEHFvVatKhaVc4jLvis9bAoD0C+PMzhD3+WR
GO30/8z3dpCLxsgNwMjsyZtlsDXmxceZuEh9Yigv73NX0/VlkvVEz3kxxVlmrl6W
r4uRjvb52Quv1x8i9wOYx6j+iHkHzMfAK0D1qH3GUGL+FcaEqd3RZkjpZo/Gy1st
cJTLzwCylBMYyj7SQ0USGMkAlG0B7jPWxhz1ul0uZkX1kXUz6w+wQvemrYGpXSkH
gJQCj+U1MWHdfHzasG3lmBtKIq7r5Ej94T2QvahvDPdm5FZfzWK30DVKhK729ozO
8YZafK1AEO9z5NC91SdINEWQGsUPVcPuUOsp5eGJk5/0YG8mVyqnsv2EoCB9ToCh
iE7+Rt3HQWwtKAUw21okDd/WuUGcgRgRKzrSFstJOrXFtQoW0sAEHOOX+KTFSTQJ
B3Dibf7qbNuiScbMpWRby38xzlU1hCs0beK59Wj/fSC/D4+YpkttwOjIB+AYAu8S
P3Y6tfdRIuuri/q+aQsdNnBiUPY8bXDz+/YrSKxbKfzyJwd+EPnxA9YVBhcr1BrN
fUjiAv1sk3HIsqNw663/PmBNrHvu+fLyURCxGmpkQcSdKBkAVIS0zSiMMqusukxz
c9/MMLgP3YohwHgOwOKzdrWtgGli0D+ipz5kcDUsIQdC4AU5GjLRygeA26OYnn38
yCSaKunS+9xn3rHKI9nU3k3ID6zRJ2PvaANBap+BhSTGRpayG0cK+wyp8zVImx6x
uU8bg4KXB6NuPSxMB4H4ao17nx7n914aZkZ3oN0g0zW8VGfFzuNjdZWPa+8CRPgp
IYyRUuDow5k97WwVOrYuGiMeL5IZRdj+dkVOG8GcpfEiAjI54IiQoKsLix6NVWLb
i1V1LpIGV6pc3FyCFQG31wTTY+U72NTUVycafeGcQB/RIy4sqgrdgInpn2oEC6i5
Py/eSPFKGoQwCjMP2CtQqgfRImGTRrQKHLj17tkH27cNfiiyi2hbs6P/SlKCNRC4
37KbeRHjsQRwDOeabNTIctxSlckf6ryXIRz+Anm0512Oa/jg4gisqdyE8vjImPqm
FpkxKNEvXqQqentwpxS29jVlKlcDdA4TRD1oTprbxVbGhew3xb8/JUkYG11MJiZ7
F/PmOGaP4pxLb66hoeZZe4x45lS+bvt5JkLSC3ceZ4ub+1vxWPth6ZgjJyEEhpIj
UbUxZK5PEcX+5fDXIQRqMghSBh3HAVTkgJ1eTCJc2806mBDIQ+hUIhaYP9moXy57
noNuiL+qLDB1pmWqHGhCkJzpiQR4uqDFzqb7dcDLuFvEa8el/MFV0khktKygAN40
Vkie4lNFL+WLcM50LYmFC79I2JgX+h9psYJ1VnfT8dzQk3SZW+UOnooHZztpOlvJ
01CiHNwIWPffoPFND09m+5YmlvkQi43h5LHMHHE+/R279UGkOdj3LwUsDMrQslDO
TNsYsW+Ckl319iH3M9esKGaURYb/yI8EChE649CYK3oRRXo8BNmdMo1m92nYcj4M
M+0fOWyhvTfGsD5EzZDMdqZZTR6wwkvyCpRO1p8tpUeS6dCXZjDol06aDtdWjkqA
XG4xlPmRKM4t5srvUpBr+lCC+l47OZzuTpa5t7tZtQiiFvkn4bILaaHCL6sOi/FJ
O7ipkxkPwBMAMWAFCl41+07n0iq6f06wMmqYoNxqHFsXa3wtAGtRIvc9nUV+ZBQr
CaRmzzk49bnKhFGATmWFvnEBtUKLjvXtwA/Xewn4UPQIJSOPs3WGUE2SwHivYCS0
N7HHvwzAy0Pi0IP9Dns6HlDeLD+SclNl9zYVICB2lSUBR5KoXv+WKymJYMfDx/iK
xzzhGd0hs4CCMuMkMfasQDTt1S09CiwIlOH1/5R5tNTLN9dm5xgJBJRc50bE2KbF
tm+91oro+oyPMq8ZHhrZkoAaSYxV1MhTrYrkufv442z2ITFLMKdDYizc9Ooqqh/O
BFn/WejgdPvclnWmX8Kp1ezJrdNsrwrYuySoVsxJk/jSk4a6nnhRB9wHem94BI6J
fODdoLkLAiWvZfWUT0RpfQORTC8KNHIlE7SNPI3mkWY+vDazPf289jk96ajwKC80
+O6dA1WUSt51sRPgNgYvzT6+r8ukQK3c6Pg4nphe5l2g5WthPntbEH24rQTNZb4h
hs8rY3siADXyjGAEx2Uz3XlNz5KqP/Gm3qQZDQIHjVGAvT5iabpHCZTOq7KA7n++
zeh53jxNIM9UaW3IlZdc8TuNRQlPpvswGMVJXWhn7+rgara73Wqv6MdYq9NBLfaX
xqhZ8obWhlh72Ips/ir10ZQsQq1sEcdLSwwnY3m1y6yMa28SVM0cr8L/CccNuU0t
Su7Aof/G0kpa3mDnDrOo++sGy01FiFPj40RKr715RZvaGOWy7FZtdR1Ot4As8fhY
qMPo6pHRmqgMLoz7snTFh4keLt66zL+TWUNjWh94adXcpNL49bpI+Z1GphbeCbhh
qXLC8osRwUUMLIXTEAb/RFKqlpMqHqP9pHVioXii8S1ciM3QbHQ8xbU0FfHdwOb6
QattIxj87m6LW48/iXT7x5jUkuNQoeLAFc8rnsYRRRefV801seS0CCBu6x2TYEz4
b+sbNgcx0FCQrCVPqZGWIuaJcgpHb/oOEUkCR00QyBLhmlp6wxVY2GnShOS+EJUO
fbEas/zM4xlnBdB3y7dIO4n8N5A37N1t15EdzWpgV5VdHIY28iEUg6zHXTW+OvBB
Mb5upb2B6Krnmojq+rKMSS0DE8i44jBB3VShrpTl+qvsXX8a2lG0SMLQnaA3WHB2
EnkyVm8pnePE6tj14ZQTCsA0aNbMLrsxxrMwrBCv6EPPB3p5uf+tHzvoAXzidxrp
O3DkY84/cF8bACkZTopVQiul/DByHNYXnuIHEtZotKlyqfxS18cJ1qJMObNO/95v
69rbBpLYpKccwpluz2s084eL53mq2KY+JuDI8u4SueWrSRWD/JPZFBmGesm3oNpe
xSs4gFikAACWNnRD8G/ARTtNWrHAsuj/ge4kMKa7wX/nlYD2WAxK3wCzaL+0e0is
jboj/JKAH6ciACqRFU+2fYBW6LlxyfAwmaupHl37pFBf/WC5o/r5gllB27sfIffc
Ii45wneK1EaL6u5F2NR7T76bimsRJ3r10N+a6tPRZq3pkUtQZn2g9+gRrEPySNuI
bEb4O+c9c9jO3Fo8B6eeZSFeNc0jhXwblX22VsUpU4bfEbeODP69KIiId8o7n7aU
9SCnQGJaTKJeBsdaQS4iHvSFdjTfkG8VFtuM6FVOTishgkQpfQhQ7yshe5chgBXS
bpXp0kozzsEBlFiDH+QHqXSg8Z9R5H72Ng7wTGx9zw5FidiHRqi3Kbto6ZlYtepL
ryeUz2U9vQcaxA8KoA8dJJXOzeNW/xtcOUJf/tsrEmDwj1b9opuj1jKdlmnfYmoZ
s/YThkrK6pGZvNokJBJtGq/PEx6zxaPayAjSaopjToYMfZgLtJ59iXbbMcSfdItO
chNpNs+ukk2nG0/3JCz0IO3fw7nT8e0Ep3PO85L06p9UzrR129TssriJzCaqbWm3
6Z/wKW+4Ft6JZVdKhiFA4ff+fjBWz+g1b6WHnm1rEVVer9lf5acu6MM7iRaATkmo
8Urnee6Oi/TQWNQ9u+73dGfEQoYYxIB1iktLRXOVZnih9qRGaGsdREsmJcC1qYGh
pIajAq8DxoUZsYN3E3iPVMG0GN/4A+x0EGBr0l34hQXqstZhEBFqmylpByOkTHEd
HA2IWqJVbUWa1FtFREhzkdtdb//dkf9wHJ2lMxEw6VoW68EgnxIB+u8w28x9dwI4
TyJKDP/DlL52/l93esX+Rn/3JKAvzJMsjhRSql2Syoro7QvDPrx0qWhejCt3ejRf
sR3U7pD/6FBa0fvzAumFXifiuAunkEFkhQkAp0z9bS8flopVrhO1spYH45Ai6pQS
YvR0j1SzmVp+7oI7OwwWZ0gBpZuf1VWSTY1tibk//DTecawLp+YXRFtjTTqSteu9
RZYmVPrJip9WlZyDfzh2s/GR+PlPl0aLqpwkZa3HJ6RcDFvXIswzK8sibo87lauz
YfA3JZ8bZW8WmqC6iJwlYFKXST803H5glnzeipngLRu6hu5q8s9KkusvuvhZABs+
YMPsH6anccFXbH2Qr7ICjSiy4EWOzX0XL0tDMNuTCYlu3a1lDhvAK+DFT6oZaII5
ILLX0Lf9FLxH0ddQ4yfG+a+VEcFjwy783K4SucmPbebcKiPcnrRnta62JVVvfMHx
7tkJ6W2qATotUB15romdxGksvrBSJr5UaPQw0dic5I7m9523a7YzbTkN5bUB/r1w
UpiEZ1VK+zbE6Qe0e6P8bkJlleb/Ppk7zd6x+guAgdXUgyBItSgOECifIFIhUCJU
WDF2/0sOPAJn2D1d/tQyVsCSE7yqVryr3PLo+OhgmdKoEX0nzB4xDW1cQ67V4Blm
QEyttpX3hbJv9LXK/Wimja6BOFWLAbkQhz82/ise1xZTFOmH5/BXp4siz8tc2kny
MaAMb3ccuEGLgLM/oyH8djFNak/udMt3IDJ4ldtM5m+DQbyCFSXS+RDG2VVWg4Sx
WoOiC1KfwoX3oIt/UKnsuA==
`protect END_PROTECTED
