`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
H5Rp2vgeTYlMNdl5DsZ1eMFkPPADu3HpQni0N98Q1cmrMfYt66MvOuZKx0k6Za/W
SnKGEwcLIRabFTxT2m+mJVpJrjhSWl6VV6fmvC6oC8wJzupucJqfmO3cdwa5sCVI
eEw3hD579P8ZDmRWTyQWe9zUk5lViFo4L9sTeSAkIUHXv+KGJDbwa4NsLl1aH+VI
`protect END_PROTECTED
