`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
f11uP3tAS38J+2XEq2c6cCXqulsLlcNL6TyIPPAS8YOeeWfpncWiNfLmLJxSx2xB
ybMBixzl+R8d3+94DXpweZZNCfUwC2LXdhU9WYyBbAP+UuuTzmlI2Y1n8DqIRxnh
l4P06cdQ6lJ2Li/E3SiItrQYG/U2s8cHm4No6Ut62S0FMc9Sjk6zfi4dU8KuL7v7
`protect END_PROTECTED
