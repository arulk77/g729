`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN5WjeAc4TE0COKFJ3A/FFNEVrgZorq5YF1EG17/Q5Xx9
qmKsT47rW+EUOmBjQTCHOKVHo6FpERyJHc4u+0qo31jHq4QXF825pFne72GKC4+u
CrhdOOL8bwANYPXPy9zCF/XdYqIrZlnFGBoOGIilHSjkFMwqE3+HTUiUr1LDo84b
hpQeRhxTY2Kp4ZfqwCosg/zTdGvPwyO7p1y/OZ7kgqsuk8BNrfJ+teOUpvc+p58Z
QbBrmDaQBZ8/C/ypQ5f0uEMUIijA6fQTKdogZ7Cvyl6ekdf9N8RHoSH94K7GJa18
AdJeXRS7DEi/fbb8gqoUvHK4mJfULXXttFtYlEXHv8B7bkE9rN6Bh+7sglFAtqDz
ewAsNOkM1tDY/C5vP5gZilUXPoC4GpmDIlLodyAcBvsZ1nCP0aeMIAX9OMRc7CwM
rRROy2wDKMXy/Snxvb3P0pYrzAbj0RzP6jO6/gBhZjrUUylhyHHFgNMF/qajd0O6
z3t3I+xDOtPWwj+zaiOyUEKyaXRVPSxyk2c6ewDk7UbYDrXhmlow4xFVeg2jm8Ss
JYBpBZsN0k4pYmkIFNHwRhgV5wHMN9fLHASfY1CQ680nGYnl7zZ+l+OvJ+CZ7z/V
E0SUbYnx3hTFUEHmPp99J0oUfxsISN3fADKjvNW67hP06PDwpRiUlD3eqCvEd7JT
GOzuTAxxWhPXmtQ157AFG4HiIGYB4q7WhFQw0azo8YTm1DA7H8XLsgpVpNDq0V37
6p6dHy3ttGOWYK+cFbRzVNBOxrJ5b/9x5YYSWzF+uuAlxWOkqEXYW3ACwVFvMSoD
gE/OMuh63CU+JVGoMXZnDEdT5s2b1oS7QMJUXJb/77bjxS6FK+/1Ler/YoZJiBnM
FzL10sOYonBmc7/XhRJqFEuxFTrm14msDnJASHwNggLXnChdopMfSu2pVTpaKNJb
o5+oZGQg1M2L3rymqH1mo/mecuLLVbc+BriiDOxg9/rcJxRg0SclXGCbMC0DOOfy
FdpF1yUkoS++ns4GgWEc6H2Axv7NRtWS0IHjHSquIF8DiTdjCJpKipFlZoBg3r7O
j7nnF4UiCkpxjVXDxDBSes8JJPvnyNDjhfAmZHTDSWs=
`protect END_PROTECTED
