`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C7dl/ZwabBouUfg/CMBCp7TXDqGNYpoyeF+Dhyawrafb
LauR8j6X9TyNRL79L/EI6RqoktThpSNalVHiAiusS9pCHiSBQIeoLtUSnN7qBanc
Vf5ggCbLJBpynaOS6bBpioNKQZPBm14+9ZbUVy4xzyzN/VBIw6eoRMLzK/EYa6+u
Lqbdu0grLKqKLqenWGQvkdkxXGz0fKcu/XpLYqhVMqtl72MvUNh2UzN0bV1zPr5v
YTKJPvaf3ncg3bh/GFdtJiOxwQD6Xje/uQgbbv9/NKp+DUKq0Q0zaV9FvXn5G7+S
sRCJPtsRyyXWC82mfdXzaXMhYTQ2vf1HT++VvCzOG3T8Li0DL0bnNtLALSoZs65K
998GpmmEMqGNjRUjyj6CTbfpspMAZ4gbf8vXzsMHC8RovkPb6nT+wbu7xjDKB5tC
JeL7C6aPmQzsBDyfZ5J8ODLTJfocO437o9Ur1uVzdl8djeQP+zZewiXsqy21PTKa
lRP+u8lUL4F/AIrrkVm++gQ0LLUlgSepBC1jwebMnCn1Izp1ddGY7jKCx7Yw0pkd
bR/j9gtwRZVOzVqc1Y6HJgv9Xu5iATmcTDpn9rP79TVEn+kbXGXQ+4cbifXe3mos
Rg0wN/oQsb6QBou7FIRAEdDxy3VuS5iP3P5jlFpPfM1AIITs9y9La/ierFzR/B1X
zWfdYvJCLiinxFMSy1n6CGXywyZcqrniLduuyCLzKpc1ZAAftMwKF7Ji/okDt12x
tbecRx/rHgq04S1BA6uozDBrxpbTjs7KmMeaFyzyIYRn2zENkw1QaBZsehQkT9vR
rQGNwaSqmh0T4bLz7siZEPD+tmHVQGN6PfmsxgE78pVB9hRfTlxdYhV2biQ2WAbS
V4f4iDXVDURHoK1fUMmPk1OFN3sws5QyW+rXUy9p80Q1l7wEN07PFkFYBhSPegXQ
yN5c1QQ8M/iuk6Ja1MijNG2SC0dVRYs5VqJnFlF1ufEISseqaFir2AQzDidPuxIv
XNwhIeh1X73RSe3e8/iPq21uDJjojIvzycqAr/wm7WpBJRaAsnUvz3PV65dbryGR
ZC2YVT2RUOhF3Qg6aEOEclAmDXfO5d77aBtWpbyCILvEwMKZ+koNwAe32+PbFwCL
YaCRr+eaq/dOkQPzT3pHCimPgX6nu9SZcCieYs8e52BB+NqDsp7LNMMuLA5yS/w0
4i1bT+b9x7xC7XM9/NmHCfm0todUxzx12fcg80eLjngzp9N1PtQ2MUcvzwIsoC/c
Z9uBpsykN+YeEtjmZrZqvPypgfx5Uq39ugw7RT1l62lAtjonZQiGYriCA19Azok1
7KFx8xqjDS7RRw1/V0ZCrv2cWW0FC2fK3sH1U73tv0QfwGPqZvLzFaeiTBG7hIht
jomy8ZxqTkikvLvKsjDVo3IryuTixxoVEnhUAIYA7qulv21H2WQnKX5wAeJzEjK/
0lY5yRL+ZaphzQsNgSQuq9UabK9V9hO3rZbyC22hDBPY7UNajyPetjqC6uMhnF9w
pZd4/8nErUEj/6ShPWRmcE/NNx0jdtqXTO2KFO8d5SxaLY8VHuSSesvY2uJYCCNt
yS/Rw+IQ8c0V3nGmNnyWx+zosQXuTWghcLSBm11B/VCxmEv2JgQ4CLFNwe9VL/5i
FP1sH1lUV/h5AZ2E2jTFFz2Ai40jao01BMnYnjYm3sXxIonHw6g0DbGd3VYKiw7c
DSGaCE9kMyLjgUWBh9FYg5SiB1AtqTQaJkoYBoCXkiWhlQym22T1m6ztMuPJWzzr
j4CXOvjqYgvuz7FJyWjzoafbyiGDKJDOWUROkvX7r+zXZ78kDd0v2qi5t+6uWTuS
LEQfXL2dgAzXX86Ugad0O4ULS0YAXmZKHy9QhEZp4RPO4Dic6H2yN0Y7pSzx4GDf
RX4obn9iADMEO/pFJEcog2+hJrKPo6o8QSG6X47FWPPF7gpOW1N0E8zBDTkOOPEj
nzcR5KqcyAjrDSLmRoaOE/LVfgeCpaeu9xt26JW9VTSgQnvDRBFZAe3dbnz6smrI
FRcfzuIz84sD5n0GAwygW+s1ueL4KK66DeaLkvN9da/BRbdOJsCsleR8adET84Kk
QIvU87mPqI4tBeWt6CN2jra+7Xn4IhPI5emRK51qbeSHr7b+kjukK4vVNhWgpJ70
uuk9zKyR+aZZtwtxBWAzcWtZIkLKHVX8DTwNRuPKOacNO4F+/4ryXm5QxdnJ7eaN
3TJ8Le4+UkkCpFN3L3H6yvzIPnl00xCKD6hQ+HTrXG68UtGOhBAAFy46iWHrAU+1
LfuURtSEHCGrV+K4Suky7QQ4ZM7Et8Mhxnm82gab20sSGc7HtGkQShLbV/R0Emhb
vrEpmNfIRZKjdDSwoJbA9NkDjui5+mOiviKene/uFIKOa6e63vdEcNcFFRXaL2EG
w2BA7CMx3SeSx1gQUQsQ69XCy7BIHODFTpWAbkfXrfbv06kCvE/9FgLKbSkI5/vo
uHP2iL4gXu88j2r4QPeavziapPOy0orpAVH4JJMxFrZ1fEtgcJbMBItXU1H6nn/9
Er+Bz1Vrgi7pywp/Bki0tvnw4dpbVvistPPSm48OZ6ek/CgBD5OXHnuC34sQGFgx
bZMd1tnOszbZ2+xxx0Lb4twR60BqzXPRBdVzT8DyAoHGXr3jMEeAO3CS0eKqljBb
UZhcjfq9culjA0CgvXA56F+iFfUcjZXBnfMGvZrgixVuoWUGrDqDo0CykHrIUO0F
IHanBvywMTNiEkPz0LFJMYjI5yy0bXGmOE+oX8Oe/5Qt2eK3ny4D9KysKSI/PWfI
asWcG7h0jQSS+nvlduMH0BB5onI+Sf7zAfKYjjDKGklVEOuhUKjQ40WmjJFTQIjV
HOBl3xH4aGlXMcxfhpOqaS9PoSEXwQ7c3PFKWGAtUSGiCmcmVcmU0kdYr0yT3gfH
y2TR6nG2kMQ8ZCprCT3Ad53cVr0DxcDdCJZ/y4kFCjKu5a4i6dcGXv+DWh/f3Wmm
nmm6X83GqTC934KCW0CLs1nb8XLa7WIuskkkkmVABvEN0l2lPderLBcvXpfeQjJD
topB2CzZPWRUj7jBZumSKFvR2CcDm6sVlZiKnZxf42vbhzJ/BkIYQ32A+d59Z1Sa
7ODF/47zFtQKvLppVcqtPSoVoHzlUX06uWcsLLx4m/SZ0qWOBQ+PwGumCqhSWW1u
8Feqmx7TkVeoxY6cOUk/4LFC49+4E6sYiBdrCvI9gTx2oz9S2pqVOPsQDx4e4BnZ
2fuHaO55B9u9WJ657pZOTR2UKdorFe4J0wSHMLkDWGH2PCfdOUheAFlbe1vu8pH7
7p7isFyHgV9SreGH591cdYquHG7OaHdsaJmPKow1kOlnAw3yatLBolp4hFb1160Z
7lhrES1WbleiASwiRdqCgX7maDgp6gojlEBOFVWDqdKkoO3BO3RJ5GOpSt0tM8aa
wXkZ3YDThdYJSX9ttuo9cUE9EtaaikzQYuEwI/FTfpWfAMgBttCz2YqljYq5iNJm
EjIVvpHNBbzpTRrIlQpyb/D3v09y3tfafdSNJ1kIRbTEx2G8O1gTzEpJgO7GQ5E6
hg5R0FBZkFtcLU4UOQ0iowdE1750pC91W73NflKyd8e5bozSzBt7y5GbftJKMRfO
5OhQNukt3yaAFmlXP3zGaizr2nhWsTOt8eE2lEmIjA/6TnrPL7p738PPNq2DMPuk
ng1qf6ZBIYrm9V7OLo36z2RVF28dOM96vhMc4UmM5wH7SFAKRQYNDzdZl63b8fSW
mK0GvD4IzRj+MG2tsaap4Go8RuzRKfGeFrtWwHvaUgzvhXMLYYAUBPeGdISi53su
ldH2EPn2YCfLkaxkaBWZarKy8n+nFJPwRP3lPtBzwQQHGi4aXF/jAfUvygJLPTTp
pSKxPViKmgnK1E7iuCvmVsmhLEy1U7AGkUxgDF7RC2vmFvMycl4i8vkfsmNInqAP
KliNX7cXk4SWY2XKbvFESZ+7kcGlGbGGPrs17Fse49n6Exh1TOYDBpdKeB/JxcWT
DhXo6BBvEPA8WLAJKvkAZ4jE4Yf1ztLM7xKB25eAtqevE6VXmivZDWooIwJPHHrq
xM9djsQpg6NNPF+2knFBMCjjtPYTO25ELsiAW2TT5gQ0pY3a1ye0lVCwbri/CS70
L3aEQrUPOSAereX2/G03dbqDl6fkTLpuSpsN+juOu/IwFFahKYSxQx2YSjfuEA8y
IEBtxTL7EcS+co2x/dkKWqJ6xyHMLD+UYuWp+GAQeS7gTq7rV0A9StYxEkgnU5T8
7HZsKYje7jHL85INLgv352Knv2tCiBlDhrNPrAzNizLZWg+Y8bsPpDg+UlkhOq6y
ogjmWg+HOOrzwImrHOXnMMa8zT4joW4uoIVfQYTRAmV+Q91EY1deT0q0LSUuCSFk
+YZwPsFBueAWG7C27vAiaV1CXRTBAwSsgJsz5I/msgVE7ewwaDtWPogRyb2AcBCN
QI15Q9dHJ+ofEk2zq9YCdFbNrEZKvZhuzFmvt3WFUl4sKMStw4UO2/b4DSFrXqyB
inYcPQK6VsImB+Xxi5/BbgKhhLSGaKZxakW0IkSPkSSRzNg2IuWWdirbIm1CyFio
HFNDuZyf05NAEZ6ML3p08iybAJC5iQxtMznYdIjxsZqnsxTuOcAYWKXx+4bZlYd7
9We3yvw0StkIEAaW1DOYDxle6iRi7l7TwTmM90nJKK4nReqyOnEnVDcGt3tA1r8p
UueTXTnGjos16ItMXvz1xw/XBMYJgMMiuMg2GdtIv9n6ZN33STa0xTSdTbaWpVTh
fAv2LcKr/BEHVogXV7dGLTQ8OfmkovMQ/RPskn7XyFmYUTkdjMVPVyQdRAwqmoXh
QgmR9Kw0WGG5k2mcrfFVjJ8BYdImJBRaWNIxo6LBFxLhX0VoCsN54PMm4LBfe1qR
W8rd0dhDPVShxw5ue4GlxrZ/KlvgJxImItUvh1Fnt5ZZ996g3ffRjfu+g6cBOpJV
i6WWribqMsLxwPPEtN1Joad743l+0ZFO5T3eMf8kKpN452ic5f8EnVCm+G/9PmFM
AzYcJfYwWun7ZiV+buyI4dem13LRDCQdxgskPmsGVzhIbyHQwwa++6xBKh0JKpV5
bZz8z4oSZeCa4xm0Yik0iQbODASic0qXwhyPuSuBjnkYs80DrMItx+yeskCHwKmn
slLtIf9OA8h+3vqk1xiSCDSYG3+x1XZVNp0hQ7OoBqBZ6zS3Fu6bYPOKNCNQy0N9
+ZuYJFrxsikceiCxK1qwMuS6UwMzLhPdYg1PA6pftoBS5ilmP12V7eHWTV0rI0r2
XB8r06SMbJcV2AfHMI21m65HlX9u8otJ3N5R32CkyT6A7LOdS4pgM9uoqm/k3tSb
XZwPkp+DnCe2RNYiROxZiyowpFHA5SSwdS0PZeH0P9TEvP901bdfHz8Q3wrjZHt9
63K3ESw87qM2OAHOnqVdHJ/S3lYECkLfkIAmdW4x9Sef3T4ZSpPWROdTAtRzeevD
vq/ZiQpIHH+EQWJmMn0xxbDNtEkKINO2Wh4gKGr++OoSLsIBgtjUHZjkMspMM4Pp
gAXkF7Ws2mh+5ZitQ/bo1L/amad+Z7TGH+Iwq1MXk1Brnl/qf+hfNE1WHpxPL8QS
MrPk5zoChg1myEbweZnNQMea3vwM8JV+9JDMH5BV5BCuHoQPdWzruYyxVyzMD18c
8S9WmGTDyob/0yRbvP+U3KXHKyXFWLvs7M3ZluA//MStV8md2Fzjm0mNXYgD05oA
bbupiqDqvN7a796NJBTJvQctOqtYMtLV8j4rfEaRNpghHJ+a8gVpOlmlVKTb1GN2
KPpTs/crg4gi4hPuCG1UeJ73lP0gavuuc7sX+DvqDBWZlZOLtpwi4oYlP4uOrp3w
dstAlAjuDmBZp2Yb1Puc639RNw7+cnELvHLII5PENBAbwioEUOVRl8HEY6H9MKkB
y7vckXFHiRSMXJbt3Wm/eV6/mRI7+3Ntzpc1WPVgytc82Cm/0Yj0ElqmTlwoPo4M
aRi3AVuMu2CgXKncN5FJESSNyRSGtb5JkYJOfunVD9JrbyDCN8n4wwD2D1YWc+aK
7AEbJt8m9qKgoHHrTHg/RRRBzuJvu79n9IQ92OjRcYyCrtVRdhDxbOzze5Q5ZjGq
eLzwMWoXd6eRdV3OSJ4cZI/35WS23XINfCcACUyuqM1C1vD4ehudgWfwCRmD76UV
cL8yZmWfRqj9jfnpDHk82HoqyQA6Y6SEcPn4VnHoj5ilAeno1laR0CpX3UW7bp5j
xzMbBLnnIBv5p6amT45vYGN+iXzR0QHmvd+74bdXJK9yJap+BKTMaP0xIKqJjNe/
xRsZw9/7KyV4r91BB4Wd3df2xOmSmD4CV305a+PAx5ULJcQmxCMq647H+CVpKy6R
RFZOBn4v2DdipcYCZZ5lM0VcyUMjMa84hcfjWWhPCypHgwhIuebYBmdKw2/1/78u
QwvMGv432UFjPw7JwTkGCPivhiZ10+sYcDcSs0TBFkdYxpAWMfP/+SgM2f56AEbh
cBL7kYVfcrMZ95ET65IzBuWlO/3XfSJOv7uXZePuYle3GY25Gg43RA8trap+koq3
bI7wz8DqG8fW6M9lUcRJeSwxwzhWmGI4aBubNZaJyLmkH1giOXTdzZMzLyM4ZIid
XyjF5M0hgkmo/ic/d46Pdh6YtP43qR3dw6INtDSTdmcd0mi2UtnENgJNPdl4qFxR
Do8rlifiRrUxYBi0Twh70+80Xtsx4mC0GeudQt2lH9JyDjFucfU/P6XtyMaDIiLY
ZlQ7+S7F0sZwih4lyVoJaR3jHIVlAM/w4F3GPJdlDqKT76HMzoTInB+ccXvURvv2
XPFUsVHLOcKjEiWzJn6b3JN8duX/1EtdA67+JoBTnzXnsXUGZj92/kGCHhXfI+v2
FoEBVnPB5im/vzGZSyfK9qSGIamzagb3QF00/JNh3yCLkyswAzoJGC6Pc5Opp+Q0
lwGoRw9MvaKPFSS6xvWhkJlhp36sS8AIm5wJtuTwDgs4B/P1AsxUoNh6R1fsMJIY
IoBcMItkdKIutFQ6zgchTAM3Q6olTThFOKkiFeHCDmlJh1unRVDyoDR6gedTzDlX
098vLpma9NXLu3dh4A6T/oSL5njyIEMsK8jwupyOcADtHlXooStgERD0NM+JpmFF
Nf1ag5Z72sEVj0V+xUk8uCadXDBQ+oWtEmqiJaLmQRzQgtU09us7XPDnly6sn1Oc
k8GYbUlPRUpywpRImooJ5/SLcgGnLSHbzZDi77nNdTWAVm3U6YKTSymsFOdNKktC
SrsLeoUmd5h92eVuPM0Tn3mZeC81ljN2iiZZ1YieQ9KWDUQdlHUOJugbDfz6URYX
6VhtUupnFicUsZJgGkh1m0Rhbmml7AqQTFezA5Qzv8c/k8k2gxbRgOj1n2JpbK14
MIRTkdIF4YW7pwy0ZgQctrSivVPoTlfsKFMk7AW/IMoPfSF/xmVwwXG5OptRdlgt
iUbhQUglsLB2Q3FyD5L/kc4UE+Usu1R9Ivb7H3WLYD7tXGhYUPpUni81pDj4rvf/
6bSiM8Am6NyBv0DmQIqX6y/OXV1bNfQCr1xhBxWffpIX4j4p6rkfsNC6Z60vmmtO
0H+U+952bmZbnpM8BYNCaGfsduBLHPVPWxo/lCWGdPYslaxWcQfSzLYubbdL6f99
39eqDUXo4yJVtyOIJ0+J3P+YHO3uGe4LmIBRNSfbo90Xtdm7ayASuGhyulqhoWf+
EV5OsWOAM57ljfycxQkC/eJSv3VmFluuxvJ+PqjgWmT4SlH9DJVQB7w2dlZy5JaL
rRlg0S95Hugkk38aDJEQN1EtzFwXm1Fek1SeX7970pvwgxAxFMhm9oYoZXmVugYY
Km1YjBRWtVT4Wk0Nd6SWgahw1Rjz7ag5RtGRBBFeRIWtwrTstqsl2YRQy844uD6c
dCWDw4KNdHX4ClvKqldh+hrls40M3PcCP9zMrYBTYhwvfJlmykDjuURvuFkT0/VO
GELzE4vKH7eNcU5iOcmuLLuFBPd0WWmUOiR5lsIHo24GDSKIJzJmT1ncosnnxVY6
ytSkXTSi0I7vvZenVB3sY79KBva5+wbL+V+a6CbvouuJyxE4qDpiJ85j6daXpazM
Ep5VCbqMa39QNEcY3Pj3NSA8NT+/ijzNc8g1hw18DpqZu7XRV1Yuc52lo4SaZWvt
lQv8+hJL7YLEew2KOaSCiTnFA0zVuK/kgcCQx49YYzpkfNaH5gfLUknx1mn7Lp4d
BH4vTHhcHNEZxbl+0/+ZaRsalapDXa57lrBy45SEKruoUwonLWrzDtfETGB06Uhe
2XzTfD/gnbAAtsBbSUepOyTCSV/aA366jaUpmLfkmifaJEuQWaLxk1m9qF8tFezA
`protect END_PROTECTED
