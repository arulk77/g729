`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNku1Odfgr+OiMX6EOrTsae7/YWIqVi+6c2ZgyTk369J
KPcbVc3T/fP73Pp1VuwmEHkr656T7FxGgo6/Yal3cYCVzMWhAsSLbxVp+DPupqBD
GUot1Jd8s/GUdDezSPAFjle+tixhf1Wkd5jB0/mMeqg0X30FNUTCjI3thzuhdwK5
gEAbZ4OC85lVnJrnT69TQcdZJ9P7Ws5CENOAXclFdIpjwul1akmvKi2T+IlqWdRn
`protect END_PROTECTED
