`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHVS5Oj3WuZWTsWbfzrs6NK2BQoPUSdkCmOsS1VJPsfH
wo6a8zpjsJWaVAqzKEcmOe+vCFVRZltqIx1YAA79Sr1zeuNEUWhPIZxcHgF+OM6j
kV8BsmiuEazQrFD2fMDVcdki9CzvznFgtFh4iW/aHuAfpwmZO1vCyI2YAp5APkRN
/buB4WaE05QmPpyGe9ZjPxrS65rlJbLp/oBC3WLuEyyw9g5Cu3Qe2gyz9/cMykoQ
OCt1lySwUfBU/JSMHzj6/6gMEBQ+Y2cVdjVnxt0Zk3zFrjYERR92AZrR1J7Apdbn
7sBYY1SnRlje/CH6XP14u5vu+H0Jf0lYoPUkLOmIo09ncWxwnQb5EIGeNRL8BS9q
Dw5CAHD7+G7+eHkx7bhhUSamRi8aOvompCab5ZLQWpEgk0Kknth07o22gMqUwogW
`protect END_PROTECTED
