`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4ykEq8asqeiZQSZs1eE/O+kreL81vL4E+mUrM4jxd9CM
cu0g8qCo159W08elQ47H9Ui+f2BO5VB+uVlEE9qmcdtW35y2fBMCCwxWl//RTR0z
PjwM8wfKT46wicY8fNUZqd5QEnvC28SJky1Dl9/ezvcfqJilMlnIdkj+NgrwiUZd
sGPVbOPIOsPBszZTUm/QGteGvPWVCY9UUGC6u0PycPv50tMvUyPay97ka9ENT02M
9bY1lx37wSc0EyfPWHfofxM4w6p8+f5+LfAU2IB2r0GOwJbt7c6/xRfRNymvhZuf
+SuYRfbvAdp6uwmp4pUXcZp8e3m9kU6VfypAjIRvQUE5o8As5VZDtFRj2+p+B4of
UoRuWDtIxRVR9cq1f+cfVtchqWuNY+RuYo2dw90Y3BxQP1pmhqbaWZCmiGbATiq/
ZHNes6eLcRb/u1EkccRrhsBIBPIAMJ8Il+2pMsmTO6KphM/8sroMAHUUhv937TXP
`protect END_PROTECTED
