library verilog;
use verilog.vl_types.all;
entity GT11_DUAL is
    generic(
        BANDGAPSEL_A    : string  := "FALSE";
        BANDGAPSEL_B    : string  := "FALSE";
        BIASRESSEL_A    : string  := "FALSE";
        BIASRESSEL_B    : string  := "FALSE";
        CCCB_ARBITRATOR_DISABLE_A: string  := "FALSE";
        CCCB_ARBITRATOR_DISABLE_B: string  := "FALSE";
        CHAN_BOND_MODE_A: string  := "NONE";
        CHAN_BOND_MODE_B: string  := "NONE";
        CHAN_BOND_ONE_SHOT_A: string  := "FALSE";
        CHAN_BOND_ONE_SHOT_B: string  := "FALSE";
        CHAN_BOND_SEQ_1_1_A: integer := 0;
        CHAN_BOND_SEQ_1_1_B: integer := 0;
        CHAN_BOND_SEQ_1_2_A: integer := 0;
        CHAN_BOND_SEQ_1_2_B: integer := 0;
        CHAN_BOND_SEQ_1_3_A: integer := 0;
        CHAN_BOND_SEQ_1_3_B: integer := 0;
        CHAN_BOND_SEQ_1_4_A: integer := 0;
        CHAN_BOND_SEQ_1_4_B: integer := 0;
        CHAN_BOND_SEQ_1_MASK_A: integer := 14;
        CHAN_BOND_SEQ_1_MASK_B: integer := 14;
        CHAN_BOND_SEQ_2_1_A: integer := 0;
        CHAN_BOND_SEQ_2_1_B: integer := 0;
        CHAN_BOND_SEQ_2_2_A: integer := 0;
        CHAN_BOND_SEQ_2_2_B: integer := 0;
        CHAN_BOND_SEQ_2_3_A: integer := 0;
        CHAN_BOND_SEQ_2_3_B: integer := 0;
        CHAN_BOND_SEQ_2_4_A: integer := 0;
        CHAN_BOND_SEQ_2_4_B: integer := 0;
        CHAN_BOND_SEQ_2_MASK_A: integer := 14;
        CHAN_BOND_SEQ_2_MASK_B: integer := 14;
        CHAN_BOND_SEQ_2_USE_A: string  := "FALSE";
        CHAN_BOND_SEQ_2_USE_B: string  := "FALSE";
        CLK_CORRECT_USE_A: string  := "FALSE";
        CLK_CORRECT_USE_B: string  := "FALSE";
        CLK_COR_8B10B_DE_A: string  := "FALSE";
        CLK_COR_8B10B_DE_B: string  := "FALSE";
        CLK_COR_SEQ_1_1_A: integer := 0;
        CLK_COR_SEQ_1_1_B: integer := 0;
        CLK_COR_SEQ_1_2_A: integer := 0;
        CLK_COR_SEQ_1_2_B: integer := 0;
        CLK_COR_SEQ_1_3_A: integer := 0;
        CLK_COR_SEQ_1_3_B: integer := 0;
        CLK_COR_SEQ_1_4_A: integer := 0;
        CLK_COR_SEQ_1_4_B: integer := 0;
        CLK_COR_SEQ_1_MASK_A: integer := 14;
        CLK_COR_SEQ_1_MASK_B: integer := 14;
        CLK_COR_SEQ_2_1_A: integer := 0;
        CLK_COR_SEQ_2_1_B: integer := 0;
        CLK_COR_SEQ_2_2_A: integer := 0;
        CLK_COR_SEQ_2_2_B: integer := 0;
        CLK_COR_SEQ_2_3_A: integer := 0;
        CLK_COR_SEQ_2_3_B: integer := 0;
        CLK_COR_SEQ_2_4_A: integer := 0;
        CLK_COR_SEQ_2_4_B: integer := 0;
        CLK_COR_SEQ_2_MASK_A: integer := 14;
        CLK_COR_SEQ_2_MASK_B: integer := 14;
        CLK_COR_SEQ_2_USE_A: string  := "FALSE";
        CLK_COR_SEQ_2_USE_B: string  := "FALSE";
        CLK_COR_SEQ_DROP_A: string  := "FALSE";
        CLK_COR_SEQ_DROP_B: string  := "FALSE";
        COMMA32_A       : string  := "FALSE";
        COMMA32_B       : string  := "FALSE";
        COMMA_10B_MASK_A: integer := 1023;
        COMMA_10B_MASK_B: integer := 1023;
        CYCLE_LIMIT_SEL_A: integer := 0;
        CYCLE_LIMIT_SEL_B: integer := 0;
        DCDR_FILTER_A   : integer := 2;
        DCDR_FILTER_B   : integer := 2;
        DEC_MCOMMA_DETECT_A: string  := "TRUE";
        DEC_MCOMMA_DETECT_B: string  := "TRUE";
        DEC_PCOMMA_DETECT_A: string  := "TRUE";
        DEC_PCOMMA_DETECT_B: string  := "TRUE";
        DEC_VALID_COMMA_ONLY_A: string  := "TRUE";
        DEC_VALID_COMMA_ONLY_B: string  := "TRUE";
        DIGRX_FWDCLK_A  : integer := 0;
        DIGRX_FWDCLK_B  : integer := 0;
        DIGRX_SYNC_MODE_A: string  := "FALSE";
        DIGRX_SYNC_MODE_B: string  := "FALSE";
        ENABLE_DCDR_A   : string  := "FALSE";
        ENABLE_DCDR_B   : string  := "FALSE";
        FDET_HYS_CAL_A  : integer := 2;
        FDET_HYS_CAL_B  : integer := 2;
        FDET_HYS_SEL_A  : integer := 4;
        FDET_HYS_SEL_B  : integer := 4;
        FDET_LCK_CAL_A  : integer := 4;
        FDET_LCK_CAL_B  : integer := 4;
        FDET_LCK_SEL_A  : integer := 1;
        FDET_LCK_SEL_B  : integer := 1;
        IREFBIASMODE_A  : integer := 3;
        IREFBIASMODE_B  : integer := 3;
        LOOPCAL_WAIT_A  : integer := 0;
        LOOPCAL_WAIT_B  : integer := 0;
        MCOMMA_32B_VALUE_A: integer := 0;
        MCOMMA_32B_VALUE_B: integer := 0;
        MCOMMA_DETECT_A : string  := "TRUE";
        MCOMMA_DETECT_B : string  := "TRUE";
        OPPOSITE_SELECT_A: string  := "FALSE";
        OPPOSITE_SELECT_B: string  := "FALSE";
        PCOMMA_32B_VALUE_A: integer := 0;
        PCOMMA_32B_VALUE_B: integer := 0;
        PCOMMA_DETECT_A : string  := "TRUE";
        PCOMMA_DETECT_B : string  := "TRUE";
        PCS_BIT_SLIP_A  : string  := "FALSE";
        PCS_BIT_SLIP_B  : string  := "FALSE";
        PMACLKENABLE_A  : string  := "TRUE";
        PMACLKENABLE_B  : string  := "TRUE";
        PMACOREPWRENABLE_A: string  := "TRUE";
        PMACOREPWRENABLE_B: string  := "TRUE";
        PMAIREFTRIM_A   : integer := 7;
        PMAIREFTRIM_B   : integer := 7;
        PMAVBGCTRL_A    : integer := 0;
        PMAVBGCTRL_B    : integer := 0;
        PMAVREFTRIM_A   : integer := 7;
        PMAVREFTRIM_B   : integer := 7;
        PMA_BIT_SLIP_A  : string  := "FALSE";
        PMA_BIT_SLIP_B  : string  := "FALSE";
        POWER_ENABLE_A  : string  := "TRUE";
        POWER_ENABLE_B  : string  := "TRUE";
        REPEATER_A      : string  := "FALSE";
        REPEATER_B      : string  := "FALSE";
        RXACTST_A       : string  := "FALSE";
        RXACTST_B       : string  := "FALSE";
        RXAFEEQ_A       : integer := 0;
        RXAFEEQ_B       : integer := 0;
        RXAFEPD_A       : string  := "FALSE";
        RXAFEPD_B       : string  := "FALSE";
        RXAFETST_A      : string  := "FALSE";
        RXAFETST_B      : string  := "FALSE";
        RXAPD_A         : string  := "FALSE";
        RXAPD_B         : string  := "FALSE";
        RXAREGCTRL_A    : integer := 0;
        RXAREGCTRL_B    : integer := 0;
        RXASYNCDIVIDE_A : integer := 3;
        RXASYNCDIVIDE_B : integer := 3;
        RXBY_32_A       : string  := "FALSE";
        RXBY_32_B       : string  := "FALSE";
        RXCDRLOS_A      : integer := 0;
        RXCDRLOS_B      : integer := 0;
        RXCLK0_FORCE_PMACLK_A: string  := "FALSE";
        RXCLK0_FORCE_PMACLK_B: string  := "FALSE";
        RXCLKMODE_A     : integer := 49;
        RXCLKMODE_B     : integer := 49;
        RXCLMODE_A      : integer := 0;
        RXCLMODE_B      : integer := 0;
        RXCMADJ_A       : integer := 1;
        RXCMADJ_B       : integer := 1;
        RXCPSEL_A       : string  := "TRUE";
        RXCPSEL_B       : string  := "TRUE";
        RXCPTST_A       : string  := "FALSE";
        RXCPTST_B       : string  := "FALSE";
        RXCRCCLOCKDOUBLE_A: string  := "FALSE";
        RXCRCCLOCKDOUBLE_B: string  := "FALSE";
        RXCRCENABLE_A   : string  := "FALSE";
        RXCRCENABLE_B   : string  := "FALSE";
        RXCRCINITVAL_A  : integer := 0;
        RXCRCINITVAL_B  : integer := 0;
        RXCRCINVERTGEN_A: string  := "FALSE";
        RXCRCINVERTGEN_B: string  := "FALSE";
        RXCRCSAMECLOCK_A: string  := "FALSE";
        RXCRCSAMECLOCK_B: string  := "FALSE";
        RXCTRL1_A       : integer := 512;
        RXCTRL1_B       : integer := 512;
        RXCYCLE_LIMIT_SEL_A: integer := 0;
        RXCYCLE_LIMIT_SEL_B: integer := 0;
        RXDATA_SEL_A    : integer := 0;
        RXDATA_SEL_B    : integer := 0;
        RXDCCOUPLE_A    : string  := "FALSE";
        RXDCCOUPLE_B    : string  := "FALSE";
        RXDIGRESET_A    : string  := "FALSE";
        RXDIGRESET_B    : string  := "FALSE";
        RXDIGRX_A       : string  := "FALSE";
        RXDIGRX_B       : string  := "FALSE";
      --RXEQ_A          : integer type with unrepresentable value!
      --RXEQ_B          : integer type with unrepresentable value!
        RXFDCAL_CLOCK_DIVIDE_A: string  := "NONE";
        RXFDCAL_CLOCK_DIVIDE_B: string  := "NONE";
        RXFDET_HYS_CAL_A: integer := 2;
        RXFDET_HYS_CAL_B: integer := 2;
        RXFDET_HYS_SEL_A: integer := 4;
        RXFDET_HYS_SEL_B: integer := 4;
        RXFDET_LCK_CAL_A: integer := 4;
        RXFDET_LCK_CAL_B: integer := 4;
        RXFDET_LCK_SEL_A: integer := 1;
        RXFDET_LCK_SEL_B: integer := 1;
        RXFECONTROL1_A  : integer := 0;
        RXFECONTROL1_B  : integer := 0;
        RXFECONTROL2_A  : integer := 0;
        RXFECONTROL2_B  : integer := 0;
        RXFETUNE_A      : integer := 1;
        RXFETUNE_B      : integer := 1;
        RXLB_A          : string  := "FALSE";
        RXLB_B          : string  := "FALSE";
        RXLKADJ_A       : integer := 0;
        RXLKADJ_B       : integer := 0;
        RXLKAPD_A       : string  := "FALSE";
        RXLKAPD_B       : string  := "FALSE";
        RXLOOPCAL_WAIT_A: integer := 0;
        RXLOOPCAL_WAIT_B: integer := 0;
        RXLOOPFILT_A    : integer := 7;
        RXLOOPFILT_B    : integer := 7;
        RXMODE_A        : integer := 0;
        RXMODE_B        : integer := 0;
        RXPDDTST_A      : string  := "TRUE";
        RXPDDTST_B      : string  := "TRUE";
        RXPD_A          : string  := "FALSE";
        RXPD_B          : string  := "FALSE";
        RXPMACLKSEL_A   : string  := "REFCLK1";
        RXPMACLKSEL_B   : string  := "REFCLK1";
        RXRCPADJ_A      : integer := 3;
        RXRCPADJ_B      : integer := 3;
        RXRCPPD_A       : string  := "FALSE";
        RXRCPPD_B       : string  := "FALSE";
        RXRECCLK1_USE_SYNC_A: string  := "FALSE";
        RXRECCLK1_USE_SYNC_B: string  := "FALSE";
        RXRIBADJ_A      : integer := 3;
        RXRIBADJ_B      : integer := 3;
        RXRPDPD_A       : string  := "FALSE";
        RXRPDPD_B       : string  := "FALSE";
        RXRSDPD_A       : string  := "FALSE";
        RXRSDPD_B       : string  := "FALSE";
        RXSLOWDOWN_CAL_A: integer := 0;
        RXSLOWDOWN_CAL_B: integer := 0;
        RXTUNE_A        : integer := 0;
        RXTUNE_B        : integer := 0;
        RXVCODAC_INIT_A : integer := 640;
        RXVCODAC_INIT_B : integer := 640;
        RXVCO_CTRL_ENABLE_A: string  := "FALSE";
        RXVCO_CTRL_ENABLE_B: string  := "FALSE";
        RX_BUFFER_USE_A : string  := "TRUE";
        RX_BUFFER_USE_B : string  := "TRUE";
        RX_CLOCK_DIVIDER_A: integer := 0;
        RX_CLOCK_DIVIDER_B: integer := 0;
        SAMPLE_8X_A     : string  := "FALSE";
        SAMPLE_8X_B     : string  := "FALSE";
        SLOWDOWN_CAL_A  : integer := 0;
        SLOWDOWN_CAL_B  : integer := 0;
        TXABPMACLKSEL_A : string  := "REFCLK1";
        TXABPMACLKSEL_B : string  := "REFCLK1";
        TXAPD_A         : string  := "FALSE";
        TXAPD_B         : string  := "FALSE";
        TXAREFBIASSEL_A : string  := "TRUE";
        TXAREFBIASSEL_B : string  := "TRUE";
        TXASYNCDIVIDE_A : integer := 3;
        TXASYNCDIVIDE_B : integer := 3;
        TXCLK0_FORCE_PMACLK_A: string  := "FALSE";
        TXCLK0_FORCE_PMACLK_B: string  := "FALSE";
        TXCLKMODE_A     : integer := 9;
        TXCLKMODE_B     : integer := 9;
        TXCLMODE_A      : integer := 0;
        TXCLMODE_B      : integer := 0;
        TXCPSEL_A       : string  := "TRUE";
        TXCPSEL_B       : string  := "TRUE";
        TXCRCCLOCKDOUBLE_A: string  := "FALSE";
        TXCRCCLOCKDOUBLE_B: string  := "FALSE";
        TXCRCENABLE_A   : string  := "FALSE";
        TXCRCENABLE_B   : string  := "FALSE";
        TXCRCINITVAL_A  : integer := 0;
        TXCRCINITVAL_B  : integer := 0;
        TXCRCINVERTGEN_A: string  := "FALSE";
        TXCRCINVERTGEN_B: string  := "FALSE";
        TXCRCSAMECLOCK_A: string  := "FALSE";
        TXCRCSAMECLOCK_B: string  := "FALSE";
        TXCTRL1_A       : integer := 512;
        TXCTRL1_B       : integer := 512;
        TXDATA_SEL_A    : integer := 0;
        TXDATA_SEL_B    : integer := 0;
        TXDAT_PRDRV_DAC_A: integer := 7;
        TXDAT_PRDRV_DAC_B: integer := 7;
        TXDAT_TAP_DAC_A : integer := 22;
        TXDAT_TAP_DAC_B : integer := 22;
        TXDIGPD_A       : string  := "FALSE";
        TXDIGPD_B       : string  := "FALSE";
        TXFDCAL_CLOCK_DIVIDE_A: string  := "NONE";
        TXFDCAL_CLOCK_DIVIDE_B: string  := "NONE";
        TXHIGHSIGNALEN_A: string  := "TRUE";
        TXHIGHSIGNALEN_B: string  := "TRUE";
        TXLOOPFILT_A    : integer := 7;
        TXLOOPFILT_B    : integer := 7;
        TXLVLSHFTPD_A   : string  := "FALSE";
        TXLVLSHFTPD_B   : string  := "FALSE";
        TXOUTCLK1_USE_SYNC_A: string  := "FALSE";
        TXOUTCLK1_USE_SYNC_B: string  := "FALSE";
        TXPD_A          : string  := "FALSE";
        TXPD_B          : string  := "FALSE";
        TXPHASESEL_A    : string  := "FALSE";
        TXPHASESEL_B    : string  := "FALSE";
        TXPOST_PRDRV_DAC_A: integer := 7;
        TXPOST_PRDRV_DAC_B: integer := 7;
        TXPOST_TAP_DAC_A: integer := 14;
        TXPOST_TAP_DAC_B: integer := 14;
        TXPOST_TAP_PD_A : string  := "TRUE";
        TXPOST_TAP_PD_B : string  := "TRUE";
        TXPRE_PRDRV_DAC_A: integer := 7;
        TXPRE_PRDRV_DAC_B: integer := 7;
        TXPRE_TAP_DAC_A : integer := 0;
        TXPRE_TAP_DAC_B : integer := 0;
        TXPRE_TAP_PD_A  : string  := "TRUE";
        TXPRE_TAP_PD_B  : string  := "TRUE";
        TXSLEWRATE_A    : string  := "FALSE";
        TXSLEWRATE_B    : string  := "FALSE";
        TXTERMTRIM_A    : integer := 12;
        TXTERMTRIM_B    : integer := 12;
        TXTUNE_A        : integer := 0;
        TXTUNE_B        : integer := 0;
        TX_BUFFER_USE_A : string  := "TRUE";
        TX_BUFFER_USE_B : string  := "TRUE";
        TX_CLOCK_DIVIDER_A: integer := 0;
        TX_CLOCK_DIVIDER_B: integer := 0;
        VCODAC_INIT_A   : integer := 640;
        VCODAC_INIT_B   : integer := 640;
        VCO_CTRL_ENABLE_A: string  := "FALSE";
        VCO_CTRL_ENABLE_B: string  := "FALSE";
        VREFBIASMODE_A  : integer := 3;
        VREFBIASMODE_B  : integer := 3;
        ALIGN_COMMA_WORD_A: integer := 4;
        ALIGN_COMMA_WORD_B: integer := 4;
        CHAN_BOND_LIMIT_A: integer := 16;
        CHAN_BOND_LIMIT_B: integer := 16;
        CHAN_BOND_SEQ_LEN_A: integer := 1;
        CHAN_BOND_SEQ_LEN_B: integer := 1;
        CLK_COR_MAX_LAT_A: integer := 48;
        CLK_COR_MAX_LAT_B: integer := 48;
        CLK_COR_MIN_LAT_A: integer := 36;
        CLK_COR_MIN_LAT_B: integer := 36;
        CLK_COR_SEQ_LEN_A: integer := 1;
        CLK_COR_SEQ_LEN_B: integer := 1;
        RXOUTDIV2SEL_A  : integer := 1;
        RXOUTDIV2SEL_B  : integer := 1;
        RXPLLNDIVSEL_A  : integer := 8;
        RXPLLNDIVSEL_B  : integer := 8;
        RXUSRDIVISOR_A  : integer := 1;
        RXUSRDIVISOR_B  : integer := 1;
        SH_CNT_MAX_A    : integer := 64;
        SH_CNT_MAX_B    : integer := 64;
        SH_INVALID_CNT_MAX_A: integer := 16;
        SH_INVALID_CNT_MAX_B: integer := 16;
        TXOUTDIV2SEL_A  : integer := 1;
        TXOUTDIV2SEL_B  : integer := 1;
        TXPLLNDIVSEL_A  : integer := 8;
        TXPLLNDIVSEL_B  : integer := 8
    );
    port(
        CHBONDOA        : out    vl_logic_vector(4 downto 0);
        CHBONDOB        : out    vl_logic_vector(4 downto 0);
        DOA             : out    vl_logic_vector(15 downto 0);
        DOB             : out    vl_logic_vector(15 downto 0);
        DRDYA           : out    vl_logic;
        DRDYB           : out    vl_logic;
        RXBUFERRA       : out    vl_logic;
        RXBUFERRB       : out    vl_logic;
        RXCALFAILA      : out    vl_logic;
        RXCALFAILB      : out    vl_logic;
        RXCHARISCOMMAA  : out    vl_logic_vector(7 downto 0);
        RXCHARISCOMMAB  : out    vl_logic_vector(7 downto 0);
        RXCHARISKA      : out    vl_logic_vector(7 downto 0);
        RXCHARISKB      : out    vl_logic_vector(7 downto 0);
        RXCOMMADETA     : out    vl_logic;
        RXCOMMADETB     : out    vl_logic;
        RXCRCOUTA       : out    vl_logic_vector(31 downto 0);
        RXCRCOUTB       : out    vl_logic_vector(31 downto 0);
        RXCYCLELIMITA   : out    vl_logic;
        RXCYCLELIMITB   : out    vl_logic;
        RXDATAA         : out    vl_logic_vector(63 downto 0);
        RXDATAB         : out    vl_logic_vector(63 downto 0);
        RXDISPERRA      : out    vl_logic_vector(7 downto 0);
        RXDISPERRB      : out    vl_logic_vector(7 downto 0);
        RXLOCKA         : out    vl_logic;
        RXLOCKB         : out    vl_logic;
        RXLOSSOFSYNCA   : out    vl_logic_vector(1 downto 0);
        RXLOSSOFSYNCB   : out    vl_logic_vector(1 downto 0);
        RXMCLKA         : out    vl_logic;
        RXMCLKB         : out    vl_logic;
        RXNOTINTABLEA   : out    vl_logic_vector(7 downto 0);
        RXNOTINTABLEB   : out    vl_logic_vector(7 downto 0);
        RXPCSHCLKOUTA   : out    vl_logic;
        RXPCSHCLKOUTB   : out    vl_logic;
        RXREALIGNA      : out    vl_logic;
        RXREALIGNB      : out    vl_logic;
        RXRECCLK1A      : out    vl_logic;
        RXRECCLK1B      : out    vl_logic;
        RXRECCLK2A      : out    vl_logic;
        RXRECCLK2B      : out    vl_logic;
        RXRUNDISPA      : out    vl_logic_vector(7 downto 0);
        RXRUNDISPB      : out    vl_logic_vector(7 downto 0);
        RXSIGDETA       : out    vl_logic;
        RXSIGDETB       : out    vl_logic;
        RXSTATUSA       : out    vl_logic_vector(5 downto 0);
        RXSTATUSB       : out    vl_logic_vector(5 downto 0);
        TX1NA           : out    vl_logic;
        TX1NB           : out    vl_logic;
        TX1PA           : out    vl_logic;
        TX1PB           : out    vl_logic;
        TXBUFERRA       : out    vl_logic;
        TXBUFERRB       : out    vl_logic;
        TXCALFAILA      : out    vl_logic;
        TXCALFAILB      : out    vl_logic;
        TXCRCOUTA       : out    vl_logic_vector(31 downto 0);
        TXCRCOUTB       : out    vl_logic_vector(31 downto 0);
        TXCYCLELIMITA   : out    vl_logic;
        TXCYCLELIMITB   : out    vl_logic;
        TXKERRA         : out    vl_logic_vector(7 downto 0);
        TXKERRB         : out    vl_logic_vector(7 downto 0);
        TXLOCKA         : out    vl_logic;
        TXLOCKB         : out    vl_logic;
        TXOUTCLK1A      : out    vl_logic;
        TXOUTCLK1B      : out    vl_logic;
        TXOUTCLK2A      : out    vl_logic;
        TXOUTCLK2B      : out    vl_logic;
        TXPCSHCLKOUTA   : out    vl_logic;
        TXPCSHCLKOUTB   : out    vl_logic;
        TXRUNDISPA      : out    vl_logic_vector(7 downto 0);
        TXRUNDISPB      : out    vl_logic_vector(7 downto 0);
        CHBONDIA        : in     vl_logic_vector(4 downto 0);
        CHBONDIB        : in     vl_logic_vector(4 downto 0);
        DADDRA          : in     vl_logic_vector(7 downto 0);
        DADDRB          : in     vl_logic_vector(7 downto 0);
        DCLKA           : in     vl_logic;
        DCLKB           : in     vl_logic;
        DENA            : in     vl_logic;
        DENB            : in     vl_logic;
        DIA             : in     vl_logic_vector(15 downto 0);
        DIB             : in     vl_logic_vector(15 downto 0);
        DWEA            : in     vl_logic;
        DWEB            : in     vl_logic;
        ENCHANSYNCA     : in     vl_logic;
        ENCHANSYNCB     : in     vl_logic;
        ENMCOMMAALIGNA  : in     vl_logic;
        ENMCOMMAALIGNB  : in     vl_logic;
        ENPCOMMAALIGNA  : in     vl_logic;
        ENPCOMMAALIGNB  : in     vl_logic;
        GREFCLKA        : in     vl_logic;
        GREFCLKB        : in     vl_logic;
        LOOPBACKA       : in     vl_logic_vector(1 downto 0);
        LOOPBACKB       : in     vl_logic_vector(1 downto 0);
        POWERDOWNA      : in     vl_logic;
        POWERDOWNB      : in     vl_logic;
        REFCLK1A        : in     vl_logic;
        REFCLK1B        : in     vl_logic;
        REFCLK2A        : in     vl_logic;
        REFCLK2B        : in     vl_logic;
        RX1NA           : in     vl_logic;
        RX1NB           : in     vl_logic;
        RX1PA           : in     vl_logic;
        RX1PB           : in     vl_logic;
        RXBLOCKSYNC64B66BUSEA: in     vl_logic;
        RXBLOCKSYNC64B66BUSEB: in     vl_logic;
        RXCLKSTABLEA    : in     vl_logic;
        RXCLKSTABLEB    : in     vl_logic;
        RXCOMMADETUSEA  : in     vl_logic;
        RXCOMMADETUSEB  : in     vl_logic;
        RXCRCCLKA       : in     vl_logic;
        RXCRCCLKB       : in     vl_logic;
        RXCRCDATAVALIDA : in     vl_logic;
        RXCRCDATAVALIDB : in     vl_logic;
        RXCRCDATAWIDTHA : in     vl_logic_vector(2 downto 0);
        RXCRCDATAWIDTHB : in     vl_logic_vector(2 downto 0);
        RXCRCINA        : in     vl_logic_vector(63 downto 0);
        RXCRCINB        : in     vl_logic_vector(63 downto 0);
        RXCRCINITA      : in     vl_logic;
        RXCRCINITB      : in     vl_logic;
        RXCRCINTCLKA    : in     vl_logic;
        RXCRCINTCLKB    : in     vl_logic;
        RXCRCPDA        : in     vl_logic;
        RXCRCPDB        : in     vl_logic;
        RXCRCRESETA     : in     vl_logic;
        RXCRCRESETB     : in     vl_logic;
        RXDATAWIDTHA    : in     vl_logic_vector(1 downto 0);
        RXDATAWIDTHB    : in     vl_logic_vector(1 downto 0);
        RXDEC64B66BUSEA : in     vl_logic;
        RXDEC64B66BUSEB : in     vl_logic;
        RXDEC8B10BUSEA  : in     vl_logic;
        RXDEC8B10BUSEB  : in     vl_logic;
        RXDESCRAM64B66BUSEA: in     vl_logic;
        RXDESCRAM64B66BUSEB: in     vl_logic;
        RXIGNOREBTFA    : in     vl_logic;
        RXIGNOREBTFB    : in     vl_logic;
        RXINTDATAWIDTHA : in     vl_logic_vector(1 downto 0);
        RXINTDATAWIDTHB : in     vl_logic_vector(1 downto 0);
        RXPMARESETA     : in     vl_logic;
        RXPMARESETB     : in     vl_logic;
        RXPOLARITYA     : in     vl_logic;
        RXPOLARITYB     : in     vl_logic;
        RXRESETA        : in     vl_logic;
        RXRESETB        : in     vl_logic;
        RXSLIDEA        : in     vl_logic;
        RXSLIDEB        : in     vl_logic;
        RXSYNCA         : in     vl_logic;
        RXSYNCB         : in     vl_logic;
        RXUSRCLK2A      : in     vl_logic;
        RXUSRCLK2B      : in     vl_logic;
        RXUSRCLKA       : in     vl_logic;
        RXUSRCLKB       : in     vl_logic;
        TXBYPASS8B10BA  : in     vl_logic_vector(7 downto 0);
        TXBYPASS8B10BB  : in     vl_logic_vector(7 downto 0);
        TXCHARDISPMODEA : in     vl_logic_vector(7 downto 0);
        TXCHARDISPMODEB : in     vl_logic_vector(7 downto 0);
        TXCHARDISPVALA  : in     vl_logic_vector(7 downto 0);
        TXCHARDISPVALB  : in     vl_logic_vector(7 downto 0);
        TXCHARISKA      : in     vl_logic_vector(7 downto 0);
        TXCHARISKB      : in     vl_logic_vector(7 downto 0);
        TXCLKSTABLEA    : in     vl_logic;
        TXCLKSTABLEB    : in     vl_logic;
        TXCRCCLKA       : in     vl_logic;
        TXCRCCLKB       : in     vl_logic;
        TXCRCDATAVALIDA : in     vl_logic;
        TXCRCDATAVALIDB : in     vl_logic;
        TXCRCDATAWIDTHA : in     vl_logic_vector(2 downto 0);
        TXCRCDATAWIDTHB : in     vl_logic_vector(2 downto 0);
        TXCRCINA        : in     vl_logic_vector(63 downto 0);
        TXCRCINB        : in     vl_logic_vector(63 downto 0);
        TXCRCINITA      : in     vl_logic;
        TXCRCINITB      : in     vl_logic;
        TXCRCINTCLKA    : in     vl_logic;
        TXCRCINTCLKB    : in     vl_logic;
        TXCRCPDA        : in     vl_logic;
        TXCRCPDB        : in     vl_logic;
        TXCRCRESETA     : in     vl_logic;
        TXCRCRESETB     : in     vl_logic;
        TXDATAA         : in     vl_logic_vector(63 downto 0);
        TXDATAB         : in     vl_logic_vector(63 downto 0);
        TXDATAWIDTHA    : in     vl_logic_vector(1 downto 0);
        TXDATAWIDTHB    : in     vl_logic_vector(1 downto 0);
        TXENC64B66BUSEA : in     vl_logic;
        TXENC64B66BUSEB : in     vl_logic;
        TXENC8B10BUSEA  : in     vl_logic;
        TXENC8B10BUSEB  : in     vl_logic;
        TXENOOBA        : in     vl_logic;
        TXENOOBB        : in     vl_logic;
        TXGEARBOX64B66BUSEA: in     vl_logic;
        TXGEARBOX64B66BUSEB: in     vl_logic;
        TXINHIBITA      : in     vl_logic;
        TXINHIBITB      : in     vl_logic;
        TXINTDATAWIDTHA : in     vl_logic_vector(1 downto 0);
        TXINTDATAWIDTHB : in     vl_logic_vector(1 downto 0);
        TXPMARESETA     : in     vl_logic;
        TXPMARESETB     : in     vl_logic;
        TXPOLARITYA     : in     vl_logic;
        TXPOLARITYB     : in     vl_logic;
        TXRESETA        : in     vl_logic;
        TXRESETB        : in     vl_logic;
        TXSCRAM64B66BUSEA: in     vl_logic;
        TXSCRAM64B66BUSEB: in     vl_logic;
        TXSYNCA         : in     vl_logic;
        TXSYNCB         : in     vl_logic;
        TXUSRCLK2A      : in     vl_logic;
        TXUSRCLK2B      : in     vl_logic;
        TXUSRCLKA       : in     vl_logic;
        TXUSRCLKB       : in     vl_logic
    );
end GT11_DUAL;
