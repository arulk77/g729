`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
f3hefSN9w0k+MPMr8O/pk/o7ajsiSxuhOs4t0XNfGLdazHFU1tbURMxRo8g2lwtJ
LZV7E29kWPhp4XNm7VWIk4bHV5ZKSqPzoEew+rUDy4uo6+FEJhEFHCq+R87+hYQ+
peGMBdxS06Zr3ur9LX4D9koWodoQk2gY3zkZ7N2qkZs=
`protect END_PROTECTED
