`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ab3t38y2wf5+qsH/48ktMCaSzgc+9Qc+kK7mooJKsXyvvngwQEMO8GZsYfK4yHDI
qaZB7CpMinfElzw220PPiHiFxp+AVlxABqCmp5tjOaCDxBa3oMw6BNF2C2lKczyn
hX0weh+WavWoUnZeL7fJDBifk8UHYSq3Gsvwjz8ACNdrKgqwU747N6uv4nu9QvJW
2DP9nw/8zpgsmSlrR6+r4P4JTPdSPcub6ZUy6tbi/1aOwKGXVj+71lr1OrFveZiv
J8M2ccrs1M0Wq0AVCTJPitI+p50kr806/MWx+wYXs2h5NEQjrOcG7xTf6o68H144
L4x9hI2e6fIYZdnaVt4TPtCfF1tdRMDJ1zkZ7CPkqygXi4syOHmW6XI6dkhB/mV0
+ZTrAunIiJzJ63HCg8rKW6yJPDxnvBYi1lv3bRK8Bttcit9x2hA7Jm7Z1hL5ofFP
+evk4JHV+VwZaPkOKLRY7dyGIKDni9nFIhVH2L8QUUo=
`protect END_PROTECTED
