`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wlweytJmmHNZ6FEcNcgJOhDGqKihZOZjh38bdIM9VGR
HB52og6+/sTsSwiD0M5U1NTlDEtkz0L/Tmmcnf1peal9+npu2av75oQYFs3W6CkV
hx3f8J8nexTkiY+3HHFJlMVLgT4BSdWowW4onhs/OwiwJKn6C3+iMXMeYGvzFYFU
rujxCmAZy+A39KIYzrNH0b5iw/hCF4EdPU3HkifluZE=
`protect END_PROTECTED
