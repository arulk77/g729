`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF45iFdLmctvdojJtjEIdBRzALE7IBrsll2lBYHK4doS
SIyHCLueyfuDbIoS9B+03mHVB0PQ0pAL3o5Zb5tBIMS9HaVtPl9zT5Wz6KJpZNr6
S0N1If43r4iInLv22WinK0WL9MrHY9WHw56VBXrry2boFia2speOP7qJlbcKVVMu
xE5hLXl0/VVeCrSybEYTZIWcaNyiqsLELvDt8epCF7XcXBJ/kVdhERYMoFf3asrh
`protect END_PROTECTED
