`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40aAHAearaFNVKpOyBA5NNsGHwXdcLl1vLYj9HtDFFX7
XOCfqPgk8rTpyH03TgRkn9U/Th8eopx/u3glafSAAq8URq9PFiOvbKWOPnLt6hhr
2jCO2KLvY5LKZ48aIAIylmKbS/MMhebMme8Xl7/ePwsGkV6lNZnDrh4IiuOZwENL
i7Jrk3a+cbcc3V5lJhU9WC5D6TBIFB8/ei32O00JmD9PmhrdhVZCfI/I5S4g9/Ul
I24nkfOoFU4lbMvAfPexFdoaIhQ6bxDV000fN+vo9lRnAaWdW+2uUcWQXh3MHnSh
UGEh7yL+pjNk7rn7WhSZXAhRnoOIi6Z+12bClFYQhPJhl7s1YPXK268ivwB0QbH4
WUb0OKv3329U9v+w2bqujw==
`protect END_PROTECTED
