`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47XE+mvuLSnmHpmc09JfW2ed7mASyOdobjo/qo5VhG2z
D//49xRTHPC94sBavPA4Ya5wfk9AEFfqmaBMApBdFqVe7Wz0vtotA91d06VP+tjs
dyL/piJS26ey3fqHYE+i5c+CM1ReBcPakWf08lyxYFoxpSUOLR9fS6bIHqJig8kW
jQe1t0bsjhck1O4XhYy8zYIKLrP7t6JBoXHzYDPt5N4kVINGwmxH7yfkNic9xzs9
2JqdDdQj2kro4JMr/k/gWrVnonRqkgKOkOu4je6rvX15DP58vTuK5xyUnmJCyHHr
WCE+omXjVMAjC2S9u39jOQ==
`protect END_PROTECTED
