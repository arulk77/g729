`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JS6Ee/OUguv3S0KjECptSLyltoFOXIovhBqInEb4HNdF/pdEDHL3aXvSL15RrKTX
qji4lO6gXh0kSIUkFi/15Tv6JEfFOQANzOwSX/LUK9scKNeRF6MicaAR1gxOX8C3
fPEWBz56H8QIVJGx+TYLafTPZC9WHNR/xLDHvAnKPEHoKcGwDlbyUaI7NYKR0o4d
c8HgL2+ZydkmPkqfpLb5aLhqB0HBuCxzxEHS9g7KgwwvCpV0BPDIUDmI/dhMJ4tb
C+IoODcdFCME/AxsSexVByA8bOpKcE8cCHrt2ZCrz7wHj2EfBjirWVrLFHM6x2nl
9el34ERifgYVKINS73BdkfuXyEwR4E/J2PxkThZ/qNr5q1ItRQ1VPzv5iG7NYkHK
N7LwblxWVQxcMmMtO1eD7vs3eO92FlR9wsTTCtATseo=
`protect END_PROTECTED
