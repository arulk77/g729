`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47T5prQYpNnmxibkhQ5tazAFhXK8q9Exp5uBBpxsVq29
LQ5hCF4LgOH6Qr3CExubtNukfZYRBe6sWQEdBe4pfgT9LvAxiBqtzzoq5KlYmP9W
MnSmdupTLNUc8qzQ1st+FnCwtr5NrF4nqdAew8VuqVRhwUG2osObFcYmbFUVd3rJ
dCxiZckDuDdJWLRwDWff7L9/3R0cQf1sZd4tv+VWZnmzuLsQSlSP6jWQHBxVgEyM
yTxMv4t7mbO9Ouu2gStfGxNf5D5J4SIPiynw4IeJPuDIooTdXUNReiThBS7buhei
BSYGX5Hd914jeiDL1GVENESjcKCY9u5A/fgtAVZawGkrTDiSp+G4EJ5IPBuIjuQF
HVPiyWcZzGm/1FZChLhg0w==
`protect END_PROTECTED
