`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDATG1GT2rdsscpwuKHp9FbmgGoJRcwf5c9d4g0hKnJN6Z
sDINlDWDR8/oM4Uc4LUWjfapK3bZguxJrerHLplaDtBFE+iDel4glL3IyWVPbi1m
LxSFYEgT3gEItvLGnRkVuQRpGRNX7KtSMuFQm3GYUDmJjh0shaShSSJXp/t/F5El
BlLG0XsYWiZHhqZkp6j5saYpwmCf/rfsZFmYD/csxQg+Cf6e+7FEaYP9xE5a4Qna
EFOMDpUJi8Z1O28s9LywzftnoBl/exoNM6RW16+UolnQgfIhFhdAna1lpreInp7T
QMpG1oW8NNvQtnCfXwfyWlrQ0Jg8C/ZzABnQ6r1+Shvc8040ASY5aK58kryFygBn
6lIggEd3Mk/ywHb54SRN+c6cFkVeeL9GXf7x7twKT5RU2Jpjc7CjczQSPbPc3IbY
FkYPZCtwG3ZSCdetXJrtEeY1biroP2fW69i3yBrDzDcOT+eZYA+v78TpW77BaFpF
XSOQ9CJ6AumZdjFY8rl5nT1emeGMU7XrGidMMVDWy0lgZdAGTwZx4C7MmHFEN5fg
yr65uxc8plz9xbKrN0gXr6hTRWtgHqPMnCLS8o4ecrP1um1PeNku/5mgvw1S0jao
ySQrTS1hAScMA/WuP0yHWY97DxuMzHsB9GZfv8/lJlfAdGanDMqmLAqNGa3FO0ji
4wpTuOoiUicaGamcHw5osonpCnrOiGIfgk91XcXJS4eM0qB3a6YVW63lDScXSi1A
TJEsWYGtnr38EMJL1r+KAjKtmFiMPDGoNbwmI5mM37XdPI4TjFJ2BUhxJmOS7xP+
VYFNYXeuRXX3RFCYjlxQ/45TUALpk2QIxLTmy+79SjwxjdfssC1gqNHhoSWmHLXd
XSSFqSiQ2HM0Z3IdHwjIcP9ZorSQ29TklEFdBeqFbF/2D6iJqSv1f/IgreP1VIzZ
nRgUycOud+QFQglXn6oHGSKFuWQi32FzxoNoILal8qt3iCb1wo+9aPeaVM6pHqjv
6cDpPoqcVOzMT5WMwapn0FV8c7HbF/KtoyLyO+BE593xGf9baWrisGmBPudHu8ZO
PniP8wY5fHyuZRfNRrJ1UYM9Diy27UEO0dTqT6urBFH0h5UZ6cumLwA9lkNtGJhW
X4VX34H//5ckZWe4TQVuzb+zTsnYrPsuuy146rmKK2rzIQRlB5BS9bk8yQvXaJda
RVnLlZ4io8Lj7HByS8btq8vOmNlWWxY6W0xQEqxTPeIB4jpGgBjKJEbrkskUrl6O
L8vY4sRcdsuDdGuVankAVSw7VZj3+8fcTP+7P13/UH0srv6pnfKvkCOHl1HZeLLN
`protect END_PROTECTED
