`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJpZWIos+mWF/9AeCWPSFM0zyjiOVEoknMMftF8T1fY0
QCoR0rWAvGp69gySKjwRCk250O3WHEOTbxmNs8DfyZternhRCzU0tzgwAzS8OTts
+NR5/Pt56WbqffhWajngwW4cfdXgjcbIfLsu96uxNz9+5lqXdjEsCmg/xgqnDpLY
9oCW+Z2t4Ngz34bZ3IzNK4KJdZt2VIE9PPiRe99tjuWk0GH4GXhECXUbgfhGvtno
wX0TdmRGLOQ+RuJK+o68cm54SZNcxMXEKmxyk+MflcQnZBYxgLIwBVwCcEY2szTv
Ye7RbA1DB/N4zfDuBhzntKS6wnOWSSTbBkdUnTmB5mRm/OkLjjSrFkZZ6cgWkMC4
/pCsObmYZbeacMiyLNCPdExuYxib5buW1FuBJAFVegxwBfKsSGaQVNuT25WVp95t
708LfTi5BQXVPEZyIcj0Qz2c2XqycvusgXtN39RrfBBwamlnsa4SFFwbe1+pNbqs
NhwuU82+vMxejUU+qiOFrUwxr8k3PgLl+2hk7tNsMkVq26XV13cFhUpJdM4Gp9oO
`protect END_PROTECTED
