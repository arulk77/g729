`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
nRscQNm4NBHBPDCfqVjd/g0ujTBE2k3wzr8/bQ7ch1D3bf5tNU++JLIVmFDz4br+
KlN7ggkV1OfsGvOsq22KgK1FKlpGRKY6Zmjs9UgKa5QbGCMBQTMVPClQBhA6S1UN
nZnwHx3lIrVKQYeE4ZYK4ZedypqAQEKW+/fkndzlWPIwEZXfpYRoABR/52bGycqa
SNpC/a1TJW47H9UYA1RiDcGV7mVqQZg1tn5pF6jc66+72gMFXGlAbJECVlWGSFkl
YnTUA5D+YbMX3N7mL/Zxg4jcsbvXaAb+IWgbBmnA+vw=
`protect END_PROTECTED
