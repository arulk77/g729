`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aWFxMIyRCReOJwSlK2VQqBQ+P6eb9RFTmS8/ku8B1mII
n7Hv3jrBxtgxToKD5QYHFD9YbGrW6VdG7DR4iZ5S1NAeCEDKQGv8wRm7i16gnPoD
Bs086k0BQvgyol5g8mJgMddDTA1FMxlvbNjxom1Wj4+IyjxW9Pa0J/G2ko+JQokf
5ElSt66stpMpQAXCYTPWwmUclH0P2+NYvvaou4AJ8Mrdc6IgW7co34xshTA1ars8
`protect END_PROTECTED
