`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveImpsW6Nol6cs77pn8Kr25B8G3TfNHy37rjL5ha8ROr0
dU3Cg5wuWqkCo8na1WzarnFTO5rHSDcm6Em+0UIrPRv52yF5I6nH53zGzU2tBHpx
0K/5GTjoebI6QNpv+1jWC8EReuDwYzTYB4tK5numg3PB19ggf4njJ5sJ5rrWCgY8
`protect END_PROTECTED
