`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
RGtwPMC7qTmGdgasTDMdDKSln42TfJ1D+noco9HVyo+LeDwdCNOdvcCU3Ae9WAbQ
dkyJulse9AKr+0Tb4p4DSa6USDKBA2uz250e7Q4Z9Qs7CakL6rbdcl6cjRCwWKxz
H2z2Y4kbKgoJg1xo01bjjZ6TQgbTp8mVHnLBexJJM1CurEGe8YvTHnnIC9jZfOTl
bWXb5fMUeXaQPKeYHcG5NeWMN0trz3X0fQFAoSuTKpvMFQ/eUU8S1FllorPie5fu
x1PO1OQYVnKgcDMCWStmtLjcAvk7aE3VkrDYS4cOMQ7LhwWT0VbT6YAMNoy7WcR6
3/jd2RUKJr+9q0ANv3djVUUr2K/9n1Z8Fsv/RLmb4jI=
`protect END_PROTECTED
