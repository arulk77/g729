`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIUZGOWE38umPiLjkPXejZBGPCOOO4XkuzxE0ofKeYN4
Q++EPuMir3NVsvkW9F0V3yA3AUTNlfZf3dCERmLoA9uxOmemgMMCJna2ovPLgY+Q
HomtuZb52F0rhc10HzEhqmSyy0aVQeu3qQsFbUcmfeg=
`protect END_PROTECTED
