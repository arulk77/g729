`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48tmBPP74+Ue7z6bOlNQLSCm7axUCpZo7hVhXBwFO20u
TGecnuucqg/MsVn/LcObF15yswZ4/5L2A9LxB7xL3Um12GNGaOoeXhNFa7wuiwc1
+X6UrSE7mMaaH0LOXJRm7yPviXMCqTJScxOQHSPnhbvHaYbO8qXur2Jn11PkTnPw
YCKINh5Lp8zgG31I/Lnfp9ZxOQBEPKy+I45hsBVTTJ3XPg9by+9YSxjkvEmDj9xf
3XiQdHHHUew7CcU49tmx7HoOk1evwnTgcSacgWAsWx2zHGUGpmQ9j98mdEwfyr2a
d01j+sVqmxRcDEsGS0OGSopznleBw3u72CwrTMe5Uu+WxQbnhE+saGp8lU0Ox7rI
hA+UBdP93WZrp5ohshfHTg==
`protect END_PROTECTED
