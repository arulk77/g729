`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveME/IBh2RtyOjsS7WyA8zxoFkbZ5n8+GldfsrEle6Nue
9vU/fzHZr7Wqj4QtYRDvLfZPkmHkgm4pyk5tN4IjqfcVC/GN0GBasBDwkBSOeT27
ViMGdNXcvKoNeliXlq2qz/jGu3tt3aS8oUNtAsXHerSiB9D8CQBjNL4aShSP6DIM
9nzlAnPXHCAvg6qVkLbVIdSaZOGl1NJfeeniTj7KHeSgupOGhmQcjGiC0iOd9VAF
+d69x8bYhngN4wJV2Sz1Sm6tKTvLR3++rdBxZOKa/gIT9ftRVvDH8J8i3HIhDYAv
2qVbkNS7NQogeXFJGGUGV0uIu8HHk+luvXAf1YC2T2X53VN3zhmURSywwv/zu1fZ
LEvtetgl1ZJcPtv0jpkDGcna95DkC/ZZV+mWDdaCpVzhqydKtxOfVf+R2lRUj1cR
yMogHPLUfvAQk99TbtlCb/ate8Ns18UdEAtCFu5u6dI1WqbDwVf5UXynphy+1ug/
6TWXHMQYWMBWP550a/CytsIdw4pNbX66aZp+M8rVGzV8NSO428CepVPu2rbv8gNx
`protect END_PROTECTED
