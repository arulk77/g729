`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ab3t38y2wf5+qsH/48ktMLarBahK+pSWDuz5QBkJQts6QJgMkOBqMLAs2JCGXjXv
pMhEElIfdkb1PQ92Ie3ipBRiZQyQSoRRjFlF7NOmUOIpvPQYnKYIqVFuLBdqwL0h
UbqJOzGOcDpuT9TgCOFpgOgyP3LFvaksphZIF9ygaEODuc/DLSFVGjarxoP/lWFc
H+GJeA6lAxrNuYa6z5Fl9gp2snrJC1Pic2qZrTAbprFOKnDjUP7iG6oHiE/HwHCI
EjJ0jJM0rPiKEcL+DIZFmRhcb+uVEf8o90y9WYuPvUIA6nY8nplsNowzMxIwa2IX
`protect END_PROTECTED
