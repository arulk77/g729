`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKtyN+OJucP4davfphms65AWBIUPQKwsAimfDTEqXN9M
VYLmmNUClqM9H4ZDjQhyuwOqo7NGW5ZcD/jbzpi/EIP8zK9dvDgCE7OE1LQTDvji
b5ZaLJTkTlfF7YpmJEC0Ae08txSAhaCroNopDblbTt3VuFQE24Ii7S6uPJXHIIZN
4/XwjiUtTHv8rMgpc/FK1K/j55EH8O6Ax10QCtAqzxuYidEEdyDwX6N0gpv7Kgbt
aPmMy9fQygU+O+aNY6Yzuw==
`protect END_PROTECTED
