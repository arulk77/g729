`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
VYOsOc83hnQRAyP4uwpF/RNqV29E7i3YvM5IFusWmc4TchoaTxoGdXqu5dWJsMRb
iwxNvEQWSU6fqbLXLXWVnpHkKSnEWxw8hldsX7XnQyC7KU/BRsDetmuZfZevbHha
tF6ne2hAR59dqRq4UNxikGayKCDzFIteoeeL2kuskcmvokW7c4wxXx111YH4Y1rO
NNk7JNqUvIpopqtrVaR8WRcmo10McMTce4yTpSjZtmPoA7E8TyIIDVfY9FQwoVuO
gCCv/M1iGQghxQlkGYUrCSAY/0FbqH7/wwEQWVumPSlvuQOUk4ltJ6vH4wmHZCvA
wNT55Uqu0ETP+8TYr/Vh13SZNkycN9C3vbzBXA1WEEs=
`protect END_PROTECTED
