`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKaZFvsgICVi9iEsuj73Faxw55Xxew93NPY5ZAoGTKw/
2B2GN2MPY3WCLe3FOshgx9t1KOmWoon1gnEcXmSsfY3DofaFLfNYVqlUztGjyNe7
ngHXlqemC63UgHel8574E14YMg5G/Pq2yNhyDrnOKflQ1ET3Z6BUlbz/kar+xFaN
0Bi81yF0ci6iN0NScNsAKuZA4GXOzj8aJ69D5bKegMAk+Jnrpz8QByyIoajPyDu1
3PAJPNCd+yQ6THeOScGK5UylqkK6TBDXu9hzkaZai4AVL/HGnlxl1td/Sn2U+Chd
`protect END_PROTECTED
