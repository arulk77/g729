`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wM0zfR5vW4k5dqWU9pT+lSNoBChLPPzPtK23YpenryG
BgiJsCKaqyOKR9L6ox6gVQ2CJ45d0SKwtwiKmyFiQqta3OlrhEkQTvL0JFZ076dT
+LWTakI7dj914oP+/qN57vwc/N160f29NXrDhYvihxknCrzGbPSM7UsVOhZT9G9p
DJsbunYKPwIccrt4sWec2tLkGsc2y9pcpS4tWxxiwWtAgY4ltuoqZFA/9CGpARdr
67HravTuiSQzA9P92lgJCwMLD0Ay2tRljDBzJ6JTx4CnrWSxCL+dFqyJbKpaLku7
XNF/f2NYKL9aI5QV39FjomAyMeIq26wBr4YtXpsTGw5AEb0TbZn3fu75rMaGUYNE
EoaJzlWi0T4rf0hZ05ozzw==
`protect END_PROTECTED
