`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zFTwxWtHalS1dXiSIV1DDOCHAnyMxAxO/ZckIWg/Kbg
I4rlk5WZAILzgICmT+40rS80qL55LzKoA873QLN0kgVauTtE2IeGYKJjyVivcVMx
svpQ+jxDHTaq8hFS85Vsw40+Q0NBRizRrjl2zgCvqV3oog/pQA//VK38X8Qx+VCR
AMtifDx0QfHvKmlsZof2HAncsuDkRZW5U0DdnQlcPV8K11rWb5InYg04NvTP4P5Y
ZLPCQiMO3gKCbrfa5n83qmH1E3hVb4tI322Bt5rYvsRypIQBdWnrjQZ7uNHzkayO
674tKMLVvYe/l7vVOKdZ9uuNsPmkBuc1v4+ngenauhqH8u9I1+v5mAUmCCwvKA/y
k7FP1HBZYzhnGUABgCpLgS1VXTnG6YkQCM27CFgtOYZNn67kDXT08k8S2RDh2VWs
A7AqWcM7anetcwk53DI5YIGYyOtL2POuwfYRoGTjxVK1fyguWkDHGPHsjgihGJEO
PDs6FCmzSpIms9/luWiBp4+g5tw42yTFuniTDbSrExJgIYv7X0CW3IOcvASbOL7/
1HM/65vxfLR7+Ah9pPGQf3FNy1DNAlnxvS8KQB12G/1d7ND+C0u/T/mnkeK7Wvz6
QZTezjH6x1Ao304lJkZWlnd7NaumFWD4mr6Vi6W9HqENjj0L0cIsopAV22APrtG+
JcwyzmEkrfFWay9l6mZem/mj2VHJRGBj0ZCEEWzRO09pelCxWK0Zrd50AxsJawJR
bT9X78qoZzkLQEKAjYganIhXXl1EeMz8vnthYFHkhAQNyOvaWIExXVwhB5GWS6Mi
9ejUuelXq/jx+pzK6zGaP7dDt78uMI2hTuQ03G5Rp108VLhpXQK8OksPMW9uXGBn
oASR5fkJOKJQZM6W9Vq7iHdgFeeuemm6W/ilGjR0ycFqiLDh2V9bUKFyE/kAfBJX
6z0KPQcvqptYKyk/OM886AjX7T6ddP/1OxrvH2GRxvM4Xqlv+7eexLKL4eGgxCEB
1gnP6u8aSzO1n6/h3Onodw2Rd+oFCLQWqk0x7cNlVbopUCENNYav1RwnzBGPfPg0
SW5HatyeaPzm2aLtjgI4hGfPfp7787pboFK9TfP/f9rMTeJHh/57TeGOTMC3zgGB
ot/Y5HZVP/FyjR5lovKXxQtBvJnT3QvKNITWcYB+owtufcrt6CUnB19fhzCyTaI5
l5sC/fprF8J8xn1Q8+sMWGgYXVdF8UvPeMcvW3ugqkpXqQ6Nppo6DdMBz8xtUu1u
MsDJilh5mjMdR3btVhYr82BvHp0YpRl8aWDduJQNxt7Na0SDQXy6GT4/sinFR8+x
b/JkN6vZ0dSFkaks1uKOWAoAclDk0fyNaEtWJvDwlWsu2Eyq4ecYR9PiwRid8io0
9Vqx6HglwIqFnbo8Twa2HWcmnUc+Zc4i3sIJJKo8A5jLyhGFcJf/9G+v0q2gW+6j
MOSFFMywwcjlUw+4qIGsLMOzEpCzYqde1S5iDvrMiKBhOiTqzttxIAv2p6HaGd2Z
Dx1e+mh3eukEbnUBVmTCGdgKnafgXY7Ia8Dm9KrP7s0c3aSx8bkXUUJSMrXPaTyn
d4tO2ZDGclGasNIr7FVj0/o2oMMtR3WKxL2OnyOrmI3B5B1kkFOnrPFX1YW9E5nI
v2xbAfjcXLyZ0sx+RSrGoDOQAtYivXQRlZD4zYuCgOCOhSq6rrWe7X+73uu3SS5x
TK4S1y6YDRPiJL9BzQy9Avig7AE8mPLzYArs5VuSwEbfb4563VuRlTh0Px5R9mHm
9j1b9hkttWZEErJhVp/qP9IeB53JAhkX8BrbxVY6VP7DDFJ2Nv0pz4ZusYz5ecke
Vy4RepqeZUJMGF418SAHdajA92ovkaYS26JlGuT3rzRn+utxBMKHRDeUQUmqi3Av
spPslgh9Y73OtjUgv924K8BkuK4HogKkNe2rntzi6wrjY454YCC5mMs/aezb4XQ3
FnQnUjVYZfYjgOkkEcMNLMts45dsXiGvNCZt/1afJENoeACxevJhEOMXMpVAMQ4Q
jOf3nSa1BcneKeRIhFx9MFkPGju0BPXids+cmivbBUft9wz9Oz+9kjMIqmQAwito
cAJ8imnoTbp78ZRWAy1YG46WjGxvwYzd9aWROQXUoNO3Xj6L5ZyDhsFiTF7GZAfv
Z8Al2MEC+5SOdYpUaSCDD51+sIa7Cgjr2cNTnWSCQ7EUBtfiy3t1k/P6XiGcWbAQ
eyHt/nzcrza03Oh658HUUpIRl8pTOWK6FDuiZSfLUyvbouN5TR85HbFgS4NNUHNa
6u5FosK0oCMX0IBZpWxc7xykceJUw62Ffp4Ome0iw1UAUXTv7Xh+nCCtWkplkqSa
cX6Ck0CfaYCb1em7cgJNzVGugSIDzHo1Tm2584J2AAuCMzLGPxN+ARUyCEcakcHH
xeT79TlHedezqzb5hVXOpDgkNtCnAFcstlgYfZ7duqRS51cK93lvF9gaf08a0E35
bD2O2b/DWYjPy7ezHByDkbQvJibiIjlD1RnF0PLpwBABSN/XLY80TEwHzdTTHTq5
al55Ms2TfsUa5bQo9D3emvv4iRZ1x6Bm3ync5TUQo3zHRWWqJTkc6kQ8e7av8cNk
I9uWlhzog0mzKEFzTaI3CjiyS2qFroI9MnDZ9ILcreXXChAn1+QQ0CaVhrWlyj25
h17UhqFJiwR1OA9AeZv2Ii03duQAQLJ/O9+JVi9phtBE9VHS1q3dFAM1Ua0YbZE3
lThnrhI6+mJCZKzK/31mF56uWF0K26amT66GKY6J/obYacDnVNjXx82Xi6zRbbTZ
h6HKLzH27HTuvfE/kX8/+zu3i5ZBzNuQJq7Ln76vvqyvvfc/FT4OXQHZICl/QVRS
/oqtNeB34DD3LZQ0xF27LGfcX+DK85kq+cCVooSq956mw4q3ioJCxaG7JOff4Z54
thmdeTKIVxJX6nyy50uUzlBKPYoRwatAD7BKV0IuX/CYG0U+kXJUrvbdsp/oa/4L
sJU8QTH2QjHpxW/aWZ8pFt0CVMg4dhScVnPWGJX1szXXJmsi6ejUPoALylfw3FFw
z6N6H5L26NPYl2W2MtbROdtA/4huM+ArphX/77R6xdo=
`protect END_PROTECTED
