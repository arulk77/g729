`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Prgb+lMGK4ankHVaNnLDqxDivhhwBb9BZNQe5ypThnENgTwfDeb4E5Z7TNY2QUJZ
VrZ09qeLT9Z9RgKfvQ+irHbs5t2HaBGaandCNOsOaEpq/ms+VffRj29zZckfswOQ
PyTpujdHyesDmcMKT0MaVQlOZBLzeyB+JYN5xQXJ5/vQxFPkt06A5roHQfXGaMTB
NTfrqM+uLAgcL+LkN49CC5/X4RzmyY5wtRKoJLAsoaSdJas4ygCLRcb93tVwRPxr
/i5SmcIwrU9hENFpq5Jslz5J8d5/4qus9kU6qvgqc1Vmb6KtU7L8KfhIT+o4pl4c
1QkeB78s0ZmZmTLFmn45NtZhoZ+vPBg/yLAFKBy5CzPZz4I7Zex7hQeA1W202zqx
`protect END_PROTECTED
