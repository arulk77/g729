`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAcOES2EaV4EJb290VIqrKlAILVgaB2byBKRWYSWJ3kdI
YDXdhgbgwSHnrtxdIahGeCWzAuUjWswYn8bMGTvGECe5lyCGHwD8OZkoJ4PEHmhk
jfrebAvv3bzy8RH9GtN9qOrFipTEuZhq3gDx6OptE8kbrUB0yYtxcnF3rVSCp2ZG
0e8VKW+xqVMOwO4kBtZIHmepaZxLY2KR7a+pKxmLv+ecbHRHY3z9zUQO0aTecVFT
MHPZACO02wDrPIDpWql/4ThZg/WwpAy/L7QIIqHQ0d+847CuXSu4ifR0YJxsfrXZ
TMDqp1rdijWjf0EOEaUMlZtTtAFyeMXWFErGblQzvAGdx2/iYokZ7QpgeHFD7RYj
k5wBnWdyxWirHR2vgbBqQOF/wPR7JRJEOSbON2qpHcNaPZ8aF+Xjj+ua92/8QWap
IJjqis5uUUOtgjvqn0AU0ViHu6HwvLQ8u+vxjOIv2Gw1OQtuU34nhCIrN3zicVvf
bTkuDU401h4Q+trEeycQZt4EKP0yzDWPXhCN1XdeMKv4Kzh1MmgNwQ2UEu9ultAH
`protect END_PROTECTED
