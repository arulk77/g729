`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4326CgMOZDYrjVHZDBxIkDGOWnGpk4zNO9RDEDsjH0Dg
9cps1v+iOa30Ask0+LcU9ImKD9tBZsAfzV814p6zqCL+mcxkDd+1LChoOOjjVwyp
Omym8eGGN7fpnMArdNWWH9hR8HEHVeWbCQsHR/QjSwKaXyRy7DYMZ16cD0a/4eLC
9LB6AltrGwEKkxCOcg6eBZv0N4gfGHAcqu8bu/lBP5awGKfLM6Ly9P3E6ItAAh4u
rdAZnfkoW4Hf6Z85NpVCkRdbuzvoJlNtk03ySsgUdvA=
`protect END_PROTECTED
