`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNye7rw4PepidgPXNq3zGk6oMSm1pQZnQoUzCQpzCdwP
SBmx0XYdDKDR2MylYfU1vBMKhlHzBSa7hXc0/ombPCKnQO49c9ism1nM45n7CnUM
BDi1rHjerwVTG7HwVm7reR56tSfNlAaHfv1JciePy7vPngyopYdQ9yPgp0dL/vGs
P9PMrEgwlCEyJKhY27nAUVnlHy5sd5ZTqMWyfnJ0hyrxC/P1x5Wtf3YIFFHmwjVN
eziKEHnNZlWpZaYPsYuB3BM91qPmItP1QxJucwoMHKLznRLFTbn/SmyMKVOXrJ9F
4VEhsStgnGgTCrMI3RVo0c1ib1yk/c/l/2MvGbhxL8vcLZNxprdlmtq5Fe3VFGuI
MxKoaOMOH3y49eRlGS86Sg==
`protect END_PROTECTED
