`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKt4dXWH8tWjpVmtXlJiEUwFPETvAEoRvuH9BJjAKEhC
XfAqBfBA7d/hTYwgIeCYsXucfV4p6QG6rn5NAesnwZ3WYsZff3/O/cMPVtlgcuZB
YWvzXn/qA1H6nVVsypBnNPb9jDCTPhR/RMHw6bswa08nFnVjm1k4DHTtYjC26lCc
COPeYh1HcaMK2SQcVaGwVTg19NNVdhhIvdTFhF825Sw56EVzBQOUwnxVcHvumo3D
`protect END_PROTECTED
