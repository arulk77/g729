`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOse84+uWOhn3tR/OBWQAxtqarakHT9IUFwLK1OX4TQC
PqQIFw/Fo6zGvmNDvPk0lE4iuKGzcVENSYeJOPpjednjaXpTrqdqscrcNiXVY+bv
nL2/6W7WL2uxF1pL68ZAT2MJ2Xs8OMScPVcBYI+AOQsXfUQ0nk41Wf3V3NwZIa/b
VgSJk5Iu58TTbsSF7ydE4Q==
`protect END_PROTECTED
