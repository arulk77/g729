`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
SzM7JWeDlmHa/ZyJpwkTw6P5ORiC1fpOuwr3lMUl5v5TaVQwuUhclYqH0V6BcpjP
B35ivEnnQ6dHGmCKopdBPtLFzsegYIQpnVC+SyUKK+O0vNjidaVtFkUgsada12vy
fNV+xXbEnhei9VdYYe8AFEQShqHgOtFu8u2kXm8vDCke/mzG5mL4teuQsLaJ1HiY
CSlODr60BtfzaZxhImgRGuKxRmJ2GMl3ZphuqLH7cRZOYz8XLNxD2fwFWyvZ/vYV
bo+YYKsQ0JWNJ7Os1Tch8GG2RWDNc3fCEKfBjSWwj/4tLZjFxIaqhVUmctWsIiWw
U4JhocFHRC3VeqvzETNuf14FnD1KvZASm1Bw6R0LmmBdVNWY4baYY/0E7VbTqEqa
BU5ouv5qS5CfwabL4iNvAr61gxHym0zz7qzEj0cefuzz8qwbSX95jv8I18RDj8hp
1bvTZP1k5s+md2yCtaxqh/8CMGpl2IPQ1er5PsUfQ5nhd2pJZ3U5FsK+ROZe4MUT
O784AwyJGdgXW8lnpZnl0p6s7VLXTO0t3cVnni7IvQKObtFpJg5X1MGFNXdUSdLH
MHA5DT/7jjLoQ/6I2bJa4gzijU34HsD77mWWwnmganQiIDE1Y7x4d7HV6VPiOtgh
RI8h7sEl5tZI8NeQ857y3Q4WM4B/6Q3nLlWETh1WfWm0c7JRge7zSv+0HkBu4D7m
/vpg3c4lH0ps51z1t9rdYkSIjS3CkstuRzqY+fm5neg+1Ky2Meg3XzDmZ9u/d/BH
n8TCbmOm4jsAUYczaVskpCskaihAIZR5vSL+8bUSJoa8bXOgFezv9e+EBN6iajbb
WeCLTjAfWh0T9BzSOQcHskvZPt+Mc1AGE77snhB5WBzYQ13S4jACqCGBaGpudJRN
bRM5PrPSIBCcBCZNhuNlVQtPhhHXn4r/7Rc+IPUhF3T6kVivOAnb3vWN/SxZxLhu
HkKWZwiZtrnE0D1nqxEvsm2dcvNBIYWIGdT+ttCXqopHV8r14wvSSIxkXchRlDgS
0JlSJoBwwfrMJRRkf3WzkVA9wG5tCZukR4n8Z3ury3cf1Iv3n/cYi8oqR+21NOlh
hVtqXt6KOXsjBBUZbGSpitrIaiZJL2sEM5BeMFkyCXuVOwHykVC/wnuvymQdPleU
wG/dVvagI+oUfeI4ANf3RlcNGGeF3/qjHBa170zUyiSdYB5rlYZE+TJN+HO1Fdgg
Go7nJUZumAq0k4JaVocjzZJLbKFK03zEGVhm7QWUGjeX18NPiGQ9t41ZDW1CXUNp
oNUpBGTBHkWY+0wKtLAOybN+9mt6zXChI3eI5GGKlDA8lgQUheNRlOK/lQYl7sZ+
+wEGvVqicsxefGIspcp7elC6E80oPN7JtzgIJrCS9vHPp+kK8hcABBdHC6yxSSHi
pfDUa2/OO9FZ0guHYiDHrC31GUQeeIpndgheNRVTTGeAht7bjHi+V01GrMck/FVk
tzrOxneYiXCUL3WPQipHvpqy89/NDO019Ce5jKeOCtX458+RGYHO+XZNSB9s+9EP
KvhKq5ga8W7nXajJ1cVoUz6HBrtLBqbQtqU9MtbUgCz8oH6a8Y3/uR02hAsZOhG9
ALJUUBCFcO59PzkhUwwXqfatdrmo+a0nyoWgqil0NXbJEb4KSL5Cdi4YmZBQ8fvu
EaZ920BkW/Xu/ITLGbpoF5sVyvGbmFeDkz40aPyRI3hCpkG34BCRMNvEq1q35Hle
IB0+Gk8maErmXobP+qdjJNyQdEhhMe/7Qm0orhRfdkN8mhDOTEXlN/DqZh32ZkfU
cbCgxw1AGP+jcwUb0ad4f0Ff6dpCyThS1ymxnEnwy+9KLlNXEVdFG3ETdxRv1ClR
sllUcgMd9WmDaGwToJn/rsLfqKMD/Yot3yAQxi8jMFTbONL4u+UoHsV9W5vSB/If
GR6RiR4scjxvnkBogHIrzyj8elgjs6WloSDl9SWLTak6Tul/03ADdZYAjY/asezi
PzvA8PMgAzCNCBz+VZJeHynk+pTNA+nRpCyjj33pi80TPnaMhA/7wzKTaon8sWCV
kfMSIiqFhKZA3BEUa0j8JukmcCsS5gPBPb7Ou+3P1u1SqLYfXpGGtOqdkXng7sU4
DzpsOyDSDUMLaCI0MPV1Gws6z9P7FldM/7lgKd7aug2asO6p3t+WMUjhzDC1y6h8
kk472FuD2k2RToWBUvDKduqYWUxSP2QM7YyI1+yNBc4zfR0xaoJdbUjJqdrJagYd
EHSYF3rDQ9JtfW4TUOmbaSs4KCA9HW8+g9Q2eB8vw6oNHCoOAM0wEr1P4edfwnVk
TlP54H3nv/KCrl5gTxZo2GAWznSvI/hH0ogrdQtfRC9xzC+N38dKQaUF/ZCbBU3v
dBeG554eKv2ktSTEIPOpPpVnaUKHfxgMhShspaefvw5Bvu5EmYkZK4ZthiN5W9g7
1DrsJqGBIIhrKCqt89hvcj4ikXbYnJEGpgE80ItM2pek+bxWWByWCOsfG3ceBnNB
ErJtpX//hfxMzShFAY9WeoXDki6PY62q2FPJoC21sW7gcWBLowOUnG7RrZ/5adHJ
O/xtthievgo+uTRou5JtGrFvvD/zMysuO/0iLEVJQkwGSo83dzee/iQk1xdEJCzB
3SmS6W5c+7G4TqYTl9zXBUT3xbyDYCZfO4J35ZkmVRz1K3GNjLqOMh7uOqZ4PMGZ
Uabq5Hgf8kFPVCCk3G+DK6NxPWFeCmWCPGXFVKsfrzgIk+GURBd35USYDU5qDcGE
AdAVXo0C6+QhbBXT3QMLw/uIlb/Psb2S43w9JbYbbWqpo/LnTCzwNmY+ZhDqw1mP
OESbJpC+BFgaI3xFYmsuuanGw2MGD1b8QogJdE3uI+ixun6+XzuOQB/5uVuRYg+w
rEU26ERy1MSYAr3F+qDTiQP+EOwh+LnofNBL3p7qn8N7M5d0nKCa36zPa3UHSGMw
oK+/KctBYUYppj2qW5n7Yavt+zLACaMMTkxLvlT05kNvkpen9DIs6k51AkCVDCsc
RS1ZICrDmMkhP6arPzzZSZ1mB5UnA1LrsFQ2f6V/IayMD22b2tL3MTKKpAdCcVNn
Oy1TCyoSUDsV8X292dRyWlNiwKh0yUZbgTEM/Sct7f2UHN/WDBFC7rutQMXe+EbG
JTRzNfw2Lg/yBwqdZBK1rshTyvwXc83H9L+gN5HXyzgmiYaUuBk7fI/rlRBLG/LF
7lT789qBJy5JA6NE96w1K50O1qL0KzCEYzdEzIkHL1EgxjGgdfY+VtTyB1zGlH6v
RDK9eR+CnsA2Cs6K3XrgEpr/3UTPlTMJR/fMs0zP6cdaUg1GT1ii2T5FtV8tidXr
kHfnjkWIbgriiLzHaKRwXT4yfA/ITqkQnTN82GYyvo8bOnGNVijaWfeOZXY7tI6M
HtjHSUEXsoM0a/oPGRYSxdRZPkDYbL17yMOTExM2KvJIQHjSenczbarHhZhOh+qw
QY/qP0UAoWk6QPq4BDFYpY2FNacMpCr/2NPxn5euL0AyHWUDl6QbPdUVjLs/WYGB
nlu4dqh/YchDR5y1ARJnJxO+w07ZP0kSJwPtFJ8vfuiasStE/beEFxpHFS881NWU
kZHHbZds+xwYEMZw0IOmLyAwdvC0N8gd+NP6B2iRicLmEeFTE5YQpU4y4kCt5BCv
r4eFSmx9tGSbCvXKqoGnLkQPdO5ZE6UqJeagbGU0GZlScFeH4zh7My5IjEf/lmDG
5pjYaOwKdHMzC417BE+l/9vxT9LZBav4eezBKUopZKNQmg4jyCKNc1UBcjxDN92B
+mrfpiqAgm6W9XmpYfi5Ok2LJtLDVvm6qJptn4qamzLt7W3kf5uF/++VT4EjR1/B
+mmsYHEp7F/KGOTTi3BeAXHcG9o0kkrXyqulDwkFrDAcPByv5aZSumkHig8xv1JB
AE4jiTPVUSNyV9z8Egu0W+hoZSkafW0vVL2Z+Sz05L+gl+PzdRp1Wepwt0ilRrs7
VMNiVCCNQfFBVedHOjHGJL9mvthIicbchVygLZgXaeDKKQ+UP8DPmMQ4GJBb0GXJ
vfiIHw7mRSbncNX0ScH2hKhsFW7c3QCeZxL4AKxzMapHuy8vRx3A4byCFVJPode6
7K7f+T4JuGZg/44/VAdRHI6uSsR1mqAm8BNccigh+UlTfSJn8QWWgzW/mHyiIgJZ
F5uQVXPLtri/o1pYPWXXR5QnFKkxOtS7PWF4zH+Zrwvya7fmDcfITbjQbGAxZamy
+IridADaVPVvrA7bxiUNa37R3dw5WoAv5CWUvzmQDCzfcKPYBX3kxcHgAfZneJfL
+YxR8QRZdjbGXc2mWD98udg73IVaR3TDIrnPjRGil3+hSCpLLGEjD+8iKIJzgAA/
J1Ab3QPMXJSyPqagcR9MWEJ1BDWAYfCuY60nwILwwsbJpFbx2eQMaNHurcXl1cqE
JDmtMtJOc65Zt9S9bbzdcx7sHqQTchW5SbGlvojmIxppkqktJDZ9Q0OHuKvv8Y32
DJz7qozXydo7y3EIB2x9BSDTBRVQkWhA1XFx7K486Dpyj2W40+B4lODbPGLMGYwp
Bi88K5K0BMZxeQwuHXEGjsww3aoL6pCYzyjNr6ezl85EWfcQVKAq8AqGq04tSTNh
fjlG6cXUT3mgg7yzdxan6pJCcRSLu0FGy76pL/iTDercerlNqeEpxgoTpVZHD8Vf
dirY9bqjF3VlywlrEPKw0pBXP9c6t+znTYW1VzAcpK00X+Vhu6xAWNBhFlktQuYw
jsGEUCG+xrNB5lFLU4krVZjHY0DLPMiIk74sln4ApG8Qf0hNBBsmtSA7BKqufNvT
26F1LpnsXES6DXYZqdIrQqNkDD6ztNcLPNK687t1OYJ02Ajy2Vg26JIal8cJ0uJh
wjOSgdKg0AhLy5hieLljv61DaPrk78yiPLX1bI0RznEh7QAKr8sm7MjN43A/wMbr
/XSKk6P2qvfy5IIqqlVGaE9086hJkhESM/vqB0y8ASqtdxk3tUwnItYbf7YgOzvl
CY5ODbLGYFgohZ3LU0x8/pDhwkLz9Fo0O5ihKRhWAsTfTHJNLs/VMAf1l8L5tNQD
YsF9TP85s+PEtKGxhuNu0mDPufGWboZ9Hlvs0+LNdP5T1Rv/Js9vKL6B1K+VMIl8
mQixA3E/HsY/TWJkvHtAD+pXgXAU0Wo5V5EcW7lnAZe3z1xob0vsBVGZkQNLICzT
ytJIIP7WuTDKMUrhztc6gnJN3VeYw9pUKdAYL8ExEDw169xJdNc1XwLOtIzx+q5X
8LMIisWSJQrcqIKmIxz3G5+gxaQpyl3IBRwVxerXjCr2Sb0ICVi+MEp9Cwzwds/e
wpBy5dpUAU+FvKqqPsieCiwVjgsyfhRJc7b+hg97QGWm5rUABfrEhpr883/33HG2
V9W8pphOixfp2Bm6urV39Usckh61MK2xQnJxNGUf6TwK3c5kVyWqHsB2tn9+iU0r
XjMBQBbr+sqFN9cS7O+3/WOjZ9zoOdzhuwTg7CcBqaR5ddAkGQoMONd5I1z3HDO1
J9vFcd9B9/jKVEgH2vKIpOV4ODsyYqjEuENGuoxfBN0xdSlr7vziChuY+G5V4p34
ZR2CaSTk0crvxcrO1gB6cBvhdj+IIJzY/Ayte7bClczN74s8SkUK8Wcp3Fbvftff
JHuC8h0qX8Fgf98nfVu4ZP3xjIjzejcai1+RfPqv8+Fl4FpaF8mBdbdjeSRrGezT
kluHFFYcJttlfojWPNqrcaKhzWuJnNHgBzHYPqhXAae9BG8CYHi6QUxUpMu2r0qw
f1UqutcGdBbsOKQvyrMygNnwCSQdDZKQuwNlJOKpWJekhL+IWMPvcAGRV/ZKQcBq
GUW+rLweGh9kUxrt43rh9TW4auP9vkSczA4hpNEih7XiscPLUgIFMLVsPxprXxSP
mujODvbgm4yAtflEOtoQwn/9+VH5p/Tkvj+vECL4mvrRPrEmQA3eVnnWbPohyn6X
50sGEVmfbRaXqW2Ta1GAWJMSqb4/bf+hZYq9oXJ4eDdruRiVBVsBShmYcmxr/Ga6
iSHg4df7O0R74gb5r8QUvHJRW9va9zN+bCGUnEX0Bu4tdAeqymBrwrBlSno00elP
/jkOvPLKmwkMkN0Ej8dEG0sdJeTtaYmS9QYspvbcvf+bH3ZlZnc5qJizk7xNbZwm
a9YDEpyov6+7vzbGZOcu1D5JK/4fw9mpOqj3V7mrGt3hhsPRvRpx4d7fzNuW50M9
Q2ra/7fZ2cXf3b2lfEA7iuk0IYb/reTzYNs2LxX9rXAnE8PU0y2QCdNEF3XGXY/G
FhIw5NyFZw9lzk2QK++UIYg2G9UC1iAprxBDNWUHkPCFadIVZEhVj4YndHFPT9ZM
OfSkVPUu8LFh1889b5SgGg7Z+Y5ulWZfBTYhZDTyGjVJTeLB87N4ee91l/Rrj/pX
LO/dolVL8hoi63H5VCVHx9W+PLPs48LyhHXtEULlUXTFSW5qjIBIOU3eEVmCnFNO
8NqmMWXWPxoO1Dy+hn32sSL4jalFPlQcDaMg0W4zOIF5JPSfTohixKJrTofN22FQ
yGP7IlYwbdnyv4lkYLLJBlh84ynKX2+et2A8z2DPawCdHuscJYhtgURnCIpxzxit
KBYqpDnd9LqF1tvfe4REXbT39r2GGHDkL8BoaL75ZMqkV/rTFJZhFbnXsxh8kYpF
JOLW4aFPqQGAnP8y0dS6UTclW2hkAWgfvtwZkuf40kVLLZHQeE14P63eODdZhxeX
hmUiO/1oSXp7TKaju9do4vU6VZM+PjJJl1HqHM1oLbgZH+b+HiOQNS+OF0yQTQhW
ne3JXLdawqPEAVcPIaZFY3+KQsBscfJ+wGHeY/nbQfgpGm0u3VKccgyEcxgvQx97
eJ04S83umKtJF275Zq6HchxAD5yh8G9CX6OdBsvRC1J37zlXGcamzU3nLgmSt2yN
aixTS8+v+4O5pswA8w85ElyL3K/xA5OJaY0tmFo65ZNcCLYDvxqHytFmAx0XAjvD
mZ7hm7LxlEgWDv5cAjZFCnYvipNaM3Sjaq9EkYoLtY5HuQXaIl8DKEC1Kdn9zrdJ
GpH5I6Su+rfLsNxq3806q40U4ILdO2aM1BNxuIyst32qqcnY67tP+oKGZCKT7ITA
jZtumft+k9mb3EsDG1dY6K4KMYuVrD/AavSKUJhEPDUxDrCyD2jd33uTwJPSfJ1r
TQg+d+FkkX8/ZZFmzXEQOjy+3pQxfeXGzMbS9VkDGzunN0QiZXEk3UUdlViN1M/0
SH137wJJqgL9cBQWQvaAnkUpqbNxETVYLZC04mQ3gnQFgGYVZDvnjO1xyGPwFeek
HFzeV8/pWwfoxfzo8MN+W1Nw+ub0PX9yh80Ss1CgfQzWSgstBvS+CKYiiZyPbMkl
9cVKGPWTIMctOkzeOVAtKH5m1SH8lN7b6zmdWTa9YzJgCifdgV8lKIYqWhtZFpum
LYMs6o+KbUyGhN7+CN0c23QvMprXLZCDSCI7xZ36QmxBlIw8EUp/SovfFPhfWAfe
De0riegKwu5fooSUliDF3Pb9lMak1mdaHrU/8woeudw4QVsh/dYQO0h9bFz13XdQ
1QCJr51PTJFykTTal4tobMgAI0oZOP4fMJaiAFkf3/jdsb2J1tmcvoAGUVzXj6EA
hHKUPanUNlRyDPJuR008e+Su0VYQxjQY2FqBI89fVp2rND7JwvFfArLeuHwCA0QL
rCuftCAPJjXlrOZ8JQgQbzFe4DOqlTFUHW3pn69Pzs0jZpzrRXWB76JuSye0HiYf
2WwQBnx64SrtWyo3J39NvYREysIYeM0mg6IAwUhD80RsEdlipYnOgA1/cxw5ujKW
0nFrELBYBxW+ryhAAdLpiGHWuWYlFgUhIdbkBX4aBtU4pgIBwi81dw1KmfNH2OKb
1XL98rhw/QWtsEPLW25MxlBvCnsK3N0rn4OzkTMsdd82G5f49mFS8m9G8Ziplo7M
ZCAaRUvEHoh8aI+y8HmFpAZ1hz/1K4pwTUlNyZwrix8YykiB28rRzTk1+bS7RRDN
olwgesOMn7ytcWmwJmv+MCJ9w4QHNb1sbl1GjDcRip9532wT2Qc+ioXNajim431u
VjdbAiINu21hwxD3iOdiWUaq+QlYsockWSnNeVp+b5Xu6/ipGV37+fPrLPZgtyuN
FE63vaKzTsInTdUTFFzKM5kMTBcWoGlEwRb25sKY4geYzWnLG8s0TMWDi/H7Vv9B
UBnX0y2HaiNM5aI8wR4xQwuwM4hRdcQWjAPJSk1YPNMqFaEBPpvrs2W0gQ3PXJZd
vg4PeRbLlWTgV/XZjovjnHi/oE/B8Vjp6Q5Wl6ABkIqc0fYv5sTOYjmyyiBwogKv
+ue2VCB6RL10v5pf5tlbmFOUZa0HRWYijtII5b/DZbygz0mtlLgTXsliWEfbaZiF
oDZouRb6MRijDfUWQb198rvMiUJphZJXJXZoWj8viKBJqq/KX5wOasevkMBiU8zx
xSf1Hk5NY81sMm3+r4rg/ey9FVmtWlji24XHDwCOucrDb2DuCkVzEL+qCbKeNIaS
LZr4deoAsiNlkBGxx20wekZ9q7V5sTc6TBpVfCTYw3gjZ4MUP0akK6CIyK3gLeSX
z65O9t14/olLiUgQRYXh2HabpT4hAs1bYC4dRN7ZHZ3M2lnXlxQRaNQ30Boz3C5H
MmX5KsDMGHD9LQQfqZrz6QrNigUwLUefBNzzLD4ewREOr0K3QDZ/IlTJxTNad4uN
qEIrZATUW3pDDxBWzqpY/6mgClendblqlaMQYNYJ+OsgR0PvMB2ZXaxh3Gb5g7dy
VCLBvHyYgN5ElwCsWbdIBij15Os2fjHK6BXAz0CJnHa2WkWdLeMTtwlSMGb0HAbV
PYAaXvuJRjcSehEqBjHK775Pv2ieXG4XtVrEt9UBykMlxg7rqcUj5ulZ36i711fe
ObbUk/lwVtMTPzL6j9GSRNng4xaatlqOUrDC8faCzeq4WUI29QKBpMgF7hK8cs6q
TLmJMA8Lr2dJn/xnJCf030I5RBUnFIFKr0CStBaEylTPrN4Xv77x596n4XKY+f5E
UekR3vhL9VQG/JQa2GsoD9o4Nw/IYAadmi7hB2ISHyd1SPTmoGnU74NOurO2Vus2
YjIxkEEhltP1OEld7ba8TwoZgVYei3RPGkbVYeeGIU8mmu1dztxwGtsVhZWBWdJc
QIQeliEjpbXaOknmXaFbH8gI31lu0jM/YAiIT03HUTH0IhKObFMp2h5cfG4cRa/P
VCikdNSI2ETCqBG86AO1PjBIgsJFkZgZTVzrsTQkvjwkcgxecRf7IGbTwobhuMns
oOgPez6w22ItvCWMD5aqX+6V6+XtUdqm/t0r5tgxd+1DkaUm0Hk59OZRox7m80Qf
D1p6jXJiAtMuBER7ND/1N3mSQOUJ2DXbIbN9q5keUBEZLq3QyQw2Uht8nOI9ibUT
C8y+MqIBDZKvcw1JRSEOyaaoqs/X1MPcIgYCqeUw+LOGaCHdJ0b7XfDgW5DDmAAy
JecHADqS9SzTvteNZwRw/9bgfh4NuR5jnn/ByCcVNPDn10figEm+4EXJtnYe0qPh
bc7LGtPNIn8gG7Wi+HnapnUysnqX4QJZZw2jLTeuLhxpD5up6/j2Muk0zSAVXmqO
gnreOm3a8SLPCkbWsImYBsfotpEp68jgbQ5UnUhF5AcyCIcJ47P7wk7fleXt7Hsj
AB5sntuVqFyhO5HDwHtj/0HDQiOvtbLQ2XnedHKqShZleHDIFd/kIgK1AH/0rPyL
gjodQcwt+bywyE6FklHIsUBUXIgvnHe+1294q83xucNgLEqoI2th443xVzVNCMlg
fCaA0+iHvdFYPpPvwf80XVrhRXTLla1kPfYZfBsGx+4DtuhhbrCUZZ0eYp9MCCkY
Gt8geyd0BWxmSLJPUeWZDSWlIE63juecDtqTpF7ANY6YKJNedGcbBUbzrTv/OhM5
pflZubKwkoJm9FCx9apZDzgUBCsk9vMFKQ/3k4l9ZZqRkl9dQwWroGbxtEsDSwEH
9woRORTQmqDvvpWeMjtJ6EhLtOTS+FUJp0hAxS7M9wUVDlIjaIZ5gS05oU/aFjik
QfnS27FZuum3o2b5QC5H0g15sfzkenBVSI5griYPB87oVQYPR4IOyAl7PXFEh35k
CvaQNPy3z75SI6zCtEhkKkNHrC2AL1QNnTODh1yB27IPsSfu60EDB5/p9sKnLmGz
AimsKUIARux+jn7NhCDImBlrp6UJSk/07oqJnORLQR4nKZ1mpVeU6bhHZ+Qk6Mws
5CXD2PwCuyERzyzfz5wqozpGGdmb80mphKnjw6maHlgFpCEi1QM2aEgFjkTFZ6Zy
klhaaunMLPBIdqniwXtEdbQMoEW4Gpt3eQesmPKcw/U2IiFJ1Fi+t2QAdW+Wi3xc
UgKQF9eYq5HAW0IZUIFtZ2lNAak6FlamlvLs2i+bDNRQj4Rntu+WLt1yUhkgI1Qy
uyNWTzSfDLx+dK8vRaXYUMATGmr1og/mUaqpYZg3h6ydYcwJNIUw1/iLKITBihqN
W4RSHYfeqwlJ0XjlX9PkU6vQR8M6C8V+Cpc0R9h2/OWrDmHR3AWeafdrhBpdhjue
mbUOx94FtKPVOj9bE2KJ7k/V42kFfBXfJE2JB8s3mTICR8J0Tr+BZPdqHG0yDBVw
7VThtlhnfmH1mf9wZIk3T1a0893cy9yQNW8gTAup5z76dLfBJO3+rSxF0CfbwNK2
7Gr4gnmCOouCFhyLOUsJ4YOoVJqx6QgC1z6DiJLrC4Zz+qz3G7iOO3Kn4G6aFyTW
K57EuZz7sOVvcH43x9omlFSiZ6sq9CbhZiiPmQ6f3A/MPepWZNjVbxzFQiXiWDOy
Vva71RDTOER8YxC6qqjrKe7uCci91gvoFpLbBUbONdSgFBsrCsO8joKidW4vwOP6
om8D/TmT20SEDx3cRUgN+VPNM0ZdTV8KVAzAlB87REfj8oIpJ6gc8OCoMp5lleMd
+dcyrxcooz8HpAcNpMNa8nwP2tuP6pDm6bxzP3InCgsmU2hWbMZVARwzoXkjHgJn
zYuj1aVZp7eApD08f1Ym7dE4KMaAiwZEdf4mIKTnl10RpFJunOdgi6WcLtFk42fi
aKU2afG3WydSI5UF1vn6HqxEYXGTWQGN3v4g5LW9J5g6x7s013KiIFHSSLs1UhZC
UcpUB+8hep1q/FILqctY0a63a/VbonB7/huYFyV0MhfGAVMM6uHS+Dz5ohHvXW7P
j5VSzdskWIandy5jZI25kf8LHTYLeNLzgIjDfyO0YnMydYjyWR1j2Tc/8vVrAtpk
Bw5nsqjNYsfnQe+ruY/EdB2/BVj+gx1RFhEX+7otZIzgRNAeLzX8uTTRGxnHc2a2
ExbbMroqxidmRHIXHSqG7Sa9fHFJRthhmbjv7adYxYDXK+xCv2hAZgL8hjvDmbJD
MUC5mjkIeJ5a+aLstVExETLFqPq0e8js68LGtAD+2SHeN4SGd6E52dzBbUNu2moD
Dymr87cMb+jFGdKFi72pIdHI8vRY7Gyk1ATtWRUN62zoA4vnfsCiRCzuI5UJ01HQ
vJU9JYe8S7sdkJNTTzr31Ob9oMkzNgeJ68KxKO0aCG+baKpKwQ0wsn/GROjCFeeY
SSXXIrI5lu3Q3vHuGH4byogCChPp0VDjDbXK7MDnU31WMW3TokR9c9gN03KueqGb
UFo29dbAcrrGhm/wtXj1HZb7A7dx081BXODSq0l7Sx67MjNXgHuPtCXb9+nVA8wo
BGrHwKk2IinvsXGRN3dYat6zDzJUWLkh2zwKNA0uX39LkXGlOVe47GmfKxgrM/hp
jNbAEZzFVVbEcqWM770qGUvXmleEr8kPQIRa9lEWWoTmrvLtxpmRez5vOtHtTTht
l4/a75akjAOIt3wv9rrTWwfS0woS0AoCfxv+a6vhkVp4UWqxwyrHj26Tr9tNqDHV
enDL3Kqr46trNbpFPaXigOQz5NUIpoahcnltQNt/LHsY6y6zvSqp2bpiam/4921l
85bp36/2gYCm+I/qYfK0D9GMiHLMQWyMtF25W4Y9ASpbEKIkTqHsdwZvbF4pGWGJ
Kv+npDeuKJMlJKrKVrqVM+xHhWHV9P+FSQjG9szq0+O5N/8rrT3/oAChcGO5fDu/
Tla7Cm/7ia81WoAltf862eSMz4COxcwB4ThFGMc3h5cvkE6Ih+PtEsnjISAD3z2j
qybunJ4Z0MTk3G45j+MWDutivSG8WjFIdww5jvMdOjwC0CIlhUAnnZZGo/7+Vpuj
2pP+hk2BvLWPQs6ltxnO0gYjCTsxw/zGnvyDfxxen2sSBH0HN8Tvpv2ZWV2vcaDs
0YS0P4Cv1TR1Zhm57fsrVdHExccJ7fluUm1o65TeY4UGoZnboPiGLk0HtyukNn9B
6IiTt9+H0VDt9jZzecu9bhX/1YaOM6jChBePIMN8DVCVY9WlwvzwfFlq0s6yUNwb
+7DcYesJXj+ZnlKxbEfm7usZXmN5zzv0kXdsL9HSfYbsAJRdrUdJ/VEH7dz2poAB
aqzXsKUh8w3bkpS7Cr19LjLlYwCFZQjclBD2mp4MVisWSk/kQs3Z8K21XJtWP4Y4
1MRzd/eHiG5Leyk9woAMendl3G+gF5o/vCWdYm7WLGqjWNzhP6d00PyetoWLyn4C
Vyw86CSZUvgSo7F7hSJ4IwoOAj3vspzW6TsjiRNjEg+bSAABLRlSwFDiXcvHU18o
EDk1YqdwqnUfmXHAuit29cnksBv2Z2mehrW893y6tTZ/729z/sUqSqdo0uorScSq
GA+TlHm144RsKjK78JZENyFW/AH7r/adPAhWRej+4xhhJN1fKgVghtrcPfFlzVtT
+LV7Fq0NnAWE9kpkE3Fyet3cybSV0sDhUlqcgnnNQCxwK/I9dGwj+txF+j6B1W0P
nQlqwaCL8tTBt3WTyi7OTo/LiKMxQW7MhTeKkSzMx6M4WnvQQnW4k0Qb7n82L7IR
dRT3ABK0CJ7N1FKBtDX3dVT1wWt41gYsAfg0fWhSFQCxEUeJQCqQsKgZtI5KrHcQ
SGby71h+/OxOJxHso/GG2PStw5d7UtDRYtQ+/CEmtwmvHvvT/VwSeqT90MekEJ60
OWxHUco67TfgaorhZ8sdVc2caUZTR3YtbAu9Y55yCHseYitFryLNbhH3HvCBbdZ+
mECC36xzYQrUDTcBpZIQxJdb3ayedr4ym2zSk4E2zg53kUoDizHqr7AZXrQlFc4y
Kon57y4oEXmR3XtfXL6z6yEVcWQWT1KbzE0n/F6KKlInIOHZ+GmfBQG9TTtaUyLR
LFaJeiBTjvMX96E8qitPJwrfCivPhIN1TtOwSlLKOSNorA53/hAQhhQqJDIXVZof
3LQsfDwNn1Yy1cQxU+NX4pGgoCSgdHs3PNK6ORYNUkf4Cb5epYCurQ1d3chuzJ9V
NYfin/z0D0Bm2pKLSIrlJZT20ottMtv4+NcDKDU0Kzu0uGwUjBF4ef1o3H5KkySX
jEbKtzoAPnZcFcgyJBgTEDNp9PdgJlRsoFjM5JtkPNYPO6jihLGvPR7fTYjxee26
0XSmbtWDi0R/bQPaxFngq7ZkSGPE3Gg+Y1xLkYiecdfvIQTPOSMKx4trZ3gYAA4O
3hWmunH+Jd9+D+rMUiSg+NtXd5v2qQE9hIL8Oc+wQE/0JeJptt7GhksgWfE25hMz
F3sYMfxQ2Xe3jZ2mgPjdl5ynnoR0tzqIJ8M0Ewiw0ueF9+ilNBeSBBo/WG5BIrnE
q1OZIBo7BTqB93KcCfKOwlRXnJOPHpI0/vMFkonQ80Rop8WPoxAijIr0+j2pacjC
924wQ5BjRvpOQyvnN755yrVsHMGYtmrJTIkNplAb+MP7B0ZUUJiNP/cBQ2xc0pkH
QJX8W+ozjAAo+2HT3EpWRVWnow2tEFgozRI08MR1y3/p48xoRiJi/Awqp47tCdup
X09SY2LajlSPygUIqXwv0yCChmFZ3mH0JrBymHrrbL0miSLEZH1kH+cMF5eRKI5a
Gv9dyXPbxoHDmyK0pfDdCv6st/MvUBG9C+0gjn24hAGyB3KNivn1ovUDJS0xGbYs
5F+RmTZkRbE58PhxH/Y9h3aOtgmU5+G1dQfW8NXvYhy8X2wRlgWN3xZ5/pHcQh6k
kgAqSwq1+6jGjjq4YaeR1/fskd6EPs3iHTuH4DG+ptPgI8l6rIPKFMI/ciK9n1ud
WP7Fu82+DIXsMKZB2tI2GUbp06GAySuL5b3747LIebYzCqJ3IZxwEwz3lpgfHpqX
UUXeHAoTrDKUC1LDeDquwGxxNdoRF4/HcoH+nW0QD6CVXrIErd9sQ+t6ef/zITOA
3VlgAMV7r0n+rkjThOH37yiZXGDF+zrrKLbbFDvAuzQFQmy/mfn1bhv0MIXKBJOR
UqqnmbQWdy6uQMyg1Yr7qnUkkJKw/JtiepPl/yntxouvJFtigtt1J0yDcW/g8mRH
T7RWJ4SGo/fjl7JVzhaHdQbvey2MXWupuzzFvHm628v/cLKTwtwwzQKpATIWvrO9
lTzgCUemya5jNkhTit4kPIlQe9mgZdNKUmOlp+e2vvy34gqdI5fc0h9pCW27WSgl
k3DFsz77UZxkFVHA08LkRcohiemz23mOy9UY0o8jxXqcxupXYr5nW2AgbhAmY/cX
iCYbch6Br+XAN+nutHdApFYK9HIXA8MOaR5kM7Ree3O8aXlg5MvWaMK9D97ewze/
qbxi6tekuA+tk6UYqarv1KU+rOvbWXzwzfjxqJffH4FCpAOl5LrGcwb6DziGK0QU
KMtnAlJNDcmCKbWN5S4PSI4QcDzuyv/g8R8UjPNrkl/YZuXJW7C2pUS59MAMr2kU
hWhJEvbEHLmbwL9C82tHZUSYWIX8EW4yDeJnmSVMGPM69NHdoi2fCoeyNcHwCIrS
5Y4QeUe2dZbXh4EaPA3wsl5jWpdagA7tF8bZjzLfuzd9PH198uwT00lXXf68OS+h
48Loc0tw0zeYYky5EWuW6d49MZwKxZ6GM3NMxgGdvGiXzoPakuOxtMir9nSiu0NQ
bMlQ3PziDp0OZqSGvzea1dm4x+WbTMDNu/AxWg+GVDKv3uF0zQN/sxyqc4hXUvDT
gibxonaqCI304bqu2HuEoFeGHPDCaWsmVyu00TslQNcQtDy+FJF1gtMkW+SDBV0e
X0zMCEHFPt8fUHMWl7KINbKMVHw6Lyqb0+mKQXDsMnYIK+JuASKhbc086PDLM/DB
/zCV5fURVUsAk3Ku8Qa62lIoAQhr6FDPoRYU0VjWW22fN4npxsmg3SdZXfb9LTuE
vGQjPIrVoDwMMQmAVtVcEsiybCOA+O7HkI64w3yVMdQrScpH/KoZb7NFM7sI0UUJ
nps6MEAVR9nPZRZ818gcdRD6hgcvTtG8kpPlfrZDaMqQJ4/m20tKlXfk5Eg5ZJTx
3xSG/EoC8fDBync28d5w4fSadMM4mxGA2qb9DfL8z8GFXNvofdZgmJ22IX/ByVGx
HzNBGH2pUkds8AWhhVexAJwCq7GwoUpBWLGMvXLDsg/LY5AlKQeNNn0Gma+vBt0X
r+fopyTH3cyNUeRLl2M5sPF45He6O3X98P1UVmejoNDmOs1359zDlsZuV702Ze3I
u0zopfseQwmXn38/AaWKLQ0O3jFdsrKn1DxvuL9dwC4fw3l+urgQ8ubb/rsMINmc
JWMfQ1qPgKijklV7ZXqiyNZ7n6O/IB50mAZD1g4CMldHKAAlQQPpAaZ68FLhkHxX
bCINp1Sl1GhG/5obVFBZGVu12N59RKDXAZtzGAX9wcn9iHU9STfCxtd7eKYj+Zlm
UKvxfMwWudoGorPJSRDsqyE7VF0Ht4ZTwLtgqN0AFgctP9uZMHF4W2LMDD3iQmpW
7KpbjZQ+4bE5cO6mCSwUzGjYwV0beFNkeMTRYNyQeVlElM7Zhb5GmoWup7Kl9J5T
nBj7jd+R8Q/YAEuj4N4QlKHyQ/PYND9Q2rW/pAjI5w1ISd3bnpkRypX6hpPLKbvl
kngMEYPpVgJcLizIhcevgTOatB1Fuop8SpOQ2n2Wn1bsuZV75FEhvvyDKqSDVIX4
j011wmBr+OlAF6BVXA4PVQjuDpkTYn6SX4Yn/ATHyZuqMIbtZhP3XN7nV1rjHl6/
L5MEpQ5pdjs1Ntuc/IqkDSI3Skg8tdRkbu/5zh5oY6/biZ1SDSBMY6+8kAcA08VQ
IQLq+F3ij/7HIXC8bK+sbL5iFkEl1NdUY95yJb0K3+J9MQQMFVV1KQCwDjJ68kCJ
zBfvrdxrEyHGN9tWUEjgOd563SoL6fnfEy4GpGoGPDXHCzGt/h0iJoFDJm74fnlK
+7cc0Tip6uSCbwn9zpV5a1vtcEN1sb3VVI1O2sIFlu0tl+JkYEIOE5d7ZTWx+eXQ
uZak+5GRok1bfvJKyZI7MvQxvUc9O0YwDN2rY91wJ8snANAnKTptgMmwq8Qw2UtY
QdNsS1SnMq4PUW9uVWN6/6l5CZkyrEHanaf6ylpP+oCGA3161HQBwwm/7lwWzBmD
6v2CxhmDsGMM/5Vm740h6m80wW80jcUmGgRvmXoXGqwbvdAsZ3UA6Fu+lLwBcVll
38AOc03/8tCTV6Gh5Yqdwt/T7Rfpq6leMairlV6lUHy2D5vm8sdS3SdtZskBqbwV
pd3C/XzdW3tyykWeSEbMGhLlJQaB9hCxFtzvdaLdZBOxwXNH3y6B6T8bo9OaPhrL
ushyMZ7j8tFYUUGk5kia36oO0kmTf24tzczV3rUR2Fs24U/62bO6dgHPcYFdNmbe
4Vh4QMF4jzuwjdpsVviD9Ny0vpJkVZxm2o2yo/YjwRbFR1Br6J1vFZCd7gkh9XQV
vSKVQ5UpTjGZJYeU3jc6peGV51vsr8l0mAbEwAgKGFbnkS5qHCV0qjegCb0oUcRo
XQWmyL3i16FVltFUYBtzFYckzS6yZYPgHvSkflnrXI9r5rk2nBRz7WtZb47hd2n6
DZdOD75B4auGYJB0wLANZo2ZaC6OEnwEUDR99qSeTvWkS3y/ggN9I3cF5Si0OkIU
i1tYpnES/twqEkDwi10kDAnZf8WxW5bHI0W+jVwAbX46Bh0UfX4j4uG/VJa5up2i
Mh10eAUTzsa6PWit5IQPomZXx2LCIJdsxNjShQRSk7njXGOFTTWNFQui9FFSkb2k
c+sCYRP6TMmCzCyLQtIih9ADdsm1lyVIoTxPn8DZ0dzJpcKLRUNBOxGHe3IWILPF
dAhNiWYwiuuwS5PJjI66N/WHjLAWZ7CgNVoA3C7UUZHQDRQA0Zape5xlZlebKvZk
JW4dJKoTU9bc9vIi5YdPlyeG8LDFfo4F3LZ41AXcJqpOAF8mfoJrxrJKjU6Yle/G
MKsGoWGzTaiif6h+Reji+5m5+ZevLkHa33mJw0l7yQuExRJrPD9liIIZew8p/i7h
a6VSbK/a16UDwhrX5iMRjWrlZ6OnFa+l6ct2sxnknQsA/r/NEYOkssDtfKQKBWpx
jVZ/DOXASnKyCuTonLr7e8d2WEO3mgklhywAN4sKmC091U9llLbyyMFehmc+8vms
TJDfSa5HMYIaS4EJzfcFTMed+Al7ZRnf/tAofIUCjw1K0YW5c8cHaUZi7UMCqovg
8iVWYKhSS0ZdMKPg7hXTADZ66IDgqlYQZUfEjRRkz9N74HAtC8qUc86d8VG5pslx
x3XqckftE5+llSX42n3JYpAU03x2FMLViBX8OtDgD7pSzwskzbdWqqYMEk9trUYx
Lf8shppKo+TA5EE94bd2/VgmoqssQu1soKL8YsERzVRhGme3SGQc3uijL/Muo7nB
Zmug3P0Tk/F6BFB0fmR0dXHVIO9jWN5JvKNZU/ZQBLLaXU5maNPNnAp08krWpymf
ASCR14lbQ0CzfKp0VYGmGUl+AsSjcM7EP/Gl5Gz/7zywozzcbd28Utgwwehi22VH
i7pXMF6P9UZxCgiqDMXEYp+AZrHgwxMxZNu1EHybEqgN5ReDuXPNJO4nIerwI0sr
oE0OJKX5VUbTL5g1kC51FCbKfmVChQjtW0COnUG87mXgGX/U1eErT0Q+nKQHmnfn
aLnwSQPc4lE+Po7LQLAuXWUoq/L/q7ygLN6u1IvDFk5i55TgUijKxfMmKKmSa00q
iCusLiXWUGOvkwGvNCEiPd3LZvmvCSl04em+8lXfcipdIHgXHc2E8l8Qam+TWPra
lNMwnEyBqjmZjK9f+ykIwrQKnK9bQBVYJSD4UKt7JqNhmqiX3oROnwIdMXcHFI88
HukKICqURsss45TWbMhsHnpPvHNDQEMsWC1hQDDjxggDD5OnEUwL2uduqZrtF786
eps1Zj2riwUlQL2Ei5ubWgyE+Sr8Y0GdJ9u5w5QecE0tWTWQXLfHNCWz4ACymqQ8
OtiAjZklgi1go2HpjMmZVTztGShJiwHVgc+/XwBaF5SpD9xinum/tGujkdK6DLY2
ZzdiUzxwt8Xs+g6dl9kJHahBQF3pI5cwZ/hmyosaWg73TXvT3E6oXRRzCb2wYUjX
oRFX/+JycM92+EHqg2Bb17QPU43vhIgO+7QpPdpK6iTUHVUtwByE1TnzJaOIYsKX
dmRLzMlydciQdHImOz3aJgvFjbq1qy9oVt/buyp5X+qkDyuiD55DiA81dM+RhlAq
sYTroyoh6k1dV2JXHU8GQaeQws0hi4AV9xjF+xWzOTcXDDuBEjxQ6REBcwNftkrf
sLdpOij/yM2JT5T+JbTIWtd5PNXEF8jD70SDNBj2Xi4ncTx0kJTTeEJtzyqAm1Tb
g9ES4MLZUmMkKOLOxt92092HUsOxXiMuSchRO5PlNvGIWFEr8fLeSlizKMy+OSvP
QXm3l/o4lE8ls+umBHkELBoopKhBty0SoMZ+4SzS5/O1WF9RE17vgOWQsB0AQ2EM
8Ou9IRPdyIuTbdUakjK679xADRnnGcoxLIqnwf36FMaJtqeJUU18fb5oK4MWXL47
JnIFhv8Nqm5SqWNK8Gjf+XLPfRH/VzkZ5QyibNs1RdEf4Tqua+IA7fpYAnxhVPQY
4mKZz9j+AbQG3vsxQBfxGi6INnpA3NpH1Py0oJJwCbbqiN8ldgnKnErki1SmOzi9
tSR/dTR2Hz02AxMhGCErJwDfcLhPRNsqPEo0pi/BqSqcVK45Q/GBJc6acYsPCeYt
Me3/NPwabtVcN488+YqfLlimfKpbhWT/5UdQeGmtUjmVI7q92yxEWDGNGGwCm9ey
sOcVxWiEzn9vW1s7BxC8oqhOdcXcKkm16hl/QvjwVJdv59Wo1bigLLGQJNKZXubf
9BpvqIfANTAfvTQ54qkCHwb2qr4E25FxFr0P9PJi0cOGIzwtkLtLRrQ7rhSJgDt5
c4cgI9HpoBFS82NCl7BYM9HXfyV5wi1xOPQn52o1e/reuS9DN/tPgt54Br2fNus6
my0JLgfR0neptSIGvBYlGMXkH6w0UYkLVsFizzJMIzF+z3Z3gF+jNY5MHj/Rh+D9
iVeBtjp9bt+21Np8tAKRxO0vfMYBPdmDSSLt8h3wNxqD6S/ka9bfLMHvRmRHSHuG
g2U4jMclEgHe4OF3EOYjxDjNyDL+Ip7voFnzig9nCv3oIoNjPzsGE1wwp/NFVlrU
aeosyxuJSW5oStWaAJhOmdAmq3E98Adv7LqctLfKRKmM2Uc1DgCINF+MMZokkjQb
Pf7IYdsdhnvv2z7uTEfeCEjcmbMx7LH4oeUXrs098dSmkSuXs7eXOCaqAQqknU30
VO+0SZrX0xH/5mua3dXbMHBpoqZrppUs28zlMXsIWX45HKqmiyznl1elBcExA2fp
B8j9iOVU/xPXFyXSd0EHWeLekYzZYFGRWQ/LYf31r/dxvqkMldrYDgpNkINW6Gh8
lajGPLHiJtDFLnjHkxk6weSvCBhRKb9iKkDFRrYYP6zsMC0R5SRtY4Os9My+jcq8
KHoVWMF4MToDcELc/Pllc7eELJajvzdMXdeQFbWcpWkw19SINXy8RmaIcOAUtTys
d2ZF2KugAIDqx9lLjhDGT6UPyaa0K0fUtm8hGTGETWZXUuV3H1VgllTh3eyH6JvP
kAM/ynLvVRQCa+WaMYg9vQhwZ1kLbRpAxkYnh80nK5MbUpxZpwIBKtO2AqtQoYJU
aMHpoG6dhLwG1Syfjt+F4LqpdFWmmzCfxRn2qmg9X5vnAf2wgRhWRZQ1l2yBYiQn
K89lnKxpWI62T5OUEgUImwUcjgBCkyvbOcJnOaK6kGnkQag84g0cqwCrm1l2GsGk
vxbp7BINUVKTNINBjNK/al2Kn3uEeRAudOQE6QUCWRkbbKVNiyHVSEKDV6ZV/OcT
9YxqunazvhMT+DLLmTKnYZnTH5XNLJMKGhC70w+0RxgZavqoCmUMYRwVwTndcYrI
hFztqF5vjKxIkyujxJ6YGZTGpY5/zJ3Y0va/cI41c73OcEF6YrEye4cStzO786mL
baQRv9DU4zTBqNHthzqFyYF/WsdmVEfBxBChA9qTz4BeZFMoT8ANyoinlCGAr6ef
PPoIO1mc+L8aVXrSRf3wjFWFGkkrcVW9nQU8OwJAxImkD5mJCz/KtcZYCKGeh9an
v6hDEtU/tTV5vcwJ9+2SVnXrTgsOt/1klucsTd6TndvOMbeOFQYIcGLay1acwem2
3RpSxoSj/eAnGgNLpN6Hd6n+2doax/Mw6LPBuQ4KjENst+7flFl0p7HcSk3YdocG
VNXICs+c8o+8l3VRP/ZDZqqZMFMzS4XbEVWI5fMpwiWJWaktHiJRVQIxhnmsGp8J
tbYD1L67tLEd8mjzm3WIVOVz3PQEyzsWwSar2aI8rN3suEzmZxMdH7U6x6NU0HgQ
debP3td2FvjtW3ExcHpgAnQID8k27gXbq1wx0cFJb+LS7/DMOcVDSAU1xHhaomqY
zGsdFK6uorFPKlDkvhKLjpLYvPTdJR8s7xCJ0CgdDPXt6kEG8t+xHxdtzI6+X9mn
oJ6kkgVMKN2XIhEtQy+GGaT1RiwLEfyv//5dG7jzK+f8X30abzCgzYwrbMS4bPuK
dq9DA+3KnMs2IhSxrhrqE+6+j08ehFh0I9KPBbRUFA1uaZqDv1ZWlRvkIFaAYseL
Fx0J1QJVWzDNRMiGc0AW0Qi/RZ2DatrG02QX0VA+9YpeWaIoBRAuRw2w2m1FT9RP
kqZKoKn5kDTJjs16U18lYzj5karK+nONH9x1XOYhv2Bm7bFFZGQ0g5frpy6nGZsa
wPOX6KaKkxcUEOeLcptMGXm+m0kOYviBYY7H0EhCr2lBy/n3U/eLGXnwN7eGO/c8
mDk1MrXKIi3pF6i0A4ir6SisjyjC/lKzmdfMljmOR9FWHgWlLCQyJxf+GSqS8JoR
rx0/LP84LkN0CV3Yj4KDSzLgfFtopPZVxk2jVpLeHt2E3QrBZ1Ti3D7tO0JGrL9K
2KCFt1vK2VCwj2F++t761ppxquR72gIUZrdU5Qfil+bWyl4TgZDJZWLPrItnquad
tSmJtXbKgfVSkAROXpC6XG2py9jgXMAgGAqXUYXVsbpJoOtIh7F1rae4PYiZO1wz
SxuAQSnWz8oKBinGi660D6OjlnvL4+4odtZsRBhvsbd+8DxBRsNT3l6rdcmx9/O2
nUwfhnFWlP1hUfVUUNsdEZHU5EmLyDIiiszjkD/s5YyDGzWR5gf6t+MeMey+AYJD
+WwtMAy6rRA1/sa6m3Rxf+3o8LIQi/sdZCU9WIG6MntoTyAjqgCcVdqMjDk/sDnE
h4MeB8bL1sZGp1cXmUMYqx2EBwzuxSE5peCyiX66UzRuL/RiDujVr0tS+wYbzBjM
gTnMnllzRVdrymn4sTx3cRuo0ckmxYAPnvgB5bRPsxyXvtf8PhE3ktlt5deElxHN
HIyzFWYzsTiuKzwqWO5CTM+Chq84JwLnkEGms0ndzK7IiJFrqn7lKa8F5b5zS6ez
DrxZ2cfEj2DBieSuj87EkONzAWHZq5rQB/L/GPEF+zw0RpnGAveApi+X+GkZg4Yl
Hjs28oXwJLA7I97zDYuzqYnHvNkvuo771a7LgQ93dcfoAbJrhFQevaAeYKt6AMAa
FtlDuHt27VRwIPW3Vm7vgKHtEg5IJyNh3PyEGEWCoBxd7uOUxyXqIcT7N1rHwG0O
ddkGXdpeqpbh/AcC2YgAxRhxyXf+0DYwenhOmSpSxSGoESW3kvjM2EVhxebSrrjr
goCiSW7vN+CSyh901A7B16p3N8yxtr/1RGNjFK7p+t8DoWoSjnNrxTsOr/DNKuaM
HMSzu03r6bJtu3ZSeoS/fEabh/CFxa91x1aaKbo9ue1rkLc4DPtuwYtCBFBKn6tb
8bFNtJacvUSVSP6zAkU84SVo31HWud5gWCZIpTRFXFqsHGdIvzEItrhiFmRrLG/K
arBWzMs6Lo32d+kN68AgM+LJRqEuVnhfLhbfW9DJ31TUC89pboOwMVcD0Ig288ri
9iH+qhgXPmZ9keZx9wCH2IuyU7DsO5XPr17SIR2vjoFTXLfWPDHepCq+CEhahbiG
2RQFp4D4pLfaxUjjIYpqsUW2uI87dpfhY8d7umV7SzOIKi22an8dnXwfSjS2J1fn
qUSjz+qnss1NdJw2DEA4kOoadDDrZcMMKuqpCFzKJY3a8e5IkKsgWpWiR7t5sCEf
gQNL5KfrTr8rjl4D81gpDb0Iu60P1p4zWsh5L+ougEJy5if+ld82aceOkTuw9RXO
WD/2mK5wbsuuq0VSA3tQM7dx2tnh/Av7L9n1Q7U4YooPTjHhxXG8G3YHYCn4gHt1
QSUeZZykm8EhxiHgSZmf9UGliruXQyXHv2kD5HnC+4Nwnbmk5uxYDkiVC0kIoF17
5VEdPmganpcYOpjZzobv7oScgVTVd0yTDvoWzwXmDukyQ7rxIVknzKzvThzj3yjo
+mK2HYsvbGTSeH5W5WMhgI+EWbKweCnrgPaARonXqSA+36YoxgKZ2eU6ezuMNSh4
CVte0FACi1b4MDRvW3cTuTNiqArzX3Sj/3JjtSKPYEM0/S9d8gOGHjNO5rNryW91
bA+3YfMZgfTvC6TFTie3hmtwnOe8rhC7cOFmFNnXZHmG1eB0GfNxXSgvnsQv+UL4
iOqHuz2d8GAvz/ujj6PH4+HrOgU2CufcNFB5+6zfEZoGMReWwal61T8YBR/1Cx30
bjEe3A5YVd/PxAtyE4aWBl9z0tu2u0FbyVCSSQJkD3xwG2NLYoHIgwWTVYVSqMws
wgmg2iFFv6c32XuF1kSIBz4eEBP/8uOkbrwRxdSvukSnwDtpQz1HbVe6J1ZMKlyl
DJg5qOU3FUtFTcayKsWsdhgD2+c6lz8wLdC2bKW3AITqdBm9S8x7hNFZpJwUuJ66
1b8Mup/jBS/2La6KF6V7mlwe0hXeCj4pJ+W+/BVBYKO4z18xwP/+QDrhuv7HuddR
4j6u1wPOpS1uNJk74/4W63LMIghjZv6pSReWIDT6i4Kfyt5xaKWj6y7q5PFgj+9U
3uVvReZABT9TuECmAejjsRP6mlHE14rU5HqRBi+MCc5dmaQfUw/Kd+6EmfbDBRwl
Cf1QmZhdfhs7+ZimXyuSUwJQ1YkAzYGU7XKfEIsDvvJ+4ZCyF+8tpu5eaRuPYQPX
eMy4eCwhztc7pdWks/aXRwjBGbPRUHDrPl32TJMjm5EdWd6d/uec2GMpdgARUx8C
MRuoSNqjUkJeA8EFrAnfLV2J9i9RdaTyo235K0VxIO9RH3BFd6sumOp8wxXPX4xJ
VvjztXM/GNy4QC27d7Cb1vEW1IanMu8iH1+xRjTHThYJGU70Y88IGjYIaW+YtYtd
bBfXpKrdfL21Cc1E/YVkSNWVB+aTMHqOaayUv8/AexpFKpMA+CPrzrngZt7ba0rP
dG6MmHFNERtyDwl/UYsUvdGK60kjEWTiNYPB3R1LnUgP0+ZReGWTl69/FwCy3ZSi
NjF73YzSiz7+W35oNCemkaC30TVKoX7LR0UGNmoTV5jjaUtFwoiwNtWPabbqpqfg
HXr6Jjq//d6ASkm0sF/N6Jyz4/PbFEbVPsvDH4oA5QN7BfCS9IGPsxBVnejId9+i
Pa7SfUJ+Cgp6Kss4dnFGrHCudV9hysKAVHhwTqYpKHYnzUNYDH0xX8sIGY37aBGf
YznZAobk5chLxxDqJquOmhnyk487sQS6HA4lErjZz9Ds/1R9lo+TbJgfbCyjsRo9
aUyfEI4zTtR3DuPuCVofim7rR1CM16SCZqEwIf8KbgcKSgeUcxNc7neAnnBaUfir
w+vJigF3X0sMc5vZKdG09YzLG5gmkOYgQtHI5ZjDtYKLPV30F08vwMNCOUmPATbB
LQ4xCkkFOdemlydeBtvyWS41RY/SnNXrJPmF7IQjdQThuduR7JUaZinq7B/q+7Sp
Jz5/sv2JQaS7OOh0U9Dlj+A9/aGyF9E3RcQ8HdwIPUQgRB27jvrTmneb3M4Ci4Z1
rEpMDdw83jRRPk7OqeZcbGGz9lgzXdYBQT3CDNQDX+EkoiXxU77qLppROS1yQpvc
Ji+ov/OXJ0D8fOqgVBachk0qo4Lny7K/tvwAW8bEKmSHxbagSY3bZxD3mtXc8vfJ
yPXGozCV4H7D0UqquFo5cS+watQxN4OLNxGkwEYew4T54r+MvymExS3NKaWREVLG
cDv9+kGB+XrBuY2lMCrgEvEiBAzaI++dF54VfdBDt397jKY623hSqQ/c835nOn7y
VfRI96Ug9VMTB7N18womcLsfvg16VN5OR4/7ApAnfYFjfz7Rcjtsr/aC//IS7Bx9
wX7LDpwmIQqeQsEPoOIWY4DmZsn82EyPKmrO40RA0zudwyIrim0d9eVebGfgq0nT
LulO6ka0TdEDHe0AcSqjQVO5MLwcW6jOxq4P4pMLLwVkbAR9ZChtdJlj/jQUAeqs
yVyjxONeyZlDXw8zba61NLiUDOFLxurwfohB5so6GzB4SwhCcaT6qTbF8Wu9kCpO
HFv41Z9PqrtDjUt8GUoZeV0TZ/vHxn1mcLxO/fCo4EVlZXNMVw8IsIcT0sZDeAxF
dXfx8G4BC5k4Bwr+tb6OEHilt6MR74SF6qkysw7vNI3MkVnLI3CXsqeW7UtW/dKi
N8j7BUk1ryAIvszjQCLKGAm0c7569YN2aL8FLurnIb7zlVLXsdO/8dV4bsfF+huv
B43RIMICStOIOVMhAxGn0yQEcmIe/rIN/lygrj6q2DAOIdpLRo4VKwflhKXuQGyx
nHOiYv0H7NtOEDhQWbE+ob5E0ScHDojXbDPW6U9i/Dbi5aFDkWzRJWwHn7vsSYKt
PFtQ6HsAg9O7yKTGXpUjFwPaSpIONOg1qiFTrd6b/ID8sAzFQ3B48qLDpwwqwlsT
qqJjURMHO6wUV3WsAAfVXeMXxgdOyMhBVP091gGBig+bkKnwKK8jPvrkdMn7zcWn
o5/OafhgKbpHHhRInWerKxRrbVzDbsgBYtpD5l8zXamhwvu650C84kdyQhd60Gq7
1O5qaaCCI5ubzerx9NSUH5SdC50MnADyQY9tPDZR1FLTLTroT1hvMJcXKbvhJmVB
pv3dgU2qleGdMp6w9s7d1wtLY+StqGravWjqkAKHtAKnDLyJo6vUJt3iYJ/jzVP+
xPy8mBO+Zqvj0pNq0l7iYXm1T9SigA51aCxgfKIZCHDxwfcEfvDx13kdvDDF5ULs
2WksVnZW819K8ILA5veTJqnCORh1lwocQzwKmNYBh1kLHKK580tsHMzveDlJZyIO
iyhXz5RO/JSipQ7u1gfjIGfGieMZBMkbypaw6t1bTvMOUIQdFArOGZ7MUajI0b1d
`protect END_PROTECTED
