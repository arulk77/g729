`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM1gvAyOzhpNxpAJu2d/g5ownmIpLplm26CnoJoFpfml
aZcvNDvPYHvfYiM+xcdwtzsAK10mddWVOAkN4nEqpA0Sgs6wWy32lICmA8NUVkQp
xXBXX/gFJi/0IaXyUjTD1E11Aiig5NCd5G5ydCYEhEhLTxV326A9MKJDZQclt3G8
yrvmKYV1kDKg9h8aBEmdQDdjrIXAoetIHDBxg1GX7uY9ODYVfsnj9d2B/kPMmaFd
mZu9UCxAwOCwlAoElYZIaW3YA5wFxlpfjCds86TrvxNZgVfK3/XdSFSUOSW1kmnX
joF6X8LHBueedJbEaMxfCWRKGtphYiKV6N9NmIlGPQLJ3URsFIVzQi6h+Fmbr/T8
FpW8h5xhSaigr6V2YvM8+qdrZYu8pvPsjDiCa5W+nBw=
`protect END_PROTECTED
