`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40YJqPNVmihZtJjiiQiDNkmTXS4c8n8WWDdcKH6bE/fM
wyr2KAMy7cDoKVn8VtWfw18/BBL7dJ9A9C8IC7DNYWrlGLBci2klFI1SdRvE+qdN
XKGYLT0tFz7hNNcai/GeJM1Ngb2WOQvYd/teoxBbmxXbQAF8iEF9jGWYNr9DmPr/
1WWvRRWq3MbXRTRBhJk87K/ngtcM1++sDUTuvrM6XE0hPD3qVaLWJjiabKiqve1o
ui6YPmmhK4vSbIHNAyCKdM9m3JWb/+LdyudbauNCSVXd+TjBqYNBbpr7/o9dhYSn
thos5e+8RTtUN6jAw56dNA==
`protect END_PROTECTED
