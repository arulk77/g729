`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
lvx6KDLQRXIsuM/b1IqqeNfiRjpIydr0KMPXj5ypeGRn8XfJY7ZAgShx05Y/J2eK
oKD8fXeQZsw0/+4BrMcnG3ujMA0LZ36yUyvqJrFGN3JFis+wNIHO/09yC0Os3TmB
+DzPWtdc/Z0suZewKQsIZmnnP18rBWzV82jceSwOtAzdprSW5nTAilAKXu64AyLh
QNy/KWyt8l8oazekGVPg5pyaPl/DnIptBTf+sxDMxR/Mmh3K+C5W3Mh4Ac1GWMer
Rn9SfPpLPsmmx6VPwM+e30XHI//xjquZJ8ZPnwIF8fWSLE51LVh5/C7kNt1wp/lX
fvVo6IUNRuUILVIjS8DCPtNrN/BqVnb9O4kVx/8XmmxRJOhoFIJW0BSArV4jTP1v
rcnwflg/+S79FRfgSjXcCkzwS5dnVUHlUOxrHtKAKeqUbQ88xLX7U3gvCSfZa2gM
PEEri9kYTloOMencb0B4nc52sHM9y0i3VJP8nGpNRDJB1GTt6RyvdaFHQl6+isdV
N0WuTbV8omG4W7pv5g6GEkrGI+F8LTLQ82FH/OO9d3VJmg1rq8PfJRo++0JvvlLn
RRSQ/id411ornNkrqXaBjfFTtWlGRuNH+kSmppJv+XGa26UeIjJ9BVZ6TBaRLo4a
+YppEliR7Lodoqq/8DSZY0Aj/Y2w0f4DkgZdi4QD1ZbDP48fa7NrsYo/qAx1XgE+
IpwkNq1vi4kTZJ3tQ7KKJwo+najYfxld68MWdVqQVepKggxVq38mebvyViLNvUpX
tubhFa8geu8hz1H7A7TOmLAbqs0tpcwiSVdU5hiT54d1P0cqb1gphnlXyApeVWJe
OH/c0AJE9R4uG3kvmnlXhs1xi3sK07y/+P9NYN4qmLUvQOVZU1EpY3tKnzJmAu26
HMYn3hGz1cC/bBc1o32qfUTwBNqM/j9AwHinGHohWns=
`protect END_PROTECTED
