`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C9W6q3aHVsqTdTXR5frG9j3gcGdAc7VwrFE0QsyZ4+ug
a2Y6zWoNW6jj606QGuSle8HuTdB83THbqZBGgeXg89AdPa9RZ3OnJ9o2KdYnc0vR
KQnJaeMFJCyPfwOGqyQ+cjWsvjOxtkWdBKoYFyaXwzhAUjRhyIhxsd0FXE6mPxTZ
MpZY9rkSnBbWwrKdA/Qps1FVvyS8I75lG+J3MewUspSpzNIf8g101pn9rHzYKz3v
UXIh+h3OsVCxkUxCG+4he/LZIJSo5pAHmb4jboTYLWOYArM6o6xuT9jNB02YbHFH
xY49UAiZH1iEiP1xBqMrJ3REgEmDK6gM4zrNZp5J1OCLcuFsTVKIIBpBi0o7aaVr
p/RnPxQ+B524QNzacK0sA/A/huTBJPtQ5bk8X0/uuQHOIt5nPealjfjYZzL9F6tn
ybABKW8BLC1l0Cuszod1GPbdx5oX3/Sho/RhqAD6zsAM+vzjhCse0yK8RvPwDPoi
iAb8ZN0INzhxHTlqiLMAX3FwtesyV33PD6EcvtEIpTMB+FGB3+0E8nqjmlkOcRjN
n8ngx4Z07bAlTg4eE4bzkm4i5Xv2VspxkR4PPC7fTj9orEOSeJ4KetX1/chKhXbx
JzLif5Dl7iykjqhk/P3WkS5QKQ1t8oyg1R9DuWmhNpOTSqR6RQ97w0eh/Wk78YG9
x9f+YuhIYFpb9l27+3k048XHIq/g4tfWeXQTWfdxqH8OqtHORlrfeae0xd/sJSIN
US1JMFoU+cEIYypxfZRbJWSznZeST7o9mRvg++zmtkUpBkHJFSQH2Ev/Fj+8+FIT
M4B4Jd058Lgn2aHWOd5a50Wc1Z4RAbMBZq90FZ/ygbEgwWL337KrsNPrw/gTwqyD
G32fJ9in/s+gMMArC046UImyCINjRESdBQ9re4TM/lySvQBcR3fllVUo9XSxLD7a
zwlR4i/hgnPLr4rINQTZeOpquNSgrp1Sm5mWsvgGjiHf+5SOOk9H05XAo5FaNjnh
xcQGhgiqLXjpEln67RSgZcA0G4CbLHwbFJKjPeVN5qsjR1fvJuHPacLuYrq1MGyL
RymP8La7xCWLSOeOwd0Aji/52+4J+4hTBVLpfFmngYRe8WMfTt2O0uSXeGT7sxk7
KF+6d8ljtMTacnrLlCXp+4pHmC9ruiFx9cAu2R6b5VYnDNMlZTwKu0/wuQ2xpox/
SsZ0JA3Wz5wKTZi/XVp6An4UpKYiq2zIxFPcizRUuACH3yZaJ9wIOSRd5n1dCGtJ
ef1bML/GEn6Y4TM29TfqdcxVcDqpuJ6elu+VxE1a9zWAPCs6iBheMSdDE0GlMy/A
GomCRJFx8soeEJ+WDH/GTZ6wgrz81/4bEih4igmte/Gs7RfppoUaSbh3hlYraEJP
kVpkvAe3MGSGoIsNJFXLg0a50S0wKpq1iPg04nsWP5DiG1xbSr7lOWgQ/eX2kuPo
Zk2EKnPlZb6pqZF1Koqlv92lArLkAF5wpcrBrUOMA16ug+CWeBLAFCBJAYXVKwKQ
4OWLNjVbuS4NTgOPKDw3CW22DQ6RrU32Zj/1aMSghOv9HyOmSclxpSFZIErcLlAP
IAltOAKgPwGYmBjl5nVef4JzDFuDTlHlurSmmYb2qlJFsyNA5T7vYSzvtHc/k9dS
wKmrIiPVHkguGUSKZiKlkYN7BekRVh/go6BvLAurngXdvaMsmKlKwFIv0S0UKexP
wZw/UbEWbIwDd66DAdK1lXs0ekAqbqPLGOcJrWA+Ybp9r+u1JkfG0PWkXG314toN
iH/CPn23tnXku6n9ieIT/OycXggTqDlu65Q/rOE5RaGGmZFrNtipHIitX+cf6ArW
+6mpLFyPh1pVcwe3bQTyF8ANNvQDECrBmjJZHvOAEuUXk2y6hxyHZhxE+8jLPEXg
PEibiH5iFOAYvN6+QzJeK5bAh1CqMrSCGMxLpUqdYb3fIzr8bj224+vv0WzUtHyS
AWKDGVXd+SWeAp8vmgT2dJU+1nxUswqSkDDHwtWG/48Je7n+jP7MAsC0fcWknnTq
atxIJxwnLqk43GS8yG7ifA==
`protect END_PROTECTED
