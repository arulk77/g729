`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD0gw8/QNlhSAVyTvMzuV5wflr6qJmYuApIWseYpVAGe
+CKxJRDZOBdjLKhBfnr+qbpb1Woy6+Lz/PE3HJGlbkv1LFnLPHVCwRtbBqUkZF31
9rjqUJXs3VCje3MfhAlauo1Rc73pR8a3EMH1z144DE0lYUUNrZwPPAhBIXutsIlT
YGuxQ/Ur6mzln6hUlalAZJHfB9ya3UgNRul9XCqnWxEa5twWCvcxnoJ2UcInMPWM
NDOst7D+ntAgKSR8ZhdfZPUafLw3OkkAqcBXD32KNIBkYkTT/7hlypI+OnH43m/r
OxGyXumVR/slqc1jyWafYvH6/hw3I8MNITrwPErjJPXJMtW/LxmXnoNB4SVxQHYj
BeathD6qcdQ+qO+TeUXerub6oRU86mndtRymSsCwRRhSoBv08X8dULJvMsoOAByS
fkGhFb+zcBc01x0Ibcq36p+2IXpv7rSzW86UmdCidhZru5pYLEaHoqVX1vctJtSJ
RqOBb0zYNQrv8HSRghVgZr+Ifakg790zMRdw8OwsypbNDsfyZdcyLX5JSsPbT7Ny
PVrQIFkEhqk0aOuNzaUmslXCf+s9fEabhSOqllKhFDqtmaEtnF69LlV0bLKBpRa+
`protect END_PROTECTED
