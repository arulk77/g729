`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
/DSTI03MToncvH0tGs5VSWvat3IMHz2zZ6J5SxanjUTUg4KJUXWTNELpl5AVCVSH
UDKlx04Rgbcqq70NMv7b2Ev+5Gw6ZMBUUC7ScaleUeGpb7W/Jp8GdFtTTn8HPLmO
M7MTZlEC54ZlhUicNx1WG5SV5ZZTaAWAHim2JPVGACqiGIWdyNGf7Q01ejT6gzbr
5Tc1ZGQrscn15apR2t2Z91uXRGOYMti6zF/kn7eQrIT4EOu24xzYSvFOKNXBxIJ8
S7nC/b7jrPGJt/WpRfd8K7b64aQH0JSC84kE1VfL9HHO2coijEfvauTz94nkstFs
40/kpi+nGZxyUACNPtzd1DOFd1OCBqYwm4jITdLg9gsz2O/e3J45zpkW+B1br9ld
vkph9buXeg6B9OQwevDoHdSc8ojbYbAK5aHtliniLuA=
`protect END_PROTECTED
