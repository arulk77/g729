`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Q6BLBpDsffMcVzIgNeYEPAyLH4KxdOnddscM+eZbWXyxP1d6ge1p3IXNg/8IhtlF
ammwIk7gplt03im97yjOceQ6efD1/ZDYZKrvxczVvY/HAFopX+soSPkZohU7QoWl
sko3kSkLOhtwipM9sFD02CFmGlmdEiMvaoY2jBLoAqg=
`protect END_PROTECTED
