`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL+3EzogHt6ZM0+WL6hGXTQAKWXOACmesD1jQP6NEomz
sMuj36fki9uqroCMMFYMJdza2yfj0sgVjRKG/p95LEuVdh8qLk+XCEwF+UQJvmI4
Hu17KAgIXIGUjKtOmfM7galT+UkeUtXZcGazcIfVB/ePPriuhKzNw2mwdYV6LA4y
Ngvi/VYppcuNdcI3cAfC8ayQwxWomUNgRjyjeJx53201asrCLXFZei0uPmbuphFm
bpPhhmdUVwpBLuQbCJlbNxIfEgN69JAynLWIvGFsRcNx0MPtMyXKAA3mOkMRSNE5
J0L1rkQJ35LCiqsFTJZVhTptSH8WCCV5CtnzyIbj/cB2giUmW+UwDn0OIglgdBZ9
V8AMh5e5A+aDOP/qXAn2kA==
`protect END_PROTECTED
