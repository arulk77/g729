`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wxCdATddDZP4IpX0QeqHRVKdXnz/00IgFGhmPEtqNYw
DIUrI7HPeX0VgXfAeY9n5xqvW/XaSQbzuTEq6TEBRCZ4ZuMAODCnyFM/Dh6mL26t
CNw7nWBBl8sV1itpGi8evIQ0cpV7kuPHrsSKtE/d2jYftMnIHT0lEm9QJtN59z1U
GW7nNPt8e6Q90goNBoJomk6JtO8qAJtEYvyrx93YuKjDgme8PFiQiVbvvtnaFSZS
cL15ElIKANOZI+udmVH1RCwXruH0eYoc42p+LDD/8W/Raw8GF0OBZJXzaAdcEoQ5
PEYyz46HOBUhZnptROKHOw==
`protect END_PROTECTED
