`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN0IIHASSNb1S7DebWqmxSh5eNtvT/jFuF0idPCPwlkA
85UEpN8QJOD92PNP+iJ8kKpGUYWeUx48/63sxSiBD6FW8GX71cP8cK9I7ZxIi+tF
xt31bUeaE5Q5FBYjNf4lFAYkHoMchflsuneTDpeMHs5kIS0bq12l4P0TaZYGzow6
j/0TayLpGSEWU4uhx10log==
`protect END_PROTECTED
