`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ab3t38y2wf5+qsH/48ktMKcyrM5QHZqIuDSb9XzhKccfBe9rLi33Rec2TvquWL1d
cD+/B6iVDp7oUjwhS6HGdQscC7hovApMrmzowCQKhogAJaQssYQWktDycOsBVYB3
EaSyZFk7AGTeMgBVbnsKcg==
`protect END_PROTECTED
