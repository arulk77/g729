`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDEUtZ2XD/EW4whv3Z8As/fW8LEPa4Q4KlzX26cN8S7o
B/UENKH+VmnqNmSoxMrtL6IMoTO5rwPO6mTr/USC/n7agvQJaSgjT/0fBHuO2emH
xZ9tofXFFmftQ+MZwMy+B3W+Mz9DrTkKN/G7+ZILZxAFfn6TBknK6YTyuVEkEoxh
9YePPgFowocBiDpn0e+3szYYxZ0mCnf/4VhsnvLjk54OK+Q9AhtveiTU+GR2mvTq
fzoemXs25LxCfIhjF1eQH7/ciMQ8/Kbw3aR7iOPHFQCkvcJOukEWwTmgSSllvysA
YbQIXNnRdR6FXmX6lMeBT5+Sxv+trcUsmJatP0S4qvdtXZWPKWOivYV9YTe5RsvC
OoesyIRYHUO63oaqG/FOww==
`protect END_PROTECTED
