`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJTq0OvbuJMH0ybm6gW0PdQ4PPZSvbBNI09AYwKZgjrm
t9t9ZKUifS6i8e09HV9sSOQ9FUHhCG9Dzt4rPNlZPrEXLSdXJ+rkrOl2ByBCgGrR
Amzv0HTtSlJP7TPXDHeVTIoAjopi1t9gnUv3VE8/smks/RJfHfzRkWHi1G6rSty0
TTxvfKuMFh+Fwz7zEkJ+KN9i5hw1i3hR16TvycDqFR9Ie4WxwTzTmWamYB/VqxCs
/+blCZjzBxjfLV/wLEtfjPqv52fyWLNQunH2MrJeP2pmloHuXQRDmMnW5phrBgMx
JWLbOM6c4vCjhZMmsExqD+SjTPz0PK5805ZvRcxB1cc6vZWnRbkvQBoUz1Vu0wqa
UINyq7j3ReAHqXUvSL68LfrOEeW8nYRehTbkT5Y4kNXiR2W+wkSFy8gGrZtVDNe9
xAl90kBUfHDU+kXokMI4Z10nXfaBegUi6KhjnejpgfOnkpg3CQNppP2VtobhYNRK
CemkGkPNNyEFbUDOIP2J5Z5dFUg7S0JeY5IaJh7weonxVfJ1RuwpEmNCQK7B2Plz
`protect END_PROTECTED
