`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD3NHGCsc6nClCQ3n3hr+bYaCio3IzxnnO99FaPbEwzy
GWi496ogDR/hetkEB/rGxQhbysbXWCV9JzowXVIOhoGsLin1DvfGPqb5eqMnZMWq
kDeTVWLFN9+a3kgYWXMDS9f+/jC33JyHo/AjEqfDCVT/gOCHhkDn8TVojLiuQdN2
jonTxRwvCc/Dka15whj2rGCDbo/Prf1NNI/eM0qSelmFPxtm6weD3pM9tUSFrEhI
Q8EvaxcDk8ZHCid07RqYLQ==
`protect END_PROTECTED
