`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
6jWCg6VntEnKgLqqj0qvdYxIPsNt7a30aQoE1jGtAYF1DgN2xgweyPxcecD6i1kV
7LBw9Ogtq2eYh67wxyNgcZ+EUj2glPTpX5aOcFByp0d4+MN+omy6VM+QY8dIvRf4
HrDMs3lI8wD6lE1BHqytBZHrEi4viCGgNXJ8OETJpiGclHKfDACdjJF3NA8vu6hd
q3v/QF6FA2mOD35lEqK4Zkq1rpeiFEHWiNyGlFViyy+AxdQkQM5890l76BoiWgre
KblwJH32VRPiLzSurRw5RqU9Wi30dNXxAPyXtr6JV8A8KmQZ1Y/TehWARpz9j1i6
qfpncCcsCoQOfiWlV4xuIJ2r7SThYFom95tGb/SDfrIG+QLhhFwJLoGtKQ+3r2YY
C3/tTxnAMl4Cp6BN1U0A4BUWXnzHifJy4LCndqozC+srdaozxt8P26STI0eXxs/D
IrmNj8epJ8EQY2v7zv61l08aczK6xuHJVCjaEyoVLaxOVJDu2HCQ/A/8vOLkaIGN
K4vJyFMYy3l7GyY2pz1oPcl/OMTqyYdGJ7yEL5steVZM7vqMB1p4GYAsjS1PY7eq
KunjbYbWMwcCEb27II6vSryw43odhouPgxYP9EtsIWcPBEnqr2V9PLoSuRy9C48M
FxExQKzAP0tenTyuRQmzDndu00L5qzBbWUG3qCOrmvucGXhKxVJ7e+hLXLX7YIZm
it+JJ1aThqzOJrRjA3I+pSYCHOuAeOI4Bs+MTvrCph/X3ZrneTjFvbKvdlAx3Ztk
FjFJmncXjzDStfIfGB7GhEKI+QbL+As10DoNu3Q2iZUAnhMHRDEP+335mlZYVrut
h7NKTtMMLdwprbcTMQbQQxqIYDAF6FABCz/15etL0B6ar7YmOrLzBInSfa+ELuCE
lCgtS5DSpJxxRtZGAlDb5kYZYbpGfoGDj38pmMXilb2Q3v6UAA4KdnOOoIPdITCi
/5h6XMe2b0Z0BwB8lGLGbj+BbcdVSmv9d/XfbOVeePr4J363jkBvYbsAtAxgZUiF
lCkhP38lK98H1AzzW7ouAN7aNfnc0EZ0NR/0J11eeth3/rCwP+M4ZTzGOseS3ky3
/GFzU3AuU1lRVbhHft9VJbb/QACofSpILvbD2pyj38KRum9HOOCxCts4YfNelM5B
JPdV41LkK7+EkES/cA/LBS0eYZ4YuU/wy1V/udeKrEK+wZunSxvaVBTDWSnEEP8T
Caqd7N23Nn3/I2N2muqabXNNUgtYp/cSVj4FovO6x7hCMRqFeYbzMsp3JPp+el5B
P2LP9On7UQzXyaT0TYIGyT37OsWwnj4MrB8a6U+Rnkvwoo08YebkTRcXoSxFG8nt
evPYej1kDgIZWxPMjIviTl/qIMTgTY0L9by5bv6uzt7h10sMrvvGLB4qcQNwDI/+
Tg9u8OqKy3jJuxpqpuRTarhJ38PkvSQUcFTXSgARWi9UfqGdHjfckVGU3yFXMXLX
ozI2DVjg1x7G1McZdyByoBiC+2o00H62JfnfzfLWXSYdEyhfWYrtQNd1VTUEgxhe
Umi6aaCVPZYDhf2z6Bp4kBor3eIFbdoFTWnichdZioRXwK8Kega7PHdY3Lh4Ztx6
aj7cMxsvL6Hp5Q83LefVtPdn7dIr6FZikZ9Zb5YQBLFnogWVMg26SKUCJx16HIgC
4LaL3a3dejQjadxBn7sjuJ+9Yne8p2yXN3vWCXwGe9u1+3OHKuJVQdffq+S951ex
2ShRIp3EgyXn6/K3eIs1p7WORZ/rZGfFfdcuyGEOgUjEEEu19tc24O1e8hcOKpEu
/3KHJB2hw9fDiLmxtdSlQI33H9tGcyQTU9Zsd5PkBj/q22Mlp3ci5sA3Cp54d2H9
lwWZATFbrS81UQiObeGuuYrk5kEYxM0V4UJDWylAasfoMnNuYuT5Hzbp0l4bm1xM
dueWCR99c4RUS1xxv7RZ7nhB13l48+GUqLVRVoZd+XeoKd2zUjrRHpT83Xbgz4f4
6ls3FucdVWVJTJCKy0n2Ml3rlmCL43kwcTmok9ZDQEa331JXhLFmjQv52QKFadg8
zk4ogSvCNLclZo6IyRBwnFzKSewhemiD1rtZUbU4rSZYZBodqGWafk8B5F8koLys
Exu/4jsMplIqxPLJcPW60iSI7Dk6jREECJXWpc52Ue0wx8h7nVnG0ipSmftrX7vx
nmMhOmRQnjXNKmmPk0hNvs+sY9Hy2YYboHvwUHwNEebBUT25RUOUBaSEBdN71B4S
fjC/vTFMHGTAzBx/5dCSNFia9t4pjlZShXapv9d8CvHLXdOoTef+xKJbPkKeC5uO
2gSYhE9WZh/lQFzCX9pvjB5bJ76ZNB4FJrAh0XXtJZpjcI7hS6YLvGfxm3++eVU5
Jnj6W1DKpV66wHxcbrOQOlmD5ENKLkXxtbG8XZHOXpQvLIYd8lKWp9VlGJw8n2Pj
U0Zo3p3Z3CbnY+lYIEzTOxZWO7OI4+kidsc4fk5cT7Qw61OdShgl7NizRcO7JE7y
Pko1iBRljZD8GJc24sLR9xyb3g4QOCS4CPGSA5yCIrm/XDaji+MMDX1QUIoFAMEj
liWtWhARLWSeBA4Cu+pSuVKZ/v4CHC1kqvTJDkHeYn9RkmsT53jQEkA4I9V1e4li
2jSEquRGcsd9CVp8r7dGosh54TTMbTGzW7SeeMtssN+uxdToW/PmaImsacBrgFVC
bwkuw0A6OCUPTuVqbr/dv8cExHoJ5DO1SRP+U5o1Hyn5kZ7BCj2oSrjayOz9pDwq
D1AEU4V8VT4yAWuFGYnA5lay8gc3uPNak5b9riE2s24=
`protect END_PROTECTED
