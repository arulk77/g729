`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C8Kc9Kj03WDXiJbRcBR+xf5FR9nk5RqW4QGvLReYc+m8
esR/3WImQ9gYjCnLKt+FRIzWFNsvzCZXtAALQDyjniM2uvtA7P7K6jdVu/q730N3
4mIkOC0WYxq/xRKOcJMvKHu0LU9wn08rkY4iD4YCfPzfVIjdqeIdeFG4e2mn9Vob
BHvPIaoGvzX1f9E892U453WdByLmHydfb9kCOZamVz1omib3TgFeqtiFzc3CBTet
2ojksL1D7NDV01bTMy6bEEUqApbRgkpAo22wCLzHs8Ruw/Xd2/0KErSBTmasflBM
mWa7Jkdp8ykLdzUx9olABke4N2M0z3uvvdi/yS6SYhpeAEf42Pr/O+5sjspOnaU5
0JssNoHQUIjyfOnsfC8G5mC1PEWFqXznydF35Rwp184+JVDLIKYtBGxmh0TRgYwv
fG1LoZ45AVpWp+AoogxyIA8tdiSCvYtIN3+b68JbU8TbynO5KgzlHMkhqxrkI3zZ
BdtHE8rntv8W8ua4egZIddabbK9Jk2BzPOvkdXBL725JkWbgkOScN4Ves8NE0UZ2
Q92FuTidBu2sSrjSVC3Xo39Iaq4L5S5VRNy4Z/3YLFwYCzMrvVZrncPg0nmm4cnz
N6yy2ed02+kZPmBXZBkyOOrewx06F3xq9w0v7WhparvXNb6N/unVnZilARkScXJ7
VAoaADjwkdauwlcFp7uvkN48JkEorPBM7+1PHBKHslyiq1H3/EVnHuiKZejfefbU
PRY+f577jCy5CxJozfMdFrW6y4mcXraNL2jChUAmLRre9BqeEe70AhUb0fdl9UJ7
ZAdeL7G01TvHX3VmcLVYwDa4lYNh+5yO8olv+XH31kVa6yNODqOKeDPERd+C+gH+
twm1XuYZLHtpZ8oJgRey/Dwd/OQ7QI1HKY8fRWMD/zZvc5v6D1tzQKQW5mxKsyGl
cFrEXLJDEpbSo5/wK8Mc7MdlL3rj7T3tJqbtdzoGtTLUSyctzQUGpkLyhsnqNZ6n
i6RqvAt9wpu+lZ2bAb2f3uPBYy9dvcwzSl5aG+pAGev/hfhUvVo+nhg+jp1LkJu9
L+k2DZ9fREwgoBAryAjSVxhaqBRHtVQgXEEssNn6CmU19mUfob+TWJiKXBp0dw6w
3XZPAvFBFqID1lvLmU9/IJxlFu7oxAjJnw4jfWxsUCc=
`protect END_PROTECTED
