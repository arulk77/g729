`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73CxL2eBvXYuNQ/3AcaIwu2m3EuCHMFGyHKVbwob5wTuT9
sZ7Yfu+kYoC/N6ynUOk281OBAdpjIzrsG3gO9FRrTL30M104gUOpcvDy0z1g395v
RxaFeQQY2quD0e5uoWc8oKRoA1OAwF1MDNAxZ7aCSJBu6k1HAumfCSBLnXJHyX48
sxzq4rKqlPXiCo+obHg9J9JDVLSLBMMdxunpzykaSi4zdOPtBDgmV8KO3v+XoFuH
yRTQvqthEx68vpUKeHtCIz9+MAkxmrGelJiqb19iqLP89lzIcoe8OafNdFgBLvM6
WH9dCBq71HhpqSBtVbEhhsxmYWHIjxd1jJfcH1sNFpLe8TfqBEOD3I0meyiCRa6p
J/c8V/0mHuD6niJ/VxolAqkEaHjIolKvw6e0vchrGXMvc5z7Ywhv6iwV9mrDNL7O
zkgQVGaYm8WxrL3+P1xUoE95182V1pqlmSTx9qRTde7WtzBWH5SnNLCN9m2vYo4k
u2acD71BsRPTASGttdqshHHGssyrRgxTrv1xFS0ctPzU851xGlnJO1ac6PsRnSn4
hLCP+4D9JcfNa5rKjysfRYRWh7LlMptHuSwVkr6esjuuJoeC9dJEK1T0zjXa6r2y
tXCQ4p48nbk5lxA8jEWlGcf8s2nwUoU1rj3AdLfn4O9Qi1ePxez09oZeYsyY+4kx
po+wQl/5gEJnIBIzQ+yfpF0CAJVCagmBVKZh5ApAkSrhMu8mIEEYtvCSossOldR5
`protect END_PROTECTED
