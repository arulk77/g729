`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
1WfGesVWTsTPbZYS1TmQ3OnoizrNkC/Ek5a9Sn85yE/gpcR5lX/i+K6bZXdZvn12
0o6vFawOv43P7lqF8hxBqYxTbjWLRdJG3MnVJ9NJiCbyg2UB9BdE1MznGzm9Qynj
XNyp0YYjrZnr756qcjyOg8LNGjrV1pEn72dMwLhvn+rGITP68/hQc//2dlgazpN+
7DxJKDGtl+A1HJzNE/wZ9NZASGgn3CwMKUlE3ZRf63eOw/o6598mA1kTZASRvQzo
olIj//hJqeO0Y5XxKiP5t2x2vkvJZ1ZajLjpZrakloQ=
`protect END_PROTECTED
