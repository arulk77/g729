`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCRI3tJX/9zUuqL/mNQBDhrXlAv1w8JoG7RkSzf+6Ais
Hh1RM2ZpSIryteIWqdz9ejO9PByhu5XzX7GzfpWWqhXJsvXAQrlKOtn1mpWlP6VL
C5f9p68fWM8MjCKvP7W/zIhnJipG2rOBGIVsrqLlMlodYvfYE0npa7xjH1JlqlRG
`protect END_PROTECTED
