`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
F3vXwhZCiUNUuC7MoAlaVHnAjyUb/oNtv/UDQ2sLHlSTVqiaZeCLTUdIOrqgXj0V
qwJjG++F0vIQvYQnJuKXACRxScIy4XLOz5sJvr9lHjRERgM9Nj5gdm9xPvhel5DV
dAFKyKWAjIunm+o6aohEBdigO6D9ZeLY0pOBUnbvNEQhBcdMkcUACXLyF43sncs7
Yk4xt7+1AnRqCm7nUbPi/dGqxXSZOB5Qj2CEwTCjY/0VhCWa/6d9hQVe+ont99uh
onkva4soNRNAYu1pq8DAuJunvH3/TcvgW6+adxhttEY=
`protect END_PROTECTED
