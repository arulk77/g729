`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xMz+Z+/Dq5GBkwijZZ3WElyRvyZ1fbGsaB+7Fa9jHuw
fZdAxav4wtKvBR15TGteerlkt0BdtnG3s87JDijqabQ1RdMXuHUldTiQ1YXrDUzo
nxI2rQlcBVgaNIuAKhpUt4vDT5jJa5BtBJHFirzhVdifeygzSBE97nDcLOKitHM9
J/mBtFnMTp82zQbjG28bqMsdfSewgu5LQgxaU+nRURHRzbhourycBiGxBvPFO//b
iXQL7Dz3RcJhuwglc5hchU8HkSHu/buvjKPD5ka/21o=
`protect END_PROTECTED
