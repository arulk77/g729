`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLoAIcsaDK2I3biH7bPGy+Z+evc+MR4kEzQmE9vRHCOX
nvv1m9nDnCLy2uEHb5IXHa2Bg/M+bzGQW4tXc5yGUwjdJYtgsp1qn8CKOKW/Yo+k
ruZvhUlKBEEmLqkiJo2LxqUeLpS0brxNK7PDROqIl+Lcogei7AhtFtH9X081zuOP
2j8bZfh2itQiyNXdWgBdsOmqhwdLQuvY9AOLvr/dP8dTmahRusXVCUyTi719XBaB
Fp/8YeHH/BZWAExDXjMX0/KAhgE+hdizDtPgtlwAYD8L7e8q6eDNLKd8wyjRO8Sd
QcEIZPot+My1tHO/T/IpGRLqqhHWPE1RDm4eWgCw1eSmV3dUFo8yJUJrKq9vcjdP
`protect END_PROTECTED
