`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHEYK3A8dphQtX4rdkBSHDCFOxD0/Zz5dXn+Up7oxn3c
c7UY41jgPBGk/5utVC+0Nr6vugwM3STTEL6703s6Bggg/Fmee0GWg+UuJNcMrfyS
6kSrvth1hw4ElsNUAMXziOY62Gdp4T8IiRLCMvZWczlPsH98wmyVT1sZtkZq9mBw
IMsBPGOZ3tU77oJv2hrz73RtHRZTw1EZa3MY2I54uFzSJjtXkRHIZDqfa6v94ACi
yb2hfQPqA7YQ0leouSSRZ9RVlBzQRRYAeszdBjsMpXhe4uLOlQ4g9ZHw326JANR3
V7BXVkAcpZ+j/UfV3IRIDd+0v9s4o8B5Y2h3TLmZUOXN0is6KabiiRltePxbz2sc
Xp8PRfBIi91GFr3qcKiAmQ==
`protect END_PROTECTED
