`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIn1sPBWj3dCnOLP1dpJpbT8QYsIkW5Ue0TvJtYNnbfD
v9nQ2L6Mj3PB/Oi+uAvwvqr/E5vWFPwKfXlXw2mypxXuyE124TsMXT49n+WPK7C1
C1KRrmjij5ep1EKwmw2EG/R83jmYNZjq5mL81TzzPHOf5Zn9LAlOOqvDJptMqpTU
a6mFiUaICPHg/ITGhIRQxwquNZTD4l1dKmsKC5cz3ptcc7uGS77upae/G7cOMsfl
0iRxVEn7hmymq7kc9hJBKYnaP3PFIqqEzRbRHcHxGbkH8l9/XyvyYEuUSFKuSBUR
NDcGmNY/bcwrzVDBRJfauVje37BQ2eMjZ4iuTJuzjccrvB2XEQMfTYELcx8SQ0Ho
QqiiTl3RDGO5OYR59yj8Fos/IvhSVduedqtoJU4FIk6b6t+ZAfLN4PV1g4EXcSuO
7FAshO9+zt/6jE+a0YSAS7wUFn+Vh3MWlbmfh3KU9qRdL/pPzKNuvqo50ZYZ596U
YyejNTubbyua6+TXcFpPH0W/3UB++1SWgcr8hMor8nBXqWhnEnuOHiAaalOQFvl6
Vo+nL7AKnfKYhgilj0jE0NsJ/zh5zdz8TiLJxeVU/Dyhrdg2hLwhjgAgKgRWqdAB
`protect END_PROTECTED
