`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
O1f6jYjJpj7Ppam/hfymDDyntkA6gXJs2SNPC8hlw/zxm8ozbk6UQ/lRfjl4mKM2
LKEFC2TdTwEREbd8/i/PFp49X7C5ElQRNWnbn9fPayNXD8RWwvJxTazAAOiymRTD
KZ2xMgDD5wfNfYS1SNiiZP7OEreuPvc/mUYMKWleJ79YAD9qwCbR6WFSv/bMo8VH
ML5CKWlechar+A2H+Z61W+g/yPcTkVYuZ+3uh2RBPALRB26AfkBOC24AE7Lzhr3a
Q8RlkeoboE7waCGpTbpWxwkwsH8F0GVsY+CYo4JizIZM+qBztTnEea3lZIn3oghg
2cXaJfdFyof6Rqc3YbMynrgUfKPvLDS9O4jM2WEDQds=
`protect END_PROTECTED
