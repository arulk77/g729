`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIekSBl+K48MqxIYvKVJd2m2uf2qLCyt6lg78CtfXWWg
3tOaQtELg4dIQW1CxXw1NoDVb9LQNWnYrnNnoG/NH8YsoOyKi2O8hFXx2eVEaia5
jNtTq2NaIqsQAC3u9XXGtaubKvhS6LdA3fGM8QYiRGAPs6U60CD0v6/p1SfcwxEB
HyknipdP9/1DJ4v2hsrtfwc0eOg3w9AWtT3KA7vcrPyovwTU/m+2SkSuuNLU24lW
5DgTk0bEh4rkvtiUW+mzkMjNxIyJLDeecZazctYIB4DW0P0IHsS3QuczmyEkQZnr
YIGK6d4axt5wJCZrXSNaAWkrTfeb2gFCBACF93I+uLxZXS5JvrSP/MD9tbe9qaZp
/x1oCZwLIRiVMdlTpj38ke11tjNJURpGnp+eA3iYj0dpjObwLGGSqCZUJ0awc9S2
eiw/ktiI+PfPj1jBSwrYUJ96tz3xxwRng5f7s03r1j+rBIdbD+iT+QyLIqnQLu/Y
V6BZtq660R1YyhtFUBTSDSjNXjSQMmb/jnz+ZWr8LkYEDFS5XuTFH09hBT52RGQr
VYvHoVZKESD0pWXDMRDTumlSmd7/CG/s3UroknZ5AYfsda+shJTt8ig8tabtwmGM
2H2zeR8Hyah9e0O3xYxF8tyjJAlH03CwlS0MOEdeh9Jf4Q+2ihjwUtH0eYvBjIHA
8Nk/DSTT8MHngWvYoDG9kgrsEAVi3PnDSipv1i4z57MyqNkCm/ouJhidU+V5n6Vz
EsySV+q13mShbquVhcaKkC7NfWnpu0YQUu7jbeJz/5btQN5D3LgnS8lAD3csRTyM
OLh+E7Zz/vU06U2MXfMYk0+5noiLeT4AsSWmjkQKDeU=
`protect END_PROTECTED
