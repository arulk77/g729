`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mgyH0ssoIxlogg9LhVIcwZuO8HPpXpST1G49JNnFLCAqsdC7QKEdpwMwbFLx4WqW
1rcRPp4Ol2mjBHQzla6mGPrEfoHZ1xo5ppEK5dv+ReTlE3vSJ6Z0aPl2rpRFZDWk
wBagLDag8tl3hWczOeg96CJGW7x625B7aWxoT8ZpfGlolJfOEG/wviOM09Chw4au
o9POy6EqKQvoi2pJvvi+0AGu7iVWex5Jg6kLf89aJo7Qm7Dm4FqhssoyZVdeaIk7
65UYy5Uk2M4IeVFCkyFSi3XNv1GCTRrMiWQUT9PU918=
`protect END_PROTECTED
