`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePCRTunVcLMZyzOwcCvTAzQy3sfwqUCQnVtq5N5cAQ62
q/EPLH8a5Tb7rskJORTTRlCy+VlZHxsYcqcgfASSXp/ypo+O806hQfIoEO4kG8ak
7gaxaHGqLDy2+3KzqtDz83eBSvWdrpc17Vz9J2PX2JSrz+6vThVgMp6Cj235Jpe3
sRz+L4WOLq1dNy26QOXPSfMA1/bsfJoJTzPp27LZQrHLOqJiLzDW+R/wjORpVNN9
/So3W4W2GNemVdy6lfkSy7FmgZghH/4h6b8b8WsNob6pOfRIWAsqqEqzxL/BNpXr
0gAkOrYcSAKehVnUbyjNC1KEEXXP67gh0TbJNwcHxqTmTCcDX/ZJuKmdBv/rsvOu
LkgbO/kBv+sZOC/Tl+bxDi0vNgGaqmnwiNE8N7gdiAXdy6zmapJBefdwLXt1L8aG
orXW0tYsPLjfGbINn/W0MzibXaMzYZOxehnEhcRg8ROXZRugW6D3IsUaZsTJ+b+l
12Y5TwsIXP5cmaocxg0UlntEkVzlSp+mkVfecz3GawCwrp96BPaRm35kLyKpCusH
mR9rw6vu4UkTXitCYzWfQoV+44RLWAQD23Bqud1IG8p1uqN2aNx/1Qa3pudue+BW
0Dh1jdIz+eHPY7C0GvPsqkzM64TK6d0hyDMgbW/44UqZh3BZHjYc3v8fhFzAvx/t
l9UzyF/uVrcvSNigOMo1ypNd07LRqZdeK2lpFzjKyrVW32e1MxhsS2JLNy2VyuWR
MkLEFSWVGa+RJxZa1BcOaDTzRRYi+BdMnz0wUO4dmu//wxD80ReYNy52ksZG5wG8
e47MoUh4DW9VZG+HztitGbw/A3+rzwNFlFLL35srPxk=
`protect END_PROTECTED
