`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4y7pn6CKnBCmRmaTkoGvWHVQpkC9YQawPCDyyvFDnpht
3Hhr/Qk21TQ1UesSiYaMTTUrG4VrGbb3QON2Z9XdyMT3e97LJ6APsPCgX2PWtHxI
bgs1Xee9CT2tr0O7MD87aJpIaN5syxju7VBsgBqB//hoHGxFbcmaseb+yiYHqdkE
c0k6JH/JeTPVAVhl8tltZn6bG0ytYdfILDhZIYxVfr/pVJS3LC7Mql5A0Hllnv7r
OKe1Rl+H2127rzsoComkYRBUEZw8aZmIee4uknzGGQNpTe80Kz7y9HvbcRhMaLtC
+yZRxhCIQ4US/uiiy7+fsUSvyeaLpPzOwzMjlIyNtF2TmuKh0NnadtcBByxNu6Sk
4vl7ALJnnW0OTWIAAv/g7qEX3CjTmFOMgDy9IfkgO9n80nkdc4qA8hPnjd5QNH3z
Vi+KAIS3gK0Yrxzr0xsqUG5nnYLhzrYIjXswdvnF604fN9o9YWvVk/KhZTsVAzOl
jSWaBa4lopMx/U4m7dvFSUzoEBYMr6EfQoJrwd2yUIUiE/AWV5mB83jwI6E2Gnwr
hnhBNlEo67WrFPUnjW1clx+A+HPpMXoUIWG4Q4TFPDaL3kk6O3CLfGJqDFJ9N/3z
`protect END_PROTECTED
