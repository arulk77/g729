`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
FZbNXoYyCRzD9PdiPwUA4j5QVwgSsFN+f8fQRFt/CE+YVsQp+mN4LzwSU3LMBpyp
TwTFx52g8ZfpgCoHmUnad3vcSxEBSeOPk01qNzs4yiw3CQQqITYM68hRQBJajkGE
bnpXtisFzfae6Pz4Sxf7wA==
`protect END_PROTECTED
