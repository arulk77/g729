`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Xx76gbuFUV5OKBBJ5cvnFndZSrxyko45W9pa1/eS0zIhZpJw4CwPN93Fkuvzr7dA
4FPeM+2vbTPU4z1u3qYhngde8Qt0iEqBuvGe5MMxPRXHq7WnBpB2wuaG9gQw2nRS
Dep48ZU4X5OMA3HeHpUuKA7fQ7dikjg1RSvAB41ix8+Z8Idc7wffqS3kNNlgNkop
`protect END_PROTECTED
