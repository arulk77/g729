`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C7z5xo7Nrux0VtqJDtYGWWTvpTAeUukoDDBRiJ+vBJJ0
eohT6KHYVLggsIBCdsIgxYbFKFIdRUZF+0npXTVsAoCFThP9hTxDWByqxEofQHXM
dxksDqH9WuouYWEBvUl0NqQx6qj92kW8qBACGxeWBEQ+cO6a6fldlxuM7z4jpByq
TAHfRnoSpiS+VQolkI1tW0WJ9Y1UVhHrdlUgSocCE00vOWaUqvQIAhaC+sP1bIVt
UQIku1uQMqZXp8Z0tec9icKQeMt36yHNKqkCmboQv06UzPg7XMg0q0uWKUTK3Ty+
oZD6hwFQRaTyigcCNykeyWVWQyLWsYavRzX+wMbW+BV9DodlOgMVM/SDQuL9fZ6y
6Ck1yYB1iJIpCX5g0wtLMzgmdM74MFx+AU/3AXHj8Ex+8CTJzMsmnRqWKO2AP2Kt
BC0jJdX2yrUoDBca7MY2AQg+TbYwJ0nqPhOYbYvOu+bwYq5m8ZOvM45ltNxwVLiH
`protect END_PROTECTED
