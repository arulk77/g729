`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
57nOEIljdjtQFfXnqnz8tvb3tooe5E7PsSGlyDpRpUTC4bCD0eTpxiDFq9FJiM7j
53UK33f3nmhfgB0avga67B1VQPjddlqzDtI0BCLzaPTndlL5kkz/pGsC2hEfPIi0
NB8xHXYQr4cRwM14ZVfYmYehP6CjoLbSI7kqIbpLfshYV5a6mCOGuCvSFanQUcSn
EYjILJZ3w6ryv3qwZphCyNY9C03pxeT4c3IcFI0TNiYGZoBcC426mkWn5ixoqmGi
cmFpke9fAUZ7EwS5J7vekndhkv7PWaffYjjdDlovG8O4FXYrMbhSNJR/8ZQ0pLhF
3rsgsfGtaBHjJLCleTngjqhutdoD2i98LaxkUTcTpId1uGoeh5mAGp5yrrKKtW0m
4X8GhrvNBtZYMeRc13oLlsiK8Bp3ptuVZZecygTXZco=
`protect END_PROTECTED
