`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
fEc6S/JlCAxWuJ4Yp+0b19dizwI/q+oE2KuBxRfZN1fKKdytsYx5BPAqZQqTzi4t
Lv05D2pcIYDGhOQtkYGd6DS14GPbhuQj7xlWyMiOLCBA7Vj4nTp0tsU4OXjMtQ8h
G7OXmrq/7FEhyGLK0epGVhFIwu/XBhXTEEEwCfgb9WiqE5Qi3H/kDJ9adrHI84ES
ET15tswQHUi0Lsh9XXeILWcCzG5zRYJ2c6A4ixWqPzZLMbn81itZlZKO+VlMndpX
crQ2WrNUTHmxlpvA2O1S6ukjMvm1sox5tkODkzpXySqgs+/uC2GOuJiZ78V6MUZv
YXBZvUyxi5lZbePkgMp/2ibDAoWL2OjuO6tRzuDd27+y3WJdy/vJyWp0y+3Yn3Lr
b5sRFohyEmCMJQHe7EqYG6U909UaO3Xyn64sCnGctYrDaNL41YYvnWpSpfbAUC3j
SN6Uu1rl9YNFQDuw0yX/cfiZhQGVomzUYmp2nQ+CkM1mxtA0XJKnd1deS8oyPYEH
Q85jGqCJcvGd/EavmKH4DLGbIinSwDAav/K4r1FSdCUt3wjVCnkw/HaLq3vvdKkD
5NVwrUv321jtufxvEHOk94QsRvOgnTO38rSlU/1b7QtNOHwok5exyY5EiuKUJEU0
j5zzCw67WwRw79tRT03MP/4jbSlUJwxAIC7edEjLej4rsE1LreTREXJ3VhD9OwEr
Fedn0bfXBIRAMVy4OxjXfNtPaUP7hGJ2iYthrTkGmHL0kfih5dljyDR45MxQ+oDa
3JEvQ9wDGv9Ypbu+F5RleRw7Stk6iU1iMIF67Q4idpl7hBl562EhXDwyB+v7xiCe
IelpOFZHr3NiwzljcJWvEYq0GuxJIHKRsxg2lGLmYelJmPRoxKTChf6XXWS0U9RZ
QtIYY6sbGUBorEJ5L6I6PkyiFRRXV57HkSaEF+a9gBFZCc1BDJWF17FfLbKdhL7U
FXLqisJ7u1XDwHL/9J0GOxCycxw/hDJaQSrR1D2oXPVN/9Cu3uZGia3ZfIK3IuYG
S1MORHdReDeSYKFfCI5FYjI0JGfN1YSlyUMe/H2yAeM7Wte9ghBvZjbJE8vUeWWG
ZfEPJX1sTFRh1Suei7QWUPf4ZPkAwTEsFxNOk6s2nYOzYEIhsp+d1jk+UhpVCtCl
izpmqyPZ5qbHQt4T9si/sWF5pHgOgCBRHmlt0gdcwe7xFTrSuEzNhT1DjR0WJmhT
Rurpzx2yzGkq5jhhuC4JQGCDiHKagQL08bgm3e7583zK/9YW472N5N5uoBECQp+B
i8SmBgbRBQayMb2uAXOgcQ==
`protect END_PROTECTED
