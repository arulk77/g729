`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Z8y5/hbzgIvOouD03txJH+/pF1LB1JofXIDlKvRRO6VKCy9zmwYxhtyCp1mHB2sw
+uL0k3w0a4NRHWu3S8feM+96ALNBnZtOTv0MkZMGvklWSrgjbljCbYMNXDY0oOlA
jkTT6zuNp1zE9dopXzmx9XCm6Q9SsA7zPUzDL9iIeVLjOjjdBNGGMbvgODvLMaML
9hhWZbjWD3MuoMrLPqzcmO0jq02ffzjUQiJ0fdtXutNWrIogRlSl/bqnj5DCRHt2
rJ5e2yDAfuLO0eS3WkzqEWS390CyMLHUcxVrwK1vDr0FnojD6DCrLDuLms8NNDwz
8gzl8ikECuaQxwOrA59u/hFvkZ+Q1XZaY2M7G/w3svZPjgE3JnstWOKQSLA9/TvZ
oHlVJkkge1IYasMftzgr3Eou6bWE1n2J9epMeM8e1zQor5CNFE0bqA4IFdEdSdua
8ydnVEjOUXXnxntwlnRmtw45Xv4mQnR2AJkAzCK6HQI8+UOqNDY1BWRU/RxGb38y
xz+D0Ehp1CCmlOLwYQc2ISZ2G/jasiL5r28ncBXKmw6//kCVBbwYNEhMHZov2TF/
fciCZ+v7gmWoW/ZLDaFZxLhEFuU7uFnGUjefgDoXnAKqdLC+rdu0prFyHN61ZTRQ
x9RoCrbAJtaJwbyzMr88sXqbXvPyjvB5PBlWP5ZGtroAIYN+1VQxEeGZciOV8Esg
WNpzFGrr/XVfZrM6lN3HElc+wnosuVC5I3RqZxOzGBn/zv26CQ+gMG6eidcsSRYW
YLBw8yFUuBNaII3F59vefuCIVgFpqwpDyHRPuCc3pjl0C9yigp4U9sbSa6WxCEhW
wwURfKWbE+uL68CrIO8j42fBkPhSLn0aR8MeKF3IVpjDU+rX9qPp1FxO7Y7gr944
ozn8ux7rr7Pfraw3eBfgqzVfsosWVyVoPP/wak+dc4wQ5YD3ABAplB7d3ylc6F+8
GdegAR41HigdC2IDpeddmOJCP3QaEtOIl51DNGE1L5fOD1tkINpSNpIKqOAVjCD/
U7GrDb0HNk0jUEM6IZmTd4CKIzl01qYXIzLn+ohGjTnTGThZs0WK8en5P4ryIaUl
CmmtwZQK1lY3Mim3e4tcn8whQin7y3hQe2/TtQNraH8VuKr9hHjcIdfNyvFjmRVf
TvWcuuSTDEChZhg1rMnqrtyrD9V3qhQKauafDoQNAD0RiK0xQu1UyQI6ptNfol64
WLNDN4iPJf8qoqBFQABr7ckfIxFWf3zUMVCxcmcEaXl2IaDh0ocZYhYyv6FTWm2g
J5/3M0O48ZHXhzLl2oqPM7itfQYQpX1XPjz/sG/6gmjqdQ9/fnyGyXg9JbbHwS5p
yA2Wlamu3n6kSo+BOugjFfNOhsVnvQEaoj/vHBUNFzTYv1J7SmYPk7tPhsVCsynB
DR11PjDlakZ+731p/aCa1xEDg+btsQm7R6xwCuF66uABvm5CTf6vzYCaafm6xzDn
kBzEPOD6u/zUkCz2J4FrKkHLAOcJtZ4WTbM0/rhnyWntyasd46gyCbKs1R2145p6
12NpNZP9zxdQimDs70xlcpS8g2MZOsx7mSH4utB71Sfv3HmX2OEE70jkWgDXcF4+
5nvr+QA5DWaFRsZggEhrXdqlSY3w3/XiGEULQ0A6dHlWlDMtpBkrHdGAgDxgDO12
dWfsOA9bfl4TTdd8TQ2kyhjr1Eq51hj4IOAD73Z5/Itn9OahH7kH39lq19tNqiAn
JnqFDEqkofjqy7eV0zqWaZVs9UUVcHg2vwBwEAL/C7o0xFY4SLL+dJraYZ+Q6ZCK
5GiZvFD6WEMBVeSIVwtuxH0HjUbryDtKqPVc9srpc3P81UCqJSgw7NPGVBcJhLkP
hX4S0Fti6VZS6SfqCA8ciNdggtfDoAPaKiPxCIHVk85WHPKDQ754+Gu73NZAc8BW
ogfiATe8jEOn+1FGCRSlK7M9lyILpmNTTuxuUDzZyJd5KFS7hDhFneXy9VOjk2uT
mRdi1zUJNoieVz8wxevPt4YIrKDfILu2wSYex93+iCVy+e2H5v2ET5s3yxndHLkp
k+M4Bwtco4g4QwXkZvvO2QWKc/D5fvrlRjCnTSKHMmaK1wEZqUCGSy7qWieoOgpU
2f8GoK8habHx/7cgwre2EgsZbAER7w4dqyV5JBTC6cmSN59H9K61FTNs3f0XndOl
suixFeVlW7aPgjSs3wyxw0230t6BiAQayU6OH4nuKXqKxk8SSQtu6THqzu5Jvijr
G0ke+h0u4+8NVvj939ffh8eM9a9hJd4bWZVmCFr+mRwdWJQRfnFIqThzsrXjD1EY
Ftvt0M6Zu8Hp9nphqoK2vsQYsU4gY7pkuL3q+CzX+gtRB1HmXwQSo+uGhJIbqEOA
OZISFHyM/WsoFVYjkiEeUH8HiNSX7auforqcAw9xETJbSvR/E2jUb8V1rNYjf+jH
dLUla+obD84qO4nsjXGWG0TH+SQla7GcsE5OKO0xsWCZM4gNA2ayLx1K0gNSwVji
tTugYi/vPf6N12W4ECX6k/Q5+YYkGiv8q8X1pmgxEzIoiZ8MTgHTTNbXVxl/Gwl6
1gCRNTyF7cUU3YTbMiOjCcUwFoo6IplFk9cNGnh3C27pQpRRzhveEhuieiwuddJU
lS5uLWLP1MxCn0kASZMTSyR9MF8g3tGMkXrozB6gVM+YU4N5+S+48b8NLeQs0fIO
3fvnFUOVTx2wFII6W+ZYLJGFzdapwyqicciQhOi7jfCOer7INibyQhlQXbXYq2EZ
gRtcvz/fjwGA9Ffu+se4RBm8WkGZSQvelr0JqHgkTL2VcBESAxv8a75y0x+L8Nzx
69TwHfEYWIbA/+jmEVH/PMO7UD4CR6x3X096FxiYPEhR5uJg1FmDlI+ZNTPHSEJs
yF2MBrxkQ3aVz5m/kr4lUuP+xRvacCvOnTCHWJmjZnlXHzMsLti8BPPlrm8vFezx
IwK7qTZ1RNdfKsHOCXBN2/b9AyulB5NqBK/THegdZFyn1/Cb2nUlQyW0IfYzdHZa
l437HSUa9Nxk4YFQa9TFEkJRah1ghGwcKVVWSLL/TsTY69euE5gnB8W4Gn+FzHc5
E7pAKif7U0ZYbEtANOVWGt/qP3+AgIzjYL62FIljhRHdvNzUfUriMZOKP88PwuLj
WFO8rtjwLqNl6aAA9X52DBaYJvZ+TC8ziGPggL8IVyftaZOR8zQ0BIsVyVmeHvlH
bUlJX915HsGBpwkW6P6tXAfBjAqnx0jh2dvyQdk8dmly7FKrHF1giEBibWhdMLrR
`protect END_PROTECTED
