`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkatu/SFBg2F9ZAVNzaG0tzz38YyxSkkquGzJEf1XsMvG
4B/aNVikTmbpcXQIJJNclT4y2+QwsFmJpy3XT8Cg9m2QBjcBQtvBSLTeqfI4cq+6
q+g5z6lGKvaf4k3ohSpu/VEmRO2fXHgUMpn5b2VbVmbnHBFcHjrPEUMa4cNiJ66B
EuMXo54/ynD7rpVpFc5JsdIa/D3FZtBCuvsyXGYWYQN02G8kd6cHI2r7c+e34AF/
IPPB3QfE8lm/CW2KgUdeyL0tZxVDk1fxVCbtjeRdWUTeS8i8O6CkKAY9b+0ZQGxC
oL1G3F3+yhzAIISuUMClMwAZj9OrYgO/Q0XX5JFnUUAvw8mljAv4T8OWIGBNUHLS
EDm8JCpC0MRRddLBVY3K+jbniRS+VJA/wYw3wLZ1t7is5bssIJ9DbB8gQqCMS4L+
WrCbcCI4EMuycHErmr2UQEgxl+awyKm6ByrApnZYCiWEmRLBNMjWtfZrU3lFvpO7
lyFaYqt91JUT6gEbQFqU0Ccka5IuT/e0rG2CL7i7TwDt78QlywCDUL18ncHRgpzx
E9BiJp7exZPBM1b5hBA8vF9Uuojd3e5RVhlzLZljOrySb8CGaKgywxxD6c1RBeU6
LW6y0tXGCIt3bVqPvO1oviwaupc75V6PLhbZPlpak9h/i2nuqPViHe/MtwZUbUfh
zJAAXxb+Wx9j8lCtZ7YPv7m5H0HWaPh4a35ei7SXYI6lhLpQTMZDbr2LjRs4n86U
igpqfK+R1nyiQ3GRlLh+IQ1gTViuguBAF8jkaWM5jZFU6e7GXQ4zO1fPtO9OPSCT
ii+POUirDIyBUo5PDHnAK5lNd4AYN8TV0TuVZAn1gXrXbd4mZHACNxRgqttyfUIe
VMrf7OUq1JpH+zNGtQhVOpDidlmcHbpb/mxOV6fOw3nH5OJ2tu28II46zxK3g7Su
kBmYywfyR95Q3ccAa4ACDKriSrpS0BBidv1+COYqnvm+bzaL7MRW3Ce4EBzfHC84
OEWDVPk2s/ypxpzrrNWoeaYBDJLniSpGgHMJgS4zZwCVg1UUYrme1NrgpFZlchsT
OL3+yIlFVC3xu2CJlzoCi1UD2PbUWVszYHCqwAZ0pK3UaAjIoun2GgJyI7oMf4wF
UzVGc5taQXsFjG6OI/eNOa9kKOB/mB+EYkqGciOVd9m/Sq825D2ogMJdh3YyFsvN
LnHQxAaOpisKRF6B/snq5RwEIXiiA+yOAnWn7fHHW7S8OnoIrIhidz6ajShEyQu0
ssScsh3WkPMJaQKH4j0ptL6pMpMeOPlt/vJ+ZD9ChGeRr6pOyklxzWZKPWtK/PDK
jwMDeC6Nd2Qu9rlYZYlMbzNTQOquybPHvw7J5YvLnB1uPU6GoEF29UxgUaUxV0Jb
fPuYs/1LBd4mTojRY4Zgcwtnu4jC4UcNsslZjpJ/MWFf6PGWBwkbVq70aJGvBs5/
m42Bumj/R7NyJomPZDjXZPYJs/yNoQquyrcvf56e4gnDvZK+Xq9Kj88nFVv671DL
FNP2JOhGUrwysSJBnwsF0MXlzm9aOn8YqLVycyz8qoV/xNPZOOUtcKehYIXzpxNU
ObKU1MJnFKEB7V4N67LbVid1YpwSVIdbszShV94qtB0CNgiyv+GKvY9+IrEa5LJn
qBnqVHeuhCa7WsyDFFmiy2f7TJ641HrnXp75OwwlY9SJs6oGIjHGC6aRVxxvdvfL
Tk0fvnu0VWd+EUj4gbaJ2nNjwPEWi5M17tqaXiqrch9HOVu9kBpp0ExEAJmehE12
poMV5qQrTJampxuUqvvrQn8FX83a3rijjd+LssA7sj7fUFv0QtWJ7BqxUxI24PQQ
sKrgDVhjRn9oCr73dOKmNamQaR7jqL4RDYkGOuy4acaRl4BWxy0F7XacA5WlHzbZ
fbUo34hXhFlsemdzaX1gegxyLcxf82ZZnprjqM3e8Z3klxB6Wc9MmBiHaHS9FaF6
pMsSI5Mwu9Qkc+h049SMJHZPqJjfSJ5/xb6pPhcphdxS/LYOe/3MYoFasmLRvdvA
yCVoyQ5MqxF43j32fUJt5GTRixiPw1D0+fkC0Xc2cE/ENoSdHWbSl6Ckah5xYH+N
zyTXv/gokMsbRY7/pSp0XMUwlaR72bdHsqJPqBB3MblfBut6JGF/BEpu8UihcCoy
RS2O6tep1ivK03WG4j1TUiuv3e5pTjok7qhnhHGgA1aC0iTKJKB6dzAAG9r3osO0
SUt0DpKfhUgzSg1HaU2fjpbzfxtlGMMTlksD8hNtPaO4C0vmsK+65vhe6okUh8yq
iF/WPKWNa7JMrrnfE//YpYZ8x647EAw3PC6s7r3aCLI=
`protect END_PROTECTED
