`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN2FgYgEypEaRhVbPpQ573QIRwK9hIWqhwweTstp01rwI
i+KyGep25OqhwPqWpc5C3II1ZaVIyaAqAWTJeN9jEJLO5r9pRK8ED+YHkGSHxtVA
XwgLc0ccWs/qcf4HyyZoU1nPloWenBHFFEj4R5X8VpDlZsWq83H+6lD2S9h6sfYx
uOFHuRD8HfhbYSIxJfch10JvY80lKQ45NF3DdhpjgcqzJ5n8708KMZMVzPgUfiIp
BDbvaYVRqZpUxl1jBEPtaJQ8Sgm/YthklXMvkXFz0pJ2kE7GPiPDC6RqWBRjC9zQ
ZvE+FY6Lymsh+L34ysnLRAf0wAnVH603KlGPlT21JgKoSt2uPgpodJ7J3Fnmvku+
U204SC6bJwyP05otisDqmUg+PS0iEsB8XjYWAWdl8rxob8MHvBIMzQIvDAazXyW4
uFiDMKfInU/SAXcxoEQ9SeM4Mo8NCUEJW3+jvqVF5yXCxgBJZghKv3TvqcipxpXZ
jl8eFubhVTawWIoW9BD6w0IrVXN3z250uP4SJTVD3ao/LZZZYp+RQqG+u2r1ViGz
kjgLiYsMSxfggh/LGMGhKLAyN98mDiwZnv5JNqD/9uFFmnZS6+QaNmC98+USmoU2
wkjI6rMNuHHpHOAX+79gJ6oFuLxg4Vcxj+VtCqnVx29rV9kX+o+x04+A6Ef1sGT5
/lYHXHDO3WJ1v/TZ2wJIJTJtEhoRHEV3g8GXO8xoDDY+V5xMAOTpz9IRHqJvZAjN
zuBBB5DIOmu3oJIuca+1Q/LdhGVkc0US4FjW2jyHRfs0ZfhKZjYr57HoskP3CJfb
RyUHER650woCZEq/ToAlbvzwcroBR7vKl5H7X5XFRwv21FyA21ZsIXosI98uyT7Q
jrsiApMYJZl40pzANScBdviq8giK6q2Kym3IqEx4BtaZp59jrgk7ktQuAA3XGXNJ
yGecXw8/D1lRxraJkL001qAwCNn2TlooHE4OD7eeNCAo9VEOcmLt032naJQxR5a+
9uxpcVbFhnC/oocZoHwiknr725qwu2kJRgTBAw60Vl56k5+PqDoa8Mqm7y5Lwt9G
jHB+lvObKmfuiZVbNfkNMsEQ4SCCH6iKarttuwpCO5X8yjcoXqWvVWYKu7r4QrpQ
issHkkZj6ohAPJidDkR2A3PsOU2TqVHDFPddkUh5BcCyfig+1Qg5D+Wqgi4S6cP4
VlQZQltW2Diw/sluDSwmSprlm1PezjvzGHC6Ac5tEVsIfHtdzTl2hKrE459ZtpN5
9PR4QBQgVMHdUaMZ5Swdk9gQSpw7y5p/ga50ZDkRlVuI5eIbalQE/kgx41SmJixA
3OmrIGAsXUT3CwTIvLmds4q2h1m/k/QnYh4aUsF991bfDj7JrOgKsonwugcCz8Mb
puc3vGvqtVauEaexosHxb5py7/0seaWp/i+nqf+59niyq4lS3sjYrOeeG5+rPxfi
Uy0KeJTnI7gozbu4Y27Dv9VWvPz1zEqD3shiJgJhLzHgSrwrWwa/ZB8u5mWx1rjA
6p9kWsFmY3xq6odwyYl9t8ykMVbf3mto+HObvx2xFN1gaLEKqEtjwaQhfoncDovR
GXqgU9DF9yoyofnnF6joNCVEjTI66C6bikM8R83QejVQmmh3fgyhLMD43cEUJ0Kt
LmMAneT2f5FwsArooOp5E/cZr66WOuWpS7aj8gDiijhG8SY78NRyd1Eq7JDJMWTt
eG9d65zm5bEt4kAv0fns3FpresSh+Wl54cVjU4FZbV7lf7DY0ZFq2rO2XXEi5u2w
3F9D89JVy21bx5AGvs1KHW/G10CyMWHvpsk+tZLi8ojbIE5mq8N1fpgwiz/eaRXK
QlmgqC1qvSgJ7NYTBCttRJ2kukbi9O4xWKLOMHvmBx/SbCU5mZk2RnYYVACU41AA
ukL0veyiVsog66YalFH7faFac3V+ZkfBceCcLKmOE71PykoKKmWRya7OoHx9A5ar
6TIngGEe06mMC12jwvyXmgYKfizc3kiS9qZ1V0UTtmaTIhiTYVNwetcKApwAwr5d
ruTs6RAX2h0YBTuzqvlzPKabphuoVQdkIATVorFJ73ECr0i3gzCqJP/e28XAwMaM
mur27QWQRmupG2CYb3ySX2PHQPug1dx/0bDrdzZWtRSF961qS5j73UlxUh+CepNL
L4RUOYVFGOajF6EYxU5YDorjrCxh11KjjqKC5Or0AZSUDYfkIn0Tr+eHkrYV8Gl8
M/x6NJtAzO316KLAsXZ9BFiYeuNt4FWLKFIujsIFK5Wq6z/YsoE0qmXacHG4qua+
nmSHEqRvFYPsb/xI6v+TIkFSqFJEUOmjTfrkHRhMdsjDwznGa4S52I86XNTGcTr0
Dis8fFrvD6eeN0VEMHHgpWLlqjuBUYJaFhiOYtN5fkyeuo6A+2ppV+xYVCKUR1Vp
Tg/BV7YXNHqYmV44UE775J4WJb0fpI3xU9fdiusOAhgjogHrg0AM770qB8dzv7wU
LtdMrMee2XZrL8P3vwSEpKo2DgAozsTQ1dmBD4T5+wHE/d82iC1lvd5unRMrA4ah
vE2e4z5ktcSKkvULOc6p/zGksjVe/5gAmMJNJCTMvTsJ7MiFPxdzwzPNtbJMKmm2
TRVhMg8EDzGdKaA9tJbSzKz21WKFPUbfAlZS5nBoahgly5qGhjhzGsKX+n+msdUw
T8udT43hz7Szaqq6zkXg+edbrlR1lK5UCoZGfK1LO/WJJgnFj0x8Nl5cJws/E6xs
6aZvACwdSYe8ALIn1HfJRBSmWksKnjZg0V9XX+7LmOn0LHkUJe+F/Tw17qh91bqN
`protect END_PROTECTED
