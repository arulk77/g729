`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMtxeSYxAgm2MwkyWlKcH732bcUr7MQkx7/WMAbCc3jJ
aNqiWvUVuqd0HkcQirc+px42uwkdDBMZ7gUdRx2GetcG/VtXi0j9oIcXPLauTEwA
B95Sb/bC+yiLS4FcLmzJMyv/yxecPtOpJVjrYebDdSoeDH0iSrBlsKe13PJoztbn
PGydQBCU2A/LNA70qU0QnkDII2ePJckc/zUSRII/S1Iu/lSvIgEtjy4wuo6tK+Y+
lSGFZzw8gvPH9zbrf+ugykLzJzB+Up8ddcXtkMuZp8QuMrsr+rO7X+epw58an1vJ
`protect END_PROTECTED
