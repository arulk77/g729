`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43CY4mbqckBEbqCOiEsZ7NU6FmAh6kGhLkywR4tScLnr
9XxsEcu3W3HUp8Zq4EX67Rt5jy/BUu6+Dmttn5eVXVpD2hnKqmIt70P9l6ZHcfKi
MCgEOzALBoduvEBVmaFoMbiDKXngBmYTHuAPHJYDTz0Nxhz67kZ/bUuMGSsq2x8A
nw25Y3glThZU+npQXBitedDTgAlNx/swxN5qvcOTZsCHfxu1rKUvT7IBz3Wkdz9l
tvtVLoN+e9//9NoQuwgWLwRF5H717Mm1QRlGUYO/FguhrokiSSjZ+booYhtc8+/d
MWGaSCm+i6YOVOtRX7kxM4dx+LMpgS4xc5KrbBy9LgeMe4iqeYXDQuDDrm1qMTjs
7GLMl2GIY/Rh1CQSbUVDXw==
`protect END_PROTECTED
