`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SX4IiUYqKQqT/itzHVRU64ggZ8UIthp9vVVqR9+1iUbO
UUhLYmvrCsCnTQ4TXRjgQtjcWIUtF+hHlVwA5LvBMfLc45ckm/3TN/TrLzaxqxx2
4kzMEyPT2Y6GWsrRktk+DQ4EsfBIl0WfRjMDTkniz1d4xA+TZ6RyIkZqd5zJNejQ
lA/jkK2DaU1iiAb9Sja1wIJw2jkhZe55nW6s0pdJzpb4TOpFaHnfqUgcSwePbbGC
WHPevxJxcaaAbLKRDYk7g/B0cYWkqCjEtRNmhNvgcOoAhXMgB3mtpA5QOs/0DEaq
n5m2stA4fGI3vvYZiVVtkrT6NBNj3uEzxcAkmusxwcdkdRDOG2mRkOEdg6kmkawT
UQDyAXg0387s0vIP+OaGqTev1Qwja9mozQEeRkyDFiGdX+/bue7qJfnFJHXdy4c7
LoYNfVebWh5qT/qStXp015zOifaqLpI88By8hvZvOAxNtnrp2rnNM3ZsVzBKs+u3
3OX31156qsVUBn1wvuk3woNpg9T5L7wnp4b+u6QGvtM5gzemc/VbvKwrQC/+spp0
qc1i8iFt0Oe041f+XYopMJQ8fPWUI9KfLJ7RIsiRgE1Nx40GYI7myWkyHnHvG2EA
gFGjCRgr61nYT7aNtE9ycvp7VLl1HCJVLZUYdfbkY+2fB7+al2tgqKpfTXA5tjVn
lKDHfnqow1eW7Onyia0A6fagJj6BzmFTsxWWg1vEFX5ZhrS9Kcsr8QeAJLpc6uQ0
nff87sdHQXNK/JVyTCi89hqz/XyyQdA9Cab7DSQtljhAhjCTAHoFeB88bQARYEbe
WR7OyrnU0yXJZYpTP8EadS9Y2jkkwNftE/kPyeC9D24wqxCkCNDogVx6/Xn/yHCR
1RHnpdGs5UC7vB5bsrRUT3fvhPXtPmsYE+3KXViP6wxG//TbQ2TZzP+E0UfRPWH9
Jw0Ew4/FqoErbomvXiZ0sw9E0e1378ramP/hqgGKSAPLAsmEUn/ZsiD1exo5Uytl
GPMl2/1no4X32DsrT5rp4Sy+ffVSGF87Q968o5oveV+gjb/OSw06lwChoukYeo0u
zV/LPX6G+SHgLy0+U0MW6cdUGNI5kIeQdSpZ8Ye+/Hcl70N5TP6sRfTBtGHS/Gcf
PziUAkF4tiXz28A0VvARrxK3EYf05X627gNc4peumxo3V88YwB2Icb/wEEzdSVTh
bEzsgjhfMtNqKgZ9DN42ZCXlEzcCr0cliPTsM9sW29L+rIk9qIro6UrLYXvD1Oas
A8Un/LxEN9axdNy7nMAXe6ZY+ol7lfz3eGh2lSrWkR7z4NNEY88GTBZbl8HGSBsA
xQbakzeY1i1rrVzoYiQvZvGZZqC/BG0zSANzEDu/Hd2yZQLfgu7JTY661PaS00XY
A3MYwUFgko8nrkWJ489IOeMSpVNFLEfVsheM3rX54DxaZRMSc05esPC6bSNo3N2k
cG7eRc/svVVVnvIAUOn3mSJbCaDCJg9/pmtCq/JFQzfGDAH7iPOdppVDchXYa2A7
Vwk5Xa3g6N5wycinJZvgPPN5rEqks2dhsa1jVRXwgW3fRKtgtv/ExQYwr775ew6S
BrThj0rlTQz1fxNvbeDudamAktWMcc/4NlMxqAs+TyHCDrprUTDp1oJiCM4M7tXG
fwLvDX/1gn34dpQDYxA3d1agIi/EdH9/BoVB/r1fICMaEWOcw8WHPQXe90mhueYG
3E4QhoM+zCqQx4ZGO3FCZms4vf8hoOPxEJ/CB+yvniqQRvkeAgEZvcZRopgSnS7e
bFTy7m/sjsXWQocQZ3VykdHn3PrAQsY1Ny4Q3wKmc3ofQes7E3WBiPR09Cy53HRl
5FSxgvgT4iAp126DxkXtFLvIYdE6zGFbrijZNEhbCGpSQaY0LPQIw6D+98BErMt3
wMWkIjgHqu7ET440pA3mnFK4XSDdiRw5BJF6P7PCzf/6CrlEwsn59WUGNfX06tol
29JzDcEwiERtZ5i0Yy5gsA==
`protect END_PROTECTED
