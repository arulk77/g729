`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/86yjwYwOifxfA0oXAAKVmX1Wb5RsXu8B4WA+jjYofy
yftqP69ArEDniXnusVhlpPmPxWQrWscvsPHSRqSj3DU7N0fDQZRKc2wEZZ2VqTqO
8Uigf1mGHYezJoNTjki4PNhuzzEOinCWRrGUFVE3yDmA4G9h12Y0Dm4DTOTHwims
WlJHHYXX0fcoCgYm1vNLRTF6c9U2PSSc6EnRYKJ3HEV/5HZ8o9FsE4UmNDYw7yoS
s3ugio30NlxjcRfGAMYPfODPEMwQRuJN6FlapRDUPP+mjBenaT+vLoHQMI/X4ONC
K9ezIfy3OHWsacA1pt7m0c98i3QeRARBd4hoLv4BxzESegZG6vm6yNBNGXXxqKoG
7xiYDRjzmkdqSbg3Mj4/8g==
`protect END_PROTECTED
