`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveH5vc0Vug5M2PKUtZ4gsvbXOMTUsgZL6ep6va/is/p/3
lIWBfX0xvKD3yQiyDoVL35l9UpUnHg+ALl2RV2vwto3uwGDz08VIGFp/gBjHLeJp
ZkLXOCRdcTohLPIkKd0OzzEyzknrTNrA0TTVO3qRr0ZPDcw3vjqEaJPALOw6Ay7C
8VFBSohZUhya3Kxfwat9aS2iEQE2isFQ/ASZhfi5ErdtQd7DdrK6NKQBni87EEZU
MSAoafMXpfzJaqmg7X18kqjJWLHlHeCwPdu/wPtuVb/SCA79AqpVGVyQTIVhpTxn
1mUldMTqd1l0YWO/snRlvDkLlt5DNabnsUQsLUa5KwLvgW4bSDA1r8QJWY1Os1JS
ieMbetx9K7DL7h/9EhCFZGpOLZNUKw2S+LDaHVQQds7L1AtQtSj1wvbbBY/DQT4l
0JvzYAP0X8fDDg/5HcI8L1lbXwzUOjKeFMaB+tscvDQ4mgwNwqb5Hu7mv7YOoXHI
6KFL8kOQ3m/UcuVjw1UE7WWX0w7QEgXDiKMLJJDcDH8XW+Ibh/XOtkNwXNWWoTY3
dcZSFcuMzWg23guqInVJCc0WPcjlTysA8AM+m8dnU4WapYOdINNPZOZX0UDly/gf
jlBdzPsttsXCqDcVNaF26gaPbQfA9N45ZUOSktxJ9X2npR2QysOj6zN4trwvniGd
dBsKH/GHq0ZJwlS2ffoj4Cu++5ePdw06IGUFy3FPYw1SSxKTaH+TzlBOXfPH6ZJx
GEWywfgHrTg9jUDvyye4nQueUGXIhMWKD40Zco5ohJ/DXDdten+77TfMLxLf8W/f
aw3rHYZuzAouUBvsuafqrjlnjlpdMVqX8ttprGT3KUk=
`protect END_PROTECTED
