`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xBkfLIojW5XRjLfUo0Ct3h6AgMm4gr2SZ7If8Zam6UP
1Hr4ULoAmjg6da8lyX+4AqC2PN53b/GTriKO1GieggfImoIGbZeKxX5K0RGB1OPC
DCLl1SBFUQ2YAvBxq/+VIVCcdZ8vzXZrvlh0v6ZcksH8SXaTNUJPYRuA744QAWjh
xgD2CWIeadS/OBHuSJGV63ofKj25VcQG8/rW5riSeeztxLlLTdnCdBV+N4JoWWZG
OQG/EFb3QJG/ornWS2hZf/ad9zIUTcmEoH5K4Ba70+kaF3QIDUMpSVxMmAs4qVli
cSjo1K5WjhHRWXTxyJmj5g==
`protect END_PROTECTED
