`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44U93OIHJlw1PTkX0ThapxuzONNt4O7u1aJeAaQ2F+Xq
a4lqW7r8LitHxezdM4BVpOaX/lXpNm7O9QWmj/EebHnnLq5RHDVgedW3h36TsmCz
8sv+OzrF2vXrB7olRDTcM2Skazm6ovQiqNxVQGGvHg2QGWYjrxHz+9+U++ZndrRK
rLZJxMG2/VmEXEfnNkGaCk8Q9WYvQ+917/k0K7J6AzH0XHsSdcqKsvPVHvshJexd
SIOTuOeTZ5AIddqAiU2wcDYp3x4wQRwH0vaY6Y9r8+xJ0swuB+SRk5G2ERZv+A9R
VXjPkp1vTIGHvpWrtW9r8Q==
`protect END_PROTECTED
