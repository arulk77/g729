`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNmaPSJcW8hvu5SJ0Nmv1JzAMEPmcSgfvNsa4vJWtTFQ
21GzLAPHGAOgYb/lT7xbHLtwWkYP6/nYqPwKM2MzYOAiA4yhUQunIFOh1LV4dHbg
9OZQdFm8s/TXEFh6eqo00BLRUOOatyKIEsf4dLOZPJUn0Orv2ft0nV2AbTYx6DGv
yda0Z2U7/1K4KVXGq980jVd/0TbW+Qulzq3dIejvFZAUY1/pxmn60wSentL7eHao
IL8RB5s3+jughGlQDRLMNGiX1SsNkYSWUiAd2l7p7dch1mS0DuEKJllMU1ijS9gU
6VF01n7hhbjXU8rNRrSz+hY+2k9Lj86Euo2mfqzIF5ukUbIxOEpEXPeidPwARMZN
+5fwAezIJH/QRWu/Cwcy+YT+LD/xBh0JJRmR5pbaSiMC08AAU7wLcGaNV9TOegxO
xMelw4qYAeCYRU1BtQTorpRqvYNfghfFLS4gf+i058QXyWmk2gJOXFl1f01x2Rj5
9VVen9wuELT4KJFEOEXX5p0K0Vrlwxvv+Q6uzYUjUoNQukwRUEWIsIkmJ/bpp39B
MDhUwweuJn5d6CzU9a3rVpByK+RBUrtlhBOp9H/b49etLKIU5frQKvWlhH/KW1Ss
4TFInxq+DaDq945dFMMpU0TDAR/ia1jzuxF5NvNxwSsYOg9LuiNzB8OXZt7BXmai
qgcR/1UtqIPjhbryq9ctpHreib3rBJIZtN+F/44NwSMoiFfGRACdCYL7gRVQi1vy
2b8j04wkdHvD/Jqb67dq95QQ5KoNlIJL0LOqGzfiC4X4g8FvF8OhlwpiVJ4/Rr33
tgqNk4MNvYEvX0MwbOq3nQRyAMu1+OsOgF935bAf89QLXqNEWSxe9wXoIaqjnHa6
bKNxykBQtsZUnngRSeEjOT3WohneyypObwJl+dYBZJMl9GcP1NUBfjW9HpaMwwyX
1AnzXtah21HzqrVSNp5/JKgNqoulODd8GB7cUqxQFWUfkxGc+CBl5Tcwa8qrWEbc
uGYeGeSv0GkvKskRur5ORlYv+wgWIiaWZHRzFJyNkgsuwrhMeMcvUN6/wrdiWJZ6
Gcze3c/GPCOr8vepnw6f370ArqljTQtgIzRe7QwOR0OUDgUVVaZDqJtpzNs5Pbp9
sXGocGYmBWo1yYs26NnHy5cQjoTQQ+5OSUHjl6Pn8xXK5WrgO+C1i39CwgdeWoKp
B9NggYHWeq4HAXTBe8rHij1T/oq++BqZrTXzSvKYO17Il/QQPQBEbhWQs4W9uNgg
XhSw8B48HKObDAN65IhsrJk9FH0tpKJd0E7ToIt6U4GFg3wOghHvJp7+9KonZ78y
F+0UoAoh8zSboAvJ8wIoUMfYs5eU6KN+Jae8dkKVTOkJfNuSG4wq7s0y6ilmmx01
KX8OuHV9++3qx00d8mk5uon/lChrz50K+hA3UnTpFawfZFfmCF7O1px+8AhnOz31
HnjmE349njZ83x3oN/66iWmUIS3SzQuUkf1EQbJv97i7mEdikPV/reVFdhCj0JOK
GUU+KACFbFSgnjJfX+IEcNNJxTg6QaRU+Derh5WQfYT3FlQSN4ojc3ZfGDn69uf1
yQWQbzH+qIjcEP0zHG7VC1/+sqeNE7G+f4lGcGal64BVdeDz3mwL2siE/V57KQ21
2T0kwQLg8aaNc7L+n15GjwnPIf7yM38SCj3CAfR098641KawHY0qARwohhFiP8ys
YkQf/ZMlNF6K8irCFXZIVfSqLocfTUULMNlrsrJhVsRv8gqCqfV0bkduD1xODSja
vIxRUhjBgIR0VSUGgVEVCnMy+puCqYUhiyoO3KnChfIowZpuXIUg7H5UKYSPWtqs
u1VAq6OuMLutK/a3oGN6Xcj6mEMFI7QY6MVKUuZnNWkLP5wA2+pboVYTQOFjMqUz
T4UMWXUTEwlYNcDuFT4tRTyyKn4a+x81EI+tzEwJhuYINnvCydypZha2Azt92t3T
wEHXwbucG598eGMvZtuHkGntTpdWvFiFGqV+E8Ld6cOqN6xnTsDjZv04HA/hxiZF
6BLmiewkTkdhfpQcDSt7g2DFMXcI4Es1Sb6TVqdeYNJOy7Q/e6WAaGslVaBaVLvg
paXP4+PzlUs8QPHV1MZkSbgB8G7D1dWXeYVfE/gtQcqMeQA2bWD2YZJZ8n6AxSwN
GyvBJO9kXOYMTcvVeFBOT2XhfIOD5w2FtqCaWUN+Eo9XQU60cAgmDdYI4OLv2JGF
U9QNEgiEV2vTpflda+Oi6EVaHQ4VQZd1W7AYXeTnzEoKW5TOqnIpyzP4As1FvDa3
wKpRcbm3DLtSLv8IfxtnGP9UvnjNTXIGlWTdXSuV0o6bEzn/fjcjnv6EwHJ3V9sZ
CrFsWtCEsuDkw2C8Mui2NztB5nBMCgAhxqiScTSyTjVhu3AroDbYrL0/OLRtQi7a
2SQsXL5jnAbMdJPDMO2gDHHnWLhFqKJUb8Q2r0vOJJ8Z2cqaEmPgsa2SJ/QxYRbo
qv5ivez2YYt9h0apxUV98r0aYq84x1bp5GNbLdROSCSQ2NlITfMWHqTynk5tQGmI
cnYYGIFXDCHNHhZlevXzX9wq9heYIkYSfo57kz5Z/1rl5rR9czicK4ef8PEdg8fz
WTitGcHuiP1109Z03AOHiRKCfgfweUBggT9Rl00RSDIpIzrPNZsV70+PC+ulJ0Xh
kt5et1kwbKgXINX9KIYtlG8ycvaeLMX/WDrM7q53vr7DrQrzBbLlzL/77D+ym7JR
bLW6+M2wopw2jgDuimM+YoV2IAGzQ3Ce11kYto0RbTDhupf8Bv0fiIqnn6WVtKrk
9L3lZZDn/e5AqChGb2ZFOOA7EgfN23iqlfOJBmRrz1vSdgKP2xCH0jo+GGtAu7Cq
OjzrkJGCuvyCY3FB/yqXVrk6TD5lb+5t5sqggFH+kCRcvhKL9Z/O/QLgq7Yll9qs
PQ9KiZ6p2bumaoDAdVAcBk3ffNcVpsjIO1shzSlrcC0EAtxliMkxrcHsRhE/CGqk
x2LnA5G+fHerfNlOjDebpMSnR0mKnyxLJ9xqiLj72TpWpbkSpQ0zTuak0Uo5x/+1
ZBpXlDv0fIK2zv28iQAIbB8bK/kQRnEey7aBRCM8yVp0TAuJPywerLKSUxMBP4K2
kQ1HMYJRwKinFUyHeyYCwdeqwL4T3d5plYAnEdkDm6cmGu8jPmJWs08ifgpBuPWD
sw8ej+vglew7yPGCi5bkO2nxui5NmsBq56XPMPRPnWsau6ZJhbcwnfP4Qh+1neGC
1UcuUKN00duUGYq3uKJS2rA0YPt6rjjUcy2RFkI9KnmrwHZlLbfEteXu3+c2pBHK
dinHce/z/ST7p5u2lWaviSJiacNL1j2DmRrw2FSposqDZj8l8DNRPwIOhe86CSKQ
WyVdJWNhp/LSDW0/STeTUxr4owBw4P7bflxIL0BYWsWKUWTZKIbrVzTEPHSL4Zjw
685QeOsv1q0IfKJJ3WLkyr0XUcaQJHvIA7Wb+ej94TrFk65X2g+Eha8SM4q3Usvp
TBzNJGp0wbghtsMDE4u7/V0RLIOT6m9o4OLzqbdIWjeD7DJtoLsmhRe89voLfQSA
nbb1wd4YpOuHCOpY7ON6XHU3tiH5wwJ5MuFo1dTaIGut1Wy19ZjMDZQfByfeovYb
EDgqKd79AxdTSEimy69BBzkL8DTyY7sgDtHmsCb6CSYrCL/DTdxIr+U9yGhfv6Uv
KK3A2JYEbsr56R0QVx1QCa8S4WA9HNTb5K1Wj5TGDKSnGZfKOZuyDmMB+nuE9+kc
Em5+hXyrddo6E1xsiBUBQccdZNZXZY5rFNcOTeLw3g27B/WC1nH6k/U4YgeYr324
ZDWsD+rn3GG6Pr75sO8OZvCNZcZPqJFGaAVHi4Os9D8riVMAWE6/eCglinAyUTv/
Y8NbvLmD0iuK55kdq3ArU3dtdvJtnFrXl8JT20aTyju6ygKudI9RyTLSRhljeCPS
5THDf6h+OpTUFbe9QwHXbcMlwGf9WhImpbGNFkmpHhFCpgthfCyb0deqLNOlay2i
kGkSKs4PidgOvgBhrnjnYNnPXKNIqDZ+mQaiY9aMOrnec7DEHTYZCQE2X293yNMK
I/aepY7iwVu9gIuypNceCHiwK90A0IjX6R17UxShv8WWiHCNE1MT1pEKJswTBojS
yrL86IT/WKBlRx/htnYlZDd1wcbktMug2YbqAFg7aAZ63Qy7EsZ8Iu01Bdmczv/N
7s/wTHXEXY1qGpJekVPzsfLtH0SQ0WSFGhs6zlCy40oykGC8tmh7TUCoiv7mYjdY
RvCrl884mskQX9QOqc0KS7utZWI590wNmjxRuYZYmSHIZLvUWSd7Ve4zPCHfIll2
Ypco5dLjpPz0xSYLvh6J34DlAddpRuFfzoQ06wloIqlrUwqNLi6RrEudts+FLTGU
CPEUWOipG4MBYopKYbwjPhfW0SrsxzkEDo630i5/jmV0zfzKWiinNNeJWZxgeH3d
tBbSKhws8CJ2Bi9kd3t9pcbBuzdADn7yluPrm7BWqCqwXGB3ajRxDXd+mDjOfaVw
n4AqInYyHFDcKmSAxxLXufShj01OuJZ6jjNftxbv3j0TwWehhVPRKqnIhzAZPYKQ
ijqj59nT9AH1bOoE63VzgVUHSICs9FvBiXhdgGKm/bUgHEWOjZTwXkf+Im9MGZ/g
89dh62euuwvLrG5Cipxy0q/c+RbCw0FWzKQMv8U+TiH2vMYg6YPpzxVHqyQrtTpx
fTj8MhyNgjoktBBXSu4vKW3X3V3AwqaJpSn5faQ8Pp8U2AHi8YbHovjNLnEomTHG
2312O/iB8rfnS8mxFGHTIIY+s+EVMsxM73cf5GZASGJPmQuvvoESpTlpx9p2hWLY
Vjl6zvvvez/sLOqaUdL5pqAXpfLof/tsXJiaZzkrhYzIkCq5D+7bI/tbTIfrolkT
Vi664EGjDR9Fx37ZXtAWMYgrPPSeC/L7FFhAkO/9emfiYKERKneueRvCL5bKo2MP
1De25pmD4YABz2c0Zj0Qup/A7RXvgcJ65phLzTq7EKFt2yXASTfy5BByvnxpCzYX
ZheMUZzETN4e3BKi+dR4xJmwEfcMJcrVQ0P+Tw1LGJGVWlKz4NNFqUB5Nh8HsYFq
VRDsY1r44TiTudROQqfau8TUtts7RuoAw/tM/R0Yc1VRDYimsH+pcPe3LIcTODXO
DQYKrVe3IEoi4JjZC134HLs13Q2ZX3MUmxdZFHm9bVtWzPTJGFbneuGKMr5Rjfhc
hjshZSL8J+KH4hPCIoz50w5mCKqf3M/njTAJzaJTHmIqajFM8aehO8xTDaTDTnaJ
32VB5udq7/qO9iHOF889TGK91WBNiY3uFvHBIj6cX/diAOHhImVqP/XZbIx2KoSI
McbOi7V3klTTVW9tGAMbY/C0k4uDpVq151hNGczpNzJW/7UQY8ejEVoMoHe7hM5F
gHwHZJw2QqbiqMu6oR9sCUo1QaRLTwKx+v30Uu1OOoQgLfcQj275Hy3/KLFD1TSr
DhRCoGIhkXCSW7DwBJsuEQ/cQpQOef43/wuwdB7g3QKdpvm+QEmC42aloEoiqn5e
AiQGyyn/MMc/eMB+E8Vgsa+cvRh9P2dW9lIkwh1IpgytKpZUGtr72D+VEMzNyKcw
wU49YvKTFNIl+xgzjQ5pwOUv4ReeWI4zZCs6fEZzLdaRKeoHJENyw6aMABygOzbR
OTyyBTY6fAeO1JOiPsMvSD3F7fRtLZB5Xs84IFt4pmriJMGvSyacWMtF65Pb2iIW
E4lBT8KK9V6o03BRdh30Em0ChECjGvb1cTZsobvp0u+CBjv43Vc1zsstJ5ZYo8ct
j8xBCGQfo+K2UR0wGQWlPfFaGOKP+LKFeXv4h9phK1vCcD2t2YhT0EnTEgPwn2wy
2DRaTinwBoOBs5p84FXl9kes0A2v2U728sq0ldjV/0P8IkGE6YhZR7yJWB3PRCCF
bF/rQw4aDx9kWLz4dpndDHViWHB4abVgSqcaBEfYChIdlrZPsxaGzWLnaSOck4G0
AZzDzVLuMYW+Cy/mFgDTgK0voRJA+ZBT89ljwE5q06yPu9kH0YhIU7lxqjkChLJh
WkZC9Q6D3C9S9veeuTaxUdaFJzU7O2N+5ztNmEynvj0YzAI1OkjJuKMStqmRL1SR
QTUBG7kpG558VPF0EZvLNSFCf3G/S0YaPKPZv4SdjAIyOV2bP0PQbrunD+tKWFAs
WlbZX1T+8tUpUU+s/46tzYszoRB5A8+uxzRFfqU8yFAiZ4+RIHvMUVyI21GlGejv
cbTGO4U6NDyquzcpZZsABMv8RKNWiAo0Tu4UJMkwzK5NXJSU97sOEupPoHp2ULnx
zC1WH7R5vAEjKF7QrvlSQUrveiaKx7YvKl3bjI6l/fYduThhCSV6aUZanvpjiKnl
M8P2MDyiF7qEcp6r/XJTuFu697zSLDWl/h4za5NAq11xu/jSUZpFWbpr0dYCoW32
3f9TrZeSDYlb5qc9FKT8KQSAsJS8piGDwyTWes4Fmt3NHNE/zfZn3RPufpWzmaLT
/wu7NHUKw97Gnv93FfxEL9piga50hz0bV8Q45qnfGmz9uujl/WQozfsut1IGyOzA
6yazsY6t+z9CLoz341v6Ttqs/X3jnr6Ob4yy+saV5KavfpyhZ39R4LigsxD8pHzK
KpNJrfkdWs2zidDZOL3TFl7KVoR8ofZZpis9x7zvceeZFeYc0Yq7dt0v4VaiWi9Z
KWfNgtDCrfczJNiN//5nGR5dlEDOxvIg36YgiKKZPyjK7vHDdYAnUCo5wSJrCXef
e448rFdY9f3nWVyyu1WjnJYy0PgwM6IpTd99m3BM0A9hdfGkALPVvYbf9+UFEHwL
jgk1HqoWhEhFoYzShhCn7t9eMg4Ejwtf+3w+OhPclLACs+6FttWulTm0CYml/flz
c6EOis/UjV6QmUUhj9v5VbwNBIJxXwVXd82s+ypxB/mBwbRFJLDDkBjDbl3cMKeX
RTxqPWOUaZ0EO/9balD6pxVkvDLRF53oCWKpapn6bLvcZnx8vZUIwtqxdiSRUiJx
gGLJrA5aG7euqv++Zt9wxLqz7dCGo+Vkv2dfZOyHCznWpeAD2hh8ZBOOoWRxIciD
jPyaqYdXTLz8hzVxlmhiSgILe1zjSlyXdE+sIdGeccfpMIXu7gyEamjS0whe8XFH
DxJ33mee/RlGsjM26TOc6OEefydZWobiL3JLIfUTxm8Z9C+zkho6UlfWJt3Fpd7x
BY5vrLYq0Rgwd3P55t3cGcygRhw3TSIlNsncpprgUdyIk4gDULkvgfZcPzRKZF67
D4cJ9sy6AIpfpmPnl8tO8v+sesHOZKEUAVq7izdKZcJX2vRGY2CDGTv/qA1vf1FX
ZQm+CAVR5oVkJIIeQ+gtd8/Jwf4mo5INAb2+28JyRguot1yYkn+i0BIoRcV2jkat
Zr2Zm3NKpdXtpMJnXiAxtdVPcMRSl/NgDLiM5Eu4l+n2E2ui3v4hQse31mEYC1dM
qRJpJKvdjrrUsOVuvVndWBaBdCzOS0Bbh5NAFP0HjTiR46KW2VYr2ujoB8lX1/c1
TTnS4HRU2tse+OW+P2R6YJ9D9UzCaNUf+7rnhqHchzkVvjB91W0fOdSc4frT845z
QrRw16aavTkQI1uB5bp0SnMJ5HV/hIalOL3j2A5luxMtPa0Sk+nIZjr+czSgYFwn
HtAhhMAP3tslzW0g85DyZssWoSQRGin+s7luC1LQ/pCGvHeyyWnzMaUmBLz4+nEx
jeFi2uvy6MbP9sz2rMI8xcYSwbS3yjep8rxYbpOQt0/V8DICMkz/d+RTGLslg2b/
q+ap/6vzl8oGVDWUQlceJ0sEUUOXuV/Ig+jgWGEPz0Z4oj6eCkADJhenVlBh3OXq
uvbSb5Gin7TfSTy7lbOL1wHp/W5VZPpDjwY5+W8bEOfbTpZ9aaPyilpeGVumYXh6
1OOqVxtlfQD2vN0YLPi5CrJDscBPK+kQmKP9Y78ExWRkCy620daEa/VS8o8VBRmY
Jgg2IZnLVhL11pfyo1PU+E5nYlA166bQkzzL0UHt1LIi3KX6nUTKBihsH+uvtUp/
Ijf4RNVbpitnIq8N04K2nAechQjJ/jDSSgQA0MesMmH/XBfqcLK1tKaqZDknwu3s
lt8baUNx80Sf/jEUKJCVGpGzen7sVdicK5jyIKnhBi3eDgI9TWoP6T8/vsj93Lby
XXyX7iwxhcMxvinCDP66ezJlOaKVkBKdu42/h1+nEp7KdG8/Mnr5guJJX3DeX6go
CmaMWzR8Z8EAJ2Qm57g1bq2g+2uV1PscMuA4rLeD3TPpxUkEHy5pMvZs1ljOQr8G
3IQrvv066VtpSppGJrUritqgey1a+kzbWMoVsvfBuzt2nsGH92Lm9+V5kqJ9Ngf8
nx4fGP5XxRs0DW0yqz1L8fsn0L0si7Np5izCdg1mrwdOnoTynY9g9Cn8BhxUYTQ0
OvekI4GvGaP2Eh4khcozxwXKOE/o2fwOw/n2vS9/60bjRSa5R9rAVnOkNQ/+aWZl
mmsEHhIs0ooQfxaw175qGHg8JszixVvpKCqeRbu+yKR7dCfJx1RCMIwyJo164Cxe
PLy15H5JRDociWYw06h/3a8N3RT6JbwOeFvmygmYhxcudp2A8JFUtyNWVewuzXVm
FC9YWr1UQuLKesWrENwz6JY5Du5RS+vwZUoFs52uZ6xFU9NIZE4dhELHFHzTwHR/
Au8IlOB0987RW2V7LaPWXLrUj4oR1FN4w3C0HREfoa7xVEgHVsBc8Rc/PrQEXIh8
S5ojMorMziEXLKMeiI5H13pzbKpEnrAvyVznkAGlcjbySF6TFezLqF0owmoiL2Si
PeNTjao3A3ZD+UKI8gDToRfp2NspIy3pwnZLymAIaJa00y/LUIN1ejMRTW3yRNCi
IYuwcwWuiVPlWLomZ3nEf9L906InnsP0SUs/DX1YHsPt2gqbGcIDhsU8m8Vo0IAQ
LxN/sZf24UpOPwum2nwfOPbyslBK9o6+iQRo+BRu+VZFgRbBrE/Gr53gW9V70J81
hzEZ2sn4APj+0Q/IaGNOf8hqTwwnkKTVVwSRFi9UYHcUclPe+zREx7ojAx3jHojt
9BWD8FZu+AnjNDefLGnRC1XP41RvwavcKhd4NMn7XPlxvUSYhh9SKkaxNp4ZqgpO
W9aBmX4SW/GHIlJDz3g/L8yuhzbDqorD+p9isPzvcND76fAHFPDE0hHSExlagbXb
bWHj75fU+URSwhPBTvdnkTO6+WeU3s4oUWoRPgwX1tyKokblurbe2TmIIjRSN9e8
CKMgrAUdJqK+ADDW82TIr7re5NEk5ErFo/Yy1JXu9qorLdOs14KUhMJJ1vqUdx8q
/hmUs1Z/TE/zypPBOrgSsRLtAK11mQHgtnn2HdofJMg3XVpjE6onFYhsAdSJ9g4U
DPDcnLUN0SAbXKnW7NU45DODTtupxzjscd13VV+UsqZZUnbW6OLX2feWmkoxkz85
/mR5tDuY1sol7sB9ervSx5Mw0Tj49qMLFomNHQCFktUuBGRPJTKxOLLS7FtcGhsq
yD8b2tkHBcrB0kgRMMcJOC9o2lQ2EtcmrXtbY9fuEJMAEmeMwJroXInqc9XXrxif
4JzLGYhUP7GmWR1lbK/s5AmVji94cgVyiA+71uNCQBE5D1jvH5eb6AxASwArCNr3
4jLYBmZIkFyxrjlXAXKX3nctjBz17DoYcKbH/UW3dUxpERba4RX3wul73wElERN5
/JaPbheUq604Y2F8yL+3Qal3lOpO0YCyuJl8vMwvLofMRmeIBgvMqv530iLGZwNq
HmE25xhDMqxf6uF/tlNRAyC98gM5FWfM/jQWIm+YS6bFaE2WG/+huAJJvupgtY0k
ShLfxa/DVYO2R6/aXEMTLtIlLTMv3qOW1qK6E8Meu+PMiX1L+L+s+2+QFB9QIKQ6
yuNJT6ZMxrLcTYdXAFqae0cCNxcpqBrO9w6IXbL7As0NDEjdlQke74JhZPze/4YS
2uMQIeKSaE50GB+fqXI60jqx23BBvNCnR0pggVqbavaoQ7b+O8wZDMMDEnnUe/2b
r3iwVmiZ++ifLutHXnRYQlor/utHsfLvCoQ4FEt//18rnvuAN3Fsos0h8t4J+hs2
yWuJQ58K4sglITZFlMxzUvbYb6e65JJvXrOejMcEEP3GOej/IiBoM+QYq6PALJcA
BFsWdm08IkC5UoyLJMO9JuInMG3NxH7GIh1REeZaWmCwf3ne9jXxEChvYaN7kPaM
csqR136bysc+sLPnHA7v9JhRwJ8VPSDPVzfqD2MQcEsiVmEv5g5BTq4aAcWpZAqp
n1hTuyYmXnCbFZbpvO2guN8H9agEAnlZJe275e+U6IV9h+wt4EIFPNPNXkX9nGE/
+KMD1XIwhi2x3tNWoh4pgCV7hsQ2uQm9Yhg1wTA7IUXJsun0gbL9nJs4dq0Tqo4+
MWtU28oeuCQ3AtwBTgQ5rhYOcpy+WWjC0K98V2SwZOpT6NO/lGr7dEOP+aG2elM8
5dG2RwwhxqU1XBbu5TEx7NcR5Z44kgAtJ5Fn0iOYijHQfUaWXAInGvK7nO/KUHSz
J8vgu2+trdCCIz4dxzHZ1qSRLFomVKt8nkt1X8edy5niobW9nwniOOZ/a6MsUYow
odvKWzS1MpxOYeCp6dIL1Wo4SJYwP6lnYSNTYVmKUO7T3WOcpDHeDOXO8eiWuFBZ
Iq+8Lii3kQG+gHR/0/eNlDvZ2Av3z4f73TkJvebBHLJ88ypw9MqkgNy25i8K2Rss
fpG5MgZpJPhrHVBk1pKUuQd64Xlq6xfNHTOzI872d7wkGVCDuXZFtRWxsYwV4fmE
2izFRbH7g6O4poGN/vtRp9J9hha8JSQH/5eh4UR1uqG+80BvwkJh3I4o6MtV+zYl
WzEFfy33xGPWrfjzvBwuStnyKSJKTWQZp/2RsxJAmntpRqzcTz12Yd3LL5Ucmmjn
MBxb8Vz2Sq64EgTtXReNxsgzUsr9NWkQwA7rTJnKuD8h/i6+rvN52NS8fLvjyRSD
gDv7pq4O2eQMAPmkvebVvmhPzoWtqtCIhEnkNJWb1OWdp9+8rTIbNqFr4CYbCj9Z
DL7S5BW9Ozkx45KV2K9a2dhfDZmbpS9zJ1LkkE5NaBxd8WjGFiPY6r58kQDhBi2P
dTD3HetG6gE8abtgx6GFpvxJ+HV1ZZGyVFqyChwfMyQ3PH1eeBKqTk3t0pxmy0u2
Jn3fjDoomDwIPhQyp4cZmmD8qdHNxvJ+GSySABf/Cc68CE2yoSBwae8sSVCAP2o2
BKJTSdYicz+/m3/MGy2FZSuQK6wTzN41mmJIiAQnRk2VwvJ/MVgsvqxS6mB8AlTO
R2g/Wgyrq5jFmBuLegX3tXcVVnzQWWOaR+z+bczjY1jwsJKMSakwT95aJzBimRGI
Ob2nyFJvbsh8tzPbJ0BJHUctVEf4Oi5HDdLib01Zxo/CNgswwMK7OeEL0zv18nLT
/U3TZILqwhvAWLbg0m4b5tgxX2oQ0zXXVPavdzhWp4Z8AaUNmS8GqLLKnIXhZOy5
1Ra4l9IGsxwS3ca1y29I38poSK2c/yQ1GeEIf57KrIqct8Qlc8PbXQvNAcGVqdDj
QdP5cavDQKNEEwTyG5/klxoLnzaQ1V/QmcQiF3XVAXsOTYo0UqpRsPv7iiYnyFPB
JBu0zPN10TVV6EB8yzMPCFUtqC58ZahYxqWMumK5YmqEcgAf5Ywmvpeg1EKCNLwa
s/R3oSUc6pJTU+mHpc5OnXLURQYqG5EbklVi3YXQPSEpWFrk674dIBuWEOOYMxLz
Od0/anG76/3Qan3rvyiMSUt0Z6vVJA/BobyZFX8lsE7+yd04OFNByaSWSa+Wmamo
LOULCWwPOwcLo/8aDjeXJUFUp0iC/k2E0Lf7l49Ha4yXBSPqS6orL1aR4qIGvDJu
+ENdIVuGvUoqwLCNFoQHhH6RG2fXOo/WJtDsjjwmZCAbUS2XLvBdHMaTHZozsCRR
kBkq+kVsE/HxIllOY01N1036rxsjaAI/YoOCm0qSEle0SD9OYEW0a2y1njkYwm37
ZW5em6x1p2t2dPYnDwDNRiAGvXhRip7Hkewzb6XH2V5Kuy2zU2bMZ4hS+UkuysHe
kNdkoupadmfUqFWqKWc/bQMltn0OTh+Bl1IBvCGZCUBU2u7XHDlHK1p/fLHP2wOX
1Yn/QS7a9in0cvsSAVijPPIhu/LRnIWr1sDWTdIO7PAJbCvl3rv9qkCZ7z6opZpL
z5Fmoy8WL92F/fPTvWNe/6qJ8cQcr0905jeUeXjXVgvi1cE8QlWn+ZqyX6tPqRvN
`protect END_PROTECTED
