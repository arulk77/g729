`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveA+0fgW4C7mX0q1fgaNromIr+mYokp6MdWSfV6KcUncN
EqGMkVLT1ftaZA8AP4hZNJ9Ewt+TSTr/iJjeHQwN5m+nYroNpD7m2DyA1oLfzEHv
OBu4kb/XcgPhBLLYIBg36xExUufZ7jBJlvFGJVtwZ+bz/Fz4XQwfSkNCiLwRuyyi
lZRU1MTwiPwkFRxWVmGAcalInhgqWr+ENowGEG6Q5EN9eaCbRo4fRDi3a3Oh2lGX
eVdkMgiWLmT92+SQ1hvhQvW2MQOuAwDeuB847XMahhaQrFpFrU2g0M6thZYhCcgw
5Uzdu2mIlaJBjF+qFS3sMqs2xHcv+J4dxNqs6x1ZZGHT/kn92YUD3wRMRk1JS1AV
9kL3aLaEWpgnKo/6sMP20Q==
`protect END_PROTECTED
