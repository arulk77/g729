`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMT2S1Xl1oLNbj0r2FurmfuHb+1yFhzNvaoVQ74qXlcF
W57SCsr4HycNQ61sUTQ33Anhvo2xiYKsgtlhG7M7jqQc/eTu5isUTinFIcT2K0rd
e1HpVir8l3lD9RTgr96e5DX+Wwk2NG53Ig/8CaXYBr8+a2hmypzDVMysWlcIitmB
aTrEIQ1pQCnrlt8fs68fUeTbedJkRCmrWP1T0kkXyEQmUyNsVYx3gyCpRUo/Adxo
LpHUXMn2bxVwEcixzGRWXwGBWypsvKsBLEIg2I8+q+zGUQw5Wc1n4nx2EcqxC/lH
6E6b/XkxrttsYO06MNO3h/giiRnE5Miq12JAekLfLQcWLgfJT6i+yjXh+szsy/PC
4WxTN44qOO3u4pWhsP7WgA==
`protect END_PROTECTED
