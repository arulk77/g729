`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44NDdO646LtBN5CwtHWfQ52Q8xzPEPbclH4ETAQbDwSU
kVzaaeLMk+BnPxlSzvkXYSwalRXPpZRd5b4r30KHIzo6VgXw3rwmctR0dxMSH4d7
ShH5FuxEvv8XXQXJa98vOiQXd8aSp2yap0mwbRLQB6IaoBeLJ8wZHQ3K33xlAiQ+
QDXxSquWHA3tC8mVO+cTGusLiDr9gw6pUckXtjNXE1yxqS4OErSpDcHwgtWIp2C5
7TkR0PKdD5jk96cZsn+poLP8kiyaPUSI0CdZs4PgciY=
`protect END_PROTECTED
