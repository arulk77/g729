`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2E8syGDBx5W17lqM3p6DI70pXTeNNzD1ltQWXCGzN7u6OzcC79K+GkwlZdqUtTsw
dPAGqdbBfFI+Z/JVxIQidTsoRmnr2b5FUrb2QIh1sRa+lGcmtbha2PqEr6ghWwKh
ZLNX1POD8ihswdHw21fFAN/3AyjCs+57s1VeaOx8LHpUQ4bbJqEI3o5IIngCGE0B
FhlBfltz4BNcdd2Hd43el+0A0vY+P3XM/Wi1ZofxLXQBTaABGDqG+DMOq3xlhmBl
HUJlCJeKuPaF7oNesaUblPmffMALbvmndHBoXnxuSjYZEiSrg5vCNo8ReF2v44P0
oLtddTSfjGFmBQH4fE1iXgD5VO+bQASc3O+IxYRdwVvQKrfvo7ObVDsAH5c+PKwn
WTX81SSrH9RGWFuhpfZOYIktNd6gtEm6RjZtnGqSPfFy6v2B8OwsofBBxg9fiv4p
mDDrSRR1j/+ER9gLfyqJ3BHGEKjeof2Kldi3QpqjEgdpnCU7nSC9S7Qyl/F2K6U8
UXkHJTXttOP9UOc+tZpPP6xqmUEmgU1MSBp0YPhrmpdmEy5dcCrFjqk3nKzNjtxV
YTbdNKzA4vz1UdyF3wUSj7HUpeqtvkgEIu4mvdkTwBBFPnKqFuJgi6zID0Y9Vi6E
`protect END_PROTECTED
