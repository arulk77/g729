`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yqCsKR2acQgxp8N3gTqEQVzHB1JsEYuLk/He3bulE5o
xVtFkY46c86Uyj5kQeNzUbtBIYVx3OyNC3EQYBFTVU7E56MAPW9GFa1xV7uOWRXW
szuih8P8LzEYN0SLVnIHLxjB4er8r0JDm7WBid8gcp0TgKTiOh9YcpaZSwmTAjPr
loR6o4MHtpM0w5Jt+/AD7J3TstPgj85xl0+VDgtOF7bDnYFj3LJRTD7lYDaUpoZQ
5IlaMekaa1s7VQTc0hio8FIgG97iWm/ymfo9/mEM5W/axhHt2MCqqiA/+cPtnkZ+
ZOiHew1XGi6+5WHr63to/APLPKrXG9MBgnkQjvMtWckiD/AoLYmQqWaUU+9oozrB
1bhFtvMv5Lm+u4FFqzmJV8nUKblP8P0+oRt+yGOp6Xa3KP9QEC2AjLqebkEUmGFh
UMMR2ABa3t/R6WRlsD2jUA==
`protect END_PROTECTED
