`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
nEvdoPW3YYjcUwmsGXV+QuQADm7gGJMFjM/5yUpMWEFxNERg4CqZ2ZJxYAC/zATC
ynyJ1eWciTy5hHwT6GZDEKaeetdU8pvBNOZseht/PKvCSe00k2Uq4GYvXPNTwm24
wnkpCpp2nwlw5G8wJ8LDUU64/Qptyh+fi+zBRxWowktH396mr2AhX3tx461eBHKm
UNSeUM9SrJja8cdhpyaynzaZwMhaEX//LZ9c2TVizR+bE6eHu11yBRxxbKcpCDdJ
KAuzZX/qjRjeDSVlK/p5P0srraDOvKP17Qk+oOqT098PrvwZSSmQhHID6gkKgznC
I1P36uaS1/dXoqUbgRWJ5uegPJI97bdmyNDViR1MDxI=
`protect END_PROTECTED
