`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGr12Ol5+iCtrjPZwi+fC0c+Rurd4K2IajF071SEFDXn
Zc2kovdv6caw6eTaAv/vheOIM3rKomk8F5DuPu7+uRGptt2bhXcUOMNx709INU+i
Ep2qrYXHoyEuY0KaCTJ5FcZ1W6Si8GTCTzZ5nImO8isXajypM59cTFrMI1EmtyOA
SWy7dMpRGjrgrmrkJ/I2N9WM4r+lGd6t+33hi29rZbGQYHCkAzpLcHAtbpf4Jk+3
`protect END_PROTECTED
