`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePHAzgJruB72XYzl2dEs/a6JwnjGocHUf8XeuDNDOEIb
Rsu2I57LxvhCJIKM+RZvSZxulH0TZ8huaNbCASBKGzSNO4v9Z11luvlAI771NlGf
LcfgmWabveEbVVlE6k45+C6nUWmEfxonlnc0goxtLpoMktuR5iJCMaIVMqMd5f67
SKyHXr17zZ8SR82F4iyiKZs00JUQAei3MwhE6RA5zMAbCbasXI8yF28LCd3Q79J0
rl8FnbgLsMIsa+Z9VROiGsZK5EQYWODGb4tCSy22DxOYMMOae9VcwLuOV8eug22M
HqMQJbobvHyGaJ+MBFtRqe2+3LEAknCMgsA3q9TBy9yPfbjWSsXl2z86FUVmI4mH
bjYeVyVpbAZgAFmjVx7RuY2Cm2aMzftkV1iKFg+Wb/it2okmaP8lNl9c6cJNFnC7
5rUSU/7l2xl9C/fw6zLLtkG9WmWObGruuuclnfc611UEknqJzg8WIuTjFXKLaQ53
t3+r2CEy44q//Us4xEj3L0S09IF/dcRrEpSHpngBbLc4dM7e47F7P3iDLckhX6LI
Pz63FQOf8+g9tjmAs7r5GNhbgiRZgpve2CaFJnm816BOvL9F7TbRQFD/ROvtcAWI
`protect END_PROTECTED
