`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveO2fnqrTfBen/+3etUuHWpXvL7gUcnSOevCxLjEtvihg
MuQ26zT3QpeYNJU/iManWTb0TXPEdFqEKtYVixCZcT2wAWAAX7hJ000MadS8ZcbG
9GOWM8WXkHpZTweIw9dSvfshpGQ/QiCxDM/joImx+nQgcsF6uxw8+PtMM5EMcJwt
KF0G1MLyGtKux+cDB87pR27Zr8f7ayHNt6irizKzN526QRvYJQI8z4F0yHNcaCts
`protect END_PROTECTED
