`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
AaxVDLtJXv5DhpU2V6JZevTobzZgoU9bml7QxCIRCwr7SeYZRj7qu/Yn/Dz0mDqI
KyZF0sAV8mSDVWKAGNqxVM0g3PMJUS9I7w9UuuUwNqngD+3a735SjH8++kdArF4j
yiN07vtn2hVKM+uOHWAeNbcFF5+hSm9yPcxomZwoj5aJPBbCssOjS1aFSkd16+Wv
W6FSTP1GA5oz9WJ/1fu0bYaZ6YE1D3r0obp1ALpKaPk+Gwz2iGm7Gz4eG5xHXkJO
blnoguz/rHbwXtDa+4eGW2PqGTqfLIag89JMRyY65DVe5C2D/XtvMgUDJDsFI8d+
USz5SkrfJ1lXnzcPBxG5kaZ+WmiEVRXGbukLn2duDj03E0iDk+UKjRWeqBjvrZjZ
ecGnBBOXb0Jzyye3zK3+EAfUNasMXYLXWrZuT65Z6u9QUsJHLVN/jnm9ueyUtqOG
nwricWp0+AMXN8RBHUXT4A==
`protect END_PROTECTED
