`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDATX8f/twJRjE6RjHRZ0rRok1DYAdI5dj1CfUiMYkzSOZ
0/QuWk/GgtnJ8LQmHBc45nUNaPdT37dP18VaQEZPatCOnzyNvFEWDJAw7iimdEwM
vnCTA4hmrB0DB5MA/80vxPg3LZeFxBECGbCC/EvogP9s6o0WIzgJ+puNu4SawY8L
kfaypbNwtzCpVFWolLLaD8CczuWiaxzEocTyU8rTZXORK+Mu3xtyrtDSy9kp8APi
I1ct2Zq3dB5T7jP43FzVW3+sTYxhHPH3vxcaEShWctT1PHG0zWYNVY1F6V7crIzf
gSv0kGXXgDGvw1WskuegN/v+h0W5F6jS7CR+wKRX50sltQbdZLv+prVJvkMaxbUu
Ha7guMS/lb8H26XoEWkkWmrBtf4EdYyLjN5z+QcoI2gDhqXfCOpQq28rK2mq1T7U
2P+iua6c97IMVCugXcfN8GvUtVkNTsezcfPrtGUX1HFVz2Aa59unRrKmmjyK11Wa
yrzPUegxgVEXiCJFH52St3zn+fz9+uJ3cKV8ruWvziB5nCR7+n1TJlU0alWzxgvr
ekfBR4/XrsWayS1mjXiumFfypz6F+n2Sg1t26W8RcoA/o/WIAnU2u2KC3E0sSzcg
Cgd2jmFaTJD9FSdYfeQFGcgKIUbPDLq6K2cK7Lp7ikGxDrd2T0dy/HLKyJFeyUb5
wrosPXO3745QrfY6DdAKmIBzpdDOBmLubfQMCMEysNOpgvNA2qYfOAsUNHSk2OTp
HeLLU2ShcNIlwXyckNLYLPiWBcBi5tNwDA2Rignp36NGh2BfoCQ0cGmsrkPmXVR1
v165iEKXE8DHa8E/P4PZVTGyQmQn/qNWX035QqhZb3YIhry4EyreiA/XFAB4jvGg
lAw8VHHKv+A24ABI7KdYPqY4Nn3FK14L1JE4McKqG8Y4HLewnooer1bPXo0fIiKv
5qd8rLCQY+bl4RVmMW3/kw4IWRsPWxsN2i8pVrLzt7EjQOFRj2ZCO3u9yxCMmVz3
546Fcbs7T5JmhO3a1Zx8U0UJGrjmB+fWo40Am8EjJABopM9xwnBo98tNh4oSJUbm
Pp0mJML0qbUHObFHbkCjZx67WjVtgZmlbnCxoSj5tgejcCPnWgsw4Gp+peFgU32e
DYp7+6pv9cJ4cdRF+bodEDS62VezvUy8ddejoPgv2LwPwnG9A+XEBiwNnteWCsNc
V+SurZ1LYH+GoTZV2kvfEqpje6pg3ZGU071DoAOAoNghYK5Oz4HuAm1AMYZeqypb
aXBj1t0hWzdoKKcGOys7pesnpC3W9qblGp5k5XolQawFcvVJeQR42IyVD88lkHY+
QsoAMc8HI1uTDjM99/8REQLjrRAT9ym6C73EZdB4gUabKD/FqHiNvfXXiKekUtk2
k+r8hBx2n8Jo+B3TKTFXpPsbNQNucy8Jal+73S2VxZ+xPNLCnh/WoBqm8uGdonvp
HaY4/+lSUDHPnOXU4LsHQMy9Kiv0r0SzDr4Yu0LmVAgbaEslJEBwYRo83i76VmES
B73j5Nd18gUp5PD3d6mZ3b9+NwN3nFtjfdo1JLYa8JYpsy9nlEl/rTTbIokvLX5F
l901wH3AIYz6hc1U0+9NVD9avYCsvRAMqpw92Xbsj9Arq0T3rhbLRWYcVoFiRiOA
XeLGFCOQM7jbIdPfUa7Ut9PMjcZDtzWs363pBOMqtBVjYnqgSLbe5dpwBlb06xYn
wkvYfPXqNUfTze/qaXwzl2ElfPMRlhyZvjOPzvs4L1nqrej7p+81SdSNaEtWjfva
yKTD11LWwLETmITbUiwkaj9pVCSQ+LMbTER5w+KoTe3z+aF9momD4XC6eCN3H6mA
P9QPP7KKoTMHvzUlmJSxRMFoMyc3cTmsZAG4+pBJfTuL8t6t/+yqyBAlocMuNAKG
ECO00DcUsDs7FIPeNXAhGOcNU4H2AWbDpIHqNE0xPo020DhVYkSivnOh1UeSNXjP
85NIWyiyMSMuwG0J04dyDFDsm7CNzLV/cwFqnwWGjMUdFcTefKMhVuccNLN4xNXi
3TmnZTGdqeEcZr4MRa3sh/irsQiWZxzLVVo3e5JD/ZPlZRqppcLPLjtrWX5F0W5H
7Z9JfurPYfCrMPgd2n1Urr25QLWkBXZg0vF7BKUI6yrIExDorJtZgAIzt8c/nYpM
dEhTAqqKVhbSDrdP1RZjMrgRjPLEA6ljS4BddVSr9yIOrkL7s0CMv4IZuYLYCByK
/zDQbd1BDYddVCR6QHsvqI6BcCAWD5AdnNXqBdQljk3944NTyiXRnuEdB34yPJdt
JQTZj0tHQyzHyAKrT7tVyku7x1ssOGVganyuQTytBG04dR5HXaadvLNC77qq2gl5
GZNrNCpTMbDrXpwzwG6qVwsnCpYRJEpvjsl8QZzQm7G3qQ2ts1Cw2OZD4f5bnZJc
VjIY2+O/kq9QmsGZrHdcWSLMDFSVfvcAord+aUwaQXtC03GsBZsZy93/G8CrTiCE
C0WWC2THJGDPMEnCqYzQqqwAgmB/D+lCA4eYVD0vtc8g2PddLitc96qoBAjQ4G48
Qi14lFuQpB8N3Yg9gpHJqOZKfws2OfMC/KuQkeT/CCkhX7Eu75PNJAuhXPPtrMwV
6FFH+OstKTBJ+RBzk1wT9RrMZs2SzaPkuNbJmffEsHtnFSCxpsqgXgrdjtmvqUVG
vy0uGvqOgX+bolVGwbdijylHFnuNFgstGCSOHb7m1bkUNBvAQUrobe/+Cc+KpJYF
KZY6NXYmPyqnUnxfqPF3OJapoMwpWui/wocDDFm0wciZekXgqMBtqXxYhcDwYedn
DuVzTSzq8xa0/TOtWuz+xCe1LtgemkpqVA0q2JrQZkqeGosjCjP4YU9oA6ruqF32
Gfr5a3143s7fzM97ZI1wyKbeyoSkXvmNfY37RUyqqFdANR4v4s1728HtgFz53LlM
MrdhDu4PJE1+zCfuvwsaoLgq42v4abnoxnQ2fwm9KPOjYkYYaBgAGGbbfohh02lC
la2Xj6j5oo3PmlkNZxYAloz04m9IR4vBiQ7XPELgQpO1fxuMgBVMQ+QfVWUL/jKa
Vac0JaKxG3XKsml93I6otRuaDr7DrwVHqYCDITaAXrjy05GFH727jpIR3Hu17wi+
9CkY4GAVX8KJwVP5El9TRp98LszKuzLKQtWy8ez+j0BL/aULlqEuOsweN53yrG8i
SHge36qMj4iaX+I4gT1+EFQxbETAK63d12fBXI1eLXSaCsxi+rRLWx5ckb9jVpoM
YXxobggbmb6Yj9ytvU//Gz7LlDnLxPvAdGMp9rIFkyuF2VvDYBMO7hh3P0CB3SR8
jSTX6Ip/5Rw6LfjMg0MciusVhh/Hw63YmW1pOvadaj2lGigXx3nsglgCgI6dJg9F
`protect END_PROTECTED
