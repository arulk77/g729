`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKIe8bN5b7KBjpMQ148b/djsDMKx0eQRqI+qlh8SE7w1
RCnmcJNOh326W6x8NXL96U/EI/f/6sllsjsi5YDYu+S7nHxSECn/ftB1LcVhotvb
5QkbxTZoNEOwZ2TYNOaPHZCLuJDEaMGR7Ixa/rDPWAqkuLW7z0v9y6dIqZGJpwI6
mzTY/Lr/M3FlbGHyQ7kleBEr7N8RrCRW3K3ONuBEgEPmhQnQL+HnaPW3d/rMgj5F
KKT5ZBy5JIfVRxLtiyAlz2kXRUZ+jmhyHh/0WZqZ8tUaQqDWI+GEbJWYHIGJKRqX
K0TGhIDm3erINLK+brgR8mK5yrVejpKQTW3YQXV+e+ufqGLkdKiLteYCbYR+Q4KD
1lGIGpjxzie2JgCe23GjaKnsMHIsEgSmv+BzgopvUzyn9BwZ+16UtueuKJT3jj3V
UQH4QZjX3vtS7CiJqJTpnGQKdYlkNYH6aA3DMuqLCXeummB17rdRHioXBTV9HWYC
RDzar1+ihfu5xjeERux6nh5HiTZ9CFKI1HGs++YWpGG0kYiH/FwR8kIXexNgYoN0
X6nIr5D9hyaJhUJK25XOC/mPxGUEmEkA5lpqr1T63ohCAaGnj7MTgRIrTAY0cY2f
frpcXai3eqin781zLj9puLUQD86fCTHxXUtdZF/qX6uz2l+IXaqj2d7OQWMNJ5HT
`protect END_PROTECTED
