`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wh3MdWUqLK2772IY1zkvGZHQwfAsONiCswbw1mV2U67
L3z5s5OaReDvOKfC6vXyLW5ZbMVPVec5kSvkSDYoskXqjneF6nn7mgs83Sjf9J3P
vVysFvl51i29Gd594HWyOATSSrIhJ5rNvzXCii0WP/tKgJIZ2ZYyFxoO7MhpRJCo
9TGqNEq2W9cjA8bfOpb4HEkeLlonpfOksclXtk+A0EQ6bEnwHWTyps1/Uo5Mg7Rw
TFC4TwOWuvWTqDMqCUl+5l3KLZgmTHmYBjFOXBidjLV0sYJNSt361p1EnakpF9fO
yS3SNeoZ2IZ8GgjGxlsVUCV2EhA9V7TxLEUAJNQxRjsFWUFOUrEtqnBM935XyMsz
162XscDhOdE5YpBO+AYi5A==
`protect END_PROTECTED
