`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEgFP02SXEsWiwGovFxqGfyMMpX2LF6GonHI566wmlrc
sBABm+FoSKz626Q/mXflqiOTbHKGWheTnXSrdyho7MRxEJoKawBHs1nqRXpG/WGg
VCpGgozzvYZ7YMwJnULo5Pe7PhEswm/VGVHRFEhtnQZy0La3JX9M/5bidSY4RrEN
ou5ffrjA/PrNP0WyAOknc43nM6NXqgp4KqyWLq636iY=
`protect END_PROTECTED
