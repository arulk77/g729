`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHY1IOT0w3Um1LH+HS97wg4sfY4zYNIAiaza5i/EqEaE
QTy62BHBp4OxapK78K6vDyrBMo+hN9Oi9eRdr7ZnX1YFCUDXJFfOrwBwQbR6o2L4
RC1lLEkYJbTEeX9OxGXFtv4qSGEmqF6nte4eJ4pM6GBg1aSJsbnBoljrDXUTKUMs
GIqVPVEqeosbr/56v4BlmQGqBZeJXU/BWN4RJHrzXsZQg63cKSv+mM0DUbawXWTR
WVJHr0kZDSVpHJITPRP/MjaVazx98Kv+OdOVR/Imcs4+GS4+pTTzDtj8KZdcolTW
5NLVScXOD8TJrzRHKlJLlEL2S1Zyh+eABoxo3DJWZLHXFP1Ngx8/LGEdSPMDmkqQ
ehmMrgribDpspL4j1HJoLl8kdddhdET7DT6MdyBpzNVMXagSZQjLouUyCHYTtOoA
09kjnni8IehxAS/NSMg3brroXhWnrSA34TRqgX74X3E=
`protect END_PROTECTED
