`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aT7wtzvHCxHEkqOBK2tRkeEu3yfi9G447DxOAKi4cPWc
TcYEvHa7KxVJwfzRzoCv9J+/+wxclM9yBjNE23oxvxcl/RQ2xCKqqvvSSF10b9pD
v50Zp0mhB2PbD+9b0GgvLAWDZrOuiEsUm/GhjURK+YyY3LcGQ6YlolRmZw7dkAl8
as3Ki7bx7t6awFJetYUkmgzbkmercgU9N0DTvhqKmZg7ZthW2Qpmh38NrY8YfZ+h
bJGJlX5UXweiqUyD8S0zuEA4jenVM8QIWWBaXc9gfp4FTd1f3Y/NAhB1K8LWcBAD
fFaJjII+2/60zVXMOJQ+PPpu9vBmuGD3ecyULm8nY+25SF9H3apqm2GLdXFIAus7
jOx2Se5lVK9W56cUcUBvhyg52tXUWPSEFZVHs5BATtRzESs6/l7D/PukuYVXyF3q
95XopGYc29QTC15HdORqwMelryt5wuMHlrCIC0LP/33r2tY1eX26QGlBcSrLt4jw
nLSYDpq6Z2DN54OdXRTu+phK0V9yrZS+X74VTFc7xqoUrCQ4qigB1O1P7ztBHYVh
dbEOvPl0VTss1scmFhZas5WWhpFpKg22XEddUcZMWdfMwbOhjtQH0GHX/J5ixeXb
kV8Ov8CN1Zxqs++wdSjeiH5EelXNAWg3xSUtR0yTlQ9sJ+ECzFYPnrhzGIcbhQVm
ALIYpjGC+GpL5jjbO0njYb7OuFy8XfAT7dVUFR5QnZtTVK2NWIdhawhKpaFFY60/
iMPG6g/qdKFm5Zdjf0NisNDLL6n/V4VR5iH1S8PKN8jNIXrXJ5AZJsugpDVo+Ntj
V94SqEhWMT0fyGWQ5d9GxEFiq25WZQ51HdA50qBSHt6KOQuOIzXtn67FxW+Fc6yC
VRC7JTwlIFp2KHnzH9VSsULOCcZgNs8StFggp1HIm5leSTeXIisTo2Oax9H0nUh5
mf2AYdTITJy/aZwFvsqiH7BlFGsuzPQGA3ygZFIjLiyEtdE6aLw+ZAR1BhotV3TN
B+qlTyQ35wf2HAT0Az+iroGN0O/h/bianbFuKueVIwQtZUQWKujzAbiNFp6wWzCy
z84BZWX0BlhTl1DeT3hFcbGS7/pQzrckGXWG4T5moc1XK1aZhsxLq2Wg9UxUGZcp
T3PFwqLD95LO/0OgijSDNU4KE10HBoimZa2RH/HrZg2bVjuQgSxP5JwnEVOR7m8s
v9NDe/IM0pW2BVclmR/1ReC5GJq3OO+bYBaDDu5cfJ9nyqCibEwWs6melh1agLkn
MJBMW98qBueNe1eTcirnajZ8cJD7dkpb4uBWCinCt2dpGm8xWKSqnO2BKr7BExB/
Sj8se5LcqWr1ME85TCBbmvmqTN7VAZr3VPWOkSddY9ab4+XGzM2pQqbb7zYCEqxU
3S8Zob/wyq4cN6+8GcQuojtLgNjkdeWum7d0dnM5dmge8UjJMvDHTHp88prE7UNr
urZSrT540gXas0LjssGrY+y9fM1hdBx/In1psNGsiXxhdqaE0rPJaRmH3JSUj0VI
2C6Ex/Q1cbzX6MWqVib7ERGB1d4yxpWLTGCw7+R/CVp9oqgCQ0vQyvelSb3bHhXW
ievNGwMig9YWbWQDBN6o085JVfmkLi/U4IpOYb/YNP0tVg+hB+oyav1iAg93eSCz
UkEPL9YofJNkyWAKsiaNEORnxJB95/+Rq5DKZ1ABclKmAnLouHsIJvAOnXEP1v6d
/HFSrabc/RAsCF0PWLQmv7joYOLZtK/jP6tKoilycJHmDAfNDM2SgZ+oCblejZxw
3Easvyq5nMi2hximuTqqPaQs9kHICmJPGJccW9p7EChFEPFtggPavaxP2SPkvlDM
dmjmAH4Ry27GfAtqvwAdICVIP0zGoEz/S1a+JVbtU8lUezai4CtOaMO5q9Do+pTF
CX5AFYakN8cc2ckCZqF4/zVIU/TtUOmJx1S/+b+cThRd7cNynmkCIrsINqCa6/F9
PSH0r0QEEOvcRTkCgYS47oPq/PPnoX2CXxUuXHxr/8vxo9PvBr4n6wr+T7OCNvJS
5fgH5+9I/SaihL8hw9h/1chO2PGWhzlGLjho7oJLnqnOpqXKksyEFJvU26fZiWXA
UL6YidFgwWxQusIMUxD/atCkB8NZU+x7jbM7jvGYDZOZl9xwyoscwB6ot9C/JdGr
P0uDol9o24BBqGhzmNZuO0OoOlIunKAMBeKXQ77nyqDs6lEV31jnVBqeCZrCo4gi
WShXFkYM7iBL3SZSu6goEqTqVeCkOi7iRr8XKA1qHLuOetknxJ1aHrwpRKvQ2/DI
oBjkiVChljn0AGt2PHoUNMRfZyyBXXVIJaeLknYJPINlI+iL+/58JdYZ2O08CaHx
LGNP75AZjMhlK5vq6wffQCJewrE2QBw5GGy+KojWNzoEAsS0tPM+1L7m3OrtH4Sc
N/z/EfNUBZSfTu50rz09Zc5oR8g7G2zo5HtUvthVmSJofH8wc4hqPi+MN5w54V8B
qoSFnuiJSDzowsxRLvD1za/yTQyd7OCgxljlKK/kaWM/7Sx3aA3GCX2Zqos1hi/E
5c2o9jxQidgzBFzzz+EaA7kFnGwRqV4akkjaVc6VZvXJytYZA6/iArrJonuvCw6r
Lx5eZ7ZJ6EdI8r/2konfSDzMAy3vl459K4AdW9SXZhINbG56zQEPDMOWJkGCGuWB
7EmjsdKtPMpp9bEsaC1m2ts42gARIRbezqy5flXVRLdCzYyfQ2NC7lW5vMrk9JtQ
57W+29f55QdSJL5fNOu1PVvCkFYF1HaCoF7Sf+76BdNUtiO7Ibn7kDDXAu1H0WxW
cPrFCgcm07KpfYrBzzoN4R3Y18vepQ+/0kHBRFDTgu/OGsIPPQNw8CIxr1xle/oQ
3eLeIubvEnF1L7stHbJz6SDmKUon6XPhwG8ZS0RUVFK/PAPlmIr/6E/LH4+II2Td
swZFkKleeC3C9uAfShtn672KD9o470K5wi4YvxoGmTRs+JuW19dGzBSzyXuc3s3B
ieirFMBA33PcGAuZffb4SwzdN4cc/CEAc7U/BIT5TZUAHiFHSBqwO3lDggOqUbFP
aU9bkA5bOvrIzPF7TKNjKZDuV3hcbYIDF1ID6Pxik9J2BkQyVkiGYmsfdjpszOEx
2gUVMG75ZaamS1bkY+8ZLf/T8X60u4l9Lc2izcNhKKqwsB/v16ypHsCITPP+MG7H
vPU5wzMiOGe/oDEGOG62s/MCIAOQH7OpnrQQXRdQKrCnzSe2sW7YXpWNjfJRZF6e
fXyY7Zp1ZKw+wjIo3qBGL+BmhjOk7HFCc3xhI8zW7ggFyRUcVu/M8Ljtbw03yKKe
JmPEOlFzFA27N4UV+UmgbMvsVdT5K6PX/ll5bA0NMtWeYbHQ6FNY7H3z7BinbkA6
GlMODIOQkVyGeqSxneby1ZdtDmZioq3rxZPOkGJaJWRHlEQtSWN0Mn6mq3+3YJvb
vWxdK8vBWBznNgE057CLhU46E6REw8mYC7l1J+7CZq0j78TlC936cxzHDFcTAw4P
NgReSJ1HbgZm/hPFe9JwZ59OgEXvHzW9VJpXV24PCcDgTPx+Ktv+S/fJ2v3XDzAk
i9fu5folUvQvLosxaN+BEJOusOEXhMx8FvpuVCSXLTz+ErMpL/RjjyCzx7RCAiR3
MtFmBrpRk+h8dFZylXhxRL58Vs8Pse0Dduw7+rVBoPR88vWgSuWZG8If6LvrIqgq
EU+nwgkxzPCXBXOnOgXHf3TqdBRi0e4DzJqukWdFs7w1C/5FfG7seUrCpErbEIPn
ya8wtC3o8djixj3d3/wV166lOm8pCLwbJ90reDc6OlTsE7HackcXKIDeASww3z5O
xhJG2FOyhJjzRNwSPxC8nmK7Y8n57KVYAnvFLMnGtK0V8Ke5vicwD6yumMHyG7f+
T76MFi0hmXzJlbWN46HvlMsOnNj/qh0vG/RYnirpOX7KrFlvzm+KKU7rmQ/3N/DV
jJ43qZojUseRDSTwaUSl3UZ2vOkMpPwfaR6MUBQh2ZPm6f96+FsnJM96sqwZnmGo
RyjVQqQHJk3uWLwxETjcrU1KRj/ykvqi/695m4s0xqaXM24eFyEC2tan7yQGESPD
R3BL8SYDUnsCYbOOo4XJbTVQusihvYXeBQk1Mefr3Yb53fwO7RHUNwjyWD8lCSwV
+npLKoVmL/Xp8Mcg5iTdieLSuvjqZ6TMjktznvDOvePHDfE0eb0CysVEwteNceBC
gKYNTB5E0VaxnLMPlLFMEhJXk0yuFUjmXI4ETh9Br8iY8Q2fLUyuYvgj9YGW0KlW
sufRC8P+JCu4BfneQABZfALvRZ+mVjtklyhVLc8l2G5xO+DYF9Cp0IZ8kLkhZSdF
XGgwfkD36Z5WO1wSOla3G2gUPT2mNyRbd9+H8Yni2mV94qOMEUCRBNQPCw2/vEOy
H4qWndT5FF6YGvOnz8eayO27Mf2yJuPF2APMxCJm1lP+H01gcK8CvYdysWd2UU9t
ePUu0iUF/FaRqelMjZyS+JBwKrFwNKlcJEDkrMjRwn5n5DbK5QBXVIhTwlEyjhvA
8eeHGWD2QW1+vi6HYYr6aA4EMdH19hfrtXCfzy5hsxRqsTo+noLWeeigLGAO4Lsz
KPBF5M4zJB8nDzN55RjT3E9bIUJwOTANCS3g8kvlDgUf6KiSJ9iwORJTUMR0V/ub
qMPZGiyzoq6fFBaHD3n3NnLGPg7ucJ0qafr/uzlIRCOsP9fcBJDJoANBIO1HWRCE
0yVA03dQQbcVD1ZxtzK5cYV7qWpid5yti4sl3+foMd2Y5hva2c89AA09k/Nlnmf/
JZUu8Z28ZzvM85pV0yZDvOMOHApRd840mKLWY3B8nRdF7HRP/6vMbrvsgsvlcsF3
5jqMoJYc1Md8mr/0GRlI+xs8JEOdtEeRY+9imAZyTz8v1H7pexEEcwGgDHiBnNXJ
YWh58sH7KxoUQKOI3G/JNFKPd9BQ2KO7I7WrcEhrYIWPAAluXsxhUDsjRZAi/zc1
329gRXUzkpxAf7MQVkllR57O2bX0Jh7z7ldmqQC+bxsWR6ntWZbat1MPStcgqlTm
GNop0BsnDUnGvyriZ2b++Z4m98CuUcyH/jtjvmeSrB68RzrEP1APYiP1w1xZpLOs
LxqecOUZd1rQNa7dkATZ4Va0JJD3Vo+3ulgWAqmsIIl98otuTnCzi6F1gg6JGBKE
Su0QZmLcCKT3PFmaW/ilmYtlP/1UqwkEul2lrMwnkPEc5yz9biEflrOlt7C0uEi7
ukGH47DrTuHJ26s7FtOfxvdonG/ZLyYc19yTDxs+3QUz995RGCdkBaU0p6dYmwMk
0+w4n2Q3a2j70s8i9y9S6LkPHMf/XTQdOa75Sh7n7SAQDHFL5BnZvOiFDGuuutfZ
W0TXqyQ6t/YiuuvaS+tMswPGDaoqc1+I+2QWUbXbeq5TFyZ/aclmNPzVYCDAvi+l
NMJtxuiLOm0kbNPvl0JZpKHvAoA3+c2j4kriqa9kxju3lgTbHchmGSx+TVV0Vcn8
1hyz0jjwx4K/6kRq2u2lge37UEj4X3se+Bah0oSr9TSXFhQSlMPb6aVUSBblLGZI
nKIbSKapgGCNsQAIHjNaR9dYY6Fy2/aHbMtn7BB30p+R6FbHfbX10xtzN5NNwIYP
63+INrYDwVgLQJdFU+Nu6jOZmH3dDYsHlvIipBaJ/AnwIvMCkfydyQLhC6CFrOum
eTcFW2Ke3pZEAKmdw9tzHx2HwIyBwpztvsqhdnZKFFRfFYJtCTescctw9ldrmU3d
SOY8aaULyEOVPlPJzvoQjY9252m7/yFXW9XGHumfwCeq27hpkTq19P85EpfGhplV
KU0lWwkld1185oEibhnZTGnkmKr4YCaXdx4pfpXpeFaoLOQsvwGXuNAN8lR3f+PY
F1S80up0t760S8Dj3Jb02g9sl4Hz/lI2BjLJTdcO3UOD4FrNulJ4s4G0Bx64wftx
2UCUbacKTQBelFZz/joarVRJM6C+sxHCCf5TUY4MX4/Ko5vpqnlcm7POpyRt4BYU
gnQXwnq/UWCSWIqK0lendFn1NbPPq8aHIYT0P1Y7bw7nHgvUpAb4EqNjxhYhxsIl
RTV9dw/NZ8imT6Ecf3L2ajIxVTwY5PyftsaIDuIvAt+JbkLgO0NWxUKwybzoMVNq
hBl9IavSTX8nZBhREiufi3nvRcg7qwnU29qIVcaOpCTAksjU7jeN7Xd4EJyDrVqH
xng8XsdqvfD4S+LjuGyAjCfnTyGpP8mrEK0HTakxlfHFrMDXLqMOS6ZkFllySf5k
tq5w/KeUReOqo+dGCoRNFl+0CNR6ZMKESFAPIcbODp0BrbdfUH9L/IrIRmP5bG83
we6YU0+WYtD6rKYsUXPM9NBH/WLGLnraax7ZlwvJ5smPSU4Cw44kqusNgUbPEst0
L1xWYYjV2yga8M90D7e3KmXI+Ek4jXg6mK2D7eRn/2NyUb0lsrosXjzZXoPQYP8j
Ezcv8ISZsE+pDps7GH3tto+eSnE4E/ZP6kCZPrLEuwT2EYKXTjU+uwKMOradtNBV
JUiS1jMy3JEE68d4Z7fOvb2tQrudfOKcdCpDiHgwivis4j67u9jj26BLBwIflaql
fm+Tkqe86Bky4XAPeKnqFRCrYc/ufnoROr470NibaDepcD0JaAWj0mMlMTuZKfpz
0KA3ofRMA6ZZwn7UzCQyptY42r9fUR7GJp518K6xqFjpKgGoq3SNxY0+af4ZFBfD
oj/XUj52VDKH1AKjzeqgFhgNHKL6VeVJ9zW5g2zThKZfyKL5MeamVlXWUrQ6jIeb
o+Htbtvws6mEzUl9wDtEQeyKJoOYb7mq2g+GpaB8MB8YPmwJzUwIr7uWQ8JOSAHo
AIMCKwyVGIPbSoxvU+XCPa8eFLJVwzvtLVfGJfDzPB6orFu/C/a7sa1ln/uPayK8
6bMqsH8nFVj/HlBpqwDSc6um3EtG90tK6VwWGT6/yycTzmHAoRJ6nYaRaShYrP0H
8FCNlRLB9EPXQoENlfVDy72zAWCYVSKvSQS3Y2Xu7TezadUZbXzB3KybrkOlq4nc
Hdu/TFKZ58cuKqGOaXDlvaIXSl8bcuCJGrTf2fzZsolLXyPbDEFOlqfG1UuFhLpt
wuIm5lPXbzEY9gpzwepgZdQSusJvgGZ5Si0r00XmhLV4C5b8tvjy5XT5Z+/N3Yz+
eTxYh1JlQTFTHwjXDpVYni4ORGM9Ep13c8ndCVuvvl6QzX9eauHTv8tZAPUvQrPG
eO/4vwRV4KdvnjZ8vYQWKcTcejSID9KIkjtkbDTEOjnZuU41WoS3iDbEWLghA3w+
E9rgPDONXVpIwpXb2XAz0zNb1CaOOUpNELEblX1+K78ngLg1i1pgQBgb0EqfIIkL
ESPQnF0+tKM5dNqNyl6zlhcDvEG0XpVBKtDk8bRp9jxHq7pUqOXr2eu2TroFbCX1
JnT8EYviAqac6AZYNxtvNFBKwT+5tSnW5xGnDeC64YSDkji0oVwU3MqdXrET/pOy
AA56gOIRvijs3JGksV0CkELjAnzIfUcbX79iTw8GLbLj7lR3x0qNzCu2I/BPhO7F
RZNdcWNF576dFmbJIn+lEJcppCMsFsod907gd3E8QFJ4YnfTpiYJBC2M7Jsl6O/A
U4UeIdUGIF10JyR7omjEdrqxUIfTDyeIjayMqBC0TsDGmOTYZUKJ3wDvLXlLjHo2
E/MLkT9Sp3O/2ryi29qIixOAxYeK2qyp1pDO8xhobG0+PlnIlnWOo7n1i5HUs90x
14z8HxNHfDP6VevMAVvx7sNgYpkzRbXu5SBxP3Ct9GngQhjndn2UwBLPHkMBULk/
EfuRu9ywr6FjglJiO5c0+SoY8XYnLsqle9RldtE/T3Do4uW8eefVSjbQm5CiwOi+
RWl6KgIWDMlPeUNPRJNNpd61+USBlm+PqsRO8CqRl7n6mwKnOzNdr08nqVtbwwdd
tDdsW8Duasg03F6AY+kzvw0JddIiCT3dHDOv+1LqXFx7oiOZKfQVm95zQx+m1cLe
IiitqmXCqYP0VTqsu42tQujtV0o4KmBHsreO1EMGzvVAd8l5M22nW/1JiI8q3pGB
VARISuQVDaWZV4GDT2ic9yhhmHPJGIKoJUv49drn8ffOibgQN0oqwZ+xJjRsihbb
sBAR+ezAS6rEB4qYLPIPzBrMWXNjVPFjKiSFpDdnqTzJMD1W3EBNimvhB3oZVgEO
Yu+T/9SqggV7c9J94Zg1BXAgh0FZyO8xRUxo+5c84DQBIlahIXHxRA06HfuyisqI
z1oZK4bJURzXpviteP/jq95jkxA9kKzFw5iYtLHbbGs4NQCd2KJZPEMmuBnRvkQO
Pucc511BqkiiNn9bJk9JCGeF307pKIiXyh9S/R/n8v0l1OiJikDY8kDmCE9P0EPk
S+aUxQ4xOM9Wbfc6dd1bVbcwndrE3UO2bb6u3ovGmQHqdKJACE6X56QEmzUuJPTJ
MmTwQJBkHutzByusXNHfyoZMFlVk9WYFP0YPJurpMEazjwwb9ev7v0YMvVAtMux+
5y7SViTLEC6fOnkFyAiFW8qDaP8vHGkaq4l3lA5i6xJ973lMUdQiCtcErA031MUL
RGUMKwF2+DN/hvUXLtbceUOSYNjsD+THDM0epY2PSgywcnJUMzjhWm2yRb4m4Idm
eV8vqOaUYJWqls2zGWNI/370Xq6m9sjMg6RFQeXmJwX7F/8H+K6Glm0JbCI5eNUV
uCXqHUC8EPGn3jUweGATr7StcEMXeO1NSMvd1P1hItfr9GoBSym6cDS7gFM/uoCO
AiVDPddNWywd635aFI31GtE4C6KOOpZC09wLMQk7sL17VTUZFd5QktWpIzWTx0ET
7zA5kB5ABmgXtXmiYfCN8172y9A4fYHOEMZXXe/wXWwGvwq6K7Ex8bQ2hNBdL2mJ
SN/Gg8pSAcdfx0XON50/fIXq5WaBSee5v5L5mjhUSVx3UGsAW5K/KDnEJjutFCfl
GYNVkmPu+cShoZ9vMEdfCKjmLEtrVkCQAgUSQilpk83XnKv6FnsxR20ztMF6euAU
y5AYcKboL8Pz1/WsQoUbj4cEH29nCYQkCm7Fvb/y68qJZ8zCJ+xce/uO2JEHjclf
ol/SHehBkYeEAaskg/CkNICm3ivHRlGyL+YrMNPkybInvxQcKAANNEbPcv3Xp9Ao
bsU5JTE0QCpMCd7jZIAFTv96njt9ndpyO8tYUuojQwbKmJYzw9ZbIbN3N8So/6iS
xQfZLXzN8Ve1K18Gp8vyB8ZSWPFryAzY8Ut0pmPkIdR2LwdO7L8e9EPUAvN/QEfN
kl945eDCaLg/+x5X5n84GzZLEOI8NGY82bONaMxD+05Vorp/Ne9s3sFZ4Kxz93Dv
JdKw6nTi6/TFO8XdxMuYNXc6NcC8QH+/gHQttsiomIwNLFCDJma0YutMgP7gKowx
Iy/4yx39/SmhCFNEsYOqUB4X4poET5QKBcIJ4msEDdoo4UwJS4fbSQAjDDvIyVAk
KOiI+yNrq5Bd5QUYDg+siJ4rJXnx3K6OY/LJnvPTHfS6YdKPtmwLsdCmIA/tPbLc
Tc9r0z/8W+Z/dnEwnTE18bKb2EYmK9+7kEeUJRQY0FOv7lEyYpwgl6wvnuitjgYy
pbta09WW2P2fBZ0W9vbkV7yx1Vrf37+QaUtYTopYVM5D3tb5aqbXCmVe/qiakL1o
JkEzDA23VSKQpP8p/Qti9Xv3m6GsAIfiOMNRexHAonZsWB+BXRGdi/ByPcp1im8v
aAVDfpa9NrxuqFZ+WUOwYknW6st9V7iMvmoXzZD8X5A6PgfiTDjD3oSAuKIAK6+J
lPhs3ToCL5hrhE1uJxkeP8LaPAeKm53jjuXt30Gucjenufj8vU5oI4ScCcktpPIT
a5KWikaESr82hHcj7xSOkxDtYqTGkKWr2yKp8ubMTK0htDBr/rRRxipoEaVh/VdZ
i+CNQVqS67E4YRt7snL+Kf9/zXMNeGLuLYMln7JPxBD21sXR6vJQ61OE/RuGTa8d
gGHDI4ccpiVm545tfMTVIlzxsc+Jq+VJEgF9V5og109MvT+3R+Dyt5o+cj4gV7Hl
VK3x0WkB8iC01kVT0d0IxC1V4yKZcuKMtZAVJzkT6YnAez13H3Hwr26lnthEmHGV
QH3aUmPPE5EOs+ziOeSmVgvo9J3U4JHI1rWeLO/OP1BI1IyVYbR4QbbSosopRP5a
+9U2IGhDiqzU1hnIE9T3PP9Q+q6tomPFj5mcObRVDYgW0p1bIQPtwLqLdnbvzUCH
xR4kVVFf0V1aY0agvNiMHnHvPVB46uFhocUNwvhpkE//bEpC4d7FBNW6wNIO+mOh
MvedbDqJSzjBlsbaRXqkC/TZCEQyTTu6CAeD3z4/Qy1nHFlm828rLklOu8XrzPrk
06+6k9HrHzR9aSbXlPmXveRyuMVY0xTLG9uzNPqxKBxGznhZG9Lq3JhIh8Ntzvon
rUvu9wZIraMMu0zXpoi9O3G7NsqwN+2DxVs4wZHs28w90hDvdGcOY8Zos4yjLSJI
l3yiewC3nzI0BuwXFABFKqtbkCGnZB8DwpzjqpRQ66X4SbZm7qPTCT5RovjNLJGe
/ONaAyQaXXjTRtjWnTVVq1/hxK8xznyfSzopWbyKldV8XAipNB0KXTKQJyyOgS2n
Jhhsa/5wuuiDZyC5RYwjPf/ivmISvDG6DkfQtptHJpmN5TfpMV7fzrHT0cpY1NHR
Rsc1WOYC0uOrkJ3pgV34n1PFyU0FfnfijndvyBa4hC+L9SMJwZ/f6YisScjQEfaz
C0R/jf8W/EEnmzhYYMg5I/nkBTZdgvr71jIFBQS6YZZRJqm7s1zDYSwUQgLO9HoI
TDg0rydBcKGabGxJjROVeh6ohjgB4A+8mgmAZ6Qsb/+hhxXufRz6IbLq8qwW+TCf
7B90k2v1A/TQtpLfxne7ND4sWXGGY1OiyRkN2nId4UAyTeYTFl2sQXOjmmbtWefK
oNYZhA2uvlEZH4tdGZLT9W5Or+y2S3RRqq+PG/gYZsaf3MlGYdiKPDnZ14qG44yq
sIkrzUxDTWnkUT371nJyxD93gPKX7d61yTotIGnla9JQhwC2HgyLfbdoz4jJKB9g
EVKC0w/2+GvmQihQXiW+hcoGObGLx5R03X5m9XmH4amLssImBGmU0+a11bI8oTsb
8IWQjNtkpvyg8DEN7C5Bq9TWUvigtSkGWCs+HV0rqk0R9QZsupUWJbELiVXpMr7O
p5HYLVt8Etx1kzGt/LHYEWDo8b2/RI/GhHRFoLj2ZS2PosFtWT5h0cyqvzSGEjAu
L6NCO3xZ8oSrZJfzrp1JGK9s/5W7Zwo1WvHO0Q9Cb3qZZlqHXhuUwepEv+ezK2QA
fjC/Hx2c2GVHk4yiOA6nyPoTz25KCC2f30gzgA+nqayRRLKmVeqiTeGG5IiTf8HY
URCMdBIWKJbrf8awslUQwyoOjFysX1DYm1glO8pWFJwqrfhXuSoKYYpSOkCJrFaN
Iz8Fxk+s7n6Ok4fBkOQfNjQ2k1FDEJz/9JquRIbB5PsRAMoBBirtnby5yvwK5m+b
N7tTxR5o6TSIRmO8xHZ3l+wCzNv2T/oE8M2a9dmGJLrF/GW3K1cyFKQUV6ebuirw
aByKX3th9LHrc68hFv14bSvdcsmb92fs/IEyKZkHga2D13J7xUx3o613IL7SH70I
4LSNdKmkZMQnYjt3VXuMA/3wR3dwD7XzJ8oke2RbdwoMCapg+Y8c9ygn6gAaf1CG
v+SpdeLPZYs++YD43GdG4VKnHNThhcBmXjQVp8KWgLcAAgY5pdAI9ho989Uageoh
HBm4bdnPrYqns2+aFFfsnLDiDHPWZgJn1XRwGs0CGsUmN7YsewqXt0irw64fTYZ3
NzZ1jC0NpgSXw1bfy2KnE/NjQ7enLKdiD6hzWmnsAU4M7E8HlDlJKknQ0wmiKBfE
EUQYWokmebBlVOKgj2MBCr24r7jgR6nNI+adWVo6sIIjwLULEHIZLmvm98mHRTFc
vfloApAxSDyi7ynBduuQwVrFMuoFkZwdij0BcrITlEfdEiugcDa38vqXVFvvmURh
iqxeRHweCRlVZKsanmt+HUK4B2lz9EBAow50jz1wXEwrwnS1tPxk4axTGsPbluv4
hlwoUcGhLadBvO4K+g2ft2oEzF7WVecick85h5vDSyjhetJ6FM83MYFSM0vlD3Vs
ZsEAonDDSde7SYdyMzXmM73X7cTM4PGgWCUm37TpNb7C7WYbArFjfjKB+QjlSJeI
vj/nt9O7dq4b7khiAaOO4/BEIGW/KKfBB+xD1rxSt+mfqyXaYm3CNqbW+a8B7Nx2
rBEW4GstCvn0s5+iqJ11HRJJmmOS7JUP90GRWNPHItiREkFmeJb3uJbWTJlySFQJ
JJ3q86T9iTn8Xi9mMzXvxbLHuBQf5euzQozUM0h6Y/TR4ccJ/7FsG6iKm28LQsv9
MM6/AmXP2/Ba8zln3yJ4+zpnC/OkyQXQq3EqySsEnN3VEeU8ZiXBN5mOpWycEIN0
x40iXXAKrryLfcJiJR/tgl/oVM/fE2YoV8mmXB+/PfSnbCvrre0S9ZvwxJIdNBKG
5GQKuu7nOo5UX7/MGaMEUazOuoSQOwMegHvNwuhxlxujx6w4FCcHKFTAQo/e19EJ
zat3ZwfgirBl2fCQ0/nCOJXDQdKozjj5Lysi2VnhSzn6UDDaCdudUlKyrLFHNy2+
Fn8gzd+JANg7AWVaGNDGNOP01+xm3hgFL3e+lQmEwJ7gkWJkwWq6GDwz2NgdxlI7
LEU//I9mOt2y8xT3JEM+/aoKKpYcQLAawHtRE3yq+g7iO2FIq9B7C9h0THv1kXx9
/GKA09iuM4K4ZBvOFAU7u4xkEzF9uaoMB4iIxzudjajzsNvexUxW6a7wqu4X4ruQ
oGT6ROBy9dZhSLBz/BNBXdey1IBF942tGnb2wITjoB4DDjipWQfBJizLI0uvULBI
azCnPx4xzNm+i788UKZZ1WRfjaggdh0p2oQEe4w0SeL/ZYS3fyyOVTfPQEd++xWE
yWZ8EN/v0AbN47xQ3bSIPjUxz6Ql4reDMe+7jqSxqiqeX6IZILP3tkJb6IiWBlEC
mpVeFJf9kRq5hBnY3Tbh3xMf+PzM/Ch+c1l41o+Hr2t4IOS6WOBAp/mgbXRYZjYe
Wm5xZK7gAJrCDK7f8CGqLyri5aS5XFnoNNBjDIR4IqeU1moaogwO7Y5TjGcb0/MH
GjFOkDJ1DPhIUmyqW7IzBGahN/ulNRkAA59KTCLH2xjSkJAck4vyDgA+ISQ8jr4+
8YoBdHEkUmddTLw/921O0mFPhLmDLlnqamzaa4t+ZTvJZnzD9AtDcMfKwd15xVRE
ARw9eyqgMLzmiib1vjj827XfodRWvLSQ58B3KheZpju1mdciGHASHIwKNbvJ1sQg
C+zGoJlDZy6jsp30C6AieWih/4aN1uc7vlj7i+ldJa4+hmj2Ia3VBJQefbaR/c7j
ngtxmeeWP3z7hafPllYgNAEzRFhF+eqOAEpXjphMSEKF3lpUk1fFXDqvvNs/fLku
D4lPLA1ZIGYK0Wj2mq+deyANE2sv92yxWXpWQVGC/ZasgDr3c4/damZl7hRpyIQr
4sUQ16VapBrTbABOFyFxPoGs90fA1glrFrhanSawPb7QUT4I3PUoa8vyz5PdZQqw
aGRRFsLyUhU8icqay6bGJrVQfMhkVR51rYMw/xdP+5M0bFtNn8/GXHTHvF6KM1Ei
8Z36SeZPYLa4YuOUBCXlaZviwMYdhczxalAWow91YKnjkpYiJ0DaJun6W6v94rcF
JmrXf/9BP82B1JvTS8x0MOfiaLV8lNcfM3z6ofMIPP7wONBHlRCFme/LHraEAkEx
hqAk1yFZ7evXpEkLoSAD+yRdQpc2QGrweyxD+ROlsh9xD14l/7UpQjv4Ouk1u1Jx
rSTuGAvgdwggczf3q6VxCMFdPPphxOTcXvj6pyPrFC73Sd2okNNqWrm9zduFalol
HiQU26X+CTMQskaaYonDvwms2Ok4hiF2lyl+6iaQNeZqxORFs2UllfrQ+2g5gdCw
PKpYl8SMj8XytidG68H1tPg9vo9V2DLS9LY26GbQfDGPw4o8yAeQpPDzrR0UPWrm
Lz0H2fafh2VXopY2Ljc5eSzqKCebP7oqFpeP54O2rBG1w10kqm4VWDSYZrHQe16U
9uDWBBznikW4tL5h3dYSlMfDk5nGev4uB3Ta7NCV1jZm76Vk0n9PqFnNwqCg2UD6
F7iRQJWZz4Fn1dV7X+L/S+bSqHoDdebjqlQgc6btZ//dRI2FXQka5SR7IDASGBoY
PPGZZF+vYyh7mu7H+GqRQGcWY3b+JE1rUHFjb7NW47R2omgrEm3e2LQ/WClFQHvm
T84NnqDhGKklOZFtzABnb4oH7EY8Q+Q3tsbXTVxBrbakEzlDgvOjyiEGSFg578kG
vzsq1E8lR7dDMuoi54jyyigblrFKeJ+Nw6mzj7RK8pvdhQcWegbC8jr7iowRjrCS
0vjxnppDqidrRyF6hqkDlYdoIkTbeWzrXW5SZ1mz5ETLzA00CnE20uw89YJ9dwJi
8JwjYRwtej5AQvHbeiolbnywTT2xJFUO+gLCIf9Ch5aTUasPwLO+oUe61f6dz/6r
dFVsJDiQDsGrGcQDSp/Ub02eLViUICLEgarDvAvNQCnwAzen9tD8FhE7kcb+m2dJ
H94kykhpafDyhITNSuGRYUy3r3mIbs/zR8s5MYJVk9a/FBB/8ySk+oy0ceEP7ccz
yJcCp5FHAnDAU+rb2dEWk9ZulowmnpSTopNiUHShHsfW0z//mljmJeY225Di8GAS
+MdOzv80fj78cysm1kZUTHMSOw/ViR55D8P+SNVk5w8z6RAXar/rCcQ3dmGK40mg
MCKH60mRrIlpH5q8P7Cne6YsmjjCEkhyInmlUfbPOft/1bJlqPzpbYy+mUEq7VTf
vGGIRIONfrBMlSPG11NY8qvvzDF538ALhURSijpMR/JA5MKx404vjfTqOUAwd7/u
bGvf7Kgeu8zdBMsIXfEaSP7XOPmCxSHZhLdcSkPuXvYPk8HFyCi4tdSOTBOtXEiZ
6zxrXn0HzHp3UQ4FDkLEOF5xUzfvZJBU2GP28XjyoLhHLKG794DntC++Yte62Xrg
hUeKg5BMJsCKXIZPeVFyvzVl+0NU48lCrczH2UcWkubJYiR2fIIy1NPsVAcH4JOh
TGBazYHd4/anKfVqZzr61xJYsvjsgcvI61oSI0W33NefUah/9WJMBJB7C5z1jUBU
o/pUXSQFx15g4yRD6LDVVXgHhy1d02i8s3cewECS3owbpXoMf4rGYg8VVJqnv4+T
98euqNEOOho+1BEKK52bNbkQF66jSgamLDQPwcjpfvyrxYrTb4dCu2Kdqaw7pv/w
5MMqkPygCFqr5SgGU4ezkS/EABG5jRzGygSiLQNHb2rDquwnaqI9U+0TdykJ+0+O
d5U1tARt+yerPH7fytbEx/pfdgJq6cyKOqwlr3zG7+evk418XcgcUY9W2Xi38WVY
Z2mb6XqqB55MTA9B4VWjttyp7Bf78TIS1gpGkdZ9dg9bu3M4tfMdGqPGxMnu0G6j
Ivmh5LFgXDXX//4F8tn+0EONS5PNXjAHugE98w2/Mta0TNy8vzE8BAg6HELXXZKB
Iqo4MRtdpk/eRSJYj09Eh/h7+kF/rUgpCgpstKHSolyDlIIwLqckdeR66nKJQd4n
KxwEhDWoTpHPgfEHz3OKxFbqaeUi+KA4nvrQro6eDSQ2cQ1e/2ePpeCeOZs9Bwr6
mbVj4ZyV9EW5y2qoyJYDg18uWkSIDHXx08j9rAcJayk9yrKlSGIoKwtHcJgfqe+A
vTDqOrZiP9bjlrfujaqgQCv/S7hzncgMRUdgbL/yIU21nzGAZf/hvvTgBzSZcSGa
vPvh8A1nPzE9tVwoHa3Q529b6fzWVDuRYU21lioPn9YoWdk+2uZ//K/7R5GBRhj8
PUgHEFlbQeik278valQNLaINKl9Bv1OjpO5xqgmyDMK0zH9qEeDn42B+3ioMt+CA
MZ6t5tilJdQIf8XQ9G5YoG6KbH3Ph0+XNh+8HN06pwI8qQPlPz6y4fGl5vyzjKdC
F7B9/foWJDoGwZNxTXB2UeoJZuFa5lZbdbZkt2IJDb5t7zBQaiaskNUm1pGQzuFf
rIhgU7N0iSSiGgEf9hP6Tb8jcLZFIX4rSL7wWfaZHs+IElDMyROPthJFJtUrkZgy
kKpRr/Gnj+fnOQFtip4uZDEDIdhAQEcqAgbKHzVVM5xh+tWPMssEXKmZLPL0mZAV
ed2B/PfH/Iu4PgcnIpZy3H3vb1DOG5RHXb+t+LR3yhuFPJp0rLaXwDOQlDgaVGIT
VbWdu+pkL/K4I80dZo/9pnQLLJg4e7BRLNtX7Ib+WtKm0pBYUA6B0ncNbmrGL3bL
YeTZ6S0ehjWuDlT1X0mbqGSYUv24rfriUO+OodCZdy007/zVPmYLkCorUlX0ZtmN
/ZJ9mLJHoto5oFnU9McDMdN5iuG+XPzBa/eltX4E1Lx2SQBbKmEBwAuxZ+IIgMgK
e+wlEsI87kivDwp6upzl7AxR0qmTeo+3e2TUFdX/9m4IzUZzupgp26vo1UdltnQc
g1GyR24gK4VhJj7uf/U3ppK8rIE3OtIMV5Imly4DzPxj5AyCKqH3br5Qg0C1Ms7A
G4jotIXNK9Ep42HDGbyqruQu12S8oLv8X8wnr1SMS8OYBbWWj8p35aWuhQPSkibn
rR/SFADUsA3stoldUPfDcBl+onr1yWG+1lvDKVe6Aem7Fg7X5/AxGTLHy83pqYqV
DS0Wnl7dWdlTdOjcmrKIpZTZ69IN87jpsOpphNXNc6XgzxLPGK7PyXtcp+sFFv8J
dxrVG+VjQ0UvFY3CWyxrox6CO9c5HZSkB72ktvI7zHz4Gwx5nvQCMrl7h81HJrN3
3HmDm485e/BYONlU2GMGlCrrjWQISx7BRzRIxxd6bc+eBmy5vXKUrwxw86G5ajzJ
ebH9OXYOA5NlR6AYe1IUkoafnf/oxdDmvrKWGulLyXGMac6tH/TYdK9QlStbk5Aa
c0EPY5Oi7esS7LX8+1EY64P5sUYqd1B5kWlngoF0AviJZX3CtFXzkXRARWdYUr/g
syTjqjVuvhDb5ElMjvx/DLiDXW+2nElu1AXMnI3ap1FyAOPM8VP/jr66osHLSZX7
IApTi1HzU7Ov/WrT7ZTdwn+KyTe6bKDeVDN53n8wqUo1pFVWagefPA8VK17D7WI9
Io3gaU5xPnq8M+a0k0GyupYk7OnFSWz2MrCI+J+1SMeMmIHmkU7eyNpPQP3Z+bl3
99sTsoDWH1+LtUPETi876/CBF3yCoDfOXn7MZIpMQpn9Vu5Zzb8moFoVm/pUUgGA
QKLgmZ1XYzkgS3Ew6foZ9WTCNNK9/5CYg14lB71Bi6RXVi6N/VuaA7G93urEztf1
XmND4CMT4q+ApXigoL3dyaiT/PbqFI3CIiOA9JgSZVjLeeDOMdqj09RjXBfHDP6f
oftwpB9tc9IHAXGoZeNmm8F8b4JpNwQO7FpKlTJ3F70sFZVzcuA+3EBbgCJ0kj6E
EEYGjgGPox0Bv2Yqg8ESEwSHnCMMrTxcgQOANyxoA3LlUo2GaDsu+NQAMydhrIr1
7PCYFG5+oixWUsZyC2l9LaxNTyiqXZ9DnhBC3Ce0HsuX41XZ4uQpLti17Ajz3y/5
/wxrXq1Xyi7BMGEsFAWQhdC59BM5brGMve0lHbbumm/l/25XiqCPsvwSH0ia/8XC
ghfAQm+B2J9fAu76GHPuodDhWY9OlM0KlBeHCS+PtB3+xLqVwnaaPqsknFGNxxCR
epExJsyTxR0s+zDk4Xf6c1YwasxkOgSZJipEsg9tckPNDRkTEpP5JOXBjFKbDfI4
fNc9s5mphTwAsAwRm662UfLjB79K1VF2oYT3lbekAWSe5FuUthWLd/f2FADk/sAs
/Y5ma0M76r0JQiYn+h1bCbxxaPiMz4vB8FE6+4JkO4zeZ4u6I0xO+mPT+99l+h1N
Rb81Q1U41+NQfNi+DWFHYpAl4bfN9x+7GA8W1ILRJtCnNokZWFwuJyUirpy93riB
DUBqXz/VuBzqEyoGLU2/fiHuwY93SF0p5nWUUqKl9qJXAqL76iStjCW/H6G1spYk
jzDy0V+1uAQzLguFaazcrzTNrYzrGHbKu5MNkBGPPl9IW2v3BSw/Uh6bEW0ZIOwK
gd2GTFd/Nlqtc5nix1PvKiNkiiZlv6K4V5I/gPwNQh7UHXNk61cOY2F19ksBI4+0
g6siWnl/FsfmAfKpYWoOGV1uF+uhEIYtOYCCLGS4LS9aNZrS0d2GgIhetjIL5jXG
/MT28QXNJPSUH2YdqcZWWrKcFdCewuSkNsaR1u/vOjiBCu0fI6ZDJM2hm7tIZzS6
dXaUTlqBPESXZVFFIfpJaNF2wu50DUW91II/GcRK7SQmhcxqRYbD/HZFI3RY+wWg
6audtdFNXnu6ujGPmA1qNV9wSLKWRWAH2a6Q/E0nHEnwvNUKQNwEmNBhU/qoPwlN
CfpcX4EyBI1Jt1UBLhbj4hOsnP5NoLUTWH+YOkAYUZ1eszj+8+FAkSb+iUEez8BW
46X/OPlY1be9Cx4QSjT3whilcCkc80NPSza2G+hy46PlMY5QSZjqyrY+yXGh330e
mFk/+C5sI84uJbOqLOmsiZFgxDnJIFC1VMpPX+bv8LZLbG35KfvH1dlHf18KRFXC
m0H4siKjerATDfq2THU6N1WJuwshQlrytlmbRFiNW4nnvgRefYxGBzMxtmIhSG7Q
0DLJ3cfqJv7kLtplBKVody6/tHcm+1aAIwT4SSTHhezsRwx8jKsoINGlDk0HitxZ
tOfOSan043EuAtpXvm5jM1OrHlK+J+P/YrQP+x2lFcpUp8uxAhWnpFIfBB5ap9c+
Uf7Lxrt4pZ4PamWnWlqGco8XEh+UxN0urTJ1JztRpXao/7D/3bqIUgSVcrt0Kao6
ERCaEBY/clzAryXlmjbS56ycx/TcBx578uDwfrmbiDXSsWzka7pQvsI7BLvBK13s
z01yV/5KrZWq+ntsysk52jXPa73Pic2sfAXwI1BPmSas77VU4tbxgK90acJVUQGg
zRV6DTwoksEtz+x81wamSUtSc7FfMRvg8FsJdUvvdlof662SAlfA2xuVGgorsGLZ
hwXINX/Se37DyFQjEC53VprWvMJgGKpUeNixmG+aNYvr3qg9dwnYc6nhjiz0vS3j
fq1wEepuN+MBxTLKowrLn3uFPNQmeInH4h3jL4qGIlPcXXaBRsdNd1F6xaIJ3qKC
vQBKz4+yYC4BiTVs4NQXowHNQZI6sp2/xvjWjCYZkGWQAV9gTPXS2sgBLMv5fkiv
S5wVEZkvpOEnGKzFsB5A6oenqIg4M2WwucVoZyAJSH88Hlprwn8XWMZFLgVaN8Xa
LdFZyTtV6xWQWT9naY1O/u8vFIT3ENRC1OOJWBrvC98TOHBjcdi+SUoHZzsdV9/k
287iKQvJzziP6PiTuOLO2qvVHVgzjVCmH7kCvl+Hb0iDJLVZAPJuJuhUqJ2cObBG
FZfFLpsdijrKXMOF3LuhvdQIqrYnDAGKiMIm3Cs6uhH5BeHLovEUarH5owsjZufj
HGQLHJ6UW4749PCG2GRqHwJzBGcR+eRgMdNcQbEWEhDya5brj209dvDmszibIofE
LDH8v0iOeOQRhgTMXh9V9tfAtCtykndkbZuCMX9Zhk2TOD6VW8Stlg5C9wgRAOPW
eI5tpyyzpJUhgmafMOfKJA9Bktzl0VKixBeNlRjh5g/aPp9DtNAFEzDEpIB6oknE
ePp2mD/XK2QIjYMDzxjaN5WIdNO6k6y/+EyAr9J5RJGQH2z/h3cKVwMV6qaf4eu2
UMZ7ygqLbSKFvtGJsasVhf7tlobHsKRDfMOZdEIre8+3tFT1+/8tC9QyUcWJmK9T
uMPmtj8WqeTGQpgsD01LPUU477XMxQcc6yOvnxNAWH7Ey999fGb+5u6qwvo+1w6m
wQVAztxquXzenw8DNovOlx0OzeLFEcidf6Yd6MkdQRy1xTEir14KTILtiN9VFP4a
XhgS/zEPQsZIUE2Iooly2qL80lDyf56EzI/XfnVXo4AphdekNutJR+3Tr0HW9ySz
5DIjiqhugVuVakAbMjUlf9MHMcGXylFnCGBetratuNo3QudY06LRGBCahtBN3hxG
wjvs/cDw/LCFeRMMPCl6aYCi5SkcxYLdZl5rCEbKJ27ruZqgs8N6HVOYffhucySD
m8HVocCnkI3PaJq8SL1r9xcPKHWw5+Y4Li8LvoohLdArrZ/0rlAXIJz23XMsyxa3
VBCSxRhiFiF2cR17fQAjt+qJmHlkEMtyd268LhxX3FGK5CO/VTnZj7gkqtUygkBD
y5z1HyxvGfPGnSdnNyMrK2/Lkv8lrjGhi4eGqyKZPsouvlIx88/JrUJDXNWAQ8J3
3l6F3qMWJ19HSllBmzvejYR6yVMftLj8Zll4+88UkZqYF85cr8a1HxnwUZ3Z4dXc
L0qk04VVHedhsVPSdIh35HoRnvrqVlE8XPtJn+58FjxB/GIDEc93y5GJ8vYv6985
P06GAj6wLlnBVkj3AHNB28f5b1fpVwAIo6PRNoWdQLFwvfDBxRxb+uS5/V/eSdKb
qETu4EOScDJ3yr7JuUJ6Hcmol+usPUACCvfclEXjHwKY+skBtiLGJw+KtprPD0Ue
3hS3duqDv787wMsFhts0e/RxZq2zWjhjBj8d3KkWW1vp12ea1Xis3PfyI6TLFI3R
oKu1I2NElx+j568X8HytQTutuVcyzRC067gZIxK4A1iaLZC9CsREQK4q10k9qAlw
C2NNLWjrYigEMeOAZmj26Bd5ZKEyHPNSiuqbB64HSKYjGAF7E7RBud2HAbFiBtIp
afx4sRkzzL82kXWa4WebXA3FdZYJZI5RQ4ifRK9ibSZxQpffZxqQyTb6rBgam1cH
BAhz6A7X4Ml57fHqzSwRrko/XL0wsG9CkaYNS5siJvMnMy0r2e9nCbqRP5vpWLqJ
PAbuXQBn+AEGxEncZPqhHy8rHLfUBX0OdXINti+qP9TPkm3X2Mavq8QA8UO3PuaO
pS3kLVXUkJ8ehQtGib3RQ66rS4/dXtZ2eYPPe3b2fInggU92Or4namjhricnTHmL
WvZ0YN8exQZvDTDt424sMwhnJPqDKO3VlkqwHwWTBVfmBDC7sCxT2OIGIxnCbTX0
zdDDpMGTy0uiCass4DwvxDPww8TCN7Mt84icERkG3+gEW0mNlvmnshc3ty9n3xQi
Ej+8FeL1+Scbt0oTLmOlnqKvxHkV/6R9FpzMZLRBjUDJhAHMWlo6D5cqR1QZpUjK
kYQ37pXSAIqo2LYSTowFEeeNhuHqRpQWR7+oUZI52aunDt5gLzNrF2vdvUBiu7S8
TuC9j+4YWF2uTbFTl620Xa6WwSMJ+sEoo/r0cWJYDaCN9BI9DJJMOnCN9foqcYJ1
JRfcLpJqZsu+1DQtHYlIytbK7SGpjK8AsqZ0wEw84gQz6dqRRG2A5YGx4eI6mtcQ
QZhWaVm45fNmxAMn3lURJDMsJt0/k31sKJVccHb/jk+DyZzwGET2S4HcK6e24OL1
c+2eFUZmXZWG7fOGIr7fw5Xr28sFojcuaozK8TscegQzMIBMaxcYpPuWk2GKVQXw
XoqdsP51aI4EjkVhgNXJJmtDUu2/9pjaGbHKG4nyhF7ub82QSmAV7PRXR1TyCiKd
zflovNAt7/2P2NjPcgIgkuvi3d9zYfWqs2KM7gmDZswh1hnXqdIhXQMyrLP91k4I
NEKiivA3L6oehJvDWbONB+LtucNRsRhuNWE4tDyIh9NNh8BrAM9UBqgBGeVWiaso
ylsyIkNnkp4SuN3fdwcZNB4GEc8XGUSsRPTNXzHLzVJ5qpd0C0l9pXdaiT2M7Eha
WqQ4I9hJrh+x+TZBkNuHiAXO91+APHfq7zkNXAAUMxzv19/cEwXsVyUI6mmqgfpW
0BuyJqzH/bQHdVJw6rqU11QXjmqvORXEraRvuhudJ5So6+yUJZYJkOxVWtxCn/p4
5cjFTU/6Qs6T63xUSWM5bX0BK+fPrZsMkOlth1AYQQgxDgB5t0oQQoME/4NQi+t/
DYavxDLWCzX3FVhmcMyHjZ+Ur0yqw+DGH/KlYPcCzmOw9mQO2fLetr+HFdR3ione
aHebgaKtmDgLXRD6sEW1zzZQQHjfFQkMkijuyAGyZHsGWgW8tmrSExb0UBzUoXO9
xLd9yah3bvSaKJ5r2as2c+SlAmSI6jTFo2Fi8TqlTbj+czyuY0Y3DLqQHydIt/Az
RC8Vmn4CnGJHECBwTCY2c5Vp2YF0PexS2mJhyCiMKx3bbGPEGWOJIa4s39L3IOXk
0d8Tc7FQU5Cw2H/53IXlxayvoI/XiFN33oNKp+VC33seuA+C8mSV7GIaZwXrgeyA
UBEylpy1gEG7dN/T/DWyYq11gTHPdN5zR0/ibzA20r0Ep1jMfIwmSoAw0clyXB+v
6m28hgxpdfzeM04KrJGOc7MWIKEsjjK4qA9gZflXj8/mx5bWzYhjbEFkjqLqePIC
Wu9VtYyxCkrIXxwZC5N48lG/jdgfOyaKZeyR0ZTjHBzcYhOvzKsnfWzojb5coPRS
hztgjysTDcJLqSMuAFz5LdbWfLE9Myt1IE1iYCYVo5kFyFk4AWnuyNrOlyHPenb5
hFKBroYTst+7DjDt6Ch4NeBrGifF5TRsw1aWoLQ9Oa25jSuNIquNh7zmtktOwgYl
+agth7nweYljc6MfME9kAjmTgmu/ilw4ftciTTxtVx49O+QGHZFXT+Pp/6eiMFNQ
0YaeOIOKThhM74Bj11zxTeMcPKQqAxNikUJ9zvMgRGg55nJpmcRnAWUHh8KdU4wF
dsOvVsOB7idhR5O6Ymznrqv8INIojNS8lhMEFBwb1xx+uA4vkFRWqZmRACcVixlF
4s9H6roc65Ouk9aCJJGK8agSghYVyYAjWnwTHupTC66H2Anoo/zR0GfGbyjVxzt4
3cM4xOiX7Wi/hE5CqJngk97f4ypFjzwN1uHtOlUMnZaeXEU0HgB7Uq6O5Ep0nzXl
kfM/ehr2tOa61H3ASRJpWQjW4D7qaWTelsb6TYq6mV1lSOMxXWOkOq9K9keeV4SE
kL+J7THbv4jHTIntUZWKXfs8IbRF+XJxau5qr9RD8OQRgztfzwhiR3qhdqSGS/4q
Zm2p2N5ZXVq/edn0FivqQzRnQXokmSOGg0IiwbQQYfflIUJKoFCHpJc7ozrG/jML
KgXCaJo0wK33iuD0XCvK+hBkk3pHRQMBKMsEnULVzIof8vBABMK4sMWXr8jt5U30
0VzuByyOQizTlICf7OREVfjShRNT2v4qMNRzH3fs1reTLb51SwxFQMB/wPvDODEH
rc5q/wp941Y61/Vu2sL39UtQ8AnRIAdytcB05Zr009lxjmVFKOtsCrbHwGxWf7zl
I2+aQwZhLqHWGvHenVf/3jRkNhw6w5dFhDOw2T7pLmD7eQXpCAYzyt2m2eDSnbuM
zyCZGtu2W5mVd43+PE+hJ3BT4KFiyWM/f4agrRlnwG8bbmAvPGkn/lZuGEGFKEJ+
1AbC1D7SVBW86xhEY89aGL7rYGjMOwozATc+GzKLEv0XFUN3g8aMsSdETgMxbFZo
frJkv9v5NmyO1djtZOsYZ1omy1tsVsgFCp3QqlhOrxCJGesH/57BqlEh0mygMqkI
duvzvkIIe2TNR3ou2A4iUIFiNV0fxs1xbRuXHuJJhbxr1iX3PbDj4o8pJfWOrxwA
+kV0Y/77AVtjYD3IGUH/6P3iuWBwqKRU5oxVy56H9itrH1rBXctAwdLChsukPg3i
k/vjdtV/Rwm8ssIlrqu6jj8t9dHmLevn4bA27Hx01cG8amO3xwiat5WcREFhdEjv
VEaRuGP9Pwl4W4BZ+jowWS4iJ2xXxwbcVLbMT8GTaYA=
`protect END_PROTECTED
