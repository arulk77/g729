`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNNjxD/0bPWuIEoTKzyKKJFTvNmeoJuv1NvPutjSfH4d
RXWd1DZbxRAZr3IvbG2ZVBv37GslOm6UQUYy/Db6B8xVbuiTH+toeDOzwpkyN3RG
YAmnU5G+VPhc4isN/9kPXnGat+1PoIN1h4tYbw2nW/1ExsfIRshq4S2+ML6nt4DB
`protect END_PROTECTED
