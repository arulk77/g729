`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aU9+7+Ug60T8kE2RpDTIV2WeSHnx7QIWeW3JTrDopq55
F/8TJcNUl1B9UB+63D7pO2I/RolbBkZ1U/ZPD+pM7Hjc/d4AxsoiS93UMwR03OnB
WOCIAlMS9Shu2VRxmv9bMFZMW3Iizu6bK3r6blds7dvw3LwoeU0hNiEP3sX2yWc0
9mk8kGP0Rij484KTx5oZALEsDyZ0HirkH2TV5seM8qzgfTRp0NoRc8JHtp9chPvl
RKHbaRSOfkiPrY/KfnesJVXkO/fKlhWRajbFEpjC0/GBlUOLENfS9Jx4wpdMcfD7
tYXc6WmhYJFLnHbnXOqdeaePUThcxyJmLXCFUHioaSAJ+3pfVhoqpi9GLqBkut8s
eSYvx3OF2Ix2zhuUHO/UdJQJ1ihsHT7T8sqa+OtSRfugGUYnLOCwXU5ZEXUBpv/z
qcz6OhATtRodh147Dj1YEZ5iSpzvm0grszz2moJzpKG1x0k+igQQ6VA1sjswWw3r
dEg3tHuOjPlkph33AiYi/Tl0Be5VjfH0myegaz5P5kvX5TnR0C21m+qbxLCZk6fv
25hoJes5131yvRp7slHHJNgF5/l1Yj1ADhBj71l6c1j6m485RgBCjHtcFpu8Jfum
ZGejrlWtZnb/EhPJeDL6Y0bOrEXNwOlvHmsSS+0AjWDnscM043WU0DVXPx0krm4u
ucK5iX1uDSdN1l/B3HiJsqhkglSXr59vXuj5qUMjOEdO9YdhQo0B+WMlM3lertUt
b1Z5sUkwmJRa26MfsJnbcW2zsjLqkmDwxUHve1lipMJoaK7MsgsKShCjxvwrHEEK
O3lgd8JF/Z+w0m58QkugfxsqfCzh1Fd95QhEzxwSyOF+RR+76FE005YmGauVChnI
qWzU9Q0HuWUA83c9WHm0UMmpe2sZ/nKwoPJB8FhuUbjS8zMagmjqn8DRUT0C/bBl
Tq7dIpbg+O7T4uEXV/mogEWrVUaj+qSijRm41Xaf66IXLzro4NgZS5vpHmsuMBqf
b4Q7B7ZqWFleWKaZEbvKLn+/qppVCvjVJfuxVRY4OBFKFTqSn4V1PpN1rRTFsmod
EICmwlaGkdUZegXX31sq9gQ+ebscZ6Z/cwfovTdasxvA9BkFAa9zvGwBfRvCBAw+
/HypCYqSyjvpEcmL5THVEHlmiqbettFqf3B4UHnSi/sf1bOSYjkvE5VJCLZai8JK
ozDNdIR7doIptNpA1yr44J1V9F/rVPnmumXceiPdxwCSmx9bcF6YNvp3jotGe7Pe
ZKl/+1SaEAqASBmL6S9SVHC+10i1Xmnb2i6btEGVqWSBV2IiissVv3DltSVPbxyb
39P3q5/jeFrc+oPGdRH0DvBh9lDEptJuFu4PLlIuMRdZbc9nJcouOJDcSwaj2/NX
wXCB3Z6tKK7TRyLAs06IK66ZzC2u7KamOgsQI8IzVi1okTKx9vPsNRkAV7RWgDNt
lVRBxYhUxyqH8x+1fDEleq/d+bYw/6xw4izkYc7bE4Nf+dKxba5MTLITDfjbn7BQ
xCbDeZLbXTGVOjrPB4YiJ6eSJVLCmHPcYDrv7uTNHrF5ApkqB7ojcAoYb3Q6vdgt
z/vkxUViIO7drRvPxmOXXoMkgCWSAZHd4cvnzUudPC6v35yWyfMiSPXVQjYYPwxn
2DpMPOoqoP903lzPtsi4iJfvX8MZEzUj13BRLm0I0PjLTXaz5mOA3eG1RK/KRZtL
t/rnGbgM4c+Ddv5EaSmdayTQ91Qi1AVtJ6W+EDK/w8+uiHiBPXAQ5kOQ0ij0xd9H
xwWht7mj12ltMSndg/+kObBSlM7kbI7tk7m/yNRos4rdlHI36xtHzkHtY8vqfmQk
GLOUFxcck4Tg2xY7wdZlpfcoKJ7tlmArLr7Zz0vgjd6KAwG0OaBDoVjgMYvGrsSd
qWbg46m7X4dPRNdPho21NvaaEqw9MrbckfyqBGFIVD+RcaV6iPOwmg5nO8bIvcOL
PvYQfNlFq7FRyM5luvT8tJ/eB+vqNGGdgRX83Olnx/K2a7VpMoXuw/7JQc+cjujJ
jTyTfWOoJZaD8lorHHLtZSPQjMTy97ABIB4Rw6vboemcyVrRxrkRWURVVgo+3nVl
fGZevy6Uv4jlEfrOe+qiITo/E5NFB92AEOn2i8Zw5TkEQBw5O1NSucnHN7zTd5i+
laOvEkxWzcuAmFc2hHdLkKu23N1sn4UF/AkMY0HPNQfCORuMh3pyTgufA1O5JXPE
YLmKsuBXgjtyf87FozkkkfsC91QdsrNR9i5LGZN22f/vhm3y7Ysk4zUZMDQWBhJV
gHYKvqpuUWOTyvBaVDVhaC2mpkNGGSo2A4hJL914BSZJRhZgd73fRbBTi2QdgH34
65epTE8op1pItxR/BDY0dC+jxN77/aVlrHG3ZOHUANTrVNg4pIePhbgzPlXkZHah
b+OCgEAncjmuSE8/av34SfmCoVOrOxM2ZuT35yolX/rwGZ0JqkzgFNCQdRbphGzf
TSsoG9RclJj5aof52TV1Cdi7CewtH0eerXMep4QrzjStUGUXfLMnTDxuEEYhg659
zZvC7YRUYhUkJuKAuPb92c6mjkoI8n7wIGhaYPX5jkjxvlFDfqxjF2JmPSlsKFRM
vVqXiLZ9MxFPSBe8aaELp45KXe5JuWCZymM7B0odATl6h1bqCE6Dt00qPNrqMSvO
byVMoWsT2f+RHYOmPVgQF58syGSXBr4WG+xpGs8/61JZA5UPWwYxgzmddTNGOH0u
KzUVkHp27hw/jalkoHezhSq5znCglW16IBp2ZIKVDDGDCfRZ9WibAtsnnI6Y4QaR
pPkGXC7LB6lt5SAXeBAZg+VwcdTdzspEh/bojrRlFpE0wOXJT+VUfOq1VRvm82P0
HA9eLhq+9nHsIlRh4P48kMl6jciOk5HBGW5T9HV2ke4REyWkhwTvL4B2tVENXh0r
hp4uUlUxZr0KY2Mlubj9nkU+wAWdlZVGhIFmwnuMIAjuBXZ6k3z6/YdTXVJ2HC2r
1CTvxW5r9MBCKQlwPv14Qr23WnXI6L0FVZBKgbxBzXcOS5m1M7ujisoLIZbO7Lm7
rdlITSngvRisoF6DCwTp5v6Jzj92eh+yd9Mads8wPSqfYeFMBp6tcz2jongGx30D
wNDimkLDe8GydmMRYavoz935jcRY50294Cwhk1RUxi+qks1r9i7S0CK9DjhhV+K2
dyg/Dyrn4SI4Zz2uMULYWxzYx2qMwB4WqO2YdeAWxwcPH0w1Rr3YovOGN/kENmf+
6nm3cNp5XPTqMNQXJT5bnuwGWvxo9HWADHY7rh+dfq/W5e5U/nF77qgX7LJB/SFW
xB46XShtmtZF/MLGnYl0+N/kNLoXJEetZLRUta92Wo9V+Kl2/CqxtqjuP5LqF535
ehfAfYgNKBICZjuRYv9VxfTD8uyMkoh45GfPaYaC6vtpKcqchH6lwsVdieMwJk2R
AplRa5CdxDjY94e+9ii9pyxS/+PLcsOJ3Q98Gzo5Yz0ykVjJDPU4XH8JVoVAWzYr
Wf2dl/6+XTdFGbXtEnMlbMid3JqP5Mw52g38XBMrilDJZbfy4usJYH21yExRQxl0
n7S3AbPQS8Q5lIa0XnW+J0r7Nr5tTB5Y5hWEdp89qcbXdIwJM5ZaqRN9/XIZcP3s
91kYdG08nVnPvmzCVcJE+WYaz3WULb5SN+AN97CK9bEmckhnB/WCUYpq9yY/Oui/
ryXNSCGfgZjcwis9nfgL4bhr/3UCn3hmQ7oIE56WMbQAPv/KQh8qVSpvr9zX2PCr
3SLNAv2V39HUxQ8Qr9oUHh/P7Xxk4zSXn+QmW7rA5qOHzaoX71cbd70RPj4aTEwk
bxwpwe3uesI2YzCWOyinQ17BTwiG9E/1W3UjSi/yVWUiLG0Ohttgl+ooe+xeWLlk
kKw4M/6zFlG2qxefzbE+7cIDruUQUVpvrl0wFi/V7v35ETbBtFQnTr7tsWxAmqw7
Os55SQsu9xEuXH7kvbPXjQarizyH2yTanUROY4YCYPr10gNOqlmorPNLQE5RexfE
eq9tU9umJWZbtS5ktpiPOvRh1cCKLW0TphfN3PGluHVBfGnC3S7zt4dTKmyjEUnA
`protect END_PROTECTED
