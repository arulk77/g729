`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
88v8mM6tMaGbYQZZ88gveawz298tLHBRtZ+1nqcbvsejtwL5NddGv0QdQ+Lcrk3K
8cNcVmsTqojrZZFxWciSyiU4fgQ3cu41W2gnIeXiJ4ikFYocvJfolbwVTfXk1ZK1
RnJJQj3nVzXapLKvCrmHB2ULvh7+TbBPsq/44lB9uD9LAFE1PMN6lIHXG0TFpN4x
b1sVya7OqcYgcySZlPJtlDFimrYuicpaZRDOWVJU/JkG/n8yf/Z2pOx5bp3zeITU
vb61Fe8T59reITU7WDOjq3O8/RTSQHi0LfuJyaWOfqudtmPbeCnpMx4Wol6AKpAS
e3Iku+SXrPSqap1HMD2OPOdpBhSPwsp+kFW+VLcwjvg=
`protect END_PROTECTED
