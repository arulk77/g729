`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIq9znfPQDlT8JvBQBxsdtqmwptcpzjJ/70i6Rshuq+6
V4bpgYnzqw1Z0Pg5XQxVuKYqDJ3cQ65D2BQKwz/yRMAlANEAx3EmfL1sKR1UTARv
ltZuqLd+iQunNuEZfiHf4dS7P8iUzN/nU/0W1F1QHhxk3iiBrjb4gCS7TMYLLISn
LvXczCnVL4XIMHIwm4eFKTh5Oi59v0zsTvCs+Ch5W3QO9agiUvZgrTcxjzxyeJEB
g2O/N3ezJs1x0Fn1lp2rbZ5lZYsR9ITWG2QjkxFB1HNSbLw8BgFewTZ1BoxqUTUW
kh3wgiVBTDS6MlgZE6kJJN24fbCkUTRo4KIXXqdkDn5IHw4xYO/Yu1/jd9/+2emf
pPSlB0L3KhaPAd0BIXOf8yog4b60w+sSJt9Jl47FvjtHglVVq5MxeoDvLbTg8H9i
`protect END_PROTECTED
