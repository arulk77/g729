`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGj9DKJjMikmLAzpu2S5E26owEnP0Z58pnJ1PFGswLwj
b1fCOY6ot4Xb+4orbAGagyU86KH62wvYJsKjMnsudgJITEb5pwEdXjhyjuJoQvdS
PChzSD5jW/ncjYb1+nHkFJ5mlgW9C/b+VYjw4LBBC16ny8y/EHHQ+GrTL0u/6WMJ
YpmlSDSn931iMx7iBgXPI7d7RpsGHwvoLppKLm608Kg4wfZaBY/PBBAREYVT6xQu
yVAyCQeRiqJNWdP5tiJIAbF9dRcTn/hPIRdgGP3tGMShBHwspLVTMCnZIo9X/aWA
93tiVbTYqopk2XSJyyNiNuvA1kGyEaB3IL0QA6qkL70UPP46onjhdf9n0vUCzIdD
niWtcPi42NKxtjqxDBOmAIppHW+lKiNO2QgsznzJShE1E8uMrIXxKE1cUrZ2XqY1
`protect END_PROTECTED
