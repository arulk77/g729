`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
KECEtLUvjZ9iVkp/KtWK61t9AjuZw0OdCRQboGBkQq7zk6FX5qiP/rgtdUbO/4xO
L/dwSnwVg3DbgqAo7obZJdAxwnhQsZn/qvFjX1i7PMoPeENV7kw4FMwDFJPQGnf7
320nrn6JGRRj6bPH7YeL7vId40KCojGfdxLnMGtEIUDKbvIQ84rAPk+Ab6sZuSNX
snxo4tKgE5oy1DYwrBI4b3+SGw/VaNM78A4vLdi3+3aNKekS0CGOc1RcyQlouecP
`protect END_PROTECTED
