`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePuymp8Y6RPOukWvRSz2n46ksz1jTNRB7dE03ecsAlJS
7Py6NMM0yU9Xn0zkx+iZGThWf7UGe9ujtgUyB2AUqPCTnNG5E2NQ+gvD+U5UFSEL
H87DxWUjNybkMyo100dZxnCZdaYHhtZeKN4nv8vlcrhII1X84wJCcje+REr+4aHo
RAywP+Zdwa36Fpcqwf/cG8mvumlYedrV2JMzawqbkxiQapaAceQ4m8AjsXF9eqwb
n43UFWIWdCJCOYmWgfPsi1n7vGzqTZ5nPtzIiku+ndsMvwr5FH1bfu7dXFOd/sV+
+5pYekLfS/JkMWHxpl9w07pBkHYrZNyOm8aL06BZcvTBc8K6YHHstBbqrAq9gUZN
ORRCuG5ZszhUnzeOnM9LsTqEcgxJY+LGjFuuX/Pk42OxVZ5bkaWvHlwH7NaiJtuZ
feMzGZywlpSEsGQaHCk6pQ==
`protect END_PROTECTED
