`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4860E6BWdfZosy2ipChkDOcay/PeyXFtDCN4BjYK2LIS
fVXGPu7oM97ZfquqZkcRb+Q5HKGYaKH7vUpzRVAQjhRPIPatL1XfljOOdldKVB0v
jvDyIDoWY5xqZl3f1mg129gBNCFT/K6z3h2NLkSpShZtjzw32X1sbYQ1+UmweJib
s45CKTEcApYtOVzaoNoXmquhQ6fWt0JHRpCoieyaAwXLtq/AEFOOtro3ek+UCqz/
RmKWgZJJd8hHdnzuXXrB3g==
`protect END_PROTECTED
