`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG6hQE99kkvMaXPOfpUwrIzrsnkRW8jyLeX7chRSuhUa
wJLt4gnjdYUYDbFLEi4IxqbwYO5EgX8xPn9GS98uQHej3ZPjo8C3bgCtstqbv/sP
Pr6z7l/Oc6sDjidelUBeG8uH88dZnH5bVioUlVqBXQGxbX5fWZfFYw1GCbgphbj2
ORs3gxy9ZajADxwgP4y/7wq2dHgzpxlUOuEK73myU5rRvHLjJ5hbQz4Kse8Y0+le
p1ivOJMy4d9+rvt3yM3qSUN5rcUILpDpwXqtCo2w/aeHbjkvYjBvWArwQX/ZqFI5
2E2eEkTs4EqJwH1oITDlK+c/YSP2aOLCxzaN7IAFJ0g6YOwvEompZLWH4bibgWSE
XYL1e5KM3JbbnQkNKL/E5dzJ2mcRANK6giJpqzbg+nbH6PhXo7O69/Q262YKYtWS
WvB2BeSS+g43e72ecTL3BkJNg85/CqnLYjkpcrv/GAJB1fyx7sj0CpcDAVEN70/v
k+LYSbgKFjAfeCMA5YobtRu9Abq+lMcyFawXKbaeCQJjlTTY0OAIAmhLA+97e6UP
9owifjsV+zCM1ACgeOWErncPUgD5wVzqKYBkgpUnrsDYetnvzuK/TsxbLXegErbl
hWFG48rcWbcb1AkfFBFoczrWPYZSb+b1q+fR5L8x4HyuNgKzCjy8KRPIgUTvRz4N
`protect END_PROTECTED
