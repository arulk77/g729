`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCLZyigf+54KTZSYJLMhTFl/YqCtxKTWSugQMExX6rYp
yqxkEHH4M5sQL6odcGb5cUk1k1DUBK04cPBz0ODi3z36pbim+/B+qCL3PyvWWcYk
Y0+UROlvqTqzAFOtR7bE2rSFpqEuqaJE9ybN2y9TDQ9ZIg1L1eUUGqxvM1fklRuk
tydwIuF8rWOCfb3k9NYUKiKI16TL9pFcuV0MVRIuQDZZhzqul8ftQep4dOayQBbH
73yOLT7jhFyBj6AOgxZEdJ/WrYxZvVvSsz/OnKhbjHSAa8bH4+UXeri6TJraJkgM
s19gASqLkyjgenmQwWY/709I+EnAYaxY/EYO+poUmDnJDxdy4/7FWs1co6bzYfXS
Qh3w3Y/7QZ3+KOnxwypYhrnwU56AyyJu8J+qj4LI4QzlcNUnINVcXID/Q5F2K1H+
ss/W4y3ci/A6p3CjPo6q9R5emqcXe6h6gFQYzbkNOXTq7DlrC0eVfkEWWphU15OE
Sa00gNwtThdw7vAo3oyJHg==
`protect END_PROTECTED
