`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLhdWhmDaew69JvdRzHrKSB2O18sgLy73NUVUZdAbRFT
jU3wnDGoaVGtPtDb6u1Qnw64I/bTxvZ5pTx+C85SZ2zvqE7PMcy7m+je1BrBBVSs
eTi1HJ4xP3b0OMXvmedyfltiKgJgDaQJcgFipmfbSLRVhK2/J8xZU+Q4Y1W3yyAW
fodK4COuBcb322BwWe+xlVboDNJX4ckr3c30DymU07DQNy/ZufeZCqlhlzCK2AiH
bgHCI85tc5WOUNkR/OdoGqCLeoYM7aK+5dk2OIyd06VSheTLQpeJ3wtFsTBLYsb2
Kkmk818z1trGsqJUYi/SJC/wCZ4z8QScFbm5mJ+CKRsPHBT4LjZ9/nqvjwbJslrt
58uTnNM9KoWhCp0gkktIk4iDiMTO4EK6ijLCugLJWtGwmNTuN/tRZW0SvcTE+k9Z
`protect END_PROTECTED
