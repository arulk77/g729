`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bHS1C/wcnHp+nSrtrzIjWuJILuHMYU4bOAu7hrtwkPn7v0LdDM4YhbUHg1zZ3zqp
Sm+BGq5umWAUqN+DVqE8R6p0LrO7QuyAfkL+g4lpSG36OfosAym8vaXFOiy0DdBA
mR8fzMxDUvELy1RglLqLeAfFJfUnJWBciG+LGx7bQyz8mbAr2C1sSKW247B+sPbX
Ba0mTe7b0BwwHYRD6ezottJXANgGdpfwX3Uv1+l+ZS9ENsFKNYOy9VsnUcyRrhk4
`protect END_PROTECTED
