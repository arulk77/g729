`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJB8lvxI+9oYUvewZi9iRLDvCjVkUcGyEiNxsYeAFOsW
uxxjRY2KJYoS7EOQmwRGoJtx4tXlnrqUMKmPx9zwZIAentaCBMYofNsBliNtPSQz
oU+fxKQHT+liUgmdnSbS4i3HyAj6WpiCqTiF8EkggzS45Tj/9hQsc3fURSHzaX4C
`protect END_PROTECTED
