`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveH7YLDizax11J0f6x4OlDaMzVqusvU5yQ8sWB6knrDgh
yYbv2dfLrPgYI4GrQ6WnKyf7NiRWPXpxPavgecFdzLx/mlloA71QaIUb9aNe15qp
fjNwy8dQQv1H9Xs9grv155cVOpabCa9gCLx1wVnsCwqPk1qj3uRWMKURK3vS1Qgq
/zUvTncS12CexaonQmcgWB4xRW39p4McssyBFBHO8dqCdTtepp9dqXdT3YzUEGaE
WUZOP5Md/jRTUtU6PycLMSJ9jvuZPTwQ7crEw7ZFFiLVeZgPG3Md4+k4qHTW04cP
e83YentkHM5+pAzLUD8jAdtgge/Reh6B2fDu8Kltu272PWkcStgkeULrMHJlp1dj
EtO6PPDiM1hKgahLUe70qGb3MLexs80aCeMDn1rKMyonzWtGInMjjfFFCT1j+XFM
QbH/XNiBd4+t9w8QQ5h/EyjlQXwkvUf8pRAfYhWa9TmvSKaPnthMM1un5apj5XWO
YwB5FTTXDIv0fkqYgfdxao53m6jiiV4I4vA61cMLgHjgv17OKQEw/jCKmqqQvXWY
`protect END_PROTECTED
