`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
MwMP8LlpH7+Wr/zP8QuTaQw1Ytjy9Os43FtBlzMmLQ1ryomogzKEM833uDvSLF7Y
zivX+W1RMFdOs/sClrehTrJyniCKLw5j+Al8UIqTAyEQK5wQVI6R2El0bNploKSW
+JKaAy1wn2RQqERfqBcurP+mMfSAHuqwsU52tKRBUdDr3evRhXhmqe6VwBMPxrdA
lY1HrrDqmTPWeWjFUp2uOydSNS7KEib6qzNwTpag+REkZ//g36k56BaWHFx/UiML
XwTbkT2nRFhvw8ntqbB9+TkqKMhX1/x5d/IX7G3eYbo=
`protect END_PROTECTED
