`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePqFaCH8n90MrXACdMPGqgV3qDZqtl+nOQmC7RuhmgUm
GpD7yKtQDs1WYUifzkb5ajTu/zWZxcJpoIXN8O9khTxsts2PsbzeRTycY76foGzd
rJ2ebeXY+7yLOnDHoFup3qJur818Dd60AlYhJ8pG3+Fuem3NjITXh/vZo/zeDgyr
561xKbvfZTMMWNcLN4PBBwc2/ckGgCpm5kc4CtP59GG516vssvireChPQl6a8J4L
i9+m7KcCELYChYmAz3hdgGYHWnhVFnlfrURNGZxNGI0p9C052xIXwR5EgB6BZ4Dd
w+g5glDR2R7/eVuSdWSUClnwr2RSN1NehT6+btv8k7Zn+8aLZSuhuej8lZAHnkHC
w/q/iI18MITgguYTEpOJmQ6aCYCCsWeNqi4l1CQtiYFCys/Q9GhM0RXLK6pxer+9
LvEjNOEXeVKSKlyeS1Od+zVb5ZhqEkrVIEJSSTtQocyWOcWP8DRVA4DZkVYFWelg
vG6WlcVRLv9HhGIKmjjCmzhUpd3jlYgGwO+pBMqLm1fWPaO2H8LHoPXIrDjY2Z6r
rajJkaxM7XqVM/8AAlhltfdcOC0q7LxxF14yVAtv/OKnAEeoDWR/tRXZXlL/vvIq
IlP9sJpCL1FOfYe48CGnC27xyli2CmaDassLtCYEuZiIsv/VGBL/1JtKsprp2XSu
Ysz60CyjqEBphYCkss7jopspK/hcliUPZ3ds7i4nS8IjL5m6C1vXn4PUlGHECgiV
ME7HkUQpbDiw1PGLna6I+6VnaYSAEp8trKn0mQTJbl4iVobacS4Z+TCRop/BGlYE
K4zL7ilCuOLH8ojkyoMPJPdmDPOv2LkSefR6a42mu3Q=
`protect END_PROTECTED
