`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
VN3cZiJB9f6xREOOK65F2lXTPoHZEb7DA/dPdlnnmBuC4hQ7tEG2ug/CRqlzdZCh
9p8TaKoyUG3r3ehAdH44MhBTnQseuNMQP8at3htuOiIWi7zaaYklOBqlorQvydPw
yfa28d5P2yQYooxkuCFru3QI33RqC3SE5jI50r5ZjgMhHuC/rkKyWkJ0Vr0q7aEO
rWHoPAB/xQRbHLNXd+vH1OcJtw+NILtOfMYWjjRMf2AIMpIYxGnTfvKNqgouc5Eh
lP85M7MAtUkvlsidzcW3U3wA0B79usczoS7mB6bGCt2mWKjPtBzQ/0HyWKzkf43T
H25oJh0Sc0jvd9xoa98NYg==
`protect END_PROTECTED
