`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
tPYgb7xueQwo7mWfzSV2D5ORdYLYD1H5V3XogSa3YwxYe49byjsqL+uHRTMXsEtn
sLRI0Dvui7kBUQc/hSmDeYsJyuXdFxmdP9d/ZOEftQBIRDqLzRqA+gU0/7ANh9Fa
dZgCurStOXEdHdMeTb1OsJMMBS7mH0seAf8ENbxXo2vYT9Py23GIGC0uM7mTWUeR
yt60dANo8qKtow2mj1DBC3vk4AuSnityYIFz8uVPKsLhiK9g0oI/0PGKerE9YiWm
RohvOiKwGzzhSb+ABM9Iw8BvW61/iJbNPNo41CX43CIQFIBeho8Oosays8x2a/3r
aCYctrSBv7TlKrsb6qJbs19uyCdnFNZSu2zAq5V6RVNqKxnwqFq4tzUyfvlP9uon
+/PzDeVo/y+ZFqGDXKbzldt/Z+0xJQ8sOW3vda8uIV4c7uYkImFZ/ONkmstnq86k
Imv0MZOlbmNaIeesVUiHCPGxvkB/0IjTImK4Hy9r6E5tkkX59SUB+bRiR1j91B5O
mCXlCeomWjwxgXqYD1xooWMgwqtNAidPH12tcQb48S5rbeqKUEMILgffMB/vRvm1
150busR0t54a3LKpHr4BRuKH9IQeAdrojY+KznZOZtUlqwlOusOQUZdyXkPF93vf
IT4LDp/C2328V1x5Bb2C8q8MXxxAhTY7/U1GdZyL1VDrrWRkPwSIZEbGLxZkcb8R
CNnKcg/t1F7ODrRX9F++qhKFdBPURlRgAig2UvX9XvDKH56rQA2hUZ3LuFEXWymn
khAw1WoGgt4cuiYTlXrGxNKc5QTcBi5HLZlU11sUmQxTWSvivpFWxrIPRVXcLIKP
r+3Mnwf7GVNpDCyZ8pszQ8HvYjJwN+89ajZJWRWbVn5rJWMHJvTsOe2uJsRLi82L
CUVnEftXkDF/T05pqDeKUeWBk/3NQBv+GJ4Ep+c1zRnNsjsotjiVPiRHIh5A8/BY
djMI0CgMrTp7mFXNwIhaWLKnSYmA1D1vpnpsX32O04q4slfe/zaKrJCfYuOGGfOH
0cDTWbLlM5TTnkbRNymWAT6H/5p/3XtibaQob/LX7g24U4Hi1NyHyIVO+aGXhXJA
huntFacxQNj1CDMRaiAadKEQnLVss8oyN03l7bTDE821vi8VjABA+hdrldOjuxvZ
iYCyoMmx+dEZOB+Peu0x4aG0rA1Xe2lrZ8+Mur98jkp/LA3VaBB4NWuqeR0r6eMQ
pSjPvk66H9vmSl+1ixwisZVQubRxS1/MHCWLWf+bBuZ1mT2/0lbkLvKogT9YqmxA
LyFvF15dH00HEOjfMx8ZycQmskRrUrtFZbBe879UM2toNCz8Abcm1c/dqJNjZK2B
TB2F8H0tEoJ2VujsWiS6BjFaUDBfzZPhaH1/2RHi+kkLTrSy94KwQPxlVFpAQflq
Kj7lfSyfbFisRw6m5GGmOmMvdrDPSdgwhlYyrRBFqKlPHUf7vh7A5dzhSIycuFHI
6YuLHs/FDhu12/DoBiNxXbm25gTUoZd0SAIqr8uDFq5+rHJl6b1JmLKFueoTwjzj
6RrsE0H3ZGApYIJ8WRf2pdlTKWazKD3IetnNX2JsSABJ8ze+1Uw3gr87KRN170kP
FkukUx4ztHJllD85rsaIZ5SUlkEG7inQL0fFF4a7xzbQIR/utU31aeFM5V8IRPlo
OzquXUPhSCX5grep6dNtmQxL5f0FjNXEuWy1mxwnB0TclSuWKN97OQouZaILp0rX
bqrKUithp45tZxFb8n37zHvTZT4lTeh3moN5nz54JY9z4tqrwxNVdm/XUF6d8YN4
IEQyEMuXGg9vG2W2Zue3cH6uxz98ZwlH6JWGbMJplqiL4FVD1B6mDRG1yZsJRM58
YtZuxLSEx9wlsW/+cA2CQ5z0tK90vCIdR8OfMEdODWhgUQ1YHBExjimz+DVqnaWz
ZK123NnQ92mPnbkEontjYL0gO+HFR4dmcKP39HGR/IneUkY1Reu4PkiES1hH1xrK
Va/ZpeosaPcUjhbaN0XlAw==
`protect END_PROTECTED
