`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4jUYkdt5VjR8oFbu7ZiLkq0XkbnqZXSJjViEZ+aan56/0w4dT794pzFaiRgvm++n
S8qwUryKduKGlzvm2G4mSxx7LmugGJrl1JEv6iUuFYsEFKcR8i+RCZ3m6lNennXU
JXXpUlfv8QdCBkJDNgVOYxCQWEQuw0S6kBw6V0s8Dx1QM56559JoQPZRJZd8zjdf
vtH9K/+Oqq7VqqBLNnTpAz+5w0Qd3+0zeqh27CqgEhFIV+Z9fXaY63ZFZ/TQITZA
`protect END_PROTECTED
