`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48dN3JIkTXNn+qVfUCFZf+IYqOKpbWIhe69hJENL5yuA
jLvGrtGQA8IsYIt724nZTJhP3N3kaev6s1XJABoDjDAXmA8v4vbRrn0kqZ7N2haC
pu1Op3PKN5XISgytdRTAL+CKFCUBOu8qZyqdLLls8gzE5FlmktDrL66S4XUg0Ctg
pBTabDTklnR8ICJ5O7OrY8PcsQVyTm5rpEWsNxHW4LaqIDsnos1rsmuTpALQNVoh
eZ/M1gzzE3j004t9QCKQJMzveIYje8gdzjxQ78FIbcbnVnOoh30GWUQUVDOSI0RZ
LhX9U+gxTVAjcZoGe/RwJg==
`protect END_PROTECTED
