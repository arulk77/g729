`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAQRzvdXoLOrIRVSO2pFDerKfGRg8wckOTUc+5bJjzxk
b+40LTuPmQKXJsdbvq59Sxrjj4ul1wKxcpUZ2JJUJndhZTUHyV5oDvFNL2LG11Zd
ys9OYNsiOG7z6e9G4eeSlwpmErAwIS+HRUwsp1JXMiirPcjG/I56NDn2U8Oanpmj
FQEep+Sr0wPaRemo9VCnKw8VO12srgyJ+tHLlOmSAJ23Zy5niYcFiSgxOgJbGQcR
XiYMVbRfVG0F6OvLM1Y1seRSZSmcJxNmikEFBydiCq7IIE4tVxRtM2EWwVpxmF5k
W4K6H6V24Eerb4D9ndNP1VyKMeyomNbaiRaKQlrprfjsSNOfzAXolKAV7HDOIRh7
hERiYVyNtVnXGXGPOHKDnbGX5lSP1mUf97Wv+aT51fREEv4pbXKTTqEusl7NhUla
9NiR5Vdmsj7GGUG++9aMbEHZB2qj0ns4xLb3/QRbDT8FsI5O9hiO+2/m4FCihqJj
`protect END_PROTECTED
