`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN5XftQqxJreJQkvz/xdv36MW3N6nJzk8qwGYmtDWJKUq
TYkF/VNZS6YY8X7QoIVRfXLCU3ha9S8GqS/JLkJXgLDUg3wYsEFUlJ0CpsGy6LhD
nqvO3KwTTRSIP62qeqGxPZFBv56C5s+RWZ8ZN6LDzoiRwQqFx/+05YEo9mK5fACr
rgVCwrJL0vdCfLVWnDUFiWqgkrWQNRlZKc1kUutE4+PlbTjOSCJGGWmRWhruBfj4
Tk5mujLe4fiZE9pfRUYL5kqV/J724yqVlTrnMhCqRZ2A19yrOZyrawWuRXUk7eU+
jFqFXKf/1rF11VsrUzcUtvmbBzpCgVgQnP6ZMnOsAC56CbqvClGQsA+Qlm3bsLmC
VN2O1dztdC4kabw7wzgWS7qf0TghHv18Xr8J6F8xAL0inXcN0s/FWWHPsQadjS5G
Sx0U8QUua6qhEt74oRZ0covg3LbdAsFE5IWbZRUwf4om/fKOeF9ynYFux68LNeKm
gHidg4VARREoMD2z+GzKw73QeRNE1etmvfvCJbOJM4XuVgIYnyEAIna7Vvq4Haq/
uXrRnPaJP5Z0vjvtk0qbWe8Z0aJsilTdZRlUEhhgCePjUOuifSGbzFQJ/MAH+hTs
XfqBbYqr4JSKXNm7rI0DSbwuWTHJU6iDWA2fD8qVyVYPEPf39tOUJ+zuDVely5MH
DymvUBwpf4d4ydznx2Va5tWiTzstYZr6VUBz/JYWoizihtW4MslbndU64qoiI0rN
767KdEb0j/xQhjqNS6/V139HTXuLZy9RMsvLq3TDnO/aFxd/phxLRQC+jM3v9Ci1
paCOIXkKb2Jhpfu6xFsPNf/eEsmUEpiAszlr9IANCqdHlkmmqs/qDQlQ6efDZf9E
adFL9Uy27WfSYCvxlds86QzdmCRONAkUHmEXk+9MooLwqjf50PxljQYHhjrg9bLm
fYaIVq7t3HVKYPMewv8XBLuDZm8AfJ4u9kJPVnER0LBlpkKL6hXthtWJxmjS0veJ
9S7sl208LtzgAMgAZSG73i0CqSH4Qa1ikrAf8AtRdWC6AZ4n5l7HECPKZeIdC3U1
/o6IPM0DIZy8S8NxG0i04kPGWI2/3NPdpA20BEhbZ13YcVf7AXs7/lSQiZHbW45K
vn2VBBzEYu2fq1BZ+3v5Cx4av7gBR1bA02Lx7z4ZwgHOobQTyJa8xyeTMsPM1j7Q
mdXPzmM7+AvYefjspPLd4jgxndyjgWdr5V4ngdP48GWrVAn85sj8n1HsWWTFUSE4
ZD245PMnJqf1N/mepk/O4JuNjR6T+CePahJWS3rslNHEgV5BSzhovPn3gMlLfqNO
4rw3zVbMg4tX7zLj1xSGa3iv0Np7nDDYQ4eOib0hDMjkHrh6r2LEowPefXrwPrIy
JWS8tO6aIOJauLc/iDFfhZNKfAcLqmT+DL6uF2R8HKISaeSXPC0GkFtrTbFHyfQv
XgRqpYtcamU2we+k+Bn/CVcme8tcD/zXCDaWncmMWnSL2FfnOFDU0Tbk2hTrOtIH
/Fn/1WmymdhY+gR+JC0K9uVylOHHtrmDSVcOLiyhBy9aEz1L8lEfsiw+fjKAxuf8
kaxUX48J3JjQRU8EX3hIX7oCWlEIY/ZVcGm0PcyCzmNYoUOGvD4Nf3Bqdgie84rs
CYXZbuxyo0g+i2mPOjOq27C/Wya7VzUAUy24XG2cXPBlSvAO6MJ0Zsv+F7HYXdJU
aBC4AIj3oOCR37mrCqaA2iIpbeEyMMLD8/gQENryopSiyli4MiUljlsMe6i5fsra
wWxdY+ld8M65vHZlmWGoMb+X9DfbWPozG3R7ByKR0JI=
`protect END_PROTECTED
