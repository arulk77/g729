`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
q+Me+nrhthd5QkbxkcKqBV2zA/PMsvrtY296MLLSe4TeXY2vXcYtQb1BZr0fUwGq
Hh5BPod8ntDIg1G8sIIJSUTZ/5wOBT2zWCcgZgZhp3CyfRR+YTSZEJ7g8QxjnTo5
d0+eGru38I8VoDVnESDvH37ygI2xNWWoYuhnP0UC0jmxI4jBCr2XeTGX+zuBt6Sz
`protect END_PROTECTED
