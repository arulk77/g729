`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
absgM0bWC51S66L5Etioy2+IGIxpJwW3GxwWwhKC6Dr1jBVcF2bvvAWHyox1l86i
7Xkj1WFLMIF4I2mU9T9R33oEawQ9p1ZrRGEozMYWauBYwGnhFz1iMau3IC04xI3b
e0rP6Fg3mZGOZRce5hupmuGVz70K4O6zlRAAcipO++DFHPo98/6aiGmzweBBIoow
+CjaxDfhiLSYIKRyyR+5afn5S+U7H3dVw2V0clNrQC2O8vzA9MDs578PRsCbiZME
XYliwpHJePeJVGwRjHdKwJh5Hn97KYmcbQlJITss4MpNxQwdD9NT7lY2APJ4BI0+
zHt4WYVtLcqYWfbW5j9MdhWtaCCDD5da6Dw9JUKdPZKGpa4SAFcgE3+VE4HIXKgz
4U159GgmiXvy0A/gzxzVk1O0vXBQY9I3AIZRxD14qR4jeQJXk+NO1WtBqIfKJM5W
/QaxG4InUJNpwUo0qTeAewpsM6OSj7U6WShc4HkHfF0pbfrHvF3bVjIrceFDzFr6
Lq/JkVv7Rj0Oh0joFfo9FzBGDW5YLCn948bdXmp3tXIjAfXc0mZx78u/c1guBm5D
O/K7vXuKu/NdNlN8VKD/IGvUH0gDvKtDVPlLE5HGe4w=
`protect END_PROTECTED
