`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLzGMa6HhMVA2Bbl1gE9KFYc9/FuAE3pBp7/kp+Fuptp
5ACn+AVRak2XQ1lo8XsgjjClBl5lH6z+MrTU+T4MPcmR+0VDIemNKHUINcawVIbP
+jM5mpbsvk99I4pZ+6JAmr2AuXRAwPAs5WNYFLihs3kpASxW9HNXTWmtEHCpNspy
REIQIr7q1pVEYt4obheVVTpki8rAcKdcsywfUnwS+tXFM5bOlbbJmqJ7jl5Ce2s/
/273GfcjuxQYfW5tYy+eYr1uwUxOlCLLZ+NKyj/ltcE4O+2Mrxei5GZAbx4ZekkU
ptjhRB1xKUwcmFQKWUhuu58K2w5Rwk8m//aAzfAIgHOF+gnO35Pu33EPyJJB9AWp
mhrNuCP3nPCwJUW37r8bJHrlET/H/r0ZJt0xMov5A+dzfwMA0QOE5xyZqq+T7QSR
yy+l9PyB+xYTvpDv+gGyck/Xn/cA5CMz+HO6qg54PZ4JySTSQUfoWn9B4r88in2F
KS1haAm3/OzU0iOgf45R7tHLLxTpIbrBqc9yhxwDCirhJjHqOhm7+KM6V4iclFF7
SOkutmZaNoI9TAT5XxGNyA==
`protect END_PROTECTED
