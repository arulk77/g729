`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOW0NFUqDGzgLnmzMlLmA36pET+QkyVCuSDXMkWcrOjZ
m49oX3owgyo8VmPDLPDQ2naQpKgzty/TAMM7Bf5DAn414fxymVoC6x9p8reZoL+p
RbS4C20cCY3d1uAM/g2jXZRP8xeyjs5JPkUGLeTDUK1zGp8QdBakYAa5xVis7yDy
mQJPkjr46XBqvJDKvAK354lDx48BeATvgONXVnHDVjMi4uAl08sx88x55WEB2yHP
SabMNMsisWK7G1c0fOlS59vT8N7GXZyVeQi5VII99aqelfqmKvLy8aQbt878qq2L
GV8nun4DfshKw1Zj8On0tj6cGNsapBpS395CfdcSeSFp65auw7F3T2p7iO7ysR9t
khxiedfZJtlHROMONjrUPuVTEMfPA8sNlHIm5Q2ll0Cx7BbEVtynOapn0aVscx7Z
fGQfowm3ihz5hak80d9+DTZZ7Oma+CXdtKBB4AR2niPothvz/DYU6xWMqgumw1Wa
EStrWPTT70ao/W8LBbdcO5aZGSWTQMipR5COiDjNHXpT/9VLkkivG1Lvn5k0Spyc
uGHNhGp595i2SRGipE9+oG0R3tBGtn8rmVJ0AOOS7GsRLdfGysHViiLJuN9p0CUf
tmvcKxow+X+Io7Rlhh9ooLJ7D6kO+tUkxYPO9WzpaqnKpRAbtAg9gACENWupVw9R
5cuAffXWyVtGwCQkvAaG9cTh23YqOPZ9xU0J6PQd8tO7PEhOyzd2h/RkH6b64GBa
jvNdN+HPuBlMF978IGIk8V9FEsqE2jGdYMCRBH/VLLNfKiWmaT9QQr8Vvm0CZk3j
gldPvhOTijERzWm2LZH63L+aHi+2VN8XqHQ7lWlElzk=
`protect END_PROTECTED
