`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAV6VuFa6KdSSGOBbPXDxV55IXFKv0cuaIXjWum1uXXoQ
ux4JxS6kP/2xYs1rETaRSLoQ0efHg5ysbfYR/5wqTJpL30GzuYwejOHzdgBEKiqN
tUce3C7C+sUnHyyVEs6qobFRnPwR7tih73L00hIDhyrfRFmnydi5ytRjxpL7uRYO
/WrAueuxBz1vq/X0XSB6zswKQeHMrfU7ogNC8cyWLhIRKffUMmGTQsXViOKiWPya
B2kl8+M4dPmiPBKWQ+Ia6hfdjP0u1ytbidH5JJjHhn/N6SyD+WFaL+iMi3Wl41nO
4oPTeDD/t7co1aq6RQAEpw4hTHPPPYoTOO/qedlvOog4eeVFhADwXBu4kfu7RX83
7vglXMNPseoIvuMRb12QITcX5StTgQ/YDpNi7ketIXA5zya7q5Xh6wKFkppwTwbJ
6YcwekJ9sKCiAWRg+SM3t8vBBh4026cb23Dx1cT72UDy+ClI/ChrABv936zFVpdL
Z9MRicN8qTa2ytlKEaR5o9IUgcYi75StwjjcK28V1T59B8GOuoZWCybEZB1bzlBu
78rLOM3c+Il1iq8ntLYG1MD7Tt1PYFAsuVeM6FSJrlVk9NC8ypNSbuIy7SqcGlcs
0xSfiNrLJcxZmEm6ApBHeRa48tXX73pv6XWVZdeM9uECrt+LwhnOwJPzqtJl7tjt
NWT4rWvDTZ2520p4z3pfJM0b08iGvo32m8CoUuvYB0Q6kDRftKCkrPoxTInMZ0j2
Rd/trtJXAtKbIHfB/Nz7HKQoXCJw7MdMDSQ1FwbltiphrfTo/3+4Ist6s/jpEpVV
yFSf7DdcUYNQvMXRrtKRzw==
`protect END_PROTECTED
