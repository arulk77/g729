`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
5Rh/ow5Zvg+X9QWyre+29xrpc6rCuyLGlNHf34WcplIBM5XS6lS8RmWiHRHvG2zc
ZJtJvHe24I0mU8aoEs1XR+xar0qhJdXZWWWWIhHpow0xRev5O7Snw3Ytn4F063Lo
/fpUo+uXsPoTbpbnnk1ijpPyg3+/zHsBh0BxpP1EWC1zSwpVoS7Hesl8eyYLT53F
G4Z0X7bLPTkTHogSkH9hNIQkYcEJp/8d/k72xwbXDihlObzHcAwMMWQxSjJjEb/X
JzicB77Yz08ashDsrZ4ALUKQ5pkUJqg2WwKWBUqb83IQLM5V0LAE2UgdqnXQv5xR
19ielHY4qI7vJaa4SKVJXenctUMSea8l5quCd7vE7mq7rN9d1vX7z55X0iWDK5Sw
eiA9vFROmPMywVTx9Qbvm37nWJ0az6w/Ddi61BqphGw/ooL9nTs9jYLOpvaUGmgo
t7cAyYX3w94M1OxNWjmcHcJMZaKbDsLd+a5lUMBzAKS1+GTEUr1fTjDgPtlXoUrN
1sMKsWkWiOurbqfAfzEjKnvdYLMQjuRbkKWqjRitfx8UFDs04QZQPqpqoBLzGytZ
yA331mShEgOXf6OeFdzyajdRa2NUmp6AlbTwHL7AYGavhbh/1z/DrmrrM06EaJYF
0bIeG6zWOhfBIlRmhEqwjg+hMvqDPumoR7s8gCv15nQAktBqqaf6/W8dDVcZOFZo
cf1Ik+YZdDyvUoNB8Lul/E5+nADx7XbRM1y3npnfJevbYv6PfSbnrezAgg0evoVs
gxbC0sHkgpM71I0S2LwkePKuQ0sgbW5WtljXfv3Li3W0lhPGWK8aCt2KKMG/JvRw
fGz+sd0FK+aI4mamHSEmUz355TuzTSF8X10dTXaoWboSciNTpynJSQOjwryqiL3R
EwpjVUuCHWhuEUHaGHs2vwtywFWYQtSp6YNWshUiZ08shE/gRQtCEUpolKxcSMLo
qIoxznAyxhGfPwlJTVSlHJLOlZNYMQqr7WAxp8L/lRNuwBldBpi/0qUMZ94OxzrP
xZSfyUEeLrw1xMJjdfAUW6CfskgndFimwWlXJnICm3koNWSLr+qi1zpR9FeElDuK
dA+DpVyxPemIqe+YylxWq24t23l3jldUThjr2oK4g6URmk5IGD5r8cTzb31BCu2H
iX0VRy2fxmjlt9M5fnUUhoqsTkCDKeoXya1qybGSkxzIiOj7Y0PepYIhZiiPjJS+
0g3afNMQDjlju2S782hSOUqgcEvo7sEmz71JDEM6N1jB8h6OGXr6pBCR2DMp6Zqt
9sjjIA/1uAGF5s4Yy00paw==
`protect END_PROTECTED
