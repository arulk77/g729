`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN7kSkP8MWgXcWRjmVpWNx8JeQnwCjR3eEtOHwEKzJEy
e16GbXkyv3LUgFvn1Vi0JpCJlFeETnTIkkDOLzbUxTY3rGxnD0x2xm6qM2u9H7+1
QthTdtLLZg8OZjLfYuFfELzCBCToQB/HaIEds0AArHNaWHBY/3M9fCZz5e3FE5xd
GjXvorlsmMLK2ZXKHHm/NulS6lhYgHcHIBAMqhjg947qbUhDwsyZ3RZm9lMhGP8+
4tQwDsT3aJg1X8f0x2svBNdCH+1onfimV6lGbqGhqmuWinzvLQAIk0Cu3E5CTjDX
us9KW/nj7680pxhsstCx3K9dwqj9Lv7GGDYwIqsu4f4hj47GlAeZm4G8O1rm2OL9
QMHDJIwdASyBTJgF1SfsgdByA20XL5PyWkMl964CIdb0SUxghmBUL6GMPJXTEIW4
O8pkNV79/+88x8U2gwTbcaN8tcyC5XE6LWFjjD8cg3dEQ4IgxOoe5M7J/jwSIx4d
QqQSzzP1FPoEGnHPctIGF47dm90F8tpBd7kEKYFjEV3OxDAvgvJvq4QpCVVdiXmJ
PAMaMypPzxqBR0O50QbrCWZfiT0gZ/qYyetlY9xbZP0bIT0409NS31j7NLE/B8Bj
M0gP1/+OM2UYMdyd5ntVRHDs7p7bfjO5QQrgOWgfn7ywizSNo/+1A/rzoeCSlm4d
tdqUvVjEf6HpwjRNvv9XD6BdWgxI9XJL5frQ4bknLPwhh+HVsckkDE4kfbTkLNBW
E/A2l9wORRntR1qcTFLgoEK0KTj2xdTW8fZENypLKkz1nPGhwB/Klyp/J4eBr4jt
NQb33oGR5JAfX4vWCmt+62I6aVmNmMckPMd5GZoA4M06t9dtM9QWOl/i+7aBa6e/
L9x6RtYTJiSYMARL6TV51wsf+hcAOgvWNhEDRxdSPWyq0zi6FpmlIrqyytG+vrvv
VwH7ixJ6EGWaaJxlKmnc21YIGyZhtBAony5PRWZVpPR7YzDxWJbp2RUo1wbl/VDo
a1Vs2rYDsnnXZTSCXI4ri759NOGNLSkdVNGNbU/ERHssC0kJ6PGUOUB9tSWlLG8y
biLfKrmpzIY/R7APMj5ZNOeTLdtvdoreEEsjqedXb8kJ0RDf0gmw5QIPZv58pz9B
ox7IehmazrRaEaxUCBbLHGFS8Tf8yU0IKWLV2bQ+IQUNsqgI/wqSiGUFSaSDbD+l
ezJhZgP/0RbMxx6/xwCn+FxkWBQsxI4mz+cnwEb/s5kHr5HRDWRRdjqOGLEDfJZk
d7pAF+xJfrsVyG0NDmJq5xCJMmJxn/sBeT6GZfD9KhDtNYqRluvgDGd/b72mhZXV
pSCEf54iErRCvHukP9r8YRgkumxVN6Hu0hEa2Z0Q4DAI88gbmJewo2SpV66Rzv/s
7sC4cEgckJEQwrcPXuWeNz0156qoWnhbuWy3IP6Jw+/EwiRPXAf9/n6BwlY4mLu/
zi1cST9TBXlaWjcaVkiy1/XtDEs6eorMZM8hvIrx4XX/b8MUZfarTYxGRbCR7VEg
oqtJTxDECOixj/dzGh53EJamFOY9I7euV7rauN9JF8Jwc4Cn6M4HeAVBakYdlsMy
CEZF2kaxaQ04p8SX1dTGBDsT96EmbyqkOfdt1WlnfSQHvazmLI+QO85Bi0r8Jy8u
9D8e1lRq/XiiBPbdQU/jIo/xviBaeQbM5Fuoa6fskzuxdzjHxfkaZsb7Qe0dSQ8Z
2wTyxDJlkaWhU0IY5Z6WnTFyn68ZBO1KfRcCff5Uwtqi8IJhCgXDPFKDhXQTbW76
PxIhbAUt3OrhZ/85eEIhPQB/1rum7nOJ1eAHYdMWpghknHa1gUkgjXKwWTGQZYxX
uCZtVWjYVfLzmmog3AQKir62Z+cc3BTZUtdIa/YzyvI4lS61kQpkvRStq1Nr3DEf
n7XP9JJINvbfyIXvyLKjXVwMbQ+8u0hOIiWmwEAwz2VwBddLgufzHeLOcTl4Wf6P
XT04zy+su1/PM4TNStg4dOaU2fSU+wp8E/uWtlW/UWavBfpkwP7lelfEPOuqIdYj
mq3BfuswbUUQ6046jmjDdbfp5lgKF8cgqvApiXaoGeRxH+9/uEhscgdEc/dyJBux
W+nZclZQ8wpHfMpCTj+YoCFcTXG8IKn96wWKFwug8C+HZ6SSDbQdzOM0uU1l2PiP
KuTlvrr++4Qf9w3s3pRJfhlXSIFt4/bsj+V7z513HcTGe08aWtU7nP+Kc92zXXCr
p2jrXBsPnM1CXcx7mDt1k47hPYKLwPt6d1xfTOvEbUaJZU1f3EqebxeZhW2/ikjC
KTWUBciZL/vAXaacGqFejv4hVzY+BMiuQ6qKSE6M0F9VEjcbLAyH3mUrJg/1Mp6M
qIUYTuLgAeSNCMQbbYkEJnwR97N25jqujNQq2SZLJgY+FZ6xN+khQrYtkXfvXFPa
E5qPAPDPpOoIDBbB7GFfwVvEyp0Svg/TP5wp1SPEeatEY0RqAGj1lRyRM5nf9NDd
k0LlwGxqk6K2T9aFI710ct2XLDHmfYN7gwCGFiG8CiFKnN9bGwBrz6DCaw/1h78h
9FSVBkTAWSkM42/by+qIwcfkznZi+68qEJb8BkMsmFqU9USUplcycQC2OVGid0mr
Jm6d4Czvx9xSt80NsoldNvawSlMOnrzG1NkYV3dSKDD1bMnRdYCjkq6tLRxjgn+c
n9o+A143VqAQ2J+JWZc5VXuAlNag9/IhYOT8LjXilC4FCrImffVhIH02Re5/m0ly
gq68DMZ4vuAZUX6BaUmBzn6jfN17zjSVacJOlbDKvbX78iy2BYv/zRTKUG5bLap8
2vI4Jo7BNwIzY+j8mxzAhTBgdRlAMAfsXhZVy3gvCOa4nhvErQIr4Rfa22wcp8iu
YiBw7YKJMNMIzhjcSj1ZdpprmWYp9Qis/XWKQwURrynxwxNCuJHq4z74mYx6Gbr8
pTYggxs0EeGqPpiuldJ2Xql5H+nrnsgSlcgFLjin4yXjuBz/ao2dtXdFyCSkkCbc
b5JmCzr34FXkn5fnze2eRUqU7c0n8Ax5zNrbC9HsacZiUgVOz/67B9MZV/61v99j
B55/pJsCI5ghTmxtXxdDvpgS7GNkVqeNB+R3lfRUQw6+2aWC/a0E4IzGC6FD+u4k
70w85UGAGSAkO4SR3f8oQejEc6qJLVJtSQbFG8dXx+NfcuK1nEa5KkgbQNjVnD4h
chkN4ZvS1oPsmJhCi3VoGUkGbyTwmQ+x8Zz4b7WdpwW/IERqV1NQyaMHY/apPiyJ
qrxpXfPvbLIsuIHEFh88F17f4lhNcILyyp2/vS5EgU+Cy8imDIr5MCyMq58IzyfV
+bTvlKi6TE9hJfbkorB7F02VuyOzxvvRzCiAQk3wLZW9Lt9c4ZSACmE+Jzk2S/Cp
AVicp52yRtVbFd2JjP/1w9ohb8M8M6zMkdVT2/5XMKRTHdqVnZksElzB3wyL3iIc
f8yVYhpqRVWI9XdMUvlyl/92W47taDNLFVjPifqFPtn61RzbQPtsIk9yxLjEkJ5o
kYUkbpHXCsUhG5sYrsNwMc+2hA+7a7ORdmD9S7kVxR2S70+TbMB28BTrobuTAPYd
cFM89nJFjMcc6m1bJN4WLfNOlvtIOXLx4w0Dxe6dHWx8ZAYQKZmT/pNdJoQWrJml
hB7LPphiF68myWVKTWh6g9RhTPTaHIvZ1jJ2uhg9IUSrFgdeKyV+vmq/x5YcECIF
1C2alyUxh9bKUkeXVXfL8WFqCmOPWEf6t6LIUydAG4fMTowqU0/TSiiQQjgJz9Ny
IP5z2Os/PBoUa9Skb9BTPYHo3+8LTwvo4RJM1iWrQZcw815HgcHr9ASRP+Q0i2At
izcq1g961roUwxpXrBa/eeKKDH8TmMmQlcCw2WDbrBECDCQ0ptg3BmhIFQNSYucQ
707/oX7f/tUshGEF3Y48DL6XOI15sY4Vpf/5Fj2UnrqoY+5HKbRB0Qjr82/Dq7qb
GCaWLWMEwXeXL2sX7m6H48+yc5ThNk+/hF++/0IWLtC1seLYBppqSFLKUh64FjEZ
UHLUQMst1vDoLxZ72FQXqhvExnSdY4/L2ETMpoKwiHGacErQnKcrWVA/fbLUTrTr
OjbJToHYCCqjzgLd7sl7Xm0EJMPJstRi8WTNQkJHs/0ChXjA89XwOLNXE5IXNePu
d07RsiLNTM3ycvt9haq4xVb1qbBDUTQYM8noQlJ5HQjXA6y5MU3dQLItb1N0chId
jHWHfSMTQajoddDwsS5e5MdDaeKWUrQehwRhxnR9hWdLxHZCqYX5ckLOcG9WaiX6
tK6MNn1/GlMGPDoQM4iuzqkw7k82xQQdmMbw6BJewtj30eqGY9UFpm7Bv9Rq8KOG
nDQ01mPdouTsNvvjtXdDxUnikXyYNm5R8wzpJioEMTQQtAa3HDNVOXpXrD4WlHyy
USjKUaIDZvVwhjwaBgRNjsguCmZWZ+U76wdOv+OfRjFNbkCrlDna4gyKOXZFrlrN
TI6P0IyuZ12sA9O94n38TalJdPW3N6qCm6zVE5nqRoc0AdRtYqAzra0Abxq05zdE
SHbKhSCqgXNLuQyK83UhAQUIqO5CFaRKjLL/P4QFs/l/HAyUOQEM08I8EJ5o3ncP
f8JbkFEpxgz56U9WCNX/wJbvGykU5luoLxwHq8Lh9VgBD7DLqIQF12SINN4yNn9F
tTOZDxk/HoXAzoeRlc8DN80uEqdZJQQwtS3rH+9WACulA++rVSPdRW3ntJjiKWp4
85hlm5Xt+uINpIlxfb4N5wxlGkuSqGg7IqOGu0xTmd/YrxsYlD1vLM0f4OszEbCF
0vTp1pJkBWWyiM/fN11lSz8Xl7mmFDxgmQg4jCM8diKtk6kDtZUC5mti4hWnP4Hx
b6Xd1U+uninsvfGRmCmvnLV4m8228IZ/GU7blprkvDdbCwVtJSEzAell363hqpOX
nOUTAqbLmsPIx1Oz4z0f8udIBttCqStf7XyNXhQHFU3PYMq6SU0HPp8i43P5b4kY
y23TM84au0sLyuhMd5gBLv0NJlL+BYvj3aBZuKFRB/P0qKB3v/hHdNWmS5qqh2Zw
OwvmoIXhmykiki9MPtORGrd344h7tt1TYUOZfCpTGKXwF+teDkhNTdNmcBpL2Q2v
YpMUqMinbfDuxxzb2WwUnIQ+khywNDId1T/9DiT9tfkWz0bKyL3QWMBmNjdO1ULa
TN9fykuny2p8rNwhmcoymKaeVi41YXEw1sfxdG5dF6h43V7W10+Bx20pQjEInRO4
GUIDqc1GO6zmv7IP82f1flwGpuJ2+D+7YOuv7C2NT7bz7VA2oSezl+M8Vt/2jb5a
a4K3UT6LTcwRUhT6YKlu8nHXl7cOsry7fj0gVXut2SIWEeVNeW6EosHvn7BfVtVi
wb8vD2K5zn7F3qvGjnkRTMhSC0Ehgnjaz2VBykKV7ietsZgvLoF2zeFSG4lGjTlI
zhWJLqM5JLnyF2YlpAUm+HAo4Z8VLTNGU6ImcnTSPHXGcwNvXWm6/QTBLVmq3Lar
kR4T/mYpfqjan459maRRXw/2BJlAI6eBcZ2t5m/e+eXBRplIum342eh71MTJ4Mi+
MVSnkiAKqi77u8bGYhwTWcNR3AY8mmYqeuqN1sLZ8mBeGIsJR8CQPQYgmZ1nD61T
oBBcyjvI1gtK57cNDzbNn1kFmLp7gs00GZB6VTrC50w7ARzM4xx+nDErvVBWTMY6
SHODdm6nDuZ7yz8GMN/5HEW7pwnJfr0TKi8NgaResDG2I2QWhoYvd/gpnvW37vR4
RFFhPB2YudZRYV9hhrkqFS8c5KCXd2WUwpF/SFuumhUd4hXPtlADydIfzk7CRdm3
zvKyUmWwkhKHTsEEndyDD7GsEV6MDYr5lFx6wDYzRPh/mdAcghCum002hKEj0VFp
L+3fN1BAOYyw8yHHPVdLi/hEEgOuXWWVG4Ehd4clh/vq8awAJRF6VyHMXIfiHdWL
saflo3WJFzWfzrGvxL7wPeshwTHe6fSCBboKIP3WmlUuxYvXCdSHC3qVwC5ScVaG
Ix/sMCDxrzQlJKqGTfbYCIbnr/sm2QpMV8IFT+dnWPJCLNjh0J7IYvTRwfyb+O8H
ue/0Zw6UAKC4cG41Fg8cyqeIqoF1QRE0tFhItNIDubwdhi9yP9MJMyS/6RBWstZR
gyV8JGXMouV5h28a49Qf10+QEeKb7TANhA7adpksm+Qr3/TYetjHDah4uOZvIYCt
La1iAop1LAv+B9M6OZ5Y6HYxPYEA3r3p+gJoauWrtbhEUFsASlUKNBaEyoRStxnx
rM4CuW1jieLqNvWMIJEQSN0mXMrsu5KFFYRGIwtsP61U1ll03Tl9R0pytW2xqsqb
DRNXUvzUgtSbo61cRmb2YKOUE32F7FP3QL2WocAyXSrML5riIstMm53Rj0lDywjh
yvdHvxuXhM4+U2TXNJ/9dmckhPc8zh0/929xnoK1yrp3LBVrDW8zj9MizW5C26ba
tIN1Jx1DMq9kFotEUZjW+ku2/2cC3zU5HtbiZy4RndzCV7MqlsouEhO1EgvBk40M
9Jo+TL9+xSY2K9xhzLG1sSfBYqz/8V01qa8rA/zMCbBqRRsFtZMA871ZA8r9DUR7
7udCDuOvxpRud7rddXpNvqUFW8NnbqOL8FnH/tQda2NE+9DR4QLTnq+4vySuSTT0
L5kZWnYyyvpr550yWE3qXJxrmD5AvVZKusHCxEaeaH315Koim83zkspFN+6GoDlq
mwufsYKRaEsdKZZkCppt2N2sUbCe1+DMKlW70trRUy1NAYTEATvv5SSvVuR5flYY
mHVuqhd2lGEy7ONvKl+phrjdojkiPuP3aWtRQ2BidygtjBv7KBIrItV9RFLrR9At
7/icVGv+0KwM/yPhyEcWtBNdsgkyirJK6tpO3BQXUuEOkb05wnAlr1MY2NA2xmMH
UsPzSe+uZ229APmxddxgC5B5La7mj/WsJhED1zdhxEFRsAKdg2bx3YxzfTISre1P
z+x4nhG7b6C2H/GcxJlvhz6RGz/QkDF0b0vLSRSRA5zZUUAioKwr0Gd5YpKWw+Eq
efwpqDRtYnHyrnIxam6qlRc9ZkHpP9d2FogfdTkIEw5lfKTu5B/q6vv15wm1FeQj
qBZjUsfznqrzCry2lcWMykjVqYFn4I8mcBF7l44IfRYwFjFYQFt04NrlKiF7TdNM
M1xR9r4GG7L1n2QsHZoM8tQ6pKC1QSyEBBT1SdqLA4y98142S8yDMpVeq3H+2TbI
N4DfPVN6wHZbNOHDayBNcwL/3BRvywk26Lqcmjq3v/G1tf/MCBHRSmQKLlEgy75Q
+Idf8QHZnrdNVQrzR249RNMmuMV8yQ+YeBl1/E0z1izJ4+btm8xh6jSrzmlNkQtq
cn2ee8ZzjAvNIeu6P1khuXo7c+U53dqWYAAoBc9bcJj5O5W5qk5gFr3mM4bbuHg4
P+V53LuOH+ItNahklKPDiaskBbrORUoulKwpJbFU/7JCt8Ao1omLHxFydLHcJZM/
UH9RdLsS1rDxl40OXWkdKcJBRFjv6cxqCkvs8CjxftQHCw0j6scXw57d7BvVXoCx
EoODpJoxq7jbmRXJ2oVDKSxRC8uW32Q4z8ddWqFGy+Z/F74xr9S1ZvRA0EhiAANN
9m5/fblJImH3rrTBEusTKSpy0kCJhCVgTDKX4pkEW6cEqKrH+JMZ6STnq/y+OApG
BmFovaXjmXPiRBmh7q74rAxrpeRdORa97LP+pmNuIZeymTCNxI1k4k8m3FMdUXlX
xd34YujHlqhHeow5KOLQ69ylykurqU4BU2fcsMn7GYDELm4n7kDZKGDP9M2ythCs
bHTtJl73lXl06bMuCYCcX9k4EfjIVyek2DgRMORw+ju3XYN/NU7y3yWu4Cx6vh5M
qagvugiTLPhhp/Lbk1yh+l4mH+zuTJPDMXf9fQyEsNkGuE3clKyn3VNdUtS/2fAI
vs23KAiq6Xat9Q3dOrIcclFMaez+ts4Axedgfxui8H+ourneWVOAHnjt1UHoHF/x
Bc0+lpOZeKfAQplvwrRl9ChW5ygHnkDkNnAJ+RRhmul2Qia59JFu4PHQ527bcPFB
z/L6qlmtKZRLZAfREkb72Hj3mjG/fu9kDOVCPnCDnQxkeoxM+PgaUQ3DKMLf065E
f/sdWLpyhDZvxLi3Cpo8QjeCbdwGNvYnB1RsmLZu+FPTskUe5s4O95o3iyG2+ihr
ru0uHl9rHrepYjiDfiUGWUtUKh8nrFAqfwNmhpWC3xE6+YmQlQDnw271D6jTVqbh
vTqaHFjg6YmfhooShU57JB1oBdExUrEBuck2LaYDlPW0R1kEM3srVEnmfrIs5NaC
O9GUYoEnJaC8dkHtet80mSowHo5JyAJ9HrM7CQav8m4VYmorV8PELc9zEAzBv5wg
xWbrcR94T3GlQ2futljEjbILkvo0W4lUWSSkuor2Nn/sK6L4nvio94v9Q7T++JgQ
v3y+sBphBzgOMzjlfEOd0fpfbwAAYaO4jimADjq+Fvd4LFI7Mnkk77kHvl7FgDbi
wFAprNiViygyaCg03x96+00+cvxzlX9LzfBJLQIkezi9Hi42pD5EikvnCKBwi0H7
8QRL/Pm49QGsShswnZoVQURrtH95lybe37aI0ROgSXfDPCy0Nuw091N+bZWxcvvd
qAe9xoczQNhkczkUEeM1LsWG4sDQD6NUaenpcDouwqz2oiFa6tp83ei2RsX/0sD4
JLuucAAI0F4cSA2s8RPn4vLJ3NuF+hYXVKFKYDEfPpUqYjbF/82DdWCUI9tXqf+5
HqlJpW8OZGd+E65lCYCyhAhQDkHxc7KNLh0LDl/XdtITRizya//uNx15YXjtgV89
eZblosM8ijAWGILI4Iuk4lNVPNZ2USBKftktm7Ezg3UwEIVFOXg6BoIITTu4Baqz
Z0hP0873Sg0ez+tBGFHUYxTbeiv2NDvInaDKhaKl09fPR+IuLw30weVXD1QBcgsa
eEtLBqcj6rWlmeiveMOanIArwIYyYhxiDMq+Ig1lYcGmP14fx6aCuCVefKq28XwC
NrALpeQsMIrpttA178Vk8+Vw149TbceOrynO6ChRXnO1zQP+i/aOIggQ3CTRAZM9
XVmsMniIuUVJ+7+am2H0eBIgGxd/dnnV4W+BDPRo3KQQ2QnCXPF35tdirTHa5rTu
y8MiWmR28w7yJkPwHDQ9M1VBUqTy9rsTSDxGf7mwjNF4CaHxdQuqfpw590tePfDk
55YbR1UQE3l4ca8g6yHpMaMVViBY2OBorpBAvKop0CHDIugo7NVDFjcUPp+1xQI4
h8OzhZ/kyU95oCphVhCUb91NnlJ3OsR9XFmTEUV4kpJv2Q1FIlojLRn2DwVQ84XG
eO0KCVgbTmAgdvQoXSkBQMdyo3Per+cuByN6PPaltErgEmRBS5/8eyOwpoa6xD58
zQ0EW6C62rthHSJMrNzelgpSZs+LSSornz+/uP9BWQrSSo9zLktF98AvNwWHN6rV
PrvCL7Dvvs1OS9jTjcxbaFSTH2CDvEY0VHxuX/O964SGpX9xgfchT/51UzRuyJ1K
U7JzLsCLhhfka+8un0Ja3mGEqaGTPntE723fEMTTixYM6Y8z0EBBZ3dJ4OngOZ/w
lOJQWzSPvKHj16q/tFrEtW45ogA8e84ePHTMEep0oRw0ztDSNCKd+L6J/dCJxRMS
Bxsa0gZ2GjA3WS2As9C90fYiwhQEX1MOPBvu36YYhAtKguKeZO/X/Tu+147rk3Sq
6aB/AZ7UJbxt4HU7zh707Gqm+Xdt8QHxzPsGH7uWOzBcUcZHQoX0Ww+Ol/kenz/i
95m1f+So4PT3H57E5aVz8V7wKS31bYEGyWF0279W3H9RF14L31cVBELMUX83gKQe
8OOt9sXMITmwZCJvdtcBdF9YTCK6dE+zE10jPnS7tAA9+xyLva6bk4AzR/L6wE9W
gg8Mw4iIkG7ilq+IPaCdm0l4MQB9DG46IB5WgXJkJokAS7Jg3/mOzCmbktwmYUlF
Pbgsai6OIz8ZeoZFFmtHpu1NjWapzl5jsIrzq8tuVmWWYYtoZfNrgA0QoD9wf0nN
yqqwCDkIolFe84a4kyZaukGkatSNzHxjdbsqySqpr8PAXtN/yDk4U4gpiYBH2sbu
W3m8jwWu2t5FDbhhM2lUPjcU1f5SG1MpQxiUDMCsk7VgMw/CAeOgxbK3IfvSs25t
t9+eKzf9ImOr6AuSkA34kynPtGsFqlwmfKriNXMH5oeqgRY6RdT4GA8vQUhVD9SW
PvxIrC1SH+FoYyH+WPOmhETRXa6vINPhOwsriy6T5kOskZddDlhqpHtkUIg4Hd/l
SHOpp9hjTMzQnRQ4cTkiNeEZ5Lf+5tAnSkU6mr2bq8ugEt+gTdD6Z34ESd9Qpu9B
IxVvVh+ytB6PFuJO7wbng67CzfYg0JuvTEdrx4KA9oAl2ZNWpPfDa3nJC++kL4hx
nTQIefvOw9iSrvrbljjyH70jnFMfmqWhNJU/Z4384xEMI6IkTKxoXotbaNe+kHPq
Favb++Ji5Bnh/n0SugnhBRqmN2V6XrzA7z+xfI6/XCuAVIuVEBUxeOS4hCxwG8yw
WHrCkOXh2bL9hPSOpoCZPnugRpi4Yluahm1BBPdOunj9kWW4nK7HamdqjrU7LEGI
RXlCvwPXAwiPeTd0QPCbTS0xfdUWNZWDD0x7DT6SX4f1YJkbEc81gyB9K/anHygs
GW2EOGeZlV0K1PXHakc5tJBkKWw+EdvEP+Txbe8+Xk5LQRbnBEyvQV1qzG5nHKG7
OGPvPMIAGcjCgfiA1g4BW1VY1o50pfjCZo5qRD86Ha3+Y5Dz8zVF8bObP/2tJxfW
ivz0Yocl9fMn/U6Rh4i3XEjzHabut+OhXAjSy4x8GbU4TOXkBVWisRxgbUdUHV0S
+6vxvV+4au+tL6DsKBb3j1uKSCSpNC6W6M6BPwqD2ahWbgkBjFAV+IECwPBdLjPA
OmOCRYAd3mDOVMahljv9SvwYLveaFsB5+Lb5U4znM6l4ZbvLlNIQqu6BVNnzDiz8
iTfn2Df9NTHBxZfF1VmonaUbTS9TZ6dZJPKZa1/8CKkn6ykrkpNKelrdJmdMNS35
khpFcaKhzYi3uwztBn9Kn2JXZZYqwUsZ/RdBmFqKs0jdy9dUaYB/6kuEO5mojTJm
TxVuGwDiPkfIkXxtRedx16ofOeeki/GjQ7uXaY1FmxYeSiGwfKU42rID7LOB91wT
Mygq5xge3YjNz0lge+zJZySsReqSND6KF5+YCp6tnzg7//BuDFfidcmPXzwTLqYr
CuPz6A6N4B+tIcjU32yQAlrcQJEm8ljLNCIw1h/7XemAMjhMHaXPoxQntAGn/rBz
a45VVqVyWKWzm8IjoQdgcNEOVB6lnwkirDvYlhqAHAbNxq9ykzoDeILRmaLc6io4
OgUEZmlVhEij+Waa/QkZo8aFP76uSClS0q/7qpY7M7CmBYRcAltLXbLWLnIU9+Sc
2gARHf3CceHz2fqhuhZbr67vhgQIXYfVR8ZRpvNczABASoN8bE4umKFB3gTqErtl
Bv29Bjn4rOiWvYcIl57UxoS8FxrD5BHtgwTAdea5zRkxQlIWqhLVbf1LTKWs/fUf
f2k4F/fpCUgS+uOV8RFS5/Qb5wY7eURLLqHQqOOFIvDacbSW0SPCS/dpYdrnFNKt
AjC8fib8pFyA14zhdKdhpuMhNK6dy/6kSnM9savMog/8Ojuk9GyNa9CtonU/lLaf
xacxWLRMka1RnUrKMWXmGZGFQm+P9I7Oo2TKW72onSpO4422m/PgEnRfw9GQpqo/
rO4XSERTVWLgQd55r8zXB+UFYbB6Nl6CEF1uDOmTRE4pN5peyxSfcmL2L0ZSHTHh
1zsJA7qZmLpQT0S68HtTZ2+mgW2/L8fUe4Sy+ArIGvrpKb6RpDcXCtUfU6iUwyAO
u/2cJQj1P7hS37ar9aJyk2F2EK9d5DVJHCYySFPSK3KM073XK6nCBrdVJzu/xlf7
pXoRa/GCneuJAZhshWKWilHIqqr9YZPUTMFzto8bfuplEWDcd7AHP065zxhCFER4
vWQF81vio1dcfPLTmMoTr3a17iR9z3MM5/cyoOS5IlrMEKgm4tiCjv5DOLN37Mri
Rv80bcIaw1krzt0c6d3NSw0JBz49v3sKuZ/h6FMflbFfWcT9l/qq29yZ9QR7KwNv
+9UaFJEJBrC+v5HsOltV6U8H75OVdoLgGq+MT2ui+f2KCFrRSUtkqoV43PWlwaVY
Svc4aaKI21ESbAYKkwsNuGr6IgVBu/M3fQnf+PXHg4LXwa0L7bAEtvoo8nS60DdL
hXlCfQBmLLsiHLG78nsevRMrrC0YwvtIdhM0jHsbNyln5evmey7VSSIyOV/x7tdz
fuJVrCI9Bc9XRZhyLjLPjqh6X+AMXf2Wuf63c1BO99qLc7wDOh2XwHmNK05vVGE+
ofYft9xmThY8BtA1Hy9dqVjCReJ1D4KDECEaHkzstMeey2OHP2tlYUpx1DjE9gIP
hX1XRC7ofqNuR3xVLME0HjVHtU0H2pddw4F5qufDLhwwDUuUMLbr351U6MY7uSt2
IBDdN5RAn0QzmsJBWSqUYg4hvK6bWEFJG3mJlfK73PekeVTasTwOaZZ14oFAmFfP
YJ/ej+gm0x3uROZTgZUIoBhq9N4XDNhPDNZbATOKX3rhg5i6jEC0Gy5JLs6rWsFA
dU74eiAbpUHZMEgFEL1/vLZBb4kgJQXvImkLzGpO9JrGEwNQJh4KI7U/DKrHN7ih
sLV4wS6YaewgArpUanZ8tXgjWjhiHrWo/NXzSrhsl8ryu8MuU2i+Yd3zAzjyJPW+
Y8u75DOgs6SxWtXYSoHJgUB6kw+MKMZeU27qHgnSrGjzL03Xei5jvUPJ+fGu/wbe
K8OwdEQH2pQvtTwd8fDCXowh9UacP/1PWnsakW8sYNSMr9R8T2ZvkG7qjm3w/4X+
sNNF7oi3cjGltbOZ3DaivtXMJt4G9rN34iF422HESaSe/BircbazzHtK00aLySVR
faZvhsyJB4wnhy++q8K5ye9D2GYsEdIR+CXpXjElQ5KL2NwQPWIuPwPyQghouWFS
j8Kgx3Yrybx22CaATXioSRrqb5RIYiZ9xOw+4OS4KXmQFV8zBlZwM+MZg2mB0k+l
Hhm0qfQXJolvqNKf1mcxRa5f+889o0I6w3+edJjk0CHJ01bSZXhb0xwjy7W3QAND
3VBayuiRUSVbKLjV3I3PECqCdJ1tRuUQz9YhlH+GR4XbFoe7/dp1YXAE9+KI7kQx
doF37Isk8C0fLdO7sAtN6Q==
`protect END_PROTECTED
