`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1adCdxlakQnoGHC6+keryNKaxc0gYcIiZlwiK20NeKQOv
82qLROREwIHO8xY2gfvKb7hWUVsjKlB8WXI2neBd7xvRfasNI2LCQUhcAePz0l+e
yOobMES+kXErnnqiWRSs6JbjsDlp5qiCvQjRuR/mQBfJxFgt1cKUJ4cWYR7X3YDW
pHWhmlb06Kz0JOLIe6waceaKJaNwvmS5F7O6SuLbYmR+4IJgj95HmlhyQUo6gVkU
a7bQrW43pryiGkb3JSnxYF7MQdeh/VC1OGrY4/Zd/t8fQCitpxCbjsIQzE1X31fp
KnWDOv2Omg9Nl31X+5nxDeYHg5UiI48vuAYuUrT893EzXCw5/OYBs8+3WF3gmtC4
Jf6h+BpsCC64ULE0yTKNFyj1j/gqdpAMSLxVQmWM5EDUjMM52mLPfqfscsWrRKp6
E+ZgtycfydIQmurZ8YG/RDwqtdEvj5JORFSDFQ+T4rlV7LbucZ2zVxlnZ6a8EN07
dar8TilumTG1lwuxVPmD1uoNYFfX8LJs//95JatbTKHwsQ/cLVDhK9icSNImB8pw
avi/PuARklfgBYi8Xr9QjuW7ak+6Tvu2FbfS7hT0Ddl2ex0HsUkYHdvwb61wZxEw
gzkUxULZJfBCtarGRZYyPfrmFMULEYoIT2PZVIqImpycur9ZzU1aliecH+4QFFhQ
`protect END_PROTECTED
