`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePPHJZM66FdIWNqp5CgTAyvayfMeLEBprTsbx0W9p2YN
/F+HOcSQkC3N75rKi2eSR7GnMt5SKSVxVk1XCdn9o1oYd5rWC6kwLVk/ln0zHto5
S2QAEsUB7ZZUT5Aduv1d2ECDzJC8X2eruannHVvc8c5ff6596r2iEVbIAfV5SM/0
HO8S9Sw4I3llHS2/hFQtRluEC5kmqbnTxMcgtal1A6JMdJkunEB6HCESLs4m9D2b
yJRdydieJ+ju3ojM6rPhVmPFlrFHf6kAfqEzWL1NWy2ZhGddAy7lsPdyloREru9v
4Q5HCcpig24azqTaTBmnwE4Tw1pbjowhiPq/vitgXgUQbn8Ubgl1a8DAr2FmsSZo
SRV3zk5DVoXN7TKCrRIl0p8U++xdeXSeiqMpZcusewLEvv4BR0Ix5TFzQK347bef
MWcQ10snXbJrY1+PL70YHn/yUlI7L7+ZHOI9S/ZKPV7+jpflZNRqXdPg/wCmOpU9
PbZ6rK3FC8ZVQQEbdLUIavdou2qe4ez+YGv2812BbsTp4d2mJakD4qPPzAQmmBPT
RSaI28wLHZaHtlf8tddm6g02zF6bcOfIxX3x80cpYFd5wA2l/DSEIZXnlYuUFHPF
I6HGqzKpNzv71Ww0gZVVD7nB40NiWe9ekcT1h7qLowSkV02OIig10u9NU2iScjdB
L1FtVDeRR9MTrQ4KEHIATxK9sTRkHFj6aDv8xWQx7NpVzSqqW/DFI0WnrrUUkRqW
iRzMzHeTSEWEM8qhVlyDcAes8AMhVijXqAdUhkC/U4ADe8OBbh9FFRYWRLtnui1f
CI9rITosWuo32Q8LgHPXNeD9r2o4GYbHx1w/iGM0B+J3JB14kfaUuP51fpBDa7GI
imV/cFPvNOzCPp5ZI1a6dBllpyiPV9cAyXowF+HME/IevXQ/SlyE4LwHeHDmFl9P
7rPo11sff5aDVk54rAfHO+EtGJ6LeF9qQX2vIXpDefBXtvswj0oTvsIUur66s/Ug
iz5o1gLeSGH82kGOGJL+4iIpBozGyPGMdd9l20sSYFV87tCWvkqgrf8IwuA/flTu
JA7XN+VIOfysVSCbX4OFPZqVL+QHnBLr6F+0UfjK+W0JJuUiaQ7PkWJCkAC/xjiJ
XWShZ3/SLNbkbxgYJGIzwzXwd22AWugZkOruav1ljtZGlByzubD6OFnD4jOWYcF6
SKJq2Xda8V/GEb/gTYAwMi1IjFi/UZwW7KuOtTLIMumtSopBgmukmT2DBdy91nlm
tTwy+xskNn5IP5wJ+m9Oq8sPpMzFQGbK1Wo0sla61jTw9JV+Z0ZeTefPLZd9LBcK
Y2zxudkxLZnao2VN9sq+bjuukskAzDlXXPhmdVIib6hwIe2PZRw/Ch4G74dA8nLx
MBo5fd794Ta2XIUsNY62UuKcJbGB/UZzj7doQm7Nkgf52cU2CnWpPlh/7/l7Lzjn
sVIcISFhlnwpaR6hF+6Dl/qRkkpbXiE9Ca/nOjPe7jxh6W+hizY1r+Vl29D1Nm34
IZWyKfMTbhtZBiC/ofLFLexmAW17QrQWpLoBXmEtbzOVthBRshAL0/wFeVvZARda
SVCQjj8a3lCwalazdXCuhRVLQWowNtgLNTSsHLhqF9Bb3cdrsltrXsm5u16KJesi
bgPeuIEZV0akeEQ4jlpt3Ucce8lWs6SMR2LWBEJq2RxTfgyGvip3y1JVF3QytJS/
9tCLdG51IUSUuKSeGPzvdDiWnrSvQTbK76QoaRuyjW9ETWsy0oUj/Y2mz1HUR7ok
cM6LE5M6UUPK7N154j3t6tClPugqYamN51ByhGJMwRaDRRc63PjaWNRE6qyT8R6R
nbY2Eg2lwSeQgESZAXedVihRab1GfitBT8YZwiBCP99LjDPtcEV3hkfsPZH8gl2K
Fa1lreY9n1k+zv2E12/vtIBWKxks4IXZDVy0vlgbhq4ySb8Rf2VC0jLsvzcrpu5A
o622b1V8NEOXbUYog3UM+XN3Tqzm8tfGgUeP3ALouUbPkYrbNDmtTFfBEVZJnNkE
oqs7JncUNj0hJW6z7NJhAQ18iT9wHiAAqUJLVAeEcxDLZmweNAyC49BxkUQqeMED
jBa1wToOo8mNrSvLn3Ljx2d4BK0XpIFj9H8LwE4d+8/0/CTBskjFgsFFyCSq7gX7
2c4T8LTpz1QFJt1BFUBmDhV6VAjozixa47JstVB9FpDW3UGUBXYZCwQgpmye+BKU
Hl1GtjdbjqfGrjwHyy/U/dneYD4Gc3MNLQPeiA0IHIgoyNqZQaXM0gm+QkAMkrUA
kvhKjRm1Nt8u4gsAglaBes0L+2+Esi1XsDGs9uRx9+uCBkbvY91Zy+9phAQ+pkGG
mSb+gu5pXMfsbW1Fg8vkZ/0ghwuhAWSz7DF2oES7ow6/3Cdbz8BjEFVy59ObXFko
8rQPT91PhBT3j4c8VaA6Vdx656bi/O34R5fz98KnovJH1WUcXCCMSV1mUXAYdFpV
CYe10pe25vDlSo2u5A0btf81cZWwUQcsQJXuy6i0YICvcGqi0MpXQ+X5C5eN+ulm
KZyDKjMP4SP2qGcL0mz2ZxfRGWEMonYG2VmkJMSaY3O5RSBlKAWBJOmRV+WvVt9k
YD/YXq6N+yk9lR3/yF+Kh8jwlPdSSU33oYpqpU6h6lQ=
`protect END_PROTECTED
