`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ziklh5axPXh3LbPFDzuwHQIJe9cGh6AlQxsB9xnVd0/Qdyix4kCP0/5uKQ0VuFHa
sDfduQUemtuAwW3gZuWVg5Q9FtZD1uNxPfOQkruU1In8AU0izQXkIAPjfo1N2fXF
YInETlbkrYa5aKSu8SlMsbwwiCyqlaTeiQ+gxmvJYkMgttMXeloDLfGhod6HBLIW
/ZsGlIDvby8WRiJ1FJUtd2Vval+o6+jIwvqFdrqqZLVvpAPtaVyjNMJUL5HpJ9EK
JvzVU60CpHQS+iMH/tm1N3T0x+0yQD/WrU9rkzlRRpHf+m0tQmEKmpuKYDukAQ+z
U5dJjaNGDYe7u3ViUoKQU7ptLmstuAWoxsuHvWAaNyk=
`protect END_PROTECTED
