`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
b5DwubE6Jls31lciL9lS8cEfXT7aQkNp0ZIX/R2bfTckebWmi1UtQrYLvNXJ4VN2
Gq/jPqo5Z4kGN8CLaQNUT2ujRIK2kXfZC8FaQtm5kq0YQnkBl/7PS7HZGbPuaVIL
e+1+FSCZgw7HMKJq/vFS819Mpdtfzodwi1bzyhiTEuWBL05JVIbhdNYzmUFnXoAw
T/JyDtK7p+ZZRpQ6KvY2H0ReTXAsaBoPd+NlNzgo8wguCsJ5NwGyKGIA3lTJ50u7
9BT7belGFw1UmDUK3Tb8hpB/5VL39r/pjybRQNhYoxH8BroCKAG/27Yok05K/7UO
d07w0DyeuomGp1J6wk9cTGqkEayqkxeKWqGvnKlZ088=
`protect END_PROTECTED
