`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
5ppREoe448u1KAlSfeSBR1y3PMtKJNnMzji0oLH6ltgTKxmg2ZLXh3pSGjwlXqPY
WX4TH1inyDrxqt9QrcyOY39BxtzlplWo/uHYEpNhrWZKcsvPNUvH5GrPSCLao9l2
MQuVdWQasqbdVycNGatqnfDVyIDZzcXDCpHQOstlrPOjHwWvp4Ip5oNaIWRBD8RC
+3+X7N0Cb9MU6fHsFxz4SN3KaGHHGtIeMPm709v+tX4MNmXDm3LYiYFkpkJd9Kao
Sm/fMYqWY0bGYpsVEPZTPuObiBsmSTA2N3juRLFLLImh29muZYR00zNO0eT90MPF
`protect END_PROTECTED
