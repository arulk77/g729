`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN1uZcgaOHVEDKb221M3QS75l/i5mInCXhEtU8ACpfYZ
Di5eXPUp6liAx98/2vsaSWDAqKio/8jRxHwzQe1Z2UtpChcb/BShXzbce/KNVsws
7ye0s9MLt66yU+VYsEfmahv3SD9HQSlyStYTLHL2PQV/YnGcYhvyjinskdSvSKzK
yOWVY7KU4Ak1C5scPdUSdhhwuKgKkgxObveh7/pNFD1sCTw/93qmrR/NzpCGBVE3
mrz5uh/F0BSUgo8l9DJRJxF88P5+DaUfkWFQTR+jUcEVINDLeSOUjGvcg4Os6Sp9
aV49+4PQGSdJRiufEmVlX5XAqZZo6eXyImMfjmw8rjlbr9IMIp8zuhcH4UQXQjkT
FnYswkEWGfEadiWsSXMU1yz2ImBSwqaytD92FmE0Sn2yzN1qO6v3C56a6v6+E3KX
O5crpQYpFqysqHzKNPM4vewBPl1e2vkbt9WPpiuuOjOGJmLMgEa3eyhg0M6qqSDW
556dzqrBkCmONHR7ztrJ1s2r7zskR4ZzyzZBoXxn4Apna19jy78HDo2TA/AaEUn3
uq3MZU93uSWoUEMo0Vm6IynYaVO8gNHVwvlX34V2lqTToF2Oz8t0VHGerLAEP+TL
4YmMKvQMoCbW/7G6LWpUiwwmx6qY7nNKV/hxf7Jw+9voAM/xA8m+8j4vLSQWLp91
JdZ5KBNNpNS5BKkpPimEIlXkHSYQkBNJs8L2cR0C2Ljtlz+2mxilosjJJ6F9xR2M
9sQUBIPtPtHTO0XCh1v4AZAu9wbj8+XELkiuZXW661vU/830K/9kER+lWFWHrKdG
mnOzuu5WTIQ0UhbinAScPjLQqbgevbNh2XDM71ot0olf2rgc4OPWy/Wmf5XUKbY/
IWthsxbHmStx/gx0GJKTqflP7CYKuFQDh8ql5IBEcKuzYpbIJDcPzPBW8zmyPl/O
niUf359mbClcvtdE7anMQQhzxMIwYrzLcAyhmDW24g5+6qYXJlcfchx3Li6vqueD
OR2vq4yXGFuzzaIPP4x/unDhLootZ0NKmeqm54Zpr9mpiBnT4bNPgRFyuRLyrEC9
BswEwVrxjCWftImAVcZUtIVP8BKZoNoIH/bICHADm7YTD/G45Uzxz7H0BvIquAhm
9MnkeMEqV+wyGpp/1OtFA91LhlATGvaZYpi1g/B0LR21N38fcaQ1BhAbrm5lhY56
mwP+RaY2j44AcJ9vgWiRyoJvj7olhU//Xp922kSHNsepwBfXbmIwe8DXSRoWC1lo
ydtI/k/MAeSsBE9TvQP7iQ==
`protect END_PROTECTED
