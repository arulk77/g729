`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4jUYkdt5VjR8oFbu7ZiLkkVXiwADe13M1V68Cq6p0utJJGgDKY+Zk/5CbIRQL0pM
lwYAZkhTbgU94ch0vHBcpK7sjUtYg3JtxCmGOQ2tcTQhInFCaJQAEIdJOSS5gtmY
K8CC/eCLnnEcEoTAMRYsW5chYi/4L0qRNfI+1v9MurZolpb9omO9Qcf3Omq2hqze
MFXsiBcfgDGIRFlVwk5hG3NYgwhUDmpQTpdllkHNnIh47G7AgzpVxfc2zmC1vxqG
`protect END_PROTECTED
