`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGdpuzBU5IhgpS6+Kzdn5wzRi4rytvnCWHyGjao5iC+e
5yrWv9Q7iGVIPpFCEBwLQS3GevvxlygfaTBOm0OYBf46BYyWphWdDr32IWRjW/W6
Eze/KTyxmQQ5SB230w1102frPMUcrDBfn+kQswnYA/Y/3RhAupTwiuYgWUWqL1Qd
e1XHZdcLR14IELxNhfLdpdajVQ5FQJ3Y1Zgi31YQSl8NehA1bldnUA6NJgPy1OBj
`protect END_PROTECTED
