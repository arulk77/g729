`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ3jr4MOVD/eDV5hFGHcSt6Vgqt8AO60fPPPbjNapgll
fpJV+gO7xNdrVVoOfkKD5aMZXsTdec3C2uN6xDe3zXSI3DNXlcD2nLeAtI4ySP+G
vUJ3+uAjzgEiVw3tD4XeXgN572cDOfp7Ev/dd8vzdm566q1wmJhwl0sYXlVGSkkt
n797vZ8R9inhX7YFtL67fZ6PP6cSPx50iSatnQoie2s1GRwib+Qjde8Jxnj5SXhF
nV5Fto0TG+upQKIrG/xsG3tTaHX/a8OZF5OYNn15Eq1kGsjS4TDzgfXokySFKzpL
klNkDyvqMAX/FM4ezc61kMAzo34WRcoKoukhJo9OQhzuw1r7LTnk+QEu1RKxdP2W
itqJhsgc/d/wANGycHxkdEOszYtSD5HRTOKZJJTt79By41ybeeUgVE0A9j7esZRM
JXq27MINzwlqckbzDxzC7mAa98MywBKNsVUclqbnogT5bk4aIyqL0SSSY5xQXkAn
YhEG31CUoPh+ORL7Ro+oNji9e1VJWuiLnD/VweNTIcaGLM2dUBJrCKQu6M/N93Qx
ZptkOxBOvvwZw4R2nrrw3DIi14xM0HKd0pe7yoNPGmQrORdSDvxshQwUmLK/NiTQ
7z37wIwj2I49biw09K00yLbGBKSjfvGZ3I7IEIEKYv8CWNbf+bSp3h2/W48nBG3o
`protect END_PROTECTED
