`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SVUMLjqoB0ZsXFHQ/SewEMOzD0pCkiPStCARExcd+/GB
Q8sT4OZtp5Nt3cOGjIYDxn15G/fNBJw42L0hqHnmurOtkgtq+Uof9v0W0Xd5tmwm
r79hzLl2KpwmGB7cLVVYEmqbaBoIZ0V1BaZShWqeaXlzgCgMcDfT4+KijrPN1Zkb
kW1OUyVsuX+8gg9nBtFkor/9NRS10LfODaMSXF7Qza5/gjq7HEMgiw4/pgD6O2rK
9zOnFcu+HTKeGgTefm7QB8rUeCZ1MqGmVezFnsXUth2i5yrf12qV66QUbbgCS/oq
9xk3T5eqBWAZdYpigU3kFsoYFRUe8XOfLLbyUH4VGNoflyKWiVOScmI9UbXhtuTw
0/s+oc8jd1MDA6qGOH9piDqeemDsAcP4SzVcCL0Egs5d83oddelKhTdy78YqGKcA
s0URxy9hC/zWymASEews5PpY2ENMMQVc6ILPtWRvTbCGhQyGNk8MCLIfyRSDKRET
/8F9rEdK5YGn5FCyvGa59b7GI5+F1r7xaz9izdtqIpJ76gXPzikEn5FlwpC8Bq7n
URvUOTCXyfv5KxTD3sC52gbFswM6SF1Kx00K6/MLlKzyDe5hmAFriRlE+cPCjMC0
iVjIWgs+n7oKOMty9T62TbQruDjIVRBYBKVAq8AY+bHhyvtEfj7ysglZNtqf/NMc
8D482+Tc0v+QUKMeiYKGANX91feeytAa2SZHhK1BmZQ59U4X75Zuw3W1B0Hu7M6M
BSS2qh3EzAytOj0h5YKD3Z9u/ctXkTXGrqKz4BA48vgZxZJ0HU+NbOohNrTXZQLj
2YVUGC/YieQeq7LgZRy45YIyy6jpWu+vOXjnU8tZtWCIuH/MMdWFxKPvS5Q/VsTQ
H2WTl9h0XkHa63iyFXxoR5IHWfW1BI0TzWjtDnYV1+nvZKM7Ewue8uIPvJy19Faw
SXLil/VN9qlrHPYCUIiHDxwQ5peRsq/aXLu3TwgXwKzAX1/gRgSmtHtdwStzcA/f
p1oUb9DVQPFvIJjo4PQpqSe+vlINp/L+KJQ4MFXMy2JTBs7sW5upXCKJYWLBH+IE
0hN2grpaQIpgOAkUDaF7x+mmhLjP2xOUFcoZpAOjW0k82CSWeDAus4KK81nNYqJ2
N3cPDu9Wy8fMtcmveH5f9AVfh+vUwdoWTY3NmrDBAbUNvknxRfgMitcHszs+Dk4G
COp4FPLufcB0bxQzBcmMRLMl02f0Ljg7WqdUjnQVHEjt/qC3RTJvqOwTSMBGmVdJ
BiR1oeri3MJrfPWW589dgeypsjcnFRhPQ360vqlknhSJeij2a/HVAVT2MBXMatPK
asDzjuL8bPUEbBRMn9+w44wmBnL/3nE5VB4NM63DeKbR1WWeAxa7qZYRoHSDneyf
PIiTj1otzjvi8g1DxqLq2NyUK6iO0MhACtd9OAEolWcgS5Ey8xOqzC1rxrPbpA/Z
Cm9G3Ii+MHiUduI20kJbOkGTNDoC4+sCWVo8xlpUF+qXzllj0uH2pI3yIA4iJABE
F7VY6WPGaeC2c2wbp2WKaL+8djTAMtd1YivXAu/dVT/x1VtYZ15Fh2oVQCigPcyW
loYaatn7QFAEi8/X/S+DOzgj3rpcVikiQ6HX4h+xxOqRugLnfH+oQ4TvZfrJTNVK
`protect END_PROTECTED
