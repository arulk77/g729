`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
WxVlRxIn5HEWDaN7aiKI0s07/SEhFUURB3JynX/cqB7CekPtaHD8eQuZ9YZH3xof
0XA+C6Zh19ivp3hX70GAkgToxgnp4H2B5TeKLrMhVLNk+V++gy2nE7Y5j54xN4AC
Fqfle+/PRGMJDUSTJDwK59v3F0nreUd13KP1kUzpEVgo7ox2GxUMxkCs4EZI0cut
WTiCrjRvQAye8rZ/l1mqOMRAq7ZGbmJrwhWJFXsgvPm4IkTe7y5RtekYvQgGm311
lGCvgrQ38fl/6q14ELpMYkd7OhuDO7pesONtkjaEq1W2qzdU1YsOjv6vPh2jjTIL
vX6D8v01Rfbe6D+auECVthh1pfqFBPOKsFyiuObvprs=
`protect END_PROTECTED
