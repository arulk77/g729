`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDvGrEtdfldngpNPTmfSHrL7aegrCiNrp6nbnTW512lL
EmGZPj+g3J+hZfHfY9R/ktK4bK53QFeSdNyYhOeqCsSdgiajpxO/+iNiwWCe9whR
DKzjmkVm3Erx3MoZs0zN/AonU8PM0/5OQqw8F40ungUnTZArW1XDtGnDf5AoKlMq
H6cGNJfzoR+NKPVNpzzTWbFzWNRs8OWwv+atYxluFq6m9Qk61P4l/o6G28FkCKi+
Vi+uzPXA4ID/ZUqhdsJwgC+tIdbzfTJpeua+bFPfZjD6i1KVrVm3UIq9CbaRL/vb
33WEdA7tMb3MmKzagaieQS96DcBS0r0xmzYpWl5kBL6loZjyPqx7y+fz57T1O4Zr
R6k4/wAAughfduymBhLkSU2iMetBF+LbfCorlf/DaYGAQ04lhtP5GUbU4rezc3/A
b/yenFrodr/V5meeq6rbv43fcX3AIUKD+kAJY7zn+Pj61tsjvduchtSI8wyDKc6k
0LM+L69xinGpyvBGh6XI8aLwVL7TwFUZOg0K5ykUhzIULHkScxKKYt8gFXZDzFOd
`protect END_PROTECTED
