`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
9hd8pvp5+EK6PDTc8LoqXedkHuzdKVrFJudr5c0oDXn/Dt8hNegnNh+dddNeevCo
XtBoF3Q94eeGOrtC3VLYP0aB9Mil3uz79ykMZsdJrBWYQD59HopTzQz6zyamxzBj
LnZ6NLzz29f+0P6eCBUUUA9I3g+0FjCXzV+vIqWJQ6VY1w7O64kQTarY4xl6Rz6K
B0bCOeRfTCUNR0O7bo6wI3bhNL+Xck5JilqcmtLp6Jiz6fvAr2nDg6bFp3WmppIh
C3HY0sLI34FTnfa6N15otG19+1a80UVd7QZ2xsz06KbxAgPiJ+NdjlWXr5uk7TgH
3Vx6P5ikbtJoOuE+Ghax7d4XFfgoIX94lI16AC2j4ek=
`protect END_PROTECTED
