`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveC3sLmrZ/36VaelVcP1KbM94fjTYpJZUvdpSVk4yc/id
mh9OsYdG8QRLcgTFZt7GpYVRELiPavMpSnBD1boD1P1ifSf5q5e9OISTwDKqVNIA
1E5aJ5nEIl88o6mQjO7mw+r3ERmNTdFMMjwIb8QsNT70ih86JCfiYJvftHeaRnra
JkBxRmPkSdhdyKCx6bPR8w==
`protect END_PROTECTED
