`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKkXE3Sc4gpLyDSV3BXt6F+T03zYeMmdzoDnboRYoTLr
gqp2yhXb2kQyVUSpKWja9ofZhjxuDIbT7Zu4Tmb1X8S9Ndqx6lgvlfz0otpOBVrq
dDiSJt68G4AA9XnKKhR1fc+K7D9c3v2ny0d4bQrs5cx9/FmDM3YCEE4AayFaffqj
p4KuYTofeMMxUcRCTDy5Mhw5hTPTK4tDCi2vz8/LJI/zaoZoHVnjzkOFZ4cP9JTq
YebsPGPHbrD6bNogHFoz8kEsQcL3Xc3LIMADC2LtxJtmf1PN8sP94X5k308b1sY1
WvIPpgID6N6WgFIIpruRRFAAy4nQuR677wuzrF8Vfq+l1gpP6ql0C7exfe1MPOwF
IoFDvwzBkfiBeV5vGOuEr1F/FWR9DAud7YFpvAQI74Bjaq4E5h74kXNVfMAvnzHC
6I9OmWurFZjx5GtnCEwqhZ/37E6tVNp7EQixtS8grRFPlZbxLg6NOeBXtkDTgw1m
+CCZtN4g4hcfk6hwLEHKfRcEVB1QTqlRL5uRzvMgYfFIbN0meFmnnuezPgVQaF4j
`protect END_PROTECTED
