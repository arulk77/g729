`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
iCviQd7gUu8n8SsX/RYoVmst65bJqzFZSEflr0S8PnSqqt6B6RRywCskwpg/c2VW
BgKYsbk1dREg0PVEcE1964thKUV/cGhX/h0npCcn0zSr8wgP2qn6+xEB7QqnWCGE
isHdXD8y7Tun4CnRLDG9rbOLpk1PW/+U1ZLrEiFacVI=
`protect END_PROTECTED
