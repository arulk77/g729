`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDnpt4FU974oobFJPlrCIQ/6D/OTU23k+Z0vY7YtmYkT
vthVolsjbahSmnlB3RFV5y0nubVsKmQpB0LcEuwn5eU94MYx7Fy7zo6XroVRsCih
onKSOLr+1phAjzLqM1uVRvIO6bRHzIQ4gYKZelKz4Jca63aMxPecNpwv2Z0KOr3h
arER0ZyW72NimbFPsOJNx7uBao9Ismjctw0GJCP48DQ=
`protect END_PROTECTED
