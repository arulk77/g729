`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aX299FOIri9nxuWDOaXTsoqKegy4StZbrsmsI5Gfa3wQ
jqfp4v8JPy7kElM8AjwccOk9ZWhOIAEV0MxZAuhb/Z8y8CSMjeuTPRHA1IXk1srO
nsjABnDRYpepcJnD6ESWbh814KmBZaT8I1J465y4Gv6NVEAG/vwg9UCLyqhq0qbv
YvEKh2EjNNk4hhSaDh6bofT/P2c1aAUlJ6hPX1bWRTPNObJ4E581F60EP2JHnxBz
F5V6UpeqxE/HVbBgdcZ4i4NQdNfxwpxdqY97m9/U8uwI9uZncspd5K/OsxDkrpWS
xXjPrK8v/8yZEIKxSX473w==
`protect END_PROTECTED
