`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEXg5nwCQAm+uZ9pbuvaLHF1Ln46isvPEyH5qBNUkN7l
Mvmm3GEV+6avXEjpWdidpEoElL7xOG2EbcAgjLQs6AhVaLaF3+8nkpo94dtVf3zL
Nm/vWRxI7Z6okXhGSTNwyrGDe9Q4zqxK2Fj2qJqhFECbu/wGK+llxan0LacmsKgR
8USXWfIwpWUlzsArqSQAyS4kNodWqaSTWk6pKN12wcuQ6tLe7dLOBXtMqy2y/xei
VQ+pJFFuhWpubgPshGAkD/TmHtN4SHyOp2+2bEWpK/zjpc6NrQwYlQctrlSS0RVK
20BnuXGGCTmFOmotlpiHt8ex9lbLm6EKrDOPWDOqrtqt0XyTPN17/sNq5mg0vkTT
+DtIMvDgYkcves2HHyhZaIDQTEYmPSfnAWrm6SHNgTG5uoUxp/R5ncG5YNknwVTx
BiGdjRQ3T2KV+am/sGNZyjjkpEoswHe2woN4bcRDvqAKZVwdvM/4bf96p4CQkuLV
gnXCvipLpYVEtUlnxsRcuBhnvJNFd6dy1DFOGCpSjm0MQwjL54dAms3oX/7XHpmN
`protect END_PROTECTED
