`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1abz/fvZGMCVXtnHwsChNZ90PLLreTezvtDkI4XHARnk1
ItFu2wSEV7gokZIYXY9i5TsavWy6ak3csqvrDnfI7AOOOxZq1Yo2vd7s3gu4lUz/
Dz8PAYkq1zKX1XH+97t8a0u+eiLOV5su1UDxJhB1sgQvLpzTKHWlciJOQoQ1ovZL
tmk7lBo8qDmIh9GGQVGxo4x46cGUW25Btbjfi+Si3oNPqLUQUCqJauHdUJZ1+i8l
WV9nlAfuALtW1K6Kb8UpbmmlMxA1bbzDDzabFCuTkW4jE9j4zIxfdaSjtBH8zebT
7vEUS3HjDiFpzd3uz1VSSRJNJBfV9NJ6+hx9P5nzgVvt/uSHh3F/QYGLXs8nIATf
7+tPZDBCJtnbY2uYHyXSNp6V+Vw+4C90ssuSWZumQelCqWY8wDSyxw4xZW+40byg
gpHh3WicRERp7XfIvEi/YuotFgK9KC5S31oOW2i8VDXBlNED2PVBGSWz5zwY8ra4
eRJvi862KPdgIXsRJLCB3YxP58E4TaA3C2SNrICPyi5AUxIROm9JfXQpDw2XZJzr
CFLV5UwDOyja+UOAz8ukVa59quBS1PnZBbjqpEHGl2rkPtYJ82x2Au7n2qDhlHgy
WoVZJ9irESHhXJyk7z4CGyBTphix8UrAJA57OIgoD6C2skYVppRMwoM3Yd7BxsGj
tJENjdM+Zg5sniW6zVlWsKEuRPu6ZjZdx79a01jTYJN3M7TIEFxV7FdDYEMCqsF1
CaiawOmoLLvhs9y1lmDGyJmB5lgImYUWkgwsvRXBKwPGJboygos4H1mzQWAAFVYz
OSO9pnYMb2e5x1P7a02jhmK09yXxmer58bb2cDkkl/cMrB8C05L/jzVoQWAWU5vK
SD7DLU5lummPSttmF1YJLZbOqcy9yFHhXrWkjyhXHHQ+hNMHRaQEUubI/rhrpHMX
x7t6kOUUZcYR8HLscbMdz+AWpZCzKQErNOdJSnVkzeDi9htGYw9NSBR1aKkNRxoe
paviDvsCQo1BKmrZnc2q0XFq6w4pC71DiXSzMjCCrqfTJeuOwHZSmSNlFZFGSyRC
kaaLy3+qjLVcIhQGPPf4S1HglORxSdr7jSJ8V8r+CjGC2Xhe11kzBI7gc7IZQuiJ
WtCQJ8WWgMhGS/6FNhwOMaQU9AidsyS+lAVm72nfHtrnsLCsr1HQSLnKilELh9hg
S3GEWjshzbufJXyWfNQms4pR+CiN9EV+VHjrrALdCHlULWHMj7fiwFW9LoHT0CU6
BBiNOKJd2DShwyeBotTkdGQgf0F0+UKRVDW5bP7QrJToEVhdehn3JiIziD0RuuPO
vkdb6PZwUN4Lka46NGl5u6jWfnrdCh690lJHL5/9XsWMlNhj5tbIW3ASfN8+yB6+
aSQ9b8jtxgUY87G9HjYuDCcZtM5VLvGCx+XNiczDL8ENSFOVjObEulcCNVAVgW5q
IXVYuZnZUZnevZHyf1aSXbXPq7rTHNu9ei5skz7XjN2yXkgC3r1HtDcTIOS12lrh
jLqe01vCyKHFPj4kvZDQ+/7aPqCOgMtmyWLlsmBR2DY=
`protect END_PROTECTED
