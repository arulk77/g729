`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBrfR8s+6ywGFgSndfGneMwCnuB6tCcFUPLxC82psU1+
UVdx/7SVHa9naRZhV5xwkijwnw5xZMTJdypVh4d3oAm7BZUegqSTx9ees8nCrHf7
WYwOFaa3lKDXq8yIw5qZgye6Kw5WKenWZv+z5qE22tg0ef8Z4J3FHCvIrvy5nNFu
C2Ckc2w6kXnB0S5up1w8KIPbYjkgWZbfgftqt+IXSx0z1qG8AOVqlSm2De8+aqVU
te9pCi+X3BPYWZsGOkhLJYamP3oln2B+1NVxS2cGVMi4b+jsCXXkf7x24dn4PG/n
bpv79hxvK0kFwbUs4GCYVfMd4LCeQcSgMxZ33ejiwxSq3Eg6lYopB+g7JjNr1kpf
oAsyDL0v7/2dZVEo3jl0lS7DHl0/aQpOCE04oRj+dcZTFnJGQr0fhSzgvTvPspVI
h4FpsmhPfg/SSVauFjCg0pwj5WoBAD9ey2T0pBhofPrhsp/sj3B87PynIWWMpJZE
UQliQEg6ucWhjiw33ypaFgWdm+1/rcp7eB+h/kJ9uYowzb8dXz99bQaGhRM8qP95
kislpM6gJNQRcCMKlpMs24m+Yznfy6nB0rBpATedck8R5V2IUh6EhhpDwb5Lnlgd
iOYKL6l7bA/NP/S486yJ51tuG2uZlyGTBpEmFrRqgPm4isOGoZTQW1DMOA4YSgyq
sXCLo0KKZSnJ3VrTg+lhj+YRy8ez/zJOZ3EAyftZXR1Vu27Q1e1SvAJH9PHDS5ZN
Atsvb5VMKkQDC5Q+gZdTLXyMDDe7UPHOYx+m8HxiQHZVHlTKJFQ67Aoa9EtUshp+
C1mr2eWKfuOEgvMU8HJbr5FHi/H1E2A0lUkKnPRovCMD/6ubruCVWiiWBsUHCzG/
MKBkUmkqcCzKgc3s+82kQjuEsMfQo6luoJ0qCUtvr1oBpIOpZneD7A+uYk74dFWb
bfzDb65x8qwgFaGcy6xbtV468DWLF7n+Z6yRmdDaA8TvnDfhE5VxmZdv8fMvt0Z3
FoFPPMCDf4fj6wzYW2oyzALPiTMdzUfUrAlzpr1QJMU=
`protect END_PROTECTED
