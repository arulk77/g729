`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aQKJvpzfOmi3y1J4cwvvq2sFxfdACM/WFYHvLpotpKrX
fL78eheaa3ewshJgIoXw9bkh2nwjgnXHrh6BC5qYvSTV+Dnruc4CtMHudKa8+0Lm
nhevUcRJo5KdjOIbwN7RNMNktUNdg38YLVWuynwnzwSTPDaw66EVsuDNyv8CJGTP
NbucHeHc9WZD65FHnhjQmRczcCCHs/niBeFCdEDf0pICDGPFm02ElXgZnmpP8MAd
0k1eEIoYn1KLfkeRG+wmaCeeszSaAcnFIfdqCFArcjT2+qqc0dzHa4skStUXleuy
XEMBuWMf8P8jDrQlQqBK4SLhnK92MJQj1iW0pY+lqt1N/fmzleyumMFei7KzLFFt
gtJbT82cKkY/+h6ldhfLb6HQDSb+0kD7KYugbMrdxyfLg5ZKi3vdAYTJ2/BnFSS8
wDPsaDW2LrFqjSG+XRVHjVL6EctSmh9eIUv8+JTC+urFeewVE+7j79G0xaU6Jie7
IZqRNuYh7GXxFMRagwXEnRWmlvQVt4EUa66FZjJZ7407H4k/Fn9vEbPfjGkd4P6I
ChhDdm58vAaJ1FlV9EaTHNgY2MggpRB7APWbzOkp/Kp8OJ39N/Zh8j1Qzp6H3Wq+
3rsJaeFuY2U0TcHPoR2xFbB2FvUeOAYdp92dT/6OWpE=
`protect END_PROTECTED
