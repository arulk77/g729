`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveA/BAUVlBV8p+9BdUl5LDdP7ZBxw82dy+0wGObcthUIh
WS76gmFkMrPbkvYaYhnGElFdfuvkKwRMgBNMf+9cz7uv3IY4WbrMma0NTlvKGzUZ
OK3LoilxFQ0YgnUJhxxNJYMtU5MZurn3yVIaz6Cv/Ck0XAOCrq5Ko4yfcCIDsKyZ
olQXm0hegstGsrNh/+l+SProjoaVxpg5+Z3kVoZrot1/FU/t6WztDYBSyZmJzF5R
PG20anclJB2Wl66rT5qen7iuGocJPcVxN9pkkFfngmPuAL7J5LYGZAKoxjsLqTw9
YC9rEg+U+4hoD2y7jV9AsAQaJlWbflyMA8GqOl3Iuantp8Fba3+0qdC9TV/1GjBc
xi76Uq82JtI3PkrIbizeIFdB1cswa/P3KlCefQ/PgTswhne229brOE1Ku1Xa8d2Y
cTUiFoK9li0q9bGSaI5b7jKV2rfWokzNLS0jvYem8956FIKubFN7WKEQCIynu3YR
NJ3uO6sg/qTvDA13CFK2HE538rGVFjyYz5iNcPlOMiyTu7/+hc3PWCNzUqzXXnDB
`protect END_PROTECTED
