`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43ADXtXh1fdOU1mPKloEYDceiywOEt6YAtbY4PWD2/97
7K9vrGmNNdvE1IHL7dRfDnSC5ehsq8FbBukWD55FJO5K33uRuYhs0bCJvyXHd5ad
Z6nPmBqEu2veMG5AhSFD0D7gyYwWwCdf+envtKFuEIx2Myh2cGQfFyHCepwWVLrs
kJXmFy97D4RZS1PbcZsfSToh6uqZLB2EMQhkVBKc5Nfn81+JMFNZ9OZmRx7zaHW7
URfhaOFTl64pUEKKngZHmrZ4ROKuvGqnAk9M+LKVDczveMxHkG5SdaY2ezHtsAyh
sq4Nu7+9fiaAZhKBD53Zct19YstYSemQpztxdupfocm8Di8MELnqHTsJ6ffjRtGM
9LG3SrIlt8qtRZ0VanjWKg==
`protect END_PROTECTED
