`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
RTf+y3IjC2sf2u0JraWEyMPugJeOHpTUE/kMQ+FVD+p1p+XyFQnCraM+DOnzDq3I
JDzhl55jf39h5gtBlo9gGFbkZdnPkQUsd8e+5GIUFzTQAXg1I8KU424fKK8Egn5S
tiFEBPOj3OC59Z4cJibVafuWVDuIsPA8MLu4PiqhmnH43KKHIzU4YSYDDb87FCeh
EmyYboNF9kBjsC3cyySfSzaYI093zbljMTeddBbJFkY=
`protect END_PROTECTED
