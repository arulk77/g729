`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wcu1nX8tSFH8zPRQlQc4Ysp1eG7ZdpBJmct92arQ5Ap
qI5t3wXdrpNthhSSZ7TK8dV2O70TgiB8hXWmtpK3HtMfLuTuPLRlPmnbqKAcMJjA
N/1hm9/ylP9r9H5mHPSSJB3PG0iXKsjoj8bmyNbgm3OO6lr/1vLBeVMyi8zpb+7j
ywwVSJ/tzCtvvPs2r/IV3fOPvS6EpxxREuM0aVQyS9gzgD8A+nD7GHnpsxmSB/P+
Gf0V4oiTexnaTEWSMCzYmpPFzTkktJvK1Z3+BfgpGe43gIcJ2aIQACYCQfCaCx3K
TBJp2R2CYVmw6o8CeUO+D1heYASbGxAaiJejD5xrpJQ/1OzvUjb+4mHCyHOk32N9
G7ppWRl0a4f+K96jlKHK+tOCOQUOkBCZWlqLZEdCHUWzQml4fCMBhkQC9LjLj9d0
fkuI0o1GuN1qoqNGjpOWNg==
`protect END_PROTECTED
