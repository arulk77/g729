`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFQ0gsufaN20sjw5J94roMoZ78hPy/qWEOs/WdX8JaEn
TgW10bX+g5Nu/E/ZsoMXv+3kVeoS+0bHkTvNYalAJ/zvZP9m3D2IEHsYiG5nqvz5
VqUAE0my6iLnDG7FLpPnn6LdXCOFMuQI5+pF2HhX8IY9MoRrYVDW+VjHvzIY8gNo
VwJkSvGod/wf4cudIVdDwmIrszNdqJkPxv0zSdvCzPxHphqzDWfiFkVhAbM6n8g9
Xy+xdmeENqp2SDts2dzg20rcEnOg5q7XZWQHNStNUlqeVorxp3Jhgw9eBAHJSKeY
X0Q4FRVtxYqEHnlyrQil12Z6VC9O0ul/JJUn1M7SEjBgFAm1JjBQxvlf5Y7pDN1R
oq8SVlHI86mmo2i4Q5bVN27mOVGJ0g5UM+8X1l5B1PnUrpk6O2mK67v5dZgInLH6
646B3vKCLhYE1iFrCMr+WYUcTEiVQREdyEYzkXdkiX4a0ctieVHVWUi1HynpmDld
1Aoa7X9RRnXd+cxRE4+YgxP8z7zos5bRYCjtUJc0zvNNbPjmJR5qgEXUaphBBJnm
eoM0/b+l6JXpvO3FynraSA==
`protect END_PROTECTED
