`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3qhwcJzrKCgmwiTyrHuOiR5lKJO03atql9jbjCVfEpl8j9q4xbcJ8Qha/ogwmBsZ
hx1ox/o5heNg7/xttAFIBA4GoWtwENQvbFlGw+y9KbBLj5ZW4n/qKFixZHl/t6AR
3/H1M5Lhpf0m8Y3Dbu1lrTDNYuFr1bYzF+LuZhTknazEWoM5wgAasNw4+/vWDJg6
u0qupiJyb22yD4BX4B+brr56XaSkxDzWMMgLx0UYo3hUYtR1uw6YuS77yNkisOuE
VoZ89wLW4Ksq+GXI0OQ4JVY6eWkzz1Zz+eM2A10OmYyecTsbMfb1UgpmYHH78peH
L+dppnGwYN01ys6xDmA49uzdQdWc4GwXQiZmZTadEJfEBB3QOShsdbb/KMRbwD+Y
9/v5wPsLjbIPIkqM7B0GFECb/ODK3XJbiZeQq+tnDxn/cI6zjzY9wb21wPYIq+KF
r7GFQE1ibAaxbKYPM52wRERePjIoBzVTMHwjuHkUFCIQYd4yzuBhPJ62Etj8Bpt+
eyaCedRsEfrdtiF1pbbrOdVuSeZBkx50/FcGQrzFurat1k5WgdkpDpIeAf51sA34
yUExVzgCBVPj5rt+KOnm0rLJXqE3knwZAYqNCHJtnZ24cb5VycBinV+wny06M2az
tB29qtConiTkzdn0erOkpFqCeoFYFlpZmMc8H/lQ8p0oht2sC4km3zVX110GzTdG
ZZQg2ZoBiog/OlWc5VVq10qk1ZLvFPyTipH1wdJnOirnpmE9FYcvlHrUUiHBprZK
KWbHSHz6KCQy4SKJmaY8d04XFp96Y5HG3P0Gx6SpXhzWvCvVrJFziXAWkDhNPBoH
P9WaAmWMtaxPTC4vloug6aJqsnIiaNICtAAFXUVVFYiN8xniMYOuOhfV5uu+6ZtE
+2IpUETsATlNzmJ5AF2WcgCJK21Kue54J3/uOV9wwZLnM9nbNYDgIiPH8PHNg0bS
FolE/1vSZnq95M3DoMfq4sXyQiNPIg7TOFF0Kt69DnIUGJgplPp3d3fGdd0Fym5t
7G99shJuEwoLxphjeQIFXjkd9D+5Opoue0GJHSAVJfWvU5q5jYZqumGJjCi0Pkts
JgsPemdwoTw77EGksUcgCydsjiPUnprRp114qtRjaosh+mOifmku9YQgAb5x+p3W
yXgSt7RjQGDcGmsYLKk9xdAXAbUPM7l0dBIMTSMx3fjC7PBaBDnCNMsbL+nkE83i
0pMtDsJm+pNeU6qSnj8A5b81eahohy4OOqzQ6d5Hlm2FXPexnZF1MzToBiQq8+0a
Kllves7tTw1HquZgTPurkpAycvBNtBFVJrmeciO009WoyszfEXE0XYV9QqxVnDbB
Ltav5QyyzZkUdnQ2x0fnYInqNGu0S/nd/yej/U/tGriImJD+V86DcJ5Mqvl7eEya
0fLoh2ZIVLev1LYjck0s5yC2DHMHUS9iB5R63gGDWwlqzoGqLDk5x4c3EqL6ekZH
brAS7HnHTJQF27Qufyw/X18M/7Nsa6HsiZAcM9XL4dngG1XsIuuBGQ+OnxnD2OTK
J4y/jOE72OdtJANlDC1M4rb0FJepkMRUrc9tTgNE5Kx4GBl7agpkFbwBnhxllJTL
yOI+qTt1AqFWROMqcgDuLrK/wlYYto3FrvHrQaJhZ+oTf519blJy5APx+3rL0uL2
`protect END_PROTECTED
