`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Rxmir7i6cRzihxysUdxjJvXQyB+Lrr7Trv3WBSQlcuIMS1a4ftBUZTf+nBAqyVMe
exMhNmNGMHyEZ7NsgBDhKqYJVG6f+xEL0z2tCYMRyp7acwiinBlkciQpcto+9KMD
Z010MkX9nVqXuON4pC6t6yKdDQoUaK1lHWFHtMkGnMgNsHoxuqUXg3Y+/v7BEEOP
utTFXX7vQoNH8U+WsLLm9MhUFSuEskf+1WmyNgdMk9g=
`protect END_PROTECTED
