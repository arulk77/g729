`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
gazXoF+o73F0ED0Ffi7YN7wsK4JoNxhIn1/fOFpgXPgJl+m74IZDuKRA2715Bkpj
dHcEYM8L7cnv4J6VPy6HUukinFNrRlTU1Uv9Wx4RxCcuoPTNcROK+B5cDW82UCtf
FVumTimA0EGNJjCRgekEiGVMTooRytMEyWHL6BcPYBF8fAC4kpVMfSL/d+L+SouI
oPB1M7fnRrP4rhwdI98X1cOO1NzbL8tBElq5L3q16TjBU2wIARs/hLAKWYP/2jPH
7JIFcFo6uL/E8scPOU+sKQ6MCN6hJXARSc8kxZF9qu0DYOMR+kDogjIyPFmnQYrD
ukS0rOmdkOoaDLpdp21vJYKh/QqPeKDHX7Y6nmOUyWgcRl01LXY8+CFFhnImBxbF
YupxLN3Lcaz4rlSqOY6nO0b+Wu3O/lCNz8HBGx6u2ZI=
`protect END_PROTECTED
