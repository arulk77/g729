`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SbY0G5H7s+INoi8hNU2ObbV//3dP9s4yQm7Nztb1aqBP
7CebIG0LvLWgly2C3oFbLPJt2gtCkzrx49muErnszZrJ/LLeOjyePC/TheCGFXgQ
zBDw+ekMzlVBzPY45aJFvD/LSRrvrC+Gz3rLn+TG2N/bC4d12Stp0Ytz7BwFTprU
AcZsqRkeoAL5D5jQ9HI9jDqzzRjCY14gHhzK7C2eQ6G7AMkfPNp6BEgGcIrmlHnz
CidOAwGhNpvDOTEij26o1E66+qsi685/UNTaiIqDsLlxBBlKjVmlpFh3aSYDMb4I
b/5ClhIzjgK5DmNLR7tD+vQkOnlqNXQR+lsjpCLlgTMLAiwAW2/bdVSXJe7BFgsk
FLB+KbNewSWGjVxR7l4F0nZC+NK+0z43/DFWzP0VWeLvxuusnolIxsdmbAmDKnvq
RefeKEy6DGoJum4ObjgcQw2WFADpLWYjTkK9Yx+i/f7iNODoR8qpSp6eMc1EUGyF
kgEwgS7Na0qlH2wXS8qpzQSEGHXc1I+aeLZeh0WHHzYcbASVTtl4MtatH91/+Es+
bMqqfqZYO+ls/HYtkn8ZKaXB7mUQqY6v+lNaCsQ44AROwGbNJ2ACWr69tqIbuzRr
r8P50AzIi8bmmiCxR+VAe8DMlu6x1h8cdkZG1tQFBUuigf2jfp5dznchBlp4hch7
V+09lgxH8A3ymFaDBUjrWdISuBGp7FLUjuTGv1oVP4Arz3Cr1Fd3t9rR2RteBkVE
WEeqRmF1bUkxfazA4qZQRCJFuQ3AVUoejg/SS4kIWTqPcvJNdXvjZa9UMM6XjNRB
1DO+vJfDxmsz+gkHXtTjPm0c3z7lUjZkZTf/ob/8CthWOgrbF4JckCYDvIc6biIl
rDGHcYay5hmd/Kcx1vwPyZYbRuSF1pE24t/dSQMyvus=
`protect END_PROTECTED
