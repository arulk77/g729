`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveH/yQOlDkY/BLUZ1SCsqlyHH81fcjF5/YT2/xcC4QJCn
wzj3rV8z/ov+tDxV5v9U2zhqrB0/AYMf0OEPhxzIytjg1SAx9Q70gJRrXjnhLyC8
WwKkXe7khxfphX3U0colU7FqJ0aHpVumHB6ftJp9QZ2LuWb1GZDiTwZB/qf2bL+l
bKyhYbtqVhFMjVyUOurur26ELbNBJYbYZ+vXf/4yyI0=
`protect END_PROTECTED
