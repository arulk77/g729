`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAS2O2Dl6vBXEJIW6+qkI303h3wkHYixRy5yHclaV03g
JfcsJ/miw9v8laq+scY0gC3NvjpiG56kHQDiLN3KIuchtMLYEC5B7E6BmFCIGb04
fMb7ckVpcfSzj3+ysSCe93VgX7tiGjV1VCgYtJgA3QAJiq/mp0Kn6cQRYEHzsRzm
2u3Mnt5yHxM3m4Ev70L4JSe42ggJK/ieq2+ZFi8TLWhUU84Gu1hwO2dYRv/PsnGo
a1rlci3Vkzk1++rtULFAqQ7VaHXPA1mg72L76LCWlIPEn+U5ut0fObt4VwvGkDtJ
OU5jQHUOl4NRQjU3BycPuMoDTp5RdYPdR8IFdz43F6tPjl1EhOi9/gDdfNpKWt1S
f9D5c0zfq+AEy6CZ7NV+O1xQjUTyzJF28rJ7uOVT2ByhuzNXeCZ+rXGk71WhmYQR
GapARcYZmJCXC9znM5uuX4WQTCzRELzwb7QnvyMnJW9zCmlUtDbuCoXx6xkS41sH
/LNGN5EiS6BxuWrfbvBWXiw8Tfj0QXsK4Jrf3XPL4o/WkLndYOaFDsINH5zfsEMB
`protect END_PROTECTED
