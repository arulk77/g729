`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGvDL5Watn8RMoY1kWf7TvOGYI3f5y87qRfNa3K8RMHI
Xcbk/1ebBRJdncdG9JqECfBdGDViID2eCOsDCOQNqiwHzAzSEgXEt98XVn0+6Ns0
RmIV+vWR6/s8I49xiWshMmeH+0l47YKGxz1rycoW2dPZt1Q0jt+tDYTNXe/Vku3H
sNLEIoFK2/ofAtl8dSIEdQfXN/DF/eXS7vLfnCBJWWaagPN4Oenk33w/0+HFRshh
MiFVKIK5NsBCAs5lDPpYKOMT2quKx4xWhF+AZCqb55C/FAtvKR7d1mjbCFbXllxg
dBDhi8PM2qCUJAS3MHkZjW3xUShsAZ3F2U0LgESZBisyDzYxL3QYCZg1IAko39nA
c2bL9YLDGfytmnRkbZ2U6OpScGYtMBVc1QbPIMgOX3I472++3f0qTcGmfxDhoQ0F
nm5Ud37EU6PfUuAS/GpIgo2hOemB3wp17pc5e8WNCtqcW8am25t2iGtIUNc1qMId
EjlDB1lEhJtiE2DUuxu4qVc6EB41k4NoAkGpK+PX+P2buz9la5CUjfBgZeyujGUA
3gU0Oh9nugv6Rwo5EziKJIeyAgLGjIduZDV27mB+t/ki/feT2/NXGL2aNKynZ2Ie
3Z2w0ktnZNHvTgxi46bj7bmwTzcvCd+38jPQX6Ep5PI6r/BCrIqG0hbqHWNitY6R
`protect END_PROTECTED
