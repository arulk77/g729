`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveE0lgbJeSsXbgcDavJcEqL25taH9y3mnTsiGhrg0p46y
PvYHynXuotuO1e0Sh+x4iiY+SUnuFAMfXXvbmQyNBfiACX64LM5lezUv2bZJEpPG
8a8zBq1GptOu3p2KmxGzMHkrxt8xyI+Dxyn+TuaOh2T+mAkjt8+wooOy2M17kmEc
mL3SBLoXEqjdz4ICdmA0ducpvcBwqqEu9j71ZN6SSFGVPCMuuc/ezPfRKGOreueY
`protect END_PROTECTED
