`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
n8Csh4XCsXs8zwwv4CljhOlEzPQxOKKdc7PUhUv2IcQbbI808Fd8qSCNwC3mutIU
4UPAFfdw9lMhN2HKOLz/hzsen4NgCMDk39uZMwurpayTVNsnCu88sWvrNwMxAT3g
NkWQHcFnKAknRoCGdXPtrnayhc6RRN4N6iLu7ZTGOZcAWMJGizQhvWauEUEUd6h/
kRIO0//JBXvCCtnip/Co4jKDVfggklI7o8j6wW/RiU1alVmdn7hQTL+HiC8hOPi2
cPu+EZjeFhuQq/AzVW85MTxp156g+5KtxOzJ3Tk0ZqQ=
`protect END_PROTECTED
