`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN3rxYNXB6LUQak6q4x7MG3YsZOG4CVdCWc9Qp8jKeKkS
QuEGjxpZyAnL+29GqAYMuI9rC/o36P2LBhWFeNoUqbedSrfWO+5V7hGOTj6ZWosY
87Z9/6I+IUQS1WTKIm3mC5rfHvIBhzkZJGvLOSqdhblBvaDNu+6dtl6CvhW5qVMS
Zcwjvx4gJN3b8G3g1c9bNFb+OMZ9P+R0QzeVSOs/Aw1oTv2UANyV+gPjp5Jm+C+d
IwNMyP+jCnwZ5lWBzLAIi4i/Y3J2F6pQnKkADZf7vi50Uhf1zThnMurzKqAVR3Xt
dLtmjhiHi1cXCodwLDBYDUkT8joiRtq8G4ZBvf7ye2mS+OMMN/A9DmJeCTgv0mR8
tvtlZ6bZZiFBCb3wi2awOtd9oltf4CVsI39djFfmQhgZsCUbnA7Cr6dFIvEM9fy/
VhdjKrCe9stNcqsvmlkaGhI6zALdT/FOtm3zApjmF1oXWqVMrjtZ4r0GQL8J3Kfy
Tkdp5DnZlESGKMQluYE9NnCK16hcgSu1xJhzypZ4Dcwy05cuGIx+bMbIRyEVXODX
+xCCR/4IyK9+sXQsai+2JXoR0Ef+qd5Kv1wSdgbs0Ee5r558CotNQJzZ5RDHBVWu
cSX7BqDnZgdRUKCaWCkn9EhBrrU2kHA9EhDR90VWUngrp9L1Q2krVH7AudD6jEqD
CEOam+Ky2c7sbx//dg/OA/Wm84MCesB2j1slaGcY3QmgE0E0P+JBfEF9MXiBvtma
lks8HmS254dQ4foIz2tKwJ1vTBxs/DyNN/8mybqnS0iME5BKqzaS7rpVlbq5UYLm
YPSgPtpbogzmBsN7SrmOthpozabMP5WSd/NcR62VEpCUh2e4rrgDMoqzP/q6PiFS
R6OXzo5KLm35H/4RbHPhHDvnSXnL8HEcXeJydmMW7DS6U578m7WTtk8SOQqZYp/A
JrKdkXBbehqpKuvi++W5riUZcpk68NkD8f0P6OXSDTE=
`protect END_PROTECTED
