`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCvWl4wBv0K2171HzCmgVzdvMD2MJriVoG2uNEcTAi7/
g7w2SOa1ZeYIo4jg1JXYpkd0aa5xMjM0Ee2xIE4RlFmG3v6MyRi2J9aO5oiaFGuz
PQpQXIdzFTxwPG6PNkbIE8zP0tQz9Jm874g5ZsmxdSxFAcB749l2RBCbvbkWT46C
/2RM8Y7oQcvzGaduaEeJbmF/XdEy6Wao55MBUrGHs6w5AOFPyzTnJj7sTsotKi4P
+ncheYvxwp61z6CAZvFR0qUxmrsOrgKS0ulYyFysLqg21YA5wAUjh8ygA/8ofMmI
WeEgPVjLl78YjrrrAwrGr4fXSKYZSHXZ0KEQAjqKz6HDFYWgSl3fF37gXdHvcV+b
jtiSTIkmK7q/ji2xvjH07aisOr+5AK0Uwt1Qd6Fpj0sKEf1gBo3/b5sQRELcCoy4
PGygCKm2bGTeH37lDrpZ/OZb0KlzrDRe6lx2k1Ctf8uLwfkS83YgwQYR8j44/pJ+
wWvjWhNrXY07xGvtaPHkPhTT1qGfZoe7LlnoI5AchkIxFpvWorKUP0EOK3QHaA0j
4Z9klmdemPFd9rbFiocr9UoVkVYOjs6gY5CgGErAncGFAHP8ud65NCKuMnNzaTLF
pTiodJKx0ZePkQ+utfBVvFHovViJQ4R0FHjPhpAjCMSYnRbVV8ih/ojFDpKYVtqo
9zOVW1OF720fZeQ/oRE6Gs1/x9+sNUUrSCaO1q3uyouauIfvHTkl71/2T/FnRNxf
SeMAKV47deuU55yJDTWKk/RRxStPhlZ4wI/i/HWl4HwtTaNNsor+UcmEeu7M1D4C
jSUlNGQatSzBC0Bpl8IymbzMKOl6npddaPnFflqUmfA=
`protect END_PROTECTED
