`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGTaDpaEf97c8c++dnKfcSGNp0PzvNYFQnw2fpb49iUv
FaAS1vYw4GdynDAjopA2X6imF5uSpGpvhUHSLrcfFq1P1X+2TjSuHK8OVPHBR7p4
WxgODdXaiWjqXmVA9v7rjyS6osre6xmcXLMkVqu/ndQ/+5UG6jWBOrtw6rnRSqho
wMxRumEtWMTWA8ldG6tGnEe4g/+kL86EM1iXdZSO8cbu8f7KizwcsYKHLUrcbmKl
z6j0yx+GtlfANTnTjIhyaXIFM2KW/+w8DgW8B5PQa+wM0LdMUnh6mWAajIsrR7c0
cfF9Ae7Zc2p4QMJqPnjqHDpVAYhWDQ9iOohzQ2yc5AsxqHGjB6tSZHR+iXe+bnGs
ng3U3t7LlCH9eCghViJkwfri4gw2erLcA233vrbcqQiNeoWGEQiznsAEowr1t5XE
fwQVao0UW47qTxZPnqHvl5/JpeF1mTDHyr00dYoZvK0sy1rzdQhV3NpwQFsFo75t
eTqR+qED6VTbWAp9dv46ov0FVjl+27XBoga2cHydTOAGJLz94rqiSdbu4YkD9wZH
g+i6Y4EYtNxIVzxnkCuspYiJmgf5wNdvgSLlpKG58sMbMNgN+zlPkoEMABthMvNH
XDq97vI8Ad2+/Pl09ah0J+IV7qqiB8wVuM1MwW5d+PMHX6SWnbTj/fny1D2MsPrQ
hgCoOTI5Fwgn7FMrlrfm67FboLDTkgZ2nIeSjNvCMuCkzmBLBgBMal6Hifk8FaVn
9UWCKdMyBaGJsFOnFgwR8CjSJqDM4jq+MnLaDxjsdBFk+bIWYtgnGNi0IXZN+L4Y
xDjmJs4UJmoIARs4ZjMgtj8yvUuhZVfGXdAyK1hKqms=
`protect END_PROTECTED
