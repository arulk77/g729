`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLwWxpnovFG2RFhZbppPHkTsVbYE3UazAs8sA6YBOTdp
krav0vzZj9rFqTPujSQDqIKc7LZLvcOTfnYqplf8i6qX1jDp0M/2jdRGapZwbTKi
ZhqyFqj1zEdik03gC6J9BuALZwZ6ZID3sT3TS0qOxXOj8xs4SuTpc7NRVxZ5VBp1
Srde4ARwwgu8w7qPSZ16ZB4oq6/fUErML1psWKzH2oRisO8nw/snFvd+08yquSSs
mRo9cWn5YOXKVfctXXlVLKIA9JGipxoA00UYKZ0vdIKNi+k4xemQ3DJf6+4716IS
iu6DcYtHodPrUG4D5h7IpJea5M1O83qK1DkipAfRlIDEIjEUipQPlqqSY3jw8kF6
bAaz8Rf81CXZ6YrO4OOtibIQStBuH+YK/lK5lkjEFFDJweR7qY8LcrjDWQCJPbqW
VNpYtOmM93ulLEHCj2D5b4VV66uN1sMLl1i3Z9stTFXLB32kdr73CuMXGjA/u99N
Q3pdHfD8sz5y80FvjEaNThsXlmZny3nXyL9ApThq+yKSiW/Gd3mAsebB8d9aNnXr
`protect END_PROTECTED
