`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43xQypioCSdr4A/J1sokHu82qS7irP/erMXn9eDHwMKF
GORHIkEPDn0CjTJ/6pBfab5WLgZAZtKfPN6jbAIr+QnDASX20wNGswGuhU5TnV8r
wFaK+qWtQ7P4M2uNrdieD22uH11Fmgie7921lEd8BEHXPJlhd+vW6wHLJl3dl9vY
uXQzEfiXrDuDr+pLXqpr3JoUHEbXBFWOVo7BZyxfXbdDiuERPl4aWwk5mLaRZE3Q
d7N/a+ZS9dUPRnMY/6XdeTjVb1J2iLDGLMus2vCtECHVkjXs3kRFlw9AFxXFLyEU
P4o/gvCECRyr2VNxvRiadE3iC5KNQN0Jr6P6L4/mnb2RSf54wJ07jPSg9cx7a0p4
y0pC0nqrMaCCv9NnGOTclQ==
`protect END_PROTECTED
