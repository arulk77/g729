`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
fBQfHQyOJdBVJuIA32YoyYFY9fwoKc0DiggCCGhsKGBQL5Uljz/m3m1eVb9gbXrL
Y1x0jKRZKo++Ed9q5SeA2icXHgTGStuTuw31IDRwA/AW40bJNPZoo/4iwE1A0DJw
jS6bNM3yk6d0SomSS3pL7qSpqRVthsgled6H42zpqUpXqyKHtO6+Nd8zNL+tvCSS
Zg45i06Y1jbhJfsDDJgqz5lXCl1bSgKlejni3pZDnnqiP04EguGyzWGIiQCpiRcE
cVXqwfX8agRYwN2pnr6FKax93gDIkR8ZeUhrbJckK5EmkieYFymzT5lZDj/IpFs7
qKrmHBFZnc8q36Kek8JEqpMHNJVOdHvHvf+MxuJ1OlQ+WuJJmt5YVteMlqFMGOIT
DAdHKnyCStsHCd97rodWiQYbx4sx6z56Ao7oFlexiUhotsTNt19om9PJYxLOr0th
qymvyfoWRHIrqpBUjsl6aCpxsNiG+3QOhVDj0k5MDfJdY24G9RRWhufYoGraC7Sp
aw3pnrYxJkFXvPz9+4RvLumZeBzGwsjieeDtZTTKMn8GB6F0xjlpn1ZSiQlyuuep
KjJYTcBGi8vhdG2gbL88Ww6+8EulvzLjdOpw1YoYgu2PQaIBozmg/Kj7I1xhK+FM
mkwlqO8fxDszc8v3UYeGIKrNgwnOo0mAdJnICrbG+zFdNrV6/tKRxbrXWeEdray5
p6c4dD6FLrEJI7KpR0xJhdClnp52Ss3hcM1JcI0D5Id8YAd7vcoHXDwhK2J9H27G
H7HuN2RgwjpQAVJu+WQ964Eh/dCpyJitjvny/QjcXCainLkpQ1lxhWaBqkoKeCa2
OzKuq8ABKHMn4vckORa5DEANRAjZ6zjYyYn8c3Qy7gR/5nxFfYAIJAJgORNO0Q0l
hcuiLm0zcaiPYfHE/pk0iWKYhjqppRhzuBeRgI5J2COTQZ99S/NGGwSJuFXQFCpK
pzlYA9R26mw0qZx9RSiPOEXbU4OPzrkkAaG1/QvCjmP6UJS5A0sCQJUJl2GUhbAR
`protect END_PROTECTED
