`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN6bOPFRF+phQSWSnzxB7A+0rHrAy+d9I+NHcfue7Wvp4
ZdATyE9qrVLIE+mHHNpW8L03sxF3yRJZpiUz4Xlx85fFCHIp2YVsYEWZF9ED8gEQ
1E5QGfQy5ss5rPz5PX+fYeXnMRdO1OZnmqA/31klfmu6f56MKRtnKBAW6V2ywxSH
DdJ2O1a85wp90dX6cBS6MRYuW/b4WBX06P9tRlQUEKZE+4AzznWH8LMxOnfVpIWD
Pna5vt/7hRW3IJQdhu5BdkIksaq1cInejAzXZQh/rv54oKv8yBW2Eb6YX8q8u7m1
9O6D3wzXA+ijtHFsVwar2TJkVKFSiWeaHGOVdgtS06x4vw6fL7bKft0++Q9XLsjw
pz6Lfvvl2Yh71LUEEKnV7XpU6fAuxTNpC7gBOebfSKWQlaik2MbIj6KGrpwuHRNl
wcCN7EKBtYemcIDCvMRrH5dXBzNGA2Dvh6Yt1QqxZ8a+4PYtRF5q0mQ6VjLTfR7+
Ta48W44q91mKMzcadZyEqvkkflVskVwHkLE/KLHqjHqh0DYSJuEF+EzJjbAqpgxO
DTCtUq7m/cTd306JlDZiJyw54xDOwzclZ2hYbNz5uEeAUK9Eahle2WuNKM2fWsan
pYMirx30lwy/GewHzvNJYtvM22bDBzzXFsrgKwUoxLwdG7xGveKjPeU1ThZc2DM4
5E4iZ2P/Dvzhi2k3LNDshetUu0pYszPfU13jVzjPlbMeC3wZrt9IboR4Nrlp7Q/D
+wB/2U+wFh2zuC+Bmtr0tvF08yFHgTM00VOEbe51yFxwlFqpoo3ivUbRGe0ZSoir
Frcv2gDQ52JZ+OaRU63M2iCi9mHz+PcZPQWFxLrOz5PfQ+6KxuzWX+fEplv97K2c
t8gjFGKHz4piNe1g0hbtF2YcGyh3w10OnHUo02Ja/y7CqqY96TaqRIW8h5Jyqehm
sIEvIyl99baDASLRJ/Ncic82ef065bJoIYA5JivV68O+q984EqMSJt+BzO4K3YB7
Dw+G6+ziNBEGgnma88NBpBpV2rr5CN5GpODwu6NmXDo1HaQmPURexMK8a9eEEMTz
bwKJwHIQEw5+Br4JtF9TFXWK86zeyVVLe6zx4t//v0qTFYXKC0Jir/Ny8I9+AuAu
s0J3DxzFFvZkAF+9M3yxFrKyYXecbVs4Pv5hEcptSYZbq6YqMPn0bTGRYb0ohvRv
hFiex/2HPdh6YnwL8p/wpt7XMrGjaQXLCADMURi2qMGqjNr2JFZjj74tWZZH3G1G
+NY9m8j2D2EVhJqBSxMqH7/dXyOZnTnGxn9VrF+Fq06tXihFFb4BW3v59k3ZlNKs
vyuWjp7FOj7kWCRh4lKmP4dAk8zOM2kSFp0/m6VtLfbC/xmEPlXgEXzqkOAcqk9F
XfUW8aNGBvVdy6FArZP7J2YN5DXvvFt6ylKB2PPOeiUySKrcnhyl/WEP51qsyCmb
4PfaFAgJTqMyXEUsK7kSZz48jQoSdXFdNBUylk5dKv0=
`protect END_PROTECTED
