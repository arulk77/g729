`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM7wBIW1gUzfz1UBxABMtZyDlQv3evq3XtCfc+y81cIo
Cgbh1K19tVUqS5CorMWIZUVxR1uKL0vWYT71Fdtifz+qNBYWmS1GOwsB1DJZyuTZ
oG7EQB1pveuOf0h9V3LEGio3WHmpi3jgGQ1yU5HYLns6RbyuI8dWbNNF3tuIeCqq
s3NnxWWmPoXfT++HL5XrqBUcAffqCvGwTIQ2tfH6avqUVAuRMEeVmgSb6GsBYTjr
S9gE0LcZGWJJ4g0hG/8x3NsDM1pV2AN/LX6Zc/952EmGIiW+XI4Epab8r0HYJx8j
VsKpuIwtFvWMfWBDlw2o6Z6b8KjXLugyC3AUaXl9DZ6jQljJaYOzDO8pZuBeh0uH
b8Nhx6HHz3yK+/KeSm0V27G9RWlkaVNoGlIwbqcxVeEmQhSlDmQJ77Gq/w4tVsFG
0g4/3eubUg2Z6G7z90FCztJUYor2VRv+kUlt4iBHURQWTLJlyOJhZEr3O4ETxhLh
wtYbpsJAYcaoIPfyE5bDOYK2x/Q8KQvWYFQ/ds76zA4rM+xby43mVEmuebxM0TKW
`protect END_PROTECTED
