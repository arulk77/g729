`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJbPEubpiXqsEc0IxCmeO3xsFj/KjPebpvJ3XGqE4M//
Uh1JckvfVz5eeRZsfiso4bQBB3rbQc/bCySekFHHlP8dulZW44QAH3dokVLYY4h4
freNLnVetKu5/oEd0t1YfPFj9jQk095+tR4jaWd04609be8GjOk0GjBzjyLgwKS6
Z1GaaVe9G2m1g2OQWn5iZ3rfwrifDuApCXPlViQxjO8uFV7Hqz1GU95K3qlpw3eE
`protect END_PROTECTED
