`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40fDEmPUaAs0o4RlTKvnDAET/QNjyrt6GDEJ/ioZMFx8
TzA+mDY8NoqMh3MYq4h+EofBtIzYe8eN0FZW+WJgfvWgD+TlWe/PGup2iyCzDNgZ
8vy7UHr5nGJKNrNL8fk22aycqu3Um6rY5sr+DW3FIpLweJk6uS/ZMU+tM9wFxi4k
5P6HJ+JbDgVVjTzf4Ltwwr398YwB/AD/c6305e8eYiCYPVauTlvBFZjfivnu8ABV
AUj1RzDbLRiXk/FgwaJB/dkpooXP2KVFTOBjajnPEhQckBMllGLiD0oK5Z902rW0
mDt6B5kPINkqOn0PpvK2DePzVWQPP8yfW3+RVXrADYAztoqsAlV4QZsahc1+YxJi
6OY3o+TGymWeDDYZItSleg==
`protect END_PROTECTED
