`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4z1NvMejhYd10qR4qiU4Cbcp98fqAsfPf5mjtejQfwpD
gBRch90k+JeHS6DMcWdVZZrjTXUp+vyKsjHLM1lr+RFEhcTkQIeum3L8ZY7xDOJJ
BkWPk4Ns01rddCAEyHgqbI7JyUZyscMDdDlj34CiPtWHJz+abLY8NQZqpzV+GmmE
snL/Z1tD45ZhkHfEJanDKLqqzLGklX1SyXP+1XqGaS+5p8YcrbZVQNqSpx9vCxbd
rl8KxkBGceGJeAMEiyWjgiuC0bgCQDedmGIibPfSAqo=
`protect END_PROTECTED
