`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJSxczrNaH7tF3NSjH1nmG6D33bEITC6UYXGmQjdYpeU
x5n348rI0/ge7dD9EuIZiTcEVVguaqNkw/6+HLPc8ZPwAPBW15RCNv4Jf8OX64DM
ccwL08vMgnvNvwqNMJm1r/zrE/e52KuTA3Se3mmxRqeXN8DtILBDDtKYlRZSpT2Z
Ii3AJTxPaqtqj5HSyUDwyREIzpnP8uRSn1epdrLDVyUTk0nMR0XeCRY67pSaMq88
LFwu9PXkC5zhE/C+Li75IFLw+5rg5SBgSfyZoWGoim/yMoW06aapjX0JQneru3tk
aPUFWW0SFR++2bpVSTkTBDiPmlILN0CO63J5uxSNubA0u2U8uwVPnFMOMQVwIgGM
nDFknD9e9mfdr5RenKCNTZdbq2fgfEvUByoWrq47+jpiv4pYrDF7/IdVM6uykzpg
j3wxXn8ukAIb8GYXu3OHmQBVxiRgsgXSlA95P0wqbC9vPy8GX6W1m0vEqlB5kSsr
`protect END_PROTECTED
