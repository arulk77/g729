`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
hBspLIeGxOiWx7k6wRrX0Pz9wMBA6dSsYzFBwqGB/6moubI4zkimkixkfoSYilwK
vqwS6ZXjngZSCvR2ZiHq3Ek3vmphsYSCkpey8M9fg2h9PfEwD7C4G4YyJ1c96usB
FMFqldS+IYvLX+J5twfnj1yhsuRg7vOwvF7t0HHmMBuVoqm9dYHWHV6XyvvwrtuX
pSGaXfwtU8v9SNO2uj9dadxyAS1ClBJpZKty2/6Dh9NCDbJJcMHa7h+db3weCpYv
b9FXP56VRPeL4Oe4oHT+orIdfJqzlYxQjYohcNuyBzZmLnt8OshIAZiQNDXIYwYR
u/pHS9J6/ZW8XZScALBhNHC50Td7SN1/HZT89hvkxuNzZbQmpxv1ZpiFMtCCVa58
b6TymNboTCKfyYVjmmoDcBTC04b/fnrNHTMYm5S1mqvDFLgTRO/SuW7O7dr+Mf4K
QP1XSRc+DstV8n8CItRtLLPbHX/Jr4SgN6lB05c7OBxnr7hAnsOR36ladLaTiqGg
tkuJIawtZFF7Sq6W4Ug8JpzzTDJtmRan3SMKD3EeI9PoVB8frvqMTnw+yogo51Im
SqrqyhF4hGZwI2uUXmefEtj/lgZgKYERDMtQ4q/hML4pjtfBN3N8m29vJ9BsuLWS
fm2jmEZreeHn4grX8LiYlNRX+cgqDRGyvDmn7Tn1OZgOcJ9nxP0KBhio1J/Kki+m
EkswVF6wUzUgSDCe/OSRRDrSfXE0MuU+BfI2awb4xoP7NqP4J0aPwVyi39Zmxqq+
HQmYIte+LAvCDa1MqAGN/kRpbNDG+G1WACIwrVJetDaC5vqf3VMyLbEeusXRFoSg
N8pWhul+05131BDJKeO9oJI9PWIGVm8GiQl2YS157qYrVs4NlxGLoAQuHtTS7a6a
0gpT6w92LeLzPaU6A7VOqycDev81Wa7AT1DrQ6yjmnmzw5LlO9v2MymcAEZHPYuN
ypEW9beaIA3Q/LKsl+cCGbi6JoDiu+WR1IeLxQat5QvRkZHAJp3LLYOntxR8VWCL
EMQjAiKaNA/ZBHTHpiC8H2ZZo5e1M9PZO3p4ZF+scLK+L5Pop+ajFy3NWbF8Ok8M
AH8JCQT4KBXM4b5a82qxDy7SGW2D5OOTg0vpXkqhRbT41iqsZPSEF57fTlALhSZJ
uZI1ByWW0n7cZkLwfdEAe8yIuNKan+zy3xYAKhNCj/gLgdEUklElbFXM0UVLk6mA
vpuq7KIG4EtsEOGFmjMv5sqmdl28oYvU9PQiIHPyX1PXwsOSAgU9oo+RzTUPcMS8
W9QyWkVCHIneUqR5X3v4XtLpr7dvcO+/SUOJJKH2gYk0Fin5HHxFVm0sV0ZYVD6a
jCLNKR9R76avGQKlYarcUg==
`protect END_PROTECTED
