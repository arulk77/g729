`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45lhNsJoBVq1tUh2iEl72+igCEKQJ8NfVtQsXHOg67hE
f0ufteZDPmGuaPSSx64M9hEgalr16gTXZIU+5l9bNi/y/3CTAHRjL1/RWOhC04wk
uFo8lVopzc69s4NMajWxB4+z2ibKc4MpFj7KvP4TREByhwznwmigQ3PFAs5BdhMV
uFI0V6BiKoZ9Ppu0KEwYFRSpQi3tTlba9ny4/JlLVF8=
`protect END_PROTECTED
