`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aWe6DUFa/9+RiSsoA7/StgtNsw30zhcRKmuU93OCStxz
YZ2iLAF1Bi9ZjSfo0SU6FgEjukcyYfGmHyDshnBg3MbQtoyKIG3bhUTAwLOG4tJu
P2egT9mUmHZOEc+svLX74qZnrXv37LLRFR8IMBLeCNsWZvXWP3fZk8iaSEHlTmL2
lalQYYQS8O+82853n5txA1XhldN7OSGu3/bHMRb6fvOaqgfZlBoJCIPSEIlQlxko
7P2/Hqnf6E5zOqadRCRURCIB9DPfSYpolC1ix0WdXYC6m82D8pwf1BLFaTItaSX2
9OwcT3XKViQcfoeAaHAoOYrsaHYSiKuHIJNQCsdJJoEBnhYF78xLHHoBvx/UX1IN
IjTDOd1f2rfUpnvVzRsTZh5mxLZs6+Z7KUxGbh6o4Ph2lNANElIxI/oLPEFvWTYy
pHwMW3W6KT0cJOvzcjUGyX6VHDYhn8+FDKS4Gtp2xbQgDa1m6ByPafEEzsLs+7bn
tX5PtxYj2OVwSvNOYh7ds2D9xDFXr6BxL4P4vb9fBT5QtakoQxebS2SzVcU8PcCO
XWz8poLn9LbftRwRnlvqsxqSP9+5Oh3qX/TanG5gLZ5rWqLdPMVLQyY59L9n6Yw7
7HjQyB8YrIIWIs6LwHMSVtWRSq/DNz68MVpru3cxbQCqYxvKN4aE+sWQD8xONk8c
N0ez6yzOfu9N5hu48OqqhZrob3pwnIczlLGlo9f4y+uCOou5Kv1xL/iMGcUikT3c
xExZYSAI1Qgqx/GyrqCPgB+FoFLxUbDKKUao7QyDas5ttkg5jo2I2ypDHpuJJrZD
Orht5kAAwm3Y7Ffmf+nBJXz5gkKMNcanE9Bqm762gGZtmZc3rLyO40cdu18Xow3e
`protect END_PROTECTED
