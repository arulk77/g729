`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ReIsWZsgy++ZoKe2Uj8E9EcN4I17R4I6ezrwxIPJuLSOv/7P/ziIgFTgxSkKiyeX
hQ3wuDDsA/rHT29tMQKlF85+kp8T6EvHfA4okpYBZ9+NL8CrMVMWUKzk+l6K8woc
tU/WFgzG6aHbIcHmMJY8YJACv5WCfL3XeLl4SytETizIGowIfzG5uQiPtFZde6Tv
DkKHCsMaeM4NvoiKDnYnnAJYTsMdVTeqnOShA7vkf/cnfGnmvoqvkld6Pcr/5pSW
JqN+Oh5nX/5onKnzK8IIgJ5g3okfB0yRqIwPy0+TXJi4CRrWoO2cRTz4eVQQkmWC
WriKO9oRsEcI536RrxU9daq3at+lZlZ0g4P94humOVs=
`protect END_PROTECTED
