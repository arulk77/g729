`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42GBXEF9Y5K5eN1x6qoC3su6z3XFp7aTAHxpw42+K6tr
yWYI2VdZfoQlulA6Ec/WNsrMFtTKTpMvTcPSKhdB83HS1lwF5SofY+SM4KKtjxgI
ENpWrKw+/p7ZCkQLk8ECUHfCcuH0KZRi6rdRn35++70WHz3dwXIpABhqAcpMZEZC
Eur78XU5rXylhXYKuat7qcX1w/qakBfCh+QULgMxBfqBi5akUWx4DBqRd1TSxqeI
w8Vwvz3dPNwy6nopTXeUf+XjR3IZFhyXZIFcm+SaB6Bgbfw7IgCLdRlqLWNogtVJ
A6Xp1TJ6iFj0mS1XvhU7NmZRgkJIGHaqWDCk641deJaIUNMLjc0ZdiX3TgGOmL8A
vsnw2QPlyQWPwbnKHVsD/Q==
`protect END_PROTECTED
