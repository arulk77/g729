`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40oJPmPxbMRWLKuz4wXGGi5sxGICuCo2UraQMwJVw1lI
ghSOi+eZW/S03xnQb/zFPa+B0RYaGYya7q4ZOfizodvQN6XxOhET/BWYewDsJFsV
QTxeE4yj0OPxag8CJxMDFSw78v7SY+OhpaHe9yBawYlds/S5G8hXL9O33IkVR/ZH
i+IYzLmqyaB373naHgWH60qXs+pKrQSzQQAyQjsdMPl4mOxc1ggeKZ6b6zehlSlO
xhe7AXoJqduVbYGm+7T/EQf3A1vHGYveOeMGGhw5fMYFNbVyA+q+FnWVt4ygag2M
OVMBkbE8uLNojsryV4zZ8A==
`protect END_PROTECTED
