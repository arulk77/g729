`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAbiBsKXHrIDcoWR7dqiZzStBlYrx+qsuwFtgVaAgRXIU
c4t8jRCVvEvjVg+foRP7qtzbg2hX4IkMWn8bpgqVljSgUppMjLYRfE6/tw5th36i
MqLmVtZFaKI60nZiQED/2c3vB2N9YGVCkSGXU1Sw6si/Ykk2PXNf0fGbbZXV1OMw
+ahZWKJYQj3Z03HHTm2jGJLihEJKRJgC8vOdo6gzAPiBLBv6TjS+i11sRwTn+CjO
tD+cjlciPrRZGRAjRguyWIqzt6az+hE37yb/KWCvt0A04xGOGxaOR2b0JJ3KOkpJ
AnFkD9yT1XNaxH2gzi7s7Lie5gdkkJPTPK1+OFhpCqJLn0PzDAyJwZCYOmcI/993
4Tk+Svut2u/u4A07gLJELNpO9wRzwISPv36ugwLUDahqCRxk7yhZqGbj86Lxl9gj
HVrYApJ7kbnexy+Aqj5rhjJPuRn0RQZ0x1/P7xmth21N0Dixqkdqnyikg8n3E7hy
3M8xCGlwVy5CPyasEaD8/+rdttguXEgefcDUqBgpjEQzMPHJOVMi6CNOa/6VrCIi
YTucgR5rfRo7L3zdGXoSWoQJw8pVRBuDk56rc7cmkYtpQESBxnNZmuWWUCXNL4nb
maD0/+1lYYc52T2akqXHllDRB6HrhHPRxmK1c1AI1PbxrQhgH/gBjUa1GbQorCIE
d7E08C0OQTLCGCdCU2HCM4E+6+62f2lVR6DHmUp/FhHcpyMNlPYq0fbTX+eLm52C
dm0hnH9sjJzxT1/KrZWTG71X4xMOsmAqrvi5CHMXh/8CXbeE05xGKQYhgJjswUfG
`protect END_PROTECTED
