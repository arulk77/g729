`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Nxn56uRcy9MaFJBTmUlYGePZi4Mt+YTiNr0ckcGITh9PEaM+j2gdk7ZIIQ9cH77p
FkvibH+Wa+DZQDyBj/YFl1bLMpdWIFL3bjVdFN4J/lixH3Tax8Wtnz/qIbWEzl/+
AYt25D8kDd8bxWMm3dsSgWDcIQuzJzSSAA0HwZgk6MPBPakno+hqycL6zsq03GXV
JmWYSjjU68HrZGDkVCrou2tTsSb+9l1ZBwAHeMKjlWXkF7hZ83cRv0cOvw6jFNr2
P4K3Wk8hNA36fzsEVEjZ0p5MEpg6mcPGzcrX+oPJuypkZzSCRRQUlQBRfywU1IHt
pDIsTYpoMhIY5OlxjPGjdgljYNY9UkJ6Dsh4OYVrrYqjNIToRY7xXvjavmsBlRgL
T9Y9R9SAHCVZTMxCzYEdLxeHfLILXQydFEHwVpHQeQSDYy0l9zQwwVhQ3jQ9yNdH
dvD/S6Y4oVvZM8kwyEDWxOg0k7Jqd6kAZzlL7wm3pnJsYgLGx9GvZ98rjnY490we
CQ25sQajOg02LCYOhGuAjn6K+8MHImRYpY/p1bObzf2f+wOzE/Y0jzwWMrAWuL58
CLb2gM3G8gKfj/Z8KD1EmWQ5ADePMVg7WoEjdrh/5BHy8AjdTswkgKzqhUt//aqo
P4wVZw1WgCalWyuX7fKJRaL2t5qwLvV19wds6wIRv3jwI1NbG+8mltcV1vqLXhlA
laLa7XoEsJHMpmV4Ob+k9EyW7F1XkRHOSUUGCvD1DcSM6oO4yJ6fqehvl1/Vnzya
oIMxtuG7ILUjUa7JxJ74qzbRPQp5q0C6Zwf7rcOiBSwUs79AINziItI6/rdr73zD
wtUkt7l6IBy+zHhdZ/2MuFvqy5LFbDFGH/+A2MuPx3dH1YA8dmxE9acPw1w8dWLB
Oe12ES442MLOkqkQnBjGcrxik0ltU9X9YDvspUOHUUbjgBj6qeTOanvKXkej7Nod
gpyq/i15q4elBnsxNhSSqe1NdZbs9+0lHGPk55DCwbMxNKR3wmthH4EssZOKz/PI
h0k8/tPHRLLev8YuVduL8Rjy68XEQtmjthB3s7wC+aOAQGWKc/wn4GgyL94NVb43
TTtufUxQeVAj/P2WGKQraUypeRj7ah+jotjCbfcdLWqyC0r4QeGiFI80icMkKli2
Tw6Abr9KJvpbP3De+gWoqkJfg8RBQ5VUI/XszVzMl4xJIWsrd/wr9tv/E6GDEjfX
76f4ykR4LJw5W/DqxncDUR+bIMsyUcKdENc65VKYcA2zbZdZngoUtJtUE+CE0O7k
/uTBQAmKAFPp2fsxcQAXzoR9YqclswrdiIgGQWNW/qlNTSgRlpqcYaGkPOsvce3j
HaEIIX7pw5wdd2yiu5CGJw==
`protect END_PROTECTED
