`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveA4pPybcNu6rEqbJhfAeDELbJPoEqKEaIhCioQi7KKJI
48Dt4JFuv0uuWbJsw+G22ed21SfJgKcC3Gno/lygBlKuL27ET3ceFOhJjdYEsny3
Zig7FgtPEtLkmbopx9JlqXNLitnGXFfrTXZ/oevtJG/Y9M7hxB4CEvjRc6hlNdio
kw9wQnaFHDCpQ6p+hHW2QA==
`protect END_PROTECTED
