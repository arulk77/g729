`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLKxXponacUx2EUaoKVNHvg73pEstCMY6d6gzVbd48nM
9IOBQUJE45qkiH/l6tiJpdL4QpPIjzn5i/zRpHvh5W0yTdS0Dzrw6LS4yt6dIhEv
2zRZgyDBJHVukBZsFXVydCZvXvwfCR2/jGGbQGHWmbtRWrgWcArxub1RcfpfCjCS
dOJmvintihZ4eEe3Ywps4xW575zQq9TCiKPhYnbkWSRxBhMZ+kAndkMbigiQnQNU
pHA9Oi15NPxbVQnnd1G2Ucqr1LnD3k09KcE1YR+C5CnLWYAUobdUAXBAX1lCpjGe
3LXpZjJDlkxoX2XDHAaExA==
`protect END_PROTECTED
