`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN7vOQiXqTFPyJ0wys5mpWQ/mmw6b1bQIo7WPBMXzjQDT
EGfYI0r4np1obsK8JbJG1c1z8QoQlL+lhwA+2nLG16ATP202i1h/IfAGQjrHqEMa
cdKjm+8ZKfwqRWbFkI/a9KoxQAa3zgod9Y/jOI841le61h3+qHozZDv4Jd06DzNz
3aUJ68oe8bUBoOWIfKLplWTiwWDlCIkQvd8hpmEHOs9UNhs7yx4anjge+H5nDwb7
aJSKzPHo2uM+h7r/F8sy97jQzRJuJP7DG4sHUHw6ylGtV/Sfft5UvGLjwJMF40De
Iogo0eqcqEDOSiyvbS8dMs+oQGkXn0kzmugzEcWIPI1wy9qht9fPCZyvC4RsdsU8
AqSrDWmsFwlvldGYAL0qrHNjBeQZej1SwZy+19H8nxIE3dK/9+AfO1dRHckPgcU8
sPIeeEtIyfgE1hofmk+J4gmOV7/R8ZgTW7uLgW87M4Y4r/aeFrEyUB1JqJbV9CxQ
Hd0pTQbkGLorYBj9v43K9HIKuRAEBp32dRXOQr+G2dZCU6V8T+cR/iVwjD9SEQYR
lcjLanHicW0xQF5e2F+NBip6LWKQlZBzYhHCY5sKldChUSqszo2xjblSoH4VxCg3
K+Xw5p/6DmePiUbFvavCZ0ZwBq0rPLE7z1DAWb9t8YZAr3SdR4YzXQpAU37vtfND
lDlPGJEsO4FGUwqRxP6DU/+Gl/FZdcStKFXVBAmDlxH0TXNj+B6l9uydl3N4m20N
OPANv34BcYAJrN9hvgKAup2we4Gxvfy+MciMRclNxKY/h+VGWbxujJ+8f+oapUU9
CSU3zg3esdGtwfswPdjJfKUgF8cr2ys26tnll0orxGEBdfjD6mYbmJ12xV+Ek7Ef
ESh3k80LXuNmwI7W6O7a5DvGYNmkhjxKALlyBhBRSdQemkN7WYd3khIRHU+hOi0q
/vr7WKuGWTYeqIH/Gkxs96aaGQHtbcHYPBt9gv/wBQmHwQeJrg5rHDP8A7pgBAcy
grJtC1zBY17hOOq37/tQimjVu69v80FUwTyVvT+kG9RArm03nTW9TZRLYzhlrTfQ
V1IcxD1yHq85AJmGdHkfASs4z3NUUYGgU+yap+kRuX1llMWCneYBxfM5fgDdAld0
Bxq/V/N+V9hqZPAebGA7Ys0GU0sPYLUybjyuu3O3AndPesFBCjeffvvSbsjNx9X8
rHUXEVjwi+p/r27x348roxgLHXTaP4bOoMIl8DhJ4WpyttKDEcAnG/Fy/+tx91+O
qU1QJciflElAUrcg8u5AMOBk8PL2YyObw2A6rzIk4kDH5HZmzv6atDXhU7Yvk9pX
Tdn7Ry3p4/IIBexcbQCcfKJrtZ5V61WbKlPr40vDBKNo2IuIlvPI+WMFoxwVvss2
4potc+QJS6ouGv+jwxR5pIsQlU1QhI9wYdC4ZOf9pgyWe0aA0mIO6609w9zuEsnz
8muflUWJWsW25MgS1eH5fhBR/lq2p+uysZluxXJB19EqY8M8tQJdGGxdrYk4UsnO
fthfhiQ86S/SY447MsZF1HQ3XLs830WTyvwEgQ5QTU9kcFlGm9vf5D9/v4AEvnqu
a45UHj8w02EpnPNNVTN5TGcn78yqPfwLugFZ+StZaw4Tms3W6EOfguWTSQMV7Hrz
6tVObwMCEKmNyA+MhYQRJIXLXIkVq9MAox1RaAHw3lTbdNTSL1Lah8aYiSYB23/1
Fng3SZz78u5ohLonzsEVv3IwNa+b1UkGc7g3Ruf/8m0JATTRN6aNfNz2e7tYreZZ
P7qXNWJ6dVF1MlTfM+E9pvtbswWJXcTzqxmyr5MNgfRzIAMI5PJ+H1Otoeq3qEBT
`protect END_PROTECTED
