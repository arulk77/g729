`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBSJUQp+wkN0ZKR6wmE7VvSgOx4DUeHpBeDybKScMNIT
c55jcCASJRnYsQbg4+AwUFgygX5CHKChJhe/ThbN1JiRcYvztwedna2UzJrL098F
MZloJi8FWUQh3WTqEqJZ+jn98yERprR4gkWWIKwggv65/7AWsKNY+MnEWaYBMwYD
gQV+zwVJWBn70v/yrN7FefYJDe3a4awPYUfj3KKubrldO5AmOnFkIH1MQwUWQ0Bp
0EJwMJtZ6DLXmnVD+vmiSQgymgFlflG9x9YA0ALddkwgPuzX+Cn8iXDce1naMqII
hYwSs6WGB54JqDJNwPi9OeeLUIyD8XR2g+wnWUX9zldwIJd9R23cYAN4SEDvzjSi
WGM26FJAaX3SOGcqJUhVe9XRh7ktp3Kdya6+0vKuSblADuynQGKbUc/rfxq5FKDK
qr27kPPK5M8Z96GCYXN+smh23UwZsXcwZMQIXiWw05LfEbj0wJichKnqVVF5yxC9
`protect END_PROTECTED
