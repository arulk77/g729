`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHtN4y0TEFcwt0JewAae64QJvqJAOIoqsD1lf+7Zimho
DgGQZuKK5wDu6TvdMWySP8OUpGua0l4I+0DKJgFdQF+vs6NbCAf8Oh1yT9c1bbeg
A+48fAXlP4HcZjhsaWhkoNtCN9ydCEXWB7eEyLxDO83QpGUIG4e0SIosh9MPPnCI
srV32tm+1oAxkRM/83qipUb0m0HzkXREz4HQCSGg+wOYkDnYflkOdoY6rt1Z2P8w
W3vYbtM9Aciodxe/eLenyGENi1DKR6ECD4fSAzaaNYrAfbFKSWdqppoTIMZ69sV8
Ple6EiD7qf5y8XlQrDLNQkhdcE2tiVjPip4abS3Xx1obEQA4gkOTOJzaMtAlMkq9
Uu++MIYm/0/WN/tv6fxDhQR0ciDhm8N2Uu8Eh1jSK03KnONMztSn7kVS5JiBJCTy
LzHViQYQzAjTpREl2d4fFA==
`protect END_PROTECTED
