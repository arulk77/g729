`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
PnmGCgnHOiYlw3h4TaZd6E3v50zce6GTLZjYr3063qe7eJ1B6JGuSGMdDKNExXk1
vIy4vkIGwMttkEFPFE7CxvCcDkUCHHQohZtZFpDFCXKOCxjrIWIoof8iPfidEqIo
4UFd+C82QZ1blrASMcJC87Y2nOuz//bGAz79Fe6I5VuSccOOoTkfxfvi/7/F6vOc
uafILNjX0RWk60YafrC4R/5MUc8/JuKuKhGC5oOmkhNPPUCcvLpLHKj35/bqU7gv
EVPm8JA5jVVMspuWxgjBeil3DSp8EyuiqXnmaOosegwMCRPWkQ2GqGdH6d8Ex76D
TEgekbXGuwbx2GJIPnVt13VqfJJ+n/+Kd4VNphAQLz/5TtQXxR8NlgF8+wYgzPHO
z8xNVnZLQJNxBaYLUtnLvSAt4nZEdFIJGZ5dPDZ95As8X9xiqS+2/W6QbRCMqTdN
tZTpxbbpMHp8trs3ubqq3iWQyRTr3nkhm8OdsakVzh8zLH3/7nm9QttqeWqllQV5
/E0n1RMBhi/rP76qXjocXhlOK9WocJ53Bi2STfBltD9JvN85UY1DwZhYs0CfHcuw
ZjjpmjL33fHM1MmQ9PWOcbMo4kaCdpqOxWrHthxScFCDMdJhImmqcgrhdjGgBLE6
bbJPY6Iy/Fe8mDuY9y5d0oR7fi3EPRi6kioPUQ8SO0FKHfbD3fONuj0MWPO5Em7M
hQ73u1SW1MsSswOg3m2KiUtTyCh1FmDJOxmhi7McI4dTSh+TvdS0aaGoxEjqBoKC
mj7KZ/Lr0BlWOhr8cgH9pRjKBr1rT8o4u8nJRnFG8IhB06OEFURRwWzhX8Mut1FR
qHnzCLIqCVbraZm6xgG7JUOEDaeuIkhxBXmcyIy1oTlUjW7JfmKg6AFuuF+fxxhD
dvzkoh3QyJAtTkEasTZGiUPZxnuN2oYdzByUYhD+ncv/ND48jHUIUVe+MGD1ngDy
TaSPJxA2v4S3grGLySRz6bSuarYv1Di0O7u5EvsJcij+N3+BzoJIDmSyHX74oDNp
9FR97rfHMjtxd4DzmlobRcJUR5/jh9jYjBJFE00BUKOasKmYM6E4dcKp7uO5z8hi
EElRsOhtghHMyflzR2pIZxQFo3y2oGEhOVX/kLHPFlA5BdBoVharIELjW72x5gsp
KHImpsLIZk9p3P7DHrN6qBEBsSQY5OohjwjUWwmTZznjnII5x9zBcySTN/MSYg2/
/P6W145NFGCccecklrUCyqKk44aGfKojnvv4v4DHlZvsHVcXuS6nG6az0WRsYYZi
YOY7bPObWIF5XAwMHJ6bfYaD9XnOlGAdegRQKt6p3cmzybOr4bqvdC/WqW5PBt1Q
OfbHLrqgfPbzNE2LQYDKxHXS/WoBAgPl1tL0zV7FZa1rS/CxYRKr+oCNc2jiPUtW
hjE+clgmu+H8Ws2dRhu2NSWx367eYFH8sznXB9U9Ub+5E66O1SuUqxG9LYorhHbi
e3fbvGrZfHjqMgsJz+l5AyBcQ6aprlFh31tQKdfuo/JhqzE+2bdX3TyTfuWR5B7R
NM7qFYxOnTB4gc6fEQO1qYGg/9pes+pf6Q67enOzRGhDQEOqJaU5IDmiHFpkUP1S
rSBly7WvQ5MEamU6ibnJE62/zup1PQ5LA5y+RI1j4H+zm/5YwCJa/RSFPTERmBnk
nGKt5EEPMUaLaXpzFWrXZlECo8BGy0ijnypgvYfHPVIJY/7UQ35EEBGEGk7Y7NL1
26z9bf4VNOPaayxBGIuLhTYeIyxogrZhYL7MusKitwT9wpoYz4hPSSblCBCD75ZL
b1HrpMi9Fer7zX+7uW9TsL85KvwFlq3lysliGQ5h2VvkeVPmzNi96GwIH9VSNpta
SSfEer2jiMTBhorYyRMSRJpriMzO3kQotxHa4OY5OqIai4naJWLpvIcPhIj1PVGr
h2nrgQboHJGNkM7dkzflp9uLoJsIfjVeGzSy3IwZR+ow3vs/dP0wC6qpZNvPR1wn
Kteyslyt9eolDa/SCyImCs2Bbupr1DW6WyDZYyIY0B9gzOJpwOPhdGU4TOTLmwQ+
tDeCvrcDHsXqu6xpG0uaz9ZGEF8o97KoeWOGjxZ4GV7V+VCOV1/ckM2j/La5xOx5
ovBHQbsgLCJso7rI5Wfz7ztxZ5U9A9cC0UEnsKJvPWPRZ3m7ksTlbSuUIGsl4sA7
+LdRt0FhK2rGtZvUs0BKLFnXPY91a9nw+4gU/eEryzvSnjrM/ADQRFZ5i8VLEE0m
2uvRvWqQiiVkQCV0bdkjLfOevNNy586sZOLgZSLTZgyhvL5CcCjHI95ubsrbOCL+
Sv5xnRxuOh7YZhuul4HSfogC3HwVBcF2YTADJ7IYybu8wSST7XkqjrMopQYLvM98
2yNs1zIF6Tvd0So+V71NFQIESUZkBKkyw+J1lotwuVDkKZXzeIMDBZ4UM/G/Ei0F
jIMu1T3Ja8mdezKrkl1QmXS7yx0wcKnGL2JGzx6+MTtLUDbFeo3LHGU+LPjNvKxq
6RyXmyrG+6X+DTidB5Y3J39Mzyk2YAfEpuA9R9pbskw111ZQ/kmGe/D0ABHiit9l
pnrwgD/TrZuQvFm7xgr7TIz67tM46uu2KZhsWv+NeR1FydA6yrY0RixQmpIF5JQT
q1NvxIGnAy0M6vW+riKKsCOGnBeO75/qTeskwORqH2H8CrHcfS4gcNH+gipdOcRA
O0CFvTs/SwMQBG72BwuRX+JtGVjJkcpUEVoz6DNLcKAlXFe0rokmSaKEsUX2vtcK
5ftLR61LqajITVgFyaoDptIW93+KktDDlBIe6nOR7HrC5SNLa/W++SIpFR4ERl0Q
RuLOH6padDMqASuI8c4Iav+NVltZfOD9jJ/25/ff4uYak9x0kaMIldwWUVSHeUp0
EUSifdW7d990A0psta7SzYn3S0LHxEAq7x5Dn0evDJF9+hxjrqiC8tS125Ikgm/k
Tzws3Wxe/0teYCTtoDxFG0mP8IOv38HLBAM3qDE0q7ED26pnIlM10TxOhr7N9FsE
Jf7raIXJiSq7v8rrHpvHLMsSh4cbHG72SGqeXv9VWIUFdFtOagr1vVgISx32E9PV
1FZWZlr0Ys4YdSCl41aJfLz6DFcr05CKi5/YlFrWrZoRp/ZrDYUOnPVGAtwo2NNd
Uc49jZo2HahA1iHTRvFbT1JMQQ7thF6WWpbQ94/UoXZnl5ZSSioVGZP62BFQRR8i
LjiG9U1Zef3b11fZ9Rs2YtnogpnvXw6xSp8hEZCdqZtHCa8CHNvgfPDdlQ+nH981
kAgbkXfPlVzltuYPSDKJFZ/JfCp+M8zsfr+QWiEZ2ALpm5haXg63uRFEDNW6p6Ep
U9+AKXdfAQcd6JnVS/yQWlKn9ySmxMQtoVavftP+0hr40jVukp7z5Km8b00qUSea
IP2PIaAb+0+oIhKMLfzYWy1pSPPSWjf4+zogg3A1ZpCxHAYTfMSuLnfcsNOLXm84
yxZU4mQDftDep29oDCe/rCho4D+/SFkQWZiEViipRldgVWvMENWP2rMVYpJ4v3Nq
tNfb/KYClwjag6zeOm3/ifgSTFaX0kjoBFhezaxdb05/ZFAUaBJsDqQ8RvtxcuA3
pKo2EEBUe/v1qx19Ixyv++IlreR6iFkzUQd25FuQSwCvn2rwV3olcjodHJJEDU42
hFs0/Qh+xrBbI2x6SjC5mYHr3foYNHDL2oS2+K+e3AhU149ivAhjV39ipgtXK8WW
dgV5TWoF9gs+zonm1rSgJp1JlWwiywcbm2rGmBDVtsXsUWfPCATx8Bzc4vNjT20k
iCLE7XT6jEAIfT44Ze2Juo33T1vQ4eZiiwa1/dDJi4bcna0cTKhn4AjkQi/FH9xB
JQm8FVWaWynGnRq5bGedKUNeol76561pl1ydAvypk6t2zg0HZJrwmQ8at1XlKqCH
uHWMYiG480s3SxXB+OzC7wdRt+dYrZR7RwO9SBgOQzreDiQXw5sQGaOvqWctEfNC
oCVtkR/Z8FHUSLnL1H4dFsaYdtxm10tOd+EFQQbAt6Qe/TlKiEhe9NOuRUCJ5sSZ
kHN4L/KVOcrYraH6o47DC9wnkmbg6Hsoc9qnC8FF+UvCwIJmtvrPYM1RutyE055P
U4LHmWwFNZDmjHD11ErnrTVhkiSudU+xFoSQM+i5YTzEB2Xlk5Bv3IF+SrK+T+By
h0VHd5tnP0ESw5LxD5i1Hqy5RWksZGbLhexZnf5OGEi89mWJgLzRimrtjPBnVXMy
zSnz9avIFmaGKlGbxA+3xdhUBknd9T8HqyAMDBqTjiIKlCC8zqD4jQc4ekFhLewP
YypbsODd5pOJ0wykOFbFKKHzwykYqLkVuwbXUorMkxtHwAgzZti2jnJiqQl5ttne
zY9pf1HHBHodDTENaKZ4q4Tr3kqETsm5UK0LQpLCs3TQormodYIdZh0wMOoT4d6D
o/txdf8pxqsN3hVpZJ2HEX1Pk0F2CNLkI9AULQ7VIP7E/XFGXhV8XIFTBziF13wP
Qwt2Jy/9o2hgVgNVUNHr2kzYQd3j6nvkOsGcTu8MAIlE4/+GxcD5KKwE+NZQHn7L
LgJJHyM+9TXrUTNFq2hTEuAcy+SuClrJaYURGiXIX/TMZkO1OCLQfQkWoy1So8F7
/VJGmrCSApxheTUykw7dFn3+doI+fNYzAn0PKs51WAd6nRvXKklkORToLkCGp7r3
1OdAIWfaEBq+aZXkBWDSEg2Kdbsgh8o1QM9Gotwhx1Fn4epsYhaA+GD3uoQrFr4o
J/su1HL+6tO9KfLkA+889BJgFTcmZRNCfmKJU9MJpu6RPp8CdilqHHEW4hcEg3F4
yl3rV30HsSseyYAUb2Hlc3P8K0r+APPQhnf6NqGKbUJqQQbYmB+dbIyVReXOIhpZ
nv5YbtnN5ZGQNPLJI/1Tml/V+wxGvtVLj+yG7TFDD+7WHCEWZuWAM4Afjtvp44sL
yFB3yYO07haqgxEbWy+hMOUndpJu+KiBi1q2L7BFHwJSHFLJO9+ao2OWTn8CZ8Tg
2enIBqoyWo1wEIbz3fuCb8aXfEbA5poHCPVsQ6xwG7NMTc56LabVwC1SYzc2AuzC
joWsmA4peOz6CCWkdnOZbViaKCUmMON/P+ZzDp7ivWWEAyFh2YX8Euh3OIy01j0F
9aGPuU8AyB1D7cJoEDf3XQCCDo18zb+wj1KdPiN89nsRtKhcwn8DyNeMj0+EdZ+c
oxKWfIm3OQy4dnu5OA2um/uX7S72UrMnwVlwZRiOrRTDm3SwClU0piZKMyxZv10U
QOoEtl9+kHbztY4POM509yYevz5canIxuWNgQwL6Cooh73aGvvV8M6FhsDvhRumg
6Jr4Dpu68uBfYvYddUw3A/w0V/Y+4FfhY4XXiMobe6kTr3gVAfk9buedf5SWdEUL
Y6v1kbSq+PzO6miL1WKs1Ct2kCbzT6uCeBJI9ecEaSq09ay/hCOxoozi3NUdRNYk
6T+mH1nZePkRRT0FGNXdAF9DSfgCkseAKT08foP9Q7lFFV2DNm32SDjil+zeoY8D
IZOCtKXQo0FFHiv3lxXZjm7OkNIVEgI5AA4lXiXDOijKaac6DRFdl60rtnshjmT1
D3dvI8l4TBlubwxN7FBsRVhVX5Y2c8WmSDNunkb+PQ8LQY71hDwhnZ/91/STA/8t
qaeoxBnNxzX5F148xO2NV4QePiRabWsKO6+DXs0dPqzlQD1Ci0ijwMwEY9XpF1b3
pGmlvl7xm3jLTEnNQ5zKwtUI3U0RPmaWTsXorT6JChjNabnW539dJRq7PvScP7wf
5zZRKeOnYbAkblspKu0PkICVKHaY4kzMnXmF+XWZ/sIEGRC5OpMC1Xvi2bafYzsD
CByAho22/70H9qmdy+brUCVHstlCPzSOs8KQ/hNB7ZcESDTS9QLEygdpJJApJEIv
JrLEViBTLS5iVKD4lxHxkS6bYonzeD1iOuz3fX4Bd+PMdBNf7k1T8njiuEK/kekZ
mKFlAWXEAQx0IoZf1UMQqha+Spi7G99swfLomgxNQ9TrdpmSPCihVIWpUKskr67G
mTBR4O68NgZudps4vqHues31Qgnm+QZkFGS3DrdbzYqvg40bpK0EgYt1MEupC6LF
jBlD3QMMt59waYnDxYifUrcSg1OnwyLGBTRARvZmVm0M+hzqfyIFDV/pACwb6/uS
BwmrmG1LGQ4LPI1Ro79pGsSOajzf+I3wCePnOMDvi53ZAAdtueSH6CTp0vmk2MYX
BsCX8tVvVAeatwJph5yq38rtWgtwKZjQhHFFJlYNaXUKEXJmylDCkXWgHp359Y75
7zrnyhZo5kqjAMtbEv9l1LpYEtrZP/XYW3s+e8TuUo5G5kHxIzSTINrL1Ym7wS2u
XDxbnjx3MtEnthpQMo0C6DLXksmrJUomsCXB10oROkfjUQ8FKkBpJRfgRbu3D52V
KHkduPLcxpMovk1sh/4UBjjfCBip1o283hcLICEp77s/8gTUkDZDrztl3lms2F6h
U9pZu7QVxusevvheTY6atg==
`protect END_PROTECTED
