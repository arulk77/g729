`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEB2s5gnT0hwCOQEmlfhJwmW3b+qXByopNE4CtFWHyDd
QOB5zNB4H0yVtQgEPI+TApW6uwJe7GS2uYpZhU3W0KyE5PgQuX/bxjRcRX93J5tl
lmJA7kmy4zx8Cweouz+CTC1//WTVbJ4sdcMODw61tt9GdvvayaYyop30bSYRkpAn
6/Zan7ubFCbeJTgIYvL7FfS64TD18o1OnFrPGbfTjuw0Pv3l68L2O8A6wlnJmXIX
33XK7J+m+scvVnUmYc0AKcjknm11A0sq3xhKz0cz+BWxtwnDS2AEzlubuec/xwWl
ABIvNHLbEHr/r75eFsedXGHtHo9nQz0HR+8Q/Ix7kWM8nS07RJBmg/yC/nMXgNVQ
7O9CFfNEhKaVcAJr90Ubcx5CjqoM5jyINE2g/FRmkJxgFsxs8WHX5KjzvOP9GXik
kTc2zNX0EJfjTIQlVz3NuljYqvDBHzxXDkpYgtMgWEfNoRl8di/jK9EejBeaZoSk
`protect END_PROTECTED
