`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGUSWYTMQsBHBQFNlbcdUPcX157Yc4HoYsbiQceNdNYb
Ui8moUiJKer7DBFT3Fj6Q8Q/DVq3XSoWIofIIDwLdo5jKCbWQy0Vtxs5wqduV3S7
WzQ3ZVWudtpaiAE5wnil9LwSd6nxnqE0TX7HO4Yo6nCJHO6AUC+ddIy2tGy12AiV
JhEHV0JLDt4OcfZRJPacK/OL9/t3PSNs5QfGcNq09VaVgYeR1W7E53j2uhglD7kJ
pwVwKzZDNE4x8fg22ZeDdeZNZ4FuHcJ3tW7hnGtCyJji8vifVrSt+K4NtkBQBmoi
mQlzdTWS2SUtwWtlDFcvbQ==
`protect END_PROTECTED
