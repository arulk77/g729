`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aT3SDVrJqx4hw6UWrkk1VdwPqDKBh3oPb/vnda6fThwU
kdY2XfcHwPHIIRXIY1rfHNqqqh6kyyXt1KMXiNjeDOzU3lsiCzlnNwrGGIhTTB/n
u3dHA6NA83erBiTPBMoyoGGI6CzepiYdM+6teNyFwrqWb9ZRN9IQy27fdbKlF9d1
neTAwvVMONTKdlKDqh1Thbnkyq4DBVYSkWJIzIfBKVPE4RcnAI/EP/3ifa+tsTTF
XgdzF6Vajqg1YqAMNZTRBVEVgYE6cN3MlsWLJB+qU0e/yUf40zMmDeIOl+Z777s5
qy/egdIQ+cCmmpzGYBqJn6R2b59DJYAiMYjUr4ULvKA9SYVFK3NC4OpzGLFPhkN1
qYshreCzA5cFjB1bIsuliUQrCwp8URFMIxQTRLRCcdktPFgDJrcj5shN9tqJIgWb
F3lztSepHJVfr7kVJGu9sMGxRR1k4C99fQViuRaOISrd7+bpvPD2B7Id1T6GT3dW
E0kpjn7OGe+IP1dsIRnNJ1YgGHVl2taGQZIVYe40JJ3G+LiRnq6dGFuMMhvP5Auq
K8QTk2i8X86da0+PQuPD78wpmjASkwG1s137MJ1EOajaJsJdQwIMX1kZFbaZ+sJy
/ThWs6lcIbTE9GqQr/CH25Q3JKp/PtdLdQw/QfxUVr+mlvDLHXSXDep9SrKHKvIo
k5lEGI+JkEYny5oaIXV8GQFxSlisO4N1DAJBPKx++Xd1xyppHjJnMTpET8J7QNiu
0YNuG5eLlo5gFBqzPckbhPMRalxGqpdonuP/7m5oyBprlboPurcX8HFedYu4tMe4
3kpCh+1kJe7YX9qILpODr9bzOZpveHzlCs02BisHOzf2r1dUsfGOYvjDEFJK72wH
56w527PZ7tNWdEq7Wa6y/8vaXMxlXqnCP9/3kRI/MN6ySM4nXxI7aaZMZMuxf8bf
K2GH/auclhJPZ5zZl5LODU6ZNahW0mI5NXIjkUUrk0bOzWi4ju4IewRQmZG21O82
sK/CQLHSITA372MYriiE1F+Obai296B4QjGCxMdzt77jBqQJ9IjWMBDBajNkWWcf
Iw+HpwaQZI00jk6sbrMJjAhTQXZHUkonYVKVnnZP9S/WMQmcA2nEVmkP28fzdsWc
RbjFtOicN/oYayxIpG4vOR6g27TjVwHZigb8hFJeWpYwpodzDshp8ZUJq5yBhL+E
/iAGAI6T+9MsVz1HT0MCZMu2EHmRGNMBYNJuz4ieoRHhyUg/1i0AJfJ7HWdYbSar
7WU8GluMXyqGMnY/+88Tp1CwtxVkMwEJdQ435yUTePUHqRWe+01UjGYPbZnKixg3
3NtMjk2MExReazEFUoUwdbBQjFKQalFWBHn309n7lTcU31CPFAsiF5xjfes5kZr5
2ODUhTpJd4u6DONC0ZJJ/IL0ziGHK+JK2NEa58glmrwNxWPyyYO05Zt308eUkdUG
92yoM/j32OvWYPOO+R4oW4le3msTQaN4FJjLPUnsWPliiMBF47QBNwWHb32K3Ago
WnBjDNHGzOwuERUhqyLx2M8aOBdo9qMtVzt+o/FwYRzjrKmqv3g/gf4YPb1bFNhk
mMqK+4o5zMWWG8PAn6/SXCApeqX94bQJHDDrdcvseFkr0G00bayt/z0yKFr0XWHh
yVuJSwiBPQ4+p2peKewJcboURAevl4I2sbLjQDxOMLR3yogR6L7BX5p9nBFkdFHK
My6qGFCSe9sJCu/Y2XSxozuWJwELH8Snu3/sspIQsTm9kHhGFbEwyMSktmDmD7eb
tqxVHQml/EMiAuIK2kZtCxSpIYKKyaMfPignEi8yb2BpZfTjWqxcCka6jsCf/PYE
ruQb3vsgiH137OgSpoFnEkFK+OVc89/yN7Rrv1bHpWJEPCbVQopPg4GIclfwKXJT
ve5a2dFFv39oxCMJUF/ASasyo1T2AwBwz7i06zqpT/YghP/pkndJeSe/WoWwDdJG
xlc1Kp98f9h+/q0RXzUgOEG5MYCMUrcSFxG08ukLE1eAokJzx/H9CGsfpCUMPUBk
Ja5lRtsYB0yL3eL0YiUwqvOnqa/xn6c0z4oovy9lq08eq/ijJLhZcTZoPiTHXDu7
SZasxPWqKewA/MYnZEj1d5eV28R3y0AYQTq1Bo/q1ubWOUM7fTPuyx6at0JK5Tds
px/Jh30Tmv6u/KjMmS8G/jMoL6AhoANA9zg1GaBfmNzKN+xal8SRQzTG6qJCQwkc
aShig73OYSK5E2MGnR8MH6L4opOmaiSui0zQmqjGfVBeY+9/IpUPHGYM1sgxuuoE
3Eax1y/mv8PZ/wrZ/u6uenfNRLcYc9i0fDx2MeOSMC1MU0aO7ZMrGqLUoFasQvLS
Uu+nYJVCF54Pawbevp4ggrS6E9m/Ti2B+ZOUNgEYl391z+xMPJm2BXf3qzs42Qos
tb3j2UVSDZ+TMFxo/CeYcEBfi4jbcyw/okuk1h90JUN1hVxLdqVgkp3AAsTX081C
RaSERewjuMPSgrvAkwA0z/LsGQXOISscDWw+SPjKP3EerapNKvs5WPIASrg/bf0I
r+0OfhcObawUW8nwGgITIR2PES2HItq8DQkT4ZrYgUXIB5zsoIt3n0jUopqhN8o2
KdtqW0AIFVWwkmMr1Y1lOTRcWMIv2sysUQxUDgVrhrORgd47o0ZVvFdJh9pSfTyC
CgIuYjiozjNczkHtr5m9qwNnu9Dcv6g+nOBPcX6o9X0fy+c1TymVzCEfRQVtuzFi
sF8gsV+742lAdVjFiArC/4WOMkoJ4losDn5HIHRD3ERUmB+9z+TWLyOYAk7KiN2I
2FSzVZSzx7x6xs5u2NxWSdYwhibjMUyqX5HqwfJIWElwsLlyY9FJi6GcoNd+7M8c
Oa92MohHHtl1Kg8qe6LhfLUiczMixkHWp5nq52JlicRVjkKuOsb4rxSDsXCOCOXI
Mwz6LxYUgYIoTILRwPKpUFaUz4yIEW+kNK05Efk2PifGpUFtLJdlK3oAiqSMBiIw
4xg6anG4ZgMohU1hOkF1DGySXIFmc0SVE/jPKx7IVlrPduK4H/7QDSCs5i/DxJNJ
6x6pKY9p0+3mvpsLHqw8tok5X5egBMuCw3yrbmN4jzneNQOQ5heGyzG2RROB89go
r+nk2Vtut+h3pmc0vF/Tcamc8/9pw4g0eRmj+wTwlgqkrryDCZa06cGv2ZY6SH3+
OqFV5+6F3gx+EoY5kX0/mYIMbmBo+zQI6eTCxOmApl339KwaAtbTM7f+TCSA8GPz
rebOG7nqMpBp6vi61cwFYC2jWwwc0RTDHni6t/XwqoBhafJDD+BL3uU0hQFWFDgP
uSU/VcpJ/KlfkHJVVmc0UIux92ZLrzN/3Rk919AKUDXgrdV3MNX7KBJgbNuXaYME
pNWa/twjRm4ISeFb1vjZTODRC65/VcfFVCQcgCkDv5FgXhOD1CW/x0gjBkEmSqGM
C5s+UgVWo12m93hghvU6AhnkWuLh90T3ThxliPmOjr9siIJBcLQj7s9jKdqeLjC+
XoqxCNhTCRnb2ofjrKfD8wDicqXr45QWnE7/ROUefyiAtl02tYx3MXOzA4uYG5wd
4m3EswsdRpQhodlv71zOYbo53vd2DNKHRiFh1O0OxY6mCwLQLWL0jRjJZ9Ha12EB
OnvTJ5MMgC866lyRsFh27I/MCHVCSeVBFq/d9j9O+sbp2zxscZqACwFpXBl8PVCQ
zzTtoqrOZQ0XTiy89YenHMQCaTCUT/40QSwxSIb0mV9kL/ooVTyd/UuxlpGXiUQ+
ljZ3Ahe4wnUI2fUx2UDCREq5RezGySbUCrahVM3z4JgSKV7AQWWVbIMqbSmQXlB7
HTDtADriw812Zg5qRRu0vjJn8WarvGdfM4f8UgzBqSai3IQGWLiiYoRKw9uXw01+
FLblrVL4mYXn10VDWcin9oh94f40wWZbztKIFfz37gjlF4zUAuP94MKvaQT3c2Gk
hJ6ufkZ+3wgCJPf+GUh2ucGkPzfLQWuJ4QDrcCQ50yhC9jI8UqA20r/Y+xGFpRD/
v1HrXshwv6ZKo1nkiwgtzKbxYhpubbYtuCJWbOMVHxQKtsofuovkF8z9FEAFX5Ob
LVdPvTYv1Mo+rVceN7LQ7EDIllRmFiyw6Mc7A0rPgGDiw+/X4m+Jxfsh9guCtNI7
5MLhsfnVu/M1YOpSPRkw9UqD3uny3tYd2H+nNjM5WsazC+2gr1Oe/OOE5hHQ+DZ0
GgWI7gwbyy0TOANeIg1wlEKFlzoEMkRadUCY/lZPbSWF0gw1fY80lqvt1dOZq42y
+NMlpWE1QIGPF4CV8rQ2d8NWMzBkpqQuJoqhzwOupGSDEUfRAaXsmYb7NKhJeQ/g
xpLaB3vNCuLfiuZlCNJkEFJ4G+/QFdSimuQzHOF2eFL/U6HmtDPwwMIcn035oXEt
Ig15uRQZ9FuxJWL+pa5QUhhSPcBfRQPndKHWbMhPG0JQQiS5O8iFuWh0+tOfkRzH
iG3oHGpzsUtGj4UxCaE/jatLCrIBeY23wrXOS3gfDqmmlv/3oa8i5kzUhvU2F+3U
rAHayy/H4yCvmHQE+AEvUQdTI0AqgtIJN0akM+13/AaTZtFkiltjkS2ZhxVyir9s
USUNWK/VAv9G+7iyMEwDzIDt822MTSABsilfWskcEK9+tg5DVNOrLkD/yh8TXcFX
WpMY8BqbO5JROHh9ld+qSIa1xVC554ITNVf2oFbrQxcETn2ujUDSanjHFSDF1cqk
BgmBEKXOOx81r9rvpbaiZwayozpc+XI441p4NERJkJD41gpCwjtwcFiZwkFyD7CR
zRiVDdUGT40akPxsSJG+C3enpBYwnYhAdeIro1xlYW/zWv2J/LDLclZSCm4YMU4H
PsL0Z6yObmJcTRkkRXYn8coAUS+p0y7f7UiigRIFO7xKszsGTyVsZ4vShWipPIzy
cS1bPsAD5z17zhCXhzKAv1vySm1rdWEv+a0cNRMeHQLbPmYvLSptvnt9yFpiNvuo
k44Gq4pJTqN7b20feE06UTfLNa9PGkBuMRCAj//91QUr1empP+FSbaKLbyW/ehFm
oZEXVeHHZrH9ygEjvpy4rMsYmGZlbTn1ke4iflIl3l0oMKkMQpFtRJ9TPk62WFH5
lAX/jtPNn+drcPeZ2dqKhdIpXSznnwVz2ljAHkWz32hWUt9TOFUzgxgzzjWqESMX
gfI7jmk1fAiqzWnkuwUd7ntdRoufKxo8hA1D58SZLhsdslJCXI5HGLYfplo8OPAz
9s7Kdz32l3T45AiUhH3lwDELRLVYFB7XzAIRjsbLBkE7K1PT6xnCtLMoSh2vmjF1
zClrXuXTvcxHOE4r4fSgXw48RFbU2SOVdnpy/7w/Hu7ehPKpj8MmexOKTjgvcMOe
IOYzrill40nw66G/vUtfQWKqKbm9vjSNXNEeI4zPsu6Qmv0MHImc33hkgXOct4ED
RmAYzGOaL5PVnO+Ui/VFUiMZBplkvgwV9bn91k0euEtxq4ppeSgZUFcBwXF2p0vH
ZSAPyhGIbs8cSwe8FdQ+OMzXYflZdACIDrQ8bV1c7C6++wGC7QOY8KG9byK1ASsN
/6CA1B+0zYLOuygOYtCUAEZpCxglknUYltKLk8RW2JjTkOHzoRGiaj9uBss/pBcv
XhHvlo1RFCOYN/K8aOw5RnRz52W89/8eJent5vlyaLV+9MaRu40sJ0uBfSj29Hl2
qysoccfRkqBZA1Ue+0fdvByGNZC8DvuG/7J3cMvzHM9oj6kQo+LN3jH3O1/E97Q2
XGZyLqRHcYySDXxKmVt+E3mgpJYhhlbCFnu8Q0aSW7IkDjt0jGk08iagRLm1ub9Y
1f9cu0s/ygO6BvnejgGkw0vpB/vdNryDBpik8uR6DiO5Gx4cNH6hTtucDzwyIopc
T96BUf5Q+7kxCSOxC4M4pyAwLz8mkWIIp0eiUA1g2TGn1albPRYbQZ7qCPntEc/r
y5rTNWeHKqSw+dgxxQ1hYCzHSe3S62qDceLfDwzb27dulfzvOO/mB5f9NM5nrWxy
hz+ZN17G/hH0llBGsdgo4jJQNs6E1Qb3Y4ExA94xiUMss/ypx/5j4G27ajP+TelD
kZCRWdH1uNnhwCq8gbx2kAM2gBejikCc/gVqIUQ8KpYrXVlANOpEYniVf+Nk5bju
7QIuV9VYrPw6EsuX8ApXsrHIjhNksO1UeZ6PD+ujIt9L8WAMTuMxp4Vd2JNhi8PM
x5sPgCWmkNvG2qtssqCnD1VbUOZVtQYHLEQlWLyp47e51JZ3KWG9q0flTQDBW79U
2DHJo3Ub5qd3tHKoL78DsL0PJOP2EbHhZe3ezM1NbLSmR7ucmPtZQg28QrvrGuLu
B/o6PYINX/aK4+07ap60YFUeUa4NWh6XqpMAci0IS0c6kINjGWLTAyB/PTscd5F9
L59XF6wDOvG2tBsOhVEr3hiI6cQiFLm1MNfDs0IJYa0TUl7zglU93JtM8MyBJdEM
X7GHNd2+yWl8L8OBtiwhjBHahVQkUEhe9Ch1AK/f9SerTyY1s7jk+UiRftDE3qIw
ahTsYNH2iInsDyukhDGHLzYhPZE5l5Ae6yUFC4eTpoLrnjiWZFp2opTDDHYi+xps
cJuv2Cce6HIidyNB/Czs8iV8QG79xXN++Y9kWpVocZGobUswZ49/EOAVGZFjcQPE
R5lPbNjRhXrkiZWI9O/VEzYHAde0Ju0Bciv1d9aUDhcFvCy3epNLVas7cX3JQWJi
yqgeW5ZOg4CVdVx5O15HArrs1xVfDEU8yq+44XuiBLhOs768LpD4m9Pq4HIMwH/H
nUuC5cUtgnHkU4Jbxe1MgaHUX7HsZHs4X6wz981FjUd+JUmq2GK/uPZJQ3u+Nf0P
Gt6EQ9+hiBqYZOR0wtcTuL/kwOSN/TGCJKFlRYcZ1g6A5lFeXgFBXumLXiYtaolh
/1TVlhcMVxH3F/IxOe4n/p9VrCslaKDBDf+OVySDu+EmAO2hope+tAHmUYsHAhce
hlmx0qyz+WwXYSGgZD9rEVRAuJ6qevJZaAAbCPJIA/4eswKc3jHTxWcy6w4iDfp5
o7Szp/Bnhtm0A2EWRP3wLDKWcouZZPWHH2dWzFDOYHo+H9lwUKWaMEAACWyohD40
85QF5paucV2nFJQWoLA9EQ28CsioXf31FWxU0DIWGJbppYqnCEeNynSHPsoATMBS
x5EMTGCuKDF+FbIlK8ceszLA5aBhhPZFnFmim6M03LP4m+3lODv4xMZpZk1KUQ/U
e+P4x8UL3wsGY3O8ozJTWfx37hvrTmgm19navcoftnUqXj1ih1H9qQIcSGApa4WJ
kO6TJiKM+S3CLhtBE4M1ZlRSO4GTJiExq0XGnOIuhS95LomHE0ueqi8WtGj6GbOo
EQNjeqMwAQpGxIkgCl4T8LlIstjUMahymxEKFIFoqrpbZFCv7XD/WzU/H15a6RQa
weYAn61yRKHOCaOy5f3SfF4JmoHih7P2iASfclG0JudFBppdkOcGxxA5fVSwdcsN
vRoTs3zmWGZ0OoVPHpr1GXc3/GOAuQlCNdMY11iJpBFMsgMTq96RjAv8UPXELYcH
8EEXux8lAoNRlAcI3iN1UBGDl6lkfetp+xRzq5bprxlw7LdzrDH6iXkVJQTAcvSz
0keiwpD6MSVt+6ApTIg61oOWMDz2beI9xdJNMk+F1z4LOKlzEenwwrd/3WzWzH1M
NNk69VdCM43tglqkT2i/GJ7M/yB3tt8YFZiAcriDEr4Yy/ksNcQlIetJdkH4zbxH
hKkMEYTrvu2piX/gVJoHHVSLyzMBmHxhtdn5h1MX3lkl81Eyhzm2Vw+a6Kt5OqjE
HfhkSBe32RTfpZqtG1SXspwvoKsfIKstk+FcvRsZnIq76+r7TiWh/pLXTYaOU5r1
uolI+niCJxnnbH1/tmLi4Fce+LUG6ZJa5lvSM8f7OY/5vnOHn/GjWhQfy5IpKGZ6
VIWLTdqYAR9lY1uKHfF9cspWuSEb4ec6tZ0mqqVp7ZaBSFLJEM10YVOuOSbNjo3r
N9Qr5wIGbg7EODI7S0NWylZiN2idJgMl2c5gtumI/YfAYwnqX/nQNqLxlW2pOIEv
QMuHxxAWUCGkiDV4eJ5Zb/vCSR3eVvvbEbxv34QfIUpb5Yjrhuex9WAVyioG+lBh
gLIZYyKbs05V3gXfQKEBCX76xYzSWlJNMHk/cTpcJ0TCxVxmJSnTFfHX2jaZDz47
iHrFWjL/poBWf+KZPCXSbOv5rTNHFJ/jD0MvMSmq+DmbX3muhNURCn9NtSB/lh9A
p4KDMFq/7hDGaZLYI0z7oDuBcTfvBzfCQtJJ7J/9MHobjbg+/V7MvS1qlRnMlpxU
gedamcDnePvUJowymOCmXlQIjjEjzmeBj40o7xQT+6W4QfurXM55P/2y1LzULEsS
0uuvyY5VjajnapdLwZ6/w/Nk4h/eKOlMULuIRxkU4v0QTxeLJdiuZ6fMcUKcVV92
9J1wnoVma/uMPoBgZ1H8g5wbTQBaHJn9miyxBb+3TANdC2eF9OMKrEvDw5Y8g76T
AjCLbe3akkD35Tj68wFLH6d2PdLJJIJ7g0A99hIEBPI+DTp0/zyv+nb4YGWdkJz0
uo1HepHTwhlCnCuC9dbtdRZTV9IIep/gy8Yx25x6SZJJUfy+FYNj6MwObifa60tk
+Nra/WcWVeqHfeqSvV4AbpcIYEAosqolLLUoSViCdm9gnPlhe/oaut/ZuJ1RHZHM
OoLNTsAsYdiooCHB/KX0ZGqs8DcnZCoSaUCdg0eCTZ5Qshp0fhi6uwZZFpx26tRL
k2ik3bIi5TtLYxWhLdcnFrpDYi90fYmhCdf1+4OlB+ms4weZZjP/BLbGm9kQC5tt
3efGuGkacr0D/u2qfvFLPEuccRq3ytV5KLBQEYVJLlreMwVQ6Jx4hD14vCLW7W5Z
g+gAZHtLe6p7g9lO8EIDGqNhp/xAfYlNtMPp8RG0of3bvI8kHXPc2CIbOy3KIe8q
0AVg7QUYAch/wQLcpTBXTtHCib+k5hQOu/+g0k2LFyNSPSRyi/u0i5ZwN9fX8XTU
D3L9Q8HzNCaABvnyypvhJ691IEpMPKH56SQdJjAFSN2hrQAEkiFwBVc61f1vOcTr
HKgvTcNv9qOgPNVXHs5bVeHYjjgcpikbWcCQSFbnMSqbw4o8+MgRSrM9wTOwM0V5
/OJLrT8sbqnjRgltkuunripTKEWVOArzTvNCxCmBP5evTRBsllbNPze2UUdlb91f
JCaeh1QwcJro6QuRI73q/GgogjExYzg3oNH9N0BOCVhVI1nz3LOMZ8EXXw68hE2S
3Flnt9QPyYxRZoYSrfroAfm4gTnJsE+Xtp0OPMPBMVfdcNMco+GGYPk2VvY7+rP7
DoiaWy9gw+p2exytgscHuST1jspuYs6uip458NzEjxzcLFbjxEy991fakVinfGkI
e+EjnF5ejooqjwyv2nt+ZkwQCJhxl+/TH/GQ214Par0BC1a8pu9ZOQivra3RctUz
HHT8WGyOJB38gswVy2ORAyraL2q6bJFqttF80dx7aerw6TWDUjNrnboPiZbZz7gv
6mqMLP+2Ws6us+L4s0KU0dcXvfyo9hedd7iFNNaGAxOJEjVEhrt/JbOIs0DQpI4C
ANZ3n32f1FCcuW3iB4aZWcP6ofl6Nl5NcaVLSBeiqf/vFY/8mlF0ZI7VkYvGIcYl
gf0HVShOWZ+ZJYCP+MmxtqXMeUQ4MPp61bNlb3A0EFYW3/ckPA5Lsv25q/oIdL0O
tpGNy3RxttmI1LLWhIgXkRvMAs+ZrNrWRYaZI/iAu/KM0TLaoz+GU9bK1oH+9U9T
rywotkejV6AgjiOuRx2RfSpUvPUX+r7er4G/IRbgQDP3wBsOyhC9XuTQymx3sRXp
mqHnYnJf4VLhzkchqb6BBj6B4NRxh1Z9Q51yUYyg6WESWwt+PexyAjNpP39hNc2d
rKkRqlhNTY5gb4WGFrtSRHq5D1RNum2A925jgrRzRld7LqFL1kRhLUmsxz3YmYZO
dE8o3DDmMD7SW+y1tR10lcWmOYMKYv9FDz2qI9pBMBsGEskJeOYchHD1MSXbGyle
NKKLvBzfLmcKKGo7xWVO5oj6jVtKSGS1LiGDr/+JIukBqZCljLjDcHGion7GFcrV
WRtzi17l0cT3SfM4qH6LsIclAaDOkrr9eSGJcCrpvrutM1AAar6XB60inmb00CQT
aMQSpFNNTPh3UtUsjPHIGIP/g0+kw6u3nKYQYyg+B03rSFJcZlbtwlsQcWer3fnw
qyNJcGK6wgUtxAVgxKC9ZuX0ih9S1DK88+RGZw+MslXBfS+QgA0ygKvxFb1+28T2
1MVOtXWuAWlVoKx+ZPmUi+KBdpfF6/ZIoEQoeIi++ai5iIGYBlbKfMe4P1IHki29
UNwJdhOqieySD2KrWVnyGCFFM+V2/fecnto66KuCIRe2CdCHOBaswcgFJfNCGpOD
drB9eSZi65+JclC8AElC8dpuhivyESH3RiZwmNxnqroOvS9FtJR4Z105sgbS7LxT
8VlG4P6yVv2rdGiPIGY3wiWI8JgSkYSlirWUMUyjvUbmPgxImzKSKc3x6ulZ5OwU
Mv19HXDJu9XZizezLlB4+Q/jNptSyqqyWACcaCkrTc2JUNx8eUb1k/kk/0u/IxSG
55jkeC3Th7VKiYlQltPnnyd8jwGr0OSqcFnHnFVpx3Ntq7sXpk8AiJNECsaJl4iZ
MwLJt1ic7018B12lNQ7VoIrVD/ZKdGSJ2/rc6Vjo08SAhCkiB8ytPvqlDFmtqSV+
wN2XXC8m/X8uJ273OvY8kXN382aFxvYO4Yx7pWG1eNHaexSQtK9eISMq8UPel0v/
DF3TW+LQorByN7GwEejhQzJshg2STE6w8nOSDzoZ23SGInQSCPNMIGYXzKQZwITp
2a2hAcIUeSGrRo37VtSxDT+3RN//z20kCyAe7nZBghymejS0eWuWy/vCdHRBPnsr
mFoUycyU8mvXUfI6zpgVdMZgRVtptPUOZ/klAJewzA1ZCI2VYI9yx30CPyew7pm/
6SUYdrcOHUubR7Lpj0xLhTIT++HhwMCxh1ZJONGt7i3N4TgS8/eRs11v/TumccL7
CrzSocoiqvunvDiPCRpBSeALZM7daI7A6T5PbY881EDm3Q95fRKN8CcT053Tyy7f
FljQRCnTWYsnWfBDeFXWmrDe3YlFNWX4tAINoMlJm19oNhNjTZepGwz7qiZCt1U9
lORAl4iQ0d5a62twgMNdmWK/6A9WiJ/IZrzbUItD/Fnwbz03DRUkxLr5QICGAkAY
i92JVsIJqRCDA/hxhppD2xxT2PMSztfZLqi6ReuUsLFFO/69RcIJKDN7kNMqh5gN
N7ODdUeN+i2hzkraVKX9zrl7d0Hu4ilooxryFVGfJ/w385zIPCK78X0kKNqKvUv9
HS92Q49LJL8GL429AH5ZIbf9XS+ivQP/r5AVwJte20Jk82ufOHlHB6IhOmB9/EhQ
yJKlZT8b7jbcMCRBgYE92lJI1oU9VQJvnPKJ9DMMzwn8slSauo8IasULxY+Jd51t
MjS4h0J75faqVv2AgKGMj0uzPXtbUNwEiyw/6foT82KBvbG7VUe2Yh4R/lN+S2OS
SU3z5ilLHjkEoJiDIkBGmCdYzVkX3oe+EbmQGeo13wpkQpE6Q4m/0UshnRASHtl8
nRA4sNnWB64J6uP4BMndweI26wxGIk3og1MYi1Bor1yzimop+3fCg5MRCEdevea1
72ZCZuGDdrOtV2DYfAaEkGUz0TpzJNvhva0JcfA/8js6EtL2rMkc1UZt0EN2NOnS
oPbf5HrRalvRitHh2kVA1rCz4I2TBEHhewnjVUDqD86nt5NSbzKMHG3og/PpKvil
hmzAVxQKH1hCA174gOiUSSdXKRBBgW67sGcRfa0MBje9oymIizSeEzZTmtpaKCo4
pP6X7GCuNSA2SlUV1GEY6oHnh7KwXvbYBY7COCsuDIH4O+ueoWUlKlrwvZ+msvwA
kfwfEG4aGSu4UO+TGOvT9/3kf2KvixxBAz99+QxgcXZfCN7KgRrvaDyokTg2t48S
HHle30nxo6JUwq8ksKlyC0jAwan21BKRh+Z7T8sWtYIxov22R/byWLWNIpZETF/e
/cIGpozbioaPAMUxkeB9woKlTn6qs8VGYekhP+5MUCY=
`protect END_PROTECTED
