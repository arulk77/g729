`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM+scDjLsdqYWIM1uWgdxSTZE2OaZzsPzAe1v9Tlx0Ik
euFpn2WB7vCvcKt2Don3pCG+3zHYtfKIwLnbhWQ2UO8M7nIc9gDINqrMow8vvqpW
244cMDt2Bp40efigeKnZSfMkPnV4Mjy/dfzmz9bn7moZAEsicTuLKCtV8F2im7Nk
0d6hzvueeOAzcNfYEtpOorOQ1gy9QNGvOLrMj5dOX6XGX3pkoI5K7JnENS2RSdwy
DbmeMK8kt8wejWSfpZoS1ZBZumVBUNY5PStOVpM8KjDBlEP30eyh/OivH3OtNQC1
lQ8QD1k9DB8+1lCnypcrG2fXzXpLP3huLsPmQzMIb5KxLU9VUfVyVlKWUviPnByr
nScfgSZOdZ1S/YkODdOwImwVIkdp1ediDOMFL3tJa2pj8m+fL8tsOBLBAIsu4jvc
oXYfeAL9FLIwEUo+whC8uAfm6XhZyKJzUSA+UGKv0FM=
`protect END_PROTECTED
