`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu497VqqLfXnFJNjskeNjZE/UrOnNQe804AhxsTyPCFjEV
wvw+u932omHOaQA6Cy84bKBVdDXaCTxGLKTKmXlb1LtIyIak2z4KGqXLEdw1HL9V
A1ptKfx8HtEFks+nDzRSAV5ONSYGYfyIpM/gmyJz2NoriMgq1OyfuN2LmHSFT6B6
Y8tq9CcD/vccI8gwCKVZ4tZtiBQGaehhHTr5FwwkNe2CrHwIi1B6+4U/DqpxTM43
75D0NxCpro55ORgMl0oMbn8cSF+gdh8tjtdMgJg7jt4M1x03n2HVM0zV+VrKYc6e
SvwwhyZ1OMylUmKwPOxvwqI8vUGTh5oj0FnWgY1InxWN2oSCcYeqbBPeaIQ9ZbVn
rxbVNehkF4bR6Vebf1+lKA==
`protect END_PROTECTED
