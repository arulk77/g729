`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNMiRWZChNIDaiB+HhD+o9gWaLe7Ccyb7HYp60cWYKKr
3+Tp7d1AFT2UrFylYNgCD42GHbqQbUYEnp5f+uywv+X4fG04FzliWGvmkMn/ZN22
39OXBKhwj4XOpPSxBC2sPNCfyEHXZrOn24n8W3E1dv2ZzwRzn7V1RrLQgKXa9kTh
jQS9sj8+AYVqtnWneiBS1nqDXkiD38P9+oSnIcx9UMRx+sKE8azArvfVDTgWlLf8
zGU5Qo3qdzs5YXtFP7DLJv8vAfIpVluLM3E+i8oGPNqag0vcunQ22T9aLRAP5aWw
MlhOPKNF8pr0ESq44wGlpdNQCvOYo+GoXZ+rUxOGkIsZsGkH9oof2fMCk9B5cL+J
PjcsVrnFB3zEUrSrEoFktwFzR/xKrRmZXwPhKKPKICJQwNfZxIENDzsWRUAuGhjB
DmMwf9mVSNiv02Xb89Y3gaFdb+1oQ7fjdD5yR2/jdtJVoRLIl5nUZDpxf/B39/rT
PoX2cjcGes5fk4e1hAm8pGrJbflN45A1XxpBN3n3VrsIPWcOd49vy4SoFIiU1fLR
77e7ErWixICCYvFnd3/4UMHclmFzE8OV11uR5iY3kyogaTHGDlEOpUZsSlbXv8wl
91C8J7oQbSdIeCyfTyLGk6e32BrennQn2rxTYTDUJ2ONyKosh4+XhacqEt65ZyDw
Is7dYT8IO6+qVDGqyNEQTLZAlcYtMdj+42JSgqk/KQftzUhmYYbn1gWCA8JEVBvg
8b6CP09LgOPa/hxy/udePG3Xb5jjByB+DIVJz+bLjF6NG1edsNwQnEjWtJCtLoD/
2C04lPJYIGOYXfYhx2/5zHIz7lB+oKsHx610PFlRT7E=
`protect END_PROTECTED
