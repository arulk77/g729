`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveERMc/Xkbtrjp/3yhuWjHNbNB/Y88zX68PbMwccrJHd1
MRDl+dXoPzwHpfLrxlbSI2/qcz5STFjFg+yrnq8KPECN20R/6xKONi1NT4Q7iUvg
ioNtF2LpHrDakwOkUZnA4W6ONBCaLkfaoOpncMDWCzGe664GdlaQy4hxdvGRGRlK
1jLxKN1eByyzU+7+aWxzAUcNWe5sZ9myssd8nD/5wyFNc87PfN0TxdawzCUF6AU6
`protect END_PROTECTED
