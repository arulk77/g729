`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCtM8Yoby6SvreXDfWiPomDa2npG9tC5OmC32sOHIBxq
gRRG+U666HSirmFpFKArkQts1jIxMd3d9HLHne/eGXx8S5mBQ4facQcpkWKvAWRc
ceGgiDfpNA6ImX3A+Blok9fHgXaLOuJ/YtwYeW+6rT0JKQqV17BUi6Li0s6f+OiB
ukTdEyd0xWhwW3zlNefP7FXZEvYhDArz4Fiinh6p+v9BGtxpfhEpz+kIKtd5n8cr
`protect END_PROTECTED
