`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SVVxL7xHNxAyV4F5MtBgEkPHyMgLH+/RWck6dkz4KYFX
fzIsA7kW+RNrk/TkJ09J+1o75rYkbJ/GTkmfwjWbqfDOILErNpncXd0KB/guc20Y
y8oKGa9K2MnIir55h8GY8nZ2birXFldG8a6C2caDX1/Pl1Kc4SYDTjFMxYWDUMC7
mItBVPhD+47hvKRtWjIx1SII0BnGrqke8KYFP/I8NwgJ1ohFaC+CxVE4RWw4FbVt
s+njNe2goMiNJ3HL4lHo4vtwjz4ihmY7aof6aW7wSEU7oATWPFjg7J/ZbUsNotvH
Ek/+wl8KYBxdDnvdmExFAqDYXAYaEoo1+6psNG2eQOgOL6EYWKTXeerG0JNPo35O
m5dnmiPRtdz9u93539LMW3NiOLODqFnFqbn1YmyjQnfa+joRUlr8mm04855e01oM
9tI+hnvslzh4150VAc4gn7ylcwU5BpInkLrDlxiVi0AYJfDmjMxNiJtMesDvxkyq
5JUEelUE9La5g3M8AvP2Z1STSBauLG7bBasqMJ9p7G41nFiE7g1mRCwM5Z7IxvMD
w/hil/756CpzU/R/N/mvCsGEpOKQtoceTQ9C8ssfvohfkTzYumFjjslrsyhsK4g+
wXOUigfpA26nbGh2PuJHYRtX1WxmzMgsMsrE0bw/9rC4FmXfDlk4vMFky5wWrIR2
KOIL40Afu2UXzzY08B+jn3XOmhBmIuBuAqilJ36x8ZuvnBJss8lLK4dqU6vGfhjH
PNe2aPn3F4wsXAhtFmXTEqCgu3cOVdpscdArzF+1ly2BxojIfeXbaz3OsYcxGZb+
oXZk/ACUeVhOgd6eUs9hRwxEtaPSen4YLZWyocW6lDKCMaz9ZUkYYErleVVhIs+b
uqswKbvLpJvTtSI1WV09e7zyd+tKzVglf9vfS40vXprslolOvclcRq5JnldIxa/x
SGju6eTjjHEKgM8mBjj0yrP+s+MJ3qmrEp7UZaARzBBjMBPZf8HmMaZMhhhlh1wI
Dm62iuEmyopOpZIKEzOG6ePa5suNC7O1F8FwJQv1cR0m+lL37/mgXESiQkMM54mU
NB22aXcRHJMOgTOHTGRvOLYy+rhTYwcb/OJdvCP96c1Hy5KpNt3eysldSXyBP8vv
4lDGPNm1lUaPedPNfctkI6ohbK98EKyfXuVQiMA11L8auVvxk8AnA2lPWkqt4hXe
3Xd1pTzBpikvyLGl1o0U1bLlv5VR6dIn5T9Ue5feZVwH5sxl9Ktjg14Pcn9hlwPm
SWOZaeaJ+SbSafwtyQ5il4KcNdGDhyE/MwI+r7eA0vbj07OkuDKrsJO1wZ9hxIJo
MVsEPuV1PhA71N1J6D2Uq9by1hO4BCaqwBhfyivSslleFSf5L3jHbQdMMqamefjK
4fGn3+qX+KK6thjoUMPRU5o+jXINRsdZWtGVDHyFbLPO0SPneDmGADdOZJwE7wHh
AIiTHMOF/RAtW33N2ygk31cAcHjK62F8Qv+I+X8MLRs81kT8ZPb38rczgSGMlURk
9ZdCls6xRPLQe66geaPMkEbXsOpWaHYnOC04fdNNPR+RCKJ3jO/TG0vsfP5QkR6X
hHef2Rr0XBxOnje+HbwHSIgqo200JTy8HzncXt4ItrMxlk4Z3cgmiwqSeH0vXpeS
nFC2WU3UOTBQgkkzEEnM1hU38Oq+simBeoljoYjAfuW7MDevLXW3+/Vg46RBxqIe
C+IgsMSMBhEnbEOfmetsA0pt2oqUeXbp92gj3zTtIBt8jGENI59tnS5zuhpbv0Dn
IMJ/RkcsKpg5V72Fz1wllF9EH3ek00MIxYQYwiqpXKVDuwU5A6NTUZGfgkO94yBz
NtlciC95Mu5pldbRNVJXvVLwPuY3vwioRFgCW0/vVpWwJ2YII4L2QPlV6YBUxgUK
Vj71U+nCT7dHSu0wg5I35yFfZ1teQ1j+34AXWcJG2wNjnKlwhvTwCGwVd/t3WTb0
KKNjaDY2OfWyreZl/JN//U2PCO/r+b/J9O0bjkvt6O/q4mI1TGZN8TGEYWRg2UE+
BsMtpIRIkH/Y39l8WDUEAWTA4BZ2K4JWa301IfsmU6UizgJ2CP++JyYeK1oVUuJj
KL+CX+/HgBXxtZHrb6QVwmErhNbdeYMS/msx0TosAclNZq7YQynNgdOAAwS7IWQV
fgRqeYvy6Z3YgzHU8Xot4EF9ZLrYZUqfTjo/J6ai4LOv3mUo4JgexiOLZtNgwkAz
Ix4/f/I3PlrCtIgc7T97wDSUfb21thYormSM2x2XI6g5amc2U6c1Z7AuXoQopWMm
FKPgo+Uqyn8P6NHm7KObAhhLPU1IaJm/RbC0K889WlLKzVekG0mcINmr8qJSKs75
A407pq0jVNtgDrrMAV7c3SdLJOutzLTJzXvfLU5h+1xBUmWLi2wch+A78aS+FFCz
5lTDI4AEb3rVS4R7XIG+AZRz9WAFevDPKp3i5vcYneVaGuAiurktky8obN/W75fz
GV+ZrhKKG3mS6+bhRpY3804uR4HBDmxWF7OKCwGh9ha8jJKotPLoO+yclRWh8MtY
MmFIInkHAVKgA5xrxYjzbHh2KdMuV2duysyCenaqOL8LXHLwFKzvmDg9niVLOENE
oHTETL1upllO2XLjgILam/GlPscJayXTWRUOo+QM7kVJOeg+YPEfkCYREtE3L8BT
kJjBtD0asV/B7Y0wwOv5hNUXZIM5VJK63ddm7TcHwKkLHuinXNfxErR0hgDovUhu
ohucR6PKkz+pyVVbTRVjmIX79EQ8WTyFTsjdZK313UqMsEfwGaOGdvRqvpdw97EV
CI4USgIkCw49EWp1qCcjyj/3brXVIJ+Djgj44SzrF+NRu/TRUEKiPW10+IInNKYE
7rxjatjf5InTEtUBT73pOjiADdUpokxl3SoTAd3F8dhPMmADj88L6+Z76L4ch6nY
0VUjkXo9tFrAKKbduUHEYXRTfed1gjiICnlyvZ06qFrIRIfFI1rwcYt98pHbppl2
thnXQiYJQTgHKgj3Llg3lGeGVNyyBc0Rhx6Qm4s0MYtTtR4mSrC5Q4IMwnZvqyIF
iVF+fo/NvS7Om6MF5JaabnpHNrxt8sJ/S0hQRuqj2D70kykLSDQ4hY0UwLz78swW
+sXPJJsaxdGZu6k46TDgjWgZj2odk6i5VBpod3c+K5KTmEcv/Nps4bl7pWwJ573s
NPWI/XtD1PbuwEzExgSSodQn5kfJoW7llpYXQCaF8xJI7HZeQY0cu3D9/ARyAw/d
8FWSGsLAa7LSTdLufZh1KsAfm646O/gSTIgOpdQiwzufQ8/THf8phA5QLsa2qHdf
sXp60VyPEcN8IJLEa0Px4ft7RoLX8xz5C+3nD/1aTsboNmb9kb+8L/UWg2e/miiz
Ttkyk0F7FgrjAdYothjQgx6rh9gtQZyL9zh+YyG26iHNsW8EmNh/FqDoCXZbWOtk
I6vViaMEhG/mCoz1r4HNvKVd7Vx9IQwTb+e6GJ3Wmd6QEVogoiDlBtic5zj7J2zt
bYA0V22isFeqKesl1MSt4N4DILRg/QaWvBh69u+U3wikJ4QAHvC0/yYRbZZ1U/1Z
doXdLducaR1Do/ayqQ+WCHemXswwPICKPGita3G6fcZ7g69YoS7Vf0nGtakJ5BWr
mmpoaqe9laCLKmx0EEEKYInpXjctKrlFNegJZ4XVKqO0Brh5tBtosc+7SuodP1MQ
FDYmXp4f9HMTQdalAkJAng8lUur8Tx7wse41aaOuMt5cItbqPDfMGCCcZWa4V03z
KPGMfm4HfD0HCyi6TOStXhFNY6Lypkwkw+pInPzWZZnw2Q0MQ8LW0sCjwld6xAx1
rlUwjDEIBkjn3FWU75mCrz/i4DUllEFjNYytY83clf0MdNJqhHWsdMFyQOEZiPxl
03Ulf58fQWfOgQf8wqsvLMKesUfGZ2RrakTb9V5ctWbPmo54Ol57xDxzgYipGG6S
NE/qf8q7UVtmGakEMCThLB2OF+tFmH14FKGOWZVdEJN2V4rDFsuNZMCqAZM9uOzn
dYnqLzdsLFd/fVq6oE2tfLm6xiRS7TATNcF7JOgQ7Zf/Twp/SrA0D134XV5vmjr/
9lKmCZW5l4B+aLKcZPnfN8kmpW2KAYdZIYx/EDN1iyos1s8O6r3J3HjnLwT1cJ+2
06Hol3+Lz0qIn72UyFfLQ5eV40ewslUiQt5BmSvr75ODYV8M+x6xpn/XI5gznZxs
zLMsumDJcTshMZZvK18yr3IbAsCDnbQG/twHZxoqadtm4tmkAgb0BWZ5yUc/QVRo
jjmZFAs1HqsQD7iTgUuSgZDag0GacXo+WQ2eo8nQ/jovZsYiU80ttxnS98CIviCf
q2/PzF/wBo/hKzCr8dvJFJwuzgOfS4xNMWmVBGGnFEn1fynP/pCA7Q+cvgKojsya
+wMoXuYVdZXXP7InQ4DdYUh91TnzHLILF7s1TGz8BWvXLvjicwdSPESJGJ9GdmXK
ipBtvhGDS365WAOmuINQKPxUUFv9bA9bBfJLiTu+q/AX6+iWfh+hFjUxqBq6aNg3
IxWYINZsvbtfg0mpX9CjYu5s0jDC6unTzjORp1J4cHCoMSFoEYnOwyeJmiOXhGi1
eXd68GWwq2s3j7Xg3IAF1XPJSsFTR/gqXniq+0T6hKFcjNt3xKdNUI0MBn/wkqNW
7APYTimoyd85SQsqLn1rrGdT6gLZXKczC1ZYkrcyJqd8LJAUnH+bgNJGyHS2BJfL
lbfaxmItE5WhR/CTTzP5sD3SPCBAcZ5Wc+L2j4hgxyF6KrzFzr2HpC2tNniw9N6L
Mt5Laly8Lv3LXLuAji7qfFEDR4WqNCWRt9Q9lNpKjqI943bA2tlONHXhKfH7CY+U
djWnBwWfBHU+1E0YJpXK2eKTKAi6fbI+Ci6QSMIdWvSDpA3i+mD5rJAfGTj6G5ls
YAC0uKkcXVe7fcO27VHVXG+JipKtWkShvxjd+6lpt5cMwG2PUQxqxnGAI1NnfkQn
x0J/ucOdmiQKzVg5sdbYOOce80rTu7sU32JeH4uOiSRKfqkLHeKedI8hqRkrBB42
Cy/wayPJE1/3Hgsc5Nb1NEW1w00qfHpGTn8rIx1IcjiePllOEVBZTtwBQL+FDZ2Y
SNvYwEgy1wt+eVIPujxPJ5o4cI7X+LtfGUXmRI++YwZOkSJ2PpEvZkmMm5UAII0W
B6tGkwb86VMe1YpJ1dS1N2popvGt4l3K57jidc8g9FrKcoGQ8s+rVFCOJWrTqvrd
eExD/WgKNVW6Qye7amgPThzAV2288nYGLrbnpyGn5NuUCvDRNW4lOQzWoZomMn+G
XyJJNQfGIKbiJxM0o38d/Hq4/yiuy2i7r/6j4MDajv1w3PigdB+Z7oeTkbOaaT1y
hor64L6O6NYrrIm/3NDm3hmZwVeGv+stqLSIpOBGr0LxLM481zDXi1hlRh4BwAgg
rf4KV09fd02oekqFutoAPZL9MXLMTpeBWfhpstZFbh4ng+DtsJhrKzzgrxLgfC1E
UWILz1UXRrpbtwLfsb9ysU/eS0yxeTnHfJ4WkvmmfK5f3dj0niv/BmcLrBUlPTfu
Mq7VffHkMZTmkAVbnLi+Hmwlr72siSX19s6XGKtoGQrVytD0H4D7XkoNO3YZ7WrV
Sl0GYv/tQwY8tDpqLU0Kt458paR67XvQk1t4FWRvix8JAWpmuf9syjO6ia48y5zD
cstgg5W5JXuagCJAziGerY3qm/Bu2cp60MTbZ6NKypqq7o1KQj56U7zYTcJZarFR
cQp5fRQg/8+fuD+IWl5oYBIw/qIlgaZp5ye+oOCkvq5jLCoj4t9ECuEwcMd4sW+c
WciwrofR/qqUkfTC3lQB0cB4bXc+p6a3uQYkd6kkwet1yKbXQXl510ximOcilBRl
v2G42ug+73eOMQ85xH+ZuuoApyA1oOuJSSo4kKielR2K/0tEo3wyrfMVL3NSLjJv
HtBYt2wzhJfF7/X6ayzsEjZXOjYvA/TXS3lnEBA16cXFMIRLWzoXmh1lcQimuZZA
9drWhM0rgXMKPVEHRTT1E+C9Ww1npbB67VFUK9veZjSD+ZCv4NDtvlbUcUL6bIp9
b44Cu8ipsmWPKgCfI7xIrDteE8QTvehtr3u1b5ZZiyJ4UF3TuvvT4fwaHuCQ3FPq
m3/CZuCmhfetv23VtbGJOZ//9PGbAU+6vdhWffL/WSm1rM8csyMEImnuwCACgs+6
k5vqRsylxfF2jU72mqc790SpV1c0w79uBsWPrQenOIYPNl8MugpmFBYAcLAzTrI3
8YE+hHf8H2KXCNtjcNkJEB21AGKPyH3hKO0655WQu18+ad1dXZwBQmDu+Hx61wsu
BHYLxJXiCbkas0tyHwJWOnl+d7Md9m+iJ0404WnmrbYhYHupX9bU+IFZNj0RQQaK
M1BM8tupT3AZQcy7SC2deeFj+uXAqsKxsCY5nzYVj7EpJyxg8ImPX4epoFpAV5X6
4d+PEq136A31wVN83309QdN81xlB2+aMJP9p1h8iA3evBClREg1Be6qcJJ66MhgA
vNDIYB+sHgaUNmZOTFYXLw0EvtkDngAkS7HZFqE75qnuffh+ZjJMM6/JGOATYY5I
LzEbUItHkuzfZ9wNuRO5M/N8nKxk7E4VDdic06yj0ALGF3SQ1IMhhP6eimvKlmuD
bO5zUqbuwA3qf039apRDUwByMQXM1V1oBi8kWvdTKqYgUszIRwjjV1nBW77k+8ZS
dT3TUWxKTJaPZe9MMFcSxSGIfUUyqcYQip11VYLLjwZHlnXWG/5C+4DhQonz6gzA
M+fR22OR5FMtTR30v8viXlI5oYox83SGFcfMSUqJy2P7yzwmtudbvvmSfoVUoteL
VaiI/EzSt2kilGvZ8BFeWV1DS3yLMQMboy4UO3CFfHeY/8mv4phjmEeLcz3283MJ
zZfJf7iQeeJN3V+UCOyjyleFjFl/ybnAB6egWXRxAu/ix7WFIFp82wCX+VY3USEs
PwPXGudF6tRuNS0aXgNpixKHo/AMezQNSzSI3ttQxkGgbBWLjo9rHdw0EOY3iLgw
9qg++RW77Il6UOfhs+h+Cu8j4LMoyeY7eUyaCgULVaJ5wfsg2+XjRy7fMD7rsC50
zI+aYSBHjKxFhZ10gvMnHelQyTIMCyHKJrSI8vC/xwl00lYz/r0auGd4P1wIZLC1
s1eVBsaNEoAOt80LqBmix0FxXRFoeSGJOsymfpNQ1YWoQ5q3FFPmTZCd6EWpBZd1
gxK71HgrUqCeVHWimA2N/SQvKNsq2vZ3ufLfyWGy2UxtKNl4eqCvM04MW3FcfUfw
6gSNl/vEgckSKUpqAM1dElOc0y5AnrZd/qZN29yQigwzAku0waLKC6/KNn9nW7Mo
EzZuV66eEcFXrbDED/a3bUY9PN01pra7N2Rx4kmttEyO2hQVTBiP4wFMFVXWzFIi
VIKhAf1CYxazY7wjReLZK/0IleOwBR5MmQJbN8b6VhylsNGcrQYmmUt8M2cHQM8n
FVAwzqIwlS2rdZBlNOElqPW/KTIrZyG2cdjOmuz6fKvNLWUcEQ+A1l7erldVox7Q
N2cZflLG4soq4Zuz7L6bTwxf93512+jV44zj8/VaexBX+x1ZrBVNFwzguEV44ueb
j1jzZkDIx1m64DtQs0bzvfcV0U6UUNCURCMr04IueTfZ185GL8nEP+YjD+vGQUyQ
8RcV+NDxxmQb+8ji+bJGBpZdp3tGmG85aBgdHaVAAYa6KeaaF2QnUkq7MQocZxuP
eey+oR2NIdgzWzYpRKs3dne/N0gG/xkpjkPfik1Cs9ay0GwRfFihmBOdk9vPahvm
CaMQN1adImCAeNEce6yNzzIz+Nro4e50F+BzGPHPR2Y0es/hyFDqdLlfNuOAZhSk
79Z7yu4zCmfbleEPzTxfhNThtZ0ewDUitk+1oSJVUHGCzGGashgxk0KS6jLGbouk
zmj2jnocWXdTYMYxNT1q6wMGEfbd0flOcb3DgACHNzBwdPT1BsatoyyHJ4v9HBL4
ByGtoTcL1w+9ce+QGr0Si77UsGHfspLSZlGLHcBd2/iz3OMVkg1YsgwfHF+BgaO/
LATAb7dlWhjgHLeTJEPF1gmS4qPTyW4VnD73qs1FWr8D9p+WAB7NVxl36unKysBx
aRAsUx/RaYGllcqp6PEcBdZqkhZoVUvTgRRYEDof1pCP1G3eB2CiDR+bi9j3ZMQa
RDw9LSPJmgDB2c2fVnPhhDwbAGYXggBCDZSPX+xx6/+3fvmzyuSdQS8AIun3pL0m
HcIJJTIrPc+6rflrwwCPnW5eRhC11dMHRE/d0ew5kuyiO0EgxfwQ23JBbRZkTa3b
FNlShblYRmd9voaFS4S9bOIlETOs7FKhmJQhYvk/RTLgsJwrectzY1O/61xVvkKD
FwOJ6LPbEfBoDGbJ365nNCqWMGYHXHzn0XPgjNV/fnR+pIfK5vlINo1OqDGykMnv
h22Ru0f3AafekwBM2vSWZrKmiN9V/O2BMGSZoy2nKRDFHkH5NjUlITyGLuaykWq5
UwX1AFdyHdHKBXlJTvG7oLF4R7cIlzuY4bSeW2NtDnBmkZOn7RlebBAcKFYs3gqf
Y1AvfoVle/B9zQoryIIQS4a6G0PR7khZMLUxBM59uvfBSFHmXvyogfHwKfrQEBcQ
ltB6QUS5xMeq3f+9gXF9oxgftgaola4x5QuT6YFOa2fUbHvf4azCKqB5IrVCQdvL
UJPf5xm+hLgQnBmDr3cmj8AP84HkkepmnJa8TiWFV4UajKjoMc1cJSp9lMo+97mA
7bjKCu5nPYgku97wJTnpAxTnd84BrwuPFMHcDd4TcO0wF9ssLCqoOUDRTZEN7yaw
k04NYSrZLraBYHoJOXlKb7qy6qwfjvSf597c4IGwoJA0vZxq4uDsiiEWR418abGQ
bZZJu8tswYDdznI4j7sqkTtZYc/seZV7NoS+/duFygxXqV24rFvBFLDHgkaSTnhv
WNduCqbHAFQvNlYD9ezrFofylTL1/zuEUvUCls3YyUxFDLQ/JKQnYlLfIrWtxgju
csZTmS+a4eN6G7JMhDIJiP7Bb32VYOLnD4c9lQxZmkHo1/GuCr50XYmP79n3sVGb
p0sw0bRrOGEsBXpIf61vY+DQIUu7lQrdHo0q7hEe6Ru5y62zocwxkNCvt1IB5LJr
vV4NvDIdT86pKEXPuL3YZZyiONrDzVFAdxH0REapjvxNGvTQYAeLnBJI4eGuRr9X
HDWr4PwRRXRKS96VqbOlFjrqKgSiAS/Dq5P5VXDvCGXpqr6Qz67gnlyOHEoVhPdy
MyNcOPzrBq3RgL+qQR+OnHLVOw0kzFtJ/MU5syjuFjnuhWdY2UE524WwFanPMtgl
74vyISQ8f+fC7+6aTbvJ1Y5oiGdHJpNM7pznuWPUS9WWuCpSALhzx/k9tB9dLoML
LuIzSvuij7OoCHEp1HuNjTon25Ab0x0QjVgl93/hnM2V98pJ7Tfz5l3RZYFXsyV6
vt5C0VTfL+qeKfYXIQQkmAkZ9mBtWyqw0rJtR8XrdbjMPMyJPAEgPfYsZ3hoH9aS
nbo13+uwPPcr2YSEetdC2d/DQ5exhZDMxck8SNkrYSb/WKWJGc6+JYKLUv5pxIT1
+9KpMk92xZnyWpJPvJgxkV4otCQVk9n6oMQLPdB4pExaQ1I/hgCL5fedMYTubYSh
H3K14fRzcfvuLojNMdaJvGb+83ltofUGnBzf0slHxvmZ9V6d2BsTkzcF48P/Kk3K
sF0Bn5B7ywUIULNCT1zE1cJR0Y3k5pRKc3j0/uDpmOS62tUkk17xJuxl89vaJ6ks
7as+Eu5ciYeoNuSlihsE599wn8E3cPGNQ97yHfLKezaVg2E5nM+CQW96zpptxHno
ApG/ibDewFqSDv0PdOmOqfVMs5Un8PjOccR9QexORz9lNb+VWguVrvkyrtZMSBBJ
r4mpOTXob97V8cOHeXag7f1r8aVKmKtTyoHh6/uW+VgTJxqNlcf5LXUkS9X6FKG5
cMPOiCMHEUDRDv8iYf1vIBFRosIkCV24rTCQMLu5dTjitGWBOMxuMSxWE/vqwC2t
AelTPa0RyG00PKl5psYiSqZBawyS6/4SRg2aFdu/f/GY2D7/Kpa7KtOYmcT3nmla
UBOx1P2oKMz7acWryiaDCje8CHyrnjdCHsFeDfLo+/fIEyRIomINsBCrr3RIjZ6N
BM+ddNXDMQYq+xuZoy7yj9tF4PcrseE/u+EgfkSHur++/mjrx/UUbak6oINy8nCa
MTqNwIi5o31BSKlxfEJUIXaw6HUwLS2rbhJudHp+1mqtBj56Q1oUkXfQkpnfcJwl
gKbFFcnkX7+B0MggtEXVNZSsNtxb41WADUnBFUCg7qFc8CWW+Tsz04ujdaqRzgd0
L64Z0vu4+EaoTbq6phER0I6vNwKi60NR3GqMjNXbMlwq0fQ/KYggtweT98Cg+IV/
BWrXi+GRtc5JPa+eaUp9oqY3X2RpYkZiAv5XE6z978bmgCAkBVUAgGA7iDxehSHx
4sOTMSlhSi8aoAG10hX+kwZShaEomk+WCUb+2CrwDblvN3Xpt7969a2wMYxUPKMI
DgUOoQ7fjU0JpAAdupMkr+wNwVkYLFH38fT/x7WGJL3xNXU2+huM8X+ZQvOmxrLl
Ctyye9/JWaaEl07St/bZIq9CGOGjGrdSa2ny4klJCMSZMhKvjCwFz4fJ1Je4t6a6
VPBmsgFDCHmsdIE2vLpSIi3A3GnCjIWai+/B4+gpbO0hKgRrFG5GvmSJF4j1WLML
JupX7vFYAJ1grtB7in9DvGnzComGNW6jkN/yVwmW8ORytVkTo8MYd5Zt2Bfs/Xdq
LOWiXBPv849ffJhPBlnBBrtzZCF0CgfsWF7TqbfDa1gDwwbkwowVRgMQeqQj2blw
jdSL2GxKe4ZrRHT8o+qPR/GhGZTZ+LAl28tpMDSWyT4OlTA8tQDDTzpfOeGN16l/
Rdo9BMg2usG3fsJ3s9zYwYebdQIA8W8CNFqiotkU21EtFIiV5bFi0UggUUaxM6Jx
LH5hZTivmmNjGsz15nGNAdGtYT4QxbSR5qhKQYRqC3iMhcp2SO/pQ0HDdYfePXD3
pyzD2bJTaDeD8/pTHVSz3P2lMmoNaGQyzfQWyPSMtxBXtab/D0nhMHRIs+V+pF+C
h8RKNafn+gyc9T/sW8Z6qhX3p7oaV8KBwxIc7nH8jkx7C6G1banBh2tTWs6SUa2j
Rw82OzbM8UmaeZl4YdhKNy7hgNWgO6nzZb9EtHqoE6v9FthQa0BwrJHbAQzGm3If
ZMbAgksV2d5cplM3JKHxZvsdIvgz6d1zZ3QLEVyrkGG1BMVd9ST5yKjTmkY0VNEB
8hMj/jZRPicOmJdgRWDpRDMMs0LB1EFJPSCsdHW3XzK1BLALBn3oPL7/bWMtyeym
uKDUQqgf1Me4cHaymrSmmQKfLGeVOPMER0b86tFOId/W3ice09ioZV2PNlsxHr1g
IWDYeDYRUFoD6+slbxYjgdFoD6L+vwrP1A69YAKGRGM41XlWZ6HCWrEUPnuk3Z8Y
vvwGNr8jHbGexh/9VNMVeqUxB6M7LSOndsev7xOT9aCZmp+KYDjJqDO6L1Czix5O
WjQ2XgFvNdfiIob2dhRSH7Z/7v/D01FJfeuTKb5CffISnTDDQh/ChPFp7mqm7iVb
H/vTD8VFzQhVXdOG6e8oRakrhJ7sSHaQb1k4m5rcTQ59LZOzjAekkVKATZ3yFEqD
zlPhGVwKGWB2V/XOokX1YpYLt1QdYjwpQEvRLSwCa/KKZFVeb0JUW/vx/orPYEXh
9HBOUI2wKw4+fb7uXgxKdeP1l+UUS8JzicgvROM0J0Gu8uxzs0XVRUiSJ+CZK8Nv
fd10wvllgCb4X+RBAXs7pYdmHcCJvDhSnyR7pzG/wXDXffo5NOnlKh2Y3pces/ow
BJwGK3crI7VP/rql8MWWxbaoqb7RAN4C8KTxtig1dWlcBbZiEIyQCWYGW3a+pQp0
TWNi5xt/wqtVn3M1VfIpro63eXgWzwowUImp/1H2HN59eqrYH08+3ioZ9nGPHJbI
Sff63I8A/VplPooKXOWZzLaTl6mm1Znxy+7CcDqO8RieVWarw56Gk6zRqM+vhYo/
/t+jIqdrKoWgEK9Vp1z7NNooOg7J8w9q8o/HcPlIC2rVsKeIpf+AgNbd8mz3h6Bw
VSlqlxWHLZ0DH3XZOKieFkK1/lhoK/VtnwPZvrQL4hMngo2hyNRVGS8MixMfKOy7
/z8Rm5J9KuPsQiJjfXmZNYFc0pV43KEsxAzd7DzliykmXGddvQDfbsBdknl8Lk7C
1hWfJq7CYFnum8AGp/369O1wAV1ATP0lDLl6vlZ0kB7sBR6cJPlE06xvpKxjxkas
o+Cp/BdBfaC16NP+qVP3rR3A3uWd/zA5hF81Fb38XRCLbhE7iEaraJyN29Wq3xoM
bxIAXxohymKNgpcY2GBsV40NB/nCSXACtl8XOCLZPBAjmgcsRJrjJVXZ1lsIpZvt
S7dGHTvEfOhxxADmpWbV3tBOr52uUfIvoS3684UxLCxKIKhcGjBs6dJDQ2qoxAhU
6RRMVSE9h6AI9HNTCi7v2ILk36K0hihOOkQ+tql/XSOxWmu/s/GFMHVSxytZ33dF
K4/fICEkAhd3xqREPLB6gSP2aQGP38alBNtTPjwbhPwj1XiDa2pfo5W6uaP7vjsS
hRzKaE5TSzOSHNSMz7iek67u+MJc6KByJnL3KJNM4AKZNe8RqFwOLncXJFcSzDc7
w4e1kit2qVmaK2eFSLCuFAgaRG9vJcjH30aQq7VyImTG2seUIGeCOYjGKk+qxt8P
PKhEk3UdndUQ9OGOrXkv9VZQNPqTNScurdUoB3vObaoIUo92a1PlJCxmL+AE/V3S
1mbZAiesIch11iAPTWUmY+UkhEYqZHbs6rnjacfMkK2h26V/kOvPzxmDf0hw3bH0
6RnFI2sseGduRA4rtW3yOiNBPLky2HYI7kJy3DO/xBxie3uKEDdCxyvSX3CcYGb5
j3mkgdUslWJHYrqMvDMCzdkKsv3kgSoZ7m/nqmgEwUxEm7BDRDwJ7C2rjDA0CCAs
5cmZpUfkzD9ksplH0eQtyk2N6lYSkPOqdJV52S4gb22V3QsJdAQO8q1V9dw2w42e
69ASEMLgbQVz2ZPDP3ygJGIgDowiWZK3e/kLQ6EG9jY6uj0/z1Q6eSz21CyeMYed
DtWzEKKwWLaUibgk0mNv0zWBqKUJyiL2H+7/QT/EBnHHfGS8DJTP+dYhj+vd0Y3v
C9Hs4gE0dj/2zEY2bzDZm20mhiEpr1RPKS/eaUPKml1jT7CwRwLVIR+bkEUS0heG
K2ih2K8uo9PSycZ7EC/jLlQ9vvLUJWjXGcXs/uaMVH82yL7mmHPmz2dQ2nIkgYuA
FUuq43w/RprOwm3eN0sHE1qsgSlcwIxlmplSPCDeryk=
`protect END_PROTECTED
