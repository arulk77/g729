`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN3uYYQY0IXDfyJlGlQUFJ08FPR+tsbEf75uq0BVqz/B
bCQTqCd2T+fkqzm/1LvEAEwGHHyCDJ3LrO8Iv2ZQ7G8a3Vi3QJXTLQTFyFVv4/1n
bg6IMOnMWVfNhmneCxPEqCK7UNVMIzTX95fGeAK1O/3e6XtYq07O6Fe0jyHJWkPa
bCw5v5ijj9z5wZbOCkH1kcsxjLS3bj8QUzVo+fddhqYXCruPt1fZVTTBn1cogAxL
P9c2hFv7s5t7h7vIpic31Wvtip0+h7S32KtplYqTwLAyn91OX4B2uIUkZ9XUF1a7
Pn9H6B3GiJlTTkzNek+RuC3cCZxH5J8iu+yQRbqLoyNYTpTRKgP2hwqfZ1Z2bs4z
BaY6NsRa3hVIFGxnJ/nvJh0h/x07oFT7NKaovjnxpe0ES4oiV6FN28/lvFdSbke7
2oq32w/OfRCM6PzYa7HIuWUMNdKcZ8MM1uvsLUHwLY38TMBw3JI2YXlFWZo4OXE0
VEYGE44+v0/MNjgMab9hN5Q2TnkDUIFQiWt0dY4PjPGZo4jxGpfph54cOgxwVRqL
kkbos7IDfYxz0rcczFaM7684DB3BPlwGxrUNIAE+AY0=
`protect END_PROTECTED
