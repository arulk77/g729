`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAvx2Yll7zKWJJcLW8aqrvK99ffU/CcNTW8bwIJC6thr
uhn4nCoGQDc3qii6lXU5GMm54m3shabPE9cWA10RV/FBfWzdfzdawvnPSqr9ihvz
gsDqS6fhFZ2/1g5MtJTYzLEfREzEGgXU7H0dxzJo9i2XXLM8bfqrW8VmYcsmAE7k
cGeyG4c7lbTWCVOz28sxVM3dXtjDLn0NMW98lDldf03z7efsiwApuHWCvoRtnvQr
sA4FFtUd3fLdJ9rl3jO5yA==
`protect END_PROTECTED
