`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
NCgXTppOC4uut3/fUHet3uxyGIi34ffkplFG+lhg76SxME9ocNR/wRChsvFna7GO
f1XzBGSzTu7rupBn9/tN9cf7zerX1CNH3w6bEgnM63SC6wr9CG0u/Z+Ij80RhM3O
L2wdr6M4XycPNHseaIrYUipQ7wkM//UyJZK5NaPU9M0OaVeujEgdxUmlqi9Pbf3a
kef3NGQw2S7dkaarU8He85Cw/oXjD75BfWiBmuXnZzvTNC01hJL1XpDUF6XL3Rhj
K4Ih7qb0cHtkjlcGaEnUtfYZ0x8ELlRMwrYR3aXnWSg8+3zW7N8AmBko4n1/agdp
Ej1GugXD1X/CJOB5B0pHlsIA5/ztZdX1PgjZ0/3dZMMr89aeRqrnu5yP1E4rWsTH
EtwlPgmFtNyFJZPwQPHNEh0mIp+OmjW65XZIbwnBGR4=
`protect END_PROTECTED
