`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mlFBzCyNIVABC0bhYTMiK/VBmX3KaxOYYxCYQkamYMqKvnC3a7zEGsmnSQGnjic5
BD2gQQORilsmjy98YJRb8uFdgnkvsv/uCn35KbmNBjESBLoP9NlB+HYcXkk0cP56
Y68GOrAn5Vb+mN/acy74gw==
`protect END_PROTECTED
