`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEVeC0576x3GhQ3qd/iDhqEyD33tUrmWT70mHAKvMUxH
TuAt54naBqY3Sitw+Eo/DNQrt+VR9c0i5eMzt2HCr2yOoWbL2HueqguoQlgCyYBs
u9Tg4VCa1UqFO0Xd/egzUx8o8Z/ZmhERLanrhLKHUsOSuhTUKl0nZKGFcXww2Oof
vpSZRzOdpzeKn3eYNubltg==
`protect END_PROTECTED
