`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49LDGAYQBGYSNuUS+LHAM16f2cuKqMv/McV/5vFUpiU3
VI71ogkdVYPu/DPz3vEw0GYcocroBBj+3CxU/+LmqYUQ8nzBp27dSqc5LYt5UInY
kPlKHtqX9EF20EE42k7T6F6BVvJdqMO/OL+0GsELK07nOqQgmA3nybLhclJMUzHj
NqFTIYS+8mR6c8rNZqdnVSwlRHHlEkRYoM2UTFvH0qBIOM4azKRCExE3UOZgD+ye
ZFo7U0XYr4zjTh/9VqSlXSw029rkQ6pUwTEjlfU3JTQ=
`protect END_PROTECTED
