`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP9C+oB1sevNQHRzpKe63tTDcdUCq++Pp5srPLgkkibO
xKYCvTtfLKPRG5gmNv0Ap+piBCG7z5jK+/xPuOljJQcQgIDc/CnNZ9NdYLF8wBsa
ijwi6UQ++9CsZ+n0Y8zdjbnJsvec2XHxZkj9GN8tQhuMANOGA22kujjSIqYANWlh
qFYG3LTMqMcw54M3huez3+OwoicIai8FIt8Gpofc7BQqMfLxDsgucoVzo/Es1wl8
UoyrHi6IQVxNELsbI2N9l/tC/8hctUiRz2zuA/IIuXFYEB4ImO1bddwSMAxkz23+
/QF6B7ppju5OXcpgX05ODDiKQejmgtxdzWvwlCmxpD7L7omn3Y92Wqeh5uinCnr2
+flMz5T/ECD6cT7+WUzuh8IspzEeTybe9Z5exw/8mJjwhTbyXH4QX4xmEn+nQGxu
NS7PP6ilN98fNi1XycW7pGhUmc75SUMVMVvyKnatSKiUCmZHLkuWgS51f8nSfYCB
G9gkMsvIvRi527oyikyHH5moY1+BzIisWdo8Gp5c2VRfwCPextVp1K7tO33dxCaj
vYZzHzYBByWl1dxRErkvLFdU9IiNNmXPFxBDTHTurIlFglY86H1W2VsbWt5akXmW
QelOLstUetSPKX2YXye+GPWDJ/WrIlOqDsa4FjHcLuRsAl9sas2T5gVGuAPWwZTP
4sWJoByX0Gn4SJvYDehurcLIeFLaeQDyzPKzGJngiPnLrboffAz7N+BImxoqoO/u
mbHtCqoYy/T1qoObhsU9FrHDLazsRgsJukK3r0dozuNyS6L9kQ6q8pcwZSxYyFxN
6blBwL9KBYCHFL3EIG0HYj0CcihJM78KhlvZTkTFcKtgP3v3dpTftBoFf4hUTat2
BwfEWxzIX1q+wZDr9t+RWlIaF4USefDRNQ/+xRU3l6PCpvo+b3/a7Fa6SX30DJ00
38NAeREd+XiKfgl7mx9oSz6PKQ/7yxSKwsdTOyHmOZ0Cz6NCwq7u36/NaKydCrNB
Wti8ZfAW9D4N87Dq4EBiCSlcqGe7iR9oCrDAR77v/3patuEXoNykj+qhY0VMPyP4
Sg1uwWRdQmiqn4gVCBH+l5MeDKg2o6ty+y0M4Jhyr3K92vk6cvS2JKHurvirXCw/
xip+9bmrVFDunNSIjZXZXO6qjJ2l2CTE3a8SHQEEVEqvX6U2StjNEDK/a/5g9Gel
hrMilEd1k97eMyaIAqGNab4ZIdC/ptvqRK33/Pkgis+ZqRAUbPLbj+eY6z/KflAz
1FpUs979jQfWd7Sik2L0ngAP3j7YNreNJZmsvZk294u6Wg25fRRzTSx3KkkPhUzB
XslAUeq00PrZLSMy9PvhWZo7H0IUEfrZ994MqSdHnQTS0XseBOBw7Rjbs61Kewdd
5L2bv8Yr7kYWVh+/KOEUw61ynoIvJG9QSBykkgpN7gMQpzebJsAhnoBpvgcUw1jW
AQtR28DMDaxdfq+10wk1GR9c5ZV8XS+8PIeQOlrq+pNj6jsJPHwyethm+Rx2UhNW
+C1okQ5XU3AbqYU4d07KUIslDr/PDZazJTFlO8KFFC/L7GdsMjQ+hhDDLNA5CKbo
Kd6bRhseEAMelLJzEME0PKCPTcxMATZQYRJXPwQ83+kqvb03S/yoF5/OtQanSIzs
BuzumFX8E+XmAxcxfnMAyQyrK2I57Em+DjKWlVpMY1uA29frKWBpnvZ9CMhJ4/yM
KBgQrclfBI3XSUHocfTVU9BRo825QUnQs6MfsnnmU2LK0QAoyEmmGMHaHYc9xsch
74DOz1Ol90gMRYI+zWQMkqpKU9a+TtK/v8XxMV2m4+cRudEXX8vx6yAhiTGwF6b9
ZdgUdCTdHCzNDqaX/fgz1zwShaa5h3D7WAyrV9pFCGBwN0M6Ikasp9OLIOf0s65E
sHYqqrucRutZEeQpKGxTJkaLkuskYe1MOeH/22jkVDbOnHprIcRif9El8vfE2An4
MQQKfLBWxZp9fr78V2n+a2WowiPsBjb3eY1BDqsp0nfxEo+GpuqjicV17+Iz4A9u
lu2jVcgKrrrCUlIu4LRjcuZY8FR0Kr/vKmM79ESu9AUntGbKCVstpb9TomVO06+P
mRnonH5l8F4ADUcwlXaolJVTh3z5G7heEBbbVoNo4gTLZ95MET1/Xo542E81nNMW
Ecmx/IfQwjQfeO7yb0asIWHqu5PAyb1Ga4eXxsCPlVLcePM5BMF6hTxp/IzlIHc/
WFtsygK/L1r9GGkLv46122q1sSzwAN9TRFWw5NqJQaHgnyNfrXoUvsSsN1tO0CLe
dNNSRoeMq3bcUreiAUHpVqhxBpwNBRdM+8onBpM49SqCwgPjfpTYsBulcUm1YOou
2UAaQIqPDeTmR+vekWyhRwLxA1MACiBXbPJ/V0yiuqasWwaMhP486MX6EFi4b4FU
drrdC9WplnzCWqnsGu8AFqvioyAhau0rqcbxZTpUg2UaL/b0DupjijCM3qKIm80K
88QFTId3Td0l/py4ogz81U88GIlDwJ5reUTsXH5yrDTdAKk/UrXeXTD3rEQ89a6h
F4vL9sll37jDPuGZtGqjtJszpOPDBsMK2hYEP5mi5mkzBCiRkdr/VuG7Hmp31YNB
RO+LD14HOu4QkyJ6n3Lg4ke7uiZdrEjv7e60IDFXiSv4doImsepjZ2KehPEQWZvM
gn8pbASbBlhiT+4EeaLT3tr7gMEgsvkNF4Sd4pNQME0=
`protect END_PROTECTED
