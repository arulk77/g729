`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aYJAuNIpVSdXWgZeluU6vX2QIIsSoEgw/3pKiDha7kAS
aUyX2UlPOY2zFLmcuXRZ1XITQEFhKsiD4KxHBei1s6G0IYLKARCQnwq0g+6uPLun
owcBGs6PT3KL03El6+LtmK/bAe6/v9lK0qH++WgMZx2idYRhdyjQQCaDE3muKX5X
7X7se7yyiTig2iBTLTjwAyGGOWjSCmn83VeaEV4gv+zbEtIfsixMFzECgkflNiTt
Im+s+OMcbVDSqeH0h1SP9rcZuVhzp/uBn7uhcpzvm9hFORFJMAx1R1o8nNrS+LxP
+91E+cD161xShJXDcdUutQv+W55s1hhJ2U+k8r01ZZKY1TLczJFowLBhYojqRCN1
qCQseBs/dHFh4scPIZpWm4SmgZxw48sE1synnrYad8c5SopiZV+dZo/yfuOia3lR
AgOL7Ekx/oxnewT8jI9s7MwD8waQsRJMrevfXqSxU3mp+EvUmjY4lbfOHPvNC4Ic
ASL+08qk6eRiWhSN7gY3IVgusuPRDgw3UyHX9xQ3JrEeU1Iw4zTPN96Hh1y1Kvd2
cr80FTuGEDo9bxsgxxkEwgfGuDXzcEmSAm+jqaLQtMC64Z/hD7qD1VKRG0cLIPwT
MfWMT3DlqwgH3CkYGaTxn26AGIX4LGnkV3eEemyngvuGeUvZPFbhk/XgmIlHV/Mj
7sGaltaXwINSfBEllB2cZkA0VV0eAbjgdO/Py0SrMIPzYfL4QngF+TckykMl5jqd
XBt8hunDMFS7JpM2m7MCTY55S3ve4FfumBOxBKOcMVXYYCMNDnwYT3alo+FdjnfU
`protect END_PROTECTED
