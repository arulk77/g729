`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yGlDbUMtvO+2oYUU+7T08HE/qYaxRVV56riG8Q52lB5
v4EEM/pLskyzCyXp49KiXUMTQCSooQDaQKrrra14auNVLc5cn5OZLpUYU97MZPwa
+Kp4/qPxwZ8MS2WEcNsPaTt6ka7O+x/MAUkMFR3ntt4dRz147b4+0fiAC17cRqF8
jwWeGo5Uy+0kDPuHrkll5fdKu4LigrHFG34wSb0DK9lITG60qUIJVtVnBUTx5d+v
429NmKQ76I98oV3CSQsB6VDe3e6O2qkV88Y4CSNpWq4UrUVBIHfuQoXHFloxeQFv
VVtDR94H10bP/tAfICGOhvv/n3n1dIBnmomqZIYuu95puZmsR9qRZ1uI8A6j4vbA
hIh+M1DYgQSNqdbTwCEEmw==
`protect END_PROTECTED
