`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47IFLHgd4N50HRrTab5z/3EIYqrFw1rYDqxPUJUli/VW
0CZ1vIZ7gUZHSHuYekXmR7zGlw9AqLYQI83ropCvUNNs6nZWBg5ByU/J4c+NVJOd
ecMSQs+U+zMscp/VVlyQyWf/plGLZwTlPyvLyp5470fTeD0kBY97ZXwUu3CgtXCb
QlqbDJrH4QjxuokfvGd4Yv5TP21BFGTuDckxpIbA4s9e0gxlP4vYkTV71tD2rvLr
vA3YUcNrLk3fzM4NjAWkegIqJqEWbhQo6RFmpLd6Qytviy/vxaIRgKO2lEn6PGmf
jAUFwswsh/IzT6MjMHvq4hKG13n9WMGilod9bsxwyHoGp/W8gqhf3WTdQx4vsEu/
ms+l1xA8PVrd7l6TUUkIxw==
`protect END_PROTECTED
