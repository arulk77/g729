`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
1LG43y7n6eeeBE+He69cfACTK8sHuj24fDCo0YJQYL8ime7PtOZW9zVK+naOkQJZ
/hOjQKjoXavOJsFCerFSHMroOBsd6X0yYZjLdZIzsKyl0waq59qR5Y7jGGsFky/q
vggoKUSJTwZ2JvuN9Uy04CALzWmjqYh4uN8qgC2CjGDMcAuEKoHrBL6t0GPxQ57y
FSx6Q0LBdVWQxdFVuThRkiALU/kUWfuDIKIByyDyh9xMJjBLSP3Up/EkuXQ7oSTw
XBuFMJKgGR1C3iZPfUBnvGQ4GTsdLz0tnPCFM7+m91CLWMio6aNB26qFAEre+m4p
ch0wcN14bz745d3WJjCQqSf48W88P3tomgknSyCXjQ0pSx8QgCRj8CHdnKUlXai9
n4qnaibzbeRTy7pmmrrligv0+SE6Pxnj+YGOjeH6OXHFWGK0A+xs3S0dOpxtykc4
wFd7vf3nMhe3aeG+euZPAh7htO9yDb5Z4kzm6DyvX6b4tRS6FPPuP7YTq7aI6edn
VM8j8+3SO8Pdc23cQluKZd4bv3jlZdtOIi4YerhQQRQqr1aiBTWmsmQIaTH6OK1/
QbnqIRVVfPDBFjOV3eD6bWLwpEGukzjrXp/j1+bOpj/lyVicFRGuSZ4HOlzwa+Pz
yZpWRyMFCHV3zn5alkHHnzRfxoFdQMaILX/m9AhcQKfYDu1zXPaV/DoYBOr32688
`protect END_PROTECTED
