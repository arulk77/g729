`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
6O+XrkSpxtumpknl80QG6wh4yz/aJ905/Yj++XA2scqP0s2OzYBQaqMjqnDppv/1
nRMFvGrTAhOAtHuMHEnP6J295Bo6jCXIci/8hIaS3SbTTg5XY29gL9pzTgXWLCdl
IhydyMd2p6EzD/Uv3vFsibKA5g906IHFCpcriBR42i0BIA64fvF+nqDAvnRHDdjx
5YFymmrUXZz4fqQtCZlIF4qiGtQXff6kKgPyhEStXdiYy4eCt6FkFeQrKSuJ/2O3
A8uqUaXaNo+6vHQacEd6tkwCKSLFhLTD9HUsdTgdYP16+zsywz8BdRQM4q/rld59
lH2XyFFRpvWE7ie3prfNtHV6WjJir0b3RaOEe1hkqoNcHd+zHQyzNYTJYuXMwgru
ckJzS6IWuKzRI4O3ouN21lBimvZyoO+8NH6LbP0C8sfvrxp0Xu8IivvzIsfu3sEm
/ZAq4NPfxaDMGFr4rMzNLgosbqHQZ8oTff4S/xHGWOVpHxym/85/RLjqQ1KfmNkC
rzfg0/CpKF8cdiF7Z8b2xTICIO0dEN6BhE9dpPOPyyiZu6+sRGeB8WV55MsJDqN/
KenNaO9Z+ad23lUk1gqPX+9+4VACajb7Z7hi+RqPk+672wJxBswx+y/ezfWlXFww
MPE7r2E7fWl9AzoyptQ9vgOyW/5I/65ChINbF1+NxKIAskudZ768j+fWr3Zt72Rp
i7navM28bWDExYRgW1ISMrkcMXOkqqp3yj6oVhVJXu/5BdJ0ZH+vsUV2kEM9QdHn
WZV60R+mHspDs35DSqXWo25aGEdvGFTKf302IXChDNOG2Hwvuahi4ho5O4QkGBoJ
`protect END_PROTECTED
