`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
36A/U5tO69wVl401zVMLLYErjFRxSnsMCvWcjXU4pj5QiFPJhw+WWzWKjBmgL32/
0y3rRSemqEFq8/xqSK24kMMSHlj/3swWInPlsSBRt3aPqCXr+hiT1rwUAF8inkSQ
gdbHc3z9ibK/sY8I6GeOl4yXx6/c1H/oQTcKkb6VTqg2Nogl5xTprLtGYw/JJWwc
53OWEhkSB/0I4srJgjRWa6IMwV2kjFt9IrGo0tQhaO4LWGXDoqfjG7w5qVDmQRoo
iKfHVeDySnrAXanYDYmGysIguDx80hgBKuOhZTc1/mACpSGaeIXoKpYD6W1/Whrs
NxOBgfzbPKjNwRCQnsEKdQu5HIBT+tRwWLkkKGzI8jk=
`protect END_PROTECTED
