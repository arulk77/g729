`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
f11uP3tAS38J+2XEq2c6cNQoqsmRKFBiCH72SFRfve/AnMxfU+7CFQnpMi/afZnM
hQ/XiooWVQO+KLY3/A8x6guXnDVtPuwNn7R6UOgq8wvvGZYzlHzW7xxYslm7GAdg
8B2foNbABgrPQO91mjqE/speJoyuDJAFJSEUjyJWg7dw1A1FAbQYnhS3WmeTCMXz
`protect END_PROTECTED
