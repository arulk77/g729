`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aWF7FwcaUTFtJVQbjpcpSNui3tUdsKg+x3sYNoDLem6a
sIIxtZp/UUPdTa5c2g9TCJjiBzOafsAFPmptngsLsqu5Li8NBawPPBf2cpNAvLaZ
a4MnRLFpZgzdpRKGnxkMOv4I36LJCJSNJiDU/4geNfywT0CjKN+9pktsZJrUttzZ
8C2cT7BZNuJH5PqcEX80FAuO8C2AIPLskTvpQ1+2s44RH+0nh/lPzJfqsM8boXsF
t21Fx4D8uBwaBYyVo9lNZlQX+gTmJeb2HNzpMyLzLUJX+fubVvk3moOu5kDKplbf
XQ7F94QQFjhov1nBo4zl3APgk7AFvV9mb4/J9FQA2a88CJo7MDsS6wL/8GIiwTTf
8DQCXPN9nUEQgLSvnV0rXaFGWuvum1RLbfN+HTFBj2A2T1ddVfv+pDSl5L15qU5x
Swghs64mBXrPqcCSVQh8rl6rjZ5PV7e/UDmRAsuvAX4nZIlL60Dkpe1aZBHt5dZ0
KV21gxeb76TGdcg02XjuOQmQoDjd7iLB2kTmdefcxWao1GmQgOkzj/F93DgLBLn5
0em5g5eceHtw+ZIYean9XmdwWJ7NuSVt4KQXYD89S3iXCo3eeESJCPNrvo0xeR/b
COFSzPmg43eXU6lsHeFPtGgyTSErF1e4eggpU2PpQkL/FpqvsZoLg5bzaNEEbYLa
fpaurQ9fFMNeVbPrV9tZ1bbgPRVPasQGqb622j2oKsdVkEtJpFnTe2opZeTrgprx
jtIaOeD0Uyt11KYRLveJokWCCqqAPt7s0bMo2GMKu+OWUpcq1EvqScVV0tAtdPLo
rdc8f7N/GS65hERPyeujCevEy1cLntKH135uAPn4Z8Y8WJkZcf1yKITqRpRPnXrt
D8KHYGoLE3qmPg3Yy+nqCp8GIZmgy3e4kkLMCjbGJWPKoftKmMUWsdOVM2Dhp7Ku
8GyHP+dKOI7toQibAlTzGLo/A+8uYeAteDUAdWd1QdyS6FSoezQY8thffUu/8cs5
ObTfqbHW+HOfrWacx0mLkv7MWCsb4K2irsmUA7c/APzyeo1x+EOP5oRDGVGrdzlr
QDWDpDIlFesG31ca+WgeQ/PWsvNnUC272AdScwjC8+2BPFVF6TenSwR1DWORZUDD
N9Sr6DcK4Kum7niY5fFpzb+0sgceLSNcbJpkh72z8gDvdUvMn0b5bFXzzFNteVQO
FZBCBZ5kCpFVTaE4AJFxA+NE2bZExHmJAux31F55R6hySXXni4fYN1fQNJWsYBV9
+n5G7c3kjHld0klS6IcsSGaUC6CawuvhNWfxrDprecea4Ff9k6y0iqXY2jX2OuTo
2o9xdnXJRcW7Yy6S9bKc1mUr7SB6jQ8NSHoD6GGB41ABWamZ8wbKquKFkEOvWsqz
4msyHJ86XtChTkfzmV7t0MlTYEFtCQntMaouda4lLSv5Q8Z5B443M7/B+jzf2z1j
PYSlFinFlHK4MCjS8snmKPBUeODtgmb1enaPmJyikl/kbBg46R+GnFNvsh0Q5FOt
DHQU7EyoFg/NVeiT4PGQ5WWRoJ4ifmdEMei9s4dpfOljt0oHQhtE3taqrVQfuzNd
U6/zWAotv6dXGgOsHMFu25MU0Oq3yplyopmcZMcyTv9xGEpVFe//nfVrtycUUy4C
qbaGqFpqvovr65XvBBt0Qt7vBpF/dhKPnq5FrSd+QSecUKFU3m7IochxttHbgLmW
99Vda0dKhEKihCrTd5NPcr1kfShkNmyYoS7nnm9ejwxOX/uwBfVAmbhdILGM2s16
QVBOlGMKN/ec3UheSa4YmhTM0uCDbXYkwwPJ0OAc0aHWIbMLSNJ1GmmFHMA8kWXU
OIvcHghVT+vStKuU3PgjIBSsAPyDkdlF6LMgYZlYfFtN0qCXSeOv1dQfLcS+5Ozn
Q0+lephAbCWNxv/dfJFeZBrXP4oFeDTomI9eBvHaWBwJt/UBOHepYbcektfAYt5Q
I+Ikj+FTF4/mTRDbmU3MOdlJw6KyZ1dam8ybpocRaciN7hvlLCeLc0owLoabHJxM
XkzZUr5Ui4HXXgf4M0VISAKpqcQcU7ViO45MJuYCPSJfI4cnTp62qAB854kFcjbw
hklPRxg7b+Ly1I81IsCmrPkPbrVZGd91fVcimcI+nON0OTz+0Z2ytZbgI8FyTCT+
zg/22BbNppS4AXqcWvjYKCzz3jTP0vrRJmbuR/5cxzkiJW10Q8WgEsdnINq/PSZE
KgiR0TJyYVOaaiT3n37Xw6ewp0/NRNo6isEv1LPDV/yHzetEJyemxyMG+XSgWFYp
BWL4cdYujM1Mj51Li2oRGNQ8Niq6twZYr1bhG5Wc77REu+e8vk6DJVYJeYnw0FXH
sBL1fA3z72Iqm32gkfBpULmeuCLfsqyh0Mo7Yn4wOtuCxM/sOChGHYDA0RvtxKh9
pEB2LKeA8w515TqxlHqxV4BVt753PWUsFSGld+7zJDIrCd7vP04eF4/Bk1Sf0p58
pJE6TC9N68fA9bkHGeJvC6hY6EPyewJrgf7M+2flXfqIZ3NwR/wrSDLVLuYncLrV
ObKJwCd4Znd9ZIYPc/WgNrSD6S7nNrneL4qrOhoZ/xzvhoS7FKmvR5s5u705EzSw
4gfyfXDmLP6ZYxo3vzGGiI3nhLxJ2i9tLuwBfUFX2gbrnbXnS+DzwWwbqGIwkF0D
gnC7YqJgW208gz2fMANCtDtykT0gYcDMiIRdv4DbC8wXGSzewq8Rl9nP3hOF6CyB
HWVSMWKUhhDQOcq23J8lH7oBcwLS7mVnfpidLlHEXjRtO6xuQKOz8iu6ZDqqpKNX
JUDn5G9uTs+OD+zNrTyEnc1apHz6VsUQ7wq6M8nAr7Jp4Y+LtUF1WHYs/qSc9xiB
PAh3BUpCLpV3dP6pHVbcPTt07o6+ZyOlkfIfwYTNBBJK4BxEOhqtJnDV4HM3oIl3
p2sYgjxR/UJ53infyyXaeaZLR+q3gs1cOClHz+8LVYvvAmxVtOtasFvAhVVZ2gx3
AhrJlxXPamRgdDUIovgVeMTOUjVhNHyRhdzFkXSERblNT7XkW/Y09TLcTmXlonLu
Ii0jmfFAVieCXRS90F6LRvXGKR6S3OyU7gxJL5iCGFoDuUsmsob8UzV8pA1j1oAQ
aTg31guNPC7vHB1/4tKQH/pqNpWsAv+uP+sOrhVUPZGpcumXKlqYtTB0Ix+n7N4V
xpKuNk47oeiqHMuqRr4sibCDj0QqawVZPSf1yPs0dlwlpTO17wU0Ab/bLyKcQZpk
ub5d87yVE3L4HugfCQ6fmN5AD/fTzpNP6JM9SKJMsaSRb5FvXwppuh4y6GCbAAhb
aAJGHn2XqyaCUGaWUBjkZfaGTowj3Q8b+unY3wBjQbpKZKF8M9ZZRHFj4oc/8ZbU
rQl4D7fj0ngByA/7m/MU5L5eurin3MlgOUNvd+5LZAT9eLeax2K4xcL5Ll3juhAD
mRUT80exNqJ2CrFh0k/cB6zXmxbPcsIoqoUcjk239vWF4HAHQkVgmAQ4ST4NFkCj
gDZEYIbundVzg5Hn5KZPkfAzBHuGVe3QiClEAaDXmjFELn6qc5na1pbTCATzSnKI
eLvG2eak+i0BPxuGNlptXgc0kX4TcgZzh9YFIDtvC1oWljqC19dsaV2W/XgDJwP0
1Cvg+fVb5OaEwK2Exa3qaySb2D8K8IwND1XgIyVkusST/6JixRB5HlZf4z9EXTN3
EAuGAIGgO9vCL8FshXJJ48qknu2l1WW4g9IvAsBEjgXuqfpC4B8Zx20WKIXbQ3+I
4Qu8Y8tCizXVwvgz8OAQfs6wuqziVSKGzqvud3RO2KAG5t2iRbLl9/o0ZYy7uvmi
hCU3w6BxqbcE06+7V/yn+dfoP9p9pcm50VsPSAhQJsDKWk9EWUKLOTvrmJJPlsvj
SIVJS0TgTis03H2XyLIbg0XPTmTspezpdujjoBkjKyHELOnhAOi+5Spzbhfau5sU
WgS1jkn6aenUCJoBxpwEtEZWbjijdthXj0Ub1mJYzJBUP17fbhVoeO9nPF1f5zIX
35+kEhKyEdMrNA+sIqEVDkwiNG8N43cYUqSUQjH8kXgfeH142KN8ZigXovhT39ZS
Y6klEgpjUPLjVV05AEVj2IcuRjTNQ+m8EIEa0hqieGM/8y7CPeBkyria7u2HsSgr
zYBELZVpQEfUQSR2cmkaC03urGzxj09dUxLdq0HeFdrTHk73Xo4DvtUlDRqcYMQn
P8QNH9BbicxKykOc9Ra/b/YIm1ZaSQ7BmiI9gFNcVVpjTX4VeSfL6iAg2+an11AY
xwPieXi+1lhF7WIGExZ+PZMkG8DZo7beXyIk/dKw3NkTWda8nIC0mfxQ7s3GVY+n
cjRw0NY/bFWKrdxKBJ+gMfdKrzuVKgAStxbfkOP/R9gZEcwglgB/oAzGtFbwEJIZ
dhglkau3/WUpbpyz8p2O8IVuRk8px/+nHSHRCZCX0GyL55e6cLpTKLr7xidBLvNw
MPqWQf0WRW2zhOvK8wkN4De8ku8xVagocqzW+NukZpOkBi+J2hSubiNfEL5IGhur
TU/F04ChNcOrMU46KHT6rgaGK8BufFj+kcH82nzwfYRPLvIelfX/Ci2if1k17UgZ
zCy8WzIMhus5W3fijL9CwAS+mh7uKeqJ4rbXVXzl+i/B2GPJtmycj2EklLnNuJsj
Pp2YRR9TqPt/1X2NTQLT0aLaBF/LSMZzBEM6Hm9qhQX6uyqF4GYga0Ph+stzwmhT
tnE+sXbl2mKKesZ8rCZb8x7rkTxONPMgricUr8E8xYbGSBP4lkVwG0WUdjkRo3uF
KJSN5mI8lunRxIhi2qJ9v4ZF/91qGg+xn1bVfShgEJUIwyilF+bg82VfQTq4qcQr
wO026U8hY/xX2bmpIDnagK8vEJzgnNnCUY66ps5SiKtgfIZYiva3MExRU523Z7vg
/y8ED+QFQN+FqhALfOynynbvGDIj36b82V5fDzfcVbOCnLfL/ESU9nGadO8XYaPq
rh59gyRfw8j/CmxVq9fti5rOi5QOYuX/JLh+s1EwFM03JlHe+RdKAAYWdUtsv5Og
YLOvLtk/9IZ1MjqQpon7cd8glmdngCFP6nINg5JXuXDwv8HtLnd3xp4Nhqlv9Ig+
dciiky+SQNTM8eW9eeWOJ85N9Ncr+qY23I4s0aVoeEqA28JY0Flu7oLz5drksyWY
xkkCnM2dnJtfH21TqloRXyoBxA1agiTy5Brh5eScoztKMlHiBlFzRNCGa1HuGaFH
UA+HufQUACffAd1xURgi8Z/2MVUzzn5IiRFy2xUpx+pD+SifMVCEuGTb04aEb/ba
WaNDu7CqosUoSHxg3XkwAR9n8DgQk+9Qd3xFf/zaLsIj1KtwmIKe5qdybu2zGnz3
uHYxM61Ofdxnxr9i5ON1jOff2MliU6tBtvA+z/tDICNacT9DALXFb8U2rxjJe8NI
gmCQjjt5B9GA/ldOJ3eYjhuWxgKLe7BPCxI1SFBLOX1qvJqj1dg2IlaKPvvrO8OJ
/Gy3GW5soEJCojqLEBeAGfdA1IS7CI2F+jBYig5gZJh9aoSeSW1vWeefsMB5jiz5
VHrXGEHpX3c6vXaTZEpMtGSAyaK5Oachtr0ueRODMU5+PN0/X84bG/3E5JFsW+if
KDfBjfrGUN28ZDcEtzGjMh5KNttTZGN5cg+iSczElKAyz/EdXgZ1l/2zh7NPPLIN
Jo5CexV6c1o4Zh8oVMpWTjPYtzgGi7Bw5hMQVS2Dixt+tAxGZpGdqeGAk2nKKzlP
cby83JFDtMN6J3O/cibHM5r60VmolcBkKzE7xC1FbLrR8XcW94j2+8YUny2leJ+V
9EWVSjptWY2PDqSWxRQnltkmqkkdJdSzej21ALgSM4CTEyWRxmpclv7ymiVDGUsA
aLyf4BQB5F0fa4FSAGrFZLq/PfGpjNpo7s7q1VsDQmfuNSQRnjp/gkz3nIl06tL3
bJQIOCIHi/3FNiLcmMF0g8r47OwdNZWYvFrolb1r/YZ7ejNvwZq8taCpFHKd/j77
m0bveAmWZVm8cw8mXm2c77s8uTGvmHZeAw/m6GQj5pFHGOFDYaOsTLzGK4nMOqLy
bnVS8DJZ/o0z1UE3vc2bTKTb277bfp/jH1m0DONTf9vbsjAahg5mn9zkWaO4VnmM
zHhn3jAar6wfcMV1xe4ayO+tO/DIycMl5uHJQDC4ZilIDwLsi71RHuG+6T36fq7L
xoD+Ke87mT5/UX5TXV6KJF8zBZhjOIShEmYbw2VNjFl58Afd0cG0j1wCn4Zst4sD
hctNxFSgKb4Xn+hclkEU705sW6gmM8muzBzOCYFwbqnuvg1upg+E011uHvb9upi7
MaK9upRjxwHJBHMhLZ5kAIxWuREwMz/1w5cU+KCE/FPqPJvDian5NVcJvzkoGrdE
05gW/UptoAOnyzbsjb7tr0QnDkEigMoCkusB7yuB2x9Ws7n6LPdOpt6sour4yxdd
xWvO/pFylzTLCQfpHFejImxWeKVAA8TEBGRlpl4VkPNU3p3PyCyo+DAWp7BTum+i
RZsNsFhgGdVPQq54DsEXC/HJh7Z3vyca8MrU8f0hfCm7npWm7JhCttFi4gvcTPgD
v1U5PUP3uY+tu4Cvz7m7+jTA+mfHYeOTV8WHvGIEbXlAhzYhmcU7rqvjH5aOVo6O
x917WyifuB3ih6oYc8I9hez+YPoGcXmSxYg6NyxbXumy9JA8AAq4jCMzdQLXgw27
zGOJWxyTzdbdvw0zJ6Bk5CdfMwm7UHWWlzYoeZ2XrTg5qaj/iXGinoVj44CzkYcL
VyQCfL4yt6lyNRYYq9JqC+TPhF9i383nmqCWPGvr0UWvNSb+bmJHt0Qk9RJNjizm
q6WJMwf2CGv17MJTiSvBbP0Gvx494Fd5sWQv9vgF7w9wOf/e8ref5+EH37XAdxzV
JEKjviW/ClClC8h4SqCrb+lHQSj7ux2kWo0wp/nvxq7oobIuqIna7gEn/oaWSGJm
Sh8qi84pEwNBoDL1DgvWTKnaIdsyCY1aObqN0uySahWA26/+ONFzs1ENN/cWqbTG
NfgTs/6ParnX2X7fsO5CiiTIq6vrY8ZnJnlXpppHMHz3uJXURutGjur2Trj0aO0C
ELSkzU0f+GeuruHaJ7/qT0YPCM14EiyD9p7x/IBzhw25i6+K8HcKuRgUhhs47XUr
/oQp/PQfQkloUARfti8oyCUS4sjgBCd3ShlerGLLY5xoPn2zJRSKLe+jGNIYY+rB
/sxCHJQTICFyETzu16q/Uu8NDqxI5r8o0n2ret5jFg7Pb8EV6ttouTQ2krQ36Lxf
znKKbzVRizSEGlJQdQlOX50rbwvhUCFBNCSFd1Of/6zhB4dN0CH84NXNlJQMH4nC
HqIM0Tr6nWXgUcg/vObQ/7/UHZ0fRS1PwTOi7wXi7qIX2kj7MbYZ+4K6WA/zJokg
U5ixgMuKD7DnU1/k9MT/l6DstzuFRsgucFA77po6nMjDUUlrWQoN6FRT7SZHgNyW
qv2BGh+suy+oiIv8e34yASmQs+l/thVykAG5nFkzZDMhchSFdxDMK1HNpN3wOx0L
jDhI119tapCacPaIAEDnAQbgTr0WkyF2eYWgjajSeYAfVfzDkSyxNCLKetZnDb0A
pSHSySVoTs34IehmCCdMYhScmkVmvzRJgeD5xKKv+cf6O+IyNDfQgjE9jnfIIu7u
9x2fmZNKMNmKuCoYMYLoqRQ5kV28brFvIYVgJLpcsimSshRdeDNaWZ6aJXF+YLc6
T6oAk8EH1vPEa8+h+Wu3Fvxd1SYT2ckr51Qzc1Bj+ZXnXHQPYllp+34KOASVJYZo
7Hxws6yPvTo3+4GyM05eS9R0FpFl1qCcucFUUo41c5FGeLVguDahLk7muZA/fczH
B/M8gI0voZXm7JlbMOsrJUPKKNBEgqITDtBLI6reAtL9NDF1cQH94xkUa2jLKxeG
RMaY8mFRxDRP6nkTaxMKH9JrkAkkll9glj9/03JM1ylKAlE17bSdP72RD5JT/sWn
mQyQDIlUl3yg/XKdTK3R0IOggv8TWjEJojvm1d+O2zK9IFaylPBXyD8BgtrJC3Ka
ceT35Aex2s/M7OO99v/b1proRoqXvkS4f8K0jjFaSsTgYukPS0TVHWcDoNh6loNM
DhQ5xMcKG3bSI0f5IRg3HYXmD2m0KQNvX3nnxONcG2r2WHT/6UI0BRWGzLdQOqh7
ms9CkY22VHZa2/c34LrL9ZdUE7ffDQxgPgYExuioRFC2a0QxoQLvfjTHJSncgGZK
Gy9/cqBzpk1doU8SDskiumr/uM3mycL6jJIDWVdyRm7+VfIB8ISdp2uNR0DJZ+ao
1qHAts/q6ywqY3W5H4MRm+d+VqW+nD6hSv8bzLrK+ofig/ILeQC9uoqaT4CXzQcX
jAj4q1t0w2J967lG/UuQrCcq0BhC38c9Z58hRZetE/+GGLv60W6+y2spju3qM9iH
N4Uod6h9B26hVLiJPUiDbPMATeq4zTXpJn8X0XTVcUPlwMTcghQnGi6/SbxTR4Rq
qEo6bE1H8rVehdTMv4ndX9YmlWUs1IBSupUUGNLpoXwytmiYYCfPAQ5RvtZhiBLU
qD/oB1lTuYai+V8eMh9ZjbBp0Y39p9BIAiaeH/RBFanet+mqgXzWpLkvjL2rr+44
HVySdIdosSIml74DBSezwUHZeskawH7GcUbbVEgKVTxftmwgC/LlF/jdVHPFZtFs
9s4p6V/p9sVRWxvWhPgSdvhLHdeqcET6XyhPC8OuO/mV8endMhiZg2pkCEMsf2c1
sL1D2bJjFPFucDvglt4/FZbBJU4jX9W2QpGy/Czm/KJX0maKImRZsipAYIOCA2sL
/Skqb90m4wTDAKWQUFmwwCMLU/7zRaq+O0Z4AI0MKAI3KJoepGuujnO0AfJk1Lrs
l4IAgXahvA1O76tmXqB5Nosu1UOKzf3/M7H0Jq4tEsiOmIhtDCcE7HnGIzXqGVxk
GbPNExlwIEbScZdEFxMj/h/xEkzBd4bbutGgSft0+pfoQBoeS7l9Il4SNcmX+CWX
BBcknR1V2vcEGIfnEChc6usw7locOcT3JSKUgkusS46QXizenq9j1CcpPFzhFNgX
8KtOowoTuthFElafUrm6ocaQfbXpn/DoKG9i2DGvoYPkHKNC6vIvVHzNz5IE4pWB
ssVXDvOIN+AXO9Quo51EdHPRvqXKDGEy4hZxA+tloSp2/EH1RiOBimk11p2wZXiZ
nx6U1iQSq410KuerVmb+If1WCCcFcfKktVKpy1uUoQaSZGLkCzZoMiDHxgK5v/pd
fKkhx0419ZNGFiGzB4IPTbWPjvHkqRSkvLuwS1zZPHn22SPwlpCroYVGOGbTzO5R
kN6vL6LMWv8R5WP/vu6OkiRKA3FiLv2aZprBg7jlENPHvDRHK25rYS91aBZS/yKE
BfgmWwG+vLgEfGSudWHrX/7e/q4AXktZXMRHjwS7pxoarHLSU7sW1zh2yX03cpXi
cORQ2JPL5N/Uqzutmdrk2pEgzhQIIMDhy7hWwBMi6JYILXEWs1uXOhlE2skZVuTQ
fKFkblDXRROGOIDLB4XDpOn0M7LhBzYF8JBVIDUXmWEVVcQXiIKV+zy3FFisFq/v
m0SbcrGnlEpykp1eILjK9piJGuWEL7INJuEFFVcIQ1Pyc7rFf/40VhEBVi9HEdLd
KBHEeFFSygu1or2I47Vck/Y3McHaAog75POZcNORZhuSBTQOHwPyW6H/ZOViYqlh
D95E0XyYSGewIlyvbuPCDr+ChQn4IlFyJ90F7Jt60sLDvkgi7+coDY7o2GP8+PiJ
daGfs27Sy0SXjA174YpewqIQLiN9Jp41vYHc8a0dJnaIpVwtOcpQWMMXu1g5iZg8
cTU0ENLiQWU9Wcr71DuebfsWpNg66qEfUxF1cy7L8FIxTtQY4u1bBeyHDYudDkz7
r7MUi/7WezuVqb7pABdoH/9ZIgllnO4FugcfLpku8+LEp5D1Ifmov5cuaSRFXPws
lWYrMjr8gHyFTmHiT5px+V2vedG3toO/S73vPCVNsiVBQi2fmSDf0c/Sar5ZFyRb
8ltgGuvqyJhc47WTkpw1J64WIE0Fq/ArlRZXj4mHJTZ0jNCKEVI5npZ6uH+C1ug5
CgtRJrlpOxsrOyiZ+H88BH9KkQvi4sAwv3vGaSzReamVzjHmM8lk4Henxt0xG+xU
J9DyP5vnQ320qsUB0GPCOq7bJqquR7tzWN/5ooMt3rxNL+FGgQTAQDZZQcVW4TRW
VVF8qsxbQtJDA1wzLumO0og7Uvlb2ItXn1ZL3XmK2vTXE2RlTc2f5W/B5v6pXlTA
O1+XBLfDvSnLTH7rtzCJbiNb9DhVtmTcVDn8dyPRClpP3W/egMH8Kvolh9Uezs6+
vkrxJdzpUcPOtkux16d5f/kzVHyhl9i7pYErmiLzOR2ZBU6CUuF4+xgzeCLvPTjc
+gMmt9fiZEsrLkdIKfkKR9fl13ZVCqAtgnVMwrUM5t5S9yEhpDrfWbaxd3rI5/8U
sli3O8vhaJMxrpWQ2Kr6R/ct5Kq/SRyhEA8rtklAO5JjdJi0R4i/0Z2/q6+gyp7F
Ms20Hcuh9irE/PnVgeXlKCcwdZRmbct8e1LCmqMgPtInqA2p2FwLjd584sIN2EoD
XIZw6OhAecmHAygr9pLdo7w+/8LLj29FwFwRGj2PGOa7WHoBe/sZiKAURzAK/JVE
yNrZi3JFnmO2jkIE4mGf4Tcji5AJ97haUjLV/SDb6dmdHVi3E9Et2PJ3eqWTMmx4
LuhMSsuZNBn1v/564Q68P5J3FFQS9jvRmgOXncOOiUa1SrsWlcs5X2o6SMJHUeoG
EJ3s2VdShnobO3bs6O1EVbw+Km7xNsMbfx1F/8loHpw35cs7RaW7CTFEoOtnDI1J
9c/f+IU7dMhS6+nXjovD8fIvF0tKEdjuIXQKCZsP/Qwo8IaOupaq9K52SV6Z7GuO
zTNi0q48VUFTS+aoJeIFxqobYGvR6NZvmY3S+SHrnfDWZgL8tNb8da91GH8RCNS6
2XpAMbBbkO4VrbitnNmJdtz+JYPRtZfSxrKW5nm0oJgbvPCOZ+kc9Kb2K3AdMRk5
U6AEbuWP3WlUb9vZ/m03U9KQK4LMLutYW5+bIKPD8MY5FjMMUL2YG6Tq/I7Nff1B
lX+B714Dnq/GV2Zww13Z7bDJqUvWMPgAU7TnDh7x/emLMsfNHr9AAvQOrWn+b5Zs
kWzdff7PrZwX4xH1X9iPXBMu29DU3/hv0X6FOYsLepjmrkpwNnQUVQVR65lUzO85
c5htKdrGfL5WqfTjpHg+q3PGMpqbwq6R+lQDpsPojQRG0zBN+uHjW5LvU9RtMVSE
wyYt8iKPP8LBF0HatxBWZa/Cm86cOXpAhJV2GpxvnZvVD84CSN7teTRtORQbfGw5
LNxQnsraFmaxGfbOLaqBr+Flbqd3tWcsHDsivfesj1fDP+fyi92HlToKKI0t3szm
nOWVP8j7d4cvqV7LgFs/0msLZLW/Fxzw4nxcqcK3Gshk5VA6zNBdMPMTfqvXjzXZ
FYvZh0/8VI1iF6dT+VXyCRjcBk4TErJsLHGjW53Bi8jILvmzNvGSHgbygy7CvXly
aLoNkpvpZvBrUhjNUHYkqWwoUMc3L848gzDQK8uwZSwlzq/nhjptA4lIP/9nvMW+
CjRAwt4vUbGgwV2YSQ1zhwGRocP584SQhWc+f++LrZQ478i3gtmGQas4LrbUHVu2
NAYnp8BIIGpsl7D9xD+4Mg2YfCJlJO43rki7kArnzIaIbwx1gBX0j0wH4ByVgHAS
S2aa5yYw3yH1uo+CqVMICOmqTGgw8EW+ZCAofjgfCk6NzyC4nXXlLWGsx7FMgK6T
uNxW6Asj+jFMbwchv0PftimTo3syUEgJkgfW4DdPUcw/+EtIMFmoYj58/7Ec53WD
PPB+OV0Hsjy/sZqpRRieOSPvZfr4cbj13yiJ1IFGV1tn1Y9rBSAc7x5y/9KKlvFA
dGm/LnS1U5UoUj2JOYXREq8+wNOPcYVWYeRNSwyfoOOd92Ta0CgY3oLz7FGy4OgS
sUYza6AmKJjnEO7ypdVK1UBlaoCl8NHTI2hIvGgYxJAlG2HLfU1Kr4wk9KFMO7Wk
8FOCnqHVs2yhoOWS28cpvfiryfjmA8jjYAjglKxQrXBiilnJYTg/KkTpOcpT+iZb
ZepHZf5aqYonlKKmpIsTDR7bOceTVD6kf63okpu53WEA75UtI5qprA6dlaJYSYV5
ruGMMsfN87X0mE9gGwA/C4rZrz9vc21YlLG78Mt71XqEUaFavwEAQ+ar00faZXC7
afwYmvTCV6vBFKUSx/0oKdI9wD0vDcqEZs+HeVJ039UUbnxfXEQNeAFtT/byDuw4
RcDqX7krkt1HqJ1fOnjFxAmGznkFJlVJN+rX9qnwstlL/OKzKkOO+vaoGrMkQzcU
A8m1T0zhVFpKhACx+gDuKQqDc8oXfQVqIe87/vNFXPlK8fcu2pLZOH1Jr3i20TrZ
lsZpUtjJQWsDaGV0E3H0gl+auuTzrDkZy20RK4BzMjCb5ESaNwo2SKaZRGOPKghy
TWu2ioI9YuIexlThZ8JvtaQmZRHmS/hUUgglYagU+2Z0cb2RG12woCYcoIM+EeHt
nVmyo8fad5dpRZZSFkcRkN50qM9FjGObl/TXQNq8M1t6bUbFRqxkWRFWHZ67z2Bt
Z1aAJ0KpPuLyNvP+fmKj4++OM8PbGkQ/J2Z6kBuqpzZ68iLuCLKSZfsepKuNjJcb
0jfYcR1ruRtTRNZ2A7VHqglydYVOFkS/3BM2WeYvJ8XnzXAy5XfUPsNTivNyFRrj
hzPz+mn01pAcTB7yGCN12ikdyKoqy2pJAkIAqDmQ7eb+5KbxELeMB68RaLe6UvzX
2dFx5OE0a8IY/N1VC7nu8nqmOy3NdkaUVExiZieoc1hMIXMBHoBL6RYsOAVAn+ZM
wcjN1AAQEZZxgE2AXgU37KC//wp1DLQ0HWFkoJZPobas1hhDEWRCxeyXJ2d+s7BJ
We64fJnFsQECHVDuGThfK7yJbyodnYItd6zBlVsnYnfaOz0gVf1w2WcV2tmaRZst
yA1J0ioN+O4JR1W3SDYnXM8Jr1FhSRpBEZrLUxVy9I3D0eyzIRXk3aPt4GyHsNdR
b0wLEHgB1XocOtgXf73v2NnWW3zg0TrPT1BNMcp0GCgW4TbbhZ5sLCxqMFbt3U3J
08ASyAro8aZX7cy/6JTziW8rLns3Jt+jKa/u7BNWdsnW9kQEJxHyoQGkdt1BhaEc
mCBOXn0rEiNBiCsbOaLErg1KffY+I9eYONpDAY0ZK4zbACF4uNxHxK7FGlAFJeuE
77PahmaON6AC81zZ9KntP1WG/Oez063zHr8CEFv0FiatcQ7+K53JmY4BOqorSjlu
R8RqFZV077xyM8CuoSozM7zFG+dugj33SHvHMy6ry8OPpCT8RIU9jyup2qntK+0R
eg8hFzdcTEYtnISCUosIrOIwwb0ZRyisEGMlpDrt+M6emnVrqNpyqZuyemY0EYnK
7TrcYAsTNQgVGOQqtvTNRYhYASwHtBLOvOlwiOZ6R9qb/W6vxMJ2aAVFvB1rEmuC
ME8ylHxeX5zFo8tyLKu4HGcCdG6r5unSLAfaHOaICcOHLzTSAsMkHfVIw4HfIoLV
ovd48DuJx/oBgK9HfJGSNlOqJsj4rFjb5G/oT0oYX8FOyr1NT343hI1GV/d9t5BL
yPwnmORK2iYeorBSBhSoJy4xw2sfoEUR4p40ULB0JbU6hQz0plYvuRFaNx7R7ik8
9vNJzAic3Z8vLmuuM/DlMyUSeQwdBonkUpVNIvLJS8foFYvslYMVPNtN5OZL0c0Z
OB3VetxHHfASRk01J9dU5wuKbA6kSgGjxvQfhLRumTRt5PUsFRya2291S/Xuy/0h
CJjW/JusW8HT6j/0jijWk95jOcbmtMlXJbtwzLLfzX1lvV6M+1WyN+FFsR7PkrKt
qqM3b55nouNObkheff9kVB+f3r57bnRKac1q53YdtHjDsJ/FQGxo84A/epLTKOrW
VUQtj2GcGF4h6vN+hLC6pKcC1IUSZ8z6M4b7qNVF7h5bVK2V7bjrf5myuQg7kTfZ
QT4WuDi0wM/lXmYoJ9xIaCtGyqJay02iJvc/BjBfpocIZf24cXQY6TRQisFlFAn1
WrC1FmB/poPHmOdtDsayRfXLqdqPi3iqCBeGKdQa9BTuoXwKmQ0XdJxaHOBXe3Eh
GkNiEjHRd2oAkKLaE5uGffza3Hlu0YGG4zRBsr2U+CfcTU0y9inm/69WBBI3Nm7o
27juBITHe+9/fEf7T+WwxfL+x+N5L5kRZv561wZ0KiDbQX02GUaUCTHenD+fTJBS
0GsYzF8CM5Y+Da4rChSNB5dlOrDPYm2RBmZ4a1C+d6JfN3y7dJm0UMAJTi8AvluK
UX4y/7TvgYaC8D1ieDvKnVUurmt0B5gKR/FWRfJZUOJ7Ah5pIMMTRBAiQr7kdMAo
zJ7rge3ffeHgf8nlhBOqT/1+Jf8ezy+BixS+XsNl6zPuzYqb0s0yYTMC34glEI5f
/Su8j0FGd365LVHxwpeW0X0ejikyTZTQHLuoFW03hBPWpeRCm92vrOGiHPJ0HHsL
pElJ6Mydvq/1Y0IsDe/ZRf/kYyg0fbfv1fX8vt8KCtZO2liZpq9Woxl5BqHqtxh0
GittF+XsuW/PTSGt4NgWRfnKm+Iwa1/XmnVsOtI4QAYgbv/XZBY81xoy9j20LY08
A+PMHGnXTYoYKBY71g5aYXirjJIi7ti7R6xKtkDdRSgdqnt7Z8ZjvIS73zoFLT6c
RphQ85lRVn6JDN9R/CGi5eQ5YAGY4QmiEQ7HimzOtqAms9KYkZDhvhA12j9n3GPK
ZcVEn+/OdW5ZJcbo9+i0rCyjT1CALFJvsO8PeSAsYyZ8J2Vj2JJR4a6z/OPg+LhR
3cFVtZ2ltPxb0efDoQcO1enBRf+80rPBgQHLe22I91i1XUX8nB9nSiCGpezqKd44
Do62/jZG+7xV4rHYCkkFAqmcokweLh3nipaz0guRIWJFYemIxSfDh2o0uwUB72Gx
dEZt0k+b7NQD7lgSCdTLTNqmEQF4YOvduMPBX/8tROuksYA075EMyF+nl+8wg3RO
hAKHyrW4b2h3iqWn2QZMMva4NHGciXxpIMRRV5Q1IsgHOEuJPq3gBz3pcKP8YDhK
Y6CO4vUHe5FUY7kXeqKRKvaKmQBTy/tFzlBVqbmVVQOnmei57voBjrZ947mWkHqp
epQS5xkFr0z5722ZjgJPTbHOrsFzxw5QMNgJaWSrAJKpw0mXs8gOcirC64g0XvNN
3MrxiSTia+3XoQp4l8UiQYApTb11dUyCAtSmEUSn9eGVRJ34oxJZpQhpBygOfntZ
yJrFfoNFOSsRCgUpNEc/J7Xz3hHZGsz7iItzmIUQ8zV8HmOYZQpWQ+baeuB5EznU
JwhaQMGETbU6yV26YKLBYpDvWoLA7qd34yw5QhvyfTno+2S8wFEJ6zENnHYqe8LN
Iu3Naa8QeOb79TBsIpZA41DM0w8Z4gDybRB62Fp7BtOFADm68MbA4GgjbUOOAbLg
ZXOLcr7PMgJZSOj+HLE3OStuAiwfOCDNLBZ/5+IMs5M0kpasTfwd/bfGoTwPN8Ro
jRI1iJv3kaTXS87YZQVocBsO+NI9EW8ZuEKP32a+xxQCucJEFILUCu4kucIwSaeL
016mnrl16l3h2zQZYYuEgAXfcpvYS+Z8ys3wtI8IZAR5PDZzxJeceH5eQL5b71Fd
TX4g092Ep3Xqh/jEL85wSu6AgqKxI8+KLmjfGIHBoUsuhOYohHYOzSOVeUkFhno0
hez/gAGDVt7jrndv04Gf8PUP03eFrlllJhywU9mhhq9sqNAiCW0lXnVhVlK3iWnB
gV0aKNWgwTndc7o0IlFRI4FjJXiBaT52w77XEBLKduVmk5tYVy7mnAYvO4ItEGk3
0GEo6ykrxDNsjwKfTi7QUoyDNLL4ewLoC8lIQeRaQWOQCwhrSgXXshIndZ2+SaoY
w0jDuZZXGZJqqtGjprhFErqkyfs9kzTDDJRPLT6j43n1jefjLD6qPv9gXOcVt1F2
UzNtkaHgaYv1cYmRZ57ivgKeS444mzv18TosBv7S0/75C42l0vmr8jBUqcuyUoOX
kVNJiV1h54S8zKbPgJtOdVjSP3wXRATEuCmv+9jjl3koMp1qrCy3PGpBtevIp/T5
4cwzsCcQCcDIcj1iYOrulKD9UZQhO7mSqlDwYhJQcY+t/sT6jIAuTFPFOSueDBLZ
Od3zpzazTBOGHrqOt81SuzSe+aKlujIyhBl5cZBEj2qKJ3ADdPqLsKIqkBKpKAGc
c5byc11tNfKFPKOPwuO9womU0ZYKheKfMZvUev07XFQ4x6LGwRGFTGdf0R1muTXy
iR51WJ9OcFnFYSMJzXYQqY4FrxDkLx3szyjM9EbZ0sbHMNgu5nQCczrG1+Pgs73M
wMLENGRlq5ePPab6EEbVA8Lqh/HPmzDGxcziO42pWe7ZyR0eAvBhauUytVvv6+yB
ESMJd5wRyebJof68P0OSeLWX+cY5WkjcsClpQAluEtcbFLLsi3gOup9Ln+yXZYFE
O5JZn6cgEqjjpJ0e9eGJ5nazdehM7/6TyqZ01LRK4zpURqtqXNYCSaK7ZDOwW2q6
ZKEyQUme2GazuCFdzA52eh0weChKqneBsiB/qpNcpq2bUcoINqPdbIp7pGfbx0Dy
a8j/ZFGhc4xd5H4+uW7gao1U81jthGLuc9rdpYxAb5XjGurtnZbhYXslvQoVVGTt
WhUpkEFQhUpERk1BPiUTaq5LWYki3Ono78+GIwhK+oocZz7I4ng72nOlIZykhdFA
R3/o1YN8isPeRx65OA4hOQfQDdNREp1u5X7D1wozbTpHZIeTQlM7vSW4byW+RA6i
MpcJuGHH5TiHXsjcPx8wZfhVbnO8BrCZezfLT+V4QyMoc4wI+3RxhnGpcMQ9j4uE
S9wUu4ILlb1Y+pJYoCkfqoT57TdFpUhvS2uOBNjcGk8BXo1iZcIPS3kB5p/atbT5
aBa7X4t0PSyrjD4+oV5oKLsHA/s24U5Tg+t4AUyAam1z34LyoxA6E2z8jiKvZS/f
mmFz+1WqC2LIBYHb0KaBrzuwxTzgYpwcwIJXlcqrQkUwa+0FvXdSs6OG3BrvCoa7
qGLiptrhrS0ro91A8ie1rvw4qfD64ddZWdd0uCu7T39e46Ta0OMExvZ9IMVq3csD
igjQeJ5H/cmkf81N6+ZgloJhu7x0ncfWeZ8xnCCquXR61ooBJ1eN1Z7o52KLiubX
Co9AR3Gq20udN+oPofrV5ZMLtxABE73VVIQH2dcrgb4HHrJlqzsut81y8ZqIk9Wz
TXspuRgcYr0yEWUaZe0eTMEKgppKJPKvpDYH0/du48+A7fInTeNvvG1A/W8ZHE67
k2jmTJ+ZIWZpxDhGiHZrtjS+BaMAEWpjaAex8E/yg9RfJqwkz8Fqdurud+gubpby
oUK3a8VVSAptqOalObFegoiLrpB7E5FqXOEiVtnGHy+595f6uKCaLF1fG6svJKqi
EY9TYf+QOmLFjJ6BKlJtXYmTD48OKcmdRcYEmUHWSR/cu/f+kImSzg/pGfQ6S9Sw
3Ukaamv/MbYv2wBriocFgV5PDpK8hvXA+Ttq2CAKbUiB5PYyKBNfuanCRCZrFToq
2CMnZBHIiygsAn8Y2eqkBhQEtcBUDcWmqF+F/UEbqtUOfKLL3VUiurZrsZ2Iv3xp
iLc35F3SnS3VV2lAmgcIkGDiuZPtXUn3zRu6OpYJrqUl9eFB572pPEYWI8lsaGBk
z76z0TIXXO3HYxkxkCtbImErPYy2yWUJkjtWCTcHCm2Kex3tH1rlG7UJsm4gRk1y
rf6d5n20aOJlD0VycVDcEr0Bd56jEsYtRLAYQQp1EOqXRTnPq0Zy6gnk+uj0TEMU
ZIvW/R4ISlysyzPIFUrLXCZr5LzGG31sSdS3SlbRpsnXA24N9amC+aBjnaqfWFqW
ZGcSvLel/OSj/4U+aGCoePLqpszRFA22s/XZOkuc5JKp+R8WaPjisi/JW2rlxG0w
45ZdbetPmyy6Qw9dQBzqqMf22XynSUywCTylJCYS1pMbegtyDpfXLE+TuXetFn7r
pc9x2ZzN+QgSc6fm1pq5tvz8qLsX83eAg0PAn4XYZ2BVacwoF6BEc9WfEn6X5caV
v4RKpKm0IwQpMhZgqetp7/c/vmK90rcwCJLZdwMQTMBnh696elhPYsqX8JSzrT3i
2fmtjSjpaQE6R51qW5NzZCFESBrkKa0D4XTGrAFd93oIuGrDaTB9zsok4dWNPfzU
r2y+mLSDLUUGLAk4TYdAyPxlN78SCtQ8PraRSJ04CEnukUJ1yXhSp3MhGIGBdUEt
F+t7WpnY/9CWfOAIDN3XfkhbltcwhJOqadHJs+1aYaSQLdTMGDxQ0mx8sE+Qc2sq
SydK667E/RtRQQPL6NqXUeq4QeYMKgKJBEbcXDrAcLgTxz8mRf8fzZGGIsHXVJ+f
7liPJNw3srsT85WRzO16hGqEnC8H5cwluSC8y2UuWNQvFp800DT631uVaNmNWkek
FqNICyU7+X7m0KKIOjSTPw9jUDrwRDVcWIEjAeTxYK4/3zL2/mUPqvpZypGitwZ/
IU1pD1bqyGAlLAy9zo7v6oHx15LZ4Vl9eCmZK2D46c0ZQGCtJyQYCigOweR6yKHT
QAmz0VL0HvTiN2P82ebIfT5f3woUyZdVoeVCZbyYqfvQhSF0fMSl2a0nsPyw2Ytl
rfgsQ+rBcX7PIckSzgTy+qugkf/OkkEFfemU5J7r82Ivw1apbMVQnmhcfIUALPNR
o3MuP7IsEW10j63U65Vlg09SvxK0/Hop95F5EhzOw8ee54GdtXKaOUd/11KUvK5Y
D8BGnqDgdtyO7YsH+gjk2BUnxseCK+Y4RHWKrwb7f72gXL4avZd2tavAYp7ZUFd6
wJ2hl/lMW4YaRbBM6DfCGZA/N3PhHfPVsxH90t/8HC9SWpf89PtJRmEG9OWY0KiU
sFOTq2e/7JcTMrKDa00/gVN42mZc8BCR9rSIWjdwyAD8XVU/9nPBSMI85HHpbC2R
PIhTWk8iZogzS0Yk7vGdbNbAKl8+J6dy5YfhnpdqmyOSPqLVOJextTVZQNS6F9jw
1JHxvK9Umzdv9Q/89UuqfB+n+P4PSzp6DvfUwhccKBs7RDQREy74n/qDM+UhpIPB
LUnxhwb2x+hTrdqqsH2W5whIBk+fjXwu/wi4gSNTypaDJxhJL96Vj203k+Y2Pg0E
CGpw4YqhwHvcOmQycAbdMDn7WtfuUZl4B1afT5HbZZuQtIypLgRY45yes9U8lnJD
4zhLerCJVjwA2QGmoe4SO65n0bsdcDxhX1QcRTfFATlMCiqJTvxG9I7EEzztH6SU
13jpOLL7k+KCs07GZTc/3cpet929P+sB8Kk5qxR6UMj00NNqnyPP7DA4iLW3nHkM
cgcEkvDTOOIKeUwW41pKUUKx/xz6EAhZw53nv0nMQrUNv/El9RaGWjswfRGd5vj5
2j8OnFmLLfEcBYbeBxU1MEh0rPLu0cm3H1GXtQvlV+KKVux9lolwb+EuqdFz1O4h
vj10RVzf8u3yuZksGq2yDM9FIR8+X1H13LdA4W2QR16x7K+/L8ik/Tbg+WJIfqvx
2SjTgeySu2F7sKLIQIpPraUNKbeAJqS1Qrc2di5pUQfC9uBpq0PU6kOKRLcZ95+o
HVnE6pJ14XWLbzZ7WIL00VO3pPklZjIauU6Dzl10ALvWgmDF0rnv4cofOsTMiRNm
sxSo1MtLfH74gxzBxRT/6Kv2nV3CARXrjFkAnT43DgojMzmoPBVD7hmkMqZDlK/1
wF/IgCRBQJnltneJ1vTmNVNtJsoNYUnykZE+S1ZvTtsFPOih/iKUgOAUntI8jqr2
T+899hhgMbi+gvUFZgmZIatTFPC8CK/RWr5egK86F6uJ9VFbJAu123/KqfmnXnuv
HpK2xZH6SStTVvYM36yQpssTjAW8C5nP8A8cA9WxcDPkbAL1x9V7gX0N3CdmKCYe
iEGKvOV+CYGBnPjXkudU2BjM49vgSJjEvgE/G3PfIwSMFjOdOetSaMafdH4uAKjv
oV8PzqmnLgGRAvEzFjFJ901cyeEifyNMBHuWLY96W1gCICu/UYiJUgPedtj3Jej8
QfOymIcRxB8Zto6JP9p5oBtrHAJrXjC0Uy2uzdaRwWDS8DD2scib1/hN5xRn50XK
Aga3FriB9yw/FW0M8G9cZTmgcfg//cKEjsN7Rh+M+fJijM22+TsK33IdHmlVKpnZ
CySUc5/cceTeQgBXqxfYtffbxTf1XXedAsWnVbLxY/M1eAw4b3LwYAu7P8UX+TDA
TIfO2hWdolTWeo6KSmcj030vT+joXU8Qt83/fM60t5bQuPUBOE+qj6wcivpvNSwT
dOXFroORavVukD++Bh1FS67k6Lpk3lZBIAgGgTA3sVO4GT9b1ADwAXQheY64zCYB
`protect END_PROTECTED
