`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveO1eVONt6ipztnbB5ycXAUhoNbMeKMeiDZDOypGNCtYx
6j1ORt9yb5tvDs+69eX9HK11OaN+Ip2uRNMyqnr7I4Xj1QrpRWoN13AbugP2zruy
VMYGu2MXu2Ohmwlm9LK1TZLjNAVC5seeVpfL+ls2prh7DqJcgHWAIMjfCl+3qojx
3yibKNu5NvEHgx9SGwVID4Fo9uS9XxhEYtedIx6GN5u5gY10mk5PZBDOdBV7UYKB
`protect END_PROTECTED
