`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
if7OW3neLerq5QTb0GME95jJuQQSN60IxjVoaWgR2Ew/Xrcji9UQY1QkKkghydkT
cfZtN0t42oskgxpOvhBiqTN/f0p1HsFQe2osutDKM0HTcHp6qcM/eEsKGjSB3w45
//jWP1sWFdcgcKRiuUtzmsHgTH96wt41Md3Yu7GYb6KSFztZGHsmGt5lVcGSCYmp
Pb4+wDVxjbch5i3PcfDXKxxoE9ye7qPVrt65gT77lnd//viLd4clO3Kvvg4YaQYK
Qepu8iXopSwsUC6wbLt18sQr6aNe+w/VqO4116ADZOtMuXKrNkqJQ+t6FXv2UryU
`protect END_PROTECTED
