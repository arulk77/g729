`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDmC9VHYs88Y79f4zRi3DR6cB6PJex7Tmx1Fxfd/hp4o
932wtFeoevJfw8cXXhm5yyEz6R90ztVZYfgce8GJL2WuQUxeg2TcJK+ABv6vWTC6
gSbP/Q6jTuYEDGpu9dL/HFkGYmxKK4mY2ntWteuWMyGcQvaTPzhGnH1Kb/YWgXiA
`protect END_PROTECTED
