`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIGVxFml1JW3MRJbjSEXqJk9DpfeIUfar+kXCSkRwtWw
nDkqMkVbCwSWQ4exR4zBx89hviimHN8h8Cybm92T/rX+7R9drnaPydl+fEB1qIQI
bNV6P9qnzRg9q31an0TXF6ON6+c3o0TyzQu4+EUPTcHH+Ybe6Z91wOUvRGvfLJEF
EDWvwYPJMLNlZZu6Jmdyu+Iie4dfs+ZYs/ILlfWSFgQISTu1ZETiMuANYkA/R8eZ
aOwqrBuDth1W8colcVkc1fois6xXd+8SjQN578KvuPZsAW8jlSQ0GhuXkznzUMHJ
KzJEuGgoazFGg3zi5Lsncas3MMiXiw/ocZL4LgKbarebZBEjzIa802UegDuICWsD
ktLD54vh6EKokQEngStQ3NV7FA5uF+scrBqCoNJ1UcIRGK4JVyWtlXzIj4s7YGid
EPnWPmImAMtvYKSMYDjgzXQ6e/gocRBBjQeTQtBJ5jUu2MArrM39lmikvytuae/m
XhP+/f6Yh/Y2AAKLKdo3LSaw7EH9vlnY4tk1OjxVMS5wXlAPbRqYs61e/c+tkx89
`protect END_PROTECTED
