`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAadB06zBOSnW+um6lf30TkPSoubAytJX7Ir6Dd5TpN4A
txH1A+/rtppIkPPsuoTGzTH6HKbJbToRSZDtrkVjTPzESLRgnbRAKqnXcSgxYlCa
rwzWpnNoqpx/5JbSGv5twpVlTfv/2FRtCHv4q4fIhoTtN2aECUMMRrLC0ErLh9jo
gD9NMCu8y3e4crVhh0+9JuE2PCZ7rurOpDyXtQzVMo5c/5tF13477SPsXb36Zrhl
S3gNAZLYyIS2k3bElQeB1m7VXXQVViqkid+OpOfPrvj79MFVM6Fa0oty8aX3mi5C
cl6NoIXe0oIKe9pJq37vcRElcuNOQ7Mncxh0gL1tyKqnX7oDiIh85FwkS9Zcv/hO
FmlN61SQ2B0r9MPhNjoxVU6fdXOPSi+XglX9Nz4VvWXk3AOQiuiJ9MjjktAqX8Mt
70M9HZZ9P0PW82WF9/Yt+J3Xo7cykJYKiFytcNGtBRRV2hk3hujnccNORLhHjxzH
xd6+/wFVCmMDXTPwQnYged+lyuMmrKRjKBV0VraKVUb7cYA0Amzd9K9A94vZEd+Q
5G4vlUtrl2XtlxZR54AyynAtQ+EfEaQZZillY2k8fbK0kiwlRsWv7ze1lMvJMesa
zho9qcF8OT0ubC406vYYz0HdXEY0AUOOnYV3/ll8UIGBQDRheaw9d1xAC5rH0oSV
F2yN/C48515Xv8jgy0n/iP6kFgOo+f5cJpumx2Zgm0EpYYZibg8rKiFPkzMIQn+L
xhpPq1gWk+bnNL9uEJSnN3PYII1hyKQX129F9rJPQ5plHtMbu4CndVJKpMPcoNIo
vcNjjViNOIrPTJreuvUJ+ZTHmgyukNk73CMfTBsJBcpBY0ieDH+Wr/kgICyPmQ7u
GxoUUxoI6wqExsS4nsuuQ3CFv/Pb4TtKwTScg14kHai1KTh+B7xQ5b675HGk1mZ/
0LJUzq4FULd9X1Lejz6zaZJh2LMVKQSwg6XWofWZu/SyJDHmCmOQhMpRq0RMAfo+
Akg9l0GJbvqXRZlaFgSo8q533n2WZhLh++4Q+5Co5tE0Au0TGf2BMcC9bHB4csUX
1MOxCkmZzGocfgeQCTxweApNXBWZ+tVE9aldQhR8HGyTRyTOclaUj94m0UuB9ngN
vFn4Z7IDwBFfEEv5oouKUUgITIa4w+4KwHayIHpGIR7sd2qJjJ76sDBlnl+71ydG
XmSLfxTxnEDlgFh5tWtPePV5ueznHvfGWYxQKfa9rcgaUt84yC9h3Hk4un7qolUm
Ksu8WvevUwCbKa5PpvziIP+nIMBZ+6HRV2gkkUQOMg4lI+L694BXApDWHMlHYgHU
S2Fi6pxvA8E+KCF+bywOqQrdkDxL7SWocs6Gqutva7vAIqP4q6Cmi2VOLrvabN2b
NNGnn9xX0JSjsUlPR0+aXmDW/K0sVdc7kdM2zaXDJyHZM506mBs7VdR0y36d6byU
vf/0bAmpAVH/xQSgKmSqkF/4b6z93gtfzc8/8KbeUOW1WdTRyyNuqLYlwWpdQSAm
RapgLVyafnUISyZxTxOlOCNPKGl1PpDrupLdQwckTdgwBZke6ziPzafDlZ5oQYE3
MLZQZM6V/kes5ky6jqxVMqrIAIiBFFMyE3oQqgoOW14FaM4mBCf+o7QGPffaCRSA
g2pK6OPoLInkMjdVBNEODN5AoTg7bSX7AMBf0L+f6zJtI5PTabh6kSqAvEJ8e/+R
i0BkSFz3iBpLHqueAR4LDa5C2X1gf7KYxASSsG/5rdYtpIRsNzTc2VPTP3SXDYbx
zNZCjlG5ZOIjYKrq7TEBk474fs8TUFZFtX+pxyw3FIbdhk1jxpkPMLhm3oXL36de
eDFZCABbWWmEoEHSSOttj/5nTOU9CHNF5fvtT6W/8v1hL0HxvCY0wDnyUSPKX3xD
URTA1ZlHbSswXAVESRI2YLj6nCjynIYXXndI8rR8w6ccci5MQlpn50scaH1/eSbW
VnToZIvH0uMXOVni5EgpLJ5G0gSZG3fIMyb3rH81g7Vg5fRnlPGRRM8uhM8uGB76
ko7ZT1MfqyyjQfgkefW0+bYp9OKlUMkpbFXnEy5GaSoqMf/kxllnFpzoLRIXurBv
sFIru2vI2UgmRYZ/BCvhPoSd0rU+2e8pO+IVeTfNVfSS4aF0vwiwGK44dPWDyjtq
epdKJlVz+zNo7N7PD1ScXih58spF2io7a23Eno13JY4194gS/+2fyzHi+0mGsLsv
jJaVMA0iyae5yWwhKQDOY0BQFLE0q0s0pAXZPdu9d0QRg5pTxleGAK2m4L/GagcW
fBw7c0e93x8rPbMc38Go9+E/hfZhpt4Ssqv5fArHm0FeS+uGukAVRdciIKZ+bZAH
ZoSnOUFGzmTSaxCDuIvdDizto2uL10GjbSMlmhtbyui4QXdLqkwceALvsrthaEJx
hL03qKMzwxB3uCEg5seX63VaIXybPQBTuLQgtQPG/03sDcfwPMYRwMkODSn8n4k5
w7mTb4qkQQPrm5oVSUi7/s289MHX2a721FFM2WtTMlExHWxqN9PRAI0WenjW7IFq
5/hOPDNtp1fiDSEnDRbo0Mgx7Riwjok0t/FuTOsPZGPDZJqP04Qs+arwL+b97e6r
inmP4c6OcsI9GIYCf1nHcy3qiLrfAY+wThXdbdILQEIHp+9pyNfZHkJOLzuDyhxQ
y70gLQI+5XZBkiVRuu84+GI20yxHq7T8VvfnQ7Rd1rtH+dd/5GX9JcZ4AXzWaMz7
8+laO3GhtkhEOC3W4+g4VWnECXe6tMQXNo3nFUG5uevm0VEi9xnvcmQt8ZOagj7v
fu0ELXf+0bh2LxFXynlAEfhkSicSjCfpjUyJKYuoPzUEDv0TMplwnPMXuYhU5jcJ
ZPNRWOyVgj/cxPw544uRv87g6B67Lo1FjRUAt7v4c3GBuxRBzdyIMxpNFSHOJubn
cbKWD9mLgCqdgp144j0QjlnQjFdAHf94CNHRi3KqQvg8Bre67ZETnVLbeCqmNQVR
UZfJ9x5/tq5bpCn2+Pz5bL0whCevlwTdn2vZTiuT5ILyokocbTw7T71WWnrumyxP
kuISHIqdujen/XLVLj48GlvdX0x5bUkpQeWAMZ7jFpXZuB32LC16HA/IUgAOkaFm
nB+0YapGYONJwX2Y1tysPFd+ewkT9zArL80+9tKJ3i45lz/JT9TUJe9K2r5qg4k3
VgJLDRYdvZeXj5q8QreXEPAoBvviuDq6TL4I+KobSJ86q8k0EDRjzbjH6Aoe2/zW
jD8lC4L3vU9lQlxg7IHyXJOwWziDuOKEx9D3DKhyj/NUGH4GN+erVt7zd3Fghh0+
tslKdZlXTP0recayVbX+gPaa1qctC7bXXsB3050hif9TtECV6qylbHAUcEWfqBTc
roJTryjyvcYBn7HEQXKSysyoYJdNnGshKmGqHAYbcuT7oPGF1IoU/5PS5qJL8XiN
Ir6NDqK6iMcYf76B8opf2qCHad8cc6Em3/3zZa4NZEjBbLf/gz3Z0ORuqSYO4h35
dgtDKCuvJRBlH5ZEXBwDpzsjO8UTucBTQ33pA/iXOSksLcxBKFUJZxeOB7KsA2+J
pmMOO/yHqIou8ev4qUTExl0C7PHueC2+qVdDG/I4ncHWyeLpBdysMq2g5YVSx2q+
tdPUwhkC4sjwKxAFVFZkLA677qCiNgjRGhZF0Tsm4scsPBDtTYE3udK3a7vYxtQj
rZy+XLdyKsaUoeHFNoCylOmrxDd/qIpSzIU3YgaMkvYBLpNnZ2ul85r9GHAH0Ag2
c6EtIQ35QCeBHrV5Xz0tLWVzKdlqUks0V3H3vNfzbuMwJf6o+Gzzcp9u2trnoKN7
u23ShZ9yPXCUTufPKx/W1aQQzjExPn0pZD5x0454j4OvSPSEeybIAQdyu6vlpcys
Iv+y4AFNsQSiSogxNpUkPuVvzxy+ciwbJyuPxvodttpFe1cFL8Xi6FLjfyctaAEZ
`protect END_PROTECTED
