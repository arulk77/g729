`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLEWKKAI3g2qF2m7lrfi8UkTE76Bx3gr/ytjVZEw5qSA
d8SRX8F/NHNYmXNk/dTwzIvnraGE2QKka2Dl0rfHY/MqnSHrGJDQVuo4IiXT3pgO
+6IqV7RmWgXwPjxWP6BgyprGGDL0lWT20l6ziU8onh+eY4hRHiIeVLoJ9HWiFeK3
+YmMc76EpJ9XDtMUsH9ZOmOojytqr+H5R9humhIdXtkyPf/FRVJ52glhFdPdNIs4
`protect END_PROTECTED
