`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48t32GWjk6KmtTOcFEQPHz/4T7RwaOAz5raDlwPXwuPH
LV1doSZ/zZfZCq+EXGy4ubfZak6H+CKyfwY40GiNJZ2N0KwbjmI3xKT23HBztJYc
3Ia2lQyjvsZ3QUnWg91dKGzv/o5eohAgo95LLFkaKH0TexyVsjksuFslH+JNXmTq
oX4MKlM3mfo8MWFXlpoqe3Ahrze6tNts51LRVaqyVMtzqOeegB5i1hCDGCB06+kO
I7ABmYGChdDP5un/lgjraj6qEBwk96qT8CMQwNviwp8dWn6LfsD7D5+WDqOyE/pq
//wPQ7tXjbzFyAdQH06+4A==
`protect END_PROTECTED
