`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46q3BRH3Mql5uG+tnS3JnOqEGgqBvxlHp9VTs1gwWDf/
zK/VddFC7KfuQ1UZXzJjJskioDXcRBFCwOBW159wdCYi9O2BsopWaC514NWNrMnu
OzvOQd0ZtaqSGrjfa3rmx7Z0WlyswWkFFc2nWinxpzq0otQpz/ei+vmIFSlvS7yK
DU7S/2xAqkX2Y4K/uQ+cNqaYy9ioNJ2U1V0EevB2KOgAGSFzNvOQt+PVOOjVC6dK
7IgZ1iZylL7LnwFmpg1TdWMk3Iyh7dSH+2r7Qvb+Lwpq1a78VxxcinpMP8JQ7p/c
+kRE4sc0vTyrfLCdW7fFdkntLZBxr/SCydAMpajHiZA+ynzwC4/C1vad65GSbVUK
STqMk0OJquWt9obJU7L00w==
`protect END_PROTECTED
