`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePJZCtUblY2w3hg7DK2NIsEvwOmSziYjdHXJpFTWcal3
k08fpMt4EiIWE81rtYREDOdCZP+0yWzUhZ6ZEbSRanF4HhtyHoz7oAuURRok7aqK
Mc5cNMiXIofJxcHFvTpbI3M+Av/isJdeBCy+MP8Z5LQOAv1mk3lbEC7GZaitJBlL
XaH3QR7IfrUTX/tubrPf9Q==
`protect END_PROTECTED
