`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
1LhUcWbiDdQOQQO6nINwgpIVNX/XNH7aIKnwjikt5Uq5Ld94WD9IFr+OtPU/4F7m
8dkPdUDHyYzkONiiFDFkqsqKErF62VOuj7VP8l+pE0NhxtSqNzVMfvlk+Bhpy2Qn
/qxNi8p7Sf50VeyYNJwSDU7nt01S0Ssj9kRLUsj8QvmYlQo3szdLtS9aAJUmN2lu
wppBwnrXM6TUdfbzWVzSL2qiMqL6L+cyjKnl9/DSfJ10YSbVRJYLBQI1a1Hodmsl
SFcwfoGxPcgFfxzRKs5yYAmLiGkSaF1FVFfE0TsRg47RAnbqdOlJlaDb4N/1bDqb
3hFki5UPwVJFujZWCo3Lw8AKvi7mdmX72mQHEIiKyvf+LDOHsWfgnvz/pxxbE6/H
Xg1kqjDr5K8crkdF5JtG2g==
`protect END_PROTECTED
