`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCMdQ55qLP6RvJIu+sZiO8Z3XXIQUTDpd4g2BPErsmd9
dYtw1GFWv5Th/8hDRU3cmFIyGZv+KMUkf3+bPKdTaxGJIK77bDv5uL7tPsC/5lHl
VM/oGiHqt+oF7aG0m1pRMFKhsa0/p+hFXNKI9DN794HWXYZz8rkOFAZsje1mY+qZ
m00jnqe0Wiv6tsQURPqlRQ==
`protect END_PROTECTED
