`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBiMqL+topeqdw6O0fJeTDL95sgi24gy6qyPGt6u80Aa
5Ec4sX6LWXmXc1dNcRumjm0LLdaQoChXV7BnsikYwrXg1uxXJQkyk/SuCK2TLOut
Yc6NpAbKmx2Ka8o0zDvD1X0LdLbjqZO//rvZIkdxAaUp5MRt0kl2h/v4qm2p3JIc
y6XyTsR5BJDJ+8ty581h3w==
`protect END_PROTECTED
