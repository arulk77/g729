`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLRsbpieP2lAPIx8On6vl5OyzYHpO9EyL54rx3zOeLz+
QZaaWnhPOA376I2zAfreh+pdbJjSmZL5eAWBm5dwk5HvINVx06N+BU93Tnc479vp
Eu26bcAVysTaLH38EbuUejYng5/5a2w8MbVLAnZmNm68HCQ3rcyzP3ZPwP3GbGS4
`protect END_PROTECTED
