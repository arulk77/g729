`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
7RWERbz/SCu29vx1yp3KRNzM7SS2Qdy4yKfitFEvNxctbekdKdohpHpBLNGLbqAD
HykwboekuW4RbqrYij4GvpFHAK/uqWAp9gOYXUsHIsztxejyjCZgypzHHSqtWjaO
/Ejpm9nlNq9vA8MS2haosw==
`protect END_PROTECTED
