`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIVBQKmYwX+Htb4g+OpZmKzsTe9wndqL/RR6hOT4cL7v
7DjXLVr3oYxSuGe5o3ry3lMTKDMgQHi0+N6xf3oRcYR4+gQNXI3JeaOuC/pHYfGr
XIZyynFUIyQveRNNQlvvOWU/Z7deVxZP8OMMZSuQLn18+7aeozilEUv6iVChXxJP
E81Mfd0Xc65CZqWC7UXQEg==
`protect END_PROTECTED
