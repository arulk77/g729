`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
5vjklJ+Q7+QLU0hoqrqG7rvxGY8f8EOKQoZ0qY16xldcELfcwOH5dlrMEBtOgEpt
v50LUhRa82F2rF7IgelX+4Irl0goSnDUZv47CDoHJKTc9AwDQXE6/zSPreH8SNuI
AhB0h5zI89+sGFuEE9jXez3Y6pjdov/r7aAUnPLalrawuKpFnK9lyjGGN2s0nLDD
WNp/lmNNJZm2x2fWa2fVqDcn2boBDQz5xtM68Oj75cIB77yaHnEtWYkr/SZo9qAt
tgJRzni3rFWWXFRwdVy3x3QFsFrkBUnUsmVZ5xZ8hRms8Wqg9QwDPhChfik7nHPS
cFfDBzqxvDF7J+Zyia0dh+wn4GET2E0WdDDyuuzY8OTVTokAGyTkQE1ZC1JdQXBw
`protect END_PROTECTED
