`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40gbpcV4NYpg4mqPJcTHGF2nr2M5Ww036BL9mzgJgNqP
2nj5y4GN+o6NhTpWjMCR1zjxu1+N/TY//ofEmr+5aC9wXByPqJ0nam8CJ4qajyM2
b7GS8zIYRGyoGRVm/FoKl8qF5XSIQa5aI2G0KPBlmpVNdEe8nDaCn5pm9lYaHihy
zymnvDHd9Y0u9Ez9ganans5JjKOke3yotR4aBZegylaslvcfraeiVa/qeQTr60sx
Mb5PFQvDUTlOv9bBAG/oA63siXNsTz4P7ltEaqIveUoaWFVH2rIFDcuv0A+1cfEN
8vBDnTyx5sd1yoqj/x+3sNDPAu1sLwyyUVpwqQ8LE1Vata8qfoBoW+yvEAo3pUMk
zz9SKAkC7dX4PFt2xkqk9w==
`protect END_PROTECTED
