`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wkRttPgdMT6s0m5RM/5cmslRqAXaFVI1m9ashE+e5EN
yEf1LAX8OZrfvFnbQySzlYV1b/HL6RORCFPP236anT+mMzcg27UwOo1AzXpkASlm
qcw8sdBz2jai7oEV5CJ+1Vwz7Btd20ymwtJ16FO+fT962IUZUZnG7GL9SVWV5yLG
7QR5ziU8cJLnXH4PwyuQgLCrX3DNJo7LYWlsyjR1klBdVE7t0ri/EWcfJmk/8g0U
tM9k/+asA/JlI+VyZUH1IgAa0ODY18jZxKTauZHS1eA+4kFBnaElTGDElK+nAGsj
kgSobJ1RKcXwXClM/X5DM9gpRs5ooGmDGWGzRUwP2Y2n/Y4mN4Ca9gStv61C40KA
5anEsF/a5jFoDqUMtdGYo+N4teUqap4POlYIOVYpU5nYq76mgcnfqVUhJgY0Y3zb
rqLk0d5wfH3ub/2QAPXDnyIRhfzazYuKsW6dzO2bFpkMSZ+ObHBKFklvFdL+n/1T
`protect END_PROTECTED
