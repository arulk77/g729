`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
dtQf5TruJyI4L8QJI2Frhv98GEsZqahn9xW0+Ffno5dcVwTMPoxlwOm+zYvm/vjA
JaUj8BaSgue9U/xEQxmltnTSb5AsPtJ2Dfhho23aAusnxBkUgtDro9+RXuZaRoF5
+4dhVj6/51r5zy6hbCaIVTDwbpXZoeB8EU24p1kQzoSjdks5gXPYtbWIG52Jwg6b
afybfKP9X099jiSNLdYGEMTK7BWLC0nBJjd2PN1iZMSIOap7ir6epGavpswUjzCj
r79HbIC+hcOrVOY0ttLJD5fhcD/gGoMDciea2w4pJapnKFBMCqUGX5tOQdjWK3Ml
BZXGg3OX6QV2bXx8K3G1/W3/VqSaNRClPDdfWUWEMx2mKCWeIP7SAL2UzzmhFKyx
RdlzU28zRuKSVL2bbF8wA6Y9rbjiefCadhFv8mhLTu8xn8IjvzuOqrE9vINLzDcR
TIr2xv5Nm9XUEnqgIfjL/RRosYgyhKh3Yq2+GoLc2Qcj7qwNbdc4NEo2R8Tjg0QY
2Ven/mROw1RiB6zl42l4y8vp/q9/Tfrx5eVUJA1a6j12roN/vrQ6TfGmTZRIWii4
MKe3HmbKsAVnDQstfe+QTg==
`protect END_PROTECTED
