`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAQyB1UjMq94xsEo1Hyxno8cbnmZMqxLyFAtyiEytkWA
o4D9FqLP7CmTOe+NPUFhkq9PfWPNMN4yRAt86W1nNmfYLoCPY1jWJmisf9wFLN7H
6kxLMeheV9IU6nybbWG5UQg9/VVnFvv6azG7nSimzW7VxXxeJAUKrHwapkKgt1pH
/NNB4rifFfBNqn5ckVvVE0S+OOhSO6CxoStoXrcaQYvVITN5f6Q0DOfSapPOYpTp
9vWNSfqTop8l+j0CFYaJwJuwaaJ2fG5VHtyWbhXDrUrHFNEVJg1naMFfN5KqAtOz
0YTTPxIylXQj2lhhU4PIGrQtMHa5fYXHAva3oyS50bpKZ/DFk4YF/PqMlQXbNiPf
nPcgfGeqf9ng4Ixiv1IiTEqVLVB5G/vU2wwSZ4PLWcgb7eO5dS0hyOTG2eFE+LuB
1w6ERP6YqGRI55ywu7aBSNaAnTOwl2fup0j2Tsks6byQd+ojloxT0thqKAansB1y
`protect END_PROTECTED
