`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
DE3/3Y/jRUXXd5MOQu9u7orLqxWuwUHk7ZFVzZiJdgkHRvxBfAKCb6v2dHRMd4La
7+Vw+HaV/DqG48XmF6+OUwatDLBySDRabLJzg/GS8YWghzl6jwPHNUEroo6LPsSB
M9knJe5c8vBu/JRkeErC7KGY8Kl/7T8oRfJEXsPGW4EjVXhyebtXxWNTC+4BXipC
WZUc4PE8hEBT/2gEeOMhUmva/oaP+hvIXi91GKI7qSLnsdt8j8cjmy9v/DcYzE3m
yy2DJLUA9yXczDX+IvkOZBNUMLYRaHDoUVmNd1SL7lr9kQa8ZDvh6RYaMiaViRtX
e4bUsKiam2GkIC3eMJeBAaqpv7VPqyH+xAaijQvYbyc=
`protect END_PROTECTED
