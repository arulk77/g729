`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN/8mDO6VSiT8g7q3GpYuayhyUGoJPPRT2A2yYrb6jwn
Bk8GnbORCA1R2ciD8Ol49SKI5NC5BSChKG1xNH0fDexXZE7iguq1MnOcQEhK+7sE
E/fsA5G7c6hF5xnT7M8JwO2PEdyjqK/Ml+WZTDXYmKTLQXtwL/5XLF6kn/VGLURs
mzM+U1Bal5DQ290f+fBEizk878Z6nfELAIkJd+IiIHX3ucfwwX4LBO3GVesCN1uD
woPY5fL91Zf/8MSpgYCqOA==
`protect END_PROTECTED
