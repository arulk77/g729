`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMbQslOMM79ImwqYnf4sxofrgMpITNiZA/6a5l7uOTrN
5Q1pT6YnRbo3HPQyiir6yqxWFotNMaw11HV5gJ9tOoNGZEUUfM1Ov99ws09ic9od
sGkC3bh3Uct/0cz8tGHF+ihdQJW0ANWX2nkm9HcTe8p4pS4yZJ2vI30BnPmhKjin
Z54UeBU4/8ZZ2gquGzd6EaAYGz3O+bKF4hVhKOF5NPUg6ExeRZb7lGyxxTAb6XC+
`protect END_PROTECTED
