`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41ObEIwbpeM3oqhOuRyfhIwwIpzN8ElYreFEkWBgLunA
tyBY33dCqkqmJ0Dg8iAkB9vv9k3BKYhCdtG95lWaPsbdTESKI6J+svy43kUjdhHs
mhMcqS9HidKuHZtw9lRBDIkduWm/0nrf2jU6QU0+x6HRO/8vVRT1JDv+MaqnDfVH
5bRQyBHptV1DWAXK6OeGvD/rQ8sFT5RgVlCX3ct4aoDyNjsBmDvfJb25ajkAlx4G
/osDHku3UlWe0D+Cx36dL7IpI5xRvitqIUdqkQW5/E8=
`protect END_PROTECTED
