`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD2bQKupNVYY6+QfFx4DHGHUZdSt/TYQD3rsQC3IJnbT
7J09gaiFp7wYrZLmXa9YEDyDeTuI95AGAI57w5YZpqBKhxVrV2ZMV3Vd3+hN/r3R
qh/iryUT1csdonCTjQmmP8oJ989Ze4mEmTbturbSbp0Z6ssRoa3so6buZqucubWw
tpgd2BxhhV4JbA+1ph3/oxSM1KyKE/K8gxUwxwiUWxbzqrf6ErHLUGowI87rAmoa
V8F9F8xhkyGQar4MeYe+wnhQ5QMChA7YwM0YTfGemLuj2hghZ+4624XySyfunNjE
X3B3jc+MpxK1siErtW2ocV8cKsluUIFRsXa3g4gDhTUvR0KzW+BPEEWucPLXfTXy
fGHxz6Gd9oIFp3KXtJ/LyaAJzn7/11AnrPIYrAsao++gKPtnWIyeR1Zuzgk1TDao
FlZlQExRUBQlGK/wsltD1+0258Qe6iLWCWuEd5sgDNNeKvlbrLhr/uGiwpzSfGzi
F6XPNVr72Mm2ux0xh25GJDW6ZKR+uciM5aNcoNAJLCBc6xHHKRSU1RDmpxCY2SGu
7TPcHFx+DxaAJHtanRTJ0w==
`protect END_PROTECTED
