`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMT04WXoaEHXgTiQo8mD/aemTWrirVg1/a0wCnJxDLvJ
kMkWcWVWEsTjGYXP3ZGaqSYPLryUz9rsQu2KTqk7kjUHMMYISSJl/k+gRCOKBxNY
N/NUQU9ukJOdvfVw/TCfV/dTqwZHkptHDxIayvka13pbC2IhY0Ft2HH7P8avCqrh
E+urr+WcNSxU4bQuUlUgZRq4ALzE/eSmeRajC25prtxaJIkXIGILexbuX0QP2t1Z
dtQZol80NUl6vA+TpnZl7uqfMNw1iu7946awHPX2maU1WZkmKIcQqi8712dcjQ6N
WLja99UY2Hvx46RSlZCNmLjLCnITVuKlri0h2nQ1nR8VDZPCo/XkDgw89gveAbCc
dBYDQ5EgBxc43iofSZtC+jsJnqBxUVg30BrBi27ehthiACNDaTLTlAaSvTPx4l/h
7xK1/DcqiIodR7W3O0kq8v0Ph/SauTcN/ZBpyb4nuga6Hl5G5euUHkicgRFY4vRi
+cmeR8Tj3Ak2sP/wC4Ygw4fEzq1IBoq67BWfrw20wMEo0TPsMzkwU1JfRZLR8knG
Cj52fwtNGPjyJLFXB1HwuvESPrQlyxZqedRM5bNC60yx5N7Fx0iH3nBOhOc5jEVl
`protect END_PROTECTED
