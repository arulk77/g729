`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveE4ThWfo+wtzV2a1rOUZqvVFCZZOXhZ470x1cC0M/C7L
u55+QbET5CCoiM/Kg/7w6PVOSqPrzE2E6257rNpLDW6BKhaFKXkrApnjWzOAVHrh
2FdvtkqIks5247Ko/Lo6uc9HbhE27Tltsqbe9ZjbjKyoxcO8Fjs13nYXA3KLuYwN
vwRgfb22QxClnp5Ji+I1Z/TQhGUL6Czi2BJQphYHtwYy5040/WnsWwWjsV9G2FKX
zem+mSg8unTsCbSwfh1Tmg8oHqvzwmJq0Z2ZA4A7Drw=
`protect END_PROTECTED
