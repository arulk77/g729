`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zMMWcW7E6L0kWAB/Pwb5NP5lgxcKb1BXQMd3+pS3Ma7
gbu57c62e1QWgxFOR9IlDlVProoK6X6wmIz3mmQhAlHdKZIBnkyTzU7zN0Qgubt4
0ylQ/YiHBfTq350fFynkT5U8V8tc5++DRwZp7VfeY6UYOtHZ8t5nNzAVPTQ4qFmC
1vVF0iVC5fk8AayTZPpXOTF2HhmEyhNoPm1de8KYjuetlCKWhCbiTEPcnNlfDRPA
kDmuyuH2A2DyZtrAcjJsOZHISFhV3/e7lRjltmeUACM=
`protect END_PROTECTED
