`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45jTvzaWMZbaBATuMgBmGs0W5mADR1sKggXhB7vmsXFP
zdZLRq1du//Nmdp5SljXyrw0gJN8O0PNy3Kde9wc/I+4Kvrz84r2As6L8W1Tv2hJ
QAR9QNV3KtX6S2Gjf+PMsZ7+OBRhxNCkzNCpsEPVLFyhpPT644KowO7MHxCj6BES
4ijsPXfjdpms2dWns19qSGq0+YCTpHmKGWanjno2hgb3bzcOT/B2dXh+GnCcRPaj
RUFrXxcObyjxKDebqoRnIDuaR6Yz3NCftC4smnzb6KI=
`protect END_PROTECTED
