`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAelr/radkaGkidrfusp+iDfR32wjH28vqG8rJVJwbK+
LhmrF6R4thPb0Qt8n92UQG91DhD0ykmOH1sA69UraoUVv1Go9EMAjyef/ZAKlfJ4
ysoweWHMXN92923ujfjdk5w9WIqH+DgvT2eSZpo3YBBw1yHsI9IsmcTcVZP67TNL
uz8FRdq8h/9BjT3NQPKXNFrKSQ4wTUwWgz29F4snlphoTUzETerdDuylA4kWm2c4
`protect END_PROTECTED
