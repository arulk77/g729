`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEeV7oa+Q0xp3bH+Z0AK+vwSksaJQZYBatHRtIXg7Cr3
sJczbvadcvpImfCBVeMU/JNXBc8OlNseXh391XBCFRRc2IPnNLKJrBf+LAVmiivR
XKkeh/kJHmCrSkHlbqSZ5A==
`protect END_PROTECTED
