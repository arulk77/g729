`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
euNHD1H/9nsKTUYP+RIu4jX89FmmlqhloKywIoG8/vqI0GZP/ZftfbHw6dy21cdu
ue6RtDl3QEPFOWzwU1qaTJ4asOPhQj5q/47KSvVVbmonbddIvVcSVR18saegQ5He
sKgHKTlBgXW+DUSvdcYyGxl24ai2qptZgPAlC2FUXPWwDphDgKHxuJQXyeeOQtUU
z4LEhxkEPHbojYDOgbQGtEed7wRzXYkNn3c05G5fgX1WZiAQDnc9yiUyXr8vDMNN
5kAG7G223KHD8qT7GWnPU2FroxHHInZdf5cCgvV+2fc/gRLNuNiR/2u+5zCBO6ld
wTaZnIRqgBn4brX1FpOup8tyVvVAdFvjQFRls3sw3u0/V5sQeQcT8wo7yJc9Vhak
/RjjWLIMk1E2IdL9ebSnabYE+KueE6fFwR4bWW8wDYmozlio5+FCzMTq6NLULX44
IZ4OoJb2arxlLUziaA1UDr6VRq4hkKFvCYpGiwE8sltN1rDN2s6X42rBIsay0Ems
6OZyVXOsBNIBo7KQUjqopsb5HVm8Y8ccewDxgQZ0J5CRUeZU0F900XAQ9nZBDk8R
tmFpa60dz2EFZOr9WNKKsjw8CfFiYwfK3hVUQBCcmtHbZG7dVDbTqYi1jCSzLuUR
TU8sN68WkMKA1JFw0W8ZnUnnM1qb7fsOrp+4lVa6cnJVFSOiaC8l+sw4Kt2M44Gk
14cs8DiQ0UAvl3JGNai2kAZXYKPHNEwQHIN3AAv/ysl+2UsadcEnH2AjLt1ptZSM
g4hGm6ltab6sc8zl2jXKrg==
`protect END_PROTECTED
