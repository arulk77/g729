`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pnyY3jxGyCgnwWklYcFi/a26A4ZXSxGQoXA0HeDiTLKxyoXrWBIv0gIUkQo0ReDO
H+VrMyxBi1f/FilmN/FI3iSfOSIfXwg3znZCW2qpyQzYhrDo/dE5llkjILgp+cnF
UA632L9blZNjgnckhcrMfEmcnyplArrK/L8jpfCk4nAZk9jhFBV5BRuAch5ocKk7
1xbyAGBsXARh6BJipvGr5z8NrM7tqd5ly1/WN5iWpLSJ0ccL5Ivhl+/ZK7wi7BP/
HkWItvbEWu2yLgX3wRWmZGNhDbHVKg/2WlYH3oKHgVH43V5/5JFOI+GmP8i6ftir
zQKUQ4CSQjYwkMg9u0CLwgpfefqzRjrSQAuIafId2gQgxxprjHm3Y2Kvf19zvYXm
`protect END_PROTECTED
