`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C8In3impixYou9IBQRQuyeWZLnR7FISS20fzqvSR7AKs
Ga6GjuWR16ajE8b0c//oEOyGE0EE+BumxmC9YjIBGMQLKsOFmrqxkJQy2W+ftY52
o5kix+DMlJmVfuokXPtkJUGzCoHHcuH2GmSRQvcHRjaC6Pk2MiwucEuEaxCq88Ay
34RlZuKnocs50BeVgxMeDbkvy8BVfD0Pj72sRZoJySgdO/7Shd1hAUH524wXo4JB
CizBtvm7v1wFZQu0k93z3OLPPfv+cLGY1KXtuDQARewTbz5/KjLekQKBevtaRkqz
hhclu1v1v9XJtm1NY+4BIwX+sVHOn2iQCpGVr7C1aSyd8uUcDbBvzdn+J5uWCgzV
3osbVCQTLq98rs37x8si1Nwg/bP0CIAjmFoyW2PVq7183asoOWMMkMd8oGYbcH7i
9aFNtoI5jFp7U8eRFrnKuyCh40n23WLhTpVtTC2n30U=
`protect END_PROTECTED
