`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
9w8B5h88nQMyf6YzAT+Nyl9BrQOPaY4GSiPVW/JP7wbltTY5dp80qNiZ7biDFqdr
48VU+O2AGhiFmgSYuokQt/5xHaKoUBB81Xgt+n08u0BCbR13sQWXP/Fv+4IFkG0q
GG8K0/wedMAn8ktntGQz9Rve+sqkHEwPtz2iNGBnjr4efpL+l3TLMM6rdDptgzMi
VSkDYwTVpQJBkPgT2nUvuXTYCFjYUPeLNN6uVjhLn3FQOgksnYykXRGxJGEahNlu
hjeDtt6hzbEg9/iROeem5bhph15LpkyB7mSctFOCt0ng2UhMyR40dGCxDfu7EyQc
WfepXuq+7jWXAECaKdCmAKhoVsTCijhmW98Wx3sX8u4=
`protect END_PROTECTED
