`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JiTcIp73gERtq2tKmKSArqJM2anUpMmJ6Mpm5ZSQYwutCAEMRww28McpS2Rmw3om
FA15qVDS8LaniDAhEiVS7hn5i5g0XdAfmDIMolDlKiRoWDzUB5b35co6FpheaYFh
nfQC1k4NYzAEaXE130EPKyeH9RizC1yjSBXqgEigw9dgLLF7fJtcAnNifIImJr3d
pAYclY1RQf9bQhGq0fwt9GemNzAaNSzqdwdyLVXdUvagC0YJM4bkDNTs4nXr7bkK
yKI59EeugK4YDoJMxHL5epIVkA6IoirJuD1PJfnPo25zhalUKDZa1l/oL1u/GlC6
lSGL/LldJEwbvxtBW3JIbkzV0Z3Li8dQI3fE4RLrBuU=
`protect END_PROTECTED
