`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGj6OKy4+jzjkigHFbtSr8Oo2ubuySBlVicsnwSVrc/G
g/9A/7yfFRz5I6ggfvzr0P9ZZUlAjYCnso9IZzJGuL3egWTgwumz2nCUxkRncEeG
r7Vzlvo67EUy452ET7XEBE1DiVNBUQJqokfOi5XCZ11h2U02x7YIZUToAA/OekA4
Cma2Uu5Dh7kDX+aLWSyiU3JSaUeS6jf1MFEY9ztxKRe6zba9pUw+qbHQUxB8o7OI
qFtRQfrNiGzLpwSKM5wXYr1pcdgB6JPpEtB0yOX9ecdUURVcIzr0dFO/o9XAkz6W
J6dUTE6sUqxbuYsDQ4zoGtXVkqVeFNAEH7jaOpJtTMsbEddOTvqpLh0Xhx7h5dyo
U7xBS/vaeh+uVYPJTCapNFgN5uahNk9/RoknyGxEMv96n3bQlzuFjZn5UuYxJY0z
9Qm3rUBf/f6XYyJT/6nP/LXvgb4VhK96Ta6PpdkQcPR7NfTDV/F6XMzialTb7WAR
SaZCsfpqzhyuM38jPhb+U/kZwLdpGuBBdH2W6C3FwPsB2cp5mbxpFsZg/e+XLWmc
eoixLV1FsCLq0DJh2fLt5o13N60hkkU8a0wo1xT83BY92Pkl4bHxVD7/yG28rGcL
6fq7US55ajDdDPYTl4wUC6nR8aSGUsDLhr1jMIyhB+XX1HQv3oswCpR7ZWuj4VKE
1B/Wb8rYB+JabO4wzXuhQbUvrKYCz2iGLgQPj5AwVlIN6e6wGm5gPXNX915yIQH2
g2C3sxilT/3RYObAsgMshAqdyLtE/IAQaBh9PNND57Cbr+M9ZZOB6jxAnvMAu/Su
rcxMuJGE2FdR/eaZHHbXsC9oUQWKWiXYkC8QWPNkxog=
`protect END_PROTECTED
