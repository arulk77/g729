`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
76sFkWaWtW2g4TUTKwVVqtFpU7DGuuDG8WZtg7tp9MEQz/4bdtGcG3VcqMQYL0rx
5P4QuXQsja8NTQTOF7OLvCbHr8+JDZMufskSBQlzTIM24C4xpJPOywznGluDHYf0
GhwRmmBuBO5RvGnE/vqZ53QetWOJ4pg/1r6zVIyToBHHFvKuVQBr3ZJVz2L38kO+
8S4xTF7opbsreFlM0eads9slRcI0ArwYARR4CzWHgCyqJOVDRB0K7GmLqXrC+WiZ
2yP/yb5KFOk9zWoK/5D0jjJckwAnd6brZAtkkK9Bzy7hBAWMO1gPS2F95PCmMrbk
3gT3Lj0HBFHHKEaqoAROYXJegNVihsoIVjN7TcZRNzHtfJ+/Yrra1QsFXu6nE437
liQPMJNHaHPCP6js1mIHPT2qZWJ8WAmQIEhTeKcN13I=
`protect END_PROTECTED
