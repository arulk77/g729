`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xA9vEj7lLWUsddqaGuhsXJ3VrOovHlCOT0rtvukTKq1
t3mh3IhSAL4ah9J6NHYFuMjmdXxD0mbOyI5Jt/OWOY2tvbLgQFDPEDWoqflf5a+E
zXf7FMe5uN2O3RRZ08csMmXcNG45VcjhYtUOXLS6Ll2nIY4z8Rs061u3pnbr3czV
21ynwi/gD/bTLES1+j6areInst7b5S7F44bND+nrF6DX547OrBUjTUJmXteXjRv1
9ZVZZDkp0HgrCsDKZ4XjzjH8T8ypBC3+UxoS0eYhnpdg1R6BiTRs0UErumGaPI34
18qH5boBEHSh2+ATW0GpSX/wZZZXDaFM2dju+2ozCHxG5IO04hoYKBrSc6C+xLJb
L+rSBv67aqj5pqjpX6ar6g==
`protect END_PROTECTED
