`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
sINtcoOXKI1doRcaqc8fkZ5Fa+vYLPOlvq9oEJQuzmFEoQgqVIfWKGboYy6R29VV
l/Ht4BkrhJU8cm3Mk2Aofe5FeH37fOFJ263dgepN1103OSNvOJkG1d9WIy82ZhOQ
8sOfWk9eTnJdvpr6Pk+gZMyPvNZ5ucNXTWbwoNc8zKeulWjrDN7M9mWwH2wzsUF2
LJ6pzm8fpHgto88B66m+gU5GwC586nhX6Xfsx3P8fJZM+Gp9/xgsY0f9SVM6GC5V
Nbeu2ealodq9LjPJ/nu5oOTfHsyEHy8ey+P9uje7VjbPzQImDmDdUwhMLU0EunYC
TgIIo+Bvduo6/7ukUhhykWxOEwQSLcAT1QnUhMxMUrxbtyDhBjcEwN153eDl229I
/aIVBuQGyIInYe4hRzg6y9O16/STejCP25aaBi/5x44dTS3kU79THb5CJRl4huHx
3qIjsaEEQOcxA4NLUBQJM8wf6haaHZ4pbgHf0Kmxuc207Mf537K/52yDxitk0PQU
B16ZwLAS0eBZ6m1GL5fkqxZ0V9w9nyeDJ5vW3ReGBddW0geFth8qitK5ve8ZGbat
RolSvSQsyQineck2OCDvLA==
`protect END_PROTECTED
