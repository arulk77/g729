`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47QaYO939KOTdbSnILlz3DT5ruHSn0Hoi13S2PrJYTj1
RpXTC/dT8C37+DueGCCyNZFj8xUKm7MkcPoAq//HMkxJgM3ddWBXW9c3w6LdyofB
Fbqs1niPA274mxEVZ58JZg3r3UZhsmpuux3ZcX80/k3haRtD7Tngj3HJFT3hS1cl
d+0HjBryVGyVXp3x5yZzmXJ8M8s65vj092R5RjhV/T1zs5AuaAjbuvhObHlgf/Ok
RTXHwR7D08kgkwJl3onxk7EapXvebtzrres53bgImetX/eAFwdM6is19n59HbZKn
1OyhoKo28lAEuaQWfsUqai/uqcqZ4SEBhNw4K7C623i+OVNBJAQEymZEPcVui6io
1jzUctLX8ysXJIb+z0NnOQ==
`protect END_PROTECTED
