`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJcdmU36WX4Rb2Rk7bua6omuKfQJkH2Kj9961Gkg1+C3
tSBauaMxz5ad0ws0suw6FhYB7ehXS43K78T6ClDJRqUKQowWJ/vtB3HVdrd3rXUQ
qFPTNw0zkHJ8lpYA0AXipWBZ4GBxSQ7DvaQMNceGWnrwmho6bQPmjNTnQt6wjuNC
`protect END_PROTECTED
