`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43Q6QN1DEPoze2DBTCSDYaxek9ODmfT8hJBsMTCuJjmE
RQr9ygoMNvA4UrdYq3O5Xp+JjM3gDvpiP/2xqEspLJWLcxDQTCYoy2sf7ZrWbmu9
Mr11HCG1jGnJJNWPvNLXAEwWdUj1Qw6+nHuVxaKoUuiIBPUWoVXy9uUejJwTEO5+
AUw14zEwf7HLG8IH3icxJOnHgM+XWeVZw7P9k0e2E6rvNUAXXdBfnIJTr0nk+Kb8
9YcIrhCB92AW/hXpZre/r+BfDnwc88vixNur+uyltMHV1nbNEdbZJRrVjutSPlfg
O08moPv7h2tockhx9bIMWvoU+NO8rXycpmR6HbRLcmLu2hxz7aJ+evPl0RmX2ZDB
AyxELX5heuMst5bAa82EUQ==
`protect END_PROTECTED
