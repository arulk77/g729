`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+DUEHLgxA1NQqxaCh78JQjGA/Rd1jM/1hOvL0zf7T16
JpxKEcrXd/f7QZML0gJclTruxiVtpGxQHIK8aCc4PQmEPZIxrVBsq5Kv6l8vu/5D
WaaHePjcwN+2BYBrN4Lkz7LyCqbfYi/rwUx+6NafdififYujKSk3ejW9oj0jN0iZ
JNWNApSUQRsuVtvBZhQKIWV8DB46g1rLt2qWX8m/ebeynuxY0Z1BTH04650SNvVE
PiozxkBvkk8fz0ffqKlpTbdUrNsKWS4ovNdOztcAZmq44IC41EsC/1M9h19uK3ru
nKa85fa1ixf8FzEx0nSU+8qGEYWACIw5AI1we+VA0mwWqD26YPnBhteW02L82Rds
MDMrOx8TEO8JIRakGUPCRQ==
`protect END_PROTECTED
