`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG4TFQDpQ6BVGIHYnoT1mzcnbxSNgy6mNHUaO4Ljv28Q
T0i6o5mwjMxvrJgPBLH8fBFvwYSq0r5dNfmyYAdNUgSzWRucJSxiHFpZfKL/X9rT
fgCDLmdM5ROa7/omUlJXxk4iJ3bEuPVLwWSO1CL+66Z8FwElmCBV0ilzPI2vMqsK
0cNkWsVWyZsXcaHz0qN3r8HsbhF4Ns1OQGWxLObXvfphsCvP/siao4mvMMCZ8PJq
K02A3nyXym9+hHAshMMMB1q/vHQcrw4CCxfR7di1LxcUg1BDejPlZfHJ9ADvuFwC
NKuq1GGmpw4YGMX6OoNcid+p7/tvQr8rrNKk94MEla/ZbKwvQGJjTKfqNcRZ6uk8
5I4v+3uAPUKzdtabnbRu4B7BnwzLzFzByM6uUpPGYTnSceYOAjWBwj9gdEe0lCje
gXjegYC3Nwjqrc50l8pCuCAPgeuBM1d6J5R8aIMqkI1ekQ6kd+dRYg3ooZ+tsB1q
vuLpSpCo7ZXxztdpB9JIxPim6LWcjbB9BWRpV4JXP2dvMydz/kIOIuEonlnmmIAY
`protect END_PROTECTED
