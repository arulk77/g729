`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCvyRjdHCVw3zs2dRaYMc5LgQ3zQYWCXv/7ra1WOO3Aa
6bKVFIgmTYOvU/W7r9J9zdK8QfMPXVND3cxGOe86xGiTSJE4IaOQBpUNgdhpWwzZ
rJzzP83Gy+o4bpg50HEmZcjxyL9AYf/8uzhlW3/TwqXiBR5WyLbk4f6qzCIFKRWd
kvSvyfrplYNCfeqyEkp7SniARrUxRMCgcjhd3N36+VduhHkDKTKKYEp4XDQYikxv
`protect END_PROTECTED
