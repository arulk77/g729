`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGkt6ZbGRjuO8TDFhTC/Lb2X8CKndTlhE0KdOQ9D3hty
13wPJBc4epzZ3Ae+131sTXz/Ut0xdedFdNqnbh4yeWYRqFBbX6S+LKMiBwIJZjxC
xAENvNYMfkUyFk4FfNb53IPlN0MP36Xrgfwmy66gKTfU7QTLpVlmnOGcLcREaS5O
aq1z4h6tDSgDbqvA1LBsgMJY96CbCG0I0FTa+FdiqIaMHYKwAvyQExyF7+eDwoCu
`protect END_PROTECTED
