`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHTVoEYkcFGVAo3tw9u1wGwCPFq537mEkeaDeR+Y1Uy7
aBU6GxjTWd4b0oPewbWWU7folYHxuhXKLRv4FmlTaIoYjDTNWu9eS1sLvu5Vje85
XzDlEW2Xb4n3mDWegIh5Vykp5VScrqmyQl7zRse+aff8NjmZGy6lGooyowSrTUkc
QbNkAZKsoTD9Wfa59aObBHlOUIgOpfbZ+Up/mZS5OtG8SGnoUHyuLp63iXmwzSXO
`protect END_PROTECTED
