`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44aFqfLTuHXxySg52qgqIrZTTu7EatjDws2IUp8jTk30
4hSjvmQhXAlQFGx5k4sUN5Yu4gdHCLeVyDEV0r5IsyrQ9YLImX10JvOenHvY1Y0O
+9K2KWo4WAXH/BLfwpqRHjccJTERT64QHmgHHPRsoUcP3J6diEwIbFzvHQH38qSu
FRds7Tfuxqxta2Q23IVfUwBaGNq22YQqUeOFQEe141KDruBItXH9DUuTMcROHYls
rtd/TIzxsarymNJ526gvS9g4M3BbFyiF1l95krV+cyrdb3VKM4TrXsCqxU0TjHZ4
9JVlbvyYOerS5fzj+bDkdg==
`protect END_PROTECTED
