`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMdpIqPY/FmPFNjDvT6KebiYBprRPYFVfsNMEXK6BPnh
tPHy92VR8PHCzN7zdOuvPeo7giG1etQXQxmAKPzd6iMteyl5yGPJM3whhHW6gWIb
b7SkTtpX3GtmUF8nrYKoE+KuIH/+hQE2Ut89KhC1hhWA/WEQoHmWQ4sjZ3OvrZg5
9iDsrhqq6vU34HvgvMnQ4w==
`protect END_PROTECTED
