`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wEyKgxYm7/yAObfGaTVQfCmXkP8nzBej4YUFECwxn4X
5pu31ntG+HWHxJiHdI2SS8arQd4O/Sd06gLulIU5r+kN1yLc3uxXNw5i/OWlXT/z
2vBs/jgDroHUTh0G/JUUvWPV/ie5raoynZKhG9ULfUcLvkpnjjHjqB7vrKa4YY4g
/aSrVnkqE/AI5HPllXMSfivDrQ3n8AYWJiVwgvawXfPkGVjowFQpaaslg9QQb7tV
eNoJmfgPanWGp8jBbBr6j5Xm5PLB+fPDHPw/IjVJyEI=
`protect END_PROTECTED
