`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMsbwSAbQFsITXRaGGhqN0CpB39rQxnlhNDdgAJQsioG
bw4497g39IOz1U8Wz3kNCPs+J0JEF3MVz+np3wwsraoSU5KXS5u6NuRWhB0cEsUQ
lX59v7LKvS/YiKgDEKrPmzSVhEB3pgzAlnMk2uIwhwpILRDke3bpnMsV+aXFVFM8
m5z87BLE7QLrfw7rNGYqhSGsPTRiiYJazXDfjVc58pbbUkOQeNm+B9TVNz5FE0bt
`protect END_PROTECTED
