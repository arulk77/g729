`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePgfb992i1ZtLexIAJCXmKU3eyKdaYpFtsH151Wb3teG
ooRYrCr5GELDtoYq7DHt/yHVOhHyjVJGeNANAwgcA0tpEKBxCcoayxmzPHiXYzTc
8oBWThD5rvPlDRC1kiDncPru2ZiHkwL7cTI8mE4SUdZn5qhXTSYBdkrfdWS3NpyT
E7KrkZNqZSYPkk4AQyS2xh9udtVtwTCghp2Im1iFFnx5TThhUSDFGHNBVEna898W
`protect END_PROTECTED
