`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42OZKUry+AuctpZlwExooZy9/ty6pwKweqf8l1Q8lTZQ
H4SMlkWx3wltr4J257ycBkBOVNQfjG0ykS1i5IzPRl6lpMSehCYZn47cO273O0og
kVMOtgNQmR/jG8JjzgN6Kx3SuF6liR6jdEizfDDBH7gaB8LI1RAoQngSjJrw1V+f
wlI8Bdz8AQ5yX8FehkHBiykCrjMwdnREo3k9vedGamI7UpQ/GlL3KPZGE7zdNzZI
dxBG4AXda0So2rMrj5zb316doi3bxvHkNL0x2JuONGo9Z07aqyv2j7iJQww6mv1P
K6rLz/yN/igExyskNhBVPKlkbB8IsY0LRKRDLQZbK4zd3Ny9zwGZD/IVX8Joc0wK
q3f1+AIXrvS2kq9E0fU64w==
`protect END_PROTECTED
