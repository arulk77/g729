`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAHIPuO25N0wLfwYKSqZ/V5qNT7gxfq32jVeFRMlEVt/
GcnVjdnC1VDT1Wqlj4nE2QNy2AwFS73Sr9Oy/kQsdKMqh91yzin+1tAob/ToU5CR
LZ6fRndWrgbykyJRdLBMztxHJea1jD5zf77JYACuOdooEfodLfTPUZ5KltFQznIJ
A0EaR8g9v/oEH/ANlSKkHiYhxeWfXNsyiNWEZWZ0S44ijlUn5SIJEcTT0oPY7wyr
`protect END_PROTECTED
