`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJkUMJYFr8wwOoY6Vf3LyiaroisNgGxcgoEIaMnXmxUv
rzK0pmQeuolrQnhJE9Y8/uBS/+Bd02ARo0809DUamqEM0gcSuUfiusO7BLiKZUrq
cyG3WHuB+wzv5eSxcwp01kUyDX+j7mO7lqfUABddzKGMA4zOaAGbkEUlw4sDu3ME
7D9HcS6rYJU1sg8teu5kIWBRHzXBZ4Gj0NdHMKp/3zRigiN+YfmIIFS57pzvnD5X
MwvXYPtkyQcWa/SbHdf4MhP3wUJJZGxEMri2pX/8hLhkSmm7H0wVJZzKzRQFGemo
C6ZJvt8/77MwU9h5JPMkBbR/L4qPz5Stmr6c1dLhSxzRXjPKgXSGlPkRgG53DIb0
6HG6+LCXuTdDN+tChHz8E9pGVeZxTiFBmE5nsV+J2JBQjq3JqhWAECEJGwr8HwfU
ANsEG7J4bvmUML+RVAkGF6h07mAUgIN0a00Y31HWXEGGBzfX8eGENurrKbJ61PpT
vYJCvpbUQrE90khUKBwCXI8mKt8AFph1lA98Sc+r6k3Sbxbt/jHR9ssb8WUsMnhz
UYQKwZmWM+R+wAp3PaiMtdYynPXZtFG916ReRvqHHOK0efJLwEIuwHGmb+s1iwaX
ChvrlrwKXl08XtQXyZU1lpMNS1yWADBb9aNkovUxudBIygpUBAIYWzDNWUPUkXaC
`protect END_PROTECTED
