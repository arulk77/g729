`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePZEf8wNxy4Xm52gPP+bH+SWL+b6T0FaL7TGKlj4Smg7
mbO3YxJgMB8nHeQo0A4nf9M97/LOGkZl6ByzYLPEU7Og4jqpqIsFQ+I2wKNutCHF
4gBep1Edzl82wRE3AwP9Wt9wRaFrpDQIA5Gy2xkCUK92hN/Ao5EkeK18mbqnHsrM
u5SuuqxARpWEQlRYbvPbuEGJqtSSbaQGANUrzl5plxJO8kItETgBCSIt9rM00S+U
xPvsGlFkBum/0MdkhSO9Mgbi0nPHh6n/zHJEFcf6X2TE9sXLKQ5lcBZ5XvJ6mcUU
05xFh70FHvtrKYg9vCUiM+VisUmpX0alXcrKLrvTtxuzG6XGwPklmMk0DkkMP33z
8H4CMh/33zMI8fmLSJrMWtOSh4RUZ+fmTlrUQbpXvxNWjpJLVDpl2gPEq79lgpJR
jlO9gLZYw1Dyk7QGzhWBDkp+/4Uq45CnuA3CuNNMj14UnCadDx4k0ox7dsSA6auU
JrJVcc/AAlB1Az938FjalYqALBYmuk32cXgXkhUiy+bB9NBaecq+x7HpoMQF2sgK
V52xnKUD4ft9ORCWDLy4rSTqtOfZX6uH0F2zzKt7XGU=
`protect END_PROTECTED
