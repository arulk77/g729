`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
dgOihEsGEmPjt66fikZMNpjrxVzwO//UjZX40zwlPkjSerzHzYSgMcW4lQOPuCTI
2sFbz+p1eGiBlVHOPo0mPzhcJtV6QswhTCpBGAmviVcRo5GZGG8xl82j6cmv35vX
36TISHsWBEQ5Gcu0xkeNCZfJsnM4iJbW/nLm3xJyNTxCrGJgh4mELhdfvoiwCvDE
y6wVZJ9D8+3ngZD8A8zmBpj+T/aTfsR5EOgAMn5PgkI1mxXSx1SomqyoXGiAk4Z6
eGRer2j0wjSHWMQfWlzs2y9L2pLXiAEHYkkEwLPbD3/voSC3m8l+LnMye+zQ16TZ
i6Sv0E3MAV5uXwfgbd1mNe+zB/5ZvoiwcLo6in2jARk=
`protect END_PROTECTED
