`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHv9FXmoS2agsrl0LXAPuHDl3eYBEgaZMHjMy2yDkbLu
Ab855K6BtdVC9ArNBggEGGX6sXFCwo95o5vG2TLnIWldVA4gppx89fiO6pX4o5qv
ea4PLItcFyKJtE80NvmsM4gpNdy2hcQ+tGqrbLjrkkS33JkBGRG1mXD0Bq0CpS5R
pPFqNE07UWwABBijTgaya2wqFE3fSdgE12rxz6V2iXg349O+Hkq5iW5Bn1TGY5Pi
qgboBJPCMoGDs3Gzue7wM2Hu9ourHk+RCFuueVtEj2ERkVJt0Vkb5BXXiKJ8RqCJ
D8tkXVU/zy+g/YYj3Coj7DOGzQAXP0GJoSfeH5xINmIrC2HwuN+fJaaKhBzLFhCe
e4vDo712OKYe1cFexR4n8U4UvI1uioengjHcZuDF1SmF3U0+1LWxmp/v/XZWvO7i
wG2uFqAwS0JhddKeejv8MjtvssSusMrHWhZoJ/QzVE9U8bDortHWceNYE6wNv3de
I5FHhqZ+2weO+0kdJy6nsU5LJx7fxpeXDDvJeePr384Kh+fxJm7qqpWMyYtXxguX
hJslP1oUd9CK8Vp1CwImJk0uEbyFMqAVbfGlkjw/LJvR/22jnzqoabGnTUuEgtrh
hvQEETgb4hfzT+/gHoWbPX1oht4iCQRidQz8paGJsy82IW8Cv31IWlaUmwPoLNBM
`protect END_PROTECTED
