`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wryOYioBO6eXYrveRSTAAEC5eusNAMkG7ovtIHgRdbE
B+vyyqHVr70R68ILPW8HRVpp/EAGismFAuExm8VHgB0yaR7ip8dzxAozJ90Gf/z7
ZeLsHHcMShKmHkiAKE6+3AlHimNoZr31/yhp7rIsA2SVEIQ72FLsz2A26A6GM8ww
nrTK9Y7okc0x3hjUSRbVBmJug42zD67NpORfb/VU3O+UFHbQh8v5UHsbVUbl1tx6
VIxYt0i5DJrlMMNo2hwW8XKCkGQKuIeF+qzYR9U0scFuTILSHFQKznqO0oVdrDno
RK2nf+E5a2MegEtNx/d8TCftpXilA3mIOLYSN+VhWuna18CaLtHoCx/wtj+MrSup
iWSkcqIwdPe2U02CKRC0CK60YZvR+ah7X8qiW1PEC6lrZ5FAhzVLTxiiaP7ock4/
3Gx6JoKKhdw0pTq7iTc7EMc0z//4Xk6JkguWoKjkpic9qB/zJW/GJLdLCg1fa8Yl
G6ho09dUNUINqpDGiDmGYVSt1Gk/cfrtEkAd9W/NqefbCaKuFMY02o1DVxYOy6TO
bfA4iEt1RsxHA5g9LJqgb/WlTwFua4jjNQgqB6VirjibU0daR3kW6oGQDMTa/jOR
f2W0rO0fLUzYif+corXX/UgESIhIWoFzSlRvUipEkCjrInaERZyW8LbzuMVuC8Lr
HP4sNwD1R5XseB8E5P2Gvyz2c05zV9podD7NVM5Z8/6t0kx/SPQSa/mEfdvroHyo
mE8yxnapefp/VTS+ISbCBQ7nALuivl6jpksW/R8DpF9A9VaEM3kOKXyvJkUs2pAv
NyM80pjzhm2w03FDw7Ddw+ITmZ+to8Pl3M7WkbuLLw78M+v6QGw9W7zKHfz4TnO3
Yb4ZuFjTnMmhYMT8wYf531YXS5x6f1EQQqX5N8GxUvn2rVmOli+SgWcOEyTNHTEL
HT3wxNeoepLh76ARcE7m+orqhflD7+NAvZzc2yFM906xGygZ1fH1EDc8Hu1mqTQD
TfZXUY1PuirvMZgQrGaVtjwaV7a4zcAeX/UGONM4qbnhRrGDOneARISzpdCN/Svd
bHcB+LP+zrBwu3jOuPFCg4cdepP36gbm6mdYXG4YtWyRXHRvG4j59QLFjj6aqFtB
eK49+7kFxq4zNr2e1G6Dr5rI3xF6uzY+ZskA9yO4sHKQuDZogRiH4JNbsSBo31tx
AVKmycYdgQUIvaCCPoXwVHHnNQCFSLnYLEtyQHtjRkuzCHo9dlXTTQJL6UPMVZow
sMgG/anAOhECwexe8wzOJ4gN9zBZ+vBAdItqYkogx9m+fsUF5nYWVG56MI7TRbPz
RKWuVIoa+hF3KITqncdkBcXe3gMFH4g56tnRmDIdTOEf9FbBbofrBDzcHkPwepPn
JI7I70tesi0Apf6o5hH2Db8UyKfNEnqkNBbSD7j55/M7CBQJIC6RqVuLZkOCmSeq
RFcN23mcCEYPHxgXLP29zp4xj4OKdO/HOnu0piao7Jw8H9sdhqNPzxcv/Jp5QFF3
dVYjWpklxdV1AVFZTXjy5PVSFGkIAJhjJvixKLEB/EttFlvAG/Mgx64YQGKgJg53
0LiT9UXOlmksriHAmxEmum6XMH2DZI6Jx6SMEyKbYTJDbGFvI1Qrv4MBUW5kl1t5
ilaPZE5NXiJo2Mvi/YAucxQdcqSuSEErpGkFoHDSagJahfHE7E2q9Eq9xB2XezVF
RUaWF/PIpSwcNWbP40Nh5Kg1M70mL+fBnWp5oraBGnWZ8ehbqfPIuhMgnNbbJoc6
LAe4od4x2FAe0gHf4OTsWBNAZltczKyf1IUcXP3o9ju6jdmE5tFUc/9ceoI0b7DW
gMmvedkrYE1cMIE6mf45ydVEZ9N5tdTF5YC3tC8U3WpKgai4J+IhMpVsfW/0oBQo
87nb49mukeB3OSYkyYwGQ+hxy54YKlRulGsfgPETFeakVeQfHpkTWG1AOoCdMzi+
ayLvXzKMXtMj4bBaN9qk8Mi4fm4m6AqjylPju0jM7eJPqMXD+vMkzu3j1TfwPjMl
VR6SA8DZlqgZIyC5PORG5d0Ajg3HV1sNPZVUT9tEcxi41m/Qm5X2OnXeokUB7Yf0
XgpcuTbcw9GXZpdUAIlgty26gwkHOUHiFFGeiKeDFK6XmmYGbLI0y5//fafPL74M
LHL8Nx3kRIaW1hN+1FxXS8+7gdU7RLD5lM5vzMykV7haWMWJ9c2iOq+Cn/z6fgAK
xL6C9vKlQNbCDbmYbazfbnTj6f4e33ZT/ZkDwudgzwyM9+Ezo462beXqbyX8drm4
dC7ITovNeuR0PJuf9WBziYPZwQKPf97bKULUq0NpxICvIFAASGIV4EvPtj+qS0CN
n7fLYdsrlIH3daVm00CIbSmOmeVgI1HWdYooi8ekoF8JP4T6tMYLfXF6g4QhGjaN
9WtA8ptXFOxnsrvYR+jGstj7pONbnaOvg+wbNPsH8qGIJFoDUiYGZSBiqliTitlO
MfoWI5n8/WxtpodSxEZ9dYAoxRXYzPxfqg7CeXs6WF7qcecZzHrJp06TSw466lal
zCiHItXFFJ4Q8ATtwhx5ZvgPZkOOw8ESDKEelliseosiICQ4Jdgrh7tgtqetqKQ1
FRkJ5yVQLvrL1zcOPPr30ElNW0MSK8L27bRvBDM9iLWq2jcmezmtH6p84crcYDaz
g2OhNjQNwDrPFjEuLbkW3ZJtxnwygiTaeTLdIwxnY9Opazzg5/pR98irGM6Yh/No
mWFfpBVVe4UH+1rqb6JZUg5xLxPOLcV4rj9kr6WHB9WttSB4V3SyHOiG3XukFmLR
D52vX4THmMw7XqvmiVnm5ikkqEnddsv61UPivVVqi480x+bXoJ6fbLWCQRldbrOZ
ilLYnP9i4JBxbXJpL+gqfZMKJuD3vEysrIxWZSdt2nrQ8xcnoWUqxFZ90fWSz76o
3oir+amiK/HIutteq9ujZg3+MfZgLjaTcGF8aC+2ekQwSl/on9NXOCLNWby4HBkT
lQjVPy+AJu8NSqZVQiwuJKZcXfaXdsTWBNcMPjUYrZ5S+JV2nhZHs1JhpJtz4M/q
tK6XV3EVfWyAzX0AykAtSGTzDHjhUahuKn2X5RRfkQVq0OLJeq669RQG47U1n/km
KHhMuzUxogk3gM1ZLF2/Y0Pz7Se95MMmlNzm1vVQo0izRPI666RxBiRXPPkkBzqU
m/AlisDPgtb9BtRl8AVXkqoJILyHtvwN0Gn1lbsZqnOX3c3OCLT8yXD9m7q223Fb
wDmxu5NSH/LbPiBI5Abpq3ABqm2/C0li1i+mJEwCYKvZQ90LMRyVnohAkOrihWsD
Pp4b1+Oa88HQLEjtZouuw95NXu0axOb7CKhHHS5PI7g8S0jh4xE+p4cUH803jpSj
/bSBZNk54o7Z0EPOzI2brik+OUuQNG4OM5X56CFb6VS+2cjNC363jKsgAEOjJYH3
QWXM0NSU9INVwUGughfsuR2PBITWODgJ4xCgFH3ymlzqYObbcqfncF1nHtxcT/Tx
KxgFN+rsVTNFo346RbzHjs/EJigKQnDgcaJ/yg68L1kndxpUDU/hAbQ2Sa+vaQBY
oz71Kdv85Pd9ruYXn+u52jxzzY7Hu0UX/jZmpt64LMA48inzlmihoDOvZG7zliyc
NEaW6svk7oRk0AygZF4st5oemHgkz5yc16kvBraBGOo/Z4UZnR16KTedRhRHibXi
yvcQuj/1czpLOkBsL+qcm1iPyphPPjkHOcB0ExxrfKmkeCM03PoL6LEwpqXJxHDW
X2phm+uquGIfR5G7auK0gkbFOIgWWJC/e2/NwvD/RKstyl+3roZmCUmAYata5Pjc
sVP3PoWVJRT7JFF71bbgN5zIrW4ztx0hYkkUVRUQGBalO5gpINzsaESHwu2lTIj+
yHbHyeTo80wFwQx/mYT1jxwMx3eQVJ6P1MZQUNKo6wk2vUfVrkLHiCD2zQzUlEF7
2MOZmX2ELp5t47czHh3M/D7lB4dEpvqbzGfEbrOBv5HqXCloj3jOfQFUv3i4l1rz
Q5AWg2r+Sz9TLTcfsjA16RhlYhu0ow333t0sW9JVcrqqzGxXx1i78S9G/G/lbmWP
UrYY17ufs3qcgMFp9LsDfzF9rH/lpugKBlWv5EMd2rNAAWIIji5/Hesnrv2dDVUs
5ZUmk/I/PNhSUre3PT6MBdBsz50JX9RanQvKKa6W9uK6efU142S0BA5PiPm+cd2S
HaKE8rT0Bg1P/vNpT6TlhKk3bH5dRTjR5RM+VK004yxb3U9U0w1SsWP0TCTFIY3z
mkE1dlcOaOdQ9BO3A3OysD04BJHpqt9X3vHvoNqB10N56QDyM+ZyiaVkJKJgJNaB
XLnnQ8Ng3Xu94osbyFaOvaLA/E4tJ8KjovGYx0P2Lnrpuv4glm52kbZ4NPF32ZPG
GQeHQU6Zb/Le1o+2iwWQ/YfqqKLXgL85JHRA2NLK68zWPtZXHxKXP2VwTQ1qtrqs
CynX+VOI/eChl8PHIhbC6l76X3o8FagokXGTw8YQcB8JUC8bV7D1WDSEU4YMK6U7
eWgCbrSJ0mjBikni4TLik2fKr8p9u07AxEfvnj0kEFBK9JHpRbWp4L/i604IZd1c
LsEeg6j9qYgZZttisTli5K0pr+GMjXpQQsigIBD6qYEniWhpbIx2xIt1jaoDIODQ
i6T5yXEd0p/RVLK+89uwFSWq1aQwluUkb0gCVWhENGmRB6GhRxAEMzrzduLVdF+p
KaPg5LncUgAGINTgcoi1tRbmTFK3TBWffzSTHLyqpDe7LyMZiQms9Ntf5q+b4CIK
eGblLKS7cZiuD9gM8ePedM1N4vkd2whfjegXIJPcgxvy8EE6yhERVLJbt09II1cV
OE818Wz30fbWJKqBgFdBRF1BAcpiWrx5YgTArnsbL3Cz7G7vk8FSp/0lqLmkVRUB
5n5PjM41Zkvg2W59t9uOuDpq0K6rf4mIibLqIUZOPrgKrfGXgoL6HnnlnWzXx8WX
fyw0JXAmlggaUu64WT02OgZEQrdXGFt7tR9I4xt/mbvQSE9qHmyt8GciYal10kPR
xncReAdU9llnCHh8fR+GR5M1PHt1AlI4ILo0sAs5qVGd43WibKDDhLtcIYXazX4T
fNzAkJ/QH2kN/jduMgLbnNtBWiYtQyZ+weEwnwJjbnUebt9mhmzW6mj+HaqBU111
Fzw1Png51S0Z7gA4S4PIFvBXr86bglPq31NUUXODej/iBOVuulANcZ0ixzFdIaGO
roL2FGwTR/+dWTrONYWzpbGyyCizgNlyuSQvAP5JhHHCSzaIhvrWCM16Lo0x25lS
s4WF15Ubz2vPWNj6k03yta4cUJvuX6cZMExjEOmSkg0k80+BYqhqqFmk7JfFaGoY
CA8atWjZgFkAC/W+NeZmF3unBeM13JttQ1oHX8609/vugi0POKQ6XoO2Vz34kaRq
lxuiaEXnqCLQtFztiS+RmW22jIZjxaKloQQiTN3tKA9NWPpWrSFl00i8/s5G9yTU
5Vv/g/l/OcIF73tpJM77THGLG6jcIQ+Hcd+1wUASyk/f1TiGgWwPn5PoBS1HYLuj
YcskhB8ZFgRBH9PkURXU2giUjM2uhxiYONncxCIu0KJ+iwZFX1EwxSK5bhCPmLW4
MF8Jnt1ENHlAOkP+6MI0NqobLl3qeQrBs5QQcmTX7wCSggS/0gNHK1ddwKIbzjl/
1cHwDQ0bImzjnuK+CO9uMCT8j172Aspd/2SxC8CXWdmPF7d+g0vR2McHD/axR+L7
e5fLdyUOZlNVY0VrMVYANOuHQyYNxE/n0MfdVsIBlVklP23mqjcXIwml+1sOIbSU
TqhBr7aGZ4TY4pHnoYQiXBwNhfUJzwJlwSqkBILO/YW08FILN7xP2tV2Z+h6oCwf
+Q5UtdZKxfVb05VwlRMvJMEBcaiwsC7EhALgutJsmTkF80BXVmNkV1rYIAw8BvFF
aStuW2Dv75/2z0ymKcya7b+jOPeVULUHoeSwm/FYFjKZncSffv95OVfGJuLC0dM0
uQcMaf2ysiVfh46ii8g637lUWpRb0/xxIFQ17T9hXPdwSjCxAjxVMvt9RPJD7q1F
qJWAZmULB+oQntoGkkcwWBFe4CzXSwVrukYWwBrjyfFXQ/iAPJ31oWgCiyuC0SxG
eAH7COzyoNYmcTwLxL9o4F0D9j8kXu/tviIHXHpyrAMXv+2KRwUhQwyXA9uDeWuX
o6zEYZWjw/PybhAnPWro2IoiXCQ9GJ8QSuDAvIRppWcuwzckBu/KkceH0kQVFZ0s
e1gnvkb9Xbldi4QePVc0gZXkGTtxgwVWWvy09dwbvX05LdxCKx9ibh36Xd69/S/R
iuSxhBLbGl8w2HlCjcvhb2WBDCbPFQl7H3oywA127OpXckNEDuptModGloreYuly
a9shuCu/q3nHr2fYou62MSoVzGBgm+5tfc6fxryD4GsmruOm79zId0KJM8e6w69t
MZS82hSuQmhTlglOhAA93uQOaobHYsyQjevqLZvTFd693/YfowbLBG/CPw9HGa4g
vtofE+hXTUjVYF7foaySNvggKflRMgBP5vlzgcaWcGUJ8Eet2fcl90B5H83RB28M
OGmnyIbfpRMeNv/Dta3Me2c48G6hnrBfyD/lBsQGiY0Bckgg/94pdBAi3cIqTQUI
TKpDynol4GtwHxAfjthRbcKLj78x21JXYewzHqVnCLW93imgW1cZEL/KGSpkw7j6
T3uxFvSgVJkWG+b1e9JR3FAtluIkUQMgv8t9zV5q80mJhHDJENoyP+akrx2YXvU0
3k7jRsAykb9jkLhks7WxTmydLyfd1Aj6HkOoVIEBBD8icd/6bhkRhgd0tg1U0XRG
UT0hRo0V9We4U5wONmAnU1G45GimvqUAC7TGz0xbP775ndaHWq9oS80MVcKsUZ6t
urqsXQuVoUI44NzbADgiMNvWirxS8cN+sGuaF0SU5X2wBpyN2r4pBf/DAJQ8WWzC
5s3XbHTrsLaDpOfcql0rPt/NKKny86leV1td1opYjEEDD15QdEZ3D0fiq8g+3U8d
b/EKMrsSTfSISp81CPZRgn71IE0luugNhh0nwToYBnBgvM1qiniNSPeDkZI1r0eV
fkeTNC23lyLZppwA7vFxMVQPPtNZLnIwOvQPrjtdziH2/SL9mHXA3rcaRhxdFuCz
o4LG9w1G4d8qIar2qqyrEj4Sb0vg7UA1HdWH6UhzaWZkCG7wZjQb601JVfD5zbgV
AlajB+1Xd8KitUruDBXS+jIqlNDx2T77kg89EZhypYSTUDBOu3e6GgSKwkzcIYws
1h0hf9YOmbyAHKeL+7p05WuF0Q3Gn3BtH4rPUtnOtLtqgVNIVdbqx5D+7m+hbRsE
4DTaNsqxN7siYjnV4Bz/zGEsfDxR4a9+MqIHWl6II4sqwETBWqqj+h2GWzZ/QTxb
GYs3NRsH8m1oPnah8Mf7bIeiwrKMBqSOyQ2h/QXiTzYRTJkwIuIAzhmp6JXqEtVD
HpKsu/HGWgo0PcPElE2jN4oMvVtU+GVbqFaTffcJyJPY8R8jS9Xy/yFql4q6mJ5q
21jLjFRYnqRfyduXoeICOMU6uOQ3pJKz+gC1B+HW8JIzOfnhphC6DbkBqRedvv8/
ix6L03NQv5QxDE6gYmk6TCtlVnnILVIT4hH32wowUHpF17VYTgQnnWCGRvNrUJ7Z
guDo7z46sdHPt5mI5QE0pxkqlUtEbRisG5RyzsZ8k8yjggbTOy+jMX7Un2jMTlSM
HTx4oPL4SAV9GIDWlkg7y0MbaIY8DXeKvci34YOyHncuAUjPZXHqfroGUFjs0L2I
XZMcN3UEbuSQkwBaW20GilUKA7ndElA53Lr1ChCzb0pSgR4yvMwN+ZBtEWqN253G
garF1NMeX42fyO873NwapDF6Fz3sZqOrI8tsofhYP9AESLBdlMqs/N0BqQCBipdM
7qPtm0vXlgXWA57RcQ3sjy4X0ujzm1DNa/IwLVrsyvPh1eSYaEayxz8NO9ZK5edn
sdUDUN3OTks8aNdaKdo7AQbhUyNro57Kn2YumgDhWbdkA8u7h91/mBy62D2/Rvb+
tDP+Xm/gA2yduZRgJHEb8BLoTaJj1qmu/7An112qkzJT0W6TcrRMGg9bB1qEDBKt
Xg3oIJQOOkEFnk1sUPsRHZLJvCaVO/vXYx01l3cKta65rtL3f4oaPegsF2l9jhSa
fixw8PcCuJ/8NCW0E6zJAuG2sA397GwfM75JJh5mP6m3hqIskcF3NJoneM+aFFO1
lmX/Ojz8l6RbctqH6BKLYg==
`protect END_PROTECTED
