`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJkL8dZKQ8U3S5qUvwtt5goCt7cBzZKYRoHRsEFLcyQO
90Ev2vwAbAvzYr4iTWbgzjocv7sAYGf8yczywbMTsXQgp/mthG4BOOGWF3JsCo+x
X4GsVcIZ3EeEmKy+l88FMJuV0WZisXZA69636Ome8ammZEPa3Ag28e60wlNGluRK
gy7bLAmyccBJ74l0bMiCag==
`protect END_PROTECTED
