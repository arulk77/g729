`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ffmyuUfKxKglsTYq5oq9AAXv0TJjWdWcm9DZiVcJFcoqttrP22+I+m1kA7gIcQW1
Gjtel/HTzZGO5OAj63XCKFcgIYhe8qsEoxwOQG1ajSNAf/XkwuqggXRiqo0AofFZ
iaGfcnAVtHdM6HqyNyFSXekLDNhl9WEu7Z6nLuiW8G763hKkuc3IlXsykHVVk2eV
`protect END_PROTECTED
