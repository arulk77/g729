`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
if7OW3neLerq5QTb0GME90uPJ/Er4YdAUV9MpDD8CQtluhwWGPxhbwTuIbgNa3cb
mbKKPzDQP00fvrJgm5OKAxx7t9SLK8iKuIhAakWs48apT1wJSWloXsxnjxvd6XQx
p/6BtCjv1d5ex2vMxwBaBn/tm/q6LHnJqB1smC8/SEfqFUWe0nqVDrMUexfl8lkv
LiilIoYITgRvkqT8z2qpCGc2wFQnsOkNfDQvuQdja3cEOLDhwY41f3Grafbwb1FA
pK6mkYnrhunCLkP8F4PUhDkkF0ojiPUzMpiCH/hkTJzUUXo0YxgzeeMRpnQpasJb
`protect END_PROTECTED
