`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOdW3GfAkl9SFyzyJmKqcIHue8+NRg7Fks9lsaFGqmYp
tZ6JIjEGa9HxgSy10UqsmXIMMzwZ8XwI6JBRI9Wfpj1kmgSlEVCsl+zxVBM6ppuh
FUlC94FsIGbzrJumqq5Gjkwn8c5eP9+8IQjPRe1bWEEDTLRf71lbRF3erV2obSyB
P/zKe5ehsdCnNMAlqY0BYQjD3VSHYDdmF5DvLcQY+ZneIHJfR1BW2NIYlBtaUvvm
+Nq2R4MQ7Vdy+aOpkS0melsj2yomhin5hFKOPZnlUAkO0IwQIo+SVZd9JxzdVsmf
bTbreylS49ulKQrA6N61QydB41ffCajhPfUbNJikEObBt+q71aswhs/DWhJtiuj2
ZlwFkBRojKx4I7IiYkrEYw==
`protect END_PROTECTED
