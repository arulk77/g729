`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
36A/U5tO69wVl401zVMLLYkGp5XsJ6kXu1cGNGMJG+3NtZXfEhKdIaJBBKacG9XS
+366Rf37NDfIg0j8FejdqJCInIF/xeOModKL+zXt63gbRBX9AEICj4VCpXQ7qOcN
v+0niE4HxbpJoJLdARpCbft8TNkCPOSKjgcg1cGdscWNneATCxQyLlgjr/CZbZEY
32GEEfSvkjBWa0P91P0YuMSWxg8dLsLiYKUaDfiE2zO0rAf5BvCc2Jbjd3nM0EsY
s2ww22C+97Ce3WMqrb7/uYQylLKt+B1TQN11yuz6ghbqMxFfs+MaqWuLj/mYza/R
ttepQe6kkvqVxXT1LuwCk+f/Sr/uK2Gw/kqfEmZrHk9tCDr5fyWByCaVvpzgEfUJ
`protect END_PROTECTED
