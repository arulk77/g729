`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKuGfFnt49BhN0mZ93LytkI757zCxsCXIB2eJBzBcjdF
Ji5+DSMmWbRvp8F2gX83SOcM2CS5VYX+3CIbIbdut4wKL2cROrHXYJlD4tSb9OY5
oWx/DZCUaOaVKaJRgkTeeqFdUrz+gFRMqSyLD778T2rmIdrNOX3/VQHQA+1yfcvm
ieDbrwc61rRTcH1tOLQf7hILuUzODqt4tIQ/YkhAPgiRZNkkVm18YyIVVDaIDvCF
ODmEWUVnpLvIVv6ud5IY4Q==
`protect END_PROTECTED
