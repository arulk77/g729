`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
S1gOT+i5hH4nUrP+CWA5IcoqBl/IGlXBvzOl8W/Enh9ovuTRxgQMXIeVXGKdi+hC
1GVy6Lj3qYLmGaRb3ceeCEJptFGnGO2kX1STFmtlxi7TSK7noWTYevJfFOhUJ8CA
`protect END_PROTECTED
