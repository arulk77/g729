`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN0natH8my5RvIW+LsaldGIGmT1PhAIauQBKXuy1adPZF
siDIZZQ6U9CV5PYYOgRUQvZPcVVA5q+TO2ZtbDtsw0BNVzhafcegwuShHEywPadv
EJfV739i2tFlLc4tqhhRPWGreQpFEp7E78Gd1R9TMdxWaIU8JTGnzwmFcCuKq9/g
hv0k9fgw+K+byky6fmnBpY+pZ4LIBp2Z8dL7+9nI7mZxOqC5+OWyFxiwehgFHkpA
Kmhi569C50AqEA+ILCBu+pvu84Guq2jWC35xQzGjrrrDnlKwG5B1l1xeahUKUDx+
bTbaFH28cepp17ho3yzy8Dl5gH2GByiXDUshwXPts5NCF+yb33vBoluvtway9dF3
h5osFBW8qBhBTAJzzHpHvaEchHlyIgtjOAYRTWDcgjHhoc+vCGUADCTIb0pzCja8
qc9uCgAuX8hOVuZUtX/0SNeLlx09N3jjmZVinZ9uGcFQvA4NwlNcLiHAUlSJHl/x
Rohb90N5Ny28QoyOilVqacv/KHZ1ZFCWuV6rwHVZ6cVYqI9T7p/Eb3jPnM0GTVp2
URcisXd7vqdx3nCrOLUaXZbHp8KAhsg8SM2wnEo0ytvUGL2+bA6iLujOc2XVQBTN
NSKUuNWKeJghkZVkfKt6DhB4XsEBC/0Tnc5u2OLnrKHpeQ5Vo0ayJJfuNW//nbXu
dDZJG79VNCaF4/DbQ8mmEJtcL4PFQXGNUevXcnJFE2lJWdtorvkC/HJe2NkoMk9t
EVsMTCbgBxTeYojZkko62caZIwu7q/yVXZp3Bjz7vyjmJOF7VqA5ykJ8iH3p6dcZ
ORcyDFT9bgfq3/zBbNibalBmoVNW00y79MLXyScRxmPJtCoyCA4FafzqzEp4J5gX
VXryNxr+Stfy6EfjNhZdSfaqVOR7YNiZfbMZSrkYGc0W0RH1E/UwVO0yfJ88+XqI
tlqulGTeex/5wf6FPVmrFjrNR9baewgUyz61Gu6TNGH5IRB6ni53g7YU9MITyaO7
YFXAWUPe6N809MGl8q7jpbgk1leDl9E35Nkegh874l5EEs27IBpGYLeMqCCcRwvs
WLcQ3Des4+c8KQU9XBcQNhc7TxrcM6CutEPtlhfmLOtb55SI5z0ITXWbgfuCt7cl
66ceHbYlLn5L/vhi/tePX3KVF9yzMft2XD5cvYPuln25A6thK2//FkuGYWMcnsuS
3WrVEuXdUM7RsvqdK2uRp7FwDz8qleMgfdAtx785hEtycQelHi8Zei4qVdMsqiuO
qGnIJNF87Sekv/KdG6YJ0rdop6WTBIJm3iDaVJd3tiMw0YQtZ36Kr+uONHV+qbJV
fgTG7Y24zOckfDy5ZQaf9BmJT9qOIAvydQ9aYrXWKBhmQWZ/Rvl2HGYT+R8ZeWN5
5JXvj8Az4nuGKnuxeMXX63tTp0y6ad0IaOfvB66rjXzm0eP4AhZsEfE/WwBtwbck
zd5yzQFuQubQwAutpOwEpMn5bifcbA74n8tXHtP3YiCYus4EC+QkQ2VAuiTUIk7V
bZlQUV9arpyESAIlqXCgzUGkWuMgfpkXXE/kVBpqXN9rLtreWwaHsD00EywWUpd3
7z36XfmGfT6TtM8/auHwTZIIvKlLAOzbTiofgDsZOFrk6ZvH+FH3sIaEwAAb4ud4
0JUnFrfp0hlxtVoCGN1KVs8fiaVzHZ84FgHSY8vmIBBxyH0zErlEdhDJWXxWxqAe
2rrfP9iA7RPdJ+xj4G4EOxsgjEtMmUkXh7Cg0Ey4dF1acSnZ+YAHFO1ZQ1GOg2wY
vSPIjIL81Oo1tkajR9GCiOKcjlr/NgpJWtRlcR69Q1Cbm0O9rgfTzbZb9xtgRNvU
URC6trqqC9kthIm/nOGzNYYsP1ubl4qulU63mUcbuBhd8Z+VHdFG9qwffLpnyu1S
SYoaWoIhgdDGubWM52WWncD8BevImRfPmKJf3r8PmxFOz2Z2ZyJ6sAdDx2ecnAVg
Idlz3Ou3yjGNFMd6zsNHe7EC2kqFjbG3TgUpbsYbt1HmJQ3TotMsDtE8PJr8Uq7u
hkEKSUWWkpotl9l/dLIHxJuEy6DyQ939MikJh3QVo5k9U1qByuUK/o5cLGk6lCN4
BCHtQy+O544bUyr97D3evQ==
`protect END_PROTECTED
