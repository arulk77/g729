`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL2UjfJ7YDDxA91xywQsX7FroifrBUIZUGE/SA7rmlVT
xR9CKVIvvC19iC/QT3TtSm92QjHykf3TClnE55P4p4RURkOhlMmNpicNiqn4QnSR
s9uztMjcdf+lMjDCU5nVntIVyIGhb//554WfXgSKpOdmaiyYKl0PypNhZ8PJw4BU
dkLIh32t4JE1NoKKwKmjy2hlK6RVXDP+ebHUUwThMrb1So893hQ0PIqP6FQa3VNY
3I/boJbgqHUgC4DF1wSiuVtqSKFDjk0noFegln2s7523FF6dC2Q79PdJBJfpixH0
FPuDOODQeC1zacspMk+8UX1IOu1oabHUcN3Gg5lTE5seGtPcrqNQVe/hLLr8GHbV
`protect END_PROTECTED
