`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkSfXivzzsFCHz84DJjk7qzEDXfOTozwk8+LDw+9ZkitL
UN9tMQtQi4bx6iFJb4A+2ixie8fs3aEgL5WYl9yw/XnwjILcPZa6fOjFPwJP9hPR
PEtnLkDotogXsdgFrNDe0HO/Zj6GdL0H0F8wZzhz27TViF7VP8hzd9mQ9GNH0Amq
tLltGZ7zx5mYmFmffU/OmWjTYqEBSjXuOz+7cOWO39nDbLmQ5KMV+JvKUNdGl0pZ
+XLzLghc1ecmlP5WAHeY0G+TmFotHPIiaFjiIvo7N7pzzBNKWj05gaoGvdc1hfxV
RjVecaG06xVoVmBfZ4z8BAxmSeSvdo8vZr9GifFtT9cYVChuus/p9/t/mmrgqwmH
0cLigwys3wD5SsA8Mx7TYTv5qxerRCwUVSyiFkAkLAoK2d2MVI4X8s8FthhzE03q
CpNVoaFs6Uk5Vuc4HKkBc5T5q5DaVh796eUEBjsdq8WSnfpn86AK936uUJ5yWz3g
YJv2mnXELwvAcNCKCQerV08YeFz2UXpNk8xkl/wBk95iHJzm5LUrAKMtnWoRXVIh
tP2VmRtqDNe6MFvLgDrqrYop3lcCOwHMQNasiTZUU9Yva38OhUROwSWwvCtoshaU
JQO2S41G8ID2FkTp3XsHA6J875D7S+CwrsGBh6dmqQ7qmhoHe6loLeB+CSxPpiWl
/XNZpI2vJwVY3nBODvFnN+l3G2xlfStLPOtHFqvTeoXe5Dflja/HwpuqVXpHQZD3
DqyHbwDXyAPcjVagpOGddEwpcX+ys0cFP3OyOlCyeVu8KN1hYUDPJ08+bhiJWeky
eXoK9rQJUoV21wAxevO02C+OWNERGi/ujrX7jEJqSj1sEPrjYZPC1BtVSNocJYhE
PFEzjVHe/Mr+OfLFwGl65f+oxhmA+70BRDrOX7REs+M=
`protect END_PROTECTED
