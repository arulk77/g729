`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47snd6JdNX5sLcVzKS9RsQnYNA6cx7wnP3Kamg6VxxHD
2192L1efBStQOiGYxqJXEmVKQnvAfaJ3hDiz42fwqmeb+JVyBKT49FWRmTMofY9C
YagGqAHCvdK5eVfNCkg4iw+nPXuISyhQAYMRPAMH1yjZhUkOGdPQf8JrAoocgZEc
PyRPgjGQy3sUWKchC1rvOkqb6dLBce7eTxMYgDC1lXy2Cpxk0H6ywCSFC45QDibx
l1WSsML1kZ1lqp8D+HoNLa0TsqyNsZghRSYeqkWUy9pLLtlxJYosSBR/YvBAuznv
ok61TbPBcQeYDT11mO9QvhJVVOKfRnNEMDRwhEpO7+yzg9USXuXwD3Lz43qH2D5w
Nqdm6T+s17A+vajjiWmkwV7HhqjmIr3CueLbLfUZ+ck7vTR8oi7s7QATm75Bp4Lk
TjOZd2sFkSh7sdJNSf+I7dq2Z7sFxF3WP7r6PBv2fwmESL+Ap7gg7iKqOkCAzQJU
`protect END_PROTECTED
