`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDATJ8At9Vgi59W++vuAkOFsuyPM/0fUF7lXSm+/vBjc0d
sfyDz2TlOlaPD/gWyA9LgEauO8He6Urf0VGlACEkWVY5npSBPN4fgrwpX7fsAXuY
YyMYph7+ao8cexkmiJ7O7fBz6rYrK8ia0ChmFT62GuxQiYfewk6yWDdsJe0x7NG2
QJz7lw6gwwc5trCp7XjORG2sY7+r0TrnuKxTpxy9PIURzEHExFlaan210nqkMdNY
nlSon09hNZZ+E28a28KPng8F4pAdnjIuxh+Nv+j+pATC0pHyhsbPZ1xGCiPXZAAe
pP3SqcP0QtvZhWkNHLiI8PO0fk90l7UWMbs+/K//Oxv+TAP/eBE3e8k2ZkE4JMNP
y7AOSFWaCT6ISsPq0uJU2SNbFd/EjwGI7d13H4q/su9SjfPJht5Iuh4KcitphYee
nIs2PnO4LNwq3u7kiKYCYYbkIOjhqVlTIeBNq3f+v1eperPo6XzLQrFRzWS5IuaK
SWGlZY2LHyxFcj3emcwylDco+0ODcGxdCbpqLDKicH5b3MbidhBejJZDDNoyI7kl
e3lBDqnzvh0XKTQuI2/3Jn+fV70IY+PnotQGpL/YxOJF/FbnQXGbaTSe8pA7UJC4
qLIpTFwXZ0TwcswCRek49naSDuzRTaTdF27oEurC+osArBgmSrms4vYo7l+TFprn
LiQYp6cixznBocn1+DMMcd+6qZfEJS6txF27cKB4Ctgeam0Bka0wqCJLXvxfCbgb
313TQh5uQgr22u1wW3eO8N4wMgcVwbqox8tC2kUyRr4ABDHX+tIE1s7+4weWxHx6
igB4dC3xNqD/T9Qd9XgaQlfztx29c4oMLu2zZpEe+1O2JH8Ka1mte3FSfhIkpR4E
d/fzidrk9zfGn+Xd1HfJ833ePgOmKs4odBcHRCYzMFpNWN6ORV4tgI0eX78wE7z3
XSxhhe42Os6JJ5/EFvysCshiuKU6SbLbCS6ihOwT3qKmNrUvDziYj012UzTiEYxg
eJ/s4F1T/sKPt0j3CLtLAiyN89foXIsmTKDOCtBqnmzrByfAa8GXnKpxQkcBf+R1
vc79KmQ9QL55OkZS9/YPKgBOgTqOZxYFAWOQea51bP2rHO6AjISIiexiHRBYghfR
aFwLpT+Gs2QNsDRQvaCLpDGVQM+2w9ePOf/BvsdmBqefN1IncPrxaJ4+GdwzbWg4
EZ7QffiktSS5qQBI9AcRTyY2g+oKqbZmrE9uNodDrSjNy3MzzFmSC9g8vpNFfILZ
jw88xM5gQaC4iXwBtFNR7N9Kp4M1Iual9y3f1nEbxL0kBh9JVnr/dISDXAfVTfAr
i6zJF8dA+4VxyIPtck4i5mQri7WAumbm4pZAEWxdj3+BQolUOnT/ziHYmurqQn4i
ZAI7wgIhlcJMHCVdXHBGHXrUReyFrXxQXupbDl3zZUu3jUhOpKs9OhrffrKuRuht
u/K7cuWCrFV0nZP7+t5FPZ63YM+1cS20TW5aKVBecwBayWLRytuC3R7C2ZuKBXt0
D/xnNK+cpH4HaH1uh0eSMfZDaa1Uq1APhvvw+mPTPVEB/oY8eIlf2qbA6ouB6EHa
iymgZ2q9+Svwk7ly+EWhNyx+ui7dS1WCv1vnDuTgUiTuV8MbwrELDiNctQalQzd5
BF67/btwxJY9MyX37WUo159XkdMHyx+YCLOTGIn2Tk2zeySuEI3qddtACorfrrjx
uHlTv8Gy5vvp+02LB7ukgtqbLB8ZAr0pXlKT00d9ShKUwmLeYt3UlCoyesKbvSAg
7ych6pcynNp1xc7fs9behIsBEbNZLN8wyaGK4rtVA/pYgXI8hNABHvouYGgrPebH
nzZcWaF5/42Cdol8cVVBaMw33wIxZaY4kSeaa6DUg3VtafZvSsNwCkGK881oi/FS
wytbS5Idc+1jGFu4LxlpFokBNuzD354xYVfrpfNuJMHbzNBvftr3h1wGGJJjNXXL
yd5/TnjK8apPodoolOO4C1TDok4j880pEPsecUie33w9/c2h5MAoiYtcwO2kbWPh
cEWhtGpDhwvls08EdeYfUkxMWSMW5RJ9OFYSgfWcRt5bBXZasnsJmE9xxFasTSuK
a7zyhIK1JNa9YL1dijKkFWtPIqYh+rolWP8lQfkqITijzoqyZ8VL041NkciWPCPU
nz8QC/b7duAYuCariY/iFyZxnYP+NMEZJhwjA8FK8YjBgLHhGoxPyMPz1AbDaCFL
sE4q9YJfMi4602AfBrGVBQOZy2UJ0SR/Jh9dVxSS7kDG+6EiUJojNx5hRPlNQlrm
V0GOf9Ys/hTkKtPTTy+BcA9MyzodJSt0WUHBzUt5ufXqe7BGUHiZwyyHUHkQRmwy
Mm8pvsFf10eOG5JVHG0dLaGrgB4/25kCtXQA9/wQKcwcVAHZoerggPISt62NegZu
xMyROQcHEEGRuOs6bl6nCn2FNeMfS1fJUO+frCHBI8s=
`protect END_PROTECTED
