`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDsymh5yDlJwzJGcJhjuF99yxoJGI8XIdNzGARONY4Yj
lgtu3pOZ6dv1RQzGcC9TM6ykfJdTOEUy+jnTdQAHR06AeSQGJSlPO1Pd49DsT1Zl
vbQY9Wujg4MoQpkEgpb2Imxihy/sXOgWN9McIc/y2fkGx/a7S7GeJcPYdK9CX+Mi
vnYsXEB8fqFxIzeO2Jg50CFxv9O8lNQwljZHnuUQbibd9FE0ddwzm8s7uftK2kKd
qnxsO3ZDKZZlcxdBSQnXN+ecdNweCfFrE0nUHkNvi0CLdseytaLrUsGQUWRfoMlZ
G73q3fXfuUkB20gfVjLr6eK+75Qql7OEsfeejBj0pcVFM0H6es8QQlhBJCXMq+9T
8o0FVkpIIMN0+Yq+XgWLkiCRkSfawIR40qozf2G5x7vlfavmCETnBPoacp/fy1Gj
eNyfkVaV+eM7zIJ2kYezQoIqwMDe5JFPh1Hirnz6Df5pZ1wSEHzKnaygU5YoIzAy
AhARhIXiqjt9+pKDSpWwvmORnw0GPxqujQH1vYEvntMAsafMofo1GaqX8Ffq3+e9
o82eYqKPVleUT/IYtdblPf1+gAJB9VS62lHmRNSpF2xiGpgMCnnRRSBNsWAFqsNA
`protect END_PROTECTED
