`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEOX+Iq3x7QLea4dFiuUNE+PtSxxn7l7VbThUV9pcXed
CFWYhVEj/GA7nIiJhkx02Bp2UBHNp9W6IAL+Ltm9qMhQ7m56F0MHbdsZyeg51izz
rdcnGGytKZnmIGFVMEL6xrscOdKuFfxWBWgQG8FQoelVlWY65he5TgeJMqfWCCz4
dMJDe1/m0cZd5mEaZASdX8I0nCh/Owe1LMGBQuuaMHP37N9iCiJbHMh8KYjiSHlu
FT/k9mMubyde5hPzhW7M/UYATP+1o3Du8tdGg4NNCq3g2Km0NaXw/IHhuj4Rb4oU
rsxs6rs0upaW/e0BjHP71P8Mt4sV9yRCAlbQgocMfljdXYfhmTdqG9wriI3D5fbb
1S0+Lr6bSAP0oQ616Xf0qg==
`protect END_PROTECTED
