`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKjVxINv955U321guDqwM+dalEVNFfecBg5/SVEOoKWZ
ZwVZD83v6PF/edUjwFRQxTJBqwUIHeIm7P0wIzL41C7xWnl04FoZQnqNLLDhlWBr
psdUZu6kBCrQvGJeq1q4cydjnBPQW4TkTQ6d8Jc0rKtT7L75LJqxodrU+zjixU52
3tgy8KU+59q4aeMnWaesUt3HBInw37d4hZoxMl4SGBnmgxerdJ8zB7NDbZX0hFnJ
jeWKCymS8a4FZFHNQha5pFIJm4nYoKk3o4biW9ZD1LcxMusA7y7C8FOzOHXJFO7v
`protect END_PROTECTED
