`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePfUZa4CHyTLmH7UTdsjBbBFSXl8gTyIAKETuaEBsBM9
4U/DIYmfP4Ar7+xeirQ+7yeZ9PLmV+zu+xD0Z7NReBiX7GHWCmoQzJ/R4yqlf0Ns
7/7M3tw8WNXRYGm2IxdE975/H9+fioGagMWTm0yq5L0mHdwK4aWfvYEl8xBiCWl+
gbtT2oXWHNoFkJL4NtdpxnWpks1YqM7zApNX6gEZp7M7z5xmsjJ9iExoGKuNXzrd
ubguwg9FM4b6b+ab8o5x0w==
`protect END_PROTECTED
