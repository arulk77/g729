`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAXgvZkTrVwz9W3qAYnyRvO+vLWYhyd+oF8AkXeinRcHU
LgABmjdpaifM3a8M0+GGjXJppQ7Lq5Z+3rfW1F2ByoRRRabLlGAvXCLrBrNqUaYh
LHsdYIKQCXjCBBCTDSOPw9f1bmzuOj2jcePyoFc5VoAdB0BIIhO1tcknMEnIe7s2
2Kz53089cNxd+4lMpxSXn7JqUu4Kq+QCdQWn2MSnUu5N4Z6UXrg6hsjbQf5gdQj5
T6NEh6J93ottLL682DNEZUXldh0QO7QJ76W4sFxJZerobc9EvQQza5/ovSP8LdRD
FI1PaPFdgbbTjApU/xJYc2m+0kbGsg+qiI2/Y/KC6ckJpNtKMz4P2Yc4XUsshS+X
AdHiDgy+2KD3oFNYQ/eoaGMlf/jho8TcPgcDQDByhFQrbDvXWDDvXncp1yZuFN8C
daU2gQhsuW7bPCmUhi8RT6U0pXadU/qd6APnm9nAv+XVvIH/CEtidW+rdMNSHfm0
DQ8A/vZb+eVV/k5qfqNqF1116KNlnU4c1TNQ/gz9vgLteCjfGDvp4o5SF3S+16G2
Qbjr5rMBg1TsM3gOtaxSFptmAzMU+EE04Cefa5byv5iP/VjKfG2Ye0IJ5FFw5hu+
XisKOkypxlFoNjJJwNzxOCX/GgEynma7/YMaV2wud6ad6E8Z/r8d1X7g09qgT96H
Oflwy2YpweNkYfkPRRtiKBn4QS6xXDUa41T0RL7Y2kskOV8g3KiZ0FLyqX7xHsbj
yDC4kfl2YRHa95oEZBDtIO+ukUdu8cGl2HPaAYRY/TllC8DwlfdBmiCDtrgFYYcq
fbOxMRWjUFXETG3LzTyovogHWqeJw3pQP6VUxRPRC7w5wq76F4FmD/sD+IDsrfAZ
ErRrnD/80rjf+uKKZjDDz3VEQ9UZuJbMvzAbrwD2mnJPRDwf/Npm6hDNnnOg0wXf
XJwGkv1Hwqko/deD4owp1eaW8Y8kcDGuK3nLHY0Jj75TA2wJQJDcotYB40ALT8WY
589AsPeCJ16e4wRkaq38D7NDerX4QUSh8ceJjt3dVRLztlGpiTWY9tboqmyygcmi
x5CGMmOwBoEvBqtRb4/PFlenkz7QxunjbYkVmXG+Du8LnUQMuPFMf4R1D5I9L18v
OMJyMZpBUL1CnLHkjrahRE4fYSh6NqiEpFFYGbuEHYJOUwyWJyRDYvVN9iuq/M6y
UO7+l7Ss8y92a5i7io8eTD2/ZL6vPB/fvW5Y7H+S+7ZLaa/ojRiJV8YS9PQVR9O7
7PZCduddRMAZ0EiCvECG/97/gjgJE76WnKClujE0KS7jpXG7wXaQRHvP1MnhcET0
b3UohGgsQFVZhYViePT5or8xA/DDCyT/7ICoFJZEr250Ndr1caxsEN5DlvI0OIhT
hFcBR76J3/JlnVLfV6LxkqNMHxuUB0sqP20zS/0WIc7Vie89489SCyA3bH3/vC1S
x4kWJ6WU8zQx1bnNAq/kJEx06pnrnd75MQLWYv4Ijg860YmsGs/UBpd4owtLNdaM
Vx3FfYh9kXTPB0MZ9BO7QL6oTsgZX/B9QPS4BZy2ahE+GunEIpfN5x7hcUpRKZJH
RtCnvd2PCAhQMfAY7/cqsqojyZfPrQ6xNihbWrTEKlAJUggJnzqsBkQ02ZM5IqWr
+2qKvI/f99pfNmpHOt4BvRVDJCaR3suNTF6SmsyLHC5ApZwc4xsFk+oaeS632hUU
efHge26JHYS4PUMdG+dZL5ubZfKz38N0G07f/BmR5ab2jnGmRl0GjMGI6pwsQm6I
AxIyySgT0w+V05tUJoYPyQ0MaBSN7L38DoHAO6oAPcv8480Sj88hFXTrQCc3sdbK
66SPPZoZavLT+jGfqB/W34cMTDnPm0KBCMM3x6Wv9Zctyo806Jf5Lb6uj/bCQh2Z
kab89aIiisRTG5kM5VJKbGIKNDtbFDLFmGcHcsIJQT96iUTcJdQjDIBbISURFnR/
XzTAQLLTN9jpIacwELJOaeZbfey++zXeos+LkwcTu3ObF7uD18qiQb8rAM2Pmymn
poRq2Rb7aWwiegoiIJwERWG7SJ5X9w+M+yKObdLUxZMrPU0HSndE1NqTMDiOzLFL
RMOqTKuTa+0lCMj1hYjfscgfJHHhFEg56wF7gQs25MclY4u1wl5BeTl2s2JGbRP+
KZdSOLov5MI1N29wNHvq0kkjcr4Z0hzeUCVgkPjebXYmZwdx7vIWc7Y8QQVRDltP
ynarD9k3MH8Oyq1QffDjjd31GGB7TLoJ2SL/XBD+Meuhc0Ko0aSKMGWGxjrWvHdH
n1PAo0WElnWvUF6Od5egIBTTm/Ww97+EInX+WBNp5df4aHayRDF7UnRKkshqZpSM
ZWI5aFZ5UR9O7605rMmTGnnq4A3/wh+EnIrP/QON3xb3gKBVGbvtfhAwBLE+V00g
vxi9xI9gR6uNg7yNLtMP3Mb+JYgaG7eszCLu6mumaePibDmu2UUsIjKdH2iUl0GH
vpXj2b/Yhjoq+7tSZ31ufz8R1C1sCsN59+RFrrl8QyydsoH142jrm+DOAStQj72E
CbgTf85LHRpo/RpgymHXjJdLRXu1/Db3oc+JgmjquAsYsSDnTbTfrZjTJ46J/lwT
71YmqAnUf3hw/8/8AXvZBYgmRKbWXE8GRrIy4y+l2bb93gzsVbjoT2Y4/PMal/+p
fuAmBY0XAprha1vWuZezibG+AKac3AVgVIZ7G4p1MgwQl/ix24wRVPQti1ja7LZ9
4VU4ZDKPNJdfFFey8uWlLxMYP7pl1p1tXJa6pbiRLtk2uUztENQOxl4LdO/c2AUx
WLHyvhpEaG8M4WDkA7frbhHuy1XBlOsf1YMkZkcPdfCwuET+cjt7w1Z0GJVL1ABb
A21cz9ObkYIxCcjN+O6dyfLYGNgNq39O2wM+FdfY/uojFHGwOVvxxQEVaPtAHT3D
Z9LBZY0rMijkYf41RXHBCnlcmt+DGfdN62ozAv5N90EiOjzWoJgxL8eCrjMXVtxq
obUwVZ1rmOomhromEtH83uWBVO3Ov9rDIQc+kBJhp+mbx6ULHm1V4p0dfdEuRh3r
r7ngmfay5SQEKfbmSdu4nwYvqTzKkXEjUlhAToT93oYcEYxlXRaw5XvtAIdqrqXq
XLX3AeSUJkCWxJNr4dDMb5kPHrXcQKP5n8ZWImbE5y1W5BpHPubC2xQavOhiU9dA
0drBoRBBK4Syx4B00T02D3dkWKzeGEdo+8VWWjndRiPF0L1RjuTigm4zneDlGkFt
31NmehuRZ4lpjATgnL9JLgNpjupMo3w2tbxTLBprNWFrjLDHA+P5umZunprU6iKk
RTGx6tfUQgO0TPnVQEWTzCByvZ9Oi45gto/EUN5m0WwuOd7Zn12VlAChkIx804u7
Z2nWzFBn7btHR7jKxAI6mBzNDJRXJsAkFGczup5A4sTKAcwCuzGBSHIMiCKtX+j7
EoTxelUOV311anJkSpGaginLqjwWAGxV2Ah54OgOZMdmho2BMSc26IfJP+lJQdDv
3MfCgtzv6HP4Tgg/fyg0wijEEQKUaPy96LSBxlZ4dgGCj+8xL1I/lciGQ2njamzB
PR1b8BR8cInVfE9CJwliiSG+CNN4mEInp17ew57fWGdagvLYfgvZ3/p01f89K/C3
GQzubDmiIudOdgtI0Y+kSt5tfmySutGg0i9dfAKTJ7Ic83wcvPWv+DWBAlcKut3R
mvvbp1An8k0FycizJU5rtNu/bjUIoDOc2zai12WimtVB3Clysqr3Q+kq6gTNhuvs
ZfbT1/hOlj56yW2ndUaBUgNHHex3Q/sQ1Yuz5ONsbOgmX3+CbLwhTNZvSdVu9twS
NM/ujnWcY6uQBGbuwFkDqM/npyuF9Ied3npTe0fQRlWRByfYbFpqeuneM6YBlD+h
fPOw9/41LrNvCMyHbzSt+irOZCv7/rUBQYI/KzZ5UbQHBFBIMte6FMJYco0sQ57l
z1/MwKlSEO8zIDtlqOJLtc0mkD34/d8YaiLH5SxXHeIB0tfSS0NxzMNrrA9jEiI4
5MMUOF0UcFAJeIan8g5B1tC8NmPfd9P4cRNySIICWwDtSDuSQjv1BYI7+NdZ32Eg
OMnT8kYsDaK+oVCDdL97/B4n53WsCKRz4oJ0XKF5tulJixgO0TlZnHq6EG7VqB3V
qBAuxFQsQ5jhqTceskFlhxHCdeIVRmf8qADfElUcr8dNeK43ccRFRbVhtpchCdvu
iGQElB9zu8UeOLB5lF3F6JyPrDqJ1A9sS/Ldnps+z/nlRqYNEfHcOZYQeUgV9qsM
IGDVqCENceYvRoypmlEr0iEK2ITiWSVM9HpLHGdMCkgFW5Ri2on2iXRHNlntGtVt
W0riMK5GWrhIs9j60rGiInSM1KGY/nWpeXVwQh2sq9gz2YJIqIr2LdJTUG+AZWRz
KjWlOxIvw7O0otiJKnubXSSB0MMuTTOk4T60rNKEvW1CVXnai5DAQnzFhA/WczUO
aGENoAwcc8QX9rl/mtkxW6EvMMbM2N6T11oPSBmszH8pg/1zvaRYJm3T1M75Hhjv
vr4VBpf+ONk93nNTsOvD2hgnyIPPjwwt3MYWvgVQn4bWI5z27SPddUjIRbrl3Wqd
bp1OgXKgFU2TpjXNfDJV/NlSw8umTKWJ1H2/FM3HffdZfRb/Pzs5wepJ7Pwng+ok
UL9QtJbavzOaZx5E1mR7Xo9RwXDKgRyp5x8vFS/lyVghfLSxVG/Q+cPe3mBGnFGm
nHfZ63DtTw5zNB2/yN6JK0gHQ9br2UujXLeiCnOZmv9ePAJCKUozB01pmTAPbrmr
69HPb0EO9NTUxegWj7CpR3yBiUqbxqesQSa6gwLzJZJFz0pqmHuOZFPn+6yvNT1O
EoLwul+2ld+ZC0LQqP/ChEEQa4ny37uySJ7u2abevF4WaqOoKkwHqpaca5w9RYBX
ZL79+qP03OUb6nhIGUHyiJGuXyWy5mQ1xjnpTWKkotHwDhZgNxGLW2AJ0PQKSn6N
4C1JmCQwWK58GO7dW5D7iUaa2ry6Eku8Hizp9vrv5LRIrO+yITaEOXdgg/mR1zIt
/sigVQ79qMzhzO8RYJQlXlvga9QtPxQv9S8o8Z9j7Eqau0BpsDsaQWnP3jnqojvK
Ov7ixCXldDi3X9F9aBlNRYgnwd38jTh1OZEggXGv1UIxd2AT9WfdS4CFClu43cHY
PmQhD7U3JL41bXFe4f0/TnZlyD4zPiiy4xEZIXPC14Oovta5TpckyZYZkuV1OUF0
iXrbvZsBU63glIM2YLO6phNAgiSpEJbk1/xAiKVjXk5u7OZQ4+s+JmfsOK2wZhZ1
4Oi31BeqQNlzbSclsPlErrG41RrajvhzYoStSP6FmaeAq8i0yG2zjuMUVVJahu3d
rDeyN3hlF1O+6WuqLjwDXiEPV0ebVnl49toCD6Pl4q7dUwRu9ZiCX8ARz0nkYJmn
v05QIRZfMxKN+L+G+JmV4MuGLYLLqGK3/c5iMhVlnVxfWDgIsmAoad35CLZjYhP3
JXrharJS2bgCoCon17y7D4Jpb1wLF+aO+Y2+ZA7DVtslyZ54cA5z9Xdhib6tCW9G
ylEkZUfZWwg3iwuc40O7Sqk6gTnJsIi+AnRfbO8beHUPKWE9cHka0bGm/3kc0K45
x5Zq267X2yYzWlhVvM3TZPfc8EGMW3IbcGpIb3BsdXoXvXf79dJT1iiKL4jVQl+W
NNuXEORFDNNd0lQWYgn+U+Qykc0fQnhLoE4hu2Q7LYcbdn4VVEx9yb7ViS3xe/3x
1juMawKgBzpdMfbudEcl5uqdx73Jaip1sNHm4CPwX6BpqZP6gllIlH7Y3fGOT5P6
As1kcDnywLNh0svs/HpJ95/ohMeMbC1rPCnadG/UADrBikZ5bPuArc0Ccd91MRMf
sp4NetJZlDe3qXcYob21+Ljq5BJ94tDegwLjmg+w3C6zwCDocSTuLa/ISsHCIrkT
MHKZuZLDHPAEvv9SmiN625fhWEsEibVcijiaDlJbe6vHwbFwikGPFCsikPshi1GF
A2BvvDJoU2kHXf5hVLBYOPawc3c6wpmLoM1ZGBpfRsTh6Z42cJ7XfX38zz/MQyjo
hBXaoxMHG9FpA5SLgBI3lMPPyOeUqSm21TIeJrlOOjuc8CSnRD9B7H+HSh6rzEjL
bjomxvwT05LNXlQhvKpP36gU0uWGQ6tTo07apJEfzRjKQApNrn8wNSph4YcQA/HV
yWQO0hqPuw+2xVpE2zGfKyeYmjOj3fhUQdPGRN14oQ1OM8FnJ2r4ArpkUBX+FbKf
OlFV0B7cgPiB7KIJeNpado9KIrlALmIDUhv92Ty14+9IhROmRRDmAia3RZjNmlyB
5fy8ZHXZIlc6JZaVOkjuo19EagiXYpBKh4BNpBaCQXSj11lLEPb56nKpnU/PEGc1
VWhBuOsjTXhK/3r51sB7/DXiUcSiXyL8EbDUCMq6otb1MOmoO2QU4YDKd+JzEWI2
ONACQMA7PNZv3fqGM4Z3sAOTBdlcgEdEEhu+1r1+QNrYm+lsjczQVxB81ScW79Ua
pchRW2aqoI6TH/4iOmSwjVzFJCvP85z/pnYQv4Saxepn6RZvq4DJQOFAullqxrGb
8OhqXyr050QB8DSUgCKGWZTvCQo/XzofMmum3lXcB5eDikKfDnn5aipOJYCvXzoI
TiZx0a0HYGoN3tHn/bafYksxmJwCe4ChOtoPYWfSxUw=
`protect END_PROTECTED
