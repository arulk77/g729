`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMPON25W072Vw59wLqJKQ2plN84bqch5z9HAYIMViQVL
7RtwqdC2A5mKdwPYhy5UOEiGFoQGR02HwFd5eUNUHrAr4eNFn+VyHRrVCV/sv2LM
rFEB5k/FXtN2xn4kBfPXUNF4nIeOEzZyX2MVzA6fR7uAyhEf81jU2aghuGJGOOm2
ckuZ4HTqm0nNFz+eK/aojxTuZXsMPuirQ5MpsCPYKDJWfjqzHFugHnDpHP61RHZz
`protect END_PROTECTED
