`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
WIh6XhPIt7tknXf9QUqbT8vUX5nxInRB47mzt8DxvNE5PSPBB6nXE8M42vCnTISE
33hqYy2nQGYBucglKCFXvIfEatz7j8vEJs8rD+dZGe97tX1Y6lcouWcALGx0IUI9
uvSK1T58J4AJGvkegmZXgv8kFD3k7yi45zh6ytmEZ72CIZaGbY0FPoWl64ktXUwO
guFHHjjXXKNO4J3rFZ0GcIA8xO4iEdYTBVt63y4iZ9QoSA2YXXr34QT4OL/aFV0n
FS6Qvjvm0XLanh5ZQTxuPDpkT++VvaX7CpdPQN1LBGD1qQPNJCg/nCb3Qgh/r37U
P9tOGsbJlsu7Paz280kq3sTSzQP1pNnVM3or+VfScbNjAAdeVYQNq/L/7SnnwNz8
OPnhyJ/ZqNBSb/HzPa8r1RP/0nXHyqSLHldteNAhObcUHqL41ssKZOvIcPHTdW3N
MS1uNbq1XETC3dJ/tOFnxD9zhP6Ds+6bZ0zzmWWoq2lJ+UER/TkURAUWmbuqkegx
acNfrWZvwO0TtR+4YhG1ZOdX2GFn8+HZLc9yMxeWQNikp8JSRgnXFp+G2nszkXxg
UXSam3eC37KhfxLXBRMHA//1WK0IMFo40XHdLnlC3eIeoFm85HT8SXPgYEFoDNIM
JIrZk3ajqXOu1hwCqokMbIgCRhVBzEFcjLYWlG0o2mOcGmLa5Pm9doTwOoApfs5O
jUPeObJQ9mlDwj+QESQ9i+9UExAtIEWBz1BIJ0PpVlQ2Hh2bnUnd7X6XsJaczITA
tk8Ll/cEyrbGmXC67jV0BRfled7M3lO+smHpIpF8qLNpFeINdiFrXvQC+jori1nO
hc7hyWAYEPHiYAK4kaa8xwOS17M1kpZ8YgNza9UpGrmEwk0pXeywYC0FLh8ur3yz
9dnDZdgllBJ94+JLMOJOB1DJTrseAfh5fb3R9eQc8I7Yd+FZZlG0R0jo+5L/+mKR
RuxFjsicjbvujPveipQkkU4H545DfmQamLHOa6mKICC2y7swztx6Cd8QCOf/tKI3
+ArCmRt4s+u9Xr2xfZpGy4OJkLn9Auu9kdnzaUbavGp9du0k5g0m8p69cdi/0seE
lj7YLfKeXwwAbrOTc/he797Ystj0e40cu65yyxTYdb2gP7vfMkIPcEH+2kjjzG9j
gh0RNTUmpMmFsR6yklCeHuP+MiRmPrD0HAa9/mNiPCC+T+7WKKnGTZxiyTfAxjlr
uVxS0Ngo6U81EaZrh6h8tUEMAWh9m2VS/jqe8X5GQQaIf3QyNb5ScWIKu4BXY+yb
596ModzdEPAd5N2NbHejM8quf2YC2qjBC+KaMk0c6eDKddlzpzNfjjQLBOpcRvF0
lX2Ez0b4MeT78TPNkW1pEULoTKI0cdnRGP4maUkpnSZ03c9cPCu21f4YBr3stXid
2LyLcka5lxtYop8RfhHdmLmbfz1zU/ftxO6lTq5e37I4AvPZyZEBY9UXGb87Kw/v
jY+6wIJY8J6JRaABLQL1Amav5DsSHhKGEolutoplw833g3qD3o6dZERuWLvBo8jf
q9wpSI/sa4YCYXBy6/2qaOaF0MmY/TIveMWy+iizrsioLmKy1W2BtRVlSQ+18udJ
Qe1NvLiPiKJl6rKVBzHqJUtyFqC4IMP/r7dBvvBaghRaTJI8TjFIyqpoEq2vZkpY
7ZFehhaeOWNMNtUmFoTbcj7McV687RRjidBuY+rtG4JiFWP9X+u7t4nRXJjvIlVO
yrPppLGyGg722zuliHgKQdUgf6XZRQ6ZFPoxkvP2D4qf3Tl2HTgHbZ+ux4myJATI
LmM1kYkf+AjBjYBn5hJqeDl4F/dSOt4KLMjnhrN4jUc1NMj2Qt/caJV2OvBWVNRS
V1iZJ1vtfLZmwrGNn+y+5Rg+I8984vGdqrTzUYmFTApZJ3J9CQNCmZX+nWe8QPKN
0KTW91xDGkXFY8B0EnN/u4Hdb1xM9aV4ih9s9vYG4iaJzZJ4fNpNipM7qD7voL5+
l5ewxs1UZopI2zGvILOfZvJQRX2Tus5Tq2/tntTsO7WdGGGi/GuROGCYMLeeORb6
8xVayJFK0D6HCn50GedIyCagX5iPganghjDdfAq2rKDw52Emz5njgC9vZqoPe4F+
O3+TSs07ieUtAtjCrTG3DA7qGs7gSiBf2o7eQs9PO8i8uFWf24xcCklLOOB494vn
zHhuW4oBRgVM+Vc79QBhjy6kMcIjCN1QEyQCy1Eexe+pyBVRDeYuSPeRxzkgklDs
GGKxWyeotivu96geqSV/57C+6+JrYTXY8xnUSOHEz0SFVxMaYxraq+4Qq41JgEQz
hKyfYKbdBRTNI+fAKSSx/Xd66Pw/V+CCLueqXYp6nADbgIUKzCLLtZvf6uTU2Dvt
g6sYeIjVLS2140746A0kmhEKh3a+IIFwngxVL083DwN2uXxgPwxvCmN/cxSJ6Uxw
Mut35JdWGTfWWrYzwdLHLhWjRaf9eKDdCHcJu3HA4DBHHK+haXm2JJkAPdtpDQ5i
G1NRRFiQl5GNDhOmsEOX8HgebW0sG853k6/bueXHw6ws13fEwO0GNnL/TlYux0U3
h8LZx/LR1qZ2tj+Ift1hftMsN93QWcHyNxr9cS81M65IWNaQu5YYttrD4P1OxiSG
rJVA0NLQCiKxq0kL0TxgKLYvHfJygcXA9J+opLDwdWEXQBMTgevI7W1cEmdJV2rc
9q07amWOC21Fr49SVewe/JWzgL2Dh7K7Xzy76zW9zHPxMltX2ddDOqvqeQ/WLJnv
c61Q0hZcWJL4pNNJ1UTj77YG57UwwLHvSHnqB1fvlWKLmxxI2w7IELtiLQnuDc87
b/FMmhF3wO601vgcQlxp7MBMr9dNmkYfK8WBvlsKlfu71preGKegBcpODVefhww3
ceZZ3K7peMYVbfEgB92WdIVtI2dBorwkgTEcod5heCXAXmGJSCCSMy2xduEv2vDF
x2LwcilD/3jN+g91NVbkl3e5W/f6GLarfC1bmDF3uIYUCAfcXlSKM7c1553vbhEt
q9Hlp6ISPmsVJG1xYakOGXe/G1cTjAll7ZvCcLdtkR8vVRpDIrZBv9c4fR0/MGE7
aNzs8Xccw8ID6DszRWUwL33Jbr292p5IWABqZxNwa5G64fH1y8JtXOJC9lgl3ir0
WDN3pQ2uu31S84TTX0VKB6A/6f6VQFmtwv/gD64AzcMjlSddNpJsXQYcT7tnlxBe
+4ottTrbSKEV4SUUTlDs8poMiDJMPcYJj82Z/Vt0ramgCeXxQVIBDosNAwLZaNBd
eDF3pvz06RSsXoBxH80F32nv19e+fbta2qeKnReMUBfo78Pi4PabsWZS+wDBxy7P
tZpaespaZ0yKJwqgl8ENnSWrcoe1pTqYlhT5kj/m3nAe6W+Mk5GlmTeIpiBm4YJ+
sQZbSZFcR1iXTgW4VrSqGcsD177DZEospK3gwMt+Y/czTHKUGlqiI706BvDSydt+
CRRMnX8qc9ooC+Ay+MPHMakp6ByYvzJiZqnNvhGIPAYTrgJ6KMFoqqjoPV8ynqig
iyry2DccBOF8CdDMFp947Sznho6G6AV6u1LTsr8HwOUyOILdrVRqhsxMnKu4UuJt
aX10nchSPiyfrU18xX2AHqCk+M721OGs00bxUQUZO4FvHPk1/ljPOg+hvPIb6HsA
ZIK8GK6eOmfQDdX3f6ZIspEohf1Hblrm8rDXBL6mSaQjvsJwwhpz1CQTOSi9f+WZ
3ru82hcZT7XeYay8FrlURZGT6Vok2eLpmqVCt4f7OOXseq4+YdHVWRvLzskOgzaS
PbCmvXluG2mYm5JKhQO8TFWeWDYwigg63bxIjDRyBMe7xuo3RXJwabdAVHU4wG8+
8LvewpzcnTm9UGEDZAktqXuwSeHic12Se3MPIts6IDfLUYeg5Vpc1ih4LQL7TGiU
gX6/jPLe+f+oOzzVG3SFF6Bufq8BiTVJn5j6zRep8h7vAQnYoL7lP0P8CqNl+kVv
eg/bwfLx2EwO0Uv4H7K7C/bImF2nkPjG7DgJdTxCaPdnOxzLHUHxrw19U7RP6TxX
Q/JjwUV//k1d8KO2WDpM7YVYfTiG5CWpxATrHc9M7gywT40MwXX4Tb7SxPba/EXG
GuvIbPO9n/zBmBDKHfkE7guoaMBplHcAjyJZItfVVK101wkx3gXFkLZIv85Z71f7
EgosKVwW4ua5Ea9oXs6W66QpG1iIza4c1zpiCESll73PIfIuu5UC/wc1nXjHNM9R
q/II/mQRHK9wDRGFzFppYsMQ7Y3vbh7MnPoQYy2wvUSmclbLfn0SygIMcTnuTZXs
hmU+/oGnto5iGfvr4jArRvxaGvv4+/bMj5mZHuUzkEYF4uWFgqQCaOunQSTj5bjn
H0D9czdiNQKsS81+oAw5L842vK9T7cLj9xTGmveEsqWICOu/hCJo5t4o0wV+MNDb
+LYOQlxbyZF5uFCJoofB9hvxUHLkVdrqUoWr9GeZFifEx144mBIh1d0Ytw+magP9
kgl89EYEo5CA26CE0JidDi6wUAzVcg+ggrnk+da6TIaSNxr7g1v0kqbC0qrWUwAa
FqjdFIjGifqIWiZnlqcQK8+C3s69fJbRBSOyL4PyyltqYZmsAiawTFDUERpfTJRf
SrM5UyVxA0TT26AbTSH8VnhOFHMmpYrwtjysOBdsRG8fXU2qgNVWKyVIVSucnALC
FdLGP8NY0IPMWnqPaWRmnufskjquwYTHY/a4m8FYNDzSW6hdL4Aqd8cov5Nh/54D
ipTptXp7Z3wJXeFQz1UEEgllooTVZvT2xioSfx5Rn0dY7B2QRb8FZtjzcbO8H38Q
F57UjgSslpY+gJGNpE9Bivi7dY9wx252bQwqDo+PtiFroRr5S+JZXSo1LsHQuDCT
z2/r/ZqtjfEiUleKd7kDuE89OhRSWi5yqFusOob14I20yaogy7N8ZL6/zJQ5lplD
BtHov0nMAeX9A7aNfRqzYrruubKbJ0DvQEgl79s4Yt5/6eAQzIcKSDaKEr2A5593
Je28csOsYKliXHAu4Tszq2qhW2vK4M4oGjD5wgaEZAO19O/qQTrky9pEUkEDtzK+
PuPtOuAw9+fQnzF4v40A9Me87IEHJFyy6Phj3e+kSYefwM3aNzPjMoIA/GpXQehB
gyNrn9zThWXMV7L8gL4Ydh2fwb5blkwk48cwTokKXAfzQyjLu44PDSP/VzFnAgyJ
NI8P6W574bJbmJ8wB2NMm8dcg3wwHIFVRNsnxlL2iB/n8ekCDpwwDWdutJcegKml
vuLzDCCwEHyrnNVjkCW8drLPaM/HmLeaCYgaVLfSp/K49A9chVqE3fyXEb68MAmf
jmvNLRkShdOsXzdoDnt/OpqJg6HmEQKko/iZf/pmBaAxz/0jOqEZf6XC363uGyrx
d5mhcbY/Y45K4X9lTbuQeJ/C0UgaZl4wPH226dzz0mlNqM2cWZGRNc41vJLNiOuN
6s5dGWB64tSM1W6bXO9Katopem05KmcHA7EThrU5RqV48WqFfso+55YKDFEw2MVr
rKj3E3BVB9QDAJYkNjAem2zzVvJ1Q3nw1atujqYVNjpbKIMkJBjz0iBE9iETxVr/
JUPWwepFjCgGB6vUbTBEGEjl5eINAuMDzyKWjoixdZ71VGSowGs0IwCXwvJvb3zS
CI+8iXJUIy3Ip4bwPky4aJUP0S+aPCkUcsplo/wqIhTnPjJZ7T6DdVuiaBWNT7lZ
nGGS71eBYPTOTSW0DlAHXtd+zgzA5efvNhu/h7RhHZyQoNXKVYILRMZ0UYEXa8DG
+LYktp+kxD8BuPsEikOOkGF89ojsX50Df++JRN5YA8fxAEpQPwny0xBBd9/sKqy6
SBwbKbz5mqlACt41xzU5djP0bog86yaEn1BrVd2MF+kPF+oD7jOt6n8o35r9Q/dB
koxT5Y6YI4pzwgKRR7FI2HRPgy+iIXhCeGG8xABc9kdFhhx+c9wf6nLIfvIqd2Lb
bcUpwKBTpZyFEpf450WHHHSn3CayC5OvD4YZQr0qQoFxqxm8ILiXfgGcXm02SeHY
v/lS6hJZ1oqdtX3REsXTXzTTdkv5pahsWaCEKVVF70OWOoAoGnP2kQnW489jTT5j
Ui4clzPq6alHlTu8be2F0UjiyAzmQgHs1isL0eRRWL2wn6/yDEydToX01Pw3yR5N
cx+3ealeom2bqzrd5J7iagvGOsKN7S3jsQbOrlT7w0vVO+2QIH136kPfyb3wbjOm
hXh83w6otZKIN9s4hRBQKj7BBPNL93m00hkxIklpCPv6TL7GOna0IjYF3LzG3G9a
QosoiJcyLPnsn+qR8XOxYxYZHrNaLz7pOYUvJ4Nw1F7sZPDKPJbile7kkyDaXcfi
V3HPjrKPN3ARGL0w2W9F37IanQH1XgV4RRwb8K3umYbCN1AhybIEdmR/qbNTQ0OM
UklRdUz/O17GdC25iqvLM6iRI5iItgH80EuTsiYlcff4o35ePal5twlWcCqjUb1V
WQVMvjKrsaNHqzfsuOZ3dbWc0+tt5Pbk9UdPKZL3hd2kN1NvKICtinlaha6Oxtdy
HSPepcY6C5PvsGvln5fK9onyxvif1Su72hT4OSdY7v0QBjx05R89OmB/aT+yJxk5
YMlHtpbtX9xzLDqWSmTEJ8yDpTXmWDdtqGBqGcJ/syN3fv9xUMa/cmVvJWbCYySQ
sNKgVpowWD+BsfUCAdfwPkYK0LsGqJTfEMXDmKpL5H1sK/018N7w+kJlqtSm69n2
JrBZ1clTnsTnIzV5Dj/hsUUcPDhEHskkLv2ikvAPnYvScsiSfrrJqB0G/7uBRn0v
+M50yMJsX9/YCmwa5RtuoCyrs4j6olH1OeuY+eZ72PDNAiKHZUhLjP5X4XPHoSBj
2dLnkWyfWSJfqPo0ky6Wju/Dx2sk3fsPNv1hNuT7OBxdTKzAzbja7KNpbvnuoaoT
iA7R2VaB44M/yB+4p7RR6OumT1d0D3ZkTfxjmygfIJYoZ25MdT9CsMI5hec13mSo
ECPNnslWpfyvc/EAbFHOUnUYIMGUOU1MSKgz4EEvXe6g/XDR2DDcJ1rbvwmq8Zp6
TZoiVdrZzQhhzCvmwD9M57DtqVm//d1dubC0NhHBrNZx791pC4IYgTKQClrCR+Jt
zFPaLjH0hCibieu6+mlUGYHaHE51YGGxI9undHuH9zyatU9g8+1ppGTrFEtbpQUL
WTXXcBKWVRmLo13FoM/DmFudMlZjKJk2g6U+oii1iH7usjZyCH0TX2aYm7W0DSCm
12DJoDgg8s/IujWYWF3QmHmzhSN6Wa/CzeryfnQPKNXzNnbcme+byxF1/788T9lW
D5vA4oZYxjlXvu69eg/KnG5owkneB2YJIAFIyumxGyRnL4fYydYjTvc4Cmux71uU
/cD2GYvCsR+aK4qWHxt1ICHp6NUFBssZDvVkuFj3BsKqdba9pIf0DvNAQiTNEo3m
v0z380eUCtz3DJXCRSUo8fy+YS6P/52mVl9JlrIli8FSTJ11J87CV7+3Jr1jHLl+
p2NOwk8AiJpVVPdiOfbM/JiZjGpRcEKbNdaMXZUSShyRK0l1/UEaUotqzoE1tzeg
dX/PYTEqnCZVTS901i8RCNs6VkH8XJtiAAPqd5EWl2vhlvh3a1z4yAqaJWer7jx2
kkQF58yHI/oC2XKLF8zWm29++Bh1LuTc039EqgaWSXX6G4Hs3hNwnuOj09yD4oA0
9XPHhMRlNECegSj7WUaTbu7lxY+ba3zo4MNHo2d8rLlsQ0bm1YNqJFMQw5AEcwq1
K0pAwRgdY7uKeHmDAK0zYe3rmGXXH+HiHy8TMXpgc4zpFHCAWtdeKs6wf4KkqTJV
WQamaDtY9piQs2jfCrum2n0O53HgwXnrONMMV1m/ZZ2OZXhMIlZ3RH4zhLr7AxOQ
U820MIf6QH92+IcwRIxIjhUu5ip+5eIuOd/it/hqB+tysW8nEsKQ4Hws2THb96xb
4JRf4LC2Opn2PPb1X3OhVionbNMM2EMpymnyCnM9+NdDGD//PtHrXb0igiGy8BZp
CzwrsGvAgUZT0r/RS5HHqvPg+/9o10D8JevKLDuXgLarIVx+MMidl1OKWYVwYWJM
ynkkgSDxWwbLW7yevhYDicDYOriZBi0iv79u5z70gRMwlMZd04sX7IUIOQwH6PiR
oOvr0x18rIH20A1DW2tikXTs8mOVNez6QHb/5zpC3Q78kFhZFHCPzyMjc/qLHF2o
kfSoUMFzv3X+ia+3mFNRxEzbqcX6bEirMz4RLPiTtO1+zy8v9t4xHhZyPZ3asu0P
oknwtuobIsCWQrux2swfkFS3+VUz9gUXVAa7LWvyGE7rMkxMPQ43XVcppF++DDNI
svc+cT7G8otmbT1rKt36gSVYTs7DUiY+S6yyewZ9jZfySAXYMndzd56QfIy2zCuM
XfcuRTBeBOLTqgnFLjJhFLwEylS/z+3BYdjAm148UypgB3s+LikpPOht+8flp35T
EbmJcWVkRNmC0F2R5ae9972mqW01ORfkQtCdltxoi6+djloCof/qjLr/iA5Btf2i
tlLZKDnPTEjproqpCJzzbqnaUPSfGsI5UcOAI7SsiLPSR4VbOrtCQ/5COhxcTg51
jl4tF5YylyvglgsKvX5OPkCC2VqkxeWI1Vi/q0CSwM2WwQ+s5Ztbb4DN0y1mri2N
mBRNxy/mIwfvBXD5mB+zsGWAMbHn6yBE7lRQieIujDbLefr+6nT3CSWThEtWqT4X
RIGKxe/aXuNUuQ2JKiAiXdN5MZpArJoY0Pip8BvtOCDj5JnKmhfNtaF2+87h1xoH
6Ye3jb0+oMZI0jpt6kvriC+AKvZxhZRwEFLuVFrTFiBLNVml03q+bQKTXG3ouA6A
nheoydjD1Kt5zrvDVm0WKB1muM4gYcUGh0ZLwVMls68MZVjASPAttSW5XtWN3zrV
/6X2UivSjBvDE3L3DSRy2Ia0nYG7DkTgYBtUv73cd+x+wwlnxSFNpgIu65cGK1Pt
31yE7jyDRMcbR2axmRsp+/BgcP6FT6PGHW78a1uK1MDNmcb1DIL8TnH+vvsV1Qk0
BucizO7FIU9iJUYYnIfxT1ud+S/xUvAxiozRDkcPln8pQBV0euYHn2W/mtKh+vg6
kZANRLXnqUxMNvm8s4QP7UGYJ4NsRFCpmzRykR/0Wtfkge4E9MB1nQjU20a3YXYv
lWm4+IpP5BWkf5fl3QP6wCj+mM4qXL0xvJfgEh97lvucM1JlCuW3ixu2SwPN/LiN
BJHTxxEQOKVbKt5zZ2JgF9WasSvJmF1Izk649JSQLsSoYChCuq5QAHBzzWekO4C9
7Z9Gtr+8zoRP84dp+8UePzMBMGGprJGZ9Rb34mPZDJiEeonc50rvVsILp6VYeN4U
4Synct2024x3+cnrln/7ixxN9B01xWCZAzaETZcA/z7mPJPlGuSes8ajTb4m9TzF
bvL1q1YkOZ6ZDcUwFSnLBupunLRP3FlQMHlBzp7SehenFfdqkI1Is9oCfnf/mkpe
9qFWt/r1BwPCHr/nX5vyz+GpbLmfpSnaFUY5BCl7Wt2IhJ29hizrUW8YqwGPWrmv
OCxrNjIpwO7U2jov9Ya7QjMOQguDamswQglS9oJK5Aw0B8kt5zm10Yu0JYx0ORRP
5sO8WEr5ndcWGHKzmN4uExp3K6sS/2MchLz+EAweExXxjLUdq0w5WWvMY0MxNzsj
dCoUSEMYl3PsDvHtSR+J0bzmqRVnfP9lqQ6kLWFvYtNPeRpieDn5qntXu5Z9SCA/
2kBOX5bvseJ4sGFD08cpIddc99TEOVzEjt6PKAat4nu9tfJUULpohrbgEWMPhAHe
OKE8Ow3wrfrtxE7Mh2fXR3tq3ie/qu7VoNcfksL5FycwcX8X0TEQcht9/s+urPda
twcEQ+fh3doqsus8xYAPJ1+fK9OpIx/QXf6+sZJ0g11ngxyOrYMVdHt8p3ROLWwl
SxA1/JGEUDdGcglJFDTPSnfsyZroJ+MHuuXafrjnlX/tL0w+g2NRlycKuamlDhuJ
P3Z3WxfEIzy2NH7SruKqV24u18dyJCoDZRJusesIT3w1YV/8DQdPBGGPNy+etsuL
mBoyqY67OxRFn/f3uzOsI27o0jQdTdFtgTId8UNzDcQ75wup3uJnvcpE0gb2OCUH
vse1/xC65c8yeHjUQK52pqB6PwQ9zgfVCsg+qzp1KWNExOPcQvMcqRSs7JJSxLaQ
JsDx+CUAvg9hc0opvdzJBEBK/LCSprpIu865oQW8o6MDZdRU6tUzjV1BCeQp3uaa
mZ31lc0DfEa3ylO+NBawiXKRI5QfW6TCSOLtl96DvXGwM8aMNs5rgauKyrvTp93+
WivR6bFAsMP57j8o5Z09YanL+GCPlwvr8X0sdjxRT3NSWCFwtNgOaTijMCSoMRhZ
VdN11N4hPd4zleSdtRpfG0h4rS45rJWKE0GvYgLlTfjchfJeb78kcbwOrIQAlTrL
HF1AiutbIEv33nlKnOJ6coZluxqmplWNrQV3tSu9fkCAThRzzfg9JZeFAfo1GHD6
m1MW0sJ5eLlIE6gYcDnMl/xuu0ybqzrWcaOCi21pFF+G5cEJTCT7iWxdfScaylr7
+fbWn1Aj0y9e20G9yRzOA8bpTCwuGZm8v05YRfzSJL0/DxmgciNeOwzI8Grzvxrx
VZsa+lN54kT5HeuTZ4iKcX1T3scbRv28bYVvEXgfZUSnRSggi4MFoconrC8BZqas
/yIEbHAMdmRtOp5BQUg4K9ka8Skp84UAd9XzaWAcOEcsEbUAbbrV3zJUdZHjP+aO
D9CI3Gp7e1gQVAPcsswgf2fBF9LwTJPRJMmG9oS8ZqL0FuFOFPuknc++YBBT0kEL
fvHJgT++oVR2VH2LfYfYaFty94dn42+oAVl3qPekYI/hhBPrVtr8q1OhW7MvoWZG
6ohgpP2Sof4+2nyy4aS5p122fwO5BHHjGhkkDkuHrHu6Rmhd78HIEGUCnW3sCcsN
y/Ih9oGR3Je0icLQi+vGnjW/3N2hjiJOk54RMdVWWHtNh0KAQ/UA0kShJcg93b4o
RD38feaP9rOVypwOxfwsMmSMT2wHOZbHAd/wUL2N+LF788x9873LXwVm1eD54MEG
X47RXEQ3PK0D/ahe5E9vvmZo9lBoRuvsaIpXsn7I+EKTVWsu3Ktb8AuxadMwlFh4
DeSueTN50YpFFWNDMf7/4UyUZ28PlZMazXfnZ4eg2nEgFjNo62Ijj1groedRjAfp
y+WhIYSATPM/6jrnullfceHo8+23f2ZI9zSqzn2rcbVQumwtv8vQT5Cp1CoImd8j
32mnsLsBcHcCdc5kydc8ARPQZFLzH13h83rZTl1DRNtGmiAe6amEw7B17UTNm1yP
Gio5mydi9Qn7UhHX3UMiSLxviOYt2+V3Gb8JJmHm6A2HEDPLncpGtfvI56pjq3z2
aFujNWHviDraf76Ue5Em8UAzSaCqx0nYL+m1i5IuvkBqtCrx6J4GbQxE2F/arF5Y
V6rXcyZPI3Mxb3peKfOoKb0pdpR2XZHhfSggwb5ANerUl3GkKBZkIOr3vBGjd9Di
erzCar+PwqW+YPItBCPbml5E2wW/iS7R1nupDzrNgrfb+DT+xiL7yrnu8uzLYqUA
R4SMtoiq84SM8TIZCBt4Q4HB72c1CEGvSrJ30UYAgfdUxTuMxMqIYC7jrv7Iiwg3
3+j3SflcYC/C+okfsOe7UtPH6spuOVulWK4Stdkmi+YLqBzEsjFhbn57AFec/eKW
gBRLhX6gREn8zx11zvgddzGgnKa99ZgCdrDte0zRTOw7xUVj4HCqSfyeyoNMVZM7
5tw6yD6O6wdyf58BsdR1vhsCJM602ko/wvH0e1ES78uwFr0VRg/VA47+Iu8Pw7hh
QSV9wxhyKOBRMtM7+/tqGbJi6oj0lq00+e1Sbv48kNZiW/7XmJG2P9ao2A+Ixa6W
RtsQl2//p4Jlc8lX+ujbmfmeuKijjuaE0HryYXntIcL+uf6zOFd5msSkU/qhXeuC
k2C8NCIkhTaKH64WaihxZmFaRz6Sk+x58vMAVFvq2238XJfI8rXgYscSio9+Zgl5
36ChkZa7jcweeY1t/6zDpMlzPf7zrYHlmn+iUWaFBhRZcIt/wTol5xLINj7Aiikh
TonRdy0p54Fda/zJfe9emJiX8xuqmnrtojj15e0tEEJbf2zBu3ZbZoPm9Sd0ddXT
2YQR7zhYxFop7mEq+IKO0qR9wox4fT4UFe8h6v3fDhCXv5H7y4Zd9fubjIHiqNdm
UxuZKcL4L7zxZt9SRj3EzJVk657U6lZtT8ZIxnf58N0En9P0lRzPZmdTGB0hOaxW
kFbyeXf1Wu0jklDpr/i8QIRK7Cs1tQCBr13jds8XzLu2lx8KnWSbvZbQLjxJxbI/
3xmNElBn0jsHU8CSzXpnXbtkqfAsJ2y/NTocyI8ef35Jm8Rk5bE1epphnSbG1TIb
brpmM6lFGN3g2tsGwxTY4YnrSJqL4mTsgUZ/ki8rC/VsU5ol62wkahGuYd0TxQjA
DMyDGXRFkrfOj2L2ctNry4OXmCh7bMpYbh6QHGzGd4p+wuAZcMDS2LRlqhKvbjcj
947mxiEKGW9bhXC2xGd8u4JrdJNUGTn98JAhw/VwOyMuiKFqb2I8JDOk/HwiokW3
C8u5m1/mQyUoaJR26+uVazce1b/tO1ZbPhNCAFDlYIhPyRF80Pb9zKxs1zyh1MU4
gvSmfzBDt9ocAn9qX2BltAiO3tKIyfDdZsONRLVnqrKToWPFn/i/yTcr6XepNgCX
w4J/P9oiQrLZHy6LIEqzyHhQN6UP+HkDGku+Xi+gbN9TBdGqMOuliFlbb/k7DXrB
dV57aHj1dX88bo2+DHPJA3O3yP1zCTbSH0VsztIolyCjl+6CMtb9Nf3pdaUPfaMf
6CMdB6vUTf9k+p61YQTEL6QOr3deqbRmwLEvZzq6F1tnPu4eXRxUOIlcYt8JZEm7
L85Ver0WQc0atUb7uTmVBzLfXADlkc2yxlz5Z2r0ReM13PekZnT6Z5MHxWxW01fd
mT9TQh5HdqJzNNNSl926Thl/5aTteKaKWGpwIaIdQt0Anbwuj6qx6yVlGz3WLeWb
phJb+9rOz9owbZ9eEUQHjnwVtL03Ogoj+iJqT6NcFr6EIYOX4bnDpdQyYTbv7rb3
8PgoJMgbEB/x3zUUMi3ZfoDa1VEBoh16SaqXcFTIoV/bqPcvAl/VyTXRBC+XmDZU
BXlFVmGRTM++iLz6+3MsvoQ9p/PI+RYV/XooO6oVLmAxvrOk31xC2+5I2Fvto7Cx
1WnCS0T1ath3LYl46yx2apwGT6W2SS/B738313hRSsRyHOUdDLeL6+17jb/JovOy
yqMfHRwkBbZF2v3fQInyIcM5MxFJlKtVJqnMw9vLFXeJvjkYWjB0FyWdzfSyB/q4
0juhBdzjZ9tRmWWLVI50y4POMxNvTE43ZAaHoXdnDVdRcTz7vD4KlfQLAPoppELv
TkUB0aKnv1msj5RREcwV+E27y9rGAy2fyD1GeiHoq4FqmSwVOulAWFHJFunazspu
DOHLrNdhsunnZA2g6QFmwGODbS7A0h7+taPT72KCb2vnCjmSOe1l0m968GJyw4q0
CVx+J+EtqK8L5jyxQ7+qWLDueHKGiBHVG6eYWrjc+KHsAn7t0fVqe68YqWJWun2+
GIGr8Twk9a3cYljnaH6WeyaACU890gjIqX4gsnbfSgxunOKIFWa9Zn6rQlRkINUZ
XskTc7JgjpcHij/MVwfED4oY1ego/oQi3xEODiVftEt/Xw0mTCWPDV3dpXHcr3ZT
LTUW3ba358Q43l7kpfvGt3RuBT3kCyMzWmrRa7H9bLoLNXG/2y9XahwYvFXvsoBM
itQb/QGL4E3HoCT4UnzIjh72Z1Re6rfhWWyP8wB/8ijWC5ywHIZzG4ff5Rtvi05S
OVjq1+DD1bkiwaLd5YevRtsSRmtV27KtavvVYo3FTHo3kOun9MqaCMozuuVDLk0X
7kBTu6F3/kIski4qkVg3TgJpjBQ19R/HmpPc3WbP5DO8EMT+JtNbjC6ZlKCNe0pA
i2+Z1p/nwcipLFjrBci6UA20lFONNP3hTwGG4oE/AHtQyEY4qDcWSms6wAzbLeS2
XpFwBJPFGCSS9yAiBbRnhzAOeVU8Jpt87nHUulrh5YbsDChzgwPmJ2hrMPT9k7FX
cFZCHo2YLFYUQhlrSbARXUSdogktat17f+fGGHIeH0NQ4miblNzZSyREQiJS4koW
BkCTkoJaC20bp4qU4RfunKx9tqfqwMGp3gAuDar8TxWoaNQPsJL6k4mqTaae3w/g
f5LJ0bTUz4MBb52SsdMYamkuOY1xMZu6bnzO/XwJLpveHE4/6Cap1ps7hUgn3+e0
tEJLyVqLAvrfyJ7DmTPeLe0Ab7v4/0ct6tu8sudBqXOURLEMgXNrvQbQkVsDC2GQ
/LMMLXjEB5nql6Bqvizvsl8ylBOlKivPsP9lBo8Oxrnrix42VaLtojBDT3vbaDEd
0wW0aYbl9pro2qSvNU6K0mXMx6aiiABH5cr2Vd2ZWD5g7P9jTuW3BZ9CNoTrD7hc
M2VMjuLpxq5Fsw63Dg/wK+VStdkLfijtxcY2vnUzF+x7/OamH4HSxRlhH26qLYnM
qRVATAqDdHaARlOTtTILt8sMny8Hm6C5ygLWz+e6tFjgltYNKOQd/eHVfMHJCAk+
KO7QuqwrDA7PfbJoQBjUUHMrbeP59MQMj2wpA6wOtoH8K0rusTOg3bxEm0kuAT/X
UToFEA0wzUhfHDNOk6iRNihP1BPgxOxWjnLddRA28eaWz2fAH1TDV7wOsuHBql5Y
PIXAERd7yYttt/SW88nG6SMf98FKkTCIQ/FsALE9XNg1D8vhabreP9asGLQOHXpR
T67A7IqkuigJW3yZvoE9Oj8j24+i727ol3JRMMMxTsLeih8NZoz71xwl+XHwtRHv
xLuCsGjTElEM+Pa82ddXkokrfPomDg1rKbH0jS/lbttKwMayGyVrCXrFm+sb66kG
lE8FMueUXyAytkq2CaZ8Q+AcxBgArTrlkd6tNPBwnB1bggBn7fzkT4FwRZBZODRR
wxcY/sFAkwQ3Pa8KjJMlkRyUPyXGMFapy5/MfrQPv39qsZCXF/yvHLyjZOY0H5NM
mKrOvJWVh90pK6620epfHxGokVYGOVwUGy3+l/Tqek3xEYcMgEBYz641/mmSuvq5
LytCHxZN5MgqxD3HQL3x7+mFbM+h1aZjlPX6ltO79kVSsTnWGto8L2Lm5BnU8nAu
q6jqeBU16PqnkFqoS4zculyYQ9oDKKngpbM/16qmdrbSiuVyR9TRpwkE5PLFDMPq
W3dpPqzAQTgNWNuevXWYGWEHY00kjmtMAUDtX+qrkCgj9mb8cnPk8rCdvWsLTk/V
+GBR+8lT6YX8mt8G0XYj5CkxONDLk90q596s9awioie6wJChN1zWZ5HEximWNz5c
xleCdHsznqWCTj8bKkbpTj/ZUZmeIID2fslR9hasxHXRuV+xlE+xxUBrPCkxKp+b
kVgUliOYIaBrYeW9WqRnUfMgjlfe1XP9KjzEVUe9kUo2gm31BIomIM/sqyg0JZbM
E0ojQX/wtX6YVlLj0yTnat8tL5uy6y1REo9dvpVHqSfqYd24eE5u4NQzISTVxZX7
c4i9B6aIjN1iWJurTcn3+8Fspgo+JekxwyZOrJsF37TEiOQynLwxtDa0s3ivEiS4
M+IA2ISz4YFSUjsugIuySfS1wfCQuc2uJAJ9DYUQ7QM2ImG/wGuxu+uDsIX49Gy+
wSc377pnCIyOmxjgUtvC0bVeYhzW43qPF9OQvswFgrY7EDLBvCEirnE1UUW3A0/E
9rE3fN6EbbCm39R+6xkDiFExSjghFybDVIzxeSJo/lFowa9uwjM2jy+y3Oe7ITqg
G5UKPF0QPhX/CEDsFL0t1OwcBsHueawukBYh0Zl607FB8KItw4znZLUMNIYQSPda
fBKcssAneLSs2akUbp48V3Wgwsf/LZyT5lFrXEyfpNVCThjAbRP1DzW73j/AdVbg
YElfc3o8YHo+QvfRjdBAsICvRA+mPO5YX3iyr8o4inw7tR6ICxhxMpF0J0I1kCo+
H75YALZX4ighmZIvC4eDOvy6MLf9oCyjYJEDiaGJu4HP18xOaPe0aZa1nyIuBjo8
42IKr5UdBppQCZHtQdhjVtNZoxzsxh2EbXso8v05Yh216wvSX6ayT6BMqToTOXhH
2EvcY515gDvIl02Z70kAmusMvlTJhxo/hAG5SUY/hmwfrkoo2iLUqeCJyhbSI0kN
ymyJWaQnHZOmucrN0OT9xgywct+RGg+wMlJRVCBjze3BB7vX1xfn32kCMhEdmvRp
PSjCd9YdP2O2D52LyKEkXfKbgXDllh3yyDmlnItkR4fLTCxaN9yHRSPRMl8110fN
aN3y1UYwKWAuRcZ1MWaBzuafVSZvBQHDjvCopSrAa/sabduzCMGP2L+KmOQTpqde
0GnldxFNapN88gFtYzAtfgk6NrG16VkdM8qMv4gtzi8P8pAP96fC/WLKipFfhL52
OiMGBeoh5p7P24jVTnVWxwy2VAiGHuW3lP9zebwTWO4k4gDfQEC+oDNt7hn+ImbZ
OAaPwRyJPmQ7vp6DIhfXhHEyB31/66Q+F+UA3fd93GQUsaMBpn/vQQzCgb8XDmwr
9n11ZkW4+aiDAw9mNazqCyOr+jNQI2VDJeFyzjOh/FAUSKWIUcAqab0mKrybY0lz
uunMhZVuaq/RkosiE3KQOVbuzblOoYtNfmuOs8MU3iyCesAs2gpJwKezlnf6faBb
Z7If7+s10CpYatAiHXAWGzEov1AHhb0p6zdhqOtyb7+/PEX828XgUSy9hwaoBsPi
EkCxT7tjeQBd0MG4UHuJr5m3LEcHMnFjBHZogcM16crGIpBkMf+Z+MQABc32rwIX
VngfMV5fJHWslgE7wt2LbK5uy8ezbhOA75A323zJ9hTvGFxWxyHIuRK5e6FGp0yi
SfpmXq03Q6fomnmp4qKMUxe+HTWAQj9uOoXwu8yealoblzvBog44kXckx56Z5F+0
VtvTyQ1P5toxwubneBLNAPI4YU1uA7LbIp/+MPVy7wsgxBmi8Z6F/IDaS0cwiHbt
R6c6VyXFqHO8k2ImNZ2iEFvOCAqnUb9TvQrpzpWAAc+x3IlRvzaHJv5tsOzHF0Fu
kH2aiai2Il0t7Zl224uthR+7caWtO5356+gDtXL7Nc07ZAk/rW2A9DNCej4sW/QG
NOPDJsGuxG5K542bp695/xeYcoBwarmZ9tiC7ck5rExJsO6DnNOPHr8v4ZkqA7nD
L0z+y1EBvvGAzb+rxfAIJJptH31fRabljAM4j+RS3HC2tF36zIdUCFO3FiHGvbsv
izh+nJdTZgiKFSJKP5JbZ/LRwldUj+ot8JAk/6gqaSVNtAKSGc21NbH/8faeS0qY
cmuoQHxBQx0AGf+btMaldHCAoxYE/ZuLO3MBR8LESKA=
`protect END_PROTECTED
