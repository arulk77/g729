`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2pjSQMqY4q/kAWGZ4WMpFfDxbuHW5pDz/rr5w4ZVW6ovPlO08nEX316XFfAZeMef
IK16cyKfaVA4+bitcPvgMtk7YmbF6tkC25Px2j6MlCnVUfvQAokEVVplckqAm7Sq
bl0I+Lv6qQqzk9wRi0i7ALEn/UKwOBm0bAHb9C3s+UvlaqmWglgvHjt62ZjQORhV
`protect END_PROTECTED
