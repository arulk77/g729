`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB5QC4McBgvctj15/Vv9delJ7bWrhImJv6v93Fr/iPwh
kMMtLVEWbzCXZW+C85sbgqPRJJtX9LXWnmvUVGMGXONzoyLPBUlmymLJ0Cx/C4PJ
Slgns1MhDlp7Z/0sPmeoJmR4rHjNScaF5at5fM8CeLNGB9pCxax2/Ed9++vB2d9C
erFuMa9w6TPxwnyi02de5vQZObP9fuDtiDQZEmmGWIgACUHw/GhNSoHrZw9npBKC
4QiEaLLvonTJjo1ERxmhiq3/FPA7RJIAB06gT0ycEuH5CjrmtO6YUIMtXBXKpLHV
7kwWpkIQKKYjuUkWr9f0aKS+8ALybXAadGEFYUnnLkQZ/J7fdTnj1cArYtealveS
Z1k+M5rwMO/Zea1E4A8rXOHmtuZxY2tRoL+c2GyXL2lrRo78xc3TCgFIBtI4e9Vm
va4L0TLEVMf83ye+dLS53+glyTAY+mF9ROcqh04u3UVECtr0O/ETNQf+evRIbtY6
IKnkf/Ay/fK/f1tHQG2TmMh3u116sEvSfWIZmwaw++E8MACSaOrKsGv6pDEFDmC4
AZiQ/7ENlCjNYst/yUWjI0nH1gpRJqMXsPhfeWMZclrDolsdOY9XRqwFpGXZDlw2
yL2Y3khBDTxxBnrsG5HdHi56tfn86e0vWSQ/Hd4XjFDIn1ZM9nHvsFPoxc3/3oPe
tSce1WPjGD9xpmMnrdu/7sbJBNwhhiO1a5n4s/6GgzSEsoJR3wuSf/klgS+BYTwZ
LQPnGGFWg4HIXi4R6rbFrJCeXgAw6/HzNaEU8VEUAcFqkL9RLstq6Rh1oPF8D6mN
gtDM0gbJg8w1hKDnZIvbXTkpgE8dbbIBWKDD42i6kZCxeKP8LyWXXUYIvyliJudB
Ux4gvMybos+k3IMxBt8ONkMpEtfVuGPdY6QzZM7Zf/YBSvItOxmNYLDWMnKxPpuu
Ekj0j054uoNZMUPlHp3hhZaO62yiEuv5rFlKKlqYENU=
`protect END_PROTECTED
