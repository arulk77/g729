`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
PfPnoOZ+UatmXSQ1diN2rtBVPvweeodOieXBhm06Xmat5HFYhpPuUUH0/Q/0BKQS
DIDnUpuro2/WVeMcaGXFpqzMLAnNiVnoz7iSkrxa95ZpGSoBSu/Ln9Yc0KwxTF0U
qrYV/Gz4ySpANbxxGDgRKQbhrWEXQBns7lzOuM0Jb8Wlm5O+pPCrMP7m/Pps48wE
owPSUiWS0/xibCCboInan/hp+wCB28Da+kSnjw70D6MKkbfYafeUCt0euFzlesd1
sKtkfPuaP3qCPO8AZbLh6YYAP2eC+aQ9PU/mNkxJF8LuXS414kDNRB73PWRJr+X/
lkx65Mj207D5CpTrtUbngNPvBPi2+j4wYn6p+W+ll1Qa89RwXlvhivdTPrQxPgH4
xvwTm5PYyRXmqyc/LPmZWpNqOGFFfCyfq7ox8Lj3qPasecx6T+ohPCGMo7leQV9x
Qa2LUnu6rmsdW4Me3jIiMoNvkU3ZodXX4gb4AP6g5ZUqbU6bBhuiQNQdIQ2osb3m
fRP0oHfF+c00gPaMKCCRdziOnfGPWUm9W4TIKnHQrUuh2Hz0oJrIt5wohU3c65Dp
EfGyDBiz58OO5xvm0Y3ts6HL/pVlOyFwuB0zqSi250BMYWGHD+TsWYsj893NPkcC
qnKVPHcMeUQmhVW5djtDYCjUU6wLD5mCikLyDf5pL+8+FZS5tnCuSFABa0UcO+zu
hEFR6AfkhhIYrQKv9Or67LBANi97izv04PKac4e8Jwou9ec+KVewTcSs+TYmtPnV
DaXr75fyqx+sc/v0Jnf0QsGkjvYoYWo25TzemFwYdnE/3zY+5r0z5GwXih1ONxua
fmXD0rMS4VWmhMyBZHi+lbTEHrql71HC5dUBu1K9uQmSo8G2eaOWs+iGbKMRurc6
+f0FueINzg8SgCyv1XQblkm/RIWdHn3Bensn2PiKbhuxy20j+d8FwuY4bkgoYrza
rFw0qughmX30EspEVR4iEW7Qfc+7/GWCQuZncWNz70Jw9WIf721U+xAN9HIs+pvh
qVclrYvHjppHZLwkz4t5yg17FVM3F0F07166XOqap/GySb1ef4ssstQXPsN6lyu6
`protect END_PROTECTED
