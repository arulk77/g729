`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
5MEtaEVWosHJcOn4uq0/ZN99CHAF+VkI9Y268IBs5oZYbLsTI0URi6oXeodC73jx
p0zXr16qkw0pS4O3tj5P1sZMwUFX565z0NUabJtFI/RPv8RTrRJ85/6no0HzXt/y
6gSP+Qg+b0sGzj41pAotEsYap8F9gmub6qBJlBY1epJ0ggKn/kkO8DcBGsRso/9k
EjVBcHl8WYEY9Uqg5zmABPv71I5Tf+Qy9iQ648olHkw0PikM3C2rT2YU6YGmJ5Kw
a7W/9JkwJ3VV3hsKcmmfKlF5oOIW552mEOpjZ/LU/6BjgJl0fyIh2+vbnrJSRj4I
PqSxP0zWuabKe2ubO1nRK8lcJShVRaQz67MQdhDDxBg=
`protect END_PROTECTED
