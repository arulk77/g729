`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aQJCjwzLlVo3fYhNmIdHW7VpIMv7jx+2RoEDTgC6jmKP
ay3lKvt7mXwOawBHepOmy4rM9pCNXV1Zi7DxvTxYAaSkM6lLnRPLLgSvhxDDmdnI
XVhRtZ86c4/trEvtSEsLKIIp4hs1gDNyfFljh3mKeZfaFqY9JBLtZwBI6ltBrqv0
GpQlvDhk07dG3DwH2CjafBKpXgF2ZMyahd0T6exV9sxqK9YLjDAUqaWux3m4FGqT
GVQFn3cCBXWgCmPgl574VyZRlkfIFMh0LUTT2ipN2ZQQd5g1R1OmJ6BariMPPiq+
0nec1Zspe755BeKhIB9dDFD4qyo7Hb4cI+KNZ+JSNpQL63Fpwfe5IComxAJb+Xnd
rrXzQtpbaMnG4h7pJMmPChps83qpidyFJ9nfHCyJLRIRAFN7ICvnPZvVBh+UXzyA
FBbW6DGnhSg7A4ZlwpaKIrQqGIgjRwBdQNta5eDwHrOf/7YJz9ndw4ZYmOYOKDyu
Epawf1JWmS/mzXpvjg01SOCXqJhRHjTI3/4ONfHk/15mRH5LJ/CoWFYoQprBOgSD
wsi7gEThRUrjjH6FjWOSd/PLoz079eElY8rPtXXHwH7jz+17D0047aVG2dDrDHdx
4hRbhBlEf0n1ODuc+n8G5sldGcfdHPYoW75yKbZdmcwJPlcM7gAE532QWwPvCWfq
rrn5vM1TbkmSYKijFy16doH9LoXiD36gKbmVpLV+c3pai/QRDOSm2T7AfPitoSz/
Dye7oJliZOhjMZg7/UXVm7Ebu3ZOXmpAAm+cfiruxMCqjMq0M5FnGQTryVQ609gl
NML4AmO7lVjkIDn0NAy+FfGi1yLmiouruzbAn3v3yjKCo1PECiJ12k/8iS9feNmV
jg8kOvvy4IQ2K472zLatvQ4B800ucW/JUwgFxK5zUewq+BT3t8saenN69l7QnlJU
VbUS8NBRgsSGwutE7ePORmpHaVc5kmL4nP5ddcSkWWUbR1tGNVYLzzjEZ+fY69lJ
/cTVrQNbtq6i9IED2l1Owqdn++oBScGrzAyBv12J4ffI0oxv2oeveyIEAkDTJdtY
9CTaFhcFDmN8LkjOpyO+GWpa1D/NEyfww2H4rPbZHZQ/vflb+6GPrAElcNVkn34P
G9TLxpLCqZqTEItLFOyuYJoioASycgdiXTgFJi9xXTm0QMM0GFpq9CYHrV+GvOUi
Vni/vuDaVAl075WjkcJ0q0WwLDiLYDuhHpZt61zfswckK15pIftGZYcHJXbxzjDa
sYNaZz8zUTDfdmcmielHqXFFyHpWaa6ldxyyAdD/ikD2ZX+ysztiDtavlan4g8iL
FfosGLY8kE1rVz3POwOwdCWf/B10Mv42IYxjLenbMFV41z1Vd4yEDtUiJIPm8Pr6
4Nyc4KbOhRoqgcz3LxQfoykk+GWjDTnhcE4BA94iNgWrbf2UnJjtfuVaSOqq0LZO
E/u+y7f3S1xSVF8Muu8B45IetinnQ06w1XBNDmtBhDGZvihKHa2vSY0PnuWNjplp
+nQSL77JlxplSE06QXcSSobyi9mKk6dqs4DN/ajM8JR3JoUH+GVIUNYvZ/SAKbzH
zG1j6xZC2grJLuTqHx/bpirnS9Iezmc1ofQmzQoQSUb50VD9C/YJaVqepFI9X2Uo
lDHVgxuf6jxZ5JdquIY+BJvL8lxWr9ccqTUtc2ya8lubkWz/zRKPbEP+aq63PE6/
/hfAA0qQ4SvlEPaK030pM6/4RpTyxbuB+haZF36KlJMo/IjHWqt3LxRIvOye9ckL
jNMeD8sxzZoFDZl7bhfIXAngtFp7+UbM4XTFOXzegBEiW7whQe1TkiBPqQiZnFFR
FW/uPCCxz+BZumZu6g3pIv0E+KaHH1lSZe9Jsyfd3CQ6khSt+tZERhlCUuVLco1q
VaBlE83cXnyDpvyhc4RsZYWhi/idMn2Yiw4YNS6Dpbii3pEcy4EfGN8La2QLP4Jx
qBN84ARSh3RLMW3At/MPJV73ewfeaz22sFaGa+Kg+lUZTT4yLdg6aSLsQW7HwSD0
zaUIbKXK2xz1zLnWDCQXArZ7kn1qggSGHXbVe9cPDw+nTkGqYis5mx1XmLbJkPz/
ifiHsKxi3VbgOfQdkmPr3A5JSz06yvnO/NhS+JspRlwQ7IJpNhJXsD8iFeOqecq3
jsEcbSmp7SQog1SjDfwPqy7oozmOSSWypeyjCv1N+Yld0JQotZb9nPP7E0OrbzBM
Pzj+bzF38GTJOWgblpPHcuDNZaOIJVVlf52amiMPzo2nGxdAqQd2iO//LQNqmQRo
EXwdbYu2ZGiJkXUz+8GsFXJlXnNAb4hvwz2TLBZxUvs4KYgPq5TRA+WeaQ16JYc1
QGQ2P/bHYwICBk+m5cMjdoZ2KY7WpaVS3s1+tmlsXxyoeBNmby0IQN+4+EosqP01
+94QEcj6PEKECuD/buv9v4w5GuCz5Day5So/VE3VsIfzmSFZA+X9qpTXM8O9WGAf
pivSNu+NCeyFsKSm01G2k9AV9QP0d0x4vYFmwlWgsw/UffzksXqiX2z7Juza06Jx
FYrxXGF/vDR8bNfmxunTrU1n3qpaVSObt2mseZCgJ3BLuJ1YYEVovHqUFmVYMNaJ
dO3cRUGd6iX9yIqM+AskmonES+giRh/IhMxf11kqGP1KKbnmxBaZwxMx4Wpn7FtQ
slhZuGG4fO78AHN0hF1EsTH1PyekSQR5Irmrw3YL3GtOCtai4HwILoBQ6+zoA65B
LFGfFu2tj+nUZhi0Nn7J1WAmq9b2/fGJxtsnJ9i59vUtHNQHEDrNHeawnH27/+iO
6TtkxqYsezGAvqQP96egLaK9sXpBdYBwWzBYUMNF7++D93mqqIAVThWJVtWe7LpN
xQVrZS2JJbQ/Sh1F/WNt21t+KAV7eueMn68y/HKiezVArLfJj6C63gb4vVt5MEDE
0bVUpGrEtiPZkL0saoMw0qFhP0NUmZxUn7iAPOKFGRhcaH6aixQ019Y7V1ByGWfA
PR0Hl3GTfOQzMta1YIlJM5ApPz2su3XRmUgD47WxixXadN7QXXuwtl42rY7iCyWz
FLe+D2kGZJwPdWYELp/H6mjWfC4FkzS3BATOUaR7hmHgkTFu0/rZLiu6bgw9zhfI
2KiKSq9F/b4IsHesujXwRuW3nCUQ8yIth3Dq35nUKxghYy6LQ2k6Yecy3+lYHFp2
GVCSRJhsEQJc0d7yhfztmYrNJ03+/XJXrbj/ljBc808VN36xeA14YJHYAmCM48ka
k3goatOBmUehu+5ZjJEusIIrI6GsGOSyk036Wum72gofqQZkYWJTJ46/sYl9UnHE
5jVQn8ozAaW2rtJ06uXFi01IswZwakLkAmp4lQGxKvoYNp8zpWgoXC8pHeLEh5pw
1T97bXhftl5623Yt9wd2Uczab7V922yL3iO4WLjE2fg9ztbnlvHCPEv4DoJnwqse
hfG31/4jKVChd/83EBB0XV/IhRk7rlWJGxMv+2CR3ZgyAscSBRn9RRruEguHG+kx
KSQ/bBli9zctjUR8jP2Dl1b1TmVOaYnEfRM2wOg1lTXvhLY2XB6PDU77NLVOEifM
l0HuGaL6CowD4Kuxm7xWNKLhyHgJx/5NsLwVs1oNghM2MhzQ+CvG1l2qRf3AfxOQ
9Ir2l+E9AO23xPHDlmdyqMW03iX1qyiWv0c1rRb5iot39y46rxvLk0KSakPGKuIv
+B2mgBkyUohHz4GVetRkjbh2clPsgcqbMJJXTXnu6YpaQuXlfDWgF53QxGq0GKBG
H1xFRrn7+piZFNVwOxlRszo+pVV3ktOMEn1QYD3KYFl2xlozdj5ljs2vxDECLOXj
a5iynm0rU4ahLBFUENsQP6Kx/faJD6eADQ1BK2XpWkUIhnhpCTR8MemVd9J0s+6R
I/8jX4DSvsKn6O6dMpDPoR6XEBPBQYWUjV4SQ89waiOYNU/+Z/fsqSKUqU7Bzdjv
/V/3rDHT8i1ncyO0W+qYw+zlJQ0tG1bhpOJHuDEufm6rWFjj/Q1DP78L5fN+5Fas
GQzDwRlNE3eIV8D30fmt46Kx42SgcxkbiPIslwT2sZHvH+ffDUU4f/OSdeabUxJf
OYMU/zXnd91ucZ8LxB3YL7Uu5DC/1coV3IVAIXjwYpqRfpTq6RH1yoAik5aqU5f3
4brOpC7UuLyugS4QAj17ZwxMBowLHalvWJLFvFaq/iLPRnsVAgR6RUqjA7hWagj5
m2xvP3H/C5G//iFJp8Pos1+ADt4SeGjLk2apz1D4rmWj2jiYt1Fsxoluiwr/t1sF
wdMXzeMHOKB/TP1S69Z65RLvvvcXYtCYqmq2Yi8/ICmUzBwuRaN8GNk+rtw+qJAL
CYB2/HvQSV/ieNy2YAA1iHNWo6cuIBz0UM499ypc+5KBJTUpln02WzzpleE9N11q
Rn9R26/0p/pYa2yAvYz6sCLVnvkSReblklzYDABL6SVvD3Q7FvWsdX12AI0kwAbu
aA90eA5snrEaBeK9x4tJXKYOQY6H2cuMJL1a+J6PGa3LpdE9iVA/Z1eelMXkmF8E
n0icxN2DDGeMwpxu/FTFooDfcctJ3H6frZAXuBlM/YI8V7ks0x2pRqXVFdMYJtJF
K1GQaao+77iu/i+kFqbYbTvrlYEEp8lvU14g3C+Oxe4fU92WzYOglNes5J8hFoow
FNY5y1P0o6jvv2pTzxOoDvCyNQU4D/+g/lTi6jrDyBLkWJZB/QMudnJ6YMCU3rx2
ihe62disqPPHN1jJv9E/OaEtQmUszUu5+eqFKDaPvc1dUK6nNzZwOes2SIGlFz9L
YOQg8kzsKPp5SVKZQoW9NAzJaYzoly9mGjfv7F4WXd4S2hsnr/553JQhjT8GlKAT
EcHKVfY5P+Tma6r0lW0ohQppXlSM0+o3R9gmB3xWuuEMNysFWnxCWOzsvpRkIbPV
6Lm/ENzXFvsidJ1UgisWLIZ6ehkP1pPdiWAQ1KT8zi55mlw4WC+5JNK3fZS2xoty
xLm8HVXjUqvpaBjs+8B8cneyE7TVHgpRXK5wLdhRQQdukJbItP3Is4YvvvNKMetl
rNXJWigmNcz2S3Fxd7zgawHZ79U/ULhj8Vvf+Onz2bCA35LwJtZEZa2r6l7Ld/Xg
fgQrzJFB4g9wi0EMLBrstUpVfT212fzT+uczudZAGV1cuMtoASJXr0OCPG9Bpzwa
E3BKB3UwBmrasWUsyHWtsn7VsvSk9umiAOj1MB+2Jo6l4ul1GCvo7YUYDtgiteg0
qcMdC9SbterYI9zTlczbRpySADFwyS9goo843J6fPWDCj1kUc+d+bYW3c0rYbtw+
LFtbnelk5Suy9GbuEx7eeM7XfTPjRZiLq999M4JX0TU9/Oq4RNhbRiDrNTRBSeMK
G1wK0/JhVtMMkhtnxfa2vk7MfFmGYHj8tKRygnyZtrBMxqI/ru0jv2wt7/79scx5
MBgBbCZ2ighymgiEpnw6VB3nATEBvz4Dmudjs7/jGzo7GGqMZl4VlsdNIX6W52DH
+sQeXa2ROQ7CuTMcvHHdFFPNpdSz/S9TyAfR8VjKWidHGTHWJyvtwJYlNnde9pXe
tUc0Nbq/3Ge0BwJkI9A37gDizm054INnpr/zffcSnnV6aPLaKJ0UKRkNknqt4YSr
/nwlP97/QZh5VJWG2+RwYJv1XKdTbyeM8dMvueMAOl8Ykpq4jHR6LKK8oB5gP4gP
7iMffd2c8HJq8zoK33J/U82RN8VdN6lgP6Tq4zEB+MSCkv7/eywli0sDkYuCSb6r
Uqi87PuoXOsJ/OvVrilSeGbr4fPThgrXb0m/j5gjp+L0r21Znv4GEUMJniQ5An/e
4d2GMh6+jv62h72tULyeq/BxyziI+kAbkbcbU6kzJoag3bdm8laZvAPM6S6rweVe
5A+3rJUIuTD7FOsjlOoNIl8B4NGZYZ3uzdlAWGX4vtE77+WgbuKfJdhDGrtkv++C
hf3H4UdQ/6DeY7xrp/PjaME7kmyzSFAhkWpUAU8JQCV7eG+Heh+liBzEBt1z1CQC
48ae5hkhwoogiSB63vRrORAd1S44LQ4mD+rCZT45ZO2ZMGZdaWwtU6NwvW6hjbF8
2w/pSdaEhrU9aRzYO32cLUGaCpIkl70x51Yrw2BvqzejkwBKTcog6Itia83TI47l
OFWzYpTL0UL7N0VzKYjRbjYpilTcZNsRkclEueMBS/vH28ee5EUx4ip7RK2T+hf5
B9X0ZwU6439ybtvxfaPrxEklmjiDpVyQfYKg8BDnBpuc1rmNILqIIqHEDAIICX+h
NRk7oob/zGepVIE8izC2eiYdcxX8PZkX1JbdtERClGSNhDaWvLw0pgmvV/kw3UvT
JHcazYq54YlNdhhoB8FnWrZ1PiUjTE6w57HlobQekud92wZiUQQWU8Puucqc41CC
vY2htspAviQv/yMITfBY6dTrCyCADBtsopVFQSuwNP3yw2SRI0Mecw/E3JVZgtjB
+Fl7pkuMhqJvSB0ro8comdXpPbbUe7sQntfGq/+UdeJrnjWRNDhNqKJajlO0nKpO
EX1ZZPPzVOs5h0Fdw4ORpP9vmFTPchBPvvRgejdlVH/BucS+KOBL8GbuEK2BBvEj
TFRRynpXw6+MdDD8y+GxleBUcWKFKeo8ad+CCsu+PD0Oiwx0FIbz0B/gzVJC+Jca
s2qGtT6b0HpwX4Lb0wnbaiPWCjAfe9lz8RCpnNBgP/6Is/7unEMO0o7jEPRekYSz
qpw6ZuWs3wboFJOq+M/uzugHxQvMxDoYN6hr/LjOgEkKboV7Eor+9ExczaRaZvlz
uEfqiiPgggw3ycaNlGvVQqDOFI/B/PIQ26gzmYuLNY7bRvewAUJjR5Ndf/KyVUGO
DVPK3e2zAS10C8wvkG0fh8m6ltVwj2R/7378hvu+LRRzcI1fXWx4gHfUZb3o+Hak
hbzemoE0xUe2/OZEETQ6vVyy4LUNWlEOp7uohl2Tn6OFI9scU9+mjb4W85jl3zmf
YJvctoNrcM5B8x7D+Oy9dimIRgwfOy4ncVT+nTixNZwG62wQmpS+p0R2kqzB4C+5
zZXTB4z5bUEfq4bCvsMRQTezAEeIhDCyZlyG0X4fqI8+TmefS3WMnhniXjqcKyz8
Fg/pGCHaeUXTKZIODzG4fpSTaFIHyNm1xRhGIuYamF2h4bgfqcdJY/O6fYqF6Evg
whNsMOdF36ISNnocEJ43YUVpmuS/7t958HgS5S0gkVdtQDQsv1FppQ2MrtmaP6Zs
nuf6YdIlM+2CnWOc7c1icHOPOOSPVwZitGrWX1pvLLTLgyRuWW8mvIThRMMytNrU
mavB9BAbav4RkDT9RMdSRukZOO6IOWWtYRRoHMm1kQW7Zt15825o3WbNhjz45o2W
Z7erN7+BgfBHYjWvkEVpGyR27+FsTzdW2I6KGskv8CfcsPktjG4LECYQBKnXrglR
Wc4IB8t118C1kBW3L95tp8rHdVTYkUZr8SD5jxBI86zspdl6kxZ8mGLLAsPHEgct
Wlh8FyZ6Mj/i/gyXybjFel0mBugnDVRpRSi5iAAWWSif7JaYiwqAenlCzzJ5xd9x
xjQAnlm493r2s5fBxykvt1hM5uJEf5N9aizlbLHf7qTlZewFy0LGGQJkFHa+eflv
DJ9jXS6HewJBxyqOOU8S7s8gNIYvVhPX+qw/8ue1XxNAqYkxXExtIHQHeHoIgx7U
UGsZxDxbCh4CJASzdb7LLFwTFGSYuyUe0p8bldH4zXBi1uyqY8hDI6Oqa03GyWmh
wdL7ubekq/BlLoasybmvY7IS0NolWpi9JTcgav1NNEhlFZa1ZZlDvs4oMywmYL1h
kT9e7VG9XuvAF5CVdpPOpeOBWmDO0EFP4m5qlKIXQoAbE4qltcYF0Vv8KhPfZOrn
4Ds6S5uOGefVCEv9iZ/eb1SeeQBRkYWve3MKT/+1OYSQrWtXt//TSc+kxMudUYJ+
T8mXrl12YSt7toVmTxuqRWQGs6OCRwqvdw+oQPi3Cidq2OJ5/MQS/NQJo/kwKA6n
4DXkDG1RRKVcbb2FIG4K7KI72magqzvssHrh2guNlHbEU3gYOguxkSrWpRbY2DJj
f2VE/C/1CNeDrEyFeQDHnIifw8oLuHr6AUUnePJrCKGK8Q/Ycz4ZSeQnWE4FvqYg
iUbOFr9oRKGoWTsyIwHjW26E/WBa1I2YrHoCV+5+xsbzczvZsuRNdPpkRsmzonxp
/xdVMvsx1iK/CDszH83hfzRBYWtky1PA2PFGo1PWEQ6iqcfJ6fMhcJBptxiN7lq+
b40tVt96Iz0JX7e0qq8n7TjSWYDZufaEq4IY494pnmbkCesWKIKvfohEOTOKgvYX
V6G5oFJR16UsRHiHhhzJFngwbG/dbCkHjLloI45GQ7tr1UlG8IXlkJsqkJlQ0b+c
0/Gz30GhvcHS+2OvS9pimqzfYx2QwXp0i+TYs3dY0U8pbxsdhSLSTnx5x8bukVoK
LInYksLqoCrZcFnfrZgh0dC7g3R6q1g4PujrQntqs8ZrHrPLigpS+6pZWRDLloO8
YPe969l4XKtR8RLjAjBA3FW36NiuGx1HszJubk6ofDcY7vCn6h8USHSk61YkTmwc
gx+byDxe3+dnZWNqB9RAi7Qt7FwQt5kwWCq66VahqCorfHs6J1L5eAmmPjBd+odK
Hil2i9SjpeD9eDzup59qa2801Mv6b0QT5t+tHJnzSibJI3TqSRlo5QEHZtpFy1iM
zc/Lk3JgnnmQ+1QkZtBiM71ZMomtz/OjP61Pgk3/r7CHBonRfrfN5WzavObb/kBG
5cIaS0J1uIe6T860naNMFnsNmJy/fENilhF651DB4T/CWx+ZvKTMWq3QEgSMOCLN
Mxd3PZNuu5AP7CO5+tZWKLzgl6UlHBPoKU4YiOSN1yiLW0ByDjh5HvMX9y0Tiq2a
T3k5JDdKf953eAG1Cchrbh4aqBE39mnzL7vPXqSxAfAC6BI8HZSTjcWYC18idmjL
K51QOguZdGBnUlHkqxwPIE0rB9iNgD91816/FVx4fa2+u9OLOYJub5sE0FkwiZLj
qXy9+LJ9LN2osSF2Aal2nM9y1VHLMJ26b4yUxp8peMrtlJ703zhavwBQpzH+JpIJ
0UFmpAiPhG7UFY8R4oPCQyg0vU8EVSW3YgsM3HDdsC20Yk9cK42BwHV3VDhnyrS1
1c+wusqS/13y0preng5BW3OlE9CDiTgNT07Wc2BliEZ4rOqgU+NeTO2C1LQwcvaa
Qhp32ERu+qr42j/NPGLTJhcrEFjK3jiWctLPrlufJ86MV4BgCW0bHcSa+PigMMBL
IEybmH5y0t+uHdPQyK5UXqEHOygJWtb3ybDkEzb+lqPhc1NCEQKpRe9E4xwJinHP
Acai6bovN7ZbbCbhp0UMwpbbd7naG0mgJlYnEudolFOZKA6SaHldkxhEcN5h66pk
S+xi/maOlsdPUP54zKYX4Nsms+rYuvim9MSSv0gdiXgXWmtyiXEj5qScnjcu7VPc
Y37jRSyxzdqOGGx2klTgAtBhijjakTRaNd5q5KPkBM6PreVx3Qk04KYlmYPQTyne
29st1OYVPvA2VuTxew//zB5DYTdP6fw8Zdx213700uu1ZJJk9I0ubwZjFQyLsY80
JXuXiy/dqyYQV1uAyCLqDoEZTzMqcsWWtIvvLm4PmUayFgM8703dlmMPGzW8orrs
r5MxJ+7/rre6r2AIKnyKNEJqpiDvnZUE9QZExhYi99BS7EFPL+ZUpQBbJrbcAKB3
18prRZIXhIfcrKMl54tCMq/GazHDva4GQtKipv7e5193sgQPeANDK4c2BgNTc2a1
BAp7wkU3u4cGa0REt3fq+onSlZhdH3owzjJ9yCD9r6p5s2i9OtDbca0+/fcgmY6E
nzrpaXl4aSaHIh0qil65VCwid4djXSiFiZf79XFW68HXaOhBZrMdT4w7ocP5BnRd
GstBAc6S1uXcdCvm5c3X9Doa1FVGDv/o2Fu+2pG1YwxYdfA4Nl1LbuG+86ErLxL8
l23giyKCHrOLG85gjZ9C5v/wRczp3UgGL6JNRgP77tS/nB7uETTL+yWZ9Jzd9GjS
+W+K06O5m4gnH5ws3NAvRVnLV2vLJalh1UCWbEKxK2B6oI0fXEPHlQzkACnpCQ2m
3FQ4pd4ENKJWUj1hsRqOMdm2mscPaC08by1/6Y3G/3NP0qW6f7/WzalSPfZ4Cn3i
mCAH/Uq6XKb+LGk3B8QmDprqxybQebLE+zWPcZe/r99rcF7bfCeog7+gITMuStf4
ViltcdX4e2xOJ81cXzAr6z/9+qcp8zJYyCe8lS9sK7bhV3zaRZZEjWDuTf6cIptI
tMx+u8S49q7Kd39JscHlIro8efiiM1eE07htev+7mihUaxfb++uoX2CV1KfmT4oT
dyENLiU79VszoY1MfZhVGR+BY3hGvI2zRyFYWTjgwqM6snhKG2z/kbVaF+VPEbdG
iGj5IYaUGvi/c61ImCh9/90rpXt1DXZe6dycCZo0GYf1pzTYviluFS+twEIuaLhN
9TYQI9SwzNV8/h7jtdsKZX2X7fVtSK0JVD+r5izukSm5I0+c6UgFlN8vcb0tzfqt
+EHOeY2GsvWghy1BDYTLeNWplv6xeo+fSwrXnMFPXUrHLHVhneHeJVHTVdm7bosm
sy9644/ElMRRzThNLkOp+Yn9ErY971DE6BHPgm9uc7E8BsPHEJ5oxwnr2oA3hJHS
3JZWurXJFvKYxvw4/dLgYZQ4xCQKaTs/iOGKYp1e3CecxAYLojzQasOKlCMcbKRI
4XQvl6hqZ0KdLAHOOXmRwkduKaQjqpec+iiEp8zu8tMbQamN92czxqpOnpA4iZNj
FjBF3HZkfesm02PF5msTnVTvUIIPCo7Y0PjVir0xugxEWBNucVL7TdlnwGnVE4Eq
LZ1kzo3/9FYZAT0ExEbVAfKnJCIwhNQAS3Wk5xkXaJcUyH0/EaaEbL66LOVRcnLa
7PIQDShUc22Qf946exeNEBSMg4OfwIQHwQd3x1q9hHW7kuQY0JEaFXs2tS/cLOAn
H57rX2nfSLeN+tEuSGouBxvfyxUEnYVZ4ukiL5OejBDLhfniVd98IpPWKfgVIBjY
wbkDA1VJc6+xaSfuv6ZE3IpVYaewiyEDjmcKF8cy79bH05glB/mr3fBl6m3svPDB
`protect END_PROTECTED
