`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHPK/xKmCbjl4yNNPH3YkJKeCuva2ZCsx0bFMmfK3huY
tPCfADTNjXqberJuxjnjiu8eNOGlIY2yhoNLl04GkUaMrd8z2juXaEQNOOUb83lf
gQJfMMY6wouH2m0tC54uuOKaJeUSLFfkJ/m1/w0gzurMaoy+MFDxyeJgjANuOTSz
8O0XMBRUCT3m8XDkEQbiForxItFoAy72sdhaSP5M5yKc5Wdz+kjKVc+8KTWHAd2m
CH2Ygy9Oey35Vww2bgAblmXkvh3v+M6WRBnxrSGutgQDhZq0/P5+de1a/A4qEI7D
0P17/eV7xcctDdqqu8r/qTkS1fpNtVcw4sGQIZAnVRblhDsVdvzhHYu4uqSKZvyi
8Lur072WpAaISP2pQccbCw==
`protect END_PROTECTED
