`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
VXCKgYp92iDLpF49RLUAY1c2nMz/PxpLSLVEJ9VTKyzLgAfnaS38olgav1lnu8h/
TELBHCVUs9iyi3rsBxKUWiXkSnWNxZEQc/UqP/YV9yK4djZw8f2CQ1kpGJeWvB5G
qdC40imea6uouFBeZBpQuRRvlrV9GRRyhhLw6EiT8KUL9FHyCyU8H7d5yxEweZ99
`protect END_PROTECTED
