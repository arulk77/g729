`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44rTESaaRgS3hphDtSWQVn2BLvF8WAg7N7NZbenNB8jD
uRzxQnNvdegq2MGXwCRrzMLDLbd9v/GXqKGtKANCXtF+l6YxIdASQ0w5O4HnyNSn
g0/fGwqprU+YWsIMPo7pDcyWjHZvGFl99vw5PGnbHRPgrI1w+tNOcDlIuKgfgZPI
91XWzsAVw8kEew0qPs+tV6mRKE8JdjDA14us/Yfsr4DWBmVi6TBNWykqGnm3V4OA
fTGH3Nn0h8uKsePZOa0WJsjt+U8gGcn0udm64IguUzMpmFOBvsazpckkiXwcWpJJ
n/MD10h+j6zCYqOTXorF+g==
`protect END_PROTECTED
