`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHl4M1bGaxSxRoDRYnbCbLbSnWB0xeo36+LeJzLuSLh9
2fMhi0ihbZ21C3Hckl+vlYmLOUXiQHH/U/PcAI3HkIpI/lr9CnBCjYxXFJxP15gh
pym58fNq2wxQZ7rdPNgITKL2qezbyJJ/iW6T0nAO45HnzOVOFSQ2gOg0GD22Qn/k
9mqg16YxxsNV12zFtHOEWlPZgldLHtUzEhCqConE8RmshAElHjXyWqULz0rgdsb6
m8oHvxTuCfwY0bbYdIt3JQ==
`protect END_PROTECTED
