`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDVavVda3RgzH0h8lNbU1OnZFkov+IPlcCWWNjhxfsqk
PULuXPEcK38O8tHC2zhT/boTC4N3/K1UQ00Nq4tYEqChRxpcW83CjP3Vl/GNbeE0
67+D01Ta1Wea685aSfNG1ppcLI3xlgzIAgFNNir0P5F3JqjWp1fQTT12uFriLwRV
THZnWYyJNspWQXEnSYDc213pNesrqd5aei4Jc9jOPoWn36ToOCk71GoOsZKlnD9W
xJrpFx01d5JFcVf/fHu8iD3+oCtuVHXGiDerDI+C3+F6aH4sfir1Aw4ehWBa9lSE
3oWjVqymnJJv1qOf/qdPrw==
`protect END_PROTECTED
