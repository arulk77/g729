`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+7rjLv42B8/ariCdeVOsJUyND1Hyd+XhNl24PoTnPPN
jZiMO8QoEaWg7Zb57iHq6kcqLOsoYrdM60d3wAKtf3LcNf0AFej3u9kzosPzfLo4
yAx1iRZoW6+ibshekw7oofRIsCqSQRS2jptmsWwsGHYvm4+4hN8pKJM1U3YqoXM2
VCq1kEkHdNoIrmLJmkLm/VW9YwzRBkJi1J3qjTVEQeW16RFUwFmvPSVlv5J4rL2T
0nh0i/IpWEDauZWkolt8YKP5Z06qvd7Uj0JvYf87B1XZqmijFZ53WSC+R0icqVZv
2FxsFzmP/+DIJ71IiUfRlF8DpvcmGGv2F/aSXF7FiQrlbNVkx8lV1ko4B0CR+ygY
VkJ4MEaIDKn0ntHPk15LFQ==
`protect END_PROTECTED
