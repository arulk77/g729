`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL227fsl1UujaRKzi+zZqTTXrELF2I3vYQBAr39dHnpm
0jtZqpK4M1hiLj1N1/dJWMUvie0fT3LAHMh8aFJlGkxPFQB2LYwDgbwVa6B3mjc3
ouQdnrae/5oFGyxawc5pmEaviPAuASxHTp25snng79Ov+I4ZzjxngRzjJVBiAR54
QQdxxpiEEji8/N8NdotdgvBlC/MBIWHoUW84CKk31OQtDw7ryJET1YO+9eHc6Bnn
SkHkNj3hWpsRAnBTiWK4bmEOzU/4LgWdw++99+mmwmE6AsAwnD4dUY0Pq26Mkb8A
VGk61/hHxW29aUujDk8dZ7oyEgAc4+XCJ3I3gxwDHgMWRnCzJmhFCOgc/7fUNkgh
vukLdGsnxw53Qo50KsN/dA==
`protect END_PROTECTED
