`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
OEqzVT8ldaECkSGtg2eL0wl3/MapKU/vklSRf/4luXETk+px5V4X2cJxc9F4yQLz
1rP3DV43mefQvkUQmChcb8/POu5e+j2/vDaN0u0ySYTcLBv5wURAB9i/Pe05JjqB
A9M18w7OiGDy6gVnhYt1iM6vwNU18JpXyRbSIv0C7YWY3ks5YbOQdgcD/jS98A+0
+J5mNxEQU0a7fmgSx0jCY8CR99oPUlAkpkuj3vcwYcmoblXd71MH8I4VpLGuJ9Os
DYazRZ1hlFWtupi1hNblkC1TppWZ2NaexKeONoyn+1kCFOCthtTjBE5h06XS18V3
6eJuJR6zAW0n4GuXF6W23BLwf5SNn/mVXdtqsu2GBw2avbBPyADBW8QjWVzH1Q3R
PJ5rE7qDAQrlFLrG2Hr9SL7sUSmweIRSVYMF/j5rypUagS/HhhXEVvR9UwGu35Wd
lCeTE5z7bhSD7AqyG6Tbkw==
`protect END_PROTECTED
