`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNzVoqiFyve/D8uxSWNmwGsT0T0L01YckAQWTRZTi3yIc
LxaN+R/KGDgNYwOkp7FdC2wtgfEDigVG21Z2+txrDCHfSO0BfnOFzRp6HzNMWwUl
2u1oEh2euDPvNTv6o3V59baPpzImjs868+NarKx4quC0wIO8dFTY0z6Oyg3q9FlR
9u3wTb5fNCuIj40QfcriQPbdBKUCvFhIuhZbVYC+KwgNGKfSL2K4j3lnhnHj5TEP
Ie0z7j2csew6JR9V0YENU6/qm3tATuqXQX0vuycWeMG55X51VdV30RznwksfHHLE
BRNQPwY34ovsdFyEyvxQMuJC/Om0Fy97I9KbwjVh66xaxZ3CpVzRxf3Wng1Fd3eJ
hsrIuL+qmBeN30e4x7gNAZFWt2D5o7x5rTzoiNcvk4qxNZXgvL/zTsfU4ILrL2nA
/Isj34kyM7FRjJr/4JK0LE5FlpbDv0hpaWc9t/54gpokxAPcQajxTOa9254fUiDi
4HCn8sv+i02iIHa1Exlkfx0DfcKUAZK4nO7ZSQpkE9Nu+Y4BHT+CFq3oPfUurC4d
Q9ylXcS5OllMirdvFZgyf/MM4twU4dUPQ8wl4kqOoWWhUC0vJe8cpZXe0/mLTQWX
mC34r/R5XSjCFNS1z1ysSuqRbdWjLYid+alKlbtJlp7XB1ha6XTrBiHp6PKaKVXk
gC3i9hy/oUr2Rs25qsxq8NjmkvuB0XpRGbvADcR1uFAWw1w3ik/XgKiOijVqlDyR
rpMLrT1neo2AWrH9+8fxmh4ij5C33BCl6G87kg6pxGhRLMWaNszhhmOhoDfHfcUI
3yhBeTaDnvFEQOzWelPVnMXh58mdwZ07/c5f+mcL3hWHi0EdBs81PoFXZQNfanrM
HuBMC5JN6/GeO0BLy+lWYcXun4xEj9XBYsLIZ4AR2en8PiCcTx1ZtqKFCdQhWtUx
p81NfRHGojxDXhz/2jEj3Q0T7yl1FYNS6rekanROYxPeKMyPjfQ8QpcDH2kyQwMZ
qfnSu2KoiBAi0tGeOAv5LNZQdHMOxcaUWRCtPsP7ycCUhHyFk9oCmJxGaJr02yvc
mNwHJK6ImMrn2ziSsXVHacs6rXv9OU5jz8PD3HTwja66o7Xp+sCbFgASsEfoaJJD
UDK2hTdYcvyQrEB5hrcifYDhXPrfIv8Z9OTebWMpLyp81CGXBneda7CX0A0j8K7/
ll1oG4gT307By/DGVgLshSJCF54QsvINvuC3XDpVC8egUpka09brBQIRF33YfhEc
t94VAyAd6tM2ZRokfbFAHUhmuqOtU97AoDwUd1JeC0YClqce71btXrpucrrCdU+j
GTFf3C+WEq4yfM40qaz0wm07To1OlD3lW5kNoh0zufbRtd0MlVlCA7nn2eee9QBd
jEica4b+ScCfFIoW850aP8lhF+VlR/igHSxR+e97OK0=
`protect END_PROTECTED
