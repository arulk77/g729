`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
BdCB4HpRyWC7sw/8ggd93Z6JwcBRs3ZdxCCtuvQygl8bscTXvCTi7e6r5YAgOn5p
tcBOxIzNmQV1EAENCXrGt5gxBHi0DMFVTFGL17c2OUhkNzkzYqZwDiYMY0VAHQf3
SUsW+GY6/XEUVXMZjqb1L7nNj+7lLqslPYRqAcBiZdvRYKaykaMjwg3TpEnDwV9L
T+VJqx8diUIIkRu7XgDRWge881BK5quV42tRwqnBJf+8+lDAZvXz2lEUVblY604L
t4HswVrGDX+BAzdPRxKsTDUnvgFedKvdpSXUOBLFJmu33siskq3hamCDHN0sxEGF
BsY0/ZTuq+dm+Ti5YajfZ4JvEo1dQIXlo4QNgeQaatU=
`protect END_PROTECTED
