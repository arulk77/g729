`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDNupqlus/az7ocQDwtxqxSaVQ60scqWfICNxumoq6e1
orLZ466uHi3HAgOmpSjcTR03/H6ynmfRMkvZon92+iPll9I3Jl1Ls5MblNlDNNP7
vvup+cS13norqKbqsBKoV9ScrUOomLOqr7zKq71itRORxGA9TW6sAwie96X0oF2B
QX1PLtRp6ajsD9OXjZPymmrfaEJCW+c++jj0uIqWbCxbvjdBUWap8+DHrGmWiq8A
0DPQBQ7/7rctrsSvmybXON6STFsZAgrs9qangcWM18+EJ9uW9kHaCqjJdRJyJVa8
/8iRkbEOgQF0tQpRzv2Bag6d/+Bk0fWiYeZt9OuFWXPUqUum2ReF8wlYKI16HI1b
Gfojoh8bukH0i0PT8C2g2QEt0kAsyrj1roldh44ELF43v0VTWLA5eKRjt8xATv88
gC+FEXxNMJQx6W2N7gG/eFIBqPZ1ZC6yfQJdXkNgp4qMEE+blxGZaHPFdpM2EurZ
/jowIhcxrdhgFhvlAim8f/sJZJn3UNTtabhKA5o0QH8cQCDPqS/UTdylFZ3W8kyr
`protect END_PROTECTED
