`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
E2oODTTWUOLakJnDyc1oevOH+DzMuoSByrpDYNUEMZ2taeemSeEpKcF2QbDQ/MMI
BbJcI5Oc/rpa93z6YpSzn/wQChCx4kiLQUNw5JsHWVAsusmP7Pnjpw2JW/84Jl7O
bO2oWzugr34sRZ+LwpXeH2D8EVVqyVkhm8KLsx4khTtmoI1+/ThkefIe1apB0Q1R
`protect END_PROTECTED
