`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4ykFOabYSqzJ6mgRZGBodW1dWJDucGIACv/RfxWCbRKC
1zjwNqkd4ia1ZP2uiOcQgIKCpmzADlDnc6HxJSWGl7BDRPMItyddLhm414ogWtGk
v8hP2M9WDwGPfWL/GprjaxOLT+UoqSZ/EfgGSdknEqSmpyopkSuX7DmPKvQnun5C
rU0Egqh/pmBXPAHDZKLgN2FoCBoWY0KCg0rFonvEp2Iomhktcy+0LqGIYC9DOD22
XwAigbd/xLHglXVs7iuPiAMhGD73+TsehBEPFLO8tOk=
`protect END_PROTECTED
