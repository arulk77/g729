`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ab3t38y2wf5+qsH/48ktMHjcP8fbKC6djy9TU7SNQlyt3OuAtYqRJJoUWDbuo/OV
qdcHRi/79/SYC76wow9HJ3W42CjaR7Tb0LV77Xsjm78aEd2mY0KFgyZYo23tGtvb
XoaiVXfI47Li7DO/7vtoqA+nyKPnZrcnncTlZqr7uUVyVleJ3desB5tQ3ipVda55
ixKmaMUr4j/Y6HopE+1Wbli8Lcm3b+A5qS3AG90lWHOPuvFUj9jDghdYgYdqTnOK
gk2afb0PYobanf8gGmQ5W1IIBU52VoNHL03QKiR068/z1I2TzxmLb65EZTPqZ5Sw
yxeJDnwKtQjHYIlCwyrxaxK0XLW8NdGJ9GuqjSyluLwd8wssqOKI1bJnz2Lx+sBn
0IbXNrtMnhWJZyncP/nnaGWNIGZFDLNKai6kezVKSAg=
`protect END_PROTECTED
