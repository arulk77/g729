`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C6zaxBH08SKPWiVYPX3nzSWa1rIpX0O/z+/X9uzV1C0m
1CI98qp/lDX5RzYnbR6mb7KzsmeYO8PpLhuo7WQsG9X2TmoCXCPyffZyZq06+yqI
Y0tOzlxQJsacylwtlBySU+v87at4DfMZpsU3S19Ghp37I3aNjtl2vE4veHBkKf7e
vW6LTq95gykc5yQ+VMywdyTGvvAzBJqnFkZZNkJcBlmyRnmAXtlm3DdgJ6E21IkJ
3XwlJv3soSVB1kOFq3fp2e82u6eR1wdRqMwQREcnGDkhFo2g148L0AClf8SMwTbF
R3mLT9qFEKJZzBopCx2W+pfchCs5ORlZKS4j0vdi/A9AbR8jQlA7ht8l29PYpkBj
jripyad74MTPgzhwm4xKAD+Q257au3hgPaBhC97zm4Pa8XKDk1ufgv/cHw7/Zon/
WPO2dfWJfKTnZTqtrBl0KrDa2vNtM6mTuOZxmDNuJBbDXhFmBpafZVosLs5A3LCc
/CCvoQcxg+o8UdHOwNJ/LwbTIt+MIkj6RlA9SKXXo9PjIxnXURj1PxraxFpgOl4n
GI1xdBIf46Vn6/PL6N9utwC9vUZrsYuMNMfqeo2dYDC9LIfAbKWQB+FwxSzA+m9b
HcUeeCrH3Rnlta8n+x2Hf/6p5Rbrv5lR/br6wyY4TEMAByqoMmphVoBgWhpXXGRF
9dybnLYNdtP3gryjMZ7WkHF5Dw8V6ydQhyfuzWeTbGxPybKvSRc6Y5Lo5vlvcKyK
wBLGq0+naVsIZmFOKdD4zxRHxIZG4XSYL+u8Me7KczU0nlU+6CjLQMAJ1ygV+pXh
Xl+kYwDGK4Yg4+QuYsjSVHzVEBMfah5Kl9DdPCXDEAv379sRDm1ebdpc0WsIC+ju
3nxPlG6J+Oia8Q59afhO500Lrz/x7ZVjlbJFcjt62nYf2P4tfMahpLUGboTNCUPj
uNjuBrBpmB0Pwv16clvY+AlMp6MzSBkSiBD8t+2Yby1wIixyvrdA1pnD2XP6zF7s
v1+2+E9mj1+/pC5VS2niTeEWnJC6LbmAwu857s9DhHgn+GNsT0GMcsT/1FKrwC/H
cA/eY2yXSc/AUnkp4B9PR5P2I9uq8LIPYoQnNDi8ryTyhRtylDXfBIajDdtrgQXb
AUhXiyPbrE0eutcv1mMefPBBV6PKv1ORQjSSdHXpWTn3tsnZnEJ62eDyXviECjQe
HhRdEh7BmANmRmUOhYD8PYU43zLKOaK+BuZ/nVn/5mgRAlcz/Uje+aKiT5PSJXxg
1RJl7dtWsw/Yp9h9iIs3KWKvqVw2MM2AF96eFxsh8XUELDoTcQ0wtNcrJX0LDj5Z
ukmozW+eaLwfWh2jWvygQS8VEgVuhbE/vx2HPG53+Eta7oPhX5Rbi5UiF26q8Eg/
W6JGaI3dz4wgg/IPbwZkEOx7+GuZfdfyj+l/U+9Vd/Z5H4M4FePWp0s7vGwt/CMa
mdjdialh1to5jS5FiASfWDLeD/km4NYMazqXxbnGHRGKWt0t1x6xB5xEbd29VdYm
TkqdVHfWBmKEYSOrkxoTeYfSeccNidLSZblMDUWIQ3F2n3t6QVpOd5jl7zcovjZo
PYBEVOoF3qiTfhN/cO3s2LcR6ktL/duBgsz7jqJxVNkIE5ubtVgWxA2y5k+k4McI
sSWgOQMWzDRHZsHMUBidfSxSwIuj2wuJK28/kESwwkTfw84D7mckg9+rKFvAVn5e
9hhrrc3wWHYlHvRNT30lxJ4gcMy6YPmJfQKQsWcADIquBcW+RqHDrx18k85DE93s
woeOfok/D6K3v9pByiPw3pDE0DSG/U8/D38YbQ3p8N4S/A2uH5dAOOCnd+GmDn2t
MxTwzuVvekQAWAkjGwjjdzIrYHRFFKQzHLn+5YBfmrgfPzlUtv31zzzNHK6tdn3v
QLlpd/mw502MrgI4jybg/3lVN+pCJFUsLtdHf0WUwIyZnJtBrEW3f/kCBJuCPVH7
`protect END_PROTECTED
