`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
AF88HjkcbhBSwVooprXY1o6zI0GxKsp/V8ODjtvTetzWWPM8is395lA27ClRN+5J
v84U2E6xe9j7AtUWpLznOPMzD08w45zjyHSCrELu10Z6k7b/FctKbJcIPPabB7hy
M3LY7/UpiQgRxFOizRd6t3l1IDKIejxJVeRRS6/2QBVGMNm83p9djUsOw/8AzotN
WJBb/WSazEWmmlJ4XXaEPkmtkfVl4J9JFcTvyW6tzG9c7ZStVB743ohKjz7kO9tE
5AXOeX+BsIa+ci2J3KaAtSWJ5r0gEPU0CzXpX9IwSK9uiTHZEmpHc8oYZ6k+Q0SJ
+ocpep28jl/EiIMQzazmzK5RDITagXxpmSRxcEFaBzBhZawkmtO8kJlz6Ev3k8qK
R4CoKCgRR2d97KfVdg4fryfKrU/pmaZW5B34n5wpYGD1m7Eji8FOCRToVZXFDrvc
ISUG8Qkn4MyWt7mv8qcpLAcAnSrDuhFvkE7RnuizdoVpO8UWh6ZdhIPxg5PP7njc
wF/40NEV6uZCocTAXl1QJFilqmuoQeW3Iwydoi0GaaDmRr4V5DmxQp8+0fGAWVXx
TxylmTeX9wGMkbJ+Zoj9L5vSL9rzqTMopEvdksko/vDkTkZNKGMRR5E5alpjHaZ1
J3hVfaO0fspZtgcquijwJA==
`protect END_PROTECTED
