`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
F9yKDVOld6yrmzcnh1mfIovORnrkj7tiDdCJbMrVO1arGiwBf89T36qtOUIKUJYx
hy/cmtKiAoy3HyLJ7hoelxVAp+pzgD5J4nA+NFjaFnUJ6jR+QKPDTTt8x2Vjxs/9
AJTN/kD5WhSetMz0c6fNM3GD43ektuYNZEH02AxBp4zACn6KgJeFDReGyFs0J7cm
gPjsxVqdQhxSyWvgL7XRAOB6XTYNSCvoNYxoRdfFIJI9/IHgBIKBCub5sHS51ePi
h0+nxjy8fYj/GUWpGIxNy3V2rG+4TKlnm9AqrnQFzsRcpc6HYpFZmcZdo3pavO3d
mABaQYmnpPb/2UjaVWGGPDctR0793stjkoyYoffykPOl9hzPLqUBb2gdC5ONxqEL
CrrTIiY++O9BOpWy00Wwdd377kqzhfpUV2/MRWOhaUMc54vvG3I3tyh3YQETB+sx
Gqvn+l0koh6mooclhsVelTrCdrjCKLgoehNfsysbZWL/wTX/gHaJYBsKQJRUFabI
40EU4g7K5FPTbIhh4kBfWAm5tvo5LdXYK6WrtSayGpeS8Nd8JyByvGoQrnGF1e7J
gG3Ykt7IJxjjNjca/rF7y1Y5h11tZeo1RE148ygdOfFgqXIU8svH2MtL5aUipNt5
UZZVlMF0fwV46cPnsg5KxDYhrN1oY6RTuSwMqI8UVLb0hLgTwYKhYw3krqL4U5wb
BYh2gW/xd1R5dcAT0wFQ01z1CsM8AEQOtoP0FXZJT1mP3Bg7Q62pSswg8WBi9DWU
`protect END_PROTECTED
