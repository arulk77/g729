`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAQKI9oiHkz60Pigt6DkKqTWW/Ej88a+MvVTqHY59YQWz
X6HzgzXfXOfcLUdiowcwSjyvijt9YhNeIG3CFfGymKDy7AkLleImcNLXJQSPQp4M
T8EzBYCBxhag8KWN0AX/Rlx+z4t2EadXRU//KCRcnPxU2vzJU+JTnoHuyHWOIZ9c
CEcoC+FjdW0H5bsbp3DviuLDExVwUJ73DEkVH0QWPhkXA1SpCSKChFpNWbRpZEvk
Mb7rW24pJcyIoOXZ3hh/hOkFxxfIha08+TkLv7lJOth+3/IVoYtIlgCDobG8qmt/
i/G5+NYmB9pxIRAa/TlSUY+AF5F0rA2lvsgh8Bbe3ysngox/TSrvYk4+hbqYzHq7
lQmpQfyL94ERC433H8DCKSKeRzp41ajsWltZiWTkHJcCh06MeVzewvW1xYPKsVx5
JXaCXof1IfLMQ9baCX+PrageZ3smvLi5wvCD7w7Tr+gkat5fFaMd4ElicwN4SkK1
Yco47ohkWNNNNiFXZWYlUtBdh2pul6wtJ6jf9C+58pT2i4YPtk9OTM20hLgVYiwz
IGq+lJVsh4fRq0Dq3wuukPmgzkv9qNm3qwvY91259AuaBQwL+u+j1rueZyfkq0iY
TD4+F1vlFr0MlMBz778dr5C2MGGQHGalZOX5Dk5JPgI1TSHTulgIMk9g3izuBxpF
2TFMulFH2YE+xFe0HMgqS8sXw/0XJEdfQtVcKhzBelsi7ojlANVB5tUxiw8sz9o5
ToBAZUugKgQheBkPY4DV2wEnbughlc0CsG0vb19W+BZz3QwY6g7mN3G+QJ5KSjwf
eG4MB9pdywgtD+Usq/hdzaoLAxwGBnp8feA1DmgDhHjwV6QMiWYIR7uP+6iS3yn5
oYoSD68tNR/9BTp7+6keix7iP4ClXL1Ef1bshxqOXxU6Ln/UPz3IMGz1CP4Ndl17
NHJk7smWj3krZgFBhFnWl/8VnRsCNNcB2izDxt7I2KjpBivUblqPqLwKWlm3N/4Q
Ea1sLmXNBpVpj1fwOv4IuNnwFnby464dvhnTo83fEGo36QrJ19/jamj/tBF8aImK
llHchkmEXWIANa9tHQUuqT2YzysDPbkO79cJle9Bw2yzeWHW49cP8JVskfoqS8tc
a+FbKJs+F+ODEQWGpD7L1WcEZOCiDd/8FDG51tPH6/FzqFPWB0dXhmddbay6B72k
Ym3LckJ36iZk7LQunOaq2Le/IcBFCLMeyfIlpsK+wnwXzjkKIQZ8AbylGnwAjIfH
HSiP1eZ8z6Vl7oH+wLKOvdgkQRx/DkdkbIlDLyoTJJHkK1cy+dzSQrEym5+Usc2h
i2nyZavfzZ26TKHz7hx5cGNHkvhvyd5vw0XcVKRAB9ab6GDwDTB//Urdgw2Vv73f
sRBus3HRWhPdmvZvGAoTTSkTSTksnr8KFRZGlq9Cl+bYEk92Xuh2cQ3HrT1lOqlg
QWQSaXKvAXTKKr49z74QTStx5Jx+B95ccN+T3hPKbDLAmL4SZlWh9ltSKUXIAwz0
GHB4HhmDmaWQg/Ds404t40wgwvxNyvVFn9y6useiqbnFwqPdb7qKmcIsVHZqNzs5
2yY2NcjE5KF2f1vZilyp5jfl/n+LvhC+Nd1IlNFw37rsdtvi5b5MWgwZt+BhMmhb
5SCl01NTjZe836edzSw2Xl7U/eYdEyJcB3U4Oy8iLn6StehXMrFHyuclCDnT5+Fy
vh23Lzht6n1UMmlSkuQpdSJuK7SMWQDSDbm8qdie7zTTfl9PpeKqIv5R68eihijp
TtfwpkgRDFM8poI9svg9hmrGNt630ZkCTBbzNhKDwpyfhphzqzr9c6DwXGkJjAjd
2a8FBy6YefCe4ZPm4tao1H08WbSK1ASESRPCFlTUEI2HrP7CVXnwJDGcrEbgsB/F
tpxv3uN6B8qeCXhvQ8Z2UuUnuvMfjAy4sl+CZvnPKsG3Jn73q+umMfK3h/O+1gWe
jk8PXBwHNnzOYU5DqewSqbmJad2LIoKK+kNrZF2qeNv9q93TBi4TDz1AwxzuMTLu
tunMn86fUcFmdeULTNg/pB31/cUISiecj7hqHztO03pwcjyqAswOsnkaBPsq8OjK
kNwwflqHHeOYNa3iAZzauKczvdT+N5TzLqQELc76UVS/3iAvbKO4g3pbUxQ2iSJy
tljMd/RmA7UjH6flWnNTGYS6Kbo27Ek0bXfxDjZEuxJUz+RDCc5sdFGQ8zMQLUKY
IKkBXpOiv0+UK779bXg2zQfjMNvEPj4MzPhtlfBgMOgnS3cDs8h4VPOfWkHLvKEv
LCzDs0K7ofsCDh5LCa61kpSXNA2SXUbAVRcnzSe7zm2QVnr2gdYjf6XWFq4/bPkG
B6QzJVC+IDOLMD+/3GQ64m7GxzKYvSx1aAnTc89CHJmgBe4mBRcu1ec9M4AgmtFq
jpLw1Kb3ENtsDeO8mq5SsGP7IEexDr1ce5mmHIIlouSCP7hgh8EVebhcvA4V91kb
4itFIM/E9Smjakw2js8BgVno9IvfY6vG1phb+7Xy3V7CnM/vD6WhOsJ0IXAJqgkT
DFdKc/RUefZvZiUH9KOOCi1YP4LHjwnruu4Fd95rFkpkXxufy6a5mXB4H51H2JEv
2YEdLkx/ZPk5alFg9+CVz1oirreK8WMgnTwA0Z9uDkt0nQbEvOo6oOp5wTQDvzUW
AsvJa7zt6T5z2X831azFMHnccH4gpFxk2sSwxglAbkxh67Tryw+zShudDbd+isPK
SDpRIMYfN7Ayjc5pRunk4UK4QsvZm9L/EFkfbJAXS+O88ZW4XFvLt6wk6eTNJw4V
UXO5mFUSVicJuWJ5TJE2pOExt8jtiG99AfMqckqTIjfm15exQVlF9jy+sOpVgjl2
Z5xhzOKbjUgwaAfTVFUHcz0imUvZwumzB2+1BKCJQVolOGjPuGxmLI4sSFhlqfXR
lMLcpXOkrgKN3ZL3l/McAyz69mz+YBRTvF+naalRsoEzTAIK5vl/MnnAsHiOsr7+
mJ/XzyXAwy3Tm714JWUNFRCg1156oA3MJqX17jLIEUXx8McqRYT0LMzpeCO8/79b
7r+CC+Fljb2CBCUu4RBn6CNH/Tbf7jjp493uPV7TLx+sjDFrL0mTtHicrjWHgL/D
`protect END_PROTECTED
