`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48ApBOLbc8e7vtsfr7+kzQ/j4g+5KwKhDs5RwAYca76c
Lp+w8YltxLMonBy/80J1PiySCx9uRj5Y9sNcJ8R49OEvosZI0gLd/Kl8cuvqxMQt
3GXeAePnbJ1F7zFlqsdfWBns+Et60ReXCHJPS4fkxAh7i0Vou7q+QV3+whgj/qHT
eU4ojbmP6zuqtXEo8ypiOG8Jt+q/diLhPq6p5EnKyPeNN4ZhaJzFuoTNUzgmPY/Z
pCvWSYjmi18EI7jZNCurw61ozeg1DoWgVXaIoeLbRARWoQPsmYN6JoKXJ57lnUO7
EiZWHIi+0v1gSxmKO29uIonop4/vSRe6RrhCgUgQLpXLGY9L7CAInvjYbPcR7vHS
Ofli+tPHkRHtPNsw3Ukkkw==
`protect END_PROTECTED
