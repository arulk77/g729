`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
FQ+UkS0/fMgU1LARBoETmJF7Ry8U7jK0NeSdWeIKkQSGiv3BMWErMVnyJafB3J9g
PWBAvBCYwASeVANYWlvS0ehcAQzrPr4gRpWHHxY3Sev+z2D5jV+52iBq6n7kgnEJ
jr0xmQ/jh/35D0yNXoEjjGtqA83yYjekwUQy/BpqCdwc61q7/8ezLj47ESeArvIs
6/jyzS4Aq+nQEp6Kebq0rsgEHN5SlEcehwt3JkK81YJJl8Z+Jvel9zb/99cTdCSH
i0MGNRmkDdhjhcweLo9tXiaDWKIJkbNMqPe29J+xQ/2d7MFRAby5v/xA4DbPHJK9
3JjS1OOJ/dYP98ijE5iSBMmSnH4lJ7qsHrzpJRlWGS5wJDabuJRC4NeaUAn6ht00
DBJiTXRWvBw8+mlkExhrcbJ0sIl7hoWuROYlMjo2+7URTe6jusZbfprDBKJwaunX
CGujD75GmyLo5AQL4qjnW8nkEUx52QzjfdYT2cZ4QLtrXeWrEd2G5FvrWvR9YhXV
vt78ejSJQFk7d0Gpa5sQ/O5K7N4RSa0IMyu2VbBhYEOpdWwEtZldjhHnTS94Tkdt
vTrtqW97xAQpMrtgehv9Cxyfcqt+F4R6nfg1aJVx2msLNanKIZgEG0iDJOqiLi/U
dIP3kUn+P7mG37HfExmDhe/Nn5AKvC56TrB/STfSgw31lAqvyxdenRiVdYLh6mMG
lNI5BgcS9sukIrjqZy8ns/BaTk2Cm96u9a35UjmOV2kZi7Ms5085Wz8OKQ2GsY3z
1El4NTffwRysvNbQn8x8s91LPnbhKtgrRf+cdtPbM8c=
`protect END_PROTECTED
