`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN7lA504NidXuF2V2fjbkq2ElG2+4PU0zD1gRKgrZgWG/
07fv77nBMTWvivWLBMVQeykxKqtH95mCz5kR+da1cyH9o9KCQW6XR+jCJYhDoPz3
gE/kXAoA565F33B2Xk/3RQtBSYoKPgIYYurn0LwVmgzwR7pUZ6qREteYbToUWmPs
HeHpVqXtC4zsNuVK5rKfDue1a9MTdWBraAUrhteA3WsGYAMbZYv17tiTK18oESIy
MYlyYzBh8wIHtbZVRbLGaZCHiQbnQO6GIl8O4pKwsI1ClzHNGWP+yutovEsZHQxw
7/4M1aCoXW3jYSzM1mG15BHLbVFyLXU3NzB2LilVqzKTr2EihyGxkYQDs37inG1n
RP/kC+1g1s+YFR1f6OsSiXyZNSAc+/wvOclEwjcauodYdq1E5VcllrI/xjLCB7+x
Zm4nkcBMHa9OWM3iikQ8HxFtE5ijP/WftQlFiWr9ttwNVEwsmMCwEeZaVQDxX0hY
ka/Mfmwk8h8R3x4abxx1BmqOqFfR/L5VESEkquKGOJx4RTtz5QgnkuZDm74XDlqY
pQlP8xCmn8/mHg8tWsgSWt9lSpDSHwI/kbQLU+fz/xsL27aasrCWdDqydpr1FNLg
vtTiuFDgCO7tv6S3CLsjC2GdeKDxsrAb9wAgA2yHwpmNM2VJJW0n5Ezwg5BNde07
ccxeWQkw+hPUYUKL3uPLfr3ViU9xuO9x+fdGNdQW0KIKabZe0xnfx9tBkwaev7Wi
`protect END_PROTECTED
