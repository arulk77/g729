`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44uu/VoBMbiJxCibZa7nQXUjtAKjKkEqmLpr/xwDEBPj
c+rzWAnR1/nF90+RddtfofYzo2FJHtyn+nb5WuOnXncROpACaDsZzi5JNDYvr/js
3QdSLFTXGMT5B5Rts4uzNLYntkci/qfUPrDd+Hmxx2aXSy+kwkOGDdwM7FLroHPr
cQmOapktlAIjPxq0ExoiQmPPUHBozm+7LVXRg66xL+i0IeW2ZWzAEaEkR7lnJumK
cOKYT66JuMbeWEM0vZ+j+M6vjmyDttvBcrM+nGaG0CwSEd9vlhLr+Ism5RKmkPq/
g9VtsMBYW/uZrlVJYXQipw==
`protect END_PROTECTED
