`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveETt+lrlXFFPu7W4xt/VbBBPlh09Ie79c8y7wesOArtZ
I2iAAIhGf+skx7ik+V8N1DE2lIuD6JZu3mn0G9PmIxyRIcuU+JlyPPewujZBgAYr
sASbYmCLImStIoC8E/ZChMRGUkamHzGQBsIJ2Q/cPiYh1cdi6a5PTZVYSplwn5Ua
dMpnFOjGCFr6YMGVPfX1nKu700fiHXfANtRHETFxd/e5umgb2PnxuVa6S9lKGWKO
Rwc8OcC8qk43+vsBvZeZ3YgwOPVsMNq2R1BmOK8Xbdf2d0rMu66okKTfFdsmzgHQ
LfDZu0CNcmPKMdS4LN/B1PpDPCq2lgU6H1VBDuEUDnlbkqW+frUj+XVBphXP14ET
GeT/dt46IFTtKDhaWTiPiA==
`protect END_PROTECTED
