`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCoePBNQ0pmvaJaqrrmU5+BVuUVvFZ5YrE0FaMz6+rqJ
OTw0lb9QQDyVb1NlDd9LYcsToJy+/qCUIFue5ROZUlwtUw8ROfjc/+xRrcWlLkjD
CTsJlw0a1ozV87V7rjFoK/Z+eTHOfLSXu1wu7aRzGyvluLbg5yg+HwUy7coLXzst
dPq0vIVwBcbZdodUrNDPMS2fq7laxhJv96jbB9oAgBHo2n/wq18kBT8HixjoM590
jX49e3ZD3gAu0yrNFwtbc0oBlieJ3mFyuFht0VhfneDbgBTyweythefKf0K85gLB
nXiALTCEhg6b634E5SDAItgotEgfSkvVCu5lUhV09bMxp/Q0wAThPrmNDW9bMY5k
rMfW6SMTszQ1t1zqeLQYn4t061weNxcPKA2eLT07aIX2XWZMyuyUqOoploGS5nEI
bU63yqjEeiwCWFVcK9/r6FLgW0kHlWz3HIs+wBFlqoSfw7ZrQwMol9YTgJC6/3Cs
yVdjmik8ImV3fEIOTpcWYPj0x6RMSh/4qP118phDgvGxgwJ3F/XeSB9XbZdznh5s
`protect END_PROTECTED
