`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveC5awrgbX19LzIAF8/oNIWbBUvYdhwWRUeKtYeyPKd+h
cQ/rLdg6D44rcuRWgK0lnwo/xtb/DXzy2EQaAuDf7Ny9vvQ8LrCRcV0DKmSr8RaZ
krgdmsOV40W3FwHYRxlb8w+tOzlzjbae/YHMA6LhK5rAGKrv53UjurxG47P4uiQS
y1sy6niRL9qAog90Cj1WqA==
`protect END_PROTECTED
