`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFjYE2vw5NcKVJG7m5xzo5OdkUYnU32kigi0VOELaAXJ
/a9dXS+PlNs7zdeRNGQlpTaZaiJSC6zNRQxyJ3vmorEYfyn+fSF+Wp4q3BupnRuL
BuuGDFN1fYM3VAMsWjp/oyB+2aekG3+4t7FOux1nzD6VQA8J/StdBNALMOl9sszN
8hpI/eK8KPcaAaGonY7fDkD5DSW+glApQ4KyyuGc6+Wk1MmXbj+eJQBN+OIfDYjX
ijVP2WHNvBX6jbofVaxvreIGDxRaowP3W5/HKQu6UCWNJrWRHZC6ckRiRTjwunOg
mP7m19kGjEs5A+3YT9KEZsrgQ9TwQgBpTWCZLsY4lTvP8+4Tfuxx/gBuQ/F8g7or
`protect END_PROTECTED
