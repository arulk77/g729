`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
W52by5FksJUdhgHLv4Ym9CG7rFPHSXJnmPDb8jLvMxfxHNfyQUXBbGQIwxcyec+U
pZBfabxDtihkk3Wdqz2JiahRqSERerw1/yhfiwOxa1ouy31oSepFxgxjUp1O5/rz
nhAYgEUxv+hX2S5MY95T6JYPN3MQqf3fgn5TIXJW5cYC+YnrgDP6HFvgrspATy00
KvnjmQyEyqIDbuwzlq4gnTm8k9W/a35SAz09NAj5li6/9iRiLzqoi2p83tMRg7BF
HP5SzuuXdRbMYgMSZIDV2C306Ag0GNwnTZcZyvq+cMKVgrSWuWOWucQlE/PYeKsW
t1DgZMhXcEmi02fqH9ADz/ApgfEjN9TAlQQwsSgtNYA1AbJ6Q0R9h1z5QYJVk6iy
8TbaneieMEU1AZVBEB9+A9hMUsRbPYqS45iK7CQqLpU=
`protect END_PROTECTED
