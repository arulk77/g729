`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
HhTR2A7mHdPZJiUoV6q9dznZw1KmVGsfz6vj7t+l52NJOJGXofzqRrpudvOaKxvp
8zeNTXmnJmWxLKwsgD2QptdPrq2YI7gn300uiVQdt2HhGpRxd5k1gMi9UjNgupDg
dIY9OyeXG8pJp+6ZcBvxG0TgZ+eZp+Is6oykyzkZ6qAi2vrCPFfNSyxzot2Kw2eX
S5+5A9V5crQsk3MWk2aRFShH0qimCXDk1mjdQFix/njwUntLrJDm9qNtPng3PFXp
KB9aKQdF4JRUOpeYpkz2VFkvE0HXz0I7xp9QI6amHzhRgr+B/rSyZ1BFXtb9TDhA
KowFoUJR+t2VomUcxLptJAiPb1k/GGvOcb5Y9OvUyef/JcF6fb1rpRM6ndQjjiMB
N3pc/SicInd6ggQOSWbO6LrRS6avyBHoXep2i5zZ/e4=
`protect END_PROTECTED
