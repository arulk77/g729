`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C+n7dhvHoGlyPfLJNbTvhxkVGJPR4zKoosuIFnnMoIsC
jeFGLtRR3XkQBBw8xUs94PSHnzhcsIp/RfVs6TA80JiZ0BhF9a48BEP/T1pgujSj
B7Q3Y4+3b61t5pTmHnlLgBeev6+OMW8i29i+FzU8FuSUh0ClZYcIQBS7E6hjpUhl
PGXTix+/rNxmt91+/VqwRGoCf3uzpgOS0mzHxineskbQCTiOUWP1hQURbCvpNBMQ
cvwigB5AJuamfsWc6whZRULkNj+Rj4fTBEdZx/rBugdsB+sNlNL844LP2SdwPP6t
fvpE6Yy0qJ25F3ccV5oleyjMvyChC2kGajtMU7/JcHn2tx08cgbutYgnSZfx/ccB
ldrysajdhjBP8gbhbmObqlkhFRg58ObcHNm4ZvQoQ041cN8kSzPnl9HGkr7P1bUu
P0cKfzN1P0O6VzQCJDRygHJIz5nE+hCdD2yAmZ2XCdDrPZ4NOOsTnMkCv8cgz+Es
W06nCYRa8nKF/Ye2TE+gyZRcxYidqdjZU+c9Qti6NI8wZe7NrOOdJHK4BEG8dM1O
eUow2uQiZGadhMIXJ5V8KGlwGB8GM09ax1EzJyxhZ8tcqKCcAI6NBWypwesTi5uT
47SVMh5+XlUx4DFZhcQaB3/eJNJNVBlTeRBUx07Zd/asFx+ILp3v4aplE/n8AW7c
Gf+UdTuwhkY2GKQDJgKCGAZi6+WjNPsRgljKeOnrs6trEOxVTSa+8JhgMoEZwh2s
7OmRvHet79fDXSGTsuyADJf0bQYrHQH5nx/OZ64FCFkQUwFHNfxKAxTZRQoi3Avf
3u2Tv58W9U6gy0gxwyxjtyiV236YvrXyVeqCP3zo2VxUN1icnHyGz3X6LqJLoTo8
y6t17ZOlwDXupc/ctl5bIsUve2MowTqH4U++4e2WdHIu00zRx29BlDL5JicrfCFK
4OiNyQNS/KRwqWFpvaL6KWLkktwVWtb4MW6cGNLlc7udo28sVBBpG0ZA3oX+5wXu
eEjISKg+3cgR68vbIJQ13LWE7oawvfzDL9zcLvqOmRiaKlgDaigOjejJHKXAi1vE
hmOEmSlfvwJK2L3/Wf0eBQKp9biIEeT8kg0kTRBqzaarQ9WGn3wwTEKtJzRR/QGx
e0EFeLRsQVuTF1TS5F3xQCLG1K51StsLj5EccwhAMWtB3BMrF09om2kS+6z8kpap
+dXXZkBm/+HPTqD6QfzyuK3EhFFWtJarZdTVjLzOUwDpepEGj/CVz1hYne2uqdkc
gIMpqakTvAhNxVkgthhCcb4xrt8vERzsvpdC5DEuXovKQ7zNvee/l1Th9LqqZ0HL
rW8yxHi2NYOZDyhcYpbm0fPV972MV1JCTk8XS3KOI1mOhMmjkf2+U6ZKA27R9rPS
jwp+m6114Eg8hyuwWzs3uE3i6QcOf9LZXszIMjHB0uu57oDeWrMALyccRDxKy0fd
7D8BZ418Q6Tw9CnrQzqK/SCEBnFSs5HHc2Fy3Ywj02efSCppNHxXOp5rCDW+xLJE
bjJp81wHnUQKsnu7ktcgSEzr+kxXc/7x+KZAsT4CVz0GVnnlIfJiG1Y1feLfstJ+
vZ13ThHG1PF44w2WRDWDzmK+w0RKZLPpS9/R3SN+508Ssiakv+A/YC3n5GC25s1H
GE/LArKHq4OynALumAjq/lEsq3TjHzApfOUzWk5gwQlvfrJOuRIuT7uVSd6Bzduw
EZvqfhFZ/3n+5ugfOMg1OZE21Tp18OGepPXy5rt3dAWezr5hmHVmaubJAzmg4meM
+P8pCQSfVm/ElBOVw8rcREASf3ahWtC0Df9T6GUNk5JrYfh/hIwarR+yB3clSTLg
P/7aJht1A2CuGQkii6O6bCuluoSDHx/R7FLyBYqIovp6s5cMPbsc8gLk51bpy9zL
fVkFQ0TCDMg9pvh5OrNACzs8onajYpXuEOMH7UjLV0OjOzR21h3kQMVHkBK297q/
CWLkB6YDik5yfYuZzgXnza9+t8Kcp32xGy7vlli59S5uE1sjiUamjYHccwri6GK2
Vqp3u+HiRAVGZ9S4LOrwEBWXGG5j3qfrlZ3eyXjp3gTNiM0q9jhD1sHeoI/6ri0d
51C7o/dMPRn895LUiSc55XNBScQv1cmWXke4eTrj2kDiltGWiUEhuXNKzmgvlaBA
I9ZFl7E+y7eqJHg4P4rgJJ4bFGGo/nv+tJWT2+B4H7hp5GYhgTzAJx6KZd3K9FQO
xLsZM7IYo9iv9TGES11LNQ+AMDXogEYEBkExOK1TGKEavmSvL3pbjHQ7LduTHvus
JNseN4BL7jxV307lRwD8TuhSKZczTCANTOeuCE6a7O1GgjNurMX0PLfI1y9sXiyw
WFwA//oJGccHI21wEGHAWhYqcOVTnel7iXi5Qp1FeGfvkJgFZBDNFv0DR7xekEcb
Z67YdJ1Jb+HQXV9YDu8oLsCHihymCvAk2Gfzl/VphkComL/QtyAo967DOd7K5tqB
LDmLyLiBImjzJM2PteH1ompHlDYXnRU9Vl1yGkEIuqSDpgU/uqGijYdebd+KZsAd
Wm4XahF3imsL6qKExChB5DhoUOhg4PL8dblSKsApZkDcHCFEZW7faNdK8p7e+W6D
k87A4l2jPmI3Dbt+zF7JEk3+RA3Qz9/+Cese2Gs7xfPCpOb4/zhhMhfJCotWyehy
0rMJRqJbRvSJApp06tJaOhhpSgzMql8KrpjdcEQG8JC10PTR0H7thZDu0vs11sy+
9F65zpW2gQejMBmJiaqG0kYOjDGKEwyfDehEpbd18Hm3+rNWnOXxIJN2/MD2drks
2ErnST7Nb7DkAnCc5B0yIIrHa9487f+L8ijd+irqPK/2DXoPoPbuZL3+8oAIyQgB
P7PXY+8C6XWfjSlNm4DSE9pXWgb7szrAAM0/78DudVItlHCeiLzHBhdGeXYjLyz0
VsTwF4YITWKju+VmayUAaZpoPtkRU7Bjwoo2Dadl2PLT/Mw2/1Zx81aS4sDZF6YD
LMLxruoMp0mOIZ4+StS11J5s5Zetls4m0wmU0EPJaMwMlUFFdZ5dbTtF+JMi6it9
INvl//QA/NALJ6eJyKz80wscbMS4qErizvQBUZXJLRzzrBdqxXbzsakjSHK5qBsR
4zYVW3nirpdYj99tXeQFyEdBmMXM5uhpWohBRQqUYUL/NYwsT/32bz0s/ZgBS1J5
jBbF2nXnJVCSJmCfwlysEdh219+NPoF+Uud+0Xuhj0gUOV530Yv8VKdtzVETdMcZ
1IKd1YImBRJRnOPhHDCHYpH7PcY50hs7LdXalS335eY0hESAJlbc5FvKng5GUkCO
`protect END_PROTECTED
