`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+ZOPyhjgpdDjYZfkxNaVr9p923T9Cb+UOVkD0QqqCCCkBm99JTQLXAgRRpNQaFlR
icJaFE46mmNx28Zg8ebpUDJmDBrdnMq6dV/Lqzr+s8e0Ja63P6d9Dchk+Zk+lxWI
KakEJTdG8jGRdAxomS6v5P3lHyMJK5JwobW9szhYQEpQfxFmzY4xGFaP5mw0rvI/
XPQ+5gnFoHtnLgIDMghQ8AtQn+ccBzMwwOg8Y5i/Y2GjZ38Ug1ykX/5dyH2N41JM
DsZyk/BJPGOkfon99uZ/n6MJMbInPsy/flGkaeT/pt+nHxFtxBd6m/tUfTlrg4V2
ju/Hn1XftEsupFshxsZze9dmAHvol7nFBhpXG3lGa1eeh9r/lwKVO8JuT5Ab06/o
uwLQH4wJyNcmxN2ydCKgOnVME22sQUYTbPLRh95hAZcC6aUQUAS06Zb2eirU+bnD
3WQVbul4jnhYUveuATXv5xpHn2OILE92p6qZxAORfc1o2Ne4+wqQFc6ZLKo9nIkv
hpuzEfA4Rzci34NdClXIJXPEYVIoTkKD+a0RJ8pycUuHqX0CqLKOTJjb+Yhgtk7W
266FBxi/shogot98ynYddnLLvmrYlwuI/t14xUv1I/761WepgiWQTuRZdTNQo0ok
Ui1r7ayjT5XFnGywnrXy5luzteJBpdBvxZD0QriSdi8AY7SW8x0JpOTSLwLXyKuE
l4d3A/1anfslqs6nl/SnKOZP9pIzC5jok2vCTKiSzsM+PZYy8h5t0PpJ+QWtMJAD
ueylAT4q8f32IHVECfU7bvjrRbUNLZX/1L6wzUCSwhVcY6y6mnzS1uIY7gUk4kPB
t2Wy8vwHrmyolgTXT3t8wQFuN3XDaRvsHIiE02wN2v8aZQCLXjEt31ikHp94D/g7
/7IVWRPau/pcxX4tpDq/JLoce/hplRyoPoh0fehbitZ0DZvj/dMvKU3/qkfEHPUS
ebf77apx9Y603FnODt3L3w==
`protect END_PROTECTED
