`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGyqU/2HEc0uzvsq5Tk9U50uI8KelTBBWc7lT2KFBnVg
QF2pBWNpIq/9pjPQ32tkRviMHWY8UNFBB9im6PpIf8AFIVRT9+S5YsQqi4F0owoD
p3NaQ1dvCaAnK2t22RFsGMA4t6192m8sa1q1QXzBDPz5Bxw19xUtwD4Tl21TZhbb
JtyQKSv9GDdGcmhtzLoKeYx+YSDk0KWimsML5mh3tddRf+iUXq5v9OqP1430ZMBo
`protect END_PROTECTED
