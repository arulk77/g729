`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
OyA67kRAp61XLnSvP5JarMkzMfm0ki+RzecuXUngooCY4wjsR5eQ2cN8hb+ltSM4
G0GxgAUkXhHn3NAtrVrey+iZIZ0uC/K8keOaOlIcbb0uyPso+HT4y65bkgSzE5S/
GeLqJAh9xV97yCKWb6LiN0u5NvKYqPcpbSZXGRytTptyhsxDcRwBD1ubIvEFNd70
Mq9tFG6uXp9TnEPaXdv2CmUqCY/iE2cpWHh/yIvbwitk9mDq5NJ/3m8NZU1YfenB
OJ00V3fRmPVB1HAUd37ELntnYKljySG+akkUVG532cRzMHTfZzKRKG6OtkRjUCVu
`protect END_PROTECTED
