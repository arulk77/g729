`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCmihxLogRxyowBQqaahjyeahuqDPho4jryd1CJXOkcK
icLm3cSuo7PwdJThWRGL8aXF6bUugPSjIibPLTWauTs0yexKqkNfJTcRByru7WMd
M6ZeS7NZyhLd3oVX8ok6zOxrtUlDNep78f/71/g6eoAwm62bd0kA9CaHw6jHcPZn
gtgZrvgJeQ7TFp+AVa7FaV9LEhctq3i/cmnZ2ThvJvT+j1FpONCvlJsct329fhAG
h0l9uqX1wuQR3CF1dPohK7gIeQhvDPhPx3zBAxxq1yOWiqe7MxfvXdnqBP/X8huj
znkfKntwDNmjAjLT49zLUZak8Kkt46VB7d/dImcHjLiYrtRXcruR9tnQ4pSFbxEn
`protect END_PROTECTED
