`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD/Wtzu6agzxKadgrl9pK0riOmPqjueUbDGhtodBsljx
6r76e5KS4Hb6QfngsfL9AM2u664CAZ7l9X6PLH2UGf8eN8HIddMHVfj3E3FSbxGR
czhaKK/poTz0uE4teBqRwzkTsP64JYhiVB4743GF1llZv/aqJbN7I668I5mCZcnZ
QQFkgTB8WBH3ph6GhEcPXhpS7hNU1LVEKuNILEsXG0V6TeUNUUfi30H7G7piYL/v
tv5KtLPmnilHq99oRksfK8y0/r3rndXqjo3jqUkZOM7bvfphFdw6UplnOh2fnApc
tkU9QvYS4iJ0WlxfYRMIDQ==
`protect END_PROTECTED
