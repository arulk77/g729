`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOmbj82rBnkvHO48VAbOIm+5/vOflqPdu6ee/ee27iQz
10O8edOpB7cUqVcML3F/nuGwTdlIh8aNh18ozwYYI/ECCR21MTADYzi/87bHb7hY
eQE10PiIXd6yGC/+mD5yYog+TyG1NFRJ8E1mcPhNOoy6dYyJu/QYiU5hA1mVIZhG
NYND3h7SL1/y7334c1Hyw5fGBU/1xzPM5L3ZkoqqbUSFvHonn7c4RKpj6j1VIQYS
3BwTO9Sl5+OeskBzlm6qxuajgsaT0pk/UeR+NBUFBaMbJp11x69M50IgMVS7tjaw
19gKBwuwbjYbxSZ9JkQVcPtN/7Tf0Qzd++nfbB5LGbqAleNe3w58+jszGPE7yCv4
`protect END_PROTECTED
