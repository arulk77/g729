`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
f11uP3tAS38J+2XEq2c6cPypemmtZ8hKHOfG/4zRT8bIkSyyGqHY6e634GROsDBe
NhWVa3zEuuP2CCtT6mpkbCXBvspnECybLLMmCzo4mH8PQTPu2nPJxmhDlvi6dWgT
diw5fPQ6N3PpBY36E8gCh6xTrR1J+cF/or86Zo7LfNgoHCmMZjVLmVomlf393Qgz
`protect END_PROTECTED
