`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
kBu6TN0hCYMTRzKUrbhWNzvAITgNMwiS5KPUmpZen75vYR6lacfC2GrA/PGLZxKQ
/kOBU7T/wWOTQkwj54ej3mPpt7rAD1ESizPLzRmrFGmNN8iexcjHU2omOzAxyU4d
h68Sde5RXExxMniv5sHmetJVC8VbqEbw0uv6iND79CHoOqRvK+W6wGfnSMfx7vxJ
PgB7mS8cC8G7duCMzVXpnflNflnG+dpNzgJ+oKdZKZSh47o33kSghMwmdt5lx0Nr
D0Qw4F3iyHSCrRFBhzyHnbWqICkBw+uG5eOufP3xpIk=
`protect END_PROTECTED
