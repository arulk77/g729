`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDde9jzrnDMhGxcF/x1HUls6FmdBAa6EKsctEnCHJkDe
EZqp3VrmXQwW8wUABXhru2wKgGJHuNJ3kj29Tt13q0/hqGKebheMUpoLGsYeFez8
OjHJivPBFPgXREuTdmf60iDSDAtEBLVOL5osMWEj4Mh/pxJGK1YHH9SbbWD9CQAj
6CIN7lFysl8hhc06txvzrg==
`protect END_PROTECTED
