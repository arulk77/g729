`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCGUcdcgkkVAl8cQ0L/gAMjHT742wcBz0O8/4kRNkGfx
e3nA6Q0B8dQgYm80az637VS8rGo0ckRXLbZ7e4EmEfpIf4r9t0wzPvTftiqA6RBq
v95iWOoXgHfkeZ5+q82fotCpd+GQuHtIXCd1n2wW1/NB7+BvWl5CEZZpbb98TFyU
gYPo0TSDEB42PbKkRywgxcIiSly5dAO9jU1WTZlSOFVwT5tCPGd4ecpPccR9y9S+
B/Cc9EFHV3gj1hxiuGwadePIawgjlbB3SBy5aoDSNYCx24ADPMb7ZYTXbrcKnc3d
`protect END_PROTECTED
