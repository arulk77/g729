`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/ke5mVxZmGT0nDRzSMSlf35cQsJJK17AoBsPjLtdz69
AOwyT0LC7zB6CfZZKjJOPF9hDDq/3AIU1pE1NCxxDKdw4rgS1GwKCXj2pT0KLogJ
IC7NrruIBWPI2v3io1kgrRrPCRVqfUOOOZHHOpy601iptMpQu6ffBWrrYxVhclhA
1b+2KkUSoa1cWmaKIPPOrr6Jd+M6YfBWdO5oJbFj3F5yCZp7iTKkLXdHjaNXwOkf
3WnQVjN8CzGs4kvBZVSkchsZvspSLe39E9I3ohU6QKQ=
`protect END_PROTECTED
