`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8ST0ZGuuvt29PaV5Ici7UBTjoZXoi7P5/HO5bvMke6vDy
vW/tvBcshKKu3/XQtrb+oh5J6BIRDJwEWqDJw66QjUoCo7jCC2pThThk7hUauZu6
QbD9bN7gu+rZNLF0t4TpR0nw+7UBd7HIhDXUGEPP/QHNOF8EA0uwjapVoI+YGDDK
R1HRlfXyeQGoE9i5GWjIrxopAhucD5IQxHqJjZ7mBKFm6pgMAM18TtqAsgMnryj9
c2nroufh9x/KWZZzKKdjBqdDmlhKDr4Gt4r0hLr84LS4fvG+lYVoiwwegTVbQ3pB
gylgjNlmg00xrq3NzJjeiyGhZhwWr0iIaK1nCzb2SVpTBG7NAfBTJ28eGw81jlsU
FqIjctAsUrYjaqGAodNnZu3lzxQDkqNqdk1YKgiWOGG0obU9hqZlfOJijNHCsnr3
/+iFh6p6lKOBwxvHeOBYxOagDw5c9KWViuqN7ybhMWRwim9MJ+w8Kw+Mt2cJcy9q
yBqsM/hqSYJKg4qN8c6mqxf6+i/iAgBxpkKkhS/3p+Cxdp3bXcyTln+/42s3Ecgs
PJTEYqk6Y+aNlSmbuIE5TuM8vORJubp18lSnGTO1phxMEUaZPD84vqBu1D/Xx3+5
BjcZ5N0XDHmFiCmVP0KTXtEzFXuKp5UFJaTEAIhx1nCDMLUq97zeR0cLeGIZjM2C
ypSQuSQvedeZYVG42mu28Lkii/Zqbp/pedDqhEIimOEJrFUoa9LtsGcN6t/ywvQD
aEq0AzVYzvWChc/f4ur730coowZEUmLLI+jdjSeumbqWk8dKcBU1/OZbJWydzak1
j5mHo4nuSpoXwyQJPO5ptWdYApubYMrmx9AyOqLxXQot3gz0WdByChayHN5Plxle
`protect END_PROTECTED
