`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBU8XBtLXda+LsMo9hqm0mEfAXV/UOlmrhtnTjgC8Xsl
v3nGCtk2hJ2rSwiqgNSYiRA+UwnvluDLShos9MGHXhVpGBgocbp69DwYJ8tJOYSB
V5R9mDuUCmjpz2V0YuTbougPj3EUDXiYPUlxJLdc1iv5y32T9uBGLjxhfnk9rILf
CkjESxUPNlAJH5BQA8vhPAV5j1S+LQzsTVl8LZlYjwR1TkwD22X/ie2k0/2G1Gdw
rcmd80axaxWIb5ukKa3RE7bZKIAm6uWWba769PX59yVFiyUD/yJWE+rL4LZfJaE2
d/V/JGniqhFASxHpDnwEXg==
`protect END_PROTECTED
