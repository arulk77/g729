`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
TigNQFGASyXVlCpbuLpwoe3ev9iqGJg+sBGN5nhWHpHerdehGlALKIik1tFhewmC
RUQ9umKe9QcEGVQucuYKk2F6tVDoTA3LvCBxLCwwLYWt2RmMzGqFwq8A7Mpw0Ci1
R6kcEnkMOih/7bWuEjgkNlDpx4PNCU4QUlA34Hy+ElbRKn5W9Epxs6sjz2Is1yAb
I4MmxD4rxhKu7TiuyKB3yv/PviZ1K/ouO8VLDtbWnLCp0SiJpnkCq31TGMf/5J3w
Jj8CTDh0qcBNbNlSNrSOWeZ0OTZxCKYolCTuOQJwTr0=
`protect END_PROTECTED
