`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMOC2LdR8xh//47YKg/ZvWDPMGK71SvzxmynU1XG8rz1
W+wiNdlsE/VklYiOobf/2GzV4ADyW0pa+3/KKRrMhVks8dgC/kVNEECFMP4oU9Ct
AMHp3KGPsA7ZcCLkJLpUmA4VLA7YyzHGy9+TVD/fHZ5ZzmVj/myc3H0sEJgoBiLz
++IGfEOjMfGqC/bVUnZviTkjU3+hnbfBVqOaqa0QccIC+i/Q9d52EF7Xjp67EDB8
oqrWwVumzgc2RKXciwZlkXbx3ihYZHaG/em0cyxo0Oem8AhchZ4W4OtAe6ZW2I8M
bx2Svbi6LRV8BTbZNIDRJoF08GxBSul1df57h2EjSM4GnzkKZIkPenWpWS0IN4Y/
22WK9CiKiVLwvGwLrqL+usNTmVjTjBrfjujpuYU+v/gbv5RtpPv+DLYCU+La/JK5
bNrS570OYWVrSKNRsXp0uZr0DJ3ZC67ntMVueJjcsgz+LijhQ00zN5VBmSyF9EoX
biorYCEtj+qp81WXUoZIkhpTHmhgiypE2rdvRmXomGT8qWplavhVxtQuOEWDmbKj
5TpwCZW3f1ET/Koyyloc058gqtkt2LmoX2sJbh64f74=
`protect END_PROTECTED
