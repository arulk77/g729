`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49JeMZX3ToOJf5IAwhw7+I2ED47cFz7uRumWb9+z9QhY
e1GpGgw+UX6MWx922R83fxu88Ur3vPUcK9y8/YRKbzzdYpqbvZk/fglqPKznPz2d
57oBcO1GwUu/LxnsNwlUAhJy9RzA5IvJx8efMCBUT2qQUGvkb5AglfgR1Xu8iaN/
zyKHP+p+ZXRXpy0fVbCN2UFVyZ3l71b2FUnYzpt47JyTgB43FJK3ZbFLtEPYt2UQ
llGm23tp9QZxSKZrw9mPIl5eBQ58lZz75qfYhuqcxL5iTrpLEE0en984aXXKxDVy
FAdPLQ6rNzYukBkHGX7a9yVwDKJOyr2sNYj7n13eOcyVxqoT/pUI54j7VKuXbHmb
eJRMzcyGG67YIUKOfLZQaQ==
`protect END_PROTECTED
