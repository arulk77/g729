`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEFcnyDsesszsUWCMT1RiAsxpMMRZIUDGyVKyo+c2GcJ
vK85fwJ6np7kY1n+e5Tr4k40YgkpLVQNNXQlXGGuLkZSH1wWTL/DNZvPfWKDYRH4
mb1zDJOlz+2A0lK0I2C4DUN9hUe2WGKKwMLYjwEj1JANMqCrRLTtOHmqy4+DP7Km
iWD6zuNbMk+6Up7KKIUguw==
`protect END_PROTECTED
