`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C4YXz77FJmjcbnitRagvzIe2aGVko7MNtVbtSN5KgPdU
ulZAjo1Ce+4kCzc0vyg8GsGhDi9ijPcD89WydtgkgHJE2HtN+AxQuZ/RNuf11Z9Z
vz+k30Ge/jBKzrIZEWrFxC9KdLH1OUWmQb4Sfjk/CEScR2PVneCrUvmOvZ6dBpi8
2jMDKr9lfcG1eeUzAu5nh/JwC+0K6Frc8GxqapRqWXOxpjz0/ccGrcI8AxJNw1nH
BUFJh2eJ/PUZ0cvKMVwxpfYqTcxCES7UJEV5siCiLjjT1LRQMIRpjh084or0scuO
X+SPrYZlZtVn+akDu/E1ANwqF4yKlktRkRhU1FNipuUt9g8CPsDzqK5WG6m8oDbj
Rww9IawJuztWviCnnWF3+zSn4VquJcx2qX3XxySJhUMJ+fQpeW1IkWUX94P7yh8q
gtMSBjXyp58Qg5uN2WbH+FMuQ+Ajh3R4NxOxRCYml5NXyGQW2CyYIXvqRi+N1Fry
sp2yC9xUexqf/P4C7Xi72MRPXZubUTi/QfklrJg0b1W4HtGRPGbD2r89cE3bUR+q
8vkLTRDjWD7lwTqPBFFUwMiiZC6McaEdIu92rvt4w1jiFIJB3MFAWdVZ2RYf+8Zm
XIaDvvfhnrkzzKw2pVWkMYDJvxOb3qo2PYCjxxsS04fJwCk+LItox5nOfBvDzox6
98xeRIl8sgSSRG9Gf8OQaJrNudYqlN3zNK/l1cGn5bT957VhHJpdbxz0qEntvwPZ
6CqeS5OC6kAUfYY8vkKewZCT5kDaJQvX/jzLzk0SjFi0nawLyR2i4fIygEjl9CUN
WdtqY7qOceFNRGqm+icgA89iqeeTOPOvrGtdioSwXeP4B/H8Q78iC1L145DqCP9o
7OeH92830quBZHTamzDCgQ==
`protect END_PROTECTED
