`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
o8nUZ3RsWZJ6ggEubvLbKT+Wj6LW7XjzmRhkSD2WWPl/+JHOJgBfdBo/N/9Om7FM
mLXjFhdI1HHY8vPGEN1PxHa26Rp8Xl4I+hkDYKvsaqbykzFa2frMvB/jTgJTFgQs
faypQ6GI1Zl8AX+QTAEyLOy103k5uNbVH3YQkwwiO22X2oWZ5jHLGDJPF+tFMLnV
aW5yiAvp6V+yutgAqqAsjZEPS72D0C2k+ks46hC2IxFGMhmr0uO4nF3yCz4ezAPG
t8xNdE7NJKb8LYJkEN7n0LVhG4op/2iS4kDp0cfAli/plcbGsmlT/7JiIBwhut5O
76eWVPWeiwDUAUpD8aChC/U7MgsMkQdLak95DCJCXTkF1wq7Yq5Yc1zyLk6ac9y3
4ooZKaG5v1W7WIlpF5Br4k5rfZ6QfwSSntmC1JCZe/Q=
`protect END_PROTECTED
