`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
whfZdEhQhIVICrvn0VMg7u+YGWKNhVfFyLYgNezCXG+2VE2a6rkCFV3Kp/+hhPJx
F7sEsOTFn3Dxf0OFbRp+G9K34scvGy7o9jSTpukbsw4z3Pdvrbkw5NuJNrTjtlXW
lzmHKHo/1G/q3IpjXMj9wCeHX060pji5Lc07b9RULlrQAQh/ayYWvW6bw12Emz/Y
fEpoe/tnkbJBav9PfHBOvhglCkaJpKK38DDBVtrqjCCKEDhuWJMfmsquI1h/+8wN
k6LSuZ/jrVBl4XDapKnMeHofFzJ8zNJ5/PlEdW4G+v2u5Nc9mDlzOLTw4YMX9exI
`protect END_PROTECTED
