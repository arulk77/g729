`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ldTs3hSJL9bXEh4Hj4qnxqfv6wMoMK4SsRBwx2Sx43uZ0OEH7asJpdM9ln9XkiaJ
fUBNWdv4tEzi7mc9c86L48j+CC9h6t4mpgD8Tl4gpGNZPLzsAo9FvL0V8smdlup2
WA4S1q+K66VMHIKrMmR3aGrgrseKWg4rZSiP/LFy/tH7q26bDSw17z+dmqWOW0Zl
g4IeJ85LxQjc0EXPcAv5bOUn1mL3koONL3Qmmnp5abQ=
`protect END_PROTECTED
