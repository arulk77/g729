`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB5sqr/JmsqhVkCm1j0f23cLiLHKPQzuTlLnyKUL5Iv4
Ye0Rmqd6JjLnq0QiSD6csd4e1k0t1Ipr8hdZNZlVoEVO2N78JWtGB95VdzvrfNm5
D/Q2lbp5qd2qa8V6v5yybfhkOc8sNcmrRgC3mY6M/iNWcE5q8dlxvMcpfe7F+YZu
4qeAftMfqB4LgiEglvEWkIoetVuzvseyAyK/6Ci2mPuRt4Sm0pTmd+ZhUa4oC0xd
xUT8dvD2lgbhORkKW0484SKz5O/mMqlWtD23MrnNmnMluTs0UMI1UQ1NRbfZGxoS
MShbJl/wDiMYpSLZcZERbY5O0eg89PmqpROBVBLiPmbRlEFieds8ucbaF2Qit/dh
cy8ui4gCcOQWhzzgBIvFs0/VuuYMW/y4yDKNUNPpU3Ati/u7XEpPnux95yl5+EHv
EGOwGaWEqd/5hPTGw2EkvtPCXrAn+Ex0RtQu/ognYeDxNS1arD9Zm6oov5tPOUTD
Pn3O71SaXwIcLcdJWoqCSkJi2dV9fc2tuOcj7b/206lmXPFsvSsdgGHFziKNcIy9
aLFYNRHFfGKwiET/8kiOlErDWkSaDeMFczfM4moZcet4vy+8kQdGznp1/EjX3V+l
QQz8ryJ8E1HlUMv5PhHV0OYnUiAmRQQqbhXAA8+3xTbGNt7ONaAr2A9mBLaPzueb
ZdR/pdwaoSE6rMoSPI2ZsqeoW/ihSjdIXmoP0M88RjZqAIk6+BWQ6QL0dBBA1bM9
Jd7Q6fzRgBTAcWzSZw8oDGnZDbX2yaOJT4ri6uFYSfRM4CKNOS8+OM7rBPsHpqZI
PpmZ8OSGfBoo07LPt8SJPTMgpNI1weYI6piL/z9jTlVdkMheD6bFcMt5j+vsFomY
Mcx6BnDvEGTATrogkhS2mPtTafVUUcMuwKEO/nV7sb7h+Fp+ckHxrX+c9ml1+wEV
2gtCP/CaP5f6RJ4b0O57yQrPbERLwFri6rMWyOaXOor+Lmew9T4qKwzRs6eyqCze
2i3pCsPDk9f33+ZdYsDsrw==
`protect END_PROTECTED
