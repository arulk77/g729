`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCRj04nETYQU+9bSQADJQiA7iuS/mrUZznKfadbHMy5L
/aPtQuGSk3md8ookKpMAXLMDcgV+ufApvhNkqgDLkzVBdslwN4iV9AbEjdCLmZOO
pVX+8tJ2kx6Eran3qVqOvLyiKIHI81ekOIRMLlWIZHu1THoFoWkoQHD/1izAAdIS
WlGkG3x17sFGVSow6LPIQ+CdcQZcBWL+Lhl0QW3yik4AsUHC1aohqDWHFAAUxppY
dl1uDD4t46gaSzN1Wan1MKWqTpo9C/P+hWVMG9JeIMko+spB7fjfPCT3o2H9VKjW
z3sescoLf4PUUb87MPA7UKTI0G4mtHt11MX3ENLrE/43fyolIfa7fNsASe1IB6qG
V4N3jC2NK3B4iPwAoA1cL3GRu3pgts6VOHUFguxiloTDnXzB2w8npsgIv197gP6y
YpDRwmZojBmxvoNWs52rGi7bdjlYgmks08sWBoob5fRnVMp2gsTlQ8IPUmaDLuAB
SPB8UwU1BVD5evUMUcLTEki7XjhaHOUdWq9W8d/N89Wp13QthoTPM95eOHCgL3+C
qTKlZqnZ//+TmJEgcTCmAOa3ShsXWiKCB+ZEo5X/xO8lIa3VO4HgMlwlRcaYGDw1
KVwYm9DJH4BY7hmj5zl4ibJQ3cMAIUMC38bcDKs9c/f497Euj7Zib98x9puK5uep
5bCYUMBDup3efuL3Gecc/Z6XxE8tlhx6KJFWESwg0wJ0q4Nghis946pkW9e3Jzl2
M7TqZxOptAygvJydHEvDOyKQcpUI7eWxxXl7fjk8DzIRG+U3iFn3/ceMtfADt0Pe
+9G9hqUPUQlmImCwYynx/pag4vj1TnEYWL/UJQy+Bm7Op0eDDm4oo1oizLC4LRGF
RjdTM8Xs/1TLHyMgLAu1Yicf5UFWL6ishMQ4E6cIEDaGngHSzSESrYVk0FJ1vdw6
w3BBdKoLqWf2V89ATLuzvg==
`protect END_PROTECTED
