`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLLgDehWIpnKyL6AdNfAh1NgZzTRGCehKlNbbGwjPT5U
CnKwhQKJTyYO5JMOTAU8k0YUdPMfU8pHLVLVZaYTFpHXxED5+G5IymUcoVBYzuTt
VrBXXT+truDDH0A4Pvx1dR8VrnE+cJ5bt/xtP5TgKatvI3jDEUisnlV8wR3bhPlI
/dcClo2FD/6xi2WZ7YaC/8/ppKpbg9ic5ZuDvEDq5tm+XsRhQrb44j5xeUnevXFh
7nnvOVdaw2UVbr7P6KRy7RSf023EYcfvdR12MdjHjkV1mocR8y76FPMc6dsTLU5f
Sj+1n4i05/OQ5Q8JTDb6rIkaBAao+QvHeHPDwEYhy97Cozas+r+9nWfgQc9VJn2b
TtCM9sNauazlwEqEf85IvTZXdNI0aHUAjGTSihsNazJEexGVGQq4kuqZImF6gdaK
cDfpkWJaZ+cuFuhrVf/24TygIQKbtOvY/c9xqEnQDxVhz40+o4x5SxnMryT7JmwF
jLHQogExmCJgKGSQesPzbulFahA4ayIzkgmDpGtqZeWZGi3djoLc+6zeCPMYkyfW
mvp9wTWTDMWnIuJcfzPY9N5FfnR/vQKcLrZHWWE6nqlOuk1xozCfTY3P5L3EuWCE
/Haf5/FokSz4Or7BDC0nOBiWuzEWPs2gilpvnv+pAzy+AX2GQzMbbrhnbwnymrYO
eqIja6Z6DeJnthM2GLfqn500OVzpP2dsHzw0gyG4NgNs2A38t+tH0FuRiBYS5JwE
AfcKwCYa0BsokiLADkHRjfECfrUvu4MGAOfVEiHgK4vBdjlyo2kHAxCkvzOsM/Pj
AdoxlxWZrPf+7POv/AyhIalqPYm9dtfmbXGUZs1m9Os=
`protect END_PROTECTED
