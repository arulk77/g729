`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLxZ9D4YmORX5V8ACcBSgH30hNDIEF6J7ghBf/918HIB
tbofxEqv//oKg5Cc4aQE9evURG3ohr7ZoxrW/hHE5Y6wfObQ1lY2aKdJfLCMwBKq
OLMfNU93yKZ6/MZzK/P4nKtEos47/9W9oTmMtFg2giFhtPmBnHbns2h2l+IzYaeT
OTXPXPBwLXqcxiZ1V9CxwQi0kTD7ANoxJ0bSdsfhx18urXBJE9RSAETfk5FC38ud
M3shZQpSoZEf8Vr/WQU0BmsyrkhIwGJDtPA4+rEEPG8SKX7Xzh0SvulGyRX0UwZv
5CblLhf9JbRNq9/4Kh0GDWJs0pyjAV3rPJ7cY5gE8VL8Tuo8RcA2htSiMEXDBjNH
HXA17uF7Ma6fZXtV2SgHhg==
`protect END_PROTECTED
