`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JkiMS/Y5+LSPtGEM1ItJQIvk9XXENztC5pUewzzEHYQNcn8a+PFJP/Kx2D9vzkIP
48obkhs2O0h/I00qz4134Ly33200YXQpcZj+i24Hta7JJWMPP8sWEoDl228NihrJ
WhfVHNyP2Z2XJVr65tv6tYTkbkcKJ+ctxx0jYh3rsmtSbY1lJ62skhd/RI/9Qpd9
oxfDYft5BFkgaD80nA79z7QMb1Q6l1MzSL3vWkzL+1yzevyB6zoCptq4p0IKm7dK
LxVBeOkL2Y5Rm8V3gyqICFV+5R8aZ8zRjooIoJ+0klv1N4ho+rkV0NAOvt0Ni2Gi
AsBgpbBf+BCOnaBhP76odptHOch7KetjeoMolfIyaCM=
`protect END_PROTECTED
