`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD2RADFSJj0X50Vm/h3DIT0L49749/LV+qXRheoPjcP+
I4179ycMB5gw9IeCZvSVfkxg3E/68XfXorm12q3g4FJckO/Bqs63K3fnwOe8/mrz
NziyzhErNDyu+0Jxl3xMMzRssMOfV9oTTOtO3kD2zGwyEBUnhf82qHE5nHCZGAxz
T8EqSPlyQxfEpRbp2X8QzIJkIlDAbPLke/OyUif4jnTkOO0qjr4/2Z1aX4tio4g0
`protect END_PROTECTED
