`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
XWXO1hTk++BpRNjmp32+BmGFRoLGgrKMGLPNfRwF4Wl7fYUKv34pt2o8weA+U0eM
jLMX1Z0GKu8m8u1obuEz3PxgxUGurrTKKoWry3MWe93Uhs5f7KgahDG0VdcP1TSI
TdWQ26J3E9lIEhmgDziTosE6eIh/tOD4ORNo4HFiGDF8nYc99us1pMTFoys/fyt+
SmesqqQJgEXhulxccfGTTn1gAEO+WtXSBkXpoKO949YBGWTuEvRJLe6r0is8e+Bd
JiYj1HOppmKJkRguBZzuXOaxA3KQ+t5EVUy/UoEZytHaMfmboE1ZwrX656DG/cBK
xl6hiAjbPePyaAuw3ij8uOd7IFD/Zj3PRviWOH4f2gwR15cQmgbEn700fGVdNP6r
lpr9My3avuPjysM/+VbBrAd9mAIUx0/aP36cry4OZH3YNjFP+/e64J72rarcyZ57
Kec5EQs0i43y3FkAPLWgZUyfpgrU9uITLi86IFwr1tY5fVymPr09Ku1Z2HZ5vZDj
WwV4009Ied/AvXEgF3Iu5DlcFLPQxLJfal+NP2d6OCBTFJ62idBruMPawvBrmQVR
LbY64Mw96+3KEKl1pgFma9UQgrE4Ic6kxwWnNHwsBd/nY3hXLzHdkyIXSOZRNwew
OMGT0thom4fSup5Sa9Clkh3z9hAv/tnJAp53s/SNjjZ9b85qSqf6aKYGjFe2Wc+R
5/tW/von01mm0ACgJN2ImAGsRrYvnNCK30XQAXESyoMldCwTfid7nTbDwIzGRNWl
/P7a4BtyfQD+M4T1RuAlizlWKzpdlnogiWxi+ll7Eo0a2m2jimu4KSvNHEallnnL
OEmuO5lcBJ42klqY9ET+J6vNkSdry3ICioc1wP53/U7mSMAJMffxLclC73KEhUwW
BoW1VThaeFK2GIyLcg/+hHC6pjGPsCC+FqV/gyv8b09t42iVS1vqoGT0oGb1z9da
8l+qbnYsaCOHKlfXwAE5XU66o7NnSuBZh6tXHr+QQQZ0HIIISPIAFiKo0kMkEsDX
12Fny8CkeDNDnYvKlfLa+l1erqRXsZ1+Vr8hzRY+o5JWfcEL4JSVSD1FkjwEKix7
DgTLa/JBfaLgOsU9UZnVWdtAeYZhPxASQgpXiwvb575A2Sn8HwspLduqK1qSwKxN
x6sHlJp8DEfJCDZAIJ+deHo5TNH165SgX0ZZqRYt6HXNpWuD4IpUaukWkGO7l+Z8
i6yDOdnVcnbBAubIFupkLrnJnAdYfqnVEM9CIjqa9BvOUDfJlshjRWy4E6GjDwr8
ox9SJc0h987J1o1jAUInhRA/UHj4vT5+El4fGmIUp31Ik+Bc59dzYgQ1wqD9/5ve
PlTcEcCPRprGzf2kGt6jOosaBfBCTR6imUiIXCNHUIFRhZlWm3zrhJnAFnZopcec
Kxxtoy3G2nlkJWkZ+19hreYwbHKteZGIwISj4aIcMxpRgXCsb0PnJfnsrxc+4Mcb
YqAlkrJA1OJP4rtg7xH1OqEZtrNZ/ynLFJIyILJOcoflZAjs0ZB/f0mULunXK83g
dmfDbm58/WzwLD8p9msycdmoNpYw1Rx8VFum8RGCvyMgnaKzs3+uaw2ImzeULBJI
870HUzBhvsoeiVuyyYT2zk0uqqjZjHw2rsHJ27JMa9e3453zkRPJHYBLC5Ycvu2R
kZTSXr4xl4IApMCxI8XqgyWO/3glL85PbaI6L5EIB6popFJ0cPpJU+0KpBtx6Xvz
0axp7A12QRmWnlRkwb8d/lwVIyFYa7qTW8QkVcNH5laje9/AUOuwvEcLgxvLSxYZ
khhZk+hEJsAIFKuE+5ziFxyxslF5CXdnfZtKLN0eLNPfhhaNYt1QljtLXca6BaZx
c95Alf9rsT9yHJtvmK3gE78uTafNoReFNhheluKc4FhehPf2vm9hBN50OuJsVKrw
HGl2+Y2PwbouhgLbaZfOF8/e6CGxoat3GN6oeidrJf8lUY8/pJzl6/PLUWP3gYAg
ZaId1czHdli41mCA10sweZwzBnekfoJlJswOBNXXswsRnAwRkFyMGNJPS1ZP1ThY
WBxG0s0FwJiuUHctg1YHoZdkU/aGqDmBMubxBqqsQr+N3jMnlT1NVk84LofI9nZ7
Q4FXShTu/NWpF9ST16+iwXxV46hOE3VK/OLfqBLUna1xCJ52ypziwV/JhTCwBvkx
8QKh166AAkbX+eG2l3BZ7Lij194UKwWEGVS446SIM1fTD/P1jniLoeOl01U2ALps
tmGGtNls4telseqd9W67YN5wk7as3qBB8h+/4GeJzGE1pRTu+nEzd7ry0BVhMR8+
h+/b05ODL1lyAB0w+44f/xPWtQfpkJxKmFpwE/f8jL0pb4MVBgrChVeJG+DxF8Kf
OKZkRq7EjMmh1LCbXoK1FhVH3E3p9VNgDlQG+G3h8e8NcxixcvZ0r6/P+nxXD/qV
tuVZYpgu3rvDYP/o3furzGEc2ZsK4OSh+IIEGJdyW1GAkY2u4eBXeIQ+0V6oyGpg
XJP/3x0zwbyU9T4AyNuqypIVXYN4BZGlTXYCsEpC0J6YHPcjPNPf/lFiB8XPB9Fv
cW4qnD8kkGAYM0OgkAnsHDI2TedRsveOjrMWy3wxEewYpmScG9RWE4VNGx2VIhIn
v46nXT1hAN0LCq5I+PDZH+YRCXAGdmDlKjk00evrvpTie0S0r3p0AxVdYak5Ljl8
BwA16Yqx3OVdik26CdH8+ouWMK59SvCvpg+WBWShwWLbQcT81lkisQSChJyfReeb
cgk7lsNQKldOXbIZx3ywK0PHO15OyT/Mg1u82ouUUMjjDFDu3BZ9+wfDcCBxSIBP
yJI/1GUuds/DD8C+Xw/aZ7YXTYed/FpdnXDJJvo/GI8/oMfCMYq6YPyT1u/0k+Bn
ugIj3m7U2g0Wwbhd8LayNP8vBRnWe9a6HoNs8zG6phBnmJvf1cSHoSp8pWy50PMv
0BJusg6mtEi523U8MZjL646y3Tz7//8TG2kmnwWQR6w1yuyURxDMlUA85liVGDFx
xdnVEVW7oBpbPgUQaLCgHvBTih6qhSH0R+QK45oCJP08i7JjBg9AQJHcTq2g+PTo
K5+qr2s29p2qzv17Igbvn90KxVSyZCyYgOVV5XYtt7KO90a009WRRbSZwsuKhSH8
fmEv2YGPeC6iKTAuQoztnjSjSECPbPt6Ga1SsiXYkyCMcRbP2Fi/CsDL2bYAc2XW
SSHbtPq0JgoOptJTgp0Qf6CoxV6F4C2Y3kUVOniIBANoLYQdGKQOaqEHv0QwHF6x
45ndZf3oHLDeEGyGHkSh8f3yzsZP8qTN4ModQY2d+IzRK6FzKeIjfwCffcpZZoOs
FZUqvxgizsiviz6tf63Lduu0N5myTN5UjHFgLIKT9l69/Mz0ZJBYdoL1jyf2AURj
xX0osi1+C8tvBFDC4ErGnquOePKFJsyWuDOh3GNekbzFh1HVYLXrEt/J0hoo6In+
qgPG/v7fMC7K+ZwQFtfJ0dUzsqmZCvAsefjlF3uT5ap0KAdz5EFLdaEg4QeA4Swr
kkS7S99Igy44UO5OKZD8uJh0gAxTfMZ3u6MqB06an/wWBk2WoPwb+xLj4y/J/BRU
Pwz+KbrJfxPle6RlkTVmNkux1fcSrsUK6S2zPpnvO5qqBtPzyyro+fA5GG6J+j2f
u/4GTtahuNkkeI5uyS9SORiXsSyuzXmkfU5JsU8eGiNSqDB6HQ7IyMTlf7BcwwzX
mZPkHHbcoQvW7A96nn1y5MQhR/H2LxuHv3HYI0vInfEjtzw8eTYGzSpt9Q19ckTA
K0Y+ZIBS8jHhkqPYLVrbSe7i+U8O9PusIxuum3KSgaQSvhVUy3FPLdAQoXO1GwFy
5lj8qROVox/LoBasX2ZI1SaaI5dcKYCLuX4deIYvSGTQaNQQ3ztr+vVB+ROZQOcp
/+7uz95OvzX9aicmZCvGPwpwIxiE8mL76rkVYxq2HvOaI9VWSwMQZekt8U9vZAzZ
D0mmA6EwxvOlR4WKJeDJTcRMkppOAgBAdtR0bZl59drAcdM9rrfNQJZku6drt8ah
kFN/VxvUKWglTHWjeGl4U8CvtlxdTTRMj36AaQF/Azorl99Yb6weS63TiXChkjAJ
qywEpuL/SZvgl+MezXFMCpupRjtvYE+VyfqeiWFg7rMmnEMXszYUxlzxsLgspjwc
+wiX1BM/MLOmrTm7KxsD167jJwJwt1skOZPutHuOESJtZmPOvW9MZtts76Yv/keh
CbuZQAIGdDuWR3gJ/CD13IU3jUIrzw6MvxpjbkqsAT/2USbc3GhJPsuKumWbeA2/
q73UK4XrLf8Mz22lXw2Uuj9bowvz9YnlhV2bF3m6hUMQ4P+xyZN3vTMzOFDsnWTL
3lCckqdwzb21yBQ/yFK7EnR6b2xUxsmXFYPypl+UbbBZXbpg4Y1oKFefJlI1cJm6
Rj8lgirN6z4sqRi6dV2YcjrvW5gdoSSUPhVRJInWFrs=
`protect END_PROTECTED
