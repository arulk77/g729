`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK0zP9D/3neYNSWIagZnjyuKCWMicxXIeqRt/ySDEe8z
NsM8fz7J+z6HdTtYBWtFr+qk+1fyPaJUqZ+5gh3MRGQlzYRq5Z1ih0KMZkNBk1QF
P/oRfDq4YolQyEKPNYraQ9lYcU9OXzQVuzz8Dz8sfL9NUKvvwA+AotTXQPPnYzCM
Sp087f6tNe5muNuae8LhkQ==
`protect END_PROTECTED
