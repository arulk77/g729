`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFRVXsYVveYlXs2X1FwBZwd4+so94pTU0NKyj6gamNdQ
UKq0hIHI+1s3kRJLrb6ihjHyRC9uapI1Lvo9Pvm9/OShDKXYlwNxnV3zZwA9l3cO
OFdWAAItLEz/eJdWWEUEb5uSZev5cd4oUU2C2lATX5v0nTsPiwcaaIy5vo+Wtm7T
Ufyg3L1mpL/7An6trDudF0XZIUpymUn8yLtMJfUu5RvxM1ngH6wqEATdhUt8cXgB
NSIMHcLL7JWckGk7bMUg44VcYLdPZIsEmeFYABPTGJOb7PHpEouOWB9X0FVDnKlH
MxW6cbI/qBkU/Ag38lecX872Kj3GVjhD4Es8QXzPA+PIYOjuHugi3iW5SCzns+D7
f+bdCiw2pvCYZ41uFXPGUA==
`protect END_PROTECTED
