`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAY53AZ0jCQItfDYzNb6DTYKqNRxPkH3/wM4OpsFTCTVm
D5+6JJlL5ibgEbaty/eXhfqckD4tsyEow6NyFB2757+S9dId0Zp+VoRhjEah6bGe
kdR5ErLZV5DlSUuWyBmDuu/qwOB53Shnk+ihIPEtI3SyxjeQXYvascrpr7grKPlw
ZyKWhla7uorYI51JWucvv4ZXnohQ1gNdRJu/Ub/RMn9ftONQM1AFpOC4vJR0dQqU
ueozF4WYe9suW+aJmbE39lzHgi4gfqDaOqUpegu11Zimqrow4LRJkSkO6PsSy/+j
XGvLC/LqL7CqFW7/48osOzClMGlH+Ir1SsjwlvIP9Jem+0cPzNf9sYV6//LXKCmr
viq+9JEKCwFUGJxnmCe1cLQbtjOyxCF52r6Jv3tpLyZTdfH9jKpcQasZms70lEsW
ogNnWqpnh5019ahfjtZWg/Wxyi8I1gjqOYSrGYJcgFOac5pp114Iq9rI5RCpP07k
cujMGU/tAEVlwHQO30yDWNap/6WXLo2ZY9m2h6wee37A1Kf3fVAYdXAC8WIX1mis
T+Wa83nUujKPgGey+h8rNEMewWS5yhewhGWZD/rkWwgef9qs2g6sEsjJEcmlnSg4
92Xsg4aG8MnEmDRTSdv8lc9fsLVBy+VflLDhql9sTlCs3RND1+RHKWaMvdmv3Iy1
rEr4GvTRVrQBAh7xWyK3cawURZ9Ah4ZVKXlaip4sx+/tLTWHEVCF+vqAs5Y4QoyW
hZ1MHr7LOJxIQDpHwLRU0eOfEDPKTG7ttI81p0QjWsaIavt7Al4BEWxR3okzcwF+
+vbkFmAkbHV5BOMZhuV4s1yL0avnsmKjHFJp8dyjZ3yNE5GTXm6euRuakcpT7EXK
eQv8GpD+x8vALU746e0EHD+GjM4jzo5c53EyP4dkzReBvAcbqtFPt5C20Gz+sxTh
ocVYJh1D6bySIoyVZsyclBIA3UC+PVIkprEBt2Ne8h3G/oThJnya94jsrMX4nRjE
RHcaP/ob5mz5tfSg2r5J8UkzJjpu+nV8MwhE/9feJJCew6r/AqzzathpffHNzdyp
tfid37rS9WZY5lgh+fQ2y45DQ0/yqRS3BpiIoE29H94LbFc30Gy1By7Qx2vRrl8A
HkIzi4u0iQBmgccRvCDHH1pqmZMmgj8GFgSivTQSifXRDq/VLbQ8C/RiF9g9VO2y
Eqz7zevRUIX03YFn3icZbWL0+j1IMl0y8QNjToBDHD0dOwWmMzW1R0mjrAdP1roa
AZEHu9+4F2KVmqknfFDGLN9mhPvpbmt4Dm97mAX1psFS8OOWrLNIWUC/YgPtbatJ
lFRmXqexkGEnh8kqQ6BdgvfxqGwVTCpMb59L8gMrz71mZ6jFPD3eirKfHDOephE4
EoGCGeHxBwnos2LoWyTMj1F2869dlR+jhM05EsLGMga34rRzimRMJ4qhgmpeysTk
UXNza4qDMaikJe6dtFiwnMXakrBXgs7FsqJiXD/ugue1ioh/u08mnKt0OsLljbko
xbM8OZLyTk1R1/QdSPBdz2GMRGFvWo2xwPJnWrV/IudgDhP3JglH5I6UpG4fcTuK
NkpT80EG/eY6OOCJFrKQ2Jh9x3DdsZgZpRwT7AOGes5owV44qqfEuaKs9wwh4+iy
GMfGT4m33eYnuHQ6/L1WHin76734MbyRrXL0LfQQaZHg1kIQYdUkuOIpfmbYIcRM
kq4x5HNTKZE8F2zmKdGv3uPtSjpW39rTI/P0uaGIEZcvMVFVK3EkLESRrNADhb4P
2te46nG4Mle5H+g2I8LNpg1ITncuSzk4+oclrN0bTVQwSBTw/fexO3jFYaaAmc1m
CQXgdti3tZV5TXejSdfOz2n+vHoI25szZr40YA2cnGQEJkTmy7Xm5HRszxGPIaLL
0uI0VR6Js5vK4x2aAIcyY6dhovUlyWik+HHy+Ks8nMH5l4+IOwsMNqpXcVV7I7gK
LcH5zvBdcWrGvl3Rb1RrvnylhGnRE20e0tqQBj2yJd6v+nDngLVFRpyV4+e97MRQ
Fu0Y6+wFpOmbz7oI8gD0FIf/zqlVsCNHGf7a3nJYwQ9d0NqjgJLBuZwXi/SdUw7F
++y9FG0IdDqW+DcbIUO4R1juorIoGyqo9VvDF25k1h/2WHBIEkfBUoFnsVGzM5xW
5gmlL92W2FH655+g8sM25CVG98CF6fOCYeqAoBQXy0UQaoO2Q2UVqKbeSZM9PlC7
UOFpN7EsqNtLWLGlS4a30yC36/o42ouHfOfrf1BK6bwl6DR6vv08DEjtrqMSGR2Z
LyyDqWlUXOP/rqhS1SH8pABJRXLWYcQlHVQFyi3y8c3EiRb/kzCqyIo8FdrNqhLB
5t3LLNNZapymHov9qsQJN569BJN/oeBodUzguO5mO1PJzZq5KQUCXQrVDjZoNJCt
Lem9hU9nmQXVvXAWPwM3H6RGNXM25DrHKax26+c2ZWvTzckgwUjYBCC+lxxCzKZ/
pqxszlyVhdTBLKsMxnN52exLm1M9XUpBI7cBOhyPlmlY562x0bZJrCnw/gs4OcwJ
uvKB+7DRd/sJt36//eA+npCuLN6utELMPRHEVmUEiPw8xlvhnhofw4uMDQc2YpC1
9XXWHTtTWCxTtntYEcFtELMbtfnsi9iLzt9Oe9qkgjp8SBCHgscQb5R2fYo3n07w
dlYKg6lnYIGrbCTlub4HW0Cma5Lm+JNizpm/pIILJSvtxi+UJTlw9eHcAmyg9UK8
`protect END_PROTECTED
