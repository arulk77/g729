`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN0u9FLD4hkSd3vlN6FHeTm7pVDLihT4hxMWIbKCg713q
ANKAcHXudD9Hj3FPek4Bh00+zXsGgeNjPMZujWZ6AmqdxdNsHRwIaDzDNJrO4hLE
caijKAs489jTq2MLUg/hj7zklWxZf9Y0Bc3EvEO7vcTDbYRF7Td18+KqwzVXZd0K
kuwjOvdyWTSVsCDsqpJHs/G4d6A0n0pZ7Qcoe2+nl65VTQf0IYuH5/OYGU2uK8fx
sH/y6TajwhK39WAJZQsdmcdBfoVRBBurgRYUOLYHWF+1rDNPg2xBowL0FwIL41ia
UTYl/WAlNu87u/LvJJYsgJivq+PbKhu4uKRI6IHURMUltiOu8uQhjV65NIi9Y5tL
UFMTCFb0tppqnRGEjyltqnMcqf8kYmiztmZvrwdrsAN8Alnx+ezvuntcAEfPsfew
JuUyxqYPqJw9udTVBi9qDC5AGB2prSj8Bqipp/GCI84gNqoTAwEbh6opdu4ACS+D
RKCxozG/AW/5JEOsNaYu1IC3kchQNV4W2fr46f733L2c27J92WOlHknfvSFFAuCW
9xRM9BwNvSMxT0KGtryajFgGSMPmRi60Dox53yvhymzQr4e7breaN9AS9xthz1qE
RKiHT+x7MwAr3qs9O7riJ2vsr7R+JOQnvCJUZX6iQV8o6usqktkiAdkXqMtVet8U
P+6wZvL5cAo+Q3dm0pXdcsoB0gqfwt4+VnAui4WlAPYOcxkaqGkz6bQpjRs7AHrz
Gz6gXjrHEFHdcozAZDtP/uLD/fTPFmbT2PbrdMZWZvRDRiiRnsCwUKrrqZr7c4NO
Ge+sH33WG1Ka5BJIhgVKJzs96nyFr7BCAnvpiJhVm5DsmSVfFqR3D7q9ktsgBigQ
JA0OkrKgmXogQdHQLiVoyf8RQfTm5HXEPMyDLAUh9eALZiFuhWtY71fJsLFtLvTf
VwgNoJU+0OuVd0zZ0eSoMku5LuGkppGDTZRoEcUmoGBhs0rlOT/s/6zGd/XbRqEP
D6Emvs+8SSS7haPEi1RKJnVYFF4CYkf0JykEFAhZWGrJuK19LI1m6jtAszPXfLDq
TCd/5f7SVLDu6wOTmTF2IhAyxy11I3RaOGgdXk6cx6h55H1jzg6ASav1GM5Bo1DB
wbXlyBkVNLg0yBz/1uCutQjX3u4wtKzuYLjgpElmkZhDVghCIVbLkcxBEinRZ0j9
4k5DfvKspkmvMWQ6AoVG7K5f6rB82KXKgKlyAtN8E/EDsIhCDCcbb5b3ScPxIts7
yYUeBGPvC8kFk4zdRf5SbIHbze/McrACFuDDw6502brtTPlIrrcPgFkVTrzkQMp6
ToPQNGHiitaZdoGlfro0sbtGcWNexrUYRKJE4g7cyEcMHqXQ8jAllVF/CL2lpz/2
tyKvXpc77kA+sqFd75vHQg==
`protect END_PROTECTED
