`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aV+aim5ZaTGlLZhb7FtJDw8OOLoK/x3v/MCHnwsXFCIM
0M2Ymewa6Thf+NupOW0WqcUIIQi/GxYyVQ60fL7AY7QIEYAsBePed78w8SmvZeeW
h6KBtAcRLg2QDXgYI0syR3aFtPq6VglhaCPIeCfzHHHwQ/oNSv8VKOL1g3qQVbgk
4J3JQSwNMn0DGtjGz2FBiUL1/Ut1RpTqNGEUtbP53RrV6edztLVBD+dyZvepi0a7
j+m5czDxpBPcDfwVl3fpNge/NiPoI1BZynMQjd+AdDqDNUW8StcL6SWuac92KkWB
CBCzM4vj5szUb1Jp/9ptUlIBl8fO8UbBEWcskoMoYvHoIXCSKL7hW1XvcGZbwuGK
+uvZ5VsAPmZeTFLu4Gs8pD1QoLy45eyJt+PRFX2dKOTWYqHiZRHItCpzrjiSI6gW
YmMkXC+WQNMKzgkSi4lwm1OHwXG/uzghnH9bIVn5sUtnAPhXLxFW1n/TUJBo8g0I
oYf5xe2XOdnxGb6q4UexOFt+txUmergpsn2aUP51qF5PiszamTtuGx2RHdP9H8SF
mRejG0wYh+9aaaPb4+4jZxl+2t/olwpBZI0UukSEh5g7V4RggdviwvQe9ennH0rU
8TufymkGQLqYvxudx5bzLzVgsF2V7uWSvhQyBTxl9yFD2ySKfuq44ZcLw9aIB+NX
Ev5xDI5+4O58Ju7x5ilSEekPBH0ksftPVUW4UI+Qf5I/yS/2ngkc+dbR2+D1f+19
68iYvbzwlEY+xrixtMy1K+Hsb5ml5+d04KPipM/48kZant6hjmxHE2YmH0x4/8iQ
I0uhtplDRkqm2o252NJ7SBVZXoXLd7iGnGD3/jX9oTJV9u7b/hlpBzyntpmqwtBv
+cDHNLiXB07eJMeFPaLYs21j45RbSI4Ow28zW7emv3kEy4ACyDNkPODD+lj+7VuC
DeRy/+5UgX81BUMtjJcZia/ksbYHHxoWUrWXKGSJQY/qu0NHenb32vq1rq1yniH3
AuYi0BeqVgQU5hAPq1Hz2a35+8DVIgbYnRkgpepdDwd/RRWNAMHbhcL5NDXEoAdt
SeTPE5yOm0b6gzE3Vl2/o35+9yy1WX6b6yfVsrGSPXolJ7rx5/X1OQDCNdhFVL8S
ZytE6MUYCtTzz4RGwO74BXNT0CjSfvQZpBH7LP4q2Ggcyju8emeRuzdMvANdWIVu
HCpxbGGkqCmoa50yKTCyLs79Bk99IYweDzYgQoS73+widMxCb9+dt07fkPwtEakp
neIUVQnCdvHuD/Vbd7LlVzS6AkRPgvvTyJkOVuXfZgsXeUdjEkBdPfuHrb824tgc
F1qdgXB27TrFBzHSsfRp/v5idhwy//UbJ11pMKsDIJbtCjfCyhLwzwVXP83ZRT61
u4G0+zcx6EqacXw3udkSeSGQv7i1XVxqinqwlsACM2OQl4g+3cp4gj0IAnI8OMJH
K+qXnAKHz6reJ04KgUxYQmlgc2vWW1IL71O7r5rkYMzr8Kt6FnMuPJaywqoBI723
COvX0d4AYTJ3U0j0LpEHE8DRfL6ObRg0HOaVWhGuAUi2ngLzHbpP984wbF4xeunX
MOCkP6VKTnF/DdSitlfgUZj1Nb9ovbvH2tJOlWPwWKSLT25/e7M/r6ZhBVMYZ4AM
vumDmVfOQIlX199ssxgpCyqC9BMoaqNKF7FO5qhd+So7VZDFYd96qdXhnoU0zKFS
6QCuKa4lOSUeLThs8mpY2zsE+zOyjW31+lEU21zpyT1sKiRmiT8LNBtJU1al2o/J
/dQdQ4b746axWoCrLT0nD8yHaCSBKvQLtO540asBBBaTlnQ8+b2QOrZS+gOT8bav
aRJxc4igq8OMZgnMEGv3G684qzdiO2SVusLQbd3rOVe9SpEg1/bgFH0sh3EOvRxG
D1PjsPNMguv0TESxvHwMXfBMy9mqOZgvDJFP6YGphq+mliWX2EIO3q7to5xlOZvu
hfmNjzVQZk5H9876dKaAIrfFx241u/lnWjamxe1YYfzpa3uI7YckBq3QxJXA7vQa
nOfLCvB3gLejcsHhmZe7Lr0ZJESP5TPs5A3g3FiOXQVz6JLpcPvjOn82+7zvpipT
xcskjIqBsWqBXGbs9r3A+AIVnIpTu4qXsNkuVbeImYvdTKDNLXHV17EiiWJU4qN0
1QxDC9CwdeiuLXKat90BCsdttM377Vx/NRgV0XnZ2osSTUzgfKWV1Q+oSUXgOJfm
WJe+qHP6nulDaqof81tj0/6Gq8kH6a2Wjww+4j1G3qWVj1OTZ15uJMX5gdJqkimm
Oxo4ORtuaVYt2r/VaLzgS5njPeaR5VBEky9qlO8Jn9METcKVzDKp9tfaU8GNlSJH
hc7LE2u0gKCqCW91AFAL+Lze1vbmyLNzRm+M1ehZR7UJtA1XvcgxkF1ySuX5/DqS
uit9VHrffj8axZ93Gzm7RnKNRuLz5KVf6FfrIIIuEP2u6XtmxPNv83hywXFTIdOv
2dY03HOG5P+0Htx4H3KKM6FX78xm1VL9NtswBdAT0AqPriYd8mXRfIuZp+be1rlN
WgyI7HzTwS1tmDwHZo/DYH6JMYE5Ve53XAkfW0JIEsSgGLmxIitcziPtXk1nscst
nqrbz3Fwu2pbTct4Hy2x1+yrkcB9WhqHW3BhNBBAYkprEKDVLMDYMHpf1ouA8kLn
SEqTCAeutk1kZy56JAaxm+03u5ZKJ9Kr+7rsQjWwh/R9lzfO6KadiT+diCuhVJF2
vR4Ym4kRAjpg8E/+lsGXGnSll5PSMpUpBZlNhkgq/XOOc/Uj4nrDtH4PCOxxGb7d
LfYj8f4Wff032xRuppCAu9dprud61a1jT6YQS8cn2RM4IIa69+TBered+ZegTaK5
jecQZUOXiL8Ba/THsQQYSnbeniYb6eHtB61vdjX1rRqXiFZzlZKKIXPaNFcVXN8e
KYK2SEKpEY6zMAOuWvHV2GyqS6A+MWYGqqNg3LFVcuf0H/ZlFnifhFcyCk1/rgx3
1IYvCNNV4aIhwXvnPoPbSKFIkIT43U499iEgbmZC7yIn/2RSGwc0hi0HYK5ZQYW0
5r7a1dLQJASDYHxXpUc4cQmBECb1U/uWIU/DQv7Wu13W/rbeFoqg1JTo9KV/jumO
FoTHnAMGP8HSnGPKOZFmvrjbORCORE2cyug91o+FYqt9SeEGD7bhXtYnXyaTcKdq
ZidLail+70+KogZK8D7G4tNftqVs4wDbXSIra+yiTtJoYz8mvL9ze8pSVYFgLhP6
bXNokGAzuZI88wYa/8LQ8zbWoJ1N3IG7+kDPVuFBUIDBrUhg7XEZKMJ2LkqTitUO
D2sk5PF1GkqmlcJFerCQRBLElr6JYToNVyXbZY2/F9GNKcfhK1/zo40qU2+nX57k
Uz2viHzFZlESkkoQLwJ3Px0e4CqIPXb5Yhcorz5hxSAFGkIPx02Sq6iYy4FUJCON
vrrFUFAteeYYklG8c/OsTkGWKa2SLx0xebzgPo3PAMrFU7o9Dpk706moD3OmAw/5
LWLZ/560ealEaeE+uObnEyAM+4bHRioKBcuKhe09+jfZ6OmNmrHdMFknJsuTkema
n0khUFIi/KFzMDF1ssLQLE6OHJOBfHX/namDmve5D8F8nNTaQMIdqmB1w2EdwqjK
43XyJwRKhYbhA5i73tQuPBZZx7V0PgI8sN5wuwuEpwteVrcwD3p3Sp+a60ada3tR
br0w0PvKoZKNz3nvAM80lHrMWFDciCFvURJAufpbkOcSrsUHeHrIqlTegAdVKzxo
/ih3EqGfpu3RPpdVTHg2ma34DGOo11i/ePwaEE91IhoqkWWaHLxBx3E3cGVJXCbt
e2Ps3D38+81y7mQUyMbBciI2e4RpIll1xrwD0blxYEmWjEHnm8xjcv49gpUduGpa
t1J6HERoSuu1+90C0duXH5r02WPMpUWWEKUJdpC+DbR68gEsImkRIn9TW83IZAtn
vxfJBLHlx/r6nEVlxrpODGfH9jFO82TAQV84GVQWqs62S9i585dWanxf/g0AcaEL
+EaFguw8FvfI8flR+A3NYuobzDLzKSSU5FpvvNtgpEvKsz9797p5v3sjFfKLmT5M
0Q5e9W7GCwFTM+pVkE8eGUg9uK6tnCeac5OMFYTwgdkHUNnO1Hie+FA4uMCD46Y0
L9fK0P5dBkqojYrC0n2NxX+KRs3ssWY4xJoCO77OUZGgMRl6p1NmW5C/ttHMuhwD
I0nlmLBKjc3qQuhjq3XJbZy0wBnZ+znI+HCeQbR42ArChUEt5kBygm8N6DW2tzm5
4cR0UJmbodVhIGF5cplVRk/F58vRIWAxOd59zcb+O6wAaRXJwljjeltc20+Q7krF
zrGADeIkr3uQ0Q965AG8HxTrvmklsZnC+DfWP1oDS4mwbhQ1yOePUzTfpCBItM44
mxiHlKI2MrqMxDlBKZTnP5b+5ahxHscuVMTIDha/EtLWc2JDljseh0T6xMGSmkxY
PhNPU731AXcuJSfvNAJ/0s7C942mvL+c3qpBxrevJ5cH9sGnDrlgd/YbPbyCugWw
U/N2PJN8M3ESXHHzw/DFWniuJIF5OMtad1YHbm4GFvdfko570AIxOYc0+dRha+U2
DDy2C05MBhT9H5+bJdEQ5TkacLLBeXFh1n3T3Cpab7ULUqhzwq55ff8VmTUt+JAO
ql+RV/tcxOezOiS5TC3bi+h1MpiI6TOX2lt3MbW/ELXO02ukj8FoQA47mAAHYqJd
FWwfF1YT6Oe4etT4iSMYY5ABReKcBg/kpzahEZB3gbax552lail8uqSy8ZB3mHQ0
ELfL6ztbKTim9Km6xOuofSMMdsDx9AhqklrXuvF8ZVxF0QuiUExL+48J03mlI//y
EjRnhy7Baz9itXI1MBbNwZ4MGbK5q/Q1kJ/PpgMBbTfBuVENPlrHFxfHWqLnvzNx
p90zv9P3WwBWYnBUY16khQXGSxGQYjFlbGyN/kxWv/FQIqzGDVG7xT4B6A7afal/
KRwGzntv5RsBEjnEfpPRfRxKuwj+ehKtcKqREeFQx2TZYrhtnineV7474S1QCvmM
UyGj+YgLCMyN7wAyaRy9ZJfWzHYwdSF81mMTDi9Z3YYJaIPIpRqtcCU8PQ1fIdmo
`protect END_PROTECTED
