`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNz7RRkSmu8dZFaeNM2Lo7uN+J5/jJPh3PUpIzsMpZKaf
c2D3BFKrRxzxTK8GTa2URNbv/iXL3lZk0fnf8fgy/2ht11b1Rwf6PdC93YyS1Ogx
ucHv+BpVftZRq8ihmbge2iWGHY79Uyjv9NqrIatE+kG6Tbu/zAK4zd0tI3COFDsM
1Gh5oy+0hbsVfkQua0tDwaqdKjRLYevJ2YVFbPb5Ei3Xg1sKS3jMyEb+00D0/wxl
jAn3XE8RNy1XGn93X6tsqY+qMvUlvhqss7yVzqTmZMjYkMxRoajKEbEpWKXi3I3m
YsDbXHYg5b2u/Quc6rQAIQhL3NErf9+glEXKojxYSiC1wuphr3et6YoOQmnfXOJF
w49fZKzv9mt0y8QGilUnos5PoILQPyiOITHTtuGwaXEAIKY6uLMx+ve1Op2Mtukw
fe4R8xQQHJREQG8bAcRFQsWTbRxxWbQRKYhz4HmELIcqofNP0zHeV1lxXLV4/ARt
Zzy2u8DFqdNV40d7KjYRGqgOkuq35JxZZMe7d0yato4XSrfJvuqN9JqidJq6dVja
TtZwV3h+xIXM6vyE14Yaq75Ebxy8W94uI7P+3v/q7m8wwYSzd7NjTVeDpwRaU7DD
q2q9JYTOX668CneXdQpzP1/D70RLh1auUhxKhXMdaheR86VJlZ0Mucj4lBRG9fGd
Z4YdiM2USf0VWFmFxSs+tTspgCEvMRoCxb0Xr40RnU39QX/I1LtU4Xak8sr3mim1
0Iqrv/6U/TWT3RxPfZjMixRAbJc9rm41Y+Ms5Evs6pflfyPo1Iujt3GN05la0KJA
7fW/YV8V8xnMXX5nH9lU+nBLSsFpMV7lq/mNntd1+/0xrLdx2sOY2e81Ed8BMFG3
AXRQ6wMEFfyktzbgtPqgvu9DyCxOdN/m+wjjN6/bv73JUTa1xQ/MT9bGPTFYihzb
aFWYqaa4i03e2U8ZNl4OQ4fZ9ZVU+nbUfgd24ciBeDrx7pz/KS1r6KpLD7EkUPjA
b8S6Zl2klUsQJL9bEXPHrEO9hCZe0vEnYmyWsNupRsfgu4nj55wAYBqrAl+36kFF
1xrE4mxPjzAt/NqN2DGj0e3QQizmFfk53jPZrafY7niPsjew88UCWas4CW8uGFSo
N1Ofy4o9j9G6INeEnMeTZgxKILQhP0pSvDf0qBc0C37VvEV/gPZ6uQZO9GlM6kKq
MtSAtNeISdTse3amWmlmuYSilz9UefSZ8OFTEXU+bxbdWgVFy9hnwjklCv7upGu/
bJ1j6hwvQLIdICWWoSmCNowkp+9p1MapHDpibNCHZGydpVeiNIqKezgFcxpxZPM2
epa2r0FuVWbr85jaGKConlovC3kz1dlx4V0WsPxSoS+ehYtQirVbLcnXXrD+4fMS
dfBPal8VKN1w/y8dfFAj8iRdkKylZ3K1ycQsWZHGLT5Whlmp5IkirfxO4MJjDdYZ
Bz96g4ACWzNY6PVjWAuWsRqWGboRm+njfK5HUibDDXtZ8Q9NrkHFAODoqgOo3S/S
OM2maUeRxXVH/JYZNJOvukdViUOPZvlda5vhUzPYk9PYmN19wQCkGuUnUAMLpnpA
P1Wi+1EZ0T/rPhfSkyHcu76LJsEX0DQYyh3CQSGjyr0OTWoeBl+/0clIBtwI0SwI
ydVW44XBnInMjoyihsdQufAG2ALsWH3ErhGwmjPX4+2pZI+5SGufV58WJspdqDK+
zV+0ciQvdJnqy6692vRqOPg4aH3R2rEM7zeF6tuVK/I49wNIEBsfnCHRRuvIpLKe
MFAh/ij2AJbvuV+BkqJN3Whh4XxI9BE8RLYu6xN8lwoDhNyYth7TAkuwYiLJJbkh
MEUDo5XeKBaPN+slnxAOBHbeTo4GyhAbVOgSDoAcVlLzA+sCPW6DS9zIEyIU/Zsz
Atp/G76lP8z/5hcGtRk8jc2k6TpwEz70nhYPdKKhK79I3XSZw3N7NCUluA2R20qH
Uz+OCb1BYz0PwDuwd0qNK6cvZiUza1PsC4i+4hjM/hRYPubeF1Zp1WaVEYYba7yh
jfinWaR1e2gjSrPsOOuAABSYak4XhdwPj9/5kc9MopY75tz0eu2R4b7c1A6gNYw4
m8Q2XVfIeFGyCpolLzwl2sAysT3+FPgwxpi3lxzAeRJMh4DybKlT8MSPiUV9cqqH
k+4GtehIOi3lgiRd+3dSijUHoUTScJNkhmVQdYGJU368ho0ky+Zs9bwQx+xkGi3M
PQT0M8HTBdX38gvJJNPwcIQVFkEuocFzCuY04ZHMdlMxlONXpc5SGvqxf/CAxSAj
KQkR2A4exY43Nkt51bBceHo4KeQVBd2YszLwvp6yHKygBt9CEdPxP4DtYmuVlTWR
OrzUK6ZrFpBPr3f0FwKsSEn4irO8kt8uiFpPKM0fMZacOclwFNQD7MfUHYC9gwwG
OI3N8iOBV4NyEV9bkma6JV1nYTXRfPGAj4Sr39bkFI8zKsGjqgvla1x5k7/ljVR4
GKu0UGd0rEuql47eWlWgcTLEtXbxIhLOOTRxk7bC1Pnadr0o3PEDakoP5dIu1kqs
NslgOhKo8RuU3W6XHanVb2zPR5gMQKP3nM+fxpX/kV+Zjq+PDGHT2lxEbqcR5SHF
DP5SDDID1diCaLD7LIqYJXw4Ldcki0CCCACokBDYNZ847SPehISlQ9GoezLWvPtA
zxgkq6Lr9Q1rQ0SX/EeSkVwHcTgNJlJtuOrSd2jN5tSOPGt16i5b6njKaFY5kOua
/MqktbYdF2POsXuLBFeQfZ9LTJia7dzskNQGIYbW3YozHT7zFpK/hixtx8mLfac6
/0XV4IVnK9o9KkF7jCdQtVA5DEJNmxDohzqcZawbQhOTFZm9Vu7N/hbPADcsYBFk
5kQyz+dBG1GRjYVIZSl+NhRYJzqmOZX15G3MvaadTgHoRdQ04qoHeEiIHDLmornD
st1bA13Ao0gG9JSnRlfsPCYUuysy60p0/TAJ6RjxgxqfS29S8kvR30zvb+5DeyVK
B6Ys6EW9pTLS/+1M+9mzvcGs0XO0/T6cwtiSNbGFbQD1+RgOcVwIPJ1c9MPBKPge
iZa0LE1yEHV3QB3/1tWJ/Xar+rIsXMtKjXbPEMpcRBK6wfWiss1OcmZeMMnp8FgA
cVLCEUPjQ84HkJwAr59wgB2dds3opXsKJDpZkAB+/golYWKvBANhwdewGHkDfrC6
F/YON8k9KinYH4v+N8R2o3UGx3q+RpZC8s7T0AcCyyk3euMQqJDW3gy+/EXsQtj1
AQoJUuY4QKeLWsXnxRhhvuJuT1MAUkD7+Yf4ZMTpZZcRubbhFSN7SI+1t30IllfV
3sb1Yaej62zxfdgW0SCXm2z/8r2N9QrnKEoRM7YEvNZbaOXpDUhQOv+0mZoKTH7r
AdrfjESmDINBjCy0oFYGBibqk2ho6QgD7dM29gK+NrTOk7E9e+yaOHNAUwNb1xDI
bStPNvUjxf69jeivJav6/rF9TBUoZsIcUxGtAJtGA0vwzeRkd8kvJ0DxTBeCanKZ
mAGDy8lngIfnFPkJ+33FeEsfomPPkd6a/0SFr1BMu61i/NKcQPwm8EUBtSp4Fdkk
/5USNERgqJTxR1fPGgtnn/bKa8R1wA1ryHq72L+s2DTdIZiWEkwab2oMdUjnafA0
2c2p6njft2DVfzWbHHURUMBVEm30m8FtZNFNKtveaHNRJ763u9ld26beE96wzUtG
KDuZR0jvw+f5i8gB7BYGMg95B+Q1ZF64Isi9JYzQROPKAsJ4jLVlEJk5uxVvOm9z
FIgZC23TMA1Njs3JORtKOVrED/Gm1+kHvyo0tYk37f57VGv2Rwu1b7br4iuN7Py6
D0XJj6nWYUIwVYg4o6WD5NpvyOcYGWNvH2aqsJeAhEY3KK4bbY8s5I2+SP4vIt/3
3uG5BnlmvFI9EkHeP9SQdWRX6GScBs9IZyxIQ/CozQXnb6VQ3Iba8l4ej0BgXrKb
ZvA4CBGJBZpasz/2WIdbHx37A+ADEpBH3QQKUVsEVgTl3xghFbAM30N9RK7xds3Z
fJMV0eh5eKRnF8eqmLI5FmWBb+ukcVpypM0mNrMieYRrcXOIDpXj14DM//oYFRVc
tzlhLCGtsBt1N0fkxvqH6STdSmo34XaOjgtZTbVvG8phNNerxM/RHT0WeTR8+SIx
VU1myw/VSzeDGfVHl/9mXKOZUbtiwSiClgJIuG1X4jZnyk01wLi2UtwruKxImLDc
1bjabXpxi/agPp2WnrxPkLKCwBDLFyEXDEZ3+PYNFQ+a5aV3SzPAQwFuxIBlyp6j
tbyaqCyXlTDG9CTq0XhrdYMiqW7VkyGvJwo+FStvS3RUg5jiQP1s+M3WI3VpWy6v
n89wVtdPc5XiIZ9bWZbpoY++X8GQodUCbugHC+D89VijXZota/4qRym8VQ9cGYFb
xnOTK9ZXj8ZkyjQ5i2Y+d/3ZmjoYbHFxI2ON/JtGX8s5UAwFEP2rppsPF4fqh2Va
kiRXPIBWT9l83tzUZNh88sgaq1SLrYQxoXPverfOoAG+qr8/LHQRjgaEGc56gpfs
EWvVjHxx/tNcD1w6wItePxFnHCzN7HaNr5e5qW8B7eQAnV3phJQoyUXyCmNrR4SL
ZRiAtcZYuFb5E39c4vrO1ZGuawFlJLgLnRvi62QOMXFx0QEoqqYVaBj38U0LHqi8
fVS1WwqbSG4r2cRjdgfMFmpnkwjDzsnYSNQD99FgS6Y5/YPvHInmpSkBglZ0qONx
z+y2M8aoNyyq8gP6L/SPx/iGt5Yx/wmc977ez6A0JZr2qwJVtPDi8HiUvpXZWPGm
Nj1TZI1udzEI6DEMfFZZmvIeiK8IDcaUJ952G9GXnbA6WDmt9tMWa+5WgJG4nR0k
OQ6lMsKrsW2gAxzQhBj3Cjb/SnAPFcV4UAG78FTseYk2BPpWQjUtBZAKpepzz7oM
ATDrKsHRJV0hxqn+05Rv0uvHl26/dWEutAjkzmhcY6PYsWEfa8/2JfWmU5X+r8wW
irdvPvW3RHqYDJlMuAyOK1G0mnpf/CELaX51nJ/Kn5UpDIoqlrOzQWUcsBXYT2qZ
XfCxHoajq8FY3AmlLg7hS4LYiCV8EIY+tYR0S8CIKXi/KzJ9zoHoo2ORdM2+gYl7
ILLUfR6c9Iw6hEEbNRqo94XCdK2GjbbhM/lvKw/C5BwblpQxKOVApo/keqk7DYqX
yblRRnBlMb0/JD9ZzYCCJEuhuYqQhg7d6MTRFIJxIUO0J/dkTc5grxt68i6SNn7E
JvC4bLFketEoR7N645v7FuSXJhRO5wEyyfScmv2sYkgwvB+SQUKZslfPQt26Qyk9
D1sZbyzXU6d6IlfsXwFG99SQ+i+l/nQwFhnnVPQ6FQpU5LUcfhmpJWM37gFHAKOQ
DtrU7S0aJGN2HLEc1gAi2AQF313RdPfPHEHgh+Zdh8uWygXir+gA/HsDRNdk0Qu7
X0OoFznEr5KRhLax8lrBryZbW0qHzNgKvTW2/pLDBy7HBkCSpZbVQ6yLo/SpukGu
g3vt8DcZnVh6wOeFzPAZjwEWSFoL6RUJAoR7nvjjygThi7f75pdoiv0JOfXDHlD0
XN7LksqRy/IfDFn0DZ4yFXDER6Cy4ePHhdM6VBnPVV8AJeYFXSg42wRUV834MlG3
76LYYB04OWYBNGQufC16Nlz2mW4+ydFMEfoS2SS3Qqrey0TGEmPIQKVPA9Dd4b0x
AZCbZsCKA2ZlZzCJIxNo1UeLRZse35CjNoCrQWBvEACcb1x6s/RxJtk1AbidJ/4Y
DO/7IOht+qfXz7ehF0b/ToXhOKh0JX+q2yqjQMA13eRQ0JPkFbrUUJCSYG43Sxcm
T0fd95imQ3w2Dodv7MLs4G82ocKajUG6MppcyiJIsCQdfxAoId2egsjJ+r9+tCJC
ezDGniGuCJc0fj6F4APlWdv7myPQdp4NdXg+RYl9zjHOrHUcgFaYuO9ZPPmA9NB5
PK+4UAkRI9OthCsbcvqslIjFqd5/Ce6UUcHEXGlTTxGNq2jWb8/EySPCcePZHQgI
98l9U4200T8ZwCa9o9wRmVaNT7zna609fRz4SrEwvA8hYirhjIyBY3uaedbgUsAD
w11sX7snXk6ROzgkuXYIFzazt99xkWxNQ6zitpO4cMVrmQnRKThfoLlYYqnTfPu+
EHmrdghbT2PJ6EkP+sfAYlGwJaq8do3quisizdsS6aksU8mwr9/YWurXL/BuHsKu
dDhaGFV+M8rnBLiAQv+P6ErjZOlIpY/tkWY4HcW78/tdJrNiVNWJL5RlW1PNiC3n
VambEz4xJbvWvF5SlzVY1+0tHMqCXHQ/+cmcHR0pZFe9co3UStXWz0rwgprNgd9G
XQdPTa+8gw4sBr07KpWLyDIbxEIiM7HT17M2opbkt53y5QpDx573Hdibv/WbKphC
np1DLZyke7fPUcQ07o4aviQ1lUvbNRV+AJF0Hjdf7UGDOV3KP5LmSQEPfKaqZ1vW
7l3rLSaKUMFMHHtF5dce1qvKWGIJrgmdidOVuHdUnRk5Wtn1TIV061qh8Hf6hP7C
15GpisWey4CW4HpCUJWC4Arw2yIeqLeEloWMw2zZJITKw/3bEgDkU3ipJNRjSUyz
3/qAGhglHxrlrKPeX1I+marW1OsuN3Yilil5PSY1IH/WtV9fegfcPvU6F0l28Owx
T3RowcGIyUqL8vvIicR/TfHp81yZUFoc9Jaj/A0Z/6r0Q0IMnvzLO9JsLbVTQ7PD
23BusKLe8P1ZzWNai20HwQ+3U1hvIPJ4HVoriH5mupQTsGNYcZbjCHsvSKNSGueS
x+Cx+vZl2cHKpHqL4/IA6TBJmQD4RgHkPEib9J2IB2t1Vry64rSJOThTp08YdjW8
aVt6LflM8qaYOvVfEqMPACJTIYRPcFq/zAlu9/l6Mct+iYtKvUOML7kvbCIiQjxT
nPi8l4DbgW9nMMeNxsG7nsyX6N/atSXpoovLnut1QzvsIqIiU3n9el5eNLs+Nmlh
qsaCK6JPhmA0vapu5PloQ721k1gQ+xUSkAkHx5+Fb9I+BLZ5vePdo8nmbeYxDW89
wQoL1vEaYGnK4ThwiUQv94J4nb4zDGoEnjO5B1mNFDn4k9wI8KuJPPgiwXqfqJj5
lnQBdFBky+6/xu0Ap+RQgDQs+AxdUNAorBJ/e0HUYnEpxhu+UsDpUDN5l7jTEB7Z
z+u7oap2K23kGXi9mxejqvCky/wlDqPfyokgkwIvQXiMv/Ote6GDtajYP1kje+3c
lygTHVKCeZWYLQbq+zoX+SLI9hJd8RQ9R1pb8n73pqzv+as97I+8tWOiBm0/JepA
e+4YKw/up3VECCpkLMrRSTOyUdLJ2GtOPw/Kq5nY8fyCJOCnhY5Ha3O0i88DHsk8
pDS8vDJNAf8qZADdVh0lmV4y4u+yVn0cxdSBBQgeeYx5rREuqyk5hOuV+wYUMSqN
COMyIDKxegYJCJpPAYISall3852VdVy12yd/QfEkKHYN5uljmWKUteaOtTWCL8n2
CopfZOUrP6hx2/VNoKzSSDRmzvaZx0AXd6+2A+U/hCjJ8sTnzPmbLWunkBR3/io5
4JnSQIEiGlbEHYoATODNbQi9WfyaKo3YVIabF1rBzNovTP7dlNOLkNz6sUz63iMt
P0k2cIvDFb9jquVpJlYHH1nTnpq+40IvqTuCgB6Qha6lxRpLXMkgJvoHxRHVkOYs
yzFRvqkpTKBwYGcPo9q3VESBshajD4+1NN5M81rjVTvpuAmgmvkKuoBh7RazSmwy
oszgvKzpAmzVOyPSRWxEfmTAMsph5UkAVJZS9j3yXDVx6EvCzTdcUp29n6ck5LYX
n2KIZLOfbxgvTVHVLzd5G+6espIwRdmP7N5wXoLIkhfXbynErgGoCBZol/5hz0Iu
bg9gSBWBk2DZjr6ZGIruzuHSoOY48m+JCgizzjA20K3oSSZMCLl8dBOtuHzvG/9d
x/Ach6lVUaNEVqAPgRB2OM1RAdH5mPZCe6ykm4hleGaYIMg5t4GssDT+0oTIj23q
rjud+rbINisbc46qJFrou6F40iQqPqr7sr7n7hgk556b3sjAI4bFRGkfgVSB9n/e
Z/8TA9/DWnyDtbFOiiEVfjjx4tY8ZFnUkNb+45zX8w9neJ/sHBHc0/Qlvj1bWuap
7Ym1rboC+TZPaNawfQXhW1Ub1ucz3mLpMgIBWVA0SsBm6W5QmmL8TSFUNAK4T5zp
3o6Mli9fBFLRIfACRvzVT1lbj2nNXXPO/j1rTQR62vxuYBSb02mxL1RYeOEGKIci
Iasy2fnhWF3OYl1Tm4/KxRc6vjqrd5glkRi/gcrn/pHlJF3blcLCPI0+kIgfZfgg
QV9eHBBvW6yEiemzZg8fvLybb1sBjjgc9OjbGAhWTFWjf1sc4Pw6gYOCRlQWNkvw
4UiSDuYBcZxuNIuq+ZRu8h/lKryydVFKjnalWTUa2yEQxtKVaiJZ0p8Jl8WeY40S
kDZgsh3n9SnjOrqRnhkswHLBsT/HyW+hS8gRWpigVq7KBzflqG5Pv02h6lo58ySl
KTiNMqMCxuJ+b83SKyGRLX0t0Uw3TqffgWtpw2EV3N8jhP4oH25kpeo9HlYtkyaw
BtvLEocaMX5X0eHEEL5NHpiB8THpFzqdYP4iViISBs1k8nnUMcWllPHUXfR2VwVB
vZ3Wb+phMkuL7fHsOuu6YcwNOfCpldINNccqoJ+mPRgB53JzXhnR9/X77T+si+xn
QCJit1V4fCGne4lG6mKvdzLQuUO2j42bqMsJHQHDakG2o43rFlJhTCidtjpRNVV8
bIus01ObDsJYBqiRop+ytw9m5Ft4EtX9bBHj4/pqX/ABs0ylyhcO9NiwhsQtEaEY
acx3R8kNWOLAGn4FGnbZ1bslRniLAlG+ldbijtwv4i6clHQPtWL0QbG6zE5/9b4t
Ieefo6kzuBvSnG+blgazU5Za1P4RWGIdPYchML6IVPi3cMaRpaLy96O6M055tF26
EzJQos7cyqJLuI702kVI5ZHitSOuiT7N7Yv3l7ro8FQ/B/ml9aT6h6UNg9GnAAYv
O/u4AE6B3EO9utNwwb/VuEaXZ0R5Let6fhJX+cZInxwsO+ngeyE9JF5UvdO9hJkh
1PbMV4NZRpR1E45yPelsuTkWiHXA6ja+4X4wj7NWNMtsVR1aK6uPmH2kfU2fFNlp
NUpn5iXrW6GiuHfu+TbuuvG5z0OeK0FLmzZqNjZJTf036b0AG1oqigNbPoQAxW5p
kzM8HCJ7VMLxQ5Cw79AgUvKwBCDRoc/w6k/jImtqfIfSb3y0gidR0gC5ZrdmTd5v
hq3mEbKHU0sggWTg+pnPr49ugLe+jSfA+8z5rUhKn1sxLRq/tCb5Z/NPpyAWTAOa
hJcMRuAV0gBuqHvfNLH9q1e5zD4AxrTXO9QuBUfSxXgAI9RX0MCDBbhKiw8jfJCi
Zvn92rTiuLMIr0/KZpKVXb9Rg7OAu4LwZD2VgeXgl2i3R6gm4FyyeaUZLELx3pLn
COSlLPUfcHfRsXZMQHIGuNYh4Kb1eNTLDay+ftjF9jU4HeLUBVQhl2K7cVKSS4W4
vbVeR2onDMqFiwACk6fqjX4bjofxUaXoLaPQ/h2yl4IjcwdD2PALjqT09IztL9Gu
bCfOlCB0xrwnwBh7NHwzBVvehQFuUFQ28F4gBNApeJYkg426ykiesg+3VEhrGcQo
rW4wyFvISyF+I/8VjNCmafyJNhkUxIKlwrgGRi/5ca8XwsRVgb9tNwwEAWBp+5nq
zfaZ21tH65pGKObpHibxSw==
`protect END_PROTECTED
