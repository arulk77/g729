`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJkhOo8cmvAxlqeqfzscdc0UbShf0nixXyz0lLU1TuT5
Mq439W7i2oQ4LOd0/xhkbGAn70CvvUjWzpNzdZXzTC0h3RjnhA3YkkMcyfl+XlWZ
iZsZyYPfRuZcAZqVRVH6ZyCduzSjEbAPklcQUyovKevm1mzqMWlR1GH9cYBWBy7B
b4kBk/H5pvlsjbh+mkJ2aW8MYlzOmKBnPhph9/tT731Yrx5F90m2bmVfTDgAUsGJ
Or0yLX9a8VyXF8ul3UhCGg==
`protect END_PROTECTED
