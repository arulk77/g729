`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLCk+67Mx1fradHQ9otM137VBnfiVyMJlSR3mLL17IJ+
CJ7+bzt4zmkrOCLjq+qxCrT/Gc1bCLKS4U8hbawLsT9Vi/UTgVXcKtpAHh7mojkK
pUJg4B2MN/isxjx9wTf2+Ln4DZ14uzHvDrcEoA/pfJPL2UcU5zv9mqXoX6KUZ/Os
2QjEYym2BF9MuELRBGFradxSlCqGkJzazLlsKhpRtyip4YPu29CZAaYD1NiWl2Jl
DrGWy3L4PkEJXCKNu1WyCaULMkYsisP7NsoViLUhkcsz3IXRNQdvaapjSO53kegi
RJLJnXi6+cZ0zC1GeAyiXYCyZL9DJdo9ranqNSeM/667QSQwbsTWFj5q1vD2RZOC
wrgjlwK9rXdw8++SGnwbElNSt3/hhPF+irMJn7Bre8jWhVi02MU5O8Akr45JSuLe
mUDcvB0ZjjlBpFbQtr9bHd/QME9lE7A6SmYAgo8Xy9g0GCJ5OxuByG2C9fJwO/0L
SrUM45Qq3DpLmm7FHnk0/kHPTCyNrgor3pqA3lxWNwPoEYNg+0jt9UtI4yn1+xW2
moZadoV99aMwyskcBXxwptQ/a3TOP3cnCSZp+upFIzw=
`protect END_PROTECTED
