`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45HlHc+4YEwpaQ/N7RnzkBZEu3dPLFna0TmBraCliv9x
8IZylc9APWiaXRGW8RdyjTZeE3nwXJ47tMlWCLLgngVOXl3PE40nUDtmD299uyxN
O0AgZdSgn1lZZDQTk2ue5H3bkFG0PHaL8slhOadVf21XF44pIXHqecDKsLxTjKbD
zO60NzJxkSk3y2ISAw8/fwy7rF7naFG5ayHrhKyFOTRgaZtwZSDgp/jCj9F6qQtQ
NCTny6KGqQY44QqhnuLWxp33voUKIVXYzkWhEfU4CJPohxe7cF3sHjk8V7mgqSis
QwI0ne1I6ZqwYwoH6xR4YtklSq6+S/VVoyVPDFO/keyAF/MqT0MnBRmovTBqQeER
qA+vgC6ou7+x/+3rT8vukA==
`protect END_PROTECTED
