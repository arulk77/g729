`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49V1JpIYJXI6CcfL9Nt9FWEOiBc2wtUI7W7N+OD/SRC1
6sNi14q4tTwDbFvHvMSF0wOocmBtq1x61wS2y9Af5J4kJM6M3JyMeifClp3P6+nl
WczRJAsBMla5vugYVR3/2xvCe6dIA//8lIqyDXYE3seqej2WE0As8GBjCvUIyAkO
9dcZ/Whjxo6bM59JMVde6MiQK9W0AF6Xq1xvbeWx000lvGhjYzgW9a1RYQRheyvI
qNwJdisqf9jUjooh0QeNAsxI6c4F1VcfJgn1TwQGfrmEB6rLmcjJgP+NaXBnK72m
YQXmAI7g03sFR3IBIGwFDBP6JZsw8W8XBz9l+z37ZuHUelkzE2N7byV8AYO5KM6F
HrnqEoMpjmVgzjFNghAh7SZo88h0wCJPj1iTRD2zrt30fM0eZnGJqmvd6D7L/lHx
6KSbrCigI/gFD1G3sNqd4upAjNn2FKhJDWdZ8xj+OEpReYlUDpTsk4m9pcXPYOoc
b+5S+TCE1ZcoRu96SdhucQ67TDgL1gP/TFFAP7ypJbL0oue/XfJWVbOnHlHn1yg0
xUDTkoVAXPKaXW6sJbCgwnl0zavwM96OMISMNr3L92KWxOXvkuZP/bgTboZaNJoG
5sRkkxrI/J+IK/qKn+2PKObkSxWekAeReC2J9xHkmA8ntnlU7hC8AMktGwyElBRQ
UKCUGHTSrDOGLVIbOaDVfvDq6lfqkgKUbMxZnm3n7yZozCAYr/MhQvUJD7NWXKQd
YlTJ/2UmS2G5ogiawJSOgOw5F8V/5iTCeLTMVdvl5WeALCgrnMut7ujQgRfRFtZK
nQ1hqobgxgb4m6JYzIIsk3nioT4cfL2YCMMjbCENb+htpyEO9vwcgSnTZGNqN7JZ
zC69HTHG0AX9lX3aYxM9Ork/P90hmh+VfsnLKA4Zh0z7yvI5YdsUR5jTU1DUEGUY
b0HsUp3JBME1noZfTrea31wgTOI29utuyFM4+UgLI8zsQp84sjqghjrEEQ6PmNdB
KxvSqoVKgpzYquAi8kaKtg==
`protect END_PROTECTED
