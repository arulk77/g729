`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFykaapq1eWH1a4MUBfQVVXl11V+1kcojPdskdyvDUVj
3Oa83OJ+qChEUQ/9YnPd/tJTGITotIAAfW5eh2rfhEG3zOURw/FoajxelW2L641b
kjnW8KkTyxU8wl86xJQbEGo+m8leZFOSgdQwtFnVPcWcY6iD6KrqXSnGGtiy6oYJ
WGdtnYB/dv+Oob4j9/RYuKfEaKX+EMdhCFFW5ksLN/Wm1cttc2clv7rLnbizRRO0
`protect END_PROTECTED
