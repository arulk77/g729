`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP/kPCTwejiMMs/BV1qfFsalDeOrJdXmAnHgCh4LbUId
7w+nh61L6ssOtDK73RiFToo1jvcoEuSYD4CeEzz9ZqZrQEHn21Oi792jig84DoWe
1jWTLkT0L38t/YUT1uE1ZUUMqMcc7YAOvA1QjbkEi121kCiRMAdmhba0C9YZhFIX
O8elz6Ud8OdUiyrNvL3zz8CdX+QYk0MvCnaXS6SnfnLLYZ/rRXayDR2OwEtgdeC+
`protect END_PROTECTED
