`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveH2pT+20Xt4TWcdtMp66dPOO2/au4U68+JkD53nv2HRA
4OSsqQjUnbmDfmWI0Ir8M0Sp4RElo05ZWbDv/6k+fGu+LPqa95Dyosj9DbWHZ0Dd
C8jst18g6o9r/J60gVAE+iDMTcLQF25aTBloiZ5mg8rjPk8cavOxO8f9t7comlSf
nFj4AHLKt6kBcoKx056IMw==
`protect END_PROTECTED
