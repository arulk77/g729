`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46Oty4oQ5kIDVn364EoncGQ1lZe7Hxwy5PIQ8KF1uyPV
WN6pV/kBwTrNEBAJCx6/H8zBB/G98vb+vPaSDt96frg4UNL/mQrcuCX5Qx+RQCQU
CNkFFhpOc6uLmXPS9FGSw/QzTUHtdsYqsSElVHoVD6V2fJOZR8v2vX5ALjTk/Zqw
lNiEkASs1evIeZwab4z7es+RylgI+HgO5nVgkH80UFk=
`protect END_PROTECTED
