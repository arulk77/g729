`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu432cMB7veHVUk2de9cS7Wt1OTrKsF9eyJY4Y7m7AYUsA
0dTcPW6tg2gxAxjonc8Df1e7gWNB6rQvXoGW72PlBbD2D/xBBPQEcg7xLV2GrPmg
lG69yqnaL9Hq+jOQW0Gxn0kstnWtjhDgnwQkn0LswyyhjuSRJnVQERW4aBBro/Dm
KwxD+WB98w0h1e9G21SARyMBZyc4/BhgpwRImz5AOc0=
`protect END_PROTECTED
