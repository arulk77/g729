`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zH/Xj67xlDoKYmwu33fQtsMSLXsY+UmJisCk56PZSQ5
H2c1dz8IeAYYOyJCLbWB+/w2rrJFK9eVWFhxbvO5frPMoDHNUljr+xNv2TTmYe3B
XthOmn28kqXfFMJl9b4kixx5mjN/yl36H2KLvdcYSNVsWAnD5fcvj0BtRkUw0nqj
pHxzcdOrWApjqkbgW0U7W8tGJd0SmuzNfIh3u9NDhwJfhj1IWATlFeUigPh6dchq
rt4t6t8kxQ2lk2Qf2cKCuCQ/p7tbgqIK9G8iLeI8sFmIpd3VAjt/0YMchykistRm
49rPyc8o9O02qrAmSpyrIWGmutpvFDOGN55AcfkvGYDlqcRH2uT/Peau8leqnWoC
rAKOu4HDxCfMdv3gE4N5vxn2nqjn7/IZQwjzUA4Aq/dzYjjz5z7CNfcHOOwHsLpN
SD+N49CWpslBYacYVk9ExuqVm4LrZ5IE3Ap7zi4fiqavIhfE1ip1YRMzlYeS8Hj2
44EF2Ev+NRMBzPCI9RLh+wcN3hEzP2N5Ysc8MI/hgGyRNwsWoBO5KlX7VErRJXGH
C5H9PUzerCrHH5ODBHBcaRU6jMzDEENWdKFczrfeJSqwQHgvJTivHDV2NGoAWsRa
luLjLbALjoh3FH9386e/wBtCNFdLyeJBwuY0BPQCDoh30GTHt0nOlq0jHZ8rLPVc
iGH3ztInnFv9QnLBGgWc9cIqWwWPYp/q82gwTDuv0kA4UpcpkREF5R5sHVZXmONF
xFmcWrbhs+66FZqopIKKRxbS5M5j4M3TCxqU5kaXw3enBmWD+y1q5b/g1h3anXj2
PEro7xhNxws+hDU8bkd8rWi0r9kavu4zwxK4na2WBYgVJcnIinebwWjoZJ7LLocQ
bWkXSw8laakU/zjNMsVTIUIxWX1+TTmplda2KUWHvRSSNgpJc9/XVldytWwzciqC
eWXYci6FpJb35D4MM9bDAO/6gNl1tZHWpK6EB+TnlLCgXMLiNWyHd2QV2Xnvm9Pz
NP4IIOY4CIs8Qo2bROgqtp0Pqje/sl7wzj5+aLOz6awzKqDVBLrfshkJTR3HTzau
RcJ2/ejZd7QzCetJiKzGS7zsM/D0I6P//99IhHLdthBQuer6RwvGjiuviLEcK67T
E95RzC/OEsi277wRo2V/uU1o5NX2X8DM81+mGBqhCbwI/DPNTlbbleeRg09uEhik
WiL/2+MpH2c45wha5rdfdEhZL0PhePXkAMmsGuG8XRVHE+Ws/XiRoNpbtlCOcL3S
6/TjWE4qLcz3ibRJW+PWuvoy+wlkdmFioJFTIYTgMS8D+qjo6gguSkadBvKziI0r
GdJBnULQ7qT4cGGcuE+qhXUV8lnooguM+sc+y4aQVOMW32NExY7hV0GuXncHVfIa
9+1xbvly8yjcK4mtPYr31r3FOutEsJovXMtci2N+jZvDRQtFVAJTqJHh4ynLHOjW
X+AS2pdWhu10Qx9JqRksIooROzDJOYPKwLtrkhu+yM5hPZU4WtdDyZH6X26VJgik
4hT8xM6MdNSw6FVdBYb7C8p06lF5TWX4a9SK6Q/wuqLZnXCjYmDb+Wq5+kSRBatK
O3366ZpF1EgNRjOMFPbuYLcpAjeUVTLA5bPiAoE5jmYfNV1OS4jsMh/0T8hkLQm0
bEDiGdQngE/rUkmkrelWgKnrbanCFxu7vWrBd/hFBrOvh5NIlbo4VeHYre3r5WOz
W7+SNTvtLduuSXoh9IaYEkPtUyNnXKAnOOVNYfqOTvAdEqu1YX1B6p1v5BGV8GdW
zeOT/8pcZTz4QQztaLTJkKrOVZfkk3BLlARyX086ynFGLtHnU74rm1/fmUFzY4Wg
lUnkYiXYzL8eyq3gMApU6dN6c3vTf1CRbI1HEgtAMglu/DdM3GQN8ddiUoBHOLcy
quPSpVeqbfWyXHTsHhL7VkOnAHyyB+Eaj5sHumeJeEg3x6mUHzLgYUgR52AtTomY
V7e7aOd/0alsXPPDfK7Pf4dXY5/LsCYTZbu+WT5wOlW/7SQHHcdAihLNhU1BMCds
AQTHhDUa1GA3gqROfk0JYaArmtYvcXRADfDXLoTbj0ne+79Qf2PRu7q4QdnUEjYs
z2DoXb9rgr/19DPnnCbdfELWb+eoPaFlD1AZ1Ed5pNwlSZWfv+q8Z+vIHkrzlicb
1C/uI0CwO7T0q9HC7t5ZVctiPl2oRzdcK5rJ0HQ00JVhFRFduUSLkYFZUJg4pBgf
qj0lcE3qENKa/4LpLN4fdJ2orU4lfwMCVSpLhiC+CWu+vJ5rh1n5vDAKxlwG2jrm
i+jti2jPNI5d5gYDAjat/Egn8vF9f3hvrno8oKiDolR9JwDlDVWAK3zHt8fF3+Gg
A19+5YBiMU9k2dWxMCWPtNj3+xbdZ70qcmTDVyjpX6WySNzoct0YSbhs/lUYMBen
FD5LvsDRr/rFnIzX+km2GgsMQUQayWBkqZmnpNrG6pqlntP1H+a1ghK+5mtmelPf
Qv2NhiKBrG8gpW0oavgYFyih36ZlIAqXeIbHj50IE1Tu9a0LsAMg0Myh/hUe6Wpi
eWq+Ck5X/EFuO+SVNCuoqvXkePZaKr2SZW4EB4pzFqnLBmp3Q2HSB7ShkQZfP8h2
hTqc1SNjj8CAyguisj37xMnYYLcFLrX1z08cSR6nu4OFIU3kKTWS6rBny6lso7d0
GviD4BYBSiWn4x71se9sCuLTuOu0UZatGZ5zXWhNNPAwrpzl+EfYaQpRmo+QTPr/
GgHu2Ci2DYm9r6PrIIJ/Y/Xo6MG2FvclbQT+tWDNqxPFAEjMqu0xWrL8H3dlTyjy
8qzFc2Z4eG7KO2KVwHll3OyvOaPOieGRM4G8iyi9ro//vpFAUZVh5xyssIP8SGwD
2Y4342bg95iQ+mU62R5ThBliiB/kxkiQuwzP9Cbm7H6WFSrnk2/ILL6UQLSSdD7E
E+DjYPhXAvfeCaUimUSSNYC83LVppvmmlM8k1XR52C7ffyi6trJP7ub9OAskeHTd
tBfBarwrRGlFDwWcLAZEgjbr3ViAVzm1ZZu/65wu1F5482f/NhBj8HvN/M/E/MGZ
Jz2yZJcgbeE5O2nKiLS3lgr5UaPmP2qQCSbDgTtPhlAjaN2KQLMALgaWb5jNagwC
MT4YHpqhplKcB4nRIvfcV9gEcbdHqNyTFxLoJyAAToHR//mxE0CewWLEFaGtDCG+
KPB8HQdtCIJnkVoj/Mr6Oy4a/G7ebtbIJvxCTtfpc4RgYz6DzwFLcvG8Qr6evj4T
QKPr6E6oZIl0vBQMWZjCPhkJ5ZWtjbg5BF6sx+vxJYHO1T9elRpZy532giwZ6bAm
dSjrkM3y+E+8VkAp0oSKF4BsqyQWRqfiyo++fTlYbxdZfu4a8h4yzp1cEn9Sf2+i
h8skV0f6/xNBymSXtnsIFC//w/F64hmVdtH9Tqs0i1Z1EZtvqtO3/exODq1kCRpa
lcR9j2V5A+4ixAwqh57YxmNMyJM2ox3j1u92GqKWOden9KyQQE/fXnLcuYiW+ago
exFH1fwE6o5WTbgw1EfVOj6NxB/lXMwPVc8rvD3r87e4/FUlhRlWvA8gZJStlE2P
HkGyaX/N0jbKsNVuvxbLq6KLK6kIwADJbRRJRVLnWB6YzRjV85cLgWHZwcVTewbf
pU/8A49i+M4Rz+cBgxrxSM6gfjvaDpnxC2nLcckBXVz4HMDPNGm2G9xzyv+INMj2
MKHUzRcCmW5di8KGIcOY2ywlNpqJvAo89RsW/4eYe0qCbr/9eypDZcdpt68ujh+1
joqSWOc5eR9vwdwZByxrrZWWFbJeFB4ViiApM4avB0U8nmnuyWQtPGI175aLTWYE
pZLxmOd/vBoG03XH6bJJq/NwEe4dTR/NiN1ioI3GS88yfzdbG9jcmP5GuOEAU0Qs
nzpdMs2OkIIvvJUMoFNjluTmYiBvwAzaWdf+2TtlZjawcaTIE+f/VA6YAc5oCT1i
eknGp5Gwep92lbuLoH9EoAowabC3G+/spilF1JQJIkVTatM55WgLrjY+OaoIEbya
PpfM3kvfIK1hDWF5nizhZ2CxeB/Naul7SFOSnY/xAPeDL17kg4ge4bies6uGUPek
PdS6z72GtDv2Z3+4O555rmQQ0p97WEsQRblPXX2TVMGkcvKyd8MP0l7lG2rrET9r
1BlkqpGTfIg6oWemE6+gyj8atF2R2uKqjLLSyR2FhP8j/fG/XEsDIDsPBf6Kl3Na
dGNRP0978wyA1D87fjciUDu6ol7y/dU9aUkUXYPfWgxXRTibFJlcIzytcZcg6HWI
gCVv3FL8G5LF2Hi/kJTnrPAguLBrDE8DJBOzt4LHGOV4ZnMgnxnUpSGzhdSAIPHF
ivzy7p1hcd6fIwsOpTAg3pjAm6bRbtt2kByNOriNwoqzGv5LTDW/C1Fb9EwmOEuL
40IX2G8BJ+VHpfZtqaXLL2UOLs++YjekTEjyHWafVFP+Jg7HEo9/Q2oU4IngcIEE
gh+OjShU0FADk0NWVj3tFZldOUKz95QOrrktCOo2j0atKGKoUbR6D2YBAwugZOOE
zh3eM4Pe5UtnSRXDhpOVewIHcdnt2ymVUqgw8caROe5FNj5Nx7Ez1YaO9NNS08+k
n0TMWourarggDpc6a6Cz1g==
`protect END_PROTECTED
