`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JK7nyQGyg26bn+7za2kuFdz0r2ibyB61VAv5oqIfBgC2Te9h2bP8YiSI7yMjmzAR
Ja+3gJHTBP8kGsX9DIPIjXcm4Cm5MWk69ov4I3TCmUmSOAsijlFAMGSkdquybhK2
z5TzGqrStsSJ4/XW7zCYPB6GJKD5ZI2iOm4rnOkH5r7qervmbJ9oPQR7/gPRTChg
ED7eCghOj+y6jd4bDnkCBkFSJLN303KVZrwp2Ce9/KSNXBXa5y0o8vHBH6OqsPK2
6NPjPCeyOaf3/lw//DwiaUI/HspbQarzuvnSOfmWXtXgoo4ma886Yqjo7ujOwinq
T6NscukRI6B+huQFdPQspwXU/lXVa0i86D/9r5l5VO4=
`protect END_PROTECTED
