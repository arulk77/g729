`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49MR8Cn3Aejgm0VA2sj22WzHr9HufVjVmQP4c4ribEtU
1ovXH0qr2fOnkRH7X/Yln+Wygmtb6Qq6cMyfBy0r/4+s9LV/t8AcCwBewa6PUnAI
4wLSZMsRQiV30dZUhyRmly6PiUwJejTjjLuOZOh6HyMVNWFUdWPR3419BgrFO/Ht
zrQaoYZ6l3JBSMCtMS+8nhFaab6rXuYaKh0jnV0Nu6Gzf2l2lOIWnZIEi+hIlzQT
67bLK+ZhgZyyoOudJZ2qgZW+ZRQbDNeZSIT7KDF3ftxReRqAGEv6SVR8+0wfoLDP
vVgcmCDbtZYHbTV7esD3DL5aDy4eorQpAZntudRgrPRLM6IpFzixWX+AkhAyElTK
VqMNb75YW5n+MnlfVsvFULXpX784c81Vjrmi23kLWjxa92rBmeukVH4qYV/+ocTl
UDdYFt02bzDAEjnI5gHTdRKm6IkTd2FMiFMQOk9UIKi3IrgVJEJdkikPXdzeT01e
`protect END_PROTECTED
