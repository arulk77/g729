`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49mQAW2JRNGcFRvYSXwJ+YqzTWHOjcUwwKlAc0F+Kyis
7YGp+Ifu71HkDe2qNnQQhg7H8a4XitaRTlAx0hYNSLVMo+N1PUQ6XaaloEkubhTh
Jh65J35O99vzAzV9O3htyi08cxXwLXUG7i0/SXPmneKYir9bb2UfKGZ/VFa+MoaV
PXH5ZRurxTmZQdTJuEmRFI1inoeW7UaxIscdkUi+Vgm4SwDmkGOE9//OxvE6DbFX
Y/HelcUeVL8zimuzpzFjD+/bwyicgX83MWy40R9VJGHb0vr2CeFmcVPJTh//oLK6
PqORHWeRKS3po7DdnJMjN6+wlTow4paXLa2PYhxhlocI2vUIT+BxiS44N+C7W7c1
FDNDdF7Wj1rNPH1Ll+Bcqg==
`protect END_PROTECTED
