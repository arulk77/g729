`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKe7bQxB3ghfqPMt/si2KgzoQyHfdWBlogK4kSiEZEZd
2i7IMJ62RJ8L3hIogxcBYgrjcoCYi9Oj7aFR8h28K9d0PxuVQuSiWVRR0y/OjG38
bBv1vsPv++bBXnwH9kqVN6tHFPfvZgZza8ZfEgtYhuZy/TjRsS9fJN/AFyA4mW5f
Qg8LSe02g1H6LGMw6lu0Vz7mAZsjL29cug4qzFkg5oNILjLHpG0WO6niiqTk16BU
BprJxETn925WSW3Ok9hGKQC8Z3Nx4t98wzLcEogLYF5XicUyZYeb7WLCpqJBSJpk
YTtTIekT2EfVENmMuW3nk9bAOYsGhXFtA7CbWXpg7z2nqKO6rNCWPbcYcubjNpO+
zsoeOFgCTGLM05hN/8XLW6Rh+zHjLdUF1JnNe11/KTV4VB4oWH6ipSGPhs4yfbJJ
vqB0h9VeB/WTLqyzSQZD4Zf37TbB5FnRksi39TkEvRFcTQdDP6sQK9r/59p6IVMk
sGghDnIL72R4dl9ZcKr1hdC3PZ4p9S0l7HLQ9uWBC1xPIGIXBEeIVo1/bfuBM8zM
WWcwmbaJr39N1qSXJs8jNF4798o71IIKIlVqUZB1ch9pMF3TZqJYkF5CgsKJ1SR0
`protect END_PROTECTED
