`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
vZok64D++n2D3c+82H/jdAnUgnchQJZp6wdDoHABZRAOUnA1rDXbdXLFzY2IzU3h
bDs4crHzEaZCIQI7WmY2BOKVZUEfA4fi/AD6dGLXSngqRFmGB8R0A+tHRbu7Xcu4
bcYYCbnJkAQ/+BMztbDHj2KcIE9lsGxNmlC2iwzAeqndXSh85zyl+uqdRg1XC2UK
uKNymV7tjJFxE0r2yZB33dNuSZCG0q1hPGBTbZ/CNT0BPU++yN5RAf0SKOfA2Jz/
A2g1jHKylRJQQSCbuGThzbc/MLABZoAlkoMatMWhfviNi2RqFV4iBobnQ63yV2V0
bFV9K7tbEAQJ2aS5/YA1QNA/5WJdzLx+qwy93wfTc5Q=
`protect END_PROTECTED
