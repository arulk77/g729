`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkaQ4bVrfzOGtVc/OCkfghQAMJ+h1j6Djl2OsM4FaMX7D
T660nr8VjNqNrhkMa5IRBzVr6onbgUmllmBaKXsaZkcNTkFN+jPPzbU1CXxdXwv3
tcXqyoiSBS0/WqD7db8pAMAI3fsGRnBs4Tj0wTPeY3mdoWgvLPBOaeLvWtP5dDxK
VXr6okBrfCti0Ow/xX6mT2LFPUWsT7D2C6HyCOeuCZ5OR9evgL/oHDm4njkY6srG
jcQiudYlvcNiTRCrCsI79EfMWNhaEQxjtOSxeepOwYF4q/lHyAiZCyLKOf/UkN0j
PPLrR32xFlQcCAapFnYc9Q0clsgq8RnaIGNgkXE0K9FMnKXRRy/hb34TTUxv+Pnb
F+PVy8+uEzLMou/U87zm6/y7p3YIEcZuKN+84ThMYsJwaFFEJ6OpKIug1u2EqWoZ
Y+PGU0D06FehacShA11sinTK3tbqS4kmHMwEt5qU5AeGyz67ZWrlKWRK8RBEksD9
sk0rvv+/wWasce5bq30cPQ2L0PE5LyMDsM7YvD56247Xc7WWwd5WXoIxCr1+/llh
xBkQl6ywYzzc2PRMxYxmjgleSmsylQXs689IrCC6BX8OQdf0qMZTXeKl6hkz1vCP
hq1/D318jQ2fNqzklfasAVM3nQZubV4uTIBXwZHH5jq+iiZIi03NN201Mt/dfgCP
J63G6r3949pVmPKVo4qQhMgrJnqnZloV/Jmf5Xega+RvVQjm+HM6R+tRRgjEXxFu
0x8KenvhwcqoD+GNr9S/VWK+GD6PB4y2mE9An0agcCGeQ6J8SXK31ZTF+hPNnCHl
mYsM/v4wFDN5AeFS2x69fSNPaofeYKR2hockDgaq4I4A8KQTWyRPdd7/XxY6ukTN
tX5X4ZurB9ufIK+JFCaznZFlnvUUFF6sy3H+Z4YNXS/XvqocyLIDC2p4CCOmKMo1
`protect END_PROTECTED
