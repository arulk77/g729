`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBZxF02/7owbGnMJ6ol+brKAWEJ/Z4R4PRG2RBvSceOw
564+3E2KBH61mPUOQX+fHaXY/k9c6Bgodxbmt2k5wmVPCEwcjkL4Krcut/2G1i68
lbZDlKjT4+tvk0QDiZs5zRES0BNgWlTzfvFXwncR2aRAGslH8LsRT9fVRAaIERtw
fhcXQ4JVL016CefM+buEMX8UKeDzsAXtq5x8sLd/x5K7uEhM9ilW4FGV+MaMfvCu
wxbj4GUhtfi2jUGTZFt/7BHsuVq9W0F2QLQqWKDOVLi3FvFFCDddYTg4NrrpN8G4
IJEKezcfxlvLLMxoFPEnxnZyVkkfHDFGrHvNJTe1lhC4m+eY84//RCl8ztDGNwIF
ePM8ps1eI9jXTaU+1AUVhDAv4k3bqX1qQF6I8bgCKZ7okYmJL3k44hJWkpnjij+v
TLJb/Z1s0/7aAmSeKqT/uoDk1F64Wo+H4yF0Y5dJOOJmQwcfDj/DT6d0IsLV1yqY
PY7I6urAM6UOG4eCpibPN2m7x2w0nNnvzeBvfA+4N3+NggVNzFuIZgi66zXp5jLR
ilBf75NYXh4p6xwzrpfu6yRNeNfyDL5hSMVhaCHUX+F6XUI9NGCZ8VQGYvEysDRK
jyShX8t96ldzDw4hVAUcxDGjU9ppj5Cv+o7KnVEKXWFRQYeoq7iQcL9Pr8LKWLoH
`protect END_PROTECTED
