`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2akHwXUoVotYVKDpWlW/3l9Bl2X6WZoWJCo2JQ9ivnl8ElA48urZqyVV7X5LT3k/
5+gqIYX6EvBmEIKLKvD4CPrQsXI9aq8pCWTuBaThFJpHx5qdXU+70C7U9jsZAGXX
TXZqW+6pGc6969CFRfl4JgdIrxuXFI88eQEiMZP9SSIaUa7BOW4PC6r+prR1xtmO
`protect END_PROTECTED
