`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
PgbIHy4OvA6S0GiQASMr1B6APzn4ikXU5Dxg7954MIViMX7lVCLWIv9VOl8nYXMW
+bcWpblEta8V93jbCYOYKS1QB2H4bHUZZhsKn/iHVHJEtaeHmHWWfDGXjAoCDeYV
QmWvnHjKRwt4Tp+UbZ4ndRhycKpdK3a5cKAf+gf5Yv6PHsJoWqGqca4w06aowJrP
u/Jh82UqwP1lusicAcZvjfJ5byHsdlagDTxQ6E3HV6JuXCg2ghBsLUZA4KRnDBff
RY1RTH1z/hJ9n0VfWTkojw0gUJn57H361Rr1ANfNsgrvQJ2GTH2bQxXIqFk9A2Ee
QECVqqQvD9YtHsHTVMS/tEGzJw6ENEqAKR1p2tMOQWyt1hScXNDpz54ge3CxVf20
pYuHvlLTbnvcmC6CEM6MQUl4wc741W4s0JvlFHUQ9943kLxTnS/QnbYH1F4BRd5/
iKzlwZFNlCclNAmRTFe8F6h82Hf0MsucwXTEd7bIf7jsLj9RYxs+vBRRoVLm5i+a
j/FqmXr7Iw3IR323DaYBoNhgMmq0prlQfC37hx5U1nlQuS/fvWAngQWZVRq52ssu
sHU3BHA8SmK/yjvOARv4woNpHwKZpQcSgUhzcYfdziN6AL/IxPakRviRNYXvNNIb
BQqVh+NyEJyqlYz8lxb+kQQZjVQT0cgXOC5Tokx7Mf0aOETbbOX2V5vnjHfN7XRW
x+nMk08qZPf/JwwIuhOrSKvxiKGjUCz1zR/FVdmTjJz1/BJjDDgrVmHZ/5s+j25u
sGbw9sGbQipR9DSwisPLv1tz3wi/NRHPR8n4SVHBuGc7hrXAGL0TOmXKilcolJt4
n0lO/u0s1xLf/vFNYBAvzNlEuu7QyifXzQ5j7L7aMAELp2pzM4JIWw0L0KYzhxWe
TkoVdhXypUNpLesVWx7CJid1F6T/V2zXqwpbbBU+4d8MrrdmPH4GfTulWudoKFfv
Vhsw6xjxk143MXKdN6rPXJLmF2PfnXFF0H347KWmpf9ERE4F3FVqFCw61CZ6jLj1
HHjFnMIrX6F5HK6f3aFIPkRpmfX7lG3YdiGUhUVvyp7ki96LNJWS9MAduv3yy/9J
c2MP7ezbPLybDNp5jys0sbayVVSwtbIsk96K8r/xi5luHWljaDl5NC43PjJxzbBI
NRFtb+9qaoFGvPC6U0q6OdAy3Kr+Tym2xODESGz1MXAh4KfqynADPF04jX9SpC4h
1lRree6xKZ9DDmzSOzkK49lLHeyuJ96tY7MhfwxCMvvszd2idAfx9cltfat1IO0x
5vbxQP4tuJUJBR71VgmFiXnurt6bzCfZP3lNDRq7KMKL5WAmP4NvbiSr7FEXlGdS
+IP4mS91b8R0HFoat4Jj6tjCJUQL/HNSVTR2AunA09CNnhNhelD5ZGRLl9B35sa7
j2lv7YiEn2XvcMSWxPhywcHkcHsf4Fa78OHIeQ3uxZilHoxpqb2Nel3RFFEEsdZK
nH45qFkJmAMdiVYb6DUvoHo08xKqvT6YY5iMmhr12avdw4DP6ZehEzMs3uLdzDJ1
qka2eZZxa2iwHiiiRwY1g77kS+kdvfnojbjvrTxiTxgVQxWriw5EE2GYI4JHhN0F
dbvAeNeImI8sBmtgLMzeokU/VZYtd1QjJnwYT2d4KrICjj90DkETgAJ8M4QPLYCc
RDOsrcRKcZnPI4sqS+FgapP1dYf+uiZbhH5Q1mVjRfEl5iJOUk63RBnUfHsatA+p
xrguYLT31I2R4BI+gqzCsqdQyYIImVqh3Ag781QeWEy4PZ0rgu0DiI4hOJS6Awuj
gbvQNXWSNLYxCysSYhi3YbtEBgakpnWmcXV2X5iBZm5N9rIY8OBWLhcw0TIm+SHD
1nydOA00RfrOhjnukb3C33kgLC2HICzN1roe2B/LrngHH8oAlKe8+vHwWm/ofszp
DWSaTklNL68Lvh15qO/hab8Akgq19iEdD4cznaW8V5kQNeN8lHzjgfNWn8nNJK5Z
Oh1+QN4VIYvmw5D29+xSmokHbii+tSkoNTpu0R4VmVqVdyPX1IXcmyztY7iaHqXk
IBL6JR+BjNVQH6g9Z70TmOxyU4HJ77cRIcu+1tRMzHVKbEnGOiYuukQYqsmICxL4
CU3qnMkN2+4BFGsbvUecx95CHwz8NkJGSpvxVNLRdJN8sVM/VQh/CvYYx5mGiNgA
sKIxrjAM80CN4TFzVxpPwF4ZUVauLku9ufL/hQ9Oeui1jR1nejCXPBryZFprTwGc
Ffmr2zGN8sE0PhmpIQ2Lc2dYiGwa55vbdZt+fwMkWSRkCs5WC2h/vFgGrQtDKOg6
iVTmFaoY//Un4q2N+zV1QPzUJvpxxiazghXXJteDlld+u8UFde6XF+jUf/CC8L1F
8fOTVLqChAMrEy4tw8gVkLEUGjq/ECilSaqRsAoxkB4zAPdOt/9/UkURX8nsFzix
A58AMuvBlA/oX0qLlfmqZuZaOmr42NosdtkekHSjhCrADmZebIlj6yYBpbDfyrjE
2i8ygrBR7q0bmRSpa2PG0czi4ryKbsexecPjS+X4qOmr810NKvUqP7vK6sutkFcc
1NtT3HUOQEq2LCEVQN7rBVJDcOaFe1MwpzFJtcYgWUR2K96KPsOSJ5F//eMQakev
9LpA+JMncrah4QSDtnaRGtWIiafBvpmoiGpCizRMdS1DOCYqQVcJkYOz+yOr+bu/
s/UkR6GNixxoJY/zAwYX1WBkBcXacY9Cd8XzKSJIpkoF+KdeooAJCVynH+AKFfAZ
5UXLY9Rrkc7zikygII2nXZA+d1Nn0sy9H1ShtG8ZS7j8U/TtXvBiwDnhKMfhOjDR
bHOrvEdsvfK04WsIewdOxeeKXIPiMUJ70xj13tN+GqdIKWZdJpFslY4Em8IusHjT
hMGKazP/JBAFbMnNhxiBqMUhzsrYYUUcGkHjYiwC4taDyxWuEpQLLV/ErsbNkrbB
rpYFtauqeInx/IFE3uEfT68s8hbi7Ea1RpZt8pjKzPGPaeq+C6Pr4cu1eccyCFt3
CIWI8pzbPVUpRj+DxIbx9GUvgSftYF/dHvXk2DTdoYppKEvIhgIQnlLzL1kImN9v
Oe4xVQBvlc7VS0+47x2BsQ1NIN9K7ByN2o1dY6YOdW5sXRA1kOSplVHLWsPOJR0D
z/l7gh9dIB6uTeqwDpK85rbyCcTTnKBfDaPUrGAUCA2lO4kIQGSI8yJlf3qz/Fos
CVAbug26WtNrZvbQa/uaXaidTiR4HSGRnvBRcEkHeUOF6MT5gI1kjYpYumLdO4fC
1srzBjuGsP3NGl1pPXYyCR9vaQW7WGHWGEjamuYdtFyqYWKNRGfieyY5Hz0Y/W7O
DjKWa00b4EgC0hJIcmeMtIZnh3UkbEf58+H0elnEI5IQepqkk8L9mtzn+62PsLBf
ZOyfmXJmjQ1tOZsOGfBgckA03fv2zTZe5jSIbxaCILFKKKQmAtv5CL4QJQLbE/ob
3gkP5WWaUXJEkhwaozikVDYoQ3C9FyfnG2mVvYKepDefKW/S0VPTqGxIraDnh8GD
ivLrJrdPtD/myk+A3s7HYd9XV1N9o1sE2ogp4eCcv0eXnNxgpzGtbtuApC4j15Ku
kHpw7oVDjQBEXVEgFlz+tA1dGOX2XaFbWUmFpnMdHD20I70YvDsL4Kg+xoC5QQ2z
DBB9VJkGd9PccOOYBd7Hq0r1/AwOD4zajibPAkTJhpT+9mbALMPHgGgWJP+DaRmm
wFtZnTNNhSWCqXGX9Cx+dyHrkqU9Lpmi5UpJKmPImbX913vY6Mwbp8yEEA4INVf9
N5ePQrU8O4oxo3uwXEu+gfReydcRQ+BFEAN10aV2vpo9xfH68VkQWGyd499CycLV
MTA6IuRtsgl69mU6p2kG5irk3kjjJ/XH7MvYIGM/X+3Z7PjlPB2tIIuPzJaufal0
MTqEqHbveBZ/aj83Bttol+eFZUq1wPA7XoTyTxJNBXwHtqxu4Nn0qgYEkTco6UX9
s6482r/dGh1h++yEKCqQsZqCBtEgvXigWZObPwgl5Z9k328ibG/t4jjW8/J2xzBF
UCKjV3sbqnb4Syyyn4XMjKkDm/A/h27WKYWBKkmceLRx8jwAjm3sqQFnj/jc7s4S
iXwD4uDBr0e1yu+nB3N8Rtyvui8wvsOednPxRfQ0kk79DEq+rZlLSbuG3UkiP2xc
Pa1Drt2wwHWDHK6lQh+ohfiV73I9Hbf7FnRKMXmxyvFxlMDeypVwyUGvkK5+SP2v
Su9lY3gE7ClzFuunZyBIZJ7RN7DofSVF6iA04pikVTfam+hS7+IcwBniEUsT8f62
4RGIL2wE7uvfRywIQv0tyBvJqIATCGfSrkmJ/N0Ye5LFoEwRQHqK/B88cg4WxG4e
enzYBMkjaAC2ET0VKCXSRCWRfGQgvpraFARfyQOSVD5kgM2dIpDWebvUvZmSREeG
KaGNi4kcRPHbwLbL/bKcUDQ0j8Tk1SRs+U/WKHkM5CGHbwik2B2T+FMN9wjOF2GV
PQKuKqlsJo+bPEOAXUwq256n37c4QVyMDCZw+uaIg9T+5dnT61Wr9vvKlOUbCj7/
MI0bsY2U/Kx6fdU+kPCLDNDYKJc6X+b863h3YD2hPXtDJmD4eSHrYKRFHVzdz2j7
PjSIhKVQBmsJ/li3xBvzyGW6ffKgl3OwLUZZDRNmrIEFvpzx1G/fXWB1RmqMJtSh
7D3gKVUQUqBa6XvBDIszoM8xh/Wi5Be3DWljNeFrzr/XXqKQyjc3W8fHhjf2jTyn
hxXBFZFy8CiUAViBBzvzI57DOUql9XJtIWvtw/8sz99ojItiOY1cSR4nyOHsaF7H
8BX2AN3yH34Aln+ztUDdQK8UMHow8S5yucdwU9u8qlU7zUHA+7VBF8Db3hXyY+Ri
4iBfp5ArG/3SpLjoaYK1ht+tkG4/Dq9zNSn+VoKZb7r4s/SnfqGusbFk1CuOCKjF
0X6bAgIs2QIg433yI3jRMUbXipLP+qvgtzmw/8rE2eVqB67e4Y/BTgJK61yXwPSX
ZuEileEsanusUBTCtu2q9W1zIFbtlI1UV+/dCLJDJ3mxU8w0os5rW7ww1mpP3NlQ
FocjGa2+GxwYXJUvsUGRByrX0qO12hCvHMbHEa0V0ow6MnxNYA7ikPs0NG2FiMfj
4iuTBCOX0auNrfNzrg25/qE2Bd1MPaO33dOeHuxAxSxiE13jV3Y3bPtKf5VYDg3G
4nWnMONDL2Oi9SjgpFsjv5Y9SWbY0YbY41qB68z4MKgMLdRw8GfendqRd7yy2ScA
7kJir7TEiygqOvLYU+am7DzxAsEOoEpMZaiLMacRYfZJ1Vlfnma3JyCchEPyQ8uu
rxOcQCzRJBKVUcFfLh78TfjmKnIGTrYwhHTw2ClrwUtcfK1Jlkhl5BuisJAhK518
GWv0al1s4UYpCypHrldWO6OvjGPFXfO/5y9LJOl9M3FIPs8zqQj0UiryNF3++GU/
Cu208jrw5t7meLaYGmY7jqHVWkfhCezWSQnXq36UEKpPLzSqAoJGXz/z/BKfYoxs
o/rwFcPnD2Ewo+bwFV3vHQ==
`protect END_PROTECTED
