`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK4QnhrV+uMgagkMJXlgCIf4JLYPtBQOxfy+tNbDG0+P
Rytj8kiZTd780iprZaVMKPxGtwOZXW3Wbf1FLcK7UPnzUkVLPytXtjTiDWd6mlCu
nN7diO3qZGMGWwu1r6M0H7PHz8hPyAIEatT2FGBKWPkr1yuMV+CewFB2sX0tDCea
iHrk8ZoTRpLCUIvf0CVKffqaZw4HFkkLMqD+suK+bvlh9JWe1kWfV6hdCyhrkmbG
KBNv4O/obYdcbBwA5RB2WOuN34F2xKRmaR7PYaOvGVqzeV69lqMEDIpuS9JzR9iH
QBl9j5Sir/Z5Q5y1d/0hpC5OPQqWGrVhlXlnwK/DSA1+o4RayQ8KSE6hi9VvNb7R
ty5nYUu3QwQ7lvFPSh0sRZTb93rgfk+mIr/09MAeULHhqIL71hg8SQkp6FvtziB/
8OyzLdbMAnCz0GRZX+pZXkCXPxqu/lgrZR/O5j/bsvZedEJls6pqxN9pnpZnT+aQ
NSGUChbhQBy259oWsYK3PETAHPrxSej2pP/Sd8A+B9QV5DP1Sr1nNX5gKP2nf7Js
kc2TRnQ1vicgPzTK4hu/6JVn5RMKVqci/SRkOHVAnWSoDUw0rVO5uq8dwZsq7rCc
`protect END_PROTECTED
