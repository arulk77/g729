`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49ED44rGCfSk12DaML7Wf9P6ypRqoWNB2NL/VUoyLnjx
hzkj/82pqWBy6ro8TJ5IAm4y1WP2GD6gHsUwwBIp93/PdVyABu9EpjyvBL4vC75B
je91PjJJDbgzWV7GNYKt7b9I40o+sKUyrJoYKmMgD6AaAMBtVfXqGQdgPJFYUR/y
EA2LGog0vYWWuRxkEXG9mIl1R9tcosodJpcBSsOK5kQ=
`protect END_PROTECTED
