`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
0AgV1H6vClQd1AVUBGcij8K/c2zaW3gL1DwOlaCF3u5R1JyQ8Bmor0DUpj7WEEqI
3xNBH6aKeWXlCIHvVQdUAwST2BO1SdtBNnKn9F5XWSJhm7xnSUZ0JX1cdOfajmeL
S7UqjkrpujBPGs1/y92PDX7OoEtyvvrP95hMxg/dsuj+4dKD2bDDw4nCSrBbKbhr
iUFJlj1MLdgvOmHwn/HTjOTWrFry4I825jqgV06Pdfmy+6+8pr/7ufbkByNlsWC9
cHqiJ7nx6K+FvMNXLSwTy18/qQpG1m42d8K4SQZXuAaWXFm1Dmyjm+bQ+jNl7h9b
C4hCYWjaGuUZwv51QVQL6ev5MQmN2f9hEz93f9LiQB5UadkwwiRyDoq4bx5iNVvN
6vFgzDLNbB0rQEuof75twGlAtBcK961rGsDjiA0aXEKu9J53MLvr9D0KJupBXutB
/i+HC6VsmReP6ZlWCprM2gMEEPJrwCncHIQ1x2st47Q=
`protect END_PROTECTED
