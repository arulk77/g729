`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3Zs34nxuOHqbFxU+ZMiusHamfgnNOx2GpKR2dU5sQzBTQVbeu0Uvzox3ttF5Qsco
rkRUIqMUYmb7LWaFrW1EueuOEdP1qKYfa7HGC+8dJr8/vaayIR+oU6Fi/DdvXqSl
Xq4+48+q+0l8JOMgT2egGjFeD8M4A1V3eG0B4ZsExe0gOY0v2TCzcTSJ1l4OR6Aj
eeqdYIZiGxJDsDjN6aQWthn0AvsAZcm+94OAZOkZcnlIKLWUCCRafkg2G97FYNbk
Cce/mYdoQJ8ayN2evHYT1rcenrjdoGayVb9II5+YyCr+kw2maYmCaiBmZBaTkiqg
OEyu4i+vOoME0Hg8KgI9hoqekyvJqdw6DUyVVySlzBcBMJXdZucjnn658R35MRIl
p+hBEikCdLxYyi2L/2zIeg==
`protect END_PROTECTED
