`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN5MNPZ+RxcSQZoLem7ZKftvAYyo8vMp2ehp+JNf/o6q0
uFOiFLhLqH+d5RHXBTgLAO/Cmof8MLDqQ9l3/VOZASC/2atlFl7v7T0SHTzDCJ00
hmvVE+WbjBS1npjgVRSQM2wLub5U42WNlU8PnuFuckF2WGkvAXKb6AjdBQtZkzv4
3/xDMgg1kJXKV1oIXut2+PteWhN4IlvXhCCNva8/1YPZ96zzPfWY8+zGRTbakoZE
WukNoV29A+7IkoInMuC8a8Fq7qZN6Gpdy6pBO1IyVjaur6dYAtwK0EXpL9Pzk0G4
EOwvNDxT9N4YaJNOCQ5OT+UBGGsuQP/EQIOZFdpoVmENkJ1GcXqvlzKvzFkwFvED
qgQ0atUjJbFa4mPhy1Fyv66K84anldCGW6T8VDKT8PMc8AOrFRvIuVXvmKRZshNB
V+cmG/mmIrOVaIGCCMrVjFssERFrma/3CsyupkskERna0KLRcsS3W7e2clYUnGJK
cSx1S8y5Ss+8ekUQy2vF5hgKHhIOkA9CgI7B8ear0222ymJchUdrOVN/UfrzrFMk
/vy/FAjIBG4Ozn7Q/gNJE9tEhSnS+mM2gFus2xUUgjg9u5JLFHE93JjBATzo2mto
fjOcx3Lm79NklBFrOnsk1KBjBVe60iUyJedVc1YZBTSoKS34FufzTvVkuAXlxbZp
zbFulrM2U2sy3c/YI5TiRvQhbD0G0frk+j8mknMc912Ijwr6MBIy+uUwYFYPRAZo
HO9lC+8P3E7UK/XQIWq+ZFQ+4dupFQpPoVOwF8eWwf29OYLp9O3XRK9Mm1vCxdqU
v7UTqHMFT8V9eYs0gxsJGEW0sSRVOrMqdH/Hui0CO6XF73ypyt2cHsHCkJxINels
AceHIFzXCPocTNQMaTBsEVXhhdB7h3LJE6qPy8gyB8J5gDa3roA/kv8W5U7fyaOl
DYatGT48/pE/q1km6WiYN4E/5aLa6qEcr8rbKlQrpAyio/MfP/A/ykVcs/qfMGPL
cuTMr4Po6/mvNdr8k10YcDsqRXEBsQ2Qi4VqrkpAox+hLrlIbP6TCkzaNkbz132l
uIGvlEiSyM8f2u+8GfYySWigVnyTJ8mfvTx/Tfe6H8inOrwLvrjpyD7NjGRldoZR
jvmfktogvxlwe99O2LiNfabAxZZ/Ya6wljci2sCOtqOgo8lzAU2Q/beegTza6Wbg
LyBIgSZkCcpIXzKSc8+5VQ==
`protect END_PROTECTED
