`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAVcutHD/j/Z3AEGK+XlhuSD9l2PyyLgY4A6tYVIbnyd
qXUJV02SICHrWPPWk8qof/USf2JMjcafhe7KwfM62DbCtiy4OSW6mVgeFBdmRvVu
2p1SuzKyPAfJao+lHnMkg9sGggxB/gNHN+O2MehUYxrXy58JCYn0BDfzvA+givoi
UYb8V4SRc+AUc1DC1LCbEPWOSjswdkWyMDnQOQkESmRqddSKbiyZO/68SAoBccyo
`protect END_PROTECTED
