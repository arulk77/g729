`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkci0QINRCK5ph4cVK5wEO0MschzEOA3Lsltwcx2U8U8A
0X8qeJHKHwAkOFC9e5rPwf8y3aEkM+6xOp1XshP/FvIv+uWqHV1XjkL1oP1dH5YW
K4oa3YexCGuCUDxS918J+z0qmqLhyREka68hvKptzRqmIC60ELcoLSqEYrpv4Hyf
ocntNSDYX4nUq0jaGHmdQW88x33Cek8RdtTvK1JluwigirYBPjbXLc78q4zU4yON
J8UZYat3BEJc9ztKzpNQTJTojPyoHGUvwHZ0LeyGmndwpDTQL6YE8Fa/IWkkXnrX
iO/BfpXqmeCW4nm0pbcYEuRiL/bu4BnH51Gj8Yn7g0lO/2A75byr0qM8+reEuvkS
VksxTVQb8kXmF2uBw64Fmann2Nb9WBH3gs/AbLuFTP/sm2VF4mKrubWnvI4CyFW8
7feLl2cBMj5SPlg9nmAVhpeIVasEap1yoWe6w9o4ATlPfB9zzaJDty744zxNIxlX
/yDwRUoTni6mgt14g+lqpUmhaPC7GZ/+SkgLYExgETQ7//UMSk5Uwj9EOZkKDr02
utYsAGruojL0Im8e7z+DIYjeqIK0X0LRd/1QmwkNMVtZZdBL6VTR1RLsE73U/wv1
+3ohC52ZspJjYGlrpRkGQHWsB7PNeZnRh0RbxEngrkCSDIPXMBcGOSvHoIoOnNfm
1wvRTMnZ1i1VZGq/Y0pjPyC1/AJ8dNQ8ZW5yddzVJQ3fIU8/3cZ/76iq18dD50Lh
erezO2uWjyfsgSgqFqsjpbZyeDP0gtrLDuatyR5C+PPJM3PQ348MoARKnycVBR+e
3quYFBO+2ky/m8i3RgebcL0TGrzi8eutxezlPCDTWu0A0pEycFpyGxIXwXUkSHNy
KTjSQ2fSrclq2AyJy02vPK/hvTRLvkyY0qtkGC9W8d5no0QJc1ih4aVOesgNOnT3
6pXBeOT3aOj9u1RdIjWIqJ0Qj06W08/XbKr+NCOMhKsLsEPdzx1lekTW/n71JyCc
glEFVS6Tnbv8saijI5q4QOrlPElv9RzCo2Ftzork0VwKM/r9dxXacjuFBSbuON4U
V7nH/DyCu7Gv7p9bbDmAu+s45laul/m+AwJCYJGjC7X0oM0CPq8G+19QrZM8c1Jc
3cSRBLVUrr4qnm+H229fD1WSXTerHAQQUOzDv+I25zpUVjrDO9/L0MoJJzXUm+PM
I2IViEH48mnKslXPsqibvxPzNtFt5V93GLF9XamZi2Ovs8EX2YOizfHePLgxlHjy
wsLGKVdS243HqixJhLsnXyEuNJa+MY14nw/X30NrJsUH/Udb49ZSTP0m9Ylj648t
51ClSrWnkvLJV3+ZUy/MuocUCjn8KuJldCdN9uAe/Sd+iG2t1AGr2NaADNvGVF/3
8+xI1+D8xx9F/gebAw3318JWRGUWBduL7E/7cz47OJfxs1dycqXJkrK9QHjbQZn1
V1u+YeoyKZVy0/+sdXZl4jP5lljdcTP0Vak+bMuRfHGmfGmENR1HPtoWW3LPTAtV
t2nKDhMqzje7HpqtSu+8xwhLjVOlyJmKiZny2Z07QlEBGEphDSfeKIZw5uQABJIL
N7e1aYruf7yQI96yA2R5+QFRVN5rQkiInQX6czEL4seJCHDnci2t7JpYp98zDsyX
GzZoY9Si9oGibURPcr5DRSxvmZrX4pbfPZxR2tbwOTZNGFVzn1veT+2meASw0f2C
qFW2hh9d1clDL0GO0iincw30comPyRBQy4JLvjr2CElIHLnwMLS9Ulkn58pZTJpY
nCAyV/ihE4teDa+hnninJlb2vBraJ1fs7PO3oay9FvOGTT9INrdDbGvcbreEFYt0
ukYVZbtLJJDzx6bb3Vq/+3Qclonzv10zoc/25TLb4NAtfxMjrUbX1DYFbYgkNTFo
wzJHbVK3E2R1sfDXmIil2ZnKn2uT9E/JncLlkuXDxhnJZABnfo+SfcB8Ik9NgNuA
VLeVZmGdfmllynEs7UK0kP5mHC6txheh+bBCWsrSto20MjZrTZzfX51uYxmeXAuJ
lt9ufVh6TlHscZG2RsNABopGnB4ERL6RzNnaeFQwwlabPqZgl7w1HRZVrXBkIyMC
cIfuEsgVrS0bF0j+z/YCTTL/CRLJqOqYkunHIrje5PnHB0OEBrkUSv/XSs7cIObW
iViEcOuaplkuHv0gnwOpgXlnR0rwPsLJt01698qolxaQO+lT6tMtAIVuJ1h/5fkK
enU+gMe32NlAALxHzrWLrG7AwIJOAiVRo1JVEVIKHBEsDEZYp536rHuHQix3FMIi
cl8jaA3c9wWHyjSUnL+xJASuGINloO6ycKIE4/S530pHwGXCYc2Z9wwX949y+p6c
uw8fcM1K8iaJqI7D8dKTCy/Nkz9uLL0fODO3hIq7iYtHQZjJpFvmGiM5Qu0yCPUu
2LbiZzKOpmhdC78lNbnpjuavzfaA6svgiR50gYv4cD0Wo1h6jpQ8QkZVgpjkAmEm
5RgHIpmpS6uxwxghaVocg2w3IyHJ0xfefIdzzUUmMGlwMW317jziAq4O22WflPQu
7TdlMNi9owl9oaE1MG8SKGJL6vB1VcYilaWyoOTn34IdNA89+KUnMlnk+1Oy4tBL
ZcbOQiYrhkWBbA439aGL39FY5ToidXfMA8GndERn9lPSiBg46NC4bkUqKkrS4cqL
AV1I+Io4bvVF1qscn940KSUxkshSXSfR3JBPdR1dx4spWNvxdfyUpmFsXengbsSr
9MMA/UhukbeQIHIuwcltQA2vfWE50IxSwn8F9KsDPeghklWGM8A/424+eAhzUCh+
0nSqVmRckYV14dRewlhnrpZ+VL5UZy0jDEaqQ/IFZKApiuaXoJtPpLKycYcDiimG
1QP/x6TXMP1dy496UEi+QWylNiOD+3pgBhU7WLmsbGixPSRbSsiP9wNuKC6KAOZX
uKzzqiwNKom772uUKWRTnFATIPsZQmUBAzRQ+m8FDkTp6UubmvK+bRPHUEAPr4ZR
orDSHg0dnmE+D6CDHPTr5Kkh2RDic5/p6G4AoohB+EmlaFuPphaCA5zrnWxYzVvu
7Ssf0IJRAUcvXSoypbZGH1Q4F5HRiy/tgvjDyYxP9HOy6T+Wioa6s6liTMGZI1HD
dZH8pi/sRJd7J7f8whXt+U8oTj5jyYGh0Do5UuA1zyyeAlJeCXfx18ERHl+9n5bS
uZD3Vo7fryD+f0leaKmYvMAUS9SpgYSPDL5yMPwJHWDQN47Od9xdPKX4H43RXhXE
2J339qMfnG7VjszR2NS6NxPs7gpZ/1U8KtOgB6r584otTp9nkyPm7DDC2D8XOlbF
4YuFolSEnSAbSXaKYKMAZmkPBcc9PMk3PBsREt3G4wUdmH7WMIF89807XQR7NSsw
VNj/7t9K6B3C1XfkexTFBDsPJXfs8/mdqu8+b/iRrlx7OJtDUDsr8mlP2pPOVp6H
WW8k2vr+LsTKTtTQVzs3VgURWnZdIRowYFv6jJ3ovVsvbHnEhZ4e4Jc8kUlahpzT
jxyK4Ij5g+ya0+oGNli4b+IHOFeOcE8Le35P/vlSBITdfCD/Z5e3G3OmcTOR3zIo
2rmJzN3ZD3vQb7uGv749iYtdQuA3Yi6Dy33YxbABhjIbhFTDt4IKaU7oig1WsmSy
j6/VM3TT0ucMA+e/yxnPolJ96Q9Cwv21ELRmF7fag7BpJT+5x+GsdxQO7y3PdiAs
0x6s2eg8bCZBRCA8lbGaGzIWE8EzJXoWZNcmnL7/6vD7DO+rbkGHSYk+6DXqZfRq
9nl/d1pUuax9Olkgasu5TwPdht4KE0ccXAg2/3x5M7+Iv8CMU35bGCMo6sBMmjBG
5x5HuGYegJQpafyLAWt2adqrGFtt4TaeQebMYLDOvsFY/UqUn0fQ4/tjJmm4ON5g
gCGOvyOPHTeSmwfa64G5dfJ6dBP8ClUUh0mrc0sNHwVcop7fXx7gLf6rLVQJgC9e
T4+8xPDit1K9BfoZ6HfxGFDhJnYbbETbof945GEGQ9qkg3+gJ+yvr1gPFsSBRYAj
vvxNqpQc3tydtrGtPE5ZkK6qynJFDF92Ng0RrZbrkjcz3eYmZY7sX6XZRclhk+3L
luQ+nxodsVE5pY3wCrjzz7+g7ZOk4IxCT20XT9x9+3w059VNtVVSfisNls+slbnZ
8xi2OK9Ho1V5gGJ/xLoMm3Y+Wn6NM3xLNnpiPTmnXShFsSLh1bhIOb1Fve+4a9Jy
/6Z7JcGwMR0hjSWkl4ZP9IINe/RWiTimZhG+2Om9ojbQi+ECHZ2x+x8gHN0Vno3/
eNBLo/c3KBgLrsr3RJ4/8eUNCibINWlMPPg1IflOmR04/9+vQzZSzAjrvICvM3Oj
WPkE/G+zspIHIbJ2fNoMgBCRjfMQM9ozK0sqiC9J67YkitxwxMZKauCCCZDRjB3f
lYXB0oz7GmRSkHfEMbtdckHecagUGvQysiWxerC2GVq2LoGG/tMUdD8Mt1/9Bp+I
ktMYQUhJdbKD++p+aLnZ0ztOfCMuXE4WfhIZ83VJBOe2bXIPxKG7VbqB4BSjcHWF
Q/fiCIDIk1KBr2wqppnmQOmZv+1XaH0BRRRgmC+8o/+Kyx/pviarjEWsrgzWLM+I
Ep4cBHf3KMkGO7sfMpX/xr1okLXX6Z1qlWqcYc8AxmTvC+lXnIHpweqx3qbQ7x9c
gdNiThaR6fSA0WLz4oiEQX9MBmWzmb50dTxgbHcNWoslgJLuefmMQgtHXkqzkiFC
di+Q5DwFbxbz5wqWJ17shXn+50ER8Yii/7FZgBtJCUFwzTeV5HLX67Om1WEea6c6
Q0UhTAcwHkQzR/GFBfP4FwqgboCQtlBtXoRpnyHczEtcDuGMxL1S+Tchhq/zyWZ9
4m1VulzRP8C2gpMzgdDANA3UtRj7H+MGu2qvM5ttnvNyyVTs3ZdSrEuy4Uo/Hafv
Yq+bP8h+4K4POa0Hf1B5IRScFJBi5rjE+Fx7e3qUASVcuk3kbpYVvkA+OPI0B6Iy
adNRnj0my4PqbTakhvAyJaioFJUAadXkmCUjm0ckZrCzhyqc7eT50gD1QzIj81ib
nmqk/v/Y3UY+HoAaOAZEsX2uAbBMmabKc8h2xO7ufI7E3WIokK7GvQaaiX56aevW
atk1zwiNS3Th/nEIct+c4jbDlt35oYC/SHeXJ5CZho/wxbJu1l9SAouG81i4OUW8
phdshDQmS28E6Y3pvn4PCHKn2WSTvwrdP5ajFVYbwSCEuxoc2+B4ZZQGOa8hT81H
ajrCo2K7KNQiz+jd6/uIkdyOpF7wKEqqxnQ82GUXPpMURHMdE4yqwE2d4BnGZ+K+
pOH+nb0HYeOCMBZyUHxpzmZvmpsAgIS415rbBPNLQXURQzMyoZTmNKmDCuBu2BhR
BTVKEzJcqkpOjRTufc+G0uO35soQqlv4WsfXlwqBTkgS2KPuu3PbpQP2XK+58MSZ
MW/hvrD7dqasq6mJr75CYqt60hePmTw2v/z3hqgssAc/eeZC3l5fXNjIpNxEwunz
HTlHiJ5xV6dndyTsrrto0YeC+q9x5BUQ2F4V13HiBqH1/qLJKtOLq+I1AIhgBaCp
nLoea212GAwAp5m3dQ8yTSXog851NHYBJ7Rj41z5vap5AMYfF26FX1cDdrTPYZXt
gaHTrbw/JNdyoIUcVS0dV9ZiD6JuxU7Shs5UC4YdwVSEGOfL0I6/cAI4Y6S4hbcI
UyVppo2kBfQEMZ5YnDQOVVBNQPPchbIut252LQGYzgLw9k7QYA/hFXG7ddwvSNBz
2t4a3yYZ0HzT/M4Ly0yilJvcrYZaKgPyxglBtc4gZddzgbbhFUJ93mnruTdpZeUE
VLudZh5X2/I7AnnE9v4WmpY5FHQ1ttvabkeqKNZ3B/WvHm+5ZCO9IFfvEeKihv50
XeTHG9jn2urEBedVsIP5OvE9Oogdva6P2RZlch81LDNMXUSR1X23d5Ooxql7sgTF
JzjHnKzYxlriZ7iWiBea/Z5AZB03l8tEshvsUwCtzxQYbgXtYgfhcv7pfupWBovL
x5c8aMAS74ZXEJ5owG6tT3KYIedewctb1W0dP5dmg1exY+V/GqIByw2K1JIwpYMT
nRWvp7qar4YHjm85zun8lOaFN7+bBnXoiFA1JVeP9b3p/vzY9rHUcPFR+TiC7kVx
dRMOq1pNPco7TebXgVUUFcXXEZWcxvjozoeax7UhwYjUgiWwz1buKGtX2qkLlxLG
Dp4Cz0ZwLBD9fixBhmIQGZigRRIBG5l6+knki6Wb2ZZ2h415Fmv0IzpiP196Lt5h
r1JRCErhZBQqgvpOZcZW8Zsz/7UcKC5WfsntWRe0e1mUlv/lgbCssytKwsYeVdw7
5lBB6EHrF6Lw1WlwsCwq9bFK4rAzNSTkG5Dcz3VObbnHsJDcinUh3OTliX/ZqXZB
/KX27JzUbVR1tu7cPJG4rdmvsgimZgJyDPnBgRMfAzI4+c4eJUREgygoWSJcBYP+
0i01cVbIAUmRjs57t7m4TEJIdpDc5wfqnbGotxO9ULoYQrb09q/+4ZE4f8MJnnCE
scBCOkRo2tO3GFgPDl1voO4Wcvp5akRzVVRwZ34IItdaUDh8XwsvmCzrcI9j4XFz
xrv/fbJbrmQeKOjxKYDhdLnIAjiQd4ry2SVh7qQ4YvVfIOC7vZrqMySS1M/3zZuU
5Fn2vtpiXh3zdHCZQdXWNKzfyteHtlAJ5Ri72842B2Q7GnKXElW4q2GwA762042x
6S/EVKL5pqK4CyoWnAio7RsQBiD2IECSj/HXGBjGBEcpCCRy8uRCOucV2hIQQ1WS
VxxLZV1zNxiLhSkcctWCCqhrPfEqunzOABSb2Cp3hNZukFws/0TfJk+qW99I0usG
`protect END_PROTECTED
