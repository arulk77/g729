`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveChYWf7RbNwMP+7j9T6kfQnnf7foG5AjE2IO/r9/sZcx
73RCEprsukgD4eymijYUqykOA0o0NBSINSQpe2W//DSldGkjkwoVqxM1ViG5LOjO
p9uq8vUSS4WuXoG+2dfq8Tzxx1xVsnuz+Fml4dif0mMQbj/AJi7ippaP5khAs55j
faHcC/zGKOtNbFEBCmFJgzw7QhD3zzDD80i5Z7NFIa0IZXQnylG9XTu+wV0dPOtt
XPSRstS35HlRXUbOkhFFBSCYp18TxRXG2L0QOTQ+x4Jex6wyLy5n+Q0jhywewb+T
dyikhnCMDezrgX26bgmckg==
`protect END_PROTECTED
