`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JT58FtwiBEKb2HZZoUPZ0IhhKXs1k9CKwE3trxugxFskclclQWEH1FmUuROyC+Mj
qnz7C+H1zbNUNEAkZEF3043g5xe7K4IEc6VOWHc5EQkvHvK2+r2/C8haPEFMCmlB
cDTOeVzjQocjWJX9YZ5cnHrGcuvyEYeFS7y8zaQsFOs=
`protect END_PROTECTED
