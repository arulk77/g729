`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
NBIlfb/a2ZgeH2lwc7OlbdHqizfLVNrFnAdaCiEm9JtNpyMjXKGwpB6vgIjklKaU
SqeHmvA6gXSRM82n1HKGM7DVNKa8KKdUAGHk+H8tUhw6vTdXKnVuBj2cT62Ucg6l
ublSG6G5d+PUt4P7ZDlDfquOuHGFPT21QwddmOxd7vMssTpGpKfFypt1gr7iPTFt
e/RboPuuaHMsjB7Vj4uRgj2hep6S5cPchNGIPawFKXaxqvpV8y/MjiW8Jbl/UlO0
F9u68KBbYRZHVtr7dcm3o24mM2U4cSQca8jGhat49jkW7fACubYxxNRYqRHiywH3
p4ffXIwyUecevTc4Gjk1ylUPrTUpWg12Sl5R/rUov/8=
`protect END_PROTECTED
