`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SfbiM9ie1HTNo68dRqd1AWq2PT/JhO3+hs4Vjjy/T7dn
hQuHtbbN90UQLH+t9hA13qOxRPXbjhOEQOEkI/n4jyCQISgX+05Wy20SKhKcOKFV
M92ALWl3UtH3khZWby45ZPEErfHjQLhzVhX2u0lEKyw69AMrAJh4S6Lp6TkMH5Tp
3C/KFGLkEmsuOGTWpC4la3USjsxKUN5pHhaptwfqovp80ItN3qe60HRl4nKELGWM
ICC9q9xo1Msj6j1D2OakJoWXwj480RgoEV5I9tYrcegu9ZUQLrSmrPQVnd8S2gO3
3/foEJ0OBBuyi4oDsx6ynyNaw5pXaQPJ0NVUWjWhhP3BqzvH7R3fU//rNKlVN96l
2lwXbNYpXiplQN27eUyUak+4QDXO7/XEXmY5nYVBTmhaA9KsCx42HydRQJvELs6U
9XTKJ6hE8MSDemG764t413XTP6ua98aNfLlwjPuymBqE7VuoPM8u56Xjbn54yfJg
B0GsgefvbQ6b8Rdv4M3B9Bvw/IKduFLLJk3kGe08gfbcVnRXzlWrljlRejFKOGqX
AxaG3YoshDm02hJgPFKC4ShHwoegiinq15/R4ur0YA0RHBeGUqajvrkoCDVbANn3
vpv5ikiaQynJ3Vbg1sYHB34F9491Ko7R6ozIMZAoswycN/nNIhHgCA7s0sZ2g5qE
Clf4R97mDKX7+y9gouU4bI91L75n1d3GfOPDwmXqjEKx7uAfPrxM2D3Reeq+jQoh
zu1aFQINpExzGaqlTEGPH8GswqS/MGNIyXjDVFYGe1suSXjB1YqYubZzxVrv705w
f+SsTqB+PEihSgTm6vNZBvGUqin9+ahAQ8LXNrFHYK7hLwGolEg90FmHLv2dlv0f
jElw1xQgMBQv7LFxBs+/rdIy5IZdmzwE+GWH7/m3T8dvgfQUjaheqxwb9Iyg2ix+
PXqYPKO2z/M3KSAAJ1nv6Lww2SLwGRplRInLVTYlYeA2V3MN7f5Mf/8xbojNaA6Q
tSJkRKuTiXi/9CAj461GahnxBq1GnW8eSOV0jQbNBkog3knqurzA2aZyyEfYo98s
qQORhdrPEJlDwaTEqUleTpULa9KVNw0bZxQXoSo92lJuKC4/lVfIkRGCYvJihjJU
h8sJZ3pkMFvf82DBqEQZ3jYspaSuvei8Eo980rE/liyYqEosuvWsYQTlF52rcApZ
wlYmJT40G1a3AXNES3UWVgZdRm7MY8X948ryTlPo/3zcPH/4alxq0aulFauJYTSA
GrkcgXAi47ux0HvP67WO2XmuJDIl7J+Pbu+/RnrsGCIwU7gUWh/voa0AU/T29RSd
acfem980pkNtvB4N86jjqFwRtnlFmxwXS0Sl1DDrHsB8ircbBm1s86khpmakZdA2
S4kPY1Ed3QvYuaBCZQc70IEYU+i9HlAfF47JyFi9kOB3kNfaBupRJPFyMav+NQzu
Z4Jnlc2a2d1prVQIg1B4pYQITrKKFCf9oF8hKOKsQRDSve8OJjPYyV7PNJOkqJOq
ntrulfLdrf8GMifCOuHhJBXQUsjMu+7rvtRo3THVAL9KOSJ9lm3WnOEOfDFdmEQB
JM5TS1CiCf+if+U1DSvX/M+T4PtQk4NtU/GKl/7qeVzBhs5h6j1effaHDolHWJN1
`protect END_PROTECTED
