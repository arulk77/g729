`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu486GwmFv5m7IKMG3ck4YcWmpBOt0UCKrINdAqwN6tWWn
LI4ZsedsbX/hHg/5ucPeBXbz3cvggIPB+yMa6+ZFcVOySlnqJgr1zc0XvCMpi5jw
oyAt1FjS0I3bCxc5/UaIq2OV5yVXOS4tpTPXjZoNKmAuVGAPc+R6/lQNMWxUva4C
iKwM33b4FsY+utNclrqFnNFKvdNn7m1YEKTRYWWRsyzqQfq+0J5rYholB+YbUaNu
JLUyDBoXawVpgKRhO0sxEFce3+1i5RgTx5tvhnmXBS7Sq/l69aw2gVqjRRJb3swr
q70aFmxEG3SdFAeDCyjkgU9NvImPnr5cNkdhQC5g574bLu8JaSOeXtzRoJe/g/0z
paEnphwkbHce96oulU+EYvpV+CmoUS7pFYrCSG6Z5uDti9y1+Lfut5bwgXHXMHyz
B+O6QY4277UrWihlX/UR220Ph6Wrh6CY+2xQyn+Fv08nhiF2pROKLDJY9/eqwP7c
`protect END_PROTECTED
