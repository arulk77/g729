`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOWxP2s1ZrAmMF4h5sKLsJr0JZyzSaYfk6dOnJareQ4U
PsuFFzp8W8ZM9xus9RAIHcF9hfBVmzquCvYHgFeK+OgNMzYTT4wmyS6pkxb5IFe6
r451XjMzVHUzXN2tCTV4KIz2a47c30RQ2NL5bwW4QhlegC9PXk2iNuGIf2uWKHqA
ZuQIQIEnXKR6oEkq65GZbWDitGZuRstRFUkx9bIftKJ0No9Xi/cTP/mr5a4jQ1Wq
BtR72ERt1YZPyHVC0V1br1ojNwiHAhXjiqSF9Q4A/sWsZ2BKP97EYfUcNAPWWXcz
3y+UpbqE9JAcDJJz6FZakg==
`protect END_PROTECTED
