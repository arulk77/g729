`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
n9h6WtB/1yTE8wOasQ7EDCMNRR5n1xWENxzJPlpdJGymb8fe/rdmGYKjkwRxgpeZ
AwhFoFpgkiAHrRDarQuB2bzPez8KTIdp4fwnWhfhnwnmO3EFZpwA9D2Y6ZCbGH37
qJFjWbPe5d0trK5f1rTKKG798IhUiAFr3rj1Cb/U6nnXLQI9q1GNz+Vze1rBd8b9
cQrPP+C68FoddtG8xfVVf3K9i3sheSutmGCJdwMQGefkITU0HXQXuSH3Ro8T1S9A
oSRta3LTaq9FGPkNBVL7OnOTY2sXdaN2S0AnNLeZOpj9LRUs/VaTRWX4CYU+xTo6
kZcyA956Tsl42JQEAga99PTT3Helpf6vgVlUUaWFr/v4AvY41QI3VECxOR2hbaFM
792T877F99hCdUwOeecdVlS/g/q2mFN7jslH+E4o+kmyOZe+HokZFd8RYMzjzSTh
xpTgtmyd8UTAvj61fwnLzZB8QkaacP5WpVpGwe/kFMTkdaXeHguM999oNmFni9pS
Vuptyvjh6L8qiYDgpz4SYr4kQLL4ShAK5llGOAL2hmXxrNk2U4DCpeX9drnT6hEX
eWlOHARkntRWsXAAYUVnCzmfQssnGwH8eLRBBDU4zzAOzKmUti0lElRh9EhJe9kX
DdWYhdqcmuYdK+eSK9JwyHoZosAVG8j8Wx/QspVHwGMso1wB6j5TykKAJorCMj5d
1Vwy/d1T9CJtNR7hWXVT3vs/SsI9X2RkUB8i4sarTxF6wETAqU4H6f54fVErJayp
e1Wm32xsh2b8joDQyqh6jmvoaIEhSw6fVimPw7bgWl0mUHXydNrajwNJBG7Pb5pQ
8P8F5iyCuVLcK6mWTO0uICZyJhOe0zLVvhbYu2VS4CkFFuohs5Hi2vqlQjUmnJlm
WFPbpUOJGfcqkUcQYGoAFnqgPKU8CojNNKRP6ITzDqTls6gvWswOUTbog4/1w/kJ
idqZ2UemKHOgU4qO3Sydrj4Ku1l/N/0X4eQ3HbA+TIoqnl4IkrXxIp8aHNRcTY+y
VdYJX/SWussrBJdYlT8hBuARUxSw8+D6CRqdOkQT9WIgZDT4u7jlfyCudds/Gr7X
s4vyfKdExxrmJal5OlamLbO2gw9vd0985YZJxx/SaS9QslsBgaRr3xb1fhRgPS8D
/nFo8qDWiRNXFWnggNfIgR0x310P4WyWWED8lcSrZRzKgaxwQBCB270xGhy4QIDk
2C7RDcT+qRvWKyTxoiNXS7cibO6w0ZSbtzkzNOU4CnvI1g/4nGuKOfxeIzeW/gav
bIC9hI5mM47Bgmlqr0dFM+HDZzhd1lL1gvAjWLCDyxu7Pn+gHJOC4B+ffJaWGF0l
XDD+IHPVa0+ld4K92sNijSKslMOL46UAWaVRXUj3Gw9O/6EBJuw918cAZsKhb+EU
TFPyoobkLYz6Vk5rOd/OnKyqW/iKoqw5XVEZgavJE3jsjr/0vG66/U0N+fAd2idh
6sq4NMQVHmRWpoW91NrxyfuRqmxDqppVf3UhW5G80Eag1q9GtGq4DLl4ziPtbe1N
U00iXKDAVskBUYv6YOi7NyK1+GvkOI/11gFSOZgacdAc0HSdKDC/5yOK8X0zfICp
XnZ8bp9w1yu3096PvmZUeMQrlv+geDRRy6DZMGDX3vqJWLWd9Fp2cElDxmqpIVDD
fesuvxW4iYJaiM8EnHxuizAjWIxZWsGuPBMgXDeHWS4FD+ULiTHCdxaaWw7XZGKh
V/oPe/Q7jq5Sk76BRT8yv/c0UeViOG5DAOMewy0ys+drhCyF9f0C/p6hy5YAGNBK
0iTJ6YfiYDbKvDi/CNhfUAT9B1o6p4sy8bxhaFyieiYwabf65QLtfvxl+VKzMUFQ
AT1UbH3zfK6TK8/4n4jwwqXxOTuYkMTV8AaZYyg1WY2asgMMu0fNooHYOZb6uNz4
GAx41lVAq54NgBwCLt/n/2maGMHdYLclMXsPAYQHZB2JzIo4GtRoPzVUd1UjnSXj
Ffo1gOAurNiWzAiTJOKj6BlpkMB6ocd/KzUiskkr7JiOt1slr3Pyl6Zv8PiOhb9J
qxaE1ZgylNHAtQCMP92rkfmca0JQ9iT+3BVfBhdgxpbLk2eLbQAXN2Aod9YB/DUP
wXet3voh1w3hu7YgsgBOjugyYwUKKAuluScmKaxo4NReyRTKbO7s/jnYPzfJ4VSu
O5t1ExP/8RNgoLAQ/HGbqxCJH5ZdcfXMqjtozbA7VYYRoHJv0pE5KqnDgbWz//16
AqR1qVJjPzZmso7+GUkAkhBohkZoU1AX3pUJym/lCGGRYuLjC8ENBrNVvhzoSSQN
1IlobcZEagPCupCMCtUMI318OhnE+iueNzcNfZUd5bY9fWyqqTOYLPKQhvogXGUB
+N1ylR7WBs2W2lMcKfTTIn274YqeSzXUmh8ApJ0DrhpdecknywaraakjVpfwtSbo
xNcCkn0TkqFBt9muZnmnQFfOpwFVuqEFGV4yqLLngSPXh5UxuV7f4Mppg6kReHck
h7Q/4H8BxBH9U911gDqDDF+3bkF7KRc/2q7wfhj1k1BU/pigChR2QmN7BiAhEw8O
IL7DMZJFAAhwB69gGxSi3Zsdd1Mnssa3saLhnMHZKg4l2lNbu0419bLwfq4MfhoY
zf+hquNWtWvotitJN/wkyma2wjnNPI0fIvB2As/kazVyYjn6KVZMal9wJtX/t+60
k5K+AR5EHbHs/lUAOc4CfcD53mqdAnSb/+mCeWliMGflQfUpg/zwV4P4A6ATgDqB
eLHDT7BNAhqyanzv6VMH1z2B9kGDxZUI4/BlPuVnLK88D3w+I5ZU2TNbgs3Q5hUT
IftEZh76XUrEVmY31Wde8/rS5QIYy8gzn883xHNHKvb0xPPmxnGpZ3LagNA8UC5W
r+ibJRE9Vz4/BmV2uC04vWqxdBMCRdK7uv0F2gPrCSVarE7hG8MUMfLz76u4Sb1D
kHRR0Qw3JkYS02/wm+oVF3/hfeEPGj4D0+fiqoMQKhaRF3PkiipKCtmv+eExbz+n
OtAGCcQUq45X/mXZs6h2xVNzFCRzycLKeG0EvuBwpZ6ONgbK6Y8sWEiwl5P0+0xQ
KMiwOutyjg+7VmeTE05tA7tuMPJkBe8RMF9I1pVdBA0z6ziO4m5n4OzgAmz/PjJA
zry9HxQ0TmSRRp8Rt3NvkwiWJAnZIEft0NtaKBGx/QDrGXUoVlVmF4KtwGrTnPlb
JS5KCia+QMxauVz8+Sw2/OHqbmnJkK8JrJsyoBjBew/iPwLDBvuFIdJglqP+Bcro
WpoweZpkwPTQ+k24PZIrNfcFckRLXi01L9im4PyCQIhH3P2Ac6ZCaTmcfWh33s9T
t6hPnah4iy7Fwyl2xPut+GSb7KB4PzZZvtybH5wnbjErSt4ChvSO3kr+WijBFjzP
TLpQQy+79PGG/gIlS5yRtRzo8Jyv8XpsDR0RD2xkkkW56Ga6E4F5sBi0JLezFp/I
sEMVAIPIWWXsEsVwVx/U2YurJmW4CQSz5f+dJ8oT+SghqY0uGkF0AbYQgs0zvQdB
4Mj9sVmO2iHyVx5xiZXoWBnGxlebVGXFHjJIzHoF3jTwyoaBDFulSz5UW5K6cDdn
CspKQ2fEDShiqAwoOwaWr9Dr+JAQZiOLrh9BoL9N1c+LGplAAkeGLSQUk4F3Cecw
falqSJ4ZYPJJea4lAzYUSF/20Rku9Objc3lcHdfUwnTPfMP3OUp0C98v9ek31mLq
QNGrHMCieR77StJ4Ba3eff+gsGtldLA+Zge6pwhnqMjukQ05IB13ttWDxiy/pyQC
xx6mT+8xu2S8VYZE/8FelDc+5JT+CqvNhruCoHGrlTpfTTYq1qUfL3HaYZEandZJ
FGWEoZM449MTd+GH5/Mbmw2u8XljIyysvBFPJFu6uMCuUpdQBgy/QNluHwe2r8BU
keRlsOLa9mlaWZyHYPcK1GCtOQjEI5v49iK7x+SymGHSD7pCcW440CZSeN9a7vmJ
9dCbr54yBmWO34RiVPFmYMKZQ4lRC2zd1CbQhQw3BI8FI+5vhvNrI0hVfEPal1Ky
vt4shCu8B/uw/kgo3PxAnD7DXZwQExnv8abtBop93KtfB+nQ+ytVMja8ZeaaxlkS
9ATlv1EfnndYl2gPsRVeUTXNgNimDgI2cOQqTiC7lawKHCn8RtqzxUbm9Ejk3rT1
xZvkoErjmgXO4SFF1qDRnKgGbUuSx8Mgzd5WMa1U9JDH2lrPs8bfPy26/sCAvY6R
YyfWaY474jGLBA1tCSnFN4pP2ZvTYkn2FmKO7zylPD0PW6F7kroqO4ytfNKAyHU5
TrOYM25UKTrZFnsvKGu+BWCmr0YqC5OEbYo6uD4PpCw=
`protect END_PROTECTED
