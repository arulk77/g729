`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLdnOo9dFQEU+pL+DAk0DkEUb0/5Cwl12zWj0gLu3qUw
g5SaH0OGI7p/dydwRC5/5Lax5Rxn/w64AiYG8jjHOO4SdeS1iDK7R9KnuE5pgy18
vpzx+xaZ+LmvYecxX6K+4ad7ZiC/JZ3McQvg3xZ2zrhM8FlWyFX6okJorT/eczpz
qvDzoIwksMSXJTyoVHyACkFfN7plgy0eRT159YGkkF7PrnPWbJ0kg17iX2AdGzsJ
`protect END_PROTECTED
