`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SZ3/G4LjY/wUuToCH2e9fgIN+K8BpLqpYufjqw72wewN
HdtG2MjuW0jT2FfjXYNxAX2qf7nuHytxBPIXu2QVdtIQe+6xLdmaBg9Fu71jTr1P
S5QQwipGwoCDTAEJmg4l6QPOZKCremakwN70RjJq6IX481p/sOOgHmoOJ9JAr9fu
c1ECi0N9FsPXSipbPvbnPr+OI7QlYxE59F/YFGkcMEbl60uJ+UztpyLB4e9XOix3
myn7fMQ53EiRe2AQdvZKrUM8VzWOMdde7nB2T/VSKbJNRgAyOTafoBRHLj5T/Jd4
r98DcfLw/JT22jRr6kxM9NbmAzLcGH6jb1T7/+u4VpPPcSJBmcKmRGQruuAMwUO5
lNVOkdpImcpm+FX0tHmxwrAVIGtLx5wvTQS/SnphtG9fdfXzJYcUCixk0yqCK4L0
rWrYS+o/dM/GScV10XOyKqT26seZd/AAoTraX8N3Vtpzwr85b1umBtaBVLpA0zji
`protect END_PROTECTED
