`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG6U4iNRFol96JgGklNXTumhU444KGstpZXHEgOoQ5gU
qIw/TCbI+aaQZZg//Ao08i9Vnlctllc/tJkLfaReE97YMAqES0RsxWHiJJ33romY
vR1LTlUJ9RrG2aNUINt8YQb6zZZSQQwiywAOZ/ARjJmve2+Lwh11qW+xDgAJaLRk
2cagaA89tcUyJeTEBisglJJ2Nw+uVxScNvgmFpNSglYsjw42SaUMYvR2/9u9aupv
ztqFfK03t7Paub12310QQtxFZc0NKMhFazlU+R9470YeGZj63JypM4S/r68JO5Bh
ABUODMHMdohFwIohY3qLXkWVXFZ1UdaPv45jzmVqnobafWNdNtANId1zCbeqOlOn
5BvfJ+ncUuucos2A2IS94xn/ITRVYjn59wrlx7cSE/CsSJOV7xCoHI80rRCjjjnO
5jo+3NU3kDa6YgmGGpPY7xPklOrK3DE1H6Ov4eFb0xZwx6z4vEUOCGufz/JT0YIn
qWYso4kAYJxj+TuBj00sxQ==
`protect END_PROTECTED
