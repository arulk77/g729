`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41Bt9/8uXv0kAou89+TpQMrSMGeUTy6DzYEKAUgdxiPz
aK2bDoRyxDx4QZaewUOKuSZL1wSvJn30lcnKKGJ0ftldQClHtDRnGKr4JH4AhXSP
NjyM2OBlSbgONiv9seo8c4B+UGppYCfyLjNVATH0Cf/J+qqOHbj5yw6q2UMwgkch
+/6iIuWXskzsAtpRFv5+WmMid9ytElfjNhb9MivXMJIz9VA5lPIQ55kiX3NbMEY1
94Ze57zPBn0ZwnR4TKikRirXZuEnHPD/ARRfLX3C7FriNtFqwuFFqXCcFAhL77Br
4PeH3Pv6SJ1+C4vlAGVSmCNbPbVv57vMHBPLye9oF7iIPc3sumSiX0r4CcVm6mdu
c2OHqoUFxX1TRFOz6EXvorSQyMCp2zPFVhqIVWM2cH6v84ZMyU7AKx9IvFq8b+2/
aDbxAhx/zGq9wkgtP082gsywS7YWIfZtc8ecYkjNNnMioWTrszikizybNfrw80w8
`protect END_PROTECTED
