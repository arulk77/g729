`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKAslCqQsREZvgoJjIgbYKdwGZCakkpvK0HCBL9gvEP2
akRNWEE/mbMFMz5mxi60tgLWphNYytLTk+S+0Yuqz5UmI3G0+qEsAw0Zas48tv0z
mJ1PLARijLdDb3ElmZTkl/HvffshQoB3LLdrnN79jhga2C2G2oVSHzzP5WHVrY+4
0RpTzZR9QpnSlO2hhJRFvELV6flhVpyrMz35cS5FhyrYcwAQNOxTzVDVb1mRKuw+
7KCYF5qHAjM78YHbB2lAlWXfjWJEnqkgx+k1aNYiKmF7H5F9oCsugxVMBHwdGmsd
PjiqDGjByWFug3WFONvOCCUbjSD78TL4A70g8VHr9UYFmsSLvdtaFXq1VUf7ARQa
B7k7Ygaj6wfAKOxBSS0LtNrRJUffTSSNsHK6npib1mytf6RVd+WrIsf9EnP9s63r
riZQVCmw2ghcvas2u96qcZRSZv8MPLLtnqRFs6YP/aoSjJ3hWl/P3V2wKRfEhcC6
rzDEJ/dHGUawVx3tsWWmenQetHIb2tH1WjNNR0cnO54+N2yazUz2BeLlKwOt9uqn
xeA/I3xtSCtcOSzXhcVcAcq/Nazs5yJqEQzlYo9NuQDslS+MFmCo1vQYkb2pkydk
pQntzpFHaN/K7iNdwbpqCiDAeafbLAV2LIWRZfNa7D0Dvx2+OloqMthbUVSz9OyQ
SF1PQsncZ9h0uteWXchPYaaO1bNIg6MDPB8YZJ+gQs38C/FusP0GxWXpHITysQhQ
AjkjK0DcfxcJpDJTOz67JypkSRiAvTJLJ1qDQwbDgoFBYOY8QLTWccLVA6u7gO1I
FC5a6qlw92ojOqV4EAax0nvdpLFNRVpaXAI2asMWcnpk8KEEoF8CmTpj80VrGnwb
qhbwWn08r9c7FA5Vx06bQRcYZRKdBnY+5opQYr5JAFxFSptuuaiKRlMBbnBfTES/
k5sd7UqCRvkWBDmno6QDl1zsxnSxB15OS0w8zgw/Ka13OnWfceL7AHKogvRUjQLV
SD6nyK/Ftm90KpPUm4QZ+mTt7N/opdrZdu8sKgztrqSxMzaiXnpVgicQ5pxoeGxX
8q7BeSPPL9HmfH3AIyfTPU1HYSb+E7L5I0Q99QLRbgxle1OstPTC5DFnqI60av8Z
DKjENQgxmueGfbkzHZkXU3J1wUp1Ck6tiiuKXs+gi3s0l6UojzGtTiDS+l0wq4Fi
MWHqlKrS06Z8sPU/TGH+7ONJtWX/inDUnFA52STX5xOaBMj4tDKtCKPBdwEbGUjj
wdtuSxJjGZtrlrBik4LukDwhKPE9lX01bZGoiEsOUjkMYcQwtkr9yOn+WhFCuUZJ
xmODuL7R+C5BtGR0UevZswWXfb0eqwEuS/IoDoW91hCjVKPWbAgIOEocCyoTeCh7
P6bKXy86McudG3tqeg6sp6KIHPFb7Q8vTmgODL1HFoBAkPdfNdUiCv6Bl5UpTyvN
r8Y0vqC/GW3IMl7SU0RHgG+FhlABgPWLsTpMgVyDGrN7omwVFLyoJfcK1fPgrXhs
f2HsETdPspNmLnUSO48LVKVn1KmvG6COLjwXiAvJWYPbO8jlYv7q+QzYdmev5LpX
mhPJuMRjq+crO+m+tdvycXv8s9ujEG8PxvQZWWFckSxTYcRIBOVVaec0BD/iscD/
LVLlPXDoImD0yoY3gjGlkdVFp5lD4WrfQmitlNQQkqjn+dTX11QiHjrdCKk+Z0Lm
A6opTRjJdvGV3UO+yaUuLX+/Ln7dE49vYjJ8Ordgnh7cd/hCCpi/MldjJ0Ra38tR
GbALAF3ykSW8CDt4fT5c593Ms1IXyq3lec7qOqigZKpzYLeUMKmGu46Gm0V719H/
PeQflSA8yg73XH0/X4jE5BU+fVKrSgbkBFkTkh336IDC5HGd7OFO7CqF+IFSpCQC
k5chjPojYlz5iIQ9PRUVxTAzTfBPH0HonXmOGvYoRoLB9ijNCxC+UWeJHrmW6oeS
B2g59VuGHdto87OTgrqFfITUwEzFT8D3BGsWvdzFVecMj4Y2SriaaYyPuBDsQpac
WC1Upox+9i5aa7niXFB0tps0fvWb1K0ThOUD3b+DJjCSGQgoiNxkxk7/tZuglDrt
HtXA9YmyOxZQlYYMGJhmrbK1bmm/ndJeNd18dQnXfBQ0cui6Lxn4Ab0moyMbGNrL
8uBw97fyKQMiHaSYEwFodkcx8Xk07UEXZhv81/bWnpWKWOiURzKUdIxdlAblWFq/
5fMmMsWwCRf9CP70s2j8uVwxRxzP78HkJs+VjIl9syssVjKmiWI6jOM7FoWosYId
UhVXb1B4+TKYaQ/Z5zgmn1Mia00Eh/OyA5ic8/5VGXvCMcLBADNibwxUbuTs84PP
VCQYjq8ZF8rW6Aic6p2qzMyhwubJWEJX8DvUvBlEkWEqfdfv5CAdBIZLo5Vy5eDm
jT0/QrSam8/opYSG6aVN8aK5sw+XdjFfDk9p8ekgssy8Y5HqurEKOaJgPAWkQHV0
`protect END_PROTECTED
