`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47fWAsKYxN1+66y4NtkK/6t3VSx1qMmbKmtw+QOqC506
Tz+brlOcXW7tvqr4JKWk5IY5Wz2KrI9fYL+416EyOra68iiIOSvHeRJKq1WzRaR9
iqaljQ2pT7z1kPvYvzoRH2uti9INjm3vniysRC3lrf4bawLA+kDs3x1iv3ysdFF+
besp8mrc2qqia+IwrFWnrWC8alKQPixOVNFKjzeR/nhjgeU6esr6k3VhJxmsx7n7
WjhdpynXX8O879kDlYVZ8aXlY+S0uGIViG2SSKTbzOLyigzIT33URXpxCpvQQDHB
TW+k+n874XlgvauKo3RK393gnB5lIratPer3YvtqjSs8Zity3eDRzZfF0NSSwzzq
wkBHOV2SyTIzuGcnCuX/EKN9nb/pZwscxn6aB4bZXjlvuq6w6uWpu2Z8JsYQykue
EGHZrw9m27DaFCG17qA+ZPPp9xvv0UD7VfwuB1+w3MLjWBcNP/hZSZjNXR7E1mQo
`protect END_PROTECTED
