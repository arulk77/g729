`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN8sNwD2Zs0Up4iuay+PJwHyfbK7s+leXzNYkLAaDmYjD
s5c8ftzv8rkh0d43l2iwerSVcyHdPbvrsvdSGcHGvTZGbd5xdIPCKdxI8eajYTJg
qFadpuM2Ba3OB5+kMakAL9AZHCohP7lFr7uZCp1mWklQ+YOHpyrhDPuXj2PL9w+p
ZOPN72F9Ks/9ZH7nukfVttwLXwgfa5F5EJoMdbyVWK62bSkR9hIUKAMrmm6bmhWf
HpthFEFrUvFWNc1uo1JZRV4Yi5iQLzzs8DWmuTHmUUbNi9BbBasrNCkgDQVkX8Go
A3OUndL0PZeRvN+eRLADbCvJQBHbkuX07xtaAvARcHuDweKLmdoMI0trH5+FZ/Io
UshE9AGrgWK4/550tISRaTVrOUKYB7IVFE10xdaZSEneA5Sn3Jp+xSSwpI62IEti
T/J3waBhhdsQdC/XZ+4Ms4aql5roS6Rq4KWl0hD9MX3SVDo+tybRe1VQfh1ofHO2
EkMqE/CiuFLQvBHbNWXz54szsF3w0vsFX2LQ6NDLmjbwKCyoABshaOaSfcIrrGQB
MKgoqiVHQMN81pfg7X01AuyNkNKe78sAtS9GcM97yqHGqY1rc4JIUkM+W7dnnuKI
9WE7pRIc9dvWPIry1WOrbxm4nnsnf8ZsVocIddb+sEynCsvECSYReUVoY23/D+zS
FNNpYkFlnOqq6KSTAX+z56tuYC0mzZAIRrUl5v1aAj4vzJXTP2u7/XrN3ihWSGIW
CpLs9KwxZhj6pczR4TlBANaj70z0v8MYu83/4xaHmTHmdD6ppQBD8g1rq547VWN+
uk+lvS+xWM6m/oOfeMsWsXXqdVOX2O0HCj9RdSwjIhlZScA6qIcSl8D0AG7G4asI
`protect END_PROTECTED
