`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLCdCjLrTkn+0MdmAXAZjn7ajU3vnnSkfimuSusmDR4O
iiURnobS769FM4PUdqxhfcvVtprirhGhhxPHlpXbvbYBmD6Fznlm+xJ7Oz99JD7L
Qw+t4ociqM6Voubql+qxTELMJJmJmHdsfAlGBG0wnW/UU0KmfcdhMIMMngqZYcM2
Lb9urbY8lFIHn6NnCFPKllmM5pLciasNrn5O6K2BKttEOfqgGv+UiJG9VtsS0VJR
hw5ROY0EIqMANyaJAyinigTAnevSb0oAi7MetFQmcafLy9rVu60G9uQaHix55kpR
OwgNiRSqg4Pip3BMPfSCFLgjvaCcN+huwf1VpFgZXwabwA9/Y6JREyZHSE9o+Ptl
Ow/NdMq8lt5Fd7kkM/c2exx28qHC9cEnZ4UFHXecI37xHlgxSCT+vPHNXl3iHFG5
zo4y3YyTNUhPG98TFyYS9jFKEt7+Fi6Oq6YP+GTTEPan40DwcBmSlYRS7QmRrx+k
uNGhx4TZCacJU9uRdv5CScGN0LTjnI6/uUAv8rjjJSV6gXuqAJ0D+nlztnsz0zql
4aLwA/yFmWY6KiapcIykE7uLc/PP6N4pndHIrafJ8kjHrgHAteS3SFkMCq8ZgSXo
`protect END_PROTECTED
