`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+SKPzw43+5M5iHZWvMI/S+nQHrtO0m2IfVYwnPmacqI
EiJf87OmSWwPJYW5xODRRS4MQy4kreWfak8dcTj4Kv2N3hLOWlemFQUPweBJWOcL
xRxOXAkbMIwxNKmbHC3yH8es8YZPmqtQOnUDxEyWMBh1ImRlcE5uwnEn3Bg6IBBQ
6oIA8FjiHqWuReAjSapq+ojldKWlBk+SnX9/uVwcvqQ=
`protect END_PROTECTED
