`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN4i7wTcprOFPPAL2hfUMF/PWS0h7X7nkMk8WBGrgj1b
bX0MZt7qK9tG54B+d2uycG9RZ9il2+Z6uB8PfP51GH6ajugsQc2c/jJSc0fGGs7a
yOpIw28t1bZAwR2a1EVhZGW1NMc1WcZaPffTjyf4sNQkEZXrRfgZKyI0BppBlGBt
0YP6icWB45nfqmKXzzlMKPL0ypVuL9lpmEkcOlHap+eb4xS2wZfseR9l/hPbIBQg
KyRvp0OBLnt46s0rBFdfqtxd1/zplGZFYUTdqtMdTOMVGHQovglxlzAGnaKkaJkX
cEKrHV2IriPBIB9A/IFgP3zXNlNTkwH7APLLchU53RvHi+Ypq9zSXFQ5r79JcVal
`protect END_PROTECTED
