`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMcRCA4XXbhUqxTI19aa0nKZ4AAKq4q3EBF5JBElYh0M
nmw378HoMZp00GcepvpUPB6NOPzRc2LTeylX8tOjmbSJ68GgaFgAIq3JzCcm/0aL
L0LiHEbeA5ESK0Y74+JP2M//77Vs+XcKlwWNcWQn7QIQvI4cgSKiQHEP/ZpMpMAv
MyDFHxqnJO1FWySpmMQ1Vg==
`protect END_PROTECTED
