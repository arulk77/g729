`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
vjVt7KXtQisEVv46ABFwvfMeb/9SXrNZDMcNJP0G8a2HOHVOfYM38OhEIgasiIlh
6gpJ4oNRxEQXv0YYxukPFMEIzD36jlcd7c0Urfl4FXtBvm2OuNg7acHRwOAQKf6z
67/0lZdlEuS64Hi5Aq07zH3PpI7sodgzlOgdG81jc98IL1usSgmh370iPe6VrIf+
DP7p+lNzZmpOuIX+M/0Cc9w+M9tP7Cy0GAk5QBpKAp5FJCxj0SBKKDaoytk/C63h
Z2ntKxoJv7XQN1Kacx5I0Id8nLBW1ve9NP/J4bH3x6in73GxuiyvkiYw4k4qCxPH
7d0yXPxC50+Gu85KB6PnQrywXJ4qM8bLFIfT8DuYhPNFBDf+XpdjJnYLlNjCfso8
efBfvHksVrQ2tMXiGEHZIN9c0IH24E507wU2r1kjVKb4dmkqv6W2WMEdavwfcEvv
KaIDNraW61koz1wRTAqfZpZKhEymgnLxqqMQNYwBsG6Cgi9q2rlzobZetr/DcShh
EFxAzrvWKlPILrOWc0dCmOAy+gPa/ObSvLqO+yOjkx7Am/QF5ivZLeVdn2uYGpdR
M4kkVMl82eAmnBxAFRceFr4dqv9sxd/FN9LaIsaTGjMLSQtv2cpX0CpJHdJ/RQjY
Ml7iNnMdq/tCmpQifW+DG7XnhyZY6Ob3vlJxUpTcduOGveGV354ma6tbe0ItLCcK
Gt8++PAyl3zwnNXGv7MLfwP6OY+VlyvP7aXR7ozJ3mPB3FefzFbFHwptfkS4ZnJn
Jfyi6btzhK2QS6vPBPcu3D+PlcPLrMK8qKwujavOL0bytc17JTqGArO0/izV6qJC
uiAG4I+5tlJZKAQiWeomBg==
`protect END_PROTECTED
