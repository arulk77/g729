`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGoBg1EhgVUXGCaNA6H27MgLqQozaLY0HqIU0EGNc5iM
Ie4RvtJT+g9qKr4sMB4758mEt/LiHDTPR8VodIEoF180RtgUJCjcYzrLAYiYtvYb
S91n093v5bNZjknIO72ekfdoydXmaT27e4ap9JgwpS1615mGoMAJBFOUgV9hVzgq
n1D4TlqQ+udaqOl6Brke1sYGpwd7gIC1srWHwFatP3Btpl/V9hSHPKcJYaDXNuh3
mIvPwR0HmPDXYs7A1CbqDFYi8A7oDR3/IbnJmT+9xzRZx+3DnGKMQJ+1zpCZOwPa
gapwulwqjRtWTv2kNZCi+oYwaVIGvkgasm0of65k5TYFRh9phAeqDvMT+9xoF9GQ
MdADkRw2jq6MJqOrPK6VtA==
`protect END_PROTECTED
