`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ7vdYMf53bk6Nx5za7maCO4s/1cv75l0EPGvNpQQVle
D70mxo70XPurLxINAnNshP3ZJCvIvkNte7b0Tx76zErDGLfp3U/GENkjIwCzJox6
KQdivxxxAg+ujzC6TC10rDJFiWyK0IYuGnCjKBiNBh4SVfAt/4WS03Gu9JySJO1r
p6dqOyM0F53s/F/BcBGhjsUUmpIe2CuDeb/WCmpOTfqb5TL088oPoYyvc0J7wYJJ
IC9JHZj6OCQCI4AgfpmS7u4FDNdEuWXBzx9+oQdrR+Iz6NfSnplb+8RATpX+viPB
E98S7t03mmpAUAoV8qBHd+2oLml5uQkiyRXLtddNggihgBA8mGH9MIHaKFGBDZR9
eKO5KcVLxIv2JnxoDR5iawdctCRjmzRTpgcjgSD+/od7KPJ98wKysbyYFw6yx3ci
7fLCaYq/+wf971vE9zttJoeCFmpEB4jZImjyy5Tx9Hs5M4LW1oY9qmbq6CBCDPop
25EQEQTG8pmvutJHlSq8mAbcSh+OaaCbCCjhzUVNS5tA5tkIWbqlrd72hCqJOnja
jzd6xh77916SrN9BCmfarYLxQCvhpfTozYdZrRrjbKmGx3523liMe5P2th1Cm38X
wxFk+dXT18UGQRDo1D0YrOI0qSg688mxZLtfWnBXJvOR28x6FckoHcbqyieyFwoy
DPWhLetoDfvv4qAVJU5ehDJPv3jRxvZzpDVFs8CHVImQDzqv50w2vzXJxZlsA0Ci
7zF4mz0HCRRg7w6g4im6id3Z6ng6XqWYa4Kv23zMNkq9SRM3E9T3gF6JQSl3JV/S
bD98NsCrDnxVKgAjQC1KI84CyrePhWx4fiOxFg3mPwyrkFnDuBguqiztPU3z2kkr
lkNC8ofEbWTv16UedfXKMdyE6kLDm3zyDRBNIpSFUVsVBiOrtnJXyvuyx2TTQWhA
E+i3hJdAV0qP2V659V6ePdxSTH7HIBps/KgMk8fWogP5OQFt+IKfHdrsrTXdYqSI
Iks3oblxecWhPFE8JgfWaSvztzrs+3d99ukoDlrITlxqn+jOHQM3cb89iX5xpVe7
CxFeZztiURGjmWpBx51XnShxCajp7iyJBe8EMFmJECojtsjs6wop/mjh9pVGoGTE
3xIlegTFkqNdtKpGmzMzXyGNAn0E8xotJIHYnEeOoA53C67CMbFPIM/Nf35NXbzh
l7eKzTWmo4F/4Fc3uLZLZPPAGRWB+0pV++Amnnok+o+KL8EqEFAAcS1W/8z3qnKb
0GJmQrfxUjbuKwvwUafR9PFsZersxpm31SLy3tagDfpSkW+uFKJE6xiAipXzs/bD
dVaupijQa8rdoE4+FsumLZsrtdct9Nh7LHv37+hKnagrd8eXJfjZc5BJFLiR3+Kz
bbfpgBA4dIGvVRk80h8TM5N1KD/0jOVwBcSP53N4CVoiqb9W67oq/l5QXBI9sdGX
4HJHCJdFdz8E8y1/WcMLhGckIeMFCoIooz2jTg29lCeqmG1zx6IbY4hN70J9spqP
WJ5Fs34bbuseaF347BDh9XAH88Rhs+vyETpA/vgk88WwfItQmLphsN+TWNbYwcxq
cMxro/72qEfr5tneZZHFXTKggwzblOJ9S/M/O5g/bFI=
`protect END_PROTECTED
