`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL8Gx1z7SNKmIMnc04bmvxWZZggvhzZbsvdiozmDi7m5
eTPo/Klm/CYl1VQdCGos+tjimB5Rnr4JqmFWhAbOpnPdPlZg20WF5RIotNhN1p5H
9KHL2DBNQzp9iQ5ZZDsCX40WylJA9tZ6pCiftzbUO5kJSwCksmFCSdXFKvnKuGq3
V+vMmSDhotrQRwSY9qMw3g==
`protect END_PROTECTED
