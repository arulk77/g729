`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDf/5UVLwYZ8HY0h4UQXAs8UlaOUItshOvtwUKN955iV
a+NpTJNEMdQxRDR+Wp/5PR3BAv0zirzJYQr6RieT5aokjMwIzzjZq3eXPMW4gybU
5s+vmPiEzGOefkG4PmAfNx+Vd5+13UFIazkkRfO05qDpzRxsoZmDs7jtc0h8O7us
AEuy9EfigjcDcOjjqDCjh7mbHCzz9iKRrzHphj6+TI8NiVdpBmLp36cm/cyH3ZQm
`protect END_PROTECTED
