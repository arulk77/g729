`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIuX0OF97b/YKtY4osgGhZITi77wr3Cpoavo5BKNpcym
DlMxwyM6KMdnPnIWZoIaZV47FsG56mqc4+iufaq707GwecbIhkbSuXsmyRSTyicV
miw6bugylVuW2ofn+stLoHMTiqkM3Cv1Xi4zs95uBnsjA00FoQZQZcutUIWVL2uz
o9NATu+PWGNeEVsNbGYKTyP6onvwq7qK5mGDLKxyfdMOUKKeHB8p3uazvBi9Eh/q
`protect END_PROTECTED
