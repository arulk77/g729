`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
72DKe5MEZSH9IT4s+0rFcHKVWkn8wtq54C28kuDRFilHO78gMyMNg4u/9kYVnl/q
5kOB07xosWHiZJ2jNMeG/ETO9/huXQ0Ay9imAcEbVGfSRWN1bQgs+jclTn3SQNs7
36sF2SbJaym+EE0Uhh2tYnaZRBHZTmcvTNJOFOMzVQNCLx7wsGNQDguJQbbnl70K
fxDmgV/wLXomCtqPO/FS304UOQO03YDSjBr+OxCIjv+cM0K1eTrF51wA40lJPvWW
xAk8wjvngehgNk5bGdaVqMfiF2oHLIysU6/CpN37+A6CHqE9BlPi1wmZXj0DNl/I
`protect END_PROTECTED
