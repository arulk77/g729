`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
PnKuLAmpR1hLOzR4ePT/K/Nw3C71DECT5WoAv2ZqCe6Iai4aD67YCWkiCvQk1t3I
W3qWIlxBGHOTEn2vtAuIAkX33Ejd5I7wYIDHMWQ9yYU5OO6aE9FcFrpVCX93SvBu
RYnsg0Ljw7oNOmyY1JSMjrQwkQT+mJ8umxSWdDxmfhypaJqteCVI1RcgTR2Wm+KU
tN/DgeaVa6whJ1EHccl7Kyr5aoEm3yopHoUKfzzod4hC3lWk0QLfio/IefSrDRFw
UDYrpuSdF2NBFhalC4Q1gmPJwjuTW3tMIoqVqapajdY=
`protect END_PROTECTED
