`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
C2xTjId+Q4RCJ9QOsBdKlo3ZQhDHhZ4y7Ht7b/5+ETc4V8NvCzcCBswJdrRdmTEl
2ViiTxgFUV3zA9XNsZYoI6ooEctT+cO8DW9dGEGJHsGd34A31P4OxyPW0SWb3wPq
ry9iUG54fHIJThUdnZ7Db7IbTHbV4q/7+aMvoSiXUoJo0lH8NYU1P3/Z/3l/NUaL
ahFGx8yKw1FrY/SIVbLbgO0P76bKAe4kOxMDSq1wxp8=
`protect END_PROTECTED
