`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
d2/TNRZa9yJNXWgw0QUTlns/PUIMVe+j4vEhU3yyhXbx5OUgNjO1H1yMSMEgD7Qb
4FQmQNnfkix6a3aEjDtxvQPQXX2HnLW6PWJ+UaXbhIF2TtIY3zxHQvlOmpUwUs9G
3vgnAcwoeVFFuHNhRez1OxEsLeBuCb8UVmtwwA9i+gHb9cguleOmedxG7xBtUc/i
nbN/FAGTRXgF0K6Fz6r0Eaq39Ym7WttmWbpG0HdYZHkjdS/iMK9XCxVhc5ZW8hVg
sXfxShkeVI9gGRhJ1CTnrvQVp5OJkJF+YNRz1DZs1HJ4NZ/ED86kz8XXJPlHF9d8
q7Am6z+K/ZDeXaONfe10IwLg6Cg6bzMi2w+kcfQxNkYNKXeWcEadqFP4vxAWVHiY
uD3fsiFU3RW5elT8PbXYFahNc3UkvSDuw1DlAaliLGaLqvZa43lNYIKjgFfciEAE
DKdffAOtAA4TzsPXBSAoBB3RG8cfYXg8ocAmbHfOWFI=
`protect END_PROTECTED
