`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGUOqs+SJp38s49qkoYnkgL+L2ijZB7Ga0Y0mH6e4/B6
ZEMIEhMJQ7zh7NTa2GBM6WM1z3mX+qhgysWatHZHPpxaihkMqWQPQn2/smZOPIic
UQ6i1DZ/EpJGjLZAPJXa3xasH9aSVXMeSbAdEPJVvQ4bwtrWC/XTywcFbN/DpiB/
1mfgLksF0KM4HHtbPSzMjLz3k1bCw8Eg2h9tjn2p7c1R5UhwMla+cHjdrvinTV/9
4ZzesGsXwQZO3aJHKjHqJas98QFAJ2Hf1RfZmKEUYYSvdDdiPqr90HM96JMqMUpO
t9ZGqY47nYFXdaRXdkO58g==
`protect END_PROTECTED
