`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43IKFu7MJ83h9VR774GsOLCy4aff8BaX/Ixqz31NbFY2
nG15xCGBBJSGKMFFYVZC+p3P0ueLfJ1JYGr3zjIaP4UZ6nuIaDL+C91C1LcCjZWj
lgR7Ta7IY5bOOmB9FU/VWr+rxg9EG/0Od6p82ybl87P5ogQO/PCW6UDOFSP0HlHb
FMzwz+BY2V1usO8D8SIePw+hTiL6X++EkxmgiV4wED1F046NNrdiZDSDJdkn9woZ
Ok6d58Cq8yKFSSet4xEQDsGaIBZo5Km2ZeBeGmUc91g=
`protect END_PROTECTED
