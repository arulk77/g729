`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLQMgU9qHFK6mA7i3FY5l8AkbCuYo1bRBNA27nJkyBzU
Xlj1BmRVF2h61FUUcj5+MQjTxIexOBKTb/ivjgyqZYfupL+JlEPacERXU5dSvcRA
l0b/c528WwCPhlx+tBnawmr/uhhk2ib28YszGCHT/lugtQZLvKiRUYfM6k0xSljB
wYVnMoq0/KTFZgW0sM7DRJ0UwRt5roJzrVxDZxrct6IRCAqlWoqp9pqscAK6xcl0
OvIAD+FC5jOiJR+PjacuG8dVvzlgE93QledTjSCETVnG1bJlcbp9RUy/FqGbl7bV
pEdbDahrmSwzZbM6gUIaWec60aY1Z5Qt+g5vU9oJQtCHIelbjwk/CJ7cpYi4vQcZ
wbvCk2/SGlyRegwcM/69Xb/T1fKP+ce/Krvg0clHofsOR5YhzAdmcradXiffIbCG
vBdX63vPxxerP/cQPC1+gfBJ3lD8/arWnTscYkDTZgpf5kFCoQpbrb2SIw59S5hR
F8P3+wLt97idlV89w/ee2qW09yct+C9oH7dpVGw7CzgfqHP/lXnnG0C4IACF5RJ5
`protect END_PROTECTED
