`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3ON6twM0bRyFDJLDX3Tyero7W+HGie3iZxF860Pdb7VAexJSpDR/c6Z2Jrrzsyzk
oery2jM839y32nH1JK5M2NYZ5cXgd1IoffGK8F430vMrzWdtcKi0pJeXDZbBRJ9z
2TNYBCnzkEyylEch4aMNyTtKA53hVgzEgbLKREkWC/1F64kwK9Bf8ZrtYIRrKMGJ
tvzkRli6S4xC4vpD7tCGog==
`protect END_PROTECTED
