`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
K5QREUDOQECbkEI3a7IRd5julGjARiNt9KSc1QXWKEoRwlOSD+CANVVpDHKuuIpe
UUqypOiPSto2V8TN3lUeqAMSIqx5GCmIewee9RVdVVFweYTHNUgwnHdIz26RLgBH
W0c4CjqmmwNya234VU9NWMtrGpT4a0odVcDafCrRmrlYMdrGW+TB9uo4I22Rjpas
clYyp1vXLpcP1remyi0B4elTnZ70apXc5H/cmMGzFKGd2zsub3DluM55s2WS7apR
ftf8bgqYOZ85B5gj4oipFlBZvD/ueI0yjqjkH8Gkefhh1faWyy4UMVd7XhkIm91e
FDwb9l4tsKxsg3HPrQZu2jDUj1CGFD7nSv0eplsXaS5aad15EKIZ9gW5dxq/IJmL
XqS2oByaS2AuSGpZNBYhlP+PHwsHXfNi5kgmSkwk29fUCEczYI5CVSbZgu3ZjPhS
raJB+rYgqtS0FlldwWC0x6eygzYJb2+dYxdqU7C54oHLAmnzFhyfUxLK4i5iv0TP
dHRyStAAb8zBdva/WzNwfQLcLSNe6liL7MxGf4YJHxO3dOSwhbrnxMm6LhP1xCr5
05ktzp2TPZtHKdyo07MSbw==
`protect END_PROTECTED
