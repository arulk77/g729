`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKv6RVhXUhmh1x0dziu9xqjLx8NWogEZEU8ucKbQO53I
lvzq6pz4wRH7hc9+48aRVVCZROWX42KaFQV5Gbxyc+D+m6duts0k5+QeFfh6KLeI
tEMSJY0A4bGkQCBtk6sFxNg3r0sYfpM3FYONnjO+WoStIOCbceGIfpXwIVrcmDPp
VhO9c/fj2Wd3kXufdBw4hg==
`protect END_PROTECTED
