`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
NxRPnlBxph6QYM2NcORKsmLTsZ/G2yI5vxkSY70LX2qHDNBET6V0AIbNBfzx4DK/
Wv2qjtnL2L4i6jaycqFIVZHiQLa32ZFgfRAgZNN0Ktlr66jOzHZ+eHyNsdPJAPB9
WBN1ySa6IgZ6QeyS7ZtoYOpamTPMxd2PTF/2KT6GWej1k6BVSHLSx/DsimRqLXmh
0jPbFfVU95qbEgEAFjcYQsbH4m5K+owzVxZ5JXle2/I=
`protect END_PROTECTED
