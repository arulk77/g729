`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKR3ol+yIyQJgp9kdkqgAlj3hE1FaqeyFJgS37RIAdym
HEearP2VwrSOh+ViNndb6Cb+yv+F5b/idWP++EXwAUMuQhyMpMDxMNIrkI707jRv
+t6viitosD9sBI+A7qNdFN8HmRM67Q8MTlLtFd5XN/8m2MflDMkrxuch7rQe2NVb
n56iwDNTK70jIKfvkrBVJw==
`protect END_PROTECTED
