`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJS1za5UNbNv7+LVSgJ3Fk8Nnnjy2oMylyJsNM9F5eMF
NMVtn0i3s3S120aIhjn/zX3YCP2BJYe23+k/GaogAAglq4rsPc8BQpZWCVILiqI/
Zg46mGemxhbC3QUf9L5wuefQk2DCR0YByWg5TH6ZATWEQlGB/ApcFvX/A38A8D60
pRdoubK+cHrVRETutziB/Ddb34dQIPHcOwiDoO7ji63ftbCOjPz5+BOdS/nF+xtZ
w8Y3K7hv90yWwxANRqL9slGb+vbjw6OU9P1lJaakup/7WduCiIWMa53G5Z7XkoEW
XXgbwanRqXC1SANhGn9RcQ==
`protect END_PROTECTED
