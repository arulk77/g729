`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMZZ3TSVDKy7d/TUDLo8RCyCNpFGfW5wk2eDzh6NnnMc
PxgKCTrlGd89hi87OTJbugpHQmX47dssMQN2dp1Zi3qAcOj51rKSBmFCGsC6RhpF
po553yhQnAPjQTydcLkmy0LO5qAgP9desSM5/t7NA6TvFuIlRDpRfGQtJgNx6w1e
Cg2Dvct4kKLqLik73+BqJg==
`protect END_PROTECTED
