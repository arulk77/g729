`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
if7OW3neLerq5QTb0GME93UThSnEFAh3/1c1OJv+xiDmL9drOhTghUA+9tIKYpnw
XjiJOdAxFuU0sdbdFn2ALlB47zev716wEpA1tCRmesADSUppKxqGMnm6AARUhMgw
v91HqvFLgDXIudvOoAJsF2sKpT0Er0zhH3YE6wLwMVkm8+rasFLDrW5T4btOCYIG
8V2j9UB51ty1Q2sG+0ZaayVj2sfkI2OPEcC+uA6YN+677RHONH2cMHcuGCNVCg5N
06U1YMp12OELtKZhJefs3vxMk3NK98iOU7dM3EfGqTqPW4tOofCO/lMqdRMJnEk+
`protect END_PROTECTED
