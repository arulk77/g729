`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Flus04vghmlYdT8S/trBMsfaMJatwXIvm5iJQheiqx6CuLFQgxs8CrgPzwBt6A6L
QpyCvHvE4K6uTC3Zgga7P6j786CTmOglR9x401LPIXRmrFAciR0JM/VvQf6lLR+d
pVFf7sBfNqzfbgHbX5auYPEKHimTzm/GumLrbpxNuatavsOPt9Y0P2KK0WqpQR0p
VWcPmgW3Cpt1YtMLq6yN13CteKhBZN57kM2HbwIAWMp2qjfIQnK4Fdm60t8N/U//
ktmUmzuawZw0dYv+hdTftan1wsJUZVAx0KS6pp+EQAY+FLpjKrQVva9dYYeQGwW9
vdwRD+wFWhl0Z9cnQVA6PDc+3AQbk48Ubgb1jgIrsziED+hL3YR0rL7Cnaxj0Lsc
RdTX3ALdI3CgDQmtmjM5ybwqXyQWr4SvmnP3KSm7OC8Y48/gMHRFJszzFysD2l8U
hRkVz2iWQmCN07BIUFRMrkKZd7ujK+IJ+MjugYa+0Af5w62hfL1bSsHlyoV7UWIr
F0zkDZfZmX3le7pURitxKvUcxRGS14MQjLslC5eZDNDyJOi2/6ccqrAvKy2hKc6/
Ehj2cAG3PAlsmh25i4ox40mK3wgNZIwjF4ZZIHlq0O9zUiQffazDfQINcj+/gSOO
DAhxJ28Cx88JX6oL4/Tic0bfCx4RPHRfyAvudPsNtKxljSTNIWOm20z1y9ijp9Vn
`protect END_PROTECTED
