`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/+/YWjgCCq5EsWiziAYzzUrl3Ekhq3v6zknIL2ZoAs1
9VNuBScfeoJfbDKYjoz2PWC/mlsiA9QeXldlGVwm29GLqWNzSpCJCjhIX3exAbrL
0RutpV6tIHBMEeegffa4RvZt03frUjVbmPRDz848/0AQ6eaf8QVcWiRPuU721bPz
r/TDT2cMKzuYBW9XL1C9EvJ1K6yZ+C2YeLHF2HddGpREbLJF8hWGl3GBe3FW6yJG
CXj517m6cFyTO+WznH82y8w0Ws7F0XSSe3ZWsWIUwZn65gZCwZZX2pKFTQAz9Qin
dbKmo9RKl+15gJ+9hxLyHA==
`protect END_PROTECTED
