`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJpjsHUBs90JPN3a9vfCBDL4EWgE1MkpmqFFC/EAQxIc
s2kXrEK6Jjy6KzWraJJ/Rkby9fv6y7DE/22d0vPItEdIzttzM5/TzLQTV2do/JFc
ZUE1a6mY4kZo3JuZHfGd0t08s+eBHSrSdfwVFCBOrLTMT3AhXjgwBiMW+R2pU2rH
jwT5mh4VdTxtOP005pYVOntK4yC+3U+qEO/7/SgV/Yh0rFNN2jwEhJfLKQ5Lg48M
+LAh+igT1p2TmWOSSYmW3rrIpnKbErHAEFfzSmpv1pCfDrXeujv3LTGaJhxNrWYo
2+t7QvcQmXrPHLkCtaFbsyECm5ogsQwJXHk9nblow/Y8DyqiEJtxZef7oGqn8+pv
kn31M3Ugj+UInq9HqcpbQsACv4RC7vjZCbUMPnJCGIliQIGLy1cKCJITGaWPJMvq
4jDzXijKQkUhPX9ZHV3Dni12liwTxENLb3wi1fAqs7ig9sGV4O37ImZhEjgGZfjX
`protect END_PROTECTED
