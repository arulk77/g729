`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveC92HytrU/l7trdMYr80b1OJvD+E12dSnZGfJnOCynxy
b4qG+enQ3aC2asH7w9JemmUSwqiIKRymMGXUhJwT4BeHC97GBEQtuFgbRE9ofU0M
L9hjh4Klc44Krg7K7Hnr56kNsVr8kBCyYOfz/rOEW9dZQStl/24jBGLeNQtjJr7B
8KFzWArWhIF9etPsd2DydB2n0f8pq+9rxvoS/WoKMSl75h91Nhls38qdDS11dXIM
`protect END_PROTECTED
