`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCPVAEV9PSkIwztO7Kjl4mHQNY4hHmotyhJ30yl/bNpX
Au3FU3YsL6gC/iVIVciZbwyZG+Ro3HJbDW83QEpTDrhG7jxDEQE70x0Ix1uTssHR
MCOmnn/URfYWr/1Mo2Oi7nIBAyJ+mcv4OR99IHl0LLAZAltya2vFw9rPzcBrkkGG
EQ0NefowxXdvJQtwaUCc66maSqGxtKHzgP12pElNzQOUbKeU52ATAZw1rPa6977K
Q6mp5F+k0U+XwnaEu8K67y8XsGWrFinNr4MiLUQFcxX70K4LrGPbHZiK50LBsoCh
mKyvbW14zye85XurPtQZmChcibOAxuPDhyphpDj4sLyxs1h2zzfDLLKPXT2BRNjR
9rtEdJcsL7omq70jxnXqB16JVz0DoM+wZcCH8mJMdj232HvGb3EJTbDzl13gjq8S
nyTmjsls6XSyCrfgwcjwaWwcSO79T5pPzvARwEG/qPwXuAZalQdXV/lPkDZq8mg3
Y9XGtJ7vY2pQgB3Gtg5AbaTlyFc5nwVu1YBvhwaO6ax9BZaKdr/HX/NxIzRFAip5
`protect END_PROTECTED
