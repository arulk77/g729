`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
//apt8M5nAr9YM4Z9a1QOUpvWVyR+XDA+9CA81HzSj0VxQ9zAxeXWdtlgssdpDDf
i9smyRNDsBoiE4xe7P2Vw9svqz0j9rUxDOBDlUnavBrRD00qAAbjILuVgRCjem/o
bFjgxshyd1ixOELJpvwJqM0vL7MsVHva8vMXboEQx7aP7LYGxBuGI+1ziOI92fQ4
dz3/Q4HeCokJDH+L26Wc7SCAn5zyYiFtZZRz4OXC4nanSQWlNIxLr6OwQubJG1v/
KuYgJS4OtSbOcjaqvgUeng6h1LnHCvg52MpA/uVJHc0=
`protect END_PROTECTED
