`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42PXmbUh5qWmsLl/9tlKqiJnN15FRJfTgcO5hacdlqK/
ndhn/2B0hx54+7gfNes27mBuNwiWAs3jTdHPmznIcmesUrdeyseIxXAJ0Mht3M94
fn2/YeKxcg8D+XTJntuCxlM9P6LKirYKtTEtISNWUDnK/UEtFHyrGWVjIB/k+Agh
FF0tK9/PL9zx+9FpL+0gp0r4h8ieVLersdeT2rorWJkrCVsyXp33eGn+3h54h/Af
hB1rlGehcgwZj0udGwZ5LXLornkePQ9daAhwno6GFwK4IpeiWBUaUssvmo3ThPrj
ggD05Mmmbdx5q8g2lDMvNA==
`protect END_PROTECTED
