`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JUxPzCvDaYvq0+PWe8TZvU1kCj59DkE4RnUv/tnwNCssFqTnRpiktrToo4a/1Wxp
RL5w6eX9luPui9HAR02Zos74iwQVV1HXz6nxhqFq2ea0lxHxiP8hmIfIdJ6YOK+G
4dYNNmCxZfwkPP9ThCRS6fvCOYCT+E6eJRAQ2J3FYoxqVTwA7yowoHBiGxnO4XRL
cAET+MVC8z6tTLAUoiNDdnGhDc8mlqX6oNL1GkheeHatv8wy9NFc2+Mb7q0toxQF
2Q4ZMUDFSDRPhZeWMCtk19tgHfyfPPUWVbeZwHS1erU=
`protect END_PROTECTED
