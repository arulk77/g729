`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFDFZx2/KES0o4vkfocuiY8Tlcu98CGounk7SlCc34vx
3ct5/CnxCtx8WSN3gkk6KKq0r8v2tebvDLnCb80FpCnT7A6ajRuBwgteJs1JKD9b
71zNycCkCzBRIh+gmn5V5N+W1//KHzG4A6aqPjJIiG0Qxf/UvUG9LCiKAZvVb/GZ
wB+D+S47UyNq8WrPERp9ADxQNotc1AOgjkhSm/eDJbvb8DAe531TASfGLzBoMra5
OLMvKJ31vb+hYswI+SZp0hzFs/k9m+H/aBcRs6+f/57JKW53kfX2D4EEM12Nrl5F
aWJT1PfM4CP+8/Vxv5dZHGvOFpWL763NkQrrIdlYfYasy9lSY1lN0t6bA/eUgkM9
Kx5TN7HyCw7xs1DKPBrXTzzvIdVivVaRKLxb6BhO+YVuqIZ7oE+ITznSKs69NToJ
xkwB1q93JlgWa6jwlVk9AcEo/JqAGt/0LAghrOaGYyj6a4IyrGRf0dEWe48NgAdX
Tkul5SnAIxtB2zzsdYZq2h6WQjTVWMvB4T//93v3JSzfikxDjGaK7ioIAFmlp8AX
xacqBkT6pVmcMaJqHvwJMVlLG8IMCCcZpXGIftcO1vUYydjjEkRqRp3KGWYcKv//
rs+XG8mo27lJlPkLdNQMa7gXGj9GihR0RNYZoL2aX5Pu3XPSL9AgZ5yu4T7++jD5
oZwpP0RI8JyCj56pyK0GYb7SeBkQj6TZ7C+FZaK+fvL/o0SDk6DdhFIqiWo3WjDZ
aCXhbXPe469jsAs5UYUKYOfl2V++rGO/MwE+1Vl6zhPyuOIZWnKqp1W2/IWYVGzd
UgBvw+a954psvtrVMg0Woap+Dogen0xODm3vLNADrqd9/P0pL9oWxPw2Csl1+QIQ
Gt8aYfFmXZA46jo05wiKlfOb2qpcKdo/BurO+JZ3oK+q2kcTo26hY21gdDm2nNzA
Dr92aHdXq+370DOhbmld7jd4Q34sjDjtVrO+3QyJbrC4hjwBP5aGjm1G+cmLOv1P
ppOojPvuBh9GqMIDDjNIkhrYFaQhLAIgoPEzbNhyNNQnQA8G6+5GndTk2heHP5N0
DEK1r0HqZWEA71HcGsiuYlk/rEpHjQzIT/alruD1bxvx91c+I45zuxDfOzoD7IxK
zu0HwsNypdLONUmRIzU4eEk1VbNsSKOH9nqIwfOuVqNWiuhaDIt7BYQcGRF+xRE1
bmjRSjXhcrrWT6hl477yYvPG6CLvt8osRqES6mZKpbLbYK2GPieaYzfbrShJuYyz
suqa5nma1oyuSjp7xRQz9C/qAESO6M5WBNSAtw8dI/NREiiH8j42McibR5Z3bGSL
iPXCR0VzMRVSrPlIKyjbSpk0Ln2LjkhbimdnHM/RTY8sDqDH7d+CjL5acl2PWbjy
XhrXZv9ujgyG5bneA6hh4pa55jeIloITagcKWJEeqFtfVcX8hXHByBGShX+0dVuk
nMuf13ghJhjCIJqSvGw5m2CnEmPdTn2oII9H6SvAhc1piwVG/EH5snmziY0aq0QF
jLITxS/zorSoVh3AeZ/yJECTiLIllX04VvjlLbr6UGdVx7NyYcZnJrJ+fwb3lknt
iiPp3wNIZwiezDvpbnYm3UuolPgzszFaKhiTrkxkRgP8YqRmf5y/8/RV8K2xfylx
PyLp2MSO3vTFUDkiGxZt82qTcxtJik4LAUOzfdPakA1IZVj9hkwkh307vNTOARbb
x6TbNNaeYV8hUmFJfz08Mhagl8eclDZ0fUKGUbCvHNsiYuY9BW10Vwy4UYygUGCg
qncvzcNq+pPJrI3tkCaofCbTClHzu7KWzRjEkMzBYrpN99o5P7rRRUIAkmfKTsb6
X83NNw2p63SvRTIOo2Miy1CLAQbr4HA0JyeNP/j2KuoszFYahPrzvJMRrsK1QUgk
e65IYJLmrxeo6W3cpPkFRpzvBynF0qHq/6Hp5YhkKu2kYlPAa6nW9R3AEnlgR2KN
PICQ8HoL6GWuyvtYfreEh1SrW7jZhlokgVEuwaJQOO7Lw69PBhn4y2yVcbip+F+z
iYoaQg0oVo44/Zcvbu8Tc793GPT+p99y98fFVXJ8BtfrZiEVZvVAMmAK+16H+z4B
1MkakD5bWDTKYWM47eYPQj7I1ouve09jr2xDNSL2BEvpl5G0FqKqluodkFZGcyh+
K0gcF9Tk+B+WadONqdPxssi9Zf3x+8RDH6PPleq5X0O1XGZMVa5dx1SHVQJWEvw0
QfqxmYtbCGDATNmrs2YZoyXTCQRmKi/eGA8kg9Be434jefrFZBMcWej23m+5bNmx
zOXx+TEAKwLLHjhkZVWjPFGShajeLkE3V2QlaCMgMy0L5KiTpYsngon3ajC7XUH5
RNhl+93iMRF2+7kYz9ibs0RsxvMrAPksqFmtVhGRFaUCPaTBA1WIAhtuzKICxg01
ofgdAOONub8kkOHeypnuFfgKrUCD3XkTahs8zFT+hGe7NZFjRRC0Agoq+5K07I07
OFdnmBv6gSntFlijnLtueIY2j2eo9n9xamhmvxQwv0+tPEYW5UY+HksP0CfaRFRK
TWGkCMi9KMbcUo/YDgztQCNym8M2NVF2OttlL3a62cOuycJjxD5MBM4l4a35TAAk
nZUq8m0i98RDpXKfVS15NQLheUh/xaN7Mw9iJDWzh076Zm0Iwmrz5aakRmwDdwJC
YHgwxpk40YDQMFEGg7UwKR2TdRTw0e8Rnilii+IxoPxoB7qOXnCcRByiShOkonCx
3J/gsrlPdacsppqCrSh8e8Mm23xRSZbDFRIScIMpdw5uEoEZSTJ9CX8ePEyP8moe
4lp0P+YDPgw+VUuukIwfcqxqxzvpNcLwMQCSpHji5LFDs1WjRNeJDPz1P83YC9Ba
PtbZcmgW231semO0Dmw89fEGMAdvdGmcsLDzEox+pBn0cWej4JSjL7Ky/uqnlSC9
ANp37/LxrTpHLgI6ejbyPTugko9VjxmFeI+aFyJP68XuvSF+9/4lxXJLvUnQWrt0
KRF3uJnrRhmv1n/AixdK/7tamTRmwZCitl+cAwGQj2BalnFMkpYPEMt0iFZwPzRy
l1GKomXRd/Iy/oWJONdrFxqr/EDrZyj9jrd2Nvo683V+jzpNNx/AGv14cVgTkvA8
4t9OaqkeSJ1xJQ4RnFTLTlzlwUsf0vr/hk1J/vHTNAQ0xu0+KQp3UCZF1rNZg7Jg
Ft+wmiRAQsLMF1Zir7K9XOmySp0l4E/Xm/Lp4SM/8w8O/zxPENXZ5jVCMQMnLO9Q
aVVSVU5odgs56UTRw0mp592/S2lHB9Nw7AmkjrD2gGTcGSYXhkcWwrG8YQ1j34sT
4aEP6AeBzB8tO2v/cgDgW6zLpmhXcQ5SFZIVQYKrOTAF4LiyXncXpXvU1xlFXw5I
P1VHKJZX/IAMs7iiERId+I/uTDzzQma8DLNE5STWZW6pM9VFoOpeGbh+5q2uVCx0
T7lvcf7HE1DcHqnzAuD2cUYaGRcu/X/ez5T3DzRyM/jKWL8aMx35R/VKtDlqL43Q
o8IIzlxFKgdjjcp65MUNiK80X+1p2Ubkhgybw3xf0cwcruG5FgGTCQSX0PZdvde1
cT9xEfqsLzqkoXN6NZ8FR1fqGAL8MVUxtpcPgk/j8HtDmqfFmn5r70oAFl6IpCaM
OS5QMthe6ugtS+1Nbzj/fwD+gLzW26KINrw5CiJcnqRGuWbCNsceFyBhs6ceepqM
yv8Dt8bZN0v9aeCy7k3vO5Le/NII2eanRneyCeQ0N8Hn32QeMyh2ZaSdRI6g0EIn
uFf/+F8Fg4VV9piY+kSyWEI5f58XPjIZIH6IfUJpBulWgo4yPOrxrPnkk6TGRuHh
mGWTPi6m4L/ryDBeJZPaBBjwuYoCQzgMTXQf3oRzWqI5h4QQxEMNZBEf/Iv2oJwm
TBvsMdb6D6+z2u2BPnRSzvFzh0EJORdbYT2dkfhwtFy9mEp+ke0J1omgTHxcn5AY
Oy19bNIunmZadelERDzM410hjCnXIQD05HlXscTwm6dk4BSA2D/FmQJ4DQQP8Z2N
TtrrLC/rS9zUzjh5t5QJlhgGLURcls2Qw9UEI4uVMTMN4nBt6JOpOG3HdpHsqd2g
qpphTdJRqI4Dfbr+n//1u8+vGvxqrS8s/EysNoJHDOjlXPBKb6eNbcsrrDdatBiQ
6UjknKvrYCOrjI27Z7uV3tudO5EK+UbFBsZW1tyH/QUtx+43hYt4QjtzajVHYDIP
K5ieYeu8nsFGA4JP0w7E108bTKu9L+BlIb2a+6dg2CmCaAuI+NJTym7YFdbR0MLh
MSGyVI2bUcj6BfyytLGtpgQkVh7TovKq45BDwjW9Ph0KvRt8gDkxBi/ZazwYk2oC
iAENT5jqXlm8lkR1/U3UZQfBmyMMwn/WyUk3GvlL7a1wy9Yh4eWgG2m67kwcziIe
fwD/IEUJfAsJIoVw/gSMRXwPnHZQM+Nguiq9sS8C7QJygz4xbCKINU5p2V1yr+Qi
OU5Hg8WK57iJzgdS/3CdK930h+KFHX9Ha7K5GcuGjJMxcA/lpuKvTcKrbV7JvDDI
q0ndpfPNOM5VW4UWyCG+vlXV3hHbwtCCQRtVFbvLcMb2yyXjAYLi0ZojL0OCi8MM
ZEQ/YumXAIIcCNyqAXqpozfZmPGGQfbhmsW1o0LXC5LeqVDYm9xeL0VVjpxpvHaR
UeczKa8MDzKlkRuYXM4Ug/jqyvWJgSFtJvQCJwe5jWqW317KdXQym98MUcq4mzgI
j1zuqO7qf22jhUyVCG7hcqNNxJLOGRBFwQe1mBDli6YP5//c6OW/U7NNSg4TAt0F
luQpqZWcDQp42/f1++FQ04DBQH6nGSQUEbAmb2zF2igrakj4/j+0mOZvSfpOXQhz
uFYQzga4zy+XZgQniD8ro86Grp9WjdJK2M7PecMCp7Ib3jz0GO1DxHIfNYvogzaO
hnc796rW5Yayj+W0d/5HzO4PFLqOC+KCMS9HuGxlzpXtnqsrR7XrcsZr5jmJOosG
ebmsuxTfKz5X0Ipj31NEd95UD0rsX/OP/8f3Z9g24dFQi1RXvajU7xJlks/PSHUz
+QPLX00zpz/LYJHn3xj/9W4i5dgGSFJqmKZlVh/137w+8jxwUjmw/RvImiyVDn5H
/VioJGIY0XJmwIRmo8x3oqSFpA7Q/dvjJSqbWv3ugcjnEJGL2cwC6HwEWOJPCqKx
Wh2HbPPSKk2b9oSM51JE6MkIKlyaNkNEkuocYg/xBuwC5EHqLru0T32g31603GvV
rrR4LD11ZKS3Wg3xmMdvKA==
`protect END_PROTECTED
