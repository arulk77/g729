`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46DQndaCiPPPyouyxsoR/yxh0dkWz7PkR2R7uGeacpd0
GIfcKSZWc5hgnYHW8tTIdkM1U4Qf2zk0r6F1j49gnpD5Uu8Iu1x65/BH+26Sc7cR
QuMUhRlOiM6Nx0dCXNO7WpUBs+PmN0TKP/C9OMgaU1c=
`protect END_PROTECTED
