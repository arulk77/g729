`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOBkducb3XKWXrWgCu5EFfdUQ8Pp+IwLDtLo19CwQs7x
/L8+d76kQ0JitH2DJLkVtS/S1RLFMy7EF/ZDJI/yH6voxEvI9O+AhaWPBzyxCtlE
d0js4C8j/+KHQ1GKG7BFwTGzF4OHLO+Rc71vf5A0lL9V06tXtmwNswcvl/KAaesY
QzIwTHyMfV3tpabFfQyYClozhVo5S+nenXXZSGAhZfW4Cb0I/bYilZDWxzvsGqIZ
AZuQYNbeZJaaotJESpwtBV4AheXJkdTXWxxEe+MDSsMi+X5AOpbLXOagblKJnjqT
13K7l9Nd3WDuH72AFDD7cuO3wAEpfjfJiYvzniGTaB6beod+24I8+Qk5FfwGTIjL
TTYEJLCUkPYPjC8aALbgOBflTQZ6tC+16RYdg/dOvngI4XiiQYeWXZs0etQDyw8h
9GkBSgjQHSHAkSYlddHKEaoUlwc8i+pshXtSotifSIozN5cajNfFEi9F6Am+HCZy
vWYf4Cfom98+qlLeAPEjA7WgD4itjPzbzeFZzyF8PRhTt4sXqtiVR2I8cmqMtSUK
`protect END_PROTECTED
