`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
S9ULEjJpr60uqp5txzyR4G5116Wm1VdLYUT5GdZUVJm0Qlbuc8bfKYsyHWmIV/p6
8IQNaU2C4MtwE+vFhQyfj3OUfHDQG4oeLMcOL5SS/sx3086wQtXnM7lKv7ycqG9O
bBUG6SPh4R7bPTejQDaQ2v2HHyVqmxkF8MgP065uM58=
`protect END_PROTECTED
