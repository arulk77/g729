`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xYtnrhP8Xb/wwNTHGIU5GwOIeQhez8y3eC+brJvxEcx
6KkeIvGj9LmLdbSZpUuQuEYxFscKs46TVo4fiqYHDYKNUjJDHa/M5hTLRKYf5UDB
7Pyk4qJ8bCeHMnf65Hx5qCbBKH+BrqVEL9JNbSB5zmVIYXU64GlKvYsM0XuvRPeN
sKveMOB/hEG5FrxvGqvqeKJgT4AXUJhe7v5lhycLWLKnicsSxPTlwc6IMhUol1sH
zW4IWmsn/tnSEu41ntxgZIjKs6DgtXplPIfnLJRtfxN/vaAO/JGq153EcaAHD8mW
xgNUxHVaKmhvjPrCDEL2SNCv9aLbFenzDwDfy+z96jk23U1OuuKp04wcTknfUajH
zXKL7ReyNAo7frN/sY+O8NrM4FqLzVWj7T/tPpw8vb+hwDaOJ9SStGzJPs+tJTYP
kjxGF8IxE+vPgZ5rgltNsg==
`protect END_PROTECTED
