`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOuBhGMuQ2xJhJUb5OreDbi0VCECPz/C+kyUIOMWO8/+
QjZxuPeZiF3lXQCZD6R6Y2VGNbkWeBJLRG7oo1FYlJUImr7QZYoFACVQAP6dRgNW
3E1+hYyk+ZkivKXwh8zFTKTQ1ZWYVJVPfN1uGdJDyPpByQOLIEp+qgfKT3GRtval
E8EotJTVdbP+t+BNee7jn3Xp5gWHN0CPRw50vF8DPEQPXhD8FbEehDV8Zdmt2Pa2
k4CRRd9+ArflFENe5wm4FHo1i9C1aj9a7KaZ5e12DGjI1nQabU6h58kfe8fNh/FD
oq9NX9koHvB/wQ71kzBwurOIZUsDDsQqhmMYqgSWT2lUoHaPrvFkvNhSS6xFaZhZ
8SxFAquL8wTvMVoyU9ThloxAmwDwRqZSg5qiKB67LS3fHnAoNI3N2pvHk9mRBmzr
XBbeKGW1KR9gjZ1nW/YCYzKVlRusTkF1U7R+1zW6IpKoxFKuizhEQZpMqJmm4BWJ
hFdg0VypJhyNCZvenInaNoi0ta2Vyou/Yj40f8Mi4ZCS28knyNV8BhL2TTZFymdJ
Vh3r/lvFu/hN1jMhLGu26YRX/iyJxizbVnZB6tbXPPakmTybwgmnkkNmA3vi6woc
+dGvT676OmKjODrG8EuiFc/MPl7p7d0YB7hm9SeLxYhgSG4OQ+Nb8wpzNSh1WBu4
O7LmFIwZE668M16mYsGW0bQzhujDs4J98xrrgD/GMUC6o/ZlGO1P57QKYX/NGbOc
mBT5PaWQ2muM7i03943j2+F/TV+WCJ1lGdh4thqeK7iVcODjvtnh4Y32YGdf46kj
s45Mh/rHMWJaA12dfTfNaHLgaSntJIn7e1IO+QDMf9fIsPDnfgT5wkRdLdstZzbg
d7433w2DL20xsqpLLWlle5SzUZPlZqGTg8YteMhSLLY2AL5JvUs3zC/Zg+asgc3M
ELl2EYjjA5bkSkTXwk0MYRTpv6v3hJ+5hT8pz4+i6yaYmQxiHGZTgpgBVEkBrBTd
BtZBv0DJooZzNuRDh4zFQfnKAj9MpHcrBL6euC7HWLPEkDOZhd+7ATOLjLnz2xip
RP2Iw4foZ1a06uXOnCgfv/+WDrfbUmYM8bgKzweZXJV6b5Bc3o+U7mkeKtLsJZug
irFTTeIsOFNTIbpwOzF6VKD9GoL2O69GxQazl0j0vshtZhxdVy8F3McgNr2mAmhc
1c9RB4YEXMIVl/TLrOGalh0u47+VOHHcHcKFOLVOW02M6hbpI+adj3ZdBvJxpVY2
BHo3fvRpzqgOLvXPhY4zw6Um1uIDxRezNG+Cm4yeL3RHP9lNnRNME8iabfI4Xfk0
E7wQA5AxcwvgEMQahCaGdE0CGvGi1rh4QKc0PUqtqIgdNdETNdcRE1mdIdNoR/+e
TWXkWmkJ50QJEIISASz2tB2vuzQHlzzlxkyK9WJ4jP26MRfabLJna8SdJaMchXqb
LR0wMuY8ZMyZFUt1et6sdhD7QySvg6E8A57DFkcAJZvkzlB9KN7WBg8M/EUXCXnE
RGJJNPECm4qLt+kQiTPoZrfxKmbzaa8I1eMuY+AXi2RbjTuws4t8/fxkuaK1vz4g
eHDsePVXRXeScN35iiA8LKUt9tqf1jq304yDsQefiYQn6Hcv5CD+0N2qTgcJkRJy
pPy4IkbZbwVxBrznUob6XJKwJhb5MzAGxKubq0qg9bt3XbQhEVNBnPm7W0VTPQMQ
LqJSkZUnIrBObfdUesAy5hm2FDP3Z5Z77PSbGvUPA7LSRxg5IO04em47FHG/Eq4v
tl6/z8+ngHoscwgOzPxqSbpHrINEiLtu2zJl11H43pciQw1rFt2PDmIzkYf1cCjm
hctzRgm7yvETJj2G+qFoxiCT07Rvz21Ztq8v10nfo70wLjdGXTgv+FAK83olh65w
3Rn2C0hO4MHQaPObtglNBtLux0HqzL1+GK/WWZ8AfhM7ODYpf9l4OsoOAefuus9/
UWqiP2ICVUKOIlgS7xqIEHy9aoFT9ZBuyvLVyfMAKzF674WaGaBpMyC9cK+6b6Il
bUbbjiig6J44JGAlWrMOXdFkxf9QzpNa6ShnWN1Qcd65fgS0KPhihxD95j9gUanQ
6SPohWTaYavnehvK2u+q0TLxnThO+BsyM0yH8WADbc/Rmk0w0zMNDjwGjCa3LqjZ
bpeJ19tLbwL2cGyXtVXobOqhA1+6h48kU7/lhp6zOV2cLgZVEczllQRNc84IJsZ5
Zj7SIq9Sz0mYDexuCxSWBVWzBGNhxKBCW/PZH/J7ZUOaYNPfbGXRkRklfmMO7VMC
0sJbmZPk+IO5kaKRG/wU5aBIdfg541KK2eEOMYjba4pz+XU53l4B7+3KBbh/DGzj
7L5AbG2lR89AgSJ8cVQ44N9GIsCJqfgw4ma3ioiQeViI3aEaEEYxS3zs2n/JkKd/
GdkHG9HeUPPnOOqNsmuF6h/Y509zPShl4oZzB1I4LnbiQL0xpCSG/UCrYUGrKYNg
XGzSQwPytUT//yvyErxQp8ctz9s/gIYaFS6cBGldouU8jW6cg4bbGr1JeIGsXtyZ
`protect END_PROTECTED
