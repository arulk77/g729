`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
0PHRBXJkLjFFwCmnhGEJZAtNF6+VLCh+XvADpuGPwez7FVLW7fpckyZM3z2u9oll
KWZbdUlIk5kcG1W7J7x12JzW4cPNLbcM4amLe1JF2P0WoXO+DSUt/fLaQkT3TfkC
We8jTrhEgGlQ/4ZSmwIlyF8Wji0nFSuwlLUjUcRcQmj6S/PL499mLuOojdfLphV9
iFbkvAWBlWm/tsy0jNP2x1Ba3wxgZoERhYXjd9fRK4X3pNQl0CzOa5kZb7ey995w
ZgFWGGnU3l+46RhCuCcKf2Rmfb3DFm4O7kz4n2iIchCCeWnQKF3ddSh41Zpk/jkB
9yhmcaSgCFSsN2Dnk/Si94mv5uNMIAiX7249Y6jtdkPLNaJqtoDgCfRq/1Ph7fiF
KBr7et/JWApM8cls2eQaWJeQDBbs4sdPd/Tb5mVK07avn5H2o8kiJQ20tcbxbr1x
H2kmX65eddr/mo0cRAMqpRJ/wOr/hX5jWyt9MDbMDx2+/KkH7wt3ClykHPoo+Arx
eQhtBoT96kZ/MuS4FiXUt05ooYPYOYS7I496dHq2Kq7rdi80uqKLtXr353wSCS12
I7CTJ+Nc9+M5j1AiAZ7RBuTL2VncRnQDXqU4D+gN18idE6cse0vpXa2mAcUnZxq2
Sb6LUdwizeeZiICQ1oipFf5XsnIxqng4guCwLQLK1YhgpwXbJsK51Soi+UguD3se
sj8HFEgf95/MjKx7MzW6q+sfwFmwmyOM4TLa5xmzLgE=
`protect END_PROTECTED
