`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48WHy06nWjtiQt3BcOroDb5piIsBFHlr5e0/KqJwhZu5
m2ABibL2nGQWeKF3tf5F+rb6R4eHYxNDh5TeWON8Ll0aGr1eI99nIbf7GXs4vy2C
VnZtLFPEYE2Fc7EKyqVfDAbUMXCpoPWf/I3mxQbJzhUv/WM9kPRiamhOPwA6VWS9
SZFK0+njW+B4PIUbumTPRmYeFuj76lKNl017D67S0bq53SIa9dp9ptn01cebLo+W
aBdp9dcUZt2FRryxgmNkld54zOPRkL06FW/cSAxQVOI4tLvAhr8LHAypPxNbnpQS
D4AlmGmvOvhGeBOZ6085aphBM+xUMUwbIzdbOxMH6mZFkAw9yCl+ckW5ELfRZ1ee
ZDrA61yP6kQoxIIWjbKKvQ==
`protect END_PROTECTED
