`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
SzbiNJ6dJ7Xx7gq2EgC60VuiycEqoOROz4hf+zi1lCxrPIFHvZgk4Bc/r7mDkNk0
z8pwXletHBfOW+iUVFAJpvrxAty1Wuc8CiGfAU77IXQBRESEVXDN/Ilo4LNAeV6R
iTfa/Fecg23dMVMZJkMMzACNZp0zURtM2Qfr9MKOO9m/UoK1Ij1m1UTzk3eF90ji
l5071CoMCyvqKpObgeOyZ8xOtqtDUVEeHTJDpl3e8bjipUQnDIoh65t4XDRBZFng
NIIE9Wd33sZSQZ6xgNtTD0HxknoLW2jln575UG+y8zQnIXkw7qudi+/rXqCS6g5s
PEYC1RWbWX+3ci6fEHF/PQX6uNXcievbpVhdaKW6hCKxlxB1FUeRGECZvxFTF/l+
gf8XjQDbsJ49Z+jSpU336v3aOjXQ+fc4SHN/Anvz8NmeRJ6IkXGFiirw4hR9rzoD
I5Z+yBLO8HTYkxwgIfrBvrRea3F8D2fvD3pQ07yS50VDU8w7Te/W0xvLbHOMUNZg
yP6tZ+zvDoRLInjG4CIKaFe5E4toaBW1AOPEFMUQC1q8LNwKVKO5J1vKLBXSrVzR
FH5Gm3r6x4u0sQEJgoxDS7PwuxtOe3i+oR3CRZWN7QP0ahWZ579k9/MTJ4nBGAvV
AH98JFLjL30GCfLsMue72LvUKkL6rBhyxmVrq0MqPqbhFa1nu69CU8Y0NQbcmJcL
AKWldmGBruF58H+U3P+McJXAtITtyQUdZ07eXVgEjcXQ2qs85Hq7jd0Q3F5syZXf
2q+y8k+pHk/ORBeob9d0IC+xbuyYITwYL8feTcGKP/Kg6cd4cO36x5EI36EPHEuF
EU7tIPRqLdYNj0sZG29vGMBjbTphicF2959n1wklC1Lwz5Jlcy9Wg7ZwqxYary8S
smZn+xkcMnOgEvwd1V4iibkwbOipB8O8TMLND1782xgs8N8qVrBck9IeRpJAXKT+
ixhGAOWOcbckV58XRB0wx2jz5CqWzI/G9/OH1qhyBLReYvhaQHVvt7qEXtTTkGTu
FJ+uDWtftxM1YLT++3ehLpHJ/KBW3V0rx2xXMcdS0UcvdTrfvI14/YO6Sx/EWpJG
+U8+WNmbopf+leZNCC3btg==
`protect END_PROTECTED
