`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45y8q2FHkFZdSykDLISl/vJW4fumPlUqB2KbFc5dzFGA
cQBoU6TF4pfMG6osFISN8Zza1uYVKtrB2dXwydGmsa3ASe27FAPVza/38xgfH1K1
4f5w0yp6cYHE3mYH/LosQ847LPGsTroEIgC5NGAwWfOj8Ks55RKLz3sSx5joZFcv
j/Xf4xyUOUXIVpQlX2wNy4RoMiU5Shoa6w25PInxh/K9J3w4KPp3LXLrWrGhiWRV
d6fBBYB4t4TK+9uWEoUnT8/qOmN0D9QyseS9/KXUJqGDk8PeLQ9oGsrTXbvte+BI
GoiXwZF97EtlYlmqEQjNUw==
`protect END_PROTECTED
