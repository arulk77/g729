`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDeT0FjE9gUD00X4JcC7djdghMfpwBFNWrEtIE/xVwvr
dzxltSd/dTFANrIw+iJzkc20tblCYmYSiGpFjuNHctE9FBNG6XmQwkOA4eFrYE3l
AaFfsmdbnBJ4BBaYROjEasUOLIvtWTBI4n3502one8e0buj7+GVloxdYj/cq9nuh
QM0kErbUxJcg5HgMlmn9ieCsr2TnJQyXrF8/DZaLBhmR1uJAiI0Ac3bx+JMKp0jg
f9ml/kZXpit8T4sBPYCSaz0tK1mznBimhCoLr94F7pKYmTx5c71l6mnn6SWFEMME
IRgh/6iKsR0ql1yw6QD8nGniEDiHQufeQkkwHQ8+K4CHRH5e2jRO6QreRevWdE50
bnNv/MhMwVP1aaC9vpICifNMOHx1PteG/N7ggf0t0bCeR4E7sFn1hBQvr7DgjFrO
nO8D4WWvEFZGnHun79GT6dNmkDGZGaplikxwQNtTKDJMIwPMbPXPVh5CTMP8/F3b
0wHeEAktTKROr/apJomGVvBUphqvqhc3jH+7REydNZRNQkIJdzkNBTVyVh0/2kZX
`protect END_PROTECTED
