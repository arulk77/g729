`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAsdsZBYWeI/HDImeskU5/mjQsrXB5EPUczpQhEuIBF9
LK+LSDdFwadff7qEfideunsRa6v+Z8xixQSMVG5CvEIqWNrNVVBhqRAAA0KKuEv8
RxLsSjI7D1WD+QjvjAouDskVc9fvraT0TFzMshIelXi0aAfDw7VGd7veSsARFP9h
3Vb4IvXtRtOgkPqBa4Pzb5eBCydQqSanDTOtj5O3CrbS+t9PNHEvg8s9xlarvq2o
K4AuhvSYhpYCGdSAikrWBQ==
`protect END_PROTECTED
