`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xxStETsKqCDhiRXP4FcU04X5bhky1hob0ygs/GEEvOJ
kNdhoiqEPK1sjoj/QM4a8BlsKtS7w8rNQrDbTrNAlkioSiBayx0VkV/FIj3x3Tq3
JmyBvIO8+qvwZ2/II7Miv894uWWb5ZtGtTyBj80w6wvPp9MIrohuHEiAf8loAZZG
Ns8kUxX2X9z6vDinKVKcQ2UKnEu6+WxFMfKFXnyuby7S6BXYs688qOXn8akrURVn
GAN/AnrNKUgEbpoyWNKLAFzMcJDu5M40CVcBawqgJAU6Mptknu562KnsBrDePd8r
p4nIsGWDh3UVQ7DabEZRvQ==
`protect END_PROTECTED
