`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/crkEwQEZ9jwIlWpTcXma3HgxLNSReF/56z/cQJvJxy
T0qE0L4hpggvDYz4TSLh0qKinFsevzFyBqGogDNp4e3/G13PrO8/JRb9dhmt6/aA
Du68dzLaWpJuxxCABMv4m0XsM0uxlSIsmbcau/XhSrfLsPnV2WdDFprdQDDz2eE8
P8EMhG+o/vkSCRXlSs+tLdJmk6pM4VBbCjHcD4m56zQecScK9Nico1YGM4yoUxVT
I9ayFVg4fZ2J6s5zQt6cxArn9rR1DD+mvChnyxpJvpzjCAnCr8e9w8VFM2U/juNY
uP2br+8uYr23ATMwPNKyZK6rCtHmIRG++AfWSf2tYyH37hoOjHtXr9AYqMGP5hK1
Wf8DhxzScqECClpvMuf8vvkF1hNtY0YlDHjqMv5y9WRefN9WdsJ9qaGGjBxdMjgP
KB2J3DaFSY3j48YdGCNL1KzzfOR7fjYqpRO0ETkpeo8SZuvqBaocnu2/oy7ncECf
yQgVpcCsE4zjzuE5uI2iCIWS1ggEleCkt5VVMbLNN6GCep+YhVuvml03wq/sgKiA
BKP8TDurp56/p4LroZRBYU4uIP/ubg3ooISyBOD8wpSw7ZcGaaYPA0vPrZb9f8K8
Hywl/A9zTb99pPkhvMkb0Uq8jRThZXaA7NZNf8eK9H55fonA2RybjqsGNL7uHuAP
3MBTozzZVR/38CqefBNlEen+D9lEt+A3HiyVNJ9Boc5DcqgMKugPCU4SIYmEL1GS
eNmQwpiBtwzPWGNlbYGNyYWSJPF3IXgLdVF1Htl0PvM96fCrjUe4MLApqqZIBF+a
`protect END_PROTECTED
