`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
V2CAtuSj8lGucKHY+qCQNoiduFDWMto4lPvr81x6lsY0VINvEy+fOr3WIrfj6KqP
/JjB6S0Uc0Ixl5AU0XlyMfZGUreu4urTa7hgBNFwDW/QRCNtLjZGwz6mHpXg+0nH
DN0BF9i76t6PpwbCIvMsDSPOg9Z2/p5AqoQFK0064IhaoBHSXQ3u7qFd0k6FSPK0
`protect END_PROTECTED
