`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4USAQy7KCLMbnYCiHWqojHNtQVQHaVeqLYPk4l9fUPb/ERtuDvDJL7ExGrchVLw8
iFBzOhqD/g0+vmHcqMgOdY8J8XiHAdqnjbuF5wY7EXQoNL8eiR2KdCnyPSN3mj5U
lR3SAyfqS5YDD0hDETR7LIm/aepNgK4qTLi3xj3HD/bj5gnNm1M/w1H7PYG45VJD
ru8UY/baPCVkDIsC+ysPOAVdh/1K+O5BXdVGkYHTYl1c21sMh6tGsob69q8fokb4
iKRHR7OjcMvsNHCxuZVd6fofZuK+2TRFntoyQL3oKh2cbGZhq193T9/VmCcLh1cg
DNwgRihNWhluufm3XwSKJtNVa8lf6xDpWoNahx3PXdx/oZmDSNlXLIfpT86O0VAM
R8xfdQ52noHpvpjFUzGWJRpEjYlXFOQfwGOTgYxPJwwfVCwFy7/tVG3M22p0EuWA
xseQHMBAPXnvHImRVRkUv/FQqiRUhHfX1lF8ngMQxdVpJjA2ZTBxfmMYTow/MPnl
oqFwscq8/HwXJqW1902LyQ==
`protect END_PROTECTED
