`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4w20NY+b1d6Q+KFwaktunjsmUceIB0p8pt/Dy4um9JZc
ejtgK53yD8RIwrnsL26nh1YXg9SN07YKtIaXHHUG/Q9t8e7PagXPqIacZVaLG9KL
hDq9Zfq5Ctl5sqoaGMIVIRgCYii/rco2pErEMPPKNKe2ZkCSaE0jPnaUIERFwz7I
p2Y8x6PaHVJeI2uXE75Vx+Qc/c/RNQvut9GIAml3xMKH/H5NQcBnngt+AjrGGlIV
BPBMMthR+pKJIcKMAuHXHxKu9IrojP3nR6I5mp1rYMZ8bnZHzHyk7/I1R50ngz5R
4K+q0TVTtN6Jox6lyhVnDRR1kl3DVzOYSpo7JthKwaH0Qc/kF8J0V0kikjXgb8Hr
HxoyvtW4RBozVCoLE93xWdYCZSsdVvnBTQB5Y7n6JZk3clywdU2XBsEGRhy9E6O6
gYQIPAbKmKTnW15FTVaz+A==
`protect END_PROTECTED
