`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNw1AUhfKt9x5YQ2wHVJUo/OGJ4uFmC/nra4SOEqy44FS
0LlU09WG2AxAY3Va6wk3J9icfqKtXjq9AQfxOrlGyotpqfuEUOlT/ZQSSyMfkV4G
sHzKiNMS2WwAgJa5AT3Uovl8VP3GhPCqfhDeF35pemoZzRVItDQqcIxfRrw3n8Tv
BxL97mldMZd+Vf5yw79e1asrK7yBTeAD3TsEIglKdRzp8/VkHyiwdc1o1bR4KyLw
684x9ngwtndIlZ/0VGbCEmYviG22ODiGf3+5dEB00E0ZXPU7jju2iJoTp7ekX8Pb
ZcXUslKa0k4oj3oYcIcHlrDZyLZ1YyTxE0dotB3bYuqi3W//v91w0QsZ84PMU9M4
X5gGOTq7CLYd+YJvaygXaOr5kuY0RsG5EAFSW+NSa+BT2Zh3CX2+rvSUJ0sPoUe2
Hi1Vl2sI/obeaB+Lz8jGdh5corQxdoiL79d85Qyf+VKRA32THUtftGD8xXaUMa72
CwqPG43wrhHsFdu8CyPuvhzMeJx3tRB8ZjJ8dWiubmRPI37m6xUNWzYBY8li24wj
`protect END_PROTECTED
