`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEyLN+pFeZabNAD5CT4FG9Hp/QZ+uUdnrR3M1iNqf55r
PvXOy5Eb720tEM3JL2Rm3R8mcftw/u56cr5eIqVY+214JUfnXewe+fNK0mGyckU7
9BX35zcekoGH9s1Ap9YcXbCsp1V4MTSc4xDABgtXTOkhZ1zY0sbxDbz8SNL3IeZz
`protect END_PROTECTED
