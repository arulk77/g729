`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePRwsfs1QclrpVTBobrxUqkfpq3yC0WcLzKIilhgjskF
03AdOZMrUAs1P/6M6lB3Ilp1/oKBIBnPHKlnqzs8+z3hiL7+uhBUXM0r3TPsgVYx
I2q1utNZpYht2EPpZ9EpVYMWPQCH2B5SmfYRCspyWkBEScnSsuxzyRQSI2++/uLP
sO0Qpu5G1j3KRJGXeubIoYtBiAFlDaxOxTEnadL22Ct+QXiw0ia8Xqz5gyuCf0eV
MjJA8rL14My3AxtGpll8eX/8hp4FsDXCmkjgQXCixpwmgUY4irHR64tUUchLDYBc
Q5NFtEt4K5mOqcg2K/7hiQ==
`protect END_PROTECTED
