`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
uCy+KOY7zLuIW7IxcPWPkQw0llatSggBOVlc5Hd2bt2x/RggMQu9arjnUhJ9uUmw
pqPvEX4kx/IhSwPnjLL9x6PgoB1w83u3l2M85p0j6cogCdoUQmBS1wMj5ss0fycf
d/zMtEc46+Qz5ukXOfrhqZAF/oTAl61ZJXXjsHc2WbRgScqOkLnPxct0yv27GAUn
lyG0c6rWlb4p6IpY2yNWaQ2gdo3l9gt7qgOFgYY3eMz2yzyHDYRgvz7Dzpce1xIx
qEe47Gpd5IvTKSiP1ZjFWc9LO413CWOwyCmb4Ws+EG/akAwBAdneAFV4anZkm9hm
aVH8cUX34H1jyxkplTmlU3wT/GYbj+WFNU4RhwIaFkAoGH+fhhs/fMiZx2Z6Z1QS
pCKAe6ohNipq2t3pPywqErfRlJecVFGS60r59H+SRKC3dSvfODrQSKyLTI7gL8IW
YGS8LZn3Kq3Vi/JLntVEUBmVFWBZEvdEcZTcS3qT8a3dBh+WtHmKDiOhEAmAAajr
EkKwXEqhT6b66tyc7W5rdTJHuJqlkLOoduUL0Y4F70puLu5qTr4rw0GVYlzYFepS
1KndSAFQYnPY2nzY8377kn7zWw6WbuQ6Z1+p+qL52Ex66MoX6D7LWfyuuIqZqBUV
zsxPJXYk1R575H5HFQHNdQ==
`protect END_PROTECTED
