`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pnyY3jxGyCgnwWklYcFi/QSm7Dj/K/FJ5kSDWWMJ/w0TWAirQpeV67gpKUtABvlt
5Z79IaTySfBx50tfGLbuckPSEa9pDsZkRpdFIzuWz2l0/BjFjPOgR974BCCaLDZ3
a+KLSXmvmgs8vO+kLLoVTwPPU9ykCszbyi5/z2bwMNgBFVrN8fgoQ4VXCMD/7n7v
XpBsTHHwWJdKqxkchBHC0X27i421GN9YWFatnMHqTp+wvw710RTM1aFO1iYFqsyd
qF8rre9QfVDSAGkQRRhHQjjratNmChHv/MN0x+P+Tk1bGyKFJwR38dtdHnyEP5Nf
obH44aJIznikuyHCiBV+Xlzj6kArZCH4s9XsT+K+ggDSZ14d4T0dDNLVmr3eHscc
`protect END_PROTECTED
