`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C8Tzk4Tf7mZw0bbUfGmK3mwpknBA3pjoe6VeQFxGjlRM
zWPyLUwD1KnvLv/yM3E94VL2kuGawbqM37vRslqIg/inZH83M42Ql2Fv9JDB8lib
rDYNwt2SUCy39qJhnU9A1vsZANFfwj+vNuWVtSmlg93/Yx/t6g1aFVwlCOS8oNMW
fv/DSq894rQWxTK1uvYHheizlkxfoTOdreD9nS4H57NWOcX6Qql5O8nHHVqD4RXn
9crIyG/Q2A6lPCgNx22iugjGHkB8D8zjhIivmBZIhjBlI3Pj2y0kwbQHVgbJmR8q
LIns2FtzOfR3SWI8eddRIA0aLNaB9RKEk0RkblN4VGe4/IXMtuHD3HVg0vI8LWxf
SHunXuY7j//gZpFc1yKyQOZuYpHZ8HN63hCD4vXYM5dMvXG1OiS9rIdtpnw4Bc8i
hPiSVU7Lh9fftlJDGZtEzYOi9WdO4H3cqAuBAhmWDI3Z1OypUwtR3QEQKFbGAmaI
83423zdEvemSAdV+oHY3vEGtiPyDFGgCTD36+5DEWs2bCr0Ry2m0p6efDcZiPrCd
cfOXPy/OapB2RfeH/8tKuM61CR/3kZY3O/HnSLwO2jLLe2aYRPpK3v9Rjum1ChvT
SCumq3Dcswq6KnE/VdvIY3VadfuZt/P8s4241KXCRbo5KDMXthHKmnXDQ5WoJCrw
JpZ9rQ+URXO1jRF1VZqj02tQUpPz6eu1eV4KfuWFwPXnulXJ3Hee+GwJEdXLaWKl
lHx8uJiw5gLW1YhWhf3hJ/k3wkWJj2VW/2STfCruzSNaSn869qTEblbHZlnfTinG
Y15us2AFFwmwHxmz/Nscwa1EiAtDcFT9Oey90cwG0tGhUID0x76SnlPcXD8kNHYY
GxyfVLKOKe1KPP7hsvxGDpupLFdUSfxfAaceLTs0htsr1KVnxr8NUgOQQiPra9ul
k0DTdQ4pxxqVT46LjAGYeUaaIPQpwtFIbT/5Gcq1cwgRPaM18v+6Dv9yXQ4h40Rj
rfVshp4slmIVMFIbV5NV2k6D2VAT7aLVlDoR5tutRs2bjqW41kR1yfIFW/n57YLT
2gD36oNLH5Ns47vwLEl6zlDDA+bGqrgbLHDqbZ1U5tX1Sb0dUn8eH0dyIJ33sl/w
s5JemqklexYNzSNpmv9wI/ojkzO8Fc+sifnIBg7EGqPpDhS7ARxbxzo6zD1OlZm2
kwauYehq8rIqSqISmNc2IcwRuGDct7KM//MCuQeZrIXQqmlIq27bWPxO6/qYtOLE
mVPyHABJarjnptUu9iN1pjZNzE/HcRVn3xBYIo3VB51RR1C3+nFsPsMmh/5PL9Xq
MIsSlyiPO5uC5Uwp4Ai2DS4H2LjCNpQiSBt1dEv0PMTBt7ZHAlx0Y+0KjekMT0Ed
xD3YYpRwCqEeZiAL2VOGf7MWkibJlnncfKMYi8Esbbtr2n86A8AWYBuBoxAO1f4e
YBjWbAq2ZV6y+pcZITrRZQQIWhiKx2BvwACKCkNXyWo7XvgRZcO8zQ2uDHxLi25l
PoX6W7EG9KyTQI2y36CanzSnS2qiDvCudk4bOodQq0dxlSGI9y+tioJvxHnsT/yj
sgGgVX4AdETbYDqFMyruLd4BdZoDBJs4A4R8PsGQ81w=
`protect END_PROTECTED
