`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1abr/mDF63EvO+ZztT3Sx3oNRSJALFellq0yT/LuhCWe3
j+Lf6JLYkI8exCatrN/fT++Hb0XNObyuNs0P0+7iY2tmaGo5x5Leln6LLcVhk3gy
z8GjaP3oWgMrbUrhXEGziSe4FAP+XXA5lXA+dTpownVhxA7zHlgwzfkO8rks5AYw
9lqF8mXre+uMXvQcHBimqbLeHu3PAImTb6BOM5HmPFQH5G31BFzG7dN06AZb4C0A
bu5Le0yEarv7eilPUyIBWCYW93/3qhQLNYInN6TJHVhJPHwIdcP8xwLxdS1y6I6n
UAO/aAZEvKPDbT+BopQzxndePwDjsewCWIcPJ5/TyxjYYzuUA28z6YdKtLimpQnw
3ukvfNfxf9v1PMsLc8j8QMDkI/rGMYkI8QsvT0VNO76q+tT4Eg/WBrGY3/QD7+7Z
JMQ/2IPXJQyITNzfhwT/AcpZT4lWW9O8e7LAdUUky4E8VG+v3fihczv2gRVsrmVC
MN15+11qbMJn9jXBL9jjZO/9ez937ja6i61yjkjuIVDUVRcHVHf5S+pH0rhwRg8S
XDD1uRlER13/EQiUtu3EuYzG86DvtkFHGV29QbUhZhsZK6eAad24PphXjlgRqK/5
udUODNBBJVk7V4yseffytUgYvjQzifM+Uy72Bfih3m6NOEI8IVZddWlLHgVcuzLt
78nrVlLx4A0ox0upECwHds3m1961DQtkeEMmK15Yk1ql8gSTy9hc+JvL6Ydrq7tb
DwvZVx4uVcUZ5eFX/BksGKQKLNEbTiLqCzlL9l+pwRIeiI6kfv3+HhRJyIWOLlOs
IFIdMdwcL97ALMQ5WwfODaqGJo4ka9c+2KdNG/4WlbZDIJ5BG+LlwGTcw9hc+4Vb
YIMFSVF5otXnsOiS3r1mcVzzW4XRiwXA8+/7jp68yS0bpWa9t1QG+tiQCSaL84bM
IFauKeJZ1UOMvAdkSJe/2uJh7Exl64uaksDKOyivpahKeWrqIs5R2Vwe7Bxd08gf
5R4JDUvDc7cx4sL+N5fjDvFyEISpvosXhPl2Zhg38GJVkgeHW7tQr71l4ABTU/aw
zD61NZj0zTVYdP92qu+zwhfYcGZPkcm1a912I3Qz5B3qpgZUO/yno9Qvp5Z1WQ+e
0BLnxoi1hXTKWmQpG7YrckJVepkQyC3G4J7IQlCRo8BAFQzNedOfqeTDGw8s4MwF
I/O/sZvWSYsXEHVKKAYzlouSvLwVyR39W+bJT/MnuM/srt2E+pHx6j3JRlNwb0lD
bXg21flz9YuzPXlM2jOsHiQMgUVJ9fR35BndgRjylUa+y7f76U77vFpBH7VGmNku
LN/iJO8eEBZgfBlJfw+NBWOPEYlWXpzuN053oC4kas4m6T2INDnVPIs/Nht/ULez
TRYjsDuf+7tNtAGjiuwJdDUEfvT1Wh9+hcDuMm5bLBaihfk7fofSdbXPOzkp2Tjw
Sdnd29Ss/IkmHJmBvQ++7Zmp/PTaSZ86QdLupuTwSNxN63Gxv7owmHfaL2ftdNFA
v5Kz8rRzlBqIMQtKweq2IsqdplLxA7ACvGxXvv0asfrLPzaab9PojvPOIz6R8fT+
5w7GWJrvkpleUdzAT89CV+LQ4x5puBRy0GU9D03eEEF5gqPhLmwZfxLtjI1/Lv/0
LNXohb9BiyfOvq4x6f1SLGxEve4fjY+JRDhyjEoEpU4wFGaYFB5imPSgk+5ijstm
jn2hOPFyZ05SJRi1/V2KjPgpmSaLXebJYswICy5wcOiENasymprTV4O6q0iE901H
sY7LQtjjses/pWaZlUOthfIVKalejNIHxOaxQZvfM0+BKw81mSvzZClsJbPy4/p6
r3FxL417wCGDQAGTu4CFZXD4W6bW/Q7WVt1JCREyXmsgUPQ19r4x582Cf92qvVT4
7AsI/r3EaNrO670fk1Ylzkrdbue3QK00VV/pNj3EKvRggtbgsbhxJGgBULuHelDx
0zRgSoIy0O3Kl6g3y4h0NSZY9+BW6UClc/klaS1/2gF6YGX4j8p88TPANQztreTh
W0e8O206uHX2f/5FFsVq6jLmnExonkVKtbU0d9AcCupFWuZgWU5EzhqEk/b7XJQ0
9hB+NPHn+sbsYXXrWG8MtWhz7HMvfPEiDfGeB896q+1N6h727xz9CbhgfpqDp5Gd
wTRjEeSirN/uOwemr5gRyqKshblOUD6N6LD8gpXoyUXfyh+JlV9sYE4LGwpOZqem
1wuj+BPU3Y6ZXSu4vQm7FQp81Tao+1U1Y1Wk4Avp9M6RUnFRRMSAfyFkvCJRBpIZ
if49ADqB3o10dMrth5Dq+f8QydtthlwEOVcs3SBJWRMZxI+LmlwNBOwzoJhYBCR1
m951e2qTB7NyKd7xKb8pFQwf9lzI11/lX0cxVLF6/WtmMn8zRC2EDoE8/CSkaEqD
eU7d8dYG0PLDYzdnYrcQSMpKyLidY/LbG/xBI/SrycXwoynkEwkOWKpLQAL2jcIs
36zxCiRz1ZpfAJRF3pL45LbKXN4jzo6zuChm8O7cPQIWOBS9/IN/Q/iUgdVfSacj
gWydHSKHdRh+lxcJk26mp8QU3LdJqCn0PbLzuCruLZJQNPFnUIB4XDY2zxYVoqdJ
2waAfR2mo+hls1TAnWkbhKEcnKKhBxVh4ai+ybbzsu7qYgGSJCxH8//mV+C+pKe8
k8Ow6K5T4YGPefcW2JapEoBQbMKDrM47tdvlGE3Tgf0ZXCArx/6ZCTEkHPYkKmAo
6GVsI9jWb3JXPzsBid+w6PQXy7oX2Nqju9kELAhuhj8Eodl4xOBHXv9669JdX2B3
+hLipFcr/eH7UrtRa4YcA9tfFKvapcTjZG9FpI08ok7DMNl2nmVVIHNH7y/HN0mg
GOHsGIWxoclEaXopF6tDxuaFA+T5qR7Iwos8bCIrjNAJgYCFqycANox6Fhg09Wk+
2XSkSVbRTyDaBWjs6vIBylLy6S7LMP4z1JpjVmnJYeDkORVy/MZnsuRWN9ZSdyab
wrNlVlem8f2iSxQvJPfUx4puTEnEwSSZaCC69ctVhQPKLUHwsScDOKHTuwIPntcF
nMqE6tIF1jeVAUKonxpLiA8SPBXtsXyE1cusdQ3zf8AXLufhyZxWSGermjMDvspf
76S6RKPyv5Dqja2ULrIjboeqErfPd2s/Li+DXgUVmj5Monsb9fhdgN+2QE6Iz8b4
kjlvfinzoK0P8tcbB/R4DeCms3vcWh8+E1vN9+pMF2hkLoOycqSZLJUd6Zvnk3oJ
0GPd0ylzypGFuoxk8a3oN4IobDOq8JtlUMWAgy98EM9ahdk7fxgIaCvkY0upHdHR
c9tA3EnigzB8Zyr8DrwsPrdiXkRiYq/KBHe0C/BwFCA4hbPiilBv/y9K6dsAcDVz
nkzN9L88JZ6Kdlvk9/fwcmg5fyAzL3jN2ZMp+jUG6d5kY6D3Q9fdTmsSm4il1IZV
3INH17ZGFsnTXD/1Ic/pWrfhYrqKPvNVIXU7zsMuTuE1xNfv5MWkjL3LmPFuvwf+
zbwY0vS/h+aac8CoMxXYQxlGh5xnF2ussUWjwy5wsnaxwx7iBN3y6T0tJ84yP4XH
i/4CWz37wy46fqyArbaoh+ppbSWk+zcFGokNkXokgBoIcFBmtBVoRbiYb2dDHUwH
wEFvpFdCFfEeArC0SVbx+wbJFSQpSQ2oWDyl9USA8cd9rER3ymFxaWxjxMuz2rux
xnm+j8j49NSXhfdd8QhX82LKiIEB4vFLww4aCyIadXPpQlFR7Rpjh7JNLpCv2Nqt
ju6pkZ0LbHC8/07X7ZgrOSwtM59UkgSesQrxIcJxxylk7EAtZ/Jza5NBgB5Ch7rC
Tns50MkCrWMb+k5eHr+znuca73fkDQ4hXUYEQe046mC6vy00E6Gp1mUL49Izn+Ew
UUZT4Ht9VDcoknTN+KJfrAj+OPG/8WmyjFR6y1TSpcalrHEHxKbzdxyG8WzqJt7v
TYXdrVJZcF1klxIAoluDEW1EchVAltwpZpbzHMq2gNWdotAQhswgCInrq8RAdb+l
Yl2JZIPeqKhSVNqldpca43dRjxj5TtDCu/DZFWaRSZTTDtjFTkGj3tGp+dF+yb+0
S9pg9Y6gFJ5S9VtaC7Lmi0dOKngvSSurMpOI1LutkSDA98soU9vgSyHL+cdUdJ31
aMAfnsJvtOrPNCO9SvGHR/0b6IYQgUtSwVuk2DwNr4/nUAcDJJyMNBfM1MvAmu9a
mRcbb7DiiGN2rB7tRj/rElRv/dFK0QutKVYfwKCyB/Nef+pY1tp8KqCBhpb8MKRr
Di0WRKhkMapYj6ik3r7UHSpuMVihGSzdV726AnENDMWrI/4vw7VuxjcsK0vsRmi9
+9/QxcbEnUy5m/lNXDuQichHx76BG3O7/z7NpY6R6E5eq/AnhaQXF8eK3/8UB7kp
aZazUdz8SEsFTiVHWPw4j71eh3mIVyKRP2CqEtTlnOv8Metap2VRcFhAJX7zbi0m
1V8uZy6P/+9v42tJlzUxXtAuyqQNfzjJtaNmHFqg7ml/YICR0HcP8TE1Vgrwu9iD
AmmhvmfUhY5eg60xn3QQbFDgvM0xYfZSuE8qm0NGQd2wBjHkABHOF5tFNDAHfS8N
I/LMSx9Kf1qSagztgCQQEK4BZ1iSC5eCD/Eg2ncJHTl4g6264T+YNW3igIaOrIFm
mZCY9ANIZwuL7TzJI73i88WZAtAj+n9BzT1yXRXXWKdS4Y+/Ntsd+2giIaL6Aw3a
lrEQ3ZFWfbqO8io359yQGpKzP9CR23+bJquInaM5zKhDGnUcyaNW3wTWNGe23NjT
9eP5Qa3kHQqArkGf/GZLfdZeL4TzimsyTFAewlolv1b0DPz33IsVfz902EMiOHRC
5Tt3+Ocr+J27jPD1XnNpaN+Bi4QxFoDSXWJZDRbczE5W+Ui/UiiYCgKxkRsuBfVP
KrJhEbPVm9RD1XjSPmCWqh+MiTRflyzSBNXDlKFKAP3MZagNKwEz/oCTtZNRFbjz
mFYu7O9gN8u2+6W5C2LKAzUg6YRULFqgOpvkUlhFt5zVmaK9QI+/8Glbug0VFdE4
ytsHdCLZcGBu3jC31ItrQENypZaoRoMFZLxQ5swujjjxRPf1rt5t5ahcyq8H1G0H
9j420W9GfhoH3KmTVMgGwKaDZOU1IaH/eGomOak7MFQtW/0LXEeHxz8BmhBGkTyt
oSygAyQzNOgZfJPcR0XRXAhvVSzJPnPu2XxT7FdqBNj8fYPBEZUA1JwRTVeUdK2R
VsqaSdetxVQIKzgSz5YthKMP8qAhcdOGljlDea1j3fgyJTiWVeFTMiEwwtZSUMFu
fJPXIGtAxE146YUfYL0k+K/b5KuXzlDwXmHUzTNg60wjbu65k97CCQN4w8YX2uF3
ICZlRsSUecebWIDEhWiX0zov9dJazR8ZbCMV2WB47tcBXrdh70N3OAzXw+y8X2Sq
GULeIUnkoPQ5V2p7djDqZiAt3wqrFzRg2SVGy+AX/iMr52i1shl7KoQ3wOhutVne
7Bb4ofvWzSsJSkGtZY52YD37zXo1Z/XfFk1NARB0nN2ANXgj5qaHxHdOXbgI2sMD
c5C6apiyHt+ugJQBtqz6FF5mfogTDzVTlZxzBYz8iaZfhuWsly3KhOZ/E75gs4F+
YNxRUIhOJDnwBUSaoFrvY3qXxtgxd+0axUJpMeIlWJGMii0Lt4XOprAuVdSXfo4S
3mW2EvtpPXiX6sU59/QM/V2QlSGzUhxa3kRPnVPBuYMj1mIJyPJed1xRcvPhMPqs
4E31uxpTM5Agch8cLPH/tLGpUuBrnhkCteMADoZW+lHvJ+R53vYaELZmCTmoW8nH
c/M8g51+u3W7EA1XeTQzFwK0IWqZGsA0GAj25zEI9ndkGOtabtAtHlFNh1H93Zw4
xiLp2nh/aw35lV8Rd1Zsw8184m8XqmeBQa9Rav1L5RlzaAAdJnxtIXME8w/tAion
6kNBpzk6krIC9I34uGrpscX0L+yxRXTdiSo4yysXka/hjefFmhqWTyigSdN62fey
kCqiPF/k5XXz9Q5cycnYCdadMcZICrRnN3H1PZwMkhBGbfLG6PI1OLjYaWa4E07G
KXGb/vlhUFxcbrnBO1XqdQTaTR5Aonaqk0G7ugO91kww26gHq8xWgrQqWShhI1A5
g3pr+1FFnEABIexVadBj8dCI3HYObL2k9vaP5rmCLMRagJ3OQ5tB0dG2EqUDJ0DN
aDRmJkK8AxO6vvEb0zPrBcCb0b+OBzFWeGRr+3vpBa6tYvat3sU3Crn14Y4Kdtjo
VWY5BLrXPXgdJ5Iuv+ZW7dwavw9pXPL2D0Ce1dIBUsmFJU12yNIHvzt4mmQExj8/
MekSnpqs7pwJuNkoij2ZLDON7WoiTFDn0dJy5k1sZJunSJCdx3maOslqTRWiYhuL
jzdJG1j6XzDd86f/hJcDUxhpBJxtHsncPdq9hlCXCjwkTeMzkMUxCb1wcJId2fJO
kppqXlACHnGuRXNrpYxwTo6Qm+7OzG8tw6mEt9dZpoiM7c/wQ3a34U5uP79Rra+b
trAcnc5/EdqizGoUYbIdVMdoVpZqlkBAn71x+z/1pAYjawAGJPJ/tbvyRIt84/bg
M5ykoru1mSwXF0jO0kbgvYPOaue6NDumBEFO63Mkh0mmIdg0W2R6BHVwFjSWtFm4
vkHbC8bZ2Q9WPSBoBcVE4VEP5kY6BxxUPk2avEE7+TLMGEZWS+Z9UYcbA2N/MFGU
XxLciVA9vJ9GAIqQmu4MCz0y2Dp8r1lLbW6C9q6E3JhozVDmGikzovdPYiQ1FZzE
MdvhA1+wdgLVo32q2Z2x+dffYo8TU8lA6bhvNI/4GKUdDZcqVKwpo10ihLUteoVW
+LGOHoVXXLjPQh91joJhl4tR7i1FlgQcJs/wpaOudtb5wmKoxEh5sqpJ1V7yj+vZ
BoCBOnnPblwjaQGob3UCGR5Zq/mzeow0CnWIpWne2eY3iQxKnphFqGl5KeU8PJOB
Rt8JxQVD/PoZP/djgG/dxiWoTBJPZiw+2mOykcn/QjfDXe2AkgnG2F2MvN1WtVsc
acTYlfaiF4oV6BYkDeUq0QWaXkTnzJh418m6piUugdWXDM/RXqeZSC0hr2n/TQm5
2MoJE6FV9eZ3mrb0qzuTU46uqGcJUfzkNTdBWBgXVzTMYGUtUcRbA5Tv8WhY8/lv
aeo5h9wwVzKh44EPWKfVp3EQKiLZi67BOt+ROy35CPx1UHEFnCPIGawV3jOJPghr
n1s36tDfk9baHOuNFXDdg2t+zZYYMra6zto/NmC8VQTpe9hFBltcVC51/QpLvZP/
5epLbSw1N+A1cBcKY/Q/RQB0FupNhSD731rg9IS/44wSk/I2MZxDDMIQVyR9FlC4
iYsHb3EvyPlS4pVI1LfLDDxxEyeuWGlh/SaucxSt+o6BZXLo/RZVSKSVy/oGT2Er
G8Dk9Pa6SWztNQGzjeIo7xa03rCGVg0aBa+IIyFBgat+jY8iHBf4xxw7EwsfB8V4
kSG2w0rYMyE8c50SfVrIPOw5ytgVRfgGZ7OswVVZ8T7ybxQcIX5WxBB4qfgqW7la
jg6uNYgleEY13/wbgHjJUPlvDhTsdZ0LpQPp+zSt5k6Uy712S66ndjnvewep8izS
+D1LeFRfnO7hO253WoufMNUrzNO2YL60cMkC4igke2VhWSpQk1jJc3CjnW3FxG4T
WZAhFslJ8kiHsd1hQGQC7uWpxny0pZ3tC6DaEvHK0f6Dw2iIuJjMPVGM4/M05vt0
rkkXY3dNHqJKE5nOIHRfrzLDCyx51RdvlCf/e4Ap90PoFwH/Q2hRtRlfz79O12bN
OWg8kFNYWaVrsbVVYoCrQuKmjLyDI33fGut9DbTmSz3/1nHwFuPY/D0LbtUkc7LY
3v+CpNTmoGwwHpoFO4yb55bKk9kx2RTDrVeBqo62fl4+krItIFpV4nM4Jf9+7DHb
UTPYwx0Hkc7pAW/rtc2dIQh4Ax4sdfyjY9m5RnBxCSfpO/ekhzxEmRBZ0vdAshkL
VkHvxKL9fFsY9lIvj3nUBu3X2Rk8TaIHLxgzzIcoUWJgFRGvoAOpNGkUXQGrT2Yc
p9uXbFel1M1wiLmMsvoH5LOhoCpxwrBlFp060ESsJ3uF5FP1BivDuGlDLzRdVwhm
2LuuL3RK1R3X44sqRrrTTt2WxewxQixKbcJezzLA2iKFogdze5qa8SwY7jpH+6Wh
ka2AZW57BLCWjaFEmeskYqxu+1sVLYGtpWW59g8IGKFm+yZ2sBlCxcWePh+7GT4X
dXMT7FXQcCtxh3RlhUCNcDkACicoz8fMZsyX2e/KWoGR5J5zlemBRHUtCyFMYWGI
KfWpFWPgYC7R4xcW5czRIIy5hED03UAQJleyD+hnU/0SsIZtZP0AV9BGWJGYjE+X
C03B5FWJ11Cav8yiRJut5E5dwHycrAjE0GJvNnSK8jkSJcZLFRDRZ7VPvXBsy67f
2S5YvNPoUOAdwu/jPvt58pMPIC6pIoNocZS4Z/yUiBqxZF4gHj2CFVDFf03Fh9zX
PPXnpwcoJ2L+Qe3gGTAn8j3/kX8kepFP2btL4C59+cIZ/V8PAuQoPbjDsiiDPhyP
7DR528EEJn6ncFG6cDQ+Yh1S5xCQh81WayDoLfvtM52jeLuo72evxYa5n3OkwwRk
rNh1oGfLCyiGpWlIdhFPIGG7bJAgRDOxr2s6td6PnLIslXZyqKBL+XOZxcoIyyCR
X3bjLt5n76vKsR1DjokhQhRo1sD4ibA3S3CU1hKjlHztpvjIiV0+gRucFWgCqLQ2
5zPx1dL0uqNYpTaUXYvx8ojQbsPKEntmMnLpGnzbLV1qjl5eZ0b9cojSoCjdk7+j
QMR0JWMMCsa35B+IphKdcJHTwqPW9pi7xLSlDsIKv9zr9WnyQA8Z+w7ZHgxgTzxV
klhXnoGdViz1kaIEAUm1wfaWTgUhnIxh3Jw+9ax6OgQdV58PTau+2HFOT5XIKelT
F1ZjAsQVGghJxHTFDR73sMb6Hp96f0gUOqehg2CT8/SEGp8F37JwMHLX0zZqZjNy
zKRkS7ot2lShMXLZgjVkeSO5dZ1cFqftVyC3zG+dwVKLuiMGZcWYlxb0jWnaNba+
BszCJy4FDchsvM/FIm2jTKnLqlVV79TLh9OrBD2ItIG/p9eMleq8GVHR8V+csbss
8yDQnBzjnFXD7E3q/TiSn7+XEoZciNMuJwN8j4W3Yov7NzZyPmHq5HRbz6HGDga9
hwOlzSoRpNDiPaeK6tPC4q8fUn58LGF82qj7DrPOP0S1sqLM0OPMPTWB4ua5jFaa
A5OnVOt2fJU4wVJOXJIeOGDf4uOtVR1RIb3h7yFg6Uvto5esbtM6RQhMY+3WoVks
mpl83uxq72r4OuatxOwnmJo5+JK4wmUa3JnMH54ILpAzuD7HRWjWHKC0yKAStLtT
2Nfdcp+jDlEnSzloAxyAuyxK3K36K4APL/CgYnw+OPn14AL3dqE/f6REPJ8bWv5g
OvYvHRwrODcahXv8eRoRAPuobWu+ehYFGJl9CpiiYQAZnVGrlmvQyTcQXuN7YJCn
BjYXbMHRfZ5aHnNUHKk/KvfMByeZ+Xui2sKLv77IzkeTsPkBUhTb9xZKIR7Le1kC
AHgQzxg7iXTZbZzRBfGd/GAZYQ6rH8QPBEy48H4Lw2pjR94PaSkQz+Bfem23EJ9o
vHu4z2PuSSjnIr0zF+wSmZz+h4tq+g20EPL35HKgG5/+iFF7S6IpRtGxTatyc22y
pG+p+BeqrAct4mCnv+Lwi6MsPAqUqSHi9UiXmuXjPvUfJRZLSdPiXzKW9g+P6hUI
1stTn0OeFj6knDUDML3h1vA18osbCFG8wDc5/CzwvyDOXr9oLOLwiJh8P2Ij4K7x
W/IsBzowYXcUpoFxXbzsx5ATvpWhOpyJ3kJ438iR9qmjzo/M6wP5a22c3PZgxnnZ
SVfqEF+MmXidKBAmNt4Nnwx1Wgc5xptBRlqKGkJSDmFgJuCa9/icDzTd7HInt4Ul
brT3i/L3pitqyJ/owsWrBYSUejoTGBwwEytad06lg1TL6W4F5ljdb3xTrahMLlhV
2spVW4uP/zT/eB3boj4plvZRCJgShH/agxyog8aF0wcvuCFb70UjJcZP8fznBSUP
92ql0dVrqUKcu9ZkyL4PGMfujjcQAtdbmL5+OTzJzSbpBsxMBnLTve4rcCxsRql5
jS+LQqpFcTBx96Np7LzCFQIJXJ/aDHAJAeWi2KIllmYL2HG/Fp3BpQmoa2lRIu2/
dpwe/8DeKd2y/GCrAGnQqsvr64mSox5a3noMGaKYQGuSaI6CZNbx9pcrrCm4a8Nd
iAnAZJqCyR1ThbNwNalMcL39c75sXssgWjgCRhI1JsRKy3cC5kw19ZZuPeZmLH5b
56fWU5bGsqtCwJbAKFUoCGaUPi65dvYZqO+On89r9ZGQDQAKrnEqplEjoW+OCZ1J
4pZopdxbOvvuWpjxkE90xc9BNQeM26GeUttJWAEn439kpBhV9qgzXMhuqOFo0fP/
5chhhAoLJCmzi+8zzGupkeMCZ5DXdlyDHVvY4Oovq0qzsXNew6iemOF1LHdI1lGT
GZc8iIOSjw9dTgOx4+JnZGQBdfzq9aoYgNRhK3Qh7CN/rkUhjQ8Jw4spmdVH95sR
OddofQn/+323X6kIc9DrteYwcMH1n1ucUxT30WU76LfJ6nvsjEJXTAZrT+D5evBl
le0iM1B0kCAugZwXx2WIGJmhqx7dTg9iR+EJZv7LRrZ9Ul9gSR2r2yJGh9VggsdR
4yh6mINdsDkHqNNgNqpbwcIdbV41vVmKkDpUBY5GsPv/9q8Z3FjxMNts3LmVFrjU
ElIa8JeeYEMTFBfO4CxEARFDWkQgDgUuxtTXQ/IiRb67mKc2aFUURaUkN6EGoF0V
RLwnAukZpwWWYz2WJE0E/HvN5qlsEKWPLIiXTxBv6QL0kudo8ith9wRhtCtysyfx
j7zS5SQeEVX4cUmYHmuHTfF9ud9EwPOX8kHlQ6q6nFWB3P19ca+/i8drHNMgWA2s
3TJvtsTs8QqvvrJj1FKc0yPXSgBoc+cZJbV6YCZqlcAshi+CidAw1/hqs0KzDOWo
OFPZv3QcvZgzpuaRhCo3tCumLki5OYQwUNJiTpAHKiTvnpWAjamNsAXzmlqFUJeB
TO8juFrVySPl1vGwWW9Kf9fm3+ECBsdiTpze3/DAXSLZHdScvq+s2541M7dsNSKT
8dH5GU/7RrJ6RXDE3iCicNVWsJc4qQjTDRaN9gaRuQqQFGLHfuaUm0OvFW9qc8Ja
zs3ZlFsNLr6auf66WBBT73egSn8BJOi7koBeIDyaGK0IXNm1BDKHxdFEzuz3l69K
r3BdfxFQgP6PKBuU102xEKtntqCaLixQKxQtTOu8OyRf9aaREPv2U8gC4kpg6jA8
UWAcd9GqpUTSh7601SKqihBdEe4DLH9B7rP+UtyYLP1BEikhQ/aBGcBrlwsW+0vU
E41Y7XevHQXBQ5dWsVL1drw6mlkZ9o4q2lyQFYeo7S9HAvMbTet+B8rrkFK84xqL
v7RWlUAtBsqPwRFU+J69dzrsVMmT97KhKR5WRclxuAy4dH2Rp21rfRf7/Yq/ua/I
iUAJVIGL0/ez6z49BUIzbyf4wqaYQtiJGdQIbguDS/xRhB+RgP25KRR6EUnqFYCi
Oxf+1Y/fVf5iZ9udlsybMetwntEEnyCrI9rpAUPVTWbkRqTRMVDZ4Ij44Wq88b9B
Oq9n809zm2zhopqwhrh739jkzHZcLkcOvlNbqOla2k0SNXY/d019uCO/2mFkMzih
YAuHRdhIAG1T1hZyBBhsCZx+qcgehrLDzp9p5F2fsn/NiWE0suaBY5uDtd2NnYvH
2l+GvKX7ddGZr//YbsjI9f/+9Fj0BHVrpLjj/H5R4JPocTQHo4kbFO6oV+zsEiX5
7Kr1uELHsb9wPa+tYOAgiK9rNAAplBEdUCC6PwTSzOeJ+Xvh71Bq21zGFbn8jxxm
v0chljEEvRXXk0TMa+zwdd0/tw9dRf2MWUrb/dONeUhxeNZq+6VJz4Gvcgt2h5mL
G24tz7VDz9BhaLqS5ffFY5+Txg8D9mO7Sj0hNkjzrKK07D0PHwavHvJ+h/aOb/sE
eRQcH9mHNb2Iyj+UiHwM+LYC5RPyWhSTh5X/cK0ZZSCUPzeuKuuqX5sw3QPNjkOW
ssO9WfKB45DiRWbwI/sLXH/X42eAqTv+DxD7mE6CxE3D7j0HbdpneTyjCa2mjYRM
3uu5dxxAyrK1je3ZvqPmfvL5yLTuukRz/UB3eJ7k9150h/hTRKK6WK6ZazZftPfG
cMbB5/mdMTPbOkl17eJ4UrAzuCtLOtEo8Ese0EaNVYxejvwz+B7zJBjBUScQd9KN
m/TXJA8gD4uqlmrsaTmm+cXqB9XPWabIb/p9God7Ev9FDLynxBbqYxgrwaH7gGnn
yatJy4R8/EuFCY+DwferOvaLw2p6EpLSWO7wlvKN+hxF4WT1QDHkb27U2TXbAvs4
8O5ee0ocwJJ2nMrApuv4zjBd+UkEBdsXDYmtlJv7aLlLxgig++ndrjEmiTKjrzKg
eOI27DGUoPytVQbQf+eS2x1ztaR60ApaxNlxtI0mzUPyjyvRYsyRJQRw5YgH8Vm6
dAtkvtw3P3Ih3e1f1HiTejZS+gjo+QN27rU6UWvfZaXcqj/oDwXt6XwO8SNKFWdT
EJB/tyTGtvJ+3Q616HV9cFU5f0GrPsFuaEVW8+KL8MhP6wbhSZXHvpKPuLj7Hjnt
fTmBYZn9P7xy1go/tZjp0iSz7qWxJRKw4HVhmB++sLgWHd2G5zYK6eLCt8fnNeOv
XQFG4ifNmmrm7LH9VGEyg0+G9pLRp8UgPw2g850RbjpjHqL/u9nGeJK+viMmBVFt
oiQnrwtobDl9ZuVD0kJ6Q0zz1Y7hK3wbVisrlpQEcLMwP7MMPZs9qRuAU65dUqW6
HhQWLc75P/7jhJBxIWNCgZ7IpTWcYnZmZCsVd9Vviv9Bf9J9mnLsvJ51xQcjKtEp
wcrJpw5b4ZWZWgF6vGhqD6SGU0999B2BletHrQ8q4mksji5DmVFxXFnCqRGGNn3y
9yeGJViWKGWPJUOPub0ia+hx095LWqHD9jF8+YHsSyseEW2QXDT4tZTLlRpaabEd
JU5PW0AynupcSA2poPHHiI/SdVNO02PugGKS62PuZee4WZNe70VU/gVyuDgP9Hla
aaAgf5Ay/WI7jvBtnEKuwvsOf6BazWeMRalOotgZUi/NpA+gukyZTxL+WfLrSpsL
QXI+VMihfRyagjsIOjJZq6M4NapoM3KU2adw3Yb5KheHmA/GmKCsgDKjTBvFxFgb
I90NV/dBRIrH0h03t6wH76UUKbFLfwRvyEWOyb9v6cwtABcrAIRdm85lJvzD3GEB
ZWM6q2AUzb1+IQmXicGfU0NYzfU6zWfl+C4I7sJUQScAXWa9sWHhMVbkn0ZntNEp
NxKl5+9ZxINzovj2kBDLfCZsZ4ULKGMbX0RLB8++T+BLhAcwtA9lJ6KVrcGbip5Z
/nUwVmlP8WwiqsCbcSnfAm9taUEaOpk7dz0+aZ5Qy7c/XMPkga75s4eUnF0eXo1h
nj6W3/dnp9hUjqrZLVUIzi1iwh79gDUJvW0OwBc2EncJmaDAsL466eYHSxYa795n
DfM6aE8NwFy6/RkJpLU7r/8pfcX8ify/8Cs0G+zT8e1bJwqrOCOmDHTRruRqZMKf
HaotXJl1nX7d/KniyyC9NnJoeehuuuj8/FpSMUd7OT1JvVwnEIkImLofzFYXOcj1
dLMwVrGIDwfR7TdWIAs7G6ZrGmAKYgiP74WvMCLcTId1wCsfooFbXb6peJion8gb
c1RGFS1zp3vZQ/4uCG4z6dR/2LeV3hocOesYmNp80q+KfsqWUwMETEKJmtYJ0+Ia
wzmfmxGHllx0qrr4GFiCofzpFbYB7PMS1wyqnNfi0J3Rz5WQ7eCPcm/hswIGZBos
xMggiCZGKRbzp2fYi/hDYiXTNh2jwXeykT6ygBP2KGeat8RpX7nZY67Sbp0j+1p6
xkMwHRQRyNIa5eJJKxmV0jtjDUJew+bwT8kS4bxL/LAiInMsV4YSdIu6Ol1fkhVe
A0jF1A5xTCUlfD3nSGQ+4XH8VIKLd6Yc2eayExjSuAwVoQ4wkmvOW15HJqpr40o4
g4oZFYNwBY4HMhkoTzgvHQEywMkkH9mwmNRRHLFxv93SmVufPhUJk5yjTOOMUwjZ
7S/6k7ZBmrQzZd9GG9QJ/T+J/3vzEYeNB1sKBIASRnQozSxqQLDLfwG6qLEBYx/M
oY9lJHWFbdrlsM2tj/ckSzEYDOSpy2RnMygn3MteWwtM+V2pR867jOzUT82CQVXO
gwvm+11tlK0uG/c6YTg61mVASPTLaXaD9amVoRpvYcZdQA8WocTFDDVoo0Wyt6QQ
/LBZrE7acTpe5XRguPWYr5mKsp2FX2DsJpnbIvNII5Dw+K5LWXlWWDoJ1iOZ/uyS
abRe5Vhh46u+Ou54iATX9BIfbPrfWEKoNPl9mUEwWM9kgBFUrwru+6RIuNcUXya0
/i4snDSdD2S7qiutYVAEl4C4ITHKmfx0cY9maePBGna5ea7B2/YSeZyAedIRgT0k
WjLggWWJT+8EAxwMp0bqntQinEo/FwcCM595bGOPX815fLcX+w3MMQcFNtZvWyXG
dEIeDaUbRowCYYaWr6/+IiqRPv4qUX1k9lN1Pq3lGT7+l8d5OaQO6mHDVPeTbKP2
u5EAJHD7oAffKXpwm4TZL5+rJn+iRzIyOPog491kfXlSfDF/6wVNj8SJvtikD8OT
BecxZdRKxd2w0IY8FX3bLRA7gJKR2SLu060Et6jLaHC6C0YsolyOMPScvqAUzLny
iXWOVG5ub9Cgi6ePXq0665l4QMTO1IRk3aR3tHO2nNhm0OhhJLWuz4w3ES5zs5pb
tUspmmDB5ZmzAeUsOuJcv3XRuDbTgnl3OEjqEoKgoW/c+IRwJqPRovHKWPxYyXGV
9xFlCgNH6rZCNy7mUOeOD0d+vF3TxxTfpMjFXLDEAh3PVY7GaN2yjH9BUHtWtkQj
RkEhwO838YnplwINaLmDeJJlgB/QW4p2Cq5zJbmwC7eyO4q6yT2Y+nOEChRjHn2J
ptgQUo1/s8e2U3hmG9opEDMXre7ZPTqeYIr+pHfoPKZugczmWpZnBQ80pDDZnEsi
ZTC8/Ab4q3MRy2I+Bu5O5GMIAgl1dm1aEbnk6dWbL3OepXOR7ZNP+qdGEjoqWy6b
JZcvNr/tYKu7cQZeiyDk70Hqys63utFWrXv+wkdOGTCA8AJdHljttLZ/tc5RVUD/
xes5dRilnb4rojz+h+KXoZEsZDE0eAbhbvmW2wohoY7zB912xPs4cH9JiuhVoAJN
N44ZYwRJSbWu3sUIiKLlKJFTKCodUHyaAKItCJR53P4iRYzvdzeb1AvHOMeIIh1H
F3itas1fNWd7SloHwfLUMzhIDrmRk/MWo9rbBdy1t/HZ/DH8/qqPMgT7L/UJxukV
ciV1tVVR37YWb2P15+Zsos0WCI9d1UYc25DDWipW+WwhuWexZ97cuZPdoPl2350W
HuQ2IG465MNQa6yfntmDti+3Z+EiGJ6A7RWJDmfthvWOi7LkT/TcjhLXrVUs3E/c
pW1LaQ+A8PWMWhzL9Zn3H1xZplLi6ieB9YYhxOCV/2M1Lg5dBRPUDIvhSDEK6YPF
/n62gZSo8BYILRFFWAHblZTD65nseWXQ96L+d91ZW/0X1N70EGQ8dnqpP4XFPEGO
/pD6WsGFven/SucRvPGedqOxA02Me4tW1MEvH2+rPIY1wB9dK5rDD/Oo1/NSjRTj
iXRwzKfHKgxsZsQlo3aoTI8SOl/ET+WMRd2nlRIu06XMUqOUlqoX2BbJtTlYythz
Iyf8Vfy6Q+KURbLiobTDhd3xakhjwxIhpWH/07f1rixlBme/0GdnOWZnD6rn7zFh
KplHcTXJkBx0xVL6OezugcuLn4zaeZSZJRwPe/PPlE58wy+bxDvsQNARGV6AnP7B
KsOWvKweCW4nrhIC3otFRm3JVDAWVxz3/ZLlm7ig9WuYxdFN/T8AAnDd6Gn/aCPE
oXn8k92CZE5xG9RG5YUB4olmZp6YKRReRxX/FPlpcBcsldZ2qZdpN7fXBa1C6D7y
6PS5IRdFY0kyywQuer1FBC9pvdFRsL3Ut9MpgPNNjARhO11/i3sddmcyidpmirMF
FjZ2GnnA46GJLqyZDEYxjI6sP+k+omGYdwr4m9zSqi+ql72O3LiLziSPnZkDci/X
IGlTM3QSpL+S7PqmVwKXUOMYZCADAKOCZKfs0RuQrsR9QdSeDqKsBsPwXn/TU6q7
/m12i+PC1VRHGeR6mNU3v5nAA8u/a5QaGO0m8tHd2jMUdfM56Z1elKA9LRAGi32G
+uLYaSk1Z1tQbQVMBY4CsbLXqmqdUjcFsuMVaa9iBjPI9jZvEKO3MuQII2NXl7oc
icpXVUHlQl0ahLGTm1NVBAVIAiAhjwNcZjdHaE1TopkGNZQ/ZyT2/6/1b/QYInnU
yNlUP7QzJofSMiIJV0X+28aKBQA3vMQqXXQ9EVpOgMYwQLOYL5g45+twP23J/ud4
DmJSlI36/ksicjsFV4MywKkFPdIyl0nTzrayQDSLgF68yXPyzNWWWgC3Jg1v8o7I
kJQafwIgN590Ko+qGAG+Y8/0lFAiIHOKl87wCzj2W4908MSCSK4tY4d7TlzGLfD3
ycadwGe2UcD1/iU5WE6DJqTdPdg/f9WPF1IPa2botspTpNBad8/c495+F2MhEjY7
11Prv9J333lofNk5+UO8qHlP7GbgUz01hCpfSbZheWHNxmwaNDd4eP+bERh8Uofq
5i7wCMAa0Vd1AcCjqVHpaimQHtwDjfBgfYGN7OpLeVeYzodQowkGSYVhkhOMQg84
MzTMIEigkhR2Xv7RlF7BLar672sZL3q/RCtTPJObZOJMOPASXy2gwIiqz67t43JR
DmE1kINDxhoYEWy1HphKEznn8Arvxxq1HSISgXRakovsqrmlRDx0AlE6D+yMl+b1
rtAYYnRSMTi+hUTrowEcaRqKPKrt1bFrKQK78bkfCHhROWavIHQKYd4GvnOgCGzB
xE/XVzmHxo0jtht2BMfPWyNmpZoRLV07lKt4vLo6EPYcBScb5xanERLR+goJIwnr
nwDHMe6e3z8JxDXkigOE0RBTgc6VODN/1ZFVsFAeo6+13cz93O53fuQe+3cj1+NS
/yXk30I6Ht/DZnS67j4rvGL8Sx5yhhAaI6bg6Ux5jq43nGyZL/3cz3Gjn2LNnxeC
VfuACJ6EzolHr3Nk+/lwiARjQ/Nu2bsxUYZh0R6gJ1lXlIqMfzbZKtS8h9HURjwW
ZkEs2SiycL7jeYvxc2C8Isbdib+GiRhKkxOnvy/VWGj+UKwiSZ18SkSAqBGKLmNf
F+BR7a8P4Rgg3ebT3M/lLmCfsDeA7NeqcpJq4bueJKBDw5I7VJOl/qg/qRoPT2DF
meIvCoiPU/ClrXLHBJAgBL5EGVpJV2eqbOcwkV6o7uewekvhrZpuXNVu6kw0sGtj
ENxcEkQVjaeeiYN7H+U1ZH1LjlzTScrifg/VBsx57PAnYf4fFLZP0zMaQ4acqKPm
2psFhlh/4RoV70XZmXPa+TKnT4LbcMR1Xs2U+4IgYKVB7FvVP/yy+YhjFIOCuOdw
fampk1+fhuyBxRKKCT03VnnGYVeHes/UAfr5LX0Knr/rwqz0zlGIqq2g07f6YVOp
d7XKZUnrXOcg+R9l2cMHP5c/wtHKRDkgjXtQx/cMIOIl/u0Rqy8AO40dud1Dyr3e
EkvZBtAPYLTsB1wzJt6rHPTNgP8vty2dvuWln3v9Jdf7biMHglw5w3BMCyNaBICU
l/fDgWwN/n78CuBZPXJbupBady8sB1sn8UAYhA1DeTIb0FTCSef+zZVmIuv8/QVh
gV4KUilPpblm3Xs8d/3LWETtc595SnG+3y5Gr9liGLW0qubzGMN0+lw4Y4RBrL3W
EcKtZzrywSPpC53Yt5WHnVHrQiN9UXRGOqOlhpc2i1gidyU19JiNsBXxQw6wlc8i
EF0l1gr0+Lgdq2/NbkoHoYkoWMIc/T6e9HpChE+QBANJiZassgj0S8ivg9XS0ahU
j44WYIavU9WDGfqlc9mwCeZrS5GleCRFoR+1R/nijOA8M49tzef7MeUAkUnanmHp
+qB82wNQ5jBY+LN23Hbsr/Va1RAUocnzrR1LP1mVLcRDqp8GKhPktf7csnJx4I6T
YseTifWxhm0JfSZBLiMlPWNy/1PJ84FujU7wl8c2StF2M0d4Oi9dx5IWkVljak0N
I9AGv6bWc0QXWGTsQ/TGiv/8zLK+eH6g/0Schsj6GiIM31zdkT5iKLL/QSZlzDiF
r/IlrmkPLuYoU+1Cu4tDmIJSYVPGWsmJuto6G/l78j/Fxw65Vc4R6HjCsCjOI9mL
xQTsjBt1Djl5eJBFyUXL2SH3jivvt4T/ldCMyL88XoSSo/4ijFmNvRUYJ//aRvnA
gCiuTL3PcFHiwpH0ucOFWqcdqnj/rvadynDTiGmxlIp+tRDX4e8Y9kCidRHWPCxe
BMjKSkXibExdY60BG1EeAhemhOxbq+nYsAvGF50j7KRQkoA+gO1v/OUeT4eozsHu
Xq+LmWUtZBuFr9n8vFOoP31cl/yJA0zzamcwJxLoqX3MC0L8VP9pc+As44OWLosy
C58Vmte9J9Tzd1ec+HtjGVGy8A3o+7QE3eVjda3YWgG5Vj8e8OG3IWX7OkioLk0X
TQ/cLZgVlyHczeO3zGpnwT0iIswOHfitdsxaDn1tpLyp3lVi/EsAeyAv8ZESbDB3
7LoAH8UqcWMscYkLaTQhI7hXQhOPCRDsLxDXsSBMAOhp5aEs3x6LTaPFNX/hrHM6
xp/XM7Da67urcBuLwXnYdEO+fIPA5yq0l/U5xt5WkoT7m7HWOMRKMgzdVjOp1kq0
nvprlfn4t3WyXQykB1l5cgysqH9p56pdMuxKHWn8GulbzKqiZxNdx1fSEiiZfpmK
PLrg6o3lWZsfg972yKefKoHZf71bsDuDxu3F0osBfYqBQ5uOhBo6XVNsSuJ3uc+b
qgKE42Co0dpVTvaWX2st3sx6BhjlVDJhaScR0VfG+ODNOm4k3aBuLHd2/lGC4ZSV
1ESU3DGPSmeQFUNEt1z6chapC/NwhN609e3e2PBOLwNO9Dq/30vMGX5KklQ6QnMB
VvWLI07rt+Dm1dmJg8peThkanREtVnMj6h7EV9/3CPlhOduJlI3O2OnsZvnWgk+k
YMDz6XiBAc/PMDow3aPD4q0Wr22Gc7oRtFSUSWyUnWLeypGXFy8QaUA5jN4w3jE9
HFezdSQQBbpeg47lhvzc4cqQe2Rf5JGdtew4heffcjsHT56wx+ltBmL+W1YPbmVs
H4CGwADekop2l42uBHzMaK5MXKIi8c0SiS12SCYmiO+HyLTGSEwGvArjMADbPI02
9wzIVoOFPbCr/ML0kzn3yUnrcbnIuWveTPtU3T9kjWZ7TiBnCE29Uo0zcOD8E8N4
lVJiYT9GJpn17gOL9fpfCRcgwMzaSaRt1nNAZWDmdEW7osirteULPNDxn4Q82AFu
XlyAL+QhujoReG7MjTMs5nvPF9gNhflMuLQEr5L5L65FQJt3+KmFk7GMV6aKlyve
FDO3XOXUzpfa43cxY2HfKUaUdRZZ/zm0/OYJpB2ESZ11TP+SFGs3Dk3Z0UY9KA2O
Xh2RRWzIV/UZoPBTFb4PpBz+3VjJgRlIQY3WgaRglVLqd97T/tnIkKqO1Roth6+x
Aq0Dt84G3IEUNNDbEI0fwdHpjNGI9OHekcn88Hg9LPlPY6zxyBcFMwLX0Qxl2Xel
0fwjSVzR4OnCXepEC0e/PH8bD/CYyVfyBUJEpvH2rSrWks/++XFvg6PHE+6dU9H7
M8Gr1g6NAXnTlyJZ8YL8EMooNzJg+XXBRyECimsKoxCXM1y1mGcXu8SAxQqIEdF4
Wqwr3cPLy6rQOibubbhikD478f9xWl6ey2pyyy2r8YM+MKbfhG9LAxnbi9jj+3Cz
00/cqvx1iOW+eqMB0AgpzfVCRQaS9q646DGRJFuqcm38oA6y/h00jG7Lm995mr4e
P0JTQRfp9r5iCMme9oiQaqYIAZW0vBh2cC2LTyMHkR9Gth6NSdHi5YLxOQy8QOrN
FEl89JFjxJvOvNPn4DxvVYGxHTSRuzFrDtb3yFc4xK6mqRQ2lMgjwsDkoIY3DR1n
WPmcHbXyILVX4o/urZ/YGAuXeTKSiT6NULZ89VKHuoQSqMdg/9KXl2m1EPveGkLR
XT5h0H1PVGwmOjp6pHMv3ohEXRRs9DZkje8zMhuoMZfmvL/dpLrUD8COfLI0aMXl
u46CdkRt49kvkbOXgz5W274ABvuzDL8G9sV/xFpY8EVyPXGv/ww5E0lPhDZII9DT
apvVJXs6omSAvxbsVLYTBlP5mqlHvjLpawIwk03qy6YrcR66Zv6hpl9JcFXn9A7c
GlHXvkD3GDRikUDh2iru7W9DAcvK4WbC50fk7J0mc6ljoMWqbFghN39LBPcV9XM3
JHxyIkq7P9rJ68MMbZuOpVLq5DEo7og9OOKM7R6ZD3mucyYo1TjS+jHaX90IhqVB
Zret1PZ+dWACrhDdKG90l1/Ew1jCM3RP4NFeRsjnpdgafQVqcN71DACAYKFFC6du
RncWykYKVCWhWdLUblmRGu986YE/8gGPKMyW9xO6q3gS5nAozzL4nhUkPpJ6W+oO
1VVCQtlWRRJyfTyw+ihrt5MbywMJ/O4STOmQFNkpIynr79UvzkMRrw9tE6aUCrtF
6y1dafllj1+NDR9i/nwtlruPzH79u2QSjYdEN6eWtckeAMYFXb1jMzK6Kpuu9rno
bdOf5Qz3+yBfvYDcBUlFSOvEPYortft+ErA09Cw6iRrwU9KOQArYVf/s03r+XkDa
ez2YlKC8/tkiJl4pArAn6LQPloFwpxzdAZZpUVtZpHtyFqWuVU5GEFGzB4trrGso
3p+A+iSDGlfVj4V77J6RIbpS/+8VzNgZJmXdjSH/uF/LsEq97PxTHkyJxU0HDj4+
D9pCHP/A8QVmuiR1JyhOEpHIfr9sZnS8jdsXc/8F3E/3EYxzqSh4gxWDX/SYdFLF
Ts/MoV3+IYDhR3MmF/0XHVcnNcS6WuWkLfLhGK2S8DoyNtBLDjlfNm6Mt0ZKzFcA
jIWMUaZbLUu+K2kr+ATipvRXr7mhpJGOtkJ+9W27M9eBQLUzNxuW9++4R5Xa0ZDf
5NlrQ6jETNpmObbhOwhMqhR0gWGJTn1GkfuWavuQkaYu/xbNceo3cckemCXjGTYH
k0QF766/6+nEa/nWQ2VYyvGl/+MW1ImHB9eSQ1NnLD5Up02F9MZIrh6N+CE7q/wI
cv6k/YJANIC/xGPZ+dXtrd3v5ei4kRdmESCU4Z7LdALcwUldLWAo8zbIRtOv0OyO
RO8g9g9jNMubwg5ch7+QkmLOKwC/gMO3oj5pw0cD1Gcyzwr9vyXenseOHUFJ66BE
995s8+beAaq0oSS1LOKLRhKB2Jzl6DabL6F5HOu33EhMCaGB3sHfNA0wQq1EO4Ua
zPMaBNB/3k3LBOhP4GnxficHmsUrGe0ym1BZ9MgSV/U+i5D6UsqKZP810TBlFTnZ
vDyfpleaTWMVKNtqsAZOU1gS6k3RfDOA6DDDQzbnpiLvHui4V1IsbVAFaTs2PF+l
Pi69iFmW3mmjStMJFDWDL4DYgcTIkNsPhNk5fBp7nuF9zukzSq2kI4nanavZNfj7
mqKY+POnLrrTpc7DS2ocuKk3xGgk0TZP1Y4InPxzwHtbztU2d0UEa1Gd2K8J8Bpx
DwBnCIqXDdHS/D41vxGJJuZx4a6TyVqrulxcUWf+d+mFFTDyk09Yt1+D9BfVrk4q
z7DXZf7lpjDVG9U3PnXSr+iqypcpZcEbGveEKaqiJHVt0mWNLG0usfko10QlkxIc
LWm4LvZYcLNgbjbPNqV1pKKHcOBdDh6zQfM+C5nhZ1FZF6xRMnHj7DU3ZW0Oeicm
wd4fMqEAxrpjl1Qu/HJgaEPpFbFr7m/OFWo8UVXmNL9tvvMec1rdOblfrzn+Pked
UiBrIR/wGIE3vI5gr/6DEC0OgDzb8cB96qeG6g/0XtAAKb0k9fhNuUPRVPQUI1Uu
RPfdUPX+kBZpvCil/ZFRnky0jTs37VJcVV53jzUyHrfYhBTdSrY5yfrnMTIkNzk4
zxUHyG60QgYVpbRSWAjhqE2jiVJz3AwmHEHmfkhiI7vqoQIkhtystIZofc6uM+bh
vvv9+Y8/IxQPY9bIxWE5gPNpEb3yRiuhMMWB/G9iFbOFcA6JLJtBa4okESoo+a/l
6LNH6/tuz8EbQfjslbrJdUNwmw1C34Tc4yQGUiTH6WWIYPCg9S4tIbhM5hv8t9pB
qN9yD2ST8RTzRP5hi5+DhEffTsGUgx8HxApak0/QTlIQasLKkIsskY5UIZnI3GuF
gIaVDOW/RjNwmkQS79aV87/Z6wW2xR9rXO4A9EA80R7UyoTZp+kb0PoGoUMFULcd
uQ2KSg7jGG+CJaCFXk67ysYSxOqGSW3y0DvqU/5yxwfqBzGUNtadboBZuvdD13VJ
ec98+TJgDhX8i/Fd8yq3vP4FEPCnhGmbri0iAXxrYFkAMY5blFMpzU/orenZ5dX7
It7KlWbqvSnu8/UghNGQMPFWGP+XZVpoYN26zeurd2f8f6mgwKGXe0IvpiBhTU1N
RYffk/hlM/JPCIw9UwmlfJHm+Zbqlnlore/F4klnPpBXeJZQYf4pS2Hxkqpxj++q
gwd5v3UOK+2L4WemArgeIVb1FeB/2OQSPbVJw3mcF0GQksk6k7QxLPsVU+ukwS9T
wrzOhyToMxeUCfhph6zqJwLeF8SYaxa8j3I4zwLfYiBbD8kEJdFjFLkK5rlbf5Oy
ByOQu/LoEmIKqb4qOz0+5wVi79wsdWynmGlgRhppLMGsKdThKUCDmk8x3oNsSnpL
hHH5m4jmj6KzoDuwsYH0AzvK4dEEfu14k/igM1chHBxxGHm/ierrY+QJV5COz8aU
2fOG6PDkoeD2xW5G3pD6+0afr396CYnmp4jiU2xNPkJK7vjPtK0v1GlFwmMXax2J
MSHxa81osupr6ZIUflvT4iTwEg2RoyZDqKM7bRXVvHSPeNbHZqKTf3gdX/qkMzzx
tpQZOUyNwY8MV0B5TJfNqgySU0+ElbtkJaoqMyd3TnIUvPe4dN0nQpJPTRq3kwhC
RzEFwsOHHHi9/rWWPOrMnXHwkY0m7dpSJDcCJ/UOCB/eGn1/8V9ZLcbVw8d6/jtj
h5KcyWQLl39dKtHHixWFkUP//BQDjdh4JGewgWYhV2ShJ1srpzA1hU8qJFxRdlJe
fHPujsrKiznnsZ45Mi9vklfSxZUoCMAtodwlx+pRXtE01I4tgYSJ1kIvIhhqf/bF
oCsLlF/85AnX2P4xemSr/gE+7gBA4BLMKjZ//UE1t6Xo1NGZl0lfrzRmrWHSOVXS
cu+9RVJaThHl+Ct4vxyEuH+BAC60/kpctn2ZcyoNtwNH0SjpJqSZVVlS7nEewaY6
TbP4HxXrHrFNoiuVkG/8tNagJP9vIV0TZPk7VcuDXNoAx+emW0jkr/uuwfOf1E9J
AcE5b9CijLEWOe88ojHeo1wa5OfebNMHJzO6xfsGBX/U1fsh5iOfd7YP9/GXhAII
TavuA2oc9ENr2PHgpQ9vlpdfQSbxPkhGGOPjBHiofsdJwBtWNOEvNwvq+HbfYFoi
7SVroWQuYqY1jnHNJ1HT4kHCb8e78hABQHQzLjXPQN4HzGaoDGjs2fgZJ+MAvJEQ
iZjgbbCMQFZ1Pi3Zw8bNch/qdyaq+1oinBozxxvDlj8nHRguQR8mbOgDfrPSjmes
RHxBEu4HQsmwL4J3Pi22KuuBcBNMlOEClIPakBg0x7KL3EckDj2uovnlkAAZL9a3
LemLcV5W7wEoHURVl8i4t9Q33mCathmA927Gcn+uZi3Xu1BLwzlgn/paxxBra6XQ
EIHydRjvh7WvbRePXK/+fTfsevzwic2fxqdQZRB3XwCuGcvlpwmlR+J3pKdH8e7Y
Eohf2rjeY7cQWrCvURNecaMMsYmQfgqc59YCz5F3M0YuOzeGU6DLbnWVT5Udi+35
EYhSVg5i9N1/G7rs+gY8RXEtzIiWtiSEz5dQTfwBmCXiBPRy4THD8HmAl87NNt/k
RpzISiyd/hw0CudKS9ZMcwLFrQht+EwYRGnLd6Bt5WOfYY4HfrJuVIQvaNARFsO7
ttwAsFVNvDjwUS+TVCXAgHTkCTS74+hHZtYzuRisSZsrCHpx90PTn24cXvPP2P9h
PThROfrIeMmr8uY/2vtMfPf0rcfwU6JlOcdvPww+Kglr9lP+htvu94CsZEenODyN
m8xDMQA/0gbDYL+2v94mgQ1J+jZnNWkHWlLNZJMLJ+NgtBygFdo8QqJIvE0xV5Sx
Uc18Q7tJjh+30vxXjSJfyuEXgMy24lw8DytJCjRyNICxe44RStwJ6tTy9Mcuv2Wk
6cozDpi7THNeDS7n3IrCs+qS/JstuLy+KYHzB51EAYjsQD6wFvjfpT/76J5q+oUO
O0NJO/K0P3LoQGy+ykazEsScm4k+CQ2ZHRXvTHs1ma5lDWBK7Nu0mjhrkDzNmorZ
zl/RvfuvYKgpzdJ8NgErynfhGfaT3HwVlyEuC9/94Cor1WpR8XR+SRyoIjbcxZsZ
nJT6EaRr4YV/zJLV/VIzwEGpAHYeUtoX8Q39bAG/hwXEnV7NvCN28Ioz5uNY0iKx
Zhtoi/s9igN+LP53Dr3OcJr6jyRmWBuIARVI47LwkZIGmJD4PUeWGMfWErWsv2bD
+AkMcjLBStkPkvi52JqyubRyPTUtq32TO6Zb3q89bfaf2noHdfeu0Qf0YZi9BmjV
srz/iN/ksEpzCkcCDkr57ixzuqMvieHCvV9qNG0b7IM+sr6UMVy1ekwe3lZyR+J2
NRwcXUWoAV74Y9PgVk6j0DGiIQSrU3PN8U2WDI6HAp9FP8bOtxSg7JByvmLEfGED
m+8IosYGz0Afmfmq/4q+1yYSr4LYzjuZPWn67pHGaDcNulmxSRkTfJMtTFefdnX7
bO5esflG6k65QPD61zKQ1ihRkIewOacECGg5MleNnPS/LZSe3nJ7O569LavexBhg
ez0u5NBrzGfNurI7VB7wEvL9hABeckt5hTE+UoYLrxAs2PXwKuPtOeBGV2yvI4wJ
tvYqHy9tHiELJS0BgbcTR1KzVhErn0JVb+jgTQE0ium7Yetq4AsEqsV8a1xJcFG1
nX78Uhb0I+tWfuKOQThMflK6UFmUo6mRU1ySvQvDdLxxguWi7TuH2AWxr+4wvbt4
A2EVhVpTkOLGFZKSr5dqeVxYjr22u7AnxiW8wczJInd750ZyXO1rTdldE//Lsga6
RomQ/Ihzr0jf+7isg0VxURG/weMWJ7IV58H2dlX6YtAWYX+hyWG6OR99QriC7WZG
6/1YPss5IPVoNAftnVfPk4BPswSI5sCsnlgfoZ487QP54Pn7+7v+gKXN/8Usf52M
BzYvFbzf0gOo8iUt3cjWmTdQL1eUlNqv5SRipzcgk9S1GillzTrrFAZs+1KgYS1M
5Qk2ELVjGGIiY/JJjqrchRxQnBEcMgm0N674S4sVJvKRQkHObxoZEU03kVyxVOEt
sxEQUUj9fyZEGwLSNzEu1CowvU0At/7SgQrMS7cfngv35WHXcxacN/Ahi1zf4FtD
UtnPLuISqB9cqq61h386OBSi0kNEIm2+aUus4DyfNhTrHc4/DsQyWqcKeRiUk8fA
DLHxN2ySGreQYQIFLm2Cl/D4QCYckGuHhO8Eh2YJzFaqI1LWqFIQV59xtoth1/09
P0kS+Fh91h4SqVDPysKX5aGqIZU4Atq7MJdL0ijYZRR7zKk7E6mIw75MQRlgU1eA
EEu10+ekZOi38fZhLACn1iTSVEG84z4lwzfb930e3LpJJwY0mbJJXNrQhr7m/9nI
1DgYOZvol6jBbzihnq2p+PvbADAMZOkdcasQDRxxBL+jJ88U9Q8XhG2DK1qKHnKs
QDzxb3zchfuIfzs3XugJyvaYkuLxSVX/e0X+/ZrVHeGVwTFyPpyYyBXQlEm6deqs
s1lBoC1YBGem5ybqU8c2tTJ1iTs0oNqAuvMj8vTTuXK0CReGIMOzghVB4dcZY7rP
S0t9LSFfT+sEAwQea+TMUEr+SXC1vrW1elawWbDLkQfOctsVidxaYWCgLwXtiF5e
kyqx9NO+IhTvaef8NdTBx84/tUZeX0z3hJn8+L9PqNbksBwfwNbuED3Y+0sHbB5g
r9YqGm0iU8J2BlQY3slSn6AnkLB7qYwapWbFZCDgHh0WeenUiTbsg38oCU3m8qyz
R6D9L8ZQjY/Y7Gb/zJg+NJeaGSnEGgsbHoQngpWWAO/8reEa8eVQmeXV9zp8kBGb
Beqth4+cDgxv4M9g4cig62dtyGf4/PhCO7yf+QQsvgD3WSRHBYhMrjZvKLz7kRgO
gucj1SpBXhiVLZIA4VwPfIXzVdraTTf9YdTHb0bZRrl+yeJJteOQhLC4hkFNb0bG
bDquifcTwhq6+hCjug/lDn5b8EzplGWGhvbJzspH8me7Mqz3LW7/aVZ2r83RUmyg
6bYdCj2cSvP+gWRSZixYRDTGOLmKQMZNfwIqarM4mUK0DT9GjPP50hs5btFy37YE
w2Nkl7QDQRuH0C5+D6HIG4AOxhLGrVTDzuhQ7oY+AiEfvpmTRvroGRyj+gEaILbz
X9WHXZcnwH9wUghCwCmDSBjV/X3BmlpPwH8Jv2r4AeLCkb4Iq7R096j9vPfglHT+
wLy6d/uPl1XFbCPlJB3Kg3juSXQOWhuo+i1iBuQoOxIXqFTd1qaXGZa51uun99OU
7CWjK/tiGc7VxGSRYRDs9UkMumLXA1Zcn4h7DnDinIXeew/bdgt1CTq1olpmBN9C
ZLLQif7SAkt2ayT0Mn0w26zgps6ItqTy6RTasagFYrDfB+LEoz8WcVgCsWRpjbHR
xxQU/tDM+FBKj7tennJ25ZayMkMB+1mZsc6pnhbrDT1fL3R6kyWTohvIJn2wBZ8g
smH9XtXR0dD5NC8BH4Axw+f0pXr0Nni+Vyd0ocJi9e5pZYVEbLJw+av2c7ZFwo2o
GyeZhPEpcEfpYSKE7kGg435k819U2zovq6ucz3eW8iXdDg7F1wQI7ymSTCDxhvqp
zSNO82111qagZd7oWvRPfGS4mHD5JaQbe5zL3JAp4jVJ5C1j2e4uKZjCLycp2llJ
iODZ0Fsxt+0wymh/AXvS26hzgpTWKDRlsc2zWJjKbROS8MAf2IyhWesFYSVZo3pj
HKa4+jdBxniV/OJEw7IrLV7RxwrQQ5tx+C09jKvnBAPDzXwUET0/loci8Ca/v8G8
TC5PGPgKODqHF4xumm9UzuiQSjiK7KDZw0cro9Q6zDo7VZy+15t1mal12QOvYJG8
ac1mIByIaS9+D/WvrLxyEJ05FC0c4ARqFEVjzp9eUgOMaP1DqpdwMYCAJMQfJVHc
Y68V6pW0b/LgQrAYdWbMBb1SH9reliBPcpEAyYbxSeNUMvPRvnjSacQcHow5syXN
b/kB5u/Zi/pcBge9eOvsLoB6dlIntwHT6JsSrzMQ5futgleqhoO9qzWzqLtlitCK
y6z7H6yPC1fUqosnZYwMUqvhH+79XiITQP2jWTYyfIWgW1HAUeacJHSItM9OUczm
sHYXKKvwO2PwWM9tYPFf1Zlkva+bBCDqTaxq22Zv8Bo/RH+dDCnpJxPhbgSh8HEG
75sUqQrNg9Fh7GRFtIoI5GZmWENepMpdwOPThsbL9R8w4w3Quf63W6LQF0MncV/T
aireNUfONkKoQmrv5Ant1OZEkcvYQTzSdX7mvv8irVbsGDPYerclwi+S65tV1tWF
R/bfIz4RuvgDrI7Ql5VNnHgRe7Q0gQD6oAUaXmBDf0chPf+DQAfHFhdy5nLuSzZF
tZ6pTkxEOZLUPpm/lxbjXikVDEC4KeuQhIaA2NdCfP+2pyCMruE5AvOUfO/JXHib
XPOW1C5LaLTmnmjhmnLpchg4F6SmIjeOhHe5yvU35Sn8kIRjzsn5SOX/k/k8Tt57
1x0/xYNIuk4lKAy4g4rmwoJuHhxdfbWca4fYcIjvBRwyR8hE7wF3pcvwKmk/krPr
NwWy5AEtTDw4vhudLtANnyEZNBTHBPGA2/NgtZEgXGlVq5HaQ4JQepbzRISLF1et
Cw7mvsruAUZRdH6NtaOMIPHZf5KzOv8xhN5ppgnTkAUGKgAtpARQKupo9WgEacOz
Q3Uf48NWCbD28w9+Kd2XX4eT7RoZaCSoViAF2cXY1jl1coJ3dU02Il7LmjjzpbA9
Pu363ZdUVucMz90Mncgn/fWOd3PfPbq4Oa4LdQ5E+9pSE0DKoaQh00oB4NrBMZfu
7NbGIgUkzTFz+HBm8t+G98p5Mn3jcHyp5i2jcUTWoKt5BTX8ho9ttSpBiAufViAB
j9T8FIdI3Tm600spWf4g0Nllyx1Ged1Z9zD6Ry38Pzi16yS8HXbjt8vJFPy/IA36
P5S5SYTMrAhCZ/45qrUDbQub0v8sWAQKJb9uH+4cW/WWfGDM4ViiPtS/PAfAAG8F
36EToZFWmTqC4+ZtzNkaVDT0t1Zc7nv6zIH8ncu1nJDT675lP7XHHKBxmbln49mw
LHIhCYKhqX6G8JgNU17/V+CqrVCJRIOL/n9gClGLIw9UMI25jb8vjQQ9qFc0LG/9
Lb7NmDWFodKKNhkb2ZhI6s38k2q3NbYct3YkCiapKYCLS2Veduq+pw98+kmuSYV+
sVLmkAsJMa/DaCwCgZIDc16MuqDzqi/HfBXSFBAvgi0NmJ8qOK4pHWaCj/pW1gvt
NkaTF+Hyl6nNTamvR2C8+HKkkDiavNw3DgwKdX+Cjn2Hh/4yHF4CrQO55v+toRf7
/gd3tXr5RfFWFuT7hRdIm6jJjlRbzaZQAaaeHbPsaeljnqTCsKJIHnKPh3b7c/HO
CPL669XcDpFZwbN2/hjU5DmLBVDY5f2aPqZUb2+LTB3LTm7QRJFJZ489etsOGY3n
aTm8mKIOPYLI1Y0GVPKtlSsX5sGlq2ilD5AGMR8JGJcO0yY5PWLHyxmlFOFj5frV
KMcEC4rcKOlaf+Sv3zVUj98H/sD/wx1rS+xw+ocsaBiAsUrai2cwKigIb6ZLCEYv
AQ2WbBUnczPCv+D+pg1OdBLicijftZ8EOszi46npVnk9VRImdtscT7sB2Qlcq5H9
1JV4NDdotIyYWg8BumxPbEF8IFSptPI2KGPNcFUH3FcNYLXRw4oMmuPxkBSf8gKP
kvMO/lIVttKz1cpohOrnE+YMzoBxy3dN5ReNxdQgaDen8mC1WivU5aCQ+c1EGX/o
mkpWJv3Cb0hZ8IVrUidPxx68lg9v2e78xzYIeY76QVqBeWDb2TUVxk2WGl8KusOP
QrN8r4tsD0c5CwdpWhu1O9ovjEAeeTgC4avXkuM3FKKrgboDts5c30TCQp1ebboE
gqzSVB43H92VwbyXGco+8bNZc76vsj9LGzioMwiujTPIZynItuqswPCnv+ruFojf
IXCDPJ+cbB5bJ+2VS4djA5aydjtzHdV97LuYG5gND3PoE1bVrRZIPqAKeA2XJy+L
8GpQ/ItV6w3tdnDwRxCWfoPSJC2m6JUKyhbeC53LNxOOGmRbUaoqXO+8DI1CYe1n
VwCtONKYgiYF8F7NGiZKuNv1aX7RIyl94q4sYb7J+I6+8DbEgwSm6k2xaxfPa17f
Eb7siNYu3UC8b0XcQmEzv9xl0EBVf3BrPzjAhlHxKFta3jjiQdDLzCyl38FmdQEh
2sLPO44ACjkgtsRXOURV++BNp6sd8D9nDpxkondR9YB4G+Oa+p5JXeYazoi+5PFe
cPk8BHCslZAKSCtGjS0a1Nyx3wyHzaGQzYSE9zV3R3nI8awtzsxR2pR6kL8tWSEr
sWUbgO7jWwoWovvUT64JtQh+01S3LZMSPBp5KDGQ8YHYXdTS1GmDtGqloSHCKr2b
OGwbInDHBvg24Vn8IdHIzZyYT352IT+2uJ7iNkg3edjbfGZ2Xut+U/BXPbSjy6Hp
r5NfO3WYrAAy3aVcVB9OVI5aTQiyriyj2FfAENfiHccLjev/OjdjmYFvzPq5XUq/
djbhZMlhNpcXPiMy3TcY0bzHVdG/4W5RxS/+xND1H9+KDxtyvM/oMH3ydagTZeer
tSUr8H7uhHcU8cHBcXCOo+NVT7NH54ZvjQghdjGhYPaG18ODuK5hTeu/Ayuo56oO
KNzIgZbqEby7GwRdk+mLHQB8wkwBUWTjZC/1qjucyjnP3Kg5YCnhrPR91YWMznis
GcDMoiOtARFSpD2vp70uJxPMWEUenIlnLVeSQK+j3D+EEx+ZTMFk/4sUQGn26V3y
eRh1xUFVPUB7F2ngh0mWnGuE2eTgCjbVQET8ZF1XtomqXeqGL+if1V7L5Nk+846C
kdPxPeD5nEGPaz390gQgQ9TH9gGMyL5SESc2egs/6Q4X/aSVvmQ8ym51rJ/nqq2h
KNaocmCSKao/GDxq8yzO1T7i9rhD1RSwl5wDV3f7jH2WBXyKNtkQtPp785hTPIio
LpEiOgam506qSP75n1E/liMP6G5PQs2zxaWUz3MNa3vCfWn+ZVbSxZXK54MWVmCJ
pP+48uVqDCdRsM4W9ZstssVnR7OlaHbTv9+Lb469U/qKMvQiwMYlWX4fEBWHnlYN
JB6P7cGUrIm5NlZB9F8dn+65ty+daJMYgIH6Fala8PO4QIpSHc6UNWTDF37j+8en
FeJD/Xg6Zrs13GqsevmTdxxNtJzh4trFaoN/M9dSjfUCMARAD1tBOHBalIeG4wyx
Q2PuErVVNEXIdOoKNq+L2tKky8VWcjdKUU2N9Y0UQE9qHyJHMJ+Jso/RpavA0yYy
CPvuw3Q1J4HGCyCIRJjzNcx7TkMmJPLSFsbaHQxAV9oKhAkbVlnmnAWnYEJ1c1/K
v/8duzRnESHgrml4+uXRrcge8Ph9ubWn65NTKkcja+zsvDyccwYF7iHkDPq3TiaW
cdAQ+yVi1gMt83zuS5+oaoSjRK+x0L+9jS0mz1ILmwwuWrZoBwqj1ZCwGhsbCLB9
Q0NCau3Q1yxus9WaxspNu2l2V5NSsgVxkbPMF/mKDG/qflT8xZMi+NyZtt+juqyE
fnVNLk+yqsKoG+ajdOqrvbQNM27g/QBcM7FoYtI+dGdAuC25cZwDOEJsMLwnF3n7
ajPVi3hDrRT1RzAlT6nmY7Ghg70Z8TmHblYgbOx+ki7XIb4oAaTAHccK89ZuYdx6
W8XFDXZxCmQ7C24AK/K1z0EnkUCxE8VBdoG+zeZl4eEXizuhb/9trQpZSU9qB73q
s8M3VPvUmyyyymH9HGI+DW3pzWMu9QE6N2zPhyfdKujaNFr/FiBWfbDq40/d5zoa
qgiRisJA33eRDqAzlwY8kCPrW4BPhBXzNX4ne2r2lT5NXonzWOJ7iDavCC5MqFGg
52jiCTCNCw8aVXNWiH9PwkGv3Ksct1iyrdFIru77P1MUsMdUf2cW0wxJjj1Mrykm
Vu1i8hMEFTFA4pcGp12DqA9RhkawS2pSPAOSceZn34sdq//0B+CIkSMTKplww/mx
QKIiV/ZyZSzQyIU9toKywJ4DVBx+Mo5XVFvQRCGi+c2IqgIP+G3lC+vO5Ahf+WTv
2RXWzp9TSuq0l+MGtrxq9w8KYA+2lipNmQX5BGaocrV6PMKLbxRRfx8wBda5XBhC
EtpbXGXWBRWyjcAfknIkHbJ5ByAKpybaK/QVSqmL8WJ4cKE/BvkkJVvcOzBSj/W6
JO9siRfaUWgVp2DydG9ZChA3K8XLbPwKHFkx0Yv55nN7Lr68jPbUnGRsEX8PwZdM
R3oWhbe3FT+CblRLfrcEj/wpxjTx0Y2S4mQDofAZD5JOtpHPtL5wcb8eRM+6LeV5
Dif/jbHJsHE9t2o1+xuUzR14KhmgqjiKkPXmhJcc6d6ib4jC0cVG0JeM0CY29opn
9yJxP+SDxvrrjL2kZVRUTCFWUuH5jM2Dtd5kVoTW9gPv2kAaImaXexHWz6PPZPFU
znlyHFqhjWFuiP+cq2tOvNUtfMeWM2ksvhSKXB0fg4XAMCKO3VhdyJhHR1Pxx0BQ
WnWZmW87RBkXm8u/Ko26s5raL+FlLBlwXuk2BYiSoFB5Gn8XqLunyRO/JOfZJzNq
HEdovqlMopAgxKFsQ9IxNUcj4/6QoyijBhrv2s7ll31PtARTvBmW6OthWS8Zb/Of
jX7q9qCB7rEXZMpghWAacLGSckWmw7cCyMi4F7cfq7sCRSWoexoSFURXz9visfQm
x62C/ZDxSfzNe9+B/PuEvojDRRLrgz7s3/kl/Et2mtTZvQmZoL7qZ02ulPe0c7Rc
ru4658L+D2j682CmJNUjsO+yEzlvdpPYu26YlZ364KkYViql5ooA+On3jrMBhCsC
pb9K15cke8TiWYs2ir9IGMMpsq3in7dzE3PoYs7KAG7yqgU3N9xUiXOfuAamFUfH
sw8YZ1PD95flVDAUYOlaryMt7vs+NYwapzBL5fusDhmNtfwKOL11BpDArirk1fw1
/KDX8z2r9oISMEZ5q61uvvexDXcqATRE5prvlA/ElWk5ak/mhp8VxxN4aHaWWZ9E
0PW65L4IzSAsWl/Omc7nWp1iixGgUN9znBDpl7ZtiOZYAKBtPQIRSk48gx1pQ61m
txsv3YNHiP5jZ4x0/9NAbBIMOWw12nR9Rp2zjoFVkeah3WsnZXs/z/YNKKVp1WRq
gKQVNo2u9EGabomJ8TWGnGUKr9atfG7ZNBS5HE8PpI4HJEMNlZ/ZwLItZ7CTNAuv
6OSOQTFa2J1s+RXQr1tRW1wUke6ATTt5p9Kn1LpoujUBy4BLGuaIOMO35pSDKSH8
YlmEBUsDW0TtAakykVVW4JHs8oW1gITX3YyIPYXZL9IhcHeb+i4Hoq58IVEN8d0V
cTRpvRb5as4ddhHbtLmQztzJ5xUzI4j16ccISkO8fvAUxTqxiXNS6qk/K7TT1uKu
fYSQ6GgLxPc7FIz5pH8pEx3Law0e44MQl9jd/u69miz+zy83F091FqKGv0kP0zKj
0JA6JRgun/tdcGzdyEW2IDruQy2a6hFOfveW/OZBSrrlOhqoI0xM5n/1PT3Sj/af
EHUfuliX/QN2ROx/zdPcRYZoZp4Q0zIDvDC8g2SF5sGH4SSyfBMaCiGX1aWCUl3Q
z4UI5bsKwU+otkF6DJrb41x3aEXtQHuKyBW832RbREMsU87Mj48MlRDoMcL0D+qc
JNrdJvvT/14aa1zjg4ZJBY0yR1FMDGEDqKgVNSS3DmKfGun9SIDiIByUodn7Ga5f
GFpztn8gQiSXM/9CUzO7woKaXdzWV8k00RZ4QROZCwuFxvJegF9Jq8qw2RjHYwet
h3qHNvir9i7ovatPriGETgbQEAxqw68UGcqA9KByUhx0JxSS1A9g0BznZJ7IkK69
Di828BMPMZXPeuGNqgQw8WmyVSmqDAHLPBOUyp/WY9X+OOohBOp+eFoI8ePDkatK
JcFLHmvDC69BsrB6/Bz+zz7Meq9/lcvxPRTlPGQhk1LRD6hLM45S7Wjsyay1W1du
mj0IGZX5JcqAz2ClPMgrKzgOzSEmcCqdLR+v8aJBzfbR6wVXv/3ITXpQp4+7XXyR
hpwuWvtkIeZHCWcRl5L3MHcAwKwXOajb7HIhIwpal7SxzXHfk0wbDzysOMtYj8CM
Lb1d0uOSJMJg7iqndhIglpHAerqZuVHAY5Ky4rY9RIJ7lmutlixoe8UFnUXm2tyE
S7FBVs4ET3Ne6sjZewCfbsDTQL82I6aO3LwQ4Z49hT//mZt2Nd6peOZGT9sFFtiw
Id25umTmegpCx/cL4H33v/Mfa1HLny9fPr7E7Few6hvWnWYMYt1wmB7ma/AX1rrO
hutgU+Lx3i4E4cjQ9ugGp8k4nMmAof65FEHe+KYFhNufP1nXsvPZB1DVbrb0QJN8
crbM1BQ98mVevS6jTXumas6piO9AHVSVofwNYf9WA+02w36VuEnn5DIjDbPyKvzz
vFpn3udbOA/hmhVyZ8DQLKvdmNkImltaPBJZP584MBfhXXm+4pLrx4MTFq5gNa9X
Yqe29oSeF2gUX9KrwSLIqLQKlJmQlqoNtknQxN1MnAeLYQEnBVNluBiq7ETQ7Qov
6OzJkZxIuh9ByxsBZsAYF9BzRpCU3l5+eS+CMd1ucX9wnNsF9iRr2n6Jn94zQ0X3
4O1QFNUk1z0We0ZfO6D9ZsoEvkpho7CEteR22NQmqdmbvqPSV+HZ/kacGpMTUI8+
YSyzb/vk0VDIL42gJORqz4c76cDroLj+1zoKXOZQssLSeN996a4BKesAKrlQ0Rv0
AAQrOpvPZkTyKEjN4TnYAmAWVtUbNR/Frv6GFyGdwW6Wx4zlFZSkAAMZg34bEXPU
f4mjE8w859X+v/iCuhTMnc5TrlHoHJJWYuX/4wGPmNi2HSoN7P+eSsKprfGtaSMI
cbQbapBf3zT3Fn03oQdFoAJ4JHBkcgTDyl6po/XE24WkOLfWT4qpZiFA7fPuiKWf
OKkbY6AMUbxqJMKgjfy0mRdf+c8sLKX1in3eR5C79h9fFQWlS2nTNplhf5rwUfdc
+K/ncJLImulI3JC3yLcylUQeIrxU9qqavqVX3hGbqYj322F4etEh8spw7vou3Iqb
S0L9bhSvVV7s6oyfb0VDy52tmpKLlnU3ONkZhutBuDfb77HypFdqqWadVwGL/Fxz
ewo4BVCVsFJNuYzHLZHC4Ss6QCnxm4tTXTa5NXEO/HsXJd7Cw2Pj60VJAosMPB1c
othKBOx0BQ15FraYan/+MzOIDDGB1rzE/ckDUZ4ydTIOz8EYLAevaA/l4KqsGB06
f7P9zXjn0v0OCnTHfAxKd9SiPjjE28C0KBlNsd0ZHDj96zwPEwhAsevqXpV9jGkg
LdOkQCqgAebOyoN4paMuJKOWieEoOSC9ICPXhWHhcnImOzpnC4/byl85l2ZbtWmi
usR3VMz9AQWNOi0w9HWTuK/B8ud6bKYyHYg86+Bz1ruiY/uBnxRG4SAnbOBxplzJ
54pVZkkdgOBH9x3qmSFbZXxlA3sLvw4aoxlwDVLTdZoO/OwseXvQ+4NN0dA57NVv
wtiEGQ6vilG784LnJjN3tA4DbqA91TF7m8el4WjjzalnR7Ht65wGzxGKQKMiG//K
PGLR6TjjlQwDMHAWDwR5Xwxjxe8TqlAo4srwO2y2iGBtoD/AZUuT6yQpXUHCUcve
8gyMDTWXKNo6YFfAfpm2MnwlMsjsycaq5lhdHKSITWz/u6hGsGOPdyZ2KSvTM2/g
tVWYi0PjClUYTddfZMLLvWBQf0LupVlndID23cctrwVXbU1Vhhks8Zrq9Diivyd4
w44wgkVRjDm6ftfq7cFPsEJSMK4jyGTVZoK+/VHqV4rZv8zxxj8MIZvKLuJqSmyf
lxS0iE0+otu7ea3eWXsA5VAArmYUb0OvjJOJTqJzVSaz0K0zE5tW9A891y4teWo/
+3LxLCC9Kg2v4Iqz9MIYQzVMXtCBP4lkdrs9+oHybEFNxOqbfqs2iJ/5EMZ+Xabk
6K8XMkibcbalEBjmZel+/dMtukNp+WhrIVDGjAh/LfXYx/xOQjLWvlE5LVFtb8KO
9FOqSceY9TWQoiUEs966/xXV7PJe+sMuMd3X1glJBp23IdTP1+Pee3NrHinRTXqJ
hXOtRnFNZM90y7lN03ytsD4TY9EuVwJbuh3z8tGs/EtPB4dgk4hEPn+GToo0e+4H
eub7lUYp28jywmwqd5KwT2itClUc2HmkMRu17W2hWbDPiu/FUmCMdIMI8AQaBZQS
mramEy5a6AfzTLwf9Q5kP5aWDsxFP6zglgxUgjeZciz2xCsHhkrpvKYauTG80bpo
pHUIWGlfrEFKBR+g1js4ApAM/Q9e38skovzBCE2WygEhO59f0MB0AnE2fqj6gK0B
OXOjchhlDqif772Vpf1kfM/2l8dj57e5bBJTfyRpGTJw0+HesIgh2giKCIsOwHcM
NP58N+xp8TG3IQ7QmK+sF/DQvpAqbUx80KcMsNUaJJxkfRiL+b+bTOLAehh/7Te5
P+fRsCEJISC33fwlXpE62vFMIzMoM1bRVwZ3LDooBbl9uNN3hYsiOikwBU/JzjSq
00VDdKA1N9qlGc6/efN+NB2eCo+ieNcTBxWg/RYyUaJ0FNPglTiYb8dS5dfnaG9/
pB4oAMIs/gfztYhMwzlTqbxABowMudVIw4cbiLpugV0nCi4v5EgCMLUPhmSLBRaD
FUmo1aznRK8kL4s1WsCYwrDKXOiJQVjjz3+xpkmX9dG3O01txpk1kXHFWgIUePng
EWr3pVEExi9OSFVzFnCGP4WVKggBGyM86rMKrwOM0Y7IFgY9rcmtYjgezQdmuYjo
SzhiqkQlhR0nDw/HESb1QqtoZLspB7aH1bo6Mg9Ac8dz/WASIwXRIBVYYfNQCFcp
QmI353w7VOo+ntLCUVm34MYNQ9iDfQXWKCa5q6op7msZqGDF1ubCGTcQ3AD9d9Y9
BhusktQcPoK6smAMr6S/szJ47YGfEtRSYepUS9kEcBVU1pv6g0r0t4KbVADwaglK
miMwLUzuyvK7UbmVTW5P1TNZqaUrbRpPIBrCY2oHZ9rdWnoM6mKzd7reHwpClPc6
pGn5SHvOboaGbOGLvu6O7W9cxpYjSwt69RNfBWbiqQF9wHtw+akhZazQil7HEs9X
q74EiV9I7M8/XUkfcQrwizR14z7n6dIQlqx814uxOToQPY84DBA2KVK/jWa19SPI
apVSQ7WK/IXlo7LtmsVtsbtv+kDWSAtimPZAlxMDTrGPtUYEIa+quXDJBdYvqWMO
cDjy0YogoKtyXgBznfiAqaPYO3c+MYwWRGw+zDRW4TFDoDkdVv/B8ILDCTu1juHF
IKbRhuAvxqpEodagqJ5V5cJ5svKGTs8tkoDsq8Dp3dFiCPb1a4ORyBd3gWrQHK4N
W8PevL/Lr8u1wTOQvPQGA9QjAHv8BE2fWyyVIk5ocA0rzOdouBHmLvJ/qS9OIb5a
gXdiW0cCDL8tfOiR27/mqCdE0wzaO1FP58tD392KhCnWcQRGyuU4fY2agRZ/4kFS
do9v7ruAhFYoiOS7dxJLZB3NzZgK2RD+7u6k3XP0r/8YlKz84s034Bi40eIPKByL
e8XfMIHT1Qu4qjj5HryEpW0Ljk2K6LtHN50oOSXsuDvAVSYzGAVU94cTvCyC+kfl
efz5nUjuwefw0gOizNbbvSOUzCY6Sl9mDuckUC6KhNheAClFCiyyk7/Q9jkvE1Fo
K6GVfF8n+5WqdlxsN6JcUkAun4TMYDp0FTFXC8I3oIXqsqW/ymRviZ9mic4cFp2y
1EChxTS4Q/qn1v3EpBOGT3dtpB+KlDLjN7xj/Lti9NhDqF6XGhF6kiq+VMjhIi1J
ZktnVze5cDZ0Qpb3N6FspeNRsFaCc7nRMG7qh54Zfr9GXTB/KKYesvr0pz4xWvmd
NLzSXUOto+AnsWK3hOOw7Kny6CkdajE1pySZWaZgfKHdH9hB2BiqG1DlYDL06Bb6
YXaYTulL7wDgFbYGuUoBbZ3fT1KXn85cf7XoQK5tGKxFxMGK3DUhzLCki3YRifbw
fNlrStdwJB17SuuwJk70mYwG0mpnbAdDjnjZZnMApusddBiGgh+lR5hwb/16nFkX
squWT6ANp5F1fQUDho32GyWspWMicu9AAsLg33I4L++oqJS7gf/rZtGIxjCk7EFf
qMTSfQC8vALGeb7iTgtTrnWnfGDW8n3jK+7uQdBl3LyWxM4pG8AIWL/52HlFKDVV
9Dmi/XxTPPYsIPrrwHIVM7PdIVUXNaMrp/mz9QYyuhOaJDnEm4h6VVi2okXrH8hk
agCstJR5+yJK4gwbfUyvUc+IBbRSBAmKu9U/ZZmJWqPugpbpJwLCTeWgmors/lCT
hK78QG5JJdJsDF+ebaMUAwOqGbf+hMNO6gmRFhVZ/4HPZhfaFENwyynL5b4Fp/z0
d1FERbPumh4RKyE9mspiljlqCCsif6XhUlai9PT3xGXgGt0K6bcPGQdc/Omao0sY
AIShL1WgmaPYDoqjJMYLoU0+o4VEjwIMM9YxfwslJvXHFh/L+Bn24Sc7vvv7EKDS
4OQYFu9FWSMOILW2RZYgnUZ/5nM/MP/lg1iEgxyapNPbFbaRLQ8Hp0fbAemwt/VO
9TxpWbJg8bNhwz+i1OEnmfq1TKmM/CzD9RzflD8/KQOTdVW/bnq6pqgEWuiylEhC
EQyP7fgcfbTm8Q2I7vIPb4OuDBZtInIQ5glvXnGcOIVjTOqu026R0vROuk4J1cRd
m23Uty3v1MsvOi2vLIfOy4FK1oVVRwRcdx6ARY/IXuOBumlve03tytTx4oPm42mL
UFy97ETdWo23JHbf/GeIaTz0xdbmfx2Aj1wqdNFNexMn22xolEUX5ENa1GwxnhOU
UCjJEhNuBhmwetZsnurrf1RxdVTuh+mgsMYydVKLkBWqW6hLg1u7QixH+xJmf3A8
Ev5b8UL3laGXxY54gqJDJo6knFrKbSLtpBFNfgTYv6zu1Lem26aoYEdXW9y2Exqt
0sLqhX7RuHBZxJnHCDlu6mv+s16Cd7s/WAPaSfuOUDifMPJdf2KO7ytsSxOVp7Fv
RG2dFFmcSOIbFXein5Epd9LVEjFVWT6NgRvhyqEZg1QpYArpCXs3DrvDaygRIfm8
ijxVGfkSW0Kpv7WUll5taU9vIIeb96auDmYVwl6nTg99D/wKKeTwZvCJkKDvxyBQ
a2zc0XScYILrAhrA4WoQPbXs4vJl+Ok+nd7xV0t8etNpt3cuntDcYxuCnyZyOnwF
ju0Pyl0x8EqQ/K+pMThXoo3Dj0IhZqgLmG0pzXLrVFm4kQ82yApyhtXBcVKATbbu
4oPL2Q1AX8+d8tzVwiayty/3KjnXRAenhYSLbRbJNZi/yfxe/uSrHP4DsxEQ3uq3
YX7j4IwsPcqJYOJztS3IWWsyAig21D/tw3FVIhnyintjRljzd6Ee3ZF7SNMPZ802
84mK6yP6sWBarpYbYggF1I2xr60NMPcNZ3LBp+SiVDL215LSLYtxAnvWOFU3mhgX
CqBTjSvfmyxTAbbdD/Ir66WUT8cm5cl4r29SLsSowUIfZXvoy3V+1I2w0JVcVfvx
qMH5rt8z7plRIKFOvZNe099xUlKhQxc5JbwhunN+w7oc1MVgm3xXhh6UNE+f+3GG
7YU5bVNQQjKl+pghPFWzrCSRtRo9q7+g60adP9lh0emdNhDEK8LJ9cBLr6BBMn0L
79xs5mYsb0xBtU82zAzVnrAUaXtzlesvrVKV6gAoZUnUkJreXOp8k2l/dzSMJXPp
vwypaH2tdqmHB+ZMIag0VaRUTB9PPGOwCc6+hy/CocBXvcfgiE8VjzDX10mgExhz
XAuKt5xBPcqFBWMyoc97ZK8pID9uhZhve+jGSqi5IiDZeGwuou0ia7mvz+FQqOcH
TGJ/+047JzZ4FU6AnpuLeRVok/W4MvjVdE/3cM1bRoAPqHq3hwXPBXZhU3k3mAmX
oPDmcUy/6I2cWsXQ5ZlXTGG6MfGQllLJO8/l4LkNAvsLUgkrqsqAud9U8F5PyDaV
2eN9dHVypb2UB8O/VleQDjZzIWGs6qIPudspo6rVe/U6uA21buKDjMGHkTXonHWd
EBVNcg3G2/hvnxO+0JFi2uOZOuFIzG1KtWOFCkdVMZMFmXXzH8f6X8CmAXVbs0kK
9qWwo2pMQn+Fh8TOKzgAseU0Zp5f7XlBYOy1MCdq3oc590Ge1cjeCBQRYvvTg8Rb
PF9nEjxnEqA8E1KVdy90k4Aen7S4Pm79h+TXJf8z5TPi/9vByvaRhw89gaFLDRqk
tjkqIGoARPBYYrcvbYRvDgLCYpLMnsg2c+O1CuOGM3atmLvpurXGQ/fMC2r1OTOj
8d4ixepqSwAAbBIzmy2BBJHLe9HtO+0L0U3yHZBNII6lTeIOLVgwb20ZuThKl1D+
qQwPWod+hqNvUqc/3eWWyqmKadLUHyGyczY8G/2yI2TassOob0LqsyEf5kvFkf5w
uTOT0GhqqX12cBIPdezF63bhRELcyPJ6c/w4AGOtl43es9VG9q2l5eRHS+jTEU8x
6RPhT/LAFnwYAPJ3g81Bc4k3eiZ3c7tQ8ZNNz7r4YWldsnA8GhZ3QiAkPZ3mzBPJ
9YdOYm/kmuG0IKT2DDUYgV6FBESsUB1CCMAsdVHm6f8/AFFORXfDb7wE0ijVV53o
JvWm5mWL1VJ6Rvs5vU4//v0K1TpYDwEyfMg7KJX7tT1L/w3FG097v1R9lnsOv70V
C+nVtdIusVLLlqFBTQDiEUlyJlqHrgo/Jmi1jhx/AVemVDQ3pC6SUyA+Mb14+6eB
rjTcCqqi14vCXimq5B8LUK5L/Y0npnD2VYvanj+ww1unYeB4IyAzSj+jcRb9yE5u
jJ4tOFhJRqILdEMJl2ID9V+uvLJ3E/5r/plPBrgc4MvVRrHZzV25ingzpVMWSsqx
w8aYyIUumoHSGsqdtCGzVUQHDVRRzV13pBHorBX50qCbL3w0vufwRuSivQrf0vJi
qECtF4uwIxF/8j6ayaKVU2vrO8KWazY1UY7/E7vmvMselDAwzLyEyTMyHayLCIxX
HW/17MhQ5LG9ucGrbDuH4zXeZyrK2ZBJXwE9o2Yy411lU6srZ0rrar9wtZn0HzGe
BZ06dKyob022wD1f/Hniyh4O/BjX1kKm1ZMwyQmF/UL3X17u4YwuTAgOZRky7wYM
HYfVToFx8vz8EGfUpzMzCqVvCH0kX6NKh3antzt4y/HIF9VYQZNRPauhiFb4WtsK
LEeANMF4j+iyCl8+yniQym41ogUOEs/wlnHpvjFmnHgmCVYoXxqO3CZYPGJFOXRi
hz2bTpj/G24inTXAG04/DP1HV+EECZUvm9jRfR5gq3CKWQoq3YIz6l+VhNyzChcN
5/m930Ufy4O68Q8J5cvLSZY+lUDbMqgFaernl8pbPgxsY/Wc5G6gkPD9QWL7fqK/
NN2RZs8ALOG+S42V8ifGTDn2Yqc6y+wzloZ68CPg5/lxd+QCKuN61pLAmQoDe4P2
ICgJ/CLN3FCVK1QFMXfBcEGnDy55Hq7bLlbJyvjV+xR+dtLTZBbXwJJ/X8OCP4cr
zVP+tIu8CKw1EZxlQ0iYHBM/H+QTPNyHKHjjU33XAfJOd45DTjEhwHwpQgTwkeAu
SLH18Zpmyu+fIfYGvHpivRbLsBzqOw3lb8SEVzz9iO92OhCGlV8tLPokLZSozRGF
bHxtGsIpc9e5I6PUfuBJ6wyZj5WuDN9gsitlBF3IjdFacqaIClZr8f+oCOrdOrs3
gnwJpUhuVwSU1b9sS1u1NzHNaP4yyc3uWyZyFOMnCtXDJiUZDWB+9oJWhuVs6YDi
qjd2B2T7GDWTT8RYPIxHcIlBtxPPqsNmF1c3DDP58bSFAjj8aRVNLAVwTxnkxZJB
QPrXh1w7Yeei3uu+FQgEAol94y4lTPPmFIMW4L1Kdx0KNltDAYlvvHg6mOnPW0w6
ngjD53djJukDibuRVWUfBBV2pb+XAIuwBVWx5vI5fYcPaTTf1Fjc65hhf3DYB1h8
1TiZrTUuANwZcBL47d1KV731zh4vphZalQSHWYk2XZhZOSlLqVHRJbSYhxAutJBS
jgay9PuiHGsdAjy6afy9Vv9yPbF827F9HidApc22T9zdTTArel9Xxhabl+bUo2/a
IKRcGU2P/W9Zp2UmlnXsFDF6aeglM95rUtV3Mi+8oA0ScrTMHDi8MsXCFaE5Ud7Q
l8GfwPr/VZQnb0D3YaIff4VIRsSPyR8vRizgsMeeT8Km7zc2znjp5XnmOOmqDWIA
cV01taVi2tFlkAoKquO51VMlPmdlfAE8xifvNhjd8Cv7cj/wDiQzCnn4jLJApEaG
jfKKeDCPDshmEfotKzEOTjek+vTsPSC1yvyhYbSwpoWd0AFyn/RGkZ7GFqeQ2Frz
Eyiw3WGKbiZO9nLKE+0/1ZzoeLkGzsjUO6vtRSnaMNeMRvc59g07RKqh0tNPDjHi
hpTtUA9NpVWKm5BnxwCabFTD/lYNhXSrEMZ0E0lJDlV//W7Azoa4ZSwuRGUva18O
b2ASU+IHorufQr9AGc73BJKMtAZ1/O31a95Yy/XpgXpFqgn4O8Omvc+0ly2JRmp/
97+Akb7BeZ6vmotJc4k4Ybffq6AJbUlqtEYPeOP4/f17wo5wFVl3ZbHkYzAQj5Qk
LVtoGdpMgecqcTJW9cJVIWO1SFLsPTT2/E5TohlWTfWNgDLim2Iw+9QXahnRvdsa
V3bZmK6GG3n1XKZpD2c+m370TvPunkYNreg+LAs83wCYMeQ9qe2xkgkW4G2tejqn
RYpyTj4qRoI320SKPgFzg+Ab9ZSTKmtcEiAO5WKtrRc8OQcYG9wylV8f7c0qfXwG
xmO+65olHV7EkDTGZOTHze97fNGhOn+N3NHdFhswxUcF/rzj9EyXCLn2nWRu4/X0
0FHlaDzPQM2BtEtWeEV9g2vCapZ83LKdZd/miu5nz+1tlQ2D9sZrQF+/tOk1pEgg
Cs/D+ADDBxk9YDO+2bSmaBqUkY6SPi4g+OESg4161TMqgGPhNrWvVblcWiCh5WpH
Eh51y+n01vNFPghCcJR9WK6wfQHnWCX+f04yHVL4WNHfIEV7M62KJThUaKo7lFEr
mOOgI2DMHf8qZle1uaAeJAavzsq57GGJ+a71R9bppPagiU8qd9bPAniq3GOHrhzy
GB2weqLSmGNYnbiLySF5RNuxvmso7dYid7z3aE/V+Yk9xQSq/sJn0wdSTzKN61A8
PeShWycqFbxxNjhb7yAmrF2Z/1m1P3Tm5ZdmQIpPeQNk3oTGf4+pUxCgHT1ry9JU
hE2jpuqdZSHqstQgcmJKwcvg65480a/mnLglb/2w0NpjPMXgpEtHd2D0PD1Bua3t
4qPomXSjIv0HE6zvlbybnG8ZTQ/zLAJLSX77QMo/10z1ah2jL0qi1hN17XfUs/qX
oLhMIN4q7GZVrViaQ7Rs3ZNN3WK2XX3bmw3W/mPRWE93Nj+oLZhsjON55vAT9MEk
t9n0ERwLotF4SLu/yu71LAFttloDo84+vGfHvdaec3UTv52Y6PD+tazyV+tpQoRt
r0pVDY/JwLat/30JbXJwKuYRZVvf804Mjpo3VVgOgGJjjG/GLiIh7/29xPCD8XQs
e5OS2zcdbyt3fe1D7cq6rFnSZjjgON6pwtkhC0qjZbzR5Zbkqf7N38m/rhscmTte
ENXeIjJ+DQ1irr+aCzFu92ZZGQaRY0zdthmynwk5gvd6pQTwM9QEXFlhNRkdHoQZ
Tl/IZoQxYSimgR1fq9MyyJOaj55jUYDPzt0pyN4XR134t4ZJediopjiG+l00hvDM
0UbOuwyej9QAnG9CBIzCSQw3yD36BtsE+se4T+bveHo0A0MUlKDkwX5XHFYsSf5c
OmuyFPyV/Zd1Kguh9PaIWD2bUXd8neNrvHxkfA201qQ4Gc2KdkwcKIA5gj8hxHQU
8U3AcCimku12Aovon9lvwVSRuAYpiqNKih9we7LvjFJ2PR2DB+8k8zGaG5+EQYt5
9nN3audSf4il2cWjEGzW4KZ2MNCf5lpWgWsp4cMhzFxOEdCFlPe2vJdguXxtAd1j
R3hWbI7DRVsZG6JUCDjRMKbT9CPS811+5b4Zb8T2MRIj06lGnsv7tQ4ljrGLIfWO
lmzmtuTN80p4KI6T09q1ZQgvH1GFpdKTKez1QLljfcNaw5Ao/KvbNVrPApe69ah8
V64FKYzQudLxy8otxWhJuXOQnff6SPLJkqELpI++7qDpNLeI+H/82MVvzriYhSxb
USNq484PARY9iAoSEMa+pxfpCyliBLGZifrxNdDW+agZ4BJAvZcB84vqymtP/jyq
F86QwL/HqLksEKggHV+HxXPVl76dM8aQ30TO8NtqSm2hM8iOzpH5Kx4MExFXFcht
qOb6WsEmpO+qg8zXcn1+ENls/oOG5qwVLvYudRESHGffEUSdKFieFIjbvZZo4y07
/aAoAU9LCkogcyY9vZb6WuRDrthT7OcEsuU3a7MPNyfSgQOeAbq1lCUyWc1UgmFd
+HhQeWEH9UzQCJf3d3wpq5otduF/ZRNFAB/2P04GT1tGaHyoj/UA1azHA6mG6uPL
9Zv6dhq/QNwwdmCW9i2/Px2tFpCohcQ9SenTBMOmPGQPh8AnbIzO+e60wRxC6gwb
yil3k+kd/1JgsTJryLK1H3amwznlrHT93mfKesjcObDxRZBy3MhZEZW6LUI+GuM3
0XGDrgZJhMcZtORNh/2RjuFtob6lmRafGnFu40LiGe5chJ6mAYW4ODTL57wlzqmH
DQEc6oPVYkokJSl0et/2J+q/keKpODfmGcfPhaPdcDaIscHMFUgkYwVrcTCO9vK0
vgdGvVoKLGGL6IOHcrdAca8tdvOHBYpXxHjxFcBEaeDfONvOXiVl+fE8UWmJIVsB
7qh1C5eqND8MYSHeZfu4CTa5WxdTpfndyoFsZ/FM2PGg/UaK09+U5AiSLlH7FTa3
tKq51f1NW3ydL1I9wNa4hrgrYrZ0Rcqe83BPpdgWRXdh+gvR5sTqQeoJZ0NyjVUJ
6yGY3W/hEPPM6BavBc1Flw1Xtnwntxds2IgeCWYLpdYsrK5o+KoBkHcbcEA+QGsz
nToUB1zjSEJbd41czlZ6LOmxZlKTFXS5xJ+Fu4beu/ax0FGC+55r4xRbZBoI3jJ+
vZYM7Z2czPFeSUhxf0A4o4hYrluuG6GXfq2cJ9qBuMvLeFS+wubekWNuA9oTTPjv
dK89TCA6iJpkkLs47Yk9VJVwqM0ogo8752dYvpAB5jLRE/v4I3emrAbTse/Nx+CS
NJGNNvZmsSGh0DCK8R/BlLEdLw33GT2zmY+echeSmDqL3a3MXk4cXYGh9orXY8F4
e8N1rQ6/XdAS54VbE9pu17VB097TKYMJdPchufWEtqwka2jIkBbcwcRDEDZcFPlX
tpMwm0ewjdo0s/q3r5Hn4BMpZL8mjmM+ACBlThfGKtZpJl5xJs1eUswzuEffJaJK
Li/40pLE0rEQr6ODBT/TXpAUFu26WU4CQo8y+rkYNaISM56jEuZcFG1Iud6LxTnA
NAIH6ownXAWf9p2P27IiVUfKBmNT6BU+InfxLY4aaYBIB2L5L5v3knHUXgprqLDc
N7lUR4RGRmewPC04GPZKGfr587TIS1PLq8mKuYkYHc3PWKfLixmIEnw9R0+Ge1XQ
tXCnmRzpsKL8JOtW0Q2ebMj4vJUSeQf0xMk+Q1EI945skSeWyJjifUoIchJesN9H
KP5lMgzcnleL+j3Uuq3SckB+CC+dk+kRmlg7EGJswJK7ZlKRrVSODRcJvYuecNwM
VCUgftLVr9B6A7qY3kVSLJeecRELYFGH2n5oC1VORTWJz7CWKQqnrL0WSAhtwMqu
f72ZbPpwhBfPpjY95rKn1RI5ojO/dvd4B928/RfrkN30rw3Esp0ZT9ZhY2PY86BS
hnBi2osR0HTfY6jgtAxwGy2gFMWSTGIZs1Lv1dIQaxs1QRrAFAfOO3FeF+vS0Ath
CugWmdka9padUoJ14xahEAQHdT78xEDpqPaQsoeyY4h+sWW3NIuVwntI0GOxXvyT
cEDqu2q3FCnv5pADUjfTk4OTaZWVhDmX35e3//oSv2/wNSoTt+ai75J1iFbKvqUP
2bDOWKGz3+7d/yDN8z/UmEDBshBAtssFog/ABthCZWfiR8CKKO9B0H7bag1xMaSX
Za7DGba5SHX2cuH7eP8H2zXPr3aJDYdb35g/KpxXyacZLimISDUtqtZEKkQ4Hw7C
oRJuyS2ZmYuwScJjM27kwUcvQtPr8mXeYurBWHZYL9hwZoXMTfjN+VcosgsRKfFj
IvoCGuMlAgJbiLPiHDn9rZkiU4k5vo1635ElAHR5tluE/pOm6YX4/YGt/77V71l8
FvCvTP2fHb+wFdgoiwOWnOR0rLirh23EM8vFZVNISAt3jx6WbuYiGDcgqYOSz/xy
/OlUJQYzCZpmd7seOpDdCvbD/d54VuVkXdj0hSDtD21t8Ct50U1FPP+xOdDziiAi
kcQyc8pL4O1MfcpatFgicr8x8wD2SpLNj2vzNXMyi2/Qz2yxZENTHTMhGTLAD5sL
b16FHOpzDZ7G5/MEmC+CxqeMMkV7cphwb34tmXWS61yEGz/pvqzjz++gvq4yxekc
3E01V1VuPcgmHGmJypIIgykZT20WCzxrds0F687gwuYXsj+Nb6/6/4RHPwMeVkyR
hpZp6IfrUSrs3/ycgBoUa36XHrzLCDk5TOp3wdroaDFa3tK6efNZI8v9GxEbCNFl
p7Zh3Jqik55qI/Qbhd4ANLS7lyeK5vC0xt1+TjAPogUMj0vWV+QGjnIHNwSZ9f4K
UgG5n5+wYv4HP/JkPKnDlSwzD9M0aDW0rhYIWoJfL2R9RXI80+6fWz9RA+vr8pUw
4W9G1oib1YqY/Ps1CR16istcmX2r67bPeGV6T5NBLKbXGW0D7xApCamy56hykvQ8
NeFSlserAA+X9HV1a51V4V3feV/btma0quMHA+HWdo6OQakbeA4RRzdOOiIIpjoK
BjM5V4LwEEkzj8YrUvXNxM7pg1FD0ITP8TSADoua5wl2FmovNwPb0a3bKP1jNEUX
afig+ZIYzTkMF2G6rJInoF5OBgecyyxcqqrI8VU3kJt0HxJdzYKlUODNuwPYlyMC
XoKsbHqH3upaIKpfEh3NVwdDivy2Inap7INrEmLOEIELajJCktnLETR1+pvOInH9
vT4EtlZV+b57V+cKvwkbmuHoHPxfeby8kIAQakNHktm7RFHOYClSajbRWzrtSGcQ
3mwm2bLyXYs3KS66FXebc0Sm8FMwH9Qsvu7FdBiujAuX+Jjf2pdpLw0HDEXPAOER
Q2rjI5pVJ5NTfT5hcECwOHqpzDxc6pq8eeMkJ61L0qv/ivB91JqNTSCX0ABr6oHo
EHijpbek5LKa63SaWqt1p1SSXOYA38/EhyY6QAgXTZj8NLf1XxWLgTCpCD54Qkkg
bJ02mS/Hevq+6saiVnb5Yfjpoqs8mlSSpGVYA7W32wElQ5vB4OL9wV7N2twHx1Dg
L0X4R91vQ8JP2841+6kgm01YzXqoDMVPdiOovdXm9QGQ9hNWxjxbqztXa6nN1/6q
ErasqMWujHGUfL3DybZr6abG3TftBTy60b8K/12PQMOtkkfk+ZxR3DEKrFw21CZw
HYX1W0Utnxlm4m5DdDO40ikCzeU9WyMx3K7pxK93Rwsq/KGSQT02lT0IbQvfs5pE
wq2tlWTEViNzujDHG6KbUk5la0otxx+FcDKhaSzfk47CpSOoyjl9g062DBZguvGu
1BrMnxgrSvTI1Zy+u+uEL9vpDzmNq57Ac+e4KOJ+AC7yKElXFGqMHdpWxvxMWZMj
rVOsWWkzGD1HtbvgnwKOyLL9VAWrayAERfkuC3lUCSb859d7Woh+fZ6lwap9jSuh
axcyv0+9ky0g2/qJWVwjoIAyKdwer+OQHdKyLzkhcyw5DoB17sHxATj1+6H7twNP
zVTnG5u5MQZzQqbNz5kfAK6t5apaeWBVOxnPoGiJG9StvyJZy5UPAobDNwAVmkFg
I9elVRjbOClngRcyaqd0Tx3mEuLm7nRpKcNHS5sZECBK3wXjCh+cAYhodWL6oPik
EgcczTXelXOsKe9EpaBTxD0tmNYtGFZQ1CNR0P7ZHIrFfI00HGnvegL9YcDnbt53
eAa6Sk+ey7lDeJLYUTR3v46ZVSaugOGPRWtUFRDf5p4aJJLiS9Z66rOTeaYEUSqY
C5BvZmbrV6btON/leVIfgyl93Zic4JBBWlwlJ3eK1IIS3bum1wxWzzFVNSVF7ZGV
pW+LxKi0ldm1V7flO2RdaPB1yPA5L5VR8ibYU6ciMr9xD12aCHaYfvpAPHxjhklc
XGMxTBiKY0UVV0O8C5DycGZZwrh71KZcKocWLRmG97bHUfVqcOKUITMTCT+brBCy
RvtzqDHloZ0h9gfdH9jdQx3wz+YNw7m1mq5aAX2clhV5bm1wBia22y+LSiMnxTk9
aNetc/bFoI+v3gUgwWMezsHZEpZCjCBOWgz+jTfNyTU0m0yZqaSehPJqyC0BQ+ak
P12lTbhl7S5C+W37BsOm3EYYj6e517zXt0n6ypxBg3QZMnEibDmSnKYpK321jR5g
d0x1voR5E4bGg0Dgji/mxQq32a2TNRLGmq/JYwAYG75Fgm9bO+ktrYMzBHlc1qjE
FBPnLg87D7JVRpbj98ogLZRUAUHn1ZvRJVR8jcOs9LjR3iluhAzpnkSULuiExxtF
xvXh9A/n8l6R8mohJLD3Tw==
`protect END_PROTECTED
