`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
eCMXS/t8U+DBdS1kmeXzB7OTxn/tpuIr9oXnO7ltEcvfpbOEM2XfstzSfyq6R/kA
WUtVFek3SxBjdpn/Aev7Ue4mP+zg2wsrcZDhQKLyfm+WOpbTFLncWiMkl19CORee
97/dFAsIAnmvncvYfXYe6NhblLSMxACRl/oGJUgg4Fd7V1oSwUj7nIQafjJZn4+H
k0CPUxa6+GuXc8aBQAjb2gV9dKO6dm+4kBppK7JO7o11DuELWHxzlxg+MLRZw1EB
fOqgtKlP0mzxZinMddsZqfr1HtEVNQuNQIhqu98t72s=
`protect END_PROTECTED
