`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Clk/OkaIFJGbGcLgfTH4s1Ba2psbJqdLf1ZdqQmyivDKSeX2GLHbXE3McGNaU13q
zMMrlAkWT0TUhqWeaGjC/bxJhyGVB7XdqU85cRUU2TLYC4FM9Oi9MsXlQWATT1gb
e9bnRic60JmjARWaPdEd8npgD9IGFBlc0/prwYOywx94OfzF1PJKwdiA5hvvdCGU
jN+B2nV8bqOvvaXj/7Q671By54avfrY7ApQT4XIJ9LVr0dm80r8Ey71ZBrqNFcK6
xzm7x/j02NWx4fF4G2ulHMdcx8fhgJDykH3oQtMweaUaX2h6qRQfHHGUt+hQdq8I
T71ozdaGNfypqT2IsGyuq1+Ckm2mucYgmNNetOpO4L2UlxQpan1uP5xT2M8YGYNz
TFjzH+Ny1TqlMhaE5mYn+4IG2tWTpH++FQaB5mYS/FFwhXJKMlU+jOXzrNOlKxo3
yke6XRba9BvDD0WZVMPe/zTqBCJrH5fFQU2C5c+V35dy8mb9kZ53/Ipez0Mlrand
GyjUvNFOoVVWQX43n6LlhO9WMHbfjqNfQ4ZvxMnT82nrUXCl6AxKYdGXOio+XdP2
UDSjI5uXQwG0hkrxsZzvtg1rXBXOhS0s4oU0SQ17c1NmJDX7JX3cUwNbIORBnw2H
laqvlEwM/0rS/fe6utvifeIkUZgXXNV9YwcJTQXqMZNQZOM/X2Vm+PC2Cu+YA8Mo
evJHyKIy4SMjhPWWSMkdG3Rf50+TKF8snhLnOtkbjjJGIwr1uevZIS3+kTBOWOuw
WgGbJ/PZLjDESGNqneAjxFDiVwfjYUc5HDUiuMNOdCbmx9DCKjXjKOXn93gGeLj2
nlAQOTUDqKkZJBZKPZEQwBM2pmdcbEcD48NyhfFnKXacVnX7YXYfVvTHQ4mSsrT4
N07r3mriOv6aUUdT8sxXFY1gD1Hw2EGr9GTiX2iUbpY=
`protect END_PROTECTED
