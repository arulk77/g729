`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDskFD73g9ZoNe5gbMA7QR2x0m8kJE7yHj+khhyNZIKa
EBRByEZRDrMalSNFjj6ng05vE6fnb18bekrdtCNArgA8JpcvtGG9BzQLQer0StS6
uqMZQMyUtWoS5vy6LWVaGgKXMp7jDEdTIf+uCpGA+Jyx92N0T8DOkD3YJE5m2HMc
irH0HLk9HGnvF7V52OtNPg==
`protect END_PROTECTED
