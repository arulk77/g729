`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEg9wyS4Aem/fYgOh5M+wyp6VMeITaXyVg+FwVPdjvqY
Lb+/JuhwFRsMNv4lVg/FIQOPDaO9egrNQjlTKZV9JXa0fG8vAzsoNpfW3xhRS22e
L+9ypHEADluhsqIOejlMjh/iVZdWsXkhHZSukyzn5N8RKguTkc2P1CmuhEBkjOwA
/FIGBBkl5OP/4S6Q1SPePtlM0Bp9RgvfwZFeQoxH2KBHl5C71lAiyn3AM1BQhNTC
qwRZr6ipMcwb3MTEyj/hfDUo9Y9bclB+4V36tg6wsDMbP9My1A+npzaatv4Xtb/e
KzxavUhMQjaOMkAP2Alf4D75TE7BOwkklxVEjdIL7swC1HPUbEv8ZoUemndiGq6c
stYixmiZE8bjewlC923H+MkF17rARALqd1tOzv2t84Fa2e1wkX8f7FdUiW/Ui59z
3KIBb43paA/BtoKAonxCvlWPTJzTufxKTv5uR9nMdFHLcm6m7uoNr/tHPvs+RHZF
gDOBJkH173IckWOkf7Vzf8aoCHn+y+8e51rMUYnvy09+fhMV040XqoJPcS3PHasf
ou1WVHyqzFgU+/PSN2U3HvR1X/U2Qwk9hQ0iCGwPKQhQV7KsNjxcstCqXblmHMeg
pz8NA6qjjxpPzOlDaV5BUUfji4qQQcOjpx+yTzNlPk8hAuSPQiJhBEHm0PlVHif0
3Ze7XoN+hqhBAx6P5DiU8v9Newy+owgxQNdJ4YUYjMkM4x85PD37Kox4K+tZrG/5
ULQ6Jsgr3QJoRMdRL5dvZ6LCD1dQoFGC93d74jx2Bnu9mf7/tYtZPJKrDAfb05Cj
0QOc3OyNAfJS0Vs9SGHT+kab7GjqINZ+a9p/pEDrrugxRKpoVAVeaBQIMRy5beau
wdre30UAihd9FLXFEeN30VSQzZBQ5Buogh3q5FzbljUCKNZZTBeL2Il3JBoJuRHB
olotE6gHasMirawz8quEykB5xZOQHl3+TYt78VLH68pdnihPg7DGqnJNh9y0af4U
FsqHwNBpGTpOjigTN7RnLlOxm+YxzX07ECHdFDpHxBitbIwecO6JokTUORB+se18
Uwq6EqsH4huzQH+8qvKpawKYJv8Ir9SGWDsiyZVMR4Z1iSmSfY6GkyzrCyCL+zgE
5hzzqSKuKMfOBUuCuqDnyf/LyX2vr5kXy+oZo7mm1kUz8ny5FAzg+utiPvBYmJI7
ixidGDhx+9m2/paMz/XFJgavh78CvIGUzB0QXB5qRdl2JOwzhT9jfHuz+oHvJbfw
v4dOWOCualB3SYbGlPC+ZhqGCttZdO+VB3H8o2dYtH//UlBgwhvXJD/4FYXOlvs9
/gsVJR9tAQ425TbaU0O5Angbyy7+cZx1G4XEtMcYdpIAvJGv1h1T4zSKtiYU0nJm
g6hqyH8edlb+cjZ660lTJu2fGyveIZpwp/zXxvuJRF+It/Nk5cssaG46ZhVggb0d
eVxgjzce4Nnp2718BK0vUCMzSyANm68DuQgwxupR2Qe7sV36TXhOy88ZBDh/6bSr
xEeWpqK58scKOt7RAwLbBYdKiVSzpxn6D6kkL3lClR4VgfE2fFAKSnPW4wijXOtH
7C3TjHdMaDOtaCPjKSmop/P4wauq5WZP10vEZpH3c3g9ky6U1D8PsGwJc32h7MBA
0T7tOlzHeu3BXwl+xN/qEwjwdLl3UAVUXqmGbRluSesi0tTD+kkNg8sHP0sKK0N6
HjH5AdwfuYJLnBJN7M5e0Ftnm9gqNrBC58efjV68UopXx9sbIiYdJW73xTVNVspX
qGczPyL92CPqSjhVhmNcwL8AJh3u7fmlefyx1fVMIUlpSzysFG1Va6D2XEqEdH+3
8db+UWnkQjtqUVaY5+RKnpFLTwVhR0ANO/BNHxYHDYKAYJiPQHt73631DYqIAkE7
PhYbyy4/LzqO7iTKVDxcw+SsJdZ0YWitPZ0qTYjoCgPbwAncT8Hijl83No46VGkL
NxhFIDNozGAKxvtvz7Gp15NMPpJ2AHgr0W7/ooReuY5rAohs3UNdqLF/rz4EUYMc
Ccqi2xKwljMu3FYVZLAL7jDa+Ulj85NDEebCw9I/xCkWaCvp4w61sVYVwy497oKP
hhjFmEy5ESEjjpS0tqM1dxgTJy6C8LN4a8Mw1gmhA6RorW94d53HvCUUEIL2PSPU
4SjxcuTvgPAOsRT5N92Fp9J9yfJDGRlP8GR/l2ewGonGzP4OPmrVxGGkDPqOZWaE
7Nrn64olDjlPKwt9W8o2tLTwScMKewGR8zTjTzktI5NdcNoUydyL5NzOrn4x/2o/
WVnQFt9XmA3XiixAF1d3PaA+oX3NDVgwJgWpRfc7RKv3Nr1qqa6kihc5KRF5sP8W
gaLxwwIhz2G5DNjzS5JRFPf3TX6smk3jg16FWjlYOvb/291V4fbrGTM5sKjwE/wb
xezHVXjVwfpgixIawLzauRfj14OcISnjCY6dgdyUrXJrLrHUMU2q2mQXNngQIYv/
WVhZnAkX+Jp6wef4exOqn4XqbeimPldRXfZynOzzWfV03n0HZ75jR1bPKV8Hvsdm
kZoJRu9xXBc2xQJ3lb0ETtqcP4TEWl1Tjhk2XYwVqs8D2WiEOZ+fXvQ3VV1M18MW
0+HX1OXhYy4jsDl2FihPX6BwdCuXV2pQIPmcRQ+vG9s5eMSyVf4MN+Oy0XUeep0y
Vs8dW2vI0I/HhG0frCnMcTRf53GnNunm+Ur9ae4XJIVDp00v1xkOnSTL4VEjwHkF
AZhd87SXvwdcMxRdC3QaSDGToJlnLsRis5uLX1EavujSfRK4eC29bZNDaqKnpS4O
O8tWzdZfEoZV2P3j6+WD16xkrbD1Pu6PGQtGHsEjMON7Qnsw9s/hhihbHsTo2VZV
AtpzWPqjydGQJNrrim3OkKyfrVSKX40xiCS6LIO9rOiqKg06Ga7rplDZXzdJ78d6
nU/2jyKJVCWf1pC2WlluFlBv2YSaV8wassOE49UlgMZq9GqF1C96lIUIP19Tgg0i
zOEDfFRv++/sRAaas7CjV/Tfrg5RZwNa4Z8wRnHJBr2ZN93T2htpzBtlSURtSLw6
RvDEO+295+qmoK4FKUhcdWM0p4wS3U/+qeBtB16KkHVDpYjKgf9miywOQRBiZs1h
F/krPacaJQwB1wEaAsFp+d7eeOUFSHtByayO3/c0Z/nVm9Ps+Q+PEZ+B55nfIxQH
9b10/EQQZhVY3Qg9OcSD8FLGOOxFWRAH70nEg/6LYBvHFd7Otsr4KLSr/wNIQuMM
qmmzlbtp6o91AhmNC+7xiuPjW5SvXgi75xj4Fv5qZDz1vw8sW558UICnrDDtC/Ly
ALmiXNYroffLFxSLs5TNQ44bNMvwkLe3tIvAsUn1zn3VsXFwGmwqhuyESFg8xfiU
8mcRoxD6EBFO9juWlPiLUx1DbNwGh0OFR5oelAWOT0u+k3Eb8pyfstC0PZA81IL7
gCMAEB/8rkaFC28xHBgiw3wqYii09xMDHbpzWwu2mHG1lrZqAiSFqMrPoE3Nv4Hg
HUrW6YC9LNSpMJvQ55Jqck1Z5vNIM6vP1FSw8QoGW8QAjogVPzx6wRzEh+XsQ+aM
fJJTaELmcXpDvl4b5XHG4mpOixFiVQRQAHqZvunqRC4qJ7z7rv0QtifIM1X/YZLk
/l8+mYnm0hLCdIIY12u1S1vUkAJShlgxD0gmycwiss1/mOyKTUovPkCTZhiVf24A
`protect END_PROTECTED
