`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47eyritd3KjAXrP+5vV+PociWXdTAOQB0TyS2JXlDA+K
aIP2RCEV5slpMR0uJslZm2VE2JpjsCVIfXmwrf9eqh7unRFZrFFdYDY/hI6M1/j2
CAbq/SyA5UKm/a5Z/oVo4QGtbCPb9alnoY9wDRMMvxT04EPTjn/jbAMjK92TVFsO
zp5gqRQ+FU9BQHDLbKfClWEq2g4HV6ZxsCBaaorQ69JUkxmLy1xwe6hXQMw1SZ9o
5KEVLE9UyoTjP0ePorzFIMGPVX/Ty2b5O7Rq5XtMtwed9ZxKrrkDX3BdqaC7M4dR
QC3mQ3an7lfZGxb+FZD6EmX/eMqbrG49n9TAKji8yL5OX3GzGM4ejcRz2cG1xUKr
ynQjvSYh2rf+YGTMEkA2mBeax0MpjVgWUiclZjL86oA49c6sYQRDQrmi4J62NLHQ
RxN2YPCnqCqh/kYQaqxrwA==
`protect END_PROTECTED
