`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Isew3HUWPPQmgTmG5B4eSvoLdtFArT8Ic7BCuar0VvStDnps9eA8ekcpGRx+Ap0/
hdu9qDhKjVSNWDT6KJiVg4HEKo/bLGvRZsti5xirurM8IA2RGXo96wf8Vf1IDMTi
ZU3m5mhFJMX1SQAtBcqSXmwCrjYvKU6jl6PQ9Njho5s2vYpC2zo3hh3l2S++Bv3X
AAfGIcP/oAXu/e4+uGq13IATziu6Zm1kiJhh299HXJzX2oUcULD3cLKeXoUqu+Hy
Gkiee/Cmbltk/e0G5WcNwMOVyYGIUdeFrLlgyerF94h34f2SCXMwmgFTnOmvmj3p
EDkJwtv4m77zeF0BjpW33Z6BmdiQGFs+oASSv6AkM2Tt//IqQbQ1145sc9We9BvC
lCi5PpmbMxdE1nMXHxfVv4w2XQfi1rZznTrIii9uPkum85LTwnSALBrDSiW/DqTP
jM0U+QgDzFT+B7jlRYVWNnPo6nODeWKvB0YJQbkm1T5S9mUStVflMx1helITSHiP
mzcsirAXciYbyVy3ar4wjw==
`protect END_PROTECTED
