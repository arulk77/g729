`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLR6hbUav+hXhXEDmOdQUwgNX2UXVD2UmPR4C7Xnx+qe
sKFq4CCKY5crPYVnBuFbYLg06gT2zqlhaB9q3stq4WB8z1/+gUbtvuK3xo8H0uR/
hqUgGw38vHRpS3rqnSNSj+ZZVvUKTSwrPi7oU/Hctj0S018k06SDBFrp344Q3EMa
O772brQdWdUhu55isJnOv+rWzyRm7LxAeO6iZuZ5BSJYyvuNPd6tU5iyS/UeMm/9
jmzyf+yv95wfVzqghElmWH8VdVK4pBU1gBuqjhDSwuFOrqcRrrtg9zId/4ezxzRY
9LFs7r5gVrpK6++SpBxQmw==
`protect END_PROTECTED
