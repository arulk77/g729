`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
BiSBYb9LoOpluNW0OYi7qNoHv90Y0LkIauLeEEn3ZgYx+yEEJw5VtLWvSNvM68Ay
j1bDOL39lLWNOzFOjxvG3x0L+OhcA3RvyUNnLZW7CfW9AOlAnCgDaGaQ1D/Gcqti
yRVPmqN14Xz/9PyVX9xRyohbUa4rZDPyGmTem5czV1TrmzYaqqfyVLVorIalxJmI
hbmG8hJjwGnqzSNAQSrZ1SCHFcwClPSjU1IP7ubFWguazEbEjIs5Xh7HwDlBsEa4
qdGktPXe9/gWRgwqf1B691i7ut3IrGZZsPcIewa0D/Mt3Wzb4PbGg0SHmFkedeNS
lPDCBz+n/YTzqS0ctf/eb+1Dje2Sl9qZub/qnTaKWJG9OAjuaLd+8vAWIGPlmyBy
vIc0Z84rCJUNn5WZAsTi3oyauUlajwNeuNDu83WkTUcB91lyg9C+X00dWnVwXUH6
L3qW2STHz4mJADZq9t0YYpvz11fIA6fD8KNOCSfXMTuzIx9q72zlrpvVb75qnbsI
6foUSjs6hxp34a+VEc4SeW72FdwdHvWARHEnipVdFZkYRYGZK65cxvqy/I0D/iyj
lp3HUCHLi/+//NVccM5ePGYNocAyTlpHXSHRS7W1UQuOhq1+SInlQeg0DvIO8XmM
hOCoQSZtaD06YBhvEkhuQY5VLwaFr3J/uUWQXnzSjOjcc2kz/p09bRuNO7HIiFtU
UreYumAdO2pYMNjEt/JI5+kydqyVMBGch8sEm5EMU9P/HwnOXI+XbMRuiDFUU+dn
FzCNCkMkS2NgzHegPe0uO/Is/Wsjypn80S0mlBIIdW3h0WZ4JzAGZ37d6N1ofO/x
XbeZMXCUAFl7uz0nKcbEuyT6rkRXENIP9jjXVnGsI6yalHvjvwg1MinytyQ+EcSd
R03uF69o85KrO98rQJrYiPTPbcyFYx8bx1ahz10HsQ8=
`protect END_PROTECTED
