`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL7IlfYf11W7z8iWDIVtQPEEFXr9SXBsgOVCEVNtQ/94
OLJlHfvdFBfiAq2tYucj7rUNvNlbaJjL4BgeaX0QrWSL4vJPmH9NZ8ZLyu5b4jz6
tqRzJR0XmT1RLGztpotpeYHQv/PCVulePTchhFDv7IGz+bj6HkPEyk0Iyv/oLuhr
BSwbQI9G+e76edQjMREk4BSCHm2OxX7DpQpkB/B2GOqsx21k6/JbOBnCCNv80BdH
Np6FR4mm0IdyTRUcmmKo2QireTw/iOLTMQAhMqpjiS2ohF5aCk8jJX7MESSzm80R
jXuPOorJQKDn1Ai27fsYHLoQhhIAFLT6+nPKLMccaJUV9pFfOPZs24Jgaik/lvO/
jMLDN8Qqvl+7s1xUSs8LjraCXLYLgSitoPss2ShvxpkqgXwUxde1B98vWtHIZ/1C
hOVuaqLFLY8rC2Nu+IfD8q9EsLYD3u/H+jzOBjXG32XJT2XvprwIbVBsOD881L2f
zDCljsWYo2mD4yjP9jW2zT39B9ebWVHVsTrKmKY9QTrqDwzleJAkkf+OpFzzlL3E
sVYfNNT5Y0cL5uDa6ImaLbsXFqq5Wnwh/Q/YXU8SCzhOYFNWVRTwM3RCSvpUYlQB
lsC+pn8wN4PXGBKzS47k5vNceeR2YVK5QcJRmWGQIz2MPSWD1OjQhqKldRU206Os
blsS8ZoMagyi9QRt9KnB4OuHzJXPHMZGQ+cyNZn1g6d5C03VrPd0ULzOOXmexSGR
PQuVm9KCitKuRhKWKbvlB0CGH3JjFTtVCoueixNjhcvmHCbIpwrpQiES0fypRUTy
WCCPZZ/QMGXYwGUcOOA6aWpVWEHXiC9b4/XhKoYaZpuFlBwQTzdt94PiPyXliNMQ
iZEdxSd+OMicIrwnaJetsbPimijY0jG8SR5EAqded5M=
`protect END_PROTECTED
