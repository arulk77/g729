`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
VJs82tVWv/4iah8ebsRrxCVhgaUym8tL6uxhO/SpA4LsXo6g9pIBcLFNKdFuJkRI
ylT003wtMtfHUXiFrmmcswJCsQR2qCL/FeoIkmnZK3RJgTNH6F2EsOWbEY/zyoGv
8T1+nSu/s4zba40PMvs0jZuDV2IwClVnrv+YEiJd5ULUBdSimTbZmWP6J0KsrJ/N
eqyfuVG2LF4UYP7gOPdR+0tEzHEXHoBwXxQLE1Np5kCIPbloVK47bP4R4BgPBQY0
oDxx/U633P8Jk5poWRld9ST0CV04pXsqEIBICwY6k3gnjrRhgqDTfYRjQpJyGJ4B
de8AyIg7nSNvVr3ivIwFcUb49yH7xEDKwmN0G1ccDNo=
`protect END_PROTECTED
