`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aV9JL22lu4aiH53IWazeRUK4KU5iCy5n4gBoZMS77kKy
sX7ZR0eQqDb21u9vSIb2cVEHqieynkNJyPsWVp17jgXtm4Td8IlMefOIY6QvbYaP
d3mUov3fUp5+xgV//pv1hFzo02OA8ITCeAFcA8Rm60CnZ4Xfi31UDCFWlCr6Y6zL
n3zIBKuBbbKBERt3qS87xTXhIWtCWIk8gCl4cki0eyVbjV58P22TDPGDEzWNWfhc
5xVfw5YnKPFfpOFkD1fX3asA3K0YBtbJIjP0Ab3j2WSzo+PdfyImaNFpsCzHsann
RDyzh/iDux8WW39HyRuJq51JIILDKOFlZ4G//E3bLz9pcLFX6G8WuJmOr/o9P02P
aGoqkkVtC16lh7oIN/TvG4m2EpUx2vo4FyjVercqGGu20nLwdNojKmPZUq62EzM4
NtwOoUY3ld159+XXqrdYIKPlgtBPDKms6ToJ5AxUHrK6t4fvtgLW7zw9KPIVJ+eU
0EuGjKiKCjWNJpnZQAIZKv/E7gW8N6dS0XKvT7YSt/rIoMtjnuRzGn5QhKgDbBsL
HwXVC75LhqcERr979WG94yOKJh9JA750hSbbFltH0Oqn3/fvpeTFgiLnyPFNxN81
hSNbv5ngY2zu4ds0uYqrQOml/mIJh53pGDmeihhpNfW1JlZgyPQegLG+ckZGRZMK
jvSvqo2oP3IRIRCQzfHBLlo8LpgyNT2XrgvW1x2NOnYt/TMFMmm92CsjsIEPerlA
Af6naQ3EY/ldC0jM+/11dJ/dEM9iU4nlLLekdlHh30nZnqKlD2J++wOfCOzK/LCX
ov1mWdYyWNjZBDO9pbr4RYB6RFdoAujU9E8YMjk8SjFlsJPtA7hGH9cYEUyvTRQX
qicStSrSHj7JkRhNyWD7csom0soZ5LY6hc7WAouwtgv0zAy5UWz6IIvJqZobUKbz
eEsZfVQL+mMlTPRm7G11G/WEqSCEsfbosMF4AVkQKuLckx+X3TIF7sAx/L6D2gUv
UYw3xLLH+orXER+LJd5cRT/sGYBQp6+Mf/9aM7AEQdU3x6y0EEuf9XhTVuk/oBn7
1mRD9p4CY8tWdt7KqqrIKLywOVkxnYYusNIabCCiTRYixxYrLfWcmfHUbQd+e5Bb
8yyZFanR870bkBVsMXzpw6SnPDeZf8OTTZF7LIZwnPbkL35VapS+SBm6ErN9yv5V
fQhcD0IbfIgdAPaJtbjgOvqZ26nqUDWgi1lNTYkL0JRca6LHVnQ6QBvhms1NQfAW
qQOosqlXvTSF2b2ClPSGgitT6vKzEHsEdt4c8c/yWXfRASYjtuJVQAK3+6sDtsLG
Me3caARxfyY2EhNdoxqCUGAdCr/2iIlkoKOUvZesmf3sM/rmww/QDeaxkWFmExCr
kFqhygCYqB6e5sVp4TIDepb1mVp3RB8bmxKrsQHbda5eXY6kEcJ8R/av6KLdnW/a
VAi8XrRvfEGinBMjtcCekPiMdbQV+DU4c8LuZP9g1GE61kBhewKf8LnhVV+hKp4M
39TcBwLB/THll2ONH/PLQ5uinI3I6ueBb2vwTsS2Kdmj48sxPrSHPLS/XqTJ/vng
t6lilrdpeg/CbcG9SAManOJ7s09KHYHDPEYdDqG8LgDzF2WxLaWULXtYFbtcn/qp
xaZZ1MpPuvJdN+f1YbzLt+/uLN2vLlG71mkDCBis8hTHDtjhQ1XKFBjP9w4B8PIe
IpfKb9Jvj2ymAD+jJ/pahkCk/l/RAm7rEh2Q6AV0Up4cTjPg+fCfjAQNIhxnDrVJ
03m87hUO8Zcg4VTIFGnuwGJodTSgzyVNy4h1P+QQaLRissCXyBG8Dh3cCqSphdgw
L3DrcnosVvgUf2OKOJ4wiV9OVPklbKkWKwGLTAGc21aHbjkSRVIM6be5VQ1X3+Sh
qVqm0QQw1cT7f474DLHd+9MhuPcvBXmd3gwUAFiEyLIPb2B7dG/VXG0E1aN+cnmJ
`protect END_PROTECTED
