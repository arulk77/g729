`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
F6nZN+Cw1gskhc7FmPL8eQgb6ZTkUu509HZFqImM92bVyqmkjICojPzKo53H3nUE
THu6uYUBinwXQhEOLJxXMg/u5x7mP6MYLcvnS1DLj/Lt5LknGHRAqP81Y0Tx9DcH
BJtJ3ls9VlB8tvZC1Qfqb+Cp88alxaWau5tNTkVbEX2pBD+ZSNo8+VUtcPnSDbVi
yHkUsNn8kvkQSESIo/w1ARt5VMQwGhWzD0gd97mxomw9ou7nCfqyXECMJgbvgJSq
HxoAPLLhV7tXuOv2QjsoGob/DEXUlyj5y7KmWFkHQArMA0F6rAeRgqRuiDjoJUg3
tyZ0Hy+YV1uw/c16RZ3BYicv15+Y19WWA7Y00Dlo6myvNPDMEi2Zok2bKttdWkzB
VpxWE2f2L67Nb9+hsy8i2LZIIzZjePcdlBg7Cx0Dk98=
`protect END_PROTECTED
