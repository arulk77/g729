`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu459MJI1qCgSGT8MwFT6F8Bapl2vkFbF7JLv4hOmsKmeQ
UpxemKR/K2kuYE0fO8aXed+hdmh1RU7m4ainW6nIw2wBODYR6/cHqZrWMaYlJREt
B9K3GWsQCWonoDhbN8XnQuCg5EyJ/xrep4/5ye9AlGiG5zRxYDu2tqjGWt9tHdcf
umMU4ZP+b6Z8F0F4sDFBIgfOzL1o4TNFlf1pGRq3dWQ=
`protect END_PROTECTED
