`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAQGHnUg7w21WpW4WFr5jKZaO0QwqozLz/SurstmrQNKh
DmNTZOCrGAdX77yweVHaH8MTJ0wMDlhRrqoCAOmAmaBEnSdElWsHsemYU+4/fRKv
rJIwBIv33XEC8ZC2pcrPK1SJqAxzS+zMT67PUkJlJGLj2BUAsi9NOmJYWAixng/i
eptyq4R38JInFuScMynhzpOKSvebhKqLM/z3/hdhbEz9atWi+oMZ0QMS4dTiTkDO
+/4ZNmT+VFqxckHVeHaTgsECEsbXvtHjqq4LQwxIzhrom/sb5/gzsth0NDMgz7WW
vYEQjBPTiV9QQ3yX0weivg6680w0xWVlv59MWpXxqz8Bir9GM+Z1XAeLt9gwWijc
rgk89uJVlDin5qBJtcu0X//F7Q0kTCvMCg9sXtKd/NldGM2HiQ5Bn/2Bz+olftC1
dD75ZGEu5Hqmy05/X6RSmr06R1nzxC00+NsXND/K0HJP8K9MJWb2NEcV+ltvXrZm
nvbtd4XV5TaEZXUPylWQvt9KsIsA+UzY5NL2hnKSPtW2rW7Gx1lbmQLojoOMD18o
ya8IzqqfnGoOuY3leRaRrXrArv+JenbFhXCXustVYkFqwkaq113yYZSg661R/4ps
+Indan+cyzAyKxS1Yg6Ia5gVSWIWkn1h6DbWY1W8dU9eKeWbHMQh3tAsOQPd8fqi
Aa2zZ6otLNlJ3ZQYOGXM7PVLLkOn4xhNBwQNaQ++ao5qIGtqTW0fvOvOSGApaFKp
Ey/3cRhectgr28RDZe29teHEUukNbtHvvilDj90nLzJtvWxXEwAZ4IstPNamzKSw
PhwDO2r0qCIerkNT2lyUjJeLEoD7+Sraph+ThuxsZeXR4gNfbvucskqPImzj5IVy
eVg1RsrJSk4TZNk8RAWqBFN7s3fhIJSO++PZAciAJHt7G1s1EZ9OIYkuaDeV3Bbo
2XtIaJn/xo17i/27MLLDfh/nvM5iZjhiFfdexH0lt23cbaS8vniTt2CTkV931QFl
eJukxJ9D+3mYYKDFOW80OlhIMrez3cRJDsrbEHY2atSWppgDNKskc3mSA4WtGFHb
O491EOXu7ekklE6TPspGr/p8UNW2vaM9k2G6LQls5QeEtob3w1kJ/AQGOJmpzYPu
Ne7fUeXrd0caZxnQZsWxW6jLmA49COocpUrteO3OjbDm+03i13GW0vbpaLmaUG16
MvX8fEXYfUlNIs8W6Q749HHp8Sp4RPZkvCTzWPQ5oeIysJaHWDHmYzMJAmH5nc0c
EI64eZiz11VjJsR0R+XvTHDRvkEdQXivSGF9IraEtaLjtLoJHFNabItqKLF7jqG/
V/2VQzKNqsjCAyh2VxZqgoqIHV0febWj07rFNzFQ+cnnbsxWameEx8SlBzJSpOtf
kxablpWK3Jlh5HIwlxQjGghDSL40TqENGmetAS6LGG0dw3x2NNx0lBuI/KQk/t4V
VkwedIDXGuF4w0HOJBIZwuMG6aqt22H0f2UmhvrmTxLPyLuozNeBZdxSf9F7OeDc
lIDj/5PIqFY7xmgZ5im728KlgR65IvxPlgcn2IzGeNou7MxVz87AVovRYVaUJJd6
kgTWqb2RbhIXp/aVKBcuSlSeE0m0zHNtkNpuyjJCj/RMp9ojGW7NjTOPbELI01Yf
IlCamGyLnDrCDuELeBS28ue46nVw0InSpwqnINTLHam/5f06lt9s+AZgvyoJ2oY/
tX3hwX/GpsHKLuhYFr/X7pfiXXqvmIaSetxag1345rAKdUC6Si1BJSRyMM5B/YJb
oF1Bc7XwvSPIZ0OyceDZ+7RIIljbL/OdQAN58kDI+n8hWhEhLzHjVxcQsDK4ObKp
d96B0/GJNbHUM07GX9dsze0ESzPhY0px44ZjbmiJopDqsEgbYyIgEzIJ0/7VsSl1
+ft0QbN7BRf0ddj+vg3QGNU10+fhJ+IqI1rGu659usSGhSqAkra+jf1MdjyIJLgB
boUO0ddv2uw+yd4j59DS/zsJBec2iBgLpibxtIs5fnf41hO6NMg/S7o6gB3AH2c8
8SH3Km1cYmv5vFtNR18gAAzTUzUZzaQ+emI7/PYrQmXNC2j6EXDbYljwfenoBWvx
MX0Ka9cH+2cWHDqeLwhZbv5agpRstO7uxjRlM/YUlMWfAwpZHezZUIH2gn6PXaPi
C6U1CqYGPXTSvCx7uF4OEnV6WfF0K2V2nEX/YMBBTTGiRx7JQQuuyIaL90/Ommcy
57kd29yz/EDFARWgBQIwfS31h/ueaMT32RTT0pyWjGO0pKRZhk/8W1SKhb3YUmpR
1DGdw6iQbf3W33myLF67XenIUOpH7JRL7iQ8kEp/gqksgIQVcWxmRjCMAkh23BGs
W05qKtlcg/n6l2gioKIoCz72flHtnQlMoskAIcZ8dPa05wGcuIj+aFkpKA52cSg1
7P1UklmRKYffNi2TYCtIXVHNPNW+Q2LaMtNnH2yb+5Fqb7YA6T0KgUGPpyDTjAVR
VPF2RobXXO5sAllDz4bJdI36XH82BZ8HeD1jNloriptWQG4NwdqTW4g5BO3RSEb5
VJPZEuK6q11FEc652fulxYbHsV/Yb+bvxxoC//gKMVNzPDHpKqh/iyRE+5DrlZCK
Ac4cG65ehS/+PVmrLuIdOMYNjDR8gV9nNrivlpmm9x2yxjx9DMWxYtenjWWGbGIK
lTKloygb0E5lkgKyf8g/kaxH4Ok0bqmMUCvXaJTmoijmsgdec9qbChMR4Ct8OeuR
PkoE+5KeLgiI7cOGUEb73dI2Q67KB7bzFJ8eTqO2y8t7KCVKO+AfzcwmJKxy1ROC
Mse3jQWVOL6OWYdJiODRKIhUMsrXRhuK+Wi9M0D+iIQA6yGipWrhtEuT0XeVlMiF
RAol+PkSm8lGgg1+5uFlhdm3dflS8/SfqYsHOIOl+UWu8Z7DTUMHzvgidNVfBgaD
gcOLKPhcQn/o3o2zsAEVmSRjymytdoc1eQWWO9st2tkTsNuu2Z1PE+emsRqSYPs+
vxu17TwdUlvrIyXm6Jg1pC0FZpDVB1i/bJNbJbENWQTg1Fcm78F5Q3Ud0QkfvOWq
ZLgAX5sy0Z26wCREuBJax0gawcAU/9KQ2L7D4svckhMMqdYRnkxn1Mdy4zhQZhaQ
jelozalfdVSWV8DV6eguynEvZ3uXPWghtbIoyBCrEZJ0j9u4EFkoJdZc+0D7g9wo
Rm1TyCiyz/Y/2jaRGVUOZTEOpxlmdC3qJCAaKmeuQa2wzz9oeVlx8IFbYoijOFXK
0aQr/WK4FXRcVPSi9O6oZw==
`protect END_PROTECTED
