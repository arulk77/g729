`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCq51fwK7cI3KJHtXpVsfsD50PYaA6XaKNN9WtXU0Hcu
jM+N1kYyqsppUNWWBHIxI1CbkVfZck8HS6KWF61kfhuEcci1UaIrl39sKBHVAq8v
lwo5gRwc3kCYlcmhtxuVwYBkQlO6x4UIkXQWSOsP1QTk2AyV5UOBGs9B8Jf3VkFF
Nj+Mds0gwfBEikh+WvyPPwvmAHQnTmYAIDu1EA+sp7TOdcVeFUcY4Qo3S1tdqspV
++6cY82x0SN0qh4U3zxuXwMj/A6PKpUTOiSZ5k7dItwPGKjMRj385g7w7R6KZJi4
LHjidtJ+5kjscdIAVhNS+TGFl5a6LEfMeVA0nMfNUg6ltkQZ61NeXH1CcLPs7c0B
tECrL9Q4Jj7fzMnqumKxO2NUyP+XfBigs99YJOqXnH33YXhdmfCbOPLNZ051XIiZ
aukUo5iIHXkCXcsxFp1w2p1wptr9FlP52ddGjNfVW2N2fNaOSGoZNQco1v55YwtZ
`protect END_PROTECTED
