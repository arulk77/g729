`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAUE24FLTVyPJ4qFT/zzms0qu0I4sNoYPsCayYpE3piV4
FP/buJEKyWXE5VlSkhlRGD32nzUyBgx7dEKtmNM2QiMAeqo144Ndh9VaDyp3J8on
EPtLARPAGQPMcAJ0dqsxE3MdgYNCXSR+w7uAwvDaQSkqO8Rs+gmsOKzI3HbPEDGr
lu8Lvc9KNeVPyyuHZW/c9xeL9trEGpLVarHreJEoPDjncWNDE2CYXcfKoTrWCbWe
gmpsHVWxtB71lCGM6QsByWoPz+wIQGVeph8Dzk/94ykBBBn8ofjrPB8oMcgTdHm4
8HUSuiDPW+y4RAl9eWXwJCtJyynQVyVYk3ZCloJYWGbLG7lknO0M+lg1+v1PJaKQ
h4PzLWubdjaA5Iv8njV8399ut1DV0WGLtYCcFtCCLxAY4bA1XqC+BMvzn0UKTBLr
pRItKl/aD0Ge/1sb9eBUJSkZ7e+xc/PB6HzPGbXsCr9zYyIdOuofb5jFUbCUPUFf
HtpPGgeIkX0XSVIJUIwz8v519WFg3u845x7ePxzHzdHexATEI4UmYD5B6FX1c4qU
kW67l05pBdJ05Cr9TyaM1Nw//keutV3xczM17qbhRvxGglGFNaiuFjz0sgB5DiIh
FJkTb4eKKWFejo5Oo1etEOlBPAr5+YDeDc/z+cLrLXJOIgcLuxv9wgQCs7sp/GES
5pLnxgqHdLjAAUUhgHsVcMbLnVVAXTnubnwfM+KbPb1PZHHENyZeR4kS/IppLQNt
XCVXxA3c3cjNltiQiLB6OGClS7pdzshxYLN+eoszpQqNfFB/Xnlr2y2sn8hRZ9ql
tMSLKva+UXBSIOiFCf+0EpwlGTcP/vs35HzVymGOAAUR/Ts9O+p4KhOyeOMGNTs7
RBm70eLq/rHNQGRMZLf3j3Ftt75Skc62m1rm7ph0V3cnA5DIun8eoLrhW64XQezE
PWOFdQseuqWd6K68XN1AP0m7RwR/TvS+ru9iYO/HJqyo3Hib0vy5aPjJdv8cDr3a
hHG5/DEVzWpTDzQZUVg7nWDB4A0fJiIDnZxlbzErM6SwLlDCxGqzYaQL518NJJH6
IkQn/xmR9O84QER626yQhoIvo2cZtHdzQuhtmUlHWCheUzwbHNVtE0hOdWK+cRmS
ipbwOVOvmWCc6bvYU1LyBM3Fhtde17EqG1FMC43pBM27v8+DlOVK7BEZhlNOn8Nj
WFDJCqAOg03ffzGKIH866F1dfxVI6bcb9GdkTm1+IlnC/nE/Jd12yHh6Yqwv9HLb
lDF9R67eTL1HWoqvA2/QXfY7B9uyaax6c+YYCcNsuljGYtZWu4ZIFf3WMHM+T+Kq
OUsIqIFFlldf02Fclb7JxB+Ew5zqQ8sIQJUIO+tjHE5Nh7O9IRzbYIpjVeA5Ulb0
0dQD8RyjbMVkFF6r9rYuYoztmwd2zEObsZbrOIqkNG/WWaJlV6KVPDg8ZpttEda+
QbOjv/A/yU5AQPcLOrztMPQB+dl+mtLIgpVvp5bMN/xV/lWur9H2K5oJ9yuBL+Wx
vb7t4IU9h4zvJ04m1dIRM4uvapmFSkIHBoQQgxzeOKRRCFvkcVhg21jGCZquAehC
kZM9mPyNqSRi0A/gRVQI5BM2L83E9fPn14ItRY0gS6S9oo4Fbnj/AexPjwUv1EcA
GP9gK9sKqHCGgEkA4MBe/xq0ByF6VmMNZ9QMUEAuoJBwilsnmt+kHaqlgkv/ulov
S+2V2Hx3N8GmoQuv93KzbLS6zzChWYlCWnMe2cpaWQEuyM36gpPSs5/FnNdCB73V
UqdspoLqWMXcpsMM3x04gWd7jaFwqlK3KtAKwZd2SA/NOZgZWmV+4w62nNQsyrsr
YWvAvVeFXSSJiGuEKpIf5lOtQU4wqEoLg7g2IIVOPAeB/HKDVNiSqekvnbHfwDVU
sShAof1RyJ3L0yoZyiuAbZdHzm9r3qFxKG7ebPDY1NdPuMeiXyzA4eCKf/YZUF6q
mtgvCEW8v2vdMQ61nRgo5XY2PneTfV5l55CmI5ETDUw2NFKrxShGVGarHlLpvsMM
5lNATHAGXhgghTHopUwnz9+kFybkRZZrlDg8ZXviX33N6RIoTqQSTAd7vk8fl7AR
pgiI59/AssoT35v9Ed7Hzpm3BrGWgSVX/rAFF9RbT1SzyG8t/qWcYXVkrCGtz9Ww
n68vP+jODBgVY8RDWi14ZsAbDxCYn+iwapj499NbzpIMFgFEkb5AgSeMa1G1S9Wc
jdeuzp16RMlU/JZPzcVj8x6y/DYo8d/Q8Eza9X8mSuaZ49xwGMDi6QQDkBJxDW4U
cCI1jCN7ycQw+WnRfT9HL1CQsneWYJm2FJtD9RwajkY3odgiBb6+uPsLxmIWYTmk
md8iYv2moiWtsITKA4r93LzyPqKaQzFrvtfFU5OoNOulHwIJGqXvGaJJcDivtNDU
LpCx1gQPLcbB+/plC2vrKrBwC8UXPcDE987K9AusvfF7k4NPJIllz1dfzgF1zHbe
oumL5cXCGPFt3DZERDKDww7a3PP6tqdT9EiqOhBh1MOi9wi1u+HLrO7uB20BC3Vh
AyQEKdfZWogjzJCxANn/jXi4zRQsMrwihi5SOQmjLemllEGvn/4+TQ+QIC/zLXJi
6bC8owR9nwdvjhI7sarL5F/22KhyrfEHn9hd1ac4ZA2J6T5YRvZ5+SSl66DLAtuP
I/XRu4EVCFx9T3POHlGkTPRhnR2m1Cnn0ITsY0jJlq0=
`protect END_PROTECTED
