`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aVcf+8iC95GdswEEwey97Dhkdkw0loL7xVItA/BR4s8V
Ld4ThJa3C6/j1vDwFilc/VhzvPcnR+4wZ4aWBLchwUpMXblwv10gCq+jAL4snnyw
mjK+94kZ1uSVCT/8qc3LGg0OaF33Ytj3RAHk1OdKmJYgXYvZWC6XCKdzLZIPA2Fp
9F+md+MzbYav2h65A+dX+NJXabzELaeDl5nW1kFrjwIulRERWdv1+Vuu8kvOfaMl
zBopdin9BEncu+H3slICJAT/zt1MgladlxpcM91negPux7Ehk4/mgwS0X9BYrHae
T4U9+mtbgm4jKBVUJEG32Rrz4jgqcjlJ1o9q4MYwbAcHQJasFiG6c7iJ7M0K/eFY
saQkMobU5iiZg80Qtd17cYhnVflgCMmaSlqUbySCHeYqns4HUsixV5XrzZjf7Tig
3Smri9sQhsxMmA89mw0E0C8FNNGQ5qvCqJf8Jjkx1aZiVSQ0+7ahkHaz6EBSNpfL
1XhRk5cVZtMUcJvKhAHdkHlBWV7jMa5L3TzwIhfDnCcMuxQL4VNEaodLhnoPoJ5A
q8hY/dI4UmGyzvfU/deFJ8z6kJHcrvHQCDZI+ec3yzU=
`protect END_PROTECTED
