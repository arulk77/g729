`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIKc2FwPnjHF0WHBBQOHJ6RE+q6a1s/IRl0yXmWf6D8l
YbvwxPCmMQkmA6K+qrmD3LQV9DL4lqFtm89uwUhvsSbhS+Vu+fIDBGz7ELfI6INF
VXj5y8ByNh2N1dLqUuTK3r/jtoMXMWnz1rBlZcsevmHC7xhZrk4ARNUrGGOF9b3W
NwBRD7F+8WJM3aBegyqwRUQ6g3FVCdNavr6VPAs4gI2OKGCqWml0opaYzkmGmpBh
r3QW4ea78Zh9GAfFdo/y4MWMmEAvS/v+agLScuE1Q/wdidm5EgmwKgVTByKlKtzY
lAeF6OJwY18J5m2dY62AwhPomt3n7uAjM/xNp3i8C677o20HFkjuDs7kAnE45Xq9
4zplKa+TYgVj4yAk58w53Rvkb1z9ahimns8JiEZ18kIkUEkHvYHIw6FMdDSzurKv
QiLp2X+51E24kgjRDmyqeLynQ6mfrai/Nx02X9D4ZWSObOBHrvKK6Gzzhi/hgJNZ
eGXlV5jm+qvGrMTj/lKyFTGLvY4EHLmAbI/SLkf3Emljtnnk2GABgkDQdGmJgRu/
K+R070A3FaiMcvUqydgjjA==
`protect END_PROTECTED
