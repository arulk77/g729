`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxke/XfQsTQB0xMOuCSzFG6UOvMd7YSDiTugNHACxDy05h
VyGjZgnnh82NnlvQ3r7OcVoExQYX5xFIhmXEvQ7EEn5roT7Woz+Bq2zsZXnlLzaA
QYI6oYPZPHyP4BPz7aECulIrFf37gOfvvii0c4NEDyk1ugliy3mWTI8EJAbu1WZp
ogTfikkiV6bRWqd79tfZzW7QEM58onJijY32v0rJG64rbw1nyforXH9FKtMr7Smu
IY4eWbUh4R1x6WgCfdrus1d9Jh0DBM6IQJHK55LV33Kk+3lfxHtg59xzopz+6HE/
o9lqxUzsJibXDlyoCaXEKo5KoBDYTfSDuba17X4Cywd9V+ajXcNXdAKW1Pywn+Mv
xtrnimCVs/G11KjZ4DGJYQ2MWuCh/yS25Vfa2dtqYBsfpsPB51mlCqsWTyBvCuWQ
8lnOEsUhnd0yC0a6CpEGIBp70D1giYStBt95P3hd787AsNjAIcNe3KTgsG1t4eJm
7xHEq+ysSDrMoZ24ScILVaulI4KEDn0Aci0rhobGOHeMySg5btAUN4bK799/zVUn
Jmhj3gDCIztjlqFJDYiNaKoGYr072QgF+1hQSJdkppClz7RyHtRjwKX8B6HpcVyc
x7ZPIG5Rs5m9/m5JjaHEnDewACBpqd2oDptWtz8ydZBQBy81WVkTn5BDK8pxMMM/
kJMg1JDlIJLRE5Bv80ZfkXMRanLgHVyDLc77uCV7FC7iIFbcLGUkfXICxMBUYKoY
sgBCNVn9ZQ7xML8ZW4W6lRyhb8Ujl0tGQOZqCzhE+axwm0NvFPXwZwP5glCX0lDd
jvL6LoX5J3IvYd8jcEk0P9Eh3TltsSURGLYKgaYhl+UOeCFDy4gle3afZuy6r/Nq
XzgWYwr40vVbIxEdz0xKcYBmqtVV+VRcVJA9z9DNJZx2bfwUxIJVA6wmHm2Lgt5a
tQ0RdBD5Cty/dAaLnbp3CUHuns2VLhfbfMhD5ltcXOz9bn0c31IrlshTWXl8baUq
OYmL1Kg8OXJpmisy+NZ+hFbLazBtGSWvb/yYnnFOQcL04e//E88MW3zFFuDYb8si
azFg2zmFadl922/1waRfeaMhzTRwoU5xtJLGipl4SzHA3vEL6qp+AHD/DhD+WFE6
kRubHZIMvLFE64N4RhPkpPM1wQjOUbva+lyKjgpQyYiweUGlnxyLtZWuVzmMbhVs
zj8CAkr9JZX1s/GdBnVrGrv0j+2dprL85S5gKOkweBi4wDjQdYcOfEMmLnZch8/+
BJ196e2vdn9B9rbUL9cHUqAHX0K8yD+4O+YhKzzmk3ougVSAJHzkvnJmypSPphFq
K8Cl05u6cVNgxKmPgbVENLrmlh94q7E6k0FMSDNFg1fWVsmtwB3uq9rPbuEv5Wkz
NsTvVnjCERrjCsi64n9JWJqsNWwF1qOBZxqnZUPRw10LUl5tIAom6kz4u9Le+jLT
3/+/k7X3/chnVgzwBKZwZZ5nr1wlIH16nyDhh8YNXSE=
`protect END_PROTECTED
