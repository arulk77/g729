`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIX26uRjIaeKaZ/RiBdbt6kcXdNcXjLiuKLVeUnnRYrE
nzWhKPoKMw2fXZJLpgzv3K4KehXACvTTLSLlodQ9PZKQsl7IGg14LPPvsw4kQhm/
A0Zh1vadWO/TgHc/F7CI9pFbvDs8ToI50IrhTU28UgjXPdDQpuqV0qjm/cYu/pCA
wvwXwxvDZ/1n7fh+EKDvCQ==
`protect END_PROTECTED
