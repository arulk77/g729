`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB0xzDhxCS+bH+mcE73FQ+7y+pZVg1U+9E4E5CxFXreo
8DCIJigWPJBhA3xi2hMwIjVGylKdIQkF0U6OT4QqoAVmgBlcEMCYpx+m97/0pP3+
+HGqLRRI3p6LAAzSgmMpMEjCpcwVEULafy3ahty0sZTpTKwqzsydgO5KFkXjrg52
kFWmL6tUVHuEDUImcVJSZkgEmmLV/sm3AoVZLup//eFJgHOOGnmCQeYXsbCElPAm
o1YcUYZYl4kR7S+ERrcVU6X77/vb8PoCPDw1rQuL9ZR1eQCuozVIm2Bi52ZwQr8B
MY2OCYbhqYS2Aza22lYX2O4YQbdM4xA4QA2rf9x2Rpsj5fR6pDLDmtiy526IseDk
QPXWs43spn/HL3oLT6usAw==
`protect END_PROTECTED
