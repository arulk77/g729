`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIO1a8iFi4SFgIzPufDibnZq3GHwmgKYJpde2DxhRdvz
IF7AmU9Zk8pvgm6D7nwg+zIhrrXSpRSdLjJOad0eyB2bZWp5zkpCCdpGRjVygi4N
O46pG3VhuJxIW6sIXCX13I/eoiBVFxIkLd0EEpYqND58ARai/RHEYiTl25t7Jrg2
33QUoqPTYRZ2dva/XvNDv0dO+XW1cy0YxrfKZDnq3eW3dVVidswsqQm6J1B936SP
HtrE2DSA5Gu2fBBBaKbiIpSTpO6Bsv3OVw7dumr4V6UPXb6FXS/tarNFMTgeuyyr
gYAjWgQLMDVcDFmOeUkIIMYL2qnOTAe9Lwh36A0k49rdRU/W9ZVlhr0psH8oYeWC
tXiDbEzgt83YmZ6QSeMqkAD0jVX0SrNVG9PPkDOFYvB59MiCYUwDJseBUkQigdoL
41uwZ0oNWcuS/ByWnc5BECoR4rP4VfI8VSiYJ0R7SnuBqfw6NEQgXxMdb+5azhs2
OmDB1h8mfzRdg2NbIPKIC31lC04+L+aDGx7ryX5ANpUFpNSM/SDog53H5TvzDuYu
`protect END_PROTECTED
