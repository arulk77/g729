`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
zPXP1ERLoOlbciZaL/U3wNriO8Aldw9mzlz8vBbTetSB3Rfx8gh4ivcbovMGTFkt
EkSRHc8RYm3HR1LVe/NvQhmBFx21YWyIfjlPakhMZBYplv1Rl0zlXjKuWyPCRshh
CUONDuxUEiIceZ2U2xhkpuOtavNbHgyJ0eHZ7rfGTIwqibDcJeh0NIVoW0tGrrg9
iHVTpaRX3urlrBdas2btcy8V7hKwJDt6/NvCl0jA0Ov4PdwMvXaoeLap+dKcCDl5
Lj/Erfob+yUBuLAZvwqncPLNI3w7+FdQwQp99WPjcZkA1wKb6gy18XF+v4WemwQk
fSZpKiidhCJWwHr5Nwm6gzyiDdBIvQcTlhIXNwmxW80hEbCG/2Iqr36YNpz1J3oW
EigPpBgxx7tTAjgbvdOhRGEH4ADDBT4DsregHmZOPzwJ4MIdGoCl4GaZDvk8eEuJ
0eMByR6M5gqRDpBzS/gauNCyqHD0jCwEWUCAw62QccE=
`protect END_PROTECTED
