`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
1DWqYZTEBJWw4OFvJrLVKF2TsJX7zl8aMGOyNZ1+s3ZLH4U2nGq5uLroTiieqOLq
JJEA2+59aRNuxi8k2DrDfJx7PBaCaPiAGyRyZ8FSXp647RfHXTql4uR62ZRMDBKw
LGz/1cstroG0goTYxHugz3wVe5LocuVyRcWxDyiTjYr1jlxPCU5lLo1r3VKGUTfo
iQzesc6g/QUZiY0EY6JtFjKGzDayU1rYn/P3SZ9+nwI=
`protect END_PROTECTED
