`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
lBkftj2DKH1qUZZ039tg2Hgk9dOg5zjIzyV8WZ2NjbX7dFMANwi5tSCa7qPYT7TD
29zNEgCxqObOqs9ZOCfA4ABHRwYl9Io1dMMs+17vRBKg/K+NvYtX5Lv95FrPHHC6
HF3Nowe7PD62uAC1vBBumfRzE0BNt51rvJAdQJcm85mG5P6xgAJnL7Yo3QvLF9rc
QJDWrt9SFxGPEaO7madtdDKOdI4BIBQpYwcFY2PjKcUUkpnnC1nujzesIyEVKcPt
yj2USgQWquvd025FtNlROh5/J675nxmHx6GTRAhwhMYvJ+y76XoiwHVtdabhbaAq
qNcTvRA7NvEZNumykZr+avk1QQ5G9gqYwWEQCGnlNo9RqA6BwND3uaNPYZd/8p9t
VEb20PuVGwJnrpoGb9PyPrJdwKAQ849HroldfAMKLFk=
`protect END_PROTECTED
