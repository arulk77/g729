`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2RtTiaLwZbJSuPbraFO4dvprLBc9dEAy5Cg5QlOCGZYIIV7ucsGRXctSLKpvqMEo
FCWTGj7wBBlU84EnSYvybLSu0I9BisDdWwdFLTTLlwaDcf/YwuFURa19wMDAhq4m
0QVwzHaNx3Rosishk8xC1M3uCzo6tvRwLjAbwSXLEfnLsPE4H+Bim2s57H8DOFVc
`protect END_PROTECTED
