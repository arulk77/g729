`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAbgV3G6L3AOINudHAeRMJx/hKmXOgLUJU+iXG+otuvXk
/zu3TlO4MqT6XtwzmaytB05VIuAAu+RD8UymytTsqLiA+MLqvCYa5VPOwnQ0Ona8
NwM8Wcs0MuaqrEkVmntaKl3b+xiy+sF5nKHQ9tUBVf8+PV100Bh8SmBZdNXfAJzW
3d9Rx9+36WFPTYAPp4xXcdz8U38hPk1fB0d7XPMt2BUZ+2nYNHpYCrhiynjvsush
qMX0VBMfMWK0VHZ57xZTX7Z5++rpmMkPBRU3YT9n6ZdUOUgeASSryY8F+WPpBofw
3c7UieTbLPgbzkf8KwQcWxTHozVu36i1ltRqIHMp8h7vmI09j5+yysMPLShb1yaz
qY5zX1nKWlQqDnQPN7FguzTjThgxEjArfWax0cODzUo6G47S/vj3ytRwJSnu6Y99
uEuqaZyC1NU5UTsQIPNK9wcaFjxgvevwcsucEAxNtGibX7Nosu6jMHb7uP8qLOOO
/FeiJGX7t+6oi0UgHCelVy5W3wvUAbjRFofkkwkb2Ah5tUeAlsoxmzLXyA9TU9TT
wOKP0B0Id653CCtCyqpZpH9j4QbIkYTm1BSjZmpZpVdYdruCGJuBBzMHnZ5DlWWs
+PkeNCxTu2pYlsexZJDxluBzgZUlhWKolagi4CIMQepB9esuN/iJ34UHspLQ8GHt
2QpOJDdMeuGYM03ZJhZRVw==
`protect END_PROTECTED
