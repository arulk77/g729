`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
actsLePZv1OPN251biLTaGzzPsKJuBxb3CzqmeYh+2O5qzOyh7wPCfPqR3a4kayq
jmKAnr5Wq5F9vS/gWF0fJK4ZPSkKHKDoQBJ9iG57XiOwQ/Dlu56uYBeHFkzJrrnm
SeAZiwS9lF31v2Lw5ZfY9ueKupMAH4hN/jUXhG9kZOutSQ9JHxaoGzXjmbBbNjsE
o3Y1v+EFy6exTM6EcULqaWuVisv0l5cNrAnDjYmb+bIWt8S4t264+txOZxujOCgF
Xi8RRHcR/Le/WGHS2KR1qYp5FVpNp86q5uv1nP9Vw3tSpqJBWR8Xgi3eKuiURul9
twy4LTpvNP/dwiJyfQhtDB7Ve8u5tv2Agx0lXCFbkgo=
`protect END_PROTECTED
