`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL8yXTOLlckASVZa83C2IVOslwMxKcQGrz40uIeycICOwf
FgVyI1gZGoHskEPbclbzYTry+6GdqQdLbRFazMv+vSgCzJyRb9DxOAb+fWfs78I0
cyZwiExoQpeEAt/kJcTh/0R0JarLaRG8PFoqdMhJyGwa1SJ2e6X274U7CQEyFV8R
Ral3L7Pw5HJqsaZ87iazgHexn9qPybBu7O7oq43xpa1SuEK+Fw56B5aDBYjmaW58
OGqTkiwURpsQNT0jhLufZJJknDRDtjAVZZRpA+KQgTolhysvxax8blqopv57HbAo
hcB9XiIo8PdqmCEI79yxn7K1ctMvC5le6PxhiEAjUeh/7t0u/K297fy1/kgX78GD
mPwq0TBbXiSa/SMLxbtV2ACnouFsu2weE7Kl50e7DolvQwvr0JrjKyoN9peEq1n5
C0u+HaJ9BHVewRF8gL45lQ==
`protect END_PROTECTED
