`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveICpKyl2ZgOCWA2dnOTogGXdSYSumEaviOxfT+mwG1cI
V69t2RlGhbtCcIDl5eviFjNhMv8ndOSr99bXmECtaRkWK904c4MgghU5SiAamX5t
ZQ0FEq8xfAPAHJTZ1ssR11B9GpTDcfvnNsJDS50IUiWayl6BF4yKAtPilnW2HXHN
Qwy364oF04L64jOtlzbDNg==
`protect END_PROTECTED
