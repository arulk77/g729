`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/s7H+kvgiuw82odZqdsTKmK+Dz83NeS6ub3yaFxojUS
dk/wc8RTWm2iyKjOtLsqekXRDlTUBazOKTIFwVgzSDnPd6CsJlxte4e1VHGa9JLc
kSqvgjfYpM4IZDS52JS6hfwOVKEuXHRPKBXcaI+9QWDmQXeo4wI6LYyZh1Wy/WfA
js1ELJ1FvVHcZQkGexyetnrQW94pPkcvxDacZQvFZIPInWPF+WKva4zjovgkVhJT
pxpUJvOSMszMxTtb71A1o42zIqvPizfwBX2IHs519jSydVYZyjPBAkgjf/F7jbbZ
+KIJBpL6FEPIQCpWsmPZPeLrz30eynjNpYvqezX5D3uFzZu0ewhQY7ymSES6v5dK
0kJNDsr6NcC6PsJvZHDq7w==
`protect END_PROTECTED
