`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2z8yBFC9JNcyZQNRBrwtFfeUfkKj56Bqqa0d2ONnhRMAKfbypFT20UUDii0HtPYQ
d91Ej7aF3/7o6iWGJqmL6Ssqw6zB93fZoyxRl0qT1D7vLmQbRieqhRRlZWBKgg8c
d2DG9RLPFk1KVAHHKxexPPsruJigV4N8ZyJblkQ+0qdToAPv1znlRP45HxgtTlsI
8uWahr/vH3phU+XA5a5ZHVt+f8bYw4yXMp/RpyF0r4i8A/hXf1xargahkQk7c5Im
fJ0rXBBWCjPQRAxAF1u6DCQmJ/sZ42TCbxNk6bARryJ5tK3CFk84p6G/vARdO6yl
B51zL2hmwhF2KxPE8lsG0vQuTok8DuNxXzsd+g34OmGTOo7FahzF5FZBpmvdCD+p
QqD64Mm4SMDbAC/ER6Uj6PTRdLcsEnLHdpWks28xxt0VCl9p33pEIzfic5vmdf9m
pY27ddD7VpAXlYLTtt9OL2JPQCEOGGYgJ+IhmIIZRdRFqgWB8QA2PTlhR7nz8uOg
lCXACQbpi59QaFiRWR/zCv8Z54JGhelOFhK2pyFTdjjVjixn81T5Kwre/ubJZmNH
Vq8DdnQId8CUI2kikjBICQsBnn/WPP7Qg432DsDLL9WI6/Br4aMBuKR7w/4rpIFa
U9+8LMOy4jKAe9sU8cZp64CLFt+ILyLEeIoBJug8MfSsReRueVLbz0uYOZll6TrJ
+jCO+8yCMmXX/sz65S1jtGOXDCSaMiIamH6FZgvzQ7JZ0obDlIsg9dMvBXWQ39M2
`protect END_PROTECTED
