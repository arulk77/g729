`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48BxSzjSydb5gSStAyT602QnRxTAzM6CDkC15BrhX1aG
sRzPW98o6BLFo8ttfp06P+XNXQevuxbtvmwujfvJAWiWSC9RCUf+q7LMJCSHxCyC
sWra1ZtkVJSK/TR+ZlSkGTp/POPTMj1XL5WpjiR/k3/oRwD4KBMu8PGB/noBh7Ol
8BKeiPXVpNPe06F3TLj8L7pNYNn/FKrPAnD/gQUrdpNpYj8xbJ7eERFtXk8R5pDC
6YL1K7cYbj/jO6bActhD+l7Tut+p3VloQlSXmvvA/iTCbqkv2zskBWlLJgn6GDMl
HpzjEZ7ZuFkpoibEZRTUAPbNWRmGnxhdMTNyyXQRktDbPGAj0y0r+5hE5sOvEy4G
ubqqoR9UEU8g4/onE0evIWXbPM+5Tlyk5mNneC51vhevn1iVDne18CBQqIRLAqtL
L2MD2dbYMkBeWkDnhtdEJKpE//XLrGlZ5bojOnmRqvgc/E7xeK05tsSVrj30Tz7E
`protect END_PROTECTED
