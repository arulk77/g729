`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bax50QrmXhkrhnhf6NIFHwyVxm9hXaiSNpcqPK2eVMbSb9wmEREuYgK1t7x9S0Le
ELBIpnW9oxzSAfiZnB/Mcz0Ajie2NEOMy9xH/jLSE8L0H7BFZie6LQR3Rqo0q4Gv
3bLtZkc53I8JDrRIVrDsrs5ri/+Cyvt4IhUP7WhCWe3mdg5uG9SVHi9p1hlhWHpl
I3dI+iBjdIbDBKRCyUMrYaxLCgJxalq+wZCq2TuE81KUE178Ef6jKbW4UUtg+KCD
CDkD4KsY9Waty5P2zjtkqp6VbRk72g+U/+2ErowTIE0=
`protect END_PROTECTED
