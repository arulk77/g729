`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4ybyBM2PvJkLA5UU/F4L+OB2YaRO8HcxrJzMtaUJuMKR
Vj0YRbwTdl1ia3io2tKVFSZjDnqZNWpGRHj8YyG8nubgbI9h+ZBdeYyjT+9ikzqI
L53WXVq8go2P+2PHLuGKQmwuLjBQzVBYBZKn35UIqBgKegC30k6evdIjK6tc5bWE
8aSjdF3uiJ8HlzgZAnu1WMYV6R9B4JELjmjTqvaOgPztszlqjkzvTaOUUsIwJR8v
r+XHC/wZx3oE+NFE8X2pAX9UJtyRtcTY5BHqJu+FMb/5UVKoFBveYdjWr843H5ip
v9EfI0pUELAm7lPPm853ndhkJ2rrLgJqBqYMTIZiwVlSdHF6dfgsRkey5YiuMGy5
6m0MxsFcsp4p1RzQq28+63QXC1jCXj2gxjxOW/yYVE1OHwG7A5dUdx65QmL+bM3h
4iuWHVnhTgP5fKqpKQmbmQ==
`protect END_PROTECTED
