`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46TEWSkHwAk8CnEepK3uJi/in9X7p+Bi8jxuD4yvQT/M
O09828v0GDgEyi5DqIheVSO8YekYve42xDKtV5aye7XbByPkQ/ip1F7TgG8UoKBU
NO1b2uQDw2sklgEgG2IQk98+S6ZnBA+YdqxiqcvOhpNKOfp5QUMxwqw3jkx3XQ/9
s/3zhdzeU5O1dj2uynoN1O/UQco/uNU5ZS7MyoV3rEovyXu+Ypl4XfAtiic+au74
YEmAx30fuqHcktpZnEw0X61wJ4ejFVh8QL1yISbckHnep9oM4S7On3uRdGmqn9e7
XYk+m1eYswjFbpTa4h+7XM5WY7lIrIfrbiquTLJRf1rhQHrV/1rJwaswY2NT+Rq1
IQg8Aiv1kH2GgPMyC5+L/A==
`protect END_PROTECTED
