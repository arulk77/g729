`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkQe74wLhP+OAsCrn7+blV83pBx7E0GxxwjwGxIp6LXST
UZWxkNvnXic5kZkaEpobiQOTJMHQWkv3oijds18lWgwuYM63URbJNBZ7uaiHFC1/
oo+GxyCZejSInLaROzWlv8Vy/6tGiBu2MObzHOeIOt7JYRtFg6eqQgBJ+dpVakoM
Ur4rkUUn38jr8XZEFb0T7dLzsNIWQT/FBX4YX78y/t/gARUZfcSpANgK2L0TQ3fY
qexJCWN4vDkm5oB8bC2Fo82pcXrjazbI/E/1NIIXSWuZwVg7UDTD/VE2SH/hyMgB
zN1ikbd+y7Qr6Jwi74QE3ZlfQ8JilUzl1cvR/5W/S5j32fr0ewdrGRSD5Z2ddFJC
Rrz3ibGKZ3MblwPX+Q/ckQmxOjcPIxFzP3k8j/lBCV3TB2c0j7ElOJ8o/HmmaWzq
zqAM5lp6z6ya2HesJu24RC1gt9KKFiuiPEJadU7ybnXJ7UFVpKD3Ek2BmwoPs60H
8DDNnJ7f3GC8nXB+aKlEQoAp40DNirN6MIrtHs6Wn11FAj4Xucqbdwv6FeNBNN/o
t5KoIU5bpXlb4C+SpWkawzAZu/ffnUOdc3H1MoF/0mvbHkHiNl6Jci6833m5b0TD
AJZ0X+nR/0z92PO6CEJCGFWc/u1/deUBPtxbgSdQzoit6N37scOTUyZje4+uYMGV
pZR8vwXKtRFu110aGr0QlJzVeuN6Ie1wlBY1CPI9VQzo0WyzfZ2MCUxO96yhB4Wn
NJmRAtWhlLx9GLRIDMErQYqqy7DyQc1qTGK60OtDSKCrmUOkZWOpdqQAzvfitmWb
K0/WPcVYhkWoBufuul5mW6N4+xq+Kb6LB7z2rxt/NmdlDofZDx1U6cn+B3mIzLt3
x2ezOeUzGZEvFNyPEYPI/+KVv7q5XZZRCMdaA8wtBI1LiWKO8K0Pr/v8VZwCfH00
3I6zukslKNhtKow5yRQqtKQFR5fOT7UNwVN64G/xBwviH2+nII20qelGiRfIsP5F
/Grvkx9KrX/8PyVjizJaHpGR7fAZcsyri84Xy0lQSRSxZUd+feJMcGNpdvTzZvbY
0aPBkDhEwiXAk5BQFD37Qw6eJC2pMszV25fZBExi3Tt+8D/eynQ4eQZngKulRLUb
NrAB5+MK1GLf2iVK0Y8Tn8/R/ovIYMPBoXYZsQGF7FHJxHrnONs0Smzrs/IIUYRL
VqIdzHnGpv25rpfMydErNTI/MpZchY4OllLAF6+hCV+FJe8bxni9MzkCNa3aqqbH
QICnAJUdRMvwRakVqjJzxyzlUXyY2Dp46lAF64BdQAT37K7RiWaKJ9jFWm3Y1VUD
fHTCnVk8qXTUV3C3COLSaSsNE97xW3GoPTS/OarOW5jLijlZexO/JHFO2XuhEscs
WJIGlZq8Gr+H0pJIkPdGJdITL0iypc8sNZ3OHo7VR3j6fBhLa5fgA2TbHd7t7c2q
jyamyzcHhbM97/ZQC0Z/EP1PdZCVf9UMuDzOkO6y4TICjfk7c+zts9FP/iddufJB
EOu6qCJPJac2tKHSuAzqI10hdMJAapEniUqSIrIuHrwa8QKRTH/2UM9Hy8JbY7B5
rzWaXpdRznf3mtZc8DKtLKxYHjxEXgZtgfgqd5jxDsWT/TioY4+KOWVmod6Pidzk
WSCCOjaYMKclv9lVgkPA5RU12gy++n9n8Kh8ZaIDCe+Vf/14obKxfHBopY3FIwf1
AOc65a+AaBZvXutZ258OH+1E4z1vYw5APpNA5OxWhklBCH/J788DLhZwHG84yYvs
wu5bfn/MrPHUGUn44WnjLfq+ohnojb4xFI7woX4cZ6B+eBjuCzHY+Ak1UJAHWIID
zEzsGmA1fq0NfT6JwbGjwerOSub+SfADOl6BDBET1z3Ks6VbUz4kfHBhMgc6vL/z
2c/2IsvJ3omK5X088exGIfDlf3FEj/JT/dcbKPr23vIx6vbDHQsdmNnXDi31aJpr
22uKQXKgEVo4VQFSMfQV99tClMKl1N0M0TNkTwfZQiAATqFSyLJldVGHbCcFRs41
bZTBCkaMACIcAAfzdQmfgCo6U7g87o8h2zRoD6lQjAh6coiruUm6pH8BA7rfpO8V
qLjQ/mzEILWUcXpiC17LlzwcmzCisilsjQP7ZwqvR/xbuxO19KYucyA0L3xrsgXa
+shb4IpAobRXFdhwkewwpeytdkEkI0WxKe1fIytnUkOdJddsbd/DbzPQ07hPViQd
G9IA3uV7XaDykjh9CQTlGO9jrR6N1RF+LRTmvBAmE87/ALyYmbgfj7cTcUne4Gbi
HlUV3AttT081xhME6DGi53x0D2CIBSju7GPgiZwE4XFWiVJZIuoHkteQg7w01r7Q
w7srI+hwIxTvcyQ3691qA9Ag/l8X6sRHlDz55912uWbwyuFcXea455pqu/Nsm6tF
c/wZXoFod/smrcS0Jn/JSI0H3YSPIxiBL2+VZRrncvKlZ1BJx4ZT9lvvgjE4cdzR
nTDGSbiHE2dG9Wmwp7mTVsZnekxN3u8ydGq64v4BKzWa4tf5xJKCVQTKm3RfQmvP
egVu060Gfvb7NofMGdcix3QSTLdz2jxq21FAmcQMsmHVO6m1suw1wFYIq3DYEJY0
sWwYTC1M9XnewEqxIaXZRq+m6CZ4wyQDli47vTZqdE889g2SVZI3S0PSIUPD7xg4
K7ELTjPZ2d3iinVzTcslavM8/rs7QFqK5HPx5CUgosCMxQh3e2SRBQeBB1k/8Ptq
`protect END_PROTECTED
