`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3cIP9E1nepUubGBK9azHi+T2Ta8gEhDRDuhlmEihAM1b9D7Z+EpgRxiKDVCs2z94
VAnKY4v4J/4958hgyFL8rCZWIi7Eey98eGYoyICJrqgD9S39Yn6PfTystGeO69Do
dFmsjy+53faM/g3Ua/nsPJR/EJfivz+Hz4xW7uly1w3frjvAOX7Lb3/rmWoPrdFF
05iGJdN01MaLS+5myoIh1wftwFHbgP+jKXhmvR3vmDoor9kTc/uDiVhKNmMRNtdo
/sx2Ps56AAE6BgZExW5P0AUrCoJAkWS4DuKjwDyfse9uFHE3zCg6ORFyHiT9e7gJ
kQV8Ew1LpBUH1l+6jkQ7BmqSCjDAMn71sSZKM/EHP5uO4W/ujb/JKEFgMdDgEc2K
k9Xvs+qhFRF234XohrneoFfVNRBvUvgm3zcaTgteMaT/WcutxH/NIuHufy1w6+KO
+UWz42U8rFEljZHVilvRI2AKgp3PA3dcUSxPE1RfSk+3SoRE4T8dieHwsPrCuuhI
o3zrWhNagjt5nuyNqaqth1YI191ZZXkLiH8VQmxsaykyB0d0hrtVC7EBroUAN6ev
LuMVd/RAtyFYkktodTM7r9zC4pnN16zJhWoWyZrHzuRaK2+hvgH9eNMi/9SLWYfN
xDHtfNkQ+jvO2YCBEc/LKNH03qT81b6E9p/iLGxG0drwGzuDHRLuZFbVQxnePCrR
Xl4Xdoegz5Z3mhHOHimPZQ2KxBKflhQxDIRiwLjZJovyh+0iPZYMBwdnR9vEDrUk
AVwr4P0EPh9Xs+pUeBL3oRKIaPnVNACuy39dJRqkkFGM5+9DZQyKBxb8y7Sc5+JD
8/Uw+/i8eirUDXKDO9AimoqCqm0woluhz+TEU70J6hrtInKeiOz2l4EG8zcTu81U
6TRY5cFJOU13VOY8rRn4Y6nDbuCN5zf5SWmSSG9oGY/+Sk4cRqknbknJGjF57Mye
ojGzqh8ZdZkhh0unZlYuLSgm8uwYBShxqFUB7E5E86S/NBAwX1uHYuCpc/bnMgI3
t1UQgTesjyPM2JhLWdourQnP5fzTDqUKdmatUyRT8X6MjvmyWUju6LwPG+/94el+
bOUTWmKWeQKksa2M5IE4Z/O8/kojufZDfgTlH5m6T0rSjJUxIYmlSCRnkNsABLrG
Pc62VScM5pHgbWyY2x1t5E42kZwIQJ58RnsTLZMO/KWYwKtJQlQ6zDqWqaYWAL6x
hm9XgfohWiVD0vPNz1aNGuhOA/qdNKDveAcdiX7rGISLmnB2/q+WuV9WPVW3NZ5F
zRlkcc3gBkDkvVaV6VhTe7CnL62Ct1Mq0Vpv9D08k1kK+lvX6rXTsRjcyJ20agtt
7w0HKa+kxevRAdWqo8VgrKL5/ZjkQaRdo2v57MzloaSFjg4K5IVOdVS/jIXIGewz
uawZdXf1ni6oq1XdVEmRbEiphe8CVEYOr1agQ9pwvf/XN5INBXIt4CmZajBUSGWY
S/ik8dNDwWN7pQEkosllND5b8S6/d74AAEgvqVlyX+1yiauJT6QA4ovVmckmBxum
LFqWTONJQMS0f041Ga2R6/wWExwwYZBwOi/o03njHvUHQbbKnDPCwtdWaKRmRoJ5
fu8MsP586iJ0oMhlzntdjeeLRQnCQ6+9r36SFhXs1V4=
`protect END_PROTECTED
