`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNX2KPDk8DxkV7uDiMNYYmfDoN7m+7TaEEBWI5cQrxrQ
uhr0rnrt+B6HMsknPE382I0lIZI3pMxoxXXcx7k1xhSJBOLJzSsKGrX+Fm36m75g
weu1BWx/+okRvhCaMnARKUbNh1Pi+bfsQX1wIt7hP5mXhqJ+qs/2Q7TP2aO2RRjS
vhSjDaRVQ2i8d62hfdIFPUDXNNkzPZGlQwdfq6rfqMTjRpds6Nv7o+q8KRbnXo4c
`protect END_PROTECTED
