`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePjHPOd8QYJ031AFH6BBCZfSaAcbBf24gfs8XywGXP4d
+f4QLiMsabL1vPnsPNZ+pUdGcAYy7Ph4iyx7zNE5tNIlEvDsMpijBARd4/4fpKWB
4X3SrE5PDXBGUsXsGjfCbCsXLreQQEt20rJQ5JNEyQ4ijQBORlvbqG7VqSlsZ4+k
HijGVB/fArHKr5lh3GyRNkvuII96Lp0MjsCj2iDOeSoiyKhFnzhLyw6XJUUvimhn
cfb1P090R5AVpl8Zc9UxNtkvE+f7L0kuQhVwzQD6sOxU7W+n2HAWlR33V/QJUZqU
pP3QCnlIgxrnaXMJI5TIbKs+6T/omwTFkvsH55W2eJ/DcQxq3UGi56tDnG07bRtv
bDFoaKk9IEstJ4zey+diTgWbbyVGHFAZWAfGxTF0EM4P1E/KJMreLCzf7VbB75C1
GWignGB1OzsgMw1VVMtoN8q64wqZ6R3xjgxgiXZrfDpVYGH8hNYVFKZdVoGRQvKp
3gpjczpayJYHJBZFkW41dmxEjB9Zr/Js2V18EoqGk+O8gyo70i6vhJ/vshklzc9+
oxuD2pz5xflgL1fcGU0K5MLgMqeGDdYKG7oGGLqM+u+TEf/6tA277pkh6QQWVAd+
VI5sKR18XicGtVg/9hTehVW7NCUACRKP7H8/aGmhNBRff58R3Kkh3cAYsUoMz3fL
zg5IHgN3SDuMn6CUMBuXl7HtOtPLjxFhSd6zO6FKTQYoG30j/baJD52L3BzVGVET
cAQEbSd4da4Cc0B8XPMGnHtghartz6hKllN6TRu3MJH/1j9roBVZnD2MM308EQzv
VaRw3PFgLlV2kCH9CxrUsTkHY9zv/KRbNSLaHiS9M+6+69ia+acNWSNT+DoEgn9K
DBIxfyrgIVjE0PYtYV64OAhFKJFz/TYTPRK7SWIDv9FJdlVLGh0qOogNv17LOxeT
n/fVAXk4DkYv4rowJbJHvMMdZXvDLQS6fTTPWFOPY8qlsCKL/ZwDg2BxicB84vdH
OiCejasZ5FEccZmexjmWlPMdL5Wm6+RCjfmeA6w7Sjv20QCUEpMXFo25Q3UgeO5X
XdaN/ytVTZ4+ufkhMExSQx+pRvdd1QvW/fL2Cg0Z2iG2eU+GMHqdDlUwr/YsQIaq
+GrXBsgtAC+lHIowxE9N1F35YWBgxljUvZqn2W8VVcQu+wZ/5dZLfRO990LxL4UU
U/Dej2uZDvpqBnUuuYKcjDdYQsOPqUXiYiL0MyQDDeVmGMfSfLa/2v4eWVBB/KAq
`protect END_PROTECTED
