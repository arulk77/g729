`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIs6Ow2ZX3ECQwEWEhtYvEhYUTTMhBK3xQYupThXoAKU
CVp+OTtrIZbQbBFrkJNK8ulLhicCGCBUQGD4pIWHb4Trh3uKWdMmHwtox7RsSwj1
RAXqsNp8x90mlXhdhLBb0sEwKkpHAHxSveHSaDqi0h1feGUg3sfjPxTTbscO5eDZ
K3K6cVGh+fEEjyRbCuFT9v3Q3ahL39zPlhwEDNhycqvafSfYoX4xOR9Yqa9zBdoY
AUB2SUGD9OPbpn+ChkWcEVvqmkqAHcsBg2zuOL5uLzX9mbBXHBU4Wpbhdhn4AKeg
lE1tGRZAFPt7WmcWZBirjst2r38NkOU6EUw2GVlsl/GGqI8ocoku+U4qMPGVhM5j
BnbaQ2hCbPco+IQqyFvi4wcL6UhqjF3LL09Yw5Yfmu2l5YX1hsHWKHDXdvF75GJE
0KoomZZw//mf/4mQ6TE4eY6l2kzzsTMEmr5r+4QHI3vQJTdXJCSyHv7OqFt2iqe1
TOfnQFJY4/LyLWaiuxJ4YssZYC+0f+//dXP3uzPEU7BQazUw3h5IngO0AoouWZiR
`protect END_PROTECTED
