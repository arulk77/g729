`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN2r5JvWp9KoOCJeXOwL5K5g2+12ZvWe9i0FWc4M6atb
6kPku5GHzDjnmX0BDUY8JPi+KjNz9liKyw5RwGz6VUXmOUN0+C411KLmEcVr5QzL
eg7apHRjk2vzqnclMGE2IE7exAES+ORJNSjIxkp7YL9t5zUDD8MhhFd2qi66e6SF
gthArpx617ON0LSM1mtz6NALWWrtqont5z3byyknT+DTSrdY3Ci0sKZXBF+rK4+5
kn+808aI6WHof0sXAF6abSxNKrJfC1swQEWk4sQREsrMNTscKFMsi6twyOl668pt
48C6mzvmm0fTcvP1rICZhA==
`protect END_PROTECTED
