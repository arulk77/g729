`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIKY0cJoSuT5DZkkXt99ZJ62CRmIkFeDFj9BPDiQw03a
xGSTJwDaccM7CZ4n6Vg2YuAOiFHtzLCLH8DylqnvRSWKDh9YlHCK1EWVIaJtkgvS
wOP/vHxNkydxPcyOpJCi6PaOlwU7eWY2cGx4Tb4edCPJm5nVVLoIFdaSF2+9Q0DP
`protect END_PROTECTED
