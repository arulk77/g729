`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Bt6nj+jpdu9Ba5Dacf/iby1gZGxU+oHMEOVwTJvYVE/wCVLdA64LLfdOV38xAX4J
g1+YPV2A/rdttKSbv7kuUE9alm/aX+35Cm7udRP2DPEFMVcFQiSZuqXv1Rvtj/l/
zIcKMp6rVURvIKUDw7vxEhPrUJX2b4Wn6D5H3E9w6BfnM6xpT7wM1ytZ69N3buOF
`protect END_PROTECTED
