`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SaAhqAVfATW2oL5XbhFINdbGEbbpzERkGhyevYDy+Bfh
qkiHZ06a++i1PoZGp7UQx7ypQ/XFWdI4VcQEntSKtBniwOI89lTW7xz4f4+lkk5J
e9ZCOTw4KD5BcCEWuoJstdNYy3kAklZyWF+30CBEZXS4jkK89JVB/H5eOPgzFho/
Qhb3IQfP+hOVCwu4qbzgAvAt6Z9UQqoL4zvUZLR+Gy5eIWwzwW63DChg0u7bd/6S
l+aNBrqQX4+egDN5MhPicLeGBv5HRGd+H2OLGpkPZtim9SoJOIi9qvyqFL2kP/7k
kvX0KiaVCvVaAKb6Ga2Smre3gchK5kxcslT/7uxYkaThzUDG88237hJzgehyF3TX
YaWmtDMhdUJbGYJekyThjYJgmgx6/wmEjrVySBGxYQEZGVyT1yaYxewgEZqMvnjU
eYxGRBQabp75MavebwcaBvAQYGrEF+CjtHmff+pWHmN1z46nWa3JMpVBPOjr0Pai
td/c9S+0ScYSRaJrgUfswCJOsclzRM3s0bN65+KfKI3Y36mMm+Q5xE/HdWQvYaOo
wfO4azKzn1SwqyvM+ohBmhVT8jBfiwndpQHB6XzeuB2lEPHiTvgVkc9fx7KK00Oo
+voGb9qDkBuiMU/Mmb2+wPWJp0m5HBtqCxCCu8NmVRX9Tzkyp/vhDE+VWWbUachh
hTJEDDjlKO2YHO7PE7kRj4nmrylN5EhV0MfaZAng0cS+ttTawEkkJLMsGpLmVtq/
Rfp8Js5yEGLJ/xE6rDiSuUM0ew0oAZ9ZIOQIcWVxrfxN6vN+sElstHkrHPaH/84b
RQ5BwKM7ozv8THHxqTl8xnUWGoko+cvXMDVbk3SOvQquV/flnwQMhpk90EPCURWk
cgoGyGtEH+ejXwxAmODQOQoPzu2JHCpw31aiMSycOAVS/VVypeOorvdaaONzD915
qmXDOgvTwK8k+rrdc4JVcgkv2SduXbwZZycitLktJnWYr47A79KEwuZ69+w0/Kpv
BsoiQiCLhZEqRks7PlwzgqOWXWa6O8aki0st3ghzW1iyMY+xr5YRDBJomS93s6Jh
G0qPYysFZe9MzYADZu+fL2//VBxyaWsgJUXyYSZBHWKtfFvY7UH2QXte+Y0wUByf
FfpO2JEXGWXsq6GrXSno7bTK+JVPtzmuqxyyPO0YjkiDDiYOwQ+uWRpoJjNmLfSN
v7tatlzivOmRBSnEm8zN90LnKxJqHr7DZ5cko47NAXqBtcTJskfPF6HG1K/MnU3E
ysQAr6bMQ10r3U+wiYHuqqOTp1+Tm/26hBZwSiRIFMQ1qcGmfnoRtcQEENjWQUSi
CfOjK1z/MFXQykgKG29aNNkdkNXaHJNdwl1Ikx1SUKlukOdrDk7Bm77SdhTtp40d
dQoKK1Q/DkTDXZkxhef2fdIVuPRrnXLCNd+z6lWzCNQWakyP9oSIX8/XfPvVoGW0
jSk87A9hR29CtR5NLGGXR6yq94mQnDuuGM1Krop88O08cmFX7lZ04fEvqU8Ep+8K
w19bXnd5/h7EPXLsNDHAQqDJSMYUPbp+XyyldIukTkvO/pyt1GjVOrkizJ6eP7xW
OGhUuYntPJ7sr5C8BLL2BTJQliK7Pe63eejK210yyzAMPP+61QXGyQu38zrwaRoF
nwEKWpzSaMg6jZcCZEXY2DieMoKrstt6k545VX2LTF+gtunyulPpsYsMs1VjrrR8
ACtcbC+ddo13rW8jYpMyCilEd8vD+y3VM3PI8En5tKERJeB7DJ/jovaCYGBr6n6b
g+O/atUCmP0UZGQIdW0fLcz28fubpRaqC4yDVsTfMjnjgwTPaMax3TQDkw9tsDbo
IFvuko5yC+AqwZnEK112Zux3bYJvh/ryc5cntsPHMoFhvMm+tlHtdQwEX+guMCXU
wSnk8JihzCy87sHxdhwBeqS5mdznJEHEoqXFQ+/2QcOMz/Ayh5SFVKqoQKMS9y3h
jg8lGOUxHJPB9zeWDKHUBVMOypmHQB1RU7JdNfikZN13/MKgkP7kNEtsOjpJeB6q
P4nHd7J/Pbt/JvavPXmdvHMxB38z2+NkIapD2Pf8ErKL/bmMO/lFZefT1bb7cEfi
iTHS5pCc7HB9Q9Q9HaWk4tBknyj4XIAFwg/6M3cuhxQLWqp/tcyT9yPaEPyQfGZh
h6DZ0huYOtszzuzlSXCbNW8LCK600DJhwcRt6W7ld3TNuEJx1UNrnHMrHX+ZrPKs
ySSEJ+F4PWi/dEqvjJ88s4MuQTxP+6SKRDu+BkEmkbJ5aMEcnax/PrhUcjMHDWKz
P4d2usBVodYksAVy6DGjZRH4x1jaXSYdC3dGoKyy9Shf49vOFvdoIo3eqhlS1trm
RHipsHzftyZ4c/oXRI53xpDk94cgKWBNM99mKCiqUHHZ16u6U5helctuCPCDFKgv
3GZj0jHVpoeG7OTdwicatoNxmpeBnpctzDFjvojIeZUWB/Td/G3ubArH5QCFyHDq
JQEE4MmhW53lC1PB/qrgt9WjOK4CVTUdLP1q1uLkRx5quxjF8WMLbb27P0MWocNg
/pAa3dIOQQFAZirhGU+TLMg5Uxe9dEC8X+BeNyjn5MYBTNQU5bdAuhypW138rN6Q
LiBXF2t9/jSeFS/QBsnrctVd5feZCmll4nlOhJ6jftFtObAbdAWI+v65wkUlhD1F
c2S+8dQhcICWYg/Gtuq692Ik35KpGS69XTH7T1g6cQn4KqIwlgVqN+tuK6aarwo7
dqqyhx3fOglFMTdrGEcMbm31wL3rm/44RppeZ/ngC0McH67g7wL6IKRm8X7exDx6
koPXL874IgWSozNv3RjLPXCo3t1fGYXHnHvynVTp20YZCqpw8WY9yWQ/6UfhWlR/
+S7dWfim/xATS/rRtyDkdQI275t9yHVI9ghZ8rsDuxuEiJP4jI3EHAtLZLnZj38K
0C5phNDPbItDq7oGw9pBgfbI9Gp1jZo+l9J1eqYC/4EukteJO3LEALszPfDRCiPP
8mo2B8BvgeC/MDMSSiQFTL+oKLEXZW1KzdzUeTKd2AZhciNXMIwU+lmmlpHDtFWZ
CbGKmHPZteHuuzbSMNCWwnxPDyPOrVh0rSYvySHgfPuuEw7FvXn2K1316W8PAxUN
itP8u8iO25f2JzJVZ4bZmi63/5xuQ7FVMU5hIa+zivQK2lImgAfDMK7cszwlPhHb
x84D26TDZ8w7P9rMQGmRatDKvrbW6ONR9sdFB561sivdxaPmshbXovAzkuuMgXcS
EgPu5XY47vDSJ9A0CM3ZZ/ZPqm2kNVrdZ0SO+AAPtNV4o7fFhiylKs7rRkrzdLX8
p4O49Y7plbgV+UslPViItq/cwaKoPQ7+8Y81dKN5ILO/TkzlmmCiClOuzbUMpaSP
2szVax7qQ0fA4MyQ6ftP1vJOkbedaUU0ZRHpj6pceNGKZUNcHx2nByLdHZ1bNv31
JttHizyIYbmyO7+9Z7PlDjR8bLVpV2X5s5EsuT13yASadXxvhKGoIIvol+YxNTjJ
HqPBsIpu15O2GVfTUdrocTvBaEGt4JYZXeGnWu31T+p1N3Aonw582zXh6gG0bEnK
kfllAvkBMymT5e2ci36K5YxB210sW1HCXfs8j2j4sMdItBYxbh4SSkZ7mQFyPvKE
wkihp9bKvEeCaDjYQVkzGxhP/WbF4iLd+6IJ8y11Pb5pUmFuqUPj7YW7yUrTlVC5
Wu8DCdH1uVq/aqHQMPGoWAmtg8u7UjtzGlGy5pYK4VdQUbAsxpOq06111+V+hUq8
q+rY3Gp3NVYuGUmzhyW/UTTAngiYC2xH2k8SGq/4qwD9ezkbRVtgeJwcmElGR1lb
OnAow8g5Lquj6HkJSzzgUpwkyt2cZWkl3JoZbVWJm5WHh5QRKJH0CZot62ADeZHP
c4uVTKN2wZEHCffonzWyBi52OR9BQ2XUFqPq5MvOyA/F304z3tX857fxGHLr7EWA
CMpganG7iPNkg8GYaU2XVKmDYeEjpiejQyehCPvb91DMAwKNfvQIOjYX8XXHezxs
Mm9mrGk7bP+oOezaky4HXsLE6KpRFGn5yluBXiXdwLUQ0ALPVC8HibimgtYkxpCp
+d/0XNb5D1v/rFRfnKlz0+TMxUYtHhEhAfT0UWOdShNEb951Lvd3PRifUEfmzzb5
O4XVVD/Umn6Ru3iDa6Kt/yu4Mby7Igog3/h5J/M0uzX74jCJOcteWDuDJBeogyoQ
QGYOxyPoPOrw2mrx17THiylpERqYwTNKD16qZLg0XyICOal8dA/Jzqywb15W9mR7
yeXNoojess1x+fJIk/NKFXrWRgmdCp+PGYuGmztA4BOZAOQ0nrpHzgjmPpSaI/NW
KKhoQrtdjEpO9zqCsmQsXmEFgOP1fvjBh3JAauVgSyYa2o5oeSfz+bDdS/0GvwGv
LcLax0Kun2DSav89DYzqKCdaBg5MhHNXtkOudEweDp+E5Pc2x4slSMJ0IfNchS5z
jPpK2qiit+ThPtN1NXSXGWT3wrWlBBfBN2qZiinSnPVvimXFwVZTP8R+y7sImU+3
4ZZmwVqHnkzDazYJfYvqmLkEXRkxjrloKAa49l7mv0Zg+Eu56McKdOco69DFtsE+
O6LPazPCZ/RW7GdS/nlkjMAVXBN+Oo7pt5GxMi6pRIQDN0ji669IpHCmTOTR5l5b
BdQcNkN9M+/mUXLlGVYZHSkCEpZ889yeMC25YBWfV6QSSCcf9j5TI0gDbnTvA04r
5PrRDaCtFi31HAC8wXzB8GbohLHjGwEjeoS6GaZV0WOl70kbW/gMfvk1XTy6PeIA
e6uvtYt5VwG/FGAIpevsHXBWuqRfEWh2HctEnTF5vTaqf7MrVHHOE2EL/dyCFAb+
bUk8RojfYimyxtP0ZEnhHWPUnLtUl6KUpDmppJh6Qt9MRb7A+tzQWNc2dKkrWLwW
yJ11maOadmKD8Z6lnXmUVBfBuGvD3QuW0Bz41kPEGZwSJCufW3Va8c2pmTvBJpCI
ihrxyT32/PhOgBGVQLe87jtFEwPRY5aNL1mpJvFOdZoHgGoaNgL5FNo0BRe3uH8b
V2SE9cCSBWOwQhK0ybRDuW0aqMmzLbwy8ywqzhSdUKgAdi6aFPyYJ8y+8WcCFjdG
Ch4pq/JEaPW5jRT+9cFIfIO8HPz6lR7cFBulHk9d+yTRwUYU1v3I9QZ0Q7cg63KA
hudlVbqgiu3GYDEg5V8kOUq+g8uIGjeI5ykUjm8UjBOjpXOUgJJud+JqDhoIgDi0
4sA6jF0/6VXSaxE0cUwLRIrI4476zPBUSQ3OVCOKMIyvWIpJxCJvsuLGqO+mWJRQ
zNvXrdkpLLrYeWd2ilwYhYmIc9lO2ZnwZR5mUjN6qPU+gZDVeXSJQdnBadKFICWI
iSCOh0OlCXrPrvIeZ6Wy0BGZEkODF3/gOuO7P9iLw+oeMl30PfxulH8wQ23RK4fg
kbHq0J+rlcWntPIrGByIsTuYwN70/7gURKZJXKqqZvbwDXlMvg5ua1zTHTZ8MSRo
isd8C8ciJaVm0FC/DxJalr2jXUm+efRwt0NIA9i1JKtsTL1E4R2JWnxlZDRgOTTF
eXOt5RFlJaetz2u8WcgvD+6DrFpCYUVbazzKdDf7ORXXSK9mAb9xRkK5+KTADv+t
PvIWX5SxstRtzGE3TR/8MsogiBCxU6AqF7gdNOi4jdYvfrLaNI2WCF5LsDdaOt9m
GT8Z89olvZEmMPHUp8moysyt0xsK2FVTWbKqKfST+O+fK+f+ygudpLA3f8bKzMj4
B3b4Wy9PFClDqKkhGKTGxEuQeOUJhOmjkssUHdmeOcJq6sWdFoAfyOG9KrXTKeCG
XSy3om+NvF84BLOiKtm9Qsh6iHC/c5YOuaBrbOq/FBT4V3ueOkNWwsmZn9EGxxgi
VkzGza3Gwdo2dnI6pyFviASooSAVDVtqNZhHoyXUdmcZeKwbxBLUrtZTh498YA6W
F1cE0+YIgAYvdcUSBGpDCq40QIClaydTJkgeoiX1nppnzjaQxCWszj+w8YBBuObo
IxywbU8FOl86INV0NOlj2FQyPW09aWOjSCKFiPGS2ddLAea/6tX9Ohd7FkO/TCOp
dZHpIco4Sp2HNsv4rUeMR2KfEHmYah89R+HnK2o8FTAKNmj3832g5Uo80bUgfo/O
/+bqdBEoDgdrRDTasDBU+Jak/QnYWdqAIETNihe/FfJOF++rOmg4flLFS408cZ5N
RJa8ZsTs4nAvmBm8W+pSD/nNR9sHM8g9ILl2/qhkuz3RXivxmTuPiWDDWmFNMDeX
ewNtwqqzvmDDdi++5uTekpf2CUmYRiFrikEKf9UisSW1oVuc7W7oLs6sFucch/08
7r9VyApYOCsHJBnoymEQGXKS0DIYtDMectB/MbfJeujBEF0GYqY+cPFkk75QY2lY
sm/O4t6PlMXdnEFSWB5VUe3c1DIgAfsAEEnTgb14A6UjHHEAi51xqH5DRUeUxlBI
ScGQJZFCJ9AruPs2hWE1ZT22WG3vHe5MFEg0QRfAo8pU9NZuUFYIgvO1q/CgDnea
srpD4/ls6LkuMD2KRXwkdFA8Noo/oXbP2Y9/9klkA+Efl3w+Su6QA9nsPumKXEsj
I8/7P53mfdZMYVjnn9dTE7PN8b7+tWFDFI5X0oRDpRqHtFOCBrumpJ+TM6Ek1qNp
HyjgK1QzXk/+AwsyYoY5av6gFmFNCk8aksHrAw9dFmeKbgQduRCUf8mb1nyNmAiE
Wbgi/w+9ix3hemtYsq+qvoPpcXweyjuVnScAFIatpMBf7ZZ8OsqHp1ihEW6QOSDO
wKh6VvPJYTDxJvJxs7n4fiJAMBf3gnvtWEDlVZKu7zdNw1Gj3rmJnHkLYCAVRb4Z
o2g4LQIEjaeWav7HixF+KA7h698K+7eTjUbIqQ8hYwGTAy14YxPyCe2B2+VN6F/p
GGquadTtGWdUsN7B5pwjaEai3MNTPEtuFLj8V7Z9hVP4uiGEK4AHGDrA4MYlCfmK
xUtZEZHm7FqZYilqQ2zcmGCqvWVZWg/r+owHAdkXliCi0oFAOwt8bsqhgoErDM6l
3iy+wEQi5z+nEPHbeGbhXi5HeJxGfsiIYVFQnG5UXYCI/NLBBRir8X1eHmHnZxrg
Z5XyDYvVAUg47hW/xY+gVHxm5kXXDStBlGOytF/T1ZNRkv3mNFco7iFdoRGUgTLZ
cZvFgKGrduJxmWap9DQROhYCo2cmbV9CAac7yen0RvpivrHXKXJAfQAVcgw5pb6H
X6hSbLEXr91p9xzBKUKwDEd0kdx43e1ivUo5Xa2KFGNsywd2mTgeYfbCjTJ/XWdG
zMviAurV/vGETlPgpNQNOMEJbY2v+PLL+MMXcHCazMmoys2EE91JZGUFhbj9Fa3q
wGd5JPoE7GUGOmLKIi1arrYxc32gFT5bwQMoMRBdLXL9/3VLbgL9IN3z8lpK90OM
H9qZGBPMS39A2jigvZUV2Q/XweAVHrLOdifyBseH9MlEg2DCW5QVU8D0fzTTR8nd
P6DDmYtWB1opqKBYfFCgl+aPFTvk4SAMzoqXkyK9a1p1E+LBM8LcjPp3+NdLySH/
CDiU8s2jPpp/sHOtzFYxBsELO8b5QpPgQXHtjY/XTX9vLOIJUpCWR40/aPlzNnhZ
4DE8lJH6wdTD5nTQtJhA6zp4YNOMfxDQ8b8Uda1sLaYlA13xHmwDKM8oFt27BPar
tm5k1Ue7N2GZeNtEWEcZRIpMLqV24G5JibXSlKvOKPSEp+7Na7Ccuws9imbYWsKa
liA5Ec67hxxO//lhrFKAZULuCygqcsCzrUl/uDlLLEFgz1k/BfoH8uHML2zFIoH2
lVWYtNoKFoROwibFuJ5Cfc4Y8CagKJv3X3zpQSKWfw2MVz9AyVFSOHxYYRnh/lGg
8oB2yMrdSSqPfFDQBUplFPw4uOjTfX2JilU044O+uCPqJFXdiN33eyCC8BtnYT2X
3vL/0SiPlhTkIZhdX3ovFHNnL8yxI5Xmbr217aV2YBzxweMEcMRb+D2nFa6o0z/8
PkIXOnBMtDanY7rpbB5kJp9jiyPMaLzAYu4mKKArh/jWpjyUbO6G+VY70c4F1pLI
QHawe/NdabfmEv2ZvE/EFC8RrsSrpLArL83wAts8lLpbYzLVleq3xUz3+LBFsISZ
55Z4hh5fDr75zDhOJIg0n/C7SzPnxrpn0Rg41SA0pWe5UtWAKgVBjezhhcAcwtDF
jNO7hHnJParsDF2DZ4mOAb8IDc/mCj5LfoLSLA7ZL8h7iz2ZCLmi7xRD9y0VRq+b
4nTDMbx6kA1/hYrIlqOFy5sQTUWg24RFwpfOXdAswNbZ52uaqb17x0o5v0BDbOIY
vVmCULyRmAKkdiC27uIwUj7Fyy0dXnbhn4ehIC0k41pzu4ZwnY0aoFKFD4/rUiuX
sezIvgXxp3oivT5BK1c8oCZ3qr1pJIGMjpehF/fIpoOykQhL+txcFtldhed3zcVV
fF59q5vXIfMEW3oQnc5i8b3bVCfjFL2eDgdCdY8NQMZv5YIjcDpWNnwSJfBWqd8L
V+DgBgh+lBQKIBaUc7Iv2ml4IPUACWTyX2muKRTOhVwQfqQJvk+sFRAwX3e8VmHW
IQnNVJgt+a58pm99d/6eoh4rtxaWMhQ/mkpu3rSI52OMENI9/u/AuNpkAy9v62HJ
Ltza6DQKRTHtARUCtK2LzB78Zg7/GVQbgGMMAtzVIS7IjXDpygAquSKRYWJkomv4
9MBjkLc+e5DZDLngOKOuMpdgctTlmfZ7ZSkybfa2gXgGoi8VPNjGm1C14ZzEE+ts
1yrKFjvdpKVBDGMpNKsaXmCRWnUREYh5KrkgLdfUCVD9/BHThMbLG6FXDzYT5q+e
iQOFG+fx0REjSxuuW/VsyXP0/QWIRKMDI0+2489OESGVrivgjFWcDJxyN813eR+1
Ag4Z8ba/3qKPNo98wvIORcgNqZDxDXmy/mSrwSPQCoOelo8/gI8xXxV4adzD5LHw
UBDBMXkowlxaAanXLU5hXLp9/Ii6Tp2muJlyx2ZIbrbrVA1YldphILGNK2vSRuLD
OgmNYwr0P0MylMKISGwTrk2qBJU9pXzOH1afb9czwEYDyFuhEzWTw2LP+btwASGT
LKGF8klr6VJDYrRN4ohfc1Q051dJ5+EkmbKMxT6kGJtFNBROJ0rKPQ/5OWp/qghT
gAME0gXjILvJb/hm8uVvC0aAlnEtNvEyYTR7zO93p6wOen0m+jR0Xyk5chY9vFOL
HrUVv50OFNaiqdjdWKQWJwwfp+Qcv6YFq+T3S/E1TEiRC9g622LheG9pSpFXxG4N
JKN5/E4dhu4rUtRE/dQ/7sXERvtw0LNTU5YUYxONwILxt7iSvgjM/aD3K2vqGwkp
jFXK64Pn3s74S4NBA+7A/DrtFCgYe1Pg1ksvvi6+3pXuxuZJ2BsVDyiV/KPjI2Pa
2H55y6tvh0d7j5XDlbTTbwI7xppnyBFq8drvcOVzXYCHprf6w6FcD0jPPqx39fKM
D4biQipGI9ExOwujQ1S4kYFgReUsAT0nytqsDGx3FfjccUfL9h/Ei8HKktfdeySL
GwWvGgf+BVg64GvH9LFz4CD5e2nj8ZQ8golgqf15Z7RlfBUVzCgog1t7iz8eOjiQ
YoKfemyxhQNkPlxIjwni6obILi6/vApgDLL8c7jJHDqCcybdSYT5y+HEDb2odEO/
cgXlyrJOdNH+6MZu2+kRChKwkeDWZww8cfmbXEqUsUeZ34WMoYC5NwWbVx4kJJtA
kJbU8lqMeqgFbrEntI2gX0S+ufkJYyt/yunpehsmZ3GP+ic+6j17zF+0FWh+GBql
2Oh6HScqA1QzZ0OrvymDzf5q0hgmA24p1GoAL6SuIP8L06ZJ3cv/hmA+ZyMVdWf0
2hiUkuPPo2Xmgiim8Iaos2ZMgNzgD7FoOiu+917VlyzExSaQYSX6ADShw+kBf+8Y
HFDiCtLKm8DtmGhWjyj+4UKGKJ9YpQ1oV1/9Oh1cy3x0+T88VtvmIXUe+onoaVD3
OxLWu9b0eMJaAYbt+8ZtpwLO5Hv45V3XVpKjHHazO4zGeYkeev1I0oRBTcR5AcQB
UO6NooULzdIsUOSKTYd/zzCNxsx4kvBNmlP7PpeHnu+TbHfOZqyUNmVN/zcYVss2
LAN84OmEfcR5qUEgQhhazbalTa1PoI24IGixHvPCzrRY8/T8MDek/BpFDP8CnDDv
vjUQ+lfcd4qrs7qofXWIr0Az0r+brKSyYZhrutMbCUTvpsbPBX9xvrr48rFaWOfe
U9J/+4gGWx7k1qkwLADwcWi9ZhZ1DoJ93sh3CD1HhbbM/sCMBSrdpQix6FBLy/y2
Ruq7faHg151vZIx5i4uIAgnc+OX8Ez/5Yo/quSepFjsl3uChAiybn0uD1Tb+6wJ/
x+Z6B8m/da4V50FzeRwrN7bChYE0EvSqMuE2lUKcMAmJsIOzx2PvjP2428Pdz1do
EQXLWasH26SUyhlylaVgG/pmsWPXht3TDORhT+gNpL0v5w+ckqNnCme24oqRVXhJ
tAIBJRDE1uEx7wNOykbkMmVQfOpd0TA+gP3iJzYQuZ1KuASdNRCp5HVOkA3fi3gS
k4uHFOPnowiqN+yNfIlGVBxQkSOlYV8go9IRGtRQ9BpIIT8gPwjjvN8dHm+j2gct
kJ+/5OSMd5Sql+6BK21yRbEfV7Zd7MdYwukxVWHlpDlXMsDoOnoQnCzZCWN+jfKl
lq3Kdp4J+R+E/P2axWdLwgDprVznZtx3sxrOuJzPVW+onoqNaQYWEBZuiZxdr+dV
STFzUEJZjDDWKYf6RqE3yvIsi+yrF/65I7mJ5uHLZZ42igflezCSK1bZn1rw61uq
67IGSEA6MY8I1lglbOIvWXUj5p0iGhBq48lPdaBIY2hNDfrQqN4odjn4bsrxaJ78
`protect END_PROTECTED
