`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHYcEholwO+1S9Qrr1MQKuBpZwMO5UtdnDaDQ+cx5BdU
mXLgsFUCJrMaUIJQtdMPqRkk2xdMbcF4Y8tsDByvf3aYfJeU+SAPJOASeVqyGhIG
tFrgCK4t3xfbysEAPr3x0vcTIOf0nqIqHJs9FhJFL407LNwtsSBKrbufARV8e+gh
mZApU+my0c9dkkyohiR/tOPU3vb879QMEBzG0lq/uq7rd/x5N/OPgIdUSIFSe7XY
S2OSaZt3g40EAaYoE+3tUHbM/NnZ8CcFoL7UkHmqG7I39rhfYZpIXedz2DLwlM+J
oTFtX3n1CT3A71DHlOFcnEpkFSr5DFUiBHdVulIqZ4/JaFyAO5t+gmRPaOqKVp6D
1X1dxFeffNCNCSAhx9zTNbx3tmMDkpqY8Z/4JUd8D/+lhIwMwQND9aBi4pHPRAoh
OrQgMCreTBCK0wbOlbVlSy4DDE7B6DnmbKuQQsqiKHp/kvPkDjRltqFwAK4HhaSc
xJh1wv13WH+IQJ3fUq40Bfoj5+Y8H+tqmKxXWMadHQ5BSeINkf+KydwbCHAttXi6
Fkhnp+TQEobhYFQcs5jHsj7siwP3+sQSSLg9mq9yQA00VcYm6NWBQj0MM60MICMt
`protect END_PROTECTED
