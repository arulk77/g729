`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49q/xg9aIUKXlWmFIsLq0m8EtllQZQOeWkjc0QMw5L95
SkhFfQp7TqFqaaVDWZ7F7Y2XehjkXCqewbrOZnbHfVck0+H8cIJdz+RduJRUtLac
AZ7Q9/A3NqiKbWTuMDa0GNFotSX+WnjpBWvif69i7PD+Cw5ZKWkn4UkPaRg9aTDI
UCERCx0dkcRtRxj69Y6cK6ho38DckA8gjHOdEI0saNk9w6WgiagbUWOJ+WF1+rXv
kmHMMC8Mj6zpKJ3gdephpZtfrHhwWAf778BwjcSbwKgXxrlci/tC3Be7EHN/oI0F
/ueleJedsDRTA9foENwreA==
`protect END_PROTECTED
