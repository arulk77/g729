`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJoBOVHYdWAobveCncHMe1P+2trwIz2p2YFTSyCXSzXu
5seziyH8PkCsZdlBJUIJ6xSRP7xOI1DJlRTvV5OMC/JYJW03i+rdiiBnpM/x7d8R
2BaAz+YYnNbuy7J0UUg9axZnqQeo/2X36fnHaPemMN4DWs7Rcd5UpC8UFyLWq6lz
cbMAU1Fr8X2Z7tMbVoEq8Vlsf3Cz3mqIfGdIqz+yOKY3A3wWUNtPkDlEsreNG6PQ
brW8KRbv9dtLXY9cq4J/9rIiWcHnVJh2gsM/MzexJW+1trKuIedCj1McZumRzQw0
KqIHqO2qCT9nAoRxRjSzDdVB8IqdAgcsV0cZBokaETOqta0MnM1lSAAIk28cPwcR
9Ro7CPP6bPA8G8NRW7ONfdoOZzZj/Rxd/AKctMtNRbwLjPZa5/HZ6SaHNVF64Q11
gP+yf/bfB8CFa73YIl2QQsggtowfHOHDTiuFk6Y4A889wxstZEeMnHfOKFZExDHN
159Strf6W1ew4Zog+j77uOKLn8aWU4Gs1Y5G6NydvGkXWt5xQWXy9wvl9j2VpUgO
HOOQZtwzE1czEmK+MGQ2YHot0fm54l6ca8D0VQMxzQNEEkhGN8hkiH1Z7L0Er29b
IifSNVVDRpEavX1DKkTV2xdzEKnCQKKAgW7ByeN4SPiui7AjK4r6hYFB05UyiOCj
W1dn8pMrq7mrzVMsm3LozCLD3VHr+XfXo/pQq3gun4sJknxiQs9u30N1UHMDdEBK
yo/1oDcZu3zsVNFIqqTACMHg8/SciDHm/ihiRObv/Lg=
`protect END_PROTECTED
