`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
plzj8p1/s8hNMpg2VQBuFvNVXfsffH0PQyRsvW283FmXQLWANo5yPZfuHWu0u54t
jCZQt5JO9m/rxiZ6+sFVzWB5BfFUBar5exgJcylvyUVbFL9s+w5bVOjeYtXtOS8X
OjKocJZGXz1bgSlnuGeg9tpCi9TdgKbC63yDh80WuUa5vnyJYoxcttKis8V1Ww5z
OzisRAb9ooWpSXi9X06LAYtFHWG21vW9TKR1WewzOCKE1YYqS8yQvWSsuNAlIlb7
wrtzoNVNGGZfhMKbdLBd47JnroXEkaLIrLw59D7jmVTIwAoMe6UyytkBePJYVjVd
OrvvcK6NRcgQQjN/c6nKBRiWF0rVMolGdmK3qrMzdoF95sBt8FfL3pEWGytuMZYw
HohdcakUqoL/YMf0WUgrPZx/+5I0nhIjd8lot4vvmz7WA1ciIU4kZIseScuCcQXq
GjZgjgn0MmTzlT5vuzvSCQ1PmVK9Rf6/9JFoj18/uWQbNZjpnaKW601BHHVx8wqD
54MiGbYrAEe8WGPq2oLNhaSFKjYY+1XOYOriT4HJGLmiSPtKdKV83SHijs+ij9Bx
LBgoJ3a1h3saOjp5sDQWyA==
`protect END_PROTECTED
