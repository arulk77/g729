`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
PA4xonFLH9Yj+OYBPzQ4boFFr+zWRBDjUYCvj84y5f2KhXgKCaof8NMPuJdbWaA1
om65IVdvbBTyfm4VWt8YZHzrBW16yhvR8qOEZdiOKtUtQ00BhmsGFYqGf8QWhNfx
7Ne+u/7K5FnEVDqXqaknVSvQkz56rjCpxMHXoJfwccg=
`protect END_PROTECTED
