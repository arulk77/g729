`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
hNbt9H+/p6u8v8tZYfV2y916gOV9WMU4JZNcwZT0z50ve5UwXBt2qxN74hvIYYvB
TsiP37u7pXAAcBrTfEIqTQ+22gyL2eZ6+/hOH54P6FyfQd+ou+SeGL+NqCZ0967A
UVt2X+nrVGq4u8f20ObAHhrXNxl3ydWq5snZs80FZ1xX64v1J39uRSSYh7EcW8Ak
Q+3wCq83bxC0YFaJ8bL6gI2qDpadlz0LazLs4MgCHgZ9MVnCpYlvCOJ7bh5dBK4I
qY9T3Bq4W8g8OG4HhGdDrhwT7gjZ4XXTEOsTcFGIm9sc73gyH7bL+DyejTjZdMtg
ft4IbIAMOrdnJ3dFMR5X0mI5vASHl6UiCiX9l0TCcQN82moPfI5Tx1zE/9au9Os8
8J/BMsMFdfqism/P93q327Pbbx/ij7inW7saXDYK+DxsWFTgbbxuXP8qpU/vzerW
VGYwGmFl9qx9pQQyMI0aPCeHgXvT9scFUt4fx8Ppju+SMxeoCxz7w1xcI8Ai5UYz
b2erfTiFJLlFhv/+WJbaeg==
`protect END_PROTECTED
