`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOpVHI8C4JCrBObDmQISd0mU+igThUadMSSJrFSm6X3e
DL0dkKoHIE4oA8ayzrlBYtUTFmSo2zX2nAeBGYVxC/cLll7i7JSsB1pos3bWB+TO
N0VFvoaWDlhk/5oRa9yDf88CbvBw7yANzitBzghUru6DC8O+zkQ6FdbSH8LawQLq
+DnHVwp5wGfFbjMy+XrpsZQqHZReTXtWu/tAUFHoYCfeKS5ocvnEnAPLTONx1xqc
yY87J2XK67H9Zii7Gy4gDBAukY0VQFUqcriTp6iWxltjovpssw04luKRCeJh7sKC
tDE+WPDQiSVJm/I63GYJnPdIz0kZgWzAZcw5l2KTOuCvdyOCrMA2yq9Iql2aMUIi
kI2KR6keLlHlRb/tm2KCbw==
`protect END_PROTECTED
