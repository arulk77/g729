`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGlE7zkP/YjWe0AgUqto5mPe92DJQmY3axapbWW59oCr
o0ZnwVyeHEDzI4QEYtsdgg7VltCpKYZfpECbtmK0c5LweGY+wigeOGsn6IULwBPL
iD8/T0192QDbqUtYvPvbpI8bnnvqM+WSDzpCq5JMEI8Jyrx9b+9SVG65ScjY7rYg
+/wFkLPlX7m/ra+oXz4P69b19xS+CpvV3zowbhwYq1SXLd4VscCkX49u816/LFCn
nysPmId1ky+RrUVIE6PaqA==
`protect END_PROTECTED
