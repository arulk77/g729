`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB4ig0C/2gb5sY2NlBQz9PYCMch24Ukhfy9WkVZwjcu2
fBdDb5Xqn28erqu8sM5YZcXo4TRqRIdc7UeEPnSeyU6eZ+JlJ5Ace3xr2CYgsBJN
4Iw8EJ1R2NAc9dO27p2lGCT5XBBKp6fDcyPjmEOXmhqsPzt9ZzgIOwe3xJCz38IJ
ZJ123foIjGqotfuTMyLPBg==
`protect END_PROTECTED
