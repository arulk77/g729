`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
1nDLHe3WoIZJLHvBF3gCK7JaC/i/OU3ltRXNwZHmCh4JcN30qSd7IPmYkzH9DGoc
2+97oCeqifq/LyzCiMsNp2OlF8FUg4SJ2IULuJvSili9gq0RK+HGOmXoYFSl9CTC
`protect END_PROTECTED
