`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aTR4DamgW6Vavh2V/TDykE6uyyNHG1MQrHQgbM8U5CDR
P1SJpWBykEShge8ZGHU2GxODMTWrT6GW5h1EzUcItdNeChx4MbCWf19xu835P6sN
h1c00TLb3I/oNwRxLW1OklP+sBOtwcpV9xgmf5SjTFmBb1kzv2EULIaS5DhExR8r
kBRC2tagUmqmypXCmOGIFRJOOsTVhn32EyrvgW7KM7RhoP1pYByI3oWpzE/Lnh4t
`protect END_PROTECTED
