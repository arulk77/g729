`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDQ8+WgHCayhnWzxlmBhnDudkGXrsbP3OFDh7RHluLE/
noQ0xAcTOioscY0wF/F5b1ICye6X5EQ8vEoDDSgKaw72P3eaIOKS8z92ryV+v7aG
G79+BxaXMVTSDXVqiBl6RDU96Gx6KIz5jzBypk3SfUP1lsdLYH7Z3yV6W+ajzM3U
ZpL0LP13yd9QsPwF+oXPUjUeFCLPHq8tIuWL95b6dKqx4wpwAx+ONtSC1gmH2Pat
`protect END_PROTECTED
