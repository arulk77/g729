`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
RVFbVOyRUulELWMROFe/Fupa/X3yNW3xO6ezZWrL4pRDntpJt0iWfZpv5b3NH6yw
KWzCD3kVR9xfCZqN34Av0pr8KSwATw1HtyhQ23hpFTpkGl3nOyCY/reoOnHpHJCF
yQr/Plq2GT+VhO6LNRDgLyiJ/haoQQaW2+m0yOnoFhgs/mjtoxARJ/Kf+l+FadoC
RvnKl8u8pfRBV1xn/Zl87E0SNZHWIPeaPF8YiYzBOebVi3PUAC6t2fAFl/EBRZB+
DX6+2IQbz9h40nYJG1Uuqa65+1z3LS0XSk0u2FE84LanI8tAl7p2qYifVvPnK49d
MUP+HarD+gdYzWza271fjNAXzPlvqYf5KKdn1ADd9oRvgGWNWnsWWxa3gasYWHUK
5gm3ZgZ6FmkuMhbrdYf08A533Oy2Jy+V9+9VMTsBDbBpD5XDeeNV+Bl8UuWp+Hfu
nDSy2NAUN96LivmZfHw0VM+nff1eFRbXScUSplBlEg7tb49v4+SbS9oFlLMJQ4yb
I75eyn1w1Yv9aVhQ/p6Ob5Vd/bp8puF8203YIZRNBFhckZ4sSN5WOzEOnYJHAziL
IZK8dql8zEXaVou2WZjnk/jF3yyg4RhJ1Ijte645du+UZRGVSfUow1K3dU3ylph2
X8ROrMECUIu1vZ+NCPIKFUqGmBBggVDtLFi4R3vCX6V01EK6sYZeRrMcLw20lD1s
CN/9rLn+Ts0ROSLNvFhE80YzowqGY6b5rU7fgvHZMehdPdSwJEPt4VdXij1AKTNP
/HURgkCMEysPITKMk7BgMQJ8zFw2D+r/yhp+pHiCZC+DkNQeNQGJIFyvY9XxysoP
ZfLVWuBabM/H0a4G0i/jv7h8MVR5rdVlmV9dXFwtJqBaDO2G563Tnlo62wWhXUlw
zXB3WPXtHl0PJ/mu7h1qgKqri+20U+K6jMqBLlKNlnprqI5pKN+GExWLqwsLvLkE
nhZ94M7Hly7YEk7heQSzttV99c+z2mLc+8DC90D7Wn2dzzrp3+bMQG2zRY2EVyR1
PbIk3k04aGBSZzxrt0LeUFuGpBswWaDgvdoPMujZXHsOkI0VFzS6xGtFvdPnG5k9
rbwy1iSVq4K7JFTGqvsH3GVhGdbhXgLqsQCtjAZFjJi5tJie2NQxMy/ZWT8Zm39J
PIadpiO3XbxTQcRqgLxbwPcCckASwDinNISfGjyP9YgUwY6vrGTw/+dPzusizB5f
i9iYwbLLQoxfxJdE8Qxz0xMQuqucvTqjGr3sKME5WCdm6k6rTUp+u5cr8TGxrHg5
l0FL4mr8bUS3XXJReMFrPtjDURfz/UD+fYD+erUpfdLUuIPO6LinuWSa6j3TfujC
DNr/SisMgYDIG3jZSQofUG/5KgQP81CG2Mz3EvlNOyGm5+LuiEO+W4/7cRjcdyvX
EYehV6C99sGhLp9rxEte0mjSTPL3N3MQZkOiW1xiO0bssYhAbJ3EvN7CAsfEWEnw
w1A0ZaX/AxBgAitFAyM0sHUwStMKkO3pauuSvuwbE7mhuzQMxWqpmo5Iangoa2VF
3vEhWOp+k7aLXd2KFLw4WBDhmkWT4xEqzHCPq/Zvtou94gJvbJtY8J7htueNRF+B
7cCUuUn0kJIoS5L3IaW7Rnfg4l4VfwoAGUOQTsDYBMpnfBt6I+h/Zf06dYmB+hJZ
v1evti8T/cPTFeKVOs5HWb5FB7IEjOkg/IrbPmiRcuHm2+f8XfYgcIbGMn46tagw
rqYLmjjC7KlMzi93xyz2CkS7jnJ7N54PJPIFflFf7lyJBW6hiH7j+z7PaPXHKCqe
Fb1f1931JKnijYWtyfuTas7XvjgQb3SDDkNPgyXyVHX9RU/NEpCosRMOwrjp5w47
5cqghaOSY7dmbSHWitr9snZE46U+BwhUwCAOk9MEzrJ6aphdhofXsc93l0fKB88p
EJiujAmBw0WdaZgdHK2kEZAd4JLRC6735RM9xHQsSkPvS0QcRrDsC4n8i5WVCZWR
rH2UaIRbACKawCnRf94liA3QWT3r/P0/nPYcu7ff/iPl86jI7QpL/oAjq9tJm8+M
BPwJD1dc6RL4u3WF/blkozvOGFQSAzDSirFeJSZEAwtpYFGLIr380Yd1eEss6n9b
Y/5li9cmhd1/RW0OHtE40vBLv5eFZx7b9oENmNMVtcgwQ+EdefA7yrW/oq6/m2LU
aw+iSTjIfz1XMiYNR+dzIdpQ3ivg003ZDNeYayQzTmyN0DtMHBt5Nmv2+sQac4ac
z/sY4NmWbwtSFmLMAXgGUBEvn+3fPa0jZQl2EBtPMQ/ojwGJR0oCdow+n5cdjLS4
kFih0VBsCu3Nf0qfF8u9vvv+ZMwypc+8SZ2wRTfONC87e6lZFOEUcO6RSBQNEmA1
f2/8tWBm3WMsxq+IScVnwA/Y4GeoVGecK2AZy6U+e8ckYgTQF+f+8yf0pBzCus/1
P56pl3OS7tlc865HYtlCGFjcQc+t58koHwCIBe9HzatIJos0L/aWjetEQA9T0RU9
N72+a1LrZ7SYtxknhG0fxsPSNMj1Uq0R8hCxir1mMhzLOOGHMcFQdeS2rg1D8aq3
/AifF6EuqDVKU97SiCjfT0US1YqJENCWj/d5EXdaXxvsK3iRuIJAubr1ftNiBp4Z
uKUBuZLyeI0EstCjGe1mZILid69KcpJKZVKvIVN5bqNixcfaKhlFEOvLPckrMMhA
YFHTgdxWaev1eak6B4v38AUCW+7erV+ZSuZP4TbNwrrXOdHlAeHqOMCCxpv9/LkM
Ou5qHMel622pfZcAlVlm6g==
`protect END_PROTECTED
