`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SSGsr7iC/cpExW8Q0OZF0xqoXeP+RzlyB1Dddo9wGaC8
e5WcVemqbIxqwpw90sv5lhYlqPsDpm1CKrhD5JLAFMXMX2/ilyNNNDmEOzEwHgAn
P5/1dI/0rg1B824HE5ORaKlsfphEsuICggyAW14twJ5cMcSLRsgPqcC4au43Flt1
EUCasIXZBLVg0I+MBEJqDHu0Qr3p//zcxzS/Kn226CtkBhVR7syc6mNrqWi0mJ6O
q1N4Wl0P0QozGhT8EfylPHmpF57NZCvtlsHGOzlRCTFtigYgpwjbMQVGBG005b2W
m2eg3zCZ2DfVaOGDklBcJ7UzV/+tUjPj504h7+oHLKxJIn4F1jnvPblrUFZtRUPW
EF+Q6hAdkrk0DW5zhRFE7HCAJeI/3lMfZGdmE1zJDOtZzBm+6E7eboKvwVrSO+8y
CZyHylatBw7s5Da30q/ojkwMOFpyVRgIwNXvU3mowa6nfhkR/sz7RXNEjZNFm95M
N/lzelsPJ4a3IxK7UAzJjekZ0Zpz8ntrf8WfV28tiMNasZpD9xXN4X9gg3ZGW32U
Sc1LgW5LfEi+f+bdjhntJEXwHBDUXU/ocDoIg0JREYcAsQrCX0sJyCMWwEPBfkUh
/xM/8FBPRW+cCLfYM6xVwHJNrGlNDwEDYvMIV6k8lLOjZXTIw5rxweOnjQq/Ggkx
LJpEpibtCE/f2OWKJHgKO8wXK4zuRx2/ptqOUGPJGAzNaM4TLMd5v0VD/ZOyq4vg
N+hsxY7ojMlf5a//f3IfZxLqfrt//IERfT8Gb4rbKJZYQJuqUL8KF0nuXSLCfqi2
Pa+SL1X08sQNSYWb4K1dWSKrsNPR1hPeXV4mDajchRXxXN6VvBp30uJO4ZWQZcVx
36H3vtK3CKEViHdqZQyvW+i+ps7tBmERxxvmMo3TvrgLFw7n3vc2kKXms5vBAAJ7
Vnrcjf88ydCgrGeLf32ahoitAovGLtG8wJTDuzqwAs7BckoAG9ea/Rk1kXEYLZdK
DbPEQvEyeeMts4kg6HEEjGTqB2XYsQ+xIVjWtPdwSgKrVGC6nVPyDc20xew74h2N
TGCaG7Z9q8mZVr/ulKyCg9nVCl03D88KjCCXVYE8thnBOAsd3RwdsUfUKeDS9NSx
NPk7NVSwT9Q2qMiQ1PCgkl1dOr9ZnEzPahhaWonPGCwH/qnj5G1kGvkAxRfllWaH
s7f9ukkWL6gnoqyP10MrmoEGYTj081XsVRMrZU/oBNLgiZnIAtvXYHW+S8SbySJU
JVKbsV6xDKYZkTwnmYdiGx3tb8psyn+7zDYV+7uCAcey0OYcKls3vOpugxZrIzFH
k1Rev8qcbgeOUFxqRlJ5AeSaGJrzCyy4+Ryad4TnR/jdFhRgrQIcTq4NYrs1swN6
Z9k7W4fNFRk6TCDeJbqqAWJ583PR3nrvuWfVm2I8r/I7R/qyVkK3IyyOb24GZyo+
OSbFuQirjvH/Borffh/1UE7yMBYsGRgfSKrDtx6acHAmPz2psrjOy7birjS5+JW3
pfLeDKmsKdCQTyMQ5MXo6Bz4Qpa3koNGvh/qMlcL8A2rzEfqzlr4neLecUV8iJ9t
YVIjH5iPylJw316tf0LM+wUsJuchQgVgIt+SF0hQ00Nf98ljQB9L2fCK1FbxMfV2
SCzSXFTCrYs7RGRHI3BaBjtY2/f0ozxsrhzyYFnnJfoBwR9qd7vJSQiIKxJcQENb
GWw1VS0iJ/+DK7JIyF3BWyUMxD76XZ0vVZ+sVhlA5Fy3uyq+wkGWOHYI/FJ30p7Z
eWRc5tV8wFtMcKavH3bux+2lxg8V8MmV4qYzA+iaEXH1nT3FOhrgXBXXPVoXc+4H
U1kRSrrtVtZWBUBQ6UesAnEf/J8vzWrRsA4dGAXNhfLAE9eQI5J1icajJdLoiXXa
cbiMUJZ48pv9uEDm9Y+3RcNXPhenKw60AjewOVwd2RPS/9h3qPtMYm9LJvJL/uiA
9fcVJXZ/on/PVIdRNWR1b5+4l8psSy6bKEfM2g0pvJGf8VYz9gvTvabUtdvK+CYK
nc5xJYphuYqYT+2jFvZyNCUAIi+pQ/ujxkHXGmnPpkfgTU+eusp4A1TWotJyc2Qw
IgQPqRdKUIUJkeMgHtvvt6I6GJVVmWmG+WRSmHwY8mRy0QhhV/HYdMaUU3dIs+iE
68aoyQO6wibmujfI97Z2dwNpTreS1+qUlyIfrw/rCQWYPcoZZjD5SWM953zEAZ46
9SA3HabOU+dw26M7u4r5FIv4um+RVwhArDF5/fN8oddt4xp1Ssi1qLB2wfjFBTuf
0/WtPu9f/g4QWLyNMkgkJjUIxCU8rStZQbTniGJMk7v25AZR/D4wP5Qx9htg/sfp
hKMMlt6tD9l2zuHLweEN/Evs7EeKqzICqqhAiNNM0jgDy1asQ/kgOhNptVN3TQh/
ZaI0hct2wAqQJX4oaP65H6hdT3HhKoqSwpMMrgju+xPvd8S97lbPwM2y+ub1jaXw
9c6QUqatc/zbNEADcYesItYlHhE+tpU1+Guag99wlxQjoUEQ0+rFSIqT7foDBHZa
9Y5XoaH5v2LoIG17pOW8e7KP4aTowBt3D4Lwn3XwJqPUPa5xEJPM7YPEBdgiYi8L
S8TSI5k3ZJ+29LTk0XLqxeFSInpBRo7IzTSseKN/jL9tLcf7QXWW0CS1WE+TbUue
utGCQo3hJjLNydJAXdRb42hNBMn7wdlq+/mWNygMjiW72ioM1Uf24rLbEQ48sPrx
f/f8zplvGjSscpfgXzb+XbXoerDD8iA/aAiNGWDC10xE/1A9+kkNbefbVvymLtbd
P1v30LrpwwrurkO4x+caqcOaEx2841pYoAXpVVKURVZn9T0Jbcx7ARigC3Q2Hm+J
8QaEaYBF+oBhVNeg9wm7kEoxUWVqXNNtR2T6xHGZk5Qz/+pGAnBmAVAATiMeHYcJ
nCtCtQh13vkOeLh5Fb5ivQVVlFGNe4a3BSs9LacNrMuJ3dr8x7jYdAM6rG5q4ALl
UVvohPk2kNWRchEIjbikesHU0jrWGJLF/rVyRjjPbbXv2ImHYr8Vjge43sdj0SFq
v66LH3B7IlzdLXL2ZZeEKhwuoKfVEarxB2P3skXAm+xLns5M8u934tVZBJcVl2Kc
hGr65h6jDbUkFzn/5N54FgkYWNAXxpn995VB9fk8Q451i53EUmtDmraOPlbB7Qgb
UDxoIYuFsHOVrgAZ5jEvYHtj+q1wsmPWaU4kaLyP6bbOpQwgQfkegrYTIAPAGXpt
iLQGUhaghKJP2mbX5dsLXlaeFtHwm16jPrMXAqmZRN7Uk1ZpjS5wsj/oQhVkOw2z
0hbI93l/WjMkCaQ1F+cfzhndJ0fkZ54SDjUlsj+Hof7tB19+9FrLV/J8PJJ8I3Zh
fQv0diRwchUg0PC1q+N5BUttiWqUNKBtxuPinX4RYrG0HWJAsmVxIM/Tq5ezsTm2
jsG5vAlWTNldamuqfpKrR8R3NmZrJg9xGILBPiLmB42dAxky1vo2iaqssdVL3oU1
gY/TTI7bekTW/ty46KO59CmUuPUfmDdS7EpWv93e3Eq4SmdXVU+zet2Cq/JGIYAM
efDW3DNwQKTMrWPv1dPlsi4DHvHvXrC+FUB2kI1IUZKp+SleVJcRREWI1uIS4q4O
CKsxMHNIoFCpvDNnrD9ShYLAQo2nLTcL1oJ6yO1XysVK+jWZIaTmfWqPg9jJQF90
iEzD7mdFWtBTR1syFsun3y9T/7zMAfPgHPO95cfR71nBETqlFTbY6CAvA0yfDbfj
XviV0PSpxlbd9iNKNHQy5OvKIdJKL+yH7b7GvAYRHwoL0d85xHkfAt3hTpmE5Ekk
ZQM1lCE55dYf+iL/j/XpA/6+s7oEDxM2EzE77mNPEtJCRq5C8BKONwk3FEScpvtW
Nxg7Zn7rJo3Q7uZc7gZ8mmFe3sSSsObMHoeR1CQzW1AuHQAurvNFU4bzKbt1lCG7
Ait/AX1dve5UfIvTuEjenq2Ag7jm/Ib36cV+XRItoNhebsB2vdEfsESUYUBsCWoD
nWNBfhBZZ2ckFaf7cncQQW5idAd096vCdcXHL92DYmNHFshNLa4B1F9bT/48GcoK
zJBmtvM0q8x3anHrKnCEuFx8zzvBJs0z0s7i5DA/LWO6LKpZWTwAkQ0af6s60FKs
mwUnmXihMQz/sPjUEi3AAYepqQeWzkFmU6rB0PNpF9fQWXeirAomJqsBcOvd2wcv
7DcMI4wWw7Ez0E+reTMGwfOb33WLcoD1e3WFZ5Mp9Py5JrINSeVMyyRHYK2K12xo
wwiNOnGvXE7S2E0pE0pTaWRlYqZRr17xyOkTCJ6jN26fhfvIZaIG0C7Hu+qbKM4y
ZRaVRoTQOZZoxRyMxxQEPsGYwgcLfWXCGM7l2BBWi70BkCNxClFBYqhhm+8pjS+Q
QmqRZUMOVvloFBaOdYCSaIQxH3k6NMYnykniW0WPFhqXF2EkeVOvtPm1rn4Cywdr
0DgIs4mHKzeIgIi7uSM4xax0Rtj35YgY+VBuTYi5X+21u3MejZ7P8E8iEJSF6mOW
JxyWi3BQ6NTnROT17dHgzppay4FQYmMy3zhMmccXoPoOKPa/AVxM2htmRQFFjCIn
dH14sGQDUPKF+j6Xs7TmMJYeX52zWSoTcCYdFnegCvtRWVFXqGrsuGtNEylv1zOI
GiaQ6vp2i4tQEp/aGY4ng9ZQtp/TLdiZ3EFKx8AefgGr5b2jaxV/YUWhsDY83KN5
bSDzP1jfmGE9W7S8v5jLKQAxvjKjxzwqdEwKEqz2wLQv1dScgVvSpD9nvlmggRNL
ex6PjO9A6cZqlTi4hNPYfqVArGUhoH6F0EyjzOIw2wKjTSYTCRQwX0UG7IC9krCU
WtwchQAXpPJyOMzvw8RB5BzneKN3Og6f3eUPA/CrXwASyInzU47RdU3roXk70H/k
b+YohKA8zIUgRWm5clZ7hg9k/953e1TmQs3fXEBd0sO85zQT0aHxDV6cjHWJ+2yp
JC44k9bIZp1b3tkUTzJJUfMeq/wzdjGFnyhKy9C/m925CEAA+gwtyTz7k8YClJ8v
uthisbJpb1qAArZoOqOpdeCDlEuSVYVhtJW6EA45aQZmDWszulHiJmaazX8YoEIc
MboOJUNO1kW/gf/FBxJb1ZXzlG49NA//LSSHn3c/cSpoI3dvlCYU+X+pFOhQSd2G
k+NDPdPVt79b5MfaYbO7/w2owVgNRiZ8u33KUb1tj/IvH/qhQiHcJC5x87/+vlU8
OxPb7MExGlKJuDA7urSWP+Yg11T7/4yZRuuftG2d/RtRqqEcuH94ENYVjN9qQjZn
VUaaQV4wD5SyHQ/S3EbP2W6CqNxnoq7R4ieKujdke5cMz8NtGGr/t9qsvsqdShTQ
lfMT1dJY0SzKEmIt30TFEdbukJeBO8V3XfhFRlxxgUXRjHLrysAf90bUskIZW8CA
7tNwghplxjwIT6Ypm7sYfrDS0GPV9rqvTVo+TNTAqZU06RwGihcrxym2v6IW0hWA
s+8nIqlOnucmi/b+9d86aUtQlAdM+jktUeR9TlyyOM4T75LUPjq9lTYPDgvTulVO
4O/4rEPuq5Uu/Bsj50yZqbqab7bcs5Lp3TOvNoRW0Wy2uY4UKXlDSeQcOE0GXRPr
KqYEWZymq7FqQm8zx4E25WiK3YrZZRizGzN7RX8t0M57Ika9IIHqyTTzZJvKjKMM
DhLQaIusZ8BEygLh7ZbcB9es7O4th+IUjP0PCJdeLSQ=
`protect END_PROTECTED
