`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pECbeUSxU8Blb91yjszL1EptaHB7St5ji0Q9+wTVCAUorPz5B8cJzHpbWNL6EL0l
cYv3clNGpfgyi8nODD32HvYPhrwxiLPhH+ywqYJEGR7PbERH/y97SPRXUkmdKmvz
WvXwYxpuGNjrHHVaN9yzYZMeLQzsz54endg8t2YcwJ8AmU0Be957JRttTn+f3dqp
26LTH2NqEj38KcoOhW5WSWA8xKL/cwfRtwwUJvX51sxkORV6aIXsNSobjPJqyMfw
jD07OWnnKCdwtwSlC6vQX4qIF83/tH9hHclyDwXYQ7qesvQC8nsMhIK4DX1RZfTx
0LZQGxUWwXcdNenME6YaozAAI3aEhXYHIKlhBOP2/KdG2++MWz2VDrRPTtAKoDEZ
leLiiy4alxo7dL8ylS73s920W9wJ/Pey0fdaf92tsr/YnKEvLDHruJmzSlSiOPZX
2XcRCMn7gQqiIA3ueOjRBzYNqqlxq/Wiu+mw7gcjpTcDc93akeY+EA7CuzEXujJH
Wkhg8jchcDIbFW5yqdzQKb+FtDZVr1gRBYE3J3OIkUO7ezho3WmSQqh1ZrS0KD8T
bP/4Vc9K72G1V/IVpEFsNoTF2z6pkPjrlgV09uzRUNDN+KbOKkERayOKG0HlMbPy
qW4xZ9oe0kfh4jvmuXLdMIALLmdHDlWtGqUFmsSI3PVKTf2U2HZxv/HX8lWctXo8
3hiEbppvPpo+uSzO35Mm/F0wUx8Xuy7f/O4VhOZsyxj8PR1mrjSHAeK83z1zA79C
7M6fFhEgk57yIAaFmaMWpeuYGpxGuOcBQS/T4jnX910d/yPOIxYWb159EoMw4iLn
O95H/Io+KROylSVQsE1NVrA3x0NwBRgFyu5854748DTFm6RYF2NvWRtKqEt3UVLo
yPYVUCzw4ihpQVREfwuDL+QYpXnMlB7QLmVgk7wwoDq0Kqci4qkHbiY4stylmozw
AE9RwiD+PgW7ROsrOaxkqawJvWhRFA8HSyqye5ujN9mnOgV4gUU5PbR2eaiZrLoi
Q2sdnjjvNEClB/2UVRVvDUFyj18oKygJM7imKZ73toCAfGjAsvyJZ5YOmsw+wAO0
1dxgT6cRmgP5mYrTxgXlzT/cqDr6gP1167B1WRf26jTZj3Oub19R1bPwnqqLyu3G
7xs4azbiytxgwAqLOQ8SOU/L9R3CszUerKXakQ/2Ipn2DvLoJ+pKabnSsKFEU8Z5
fG/w6hzDqs7XitKl1CMgOWugzHV5AIordEOm3LeARZIeaMOAL7XX0S82wguucvqw
ZqmeECIWqd0mXn0mSBkaNhqYfZrU2YEQT9p9LKBNIlKpnTXLmkn0hGFx2zzkk0L1
x4IYVrTm1OoF4UyUIKJNnHGaWMay4k9k8dDGNrqc/oTn+m7cl0IuHlIgMeN1mo/G
ZOnsb2z8lXcmnVytBpkQ+Jxeb6kdJdcpynRMtY36/XKxdn0D6bPi1fKzFOftk0sR
1lb8snrvpkBr7ZoURgELgh99ZBvMUQz7H/29pGCRfQ45VNAnk6wN2Rtz2jtMgQ0T
Wzln+4DEcGyccbt6PhfJDl49KdrxEsBNZSsThCTgjVfHoCxPxHjS0LpssxEjtgOj
pthY9mMw6PaVYVtdjyKThe4bwpxcIbyMNJpkrGbcVT65W9DknavXu6YFYv5GpZ0x
olWvO32ecofL22gBViQlOQsP7x4GhK05/vy5MhmtFjjeWPoQfLUA18SZBy6esoKg
XzZiEXmyWNNifFWGqxpTHz4xIBTqBRz2PGjRjwFx0N5/w932kWre+Vi2+kdcp1mP
hHYP7wrh8tJVnEA/vw1te0iYr/ny54KOcL6Y4SwHB5tY4lr1fV2Y85qiwTMVLQF5
Yd568bQqp8GQakHBWY2uR8hKCr1J0qw3hyajxT9trCkLFbMcds+mc7jlOHSydb7t
LUt4Hflh3K0IRmJxevTOUlDEjWaA63xtfNeRcFXryhfQ5U3/rrU/LnoDfFdrGzd5
d5D2IBZgcNAc4h+zTGMw59NQPFWhDJ4xiYsKmHHX+GiQ2B8wDz+UnGSR825SLnqD
/zSw/d/MCLXiYqHmsD3n3ICKsSV1sqnB4WgeqRAi+V8AeKEHifXDSE2qX8Sioe6B
JMOyt1dUoZuW2m7DJjGhVrhngS/Z+G5wgEzm8aPvnfrB6ZTmLUxrVmWBSluhvlWA
6cqD6tgx5xTe9Ke0ldDkuKSFry/AJ+3YRH7Vum7pfQ0JiZi44xH6q7yvA+BgPNjh
TDEWR9ACvYgkLXCmAgOZRIrUtPBT8S84rKcDmC9pPrPewYONitJInt2vMWinAuIi
Vh+T+boSbcjLzIfrcvy8aXGADcRtPn7qCE6uGQvu+FYnyJredLLawNo+kXEmgk2r
cpDGYPb9m33r6C4BCEeDXWyVsmxBKj9/VfGDDuMULm/xy9m6CiOlcoOkU1xG/pPP
yhMnoqtR8kNOdOK7so77XPJADAqhm1vrfFtRl+KP2Pv33XH4/fTkZe4ASyTRvyHQ
OfAu+04NpCv1oy0Y7LAByckTzvtqBK0s0WmVKEcR44GDtv98qDPOLE2oJh7qjMHe
OUhoUoyYtyPUrtX5oXSv2Dfr9QAVZP3fa7AhMqzNwxR88CNuzuPELxmJwUVEMydH
mOEQ6fACfEOWoOfceRSGRRKkKyz0OsFzTdah+ZBoK/+eEORc2ePqBQ9QCqpBjcML
9HxTPtyPSJJSNPQ3I+jjnhjD2gQ/GcghnUYtCCw3rwTmdMJN+cgzySsE/DyX9SZj
3kOPIMdPpZOT/WyWtbt6ru824AknkUGvL6aypQu5maSp8+AFV1JItPzg6McFDia9
y3tJLyDVomfkqe77nqTso0IB4FPRRwqdWfaKfX4jRiKnjBJbMPDtnUKD3Ya0mHTD
gBi9xDD+0M9/+xfIFADQlxQjGeN6u/GYJvFlkbdg502vqVaYrC+Gz1PsX63MYPjL
CLXJDSJ/lCuJV6a//OyND40zC4d6p6MzcpnkLKguR7+iMyfiSUGUpYf1XqgHAKyw
tKxs7106I7DreIHCiGzN2OGF/h1XQjxXb7tgd//fTFk7Wtwon2NF1Rj7Yfls9hiZ
pLoSwTo6R3c3Eif/9henzm5uSkyCcME5ItuuT7hlYLN5R/+ScaPgoTPr+zap/b7o
kyuVeN5nc/G4cWE6QgKH7tKye3lUB9B5LaIG8w1Z3DfLx54muEGMbJ4EOibfCcT/
Pbzpbw0nQ7rKVSk0OBje68JppDkYehDDJveR94qzg23n7F+UT7WNLSZhO+FlkIde
QU2FSoLBVh83HwTdCVL+3ApD4os4+wemiKuQMYIa93141XGjmJCP5wm1XU/UqVjt
XXqGcr2bB3eM/WyXN9ANCN6lBNmxAuMCHbsNaqkACDaUBbNUubYQw4Hg7KHuZ1FX
sHL013axNOZFN6WnTBYsZunYPsSi7dbhOYkHziVv6KjI9Bxg0z8gRNS1awEAF1Qi
LJ9CmPCBx/bdftqnqSHm/ik32AKl/tb+kqdsjEdiHlvRMliPhZ1qknZLYuv6nVKe
39hlezlmHnHLsMpKeejoJI/5gHEbHzM0ALK6m/eZFhLFK/rU2xZY0F/V6DbRtK9H
lpfR1w7ZZ15VkSV9ZlN5ut1psdgmr0Jzg6UCeQnPcbH6lMSOnq6pSo+fjDZVpmt6
toTBH7AqVmkdVkUjvfulPuzD2K8SG6zkKHuAZ+oASAGbTkqgF06QQwzfTP5sUUQ1
4LDim0JXyW6+d+cAZpAo1bB2+v5vtCOJ/JsN5Jg8lnyU0f1GPogDcdo5BInSFPjZ
Qm5Fi1RvZd2e8+S6r5P43poZkzVIyOHN7asgimoOm7A0VTHjqO+ZGMk37Wni1bmd
D6h6SmR/lW60SSi4INr7y5sxDZXlQyV8mC6jOKUvLMFQydKcycrCvVEB/jLhl+ry
7NX2X8t8+TrpAlUDCqwttASg1B/1P0QIP5Ic4bT0Y9svY0fCFR1VlnMXbWBtAlF3
JPT8Tne6xZiu86ZIAOFYGdD4vEAQ+dmf4dTwfT17nQx0mM/9UoJuClGIpQx/nI4V
TvNrj8UTtKy5x4FnvlMM4YhEQNgpYS7QkInIHz9KhdamO6JniNnKkBIur0nBnWM4
muAseV/TABjgeXwv0vMyCzSKmET7iTQd5gDHdWwz5daEgbG1WmcyNzyl43UfVL/z
7lIdJCZtrv6auTdWlhP8ep8JSS1QzBMh5hZYxjavLBiRJ5Redx54qxpuS7jx3jhL
dfMnQPYf+RxwWYQ4vsOPKucdQ+Zl3NSGltDfK0x9r93RaG84B1eDMhqqLw9YwYcL
DNyNITUNhR4OaiJh5SHLkqZ6I/10A0XxnwAFtSAClRjtblOhFwyOBuFulPhbcY33
Ag6T7ZlhSxk7+mYblJoxdOrwLT6uepDEOO80u8bXGb2FCNBUz6PVwtbqe/WUJHro
yNr+V+sztLku4Wk/ev9S6FnH9OHfITLDOkGSP8s4XEdlquiGVBBRk0uC1zEk7MJR
+lTBKrAx65l/cYMmg9CgdWrW4sYvbTjSvBiZZjZPs5xrujgZ0cPUeQ26waWmeImp
KuVpXNC6qMnoWm9J5Y6meETS71NECIjaa2MqFiS5M60/hXepPPggsf/tGP+TrGdk
YQNlEOXmvrahCubkH5z9baHGGT1VfA78+WGnbJLjU+49m7CHrP9K85z2JZRjvUfp
2QJuW/rw/fZiTkKorJF92k2u5AofQUD4aeTCY+WvBZ1drZqnOq0YorIji1+sHsPT
7WatU+8fJ7GDTUjEZlYiipYOfMOdwCRTTnu5UQvhEPeRGlrXPbpHZ4n3tGFrwais
bePtrP7/wMOG0dIpgzihO6gttYLVGzDi4/nlP2oqaHblXTsy/K1FhZtPMEZ+i8Ht
ytQ/Zm9zCg61EPSlMAEf+0BPnyqHTZlhjUkaLbmGNPrEgN+Q1aPdve2glRcDUmmQ
gPHEt68/HFes3xBV8qiccobaNFVM71Wv7RQXpLEv7ZGNwigDiXDQw0ykjJ3r2Qp7
zZKdYM+SHCvIsPxCa++WUkSkKRL16ZLeTspGdM/+VeAI4v67hCyo5AXoai4ybDtf
+6r8HWvKfMb/qKIy6yOpxsiXX1BD/3aGc+7odXG2s7J8OLQRe0YSyb2Ib43zqNCz
unpsw0StiOVBNJksfCVRqBvWEdcCYEgnR6E0ICFS0nMfT4hEGVmy5facEDAhKcpr
r8Vbj8m7bV+Sf+Cr1qf0QAbObRQfTEq5IC7fnvYSIuP/m7RJ/fP70sbIgMjAU/fZ
gHA93J8jQvG1B0zViBACGoHDxmEmC8r6wSZux7V/WXFgbC70AOWcN6EuiMpu8ZYk
oeGS+MXm5rDm02b5RTp8zsIftSsMRCD7F0e7dC94UXnbua4M9BQRMB+3s8pfYo+g
M3gq4Ds/09dThfZ7YIf4JY4La+wqMGCjbJxkULubq8/DA93iHoRe9SIGY1VGX81F
WRPKLUtTTQi16CxEi5CUhk9EONKl2JJAcEfzAnEyhY6q8a9dchYSxxRQG0x/Y4Ic
8b9n0dxMkvtRB1gZuPdwUHID8ojnlIN+7O+QKgllvV28kxkYbWnbSN5eN0kfgQ2t
xGfPuU7/0k4JP2vJ66DlRgF1HM4phv4Z1Gv9Ht7Xq+XzICtrC6V1wKPkSZFx+fDb
vxPzF9VwBya0bXDPYldsnkuBSc45+wlHMMNhz4XTzjlgiZKy6RHM0hNFbS2vkGtK
N2WGoLgnbiAkmiL5oU0NwYg7BaH5tq+9vr0lvPq2NsbDZDysQWvL1gz8shl/8Kaf
/AqMWVZf5uD0vZIJMnfsIzjSld1lwhWk1jarvr84I/D3uwqzaVl5eZTva6Ublpyf
PHsCrchG47pl461oS7kpXh3633IA1kZAftaWjza14aTTS4znGMjrAurQb8VDGf5/
syigEingNmH/MCVFK46FcCtUSsJIsmRmVy6DmFAUhoFhAW9dQG3vMvewVcZZWgcv
I0SfMpaj6uKHHotwCDjn9qHAx9IRKDwKZ0tVejmcPeJ+m//AFcGGwHIHPWRP/W62
JIjsls/Sfi7UtrmItd04mEAi4hPtmOk68Dpq8xvwYgrmXGeNTHp6evrr00HCvXlJ
6OLD7BUsWfWO1zr0ad93lVWymqPJrlBCQ+3s6jYzadCIcQYSy40jqAISB69xQ+v5
zkxQKIv9OCm1CfCwkUyl2CuhDcYzATH48UrTqDfO9/LL7+cpB/K/9whtBLAsVQsK
fzUQAq9R+E57/MXOdNhBRL1hwVbfoPs0aQzVdJwCQ8bK3s0gTpt34gVgDyMCVoBg
bwqM5R8Z2m3TfiNoWmaeOM3anCzo11P1O92zejy/ghS8s40zImUQcVfr83FOtsGN
i6XEYPvunnd98aA/u6z0HZCQw1dELn9aHA7g7hk+oNPTpEkUooymMJCKK0/24dhJ
Lux2FKk4sUWMJq/jXAA946FxrDpPdgH3i9QQYNQRWl7OQh07Hy0Yfqt4YPTlbPGH
A1CAvafj+7gOWRcBDO7pGZ6IhUZAgeEA+ak/T9DVMXxRJSReqfa4rAOiy7n0mwNq
uKcF896Qg4370i1YGvCVVyIIF+sW03tgAbVhAsD/PsTN9AgDH85nYBM7X1KCy6Nb
zOjoeMJtwKlR2AX9f8VzgVGBgwO/KRYU3gU7LHqyGKnytKoD7xzn5SGEBJCkIss4
VAy1Bmk2rA4pRrCNczAw22BW+M5Ro/mbolCXMhV6/lkaBRqh22Sm1njgQ7+hExzs
vRkiYeCx227xVc8VPDzfaVHkpprnPh/M5qaIWe9cASzEW+LJM2zxVewEMtvLiOgk
IF5tSPk/ptLcUchJ/o3OW9ZK5huIqZUld6uNf5xFJ1amwZ3uiV+v9Tm1dF8ezQE1
N1aWugVNnP9dGhEJw/+ZDuMW9e30cZkmW0ywQ8nTt6gB8HC8Azd0YCQSl9Nx7h2m
F9lWdqOKW7Weva78fv9kk/4Rxb5dvAs0dSvrJiTJ68RxNjBy8DU0fxX/ebHNl9w3
JcXvYU9JjpvTPzNs2v/H2FB4CyJ5mIDSmqtXCfRKA+vLQUKgq+wzUDtHspcul5gl
9bvY1M8YLdXJQdzPlpCtwxTjF62yqd4y+9m6RSAS2zcrB/nQjNkyZlu4Xk5egZGC
j8KrAoFvxgrx4iLeU9W5WQLvqsO1ODoKpdtQSZsYvWAdYEmW3AZec1VWFPGJTVdA
Sd0RUiVP8tk0hqDE5QVZHERrBmuE3RexA2uZoaY4NLbdXsD5LUAHlK8F0kNs2sie
yM0HgGSdlgm12hI58KkxBsWqz9jPR5kPNLTP++doz80dGoqDkBiww3ReeIYUZe+t
VmBCin011yBE/F+pF18kWJ223QjmQeWeitXR9qNwSnl1zJtSVEJciUbIiT/A6dMO
FsEUrXsFmn963aoBD4WG1vWNsKdNZ0lDSF4i4Bq6VUABLMmvrJqY9eUXEjkBzjxf
gBw5GO76gd19WNHVGkEwz6FxArstDdy4e0L1RdBHoY/xPmvE4mhzINaCHUU+9ZvM
kDT6OB5CasQE3+ouJJ5eEGOKchxTLKzRSj3CEp9SF3dgK1nxazCvMSRwFNpAG3pU
qqgXwpCqsMhYOhbvfCzUGV1iugkMU5ngCW/LMenIzAW2+o48pLEkDsikTATVlTzN
fT/L441L1WepfHIjxa0Ds+iby5zkW7hCDyX5AyNi294NSr1uBZfhHHAY1i4giaOW
sPXq2m13wojssCrR5G/wljUKCOT8LKOt5eX1tL51tE09uTb5nM/b56qXTghouteV
zvCmuTOUJzEtiPxoSFO/OQHPQ+jMdDtQX6DBpSoTbPY6VrStDlYAKvmF+eTgeiNB
iKepvkihsIuV/blzGXBC07KOguWdbPtZyqn5V7hn/1km15SyaYz6h9ZMrqz7OZ55
YSluiktkgHkwxfcYoyn0+h9bEelyHbPlckhJl6eKpnNkkhewU2gyLCPJWT5D4Z6u
Ff/JLZCppysfbfMxMwoLZLpKEqu9nkBs9ZmQzrz87g5Xj96gd1dudjjFMtVTvWkC
djhxKBvhNiprJGJqqLE8l+0DO/9LPxMbV8z5qYrkNUW+JPue1WY/cTGpRyjVk9F2
QQTTQwvXR2CfSPM5XKBO4Zi2VG/km5Qp109WYTWj4nY50gOU3rsTGkR1dQpHpGLS
ZvDfJm4AfsH0AD9H8ZkNQeuXHx81SLO/45SXeF6a/giFHtnKczoA5M3UnZcbsHJ4
BkMUfziYX2qkn2grl/dycXJey6a2ZY0WlUGRsRqRsmrvqF2zO1vcxCrb0MAfCmeA
YaAdtIak/ddM47dtgOLq1aGSTIHuwy4voXDG1eJaprt93DRNICd1LPDF4xnfUaD7
/bMmAYvTGYxTijvrOwft4hvuALGLbeAufr1VWxede+pelQCsin5Ade2+YpOP1q6g
JsoAluq3xi8m9bNb813djgktkLIRmbjFCVOiw1Yy6S7SwEQr5AvN7t8mK7oAqCNK
v5l2Tg486MK5yXtxWqbuuyDcdgjia6a2U+1o9tRYoTHrP+XOpKZQIB/g1Ab/YZ4A
Xz+pImmV0mBDA8PDVqX41PoXSu1TBb3tOnzUm0F5ZJHkZyetCP8/mY/B8qe+FQLB
pFrjfVz7mrZPpFcPy5Ri7uGG8rvnqDswYaWLZefEFVS4LwMctlBsfjcqf4BGU2vx
io5RTN/U9BOl8NXriEGJfYJyQNDYr3ALb1sw/stkiG+LL8tWBOoeeJERiZbIqnUD
TefiDLYs0+mfSK352G+MlkLtIJ1QfanabemeSvARjF1bnJI0oySNf2kCRI2Vvsvf
HTwXTBck5cSeiMJKdMVI2QHe8EjeLca1g2F9Y+qSykdNyKugH8AKUUbx7EldHLda
NLtXvV31W28Qdct68fMpIaasPgBl+zTpmuA4jBTw+BXXMA+oya6MWEk6qM1B5YCh
9hlp12hyykVa9NocYb4sVcNN4ufjf0j2BMCUqJO7fZTmZmO8510S3JkSPa2h9tV+
QlJLHnPNJJZHeF8v2lSdA0zsw2pSmZudymfG7grkSijmKICAnJYj7lOjbj7LnXZP
I9kPx3rIP/uD8AAr8+kqaTiSQpcMeilgwjYTfzVQ9PqaUxLVqWQ4rBnJayDZVxu8
9J9/xPMwrnlaKtr3yyj0+fRUWpeNm5cxBoLVhX97BMcq8fQYGKWEZj0AjL0tPXJw
VCXiPn4XvAUWCRy3PPHxCdyjBBPl7y3G2/D4WUdDBdIsiPXO2czD+/5g3WdjkHFJ
NG7jXVuzQTtSGc5vbpiSugI9Ih0cyE0YqXyMjFVODFvB/+VYrEVzMHf7IaZYDTLR
WybqwMVUcHyamaCzw9Ob2n6TqEPO4ecgYsKZtkpR63bsU6RP5DFabeWRnyMf3u17
4pldhfPJ/xfVWUHuoQH07mSkb7nvTnYD0/2CijsCzvHJhowGqer1FcNv1ByBsm8u
ayXMfDqt95WLzxIYxTPFhgI6zveeJTOZsXKeIRSD5UbzUkqpvd/elJi1s1X9JIwS
Y7D9+ngf5CIrseJvxxGaKXrwsIO/BWXR81RVYjpCl5TKtKuSRrd37ALk+bViCgTw
ejDnJVskMofPyfPk5co4SKFvir5aZWlv9klGStY/ia3BHzC2K1i0Ht7HVt6Q2AWe
JsXezCi78JrWf771vIqk/Gq/NfruJy5GHk0AT6uv7WtwZ3WrcYoEbc2lkQ5w0F1G
TrZew/Ql/7f2vF1V2eA/4eAsokhIp4ORXLiVoH7gv8lfnpGJS/Uogjn6R2ZxTDdi
v8sWrQWyIhz+OJgJqV9UT7cbGofhRk2wNSMwR3aFsOQOq/t0K/f32t3ucQ1hACUK
WaotY2Fba595Mk07ipaqn9MaliR3R9923E9J5XGLVFad8BjXWSW0mADCN7MDeFp7
w1Oppi3kJ/uSfChtZL6iyITfw7MTt3dmSXKyM/LfCNFjxlWqCdzCHO/ZxrQYWWod
WroPMUnViMUGyG+Bm04aiqrJIuUuK6zMCRVGwTHNAZkZGy43zIQzGAe8bMC5LuRw
V0dGg9DqhqEuFz5EaUWJKUhx8T57hl6HRVX9oygKb72YZv5WhErR12yzh+Uvabbe
BDlnYIXFZkqv+9iyeZo0EyDOj1uyEPoEn+l6UF5UCjXtAOsG/zuR2x5IwctogsD9
pyHv3Jeg0cp/BufjrutBkSGesEOvN0ZksfhwHrya4kL6A47yv4hfqOlRz43RtLWz
T5/dwU1P73jrHq0XN2jDkTCXASwE96ZaYZ/cho4WjhM89waGFW3qizJn7z3TEZFf
/qCATM8POeYQsFDrtdjrYxvC9FowZYi4xuD+gHawhnlfK5nXWWhRENT3SFDHRsut
V6xrNDF8qaae0bBGc6BUAbVGx9lzjfhgTYqonaJaZdKGgW8n1/f+VrJcpjEf7+Qo
RfKA2MxLEQxigr/EBgPztmVHJI3N2iVw9D8fejSqcxAnkzUD4lf7GC4rT51tIbpK
7CsXkf65sGv4os9xspuLzSvignXEIDJVZndkSoCekZgzuqi7CJzHyLgc+uGP0av+
VKMrtrnzJaK3z1vlWhHGcRh9ZzOb/33WYyqDYUh0/p9s/Jq5vVLv1iuk8ynA0TqH
F4IsM9NagrUl2mYkOUymw2QPz6QfLaH/uDuEuxJyrEyRqEXOEOQSzH0qeh9HRstU
PIwDg943rrBHfR2WQRzGWcgXt4Ag1iJ8X7NgJyeZiQEY/9wi5A1Z/5PiEwGuAxTQ
6LdJHwShTBSJ2/hcbBZvVUDqmS0kQ3oE3zCBDIEMU587H/XJzBWiOsr4ixSZciT9
7VK+dlws9yGiWMCE3QC3F94d7IWEkFo38nZy9OOVpoLlN3ihvGeuGAhoiZYFqswA
w5m+h5LmAD5UR3nYUd5WNWr/XuXEPP7A1q4XHoAOMH2d/E8GquNlGJ4PqAF5IrYo
g1RtnnkQEDFDD78tFzfLVpisPLG9w53rTCYUX1Hrqq27SOYo3Lx/r9fzYJFQ4F8z
m5aPGNgL+cWV1lhbdIRRf51fgBsNR1gNmAwhuTIzoIxTWXnqNW7m/VB8addKm7tp
hRaUmRapyZ9PF9LpdOWx5A1sMm+DZ94SG7MU+AWKPPK6K5Ctb1kBodDgCnruA4HD
hP5KkFjWPEhsS+AjcYbVRdi4mxgFkNbcAm1YdoVA7hS7d6qdp0deejXT1VLhNdFy
zW/idHgJKGBfOOoBLM5mo3UKGJlBrWnTOAWK7ezThd0/9CapRrkihvmy5E/J21eJ
PiNX+7WKgSGUiMj2nMEdCFuaEvJ58ikd11e9M3uf2T1ClAhCdl0oRQI/2X04AZ5i
95hggACbttL24pbafZrmgD1AZillIAF3J9tdZK8u9BRUwL37ZEAJrA1Gwud2jxiR
zU7rImp3PfBeohehayy0EOEbRRgRzq/bvCEEKVjpr+Zu9jfw6JiDNxvxqKZHTdeZ
WsMWdfqZpqqEEs5OKdp9ti167BNl79j3veL4cJe3xSw1RQpdol1LwnRSClIbANVf
G3D86qyAXH5t5n3CeYpsVS57e9WVfG+UeJvTGq5clqUAsWx2Dk+rOkUjcHhuWR4o
RRj9uCqeTE5ZOB0mKjSqi4cyWPNfskFreeOPBoYhKwKwx3banDp0nmuKcphJgtI7
RnHcAqEAYq9VE0H+8k5L20VGxbrTC+RGcQlXHwL0sBwlRvwcdpFlfpIKQAJTRHVI
dCpOeJM/NH9TS/MTfGlnM3d8bf+ksUyzKzUYe9l/0rFfCyYMw4BXjvadfqSnxgMn
9K38qfiS9nrIwP2+104/alsvKKbz9FCOndzzD1CvrqPcnrA5h0ejUKLpZ16BRNAK
dhVsKdtOzeVwR6vL0s0EIX1fnqoquNKZcu1uT53YryAWOcZG1sokpyb1+ZLLF2zT
PDxsly+3ST8u+Ecni8uBpP/W6pCII9WzW4lie1G5r0CoqZNkI1jh8ZUcK5WEjzQo
/ZwgscASbJJZMdAFY+/Jlx/fF3w9et634opAxiIvnxLpbhiVeWohgYxXtznyk/yQ
Tyccnl3/may8Vp5za+6LWz0vYa8octw1OTKnFoO5RpbmCbSKF+YaZOXOy4846i4j
t7HDrFuFQoWhDahseMOeXMkrEEE/x++aa2jD8J3iuG0Rp+lZ3bGB4Utr4XpWKQA/
ZOJ2v57ab6d/cwThlor0z3W4J/15VszYNDccHIeMRBfUWsyCa8tg9+TGzDEt8aiR
xzZgdh7FPNB7xsy0YEqGfjlbMvWY9pF8PgbLxKTXGFBXAODPQr2aPE042tuVF1IR
Qxdj111uX3YgSEz6ywWm1ZgKH3xNgmzPaPEGOIia4SBboMs3wVLp7pLfn3qqMpvA
QbQEUXBRTEKkUJm7DrwPpfh21q4Trg4A72LzRoVcY2zDWCQTdNDKmQ5QJtob9V77
smB30P4flvfce+4zUJ9JRHTSEPB683y18GzDrelExvd28998PA5CELF/nvTJuPNE
gsH3paRjsrEBC8LrnCvTqqElnD+B2qfhCekq07/7J2HImNZtIU2K5Q4y3CQ5bXcX
x3de8MBc5uUIkhYhB4nYJ9Wtl9eJb+D6Jd+oqeTcAjJ5Fl7kIc7KQ6yNPFv7w25C
Y3ZbrC5N0QQ+G7Y67yZXMwC/qGUc9KAEExOPeijqMAaVpJ7Jxz9MJWbOkNhcEZ7C
9QViSSSnfwAkNSEIKfe7c3C2mtEofYv5IPMxQsgxCkIIWGuJ0q13sETr8KtO+6NX
GxBSGVYKMj6uy6n1Tc5VE+bR0c3rfhfZRT6v6WGazj/kE9+yNFP688qY8rtq5TnO
6A5mIV4jxSYzi6VbRJDUHoeGqfOdjhILpBh6LzbIR34LZZYyB1qxp2kqlKtR0EDL
CGwjT6eKv4holZXlIe3rhugNXC8GF8A72SpV7s0BTkEB6TLbpDtYkLUk3KN/P/KB
xGS8BbSgZgMXweEbXmXtJkYnReqo16tD/ZqLSctM3eIib2MKSK+DJ2z4ucrf2Fne
+GvYUaVen66zQO2oS5ij/yYrpNbkqFWb2qlI7I8+ieiT4PjmaUcpg5huAW42j5+e
fZRV8D8DtqhjYnHyjC6+fYnEtfE1u9ulrmEcvPxC/zCxb2IjD/4ZmAdY3PO0qs5U
4uS2GXg3Dx+RzPNvq5m+ptPg5YscT0pD62qmN6NJqH+n+NI/Q2VZl7JqowOI+HB4
AjTWMZgRfgGagIr2j5i5aWXokB23XXrZiwzrZC3ABPmOugkIIjLFcg8UBRcdxcjw
ili3M95fIXIqA1lxRdyvIpHDsdn3+5MPVej4xRZFD3GLR5B+7T2Rj23msAPkaMDr
C19mQ26hxabvBX0Och4go8PsG5QZTtPIcG57RRheTnT9/XsU7ojPcstlPC1lqPeZ
u0MPdUf7GX2pl0qsFLFYyy/Q+6+FO+hrEuwN1mZ4Bvl01Xos+S36trtmlKPN0ep8
BHzj3NosYJVrfNNGTuW+UToulUOm66kTUpO8YA1MSueTaf7zZLvgyk1wxi4MOzaC
OmGBn+iWEswFCLok8sreFMBfYPOcdo4a2PGRFQpfSHxrknHEFlNvcfdU70tiwa5L
RrFGAV2Lhe8tNKaO3Qdwc97S+sPMSPskNNeIL8IY1vKRIbYFXVEDmHR7Kf8d8z3A
ES33zfKAimMzZlwcRvEAoOeP1ztuxtHClbsmq7sK/4xWCmRai/WsRdWqyLHzKqn9
mZHQpjnJquPdkQlp78HMu/sQGneGdwcNIXluyr/maQsmY4JoSltZiger3uc083TQ
o9ZXk6Gyrrf8eNYnIJR5sQCtMjko5bypq1Tf82oOdKiNzafXKxfdsW4n2Csz6ddU
F7qcvkgwsRL38CQ1OZK7DX6C/ULRhI5P/uDqJTeYE3Rgkmn7XInlqG5tGcNp8elA
vRDwV5lObklkL0f/Z6Ksjb4h/YukDc+A5wtqPQSlj+o=
`protect END_PROTECTED
