`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBL5abLACgizXIhN4r6HmT4tS2REbOxSjx/fbYDCKnw2
L35hSZGR2ymxsKYFGALcr4/zdlVWV95loC7a5YlZ6lCPjJtEaSwPr+xmzRiBke26
6b9aAuY+1PmoKkXE/bxdk7VJ+FnaBvhl+jjEnXUm5X0N1s+5OAiC5LwE7/XkCZHP
9yWPYmM5A0x5gFt1hMhBpKFHZJktBs3GsV5Ytt5QN3t819LGPTA4LePTuLF5kQut
hXzNqy7rqdYlj8/ieyK0I1zQSqscgAoVqnVJdBbUMbbMg2euYAnbJ9Ui5O8mIX+r
HgS7SzAktMHkR1nakXWBgUpWxD01y4ihIbINZB/mBejMqo4aUqerJyRJxe5xIr6V
YWu7jLlLBYo/lszOqL5bgHO4fSr1CSqtmzgsfSvs1MtDAsIJOerJfB9kLM3wIO9m
ZOIYWQbW/MD0mWUl1ZYTX+DELM2JCwealbyFpsi+a64KJqVLeA6LVXUpNp9ILJQZ
eJq6/3FXlCr2bfbS9b4WcwYzVWwTBg/gX+aO9wTk3UrANo7cjDv6nD1gdqtsripv
ONcPEWaTx00tlCtVOtCtaoZPMm0iZRWpoHuD1crsOdf3HWj/ckHltOnShOZQw9mt
RGT9Kgs17Cn15NnbRvi4e4W6n6fXp6eLLI+CdYflajLBupQdq5IvRxLcflxZEJT6
5Noj8myV3GnPrURwgviePq8NOEBaxjHjxTceorWF0C0=
`protect END_PROTECTED
