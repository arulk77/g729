`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73CxoAUU5mHdwM7onnmCdbLMwQBUS/Vkjx0lQNL/QzCgiY
dQKaCYRIWezs9rL7VjRTvtyMx172ifCb9kOk2GbHAAw8v/ltaKtXp9c93px3GCg2
tXhkSCLIGk9RU8deRFMdQkW47a4/upmt2RDvqcnWtTsEBHBoXgc6WqIw9bLe9ZU+
bzvHIkc9B7evg4D82X4blKWnuEu3P2Sjl8iuSPLVEuVGAEfW911bsv+1Ob6SeM6M
qB9l65aBQ9sdoy6kan1giEvpr2dP16pJ/+zV4+L5iyC7GjhZ1Jxu9FoCMJrbxLOs
BB2fuFStT99xfr39rn5wchm6SCsv7UGc6RHAGoMSeOh+5bbaiLWif5UltVXElxgc
nHBLMBLd174uSS+qi8FFpOvpvir6wuULfk4+o4Dzrq0NX9Ko0chIum2TZTbNIx+C
mfd0pMRIX9zx+nvtsW7apaYQINBGNNd009VDnzjxow0TaI47IEVehQrRMm+HtHdx
OoCkvha9jB35pI9UPSXxM+DQXiVLsX/a9dMn6/tkyfETOPZ8OyNXJL9qunrPuhYQ
6/FB5fDDlIei0twPqx6PZpOzEUtJo3YxNo+h1WvR8uVI0NlodtMAzh7uPqGttr4w
6bwReKX5OEuK1mfikCUGbVwhoozHiU3uaV1KfMRuwrxFBPbL8uoarmuAZe7nWEh9
TmgUQTORGrjCTZfUqhHkr47vFVBuzDSF8HlWfLvDlQOx8k8OJ9x6NwyHIKgQNBn3
z0lkLHiOc46gi5QuDEpI6kVkqxCn5D+dl/uJQDBLz7QDLOIs6qSXUO6pfMMGXRPG
a0iS7TP0lJQE7sBf3mw369Qd5wzAijJoYdnKVRTHik2kX6Oeqmvdc9w+3S2WUgXH
yrVypLnpSF21QPEzkHwEYpMsp1c3QKPv9nlYswzsGJro7N7hYrNjSChYPs9+vLZd
1ofT+wGxo8Od2y+uPY1RoqOu/+dxoX3VmPuL9Ismx1mlolLt7/pWj6bDSnAZpNk0
1Xc6HF9/ME2jGRAJf4vVDEUNLcfFBiw5uYNAiihIKEtCX0XgbIFe18SB/o91MGQF
F4ClxlHR4ePFMSOVWcWvlSvAR2P5C+lCTio9kaYu/mlBp/UvcwODm08LizXHP3mP
j+gaEi9mJiTUlGIKa92Wead0z9vy73BTDMf3+XCv7dFBgu+7By8gzNNLTuq198s5
IjISelmTtR/99ICU1/y1iAmj5FpeDjvSvrsza8EJT0fJEp3XVZsJyCyooXOewrRE
GPSWjb4wIgiXPHclqs8Bv1XLJCkoQORDW3pBwiAzoDdGMMMQ1+sAoA+v5tgKaWlN
3QjTESPya+/gMDMdCiSqbdwM0sBYfFuATTVLfjvpH14fpAXb46A9DCKccaMLtM5r
YCzhxml4fOdTsWMdnjZuP44HDyjBPHqqoBJ+XT9fi/BgfUA7wJ2Hntu4UT+oc1eL
BE1ko+Nuari22PH86GppV6hCEMSXYJu9qIe++L2+CpySJygv0wNAFWvHsSaroaas
0Vu0pev8OWqP6rqz6CoM44eEvFzkVuWewGNzgcg6KOjP2INbb0zfJzde/cMsKd5A
j7Zp1D9wHPOqV5ZHshCiSzefClYJSHJsVhBkdGAmrsoBsLj4NpkOe37QIyRNbYM4
7OpZN4YTb03s+aaa1fJmVjBwgyi2QGK44t/qJv9x0vHRRsRFZ+LUuK1vp04Sx8VC
zmKEhlfdNLN3+3A1Ob6NDIqu2OPxjqWjBhqa9QD050QlKtVzeFb53ZqHAILZw9Lu
YYtWR9xg561mn09TsPHtt9ZzXNq5OIlIS6IR/nv2TC4tKVa9PeIQXUP3ebSU5tr0
kTXu9DY77cmefe8A6CEuA6ot+nU3tLS75Zwd5orSZTPdczMv33uag+A3e1StAhOn
W8hQ+CgnzbN+7lpMNSdS5UGEcoXw0s+oOXbH5b38+IGr/Y3Ff4peuKx+R9adaBM/
2uQ8F/LACDCv5w+U3aF3G1D3PCo1OoBo0u+3iD69OYZL3ywMPZuaqMkscBm98klE
tpM5wamLJz61//mS/nGG7mymCeVg4Bt+OIULhPzrAI3UqcdNqB/nSOEwUx+jt5Ne
BeDR0yu9wPe2wUbFoVFp0nsHGHD/RxeXaAyJOujet3TX/FBlgEmjfJBnxZofSweO
X1BVIOLGaplntuY5HtwU7sFYQIWmxD+cu1FAHJpDOCXOuIqPSmMLDdp4sU2ql3XQ
QiN55fO5aZaSbdqKR+mO2xAs2nbon6YrThVWd43aJ+e8YVQIbf3YD5IKq2l+WdLu
G7KsBSHmflGb7cKa7TM0L39g3o2ll1MUSoplxSD0omcEFN/6wLfuxEtDXYzdddqH
hcl6TE4/VxajLvc0shcnJfCF33Ba8gpVVQDvIGBaKSaMasaAqDacOEA1Ji/icA0P
Fg08ETmfDcjiZiEFpI3hzIb1vE2bMu4orvKLlJH+P5tEAd7X2YjobGTuLS0clvkY
qMLQ9HedOGNdCvarRCWjv2KmYlkatk4YpVsK12Zv6pGEgv6utcNrgT0fBdTQMDao
pvMYweNgugLKII1wvFgbM/JR9OlEjV5374ifui3kxu5kZDYjfg5/LO904p7PzQNM
klCULZFWHJ71DDIMxS7SBdhYhPUS+y6fAL8huDxJjj6kKCVi9v9rwl02T6xLNpiD
Nji/I4TLncSJxsebuqHH6WriHdIYtODvaY3Q42f9nPmpktEbQ6N9xAiSwnEJc10O
+L4GzUH5QvqhywbTkUy39RgXJRPW0Pv5dAgC1UJq/VzxpkNQiWD4h+5CSgJ0DYtz
JnsEATpOBVHUxEZSq8r6Q1sT8sfdzU39ENDNZVEkMua7VgdGnKt37LkUjsVwSYxY
ZSnIQVMLLFCY1yCgIlh3dvjZxypm04HjC50b5TpLuauaSDJ654ad0pajWPCxbKin
/Oh6fakr7Uhzjyd5ILIZWF5X7MWLETz/z4sDDPE6rkF5iQTSKvAtBp8co78D4NKF
dqV154osTzTDr6TDcsitocnOBLw03LljuF7YUBf31sQO6FBqoMQt3gXZYWagxB9j
B742UVVbm1+5bVNss+vFyLQ2jdI7TjCJK2BZ/Ai51WuXcMjXffj6YJ289Om7EjKp
D/8MA0vxjiABv46bVyQW5KG0m2e04+/QYHK+lZPS47AQO+5wVHCGs4LM7SdIGyXo
nR3dK0XKyWxA1JU9L9KluBaEoiKk6UijGWsn/X+DibwV8YUtBK66BMEwicxxUzmR
1cA7pfoCU1FMZrV3Y/UlXaxCL0LbNXU2+7r25iYZxE/2OQglBLbaBUVg6mdzTysi
9FpCEsJ1Wz1HNx3J37OoIqzyz8xWRZSLN2CCtmQywfw+0EHlYcEBesByb/cGBpGW
ceBKfIHlJeHS4xChsZ+eBydqRN/g7b2HGkOgtSKvVa2EKO6dRjAmZiDTn5oUfW/P
lj5hV+35K/WAclAmq8b8QJZCGMmc7z2yRtJZ+18uQU3qamMrfOgBvrpySsWELwd5
RTA4fC0/wjr13ROqRUmmf2pdFdNNt84LJrStWRtqOnuoI8CmiwKdWZ9160sCpGdU
vlz/Uc/Yci4rHHdlk5kfh0HYkSbR8TWUo/Fgc6NMWuzjDNsJMUgVY1OJGNHNvOCN
+yg4rMPp3/aSPmynYNrKJskDusswhbtC/3i8e1eSmvSEHZHEs9/ni62DFM2l4Xxc
t0LMVWcU7BJtK1i9Zsdcr7/CHC6dX8h95Y3KWWdHISBvh+smHKFMD61bT4qEtBCn
lhTND4GMoGSLvU2K3NM+nnXusfzP79Y9cATNRnmMUpaCoCQHfCg9dIw0Vmzsf2BG
Pt+1iSqvsAXEJRPdk8nqqvAugLfGJmx8jZXaEWl4K5Jo/jaMTaErh4PnfJFv3lx9
aNVAVKjSo594KLvuUXm/iw7H+tdNMfE1rx84bU9IBdBCPV+gMdHahljRK7nvQpiI
EulwIQrrwjW1Gn7SQzsDmJ67/512jeRJr+qW1GCAuHUhpH2/mOjdGeOw7/9Ce0et
633KkHNuhekBrtoCgFp3W09tUkmzMTYu7XFNuHp3/pKji2UcQlrgD2fRah7krOZB
hUR23EORDeZmRnU0HqeZSxlts7dmK7mGxgDSBWijmCDGrC8RKVGbaygOK2UnqKzL
D0IF3L/hiZsMVQRboiOcF20qZ2fH6kJPu22s0Kh+DLMd4rSMyiNj9E/a9PvAUi/w
1Q3gRo/BOi5RvIVNjGpLpaFq18f0Ccd38pSfTr0YvY4=
`protect END_PROTECTED
