`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePelUWVjzFUEORLu/VLhfnJZIc9kuXBV3tk2E230O/rn
uARAx7OAdYIfQ6DGCatOvZSTe9sVw3acHty34VclkOYT82RBG6NB7oLwXhKAswOx
N/Apdo6liFYh3vrpAFaYrChg+O1KfKPMAFaUxeu8VvRJ4cMq7VnVAXXOY7pLSUaJ
5antj060atX7wR2LLbKFKO2ExhMrlVRwghXHduQmQbSSwHNuLp66007BjoCaZU+9
UYCfMqgTkZQXzpgZZpwTUOJTmVjnfJgtPQ+l7S0OcpnB4FGFu0suew4A1ax7Tbs5
5oLdHgw6W+dAMUQ9smZGqBEUBU2QV0IviptDozJjNYXG9lap7N/BKmt8ATRpWsUf
bo+9G2j80X871l3dMZX/Tpi6w9mgkwaQbQGVNjwsgeE=
`protect END_PROTECTED
