`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAVd9ZtT1BbDv0qZ4duslFGPvPvD5Nyh0l+/v9CS2ySJD
7E1IF+PP25vfgoNR3PFAnCWT3pT56fuTiVQG+xQ4VXFrfYenoZENeAPYJHa8Ujlg
Vk2ucQBXcbtf2ORh7IF4QmdC0K35qta0gUvtCUKlCptRUwklmsD2zcKd9i/Mt68Q
FaOQl079P0KrRYxI8R7rPu8WDgjE9YBr331GTStnE1pB1NHUaplK5NSHl260z+es
Y037hcGS2WWsbV3MPzDf7DVRnMvCKlgitdaE9kKBTryXknv9Sj9ybVUoi6tjUDIq
Vata0ZM/U/ZUwUDsnGrjRi2UATej+fZ29rANtJbY2gyF+Ow1kgQh6fBgLfNV2R0K
lgV4am5eMyjhYHxVQzOohwmnifWMIRjqFGQgJlwi9+p0swiAPbvI+nKi+Ba25VkO
89/whGyCqLF6MVbT9bdLJD321A3sS9LAnEdE5wOJvmI5nm1gauv6m58H8brutrqg
UFk6mkG685VRAY3J9iE6eXmRYa0Zc0luooojEnDZRgWbcmN6yIp4HRbzEhXV/tlt
TPRla66luM9k/7kNDLjGun7oVplrxkFkYcXZ7CrEc/RL3xT67FVjQ0leogXr+LMs
6l5Qm6hCgResnfSkCkSXOIq95jHdYBDs3AgURaxrq1T+yrmhHKVAG1PX4tIa2qCr
MDSZmunWrH0ttY5SbFKAAnS0vGmGWX9z1P72N3HvhK/Yq/9daIvITANLaBVEhw1l
mLBaDq58GxWCX0mN2QLEum1fHOpN96QUVgV+UdxzfMKj6v1s86qS1pz+o6VIgizp
Z5eKvGtYJ1VcSQmtK/LCiQ4YhVnA/3QpL2ws9m8if/lQCuISvqTXn1yUHFnE+omZ
MEA7cgNiBTGdcA7ZlJ10jmCLzTx+bJkiHGlzytb8X0pHWfMe5aNFu4Hx4SIoEuHN
1DwTinGuXtrcpRjiXoFeB7RSxflq5xI3WKROw7HnlUTVuZNGzqCnjBv1MJ4qDqq5
FMlQGay2FiPH6RxGACAF/EyQWWpH2qJ22VVr697S7XABdEVGQMGtLkoumyO7tQW4
HKvHhEHgMo5cnRDyod+sLTqnZxhCoxIkXUsjD3+b65JEwqEyJLpEkh57rhATU7CR
5yPGQDvh4zRjwcKYZ9y+/aiwvnXHS7T4wSCCCXF3ZGWusrw4vBmj7scPFlUYrgDB
mgGG+g9oYlCsY3Vf+WklNOkBnTqk8qKVr3RXT0gsZyqEMABrVEzqhzXU9lG3NTOF
auP/4BqjUbRHo4HcpIpLn+TJpdhC4gl4OAF+p2mE0K5pQMhHfBEGxMjiDOVgtFGh
7SNK0OAirmhyaP0jallerL6v9eD0v8xpN+8C+BPDLX+ZhMTTSVxEsq2eQlXczt+F
2w072dKuFPFRmfHi17G2jOwYUjj/A0cIX1JM9B1/F/5Hjz6x7utzEJta+jWbmtn9
VZa8xbdlXeZTELwVuxbiXzCKIxjj2L/y6KfWOTuFZSSQ+EqwTIVi17UQdMIA/9MP
VIvPYLr2RgJcji530h2kk4WYpO86t0LHFDycG7IZLJoA1pdo0N/RrKWPu/emtt/W
3JxpaLHpy+xGscsPZNIjNuHSobHhftNo9IZeYKb6rjrQ21afoRsuXtvdWZxrhFUU
22GeE7CoyPtqg3cBXm8uIkidGbrex3OrnVQvOAFogzB7mn/oRot96xPOycSXMHJt
+11Jfkm2IgxXRgXF69Apnb4+KWDjoGUuosMzP/kUkijjO3Hdclv0mT6eQrw0mIcC
+VFd8MlHLRqoKqnwaLu3/+2UegKY7sS2dmBU6nGlxxaujHOFtXHadjTiOf5aXuIL
NiN/AAtvzYs0li9DcHaFHEax9CsTlftcCuuqqR0m5enRcDaaYxFW6WfoIXeqISBm
Dw+Ua5g94sXxtjimz/XSNd2vcZIgXWrwCHfdREr15r82CsLqEwhJWGW5i/GYo0Ca
r1gQrMk0pKhylLd+pvr6d7H9jyq6ohBgWgAbyAmjXH38ibA89XpK8pXVhDIsS3IG
SrOT53pyma9qLbN+xsw1DFuUctCfiWusgc/DFuR7Esis7AvzTmznIDb7vN3CqHJa
gGFl6ErvocCUnxWimv/O8hTfIOb83+YTkcdlMNxcIMkIgo1ShgNmAjKRYEt6QW4E
B/5Jl1AY4PQmgzV7LNW4nfwXUeWJvV/COJQKJ8u63ChHiUuIEKv3bmUSG2F6oknK
o9DOZnXGyxOHbr35B+5Ira8DQ5iWeuj5unLDV6WBiLxUiyyIh7yFWw1gGkntKT7N
lTVojmxyFgRJKJsCRP/OqkVgE37i9V4q1i/LFVGWi2kqof+EqXonUNMFVQmlB8vm
U6VLExLJEBe4UkmVzPKFoUbGk6WJnZenWRpvGrAZxtpIL0BgeubgHcNAyT3ursSo
QVmsKoe6ODFe12HDF0ko3MZnlExji26EiH1SNcE1CZZYNXa8dmGFqhZOFz7wlVDD
okGUrYD6iGNmB0YECB51hRktHFoneDgnzechmUpKf64B3dlof3NGH/kAqBeFb24L
fvmtakUdVCu4lB5zvi53egvpcdOnWUrTfUGsImPMrGPGsVAx52bHGMiy1NlxH7NK
CQUt9lc31sVtwv0rE/YPpDLN94DTL1infA+Qzpld+Tb0ew2jta8UXuyR9svPqOjg
aBbE6gsedJpieAEpqIwY96EO5v3kYaI5EYUqNueZ/glUxcSWagt5hor0MyT/GC83
2vQS3XIAfR2/D150pfvsumspguDgtrHlpF291CRMbewVZoiqgGDhqROrfmrTKcEq
1PI2PBXrLnIL76B+6m1hpCf0NBSYjHREliwBZp2ymrk=
`protect END_PROTECTED
