`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
scWAwqOJbVh1wRuJbrViGV3n41RSFHWzm3iqCLuZ3Jc3cIl6xn9L5OBFjB0AL4Zf
BCltNcpqcj4iFAmDO309Xi+OSEMBgiwM2GQ2PHe1OWCvfM1gcZCZ22o83DHIwFyF
1MLNsil/4O2zWESLmXKU/N52wmpS2QrwJXP67MMX+Kl1d/qz0GNIQagxmm/1de15
`protect END_PROTECTED
