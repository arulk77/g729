`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zkh5k6EQkHFx/zhgfcQtFAoCt9+Lzc6vdOSrkLeG4Qa
hoWC2LUU7+75XBFGcvWAmnn5zlnpVtqjL1IAnnci4FTiP4uWzRyu6Jzi4eVQ43f9
kJLOdeWlAgaO96BVSsUCx0w8xWbMe4q2JI2GOXfw3KVJWE7n+13vjL5ZQa/pI21O
cs31+aoNW8sS8uJZ7/nv5prdKaHxTaNoSA2rtoiESSNXbVZANehEXoxgTBHvpWww
qKXo2Am+SfGSNm+8cjoFiPiNjX+P29wq+Eb6EhOf/OW89ZuwFyQ4L4MG6C0drZ+0
TympfTsrrz/Ec4TWTrZ2T9nuIM14JpLLzZOfrnE/yyiAIZiUs41QlIHZBQ/zYQE5
ZiAN3dLNcqVm2jmf5q+sXQ==
`protect END_PROTECTED
