`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGdy7aYVFC+l42WLkh0ADdshKNesejs6MLsEa0WMCOTR
/OxGDZ+up8sj9JqlYITJ/NKZ+QXgqegJwxMO5sbs+QwabL4ByYpVb/xAK8bhaAjf
bxhSOSAbSzXwMNMIO5i0uvUDF6pWpEp6JbfdZGL/C45QUTgXY6+ITDjL7+8+ZxMg
T7Q9Xqg5Gpwq0Hax5na9A+37R/5vuuvQ9tMAyOkkgXlta0O/YNrYm5VCo+xBRbVP
pKu0B+YDDM0nD9e4JpIvApSB5mlBFH9ZKR2mNI8npeEHUlqKpqYYZuyuL1OWoZH8
SCkI1CSibRqBwM2n3kKBNj0eRlxKisufoNyhI0ZFKp4pQ9ZscHO7byO5W1xN/1ZE
DzZ3gGQvIfj+P1DFFJbJXXptUiw+jKDL9iSuAssmzmN559QTSBcK11jCV4Eug95H
eTZd3aGdpqqUOA51P89fmujMdHwEItgTBduWvtaWXGGD+OqQNP4kSJai8KMwe27l
`protect END_PROTECTED
