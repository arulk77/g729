`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG7iY1gupGAWxSWS5D6q2ihIcoHzNrIXW/39pM+nHYVz
q6iowcqko6LKnrShl3H3LgCAbAfqu8ozUjFkR56n1qGIFA073EuNnQ2dTCHFZm3e
+KvctIT20vjUsxTUIM9lVYLORVO1Ol9mLwPcuKWNCdvmhioXvevJd99wruPCGLlY
z6j+/PHVABMKBpLMVPIV2iNq9RRl1qW0CRUB62vfc5A/f7pf2qV3j3RSfp6/Ut0B
`protect END_PROTECTED
