`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
f11uP3tAS38J+2XEq2c6cOrEPRabbgkmqmMq+8HlfQR1pQwuZ40t5mbrLrB9gFtw
9fbsy4o9rbKrCR7W3zBEBM7Bk0/miLdXwdcDRlrZ2cunHIz35kcSK+w0zTmUrhWk
5Mmtlw9iiE8dym6piEMCJdwuZfegsjK6i80pLUinJFkE4M4w3votOlXFdsKRAoGU
`protect END_PROTECTED
