`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIl3iIlcDE66RIAtQv1MtW5HRiFubz4RiY7SlyBUJet+
dX2wP51xmVIPtaSXDHaTdPY7uaKaJ54sYtnHc3AfaYfw0YGqXjoE92e4Z08W5KgH
os1D8ivM+553ty5BCywCW+hNnibfUKW4/B5EpqfiHxQphUBGX5isqH6eqwKfyH9g
ShKiH+rcQLwpnZthtiy9G+zvvvzYkPFafiW3UTUjkEcRn6o6t4wwXVvQLac/RWXQ
xLQOhUWHW+UAdGEoQ56nXLXi42zRZuQ9gpD6ycDyWHAzoRYd+zh1WDVajcOPoHNL
Fn/i8eqXBjZrGnioxD1AY9Xnt3p/qQxk2YWBbT5LE3yh2ztZ0bHvhS/5pBamgiKH
1JWRhU3v7JIrpGJ52OL5kYLAx0sTWHjekmI6e1x54jHEztDIoI/CavTUwq4MDC1V
9RUnFe8hgI2KazG2am8GwMhsPfTbYUkLQ56EkyGjhY0AjX1yIKsu84gxGayIFxcL
iPC9LQI3I69eOpnE0d1pifywzepzDwE2jyNtOmEYIGogVMdwEMa+4XZbeS5Cxisa
`protect END_PROTECTED
