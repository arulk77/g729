`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN8jUEJRnJ6q9ddMvbxpGeHvV03s1uMmAbR7wZRTpoSU2
b0stid+lGToXGJShns5S/CnJaxfgEV3E3G+Ls7L4oF4D8UNdHB/ssPGxrIDQi7HS
uyQbCS0X8nslyGNgdk/plU1vRQNNBpgRvyWMTVsqKuDNnOjpiFvI7jzwKbNQpyty
PmccYS3rqS3vDgqbOnRL1dYf2mSCZYHPmg2KfKoJlUTLIbB6PW/7YQEoFKNNjt3t
UypESpLVHN2DdZPIqHspxv1TSphZ00TrsKFrHhxwsfVnT1AWkNi5fcspc3KaRyGZ
PWulJBo21Adh6evOIM3DKWvxcN+EqAa7Fcwsedi22QDjC3H6Hiw7/lyN7Sn0OgYc
YrUI1CDi6JWEDBugdz7rOnkHKfDfdgud/r1UipUvwi80FSg/2MEubJmaMPzeM3Nj
xFvO0HJbMIDXdCzoNL+VBkT9/mD8OZOd4FrhGfbdd/GFlxldt8dN663u6+psgYM2
CA0FCkNNCrmh+/V3xjeMkM9GC3tn2haJmwT0WyvoV/0sk8R0/ejWtKZY3jvsvi88
E4a6/8zoJAYf9yqewHkmAdC9F1mbKC0DvEPAB1p7bLfVrl3FOE+nClRcOtiwxKQl
peLjZRSA9O4SL8f+QNO0dYu2J7/Eu0JbDzYD1CktJEFID+AzvQm8rkJtIN6vvVH+
6zTdT29XuWjlM9d63W1qggH36t0dQps27UaKd9VDNTzLAu/eFL6gPbqON/fC6fea
aJkEjttQbtSAf9t2wuxjb2pyxSP1eSBnsFRt7cwLk+Ct4OrKbf4ItPmj3tTluNRB
R7yPSfMHj0meIvirTc6X4IbmrgIR4YFR3SGYxnrF6J6hcmGIIIV6UIaJ9Vr/S3Uh
XfRmZZAk4TH2XiGrqx1xWKaTYkJLs+AMH2FQUYYU2jpIOA1JH0u0hDnH1OR4eatO
7yLMYT4XgaYvX35Uu3bcDOssiOmqk4UQ2aXKF9zv5eXRFtjiJoyViGgZb0mj/y7z
lMo11MGXnuxDnhwmPJCgBgb3qOpnTyypLIJ07zSVtw+nBXjfihk7fXoY9p9gEzn/
vAfrtJYpGuiv5dErX0h+J03j8Xjjb5eeHyXWJM0OiE9+u0+skq8W0c30mfL1BVAC
DxodUlp1zXr7iLf2dfpW1H/1b/bgGVz6J5jq4/lz63yBHNaNePl1DCCuCsPCSBcu
FyFgmfsOwlFSlJB7moxHeJfVWyBPurgUL2WOYuzt5s9gBzgfKGrFK1MBJtNEg63F
CMQ+y8UEdN4CkrKNiTZ4RBN05mD6fWEazyBA/qhQYJCx3GULkxyhJiMaWBSwhs6j
eTXpnCPMYb+dGcQUBbA4qpF6TixG6BvuBq6CQDO8aAeXSo8nre1e5SRHy0wGHbBU
CT6lCr9QvWjTyTaTceJYcCI0EzOzFgMaje0T93apUiLLn1QrhGwNqpruKzwKH7kT
95UVxCSbXV2pnWOkQUpoIX0k9JwSG8e6m4Q+zh9/TUOAs7YRdsdWEPZWxI0i+7gB
SfEM5viIk5G8zKAT7dwXmPVEAp/3rX8BVYjoS9hT2s9aeEfOCZJlHg5gEFpOMAMA
mCvh/HQAVCgx1O78uOMMTBL/LUZwJhmzmd3ohZpbC4/xkNGlNR9jn/OjXpLa4TEY
plmhtuoVlxpGHZlfg9U+9mSdX70EGkwkyx+mz07P6z0RLqFstfFyOgrJbvNfYnoL
rsv5vLXqQQY1k7BaElpt6ZHIzCGClRr8Fl04nXxz7LTZBpIaY1bkqP81GoyBaQsb
RZDCRtP+7rKxmT6mWH4UnA00PFM4cveUDjtEucUgco5qRTFmeA1vFzpXwKwAruS8
uF6SwxIWCxQVI7VuMgac594qVg/vHcgZP/qjQsHt5XnUDN82jqJYSMGPvN+RXuiF
DP9SBF5S4pVcc+ULu+K4dh4V1NAHduMR/FsrPNWpKCbAadY6u/2PsaJoGiYbabhU
nOMx9e0tgv8yrI/wcVaiYegcW2D22Uyv8t/PLK45Sj1A9s9HvGEdfQopqJ//Db4X
iOJ1+hbOrzrlR1ttRGqcTH3NP/XP9AcxPQ4mcsnE8Y0Q9yTnC95PvYFyVqItvrQd
63f5q6zQiN9LeWNZkn2/7zZw+ZTUg832haUZlqFlaxyYBozFtPOZDrysOos5/30n
p6Ob04vWUBYns6RBWmVHKg/0oa2ViFjsaF60juPQyV9ZgeOrH9J5al/ytllRsk3p
Y8k5h11pnZaTS1tmmKYAC+4KHiEClG/qasaOq30ljHtcZ5L9oiN7UHS1FUjrym4R
/b7Er404LTDSxkf4vASa6CfUQxh+2jHD64l7unJ3y4flex0viCXR3CZKARQc6n1P
63yMTYHnfwT0eEpbzkTJQJZ53aV/pKMoWHZle+MfiUAevIgynOmfyY+v/TyP32Qo
L3j265YrrRRue4HBPBMQBYJrt0fboqhdCzXJbejTEuFPRYnn9pC9eF1v6kv2s8Q1
tQhJajq57cn98SrHM9x+0c3IgSZmGafdC3bFa6N4Ky8kp3kJYT4+zJNrrfa5nD8q
TSAHieM9l4tdGqpvCuvt8EvqMgDsUWvzrBY8O/0mYmXO7/YxByGKFGLkL7o691G5
L9a35XebIIsH+LkYUUe35UcZSm4F0jV6LcC+4qdrO+COXca/oc+zKeU8GXysEkfM
uP7bV1vpIm4HPpeCW84qrjwrD64SQ+efd2wgamDNscqE9avlt8ThXzhKqkzS+Kra
fkuJU+Le2aCHGJHYJDVRraUSudX3YxE0gBQAaLFtVZuVfTYVsFvWoUTbIs2yX+Sf
ufzzin4PWqHjMEzqtUnAoeU6vKfVxzPUXR7PwArUSYWM2SVYoHfHy3+2LFKp1jaP
1Hg3XgdHNIrBKyEvKuaN7BqrR9spksww9tUvDe1/ccVPZD0TgNga4MDUb+wJQQGc
x1lNDgXXEuDmG4TzOKWjihT43OAXdEAT2bfNu7OYQEd+gkAxNldtnY1Uq0OhtCdO
z2w9PgXXIoQJ8KKJIEe5jT4G4Bgiriq0hmPGkZxp4bB5RPwOIkM+s/byAXPkzd7Q
knC493jNVdZinrWe/MC0P1ZeEYx8FJ88RHkSJ2U0p7/eN7dNKNEvpRNM5VNGE9kA
vvbxJoLYnaskpZSZXl/x4hqzZTi/4l9aW5YOzJA36xSny+JxdXVIZfZCX2M8HcGK
UCVYlwry/SZqOswg6mqQ9Z0XmSeTFuA1Oo7hicdd/ft7eOiPkJGg5QvTmEsV1vPs
Mf8i4CQuQQaYDgBz/RaQkUGu/5eYe1vKWIIuw+Esk/IUYkgOz2Ap4kgliBJgUofd
TR5vfX+bXdBUT+30B7Hhvsz/xh7pxVYfCzac0MD31hT07SHZCdT8M80Mohj4wFKU
WpjdpARAeXF9ekcIKeGrQjmswbymh2DfA8e2g3SduEglosuyafty6hunXBoN6mnd
WKIZy2tpHgOD1RZB0eIuR7wPVr21v5Gd4d8GJBjZnDjwhr/atxClkx9UY1DjC7It
Ivq6XxBk4a6PfodLFL28dTF6m1MTpxG3baypGx7OXCc3Tpq7XLX4TBrs19AttyfT
fc5xPqj5DaLJl3PtbFW1fC4M9maVDc5Xd9P2SquCwzvZ55PEN4jai6vz48X7j87r
EI3fTt/h2h3lQEeEwzgQbi/1Wg+sa0265rzEPPutV85UF6wFVjRVuNZM3ToNGrHD
F7lTjEnVQV08lNU8+H6rvq3llZOnHXkxdA8kWgqirL0RFI+ydd63mt7XQfB06aPA
XfOL/tgL4wSgpekNMcU/qR+uXAWEkOspygRVVWTjR4SHO1Nq/enBmVyo2QBy+sD4
FPWATWs3TKbUrAQSCLsZB+kZp5rphvB/DkuPbr1Rc77qcPJ1v3TRjXwBxcJwp2q7
SkfbuPoIbBOx5Ndn0Q4wynsiit+Fm0v0Gztvxsv29BlnGZhcSJQQEH63tkBgZEE+
KRNA/2e6Ss7JzQnZMb7MEsY8+RbWrFPNtxumLpz7nX1+XYwJVnbfRIFuMk1k7IZn
PnyrMNGfAQzHOgrUKxdz+o8sX3fLfnnZhl7MjKqSmnuaGr4eKTpRO7YUHiVRx/I5
mmwRPAuq94I7nS8MVkYRCHpB9d2fu+1wWhJrICU5X8CMxG37+pqOE4Csb/KDrznP
LgGYih6pr4ywUYvS3AiwfO8rIYQAEiHCuzPp+gE9y8hZtVw2tsMAiSkV9kFncSYS
ECEeGc5ooieAE9rh12soGLfNB1BBl9qggeVQFruM3KrBU3QxeGimConeSB0/ZCEW
i9pbRSAPWKLzvpZ6GbuzATTd2jDAadBywU6XGxf9Zt2Qh9F+xiVZQ75lMN69Vb8A
FlxzUshQv7i+uJCuS5MrB7mMqDbSj10N72kY5695+fq6Iluh5YHH0Z0glm/FIcSI
Ah+W1D0C238s4ETfKKQZdPwuGcwm59KEScmiqpKcxmwpk4TaSOyvOBff5gqI4Ij9
v04/3s0s8bfzdJ5H5UFAtudsG6xMb97wL5orKuL6+hThNhOWzFK8DNvSWWP3I+D7
Q18GyifxNgsaOx1A0BN/AHvpRp9Gw9LY4jFZKt3I2TwVEfZ4s1MSxxf9rYGgY9ml
jz2QwDpn+boCm/IIU7qYP33kJLEWqL9LSHT/kNPtbgLhVyYYZ9/BEmDTwRAK3tCi
/NHk5k/MTWw0ZHeFV+ufdQI0fbRRwTQbEUGP3PkDMGSFUqjfhFitEDgH47h5IvtJ
S8J6UpJ6YisP2dNQAC6DCwxZ03TQW0emLAcJ5bY/6d4uV3ZlvPvRAO3M4d/NCDYI
seCMhIYKEbYi/tbqrOnQf59PSN9KDBX6ScUXZeSbtrHm6EiyjIc+5xu7MQS3be3s
htEguaKTz+S7HKt0gz72K187yCBTCFPDZn5FtVU+YoTLZJ/TJWiDFIdyaHCn4qMj
9bxcWlj6LfQJOqfyVmG13ABELrrzOz5b712qb32wwl1co52P1RWbDkHpZgezDwkF
QCqMFHDkjQjw4sYj1/XSK/cyAMxg7as0VSGyZ/JwWLf05Km6l3Q+68HZC6d8V9bR
E2sj8PzFLQDWJstND/MI+7QHGvL+y/In8hB5BnmYgzqcBzAWJTaZePlhaMFFQCeJ
WYJm0Sdhv+KXisASvk09lQMvWIqBamxIe+0oNp6AJZB3QRIxgHkpuBjz1cReu2Fj
kGjCF+rNX9zHiPL1INd5BNorS5fJ1FEifPD1m+KvUbRF0yzhn+mop1fzO0eA6t8K
cLVoc0EvY0BwC1TFkMJKM0m9OkciBtAt8YvYVDq7GzTAwofJXMx7Yf10GshOPbjj
Nbc0QkUQdI7fr//e2vMS8cgYZ/9X0NIks2g686/keuaYhOsASCZCge7eURfetqab
mLVby/GOI0BdHwi7DsK79cR9SONSp04QsuENGtPkuHrWUJzn52sTBj+0gpoEkCUo
AfwHWlNIzPxHxCLsAJ03/gT2qYowEU8sDdqxJP+7R4fKvVAzGc0dwZNTmNXH7iM2
6ZHQtMt5hmh3IClEbsS30TglrbUwd6CLzdKSMFnebR55dxR51jaKhZbp5IDEwlQV
o+lEi61BBvpmfHldPjDo3ntyVt6qGk+x8o29TWOjsMPTm8/oFS6kMs6oRTYQqnXl
GcSYkOjhaVzRGgN800BBh6widxqaZ5gokx8lzMbqjjXVylT9n63H1t5WX3FMZ5eC
hIlveGk7Py7xvuaFPClOAsl4ukpwRRWzoDhIg8fjMRnOrXo3EO67Y7Mm9imCEzcN
4bW+a9fyqvg5A/Z4YQeGtNV4Ty2Re2ITPaCdAwPMX5WQdbR9HPgHXVFtPwEwTPGx
wvPttd40gW9GyUc8Wp0woZRO+42GTTpSO19lVcsk/fTFnt3+6MJXS7rWuOIBybto
R5oOlcfi5s28vY9VFLm+pabeXmUzOksO+up8xm/gI9nbzySwtc+/B+ZZsOcBOH/O
IMQ/S/799ACESp62Tp38iB7fWfdeM+yKYmSFMnFfTjoOy9q9FocEMtCxvi60LHF8
IZD8WtQXX7IyKhNZv04fD2yBeJvpHiq09/aEQGr/5/4HO85VUbhNhv6V4LDo5xkr
M/IesZGepMwRwhTpH94eJEq8hR/WpIlHXg9tzFn+FCun5QqArtlmxGqodYJmKVpG
rBPstuWj2lDwxBpsOw14nCV6b3OI4c/+7OK9PUHr2qAqKeT8oulIVL1MYWpv/QHC
G+oFMboJRNYMeWoBisFUhvet585hvRRbJwTwZz9ZS/tkBcxw/sym5BBIzje/et+R
pmnM3OrTbWmGDdkvi9JNyMoclJKMxgnphRy56xd8k2GvhuyXFqJiu0w86iu6XLlx
L+TW2mMpDk3l+nsQbGNYh8ltfdBjUZ9xiWCSDCoUj/colq2sh/dW8dkYdGtOiLnY
XgQoOIo/S7wtYUgcFRZdOJzOPrjYpqPRgu08wm6wEKR1NunJo006+hQiomQlNva/
4S9UyZBZuAUVeTsQj4/g7bduQuj0EJn1Dj0H6O9b50Z3im5KZa+zisydGWYK3Gfp
XK4O98BeFdCKMBkzRJ52qim74+8q4jBCSiYDX2Hg2xDKvZCPswmsJaNH+edB+Oqm
WOLZW66eQSXXJlizknWbPIDMxL2oZI/FHVa4naGby9E/2fNcHKbnwpuQ65yShCfw
EyWmr/cTXaRlRZ3NLV87MXejodQPuI971mQ+zKhrQDkLQaLhoZthu23K+JZ388Bi
IqgPol1AQsj8BTEkjJxPzv9tfcahaDDNq7pDFB+Skt90exiQq+vNps3cuoty+rub
HYZTfCfDZzW5EO+ua1E5e47sHhgJZ2bogqmV74t9k0GBXDQr1i4Z2gjwEW42+wq6
eMvkQW0STW3BXwVrhKdkDU1SQ/NW7JGDzRJrYuKW7+GVwC8U3f0EZSHVOGa8t6jN
T91p+IpQkb4kNLMZHwBt2rhqa+tMHWDhNqO07XRIC82sbsqIz1In9JienvXG7NhK
39wlhXDa3ewnp7sYw/n6SdhoXuj+hMalDgoYxNFlmRTnYQVNMhykWC68fGLu7ZOZ
iD28qU9mW68A0Dm/GdOygJMeH7tOPOJACyCVp9hZTDfKbv964w5z64mS6l56a0SR
HP2RFEAtQ9OwBp5DVt0ri5B644ofZ5BVc7dmI5UDAY6ntJu9VFdI26EmMskhmmP5
zqUSltV1shKaQQbfjUvI6llFRo7La+JgLF+d/mA5o0ju+v8Ww9eT2wkD654mZku/
9NlaZZCHJxfvlAbVOFeCoKVZSwmvvZlGdTCmd8PrC3k/uPVZrZICRvnX/qJsQmeM
HJA+WaMAIi7Nh5FxiN7ITz5vctydOCzSHVNiaU5rlwi4mq08OGv7Ht/n9q3hKNfN
Hq8esAMGs8C5/PW2HqEG311pcm+keDdI6XrZqWopX+K5qWi8K2db4r5M8nwu4672
AR7q/3QRhrvxFdrObSDgStPQHRktPJQXZLUFBz6gOIFokDcl4t4J6AMzYlow1pRw
hIPVDMWd1zicY3D5QqduK1NYQR99bMUJkbOBl7t8jBSRF5n96JOGR3faQ63MzEcn
etJI3brLVmE9jTew8AeyPBg3O9YOOwk6QeeYgoGWNLI5EoC00JAMO3MHToWcKqaB
TfR67Ht0R/gXlD1E9TNClZNajyxy+4UTAExxBFAQHVn0xJ7PobZ5oTUA70M7Ydzb
0ykmMLG9ncGmoqLjv4QlCCwApF5pjWqBtG1v7y7p3KRd9+fQmEhPGxj/ttBVcWGR
9/n+Qs8ftWUQQip7iTzt8TAtPJ+DBFCJp4BYMFUlQDHwik4tQ0UccI+0R25jQNEf
TKoarI7Y5KnpBB5IBJ3L84rjFkxkiMyr8ebZnTAwpFciahzpMT+kOLwkCv23Xosl
P+ZaoPT9NLcT5wqRjgcj/Mls/M5GeM1XCbqHa0FhqivAjIaS8HtN52CsdmeAe6PZ
W3W6tYQIB23f7qrHIJXhAN2kcKEii95hMx1f5g1SnU809h3yZr0qvAtfIRYJ7bea
RU2N3O85aI9UFeAnxLTXfJ6PN0mvpQNGq/dZwsd7DlqFyhEz+cYigShrXX9nfd/O
cH8nfSsrd3zfEDIcuI35xczI/WlBBwKWuE8kvIxafEcQu3IATiZf7ZKjjs4VCyiG
zDVlWG+AhVWsaVJ+I1IRCFMd/e8gUNNrVzdwH/AJUrjnZGFoQbIJKuu+jIYR9wL6
neU6sKjZoB3oQgln4j3LE53Tc2vvMm50pynUkRotBYpz6L84hClpy6WLEAn6rho6
ORXsQPuTgvh7gZqhHugPKA0z0nGazba1+Z4NeNwykJ6ZHif0zr1Y6AJseuByxOuD
sIpz8L8aSqxuXY4z9H6wa5khnRZTToZInKabvX6uHkjbXiu6MizVLSDMPiwlMM8T
XBrxIBpXpNoIV6bqDHWhydSeFGiRbiO8Pc4YSyxmm/XYpr2fikF0qd3SOnv1521f
zpllI7WWX3ixZebymu0YCSaztCztUk4aG4+QKxvIEf1PqsZIzdMDCPWMgH4mfLMy
OC9l/+djDg5VGECSv2vjlzswpr42otXLhHI5c/8X4KER/45U0w+3Hl58xaCRE465
3Ol5nbzcRSwWjPd8x27qlZTHeKeD5Zn0vTSZQxwHszATy3hH41npEbrVwHJNXTPR
tr2jCCGrslpj3ipfpIi030SMnD9LfwEtiyDU0aAb0VnePctVqnOR7awhclGB6sMW
Xj0HJQtw7nlStfMZ12wDj4RGe+fYLks7qVGlAIIMCesINVtsxJEkydbpBJpZsS9g
AvLQM4U/915YCiHUxORAFxrilxoDTNB9efT75j2xpiIyxIVXdaCMj70eDkQ7pfJI
YESPj3JP8y/QQ+ULolubuuHhihsQK0TN2oe9WZMC+0Pd9srDz+8cuABAYZeJL7AA
AKtQJ5K2iGm1DPbBikr4EZdYrXOL7dSNzTC2hnD3wXtS7eX2OyvPGZgFkgk/VCyy
6VkA/gal88ozgiPApBhYcF31s3KrkGoFW6HEuNe7cxsuZtsDFbnxbP8C04Pe5jSM
UUubo2Z/nxhdxg/MLZH33Uksyyr54db6yi4wE5uf/MoaCJaYICm5oY2VGS+mwl9+
sEYm2lShU4YQ4+VEnrWRSz/Vw13i5V/H2T3jBWMgXRYLzr4Ak+Lmv57zy36WfGFk
yDA3+aXw4OVF5SK1UTj/P1+OdO86QumV4sOfrqp6np5He7IF5dO0t4uwmaXxJcd9
3u3PmANRAt5xXFfuskc1trayIAMHFGnAr1x4RkiJJxJ//LIKvJgYHAO1FWGm6k90
/MCibkHn6nzgTvkJNekzQtF03HERh8FWBQnZODAPEMZkbvBDuB/r0sREGes3TJJm
5UOpcZeourgaSRqUnCh7ikxwGdDkbKVDrgmFV8mNPVWvX0vb/cbGaajfvTNDroHZ
rICSg9clpCluygMQ+q+SJYXBOj78lnXeC9XQprjpfqya64d3SS1Bf0UWAW4TspdE
G8NiB5r6MZ+uoKQkMN+O3LWhj/k4FVzRwAeNJK8dvvXIr6XhBonFnqJhy5ruo++z
FhagBMPIZL5o7yaF0efBD45GtGp6pJP5rV0EYAnwQ2XA2JfGLvmVQEOHyYqZER2p
P9r2gQ7q0Tg68FNPdKmMPYleJye3UT2+VbRat5EkTuDCUqZb0rz0S5WSDVkv1g6u
jYy2NGJ2ty1ScnagE80uaoSLi8a0vjIFt+Vjzi/alKqyFx4WpE5mD0IFQkERpsuI
YQ+mafoVgO3vwsz84Oq0ElqZB/2L8Ic/dgHi0Sq5lCnoELcev7c139ecIjzi3tlT
Pl87bMKBNFY5bEy9UBKc2Q4fmfcWTgKnyLzcsI9a8n/I5YbpE726JgN4Xk7LZuQ9
Ycapim7qMu7xTtTq0zk3hZaLKh0cl9287Eb0/bTdXbgDlA66wrxJhYW0y/Aawbmy
b+AlEg4x2xSrvW4BX7B64l+GnCETE/4kq6u3SgUsKSdfFEWlmunFy2AWfFspzknR
IGF1b4Rg9J8BGjjp1HRu4EKyJuw5hscKvYZCOtTnAZebWtpOu3kbD6OS6IwtSaml
WW7uQS+pUOEby+hjO+g5FpEAPW0vEfvVHt5EtOABwSN0lT2FWyA/Axy2UwWeSp6r
5034Y0EotwB+83b8Zel6fGxLOd9rqfJEk9BV6mUzUiQ/E3SneCUO5uZYML2gzL3Q
HtejEUciCdhVo5MI3LUHWZZhnfy0DqTrjdT4445RaL50caYQhduK2JFaC78wVkSd
Mw3dkV6TJzy5zdgoFbpWTpQ2Q8yDNS4R1nTJd0qXeQFD/tGo71pU5D5qMV1QLgCv
T0qGVxUxfcz42xIh9Vpeg7ts3tqiwXfiZhxLGjHQJewKViZoLCsj0pyHSCqlqKFW
R9lbSCU1sty24BaRvKNk4oACtdzRfRMlQ4l0BXjRqqR6pXI8HIOoFaq+zBv4Z1Ve
g0141bpiLhXqqWmfsdo7QAMYJ0/qvIOoUCszqCV/wS5rSZ3qB6bt/h6an6+IkjNb
MZanAb++E4L90HmcH/7ubEOL4FaJ1zH5TB4ylsfrWBrS+n2sAWzQJjxUC9uhABVY
Pw4wHGSbpQsxZsKuT99DM0t0CZsMNaiItw8v138IkosH6NYUnd95Cktq1W8UOt8s
TkxqUM1cDQCUGTdz/4ogx5tZyt6V83FFonbfl/1gy59LCy7qqJJzNEb1QKvOWcyg
GnNpMB8WmoPuvQz+YR4AKg40dtcOu9YBMhrN0RnBO79s8GsQslbBchU5mrG+t0Aq
UXfFWeRiLycdH0JzNypWZ5wL3zLxhs0HyYJQ8H8gOC1MIyobudeB0Kii6fY3VXqC
YwXzOzaneyxDwRXZBhQ/MyjHARCOK+RgYWU5Xu+fjkIm7gyzgRSBtGTj3UOyPKqL
0gdghg/1M+0XTK2FKbr7v9RSJcvIN6THfPsGMRk40NsCneNICIVntWITIJ/5kUA6
us+eeuCFBzB4mL5hHRsU5IqDDcTjDrz6wVfjWs2UMWz5xom50V30ok07ibbp0yiM
PUDOwVfo7L6Prkhq2QmW/0egqGwwICgE0D2smm35YKjXCjdyTEzQl6OTl6lbVTzp
xMIDc12fpI4Mqz+fPWNCxfjqQ6f/4sb8uRUQEBlrH07loT/dclGapAxvwSwcoxY3
L8Vouf1p5U2xbys0d4W57n2mznycJhsWrql/AgWWK4L2K5jrgH7SMcUoMazy5NwD
nl5F3WNMGDCIfn/zzKz089RaPh4CNyhJqp0nscEO0OIt7AYqjuPxKbYKD3z8JJjW
CRmPecIewgbQShnPZ58UR0+7jkuFlA5/7m4STVDbEO7ypi1xtFTv6vcrrBB+QpiU
JQGQQgwVFNBBDzljZFPlEYRP+B034SXLhsuG5CNVRhZTQc1opEqDPHPEEEXC+yIF
scbdkNTMI6UBN2CK0kRsvm7MvzNjmzgYqOWfskJFCUpBEv1hS4ryqPeiZgLDJMOL
KhFrrVJKIU9cHc2UyanGMNxxG4QyeA9MtYaxz4t+4rGkIlqjf/ybbl48CdHo09Vk
kk1p8pttqejXI96CjxDm7frGHx6LK8WHnWMKdygQCM9zjRiR8HkgTK/t8CLR4NhR
ZKC+7IBPa6lQqe2ycSbNtnMdwKMytjzgTxagtkwQaGa+R0KON9bDOanYqomOMFWv
x9A7a2bXSFtgBGYW206cQYBWkvl2iTnLSpEdWnEzkRzZ0EsXGGaURw7ysiNHKs/n
OW3N80GUyWePbt26T3+kdC4b4hFVn0nw88OIfdMyEw8S2wRpFyDfPnoQ/aUWEvNE
+vYoLC0hYvqEVuO4mcVjOydwnjF6qg6ep6t2f0/PAkQAJnR08wU/7InKpZrOEmfY
hWHcDR969ZaU2YCcd43bxOKhlS9YoebbVYyRb1FSpHkSYrZ5H4Lh7/ES/kfSzeMl
SH0JPln2cGdKfZ4LQbpDk2h9b5yfcMXyGPMc/rYr6GyyWn5tWithlB9rBoM5wDob
UYTGdDgj6x60EcWa+rIjW3rAogBjR8oAJUViYF95eqCTyPOHv+R1VJvAWVMMQs7N
+Nu7BrfauDt1C+oM2d+tTQQgtJT3or6I01CFDMyJe77fFr0M5TFXZTbt4WBW/mnx
AFKmpPaY9c4D8BEMIsOQac/QvKR2Hy9qNUWHASxtHCZmgb/QU8rFORgBgnOH7agv
Yc1v5B39w1bmGd71hauNIA/2/Lj5MamaTXytCRbqRdSgPvbVx2HQc0u+KtPPRpTE
W1t+XOqpEHtyrnp9igQZE3zWW1bMKAQHiba6F+EJeQfZGlO/zQ4ddrRvX4UFiXW5
wQBLb/Mj/2HNk/finE7D+15NQ4nHw9HT4idGu6Kam++P9vAYeOg693EZFmLQAPQY
h+AYimoktBHngZ4e6OT86BnFFr9PonqqoVyqOoJKRyDRyOjojn1/lbdw1uQENQyD
Yv2svCGJg0r1RPkYfj1Rbs8HRNF5gO9PHEayFBRiwGA9EOSIV8J/7TKt/evIwRLN
N44KkOnDEW27IdL+Vf0fVA2IvB7uVba1E2quua1k/66r1EvlUFL+sN7W4HRqlMR/
4sKWKFLnqvHwYN+K1azu6gM5bTdJ+UcuVzo0x9AxJUbQhvs0GEYAihzvJ17kCOVj
GqMP8iVMQ2O+la7DnydJJrMyY7OWVRgPTKaTNKdvxP4kOpYNQqczuEj2vaHKjFkt
L/FtYHs5fMbLhsGPlMprU9gq/m+jBtsvjVncsvzcHVJ1+OVczPBgPr1yoY47eT72
Ssrfzlvbp8bUaR/MUro7O1kM0+6B89YiwXBx7hA3D2x4MKWf8FS4lg3UG9XEkcCM
isrcvOyHmPJeaAaZlUBFsDrWSVwYcendQ/SD0kw31c+JzJvd/Mp4XIFIKmYi+g9A
1XWnTy8HnxmbYjKDaDNDdx2gXtRYKtuGm9dnQZ09bLhXLVNQwMnoGoeeTUJ/F+Zh
AEYz0cBm6YnUVECKcDdPvl+4SR7X4lTGQjPtpBSWFh7mZiX+DWcRTgAa6ksGcE1b
gpKwGe/bzbtLlscMYb3OnXZOXLZKC5ULLai8g5jHj7haaBvadFyczs2XUibjEsA9
cYu5JR2l9ivO1u3j4NR0i1mxTDjacazN6bYBFTjyWLdXn4zDgoVIpJOstxeWNTIU
ZyT7wekigOM7rVC1WcTDBJyExWNt0riI+qKq7wqsLDc8FPt6Cv1OtnPqwilGKeL5
qKvXaN622uzPjEIQwIui7z+Twb2mlWS2H81jJmRiHnynMQ9GcCX9+yBD1O5UiAVo
+xBbBCDFtMOxAbKEebjIAbI9GTYzIYgQSaU4iOWvu/kPg54qDcXnhihn3wv8V9QR
Q9pDMYyCMk/NZLiEG6wYkgKvPLyX3SlMumbnu4ufpa5r06CRy4qs/wF6+BX3vZ0e
eiSdFz+MVQBSR32Hb/wctDhX7pMDxey0Z0ceBfz/+Mwfunvo2bGWG1jDOh1AG5tP
uba8LDaPYbMpdSTXQL63+Bkr/1NAF6IcV8gcIKwBS6bN1vEzHcyzHsCccjXCGHzV
wpg3pe5XGRFiWsH9IG1SsgF+1Zpj3+v2fOmjiLNEm9j7uSp25CvCyoFvJtYeISOo
yiYxUwJITYKz3x+xivyL0Rw4yR5xZjhNuPuxkRAdLHaAntO4jn/Shau/HGuQ67DB
U3QI5eHhmaKBlfDP/rtpAwNRQhUo+wCX2VkzTeZ9/a/bICeMx0okFG5MPeGNeIjW
OWPMC4IGLR2mpZPnjzB5jJijeeEQ+UKUKzDlY85/hG3EebfMN+eRBaPucb2XkqNT
AYV9uPXl4dtuk33WPYc3WvVcnWVQYuBF3pk2zqCLQYoVL/wHtNQEYdTRFHYbGcmf
IAXpNlXUatcff43wJ0sPqsDIvdA0OGI5k+fb8MLPhll2wxubXWcxaUe2nA/0MHTD
Bi9vmFiaH8gM8ZE5QFYAUk96AS71wLeKVdx2oQEoQDI5rCWekPDzzATeOR37+p5K
zXCe5Jvt7x0ORjLKtg1JxCN2IBvDz6m8d9A7jh8PAtUyah2CZzwbrZ80iyEcdQb7
E6m+Eb9xZ1HuK9TfGUzI2yCoj01lfGDng/HgQRIZwJVMDGmILPhmWuBB2YY81AEa
WSGegvKmeglnTLHpnVrIEwdP5LskCMovkAbBrnzI6mAHLILaRAguQZ7jsY1lQIbO
R10SX8C++NQRWAJqOxc6q9mfYBFtHAnpGZKoaaupEduD7QalVtcYYJwKdFQCksPn
DA7t3xRMIs0eP7Q+tNKeD1xfhmnGn6TWAQZhXv2lvTYBw5B54nk1Xw+/f5fVbIRG
pSWTUWmfxP863JJQV3OgHqrE6TFc6+ws5o7x8Pv2ZjXgkL2i2kb2flF2qPQDyzJh
BslF5Tz2Wf2PX2+z+iKOtosyLgDNTM2bnKMRDHCb8jXtKHNU8lDLci7Rxc4ABiy/
EZGPrgS8vXacTjGWUx+qK7/I+4p1fgjWmLWpZHZxHozlCEjdoov0qzUblRl7tk2E
8aWDmDvV0+HTvs32H2UAb5ewJ7dOsw74WCJBJWudr4R6giUR/82UqgeUKTmkde1m
Mr4WYmbdmumnoJjNHVKzI1zztxguN8yf0L4ckY5yhScMhoUr6M6g9O7UFyZom6nC
0dHEwuRUGrI8p7qQgWrGgFnZCDbg+nbACUTrG2Dw4RBLnRPSWKepiYIDZuL0lwW0
6EqY4OloxYEBQ1JTauM6RnRdl6oFD4p1vJwPc5Kk8N5oiChmfX5kPi1GwIkp+Rbz
4jhZ20xVeNTxOOdRp4uUxejZsCNNx7kMAH8w+d6RdfRymdFjmDcRE/YV8KDvTpqU
cBvPIkOtUhzPkPYt+L6gGfd6cLJjw9KF9sGx4s+AHY/POF5rBgh7drIyFF564rmf
HaJmjHmIwcvGsuwJ1A2sJksYaIy/RqODNuDgVmOQef+yaH5Ferz9blEKiRjh3sio
yvqtMKv2AeWmVGq8t2zqfFZxhHREx0J12HpTqxdC1Nn5D19dZw5d8d1RwwTr5suT
Q2TFsc3YiBTm0b6T8HfhF90bHjWsTTuaih5eSeFkIQ4emTINevxVwdB1VSpT3hOf
rFUIrjGo6De1mLKoLXVASd5in+X+XHKvy6oplUMAeWTe034l5OEBCCd336oyUObT
dHQTsvLs72/6RGpERBmZTm/sWIgwuiqm0yguf8b4miejuPKKq7QveD3VpUE1YKGy
rOjWHjrxwAtIjoLO1BObnqzOCYU7RGVL39pXdsZIs0ZUOH+EERt7aa6IjI+UAdZ0
OdhU3o54psVSCWoZHgDNYaaYehDKw9tcIkyzhG9wDb3volznboydlKpSn6r2N6HV
CAB+CJ/ZNAyNJC90753JIkVl5tENwZopZ4Q0kKmMWatTJaTz4U0Ys4BD0YjAf2z/
QfUvcUVBZtu6NVtrawC68/BJtBz167bvd8sd9vL5v+YSgJ1/MmbPtJW9GLIQOAie
arCCtxfNq//tUV8bGAAfNwf04p+H8LhDWJP2VbCJ4wxxwiG/DCa09itmMAyM6nOi
rTynKOFivULtI4Wwk+5wx7SlQVhzlsy8NSoUL+XMnU84XkMl5t6urInIU6DOcUW8
BeTnZtVfSJTGl/L8KLwWiXAGJOgs1HlSpFEgKs2tu5MBsFazifyTgo3CERoq/bEb
eqK4t1Meo00Tc3YLmDeckqumuQ6D+uoEWgzQVhMD0nun13A2behPLZs2tSoqvVP9
tw93cY0Djm7Rf7wlVsYfIyZzCYF/UruH6WtU0EJVJ+uJCbc6VAvj/XGUYV42eFp+
oVXeluQijuoiFdgW8dvi8DJZibwHmZdaPnyVm8s/LkAcZNyaZH6e4OsgPrSWLzE+
Wn+Tjz86cHyKZTHIPw72s+bPOuqsY8sCUVid0lPdQfXMEXhIgI8ISlLD6hnD9WZf
kdoPLWYiC5g58Te1ej9BEh4z6HXpAnYcYY3Hz0cjOnRr7jAvdX8uPgX7xvLU0HcC
/cLHMqemDp0TEix701uFlMeInWsc3O3rm7xxxZ2GqgVIAAJxVqTFnE5LfWbrd9Xp
QOFCz1C4JW4QAR72DWWbRw7CGBXfoDYbxyUnuLIavtxmpe+iCf9tkQ8FJL8m8yMS
I1zMj+uHIrj+PTmRcXZC9eenokq/TXQvXOgPT5c7S2kzWHGfmg8GgygO89PnQKOG
ScX0ZN8/rrbnCgK+H2+wfodHiPEl3zVRsrNciADgQP9fqBSNuRyguvjAHNnlrhID
Sv3J189y66XeFk7VFRj5mWIvWIDwqS9hwtg5oDVZtak2WKvvhd/kiB1NaFxKZGvc
4lri5GcJLNfw+99bsSMCWzjcrjQNiFlg5/Ru5Lf/NPUuHd285HOecnrFlijaUHwO
H4ny8yoLM4FelaUeOjfn64Ap9I5QIAV7ojBjxGWlSRtrQputuAxk9K7YeRy8++o4
pbBmjSmOMnF2gIraLFt8ylo7huV3HTPZjlESzDUwoGR01SsyZ+ED6sbQkC7/8zOy
3IkhqiKQiFsSik0W4b0Y6Zg1AGcrdCWdmtDQno9g/NuEV6oMeCuQ5a/knti84aUI
6L3Hiax4YV1snYilnvvSqeRcE1RFlRILjkhMKWwK9kgsiD/NeqeaMwHfgSMvybLS
hDESKZfanz9br9uWpgyg34xKA+2wgoSWt+zk2hLC53GMPHCvP1qFgkv6fup63htS
jdS4RStNt/oLDtYTFRcGez6KDBZj7GLuG5BHyQilzECfVdPgLTlkKGnAyY8HR/uc
DiYbc5eFX0AYwk/H+yYu0wS/DhE7ZwZ1z66LjXxaa39/Llo7S/vMr2mM6JDzFleE
sZlgJyCcGR/7B71+vvl8HE5A5C8iwO1PY8Ja12LVRb5Qt17KSkT4IxJ8AE26JmTy
BcO71tCTqx40x8isyIn7KG+3k4p9VYbQfKtuV8ackpdNGPQCVtTLn09Y7E9JH91W
KERRw97ZShnGOemjeNpLH1zTaPJkY9mBA0laODKcifsEaySZkcraYpyaPOvSHYsr
HplgBRsiAoB3a8ve8ty/UyemneXszLxP+MJDqAqo5UuJk1Dvr0P+/Kqavb6ZyV67
jBYsYP7PP4WaReYsoEZz1iyogBfD/Od4yuD+sk2yQgNMtl+VDb8+NY60jaQ0gWk/
+IY8rRsHuQ7owDqsCVZY+RCRAx2q8a8PD7vpxmOwQs74uWhgfCqwLIut3LdtDXoa
GyzbWqppoU0KoKYswCcjH7WOzmy/WwnjRZlTYF2+FdPQva+3VfBj55/NCV1UQ1Ce
0WzXUdJ9JreLC7uq/0e1gl8aTryzbNwxcGtffHxOmmixUna4MnF3sUXsON8vZjKo
4yQXJJjTvaQEhsxv6egXXKXbbz779s5dGY0j7shThl6ExBEmgx+pddSfwE+TAVgy
8uoekuyra6AzegItROY360iYLgFRldyZ3t3c6r261VHY0VlMTvLrrO3bmnjv7B+3
9fwsdd6OsdBqElAbTF5wby8PscXtQZSl6/+/CBgbo3QSiKlQjEzyhA9S6L7WnYf6
4dJttlt9xtz9x9UStfgMyMIzzMFpdQq3IuKP0Fjkg3/pbpvkRV4BZAyVbtM6J2fc
bkjlrh/Xm1PfUtn7dUXBji1GAdnWcJjkDDnJj+1rumJlGap/9/MQCgK2/PMWPZ1g
YCR8atY6TBRXd2IsKA5kUVlxSIeby1PA4LBau55vcWGCwj6pSz8mjbBtf6C/vcCW
VaGat/hJCcXGhKLkH7k1xxMHMuzHAtk6XytqwKbNFbbuz4coFyxw2ATdd6cwrYHm
hZ+cqXY9FyDKG9fYh4xZ8w3VaAR3mMtVceTNFrji7TNUxxDjKG6rWJgC7mV378iR
S4/SUcMAJhS3FdkIeQ1P8dHdw+bw07uPekJEODyfFGCzzVZGgaPy74Px685LZ0ZF
bm7s2tBADlWbSKOuGdjPKM1w+E5WxK+5Pa79w5dy1l40sPTsRTXK0mZJyDJFC4bE
M5rc0saDhgseAk00vJb0cEHyFyQHnFEBqswBln7QSBO+wziCY8ZZFyZQBTYvCCx8
u3kmPEKfc9w4UXE5w9V3Cmf7QZHssr1s1QqagtpDfHqFLs2oMPzHmlebmjuqnVKr
sSLJ744m0pPYHoZDtiDDFHETK6rHQqlI3qXN2DR/WEVSgNEwVzHOu5qQjxLoSO0Q
i/8FGKR8kLUtTygSrdifHf98Cl+8fwPPgQZUBSgbAfaTyVud5AUz2cc2Uz7ni1cX
fl2YaGs1Ni8gIaXYC2e2bSXebWjkORqvZbWfa7ZFY9eaBGgWDRsH2/yVfFBR8Juo
/iESI3OaDZxw5Yj1caB1tOkVqCQ+oCJBV67cOR72vclKb4fIdeqIGqglyPDUZHSY
ycH5l0bQD9Dmo17X47hhTf1rHLajUTBrjU7p2BK5qH5f0aOlGHrvSkdxwZr4funv
zaPJNCvAb/X94VLAaFyqPaaD/3YdsH60a9mSREE2kMzr0tqmPQgNYMnSv7w4OpqD
Q4rcqpFs8xMvykax5zglLCrX+wNaoNe4Hn7VoJTDTjLEdNJ+RQ6J5hM786FtrHpW
OkLiPdfvZtKOZtxcU5BmLEG6HMHILcgGVpxUqJRVO8MKXYx9+QfvT99IwUg8qEuv
hMUDE1xzz3tMs+DuKQEwb1PPyiGd93XmD2t6MhaAV2aFxakMAYbynJ1uphPri+Ri
S7M+pDQd7O1bzTMPJJFLpKU0G8JW0tSF/sORe3qtuJpmsie53eP5Qa032z0QKesy
yF899SvoojGhW/swtCoaFyb4JG1HdxfCZRlHk5jHSHW2W1Kdg4iaWP1B8vdQjscP
spWHaxMGePkaGwoEk4DmXW5x6Ls16pjarSsVZIUwilwAOO/71pVthKo4UQitgqhi
5V1426yqorBjj7MYZemusJlycd0taOgutEC2Q2i7YeTixz89GKaIpn/YtfjNLh6Z
/rVxDsWdLhq9rcoMexxxBJMlTqp8xi5oGE+4SzR35lHuj6FADccuMVe2munNpsBK
zMWAeSAXTViWbFlw9LycYOX5WpoUCCxbzFv/brxMdGEM60rdzZBmjV7p0BkybtMP
vidUf1anxJwEniEVeiQx45ekutwkuXypl6NaFNOofI3pL177hlPeVoqHh7y8HKfn
cXF/Q8wi/hESX0F9M368bVaw//FlAi6hUfJ5HcqsADJCXpnTNYerT/i5isSwMfst
enK9sNv2iJSRaQozcIDi+DjtK5Td/xQRvwNYu6KuFVxaNFB0iCJDMY7kXR3lnsxZ
0cq9iISp+CHyUFfalc/jL193/ttw+OhRkJls0EaKx285BNxUisDO5jzGTNuTZREe
V5Vjo6vUbep38ImB7WTQRzrE/Lrb8IpbUxrFq/FBi7+uqPoetbL8UI758xuN7f/9
cgR8WxV5yHZNuFnzE7lXdY+o0ThKykZY0V1vFuVoiCP9yS/eYO5wYsnsWrU3pKr5
TaYwabSyXgh8fA4ca+SC5DvMMDKS9QyCTth3WR/Fx0Dqrqvup4Aim//82wYWNr6+
G/O67+D1Hfg46G9OvKSVY1n/EmIftnX9qapbXAOo6W98Pf8Am9+FqMcACnWSRWiY
ZhaKDLQ2Eu3DgSwHeIj1q8wrEIoRG6pZU82QvrGdUwEW9lkrZPCap+sRjTpGSxGF
wEpgolZO2hKWBD7VMxmeqeLWUPCBaCm6sKYLS/XeleYcn2Um699JmmoqSLlacXnG
z7CMSoSt3TXRbRclbsH1r0EQmxDofouu1+si2G1pBFjk5IhqX3lhvwvs2rqkGSuv
n3L+1oX3X7tPS+NfRvvxpikqWO+Tgz3OqU2fxb4QbKnNFKlhjwGpctNReLbzSCpW
3GGjF0xOFDqmDCF5DVxFOsGSCvOWS9+p8wrw9v2FBOP9s0+E3aegJ8A4fvJkv+PI
JKAnwbvL1GRI6U5iiUA9AyJCcrLT0ISqWk0HKxIiGdXy/2R7iaDLlggKecSYrkdA
CaKlwqPU0QwcXc/cpaZWqOGJMQjp+7gRpRL/fTI/7gHCYMTjngQJGsJf94arXUVY
NraEtpFWDc3mSI4V2y6uWDLKgWukbtJGP9YuyGllGVFUcGe1IivHamvGqLlJagps
gGgU5l4ed1JyfhLFG+oids9PkO/S/uzudaaCZUDUIaeUVg23gHB0AkDknu/4fUXr
gtp0SVNA2U10Ta0G7+ZOAuh5zreZDR0zLKWoUULzAA6sPpN4xfiRNBqpDZsUa8Xk
DsTmmQv2YKxNFYqUy5tWO+ejy1liPdej6DPOu+Em9vHa529fyXZRudiDefOVv0KY
oX/JOkVZqP/dwW5SdXoPpyyM3NMnZ57CRzzoE3jPYdR6zlVpEDRcF9QrHSf5ckd1
uNzut/ehkdlIZZlTf9p9iMPrK/lj8Q97MKz7+eP5vb5Z/77aemdO96013InP6oZB
HqgiJRX3kye9yHWa5oZrQAReMxtYm5SDUzPkl8F9O7A7f/VxLkQzQcT69H2t/rtV
fBprivrPLODO+dZb2Df8+JORqYjJdfOIs9M+EE4SHeImxBj/6gVk6qFmb2PJoW5P
7eJjtzT/LxX00xFYQR4c7QzvesoP1cEhnhXKpZLqxieomaHvfhk+sx9UX3Kl66nG
OGXso81Wsk898HfXWn5qLmcNdDeWfpSTaQRyPvGEl6JbChKu5StPlQJCulnogaSo
ye2MEisV51ouj6RocU6qPv0hWUQ2Bs/1NaeNh8fy11y1q68wHDD7R+N+xkPg5F1A
cwYP7KYn9a6ihXU4wzulF3ggTl+lbdbLFta/F8bXeunE1YWpqBnSHGQCP7iM/U7l
w+aufNrFOKmkJ5DBHP5EhlCKtmKSgZ27VuoN6x93ldXbwv0jqsVEk42R9KM3+Bfj
NMO6ePNm+7usPhv3F0FgJUvNBPEV81huB+Hcm92TB+rV0Yq6tibmFSbkGhh22xHs
KfevOZsqmWybPCnstU/0mTntW7n6qObSlwj9nXpM9MwKfIBXcuZpVsyWcFK6t9zM
34FFMFA6/J0t0KKsnDQNYImNwKJW3qoQmS3B47tVo0UK/hcvkM20lxMZcOMdmRpv
/UC+fUqDjRrBXE+Z8YPQ3iT7KdEClZRD+ldb2AqIeV8PsQjd5rj4pOvPwxHNdEjv
maj7YDaXKML3uW9qtm6lUD/xTEfAKZXKbKNiPaavMeWSErKd1a+A3+N4NYxNOxXN
2h1Qc5Y2zjTLtozJuR4XQqlMiuqr29kf17FEA1N3yVTkARGkBFYqxrUyH/IFCliD
Z0z0+rsDZd0KwhWsw56KBwM90K2egRe2tLKWdlTNQRoa5q8HffzPGhneY9y6ReLE
jZEYmHMaP6uMBX94IhumYuHLtqyULpgO4O/rxhrrJqYP2MEFJqZGwC7UNzF0qW5A
KjTqAL+dN/WCl5Yl2ZODdjbDPJU668KBZHGZt+wk/J6DUAusWU9YFH8ROvdOHg4V
8AfbvF1DrHhv+8bSv3OF/KnRMfpqEU0hzqqr05S374tnbq1rpuDr0jg97jcLYxUR
vuVwkTYPZ63/wWr2o6GxniUvAtitupXOc1WTEUkGIBlhd6a/IFeO222rKd4eFzSz
VqzuFJjIUXGK2koPUZGC/ahQPnToykTo1N30xddLx+9cQAv4Rejcs3VrRnxdJTqJ
qN/QC8AzhTz7WkFvWsKvLuGPsvkQ80ZonM4htdi7+Nwga0uHFEwIqTtbaqtBelzr
wAdOIEkBP4FpnJmM/8SO/YGKekilwQZ85xt37/WmCgRI5uBU3OeTCfOawUaAi+MA
urbSKCvOglaMR8Y9EJ7tk/MvJl8C9qbWH48tUepHIj+QHFis5yjZg60s0nRcP8pO
RxlARHr0rsYvSYq6M8oQel0742T7usFl/XB5o1uicvLPNcu9DqQoRxiJ7AWMNsAA
gip1jwC7KL/r/RqdU8s60T9TFiUkwZ6MUx2p5DkPRpCjbQDCqlWpgsEGQQtTdg1V
JNzb3/YfZpBNLYt8LnSr5aAFJ+uBXfKwfnmM5bVDe+6x0ZYJwWg/+tjuYxj9LDGo
fwbrXic++e0i1VCFhuCEqcbUtJNielJpu6+IpVF/ID95d+CEXwCr4dgOwMYFxMPh
zXjs3EUVIoTSu3Ev/SFOcjIBADl7Y4ZsxT2wYgAF6FIPbowcJ9y04mLb3kKVqoDb
oTKnsQwqqfIJYw2vezuo/guhv7l7a7Xj/5RrK1icn860qBHUz935C66K2EypxXi6
xYri35baHfxD/nLoohK3ipjuWtofvz9ARbjx++W+63IdWz7SRXoSBPjAD9e1KXWI
YOhL4fH1yDSSAqNcNy7EAj50z+oFr0bXyNgWJ6Feo+vfQtBQ4Q5W1g80ZGKk+IRo
kKw1IajKdgcToOh2UmcziZtFMp9PzjlI8Pncz8VvJwgSPyJZJYpqQqASVeKj72k1
j1uGRfu+JX7XipNRJ4hCdfl6Zf46XS6DieM2CKNF0zjTpDj3tUqgqc9+PHAhKKom
wC+hdjHUa9TGECQ0nJ3IGbbJdO0GRTvYooQDpJltXFMVdlsb8yz5Sz7ZbVs2ETST
KHaq+8bYtoeMRXPc3XJnQpp1un+qKZ+BfcGqSogwEGEvr6O+CgWoBPW3m0O0yUER
WxKFseAlYHhNSP3+uRSkaud0icF2XhJpV40iSdDpzdibMEcU+Pp4VcW7iHHxQkPY
88ht6x3MMDMkr4Iq+JvLxGr6yslhaNSZcaslNX0GEvVpopfohKm5CLA986ElO235
h8l9ljqHAc8kLlnqX9rTKQeVsJaIonf9A1kWkLocW06/tCuQrLkfKYfRC4E5lFNM
SRhyZK+TT3ku5Hx296MVabu1k9v0kM7a+g0xhfAaoUeBNqsQp0cYr3Wp/Oosbhaj
kWfoBzXHs/V4DPesG3/EzyeJIIyPaEoc16h1HuDBSY31oWhxhL7AZlqLOYnDII1T
65wTzoSZG9WVINWF3uOdzJBT71KFHygptotelZjynxczbye5ZBDp3YBBC6+78j/J
X45CgjH1BjH/iPgxGTNKQyldJrF9yT85oHNzf+TShKjgbaMOpWF2vD0i5Do+j1j0
bnu0dtNZBYJD1mULaGN1HWpKAkCWImj0m01enH0d09bG5jESpxiFP7TZuDB1Xflk
A/Sq0xBYPrPdgPtZGOka+5RAGx//rC/RV7S7zubm+a7lsj0JKPyPa+xm4b+dEmyt
OTR6PLLzioXMFipjpiEyNYvztjhNX8LWHX8u/v2RmiCU/oUoaX1/UvJw3PvTOcJs
0eDqUfuOxgy0ReaPdDmtttpdAW6A7QTA/hv6t2FQXpj35Iy02in3f9a1vhaIo+Wq
aSTqAi6CHRmRiR3o90usE+dp+DWclpUmvpu0wc2XvmjvvOEk49LevAISe43VlemM
lQVNa9uYfougk2ONpzgkXndpGAmw47RbcEp2GK9tK9TVOcjYsGdWomGGocj0YTrc
j1aDcr3filHPAv3ZtCeR9wR9YMde5fsK5W7zqYpoLs/tvipjLcgpJNEAyrPfd0lZ
dUQGCVsGRK9mO9FWFL2J3iKJ8Crp12fTP71dcHbocGpA8xCcl4JceOLf1hLoZR1X
6Q0vPWTLtfQE2IsY/sBg4Jjyj90HszIjJtlex9VVzKlcX4cFr3cyWY/v2e5hfgF5
EWu4ZbTlRdkopyYEkGyKCGxDajbv2aTXhZFVnVe8reUP+FaMfTs8tKvh38ioBNjC
4drxspWGl6OXSW/f4nkwBltN6TMnaqjGLTScJ46h+oRiugC4VnoI+17XMyGCfK2G
+SDbk2CS9r8APER9rh5ijhN/BhBMSnJUcMqMnmYOaAPQsljse1kUqUT2NXjQCxkR
NpRfXUkJTNu9NXaB939BggTl0ehrxB23Zr3aYN6ocM1icewnTh4DFYYuA2/B9rGL
Y/E5WUjDizrN7ES0KMjVTZLzlUTJBoHo3tBmm7YA20EZxqUw7Wf9ZOc2HisSSIRU
M2mmL5I7hajDR6BPHNbyGrHzVuBp0vErW1y+hRQkU1GN+a4f+2SEC3vECPiPvQt/
LwPm40zhNQAANt08Tg5E7EDzYvDfg1E5d8sNXEp165IXxUa77Bkq+iq6rdOOAeZa
0/Q+2fP/U4C1dPEfF2ShmK6SwogPy1R2PzCbFdEIlWTUM0020ME5SGQGlMTDVc+Z
Zu8UIF6d2xiJFUKHGHiSOuGuqk0TnIMq8d0VgdR/MOe+fStRF+TmuoyKAJWkkMRw
3XvRCqHpJ6RG8+RbFCNcLBjIUt4sk6s72GWIhYb69CCPqlrFTeoFEpYim5UQbCnn
jTvxjguRnTrNdcZ8Z6L6jKK7N73smcv58DrPEGOL9dQnxKyFGPqITnM3e/pUOEmT
/FtnZIqo/0C3mOeQunKRkx4JVbl7396tJwLcxQDQ1cUYOaNL1U8CmYZTCVFNOfki
SV69fEoYZ2FNZLcMdc/PI+A6Mc5B11Cbb2AbgykgQhbFd12AaKAYnt+cWmS4HBEJ
5BRzo3aAbIkna89+5eblQZlfQCgXl9febCsET8K9FuJzeobsaMtJftdtsgXSOI8X
KFISRRRnr2+tTmILIfVFBgCRKcxGWqABj7WkwolBNKE7PWKZrcNIFr6Mt0TFHymt
hZRo3F9Rs9U5fDxAIxp5K+E7uRgAOgTX47bGRwBbci8HT1SDvHNzvg6DDU/N2YCc
3zrVOvLTQPiFd47cv4fMKTHsIcPI8FVCSHTFLXqJ6f6qG4+qgwS51D0ldkM09dC1
ryv1o27QlkzoPKBvLItjTKTCQWW67QVRHu6VBu3a7DUqGCgYmc68n5+0jJu6Mhzu
dcmwxxWyxBTQeQOzry6a5HIQ1loyWAvg69KZxY/9SGMthMhJefSNMnO3Z1VfuPNe
dme0VEh0FP6YpoB4AZlc/9cz/POQSBI6mXHMXE0KsOjxKZpW9A0KcMrwKhNgbWJD
II5yqRdRcwY7mtXCqsPLyT28mREUAn1JAHfmZBNaqKMzy8Of+6R3fLulfjjQsaPW
hE3Ax9+otxzCp46nrmPQ/Am9/GXm/f1rnUUTSOnfbE91W9GBCXYu/f6nIpQWjryo
oPC6NuTDGmZwhazGXRS2GJvhkKnUq2UNDpX08mX9o/DbcWxUeUCvo+YDSJALcW/i
pzs83vb+q5EgyRHsIEkK9zSPG8xqbnHQcMgPpAtP952Z5nkx6BRLj/Ya8m4vvpHw
GUUdvW3Pgieh9FdRKaIYAivaoevfhaAErramYMeUtx2UUF5a0kow79dt+R3srlEi
A+FniBPSVTAF6kpXyuKSoTZqt+lnl1u+ZBUD86pssBGFJi+SvU4wk1BpaOX1M5Zb
n7zRU/qJ3BBIAiUAW1Vswbe0CFkcL61v/rWdC0q9S2ArF2p9iKEnn7aZWoE+vq/K
dfGO2+LFbknUX2zjCZpOQZzmdIYLQy7ruDtYd8Vn1eePrPkTLxbxmIhbIgFjlrIs
w+fkRgfvLZxOpRlXzrxZAQIzPscsQMoZbYbx4Ohd0xjqtLtgUayBBmcPslo39laS
PNjA5jwgO8uucR+V37lPCtjTANG/D7p/bECZgEFpe0IK/YbSR5sLrUT+ixMPSWVj
dpIZ/kSWMh8byj4RHMy2iYzlbRnahYbX5UOmdVhhm5LHmeiqw/MGm57cpMn3htxe
tlcRFiCHbq4bTGUnqkBWvsiBEVIV2Ym3njIicQU7Ijb0uXQ72qot416L8qJmFYwQ
HCMu3hv6kb8mziEMEBlzHMJHU9i1V6K4ms29pHuUixWSQlegxfmP0vILwaT6/bSU
nh931kHwHXkOWn9H5gLFsD1dHyIaV27kd1Lr1d2UIn1g6tL3MZNrWhh5ETPza8yQ
rJvy9Ktj/hP3e/96+MM/RiuDPmxRnzngsBa97FWm2T/Y95Y0xfbvnlbYAyx2KHYT
e2IU8veO8JQ8pAECYdTMWGrChOVNrn9t6JFIhY5fx9OcKRn3WmlvtzJ+vbOpT0UC
AOamK0ItEq8xdjAyh9F/SjqnKDTPFOzYTfW2970QMqs4/F5Sf3Q2lMVTpD/HF8ud
+ErhQ6Kysp0AdQbvq6WOmng5HPnmUDnrraH3nBsCD7jWP3NlG3eFzwmoFHb8bdwI
MPLbjBPMSfpkqUXjo1t+De3NS2a4Cg8+B93Kis5y/X4EqJkT6V9yFsv3C3R2YoEi
LwzTahLFIXgj4sL6EK9CnPpvLOh2BvgqML1uG/z+DLtfaYQfLqy7DHKSQ9lh2iHD
YSLlvSw4YYb+zOnN12w4XDA+6RLAZXuOIn4rXWI6ynlh4sX4G0FUEPGplrUZwXGL
3AwnYgXbWSTgbE8GcIwScuC8cRSlobGxaY2/tJYxI0VsJKRw5Tlq9/yT5ZaRJF8d
zQqSsmhk65B0EwESjxSyxipXm/hmWkKJ05kGSq+boZM1yeirhLVNrpqGsL5UJwPl
nGgPeHUSU/KFtGrAnvxYiT0tlslDhWlKToTQcUm6AEhaCxptGK8CslAo1Ubu7aGg
Qx5DtODgpjmbbHSS9rpf5EpgrVQt/dKfw3mUJ5Uk6qe394Lk1TVkANzISKJK2DRc
r5jVTjl+sRo+FIQd3SCT5OuMQYGGKOwNDr144LcNA5rl4scCOoSBPk6vKm1A8MFo
Xo3nlKeIATN9LLzP5WLn+5DU08DSsRkA8y+JTX9SyjFCzEV4VzfvsH7NnD2uZVKK
wgN0oydcfBOPqDRZXc/4E8gtqvNrO52IjPcaiQNlMDfP6AzDbEQtljhQ2Lk4Np5E
IfBVVIor/HcD2WbcvttqllWtTDvDLEXnUl+7hBghhMTX0P6AgZoGWQa2QCavsvDK
jI0PDTj/Ew8BtjiQ1ZwJs6H/TOKAZvppI0+AtZwpm+bhbGrvV9wGZi8PxPajOZta
RQDTRaWGJXmirtrXDh9JBd6YUzdDve7LkWWtRza45RJR8CSkZ2c6zUJ3UUmux5TR
2nlOgcm2mfP3x6rkknNHDlkDOn6m8I4rcQVGGHTRGaI4ldVix64+F1cslMkoMPjP
yS9MBtrs2J6zI0HghbT1WwgdxuxvA88uiCZVKm3dmdRf7Kj88AqUQKPGZsYyRarI
ZNm7Bi6Qj7EvYBXz5zvcVExleC4+8pN25lMbZ0W8ey/eTwb0xJsfrsAApgqbTcer
Gj/bhGSr/HV/ZXWgP6i2H1U9dY258Saa2My/3rh7LfHPIDmAtOnysuCSvmheb39a
zfKtFbGaP+snSqu8EZr5PLxGdLFIT1T0UZfX+6Ty2baO8RTuLBlJKV8lA3LVvbLt
f+B0TO/Ao9kE40aN4O/5aeF02nIDJIjyqaOSkxKLyUzb9gkuRM8ortpylQ2k2EA0
BKIT2HFzwEN1hqVa/lvqJnHSZaKFgyVqpxRoeKk1vOqqojV9Xy++lDraZnNHhC1u
fV5DCBc9iw+nTr1zn17Y60ewHb9vme/7vjL79nGDsx0RpKrBEq2bB1S0zi/gtpWa
btA8SUOrS1x5Mgh6+nKPlhSdnQyTK74/y07UOlvDO+1V0s8Rd5RNcGQhJeuibpAX
rFJNgmonlqLh6KN7n3Xbi8jcksCXZUFMK/QYv32O5cv1qgS8CqPU7UqY/MX4BFxd
CBCN74nc/gXWFlssXVFwHr/X9JeWRbqx69/o1uH+dW+e97WMLEJVmujHO2lIpZ6V
9d8oMPK3zg+djiiYTP4qRWAv8/d5CBdnAgixK1+AMsIvxTmH8ZWAdPMSDPqHmIhN
2WbGGnAp8j22akiKc8d/XMX6zNJ6qz/GRsCuQyWleLOm29gOcjnR8Zzh2b447cKq
uMeW4XsKcHT7BndfYy5ANx0i8R6u4bfjUH2yYHsZTfV3RLRDihawy4l2TZOfGZ9R
svrwMHvi/i7pnMAO0X8snC6SbLCkS3ig5EWK/E28rBlGBnN3pZidyyPoTESekzaj
yjKn9nzd294FBUqoA1GxXuQroeyua7DlPlyidV9LGac2wqIKTq5NMTaAJgJDB/VH
J1xEy+JZKYxeDVly65tsTH1niHx0pRIsh6yOn5Vlnf490JpgyYjXzQPzmgSJiJHj
udcDRILS7dRI3Jw2l/FVN0qYKgSl0SKQAhrfeXtf+4JE+z28QUMCtqYt3jgAmHAQ
mv98s1baOxPxWnZ5kbyP38cOCQ05d9O3SLPIK4kvlVyek4BViOKX0WlrQrPMcqAD
xk/ZX8nfZOHg3QD70Jki0c2iq81IcobvIPdgTNBfaYz/uXm5spO2eF9RdUd//1cn
jl7LYWjOzrMHpu8gNSg1sPblO0QKvPA9zRxebRh7CvNwJns/BBJmvqZa57gGZilq
KCb4Y9BereKDEnj36/qmwLaMazDdQEP/zeJMelmjN+w5E6FfPcCeBIrEE19wlQuR
xLxT1RP+0COxcGhqL8tXvSZ2nT3iFK1Nj6mKUJcjlcH9kaP9Yl8rCXhzZVZPzaXW
igj1O8RpgFQ766FhYrCmcjsVuze+EDhlJMxWq5Ut2mSek/ufQtdtJHbXmfuodWqL
3L8AQPX0Jsc2NfctSO6EbmmHJZF0fhZvuz4flEbb4Biz+ErdzrqhMsCuZ+FPKNOj
+ozqi3TnMn3RjdwsSLCcnSV4LRu+VK/bwZ4TcQcP1wxNo+i594H/c6Gvls+MadqJ
gFOPrTWR2FPnLzJZlVh0qi6x6OsiRQV4pWKCNi258tML/ZQnpN1tmpvTTP0tkezQ
50fyNmgpxXsGwSr2rhM5/ts6p2xJvR7CZ3iFc8FdY6FlW3Em32ATTh8tE1jQzYzt
nmWhXC/ADqcurjhnQB8SwAJe5Mig4QTSagny2IGcul/6lx/1zJ0Lb2tBM8lp0n8x
1XrU/0g5YPDIU3/umTbQJ5Rv88alXQEObU56BbmrNZiskbMNF3FFyO12Ez35oxcK
UhmnKlUkc+V1onrW7sibvBXk0y+VoO1/pP+w2uunvyBRZqUCg336DXCV8BNt0Vbr
tCJUxT5JaDm3ojhXIAZ6uMVPejAaVr+oIHHIkklnhOJpbOiKCvcKSrl2URdXws/0
2rhfab3pYhfPXHPH1XAo3saXaLgitdDT71Yv+bZ7LRE5gnzS5/C19xwmsKU4hGhS
Thc3AN4H7RaDAcQfmXIvByYw3urqjKXKELWID5NYM1rYXut8vllm3KiKJ8toKkZv
ri8Au63pOXgScrwHXutC9N/6KXUwYSUgw7iHDLu3EUVicJQ9XMg932vysp5MhkYa
C1iKK6MoJ6SSmQV+XWB/5AnNY4IZlGwmN7qwqfYdrgOWNubXelDy9s8yMf6+pHEO
wYVbynbvahnwX8lMW4QP3006/GwpCUkQPYPk4vK4aA+BguVWZa462rWpwIk0NeC2
0BIVL/GH7zC/0KR8KWdtpk1U48BBROw4nwmeGwKh3Y2qDQWStWbhoHsnml9UzC5L
bDdiKu1AyHyKOzi/+l3xbeSjh7JtYhS/gf3yiYULIibJ9Z+O3J9u/5MlF4uikCTH
fjKDBdvCRWtXvNl0pya7K9TU8LvuaQ55Lzv2pD4Ef85SeD9YcL7U8dv2Xbfhe1Es
rXzC2vTY904H8BYOPNYPU4fP3PYvbkVzvdTxi5Ddbu2xtVrRu+ZwF67nestZ2+M1
+b96v4YBew9HMru9AnWiN0S4y8Shn8XP1pyV+XRZ4UYBkZE0JcjBONc783SdjY0/
zJj2Pda2k70F8jmHBhPuqKg10XkIJemp1kYjEaRPPWZOeJ59j3evPFQJBtXw70s3
zOQJ6E2hlNnmQ2hecYqyaWkNfBHsBPH1SG8GQhJ94kuxfB+BWgAmgMNdB8rcsxdN
hqTvtnuA1bZf5yYHNTU9IDdv5X7aYKe68cChWTdBA3/eLxFv7can8Z2K2QUttTfo
pXD+QFm6/36oQVVth3THAm1ErSRjARVu7NwCeAj8tSsaEi35UKhmVTNN4W9VySdw
d1WITMsvwkYPlM925ulRUw==
`protect END_PROTECTED
