`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SfcogmfsSbFpR6PZuwDtmnnz9N9/5cVZ+ZhZMZzGrprR
I4jhgvpb790L9RJr9ZgsCvCid0BR5bYnO+gD/ACJTzBKvFTSWsPpGm03euU1RTNj
23Jz/isyxs/mSWPARCN1a42FfbgRPqJ+1njz1djXTMxkO9nuWVIGhkSG99Fp7UDG
2DU4KrxeC8JcynU0BNop+Cd6RaCConbIxYtyMRxBlPVnZUXH0iUkkYZUBhB0pxjz
5Fk9rkerSiaF/SaqGBQJk0kLuD0njoeomPKtjOm77Sw8QWpBkkfAgGL97qX8XCBV
oXX0bU3Ms/NvDWQlP7woprRZHuQwheo9r0NqaO2ZZfDPP+/hhAOJEpFKuiEDdl5w
XFxhxjBRmKvv0L2kELsyaOwegnoUhY/+pK7+826w85K//Zk/u3sIZqEnmVJGR53j
2oF0FMIlML74Bu7mw04+Ki3oSKGCNO8N6yFFCptb6ii1VVkJ62ZAOIdwiqB3nAyl
8ehnvADetItm6cXXQLb5RGC3XdoN0653lRgXyjxjLEN6yBwCtlAxLytJDt5lcKzM
hJdT5E5k26deK1u+ItrlpBRe/g3ErzPuvyLA2UG3/W/yYvZSLbmHwUVlacT3Qleg
jJx3DPXggKyib4YbYwfeXjeoprnLZ1/JGZTWRu84/KUUKwLC4FEK9vvD6p4yqp6w
NOhQqyB6lnh9vEZ2MGe6zygPer6uEe3QG9gq6Ki9H2mYSSp1u4JwoPb1fOEfzLM8
e0vyhDcmLojA5sD9Y/ZuEWU1BKlbZ25sTT/Il4KM5bWklMtgSruJHeLkf07FIlbF
DdNxG7oKStj+7Mmu+nuec0PMrs3Qe4waGVhcznWtPjYAIIcRgSdPUTKPKOGqTKXo
Pd5arJ1CS8Jx1g5k4AXnZ1+6X0sTATqMNS6Y1hjTLycCkZH0nbzYBVF0385DQ2hd
zuCRNLzUUhMZnWR7Gbp4GKj47CoDE43BaTSP8yIKvkUVOvRw+IddeatiXDBzCdrR
spoK1hYHDN0exntW6iqfmkgNKTyFv3Xr8BGRdKhrPJk9h+CLfb36rDTDV1co4g6y
d4j4CpK51KnrZzdmelvnHlGrfcpmFJ6hVkfDREY20JkvUtl3sxjOQygKv6jpm8/Q
nJPPa/e0aKeyNhlyffk6mChNW/0hsAMtcB73xzSN4WHYZ6p5x/Z0XKiCKpSyrpg/
Aqnh9hKrJsXjE6L1H6hBA13L56vtS84KN1E1ynJQF1iDtIZc6TnVyMceR/C1MoW7
hlxqwUMZ/PzfVM1EClbGEdaD+lVC44VtKvmCmCV9PPBi8hHPFdsfQxJl72CfGhdZ
SuIPlz5+sf7+ShyZQCpRaioU5zydvPvLVsLOn9uUk1YnWSAUU7cEiNUnBa7peARb
/+9Xau/wb/B97mzsCts5irKbUdkLSt/rTMSzAbaIRSi1Xgb8ZfKD1yww18OBbHMx
cn+k3xomEcm7p+FnSBiD3MiRqwP1RK8YY3bhdsRhLGXVAG1xdn89Ce6goBhQto+g
H3FB0E+j6BQObC6TxaQpgxylVvT7sN97PToIoV74zt0VghXuXUSwHRXshEz/ZOiY
CbeR68U2VqcBndtYlyyeP5kYzTL6rCAq7aezz0/FExlBwCERZKUUZDAZOvAPjivf
QY+euwh5dfsdYTpzNFbPAE/jIMSNYz8JK2f9Rp1jTOmCpdyaS8tc3lsH4SYVn3Y9
uZDR6dbnRlIPTUe3xSzZu52WDvhrDI9Z8kKrpT2+tCDB5pS9NOAx0ldnrAkAug+d
yUX1VaxWi8EuP5rxuSCKriqVPRqeZzeABgBO4CaSSsZ0aY7s8Vnwj04bxRSZVJeh
qoHOuPHqX6cKH07wOrAswq0OgqKtIaVofgnaQWCoXHuJmiOWeLvpCGHlGRRx85/9
7XvI9LT2IG8BofXJbdQhsRorUS821+SjGysnSLrrvitp6gW6IdHhsCf6Fd9MsWRr
RJ9w516/m9S/+gyi2Y7ku3KtdkeY5xmflMmMsfGIEWS0KIUrdIksoWnRrAee9b8D
gP9GOZG/GKb0LQanc1J8DjeI49mDICcG8aaDMB79RH0uEDEbzgTQhZAyhjZRbxZR
344IsqHBfrNFFaKJbt8wTC3o/xuoijeQtiqjegHBN3PgHi3gfuTBtCkDlV5Uvxy9
JgzRoefd/p+aQH5ZpxppF5Z0mmSWuOzYWF6rdcWX+iIcRgKs06ZXi4u8rssIb9y1
2/Foy/gaRdjJRqvptj75P4HFCAOnSjJ+uvTXdtARToPIbAklTmX3MNJFsWqjaz3z
nuS8towjHPQkuWGXbuQJ2+PS4kXkJKbFSJqbthnY7v1iqBA6kuVN8XorKv44F+D0
udw+eJLrX+4vWn25JKolwflTtaircLInUj/1eVggv48cCP+6cY7IDfpfV335kG7m
CXhwFzo8SMtIZPCVIvdp5+l7+xWY8qfhCUb9Gl3RtyOWZIDjim/3xjLewQYpSoxK
lt/HnTkbUbA29H2Lj1D23/j4TKs/D4SAIHxr4tH8n9Iddx9ufPnKhfEs7Lz32oRN
vtXtzSH9KejlRZdXyupNoQ3qvl7k0Fvj1CbcaZjU4TZ/eh1ZjXyDIYXWUrnwiHe0
48hYjI/3hj89TbWSqIpZZbQb0qppArSCfMPIL8LCCLphuQPgyigENh4xzziXQD3B
PH6jrhx25pW8TEB7rF0VnK7KZOTFFBMtVt8cUemlXUfqH0P+FiqT84Hxbf7Uw1jC
gcW9L9KwJ9yoNhSMPOUKjsT/6al4DhvPD0qUojF0455eEEUFjB0E2LERr8KP3PJP
nAkk9OLwVW588msnrLKYVw==
`protect END_PROTECTED
