`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
wjO5Jt5+pm3XX6KVgsTCzCRDgAOAC/MsmswYBD9cMN21tEgOoD8XJx4dmZAQNR7n
Ba80ul5SAsy6dc9heFA5sojkJy3VduXBgbkbVT+vjQ6CYfoU3c2bdNi4IDiV3XXq
OVqORnYyRDWN5PRwKUG3Px6Nwrw/ys5a6+/G2EnqwrgJdu/oNf3EltxT6cKCmV60
j2fJ3Rltx9+qT3fyBDxi5L7HbaCzA8C0Ak8lyFm+hAjQmpgpTdXvKZu2XRT/z2sb
nIbNgWWt3sJcVkDVOmIQGKzzBugfZtRJNEsvKe9a8KQ=
`protect END_PROTECTED
