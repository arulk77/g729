`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
B+V58Rbofy6+7bX0q8pHkrThMKOmjYuAgoYDVEwxV/RMUjZvCmiQvQhrUNdezb2s
SMYMXl38QMNwNwf2/4IFRZpynq3rYHQzVPdic52uaq5iCogzyMWYHVOxtlAgyQk4
i0J4Qujs/XDFDzQc+3n9lZp1jtGci0RLXaVY1/zYp4RQpm1M7q+2fPbRHlnnoefm
PDeN29gFRAtx8la5HGLBgof2kSSpf6BK6dMcgvvswpn/EFoyvBwwIzxeMZ/iFpf2
HzMLyuhtgASYmDVLs3GYGNRmiubvuDgxCRtv6G7kzws=
`protect END_PROTECTED
