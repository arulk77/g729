`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/i6NftxVpfSg7MdufdZr4F/vL2h5aEI1HLDJiKA5+SJ
HB1I8gFMMnnGBmlTXB7Cy8kceSttgyDRTIAw2BPCMWGWtrEoJfLnNhx0lQhkiS9Y
q0GIQirKq8/SX1gUIJFlVpf1704yMLo3wPN2ekK8gDPF7P/tfJg5wpAJTkpjIv+K
hOHAwQREEGgd95DxuaN8CgTPuJmU3yiv94Uedh9zvDd08L8105aE4CaMCR5TdS18
N/aJU2LWilf6qCZ/UvCaHzoNpCBG1f8Mb7J46ROSHXg4qOlg2i/UT6WhmEF6HBg7
bMv3XRpHh75oRLbk0J/lERv8jxiVUZxGbQDCvoXzsn1JrhUIcEqvdT25FJhXb8L4
hax+QUBOoZA/krMPaaswZBbFUpC9NMeGFXqXY25rxDISgleh301wF9o1h+jt6GPV
G4pdp3skxSbs2pDS2VHK54yiS7WldUsb28LDDs/XCRZ6pMhEk7ki1fdatP881iic
`protect END_PROTECTED
