`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAb7Zg4C3BSHeuJy1mRtKHaRGomtR4eB2cdywUTkWIvov
fPGqxfbXywyIXy7DGpDhyfOVzf9B+N0W5RXzQ2isqQgMWLeBqeHcU7sKBRFVFFUv
F4px86UwBjRdBhXsTMGSmzAweY3Jp3k7LHps/Pmn9PbhIwuVH8q/8yf4Dbn7Al8I
ruHgsKk9oG5/LE0FsA2hlgx1hJEHmUWP7TsHxtW0u+arVxhkj8e2RYHgNMPMCTCr
QGZu5uEW6VXSqTiYGtZzFzgXQXSJ5BlWEOeP5AzTXyynsguwwwbxA1EtnFwp2Zb4
ifOvfNqfMrq06C0s/8k2SeJY5J1x1WyDPH6pAWeJfPfzoHsMAUt76hUVdfY12rTF
uYVambxzcZZsjcLkwIksqge513Y5wuXJWhxBFozYqEmoa1bYI7HcMV+hqHP8wgkm
SqwycH5eUc5jl0x+ZcHwapx+1Zz/oRhRAhZ0FSObtfkAAfoOS5/Ed7wOSozzm+kk
eu9vfktgEa0P7iy50Gp6Y2mHLJxB+Pq2hS3iMU272Xqgx59euFL8DvSPwstFQ9o8
RXQoxDIHU8tlOEI3RIVWmqTXaLn7bkSKzHuNK2tpJLeriN8dRYFgXKV4skTMtdb7
OGI+vvvKKSvIlBVlqdIZbOGL4wHMv10bDjy0e6/xyJtHlq9n7XGX8vT7BwhGCPdU
HO8nkhSD+Nh+DJijiDDJB7qRmGkfpAHfxQUZRy3pWDbc1Sx568EsntLeQHeMTc+T
y5MmM+nXQw1bh3GSxLTxoJvgHTr58yhOEIP0ESiUYdUiNvPflqA0FNHPw3A0v+kD
OkehY+0qGqWWCFoC3oflITpbSX3fQGaVgBlDPHK3tHc/Hjpm1iCiNU39sJCx/Oe8
6S7xy3++ZkIydySOZGPnYNcqkdYGJACs9pub5Kb/s9Ijey0oWV7NPmigzcHkue/a
nkifMQDD7BDrM+0vl0ew0QnWfG2BHm1JaPxvKzeVmg7G6MHN33pRtLQZftvrDLpm
RxTydstwuR3UGR5m7UKuoArBWocMJeS7SXeu2ZyTTptk9NeOovGO+psvNR8iIbpB
5By6e8y+6Gz4yu785n62L1/1SWkbPm10EbcMSR1svewq05VOLkgaLGbcMeKAMlWK
edUsHzi/Jrpc8IEbGUfSBVOLOEfH3l8NufjNm+tpg8nE8R9N/I7Pj8buR++1lz7N
K1wrMuEr5bfR5xJPxED2ddpEtHgqDf+87KCmyXo/L1/4Nb2gz3ndslwhKXvawC77
FpzUbPuCH+w3wTHeIiL367ZG//qKwdB0lfyWAVnSQ/DlUQhTAe+gxqlTfep9Uyya
5YZf78BotW6PQ46Akws7S5jmnTI2jUc9OFJhiNWsnuAMgBinP3+ItUjjw9Qjov0K
ItoLYP8C9hQL2hf3RJO/lYMyX27nu0VJKP2SBmak2agLXTYnFRt+dGH9iSdGexLw
kBvRQXg9YYefMt3RCJEg7zvsJMiYOZAvRTj9FrMEJRq4HqHpWVKuGnUPMX4Qx52w
7jR9A8+SQ4L+PHL4Oe5Zp979voxNBZcu2XIM9+hApyD+q1wZEjwH5jB/axZviJwv
nD+KKfhzFI0YDCwJVg2EkiQlkOGIkH88hp8d77rzYUaUUoSWHIAyU6qdx2fm9O4/
ow9XWno14BS8sFaOxRWkw79daWdlvCQlKmSUXAJhLgDZdMJZHpY7vzPHiou/bPOq
wsBwO8SkJlolz+odxR3qY7vXtSHI/90GsLqsxL5xjF0hRSvryoGYR1b5ahRGzVPg
Wqh0CJU+QcvvlptqrtUfgfsKZGHhiP1j87QE55s31e3/Wai6k5/Ohw/4l1Nlkge4
eXuLBmozXTDGQFehzuK+wkUjgoCSnrLJ167ne69mLKoWLrYCTaE6+5KFYkTxXct7
PtQdv2rc+PeXZ6QbMxR3U1amtjzDHcXQYxjpZNhtRuKGt5BEuORs/30L5g2tURwe
/3ITxFfWuRqqq7ot/k00S9+WwsoJhfY8YKTwdSbcvN/w6/F2dnQGJHJjIQloXlC4
F6UhjPJLplmaDhyiDWpkRxJ3J3cP3jfANEqiNrdW/RweFdH9FJlN1k5Vx+8cWWpW
tbwjaNYFNO4QO+EiVFcVPoX037q8XHJY064a6f5xkFJ8cu/LI/YDaCcpLz7ksklk
2o6QTEpmp2HNNyYCF9InMsBBVVBZrQTQx4jn+wV3EYWEcTFzSCb35b8mksYhebRK
R0UI3dEm6O/3YEM+tTEvn2FT7hLEL4f0yAx0og0ldPuxH+NRNzQ2+dl2KeZoz+dg
qK/vx/YFhlKbmCW/mkjFQT8TJBqlGfbIGpa/bv23h7Ct+NyTFHyu7l6rZ/XtOShe
`protect END_PROTECTED
