`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yWpFLYwldw4O1Hz/g4NsEa67wiLPJwgJpvSdJBVeGMi
gQ26Grsw4/AfRlbGj9Zj0y3vR4r8sS87sj5BwOuZAkFoYL/e0wXdNwKAV+/RI2By
gA9wtWxSe6uxqthy5bSNwLq7ycSYn95FN56dTnBpSh4=
`protect END_PROTECTED
