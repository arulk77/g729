`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
UbF+5/ypEU/WQYmzAeQamMf/siJUFpzjgunlvTryYpXKWsYu+f2vjZ/vmVwJ9sHD
Oa0VBFFbwVrjTEa7tPu5EJckJc7yBIdD8MvReULUX6Tx+aMurvgrXNskw2q4ST7G
ll+EceXz9HOQH7vyXLXUcFjhl5G8XgGjbAQ6+IBt2TnUEWa6m63wP8lwGc1HDyN4
iYmNETuhmsD/nGAIItS4SjVZusi8KNjtT2Kg+XTSvfwqL6yiRn8eCVo4VdP4psq4
vqbAKh6sd3stJGSo1TgsqzRgxJeSvvTl9eb4D4LUlgkU0vBRN3qDC1TMc9agjbxf
Qe2zo1Q9lbNHJyIKhrSrESvXxpuNGKBoD6n4S823BrVyY1zOrIb2qhDZYMK/PN/q
1S5bHlQZTneGcMQ4NR7skA==
`protect END_PROTECTED
