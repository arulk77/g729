`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAZpw+zEwUtHd67prbXriR/SiY6SDlgUkXTONcUxLBlMv
RwELY/k31wdDsYAeOkaBQxp2PPm7T1EIfCgusxjTc51ECLCSpd+Af3QzXV8ePOwl
mKTUs11fKw0U8o6ka2ZvmubTq126YNTX2UN1dV30XYgqSOIhBobEGtXUhb5HV7cI
q3CAahnQNDWKaMsyl7B6NXeuidXOrOrJUo3MlmcgdMAAKHKUGz/NaYZ999Mud4cZ
l/9+HKpfIejrMHmjp+qGnD4oOaUgGmQVlmRI3k4mmk2RPPx9xWW8s17UW2wiu+0g
FcQxsWA890fr3xDp9f8sOwpbm4Kx002ORnyjXoc+NR9j4pDTF6uxP71ms56AHTsO
7NB9VzhkYjHjUmkgsslJNOyqzU4iAvDSaMYOIHbd/LvLV6ct4FjNGVLF3MaxNAHg
3DHmfps1THRwaP6i44hSvPJNww3oohY6aybPsiPJGFe9QWTKyff6LVO6tHyRUJkp
5FCA0856/a9jYcR5QdqAFg==
`protect END_PROTECTED
