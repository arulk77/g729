`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44R7CQ46pSrW3S4xonrqvN3gOsIs5YaY4IFNyO0EsrIL
5Cgdayly3SBHNE4lKq9w0M6ATkLDwbbStIi2CYeP7DIO4AGrkj33Wwwu3kLHLFt7
B6l3F1EqRfGGMPKI6XKFzmfYH18T+RvFZYCkrsrQHbt6tSeyfvIzRNdAJNOK7ohP
tOb5Mk3WKviZwDfFbDH0IL47sfuRURZblNFV0NZY90GOnfZolyN164cMu0+fOJuD
9XHq397z+6j0oCQpmXGlt+YEDOr84Yppxq7ttY/oPKqFBCmJr05oOQixb0rKFsAG
B0lZEy4mzpd/EowyX4FIn4GIFrOm6/fSpfdqmPgc8xU/Tle/HH8vcWSPtfbW7x5N
23c5buQVtxgzTHgUFVF+ttJabWkR4aCqdSZq5wcr00Ewsygh8GZh7HdIqtrLGnL+
z1fq4kwrbkh3cMe3aixfq9U1Vx2sCK1KPrXG9agytWunBxbGrMuP41Vw62etDVfy
`protect END_PROTECTED
