`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
FqiwodPoziC1xbJQy6ZtJh03NgSceL5b7L8YIVYXmob4egIA77NPJns+JN5caf76
I2YxUDwG/sG+KZGo4Oe75eb3/JSqG1XA+Hz5w24t7epE6jepd1QwKm1A5ZiVW+5n
R6HFCrwL/RfhRnsJuVWDAeQMuvgyQqvzd4k8MTlstNEA3fvkSHbhlsyooZu18Zd4
E6mE1rCAC6PYBYwQgaYgKbPPpwMC0C2S+fZ2qkrYQ9ah0ZIcdJ94VTvkyrG9V9lE
aupaAt8uXHk06Ft2T/ADVeZh4VkpcJNbNNGpEDtPEkeK2QrRN38bwO+0NZ6dsIBS
rOGlkORi33c8Y5+zUepvypVf7/AB7Bt8OyJsCbpen5POJO79xUW3NgCqRbQRmDFf
gaMl+EllCPClG3/OFiAif1V0R/vCy7sOCBKe5AVH89yZn73xMtNhJENUPHFDPOdV
j4WAyNJNapB8VsIXav3T1yde+KOIPKZPnTNNMbdJ/0w9fLY8tINlNtKAYKUuBL4c
eBXPNt5C1KeXMEuiijZVQLNjNvOOKie7HZYl4gaXAA90gzIYvysOyb0x/SY+ZKju
ZQes+XouYRUDm+CSayM1354f7lHLJFkt73IwWfby5GJb3ItwgFTU46QXTu8CD/KD
9iBmdwF5kB7U5OjX2AujhGjLR51inAXHlkYiFsV5F2kWp29wTBf8QS58Ai/b1vZ/
9BhkhfOaekBguQhGvTIHBEnuwa+xmEFd+16dZM+B0k6rA8TXvyXktO7CZQMC54k0
JeDqjyv6sXm/Zmqs2BLxjxyCIdh+FAVqjiyshUhJX4y+CVW+/+Jj3UmUVg9pVf04
uxuBfxniK2as3Us+p1HTzSz1migoK0x9zl2QsrLfX5DAS1lial1u0/PR29FHQYW+
D79b6avKR8g2nJWaJLROJIQkp53wjknfzOTykzwhPXkjjTWLLoFyCcb4E0eKCnce
ThARfORJgV9A3xfJBy+AFRZFchVeS06PHtDF5FHL02vQwrAgcOU+I8NVv2Feb2PU
Qld/4vKOHbURLzlSLVbCEsMEdCIrjswPNXkbHVH5SJIdq1wroTWJpDCCgo6f3rec
e6JvzJyTJbM0KzK4DXDllxoJZLq8B65k+knguNH8dUfwObBRwgclWk1oCHWDMjWy
oxEw+7C2fJglS4bwdhJBmDgcHIYPPdat1uKycp3UDX3bM3Iq9ue+bv08Ew6+5xpz
8jYA1SOUV+n5L6SAjNe8yx7l4clTkYpeXvbxbWAksec9K/1rtoGem/AyNdPeQ/bl
KYOpjvmSBDWlfZ7JcAVhqjl2kvHoYSIwYOp+MsVGE/IjmczGfBxmuoS9TvaqVVBo
LtwLmA5310Znb+MEXVOJ1JVHZbU1K4k8E724XQAnN+p0Y8KhVaBgKjQmRHyBuEHw
SXuIqn821Ta8eK39JUgeOVD6hjukViQETqjofnANENdnngyVnP8JTjENWiQG6In0
KPykPWHhIdqVlAjdzIevKsvgQ+i8klguepqqz92gISm9sp+q0Pxc6cHEOnP4dTMk
DZ+sNRrHUIJ4gs5No+8SB+CQXsRSlSzt9DTtMmtz5XtIPtiWzrFw3yZFQTz4THPp
`protect END_PROTECTED
