`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu477cmWE/nSerVFsexkXgs47BsUA6oNx/b5bW50sE+hcp
SibeHIcmdUaR+EIbwn7ImkrVWYEmM/IVdRcyKsIkgGMJdGJmbhafQD/J/4L1Y3Uc
YY8bAGdPD4bAfGMB2oflNo3qcjyXhoCOG6kIwGG/39I4loLs4NHmxWmgtbK4hISj
wA0suKmGzhDQSuQA2hjd56NWAw+kW0iW1d6O50f6ltTK1nvbA8yMbNniTwREW45g
yO32+8YgBMR1aTNZxRlybd2TmHeMoatz74m3+4F74f1Sd/yvTS406WBZXYHYZtUJ
mZlop53WHuzQDwXnajDK9g==
`protect END_PROTECTED
