`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/UtEt+7O4XAc2J8hy80kMcxo520O0lGzRwHB5Iml2x9
1Nsj6zTLGOU9cZSJS7IMAxd7C9PBMHrnMZAt2f6x9K6O3eNaiYDlrcHoO24Kjkwd
p+7UzyAB+k+cguFyVAD/+AF6CzQhcE+miMrqGtD7UKAZQAGwIB7F4ECY5d1f1bJu
gQy5N4uQX7z/q55z5WeS5j01NXgUMnaIYMYMoHrhb3B06sPEfRzC1eUf7DWy+t4+
Bwm/Tx7gwMO2ztDRyuvQizGmUq/SCo0gZObTkMzuDHyUCb0xVUjzKQGrHXgukioI
F+A9Sdecops+IgtdeQqQWw==
`protect END_PROTECTED
