`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOvfZRLWgLnPkqYIPKwET1mH+IC3zXZnIrPMh6Rxow2N
H2guuM56LTbX3go7XQ9Qv3+PW+1RCbiSGX8o4bwN3x/bClTKzOVnx7c5XTkUzPlI
CY4UFIRcNncrZH04cdkVMmVrmig09owmNgPcPeqdRebtAAELn/nYNPKK33UYVe2R
5j6/p37VR4tq65oQUO+3WxRepfyGWrfj9mv5YkKz0cfc71nWMb320UPIMELflRbb
`protect END_PROTECTED
