`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAuBzcZzLGG31bTSWsVFSOQf33WhX09zzURFLZ0maSoP
YEH4MUqUq8zcDOoDhhNvi2lYEp4U89I41/8qU/l18EmcK/Kfm2RoibzoQuMQ/APx
YErH3M61FPB2xtCuP7IkE8kNCra4N83WfjF4XP7LPSjHbgOR/97DQbKh4QKYJvzR
sGXb7GlI1VENT+H0GGdTU/osGt8OLrriuo5NoSASoK3Ff4qxselVomJJ3NEjWHMH
eo5DXUngfa9YhPeCrj1FFK3TWILFQ/juFCHy1KQRTN7fgj+kpJQ6Oxt2b7uqiFwI
wPUuHlKQJirH37esNM7EUg==
`protect END_PROTECTED
