`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKN2hr9oafgP7Z96DNdQJdzUfdPH6/li3kAVMBfc3Y0b
Q2cP1EeqH7535/wEz7iOId+QwsGGO410Y93u+yEBoUsPRXIKANeTDKXO30JfNuhU
moryrtr1oW+LlGZnQr+QMc0s7rIdHZ7FuB22Dr9uhAcCqv8HSeWVeNhYCzcbcSq0
GKRJotIq1HjFnMwTDAbA/KRPHOi6q/NJ5DJefAZ62qdyBBW1ftfsu1tUR+NuVxRH
C79YMBTqUzwAX3MQ86iarDIZnNEwY0UdeLCAk9zGMeoQV8x628qFXtmr0mqEEIyC
LOL5HGLSWX11nrZZkn5ocr44yLuAoBZeoJNm5FxiIVVPuxgRCTYHCkjxrDMql0M7
`protect END_PROTECTED
