`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu477vTQ+3Y42PAB/6qZF6HMyXqxuMxy8MuWlr2EFs6pqt
4mz9IP0QOIn8lnB12BphONpP7nonpCMbnfzBjVFVTVR+IE2+Ehs2EjYv+X/Z7k1c
d3365BIjRWyMzn0SzP9kzTJdkKFdey62Cw9L0JTaN/V6Z74N/zMG03S6nI7djzHI
1Ge3e+Qntany2qjJFDbYuA==
`protect END_PROTECTED
