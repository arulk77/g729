`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ySFxCiSJ1zUxT7rJjrxHR1pJr7KCw8uNQt1wXR2TuHRaDzFPTW8iUbRPacoTmV0R
o/u5VVxjhTcy/VxXd1hR33RPTchNzA3Urc2iobDZODB3XosM0CUUzIHxcp1HxQaF
Aq2efnVBLJw53q3DZPdS+ZBvfGIzGbGE6kS9lH0YnoXu3qKXVVNuIpX9s92QCwYF
y9BKEpPi9QlayzpmC44np1uDGueMNWkBSK00K1yU0XL9i7TdS2IbWwYcxXx2j2Fa
NWYgv5o0TLBycpJDrWEE4Es5VlM82PNRwacncmF9OSXYPQ2CNDeZYPgeZGKIbQda
NMgjh6sWeOxSxujWtEQ1O4JtoygQf7gzOdqo/CfzZD0KxZPZjWFBMpMpjJiBQKoD
oTG6zpbf7nWfIosg/X7pSWo8bZxyhnTIRtxwN5VyZ3S5TVSD6orJUuRGoZugcqVJ
Oi/j0gseaFQqABZ9lU1lPQNlbar14DbtJXI7hPXGgfISM7NMQhL+O3iMGR19mq7G
lGLX4PDh0VcuVqx5JVuPbzLCIKyJosYbFTf5k2/D0aOUh7eaPsmS+V1Z8ZHG5ram
czvv7vFgUXsQCOvK+ZwhWXgFlMsi8qk+spLJaWddVS4II9td7DaDtjHSI+dCioko
tYpjekZVJAz/co074q+wYCKj5JM/H2gcVXmJvQnuj2wJau+k32mNEHsR/8niKUmY
d96UP3C6YM9a0lcRRqK4RkHY/S8QXqwIAwi1EKHsr3f3xGOO3be+ppodzKSXnwkr
T9KAjp41bbaxQ0ZREKadLningfWVVtuQUCQh95cdi2sLMcWnJZaP1pirmwpyl5E/
/gJOprRqbCZc8BI+8H/BMwPHYwt1duwQyG2xyK9CPjMq0VOLSFoUVNclr/yPk/U7
emQO1OJii90nWrFjizERzVdil3ITf3SUJIg9uHSUxRJwejDGKdKm6Xt7GkCxEiDd
qSKYlvI3d+ZzKlTa7H+9sq1oAqeEGY0xVdPAG7tZ7n4=
`protect END_PROTECTED
