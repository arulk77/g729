`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43XJzz1dLWtEtOItb6uwzHagtmAImI6WFg2YjhZUN9cm
TOZQPRMDq2z0tuUFpxb7e+Ry2NiYxzrCUE43Q5PZfYulZZRQrlyAe/Dp/XJRJUXm
3EhQo45nZDs0wmRnm8DHOYndoNB8Nr1+RTrKuAQaKVykDmpIiZ9Kcnpe6pC9CVG/
GjKvlH0+WnbT90UXPTs8iE/mqh90rhzy7eqqBqQ+m0J3xeEBfWPzJpoZhAdKXoSp
ZHmCc9SElP5IJU+vG/aZPoHEnrj/Myp8gWzV1AH1dfmCmKGZD2sC4pF3MrUE6PMC
MacQxFKCJ7jGb5WeiUILIsMv9MCPd2OKZ+4OCS7293ksBaqoHRIvr2UYvzSYdoNm
dYLF/XM7fpXjzEYN9TCNYQ==
`protect END_PROTECTED
