`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48vKUxNwoUvSAp2Vg5ASY++MWhmszEJ63JE1eu7TMYWw
QHZEOW8q9Tlg3r+7FqxD6If2y/TvLqQZbSZKTKOg22B8S2urWHSvhZxszO7Aqh7w
oOhlnSwYXsOvFxUoUCGf1BSzzfK7Yc1t455TItDuFkHk+nBL18ABNwRjklW4bhID
NLwIk41Iat79Hsn8bAIcnA/UAN+/f36MXmWn5yBmvE83qK8UtxinxO5VqvZZ6oMj
o0JO/hydK6Vn/jNKV5C624Vu6YvRw/TB3Q4ECB8PhtE8+mjv7qxRAlsjNDmnZDde
OkRUbXrtvrnXGKwU7WzdjP0E94TX/YztqbZhM1mJaAPqbW1+4e8Mei0Q8qb6Sin7
dlbJvX3qIBHy3P3CTjyo+Q==
`protect END_PROTECTED
