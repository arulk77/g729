`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGCrIynsy/kOq5jv5ZGZp4moGg91P6Gy4Uy9ACaax2ZT
Vbqz+hcbAXyQZSs2Vl9H3pjzBAqDmps7P6RnosnrBgrAS+15cLt6v/6wlRdY8Ea0
jj84+I6JEwIv0lGkZSredYaxz8W1juI5v2NjHcbDrJi0AnB8E8qam5QIpzBliCww
dM1y0iT8WNMeizS33FSdU3XRqCqg3KuLpqQExInBZ1KmaMyyYlt6rrlKbUr5Q8hE
xeTDZYRvM+Y/AsPXSP4KZRttr9XXfIh8griv1rgtCOSYhVJ2tIe5onvAj43B/9Wp
TkZmg+bXNzMF9HPrBbl8yh15ZrvWt1Lpd/iXyx/t4VceOdYi3J080j5qh8NGqMm2
gmd0lwXkHb3bQbJa/7s8QN+s3d8e4c1A3DpYb8lB3ML+J6m5//y1PRRwjUM0jLhl
KvxS/W66nf6zDDLZM5b4L5Ciq+Sg3vLSpSRW6s3JFdLpMeKQmfF08b+5p5oCvz0E
`protect END_PROTECTED
