`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/ha0pgbcoJoyT66PnVHJNz2Ia0Q+jeIJtsVb1EBWClx
c9111wWVPlOhb2O+C2WJkSbZcqWaKwXMXh6Q0kdeSufSgfAGTRWBLQt9Swpaw4Ic
WNnpkd1pmWPoQZU574EFTHVo9SEHeSQw2Pb/QNRki5j4asEwJwiq4JqCmWAaW/pw
VScZLrxnAxBfFNQqHlCsxL3hgICZ7AdC1UuhBZ302nmCdd7pHLGJ/N9YmqNpOyXG
bPrE9s9vFKQOCA3+4XjFoPwBSwvD78/3ohwqYizgPmU4ZpxdG/1l7iSp08JgzWsd
QVvyDWLz+39ctLI7pqxppFaW6Ba97dugMUs9CiBN6yDhoC6Nh1jcQozcLOLD0YE9
ZKfHZrJ6LiUTg50VzaT3qXlCapLFeD7zeRZVQxHJ+xADTQtwNo7pr47jabxeR8+c
IvUL4HnV87rrK3PjY0gWQdImxaPWWrSzOVyM7YsRty7M7gZikXRX3qWxqVlN1nVp
SOiUj+BoBM7gHq6iwY/C1qrtA2zhBGc2rzd2MYVUaDPh5024qXrDYrYNeysaxmy0
8fk0E2mrfs4Xi1N2geD/3Sg5YZhI6ZHMFAQ8GtUMNXWUsCFqgod2sFkWCI6N4qNm
2Snslhty793Cac3b8vHb6z2PmSBqtrrE8R8ydvAMMbFQ2ciay75+STvDDF/NgCVK
4ZRqNy/qn/iBTjBhrKDMXWQE02zo7KxupqE5PSYaF/1Ed2wvdCQBJoCJ4WvYU9uk
i3FfvjmwnnwPSTVAUKtruCqluZ0p8Mak4WXD66x/y07/iDf5SzwqvAVeJSs+ZvBq
Lp97nlpVBXgoZMRXpS61G5wfm2lkuVyhDEpD8GwY5QunyVjk4cwy4Q00/Nh1g9vN
NKnnne+sE8pAT9Lr4oBGzANwlTGtE/C5x0/qtw8eFPp12bF5ylL9jT8EUwMhZaTw
4rg1c7iFwUGvTsgeW9wWG5KKicIb0hbqN3BRBZo0JoZZoOa+4+EGFEElCXHRgtm3
j3KuoLOUiBaH1ns/j6pCtsGm7PneqjMikwx23bWWTBBkixkYj2bJDFvdBXrFp6Bq
5A5zM0faKtnsiKfIIQvp3hFpvI8JwFQpbl54tgzCXVFtREQMUWsEG6fdYM1JUSYV
tDOcWb1k/SHRSrSBAmbclUmzUGj0/kBvOHJB5POtdSa9PzJ+Y1co782QDAiSRqdv
YRxM6/nSVtgHtgDVNVb5EgdppWbAsOkTWbyoreMDOEY8G0tDFwy64tT//pWTsEqj
1it0NE8IHWdSmmiShXgg1hDBmmTn6TpN5iFrzR06+RBEp4pF373mcxEn4EcfhMO2
jYw4nIr9BTY8DJbrwoRY91kOqGQ68Iw/3TKRsL+xmU+BehMH2JPc8BUKACzWNOWl
CgsYSwAFZLRdeiRJZLNBqpAqX89WcgAWAaf7AAbmGb8Hudui6Em0EiGelJsc48fK
OVhXjR3zxuwmPA+ceJ9eGWp2uZKIGFFCXrBH+oNAMHXKssI6HaMe4HmOLWlRV2h5
EimKe8kBGvG3vC0dCgkti8efq5BwL9EYLc9OW68HWO2eSkcpAZDj7AG0la0h86MD
0YWNZ9zTU1AiygI4Yrv3rlxEdPFFSS8B7taVt/Ia15gPwmz/RCNkprOe5Ew91B6B
o+C7u8BmSuVv5AtcCIx2LwGe20e3qbmio8k2HV1NyQZaC580o29FkBIPzIG7+CJ7
t111C0xDp+T9tVv3xwrEaL4jpAbjAEJj4up5RfJXEA/W8u+pewtaoFmzTNSgLXqd
OKa6/sRGfgPDWAHvpYh0FmOaw91qtYZXD7z36bxQoDUzqBnt4vU2iru5NbtymIzb
ka5QBuAbkBcgNF7vbfAnhiKlSFgHVh9FUBChTJzKZqDTV0vsclQpe32HYc03rpPL
sRtPPaPpMdpJ1wIQcvBqhYYFiv60RSCTJSTee/NoCDnCSY0HZBNp2cEjpb6iCCiL
ARfvWuAu+vYNyqVG1gu/beGAW57tZd9jWPFW5kICWctqNuA4RoGCuce2rroO9N4p
JGo7lcr/dohRevqnYVKqSsv3xVC1CJoqpBK2wvDnUS1Pnvg+Pcx4OjT8fh6hktq0
aopgBt6MD/dAizPglc0cYuHOL4qjkgkjt5QEYjxuaKDZBSJdsTqJQQjqzHWSj+0A
P4JdzG3afy489a3B/VL73ziq9K3gAXX+grJzBgsnea//l7s2xMw1U+bnm9IVk4dF
OMF9+TO0nzHUL/upXyTd47KTXynaU9RSoyTGgMZw1vOKboStWr5/xRDv3dGMzA+D
ZKJhaEO8/WiOXO/uf87ozvQ6ZZsPWM97dEbHL2M+GjQF1sSQcxA4iLn+gXSnC8lL
gRT4G5MZ+MzqXlsxLpIjAt6rUVk9Y8liNAn/T1eTB1aY9+XpiYspLtGYpKG4rdFO
I2q1sSe++RywDTfH1H1ZJdk+MvN0Cc9Eosh7SSoH3gu2ce3SOOfwiqqNCSS4RzSX
QrsVu8hgnCDpkD41pEUzAsGErKjyOEuv1b+wAyyiIkmShwrTXBejuldfsb6WbNfY
VkstXSXJye0jeF0uF3HIX7yH8K5M2UOho0/N1ipFv7/XP86TSrzr2WZamMles8vh
ikcfdvGCwUKB4+2tFh4p69rneVjWCIf2viGPPQa1quVtMyVb6rRqzshP9IWUuLSl
O6GHQ5PyDacHxFrFMwulCtZnrxKF3agm2mMAAp0sLg5YdoCfcZ71KpIm16XA9Cz5
owsL7XkbUP6H+QNWGOn2fIZGPIFN0iCtPmtNsu5IpxApRoWoPqjnwFqzSVFpvdnz
HdSZw7hsWC7rRzuwEnZbCmVaOGzJw3zOZIBicVGWR1+1XZddsu0NPQkTvnCKkMvj
Xsb/5sVnvOYyH2bPvKHexFnz6E9kTo3CMwsHPwrQknU3e6A4MnJYnzNSv8louz8c
nZIG3viKXhpF6bH6bx+EIQmyIgriXLhtDXIE1/zgIAYye+EC21E4RON4qBjquWVw
ji1/01XeT+XLECjPPe4+7g==
`protect END_PROTECTED
