`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
CWM92oPwiItjYhO/ecrBjEpIPSvugTCxpMx3fJ55zx8t9AqrHeXzx4S87o2L0Dhy
jBkLUPahIvml7HcqXhQRyk/9VcGYoNWNGR7ZbAGG17dIldYm5wuN+i1CvIPBzlQY
`protect END_PROTECTED
