`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Hn+o/wABvOtt9nMttJt/DoiDto0f5+JGskxAxby0uKdWdKkFl47E8Ba0Cqg9sEea
kMBL3KXTOBVzdA5ePsmYt/DMdSDcp/uQGy95xhJU+SxPM3aylUnTsTF9HtyCSeeu
26nAGz3ru4BFXO3zcreuHOnFzcjzIozg6m4uQuAllaMOFteOJxC4I7WkzBJ7b2vC
5k4sfzK2DipN34ukI4Z5L5pcas6/N8kOkS31BYYNpi8QoOLJgKs5qJ6BrAjW7540
`protect END_PROTECTED
