`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFg4UucmojGTU71fNwTGRlF3sHcOWGDvg5Dwh8h1CXKZ
6AM86sm0fa5CzrTUR+zi5bzK+KL0xU5HsvdmovoInOu2x7tpzODZV03z5cUJos6m
RNswnlwBqsAWBe/N2I3BTeTQZYPw2TM/kY1GUpLxuU+9LeIpBgO1r6QRugQtRI50
X7XW0eGE5IMiL52J5Usua6M6sM9IZ+Fk+O9mxsQGr8cFx6+5YOw+hCBWNEgvajF+
XLNn5yIWBioOR+H7vV6A/5m18FQz0VHJoElxn5iFcJmHzwKr6ooKbLZmnsmVVjJG
8c65WTNXBHn6vr+4Q9p6sfgQzISYKmWMmsdKXsdkBVMV8Wej1ZVMVpeVkzzt90eG
2rePXusoVlZ9PHbKkIjPmNmCWMHuyIwNEnEwIl8yQu0Q5z3OZX+4z4GNHTFOxYhW
DEg1dWiphESZhq1rGEz0V+USQdUt2G0q+AFqy+5+49HrKxqf7uICnz6RJAv+boo/
nbIcQejrQnT0pJgaN54FUsAZAYPvJib58uXgyzfkfO2Nao1vlXjIYOrA9mV8ZJPY
`protect END_PROTECTED
