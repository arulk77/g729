`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAVVJapC1AvPqqA7pYm5Kt5DWmyxS0PYjDwlcc302GpBf
LQpcU4dlBpPz1A1sRLvq0aXAyybnAfCEUFhtORtTfODnOhsinvJfW1N2Ek6msTX2
Zv/9WlpPuU1Q+ZO1UTOy8i01ZpuUPWAjY53hkBlsatvpnuZ6RxrQBQVo9ifdvmW8
GDYOtElFnL0O6g1QDMr66xR9QCfWDVv1HIgUxQlLOn/xzyzClO2PF/me3JM8t2G0
RCJJLtR5pEGfYQlREStH9abx79qQFKMQjC/lqpWxk6FueKWoVl4G661LNuEBVfBs
XP+VlxEHGmFb1PKBp08J9lxV5/PuJXJULCVMIpzwzIGT9tKdXrW9/MCBuljROqWg
lCbaNKsrPU3vt14wEGKHxfsLKvqbsjnXoqhBCIVZXIaS64fpgAo+PZRgRQw8CLZo
r4gf1wu1dS7TbWOvVexUOrZpiYD8eDQ/aW8G0dVsEBYnloTNGHBXJxbVxa3X7HdA
l9uj3HTqHH5g16neFaftmnHRO3ZwslcJ7WuyLWdGdZzfOk9Li2P2LudLr9aR9WIX
Llqe6mtm0pI+RhpdM2RLqiEHY1Y3rygTwKISMvS6UtBYW0NDsyWzBOSDp+h+zCEx
5farABv89ddwGA6bySvWUQkSpQsMKrDrHubSwDhXA+H/2BzwdfGI1mrDMa/pihix
efToGaab2G28dxG1vSJdbAi4wMpKJZ84nD5nKt6jgcO0VHxpW1bcbYp1UHZiuv8j
0f9RqhGKgrjh7eOm0Yji9cEKc8UAW/+18SWzFyNvR8BeN9LDzxlfcxqPSwqu+7q9
82u/pvUbHgNG8psN1Go6LiZIjgCPEs8bWgXlAc5mWqFoLo+bSb1WCS/qK0+0Z3be
YWIj/Zlxf89I95XbefBhW88i5PFZ4vtjvtZJjnvzOtnuubJqksLH2FXuV1uLkPCk
/PpaENBce0eW9uDfE/4xHh/N0GUD75uXddpWGeZJNACtqvNk1bfflFxiZtcN8l4j
GaZhoT6+8a68euKslVrhQEZ0vk0wFYz5dkVuLnViyM6ckb2jGBx/L7aaHnT7NkVT
Gw0UTl2SzPrLwV7Te+SXG7DQBuFi8YAIa7t9tA8PGuFYMxEak4mkJDBnj5FE1ddj
xA3y3VmOGs7z0uVir4R/x9Uo0u8BltPXMd8nBSM4Blc8L0tEbgrPfeDbBgf+LK5h
RD+2JyXGXeyMh7fTSGsQi/DKhX8LDych+oXfFqVjU4Hz9l3uso61MkK9VoG4GilK
ZyQJRWJFmnBeRNdABXOLBtBppQ8RLezC4NWcaUuT5A4yh17Aiqc+SDiFlpjyFvzn
RWoKY2djjC7sGpTrkoeSdr9sNAkbAuuA4HSQoq1vHgvkF5JsD0GioRIZyuFSinBR
IfbEywxKQx4wmiVpejj2PYZV4dF761hS2vl75TFRlymvOaM/twumeCDL5XOliauX
1ITXJKQh1u2oLP+hYr+rnke+rv39me1iR7uvJzQLbeMvNTPO380DOfnG+pRgD3+Y
/NE4HXud9CX7uU+UkSCRVu7QBZvUlN3nqTcHTzL3urDW8fUUO2eK1G2ugEmgJlvZ
J6Llb1hpSeYCasyQJRCLxpbrNr0mPh99GspqVidVE/7W1l0QH0HSFC0XdOCTc2vT
sw7ZVBswBD14+iYc8OikkYpHQKSZIY9QxG2AMe/DsR3ZxhSyROztl58bvcFZFly1
KjKVw14GRs+lCaeHbnsexJsq62AVwpj+2RRY9ViZEceuuGw1vKqra+E+Z/T30U16
1c20cI5Z5STUGI16Kmlpu8yVAchSrvNAMNqXLHF26BGhlFMNa/d3VsAoGbz2U4h1
fEHdp281Aywpf5qkf5YlDMYo8pxfrk+EEJ5XYOWjAkGodHX4W8/F4gyNgsLmL3GW
xdP316cF5abs/QB47T3w8DWTGk4YjqPptSiFuJuA7N3oZYCPYZWnI85abRVIsud2
zOz8XFS07LmSv4s6ubi2mpQzcF2/iTHIqf60sODmbzRTWG0alwcon8/kXePdu640
FRt4uHNkX4NfBtcquMR2OHDUMCLT7PgAWo3peu4xnadC3SBSPAtRl3eFoEcZacuX
HCIoMyXNk+08ml4P6mMv1lbOD0xubJ2nAfCh4XJa0Hx93E2tbXt6hHT2EZaYLi/z
6SjZAM6gLOAvRBP8e/hkebmBJFGV7FQ/1IC+NOT1fw5o+3/QPoZV1BU8n+4DPMXw
3Pj/SJigicq0Yceu+SOdnpzPfccEK5wGSqQMGcNJeNtqfr5czBgL3pYXgVFrN5x9
hG9NUVgm7HwmbZcgWIc9fPtQ5mE/WLdQRDcFTnDVM4D3YoS9XZrynj7awf6D4c7m
S2zsF01PLlXe/6mt4KAkuld3qlmpmmEwdyktX8CULX/BRLa3Jl0SSo3j24Cro5Fo
NmCUtNnAYNWFPUiQq1kUmUtho5mDjB6SOGmU18A7+EOM322ScllcpHUe14rjLzgq
40OUSOkOAKc3exuAE+NFxrKeKfgYmzUsQuuAHI5vg/4uRqmJrEUHb4HU+Xgiy9ek
sIZbnhq2FyM4YBAlqQLlDGdxa+gRxEf5AjktEMN177C0ZDjtTG7FTbtgpZVMsKGo
6E2jLj1Ih2ZyrhhtPrsWgEsT/wvCSQRUPRx64cXzXsCTeDeP8vl3q+vjdfgW+iyu
53ZDQbMknuYy5arhKd4Dm+6XN2kk5osfTwSX2nBIsFVwtfq1T1VU/yjqUzhT/HQ4
hFi55P1aS/fLdVp8JgtnsfvJqiaWd+6E68UIdC30/VILDchd29XQuQNBwlFlIO2v
qhEIzTaoo9X5Kd4EWHuQ5bnZWm4QXguXjnLeG0XC098XnCt2EZ3wTz0ZWXWM3UO4
BYgiQfPxxHVkRPE5j4G7ZJlgCCqgMsytLLC57ejkLerLpvON0mBtpuMN2GmscaFD
irS/TKnRzTF14065n/XIINkKDSsD0eZqO9h/hAn5w+ObA9PIo3baKWIsHTDDcqVl
Y2PkznpII45dKlHwVcFSYrPtQ6D37qo6kctSumVMWItfx3ZqyViuwyLj3H1zhwpg
EjRMaNv+3wwFyL/v2e76pfs9BAncHDjq/D3tKsq3tzsdSWoIPc1Fu6uhW3Mq8zlm
AJQJ0hGbSzLZJDraqR59ROihW+/HS6MHKPZATYV0E2YPsG16esuvDVhHQhpOlQeR
udme4/4fcQScEfc0joMrjOtrr42UXQNMiO5UE1+rUDoNCuSi7CgPvtlvnDeako1F
MTjC0Hm2HjiDZHU0UU0VDO8mWc6EtqNkrchxF0KsZVcPrgWJ434kRDu0zFroCufI
wOHVfK6YeTgvIMFPJ1r/4XiQMMae2Gdn9TxNJA1cm1jv0+QqpJjOtUIrcD44vDTg
rIrTpD1opXaHZyw/BkiLzlhrqLLCKMvVA0nPf4nvOlSKFFqh090yJMd3GdxnxkP0
y090ztr+jXxw6jZJltJYYgGVRxbTBJKqMLAy5QHjfOg37kize0mxBHTk1qD3+f6o
m1pdtN4d4FTbdez42u5FGy4ljRilPGdT5zHH7MMF2kiiucn2c6DcJlrFYvjSlPtd
+MJe/TQKmZBquOjeR96tm6wzNG3PKsnF4OybrHmdpatql8su3oXXJU4+Nbj22uqu
lVsGn89wLgWPgSKZ0qsoPjjxvkIygghOnXtaRDpqYP1gTr8X7BEwPxzF/SM/1Dsc
jYdxTyMzR5lDuE5ydBnv9fqSFChKH0+lY53NlR+q5uBuQmA7O1aEt3JBE8ubcgUI
6yLiFlJPxTgPCThVW7skMqje8CKG+4yRps8c5i/TwIySISpYSy4E2wxDEliRdzrA
PisSVdPMJ9TypbQKNDlBDBEh7sNYzP59Sce85u2Fwe5bRB69/KnZFIBGDak4IZDA
X4TdlnxnMZC1jvFgDYFiw5GzFuYidZQHhuRtasS9g36FJrUY0Vj3yk98toQhwsnQ
JA8o4WXpPE+2J8ZUvZ7dCtcJkGYWT4MkITQNJxsz+aUtX0cJ0n7aTpAXNApFd7yA
slD6ipMOuKl2k0p2iXnzhJ42yMrQ7DpktSOqzqNkcURvLZlmEpZeYJEQsQQwMyJ+
LDeGk5D8H+UTjV+laJ6B06GB53c+gDrA6+va09pyrMQ1ZOGE7d7Ri7OSFfaRljbJ
A2R2nwIsy5UOUhgTsAMcVdic8TpnkBulo3EQB1gsJKlD+SF14QIDSxagcqsMcrbj
KeRWGLb1T0f4AY2v1AZSAgHU5pboa9T7eUHVNCeswoBv0ei1GELugoVxyvxoRqZP
53SdwM3Ys1FtDrql327vS6grV8eukXt9F0xp5DKrJ3mmTjYTAM2lhNOZHWPvlBIu
CZJx5nwaBjtWUfcH3iVNKqoDxuWS08ELjKmNLobXMxRwnZyDmmUL+X0EQqHRtye9
EJfWzX43zJFaS7NVUjquP1q6ZPbawX760N+jawg3bauS8TIHZ2V6MdQriTXJz3YI
p81wSGlW8pF3xpJOsQeSsmxLAktbUUKi164NsL1mHl0lvzdQdHbFGVgy+hT2wtKl
ttjAqU6PxulgSFQSZjiCt6Iffqdnpn8Mscsp3y+45yfPUgHNvudcsltXKCWwqB+a
CjB+1DKSDepgbk3HkkagSTaAZk4/LSVmNzge9O9jdtzhU0DYINLX5jpszWNCEtbu
x3SgxgwixDpV7BASjExrV7EDKN6rlXvp2PM4fSx1qfN5rrmZRdKJvETDbMer129U
5+OYx/8hsgOf+N7ryHga/58rWNmbva7wGgg/p37uyE8m6n3RwAhaBczpoxVDjqT2
qStPuV6tDxwS3ycug1NU49sT1bTe6nqNAHsAyYLqmX05v12qo6HyRgnyVxbYr/Vj
2cnFQhvthEfEk3Zo5mCRt/G9xxWo6wYZKDkYB/3Zxfw/QFz7xvbs/+B+8teuE/IG
XbxwC0WT0YxhZ7pK59PAgmn/MyGSmQ1dc4sxDuL2GlxFP+oVYKa7sMDDUJ49x4v2
cagy/dhW8Z3jcndwPadaGtGPmG4Sj4TMUo4TXy68ZRjYRLCXuF1Uw1dZWJ7skXIj
tROiaswHFlpevCvKS8+n11db5Afstax7t9gH228sdFobDQOmjUCVMwDP4yKfgLoT
uZPZ2gEjzYGCazEQ0M4rP94gAm3UhKfnh6xF3qkPUkmpQ3kleRqSmIaOe/bSAf67
ENSlOq9WpsWXFx8OCalD+cw2NYpw1ZjHV9tQ+ck/gcmcWHbhxyW7PIMj/67tDn+R
pzbcITsDJxaxCPDBBCRqdzRbGLMkZIouDNfzMvqvSBNhVC92iHoF0bZltnUnNSY+
20SuRsVx1KZ5hJAEcIki8ORPX1GBxPhyOPjp35Kz2ztawiI3L8cgEVJlzS3/spHz
8tKMqXDl+uG14StOcH7RpDLcq0v/fEhDciLPUWc2sy5Luxv3WqX9g6DCwtt3dAK7
Xix2hCIi5OyhqRXPrKgM68Iq/G0aEgYNbi8fpHMgkKrZrGPAP4uBjKqPPjxhDF7Q
cM6QOA+vIcebxzRcOI+T+9UsX1G+YJFPdgU73Ac3i9Xc5ThnLlRTVEbK6TRZOBeZ
n9okGet/uaKF5d6TQnBcyo9wFLghKQ+bN43fvPHEAs06rqW+2SSY1mYlw8X+NzL1
1rl21PG7QMY5qxx/sXrmR3YhHPyz2B03lfCEjh9opfbZeVDd6ylwpRFwPfmFPV3Q
x1/surGokoqkS4RY5hTmxfV2KUjBjx+Wr1YScJD4uD8BIzthCbWP32VVfegGxkyO
gJgane8MUw+CLbLnP0QWLCQQz2RRCZJkW81vX5dhoOLZhLRd4296DlMcdTkoqOLI
nvxTwijEtykmJrHs14Tpo2D73+ckXX4gr3FkSSlIO7ZmAzg00qZ5dXohkhFr9Smd
4m/zSFLGfHa2VdKN7DTjFDtUyDhW55iCbD5GqS05XPpPjnl7TlwsjQbkUsFPbJNU
PoA6Jvz4hTLYZ8W7XkH/aqPFwp2A1+cYdOOM1+NfiulmKk2Bph9A4YeGhlB7ivfc
FMnwW4wYkkbK3gjobdB4Mcqgx1M+AL05oQ1GZA8geBVrbB1MNpjwk3SfXwKpz26V
j7XHxBnFmxRzh3PynipctiAYfox89dHjOha0xbzKsc+7liWJcbnRXVa8xUXvCauA
Xcuv+n4V633iBlsGbbl8KWeIp8O0L+Cke+UEipRgoxOePALqYyg8KXoO9RyuFeRh
wsQ2M2fRTrAa8oApEZkonupVCEs6T5akHge/dQomvXv8UYGS63UbGDnWU4LfntLK
iH3ZlRnLn29W8nFouSOrs1fOFDNle04zrdpIfzPIlCBCiz8Nrd4lRGxBcQVzejzX
N12tYusMtye5pJ94G8wkJ2Vwa6PO2LMwIiM5p+/iD/ldqKtv0vDloXF7WSTb7iXl
PF1N/ofBwYWXy7G9KMKeP5D81Y5cytslzGONtRuM8/Xmw/1ivaaP3jGzUmMpZgbG
esHuJqFxftDDyBaUEt8O5CH2vbVlUc3204o1nC0EOSoUr88ik9Et7gzpvirAvmWx
WL0m1Z6JuVHoLXDHkA64+8rhk+H9ZGzOfm6dJsC+zlZrvDU1LMGVaY83o1kzS0vk
Sz31PHl/eDOqABNZ5akIL1EmWxbLQ5dU/xOkFThJpa0yogbd09X/SO1YZkK3LOkH
Un+H7EThhmT2X7D7vjlPSpyd6P1sWxQofz35rkqtK4QuILCnRZKrfAdlICXynMWP
bKBfg1T9ymfSw7hKtZ1uo4Ab0bQOIX3POodzr0bo1Iqj+DQ+Jncp3HlGsixyHZPf
PIUTjnWI936UpRGxut+ds1fP1XwrUHTzlrkKKCnSt5a4Hi8y4QtLb0qK7APXxNil
tzerAVwAT2YOwT877qtzbP97vIvr3Io+nbOr41LtGCe3oUlHkkc8Ui1fZRv/jymB
VvbIVk7E4zmmBhoukuwcDtaZED1Tf5SY+0RL34VvMIpB4KmZiCJLtjMnTf48VKf2
kUhnlJCP2gEGubPFbeqWzUB0Qdg80TSmlJMzA9WYST2oSf+XCUSeoSuLXpSgQlNW
tYQYSxf4TVhi6MqyWxkZrN/b2toWolTg5Kaep2KzUN9dgFN3j7lFdXiKnOnoSAKO
h8zmNpttSBW59TTTJ8rOEZVBmENZU3naj+IwxAR3TNIVD4zEgoGJcE+j1pRhS0hj
oOfubEC/8CcZhPPMBEQOmbv4+Z4vp2SVoo4fIbCH47/554SGSe2jNDC2/Dmh5iLv
ro1tJdYVElzsa/pwyuBW13+WxHDaF8R/h56eYzI9xLvv/rY+E0IB3xVhSw6bYOXg
MQMtiWB4WAV9yYh5P1zDWb48zPz1cbjWgol7buFytvsc05oBTsPGX4+lWsAT9pam
v8OmuM17kGUxGmXYwQnUtBOCaG/7Dfe7btMw54PmS4Z6lZg2Do2YYMrdxGwxXmRH
x9OQ893oe/RdhXGQSahLyM8Jjn4nQWXRSl35B5L3CZvFkkByb9Wy5WH/Zw3OsxW2
KopAXSUpniJ6klW0Km3+nTnCaZz0ZMuYvsfy/z2Gw5EMK9XL1mOq3FFd7RWZQGrz
mAaE6XAOpo1R25B+Q+LITN1BUYRaf0vp3FICs099gyXjshjDsTneqiBbzAKuVQ/O
IsXbw9yy3XF8ZQl2gN5KryD934pT/FYEsHYXdHr97VnNPQP360GteKVlHJYRrHzH
uC60hQUZcjN1gOiWm8Jgfihqs5BtaYl5oXnha3POe12CuhVdGphGfGfP0YOx5ypE
yVxHD+4gHjXjY5pR9ABADn/MM/UuqYCm2k7y2BsgIgpOdOkckNsCbgn76JdAKvEi
RxVUjz6cbbfVQr/EOP9u7xGG/1Cm+nCkOd4ELlG2HrTr5sHrJHq5IXau5mNUd+Bc
63BGXBDWbnI655WR+3VyQibMtEq7TjBqV5vwAdY8JDC+RWRrMsXXesxlrVl7xro9
ehDIsnVZFgMHRvi4zKPiCo4OKVQJWX4hqgF/h46pKUOCjkSnWd1qBnV5WiVZTdKa
lJWYCVKsLo5pDiKHpW4S5fiKku+f0kFUZDubu5i14yMrni1vTC6ZBi5LWgzqu4uL
dbU6Xb7PiRDaiUR9gdfo0XOFYK0lxSG8Qhsr473YWtkKM5NPcT7ZeqxnwwsUFdSF
4GzW7gQdmegHmUDgGE1UoU+VtknhxxDJbahYhLwcnPsmoFAkubc04276a+XZy8ry
41gWeVEGGiXvVcMPlC67nyy/JBmsfbQxt+AxKXr1WPnRGQgjz74L1yjw//AECnUq
JUIIFUOLyPRxJzX6rGqvnE9qQjutHlj7p7yeH2UNdjtemE6e5rJuyRvXPQVeTViv
g957QpPqyW8HiP+qE2617AbCkUa8JGwevUKdjYmvZJ469TYk6rcUlOGMqi7/O8Ho
FkwnCUOIphxT+nwNTECm4j7maaKjCWWS0sZQVEceUyZhkUayR38xxxaE0vSaHtq/
jBhCXNdvbU0xbSxVaybg2XIrr4ciBGJQ7/4O3ecrbdfU/gLkVYoW2HiDPM7Ebt6E
+lOcF6shj7yBxreybRIz4P0Fo8EwqMH6tkM5xRW8SJHjQltITi687aPJZnrhbuXQ
prubySQPtyg88rbRtrnfsZzLTwTcdTFUL9JhuXlivgA=
`protect END_PROTECTED
