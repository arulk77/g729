`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBWBmK8fJ1CO3n2fZPtbcBGKMW4P/u5JN1grjXHHpEpe
+ij+E+nCS/DhiyjijuuJbgLZcCxQHyDcmdSadtgRMq0KFQVU7P1LDEmij/dRuRrb
Yb6bEwYb7abFY5FAylI6CW0pEwtboEaZ5XyBL5o215wNc+TaYp/bS09H7qqtxl5Y
ceVTE/d/Yi4W780KA9kUxQ==
`protect END_PROTECTED
