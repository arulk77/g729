`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNKw3gSgbeVXHFdUK8RzecU3dalUU6kfXZEq+TNOcmRL
4nWcqz10ZioE8/mSvx8vib1wFlHD9unItGr0iu4wKI3GhEyHMw7VLcInHdXphYAR
p9Ud5Ra5RwrnYTbuLEVZTv7m+v75D58OIwcKar/yZKXvaG+RcA03l7zZS+mfWYDk
0D0M1EV3sDT1+yTyHUBtcvNWTOeMVDS5AD6Uw97CfOJ1KyNfqldZJnblILJdDvhS
HU8IkcjTE2yP0t/SAV+tcvViEYD0mjskMUHNjkW4Z6g3VDsJjErtvZX7FGvgQ0mb
UGnUoZdm5R/MubVhAMt1Uw==
`protect END_PROTECTED
