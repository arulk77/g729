`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKpz6lK+9mWLcP+y8xGV5uN/ARQ72whaFESqXD+sgpC+
MYpX+t4nW8PFUoK7GGOYyrH5PZuR0o8H9cv7tW52dUEfBrjf2QV0/of6IYyy3/kN
1boy4SDuF/VfBSCpC2o6zCLa9m15GpYbgz1XdqLSLF9TazcRk6VriQnSjXP3jODs
0KOmpSoiC4QM5lkbBzy1I+y5lccoD8PT7r0L0mN002WiE86R7DLVNiTpMeDAbksq
`protect END_PROTECTED
