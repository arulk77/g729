`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKi1B8ucDM1WWknLi8HXs7mujdEZkTqAuB3+axODvUY9
a9br6+BZnF2yTe12XLe8B5AaBFoenEDRq/mjJ9J9+rSDbbu5xVkpUf5WAzlxYoiT
m1Xa6vsXy+0MfEsqlY2gjupihAKnyekUHyYmwSeKhpcTZXRNZYX1T+oS/2yNBhnw
OnQeLObrVMYoAT1hkdpBsFZ8kxRRfgP1Z8pyfY9tOc/t0+gFOsI0xQ4hD08kuXkA
`protect END_PROTECTED
