`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SUf49RDPlqTNnzXtVVgPD5MX2oloFb+2rcgLgu7prCSc
6Kg9HzkWvF3YcHt3E0/LFcXE7fojIu4Wssi6+ZB2Mp77gczyUpWHqjuB9OdcAbxH
1H9mPrTyHN1yKL1obryXHE6eVmX/psP2jVUnlLqizBVyR/bLTXZvFOLpHcBNcYVv
aQBZNmUY7uF/a0sn0+lA6OR0txmqSwzk2kq9wB+ENGqQy5kAxpElUK1RReNLfsVA
0Sk4yZn/LKwhe82Pff6N2ReYhJ60rfqRvbaCkWiy5De70ddTps0/0EfMMxruXtJo
bWyCgIZp4mNLrcDJj5EzT7nGU6c47nsskG9PukJDzRH5SKcMOgDdxOl7n7Tl7PzE
61FruvAiLc1SXNFePfoVVsfn+7tXzZ+tTylDjzFy6l1maQh5MITYCUzZQN2x58Ce
OSQiQJL9t9uMzS8ZqCPCS9xAE8JDG/XQ+Jor+GyihpRmrbO9p69djE+WPD6iTB0H
wbQD+eOowp2L9cWeynXvEwx31/YHb9mN2KlZOw4zMmIcNDg8ExzoXfJ+6QERxDUE
+BTeK06vqp4lDVDYIxj6UUGW9krzYDOh3jM022u/MOU/uggrJi0G3I12aBMDSWpp
cvLkcvP2otR/xEYUzIxm01E+tVdcbSBV9GY+wKTVr+gEY1HDH1eGi9yiICJueqDS
PEs2ZEGbBbOP4dMVx8zt/h2r/o/wd5QbcXJSY0Pifcs9czqzzLUerTUMAuOudU4I
eDLya2050qYeN2YNd2hf99bSqFGkLxqCZ4c98XTbgwOEuizyUIh4j/SLcLHzq/fG
QTvx71/J2N/8gznOlgLYMw9ynbaS6kOuV5qH1rXjUPJucfi2Qn1GWCh1p7pfs2Tm
ASPljfCreFVXU2a7MCFBFqw+IIARTav5uSFi+/OQC1Hc+TCYWXOEZmnUF/JlVKxS
Hr/lmyO3ozeIgPT0zsPuXJvBPGB5DB2Rg4bAUs/UVulawoz4JLG9VBIURTNdLdzR
+SbPRlGbEO6JlYe8+ZBE9L7oXjJyCRk330TNUckRJ+1848hEFU/M8HPWgp6MCcJL
EPxb70U70hJxHvLpWaFLJUz+5p8exRN6O6cy9yBWlfCr1STy/aWDNnzvwKWCTAC9
IsT7pA1KwBUqXONJVtIl15xHQDGG0jzmEnxKckxKkhuqt5zDpMyoOSpdncCfMhap
fWub2E9q8PXvGFzPDMjB05EtAplssmdWhAiHEp5Bfq+fuJijtHlb+cHNlRasHFOG
bLamDAkppqSzshVJ4O8xT95uCAmv9ss30oCW3jJsYR1/nrWM6Za0gfuvJ9OlJO1G
jwIFmfHTLGr6+HosVui+wn6kot7YNKP32IITdDBaHVsVA1faz/cr3wbMpbD7BjRm
Tfv+qyi5M4SC/La/GiGFJGovlYaFIYCzqDjh9DH+Ddxe/FkRtWE2TIFELFnH0HbH
bclYGlBIWHqJjWvKN/AdgTddv96tl2VWUdWSgcoMkKE=
`protect END_PROTECTED
