`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFrDjXIpaMl9sHBJ7NGiTdwM4xEMn8l7bqjxQ3eZffsB
CIwV0Cpeis6eRAKbhkXjjLEr+yPLROsp+j/gIz/EbVZCVq/1wydS6qqXAeB08A65
2sItH4jdP2FpLnrrRERTRRUI+40w/3PlWT/PF+fPJ7BljmXxS30jcYxRJtnLBcmF
cEhZyv3eI8hUptgXfCOlEnK3unZMvpCo3TuMtdJYl/YkzUd9ph+NHrQjwFA9mRuu
nssg+5xhlL+HWsQuLglSsa8Um6O2cYVVLVVpFkCZK+u5jO4DzKTCRvKHGvjiB6xi
pHUu5rP5RMHTAFhV1kEZ4uBMOEbTlEscngdj6ePu9Upea0XxQuk+KvSw918PgYoM
1INN/kc0gnekEDWPMk7OP4akf6d3XJtuH+28HJpRfN35BkMo8FG2AF8oEZ5rzE/e
kpcv9wrzzy5rf1DCECGtrjH/fyKwnjUor/Nu0WyV4jqLMyazq+0vrHnehOfO6H1V
ol8jgJkSPYaQ6JRo6oDB4ZtVttVsNy3Yyi/RuDqm8FRwWSS4vCkaZyH9rNtM2230
sSGrS1W5ufGG9BRpgE4Dag1PleSDtcUcZi2f+dK7p/2lkf+MP+nTiSbEoJ9fdLl6
pW1iRhP9RqVB7sycKK49hDJ5T7NOtFblDvwbo6bW1MrMPKGst6QYVQX98nrZYMHL
o32ud+vyj8w5e6RBwnNMIVExsEcxV/zBwJBn+P6PLv2YoaQyDQiDnPtUBswlx904
fPi+yS6V9yLZ8Ai0/GAojGnYCqC1kbirEavYWKrdHNCbS2f3TLN8syY5prC6/xv4
9dSL2uBRKyZeoi4mEE5VVeuZCg/xx4bexLuCGji9QNjazrVqogHCYiBaIAhwNIri
lnXFEyRq1gO90AOvwtkvffWBNb+6MjG5COVALDMdjBc4Hqashciaj/REwsGalCUo
M9vav5/Mo+++DaJpyybqkV73VFVYJLfYYlQq3sCIhcQLQJm4O7CFuVHB2ft3cwxv
mPjiEiGzsrTVK5+ypwTn3itDWu9RQO03oCrhNNvb2nZAVcc6x0hTQMlDnGa+gJwt
PxE1kfC+3DS64MThwMotAQOJ7gS+CrrV082BSETqPW2fvnSc3KYwqFZAEvfM2kOM
F2/QQBWDZEb2PDGhfkUeiV4knXF7xpvZplPS1NL4Z3kEf7REgnNVlF8FZj6BBq2d
iAFzkdAqL7VwY9twS9vCpBWmVAB4ST0Wco/4fu8KgBQtx6TCG0RedzL5sZkIXZpV
vUIZUqZGniOpwU/pQkTllWAt/+1M2Ywu5FgXjkjeU2zkXlcK4M437/Gba0fmGlVd
wYUNcQUqaPhNRKwlJcUEN3ES/iCOhM/1YnroqiCOj9g7Pxn9MqL9nLP9QxZSxOJy
lj4DzFqAWSx5J+D0C4TWnMosCiS3U+R3Jda0mg+KhfV1TMf+eXyqsT4Z+g3ziUrx
3lZlM2cR+JVR1etkDMk555oUihUX5LwDsOzzyNjCaQzxD8XkgpM813drsef3HGMl
yBKaIgfe1UHOrMrqaJAITtJaPdhX18Ei2g/nprB4sJ3VpMjQJDyhIUDQ15+c/Uzb
G9TV6VeeWcCSxQIMuK7S+8FHhKaduqoL4rr5Y/zOVPYJb9uSPk2OzvaTN2oDGUs+
e05vfgqosAnedIjZbdLIsC5IZcZ79HMcj6lW5nt417otoEPsNRb49f0T0aEc4+2p
B8GLAk8PqrAs7pO61ToxsqmVjym2EhynITHv40iYVNV3nb4TDwvGgbqFWktZ5R8T
mp8jLT1AmBua+VHnAqof+wcGerLOZ2AjLuCdk49cl54O0myIXyYnCmqWfTRmCCfK
fBPoKqOUf664teHgsSLhQDy/LyY2KeLAAIg5QaOQHCmhYw8X3XhppgshqgJMvhWm
Nwu8c15oxmwSgQ7CfJ+9NTRzw6ykvnWLxZGTsnZzx/+kRA7MomM7E8epA7j7acSr
uyposibNopu6mdZ88I66K12Pv+wcp+xNcPhJMuvXadyWxT4AgGEvjFhSOc3kmHO8
t9HVt1Ah4e7qgWwQhWgEeEMAQDA74kPdU3HlQUemhmyqpEBYGu3NVwsxuIWEWrmB
LgsPda57tDEMB9c197CElxSBO4Ed7JH8IKI6McmXeoO8DsxHCZwYoaOxVVOZMuRm
7sUJ4X2HoLZxvQasnKedkt/oaCiX7OJRypm5l6tvfI0/Jb3+BuTfCAdyO3cGhXH6
fxzgItz9r6wcxBuz7T4iJNtixJwtPY6CaLpYDVw8OYl3iT64D9FRFckg7shBuzFm
HArPb/8n+GSTVaAtqGClgIAmolRenpZhMVXlQzc2uMsFY3ZsAYttFv0DqHKkh0L+
3hCFY+1l5K5J+M4DHD5lWYgydsCCOopvYbnbLoI+9TzAq34oC6D2qIduBq0lPk8h
OCpZVK1Ul2Md+ZBGTX74UKezqT/5NsPcA8GaiwjxChe5BxIhkryTBK+bBPXyBEEv
sLXFC50K5x5/VIth99wwdv3BbAXk9UczbGxx1SRzXPLO9tpOk3Deo1VG6VZ7vdmx
1scND4kN+cSFwSVdps+3/pj2Mnqk1XZcS0vVx1ZmktZihTnWtO5yxlyLevZZ4YxZ
5vQ7QlfW/tnbd6cs7ZYpZaV2B20dkmz2D+Wgtr6koHtdP5mOJBjzafney5pskE61
2K0rqu9of1zs8hs3KtubgdKpIZbpviO0lQyPct1Kt/EgMgJszlWYQDo4zi/A7ck/
UHIyucDk0wkdsS2OxnQDf9vipbGD8v7YTMQqxMm1JkFFUlJYgX9Daq0K6zfR2vHI
PrIL+QIF/0A2iauaKFI2dQZm3XdXSakNlK97lud9Hr/qIQcLmfMeFFyHICOshfU7
5TouZmeKmbLifHjtm91P4Hqgg9VE3v15XRgkmpYRLb2oVavJKCx9UQq2buH+eSQz
Y1q+HYPnMtQffduysXP+CaKabwBQmYECRWTL7yN3JKX5sO82z16sUYwp5pedHnzD
hWoeXBGshW8qEsQ4T/zawhtniRB/Gwm9F0E40Jc9H9YiJM41wiv951uzJ274OBoB
VVK92EMZbTe3sJ0WIoHRQnia0Vp/XhUrG0WOPXWKcAsyxiTzIQExQc8o55GPm/Ui
oihxq0RYRq01khvS89mDZu5AsyTn7+9HHLjw3BMzl629ABQCqy6Xk0FenGwcm0qU
2rvYIyT76U1uUntcFn8MjcsUEL0taYHyu73MMeN+soTzgoZLiJmgo58guJhX6x+K
UAgAPaxJBVFxiODCPnOtHqeK4BgNfU7XBExm3bENlEUqxbBP4EAIktQsiwfxklm5
2mMxOBc4ZSKyLpXXgdjOldtYHdX2HHl+MU2wcYjmoVNfM7ovRsbM+7tmtJRTS9fU
535NlLjcWqsFuOU1ZU5L5EFtclz2UMWV9nQQm1z1/LcFo4/pCfidE6kCVhUxPo8v
Ldhj9BJe3mHHovc6DpQIbF1Urgi9b+Kna7K779+tgH8nmfWS/PtntEsTGw8GY30x
5YFQHvXh1dzVMqwb/FykpUR094TzdNVtGCv6C9EmAm0wQusv4pQcNGbQqEJkDfJm
orz8Yxcr/vTVK4+aoT6ahJRr8VD5LLay5o6gmgw+36CiwpfWZZxjjtTYAp0xQYzw
GT9j48ZslRZ6mFZR8QPB62/4bc2BTr3GDN+yNiKEgg/k8H/AGL/uoECURrSqDJoh
e92NOReMltNx4DUpScmmnbn/3fcsiWuNWFVL156/YSQsdg0SoD8ishTdEjwDyZR/
bPbd2skFgDB4RwcGT7qgzqwvX71ekwvYFviXWuXWR3/rwJI8DopCcJDBNTEVFgQQ
Sj+1YDQ+DgalWUC+Bl3rNCuU1eTmhl1AnayblNIo0yp69XOoOiz12723AIN4d5eu
rBU+5cFmoa5IO5XRiRu1VyjHPTi7R101fqOadye7pjim007gSi/Wp/AOGJfLL2CI
qKt2dwvdP+NizbiJ5Tbx8jwZ8NqLnSmgdQA9aN2NzzhghJeE8QEU08iH3X+Q+I42
dxZW73FFh/RFcEpQCtQUUdfAAArSwSyuc3u36eoR+xS22GijXJuS9SP6VOS+39Jo
CG6jN+cVxOhFJPE/2s24VFknpaSd13opPdhODTVxJa5akzyvMd35Fq0xwDqd7kKq
Pr1DFxA7OtJdb1qLgkEisnORpaR/3TFXuNpy1aYJ2jGtoh+k/0Le/vcqBs9nP8XV
lskjZU9kdCN7BHjmMkGcWpSFhqLHa0Upeva8KSA/kspEdJE0h/XvN3sX/tjjTrhQ
8cPd1yIaEPE2KXY6Z+RTk4rkf1PA/WgkcPf9PF9uvAwKq3jSl3lXwuLspPJxrOOB
0AIkGauQfrQEK3S7z18AZdaLozFzUXQW9SvWgiii9DWsZTDvCtH/JPDX+GYTezmU
tIVlXJx712eflGHFphfFSrKGkQwLKrKsH8XVqLjHbMuFtsPRZN35L2H8gIV1I4s+
HAU1Qzym18/RDNS8fdj0mNLwkpxi5bnyZIkW8ffAh7M0ioD7dce8oOjXiSOBr2dW
muHhUEAae/StyPZB/e6MTMkvfHCJwmADfe0yx/dYvS/hUPv1j/3tAZHWSGFzAmcl
RCisaLakBDekKmgcvrGTA8wlPIDh9JVBURVk6+Z2LGaNJXaHyRec1FTuM+mmXcKO
KcCZcj0nnvT3yBXdRvXAOlhMpXKfHivBSc3y2haRY3FRFqsqyHqjm6syqwEGUrCC
idFBIoEZC0ypnXXWVnF+gy1nqHrFNZPRpHvEen0m+C+tsBz1hT39/797zguKc2Fa
rITVVrxNJprKajpv6VvVtbWjmVzSRSbI8jfZ2a3CD8To1Rq5FIJrRs7r2IMIssi4
ydfXUqD1DzfLKPyQCq9DCKMSQ1pJzmR0Q0ag7zeRdxUve3i8X4lVI8mWjiX9CnvF
LrX4WmXGvOoWTBXPGnE9No191hBECjiScpvl1gx8AJusiWn83hNZdAbQmlDCnG/O
PUe6JneTgMQP7mAIbDQM33Czn4qvD4NsVgwo87qG85rf2mHiYjPm4Ppoy5R6/s7E
mKW8asC80utNadxLZeinu/g0syiU+7mUh1S3SiSzJbME7kjWquiEfDSJ6xHaZEs9
+9GQhhMGo/W2iQA3a/1fBm86KgR0D3WOMVG9oe+wHaxRXNGSxf4IWr/54qpPCEVf
ZlNdV8cQPo0JKg/ftsZ1ZioQW7CRSBRoi8OwM83lYhCx1bykJnD2mZIP05cl5pMc
7++g/bnTh/G9uaPfIvlFKutwV/k3GJukw3mGW4bReEwoe9KIVPqsjMjYTjzwNZjM
csMoBoy0ZIxg+U6RPl/2h2frNFos/DYrk1UBe/4nalyfUptEBSMs792B8N254NK0
dAE76pNO3kJMXfShCqaTvWklpobZ9cmQagLsnBPbpS7cJHRL1hk1S/In2V3f9PMe
a0RFzIoYiEd0vCeBHmwKtFV/0a+4+0Z3cIUorvbaTYUwOXLt+P47/VBXkM3WottL
Ptv4HUuk0+P+aGvFi15Wy+rHrTNaDmASJhlX7qcEnDm8R6w/VfXLbnfC0TEO2jkH
flkvJJ+BAJv6G2SNyL5591L1Qaofv33iwnw/uu5JkJO0NqbafbP/zaqOZRi9VvGH
RurzufdnJbqk2BpTCQG/KDsBeU15RG0LFfo3ryJHArEdxwPSF8BOQji7FgVB9UvQ
IJ6ax0cmn6PL1psPwOfNIFOpL/Bfu+Vo8WYMxdDaTQ8gCa4I47a/e7mQdQVbleZc
aEj0AouCKGYKQbiKfZV6RaATinzcbEkzJtuyOEhdY6STnlS4HOC/N4ABJ1sCiYpv
DHcMxVP3XPorVtFY55N0Vb3qjYEeA+cx830WcAV50FpHughaX4rPDwivTXkxkUcl
eNsVL4nZUH0eZVmu9j2aaXpi71ZaqUEwz7EVrQ04OxnkM7JPOLcrVccIR/TOlTH1
KamFD346GuCeIMKsqnsQp75/Sw+sop87qqCxzBrwWcg+jYc19oJzAvGZp4mfokwX
P3AsYzmibSBK7JPYlYN9fybWVEvyofHtbLO4FIIWYFfE+sQ9FtPJyhcfuby3AAfc
unvXpNvSxiqOabCI+mmT2fJx3A46+efA1PuAEriFxajCFf/SsY0HTnkFEe5hZQBi
dTUpJ9nONiqB4st2CSAEv7xw49XLiuZ3is8nrv5vWT5dFjTHVx9cuoAbi1HQiSqA
egCfXlWXCvx1W3VHdUfOrsO0e7jh0r1tPN19L06igtoinGao/9YNjnLna11DsPJw
h9ZTAoVAZu13l/iCUHLPzRPylXkZV2Fx2tjJ84dnU4N8UQkUAM5mwEiINuBy4Glh
cW5I7hkn3buMYIx/8hbgypfVEUCHkpNZkNyArxksZDNVTo4RDH9o3hS1Ivq5UUcs
cxvD92HxXKLy19lTD2O6OB4mRYy/4ull0EfpvMMRjDqWgTfTrmj83NcQ0jHcoLIB
aSmnxZM69mkP34sNtrB3p+OCADK5fxWK1omLov9hOTljJlrLrUTpH+Zo0he8osgB
Juk7G0x/8DIBAvQi2s4G4Y1QPOKnuhHyM2x6/3oYBoFDVh/V1n2SnMZFs0iZghPL
vZQ4UjGAkTg/mPIFBZUr5x6ZeiIbS2ZjHYvnVphLdcOg4s10E64qUX+lEL49R+Gb
IZq/nDwOwsnK1xwI1ZKhEsvP6oQU/pxYd7dqjQLvZaO1ORNp/iyeN+4p57IZ8zHw
yXSWgyWLZNPIHASme5Lus9k+bueA8lPn6ZYZLg/xEbKI4zghpAi+KLy/kGmXAkPf
2sdxb0uTU4qvHEsmgzyCcP4OTKZSUx3dRbWW14x3PjIL0ikFIBJHAtiGLtxANLX5
QTj7UPxLO9EBdlUP+vn5lZG1F0sk0P+rOn3ABGMTUcvS+zZ/MUghiaIQSKHUthgU
1Vhman8ovKs3bsBUV7fsIUFeA/GHFo1vPONq+r+zQu3NySoSJH+Q6eix9L42Tpun
OsI+GsiABUg1Pp9inPVkZz2xFaEUVZPF6dDrlTammIuM7ODNnOykw1NmopDGIkUH
c6hdy/OYA08g7oJrc6ai4ktrGdQLYX+jpSkySS0JYm/Iwh6+fXeUupQzP6yaGQ+l
BdeFZ9EakhFzS9ZKJUY/bIb3Sz/BjKyce4faemey4v0Ux/pC+B/ogEiKYe4kOB7u
F2H9JfElSnh2/1/ZavIz23J7C22ec1BwLGBmgOgkPVp2SPW5n28HpL9P6nDbUkVE
5HPlvvKPrmoWPAd8lkjsMAMMkEn+t/gfhwKkULp2G5zPQhu0HfKKlq36wjeWATi0
BvIlLov949yIXi1GXL87TgzHQ4cxKz54u0/ZfqJYmDWaSedARYrzKvT/CXA9y26s
IcUs2SkHy6rBTluZ4SRkSgJn0vgxxaF3blDep7n2+gX+ZUqLoiD0eYNDh7ukWkLM
sFm1Gj9L1Um87YWH286n/JcA0tZZjTqQY3Iqp7zZgNECJZjXEnlyh96LhemIzmyn
N1I5a7Hfku0nUR8bhq3axy/EyBAzYAs8vQPCdyQCz4qjXQJj4bDIDRGcJMGf0Imz
bCDzkiFqsSt/dKaUhV8kLeYmijPgturpRnM4mSXvTwwiR1RrvvT6N6a/0415fruZ
9tJbbL2MSdGKoYObskC91RuEy5Wets9XCfTKKXZOpqDEu9iGZBeqG3Ndsv4xDVVO
M+KSdab7dIdnvH6oCxdLlZD0Dfnok1D5ZV5+I4bWgldQCX8qnRYTkTzPylXZm6WS
5yuDUIA8gMMKEh7HiVMc2l7HxFSH3gmvO51qFhKua7+623roi4lS1rgslWbkQcFW
VlllCb3Fcr90s05q58bfxVGaH4Jx3KxBHjuGI+EVZ9Jh+eRKcdaHcScg32pqATXV
cCTNDg843CNI4t6cikGPESTRwypfz3UhM0WrmaJg+r+EJdr/xXmL0G8zD1P/vw0I
MtTN4AZLVmEcJIWis7sxaj6hvY9QEsC58QEuejPNbBhIR42UoJg2iSv/1ZYRzYc2
ZrOYkfhkiyuYprYomhyxF3CsrDOolsA7Gz13UqY/+u7YjLVn0go6rbSntUXAtRAa
H1FHNJ4VVlrAQruGtg58T6GHnduDXyhUx2jIchoLUok+eV8owWknCN+6oI2SJ3NS
Qpn1sdEpz3+5PJCZu+NvcgnpbySGzHD7GlnEXJGHkX4UA4Fi8UseVgOlCqCpmMJT
vz3T2WejVyQG+TdM8rkchjrKe6suwUvaWintDznOLh6N45rlxLhQyi+vhVFyR4aR
GgixFUosdkkCtaYaPm/W1+x6t2YdwBGqAXwlnGUM/ilnBmwKqMKntzQ0dnOpzkhY
+x7ihQOXC/Beg8UWjEeJZ6bt0wItO3My4RLcyTESiM7OvJ6nVlTccZ07rriBFNSt
Rim0sbfuJrHLzAxuysJ+YqpJ5aoZb8RWUDD7MqXUUd7dZejlaQmX59HCBon73SUf
2/fegk4V8Nu6YwxIJUwtvSvu/w8xUEqLEgWaDSG+ubamGP5xES53sqLqaEVsgFiL
1AvKj2V3KL/o3ALSZkiSd8U2y+nIj/lK9B6O8D6ZYfwayL9jVcjJdZBOzvPb/0Wk
l+Q10JARG65S1oqtlDvR3XuNiZ2D6jarLifWMf9NYmPAa6MHWlZdzaEAvpiit5ZQ
hEtsUFTzv/pBXYymF8HCaT3N+TXl3oIqJGCHUR1CvOJ1ZB+Me+cSgFJWvIBgvSxf
SC0nuQcPUPmeNOnzDl7nZ1SBVwj8S068Ze2tIXjMsJMEsbCKuColyncTE18q+lKY
`protect END_PROTECTED
