`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCCt9tO2cuw4+DpF2gG+Syo7zzjMgeNGsMreF+yej7KS
WmVPhphY6XUijWP+VL2HiDPQriZa1czXE9rZYJ5OkpGdnOpuseOBwSFI8qnS8NiT
xAF+yw6XbcidIBHWTV8+VqYvABvNH73u9B9uvhty8a/U3Vr86uqTSjLZMAARtWhu
0S6k8ogrkm6uUt/jWyKW8yzeS9+on34cycn9KmX11eVm2nU+8Ac2Uzj5LsJWXLOb
UgTPqJmw8+IwWKWMT9diPO0VftlS+xypTJRvJEgX6pu+9YOIg/PGSyMt1/j5cdeJ
Hfls3yJtMyF4FMiFcMqPbJGfgzTV5ohL7zZ7lqyUfzXhf8AOhu4vAJ09R+EcfvF1
Uq47cyvLC93KqppyQZLVGm2VLRJKuiZ8hN/QHuNVK311lcfOVDwj9AFub6GHLlww
T7xgmcJlrRXtAVFVaMQ8GbBTqzCc9MgLsN7IV3l2Z8sIo+vWpDGxb+UfLMM7E9dm
37+vDNXuPxyt2xjeeBmFcttTa+ZjSynXbDLOQMzt44XLSZUvEMEh/wre3lc74nt4
uL2diaRQ/Satghi/4ygocAojPjpoERS9ipo5aBmYxo2SP/hAF+lvqWFCS2aCpOqb
H9CZt3BYMQwQz+X4QTHSp2A2Bg5swzrRVkFX1jij62j+7MFtWlMOxKRNKqvV39oO
`protect END_PROTECTED
