`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL80cg7ccc7VA0Vfd5V0HbNk9RVdmHCEP6pXL8wQ7fdHx6
OoOBqjNNkuAViVFGr39I7XNFPcnHYhsW1+wJ9+CayEHukFE0Ns+w7Akkv7tTqIVR
FxFqQj4Lg63EBWgCiO2Xc6PUWVSzhziCtJiIaE9fzxs1fjBZuCoY4YiM/Y0w+Sq0
0SXY8dxKSoXgnwpBWAi1TSMDBYBxAZ0TOlOo9aP4HdtRZ3b1QveP9im1iFEcrn+6
+JV1xzvbBQSxtmwZHW9QQtgApPMj/IxjIcoAhq0twn968H0AcCOdnn42tTXiCxaH
K+RA1uNaWF6IzR35nuyEjqV5i7mVFhqXnJdUvqI4lXtm1WUUPykZUmCQTSyaQtSR
DU4TIJMlgx6kuY5EEasq6PszGSWAG6qt//BsaCD2qcmx3qG1Px92YFRbNvQsieyO
9IYXqcuCJeH37eeuo/KuD17OqIzB6CNsh83nmU0KIxsMam6CpIbXeh0Xv8qRvgep
sbFWnW+Om3vdFXHBqMaL+25rMgkQUsd2dXKTtv4X7Vfe5/Up3fPMo7jVoq4kK5AW
4NFAO64GgQcTYMZbulGBjc9wsnuYvV/xhl5+lfjKo+bU92rj8zx9sn2BF07DWw9C
VVwCYRCAfy0HCfHgvHPnVIrDZD34DPkw9Y3ECelZ7bF3ES+vHx/ghCKSD1XywbKm
8zF8A9cvap8X5OlD1G42jBGnjg4VP+cIJSdAf982KrQCdW/rLuZEIF8Q819Mjr49
WSGQ4trvc4ny2Moq6RGVNjYZF7ybJXr2WAX7Ut351aQmXjBT8nrV9Cu+o36hEnfz
IcfzrLK7OMATVVejtoYQPZOsMIYZXLxtSLRCqDhxmUKNOwzNSeaVzB64KQ6kmD5m
iPpcKhgaMF04KJIBiLe2YL1laP+CpfV+qPnAcJ4xDnid3gWBpvnA9qPOd3QEJp/L
OiTkcddXD9tJw26k82PxWTSpqyTNbAM6E5WeUpM/H7kv9TN6AwQj6MzMjSvl/oRZ
+iUpP61oj2Lq+DphTbUooDJ3GW4W1J3DeyOq9Zr6j/EJ1zQ4LodlhPNQ8wDzSRQd
TSKwQHbF8shze1KrIEeLQYM1HHMrjEcfQwPP6F46mz6074wb1p6cwp2oWhGk5TPW
a0bw/p6B6YHF+y0bdN7uzw==
`protect END_PROTECTED
