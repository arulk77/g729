`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
vA2bw0G7sNzIbwOhYLHxmnO2QDBG7Zb5b0PBOmGDJFvx8z2AC7LFc8AaYuOKTKrS
h25Kl5p9z13MKhcrtTA2OjWKrjvlLt3x9Bn+/jBACucQw9a/ZmSslIYVWcnKBjZI
HmTEJfXr9wvNpAzJUKSEAC97neIZ8madYX/n7UmCdZ2WO2R/TUfYbey60o2bY8tO
`protect END_PROTECTED
