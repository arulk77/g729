`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNTPXt1BuSa4OWmBDyTboH/8DmPs4wsLaZz3mFmy66Q6
n188M5VWlsbEkP35NgfLL1B8A7GF+bVoUDLPIGRKW+UaUAQkfEz496mE6CDCkGGT
vAatIwpgfX6j45I/ITywv9INsVLmFdqqHvuKw6rjMehFjmMRQWoalE63DLqwGSQW
1c513byW5J+CZzvNH/y+EB63Nwo+Q53i/3OhDvAllcquV/BexIT9zP4Sd/TQ2V7d
l8VBXlPQZ2+iPbsvDeDKgTUf88XyOXFvTOw3WmR5z73iU7mEqqhaEk9LxarXDkiO
ozhjSbMZhuO+0oYDtOKRB/WPKVsG90UMKVW6HSmAQv4aZP66ORF0rNDltIK0ir68
a3IyUc0yr5ALK1v65TuT5dxbjQNh0OUuLWnBlSNfbmyOskCVnLOpuB31LOXj73Mi
AKneWdQxTbaWxOsO/ZbUMCNGqinzePeULD3hWrDt2xX8qfWbS/c5rAdYPENF4z/O
R4Pqc9D1J4SDsNVDS1ODeEiFfQiXxaSsq1Ry3vUJ+to230IozTLF9DcgGCwNnVw+
n3m2hRYB7O9/WTrhHEtZa+yGeY93uBK+r987lyzmYxMqvLgJ7CG/FVw27cBwPgxV
NyLJXpFl1WzYxSKfr34dPwFVU86YRctOzSxH7QfHDCofQyLnLAKoLfExn+B4mPVM
`protect END_PROTECTED
