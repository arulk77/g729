`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
e2pSC3Zo4uvMUhxtJOIuWu3LOUlqsKJxAo+0hSfVdEZRbIxSPHOQViTVXcM4gX1R
ccrx4D96cDhU9MJjAF0rzq8q2dFYjPVBGYAOP2bIz7v/JsqK4oHoSFxBKPYC3fUm
ct/eCj9iZvLikUzIl+zwlJn8FEzsSz0lL3GHone6jd450QpxA61CReNQ3CZqWVap
zHKwxG8zwA2l95eIjGG8XRY5jjGRfsbgMXXpgu5LE+H//y0oq2c64kdWRjkv/3Rs
AFtmGmcKSMEZ6JUw/Iq5CDr277CApdr8zqoApFLgcXcqdeS5/coq0mlYG+MX4/Yd
iQ3HLY/O9DZo1U5oeGVThSQzL11TQZ0JkQuTv3cFzJcM0Uzvuog+xil18c7tq640
LEQfzyp/qdgSpxoM5sioHXAhnsxJ5ZXjqwzk7qYMSH8/SRbDguTuwO10+xDNnCkK
+Ek7999fxE/oiZKkGL8E4Cuk/LmVfm1dKCdPdAK5cDZ+e+H/7OW4+GytlaZxs3g0
L9pqRTfGQkGWD+vcvK4BexRF3ScGTC4U883ogg9H6hjvBOLt1irjbbnrX7NC9w3W
zXrHaIIIDoFSIyCdhuZ76g==
`protect END_PROTECTED
