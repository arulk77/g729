`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN0Tmp221VXIvsbEgzXJfyg+vmb2MfYyhPUCzDTLH8w0Q
WNpeex1EM6ICl+IBw53FRZrqJOmscgv02z92ngOMrNRYz1KDTc5Vd2caJJgv3aFb
aabwWNaIPV00zLJ6qL+y7P791GhXstVqVqe/Gc655mxAfXMj3kC3Gi9XEMFM8nHd
fWDqT75LS9N+JT8ZwXiMZHtDO9YKGFqVPa+FjNYNF/T2lentCTwT+ksFj1O6qH6D
JyNap/e5cAnrAzCfEFU9ol+IF4WVeDAV+dP8TUL1kfRkEH7nZqDZEAtLkG0bLePN
hmsmZtfGMs3dAtRwLyZa4bQUe4j+gBXNH3qIeUoCfuOyf//d3NrmDzPi6Qn1k8op
sOYJGlodKZEw0+E+hRTzerMpYMSg5fMgHn/NVviABRxfqUEvZb4Auyo4gCnAB0Qi
kEHD0tL68jOn5JuWrnpLi2SctIOHczrR8FxhRGhAnnYvrT4c1qqJOmA5BlU1EnlX
OI4RTeVKrlpbzUecFZBblVl5+7jHJ8QWmGyId+WhpX4L32M26+4eEJUADrH8QVUB
faEgaRNgRhLV+m5GIi65hf2dtf95vD+rw2LmrXIYxmS2Sr72mP19MTz3XcGdU/qQ
CMCtixLk6mETgfmthKqxKwrQ+8T+XWudkkzvxI1AuRmXy1RUupWXCOhwcZmsSzgu
cGTJB9HNwYXKtAIvauhlGfXYWnKs8Z1/o0J1Bnc1eZS3iilqD5ujDFez0NIPWVy3
ZWzIKtykYr5Yfom0YGJ9LouhoqN5RLR9nvk2RiorD2BXw9gVL9ddrHHhgJyVJuh6
Ip3iv9rFCa1dcZF4cmJ+IEh5oQNa/Ad4dClCHXeATHXacO1vRwZdvOJGQLqGLM7C
+i+7IYhrBF1iYoJP/v0UxpIKe2s36kVWuhYLZN8KrcsTHIMSrJjUIo4fJWZH+SoS
VgyTvSwzgBSRBmJRTsLrX8yaA5CrotQrJp79A+cj8+I+kiFGE6O2iQw3wBokLaiB
rDOiDSHbN6IzF380itF13Vbu7BHV7bp0DSg6Vna20P6iPs3un6DytsS24YYzoXSM
UyK+Rk68Jbe/z1RITjhj2bycOg8qakiq+Xgqn6hgLCmraxRaP9cCPhNE3zDILB8r
WjHZFdxG8kqgnUyoET/kYIMYQj9h54U/Mq5Qg9hILqv4tc44fcfEn453zsRLXpRE
Nzj0Fz8tL3d1VWibIOh2FnXnp0XWfg3zaGXB2eeuzNXVRlnpmQAPgSnTs/WY7dDq
fsqAElaI2ClGPrlcfXFxTgy0x6yBliKqeKxjaHElYPqFY+0ODCWZM4ZHJUUq/wD2
bHN1fmkus3JBRTqF+ae5pzdCTqgtv2+vZz/Bv/NMMGCldZ3pHKxJWtjub9of5ezN
wPgmPjalv9lgEKC5deS4uDJJZecPJR1TrfhLksVtFRryrsMQ4rEPkkOwbpZjzeJB
EqhEqPRtP1Z2Xx50/C7p0VMFiIZxuLq4QowiUZCwYNgdCm8L37JwDIakHHo+mt0c
d8YLMfKArnf/pNqVNTTs+Ior96epPUhCBpeODuucju6PP/rnm+yrx0pdkMIJEaoJ
Zi/ui8GCQIHM4jCAw9kz14wfLwrIf4dr+yfaE4lm2A7QNFTJF6nn1PIMVR3b9kbL
V6NRMv85pM0sqprOw3IRusgu0pCODl9OiMOn0sXAOnnF9TFGuJiBeJbt3WaxXYMS
Df3wGFqzrQYT0OpnrGwsZ/QzoSyxlA9SPEm9DG9wKm5HtTH+a8LowsqulnRnG+3T
yyWYlSqxmWyctLD6Yi6b1wJQYH2x7rc25QtIFLeIY/z4bc0Dk2uq6xB4elXNGLSR
OqilwUm2VPdcYhp/TjtQKMz49ngSGwsVHDsgjPdGqwngx4VNOnrRILZ4gJyq16hZ
XkYMOFqKjFA7jtc6+3gFGQwLfY2EMsVFUoiFLxRzRU1+MTmkjSycOWy6VCSqRfgG
7SzGHvSaneiKkVXSauAqq2VeaZ/JSl7EEJ3WmGvC8mXGKN6bwqzpz7thd6oD6Z7x
i6ecEh1LODe+/9n/k/8kKm8yRyWjSgCtg74ban2sv0FYLMtU9+ncRvuKUPIATfuU
I/4l2RBBR4SHpT9dJrN2mT1NVqj2ABc3GahTEnkwmhh2MPALXhcMXKUd0KFR7rCX
UIORaDNajJbP2w5riPIXL65I2egjEB5GgoeJACIIpAMQ7qyUPcyjBe7jcPdaXVv9
Bk6ARKvHX6VfuXPr7BbGMy4HGhjsokIvmJq8m19epfH2RaJqcRUsUkhzaF8q91li
M/bjs5lweflTtrYNRopvMRr/8fC1Acfyzb2lpumsmP3SmgSPk/uQPbidhC5/CBeJ
tlnl3JLHnVciFiwPzwRE0fDZVIGxZjTrDmDfVll+Mb5ttsDjA7CmNIm+PQgSZc+e
LE9ULWw2nA+/dGDrZXgabsDGxVEab4mUOhbTDUAAOnnB9cA6kTujC2xgw332qnej
U6aGHoJTqRPejw+9vrYUzdd8NkADOiX47r/6phx71dE7OlWzXN47sHjCgtvfJQmB
EtC7hEgZAAI3+OprpiB5doJIDIXtWsFLuChrrWXOFIVsgf/165SGEs06veBcSIX2
D0JxpQKpibyYJO7XNIAyr5nuo/yaRsxmXmLR69w/iQFFZCorAjYatVHdow95FzXE
T1dSiWe5pPkuFtzhBRjC7XmvOpGu9JrbJcrO8UyK4Xzxmi5slukjJlV4FUYOH024
DdTY/U7l3RfrPfcIs/wsMDJCFNbY0+GoyPwD+PGALmW/4FZijpEyHjuJj9HkeBKw
jEuD7NYi1xwZqpB39wjxShb+RX8hWWKCvhXfXePvyUcmZVO/ZWMIgKsyqbeLovlg
6IQ+My/DIPawT2/nAN2R8j/2vBx7valDVwZEnPtTdBSmaVo+3ajqKiy+MVH3OCBw
BvrKk+FUkddW9WpnJAk2pnjeUq5qj7mRhHKt6covF8YcCZrJFBuCrFB1L9x/YlXL
`protect END_PROTECTED
