`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePQiJ+DAEV8u1in3bw8nSJr8pxQQfwz4OWjnYpAxHce+
NxkpdY8O6IbmfEn5RCpS/fJ0oiewPGe3GyGuBMLpcTY5B7qGjlJ8LVdsRfHWREbY
MPIZYOFR4JGV6cSQTxhybI0N9r07s9zlC3uznLkjpYeYESf0uRfDRpLOq15KcGOm
UvXwvHju0syl0FcQqtxb321Shoi+LstXd7ZhYc3YukIFkKNfl+hBgmiViB+DMCiU
lxaAfY0f2WJj4swUjP8sRIdSsapC0+HrxfhI85eG0cIqSLvQsbyi8pgtYm9+3ppL
LdZmoR7o9/5rK/bwI7QWbmB0P0vMDLhKdjFbV1sItEmTRnb5rMCeAn8126gEU3t8
nVqoCjj/b2oYFAAD4wo+1Qs5+PE8s8wVzB9WMW3X5nwfPqy4MYaU6FpCTlUzf0q+
JWZci8+qfPn2vemCHWG+8ZEuVeHFy8l+Mg/Ctl5nEb5Q6N3yKKH24TQJXCqSPNnb
a7EC9xUVdW3cz3ZazGG/BQmGX3HNvbeeSxz44YcXj/pS8gSbAbhNI+IGBpORwT7a
80i9nHnGFA4vjs5kDe7uGW5ibH2DqKOBcNoJxxGkowiOLMOWbLas/HPWSv+YBFx3
6j7X0XRWIUCXui6SuF4yE4RsbyH/Ic7vavh0YuBAR+1l01pLeYllvOLWe54cUJoW
TgG7Sd3ss5NlPoArJNFGLPQ1AEz4U5/JwYEdvOy45rJv6cyZ6WXE7d0hxPW8VA32
XDs8OZpMk/8OFwh3adezQ1kY29bdBvt+SK4ukfCOIFtoa3axCs8yuj+9RVZ6cd9v
lNu6N0FD9TgK/nuZdqOISw==
`protect END_PROTECTED
