`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNxZKZaJFMa3CmbKWZqGBkiF8vH5V+9nxRaRJgbqXWght
Fxqu/eN+piJSSG8ALSDngS1VwI70N4gybDVfyg9UX7TRawSbOB1+eLyLB8ehNIQP
DjjU2xLLnqtn1HJaEKfd73CMq3yu6y0FVjgOSi7bcUyYEpcxXKycfUXftXo/Z1qB
ZOr5pJUEoW3nXAa4li5sdq+A2HcIgHYSCZj+X/mYPrqsIm1JYTrkWFbZRg/FasMQ
UEpMLHIXpeNzxjhqQJG8JCRlUFhaRefkpv8NccdUqaBz0+rv0UHF7YYMbthfR8Xw
oDtVd8lD5BLQtQhhyoecjTZ13nS9FVS79h4VGdGddxqt0OOq4Ywiqis8V/T9as7T
3UY2M1GSpknno+qUuhTh/w9o8qD5Q1Odp6Tl/Gm7p9tRgwW+hwapk8wG1efY2YKW
rs9EiqDqlTWMcWRbWQHnKPa4Y7HbuqklscGY1Q3hvZLQcR016x6cUUeVHOQP/3r4
2Az4u6ZcPG8pFwj0GIh7sFhwujVHt5OdaVrjgY36GC/anLHPMKH52h92d/hYJHkd
4W54aC47CwsdwgYbzjI+F9qXVTmQEzzJiGpBguyo91DigkqNNnHnKqOT78Au/z8y
DrncsX5LynLEBEKKcGkWovp+gtGOR1YZ0LHGFf5X/3jjRiM6eQxGA5ru4kg5a3cN
MalZSjwYaM+C/unDL6baZIQoAAO9/h9/HRb5ECwGD99+GSQ3MmLxE7zN7DBL+FbP
ICNXQ44FDzESVciCgjpHztkpJm3XAWDY6WPrWZ3JHmLSFDIFYpIZGJ4p/9Pd/jNR
xag/rhcn5pVMrBmokvSLM99i5W4GupN9sPZ0JImysYeN+2ySYrG8mKqiyxjo0Xb8
U8x1JerkpF2cJkk5KlhfsXKmTwR7gNiBrR7i/nmFM/LsSbhdKvuFiAxME9OgJcFc
cFNJTHPkQ6dJFgbHGSwOyzBo3dmaUeqsViUDP25nBa9Jx4EzXf5Zw2/2b/3eoc0w
mzp/uhHLVqbpcnc/VpgbBUrx+5YAbRXKqcEQ0tH3YTqX4JpIJVRYd5DUV6C/2FOB
WeG7+XT/8wbz3cwO+u+c6TCd4M3LwtplAsHqnbBJl4E8txjRi8Kxr066RnHUtPj4
zjpLWquKMBzpJKjSb+Cp8dEEe/+AZAFUoTomyNL3InrrbCb8hwM8PvHK8XWGHpgB
W3aVm2GwJY40RZW3ZelDJxff7uamSKO1AmT9KTDtow4OX5GMVyYT7Ks6YNYbE1qV
HVcW21YNiaeSVHzO3IlEZKeuu2uvUlagtPACmiyLTfKCB1mrYN3SXsDonqDky0ey
4IUGCxBeu+Pg1tJEO/jC0sy9yEITj+/ca4wTFJGVeoIfbInbZelhx31RNbU/Bh7Z
FUbzDNbEuT7FTrOdo7/71VQ49njy36OhGQTJHV5BrjGzAw+c3RzfbiY6q3EgkEZ0
aVChH/m2LZ1TDSl2GPfZFa4LROrOdIsaPYVtQSJijeIVVzdlHWBJRGD/BaruKfbP
Vn5SfBO3sSuWlin80WS2qXPMyr64DUFTL6hOy0YSt9/ipPPWW8XqCnEUdnfvUUWp
UwS74qC5psZPglV3D6W12J2WWpsXfRr2hjEx9pDrWsRai02ODAW9kZo+WyMHIh03
jpPZyqRoih2r40WVNQKLhVRQjLR3st8LECaJKsWsJg3b9m4xAvoxNBQeuaYtkWA+
6wUs3gGPEUFVFM2dWYA4ho26dWnX+609A0r8ySnegTcelkfP1figWD/GoKuorBh/
iWfFPPvt+2QpTdqxF+XyB2SwRpy5GNXRL9bysBUc3hYjkQGo4ITTgyXotV2+gDv4
cv/bbBUU6ubPalArQvkDMfT35utk5jlP+pAYrbqp2Yj84rLGo+pG5k4k0nsPecys
QmIfyaeRu8JxyAW/xHUQafmWxupBHfguMW7oElRfRDs+16z6Ne2kN0If/xT74tP9
IsOd1GWuG+INIm/AAIZj2LMuBwjNiH4aZE7V28aJYo7g5LE1oigDAZDLLd+8yNWK
1SE0eNGGLP39SwoM7tLYQN/TMoQuN16Nd8gv/VV0NncZknYeuCH+/lbkhLAfQMda
eQlzAbw7ekMMFK5y7PJlkv8WVsA+rLWegUAbGZ8ccy1GWCwhkcQe6qWnmGD9h3+0
rEcftjGfzndHr0WaI1gX1ocorUbdp8CZFhw0RpBga/u7wVYHqx+lRMET0kqI4YuK
oT+NYG9EEGMnwoqwp75sn38Dg6szgJ1/uGF+nTePF+4EymKey/0R1k7IB1xUuk2n
fZ9N5O51KcBRuBnSdshpXGFRu5mrPMZsn2R38fMi0IC2HL/g5AACrn2Ql3Wv7cy2
N9IXaLtI526RGwfgDh4NiEblOL3D962uf8Ifc5qVkDuYoYJsmJ1MsZxu3WzbrhNg
sCKkBUNthb0LdpKP2reIUIgkGcjeuvQYyH4Amaf9dnhwoBF2Lk9fjVxv0X/+6O8C
BLIMzN/vjpCwZ5QbZFzVCgbvR5LM2uERygugSmjo5WoHKxQ+LeeKYJHRl2GmlwtI
2dVceCkQV1qT+7edomA1Xy+dNTWQAPErpl93ZEMhxc+XK4qGu6LsOVF/0AEshuqk
xLixxPki0q19BIMP8zYdaTXKYLnJ6oTQIJMCjIuw3cpA2u4wa+qpdJxb/4swar8j
GVwDPu1NAvDtkdlbN5B+bxwm4q38/vBXmH0BPbjeru+2mfKN3zGU/+iwMpWC1czg
VdckLsL7RT7ah3JP2bQAQgXnw6kFOnJuQae0CHhB02/YgUtTR3SAKFpSNAHWmxeZ
+DNT33Xc7nkXLiuIi/1hauXMiIIRJfOq/5enkhI7UoglPbDr4WFnmGq5jjx6NDhf
kMBwXP+8gQml1AsxjpS8sjpSuJ8nTIvs8syLl0o7Z5qJswT/Y+FTpkKf2yS2XloB
R+0nbOgb2OcBq55Y1e8/1OK7/wqGKeJFLcsba7kZwOK6WJxR5QAFK/UNgggs5ryb
89/KaloZFn7Icvp4iifuH+3G0ZsyTmWzKtGyR2qihSJWMOTCrA/Vgf8CfLhQGcQa
anofoahPempbxRPnWWzGXqO7J42B3Meow1UHz/dMASzsmhL9vfx4EyboQ435mEhU
mmJQjkv5j0ohYSZ7/7maUzXBjZKnR3r5XO/K6KLVcSlsu+6movUt0B9w22Lr2Ekb
yCsoqmDr8qxVHvtylAsEqKhwzffjdz9Y1Zfj5FjX+GY=
`protect END_PROTECTED
