`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAU44SkqKIwVqDuUbkkCoLrEa/EsL5a00o2qDpMknWvh
RWriKt3eg5GxesNnH9EA0GWYZbRDwnmC9CXtrkQtvxCkqTQvAy/uTJ9cyotO9eNW
yI2Pr3DKdjJkb150Bf9D+t1o3zzJqSFgzkdoBGBl7+kYnj2CddGr/0B2k5lbVhUZ
kH2QA0HQ/fnr4vDnAmTSs52TK2M1jiOAwH0Lb5xmFtdTXreQNlhUqyojKnfLe1Hv
`protect END_PROTECTED
