`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+/CrJ4VLaaSm6uTqSTf353SVORMBeD/6++S0ZI9c36y
8KiY2Vj7PO5YlMDasEajsnH1oFmoYQxP+V+D3RMSJ8V8Qp3bemRhUrto9MrSeZJa
Yo3jjmvsgI8xebU7aHVVfcNqV+zhG47PpvUIqJvwSQC1MFASZriczkWTYe/EMNwR
U0c3mefns4WhAzzMJWpnJ7gEKsR8Qz+QNfGEp19EWJ4IjBLQaWCjigobgzKZL8Sb
hy3RmlRjuxL0HjsTAPBzpwx5iQdnOJ7nWkq/uo5eRTflG4c70KbZCci7XP8UlH+Q
IZguZKb+pW7qi2E4CQDSvg==
`protect END_PROTECTED
