`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMAm1Pzvw5rzB45/szG3RzcsV+xn+0cSBSNBIrdDdyFm
ZFM0ouDuo4iAtY4a+hA8OqIsgQBOYktI7c6XVx+Y+ynMEDZbGWnk4fP8Y/abMfx7
zJzLV3cYE+UjyMJGssLCBAMKke0qfjb5MmDvEcgZPwBzu0PBFYA7FDr7WDvZXt9O
P//lLmckgpqst55FAQV5jSgGXddym6KvynoJJOwphAwm3gPxbUdlVw6CgDO/BKPH
MJYizhaTDWLr2Ecje51QAO8sItrzJij9L3ST2CfEic/aSCbmXpdZtpnVrO+kt96R
qTpS+jKRPinV0ncwnl0CODbo1jAdtZZHA6wOeq0Ve5ZdJeWJfbhmvNd8V+oFWIic
bIw6uV9HbedJ0nYmKfA/wZqHI7fMx/NA8nAdqEcvKGpzbsPf9lDDO1oWwUg313ry
zAP4s1rxlkPpDM9BxeZsxbAc/K+6vNNse17JSlxUVTb/DvHh0pbZx4qrc2uxiVoW
bX5eRh8ILOc6/+11I5+TCAQOJ61TJeNUKBOh9uGQMB6HNEFIPMps2bfnZOdb3XgO
iYVLSYpcJ0lIz4UQbABnYeeMfTmNzt7hQWmuoyAEO+Tem2Y90z+bToJ5w/gmocPS
XAVT/popKFGUfBVr1m0DU20ACPEtZLmXZmzJvRdkpGr1njyfUcywBD3Wh7gCWXud
`protect END_PROTECTED
