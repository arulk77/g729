`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
CXDo269tkFVLssJhCUcbkcERvk8KZYNGzTiWZTusvAho/lFyFtqVtOgqyqx7U82A
/ypzr2LKt/tKFAV40gOim0ZPuS0dDRtA8lfjOVFi6jMovYfJA3hyylbSnGhR+/Zl
Qj7eYDMZs8MdHJI/eZWvuzbPeh+n8gPz/7fYTDvn+4r7S2J0iqxzxAlXbFRNOp+q
`protect END_PROTECTED
