`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1adrsQW1yp24PxVlPy2x64P41w46x8r4KCnMGkfHC4EV7
0dGNybpbg0tebryAnie22o13GU89LpZSUw8WODxMM4VYOyd7Giz/XAx+3uP/SGFt
9TadHlZli46+d4CjK1oKdVlK1cgifz0DYG3M1iVsnH20Fj9TvgNaIAx1+1rSq7sB
f+E8uFFeYbTpKuQEIOBnGLKgH3JJRoyjMrv5dVg/oprPqjaqVRLne+qe/0ZLirDh
`protect END_PROTECTED
