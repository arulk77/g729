`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIECeVQHVEZ1/y+hv3syvRGOLXQKPWmdnux3OveVeYwB
Qix5ZbPxurZULYKD1lLQ36P1DgKfB18+tNXGM2A40jdx76n0ML3MqY60jf5l7K6z
Dgmj7ZI8b9G/ndtbQT5vi4eckl5834+B22GbkvyocdO0KiX6GNDw7YsjzcH39WDh
9ZpXImElp8HPZeePPHqJtg==
`protect END_PROTECTED
