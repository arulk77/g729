`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ5y4VBoUqiFfMJKqutjs2Ea15ODJF3vw6D4uHVN/YG1
nAUzQroYnrOahGxWl4KXjFkgfgVSI7+/mR7O+IK1EcTZOl7e41PqFrlQuPCqe06z
YZ2bVifrTpuh6ADY72HmMuffPzrrM5mUuV9QWor2xy73i/UBRpQ0LvHozyhl16Oh
NpfOhYoKDhDrbOC/a9KKPG8cfPKpSNawhxONnPTrvAewJsKTQxHhIASfZemYRcji
3uLkbYhyXYEoMoULczl7daPvr1HyeMPDEPo6qv17VjBLlXBezeXZD8Uu6zHtLLjD
zcVMk1F0uPKp4J93JZGu2NHZ2Zb4ZPseEpJyLHDn1TaCDZpS+e/o4FhRqrw4+cDq
1YmN37bp1A332M4JnoW6UQ==
`protect END_PROTECTED
