`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDPLoCMeGJoZPHSOwhHRtvs2BuGuBBzttzhaq+/oL4Dv
yWgBMnW2VmVGqIw94/wCAD4RGShFESStGRMtfIuR+AeHDua3wKDZBir01ZURj446
ymGS/TKsTvm4zEE+uQHVYeMU8PSzhzaK7YgxQwgLSd5hvYdwQwvEC/juem/rMUVj
hfAuIBW4oVoJYEpsZEzDVtFiMutHFqrLFDRhJpHVVEa2Uj5EfTdGuglAVwbKjbiW
KN8ukv7BhJl4zYjBnyoF3wW6AhCdR3SaBHTvLN36WygVn56J+niemro/FRd96FKp
TnK70AwwayMdHvVsk0OiOTKTdYfdBcL7/74m/APfyLxY/OuYxZDumzERkAW6otho
iAA0XxiLvXYXC/jKvU/OY7BjHbMU18Fs7rFz9PFNUBF7/QKUr7OPQqif730Ljbx4
48TxzyS6Mt8HMSp/9fqKCw==
`protect END_PROTECTED
