`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN1VYKqlPRNqLJxPSVtbemCCUDlX3wmweDsagzjZ0y93G
V04gmWUq5Yl0ma9JhsmO+ZkqIpQeJJ4Z9kKU3FfR0DTG5CW2rlK/rWmBlbr5iLeO
LXXgC9OTuFdLC9kGpnwnL5bq7AgYTvjVfNn4bCEAddlPz9hWWuBzgOLqdhzhOLRi
TGiUKfoyv4rQACeH7dGzTxWSxvR7PZ/EWBGvFwJbvf+QuRf/4TMVC3bC6cl4MFDG
rg52uspw8XhK34RRjJfAcq2x7pBKQj5B1dEvnMi84ZjO5tyAmotV+AW3f6RMyhd4
AY2YXa0O8/J0jxqLANks1KtI56esr9gURcZ/dBU8t6mbpo1T9G5DAAXFDKkULb2i
LNxTNbRYtkx/Lq2z+rl3axreAjcj+ciZditAVdV8QFqewY6kmrRuRBN/GteJrnlo
wWDgYXdgXTnTdCVT8GxY6Bqj0impo16VGGP8yYtJr8h6vZGIvGvCYkODeTqz1ZHu
`protect END_PROTECTED
