`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47feZ7G0qXcTAaxGwU9jah+YxXFRN+AnamumVfl/nup4
3Qf2Mp73RiDEWo9qtxCEHpVL8UdpZ5obM0XAXsAB8AOaNuWw/KdNWxN0OAQEgY1s
ZaeEelMQiJSP3FmvfuRA6lvnD//7t5b8n6L3qUpuNK1c85QlTeC3tnk2T9iS9vjU
TY0UEGtH8s9+DtFAJ2PbHtMRjA7Tw6pdhpuB/CccXAQ=
`protect END_PROTECTED
