`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIK/ue5rCNl1ItxG4vpU+cukQFRzIiFBKOPIv4BzW0t4
fboHroGt9zZEOvBXy3WBX0v7eQCYIRqr0Lv1L1nhP2PCRoZhUi/0mWnq/0s1+25i
BBqnZqF0GN5DJr7+ykky453or5rQD52S3wbypV7UFJxp6hsIwKfT8CzSkmcSRtFx
RX+AZLZ5+4QNlg0f5iXre9PiHCtM/y2TxqBYeApbdzHF1LCFrP35hsPmlvLl0Q6s
2GcdxeRWGPGs3vPILA59oK3iOWlDzIVPW61wZdaZ85YFF9KW3FZtSxxLHSj8Ieh5
pNUS6wwADI1i3TMY4+6mcKLPB6xl3zxhhvCS/Uw8wqelOJ6yzva0UzdpfZj1UZG1
`protect END_PROTECTED
