`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN/hdiXzPnkg4/zPu+NXNI2V4FAtgYscBKsiTHvrqoHE8
LRzr+GtdWCvIoWWYt3jm3BZkffsWW503TK5DR/zUtOSFRbSaEV0p+2xTicUY+Tz5
0lCXdiWInzrr8aI+fysOCuVaV1zSX4kvAa+gYjgGM1KSczElQKf+CAH0bDhDrvoI
FMfhvKG4QWqSBGTQCBVzrwP2cMvM8+fQCCJDGVrQ7cO5009CA3U3jl7WzR/FsJJT
muJk4RqsRA1TLbYUfIkRwVmbRwWGg4HeQKLJaojaPS24ZbOqWTsgNPXirkdZbrP9
byA02Gig3l8acARhry4kA+U6D6ZQr/1leaxuPROuqkEbwsqUk9u7oWsfMUQG3FHx
yZ19frkiKRsougwBosZwEnPK+UtjCAoXvPADN27MIux18rPojQDtY257l2S0n+k1
qxOvxg5s7hVAcV2nXhjsS1pHiCdfo0+vnjeAVx8HZVhetXxtFFMbcXPa/ZwMhRmj
e/SA5F9PYuJXXR9x6d0AD5s1b6n0M1+nFgUwl3D6GdlyE9Rkrok/rIt81Q0cldoV
c5lV0X45rxd2klNTiur2lqDqPeyNpnP52PD1RxDYypD7j9i0YvTVegHH+suZCwM9
k2H50DWRtT2bSWAK65omJ39imsBzRfIaj0Sm9EdrcI5w5rEAWtnlSue+rUsBcKoR
WRbSH1NXNginRt1OpO+XBOo0K8TgKnGWR9Z4QZG8G0WdrNd+/8NBYJuioec0g+2o
TBuHjevkUgBhnTZfJFrcSNzxnjFTai6qqAW1RELrEhRdkOWQPabB3ruFDVqRbc6X
26/DN5eNqX8w0zW442G1DiAW+kYUCvf33v7GhtMYZfzy+FG9k454VSfrfOg5yRoE
bJquEcMO7eEPKyy/y0fO14vR9A0ag5//o4LhK1qiHlgJIDFovES4viazd7V+Ge4E
MN2lphX7Pc65mejlWct1FwcOsYw97FhE2lfgkwO2tUDzAw0S0ZU5Xd5mpN0yTmRv
FqlcFbyijd1hT3/q6hq5qrQnIhfitnVKltq7dGJzt2bdJuYMiBsBiYbemQThTfmv
umynOXIhq5jkN8Axck1teMdTnllgvWeKySYjunGEqYpKcvm3nBj7zey/z+ha7mDX
KMs2ID/TFtkciBN1+AhUO9QA5w04ImcIDGTaI0XFFqQdci/nxJWmjMptYiwlbk62
AKkvYDhFyiuw8F1UYNQ9ZJ3d3z3j6SchVBHGdTdSxJGcnFtZtOMWbzS9T9fcTGSv
ktDmr4UQOtKemEmFyZCMIKoMWgt9cGdaqqKETIP388EZBNJxxgqgmh7ynM3QnCDT
y8XuOmysrPOmQHPbNovpr3LKsntKb6AhVVY60MowCTmFrgnjnfPL13qfxDFFaYPO
JRHqjWfQVPSkTWPULU+hzrrwf/IyKksZkxuEUn1Wb1Cln9Xq5MFsCiAYdjCf4OCv
qTVvS7ixceFrBS/KP5CNm2q+nyXwbWsRo8mOZKOL1h057fB30fbgcjxqkafqK9Ok
7nmUevKi/jmULLH6lUtESD9opNaRU9sspbdAA3VyCTc954TTli1FfVIHCWCnOzAa
cCtpyAZBC5WOkarc/60yKX7ejN+r7FBcLgMwAPpUgN7PjwsSj18D7Ld7z0TuHZ82
CrTojN2nRZqoPJdek3NJZf3fR1ENeF+dPhIdYG55Evvo6UlejxiBb5HibhhZLWIC
1OM4aWSIqURI/zdne6mQKnYEH5w+XpsanT5xn6TOABNvfvZNt6/sU7yVBOHBcRD8
6jtOTpPMaBw/1XZcHo2g6RkCStHrAMCZPcuY+sky8b87TM02aISqQcHu8dV0O7yb
6W0+I3OFxljioAV+wZjRV9gUebxQWFxmINekGs0i7GgEqtpmIBQy2j6xZYlb+WCB
t6pzXYWHyQYKx8AcsAbl4Uc5c1czsPhQvGoYV38w+ArZ/q1eSlYEZXs2BWgLYju+
kZxqDwBTqvkxpe7r/l54wXjocx3I4um2Bl0Ypkg/wJ7go0l7VzjLfTt0K9g6mzgX
UM2DtviTuxUXe0cCMyiy7+sAcuoHWHZ+5mOXz8JmvvN8WBYZvDhuMGvuXZYwkAXB
WLjPC9iFMIs4f8+hk3aMcZGyr2zv6Wt9U++Uzi6bwUmxM07RzqN6TL9DzdYIRuDU
TTaNPBYfD+LFQYIi6xwu6Cze/YMCfgNdtOCOG0Bf9aK+vlocRW7b3Js5KDsnJhcS
/m7o1mAEY7nlJDC1RzXwx6WPsXKvc+JFwtQApON6arGw/n7scL1bjlViLt31SWKy
cXYgbFeArjB1ofPeifTx5tUtkfISUawWceJByPG7X94AHuJve6a3+cRFj/QOvcDn
QpVhzSQKVSOFQmZ8yjMrWzPWzfzM47E9Ynsi7WEAYlPX4wZ6T8sSkN90lfoEANky
8nFILHkHeN4Sjj+Ty9tY82Q+newe7RLamkhM5ULBK1TNJ3+B2z+QJzFaNwF6QHoh
IJLkEps3Lpw1pfnLQ8AKuj/fWxaKcr3j6wPMN+nnBYLYv3JvwMDd7JrOIN3Lebtk
P7Zu2oPySA2/NlIaOp0QsoeTV0ncfUKfzPMKfbWxB4EtYSDC+l/9HMGLdv0inb55
FMDxInpgzzy8tAVNSlV1ecv7AbUK4Ldw6JnORvX//A9WnDbET5HTXrBp+COMjkaT
rwP4+KcLg3TAhBZqLwUL6f8Jnq4MOFT2bojZF5/LhubXfmdeQhKU2+kvMtjmnPUZ
DMa9hGj8KBWCXsZF2joirDlegtMQFyBnUetxK6R96Yi4q3YHZA4jZwokPKRBvHPE
ZjO2j/KJLcIpZHaZsWGBxcKZ3AKlsYH7dwq6Yoa3RU5kOD7BVnTgpidS4r5AqbNe
bFgGcrimFcwHirsExl1J/GB2tDRbD28dmC20t5YxA0duWnUiMFfcRRvDD432e765
OEAuokBPajh6qguuS07VUQlc8JLTBu793Qw9LMWFCDxJp2FdoyOEiCkzBiMD5ZTi
J6iSul8FOo5OcRO4cR6Ac2Ie/3sB08+vgkNUoHHPN3hv34QMu2py5RDPtCO6AEt9
CDeVtckg0jr32y+ZMLGvlRxDz214wcAwcWqIXJ7YfBJQs++fWFyfBLVDclA/+KQ0
6SUnMOyLLTCpBVuSbu1Rq0cXSMgvKwJo70pKGShcUgvtRa61KF03MlGC6H032V7V
PXHu5E7ZEAPMOC7UmjIN/VTLdJSpb5sAhzRjJ5N/ce3E5X4NR7qOavBIUoJe05xB
TY2Mtja7O1eahZPQszyhyImW7e0seWKhHrIn/6g2MJNx9399ecpvDihkkLbS8dQ9
312PV7w1onRwrmW+Vut2s16BPqFfiJtujiLQCKAQ3VV5bZkBqtYPbvx94/iNVws/
ApPmJ9NxCW/eJdqIyizIJ+4ykKzSLyB0q2axMWc2fCUAzrhfF9fVJUbMFK9cBXyw
+pM30lMn25lKMoa3m93c9bISG7zYvER7WItpPhaSK/PnJ8hptroNqD4ObOiULqj7
84NxB/mS9ufa+PIJP+arONtTsyvlLaDPcXn1Pk//pmkk5RTgIgwNoHmdV43wJmPc
kZjr27KPGAl/5IdFDI/8fZL1ZRW4eQgpJrOjkzpjnZsIH3JQccJ//r5nPXWJHlnt
7ORjbCKC2iIfWl5R224u/aT9gJSWHbxGcOq2RblvXBY7lqY29k3cD5I6S6I8Xzti
fFnWIEYKDvE87xpqN4lIngC0UzS2uUiWo7zqVkFsoNUJ3WOAQrC7lERb+k1pl8r6
CoQWN7FyBm8p2F835PxKtleW99oe1KSPuklRPw8oUw9f9atNJiDcGx+DqDPfTM4p
QU55DAm/opKbpmahkwAAiUczgd+zfim2/ZXXsZkJqIfJ4RIl/pqrClLkyZYnjsbJ
lLoGGbTh8304XZaxRSu90l5FVX/yrFmt4P6ODiIWqsPAyKCHCXDjeF2l86hmoTB0
JYGTjSHQrlG6XTgvS2e108hRZZjdh5S3CxAd1aw6zqkLWMnVXoNmmcaQXB+3WELW
dSntq18Fkl/hcCf318vuuHZ6XFim+hq/zuJwdXo3XjS/lFfwJL8IW7iozc1nmrLE
k0ypgdArO+6+5/GsCVkRqKTjdkElgI2SYv8IPiCVe7IYKwvX15G472iYGzhOEEjZ
xzww8+u4qK05URUWcp+kFNxKOvpE5uRALvwyypsBsRHvYgmKKQondbeLLRM41ygj
3twOzd8l4l/x8aJJJWhFjFHUI6ccmia7fBa+HeKakinmIyoOsWPHH3/wssSfMj0k
ws2qUBPmxBjyXveMGkBxA4clYovUjG47whWbXcYwsQ31spI1pEzmIwX8+Vunnop8
Ih14r6nbODZhAOkJjAHjyvoxbWeLY1H3ec3JMv9C9oRs3ZTZOwjqp3osFsRXk1AO
8d0+aRklBG60H7AtCIEa+Zt2BQiVVRkSt+pLJ8CQcJkelYu1NWoAyZ/jum61H3dh
XGWAA1cJgrjizUeoitu7BMgDOgsJ6OlMnhjq6ahimymHGH9hzLTR2VV4SIGojwoV
hR1xh0gX0z0rxuCVdxACEXivrgjAVqHR4KQW/kFUsOmyTi8yHD1Ynlo9EqVvXGHP
z1w5Y6bi8XRQsG+VL60xvleHeCp3FLK7G8X82z660KFcy6h4PZkTZpfsVU2p0Rp4
2TsYoeQsjw088j5LW4QDdPiHxCFqPrCjWir7haThNXTmcjkHM2lVdUEn2l6ticiO
H9cfj2M1lXf+lnHBzgWRgSLorRhCgbQHqIkIqrnS0ve9t7aOAe6glaT9d3AxkBjp
ToqwpOAH8t5JuOYS2C731xrLiRQaWHAOPWyLr+cCn1dGSF1yPOxMaLnf1tw+Hvs1
CFnp4p1m4nAsLfVq+aSy4WKVF72NvW4o9na5uF2MNA91EibU1fS15BIRpbHIkW7v
5N3aSWpLBJuxbDt9UHuVLmkDQ/PfdmTo5B42vwaaay1O/MK1gqZhEFDz4EqcngyC
oefj3efzRB9yjqsvB+d76bVY/QlxsB/SAdJc6VDEAfA9jCCq/aWo9BUG2S5ncmT4
CoSEhiQn86FvF+M7wSz7OHmdgDODxu2IlXql7F+lv5PEMrQrdA1lDhq9QNx2qHU2
lmTu/kWRbWQtpEULc81ZfdR2VcwI201khH5ia6LfCks1mMa3u/5DlRo+sraWHLrZ
44jY+qFEDhsNAoHHtxO21hGSq9jfN0/6+zjA8lIjx4DRjQzsdvoewHytM/0oQyuC
x+od/f0z4KySXixxstbfPNgxY3HQvSaqjBMK4FhRKAFHB+SYaGzW5sG9v75kn8I5
owC3RH0k0dJcUYdoiGzXhDxCISzfJcc02+xDmoUtG++NDRJzD7rHy7IjWGVIGVkn
M1AIw5OksEmt6vcmNOdKw5UGghlR5yZR7fJrOHZRqPM9w63dqq2fEQg+ZJ/98SaL
wjHpjdj4IXtfj0siDg+lIHKJqDulV9l9IPJ6HG4i8sLxtL1Espov98a0LbKtBTD9
Rb9kWJFTl2+Hv9H+TTYcByObXBrulCnPnEv1W/i5N2cN/srDBuBIY2o4Ri/dEnuq
RTQKDbm1uhSQgwwAHXX6Fcvut/1+cYDF7ir/yxW/7NAZcbPK+tO+Byira0Dur3jI
rJxDaVqd5SueHuPQpZKOM9/7VGTgvc4tYs5HyZJ+UxdxdthwDSADDDDSG1BCifd3
gYMPmkYoLKx5U256uhrdf6mNmoTsTpUxXaDOVvsxC+N9jsTtFbw5d5WR0pi3g2Vl
g2VLY2HrbTjiMXm5COMFaTlemALdbLJ2ELu+fe1G7a9aVy7q8bnrosRxClz8uIh6
O1qdcVNCkjorBYhCcmSuz0WPzoV6mAfDdUUnHHqOIvPu4Nv4LDriyKs1geYcyN/7
dQRX9gXki7s2vBhuyMzYszSEpAJgp7rJeorXOJngM/Nj88UPIygl4Kq03Xpc5T6h
7Zpj5Ygn48GQgxuadbkR8hVN5svU9zzEKZZE3sbfR6Q0JRD4KcXpgiEkj0qb9IeK
Ql+r+HBTn1WnwmPHf3v/7MndDO+ZbgnMClMJvomKGqpYWvrftKCEmkorSHAGkOpB
br8YmeKcJ7fgpXZeTf+K9GyTOU9bO8OmWMyU8sCl5Bp+ykEu98jdJn3PhcErAuNW
IXtaeIQ/Elg5psChGeC/wX8mRGPfH49wx60Yk40WzqkmzKXOeD1wFrGKjg2SrZxA
uLfsj0PnpeGQSOQyI38r1GDkV2LKd2voOIJZ7xwFSM6C1rjoQE+qWSDvxxmFA7nB
CLonjpFjfucrQTiTlx3k8SCK6gW9cKuAnD+cabMfqw0vdWXVLskavALXJa33SxCg
mfSPUmwxVOONMuyE82rBkmUC5yzPB6YaNuoJMXa+IsEJuZ6LwZbSPK6Sf+GZ+4Fi
TulWUEN9RyWtRMBKDiZQ+n9CDPPLnzy7JwIjbx4El+3d6B3WIcdyL4JfZo36G98t
bfPGH+XQKmlylN8N9dLkpq7czdNaMwtPAeDxR88eeNALmcQViZcNq9SYvGaMsRBy
RImAiMduTePI/jKrYmrn5x5afsfNljWd3ksPkBky9y9Dnj1WCZFMoJML3hDAzn/V
yczoe1kNemOw6WU91O6yL26fcSx+hzpQWEz/8Z4pbPTGhoTBC2c287lGImgPCC+/
HUchl9g2jEZ3ereqBVDZInRfGhRCGiP7cKqBV3caYuqZFeLGTwpEhnj7tDMbPB15
6EF5sU3D96ETtznoo83CMbPFJurNgOZy+6nFwCHpVJpIxUy2kcAY26BW2d1LgBjL
l+5dW0blpwvLd7eIgaqbQl07UpNzhhJ/AMBr1J3oeDKmadoT9vrliZ7ju9Xo8+ow
r0FMfRfp8ePYYVW6tjuaJaPi6YANNU/AECsWxy4NcCrFDnEoI3G5Sd93sHl9SVZu
6+ol8xnglSRKw97EG4OuvLeyH1dEd3zv++1CGd4k2yaKrXkecOsV8PWUlK52ThhE
yUE0TPRfhtBZzZdUEV9nxG1bPW0sMED6Qj7QRSc6mEkUTBLdV88jd8sQLyEzqE7K
1eswwIkCJC3drFCunfxFNpowTU6t9qc3GjeKeHgokxGNpBeYU/igNTADtHZPiL8J
/B7kvUotbfeUdD5+/i1lIElU5LeketkJYy+PSJsuQI/HeDK3OH3t9raDowYrE/Dq
+3zcMatd//nm50OidjevH/5vFnJCSxijmS98SFWS2FsANnEG+okTUbqCOtXYvZ8g
Q7wAOkFgHnNJk5S646Bxij1Mmie+j56zrk+X2rJueJ6DJCjzi/Do8OIjBCcEeJ3C
uOr3h62i0oivhqTRKNZcVJdRGxa3JlMDDOZHv7PtPaMAwuumw27DE+I6Q8TC0qvH
gnZGDQRdNiXJH/n8xfOf/4/LPphTxEdNRX93t7eOdSlF9UYsHXrLkb9U/0gw5E31
JnsnR/QB+UkPFZHRwrsFW/dSQGbLNwIffrts+xngwbCNZzdg5tRQPl5Yfi7LmMbh
dFemj+eXoTbX59rl8ZNDlKOeaBEJIas4PBrw66fqf0plPgv3sauaPh77LW1TfBDb
70TOxiJJYEbT8BbNcDm94lIeSc1LW1MYws362QfoL1pg/dzfmxsvF1XtacFqgLdM
5TQrFEQmhYamogJ9f2aUU/nzZZtkhP9jqjCn1D4HrbRi1yAILFy/kqZ8xYZVwvqc
UpsUxJQqPSbnCVlwYxE1cDHItJc5dY9neyvQ8/JBvM9YH1/N47oJ61hO8/fYge5J
2ZVOGtJplSL2mSFlC8AxSHEQWRX+DIhiPSb/uBJSJSGEqfUIux5x78odyDvcZXo+
INr/LNkb/3Q20tvwEUY12ObFX8bPAjgtyzWnQpJUWVa9gE96W2wRGHnJOmWOQxP6
4AJSIe/I0FuT/B/XtaVlnxHlo5gqLEH7XIv9WyssRmoAu4vN+w4b4e5uiToHVGU9
B2Wb2cddZAkpKxkoEB2T2iYgKG5LGnbNkuIckq7aD7i9Hk/JZtepVV9AgRfcapq7
jBhchP/gttAKSTlwxzPScik/IEhQoEGqdlGPUJz+0gLtxonYiSuhBS3HJwXSo4qu
koUwVZL8j54wXd294dPEvfwvEPECFeOXrVt8KhRhbzya8yoNZNVeLuhUH6CbtSNM
mVtSdgqDGh6xeS7ALBbZGwJrMeeXQsWj+NNwdIu57ijvwsJj3/oMEes66nvC18xv
JPFmgO+FDnUeJ3OBSvVyJrGRkfoWYZRJV9ILFoeGEXrAZg9YMUVtHpUTodzduGS5
0paOw564BX7nj/foCywMP+kGqfCqnFd2NrkBmarRBQf2vAGQkK0xWQLPWwpQjzRn
mKF90SCV6yY3AbHOHuIShyueG1xBP7W+zzCuAinaDtUv+XG3h+Y9jabI7G/fuo+p
BzzK9LTe89b2FnzAkA5vJ3Tlqmh43ydFd3xxbQ47Y7aaIJuCxzHlyOgylufZBk73
ZYQIFc2nADyD4yjtf/7C/x/ldeyfDNhb5Zhwo7+sTOiU/8Iot8sjegmx/hwqQFUe
z82JFmTkZu4wOpU/EmZc4fai0QVngS7wPPupvVUz3MjTVxuuMf7hklfP4Tkw49bF
JHpVllbqsOQRpHlX//BlfMmA6zMgvJaP9kl3+ycRA6i9aV2gr5jOtL7hflB3391L
vrwl3CwAMrFLag54F2LbmmAzlS03/Lm8cqo7Uld4KvcuaF99GtChjEB15rSy7r7w
halk4Oav2D2Q9JOb/o3gjLyJD4hgfa3zeA+Q+RuNxy6QVkIKvctn3/2bzMj9Z17L
Oixi5SdWuVltDHbYQ6h0Kzh6Ob/AGv+KqEFUEcgLCv450WH+LkAlpp49G8LTS3by
efFv/7Sdill4BN+zVgeYhW/fbUHuaWlS7SrvJ7wr4eVmwy1SvKLuk7WOel1cNa4X
EUqy6DJOqw243X67AT4U/94FSjJ4WaTGUyYJ85zYPfZGCrhqzL0iMQtyiZV1MDBi
b5gnvWZKPVPowmtV18As7YbV4NhLFNyT5A75XqaZ6Wyfi7InwsUe8+0bxM/iAV/V
imH9a7R8xXOJWBppHmISWmNTf74HPCFGzVxa5phyPhsCFeseI+S9WMqM3qr9dQ62
tEMm4AhzQAaIkJ8HpsNE+I6uA0MA7zJXZdvNCBFomQTxJUEML74aR5gogEPP7rbG
FQpKNb2dt1CKvSBYnjMJVr8JHaWoVF8XRKOeEVuueyGhsKNpnneuaoEBBuq6G4NF
f3SFFuksr/DC1g0pMiar3wyxN9l3OpebE5xLE5w8VjjYhJFj5tk9LlLE0oZnVIH5
zyoU97TUz0NDEu0WOi1fGdVju9h/EiS/6DMdcQH4wOud71nJqdiNChlWxE4evz1k
D3xdO+11el3k8v3n4GplcGuctzenYYOZtOs/KNmQT3Yzbfh3Av7UiCJdZpVaPC59
iw4/kxAXVwsYvQxJZX+OeqzZlWHEY/A9PztadKRkci3cL1op0/s6kh/Wpbhwkvqh
BrYCFSzOkEc/JiLu9P904iGdm4aJAtub90Q5aFuyWpeoYkrXHKYMpgWtKTfFl89T
pe8nymO3qVLF+CLOmKPmiqkXd2PV7hsogMibZe9flXzCIlq+uUltSf2UYLk1T8KO
z5nqqT/njFLGY4etOHYKd6Ia/r77VbO4b264wYo/WGhle5J80+1GobCPLC3wq8nD
vUeFUq8budtIzaXCxnIOa14mbbtgUOCW+S7ssCsmsrE22kh6QAtWXlYhCqisvbgw
X1cerZhH3RPGYwA/W2pydnvOZ628+j3lt5xM8140aUoyS0QALyA4PFxKp0zD/VOL
U6KcCYOvKyx8Aoti5vOKfIEICXfnP8FdVjL8qtYzeRi5CgeQVAWwuTNLxpvRSbem
/IOUakdCsT4x2cHvdgGi93Xvgsp9iMmFot29GoPVEnqFZuFavTLj6Kgh9OtIeBuQ
LFNZt4wYvtTNOBA9KslpNcJ2nohKbsly8GmJx6hL/Jdyu9a/BopUpGSei55ow3Cn
FyaTy0wHUgDM+rDKwoxpnUG/00EI3Y0DM4vmAlahKkmJhzzqCDcSjfP9/sVsXq2z
eHw5u78pyABXgz1ZpWwGtA6Wui5/EX2gkoV5KxO+DU95mfdaxNMXOqCXO29RhWpU
STK1FRGWf9F6EAkIPxNBeeuNjo7QPiSqm7MptkuW+Bo5iny8VAlGgxCtDzjMVHvg
SyFTLY2sdfRSJssmk731myoo8540WvmVZkDLtN/oEFXcnxOIpIxmEKcel1XO/a3a
+X/9DzthnLShI35xPu40Qd4b+xXVM21J3CyIOXtds5WerVr7EuGEKwv0wR6ZfprD
TdFx0pJ9/MFruMkxkbMoFh4Eqcb29K7orF5AWXMgSo6imPy19duzxoOhRxQD1ifU
dzDQoGPD1rXhNYlP/hFgskiAwpGaGOheKaVr2ZpumuF9rM578AghoctA9p/CROi5
QnhYG5aK+IuTY+Ss8cxxhf9Zaqnfs1h4bQgQNccQo+oBHqh14mGOqycGyxLKTEyp
SfnBUQ7XiG2fbs89J3K0VrjKK9FKNnilIPVF9ggg+MaEfEPiwo9N7X8xYvwpYWBv
y3yNxZIPUPwdJlPyAL7A8WsphkBQc7aEYMiO4FEWziLAYEJH3nMb1MwY+dekC2mY
We9bO5CDQECF+bj4heVWTAZhtEurZQjHUjZcov5R8GEfYQXYV2nA9NbHp7V7dOrr
plWiuNmlZIx5Xq/pmm13eg4NjKty7oziRlVA4zgOJtvSMc12Q/aITi7mhJNfskCd
pYVXIC4hPN2ILlD9t5VJn/HPutvOojrXaM8mmx3TOAXX2C/QYtlwQ1KdkeIk2mvt
y3NuCKX4SFpBOE1lXZRvN6azqYxSPaoyS28/KyjEF9qtUkMOFt6cyph8Zlses5rD
afq8ZEGrc0FpFwd7PBCLyhGBkQd7LPghtY8crP7hYxATJrhDK6qCKGMiAIxjBOzg
3ZhNWlYSU5FwxEwGb2k6Pa0aHWUN87FudfxqjbbOs3XDV/HN7KTetH6Li/fQoGGf
8dRxrGth5t0a3iI8ja5ggs3nvBg0+Xq4bbPUcI4LeRmORfuUcaUUzcKHfXI44fzC
S4w0GZGc71OVtdcXxO7s03n0MaOiAlyDSx8onbLeEY0y3u89sFau84efO8OWvOLh
LfQGG4yTxvMLPYEphgxAtV6JpchAzywok+d1XUg5Aj5h0G2mg1Mztr8OnDYO7jes
NKab2GbkI5vLAPbUhn5ctno8EhXioelnii1d39L5KIEqBrREQ8qMtYkaNSoqo58T
rfk+gK4ygKLw8eaJvtgDuJnyDn3hygsufAj12bs3Vksl3wnBY+6zPLksC9N410uM
qhzlhyo7e5gD84SjvUvSko9mCdmf0wOq7t9yr1R5ojECa9H2sYFyO4xcqNOgnrgU
1sHaHsgLAM1eXg+ufJQR6WNpB9NqjxMrLtFclr9V8eE6odjOl5jbvDZUoNTLu/Oa
XVxgoT5i1XHmUQJ4kduK22jPwIDPAPokjz2b8Q0/E9IusZI+XrqmhLp8nQ2I2oMG
H1Wt7ENVp3it3mgvAx+lXwrV9Dw7+Kqn2gFXJqBrJLakvbPyEVGmrscCMaRNdey7
riGdmd1UmsF/FAl0RBhqAE+4fe/m7c66GP+0WjMbrSjXJ9HVUEwECQwGbn92Ay+i
a1MNlhF+/3qQavBc8rKWeub4F57LSkwv+Hhll3Fv4+WYmisNsGCK4cX2ZZmBIRaE
ONVEFAYfbYqO6Rmim2BWVxTRfdw/4+EeSfrEqaWN1s6eRyaHsSeuMnV5L9QhWw4n
t4A9CREjWgCpMmyNVSvsNi2P73/VP94vGKqCOPJ+eO9Cz2v0yfzKwbPL/PrqWxfF
ihf6OKCTAibed2/CYMiHqUYPvWnxXez0nngX2gtCcuR/PnjRIcP5nn7ZyZXrtKP0
M6bY43QBEQ/HFqwKxO4oYCoCsPJiIJvMwYEoAvXxAKZXfpg/Tl4ijQ7bTM19AoSs
5nYTMNFlDhFpaiSgFDwDwNNGLbfoeU3o9v/1RP7KY3eh6Mtn3QIO2lztR31ZmyZQ
sszTxntpcOeJGxLy3BwGBLo9KdD7NA3LjK9rRzvYX3Lhe/ZhrRIcyckeaL5IrDoH
44hqohB0l9+356yUib1PwnYp1EZf+TiPCBlN/vfkby5TiF+vXiQOFRPsqk0FCc7d
HqoJ0rIPxUOqxoN+YTVb4KON+kR4uqrJrY4LqR8Rpn7mp+x11tBLHDqMC8ARX1wg
K1e4E+pvNZTALQnC3W9Tu4G9HWsJ0mOybj5ydzvbxgV6w2F2BqPSR95LynyFyA6S
2sbNLC31adA/0qL3VAX4ZQM4VRn4ClOUTGxleFFZOHDrXOr6htv55kw/WqCYHOvQ
WSYNOC7Sj0ZdT/Psirjj+vlKN2gL+naqYj7WpcwW2C3xnRWdESBQs69Rjh8LlZSB
4Dy0cQRKeyN73WnSvDosxaFGgJEx0cUaTtMhdlXMgzFjOzErDdB0SVeaGu2VVEqa
HsT79nmEHUbgbEXDU/+la4mHx5vSjJWgqDBa/v8MDAM6/WBhzTD/V0H80BFGU3pJ
c6QD1n8IhQgFR7dH7ySAex/h+0FzdfVN4cAe9MQvvQyTIOyeA2ROJPVSvv3CvGTR
7lWd+s4qt5MDcqcR72NMIyFzhSMNsgJDnMzpiWD8yefJDk/mdIwHHEBwd23kOWYl
xC8xqqL9yGHjXaqejCDxZ4z3m9j5TCFzYFMaZetq1Y0xxUnykNqHxOSpAFfzBHhs
DkCSiH4RQ1aSbtkFASr+i7Nq8jL8+IxhYaYgHVIgURTcEF12LIZxN95NuTNS0vwc
VhBxXi9yebYa70Uc2Laxvh353s15LiWsdg7hccDDz4JPCZNFRBjEFznZp0nYYRSX
uTJnVkeU9UT0gLgv9yi0/e7WpcDYhpjwDPvlOFXjCZk=
`protect END_PROTECTED
