`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG+VS03i4tA1HKGVn+M/HxxJnk1jzqDeb5i83SRsSoYE
766PSFxDbKI90psPtSuwFMWvaq+Sjp6XKzc4oIqAcu8L3hFBjUIgGZfbjgNI+6pI
NYI4TKhRzklxWp+Uj5mdhH4DbbEFAKuyycQuwjowGP69+c3DuI8fArSYekcyAXo+
EPCDATD2PogPVTCCQqgqqQ1Th80I0G6+UR0caJ4jV7NdAiX3msc0LrEaaGKz6F2W
`protect END_PROTECTED
