`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePbYhKxgJqHJfjgP7MXbsJYChwseBUetFgnTnq9mUEls
rwKyuUD6FhRgMrdj0ax5i/ofBOuQwKVknc5cCzsyVWSx0n0agtSJMLlreBMsIr7b
rVekfQymchxXxPJn9sLYxVX8JICTOYrxSVP4teaWdsfjYsAPLqF8YUSEfReVlImm
QExQvykyyxXCLs22S712TaDmKBcp3zoShoE/5jFrgIJAEoMbIBnAsLiTMLxOio3D
F0QQM3FXIN6MRIkgeri9jy5KFJvn9DyYSeXRvK3UO6FGXz9R1Y/t8+SKd9f9OR+N
nbsqIVbwrIH89Al7Do9kE5y+lE97YQWSIfoWKPGkPXssU4FQfO0oX/QS1mcvFqLS
bGRwl7P+RpvWvaaj5qs522EWNXtOoJUSNKZbsCFS8J/62KOeR4DRS/+S8VPb0PaX
Ea09WNeSD1D5fV8ZL7Or+u1P7zNMXPy242bwUlEz0NHtmTzO3LW3jL2GdSNc3aEb
8zdGzY2szVDbkg4C5mDBXu9NZLKbkB5T4kDdZhfMEtIp14L7y8jxNbOrHRzIlFPS
T7Llge84cKKp7wSJo+95EA==
`protect END_PROTECTED
