`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHXbB3kTQ9M1UaRKs9hehQEHN3H8wt/H+r9O4HkPSrNL
NS8J3TH+eFbV3JCzXY/zVTSOpK+6v8bRR/8+0Tgx9WmyNtdhvUsOTQixSyFYLXzp
+T7QYEYwekOD0QIHoG/FrupPxkL029jxmfRb83Rgi1AOkxtyqlJ1buWWHL9DdStZ
K9UAaclAhvIQO8xqv3lOvl/PGF1pbo8LFPNHKUEprm+iXzG+pLzSwEqDjz2wb8ti
6xDGjFuqm1l3meEjI/LCAAtyqj1xIbFFr60AyxBWzH+KMJS4D4e69zdcb8Vpspt9
druEXTSkRI0pwDpqtITcH2QtfyDVLD65T7GdJ9Fgp2h7IyAJiiFxnQ058V8tZhgh
vU8yzoX4yjNq3JHG9Prpnk7Jqnatae7RuoLLYLfva86f9LNGDT7ozWtGIX9DsmZe
T+RKJH6yzxY/PIMRb94bpeLInPfTlsT/QUMYno9vOZ/VHGR+DI4zuw+BYlmEQRZT
`protect END_PROTECTED
