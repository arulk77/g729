`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveApO/6ltL29YC/BiVzzhwWQrH5wYO4ilO3nATexSAmaf
vwnZVOnqJANgKb8m+ymdzBsrHyi/i/5r7oI5rOcY7Ladjr2uJj4G6+h9YQwEiQOY
yNoNoKHPlhOlEOKCrouraiLUiscVFQp8pv19u9ZcQ2v40S5u7lw1F4fiBJux1/5Z
1XZqn4dP2Gq1MrcTTv9v4njyPGmOKdF3r0s4aOgZzAd6JgQmBNKrNK5kczk7AzxH
njpdn7+za24Jc2vQfDC2yWbIh6TOvBGMA6e5yvQV4ttuGEpWzPMrvMmEUc5rCHkA
+4IaGjJ8Ev8TjcNNh2wvGw==
`protect END_PROTECTED
