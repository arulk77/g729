`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAZCCkmIpB2VIpcdBy77zJywjgdQJEJ0hVD9C6WlI37eV
E1NNxTjxhZ3b+OCHYFqRYSJ7jM8Vjz2nXO2MLPao6K49qJi6QNRanXwDZwdFne0a
vPKGoiV3wBMHNb/FhM1L4WqHfo/oiuwVixypzRxvvTSgm0uTAdS3U5d2oLhBh+di
9B9o7CamOPrVIe4pKlllKw4DZsNvW3kmiyYnVLCA1OxPH73LvnyM+5F4aTOIc8zo
n2tMR/8HUpedx0XBdJcj4NKYfhlG2tFIbj7rejxfNeRhZUb3GyusXBnaHHiONRRL
5Rryoc1/jmOpBKQEyTFicTk/J96fTTxbT+d/G4aS2PnaiiAJxRbu8KBjTFWahPGn
khG/EZz5uxiW7GoziyCjcS8sIoA/7Q0rBMZsVB6ultbIoLxv9GaEhZj2QRABulhj
tdl6skYtdtlo0/XtmfdxpSJGH0141GYK1cUlSs6yaHT3jXNUEP/psAlpcUndJlsd
9HmkYkHXVHqfCb9bwDv0u75xZzG9jd1RUfeftt9wirS2y2A1UkCaBbgImXDQTEbY
UUEY5mhn36q6FOaovmiT4nszlyPdhw4W6DydpZsLTHW+1laq2kO+86F9uT6H8oaz
pZqb/J56Ryaok5I4R6c5hzKQQc8X2FSz7E78e0p9BKBe1v6Y9sLa73YrB0jrKoQ/
fIv0zLYSEzfocw/tnWpB+OHoykcZV79gDOL6GxUaynB9gflp9dd5pEg90gAO9gX2
Aulp2IHHFqmsWgW5SQwzSJhPiRyA6chuDOHgfxWKPdGA0TPlU2WUQMRPVj/GAxjv
6hPCEpNP4ZfXT3J+EgZJyIVkLRbLehKbhzVoPSBFlp2svEMBuo6WzRqmEFTA/gHp
r4UCeLRWP7GWipPeopYClWR+vmYwq5N0eY+jTO6c77BokhC7Q0vH5Cq8YDLglzGR
uFvu8nfp98ZkeUNdZ3Byuw==
`protect END_PROTECTED
