`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAUtbRIunVmBmFBnxDEZKqHRogWnopIIiroAObsYbiLk1
+Hh1QxAWU65EWJN4sAjOv45yuwXEigmWiLdT0IrhHXlPxvZk9C9gw8Q8Q0NSRYvH
rq2c2Uo3jHiJx/sh/tXUM9t6m84gHX023lKlTBAmEPx4eALwCs3kNfElk5p1sxfj
gF2X/B1tHxoScnokGGg5WdliZtecs71pxM1fCPF3aodrvTlWFhxoW+KAm7dOYhyo
h8fTnGxB8ryCPS90cUeKJ9TeC7BOrmpSVp0vblpyysbV+LkyJGnnfCpJGlHeQQyv
VcTo1pBr5xXUyDPqSM0AvfbF6Mcf5dGo13mKatH2V/v1tLG7Nya4Gcl0kwYNYebN
RSS4dfkGF585JTK/KBduCrEAiDkxSjpT9oK0h648D+leHbE02976OCAgLqWqZvbd
jFKlR7jGeR/IFFlUFWLXiJHjD4O9aw2Zhye5jaIBytMP96Ey4XuzVCvftd6ccdeL
z+MqyfZZTe/i4p85+0HGOk1esqYtxMUtwoqZQ3cq3+C+b3iDKSjSiEQmRYAEz1FQ
uZ5D5nrtHsc8Se23AuP5P2wk4JCowDrXWKjl0nMrVeCsgyvpHNuzoR/dHkYZ/CC6
BfCjnHveByBViah+G1gORXZutxDRGdVKGj++Vx6m5inXHIYDwgeZqg5ml0Vyk2/w
+YYoV87bJv4mv5YA4I+JN9sd88ZpTKPDNLsg3IFeK6hxGLlxpkLD9U9SocvF0shZ
rKpoqC2Nl0y9YEpMHMcCFZREo36aXhsC1kSobnetDRNtlQdrhw706L3NBhtI8A7Z
hhjQDnZMudvrw26lv3UrmLu4jGD+Ugk8+lqPzdUeK1atGjOry2/EJqLUH/fJJME4
BGOHMQm3J3JH2+CG/Wcq7NQLHwyxuoiDac+oNsAIJwJORMxzYQvwvW3frx0QA6Fo
lCd/7tum6PCoCkl320p0cGv0jGggJTtDNhPRR8fJrmPkFy71FxbN03f8A9G5Sirw
ubNaPpyWbAulwiFOaV+bg+rE/wBrVLP57U2kQ0nP+SoUT8bXCTlTUjH23xv8DGIs
wLGc1s2qpITuJ4jpFas9Z7rOEUom5Op+Nq7XCEUdpj1ZMZqt76L4OaZh56lnb1pc
W8oFV293bIwlCm2JQ3gHzCZ3nM3LO488AbwuimCzP79tg3iXZOWxzVlO9DylBuIS
f9IWxbnOETttBj9jN6PtKBHVOr+rur0adj/RIvnDeyrk8aJKV+UWLDNt+gozFlgT
jSuRxCtfYttMvDqOP1SUNV3dH8Xe+mI10pNHg0eKrCycNhtI9124vO5be7tXhYzV
wtKw+A/mPHRTVfxQ/N5LmTcM2Dj7THxzk3puMCp9AFYnKvyCguBhtiOhgns6iOu3
mlBvVTKzqAyTdy1CJnNcTFJCAVrxoC0DAYIwKNkPR3ndCEmQksUqCbnohd7ylQ7m
BCnJA7kJ2VzJ2pm13TzgakVPGLty8DcdpNAkml/ZwWfgB5n1XxdaLG/JyCkLwHBy
991lZPA1LxpE2iSjjtfgBrIpgSzXfWCh6DnHRt/nqcDzg7lV4YygxIY+fMOu9C6x
YsnugUqMPsW9IQE2Fp2DMtbC4m3RZ3g2ZAjBG0FRnvt8/42xC0a2qReY4piZImAP
NBPVHTWHiqs0koKba/LHFs4BFlSBoxSAWzOgLMcu9oP0gtRUtvj3HMcpPuBDZvkS
Yf/moCSD5twApLU7OxEPnHsO6inFTXMdWtpArwqB4Fu0Px7amKVIPOF/keldN55r
7sbtcROUw45WxMckzsiQNAOlh5JBT3F01bvZzVfhWZroc2b8EpvnilnSBNNgIAv0
cYiIRhOk8JLD0icHSqM8LaVyrahkzekVO5F9u0GgNzZ+yK9yG/gaAZ0qOc6KO7VM
TmJODTAEAv7ceoFeWrqA5br37RMYqMOJB9/kwGBV4j722KJVekzFgzSqqdXrggT8
p9yaalloGekowAWJGmsJv9WQpIK+5k0rp9dOOHprw0LR0QcbWEEz1QR87p2xN4ur
LSmNcv4tx3NzrgHJMm5MMhyfJCypd2kgkPRBm72Ky7qENkTzjFYL0XZC/4uHHS97
jna5YlPyPNYuO8hdmuTwjmciw4XZOzyqv+12VpO1yfWTd8vj2qTT6hO1TUnpxfrG
T+OJ2TB5qckz8tfJkj/1kNoIrW9w4ub01YfSGqw+hScuxj+WquWFNXsEV0RGwSa8
ZY3dwqKDK7Nzn7Eepg2PASAvl/5o8pZOZDnLlH4wMDWiqZ2o1fRUMidfq2Nr/Y6+
S6ZXnnNBhO1FTNTvsEh3UWjrBJUZJ18yThPPaDuLQY3XJThlZbCF939jj0wRnLSV
/tJ1mT52ybmU2FCKX9ls0KxfSt90Xrv4zdnpVNm1XiB/lUiqqyyTGU9pulQ+TUwf
AfhPV19LIMj2zrgBReqyJV3FtAFkRg7B5EvD4MCjuVJGPdlV6cOYOZJfu0XtLsJk
4EiCngiwP6ZnzMdVlriJekrsFIj4bJf8mZRfPvCk2/hVp0G+Z+x/8rWrEbNH0OS8
9zB1N6jnpox4dNsONxuCmnTjJHawvA18fqAVj9i5x5jsvjoUW3imzVtE/Ibpczfn
ekygeszT9CgCipNO8sfwZVqhsEl8IL47WmFr2tuEzu/++xfnJdUXHDCqv3qVJnbn
8XyA7F0L1A4AwJ1ck6TppeIacRv+Ss5JGT/cDm3Fp9LWY6ZA1Av3KvpzixyDO7IS
p5bgDffg+XIQwcgA19MHOOmFhnQKBmCVCk/UlcG5pVGoVFntOMqRiPE8Ed1cVIoR
eaJYQf/lSFsshjXbOkhaDKCdP7i7l17NM2furDd8Wfl/331tbSmV7utT6zBCl1e5
k5TjzBQAVop1eNTnnSzatdUJwSdj/lTUqcbjgko5YLtIG8mfCtkF0kdPo6IzJ0oR
U8v//kMysAvCE4yzwhnnM5y68APkKzE11SF2ZdTwF5pnlNPtms1CERHl0aElm2vu
/VXGb9o5zGfwt1cPmbJjzT5ZRWdJ56LkNz1il1S6LiXzBt2iuczCwwS40ElkqZHc
WXeikKF5Sy4Ajwm4/UCTSytoWKxejrQVqoy7mIZwgym8SSbChQlvJdDmStcVh7W6
YkWx0CDbI+rEca8aeHoxbd6tmR2sQwOfCgZJubqBjYJZe9kR7P+r03iWtCLmyomC
biPz7Z2mTPWPphm76Kchmn8Oap43iDL4FlrsH5EGYrmHNkD1TWd99S9ArqqpnhTo
47RFsYiks70HwRFKFJ03UD+sqCeDXMVwWpccJXgRrhWxPHyNaj5dXADT+VlURsTu
q0zzzl3p3H8G9fYv599u5UKBsAJgq4jmxJ04WTxcIMtgBnLRWpDrYKs/3FUjz8q4
/+0miuyKbOOBeTjO/nOB/nvafZToSYKm6zCZKjj8d+KgqXXeJzBKpP6hG+PlioBh
z7dBwv4ntKthbGZ/a84DjcNdPa4FjIHOF7lZ2Pp/lKAA5DRaCsGkPZXyEZgS0nVz
u/VgZ6aVIRmE8BOxiVxRLBNy3Ba3SThX2eLnRixrdR4RJvQd2PO3yoBlQzYL7LXf
NzLW3VQFv2C5IsWlr2GORKdfsccMjeoyOlOtT4x06UAjAFLcWqK7SwdD7nPso01F
VpTHH4lcehIDYVR6FZg8woB9lZLHGmSPGLxGydnHbUMRDotfeU6UmdCiZdQ3lbSh
fkZ/inj9WuXdg6bKh8TfpGIc/UB36IhUIvKid7xAJVEs8GFV821kQNfpLKeJCrA0
wh5CWONyokA113p1tMcQ/Tx3KuyWMhb7GwVYEpouQ35YOl7nBq1GFGzwzYvF592v
iTK5WTdRQeQA4Nn91UJzVcO0H9Eq2tk8u04kIhrn42RlXmUi1L/5HgvXNXz9U5X3
V/pG7yOodOmMazVWDIJgZI7Gl/UGabwfQHA+fpiTmZaEiWE1IdWvuzpNhMRf0XUn
eg8cLadjqixWTRfBUYTun0dctSazd2jSnfpMmaKjGWno16+cqc8xR+nPq8SghIq7
Ekn28iL5mmc6L/RZFMhaDJE1b8ho3dyb8bmkxmWP/KwMowd4WEhZu2ZaoDggy2mf
lHlHJHACmFIuqn98C5pLLkftsmmj6gcNMZJaCy6iU9vCMB4hgyhXnUsjMVqezHaJ
omSo+zmJUZCckYH8HSNUmZNOb69CRgWMFNVxMcP3g2NjxrNY8wWHlBDWk13f5R2k
0x7usV/2XhjhUIPTkQB4AGZZETsnabF0bQFRrd6vP0nMpGzOViI46rNMq3/PFTi5
yaC6ZNqpifvMnpOImzSsvDioKn5XatH6eLJGhQEU6ZYJwtKk3uIWeRbZFH9TOOfX
xxpcFXNlY1/Jbi11+BfRoKor8UbRJuFtAySEFaDWU/KqlVYPaDeWknfQD68h3REI
inWObptSTxRQoEtPslq4B7KTY1WQ9no6XzLZcLondogs7fBolUXeXj1gNk0/mWWl
UI6VE+dmCl5Yv8NyZeRoAVuTYRaJ7fgsePWTkOY/wlwhyPaSNvYbSYZnC6VGEcly
cGNfdQiqfHw9y1gbBiJcvflAEFjmkdi39GHEkaNS0ww1RsPqvH2Pq69QSlCSYH7K
gYPelmfMPJ/ARNxXhiMVF4+H9WQ1rO/2k8+O957E2PwSuNfDoj0tbQBmd2Prey31
CLd9bFJGzT29O2koJC2gAYjeS5C0k+ahr7wqQ9qyb5o4ZGkmUz6rwahCyn1kDHmW
yBk6av4lBeqvISQ3INEffi42dgJkL/th498OzIlSFdU7zpv1PJL9bvzRtrk0Wvze
2FUQdIOILIlRn7lNa6EJXLV41fZKIggpJtXwhDEmKzKAn3pxrCkHDlTiWqWx2HaC
XDCQSA1Tyo9JZE/0lkAKo+h/gDsxMhhLtKdjl55nGg3N/yMpqHrNSm17etTW3lVW
qGeDtlH7547rcHuIC1tZrD2cF3lUVxM5JE0jX0Yg1qt2OLkHHZ6MN99y3CMJ8LmE
2D9U3l8mqddPg+tprSkbUOPeu64aGirhqJ/Z4kaAlUaULimMHObUKeGuTOhXIO6p
q2WS/YzQsi5UzzP8Job/97KdSqcl3UK02vYSgWHxz01kwXSneP9vtQxr8210khTL
7LrXe52XZ2992s6bIs5rblwsf2iEiMgNGhWExXj5XW+408e3NXQWrHXo8PtcTt8j
m9R9PbIAfPukf3iCsnxGOgCuzHtZlp3V8W0/iSrzEH5M0moTvqCfM+qT69VZaelj
yMC9tVHDug0YZ+/W9QWP9as76BarPgbTePztkwG6HnyeX+7JsVvNozlGOk9Mr9hV
fgFTh7tbjZeKzPCPSbQa23J1g7pAQM8S4lZqC/Tl1Zut47faTyIVc5o+vSavZqon
5syW1YMqX1Cc+eFSDz66FiUV81fjiVYDsLXYsoJYerjnFVu2Zr7Y9Uai9ljOgO8d
GKq3PZrY7imo2OR0vOAIFyUAH7RcSP8DTGufiRfWCdrM/9umAl8/866sgT0DeCCx
cj4sBRtyirm+7r5LNOmmQeiqD0ONMyk8L03oNu7qZ8Q5Exd5CzILuKQDUlMs8+rr
RfoF90Fadjfu5EGOBBD3jMwuQc4hNKGYiiKcb8DlpSu1aq2s1Sb2CVx2EKrfgt1d
N/wpA90mzXwAHYWoLHuRDQ4tP4CDxAPghnM9id0ckXGjZGPEJev0344RFrSBzS9C
Pid3Wr1s6UcoBumGDkRNu9FNU6k7YDHLCLyaxjMpwbQ2FgoXvmYA1n4lC4H6XHQP
yDn52+59t1XFZmmuebgk0yfutVWx80cx/9ejO5Wq3ZHvwfrheAdlxwPXxOLjBJqe
or2Dcx43kjsmUTjgREXDbu3JuVbgRd6ylXNbAhZE+spCRPv4b1fDYOWYh/pW3O3J
UK+sTvHF0vU40VqHXwP7fEgUeyAefWyfd+LXOkl8CX3OfecJSUt3t+BhMC+sxtus
wb+OJfK5aCUWyV6LMWixOrn3HOnaYe4bsvLXRx/xJnkjZjt8MNk6MhlRT6y7iSUV
s7DNC/uLHg6JafS7Ll5cinIPuQiAOgTLamz02E9Z/jSUzwCcLvrvtsvB2BT3QUiP
n3yxYi8aDe4lkfJ+J4yvG1fdyln6qof0d8y0TEIKlqVcO7CpX3awxjmbaj49FWeU
0qrwsxuThNPdUCKHrnKV2TKKrOn1HGZ5jyp1FgMXjOQQjxWE/ubPXVsCkY8bS810
wvMA6/aLpWPRkdYscsID75e/so/H9uBYswXktf3Z0CrKd5PrI6X4DqsuRSiV7XVx
44lCIE1lskGPkEpvSgTf77QwWUkZTL84GQjFgecpXct03LOBvhVW8uE2/pMNxo1w
CqgF9uBvsgQLENWtD/4In6FBtYasvrizsLzU2jQxszaVYeW0tji/FbedrhNMeAeT
jrOuEY4DrNUZYdqgw4Sq9t4qvTtmCxJhU6HxsRRrMyRMKOw7kwM0ilf+xwrnq1lb
nSHGIb4aRwy7D5pCOZsnkSjgK1i0MSGHBMLOySbuqFvXmym1d73QnbLm6hZGL3ay
fYKNA/QGeQ4ct7bDJVrHRduduvaO1NOOxpLeKd5aqPY2nUQKGwSAYmfuQKnZIKuu
wm0YX2Degn2rz4k/f4khoL2dSiL6R9cdFAje2/YHbBVFCdHXawGNL1Meun3qEiDB
UMBZ6TBSisHEBhBy+6L+rPcxZIjNpIkGN66SSbUCNaFKuehW3JkIahC7CwOaCC6i
rfpxYt44f6yBYukc0/CkZ1rCsnE0JmW8Jztx2Xlo45qarWYqMJUDO7En+flJlGQ0
e6ihDCvoNud5G8GfPHKwyAV+0EKLQSnZ0JwHgeqalQLDDhtIBva9AMPVzAgpoCi6
HVt9lalUY9isy7/CGYYyeyxjlBdPWUtXVTw+L9FEoHPek+jinbL84CpEmIh7yFLI
5BySH6hFdhgbBljfs6AIr7CDuirB/WQEYt4K9MA6dsktKQlQjYxqS6EsnWbYE40p
FMhm5BIJz/eKLCfkjAQQGyOQ476/NVE0NdIgIvWAggcRUg1UmuVzWsrNIDFlHjU7
rl1U2snpULpecwNzfSZoDqvsafX/TELjJ9os5mtiVtexfAoPHDcDgYesZ4IkOb2z
qOKKFzJwlUUDS82Iyfhb8q0i0cCL9dA/6mAX5bSYiYyVYVJBPq5qMoAy0sSE6Ao6
U8/kkg51OeDXqQE9DdDlZVQ9rHjy1hmbOffLCzjJ4RiPc753bIp2WdBmdy2cIgxs
k8c8Xc7nQNiRAvEEZv/Y41qx2/Zswd539rF/S5PaT/3YywfBLEsg2HqJWngk0r5u
XM4mY03n/GWxPSOKjXWmLVGW7LgpF66rjf7sDCyQOTqNF8sNn05lBqEeaUFW8xob
YXGguRkMFyyMtEDof0f99V4K7FlAbXjOoGfZcaXJfUgWRXM8CV2NFcctqPYq2TXe
N7hm5POBdHom4H7KcZC20964gIx5dYEWk8WW8kdUlQ2na1Q2t2vQeZD5F0VC+mMa
Mcd6flg0D0ir2JkKkGcsV7wNvPBHc4mCj/JWivM9ruvsUvIpF2MjY3ev6uLMXE+k
9S9wgNA1Bq+cRcBiJULrW0BUMEM6baxXMyeMhvfVd24/0HrmF3T9O4Nra4lsppGa
jgkXB69LQkofkZ2IK85s+AaLROrhu1CGBn1lXr4Z9AS6tbXRisI5OJsJ0uLhpAAv
O/5CqzVjKuV2Qx3eAI8twdE+5+7rFdwp9awLUvMQfwqTSVIXbwN3KLeCfjTNmUcA
NjXX8IcNL6rKFD+ulEU5E+6ydCehrfDUaclUOSb0dMrU+PvlM1p62CBwxOVLnzOU
fV4VvSZS6lnOoTKdDm7Ygf4nmwRR6LExNfbrhN5TcayGZJtr/N8Drr3yVZrOJQBL
ZDuxP1aiwbTG/1d/PgByEbXllWseN34nYX0nyZ/Kc+NweBf6a8EHf206eBKGS041
fL/LrmAxwRCOlrt9nm32kuMgN3q0q4Ejqh7kF35Kaq3UOpqUX5diTujYOVTD4CNS
xuLKLajVQX551n8PZC2G1VmoayXGgCkUk/4+pvdhVxZLlvcLHpayToxvJsrqaQqF
5RgoUAEdrUqwPYuMyN6rVPSYOy9B3vlwjQGyMIEFOvb2/fGUfcfqtZFvyGc5cMn6
stgliYhvtm7XRojwQeUxrBDGxv+9R+ji78HGAl81h4uPTgLR5kuD2cznFSfb7oIz
cyfFGECnNwHUHvxPny7hFbWXsfY/XJg6yLP6oqdivI6K8ovbVt+btLvWcy+B41Lc
iwLI5aSl3EfXZ6cfWTyXLV3sTYv6DmX+r5/fnSTRISBXWr934rJuTSO3g9Z5axuY
DGV4OSJb2hYcY15dGVsgoGBh46Yukd1IzvU0JdDcYHWGSkTmPfwbEX8WqmDFVJ3n
5BPJ3hrYEG+9eJcUwpb8o3MYZB0aPaCRlluAEWhUVP3wZfHdk5p+0W6BQ+VZklxQ
0p6LhNj2NqLBKcrpyjVDxpO8yhx9VXbinBemHKxBZT948AxLye7OIvSWuM9aP7NZ
J8l6ksFUIAKuzbJsk4qY47BnHwKu9zqP+BsNczGuWoOfEswGPYCKp7B2DJmfPhG4
Cv+EkCzPKwFVrw43WH9J6s60OQuG57+sveCnS2cKH7lVTMbdGEXZ9NcF75w5H6cg
Bl7pqhdWzhUPb0atGHJwodtWkAZFSLELI+H64ErLRCcBbflzuy+NxjVbtDCnDwgN
RYwVpD5AoUEmnVSfSvhniqiZfNMuiUeGsd5ZQ0xNy80w31KTpQIuZnZpzlmwIujK
22IBuyryA5+40HtRWyYgW9IMmH3Gubk9CnRtO4POwQ+awPWO7PI2HcT+G42gPwob
M4cgANtK7RY3YfwdnX19Xzkxiv2KLgUTkzDPfmxKFDHqVtLXJDUqK5NOheHBtoEN
i9s18ZEN/TWdURrqeqojoBNsU+UVojzruspqEo3R3QUbz07RKE2KGl0/VuU79GY/
LEUCgnvYMrqm0cZlDB+UE8ygfd1kWMUrn9oogC2q7LhaRlellukBvj0LZnOQHAB3
y2bp/GHIJGqIDvkXWfLf40i41xzr2cwWgvsJQ79dy2LCHnUqd0c62qFhHM6JalNW
E/k3sADUuVYfytHLG4T9251bwFGaorvSS7o3ss0q0223cjfcMMZ1lOTfKlGjcB6t
Dk7sjqxBLfMJQRk56sHIXhkF2fh+JeIcIYucZz6GV1XVJX/fZ3Qki/Z4v8OlARl9
PHuV5/amHPZkm3FmDIRM0AOumwTEa99Yc4Br2UGY+tSfU1bnU9Nl23VxtYZxX7Ux
cwbbWwBdkG3GNRX2PGWRw5LOj+Sjl87dET9IWk3jcKKvISjCz4mpwBQ0QbcS0D4L
oCiTNsExgI+VpL2Zm64UnBb/kOcaUotvDP4GlvL3/BOIOg6vHmPAy9pc+PtpJ93+
ulY8PU2RARdeEupXs/AwRlUohHLs9WLtSF3Kbh4kmZQC7yIz0w7xx+mbZpF0K+Es
hZ4d79hCiTjHffbhu46BkSMXZ8rEHlCbw8ZCgGTKz4h9bko+y3CDP7fXR1/7HuYC
vcHWf+P4burTMO6jzHo/uVBnNxwjr8cjRKyunefQmEs8Y07RTH1U6Bm/2ot+Lsi/
1kzwKpPmbxAz4Hsfq9vC2h5Sy6LD3MQhaIVmmjYJ52eHpKht/0gjMJGKv/gEFb53
z7vQd5V5F1z8oMKddtWSwbo5nj91d1Q4RGwSegfO9B1sq9WGi5//vM1RdYSaSlaM
8mwYIeCpzP5SbzEL8Mu7iQ7v+gaBpfaFwPsW/T3C/7wVuaHgIzl0k+m2t3Mk3hj+
wvygdiKWmIsMfOgaOEYZwR30M2pxiwBDJ8hla8taGWtyy5c2u1k0FT7DG0h53jxz
8yjzH+qqrJu0NvKQdbxzdBudgV6x54AGCMbjWPgea3GEU0u1kH3D89f/cPH/biv/
carLpoRtIlMVI9r5ik/bb0/BhsVtx0DGDcnMrrjJzfRZ25ciHSb+yWGRYRGCPX+E
owCHtoY/jZBZZJSm8YmGg4Hk+whBAZui8c9pHS8y7J9YnOkEZUw+b4wz3V0LSJN+
vZheRUfK5cN22g/Ibh4ayOU6jfwa/S90mzXtmT6+qfsbCuaFaUZ7gKSlWRZAyhY4
boDrsS/RykEa13ts7nqHwPP8QqnUe9yCWrSY5ih9z2K3m1SUIaO6EbyxwS44uaZJ
f342d6MgC6s5lJ5ZyKV7ek/zaPzQH8X/5y5DxRNRKiJfXX9G/AE/dQYe4NVKFKF2
feJpABP3BabYrve6wTRPSSmd2XVeWoxUpfLgTvRXrpg22s8F3yoibhRBRsC5PhHg
pK7wE9Qh6EZ+qpYeyijU4omTrSOPL5PbgBei0hcJP7teFf6TSsP8kAUD5JPn9lwU
o0yvMM7qQuxuSh06t2hyWD1UbhsoN6uJeXZ/OLlZSHZyWDtRf9VOznSBpbB9XjuJ
TkCDHYCt0DMO//Q3/XReAO6yTmD3P8l8i/WjeVumvaH7c42iVr9NmtGbA6VuNbU0
EEvsYb3MCYU9y4ai1H1N4ZeDmkb9eDvKwsin77K7DO9vb2CiBZqn2yM6q0/iFndA
FHXaFzQXz+sNiAv5zlse0gYcRUtgVteyAntoFAKIniWCX55OEM9Uzlwbzi4hQc2m
wh15WeDAQsEnCza4Lxjattuv/MQPl0+gTkTMkh/L9refm4YZ121U5VWVZykkGe6q
qUrDz5P+ltzZrAbUAI+FWehjMa1e35wOD55ssc/JGEmalM3jpK4bPdRpT6GPGh18
zf8dvEzX8z4hX8vjI/6BMCaPz3s6wZtzi7e6dlVAHas6aCTfi6qgrSz9oMw6OkzC
XJWoSX2NorHrijLv+h7qgwEc8zAxiMPlTEH25eOEepAebfIVcY6PMvFe8f9twupy
A+VIxh6blvh2al69cvVZrZzQfsH4eOG5lSMTJTTSqACDVBZ144DFUpv9JlcRX69x
qmpMRMfz/Kngw13wwfWY/M9lpZwlLK9WQarPnJkV9uX7J/IWoYVgDMoRIMN3Elau
iTJjlZkpKcFe7JL9vLyVOgs/8dMU9OwfvM4Bh4nQ1U4y2scQRC/BvLQFSUTbLnK+
bznA/3zUpSxk0B125uzb35fzLjc9GpGgZhAz9eHDNWb9JUfABdv8xmiB0OVTW6GX
6gNTM6DzJpEUv1CoTbRPBLGnmPECuhzLq02+q6p8nAycMYIvrSWlRAdHWdd1Tujo
6T6UQH7cgWV7ft1DC/z8VWMr6Evtnrwcg3ORaJVrCn2vKyQYLT58DGPjsK08QmPo
E9OVbv7NCdSA0i1SryZUNG9bZSNnx9KxkR2VGL4k6Kn5cxuC1bkmPPQgHoiwuHiy
g9XxoZg2Eee3jsCv5hzsBPSojveu3vS1lX4jtAQmDzIXLRha+UzWFLGfXdGSc0XO
qDsc+0/EY/4kT8louFPb/eP2tn5ReHnLxr2TtaxVH2bdySfWg1rf0hGi/4dQo4hG
k5Nsds2Oscw8DRae3f38PhilCEdQjISB4CBLamCH108nuHp9iRAsH7j0oQ4Bh/qd
zUBrio8oScTnuoYsUtrXlu5WHEqkFztDRMc2/tRCyckXyz1TA/yRB/TJyXzxWDCY
aGKAYEwWc28hzfonBqe8rALBwPImGjHgJaUQxZxTq1V11A6EVgSKI1MBQ/W8nLvq
mFnaeOEIFxkisq6FaZFdBw4Mo685XvCXZiv1VhXqljSSRp5ioXu0ZJ0A88yocIgI
QPgRFu0RwEfc8DeQcnCLtONkYUVNrdG93hTvpTCazOlG2KTANqBMqPBGC110tPoL
F0655PpZYJ7taCqQYSGj6ONf3dL/D/5R5kx4oqApvrzeQzYeQiIp78gnKqF/xI4L
KOiBtZkMHwSjDQoH28Ffoak1m+EwWLuQtZasPwzv32HNNO4HYl8qAKIh5npia1JA
zX+XOHF156fLYqRKLzbl3bZX4/bjGp/+DUJrBESQd/GSMvuslehaJzHUXQ2fXp4R
fj5Um3sJoUDbfbYh7mmM/koerWj+ocNK/+K+4N04Y6Y1V2L8Qdy1A0na3SDLyGhY
rgcdJf/LGTykcSqpo9f1Dr5S9xkdiIDoCiyikymk3vDgMu3sBMPd4OiU/nL3pzBH
M4X3dkaXnwIB79JRmB998/juDdD9nP6rwTcfyLewpzlN6m9xPyHza0FkmppZGUMi
RzC8zHy0PJZcgJNO/fmGaF4B95TsoIO93xFTFxxinmh7KDDwot5SusLnaRw8a8Vc
GYv/S+dAAS+Gt3fDwjQIGGat3Hr8SowcwXFlcP1dV3FrthE/er5zmVkf/zrMpUgM
f0pnCq4ujn2ZcGuk6CJJOlsmAIULvEApp9CpmDZB1bYyhwjRWGcCG5FzT7AnT3hq
NTGDoauCs27eKJ5FiGqHZvg+q6MYjoz4jc132nIi6dDsU0VN4dqRTdsnNnmC5aom
Qx2bhv5hTHwCBoZOXCn7OmweWeqg7hc/pF7acGYYwQwxkk9Ocq+K6+9aRIeuUkKJ
3g7EDhbJyUejiWQiCbdSPgUz59j8tRW3Pw34Zrb7VPfaKOLiCf3FWw85EIBNRZyg
lQvloMvv01GYjxAUw08im8YFM6cElGMINHitlYbahP+iS50PS6jkSWspVyvQxs7o
h7f8msZSTc7/058IRvgy1SXpBhJ/TyEfGaf9qX7qWCqSPD9hSTjxiM5GBtP2NOgJ
PFOleS+mXSIB5XCW160Olq2m+qe1mMLBQVd3VUt0IYQQ/GrvQqBiRoU4qVXkZ2Yd
2GvAkmGO92juFSGHfI9nIURJyyXtCh2tdC8SEBaq7jFEprpxbn9YR45DnfTfYKMn
xgTYU++EQ8i9/f7SlHDcYGYR+yzVJIftEPDdeIwmh7fwE5tALwQ/0br3FWjMGLuI
G/jyCQEUq1lj5mL4QXrt/6FErMSkDFu56Mv97ErfAF+LEnMP/dCe/uHS9BH15FkT
xdqX3h8JcuYAMlkLZUs0hbKWRbZ3R56r/hBW448DtBaZPCT8S0e1IHNNLr4vTUMB
9KwqYn8WwNnFB8OrB4DA4Omb5aRz5Q9V6GE59+QiRxDWo2lkxFAThVM2z1+hNml+
/86PnMR5SUvl0+tlXaK0qSRwrsiKCUWGy16vyB6VUHropJ2fuusiLhFTSUVYcH7K
4Od1Khfdzhk2Xf+HirNvxj+gdIhcFRI5ROzVF/XPjUGRjp7eOb4OB/GEG9nKPmCh
k8jIvPWcPRduOumIs6HQD0eF0KWWHRiP6xrk7M+cdwiKApG4BiM2+tgrtIFCYNJb
fG86LGUwuQXKE4EbWvxw+yvPmO00lwUi8WVl8KSkCAQsdI5pdyyUTbVaMqNSQgfO
/rpUYGPlUmEXnvRwz+uw+PSdKn8kK2qaX6il9yIBfvHgj8x/s9ihyiD2OKYFZbTZ
YFw8JbYN0jogUrMlG0Jj6s4TcEek8iIq+jYKnFbMG4I/T2JeeLVWPChg+19TIVq0
oxJvla8O3c6A9dbx4D1+TUuhJjm3R3BOLAH3ocJFMHLuyWj8ymmBN0rwsEAH7C3G
gmpGc9/zQ0N1EP4VjnidX/Xjb63wYknPbm4PA30mucHkx9Zu27r+IhPbgTNTqNRx
6/gWrEF9r8KQWTQFUNSihAyT4M6ePYxV4u7IiH44yHLkoHrA1vvZDuXm7mwxyH+F
6mWcKzak1B1B0jCi7TSPYMpKtyUNEQ8gbKE3DEevsZ1B7I1fR41D8m9NjD4cw0Gl
6Zs/hCvUTIlgY/5Bpsipa4clM+Ytngla3S9TAPs87htR3G4kQlDwrBe5I9HE/f9w
+kl8y+IBE6/zUj2FDOKx9/fN7kyqtAc8ZsaVc12xdgFAc78aBABD1cKVeE11ZNWq
8WtvYnXa9fepCIYtQ5erxKsJ0PSMt/0kQQQDyJnWstd9ZKZd2dv3oskXzTGOXqP7
aiRzKHw7dE996ZW14RGnlObF7e26HNPid1m0sXAbH4j4iHxFYsqc8SiJH1EUtSrR
FhxAeBvCwR1VWzaNpcdoLxhkVBK88Q0NUIzN/6fj548gET1Xr0SkGNaMEhGEbQD7
0QL6X9c2HYGquex6fjcwi2chwtWLRVaLmhSUKJ3UMfe4+PR4ahPAAEqOobUKPzYB
uXQr9grmEQ+8XHoFeu/Y6Y/TNayipgBVWlSJVQSijzKNYQ2mi4q1lBf7GMDeNtGi
5/9AEc9Dp2E01cgpDuQ6NSZmZ88vOIFQPWKryggoyA9FC5cURTAF414cjj+G8t+L
2Lgc7ToKqsrg2JhNFoIbwW/iKetYz7gJxzdOiLoUcL0iwBTCi5Mr0m7cpx/1s/MG
WG/jLKWM4b4CtR3VN7JQHKCYFOUeJ+wincWabv8v9C6sCe2nIpx1DLEONjX5nBCz
dbNEZYxEumUTuggFk7ccEYjO6fpfiOrkgxFhnoz/HWWKDYNtPLQV1SOAxHKw+psV
mQBWP3Hyg0VUaVUCjxoICMj/eNJ4lqF5jY/W+tLTZDfsWhEcbi8QCA9rbxLMHxra
B8FyuKTR5TFS+joyiqOn/tGlYmc1K193ECylL1b8Hd0tiM1OTWq6Uq6EyfPJ1E7x
I8ExnsknbwO+m65BAZ1qfnHXSOsExysK/dfOupfDsuzwj+m5YlUruQQ8ksGN4lO+
puG9d6yL9a1lhq4GFriSClwYP/6QvM8ogyG8g2FpwysY09wvNnRo0T7Gr4xzKT1f
B4hHxR1FO/NwdWFuKogyBmbZJ7NGQwq+AwsVHhgJ4s/O/8eFqY0rkysfHOxF3bXo
QkZX5q3v52kY4a+euv9oPXrirgttEnhf6kUwhS2t52MUuT6x7yiixxhf9cmMd5wA
9HpapVnIwvgIefd2F/eMRL5V69vWEP3e1qZFYZvxSCeuP5Rq3hyVgq4/p/cNmpr5
+mixxGD4vgEVk/IQ4CdFAVjzkX0g4te5Ed+7gu6loWW/gcV62zzo+ZzdDnQvOq+9
hN3g9eTfY2RXS1rAYoVWAOtUu0C0+DPnX0IXycmTdo+1UpSB0za82ixgxVD2nDiD
9D2bgSAj2GnySSg2sGbzE/sl8ZbfPBFkJtDmDn9PM7Vtj4RRSC6eb0fWJ+aniMfK
JUfDGSlqehd7Sp1Kh6lBNAVGgFAwgZAU2o+HN4susq8W8jjZ3YZJPUDFu/R0ee2v
Tm0IoNVVqrPkgcKqLYEDhkOe/yEYa6w74+pUW3/00N86zFqD/thU7l7AHAHV5zoA
Q7VRHUyrYKT/btlAt51rs7Txk47j0Imn47jucAnMz2r8opOvPeMSPUlTF2OwFDrp
Og2/yzcTNlqNCd0stegYsNhum92t/fxpuPOwgfFp2dVreQpnSPoDgoI8uHNXykKH
6o7R31lhHkr7RTkxDQmaSWBsaumG2Y46haFqUz4EpfVB/RghE8L0PWefhQVgF0e5
Hfp8FNC9aEl8+zLZLAPtOIsAJxPhEhULaS7k4++qx+9IhH8ifHhDg7rGhZBkPosD
6IlYP6+4HDe951xrzNS++5YpLGxSmTXElTtKUqIARuYNepufT3CvxbQk79tnoeUw
tHzA5hKZwTtWbZmZnQrN17Ppx1q7H0aL7oOJi2MhizUDW+mbtFNN5j1rpGwXHye+
XNLB080pMnvphOjy7IQndZPnzYjztpSqLiIJiiUNM2JppdL4otpmnibD5dKvCxxO
qogyIE53ej3cHn/+M1V/PI/dy81tqU9RBKKYfcIOj5ofugF9WKxPTWzLR2nuFpFy
LJb7nWJa5TbY8sJGl79SNp5UbqFRRBboM/6uiVFF0PoAm7jKqQ4hzfNbyzLQNl0V
QIcbJWuI2eoEVZGWzczfyl+MlGlxgbfDE57GmAQtKA7k6pVOCVIV+QnaYBS1cz0w
3KxGE+FzgGekm4KLVKdl3NGr8OWc2fFTsHdNeIuSdtymR3yR7xVtc6dtjP1m0kxN
9nvHUVwm9bh1n1rw9oqxzbd/m6pAVVPG72yi8gp2NMxk0pbD2K0XsYry4nc8q2J5
OWfd2ma0dUUtv/mAQIL3LHbUFavN0JkL+iRnuf0jO4wE3Fu2pi8hdKoubm+tYvRa
pvKE7H646/SB1kz+6sSgeyBGsehspn3h6h94RyBYg6wv8L5SXvwDIkyN6pn0sPdL
qAmufx04O8XWDUdM3Cqbunnkx6mKjFydKR8LyROT8NAcQiB3uQ+8y4bV2ACl/FU4
he/Ep5VQIp91ocB82VkgRlPmssc5I0Jir3TasuuTC4T1FLj8ZM9/xw0YZ+2ZQfB3
F6ob6rrqwC1vKjfG8lytpWnDTE9DNqQ+rVGxXblKjCYfr/BsntRIE3s8aMH59Oi7
kKHlsfkJjAY2GYLAxvNFVkV8oLyJDCwK1FrPA9hH9vpnr2Ww3XE4I7k3em36WAMJ
B2jbsfe2GTZGArk4IXh7iJcUW0dqdzgkv0irB5aRHX6W2Cberj1uzw3wy/mbiLBW
cE1TR7rtB0d/yauCMNfenhYwMcgR1R1klIlXcdwrxW8b4ckJzVybV3lccK92fjDk
1fdO8I0LnM7VO/8DnKp05nj+vSKnLEJ6mj/Ri65c5TiurLderz6cJqblqIzhBz36
QauR2QCz+FbX/tOhsAKzYctcLOeZY40Ts8xzPF0zIhbnaJZY6RQD6g6Wcw03YloK
S/Ta4OZXGKfmy0jg+gT5gTLFmN5dGzWrJu+r0YTOYR5LycNrQEgAzcTSFnXcoYoQ
i9xSHQu7eb6TB3EH87WPmKXG0IQZ6k5tKbt+6IJt0LIs1FVVqTUeoANNaghUybp0
ssR8lgP8PD7NvzAj5iwd4sgWD0Wz00AFe20whHqdQDkssFUEPFZO45sKMzqlt45/
yaUch5tp7KpOBDRejYfhpgn0jNLzto8PEXd14VsD83ueXHUujZkWdN7jRV4/HCBM
0Z6BXFtW/Nf0mHPB1eP2yl8E+yswGjwgxELsD+WR20ixgSrI+MdNmw9xGceZqHt4
4Nl2XZ0WOm/4Ti0CIAUROd0Z22Fa/NEVwR7Xtbp9e7NwRziPm/J4ASb7ZuII5SvH
9Jf4+amu1Hq40ehNLDZtDdGrrdKvNrBpsHBgbzpJlByF+uilnAiNDBBbvTIXD/3y
gcIPJuwALV3wLAVIRBrDKzsrMAdllDYd66svSg1AopRc55Y6B7vutWTisNW4CcsX
K4y8J02H+VbbV/+ARQefLyBE7TDowr/E3w9jl2uUS66Fw0m6bBkHjMlyP6ngALu4
NAGu+ziQRXZx/VI3MNRm+j1D7fV0id/4EGeywdNwcN1JKRNa08FNXltsAlo0RsVi
sArmjSLAQ+O8icXlRpOCYs9ED4ftToF1be/lr1xfoGbfiUd+3TE73W6L7/q/lZa5
+XmB4+kgItzQSjubf4vuCq7l8tCiYQwQezYOHzHwFBMusc3mNYM/CwbQhYA6yq3F
GInk697I3yi1d4O5pyUDohDNlXfUpXUc9RDmiwyUbaVkCQZi4xRFnYLdxPy3tXh8
EZZPYtWtcQl9PGzkelYpfEZi9BVhZme3twR+g/sL9Ign1Q2mNqQ8/+p4hdxdFDKy
KsUrSUc1fQ70AuQyPoEkgS0064xvGtFbio7lDKq96wknuRA4fQBLLybSkc9Jw6yw
gOPmT59EzxosvmWWGAPJMaAYkq6/qHJhW9Dr8hD3DMX+Y8kZWyGMn8sRcRySgh5k
uGQgWLl5OESnGWRcIc5m01QXOYa8dy5KL9Qg4I80PBmzm3suBRZ2Ar7p+RiIck9I
cwRpyhD2oMov+bzLkHHhxSAXFnwEBmDOYhCxQULc7vQdnT+825xiC5xoUnBFNqZv
7mrRGh5ZP7JUyHGGnV2qQvycflD6dVM8FPe8v4h9SqEfxg2x8hw0mxCmXLlig9t1
+Rle1hBjv9w6aTly1j0QkdUgo2slRcwAqbdiTRimqMlNzYZbmOurG6KzxQLwsF7k
880OyKA5xqkKTtR0iiaqXG2OVOX3jtywpHMvfdEcISxY1GfzNzd5twwb+b/FcXqQ
ceG25qaEkP9upsUMuQjxTDqCjcjeSG3P0J2+iOcblhZenPbbwfUGBsLbAGk5lIrE
Hhmtkhx9n878ZXjH43xNgjW9GlMsKGortXdJjX6rVlcYekWTwXBvbZuzoyDQiiBJ
p/nYi7cvBmvTdAq87uyn4RkS8achVRVLlmvSVTNTML9UzPJf4pram/TuQteC8lmS
mVJFW6AK7buHhiKmdq2n7gfUXvhwckV7mMdkTJZevM7wWbAYFNHvVXXu6jHPi2Xv
Eq5Uxg0LU3v5R5iqL1glb8VYArFWporgw8wOA+zR3zhmTyvdvLW6A6mpWC8Erwck
PXUgHGJMyAUGew0HIAHJo99XGQnhvvhdcQopqTqyrTiyRL2pubFulM4eYV13d3BJ
m2KpcUjeQM/oM8pvUfUfoz5+dPyUPWUQzgmNXDYaPpMkkxML3sD5JeKa5ezvWPCB
kaE9JJ8Stw8MgzkSFZcEbZFbpmw5FwU1OkP+w64+2ddlTLqXKFusi6eN6CuF3dFP
pZStYOWFMjOoFwXojmqz51q5hvEcceir4ADmb8TUNV4QQIBqt4sPsIZahoiYl9Nn
5zkRwK+LmuzvYbeJmXk0TUMBAVbFpVfpV76/oswzSJPHqNUO6FjRyMl7h1XkY/p8
bom3A4IEJiDSMyyBxhuUgdw/LerjWn9UMldnNwk3249jj771NHa/WszsEslDCm0k
4JqqMOBbzrQ4B97URZAWdt2yyFZQ2VWj54+iWGOWZ1LYCee9t/w9dusBVnShiVHr
1QuxI8U206CRA3FNlpobOfsDNmDBkh8wICaF2k0kTo7P13Yn+JcN4/ZIKsm9syKX
uGQg7S0QlZ+2RQclvudekPjC76CEXUA1kBUjHPd6gKn1zKK/oYQnjB+Mk7TCIYre
K6StM7M9mdP0eDqVDNQEtUx4q3sMWR3Rj7uJPdH54Vfc+zAa1ZtFdvfWk//IR5xg
rU9VZMyk+BKFToUyvPy44SuduCGZ/S1SGfYUvF+00psBrYtP0JFwYRGu7+VLmnPK
qa1pe5FBFo1QiroLWkcR0zWWa5eaqv8snGNOzpNjf+Af7SfUy1qHAaoYJRqqyfTY
qCffjoKnZ6EqOUiAYhMc+7YilHjUjTVqdM5Mki1bWtkuvugOdHTZlTWabcatB79h
61daEEPxOW+zIvviNry1+x1h3sb/gsDM7GXplYMNOI2dQApDdBoMInbMx7cR4KNp
wUwD/dbv8E6VxKRZn49ZU26lJrcGPf4DtCln3WQUZDxUjHCh617xmk10Sf6m1Tgu
+HzQx29DBVu7iQlXY0Lrh8GKFUwSCqECmB613d5td/tX4/4DjpV/38np/8Eec+rq
+Y3KuBjECVCgZ7m0emu/KLmcV3ImRro3URvKLTK0akeNDoprvmkypDkgfiZr5ITZ
KurlN95IMTxyaHpz4Yw9pY4QNfTOMJMeTT0udvpqoWsu4TH+IlfV8KeCT5Tw+ert
XxdD9lw3NACrx0sPAziOKI1R98kr610U9VmWrinewkbk5Zl2m3qLK6GjeMSCt+sX
gkWoegcodmHafVIwlOg07XB4/61FNtHmRDX0lz3SRnO/L4ArZSb3bJKjsWUDHuUs
UhbAKmR3hudHBA3KoIsS8Y19i195Yw+MSG/h5NouPBI3AeCXoPybjRJEdmTrq87E
qchQYkBH8uL5VO5dmay5UNgSjS6iF9W208T/Xpta68kmrFeleo05bu/JfT3r+Vyl
3yYDUxa5VtBb3EZ1x5E+bp11Q911ncMA94NQjmQTveFOHmqezNFZavXy1kmB7QcT
cbJufBzWedBRYOT6UWDj+hs88doanW4zVvj4AXBcGIXx8u/9rNYcAfko+lhgAsqO
aJfTHuDjW3hbp+8kJ/+TDoj95oG0wht9bTjCHgeg0vKMsVPJta1kLEou5zJfeuTh
EVWQxE6SwIvAl9GySQJXrRWA1GMWlUzBGToMlqcwKi48jIt/kGfUvKvgxX7AWs55
1CoEfRHldX20L5s149Wfc6z2l0GxYtFCCfDamxMDO1wpnSPvcp+HAo9nSaKe0Re2
eUHfijIH+Xd+ReDGG4PDGYk/quVZ2iOWE98Vf0mL1aa1T13AvWnWmkRzvPrRloP9
X0J8Yckr6idj6muJUnnIs41o3vYoLKRg7rllQ6k+AxmPBjlotpunhyzAb5WWOw64
EWnyoYG51sPu+A88+p1sNlNaN94xkTIcngS659GKyJEBH67Rq2/uLUkM/y1RPNHv
wUiClAYsc9Re1VOPA5EMNZBiyMCpdnY4ucn5AFGDeoTfkC4lUTzPoylwoXZnnsxW
jaSVZoSbNdUVutfRUQFFb04aNn/nww5byJi/cydsWbjrnm1+7RNlj3eSKI/jM+nk
DYeR+gIj0l7aNaIRQvow7fvOoEy+fFf7lLMOurN6Is6YsugS2YkYwMVnR+7MgARq
4U4RZIODX6Dwg/hLXCGjOaWaSfj+wnhb3WxSejaka0DS2WkHpghzTtLc9hGYGDrK
MhK8Q0GI2RwwI1VXZKkGZ+O/wXnhjE/weL3g2qbzdUPBjbMgeJJpJUgOq9MelO9i
rOlyLyZQCNM6+YOSNOU6kSwBCodz3aWNQQ/YKRiRIKi9Nd9jwzGxP2xAjTuSRK7g
8Fj4RO89TA/fUAGJl+BDP7Avcn9KM+m4V2kdRwlSVYsD4ASah1wsgduRCWKvAiqm
MQCHBnQuauLO93D3sIasbrbEGnMFg5xei3Lcg1fjavxOPLYxJR8L+nkDESiKzlG8
/sWJTGDmVk1yCgnwIjB0rmC8kwVivvP3SxxUtotFrJLQM/URw2SGo2othGfPP6nc
tj66wWS7Q3ii5vKesM3TRXY6AmWmTIb1DWqFyJRmR6zu/lK1oAlCMB5cGx6ckFvH
EnCZsuraN1ZGJqpK9Z88tK2IEHa+VXey7KUlVsjQGq2Dh2a6Fx2InV3c/T3Pt33P
v92lj+wF8lRPXRuPbqOGQP9fd7t/LvEp9+O69A9ZwXcTdyMRRck+SsTRfNT1mHHb
MNxtsTwQUYeJaVA3sBi7O2HDML+nA1a2l4AR4M4zLBCO3jzH/VCDNRnPCzLJW2tF
0DQHZ2eOG/q33QpUfQltbp1VR9qn/O12/sxayOQ9LVfx85etRZgoMTlGnattQQ4n
bEdLBrbLC7V9eWhHlHINAQ2+mZihouEOnFZe2d6dwz0GpanZZkuM2drloUOhQKvO
ovv0YJGGY/Hpd2hqzS09i9uPAtZ4EeI15UFa9mSrhRd00GtaK50hrwt6EvhKTSPY
TesBIv32k7T0YphYJPVwuCDTKdcb+un+o/ihDSFC97A=
`protect END_PROTECTED
