`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMppq6J0XBblzXCQi7cGCuvZOBsoE1dzRzDzjRNJvni9
yMY0r9HnZlS8QX+8Brd/FRMkCIeKNGZ6QOBp5Co8wvL5IvAhNZfupTgRHf5jM7SX
F0+w+fyHG02btZx6bUH5XWJk3fi4MDgX3yyynu1W2KTGm+BfCwEuZit0549AswjB
`protect END_PROTECTED
