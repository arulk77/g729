`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yhrTyGV3B3SwHZP2HXOW7MQkY2Bb7v208QIALkEaGXT
e8ynLL8oFcJNgTrkEEUZ5OJnwEEWfbGcM6BRdQSQ5rAnfPOReuXj/XiCjIWWK+xv
RbNeWXEC6s2G1tQ2rl1CphSV/TbBygRyI1rNCn5zsFd8MBIAXqSFex71G30ja/Mj
sIUZFku7Ja20BBri4jgTvO/dde0WbrcNes9LSdvIqpRlx5qM3CSWWXj6MhmDXLlh
0b7jAEudvlNVN1z0v8PO02BC2GzXaOO2OHk3dVGdTgIebMEUkaCJYuShtnUqJcP3
YVBpT6lmUPlRlIr01odnP5UQGI8aKFmFW18TL/P601odEPb8ydemtuAd7Q0oGzWX
Afu3B7YgechYNXI9JHp5W0U/biuHOTMApgV7qxG5VIIw/EiCj8Tb7NyxdC6nphe0
3LHOY5tU01fMTQT3aZvqjQ==
`protect END_PROTECTED
