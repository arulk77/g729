`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNzDr/0nD1X1lNWO+ueXmK9hapdOW+i3y3apNuqGt1aYm
9qAx0ijTHEQOgxO/exzsH6zbB+ehoEccnaSlIQGmUfdIMkgGVs1J8ztZctZE2NZQ
+nuCP6et2Mqq3yCPj9ItQLEhmKRAexfLzjAZpdzOfqzO7GR6WS1nMkUg2GtNFuyM
ybyJjFfTXNq4xSpceU7FHgDHU8PQpQPjzm3uN6WaEKBH5PCORpIts00YlfdyQSPI
9fpthCnDgTOeNm+T6naDwO6+gZxUk9Leu+y1wM6scbKNiBgQbDBr9R5Qnn60wo02
sFVfMQw4f9q11Al1aowml+1Yeo06TyhLg1+IQ6VjtMI7pfprOtYt1gYUDk2BFRY8
70KIJyafgQJWessBHD0z5B8jmU8qY8m8d/m33aVu70kA4ppDDEuetHpnAcOQ0yL0
d6CZzmGLYpgOkZtFXuxX9YAPdxGco9MyH0mAI5lHGp5UUys64Mc+dBf8lqKaxs2+
S1vrlKrA7fnI7gynniHP1VWyV6BrlylVXN3t77z2ue7fQXJlrP5N1j5VNM+AX6D0
afZr/ek4lHvUIXEfm4aOy/fzPmsZnIkdDRVhay3R8sz7vlD4xPDS3Ly9HRHqpVEw
XuWw7PYVE8a6Fd++dpk2ZzOfAJ2mpq55nt1ClMkQpFUBhq57Ueyp3oSLup4bHDd/
JzP9IJami4mDz/XbcYQQoh8XbF5LzrHMuRulyaSJuiszgrefpuPzGiCjP3s2wVrX
LoIfOYqSX26SMxh5JqBymMbgiuvwcZLTwaz0s+PfCy/BlBJe4eWHw9WE2G0HnRcX
hKr+cT0E/YgNHnXFQ6P3PGnVNU1ofSjwN1r2+vALG3TkLd/R/kWKB3mDhDrUSlKt
Yq78WR8VWO1RIEIdW31Nnf2O0BVMZSUjvYGfcfy+FNt1dd2RvPQ3je99cN5ffObI
pavr7NH4JBYHnp3K0dxkNfQ/ED0N/WnCKJg0rBx+i6e1x76dilPoNB/YH2i1ASsm
Ly86SqcPjfK9e3JX72DOivEwpRktHarY9Jx+3IE/dJZsyAY8TT8xGf3fCT9S1uan
dhhF2TsVimRNFz6MK+isn9eIqJv1qs4J/e7ue8XlaK1n/QeFbhFmsosz4eQOYFtb
vaxAfQV4uDOFcKI9kKUqManrunVTsac47Q859aRhz7+UYV8A3Pd27cLisz21WH5U
MW256J9bHbgp42+/lvQtT/PeYafaVDchc1MSOgR0BST6SnvHBqBO8iyB9ZWlEsRs
tTF8kfZmIHwbxiN8fLe4I6LaiHUZoz/MMZArGOOndB1ebSXwYQB1PI9B4Js3sDa2
A7eUHzCOwE7EmvhHDZlP+IGhZKNLbAaB081MaBImAYTZVEt9CXH1kGYkdNw/DTDw
9e/+rgWUz8p3ZzF1atwBIw4D2v3YWixzTFULq5NcnxTOrpKAVAzDWxpXYNS/5kk+
oSVee6fm32gUl5Y2CTD9brefUEScDwyNQLIWEb1jJ8UBHvWuuu+vHIFXjYROjj4w
dhHSwer6XJ93ctREpLwPQ7sJZ751YYhVrUE/OzRb+SL9k29RpE+ACVyARLR5t5Sa
E+GHjN0Dtc4SFtgW+96SlVITtnv2q6Ord6/2IPA9qSyzC5ThsjIwm+ZvZ86LP4Pb
EirEAh6cCIM9CNOapwMocTIh0GGX6h3AJNGAxyhTTBo90Cr6kDLPsYYKxrGHEYdu
YOF59FaEAxDLnRp6OqOB5OJpTCliiZ9x932KbbVzJSrtGDME8kkrumyMwgBTqy/R
sTasq1lKvqAtPYtrdfoB40UiEKLzCsyR9C2QFn7OK5fnWNhfn+jV58Ewu6ZJvWeG
TyqbmGFl3a1bL0Km+j/hs/sDdqe71RVhcVxb6pU0HzrtrmdjidgaJAtYyQ1UBE3+
gfA9i9lrA/slmV1QAEhJBFxramoCfWPWlgB9yH2rz48amstVloVcBX+wL1p+zitp
gnV7yc49AaEOab0/kEFLa+PqJSpseMqMgimV0aIeH3IwAUXo79PkXAGdKSWEp84v
JJKqIblkXZp3LcxHoZ7IuL14xhN9GiFTLqcPIUkPE7lnWog8IGFmkuOgyJRmLvFt
LGKV6Fe0NJOwdvb+i11rLelP0tN1OrASc2FHAoo9JEeRD/sBAowhw6gQad25NRmK
mjYY0GzaAihcJSKW0Xu4UtgyG63N0qg/JVlNMcukgPfOstxz1Sl2kbnWgGAVb8LL
DBD5wfUxn3Ndu/oBZoViRYGoUfDljRf3VxpgKrtrtyE6/CiU/TIXqt6TmK/d44fd
AjuzCyFku15VBtXenmj7F9V7is4NPzO0BBueGS45sdAxBLjx7ZCagWoHMs7EFfCZ
ht0JJ5TYI6rzcPZvp7Zatti55uKdRINoUNLJavZFNCe/OjT1DgfEp4S3G4ydVLME
5NnMT1+jne8kCa8wmDUdNv7L1W7E8xSXyLXFxP4EjrMbKfvmRa08LiF1g3di2wcM
gmjoU4XgBxCXz455mVxRANiRA/FrVcySeyUGsOUVNFMTolvR9G9PuJ3egXyaLdW8
BrfTj9fMY5ipk5tK/fVjn+VDYFgADnUsNh3ZVQWXQTc4xRLGsm2Yn/gxOvkF5Dpy
k9plnl0+kgXJ1MKqCuVKX2QX/MErsbMEWWHwZj0S2hLOqkudxKGPAq3mLJyCdhXB
rZN8l4hEUxCVbb064eF7CHayI8gMI+P+DkCeX6CTJC66Oad0VVkROK32TEPG6cxu
CFJ9phAM5DP+pCYTHkWxbPu/8qW8lUcD3vbY6MqAPCzQg3/7MJCYw9mLn2m8oZ6Y
lrd+FdqMY8zwCII5RcUgc2eGOCNssGLaCUjW+YgntKfNX4vn6g6ceQXFloofh/QF
oQdxD0G3eMnMr4Y06hiTxEsuPJOqmxjCYwzwcpnsQ9UnlIB1Ey/BPnxvI43PeISJ
RFN97ahOAh/yTBr1PDAqpiMDT4EJCh5CzrntHIWytg0QPfrJfS0f8JJkp9ERvf4r
+cKH0EIn9d8P04zjoI2RW1VjRmKOdz3qgE6i3X4vCnMWwZ8qIkaTA3KV03KD6VD1
jGSju8wtogueAN1P97KnN+yNoPj8GCAnGNKq8Do8j33FiLf9gddwTvbiYCW3xPfE
jicnMxbPoh/wzcW/4T4B4IYCjL0VsQc/tqblmZxwFczezfzDcZVRT+YLOePxRAKb
wd0tPsWeg/8ntFuYaSBUAGDd5Dpk99z8neDIjRmol0AQwf3MxNcjP4Wul339/89S
Q9azmoTuIu47Ma8EWbs/2QNp3qNaZNR7GilYP3nyNXiaLJ/ieEknu77PqxKWTzfH
JXNThv+7WI8YThDw6x77dzPG1ZjNWP4Y6MO4g+SASoVduArNjOcME7l6H9mbqcv7
Qp2NaNuBny7aZyd2gKlmm6YaOQ++7hXiDI8gWWQXQfLiZZRPpg1loWn3kCNjftJv
UFAPdzqW8YX3i9JP0EiJjB1K0MCrBgP041grkIxEuWlrDY3ZaGQmDWUv9KHST1zU
8iRd/LNy8BQHmp/1y6BGIbd5K0eX780VL/exqYlxYd/2yA8lCrAuglRMIQuBL0W3
rz1LqaOLWy5l2X8XyvVsO+cEgHjqODRzBWWT7ddVUD46QecuG0LAxaNYjamW1FQ7
0fZkhaaGij1DZfZaSGz/EgG+b60yykrr82qTnlH5zA2chBc8R/HJ0pQUTsbH+iTL
pdpx/WLlFmW9EK41Ee8rQ+YtgRgDGUyUGyeuOzSBcGvaDQnDT2XDbZdt/NNc1yce
U8WJmOZvqhluCezaMLEXGLQqoQ18K0Xjq+pv+BWG163nwghhRxAXiKuCm11eZRkf
RXu7A9OzVd4gTzMeNmMlOH8LxzufwTylBZuAdc4GqWgZs6fBW3Owp0JNi55C3YcA
9GV9OOfNMaegZy8zPLb5iRq/eMfJEjENw3zvsnx3dFNeLSIaUWYMoxcQ+EtKBdQ5
qIt9fBQerNY/68TtUl9AsZetotkMjdytDR2ErSdkX4NNXJKg9wn/J7ZThCU/hOvX
rteyHuTyjrChMDZLPf6XCIUkAN35GKj7uwK82J6hrkHQKJtjwRS+eQ6k1f6+3Izz
let0vu2Av0/Js0ObO2VCZOddwxYHIBjemXj9chH2Iv76xo68c9g7ppQijzDW5XW/
fUNlxJUjfG4E1EMYmFqgSSv9zditQ+Maz4IzFcBCYyoeBRUhI3cneWeD0rB7EaaA
teOS0rMk5epfwgCLO6FSb0oW8rGfyrNYLukqowY5GqApzFAhDYCfy+33CzUgX17h
IYnNB+v8mNzzB1HQ7qY9u+GY1dVxGwyK38QNvTrNsi8dnoYFxqdpOfEI2f0P/nmo
eER9qTHqW9HpWVJ0hNiW0VkQ93DdlxlnQDU6bJPkvBkAofq3Bc0BTApcfUP4fnOd
EK7/G/PxYbXccrpAb0ke8NUlaVVivr4ahjwssZY37811ndONlCpyEXr8De2is7M/
YXofN8jIFM9hldgAbFo5GIA6FqmJe4OvpcoF3CcQU9F1X0iU4Nkv/J4abi/R5Szx
ZN/n9fvW4DHpl5KmdY+N59s7ZU3gydAF1xwjFVY3VGRlM3t7Vw669CSO58AX2WSw
aA8Wrzff1u46vi45jt5xUj7RxXU7/4AonzbGwVBT7kfTEXdyY80UJY8vbPOHshTu
zsD74zjG6A3dNLH3uFrdbEhLUyFgYt5RnHGgjWdD3xJdr1UmcsHoB4ZIBLN1HvvX
pmJzQwnXG1kt20kAUSgEfhDcPD2Sc6EU+9EyeCQpt1ZUns50J7loXFOjHeiu1+TH
zL9AsbKmq4irkrSh8FB5Pg8HnUK5nBUlHJTIjnCnDbK86AQEU0t819nzK28sUhOv
x7V9b41Eu10vSexkBWqS2ALf/HIhzwLH5sEyv95z3PxHK586UU5KXjSIH/JoHnuc
fS6kh9AhO2zNdtCzAoCc+vcwuEDile3/lBm+2Dsp18WwHjVxqGithOtSpyo2UHcY
RdhqKVXQq2yHSxtTTpbuhoRi1zCZPgIEhdDeNmYFwfUvkuTf1nJzAK6X8ICV+k19
q9KdCXrZp53jB6akptxtZJ1A7a/012+Ih2tZIMPW4A7w9bs6nwCKTiia2EuCJoQI
zW5ZMqmTSLBroTQgBq+jP34phX9LzOv0iwLYDN2kgm9A0fJ4yKwyW46RXXaWKHPi
j4JjYkV9hkRQr7jiOPP+LecGgCaRzqOysAU2IMDkLr8fU4kgW99gmJIQBWuf9gqO
R0tXhSR1x2LAr6ruzEyRgHykMiIlykIs18X02I2rn7ontODiON1/06CGqptokzXw
aLjCzby7Ktr8Y6Ul/GsrGchfKq+3wHeHDqW6dgYVbD3ZIi/66KdP0VxPfIw7QEQl
jX+ir9IWn6TCU0BtbPXqprkFHJH+mZYhETK50iJhmMsYspgHzG5MVtmCPpOiZghs
Gp5+aeNq9L8GK57kX8XopjRV1947BbBVgR1szWDTGS1Hhw580BZV7p9TcgcZVDce
tCNnkd2L7RE025ctb49jdyBiXyjUfsKWw1ljtmHrEFDna4eVBYnQT1g9edVC5vdZ
MZ85b5OC8pMkgYilUCwYV8IHRS6hXFXTtlnRfie41IKZplnE6AmvwuIKlmeAb3UF
2wA10mg25HWJInezfXRoTw0uU+R7pfBHMZ7FLumDcJv9HjL1zJ3AO/lgtrwKUb56
ehybVhucq8HG5fFRt9rYnCneKIb5v29K/b2qTTnRrkhoP1DX/0yfW9Z9RRT0AJON
bZX6GwBRgzw/iuzxgfc0pdIPUDwEkW8oIVTPnkSuMinh+k0UHOlvcA1I1t1HS6YU
qCwyWV41CIhF3RjJio1etFKaWFbCTUznzRstfTOBsimYEqg+/+qRmFNxVOt2+YwB
mhqY8VdqkHvh8K0grWsyfRjY0ZnAmi4p6ylkKixyAL3rs/asPYwgekEW5vvCLRqM
JFddffLpLvSG3kO0tz8rdo5UiO/ZjZu7pOWpZXDHanx4tWh6GMuRCgU3opJNfMkB
M1k1p/FnhVPHslMRNOvL+NhAfmkC5MXSa68efbDNHmvvis5oAWcgTP1LrmZFL2vy
wZkDY4LU1NjLUPwm7BjJhJoDasBgTIFQ39oXqLGPtlqJQLPeCnK0ZT5WmKTpqBkw
8pfoIE0J82QpnmhXALachxhHRBSCh3VIAdOrMQmaCP4qkhW6sLApNEelDvRlR27h
cnSdaqVgEqiVrnffchajj4trqjcUhJ+4NPj4yhuuZZFpNnuDV9bwOsb7uyT4rsi4
PMiyKy5x5NFBotSm3DXL3LW1woiREtzOgSUI7bctq6RDGpGJh6DAbRaGDE/KcwKy
UbPA4OWa0ZzQv3IC0jKTY5Ln8c0tQ+wrdTIKHLv1W7RZEGYwCSgrB6MGspIQRirW
RS2i+waslaNGgB3ZcFJ2tiPz75EkdY/a3olP0XXIzXd37Ma6hOYnyAg3/E/QhkWR
EdkxRxPJ4WNt+p/fCPdavitdQfYfoWGmYZfNOpsV5PtsHXrj0U5E4BZIhyq+53lK
GqQjlJcjDhTy8S1Zb6mkme88yu150GEpa3hrv+Rma2IVoEL7dNacoRA2+nWqGu65
F6lMHBlvbql0rxs7nhMysMdlIak2/Bg0siQWO0buRZeZwWLfRgeh58tJnBt/DJGR
WTHXZr9v6sTZOXPejyui4scSH1Z9x6Idof1y8aH0cqknGYak7gFDhbvynO/MMKbJ
wkIucuvwcnUl/WI1AEBfAC4IMcl/5VutSOHqD8wbjr03W0w0c7wA+L/vaTPq39zV
4A/m7I5ikrXCSqTLEeXSaNrZNfp5XQtjk3TTlDwQ5vcecY+fkpv+Y1SIwIh8hls6
+2ILbaC+Yig2by/ezHWKwY02gxSIBeUc1Id+deZtZzZ+CCcYZt7puPVL2+hGtSKR
wH1vQ8GslIBhzAz2LTU+DN17Ty4yVWY96idGp9PBjrQg2ndduVbPhlGH/aFvxNM9
jLnpdGrWz+gbW1In/KC7wWqqb4HRHvoXr28U4BlXxtTLZYK7fKTx6oougJ6P+27X
2HUx7Xdik/aRmE/mQhuKebHr21cqMLU8SwmwAoI/shS3SGrFEvBg4m4M7PBBXY8j
TTcH6NRq9gMwkRDqoBZW/MxhVflVNh1hjvW7KC3++syeWnRHAqxg4yjPRSHe0mq2
/WgWhVV5lORiJSs9pbqnS8lstTb5RQdauvfN7rRtWVlxUXcvr1X35+OMoSq+yrTf
S8cnRiwnGPD91DkyUAAPM44Eq4gpCHh9aw65QgA6qBumJcS1po6xI+XCmvsVq9DH
TK56RUs6CZa9X3VWC+NF8ZoTJGTyMDRaZh01CCu0cm69IA9ge1HPtaWTqG3U1G+0
Tu8XeGzqnIsDnxu4evyfqu2lnLFMJ8RCPqx49a0KUbovvuRgznqgbPyzGk9titlq
zyvGNnUWHySRYMP3bf5uOTdjADbC9TvjtQptS+UtJtgcgTnXPJPLdCUAn5nXeCI3
VRYo33HUcwvO02HLQGodQV/SFx761CgOKYq6WX5ZhxAMQNGcqYIlRjaVpAKu3T8E
MLZ0AtuE88SUm1gUqlNtnFZGS5scWD6eqdr49gryV+M3CCUcl9F0a/uq+NrlI7vx
u+VmgVeMtxqEXzA3bsRJ0Yst4d1T9ec+KA6GxqUaBUgLJYj1JKNiLUX8OBYbA5mc
1mKmMMhPV2pnTbpfm9yRKP2SIE5wk/dMYmJ2p/F0O8EskLyjDNodd7yuXhWVwdy0
Aw3faOMpfflGyiSiWWwkULSG77upuDh4sa6c+2P5NQ/z3xMacLsypz2VtwYVHSNS
uxVrZTHQG4DbDBBHD8fojKaPvjdk3spC6rHOY+q2n4KjPsAqUj+OJn/QIcXihurt
TQva6gAX6NC7vA6pEGG/vhqzFZoVYzN5z4fpMb6tEyUaCDbBD/uKjwJRCbhxzv+9
cdPv4o9lzxHFus20STpyyk2JSIohtXKZjK96qqIOT9l2fX7FThYuX4DAaY+oa9K4
hfea2B2tGyzDsr590gciFXMPgRftynBxhO6cWjCY3sohMESh2SIAMy/GLdp8pn9o
VTNoAxWt04EOTQBUQYAWogeLyadOVEaPeds13zopbcoieBpH1vNHPBFMhKpdCwgj
osNdGRzQy2/enk9V9e4wQFZHz6Ola3SzCrjVOt/ckIuiqOx/VVe27peaQCAupWyd
w0ElKgG2JO6VU0Uqku37l/Q/UNtHBnlHN0CuqzBjqg+a9SmSCCnWfvePjdfUVd48
o5Wa2VDhz2IqxPdMlChVGLMoCn3m/EKdaQQC710pN45jznvelKblQXTsVwmJ3nZF
0LtPEY6gVlk91bzEaESmqmlucqYgM51izTPAMHeeXn9WpsWjMHordfnl5yE0r8zj
Ay90w75VIUl0Fbdka2GTAed+gktP8W1RUBD53CADlkLkFe7k4aEQphs7KUJ9kOwD
sKx6WCFFpPU0n28JsQ72h/IIR9hMfNC7ZKAVx9wYclWZRB3vEcJCGFGfyIrGwoLD
skVple/aT3CGBVTYNfYP3SGAD3DCdGaL9d8pW36Fi7eHx/1NPIQGJlpWnzTca4S0
TkEPZOvretHKpthg4QkJ3bNYlHVBh2uUAB9VUh/twARlM9M8uzjiXC7BSif8hakE
8yqSBR8eazFRwRtnb3g2UoGHkaW9T12p7zg5xsvTP4V1SXFA0yuV8BkXRLhAzSIl
3Mbr34yuFVGdAA/WovTxVvPaFFNHOui5niRZzp6SOO0tLxBB3I0q2KojAvsTaD7V
wa8OLQ6BEJTbPJuzCnI/B695hXf/0qn1abxE/jwn9+UGTOg8o7hlPQtR1Qkuqu8k
vyeeCJ1PtP4YbzQ+wo8xfOpCN2tVO7+eD9h+8cHkDIR15vvNU+rpMwRFiHJy4MOx
8vjacreDpMjHJ1E1Sk9kPTMRRvIeUPNeTvooyLyAGeed2xrYK/ykEl0Tvl2IP+Ne
RAfZv2Ln25HkO27z0R2UYXlVOYm+rKDBZEUvmOLnacSxTrwPYBxaAc9zXJgPKfr4
0y8vEsBxSy9UlKHiNMgB8oZPyk/15ASUXEem7yk+vosIcv8qY5hxDw0eW5PuMQGy
mB42Nww3hBIO6entOI/KV0NyXlLIWs9B//uq67ZeLsoaJe2wU1TRK5XX6N0IMdgQ
eW+gji2H2yKlgzbkfPaEdF1073mfrfpKTvsu49InEHS89/ARgjdc9LaV9nqpGOLY
sy4a4lLu0T4x81/Blka8MhBxjw7fEd4kw6AVzTr6Yf8cDcftZcaLwSyYY5JRQDOH
c7XdGxHpdpuPS8VuRfNDGNANvr0GX/5TZT82zGFI/Iah9i1vAa/GLIrf3U3C0jv9
2AJxU25z1hzC4Zx/MuFJz8ORvQkufUs721M4hYC8yGCgo6U0dQma8UuSBofrJyJm
X7nf4jVGcV6zbRhd9/GlSA2i1bcz/59HhTi8QEca9PAjjHaBdNe/J01whmJ19Noh
GQWz7W+J4G0WMw++bfwYXwKDd4kRACIAsx97yW6+j4sXpe7wSAEL6OQXLe0Zcc2m
6yJ4cIyKF9R14rbTeGAp+unjJBpSyxwIlhaglBftZH0OhFI1q5A2wUWrHcG5joAB
x/1hRuquwC/847orxxBDXhZzSXefBc/G6J30W4qnvQWWO5KDuL8OEVV2kIVwuQti
e3Rt//ePKO/m67Tw583cXfImxzaeP4QGJaqab/IEiSXtneORFupqUUYRepCVfrYX
vcDWUhSBMvchTYBh5uuGLcrYA37wv1bGQ8wDNoo3CETGdBvb+doRe4drTniSI/MQ
7R/Fh2rC24wgvSjq/XP0CgJJrTQa4DzqoazIJmR+whCFrQGAM1P0Lwdilf2nrfkq
TpuK0jJGuKRb3l70yBEf9ALyGnwVJ2UPq2eqC21v6bIj0UOSGjA1uQJrXMTNGdrL
PLCkWnzzOEpHZT5OdiisbuLyGbogovFoX69g6pQiE7GyBiCxg25efQW6qE+dmxys
Z6pi5Ll4+ulPd9PXcW5DcQyEwQU6Mp4fD78JYWedohz3Hw/illSB2+0CGJKs4++O
kFGvY9StTJBjndemMkFmjorNViQey/V0OsCdAHgdhsZJIxfdRZLdc9mxOARIn6BZ
+rhVIrA+00gur8uO8lhi4UyRYGMSYLQb7u4/U0Z3zs23xylMQg7GjN/e52pJraZX
oagdb1kcsq3slZCsRmpaYTqCVIg8gqKbwAOAdELnf5fxTPSykl9b7kNjTZYbGsAQ
mjs3NNJWwxx9+ZFD9U5hozA81TVu59yM9/Tn6pCAuNcZTzo06yh172xwJ5kaNKbs
AOTkDE9TYFqaXC2X65gCva4DIPANlTnAHsNmRzP+ZuX+xEMPWEoRfo4o483J2tU+
LY4rGPmnCVWnDfMPRatPRKhVB+6c+Srp5rtlm8Qdetv/IkCu6IljOrN+5aWJZ0jb
c2SI7cJixxbI0lrDLvURecvMpE7qZNA77MHaarvXSlzT1JUxBn0iu114FXG3PplC
QeI1Jb/7iFv142ggJaxGs+J2yTGy/YGAi5/LGItm5ISYyxbF7G+FlucFEMhSUjBl
LrsfqFeFxwTQjWPhCejzBZKOQT6puxS5m+I6Ul8vejCH+ZCL1ymNOZuyyC7I3IPr
ke+B+Ca6gii5sSPSBXzd3kCy6KPtxNS7vGw5m/sb/ikNQiXtxFLA+pK+PO24PaGZ
8azAqt/gZ9HCAfZIDeRy8LRm2gCV+hJ2shAC1kK7xwU6/ffOGfDOCDi87mgWe3of
lVQ3StecQoyzcjS4yAeTshgANIy4uv3HEizuZLgZnbTKl/b9XumphWXa0SJaVhz3
1F9Ur8WZ+mNKXnDiuN1C7IiwF2KeK6i4/Vvm/LGlMle28PIaVPzTyC2abGQ6sv7c
p/OtlqUPcqfZnSz64yiViKns10jxOAvObkyvQ/oBo5Mw8+F+RjGzPgXlyQLNkKIr
3n2IiNX+hm13awYAZU1nOf+Y0Txp5p/PruwlYD2r77W3wcOytSsSHS63u236evgI
rGFVmm2LuC+7gkLdc844/yxtmi8GxZR3IX5hYhoz5AWJct46lymgXZz2/yw/3pd1
6mXIP1rcYQYl0KioHdUkOyQ/LktjHBQZmjOPg/ygS+5lGBbPkoVCtfXVhA1aY3kd
CEXyQfIcVPyFCZPw3aUK9475Y44AQuN7SUmEXDQjPj1zOWKJypMBjm07J28k/6ib
UnGzQRsiM8rGE8FyIvr0J1tRT8YN3r3X/wHtIcxrkajm/EBrrffi76thW/eNCt4Z
x9Sg+pBFrJU9nSK8XyxtsSuqLbnrRAa7mON8hh23kjlLxAjhBcUj2v52420llLXC
k04y+I2nTqfgO6PmOdr8eF/7jfOwxLyA6WH1eQqf3fxg3kWwiQWt96kbetPCTHDc
Dq1fro6iIww+aX+SiTwl20bz6kiN7PubwX0N7Pd8vebCUCRfOB0F6UefSlkXHn6x
lrDjR3u3VQQmOj++5jpbr49b8DnhCDgmv2QIQH3umxlKCbrAqwiYFWImHQi4Lqvs
O5Ggd6zmvDBOgwLlW0hFUMdn9VNGBi5dY7g+2jCZGhss5PZzFY+RFeq9HruN6kdX
6aMPI9ynXKg0Hn2jlHB8Vv9aVpuljJAVYiE0NFBnPXMLKW2VDkf2e2wuu+YppCp9
bfD+La66+mTl+Q5Wh1WjyF75JmYcZDvp8p7H2BbPqWKxB4u5oOT71f4ffd0GcUGE
LeIMCHeH9jSYd0Vso5vyIRDzCeB9OC7+vzx31lPih2Wx7e8vDEF7ubkcRlq2CEuD
2NAhjZhz+N0LZ4YneeRlRvpgW+NfILreK8AFKk7IFK2lrxex9zTMum4nTI9tdWqg
I49Fe22k3VnRaAUOU52zyTpSA5M0mC2lk27MYnRSB8AVf44Ztt0Mcl6faFQUoXeA
YNRKtEAKxGCz4hPUJwompvmXhglmJ0NRlMfQrAXahEvMxq2mkNBNSnbw+E1B7w9e
Nu1DHq+zObNmJWEt8BXnN4+BqLKgQioKJxNksxK0AUoJXL7+fe0PW+TvnqyURw46
whfPe4TuBJ9GjJiEdpgMoNZ1oXSf5z+qcGaeavGTbjUDHHlbavS5bESIPNDXhlcM
6x7CIVuJwWtVLU1WkSkbeJnz2pCHaR69z4hin9QN/7lLjiJC+KLgkOXFvKvPLh+n
wnZAGLWVBgh0odcMWyjVF/JW9Q8JvDeh4l2TeiF0+EQ05/5SkRS9wKW1VJSrGf9E
o849s54Bu1B7uTPtWCr+zi7hOQgP2UTxxuFSA+KWOtj+bMrb8+kzkolcvJWUbK8m
phFccvHibGCp4ZJJJo4W2oAGYd46IQKLA0F8HzOW02x9UzSSm7hbz6fWTLx+LBEe
9GdoFZ11ZBgnga5bpECheOE/pR6mNnHZ2Ah+MeY2IM8utixxNy3SCZD/NrXR6ihu
PRcAEwtpuC9KREq1yB0QR2Aw3fvsFint5iQAsvLDMpQ2U0nhiWgRth73i+dBD7z1
E694DTPnYTn0YDrdSXekhSdBb0+gVzan2KvufoGl7nTsLUIKEDfYXZdnmfWfhKwP
G2IJYIkxJnvhvZOQix6Urgsw7zjyMZk+GlK4h39KZ7CilbNUM4vYCMv7JAXiZyC1
q7pzYFa5HHj53T2ejDmCX/Ca3wIxQXy/fnSPi2D5xIymrFEW/rN0m4VVaqP+2dKx
OqEnuabpjfLppk6xVSXHkyCSn3uvLdynT1tTv7QrlM3okXpNroHNbKtc1/0dTFEh
X4/mxIA/nCXz2YxsBe/xMfM+RQH5FmCaahdkdxqpKyaPEEOqQt/jmbyAj3gCe5Ij
41m1/tMJ1rYhdjbmvKHa3+4d9p8bhmR9f0zo2O8haeco/nuz/IjV1UR1TSy0V/SQ
dERE4eOKA4VvBre2MNAdBmG4mglbVqlQhrem9Tfah/CK0o/pgF5pspGyB+zjDSsU
2/1JB1FcOs4Ul3CdnPv+j+Qz2eWuq1Z0Nj10xCvcRMvj6q4gjMERnkI/puuaMuGo
pRCf7eCaSlfgRsiBrFHQ2mh5Jd5cNPcYRq7u8B78MBztlVLnop6WMkTJLMGItO20
sHNTkyI2+vj83EBOV+zr9YhTIrV5llTo/LTb8uxjeaQwM+7ZbVkoUm8T7dIMv1xo
pcBsgtxTwZcaGAuTJ5X1VRVXGqopdIdF83b6Q0rgzeB/51ppDahX8fI9sLroT3G0
BnXv4jRhWjxn9r3CYLXXzxevKqINbQ1msuGJM0ZGWpv3PUDSPLUHgqoXov4/8Pcx
pqRdKJk0wOKB1e/mEuEvzipIiNtDaZrAqK1kHmyvOXQU02FygaGPDxl86xrC90Oj
ZQFV0qG6+t13lM46Ul2YHC4r0TkAmfPYTKduPAU2VALzdO3Jqe4W4RHCqiwR1IX/
VD/FnnjxDbfW70mI1MzDXJY+LtcwcTOYxfDuf5Qqn8hv0rg4Ttbmc+5fhcbBw3SV
c8XLDHS+hStQiYXz61aa/C4U1QAnYgVT9YF+13aNtJLA2L2zZNP7YXv5ljLwZsQc
JM21ISJOHWqFVRK6+RlQJzvRA1B5OZZR6K2J9Y+38nQA93+7sslyh0TjEsB9ofj6
H4oMcldWtIrMCpmfC3Le7UttM1dE9a/i4msCyGnE0+H5pNH/wmusTpc/Z5NMM1u/
tJ5hotJ4ID6OUVYkhBhK6oXxawTEm51PKpcyEBUEHuOgHdnKJ1RjhYEEhTzAcNW9
KXZIzZnxC6LXewVAoOoL6FTR0S4PgxcYmaB5HY8zCXtAn5C9q+z6+SQH/fT+TXu4
6zXHDluBvloaD+v5CQRn5lOCpk7NCljmbpPGDyY+STVEAzsCOUTnAmL9SAe6xqb6
zv6MFd8WDTQcSKxGGEocb37W6jLpSXE0yaHhzwh25vRADXHXHZ5swa3GQpmPMplS
YQuE4XJLd9dT/0xhVYKxTp6rghT4vHx1c/RdXZckWAVsEhDp2X1yrc7DgXdp6pFl
/RLqGjyossOp93Hka/pLuUyjMcpcvnts0XJ1v3SpNYxvtIjApuonSssEvqQgd0Oz
d6YewdqZzLKE4vxDcKEkPCC0ioecRnfYizPVoYOeD9z+lZBHXjb49R0+t0pVUGmu
hm25o8koj14XA9GC7mqVhdPifsuQ/qVeIjmq4jNrBTN39K7+BQI9cj+S7yrcV2KY
NWcDRo96IDPjW3cwmjD5V4SLbqEb9uWwdFpTeEV14fZSvO5mXsz3a6gpYGRGo9fs
G71mEQVIGOHvGDR0ACzNNE92YTcPujSuYB55NobxqQmknSms2mRpfPBXeQUs5kk5
WHtATWx2jZpqzOEUwkLUXeALDKQL83ZiTZsw2J9JTzUMtd6qJtiecpU9ob6vMEck
BOeLS2+esGRuSFlqswr+zeTXOvDfT2QrCzZbqSxtNu/YQiM7YOdSzGJfIEk9x/p3
FcIr+cJSNNVnzQpEk+dD5L7GFx4n9a+6eKRP4SHSKvozJmXLQ50H5JKhkSEhlB3g
o7vvKwL7H/l5i74rfL1jK5YiVhX+ZEFgLcq2mSmXtxlVsFxnypgycOqW5Dt0UvnA
Uf3nTKj7/nmUed8X1AJ69emBATkbLMn7txKRD37JsQ225+pAzKF6Mab1zo1EmqaM
4H1byxNglYv/BfjIqhvkv4WIb39CFOCO0yeXoSPEGDwqX9m5lPvaq3oteHSJ8Tvo
0fsRiJoLo6BbTemYaqxKVVOsSFHYXMkWsMhrDSm7M1sCl0HVemwwQKm8p/srNm5/
WmVV3PxpdbxSbdUUz9U6/y8zYcUJDO6ElA6ElVkQy18leYAiDVCDI2vD3mSYOjvL
IQMswYT5afuvhycOXV7z4VTyzEg4wbNLEETBDhtmxwN8uJnXk+cpstn4hHy7bslO
M15fwuxNcZBWHubZNzuDOec9wID837kQIJQm0flqCFhh29ALBaPHdrodAD/24WMS
4LmHL0maMajhj8VB+JQulFTppD0CZws/agVXbCLDwcVkfbTrKYDnr/y5my7pfCGm
JL9CPJe9M/XQYisRR1HB/usncCqGVzhdPZ6I0umvIFL25N6mfdRJ7Q3JLXMXN/tu
IUjRF0w1jYEONmkkIlHaCcFW6WcGuMbHMfRM4GThs2rR301TI9D4vUGN/AZHiyxB
pePZMO0aERjCPTzrGw6WpWyBCWHEp7CvLFskJVaMJ14gKGqzNnH3aFRbahTg7tD0
qE2k0x1LPRskSnhVjp5JSKEeCp/wDYmgOaeBRIq9rceZCP7fAHQqLIzW5cxga+q8
IF5nXzQCGT7Z0uZErCAXDKhuTEKn1T0xeYPp0HLGsEBb8mMztYnbRf+SLGF8BgLQ
bm2/fMjh7fbelj+L2oqJ9+MUU1FCr+dB9oH5Hsw6+b8KjGcaVwsqk/7jYPe09/6l
wJBg+yGv8mGpH5okAY4NEzRNQ/Ss7coflnLxD7Yi4f+MpMP7Qi3Tyx5JT0r2BVri
tOnMGOplxgeK3CQbBl3QXnRx3oLPdK4atwAUifxEn8ZrsYjp8jG/a9Zv3GHKQwhF
YR+oxzEeavdyCjr0FHqlhcuaxfcMqAZVxBe+aaZUCHtdXZQzELMEWYSoP0HH1nIX
muhtr3DEvzJhLDfhXaACOf70bZy0m5WblsJVt1G/dnhyWiHNfdz5G4/XV+D3hEL2
pZG5AVh7qYmUQHOplWcr3D+4iqfK5U9YhW6TrQ6V1XlgkPXz7sI9c8mtTsyJQdre
m63874wNev49Uqfe0uFa7Ajxj2YxWdBW01BhUC3z3E/5qztS0eEQT12AA+4INUkt
W0NNCkJsD0EjEPdfK9cbN4KtoNj3pVXksZJdu1C5fiKdTcMunLu5z3EIzAs6628i
T3MWEZNfJTm6U0r85N3B3BN4qeEL82jQBfScCiit6J0jykobc1+emTTHKy6jCWN9
46CZu+bH4ZigGSNoS+zXnzhxzNWRssN5+/4X9k0jKT73vn4FeWiU9y9rOmaPBcFJ
vj+PyjgXahPGH2dzFQ2RY/DncxTtixLDtegLwxQdM+XXcCiX/v7bHLjnEH4lZU14
SKyCTvR9Zu1EjIFh7OQoAvlhmoxURLM16XWfGlCncdqrvq9cL8tRx+h9IbO1lR3b
wJV+mU1wd0KU+N3a0ga/W9U2ub5wyyVonMMn6MOO5yKD/FEVEmcyAeisG5S0MfoG
WfdqgOl3Bfnk1IoyXydKHD4sfmKm/wsKS7MDTrS2qI0MDXWcdGrIACyOb/Ab6+6h
bDWre8iU3B5XP+eztoffvC7BbODP8HdOGecIdrac1HZl1jxq2G109SWHVdt/YnWy
5j9tB/WgAUAtkE5sax4ZPObTQdAdVE9cXW7P4dYAFRCPAWNBqsBmxPsC1XBR4vAL
+eqMDXLS8cd+CH2D66MixxNWX+Wq+dEOmB0quQIMN42EkmNZNYJ0sIwKZ+qMVmFt
0SdD9LQxJSQ/TV/IuwisKaXp4AsEMj5SZqcVrWMnQuxD0bxmUO+CRsA6lpKh259i
YSlfB77TTPG7vJf2iwjhDhs9Ar7KDVD823UIdhlCtwOIZiHFLfvlS/Jaw+YmpPWi
wrQdASajxCcnDaw0YTx/xxij2SJdK8hxbFKwVFTlp0Qf+07HW+Xw4ZmrlwvmQnNk
0ZrWKKjAhIP0hspOlSwSHXSh+Z4Lbt0KPG0c3uEE61yjFqkRBzamK9GCdpve0iBq
3l0t9kLqyb0/i1AndI8ZpTX9yqs9A6VpsHC5qWnwgiJvBNIg+YCP5Rt86QQsq7V9
mSeAVinHvEKQ1AFOVxRblnO4fzGzJi7ukYYOi86rA+jz1MUUUZWSmnlZvM4zsSc4
m54zBM3+sdkUNtM2SIkP1NqOxDjemZwSeusmsR2HrkUS3qoBKPBEd4ctTAMCyaX8
G/WpKZ+sqr5HnZSZVtz50/NGUV1nHqTfS5jtdrPS5NHFZ/60NXkLV6w+bhA85kpk
DMeT+S3xVE2rCMqrwOTkqGupNzUTxs4RtVrHPKwh8xTg/Fh4nvZZ3WKm4TBBr/+w
FwlJpYFoUBpmjuq+JUPwZIBp2i9/iAZqmzTWJsgHoQjQ9/PoH3MX/J8Whk8TsJrM
3oij+TpFRFvAaJ8zBin3OIG+QtSC14vuU7gSlcrZ9dEdbv4uwahNyepCy1mj+Aok
1xqKLuRqRSGKGUd8Fii3HlhmKWBveoJ2L8uxNPbZ8X5RYoNzBZXn3ZLOoZcD+5tA
kIOCCGcPvpnw2xhGfH4MvKxFzYXMgDT/YrETnI/Hmd8CXTRo2OnWGrUjs+BT3X2v
j7Y/HKmYcQ38HhE2Yb/YaSA1MSvNi/ewYnqmdJxvY/o/AOxP5O8hbLl0T0JbcKJP
YWPbjy+N7+PRPZD8ELGo0hfhvC07NFwUzL7epqhE6boCNRqEhidF+DgTtaG06bnn
dvxVqIhawfRFQY2Wl9aOoDghja7wLVWetLBeTEn3v4GZK/hgM+5d0+j0q6zUbMoP
WQTggzRMlNmnGnITPv8rJPoSpesAReD1OSpED9/llQnzITSy3pLJmgKZWLqxGPG1
t9Zg93IvOjI9Vwdrn+PjtKXqVd0GN9eZNwtAm1bIrK5ZTJHxEmSfLfQLFNtbILpy
Tg+Q2qzpEX1W6aJkJ6PJy4NJvdPtcd1rHo1jP8nV7ri51lP8kUptBuIp+2mLP9RN
i1j7IZMSfticfvuEGKubpVlTQVcXLqJ2j0qAd/oLbHpTbtGB34GWd1w1RBAjs3JP
CUOkYCoRCa2ZJQLXL9etJLcJa9eU+UPyA2AuLkZ/T6mHyfAA16B6P+1T4EIlVG3k
k/TCX31BRHuOlz74ccdoyuao5XVY0dA+2CYFM7bLkYm1chcOXfBl5rJw+hAgTR6v
bdyKjj1jDlzz1NdEDqwF113Q9WjJ0XYLLweJIuYlg34j7Dll13UrioCIzLNXBwZe
SAGKLzyf8QHq81vCZceQH9B34F+xk3CyaxJR8WbFTpUI8nnTNT81P52VVQ9Qet/z
cwRhFxkQ/eGurIi8UJFBeDMcsjS4buh5cGhQIuvVQwBzb8s9ipGrQX1Vcw9oH52F
oMxdGOatCufpCzNTpZ5Z4+tEJu8Ra/Y03OHZDkEWV9FBlsCOyMQr40lecMXmRczR
FQzY9+SdLQhADUkowLKSSEoPdDNv3nhJ8OuGKfkFodUPUK6aEBuvr1gUd9YvAxp0
ARLrl0SZBB3C5qgWAJlP3NtXQ+lrhoYACH/8RSY9o4yOtOMVUYsN+53was+U1gzY
YlDlOzP0qG0bnQrxkMHZ3t67QpQ4QBQxS8dEsCZOhsRTzkl+E9hrWBfkjPseedFj
r5JxP10pFe4JPK7OpGpVAeKY/VXyVAft2PnqJ/eCBQ3p5cdoq22sS+FQ54tg2uLN
rgf5r1VnIx6mZY1tuGdQmFnn11OTHe66mUTMCvn2r086jnIFMWPKMXN3APsekMlk
8meZgv+3wJHUU55a3Z9nyawHyFQY9A0+Obli+uYhkQJE1SLeBXMPfe+kLvC7hv9G
Y2xQhOnaMHX1x8hTjNz2NhfS1XQDOlNTYNViYI/OR8RDEJY6xmAr9nIfTnfkAiJQ
i+nSjyEdEWpP2ZQf9R8yvKWAsMQS2OA9L9IXfeGOKrkiOvgaE9WtZ5Q4PfQgqSx0
5qBE3do+6PNVNOe6UPsNwQYOt+eWvcP0I0sj/R4/L0RH8j8Co541aDiTQ2qeXEmG
wwALU1l/vIhlHilWHLU3d2a3gSUHBMaJVRZWP/Iz2dWWm0VGoGt4VDjE1le8uQiO
nVFpwUaEY2oqFYzg4R1VIWo4HP8C8OAfbWLKhnNkT1HUzgX6ETlCnBUBMQTPrTHC
n1Q9bxa+B6LRZahmk6oD9kJfSB14TdpyZU9nLKboR8dKnuvTytKiHtipy3NzBwlU
BD7rMA4dqTV9n5IY9Ebu+CjRm8aB+PTTimSSq2FqnJCpMLE1UaS8XNpyZsqEcung
4c25e5aL8rgADPlMqVwnRk5oA+zY7Cnhx/92BE4cIBZb/4545xfrzuVsXsQSGklb
X3wHsmKryN+Cey2rLH+qzDuMTUYgt6GLLUxGPOWZTP4hW/5k8eLws5Ewn+xf/wyY
s1TQeI54kejKWQs46xbINfMFE/7MRRyFR7AGHs2p+AOrovMTCRr+yTztqh148WIc
FmwQKaFHz5s53OLLf8us456eiy/bKgztu+OJho7fBP3YF1mznpWlkpBex4arXwCA
nBxhTdMpCBex+B+DFGFBGGtbtVcnGB7kqbmCW7tfJoB2U2q1y0tK2IV+zfOx7YcI
rA8x2Q0zMqRzLOkx7a6ilsbVGxjjOxibNue2UNwKIFLgAjZdh57sBQ0XK0tDx5vw
dQV4TBp3ZjkcP7UIA0prdWuU3SEKZQhhvz5oDgH4gpQChXw3y+v+vGefYU3tZ6Uh
o5H9F2V38w9zfWJIcGHpcjP8QoU0pbEcjjqGOXFRK/XAxbbFYLhGL6UAdIKPPKpm
o8RdC31+J5XSKfiqLJRxfXxjiD/wyHIFEa9WlXd/pUIGVVPz1Nhm9UT0QItv47Me
kpzByPb7YBshKXNRMg23H95nhamZUCJ2bmgn4XwYR50=
`protect END_PROTECTED
