`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
0aLW/jphtwXMPpu6MntEV0BRJTVOaUqXhuzkuKqFEoG/teqECXC8t+Fgkacv9GY6
OIoPp/mYrvR4ngXwttLWjjfYyAcsIAmWHJLyWyOdlHXFAwtgdmL66t+r0am9cUEn
HtIRwIq7FCnfSB1L71zhLyj8xGUrjxUAfo1R/99VccepWJn20qPuzW1OTB+bULbl
WEMhv5Gp3yTavqin9aRNVT2Xkq0rDA7l07i4QhcaAlFJj57MSEXu5jNggPSx8NE1
n90SUqctlSqRYMs1PLbLEzrslL8qoFQ7Wush28X9hHgEL0Uv0Kx4NU3RBxRYzKvF
ZHVXfMgSs6I3o0wsh5W3P/LFsWxLbPu2OobBY0V4uJzEC/3v5o29dR9EK+jxfdQy
v0rH0+iuYo7IBfa7A130k6KdNsmKe4GMQ9uLIXbh+wyXM40LUalT5N417deQCRs0
N7MCVRPh+5xUsLxavS/zy9Rnec8yGzh1hPiydxPat/j3zzS1Vgh5yhwaRSx7hkFl
O0aQTA9NP15hn6v30qKan1SM8laP4JRnwxlO8oe1TkBcAHUVYDmmD6z3nZS0B/sA
1H9nAm7PVfl0QBpHHYmSxw==
`protect END_PROTECTED
