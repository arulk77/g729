`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLcQlijkXL3PFA9tTDy4Mo+mIV3bVYNrKNFdJmLYGHRA
gne2zVC8kIZpklDsw674K+7kdUEgjuK2nsorRGk4raCWkT1vaBJWu57Vbb32oNxo
dYwFMyODZAu9hc0W4O4C0qSJDwZCkvYWlaXz1jYbOIVnGscAac9q60H9BTYDwlFe
o6zjjlxzL4FmtfSkUZTrt8ZvWNTpei6aI4tRKhpXyYT4w/qGLsmOk/cxkn/srxQ3
gXboplfyfQjeRfDD3wdWt4xBXilJeHuOeiWO878Zoq0+lWh0ex56Us/GToFL3RO4
YMedI+uu9C2Vvkn5HSs4FjclKtOEJLDxA/jP2JZACALNgxqFElC0iEeKmBXfyAmN
fZKDKNHsTiJ6f0UCBWeaXo364r9eA4iGgBQidMLfyPxLXfurrmiPPzJlnDS5Nqay
KfZs3395YG/8iKwzkqXm74/0/4MFxzs+JDrA/5L0mcVqs6Uvi5yTmj++bfTQIZIE
OHbKqKwU8NPj66qUl3TNN1a4v58rUikofSHVn3KHd/r9J1FBBTs5NkT7CikQQvsZ
gQXq9jxlsAEeVxFW6Se8rzrHkQxbAj+RGB65jBt7vUtPdlGkSbF2xCZlM0SpqmD6
B7z4seLCSRPcpW5WFefltB9yvJHINFG6l5595kXpJp2txKsEtOUQ+XOrIr4MamXi
vJPYVs7/VwiKum83CPKV8ieKnTIVIpLnS5IYHLuS///y9GLc4dlculfrudJJfxXd
CA3/nkANX6x+qtcJLzAJjr5uGYHlJFrkaqyKUuGVT6kK7ZnVFostNcNtUmPdopHF
yW8cqJJGvYIRBSkZnDwPTPXUtjoef1c0Jvh4JyVYNKfVTjveRsEIGRDBzjMsZr2N
ifYl6e9QUNOsGdqmaCZbLN7fZWzsgTVZBcrWWDFgLnUGyGFvR8bRDoVSCGngTmRp
0vljcRJ2qA1rAIaQMt1zkKjUcPXqAAtOlJQtqYj0um6k05uBsbGmtTBI7sLD4O00
5pxIS5lMOCLQ93nReLPFjp7nYThQ5cIYmX7/7bcDApylI5qBxvegdZFuAQwDAg3n
cZom2RY9YnZCsjQyH4KAS4So/NH0wQSpczr1q+Dnzk8=
`protect END_PROTECTED
