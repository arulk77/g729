`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4w1KgcrgHqqUC+QJoicG80F9LvBLcqmSZ/zLOYHkhRTJ
MZ1H5en5KC0iuT6iK2wVCT0To/m4LqmM5Va6YAA0s5znE/15+r1Lp0x3GaJJl3Mr
E3Yn37bFfgdNXXgtESs/BOBxUQn+GT+vSlCmExjCKSrg0qkeOT9Nr4a1uP5Lhn3U
mefUuw8cwTzCl2CFuszjCCKAKDKwtXN310NZ+zRokGY3mPuZEu1c1wy7HojtM1PK
/E4QIwmWRFzJBGyQlKmYzdqYKjOkpBp3SmrL+NVrf6grW6ea7p2MbtCHpPtkjIj5
vmkuPHJD2y6ZMPCYHqxyBQ==
`protect END_PROTECTED
