`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN0PIjmxEGi4KINUv9GzZMdCeoW+MCMpRR4bk75CFRjB4
tQ7jG/CzKfflghwHAFJEqpl7Jp/gEs7zKZmJja/ALTUd1/6rzj5e34JtNNxn9ckX
pbCcsaMKOSBFqkPEi785cO1thvNvgC7I7GWsJyg8AGD2o+VNXkSMbFcysUTIwNay
N8ItULCE6FHUwt9YDdJdnxVMRYXCLOyFxIoTUxh1GIqgYxqMQ68jsZRhBEjxDgI1
TKKlj/B5J1jnxNgPWiARgdnSCbTlPMdRGvRLpkYaWC5sMc1MlP6imAU3rWxCo2wM
uX2SRNJYVqCbjFSEOLjEo7flD0yZJiqnYM0G6/tWBLcZLiqsXDEtVX+OqyIvTZ2G
r1Ma38wRZNtH5c7xS71Ck4Blfb2J67v1J4GZ9WKmaoqwZM9WAYEx1G9MUO6OxfmN
eI38DzYSgM3NDf10QXtr34B2qCPLgRFZt8dXg1lOZ2ZeqxTKaaAhZAyOzAzPkw+7
TWXHqTPyETjBq6fgNUtbZBbiftdTDqYOWswtNMb77WCkZLwRwBbY5Kz8HRmbqVG7
xne4bFlj8GqyNlVEyWn858b/Q8D0fmLR1WGwNv6SKV52gORGgVk2w55l4/o+s0pF
QzrXO7cG+2P4hmKq2uQPrgws6y+uRQiAwJsKYLyFfaOgCmn2DN4t2fGlEsMIGadK
j2BCJJQ7VsR2uwBG/hm10ps/lWPbQ1lg02GfkDahM3EV8rRN2GkBO6rPn5xtnKmb
J83Blbu4Qm9rzrYAJ4IZGXzrTL/yp1gNoQ4MoNT8pKNQzlSSk8YpHVBcmJt0hwaV
5Xb5SiKuo4tGAnlYErMljZF4WQsWy5WBkqZ3M0FfH9nB7WoiBDk9kxGfkkDZyseX
0HkxbJZ9DpMh01a7wZe3SE3rKEWOMEn8b/40Fm52BAlgQnNFo+F/Et3gcTkoix6h
YhLG0mULVU0IygRqjbFYsN99oDDM46TE525QD2B1c++XbhNM04PrWrmM1QINifTk
x1YKMW8yyImkWy9AnBeMyfTA25wmf92w0IEz90lEzJb4YApG/iZEgBXUz2PewYiq
nbR0lTL6ol/8AD8c6SZyKXmws7V3v8xntpMzceoLuuTD82nPh97oSv51clSibgbQ
RReRBj1WvG5Bai0i5rC//8G87219Xz3jeJqEu/J3NoVQ8gBS4lpmla+OAdlqNCGl
peNZ6Vr/esetwcXYt49be1A+eMnSmXpFGQSQjZsBeLV7Z733M4VN6QoFNxV6T9/6
MHZLsWZVLkwJFUKgKpY5pCiPZMnc8Q29H7RWkdcqR0b7aKn0UsksqxPBcykQUUGv
afRL0UjlQcMxrYDMM1CLtJDDihs/M60z2TKcRQMcrzribV7Xhf7NTGv9LGfyiaHF
OsLTOIcgzn8r3OB/otFbOHQ97a2AFxHJJ9XstUOmAwY7e8WChXh5ZKqdZvB89vGS
DzJkFUs8yhCPEvf5/NlOcgFwHIFBILDuiHj6BAoiHT4CBlrhy+btsiiezKH4aR9T
EESrDMWHFbhWN5tyvxL+xkUwA51GaAoGCLjePK6It/gZvt5lWCKAPrJq+UGAuJjp
P9txkrayS0w3wt9MZxmgSMEac6xuwERWhddWp0WEfKWui+EGyyblinbRLhJmuuob
47DFwDYC8wE6EVJ09jD0giVOcf7IuUAIV0i32NdeQRnC8JTquktPwQBxyaJ31oSu
Aal1WEf6YgYhEH6SFL7nt9XlzgMENmbX6qWtTYuEa7ik3au9xsJcPgjNHB3CE0A9
/bjWAwaCjFf/U9s1KtAb2C2G4R9DLqovp9EcQQjOopH48z7qMGKDKCP3Z3KkEODY
IiwjyTe3Xzv8eMj7hIqplKxwGNOV3V23GLZhJ7MDhzP8B6jX9v+mTu95JUuTtK43
LlxbdB+wzRMUI6Xxp1pPPju8T8JQbeL69s9I8MEEX828oKf6zHtZiLV2bJ8vCKcn
EefY6+e1tOSrwNa1eGN9N7m8lCeKedlFhhDnvRy0VuLqG14pqvREufmbPlUVkuS0
f0OHfKADp15g6uh90aAKGcIaSUnnhymZmy4h6O/A6oWFiIdwuFyDD7OgwEZa8t1Y
2+8H4kyRdoE7z6i3CljlQpXD4/K7l06bA/kVxxcw7tJ7w91xczzNWDs5VAgk4/jY
k+30SZGVWVOD6vnx6YbI9zIkXTE/+9n2Y42FuHcZ51onSKHJtUMKjtp6E5tBVSZR
2/p8r2SnZ7RuUDHdl/hyKCti5JBtR5h0C/e80wWFu0lgdiCthWzq3VDwfN5xsutR
`protect END_PROTECTED
