`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SXhvrlnf06YSxUO5TItOxRjeYOATatt1K5Qf4z5tslpA
L4AOb7WI56U3vtjq/97Rf2Nx2XwoFVSbvcKPo25jp8Y7+N1SsakxfAWvKs5Xo7Id
hgCQfqka8eTd+LsydyqtMld4en7eCZhezMfUTTnY5uNMJ7NhG29quPFrq2Ht+UQQ
`protect END_PROTECTED
