`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mlFBzCyNIVABC0bhYTMiK8lmmfQpY2aMbnwlWKiKsr7jQrgd5dp+uzRoLcwEzYSX
SLyioa4zfyG3sU4oLM3EpZMnbQCCGnEDNAS83zVkxhARx3sHlUpkAyFXBANy/YQ/
0RkU4mIvmh3Zh+pURlBlXRF7MCqMmeLhb4xyBO4X3p/6CnaQgDbzaKtzrmTYx8Fu
wIG3hAuvhJ0Op/uXFlVSTw==
`protect END_PROTECTED
