`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
n+Bw30caipeEjsnuwHpHRJND7P4UcOyKjMjUGvn4LGKgc2pgXpxyf4d96AMYHx1D
4oAtC8psbIqsW3EQSBmotvR+RYSbgY3n7YFO6LLDg8/m1SbKDElNAPNsPoH04ldb
RyJ/b8iS1NFNcdUy1Yj1I29XZdzPJpzTYiHs1yMD0+NGQiZFmm09DpXNAhEBPqCg
IFVfuza6wCYVOO3GzNvN10yjG+dHM0kmJwFriAMMoAYtIlz+B4THV3Qsn4xKzmNL
9+4U3iDeM/+vDDkZx7vyvpbWuiMLNZpJlmscupypd3w4sKiINpOw45+SD4vj6Otr
oNAZAc0rY8vkfEYe+HQ1PO4NsU2d58P6MQ7PSk+MMZ8jhBe+ZwejdaJPEgYt4JcG
6q67UDYtgQvuh3RYiWjGJSKO5YGQL2dO1wxC7eGYE1ChVv5SpvmLrX6YqZnqIItR
d3/owuf8ZAnNpmAzRddudS/Br0Y6M/5Zr5/98U79JezIxXs4q46C0c2yB0wx5r64
AJBA4xnYCAYtYqHeazQ1Lws+P/SRsgaKhd65RjpmUDa3WyFpO1Zf4N/thWIqh9Dn
hID4D4rBjPW3Gi3BW/rzXdIO94eigZswj5OCq+xq1HWh33JmvQK7jIgodKdaDmCy
`protect END_PROTECTED
