`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJcNGUbhvuXYt3sdZiL4PG8AUTnSgd8juGj36UEAM4TL
M8u2v55pAUMTnPPV+GMOanV65imO8FS4QFleO9FTYdzoISrrUq54nWYol2K4vPC3
2ApjYm42aJl+TBaT1wyJ1gBoRz/XvgYH5t4GIIB7HeqT8+xe8ovpHumjw7GCUMq9
7fysFg+kkHAbDr3F2EXq7HtyqSWwbaLuUAu5L5tT4USqwdArkMkSjQty0ZgjrCMG
prlR/AgVpd26JVcYcNGqWA==
`protect END_PROTECTED
