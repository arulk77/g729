`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
piQvLyyAErZ8hxmhUW+2bX11UrAh3/17olYhLPx0WyJf3mDDFJfhrx74ME2515FL
qoGYodd2/ZOvhbjV4X0dmHadcLTCi+F5B4uDNInJlAsusUciGslSfGTe6GNzZqV9
+xeSiiksDIUF5h1m7cG9ZqXy0SDJ+7eS4u5Eyh3GbC07Hzgumd9sBo/cQXIWCgxM
npCtYCsxfRII7m1tsXb7diSbjdotvwGY0YpREMEtNhD6LXA8cdy4GGw6+RyEKp/i
DNrvU8GxaMRbA6Nmvrg5XwPtgUe6nymIn6JoYI1iI7RnV1Yuus/aWByhzSRiAJqj
WsXzPyTrSZQBhv0pxAaXu2YxWH3fhS/HcWBiSq5F3oabFKdxt6p4QA//txJcHdRA
eTmMZEi/ppukR7U1HBcHBR19otZ8aa59eR9snuwUg83bNGtKB3Pjn14o0zKhau+k
rTZlooet8DK29YWHkEFPVeG1m/wKIyKfW6PHVnjbo3+E74RH5YeQqJOjAUGMNM1M
QYYhkR3dHTcJzGnzwIzEIFE7Uv0MzZg1loHPHig4qWKEUFaKWlq+nF8pGORt5PQs
34KSGfABhs7roFbK4knhjk2Ti3bOLX5bdD7zb9uiVImJzP/mntTMZBJik6hEM6LI
2I04udda/oiW8n2KJV2oTCv1idEl9nbeuo5lrw1fLjYphETQrUGc0WtKFm6dB9xC
/4ZaIK73wsXp+DwkSlLDuM1G9HHU96Ev3DO0VSPIxkL3Vdts4+Jyjbirsk70L89q
Ry7VwL/iq53uJDWkjDB5YqMeY4N+e9bqjvjqIkD2R/hQwWXx1Jt6pbv9uvzIQek+
zVfWapB/Ezsxi9FDktyOEWbEsXkX+oekQ2G7L9agZ/Bb6bKu/YTOlzoDSo0lLA/z
4OFDBSKhhiT3mpRhW5a3skstYR7d8xqnJOvvpqQf9tYuzTnKcgHfqcVceVv1G/J8
2PILXUzTcSSKTsY9Vfid2nf37en+eumMB2qC6mulvRpqzNJe4l+dzWdMAR/FzuD+
MD8ZVfpt5G7+pLrbIO3o/IfcVJU8M3dqs7CUEdX/Tc7tKfeDDTCIdhQdNV9iq1ON
f8tYLDKpLss5/sKr63mHbTrUxhEmxCXNz6hw4K/8mZz8yqFEiJRQzxfmxNY0MXgZ
CzZIRAGPaLDjcFvdKA1mW5MSg71T/Pm4iuQRzgw/vRtiPVNzh8ArepfNN/Uf4Gq2
H/Ia6biqf1v6q9FTIGwTsDwqUmJYKYUsjvb6A3mr60rK33a0eHjbG2NtqKE/tCp8
y6sb1Y/eqaABWBKSwbhm+gfPNn4zS8eUGH37WPloEL7O2KipjgPdCVaM716KqMxk
7lznkiyTJwwHUPVvPVuvF13/GWmelFeuukY0leuQWO9m5Awoso3lLjX2Ej+WjIuM
si0kY7tcydcG0cJ2cmC7rdbHVhuz88VMYkJ86JJXMO0MV1GJBzRqJeKPVzG5HVVJ
VbhCnJ1lAQxEqpZmlHNc00klTF837fyhD8XchqQhwaQdAtUQcmBSFneuOS69h16p
wBnnFVMhIJ2nmCvXXsiHP79H3/FqNEDPyjpEWzJajgcoQ0hxFnbcI5cqUwFxUMIk
txB3UBFwsYgK+VTgEe3C34QqDhUTzCMjNx5LJdffrXHPdNS9+BfrbF7HvFuUtEym
3CNIzMilhaGJOlRXuVxJR3J8WAK/Z1z+ioxkuYUrGT3UiUXyCO8Rz80UpV87iWyX
aC+Kfv2TvxeeMuqTjGQ/ZSWQ1ox5xYdpCXg1JGC8fWJY63Nsx2kNpe6jCkSd47+g
eansYz/2VfIPlLeTQnHC64+BkR5lOlNWGog4LcxJms0lBKrKz0pYZBvgoJPwb2Pm
Iz18A2oGIicL0/onCbbVVjASMu0zKlzXeQf0Cqq0IFoUfihSQNXsA5ZGPARwJ5ey
MfnVK4A1hLLVu4f0JsyeMkgB3kHyE6gSQT5cjpbeewPUqwtn+Z+rB9tdgOtlgavC
4qwjSmt9dGlRTOj9eYDKhhXLHRa7fSEDMP1DaYrH9aIulhy5l3C130BSndZf2aUQ
btqOvLX2f5Bcr5utWrvI42KADok+Rty2j+zPacjFplPJcpNISrV6HydSwStmv0/N
sVQQKWTDv96YeAEJPVnmC6QqGIc+PslI098We1UI2yB1x/o79OSZpmpmLSBZ7CU8
3ukxvaiFHYWYwdutY+WxMZoC2lDCAaepgbwYSjc13b84Fxlk+kcgVn2RZAUduXDZ
YnJPteRK8k0txlVBqKjyWIyiXyans9fsUoopCF5X5Xox5qDhu9Royf/Nh16YrJjn
0Jt4YFwoVtgXdd0gY/UybEmNL6QHw3VYB9aN0x0Er1pNJSc4WtOECJAmQkTwf6yF
ix3iNTqYDbRCTcplYSIaOw==
`protect END_PROTECTED
