`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePEU4lu4hK/1jkqCyPDfGTpYWgQaootiEuf83l2f10zW
Ntio6PHXxJXGFQ0OEmIx07e5XUdFzeC0QEIZIT+fkPLU3eOv/FNXbEuemX1kkwT4
qIDAp9rzU/f7z9+JyiwdGR2Cx77Y291WOa46mzFkrqwHRqiqvoOtnssA3hZs7jF4
`protect END_PROTECTED
