`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yUZbGY/fUeiz0HeOnUz3p3GO4q0JuanyBpyiBunpzWL
UY381QFP25xoAY6pZojJCDKcGzCWT5rzZbnzb1FWpM7fonKRN5Qib3SqiYlD3meA
mCC60G4kh4mjxwPi0yf6H+Hki9aH+t+XGxdnNF5isezX84CY/6E+fvRC5247U4AP
7Nc4f3/RIcczO8x6u0qtlL0TK05xB7mBLBwanHE6i8cIDJPHbJDrsIp2vwV8ySXz
wXfCqcOUDHGX4WqgRs2kZVf+RxrvMPePewmYis69ycV6258E2/SviylX3kUEVOw0
+gscjWV9HKp/dFXoSxSQhRmWVCAGleQQu+J4EPrWJ8cWgBF2DJlEP3/QXK47u0EG
9Im4odzoW4XjysQPQEGTcTaCFgr/BmGjyZzoCkiJStCgqeyUZZKTuSLXSuOHhS/n
JIJGTYMM2YfPf/rAv32hyw==
`protect END_PROTECTED
