`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAV9ujZWgS47k6k4OgB8U5KcagX0FafW4XMz6mNk7WX+D
PTaDmiiISsEp3kKcW1rIvaq1/RkfVeOh3vdwA7OVKfas0bazWUaAnJsfXFTngHQL
Eb6GN2mP6pk3li8FxHasCTAnrUb/LctthNpqko02csNdh5ra/oVM6r0cV3kAzUAj
+YsAnyTJw8FCyGrzBI47PAmxgvTGqhBGPPdZKT55OD0hzEhsLgWCk/XCg+gSWcDh
KDDlBy3xUk2NGRjv/3FUiW5ZiDNmcyVs8/KzL1oifPOcBD/7MaJID1MlzGJivfTV
EWGLGhaU5CUV+/KHcMuxf2Vg1H9ccDbVlPxajcvHQYHrI8i/LvADhGX9AbXVKPCH
VfyGBduRotXkfVa9ZKmWyYFBTI+ZetSfK7VS1Wtcbq4bMPLUPh9nPQQh5wYjxTiW
U5cczcVLqu+QjxW7xa2jbzDXD0+CNRSfOX5fACa42jIN2qVbf9JtRDx8BeTn0iG9
4vtxUeRRkAJC133xa/nDz0N/Ujs1+dB85g5zzSZkO9cjuMct2OICCgJF72FX2KmT
yUrHY+hwEmDkifWGGTdJqcBDPPvWefZg6FJZiqA4oeAH0dEDRZiNPZCibRLY+/Jg
azgE7LXDilrpWF7IR8VqQ8rMj3o9jjx0g9OVcEnPMARjPsnkQncZYHCQZVR17mOY
zcvMBxBS2JWtRMlWqksy3Wx5Hof6pxtFuwghCHWKJNg=
`protect END_PROTECTED
