`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
obhtXt4WR52I7DxxjGC9EP8PzGWJebm+90l/RUf5AD20KGyBxVYhF0w71u3bAYO9
mdxcdHTyShe7c0ZNRJe2kwphdxggdSDN77azhEyjBq3bgvn8dK+o2p1AFmhGwho7
FFObJC9UtoPh/KTo6MTShkD8tqiPV1XFAivDHalTfgE/CjfFkzjLWKaUtU2QGAM6
aFeXgf4FLRuFmaYz2W4GaO1mdeeAP47AX22Lx3/qbX0K13pp0zJcPbQl1wSOknUW
aUZZRlMWzBk3PzyA7bbxQvSg3Fm6NTT5QBfP3wNA+yCgPlZeuNiNE7+qxW0GKE15
rm9BSyxdVHk0WiI1JdNntTm1kaauLEateBFxzk6Ul8YT9oC/OgTslYxUwX1INRwl
pUcEaabGAYlDduCY2j75ElUa4FnN+v9kQdYT35fS/25/yi9Y14QxwTGakKjbafP3
P3JsOMlsuM9zNNhCn70pGt0iohn6eiVAOzrxEHvg+98c0D80l7FiHHcppvUS6fwG
/eCKx2T9UCSMPTSvJKb0NJCFS01DMn/Bqrg7kvFE1iWTr7sky+8MhldDxXvUvXRN
vw4QioPe2zCqOTMBnYnKERlPHH0cBQArH2ziB3EuFesSuMaPRHLZawxgO9giLlk/
/u/AwxBbk4KYOo1tf8StRQs7+ngrCvUcJ/a3XC9u6UYyHoEodw8cSIOBEGMrXRy9
oyzKaX4tHeEjkcj855QxzM94mL3PC66MGNLQv4wxDWA4Q8ghWgV//GaybP89v8Jl
PX98JioGxioC6d0NT/VeSHW/41Jtv7nFTArx231tZbiFf+obnOA4vgkLsK6yQgwp
ejH8a8VTstwFzYhOiO9+Nx4XUz1uFLhqPrAbv3jRV9rWLKtXYyuCBgvyeVma70p4
GW8uYXINKi7eIh1EJalAxeYtIdKJVOJxAJ25cvd3okPeQWnDEVRCPAzueKN4pwUq
lbVAocrHUCSs6FUXN6Q8pqyRK68PVlfrJdr4mbfhvb8JHi0aX1iZuAFXjMciWp5m
DtvCnMN5NPbZwNGMFrXVgftmVf9Dr6Q97h7jc/FMj2v5mi2NK8UTeLr8Ts7F2j2X
yQEyEMefswMF2TsICcfpJoaQbOh2pQG4c+wx4gyV4sX56ojt21aX+2Ql5oiLryO/
H0cOqKqxx4xjObuVq8l6l1D78a6xFtO5QWEVRNsZiU/IYNjzBEfpvwOQd+if9do8
9MNCHqJvQ1r1MHKjqaRQOZsQD4ybdOAR3Y3YDPyFCiSeYJEhWzEyn4NsLMHR9CfW
s9iw1aRsRSCbn0rpD2Jz9UxMmX4Y7an9HelpxK+56w/sqRa7dtNB+MjHqHmTSmC+
nbYtTNc1IFNWbWnLDCMnZ/GfDsFB5xszDcMNfnNg3uaDdX9KCG4TtcivQLMTjWmX
FbkV7UtCrNgv5PovxO/c+0cVIRjfYmuppsdZ7Amnmjiqmo7Nfvr9t+8EHsdP/eqW
30oHbmhCT08srmtPpby0ZXJns9K9KamOuX5ox4M1WXR/aKEgsXUCZP695h77gqme
2mkaSQs9vrjaOgsP768RN0k2aabkW/6zLNC/Dhay9R2LNritdnQHQdHOcYe6Xqm9
mL5Ql6DY5QABLGSioslwqnjFlMl+hZGPESiE1AbGEZ8jM9GbR+8GsUJSsAypkAGD
QI0I3AhK4Gv4r/DIx4Wz5/ZKa2Hbxc3v6MX2mCBUWEmwsFEGsg8eMKy9C8VYcPYN
3gHdX26qRCtVyl9NSZ7RbVsfOYOPWrovSMUVGrbbUuoEupymQsnBym+W4VqVa1RG
lAVNh865kXoQCvSg2SWxpRG9o2po6Mks6/yIa6nKDT4mP1sPN4r/DPcSJYrQ9SC4
LzIhw+vMS60MUw5qZj+1VZMED48I3AdsX79pSVND/XLrPoi4pDLHI0EI1OPvhKlW
wOTDv84Nb+PkQNZpEJ5csJb9sFB21A0S7eFFfK2/+EJVFoLSHlCXdupaHbulBYHx
6L/DzNByrV3m7k5Ujk2oZ6jtfIHv1B7aubcKY8OVY+L5sRmDEMD0SQ0spraGH79S
V3SL77psDHu26ItjK84GNHUdIj4bIKe9iPipMhaRysWRQqNwfCztJZsER9bkc/9X
vLx2hfvgqE7rmuakngqjG0RcWA8HzFI1LorxLedjTkaxWpkZLvgQBDJRhKwFKWC/
vAwCKQyyN5fS9jVwiJ+1SET2kjPcoyZiB01HDANQNMUx2PSLNo+dFH9Z8GUscIWh
IfLy0MWatHWXnRExydoMRYHY569fhj0vE7ISYcBme7RMpCC9gx1sWPvvUAAlQXQT
ve5yqWZUtbtcBQMkchIaHaSinwFbqhiZY+7CnLeJjzzGN00qarS81vRORkzLqQ98
lgjVIl3zJSQpZD2K5BHt58oi0M5lUlrxpaQGUUoNvPYTmhILNut/NKuCT4yMPA1u
6xZEU3jgMje4lzemA4CRW+7aatruazUxV9TDjPVzqzOaxpaJUqg1ZznecBVYoPKq
8+OIjFRgckrWeBmu8FMgOXvwiOoY6lKHcjroEclM0kM42hmYnIvB4spen5j4hWFi
WKrGspQQnSJ6OhOJh9eMtQ==
`protect END_PROTECTED
