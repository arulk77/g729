`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ca4tm977cT3oSMCiIrgms3kFl/0IiesNw5n2oerSMu7CnCO8/bN2M+5UsgMnZo38
oTqFd9LlKPcWyp8gp9Y7+kex3BBRjGHerbNYKcqjwpT55vxOPozurWsoQ99gQNj2
ALZgXIVxmzkljkm6cyWIT0lBHZzPqm2yri9nBxz/padp1OdBWUGEvTKWwVl8yf1p
u9GrpnvM/gGnwJY3jF+EmPnT9qv2VaWIC71HCYaM8DVTyH+yaeBg9Ag46VAbMYLM
glYIfyD/sLy97N3F/rQEVVJ3NhJKEOLNha3W03d1mb+zUts21uKXmbZUObsddzFB
TrBeQ4/9c0C9eKdrDzrPkXHjWAdd8/lKp2TRN8BPtJL3hk5infhfuVbfflmm2FIU
XmPbhqvyZZkL+CAmLrUpqFid9CNeNtj05dZT5gy2ooVeeg1sJU7SzBs7MVwByKWu
jtLGLl6rda3A4f7kDZn+WXiw5c1q9iBAMkz3k2y+j931pYK1HSeCB3cNQebmdgOJ
8AFdQ5JE48oNSU8oYRYOL7YMXm9yQqJdkCRx9UkJDsdNw50oDtlPQ2VoEaWpD39w
Ez1Lim9gyXyM6bz8slubEVsdXiD34V+2HxPZ9JH7ZUaweIsbcyPIdXQxE4nb+J5b
Lt1Om2lWwuCvqaE6ik0odU/hKlBMOKis0/m9pR18VAKR7HLfWVdxGZw1ngSxP1aP
WvXFWS2Lb4H6CO1taI7Uwy6JhE2YzLz9yCrrP/IDlU6hzBdv5jkgMbQ/YpVScrtz
S3omKcmOQzyi6zqOM2Eb5b8WqCAbvKs3DuYkVRUsEzIP22RSI44qLcqnI7eIB2S+
v8FNUvg3OWWOvggzeDs844SlOj2JUno0bGtdirsU+3VeFwcafq5a2xKFCM8u33rQ
7tKxOpKxizj1o+f3O5mRB8rHOpAZEDmc4Zdd6mhmV8Iwda71+EqCPcAY0CrhEaxj
Xn4Imyu8pSnH89zxAEK9Aw==
`protect END_PROTECTED
