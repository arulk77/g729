`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJopsx2DfMwh6gg7bbWtSDXqUIgsB5HJOOux3NzOXMbf
OZYAyFz96yH6Wx/QUgfPlh+9mQ3mRuZ2SpZHYXWPM4nxQR4tt2n1gaf3Fijzduvg
HvCBrZo6oRrZxEOhrhMtFEg5i2b7Pl5O1tg9ezBv6ox2cxtXBHLdaEWlx+i17jjA
HlkAo+JZVJd5zEa240dshjQukzPXquVrIx59VVyMrIxTNy2fEFmUrpeY7z3tY9BW
8G0DjP80jTGmHc+oNP/I+ZaOP/6YTBI0jdFB+NDmMCxEnVV81IV74HbGsNqij25J
w9R+J9GjynSKNBvnROXSNbl1yxPPtLv42bEPJ6bikN3j3hjFfCk+RoLjG3YQgRxN
N3/sew2/FDHYa3KgN/kyMnAt2JkAXY2E7b4pQotiAwtNl2Wmqwy7NcITpORoycZY
fs3VGEgfNeJPkekTbuUWVkNNA2u8ZrLgJB+NgR+9wQJ7xWTEP1RdMF3gmCNw5PK6
D3i/wfnQyEWCVLUhu5vgTcX9yeSqyeSv4w8fkKLh+eGp0q25L2i6m3GlWzGqxBTo
eK3CFA46XNTn465R1p4gzQ==
`protect END_PROTECTED
