`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48R18Jn3n8hVhnOLPfVWtoUqqUYftDUvCffTXlpfy2Ok
ObpRkeKnJtxrqQ9pYSLrnowmIXutaK8qkd9975+VsMKma0Yn8bHcfBr+e1WNPUuK
Q+zpAapqlF/i5enw8JQuy9hMANJfnpFItJMOQGeS0Q/RN+RQN7vKd2x+WAj8UCyZ
x8prxO0SeGvc2hSC5FWOckfWJAPPHIFabz2pNDEziQlg+Fh1Z3Hk8weNniyH+ODM
kznelC5injzV6MjjbStmvBCuXblRV9b7UiOqzSiqCgO8imO8XoFD3mbuLHzU3s2A
i9ZUPx9aagrDa6BndAT1ng==
`protect END_PROTECTED
