`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN/C3khs9B1Uht5ec/sqb0/B0ihebvx9kUccAPAOG/a0
P0y/RWRocziOzZARM2tCfmwKTFQN6WdyS9gjyjzdSV6Jj1eYFgKa28hrP30nDm5O
DB7ECr8aqHy1Xn0lAk/5MOgO1qOgsBQ+fePXdUu5Qk2L9eggXpkyY1NWhCF78wfU
ObUCvnWkJ9LakkGH47FTnLsY8EixKh6TH/4FnxkJYEQYMqDOX+ODaCI2TXkibkPj
dc1OPs6JMh+6naOXZIkCucUkaCgFS75k/UlZslgGEitIOPzoS7IJnSO1Usf27Mbw
j3LbAwxeMEmIOKHt5Gzke6/HBah5k2SfLALnwVqXYTNWt8UvwxMXP8RFCRiQ7ErX
bH67A4QSnTwgcaSr0oYaodCRKOsQ+RO35DZjkoguCXeWhz8kXWmpBWewBJa4FMAt
1T0lKCsSlfoYgOxgNLR6dmMs2oUfe9m3gS0skQm6H+vheV2WifSjDMwJwZdzLvu+
zdRMl17DQ9lAodaEwcv/a5BdgXTm4mBB1ajYfqnCc2kUDoRHlxHWnD3LmLi04+O8
8PEUD0fMXFztuL6INfEVNGnbYRNnYyxwsyJJlQCjSbi4rjF/n1aXjUtIY8s1lTvr
19iXHAWrDR1EJdyvvyph8Kzsg9HLC1BB2RPsYmu4Vv/YcqHPHksuekEZJbP5T4Qw
jsIWOptVIh4PSC6OYMPShouiUKswvDC+yV7i1WTLECBONYmoXgOqp2+njkCeXKL1
s/lNXd1SIYcOthidn+MIMqLYBGjpHofDaJLIQ8oSSYrENKS+pQF9IKl9gpl5whNP
ZDfi4gOILek1QazZX93fd3iHS8U0RF1nwPvJhxhtbxY=
`protect END_PROTECTED
