`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44Pmdc69L7USKbZT9qwi6Cs0b+aB5wFQojh/C8qog3WT
2Duh4wOjqdOurBOP5XwwNsK624V9cEJWsX1axFDTfLrG0ffzOsB6e+VvLVwRUyZL
pqMFdvox4RPmt6nEa/nSncARoD4XTqPwdoQGzXhCuKurOlLt7VKPZMyX45TSXlbE
GEyF8ogVyK4ESq0W5pSYRPYfGmWiZHduPeWOfAiJ1DNrV2UXwweuhFTAA19OnU8v
tWzJOl5KLGiCG2W6i397f8EifoWzyZwvPXzimjhtGZ4eHpIyI5nCFf+pgw0CiQQv
YJt9oXIofHw7MjoQOysfGJ3pmUdFMisZNi4YPcxTYtXSmcz5AKYdoxq1YwtXWsXI
i4DLW9cDJNYN13lhFOdTCg==
`protect END_PROTECTED
