`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Na4wYWfETWm5hYPPBogd/pgMXclrr5lhpPmSDiwMErMYS/a295cq1cmMgB+HG4U8
1hZ+hQtNucm28JtnKpy86On+q15yUl5fusjekEeV1kj5lwHnuoHqfEHulj5/Qkx4
T6KQ9EOAqD52CZcc1ev6Tcc0V4E1MzVL1MldEjZ+y2KH76JL0Qkb3VIqXDMon67Y
AMCP5dZbjZ/mjQRpcPak2rvw73VImejHTr0ZQ6XMHCLMcZjv+f93M9Nwv28Yb99u
IEoMTEIyr/PEb4MU+l/9SuQrISx1wb2o+7/jIi2iGb4cB0lL0C6z9wPHq8YgBqF2
ATOtVx2yDb9WC6HxXIU+JNiLaZhLh5H1qNmCuBqjwDaz77xvDHr/o4FEae8USnHU
`protect END_PROTECTED
