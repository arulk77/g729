`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
W52by5FksJUdhgHLv4Ym9EKjlA92z7B327MLSGlHSsEMN29eRNUxXKTLR5chC9Cc
ndTQFL66DbJeCFA84V8uISLIHvOoR3vOs7gAh0IBcFX/p+Ir6BRvr6kVB/mLl+2G
oduNT2/gpZE0NNJ79tH344O/OTlRODXkAhMK9FMPP+0s3TS3A2SCV8xUN/4ahTXs
Z/CPSIokui7f/DnpCMRsYBiaE/OV2+Z2NjZijesrukYgefgnjMPw/Eb3K9i3tBzr
JiEP2swy5M9iR96HkOaCXi3kZ8fhhu7DX0Bq5NUE5uQ2aO+ULMKYf/tHOgTSXKi8
oSHT4WrpTs/AhU3+EwlvC+vmgxOvHUUO5oVKc/VcwTZjgkDQtPkBvH4VPYIIsN6Y
BpaoLH0DC1Jxw19Jj7t/Do38bcnvks7E0Qt6Oo8r23I=
`protect END_PROTECTED
