`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
CVPz7U0o9IqJbDibbdLvIYx1zx/wtn//ZgKjPaeZ1z/zQrHeps3Fa9CZYNfLaa91
fkyAidCig9zfeViJ7JiGLzTbBb42CT9k6+Qv5qkai8c8CprtPV3a2h7SzHktBeuw
+MaOaZflIPptnWnDdBdLebyIXQVJ/zrspyVVO8dBqYI3MsbUlmD4VfSIXQto0QLo
6rCvY0atPpwYRVTu+te9PK9wJz0HHZjlYTv9OI9cs0PT3ihs/UfvQ5AhQmC58OKe
ZnOlIlvNK4oeYDedDkoIvAHW94mAI2EdDoqgDkXovgxc3w3maFeC32N+LaLuF1uv
v6HpcSNFBIXtc4+eadXDKm6kXuMApafymd92d/I9CP4RwHLn6WQzhPMDT+Dp2CBX
MonqASto2+3yfNv02g+XHXjZm3u6RHyfsMJpD5IwDY2UkCZqm/2mNOSvBUhVy9Gn
auHw1G88wjHxdnZCT+WyQijBaNKDV0NVm7j9+0BqjlBktnDloKvMbx+moy5jm3gK
2yjxneYpWuW03J8bQuzDtCCIGCiNAXp0YkOy2G8Shje+FiIkXbo82rd2VBeEfhYn
/tDCheROsmtxaV/+8gRflShlDdcdMdWEMj2oGNLqeuEZwxtgbPAOpjDKdRWRP3xi
fndN4l0dcmihJyGTTBm/one3C9d9gcODksQMPl9UVdJGw1ju6GaRtg590yq4u8Dz
LZ5r7055/QCv6OSm++bfuUVpK1wT3qQllEc7Ho+MZqkEpZ0Z5Tg/OV2VtEpyeDxH
Q2cpJIsqqZVonQ420MKr6NLS+7BlmIfNPkAVth/b1EAZgdYN/DeduB5LNApJgXQr
mTVR1irofV2+Ok2gx61x8AVvPe0+rqXuWcdjwGqg5Aoi6mgZ8/Tz2bc1pxj8baN1
ZVKX4bM9+LYJasOtZBl3QPxcg+QTT3kcEUPQDCz/I4XqfduF0mxqAQLS+DN5XeNW
nD9PGsVYYe5qUPnTan1ln9eTTwU/6STIrjc/6htDWdsDOiI59iNN7XlCf+tPL9Vw
8ikWd4waXs1129tpZfVeLSvdY92IggpUpVHj7ZfY5/Za0P82BcV8rxf2wMxbJ5l4
duIK6XW7+jAn0A0EA0OJVwyslj5c83gpDw69Yr1GJcgztb6q4Tu7ZXN8mJXV5lQX
kC7jG6S5gZydtIRZkwSel1TPARkOvioMvZaHdhK9FVHPGaatPak+xo/8MDb2hSRO
BCdGigQAgWig3tM0r0LkuFL9SZmXx6a3bF9576mbLme78DLmSn3NGKAlb4tB9dvO
Lpq4GhPpaRDsS7EiwFm1AjW8rYQwgHfIekWIoEjenn5PDEVfeNMqiqY7fMiwpN+1
GSlj72k3Katu+/AO8OYlkdSd2Z1j+QwkEez+0ftMYM6Zt7Re5hiqYGHvBSb1I1ln
eWzkxnX93427YNlZM2AwBP+BzRW7vNwSW0nSFiHGS0VQZwmj1soy9ev2GOaX9d7g
UifsdgAgc6HIakh5P3aOZZ5+rbCXXvHc3ChHvcOKugeniOXrUqin4QtSKdqGckIC
VdGhpRrNV6JI0j90/rtde8psd3J+fcxqHE0i/I+WQ/ABuGaJl4Bb5ZWG+PYIR+wx
`protect END_PROTECTED
