`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44jbn8d4UeZGxrdUo8D/LbJRSW9Vv2O6DJlsdGEnbRg3
eLRl3P34QG590tEbAws04qDRG/E4fZeMeptmlhvYJl3rMhkOg9c6hma47Vb025uc
SHqJ+78DA4UgEgBwBJMRQ9rPBapT2vGqnkbbvr6XynDFPzFVj4kr8ZmM1pg2PQl/
MUpPMTaDcKgES+SQyADhYAY33CV7Ox4s0i5OLq5VfhuBrdX06MgKcOwMc9bLHWWl
zavghNeAc3W/lwa+WcLmtromb29DfQk3G48FHbLai58=
`protect END_PROTECTED
