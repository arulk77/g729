`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN8A5kvWl1tLpoJ6TviyBtAPVYdTAzRfCChzZwMvd4/Tq
nKvwIFS7yLXDgzAZDZvmno6BFk2I8LtJ/M6Vsd5SwwdUrYNvErA4R0TaSx8UHZrW
tRWzqvXndWUS2CvVQ2f47QnEJX/HS669Q6cgP4ItGvtqFMF3X+FGUKFb3JabP9JS
gl0FE7A7WnsEeKbiEUiqYHQ5BBHfD5wStc1zHo1hhLUyL3BKeOv1+J8d6RKCFNld
LJwGvFnTsEjlDEqn6J7sT2Mlk9nagq+wYoTdRLBk8OYa7juyrAEvGaQSwR7bGEEU
w2wSXtX3gGuPxdCDTd7cU0Ff57PZdXBQ5K74Enrs4WcdqwCZT5iG94Fo+0BgswVT
4lRiOU1MRmMypC10EwEOV08sdw9untf90tH7NfJy3nR8ZJzXnhnHcfEbJuZUMLjE
iord7kwTbDI8nXBXxnzDaDgsyCNAr+ACeXsB/+Tut3tXpGg11j4wsaL0Q/7KVu1E
7QvlJr7J1RayvEcuszhd8rAejqIvtdZi8+xBvbMRu6VAL4J/vM5ZycbO+hnwZGYQ
JRLWq6fMtfw2pwB82fZz4cRM8RKbqo2j7XJRMwPLuO/9uutWwW+IM/CsaewEKOKT
laNjbtmbGaU8676OhNCS3tTwB/ZUBWy7WuXwQlrto5JlSB+FGRKivaLCD538mUYS
acdRbjwDLsQaN823+PK5j6ix4DSJIkBO+DVDaz/k69+OP314f8gpdUsJfjgFExjt
HFyi+6kwWA69OGpABGU1H2tFRuqePGRs8tmTs74WoWnHTVQis2BQ02twgaB4jnA1
EFHY+TpW/lOm52U4r30fcsmQ4JPuJDzU3+FtI2PY18JAhJwR0nOHU4jKGBXzopJj
pPTLdXC2NnaHt/H4QKwuv9kvVZn48QWWqtcqp4CEIqOekJ+noPTdks2eZnVpJ3d7
Ag6uXW1nysKPV9j5svDBSY243ZRik4nKJ5NUpSgao4J29NBilnBPixs3qva2zvNw
8RtaiJkLJL/S7k8e4vXSU5tJIMPgWqb0tNGJmWwRqEqSY+mBgXDxmTTbSkomgsj+
ZnCc5KXEs9/EHd89LgT6HARH2SPNIJKYuZi70ouJpnQO7xnziVOkMJo1Ou9DFUIo
qQVpyPwDAE9rGBEJgSTIG7s8KlfitwHyRLVSUGdIU+aaN/CrXXPhUM2BImJd7r0z
ANkyjChQS4uqcr/pV2tzQurlP/3qs1NkUHJ5l7Q/2NBPRRSB+cW5N+CoQjHYhceX
cUSI5FKp6oEMYJn8v89m65yLxLBX5kVjQvbafAo56osUlYrLs5OrdXptjHR86qD1
dxk3V8Qt/7pjVUrL3/yHbajXT52x8IL6HWA/thCG/QzGpX2JQTfYxSThIPnXpKgz
bfPHSbwmfSeSzlnTA/IQrJ5QARFdeL3L5RrEtvoq3JJsVO979UaIeSxh7vSptP4Y
2dtFm0UcxMkZCEiOpb+0Ee9c3w8o1sBBwqV4+Q2tFoWC5Uy9/B6v0B7vlSi4E5uF
NyRV/y6IrR+UjQhL4nm/50OC4VETOxRdqDJPyq1Gk4W609lbQncRBZmAh66+jBb8
QKt0JHG+IEGsjDhejHfjdrTPKPtmdntm4A2vpQx8glLimHxylV0AP6BcIQ21MhQZ
c2DfLMdulw8oxrllb2JLLFgAGQ6AVGIzt1ebsVnHObgQbrnuUuBziYAPPqX8CLfx
WH1uUQTLtAZzOVOc9Yklx6miVQfZlDQL6biDOooNaTnHep8HTO5yNKv5uJKUe+Im
gTBSzrYfsMJoldbakcbJhebsrpCN8t/GutMaSZycxqTDZW8dI0phqdn34eLbud25
g3cGEA8G7l5ViUEnuUuVn+5Vhk0nGyzN0WNbMHcvYS/3LGLzcH+edlH2CKf1cVAe
shIwQpzbwG1g+A6RwPJ2vuHvKGpdQZaQPOt3+7vhw8CgwvowoIVuBhvzXS/8QRDH
k78cJTpOt3pmFZtygHCpntC10pf73iSb79C5IExgEuflVY9V8upF1Lv4HbNO1x6U
N5yhRP+px/PDj4zOi8r2H/vRROByfHNSB2dfRlyu7cEAixnY2C9JdtXE2utHNv+1
eNOL+rJpNi7HeXbP56rDVyEcvrGZX4qh4eY6ZHq9UeEd/vtCqkSsaOcPG3WQeRCd
850u2KL+AseKqqHAmlJ36J4+wCx1oa8X3nCCkBGJNGzYvAK0+L9e8jWicbIPCrdB
eM/m0vc8TuirsuAPxHTwYZLnqavZ8sCNYPCdcJrA8Xt5JZiNUjVOL2d9cvfNhsEy
C0v3kMqtcVASO72GwNHzvdsgtYpImWqqnx9z7aRog5R51o+z6qkwGc3AfrPbbYGJ
XMPgHLTZjYkuGzzJYld5LcfbTQqlicYU08xkFEvD3WFAi0dwkuFcySaCImcxkyje
5+w4JXCOjlttkyYuM9yLbmnRYo5xuguCJb6CW/DszoGHtI5zNA8tiHuGkQTcj5h9
q2QeCOdRE+4AMhbCSBURHyvaTxc4enyKqyotxlOJfWYGoUbFtavUrJJq10KYtHaN
0f+L3QcQx3VR1tgafocIJNPT4HZRv3bzBJVsPQ0x4dtVlAU7mesNdRH5uWcfsTGV
DN6M+BI9aWphG/ytSQJPrfywic4NQWgNVxfjUk1c+iquIbsd4quuxFWOBBf3JWP1
6EZywSU2wJmcmN8trJlZh7ai5I2DSeR2jP3ofMEkM2nzn44aBSIyr/J8Rwvg8uhm
iFbgZ8f/8DXityDDul1/I/pTgZQTyYle6zZDFQZdrivxnDUt8BblQS2U8HDdRzli
6vEZdz4rZzSfUZeSnuJ2zQGqARVJw4Wt9IYkCeTECRpQVdvOhhT6G73EfYH1kafh
LuVimibctdVD0XbRn8VI8dQ+TqmrCbY+7Lf1nHK8H77jdJqar8n2NTmLthgtGNrU
lHGle8To/DdgTteftAdZpXzZXUiRLBID3pCKUnemrb6UnekRmXM0Ni3Q4SU1gzrF
GlePuw3rQn4my596tIQ0dtP2SzTQZFb2qm/GNeDfuCBuWhXoqRV7LitUh+/EE0lt
qqjClVx2GRszo+IUc6dmzHqbHmbCdRkkUYZ7Qo6BExiwU6dYRCWZRjhRe/ZH4VvO
KTG23BfjpOoheaMwTjBEeyNL2wW9U/UQx8iKRtaXnxXp37jry6CJ/OKOLwVsYQMA
/aL/OhHbz5fmQU7wxkxKcDtn8esEnB1CfEykf3jHKZVjWHnLPCKIqyjeXAJCTJH/
27weJ4/Ck5BGdMI0wWJAfO5hz3b6kwBFAbWQvNrBNqw2CaEE2Czlx954ArNV/B7/
J+xjBYbHEJJJ3ZzQdqrDNsl5EUyK3ZlXH9i73YweAM9iQPzGFF0I+ixeyVIMVRlH
unfzPldg8tFhteMHFOhu4OHNcNUMd5SETefb8oREWl1hY1ctSZdxaZguB1QBNJXE
yh2TqukNb5irlLu+6Kuws6O+BEFKFuvrKFYNqjazdmCNMLGUCZ/304TXA8qODmDH
YbhhWadZsSnDmZTl88auNnlVD4wUsCqfhIp5si7fcHimrpw1mngIXs3u1sRhlmma
GLdZeNdVPahV1rvdgUxiYgRgxdv4uYhHd5E3E38GinnXN62IQc8t2/mx/1yJkX74
`protect END_PROTECTED
