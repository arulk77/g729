`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
kBIlk0Q4gBrIQIeRSz9a7xkt4MHU3b6vmZtjGkAc/ncBnYGIOBE7PKWjfWAnRw3l
xIdCvogm+sOFRzOm7KA3WNwbdZ+iPdXFPLzFuD40F+pRcJbcJeqqf3j2pzo5cqWB
Pq1c8IAfFHonAxjRwi0IzC5I4nVxh8VBx1AcpwJF2GwbAxjN/hc2Sdg2Y3kHWJ7k
ynDNox78C85jDrt52L0QxF9b+2gveev/+l0xIwnq/0eQ96agZUhFLR6qXOiTCAe9
2NUCVgO8W1mIvPuB65F607A9F98owA9OBuYFnA4/yjwAyWZFfEt4fP16qxcpEtQm
la63kpqrQe/Q7Lbksn8hJ+TG56tsxLIBSWGQV7xog5m76ueNZaCF8srR7mpgcYjl
gcGVQN/P9+T0hfdN3hl7REZ8Dgwd5NnLuAHCoyH6RdKUYYRWY/keVJ5xJArGUXtW
hpoElIEFmhNJmh7SzPZa76mf+Bz3IvLMDzfDqoE546CwYslp08C5AMh/pOU2x1yn
YaCI2G9QRr1YK22wAnFPaipCzK0L641XZdQA5cITXdqlJ37TF/8UajxVCt8yjrbE
VsJNjTAwBL8gEN7ks7Mhe+d5ybyAP+rt/wjwgDCgmlN8kgLjWwHPaGi48qVWznMp
s0/zKim2BaU0V3KRYjCrIBIC3xd+IY9wMEU1LC/p6kStCN8s0cWq49otlq+vpbYU
2PLHsH3o+BvSz5wO+d4tChxFum9bkqYgstc0/tir/IBZcEwefdgsryDVB938LNCc
VpFFhVeSTU7yUs4q/OIr9epbAiMpTxVqj3u7SWYvwNZH0m8AvVCcxGRtHftqUPLb
3wPsW5eV0EUiHDIewBWLsb5TGBV4y58+364N+zmynnQMgHNvZgC/1MUQq32ea6ma
EN4icupn35J9t//fVcfI2mEyjHOcgcZWSvlhqmFl4zJiWfI1eUNIICFgGPuGt5s+
TCKqCJNLnYXTlKHxoL6jXTvJKAlRp4jGEMLJGVr/h0i7O3owKLvZs4goPnJ7VPO1
6hlJ7FhvzgmY/+deQvvidregWejv2pOqn+iosGvkxTzy5MRDxQf7kMQznAEPrH4j
XGox57MS548Txq4ISxe3rel84kp7QfdZuNlRs3CFxQZVJZp4RRjJqUmkPRBUBqBy
74Q19F7BYcOjNDxR6+jC6i7XjR2nNJ2bQKz7wvcHJkfXmiGuRey2ESLTU7mZy+Ep
+vZogxpuFWyr0qOROsxKy8NZt2/0s2YNAMxmRZi9Jlzjkg2v0m6r1LDrfnp437sj
YD9GXC74HZQR76a0lEFSnFurfkTYIX53Jx6y8o/Dhw0OGF956ncLxjFvCH1+vYSq
J6umnBx5PmJZWEmIVrrUluGK6KfzyIQliKoKGc8Ly63lHEa4oG6h9eq4QT4y4cLV
zG4K7n92iM13SUea2jDkBhvabHqPTjxIJH5vjxfTf4LpoTlFbb8F3BXKMdgYbNYE
ApBhnMz+7Kql7L0r+Z/W4GJq7H4Fe6QJgo+TKItlcKCvruAvKKgk5i7kDIFDEPhH
SG1Oua5Ln3JpxyB8wJPeb7oOLpZALhIyVoSP8zrmscDiYxzmHE1NbWu1WJTo1qd/
xPVjRJ5kpiDyMaZOw6oHAJKpNq5X5ujlsq0lWdzQwVln7yIW3t4OotDSmpwpsrTI
BV5X160oxY9q0mltX6YIbgy9Monc9m+11mwRfxRyRZ3sgRljSerBPQY+AFVWQwD5
mge7YPZAFs8LccyjwPyn7JJaI2j+aOz4GbWK34V9XNpkhigXSBNqIxM/tW8vSIL7
evbM9vk/UMIfnBl+IRdYChCAXSjCEwAgBeKnYgpweD9Z0bQEsnuFj2gpWJcrsWyE
s4AldBK/4yqJCXrsFgHzpCwQWWhH/uPGCDi92u6IFec+AX3wrvxbJi7DlokFCIjo
fQ2eqMkzyuKTcqYtUR7bsRcvwwGAvd9CIS3vxu3WqufyNK8WHt3C7VgAOzEnPYeE
8F+2r6heEtrHD0A06dDpNYNsBVCHA/+jFGlDPboif5vVN+llzk0SF/byjWokEY4S
DKv7fzRnnr0+To+CHGjmF5p9PVFsujZ4q937rwbtGLDkXrPrlQmij49/hKvPR4ZE
Pdi4MHD4Q2qIwnpY5cAfJqtlY1W1CZLPtvBuVHtJkqsd2d11iJFz0m9e/jR8wlEy
AHCDue8UpGVzJMfdupXXjv0Ec6h2sh4uGw87QmjD8v2NHwRIGUonHhX5K5aISEyK
PZdkRLG1p4SHCHw/l3GKl867/zfsRNlx58fANMjtMiEac7MtRz5+WjI/R7+3Vc1z
YxrF7y0MCmjyXn4LY+AbYbuk7R7Fm0uv/QGTbHKk2w+qeIbosCaBlqGM8rvhdgSF
3ZBm8J0JYfQu34PLCh3WFWoAolhmNyfQhRneA/N+2OtQsgxRwPbhtGSVbosNfCrl
0n8No7d9A2AhswdwqsBQnMZe6y0ElxUwWZiTLY+tcltbVodZ8xDgPrloWvbWSNk7
FFUD5Q/bgWyyxipjr2bdyv1OBk9Suhn5072ET3ppUoRZza+B6DXec3AW17mSfWpk
aSKbMOpvUOrILc9ZTloJCTvzH/wIKDwsiKS18WCmG/scLCh7FwE02bwKD1Nd63s0
HxjUequQDJtirovxjLIWbLPveU/LyLwWn3Aaox1tzE84LcqK1NpADBA42jxsdNTl
2+ud02oeC3NfZnMBijzajci9bvRmRcFp2raFcuQLPmfBrf82fPzRGGBmByCa8buU
e3drB5VLv7CxJ8RQjvbQmJPsGbNkSCkc9LnL193I+ZhFvCkidbxgNdTWzc3mKccq
dNHYHktYFBEVcViFvMTGV0+mB4YmkNxFqcSm8rGKGqTOkFCt18WGptxmWxvWrpWe
MKvHA8jyt75GxM9yVHJ71mvi/gnWMD8XGxxzuLqlpvcrJaJ1ExGki7yVM1NhdJGf
ihP87JLGDBk2rJTtBBflbkbhd3KhQwrE6pJ/Wimbv0YdJYA8AdbwtMTE8OC319ki
X3um/rbUUtxcCniMBRQZMmQOPv28YcUCa0dZQ01VVtNWrhCMCNpre/klsbgywfmW
wf17EbuWnJ+qUBs4Y1fu5iQOKVrC6/vbVuaI7vta0iKGK4Z42x41D0v41ToL/vI3
gQoUp8RDBLGNRRYnmt0tixHClsWDbb+XxBxUfJujH+EbgnefU22i4H7nPjc2LZUF
ka/F2UjgWvFD/ODKnCuaCDoXtkB/tKVgpTTp0H7kCzXslRE3+4emg6iJAK9RZttw
a8PBKajBdikKGnN8gmm7OpqQr2VzeVrX7iGWgC6aRcyDa81TpdRgH8z6R6/pf5M7
6mr/qpyJ6n5Q2/Y6MmUU3scImbZJnnS5H0Wxu05r0seXEiv9rbO+dCGsqInXqVjb
CjnJ2dP9vU3HiDX9LMwuDVCBmOLk/50cmGDGNPpYwJ7a7hHAIHZ0jtK/6CiZDLFj
H8Xt7F9hhrXnT7eDf4tn6CuUQY6HzJwCThY9txCUDtRdQSQS5wORHTkEDNIS8av5
PHPEPho9sqJDNiB2QOcsOOPSgjT+lb+rgW4gn8cG+3zw7LKaTJ5wQU4xLXYrGKCZ
fpSwtJS+Vepx4iuGH9kZSebHV+RMZoG+chGqlX9b4KU9x7B7wqroo5jG3J0DfYa9
6ekoCOsNz/JJkNxkKWqiUab29p+XErA0A0e0dyUgp57seY/xsfjGCWc/lPSdDDmv
p2I8Urvo0x+0rmNupJJA+Bd1KTxiYfpLw6GMHjZnN1N+LpTFwJim6PpxH+rWOWMg
uXFpMCcDn3Wrx/TwrgaRB7LgQaQEm3xB0ImtrNNEaYyrfjv5mRZWkscSfRu/yKl8
4Cf2lpTrED/VO8QxBe/osgKmFXP1MiDtv5YpRVjJVS+jX/bD/LZ7LI0pU/QQ35fB
aq90/miSAiiu/v1/GofondygOlF3Ua+Xv+qI7xaFe1okEPBSLGcEapPsDQxFmFT/
AasoM+QMPgBPIC40dOq/QJ5R3UwWpWRJd7bBXLemDsceu8EYn80dUEZbd8JgrA6Y
ZVN2dOy7EszIDGqouQ54nvXonMEyKupMaCqHcu22lEbobaNIldVIDGWqsCci41E6
yd1+no4clSiNdzErewJzhYNSbm+tzqbPDaM9MpvTHM7OJnGytMbbF+L98vJcQQVN
0RWeDTDWWXdSL63Ip6TS8PcM+vlkZO1dOBCYn+3XUS3DBN7dCs/HX74ErV9tDnfK
szvinVmRAIFEjkenMHIbo3IxFdhdB345Wn4KhgE2Nqgfb+3D51+Qw5K6GoRnhQFx
UX01VANZyUNUdiz1keD+ddXSfdSrY0oOcct6MKEfDVbpyLoWNAcnOM28dtzLygjn
juqyejdrMnwhVYJV+md8EeaknXNrVkK3dUCQt4DI8zH37IyRYZyGeBDSKmrt1EnZ
keYsjqP892pICykXTLAdDWwzccd6t2x97InHYge8chAkSckNjL+tJySqmO3eoDxJ
2i77GykWw8Bky/dipyNQlXrhs573Dx4/QLD+kx8FZKAFOV/SU4OKhEQPnJ631ruQ
/Vq4tJflIwp8s1yh+4p4gbSsv2PGyq4Qc+kbwAH9FVa7UlfZdqaXy0AAekOt6oOU
9qpAcFrNmmcWTVsrdR7R3CCU0BFP89h2SaPFXZuItH0f+mRpcQnLXNvQrZZHSEwe
R4smVcvXARv+uqwkqgJNgNsyrnOpP+C4sYpoU+OSIR8BVvrwjjgEmQQrzCqcrvvo
8fl3ntWMGlsdeXEvugEXvVgfoBykUF3iB/5eL0bc8FS/XH2oXhBWeZGSWcIJ2gL3
9pExhb2ulhnzYjkD87khCBQyEQTwxBAtjgli+uOihUKuPWYeuulheaRGBvn0igYo
YJelQF0/ETE4wzV1eVcScKuERvFJRShXtX+SNLOKkmDKYqBx/JMngP6qLCLZXLb/
u2xDhDKJmxFKN73oGAY6NgqxVkJidy6IdyIQpV2ofktRPs3mLzz3pVrauUC/UAuM
2BFEB++uXqqqTmlhzPXL+tCLS4Wz6o4p+hDWGeziLkShVgNf2xxW8LYsQJxRs1DK
4q5yAdU4nIrZzFqswS0gJpSTVLOpPcRtnXTnjzcRV7T6n78a68oSuVD0v+m1mosE
seP9L42wbsvIjIFru8O+nMb4VY31y8GsIoJ9i66ALExa5qjR1krBrQRYEE03qskm
YAGH5SGZe54d5SKioCL5lBZ3HBrkNNWoUNlhgiidzXkwF0c2k6AvOx4R89DB+2rM
EQNEafHif9TdnheypFtZ0bz/VNU64gzP8pNQLN836vBbTJNKuwLl4cWMftG40TKJ
puseozOYf71icIHJp52hdt/lLapu0Ku0mNTn2IxFB4jnfePS5EX39Pt0QSaEijPk
sOU5ss/PlOkyny8Lk9GYGa7FxJvYDR6aev8+AjHvDglZ9rV+aGxKv5UGN318l0Vc
bfjTaJbIQZqRxVxotC4Hf7pxR7mFAHMt4PR67gZzQDbPvD+pNYqQl6mLGVEBAuLz
8aOmZQq50tqvNCvK36XyR/MbRjFSMWVz4FUTBJ9I5lc86YF+8JCV3b4obIGNqLjw
r8mV/16uCs7gZdcx2YIEWC1XiiNJtXhk2YLLYd5ceYvt4JN+v5uppR0WWXmbzfTJ
PZtwrBZEXKK32M9JZOB7BN7nv4Z+zm/RE5AYll5e/wbYJajLJcc2mIqV0gTrKIfZ
XOnBMyWxRZqiLSDngAEP46FOGHZ9n4cvM1POSXITVx3HRzYcsch5GIe8xdQPbgNA
CLhikZeQGxi6PtdGJm11F67ZSz8b2iS/5CK/EY0wHC44uA5W0oe8dL87Y0kq8FaM
QVMdLblnsdTIfRhLo4/TDNtgnvVYQ+jFzkcWuGqTv/JXWBCTQ/npmPcv1fdiVUjt
JDbEYWXr/ONaV+NO8XUxrzzA6esozMNdIiIkFuChUtMw5FMSx+s+fTIZFCStxsFG
yH1ovaGvgdzuQJwh9FiW2f+LUG6HE9ZahpUIyhGRlG1ZvB2eH7VkGkjsi/OLCwjm
qgrfCywWDm5cXiY6nrYBG0imwS8JMyNfW1Djn6UtL4mrB0oRHjOoAgMKg6Ef/ite
7zV0T+zGkrnD+ocPC4+yyJvjibEDX/47rhQFwdUL5GRJ/tMXnUjbZfvZXDWYhUTF
MbUBYC8srzimVdTN1JgEbZf6LrfvD07S+gU719cpxld89in6zjrtiUVzoYL9NGAu
4jFKnjqOWGp85kL855u9R/iA4wxKVOGRQrIyGWNZr4GsWDC1NL29hlf0UQNuSLQC
+mA4rztc5D1AXAq2SQDl4AqT9Q/uXZF3QS7ChptRW8VLKNzMVzhOz12dGvFCJFcc
+RyytCky/1fln7gIH5sHJYHU4obabyZmwP6+M9Nh9q/riM6E4bQy9noBMmREROMJ
ngD3uvlbTZFe49uSmceGtRsh97BfNZ9pdAVOPaY/jORaNOAQV9ebg+S38ddfi+nV
2Gqz4EwRuv5E4QI+UYywkNiq9pJKp1iyV2IYdLn/xVPigcct/kcPoZSJmeCFkx8E
JyfWNpWRgmKDktk2k7y0dOnICkV1bN0vYmGggGUtroOfFuKUxqgbjXkMGDpNsL9S
PR/wPd33m9FdgGmB7BQdds5NyQvxzE5JAzKEf1Brkv5uoX99ue5PlP4B2A787nfO
e7lFo96CcUqi97LzDFOfMuB10vgfTZuOw1UyaFOm28vuzQeAcNe1Mtuh5EOZBmRy
mUCbLr4qS3yTWtjZRD0Liaobr1xbzSti2cNao1J6BiiQJBsrOxLpylqTTqCNLSbt
TU2QQX14HvdQqRUtwviloiTFYJ2UAjRMWF6Xsoy2+QWF0jTxHnsEk3oVyvDfeYCD
aXBnMajcWwDqTCNseckADm6MzdEdxUFt/ELS6qMnMH7HyeuWE2bmGWEP1wxMA3p/
zjckNLuz8Xt7lK9GM2MmmocMhhyj5rgP2u8WC2X+OdezDoBjpEWwI/98m0h8w1JC
d0gXNsouKM54WOrizf/Cpks75blSlQGu2QR+ofw1zjiPiDCsDIGFfloQ/tPnx/DC
96373EeGzFYzbwmgFU7lcvOERd9pd3546L+kTYqi9Qgy4oc2SNmXj5tvoX4fYnT8
2oxDLPZUZR+G7MN9lQNzZWnrb7lXy5PkjddAEQzxAki2HlsUI0jSW0VSdeYlukfB
tQXSZPgR8LSIUfAx+3J5q2cSQOe+B4MUcjG37r91eANq9dm1M2FOmQzCGpuJPESZ
2c0S+qPVjgLuz+TC4Z/2AyAour4Edfhrypy35vfZKg1PW7muR8CdhzeN+iem0VkK
Dc+A2l3PBUQCyTZFU5URAsSb7PaGVLiMXbYIyuTYPCqJTwQ5Sb2FQdttJNHdI1wb
VjO8ysrVwYFtAWAPZ8MBFLiafHzOlhO96rLRGb8O6yovMdbv+yLpPGkVvbUzKbUS
HZ9xSFyiuQfN2uer7BzJTdcMiqvjejRvKzoaBAZ5pX7oglOAMz2cvWsfCK0McbJ1
Fmj2WnsHN8fKVOU3eLOuwQoC6cnigWmaMFR7PG6Jl+bpm78liYVRb9Ewx4511gFn
V5vKJd/WUMZ2YswFSmycMYGy7lZfGa/XyFLkDGHGA6Dwg475E1mwCpGRfILQYN/d
zJhQRO9YMFTz+6Sc2zGRmA3upDL1qQLQBiVmBPZUpk6WbEnDqjg/9U+IzRui3fab
MMEqQf0VdfVk5uWk3TMz5cDs/TsdlLYOqH9T6NQXrolZJHw1cFG9LBb98xQXhr2a
4wSHNt3wWNx4S3RsZ2QQCeYP9MWl7Vg9GKAS+VsB6VGeJKuONiM7A+j6Rrchqlw+
SzDC4WrcQvwkbG7eBETfyUxXDTWmmWeHJT9IHQVrQ44Xd7o8BYDRBN9hsFYrjLi/
VNR8KEqumCFx88b9Etp054Fg0VDGyq/PHfhdewWsFRDeW4ACY419GBslEzf0SfhR
rI4Fd96ogHPebbnGnLzobBHtK8Yw98Wa5ftmrLDAHvInl5vbOG1BUfYyKCnEgs1S
KswJnlW/rKO85zprwHIKcl7TD+f+UaC5zyws2Ubo+XEYEE76/aHIaMOBk0PiHqTp
IFA+SNz2X9hDgNQyfmhGtLeu0jDmAodGfw96Llb3dAVzwfbgOZvVC2CW+0BCJBBe
S7AejbzfaPEu3jWgoNZJ/bPL3Vr2KqvYiJW6mmn054t7ZJztoprox6ORg72hKeCO
MHYj/DuOoeQZtOLymvV0pEmNxuBISomZYl1kFqkNl1HWXgKIf4iIR2HyZhdBxFzd
PZ+bWpTdxbhrknJkHD/mrsvlTvpENEX2/cBRQANavJSvzYqw/RerbequQTEIQE6z
ZGXg0WC9rom97Wf/MFTVlOl1sT3WRPNTnUmT/HLceZRlndyFABLhJyk+Tco7ZF4H
qUVZ5laYiYS1L4pw0mgiBPhcwYsZTLKNS1R3wV5hjQf0zarwmzmFESVkaUz5za2i
MUK2ilErX3IOLf7zXK6amE5lqz/wk3Yaxc/QWOy92OWACjBpzNUnWblA/HiZ7ruf
uh65+8TfZ15JzEFZPomznXe2RZCr9nz+u0rw3/muMN/xy6MLbHw7zRINAsCEjpTZ
RTKtXF2a1WsRye5EOyaJ79uNvygF8v7OKn8NFl5qhBZEFsCjOxnLzflzHKaoUBXY
49A14kYN4uE1VrFIQTjF2FfDIZEb50Uni/khveDaA52bMiXs+bQ2oTxFqJjDZkVa
83gakZyJxEwxkrlLOEf2w6ZW7/yyYeNB4TwwWJsDVgMnUI9+PKpDkj/sFobczl6M
N7vVH+RrkQDwUbWX6jlvJQNr+QBf8uDsk3awB7VrcuYSyszhJiGjdFTiU3iLEkvr
LhUSZOxsi7pu/mu2p3YCspqZl+o+MxnHdynzqfG1oZ+YWhgHeIPOiflttOVUzjMI
gfd2EQ4xuk69uPxidsGBOoTNIiHzg3ouIKC+uh/kyvNm8NRUM1MyfhNI3nhcX19P
JI4wfI04N9re53n6wG0CpeptTdw86RkzBZF5NNMiV7RqYs8UvNhmsIN5HyOjRk6V
9w8gsAvUUq4DN9yexMaeiG+ULbjmj9O5ym8Rn0C8EIuNPKoq10r/OC9lUiqExMAS
UezhsZxuE5ZLHn2+pjcdQI8lfwcAK/PrjflfiyiMcb6v+D7UiPQh1ngQ5zeEvX1I
EDE+P28/VdulfY06/fz9CxY8RQqhxOVsHHK1yatDLmgfulxH1VygcE+q/mo3Drb2
7OjwayNXVv08cJit450+PDRa7KX2+KxUh11tujS2Qk9nwURBXDPKD1z1zvHG6rJS
ZzGn6vQocHTdwglH8Dri3JN4sGG39lEzP3gs7hX2GzMyfIqF1q72tKYlSaQh656S
PAcV8VVJ6hhVG8oUjF3muxY+nZeukxJ+kch1HCvNWsQE1UwYkISN/EqOJqvdlJNI
CiYup8aGHupJTkEFwALksnfxM3Hh+9YQeGR7tun5L1uP/5d9RVTRLSX837sF+LOg
2jF0M36n5yNObdbki1LQ03OgE2EKDyebktOrz8/8LkD+WJPUxy8TrGZ+9ojydIOj
VvEJKbVrqMs6xnT1YoAdfOrPbpjjfKbgc250e5VogRcSErfuOAlnGZKRQbvrXMLM
Iv6OfWQpUlXuPsc8w0JgeFlHGs47HlwHec8Z8c2nWt+vOvabzVgiahdkM7A0CVCe
X710hSYKtYFrwvV5yqXAgH+rJ5T8HpPLdUQo54Y3udT1GFQPk+b1yA84CLcAdbvT
J5UxZT9UDpFk/p/0cdC/0PZhz9ky8RqsnQXaBGpoK6UJolg28g4voVIoT6tHv5HP
BjxgAWcNms2dYKQoeb6PlWU12JjcW8Gk5tpnyRCovgf4Fr8xcfp7wPr+z7QZVmdn
oN5BmeF9Rp0om/8YPq8XMgzklNrw3b7nfAyfFErpUtaFjh9WUixlO8/5vELNeHhj
2bBQE1iNdszLCY3Jhx5NUc6nrZ2IAHUrsHl0Vm0qGeZuIYnT058MUWTLq4188Du+
W+KotJeFNRRd8bqfEr6cxwee5TWcLAD0MbCOzmsBZP90Cd6gA25TN+m2TF0sJ3yg
ArgLG/9Aq9mOU4SP7so1RvngDYuHiGb8ErWAiOOvkp7eaBXvKbhaylYPyd0Q9ozF
qsb5GVPgWpamVG6JpHZZ3a+RXIQ/LJbaF6X3Cl3UuD1gLAhZr4FG5Y3TNo9BA3iy
oknVLIrCjCTy5Zu8DGmDf3Xpb6HdKO8QoK+Z4U7Jeg8O3xw3njInzgmAUC+SWFuU
zDDZuGPRqCgmsZvMJBgH0okmwmmo9VT/1HZSveuj0+gaYjm8Sml2r7NWVpOk5Z/q
x/VFil6+EsGcCOqNKjnXatovp3WjNyhdvnwA1iNKca9jPGwC5VkwdRISy3LE4N7M
tpvHVTPyZvgffq5SkdYTeXAhmbqk3isGdrKccQe5167Ahk6mB4Xi2XXDKofIDe+v
WOgp4dWkDFz7Rv/YGzRHdYtwLaSbAJcvYOiwMgrN0mbeoeiFrDhJcoBMznA2AKcq
p6VObAlvDkLOPvk7NOr4ODt0L8xI9KvM2uShB3ndedzu8PkLdsOg+7RQFX8yBVev
RRiws5tk4MOmuv2Lr+qXHYSlcISG4o+8ZAKA0yr4n9K4wZgmhiE3SXWGtxd28Qaj
lbwCaQhGWeP65qlndBI0GuliOoTFcGys0VRNjMhqt4JC3bPQRJQ3d5+wNhYbO7KN
1RU7gm4fkpaZ+Swnph7KxCX2NQxhsI/LJFTkPkmGklHi390xqnQsKSxMUIC8DZ+/
JZN5UQjtHpOgWscBeghficcz9XdHVHLXIg9cRG1CwOn496mPNWHGrJcuOMDYjOxM
jc8yS7odbaciu8SkJ6objmm9BXkPwMai4O6sagXAQlSa42zQPc8QQ5B1Vc1o9Sgc
A+RK/O8ZuHDOTmhDL5kEJHi/yxqtMvpwrnQp2nVfULQzP7pwikK1aeU3VO6z+FGp
EK18bUVBJIK7FncPshWj/fxK4gKx1rekKhDVSJirXkDOP68HSU4we/XgCtjd4FEn
WXzpxKDkLInE/JGMet75H0FAGlhPvYwiA24mWBfkUTU2PQ5+tKTs4Wikcb5f8nWg
MO4ZAqG2JCy4sd6Nz01ffA==
`protect END_PROTECTED
