`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
/ZI0J0XsCvMJbxqbWJpuOlRp7RYwPiU3iOrw3OLgGWgPIwyvH+giBMMBYNwd/pqp
XRw3Khy+Y12RfsbpBlol+Pu4Gsz9w79oyRs8naVOuuRY70A6357rdkk4suH0j+4t
G8U+sbFkUkBtjNjcEf2RIKQ0SnKg7KJCUd6px6U02brXKhz3GfcXE3FVI1kDehNL
pQO7M1D5ugryjyMfu9AVn0audpAOVSGysX7EiWuyzixbUqlGEdcVQiRSaCHeRE8/
W4QaNlzVG4+WpaTMlu+IO54Z5JeN46jkYyVk2OZLWEV/m1lufYkAum/tSJlT0Jlv
`protect END_PROTECTED
