`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePj3BTsFTcSzsDScIy49KclGpFDDO8TYqBtzfmgcaOQH
AZEym32aDiezngnD/a8wcSU2loNalRbrnDAQw0dbqpQJnnM4R4m+DvuHSyL1iOLo
VRG3VbsfBK0s7LBY+qwv3VmOdn3BAm+E2Y15EHKkboa43cD1flDhlE36moBXPR4Y
pTSU6iIIik2Yu3dDrbU6rPiDFzs7wVOJ6LHCQ+DIzn9xW07K1RMDynydJQc86V0o
hRgo8Q6//E8qXHW79T6P8HQN6yOfuEpJhgact3VOh4lvSPBYg19pTPcq0zinOK3A
+4iPKOIksi0qYnWCfQCnVzZOUAfbUjOVjn0JmxeJkjANprqJf/7vF2nRn6r/1PMN
W2IGdmYgO5s8HuGdAhGcqx9HbZNQ2FyNjBDsfpfKe3ogrWVfrmzzfPu8fJHyu7GB
he8GCHOWnUBCscoUOE0VewJOGxErZiyqVMJeH8t+iFAed+xncDprE9RSoUn7J2Mi
`protect END_PROTECTED
