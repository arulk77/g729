`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAQtn/GSkJc1bEPPrl1677kD+iJJSJzyEitxxhbws0SJ9
K4UPw6RoT7rXgaCL5rs6uaJZ/cobmqCMLRQu4n7smVE0RT57b4SENXg/8IfyhAGy
AvYA0CfPbKsxWb4wwBPcMI7Zgop5p5NKWDawwLxbwRqITvT70ctqTSeVlLQwm5Ou
8bViywisbW7uYmPEb/XGFPN0KQ9M+OQ6coIFy3DoaOHaTA0tcMqOoJ0VrP9IRtDr
elzLWfDdP7ZyyB3DAE1+xh734f5bqPd9TEF0tUMYPUf63F1va40MovUrhJjFsACa
bmFihr0IR4n70MOFmUZeMN86myhKS81GFYg+lHCbAnQDB4Kr2LbtsL78GBhz82iF
yBBBN1vBVNiw2z3tIfntJnUJHynTEGECTzopyP8nEiGciSjE88HltGvzgKveZcjT
7vKXySk1Uh1csPA+EPOvkDrjZ6zAjAqfpV8yEOSLnmjx8vSW9cdy+jnQgRfptngj
yTKtAnQfhlsboXNbUdUf/OF0+Ah4k/VexxG3cFvior2oMvGEPm1YWrEAewLgFkug
ItNQ7H6zAr1jMxbo0elQ0M5Kb0yX5r9+r62yzlrZCXb49qZSXyv9BEJ1IExrAaVM
C0AQKsosoRqsUS622ihTaY6TadvWx2lBh6TNwfqojP1P7IA5TbX7ay5B26+SoCHR
L0D6qtWnfaqs0UDy13n5ykWFLbD2BcEkRZGuZVgad58aIn0ZTqVO/SOUE8Xk/vxV
MjjO2mGKt8hOviaiUr8Z8ZJWOmm//ACvtDaSAqKm4K0jIncoTFRo/YnG6ka2mjsN
7foUTN5z8n7pAqmKbh5qmw==
`protect END_PROTECTED
