`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHme9xMkW3Oc4QjR0F2d/Pn9LhB7sAfWYLYDyaEt8bm5
hbBKGwm/NJdURWwcrCW1hfllz1AqgXZy2VTs6Z+P43BH4/iYtDNn8hDpXaqOmNpK
tGFTgNt6H5E8A+VrXvjfUVYD2iRxw4mJ/TnMZLh9piAVNWkxN28Irv2TfNDc3W2F
yr778stC2kuyvyUbI5JwgA==
`protect END_PROTECTED
