`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SV7zW6bzZSALuY9OnGzJKtckOnRwwz1oD8nCSLvfFCEs
VQ9e2PW1zsCZO6hEzmYJTP9GtEo6+fbfBou0Dif7U/Y/ilcjpKx1hMUjxh43I471
WCjoQWCUrxYX+SraEy+7nsxpfYnfZEHGOMVCrsWVTj2R5ON0TZNkRbxHyB6Md7tZ
AgJ9kS8yAv5EaYDpyoQxVzNePSuifptJQLTyyRb17hvRLICnVVi/+YpBbeir9gLM
aWI6iB6345k8IlhZuNv7z/hUgaFEc2whYicJ31z/D5nhzDxIHs5+/7BD08Qeq4RY
Bam7/P9w8msQ5xtp1sjzI2DEy0+XCSLnjOldSOwSOg40+nZtN5un1jZG6uhUMASk
AgkH6OFinRT9jwnaPXkHElzNTaUjlnLQAPh+WtfykQIzF3+fVI8tua79fQXdz4AR
n5q68rz2VxeaTmiG/FlZm6K5FDmkSmVox+XUWcs4KX6xboimKDhwDZeaHr2oHTVF
SOnUF4a7BwUkijmSrTXKXotilGF/o/QTh7PAszsdTdONMrdKYDfFWmvZxLT+Bw2t
R6ebFvOf1jRF8rzEyH/tftb/Jy48F9oe6yNzYKTDIB0HLrPxJjhIBMIrTWSMKkMT
46XuQ5oRwIvI3e/eHcZntQJo5SsEKCJsxjbfynooj19ExRwTZCVOIUDgMqEVjNDa
AwDINgtmKd9yd3PIcLnFkwya0W7IWHJnby/PxY+wcHwlTCqV9TiXZNP+DrlBWZLw
QBKpfLBG4nNW01Lf0wpsbuEP3dqs/ngi1gYV09V/vT6ZLXBIv3jwlkO6jV71uXc+
qyIjFMHUP2wUWK4GAV6A0+IPSySBZjzEOblIhH152XZOTyD88U4pUsSTlWbC2QZ+
B6slsWctzjsEUNjr4w23JHu0IJEdkPgBx9Ib8YdNamN2BezDTEIHWuoMqPwBpftO
BwHPqrk3+aOG25UqNrdoe4T5vXPt0K2wRC+t7DJr2hXaFVP60vfsk8Mvk8bPZGZX
nymFQ1bHmEOYH10t0SEiKqD7azgB3bz8ZRYCRsJDRlhnSmMriRfY99b0T0RYv62+
geaZaYqI3nzqlKMDRHLfv8Acut/ddxcSdGtI4DAgXMSVFqa670Re7dnfiPF8pO2L
bcV036v7JTpBS7N1OkCQoeYgDqh7Q3hu86FpHcddjextd+XZDXCxfSbZKZGsq/lR
pCnYuV/dnVFW5YJ7M5l4T33Fk0ayRgI/ywbhKSyMyGiEMkxGDwo5piUBUbgBbRUi
8aBa8wBUyzJiOfabATZhNR3pH43JwHPejqknYfmn35TsZvdraykI7vaJzS5aXEHu
beYTFJV/WXfEYkrq8KhdcB/D6Ycynm6VV1OVToy2bxKmnBoUBef9xPfQWUBHsDUj
CLo/Dab0lS4Cc6JVie+pZsKUv4MZ1QWdn/rfWDLiEujAjP+WkP9CEca6QbYLIzXr
GLtNeBKz6PM5vOFMbzW4xp6fc/xYOpR27aGNrjWNILVmiwraplNJyDB/5x+2NGGv
kvwllDqyPfCMz4zMmUu7qMf8g3QPmCKuxaBviNQh8PG2StqlL/oeLf5KhpAMDQBC
oFC2axkUh+eYmx7XT+0ef+BIaUXWmSDSwUvMtsgaFD4XHmAe7YN2vzXGVAQoVFTx
Q1ztx1BiKmlPVVUjllLwit0jTLKt9UpAI/+rKXPDyxdMOkvtWPNnhYD/BE4GdubU
7SARc+WN+sDIlKc9ZeXvIXB/FUNeSaOdBj00CM1IVXd7kb0+xnGngTiQsWdk2pFk
uWSIRWQvzxtgOkFEfNa5W4wlLxjng0twHJMcPfArj4YcWuSZGGck387c6oRTxsR8
mTBrFevwTwTMuE2+PYzeiw==
`protect END_PROTECTED
