`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN8fKmOcFlum9QsdYeNmmSSc3NUWtTa78sgJWt7tv2fW
kP33ilsikt75ll4+N9I920qA7nzuCNXUkhQRchizDc2nsgTNKGphfusvB01o6rUx
2qlC1/MbJQQIJTUV12/0YYmixpFpwMPTYg9s0fN9yp9bdU0bD0Zn/J4FtMLxwY/W
B61y6x4eZtqWXdVZmZ9ZOBYI+dxYPb6/uROLun4JUuoU+2Tab5uBpaTgKA4BmYkE
tY72Ki9Zpc05Blbr8Rb1xfzMbEsXNRbzkM0KThjH4r5RzOH9lDp+g0pOJYOHMBz+
`protect END_PROTECTED
