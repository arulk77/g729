`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+h/SPN1IPUBy0a0Hu0P9ejazGVVW0niIdn/pLny9FeA
gorvRXvIkG5Ys2XqrmMlqOyW+4WzjG8CPBxlSz9XMfFOZWq+xX2h6Bn3DkPitQL6
/PhqFumgMj80V+UzdmW8wLhZHlVLbclXfSBGP0nlyMR9pL2812I6vBfBpOsqpzFE
4mW/vY78vfpZBdibtDpwx4yC4eVBDBYksHubB5lQ2YZt0/OvxgpzJJy/cSKcqdwV
CD/7tzldhaUnHiB6e4zJyqAdgHfxLZWy8cbqVGHSG9o=
`protect END_PROTECTED
