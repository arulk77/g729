`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu447ngNg7lDwFAqJBKrIWBZPz9ww8/I7gz2MJ04xmhIQd
LwSuLMDaDxTZxyp5tazsYaiYcy2WqMcFxdOoRz/7ZYEN/bgc620IQ1H7GtklSjpQ
QX8kHwYEpTs+5lTR+GTViqcEeeDwlCshbPWWVF5YqY++NJoAI/aVENwnP/zw68Mk
Umct+u/NshZ5XlET90UMJXpUN2kT51gPGg4ZXR3/rSMe+hgIsnCPnOxOwBfOhVe9
5oPNUHGgyNaB8F4lwGBLGHIYuH5h05YlqHLzP2RB+QQiCCc3+4edvRztPoD86I1U
8GF0XF+NFx/jeA73vVpE0A==
`protect END_PROTECTED
