`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG1SKVxwQJwgNvsu0GiZE+jGfZo1ag5GU0NF72Wburd3
PXR8erkpnke6pwD0JKWHumjQ3nt6jA1UPQRGgj067cQ2e7wW0EA/yvRuM8WF8HK2
8h0sSAsWmKJ6K7W9psMk9U+QvKoe+RU/qoJu8B4aRN9lc9UOiz933/lmyvZ9jaWo
`protect END_PROTECTED
