`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
1fbfiBNS4dcNIs9fSZnFuwmeUiBFpBdfAGfALCvObio3Ryrf1VCHhQw+fY93DkTS
trs3w3TRCMsv0iELfWlTWBTHBAh5w21++U0EnnP9JkZBCzgVSC+7RGIWKJ1AAUP9
o2y/cTF4iExpcacITbzrThalmAlIR8PRAu4vr9MewfOB65NzcsjowZQXitaSDQPF
nd7l6DON3/SdL96ErcBb7NiX43B793K8P41CWM32MVgTI0X10AqUnUHrPayRXi3j
ZTxA0qSfq6PJdCm5airAPeMCF/0C8lQGiMuvczB0mB3Cv8WR//nr3M4/QgbNVFjw
rf9lJbm4zM1Emi3A8z2sciDqUDECehtui9uMAUgLUvM32Wn6O6Qod3ytSkRfAj8b
OEwd3eVD3UIcKL+y8MtErKJqIZm+XTGLHisxyOgDVosBhrNXi2yUGOrQXV8IrHN2
KpMgbRV61kSl/UdhKaFL6/XN/dysperjQQ5rDbez7iD17P08Dfxjz4omGs7iMj6P
/yJhJwWnGg3R1KwI4YmzUmLd9wjY7pvyiqDpCQOCb0/ylR7CBQz2gojfvHDFW2uQ
wBTM3QNHNM3rdXb8vB19aUvDlcxM7AdnQP4rBr0lGxpEwjwVzZkDIS5punUMq+9K
SFcWZ5ZpvsYxUgCxSgRSae33AKjC9kpySxzlnDkATH5EYiJDBzp5hx1Bmg463emv
ZwPKAH/sgsegxSB5xl22bJsT2LJyte7sHLm6B3P1jdun+geuEWCrbhSukkAeD2+w
OV22UTadQdfbcWhX2GpENN6VVAWufacuZUxKEuZ28hC7xXEtpmcj6HbOZ9VCHxRm
um8laOet6lp9oG0AXIY57w==
`protect END_PROTECTED
