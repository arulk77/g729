`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
8nBJ3pbIPff1Cqd3INwlWoTIxIkQlN0qlTwLg4hU1idOVhiyzsM2XfnuI/ANmWra
4z607MJUolYgvFnVvGKYFXnbIzDN8bhaLJSkbB8OiKF+JgJ12cU2IH9fC9n+TRil
pA5r6gxsFITd6iC6P91Cpc9cYFu4BzzDDvkjht92W6VSpkChOEWcxfitGqtY+5E/
T1jnHx+vyQ6z0kTlVtuNWxqtkkvvdbF+TmGvSHMbRC2uw0tJMWeVop8ot7IyvZyP
VXCBm79vb2kHkmaMt1X8eq/zfJ+kAchKur+gjJwoc5OVeMrNJsL4+gXFNv49XRD/
cvMar7chOgeYKdB5ruzPwJE/y84DnNKrkk50v07UlmDDQ1WCC4LuVv/mFPEYDjQe
uQwYwx4Qnjjz+V5SS69zYqs3WiDR5zbjaZ9Q3JcczbK0B1VUF/zro1CFYCqX55wS
mabAhmMXWjnmPegVeG3n5NxRHozvJTThsqJCQ4rMvIyziVgccPxrxncuLJdW/S/p
uk7uKVsIRNPZqTTVlb86xnxBUdk0crrhFna3R+RREoiH0+uvS1dk9kBY9/lsmX0O
CytT3OJaZTnY8NOhDQ5D9mQL28EwuY5oz87NGCdWhkOtat1EgjxCaMwwR1lm/Whi
9Scehzac7Cz/xNYhBfSVFA0dWBlsfNWS63uzw1qBpAOQ4zzdkZKt0IeCxa/hpU5s
VoMZDZDwmumCvjX5ByvF5TE9B1lJd1MvmBS80La4Y04U225HXboV9RdgoMFO2/E+
4x/zFdVeVa1I5/yCKMKcxasfOATz/VnwlvT+3RUuxnS1VpCUYDovLCr1Ar5RPgSX
z1F+dmyvFfNs+xWor1UARQ0+i6AX3nz49WAdKg08Hsmrx7r50oc3LwRVBsyQbnUe
qrIhzUvP9RA+0w0Ud3+BhnRkOOdqfmFVo8VN+qJH127KN4/Krm99q/kErJqGOyLk
xrOXrQvVuMX/Xro1QVAdeHbkXaw3inDMpifisd/9yA+YJbtY8zGYFcyDMRBRd5Ro
409MZIq5gUTZd5/R9fFFAc4AIVjElPzUu/jPEgOcvrP1frFQBUw7xfqIX3GhxVHY
VCqzA1Nh8vNLyGQavvLGEIe2htuNK8AP0Vcc2T3Vmrl5PJjLVfXxLmwMgSaGnurJ
qS1H7UV06azUSevRIMkenStL3YYlrTyvZ8w7ryytb74=
`protect END_PROTECTED
