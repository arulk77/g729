`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
FeodjPb8q1Je1RN7ZnRnf6ucxFn31j0+Pf+QZgfpPZW2pT+nLLLUM9TMD/ml4a2r
AIJxz0KouUsPcocUonQZCl73t21pXUXgbuQkB7BhkNerfvhoOK77neiyiMyZd7ZG
k/haCetCOi5uxbqx6DqQlXBV9Ehu/cXWbsekaMMJl+vMfUYaWFuENfIbQNY+7ho2
mSM7uJfybPUawYxyUz7t5xEL+6OzdhrLfzEIKCG8BO48UFJFpReIiEr7hX8WsACm
9WdosiP8QvJ3NHgDPwDoyL1QbMiUEKo9oJgMXcn0Md9r7dkN/BuyaAOWnRL1yNnl
3VK7q6nPioGGT8+bbAzjOd2Bpvwh3ZKrTD/KK6HOg+fYJpYiWm2hm1IbN6Oc+JKs
QGzMPrtI9fRQHDpOJSQvnduf2o3JMgRJNBwG//Z1jHoedMCn9CvQeSbHQ0WiYFFn
xVuBsFjnhQoO6Nxc3RPZOxN511yZlZKN8wMOVf91Bfi1AFevryxSYOM5OkQrkjxb
hNvlgG5lxCrOChhZHZDGtIPSLp3Th72I8+Xd7dbg30kUxeNwc8ytLXs8J8WSbzeP
TdKT4bzaRa1A2oPMTEURHgAKws0Bbe9gZTBRuGxOVdVY68s1htXj/5Odxqzdvovv
n8z3Uvi2StpQPzhRlvUsG43nVmwT3MLWj2LRKyIE3NASokA1LqPLHRWMlbvYbEez
fYbwtmpdK19q+/OoYgsDJlBzDYWll6lsx1y/EsTk6o/zgwTeyrQWDkrjnrSc97j0
1giQa8OFdajgXQzTk++R40f/74+LfRo+dVVr69P2DLpmeEFFv9ClQaz3VP1vzmuX
ebGZKhHd3figj43zSKWM2culSWzCtYoeNSSo5GuQE5qzjBmWSSLwyUJkznFLv9NN
2sN3CR/04vFTTwgVJXxzUeNwMgn4jWCy66fdWEZlTAMQ8N3Tbq0f9r82mVljCdJn
CyKsyCyF6vtkQSZ8115S5zFcLZwD+g5thMOsmHysY3IfM/5lr2e17+PE7AMrGMcQ
lGST3Qe8jl+cNN+klEEtsjL264KsyX+2RPRs84zy/FMDabf8XdR6/1i5WqKSq1fr
x3174F3xWL8Q5dcFM4lZjBbV36lj5KjLg8ntudZNv/mOhv0jxToTzFKedkrGHaUe
ZGmW6/eyncg061tAlyoixA6W90rsCNVYEH+JTlAFbl3SAnz0Q1mHikz054g4p++J
ceosTtFNCZ5L6TuOouPnHZYFEOQmwak5ponVlnMY/2mfDm7ZJoYuPec7pJtYZumv
QdooRKaqyWW0o6td/NCPHruRqXZS9v2u4TgzdzaHxs0BhF9Kri5fNUWIOwupxsfl
V1uelVW5ztQrGYCeSJm17TcdmRufzegvRmce0Eed4gCDqzv4h2r3x786QpBnxWOc
sbCTF669RKHGiP8UyU9WNehFzmcwhHaTSVF3bA+UOwVPzH3Oq+Olyb3iBOBnegk4
C7aBR6Zc9zRfTqMYOU/ySYZxDePRAjsJJCiLAPU4dMvtHQbQJ10ngrykOHyAmhCN
p0Tcah1cTGj+1exz+kXw18AxmjV48XbXyltEqJAlyyHAyCTP1v/vLuftn/CaLc7L
bx+P6nhvycBVLHXyYBk+LINPorMFJXx1rDuTqjf6Y6XEstJ7w49AMEeHM7uZMSuL
nsDlQjLatFt2hF7/MZuMv/H45MBYjo5rj13+S7rkyehRnnD8xRNSzDDaBEsNA5bK
UUWZsercyG1HTcBEPQ5Nym5DlKoyR9nVIPJHbmU6f+87mmcVL2TUufmt1KuEk/sh
KFhcs31bpG0SyaWLJCOfI+oAdhQB+HLLV1i7yMRgm++DPUOJyzu6z9crHuSPiuxl
AMlhqKde8dSLC4fYqenl6ZtawypdBprgwYcv7G6M8IAZ44Ossm93JS8t+pd/LD6m
`protect END_PROTECTED
