`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42dMjsi3gEADKrwQ3qgSD5FsQBqAHvKFSBlZQvy+Pe8E
h81YjxZBxvwNALYA/a3vLjVM1DktCLQSUMbPa4nkqzam7f71ndnnldUGmzFJ0UBX
1l/3+okp5dxahJDYKwWcJtHhpIRW/fIR2bIsvbhdYEPfljDUMh9EN3m6Kjpt20JC
nNhRa4UMUTZ2pg7TxoK6YvYci8Jx0SUeMM+z52c8X5NhPxbRwntnzcWliOcxPTMb
y0mX6YvTCWAbGhSOdIGs8hHC/3cb1IqV6OjMqJyG5I0=
`protect END_PROTECTED
