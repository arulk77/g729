`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
NbrrI5NjmZsh8bPmF42w9EvV7TlCY6OqifAUE36Jv0pbnS4Wv/rvKUEAOLZuUYTH
Z6mOlLrp1WiJSNvIUmuqnTeMvpu6/r8X4JqD0dbgilLWf2wLZRQ86ASrbubCv3xj
HKI+kslOMNNCtlx6aF3TKIDXhYNbhmq87i13I86KS8zMuL+b3NrxX6UC7vYvAMsz
g7W6z94ON2bqmQ/+yR3jhX+B4cZAz6oVdy/5mB1LwoVB3SHnLcfn5nROe0t1mwx4
LnyeE/0qqEBoZre8J4OHJgdwH41PiasrOfgUBFDl45o=
`protect END_PROTECTED
