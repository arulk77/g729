`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4yDsartayYGt6r1wvVec646R/yVIFIJNi+NG4Ukq9ZW2Frti6h75JhXtdAXGytf0
GU+821y9zLCrbeilEBHI39DE6F0bXX0e+ittVkyL92p7apd5rWN0/QEzGrz/6B4P
LfXvzNbJN6AEXbOKhFOxTS6UR69DoZrMU5UIN8EQk5oRtdMLKN+YK/WZ2Pp50SLz
jdBy8fz0Rjo5662nE18JnhFCwpO9BBvzgDkSCCWyuVr3vj4weXJ2mbNBhiDyLJrr
N5BeS/PxxyUbqR6/XwhqP3VW1FIS9r2E3d7NM9MSG4uFTvqVIxlncvONA6PgysmF
8KlpHB8LR47CaBr1arJJQSVT+nwpaY8T2wzIFKlMumUPuXrX+mMHXC4fDZhE3qlK
EA0i65K8UgBuhjtnxR/PapoNvCQJVHZbzxD1So6uITzi6gngTV8XJSGuJaEHERdW
5M56FyCL5jP4H6iErmRl1nocHZwmWIp4UVs1Bs3vmWiI4gGzV8JZpNo2hFFH4ilq
FA0w3WH8Ng4EjyF3Ly7ZgZffW8gQ0TXWLr4C4k4x6hp28pIwcrimSvDirvEB1frJ
34CzYnr85xpztCwHCFfsmg==
`protect END_PROTECTED
