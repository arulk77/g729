`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QNsPahXRFAKX1XBsryS+TbuTk8dwzWyucPB+iYc34to/DjPUWT8gTKOxFf9J+Pzy
FN3ubsAE1pH0CZpwkMrlyskDs8E/oIAgMseKojLeHtmnFIvilwclz/VK3lx2LFjL
Yo/uOlll4/2JlmlIUR2fgzP5uc0DwNIfc2XXpx4KWFeCztDHqi793iJxl414hIlc
6RbYQEetqzuJLJr622ESg7hwovWLoIPNPVkI+/OYF2CvbiydlN/T8OvT2BjEp2n8
pKgPh+rB3OQjlnRImLgEXKHfP7PDlbWXmj3XhgO2pBuz2kHqLR2Mb38I6ZwPTKC4
l9i8m8DIcpdck/6SqQvSwgXHdkQdy5OGqAG7odPpdJ8=
`protect END_PROTECTED
