`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePY01cO5kUR1tztY/toxTk3DxSw//HyMTm49e2J5wfMo
apb6wbN9yeEQ6QAW4IStatUq+0d2DCGA7V90f0ieQ/MQdO0R62sFCl2Wq8Embrl9
vx4RG0C5U8eH+dgClnejTiUEs4jMTM0/Awu5e5TXwPg9yJUheBEF6iCDbTowYeeP
IvY6XZWncRrxgtazMHB9SNzZ5i8rfqW+XnpL+2zyFILZlt09bK3qQAYoituphaQ8
52V12Ur0eL2kD8uhYBay5k0Rh08AyewwvHUFqCcC9Fq02Ez8FDKIUgCkRSxy/J4r
F038NvfK3MdBD731O4gEyA==
`protect END_PROTECTED
