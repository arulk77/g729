`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHZKPcAs/Y1k3sOEFk4m2Gnd+4rLFwiIc4rujdkd2Sdi
kkD3epbzNfrtaQZTtLf8WUrhK8waniey9YB8kyq/BW94yFqaLe9UvKUzn+TGyRZY
qgQVTzIPDbTA01mYkxhg/rEkVsmL9I1m1Z6NFEYnplotgbEJqngLh5Zd0XUS+20v
OmKnUul8axdBhRtefo8dNdrc3+9mNgb2WEm1VO9ho7MWSrQrc34anfo958rlG2Tz
7DtWow2sfzOJnoukw8oxvWUFLfcsh59DuIGfE89+UfbbyniY+2XxdsQqrip+0e2a
hjl705N0w8KgQFzmLyYLEMn2iT8iy5nBLq5QMxKUS9uxzstkylKIbiq7dzdttu+J
rCT/oND4PkykEjBCzzvdQA==
`protect END_PROTECTED
