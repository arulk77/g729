`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBUbAZ2Wit4JYVZG2nWJigqlThrwiFa/y8j1K7YYzej/
akvEOasTrOTGjDTXCnggMTBLEtemZ3bbItWnVt7ajvndhTst+zGkldiMhr6f31zJ
wliwL9MLaSN6atJGnqn+dt2ZoCiEigm+ClZEM9zqZ6E+hHDqZiLqd3GfTJBC3zfn
XKICWdi5rn92wpEtDQp3O+iFzjab/hYpUmccrvUrGuEtZ1lhYXY3zoT8H3VC68OE
ZvbQgU6afswbgULlbCMoxWl5+Unyb6Zpi55gMMa+djj8TQ1t+6j1JYMr67XBRGbF
0Z3x+eBGplx9WXgnIeVkWGdrkGo6FxojucyCYrycYlvmuVeQd1B4cxDxFU+JsA66
pnQJrUu7YtRStJjgfbFk4py/ZvD7sIU/s4R646YnDh/wimMnuLrhi+hdVHTGE5dG
gaPGwKOeTTtJohFkRTU9XVrCZ5ap5aPxF38jzo5PLZc=
`protect END_PROTECTED
