`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHhjPTmugqTpdFUHiVxsx7x4LTUovBGxVIM91pPVDvkb
qPALCxVDHDxuD2o/kdkgCpDneFNx6eT+ITgxwx4KSexHkiMiIn6RUPzuWg6Mvu90
5vHvWJOfIRcby3QHQhjGTCGLaHYUdR/HHYyLVkmCKBcsllonr41xpYJrKb2mnAHE
I/qbvPSqzDADOayWhDGUXjqAnorf7J9Mq4aLolYMOEYKVA/jchv2huzulhrYJ4uY
yJTGI9U4t14fL0mUSPUn9OFp5yV0LQ7UHIfX05UeJfIM7i7wQYyFEwA1CMn6UxLo
4JrCZlYvDQaZ1OiPgmEnTz0WRXUVue9OVfm8MyDKVe+jSdAySKiIVl1KFh8VfanE
3Ls9kku/Iaj4TQkctD4Ob4JjGXClQwvHdpE/W++RhAcNpJPjlNxr9/XG9Rr+pIbO
cI3uTc/iSrS+z+0n7YOKAfJisJhwCvH6esJkp0AZMmJEJQYqTo6kWxaifkjp+/FM
d1cjG8ON6J14IOICincxyuo1wyDxCrxVAKi7QSbZS3TFANvf1UtdV6v9yZ/ol0V7
`protect END_PROTECTED
