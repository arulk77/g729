`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zxUmxZ97ggZxwuicrtW15dY90e0p79H4DRRR5Gflzrs
17S4yMJybFwvwIs1HZvsZoelJJ3205jnYJAxYXBpM0pkgZveIQPPqVdbpGw0mknu
yxmH+yhco9coCyKkIMgcNfdJAylRwV8LmFTByJ4GkhV7LJT8DTSTdfFCTktScfDF
iKJZULfa2l4HR8JK3Qkqw3s1M8kv9tZRuU/7rmVgmuJaNC27Byj75sslJy4vkZzm
WsxBPPzZalpeSjrIEyfqNNoXLBIW4ZyiHc2fHpLfxMw3OwBOCV9EgR1Z2i+7FSRm
z7K/WesM8CXIykJC7Sdb3vgx3JKRkViMyEqIHCrly7Xf+TR99XFQ9m6FUrP1FNXJ
27t4C8htiQK84S6h3MZmgg==
`protect END_PROTECTED
