`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2UytfxBgO+vVPYweFSR9AG5JFf136hs6uivZpYjF2exg5cdcOdGUSpCfDx33H8gx
0cD+6WDJK/Wt92qA9ES+PxGUBusdoblLNIPmVL0EmsC6mXejIi7BTWxoOiKjdxv0
reeBUgZCOiW2yHwh6KCTaAMUkheO9TxJ2QDe+GPj9uDU3jzthhwE7CyCSCdahOBp
06rPERulRiRS7VKLOYxMZq4HomICnYaXzkYsng2I7FrQdPn2KkXCam+Z/+Ayq5Lb
5QwkD1AwFlgNQxcjjEpKNk0Byn7NKSUgMpciGu9N+e0=
`protect END_PROTECTED
