`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIjrZd3JlG0dMiGoCOd3JV6UB0QpnCOblncVnkdnO0yu
CCcJ/5yy/krWIPqTglToYhMmWi1b8OaZb8Jj0aygMO9wR4uI10yvZ46eKcYqtxjv
GDRl/isdCmt+Rg7yD+vXMq+WbMYzyvWIrgfkNsNgF45B6RgTrmgVSJyg9lST/IrH
RwUQXzcT0ymBUzQZetxt8NJtFSQWSogR/vdb/GF/VvGSPuqz6pq8eN+0F3P5xIml
O6jBp2ovlO3rYRmvElrxEYwy+PjB+1N1nb9gNGixRSuxUu/fjRHUgg22cj/DKHXP
6hUQDqWhBVv3MYYqc1eYj3n45/qM3h9yPzu4cuoWTkDZhyTGsLIiz/khG4gLruzi
kweuUL6H+vFdOQdFk1cZuDGmbbEiezq1j3A8FEJfg4JzLUqhpIJbfCE5/QStKp4p
uIyUFQOMftycmMZOqaiSY/+9Oj1V7nUEUuJUHPcEEfzDStepcSASJspymkmWv13V
`protect END_PROTECTED
