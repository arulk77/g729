`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4z3VuFlywRmt0qaprVWIhnTekU6kfKvMaP6To3RIrPpx
zOtCCv9X1J9vgYmS7dC8JaHvdONsOZVsr1OdYLkdo9DhiUR3rtCCalU44wrJ+ktC
G99RMa/YiltSfP2DMs5/XQJ/5Lx5MANdGKKhIH57X/7FHFeBCZt5uiwpp9NZvtp6
ONU+3TR8MAOwlPQapzqc725+FAsCVnc6yoAtaKXHkUk5ElujCuwV0WKOw+wzQBBb
q9KEIQIeVAjQTGWkrnCGCKJyw7kQFuK76726yOAk9og=
`protect END_PROTECTED
