`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
WhoQgZpoQIasuZDztIsmKuCjCrckL3kFp/lcXHcXA+qpEMUs3PWI8KGS4KnKJShM
1gClkkkiGVCSmLTtqSQGsQrZ2141QiAfRGRPDSraHjINHqfbHPXtYVdOGTRt3w9a
jrdE5F8JQqiBEcptBkMLbuW4n9Em8F37/MJpgz0GWtqgK0GPjrXvbgEhUeHdrhSr
yADk3gfGBJwYHDxVDFcgX7wj/ZuarhJwI5NBvjjI1Ly5F5AamO7eFh7QGIJp00Wg
EMJztsWRR7sPN2ZWTsr/11IVObiiSsLXAPIetdz0hU00XEutb0sfPvvYDCuel71O
3pRknDyw5PeueXE055JcixfylH2FgE7KagExFlCCrnMQTVcOBZioy1jP9PPTj3cL
uISxEoz9xPqzHE0L2T5L/H13j8M+gaQD3bRRV3wp/NdIyKnmOHB94qI2Fd6uiOUk
XiQPnGMjVTsWZqMLjWF0fP7oCWyAbnv7Fd04MyRYR5bk00ezr2m7hq/QEAz3GZwP
XvW1IYUYW25gieGExFEJXg==
`protect END_PROTECTED
