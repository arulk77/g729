`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
avdSWSrKIzQSsX+7ITa+SYQnruo3OixA3q1+QAnqLix4sTf2O94u/c94eRexd+qC
63acx/wTAfmpYB7IMMbidhMPwxvPOWqSO8Co/MSaVw1h85YMTiLbKZt5qhjJLKMU
emELCWkIvXesG+XP3y9UXoLf1IAGo8v7suZ7AmbGsMVjhchnvKHpuH76vL3PH4i6
QfLpUTlQQeQo2of/pGrgNNAKzWl7Xa7wMqDtBsKtgcKmGhCjmYLoXELWaJSA6Kga
H67NLM3G5/dwgVnjd3DeqsykUjyqzVmrYwHxqanyHZaFvDlTe1PMLnwjL7JB3qUo
MwaODtkXvjMEOhU8OC/5Bi8sgbQqMgIxb7UfmZGPfACF0uKCvObpxU/TpjghLTYd
ltix8zIXQ2gLserXi9zWQvLrhgqfHjYCGM2C2jERZB+OSJLY7dwpK100tTo76h9+
SWFnKww61nsfgyfsRpnX2G93yhq7Wo0ei/2QCZYAxNMVk+2rSL6XZq84JgJ4UJhl
+92hQMLYRXFS5+hr9lwBRhHpJ7oObZPqkoyjoe1bHoKKpdk+0M5wHj9jEXJvV2aq
JKOQrJAow2Oza5BLYk8YCtWMBI8cpoeKCGSVABcXvXR6L8O8P8ndCPsnKnz/GANQ
L2onoTmrT7QMuIQ5W1hDCvMWGmZpsT9DWEg/ZNb6hOBaga3GidBwcqJdwj1xeQn0
jexpoU6zaL/zTcqxVwSfuh7+AnUtYysWKcmQ4G//lsd8bWbIHxSgwyl6S7mCoxex
ghGvQTwnmsl+hV+BggFtlPBsT/9U64Nxb9QzuMvtJklSO1q7qwxdB3+FxgztOKgg
J2Oaw438XpFGyYfHNlN6y4Y9Y5SUar80kpykJ3WGKYED9VCFqIMlDP0PIld16M9l
WFv7UPRUGqTI8Rg0o8glPoVIMI9GFlQIrYutqQnqvbafc2rG5Es5wuJ+WyVH/oTE
9giCj+xGmFPsXfJNwYeSCcnmNK3meVUMm+V6eVmqOoFTc37+/lvbzTNNLnzhDkEE
Gya4Uxs+Bi4rbI2JnfIJXZrhgyMIbxUaZRD2f9tEVe0AzW+WQyVOF1Z93C+EMPg6
/G9wjL9xvuTzwTsyCQKdN0M+IzN3sHdZhcNz/2QcxSrY3PU/0H8PTwDnF6NDhgGT
+YTwgQ3IvUfV4RuEp6Uw6Kb03x1uKTL8w9FbBrGmOyUmO+S+jkKRiHXzxfSXD42v
Y9NLETKW29QgO9TmzogqTFUlR5ZCIZofgo9eMFv8u+NkiJjFIz6n2ghCtfRBlynf
TD2XMmIEkK5y6CkWoJRJ7g+5NJphGbyxi7H0mSb5BHDlBdKQjOK1dg5tFxlQ1E85
rDzFw4KeG1ksvWD8+RVdoOu6PIxqffZI8SV7tuIzB6t09VdkmHGS+5FbbKQy1Gmm
coBbtKg5GdSKJ29VGPEEmA7tlCrtfi/CaUVU5TzilTotZdrQLIKeZtJu1dKl3un0
rOmusj31Gu1qrvhk89YpAzc+DsOwV8ew72WFoeTFkmcWOIGcECCIJ7lUHUjs2VwL
XnvpEjWHIvbI27YURiiZJYLTAu0aECOyUVwG5h+goRci/JEhf+qKIjbMbvKtq0x/
3h/QBX5zzuH77ePCBkcozqpLtxAH7L/NFnWF4HLzs97uuNlLbnnS9RieeibDO4Gu
JS22bfMnETgxhlVF0YRE6mpO/8cKLluxnimD72hNc6ZsXX6K1ptTi3pQFM38VLKA
6ybX9N378YrXr82G0t79XD819Qc1AGNGCglcCirlJvvezSOBVc1iMTY5sJm928iW
`protect END_PROTECTED
