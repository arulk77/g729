`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zZrh3+NrjQ5nxOnC6T9c+/7cTWDwdHdd16+Af2xKsZy
OVwwMm1AiS8L0dpHfZIW66oJtg5DbXTiGCrPVzBN510laX3RI0eDIfP1Vutz3WDD
O0ynlgiSjFpF0L7WWbg8duFX3QEaQ0r7C/SNjVRx6yxXN2YepAeQ3ILNwCyW25/L
NCQDrbig0Np1C635Ij+JISs7bw1z1renntpDAHJwtpOHKX1Cyd8ysrDLbJUV4eEz
5s8rotuQIXnYjBDGuFccRtZMoPvXVhCYj91W5usx26lTtOeUjhd4+tyByGL8wM5i
czDEl6J0652OZUrE5TY0aSi0fj5cjXu+HhwSTY65qHHCjROv/qn8N6HVoaV31NQG
3Yo5Jty+kSFwUoJqgtVLJg==
`protect END_PROTECTED
