`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDj+t/4mhrS+h5KUz7iR6hKM8BYhLUhIpOqCTqq8KYaS
JqSUGZ/sIgXZbjvl+HSYUrzMGwUe0HxocTrJz57e9rCsGfQPUFT+YHMgWjCcDEmv
dsBkHTCpjhhuMT+/nWil4UDpkEGrZfsL84Ug48m7qr/wCgKN7XU0NnLurCQOjIUl
HOnRenoK3RIKZqbLywTlaSTB2g+eCdUGw361JGXIjZm7eBZtayzUw8MyAdRRz8Ls
A1uyzNpKyrzYkC7LfxygfwhNyV584KW6dkv6j4n8FJjufVu4b7hUEpVOHceS47fZ
HZIGjThAkPNvozJpRKOQKwvEqvcD2od+Gxq2Ff4QhDPKoUr2ca5IK9SW4ZnyNWe/
EE9TBn+YEZeDR5aUpqK1g5PmnpWBa8nz26Ph50p7anySqwJpNNaklrO/bZk9s96h
SFmyWUSF+ySKusYRucIzcIXdRFGPqU9jMy3uj46J1vXVznX8hSnZw+N9wemlKaVM
cgh9LOLKfeqrJwrDLrZlB2Dg+DFAQUj+uHqK5X+IpZhdOzXgyslioG5ktkfE0pJl
6kY7EEO4MZFJTU/8TAvoSgAY5PMgAFNAJhX545m6fwsQtLGWOYJocQ3vwWKN0Z3Y
/3Z1UNK+1kCxx+mQFy26/Q8hWt0inyNZ5MbkQEPUwcF0UsFt80Xn+6lrF8U/QU8P
`protect END_PROTECTED
