`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePVebJ5mmnurtXlxIadlojjec3FyQWRsX3ratMp+nU21
wLjJy4h6Y0ZYUvA2EnIc/+WJd7PzLTTDyGz2wxkU27p5dSq3k5nkAbD+ZTmxLrXU
fD/08K4hoh7zZq1uPeypYKmGda81KLk43MjPe//NBL23Au8nG7yzQQZ14lnA/3+G
DDIAC4M2P7BUwgKCQSiM1tIDjJjWseB3mKYbBU2IwAK9JfZpfoLJ63tIqm5rh4yt
uXhU7tPFyPppbejh1P/Rsw==
`protect END_PROTECTED
