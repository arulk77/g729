`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wBLSjbfoUi87/GTtUbXYdHwmNBZbUd3XHhhtQfRwsJc
v2Zwm3AWprJsVPaWiu4Ay/kBWDOJCKW+pogAfegwsLj6lzQcuYDV6gvfXnvNcJkD
mPTkL3ERW4vIye+BK82cyW5403PsLDSQLC0QaHOKbA/PqraMZH7mH0EyekRp/ik3
JNLF+NcWSMxoCdfkyKzFUorWylsfcuUm2uCVzcg+uG0=
`protect END_PROTECTED
