`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
zs3hFOk0Qg+QQ+T4842qtajNPut67tRzfMLC7fTwx1ymuRTDy4Tu9XXEqVIW+dEk
svxspqcOJkAPQ8Gi0XJ5R7UC0OpHBJRyhuhTRECllJOE9Yoh47spcMY6X/hb58Xl
wzXHO1OUNT4mknGdt/53JgOUVWoNw/PQyyt9aCUsia0rqb9z4OohL4bOFNl0K7t1
bAMPcnB0fxtD9U4pItJPGFvibFDLKmCFSiHjxEBhtdjetYhcqANNCO9mWYpd5/tS
llSGnu97Fu6BvvY7raDnR/VGzlYGwe+mWzLpf8tnbkuCONjoS4dNbgiNcJM+OWj9
XVqA4B8d746Td9VkA6FQeEuvhA9SpCFHMjE43qYA8zw=
`protect END_PROTECTED
