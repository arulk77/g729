`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFJEfCUYHlRqzKpxzZtrXIzp9YyE7ijlHy2GqgiWqyQ1
nDU730nddxtkfFM9qi7dYTMuUyghADngT8KO62W3pRXM4jJRV7i9+rDkUji90OJn
5r+C1nz4/u50WmRIB5mG8DaL+QaYaScNSga6DePYy0zXxKzXYsSC5OcnhV653hCW
2gVs36lIDgrxwOMSt8YMshaIAfNYeMMlHOPn92Krb2K7RWzB8TAqqUepRKoSRakE
hoT7YZMGiwXCe0O3HlpVB5d/VLm1PIllpR2tJGyjAqMSPE7Dk7Qix1b32nhkbOT1
Cx9SoG4/q+TPG+tqW7UCug==
`protect END_PROTECTED
