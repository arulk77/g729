`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB1SLIMjjDioGP0XFKkp2Mm/KYPvJdFG+Epm0nRHl4s9
BcQKtV5cIFLtW32obOyO77F/hz+YVxevH6/B4mg4XpinBYNY6mjlfs1ux3vGeHC0
Zz0duGLOV5HPQB6RpOkqsfZE+OvOMYoTUXfnDaO7dZWfS2xF1U4ztiBh/o/fl8bp
wzQjc0cL2VgghmO8DGvCUcQQXm2kXGbulXfLzIacalOT70UqwRdjaHT6n0xPxwsh
kKktbZ4OMJTuz1qE0Y/hQv1qpNeRL7hdRoZ8AAZ9nYqw8/J0e43B/IvQd47X76i0
yVnD3PGklymYGwPrtDeVcEYQYXsfG7501a6dxstSbuYScreuqZ0wcVZ1mLHIDCBl
4bbUHx6gDOL0NxtenuwoY4RwAaEcR6knlRElH2oDiYebBMk384baHgTpFmBuoqK6
t7hE9frr3kCZ1/SHv150MQX5n7JjlDgxtM9fzNr/oeJswGUq6mZxuXtHrEI7TDtx
uBWayIcjBXOpd4dSirXdsz3C0nbR6yCxDo0bsb+Oe3pzQsmM6KpbqsmbplqoXwWP
MxGBoXOZoFUTsMsKyiPRS7+Nx4ZVGasWA8tVDzKht6HYVeOjytSPoK0OwNexeowK
EJwSvSGEILvaQBrvaUQVlfFWuADjfNmyGJagJOYPggahWUjAXN4pGqEZdjijKML/
QGa0mFHocHSoxVLlLXpHzfY79fWDhCS4DQfRBrNyQhUk5xKVk9ENSiLpxdQ89D4F
q2b9rB/KwQXotCjL+DuqZ3cQufmf/0qJjK34o+eZ7bfxCCsfA+EmC+z1dpxOMZYi
/DITTufAdpGjSb1F7HWoNdRTKqSpx7EZmMYsuRa005DM4+M/8rRWHlhna49WRdz+
fWBiQOBXojuJprldeg4bSQ+aQsnZ5oicJ7NkUwG6ij4IzIejHYDc2gC8F5hfzRZ6
bJst4oZdA7NUIb7LXglW9degdlEr1xA/qGhTPgoyzK/uvwbZb7Q+YMWJWQ8nW/mI
sHS+4lzYZvGXmvY9fWnwxX3Lvar4J7X7TAhsxdIAVjdDHwnX6vzuDEKTElKTcOxA
/efhdQR8/uVVr8ZS1cFVkk+cMGRWlDRWps0t0vgyBik=
`protect END_PROTECTED
