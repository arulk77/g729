`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOm5ZhWUEj/KtPyLGwLQhGcW42vjQBIdaqSONyCqANPD
g2sTgwOyNQAX9lzw6RHsAiNBCXqwBpAAf5LO96PpVdU4T4S7wuYHjHiRa2LRAupL
CGu65xS0dGI3KSU9Uh4wcbKm4h4bLApXKcpUJYPTsY+bDgJQDDcLxF36H0Ix71ii
NrCYopyWacHX/blXmxBxwA==
`protect END_PROTECTED
