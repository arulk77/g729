`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAp+LAIilR1HyIAETzUO/UUj1GIVRwm9rjHvrboZT9W9
OiWN56OwxTq/k+wUkQoIQCt3sOMED86rzSANma5LKQ4aeWcBGfZk0y2Kqd905G5n
yAOG1W+KyyzV0/WDCwV3/xVb2angWWQlIodBCvnm/kx+MoDNgcSPtQmTYP+/TI1Y
CFV+2DtnoKA0zOKLdv4cffGrgQJRGui0ikuubaWBS1rm6iGDxbS+S6c7+tQGXjoj
/1N80pZypXRIasz/PHVG7w==
`protect END_PROTECTED
