`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJWOQrM2q0ctl/LOjnn2WAd13LMq5LZwwTbDxa3TqW2p
CxiIrkpwzaHfyZ79NiraEhVjKgJ8AscAmIFuB5jat2QimSYjb2KhH5xf5B7ugIq+
j6/KimF2J4tW6PhIFZAGxR1ayS8AyKFpuRJQEkvtaz7eXGvhmnT4oQrt7XEVxgzI
YrwnYWnfhCy65bneK0kDgHu0Mg4Nsaq09Di2KPMY+6ypL6uAEZJAcU6BPCt1L6d8
`protect END_PROTECTED
