`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP0XcmlShS17ggpdBxmyntqm7+ByNxusX0eC1er+0Yc4
onFmJqWvFW44Et0i0xCrwM+LpZzOBHCzLFFN9+qMRBpHyYqhbJpRLufmu8xTlYGv
C+BXGawyoA+/CYn8sbEivr/ZstTa2ovTxu5lWtHGwdMXuNpQP9I/Hi1XXbnlqF6c
OlsJFSjuc6PWKQl0onkX8otWiRbsrWaevNGHVtnNOm6GbE2OfOvOIJtaoSAg49N6
DSIWegsU3cZg4tGuYgL9Atiuw9/EFqF4iAJYo0/cYb9T9qfpcSBTn8+xIR1NiJ/G
qsoYcAagbsu+NFK3jXV9/g+VIvUKbjvQBZzAjSaVivPwyTuWBhmz4mtklvB1Mp64
`protect END_PROTECTED
