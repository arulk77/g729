`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHKDuVIYpIBGut6/icm4TGF1JSbZ1MAREUpBGW9+wO9L
Eyu2PkljYIlBOtW/zfCTpZtZp3LbnX8GIWKL7+IM5lBYm2Gs1qaDxMymtjnfT5qL
SSb9NKDgWLBbxwH9QJee1FSTN5EObseN9Yp/SNav5hQU0b3JbIfnKkOtOjMpjTqw
IOSMSJSsaWbxDpUvyr1zLulRp8UB2A5VsTdVfIvcs0c6Gua/jdtmFy0jYs+Lz7+1
`protect END_PROTECTED
