`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4ywekIi+Vg143q11KTOKRMcLnw76NBTO3UNfJO+0smUW
owHlalKHpjBPF7tSJw+iWyOtWjTu9pqLt1ntNMDLttyrJh4VjHdtkU55QkWODznG
RYD8FBM59bq+SVMjWiUVGDi88+QweUW3KeHfjX98ZlI0Qc97t+HJqpfxYuRP/Anc
hj7CFsLBhKyB35146bvhweChFlnXjpfXM8A0sHGbxcFurk3D+PyFywOe5HAZbcB/
xXRfFPVvBt7MFLX12SvWOdNaohhhactNJ4vHphb/kmndT9uO950hFQaqjyD1OhoQ
cB9K7w7D/lDZv+XKeI5b8GYZOwDdKa26006yd3sioQauD+Vip3JPIssCe5/F+czL
XnepktaBaG7dUGH2nG9tGQ==
`protect END_PROTECTED
