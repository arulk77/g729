`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOuvxwkz52RZlZgaDq0OSv47iGnhsft9kX1PuI8irppO
kxDx7pFlwX9MM3qxAAD6+nUZp2XJcbeg5XDmOkFDfzAp9KA0NgeBB/1OKfEI7lqK
YlgPRPXNxoXuRLkH2zJ3UxW7xzHM+OLkk+DgyYVak/b3r+DW9RezXRzXrIQXMsgV
a2YIrk63NnWfaen+EWFbuY/SssC4qRcP7G2zHDvRKse0qssMwV2IGpDchMVIgaZb
ElJ1HBDxRYl8/fRXK4Tyw4yeiD4CFycrDUD6eOvZEpLP8O2nUoM1aixOxWaW13Uf
z937U6l+V8f23eyqVGmco+5URihO5X6uTvc+G8miTyPkkFOPgIoIfXwGgbhtFEvZ
S42GqciFfteZcIb+2/4zxvtFUklH5bDuSM9Wp3FyGcItJkAL/rPBX9bets4aB7vE
3X9+NyL+Y14elYBfPK6TK80k+0PTv+H+ORE8T0KX34gJ1xDEDt+UlKrzhrT8/n4x
A3MrsvMEjmSzxrE5P0d2W6Z4gXzclFKqgoA4OS2OBhl6y/GDWQAQNmj0gtmlQ3tw
eH2C/kpY/C1Eo6cu2Q8K3QeGenM7vqtskQRIXVPPQTEMYbOxqmuLywvrTFNHBgLG
pOw0RLwbO3/xhmRi+DHWtWbJnduuqc7wcCtt80OJTRrku+2+0EouHI0DxQXb1CwH
EVNSVGnqPGePClw+QblNW2wFT3u4b5iWMqh3TkLFHCPXJAyY2gsr7U+lnR1sBvMF
XPhQXaDYajodYCrMB9c/h8qPC88rc8faf3iOlsTJyzxaLRCQepTrYwG419f/oYZV
CjS5EWOvzBz5pb0a+tgiC3dZeX40MpbptaQfC/fuaebssVUgt1ECUtuFj4m/Tsiv
2w9ddKrlIvmVKGJxO5zERpBYlogKsKt6C1U+yq3DJ1+ChFCFtOW6JzNOsNeAlqM5
PKE+dqptA8NU/sD78WwbXGHkDW/edFB/C7/pH3Jk4RQ3VXQi5KzlTScZ2/pvUVkp
FrmYl4UXVacYtmQesJ689Q==
`protect END_PROTECTED
