`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C0pAiQa7AAAVr3ZGcCRbL0Rv5P8HYsqM5CpCiHXrCzFK
8FrmbgTIaNR/AMRLaax0fKNEu5aVOLfbqj9zndhhbCyLx/W96rnl3qDGvVdVgq5o
7A61Gpw32yjys317orN+aS8lYtvmBPneRZt2uAGBGB/XACBN5VrCKWTNVAnukJUG
/85wdZ/Wo92N8odSQ4ENrcm7Yz3PflV1PpEkYAvALj0NHaXDNuu6oOvUuwsjz0KR
8fROqB2fhe2ycXZvnk01VKsK6dZ8+hVUKzeDophf95Bbal0Xu2mfvhpsY0U01DUN
7zrGG5jRVHG0fHOZVHfq7KaAWV0c3/kgBjCXCHn/Mcmq9VCdVpaLMho9aa2XrTx3
LsLxFFcvutmWL/UhlIMuTdUw3Wr2JX/c4eDREswcOu0JmOc8v0yOibqzBHYDg8RS
`protect END_PROTECTED
