`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNyUKohuwP+yg6xHtkRm3GqQ461MxOOXRfFi78elsZP8U
bCwTU9ni7y4ZuvRiZnVPzUXkoEYQNwdhu2JuJDDwIxeNFQAfrTQ9niORc6o5TWHa
568iG/8lTuRjZEIrVT/ADLKzW7mGDVVT9Rv63a2o+E00CdsWUTWDag1Szj7M5L26
bv898VXOJsfMxyRAxcVicj7XmZ+v1kBfyzA0x+/4qTlmsDY0gtiSFEBWpNsPxN53
GfAY2mj5kt8CGX/EeomABuwkXGI3htYCGOorL0j3NWorrHDUU1HWZ4Wlfs7Xm0La
qkNsljuquPg+m8rw6iJW0Nl/Xih4BTE4QT4OrWGx2kXB25TYnQR5iLqBm4taRtu+
2DNGSJlfIUqIMmIwNQfxnLhXsjMqvJqlPVciltRxDK0/y6yb+e0GQeth18Z/Yy+T
VhP+YJp3tZzgfhzHWvaz7iDJMsbfkok1MgQ7mtn1vNmoDS5npMWb5bkuzsLrOdbT
JtJJkIz8l0417UUJmRKE8HKMtaeT4hIIyZqpveQmiwM/7NsR5DoOblwABWr8X+vw
EPqvSr9L2sgKZHY2/QdmayxGDt3wzv6iO8J6q2S3JkGrv5Sa0hFec5drEpvtc7uX
nkCQcMY2XOMc7iNVh6Ej7PUNczwWbuHz3zy971Ps3fR7Aq3tsCEvpoz0uqKROHTi
Vvorb167TaevDbxthRvQ2cOzrmqgZsrUDlj+a3wyDEpLLmTRAX76xQ1yu09kYJHt
wszzuhUatNv50LIigcmUqVzYZyNVNvO9+AXVAecebNO3G+1/r0t1AOEL6nQ0WjiP
95dPdHV1phE0tn0e+VC6/6kJDQ4vZcD2lwNYzTK22uaulwvyXgRQ0i6ezyrOHnUG
K6nbBKFXU5uRHQkQi5upWGF3aLwWqsZnFIfkRb6lltbtHDL6eY+7m5LUmDNrJyrx
H8rQGPVfgYHZlTbJZDEb9Q/Fsz8WErr40jHvFSbFXRJffc8IbSelUPD9AYtBHw9g
pKUz0m3/+0Vk68L5O9d7Es54ku6yRcIBZFO75YczmZC1/Y2oomV/TftK3HrUIh2m
USiKDj8aj8KV0tffkuycSvcYfejEEnLtCGR0CuDX3n1n74v0FqgXWv17apfwEgN4
UB6IZOB/3ih/ckTwqzh1nspAuzsq9iMBQOfSvTeUaTvD8G6wWRdQgbzfCdENK06k
Jp/yW6z/uOp4WY515AsWjQxwCHffw6sELDbV7rQgSp/Hp6u8jR9OSmFDg8CK5f+W
YVlRw4dg0ojyQ5ZOtxrhqp4HZvvWtLg+x7HTS2akVnTb9sxspgoGL98OChlypu+6
Xf6/qPDxVSstPk7Ze2A3xVlAqbk6BX+UHMmVBJFECVPBNdhmvWVZxuNZXd7yMlyI
taVp0yq/DWLicMk7kt2lEUcgMCkRaYf2LJcOoB3MZHBTHSqaGrO2L5+j7a3ty1D6
nzb/S+p41ibEsR170++E8CQgav0KAWoyaAjbjbGO4WpNGVm/8oxPjJ4M5mIAjZqE
dMwbePymdjewfsASQQr08KwaiSkc1obhheGmTpnQgBD1tObe9/7RVRHMf0RVKsMp
wxnDeQqJfW50yjzd2ZOgH57d/uYmCewy2Y2/h8rN1lAxgdQ2hcRU1xYEM6vZRSE6
7o8rf9tfvDJZEFu496mYiAC7LWLQvPSGSzloScwd07JXqiFhEz4ZYU5m3M8QdVqS
/JcKMzp9JYYJrhsmNqW3mAn/AYr0+W5u71cxljP+UAbvFI5hmlhqNe8xNdbqBvrv
7seZAidT5J+uKdgizJsGMh71NI+FIC/KeTHjcCmDZcNO6NG3CN694MlXjNlu+D9I
d/3QTpa3ekeb28OUhLA4xtp5Bq3HaFHwfytpoSWsd40rTbLXeA/mrQk2fs3biPx+
zKCSp7cjgr6mQjZgnGep3fXSvAIW03plo2wN5WR2TswqUEQlC4Hv5YOH9LAWDHe7
yUR91xiqkoujEwJ4d9/I9Nj1Z8ljQDjGfnxhg8kGA0cpozKFgJn1nzqWmDN5t/7J
gttZ17p6D4hnVpDLYtHbFh6nQIczVLhvJLjDET3i7PmDwTvHbG4rdX4G+1C28SK0
1xbqVl2z24KxZaqwJAnEbWX1CGqbpQTqcmwTdEr/rSvE9vYAsOzhzBgC/lJd0a5R
ivpoaMOdEoCKvfMtvLKg/YkHJ00fDnRF2n6TRlcV7sO0yG8hEYs/1ZnQXQK5OyVt
fUN8W1J4biqEoUbKfLibN0ji77aPQAZ+yMD4h9/ohF2Vn/WlLIZknWFDi0UNtbZO
HDJh8Rqtd16RpCT9ncls7329GSHq7TV+kwP/VtIcKlapi1lj5Q4pfQcpyYGdz3GR
XGiUyHsfX/dP4FMot22+yt55YpxaAX+lZQYKRyww2pBr7lOqQEoN/iIsixevZ5xV
Dz0t/QlH2xvPjw5zfTI+bnx8GSRplK0XxxdAZP1VAs436zUmZdsC59s63JdJa3Cd
1x1xbbLAfAVnl6qK6UtThv/KJoL1au3Dgr9EwDHMTx84lZYFkpNF5tUXrm5XcUJQ
ZB58fesPTE2iOcbDaAXkrtOgRsm+UKa7dQZWRgHe0QB/WdxRA3mwNNiq6iHk2tyg
XqYRoBOhnVaePF6NDmxLnanC78jZS7jpKiE3jGKP3eGGtfSScEkQssE1e5uS57YB
LmAnhw5ZLBNnja03yrsm5eV8Fpa6Bt1IxWzjCIjE3PqFRd+wob3/ltaADSK5lFHx
aLUsr2KQxoyt67cdJwngZqxD3ehBn4gCrVbeDamgaUBbsYOkhKw3beiQcbveanOY
oGXKp4zF09Mlkq4tOj0GyTsi2xm6bIAWmkC5DNc8tTvgnb0GqUC1iRw3iyGvQsy+
5uXvVy4poTcLLrGJaddYWSRfE1yac0YPHniXpWh2EXyiZqg/PLMxUwI7ac48xr1N
KI22x9fugJwejNElfbEEVrDJ25dY3kjVmoeYEQnC1X7JSdMN8tzIfjRZNn6Jy3kl
Jfxa8Z8h7HoS63x4NVz6G2kQBLDLI38wMgzt1+EiJUbXmD55u08kZqfSm2s9tQ8o
m3lKS2JfiETAvE4V1vY/o7GEB/OcwGMDSTIg03gFkIMelDM18V6+FVzuw6z9EVqD
uL4f9I5LzBLVUYwb8/54qP3VrfbPy1WyuPfd8vXoi1uvc8yb+s/eazP7cPrRUFml
JUCioJVUi+RjZeq+4EHtI40G5x4vQuSH/Rdt++rsAaVotzXVh5/HZTnNoYczgcnD
jLTEsbCmFLN8QEspTqtRzuiFppLwic60vBlglqISHig3gQ68ovuwG83Ah1E1ICLX
EP64OL3GB20Jp6E11nO8AdvJ4IkZJMPeNJZxOPi4JKbWTg1i0t47OmdUn1PD1roM
j9lhptUazi6njknf7A3MAHNuJgt9PXZNVeXXl+wYfVU5X4MUkrQLoiYNeimAgSlf
5iVjCEyEa5dL3c5Ze5KnHnckX7RJJkde+iitvPTPAvhi+UFolXfDBACznyajdzfV
pisFEJxAh5blJ8C7UsM/dYy3CHX7kB2+0/4MuCxQO7S5yKI2j8d7ZCteXXSpaja3
GOvNP2AAln+c4Dw+C73NvpB5HSyz0D6WeCrmmA5BTEFFTts6QPHxa48D6DmjvCl3
NStiQnbPMzlbExL9KwR44+3wJGReAvLlwsVsABZF6TjBq02QlgWRMUTBcx5NijOU
Q8/6um2jH30aaO/+kzdFOYZOCdwOpvE/LBydFGF3RI4b1xPw5AcPCM7Xfwn1lEyM
EthYfxFDhNCCXKro06k76TAwoGm5W+pFFUfn+zANLyDcwmSl3OmParLcZhelTqiZ
aBTjb6aW1J8U79p4hlUU0VjYcxFW2MqeWgzD88kQigWIhC9Ie6ajFePApzLEZhVP
VyPdACPqFQoCSHL/Ha9YS1mqkC5jDECTb1ca/EARYxTvHJJZmy5L+Rzmawhs+Vf3
jxKB/11xAgibou81ky5J8TF1DLtKMD8Y0SrTfp9/JGhOZJk1nME9b/jRwhz54duV
MMP1s/NSRn9eoHVs5U7csbmvGDWyKsBePXrXpxSFY7icPEZhSDX3eKKYU4LbErKZ
KyFV4UPl5oe9LQPxVytv1hdZd3hepzRI0+dGtWwFelbu8K1WTnN37ykA0kQmYh6y
`protect END_PROTECTED
