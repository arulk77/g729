`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40SKADutt3UIN4OTRW8Q4lKY0bp80MpkoUYM47pObSf7
QcgyASCnduy0VzSYpjLn2IEajNRL4OM3Cxvdn63aj3gKFhx2fb84iPQxe33cnmfK
mUWIk/2F/7yOqO+pp1B4iZ4PkYEMcp7DbcwIhFx8zw3F84/g+bV0KSKP6ufPsajw
6RHjbM7ZadASuIeGhg7xHvY2MO1DUAWzQcyBoFPm0K4Y3eKxuP18b37jIb1SrbHV
RUWwpOSl2cAOW5d5qeXOwnAckPh1Lq3UctKfKyn6AXgavQj7W10ka64uJcz+OrIT
/g7Kp/tho5m5j+z1+LDb+0WfzVuG/RoYTL+Wu9Z4XaUKUfE5wQlnm3LErdU6t3rR
mNdECYepG0kqAdyx1X55+g==
`protect END_PROTECTED
