`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBd/VlVXTKyBEHqM9EqeSt8v6FkLof1/Hp1K0IclbqDh
rwcne/rd5RYxJW7dzOk7RBfELmxTDRBXHaqpTEQw+BP/z/wBmCjOVRjuOsCMzcAs
sEIBKzAx8MhJAWlKruE499bFGdL7MUtwVy+IYG+HctBmBGMgcIDQ4UDKgjB9s9y1
X9MG17VtfTLr0RJx9O8ajdf6a7tOuPVtgv/C+coLvTO5ix2x3vYTaTDoAQHnpAmX
bhZ5ck7fbK0XqlQ7mmYs2L2/NLmahzl12zuXxWLFAbP0Z9/fhiyeBWQ46TWZD9kc
77s1FiYSFQZREWxRmzwNwyVEmDBNHHSJIxRBDqFCfOe2WRuv6zqxU3RARpGsnNd8
zFSj3wuSzO8QzH6ASYx9K176I1jhgOHfn3o+N3icoW2pg7sJ4SiSoBI9nl1q3BN3
rTwAYPlKVMPwEHXpfAikF4Pb3tbbgKyoGr+fIs651+XPbW0NUdtuh06NKsL35skE
O8wQ6Iw8NSv+GDGsQOlNwaaDsx2c37pmLtMrHur493cnSkHIWmDiQfdZ6NZUXbPu
cg6HFHPz5LHoN+dK8uI5KwHAPzUbBsbyXi6CQdn9KD7QCievESMfX9yuCS+yYz4z
GEs3JKesLGd3YeVLijaq1ECCd+qW81m8ONBbAxx5i752saYg54dWgoqIKY7v/vkB
Vcnn+tqeurWOMb1I0PEXtAZ12YUKtwKI6ZZiRY/yVQz38yx6jyp6LejC+jVR87/m
zsewphflV0Lf0hSWGzmeXzZm1Pz6oufKlAHq9w6raq9JOy3bL4Isy/rEz6QUZDqg
PFHTQT+zELIga6ZVANlfW+YlhD1frIV/Hkc59BFVJkM=
`protect END_PROTECTED
