`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIk61rpOzwqSzOnmKST0Xs2qBvhQE8tkClQ6/7wqOUkO
4m0kwxeujqv0bljWKGCs8pwlo6SBvHKTOMgahcuwo5eqSUfSIWGs0abAfxFJE3PM
BQ1dbqM+1RyJwFLx3Ya1MAiJnaduAArFpJWPNmUXSNHSQuJD8R6fYm15RQJcilTB
`protect END_PROTECTED
