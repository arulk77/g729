`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yIG/41JUkRbYytf7/ulpcXuq9xiYxvdLEYiR/InqjTb
+KXyPHP+ykLfzMRcbWbw8OSmOy3VjR/2BiUe3NrpWeNRYWDqskKBR2JZ9mk4hiWD
VM9VmIpSHsMo+MLKjdDXq5SRVmC771E1JTFzAJD+AOGhjYDwXTpSS3VKZXyiIKrU
n1+Ug3un3uqomEbtm/pj2DaQpqNxZPw9bxwd+MAsQ/famXzgpy/Bc87xOqCLG7/5
UGAOdJxyjh0CAoOwe29rINcftJpjfGN2fgbf6cLamDEZTo4A73YNe3AgYZnYsaYA
TlCGc83HVRUosNt0ryjElcXffiTwjqKi/dMepSA3HxMWZ/REqVBmBCmhEsg4XDHu
0C7UNsaeLf1/wc+UY9LC4pvjBlSDVb6eHJHkTM/KjwbEOAB80K2ja1owEgG1mpv9
rRh0zv6iPzO6qg6VKoW8SIYU4tJjLS8iHZhN8oRg7SFB0CTpIHbQyFnUGEeuP8zi
`protect END_PROTECTED
