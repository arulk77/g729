`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aRVV8mb4HTpuhTCVGqGP5VqfomHSOxVOQz9onZuupg9e
cZ0WCw91aWUeH4Vp2u2X/t6anW8e7+FwGvdzsS/ZyZ6QKHh6AzDroY7cT0Poev3r
yw2DQG8wp7iTx6wAC0cJxmWkRlJocsGqqMQodIZ9B06oaWncR529WuG5Ne+S6DXS
sUDENoUZOdwLOJnAqh4bJxN7VknRj3yvDMTPDmZzM4+R9+Y/MH+UA6dpoUiYG0fs
Kb79Lp2rQtA3Z2BfCtsvgnA/fpzsDouwhhKh77fashD/zAeshN8PMGrSq4O50tb2
PgXLNlTBttq7YllpFhcSLaFt5zh/z4s6xlt9ZcmbTzP7X2j6CWhQWgbWL7jpSLu0
6W0vFle+niUKOUVM05Qd/P9mAOqTfiW8dc8c+teaeabq/PZGsGe2Je0agL0Gd6H3
GSGbzJGVwfgpjcRl1yt0smF3cSxW3TnBoSG/xNDI8Q2b9Oc0mmgiRiNygLS3onvx
CwPwKTWzKxUsiuS9WeUR9kZ/vP/1WMk3iqyhSxsT1s/lSStM0oE8+eO3AyKxUMym
Ajec9rWKtuwxQcYrtY4F6VUfmsS4hHcbNIy0gPz7kG8w3kwZv0lmraM1CvHxSayI
l4ZpeoRi+vQJMAnNJceu0w5A1q1mCt4ADR3RAhdswcLLrSblHNjUS++Fe335Tqic
SKs3DzO0+uvYk4E7JgW5ULSiyV7oM/FoDTM644lpE1Vglck98VmfjdzWylvRwb0J
JTj8vcm6LiDr1IqZZZkKUja5Tc0dGv80Gen/OWKBENqB2gZ3aHXHjrSpal/EFsjP
V+t0W7WIvI/E/b5Ln93ImRCLcvKCVU8lp2DYwS5PgK+uPheLrjG9MQsGn0Q9+mFZ
zQEo6ud3szpjMKBzuvjYJg==
`protect END_PROTECTED
