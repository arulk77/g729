`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/JWQ+0d2CUcxHd9Aw7fvqArfaYEqhe9O/zdJrrwJexn
IA4T4ajINxR5Sq3+VT1wO+wKKzCFFZu3Eqc4osnu1trluJBGeMbP8wHDuFSb/F30
Vd/GyO+7ExBLnsWubn9P3/Xl8J/Pi1iX/SjCs9cTasG/b2tPZpQYMG8A8ePgUmyF
0MPTuxZCNhKiicQkqL3aRBciFUVtqVTB7EpkyikWiMVTmB+hSUnJaSi7b38x8u9d
oUJxqA73aUiiLJb7K1JVu1vLmkGvBcTn4NhdoIUALcz8PRePK0LLywpkoi+g3vD7
oTAjcSRB619aRO6+k3tsTUIpKgsgFUL2TrrnUkq9u53QrG74/3zsBO+yeh0Dq84E
42jcZq7/q/SqUUGrqDnAFg==
`protect END_PROTECTED
