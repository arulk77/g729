`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu458El/1xDHBDQnBb2T+KgPecW4+RFDkazxdqu5x74Ks5
0g/P1goL6G7I5+VKzdZPtv9mOPz6x6wrQ/bhoxA/I6YApePQ/SmfbJjyBr8l8jWO
LLM7tSGiN8zcKk7fZRWklnmzwiAWn0rrnnC7cudK+48=
`protect END_PROTECTED
