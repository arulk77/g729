`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
fpoT63MvNicMAFrTT9jSJLbJmmFhzihcZ6K0ELqKERIpHm73+qx5rYw9MyLhqXmC
lU7JJRnftMhGRG7lvCVHQuRGk+acHO3rp1npc61eMiUwuHbo0fkVsskqxFmW1l4V
pCRyL14+9W2mOTJ05pEth4zx4xAQmWZi7Er3uZW08NgJyyae3BsnRgikJjjOIe2d
9k8ayyNJvpUaFkFP1sLO+EdhqEOXPYCCIu4HgtOhZI1Y3EwaqhE+WnWBghOsFgvE
l2fWHWdbu6V+8C0coAC89/ee2ZGISJviORpP+8MuxoXXDa7U66+r4Z8/+QZD2wPm
xT1H1hkhOqgDLPqxxLTbmBgXxNOYk7pVoas69XEKOtaBP4M0zFtv32qtkyM66454
RpS9QqhuZZjPjOqckI1Yr10ICuY9D84Mo7TGQN1gkH+i2naiuNMlUvPiLDE0M/Bb
x0d7DviYk1ci/+vxva3vJFCiidyxJRl8qvTp5cwtBaFtwjFWrbVKrGxiYMFg4Ecc
Vwwi1DWG601sZf06tgFVNsJ/C3W/Ha0Yeo5ndZr+A/gGLT1ZE8iUwbytQhJW30C7
EtxoYE6L0hQafUa0ocGtXTsvQxK3s5paBybSB87i+vG+OxUp6vbGkiOUZ+oQJnaU
XjIYV00vQQ7NFJp8zJI1akVnaCokqdXxKr18x7gPL8mbreGx1NTl/iXQoUK274cR
kwpeWE0rIqAGDQRDHcSacBeg5AmJQVmjsVkmCd10WdOO69XPHwIsR9kgg41b/wpB
p6Mb4UhSIzZPhyvjRP5lUTJsZYY15U9dgV0wtWifaNbZh+o0bc9XB4Oe98PW5j54
2BbZpv5l8UzV2G7NHFOeac52Kbd98og4/aFQCeOK/cwW6OGV8rKbI7WxFIhumui6
BWnNXKhcraZiH4cV7+4Cz4S8wX6LrHBu79lXzpou81utIzBq+8wFunA/HqWvl6Ug
4zE8YESK4VoSz2JecJMFfXPBDlooAfEq+HD7hDK8QYneCU7GIzkF/cfuiXN1pscf
T2lXMDqT1nAxqK38iDUf9vao9zQFSigWBL0snXhVA1rCrc7usIocTwU0qmoNXhhR
YzXd1qu51xbRPLZyyDrwnlU6sxFhA8SqLe1TaPb8LSD2ZdpbuhfaYWZWLBX1DvyJ
Y46IKc1nZdZOO1vd6bgYuES3wDBsRW6VzinFBoReIvtttd575xpua8ElK3U8MYC5
HCI1nCsvXie+KLeNaKE2z3vp5S7mDCivJUK8swjZbvU=
`protect END_PROTECTED
