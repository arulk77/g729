`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGp7dRZrG+p/RopGScK/h/GUDUx6z0ktBJhdQzPajKr/
GsEm09BwvaF0Bw8z3jH+4A8WG/Fi/9QswB7ryaNLxJ7yja775LYEARoqF3iohxJI
C7VaXUzsgUV3Ijn7nfJ0og9OXHlKMaKdykQlACdjNzdKAXtn/FPg3Vf5pa+rxjl+
wF0oAdcREVzo27za5k5yvXD25YQ9Qwt8KtvE6cnGD81cszJALWHA2s1kuScpYgUh
mDORW45TyxXuLRbFTK5REVmClRAggjp2j4+KVsnlzpZGv7D/+3oYDYY6t5bYLQfT
t9/HE5LyiBK6IWR/Kjm5ZkBpTjr8lq5cTmUVXF0KhPzD/2BIyC96fPmr+v+BPoCS
LKt+OoH/Zqr6uMv08Cc2s7KAMNi2mCG2EioTue82TXMWuz4HwscWeRaGzQVeEpUr
aGP7SmJ1M5OFyW35VBObjBD4f5mpne/o5oDjYRuPF1Ow9JNsOUrcyrrD+9cl+Ev7
/6YxF2zJje2q5eHos5g140DZ3/Jr2w802DBNdrmLuQX1qRjwCOKuAevdSEO++8Us
mOWEbdCZ6ler0/do4RzOe9KkX9ThVzvzCBh2jjAdEYvMPi0wAGmX22xifCYAnmyF
`protect END_PROTECTED
