`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
e8gyQamJfhV48Sm0bomBEzF3PH2vJEtbfPj17WchJ2TounOq8+bGIUDnExcmUAdG
1sa2ueNWl3ZuHCq7xn/kuFqw1JXHiOtL6mjQ/oBS9/ev7B6VUn28G3UURhl1iXOW
7fdz4ybLBSQo1c1MT3J+dsMlGcTGNW8K6uXYEOlWnBhHMc61heGZxL3/HzfNLqRp
SSQyqqSoMnHVGgCHMC/7netTqrDr91rW9Fw+/GXGUBMQc/6CbJFXDHsWnFDZURSv
y5VetviVNeKow26ZBdiESqLLlkb4Yn5Lo6TISeUuDfmHPRfjjB52BzzccnvMAGln
qryqGcdEiWabaQf7grZaUAYq2lukyfRPGloghblly9srteodzjH2QJcvgo+xYxct
x/tx3WaWrRXl/rB/Rlt7xTsV2b6NUvA0+blY1NbMisna46zpBjO+vnvTEKrlC9Yc
JB+5B0x5QjOAUFxU2ufPw2tuha6puN6NYQaPdZKwFDe/WA28O3bAqypNaJKS7VeD
2pvzDGTzVSE4KZ2riX6kjk7igIPioEaeVX43yOg9beVQ/fEV5P5DGLKd/MHVV7Bv
hFKGpCaZjSa2iIxy24o5uLx8m7gIcIhrfC/DX8PMNzdBKHPG2soKVZJf736m3JXX
9Q7yFk9Ugc8alWexPUu9X1Y6CtSJryZYChCAYSX6eBR8lqWfyFdDuous97Tfa/t4
8hQpLlhzQbVUufhI1oXWKWarcfbIOlERW/mjZc1Qg4bOc5pFvDFd5aQ5AQH8qiDV
9T89ipez4Wr5vrWIzbJmMxz2h2NLHCZ/4Y5DxpleikRBRChB3Bj/k9Kxl/0PziA6
rSaRnhJPu0BlAhjlVqZK67nodauG78+hlxjnS7PqlNHCSpKv8+PLXNSrY53DiQ/b
LSQdIdHhfsoEXGLqBFK7bl+XOv4HVJtbGIF+8dKPG6KJeATwDsY/82CW07JIhyJg
a/RmkMrEOK9kclnSeLAz5qNi4vV5LrPBDDK0jSBAvZO6BqN7i3hI271zSeAIcSaU
Grv+3GdTltnm13XTQa/+W0Qcb06xXp1vxsk15jKikrotKx5LwiZK9CzSwF/OVw51
M/8o/W4KIwCdSxJkj5SwQcjqBdEdsU6Csj701BhmdBKGa3kgSMwFvyR/mh6qn0RK
Y//Fp/wn9Pv00FQ625ewM8CgPMwHLa6KoiL0hum9cTwEki8hBOqClgwtTvVLHQQ2
ZXXyA3zURtnIlbgT0HyLh7UDQKrKjzvHHW5KwHgVgOfHcxJ2dlSOAhua/a9RxIfF
qq/rm6kMr429oUilcmjpZDRwIS8cS6lvORfKIMrUH5CKxo8r6+Q2JrxNQcBfykus
HG744YrQjq41PHkTl8SEC6DVahZk1xRQ7Rtq59jNmlM=
`protect END_PROTECTED
