`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
72DKe5MEZSH9IT4s+0rFcFzjEM/E+PwcnwPMnYOjQdCKfWP83R5Ifd0yTD0m+jt5
TpPUv86jcbCYpJ9ToYxuzmzKgWAdfkC9OEOoWGmnO1o3Z3Xqxywvs7wyRyybgj/T
IFTd0xYHbdGQb0SpJ+xXZ+OOHbXDdUZ9KpkcPEhJI6ux6I10EVsnjiUhB9oHKy+q
5OMoriKsjm0fonrPH0m9SUjRyOxE6CDGMr9M7J19iFpoNYhu6kvj2yp80FBw10Nx
M+d135uXqy23blg2AZ8qpsxvvzNqjjfHhFLKeBD2taoxhytX7VIfHo3mRv88Ksrz
j+EJo/oV1vZu8bkuonl3m0AqYHXg824693Mnrk3OasfV9vFd7NJzr7f7zMYKGelc
`protect END_PROTECTED
