`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/Uqf53bJlmtz7ArxlQTJ5qxKIBlaDlH9WBhrHrXxY0Q
H2zeq2Q2Zf/VNU2+0H1YB1FdakG9MYBPTz9urYK4IH6J+zWCc/IGeYhAjb2i9biw
/Kp/AIoMkVzLZ1dYblIaUa28FZXdDzI9vaZthAkwgNF9L/fXDVESUNaS81OcQkgB
77owG24RlfKEbdRrH4jmSfUeyl50N4A/KlbnQqsVFVx/Uu+YmZABfMNGRJWyCHs4
5PYh/xatcNbgJgaiGiwKTLpLIadtXEzRiP4xrQbZqq0bEKjPHiK7EF8d0C6jq1hV
H/uiVK3PZpfV7WNyo6VGB5T8lGdQlIHgh0pMCQpUi9GhjzzHbe26J/vtKATt+P70
U5Iicvc74HF+HoWcEagE0w==
`protect END_PROTECTED
