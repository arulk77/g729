`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
G3pNAl4JAwU29WxYVMUGdJ7NpcpOvgoRolugsG4KBh6Djs70uyghVYHknHgPCKkH
Z4WjKuxxyyeIV/+VvlEQWlwEUmYbJ64wdPdY2Y9N+B8CvBnvzFoW9jlwCuR7eHP3
GkF9JD8xG8UMMK1iHFKy3EbLehra2LJu4QV4BNzSVXmeE9+BqNCjQwF2yfl+P3wt
rIAbM3jaCM7m5VOrtKR6iW3/Ls+QHvH4oMNcQgsZwf6rG/7uiLZqzRIlxg6j0Ms9
RjcCASFpM40NDY4oyA85e7EsjbGOOiKFB99Lp9lYVtSc9+RJNGpwlwozePG4TqwZ
rJADZqMY+IEm3pjGCMYgEaKpIdLyuqaAwCmP39nbBQ0=
`protect END_PROTECTED
