`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKQ/ZMpNFTuoZMFmpqp7q3rXPRqgnaCAw74xC9UlKepk
a9ttkmt5u+EKOAINus2i4vU81fR0eZkHhYNpi6pVKK+7Zb0gzeYlMWMvT4bc7PPg
9ujTvpTdY5Bwgu7m14ygeWhPVz6eXV6vU2d349RKvHZuNfIwcz30mux5+qg7gnW4
BYJ64MF1oWuAH+Ykdi29BGVdnnXv7kixD/VIkejX/YlL11nMpFJ+TmL9nhZGotOE
`protect END_PROTECTED
