`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGMHAWHNadBgBq/lEWxKOziktwIAjWs0QiDfBGo3wXdM
xleU/CcdDlch/TiT+HSiiRGN8Q3yo9SH9MB8pfrXHwq6BrFD9+4D2hoepAZvXj8Y
iR0vKmnWzDhIRvBHgr3LKSzP5IdA30QlRvmKFzpqnyfSwsZprR7T/uTXWC6Yqsko
MTsmZJSB76yGYFxLssyMXrbINNH0Ajll8SO38r3XElecuuwMmX5MZZkUu64lexFa
66cUBYCLvgZbc1ehJQhaSK58JAvsvTXwzV3VBkNyQS4MOGpAnU4HQf8ktjWJrv1n
yyVoyTqIba4AO43rd0mCnA==
`protect END_PROTECTED
