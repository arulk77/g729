`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLb2nmHk5y/8DXoktke6n0JFECk3UdeXhgtndRgsIPTK
kb1ikqke92gPx9FEaJ8ZNTMaRS1jWwL52xfeS6/VfSOF7GL7QSCid8nHjsAsZ2yo
PyjJT55qQnYGzVfYK0ImnEGm4PX7XR67NqHoPVCJBUHWB9kTACRpWe1EzTc29jCh
Z3LEsUDWtuMt9D3+N5d+hekEFzAi6O2d6Besht+h66qZoLwCL74/F80pKbMV5bmm
GCd2CnoTuttWPVwakwfKCsTETOOqEU2+wcd0raMer4bg7Q9A1YkJNpYhkDO4wAC4
18BffirLqqJBiTJW6pez0tQ0qZTbhN2hbhPh+qm1wjt47sHXJbsx7ZCMiBnMn07I
B7wG1AruqGthrI1B4fvWFg==
`protect END_PROTECTED
