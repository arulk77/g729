`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/3bIw8e68M3frTXanCdPMik/p66sePBe42R1mpn+YCS
NxZkils5G5QJiEC6ONllJvHLhQ/rHIHeJpq2Zdvg9eXQPxk6b7TYLNZRyRYHFP+1
OfQTfgo4e9Bprcr4QxqboDEImL8aqKFDq66T79APyphtFVAUAAQOQdObRPJ385T5
iR3bqO4onq2J/OZ8K+/0o7ZF9gq1RrOQad9+GAc/CCZK4siQ5Bo6xSZDDCxBbXuH
KoO28Q5qfaPXdc4aCr6h9Q0JTAmUoLrh5F9tyilCSQSI6dmWJ17DIBuE1dGFkfsS
MoJ2V7LRBnGOP7WqEAQdGCd33XyG0FS+rIacOz8o2877LLMnM44hzrVWXoS3+331
Y4afybuFhkpEI7s3dckXfngDWZF6poUes8DAlF6t7gg4+oihKucFShbwSwBHvoMh
JRtkrRmRSvn7av5Ib9VWZAwWoRqxa+UsbFhwwQ5Aynqf1KY5fRSJVm5qgZQL3dO+
`protect END_PROTECTED
