`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C0RmDdcVb9lbn7/Z/kQ/2F1jKGBpKAT12Prk5rASnusR
nBsSCL7lv+f62leU6pB5keSf5pgSHyx8MhLnoPFUA2xCoP1oX05CLd/+VlS9/T01
ROHVhiQFY9bhvM3gGAkCPn3qFa1TkpYP86DI+CDy1qwDn5yJhwbv55KESHuhkekS
i0vD9uaDKQCsSQ4yCLVyY92Dur3cFUnpWF9PPSyzRSoh6enSaLFHAKI/r56TW7Aw
1NmZ16FVWJUCxUKakEL8ihV267BgOEu2zFq5lApm1Y0kB8HI80dxOnynP6ARGU2z
TR49gDHbFydWbGJgYm+NTGde1R+S6iMSjOcL1p+Ag+GZEcy4fy6eeMfpGJKoylU7
Z3o7sul3XXPL+9eQgMt8YKj6sqE68VRFeZL4XnUDwI3S+Jk+eeDr4FbZiJeDTyLf
ioR3e5B0roez7dAHbCxBhw9N/FhdowmhITGfBlcYfYpDRzjalG5cEb77Ysk34cQh
UtT5pQtp+3oz53zyYoANet76rBqXxlfK283wMQj7YEfS8bqkTayzdhs/bBQi+AKM
DoN5ZN0X2a7FkUjabO4u7QcT0WGsPl6mx4hCa53NeBlyFiLOtpZpyNDzS8W+b++U
jtwAO/viec9at8toOm+uKASxU6SQYJZ6nzchmyMx6NWCKbbZunaTcBhjxFqfNvNL
357yRudXz+7DBKPF3J+pulLNRCNQvpwaXBR0KxAZhXuQ8h1U23mhWiR3uibt5E6M
eRGNDPJK+WCs0ShjWlJ9djVQ8ZQfb6RLsEWgbwHR41qco5uXAqrsMokqfJqylcEd
tiXFETr/LU4G3RDddFR1jvteXh2Sl4al+U3ZxrFeOW7C4m1Wo3Cr60kk0YrpJuX4
`protect END_PROTECTED
