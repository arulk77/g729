`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
1ZXOfiQOXcAuRySHa6edt+I8mwM2H6/Ndw6raartVNFcdeTKgYrBrvZCZuq4yuUH
oaS2nTd2MaYYVW2+lvP6DV9nmmQbD3Mzqu9ejAesEPJ+BZ6CwWrPsODG8n1dxv2g
zMhu1hnDj2KBYSXUh14+xqzdummrliw7yC5OvFjqqa1gupws2GSPuT857/32O8Ja
Y0RVW0kAa6ZAb8xikv6ZP/k1CyiiInZb7z6Y4QUFk5x+6gKILavmbxxk/xB9fN1P
Y6tmHXBAbotTyow1O8pjjysrT4stqNkoUGYhyE15uIY=
`protect END_PROTECTED
