`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG43fL1AEpxNPzDgaEzBQZ8N6QlbV55wEc0Ms+37Jj13
Yyk3F6IkTDF88fe2vha98GqKeRMAmjWFylaCpwoBAu4jhK/9ab4Bu5oMTKP+M0rm
48NwjakpkPcz3Tn3Ts7pYfngjHTktmMA9U4yEYzdp/NJSZFcSTQlbIxB5n0YSfVf
6VStZn2kP5qjwohJ3x5ShBH3oFlw0wO5PrDSeQlMC8W6P/l1QO9PaaIjSHv5C8DS
ZFYkpPNsaNomJrm7eTRjddiXcSujHp1pTDXHiihhM4K8DyxXG0kGHSHBRcgDbWLq
oWke/8UStNrTp1OVkcvKk9nC9iASoUHjDZDwOWYb7bU9Jwv4U51PSE7MVBeAnnio
Oi/DUvZZtcPkpxkNyBzBu6kwxaj77f7waB8ZYjHiSwD99ExT7nTqZ7aQ/85jzgio
nzD0G9Po5rv/hYYgKRPg3OMtXCps80ZkAMCakScoyt+23QOUf8fjOdfaEd8zA+n1
`protect END_PROTECTED
