`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/p2IqJUhTJApTBWfSsPMku6shV/J0vn2fUBOz5aYeZO
kmbO6u5KTSr6bHnoBEJddWUyUtvsf7s8KAW6mY8RAhiIygXAVUTmdqgHc1hRvbjt
5EiDtlXFyQMlIfh24pRNPVmkqb2PCf3F0VX3ikteHsA=
`protect END_PROTECTED
