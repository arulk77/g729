`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNRmhqCVVCwZoBG4DaC1c3Bg76IrRThw74KURJ3w1f8h
cvArHyo1zD+fNY3uuO9NobPuMZItyxaedVfYddjqVh+gvQvDxYWO+OlXXeANfPb7
cY1q2w/50/fOnyYoOprNJqJSbwmD3vHAV22rRyg0AR5iaVznfu7zlSOpP93Gxk3p
Y5RMY5ZShGfxSML4iKA0Do+yaEjVD+xhb81pOGgU201CsEoLu98HZJbvk84NOuQV
POB43iuHzBKErMuukS15Lh9VYt+wHEUACcn96l2yEq7QD4knaaPZkdd0973sTE0b
Ew+xQSsvrellTMq11YxKEpdHlff6ewR4B+PM4A69GqKct6Meh5EU0hR8X8jkcFJ2
1qmcpIHek/SUCtfwU0fLHg==
`protect END_PROTECTED
