`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
/kZjYp7H7zzPZlf5MiEXpz/1i1TMaq3aEYss8kzdPmPxYHW5mLpRTGgb+Wnb1Iyz
J0xyCpp2YUM9hSsn/mOfV99BMV+BEJnOYEFMX4MbRjTHwZdkojUHxsbuRJnJe8Y7
4xV0MVwWz7DSNuEtBw2HTlsvxpBGGNXJ0Wa3h2tIKTRpoCyVGoUHxiUGdhBQZQjP
hW+5gRpttoXIlXvjjJwrp5p8zN0wQ7evAecY+EQAPzYntVQbpHdxO20sMi6aEc/B
eLCddiZkdEo0GwvTSSRsuIhKpbWLOHwBPUXSWPqaBrb2hd4rxSCoFLjuSeLwX0X4
hnsh2X+5Y1K9DFRRsBFMUxeFYU4VbFP8vAa2TLSmJTvHwq3P3MG4IEz0LO/iTFfp
zybE8Ifn1s/Vasn69YrrHfa0rt9XJNgHyubi+j6VjZ2pYssvU8Mmcg03PO21QBy0
oFcm2262+4qa3MsHNGf/vVFyTrKtwj6oRLga1z6w84Lznj03O5cevUE9WiUYxAHK
HkGVtkCVvv46llB6F4pXZVJRqRTkBFUlTBIDw+MzkR6MEq7/FGDOrkSKpJpyQgyc
Lyk7vrEaQukQDiDBygJ6s6TDRtfgN/sGHWwPbhX+s0hhunlUkifv2v+YF25pJDVq
9uWfskddduxzCgTmg91P8ZVfrViV1D7IOz/y1gKI6+nP7HH0rgVXO3mWphP5J6GX
xk2meoPCm5AXP/n4WaR+xpXEAHFYsQTA0XJOlZZs97fyTf93wHdcTLa37JSPQVbV
ECfPmu9GoHQW9LazjV+vQP+xMfBluI3LC8ia4UdPGDP01YyfBVRCJ/ttb9hR5Pun
onuXYxnljy3J0X6kDJbYTJbNk40FCAflrWum19Ju2XA1FqqzROBdeQ3jDppN4teQ
kx/R2w4wB4jS096Lb0zhgnAdq5X91roEQ762f2QHFpa4dSoZdGUiKUtQTO50HpbJ
fwkCB6EazudwP+Ad+ST4GJZ7oHchW1rg8mN+5kXyVjOma0tl295CgKcwDWD2Qb1i
MAzww/XX4VDIAzjhCgpjEhr2MyKIyBFN2123jNObHgxKDNKxvHEntKrWK1SLM2GK
RqOs6+culpRrVyHPjzB10NdYNry+b9m9xCeackTTjCxJ+BnvZSKQdHMZCVklnFOh
+uRyIZHZ7uPDJKkqbH7fect3nC6oVbyy0UNJdnCiQJfqjJoJTwNKKN4927wvMgXO
f5rsvj85Hp/EN0JSsBnl8qHXNGnVEDRI6YFLb6qYbjTan5/IOIVhWwA1bqICK/kM
o0D8Y4nTu2xVQv1sU6T6ya9CMQtLv8N211/zScCxLgjsaTSQ3DNAd/aYxsyPAgZf
ClfId41VpKInuQF2vgdbZxkB9kC6e6UtT+DdrxxSftyqvSVsZCNasWT02pZ1VFRh
n4oxyeFlBKB3WHKcPtTQAtoBbwwHKoUoiQlI/chYeW9rJqc3K/lO5AqWXaMFcYLR
mVRyhatwXNMOGf0c68r/z+bP17f30isO7cyXRqUh9mYAQ97aSEREGyBFVdkkFCPn
wIz/i6SwhHk9d7fq2m4q6OgERChBVbZTDTQ1qm+F8UgfvL0PM2dGoRsCFCailhT0
9iafMNA1JhbG/gGgDHvaRwflkmYuphB33vsFgFEuslkcEq+baEzh5AKT4dTVEATX
Ait0n9/b4enGXQEq9Y+AOn2qTiS8XcU1q58+ls1t28BLyvlcifybTCwX8ZskJ8DU
eozZtQ+z45sUSUdACKAdeSiR4VQUjHXqEVc2/+SVQV4xBl9vPZqMxAgJ0Na1dkhH
bSKziBqqZFz8iHy3rRM3mpLc9aLxvfm60WHYB7nwQp12F7BGdx+kEU3Ub5sSsf3L
daFrFzUlsOGmyZZUxGElmIj2Ez/f/7uWNySCt2eK3YTIW4xZvV9WppUzo48LUHf8
x8Z2p0x8ih4jf+5+kfpy08s3h3ADXFXqIZd3TCKvLnIgVlF11VUGQIfFARVNw9xB
d6U4Wo9kYllT1slhIM+Da6S53GkgqXsbvd8I2YWEUYo=
`protect END_PROTECTED
