`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49pAjALp4pRbOpFN8E1Bwe9xXlKJEv2WoWddV6IlKKxx
uLvHLGd/gri2OQBKl9ZAL2cna0ZZgkShliGlrhKaS18CBY4fbWSCwRq7T83RuzZx
POD5U8m1O+zbw83CjYq4D4bTeAVjPA/oKZFpYN2HEUpLY+R25DefSos0nI0KKuG0
lsPo+xoeb4THLtrjFwts8V5vOkw4HAqmOxl6C0uoQW18EtLyrv3P5oSdCT+kGsfp
ZCxrnGSLb87PFxkblsNK2a/UlSVRMGDSU/OdRnX7PqRbePTrlY7Rw4fZrChB9nRZ
BpxOFJCYFhE3BAgfovk3zw==
`protect END_PROTECTED
