`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGOYKckNEMjebug4W/xgYB8C+qdPdjHWoqAB+8QqeAP+
faZOr/PcLE7/CY3Mhe+wzmoIO2PjbjJy7Jz8dv8EGQQSvGj3v99iTSDpMVjGrG8J
1EsI8N1MSQoyFV1c/3ViiOph2eIttvghEZrqbElW5hL/Kj/QFlPJoS47iTQjeCC7
6wgQoQVUWtBpHzoQJb25L2QAiK3XRtPdlDhq9cRGORMqLXrGTgyPnuFKIdSV50DZ
EwmOR42nd7JGTL2sTLHQRj6n9C+VqKb3cbCWO3rZPvleXcJUFbp4oYRPriMPxONd
3xPzF5Zy+DaJst2zQ4zD8NfZoA+mSYrJOI/nyVGwxa4qQh0gAqAkfKsrhGdaqRiY
Is5+n+H13yUtBxqOWZzIGeXjjYHXut9F+rIZ0rAYZRyhAVVnLd0XCn9mpnmxg+k0
ORmUNnqO2YEkC1JLI4gLxr2OAZEXudGfKUGwKQkTz7YK/mLt491y/vLGUKZXnQ3h
/kxp2xE0UtYyKHMcn+n2RcFx5mCRLnpxVSYw1inw9sqlxQ8tESu5QIJ4lipG8dzw
tA/kWmoXL9B4wug3eN5ZaQ==
`protect END_PROTECTED
