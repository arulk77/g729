`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
a6+eQ1Q4FHg60/edNwwzUcXds/4aZ3xV7FVprhViXQdMBaWM4tzPCsqd4Ja5CMZZ
xs/o+WFmimrOAS+6I4rrdCzVMXg1pvyWjwUzjNHn+MIUpHze58T5KQzCvizFtD1q
lqtHxQLgS6wTDRUeUYlRwTMdj8nwkNvDZW1zAtpZ5oz5IYipNAwl92gSjH9zzkoi
Ygk5yR64TCuDGSlMqynSseqSxfEHjdkA5UfDbp/ghxzLAjxeVBhdw3aM9BplgMtH
mUcLEStBWr/oJq/+nQ/k4KQMmEZWT7VRIUM7hDFCA+4=
`protect END_PROTECTED
