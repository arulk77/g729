`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Np1IoYBS/BpFRb55oXC2VTp3To5w7F9hi08djlzQwf0KNqImoZbMbkQXtFofN/mN
Z3jRUfv7c35KMk9ZufDkMx7y9aT8S0GGrSCP9vNSbtGvdBWVWdxN6pTzxKO/t4Y0
MfQiVejccp8DNcWnfsdJHv+oXtM1ov22P2x8kUm37V5wq8TNjCUfGWo13OU9YnMl
`protect END_PROTECTED
