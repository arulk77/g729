`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM3B2GP+OwkVV5pJLZe0U+QgqhKd4jcD6n0JRkrHutA2
vnyZ4Z9x1t7zWZpRKizgv+94g9t0b1sAQImvQfLaY1OdXFLkCJ/X8pEedVibDiae
ekaO63kTItYie+5Pxm3skirwwcHZ7AwjvM4eIRNVVj4qQGUWlLc3sFz07VbEQdIR
GJV85Iumx7XW+9YCQv4wj5BE2OSumh2l8lNnjP7Zwrzkgrb52vqXDjE354VA+zW0
Hysn9lAdbmFx/7UofC77q0PK6sq2Xz50dDF/2GkciGKp+U2TP4EKJBvgZNXDHai+
is0QmZxYoEyHVaNie1zYNma7o1aSHGXGeMI2ypMpwHVZzYR7MGsUK9NZ6WjTryBy
SSR4Lr8RQjUrOt6OdpMJf/UVqFoW+0AEetIRrZ52eQPCpr3ziUfL5kGbWzp7+YYz
o1vJn3bauyFUxKTb6lIcoAf4mlXIC6iGkyv18nXuGLCoV+fGHgPYNyBt33GO8H7x
Dn8CLv3EF1Axmkv5h2OYmFcnOr2opzr2Db77KUbtynqWe8KrQ0Sl+llBeX2L/kE1
`protect END_PROTECTED
