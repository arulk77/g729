`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
xKrsOKeLg+NtToXIt8oeCttOPOLiBJkphCWywyeKmNJEqZFsu9LVC8ySwimNUmkB
GyClwvB6OuczjPIKCUYMNaW/k1Hfdpiz6AHAnxbaQMw67IES8hIfJA3+oITbAC4m
iOfBwuxzCxTQ02VLTdi3SL+PlsFuFEUWuvjA7sYDHq45drcHVnUkZIhVJpbHbxuh
TkXN52gTZ71iUTHgwRSLzhlcnFhz+QAG9DlZNSVboMEK15pBU8brZ8quDIIpj887
GlBN8ERh31NEZHZD9amq54xUD6gDCNrcJYLavdO0LwJQzaDNwOGVVBD+YdhLyNTG
7ay6Vwo1ZklQHYooSD2LaDsXkTK5qufHBotxF7UffR/aJMQ+Fz+Ipnu0oL1TvPoQ
+t07IVV0994xHq01tJtZ2GcddyLhe2GaEXqpXqAVXQalyOKmW21UyMKEx84GtIZc
CihbMUAd1mrzMCalkPgOKzIRNxeJ94WoiceKNWI7N7T9SZeRG6fxCUDoomaEPtsX
zhdzHztKxNi1IsXSQSyP8LtAIWjchb9bbYSAth4X0QrofVvD3Kj0FPPhpPcY74ls
udYWoEB2HU7x48RiQMwWng==
`protect END_PROTECTED
