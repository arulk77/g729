`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
r0X1v5Kou5RmZz33Pmr4Hc1TWGQS+c4I1ItnqjttPkTxhuVU4sVF9Ar215tb4BZf
FV5WWntGHnhzBOdAuuq1qHfrbFSuvohcf2sqZi3oQ0J4bWvolP9rK1HbWbO8Gvh9
gVtYlDGt/o9of4b+Irxppu57xkJoWMFR38mskiYK5WutqOFD1na34+aLNU6asCOO
rhufxbsolsDhe3TWLQVJp07P+FVcXieHown0W0NqGThZGn7NuWYpI37QWursFzSE
+HdUM/2f+QSt1WaCiDKTvo9nEyTIOR2Kz1nn4uzHYTgucZgzIRqfRYBq7WSU2DN0
/+EoubF+TRS1ZrBarLmts4exbkIysQnUchwO+6SQc4o=
`protect END_PROTECTED
