`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFewCTXc3fi37v6RncnOEptYaCsPT/iFSr3WC//zOKYu
SB47KETULwmsUOranMfdtUKTWVZ333VSBBfLBM0hKCMkkPgzSBXyYRf1Ch69mD7G
xs85uAT8QQbNuLa02fpkMklAKZ4M80nCS5GiJ5q91kAf8hlgsPu+aCgnj06XYRex
QirJUL2muHW3/ib16kJFRA==
`protect END_PROTECTED
