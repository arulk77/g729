`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOxlwh1Oy5IgoxsfQWi0We+U0JqXGRnj39vu32wUetkN
K+M+SaGvgAFcR2xllpCaJQlHN+jMD/oIjCpzmNOUT9i/Z1uIxvW6JNEtL0+gJJbp
U1TMiJUiRttGLtlUXuaF4ZIUwUPTXtS8Hdqc3/qRwyhE+d967g4iAFY0kWFthszN
`protect END_PROTECTED
