`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
VkGEY6dZXzFZ5gjJOqAK8MX5Y7q6qVt02bJWgaVVmltiPYK6TFdGGd6gyzas0S6N
LJS9havCZPHKgSTqWdAOROFgm8DQ9n3EDd2NqX1gn3nkJugs4Ign4whNRnFbaUtq
EyGo9AvsuCpN4ZQEaErvarrN1LY+yyca6zTi0xzWcRz3XoZf/kIyzv8qeNMWEywy
Ez+j5m2Dif737C5qqo2s2o4N+0t51wBbSgq8JMYVF5nrTjE295qgXi6BjQmLC/sv
TMj9tqKwNdLSyj9HpaJ4zy6b/Co8wnj9PpeTrJOgpjSVGrT/DdOI9qyCDNeSc/e7
65LSg6SzAVSv4/8fqVMTogUc/uY70Jhh1cJSrg7JAgE=
`protect END_PROTECTED
