`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SaLsvCBcOWfmrbA3uKIIi3RZ9VIjeNp6DpUz4Te5471n
kLOgvQ8qldLx+Atw9JAzwquRs3d17qbVGySAWZ87HwKOkyqcjzhcXR4pdZYcOms+
xiyd4+DPROw2X2jXGtJ3k10DAMZa8PX08ejDlXAV7PpafzHfd7Zk3T2EgM+QhyJQ
apKbWpA+cHJa70RHuQhIvm1YCPme43z9q9EHsutrOiQ+FtrQ+G/HK4tF52wYk5e3
6e/WmWhoDkI7/XGfmyWXNJKD1c2zowLhB6V7fNKn/qKxQxSOuJu2gbouZG+fukv2
xTdYxRYSp4GO1EbRWXFKIBtBWzzlDdKY+5faIuAtcp/CFFhgQW1yXXMbDG+hYzSB
11oFONKTz3ThVsg9PwOTA0Nn0uG3QoJJm3XDdrQHI0JinDHJTAwSWBBbscySYeGJ
H8WuUg4qtn7lhdgRM6OxIn1zoNlaQARRoDcWLmEhaV/bhb+C4jw+zofUQUtntH2M
RbTe3UL4+WVDWDKA6IC3ddZ34V4KcWZc7ZB+hRlcvgq0lSNTU0xXRdU1hVgkRveX
wnmQ1aFKaAlrJPGQWoRQaWXKNe9OdPFQqFU/IlYQ5ho5w0N9PoKI/J1U0UL5EsHi
xQsjrrfMknDaYUu62mfroeF9qtMzWtVKywWsgNMoXRlAw9q+B98962Hs+MaU3vPm
CHD93oLvySDtYVfWMNBQg2BR2+PB00eU4kUMiAJ6PqW/m9sK1QdZpIPEC/4y8hmt
B4L8hPGUlAyFVXKPmfuPQZbjKeZPTRVfTSbnXmmkIExoakPVtY+BEte4YRjydxuP
aGK/5erj06uirIFa7OT2rgE4zBa/V+3bOoSTl3RWgqbn1VQRoG2hJR9sNXQptfdB
3Bxf0J9VHTY+sYt9JqX1BTeZHp0hl76nN1paFHxshaBj5hFAzqVLrmdC0qfdN3Mi
mPty3aDfD/gDirSZbzRprthDC1EYn61MmZrvCkaiWgc0aE6NzT1VMoAiUCKsW1zx
z/aioUDt0J1mhWJaDQcUDjrkf1T/GjqJGgb70Zzd2rSTXvlrpX25XQo6MEBbi12J
vQIk7aApeL6jUF6cZRp5m7H+8mgCsINOYPte7W5drDUu0gu9mlJeNJB8YY8byIm2
xWiWKLtXxq/rt3doG7DJ4cepiDKtIYjEQlcCV7XynqDkinDov6c7XTZqXgEsWkRl
EYWdRuNQD+TUw9Y1sc/nD8IZdWx0jmlJ3NmILebuiihRbOEfNt9IKx28b6hBL8o6
1nVszjwsaMRF70M2q18Mt+RcNjoLFnLbaoSVVDGAwbmyQ0TjM0jGEZccLaTSznd/
94XvYYl2aZ+VyE4+DtVaM9Jdz5Dn5HsQErdqTaPK/WCBnZ3okJfe7oONgcvSe+b2
Nu8TRomu20YWrzXXUle+0e5Dw8cmJkRVJymURp+MFxb1ccjwubgu72/KaghMdukC
4IeYYvxn+68CWdt3XEVFk/46YT4CFGC9aNo0p0HSRA4=
`protect END_PROTECTED
