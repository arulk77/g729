`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePLWydByHfo1hX3hhLLE01+hCwhatjktmLupQtDMoMRI
g4PaqUSet5U8qusgg45OphWV3rROMipKygJyrCEpkaRfddwNKHhcQuV2KopylXir
FQk0nWjD9faEv5rzzhsnqjg8XiAMCUUkcfBFwMMBqRGEY2kdeIabCvihQIpPj6jr
`protect END_PROTECTED
