`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xd2GhrXJAZSZPNtNWH92oLwDFudOgy4MWT0lgI5MnKZ
PINlrP/rtOGiawqQmBuQdE+nlJ3LjIjuRUExR9KMttaIZvEKYBJ/lxlQqf712S9A
sobUV97YIZT/Xn8Y7WONpW6qh9c1JTVY9zDHbRIkK/btkqbbLjYKA8rKUniGoqCX
8ZQ9rpTze2LKZNBcgmMuNrKinEiBBEQ+aouHIlFRVCDdobVz0QpE/5rbP9rEi9lA
vVrVWztgBL6anErLBkvDflJbbTtwSQnABt45Kp5mAAzGOSpgtDHKEdtX0o/8zrFj
fGCHP+jgVIjJjAHPtWNxrA==
`protect END_PROTECTED
