`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
FpWjg00nHj+Y4V4msWxQJ3f8mVCFduQnaOZqizNm4xaQPjUTU9aD2wqt2Z/h03Cn
CsRfRYM8swZjherrganALzRpJ/oruXlXymo//Lg1+tY2TYlgWt6xODvrPYC4gTey
Vchn2P+PTRhOyj6xFghYq0MRBeO1J0kUK3fouIJT4JU=
`protect END_PROTECTED
