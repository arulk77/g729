`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/3s/aRsrkBNKTzU8eT4bmeZGO/o9hxXZyr1gzTa8w6l
qNpVkcXCYPIOKGn3oKE/aOma71vsszPwxnZfZj3s1BDj1vw2jL57MwQGjHW2eVOR
M/Q7CPGCGI90rGx2ugMvCFOXF0DMv04j/gfK6oi+umswNkhiJHBxmGVeK53lTmY2
fpg4ntKZgnuNkNH+Q8chgHENjpTd9++hS83l2pyT/nua/XWyk1GDZb6BWe/ib/jr
2qjLDDCDd6wDSiZnd3KI6SWc7cUh0ZnGAWgIe8eJhHnArmd/vyH9vaSI9JSJiLV5
qGbSdxwYyNTI7vZ6YDZ6l6g6dyuuX0e1HdZL/KhQvKmX7UgCIAS4vz/Pmf0NFbuE
2v+L01jtZVXDVww7hsX5RQ==
`protect END_PROTECTED
