`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEcSPfSeiOLoZmfcqEm9ptrvf2Ap5dNbnk2Qhx1PA49I
Y8uVv0LU85iPdDps5kk5s9gRW22RWdKj7XZJOlSiE9QTZOKzzsRJaK8uUO7eFPCg
5G71knyw845CMR71mLx2/2PzpD46CpaEe2yCG+Lf5XI8tnzmqZHPISGndsvbLB0v
6bvXSpYR2/DDmUuR71/SIqTOXeHStfrvmNflRkAcMkFaK86qI/UtDKYGwqFS8+pY
`protect END_PROTECTED
