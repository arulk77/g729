`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wQ9JqIfU5QSaudnn/KhuCV7XX5TMhbe/UdJU6HJOlc0
NnFvzGz7SIKZd11amO7qPtk83JKl4txWtsX7EPHNL7lMu3RmMkUB0HUm+ESKBn29
248Mw9D2y9YZ+baa5QtRfx8iUPb9MhYgiygBaT+8GKUrZbyJwTLI4MdUr07W/aa0
NXwUlPKlMYmY87rl0pD9XZskxmcFWQiiTFzfm5yPXYUYhapeYz2v8tZRvWhn3ko7
fFjcxJrl+UAQCEvmUeBh0s6lhg2enGujlRptxI7/HGmSIrATbUKBT5DCbLG3aDMB
gqtpo5A9DKuoEfLbQdA8fQ==
`protect END_PROTECTED
