`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCUsjLInEAuov/8gF2mlmEpdNfwmOJ5Pyh+CP+iON5uu
bQG6O0tvA63mInk51P2dCWWJT3RKxu3nQSx5ZsBC5Ek+Bt97Yv6xSmM98KCnBznD
yfk7lC4rRtKbXFN7plivIMcWf7orBiQ6P8OYixyc53dmm+So8dxenBWgHYYfHWzu
QjZJxOSmozTcKomlACde/V4RbwrJjhJKE5oHfRNk/NtQtpd8bKTaKRmowKE2YMHI
IbK/VegWeXCNxfwuvvk0KyI52NkzMd9KpO8TwEU02HghCE0ksZhQEeDBeDG+1Xsa
3/0dRUsfzCJDRwZwRtE+wAmQGP7GTgIOb47E8ViYNP6Ollpb7yIOnGxhRjdrOK4Y
hNAMn6B7skTUI/0XaMmv5BuLJZ3aLSTLVm/e5WLaVzz4DRvZqKU2Lu2rcl6WlKe3
leLzQ/zETLMgviT1JOeYY9ZskofrwbKP/YGplyKYlll3cfqTxKujSsPJq/FPj+7Q
6Ve8r/1lUG0W72zHO3PKXg5faXH2SkIXeW5+QWML6LEKzb+XkPQqz8DkHjXM65gD
4RvAEAtn4m8eBMTPmXgl02V7WjmK9gjqF3PbsJFRP6ZhRtrXzFBYijd1PrmDbHwo
o8TnV3l8s9O/UShIbIaewsuypth8xHvrU80+YKehyzx1w92C3nDQbZ0za8o0eP0V
`protect END_PROTECTED
