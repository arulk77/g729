`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePuT4EJ0k1dRGXd8pVnnzm6JZrNXBDQ8qB8nYJxlLz4C
a+sDrr3hwUGD3a2mRwMNPstdogdsCmfrUAzvY0+/UQtP+way+FSPdVwbWfR6QhH5
umF5/NrL/z/B9LMPcEJjlo9SKDY2y0EdmNqiy2z3rFr/LfPUXeEXKMAxUHmWyNm0
KyItnTlYdwuBOfZC+Cp5hahEZSxallqKBIcZlziV0t3jMbar1dWXtKbHx+m/Bbwd
pr+AexQOeKSk4OFgTq7SCzQznahs6o2CW/vjaEko5m682g98wPEJ213BnbqxDB8p
+kGBv4KaVnnbhMqqiLKkc05lq6I1EreWKFzLF1WtNp6Lf4EbjzSe3H5OEQFm6nsL
`protect END_PROTECTED
