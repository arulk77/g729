`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF5JRcfLHk4EiawThVAaRdeCslbF9UU0C93uKK2ke07G
iUXMAkpaG1VerV4UqXXoy2Oi4Fwpx0gzWwoDuPUNOf9uK6U5LF+W+uwej6u1JI1z
qnRXWZfntyWjQBlF1SH6WNY/kQAi8Ll1XOPuvPM2HrfLIDTWepG3dmI9Y+zflPqh
1H/QuLdoWOh+O95nU3y31Z86kj/afhqtekeTZBn5kZ7l6TMMDUSr7lqnvJpfi2xk
gemqwlf/TWIzEqHjeLXLL251HdSKdYSKUw9CNup0MVmwfMhlmmPWdX5TaVcw7pu/
`protect END_PROTECTED
