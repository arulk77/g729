`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4ynHBiW6Dg5hsSv0qfsN8gl4NlPtXKxICfJ+NgsSbWqL
8EwAQRZiFMeui6fQyck1ZRXEyvfKGAeIMwEgJg2jKJqPbLrZJDUB3U30bqoD5Owm
PdnBPVvgAkTmdbJcYUhQzGKfCrthM2aAUZ60Cuzg+yYXeO82eFER1tLGMalIOSsM
lIJlHLTHyj/Z0fK8PAxnSh0lvrQeifeG2wVRrK0Ly7+qHRlQeu6P3Zexn0hXxsao
CtTo+oAKWo/8wGmnS7MVUpEH1jAqpsEncciRcW9XqGY=
`protect END_PROTECTED
