`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ivPSkf9kJsCdwbzrleB2MLqB2+jm9ELrQYnYbhfKDEExYbdxiYV9Hp1uaN5OIMti
euyvw5Eri9psUNKwQwSekcRHlfDADm98BybPGZD1+iEMb+W1JHSrf+ACb1d4pKDH
eVhvqwfZ4T4qF0SyRHpQZOQFP4NIAAae7T7g2HMpZF6rYhjcqgA3wvE5AWdyahW/
6t/lCvr69fohHcafA8wqYtMR+GaZmBV1u5sKnmvbOZ7cHHJ3BYU/O1qfkB20l8LN
+nApj5eEGOI4+zf9rSeAe4bvF9Ns7G6JmShB7gqS3RxBRzuOUAcTHw8xvk98Bozl
PdZSKQb5KFn29pzsqZMbRFHm983b9uQJ752jSlI0ni2RHjXFtdQsOOmMraZ5cG4H
tRygwT2pSLVlMfF4Lxh4LKUCkBMNX2MOd9QdmD7GPxE4zaLvaqLlOwf632fQ9etw
T6BXsG+1gyRr1D0dqHuSNxagywv+MkOy0zm/gWoxUG6MrWOFDeoIGjRbpya3pcH/
0HjZpfmN+putm08atUY55w==
`protect END_PROTECTED
