`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4z0N2QvlmWXrJBBCNfySZF5JXLj68g8OJFCQovTEMusU
2UvbfmZH2evViGnjYEWCBmlbCQkENS6cYqdCsSJXqhqkKJuaAfuQL/kOAUDZlCEW
+FT58BbJoh1vmJAYoFXIpGCXqW6Zy0Oe4Jd9q7Fd2PBeWjHHCbCH4UAEgef2nRgd
rCTC8opxqKjV96qfJXIBUT76lM8vwIb1Ges/QHoZY7g=
`protect END_PROTECTED
