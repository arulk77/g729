`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
yJsvB706hRM6n00woaZm2LpMfomjAdEMSNtJdqpw+ERmrA2dDL1GXi7HRphC6XFt
yFo7zZ5LUafc3XY9PU6kMEycD24K+Flw93RbtwVPcmvW3bMPJiK8EKIvMtW8Lev+
pY0XyBBqhr2bBYJ+Q0ElLemf09p68y+EI05s9T2wPsPqbvtmJFxwRoZKmkSKBH4V
+fx7NqhQT4ycGZentd2QoIIiVgIN5jQNxNFgFCD2KVrG20MVF0B5RZYEvtG7GlTO
Sj80M3QdeR++8wjd2nNsBcqEhZ3xIHYHtgpOt2CDm9U=
`protect END_PROTECTED
