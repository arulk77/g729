`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43HTAPvOiq5K7JCgPhdUWiUtDliva8Z/09NlUnSX1Kj0
kzV0y8ejZ0LCc+f/3AOMmpWTsIcPkCojPKBvWX5zHmvznKfPvaB1JUvmhqTch+C8
5L454gwp6s2d+UFwLBC/MdOAjoDg1E3BaU2uT3sR+FMXIpRRxBu/4bXXWE1c6oo/
3whPtYz5UgNPQu2m61LJFbcwE78XFGabRlC3EQNrJjLzqTL++dVJSAHqfmVYWxHk
P2NBVUZ0DMEBtcuHoKim1v1taoBZ2rXW31E7u0dOjkupv27C5RluvhtsAGaRBXpQ
5DuHLJLXW/cdPbPuh4o3scaxKQWuPf0OH5cReD/s3i6wsOY79+wUm/Ha3mxTuGX9
AqZb6AvPrsf+ufsgUqjrv5PUfBdflZaEhngtxrFzahGBvF+GbwFYKrQE5SJGrOs4
i+/DkqsgcvmYlFwxzA/Umw==
`protect END_PROTECTED
