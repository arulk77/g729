`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41aoPgj4iyARQyowBjJ4+Xul9UCORE9L9/CrUOXl2fIg
0MBUKAv58a0TjiEj/LXbrgKjx810LS0F2gngeKGZnRTD0hAcDVVaPHJSjwaIT7n/
2P8gSi930uUld7acbnYdU/kjsTb/WQLqsyrAAMRU5o21E1Wa65Cvza8P55xaf5ri
plCFhJiwsGYUzLJk8qHi8JtPT5L7UKdnd4an7IXKrDeAFXpXz5tGVUg4X/TschnO
jM8YpEPn80DYGy4digttPuv0Xeiytt9lFrGKduJtoIeS/FPHRsvRaLj2k23h+gly
0YBiAsWB6dwuRYO1UwwhqCzV6ekJ6OMCH1msbwZm13FCZkU6yNiZ7+PxloLIDuAk
Dk/jnqpX+laQ9/XzQ5RWjqnCHwLhuACRpwUqxIu+/575UoVDHypHrNDEw9tGyHq+
l2oflNl2I2+F/e6G6M8epg==
`protect END_PROTECTED
