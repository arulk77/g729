`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNyWy+jCOS3h+hphllOOeg7l3qcButealHB4wYm0h7nf
8OSaA6v1PxekDPVP4eHjWakKotTP+mi/uYULcMG8LERVzS6H/QkCGyMKO9iABLdP
va5h604h2C/32chSgNQ8fhpX85M2MbTibqGg0SvGqabL+/FWzhQes+Rl0jtKyO+V
KqRwu9BVkPFOC67ADda0yffc82LqZDr3yMJTBM2OOVG1dxYOcvfj/JCG+G4LeuV1
CtdLushpWHAzvSVQaLK0RUxB9DXKrNWATPtdNp98yVmMd+8FBPUXeeKjBSCoK3k1
d9L8YhzdSY+m2VRxiW+hcyFChQ1390rmDiIJ7B2sC7cH6i3P9Piey2ntoT4EekV9
kAZy0TF49GKu5ntVzAhz0w==
`protect END_PROTECTED
