`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEbObqvWpTX3NFdCu2pO3xUtXiZ/2p2wh3Qjhhpm4tuc
TG2fhuDQiqkbtGj3NQN7CKsU4mutatscocCAeXMIEAYCVS2nb5GUhrKzy4vW6iQ0
8zN/PXMwfZus2qukih+2xdrh7XQM+RiGpI7/TWLqBXlwJMfd11mxMnF1hSm9XI1f
iOqisre2aSD4I/qyy1u3Kw==
`protect END_PROTECTED
