`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAQfVz7PHX7lrxJaDB1VHEHab1XcCLo0lPZBUA/kd8ZVE
50ESBslTow4S09zTA7GrrX54wUo6hp3mh1ShQnFypt0OIQCNJy7o6eudzDrDG6lN
0r6tlSbLlH0w5BaApjao3IV0ySuKZhBSMcJObDwKAZbWZpIqpj/nv3YdJvyNQ+Hy
CDL+snHs8eP73lsDueQ8u44t41+egcFbmku4vKKET+LH2gBtTsggX4FuejhUAmQR
fjLidAEYqYj5WVkB7ELVUnuAOrz7fodyXIwsf0XpBBN+tcpT7Z2yCCBedc2wikUn
Os+LUQ5kJs9idPjaO4lUvyIHhNVliIb5ALLKCSN/ej3MFG/aGgoBbINwuyRtuGTz
nzeZOn4ASXYy7VAb8oOR7xIPaP6K19dc93+lEpFujhKZ5zBNHuDsCUYjcuyKJBCX
UZBcjqkOEm14AcYU+Fj23RcV5bd2NHHRzo54MTgoUmWtGQ0DNvknqS9m5CLzXGxo
uXwC0RzGJp+Fv4mfJbloNboVuMVkD8zfbp8tlwrYPoxPtvsV8BR8ETY7XD2X4hLq
KLx0TVVl1qi76ZdaikuPsd2yMk+uPYosZU0Yqu9z0a6hJHoycq7nPmiuKOJJgZ/n
e1QtW6LAW9/2gG0jQUwMUP8YRi3F5uSrrK5yL0iGhrsVLAVoJ4uGG9euEP2TcV1Q
z6UsdkMiRShR3q5J+9/SjJjkpi2ZfDhPBtIIeYdHQO21Rrdw6/bJ5lsVkKSSQ+MK
IgqQFmRek+eJr9cCtLpJ1PObOYGlxMBvxLdWordZkIy5Ec5t1tbHJXtagBV+5f8g
psC+WujOPWK9Ie13pdz30mCU0XEyJNqF/RgAqCMF0f/9lKFUVtbGhcdd8IUIJIVF
lS93emHQ71mrS8ZhkSA+toy/BJDvSAsvxLmJri6N15RtlFVCXO0E1LxFjNi0+ZgE
v7uHmUV/Vf8YheJchVU9Feo8LfHcPWO/ExcIiEdOafjmEAjfs1fa7BRRuTwVzLs2
X3pScZyQSyvLTfnh1ihE7xzVcZ4LM/RCu2n6uwkLnvcHFuNW/9m6IWbkWpkE35uE
nPJt6PpVWAHAvel0a520grqLhM2JOueZgJQ/yUoXYO6kZuu361JwVu5iAY0jRaEb
pUl01NjZbo5jHG/L2pEm+IJEWo4v6SIbcJnkjpbnHbxKHYO5NsKmYWX994ceWj4N
xLaPqI02cHPpRspY4ziC4OBRcx+mDf86ghbpyKbeiNKQMolpQKHwqTphwBla47Rm
RDdAKTeHieDtjmBeL9JfYe9RpeMPYi8iSaKY/+2hLbtUWhRvqs0N1Q92b7mjvvjN
xlLeZ/WBIYPRibexiSb7NuVgln1QzfoJTDcpQ50aRqAL/txvlMJ8FgpdaRJ3NYfg
TwmHihmVe3szP0p0ot6ULdOf5uK6LJhyrQZKUFqHuOIkFHMkbrJi4N9Q7d+wokrw
uPzS86HjSAt9gAqPr4aUI/84fu07gDE23hnGxozYkkp+DUIkWsymBKBnMpsGpHxO
XlEFkmCpO9/4wnwVMYfFTs0/IT91Elro7rgJRmQTgG3RBQduFeTmxg8QgRDS2g2r
`protect END_PROTECTED
