`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QtF7Sp/pUn2aisH26xDXjf3CsA8sFb79iIR1yzMfdoZ/sXkvFqejlOG1721obfCc
4BryouoLeVAKDwj66OAqaAhWHXci0zW1D7u85fd7ZWBg0ksy2IUlYaSvBLCnzcEO
aKFNal7+uu2TISJxpEClD4N5KBEQW+LLcx1bte79910=
`protect END_PROTECTED
