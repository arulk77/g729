`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN1qhFxrgwrL8UK4FRq53fDcmzLTdkumm/t25Vb1450RI
QA0rZVvcKyMeto9JondPDxHaqAJHF4WWFGY2yhFV+8N+2lIui8Rj/DUcyjZ61Sy/
maAyMbK7I3GAzOcNQS5mlZeNdJzMzMdpvkZc+C027LPGedANOTyKMHxnLRWvPpAz
KmuMR/TG08PJB9NIjwwtQYxp0d3PHcv7Tbzks/UIIeYkUC4RDI9g3hFktVqgjJNG
yy0fIr+KRWPrd6KvEnr+RnY0gAUQai3PlJF9J6M1895kv+Clpi41LcLVcaJDQkYF
sU6hyY/Q29P84JeYlr7JF4mzXRDdo5cuxJbrv35JQ8MzDaTsYQ6v3r/QxMzJinZZ
mohvDIPLncga3ChV7xBHMgN/rML24YWobDa/Qph05uUKSrrZxWPl7ANT3tVGb9Fq
6zRaZvuYc7D27qS+BkVjrp2VPfbSXHqmSR8gs89JRBj4kZsr0vpNeaw7G4OuKewJ
dzV/ICeZZC/MX5ftMqU0By4rCI1B1LBrpaPsr/X0zvduQZv8GpaOFlqd2iLaAW0i
SR/pKhlktdKblhCEPZI56mOqP0bL3uxFYul+WSkcVxIKKZwD1qSe5S24IKDJ7P8R
Kh8gGfBIul42VqbE2ObZCImzKtIoePG3NgdJL26J16jPsUkn4oKavo+zjzLu38HZ
RjArESrjOLuFKhrruUsTMr9U738+65G9k1MTuIkrCOrGbK0ftJfanl+WlFyoiYOf
hpR5UNvuZN2LjsaEp++vFz07bN5XBOgF9ia45sUO0+Ger8Tltz9kgevGLPltVH+3
g8clG9FSSpfi75mjoaBaA6GNrnKz4MYwI5l62E9ij7VelzL5+mH2s0wvH6wNNQwf
k1vOAeafBeQufiLNrzqjiZzCeY1YHQeR3mADjkvbMFQtRBTzYfpudFJSa2oJkS2N
UeRu8QBnsrCOuuSfES1vyENeK2MgPeqsJCiV733M1L6I9eDLaGTNMk6m+UF5RB6n
TS9P2f1NGmBfCU7uNxJ08M4ZhrtOyIWUEFYGWewxqymVvxce+EpucAgAyecub/3N
eBNoCjr5LVn2EVoGFlReOse7cVQKpJF6HN6xFIKb+IRuAj4wvxqeAoekDuSq832P
KDBBbaoL+DHLULhE8yUaHgwzT8eBoGtTxHj4TXIs5jSfY/uw+ee4g20U7rqTtqbQ
o0bPPyrgHxrx68d5CFge3qUxrD5Ye1flyAWRMMbioBKPQ+n4xuC/vLuSos9StEh5
ibNhzvMS9L0vpu0PoAUMeLRqyOS4sWKNs0Uyg05r+4OlDR6wEsMKwWzDOqK6Z0XR
f2xEdVHBOYM7IIXdAmC4Esu/RM1NhmOBcJlMMeF9F8udLHPAt0+ki48kONBq63VN
q4GyO50kgUpst6yY3+mpGkC54sB1kVJRQ4fZNknh1RuVGITAXjCfcNv69lLOXRW8
Lz6VWhmO64HBaDQu8Fi88G/URhd1lqg1lTTHtBr+vDDGsSsp7X0ArU8N84LRWeDw
rRXhiK/p5sknvVgcxGAHWSRA7HsEOxipGdFfHnS2BgHvL1nBy4xr70b65nAmNKlG
uv0Wnxz1yeSZReZiJLi8m+X99wUTjlHms6PlIEGaWYSFwxOKNMAC0JhfV92i3gj1
kKlf6KoBxosJDjW/WOFDQee0SQfsF/7RRNOoPsOGzPE8+3ASUF/2P5sSju7XCFpO
VKbB0MfM3fBnHbioyf+K6M7me5RtLdtexsT9OyRPsNcRkK3Kj6nu9zDaz3TzdH8x
ePgNCBb19Sk2qLi+swFtnS13QKgZOFO37rSP0jxvOblv2hiRFVmHnctcIaXLx6Kf
suuRIQGseZ5ZwvOUaCf4G+eNNYetFSuLed2gvXRXjR9vzN1F9vQkAnm7DOuqawT0
yNf6d9u2Huph0dCA29jfv5YDQODmGhDyChAezJJGi3ZkJQVEpdpNl7USHZyqVvr3
cGlOyoSEPyIqSiejvWKivFXseT5FrOPbyhJtXKEKBLKMhkNIiv3UUUXwJRPxXJ1v
PsP7MJfbUjonhTvyED14fn/VJpxzx+7pnTomQn5y2Ae/WUn+w2evGR31hxmoJBtg
owiVzaXfqERW7nU3ZPo1FrVq1sz0q+D67dwrekf0bUNVh/OPl4lfscxbe7oiUFHP
y3+4l2ZZSbwza+qu31ThdC0eQ9G4k5TGrtO9ZA9Z0RTZoUL+xc4FnxN1Quox8n3b
QWh0QTq7Nc+MS8jzMs7ZZb2Z2D9XDkkjTBFmXMAOtoq9LywAiRXhGdgxezldHwde
YfTSfELcXhz4x+egA7rn9uUuDMtrcFhZ/kY5T2+QIf3P90nIhT2XyXFWNKyyafi4
0vwU7w3/powGkhyR2Fy9FjCma3Gtm3uq7+2WDTZFoeWjJO6UdCWGrbJ5M+zsLNZA
NpJrJEjCzQkgCtUVs8wsZggHyoBqiy/UMgKdIHbMzQf52Nfb7mK4JAUmKpis6ThB
s+++IgqFzLiFdn7crC89WZpeNO86M+k0WFgkss/Sp8EyvbnRU/+fPhrkd2DmdTXK
k9NgtApwh2E6mqsbFFjbQl/91GZJtl/ANslpXtkx/05zm5T4p6FEbFjmU3mg2EJy
nMN64FMFLQrSOP7vY+VD4e+1h+6xMzf0a1XkYp8jjv9h3vagRowZH6qrhAcQTnG+
6O+96EEbhgwuEsuMr+wBYpx+xWYcAq7J1rPLkFWKUVn5Ce04zxvQwLYxzfG+IkFn
LkZu1T/TZ+QCEOSkB9dh4xDbxNqoQqxH0sugktbfUH3pdupY5y5GebYNFhLUYDTV
dlSPEbTaxDXK0sCIusAOAG9GBITVNZCWQ3XgW08jJRJocfwjEksplnybIPOSjs8N
t7WatjC6t27Y9o8rucv8+ZtT4dLqyEAzHDaUwsenOZW8gcj+wkK/QAu7w/NzFs8+
g3dbjB+DAzstm0erwjvGzJSRaxzmjuPg+bfb3eE0bANkCc86em3uNG7aEKBdRnZZ
dFwEdygDPGwXkS/VN3QsXrnVMJtU9gngLHTtsnkaRQ8eDakwiDHqOY3ZZ3teTx0/
H9K6l4Ndt/FCVgZT4xPwoFWsgr5OPLwBDWLI8+B4NUXCEY7+e3E5pMfy8eRC/gDD
B8glxqUp+SK/GT17dVpxs9FcsDghTiUQvY0HGDOUZ/MLvqpVIfHYguz32rzO5YME
wDKZnMy5mJfXnzGy12trNpDqpLpyB6wBYmAzrf9wUW4uLIPpY/vMgix/j7ARKbWv
+Q5hqhYa5SskCUlXsXttOCR+hVuTe+CYO5V9rkQGCFQtHkVX/jo1L+s6gva8Gwg6
ZQXdmsPdGZrs1Yk6bzLlZeuYTP9Ir8Z1FqvxNHKoqfPExUGu5Eukj+0ChFQJe/wS
vzgTIQ3b81hHTLBmd0oHRpooRKyIZtVZOCsUQJ19GlLo5v6llNIwiV7mkm5S+JfQ
gLQs/MFLh0v4Jn8A9DYZqLcMuLShRXz8RnGOOwq75OPdk3gvtLfgD/XV/J+D1yOW
k4GmFlOlUcpKBY7cXb5dE3sA4jVlSmYqYwZ6x4TvSerXKbgjG8P4chnllTbx3eSA
YGXUUwCkRly5DufjmMu224hG8VQLLgkU97bLP90SIx++P67qxPjNwGFBFO8OviMa
r/l+2iJdZav7DRh198WPagc2Xv+urQLkixbfDTS2Te7Pz9d4XU0MSZm2kFd1am2p
dLuhFnWanZkbwiJbGT6oOqpc5TSOcEJlJ1Q2njzR2PaO14XXXjNJIUqR/o9R1uZB
CJsTShBzKDcSsYgS8roMU3jvep2XDvPCmvjbr3P9ZyYrsy3uzCjJYoeP0mRAfbrJ
XV3OsOKqpymd4TGxpzH5tphNZuCH5p/1+ivrd677xyoyJeKgVaS1UIF/baLmwaIz
0G938IvXBRjIagk/WEAJ3XGHmoXpQnq77rNpj7TBWONr3eKRMMYcZoUeva5gDNKo
m1SJ50nCIYBntaIOwSmjBlI1PE1b2G7E2G17snalBQk03BvGIRNSZUIPGfB8qZAr
nXtNG0tgb5JHSczU6yno9MId3pG54a54vfZLFstc7QvsAX0CsQWDIvkBEWWaHY5F
+oDsSUKhhqe2gx+h57YqPJbt/dq8M3fmPBynCkYys/lrkzUKpW2NcJAg6KSQl9gV
zcvFLvXuGSajKjC0NFlE5dtjnAqaJPrBahHPpyBzlJaXDdEE7rmtJZaUcsFA0JQj
bLpXiLMHOHpvKYUKBMGxDzATE0Q9ki+fSQx9Js1m2p0389wxlmeaAZ1+uvfQkakS
xJp+U2zPnLlNr9FYkixAkL0QiG0KRclmbRbSlLJrNYK4UXGlQ5+vJizhPHmoX6JR
cl9fimKesdQXgQNsd35mOX8DqeQSbD4ifRP2XNRMMvTQwTVeEqvxaVq1+5umo11P
IsqGQ35/knjDqlM1dod5uJpPQzP+xiiVzIJvJXwkY5xhCN7S5Kd/mrHIn3s5dol7
jVKPIMlKWSLucxwb7YijrasWdcl/C23ImBJgU/PM+5fAoy7wo3Yf89aNpLG8HKw6
3a7bo8VsgbM37+sPKn/UqUlr+nlZ7+hr8RCgB6uNY2Om/4ybAK5JyUj77WshPg3w
mS8dVMrgMqRMb8/xBtwUqzMiiWganuQA5+m+gsbeFf4caE5vXeqqu0zH5/4lmFJ2
T4yzuqoebw4ynUo4KyoN+BeO9Zn/Cd9uf7UbPRIRXB4g1QkRiE/yiJHXaBW6g52j
yVu16GxqhbROVu5Odli5iVD9K8xMIOrdNkUujNH1WDJCx+i1M7MeZUKoPzfl4qNJ
U6M/gw4p73j7IxJf/pcpev3tFjbc1TwkfPDeOvl+VHL3GaynVkDE9whsKZxfkkpD
jDvWwoaGONSLhhztz8UZfLhmvyJgeBYHJUpofUwQYxgpCbQp4RtkT1WTotUlaMut
w8ZVUY7JgfReDl+JeWFBZBGBO2DZ1uwIfVeOKPR2A6XyqRWTKOe7piD7vlAYXNmq
48G/vAWGtg8RPk8e9WwpcEVg40b8SMKDHbpHvOI/OOKRiLp2wWlTMBnZx41Lhay4
Ye/sN83kx7ZvXQzJrNwL9lALsJbxHlr0osJ2TmIbBiWDT8085N3K+GhHkm7HwkAM
2VXyhdT4fJW87xHkLPHa8Rcu318XrS5ki2sZfSHGSDtSZ+shOUrDx5dR9n48Vw5i
Z9W8kR77LfR7g8LhTCz+BNYt1kMRWvrPqlQ2m+6VlJqM9jM72gc9kei/6Qk37puZ
uVQ8boEi5fccL/WM+pCwVM6f9aWQnRovRHg0sKVwnSOqnFYk0So/5DJvGt0Yb45n
uoTzdtuNvjXsrP7uelU+Ona7nq4vxafZOTU+26b0OnuTMkWDaQzUh5s0RChKxXBv
2ee1frVDHHFr99qcqfo8VmLfLjKbbyWQsxcWLx5IxJZxJiA/pfhZ8OO78YDYNyV4
8Ca4PMuU2xxbE5kKWHGiUcBfZU1tfAjNksoA+URqj1SYmR7HB/w2Odd4AfzbcwM3
oRbRQIab/sbTxTImxZNfHa5wzz5LSY6r6mIPpY21cTC+V8AA7fhCjx744ad08AsU
BOefpYZ/NB+vwWrKwg0E4i/p1FfvQfEbrtwsM3cszcA/gogqrF32ukvcEEghKAK2
9yj8fW7dtppeWH4wRgFIYN1McqtjK3vVQH/hf+80oVFEBltReFgwF5O6H98Aj8Or
Qk4Xx9eexAtxompmv8h8MMMEVQ2Wt15jWKxHDPctRvDypfJyfDR7y4CBdLNTHdtj
N2zEARLikNCwiKh1u/ZhyFfZIaYAk+QggkbB/gvMWQ5ejaqLplZwDbqcCvNJBId7
XBP92iYWz/BFiMMm+KIoiGIMv2JThV7aPPMs4BE8/7NZigxfdjmMenrxcbwkwSSF
dNjqKgOoesztOhjdPYSvcqsykFn/xdshd9U9mewjrI3G7Kdunm0qAyzLoU6xaSxi
KEO9WdwnV3IDL1fYdyybtuC0DgIl4zid0x6N+8rM3SRGc+w4V9rNL43XkZp9d2/H
APww7lvPuOo6p/e8oRLG7B+PJ6r3YhQ2GcS20D+BEsjADPs/sX52PJgeaBEiUUgm
0MsorG18EedZFV8MTgPl2O7IDN32rQbtoaAPNob5WBIisxGyf56v8VhcjmsE+SEK
HnfRPH/x66s+86/oc/4iR4t0C8QWHEMO0x5cyQwZQSEUiTPC9+R9OgJocVFjSBMB
yPg8kmuWdl4N9UA7OzUdcrflAS9GHQGPnefLjPuMQjTLsAMmCJHGioOH5Dzh4tnF
zZnptY18lT0XfTGMV3SmoLgLWEu4AzAFwZka3BgfNYZ684XbFsRx9UXuovfZZ6Qe
1aRqghcB7udtsFduYdZnCao4H2dc7mW09krl/pyWjdaNCMd6OWHDk8T12S/LR4Q0
aB4OYMumF1ch9A+Z224qsK2txHiOmiwFP2sqiV+yjAQlc+7AiiDjH8GDHXcYS20S
bIGn5q64jAzmfd1D47EieqnxbdvFmzN9QbarFelzTvPmHjIhIQeodgDSCzo/CA92
+2Qv9ibmaMNiOEtzGDbpgPgfH9B4xi1PrWKE11Z2Ni/FJrMoHsBKtG0BmGaVCeGs
qUVFvCR03H/J/C6WkpGrL4xmou9+EmQScYl9zJcZIUK6PaJ9L+rFL1dQHN+Oe2yj
R61LtR128FtyZUz/3P7rr0oSrVK9YwqQbCrvFWjEznTr2Oj+nuuNP+D2uNUsCEBd
bUlwf4MSzgJvSieAA8lw0CSObfGA/+iS3uEjsOEQ5YDlCwRGhJeuDiBCPA6Jgrcd
svPqRKhPb7E/+sFxbkpVDDIamCb+K38E5lGrwC2vRen32Cma00i/fsptKp2QuPYk
Ubxp2QR/WT+zV6N56rwy7qWsajqBrofLSb1mUe7NH6Dk1TowOZ7aw19QMz01Rpdf
lJmpuR876IP5AvKewoLKQ2JEa4Jtjo6Ypa0oHQ3Omd5DhQXJddaFyqJ23sHrBo5Q
uLI5mwoHMORHhIObhkWCDaLME1NeIEOpxRFXbmwi2pK4CT5pneX8l+RLl/Am1CJT
lv005TqJ6GS8EIzbbp+GFNmd3NkyMcBmnPDtm4++e4/8cGeZ5IrumXoe+Ff0iub7
XigAriwUraSDq0og7S4jn1NN+QfKc8fnpJIFPnj4bzPHa6kZWzmr+ms0ra7Oo9cp
qMdHq5/nQxNO9T2+etKEXywG7lQiUB6SWpeU1XQ/u/n48kIbIynejfiq3kNjd3KZ
WecS6AT7JCBNhICVLvVWQqQJwRlFse7ui+4Ve7MuCjsYGbJgYYqsjcz7T/wzzfAx
7Z6hf3j0bLWa7+g2PUq52xVI5+Q9X0CtJwQhiioBM56pun976VSGg6G3CbJZhNUR
FvJbRvs1Omzhah16Sa5vqae2WETTewZLmSfTyYF0q+cRv1YbfXu4PTGuYhXzSQdW
zzK2ce8LQsWeeLHLp3Mq97H4sALm3VQir1ovFlY7pbf4vOqDh5AoibNOhPHIkn5s
t4APDIALeZY8wD7AiHaep16CMrrp5jKIX+LrgbGFFZosyTJ7twbQJ9lpQrWgjQZ9
LKO/IvX2mrza9WvUvoYoMygTYAWh8QHXeQFRiS/OWIeGeGKmvDfHuQVCkJbh5FuY
Z3vPhHzNZNAPeCPh7IDYQX9PPy3yo5TmzlaN/XwamMal5GobA9HMc8ph/MNaovP/
4scc5C5EJjbbb3UR7rRBW7iwMcrhT0XdeDPRGfMsDNe+VWoyEIv4Hev6MCT7q8gH
TIfjZqp6uOZXJuEVZA8F/nsKVQL9J6llwsJ5Pw04iiaQoHRHXC/BR+uSAFJz8V+a
27h9bZXswn/NTEPnIEtBJy5tpErsnTb9Pm++WOT9UQYJ/0szxnqv+wtAksbeKvtz
69xZcV2wEbyG8N8xvU//S8Y0txqlEnnzTDGBkLp68dSrYGihktUzqg+Oa2J1ma71
ac7iIzAFk3x2qfocLa80UC6d8WujcDa9Kv0RJrtMbNm2fNOLpjz+dD1oOs+dxHVi
4MqoZTQHsbeOh3AphYiXUr8MTcF5TAjP7zzmnJJw7aa1Y46611/vfoowKY997n/x
77bagXkyUXN9wqZXBBuQqeqXzNjkEMKV7KYk580VRG9rVhw+M9k2cdFsTdxkTLXO
9rKpNtOjNyGWFw164MNU0kTRNURvx/zB39kKjUgq5F3pi6Vx/YSSetFrhN0oUYn2
IxVPWPcF1uL1ywUoDKByEjizgSwU4cPGwFySnicwtd64eIKU9zdZWsL5ZadgldF1
AqSRH+tJNTjuWNibTb9B0KYQfdAgOSZQ2+0REWCYRuYxKAuakOlemf+3RiRzuRpt
0vBnPVYanbY5exTeKLy02WI+nCyAC8ixT4p3E3+axHjf1Z1w3+Chp0LvjF4z58hj
Z3njzynyQVyVHoPZZTyNkTu5SuW3TljdHLkMxr/cVBZjmhL8xL1RHIUF+lKu0bFi
9QaYDjoERb4+hWU3Faff4qGVqY7MwiHTBv9BG6cNQzbmt/fJ1qvluKWNPppoX0W0
MrcU9s6mlrM8+LEB/CcO2Nnnh03yASS8yTDbxGKYMF0QEkayLtnzsTgmurJ0bvp1
r2XnpPPyCLHqGzJ5yy5XUdPh6mTN6acvxbFtjT9JAK3OjIdjBTrKxmmUHiLf8RtK
YQXipF7oV+2mtMEztjq33c2NnNSsfX1wIycxjczs00qDnl0FQZH6JvieYigujrtq
j/5o2q74tu5KeligjWHuXpnnC2MGp//60fPR+uUAqghR8JbY1pE6h6970SMparPR
O0LVVYxt5SDFqaajMCs1jmx63h0OQDInakc9hvWEhnboBC0MElynPFZ1mpdg2s0c
cGkjwIdG2x9KEQudUoRW4hmZccHTDtPuc/RsNa6Wexwk880jJUeEcL0lFdmBCbGe
LgS5kMm+HFPu/LsqENsZb54XI69qFjwyxJZfThW4bRQsU8cdygECyoZZsflLvmz2
0K0zLlFZI38vpDF/ddWc8ySrQDB7uxQFazENUq9vETefz9l0MUvQWt/rIgo+2ToP
ncyIR1gesKfgy0YnUx/OpwKTr2FudJ+wo+XsgEi3xg5jKfOtHNQW51PD5IeRnB+i
AWrDqmqGgGZ2rB6K9XJuqHfEhQL+Qs+aURLFgV+1LkR/a6dNCOBKVJsinkg/Rqoq
9LRCM3A4GzYpDoZqhGvYf1L6GQZOBYocXavn5vufwX0+1Eojx1dIsJcJeW4g4rSl
3DmGq3IodQLlv7oRHAVGffO3XW7oU2B54m20F575O7Vk8HEWPOCli40m6dX7ViXh
CiUnDiYWcanIM7ZyDPf+an9iP/UCx+xqvoL6BeRIjbyOpldSsthv5jMQdit7bPIz
MUWbHgO638UP1nSkXWxqvA7xSWPhBEwEX/S705h5ygXXrFu0rHqtfquFJddVO0lB
EUSMwUm3rSVk/oZ9CsxjYilJY5meLSttYZyv2e3u9uFctTxLilyLn+Tw4rhgahEX
o4dT0INLyRQeFM9fWSnhn2/hLXlT5ElkokDCX4Y/p3vRGS7qX2XVhUI0YJmh13La
8YRyR/+LdPnMPAJz1orBeHJR88GJl/cXHoewetDdfW2okku03RlzBYEr6FezA5l0
pVZJ6VLaHsFNB1ib2XYCisnLzwteyDmMbSRn7RtTdyelzi8+EHEcd/khUBlLzYxM
IzRfY4S+2u3olS2kY4Uq6HfVkgwCMz2sjsv4EgBBxK//XgZxjR9r9gXFghDTVcCc
Gx0KNmmtw/ev80jAHLsD3eVdSlplRldu+GHy12pW7CT3Tm+7H1Hy9P1Ci7AiCArb
DJPpA7OVde0oEkd5sDMJ1HGIa9hWt1AdPAw7Aglk5UZAm5GfC9mSrPe4VGDdFLuz
zZQbuh/WJL5HsROeonGhxQ2ta7yam/TKpMpzAoqqnwYwvql0sqLmb8oae5fn4r29
5weOXsICIYiJCiyYn1R0PxpH0RqiPhPbCEhiwtpZimHofKqDP8E2TC7ScRMZCYSN
GumiTxv7vEbUrBXvnOWzoGVfOe5QWTR5xysZDpwZxlEu2625GvXFbB0/d/4v96Lu
YQyAR+frxE8yti07QEqMqj4XO5MkRreYEb/urE8aiTKSCBbBLcC26jveep1Kq/Be
Bbr304uXJXAvI5o3w1cuobqJTgHEIclwoBEPAtDphrZFt7PfiMrgHveIVimy8/fl
RFq/5KXxVy6bArbd7thiEO17+snHUbqEkKEeCeM6g2JRFgIqRJUNgdlJJ4dFkS/J
KXrtFJHsQ5hZrx75ToXKwhDsEeryrd//g7D8zDCJ4bTEvTFb60EJvDQ90Abl0Vt0
QHvbW46MgmYVzzQHPFDap1houJx0AruHoH2v3QbKQYh8GXnuJCH5hYN9V0QZ/aLE
DvAAfUxVzGtgoGL8/bMfvrqtGKaJIIFO3J2kcZZ5zsvXJpDZXFjWc1vDTi9NbdJD
65zOBnKzbDWG8CTgG4NqzYXhyF7zJUAB51ZDXvls/cnzfj6VsqHZbzNbrljMZ8Hh
wbJFUkqu+OdAvLFVPCyqNNtpbSs+7E2VisXcjcCNiQLolF3ALhjtUmZlvyVBc+1E
TOGu0+N2W/MMJjejT5zMa2cUoiM2Oe2V0uvcMbCWYi5Uj+Ww+uq7TE8W67yx7nKL
mp+9FrJUb+qvBW4w1cGBdFuTIqxoRS8pZC4+XhDxWS4CTZs0v8v5MWhDvK9d9nTS
oFWGSBYGHYRzJa0mm090YdcJ1oL+sWSQMlrQkyxhf3UkYVQu4evXThDOh2BvVqFd
22u+yydCEVn063Bl18de1qjhksSuHMmGALsVZP9ovmKEgphyNbigQAvMo9bQnU8F
KsKlOjoKPI0Oi5bidO1jEfj/bOivi384Hrid2c0B1qK3/V3lI+6nYrZUi1biX3pU
b8fxzYUZyv4NDLdkbyFO/PtEx1vNzdAONjgiNTf/es3cbcnWWzwflQujr0kH3dbq
vQPiybOrhpZmkiuhwdmUmmvK7ZR2ruPlDEX76jMYugyP64UBY5lKkHvT+y3Cd39E
80KWWx1UWo+hrWsCg8OCGsQk6kmmSZZJBQCz/hoar/YEyUCrowZZ4vgMXlVw4xII
1SvYdQSw+J3A0KHaWxOB3+yGO+HdGwOgHOq3KdyuhseCr74B1Dnw6GloyHjGfDll
QwUfBKW/qvHvqcbudekK6+Rq5f4cKAIDddwLkzCMS7B9dmQno+oABZYDGUo8n4Wj
rSkC567aU58RRyFFVikWFc84GpbJEtVwto/VQC2kIuCz0zTFiL84zWFyhKrKCwCn
S/cj38zsW97Ch7bcnlB4fku0CastTsmCJi81xYBjOkuIzfUH3hHBQuJGh4GfEEOe
7ZKTh3mOZmx3KiLqb9Jrqq16AEwng5Tazk5FS3L+XOg1txJl9YrOyhNSxGnv+S0i
Q6WMiGbv3kjbh/qlWSIrmacHAQ1dUS+0a4ZkViyhkC6rcn0nE6wdkOXvbqmv97NK
7VqlZTIpwYdW2Un97cZ2AXgmzx30RA+G1l+6Il4r05HTAuFlkMv9xrO6PMEAPMEw
8CQyIn9YUgwrsun1Dzf8y/L0O93sQjYYZhjRvpTeJMtLxuQSoBYfK4Mqv0ml1T7e
CmLCqiVLkytvp8IVRQUUoTzt3TUuWrciLnSJ+ubsIZz70Ipnlz5J0DV0zs4XL4v7
NPBzUKY8lp3gKzHXnRiRUTVZo+BL/Z6bC1B19xdPvMYI7m2+i3El7TIs87SacwwH
pGvSLiVwqL1XIYTCZLuWG9i2nyH/Xi9iqX9qovZBNUFZjdJT4UHKRPHL14ZcxfBn
bGls1576xlnTe6Q6mgA6UpzTUBeRJIZgHqOf8LBUwQoZ6SiI5G96cyQooU/58T33
Yrbi2+H9q864ZLPZ4DCDzx3K8Ns5FK1tw7QXnvMsbrH/DSo6FzTSzjAVpx9SIuTt
KrB+zUAlpx7dBU+viAsxmZc2QvOgIGe9L/kxwGsFNjvTtZzCp6/iRr2YTwNFpQc1
VNtPc1L8JChBEt3lYBdHP/Pn9MSMJsj+Mea0iDX3/vnU8uLb3TLTW72/tMnscddm
K1v7JILZIF5L2C6cbMbkhlI/j6UAVZjqaKIdK+28UED7ZdlMSYApzvcVEpxdQfbe
v0TP2ahWy5y6Xj1R7cHoo5yBStUaVg+toreQLbmLqNx+LTH/T0CfGIRevBwoPpOt
8SEX1M02QzSep4VtbrX5N4/yjpt+OnmEWkjOuDDXRvZsrQdGlSwkEHd6J2/fid9G
6Em/gz2NLje8IQBqyo7miFBgdniApa/0f9Bb0A3pGUFemfQZVmgg5NpABedYWAyp
vCFBWZZBP2HN9CeLeXmgRdw0X44UKVLUWnh5f1ijGHT1Gmv/1xyJjL4ddZVy46a1
SVQKdDEwP11VNaQFa1B7bfI0Fg3gu5ZYPvmK0u/rau+FWXjVCdNJqg7xI3QFab52
ftWFPIG1Gbw3KjR6XCZPYpi/rkkrGBhal5bH2w2l9qp+3e6Skb1t6m5BSZtlGgFl
Fbj8BviZZCTGEfuqDqFEl6ZshJIEYIgrNPT10WQrJunJx1oXSgzZ8Txod96ADlPR
NAY86Kzmo4jMCuDto9+tqs2jWXW1cS4eVu60BStU6CtyFDkMqMgbz9E3G5bquh8U
oAP2sVcqSt/GOQB9KKHUsm8xeMfPyapM5cn5F7f+0DOYpdLO6jNzZkfZ819uBlJB
5UDUmJB8xg+MGr4zqvyWwUlmioSAFwhA2lSy68Cnj5TRvMjn2UTmXhWDQuHjvndt
x5+Qheye5UafZEtwNb3T4wrYZMEilLL7YKWz9TLF1iTjPRojoRhKE0vdG2sLh7Q6
bKI6Myl3vh8jjzJ2Qn8/pXCitVd0BVHA2c2j/AtDrZJvyZ1WESd2m6Lxu2kmqh6P
5EdCBJWPEQvftx37aFusmeSmqY9Q+Yx0VdVImGZnPvgXLG/BiTqSJVMQbHCSqBU5
QcnC0CC/x2AXZtPAlOdg40OnebB7zBDZus2qUQiKFfqUMndcGezvDQnYfxL2ZCIj
hfvynMtaTKvKNioJoSNwTkQnp04JvMioXy3fM50v9JIyF4PkDpVoQPV8+/E1HT44
57hxa6sMMJMoieYI2I68HKNy/n1+sqVjiUCcb3rZ4TbWfaDW7z598Eth2vpLT9KK
dFYTb4mTnN5N249uy+N9CMT0D6WwRns8hdMfpCcKKPXT8E1rXMkT4zmgxl2qJp00
Mo5QQ9j8qGZ1ku1vxLewfjuTQVqxJvcAI1qMdG1AZyGqhD7kGOM6PLIQBdmw0XpE
JL53eeTS8PqBb4F2t34+MUufoCD628zYwQhq11zl+mOWGC03q/p9awcXcSQBw1fG
uCFQJrAMNAtI12lFQFlcIsC2hlA0eeoqM7p3R6Qz3Gsq/Omry4CkADlMy9sxtNfY
oO2g1VY7zrN46SF493za3L8RO3KDjl+cFv/5czkX/JVIYaNYekRvcY1LQu5yVWxu
pMsHsk5tsVb9RKQkg5c9FtKolgNhYGBds43nW+KHr4Gh8m7NrBx/GFb0dfIdKufL
syif9o3Ek5iOqw/xEe6aX63JrSzs920I9E2DZLtmRv8lzRzUlaK0K/YWJhl8H+l4
k/ePCxEChWhBTXdpW4iK6QVwsPyWJTJrV7meimIdV2vmkOZh2c6kmWB6onvyAQLT
SF3oGK2O6l3JQSEsT8n5aHfDv/HvCtMhHye28KjsFdmzpvUt1DkUcjyrOAlhrRIh
N0rlUV6/yvhT2AjeRff1SyyUEHSUkPDf3BB4jtoxrm3O8y+XR1bVAMTbbny3vEK3
FndN4AtUAFbbIK9j635LJdlrtOZokqQdJ0cyHP/N1eFYpAq5WN2k/ZOGyz9uyd8W
PvYiN43yICpxK9qJzR4ecjVuy2u0r2eB++qUfmpNU/ixDbMLnA86ZVxAWrM417PT
0BCdlA4yDhSkIVo27dc2c6DbCBvHYn0khSmj+CN8780BhmrAyMNWYIjCUlod9q0V
Sb1v7PXlWWZ0hguJYKS/8l9FbEnmfxRkVQXe0p9T4g9vRKSz/pqocs67CdAX1IbJ
r1aMEjLGveDLHU0Lj5l/FUYjDSDipZ3sjsmtLtdue+FvouihKBrJ/hCG8UPg01pB
IOnUqvw1rhEsyowzYEvBXfkYDyvpRZqnwExAEJbmuaYnnyAWoAWlDr9bwbzhHhcC
/pxl7D/Sz+p6NJF85/vdUHSt4Izji+ftCb048EzT0/mz6KxKaOnZvug3TafJI4/S
8W+9X6eps0tyeLMgQbKIU/BaxbKj3YjkNvwRDmiAN7oVtBO3pNM8a8EZ5QPLnAo3
m96dDA5TY2M1d4rkKm+qiWyD7PzZL87Fse1tznGW8XsceuvCBB+GjlNi3Xq1t9Yr
eHbZUpZZCcmDVhhJjBUmwaf1gvbjEEvIVASTmJTDnJ3eyoZHMlKWIqUP1TmbfI5E
zrLeepazBQKGWSXKBrT8jcHSFD4iKk0BrRsfj20A84V3US/DcBYFouZ1g9Og3GM1
srBXPuha5WlmJXGG/qFEk12Kv4IzIZzJhEihGvfk8ZByf/ZaXgHXzPSUJGi70ynt
4n+tAOoUGy0EiaC/LxUt//hbKczaxkXpzcqX9KkeqfCF4yR6ANfccwXrF6U3deKO
zHkl1n/a7p0kbBZFqaPMT1GcKMmxpKlBsaw4lpXe6fFwdfU4fTgWdUAx7j9wFcSi
xDye9/DXTXZrzWQgeo2iVtes5wRSOFfyGfTiCC0iBd4vW/utp0FtO3RdMRCkuuoo
QBM+HjH+O6RobR8kmC8AVzasLpEkjvQ7YkgoWO/Cpc0qYoE60BI1FvtYCnF/17lB
OKSvrYlMRq2Vl9x5/DtguH57lExo4CGWDMxhF5YkD2eyI6ZITN0QNWaoSEgpgKbk
UBpRaa2TieSelRDxiqmEMn1IMIFgSPJ6XUYcChgU4UIQKkJ6sJrhUlf2At0/6toM
V5Qhy3tiQa5hMcSEwg6mjVXcLW7yjUNOzc4HkAdfpu2WsPoL6LVvZjUA+D7YoCnE
3vWZX2KOUpoI2pyDPyG+QxOmTMqEKyS7SoLsrn2/ncTkRJSMUQwHEGdByjVNWJPT
XocAhDMWVoWbhT+zzc+VOodvBRpDLvDur05djNI8ZgYymZmeX1vG+9lp6NRZPKKC
KxZCbrXnYk+B4d6fwr26mEEsASfc/9bGDh1KXq3k9h0xB7DadszdmLuzSSeWibTC
30NJhkCKxdVyL0+uH02mr+SiaNPXZHMMXhHOZhgPvW4PsR02JLhsEkQkY4B1PAUZ
RWceZW2lS5Nj+CqXBoamEGFk8OsxXmiYMTMla6KkRLn9jBrXDx6Ig8UH+7rzb6XH
+BoSc5ZrgtZpPtpqMCXklr0KR9R7f66mi2f0w531W7tcrg0gLHV8xy6vK7tU1zPQ
969jQAvEC231fuYoE9ZqCxqE7FkWS/myPIyDG1Yi097jQmX0pkLpbdSK8goQpJyV
p+K6zhFCy8ou+dYtazDQPHG4Z0nS0Xkxwedo2Ir3ei1GwBDpP0dhFS2gCFf3jdJh
w2cp7WZkq9WlAJHAkBetVPXPi8IqU/8xrIAO0OGLWle5rFst5V0dMzemgDLbO+C5
yBgEj82ziz/dKfEDRWtiMCo/OTouwiwAQj3h1O/XdWHZk19ZZzIJPnt4//clb62Z
cvzvV7jfqc0R+P50+5H2HI5pB8NKESErIwqTCPuudhB+fDhcb/3P2DSEjcdm2jBq
D0feaTunL5DqUrRKaUN2sLkEiFppiOTnKVdud/g84RQzo20vFVw44ajnjec7wB35
Uk0CmWosRastHFChuof9eF9vSUpihYKqfPHVViuEDy5Y/hAt4V9PLUgfip16zRHo
iYXpR6zAxo6okd25amm/AmQx9wGBbtTN1vvro8b9/JqdLwQorode4gMEPBY78F4f
qMlBk0xPP2j7zi2sKJbwN/+wUpPf9l7DPc1+YeCfbZmI0Z/ANjRR5K8tVzEK8G0M
4OOGwvfSiR59MhtnVnUG/oWYSpqFDDeMHJnjunFaY8nMDzAgA6A2W1B09VxPCopn
99uWeUjPGKAqNReQjLimcpJd3jCsLRZaCyAO/fv1FSTN3t2cdyHSBboDvYdZo8Rn
ndI7VQTA1WI7t38f78J1JaPPVCxOQdwhUWM+joV0+jTKZ+LIg/10bo82PDQtmxJZ
rzu9RO+GfiEYsJOsTMv04ySndU/aVwd8CJ8A9BZxhEOgFQhj2/SZwGPHSQttAXRk
VLSDYzjV8S2y2ngdh9ZXL3ZYabCZmhhSZbd4vUSnNMrP10abZTYS8WTP+pWonAVl
U0kz6aV+OiYuVPTduU0iIBF5hT7jzkwRcQIxtWZW7w3frojTIgjBPvjykuoTpi9X
Gkj/DAEzbrQjUV4n0AqUncEIFt6CVwTA21qWiT1LIhMUAKJjweOJHc2wU6G/3E1c
/L3hO3ffQFl52UQZVwJHa05FdmhXl20UYxX4Axn8mtiEn2l0MSCaRD3EBSFr60UZ
pLvhdqnj5phcPD+9oeASxFrG+wS4XbXiL3X2ses8QTYmFTL1PA2t5M8/FAjyn016
ThUkSzxR49DtE78zRn8KdR7nJOhq5Gx7mER253UaNmeoYtGRadZcKc1bPOu1yz6I
c0mm7Nfo91W7NdzInA4j4YbmtCxwjB7v3J/OrsCpGwvUKwOr12sBvbXZq+hzPHU6
P1bnH/8mkCMpGy4Tfoy6ltb/vRjaxv8jO/Cnu9cqKGqffZiTveW0fThpbpGWTJAy
auFuFYF2LU4SbwRLb6W1Ddcc7ykqLtndUBAc63o4ka9FpYat3ig3lMYDCB3awdOL
xAcH5Sko55U8dNViST18yWrr43WtavaBFnP4BZ9n8402OPjs9PTzTFedyjl3rgT2
GSatOqOMmCeLfOPNV/p21PXbNDF9Wr8fiX/d2FfBvBcDRaJIH+7Fk3GmLTzuYMVi
LoNbwzWaz2axPJBdplOmyUApft0rHF42b4cqsUkmn/nOzljoNCXcXGoYO13AKRRB
U0o20EgJ/Apnw/1mmRQsa+0C6X3paPWfU1Dq9rN74k3bQwi8ahIJhpicSNG9osm3
qJq/M6f2PmoWdDckCOAN530/N00L7mvpj78ZDC3jN0tIrnB3pSgq8wMHNAdORWzn
JbEWzOE1bX+3j6va1ys3J9pHYhnUraHHEamIqIWBfajLrpJTgyPm4myP6vraye3k
5bbN2D/+Ia12nIRBbxYnLfy+bfxB8F9CicyQHpOWl1zHKYFqEtYjpXXg5ftu39vo
kBsVf7pxg2mls7P+hii5iDCRn62HG33E4p40BIVjvLk4kPe1/yPag3WAXwbPYdEY
Ria60uhKmkQZ5Ld3nPx6Te5cmpgs6x247DvuYfocPMlkzcBH0QCYbBYYYV+DVyuk
44F1QKGtu4xnttjb5s9lC+KRJIjNbLTn3DSiw6d7HeFbTPocOZrOPtM+VT51MM7+
8bGtA3qNwGQaRQK1DzBEEuBOioGQmEVEXay9ypvBY3sUD2Ne0orRupS6xuSmCshq
X61hEffvoXOQ8jLViEustl3Fv/mAAJrYaZpE8XQnzAFOo0YJZQ93rvgOqZH2flp3
5/Sb8rRNsW5WWwZYBtLDiYJjE1wdKc6cJrhD+y4nRTmoxmA5sR1DDsD+G7jw5h4G
HRx8hu4TGDocuEPPdlMbEzUACrBrBc44NU97aaOnoqjLvPfpTAw6S7VJbf1Z2sUL
KaQ1/AgXC8mxuSLuM5l9gKEeVviB9SCMSlSpqg5uUraA2qlhR2XZ3T++L9WzV3fO
ozdyRuUA0Lb4UNCZa6hXG9YdU6gOfv3M41rTZ96eePaaoO7Sv1mAuIU335hawzyO
sBQwNCoBXS7Bk2hlO8gZHPfGmqLnWS0Yhbteg35u+n4ZagMFBpDoqrwe+vB2sVVU
Xa46Ezl9kf6QiayNlGb6pxa3Qd4VXSweSZVyDVMwBG6bU/PThR9u86LngA6id588
aw1GVMMUKf0uRCsxh6dBkhIxeyFtkAYf4NrbSGHbw/AuZyU7gnn7x0217e3SALa2
Sngo6HSsLq6yg2zf5MapYBbyOCj5ynVl2i6BNHgiO1nC+mr36yRxzkdpXYPVsjhx
w8wUQlhLeQqjktx6u4lctdXoVzDqyl/AN8Q8A5nu14xIieyD2Ise46cL3Gb/gPMA
cQeN7EvHoMvQGcw3MHtdts/lYhPF7ouIp9PDVbJnPQGpV41WFL17CQyF/b8M7wbW
CfcYpoY4iADM1Pt2mAyopGPYRpypuGOwPWkQZQHmfGeyVgjvIND259lqMo/UFLbz
0JWhZtFVGhoX6dDuROKDhsNVmxHqFqgYasirXXF9t6IXxMg2EexdwZy1tfdaVuQE
GYO7xQLUJg/apgTNSvnUK1RDwnmi7N2SMvLU0J8XpI/6xrHmLqYq6dKMQtt0q819
9bT7cRLmvCH7ioypv3RYKr7O2K8ngFR1B9X5mcqN4hA3VgFxtTYe6pssMQFlmZso
8xG9OZo7PiSO66zTdHZV2LcNuI3uLMUtJLLsNFNH4+SCGeBFNVt+FYcaH+fKn+ir
wiHEoFeOvy4wmdm1YdC6k4L+s43eSZSw95MBSVdsh93DGvZsjiNg1YZ16JNZqSjD
BZG/hYsjIQMZG4oVo5wJd7a70NcY2hKy9ybcwET+6dav9pCP8L7Lkj2tqng/vLGm
acHBsAcSnZKCY4d/R51JpiVX1YHT+nCHXeJmX2i+KpPkLJJCdrz1hHRyrb5woSkH
/YzUFjxcJJM4jwUEf5E+ILQCtNCna93o7AiINu73F71xNKQLE9D0c1uX6vvoBwhj
G6cTaTzanQhqlK5ySct9Scp3OsSGHehUYK6Umfmom3mP2poCP9RlEc1JpWNBDFto
YBv2IYyBUdwKKT5XESvDktJWw/0mz7rgmOwe5bjL+7VsxjgRkCrUEm/Gy0zwCmdK
8TLAbHhr3HAf354J9SN1q+Z7enFttseSwFiawNk7GtScPdMidGb+hsFQwfL1kqtJ
Bo4TTA6lQhj3XPoqasZ5XRrQ44EcQZRSS1R9ShNjgiVnfdUndd1m4SXwqiB5L7jW
yheeFlkZNyTAA0wVcgQMT1a4uONIaAZPEJC5obrNPmoSsosTMUtkcujQzJco+Hwb
5rVD+r0mRD0uAKCrAbvvuPf8Q19XAJbeq+/xmugiNJ800P651m2T/jcL/7mFeoKt
3HpYbPT4WNGFLziY9NUtVl30BXE+umb2MqMMqj+rZDhlIl6uTMLwV2nTHTVCIkl9
1mUelhW8TarOkciukqhPTeuPmN+8IzI8MtRLLA4tkIL4J0DdFYvO5UWyl9tpNfW5
t4vyiuvhm3QE7SeXrCoI0W9VEhATvGcueL+QETcKVhPw6s9IKHCEqXF5O7zYJSf5
nrh+UPB8t+1AiXFwk1ZDHoaEKWrdWranK64bp77bWRATqT8qDcHlSDITPdiAKRdy
Fwks2Oppq4quyl7R9aqJ2hlNo5bHWx8zqG8uMeFOSqiAAfbDQTgsi48iMqv1nQR1
RTy5k9KLrYiowHWPdJgQXzOFcflumu9JF7orNXzuKrCNWgHEdwDKYPkxSr/s7X1R
StSJRJEAEeIXGaL7IdrZjjBB1sTNdMaWDEad95zgAJiEJTEuRbZdOpvFVFvbA6Yr
o0h60+gN7vtgcUZ2XDIyG8Kg9S89l42L+rlnXlA1uWBwtN7wUgINqG3KVWclLULs
8A3QEcPiha8h0rwhpcWQuJhnCxwc9WhMuPUhU660F7vkkbsGBm2k7Wg38FEb/RTC
wyM+Kc4quNFXFD4VN6GZC4d6/r88Cr6FO+/m0Qfst5Lz2gFVOSXjfSWY+LErwYjj
Qt6l9s2WoZSmRaBUmdyJYOsOj5gNJsQu3VYz6x31epohZxEB+yApFCTMHsIAJ/S/
FlskiVasJDcXzb1AbUoJ1stpQi5UsnMl/4OWMeaHaeg2qXVo6ht2PzaQfKRw5sWO
pp2F4iHWgbIGSyHU+EjHvh+l1KEASozfnaz57OyBWVpGzzGm+IWAE32dSUs1gju3
Iqri6I26p5FKfc47DuJ2bz6Mynv6AVgBtze+0ym85lpXPRF9aBfMdHWLd5wcV6NH
ShCZmrLDhMuXlPFDf1J9M21fmhsNni/XwlZNC9zOfzGUm0Jd5I3mL09WqUEI7SAg
AABapNewfekPDrYgDyAsPOF/EqHMB24XnrUGaEKd2a0eBFYeePg1hwlqvRCT3dqn
Pgap/3pvzQhWga964foKKazWalagODz7vrYhhook6pVprmkvR6twlZ3Z8z2YVceU
1UdE+f9onn64pGiKBpFIVeVeQhLVi9aRAVlEtTfxNhYE9Fj7n+x0JDbzbq7oE+eh
c++w3EjbBORXpPIYn+dIvtlIqUCTITHbZqqkB0EbApExmTgz5gpoR9yXHRO/wceI
Y7oCNOWm0twdyD3xmqESZZrRVnlfYhUflRcR3aWe4rDIZ7fBuMY3USex7SJ2Ehi0
8wGmVd8FbAE2L2mwbhwBBIDjMEpZJ2ybXM2tE7pigKzC5A7aKAV9GsOMp0YBj0K3
STfK+uQwhQFK3JgQ6feS4Wz6IDP5hnF8n99Q9QJDFBjiYuihLXiMHFzI5f1RPxow
ZHj8cf1RvU5NsgVIqrR4pJK86RFtjhhoNzXlBY37LETFupUpa0fkAT1tUlu1wXGO
yZ3h2Zw60V3xZMXviKKdx7YNvc7hLQpRzqdv7IZb9DuxT7eqSxxmRdjU+SJP5MJ/
iRosIVvGQunmiRGOIOOfRg8tauNbwsp1am0a8qXQKn+YOybdByjybN0KL0dZvYJj
wqON+LuwX4aM5nclvMQA0eYGhvDNv3JPBgvk7OzG0ecti1oAva9iHkCp4nwGdjDS
BxLkrCkmHrPrpCR35xqOBAWJ0PIeo7wJeXKhojuSN3WY7lUFDw+qGmgL5rGk6Uci
1/LWbi1rP9WuAt7qS76iCrpaicQhf4Zqgm+fzBvbmAumI9uayepLY+SF0Irc/n/b
R1//KR6h2mpdEVrfwDBpg3PTPNSyR/3XQsyr5sTpHbvQ8tDUGxyw1qEY487K4sjH
KKilPZw1HEcmm/3swCgJEp2Z1wvzAznplA23tBR6h9m9RtAHuWylA4FiJUx0BDBd
beH7veA0W2MmIm45YXmIMBJ8Qp/dw0c6P5SlWc+Beq66FVltWUSgiteTgDa3cT/i
pPlB42mJqYh4gkj0KxvUeh1mfNVNpkdF1kfef2m1QMlhtzJTfMNvJsXyhpk7bCCd
VYeo1sHbqQWy2an8sqmVDXE0gysjBcTTnIL1pTFSydyH4H+ImiLiuinX1VLCz9eP
Wf8Nd7UYWxguv2Y6NcgOS9QrbiMXKgHBn6SLTJAuEz6VAq9nK1d5T7zFmufdat7F
L96xGdGrqCem1eEukxg47HpJMH/wtKmmpQrx2jgbiBTk66IJTQeABBfZWKwIj9Rf
s6X88kCToQjTcvUUIh7Twdyql42Gi6vxyw943haN0J9i+r1fPWJ2QyVxaz/ovtEf
LqDmd+m82G6Uje3/dudmTn596j7YW6MIIJF+r/lBHlESM4Gn5mwFeYQnDl8AsfWT
/W2p6O3OSSUAlF87GrK9avCbOy8vrCJe3Wf9u/Kr2P2MmnTCwZ+NySWCEUL2FzNZ
5c2dgweuQdjoJG0V9nQEEIqKTKjnzkcGKeFSlRWqQlzd6ptNZK6dHsi06rs6wLBU
RcqDSmvT8d1IKWTjgaTx7FypInUeG0Bo+AHlYut99n9xMt3sdYemdUPEUYMgXMmb
yzJQXrggqog3VnCXt+eTc2pwNMD3k+8hPbPjPxsI7FFScOVwGBYyChnD5qDEJRrZ
wmMNjIDK1fQGVX3kg/RoPARsIn5AcTUNbyi9osjVbwM6w5sAjwsc7XSCZwJrmPaa
yDd49iOcBSCHq4YZRZVXd+Rx5UIqQRdJmnM3hlODzdzuwUdgENib+J+i0PD8wWeh
/XcPX0sJguFtgDdAK8aXJPgf7JcLBmKJ1Y2xrSaqjG0knrQniWa52EPS/Mk0prdI
m/U10JUFjazUEUBWJAzuhv7TW1ESk5lwHKqS4xtmpBFk3dTxbCkjLUgk+MbpQaPv
1CqleBW16gy9ChCis9VMxhj9MkxjqJKNtKXAwE2YymwKKrUbGVG1kQjpTJ8mSf8i
Z8yGmBONyatIMA+nkSNqH+am4j1u8mucMlK+IfiKl/7ujFz4xQvagJezop3eEkKG
E0e8A9dVDuSS/R2ufa1JqNJju4fuIxUdUHd8vO/QxbnOg//w7JAdswkShCjzosNt
i4Iuvo+rZWTv2L1k8j9N+ldKZM7C95pgOU74oKSSGvk2pZjQ3CVHVAd6f3nRKjjR
rP6myQuxo4KjaztE1KTGaD03wN2TEQAl0Z7cKKZUoa5JfRcpgXDjAAm9ItCjh2sY
B4tyMKLESQfEAtbYj2P/E1K0QwAuN6/pP3rEQkTivrWv/jy94l9Lxh+ccDBUp19F
ksMP3BoWElR1454k5IbdRV40O414glOjyJ+jypHyT78EM6kCR2XX/ulzJUYV/6oO
3+yTZwaj+o7QrjewG/glmIXItSd7bWuUBc8RkIpX/9i0E1jM3VgbQKH2lslq2AE7
9BsCdA4EnD4wq1nGV87EHoPftMq9a7e5IHFHUZBphmI1qt2Zi+cvksNkid5OyywM
m7n4fIjHVm/SK4Ogwx91+jA56ezglcutCbg4d1pLjFHiw1WtmOb8z9SmuvQgZ3Ro
G953rLymrihJHJZc/SoOyZL11nrpF+wMpAKEY4/SBRt9pVYbjiB3S9QpCTuoTqnf
ViFJZ+sbs5q2UADi2tgFia42nZw5R+CX2L3bYbkG6iEX2RkY5o4ChAz8LJCFXiPS
fJpVfGElkQ5Lg24TOmtks+wCYeEL7wh0NBRgB+z4eAV47935PdlhdfYvcjYmdaVz
neDC0K1XDA5HWzvqoM9445Kd1lUGeeaJblg0gvEpHPzp84qwkmahyzki3lpw6ACx
7Yb/1Vh0SY137wgPIZGTz2PPXa9jwVbL1gNTof6bcdpn/KKKFz6DBjSaIfshA/Ac
QDj8ZX+r9eLw7RAMHQ4dFg/bAOcF/DbLOKrbKahIapmw3cEG+kt9IbSXNBx3bExx
IA1r8ih3HmxovLkxSb93wxMyhP9Wq4T/nGKSFC48PtpD7vxAXDQuFphAqH9kd474
VuPS5YUEkby3FHmoqK3NCGj4kkbDNkHmla5eh5qK8tEzIrDlsWa6pHoZ3v5XyE7n
nmZdeX134PuMh8lH3akW3WFWruuJbFKJAj5EcaQ58RjBYaYh3Xro57nP4AqCCrPv
qpwE9OP48IIrsxm87ms5aWccsdTLXDQUm3srQrGUaWUQrYOEIQMcV5h7QY/i30AV
0MTPD/Hr/jwvi5DXkutmbmPyxSn7mXER7hPh+TP7cPvqPFnB/TyRfLslLUy7CVlH
HWuxi5x4R/PlLuzsSu7m6iElz2xUb+fA5mY/Nl0f+DtI59Vi4H4e9JYVNj8Of5Jg
p5wvHlrc12PBfHtW2oPmpyBV3OoIDRHHq+bpeJ5WKkMTU7Xs9hkbDkyGp5qShGCQ
Gis2SaYThy5cTqi99kjVikUzclCEWWKulFVYv7J0iIoT6St2Pfce4MTxw2PBSepH
U34zgsWg6PuX+zzSYuP58s6iq0WAU7u9gka6nLFGgESThT95TDrDnJfYa4pUpboa
mrCPmb843eo3GOgXWZJDqIIyhySD1L8x+lBbYhqcVrKep0QRlsJ+Tnuk/iGkOgML
YSWxH5GFo+Udaopbk545VkxtNRN/3KKDuhV+GHfJPkMgDpTc7EQeMGNOOs/NSnru
H2oWecYWVT3YoqyrhWumBdOSlRJrhuZL28Nuox3NBN2sa7Fstf+/6PVMrMws+Ff9
n0zXYny0yghornScQV9SKHTHjcAxUgFsn62kJgwjvtKblrZ0m+Jh9V/PKKpL23jW
4pLFZQnVsIpfnDRCOYT+ZTbEO+Lh7vkAORt/etgwOGskwAj/2xx1bJzTau650flr
/tQFND9kem4mD4MeBT3YFl6Ym+nmSlBeGRw31lv135L/o7j8k+W407lph7+9p8g2
sBmAIYfj4IOdP7boLgvkkdIUfIM1WI0XGJU1Ha0JQtaReUuEhtbxLqcsAsaeDOiv
lGzkPXJ3bUPDxfjjgYxKFuVpf0/PpP+wgWNK+0QkTh9Y2b4q0w9TsRrjdoR7Arch
Y/0G6UPWIUFIC8EhyotdpkYeD9+r8eSHKfTBHxit4al9JfRwBFJ8XdY6tIEkHwBA
mwvhYztovtMY7+/5S3zb5bodX2jUUl4+94anWlKxm15Zm3Wb4myX2J4mGJMV/qFg
SeLXfed+nZikbH1c0QVEbXjVpIiEZKsCoAAj0sas2Q1cAOgThnKGwvQwCZn1S3Fh
7EaO68BzRJ0cq0TdYj0WgJS9vgNLBRXPCQM+lqxMfpIqYDrL1udlOiDG5hAR7dLI
6FuvR/HuRwzfc/NTNnvYQS3XAQtT5XBhyF0jr8C8rt1ZBGaYUwuaUyGeXHD1L2od
X3ygX0el9HH1SYN1eBsF4/Q+h9gy4KnRGKoWGxjxro87vaDSU6FQU/hRhYEMCqu7
d9nZrWi1voRiBOnjqRae0DPHLhQiZQpiD5WJS/xdmWC0vbGjqVojGLK19geNEqEm
HjOzJDdMnansT/0+o5E5vCiOQz77wMDWj4bX8PG4MJa5hV7xVZxkeJdrokf2LN8A
hiL8lyppJoQT9Ws6L3yXPEnUaS5r5EICuyxM2YFn373LX2EGKr7W4wkqzVIcaBTV
WuBgsBJCc2iv6DKy/9umw93Iy5fcTSQoAR8mv4Ciwfpr6SorVmH7OBdcy3dCh7Er
WC9YUyBn46ZQKk5WmMOCyDr/9tlo4n71Bx4AQWLU+iemr/DW/cgcrMniHqqwk73u
NfdAPXUn6+5uI7TkAIEXNfL2zxupSb7RC5q3n3Un1JOBb6QtWsRtB48ipHagK/em
N3j9xk1ZG+iLg29nKWkmwTdb4EuBhW2gjjLA9vVpVhilhaYSm37w4jHdXjiShjW0
DULldqcdWx15W1UpWocpzuvi2st8ufkR5SWs5zdXrH6BWX3KTZQ8+JafGyPIUHpG
kZxwXlgPz1ZVxT84d/j4iVo2eXtHKJH7ZDdX290k2X24bEt5aygIKRsF0kbES/Nk
4cxmP0zZZMQMzu2MbuqxJ1cwkNCCdAhqQSR0kf4TrkEdv9oeTXewF7+3njyLWGJI
mu9l+YlxXL6vg29lR3yFKu1UdqNKxwl/yU6pROMQBCr6xPTdFQdM6+mPFgkUY3rO
gxodo2hBo6u6Zq4+mshdmSZ+vibXvVnum7fylJw2TcJWu0db7e0ECvpXOs49JJsS
Jmzv3NHbsIpOFkgpFHqLTr+rcWlvYrLj0F8mXiu6ZFjf0Q1GTnODsayfWYcXeuty
F6A5Dg1DjzzGEHohlhx8WWb5N4V1+58h29d8KF/aip4gg220x3Cs71vGqaghUpgN
GL1fUJyTQRYg2qWKVMQCpGZF88an4RCzFBZQxCzAVfkH5zyvgxaoW4e+0jWPfpED
9pN1N3lJsPZlqPJ/JowJ+HhbhOjuzRbwHuEfImfJ6EJvzD6Knn3Zt+bXMTCDhJ8s
vmcpAmh4iIg/bKCK6eyMuqgUn/VHtJmsNnjdHRSKK/70vBo0g+HQNo18tiUx+5KA
i2vi4Ci2JBMSyGD+lnCk1VSHlQPAhlsBkrr7meoS+83mVqCod6O0zkHHk8XYF2AD
2ohtRkdyzmFSLCt7QQJ+1/SPOSq8dRKw2eyD4YCfr8G2ip6A5vvlJ4cWYT9j7eIs
IoOrtXrYI3RThLJZmsm+bBrQ/Qrcb/4nARGaXfxTT0tpuVDx9NdZegrIv6k6BGKF
uQk3VcfpI16Dhbqe0jWsQ3YIxFojwkBkICW/z3Vxn3SQ+ma/jqVzwAypP/JwYIjo
UFkb9xB9iLgkREJXQgfjamOChcbepnoR3bxDWdvyaWh6s1OnltV276rYppQpu5Wa
fqSMfzqsGTEwxPn9m0GZEBeba6lfVfnVgZlMLDpxVW6cymY79ieUNXmlYriUqnjH
2DgjNp0o1pIbd85XHF6UsHwYtbIhDu04xrxsSuPdBo0Yv1fnqU5LG8iSgsWjFGuu
HUOPn0Cgn2xSwSkV5QrVZiic9ABHKak39g3TcmWi8QE3b6ZYKQwcAR0KRYXgx1TA
nqRaywANfjgAUGOErpb5Ks9p55i1rZQaBwl51brtcPc84LmQUrofcSqKs7qp6iLC
yqZPFQCUuhnhKJAXcNE5rTvFVZ8CN4BcIPFKCT3PSPRiQhu1dqGlO9/T/nPNUR04
ZC7KIrraaY2+CbM84BD5ujoHWnEm185tOq+TZIy9b6f2q6Li5tWizJiezdFuJVuj
qgtcvJ5VqmOZ6LyG8aIFSltxoediEH7OV/CMJAkRFBu7QkZFpB210tMbcca4yWyS
Tw7Qh2+WferX7hehNi2EeeQzMgc0TIB92j8jTDw6pK09Q4NQE1OO2T+VeBDbbJDu
/40lYCtElEbwaBJ/wuwSD6G/xcd4UxHgk48h3eCca3Ys9WEi/HqAa5ulKxZmIBTo
iLmAsLyuQgQXB3ObcgCYSP8ig1aLiKP8bkd1nmfKZ6G2BLCEY3p94T4e5ZoxLuGf
rwzFv2QuxsTaqVyoMxb02t2hGnvpomGWVMU5txpQ8hcMPxBeU+KlAs3z3BAgej+i
lrntqBw0gPEz8o6GI+DuwvUe65pOAqxRqv5Y0o1RFhw62b76XxnVQgupmclTbe8j
k6nALOdgJAtWcv5pXxS4tVS5d7zkYDcUdu3h6lcSD9DV6wg0S9HfUxFDw9ciweRD
Kg7UqCPjH9qOpSoLe0ELPo71IlnsbbL8byFm2sVa948YZNgKVbmdMjqVeGnM+rqY
GaBXA38COxxLMz3XlqicNztUVngk24HoGk1GDX7ZviHs4LPznwBa8cUH3ehxDCRQ
ExdupFQmIm03zaOKo4WJ8x6K8WTByNM40/I0PAiUctyAFpctR68YzaN3iNiXIMgf
uef1AUxo9Kmby9O3I8n+2xbUo2D+5VeiYDHBiq2nWF7FbOEfDRj4YsVmAnKBJFRL
JhcO99ocJNMY6nqUf1UAYk/KmmiPat4WSVzFD/wbIDlLxh108SKnpup//lROJIK1
XbVOy3zZSMpOAVwhttqaXoQy3eWii4lPI8OfwO/ZfuiMwsv9a3N1ayQFNQuSNl+d
r3lE00U1UOz6oFcQBEwPRiL7JQCYSfZrXTXeBhq5vxzXgqH1nHPBwoq8h9adE4Cy
o5MicTu6OE9ulQCqZCetlUlAiUpfrJI+oU3i/SF+/6X2QXkAX5Y0KgvdzfGwHDwt
wVzXrfWGzl1H8+euKT7StPWZEKDeCPGMw8LhsnnFvm51gMrQMyZw/ydad4DtyylG
9lK+z4aIU1BO4g2rRSJIQw+Lof3yRGkZJKKF0ZQdVekhSoZmf5HerO9USr2pMrfk
BCM+LISq5aJiMUMBocQ+3Fap8ILurlw5794Fou0H2O3qP2Pg2EECh+NK00j+G0uw
GYOWuEEO8tYQA4jhfjpaLgJV9rPC2FqjA/jebhbvyt5tR2Ye7RdN9v4l4XZB6ibx
51aMPN6X2IqXGNldsTGbvOUwads6Gi+6MPzhtCUQmfNijHexMXvcYDgSYY8ENp99
2vopPlQTMT0E/WSRXygylDmMsicGznCXY+p+wz3yrCQpLqiupeBwrKZZtKi7xNzV
be9tGvmpVB6MbjGwP1XkZuCZfG3ifAsQJxL5dthBYRQpMeSbMDnJ6MnRVW39JrWR
jN151Q3yb9a8N098KvTgAm44NiG+JaUZHao6GdA9Wxxs9tx+QttWkD2mhR34BlgF
IldkdZNi4worPUhobbNIsE8RCubhLASsYxrNNP4i4EVf0LPi/nHyLTW0mRbdHtFY
SboQIyAqBk4RWu7tHu0NtczXoM+XMFq4OGK6TtegwLGM34fXbiC1sKyRY2D4qNA8
uZDc9qWPi+2Ekw0ctBZVFtEoolncw7mbsjMeq8u5hiHFvVNWGVjrRYuvtSMvaiUn
vNEkb1HsT95D53Cm1qdGTdnG3vQ8/klmpvq7xXSJVkcvJtcfptcUJ+cBkc8/GgNH
e987VmYumdD8PkqJgNp/9IW+o4DItB8bC3Eodct8b9QkxF+CLrOltyv8yhkQwvcB
HbZeiRkN//cRZTPAY5vCWpxXxabU3Ap+SUkT6/3R3B9vTWH5R5Z8jDpgrPBsjQ4U
O9PEuwBucom1Dxl4igUhiT/9qgcuVWE4zJkuN5xKOjfcw9E1ZsDqwI5kgMWoaD+r
zPe6GOyo+nL53+p4SmrDFhoWkzx6xPXKlDfuPihJugkkjSx42PoQG66xXvx0lwlo
gtP/lGcP5xSU+nn1vUw71EHg8KCRaXezTnzcP4yq7vLkVhV28VmGJKOxaeyz08w+
R2+do83bSPFqGWhQcTnvBUO4T42OfaK6ei2AmelzSrzjZeJTHjsXKs+CUap160ug
5SphojJ9YYCUw7w+GDvdbtdQv+98AvFYfVSzl7u+Z3JSS303y2hQeYqrzz0pcglr
NzI1y8DwufQLdmUiMnIr7jydObcHYCu7jgtvFGJpfg6Bfb7YLtpbebv8Evjk+k6m
yYJqnm8p+LLpkXcKc2ayd8+ZnKROFzm5JGDgO5C5afaieS6w4RYLYn7ZVJz773gh
jk8oROZDe2o6P+dEKADtMFZoqld7E0Rxa3zUxDj34su4d5Wai5Gj3g7oC639PQGe
D2xJ1WMJ8+z8sabbm2Q1nkHQwASKwLRM/3csTWbEFuXDKl70uz8hEJc6UK4IKp2K
szC+0vpFZ26iab0XnLDQ67J15NtufSzh0DglA2cFl1DIWHKmOWNhRC+lSsxojKGy
z58AXmLYyWZxaXeMCDxqXrLQCyhlNV9HUn4BfLG0jlXmtbWP2Gy/heQGXs80l4GE
mZiXTFKL+VHbWLHMe8kHRQvnKqwgWxeCzMZfKMkWVzdgU5X4cbZdUJRYb9T1BLGa
fILEj64yoKpI0QqyD9cSNrsoO94QxW2piDMri1uOUM0r1rozSS5Oc/FnGnxu8506
4jcltvzbTfj2ZAF3SXJOwbMItpY39FeIhOigUOJ9BiKzqZYsmVbEeX/fVMTa3oQx
Qw1VSIsIavvTDCmWa2qSm46YFUwb1xenNrzMHwqSFmhawYpcPXAOCWqL6g0uOwiq
EWGd0stLrGbY6LQgHW9RDgaePlYDIflTw7eTvweoqqEB6NnUHfK+6uv2XOWS3ziQ
DpZdepAF2uCiiYtGI6xb0xgEVgSs9hv/w3pJUW2gRM8eIn+ZakRcVsgnYmJaONZ8
gC1ypiBLzuWMeLZUjgYiE3C2c4sxZeKmmdGWo7UPiEskbuqowlKsmpSnqUsiIdmg
LE3NAkQQCjKGPF1vgZPTX0PTR9Xtgr44FMC5YujvjATVAgwOnee2g4f2V8GRG8+R
UCLqVwgq7g/b7BABgpKbkMgSQu+8T+qTfXYNFtB5Ls05bZNUvB9fwLy3+eiGSjxS
Do6ZTQg9iz8xOrnrJr/QF1ymetX/Jgi42S78QZvp1pN3Tg5IFn2Z88ua65Ot4JkH
802gBlMt9JSz/3PX4mKV01IwgnCfwvhhswHteo7/LkCf/HHZSc8fdAGSje7V50c7
+5ltJ1Bj/SISh90ydabLfm/DDnLJp/aIcgn16GrMu52BdLcPoCVoc9InIs0F3qCR
XYg9BD42lK+BBv4/eN1ufjhTsGIzkZwJ1jljdZzlwlmy/LgqEtUFkTbDIjgXtMgt
6hEfG0im9Jf8tVPt3vLRB00mo7LMbGDVEhkDgfkV7FDN29NhblQxWlvQi3kw0ikz
AlovP3Qsy6kZp5kznJh8WLCFYAwJ7Bu9AgAt+smlys7WO9754H3iJWxluv+CC1Jj
PapTAA34dygx4L2dCe3ZBU8Ucb5BmEFaDUWT1QVNIHHmXuBox5bGtU8/4NUjCPYF
zWoNx8Z6gwX3vbe03adNmYw2kGhGh0JGsycEMkaT0+4R8eXDL50/weMbQFQNU63P
QLX8wrlvbdJlpJcxLdfpdUSq2GY2U3XV8JYqnOKgzmcNv3R/McQHwP85IQE8E/O7
vx7GxqJywXfQyNBWgAeUknytBUzLgy9RAIzHCM1dDY5HGP3dEFujJT7CAGKrS7kH
efTsvPjfrFbqwbHXGRD9z3KNkiZomKGuOaunV3AlrQbCsDzyx5f/E/B5UdRrNGtk
zPmBDXlx8SiuhBda1F5FXgPHRX11sHV9n0HyHcr9o1BX5jBVCJNrkPRc+C2tE0r5
xwP4i7NWpSw8v85hvxKfnafQhtffV1m3zMQodNeGpxQEDoua5DPjiROd/3ypkri7
FcOf5uDrO5dphVT4vUTLU61wXOB/0Pj/RwQUXZ/G6dZH+t4Mi/61LJC2kG3AoKzV
C4SEbBtbDXVish52AKdXHxYVWb2Qs2jvotBMaWVh+UWuGlBKyE3oltz4hxNmbS0t
qyu8eGdWlLIoliA99kj+tWaVPhm/vXdgA2KYpArXGv3UVUbEVHlWnk+U5diCkCWr
LRPJydPXteyQ9WmRQMC5jZBlsnY7Rh2wt6/D061ZhlQsYd2SXrzQqnlsa2Q/hBDn
9/Qxfzep6/ugP7GfPnF91hN6qExOIdg+0rSgAH3zHw1SxyH3vn7h7dU8Atb0gcHZ
5LZMDZX0KZAe6/Z3leO8MF5LRnH2bNYbMIIcFRv/pnU1LwdO9vf01sWsXUm+tV36
+131lA9HZGRfWRdmHzSmoAOgm+RlRMkI/9n7ZV4NE7dkyxAO1c8Ygm4G3opVIDVx
/PgXsrEe05ytMx/2CiNBH7/84vluixjLWIGuyWEuijJ9P6bmAfgNR3NWRaunl1D+
sBi7mBsgBiYKBAmaBiohKH3Pb4sAwsdGRsGgQSNVhkVY0khG4juWVzXWSLT9ONGw
XRdzQxXiAGA16q4bQ5cPTfeW2uOYk+6brpQ++z5W57LCBeKgZ8qZWOKakAHuURYC
Y9A0mJPcPf4hwM2lVp+2yDda0uexFaqyeUNw+cvpgYi5UNppk25U1miXeUSaoHaU
SXyW4KrTQR0DAS1rpDuX9SUjANzWgvW1UFHbjLkCOvdjz/J36fKquhd9Xuh8GoAg
jkLjMM6ZyPSKpchhkNVfKPZnLDQ5GLhViF43mPAUVKLmbc1BsjC8iGv41z6m7KUi
/SjzbQKN0BHl3wyElB6DpJUY9jRGKsMJzbjMLAFponTWStmWrqr6cuHMu3NtrZUB
HYdVzzpMW5j1FxZBKHQcRMCyyBjTxphU2W9ZVQyzXzr4YSVSYl2B8fx5Law0qvFa
kYZAfgTYr0T4+pb8/BUpPWczyBpNUkQOnEuPGfbIa8vm4Zh7vgBKHVrz5vD+SsPY
NCPxPhMecMy0UGEbzftghytKFLKj3xNPmOz/NW0VF76F/OdCjW1erKQp83JBXOYF
LyF+6395wzcHuLewZWMb8WvVzvfwkLNRF1PZkyr37tOcGzGjjs8dJlRmSD36Mgc2
+bsEg6iWF/iLITWCQLYVhkuXbMKRs0nYcAj7Ju5QeJKWCwwYJjkNEfb/XsGRN69l
K8vgwnWreSTbFuKfgp+R9fwhIRwmtieQKPYidBavhK7MIt0FNnNwqdNaWyd8ElZp
iUMjZhBibbtOEVNOXojA4rEziBQV3CLou9r6Hx3QAhO3KR54qApWTi2jjHkVEVL9
AqIWMlTQs/UKBXL8sVgZvtHXA6nlHkpj+V0U+nu4zSNL9054O7JSKb03AvEwJn3C
RNhppnCL1ZRBgOtCL8B79lw1YJa0NN/nqgH+PFBEZ9/ApO6eM4Soa9rxlD6SeIgf
IhrNb0XXjXiVe+ZBHS7Turf3mvFj5lU2C//JC3wMGEDM1ILsniEMHiDWjRlInCkQ
RKO9xb6MIiu8PpI3ipsq+EFH/7PNYdkIRXUpZPkQNUzN1A98WEIMSfIssCMR+buZ
Pgro/GC3xxykZFxXhV38KYqd2KiG7E6broEWqwv7Jf/I93ex+CJUx/xLIzruJIK1
E1VICYGTyPbP19ml4Ri77J6c9vNUFDpCFQYOqkG/7G0AIHMu/RJLU6ZUN2QPIZjh
TZ2q1eVHihp7dMYuIDjVlaC6e7pzVxUF4abr1/vpXWCjbzEhncXVqyaJDjV2eT9p
T9QSMwDeoTV8ywl4FFQ602rVSolusDPf6c9Hb2AdklWKo4C79dfWTTnj7KBMn6v2
YFgVz6WsmPi0fGg3mWk4BO8NfM0oXOfeIBW+R8DtZgt6E9X4x5mW87oPVoutELjF
Q97MpfwD8KXKgXvmNyjAV9IUD/tdofNaL2GgJ74aoginpPQuou5Vt7IQogbDeIHu
P1T0pq9Ttm2h8o3i6DVE4eUFtNzRuZjRzuatIM3omaVumAMbQcfm3VqTd6CZ8pMX
v054UT0cIrQGnP28fELQPCw+Jy6xh+o2u1tPlDVRcYs7/ax9R/JNiopK8H1JccCA
siNVw7d8wJKkxSB+n2pqk3IScQQWsYJYVnDToAu5PEgFRFrhZQ9KZa0NRVG/VTdY
7PsI8+O9IZFwhM6n67PoeC2cgXoW4ttCZf9mvgpyRyhq6SlcU23mswenIbvKxxB+
cMi9IYxIwn9DWG4bflrDqEvLtQ1ullQMOyYXgcUugPQ0/lIkxGXJnYexBsr9oL3m
7EA+92gdRbVxKPbIYW5qceqff85ArQi5QfVciOwXf/8nxxSRJPpTIsKDlJ/vz0VD
9Or4nSFyWRTZY0pj667yZPHug9mqn6IHeAHuLPBmns2XEuvp4FNDwkuMfEKOH3vL
S8z/8DyfuzXZKCrnRrkGGUAFCXXplCEMnYmdDpfDirjcveGfyW/0HPsWqD0sKAyq
avNJU21OQNY9VtMCfSKoJQPJ30FG2l6KWj2GlKtSNbgVVqIOBO1TloqWvdeWsz9g
00SXG6fq47guZxLh27mbnyDd6MHxsfWcHSKqIVIu6Ev9pPVj9KOv4gOzAzKXWfxi
gmL1T7hAVBrXJLzkj9S2m4A0wzG+A204Ok65KLZn2GpwtfeQ4mtjLw6yUVuBS2Kl
+Q9A3z3NtYFgIUx6C7rwOjyuNH0RHz3Y3x5YxBbpcsPDvqhH+yM5DjBmbUkiwwC5
v6t5ghcJcwXwZpQ6TuvkDit372RHezWAzFPTvEJpEsHfMTTxbVgsf8+jmAM5FEWT
56+qbEClngjXD1dcsqaEfebMO4dlLT+EwBT6lDsqqQjdmFryFI7r6EbTpGVJfm0H
LfKNAClqX4B0iEW/xt6vP8fvx8VRxwk+vGY6PTauftrEBrzjfWLGmMwdKUe7o8I4
8IhEQpY/KtJ0fdticxz86pOZeFpH2fyjCBHLwd/YobsY9ulKCCBgzJjvk5nFv1jR
EVJ0tNYXcsw6eT7jG4xEplGLlWzgjQIhue7iPfgUkj2OBCwj/ffBdtTYpvSPQgVJ
VVC3XZ2QHBSThoc+NXeBbbA7FI9WN7PIQV2Syjj32XCNzZ3/Xhcrw1hJv6Yb605M
gBch6LtLS4kecotaqoDTHJ9HPoNtsqKOTPJwZwqG4TGxRGRSJLSuwp0XHKEBVqO4
zXZVJV4Li6FoItuMAvHTI1joZ4N8VIksBKrbgk/b3eaiyTYL4o0moo/xxdxJP/md
EFry8w71aqLTcM1OzZohCggMV0m1NLr3u9dW/D0yzbMpPHN/W/Z39zFmaJ9FQO5k
eaYSwHi6vKk+yU54leZ8jdf+w52JGZBVefb1H7TRzJnf5fNz8yQS0iaJUFiu0Pou
i+lVfCm3EsIvX1b7I7ka3mfyz207/YQIyID5w1ppGRqbNPg3+zA/pCXCtnPDKiKo
j2gpeiAU+xmwf1ctscFXoxKXWx1jwRUP1wvhTf/8D2IJUs113RBwREUh8/8d242Y
bGdgJjJwjhcg6BjQ+LINpSvt1JZKnhgF4vRtDFDot5Rd6Hy4RlzqcxCKX2ViF2X6
quz/5roSs5N0qPkoFQoo8mYHXTLe8NV6DBjzaHFpkI6dmFsMZH6BTu/ih62MpeIJ
i1iSyewriz4jE5ZDNUorAz7dI715pry1q6sr29o9z1b6ouubHdK/lMfxQtS0+Rw8
VRCFSpwRLwL0wlu3XhngMqvrUzeavTN7V79zKbFY0+bhH6Kj9la09Af0Rn9/NYrD
XB4PCwkYAWQOLyXzKnEQtzpCOt8hdvgMxscmeeOKZ/dlHZ8OAB0av/sCioodJYU1
Xpq9y430HvX7y2wo/HJbVOKt01BuecAkyVRUvCrGs/JpFFK30oEaLqybST03B8iY
8SZ0FqNQH2+X5hyAczUJLVWljRUZzcGCgVwHowxdKNOzfHCn4Y0ydqAYFTUe8BW9
sOZMxTqIDZOFt9gd2KbmPTaq3VPP5RB6EUoZ7RAmjhXz/6r5MzN/3suMDCEhoP6E
Q08jzyej89TxWlOjx8UNHIE6I0dLuyBNrVM8c+663+v+Kcdj+K8LrWCe0uW/Eri5
vIid9tuN7hNe1FI3hRAIBChYlHULdWHnEE38qDWfmPE+2ZMoc1CXKXXRRcD/5Uco
RiwIaZoP1jTu3AScVXbI1wYWp8KF1e+uhpsF3LNTDiQHb6mf7LNO1euYfzKETn/0
YAv5++uhwdp6o192Elj5PXDub8+bI+AR2kEkSFfAcxSxVVtif9jN7clXs2W9T3tN
83njJtD/3JImuxaHZqczO2CMsPRv62NuVG/VsPOSRi0GrSKo/MXy0e/a/mnsM31A
hjCpeRpleiiCi7kIlaFSvWPhIb3Pgmbhi3KIWKF3iPeaFJEc6B+iBkHKzVZBB9W1
i0x5kpmmitlvoojoSZXwUXpwoxjyDkX48MKA14Np47cjOg2OzuDrtBH/2o60LcON
Lp/gKBT6sFweHRLQiZkXdRl4FTrB4DX6DMQgofJxDPkMm2x8NVsmYFiPsB3Nwvfo
cYei6/Cza+HL8OZ09fK9Jd8sYB2iy9u/HbWp3R7BXvapiUhMGjMiObmqcmKtpTA7
tp2/8D+cL0Mez6rH3NrnF4txIrGPtusIKHjIls4URIbShyiggux4b+ajS25DuLuZ
U6bsZ0RpqriVhnp5W+28/Xe7h2i43l7mz8SzZb2jZAFJVmCOZgxuj0Y/fWbZLuKC
L20aDoRvousJzQQSkBIlEJPb2SUDrAzmkZ+A1HeaavygDDyi5m72X6iT0vk1xwfz
3GLQaADNP8OyGqVMJkjvXwufAsb9Eh3AXe2yYxr2XLO+4+KNiMLEE/oykxz/aOHH
dG0lp28zGeikvbho9ekCZWNeQInP83uqsQQ7vcQZxTLcGVwPoOs/a2q0o+ddbJCY
0siNYUxw7ARQ+UnGDDwX71z43wMLcJqFwuGQrIHoqcyzZ4gwQ6GTLfffks9z1msL
NaQnqt9PM4tPNwPE2l8mOj7BAuehPndZfd1HCh+hRAcMOjOtbM0yafcJxRM1bNe1
CPtOSodjAoENZYOOvf7Wh5lYAfL2ZA0rKFq3NIOF82Jo7d2UTplufZD8EbIS/K88
jx94y//OM5GJ8cbL1Jq2OiiqO66x6UAvTHqPaZRMbgA2wEgSVtfQeMAUw9uN0FKK
U+Iu33MPZOX7pbD6tCdPlhSlBzyqPE6S+NWkKMM5UcqldiSx3uf4wHu9tGJ59Yjq
jOlCDe68i+1SdUhh6PNINGqEK+tk691vWoRYMhkBMYsqb4nmLW2tXE6RdpZvmtTm
YuB4VL3KbYwLfY0Y4uFxf1XXosUe+oud4bNEa460CpRU2kzAqNy0RsP4uAruOtoS
ePa/wUia7/cMqQs/cofN0YcBP3OMAhXk4JzqY0ZijAXTvD3EwHU7jKA6IFJsgbJe
Bzvy0PKW8uM/l+OwNsbNO4WgPhJsVZ55LHbmT3WqkRAQNyEV8OdhjKgDxpem92bj
U6M4b05adSVmBIgkIXUDPCb1pGqpKk92l3NP0pZHngSPm7dYla6UPppYK+swafBc
JRBNOkaOVhJxSlcRJzOP1byg6E7LWdWGJvQ6RoG2HQHKnmEfVV09/hw+n5eAPdgH
iQmXlA93aIVLYmEcrw1qho2vUB3wBrxMN9gUWbCMMni3lc52De6o3aSUcYVSvAaa
CzNDG95sfm+PRzxh75I3bST++NG7WLTsGiYxGkZDIww8ZK7Mtm+d7K/bvEs1zbc+
vggWkxP3L2CWEJyOSt1X0JAlhP3O9C3whn0XnvpNSckl8usg+jVQfcUSDG4BTbfc
9O0h0vVYi0X45um5j3oJXfvcSxoCmae/HJVLY6rt/RIvCgwYYVctbbIg3EWlvDPN
RZQv9BxAQSaTFhmopFKvz4LXugr8ZSguo2SlEBJAiDLWC92fH1/e21Yc1H+d7fHI
EM/cGrRmJeF0SyhgUKlmGyI4LI9kYOz3ZBdVpGgXWtsfNxEiTab7TstuieyNGJv5
rFGZFxxI4IL+DsF25rSRx8fMRgWRVBIp1u8gIDIMHtR3/0AdEnFOqNlFsWJkQ3Rf
s7/+YT4y/mZNusL9cxx4d+ywMoiKkgI/+pkaaFYm6npX87SXvNrV/OlkRAh7qzXW
VVkvYKAF6VZEW1SJfkrZRsJlAs3LBO1W7IQOhyUbHRMKqZcRpaAxTyd0pvDVPLxT
8DeqezJ0lhZkhafEg3xWVfgxQutwERXaCmvL6nx1QRAtwDGPHE3cL+y8UFBGc1ol
iWbKTen13SZH5qO2bhbi4syB1wY48wA1+8FLFVavb+FZw2422y7uPeiLCx8Ujdbp
K6mmjRHFwkTnO7ZGIvp9M2csRoti1CSyXQuOeGXY9/gdiMj1ehlcXBxbD8DlUv/3
8MTzXJqf898pnqAOPS9McYE2YKr+2cQ/8tjT9M2oU+tvgLHoaKSAvHCsf/brweON
wpNMCHVB8TrT887rcNpPvhpaJZNoMBEocHds/iWVwEia2MZuQTn/gHeRCPwgatpg
se+NCT93GB9opz48GcPXNR8uRM2oLA9uJUoOenYYXLPCEczgECqSFOUhESPKm0ZZ
A+gQnSgEp4ttkG8WWteHWf64Ys0OTMQ+MZxyA87ne8onSawBdhdWeSkl+HTLAIAF
81fuHmGel2bnSm4uboXq/NNJDKGmNLDCbXZPpUSZ1NB5Axt7kjH51VcnXx4Kx4lt
qJ0FGx5sY9eLzjg9yYbuhB8hO3BobzPfFgB8Yy3BKreswNgJdM74r8Fi4HtREjVL
DFGG8rzH+2MLYUgjaUF4dVCNlFaso3GqJ+eSS8apZMDnkFXdrZkAa9oVPEwLpzB1
g1MctFeegVXG22khqYdtviJLEoo1Icb6sCC+a4n8/SlIUhiCN0qEsJb0eJlWJBWj
MghC5yfV07mRvN4/u4YrJGpCTTAdmmwi4lrak01w/iD3JocLYZOjt3QH5UPREjx6
DvAtIdeMvWpR1aqs0J3F2Q1iLqLcw7W1XhgpSEnSBXl5/81++ic2Cuct3sZnBc+4
XkzKLylCFr/g2eFy0sahVG70xcfdiMQNbRSF7uid0owdmEKwDwLoe8AYCNgEmqsc
Bj7xKCWLuPaoDeldEJZVze6G1T0TzxMfG6vU8ROA/0t4O0pcxnZwg9DQv21TjEbZ
eaesqIk2isP9nXzC90fnBlwJ+a2NVy1Hbv7USl7VV/RY9T6wsO+k4uRDKnbu35uM
eQLgZhMyMOdxAh5L8efDfyWntAQh/rd4cnqcQJRsW6ERBe0Wj+hbveeSo9na3HZg
bEfbLHAwGQ4IH1yI6xhlgAXinu+IDMhrm0nOXZGZ+BTt7Bujh9VV8+hlhLkUTA7H
OFYXf4oDhIZsmDJZ5uEsPxSFYBdYGDWMC5VGoEOTu20nQPDh0Soi93XPsyACP9u4
KSYm95xy2GEFXVnkWgSx2r2xXCsiFV6koFUDvFQmwUYq+6Hinoo36abC7DlQ3nsg
Uj6MX87IR4UeNZz2UtX/iVpaFopiCI+Wjobmq7mpgkdt438VPso+1bY8xDAT6cZx
vSxHbLhbdELWNlAbf3Hhyj2mA5qCPsJfhctgMMtrELtLQmtkMjgGsI6Q9AOJ/lHA
w+4GPMlcNJS7G7wMBCqWwp8k/ceqj7D8gyFZvIakbw4IQLZ9ikProoCz64kS+hCF
eiPPs8gtJLym5Hk7oQaptpl3SmrkWJKRa5B+SZmRzsfSB55rkzQoY9/IY6/Eaxr2
CKleA2ajlG4e2imX2mmW/j3UAupZUPYDGq5BQeo7O9NHZJvpxp8pZ2qPscV45RMl
QNmEHbBt6uKTR5U5wHo8WtL/oLOl79nZDJRxnjgykEUrzZBrzZyMc9Av+30fqP3J
ZMWdJWOhxZByL6TfpRgsHXzS7OqUXIm9jqqhVlpvbwuNNIXOimQZkYVahKXaQjBk
B+RnD7Orh4hsVkJWiKTRN6JbXQpSN3FISYh+ficyP428hptdt/EywMf0ltL8x+4M
UThog7ieE2ZYgm3NPDhK21IJMCb7nA9MR04Eh0Nuzwq+JjzrL+Pzj9Un8q90qpla
P6xCnvlgSyaGRUuGZ72nyLhUaEsNZARFjCxlkJuKtuYpzik2GGB4IYBB6WhUiZfV
WnLSFLsJKbSdIqj/ImT6cySPFoMSi7CjzUsRWXZ6LOjpBdx1jW4XNRjcdlLuCoLY
gzbKvwZN/EIyuMhRocyMA/5MoFhY2zJKRepLmtyHJYCBqZDVKHV473E7AhIAXB2e
OuMuTY0jCk+actgYCxV0XWE39DVCA1Dqda7Vl4Ibq1FGjFaFvIHP1EjSwflcigva
JeuwAvGPc8arnOjZCoefTR6WS6SsW9yriS5kjAIiCfY8EPB5c4aZiHpAd56qYd8H
1o/D7DjgM4G9hmPPg/p9NUc8C4mtAGmJkVYCcq/pMzTcduGmKM3CSYMXs+cM061b
U335PTWPBEa/XgcSC9NqEv0AZCIw1bIe4z11ziMsT6kw4UpXYblDpzO/ynFUwNcQ
PBle2/8H7r/bmniAFqxAjqcthNHo3LRvlrGw31hdI5feUGcmUuvu9AXNrZgKYD9k
TB2QwjRKC/CJMuOfFuAYRmGbonPQ8serEMh9UKrelJaGeJYOEsrHFBtPKVpQLcic
kCmMqATw7KUQYj7BvzAwuuIrIop8Mxl8y8+zaqGv1QvzcYfE4L4I5QxZiVy2FS5W
eIuMILOlaHJ3ufc8dYD91QzXB0Jahd1M1MsPwiXyqXFc63tz+RttOZ3uFJ53xkdU
Rs6wvSfkjSu45hYGBLNSzE3Up8xHvVQlY5Giu0rxzESznhgehQjg2DLp0XSM9/yu
sA9COHS8xITitg4qIV6w6cmnqXcxGsVp4FcXVDvOWEGJ3HtMn8p32pQ6WT8tdDoW
zwh0ks6eoW9GiWJz2WfOenk0aVX6+W0mtnNWLnJ0j7X85Y/60hA4YDshZyOB1DSn
YOwn+2YAk/kJWMDCR3jL6wKqvo02RrwYEEnpT8XriuYrQ+nB9uL18g91qmfTwgQ0
7MSDQvIk1ULM+2LL/F/rpkW6F/tMOB7+UqvOgZumTvAO/QPCzrZIbdxLbVt6vOjJ
bV5448NMbTmHaJAGVNUOR3ZBdEy4eAGR1T+5BfN/a4pLsGxqWbCXVsz7nOqsgGnr
hThtsb5qoPA9zGbXsv6zWvZiEhVt/soXUHdfLFJKPorEv4F9vhlCV+TaSMAsk3QK
4vG2TEde9xq1TWJtrsgo2LIXhx8KSzKAVHb/e0b8bDDS/oXNqLmerDiK6FTdc0IQ
pHRwKRzwW736OovNOwDvs+h5o5edJCTCSaNGgMn1Mc65LZ3fK5qzh3LRnhlBE8QI
YmxjWxbO3mXdeKPuwMdUUNjsELE07F2ZTsZUZPRjNieK9MHDeZL3kUCZ4mTyrn1e
rRe3dmytmeHY5JXfNNxR1MRdeRynhf9rQ0TxRkdz4qnu03fquNH0ypiAv04deR+l
DgO8Wf5tV4jgLjPASIRW7TDGQpIX9H+hxAarQu/q+j9hgWH2IAU9K3vtFrPh9LAk
IKGhlhl3sZt2H8M0TNY8PqrfpSPK3aevGOFvtVNIAed693Wa+fIeWWKyWYUjy5HA
RP5fxXrKiz45PXAFWicKriq7aKHARH0od2FeDir7FOtj2XFriQ0UR3sNxQhqglBl
YU5O2Yyl1Dobsm+fU/fRN1MnWVSCVLp1PEV9zb2Q0Yx1R4O9r7YzrvexMWnLH82V
0sj45Vut4jilKylJezpQ5YIFcMBCVw+TBM30OwQ3DxqwY4+m6RrbwJ9buAIJ9ZxE
3v4vCQtUQoVd5p5cTMblJrormZIhnpjXZeoxVqXD7wIzxYv+mMBfVtzy0gkGxGFg
TjYM6uZKS8GyFgw16tKmOhdLGuuxRyQOCarmsjNjpiSqxcapUq0MAt/yBjO6POf0
jfGq5HoDfDx1zFXbBvs1IF3q3ycooSr1Nln/zGJ7zv/7Z8K9aWUcvI9MG9/qAGmg
NDq63SvEwAN7iSLzJNUd8eeclTi7vrspgLPj2k0j+gsO1aL1n/9RHX3cwhFgen1h
iYJYlYA/FM7boxfT7zg7H+C4gWYLJm/x547VtAbH2jgoUIq2V6KaeIiCvHA0ihpW
OaYLbnOSF/48+jkXvRbOTg1LenGhtyMHJG1rJwztAWDXFZe8FNrq1CwKSwEsHS+r
4MA/2ghKsJiZbi0AugXzX9/H8Fu5uEMcws7H6Uhj2J1PglpprRVPo7UzCRr2V4Et
9cl73uGLkXCuzOza9bRVnTfGaK/WhnkV5qv9rW2NjSQZYtwXSFNLSheb8YXYcnDO
LzmS/tq2QPDs0BJrfk0Hqwg0Wy4SyHuUh8qvZn8UO6p35QDYSbiNTvwwvCGLvfIY
3wiNd8AYnItZB+OaZn0r9a8AdmUp2x9+WkpQMaZ9qVi9qseA4Bi/jVMg38HFQTT5
ha4gvD2JOJaZNpD02fgcrcbkCU12mWlcLVRz9gASQYG0WQiiaGkamPoAAS/xR5RO
bA8SWmRtHs33044scD0tM7VF5ZaX2UztUuMl+2ttifVabe9rJo/d8++bpLZC0CoS
b2h0pnrK5SFsiHzdVtad5UDx5CftsD5O8HpbbJSZTzzZFnGvPgle10MUy0qWMMfQ
/RQlijSRN3ANIh7OXGLEXvGrTgFkwwNiti+ZirLLSNYDcQjeH2YDDQYBVTWiJ1HA
s9jUn2Ex7hcRpJxzm2YL8qgLp7Mw+h0lDLkj3b9adzaBH2J2TYDSwwwGTp9MMFX+
54K8S8EhsvhgMa8rH1uIgRxR4cOv67EbVRhHjSBLY/YDpgTZnQgEMYG+7itaZ5ZS
hNT1+tYrPc9xm+1PwOwWYvUbkyPO+F+yTsJj16zzw+R96jRpvKw2QRKnvHxKyknO
FlBrQMEpJkDoxtRQgPMwxkiFoLAcz9iJMBMB/IIQpUq015pcjlq5CJDSul0GisUJ
8tB93hmetso4QY8YuhmQO+l+vVFzbvOHaFKIdJqlol2KYxBzUVkM/5jVunf38HdW
hod1sAdbttqn0sDfnqcHdFdTOPdEv5IkZkqyh4uFti/yx5/pZBh4EwR6VY0BrnV7
VUSl8f+vL8enzOGqE5I+80/Ttd4k2SJtMNkqs7qlqV3/EUM3+lRXumOlMY+3KQ0v
K4LDfsRPl51YQbBKboTzrUMGfMoSOB2H4iiZxoVuhb/ahkuWzlx111I5jBfSPd4/
th22ppZJoVy5+d9aQOcifdJO6UrZSIxtGrjMWn5byhX7jPiGUaMJWZvAFEzbQBkB
wpqKuysjV4cwY4mTWprgi2KefjjMgYyOBYe+955XgLxVsFTfxUqgKC1RRMTb4qU7
6M6reDhKaeFukQM9KBHAGR4QR9sHoedJ8CTirWYkCIhx0An4GZ/pxbnag0JEbk/o
XdBEkE0vKf/9Dh+WiuivGzimuQfyUExep9Xm5QPAXVdTujBqdUwrp/0jsbEFjHL0
udXBdQLWFSTD6oTKB/4cJ1pnKK/dk8OT8lkd+i7na0ak9KxbWKchir9nNlPcIXrw
/q0df5i4kWt4le18Oq1TVvXS3UdEWzskc5viC9/1FB/OBKwFjeMLtWC1/S8+qVNT
X2y+wuEE46L8PK62xsklSzQbCBr1xUeaT5KWdM+XV2/WyIIXusO6XkQGtSFLJGSH
SrToa59Rug2f0VH9LpNHyQrfFwnr7NkWV6TVM5EY50RvIzOfZ0CR4VEdYS6FaUFN
o0JhgPpogQ8UIfFQHJPccLYfxXnAQgr/7wQ4KFXhvDGYW7vJUCkWobezD8mUJmhB
6oi+a8arL+1qPTVLTjGQFuy8EXup8tMh59k5FFtizzcm55FHmw25yYRPXyluU63n
WuJqgOhZrtkKBgjBBHfFdUT7EBkNrrvsjHmNDUKkDA5c/cDDIOC4mMteoYq6jRoa
5BBbdD0bbtYgMhpoiGOdns0uxm9gg+83vzs6BAQkVj9aKoLGUWgRFpJ7TDuIUOSp
xIdll3F4d0zY9FxaJIYLAi/8WfyV+DJ5re5gkmgNJR9EGkmyxpgY0vbwVIqrf64X
RO6YdjF2qUKnsSUrVzfqYr4PZTaQiz6ex2CcVH1qXZkV356LqI+SU/2RP5n4IUyH
F1D1RjZJwv4WtrDDJhMjLMiZsndAz5wcY3fVmTG6/6s46OrommOLz7F2uxyn7Fbw
KRRk0IFc2N2qB0gLK4xpuXZ2PJMT4NtuMbRbmyGGJKfZ2aIpGIpw1C6ocs95nYIR
t0kqdHjx+bs03NWGMXbWuQkZuJiI4rZ/JiPazY4Jt7OxpDf7i60iu4eJE0eYEyVa
U8cC9kzqWmvOvG4ZnqS8LDtErc4S+CZbna1iw1fnnf19uNCpZchXHpmzUhgazmua
mo7Hfy/ZubbOkS1WoTvtLcMUZxqrYxwdUezJChKlzczBotd/zIk33XgwaIKrN2Ib
29h2V3Xdy5aGve+N6VQbhtG4jY7McMUE45/JNq1+LTldNN1a/KeThTXiBJXN5qQ1
rR1+CH28uK+lErmyseeB+xX5d7kkiM3ykkvMCkGWiJgorPGOfFUgy+O7lgzkdltd
oncgixU4tSKLwlhUof7VVL0kmtiSZjkjo6RljGQdCGuNt0pywPWTQR76HwrI/BU0
g8r8cGZwyDlPajKvq/8A2Zm6DNC1oj2js491I0LmiUrMjVZmOn7KphqClBzacV+K
47FW+HA8KlG6tY0l2CoWtEMjkuUggZvz0xb0Hn15iNbIikh6XW290yG204Pq4Hj6
mNEIZmj6ncyyEzS677cuLz1+UHVxfV8JFD2FXt/zbUxLbBQ9Q3PKEMMA45cfLypd
/udhmQTEh0mfvMrAA3CEn1ViSXGyX48DozjI0zKR2tSsNIHOv9XzOiOzdHrmyIqW
9vm2Qe+OvS2Tzro24hb6/R7xZQ+G0wPQCW1tV6vXcLILmUpn3I52sAZuWidl7gzr
FnTZFimRK1mUlVcHHLoxuErrmFo+Hu2XBPa5pusC9ii35G4R+056hng2kaRWdjJa
USebrfF4EsYBPg6CjFQ5Ds6lLAFu7EljByjR5eJZMVKjSuWOEXR5jPIWVSl1WTZ6
qJwn/r61N5wFT+JNS3v3V91EbSMXB463dM3lFCawQcpglvHjUKgwTTH6t7l9y2c7
z+wMkSEuRAwuYKOSRc6vZDEIe3L0nkCcP9xUVDQZufBISsa8Cyurq2oD3d+SBJdU
CDCh5IK5VRj4aqOrakEuUCoagA1NmjZipTO24LER/DxVjjnnP5rm3WJEfppbMwv3
3gwFwwNOUtS0UCgF9+C1jx19x/wHcRZTH89/MBBYF8oPs+NiBsTrl7q6wo+DqC2Z
XQe8KM/A9teFeArRnFQVw4JU6fcuXBa/WsujNtUSChAtU6mCDJ6f7poPWMtdQ/3S
4iDL0Sspa45jRUFZoXSvhhnR/rgsKWhjkPwix1CvHYpbSlVn27ACpKFI+kXpGaiy
a3GbLdCo7ZBMmVKTh8jrqdxGVBSCxH5cIfGXvsay1d4OEepO4OcaEXaLS+xS3IqV
AbSf9hqnz634/0/JiS5ZqDnpowPVcbJoirrdFPtoPLosoi0t+KgR2o8or0AMjOwQ
EARL/yD0y81tXAnTBCQfW6om6e4IbeHmY7WT1az34JFkIkKTjcSORFlQtSTU7YYm
WSIpPM7leozYQwp5IJ/3KkI9tQqWaxRWUPG8L3CEREGjldG6I4MMeGzOXd2np+uA
LQrjOHW9ezBu9o/XLa83drLAmwMvKPL9yvGUHI7zUWb3+jAhSv9i0sDVc9cHcKBg
izajSPtv0LfZ89aHtnEVbdDN5gQwJ/WaxKKyDs5rpgM8TsagidYNszI1xjD97nTA
nAvzXozsoLDb/XvoGhofV1siCOZMLe/KxL4Z0F6YtRSws5AYfNQfbfVo0swCBMRH
CKLtVFHA/2Y0nstk0LaXmM3IMX6CuAROyCMvR/spu0YhTLAde/AU7BhGtRU4rJGY
It37FiTMoQb/EzWgE2lTVHzbvHaKt+I/P10iez7eKBQi/A7YJe3RzOe+IGQQqUpy
Hm3mtoS2cZgMdM4QtHLykJ6B/YJnZ2QL72+DxvkPZ3fozakdm6xPuNCUZ5KjBG02
FG3Y4YI3WXeZepFao2SpyB9RsuMSK8C4oQQcuA5ucvIKFbhOeef4Kr/Rwv04JrVK
9qBG3c7GrVHjK6k0vDjcH1o5LAKcky9nBAiP+k8MQI0YX6xnb7fOGduYK67KFMaa
dQxW+owjGX2PaC8ymWqiO2NwexWAU2ntSqhqig7IVZsSmk19QXDWgeYu5cg9XOKX
Aty0JcHpK1z89PhlTqZx67u3JNB2A7G91FFln2Hu1QRFjZ3YyCdzJRH8BIX3l2U5
SRH5AfI5+PXFokS/agWIVsC+7PcXBQrCSgvM4HWricYbjppDjbu7EF5Sclc3fd4H
OGCpcLGbS8UcYdtUaM7qRldYnggiUjFdHALRLiNU2nn3FWABmCthk1boFv2hyqcj
vfjolHdBd2Nn7x6vSF88sGb65wRMMsbgD4aLmdhu3sIsmxpdguUuqp4EzO3mXxQo
E/OW6aD6pmBV94+3bq/ZmY0s7iRWS59GG+Hn4qmyixfZ76DAD9fJfIqWqxth8D0i
ntxZ1TVTgXAy23g8jVHQBsSGVRJqp4i5a+9TWqjb7wH3FvRGtp0LefTjUhzu8w/f
GJS1BLxnzjJ3Z74maPRmknWXClRmS+wUKXyLu0pFSB/gwDjkMyuy+UHt/JzoahwT
D6+XPggW/18FkbgSvK1shqP/Pyzs6tAR3piFkn+qTkNpZxKDW/lLei899rIFqSag
INqA/2rpAo3m4i0YZdiPui/8btEuQRMLgtLXSq6hO+WcSxnRcoFGbqAeQCKqfwRr
c8tNT4F4tzNkpVHKqaMG0fllsCnolbm9Xs4iFwfTFlJ9nVktWXXHHx6Vq43vg1gY
hAfbXSjeldkTukTMChRd+girXOEDr0rk1mHnc5epkgKjMm0WnfMLFJABHoZsZgNK
QspqQRHUPmsegU0DUg+Gr2lhTz1K//+277LAPcZkBStQ6dm2Ab8h2XM+dsfjleKX
X+HG8Kp7obtw/Z4pDUPivVtLn28MjZzWpE9Pwj/MdVFS8suYBCvrJR+FQCzXJv8/
T+VMVLyYm6UCUqlc0ghP3WC6KFGymubmk3z2nUusZ/j7yXZApm5K+NvhmyC3XEfl
PVXmpRd68OYbVwe9D0YreLXI3a2g5hMYoBKX+DY+1WmNrCIrQueyzOCmpMwJ1GSX
pOgg5V3U37ds7tnCnu6thrnB9YzcUlbRfVLyYSB3r8Neox2mcDDXxXgLrHn6mDjT
hHJcFzpykOgMgiEHCSkd09I5LWZbS066OQ9yeGPJqLULHlQiICpYiKSzF8u6kC29
E9GXbam3mJRmE7XXlKFB6kmQSIutDEbAt9uUGSvdpKvMciAWTVgfjLXLPK0Gka+i
yrQnvsg/dNpOP2IvIGdgyIP9MBRKE5zye6g9e7ptHnOflLu+rvHLLH/6REVoVp4i
Rcqewu+H5R7q+v8EPa1xKctv+58aJVKFzNOXdShC5Hhz+CBCo2QUsJ50oXtwRG5D
rlBApCSgK5Z6FzubUTIU6i04luXl99h7bc9Hb4Mf8q6BZMSyyylypyh2/Xvq8mm+
baVzSxwJwCvGiu3uWve3JVsHHU9oN7eU6fDtdS1jp2nSM6R9Mw2ToWR44bhbJHQA
cSeLGsIF2r2mN7Cj0DP4li6KPeBeVDjJ+pXRa/ua1TTxdk1YSzh39kT3NzHs1MFL
FW4225BAQPYq/KMzFcM4KSl8f51fQJNAnmOWogqYpaTcEYnEPe54gQCX5Pg+r91X
tvXcfC2/ZKU1N0Ok4JEoF0LiqBbd+Q0NAVlFPdeMvWvzNrLnPYUeNbn5JaKqZj/g
E60p4a/XzbU82gGFqlnahL6PwaVwEDmCu7kjgvCtTmbd4tcUJV0sUJ54n9YyEEWo
eBJRomowZjludzSz4+Sn7WvLd5QTQ7jRWmP0ye4VbW43xxP0qTAufsbryoRSmezf
SVf0ZIbLsRSQe0KTAYtRYQ+3k2CGec1fyC71Q9sWf3P8PEVgeOMx4V88mBxbq1OS
rvmn0JKwA2OEX8dP8IlDoq92OCVmZLNXVgnbLj8I289UYmz0hVMEOvH0GMB1bP4j
5F/ounmErcXHnecS/zfuDipeQwhwR3y5VN1DzQqyT73iItT/IVCwISbjGMjPtPqf
zj8L7ItAJ2Mj4aRQQ6OJH93nTtAWbbE2q283Lzu4g1NpM7x8OVfOEoaB0FZoBz51
vqpApn7a1MCUxkHOLNK1eRvVOtnqpwqwlG9DNoI5hylLJE5MFOG0hDihJZbsl9Fr
BN0DqYMy4gPJoTtGN51DEhptYD1YBchI3FdNY8ZbwsABlSmoMVjomfXan994WKEb
i3NkT46loNqv1mXCzM9x/6P/rhWvXC7vk4OEK4zAH7f8mzrBRP5sNUDXazqNLzAe
57NbSxdehbU7uRah6RwHNIgPMMsfFV2cN8i+oJuV4Wa2eduvJ6xaya8lCXLND/2u
eHzPelWSO/exuokkqQvVXHvuRHdf2CVMxi00LbiVzdwWXoyAs96JdrHB+X3p2vKd
fjJ4un8KKlwrukB92KYWhqeGBrRbcahiGFshbaTqjtVx463KyIFfq4khGHIZcEEZ
Uue31EEELtyfD3ix5htiSKEJFMBNN34XdjXINIptFR5xHCHVLsV8nrwwimAapkJS
D+5AzBu4GXftGb7+u0kw9i9RmVctsAE2iflVJ/hl2dFBlG1Q0uCQLsuROW+5HOUK
ZByo4srgyQNk0yQ4I6NZd3rxqYz7SJdjFql1pMrSO6UATy9K/FMj/z8RErQB3gLO
b2Eft2uSNMagXD2Y93q4UTnl51RJI+oHKW6StO2vX8uu1gsT6p3x0rWe2tMW9Z89
Fb8v045/wQjQF5OiPNx6Lesg6IHvRIVRy0vh2eyd7HxWlfNOUVHSIPbW92svu9p4
hiMTup2dIaPZTr7PO38M6UMKrE4y4DK4MZuNfKit4L0R3B0uxI8Lt3D/5sHI4eij
878Ub3ozG7s/F7f0hwNIf0/MzTNspUD5IDkoreu8wMZbetvG+yoLahqR89yr7uQ/
ekwNlTTXJN1ydEw2JV2SUIUWVd8cJAo9XNaThC8DT82dq7oTN728xcvNErgJXM4O
PosrMa4+7D0QZeAfydPOzWCJswHKCRtlA7N3rXdPqUr2stAKP0SGwF7beb9xW7bj
E4xR8xA3yC38f4G1TuKn8oLH34IEQ/aOX3DwL1sExcpmriEcj1nzBbBk/SOnNjnQ
834mgE3PpI8kLY++bXDONA==
`protect END_PROTECTED
