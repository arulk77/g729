`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
CJgK6tOpMOY/hOysRG97HyrX+fSpgDJL2xVDZghbprMxn0kBD+1qhwFhjORa2PTr
8nELS6u/PsGTvYXWFSR8kIt0ENcruAKs5rhnYQf0ujinG6lfg4mApjJcIJ5l+jOB
FegaofPB00Q0bZCnzEkOUSDpKvAVlr4D8xUAQ2xm86/EhNQk5yp/7uvR3EM1hSXn
BbrL6YsfwexBIQrmY7G8r68Xeba8yG6a6VR5Eq78BBDASKohnpDcDOJXJiWRv5+8
KdNZKLnYQ3AdKIIF1RYghwVBev5sMrKMTPV4H8NZRnYC8ROSlXsoaGojLxcsIYCy
j+24HEUXtM/FKQWyukF1n5AD9RNqy8BUs+baeJPB82ZAcThpCVrBOSQg66t9C80x
PJtyXAqd04zWnqDUM5RvV0QapredOpVG6sDwLmQVAWp/Gz6PWf24MAn3mf5IqKYz
nrt35SfQayqvz+DT4FUM+rTaYN0H5fdVx4dYxhKnNEqF4WmtrAGHPwkkTFY0rSqP
QeUyjw6pcJtIk5tU67CJgV95KD4QaZmClQTGLg72og3xELVan0+iPnucU2Xn4zAp
d6oHTLsvhjvtjRcEP1qOs13InPnuoMnVbiyf+6GcmTwa/Xd4D2hCCCeipVZtxrTs
afmtjIc8MtdFqYwpSEYdPnJICJ6cVYtMb/6Mbx5EPOkt6WwwVnpi1fej7LqCxhix
zIko5P6ZRYI+7rycC4L7e2ZzDiYMOiohNH6In2YYD3ng+uP6Rm10nd70LyTmkwtJ
wfMcAM/3bSYwEmiN0hx+zLzcUSKiLcluP/aN+auUsinHlZ8OF6bK+RDPsCoL3xh3
WKCy3oAP45vn9c6p//5R92Fm29/CDL7CpYGqnt/0MGvzkLRV8AuhoqHQQ1DxPMey
bAaiqUV0PnxuATJoZjtmqQz9KJQKMFK2f/HoR6WCfqla8Z+E+ETJ7IMn4k9MyZJJ
qoV27iBKDh/Cd7a3B5DSczKwZ+vZdipyk322ecVwRVLP7B8B7h5YbmI/g2vZDRa8
91DIrRE5ifVbmIveZLexHlF5X4BpTn9AEDgFg1wg/4YvfIxEzv7He3k/CCP2WKXB
k4rcf5gDe9Bry5ZAIsltQBC9w+hD/W0Fhb17ACBTbzIn8jm5DW3sBvRChuxSJdJV
ujj939/0PFpXTsWEDOoBMhNEePFQtL5uf+f6Hc25zp1sDIIH5E80r8vR6lCabg07
K5PR/+mnRjhZx5zMQK3iNTZuZb6Mvz3chaQuQYDcske6W5QNjSQeIT3D1Qj4ePmE
Zj/zjLKeFRB2ECCEVq+rzRW+GnvAHv8NBbUg7vRcIQ04bniZB1d/lAzErCNZT1RT
er4/lSxCYKhtcovbBM6+PV3wHkqm7hr/c59VVZPLOMp1O0T3sVSh/oPjRWgnghkQ
Xn9XP6UPV8dTDhUcvgAABjiP2OdpD1oqnvIw2aEk/OMxQiXfPF9UH28Tm9PvLjeh
FlW9UYkNAljG6shc2pjGyFe1pHTmC/7sz7+nWferFzCvBeOmRFjqWI1QhMrTgYaG
BaAcdIw39i8SIs3BbsBc1D2HkFWbALqfmORbGPovy+0lTzsF5kdDMh5j5mMNpO8/
`protect END_PROTECTED
