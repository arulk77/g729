`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNlEW1GfjOnaFs7Pzj4groYP2z3xIPz5IA5LIEKhdj+O
Lk/En6/N3p2C3ZZaDesidQvyLigZxodBwjSmNUFDSdM52Quv2aNPDuY2wD0QIoXL
p7n7Hp9yT8UyO/EThJShIV1WkVMEZFt59sx5XxtlEQeHGRioFkISCh9PgJcvvwMD
vA98UnFXsJW8YZAUs9N8L+pnv5lZeLt9YmRJovMJNJ8pUzFu5CZaM6KkZVVLOhUv
KjoM6N9MbR6bjUYdncKcXm551upHL2M340+oB9rcfWi5vYcD53A5qnUCvyMr8JZ0
lYDS3FD5NF3Z7uZpGi6TIiio8AFJoK7cKCjgneFnaiwV82M5V0f7N/MJOGmFz6bV
RpO2MkqXfTWaOZZDX+QXl1SSd2FhFutCoR7XpV0e3h4hSJY2B2FSI2YIGckDxM7E
YNpDEjERZjvPbA5odq//KMhVLsxftOOYeQ7RxKxWLegoWWL5tjW3VzWIMWBg4EmG
vyXCUvCnZs1/bD85hDAsRe1ulKPI3g028J21crzawgfZ5Wj9Fp+MMWtW7S0IGkvQ
`protect END_PROTECTED
