`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHopNKiuVeN/Akn6Tbq1EBX5ZmcUFcuVv+x7LiTJQI1j
n59Gzx55zEOr5MQEMEQgo+b+/iS8CtCZju8T5aWz3EHyauODhSHHME/ONgd1/c1P
Kwkydz1kwPNtl9b6FhjfzKYr44mjZSaNz8GeSNHlOUFFU+ZeizrHv9omGuwXl8+Y
DUnr9o2LwnHVu3twxfle6cietgEFy2iwrHRmBWzI7sZ/ne1kEIIzOe2rDlgjYe9C
t3IeWR29/pxnAaPVHBs98Z3trddBq8m5L/0kIXIhSF9D2Puq1HVsdn63Q6PrtmDU
K0/zWJdrJJXiFRToVjvO/jDlS9CGAAA4C79TB8HrD43s/VJTL3kK0/5eMloH/mKP
DR6hpDvLd0lz9Ip+fLsbubhA/hNf2tb0ZIiLDN5z+e+9Dt9ZCUdVxP4NXAK+sPAo
hLx/Z7Yt175gXNaY3xf9qF2ej5in4IJK3FG5BZGHZLYtqM32GnbC44BJ7O4acY+w
IU6cA2RqjkDXtZ57LKIVvsd7YGAGFtefq+0ykDjrxls1fMKDJs9VGu5+f+ie5tH2
`protect END_PROTECTED
