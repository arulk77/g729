`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFQzA/MfL1oXyQbMO5CmkmdmaTPJ/HXRLZaz9eE/D70+
Ipr46tWGNA5CJ6wJ+pSGi9HUH/99iEN7D/BtgB1FkSKn/3wmzX0adDIXxLZDUTRv
uRqrgK0fsIdyFh/o263YktxMN/VP5AVmxxefZaFzy+L0So302wi/LirOBXseDwl4
DtIXL+bVeSphMgbLmI4uGfMzr/KCzOKdlDkjGasC0xvUZJ7eeTXjuD+GofxcDF8I
R4lKum/YVCt0We/YCG9nP7/JyYyqD1wGGk7e02vxjVwLlvc6qGlfizLPxcv15nGu
lQVwSz04MJ7uuagFSDQWw0DJnGzekup6f+LdbLm9u/UkXZ0jeMk3pl5PhSMcZTDk
xk6tO205XIOaoRbzNGeSMupakigy1YPoNM3wQC7KtNnW6CQL3+9GfP58yOsDZkWU
depajxsbQS/+5yDOst01f8NjK3uKLht9PexJZhyC6Yu5YZj04K0uzNZGrJPRM6ZB
h8se3u5XaqmB9ES979OOEweORzi0bCnUQtw+zlzom+G17PvPQ0wm0JB/vn8WjO0y
pq/84LRqpc2GV3p7sFn1qXr03WZVz4fZqSQpqlcZdJUg6k8WH/Gs4MZjytce8gdg
CEBB8kFQweKtY4abxLfH8puaGFpx4SPCIHPnqz87wKrbm2853VLbPhmW06Im9c27
wdYLbSGaAvZsfgVDJcHGeQUkb7kk8ZxJjvfuAeCsO3LAJQy1W8f3KV0MfJU42Wk9
dIkGVM3HvcdfmFFTdCgXQoa48ONf1v2zrPvWbp/cdJmLN4MkOgUyQMQw80dXWtYP
nYrgW4Enddq6phUlGCw/59CibkxbvgN1qIMhp2ZnkIY=
`protect END_PROTECTED
