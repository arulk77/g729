`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL4cpJ8heo3j3SgfkImJYjcmh84B96TFTCyz25zmjghC
iEPeDWmZMZdpp8q9KEqDEJDPI+raAu5hWASbW0vQEgdlhcwsi0s0Rlbu193LIZ4Z
6vCg1XwSWfonuyjisQsJoorFx/GjE4KIn8oY+dejKKXUxsKPmBYzik1SJ8L5WJRM
w+5//tdwtGEYwDpAwhKm5wMcfIaeKXhLSoUqgo1zfO11+nPuPq3Z25bfTMOVXx4m
jrmy1E4H12npp0zrxPwCn4688D/714OZ4aFSbrDKA0LogDjLMltvHY7zS3ZMCMTd
uj+dgKbNPWKepCuWF4An6rO84Uc69chdIuTcx/SELU1hSvru2uamkcOlTY2gojYo
WaciUpECGO7I3Ow99LaZmD5T1bRdjDQ0cELoNW2LMUyz5yzn4yAwpI+tqTP2NJaZ
`protect END_PROTECTED
