`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEE1IAwcci0latksqLkPfFtv9x5C89mkqNmU+NdQY3Ue
TDYiEsaK+0Adj4HP5T7jeFj+vPwGf9yo9jawZdJy+KKscPjVGOuIurhMhJUi4axA
wIpMSiTD9UyZT92c0iJeAKmx1E5uEn0zfpHrQg4LSk0MvOcZlkxXLnqNojFT3IQ0
tBdax5vfjhZVTGIr7hnACMzzX7VzKh74kTx8Gw6M+jSwa4UGvindXjY8kTdll8pv
FXT+eQpg7JQxgqUWg4LZGTdj//T71PAsklLyrizCS+i9gigUQoHIbaAHmVgf2Q/s
C/7k4TW3XMq1URL2Fifl7bfKAHOYh0oVC+bbo6+iEcJk1kXG2oO9nPHFFQmk5zE1
e22kM/N2O1swLdI3/J/JWDNH50aupGiXahXDH4tVdGjECB6n7YOmao7KsCMPV32x
YpELhMcJo0PBghXwYk04RsopW7P1bNt11nbnWFDhol6J7zE1jSdsBWvtOjBqzOIK
VNkRKGRwTouVEyNjBb3uVSaIJCt1s1k9C0zrRjG/2kXZeLJtWDG7NfRorS0YmYCK
/DmpYeRTvtwlwEsJNyG44ScofnHCt163B48YqikXf9Q=
`protect END_PROTECTED
