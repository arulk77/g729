`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLVmxNpCezQsoFrmnWSD8OLhfJufjysYQrkqB9urIl6t
3vnG34HShahElBLnwVJYGx3yXExnvILMHgDUiFM4W9p+aqmxjKvA8a+bUQB6WzeZ
aihv4UNfoVqWvR/AqXwf01E5/tiV65oOY/XvVZ154Reain3kfMzvyszjgohhtunV
imVJOJ5/S9pk7iTxauZDGX5+S0kVmA5NwRqMuxKzC00y4VmG0/+EFazRm6tcD+DG
iEE9xIf5H4pjWXIp3+lqC8lqZzJHaB7TFlkblAUQc2VeshCqWfp86ifqLPpnSlhu
YRtdPbBgR/T6cRtrxl+FqPg582so9ire8z6I58IBplrblxYwYF9ax0IBFHpmC2qV
XAU8q26OTWa8216MyOoRl9HHEjwsqqUONkFKMyTS/biba0B0PotCHSaGVEbks1vU
LGaHdVBcym8vc8mOGm9/z9x4rbXnlbbNOIN3hYilsbNVO/lUEI+e7hw68i/xr/HF
Otg7u0zb5mRJBf0fjaboOtJN4AvHkz1ySCSDbaGqHm7uNzL2YUzDKO+rRTkHU84g
`protect END_PROTECTED
