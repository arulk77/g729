`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePNIUancy5Anlv1ISavZi34AV4qshUXZrDEe34iZDd9v
/p1waxPBaYrihyHRiVWK33Su1nAtxtesGmIJAQVAre+ke0ANCCR791+qjwAeifMz
SmwdQHDdAqtooDpZQR3gvBUdRhRXGcVm5r8T1LyD+c93hBLhsmwbt3IBXO7v6w5h
SzQz2M1s7wLHljMCUE1Zh4/QVS0fUD3IguRvnI/YATN8sm/OUUsQJxcuDuXdVHhW
jBy9LvJxIt8zfIl/bt+FWDTysa50q5yKYU92sGzv+05QU3CR+SUdnzWUxjBLtShI
BsdzQmEitbgjez1Pq47bfA==
`protect END_PROTECTED
