`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEPrngxhsks5Eo26tJBnwctHhTiYEH6YRcs/cIAI1cAw
YCD2w4v/6rJkoD5KvX3Zqbzg1EaEQgJWSAXt8ji+SbXbZconlUwQUJCjsjrb+tfB
VWJntepNG2k0BoXi2Sx5id+4RGwmPz1R3B97lb3cJsF+csQE98fR3X1jLxz6Uqch
NIkLW18qzg7xlp1LSeDb3tpcYelkgZogPmh7r91GF1IHb4aFxIhZNePben9uHMkq
gb4uiUVblzhm+cXxNY0Rq3Ls+BpIQAs8huMd3XVN6RjwG1M4NHfd1NXiXjNXkftI
aBL/8ipDC2zFiKFDSr8vPKqVMnAmFFjP9/Cf9oASwWuebIIRVItd1p6fxDFFQ9nw
pScxgOSoLypUZwmiZb+01tN5zOgcr/9H/S9Yzyj+08BozWr+3voqLUmuB++p+D2u
PtVOdQPLRNEXYnNocX1xAhWIzinK98clovCarANCI+3A1F9C5YD1dM+Vu5TCCQ9i
gBowGCdhrocbcJ+FIHA58JwUIGXWDSK06itxK49pu/Mh6L3PiQlog/WE0K03sOY4
q3NvreP0zfXvqTD3Jlxn0KeZR7s7QPiNywEDsShCF8YwKFNgJWboJnbPD1e/Rhwb
BkmK1tY5Q/+MBFGbeok/nX4N5yq+lcZN8X5fPr7fiw1wQZT+yJ05et+OzZM1hA8Z
Ika+61ENGCBYWUYWkFaoVjnHPMwb2SUs+5OUmjzoHXqA3qDviA095wEm7Kt9caPE
9YivIY3IXoLuQRSikDTW7Q3jWo9EDudMacO44RjN2fzn2sslYLlYWAeWbK01zs7O
QnMUDse7AjvQpJIMAzpWPK9hiSdlyNKO3STTUDQLitLrGhIartb9rBq+X4ZulrX5
kjbbNUggHE29N181/ufa+x3akiSpKv48RBqi+3V+7k+mUcQpSaUMNMZXtqsR8Vuh
OPR4nqz8CCGPRD6OTCiNboNBC+DneryoKQ5p0QPlfSuV5JS0N4Vn6JQEGr8Howxm
sxUO/y/LtE3sqrOevnE/Xr7xq6z0BGJIrOmW828xmwc4ExlboukAZJpLXQB2PcWG
aNygZprahE0IdX123pijWVXXVMJDOuCo9lSG6QijqSra8RMvdMiDMQ7R8jmy3reg
Ygx/U15NheuN20cI5zEaR76OluQ1TInYus4fzr40C0dn9qmY0LP04ylTN/Uy183c
nbZAGl6euPyOJT6s1elFIiRpeMKsfniU9QN+wyrGKi31cXurt/wkF/P4gBNXAcbw
+n/Awq20qcXaTSwM9LdjOZT6wBsuwlaBl9a6WBsGuNGwVjMeg0V+NkYvNs/i7VPb
pd1InFIoiOSHXwofbhZbpLVmJWfRKOImeXlRY9vPot0esvOE6OAUzHzSD1YWZWmU
4Q6QapluxV5k8NCf2v+UhYJg7UJGvHpa9LW3kwo+Nq16XckxK+jtUMFNIitsTB2j
aa9Rcnf9cOomq2W9GD/UpdU0upv79g4sruDfW8KW622JDDa2wbydnXx56UyAXcU6
LntbnUWiPH1BLEZcHLO7hUXzZanl+Iq0ArwI0/ioOzPi8sazHihZvwmum67W2qxp
2rM5KeNkiuFVkDa/9kha/Bb8KouMUWeKiModZbHQe46i0tqodDw5s4N4GnwpSPFg
DChBghogY/GGhrHpxqkOCcjOfZPSsed2eZiXq0UsBZrUTKd2C51H9GeJ+JwlXnVq
fFH9ogBzU+R/UzgleDiRJzx4e4kKOLq3H3DQTATO3AoW2stjZ7ZE/2aMnegDG+QE
fSUmZdg8fahBjQaBgHIAty/ZPU3/ZEtGI/Wjg6TLekjME4+z/k5uOYguC0fPt2sW
GOSgRPH3+Fw2T85MNYbV7gL9sIFgfR4GUfcewOUD7nCq2kwS9TcDsUIglVoZS65E
DID3II9G3+qWmaY5Ha8u/xXFMSDBkWw34iSFQmO8FD9R7y0K/br4UrSmF2PXu/X2
YErVqi76g9p0P6LFqyP9sy8Y6sf7qxWZgsrVAst/BCZeNucMV40XZqrzrdE/etko
T5Nhl5z9IjXKT/T5Nrl5d9rPhkcxbt41fO5c+Lipp3adXe4nOPYTVesx9WrEztCr
mDV+ZeeKxbI42AEYO2eaVF6jTqnipHorjfME2DoKvma/13IrLS2lp0j+3qahM7CJ
6Y3pwHC2xyd1ltWmJVa1tbTM4z1tadAX/DSr5XRWrCBJ/9Yza80jiwnYRAQbpNQb
LVFT7Nm+DhzGwlFrDlVAtECCDz/WKW7d/rgOrHf0eRhaogQ4bvfqf1XX7ZBgUbOS
sZdh53tElu+9qspKVPnBO1jd8b9MQ/DVoeUWLK3gcFmBn/43rLlGZmDSmRuN7f9k
6CAAbS+N2zYQeeK4MbWs//aj7suFsWdg5N+CucWZxhtP3afUOHSKbG7OZqgZB1J/
HtWDDlM8HSqIAwPP/KslFkHKlTMOrZxanT2ZvYCQhpgQPp5ZX7c/rCTeHxVx6l/A
1NQco0vJhVy3HJLTH6/FYCUvZ5kKLOAsB+fAnrEI/vZgf8NCIL69qFWbgYFkXGmQ
sQvDw7IcOZqtQFDbWzK4P6fLc9jLOE/IpWOTh0QtiauiVhd2cwBFcSs+/4J+auc/
lyPqnzDcEOSjHV2KkWBBr/+LNf2lElCehLkpimdO/2ooOxwnm8TG9K+rRdIP/HN1
hRBCC1Of8EjIqPlpoNqcPv5D6gFQBpjNOlAB9+VEVsEXSGujw3Nr2puf7qAN9dAV
fsXB8+QRdAoZ5QCKGbWo74rJ/3quI6Zq1t6LFAvmpE0I6enhaF8EsG5uClZSX582
hfnsRtCeIEHvdaleDoebrGZZuIE5vxkZy5KP/VdyfwCWYMqVTUet/eLrArBwAWkH
B61FC6DhyVKyLFD/p/6H5ciS1NYgMOUIiD++G0DsV1cVs7NSHK5E2hbole6jgW81
U9plfSigxznUVkImAW8vZUpq/CNZgFfhB1LCxVZF6Gtk/y2k5OTriVyjGG/1bXt0
GBVVzn0x2yeVHJo+Q8eYgBYWA+s1+NH3lE6FQBCM+m8M9eAsTaW5UeY9HjzsDMuK
BBVKdP3tRAPBkH5dbI4WxBFz+F8e1YUoyErx/rkPot0Q8mls8QH2JQsvaNL84y0L
7fn1o7L4M1+yko1cBCLJqhjWsrvLnTy0dWAr6MtC6tcoUdF9vuRAeQe7S5GlCfVN
RQ/+WoZfPc1QuJf6QhALFZA7u44G2Kv/ARmM1nbwwJnFt70Ia5SIMmBcbPthed/S
rqERMFFjYa4fugmeWCblPuJu+XCNS0qgi27fTmTvSYNrqVf/kvxkyIHR/NFZXFAH
9pzaONcvWmNGn3MfEYRJePobc2YtoILcU4otWQp4kvxuvhka/9ZB3nn7FS2jCb+g
tkYKnRJFXTWRxS8+3z4JR9T0E4Anb+W78YNZiMcrx6H4q5SuPVuBTtAyj+wdASLP
fW2X1iBaiH6TTx+40l5jC0bjnugvggtaHMGslmcr4bDHk7kGUmJD67CyrqhaEK8T
i0CZnT9uHk1D6TcQvfxnwwAkHoLxk+wyrFcSvthWavh9qQVNlSbKjAeW7Gv5eAwN
V2bxUqre5H67HGKSLpSZ8Fqne8ug0lxIik2N06paz0K6szsfcws+W6jiKxtcrceg
sbHf3sSaGJaIHeijRD2wYqG3iA4a7LyH31ZhlxPZr3epSYhCM3ZwCuD1dG3xCTga
FCXH90dQ2WRIUbU7SroXjzdrfYGhHAzED0Vq49W1cvuNk+PZ16b7u+j+tLdxhTaa
Qvywp14VpWxxiUxYC7LBKa8BhPOojCZu5x34rNLUbI03wdKRy5JtdTx/NiSPQz2B
liJtkpGFUanklo2sbanBKdmdJmJIvwttKDFAuaA91fGN6unN/LuykMxV651jPnwo
8xZfN00wUxD5rQ5HprV8v2/EajuyvTAMo1w4WTEqlcAEsdCX7F2KFecGpqMoegB2
C+XDT5jnzcf2QPgryMqePAfOrBjMWmeKGpc5O/VtIQkf7zq3D9KRHVV3SVI0P7vl
ztBUXL1bk35axU90WxnlBNyi1a4Np7aq98QTJTWf+OCy8psEMbGLr541OC84be9f
DZ3R/0pdQ5fwsf+/3FIwuN7RbMWNbJek3ksFC/1zeBx3kOGY1KzozjhFvEqgcqwd
PE8o2JsQlpfDi4o/DjScPHvm++zM4EekeuCmbFxCV6gHgC14AnygQfE3Jm3NCreW
TtUiDTltna9l7gPAfLfmtiv/2oJK9hrnvQbop5DIAKrqlz9vabnuVRvKAoDkOX0u
DOcUwifwHGXk0zDrpRsIjJUQxtLkRaSQjVN2oDFNK2oPF8ZutVEA/xsez4bGg+1m
vnjcVG9RZhqSSYhYkzkWJf3sdh3NodBzVS+B8NFMXK7dGFpSJAiezPqrNy+x8Lb3
bEmpQ67r4DHM8gduZQN/pXqgV468EjwS6Ti87UiQHP6rDn/yDqUO8DRei4woEWq4
ZKfbAvcBMdiMI3kmhx1DQZClk8ywTzooNTkGLQ43Fo2+03udoJuZd/4+wqZ6btnk
jHICSkDcUhYpLl2QeFcOXSdpwrRIVD3/6Z2pa7Gx8vG6HkdtIGH1KRBhW04EZgTT
ktfUb+Cdq9GNhIrsuQYgmLoeYA72lFTHGGIgD8N6kybSkZXc7LpGv0NMqE+EkY9M
nvTKVCimMk9LIgL9sOFeJe93epUamSFmC2p4Urh/FzM6aXGwaLWz7Dhb9gaMjX9y
HiT6n2A/7UyZQ3ovV7pvyd1ott4+JzfVJtfKwvXMoWyXKBji31L14Amm15ZwP1uX
tAVUMqj/BaFyOEagIlfnJ9Sx6AJPk9wmxfd5yArVtOfsV3dY3XUstK3IYi+bylWW
8Ds9yh2FR0IdXXg3GsOZaT7lDzz5P56YufxHdHov3gEzCFU7SgDZn9leAkqJGhmW
Jh/1iodnjS/aEFa4b1v+6zjj9TSCn3ade2J9g0ljWyjwgtDCgLrbistdU0XMx+4O
piZKxy8zKIGQHajFib2Os/iCjXC8IhDIa9c7u7x6ZZaNTiLrgk7meC0SPeqQmciJ
q1bq5fxin9oLljJ8Iq/1mlP6z+46pYEXbn64ujWnJTJoluauJiZk75tClqvh+8G5
DxjrzMcj1SCwbjc742g4q2Jc21xexsWMo/Gt9PJbJHE/cMCaP101nC4vKRlA6L4M
TgsvFDM0OgAWN4TUNAV7vaZd8Z1+8QjLQgusBy3CM4O9ZjohwgIzTZTCieabMPVI
5W1otM8RFhvM7JmcDeYD8Qbxzo5nELxlcxoQqDnlKkxyqyfeIv5FQX20kOEL4TPN
jAtDXaKUtFHllZPUoOW/IeqGlE7YmwBYgync/5v23TvuhjNj98xp099CZYg3wKdo
q9bS5KfAqlM6FCkDlhwQcaTn9qCxKCaPcVlHbLOuPDz5uHc670FJkgIQYve3PqDT
w4D1zKly/Gdm/QAKOuC8gN9txlUrYr8w0iPd+Qj4weuVdIS45ABGUTps9yaIOrdM
N+j2ZSjk/oEdxBAaAI0cquvn1Ad+iByPaeWc8elNWn33GkPrWPmjz+TFz8vfdjRz
fElnskL6v9UeP0DPH/68ovt8WMKmcmeKRQ1JVL5eEzZpja/5JzfuBuS3gBbIz1x5
sWn/CDnOnY5+kS3asej18/1sO+mfzOwNMl7kvp0zw3FuxJxqlH5NaxNu2asorXWQ
UUBlMS+D5UfKvkhWSWj7UMRiGRsmKytGN9eb0VccGcoKIGGpN5/aqsDDHT4QIKkz
8w1pVv400pcktboeKIV2bDNXktLW9iPBF9cyyiDrRfnAUfj1/oSjbI2l5bRfZ8Cs
haqIKnlSeSOALNQYQRTTv6c6hfYBp6WITV+MY0kdBVrSwbKpKywYZbpcnNpai6SD
NP3/O9IJrybkbbOsNvFtD1JsPuaSYSLeorCVnhPPieGGh+SpC8psRyibimTvyc0y
ZiPrhnWeiArhUojJ262pdLun+ZbgZ+VHgrGA561KRUlCKp0Em+MBravH/qm/vfkL
XvxJqktdWRZyGHNeW0SCFSii9m6qmpq9noe9QVt4rJNoIXp6CxRfJHOyxqTD6QEx
jSnpyYse8Kp6tUXHVSar0fMGIyUojfcn/T97hwtBFazHvG1UBIAQe/J4Ge+y6Fmw
LvYjy+LkjgysG+RtocQRdyuoU/gQu3hMrMPYQtKVOg41kUeQyHOD6RvX4JgBl5vx
rk/2yY2N2Dk+Cd3aNLAcQCs5W4Gr75lVl/0sgjeu+ldFOVwmOjD9LAHKVMUF1N2q
4kPON/uAf757au62nHYRV5D0EdMqXgSUTmeGwpelB0MN5Ysk/yKkwjMJcGqbVOn6
mG+nfb9UvUqHCPSFFvfRzXLYJiSIzIibIB7eR9EdnuV5l7f30VpjP3fJnxPIPZtC
BMd6Htngk0+DVAqdffQwZ0WNTzP29PT7FUDufA6gBn5KNc3Eh8Ikfgtw00gPAGv5
taWznVAwG0hNhfWOPAjQJYz32thO6VtkWg8kylb3gqfGFVOzFkjTn29QPkt51jgE
TQfOsocAgjZDiLA3CFfUik21/2D1Zn8FrIwXXAP4VojNWe2jiLkT1bG+KTWrleT2
SmjIwq4TchhFBenPZU8bUaFcxWYEED7ZyS2q8CkNQa8bzIRH09TW+RDx9zFlg5jm
ULHW27t2LqXVNVtexcN1rA7rGqT25ssmMmB5sQipwK8DfZGDvYQzDc+FySOasVEv
RKx8Ycc8e6NhswbUksZoN+WpPM+hqnQ57mnTkDcRRaxItxzcmX3sTg2FM7wG4r9m
zdcsAcp37ZAstBpty2GOZrWlU+0I5uVpSkIeCN1fzVYb8UHo4Nqqps1tSYenyYMi
UfEqk+MSdvnF1EjWo5xB4KsuxPsER4PUYnF6dUDCd0nOkSG7gz5+Dw/LWpSl44AO
vpDTBQGMNc9GGvr5v9uJww==
`protect END_PROTECTED
