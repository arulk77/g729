`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveABRZxTVCcL29//j22TaeIIuYV9pEJ1iF2fCy8g0EI8J
uO75v2dG2K6SVzgvXWrAjjHBrjgk8et6CKpzcQETsKQ7x9H0g9rM2O1iWg5EgTLw
a2/gpIRFWJCDEixqOYyWEwcoJ6EXhDLawyDtwPyKjGrT32e3JWCuhr3e8w4Ov+r8
`protect END_PROTECTED
