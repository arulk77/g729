`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJZswDB6XXdvkvCpKP24DsHKUA5rpkakaG61FonpPBkw
oLTYZAz6DAyq7CkRwGMWG34gGgTA7riN/6A/A07FsXEGT3qrFB78Tn4R5/SIkqSp
rPPLu/gwfxuthcDJvmFaaxLJi45HPJxwWOH3xm8edx0Je4XMvFU/j3a43oINorR2
hh3vxTZji0U6IbWyRUafgKwTvqfJUKvQC6DQvXy3l12TPs5qdXL0doot9LUNeoi9
B+dO6ySfnPK65bgOUwqm+ySHBWGpsELL6AnIlxTDRHsYYNFic3kgZZBUAn1574FO
lVIOe7+4FtXaYmnfy2FZnw==
`protect END_PROTECTED
