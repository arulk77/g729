`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKIrhGvuIq0ZpT9cl0X2zdEK+ci3J7Xfs+RHjYAZULdL
WTW9oB6xBsJGuCZfZpFIqEPArQ0XFmKYcYu+d/VnZH5HMYO9LctTAcXiVpemUiqs
yFQtLo7z4o5gPDobnjwZitsrgvoZgEEdNkirYEliTXFCD2wZmeju8EuL330z28k8
OIdczH16NgzhpjIyhDyqoIQqhIqc9prpi/dWWPRrKqWX3q/WpZb396nO5CDcskEw
V2QqG3u2Fli3MjQwqCSI1w==
`protect END_PROTECTED
