`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
CXDo269tkFVLssJhCUcbkQVCW0Q2GZLPBRYpY40Vb/BJyhD74Y9cBveY7guPocjL
AFZt7Bohm0XEBK46OqMkLQezYrR4OpJjJjnm0rMdhwVmnkmxfqBD1+9DUecXpcJz
+ed5bkfhgFd3pq2gJi+tnrZMrsp56hI7dGgGZtuxcxcdSLwriW+EF9O4u1ua0uDI
`protect END_PROTECTED
