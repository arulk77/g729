`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAB8C/7yaG79PtY5AuGsfx4kTbKB4U62INbqaaFXyxOJ
EWpX2ZOYa+RMAVHpOMvpM7/Lqr1x5h1G4T0zS/ia/tPPWyHSXc0Tj5NtHu9x41Vc
Bi2zyU3a4N4Ylg3E9SVmS80vfAypxQyL6N3yVaye2M2kND9bpOf5tWWuRdCIi3Ik
uJGqSfQKirzaR0r7i0Ob+5zV3zKBFDhUyRgRNoNtTF8KWC7XabFeKvC0Z0oxcpfQ
vQ7uo5lBttxWHTXp8+IWb3oUxdeUhvYKVmLlG3I2P8GchECZu/qTIX0BoxXZbWYG
UKSF6RyPJGoL2/XNJTmOvGgstwacVKLr611Rrn1ad1JrA7ZTkx+YL4036S4/OGz8
klxYgJrLs3TseLeCVFDsYxNoPdIFHEJX8w3HX1/1iFOEejCPzeMUsHXgDUvMpGQr
squerlNHZhPLiYNkmPiQ8g==
`protect END_PROTECTED
