`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN/HtHME5zkJa0BhVXQIItIddtLsVBoNLJnJ3hWXGTMeQ
SdWkXsZDdpLrb/mmZw149pQBHJxtAMXb0HYacyjHp4V/DQtxTehE1MT2wJY3SFxr
Y5jEkiiFdE+BppCvzuv3s4CMxEaCRplT8GBxn+D0h8yQudT4aImGwJkL0iWJeEq7
jM7jnHIWAXFlhlnFX44HtFCO3a7xfFTaPqHi4qW5l2hDmW1Hm/46nveF4I2bfeEX
uQ8RJcpPlygE+0FEiNHB+atd1EUjNOKqGMND2927z3Tb2MIxJ9aPojvXd0vuIFT+
Oqvr+Nj2Jxme6CT+Hm6oiA==
`protect END_PROTECTED
