`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu457ijOd7XvyQiX0Q707GjnD9ZlFcorx59TjggAGS7KvN
d3eXd3oPY3Qd1FKaJNfJKZFL0lwSWcnCXSMSaSL66Qp2EOd4fX+X8EkYNV9tsGDM
mFGmx+6TmIKX6+61CRQOq+KqriSAc5IlMWVpRgG24ZYw1deIG6H7UufD+WPQVYPe
tQmV6DEjVm0I96qSS1giyv7X55bJEcE5BrzxstbaYx8=
`protect END_PROTECTED
