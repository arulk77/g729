`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
if7OW3neLerq5QTb0GME98yuLI9XqqbcGcOXwYVmJJ9KXq8tA97lclKsF6ppkc0r
o3H6aogkkcyB1RiD9hvcWGZ4JdPbsNj0HEgaGMr3SJT6BGI/pFLFPE9WQemlkc5R
bzLhYOS0XtM8mebDxSQeXvE7Tojm2mx6pJu+9ftqRQeopCPTg3rGOyFiSDeLqkIL
QYmIUOBXDzkfYewxdcMiXXznKZY5E2aiG/fsofEUig8cUHBJ9brpjr305dK/uuQL
mMGPKrMjFdtQdg8jlmXVhqPLS3gH83EBperq/oSJs/u/5mXHHgFEBR8qCbQ0ZIXN
43iacmWrSJS8I9pv6XxELSvUmT/Y9kZZUKwuZJpvVNWO5ZXW4Kq3mgeBOckVi2Lc
`protect END_PROTECTED
