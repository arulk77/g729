`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47vjs6N6MM1flsxP7k9NtPJUVDttvQbsdzXKixx4loHu
34afDMYLFaH8RxbFVfnYsOQlCpUrHPwcJS3oGRNVnwW25YqfdZonjLsiN2CMpy/K
yjp7tkcuA03AW9hfwVTN4uJFfYbDTZzvOQ9GnFHInOvTsk89ANHF7wVchZvt3CBo
ffScMF4BHvjoNam0F6+OBzDq7wGbsB5pyFDyEnm9BXP5In7WJbT5gYjqReh0RarU
97u7ARVkClJjnmQ5fptVyuy/EAnCCP53p9ISs2uu3feK3PcL8LJ6P6VWmHNjrdKA
zpZFm3fWS0TE4wCjJWjoRA==
`protect END_PROTECTED
