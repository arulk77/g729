`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3xrhPPuwiiP24qDNjNYfK+KP9JuJEIzMYfVzJQJzgXPHAyQeQi2L1okEwvCvjt/v
iDL/dR0NNPLdkr+putkZ2M18KcQ0HKpjnDqI1eOcDOl8+ZmkjfIL0/mMqXPAXMsf
L0a+Olmg1Aa3NJ53ldbK2yaH2ui3WQ32JaXUPtMG1FactDGMI1/0iwo+8KoY9RMM
WH/5b3lwr3lHIk/Qh28wXTde+bhvXkP494AkiErkY0fQsGRsEwQhMaFTUnH8nr0P
spv2pGDVJ0jX2MzPHYzhJvFX73aXq2ahB5XuT7+vQ0HHQNrQTasrdu7R1qvQqoVX
HaT2Njsdxs03czC9PX/E26QZvJPRxqcR6cO6+06uoMY=
`protect END_PROTECTED
