`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN9NxAwZ7wTzCDl1vGJtc4cl4mpJO5/P9NwqcJhgOkPH8
bMq7yuqrtDWuqGCXp0wGImHeUVtywM5Por9SoE7BtCnSgZJmsJO2fZ1l2q8ZZvH8
A7Q4lVdFAnYurp1lEZkKX8qyZq9wAEW2hies8uOvzrtfq8kHkE4u5Hj34zdKnYT5
GPffavNUzF+GvqPZ7mR6vG9loLV6sprecFNkbGq/pgYbBzP0/JnegM2w7hXqhsLN
fqmok8tiKV3ob7Lz3J0gYpzrjOfMHG1QaBe6huIbhhh7c5sNSo6yxfCRz3/F9O2n
Em3j6j5HcSXVdXQUwXJ8c3Hd1I2204+GNtHY3qS00VZ+BdRFZtGORguO8wVAmmaZ
PITPB7TjZAfOwbX50ROR6gC5WgHa5E25OO9mvHOk6MDi4RvtY2SzZLxyAFwBOFPi
dlYc+46tiTnksk2vx+ZFHPOqwzVXEzcd/PCnivXwN7vKoGSMxGgnqqMaAi5JJku1
`protect END_PROTECTED
