`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
eBQIYjsMiYLvDr+L3cCtVWbpUeHS551/kpORXHbXUwQo0J2pDurCpvVIrW7c6sl9
YM8Q55m5Pw3Ws+5nAbCwEOBrK6DBsBGAnk7zLYQTOGgIbXTCkDDZk0ruBKdXpTgO
KzF8TjP84H5xDdaDdjXFjyQpFmwGFF/rrKdA+nJjUti5TcjrJu27RQAkCUe/usNR
I0MNnlQWCZcz2Z37PhmVLUCZTLPyjBTcloj+R+LIMeRFFeyAcbiZxMxBDxUcRTpK
yUDt7gx02X7142npTF082Tm55IdwqO9z/hVwLeoct8MvTsoqH17P4WNvJAFY8+mD
`protect END_PROTECTED
