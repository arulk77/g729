`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
AGSlDU3wWOO+vONDPw8VkMNDeHqnRcPulJk+gBK3W4ToCMvyzuPaB8OcERWBP/lf
bDoT5ixE6HV8IvfTxuASHiMQyCRNZw5Km/216qPSUewsTF1NixL/yKntOSD5yY7g
W/UYrUnEETEh9+rrJTzPcTtVmPXGRJ+I+mryJBiSY7haM0RsbODPOTxhYOZlD2rj
zvYaI86F73fPQruYZdLNZ3KQTwv2/rpzIuYQu71pJbxnWHuf9VhrWrhAwdQ7I1rJ
byJh3+/oWqhk2JvP6PEhmES5c75cN4dssT/5iLB7D6KQ62/6luW9O261atG/yZ/H
E13d1PlR52xrnIG9iyOmnKut6FVybiw9maTlzQ9FRG0qxPpZR5tTEHKEBlvqpk6K
Pb6xNqiGASStzboUzKfCuEfJWkxrvUkEK5soqYHAM5S5Ds5T64rsFltj/IHWnEUQ
iLHjkwcZ4hvuDNSDzTkgIlt5KPnFyOmf/yU8qu42EBO5Rfx/YKV7LbwbkUGl4z+r
IcqosnMnpxtAtID8t2nJlPUahX1JrnWoZdwVO1KvOWc1h653RbHtMpHOIYPBpvwe
FfrwrPWwScChfXP7u52q/vZ2h5OpuL8Qg8ZzR5iJYyfBbRlsOR0hN8bgdBn06oeU
MDJCowKU02xUafo85mKgxd/GRw861VTVO6iiafBMkndg9i9HTn0soDuOK0Gd6owk
Hah1MEiET32y6lfiqxkE3o6BFRZireGgSWvo7Jwc7191bOocxYxMISCPUq9gV6RC
tcJ3lOHsV5iIRf0AVjQ8gNXDYa5/VyOgSuh13Vwqy0dJ1SL94/tdKyqdMeFpQPVG
ITiNnYhRbxcOUPn5cAelr7kotO+OaGEksn31+BvNyxdqUVTbkYNpLRgsXbcLmg2R
95IXt7G/XrrmnQI/v6DNMH7Wp8mF8LBqkVC1yGQQp5Z63081zSYgn4edcXb19+Zv
cPjEI7WZyBZBVpMKKcxxFG5EqFjCNAxkeW2rUkIVWGkLqvDzp2xARPEtLKRhDWN0
24aXP0mgYC1smM134DyrL3CgYWaB2Xn0jA94fwEzCpWcOl1YNwHDAafAdrRyprcg
rYeuu4FcGjtyWotUr8ga3HPpUeGIDPgvQBot+wHRSs/MwQvvjQGOA+ZwtaGA3fb6
gzN0EAXnE4WT1P3Y3uRqruHjqRZ6yI1+jhKc6L+pnYHaoQulK8AnNm/N6/Ek97Jc
2XReMOl6xSQbashWeTs0CR7S7CRkD6EPRwaJbKj3NFsqVCKXKz+/hM2VXY5EOMkl
rTTHunzo/GN6GPH0aULvooHv/5XA0nrh0fgDkdK1TmjBXxtkzGEmMcpsORduGwV0
eUDtxaIq32gPnnFkhe/FzGbPnK1zqfqp+k+8CiFNttXvLmsz8nyejmmycc4Oh+wE
F/93miu50MnGRLLiaWFgCJMcKsJvApi79xAqQj+UvVy2gOWOp0RB1ml1/zxiInHd
7L8fP1AQr8HVZdddJZMCjXJvCgFi9q51nyzy/v85aCFekqe0B287H691BxdWa+6O
cbcqyYNJWU8QQvwQxZJv7v+HNj6sK23ugoRjQFXQBVJLAF0k9AdEYWDIA6JoGfid
Vw3bJh7z3xXyZ7Hk4YoAwTpkRGaowDfrMjsxti+4la64wVyFfplN7wkT8gJF6ArA
HIg6NGZ56wNgjpyV9r2SK9aixNAGs8DH6SSha8NEFzDbxvACbfkQtHBDfLzLzSeD
q/pFS7xRXXRzqV9rrkEBBCSmtBS1R11pHjhI2u7b9242TwDARc+miGulI1yYANKv
QPBPnJwWd3N+GeIODtuRuRizLbma3VFwxUvGfOZS/T51xpXVdPnCoqBkoJv3DEO6
nthNK3r4nXTY9JbhTNLBgKl2pxPN0QCXKzT3GhqB+lu2m/0rA7+m+YwcqeT2uAUA
YfX93DnMr3Uu9bAlHzJ/aiIFKdlO89u7YgpHIKyr0WqDOzW3uIA40uIepd8umIOV
6MCMsJXPyQwVV3c6BYS95w0aDuXkKzMKkOT7jGu28MK3QqXyg2cWe7CcIj+IcGmz
VIPj75CF8ds1Fh+/rnAaAIOwrKA7wcTQ2+TtUcbHe1g=
`protect END_PROTECTED
