`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveE14kkXI2d3v5EEvPmKEtdDy1/HpyE6ROJDymO687/DR
jNUYDhm5tLUWrchxP76NE+LD0K6laGL+CNfZT72noib0audo+4S5k4rkjOXMGzUL
rJ/+vL1wF+FQgSy/aw43GC4qPm9/iQTDsZGDz6/zErDk/9ubMJBYNwvC+B8Vxbct
j4HXYWYiqYOlsnzOOgRBHb9lfwRU8dseudKLKjouLo6VFQK056yUVL7gFXNb9A7c
XVGzdE7gx6VO68VjDbYKz01z2ytx44x1V/4g/MQDisGWbimRuhKbDW9osgRIvT7i
yMh2JetFygwEtshBaGe83sN5yjmO+oG4upaviTPx9HnPjeCghsOufC0u5kxg8r2a
4eYgTPzNbAMdp3yI63uThps8Up0H/5mLOGQP74oSEJVwasAZURkEkltnO3lMdrgZ
npzs5QpH3fPgSfiQE40KsMS972x6QJUDG4mqtfYWrOXBCYecuJzn4lwhi5+6/1zg
0fjcMBHL6nMxMqZGIQi0N/q5S0NZC7Qagz085Kt9u2ZQZ58nBJvDRuAUyMSYrIkk
qKSKaGxsPADN/0C60o5sJEyFLKQdipndZW1UEnMUfqCpg02f513A309IDqDa4fVW
5aIWRzwpkRHYa0EKS8rw9lUQi8ooJbmXghu3/uGacTXGz+xnaGBVuN3cxy7ux3B4
npFA6GKIrYnQLyI5iAZgncJxHj3RteuDN0slJGoMahVEEUbxoXNXl1MWxZfengHQ
+DM+JGV82IO0zKpayyi1w3hHIjY+Mfy7i8B+ycyaMyrGqeoHAx7g5pVQeFYtl/Ig
IhjNLTuFyvmJ4kgvBbzPHPudPEhRSXYWU6wUp4yzqb8=
`protect END_PROTECTED
