`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKW3e0nM/vyBRCpi0SZqK+PmISV9gtD2bM75hved/mVi
NJI+k+YniO3JooxLQn0sWxYcozyqcHy5LfiDxbr7EW4pPQeOpVEiTqbvUR8Yo3xP
WHa6OsWbQd/yawI/3KSnrV/e2YDtGXw47D9D34VFFKV5TYHt5I1828fQoMg1HCdI
p2e6cPPD6cyelUZSHLg2FjpRGUMcZWtPf+X6horGY/2KZfwO6shlVfG24/XNJl1o
`protect END_PROTECTED
