`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xPkvSHgiTDn98F3S0id/z5layGcYi6oW7kmkrIxSBPT
uP1YRWvw+kUak6oq7jsHLG1EIzAm73aOBUXiaeoHwuvA/BpxaHXmWda+yU4sBIJF
vXz3cU8HQSS6RPp3izzWeRdEqrtoWQAwGRS8Uh1sutCT/B/90GqysYkwLN+HVvWo
ljfDfkaeOQNv9sM15KeGcGBXHxNixELkAbKaHcJeIK7v4hX9L5OAmMKFdeoAOH/L
XSWiBGy5XCihWzx0YzSjV8nCnThaQlYb4z6WfvWLSulSMelA4KSF9BYQ8v6OtQ0N
FHp8s3WjhrU435hGPp2Uxg==
`protect END_PROTECTED
