`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCJAhPqLXVfpmEYFAJu83BE4+X9ypZD5YRItVyeRtgKs
GP1z6ikoDYS/aKC2P2rf+pDqZqMElOrNJYe0tSefI4rAxDRSuMa1UuL9SuRfmsbO
PRWdi/1M2J3O83rVy38GG7+ja/vIQ1GBXl/kmKlbTdLx2/p5TeJoa8JD/YluXrtw
M8OHE8N/J+N4KfodhErxuLKP/1z8dg6Uh4lQ5w475jQHVgrJYIADk9MU6bslLkgo
cgGDE+blzIAWwWsuh903Pz+rYdKdNxEvQVHdYQW3h7VxrCqSwAmzUUE9sjOoIvFs
F1Kw2e/ZIIlDCigIagNvFlYQnKfM7QI6CySVo1iSwl1z0BoFLC2ZRGmL8uk1VOPC
LFVvdx/Zqkn/f2jiXZZMzzd8/SnZwDLI9Zoy7YWcuJ0DaUA98Ni/SgVIjGBtP1TN
CtZkJuxYLl/CahF4dUqKibB4iHxkYp8sXKCVQF5P86gWf5A2ArtAeLYBQk0ugesy
muqHNZJRFzbKEFDfiIpYlHHOAEZw2RCInDrX8YCJWKeMx/A3nXR459iNB2ar0mnT
Jcq9r4+uudX+jMFQMm0TyBkJAMRTxwpYB0Z1rqn0OqXUDVQvrxvyo+9hi3wDtjR9
jPFXJhdnMb/FeZ5ay/71qR4CHgczkObXcUyxBu93Hk0qEk43wT2vRFG+4SmEDOnh
FKFerVuTNStknDx6MyleZjMOeyOgw7Bb58FbDqnQp68zzL5Ee8F/HqZt8y7quk+a
vuFpsmkjtSs+Ys171bmdPZUTZpNLel7FMOIXIOClEwmR0tmY6CLnA7bZD2CVGlIQ
oJVncyIXZqZMtwIE8q9NYeXGdJD6Dtorqp2TmzaOFfiOr8JlYeQ7lolTLpwg7vf8
6kwss2own4LMAB4cMgpsYR7FIQ69yox/qQ2EJ1xEY8Lu/d+JmWdcbDzXA3HjruXc
mAUMpQpaM835GrJehrT0hMpGlsuuf3WHZ9fy8DWW+KP7fUmmy47eSZa3sm7hQCeX
kF9qdXyoF/3a+WphuCWUPkARBA04hJ0tHQMBvHYohAoo7BFIs3C7oKckhuJShItm
GVmReUHtXCE2x/AeXAoad+kK5M/2ra9X38p5oOxFjmlj0vglIJzl3ujHfmHxj9Bz
vJbxvQ11h5H2rFhuTSd6KawdpfRWkJDaQaVpHnKkYeGOXrf8GE7TW13sODx9nXXK
w6rHTK+ce7ydFRTLjh78oMOku9r9Dw8wWd75CNUCY5pHbWjUDJEa/vDnP+7/65A1
eDOKgJa3MMQGhXL//Lvs6IyBQT57XbILAYzxCLseL29ABLshIf4FYKXOYRRAPSxl
x0O0sSsF8X7dSHEH+Pz/I8VdKyG2ULnuB1FaaR1WC2unxLxQH228dWHZ+gbgIKJ7
OxIB4SYzoN+IIUm5jypz4zY69sBKhcTlIC3Ngeo1rTUCDwjRHaVyCEBrgDSEv2bX
FM9lOX/WmqDIB7RRNnS/YF5yNUZXs9dPElZyNfS0ZVTaYOcfzXtVY+JEGod/14fS
GAdlVoF4ydHb1oqu+wiI+QTiXmO81WrlUNXrJsGtkH1Eo/QEbKHK5YZ+z/tNEFZc
Kpf1lvGpHGV2yXvkwHeUjPnXkJTWylQwKpsoLI30msypHfrevpP9XMKwb5Z8MVHL
nqKUqr8dlPf1Ps+u0H7FdBuRZLGbnm11V/bAwqNRUV1DueMHOh+psYbFpFgvD0Vh
2bIQgV89ZI0f+/2QOOKjNSDpqiq/hX6OYfmfMVIcoYISCx5CU7fZapGdzIik+uFy
enf0q9w9+NpRI4yS5BJtgFqxGWvLJx/D2cOmp9xI4YtGcPhvckC5e5Qy/wSgSVg0
B4pcx94USfuWeUdEsrMZRNqY/bGELWnPEhYjJpsiAMghNcKpS+bvaOonKuc2PtoB
6OunhLq+VT4WilYMmjsi/ocws4VE/a6dwrQdY0Dw+N1l27e5OOKz5U2hmtwmubE5
G8ZNc+3aYeajBAqpGUrwi9fb9bOrx+85rC/9nYT0U3/YXE3XBaYgZigUqYuPcn/n
Xd1gDBtFu8dxrkpGYfbBJUTAlAHVwbwm2riGkLTbVVZTBPqLmaLSPhYI8tyg2z5c
xCIseV1a+fXMkfoGgVNsT8fW/0QLI5YK+1QgjkwmcVJcaz0c0Xeab7se+KJfMo9L
3Mb/2jlup5Rb7rMkR0ZogLeqIytExDM+ZICXAMUspEcZWXtPAQo+qFzsB/Hv+fky
O9tT6Y8yHcOzY43lZc7nEHsRQhPTTBaGqIShzHKF1JiyYuFjBPWKHikUJRTNGqIH
hthDbk31E7nlCbn9SFRdCDGkD9k/kkJqJzv6iRixzSFOnQZ7wYnskfx6rjNGJnAZ
5Nxx1asPZqZzNB4mRskKka7IJgoJcXblGVzAb1QLODVkW3v8M+ZNlreOoCqn9wM9
KzvXkxUC3kqTlJVwDSWsd/YwkIuqCogIXso3pUVvR5FFEYD/7lGOq4IKFemp/MvK
ysy2RwUJ/Ld8/buiHmsDKetL8ioiCCKSl787JBHR2MA5rA/M3YyFOVAskdGAjq2+
V6CzKd6cXqCKg6YPqLmswq43j0E9plaUJOy0ecX9g4eENeQXkUbhlwZ2UN0sNSei
47RbfizvgABxSg6iGMmgAxpnQ157D2+YNdIEJZIz0YCsNiXrOlvW+3MTexg7OKDu
naZVA3SFP9j8sgeWgQfjYHiP0+SsESPS1OjoxwnSKWWTkDYz7pLQPijtqUPBb/rT
thhwSUtwDpmH/j/fbzvfAxpLuxqIMLcAbBc+aAuGm4HPMtfqKRvPdzoJOsEAdGF/
4eBXEoUqUCPy+zgOtKKE//6i/zRHsO7xugWUg2EnQYnNJ/IPwGF6Q/FXuMtLCQKX
njax3TUKJdEcq+hdAtmUM+/jpLiHQxO/opgmwFgSVF6NL/Vg2nugLRykHdi+TEzz
CIcOZPp4oI+x7OSDgkWKMX8f0BZM7H4pEYveJQDw0ao6zArwmkOYws6Fs23QwGml
B9y3/c78Mx1HWvyJV8XzFGt1I7/5IO3MUuNkDPgcrjh/movGs9Lbzb7QW4LOWbK/
icWn6QU25OmqC9uKbTo+OPufLa16I5smlso8SGize9vLlDlNm+WyQ4g/eSmdXz0i
v+xl2lL2Q8rA3rEMXcf/oBNxl8G+Sd7aePIGyu4ZtqmTrcYfQcAOqmcyc5KzAZwx
NwvjfkMNX7/u9l7GHI8WUvHv/Po37/1s7X5+KNuzXHzleh8QhCSB8kGg0bYxsLEv
SZBo4NoShMqaaxIVHRGwytWvwqrGpexwbSWeIrFnfMj9yTPvwHX+a6L8T11S/zAk
KKCujGAlkkF7YSUdAkgK7/OoUm7wM0mrh9K1yoTWFWg+R1jbRreMoBHd8uHsuP3A
dMENGOYsGPPspmmeK1JGUOmeoJ7ZyopID5sKuQOxHdEz/vB+WH+M3Uaqv78EP6UB
4xg/J2CfomczyGMpYo8XbHGIj2rw24q6BW0pz/WXhQce7jb+T+MmyI/CW79Y9MjK
iC1Ad/figw2HzCYnpG+bY0XEWh5xy72E6cgw18ClI3erSDmxMDRSyRnZWiXkwY5O
VK16q5kuZN6ys7kq4xOjFMHhK6XyBIkx45Zufw2TtSCWUMXT3gyS1tqkFWs+efC4
iqLrX/co/W5Dzp8AmOLNSy/lQqo+ukKn5NJCuTR7adkLRmeVWSV7YQ9YfXP1Nv+t
jvZmF+zGIrj2v6LzPz6bO7iC9DxMlMWDzOxAvvB7xPTUK+XqYDLo6bIXhQiXA9Qk
1sScSgEbctKZm3GId5qpGrbBSL/3N2FQfVdCbSD/4Do+V1uip31KemlBaOumTVUn
ADEcEKS/GwUIb28EJHQz2vrcL72A59HkhdkYUy/+luVGNjirV7r+hUHGwoizR/du
dTmTO+bDmHJCwhrYXKP075DC9eiHX7ZxIKehda1wn+G3sSa5zRvvsIOoWQH9VgvK
dB5+TbuL9JO5uoMgt/sz1DxPU3IC83fM/8NA8ua8EqG51kfe0dIbEeMdHG7z9bBB
TEsUFuCGiYWvgnVSJMk1ddsO8SF5cYzom54UTxoeqRPkm9LBPy5NfjZ5V9OhXt5n
/xR68Y/3ltfqU7QQyilou4esP8+bG/CwQKt/IBsxMYLHHykBKbOZKEvg49vY2zAF
2VZfX+czo8SBhD7XVumW0HuV57PF5d7xXpOrY/ED/sIKi2WItDR2OtnCLDTphAQg
tJSD4qqmUWQuFE55VCII3Lr3rRQgSnP6gZFMH0EGAtAiYA8ree0Uq0eK3T9XXbFY
UQBWiRY8VrF5xOXHN+4+Bi5HU9Wur1lpGhS2rJaQ1VZ7uxbtqY8EgHyT08OCCeZf
wwjhvJfV6WxeS4q+pAz99n9kobzfiZZnzaEg7vQpntnmNjaBZJl+0LSvr3m595sg
I2K2aMqgEyte9YsSwSm81dZo+efHd38WYG3VllsoU8yVxMnI9vk6FkYsqLN1rcI7
l+/SvAByZNQJe6wbLtnAPnlv/FowkCvP4PYbFcL0qxVJ0DA+YVhBsv4ac18UvAET
rmQhGi+TJkHLqOi4dR+6a1AWdjiYdtMJGvzmAof3rBsiyJHSrKheVuuLGjfyxnFk
MP5L6AtLQLT8AyJiwWKmpVRJLs4hf0yJ9GnU1scptIc0dHUWKQ89D3k3vK27PDpl
MydLNNJSNn95yl5qQXxosJQ6Vetn0xjEq0fxrXtoB5DwRbFHl1CkDO1NDydFOajI
FEoFTtT7vsYQqeHqJ6H08OTbiP8g7SdMPabuZB5YggzhKTshQ5XMKbd8aoMGnKsO
MVKTRL2PCW3S4X6LaCemXQulLp9woVqtlhieGHv9geE69o12QbLF5j0j9yyONQiO
ARdGr4cV/U3MyBlG6xRLaq7L9bqCXC6Czqa/eBExUm+0dcDN3nPVLZcyV57s/pe+
3dDYlnDP2+Z2bl0d/NLQn0/vDld3hfgN21PDqxkgvIjAZitMcHsdz9jXkQww16HD
IU/iyAqgqVoGNwNs6+cpVw6pg2xLPK6PuAaKtL8W5eNqGPNrQ4YynasDS5lNWE1W
1X0cF5jjO60qzjNB1LSolyz5OXdLc651e2qcf3gwpqfIt7kLHJjKmHbL0NG1M+mB
3ooKSQZtE21hWIL/kfELh2EGEEleYM4JGN8plfThJhKD37Y7zLhTORYwrFtqUWZa
nbCfrdiog2xw6maoWU/EQ/fajuTY6bzd6+NTPObIxCuQ+AgIF8TL8EjQW62ELN90
ViPpYIP7FoIia/9E+Oj7MtRPPTCZLkQEIrU6QDw18Y48TvNPtHs8nkHdhBnxtjld
wq3/8ThjDoVC0CJjwuvb+A==
`protect END_PROTECTED
