`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43W2SyqYa/VI92E0ttpV4lXKbs7om3ycPqzsphrVHx6m
L8TM/ejBAn8IG8oOtNefDtneiNM6xagPpNwS5huiH6BgMcw0HxWSoZ2vkIZ7HFWc
qkY+GQRmbH+JEwb4unK/c5P9C01b8ALO70kJEzhhFtdL4MQAkghgZLLfPfBEr3Oa
N/EmFk47tvsGTI9Fa8n2kBvNYi/voZxzjWHqPKGSeU3kGugil/9lm8QK2mIRaFGo
9WhoLivVWh1CLJwwuP9Y9i1nLfM8QcPiKK6MJSAbDVzB7aleZ/Gx2Q2LVUZKshI5
jYYVcYadzchT2CSBuoI8a+wxNLq7GpNBJkjruk1k49beXnbm6lkfz3SWezEWVsD/
2R6x82geXhxfFrb77mFRUfqVrP/gQR+eDKz7bjLJXzo7EyHBGuGTO0tPvycbg5KW
akVTpP6ZeHCX86Sf3foCDQ==
`protect END_PROTECTED
