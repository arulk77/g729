`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI2mH3GPgo2WLUV3hcY6/16E+AfeuAbVW6+ZpSJBpdQN
JFeu1kOI9X8/6xWnRCEJnEHwDcrmUpJYd2eAMgNss7oaJR3e5sdnrVXkIctDHWCE
fbjipcFa/cYPi19NxsAOsgtn5lNSHvI48jeyNmObEY4smSq0zSpu7QkKJf4ceJIL
jMbM5YpPOEqr4V1ir0pr2q3vTIoCh5dqD9LWh1n65V4Lxnm4uqwmHs2OHkH3Klds
`protect END_PROTECTED
