`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCDlzd+ZCQDEmq47h/HCG9fhTKuv9X/iqlxqz+/06tR2
6UbsTfRvx0EaTPvkI8RVGpTK3NQuQWtg8Yf2ZvSHZ2IGzXN4ikVyy62p3t0WCdZH
7L5RTloavCPev1AcisDkV9J/3qXk0n/y9IKhQKxoSp4q4RN2iEp/Yy5Qy5AiwM+R
48KBJ0nt/YzLFGTIBOPPv7/T07LE80+nj1zFAt1fP6HVueWCATUFOTWybEJ4TQ/q
p0AwuniPlvUOgIw3uQmE4HnMCGnQxj4T4XrKz8KbPYz/aHfkW2o8AoBrtqMgu/Xd
4w9PXTKFp7PfIAeKY1RNRA==
`protect END_PROTECTED
