`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45r6iipdcprM9HlFfqaLX8U6zFAB+SqVGkSg2CqSNyEw
yvrTE279GaXZrJhfdCW4Q1hj1MzJM+QfZDHOVekHW/NuVcsQz97ePiF681mIq57+
jAcCPzkkguiXKOaQPSrNaYBy12SpMnFW2yYFZD8nVJFwk2KH1hdZZGLbQTKE+FnA
sc3OVn9YAdURnLq26z9+5/dN0hWemNYDLUGGgCGTPYTe45wwnFPYgSR3kOBjb/US
aR4J8lwXNFHMoUHSyoVHqabR1ysAj9Jg/t/ikPAuakVDd1YEE1/lDUWlEd96XPhK
ZW62FNB1FxKfRn2SDoz8wHf7LuIavkpZQKeiMVvCVkf7RHq8qgQRwy5q2oHRzUQ+
6/xDb5+un1c+KS7ceB9YSKXKTbMFu1hB2Bk8XpMKfUQoTW8xmzIMDVfgQX2+sbQ/
VW/Aap5q+AJIIIoQLKKzbQ==
`protect END_PROTECTED
