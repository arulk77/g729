`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIuH7sRNhO17WH3GVpe2K4hJ5RBqy3N+yuVHA3/M/US/
9ZAQVKh+cSD0P9JT7eDzhsJXGmVnUw6pYKXzSeXm6wl1tkqVBHsp5vpw1wiSeAv9
h/pNX5Ty6ArIRWfrE1D2hKRx1I0XiQRPM6GtHVvctGEq13h88W7c7utrTjFlldGY
z91gd/Elg4CV5mMFYoNF7tfrAq0SmiiL5/jI/aSS6uPS+xv3MUZBdPuPSvy55sS9
dtk3jh7cAp6yh/YUHWQfBkTvZ6MIdmylQ+PWtzwhByShU4nCwQieX2zXBNSVaj5L
Yc3ShWs3vjvE6kFGc1fqU3YxeP/mtCCkVdPDSkqfF0sYbQblK8OEOY49RVU12Pov
`protect END_PROTECTED
