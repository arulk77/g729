`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3ON6twM0bRyFDJLDX3TyepeGka2HQHvneVhN7DcZvAXi6IGhGVGg3MPBVBktKVDO
jNxSnKtZUQfHygLzLmxSQGZP75olshEnYwreum5POBpLlqltDEtiOmPh071DTE29
0+KYEB3guHJWanBoemZ5PQpJXY39Tn4h9aGt5FWYxFXEpQUjXtU77p/3BF3Y6G8s
wBN/9lZPq+HiBZlxsJZ0nQ==
`protect END_PROTECTED
