`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
xRaK4SukZthoeRVHIWvJQkfk2njl6Mj3lGkbjmEcqxFMlSe6VmV337v5XGYlxCIL
pC7da2s0EGjJurrCplL9EDC/XFWi5whXabxtdz2eDT/CTzPzpSAFiIXIcofHDuUD
cqczTTn7dE3QN58XdU0oxkGYtJzYGjmHY8wx49cPpR8bgCvcUy6IhekHa4PRfnV9
FwDmDNjf0qf6Ku6H5B1fOwORjdF6msjmEbGbj3ciVKhnNuBNAbR0y8v12hDcWr1h
p1Qq//yXjQvxa29fh9LHZhqrIVOjjxZ9uicUtoNA+Bg=
`protect END_PROTECTED
