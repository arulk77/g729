`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFpIRyCVyG2HlmZbAVaLrHRIRlU6mriWYgqnOufBQCLE
CuPNCgurJG1AWD8OsTnlSMzzPp1NM5EPdzaMUGeDiXMCsykgrNubqvIAHxRxOdIg
McewbdE4rsYFqii6f1bCrYSNsZ4llw89+FEHgl0FSQvtIlVOhYwUecJ8HHIUM15X
XWmJ0ucPmnErISjkX2PSA7FgJaExutx8ARRp51ahv4fyi3AfiUPQwlh7Rzkewo6s
`protect END_PROTECTED
