`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
lCp16FjWiK6YWTvZkwyzTHzGMZJqloux5TQH5iantSjIqcPnxSVXiXUs20A6Luy2
QG8EoTbZDv0YnYH45CKxT4RJUS49bqOjcQAqoWQHZERppEh1wkBYchEZoERO+AiY
jJCalCaTLOab4HAEJfgXGZjTGmIsr8NDopGV8FDhbXEfblZBeI0fbVw3dIPVBhRT
pN/dujfeU0OftnJSsmgr1GHjckTYBHGY5QYv8K6a7u1K9eeDqhjGnl6URT0yxYlL
`protect END_PROTECTED
