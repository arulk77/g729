`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
01mlPqm7ZEZm6Qw/zjYfs99ZxS54CBzUGVQ5lDpLEyl6cF//rDcFiFmimV0Qkoqg
KzMbLsFcyX5WBtmku4HrMob20I8U+J1Bc8qPpj8k5G/N2Vzi2eX1luIfkqc2gzjR
y6tHUkHU0ZdRUlco3Ahz51sJOxaEUWetMrEOd2zfnHcfOk1utF8GAuFPt3USZ1IP
lMCvuaz0A/w4v7iVeLtaIxe4sMYHoM6awfRW3q7UsQAAU5LaVAd2q07Y1mLkA8jS
`protect END_PROTECTED
