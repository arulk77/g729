`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePoYoTHo9cejtVuGS4mlzdGLLrn0LxpjxStjQd64oNby
1cfoQ21DqTQ55uN0RaOd0jVdVZL0vvnhufAc8BgJZwE1h0Kre+fICfN5a3eRWsf2
4og9mrbqqVFDsekj30zQar+9l7bu1eKrhWTtX48kRzUhG3scwIDyD4dqSHhi0InZ
qf2wPu9JkAolQZrC20raA/jfrGv0t9MrsdIuJEspZN0Fd6wEWjd6hJ6lPKHnKozD
`protect END_PROTECTED
