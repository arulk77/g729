`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
W52by5FksJUdhgHLv4Ym9G0p/jh2aE5+R9kYbHOi00hDcXybKKz/sk3zIuLQdsNW
/uKaYJYGVBy7FTziY8nnNQV2j3erabM52FgLlUZR5sbTIOdqYUDsQHEvgqB36C3k
EpejjAGkGID54TOWD7UxBytvl5ZNmIgGLyx0+kMWs/XbgjHMB03GRaNJ3hsdMXrZ
njdT1a/4z0bUWKCNs0BT0GP5Y5rIiR4H3TvwnDYfwlONI7JNRtgfigAEgHFP0/Lz
iwDir7jK/0kzCqHYE8GfJeEfsj24teTUmteysiYhGwNC46ArxA8Nr6aHKvg/5LbB
`protect END_PROTECTED
