`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
xlspNqjRY1BLhNC6crCjPr/jbRUdksTT1SoHhKgKGau0R0WACO/SCpgpfxSnQG4G
IOi+gekxl1AG89edcuoBLKXhvmPtItifndcH5fFcrVeIOv/C8bBv7FUKYdxwAAh1
BkcaHPbl7qT8ltB+sW2xargjmkbMh5j+1W2QrpeNpw4rCU5nFerqj21J8PlKi7v/
hjkznbPPSRwmJ5KMECSvS0uhurRwaZVmFbux9olR+ESVJPUChEVatTSLNgIL7kxx
qzMdd/yQfR+d4p2dYyz1C2P+2/ZXw2s1G83d1GNhNSk=
`protect END_PROTECTED
