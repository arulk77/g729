`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI+pyw5GSaBXN7OWHC0I1TThntQUAAduEYhLBTAyHcnP
jCKTtvNxH3UMDdPmfvTmLiNKcJOiFLyTs8lGC80iu7/S81qHmiZRqEBM0etXlY96
9NF24uWZk5ltGiD4YPWTxL4+mreNXLLzF7115OhA/Y1U2IBbNMbV7rFDjZO4x2ts
kUuZwy1jd08X429Liq7S6Vd8k9IZGCjENiFzSDtiS3b6mv+ygOUKjLio9oyXbaWK
5MdVp4rnvfo03ePXouHN/tWWguAz+RHJAA8FKK3KK9cPifLWH/lM1r7Etqq1RefF
10UoSXsJLNTFO4pCLxTIIHpHRF9RJrKGTdJ5DO8GwYzLN03ePuEqpbTJsLUyn81k
X+wNZsHY+bpZv9bqjekyAVrj117hgI1czqEzYjBE9mzog15Ym5did++pO3w1MjcN
mrXK+fDk+0aKBDI3JFZa5wqr03nW++ZRB3i6MZTgeYjbHwae0Pj3xxiwc3wsfZEY
Mz9Pgh9ceiROK6JIBDHN0HmMFCLldBiWBbtR3mP3HAdf8uEnKV9YOTd6DUTmb0fp
adtZP5EuLqAxOFmWv223UKoF1jNV7HAZCgeDRbXeOccGQ9Uj7bhNc3fVAg0k2tdz
bzwgvuIwokcvKck6ljtUjm3BRVGcwzrYSP/yMMuH6gSZFMsk9aqNEZJVmA0qTFaj
8hKTNtNIhTqd9dMM9GYBrFGeiNZKZG+qG7IoV2x2ykv0ZtCB0vSRAoKJ9rwmIUzN
1A3utsdv/0EtMdWKRsaxsh1mGJY0XvBaqafo+rjPSeQAbNRWK7MHLLHqQUlR4YlV
`protect END_PROTECTED
