`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDATuOubTEak0Jhc+j+ohExLsU6bECny2nEQ463nII504H
SBnujpd2lBtAFXEwYl7mpfw7XZSpWy3DcHqCFzBRXjG9c/wWtLMpfVf3vAHJYKpG
A56TGs09nAYQHlxEh0lEMXz6eFWbHgmoD2oI9edcZ4EtKOmLhtr010bJkQ3XbMg0
PbUaTsinN2ZotjZKdz+c82N45UovKz98FI3/WrQBugavAn/L7jPIvr182LclfDog
GahYhck69Sgcp8Gk2Pi6snR3IlOclZVG8Kd8JGzi8vhtO/cFd/hQECezrC9VGTsT
iquGrvgbAUZk/FLaQStto+63g02zk8DYnqAg7J6WemjTplVFAU5P+6ZZ8QRzYJOm
v8ZJLnNaD8NDC05JqtYC/b+AI1HM7bX+OrQn73fo73xDr+rYJ/YpirQd6TybUFAp
fd35jY8cnp5U4cQ9uLshJ0SUCcEwEpHJERdl7AuYQns+zED+9N64qfKHmnqyQrJP
fFM6skevcQ5oT2kcsRNXV8KnYjtwsJMNJ9dDEe7iLT32YAzJPFw90PqXO+cxSHsG
l7sRmy3Z+XHSLua6O1gXnJa1/XN3/50/sLzBXbGoVkfReq+CJMKlKcMmUmk2YRs1
sdBcIrl8vGdNg9uqdEZOxFV+LgXGJ/TjrPjuHLJuELcuTxNBA/+pbYLiUOmhVQmU
y7888WmVJ5m5ypkShp2DbjzI9ze6PSKcPuAwAMdrQx0Bka/QH9dSPMU2F57pX9lj
7Bva+MwiIILYEgmpYn0HAzqD4wwjcc0SCHeAzsiHK8NkFmtWS35Z61+82DQ37U8m
W4x1DRJoDMb6pH+QX5aEj5waUD8zYjHmhKTdh//crHKASlnUyyjzoBpVrIkqB5iT
7NM5qM7rAoMdA6fI4SFJPqBY4zBgKC9YjQLC8w1VQbV3ortOVxcTfh1GyzY0pEi4
N66nCuulwoCFc6cKE9mhINkrPaGxPRGcoBjzQI9Yulou6eYsHHiytu304HS+cAWb
LZ0+alU6zAmRg/6gImV4Bm/5+8rdQwZimOuYoHPruD57pS2GTnQ0H6RQYpKelRmh
KXOgDjyGQ2i5veyO36ynU1rIDZjQQW81I4O4ze15TssfM5dZvzkQ/fij6hjSqfS+
Xd97Enbc7J+uTL2AESyGg8gl6N+UUpuk4weCq8ZqpxziYrLkh8TB4fhFhN9HbhXe
ELUT4NQ0HUUxDGbSXGvQzLeDTr0gCJ/dINXT7/BWXN3dStgI4fNY4B6B7UhoBZy8
gI0diyjDvRXqx9Qnibux6++4A+AQlFTH3R74d4NVq11NBuY7wuhdCV7xxwVmEx7L
jhV5kDapkTnYZgcs+7T0HYC/+OPhYwiUqweSsLJrXLYdcUHndcX75xsxvYzWLeZO
mA0XywfZIY1HkSzDJMucOy35eNA/qth1thJJaTqXVjBriFN6v/ErzxEQMINrrmWE
YbgDo1ogK/pdw7fucA9ZOGGunUJf09IXbV/zSsAM1Jc5HQ0vd0j2Kk7HgKLVdlE+
fOMxaNqFAn4OKgG1gKn9X1Azz3eT3hM3Vt/3BbtNIbrXtIWG+ubfdq9+H497y9/S
BaRbuAqLUsWiYYRK2OWVZfSCsjV0eWJTvvw/jY6BrnPDtwtLCCIXAEbDt2a35SnE
bZO5uNDkn4FL4RQ27ARosIp5aWQhsv3lFi7n+OyxOV0JIv/7NrssHwhlDjVIWzGY
U0KVFTDQnrT0lBhNCrY4EHyWaUCI4zCl2/iKXZfhjV/I7GRPmR0bs2kFE7xtNcSZ
pnA8iePVfIXS9gamWNlbGyHFncvrhqsOq9WBXqsMUoSkyMWQR/2RUZQdpnUVUytA
aUoDaXg9rYiMG3RbxiZi0ij4trUBP0L8+S/Ke2XoFHWaJKBoVvMm9fqUHBaNuWI8
H+xowoJDnZdH0TmInAhPTouGqymQaa1F2uiHtyHV3TTDpUq/VRu9lwhaMeMUB5l9
vTQsuMT/y48L5Bvf40hZuQccZCjcU6kuC4tbio4frzwTNGtmB2qtUUsmJCBqUDNu
jlLohlo0bNzk2RaJBcb00Za/7FTeLWr8zD4cafaxjwZRJUUjBvyScYDvofX715h9
b1BB6aBf9Si4RCadUtCEKtvX+t8m+B9aCxn3raVvfV3x7emsqBZPr4jyD8ObpBLF
GoU8jMISN3oMXh1Au2uerNTR0mX0D2W4aRBAI8sc1NtZDvPVDd2W1+R1uXhgRbu6
3th86uFbY/JuQXv6ZP5Z/f5WzBkaEN27XL0E7tGCd7TDQh7afLUjgXuxLfa/peNs
H7VndV18EHasqFNB5yb2zkq7XZUJ2kFCAOdnKb/hkpI0eZ4T03MDuM+LegbAxQer
+dEHb4suJiZVoAj+JNRBV29idyeQPigwnWbOu5AYTjZ/alFL1GILx0bKeClyMqTm
6iZWwN1gZHfDJ7XjACliEEl+2lYkZoApZrtFxdnsRKqFFfbqcJNpnIg/7DJdxH2b
JRvEwBH0jZtIMEWt643aaolrkLIYPbObbRVqaeNZVSKARCq0CQNR98inhfZAPzsU
6ZGsJz35u1RnKO9wT1QKYAjxOExAmqyIiKP/u9Dj1OatlXALM/lo3H20o2GdAyUQ
tH3fR3mJIPRV9NRfDjQCvhdNqIzp3UC1mANphSu/fLKmbqwr1lYyOrumbS+cBF8y
/v8tHW8hglCiKV6czZ6mYxW1EV5pNkwDwmZ5rGtXBZTrtDNFNnTgXgdLCothzizT
4vJuuA5ZCAlDzkzcpBW4gzxpWZY3J5OYVaeJ5dhTVkgGK1nV0CokJatxU86dAT8C
FtHxxkUU7Zkx6sqJvKeHwg+DiS1R5uXMz49xm9Cf12KcX3DqR6t3c4J6np8+2eYt
pzbkgeyFoKE0FqgzBZWS0NciinU5d5tnTBrYHKf5sPuFF4SJ4vLDwILWZecNqQ/A
H3vOewuO8IEim+Oottu/s6gXqwSrQPzM69JvCgnxq3Be1KfGjbOK9LItFfoQQAYe
zkC56LouM/YXh3iiV5VHh5g1h+8CyxVOrGjEVSr09Q/wBHFFVtCjINOqhXTDsoKY
uPK4wdqlAwf9/D0PcD76r0yV7OsQ1aba+lqSbjkVqCJkfkoqj1TVfsvhWNOxY9bq
ZoPNTdgmhDnFQIBkUDCMlJzrG4PG5btRLdstQIQ584IeGtDuXE8+s+3pu8xaVNA7
bj5spMUEQawmmmYJ85aa7Dmql7UXnm3YVfaBBOjgPeXXrh+kkJRNXSTvPTLLLq7A
GJ07Z/R78vHptmDOiaTApDBqdD9t7OJcJnhFfU/DEc0hztcMx0Ei/ltgNAg7XmfQ
NIRtP4vQdCArfPXFKza2i4V0VTn/Bun6e6ZzaSbagKq15H8mq6LdmRSQ7auJ7A1r
R0dj5h6p+sS21LSq9S7JMxfsqN++xNjr9e/t5nB/y6kwEtwcEwBaopksKRuGi8LY
fTNlTPR2tLrGxyvmpekd7uVwO62loUDGtdY0XFImHZspsNUr1/WIU1ixZijTYSBz
qSwHVlV29WdGBbmzfvoYmoT3uaiY5mr4HeWVDOgj++ABuWUclmEk52a+db2ccQcI
+ljUS+vQJy4pPNBCXHwl5o1EHPbsBGFEMCTIJTU097w+z9u6ytovSJB6/YkLFRdS
lfZHPd62iUSJ3eFtqAPV2A/DpXiMCi02uMSXdXQI9mzlTSQ1wObNEHat61Pn6K+O
mo7UciKI9VjM4BRz+74F9AdTdTgmGSXMJ/XvgqPwnZXhVE0or1jHtIP93Njvi1W3
jKm8roK20nfSB1IbE94b2NfyTe7Eq1J46pS1R1KjVFTRPR7BWC2joABR/VeqeE/1
CwylI/YUke+MQ7afJsNnlqs2xHbsYCNjCvdlC6Jx5PdDlIId0E46qZKIBvGd7UzZ
BBb2Np9nDwPDmGkVkQloCgw/T9z/3tDHjPCzlG1uTBEdqL+gk9AE1ehrQKZl2iNm
H3kWpUpp5KaP110+G5+aLP/JtG3yiaShvlGT5451MwM2kZ75fqfTaFOTzZRacUTi
0kTMPasTAbCq6X9zhn3G84kGQFAruOH7hiKVzyU7mVChgh5KEdZ9Mmw+jbtqGz5W
nXnfiINFJW9pDtIKxgsS2qtNVqXu5Z9RS4B1pVEa5uSwyetKqBRrruLIQCRTAx1g
1cgDe3GQtPTZpdJe8EtfG5PYmUyDEfX7aPhnkU61qLH6ibO2QmbWcgEsfSZESq64
DOQinT/1zNeFKxoqA4MyR/U07GOaoXU+yBJXQwUKOHl/SQv3uOtNoLy3AdwkTgLo
WIcP9A1Dv2BxtyBZ54dZWQYwh3nMAd+VFc5SNMJI8RCcLSmh5EqDyGIJdNV3JkXz
l4/a0dtwqc1N5z1ooYNXr9bF0tYtBA0oiMtGxzruF/+7/JyPCstLgrwvaB64lJY+
EpqQK1Zlm1MdnkAf/I0F2Gtk6sEkEHTaqIhjSSlpOSBNGOmRcFfrwfNhL+83/Jq4
zAghyJT98MTVEWBrfhrvepJP3lXlWAgxhgdB8MlPyWmAtvGPSnKLIk3bbhX9K62I
CeUGzps1CwLVodjtmjoqeYZwgDUyaY30zDr/3uu9l2HuzmsxuLaFe7JtN9JUn3A7
+FB1X14aaN9wV+3jxtusobQ/BiHYDTKaUqMbLLX0wUarLxNnDTqvGNzVfuN3nLxv
iJp3LMbsfzTqB+ilHtxTdf8gcc7cmapMAG2hCyeaDEqFOLrGUyb4nFHPaVIYoWpF
eKh8IAZAZN6r5I879asbp/GgIbjE7uvAGJas7EMrWfwt/DR28OkiMfXa/lhCRWUD
7MSln+tjgRYsUPOSKyxCD+sBc0ggObMZ6aGN8WaH9eOksNrI8ByHRDYDjI1JXveG
kziBhkhvERYOj7dVr6wh13Epzc14+Nv8T6PVp6hLL+H+de5QyTMVeYuMs0qH0oLN
12Qd+4GjFldZW2YIYyWNfnhhdrk8QHXDwGDHsISY0eepwIiS41vcFeKesrP6IoEC
xJx3gCndq91IR8jhpa8jAYD9y+4hDnZO21qWi0Isi3NkfBOfueit2d53kYmhuEQc
Tol6Xpdk7GZmXVx6iInTffD07sBxZWC454HDQPWFr2Dp+tmdGVyKKmjxCwhSlBls
UHm2MGpG67bal8Vd3ByUOzEnO1rJ4uabxVcCA/cJb3brToXUXwcXEu8HW44HRksX
iXjAfh1cZk0RWg+V96UvRTQ1hzpk5CF4ridZtnyPPQ8q+2NxUQWuC5Q8h0RH+G+D
ajHlL9CWW1ed7C60XIvvwrGxzHHNhBHnv9d83lnBBwooXMzauQHcnNXVdp0XImhx
uI9aAcFIKA9uX1Jo7syKTgT8byRtBllYDFBZ1NNJ+KN/0/olXJtwpWHp5utkLfJT
DG2IP5jPEQZkUJnyAu0ak5q/tVJ1TFlkfR8CpqC2Kr0m5NTJ1m/LNDjPaHxeiP3x
0WzoMTNG4wFhDiF6pTt4JRI0tWR4iFTqrO2k93rqeKw6kEnIR6jztpAgbG+jw65X
C1O9s+E612OMGoyOYaHeq/uMxrEPS88kXomM2d6kulxpw0Gj1rQeGOTwc3dxv+Dj
Xi0n9in5asq9stjitM6wW69uNz07A8iGQp0kBZip0Vx7KSQGu9Jv/YRTL2gdidlb
AD4jgeMP4WkPM7PFtWQRSVI355p2iBqmX8dnKDZuyx/TfnCUHNxOYe3aB3cpb/xw
UjwNd64XDgfUmYQffR9uO4d+sL68m5lUNaAHlTZ7I2uUCND9TBOBATiUa59QUfY0
S1GFGA5FETdNHsFETatLborCJbyhMQku/En0aEyvFbPUibrrHtI3S6WY5B5mpqmR
3Xz0YZwOi/Y7LGiqRiXJZEF41XgYk6rs2F613qsBB3M6anLpTG9aV+tuJhsE8IVx
hD8OUDgIGzsijWGHNf8Nq9d80jbJy6AXuMgA4yHpZ1mFP9cS05BUzKupseEfYF5l
OjzEChPZm19DsHYH6DRvfCLHRF1Um/pf3unl8fciwCgf5JvHzPsqrAIljekU3EiJ
9mGSntOeqIB/p2E3jMZRpBnjJ8nLRdBkcK65gP/lGrv+EqhhZmwUpKZJNUaR16SF
8EsixlGPLmn32y6vd+0DrnzpZ/gzitLchuf8xOQWxA1XIcGgcy14D8CpNGJHi3ol
dSi59sICM2a09bLnUBaeKn0e88oBIIhBetUUgMo61dEhYJK///q4AJUykbw5B+9O
cBqeESsF0EECPZeUpQvX5nJ9zsVOivQ5MgA1jA3X5iphLWYlWe2FUrCiHm3c9CoB
w0z3bHV7/VG0yz4CPzRp/Mkm/tI6XH3T/Bs0hAoboOKk6Dr7YQmlrHLTWW6pzDpz
1cS4apsUt1JMXn1VEbmLsk3NPU5EAVA8G5cdtenRB2M1GJem9VdevBR63MHrORMP
514UO1WP3evSGohz8U+ku/jmUl9HyHgrRJPPwDHEZrjM7n0KypkyrcFRLBCNyzIQ
eMwFl6n/tSJ3yWpkGESBHPkp5XOrGOKIa06k66tQ9hyG1cjJrY9V5+arzbIHmGNa
niWzQVQB36cnpZfKZA30yHG/GmAG+WsJZCmUCJwezTfLFUY7WJ5pCwqmyt0npKxy
WSaTWPIufNvTWtXQB4kEwO2/Sb3X6RB4M8j2AgxXIYohsr/KbgW98ZDCs62aZ7RV
GyamS4o8Ik4L6dHgKcPgaOapAUiIhltYHMXX2hW3g/ghgiaXjLRsQMPQ8ssux+62
nj22Ikd5G1pvYsFG3/g/OupyNUenO5G0b+XjfMmdLzBgp/bvqzez6K4NNRNCZ2G/
//hye8630+NNrV2f6CF21gqsZfldgSHCm72tP3H4LA6GSfo8INdbMYfiAhVeubY3
WK0P9ZfgNg9dQo/GZ1Ta3J2apCAwOqSXh2yTaGMtGKEhdBNOnRfTtPRMLRLy16ql
KArr1Xy9TKOeIpUmrDKv+tf0MU00M0LPPtOjx2/BFEXC/3cV8oMOiQ03mXVQzDPl
SxQlBifyPxb9OEXvsVuXr879wycGCwM3mwiYXY96tASSy6+4UVVeU6BZPVq0Dv8O
6+l56nPya+J2Iy/lCsxERhvWK2VOyvuQM5kDeLChvHlENT/HKKnjOngiJkjl34se
6K1ZQ8N2Kuru3KFAqpRMn1M6Ob+hwTYM+IWSHfxglVw55hKNpOtXIEUeYUzagB8h
GodEbbHNmwEnXuXup5nShpviSrCj7HWHhsW+8ZKPFvfTl/DKzoHaMjK+6h0mldep
E8JbyKXkxM05f3ITCpxwRNj6UFTjXGjIy4smGBHqntUaIV4miomygyog7lMewTRm
Sv8d4gPLXhrjMl90mplbMUzidG2QWN3QhwQf6kllADUQUVQcqnTHRjAlnRHBPXo7
HOQ09BiDRJ4df8EKVNsIpBy9dzUhf5k5m7MGsuF12vC0K/azXwR/eqdsLC9RZJ8k
lxDdvMntZlnAV2Ojw6xGQt2175f7UuwLUOJKhjT3+40TiwDB77GGByh+K5U7zvgH
oqPBuO5wDncZAn9Nwi7hzV6CMe8zI0pyWDXSkq5sdqR1UYPReYXhAxWX+24WZg1C
50oMjmnu5xyP2ADDipwuC+TuLNlph11kqqnCJD7qPHHKr6GxNwgctg+iKnknNjbr
gU0/Int4jwtUdvV24IE9TvFLRyKeKubMNO2s2KhBYZMPC2dpz9tjL0CV/qsfKAvm
SNXAzo8BBYgMPxUvGiGERJipBcyhcAOD5xMuSYihzAKfykx9QiOe/5jHW+z06m/I
OqpHEaVNUoOyCoHiPqIO6g2IMsbb/JXdZth/tiHoheiGHNrY57elMNT9gGnAvYak
HFufW8NIyxLd+NkHS4H5RP1MXoZWg6cuBXM4UBKPa0muzvgZJtv2ejyEBz497+6Z
qG7WBXeDseRFxV8AVgcOL4kZNk7hQvuE+k/nDiWrTrwYlhsC3l86IZsGlFPalKLw
mr+ZKL0bdJmTGbQ7XR/1WlxlxYXgumKDupasJ+nH3Qb3+9VA78JzN1k1Fr2v6eX7
IkW229UaY86O7J3yOcLkDOg0u0tTkun6LK6mrRSPqU0sfi0JbTXasuQOZCz3Bbx4
0U8FVuGhblMzaBfwoK2a3SpVA+/lIj/SNRKejLl+RuvQwm/DATy+dvxuHkDlbdTF
gFGJA93EUjcJSIY7TNHFKwMZyv4sVEFJuunrCbuH+ZNnhyrnJ3dUGahctid2ftb1
vSJL32Bv+irFxwM69Au50p3ZccjSxPwDqA2LpXUWrbatp7Ld/FPEs9/nc1bTQYv5
gxmmMuUFbevKeZGzLradlQHjCG9xekgwkOth3PLD8qHeX2XPeGNMDkUEt0YzZLll
22f3L+Nqoh1QnuHqRiCRyea0ijTrl08V2xDtOvTq+jERi4c0MJzitpEOQushrKmh
YRDASXMZWPkiY99TQdGpK11usMK+YiFEf4uaeA+QN94VTxwgQ3mimWpwex71IJyv
KiNBIEGSOm3sDqnk+7ITjL/ewQUgeUMra64L5QI3U9xBnyQTc9wOF7qtMJ5BUA0u
4g48dsh6g8DvcXUc4wRNbrFxU3OPKPs7kxLkEXaYyOvNdHuHQto5/3JuLC/wUQtg
afXCeMdlM2HoRfGhNTVXCoxsI/0u3b/rCmIkzehpHWNYItVjoMcJ+JnEib9Og9+L
2mrxRXXwanlndw45HDywQULgZ6qzboVrKXC+k9y7pppoM/SJBgcZzgM462jSN/SY
e+a5rWJt78/xyblPOlzmrrz5jo9dJn+EkFNCgez7p5g3LBtOTEFaIRGkdPA11Bnb
Kj3Bs1X4ZNJvFFLWAcqUSDgyuZ0hAftPdcPbbRaYuiJpv4bvQQmVbo2krsPZ9PYH
ekIUg0c37dRpk3lt2kFd8enCcilSfOayuA4VNbIy6lwVFHYGtgBfXKuqnoB4tjLp
Gpc5vCEy/JgrGinChkXduNaRi3ZasijMi7foXHAkSgHRIjbLDFtzjXaOd9zEqwus
Dtg6D5YntspPi6WYU5BiEa8uuNgE1yKHBOYqp5Vwhz6bvC+jXxgYfabgzd4YBIX+
V7AV8wn9gFUPhfNPXUy3Ty2iiLo39p9WgAO/OI4E4641xlq5LXj13dbUavw/1zYc
Q1RJla+YeU0WRmpDOXalign2dVhp1bl9KWKIIKfq86t8KuS69fbLi3+v7AfK7oKI
WVvIRJKZvopcnrHPsEdxB3bGgmGYYYJyIVWKPPFcj1CmwqC7aQAH9iiNn1zNDmvp
rdWpi6JVR3vPug4HV2ufZ2n9l+iZlSNdGaliwTlDTSyNqSRSvwqdo4IQMtW2MTFA
3zg/8I8ad4LVQdPP4sCPxXo85CS7SkrKqG6Fl5FGr5H6Yne9fZlDJ4Aqhf+pX9xN
1a0IE81kvVFSrHiVxMWNEl3Lt9SNMaJyQScDdLIX07ZNX3ivip711LgwMWD0gUkv
e+xIDnToQGmLZL6Wa3fIUT4JydtKBwUjI475JQXrTatwgwEzjWkNz9yvlV1Zy2/V
y1ifS0I4v1IaHBFRDReuJwmrbHtyaWEoMd4ESbCBA+6Vx4v51zYLsR70C5OA+wyq
FQ5VowjzFVC2Iyq+dBLeveV0DGeBpsSWRJveMBNEnTQTaaiKiiFRbWX1dERKPX+7
LnalpLNuqV4/UlEfYjK7gMzKBbuONQxJ4j6b+Y85hDU/C0wOecrUFv3OfmM5lXKn
5dhbYdmOftsxekbkLhf+7MkoD+2K/9IvEGUP/Kkzy99TR8/pEz/SGiRck1C6qQfG
fZoRX0rN7erywnOjg/wc20D2tbIZr0oRHJt1PP8Dl6hSMVCC2VZX1Uo2fBrI3h2L
mePhewrFOyvN1mDFglm14/YRXPrT8k0mqBnVw8dxkt0Th+Uzj4Wxu1cfhUib4ozS
b4arYHTRAAAPtUWkbmSW3NqBdpuAXUYj8aRWSLjXf/Axa3ddC4LoTWihhKdlRLrX
ZpFuRADCreBv/+6JHnCVbQMgGk5sIDKAX40voNquNpH+duty4+vt3SW1TZMezOWL
eyok9IfuzoGhmaLQRVI0BcVhDd/+Sf9+uNiHx9Wto3uhHTRVxifqcB11rkoOTfxH
lKPhX1ESClb+zUs5rUESd0Iz1ZE1xe5pV9lNU2oEXSGVpZf5TA2z1+ND6HRuunMv
okm7nf59uY+7btNm8KidFE6FxQVEHlk+47P+ecQHVIH6QGeIXxLrz+aGuD0ueixM
amFC26d1GYeYqkttuRuVYha+ECBlPnxSDPOgjtb5QAF9ZUTdCw4WNSQatWg3Ju7v
0RzRNSDcPL393ISlNuS3LC6AsWZHZ4fuQWU5yf5OTZc1JA+ZG/oLxcfYcA1vy5AV
eEXzy2E1yFc5PKZCjKf9Ef8RYT4c0Tio+ToU8Y7vh5D7l59NrAq0iohg15OBsbBn
PxXnhDvhPRt6/ocANqDJ2mo8XRVXlgy/K0SZMW/Q1lDHZ9SiVPMwTxO1b36xhwnL
ZzkQkC7rZjP0PlXS6zXi9by/aQsvVtm4hMOR8URW5fDcIkiLM8dxCfXaa6JY1g5P
gjwAzrbbkf+MHziKlQW/h7PGRLciB5+fw179OEYzTK24gRBX/kOiJXQScr7VIHpq
I2QKNKVf4Ofq9mK/KtUwrOClAqR5IM2RwmThiTXoIqGHk0RUT5nf1tiwBE+NeDIq
sIIhXNoif5kbeAszSY1nqTyCpXxoZdJIHybtIeWnh2EdEVipNBBxlpGUUGjmxgiS
mUthiO0qVG+SgzCX72WOwkplF5TwmHs7n8hI5WTyL5mJoZr5Gyrz+1GhNxEdov26
fisE3xT4Qd9fXENU2zMlBd+2/5MER+gLKuATwV1vuLW8XoSsccGC3zK30c93z8ec
718rrNWXpbWGnTbTXfwWX3kPJOgkhB6minGOuBsbuUR7cnteLQcWSC3Yeo/GNo69
KXSmi025t14nwfKKxgMH8XKKfo8Hjsy01mS0qWsCKT2AM6B+ODYew/hWsi0fHlBb
cTRu2W6GHVo7So3ZkcHjHE7bQnKsSa2QA0NBFalbTUXxexfydPgtm4eMlVoGFcJi
9XonbDtXwO3p05jSh8qFfQrKuh0MFSTvfIee4i+JPidKuOogjZ+USFNxDLc3Nmyq
J6xI65IVzkeoGpXmejC94KXELwxEKIYMNpWDWZfAFBBQJYslLaWaIoUJaQn8nP4W
41S6YQDYeemPwCvefh/hvngODFLg2oI9JCrMB55BaPNcLJlocImpa9w3a+HrRTp1
Uib8pMIZ1zMe7RkSOzkDpFqeA9D31ZX+eh1HQcyQieygZkYHEG8YVCAiF9ZTftl8
nQdzM+iY7UzMhdJMH7PlD7BZhRjip5atUI3ZCN1GNYqQNRd9ooJ5+wQYRLuBvtNx
LJPz2EZf/jhtxIkE/Lr0xtgpf6sK5TAu4pHcs8fs9RB0CV/vwVArTRNuvNbbeL4A
Quk5QBgFbFz6r/mTRmGhaXTwSArqkgwv0B/2VaPMx+CV8Qdot+9QGrUkKg+pfqDn
h6N0TurBzWqPHnosd/MiqpJsXNTEcexcNlDiFoZGi4PBtEkLWzVc30nm0m9DTK1j
db07BmjrosIY9x6wRI88YjEi+5mMZ8Gg1UKyDewmawgFigSFTs9bxbwWC+rOJ7wD
+G/vqK8b0H93Q7oTwxcOa5hUy0SngDvjpJy7zw8JcquHRnpfPWy4cMfl3GdqSPNf
BJbrsqQX//eiTR+lJlCntJ0G0nztPN60wm7LBnEAN2xIRP8FYm4KpvLFfu1hfFaI
td7fJJs9AWslbxAAi9X0UfvJhABy02Jz3DRTZBojlDG1ieF3HM4ZRSvbeZ0m+pya
7g+AQ4ZwS0v4wgRA7blJ0FN1VKL/a2vfZICDbGCSJE8W+GFAgO47a0rknqyHZPF6
f5xohzd/s4RBx99K81EfvRbiaWoamIwfWkxxiVZlSHl+XI4+D/PUs8pfyjyNqdo1
oKeDgt8hiiOERs3/WseBlu1goA1SHMaXFZTDxO45u5Mk6+fWGs8b8SGpC82RbRNs
4d/JpA3md2L9pBjHNL6e745AFvBlBCWBndXEJ0p3dlR0JoPYUL8KaVFEEulqld5Z
gVuhoO80E3IX5GstnSKp9uQq9mbpDqH5Zh+oJgxjx7zA7ChJOFkbHhVHj0aXhD8C
cTq6yZzZULbMll2H1dKoDJhS5za0t0VXeLWX9sOviTZBmXx6I9svEJWRqRIPSqxc
dJg41TyaZ50j+25KRCs3afTLZhIM3wkCNfFRk2uNN7ntRi98eC+Yn79d31wmnFEJ
57VgPwYe0ge2VOc0aLyUDe3YJPKY57qigLWhUMIeO0lsRoaTBmv66+dvuOd3FbhG
QJsa2LzepLZjyk1gUfbda98czk6gSodVjmbd9AYVx+/ZKP4OZ8h68Df5laVX3WR7
Vld7r+X8aRJAZ0xWP6jG6bwI8HedJI2LmB/8ErtkHcRbjca7ewHlblWsGxq+lLpp
s+VWXLvaMCtXY2IY5lMO57WeFlc0u+CZ4lf6nQ5FX/9MymHBKoWmx2ki7V/DxmZ1
1wN7owYyULUAIf3IQH7wR7gJPZLwiJrHIZi+rz6NKiQrA1NmmiJRLBs3CRjGyn/3
2qof+tNXjsHbWfkDAOP1s+ggf0xbNgrpWOHuCoewWvMCPAjMkBdlUfVBxtfLePx3
5LOOdSOA9hgAlSq0Wp2zP1g1dToZAce5CYDosGLrq1jxZSw47hbZqjCKkYAm8K3Y
nV03XEbvyjcFwiGHoaVemSdQbVnkigDlKMwFg3dl7wA7xEzpG52Q/XhHOBLApPgS
s6G3L1qbHtSrQzfNFG2BObc+56rAbz9c2bYy5Bv/0M5j5EZVx7ySqdP0vWNbF1es
63J2Y1gxVCK6/LRcUyn/y5+vedMZSprvSsAB8fcYuahphO/zTv3ONuC1gUBnD9C2
Km+ZICXJpaTJTYgBIYjNBZL6LuoswN/pGtCp5GWlySdp4gUS9lGAjoTZ6KIm64SO
Xa2wYMQyQBaAeAeuw2ltNHkBlRC+PFAtfyEltIqoNzhIMAuBzppCDuKLwgge6MFN
qhJCN+Ny3hjvcNVS4cVJIdJNVeWaOnHAJeA1P3aFT7yCCWgunxzy17WfAOwhSGor
+wjRTDJh1ivV+4a4Sl1H6YmODjYC7Ggwt1M4mWA2tafJuOqU2fC1DDU9I7X1bxEu
a4ZYIS1r+eqO6sw/sWTZ6zjfZbMW4YW9iCVESH27e8JSv780Brj30bwsvysqveSc
BONCqbXmyeBYRi9w4d7tTtiqsJq7TM4XUPnSie1qBnl7UM4uLgQBhxuqn/e4am2I
bPQ+S1xj0CE/YGUqx464YxV0ItZPVcl2udboYSfv4QOvQNJmbkFW6LbMH0gf+DOK
D2Qs51Opad4nlDq6ukIfK7Sd9R3gDQyfPa0QG8Db3kTEfKee0u5DpSXZn/S1BNL6
np5m/depbqT9jCDzPKp98RzbFBzcHwam7AzmMaBv4HMN9kQxNbMZji4XBKscj8ho
nVNvCz+yLcE0zynnfmNLm7lI08vQ8dwfIPLSjzMKIbIf8MOlWcrrvpF5HwVxNwfc
ffUBSonvweDQicBM4VJGczSJBlryLlZwwhBl/ajVbTtQAG6TIzobiJZvdybgD/Ga
lF9FueZvxBDXECCNdWNLWaXirWxWRkq49Dr6+imK5TIVGXkK34bQaGcfNWl/3HHB
rOm5gqiZ3+bSnRzWm6aryPj17/nLBiWDVJ2XpEkeFdqVa/2vWJQeL+b2DlggAQFu
WXIroSsIdy5vy9kTy7tbSpUJCz8QPu0nH1dp7iahShKPBOgVQsZG9eQFrmEP/wgx
DcjM/23hRfF9b4OrJyNj+EWgYI1K5QReUIK9hyGxvKerH+ysdRAM8AM2CNxVKWyl
V6L7/2eY1RwxYvyYhvgNNuxsAzoPZ/RTRQHBWgOn3ty0UXR3j0G6GvQj7Y7fc8jk
wiAfZ35eFH8enOJSAeal5FIK+3oXQjkT6o2y1ICzN1gZwm2epvOwuM7dZpDgDtvt
TKDnCYW9fFVdHUogWDyFoJBgQNgf08kHOM2GhuEWP+VnPyA7AE2tN+pMIUHb55Q3
XjPpAijmaBiSTXwQ/ATaqIB7zJzyQmx0gBPWBdwIRZ0RJY5r8YLGJjyVhEQvoSwm
mdHqXUUNk5T9H2mKtgptW1+uY9HFOxlXZ+zH4DyZYudX/9Npd/0lYlJsKYoBiUOd
ZGsx61uRpUVRfOhJrzn3ifgRkx93AeK0Xp5zcKoFdKxs/eMsDNQdRX2VIoX8nHSU
9lpTvygCVst7uu0OXIvyM7snQrsUE6ZLAD2uY5YIU9uIgX+imEFLzmZNBAz3IXxG
+T05PGrNoxWEmCWC3+22KM78NECHLh8VygrYCSRl0mU/ekv/GnG2w5ejIumPIKyD
P7iP2SJXSG8YIJR4TXwpoK5otv75DNWbB1befGlGhUjD4WeTQypugeVU36pogiHI
+T6OAqefg2ZJvUvzQ6l/kr4M8AKq4Vczq9tjqRKOBzHhkmtHjOz94kTM7P5hegZY
rRryzXUBICuE3cS3M/vXfwI7KpxxjPYuiiY2pGDrwh6t8+6yN3SKhsh6DaPiPGvL
kIwGxbapA6UeSSoaj8mzlE6A2Nt2sqOG5RyiLSMBPBovHuWpAPqi8Ees1LJ+naWn
E91xrd5lT7OrfSO/CyybtwzpOLsW1EJFhVW1oud3fQ0KnNCLT55aghm21O6Ic+91
PROejyT/OJ8R5tYHyzbyC/H8aVTfKgckXgmMqhyO+YlJqGfsqQ8Jl16VqJwGYjgp
CFg5ofVJvopv1yToiuwzbPMlVeww62ttsCDaHaDKmZkXg5b1exZy6yOS0vK7CouW
ikuELvjwAAhHWUNtPQkfqMQUkUZ3IfSo+e4pX8aPo5HW6f/Jd+UYDJPFtBfsFZk2
Qr5Hl8ugY9sXYCFyRgOJTfmneDUX4Pv6ZYj2nevl8A7SRnAP9PPbin2K4G3iMI/X
3UzD2awuSVUtAsDvZC1iwHFHjFwIUr8erqa17Xc8q9l/iHfW/v15xm0/m7YTI6t7
dTJU9YaILo7SfDJ9KPS8gJZiiQPcJxC7WP9hOwuEu1oF2E+8TDwYTN8V8Z7pggyd
cEAdAPutKCLikBsA8EenvwMsgVXMadk9W9yBtPPeTQsqsfz0gFLN1+P30kSGLe6G
jaTUVMGweAsPIBWwZ//NWD2o6/tDuZmQ2kPW+M1jQp96PWC2ep9dUOd6Q+4SM9I3
+2jVzxwArRCAdMBWmzAgtgq82B5/shekbG9cwGcxm6O1yQusjX+gB7ceSxBZB7/w
Rh4aVw6UIzvI12jLQaxKPrtMI4x2QQOXPUoQFdHHfITdPtBmQxuwj/KMSsyjLvwI
0DP/YK2R8qI2FsXNZRCtDfrT2Q5pNFH0S1FQJm5gfitq/cQ+rtGL+sElS68Vuxia
S4fQWS7iaz8Ky7c8ZCyhfk1PSNsXHsJAHno2igI8B0achaKcQsaCrRKWgyopmFcw
5JaZz/eCTvVzv01LHKReiCNsDGli9CloGFHuxeTk2iICXJa4aO3uf59eLFEhRLSY
uxiZOs7uAwxIxp3gq6+UNj2V/sPNp6a9i13BQHErhUm1NOoVZeVNEL1O4I3SL3Sr
Cwfa/TZInwmIr1C7f5yMTi6mcKF/6rP8FRj7Qqf2GckuSo1bLIDoKvoWkcAK3oTZ
GSIvb6Ul2nVk2tbVGos98TiD2OZV4VNyj+CLfgfqFRmtnqJ9QTSKIwkwAZsuKJiK
t5vr3NSh3raD7jfXczamkpgxRF67KUL7QCJde3zBmm5lP89Cmw5zEKplJBcdbjBT
XUxIVUukcgufyn0Q737HZ6PKZzu1jebNgL8oMuq9jsAyyOf4BvGqJMRcUO/WCOvQ
7M4oBM7oqcmtLpfFLS/OXr6+hJbB+wKVasadSLNP8icboacnkkRG/uAD5kTrHK1m
RPA5acuplIKMRG10FTX2fmXa+wNr5DAcNfkpaT1xsBTkAWB0NyMceU6nqLs+5PoS
PtKy3weQuXguiQHJ3mJFulyfBmdgxeNxyulBwexbHCEPnIYaSA4bU1jggiGTU+14
Vy1LoeDlGHrGMk28z7CGanD4GVxCR4bo26gG5GGU1ilhus0r22JbzecHPVj3Mk2C
LaOJ5VYXTr3ihUSZXOvrcED0Xidcu2vehn2/wKGukYM3dwc12h0ct3ew265h/4Di
Ml8CemjQKN45elXix89H2LfsNb2a/mxkSWXrUOsH+r/GBy5sRmRJOoXOwO7Ns6Rk
y7Hb9cQ0uoU51AJfNfbi9UykjS2I8yoIolYlL0wl0q9hRF0a9gFTE1Uh9EREvVMA
gcm72LNF/YnUWTspFPNOLa9mTVJzwbQd3n0w8r/uEhvS94KFdCwchb+snOw1YLIx
vEC69latrJkTPUUTyj1neKIX39R6rdPPAGJtE1bM0fmGgZ/B/mh4oc5QaY1lin49
gsNt8tEB/rJ6/LECdh670DyPO5ZCIGJhzBKmuzpIt4kmUcSalgfcEwces9ZQm+Av
JM+xcQYHSy3zcqe6ZwRqJnfCuNWfZzTM4bVUvo0MLm58O506NKeW7H3EzZxtskXa
PRQB0KeOKNxTpTj/18hSUHATav30b0N1MXpeifGcm7i1JuI83Q5iLYkgvhF/dOoJ
KhxpgwSay30ESh4F20hHnz/XeM10x5/FrzKK+gf0vHjlOOqEhR7Obl+KX6rrwqi0
BkzYTpLmyorN+QEtob2scWzi+U3FEWV2n0LUkocwLYrwfeLzKm6NKT/z8yd40jqW
HYMdg1F2wFLYmwGgjwE8RkLxD+fPK6gn79aagPBkSMD/67XgSfmFjB73y5ol3wnW
k+V2mXHXkwy1XwBdROqiMug+wuJvpQI3U+17oP2h1U8L0VUQQNN1JG1eP32yDyM6
CmOyJy9hO/DDWQZJsQxr7i8g1+Sc776jV5pFho/ugO4zAL7Ts/BbyQKHFZiQD9nU
n+Z4SPi8S1L5X3T3Ik853mq2e77GtlGua5X8SB1G6s6zCrc2sZiuFbCIfpCR3SNp
++mKdPKTZw7bAyUosghFUROCpR1RgCePvX5IDyEsTsCXmXSxV/+JUKE3yoUlIYsh
8zRWlPHDbv+/uYOZhyYXDwahCLrrdEoWeH3c7AQW/clZfgFu4IFdnWz/zhV61Jqs
GUK1rK6+DjqQlemTW7SYaD5f/MS6lZgf27L8qTgA5e0FAt1yz5VRPxjIlZ2WKKGa
0wueWEeEfqb8uV73x9CFl4CQCo0l/422JalGBg71l54DELXmtiSB/H4Rs30nd3Pg
QTXLHxawoZUe4PN8JlqvhsCEnE4RTsruRY23VhAlRLUAWZJq0LStipPGIup/Hbwa
pGWUSzu0yoZlNWt4hHUWZmypqHX/4vpzc6vHdZeKBJ+Rq4aiBfsGf5MMO89llmLQ
nJI5+porqAERcB575ZDqxWHRZtNAx0WLPYXNZX68HiDUCedMb+/dOo8Cp80/7eMs
oGAfg1pr9TIDSH/exAbUOHaUbYd33Ugtlgi+E4hsK1AOhJDixHrh9j7ECl68nYmf
fOv8iiarW0z07DZXX6qKl0qc2d1UapSZHYCJw0hNQ5iC4sQww5luy3V4oDoAB2+W
XZU9NXf5oCTDHBLXdmOVsC0HQJQd2otFbDrhotg7ppNuogXsHJdKDH6eeObiMosk
9Cdf7CFDE+kEq3x4ybNKyRduhcDlV5wD1j6cACTqyy1V5SY8bO+NaIo2JFRdj7wP
G5CxwBp+IBtGor/QUBitPk3QpmdJtQhnO+2SgQrZ0aHnwI2wZyn5fLTAafi2zz5e
aPIJSX8hkmHpH6DZvXsVqbhYoAuCJDht0cihjRF5P847pl921eukHxlQVnNnra+c
hJIps4XrOnJBTli7rlWtgvWSyHMrdaffMz+Vw/srgI6V2/kuZxPNiAbjF/Vtoyke
hsVnLz1P5uP/FrnbHv3XXNxb+36X+dcmys+NXn+g54x3Ch1Oywzpg1+iSL99vn/W
lZNc8rVzMjzkgaeCgKVR3RmJJ+WeYOo5V0PJTEjZPMY0qqTWAjtIOYkuDD4g/GJf
F/XDU8OAmlecbAZp8ummzsRsE1gR4zLMcE/1P1VDPhxPHw1nEKiKVN8lJz6A2ek8
syswXmfWVxvQsKnXTiEQuBv+LS1xDbFWSiM5sSupmXNRrhd8D1Y6KFXKaCNE8/Qq
aUzIZR0nJjFaMpgEiRDNtysSqIbbfzjvpEtDt8xbLlPGKBWqGOZa54xddvaaRo/G
9uwo+675bye6Zj3BsxXcVkRsaB1BDgFBkOJ4xCwn8KNtptKj40hPDR+/fyn0zubq
SEHFOpRdUnNH9kOF3WRXj+U9+iqfl5M9pQ/Y2SFgDqAgUK250fbYG24RKzBZjS53
VWQia0KAYc28ax2MmB93k3iFHICBAduLTirwI/xP/l5t3CsHk56rFEulqVbO2rH1
00ieQmTkbO9HVQp+r14TDos4YsvTBQkYKxA+XmCDiSwtMVe+xI/3zO8db2G+PpIV
QXBL/pTAeFFT7v1AkKmBvgRLJxAFAkwVEoH1gwgMzH/ABR+1erGlQWwHAynBOvQr
8jhMjOzzbltJoflOq7VqPkUKRt6H0yMgu/bkVlNQreeOjnsafLXXPX+rxpuhmKY5
7bIM15xeq0ZabwRyXpOWjgs6TK/AQfSqrOQzw0kD5L6URrcrPPk6ZRDGi8cFCHXP
8RB2gCxV4P29fVzDj32nrYdvlSmddk+9AiYtm/l/5XNCHeO+7MKs9HLgpPbwHIHZ
RulXusksO6uU3gpVrcIZXq75Re9YxZHBpSaLiNReJoVJs4gAW/b3qiOaE2uDJ6Z9
KJ8POG0JdZsav5vjYZKGJ6uLANKYvRNBoRocZHusyiejIdHC/eE/J0NCbyFkMWED
P4DVYE5DHRgLNKe16SJ2U/cY7e6xntbUkxDklhz9FrqH0jiTRvZvP5sHWbSLH+AY
WgrzY5N1zeey4Qate/9hpcWlKJMA+VTzlamgJQY97h8GibKHh40OZA7Ac8f/fqYL
KlQX+3dnQRpIaZ+/8gIuy0Isb0r0EeGEXj1wSVj7SJP56d8WPsix0HVYWFYn/tXu
rOLY0x69xkDUBhZ+jrkqQ1TMHSC0d8ONkJSEXPd2wJQXwuNlnePMfD7qc8/2lfIt
+xJjAqU9n3TPcaVkSk1P7gsZSj6WWIngcT/kAIJDTwgpfwtAC9as3MR7cGSncCGe
Bzp+gkt4C+U6C4Id1E9vkLyTeVRZNuP5uQwj/WFeQwWX4imnLDhgpKFmoD3wlX4R
0S1HxPSFnC5DE/5ehir4nhLpBGaHEkEB1FCT/aJp/Cck8rylqLnirlErQpGP8Iap
QYcOmquerkrvXBLg3ejY0slMYpQtUcVT5BeWHDp9ytatVNS5re0ZkTRHtrOdtnM2
TpJA8gTxV6XCRNeZ0PvzlbkVHbe0zyC2XGAfkUGyAb0PyZ84OiJiin+6cyOTy3e1
fjKCAj6+y9KeFhlVJ73j0PTp1roxXhiuR9PFFxJfYsgcxHtY/hW1mKu1w17c9v6b
+TJCxgEi1DWt6iA5FH6/xVhOsH4PSph6Z1ZgaboiBQOg9SRzWZm/fWutMzdjCRkT
FsCyTX/GyhmWFT+WD/FrA/Pd7JEDyfPgbTwhrXHiBp8gOArlv0KEnerQGxb/KkOH
uTO4XsFGvEYeDmkn/GhJryWzXZiJAoJWWT5Os3Zl6sj1chHmXxas30SQUWDl5YlJ
jEkl1hj0EBTHO3yX9foCDGkzIPOFE4IoWDdrug+XuX02UO2qn2JVf8zv0rrXxqJn
g9wiTOClSismfpMUdkatN6C0TCm+xrIA/eCa1v3xCFLQhRD3ev172sQgPh+KMwhN
wGVTA09RrSeGSTQnVlOP3OUz3VWPRKal3O7LODyEmoNoLbgHrS34ph7FJbl6SzQb
uClRjCvPOmdqZS4K/eoFFz8Qs8DYjdMhyqFSeqJAr5ruKd4Szpw5oda+x4Knqwxc
hFdPlkfRd6Jd5n/H2wRI1g/9Dx3d4VUIqQzE6oTEnJCxM+H9MAemDXhnau+s1ih7
rWhV1catT4F3X3YeY3TCBA5DhX+uPZliVkagrRFGJfmixcs5/WsXVohdS/Xw37kn
cD1oA2qK69+h+67ZH9JX2rIstxc4rtmiojxZDpl7Gin6nzNEVgXfKwx8sLGJvStp
DCROv5EIpD4CQtZNBkPq3+INYTcof9jCDjY/TsgL1918C2+b7ZrH2lIORtplY6zo
BczZI+aecUQgCcYajl6wqn0D6cE6TFa6s9eHRahVTu9DCFpX7qDzc9Ba5R/05/Cp
T/JVKs3SgvC/S362+SjeieCbNpbuJKLwzm+iQWwpuoeekUA4mO+jZOftMI36Fywk
JXGTyZ8Md4b1U2gEceQ2IdDRIkHMK4HC9btbgW614KEQOG6BE37MIzYJ75OhfOzc
QkU/sN87q9xudvzvEQ77eams0Tx2m3WGzasaAHhxvn0S0U1bcbv5qX4h2cPuTICQ
lW0ohb9o6dGA5Jf8ssdDY+nmbq4lBbG81VQgBrKZnptq4115WIOldGGnPcFm1dl4
DkaW67vNjI10Gzn3yn2hxoUqmQWvFgbSsNNEI+4fdYACjtlrpO20ILyRXPpVIDnb
yTLdVOaS2l2pVCSC2KUnPZ96kbJ90Hbv9DsQdM/92I5o5//BktJxHr9v23zddVI9
LfMEW4EVNDXo397t2ge85LQb7X56f+2ScbQB5Y0PsCL1UolvICXTl0ybtlVdtXD0
mNIJd/houIlA6rpldD6csoC/hvgmUvbYZfqvIhbVtn2QOxcTgZKbcAbO0H1cDTUs
LSIgyUCXfz9clT/ykFSssJTML4motTDg6lnh+BrTmHkHH461jaLcA/nvA48CaN8h
W+KVDpucc+fC8e69pVR54DJvO/otqb6ZVoyvvH1RA7JE5Z3fQ487iXHp3hRHjH1N
5DH3zqJcXemNx7Zaul+xEqcJGSkbIDCmX8GVydjSwdrA3izmJonl+i2J4o3FqWnK
1tL+kwPBuNfVgAlmxY7fg16wAnvQSD9jXXYkiFgXSQGWVWpE9ItIsyknjyYkJlMl
eacrgQeet9UdTrRy/yv/jJjeLeHAGz6a/jUWvy3U1QxvbnHEQkQYPXAZTmi127oD
0idbIsw7QWzLbLpKHTKwAX+BrOndNmPCKJEsoKSWba/cANwW0isI1iT0qz7Y/N3l
Z5T5gX533X1b3F4YFHiLBDMjA7zhm95wlH0bv1UqydciuLIHspxh3Jnm9r+v16hF
Yrw9owXk6hVTYBxATnCz8bWlSgQWoMOvjslyK1uEsahVD+7L+QpVYqLFx1HKs426
yCJK75cO1DKSTxfC/+4CWD+8TuOSFJUD5XOFSsKS/4GnM3JjfnoDcRjduxTPV6Bz
04XUXHGy/zmv7rXm9A++369TODgokjPacPO04kEvrpxJ8ZgAAJimRFcD7LK/Vp4/
/doJiCjmPjWKA4/BEtGIwbBcooFhEAmuICLacpuknw19o5KmZmvXV8QxuvqrKsxE
aWQ2YixvAB+jMzTpwyXKD0xrXZZZTvuxKvXZEgHzngnvya7/3Jek1Ny5QQ6Kgx0X
GMifGqf4HNJdoIeAUjnBXKkk4W/7Jm895W54h3iMAE+95yYmc759TCBbrn3/bfvV
VvSc7Ga2+dOP9Nc2JPIS6iSjtmpFdSd9h4XMLV2+gYo9DGUK2KlnBbBM670Glxqn
MgViddNmAZawz7UU7KrqLdBxW7noUc30XVyKBbRmVhNl71nfVOdQ2niuf2Vnpx4O
d3URbooUXiJLpU0NHxovrNNLtYXpt4R/ezl59qNKA7KW4pPHC7o/nA1n/V00SorE
FLVZR12DrVeq3qoqkFpCcjoM+7Z4LHDmhXSClRfG8Zutr1N9A+N/PiBTuLtsC9/8
cnU+guo65cpF8LOrQefq0ZKJx+H4567tyZLgNBVAqPBPU6rTQWmXc7nJj4jmze7K
9xNMpLVp5EVTZt3uTOVLEK45UbCQF+nt8I3P/Llugz74kNp42EFamoyFhmSFv/7T
lomNjze6lAZl0PJ3cDbjoidwwo/OiEW5jpFdSLYajDELwiDnBRZnbOXDWobY5Tm1
P7VWPiYa+xkw4TgxpxFQ5VtVGsppvS0rAtSRpUORarNsMvHtOlLGfb8kX/dIiVsV
z2NrZWndH0XYXbNGotjOzxgZVwtdrG+jIv3PtMt7eOpQNSrcSJSPMGvVU/JvtHZd
A0SDl75k4B/bbJCa74ZxGvyGd+uRRxm+XdbQjHfTH3qdXfs5h93t8pYHFmhmJUeS
GautbgIgLlNTgRAXqMmGEq1/COpcmYTZ/mv1X2it9449DkK1G9Sq2MmoGZwMkc/P
PREIgnWM+TxmTBNP9rO1NJuBq3RpEDGmLPRzxuT45eTI+6RD44ZcAGs0SiONH0iQ
HYh57KCLjgcyunI18GNJqNjZ4OPxtFjZ3eQCQzSoeAusYBIdP6RUea/2DqiUSMOt
XGTfI8C1cu7J7SOS5xAXQHLD3FK1TPdbRR0GhaR24O/bjjyhrkM09Z23m0mQAbxA
pCA7eFfnGzC5xWcj1wtyyNLuGkOiP/K3Nytt2tcw27eX+vaVC5cnO9ROIq3WDBGq
xRU+ytf6QGB5a078ASFWJ/lk6FW3Ob3Gx9VFQUaK4xrC8cRTBZJuDoRFrMEExjQZ
Vu0bcoEtm8/UIL0166VtYOxtQmCFVg3NbztY+JD13kLxU+j7enksKw4UdsJ99s9a
qEvIsSSiywBO/lsWmBChcOX6Hany/tg5zyvQll+XDUbn3HaQ6eKBQ0xBl5zqIGBR
YW1dgyq3AAoms0Oxl0y3eB3PNXqVbOLyjQgnyLUsXVrVCnKBHvKUmysZso33vvti
8zuQe3bPfjUBetu6iTztz4lsmuaj6odnUHie04KcOz/nfFHJNidVkYtFWe5jPm0+
sROLspQ8FC2+FQHnIur7lfcxXhswitntD3LKp+Nnb2qyYtcyV2RArz2cueakW/bI
8AxjoRjthE6iZk8pbgnU5WatIVLopoz17pc348Db8xTU4CGTF53/7zv1QX1S5IpZ
zjl5ahN5YGD9v7eg7P8CuJ75C3v3Dci/XH14eFs8q/ITqB6Ps5QKHoMKcNdJAan/
irGLcdnKizmQcdN1W067dldw59tJ+eWDy1Gx6IoJmISwKd+r1yQP5kg48byzp4vP
j9BWR4LHhF9sirR2AMmC+RbZPneMnfvWuqVYFLdL4FvnzU5vckPJlKm8/X56FkU6
QZPzN1kEM6EUx9HFZIMh/0TM+cmFsoqJl8Fc0fK//VNql+vb/Ro46vbM71pBq6cU
kOuo2YW3F0muTs+dOCWPiRQArU5SVrVIOQKxyaX9elvNLRfFa5Q2AV8lCXy8Pyoy
BwD6guO0tdO6XaDV4aGToYZzoHIQqaRWTmgPC6ZL6j4PiCLjAZ0mfx0WeaSHT4xy
OlYpR4e+ouoNgpTjJkfbSukXfVZI/TZcgMJ2A9+J7Ah4YlN2kUQD6Gw6KfwEsuEQ
+RPo0/gmej1bOmSbmEbcict4+R0fVuJDQ0s6oxxOR+/KO1hF1FAdLJg8hxONnEdv
MPhNyBlaDKOB+UkSEE64s//uJsj9vLlCGOYBKVw4ItVBUTpsXy0R6T1xgcckZ2JG
jw9eJejcZtMMMYWMZT261npcYl2KEAsKc/sAR7Zx4B2sqT5bYPNdQ2ytnQN9CYN6
3zgY4UmilZ4AsV401S83u6p/7Xw58BDvBW9XFbAwoLlKRJC9hI0gG4gRG6id/4UG
cDUxBCUh/79a/ayjTASiDTV54hofXvb5r8DFECI9VWUO4qDUQvyjanzj5XmyV0C4
Yk/gFQw300D+ji2LBAEfGVAJr4bCQgcvIUoNPvcBQijDipKfsgr2k0o8ECgrpCmE
Z2COUfn39MrHeI+rRxlEKNawabjpXVdefIn2mXoffLGyrVzWbn1CnqX4DKmlwNAz
tAZO2HlOfkXznxwQKAfRkvQ9YY0EnXGB5I103b+E6L32pQy+aLjDiiEAWD38xyZW
xNE0k0jFHGSB+4vSCkk8yMO95wjxrOpiu/wM58a5izluy9yGLaA7nvRMwrw3Cuuo
gWNLnHDe6VhxnnnAnWCkrmRiEG5Vmyv9AY//bIPS1Txwj0Y5cbtDAWphNs57hvfK
ys6/PhKjYdRq4F+ciyxSn4HuVZ3MAJo7epGwaJb2yMXjwa3D6rZx2DAZBYiHDGwt
buFe+3dp7I7cF2BIfSn7EbxpdD5B94dn7olEQFIutr2AILV2BfEe3OFIcl4ckuyl
2g2m3sIOQYu1/UZgbDuwY0qH8skIdXrcV/FcsGM9VV/YA4oQO8hjz8DXOMRpvcCU
c8k6VPKcc2epp1adtuVoRkS7LT1ENFYpZHUlw5eJVdDMfqsCFIHp2CtcdY5IrWJJ
xrLtAC2wPRMdZJ6XDLfhnp/i+jIWnTAFg4WG8S8Ge8Ny/bzEm7emqoUVi96sQ9QM
hw97GRQF1lqSTZheQCPSwMwRYM66zeNKCKS56Qj3QUw/IXMzAobjqy8+peTa8ZvI
77uuY9s2ViKh4hLy7uUvRIvnO6ZvtgommSxGdCspOIruXBUAglSBP/EHirXWCXg2
ShFKhARqhnskki/iBAz/jDDQkEwKP89vWLPSJYgJMv5pHEM1I1lAlDZKUxPRL3wY
mQ3jeXG2ewUQp2JzZrI4UYx9cWByR/772yJtxv4ShLKYqJc2VcEkTb7Tl7CsO5E6
9RCZ/g3BoQNOFfMqJfyx94BqZ4bQQpUhfg3QrkalCwbYU5wCwKQ3zLfXWoL/KQzv
erKtuco3IUJUhcrlcvpZWWZ3aDB6WrVGD8JbsYvGPR1c4kojv08NfOx2KkaKiQCX
tqMtl4GK+QlappVQd7yiQQAKZBS7+s/t37Nw6XkwtlE/CpURYO+q9YveQHUW6r50
LEP/awbfZJ6OPDavPjbY5Fj163nxKA5myno6ZxS/kCejuhcMr9H094cy0VwRVdXr
Mz6JAi1LPoxXrkV2Xbq8fzEnBYsOteZr7nIGcuq0/sSj3Vm78XBK1knkND6NxK3v
wvhIxzuMJTMwsfujmn/DelOqbg2KY5nirm3oW+o10rYvYH+/gkpMvGxeBkdQfwMB
qZAJCkX8fOG5tSLs8PD1WZWdNlS3++tQ6g+68vmKXLDR3yoDOu2GVyaZnOH4zEbY
Z9seyDgS9o+EcCNb7Dwnb4ZvnIcAxMikHlFUBnB8NOoSR8l5sHwhjrHz3pZC+g6P
v8ZaadNUXezKHXB8hoxwKHmYWygoo28821sCE9hfWgdrhhVvkGiU/0y3rFu5xUeX
MK7GcOxIkMKM/NQh5vYu+1m1o3ImuVs0xJssZKRPeeI/9gHAT0iycthg2j3bfIwK
O0rVChc2mdI87j4apMJKim1AF2N2wP8eldnJ7oD9u++bmsupcPYwmSs0n0CHzTD4
p9xBduw5sHY2KcW4hDqcwlSatXpYhMHQJVpAutfQ9dYVoCRJfhAy2Ae49Zf2ILuP
crTAHKK6AV0PTNUnwndku012PWyIoOx99E1Qn/peCTeE+R6SaW/jL+kEvanTPPTu
pRdFQkgXGIQfo23eEIwfeua0CpSpaU5etaF+IeAm35NA0jGE08Ig0EkDWDWhBu7d
7WyfSIAhR+Flil84be370RAydtJ4nVnznsBztYHew7nHdEsUJQ1iLeUM9aq53B0J
Eq2OMbiXsXQJ4hLyhlq6+9QGzAzlCh/2+ttEkFc83ikOBMViWq0Km149t830KY+3
D/kqimU+2bOdscmI+pJjQ09EjM7/L/xt7eWspiodD/AjRRS4ntlVt+RDPHKNgi0H
HAam5/htyGR0xozMS1Ke+BVxgoVDApTel+h7XgDAZN1mCTWpbZlUIcSlGXBtM+3b
pnR+x23+9P7E1DOncaqzv7uA4AwDIFHSwTrjjF6iF+TvJkPkKdQWixXPqYu2nJzw
5MH6nBx/3HxQRhbOPMpmuOdT6uxQNrGKbTlgJ5GA8DchzBygZ1/RfdVesyE+XDnC
n7voOT8pGRhWAIIIMi0wTuXhE2skYg2GAlinOSMg920CGB61xTpjtqhsilpnvL+j
yHzc45as5Z8E2RbdeHrn1hTiQBJNd9a1X93ow3lGKo8ifEW1AHXk3iGw2ZSazE9A
LmUJa6oBpA43PUIPjH8s+N06Q/90mnlcg9KK93uKSTcFgNlh+LLuHQ6tOkPfHPEI
zcxm5QptZura2pypTf7bMkz/4+bwWX6V1ClcxNN66Bcm6d0q5JISrD282z+cd8td
XZqWXAx5ff0rk7tFAIZ2xyndvnTE7B7ttZTjmX/ED92RqCYnPqzuSIxxgpWImWjT
Ph7thN7Zt3gj3iQYkCyAp0yFfxil9XJHypSZJ7EtBXFV/wfPuvLZyJRI2lZfap0a
1z9hSTJy6LiIUvmZa8cnG886m7YEdt9nuq7vFS+RxhBvG5TsDwVpSW234tJFiZaj
/Ku6QQUr4kj6ssOFDmMjdHkDGYzZcAMVZ56i12iHOo7IGlG0GV5GhSzp6/FPKbCQ
PmG8qMBjDm0BI+Uttzc8BoEU85D8AY1YHgm5OUYpQE4bT3RAarks9cj9Q7Yao8+N
icdyk8h4EMFcKBXw7/q+Ok9d1enUjPJGV7x4NBMxs88nx+3ptJz8yFZpQctWVljM
MegrKV2nPgiw6r2Y3jzd0PCqWsASup9JJvYWrYJwBeQAiAZUbKzspmf1dhcV8AsF
t2IbRy3lv8MQ5PgzTK6F+rnrgOcm3mRD3IEcDtiUWzjtfieCqMNGwNJdBBnbYpdM
XTb+sTh2eKPy3kL578ylYCk12ZreQLWm1oV+aPEjJqnhxyw2eH3Po5nBy0UuPZyq
wqr45lbxBR6C3VEoXhXMgJZzKZVL8pkLS1egCwu621ktcqEyReJVdR2p/LX/iOBI
RUYJEY4qhzEoSud4XJ/wgGBTzZOMX7voEczH0Bbx3Ik70+UuUl//82AFKDR3SyN0
WgPzceXhXYd5U1Rr1zqfrQ5/huXpX2MvCc7YwOpkNNqH3S+Yz5eiaotIbl0KA7Hn
mtTdoDl6mREKYFknIrs4XM+yyB7i1ot08JPmApJolexQOE2F1dMen4bj3VNjuGun
c3If2kRtD9XD34OTANDWuJI9fGyZkNxTPWeHGY7OyLjdr/y67veXRZM7k58noGfz
n80ExbR+aqi1+ovbxDKxyqMM41tz05WkULxyJtSN50hUjxYPV3Wz5vwCA3W6Mb2p
ub7z9VIgGr/r5Dw+RZX25mghnf2moLdOgWTaXfX1gUWTIgG+5w3b4ayZe3/Vvf2d
WZRGh/87ql8kR50CQ2iOBxa003v0qO8TyL1Ey6DRwoaLaHpzAR7QYjqEnYiIvH4q
0tgy9xFgfo4TFv/7hBeqfgXx3JBJgqgzbB2ZsInWCr8FCMXD6Ab5kq7Ns+BzCeeb
fsOi+xjgxpTs5fRLR1xtVfnzunLuz+C/b9hN0N8PjzI3K3L8y13Qn3TRMZ+fZium
3V0wAk5Vs6Sf7zjcMibJtnN3jZY8LW4/kGo6EKVCp+XsnaAPmq7rQBQ6ihVaaINw
rD09KyOu9blhrP5WEOAj/tcVAR7ySdH+t6+MTKv3HaJ683Nsj1KVTdRVMQ1Lvv2g
Tt1Uo+Qm61qDJUJWt3PVp2PRyIXJMXt4Wr9w1hWmQRzBoqEL3wM6uAi/peRsvZ7Z
J1Lg7c7aBFPR+sZLQIWWZY9rGJQ3U2OCmASMtFls7wCIEhlQZQy8q/6W5QEew3C0
Pg5zfSn9kdI+yfGN4VRg0lQ07p8AdmuK6qwJbDgaQLGNKS7o7tqAZ1jSoMZmNWYA
roUAuCvyPnEAIGLl9kJmT9siyAupqnQ1XZRh55mPBpxXe09A2G6MdJqnzbDOfg5p
Ekd1eyJAZLAxnubVN3W2cUK3tb03eg0xWiXLa9tS8+gIXq/YJJxbQHqVqPJtFdP9
IU5lnh1lPHROvUKUKdTAtMuiqQWWwgy3ZnDZshQPuCnOPrKACoeQpwWE2tqOmYJq
aDDxMtbAxJ78Ujl6uBj6yKkHVIsZxLPeIj+uVqk4enrYv2FIhIsQsd0xMKCiqvId
+q3mAY5pcyJasb/ub3HMsm4Pjho1vYdvdaAlqBCU1R7R0cTnD2DtAQAvx+63rGI/
C0OleNi3q4rbR7YPiNAcqGMVDRBrAUFl+eWkHxzWMLJ/u/J914SB0//PW8d8OijY
kU25Hj6cnpeGBlZUma2+EigT6nj5hkfCwiO4I3TM0mqtnLR68+TibVDXIShPySJ/
j/3MvswowlyZHaCgELssQSofYrbRosmIUNRspd8D2KipLpJfIrGmGPKs/DWKPIQf
iFmOktXauJO1UJisUISaqAPar1wY2o48xKR5qlPEMusdBar9/zgFFQyulX3uKUHe
ZwOYMgR9Y4ZWCbO8pZue7v5NEEd/y4MO/2tUBq0TmTz3U9mdjudCc9gVizCqUhdo
YYlrzlp7X7rkMPExUCYqMB8Q2VF8WmtkrqO39HUFEO7prDVKs3e/+pR7GxdphUsr
SaTqE8U2Qbimfut+AdWJlJHiqG8/Ls3Gr3FF7dL1JftfK4/JJNz9nrCDkCkzNP3M
7Rq9gVAGlXm6x0vowkQ/xWpVBGP3OhbfaLb/B826aRh2kI5nspORTTp+yzq1br6O
kyC2g21F1eU0iwHeK+jbajF4Y2mQ6aL/GDMCkqe7kqCC9e0PHrVfTClXGLMVHamK
LFMwoGVjumRG6mwd2zvGbtPU9gKgnK8br8hC9dn2oDrjDgZm/UBrs87iTQnwDE8m
8vSIC7w4vkTWpwya8orF59N+mVVmFnWsHgk2vQdlKwea0qt6s7JuO8Vty3wJSbHP
p36FbzDhUBgngcae9R+obUcl5T7xx563+XH6elVfA3xstIS57JpRlvwThgtgv7DH
hI9Zl6d8kaCvCJmrF7/OAJG58/f+TEiUStK2szqD+Inoy2zsSIKGBFTzU/8cO8cc
Sw7R6YMJvcKVFLzdOXeY7OhOYYpcRVyvnzaAAtEikRcPNFt22MXpgne/qDik+trk
fGizKjTmlHT/UQyow4p3EgYnp6YTwEJup1BSh/ErUvPAQm3UoARWzgjAds5DuCFq
H5SKYYDK90Mg1ZJiV4qppIuakassNPSsptzxU964+2VNJNCs9twSpVJF85HUBD1G
BdHXpcP+WHwRbY9mtaQ8k53VVilu1fkizdtHoprLE87OcznujnB2neTzlz6N54Jx
JCoWvHsPtdsl9OYnS/h3Ii+a10G1ya7SR4mXyj0Yp66uLLCfmZUAMrY6ivY0jFEq
TaSTTFBXhaAE9ZoK1mhfyJeSCWVGyb2Etvv6OU62CF3SWS+x6qofQmXEToBBNouJ
S0LhitFPM4SrZtkwSwbm7ml/PuU7CK4m/CP4Sya60Y2NvWIsfLtc0eHI+kedKpFi
jqqvkSRVIIkX7yxpbkvXyTZ9C+8PJJZAc1e8f3sLb6lwsABEviNAvhF0dimJ+SMk
Ok9Qr9wkPavj73gBJB7VL0Ir6klo3Pa8xoVbM9X61OrF953Yo6k0Y0eI2rqOSk6P
/iwoA140fZYbySSG7LH8V4EtyvFo6crpSD/rj+SEBub2MxPHQTxpbn4XB+VbTkO1
ULz+cmJlF6+bI7Td96UZHBHAy8IzjCUsg6iFL3W53UtXATLlOP70Tw93JyDId1Pk
1j3zNPBtNZzhd8/uML4G5ic//W0opdLghrK56Rn37b/jdnVvQ12y0Sdes+ONtfBU
maeEaKjBku8AP4TAI2+a4Sv4+Gn5bv6ztkNDj5/KrzBjt0EfGZCAoYsEpfLE+KQC
/r3/WgOSxBBimojL0mVZiWw3TXCGGr60LE5VXMofA4Ug1RcPXQS0ph6c9jGfC864
9JSS2QKMFfT1e3wgDFGdh9O4cEo9bibmV6BrUhWIdnZBEOpg4qHvX7cqQGAA/6uJ
LcUpJtkVLWxyN4rEE1Eawc1CPNs1D/8RUVQ2bFPLy0heQiMO842NdD53oi5hKq/O
9ElYQ7qcb9xDbCPzT3eemQK17mMH8f/4QfdPE/jYP9N7XzZhjlRPk3CUxn4fcoAg
5hKCUc0bhWUxNKGlW2inRxouv6x59Fqso+lrbkadQpGQFfoQy9WAJJodewe09IgP
nbLJpjaK/9GYWqwZxjUDPY4NQ28TVr1fetwEXp3UyJeheA3dF0auH8nyQDOXvNwO
77ixjw8ZyBzEZHO6F6qPYs3ytRuxVKb9QuzimB7bML6n4lZovBQDpP73Z6UB24fc
/K6tiLmBv2Bgf7RwTQwqDg51UObtsHlthxLK+J4fCyNlAlpIluv9mY4UJnpI3L7l
IA1c3gs7CFOLT6WfE39W7M/id5gzUOTmfkqSTBTuOazWZxzBtzpFRJ82A+IPRE67
oHne0ARuBKR4b9mGCm1x61cbO/H1wqUyJTnjq6oPxc5zj+9XFQ+4CY/dijZiiRXM
WsScNrXEdrqLgkPQWA8Q6EJPOmmkrm2pKKly8/uW5/UxbI4UlxtQQbfR/s1kUn5f
2q2O1w9NSaxZO+byW1Y5imzr7skcll6KWpyFfReCcH91+9W+xd7bpS4cQLdAP50U
xTNafimpHQ2Z6zNpDPVsJawQ3Rh6T5BLnVpZJHmELErbf1gLS33eGP55ZTMlzVIr
4iuqqy6TTomHbNLyC2yVlaUDGlFOxFZf5BUYlKiD5PRuJCflQwKNcbRjIISRznvr
oiwu3sppbS9UnyzCyfbAsOTHLxRQyYWzA16tyZW637/toCeeBouakZv0IEkOxOPR
FtScZhNsvxzK3QK7CvXizIiPpDsRp23w+bppi8S2g+50JP4LmQSBwyStRIUkMK2j
k7GsV++TnAdouL18CoMvAAKh3NFDHBWa2AguWRbibZSoSZ0wunQyNyNIHF50+rN3
41vKeEXb6facdOeCa1szsw8DrXws/010i1yJRgUig7R9Gg9z5H/wIhaDfWnmXiYn
MJhumQGASJg8w3J/vmvf5MTaUXqhObMq6DV38zjIxAvS1X1f07RefPSI64ztgNab
odD1t++xdJ6503e3v46V091MiXDV0KYZbxG3ci6JcKY2r/xPzgMRGJ31Gu1ZU+El
OPc/CX9CiRLK5BuJPizcACPxyN8904XLIqBC944KfEGgcT5qaZlxsLProdtFnOGe
7uCC25nVns/ajFBpMMhRzxYyTEBh1050qfHtqEEPu0ZsROojPlw1AvehNrdH3oyv
I9J46zJPB9agiTSpUUdEv+SNuU5ql3z8rWrXNkRdRafGo+mMeZoOpd7Eth1pRY5i
QqvVVvPPJYIrMRgboT5P6L74mULH7ImD9dKlzo2jL1bacdqBmn0x7qqUeZl0qs90
TJ8562hDwRTmOx+3Jw84x637ftXI5TH/IuuGgvs96835eZ9NFuKMhDlr+dtBrS3L
cL283jM3uDkyr1G8n1FZU91EiVVH1uQV9R/zNKf8Jfmy+d9VJN0qojtXoYghGBXs
PtJQmhU9qf5lvMZZd1D7N92LpJQzBH8lfA5OJ51BX1abFYfbxhCs6l+8/h35KcTR
sOwO5YM9Oh1iplZj6vgDOlONhuKHnuRapBVlPtCtlM50jGGJZ6ov7MjxM+TVS6P+
Gh8lpcbxPZ6XC7OzjczurmroYgcnCQ3syQHIyKGkxLcCqeq+k9njR4UeFFguyAdn
9QGuQE21uxRjzAGlmQl2qG/avvwx6+hrDzo9CJbKcngaY4P7hhfX4eYFB+BLKeBV
wux/PzWJKv4Y0ihZafeS+j88gtpc3Cpjpt+nPQrMUwziVbhSLi7kBkC2KpifceUT
ov8t2+APS0qgsrq1UXc+hYfZLV+SL2k/D3fr1qLB3lefGUZMRBrF6lgZfIXyPKfY
PKxIVFzlzPEkSnMHvZ7wwRuBghn36DfKTVKPhx0N+mR6drMHKp2OVIoJmmR8N4jI
d+eo8KnDQsEdYdlkPBUnlkXJ+LdUX8azbrRZg0QDBQmma91LEm+9oj1phuqpm6N+
hlKZzK9vCG8gDBrf6sRS8Iia3TzBr5jj3cUwo4ndECODl10/bOuGtCusEkE4dyzM
uNZXUfzPt8OSTbGdHDrNi7bbQJdNbllKZ1NrCUr6CP+pPFHENUj8pLOxjd6xQSaN
dlaMJ34AXlhpyQZmbbnIuLLYrkrDp3JyRzH2ymHWL48aR/CFz0a6q7xB0HHONaLw
vDOKXpaC+H9mucEwJCEXweIl8vTnINY7EQsTcKg3APLWLdKYZ5OmZLqt1hZ3gFS4
qSObYlfYb7cS0E2QSs0XMnPR6JSshppxzNXAl33IFOyALR9ztbUuBgecl1yhF6AS
XB4YdzfsEmeih669jTbWeMGwoZshgJqIJWdmqIUSuFxsHyRYUeqSUZ+jk0m90Khv
QhJ83b2HVNQx2Wc+FiOjEiPAu5dyAHTYwiNIrahKG/z/xi24cOR1VpKOWvuiCOeb
04AMOw6vdaRl4v3sF/nsmMFeiMbmzGy9EMLBB35tf2ymI2K4+ywxnF0h/3qKImAd
yUUb+8t/P5dK4wqGDcw65t/4zbdKW1VIxq4emsKLP0h5bJ5L6vTEwFilpPaAZrI8
hAe0Yyf/Iu9lJzPwQcSgNXqsBi+fUlJafzu8dz1s/BbCbVUkyRzyXMju1LRK1UZN
XwhEg+GKd0qtCfPAPWnmwEKZN+v/Gb7p4o+YLyFhxeSwlMHX+mTGHOQ/6wcNiaNy
q2JarU1AsgzvFGtzuRSit66+Igzg9KItldwvTOKcvvs42Y+NqwPGLCOA9o2NnEeN
tq/ArptMCxk15lLdo9qoUzZvi+lHrGoZ2xGDPmjycXueP76uayYTPNwv+t0ccuba
etow0yX6gwDe1ahnEk5wMWtJ687QqJdPNZYdcxcwsNUWNc28MWjRnTqhxHZDJFWv
IUj66CPNVhKk83+vsslZwNoj96IuZhkxEAW2CbuEWPjHofTuvUhJLYyBQ52tWfvs
dZNRrKbxWj79r6p8EPn7Z2oEC2wyFgoEziaCsPBgXxxxXB9rTmCUPAK2iPdxrNPj
VokPTb1vu8W04QGTfv3nzkPF25sMghpz/a6AWdjPoI/M1O2Mub7/UXk7iLHMcLvh
p6Bwkvaj5hxtnybwFWOfy137Juj7VFLK5aDBZtBDE+70nVD3jI1RrcQKkWZIl00l
QnmSwk0/oARLZHrGA8/S4j9ttsvujioR2Lja9m+xz4kqFmfyJf3cpDNL2OI4/vAy
9BilGqixJ5qbdiy0lLyTAy6ekDZM7upoW5gOLTF9b1D5nfUZKS1HgYfwFAInAdIN
qRIfpw770EPvobuJCSvrGq2ZF6ucB3mNIzL8U0+uhqPK2nxWp1Nd0ezjhHfkExOC
7KSYf2Jy9IkpG3gxOgYla1bhMzsSRW1Wccn063GEm8cmlD+ddQED/cE2s8de0O2d
fsw5VwI8PHBuYiNCIdGV8NSYyfGiQV+ACvIhEUX8hvahBCkcZvGdGr2ytch7PrhI
BfhYEGiA7qvKFbSN7an9qHpW2aznHkR7tU9IanS+4pUdQYFORMZ4LkBs6dguiEYE
OVjf7r4/AfC0FUe82ROlkBmbwzH5WvECzi8AWghdJKW9s53fkUjwlghnwBByLO86
foJwTJV4br3DuWH04x65kcKHYgIu1r97Z3Pnr/wefNbjlnZ+EDcCUVhB23GFKORf
5ckcbbp3/ALVKVgvP5cHhQTF8rdSu331Wdx8YryLnRzZKLVYlUFZywhUeXyE18pW
m3rvQNa1QLeU3MjiSbzDgnFEJteMWcVQ0NF8nLnRNSXo5kr9U0vzuRMU0Bl4zY56
h5DSIoTdcrr5NENepj2mVu0JSvm2vg+dhvXMMGPTrs1eXJA5EXYwhC2qd1wn3NDN
ng+bo4cSWjX6yfaOkjegqlVqGnhP29/atkLOml0k/X0/BDR8O1jjjjsazHBJoIOa
dlCYaQh9EyWTqXztIJEOPb2+6iDhcVdItPoETOW+HvgFor9ByrAcsv/75gEHPdrA
pxFTJKoY+cbW9gUOy8U5sqbz/zTwz1DBRfrrXaEdDfPCtEqVX7UAhzmjK2wNGx2L
qVsA43NF5GK5sx8GWSIPDzFNm5V09+fzLyWr/m0kakFQyuf3U5Fcy6ogIuTEofqd
mU6srV1RLpC+U7PUFBPf3fvWEwAN8kPl0dP2YAFznsaOPc6plhg7Gn4H1uS08n6N
ftYf9om4WBueXzoNnBWdyk0wxyoCpainTsb9NkPWwjPycg9j6LVbe+1XYvRbtdXc
gHc4uffSydfQnHvFxuwTNZxpq1JquqkEGcWDlMsk1hXiy5rtuz6w8dDBxlt2N7d8
hYoimknMMmCtuBX/gnBD/SlqwoLhraZfPqnxhew3tdKHovPASdv9ht1ODzOOhcNT
UeSuIia2aTjfdRumSzIKjjCJH33siSJ1GHwKnnpJbFp35Do8dn3XyLIMnFAkYXV2
2DtD006RHYF3HZgxSTd5MmCb/S/rs1JcJZy9q3K1TqF6LFtV+upcZgz+o5RJkQPo
zLvzTSnPau/VPHGQSuSLaOs7DQ0aa53uV4xXtPRiF+6X5u/VwyGnrJJlzq7WPz+3
XNYYvn0lTOqEo/0VZoGF5D7/Jh0gg0SvP02Ksj8iXm3Dnh2yor5xH6uI9ScqqvTI
qgQQsR5ZFcQWBeKs7prsuhcGXw4Z7aHLuuNE+h1ZTl3kMzuxqQRPp+LoqhNaO9YI
rvJK3lhC5aJznv2GW6sR6jplJGVvlksG8h4SmZ959tlU4FDLbD7uyZit8YZn+qeS
MmXYdzbpeHeIAU/4YdWpfVr5a01oIyPUGcnr7Cmi0uhjiqMUK9K4uJFqlG1hd+sk
uk2O/TAom8m4keORPepsNbA+mDwY5CH/zWdJ7rxwzKdzatxB75Jpamk+KGYXIyXV
dSOmv1SIYm475wP3ZPep1sBK/sF0vY3HIdlJFUC7X/kw7+xh4ptjedJ5+gqkHtDP
4QcEtrHiWZ4cpQlSQN9X0X53KLWz9QLk87ns4F1HdMfmwUQJDsSYBDhqHc1kc2//
TK/b9UA9lsv7xy4XC8KgHqVWVgu4n0ZOuPBQsBgV35LaxoODUkJNST1cM0k/XHkf
gsn89tIJs0y0/ocyet51pBlHUP5TyVth/jFthvbJVDuHvzrysRFME81sAEB7GKNP
T2Cqyl8JKznFzTz04z+7HQcgFAC1WpZOeci2Pc4Kb6DpIRCgZPKAs7aPBjDP4JQh
M1Wt1A0kuN/f5dL/ppmZ38sbe4/r6yyW/1GmfEwSGfSax0OgNLfpf5vgHS9duwE4
cCKrweIj/vLaCDrZhkvjKDSeofMqSPiKZ4zsfzg9ugDo+VfNDgh6GlR9aFvViTOF
3IATj/7uAX7ZpVQ8FeibuiQ9hknT7DrqMo//j7qvYBD7eZcjrL2tLnivSq+cJP1D
zvOnnJOVSpHJ0e8HlY8xSs76poAZYIHtOOvY1n1VFWVCe9apTyibzlrWZkxlbqmO
Sqgp4DFRXYSGHz6LXwEphaphAihHiJ5gCZwcgFp+dTQJDO9winkUBeFJP4C3yIRg
XsFh5VIxGOkjcKWESoD/pU+tAYKFX4/O+HpWoV4FEdjYe87xh4rMtrGnxznPZmpT
vusC/E5J9JEsIoLNY2PPHuKM9qlXtki9ciT0SvJ7dkGJlN/9PH7jZdB7LAUYvWi/
Tm1kj7Y7oDdobm8yMspVvcvm4uJuy0/NUcax58S0Av2ewpr+2gxUgR/tW7V/VvW5
KJToFJ2YWhr7V75xgy5nIgvlqS6ZZazOcYxBuBHLosDt6t2qxf4HZlpSHHnR58ZD
jN4jaKO0PPcVJxCLz2ewS9tLFFgrASnXss+bBm34iSLVlLQCbAc2Nt1hRxgBqbKB
n0Ddd1qf3t6VWTQEpCxdHBcwj5ed4O5yGN6HsdfTri7/SJIG/Nkc3nTo8L96nuaj
CLJFNhNgU02Kvjv5gyjVQ322D4qVvYgAmKap6qJBT2/rBIHAifwVozPtJ+FQtf5n
sBECi4sFUXzTrs+CEppjp2oTwJLRIhegDanSNep4Ch334q58AqE4hQaCyJTs3nBg
ZplQ0dIr1DPNJgrp/mwxerXVRXieOgAEI62OUPS4Wh8uqh66j6bn0COOE8nYKCCZ
QAcgBeW/kBGLIfKJQS8qfYBH2TFrf++QzZfey5nDTnENR2jg/C7Xa92D8RbOvP4f
/4NHR59/a4e1ouC7uBT/BfTUlQZOqYDVpm3Jx020+Jy1STur8LoAN1hp3qTmsQ6H
A7MrPFy8Mr9pc5VVvvSkCy6e56GodwYP4+fq9dwXvhzJgnqrLDU3YX8z3Tt6McpS
A++tQdlwtylToCY9C6pn9ThM0ROrXsUSVEz7ApDTT63aR8iUy0hN8p88r7ibFz0k
hLDiTgUava3J/4T3+htYFh31bIFPelDGbyfI7X5952NP11+nperywPNTlnIj9cvr
BqNIjF7NG5tlE/mznHy0kCxnEvwvJs8s0Ojg0BKN5YMXSBKnjRaRIM4rLVOweYsa
76nQTMszMQ1V4V0uXb+wdP722TTpS69H8VSHNz5qQuCTK8htcpTufbpZxW/mDO0B
Qr6XasLWDhWMzFVqD87Tn4RWVKjHqHVBAEVcudQzSWvD14w0+eIOopKXFGDBrR+0
cujnunjy+4+w6t6eSUVyCh4eeEmpj9zDNF6oqNIbs+0KhSOCCl7ePLr3m9+WphGr
CMkK7hfjnNYIrjzwtAQf14KfN0zJEG5Qn5XgbBb+nezzqitx3VMqbryMYTxJQvHX
MPf3P+x0sLVMkiVWr0X2S6JDY+no+Vi96JIX0RhOLgVThuay5V+5gTfjB3gkod+w
0EVYaxi4c+CgqOhjl6FEfs3/o7VgMV14sbIfqwaR1R/gaWYOpgVPfp6pjC4B0nJX
JVddQkXfexjxLNZQtX/q/5m2vLAAEttSHdxpiJASMNaGGGmp7Yd4Il2Q2Toa3Stw
Ml+wNlYdrSR8Qg7KqdICwqrld5szw8rZZcmmoGv2XDAGwkVdRdWgsn1yK8zHMINp
I+qOI4bRoaiMoUmtIm9/iLtAFsMAdvX5zMGMMlw+N591CtX9rE7RgOe3QqwLOQAn
W6iEFsxArybAyOWfIbtZ94m6CV0Ne3I0OvhzBY6tAQqZKEzR6hq719zbmwvOBb/N
ECmATPJdApFB59onfqu/iWzCU3B69V30uoRJuEt2bRZZcaQ+YtK6nva1VR9G65/m
I8DS7dhAzmccDpGDiY2lwAC6Gzh6z2PUcxOsR7Hr1+Swxl+wefv7JxA8taJl0/9s
A1yBNU8XUTtV2s5ElRBSyvgBH72Oj1GPq1HjKqsu8DFYWWsXS6pvDKBYtaUpAEgr
bPqrJhdcfNSv4f/Kk3c00ZxfxY+6sr4NyPUn9bPnorRThXhANdmyJOp4zHUruDlA
1+zCxiofyuMwjuIQwbT7QSDfMIKrERcfQBovF6vw7tCRhzJI2VRBumtAEU1vcKde
OP1CaHbxXhnepm4nxVInOcorvQaC7U2vYzuI72In+wOu7w4TmIIUz+4kIsfHwZGm
4AQT9u3YnnPD3KXUDBZRVwWSUQoF7dtVPD+q2teamO7PhqvnSqazz2TWeEoDliA8
8qs2qEC8IKscqI5D8lDR3diD62OZU1HHfCs89NBUvL8b9U9383Xl/wa0UeE9SUEe
NT+WJpcV3Ti/o/ydCZf+5T8dMkeOdbbbUJf9+c1mvlr/teRqg7xygvysieJ2HbpC
TMX3m/ChVm/drjIwZ6aYQUavIGCmfqHFIKXWJX0f26d5xXfoNTXeDLQSKCD+NKPL
LZXtEs9EMn/njg6puuxoSxJMg8/VjD963IvmPAb659c/C1a4rKe5Y4nvrQRdfVBd
DF6n4P8rC3u7ApWw7LTF5I7dcnI7QMDzMPPdegFnnoBvqNhr7gr+6k4Rme1E0gOc
QYV1wkbUgd/gJNA0zJYeWL6Ip3Q4MVBWaKi/1SGvwyNYiZ0Bo3r8VVACMPXv9utC
mf4DNFGSHSAwopQn7gmdNXdndBp2sB2NVfGedmZxLxcrks7QRCwGEXkBluLNCLWu
KdOb875i9RLuKVVuYHSgcKN3ht7Hc/VBH1javCY7acVrBU1rczgEGFZxs5U92dgh
MIxjKjDklw8dixg27+X0oxE1ywxQyYCw+geZrnTtfYbd24Xw+ZtEz1iAuUYC1clD
e9d0AdUr/Z/93qW+EZKMe+Pe1rkwdkmsDxl72cYIgiP3Uzw8+5eyhfedcfeBjp64
wZkswmUMeyEiPv6M72vESbsjYlU2Q3CA/RvPup1tjMcszaDd3sSuAWqvAedTenpD
21ymRea8j6fcZQ96A3r+MtlWf3Cj91MZyh5feAC5yaRrb6cbQjV+TXXsGrXng0+X
nF7e7ysRlS1v+T2b+9B5lC9kF395QL6rMByTgi7rdriJSqmtL5dlD9SsGOuN1IAG
2m5j+Spkog0JHHV//BKg6Z6rWKw6GSjR4oxVmUywNonL3cFioqAFK4jm6VGPim4J
OaidBCAe9uLJTR2mydRzr2OlQz4yXp1Iq2IP+EW8x0ZK+ht8o5FuxE6Zbvh9OD2B
92DNoGnI6UMJq/fSmlQPCT92hDC65+TKGJz3qHPk6RZp9a9meRrCSuRDo/UcQTc5
LkzSHgzl66o0OwIY0XVDByT9x98baNKjDiXqTNw8vEShAMkJLdMkfvCyVo2oo2Io
I4ielw5SSwzyrwT9qr73Wf6hOsDYocVb6bMC4RRMcw57hUZKl1Fj45pDmsYGzT5O
0lEjh3AHU/xtKszTFtlVunYQWfVIXf+TbcE2sFBhHaAjiM8mKwehCaw1gKrBIGlw
dCOB34dME2alCjPdHnjz6K9Ci2pKN56/GS3QLYLnGjrNGr+HLcKadve+bpiYqSqR
6YLejR20+5cRQRwuKwn8QPel3dFivaBkI0Wstd+dq2w0EXD1W+pFzZyVJ1VWLUId
B9F6sNKS2oHgk+iH46LXgwXwJtlz9VtpHygD2ZbE0s4lB5GEQHEDlSBoYrTz8Bn5
13yqkQH56pxbUiNfextzPi3AayEBn/kqNhhO1zYJb/vPVnCiZGdqiJ3ps4bl7jR1
irEf/hTVaQWQC1ZBhV0A2Bwrv/b+4twqK0d50Bh4UagShS24Toz92Ew8Y7f14zaK
zbXpP9X3XQ8xE84ANRCm2ZwyDEhxl0cteSuv4VULZ4rJ7ajuenqrbJh+t3wN0I2N
ufRQJAa02QILq2f6vfHMfrPzUk8AMf1OykRv3ormDlq2oNOgqzO3CXlaApSi2px3
8Kb/AgXLOCKRDg0zXWVEel2WEsV18WxJihB/OZW2IGpoukwdiApbZQ7B6wopP+wI
J2UZxbibqgPWmQK5hwZTMEvRFuuuLNwXTDqHvvjdNNnE0Sy5nfS/VL9Z+so+udQq
+oTkh3YH3zO9jxc89Fb9/fK60ZJp9ctV6P6HAGgXHn6230JoERaFIaghwWXAX2Am
6ReIwPb4Mk2H+wgWXdjEMAlI1hZ1hKYWffeyMF1Y9iJX1OlIVZ+u4sxNh6YDbMs7
Yg3Z4oQ85UfeKxsuugh6yC2xwLAYUuEd0MgSOEx8oeGxdfIN2n7X/5m6IiDHMeOw
Fduhwi5u0/aIYd8cxtjfPJOCrwFDf1aabm4J7It7xBsGhvxwWcDU8Ac6E3IXGo/H
G3tJoz1vKOxBgSZk5QGZToqCKOhFVQu3aSqClYOpQ0901Gd2VbiVOLfRC59D/uIo
Nh55n4c4IH90Bav4xXK3Xe5giMcSw8TAY1xPaxJpCths1IIVLUXEhYz1YHRJSZwJ
fO8T5tbrOYDLXzKyjxJ7ucWBTE3CTAFMUU9Q9BcgDidisKMQYin6aRxxt+iyEKpn
I0sNyAbXfgF38n3bm+YyAfvmYKlrSf8FdicuuHF3CcCpVSB0sCbj9g5TH9Bn0ns2
73OxACacDRFmmoF8h4bZadEpB277yPm3As76NiAcI1pkEf7FsP/q9rbMFnQGixXe
EewD77kyhPmZ8FdOREIQNJrP9fgIy0DHPeFHaK/dFDGcEZF1smhMlc3Eofd6g5Ps
Dw08D1TVn3bd/uxRz92z7wRlWyysEGfaxtlBwlr3Jlz/HQTV+3iA2fD9R3rirMom
6MBrtLnxlNlUqeemtemWiLX2QlwrlpFr7EetfI+X0RSyl2UmC1egqS+q4NUlvKJy
M6YyhYQWmUbuUBd0NTDC7Se2tNWzDB79a0lzexMPOx+ypDEEm8LoB+m9wueGITFf
hWRHaRDuBlL/iS035xW0xBJpS+2GnO4Naf3rrq2dAwrSPRWiKENb5hBkL2EoxGCW
PdMi80bbQIC5YuHXD6LIzUd0+1gAKOvZ6tTzPZ9uCf8evvl/0lgOPe99bhUpFgH8
KLDcdYy7OJc6tGsn7eGOyHRaRaEEj2KwuN9scqkzMUjVRDcxkF1yS8UtpCOLX+lX
YQu38XvlaHXsO1w2aszsmi3CyvYBeXLXsBZbnvKyjcdgCivbH7bcKIYItYXl4tDs
ZoVABKYpl6wJRcJNgKmv3SbASevH4ftYBFuYi4DuB2BtfLjWkMDTBxluPHR5Xy9I
3ZOUDVTpErOeR8NDzZDaYL/1YMvtHsPfz278ao7YE6q4XdV2konAcYlhWqC3c9B/
51s0ECunzQhhVq02F9jd3fpN3k93gxCVsbgzk28z1HytaSvbHUw/c9/0Ww9b/p/9
2vlN/sHZe0NJuVAkWpk4EnI9nX/4YOwu8Eu+gQw16jC+MtK9Ac8NCatbGtwkOLJG
KSe/yMEi16ClTn6+mr1ruORMJ5hRAljOIc6OR9jXUYYHP0AIA+1EGjdvPWfui8Ly
i9WasRGJKzKFmqKv/zlXIO3k4wCabc1MXJItLrm5E70sofw0Hhs5+sceWRtH86IH
JKcQ6fkTVV51FA28jAyAVG4QD50AR2Xtc26SToFeS3d51uRNYaiOx3MZcOB3wEgI
1XTRMirwHedvgmEFbSp7AY0wEFbPsKw/t2Fr4N6/1CRE2VDgvnocYd4TiuXIcmfF
fCWEhbS3hFoVud0r29NSzCTmIHSWY1B1xskdfjG9slcvhUNVSjmE06h11XToc3XD
gWtId3BmyaNygL6tVFJUYsKU12HNisuQvj3hDj2DT36tXYV+mGzKz+3Db4HDkiqv
+zdveDxAsyvHJg5tmaspnXl2y+TibaJgEMMBHkqT4OOjfxBHRCOFUJ7vP6E4BOpi
8PW0K6JhRatyQk8HaqIGJkAm71V+k2IUTMWZs3xfzSCCQ5jtXCeAVAlahCXXMVzW
SE/kcccHCBLLkCI6G1QJ1AuLlfNG8Web1JjSXsJZ3EWR+f2IZybmfUOqu4O4BXk4
q2kysAdfS3iJW5Ejso/IdLWuZGF+25Cs9tTjvLD9w4lwomxdRhIh0X0zsVobkFjG
4TdiVtuBDOrpMrnceClAUUV5dlus0vvfVLWPLjOvw1JUQZE1//vm28g+2K3G7VTi
omJVEQkQ+NXxygpHzUA2IXwJe6F5qPLXIEe+cG/RITJDacZKfmjo1GOyx0Vjhbkc
aSOWc2xl5tYZU7jQMrInnLUWevyR4s6WtHi4DpkSO3XKdeKRGu6slGrrpS0tbMTM
HqEyR/N0qpWAS5m5vsNqlhMR6NS8joi9wh8ibNQ1u2qZeWnyWlTPBAFVuF+zKAe5
QovL/2CtRsaJzp0AGEEtqJ8XIKLgB0A2n3TCpsdxvZnDXcvZbt94gxO/RV4iCMk5
4Uw41yNqGT58CNdP4DvxlHNZllSlW6u73bGO3/khHqIXwcZEfMUAPGpAPDdgkxvI
BXKmZ3nistMXbxFSEFOP8lL36TulywJhBOx67L5rCiiZpDHiwFuF8atYAOV+AW9a
YKL8JCtbzE8ZiPLADQGGjC6QjD7+klAW6xveKgu7nPNHHxTwE3KSPSkobTV5Qdr7
fugO7LfqMUQ4ISoL9jtgy91qJ9/Sf8ZktITp1VGSm6Z4chQ8EOy/c8qwEm4Q6IR2
CRFRVR9/NT96uYrIlrhF7X/ANkG23KSXjW7zc0ziK5B885lifZk5UugSYKU44Gsw
I7fvijAKNW7Jhb8HaAsswSCCvRITGxElX1KvlTOamKFL25DiJm98H/QEbcQrkjO3
QnrpI1RK3OPjwQuIFpfi064UwdvvHetEcmJWHU9ScUz1mEnDYGCEuAHleVbIJB9l
Z7tJXymLcr20vdzI2MhPopd6R66ZCZw27r0BBjiIJObeFcSYw1xDvT707YankUa5
9HkcD4EcGoxjZ7u+qszo3dyFf641nNV+E5D3G6jxtdGzuGZKV3rYy5uH9Tsex9AL
RIeVrJT/XBmYqFS9lWXwDbErKBpe/6sKk196jmOoyaholXOx2Us+PmK0Ewyd/Ev4
iqBNny4eyENXYjKbNsh4IBt0YvMQRiBS6Q3C+SrqBuZO6wnsSb629lg3dqZvlOrx
SZnduf95FJOrVDihoU4IFA6XZQe3NYPtyneJ3BsqJHHz/xnBt20/Fhp1+G23rhIk
6yCrZH6JkZ1RZzC+E4VcdaT7oAq1sMnkNa7zwIyJsmaPqq61pyQi3yD1boDWB9bF
biHoSkguj6kT6bqVR1/dEgjKkSzf/+5kHKBbBjPAn9lFdvFcOHt8B0xnPln41hla
Swc5gTKNrYwSIDq2bAEfnXNYBUaU2qCtCIMVnScH2LBGkxxPEJBdsYPYy8Ve7U0M
bh8Y9RQjPV8ZMAEvpiBB1Q9J8nN5uASsAtxDiyEQFFVn18cnXuKsG4/CorQwq4wM
+YQu9IKRWXsITME6ufhWRGSysJLKhKSuqNEMdauWUbhVIc+h/JIJIQR24bWlscYT
dULamVRGoKZj8ZDd1C2Rnx0wKFNGr/j+TDCmw/F0NhD/LFZHKuXej7NoNkZ3T+th
gjDH1dfmBGk9XX12Wm0lr2DD/VqOVihjNMMgyqEpActVqRcCs5vzvTLq15cUm/q8
r4xgV5R7j16Qk3cKBfCHKRYJjpHWgRoOyaOp3mzKGclWTadyR96cJn1vI3b0I4Ui
1nrZe+0c437mZYoNA1jylutXtozCb2yqgBUtoGlhpgwNyhXbacwVbp0K0KQzJhmV
CLb09174o3p3hp2frDub2N4YZH/aE7rVTyXBChxC2uIqYbI0CDjYgTn5OnfAUabX
LJBT19mvx1RVkK1U4/WWqyI/eOtQXQEDEiJ2g8D6nxlPPfZ8Da5Kk5rFOy65Lmw2
lmHaOiRR3Qu2tM7eV+uNRpj8InIkbgW2+oLl3CaRJTbsA2MGTAgPdYRsT1LCMjFW
hEzjy1JFUAIPXDGfoql8PG62jqz/x0L+o7jwhl1jwu6yfwGSH1SOm4qxyQ8l+IaB
YOUI6gd3tnqC3IfdlfMZZ/9rX+t27NNnKc3MgS8fLDjkUu+6MFtgWP3A+0zq02K6
vF+lDUjLOBIhJ9vXbaugf0GtHVIKZprzGLC7Q2CTYWVa6EGY8cQcCbkq+iqlDjIk
XTqZqDal6P6rAh7iwooUIdq6+b35F5MFIW5SP8tQMhmlrJAFSHRwoKAPn4hMa3k8
HlNzPVzK61PElQPw4g2ColS4wDl6zwOeyMugSdEBQyNoeCyN0OSWBwah5VwO+IVC
3iI78x4/pKkVKnYorwSMSWIJe+ZGoJqm47weejMfU5xPNo/YGFQ362LRTB8xsG6l
RRcWGAhhYtBeap92ugNwkXx1cvfpAAlVps1Zz3iJ6GcZqlzxgpmw4LR8irILPvYI
EZjNvVFlUcnYJJ5rivP62P9d9d8aJAL0T16RE1XUgLet1KVAJg3r+fFaGyPNE5YK
5y5gzzi22rVKwNoTKW205Y3Xe21ijkdfAv4D1oS4IcHTl/Gr32mxvdQSrP7AJQUq
Cu5aD6YG/1NVFMCCxVjYDlUChEeDyB4ILc0KoOVMArzXHT/yvN6j3tYrMUvBnVkp
IgCQKBrH6q7kUTcF4pyhCKGj6UjMzg3JbN1oBxYtjfk3pZgHuxP05rrvs8buvSNL
3Pt04hOw+3iLMXD7WBZCPeGw+fB56Iru0o2peayOiNVyxLcu/wdGvnnsQD3w6QM/
CoVS3ObIUkgzNltth3N/c9CEjlhjN81H38Csk5E4+xKEMP16i4TtmCzR+kPT1PA4
vTJUx/mY8BDSBrh9+2dsWqVq28iy5TkAY0xgtkcafovtETvxLjAi+3MSoj6lO60t
wiXFl6y/4chMwir9Ka/RMLr9fq3NJE1+uJQ04zyc3QlH6dGgvBlwvfyAvJrdSfYq
xDW5NTVObzicU6kne8o6qEN9rDvmEXTnJ0s/PRaaeQhl5Y4A95m6Gx8ctIUJuErA
7O/6ouubqy97rm9IFJfmmGQtH+jcWNhdkkTi4IqjdIzPL0H9th+ygpVuqSc5RhYr
adz+w87l8bCXDYAsBWZIH5Wh1tArKK/afk4664zb2sWFYR0AhmT91ikV2EPACF2S
nLF9fzyL6Onuvb/+bEA10wpJ9OUqwxshKiuVmAgZrCqzn+wV+nXHCSVL/Ak0Yu0I
jv7K+HnopLFv8F+A41SXIPsY9lFXzTy2gMWws1sFY23p4EoUTcegr3G2eQUTC2ZL
5ad5lohcKYkyronoVpR0JAohbAwo/tETseBsSHLOWGysj6VyIQVnZ4dmFaqVe3UA
jsEfc6/j4cNp8Meq7CU8V1yv93CwY3Ba1R/peVIqAWI/VqHEktM55xmuGa50LG8a
g4ANeJnZd8jDRM2zoqLzHHl8JQNZ25JnG8fiNMXhLnfPwOfR4L0pr+RuFI0w1Tst
fD6TygavKsqzDVHkKiflG4Iwf7pA4ZPzg3WAGgRCDbbXdDFjfceCH2/ziCS4op88
3S/9JDBHqPrelW/HGO+W9GKUQTU2u/PFtqgL0O7ScB+W66A+sGfDP/3OA5jaJQGj
xOF6M4RjJdkF8ElSVO7pohgtmFX1f3Z6FOFqXF92GFnzhEmRKvyPxnvKdW5UHYXq
8tK89/IidsuKEfAFKiZFyRkgqtPozgg2W5QVAVUZUzzHrC3T8qYt6AQhq63cXcub
SIw7rJR38mAmPCEo3uEVpIcMt79QJ1FMz8RLXn7E7UvESEvkL8tOBEpqPpjQQUDn
hakAGq3GH0h2JldDex8tU/BcBexUrHYXjsoj2mKOwdlkYtQx9kXHwQ8hnob7GUqa
oXi+WPKWy7eB6RtVWpXseypiU8SgxNXbkS8OJcMxNvHvHDyn2eJtCIWPZl48Hnrp
+DzisPnYVNEQ22fjULdKtClxjfXNDpfmGIbJ41ipLlhrJVROd8yAH0FOfmt0rKvh
qsysWzjpJ1IkrHehof78dPF+mI8OKFdc0hOWoCiM6qAl9ZWtEZ9d6zesckqz3Yci
8s7nBtuLxt5di6BPel+t/6wGUXaHzofO9ICkE8hhnyAt7+yW0RLYPXagln01HxIO
G1GFfn/3HCfbkcFfuspjnve6G/fQfMf22kZKYWmJBPRC6xtb54hMOjYonBO2Qw1z
9ovZWIXyAW0sdwf8MPt/x5riRhHf+MIMCd+9hDEOpioFI7cnpCPGI4EmtvwYfR9Q
baQ3IF62AZBda/R8ljupiU/Wn/VcZdlW7ONtiVxSFvXSS3zykQF1QCUTl4UVXej+
9yBBIJGwrYnao7i77RGSLn6VnoJAlJEIDOsn5oFnWof8NZFwmxhAlP7B6d5FIolR
Wzx/cKt35U1GWow/zhSLvp2M3oZ8tSLebggBq/S53mlEAYksKmykxGwSwElfpJYR
1wPg0ANknMKtQPDw2UtaBVm9G90bXUHi0oQ8nel5pEJiCm4mflUFJrqXfZA69Syf
tx2uZlycPOzcwshthtunesIc4J3v0lkJat0Q0BBYrsNZjkuk0tYQBJv06ybU8974
BFSXWKUk3vs2ezbyO12ZlAZyUl5NhqLTi2Uvta9AB0azA+Xmae/55Ygnpw1Afk8+
rB+Evuwx8Cx3LPWShmul7KzNfoflXWHBgymeE0CNLxhqnx42qN9Tddc1+C4IXUsB
8l9QqZrCIlG5srjqd73AcTISzWAb6gGxkYEp2RG5gNPyGSktjZcXyxJbzNB9N7VO
UkapGpKie3UCZhYfHBBFesuauTZge4R86zivss7TLJI1LQPXiAGrNfSv9uWySxHx
ChaCruaGM+iqXpm5O4A0RxQDQEl3XbxMLXz+TB8vAqdcXqKpy1Fntl4n6k+Lsjo/
+OEOAUu/WBq7ut7y5IQcojYtO2iorGmOrPAjYquxZ7qp2Xc11TJCVkdqll6jlWJC
A2rvYI5H2+7ud5pYrLFuGL7oep4vmEqiB6ttqCam7ddUKBlmGJjQdH6R3tSoJgmm
8cSl6KRq36iHhW1AiYTt8TDH0CT9hDVD39+1hRgQGbCk7ECMs2XX9JEtKRvFMlL7
toRm5Tf8OG8ib6bHIBF457y9HZsTlLBTztl+/GHE83ehYrny9Q1LV1UnKVLgTOX+
oquKdjHeV3FOFuqlFONrG/CDZ9aW74BF0njQryckOfrlgnsD1cxgtVd6wayQfwiI
DYkP8xQB0YJxh5gpm6bsycyHNzOVn+y2Kht5uXeTK9moUK+7eq2g/lhZ6IF04ZTs
tuquu8jw/ZRX5uB8CjFeZsteC3hrEN/ruKux3iWNFxnSmyEptqFlN2aVba9KhmV5
9h2q/RV1aEFg7Tzy2Kyh7YhN0oUhpQ9/JGSUEdKux50iqLrEwhU9fuO+xlj2tKa/
3pV4FwVN8BdF2NJENpUoy9fkGXMhkiJZzOZMuAStGtbN6tuHlC0wn8Pn7JILGxOz
znanYkm9NXeyOPKWvM9F2YE953cePFvwC27vt6VoAvtbTbH+bZ08Zwg/2xfHwz6N
nCzhHjR2pVwOIp4iTKTC4tgVJW8HU2s+yG/SP6hww/qYnwhArj40yL3Y21HyWKHE
sYhkICT2VNpwC81G18+V1WTxBcnNuQmBapgTHEECMF+bJ7lH14YHTEWCY/g+L6kU
fcX4HoiM8REYMg3DF63Ev6p9QbyrOfFN1eoDT2ElSpI6duekYhl352YPtEkM1qc2
3zlyIQkh9LbHbSxvudAhhILcp8+6W8iPFyr0WHT5rJP7O7YdXIHdRzpIgC9BlDCG
/L8azGZ9yZCgabEOdSWjBdzKqMwAAgZLODmEIKzZwNmoKtCi5sYsUDpWt7iI9QBV
0D55xA9WnJWwJiEKKKHK/lcvU1YG+6+bIVpfHdImUvkQSQHuG5ugiKSKpjhX06if
GumEAT3RDC3IPMDZovW5dSYUkrwjjDPRRuEX7sl4Pj+z8mLCx7SfavErqotlZL+U
IuoYPDdF08CWhYNeVSWK4eHvzsQcsekrJOKdE50nU4ANcEvuv0LA1LAY7NDWpftw
bCqq457kZQ+sCUGQrnncG/8nmgZqWEkxISHAxJm47NX+GmhovQGH1J3O/QdOw+At
Ai8XQdcAiUBlctDKVA2lZ6OQzO2nw1fdrNOtgJuOpHqsvZGbNs/46juGwC2K6qcT
FFbtXCP4CIw+Wu3fAQROxvyIYXvftVsDDpC1PLKC44F8kFwk0UqZXWwQpA+DjTlC
EhaI06SpeHUB1vvKzImqDQotLbaC2qbhkzH9m0yf5eti071uHlwLqaQfhC2iM4mi
hvgMAdj3UsbnZpblh8GZBL3BW8hKYnSNsLrOAeoK57j2zgZ/6M37DQ+G3U5Lyc1y
yoK3GWmKTV9k+iGox9lKlh/OXMuhPrcf0la4ZzjDUIP8ILGMl4fz4O3ZkXgFoEB2
WUueV2b19Mi84ZrMDyPP/QHKZyOyfQoXDT1fSNKYSxrLQjegUhVjFwt/euweIoO/
sQ+nDS3h4LnRUK5wss4L9+koL5DBPmb5CZSCMQkJO/2Sj+J+GRpdT17IyK1p6JMS
ueId+3zSy58P8FkpwipAtFcVlx6YvKOsp/DPZP2ReYQPzWW/YlSX/zc18AqtH5an
6/OjuB4jh2dwWww6iFa+EQu6encIyzOCkQinKzIRnSNRj0yKnmKHRBuNHn1J6ZKw
wvm7E+HtDYhYsHA96eNfxByz4yqtcbNTJpxdZEDDvCUYZ2VVWudOerD8vsJhesh/
LCdY6DbOiB3W1eXqb8ihbZ6eTIv+4gw6o5Z6/+QF1zBwqDbrxl4G4Du8mv2LPx6F
paGDbGsRn9scELbuJulvyckcxfeCee5mxOUh3a/JZdlKrr6AzUb0jSiKnYb7v1TB
PKsto7RylvpQiBUXAmOnTPcc98yNXAfM1QYmS2MUFsm+XKzvu+XMASPwPu7bzx3s
3ItLrRzFTvo8kWiCmFh/vO3pAIbLkF3CSrSP+hg6bnQS5yUNRisdDqXFN7DoVqbZ
Op19RP7XOEApdws93sthqq9uHsT1cICIuTrILwr8kIgkjTKFFZrdCG505MVvYMZT
rbvewFpCHtAfvHZufp3rKZQtaHxvoi4gxMy6zrEzIjMWfJDVLfHostIn6ZJo89KY
nkXQbZFuiIujYUp2X3M5qd5DSGbqRyPpJDK4Vg8AaSqDQBj99EF/KU27WurfaYKr
0fNcsEfZloPINFlOuwnzz62vdNKC0OTHOX097uPeXZhbj912lC777DHWk6SHCtK5
8msf3oV/ZjFkaU9ufmDT3M0LaZS/QcSgA9zlXGXDAimuYphK8Ci7RcNXBKvhLBt5
+GN7+hs492ATFY9IW+eKhHie/CO7WNnFy/Ul1+AzPgLa3raPlG9QhcHjy4VkXtvg
FwTZQDRqAWcdMStDNx/IU3e2+/kn817ormiBBJJa7rwFa8EZUHESOTho2PzkzGa2
sBucu30evsl3XNJnXb99XKImCkPJPy3aaXPWE2DYbmPGW4XQC+omMxG3Vs+kIsvN
gGqa/hC4jKmcE9elJP/o1xNSnZ6hpaM/fmwY4xcBIvPcGs4bnmBalQlWQ3Yz5fWv
CBC3eegi17mkEkuXXCv8EfKgaRGYSAtbJN5Jithc7WE2z+vt4t4Fa0v+TdOikWye
GIIUfNwbnrNvqFpa02oFS1IsdR51lc1GkTUup50pvegR29ohbvoNXhRttUHJ3Nvc
FKPynytkvw7ROoHxODQHpZWBKZtk2ibDNWv7as2GlebW+pT8YT4pRTLn/ecCo9LV
j5EftsQ5O7x3FRB7KjdJy7DjIvnMu3N8pwymlJkYnrack77j98wnD9/c4tOQOafW
sISIdr4RT4dMeC4WVpkBk/u3iONVbCHkLh0buc4uC1Jw5bzkBLtqhnruVNZlMWOL
w3PMC5RD/02IqzppU1kOmu4r0RwVv4rI3jSjJICWvji/brISEhg3S7V2goLZU5BB
29DmlPcX3kDWCkRUn2d/E/2Klqw95sqKg97ahK08b4byv9iNzBJ6/JoYcIhBYIYW
LYSRJFYZHszNB5Jr6k7Pv9ilAGW/yrSFDo9AcSNzXE/p9iraNrqIVOC+nBdHcZSF
N6aC5ga/kKmu0v7Cl0K6RCtN1kHQvGZKaEmAz+gAcpay/NJ0jHJR51q/u1/i6Z/J
9oT6MOa+/nWgaJpYhScCPBOQ19ebO3wudNeufPZNqhXw/9zTEQNf/le/E2oN6Wnz
JqmIK1uIOKhWYJwqqiQeFG7S2MQPP7m1Cn1ccVVxfpee0vINRbe2UchlILDbMuCR
3G2sUYdOx7x7BGO2uTEfyOgknRqIhPUhAJ0rCwuO6vqfuQLqft0jS14fqseW4xmz
reYXFOIIt3jTB0CP5Ac1IvMsVl6k+NCQ8gz7QaeclGHUVhhFPqv36Z0DkaxK81b4
2Ga+doOdFA09dcOil8zPRzk8OlcVyNyn6exZwBfr4Z3xJLYxgLyiqFGIwyMtGCYt
bHeZVdUc4McRsCTsUi5og1H5eA6K69LIiqZX/zuzhtwkgTa3U+8hTdyL4clGhVj5
DpHfzEY3PxKh6bPcujOz1EpEE4ifOj6gp+oIL2jsMvH6vyy2UomB7ztgkaPVRmio
gaLXdm4oGqTNUwdHXHqW4Q+t4N4liJy09GZMcr8/NaOlM9AicZKbMmJOOtXTMElb
1RQkoN8A508koT73/hRU4kad4jo4J+mUiFLk+yEzRWqwVqQJ+GAjNwUdFtKv1kRp
gjLwBCy75BlGFmyPsIsDl5Znmw6FSYBFAPT9Y1SlHEA22+dnr3dd+iWy7apMR8uS
IscX7Ock+qIt+84SortHVw5ZDIjhiZdDWWWZXe0NzIgwFCHnkbXdam/E9hz0ZXGF
sjQCR0pD64eKrleKVzlspfVShhrs73qk3lN37g7FbtYFDOUHXE6O9Wy1cCZbn7c0
I0XVZ5g2qj7Sg7eeLjB+n0WvMy7oTXiAEuQcPsJ50V0d5C9VaCwid5pwu1WCLR/s
Sae+xQiB4LtEWzZL4OLsmjPa+Gq3tdasuhQRvh/674RKTJAaOibuiRUboTA3gKfE
/5j+ECLnJz29LbgEm4u09bajdEzm0khSfbyG9MP3+uhcYzwP6ficwS84OR9SU6Em
rJXN6CoChuZDyQmmd3toS7JgIXJpUWYO14me2ZqIuf0lOGjaXyMHk03hxOHKLCvi
2OP33kpzpQ7Trozq8UdAlVOr22HhGGjSvOFZ1EK54H4EvKAFgVAh28gTZ5/UVN5B
Jzt0R3qj7/+NVOziW5XBKAqSeNF7jGBmaWbud+6aN6HpRwYkrs09eypWVFLNpXKQ
EaJ6YCymj0Za0PXocxssCoalSMeiSiuvnb/yIiFlnGu2gTSlLYsiMAH38MkjqsT3
1C+UFLcWSP+KFLzjP5vAUgsxUqHYK6OI4w/UBRKUajDxT9vEkH1xYalS2qOJofZl
/79zOsHHX/J+o3lTd3hyS2mSJ1JnytHuqvjyXog8OC6CDfFHomSw9VJNIZx/sl92
nZCkGQS55VgUM04T0eeqvKO8L8W1poetqo8sXmNnmxYr4wNYeYePDm4ZvX1repQQ
aobac1kLwtXcpeaz5qNTgggD3r/2hEoaecCKKICyg0cIMZwa4d1qg8gwSf67c9kj
NLiTV7fHNM2BW/jgDfJGHcqv0cboI7aA9TOpviDgzBfjRxjlmo1QTCj3bDi8XASh
POLHjkBIBEZNdAapxen1n7ZxMI4Qjg9g6clF9fRJQLUxTqtuu0/DGTa0uvI9yTU8
uuL5paaXcUeyHdm4tdJCpk3ZTAyjyvWZV1MSeSPdGEqAqcA7UYCr81BXsK43YtAh
sSq7JFaa39guIpJaI6FZLhmLQV96fTu4GVXHlLWvgNy/ZY01xFtf/JtGCwJ4+suo
IuCvFOdEfROE6+XU+hb/RlYgtOkDuurHIYeEVRKrkvZoSPYp1WdLYcCjOBI2PFV1
eWb8YPICwk4wdKNTfOZWN+n9LxvV7uAHmBUZl6PjQsNEHdLEbJXVX/I+r4cUHoo5
87y+fdJBhSf4BOYy9N2uFDiP26xrVKYMKCtoJKv8FfX2V+m5l8pO82ouBpidjuWP
F3wXcFuWlJak3EZ8uto+aTdB3qK65iEDTSsYmZ0EbIXaNS8B2z2ucV25FZprsWqf
R/cpGK3Qj9C4T4HzO9jP3InHZGbg4RwcQiGDQDsauifiTmjB+o1JqwHTIuJ2MiRG
FVQA+veT1EGJuYEGN5uGAtQhlszDUtxEhhSAcRj18Ox7zHzgravJibMuVlzeSBoX
1eVzKjipLo9tm5GjsowwjlJA/nciSUT5kjd490CN3ujaIkACXbxI+0ecW+i3EWtg
AUDKXjgFsMeDXnUgj4krzZp6JO9mukF+5c7X66AwrMqsRwLB0fBQmAdu/5Oa8MaA
rME3DEyXxgmV2xhV/ruSUiIpCXE6qCR9VYmJrHZOdTM1lm6s+HOLsN3wt+b41TYd
VNIqdvAxSAJUmp7LhcU7iw+Q8DuIkRZzCYydSqD2MFwh9vV3g5rd0NEh1OSwmvKM
keTzBiOC1cm+WfZmi+T+mCbalLWW8bwxOiVqij3+mKq9Lq5ntqNneub2jQcRxh/l
pAFO4Ez+kHqG3CkeheUI119N2sVzH8bRGcdQhXv49qeGufUVNi0PUn9vQS9rblu0
M/FWSMxNB+2r2bm8agkQQTwom8pBkB0D/9ddalumrlhvjsReeEIIQJQQB1mLpKvE
/T8QiJ+wQ4R6ndUjoPS7h/QsgpXBDddJdc5WsNJ7UcHg5QPFkbhfc3w8q/RRT5GP
fnLpz6gLp92a4cHHfc9Etza0H94ARncLWTgJyWOXkw+J/Z/yJHLyEPvJ4epHXE4+
5QUvcYI4qixCo/yaskIhJdwKVTMqAZWM9kNNhppUBYUCN/CqjadPM4J3HLnN5jdf
8JDCICSD/VW9NHwDd64Fxcfe530tJBnkd44L4C5OU0CVAJficivF1RtLsuoMLN65
2b+R2xNz1Z0r25OiOJW8Y0DLRdder2cNvZRWcCzVPFzW6KYd4miIYHgq5A3KI9Ff
D+CHvYMURBNB+KZ7NO8YrQKatS7meH3WY5K1gVJZxmV2WebB0ag/gb4WA0AYxKYv
VDMO6dCaF8tfvrrjNE+7WlSKzguH3v/TMAEEbiIfKgBOUApJ5SfFjZs+SQoc+ilL
eRTwv9nA7mXHD/Gses1/pO1628bTjmbHn+/I4ZIw+7jQXd+F/PRvRF21Hm2Oyfq8
grAfZWOxipfg7phh37spqrJXfZuFzs/SgtEeorI/pKFrZ9UhFe6r4v1o6MayAzgo
QoEtk6CVQfkCyaY6J9kx7rI2CvWLXRQ612YVWNDdyXXBrizypmXnV+fcpGrvPKQH
9j21KMVK7B/qK/n2vaK0pcMZlBEQAMIoLQJO0bbyZeeHCUh0bE8HpXvIsVJxwQkk
oH5uKwBn3zymuw9W7fvWcCgANYhJAU3/bBtepfqO2Y4pYrDyK8qAbQib7pvBnbfD
5Pd/QFF4c743VNV/c9ynM/nPpnAvIDGC6q+3KSIiAIq1V8Dg0AnojqpiPoeEaMj3
I4MjZ3dtR5iwWtdJHeLWSIaevVO3c19BZw58hnVdINIja6d1DmE1V4PYSI2JhiiK
QVw04kVO0D5aJ0n1/SBYhTUnnDSxMSaGCzESlETXXioSNYBzMQmB6JdHzP2OGAV9
D0BDmlMs3C1pEfmmCcRjlzgO/G+GFFD6sEjz768WHLVmIu6PdY7LqHwSrOdLGAjb
L7yR9qQ9TaccICeND480T1FhqSr9e+KE33Gupx0DbrRT1a19tbsnQoPFeyqfAXbd
V0hIxiaw1KvybUZ5MMLkNGKuk4GQhdQnAClvSonIYQC9mqSUDNtQMAgxxMRFi30Z
mH3/RoJHcxJtaw/Kqaaah/6nqkqFIJDPogsUGi0StBCogiBvRbspEcgauqgLqaF0
FHKsn1wwsq4LRA8li7L7rIF1Tg9xPSgIOcAcxIoTryqo3ZZM00kwZDElKNCM2b09
M0/v2frB//viXpSRIOQ8NMoxXLXUS20yru9xA3vZN2HYmaYTMOIWhqZs0wgT9XG0
93MMqNETXLOzG7juHXY0KsCtxz0z5whbqpUdYnkfRW/o9GEke+jp4WpIrRkS6YNy
rvZTdXPZQx62GnuC6dqddMN5bZskuFWKXfVmROgoqY2UfGbfIRXWEZCb9Tlh7USX
DW914NLi928My8TY6xpHoCLFn0hA9xsazUrrxrDabvwwZap6ZjTRnuKbMWWIvqkf
EzL8GJHPzDywj0aBfRyqiyUH//R7nhY7LdOy3FWZqQlvw6vl7fJ3bikXTc2St2rW
qxWC489her5yTJQUYeNys/r/qciQuhpBQJ6slHCvUZ213psgCeqIoISjE+bmmcgX
rSvTLDC4k34V+pquzyJ+vdOgAwqFD6kVi5AZzGV+aNt8nBhAH7d3sVB/+doGTZpl
AGo7Hxhrb0hInRFQBAMwj/hRr4qGz7pMe/o78jK1woppfeReehYER4BhM0dAz0s5
FgGj5k8pwPPNbD9i/qiS8JjmTO8kelQu9V1TB/DVgs2vbD/w0ntTDWd7/Hk51r98
+lfsp93n0Q3fgehHEZdZkLm7p1nSQaIXQ4tdbGRAb4pQBqkPnIUlwCYEF6EhO/hT
8oQGnxaHABj0vZmtw8kwb8fSMJxJWtqDyaXr4gp8j1WyVhr9bsnloJFmOm5zyQgd
Fw5KxWxeCZckLJt+MoBzH6dS+JRGBMj4NqUknoqClPUFQ8yi4s4NEcMD25ZYeIQC
OHBHq+MgOkMPz0FMDalx2pcgYB1Yoq01aSD3zZinNgOjAdyWFhDvOFmAQUqXwO0J
j0EXkWWYm2paWlm1s+2uWY99lmq2aI8Ls+lu/VGdPRGP4PxwCJwESFseLGnOIb+N
zr9fk8WQZo0uaRCve+Sy8Mza721EGLBmPCqXo3FCnICPNfbsqnNW7u13dVS0XZRo
THo5uPsaGMiZmeL9ed0nDj8LxQPzRh6r+AfJ33ZvWDZeabp0Ssz+w34mrqgQr1wP
oTLvigqpGFWqUQR7Z72MTQ==
`protect END_PROTECTED
