`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLcPNcEgLEIn0UKDDHqvPt1d5ycOrlm5qA0tkDVwGWR3
zsfKvZ7EaJzO8UoP3W/Jkb7AelaxklFkW+Nbi/0RBGKjTiqfu4iW2gUOyhVJFn9b
CZ9grT48kQpKKuTkwkgWBlZFnCR8vfg4mPyDs0WpQXy5ofh1AjCwO3ulkmuOFV3G
SQXOtWcCweWJsHkWjdgjHL4rzwoYGSTMB6GER2tq5Dos/+/zEoFA73ZXaVBWx24d
/lkwFiQe32Zwr5HEyIHfA5qNirA3GZ12y/afCiJPZUCAW7uiQcQ//beObt/6S07N
/SRag2hdZIW5gdWnIeqqxzT1ELpZHiCQCvvpjBUcC05JHXh7HAHXQ2kzVnASdg2l
PHXEUagIhEhGZHytDVhSDh6kCWIv8gsHwF5PiboOtMs0Xt4XE1jhl79MtyyG/CVQ
1+ETqPVlfR7KF0fMU9kU/eeQ1LvzS0oWglXU0EqhXNqKfEAwdvTsAEZmQIx9wlW1
T9VnYq72eQnN8HXsaXCPJlIED/zjBNGlJnRXA25Q0b6xixi3l1e8MaB6RF88RL3D
ERqC58w+B71+CY6xyIFjH2ymvhlvA9wO94XgrUzJW9J5w91HJhT11Y+RVqBn6/H5
Rs622JPsrs4oOONwFxusPxabitbRGpUudIFm8BBeLX/r7kTlJVUPac5HJohSNPuz
`protect END_PROTECTED
