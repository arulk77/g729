`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNxewl/XTver4X8MbtVVswQ/KW5Hr9aa0mWU+qvAycnaH
n7sbsdgoWhGRnzVyKL5xLVM/BCLSzstldbopEGUBNAkwmdncMd25drdAognbaw4W
wgw6K1upapnsZxgZwIQ57fhSSJ0xnTPHhf3pvEaLvK6KgvDBO8Lkf4upPft2sQpq
/7jxQzXyl/FmJ3XCNVWtrKVzXU9NSPTr/LOW2ijyjoJrJ79HwBgC+0LTNPsPIgnU
`protect END_PROTECTED
