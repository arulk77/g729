`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48gHVyKCRSSSmOQjNPBwYkspcer6wrOjybU4GMYp0wmj
rM6/Luxt4f3v+iFycIpVrcPBSLVQmNFHLQg3niEmveqfEjg2wkbqk0gfyGJSyC9y
M76N9SpPLFmm+JbzrpIaU5PX5IWSUcI88vCY/13H265ZGbjr7119eHzEbD2BP9z6
wDfr+zpSIw3fkauGTEqOjI87cYUvlg3IwR2L24FwZvQ=
`protect END_PROTECTED
