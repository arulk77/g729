`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKRVxXNgpb+DiI4ihYhJL1EMeAlTPg80vbsm5ARyyQwa
UmlBTAqKMzshUK6BP+ofGFyxrKqq9Iv6lbdG8Pjp2a5oFDibCXV1mbVFrpTXWoFt
66/ZX9hoGrWG2SapEoRwhtQAe1xJpiHGjZVWyjEVn/7wWQThCsxhoj0EUlzdEJTu
N39/bYeTSP51fR9uqJ63CxwNY6OFdU9N98HDcjXVqt1EFwwOhErKCfrwnSKH6OuM
I6AMACcOE5Hk6e2+RkddHw==
`protect END_PROTECTED
