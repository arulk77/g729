`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJdmUjoPZ8MY4hZhLHEVVw0LhLNIIWvoUiMzY24KkLmf
PJAiqJCT2CSmoaVwjXuTVBCds8VYjeGgVlWtrUgKoylyWxvqNZ2jv8irD7ANDSQ9
oKfrwX6lCgSB8dctyiDwKvEpe+v35/6hCVKodIGtLKsqgJNCwR76XzB/fTgkX7lN
0q1WuLx48P9hT+BNJWEHl5YfE1BxGarjT1v8fh/bMQR0NcITkivwhtjaE6H9A5qI
N2gbRqM7clM/xYxxT9v+OhEc37xDVA3L509QoqSak4A9mxJ4K//U6imt1ZLrIreY
T4oz1BIvD1iD+4SyF/RR5c+eXzXp90lWng/OaS5BMUzwY4NRxZgbFvMiWMf4u8pW
tP7xkWS1OtEEJIYCGdUZf64wKNdI1jiUEw6mhT8SY+9bdzKSwkH07TUy3RPRY1sv
`protect END_PROTECTED
