`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QNw40IqJrFvY2E8HYWz+j+ejpl5znwHQiATOEHBgKp7Vq0ylx83xng8zt0NWLt4p
h7fbuVne8aL2yQha26uEvwr+lt979JUTqIZOdKkjVV3ycJuLVFu1gQSVi2RbHQLh
xYdy+hzqbsQVJvD6hcRlZ6QMdiTKtG40ZavrQr/Pe2I6HVJCHY2g6+ZhZv2g4qLi
`protect END_PROTECTED
