`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
y0FlEGa0GaPgVOqOrTGoL1ZjTRqSTY998TLAHnvQ61tsIHkOnwvcGPDlRJPh3qgL
CLPzeM0kD2eHRO/yOMtzgt95FlqmxKFTW9iWiTvoYCRospab2tvydT/JVzvqSyxR
ZokkhxZKvPdUdqPDb/3TQirypxFluEWaKbhkbitrNqiWiyhwT1jEt5JbnrJKJIqv
kUxW/T1LewM2JK2/saL00OCfn/U/Uiy3bxx0hz0qIseuHrmAUyzn3g3pgITQN1/O
j8pbTtkVQkqEiRxnBXPk7HqGc3NniP6AbV+oKaSxYoxvTU676w+AOTGH16kV/QwR
zqGNpmTKRkirWRT/1e5jHADgtpGuJytZuAAGbPOKE7+mknA/CkZtGh6ee9lAl7OC
m2bVSGZhZPKX4BzSOhOdpHCLcl+QPgD/e6Cp+yRPjlPW5oj68+qoyGIGA96s97th
xg4LXsdDO7qdR2M6ozX74w==
`protect END_PROTECTED
