`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJWyWpYkMrgQLhf4ukkHYB/P6WrfSBS8Tx+iz/cbigX6
9VKOYZxq2/kZeLlqHSeZ2t1kiy28modr1YTASlXoymDUIDOY5D+TWlytUf/V0AX4
sDfRWI581Vi7HFxGJ4+fpYtP8/B0xBrndYRL8XA4Acm5JJ7kfs7gYWduEarcrQqa
AOMEAiC/lhgN/JGd4qNYRg==
`protect END_PROTECTED
