`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKtoLeOO29ewr+WNTG4AIbPuuAyDpNaz3jZxgnu8eo8d
OVljJSkTsslvWTELcttKSEP9Ib2uaUeTY94O7rE74E6BL7blXOYU9mB4adUWh9/L
iP1ENpcq/7c2cAsNiUj49SiFX4idcQcxFjmdKG9TNJ8Fdwk/AfnSl/VzjJSvnlOn
mHbuhXf6dqnk1DJdoKJXfjJf1d3tfZKo0cHEZ7aG0SXICRoKvStTNwyxE0g3rrZH
s83KXcwFof7DeDt/5FevDWwdXW4z1nuLNS2oc3ByeLjkCclRxxIJc7Sf8ZIwwswR
itjzTnUHUrITPO+Kq4SdY2hqLXdzy5kmZVAj070JqvLJBkiYKpGmjJrA0gWWOmbv
1DW5DElSsXKA44X2snk7fKx7AgRE5NOuXirl8I27Eg4He4lWlNy6zc5r2S/pfzaW
ql4mEOkSf2tUlV5rXGJajrQD3ax4fOp+RIqs5+GlN+Opcfp3djGbsQF4CVhsPeZA
ntE1t5hSO460H4lQkT5mDezagficupy42Adq5bD0iFI8OZFRcqMtaievyfowpqdd
IgIV9fPF9QfTdwj9Aym1IA==
`protect END_PROTECTED
