`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMdZ2flhiMj8wF+3uJw2EnQjymntV1EtkAcE6OJAgdW0
GRyqS3ui8XCVtngUWr4TDNA4lN+P+nrZ96rzyhRKT1odSaIrPdKERpKiguwquCtz
yNOiuBXu/9mBPtP0O3N+9apDp9CATdsOLeUjnN/v4/V+mUBWotSKVLFYcU/cVlLz
w4chz7lkpgHkPbH0cCVLdcnun/3sT6t0/0UcPN4p39PzqyCXiH99c4jOOBaWr4Wk
`protect END_PROTECTED
