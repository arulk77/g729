`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zjZQp42f/niJhsPNcyVq9oOdBR8fl/rqHZiGkVA2GXW
D2d03nOBr5bxksqI5WBVkJHJkdmiT8Tjqats7ZhykA24ZgTarc9oo0Paek/ie7mf
HceqgTT5cTu5HBZbp4SQBzlQqwjVu8VbHWXiJEx5BP2HTJTL6P8Shdj9rwo6U3M6
oFdKN8OcyHsROvLKjTTF4tCuCaC46Ym6Ow7mzEa0MEfLz1XzkldL87aVraYchQAt
z0vDDY4U4LWySjR1s5z6GMCr8gpc7b4U1IJZE44E8a4=
`protect END_PROTECTED
