`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4z6k26ge/xjjIAjMw5cKXmy6REOpv/W6PbQf/Knhw79Q
cOfa9crhcZ87zOFiisJ1yxAt3pBHK0s/ABtD+8DcYnpS+uKmLJ3JucXQ5RfUpcmE
zpb+yq4fKkYgrYqZPL7iu+LJMJff7GjmxL93SnedSvHdCtFRAqT6p5IywJ+B79mY
ixGZDv2aaPfocq+b77JY+1X5RQBgJdbwJj1DYEtND0w=
`protect END_PROTECTED
