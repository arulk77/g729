`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45phzti7pWlPp/vvKcrG+6+Lx7gm8cOMHwd+fpVZBSdc
BwndrsYOM1VABCgkoK6MhTrArerPXLssZWPm6u07g94OpzZYcoPcYKgW1rPKpm4m
BXR8qYfdKBSf2QqOnHbPdnN+QQSP4tdKb7ohapN32GLxOG7dt8T/kkk/PCH0U0Iz
Sn4vkysIXQN/M1TpIP/6xI3JVfrbcB3Yr07LFmxBaeRt5WEO12YjKtYydblImkz3
vMXpaphc+fmm4JNldcYn2Yey0h7ubnvHcY5SglO5nvsMb1rrp2eyS1UOh8Yr4PXo
u0vTa+8nRIl92hzQT0VEFBqtKUytkLSYBHdaUGV7MUjbFr26/ZCHHwW8085cLD5H
Qzmrc+rfV/R+iskj3gTtshnF7QRJMcODFCowfFcAJE1qD7gl6+fTL09y2DKZrBjT
QSS2PuZGafqCOQLHRz0RQM+nYsKFpsmid9q5NKcKVvdHXrUT+IVjfXT0etU5hyLt
DJRXT45RBgmrtnMWqdGNZ+Ci4nlFCDful7sD+4kGZbyOFPgOEHh9kcBWiQ/9rhhl
tkQ8mKRebxX4/1MT1XlHY0UxztwRHRU6rcYBo/TrdKGWe2GAt9b9g0F7rQWdT7o1
YF7pLBdvAo0bFOEO1IExd/4Cdax+MqVJLiTRKW6+Fq/2GZ8JnhZribIT19TZyQOn
lOZ2PIIIfYCb8QJ5OptWP9Yu+JXYVoBMAyfUBt0whhKvofYUsRIAU5+KDUjA6MrH
4n/9nXptjxP5ccExygIOJHeDwDPRUvOPcVk4jwaW3SNH9Edxan0MOfj8BSgvIYsd
wxwk2W8U3yYY3tYBbDXukM5RDPiiP7L2dF+2LdBNnrn3uxIWSlo3+7zbfCPw6LtW
H4egF0a4CJ+HZod2bUa1ThxYzSxy+3mjhrNYaYn1y9QLlg0DE/vFb2rtJiQjccwt
ooHa8DQ1g9FBPw+j1jfBCqStOeDAgiRgilDueEu8R18YT9KAeVa4Iiaq8rTwVJgl
0S17V5xrHAmojX62OjfPpiMH82ealZyyeTPcQjeuxGM00qamaZAk7QXpLXhfr9Mb
//yUeQMfJCylkBt6dp8yvHnkwyzZPyGPah7rt8CQcetG+mch2ihpnCQvZHr6ws/G
kik76cNd/FhQ3t8PM2Cgc0VzSLj1lg/VnkYqJzeZPvcPawOjSGHGcZNxIkvx8lXz
`protect END_PROTECTED
