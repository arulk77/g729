`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveE3AP2Dll/ujVXygHaxzmLuIil1K2lAtkzMcClmR3r4/
Xa8NOTuUS1ASaeF4p3NVR/vyBDtVtGpQhWo3vOqIRDo/TuKQSe58i4CiN0amfOJ8
kZavgD5tTCDFocqO19fQAMaXBsBeQgW4lUA2R6yKGrG7QBfOGZBltzBLoiW1iLcv
TgvzVZJxcs/tuc+/gbQn/g2danJ6PtffQZ/GdZa397jr6fOolABZ0ksRG3fPSUmb
8EbJllacxj2te9wEc4P0IUKA6PJfqPEge+IG1OXK06zxt5FhDREynUd1Rtrkir3/
Z0iRvwnpYaQKTviP1V8X2G4hyGA2eAX4Z3vwYepLXf71/etUdtG7mIQ3/TA7AwzK
`protect END_PROTECTED
