`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNJQNz4lkRiHJ20L67knFNStBzelyH2INcbawvxt0S5B
yBPsxJe0nlTK21b7o1qCZoNMOGx2Ke6W1Y2sTuFzE0lqpsp6QsRkhlNxDJxwyBRm
urI9PCPSIxFfV0jIYjhORxddxjZRT0VnMf+Czl1qG+/hpBIJ3XNEd5KIUZzrp0tJ
tj3xHKqR7x31ZiRc6vH+M/5pK8VAbsrz8EeHHF3Y54SUqQqifCzeF0RVWYE9eYRy
hBUHSugBva7KGnl2pyLdgQ==
`protect END_PROTECTED
