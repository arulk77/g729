`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xtFI5G9gWLL6mElMo5br+fsGkVrzNN2p6tt+5pp72/h
i8hHv98/I1L9m1va1Me9MwH8qFKw+E0fb7CnhtV2MSg3cTQ1ui6Gf8i38iNpEgv/
okD1TpYI3ucrAgiNbCa5GP8Vj/s5VCtcgbRk9Rxaweff+4a8DfJf+zAaxwzC+0Ni
9ezlqdobMZvUe015Nr3rsd6zfksQO9lYZMfUjs8liRi7/vYSsblt147j8kED1ZOp
1//7Crr23n4gYKhVzyv1oCggZdGrBl9jAVGncH4mihsIJMW/K4YEoXGvI0AfIAOv
voj8w9vMm75EDHAK70Fe7o953f7+i5aXhorLL0+9IgmEn/pZcrNgqX/3caIE8p6N
GwylFaP3UIs1I+3tAOYwDQ==
`protect END_PROTECTED
