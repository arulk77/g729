`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLnQjQjb2jPaki742RX8mpveSEXs/9gVKzx+zAfYB1oC
WQxZph9xVy7LBdS1oim4WuahIZyyFL1Lh5hYMAGRhmmeFV31SxWi6XHThHMnFxNI
FxnoHvmL9MbcJRhCSdJLluiGbiGK1PlNiBgZ7NbEdDpp65SBybTCuEOct1tnkRDQ
cic2uj2vav5qakte0uo/BgFZ61cZlvTaut6uF+pv7QkF6AKr3T5gV4r39aJ8PJK1
PvGyHfvDBeITh7tsqjZSPOVzzQ0TMhILDiabnHnUwXDnhpz86jf1Mj41qEB/otbI
xX3cRVU1PQwXKB4ncOX76g8ClRu9uQPbd/miBXP8I8i3wqxWBkBMjmilKLktR+Dl
idjfiQCiNPS1EkfwOGc6+aW2xW96ba4wzbrqIYh1X6a5kjBj3yWwym0UI55vEXzA
Eh3jmvdEwMimTYl+obwsabtVG37suxR8WoDiPRmVh2wkfQJbyR65sbTK6y7dlmiz
J+0it+iYfUMLemlqBrbas+PkoLW9q1FGfycIj7amwE6a8zkxL03ScHtcEyKaJMDj
ipcuGDBsf+7e49pTA4iRBA==
`protect END_PROTECTED
