`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44inMVFpgpER+rSVHIIB8fk2xIq2qfeVm/8zp+HTT75G
lzXSpiSZ29wHP0h8fsUf+e2248GDZ4KM/Nk6/OtGi2doa36NLL4ARoDwhPNkiR08
6kchnFgO4MtHZBhCaYfAAGpxJgqE37Vw1W+xX2Jd6MtYXOK3C2bcQWiyxZzS2TQ5
0DxQHWnXg01dpN9uBUKxfBna24IKce30cewbfNi1I+k0BsBbmjq9KFDm4s09+R8m
Y3VJsU0tSMTbndLoZtRAtbdD9pU4CN4PVfN87nM2TWNstSCsGQ60cqY64iQt1yWT
HPT+CPwhVoHirJvfk4uaHVZd1RRNoNeiaflhuVLUPwJaTNtpaCMKMNGKp+USnRKA
WOi2A9qTaEjubLkOCwQB1Q==
`protect END_PROTECTED
