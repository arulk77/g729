`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJnXml1mOGp9Hkj910GkN7XK3uBPK0cVDe+gzwhYTzWM
C1YzNy5EyEN2j7TxdtJpmvHEuG3Z5w+kHYlxRfxEmj/ZmX2XkGmRBqXukxM0CiwI
Y1jPJd2b8HZsBEfg892/0pdR5baVuTXfPWmNj5FEq4F561bRcKTKTlWqRNixMS+f
9i0tI1xvYBOwFqVEfmISLK7WWxQEAejwahKHWUNxPuP88otiwe8f7sCXe0BBWQUM
zhopY3Q1jODaPwaHGz4CnHPPAA3LNQv/fwVqS6q1qgkVTfc81I9HP2Fc7rbZ1vc2
4heaqDJkYE85ardZdCS3QwXfI41m4Uq7Y5CkiNwe5zy1B4zKLNCdF2wz/cFdGBDV
Prr5oTuCXU4sb+5//x0q1vSeqD3s6GlFFhmehSsQpWkAxGu5UZ10riQftBGpdtHx
tpOsjrBbDH8tb/IREI34FgNRv2jwKuKekI03Jw4vKczGaseznZSXXi39P0SlT8vo
tC0dbizwClxHMAQezYnbA1TV0M8FnMu1Z5rr9nQ+/0cOYv/f7sPlCSOR9d+ql8cs
X87/NCjVh9QEtqWrztdkN9Qh5PAtyXBH1yIqG1lypUN0blwO5iFMy6LzortPYAj5
DC6rpliYtFikTy5l1SdV/HCMjdm6Mp/7keMFhEi/Fxjk8S2Ta8sKtXG/AeiFGQNA
kDxfOmsv/f44NR7kRsMBsCom5A25uE0kQn3sNwpiwzas82cuGzg9DMfmW6did+cH
MmBBU7MSsB+iRwQTouDcP3/IzhndNFi0O4NPTqRySaFoMrLlKX9N3ogIOzleNlAw
HKg98kLxKsdYeZ8SADYIruEOklcbQqCnFFEQAWJIa14=
`protect END_PROTECTED
