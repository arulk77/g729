`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDfMMl3D8Rd10tzypY7xO+EvTdwO6A+Up4IJC58ay4nf
NwzvnGSPefE23yRX6jajs/kEfkFqXKLckbJMz+jPEna8DBbkSy1j9AAYsOCwF+Jv
bTN5g1KFwU/HoaXvdwiz601pSDA97oa8JNepb8Gc+K4tqr9yxjmkOW3zO3uXQz0U
uDH6OogIXDvNpI8u+2iQ+tfLjShU6fD7zoHVBIcrmgxL/97u/VNNbVem4ya/tbF+
wrr/Fr1S173LqR+hEujHc2wPdpS+2idZHkR+k16HyJxTbcC0t8/7/XS6BcxHgAHs
1NzadcqGNcqKnkVemHN5XvlI+QEgsTUe4TjIQ5lDxnm7gvbDncWYeEsw3zUaB3Yt
sDqUwAzWR90/tB5wKXNl8RT2vB5PNKP2JG9LYJ1D5X0BbpAlIeZctfWwf445N7OR
vE12AJMhM4sMB6uKAExycsD7ELRD5S3b9Gh+qyAUn/o18rq3ONBM8JAA6tpd1gyi
0Pke1uV22ZofgClva4miziW0CBLX3P8MEKT92U2yZJFk5ArSEBskfB3JB7U4oV7s
`protect END_PROTECTED
