`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHi/QEobuDjrzsiXDEM+MXyhFT6j9ajb8pV/SQrBDvcs
bIeWNbfua4JP/jN2AV9wRQZMR6ehHYnTEDQpWy5J4Y5CrDKk8E+w0T5NQ2+Tl21U
y6jkQVH5qBRlsvhbb/SYeMXg82Gh96bvzLI7kHhuoQPlcPnKoEx1dkgqgl6IXWI0
dBi/U3eFQGVkRKZI5N8ajGySWvFH2EPEiwAgFaQOezwzhQ/zD8OCqfLOX8a/RXfE
ROe3nsmr4jK8u/6rv87jOdCzxhdiLN7VdrpVofMc3Ebr/jxdTcLKZk6qwnMl5wgB
yAxoaFVcZxhxGRigzmD0w1MZWGrvHHSfTVsyXYmy1z864Y4z35rzXBQJQlKN1pF9
tcNYhVozpL+0jbb/MPflzpzft03YYj4kIeyx2ZYXARvgOo+82iAEWHT+FlhMHI0V
eUCkFHg6bFlUpMfNxOtHRy7zml/NuutdTbNfbmca3TNWmUvoE1e84OGIF6hvISGy
LZJJOr3h4GgIDxq2sWKYJ5fd5J+7R0NHPe2G4cweQ9PGp09PKth8QUslD3V/q0BF
dTCLwao09FIzknq7sAalDZY5JaevVaH02FdtLT1Sv379T5bUJ7enxktmJDpH2Evk
qfyH0/ezftXcmal6SHMJkWfq3BIjrig2XImi6PSQWlTkc6xke2u2Fy93XYR/Qmtz
`protect END_PROTECTED
