`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
l1hCsWRrO15B82/62mxt3/Ek6PfEu/4L8a3K1T+lTwta5VMqcKYGc43DD6FmpWkP
5sryKuMsADPzGUdonnj++HDCyRoO7fB/fw3BApFq82ip5iG3QKnzr9w17/eR3vCn
gKKWLUdBU0V7rd+Wthgg7kzIZl7HDzb43qxNdiLudR1YC1zAg0GmPyh/pDw/f9K2
DzlJdHzp2iCa7Q2SwmSJBYIDl6902u3lezL6zmqwuLi+t8OgUT8wmXVcLUx1GDFA
828NEZ/RQP8D8UAYZ8zHibJEaQXlkCbFmmL09qmkdr9hoQJAcldG8xqUUbYAvrhm
4ANeahxRNMBmbfyKiZ4NdN8VIHXcGarKGwbx+kXTNuc=
`protect END_PROTECTED
