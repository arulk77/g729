`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
0+OAdpuXHm3CIv5sgFc8o89UAEAq3JQj7RY2TBT/dSXi3Q5JqBbB2PYOwEQD783J
F3JeL2WirGo7SpSJ8O2sY0NPN1P3nyHrIfuFWVO9QyZMvRURYiVvEwumorVLnqqQ
rn5MXzL6v/zrlmtzLZWlRN9+zV3TCeOmY/cRhFHU5riXZW8Om1NWbeXY6PvPIOsH
excPStSaBZTt+uZ6j7ADjD697hHtNQy9pecTsOFsXQMqakT+fIiAzP0Elwo2MXGv
mFUeOwJzgzC87nvtNfHPMKU6yoX3WAItoeSwEq/4NFvvROviha4WVU4sbwqxsHyt
tOfa8ilNP89j3Q8D66UfZNlQDIxUk6LUTke6XLKBUGOByNTq8haN9AcUXPc6wKx+
rmuLWmG4BikZYqBQRunnmnTegwMGn3YS9uB/BumkpOsxCGUgoG5YjGthKqtDXF/V
PyVvAjLmRZ4YU9e1n0AtePyUGvrG9RJ4NyM32wim2HFawrSiueHdOMEWpm3wfNMg
sFsu0jTJYrL7Gs61tUA0UBEuFO7yl/x2BcaqibBzmKk9Nvv0SCy6eeR7nBvUq3m1
3jWHHBz5U4wk0fCqmYpECA==
`protect END_PROTECTED
