`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zRtNRdqj6zhoghNjrBVPfmzZuYvQET4SoDzzRTYSwhm
MsPJ7o4uR3WyhAeK2XsOIoKTBuTgIF8KWDCNDFkGNWsRSgrimWvtv26TNa7EcXZf
98aBGU+4fSNIe0Equep4Wv7WlcCJGPYAl0r0mH88uj2Wkov3pGGHMJfzLYvNd/JW
VMY+nYV0mORgE/yy4k46xRZT2eqjeVPtG4LJMBIy/8UIUkpcKP7wcqKFDYrxR2qe
UJL9q00bKQr+Pb00E0LsZxKs9GyviSYmqm7M2a5mDMCAbqKNDeVSxxsT21I/9Anj
Ne7gJ6pABC9MyLfy0v+DmEG8aFacOB4v/DNmOM2gap/EqpCfy/t4mjbFto1Plx9V
x7/ml6dDYsp5I694Q3YOILPWuPNOv9RwA3IK19Y8QfLMT7Nn/e1FW5o0LULIA3KE
9OFvAL41+7/Y+gtePTU86PXl6z6HGkZEvnOcZdebe5T4GNhYtMFwZbbkhSUn7OiT
`protect END_PROTECTED
