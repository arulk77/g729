`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOgXMcQZr3l4ZOb/64Twr9FPjXFbNNSQTddmDmDyJtcH
o45tDEh/02tQ2UfJIfe4Zuny5TRvmvS0U285ZVkrbG8mAlp705DQxARKbMslCDzd
ayAcoraOaghRMs59VgiAUZtGG5CZTIKU7cdNKOOsSyVB/RZoX/0wb+wzNu+hq44Q
Myjnb71wNfh+JkYtVl+nsCn8jfIjUJ0eVfrQpek39bOxK8VpK5YK103F/ConI2Wr
Q9m89RCoQGpTuXDeWFlfAS/k9Et+glv32N01UuXYELMez/rqp4LW4fr0h4RNyyJT
u+uGyISZgPA79ryNuS9cvKrCs4oNW2D1vwxpUgh0Wt0LiBqtgqOTGkuOZm7G1sqZ
J4R2m+6FVXZjdXEpgLCiU2lyD9168IWeN/WiVGk/0Ji4CTRDWQPVkUPXfo1cx/gL
z6SINoXUBiyzdnwVqtEdyO14ZC9sR/2B8GGeA4s7bbH0UDCJxdrFtDQ3sySPgImo
CdXuNatpX79qe7hnmJ9GZv2+Zwoq7YNiVP45TScMEGvf6/xM9M2a58USXTjJ6Hs0
`protect END_PROTECTED
