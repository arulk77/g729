`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aX2XbRraSBGIZRNcI5uftozYC6SImq+lQuqblWwBMhOJ
3LeLMHlrmSlQQMjgwfhqTdAwJ+sbOZ0RPFLlexjuz/BJZXRmV+mXCmGjzQI/1B13
RTC5PaE9dcMuNkpmpQ7l1UEQtnIdo8YiUCtjyqAEBa6poemSxB6Qb0gr/epE370E
kmCMDt+UmFv+lLBUaTr4V3dEdYe+9RBmzL7kb7sj9J+545iW9ar/CrYSG08kWLz+
Aj7ZWHfEVKaOM5q14/FyDkT39q06tIXeI2yEmLNfEb5oFlAQQaZEbTPHbrEsgeUo
z1JoCU+emn4I3KWMiRV7XWeACBSMJ1H1G+ribYryBVNuIPf24XeMbrrzpe1k+rpK
EWAIEbjhaCaFBe+1Z7L6ZohOC7DCrluub1swLsTIF6VqUd6WMERrtlQzePSZ9nQ9
Rx4YSSKZiguF+GWser3JvjLRAINVhFBSsC5uikv0VQiRxzsL7lgzTv8QV64O6D7b
z94fTVh9kwxsOLKF5wV/orYQ2dGgDYsMapFSCfVb3k+9kJyl5oHHZJqMDQyN+3du
Yc1bRzOCHrsrt3+VkYwdXhdMbulSmTSF6K9N3b7ytYPzOG6FM2H+l8pUgnLYp+00
ZsuwF25jgIqe5hkR1ryUHFE0QKB+7un1VciJXVINAmbi/8JmpyouZBmAf2gypqdT
VjiTg1ZXbaTsjBIHVad/lkuNCmjCYzZDTYGrgR+rmFoypb35sWVzLT7hfiBBYTGj
pzn73yPTX0MnxY4+zbT7/oo23nQ71SMqtS0aNsGsh8V6RARUr9LZ6Uzos/x5Jd7x
pIfK+HOuVx4JgHb3HY9ivcwgzvVWwZiNGex5CrrF71Ioi1QyBtrvvk8t0PImrT3b
X2H/rgZO7xTAg32aVsXQ+2eMiOZ61fouCT323MIyJzJEYBpsmTOBW8VeEtEDScWM
o1g+K4GiJXpRW8RTeFCorqsFu0CaS8VIUQHKhJaq4h8ILm3pbG4OOMOhkm5ovM+f
QLfFX86efiwC7dJyXE5VlqdpgpX/+Z+MS3FYDDIv+XZmQ0EVC5C5o4AgO9IQ6GhQ
yN9geq7/Fzf+JFlfp/zfgvr5f4eGW1FmD6+yKDsX+x3mjaddE5s4KMpB1ymFQKgt
Ziq0tOVo5w1Fc++rbHLY6YdfI6+Na7x5UToHvGoL467WK0Gai0HP5b8zc4+eO5Gi
gord+g1CjGDI6kmmgVeTlylCwaW6Qs/3uPEvme6bjjmECjtAfI6fTbrTeytLoLDz
O6yu3M1o7dWzNBxyuBN53/wJK6vfRGcPZotI5mQKiXp9WfPDvYJZWZHXz0JjMHcu
AN27AOd+5DelcKvDtE9iIH5DupHRq1KN85D5xOd+xPTDcIcW+Uc2dsRBqcmkur+J
WCUjC9NTvdMAP2YIyJ0MHs2/qyOP4S84393pzwSFvpEo2yeZ5rzk6HYTOUVlqRy9
xok1OtXVYMlVCwfVUJ9+fo0Or/YEW5QNRaOfiz+egLoO0qS3LQ+zJPIYAX2ElXny
q9r8U/8MfG2Vk273TK+peIhuUytOAfzNcuwBs5NxDz83KfNGAdpAaYsyN4slawqU
bIvqsVQx5JwoGXQuFnAGD2kXYuIRHdjvQGCMZm6gTPPtheebVv7gJwELExkXzMbG
C67MmBDCQMWMvSd6U308O5sepOO2xyXiYprjclDVse5n/QapEib+um6y8I/ezz+r
Yzzs/xEk4UlZ6LXR7EHhCWF/qxQgIA9Si3IxWtL0wUzstHZYy/srDH4dfbQMQstE
MXpAop+YOoLxFKR2o1csQF3Lxddq2LM6shwWYGT5HwSgmVZuJwb+rQdZw3OSluJX
9Ll3+dPgpFnpWWiIBMTJVBCRJrDGnV3WS4Ad3MJs/e60zU6xWI73ThpH96AT640D
YTIAH9zwoX9miFXeoVEUsw089NcCQfSIwfOOquUHjsAV3qV62EhSkvSlg/z6g2Gf
SyRqsQcrBolmTFOVsku3X7a/63nudVB+yBPzOa0K6kpFjhGZXBBx6shZscMz1lAo
Q3hgxfStdi7uREZtCeFIFYcPn/5/Yk2Ya7Qr9JaZJ8n9d+YLzYeB4DeXctOxi9EN
j0Z21TK2eTroAtT0x5E3lp/MtJxXa8fcKnu3UHxeYpTt3gX8HI9/1q98g16tisXp
dKY0VvyIliU5ZiPSygRA4oeHiK4VlYwWpJd2+uRHlu+2zu7NiJrve5AOPIydHo41
zALTohFi+Gvc5jisow3NGO6tWXdOu4hw7wMZHNS5vwgqlbK8ILoGlewN6GCNISWk
BvvyzeGAHwY3YhpZcC4LGokZ/E6UCoiJsfqb/0t7/TRUtJTv7obP/4ZHuJNyAkNz
UyW0H5xR6jTB1W0HWG7nVtMnG7TiPcD7BPLtX2df+78HSMIoKZBeza3x4Sil055q
LMBze0LnS00ggAq2IiSruPov7gpQUyN65dz/vZyrY/mEdWc5HVhYW40cNGIVoQ7e
qLU7zkAiGH+GCyE8AtV8/pDOKD9mJBd7fqlEecKNQBUv5vJkRfCg3/uMWz6b+CLp
8jMhxDXx7CQgbfFdNGhT4u4+I7vDXdf4JBcO2yhi15OpG88BEy930/nTGAE7gw0H
SrLzyIbicio3b/ED70CuuC9IH/4PvYvv+1OYAI6MrtzIHgpEnvL1Od1/+qQuUydB
vbFWGEBl59PVAwTDA/S8DVHMlfPK/8wkkV0l9K0frhLQlHgcZiOSNiba8Kxy71oE
Hk1bg8rrLOjD+8D40moS+uUBMmmbWz4yicBov0hcsL6BztJqanUlJStC+l6DKk18
FhAzQ/m5OQ6XS6HCnC+0y8obu7I4vZBEw6HbXIODiRsRnbiXU0u+UiavMOzfMaen
pkT9RUjD7XZ7z4y9mJJ0TC+YrUB43UNx0paBztCLkT0ZiSP09gfrhj9D5cPC5rOS
X7Y8e/83GtO6wFzsmfxmuY1GkOS5zjNiCry7wk2OxybuX18w0m2oL7vNjzSJDzBl
vu2s3gLA2GYSOXQBQn7xfqLpZcmNeSpm0XY5pgtbSE4hxbfBwwAmmZJbsKx8Kbx6
q0BfcjKTMQdU9u5/RB+2ydMwqmqUOFRiFeAXJjcT2SNF3XNqzoy3aNuylaA1d8ju
rYhw3xSQGiVr+poSLgEbOKGr9UHi1P9E90IVVM0QW17eaCVwgPqTIdcYcjcbWXJS
xjgkY8m5tdaEVVVnhtyfHm3ROT18nzy2Ai9Nv9QIDAA7GwYP4pQxstvu/9DDAreP
e8iXvHc8ztp+g0epnfj5OsZkNJMMt67Vqsqqd8EyWr3ueRnCppNJcPQ4DizwCwsa
p9bMVB7mSm9SwP0x7OHzsOWutWCOh7vjPwq2riyKHKFH703uEOYugqBVt88MDlFL
8vhkkho5L88vMcAMCyiFtyugmG5wbVSd8iUg7t8XHldIBt3/rDjVHPZOetN1Sjlj
kF6lSRBRoioY6G8X++2LfxGnS+Aa3yMwmlpjaHJF4JQ84hHOVz/mQWiNhBBdL2ak
U8sh/nyvcgL+CQmU8n6rp5ezdySIWHZFGLxnt95lZWS1ZPXEEoqQLS0c2A3E+s0d
WdjW+J5OGmhuHItmTYQVL/yKEIbWD6VB+yVVgYN/6qrk4Zmo15sDZxlSVUoljX/a
xUkswehpUDwaOj7rvC2Vb3fvnk2Q5A5naXEHtTKQjpzshouJpha4esQeWu1vfrP3
GovYw3zJwieJdz4Lt/q2JTjX/Qzc+Rnt/SN3pdzw9dUD8IYP5mecFS9jOctgydtE
8sXMXhI5A+u3p+QczZmgu74UlQfBeTQ0LJemeTYctCEIW1DMJR1rbnxSXME3K0D5
+fAUMTC935qfBrfADgWHdRl/sGYp547JRHYGDhgG47JNE3DO5utFHn0/knBBGDt4
KL5hwiORni5IbxKntHJjyh7hMEpnKAjN8ZxnHh/1hEaGoESvHO5kxCJS71d70A6Y
JEILzAOrRc3RmA9Zt9LSQ7froW2NlCuJI0L18MLphA1l+CxJl5LtSIqqgEb32INO
zTNLQISefQLgTy1RS2QmgA==
`protect END_PROTECTED
