`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFDk1taltUl1DUjYWK1MiLScD+1okkNEwRaDbPeVt2/T
FHbTT7cAH5Yt00lURuETZ2HoP+PRdTq6YylSXmh1+fZwD/l5Y584O4QcUO8NOphY
QZ5rEMpelzvyFurmagBgT3A1AMD9Y4n6v6xUtucGcepI9RLWzDA3ySX/X4k/KibY
PQyF97pklaTs/3hZPJMtBucNUrVtZlcrOBVq7M3fl4Ah7nF9ln7fw7cElaHTZlHO
wgEQ5a5qE3dZSDBwJGhaYqpzXsK69VSkC1wrIeoT0xoMfl5cqubMbVZiwky4v1/2
wC9n3xKiKABQ2+sZ/lKVLj7dPY9r7Gu+CCFHoFUuYnp1uUo1YzhHjyXEQ6i1EOls
CCRrz8s0JUeiayoJfACdHLq0tpcCqKMj6hMCOWmUHjcOPP7hC7zTe5DkiaLMysQv
2eJ+EDRsr5cmqvxBNl8cjK/thZEAVRiogWdA4KJNMOrK8AJOwlaepcAvYWeTnzLG
`protect END_PROTECTED
