`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
KO55B3Tl404HJOsoUX46GdMtfi9D/4qBq/3yqr6ZjxRY5QbtOw4+LeN04HwU9PNi
harGWy1HnAbHk5AoDk+EvzURM9YT09P4RaeLiP8+mvgBviihHB/v1WHBq80uNTgD
DkTSit/U4qaqPxrsdamEzl9j/mPo3DRXNiUtB16FM4DKSwjZk6nD98WmuRWX2k+h
NcgntAxgOFQYuZnNoTRGUy9rgXQt7IgxUYQnqRSRrKDZfaOTb3bknLeEcu5/s9Er
/Cla6GEfOMFqM0sq/2ODZNZWb5iqo4SYh7DN2wC8t8zkBx+oqFI/I2W/9rTOiaZs
CB2qM2d9Mf+AXjLPqCghYvbt54u0Arop3yVYm0+uQiwjf/FPMX3zWc6HrWKpSAKb
72I1KmzoMHrFkoNNVOlIRV+iTkuGjqaV8nqmriFfDWTeAQwdcfQSR66nC94vr0oP
2ov76VqIlhY3MxWqy9A4UyPvGvdsjKWnrlepEjUjihI=
`protect END_PROTECTED
