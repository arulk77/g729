`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47bHmEtirgeemY6D47/C8K9roI4qj+QxJZQl03Ikj96w
+SqMm4bsR1f/Qydd7u4T5eCrI7WDsi7xKaymizb/NrBukZG8cQzOkrA7S/GQfTuv
VUDBZkBQXdBZXQJcSK9CiHjdXJvnLif6BlVdlJWhlo6s4BfU4E49bLXxBOX/eFSA
rXDgG3zFUBMGqfzfhettW9GD1+IAZ1FASuXEd4VOV62BIy8+3f1ELSJnmgX7L4vH
4JokQmjW9ZMiaCdMlW9lUnu9u3rkTKI0O6jD39HnSdUA2l89kGgH+UU3fHZe9xX3
XmF4lXmZxBHVTThGL5pgn5ZvoZvg03ubXweiCtkhmIG6VjiPMxyvK5/W07USd6E4
T4JRm2fWkPg5aeqMKE9O6g==
`protect END_PROTECTED
