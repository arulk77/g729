`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEHYnnrENinRD7dMPprUgSA1AY3b6w5Fg44qL31UHD6Q
2EbB1q349bZLb9Ln/r502qHSoOlasHy7ul5XJlikWblGfq+E+WJMEhkGMtEDkt1q
Ds4PRvoZOVpGgsJ6U5aM/UsrwseR8GEP46xQaG4pOtNUZqqMtlFtC9OHkGEsoObA
PbDSjIv2+9hsNJjFqPEAFkHZ62kB0q5goCusvWAA3H5z/qv8eAd8umkr/6iaX5Te
+/5RvgkWD8avdfp4ZNkrwQR+rU414XfpJfKpTPTYPQ54g7sjC5bDCI/T8gPt2/S8
I3qSG28vtzxPHxmAPvpJiYveEVDX5Mm593byK6IMYkQKz1CjwGhM0rVeWFLJkh/N
RscxrlESX6/BtVdCXZR1wlCrfTOOeC+uKv7yK3DjTvxVgK8VisXvmyiBgaqNZ/Dw
QXniBc/m8B+pJru6jirqilbLd276ipUfMdvxrWOkBaSb/cuCa+6grUUtcELRnPT+
BRr62a4LDxAFTIKUg1tPZprhoobpdYG7NDdGHnnqdWSYxyLLt35JMvzXcGbaYobg
`protect END_PROTECTED
