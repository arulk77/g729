`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD6rUzoaCeTvinXheApTxWUJrJKs1txeqNW0Gz/RvGq5
M2hRRs/PQAT4eWyFv895G6yQNht8TuVTmZ1Y6IpI5cRrrj8husfp7Ft+FDbzpYdY
Z1r2XNFm9tNiWXUh2vzbGp2EPR4W2NlCARQaAUwr6y3SptjB7vhbNXxZRoBrTM5e
zSi7J4kS+LwDFvmV8FDBFasNx+JrUrgwFgiu4By9Wdf/j0lubhL0rw1hkDNY3SJf
F2d8v5Vq7xEDhhGKTBI0JhCekPFaW/F3tN4XYrVMehq+bEphAxDFFLbPkPqK3cx9
0r0xXExTkTaF0XkUjEQX3I1bAhOmpvd1QomtZLo1oo2hMs58c3j5HO0YHXt+8ZIL
M6/bNE+X5RGYzNBsAY3LUbaLqc3Se9Nc/Vowv+7Fch4vyARLhOsssb8rA+hODcNu
PAddYXfLw3ojNCFqrXXoeiFSXi+rl6+nZY8ifgh0xG9VLJT3H8H980LPN/kpG2wy
TASLxv5L6WqPvBUgavnT2+xL481UQNQo3jfY4N380AvANRjxOcXtu+IxI/IcEQKm
dwxyFTFHJ3tt6Key8IVsU5v1+tAaOYVfLOoWOMICye/iE/VY8E+9CcLp7dxGvl2m
2ESl453/KWYctNfx8CZzOw==
`protect END_PROTECTED
