`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xgR6w+9eOxsJfEeUhndFClHtaAgmDHAxekIgpWNYDsV
/JbJaqEFL/aqsi1iwoS4AGHpcxTqO08UbTmjRVCyh+CHDOKI6camiYb5vjgSEPUb
7UIQBmCEVyKt2UTNIbKniP5B0KfCB6m9xWqJjLCCLi/0OgdjJ0vD2eYNh0bM5AaU
17wV1FOiNhLSFvaDXTYypqNOw476M3r6H0uYUVRQxEits6ezZqVQG3AXDuMJ5DZP
4YJICvGZZvdsVxpzl5MJmrvcSXrZWoelxoofh8Hu0TQ=
`protect END_PROTECTED
