`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM7suqex5Xhglk3aayLf9EfZTYG7g8MNGop+oQ033rrP
MZmQVYmQq0ctfkFgGMQiKw0GfN2w1cB7z5BXYCxq99c8PcsmNnZ7edXnp5G4HSVd
wB9NvdAbexdLnt4YV/pTgCqRoH6XO0bD74LX92RfQ4zx/0FVRbfB6CNR9uK0+ioa
yUdlu7eDkLQvoSUijtkBk/Z/M9FmCQyBwNG/J9DYnm+DljAJ5NEqkir6V++G2FHb
U1bapKVb7fefi7ZOtMnd44HW6y3IakN843how+hQDSD4ozDo6PyXJxLT41mXslyx
u/Az/VG1u+6nIcOC360pYn2ZNZR0VvH8cUCVXHcx6MG6+HkMQRlkx0B3SUaJGTJW
n977P84rqicjbdZ1NNy1vQ==
`protect END_PROTECTED
