`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAza7GRXYQ0zI5KPCqsNeyFk2J0Zo6ju3/jJEYaDYfEE
ypEtzO5TMOSZ9dO6JmM5CgfvgyGFyBHr1RDz8neSn+64sqNBd0TaQDVsP99NOFab
NwH3ghMBbgqHEETN88U+g6IXkJrL6jN1aN63zu34cDG3dXrWcGZf1rZNFf03lnFk
QrR/l5b0ARpsl4rd8PvQ9g==
`protect END_PROTECTED
