`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49nbh+jThbbWaQE23/2HXA23p+tyLtMNcDZgZtFD7U+f
jtrBnqkyowuZBMNAs8/x6dozsssotWpP8v0gEPEdl9l5yeyXTLctcduPaQSu90eI
HMccEfjdtD0+mC+5NO6n2JXgNv5pYnIYiUECx/lT8B0fYN2nwU5a1Aw9heNFbnRS
fANOPmPLohW98UHu2FRmIHf/4CVtlIcNWwwa6HXde0y5lJIBGkQ0MwUbIT6LhfUx
XJvXqgLafoLEb/OtnHwvtOL5IAuxvK1v+PlkUm7sIMN/PGRlkLy1JJ2Tjnl/yDUs
BekmyLp4P38jwiKKMzkJ1A==
`protect END_PROTECTED
