`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDE5MB3+sQbfvQx5ZORnJj58IOrui/WWOySjdz3u9wZl
V9vJncs9HdI+06ZV59jIMBsOBsX18XIuCAwzLpYu1BB7BCsh4hkuFmmamiLI+rzw
jJVLeuO3ZsgHYZlnaOW8kMR6xb1fUKjfgQyXYeI/beYCCHWHS77l1ZsjaWFDYK53
13dM5YRo8yxNekWNfXWgfXEdmTnNdMUJCBhPoEbehAHIQFXCwHCItgwIyec7FVGT
lyReUAJdHFpIeM07CyM2x8oG+NrR5WohZzIOYq4m1kKSHFgwwf96JUtJVZgZ7REV
5yELcBN/p3G8P5hjkAxcD6ApS03qLHSB5t3NLVZxkUBqUQ1u/q5+0v0CUSkYBOij
g5sDLYinR1SE6/IuvJYthFMDSY57UvQysmuMoqItbXX5xQq6dy8Dg2Uz/qS0ZMyW
1zF9W7W8gWEVrQTMlXJMwfEDi/76Ze3WajIEMRuBEygNbLKzFusWNJlioRT1iiHn
syx278HV8VXja7l6ZKCspymdm/Rlow7bOR9Hv7e3Mrc8+FFxjbQGzUuB6zojq83S
SxgbMgh8mNgCLgaUU2cIHu08PCZYNXnKxiAH/fTZkGXPrxQ+jYNw65HyTMCT9fuz
Svxy7fpHnm+qjEPuqN4PzD01QLQ4RmgoAb03NUo7DV4XtUPk9Y9Hwnyw/Kq6irnp
`protect END_PROTECTED
