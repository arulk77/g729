`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bla5a5hLfJvGEeSdKAWQ5b11XTBHnFqBDxgY+GStcUu4NJKuKNYNvLw2wG9zx2Br
DyWll2uhIokv3gLhz8Z0m1X6e+vwsFvOl2Pin8u2L9tnhK71eaWls8yiZClvPegt
Xf5gK2VrQoau4A5dYW2ntlXEfyjaBoymZt/mC+6fgTkBoK8FnLKYkQf6pZJT23+N
`protect END_PROTECTED
