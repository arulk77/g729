`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK7YYNwFgb1bwZXLwa7Jl2JzhXeK4jyXfBhT4XzPKjlp
zZ4D29qoAZJybwTkI6wdZ0D1C7UB2TmRE+Z9uNlNnH5XxOtBxOCK1xGSqHoDp36T
RxvuDme4GEMUbXlf7soVm6yY+NCa8I00HMnvl2ozrfqpKgwUFRjgUu+f0DrvTb3y
IwIlN5skQwV23N5adzsK9A74ylNVwmxCmIyU6+OX1kV4kffb2iC58jZcjAVE0UB4
`protect END_PROTECTED
