`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aXYEhgnBhX59PJTMMBxsKKmfH8m5cYz/K9mFKNA1LkFk
edHVBSVFwIsDLCxmyOtdiDTwKU6EQ+jEdOPN2rvK4ncbf642FpVnPeiCQSKO2Qp8
Xbdu1FaCj8ID7SPyE0dhaRK3TpMcMI2sdXYk8szgtkeNZtnVV1LmX1n0jmOGtpRi
6Jrf/P7sY26pvfQ1WVFR0RhGuAeZgwd6N9KK6wMym/j/QDnO9ar0maWxMz1q2Vs4
6pprZi1XDt2swodecqAnOPdEPtFTyPu5Fp5qCr++5WZpudEgTmwFJhiOquHT/Y6r
iI0KMK8ipkihwKuDPOU80wargtzqgXdgebs3j8Crzs+tDmAaRXYMqcpds152udj2
xWZDDYd776wbIj6rmunQy25ucNqEyIIvVrwah1M6+V9P4KkxzjJSMVvALuy60Uk8
5ZxxBAgxW8/34RTiCY1Avu8DOqxB5dcUIDYK2wmOwwn0tgTygFIfyketeMmyAoRJ
6NkdkUi13mWOCDqLSMO55OianGPTbBqQaAq3HytULAmt9XWQxYt54OLcUy9KO4dX
B5vkj8i33GHiZYv81PFlWY3VfOOdhMeRgpzqKKPCgk1H9N2ZayvACDVGWOPVcRTu
xGfEtzYkjKDi9QEQ01cpWEqaBUNnwXIcN6dGvGJsR3I=
`protect END_PROTECTED
