`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
6FI6xWPyvBjGtLhF6OW1uqDS4W70X8MVdWdlHfuoZP2IxwqG9k/b1wBZed/y01oJ
nJXPRpPc0RCUrV5EmGDDWtjCHBd90U70KCg+iswCp9KCpLbK1rHs4rAFvkkcK+iL
LCGddOCxG0CAdPf2sloKacg7xasi29NmADh24vmRyEk=
`protect END_PROTECTED
