`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK3MCgrOtGqwV++rqvYzpoqtdOJ/Iztkc7kKkTugJvdc
abAx3VwVKV4LRy7Q1KmrlXIHoKWT1Df6AM/OczsEqRaoIoeRB1ln98TMVlwo2Y5J
nkOnstNxIjGy9JeLovMrtM1v+vxk4JxBt2OoqgdPaLQlaz3XT2PNCmXptKwDEH1L
04A9Suq5xrpQpUkcDaDw3tc+dd4gvTNldztfx9i+sWXpI8yo5y+3pb5Z4ylmcKit
ZK5d/Xs2yqcumgN9LYtbzX1ygGkxMTM4XGv+9t8uN6fuAvry7o7MwiEoOOszwFpc
KxUHuOKIkIkfrbuBnwIgDJvZ9a3FkQh9EsH/ndNyoeySIpo2qtxxGKqQnbEm31ei
008o0Ipv5ThpsSN01nLt7wp734fAKcUNd3JMCkYDFs8qV+c4snrfXK+tzQPwOMIx
TDSg+pROAd1oI9A2iphlNz9SEAsBYc8MJH+wSUkqorSXPd6t9NdwKwklwR2YvBfZ
ZGCZ4Fi+miM+k9O23bygEg==
`protect END_PROTECTED
