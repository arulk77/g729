`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLaC1auRLZ5Xh0uUnzoW14+Q+7RK/JDmqdE/Yx+uJ1f3
R0Jbo1p67wkrNurCP/JR/UZQr6IKZK+IjBLQ375tQtm8NjkEFw085nw2tJ2wMtDq
JmNp9NAnN8VJq1sWxJG8J2NvO/uAsIeE8l3F9/59XFHAKPi0wTxZVP8Mj6jBeAqx
vsMXbYEEjWzzY3ae8WRwqOnCgHNMCJI0sLQfvwi4YhBVWWw/jsT4XfM//s2Yey5E
IsBHCn6g51sVcBOqHwuu4hWsFr2D2MO0a67JaIUdOheiUeZKxPJWy5Gt2RqtXTTO
56FULVkMm4HrSphU0ES+RpRlRsLYjzVek3jQFdDsouGZGvMpRzCFggUo03L4ESNY
SjNM3txNWPq8CGTgi+8MmsssURbAV0bCquTFQpfa4UKOYRcY8ci6Z+ni2VGbvL0n
bxYQd5YcuNp8TypCpgeEBCk7uicJGbTWcLrWX1IgaFwL1ghxNMm3zbNFAGtCfuec
`protect END_PROTECTED
