`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ1t6tRbPj3kfvhlecaZLcsU7HEPPs7sUce0Ttcp1J3z
i3rpe8y3s8FolAXZFiN236BtbGBNWCypwlnFeJxA6Znecl5nL+dtBVHSLHs1rsiy
ucdBRP+U8LavClgavLhc9ozTZFn4Sy7W05hmbpqOdxdCUbRHUaMfzE/sl3LPqnlV
hg/dCjWh3rCTCS4GXym/2fvA4Lo9ZiW47Wkg7JEHH0fZ0knU3QR0oKjpdkoifWFW
SaQ41E3ePspggkmbOXrQdmPZYi9wmQRqpN62EYcnJSqQXrpeFbilzL5A9JQhUD3q
AurHqUZqiL51mc2bO8hxpCXQcd/8ieYJ8UA6Ve2+Qqi/gcI4AvYZmZBdj+pevZb3
tk38SCklMgl0oRV/NGi4TDOHOChI8HxOWqTPEHGtTSAbHLvqc1W+TpBzw0IiVjbb
hH6IlQ13YStBwR0HLh8NW7d+VWhPUMS+tnAIAW3fq3MAremwzDHEAjX5V1QLtbPt
m3VuA30QNxFBgpDxZO8xcV0itTgfHarKYn8Nk32s8/vPn4yHX3c1Dx7dTKXqtqoj
gH6dGHeFIYX0u88wE/ba2nKsHK7mpRg8srXrFnDOHm+si5XoN1SpHBF669a6gc6z
`protect END_PROTECTED
