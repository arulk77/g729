`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
1/PAdzyz277JjC0tVFX8DuRiQIRCLfKvACOIMrV96npNJj41AlkHPQExLFZ1M0iP
56qJdSgVSI8rf1MpiCANEESFiWm9AerYqwuydBQxGT8GTj2wHpEHM1N5wLaVRKZD
EbQlm5cuZujKbL3Bz6//ddyFe5/C+RpwrK0lR67D9KlNoOlS6sMr/geEjs0ZogOo
gNmGEeM907fEBUuYo5T4FL84i2fUTnU1tFp4cjTMRsoq5f8swjoqyKLeBtybWhVS
FzjoKH0ptVnW7s33Bt0NVgRdKxdy0JAPUSIZ12w1LJs=
`protect END_PROTECTED
