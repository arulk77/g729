`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveECw8kuywkxylrGP0PbWnG+0zS0PPDDZl1GRPwb8YJDk
8EnObomnpAEyzghm4dVXT1U8mKbkOWUFC7NKR+32BtQtHcfERrRsN5yep2qYZ/yd
DJgSM7c51AiE5X83+rfMV8X5M9IEJUWS6iv20n4hPJm7EpYR9+vZoTW9QqIsWBW7
4z5fJn9uDTtvwgSNiBzN+CGX0khQio8ETJgtol5sh2bRJh4tHgGZY5p7Y6GTXco/
d7pXPx2toehb1NYpXnwWGA==
`protect END_PROTECTED
