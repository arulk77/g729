`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SbBOhECGTNRYQie4oQJrBQ1lNj8URmPCPYTNAwkIewq6
HVZeHTf+mZ+L3MoO0OYPaiZgwklKtMDSKPoSVzQnvvrSvxxajTY+87bw7OH+4y1U
RLsSBgirMo87xVlx5hmLl5HRzcXG3mIgsQfclboiwlLk3+s8wJSTKEdUQJdE/NkS
S01c2yNCogFN60dJ4KchwG0A9njqC3lgQbE7owuevlg1AdwEw+CmmTmteKlhr0+5
2LSJBpIBEc/IiHCwdUIRN+MdkG+RjofKCXX0cQy2/vnhs9A/f9orX9jQbqg5PxlB
dKv9OiSN/cVOaV+6PKEKExqEy4NxztGpMZcmENTztAJ0Pi4bKT3o/AKkEf2jCI7o
sJKPDBPFiAjPiOlqeNvPRCwmO4TobYRpMiLyul5X25x1f48NJifaAShdwqRiPGoK
taZl5e3w4lhaUxnKAh2fcS2VBGqlm9iciAEogqD+sfYY1dnwpNP0EIMhScQ5MD5Z
ngOzgJF5ZY3VQ4WWYiyNI9JzW5l4U2KZSHX2MkqmpXnwIdu8RNQysCikHuk9rgub
qvds8j996luJMbgfklDZB3erXDFE/1mhoUf3vkVuuuDBV60sJ+uyXBF6M0CBscGc
mwPm+zwz0ek+UOgdXDey/b4tRe0z76vBnn9+w24gCEEu/ax3OejZm8GFYgw2SvSa
2AItiKwMjObYq0zD50eKtVMUSRCPhSAF2uELP7aVGQhG1ujQK+OZ8FND1IWcoHwG
n8J0YPvdE9W5kdqhVkiChCGYSldzFPyNKbeSJ+u5pwfX3gKn1nuTuULRkgJJb3JP
/qDQIanxOTXx8Kr9etMnRBEwyarnSNx9dL8AiXo741Eim6V/snj+8gDO4w98lQTl
7676YOJrv8YCX5o7cbFU8sJgsf85giaXPIDowQOpFY3+cgyLzGUtIsNS+84Az8sa
cz7iZ9/pwiDuhUqCkNqJiwxpGb+Aw4P7ytkROgontGSfDsbV+GZ5kp4zlkLM9wdF
idNHOssl7s2Ao9TmsnT1vNd1lz4jplD8VofJV+0NeelBKlgHNUYsinw8ViexBQI0
mewQ4/6CXpBH8gzgUPKuRwCxK9tkZPLS1iRu8ntvvI0qP8ezPMZDYKjJoVirTbt5
7Gkhg83I5osr580kGgRVUk/oCbtCHjBFipr4z7oIA3S7WHyenS2SQyhh7ON+Xx/d
5tLcMOAFv2uoLiGoBgo9Z5JEWkar8rNwkFsO15kHcTRnlEXrS850Q2mMn1R2LiO2
rL/2hjdpbHrZ5JmC9H68lgng9gHWV1212sGuCWJfh0GRSeGbfJt/PXcuTafhJeXF
i4BXI6rhJSflzIx5ypeN76vamkJFfY/fs/JL47R3v61jLqr+EqHIeYjxvxwgKheD
/6PolIR6vuyeFo1UJrdCrJ2QI2yqIjpJ8U9HHQBJdq7VSuLoETOj6dunHw2w8cQW
fBEZGtTtyT+1URXd10KAO4aPWJA9iUmY8zDMpEWR72FKIRVIEC7LrDZv0PQRClqY
PFcqiopA2EwGMpuQpk8ox7As+wvpCWhl97NHDhl/gcCOdno4g4eZjMjrknGLmMl2
Ys5tRiNNaJT14Gk2ISSF+X6Xsn5UGH1Bzpt3Ve+MRwkND76h0eJwdCF0FIUXb16d
ipxk58/ISIbNLWmjQm/++3Xv8ubQdqtVYYo/ad8otpa0jIHUKr4GiN0VfaN0od5R
au0xwmIuBVVTqxUaVIl8Yc52TXJ4Dsi/uvNbNYmcszD5sA81jtIfzXT3zsCEI+px
Y6aQX9ferOJ4upowSHO87ZE1BcMjugJ+MmQyTGreamZZxHSn1+WuN935BJaztY4w
rptV/16mzFmsk2QkkY3ErQUOgWJrhU8ztr5J543hIvT9oYQ5mrOBeoUt1iLkoqAF
bWks+y93ArCGtHWKo8KUpjJU4xbFLsWsRb/kmQe0jJhY4oeXylSm5QJKukqPRxsZ
YJ5/cfycc+vRs4LZ8hJxYLAxeA1RMU4Kk0XzqGTZeYwxzAz6hNJ3U9kLFrs2G6Iz
mIN+bOMadmHQl8k1SHdVW4fuEoON8ZqQuMUaWJfxeoL1eGNTdeAlL0y5/mJYYKYa
hzatDSOrvQfwRcAQYfk6Xi1Z2cs9oNdz/PAdD8ckTR59pMFRZbt7YXmIqAMRgf1L
ioxuHQmVtDkUodLFac6v37pyGNvz6OG0++pEuB9dolZWvRQEMZhgdhAiFbG5g9e+
OkxTx81cVodIoaa95QyeS/gawJJ3VcoJqmcm3StA+s1JWox1UUnhJv0yjrW5GTX7
qE9bjPq8+RHVLsVKnq9japISBXFue8qEMD1u2LQC/ozwyJAorYo5TZtH79mkAIct
EQQ1kNr2as/FEfFCqHXaRGBsmC+2dNzL1W6s1L3V3HhYy3iuWP0XMDaMFaIDEA5o
baL6+7xcAs6OWY6K0HNQaImpvMUDcctsqFBRE0a/CcBvcTr9TSSqrysqmwZpoWn3
LZQfRJOlPcHV75+d37TvzkPBn0vn0bEgWB7PrvPnv3rEL96bePS3dCBC1RiX8Ls9
t4p/9pU/pMxEc+XKqOFGw+IcBpQoSzIsrkMdDRsHGBYKP27MzJIEThcH0hRaP4p9
MwlNGC4XjKnJAe7XL3w8Z6BioaReEdNguWHyqrKjQmX/7thtEqb3M8d0LP5uF0F/
5Xa+m/YJZvgvkOiztkZbyuqHDLTERlgeXulHjSBQUxlNJfjJ3jYrSyeTNRKe4VbG
5VB7ZjceUpve8gFvr6Azs0riQ7rNzrFk2eQ2+bw6XtoH8Vt7ut2GmWGJiFKg4hOD
vewopzESefNJh4NT3X99SYHj8RA/ct34hQL21ottfXixhtbd9iN8xc4YMd7lfiUS
S2v0Xot9O6HfCgiPebW+30rtqhgxXx86hZf++RFW+PJ+MPU1Q/+tz9H2RbfNqwCp
6uS/F/5IXxD82n1PdVfOeWOIbDQeBFvxp5bt8gZ7PTxXCcL/c94puSWkmVwLaQhV
5o0d4Lw3l9t2+neCOQvrNLLSVGh7Cj9pJjPXlOvxz9cXyFv8hGM+IvmZGFMTVo77
jQ6Y2yW/I5V9W9qzNiPu9KLftn4S2dORpIicGHJ3F9d0TQ/LlKZjWlTJJnMVA+2N
kBB0A9ef2zvhwNnc4XCpbgJnMdLluMZLUth3Xw1z/yN6cWYfET0AqWdXVqQSB5W5
IhWFJPdGo5uOkyw/t5lIp5OtZgLZh2rIcZYp2Oodx4fgUcr3u0O8MTMTncDebkVl
nq6ecUAqWWQ9V8iMeesVG5EI+A7ttB0syXi4ToFoMIaP463xvsVIK0XEUteLzayK
RqV4TJ+xTf/Gr0TEX9C1AlNthBKp2YuVOhxm3apPj6/tRKWXk5gSy4ig+CvDE+Qs
SImUQSGKjz0cw6uRKmeHLY//mjZ6HdU9ZnLCO4koi8IatVIFSu6O89AXoOVEPbew
xZ9I6GiHk9H5FWCDizUwkw6+y2o3QR4dXsadTx3kWJZzqc+PYSEJbB4C3Q654rWA
9saJwCjP3kLgKrlKuTDq0x5+X4s+jyLHldGQB8Fn6w4lzzTM4mgyAtu5aeHwA25h
J7tgftFh5LJg1gfeEbbzeJFOr83drROWrCQb1HJPh1MdY142Q1m8DKRcLP9nQlYp
14q3zaP5QyNc8fB0pKRjoTAoJX5NWuUyhfDxSMBeQgS/Mhd1kGNI7BrN5DTppvb/
P/0RqDsqNBP/5o5NTffToOHLVHfd077EsqkoeWMBn3OH0pZEmiE5jUrqS2Q3WF0R
v4kN7mg0/fpTMxGmBo2ry25c8ZS8bRnRT7Om5WZptOzUt0YtXrfNUD5/Mozknppe
lAcihTtd8ELA/vjZqDvj8NspDbdd7wF9AuNQbhex4jqZOQbqB1h/8StsOr60WGvq
fr9G5Koq3U3vQ5nDRJFGtuOHh6XPaJJQ0r2cn6QU+2c8EStOu/cK0VAXUSAGgQ7h
dsbbQnL7RmnTvosumO7UNuNv0VeeZ9Aqtl+FT+RSh7o+HitUqN2bF770Q2y3A6Gl
6PisQFeNsUh3IlTEMXVArsTxle9SDMc08vjb6STddRNCHDh/oU9SpQltzh9o5FYi
QzHY3WlhubdBs5StZDdBbSWLWwLb5CDtR3nKEW24S+b9xXWjS9uVFSYIkwH/6AGU
sV0tBT7CA60x2R7+6aTF9MzeTargNtOzJP+LGY/lskL8jGLEifWhar9amliQaG1q
kwBge7w5HsgYCWQlmXrc5P8jEo0OjyaFiAcffBfI+IPc4FzkHNfIVImbZeNSFen4
6clDPw68/L0oykxkeAg7AWUx2UfZKIzsPYQVu4niuLE9l3NLCwQxsu2fB3DTNLHw
xw3RzBc8RA8QtxkR96fyvtysDLfExSR7Plgorxmuu1uhtVD2M8sCiaEzOQjt7X4c
fvBrkQhhuh3VliTREXmZ+n1FW0kBuqKKaoHkkaSEaAr+WHjqsq/J5P89KKZSI3rc
aO7jyT2LT6sS3B/xhs5ub9Gzcf1n/HZqZRWj6M6Va7aPODyiW7N5pC1VlgXCyydz
pR+t2DcrdIjw/l5+OkvUSOi+Q9Xp85oaFR87o2Oar79uj7xrUDnNuTkfZFvlmoPJ
ZRvLaGx7GqQBZtVrfCobXGfIr7+w8pz/zoqbOe7Qy9WpkSGm1uwLSas7lRGxhL21
9a666vdoUesnRyCKQYHIO6mV6RE+T3VoNRiL3kyERFS7JShWJSKnCKJk4q7veDIx
YNvBzVbIgMzzk5dpjStiXqtfFPTDPkz+dXKAkgZAKFC6O22/iQ++5X8Oa4GLy+YK
mUa/btaLBzGbfaEOIi+BVduuDhcX3NoaBg696jWquGlJLIchhPff63seQKKhtyaw
k+e8lFMljqqc1AuVw0TvwmamLGuXW44trTs8RgweXSHKsY9cmKMo0+Pf9SwjIRh7
9t/KTxN/jcYFL3rkNGZ7B8HIUpwwD5CGxROShydIaoLijaZSW4Bey+ditXxoG841
hAZetPcUv0XRgE5SiFkjQJD4mRL8e09GXb2RoeaeWPqRdZcKCa333ufY739axK3s
mI6i04ooHgnk9TEn8orH2BzSMiRKPcGqyRKdViZU87ped7gqv1RvE2kQlIzgRuT1
jDCGL690H+X7hg5eBxbxNJVnc72qRBQmDJsxhtXdncRk6FQNzgWQBvVwEw9Ok4Jb
6JRbPYQ6Iz08o0qdtBUOMzfeSQ1YQKeDx6EMnFpYhk31mZyD0ldfJgW/xvKItHmQ
KsgeeKnCT385ZLQT7xYHOPGKZJbnKBU28oJ7waYf+7HtGqHV7BJI4oWOvAxCwUYW
nAvvqvzNnzgAGBadD6C3gQ2+39bMrX6G5Hd64VkxGoZtNPcZS6t6dPgCmsMtjdew
Ldp/wD7xBYXiAKgRUUlZ/OM36kFPksHjp6e2fFEIenUx50wFi+JPwJnlZ95rMxZI
00aTqd0rtZTJpWwLvoMJJfyGza6eWI8myBWYU5NHNk7qA8wR/thDShq47jH4pTqp
TBrkp68ji6dqZQBYDbkQh2iOje2P4rl0lZpmDsAH3zS65gj2Azgm8cYMe7r8y+Oe
fFyJhMiCVSO4Wsgrk2/nPfXjbTinrxNePLrtkA3FlLeUeiLluleL2NI4/FkUaKfX
rEu+QvECkXaSv6BHtlS4p0uV9HQOcxg9VrlGQzV60cZiyGNlZI3eIDjNlklcUBfH
zltS1oQsTX7161nhiWjHB4wGLV2UVH2k5zsYF7Gt2rBst1rrB0Yzcv0fJnTJEz5v
AhVC3O2pSaYvoW1F8kknrQOUTX4+i/oPAk/SKXqux6Nx5O4sX+mEAzHRvtINoFTk
OS77aBsVWo2j2HdOnodnQdEe4lGUeJ89/STYY1CqvHv7WNXCPihC8vjRxbWc/+dA
FsLa1YADgBt+EMd9swautd5cGYVTGJWKK8D6eM1CGLKDXUhUDwN3voPvyA6l2ohd
0UA/VGPJ7Fl55s3H/ElRfsWaULMFR143+vy5xBnLgeSReMlPAUsbTAIPtRAmyqV7
oizeIrVsEtpmttJJYeoFxG6EKH9Lj8Tub8oawcXQlUPyY8iqhUNPyJEqLdiFwlfw
iNbOmmpq5Ts9QkN8NmbTbmuUXnM3bPHTUthBpCyHKf6+80QsuofSD39Cgs3GdSMm
LNkcKb/wa0kKc9QYjqY0tnsLgty4bYqyi1lX1JeKIYZ5ndszcBesXqWOQTsXl3Hr
n9SUP+8XSiQynT3+2m5V8au76xxeHdfuxzola2J6hcdFaYhDmVCSXaHzJ6F2rq79
kord/SlVqiFGnIkowjXOQjLOJFMUY3sKqhHA+fgiCdoQ6tUSKJsl9zQKQtf67qob
1QpA6/E3o5Vjf/Kl9ENCW4K0t9/Pry0JBsdX6L+M8RFncp0KyrAusggzjjIcMAun
`protect END_PROTECTED
