`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
LVK5YfpYl1m11E+jlNVT8VqRVQ51dqPyFmFP2NiXfTBsfmdrYqU3gKqh69332ps2
+GJQBD+Jnh+pn2J5b/YS6cxqgd7PZBAeujTb20UzyMzdaZCVqpaxfq2jBFMURKAO
16alRzo9QxArwXCASBFDgDKNi2CVBu8VyYaQ6gDuB3ljr3PTWuJltRePWCSwNXE8
7VpAyAdfRwEFyYb+EMO15iqwxw7Gv2PvYfTepy4XxX7sMmQQ5+n6oJAHhMOuakRa
ul7aSV3VEbgjGnP+8iUzlW+8VVH69DKloIo0K11CowE=
`protect END_PROTECTED
