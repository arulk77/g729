`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43Ed51dOCws7w1JT1txNFsPOMvATZZU3c4qsKVZ3HQs4
epg28Y4Blht38pDqenJJr4/FC5OpQMtJDAKgdqSoCIh6rHgMYJFHtgHEUz3mViNH
t+7EjQ8wFKniRaOoPVG/mGCQQxEtR3a2nn7peOkAwPW4y+oYI3LezLShXjbIPeyO
8cJ3/NhM5kZvxqhYOD0OxPNLMtFsg0wdaasqbpv/6xmfiSQUE+klQ/VKk0svxGUH
QrfY7HT5FqNv8itGnwU9Xj6/nrq67FiRdyRRWF3bNgKHT/IA3NTXkR0l3I8uQ1qu
unCmFoBETBU16m4v8oQpupcaW4MjfMBx3ZYFko/Evy/ZZ0+YUCxdiFj0R1/q/FDi
pm89J8Ct6iWXJ7oVXbhJhg==
`protect END_PROTECTED
