`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGWEHKT5MGZAsX+dGzFwbXPZV/6DBVVIEqWaKtCa/TJD
Z5ANVCLFmoAXzC9Ech/PngjRpNQeutzU0OBl2MgCA0vj/ZlhxjFTc0vROSN6f8f+
dbLNJgeL0dud3+uz5HKXeJ8j69OcHRGrfDaARFRL3ExrRod2E1UNYIrrEROX6AXr
l6BGi/cl+ifbEIP3bPX5BA==
`protect END_PROTECTED
