`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCa/AFxyDd67T2jFuAy0YS0FIhmiNMcB6peKBCbdocJt
B3UHNSC3Et5m8oqc686qfWB0kaWMj+b+zUV4iF0DLFd6+iL5rpWF1O23Pj0NCwux
voW1Quo5SFMTiep+tKYRkXbvNyfhBWa51rNosagl0SqSZEbsExMOKQq5+7URqL98
sNeK6nWlJU67I2Yfn4gJULONFmjabO4j8qD3hEBh+cL5EOf1ovsXhTWsmeN8TKGB
`protect END_PROTECTED
