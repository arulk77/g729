`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
if7OW3neLerq5QTb0GME9yStN3cZ3qrijoxCm8vuEhvOfVzmvZ6nYy8zTJXysSsD
u9AIDCwFizY4D4k1UzKwg0MO9pxyEo1yYJTe1Y+7ExxUJf6+g6btroKk3sXklwga
2JttRFL6xAPG9v4qWerj9zvy7AMFN1PXNWzcD8nGxz4OvbdnLhdhiBOjlY+v93jF
x4iiQEjKCWFd8a9AOOEBioKSid1eD8f0x6B1A+TWbYlzyLDQVhKTC6ptb6vCkfPf
VxVEb5mwB+InjwXNmfIoKhZXEhJ1fLu6JSg8RH43MmEvYbZnnWBeN8F8KCbkw4r7
fCDMLTjLNebEihIqRglEDwQJ9IaJxkEUUNzBbkP9A3hHva151rOaiUbeIkv/RIzh
`protect END_PROTECTED
