`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIl/fOcQ3Wv4AxkJyrzYmOhe6zP/JwGbrXY+LCZZHljO
NT1mdve/YeY466Z3gY1MDFeV8pPDxVAZ8KhV5/FemIVxIMVTTOeIzJq5DPsz1kpI
dmFOgroNzF4jR/UAunsenm2TxueibxjaWSUfSehzMT9FM77A1SbiAsvXAHdmmOe3
yVXQD5ySMpipFRUJYVRXfwLHzHbC/kFrwBnaVyNxAdb3YIWnzSZRmQqPFkllI1PG
eG3RXNDMDoeAxJVH7z9beA==
`protect END_PROTECTED
