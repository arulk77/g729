`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45n3pwCEUP6xRf+7jnByE3g08oO+DKEmTfvBXEJbz1UC
+YycxSsfSdVLsQPiez4101s/DW8aUPA9GbBOCL2gKttayKyWEiTnxEfXxISNEoI9
DsZn435xS9anYm/2rghVd5D5hduk8Pgy7FCeCv/0WLvLWTyvT55xuhOlW+bTIXhv
TbQ3Yb0Rrq9jBx+XX+MTL7cuKTlTfEmhpFwjml2KShZkq2LXCD+JzXHUNvKQvwK9
GWktTepibOtTFvKcTbOj9aAFt3O8WniguP36lUImoFM=
`protect END_PROTECTED
