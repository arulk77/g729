`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOz6AVWxwLRlAFAP69pZeU8ZgRW5/hqh4lzgfVPvGdcK
a34EFA9AhRm9uHAxhSya0AgbfIy/4zCyYFrRkkfq/H0PdU9Xt1L4rjGav/JD8ib8
BvLqXvyv+5anrYRLg6b9mG6FjkMcfpfpAZwEEekmoVpqmFDIQ4yftfC1WH8cRd1A
It6sI81P8R5eu/6RRu2HIgAgpW3rx4gu94I5D5i9RydiDDq1heoAfXnJoJMp+73F
zL/WjUCxRgqH9wlDc2TVIKCDKc2fzNC6Vl5owDysFuqwpPrMjwFaamxAZpxZfjpY
KdGVxD29L2H25Seb/Ym4X+xNn3nfQwbB51D9aw043PKuyKjiiSckToC9lKTcu9rj
PixpwiO/eb4BfNKjI/+E5H05drkQQ3lvVDgq73JN+DlaeeF8B0a1TIsrmJqV/R7d
ocDcjtgkyuSe2YZOzdkaIPfBJ+asO8ugNskop6uvw3XkrY45P6NLBcK1EPhT3VLs
4i6flKZ4ngBj95MdYnH+8M6iQymZB854I1WWaU8ELtTAbQWc7fA5fYkJbGKIZAtO
`protect END_PROTECTED
