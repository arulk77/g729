`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
SxlBAyW+2170weCf7zjfWm26gfzOCWkEhK46grNNQj6sk8gxD7aQznnp65VN4ohG
mMZK0kzknp433fBmm+wJ0a0tj1PxHeT9T3ErKHRK7+RCjXIzGep+bOIGmOoCca7q
rssS8gC8hPqlu+AK31jjtKI/58aZX/nBQJ35mX0EAreyAp18zOL/ZAH/jwdYbayF
lePQjLI89bc6FZ6SDrg/AuHoRou2B78cAO5CUuw2iSYpgGL83QIBbi5vY6+QthiV
54451PSqUBvgqvWPEhroGRahOeXjB4AMOMj7hWRjxfzkxPDZobo81dJ0rSUEAfyK
3hNiI3C7/sLC01zlU1TKfd/vWXMzS3hWe3fHYxhs/fCRwS18OOkc/VCuIs/GuLHh
qv/FajtnXf/7YbXwNz4VQ8o+c4b9qvTxm8RolRHuH7VhbGO5DvFnd8qjMoxD3iCJ
MOObpHnMt6T5TFT+bPIFon5u7vt9lLh6zMlq5lYiGZMPXtbRIN7CDrWgZ8DRfjuo
jf2Csi6jo50BTTZCiZOouuxnR6bJaF6Wfw3XgVkxtKIjJ6vtKYpD+Mk6OYQI4hdY
tp2JwebdO2PicMcpJPJMLWKd0RdUvH+V45KAnYkqM7h416W5Bl75Q+dSdSsgJwPB
z/SC+y9ySKJ7oQFVgpUMQqE163RqA0buGvwGOJy6k/7ZUSWg59NLbadeLafq3FKk
ZdaAqc9c6r3k+Vgz7LcnsRbbJlNNhGk3UM1ib3c24LxDWy9Z/+2OAXz9Cq+3Karz
i1WlSQlTY2OtpYIb5CifuraxstHWOYnBf4JJNsFwOMMypsZJN/Xb+xvsJwtTPoSw
RS5wh8IGz/81q+umd8liiEg8qMO5CcS+r5ulmraQRnY=
`protect END_PROTECTED
