`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveICJmZr1H+K41CazIFewjIIQzUc68dNNgE4XaaWUyvWl
uLFdrQfEC6Coq5HCRE/j0CcWhCjPRQc1L3NktgSfQolaAONSLY5xTm6xKvFrx3Cw
7mQt2FL3pGwiksKsbcd/N5W7MOAghH3E+fEK1Po4betuvmol4GCCjB7vCoYYquiQ
Iv7YfEwI6OIApbiFsp2qtUAtiAx/wWjtigcMGEehdZ7mMHLFIMo1puGeAHfWwVtp
RjvZgFkViULioaa9V5QaMRmaaPa6qFGoE4vwM51NAJi67H4BL0yc3YS5GDPwqsb3
WpsYVkkErestikDXXVqqyA==
`protect END_PROTECTED
