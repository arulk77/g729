`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFqJoP8BKtNKKh35t24rOMtvO7wkcaxE4oezjFFk+QgS
FDXF9lQ2HXx+yUxQqm7taU+oNHzbJsJg70WIhyi0LUaDoZF8oY9GQPVY6XsULYfK
bMkhfKrkd80YCNeeBLdKqbHbd3Mp/IGT87iup3y6SmLLGNtFow9UQwiJbb30Wkqi
Y/DVbQ9eqZ4Nch68R8XqD5LbgnDKj0HpwFjH4LHE8cIPtipDM5CBKDHRKvVqEPHH
UMqH+JxFRI3VASQIHBfqYS6jnuH8IWBZDqpg6LefxE+536zL7YXsChQn2DPrgxIB
ndZnmGVNuLy7hmsCffzVAq+YB3Ou+46aGh6mb0C1FffdZKYFwq2h+FYNVA+Fl3zv
x25+t7eEOLAC4hmKvw6xdr4WsBHf+MkzJVW7vMfh7IrbUsaq0xlN00A/M334El3U
0+yAvIMxScAls93rWWu2svnAl33oKzvM3UX0czadoobuzYzWcygg+SgQqXEmG4N9
KNJ/+ZfxZ/xu+/MFJM8qE/cCHWDqnAdytZbo8n8dbcu0y+/0UeDWjN+TSM6rlbB2
X5+N+VWb/BG+eFgbu4e2a/eCACplXyZMuFjmAS88CQryy9MhVxc2kCXxraaArMBV
P/yncc7IAcPJzvxZYsSI6AYsI+mp2dQ7+IjgP9HRu0/u8sRxVwb00uiuoL0ivgQE
`protect END_PROTECTED
