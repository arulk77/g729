`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
PXDphy6TzYfl7WKPx7J2dw/fjD20iJNewt2mbw1yVJ0kN+K1QAtf2c+ivRxNipCL
YBiOIakrk8dtGF/mPoo13MgALyu1/e0h9hsTb5s9OpHTXee9sJi9bmWr5lRNqzhO
19LVsTpHXSFgpY+fFnRTe9B2jFdFRRG+dOYEMelc06i1Py/eBojpKv/+UR/icGVW
FUSjRFi7qikTYW9kKrzSPTlxfVXQ0OC/eBi2RycIlRgSN6JVo+bAaChVTcrwrSHk
VCdSgGgOSpKn8wrZIJd3pamWZOVyKQQQIhuZjtbvMwf4O8ObyvYZMQ2Jo6TdD6dj
ag+CkGL92FMJX+dD8DlYJl5kp+ulHcHQqo57asNzvA4=
`protect END_PROTECTED
