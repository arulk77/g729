`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu432gRRcvEgr6XwCP1VmLyUA6O7Pz6LR7m91yKoQIR6qP
wyZ6600TDeNoF7NYlIfGxGQYaK9/k+g5sFO/QsyJ8Uxs7iie0gMZteIKb4VwJrMM
0fttUof9ZpTMghgnzdpnCg11CjnMIdzNV5ScGEkE5CPtEMt2KWPucysP/cY7V3Gm
0X+m9yMUmKiyQGfof079AQOqKgWg3k5YjBZuuNwu2dYTpO3app5oPKQqs1fNV6ci
R3MnY0fWHVMSjuRfnjpL/x4mfQXoDYUQ88XSktJJQDI0VTEbd2OELjEzs1o/RppH
hRiP0E5H58F1OGiE7dllAd1isCmSBpsj3MfH3vII/Ee4D9pFeM35ThqcAI6uIEW/
MJDgvFrNi6yKuEmzwUC+KN1CaxEAE+BU6PL2pNnNCRWM/ZNOJejHM1IzXSXlYv4X
DhG20A03prZfd4AM9Tg8NaAbgwEADoBHBqAm/rpoaJjiMl50Va6apSlzQQ25+BYt
jP96zS6IfkqFZ1d5KJMB0oRB8wxUzH2BDWl5+PvXvZDAQaVuNpIEhSHLxtNSxF9n
cb9sWrao8a+LtPARDZvcFVb41jATkDiM+pjVMrcnQ/9osgUqlQV/vJOHvlwWAE6D
fM7KcYK7Owate82Rs0jsOc+GCrNTLV4puWZGIKzskoLLDbcAic/qJ+QrQ7x/ArnZ
dJ0MZZ1cLjYo15WeyF9KTP1aItN5a3WAEQJSTh1amjk=
`protect END_PROTECTED
