`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
r4f18uklpWYn42Z9djpzohYupJNIfkl+bFkjWt6Tc8MnHho92EufsrtXAorSZI3m
zttlWbLhVvzaLQxbL5f0nyseCyxIIKvqLuWt9IT1Vy8kBO0Eq6ephzJFhMAi/s61
JBuiT0lxO7DEsJGnScNqy3vIem/jksWSY89VrhCrw54vtPn2J8YpS11P7WlLewyQ
i8SXj2u7vkT3yx6aVQjrhQzzrVJ0eIQlnXWoAKT0EEB2+f8K8vWq5WUd2JxG9ez2
X9Mg0hfWOkbOoroYJ5vkXL7JWqLgM0Tuh5ODP5BgpSFC0vQFVCp4O/4i59icwTV/
Kh7bQRbo3eoglOZWNziSGoS/IWC3B53gOMj3lSFODQWLjEgPSGUmwDzF+uReRfDr
TLkvPySYxXzsi0AGRiD5TGDHhTE979Sc9qCnJcLR/hbSP59X0cmbial8ihROsYr8
B7c5DLsdC0okJvXG0ukGQZ8wVjWge+FMEMZRN1189/JJnmvTORdNQqr1i1ipDAeI
N48Rp+u89QKI4HFn/M6gXQ==
`protect END_PROTECTED
