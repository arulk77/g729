`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGdAVF8hhoxPBJvzvMoNXnIJvJMRu3uv/urueonfkVKp
Evmd4YrvYMG7AId8KpqIbCh7xQnxqgwUM4gg2f9TdQWkjq81L5g/Pvuo6kMlDa5i
K354Z2cER5fQkj7stlqGfUAxFBqNMFQ3DpLpOOyPeFztOXP4zIyHQ3DUrM0D27MU
M9YdAE+6mqhKKngruSYcVIJfORlK5bPlH66dOJ9i5hNUKevl8djX1rNQKrhnex8Z
g9zwsEXNogSYbTiQbvHMt4XJtbBt44ghPVcmHAjdNa0fV+tdA/mDaJzhSlpq8b3a
rVBenNcqbgTlx9Y6/Zb/pGz8HXjoPIc9huOIZDvXJNDxJ7j4zoDSgu0BV1muMtRJ
bRkhxvSCrWwTQoAyXwhuNxT+/Q38/9CJNuox/PwmlPcCRJ7ntogzEQUUoDOaWI7L
FnBl2CLnckY4mXQltRHp/p+59FBpqywwg8dDUm8UAkMimmgirJrOUeE8RbNsglgK
kTM5ESrr3Yg8o+VjDHT5L/llXqDWf19+6pFi9ERyQ9dtnpBGzvmWzF/xxiWAY70F
zLYESwtN5Z788xjdS1Uzq1aCycJObRib/E49jLbpq1I9oYSyXMjuXdVluClSxZMd
Q1a1R4sBAuX4NgWd4pmMRDavTPZUAINQwL0fDhi/2m8MRnrD4pBYdr4wzaTdUxUB
mQIbPzoZ+p8ZuMG46jaffrxKbYLLx1PBOoSxIeCMdtjVXDSYAWjLb2axyWO+6qB2
PGe4iY4qSGTWUFfoZZ2j5DMQmygT3emV8beLhv41WdRtF2beBZLlakQJ5mUhVnse
HF6dW/uYXDXWV6xV+dMslR/z3+pWGXPjetYd59RUQ35ZKHYP6iKoDmQJlA2OxTNc
4wk1mEjKyGed/+l4zBFkBppCgpolK5pJ2y18k07YGzEJPOBk7GXv7JKSwH9XUSPz
MvSL/SnlNrQmjs6iZt3mJX1LSkRohKJsf18ZggtXcoE0OnUc3wBs6VG1gnhDmwCV
n6O9UVi8bU8Yn9Fm/4k7EvS1Kh9rRv8VNzz8rGdzxx0hsBQCPdrcwKxdQ526je7U
3DE8yNdRIJzah7cJC9PSHcuG1YjFk7Zsl6h7rh6C+arEgDATtez+sfe6TaurzpIh
CgupWwQ9F2zyYouxxBYE2w==
`protect END_PROTECTED
