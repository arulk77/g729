`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBPka1FNaNirEM2tl9ZLYKntCm+9WmtWcwiYGyIL3WFu
GUO9pQ/rj8CTDXfjyrZFry44ar5weUMFFjO7pEU6MevLSRe6uJKCV0NQcApAW3O9
xxsR2BMZ6K13b2RHPlVb3+dhgWlBHsZPRkeCoSJPemBeuq8N6YEDLf40i6kIba/t
upl4Vwds1bpB8q9NgyX7LhovzjUFytRnWXwbVn27YvOO2uG43NYxs20A4E/BWNVS
c4BvljN0L67j98ovbFpL4i2uwQ6gFG21qDhH/xFpJbxA+X8fZDvVgoahScT0ipVG
UsiLv0ARjS5J4URQAWOGnb5xHn8QHlgSMqSNS6bhyB+HgZqKPZUmyBG3QFB6ybTm
TGMkCKw0vXs0Kl8SEMnN1a4vA27ar1zK/NFARAW57W0qcQX4w3xcb7KowkE9cocB
STuDni+20Kxyfvra7FB7e3tO1kYmlSFENb64UPULR9+fsUfY9LVjZdrCQ/MDZ68j
zJtMnIwRE7bydeEnU94Cr4uNjoi9t0tae6DKzDI+0CMIhqMYB9uyXD6UXSB/KpC/
`protect END_PROTECTED
