`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEegqu/Kvwnrrron3rhXIxtrCrGlJ9u76fb28fRR5KB5
qg6Sn/t4/Rq3QFFUIZUWdmzK/A2Wbt0RApSFc9/9SNzIOeUewFrzYRlMKlSNwRNM
mrPl42ploo/RuFou0ggETkckZP8rF2cpaTffjKom3vdrNBzZ6i03M3IPFcGnPEu6
S1ufIX8LvFRH7ddFQOW4zNuzW6EF6tsEoomh6MQW1s7xO7Tt2oLRN2U3NoRgdAyP
+YKhNt2AX1Iul1vsyvKB+Rgmay1HPkBmAMkhvcMgsu6xEWrNKjyF6UlvtSPRcki+
JtMLdqpYej4n/S7cGYmVtdb9dqrMItdZ97ZsbveGDcD6JT/xSnU2ee1JEEHrboIK
LZ9taSYaeYUrKsVy3NhMtQn59gmekbVN461xnrarcqzGjPP4qghgHpKC9y5dciVW
XBgSqVf4qyc+U3sy0LGJ+frBEstmZJI75b6EbkMdoTgj6C3fxF1pusOYTf0/+Vgx
itpYfi+Xb7RUq6Y+/MJCBfJO14M4X/PWry6uJL4GiQj+Lvn50aLSfm8u7bsgBw9R
G/CR0iTHkpoh6TdWH5FhAg==
`protect END_PROTECTED
