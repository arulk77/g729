`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42akHXUa4I3Qwod93k/bnpw+0Uj9LS9r2FW0nV0oTjl5
M1HPkgto29JyHJRVHnn639CyPk64VjjFz0omUi8RYf7zrxcqXqYY/wW/sVoIqza0
qHJ1xX07VuXrxo982L7msA6TjYCgNkdOzwaffBdirqXnS/G3O0MBVbHNQhwZ+fum
tgfSgjdBMePSBmTg0B6Aeq/iLPyBkcUQ5l7Oq62BPLZnu7FsxZZC3XAWVokZhbJ5
Rt4X+cpjST6V2Lx/SuCvcjwnQqZ7Gthh1bG64A4AfxkiQ9+rkl+kCNK7ofeBqZdl
W3HmVIlUyp7Tv+ADxOOHcw==
`protect END_PROTECTED
