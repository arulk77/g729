`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveC+fzb4+RlrKbLJOXoLm0vFQD91oqctRIPJd3tCQ/LIo
cCu7Sy0s5fse5LwKCWssVwTv41EtKy9u4b4B2nNcvDM/4LwggZdKI7+22LFZFR50
mCiE/HLxwkX58t5kFoKJ29efZft/lA63N1ILTzhARK/uTtG89yKHsugRyY+CZkns
tJl4bZGm1v6w13Af429dIR3Ib3hKoRXbwrWHWdjICj1kdE9Fy/i6lse2P4yezjjK
npy2Cs9v3C68KrPrA7iVmpM9sER5+705Tt7GV6jWCI9HGHUMhKuDS/MpLJ+79n6h
CnRr/JOgJ8UOjLAswoVJ7r8jVtr2Ih3OxSEQaounMBQqxlI72CjcsOa0loq3KVg8
SGGM2Txm/8TM/tCvS2qZ73mk7TNWko4Oz2qjuFXBUE0=
`protect END_PROTECTED
