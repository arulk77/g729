`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePruqGg4jfFx67uhB0dWIQdi5YficUxzYYDz43/BmQMQ
c4+sP3t56o56cavNRKVZ+b7kqRDBmaG7wQlalQzL0qcWyXfRoFyY+HUT7rsCb6wy
anpwOeDg3/LUzBa+Wfv7qu1J0UfMoJBjE6cGsxg9oBZLm6p7uUq/pR5SMGXz+d3C
+DY4VNoEH51/1oQBdqXrf9w6XkGKXEN1/VKCXNuQoejbc9hZrClr7aTcvU8VwGCp
PRhBPp4pDViMQPwL/tCK2fRD43Xvjd4WWGcQU+Vx0Yri0ngRByvCf5WdaeFIedXl
xa5VQbrFB8r2927iyYjeZg==
`protect END_PROTECTED
