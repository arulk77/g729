`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47gmVhQQMc/uwScFeOFh2pcP3PucevY5m915+auIsID8
Wg3k23IlgRLCKknyUWiWOsR+eBZ6Ml9J576Gk/ZwmfIOFep/QFhQ0K+q+TB6WrJ/
nfhrroIqoLGz+Okft11bwBqHlTgtYfA/1p1cHfemXxdlgcgM/ahNkgvf9QjbFVYl
PRa2xgsbBwJ9iIzw42bNfAIQf45DR7qmutdbIRraiiDXE7IE03glPqzcoayMz+Pt
nxL+WhmjV1Bj7mVksH6u3Bbr1UHHQQmYIllAr27DQ3vSCdH3Ak30SoWjfZBDs2ki
YzJi3pTWgL/trr8DvgCQbm1Q3ON2K+2nBdPrm8Jxq/1RU9Cq3EoWayrMV9CbxFQ6
5xjTa5D3hTiddG7ip5DJ2w==
`protect END_PROTECTED
