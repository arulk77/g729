`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
7d04v6mXxif7TTOwRQ3rSbphfzmc80E8uNsUxcDJaFwQz6nGOYrT0fn4sYKhZw4n
zxwpe5GWZjbFRLnrRh9rirJWhYvb0jnkVNbf/wb2BQPDUXYuo/vSVKqt/NRMqzgy
cpw6hiR7cl4EMrIhY0PwQ2qHNryha3SzU9N6c+Ml6GkIYc7YQiXG+D0ZNDGpLU+8
dBVeuza5VcBG0RgdGTTGj4+rIWdFf2SirbVv3LLglgybkV3W8KHy7uzwuhKXTrMI
E/HkLQF9eF3j/g5gMaaRJ00BvWeagcSGRUggQ0hl4SE=
`protect END_PROTECTED
