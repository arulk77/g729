`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDpCddaLnEV4D5y4wZs/wAc5CS22RYdQtrGnOMWYWbkl
dBrCflbYlkYyOoXQ6ILFraiMPECQz/JaxinpwJ3i4P/+RrYXDEF002qSDm0pkPsZ
KUl9YhdAlnzUlqoN/mhUarzXXZYom4wv5D2djqTLSAsm9VAeqVYmkkFPbXMh4mJx
+rPBUIwzY/GGUNKwnjEiS9XronnsNwr6BQPA3zBfDFOPrrCAjcUlkK/WFoPUbykS
TK/W8Nxo8wA27w406nDXGdDqPJIZVEWi316p4wexN9WelekiHyuns4G9/eg32BkS
s2M53PQEATR9lY7oNTtREMrpTJUwBTEV4IBXxS7Cc8ZvbzYHdiVByc1MtmqKXM7S
KOoeOf9UV8Pnl3uTA7gwpG4/AoLMJOl6LM/7kzLWAC1IKaTqfe5MPoe9BRKYoAI6
ITzI4M2Zr/350fVFHRQpw7TJJ/gJDy74LYug2kHNCpZyzHsUTkw8JB8GSiPeE8ek
8GnrxJ34dF7mOofglgTLFArizbZbivtVNYUPQS2b7+QG4Dr/KxR1VfJBKeoA6HN1
gNnldxmGuW2kIMIRksJylqtRZHAJgNcUyzfwbPDO3sxFMAhVyFn+s3pl9CVmtBd0
YEigTX+n19F9UKI56Rle14SudYo+QHAgz/m62/k9Tji4uJs2p86DCTQucSlS5EJo
D10g5QJDIJH6osWVYUWG3W+ZGFcTQypDFshoF+/7SaN7uWkiW8cutGivBLPz1M2m
NtmmAD/Q6Wsrfp52JVBlegH5PteUrLqf4xlzLHRMoPjuaD/0/FixTmc6FBhZdwlJ
FPRJynvtlaOw4TCJD/VpbCmNfsOv571zZ66ndQ2Ng2o=
`protect END_PROTECTED
