`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePsHlD0luiZx0tSbWo2wcuxGpOR6VRiDRfMbEuYHIKpu
eHvENPO9FdV4hP8L1WOzq73t9C4DS4/Zrv30NLKYXllypO6fGblfUzMJ64j3tKlH
XPvl3aXUpEv5EOWFwUtcH9oxY+kANRL311zxZqPzyVG2h1LRXbTThsJtH156FM3G
sphTtRefRp3nxuXUOS84P4Jtm6U0vroShTbtFYix9doph4T7rz8gkIMKe/S9EadW
xJBNzLLjdGYTqL/VVRswVbsBnB9AtXzHWsvv3Yhxj0ttBbDqbfiXCbDaEFyOwBgt
QqMK6LThU2M5+3vlpC6PwpBx2YOGAxrYxhSYLYpBEfUvvV4SU6Pb7KBJlfVzsQ0f
XnxOCu6wl2zpV2m0AOqeJg==
`protect END_PROTECTED
