`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLMu2M3+vBxfkN3ijByml6CyRJV/Y5VD6o4jWqXmBYie
vKAdQaX/5QX2TxgWhvwVme+Hk4ec/CgfiQTm/ba1G7pk/t1JvVJehiliuY78eKBQ
5hAwh7VlkAR6dLyzqxK6bku5q+CPudfI0B72XmrbaE+n0kcsTz0tNmS4o9ARWxrW
cwRTHpFx0I8fApb9ZtMlwDuOXa6dH1uYHIxy/A/edJ0bV5VUdYd9Dw+TwLm3cs3o
`protect END_PROTECTED
