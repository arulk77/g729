`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIRLC3PRu6hxHVO3E4d+ynmMc+6tMG+XHnLrfP6/Umht
zLggnEeUp3yrEnCylzP40P1+604dqmlsuIQLaNvQu+ejz93BlNyT2jiukPS/T1Tl
ATtl9RHBXEiUD4xP4TvHWnV4GTJNJzR+U3FGmLWRyvOVvx5FX8JGCYlHzjuHzMtI
G0/5e+w6Imrugj//woQxHPEwmruedphgQc8niMyvXQWjtfvMn9+skEAaBWpNyN0M
`protect END_PROTECTED
