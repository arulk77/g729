`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
omjSrIRAdLq5UCukYjKnmETLn07+Q9CFjWXa1quOxjLdKO84qgDQU21vZnd/gBnO
B9EFSqx9zh9H4zuhuJdkuIudiDk9M6HWFwaZF7q6acN0mDioosSZV/bz3JZXryd0
nQ3B+Uajt0EMadnnIjcbSMl5kuUbv9y/X1DqdODm3XboW5aN5WcwRj8qX42mQrjQ
uRo7JR4bzHMge9JusY4+tm5y/ZPO6cUunDhz4Rqf+Jpo5CmYuszdiTflwVHokl7u
/JMwpGe+nlLbA1Pi95N/TphKCSzefeRZmqvu/gsTrwo=
`protect END_PROTECTED
