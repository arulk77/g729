`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveALhBzdtVZ2usdtFV7BXJhQ2/sOASqKzxWsrHSE6pP1q
WqqJfPDp6/ugd8zLJVCC1WECI0mDyJxw/oYiifrQQEPLqlzIJ9TaUjf9I2+WFeUC
Cg5GF0U3CldKBj4oYNh8dwisj+EO8Z5HR9RahcaFb9lOj7QjVOTNFL0KHfCGImC8
9/9up09ZvbkOKYohgO/bWph5RZQHaFfCxXco3YJT636anXGMzS7KA8E19Q4L7HQ6
FxOECVjy+7fVg/6TPrtQeGxVLgRZzLiEZXAGKtaVngC3bxuwYM9Kt6T24xNwnRvK
zYC0xHrQLIj/QMMvSvyXfyEvIkNBj0r5GuvNs2f/AeN0UvjbtM01h0KNyPSgcQsY
7z1txAVXmGF3TItauCb9mMEZ9oWoxEDB2/SQ4NLF+etN61y3HB3+i3bwN1/Gf/kI
NHOvqe5RA0pPjvBvqrzauN9BuR/BU0xK+L55DCOX2ugyG/eNsp0i29JwckUs2bB6
jTIttHrYJgXc9/ULBg7eoRUKMIIVnAm9FOWM4e2EA8XCuCtcfwPEl4ih/A5x/MWp
`protect END_PROTECTED
