`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCnOqW6SPUc41BZLuIw0qum55WYKyTqFgkd4clgtmB32
uPf62eLFBCliZdAL4fpgEvjiat12jM7GQExYEN9ldli3rSJWX/NZ08LPPiHqLUL7
b/izbF7AFqDwm/7vLxKIakGkZs6EQdW1ej2BbkhAshUPB38z6v4Ldd+T3Ut/gDkh
KkVQwZkx32HN4chLkkub+tkZuBT16PBKuFEzr0Kz/qHJ7ll/ZAfs3IsrLp8qZokJ
Wkxg53AIlj7+XJNb9Kh7UU36Ry+RSW8+gT0D5OXV8JHvbK4Yx3/uorbsM7TuwOYb
KFTWrtGbr7Obk66GZs8mbdx7bysyjcjQM6YIRVlK0jLtbzwVDvEFVz9L+cEYL9cm
CsjHPk6L2/DKkYeKsSehYad3TX66kWYVGKGbHJw/YrdIvIhPAoFJNy8X0xVpPP8E
E4YvEL9WbMj97mI/1X9VFYkh4ZvygvzRp2Yi6Pc5Hlp1J00oZD1ECrmZc5mjx2dt
qvTcWxVBCcg4if8rAccNpveggNkwrbjCtwboljLYUhtPTD8W1CWKrcxDa1wZFsPF
VKEtUgm2pxAReBEtVNU0QW+n/CGwJ8NIsY0FRqW2mug=
`protect END_PROTECTED
