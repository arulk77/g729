`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOkxf2koReeZbfCb4FiufI34wN9lKW5Gv/g8B6pcnFfJ
CHlyZOB0hcdFE9VDGqvoYKvXwDTAwqcnawKCU821JvFkpzFkniop5aaVwRhTFvU5
5aHs0xEO8RkMveSznaCl4+C3QZWeb9uKmK9eyxKAm4f66ef+e01QlE0W0muYOY0B
Z94qhz/o4FPSdn2z+N21rO6BFVCnhqiFtDcSCXKTumHrxtsLLzpVgXAInPSySRo2
Wpf3hMiXmYtQDqqGNuvZyamiEj0sI87QAi8WPTdmfk4YZoHgVzEma+qas0EFniuD
lzK8SyC1Xx2vKrww/ZxPI0tlIAUPM9F/qaOG+4sbVlyC3TyconE+VXClTB8umkaU
p87E+MV9gFDfhrb8gEs0GY5T27XUKXd8Jwjn+qh8ky0hbLAyW77Nose46oH/np2C
cGLFXlVaZFDnb4jNMwLbhqycmQahemg7qKyGpHcxiDVjPhid6emskYshve6OhPlk
QloZ1PCoDUUkPXRtd1lakpCV4ANifqvRH3Xiv8FfWfFsk0pf4S3gkCionD/wKMk/
hIDdOAKM5LYfbaocwpsL1dRUPQS7VVkdcKBFT5aZ6yya7Xlk/CvNEQUmuKGqnEdj
JedcjW5YDAnUoVfyKzIyOL2GzINk7kHqk9r4IQ8vBUY9zP3tkRzPTX1FWPIrAbFq
uG16GmUsZO26sJVW50fDpeyLGlXJI3LumAguzwg0jacBob3YuHz8y/3RLF2PBG0h
Q658aY8SDPTC26LW58f4DbTIp8yUhuQr83NOHnUpnkp16M01utkG3wD4URCtPo9G
+r+rUoKFSW4rLdcZO5fwm6av35o2krpACTJoBlpFzcsxAVfggqcqdMo8RSBjiSDO
jFTizCm6q35+cOY+SxEPbO4BnqJlIhJ33Cmt8p6W9nPMoJ+etdkGKY5sLMd1E4cx
incEUMxaP92Fmp2Tj82Fzu0+6taXs4K5rJ+Uid7xkaQLMr29Oeq6MTn6iN0WmTBr
ISv4szLfmJ++Q+1YItdcP6t66zRiZ4ISUCB+usKRD0t0FqtExYOpOFwFU1c3BEbL
mjCEdRc0aFEagQ72avavRg==
`protect END_PROTECTED
