`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePa+RIrTyvULVqXazYoR8mtlokaIQLoHsgnkslZU6fhM
w3QV8mGpPpnUAb2JOi2/xEURX/Npn2GHtCmIIvVPGh/DSRJVsWQS/4fo31P7nhM/
MDANPe2zhAB+V3Xv76iUxXh4Wu03T/h/iUOIusMMslI5tJ28lD96xG7jEMkmndTX
SVCSompeS6d3kNfkHXgOJCu1mx0eobwXwxznqQDZU5BqVtQ6W+ULVpsAsH+nXDDK
DNJn5PsgyNT6ZzWUc/0J5R44rgovA/IA5uetIq5zjJ5G/mNzx/sl/uw4TfNTyuy7
0ZRSH1yGkolujXo5HPzH4xiaybgxQBMRY1jF5Vcj26rio4lPxCt9X7nm2FaH+Xxi
PxsXVlh9vt5IRfa00AQ8qKxERItOuKQSvdg8gja8/3h2PVE2N4bY/VxiXxrZxggz
LNM8DLTsUIDEXmf/oKUPv2iUyGX4j2qUKpruQUeVdFSWBNdGxS1OyYYWdM+j46+V
en/g4asJVjks6aTSuMFI6fs0vMr/zk3GgRk4xvrPG90Q/ja9ovJ91tnJhZeXqrHP
`protect END_PROTECTED
