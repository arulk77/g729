`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMMsxOpUbnLVJ4Vf03KPPO3yrVDndJ/0BGxArtNJoZzm
SrWdfJc3jhYkshx0miLu+bdUqIzdrFqnK4YVkxU3hRkMfR1eMSPJrsRzSRli5bk9
I6G7APtsky7tzXmH+arlE7sk9MbLAc+NQrKUvgWSNo9PJVaUxsJNCn81IGMrgPiF
ctZ1h+RUAOi2+NljSzzlmgsF0f1Y4ylVVN/7ZG9syeq0G5YyYLVYyRkKCgvyc/2O
5MF3OxyFUfBCP0fe1XUtjF1BkKeQfabdYca/I5TmETyzKDFWiPVF8aym+2QONDF1
fhv9J5F3c+p40dXBshPq0UKEKMeKx3zej4Lo/Mvnn79cQb6YYb5z3OFAb99oeuch
xG1PCR7V0AFOS5qyq0oHpzAX40gzXYaW64Hg6N2xnWttgvX3uaA06Qq4TqWkygjZ
a8NujDrAVHGnkDk0W0hNzkhgHxQwHf0sjjE2+ATe7DayLYCWz+5+5ONHTXU0C343
H2N00TaaJ5rvwf7YSVX4L0ASjzkwQeJejuqC47ZdbFL7vVuiPEBbTVI6xoAJJwvO
`protect END_PROTECTED
