`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46FRKKuH8OcAP0A1fWdTlbcDNo9kAdvLo2Cf9Dc2RH61
BpI/NuzrxzQHlEfzWqG/AnlnhM7gwxIE9WWV+4DXFm/W842YpgcJdpCaCR3fmQxq
Gx38tiIBngbhnofmj4kVw30TUHFc3VX2c+eO4z7vFzdJWvdLa+7CYyOQFfVzOZEF
GA5hoEVRXoZBPSKNFnAdEfDQAd84iuknc0Z+by/gRrvkpZDjGWRMg3fqCqL4b35z
OIMuNFsN7ThxCf5hC1AWxtCvbxAVE+iUrJdYS8Eao3jpNjO1AlhUXlWHza3i+a2J
eqkuuLQbS2EDNxcAVpJg6biX+SJbc1KAtCnSVUcqQULjZnVDUK8Yg3/NHW5yuJx4
W1Fhbm2xXcGgCokvQ+SJ+w==
`protect END_PROTECTED
