`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C0LBhMcx0aPI28a1iUmSkY443Gk5yltG/6L7awVWtzFF
As15RD48XZHirWMsDeRndSGjXhPEShUfc1SPUPMXQ7DvszE6XfW1cu97pqnNqal/
EwLjQ/GI740GlnAd5OYwnh5p+TdRe827fivJ7D6U1YNMUX9ul2enYZ4FM9RPiIL4
RDgVBw2ug9fBHbuqeefRLvA/kL7iZ86HJt/CqF5AG3+4Z7U49Vw1OzjECqfxxOfv
HEbG+rzkc5lHCPZgOzXpr2EfWGKu/emzm01To+UQU/z/TIXCMbHlxZm/m5EDJOoz
Ea5CegPwXKVZht0gZC1pN5uB3HQ/BDi5IbQ86DWybaXH8oNbFUU3eySzgnDHDtF/
8BXmbvA3lHLr+58ifycDHgBpdiXNVNxJUlCxJrTDFpgtEO+8rf8sfCu/zeiYCVpD
y/CCRz3AsZQxA5LHgwVtHQf4u/AtQDxjGyw0wYtVew1rq5/xB7VUuqFTpGTQD0+j
iFlYp9sQfVOhzmrLU3rDDvQdN1c2gTLqLykSLs8J+2iP2kE/hRrH8rHuKph/tCup
avSBhlqBhl0Vdna4UTooWuxAe0nS087xqiWKMioR15NAjX90KQACGToCaAXMiu/B
s8j9kVkxZeB6ZAOrDjU9gAOIzMIm84tePbOPOtD3RU4/wkQuR0qpsMQLPph2OA6T
TWs4fCV5QBJEzNkbj2djn9yDdPeAyCv/pXTJIher/8vFbGSw3lCMWdZhLWYxe1y/
`protect END_PROTECTED
