`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCoYgGxFaQnLNK2rCrzL+jqFca7ITOYB1djmXsUFID8z
iTtrUn//2vjg5Ct3EXlIVsrxLDHS2P7IVGqkk+C/Y4X5i80TI1s9BaZSMSrGr+5C
PIv/+OsDXZ0xiGerj2JuL5MPN/3X8mFp5h+8EbEqyNe0sClR8+XycP9rzaNbNoCE
XdLCnwkHFFXxDgfxVhIlV7rMTs2FnxIcN9J2ICRCPaR6TdxB2aJwTvOVjJ/ePmIA
DVm29KQnVsIkV+DWz3EUFi7rmIF/wCPu5ROuuAEYJugROqsgRi3aJ8a94h90h8U9
SecsmG4p8CQhBVKG2LGA0g==
`protect END_PROTECTED
