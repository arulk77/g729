`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAbMDYGBQDj3SsWHEHUZZaTVp7/r99yNFIuy6WCMUNRE0
KlcdOefn8cVNriWMK3G1ftkGQUXLW2oMGzZ0A9oKcA2evhx+2mM7zJwsO1OEUHBP
OXYEpZ82qE0ZxeucwfjToVdnwH3pYWIDdTNOtOYMYlW7U0/TuZVy5BaTqxAx+PB+
HXT83FNgzNv/QYLT6j/FrUDCrOs3srazLV775AW8SB8qE/CUHLTAhcYBI2vwPrB+
/TSegcHljXyuexmLSAAK72yGhQZoWehHRhDqhbMszMN9PN6UFXu8Z5HVYAA+ahjX
UFcMR0h7spWNAmC6EVRKJ2Hqzyn/0lu4+3sQEg+wqX5qQ463CdC+cmzzOw9PhLOI
wa4Gg73YKFYU03j1bXg04ve+bBGpKhyhkwqqzZ+s+WdMPRVuZHFJM++y/rIWG175
qh/jbovJvpbza6zHOM9XNIPt95rS/rkIM90AatVyFeW+/2+yV7kyPIv+Nz9o+OLm
hMNaWApWF59O0Nf2y9wWhnpme93bBtinqMM0jH+qvshds3vnWvIdaCTXRnBycQXF
Cq9W7TB4yhFjgP9vozsJHdRmkqjG5kbAbX+0kA1JIF1TNxcj7f6+o0QP47qTT3zZ
jnUvbvM3KEXP+2SLbac+I/D4wFmV2KBT/FrFi1/Aljd7dnE4Vggvw6GE9rLKELBz
v64L8+tOf8Ju3N4E3WCCtAOPASA0mHh8uSYwKpihOWaI021A8mPD913rxpn0fkGN
rmqdTbIslOBH8uNc5/Pl9OhTTosoCzi8B2qp5Punu5EKYA/YVMbKNyzOKjEQs4fc
xq3aw519uvabgIuZN4q3X7Igwd/iToiewyVMjzYmDCgJnPGJLK17f7hcS25JVMeL
/4DKnRxnVVJZMbs4uNep00/3cIgs/i6sGwo/OOEWyjcmGvWN/XfXuk0FVK1HteFv
46BnMMLjgKq2IgM99xCZmdu9XxHGpG12UljU6ZncnobkNUKoprTM37+y5V0er4Yp
5KbVl5r0KYLSCGqASn1Gy1F1QMktOSroRCqEm4w0ly4LNzY/c+Tq22l/5E7KPMIx
wmi520bfmeBE5ddkbmtuvoeRFv/RbT66qsMjmgqQXNjRSg87q3BFMblpw3a/JSZj
s1A5eGo3i8OlVANiHt2LqKt3WbDbAeph7A9hV3ju9+LT6AKgjzv+y8eDraOkrLHM
ar0fCDLEAeKPHuZsngXco24HqgVOGbOfp4bh4OriFVv+tqSRvG8AtSp70NEqbjbN
0XhyR/Wo/5Vythwyg9CuKJwlq9yKtPoBf5HPk8pkabZhyGC96zmZ80LUSYk9qvtv
F3Jugl5q30pmMTg0UhGCXvkLBKX+1I6obRWwh7aKOJWNd6DPILzWVmt355hyXGbO
2yRQEpJuSX6CRqj8f46ZcKn5OwrCzJRBwqm7N4L9c69DqDZbuMAsdVX3MvbipFOy
BREVeNecMd54rxNszUhgU6oszcPrzbhAzGWFCt8lRt94LWIEJysa6uMTyQG7f2na
znFmTX22gpzNE4nXMj7Vu+rLHUodhYC8v5tpm3HoQTsoGH+iJUUXzGmbOm+zUzKv
bG6Su468KCe6edW/tmUtZNok8tIAC79Lzc/jaqZb26yWrcCn91AzdoG3xRPPmYmU
dNFFKRnEa9GuIYHu/gCQxauyLDexBqR4Psic1wwhkweC6z+cGvgWtTzEqvK6TcK3
Yd+6sBakukaqqxruAPXOzOTfMbSMEy7BtNwdhL1B2Ufo42l0pHJkWn8RzRwgGAec
oeZlm1w6H9yuyIlp3npfdswJyjtmBdEvzVgEFR7W29sBuJS6suioGt41GV0IMdUa
lPhD1bgp81IvPm554H6K/zHMkO37CFPsm1ESA1IicHTMPLGnwLI9rCxeE66QObsK
apicKMRR3iLgPGqQiLTrHGQrvmQwWMxRSYEMHG6LUwkDV+8EeU05h3zjvg8JaCiD
0XAqY2nkRoXrgYAHEx8ZrBCHPFYTkLu6P7awaxhUnEpaAT13zyexDo4xTGNrxBLi
cbbeiqu5Hqh/hql/+WNu5DLg17rCCrG+pVZr89Ow7ZFKsNRBmRhc3dkoC0OQzJOQ
qKf3zXuf8Pwc/Ta80D6Xi1U6nnEk1TfbtVkGwAvuF0qmhFEVWiDzJpQgNN0Kdkse
4BqAEOdsjWnnRpmaPnwMD0+yWYPLUc7JHxyMx+UyR2NZlTjD9FpNx4G9vuob07ew
a8nY5u+uw9MlePxdY4WfVwzG3nGFVuMMBwpqecAs9sM/kEFxmK3qVLLKqNr76174
3ZMeMFnhsZIpkAPk05vOEYTalkbnxe7KjnUm7Dqya77ZlA1HAUThqbKvs/Wmlinq
KoxS626XV78JDbfX++iSfxByyliZh45YPV1zS135MwsmyrjU2B/hq/x98GYmqNEA
9wv+gtE8+f4v8QwsGWUazayXHcswoqyRHGv/uhTQO/VxyQ/q77J1ZFlHpF1itTMz
D3kT3TC9WdloiXHllrVThezEd7bNCw/+fyGTeqXBx38AXth9dAHmhTvPxkTm25V3
zRNDQZrjx59znoJCMT1F6WT8Qd3biWnlsfaPbPSr0Q6D0zeSA2zUl2IEX86zb3Dl
18vxclmGoyf8eFGA8xTEpEMJQdgd7ErqykWj6jYQBeXIec1GDoyIu5ILfqL+WtaU
ooH5trGgC0YlnbYvPSseohrPX5X1yDtVi2Lrt4MdG8iPiiMnhr4i9rn8lzcCsAus
DoJgxw05r/R0t9NNm4DFXaBhb5oKziaWlnvDBy4y1hqLLSNwLoaC0DPVYtqcGzFt
2dMk/NC4kkkuMvMXvwADJXfsAFEHYk84kuqdImaP1NPGnvtsXEdS3bsdOrj9Nwqi
Z0TRHOOBCkWqUfF+xx6fJkqqofOGoBr26vtfQPeEnVqNaNfJktxCDbBHr1BKoHSh
NWyg5QI4rq0+nkOKhMpEhnCqv23wMROa4LzhlyRqvtnvf5hwjVXWRcfAbFISrx2t
Waibss5gacS8j8IsdjyWdwF79RgcdKLo/iGjNUQa85a+MfNeTsoJCZPm7oYd6suF
fLsCZFhSC+i1CIe7solAu6N0jeBp/tbA1WbXCaXitn6YQkbmUD1krBhqavXc+L7b
iIvBhPmDweKmuKZDrZ/0/H2QMkdvl/9DDx9g3dsN85SJ68jl7OUpijdqEX0DwPI2
w1bOhc9OBmcea0bce49ELwDRwxb2P1MtxW6auEQyxt5P6jWzAd9S0IT3Hd36kTBu
M7GewuVk0ONWujW4MvGf36mY+QKi5fvmn7/CB6xsMdHZb2Kao+w7aAUHDucZkh3V
RXJMYznHtEWEAqzums5fSSXNrByJreMT1vK+/ISk+hjNRDLnfpLRtfI1+6/j8C4E
cEiNrwTt8ctvObg0f0v1WaVoXlnFjWkWE96WNwLe4cI8GLpQIBTCwx2LTytK2nQm
Hfiy9ZS4Wc7uQh/7D7UW9jkHOQXf0tRmklrxM7QLRun4pHfDyijlcIg4MarmkLkr
Wgmk0LbVeWMx+04+FwhPxP+zzgUFx36jt0V6DLAFtHeM6ltFEwb3froUK5tIIA7Y
bE9jG87hcPbIWeLHP8Sx6S3kS9KxQ3mIRP/CX3dM3WT1e5RNI79842fBV/hYYaO+
Nd0CN/eY8CXM0YCNNwSTv8/fq9TbJhGahYKkrwb+ZpSZyW9qAaflme5mtNRXBwuZ
HBaGKeOO7X5KqNTVJzd7xXOsyIGJgTZ5xDmMnqRK/cj8YH2hqlqTvH358wzx3h8u
4kswuaOeL1aoupsXIL6YAOtjpeToWnzVb7EBDw9Fjy8MsOJZqq+gqAbj1H2E6/b9
rQljavQXwetSzc5P1kE7KeKj2392IujsohfHA81bOHrxmoXKkWODvAZS2EFqfbky
5I8iD+UVpQ9RE7CoWrJacdbPyjwHyn3MIqcvDE74sAk0PGt6dCNE6j0+QgRK+Ekw
4QFu6FmOGcOpn6pSRiIKFdz5FHwi9Bb5cYwad5AsyLVGNJZ5OcCCnC0G8tjhfVBy
EJlovmMRg/0cyWAjW8JZ6pgl6w4CFtmbOFDmIs8eLbyAEl1/YUfGx0ufzHtyCgTj
4l6Eczc9yoldN3J5fmipSjmH5vf7lBp0v9VCxpzLsSNwa4qnQvpC+qTqn+fmASwW
W6zBqY7tOwz5w5HdkLz6whktLyu3VMZj7L0XDMoXuj4AkUjVVmFG+XEX4GpDmDb9
wM3D+XlXtKSRlz8XX7yM+eKpEuTGwRAYcJBcWGxdpgSFi4FAKUoXLnLs6Cgigwzh
1ES7CAYxc1Z5OwoQVNydJF7rY7B8g5EOsILumI9x6lgUMMPloGWmFvOzM48ywKQs
TjJTGfv3mEnT9zTsiCpJVwUSxDPVoLq67eXOkAZheODUfp4DkhI0spd8xn94I6Jo
kfHPQV8eqO6k0C1AsmacGSAmxOOtPrzY7frGTda5iXo48jSihQ9lPRbXrnn/Ashu
Ct1or2n1MxpLw9kd/EzdC50jEwMDf4Ig9AE9Hs8tNeWjPybHtzoUApEdZZpDQiqR
shAjmFh5inSzRpb+2GiCUQopLgmu1o4RPsxsIJ2r2lJ4UERUcQmbJCMp9tJdwv0p
4/kN5A/HQkmNKKkmn7JJ6zTnYLI5tzkmkrE7lh7XUm6tz9aZmDEDLOUARAYy9+7c
CSDpZeIqjSsQEPtJjaQZPt1s9eV4cspoXROxw8TNv2eOOaPumF4533uuteNen/J9
o7qeW/CTS7v9QG46l+yr5GQ86MOyUnz3dwTcgVSZE1Sm3T5qL9tQIIivvxJS6vrg
BB+9KmThsYO7ZSAQg60/Qywv+oBu80CtBjqhqp90tE6frTNJmbhBz+QkHsuiqd9m
SsS32pU6CyB8ILEL52+yhbJpAMGrCwA/pxheqeVUY4G53CcMd3vsJ3/7G/FZ6AFy
rhdOpwoEQDDJeGEsRs0qCIegigW5yJCZBs3pcsX3lsqDgsF7cbKDIJVVyIwHRKy8
wvZjRsKOYu5U42unO6hBmCMXw79cVmKMqcyLN6QJGjdEIlfZ16skWi8WSI//BX0P
uIwgK4TE0b9nwJKPgRXVWLBuuZll1yR20UWOXx0Vy/P9mfLv9hn+CcYAWrhg9xNT
Zus6y6jY1ZrjClRoNmGs9rSDM/C7hfXkJJ53dTV/G2rBBv5qmplmJEeMkXUeQnNa
K0OXOXkmB+3gF1POIN0nSMTRRWkyEc2R3hD0GeG5AJIL1yFMaG0Lq1NvQ+xfsZoS
xhTcAwcid2aKTzXw0uxXp0nZopCNCVEsG+7RWoPg1cjd0UuNQLj1jTnt00OboFls
f85xm32jNQQ7H6XKF44+CPgIKX5xZfFMLol+K6AmlW9jlLien75B5OYTb46zEUJu
SRqGHvoiOWxoU4B/uTAPhq6f91PHDykrWxOBpjxMeMUB7GIIBnZApK/RErZgluC8
7Hp1d3n/wY4h1QaYhkDumDGhBmNhnHviuZOQPnN/capjSj9WJEyZ3lYIXYNLCD2B
rijYZJktznUi5+WbTvDzMNkDZIyPzjoZhkLtBNOuhgFLfsaUc483cRIdbnDdr2Uc
XnAGY7W192TwXEnh1XcnNcWxFQkX6whE8JW4M4WzznLSbGuONXCuybctHb5uIkbE
PVI+YzGZA4UMImBLF04s3Xmq+tR7otJBRo1VuGN+YHdthJMM3y3PxxJaVzV3pQ0f
LV2pqBpwHjcfnBUEnitgh8AMnVkue/j7YahP+q4FngTCpW/mJPx4aF/FJ9U48yg7
sNq9wFOQInQVUArmE4+oBuVBO8guY3xIJWug8Cii9DyK2I2S+VkqYo2tvV1HD2Em
niNyz66w2bVZAJ4qW6QLc+0cRYEVaW+hpRjS1kDjdnMxILiTYiuzpNjoscu36MhM
tUSziDU9JTQNdQMseUFvEk9ziSCIRmYxfScIlDYig0pgW28AGAcISLJ3SPEtOPUq
XxZFwF1B+UBPf+zCWy+iqzSn0r6PtITl73ukUo6C17bFhG9D10E++tWo0rnaQ0lt
Bj3uaXpiO86sOvs+rg1/SHGmlvCT+DnMdxcc2IP4tXiWNsKQgsmKLLhK+BsxLjDz
/Fd4IcBE1EUCdxO3Lsji9mP/D0l5FU6f/eg4lL4drc3z2W2ZO5WlVQQOqkfOvQwI
nQs3jzpQXHg6NhdMAS3AqoQOfeK0aceq58cCDbbUmc+t9uRNUXcxYD3fg8K80mXY
Cl5Z2RaUMhJh23H5CXz1PqHdThTZpHlG2vG7SH1n4ID5t2eMKR+eA5D1THExJGcy
Ut2KIXrAEDHM3eLRQZOAYSJz3KBhOqLrpRmg0/6Kpmx4F7FxkT+5/Rk0aD5LbK/f
aiYqtO9WHUB/huqUllhGvjlU4OhZZa+u5BWCGlw37kXdgQDBetgrHZ828r0QCALB
+3VeGPAEI2uyECMpEQOFDvrE6RGXknKBHUc9lTIlwAkEX63AAVuZjm1iQ4hhSadW
DEkcDpnu+yKDvXVcLtZGaN9YRZJL8m8a7jvYk9EP7pVQpFBm69wgTApDTMksGE2z
EziAsJWHtrOAmBFR7+2dsFEe6GKvvuUGyRUXCFC78ossOfU7cRFJ+qQjumwHGOxS
gEuBWZYZeSp0TJ9V4QOhqv4JS+3uG1UZG5z/3mCuuCGvTMUtR4p/w2F6U9yD0jBS
YEjha82MxJv3G7NC6DA8e24ITvUlQJbYZvhrLF+EV0I36bDFKTum7lZQyflsktSr
+ScSx29Y+A4sXMxrfEl8LITgSrT+P3ulZC4lYJ8Jq1p4I1GoN1Z4s4s03aqZB+mm
I21U13WwCtiwrQUsyZCoNSUvr0gWSiy4ZGyKzfLxg/dPJM95jn+zZnem+WHTdWzZ
CYf1HVT3DBHN71/NUwWdLCRYDc3NjHzCH4A2M8rRVce5/s7L9DFBwA40CJGGAd9U
6q5Td/6V5qc5L5Sp39U4oEafpAJrKN4wWo2U8xr7gpFmVdX8DnN8klpH1Astg5KU
x03O6ilDYr1/AW8psFUQdnl8O2jPkGrnVWXg/C7tRvsjYF4dcS+pkrvTB1jhEGEp
VrDufyacDued8O7/SYXGbrpzFS/rg3Ei7tIew9u1E9qxZSV4TqBEO6jd5FeTUE/z
UwUFXgHgoKVmkXyXWssRoUhwEm7QmSWbOxJ0YomyCdBUvN+ipsScRq4lvL91iZwR
jvNo0l30XlIJx7dkHcNLnuZPySuuoktSLlRsbCLk7MK8LfmLZTu8/+nJly7un3R2
K0o3DkdoiOlDXe3rD+45BvWODa+AoE4/Vb2GAZetqT2Uy1wBp0Kra2yxnprm4edQ
1BzJAl+JvTKJ5JvyLnqPmKyyLaz8O6XTo4dR2erP7lNzMeckuVkQiPXPd8pBFQIN
yub+q4FnxHl4eHNEApL+9qLEXr4/QXbbog6+EyhKCQU/hvRY/ZZPom8UvT3IlmYd
uU/uDJUEr4FzWWLUIzZ9O5Qdfxfg6zkG/Hrf/GeLW+jWg3lheZWOVNLRuZwMFmk4
yOI5QTS5AxT0CEIEMlkv6IdmSGYxJDfU5wfwNmYGxjnqSqmuKJKz2vVJppkvch+0
zw9Yyqsngxz5KhSlrwRoFWTyvoylMnb+XfFqeyq61takkiG4wXWpU56xfkF/3jkY
fGxymr/Ps2QifhwkIA1WJRTsYAeQOIBXu096tsHBHI89oJLbWCsVKE0JoIBM5pX/
bRwLufpa6rGuiK6XuNfWsWLX6WraLwdn5MJv813zO1ATOx1r8N/foBYLtxbo+G5W
FZyUxQuQWfQWoT9o/K3cQDQNAcRt/ZtRH6lLpm6K5qiqEd0Bli9HEQkorWnFmbnp
ofGNAytK0lxd8IP4pw/GyIx7ubMAeG3nBx9HwtAMMed+uhyriExYlvlqqbOq1JbH
qDxtNuTIp1zmhmQeqB9tgZVE+REppI845RPx3tR08h7oiGYKnfEtV85ZPv/RZM9z
HjUM6HlkrKUXMhoqDxMQaq1ZaZ992CTno0GmIrXAsQ9SFvsSNYeNc9CV9nnkXyOv
W7s4PyZqK6K0VgEVhDeCw2RInsHDrP/QPl0dndNTQllyV5L6+t+UlzcTaJ95mz/l
U6qPTsRBG0mLD7daDCdWqXqNYxmJmXJKMt6hPr2HDEg2XMFLPN+BmNTNmp2v81Fu
0tKuCOjje37VFr8uWwyXXNakKDBxkTCP38DBhk7mr0BAcl4qqSNWdwVGsXqX7TPv
1FEspFOKD+Q61OgFOnJ4RtEOgEu6Rc57+cQWznR1uNcBK49k4R61Jo75rTnhIYK3
KEJJ+sTwXb31mergo6AYyKoB2zFAps78WoFUlpN5mYfxSIuyPJ8MzdK8VXydbDBF
JP8yrZByuUfWkvaTc4C8iziz8si6tJ95gNeNP5rQxmr2RVP8jGiWLV5880fREw3F
ObAu17PRK/DTZPuZyQ2ipDl9u3oKtCjrH0tJxihUzcL+plZ4APF3pQL9xDVdatF7
F/4ZuQfhYD3QxZ8mg6SdbZ4k/VSfQorx+6S/ibb8nrBX3XonLfMI/l9WB8Z+DjJ1
tGL23RHgsRcQKh/MoGeS6Qvkfosz9QqGTWbOjcVN/PIbWjVrThUNjJbWj3DqgdzO
SRkwxC/OwEYOkHGbRFk87wLLZwyNowi/++A6LMwCAzF7Dqe8zM0AciwIRi2PQNQj
S6nGMScBKBPdg+Dw3QVy9ZFYEjf2jMtS4EY5+zFPQR3t5jrlEHo8C07c/F4IKZLz
ysvAtHK56iChG3lsAXS8g/OFkGNW6qPkBiUMbevQoFbO9suSroyy0nbl/hdNd5dA
ET9xldFMEd2ikpxpjhDb9IYs8HZYB9AI+mvYfdIdZNRgwpR7/0kDzCmF9zj9Jwjq
VlPfYoHya8OxSuMCN2h9TMlc4+Tf7WGxL34BTsRIvCwkgCn+yMe1vwxVirCkQ62M
szmV7K4+fgNBxoM3IP7Sqcue7gDyGJvursBRTlxB4UqseTSKoLQRYFMEEhNdaUbw
dA8UonnJzOkppABcAm2AZ4QIS8L1wOffpYbSvBzM53fV9ftzyBZYdRTDMjlTyR/p
3gvYTpO5iY+BE/gKTkvJFjoOlOK4cXlKDJ1bUZ8jFHN9VWuF5Ai8QFHx/zvpP5D2
ttmZe/n7DVqqiHmdyHJmxIKUFjo6JxMtL5x208whhkwKoo9P2PtNAO77PDg8UBg9
axHi/c0TpSwoHH6DGWuEiKe/bEWPiP50W1zPgwWtatGaOjDUGdpCCloy7zRiMTHR
lWvC8PYnVbRabHn/KTPhYAUJ0c4Ga/XSwXdqwcJ9o5mVu1Be9SfUf28rM3m3m8xH
vxDhffj5E3V55EOSAlXz7Pmk87gny3MX3X1dh82U1m3XVzqOvo/DmcXZzkNRt3B3
/9eze9xDj39klxzfujnxeojVTdg2vtD7KFu4YkixFbDdIZsC0PpQepLfEEe2wvOf
S7IEsLRtv7Hk4laTEWYEvXO5ou/RBhC4Qd8Fi4lddFm95AFpyH1ojIaQuvZwdaXY
el6ci1ynN/kVR8ZsbuUKI/Fd1XZn7pk+OL6weP2pvOx8VdASDBG/fazNHgcOVauD
B6EpWy/ZaU1NtK6bnPtab9f2HJbBweCxjYL7LGZnmtFeN2l4Dqcu9LEVxWdve8/6
bKfrz2nXkvfxdUDNUU8R+hmfIdjApMUm283168PmblFRanE2KbVHwXv22huJuOiJ
+/8UHMIZHP59mqZ9DLbHX4zYol2a8u86QYi1gd3ch4XAEyLXtAkx2ku5GbGJHWOu
bh1JKYAx3VvRoNS+5bscHEZSgZbaTaFWUMldWex/z5c7YjtdoiGTMVhaqAKAkgLz
lgSXaNXuSQdtDORZJRcZMIFEiGTVyIVIubBN4UW4ujhKlw0zksGaREGo8eXkqNY1
Nt4unnpKCPwxUeGwOS2g64IlFZKYAEm6ytSSHeg/zWd0iDyqNDNyM179tftlpGk6
2iEJXPKdjUrW492ay7quNHuyoPN+D2vs7dZnEuuNCjIVsBhnmHYG16U76RY14e2t
06QH060a6nZYpFJgLSxuA50MGmNc0t6tTSY5KLajxMQNjhDcrditJfsxk1fC/tzV
UEgx61IUUE04zrcBogKmQVWebElMWAxgy+wRvEPAcICR0E9h4j099ag6e6Evl+Nl
UL6/MYpfzKctkJQ88KYixjo87LjHGqJlT6gtigfXu6XE9tnBsyfg4QPj4qFTtvBT
Gs+KeNqubbnJe+TaaeAARyk/mslf5OC3nv38por72+uH1Egy6OEEfPuXz5RJlMcx
aXE5NRCN+UV2KLySEPz+kjTFO61btDlDpGFIIpNc7tkPAiqKcJCrNlhhDy62OWNe
mi8pf30/f+j2o5wijZ8xOYSU9bXebkcuIB+yUSVV14DsbMQY1mR9skkKj02Ul3bl
UAZDzeYVY7j5B+WBG14RE7zmgG0crqgL+rqQG7PQRRpuptkxz+Wiemeocp1I12GP
XzuAhzXJB9q6ERR6L59R/4h8Lm/UnstsoSIvPggA0rK3g2c+gQmXaEgxK2R9Q+qq
rdR0v+zBmgZIhPceQUCu5Q22C3AjKSCEkb2QYZHCuB1FAnLyMzn5/x8LOGwvD+lg
QbrNBFsEEKjNmS8pcpTM6UwzJ8qB+GjJ7sSWfL7qji0NRV1KT/VVeU2MXAJujal3
2Oh/wxaOEhdeLxbqIg42sCnbs5a8kRip0RNEw12DsaQU0JbApekt/enjLe/aDnYn
ppZm4qSDMYPTLELxMAR8invl30At8wOZ9n8PnUShk39rBYEKfQt0kwJug+JmBbT5
kA70UNTkCNzoGTRN0vqe28vdmG1ILBPerfP8IewGIc1VyqOPkVW4FcrdVWBcA8L/
fyPM+nfDkoYPMO2holGCdqJwUraNNkaw/ckfILJ2SUQ1qRsCRASBKgV75rwSKHtI
mSsEYKg1U+wQ/YCR8xpMm0a6uEZdtT8VK7RvrSOo6henBQwDrFB534oF6se/Tfl7
gqhk17R5HzOYWOD/ragJ6unRhQWq6kmrzXI2bTcrcjme1dSp0zvoootsl1VqB1K6
HQ7nePyGrXYXEIvVV5VruAEIA6TAfRJUVUUJBd5POF1ktr9dcsz/hv4uteskqD0j
jqD/6C8y3WBIqQy3/mlp1kJ11aWGF2Si9PYdACx9/QMXEYV9MhbxN6n4/Yq1gspq
uWEJZOGuOr2/Fc7PRtMxXfUv1/o6wg4b5b1aGkVEpfX5e7Z9PyRuwEGjRuTI/6UA
pAncVFIikaRaBh6f8bP/L6gDss1qItFZj66xeJOPy0YS4GxGteJsdt9iZZzl/Lxf
DZprT77OqBjhk5T9YMcNvNkZkNgpQqTVIjD6qzn6HD92Gi0aiWb4CJBZ+cVrQlZq
bcwoZ3sOOqoNFbK00VZ95ZoOlWgze+HR8peM00JI37R9l93HdvBkKR9eXy0FMkJY
YsUSD90C+xW7O3ZBvftpK1VeTaOG+BKj+2RkDNCeYGU9dIPGKRqAixvVFHdzqJGQ
OR8p4cWfwGJz4yEQEOn0Mc8bWRynH53n9f+raURRH3eCMGPsGll3dfnPJqCDt+Uo
jJBtle3+rmMjsYonDpulClDT+26SxI9Pq7fa62bcUyNzfH95MROvqIaKUWvxlxFl
aTTi0y0Nj/xZ1sZeup+PWMQFOrC9YBMCGet9cH9bBPFFcYRjtwX/Hy+EL3SpaCAI
wiwz1ZUToWD3jVZ8bEajZ/eiZSAfGCtaeaztRxQcX6gyt8HI5A4tm9l9OHDOJY8G
zgSUlFFIyLjAMQAEAN2nhfsZ+jHkpdi9czBywWjelLYNL+tosQLWqeFFqu6Ot5vJ
k2E1v6+9ObTR65WWvCzWkT52gzxd8Vp4v6y392OPAeH07KcFJmQ9ldAka6KZJJtj
JI3omSnL4gYRemzrY9t4bHdVrjzykjGAsyL1GrpumrIDUaEARgtQ0XkWeaB2t7+0
VMe6iD3SZyocjWfMCCxzVEbTTa6CgZwpMpJL/T3AGja1NxIkJNvPHSZbpbhplWLi
Og1Q86vnUoizQqbGO7Zq+nm3hrCB4yXfYf0V1LU/vC15jH150lVbJbFDXCfOGBAp
6UAmjGKfdmVf5KKOQXdTNWqticuPmQXlbQj/hbBMPDWSIWqJ/xj9k2ON6DMh9+El
sHNqr75imHxIPHTCICZyESblobz0571F/hNoRo5duTCSwoS6MX7yQiM3ijfpN9mv
2NoQXM5hXXhjam5iT1etzwywVMi8trn7B7aUMetmmgkdkoYVOOVMDZu14Qc7ZqbU
fty8ZupVyvu9lDf5Guuy/H8DV4V008qRiiuHmqdVyLXGqwzAn7G8NOsTtwr7k+AY
ieJ6EVGyIfLF0rdBb02Uh0NhfsDxUZnVzZ8mDl2xfZ45SKX+Bept0qcFVq1JbwFe
7rtWkD13C0mhR1YMcu/jPl/tjwGR62JSW9NSpA3jdHlhM8Y79r1YVTvDtGdWcp7/
q8ggMPYgEwyfBz7fvRNUbLXQGSj8E6YmTgJvRfET+xgETm05x3/+l39OrjO3izRi
1ogi2BwmyBDQgaxRGdx3oPfOHBo1T/pnwuGjpCgazK4CIHOdvcfkCPECGxGr4rFW
n0qah6UOAjIxsprbbLgsKohHpEvBshE1egLWDHMlEMIof52WdjOCM5T55jo05yBc
wi/4wEGsIa0EmsmFu30ilQ5YT+N65r6ldecelY/r+JGwnoeG4GwXoFGqEP93MPTH
hMdBnjc4N5mZaN3NIIogLNORuIhAFZY2u4DZ41B/8TSYHZrwOKTaBSU4gadm9r8w
sP1lQqnOpLNhRoj+ASShTqasRdMIS3Lbf4vcAnRPOm/aIYRxFgneLZpNEAXXN/CT
5WpWKtWcSwS4LKeqftCkx9Go81JX9oIpG/XNoWXVJxw89+dbLzd7wMf+JaMtE7Mc
dbxFYeNyY1QKg3OtjsBUoMkBtaEUYp4ImCqMfLvio5nrQ+/P207+3vDv02QZxmu1
hsf2PtHF1/6sk9atECFDHtFvPMmYtA+A/JeTG6olbNNyiN3Llk/0i/Z7qN18pmk3
KtklkaR6vLXdjltKJOEMx43dHqpnfJi+ubKyy5jmJYtDjxzYrkJELLxuGiguHEB1
WelAP6Si54pjU0LR27dZEkQvYj+8dUu+RxJJ3RB7BslOci4+38a9OruiIQrU/3gD
ETJOSAI9cYgQgwTBWjRn1H8hI5bcKOic1erzxAFVaj2IvBRceIKgzGFe5WBRazl/
8+KNFuWOdLEI8M+VmByBOCCmQvJOBp2vpF+cTxRHyNH0ftdVmjZdB/6WcuFmHarD
PPGa/itx9aFSnHQqyDtorC3NOg03sbxIg/nuFyNZao8W+ZO006af/bY75Pbc0d7D
XiYUTZ8uk0JcWYVV7xXUKckTOePC32jjK05Fyh312a10JiE0Ib909SesaDdV6E5L
XUOj4r6E4GHKdCr8Bf1g7spDbE8oDwfH2+L9sNeN3X0JXukO22fQWzNv+Q0q6+vT
v8dT1xw5H1qshRgyLams28yVnBW4SFe3zlSyzmYY8MweI06hLpYU+GeSHROOJC4U
Cg4aIp4e5+U+np4MucWeLGJ6FnJPdAqEFgwWJ1HvzGQRLFTtxl5P1Io3BxLxj9Bb
uUhJabpOROxzUiQndBWMftJr5+h4ft0Px1YwRWBnspI6MjMEImDj9iCxCSCTH7cw
ZNJ7OkRKRCXi81KBakWj1wmI/nKb572uTIG9lQ93QmEKqQqHfoBZbCDZum5TIYdJ
VrE2+s+LoTtRZFG+IQvTkm/wYH3BilDmnC+6DrSE6/nUeSukbBT8XuuozSFbimxa
xdyR0YzpopvrES5Fm/5+QDhkUWruR0pchzDkQ122WT6XoA0+9GwyvY3T5mcP+b3N
dtKDF8bQbY91qW+tdvv4CkC6l0lKvG/xhNPGdW3zdi/wq9UN8J0+FFS4CUlz9i/i
EKWZmeW3gMudiSBMszVA1d+MG13BuA4Mx82S2TrNG73IH4jgPP2NDoLhuI8JX0SY
JCYJtQ7cYtENfrT3NJ+OLFuC+C3YcGRZJ6Bg4KvUBLeIFH5SczYnDAv6WXVUXkB9
EbmTnPKT+ZWe2TQKruA5NuR8/wJzQ+4tL+GidY/SrbnBka+suK+RMMgDHJcHHEiK
TUyRfWYShDoFk1Sq3kgOIxPHqsSVm01OGFUfGhWZ5+s4pbRnI1/lpf457vngxKp5
bY7Ra6whLLGBULard8Zq9CpJgDn7VxaJmGfpoaU3Wg8qzdT5WzMih/u+7AvsqfOT
gyqZP6ifTBXWiD4bvBKGcwZyLQ6Ms/hPESEOCDfySUlw5LqXRmZYym831yJ2Yw67
FxQOncfrLUnmO0I1crnRuyjm2N1krvmz1jsC5OioW/4GhVF9EbemWKllS49GUI/b
5EuGN+xxoQ0WK/JHWxUsVaSPYa/21FIzxmsaoT5G6u0lZPH9INrAD1BFbeyv4svQ
ZJigtOPw6HJ0JTZcQRSPMvpJNSTIecTlZs/zT1W4siT6at9yLdPPGIsSFLfn+k66
OeoHwWq+QPt9HV7A341txOlMtRVM4v6TIIzjVQUjIOwSFVaBPVvoM9u3eKd1lfUd
FIONQtQvv1GTndAjzMvZzKmvCR/bpL9Uqu2rK0+514A5gbrldlGNwQ5NSttmwdZg
P4FIaq7MmiM/Im7TpEYqlpc7Ow/Pxln/VulcHKagz+4wXzQvmE03Y5URG+svncOj
9erw1eQqfAQO5dDohUWMgN+jhIaWT1DsBeFWUZycRMEdnOgNDTKPmUdlCAQt77Yi
tnBMSo6XOjf3fBnz14lUDSw9gUvxHG2VO7u1kBZ2nhcoMfaZjr+w2lLXS/NeK4KS
hMC7lGsD0v9SIsbgLtC4Wjw7JFrCiKPTz2prNSEXjAZgVkk4ovCdrXV69S/4jZYZ
0vBgWzFragxhtCbPgYSHQhmRqCRBFFuEwnPPxur4EHjjtA5Qj4LuiLhAihx6pqMO
TCSFgxvMkcutsPVd2XJNZs1Y8lZiXtKifQ8uAHWBVjQhu1quYY8aU/U9OMCiuV8z
v4wXdQdGA9PRpP8A6mYiDm9f5/9vSwpWKl8CFtalRR0DOLhPjmYF18s5Mws3nhcm
rziY7o/HMXSWAqi4LMGmjMzVMsXw7CN1NOH7BEe+4gGmdAbcoHFF5jsvup1UY9g1
MYv4maEvkHRqTMGlgcklp/PVt2KiZg5z2sVYHbzwjdb2c0/yR0tgRvrAAHWoten5
2X7q9y792itZ1LpGl6VagkWCyoDMugt0HBoEPjgk42jp4Qcq5EIf40MRkzPKNlQm
TiICMFmY10AjionJKPN3n2b2KheBPGNpKSEKttps6h2Cht3J34We+MTPuj5jiU2Y
OMG9CpujPOxyGeoz5EECjhB3atgenz3bshJ78Y+mI9aDWk0LhJgyFL47nsd4xHpB
rcs7UYNOABpa3310RkPPqtc5D0xbboqWSaUvFK0S1IV8KLCsL3FiSkGGwAz5XsrB
U0VbUy4Tv8VCoOXO/zIjV3yOSb2ngfzm8AoLB66pFTRKS9HBdp9CSqAOJAUS6QLG
cvBQ/f+S3pmfhs1bHDRThXzc1YmqwSGjwbD5rfuytp2vuBWo1jB+3o6O/Fwrs/6/
iyxSN48aeBb/dt5y8hu2rCbmb5oZPPNOEZ3SUHDxO/Bm4RsuZFyVmqwBqVrlXGkf
n2t4y54Z67/GjgLeTNGfXre7FVjyxLrG7+La7gzabsGi1aYkpkZT2juoQatUTnzi
tNjZj+fnphqx+jjWGqdEFmZRaGTWQLC6mw9c1ajrM5uvBzdzZVqZlNiTr580cvci
HWCWN8+KVyh2/g9RGrm+M1A2BrboIVHjKKWbrEqqvroNbvQ6Fc8us29RULG5No+I
TNY+6pAJqWCZKqYKKrfFs8oDIO8sDK6qCqq9j3ULGAlSTFds+ZYvxKR2sYKlb0a1
Tifi2aRjNI7oo89x5Xxcos0Wwu/cJPRP5ZrxH+dQ3q/1jz1AWsCTU37RXfVJ+Klm
3dbDf8DRRHgGUhXHg3DPyM7a5iqwpYuGP39Ywnx9KutGxmh7Q1v8LTC3X/MA/LxV
IC1jcYSx+OrX0Oml70c5YF5NBdqTZCjUmv3pF2aIViHqvyNf7unaMIeCcxt59+6b
lxMqlTIA0ltn8000Ikv54ehGQsmuXalksrYGZJPafywNMj34OFf2ue73irdfNnOI
EAM5O+YhnH0Ums0AlxhdGQOw7jSAH0exS3Dq1/1AqFLO+UZehh/jgZnqW7ZZ48A4
g2DhDolIrZgLkj/tMTPky+yhd7BSL1uZIDqgZL3xwH5fb5DT7isoIFl1PQeB9gH2
Tspb1lb8roGEpvQ0YezbRR31if5cnMg9mYUhMAwersKP9F/C0Zdxm1wqItQsk2G+
2Ai72SnhOq+fhqe4SZGi4Xqhld/OzuKMsHoO9TikUVoslZE1Jc1LdwqkFNk+0Fwh
QvC2ZlRyKsauvBE5rg401Yo5rIcTLycGf6KeFkttRm7s3iFwYA4JilQLcmP/d/x2
JidCOEVVYB1AltlWFv41HxRxyOs/6wGZ+mY87K1Xrs5Fwwo3w251OXC5pScEMXzM
qyj7gshauhje+2OfKyvfrf0pdsKYZAxM0LQ8Z5Yq0uA7FSTlJ+vm54v5r9OIH2tQ
FJfRe0EZNET06X1Q0Fj5oBA5NNckUzt7ZWZ4akase03sWWvk2z6Reau2t2OQjbA4
+SQBWohIBXrwA0BbfsrHKCujL04vEwcDwN9uWOebgB/W9RnJ5mT7hephLBF0Fogz
b9UPzb9ePHX6vzhGbI7agnpG4V7f2uL1bY9UmiESzBacR5mOUrlwUDiRrrrfJiu0
NM9z5Pt3bVK2BGdeTMR21GDOCewYw3zWcVMa5CjF+40r1yde/ZoNegGW2hAPKZ8F
5U/vZ7jN+OuGgCvBJiULSmAKiOIrHJl7ula14i75IdZCGkBLejdrKCUDW1yQAlyA
zLwC7Je/9Jip1YaegUyCVnJyfvTrSmSJYatnQ0aNpxD703X/b8fFU6w621ZN0lsV
DKwv6Q/7DgTggo8Ut0cSgVYgTWFEgF5JcktHpKyRYMkMXDPoc18Q/+ZEBF/zad4P
DomtaSwE50fSat1LzAUrxXdWjjY6OxOZYkFSq8DxI7ClS07NGiZdn/CytLcGD6MT
fyNgBsGcdD00+dTAR3n9DOEyr6YVF+Ms1x6+FyO68LKOkXJAslhoJoPMRKM19q3b
UQ7y/vDwBKkyiW/ZD5RQmir34bfpOq/zsBpT/EpnC1cbldoHp0ebrG3LRw0FiHO7
G9FvJinCHuzsmWPxP97SPC5SYMbw56okunKRhYF6tZrFaw6CQXqPSzeEFQClZQkM
fPOw6JtRj6pV9aVP5hR0jVdg0bg288S0sc6bGurmyr/cR+P2eYM8AtO4Y1kvOtFs
uWMWOaJOQtZNTOiU0kizlWR1Zm9wacPNC6VmABOtZWMw/q31aOVv1/2RuS75x2M3
pULXc/W/zyDeBi9v6f0X8dqb2u8WL8qrf4MPGw4DSyUouMjV1n+HQwW3pmAXZVnz
v4A2c0DqU+YTtMHFuCCcfOu9ISmnkWp5NcB75EmKDbCJ4Ihf+mW3niGCzXDVH0hX
RESmiCAHUKpIkUPIfH68vUt3I3/Ga28RRKLAVB/CoMMRVvunDPDIMjFJgka/1nEx
MeyjSCDJblTY2e85CvKojA46JbQBps7Eafh1MXiiz+VJFwrz5+ptIoe16VMVAMxC
Xpf4CAE7SSx2NVcZ4VDOnf4JUjttc9wyAI/Fr6XFQPfyqzPefvyPzuTW8ZMaBkyL
2O+djF1bIiEppxB6PD/z+egkRj7+lpcQk7AksbGeDt9F3FxdzqnInuAvMbDX7ZPy
rq+75hX/vMMuVK2uYHnzC6gCcCGMfaE9vCtk6QSzTPQwreiEEN9Rz1aPtJ7xRii5
jhzU7mdG3yid8SNlIWkCHS0OYmHxLn9HnteyjiW4ndFvzlZcRqGaWmnnOR7zsXWl
h5i94OWf0Dc4No6/5NvCoXoZDvwWtdwF6P0S4JEp9FV2iB/pZD9Xltve7M/AiAi9
61x16s/HrtZZLdNqhRz0Pxd69Mu7GomucpSEsmJNrtZ0+kHXdORmVBJAFCChj1jJ
1h4Qk+F2TGUmX04icws6HdCogN7f5jkfVFao/rUaId/4/jB7q1p9aIzehZ/gLiX+
N0aSeZy/dowBsbyxTHJdhoIJraJELIpK8VhPGesk7Kj3sKOnTHQzrZjJiYXM0QbE
IzNYE/29HJV0JqIKwdLcnWCunmWb6KxRgeV4hEQQb/9PCFGCvW8LjRTKjIG1nBOy
sN9ENcRNzOf8oLebawvELB3Y6iAwni/3HjVzzMdiJlbIeYvFGmjwmkCM4GGWlY/0
iLiYBmRQ0qEbk//7+9ZH1ya9kym1lIgULVkA9LqDKMuMskenwk6ijxxB2ihWOtKY
+TSxHqIsn5LKVQIO+3WrtB+uniONYbyzUj039tBVEdYowtXXu1njpREAaOBROT4J
8Ty1qeQnaL6n/ytPKTVJ2j8Z4jki1GB10kSB0dcb2wrKlzolT1yqM6yjoKmYBYGs
y6Unw49e599NBc20vkXYK00JSAebH/0GAzRZhFe7HVYgeBTZCZC7ciafr15D2RXf
/czfUh7FNHSaNbxEuBxfjkUlrrA4e4SGUfSMZPqs2BQxv/2Tpf1wT/2tFe1wBtzc
tHqkwwzC/KHZZ52PZfR759BTfiBjNnze4eYYX4cENVml00mhhan7fiTYW3hYMQ1d
XSf7RgrrK+ORLf+vLJHGbWmrn5A45Qd7fsGh2Ew7lrEaU69sO4s2BbiWZmb5VA3K
7BUzGYMS/0oEpGpE2Xu/8f8pAUQaNWv7krNPl79S7gF92XYxQdIymxdZrNSo9Ev+
XY9yCQH9T1pUEYIi1tDu1GOtsZdgiEWfIkUCA/JUlOa1P9KH0kyNngx2RkjKcNA9
/299dOaUY3LPlnb7x/W1n6+dlVaEV5swju6flbaSQX65mi/PH+MOycB/FWBoLVrb
9ibLrr7/8cp8As5eTnuanGBCKfO2z3cgqovOdiTmcbuG5k3gEleK6dHDF9NPbonf
5Ga1YTqWlr9M9Dds1luIy3W384J3Db49QY0nWJ0i8L1wQggsmQRk+TivQbD9WEUh
pn1yTYHj3KDrW6yYbNlCEsWVql1NL2n+7AR6YT/M273lhilVM7Ro6Yifh7mCXNDA
zkAmBkfK7g2o6/DcIekeYLAJ4UHwcn3HjHNvgKMi7UkN5vyj1rXsxoRluVmymyB7
UNpYOzZoGye2Z9upSsSgXJ4cNKH4rG5f968xJTfr+avaDAOQinEnwaQLpUPQA9jV
az5Ldwx9Lj4TjiERQcZdHgmI+9VoPf7TC0jyHMfhhCCfXxnGAXSb4iY0YqBZ64uY
5iBi/sUHQMFbdkFmU5Jab26CX9ULSwDEoVd2YBD+vAdEwrA7vYf7QmqabLuw8sSZ
5iadN/TazQWuxliYJfDkynKALGnvuQRzq3HfzJ5+VWZvDp7k8trUkCidT9AKKbU4
qto2hb5ju0+Mwh5XCT4T7Rf89qeP5UDnS88DjbsWF8ZM7zjSFPdQ1EEyZ9mPKSzm
iV4sHafJzpJr1k5tZoGFAsqP4UEbkflnOpePHkFfHpjp6ttY0hZQ0Jbk0/8OJ7bT
xVMYBrCKUg8kW9Cqt72R7C7bckr/kJ23baqq85OEtM98hM+s69+ji6SKcCNZEjVa
3zxxkr+/4yypA6WLohCDyXDiPMHtuakuB5lhjEL4WRUlWrCR/otCKBtr23BcW50Z
17BZua00sbC+MViLi2zicc6EKcrvJWVFDyYrWOrQoyPGRY//ZGH445H0UjosgGbF
68yyQhO/8Vi5kfp83vfPkft7sQE7bA53QBntGd78P4FDVfZj6C4FfTxdUtQRcnzS
1AmqwLtxA2Bc8MfrU/oic93566AHValCcaIAOpjrPu0iTo4WdOFDuCAbM3sQoAgj
T0LRQQoKp2U1/KUS7Z4Le7MUC937u/XCHS9m8qCPKL2X3aiUWElBF3V5Zs8o/2ua
tbRsCx+IUyLVmA7YdWw4gkr7S4ofijsbo1lPi92oSED4JJZRi+wNDS/1rv/tlGsS
5L7lxMuXD8xueWMha7JfPq2+HvMZit+ndt4EkviXhuXjPiq30maPj2ZaqnYqH1yM
2qZbpT7xXfv5Ex9NenRZMYgU3DDwhoI1tjyQMN1C+fPXf3qnCULfvtvFOI6Wu2+Q
VTQy5G7ImhsRiCEM4H15PNCyEfRuZ+ItS30EpndVxQ7/VYlKX0t09lUdO05My3CV
M56KnI4n8driyUKJ6/iyhRLIBsCqclo3FFrxIAVavO16cr6lH3iEniXK7ys3OKLQ
tm9pFpcnEJ+2VesW3xi6VZMhhgHkKLeWecg8uURAgiqi+CE8bQmH/slmZV9q2edf
VsXgZWe1508EYKnnTrG2KHb4g8XX1cC6EXKRCLGHfs6k4DakEgaRUA5xQPJaCU2R
38J6GtXn91qnoMuyzjjocgUuOaIvB1Tps5KXvSU6o7yDM3viL1m7fHMsxIGBrnMP
VNBbw5264myo2/lw8gSMHqRyQ6xku1aVUd8tcBDtKeBycJOayJ+DKDTwLaiYZhfZ
IMvduUi/kEjVdbZiUUKLEPf054LZR4F/HS3qyCBUpCanQ6In6fRSglc7X5GZKJv3
FDtxe1yTxddtZyIy4EQ3hWEK5h8idLPTZOqY9alJfgX/itdPz2jGk05Gczt2UsmB
O8S1YuUYxuNcPkr5vBzyTp73NLIsOpDM1K4TcgDRGcjWOtHwLn0dukludBZ5CXX5
51M+7+ud4Tq7fYsLqFGpdQvJ8/ZJTe+IxIwAyRGmTd8D6Fu3QrPDZBIPqe1j0r3x
lu/1XcwPBW4zLxWxM0iXskMdN5CQJf6Fugh3fNGfH6yt+iVIyOEan3n/rTgj0I1u
sA88EqxBO185HRmSBvKVxq8/k3/D1dcrEXQttihrHNJFE10iJYI8y24wiOVw/O8g
zGVAq03kHYI/Vfp/uYe4gVoKsMauQlRw9/4wyuEtKF45KT3XlYt7ODNNztiUjlGT
fScqL5H1BsP5kl/+H50zHEfDeZUAdE90L6ued3TkcpWLIqQgUajy/Wn4mPej4gJc
TwdPePf4QK3GLNOdFiOpBH/Xqc/1VXmFZQRZHR5f2dipREKUY/tUse5LYy9VD556
MD+6kHK2vhKW+5f/EKEfH6f3zBqnabKOx5u/evAr0xFfayJMcKjVBblBmiq34nfg
9T5WTKfMl9mz8o2tOGBX9HgwhvYZ7PxcP1vfMVyQCr8d80C2eJV1FHJVnGBaCL1I
eLcd+xxO4NoH3LtXB4Q/0/um9SJ+XsaldJ63QTLEpradAVWiCJoqnLgxE8obuzPu
ZBnFNH0+exIYZyu9V6jB2njD9JK8ejbKW/oQcRmWPrhWABrkmQLr2GRHzkjz54CU
RqV0bqqPxy7IMoA+NS7Tv9OIbu0uI5qf3cSUXfvV8xCq295ll7C4jiFsowDO3dKh
zmDegrQ79qt4bmoxHBVCm4hgp7yfuO/spjY/r9RvF2yQwX2EODZFBV2+Kzx0YooB
5Aukr5lQcFB0qnNpvgF3KC3+tAx5xzG+P58jaCcklxH2+2Ar7xjtZsawIaZI+bki
1oHFh+hpDJPaYEfVgB34bHOPo7+CYt3YJeAu7Gih7W/alxH56yMXmxfdnkfuEKfz
5qhyvOhtY9GBr9PpVOOyd118T5727pTyZCGOubdco0QqMk1VmXyk0Z0W9z7EOiSI
5PbbccCcBRW5NURXdeXKxO4N9k1POXs2AdP08Xp52lpuFHaOsbP1gfOYrp+4hYki
yA8L4xtKhbQ1NwDtoL2Bc1XkhQTHh8PeBKd9yU3HWtvo+0HLBLYE3NVol6dq4a7N
H1wzCEIBASz/2eOekJBgtuZBW0XgZXMcnkyXFib0UyHcRJrsjem0mZApb8CsY7MA
RgCyDbfaKXILBq/TBqssS3T59ytyxIYQVDCAR3bQc//IYQPYM7Lv59MVYSA+8As4
wrmB4bOcEZCX8xZY9L714HItX9Sl5Fm/JjIye3wnm8+22Vu8l7pS78+iwYn1Rm7Z
X0/Pa2e42UMZGSNjsefJVIkpb6YXRmIz/6622aL9IueL9DgIRh19eYoR+rO/8E+2
0L+lS0l6Ri/FvzBs36IrvxyZHAEluVqnrYWIXLFuyDXhAUeU7o5u5CXD15vAOEHk
00p+ohvlkFMYSu7ZLztoyhZ1vxtudNlB24Q41HEQX+/L5cP4oAs+B4m8VnMybxVX
tQjoWFDFtkUfTyTnxHfnIj5OlPUs2N5gsrUzwv+5bEznFPg4gSYttibGDY2KBEOG
YBhSzg1/SMiT1NBmW6LblQDharWm6sdmYQJlJX0yWaDWADjz/0fMadZgPyfrGJLC
wSoQSIM/DdGi+WjRFfMJWL0LBCFuThtvwSE2J21iiTy3LRMHO8YoWhrOcm9oyYna
2z6oZ9JBJmix5j77D4TSY8Czd7pyRdkgFGcjDotnk9yICGX1mFV5wIji9mPUyN9K
NrvfbiijOX58Ks9mLjk1z+SuWYtZNrleaKyufoEETQ7RngqvWJ/uTZJ5OiVpVnMi
kRlscT6s9pQkVRMFyH4MRyGLdx+l7F+PFy9ljQKZ2iPHoCALYlhI7etTgeeYhAk2
h82TdFw3pBXDc3yC04a3CyIEWCC+IE0ADOFbvaH+5lx+fGfzI61yGtBEelGw0hPn
sBYcg+QMOW3qJSY+/yJPmrnmzYx/nliAEm6hLo0yd1PHT94ayR5LPYDdlgRtGvOs
vtV/aP4SAFqGJyjaXlSkh+tFFcQZhXnGOZnR1Yo+PQbCvekkWr3I1NhqgHRCg9Vo
fJUVr5Gmi9zl7uC4pQpeh446ZUHIgAX7jZgBWAnhdm434DTjnoXVZ93scf1RmME9
SB4JspcAmBnDL4kGtpmxS52ehBFVu3SC3e49+REM8nuijF9Cu7hpmLxl5AxDC7F+
m3evfC5j4thvPPOJhEmyL/r03FhnjvNwK4AXfPEWI6j5oopiZ9agqfDKQKnVaw/2
U9nY6uuUCSVKeA9kWDyb9CdZa1zCFpPEiDd2ulFWw5hC3mQilw67vmG8WxmGxMad
Q/HCFRdgKxGZkYPEz0wvCjO6ql//SjLAULTkG3TZVAe/dojamZ24ntEEBQsojsdE
mVAU1ZHMS6vguSqSCIgG4172Devr7EjqqdHcRwqxC2LhaVpD4d31tQilpCOue3c0
WJYmG0uaFpmxgQDV7+J0DbBx4ApDlsVVmEzV5mV4uFAWvJxijCIu94A03ffM6saC
9GHOM/VNvmSNwS6ipn19C11jooEDPxkAJuA7O0WDPJhWYdAGesf1MY4QyATf9SCG
rT+whVpYtLdkDlIsxQtzq3yo1AUkl7MCES6OPe/jhKOcSDEOJw2RklprtuA8Z7NK
CAp2zcIKFae+YSofVxgFGo6dyYXBtvzPgV0FhpjV4AzMVndq0X7zno/UmNinPkb5
N6niOt46SSeVthxzTx+aOUev4N88EIFsF0lj0eR1Yrimf8g6QpCXLMMMU3m1ULzE
daO1bzUl/1dx5Ew6sBSUPFgKSWjQz00aa6Hx3bsl+Fsp9+NaXcK+aiR6kZ6x5bvt
MI10xYDCIgGGsMVWJ12rS4Cjbzgu6PheW7uSSTPzgZczaoRxhVG1/kLrhi5U8OHA
ZdhEHSecO9zVvnFL5BwlgqlbJM/aTuiha0pqZyzU7aD1EKqfNJArxfPYN9ShLNCV
8ZG+jH5HlLdXa5fT6HpK0KhCpS1TyqIsB4tPn1iZC/m9WmUT/jft2MokbVgN5nUX
0UI8rteH4vaFOiAAzlx1UfWtHDurfLPzuGFd2fbDRCI8FqrSEpB87vLbl8DXSqwk
tDuT5hrwBA4fQ5OSpee4iHW4Kcu7T8/vfbSJEsl+v2zsI9QE3wMD+9pbdeH72z4E
qo1QxI6HUsf1nQBfLqF+OV0hMiNQjTUv1BWRamocmjXOwfKqb2MCp/C1F3/OXeFQ
BIZLlLU87nq42WX7N5KWqRQCEpQMeb3PrP2zyLzmJKZzHLYMzCXA/eHbE882VR1i
XLIt/vNI5c7lZUTNbD35wpH6F90BBORfE5BhlIEz1Nw8sgBV+UKLb6BlT+8uQW9+
LVuPMcjSDSdJTsH1I9ZvXtENpRCL+yoaS8Fb8l1JvU35ZfayuVT8HPUZvaGBo4CC
oX26e3XI+sYzKbfDnHdS1Z4Tef8Ltu7VsZ5e1Rzrt0DWN7iONafpjF+u75GCiNR7
KyYMNpXwZCewQ2Ohip8BKhymOVrw5JngclaZ591+YMAT0uexPp1mo1E/SOpFnGj4
3n/KsfCm6HEVzdiyilof+Bb7rdObVbtao2mqdItUEl94KvwKER0QmA2O2Hhrt7fG
O2BKmB9vuOtGNwG2UL/IfewIoHWVBuL7frklirpnNppjqt3toxQcVmChjuxZ3cyS
7Sl3PwWOWGVHKRYwC81haagBe7nqVEWwWtv8pK+AQ4bxZC+1+OzPSPptD7Oot0Wk
KatfU7NA5pnVweJ+ajJYN9vxt80LkabI4JPHP/QRLyFq2HDskiIS1JvH5TjwOfT+
tXB8pfycnJjd84A2u5CzOVW4Yh+xlZh5rFLWzJ+MtthWLeFMUoKicjrjDnXWqZa+
6TL8Gaaz2p5hgcdSPkChCLmpuXOKgaJsErEBDjvl31SmXcmnk4Da1axO1zHYKqpr
lMq+jLWpiXnfDCiVa2EGo30VtELNZOdBCPcCvb4CE0mKtw0bTGtnx9qTaDiwtAN7
C2wF+wFI9ESrez2nVi/wugTz/6+fiag4aoxO+7qviG5rAbOzLbQtWDIzlfh5kMmP
1iXPad0VFyKEHH71Ge4rrdGaZiwPBcqOibPJF6J6Q5bcFS7dXvalrgvEMDf3qzXh
00wtWrnmQRr/i9A4IuC/LMSQKqSnDJldS5IyJWb7E6ikHldxxs1zVsRgRAvU4kNt
hXKdxKzpA+Auh2PWctF9ync9beYFLjPV9hWXNpN3PY/rA8rKki1Ig6TxGCxDkLd3
Ao+GbAPc+SI4UcnMMEn6AvlznRAS9hdqUgDIt1Hpa+2P9R4wHE9GsFPmB0msLmmR
KEBbV+rsawifZwZGzp0V1aJhl7Nc6HgSqacZMohONy95W8DmiIhqjR/kUOTNRXFh
Pq2sOYIDuERlXJdiHIGShjv0gQ5fwJL9j+1aQgxpoBzkwY0lyuRJ62wE0oNCyUsc
cHpR2OKk3RYlX970lZDxiUjrg5yt0ZLvWMPCeX1u0GTwLBJIkclVtEoA6NFLKy6q
Kg1qMFKGQ02vf5tsM6SAHtj4W0ZXQQ/QFwWzFrzKK68Gi2BwVUnoH6jWGxNLV94C
OeJH8kClNgN396gvg29LUANgZEQ4bwEBMUiqyLLxWXsXfs+q5JPxLFM75gYQ5DQe
XDeykmoctFA4/L4YZ/hfktU8iAY5Ng8gWTDa/2GeusfgAR44F2hIE/+SOGbc4pZK
KRieNdy9lyuCYJSVz672BVW3O4p/wAXLQqKJee8XzGGRV+LUnRl1hCsfEvwWNPCU
S04XW8IPOr+f6SWVkoc3TL6avwGhoP9ca5HNiHIo9H9ssOV16Fzo1/xcdIDf1cPn
x5faaLulK2r9lHGAT2tBomGb064JRxJhGvC2Bpu3bh0SUARPwa4wHdHES++T/Ny6
3pDKcV81slVzH+enG1DVyug0dnf0lKudw35m/UWTwmG8dIqaOOUUSo7w6Hf1jENG
9pcjOUMIj2BiRmkIw1cfo/nFk37RIELVOc1/+7DHOzzcy4I9opaxM2H4uOj1F+Fz
N4AheCWGhiAOLn59Cv2yDT6D+moaE376kSXEvnU251ha6Mp6Cpf9Gj0ydKJ0HOuu
xh4l235fKNhfZvra6ai3rtFOmlpFn77whFV2lT85eXmpM3J34Z3vovTBxDE91Fke
mx6a1l5ma7LUaczqi/cPBFQhIm4QGhwSxxJPuv0V2bmkiR7TVJlG6pBU/zs4Q9Yp
gU6uWMQ8alEIUnPif3TEJ2juWs0kUBrdd+H4JI4sxi7eIOW9gZnapYNEHwpKo79w
GZbZ/QTSiu7FQ3jks1FaYu74JaKwI0rT2Mud5DhH7mbIlzCG4j3ETn9AD/A4jEOv
SIscdMTC98hI4iUczsnOg218IIotl3AkzF2Vn7ZabWbB53n/5rYpUjkV0Zx8ZCdq
k5eeSjcA6H6oSRw7FF924EGytrujsPACYNNsRk+tIA7Xvq5DUO10RkUbaG2QqZB1
b3YX8+GC7ZUf3/pKvUi2xHT9noiAAYDSI7d+HxosE+b3y2kL/r/n/kEALkzb0UsP
3tUSxVyI8afj/lnxzCzah+XNhEUfkPw5d+qcUs7y5z+3U46r8CgEaJHQ5peOO8nj
YIpcNNO1+GjQ389Fse8WG6R22mbGwPonzvjNRrVRL/g5FLlEwAsYmRfLSkYeiMJP
BkudXhL4U6ICPWdRyCkN40RGSOJ2C5MeDEM1GqUEAnVaQAZWvrXi2aG6yKBoZA2t
d/Ks8Du0k85A6euwocGFjLk1Jes/RObKuL4zEikf86iJ4WId0MnEaRBzneMxLIw0
g+1EETKbP59EgAWtQUbVyJzvDJsKj0ua4dssjbudzvZEc0EAhR2DJY2jpPk/MGQR
xSWtsRs1FG8wdH5fJ92phaXz9aBUddfpHR8JoUdXT59embRsiIeKZIq8zZFXQC/v
O4SBCXAqTFVA/RujHAJxyiDyAm+0FX4MDwyxUPtOkR6m0nM+/tX4PznQD5q0X6Au
JqlHJm6+xG63YbClWqn5nG1vWRjPjUQ7fEG+O+4x109iiL2qnhTIg9+274QRWpKU
frWMCxjxQPl446Zyr22w3eTc+OPssX9iAbVB5LC04YQU6TkiNruZshLiqGPoHxG0
DxU4QzS4u/hmHfo95QVjCcM8xfvCYmPt3B18nXxXyHfAZGuZCpFBCMln0pkUAZdZ
DC1/07xPbQzDEqfzd+TwWFApa6Fv988KK3fWTcWOhCnx7u0AJXkBfYs2WVcDrtXx
OtY4xjx7CxshpnjEUSVSjwI4jNwExGfIcne8QJsFP53BcZyiHCGp2BGpgu8axxmo
PH3lUe5swrJVOrh3yHnq5T6TSkpF0BpqDIuNuoVIdYXqWLxIoUwlmqqH1+HS6m1+
UTeUxbb7X2LXaCcfsdAEPcSaFPTBex+wb6L2a/J6OSkNW7JpamJt9gxIbDvHZLY9
scuy0Cv+p1Y9K+B7zy5XLFonVv2h/U21Y8F79dlYGSWlnS0xs7GWeP700nxxa0Ju
Gy64UW5de36JOZggWeEpfJDA/N3LxBzT1Lj8RTbcAfa/ETL7EtFBywRZKRNvmggK
olRrVmcgSTlNjZMelGEsB1XRwvSywiYSq7Q7l+xC1Z0FLGN6ieK94rBoApJz7M0V
IeAHgxJIQV5jsjFpNvEPPqoCVH2zuWWzAw2Aif88r5aSEuFmbKILLh7XN7j+EdAL
4XxeyoBvNtNeb7DlmIpI9Qbgpn6Th4dB5bryqmav0A+o43nWa4KodCaZhFi9KPMC
8ySB6c4bUxFx8bd+et36ZlzsbnXoe9lMW34um7NQ33buogSSBXdszmpK/VDVtwW/
rfa9CCDjJg9INyH9kXZJfmBBZCo8vmP70G1RLjiyIeuz0qmvjLRwk2r0lJf/oBOO
jNUitknPCd/3Jn98zsJGs88e6zEPXIexop9iQN7mDJv62xS+XjO6FShT5GxICDr/
zIQFhMpp+4nSqNHwRmA3n4wy/xRU9FSAk2Jtaw2Te2INmrwXTx6EM1PAYaZKtrnU
tfoQML9vJ7xBVkQOrMasz/KLW9LbfIMqlJa4uaXL8xigYtDNWFYUvNRDWjQRy0QD
hbY6jY7fghhjhPE09hsU5E3tNXQSVCTL/EG2k+/L3oJvqmUmHmEWEwOJJRut1j2J
CLk1LKqyJibgbK2e9gvGH4EAdUWUISThxD5apR28RWLMHqCMyZueBZCPf6SahTwd
DU9iySL087ZHzmoPuOCjYpHwO+roRtm68mVjkJweWeMWL3HT98vWiaFWFc7mEF5p
CwHvjVNBGLJJlsQAqI9PFWrx0w02zynPsw7ILueEkmBnqrDuvaQ6xNLj3neBS6FK
wjdmcDrX01T9Hw+AoLloecHvYt8cGh/jlzPAHbs/b/hQhvuKzuumdXlAalDeqIJL
9UHBWD5uonnc2alf3R3htVzMg7PBcGAYUjcg7gFdPOVFklYOGUTjCuAFy3Uz39b3
gad4RbsI0cUtsJKOdKbutoqTTO/cLkZkR4HZ8ubuQNNtJAkgNFuyT3f69QAkeDy6
wSVU9b2wfmZtb4GEtaqSFnVt0ldEl1KKT8+KRU0KAqiEDiVQYlAkrYCdsM2ASkYi
r2Nt8ClCsWdYfpyAuQ/Sz18NvQ0aVDgpfuMrEsOFH1ud5Smqw+tvrCOGpupVKWMi
xRpexYds236bQFfnSxlSNdg+Sb0v4ypoxY5jcgCe0mAwN3l2oJeNTCT7olcOWXkU
2oxtLy4TA6VSjMwNyeV3gwZXQzj+2dD+WZfiycOp1VFZOMNTwLgOqhl62GShqyeT
Whd0GBbTDw7Xng5j8JYpQ1lAIi4p7tbhh+0GUkIUgzblWwZLciXda9BMFdi2fLPk
J2PzHUwWyYb7JEx0P0MZ/TVTTADq9gFqnoQSP1lygVlKCkcY5dQ4476RoVkdlCkW
Uxxwc3yJNr+R76tIVGcgv460lE8IM5LeQIvv1K4EL5WxtL3Lmgf0JrPH9Bc56Q9h
VpbqDBL6nbF3QKh49+wvetbNrHVvgbjD1vV8eRrLnh7hWVxTtwTVjhRCTHgtGsw4
RCK4UWjj+TLTv4HK+WGXKDigMxgUNal7TMuu0JXNJKULOOTkd3IdefU/GkB5WbYi
lXFnk7qaH7pRcxg41HM8P5dA8qjzWXmZZxGO/87y+2eqXRJNe5j97dOngEesR4aF
2PB4fD6+rR4CIu6l81Eqvc5XgdEU86OMlIqwQbjEDr9ZRHtl5hIMZF71GUYvbno5
CAm6IVGeB+2UjGfRgmZdAPfSNWSSAa3SxdIHNAnn/EsCU1PGSt7Ub9Xw21/Rlhgw
NViln7D/X2xOQRTlnMepF3CPqnf5gHio1ZcnHzRGFsq3aAizkDwiUpJI+zsRmf6A
+5uvtCjdnmB8J/iJHjpz0Tl4KduICBzEPwJhm2oO/tl+eYE12J5sFuek/6UfGMUU
CFjmMng1I6YAtW4wP1opSwQMdjlGkNAgfldu/aT+UxzsD3zROJfiOrAIlwlONEUr
TREOf+KVqkT85++PfLctBHGzolVf+tfkIZfSoL9vHbg+U1kGdTc24I5knrbVIPJL
U9ACq3TP8fF9R7Lga4lVdobQ1d5cpz+SkYOJx3p7Vt4DbIUpC+MgobsTAgbXXIZh
6b3FwzJYd8s7yENkGZMBi743sTYuKKxnM09jm51mD41YIatrOnjy6n4gn1MUwIa7
FybfX24Es0EnuxZ8eYuSLTD9QG8OD1GeSofdUHKVSqfQN2b8DQ15E2W1qXBiAFo7
uQ6SHrFacMVr3KKZHbUWFQKu9UDGB2IHJB4hR/X22FUy9e+W3pBQt+/mYGjIodSY
jCNXRe9q1sYpupY4reO3vwcJ8Lr6JPhUSF3cmcQ7nofpBJUmabGjNEEbMf9kbYHc
s/RLK36i2lZRskB8umwXyp7r2sSMi1ohAbhvfnZVyZuh5F1S/+TV368ShZVgHW5x
Vjn86RTXlnXuq+kSJOKtXISy2RDh/NIcJuzny37UI8pHcq/ab69vImkFs1V8N35q
lA1h21a+BuUIqk+psxWupkHwAIzcy7YANFCCt0DTeF+gaMYZSH9rWGbFVNhmu7Ms
mIuWdcixh7acnODcuOtIeYVWDVmmrEnu8rx60m1Vu2MPKdxaEu9qJDpjGf4o7n+R
MIIoet1JbuKXsKG2KakGTx7RnA+bXguKjSugW7wO/QLZfExtrrT1aR1gPTxSg8jn
RsPdMa7I0TEN5YtHFqViVBe3XqaIhzLKoA8QMFiza2NfAksQMs1Ff6t6rXxsgShM
ta5ZCDDR3D99dLrMmk0XUlDVyTzW7cAWeC+tF2hFgVnJ/q1IPpRyuKzCOmzocwht
0zrXEPAgSdeQrfoutB5Beh7k7vUIKT4MX/Ms8p8wGm6YlJQImh05ms5jxu+xu9Ra
8guts11Mc2cMrS3f8ynPfzhsoO8CF/QoKc1g2q6mPvxnDwCwCv9Gl3nzwhowkFZI
VIbbWFh9PkADUufTP1KpD6AQFlejwUcLV3dZ7l9Bt/NqmqyFANj7VanmKhzAGwQZ
hx9XGpMf38MVA74qM70IoiVIe9Y7BsvCO+c0MEOf6IaAtYA2L6Rqju4bXnGg+5iX
L1ZqBeNq0mmHILVVLNpKJoVYfuFBQMRXTLKwnHvAbNMm1RFHERAHKi/tetmDb57c
u83w7bayiHJ0OwKkZmQs2JCBf0KHe9nEITNMwnE0RqhuOVakpZIMRX3xci7PVoxc
PTrkqqWpcbdzCrXPNSSNpgJB3kvTp+XZY2iLAPEb6GoA8YrEgrOdOaZ6FU73E2Vd
bhlAk3pBUmErtQbIKYJytLPG9/j36oax5E4VML2pVmkeWWfeb0UIuHbhTeZrnepp
+hZPVch4s7djwUseQY+WtJ8aWVJb/ySYmQN3HjHPLi4yMuwO8pXsAwODabffFZLX
N6gRfthIFd0SoHP8eMm/eWytTB1ed2Ltj3F9wpo04urSOARdh3AqVe/HMjLYNU+k
Wg1a56Vpz8U1fvKjZAuMHy/pHWD4+hz5hNg2cF9yDJZyPEcUTt/dMPLJ1CskHfLq
mF5/2a6DKwOnhHthy6VfuN3ahrwifqflNKb0A4bPqG4ekear1wnhkk7LpkFByiAg
HGtfeMaGRRML+D/IOEuQuRGRfg6JBpqYkLnToXnK8rfG4L2dWJRJ7Pf8wiqTVbQO
WYEF6qQS/nZu838VYWJ5NYH7zVphdbkyNxQUyaYrliY+6Rbo5kK6PhDM90RzDx25
2D0c1BKYo7ftueW3AOG082so1gwG3cf4Fdt+DC4g8zCrnYHDhsOlRKHRm1t4NZe4
AElpcBimwb9aEqseWB12Td5YV+B62eDisv/jtYGJw6HBF1cM8i4pvlc1w6S7RNp2
3u0tCxcTKTZ5Mw2PbHOFiH6lhb/xI7lHlPRDaJXv+mw3vkdu98gpRimjD6FjJ1pl
7Ht2b6JFzn/MkDUzNXXCXGF6Sg0CJQ9AIBXUKij4PG2VH+XHWiQLBdjvk2S9jFus
E+wzZlfhSizA003PdA2DZP1HttmUf3T/B07f8POf+sNRVw+ZCZMbsqtha4L+Refy
uGE/dxzbbJPQdjeoz/Z6rIQYoR6e6j6c3TaigC9XiaoP0VdPjtBaS+SyvFJRV+Vt
IRYLbKpTmkIrVRO0E+Q8HUEiCFBFvZU2t9Xuq8IK5KfLRUK279VG6U1durGdjnPd
xlat1LQ2oy61HwlIrg2QrWUbQtInKQhLjGhfQFwL3TsVW+Mk/tHb4yf4U/mULWBa
1y0lJsAJSFf7RYPler5Gh6UltxVKZkyjI7FfmXrzyinSP/2uCDr1JQHC4ONOQE3H
6EQmq5J4BH6l0EoPOtbOe5036iByjcd39a/eaDitaLIxXxRKZAx9ecLr5zi51b1J
rJkkQ2XHm2r0AhMhDbGCefUcSmdtbrIw+TakUF8UMBGOPlfZZwPlZ/KdVhgXQJ91
ZqJ0MjwndbhsCIdq16SnmvQLN0vjxm/TbkLvQEf1qGKR7vIVtofcYz/Sg2Gubqr8
xgdEzNjKm/Elsywm9uH8NNKMUBTPWBFu/lECg5zcnfF7BnFdpGEB2+Hbx7tiYLka
L+qZh+4KSiG48WiS+UTZN3+28HZQ5U/nFeQXBWnEuxuNHVCnaMd0Qf1CrpD9R3Mv
t9PURq0pBe3eW9JDrwinIFIrmoak2JjsMRjTjvxsIy3+g7kJRc33z4rRNwCI1XCO
DlEKRHiiVmfjVu6ijvMsUmaxt6SiHOqyiCoZiWaDYcI+uOJX9cXwvn75EqpF7qXy
zgMJ4ldj7KLbvbQZelCjpBgvjzxQjReDfM6zpMZnoxSSd1A9SnnBPI6zyeDNUJr1
uGPFYdU3XvTKzoOnvv/E7RWtsfyTICNUYdEAUAqkQ6nKqXQ/IOuZ/aSW+bRRNO8m
NAfKPnPTVz8EHqnIuIBH/Ww1UKSEKZoSSBtpuqRtP+kP0eKxT/wOS0N3IK9evrZy
KkQWnNWf2iVUjruiQMS2odoH6nFglVFT00AkFYDnhNU5DgcQASS+1rTJI9vtISlO
F5XjL/mcFzJ118hfHAF6P7b4uxMauCgbIoOOTRc+i9EKxvzsdPmVA+nyrPn8Q5hi
/HiSPGq7mOsgyVuYZ/Ez0xVi+IZlSDoIqBBhbM4xdo9rN1qtpxcdsdPWRBZshMAR
I3gZcMIRBW0zIZzhfj/dJigRv6N4k3SgBlFSVmA/NwqxHVzCUNaJpGdzaeyyyFSd
5NFYhlOYx8nfIQ8MetOCjiOCNrTBeSlJqpKLgyqIleKVKXLtZTsa+jxqwmQVPgQ1
w0ixrmmosqf3o3mSDFANvtJe+CVPhblik1bQPjn2DowSl+ToL4QPXb+f/dWA/jmb
QW1GXf1BwFGcZIcwXM8DIAYvIxXqbkTUTZfiQXyV8W+yEmpI6YkOMSnd19UArUZO
v0wSPfKEOaH4KFH8FHWO6yRwNzdTu+h3oLfG69NsZM6te76bjiAF7GjaEV0qDFoz
uhAWUUZx+AAt0wtZniwgOQ7TfUkXjjzwgwGTSZKtzlmyTkx4AiH3CVw2TpZIK17H
aBJOk51qrbQWdCOoyQXaHhsvk1BIAmscspFMI8fK1RKk0d62n3DJ1WGpzXlGM9Ye
EoQLA0wget93ntCkVn6vzDwHTrLTEl3ZZ1nlgM5oD/E/Gg0Db/MCkbfI7oRjYqaJ
yCzj4nPMdq8pCnSEjs7P11KyvpWXRIXgiZ7kwcoMgzaiRZTUdCylF09XvlyrHrxL
bt1KKNuKiq9WJ58mC+p/0TJ7RyrhOjKB+N51QPBVEByPvrnXjAl7nGa2OH2Hqnhe
viV6V0KuMe7rJKowcdJnoPCvZOl4taBGJLpZrnopSjVEdnWCwpQXrZZyMprnAH57
OlbaPgO2oExHUh5oivOlgLs0BW9y8aK1mZcZ9YwLEmc4cQkiVt4NKZX+SAOSkiHz
GS9XHZQXy7xHcXv7wMzhMYbFMtdITDA2S2tsWlvOhCPmB2ogjxquxsUOjt2a/npe
3xTN3kBXvbMgXvWwIXeU+jzkVvnL+ZduxKZuglRq74k3cep1/0WYXoP6QdyuPqW/
gDsNT9JwbMkMdB05ol043x7mIheRk6zp671vSmVue/TO3YOqcLnDyfPBUR9pyNC2
+dNFydX9WrYsm8aYK+GE+BQ//1ZntCGr+m8qGcpAKHTpk2qnGdWDlVu1Al7hXXhl
xO/auYnzP+IJ6BSCV3Bne7NzUBz250YZn7AcOdBm9adKa8jnwVKzrgtvYzuhWfvf
DG7kvwSFESTiP2nprU3neV4J9UR/y0/xU29jmR7tbKoCerXgfZ43pyOhR4tGniAJ
vStYJNVQVrHCFjIO9itcYSD+HaDFtpAajABKftvWRwREzBe5YCmagpTsUDLmK7jt
2/10uB5jxmPwA62e6hWv872axDpN6ILD9/9ls5tHxE7UxdW+4OiJs4Hqjn2RvdLE
HWa9RIvkZLPMIzQLiJ3Hckj1eRLvSGFZX6FQ8zHqnOqlDrjioqYYVABF0meJk6ZG
FL68TwN9DSRpAdad625x/gOvUl+8+DSkJvhcewuowCK4vqvqHh6LNwLcREkLkQ8h
0HM7natjUXKVutxVPc3HdXrJ+nrQKJX9VySZZD4OR8f3nZzztXyGUPkgfTWn1TXf
jwR+QqiAaRJ5adKsX7LFalGDv3B5QN+RJlqwoxyFE9iMBU9tWJFqnmB89JJ8QB+z
hm0MTewDZKrmnBi+oxJHFKaF/YNjaY0T+1+zFyJMbRSR23wxr4/uWLe74SvHt1cB
Kfyc22fv4/O2ZDvlezoPzCAzHagEYnTAG8+mr1Ic+XkXkY9nPaRTzFsCjrVa2ig9
a9qsiVwemUM3n//hVBFNjd1+W3nG2GRIOvom6WtLUdP7ygmLqQk48Kx4JLGN9C14
g/ZDzM3v7/ZHjmddTftXWg87Lkn41DtvKSXGow7uq/pP68uiIQpddzvemnZVtsaN
+UtZTcU8SPLUJSAtMxZwXILFb2uMw1ZzyFUNxSH1RpsTokp9RxMr51FAt/4pAKzs
095u8qQM8CH3IVuIi5rXu4ERnG3UA5DcLLzo8F+Bu9s1FuqFHpYO/iAVRZm0Ffb8
etX8FMuxiFj4GKmBYjuMDI9FS/p8ywRe5LYQZzATlF5Y0Ti9TJ0JXd2DjpGcSsRL
NYz7ZbBkAvLq6Wmk3L37IOXyAlqnKvPxYiOzXc5K3EjH+MtvyuYc5pgJGNdeJKsy
QvWY33CTvpdS7MgNXjxVlKQsMXRxIHo9MJVor2eGVofY1l0ubL7pWH1gCrq+eiTw
dsdaBZPnIwJpPvkmaR5WUD15Y2Icb0/jGZ+QmfMlg2Ro8qJM+WynfNEH8fWYXDc6
RmXBNC5TbdUD7sDj71daAGAbDYLwa0PoCO8r67gC3Gnb+u41J5/1RsSsydxDGFlT
z+TGGk06I9n0JREgltOudBqQEvBruealQsy3yvVDKaZN/PlnBnH1Lu2KoEyH6C7W
woVFXiuulehFThvqezCKKvaFFLlES2P1tTR2boi8dIotBpXnE+TBiZ4diYkqTq8P
I8q56E0X0eJhlIaHN3yBtw2HKGfUaAjQyE9kTxProkkbOZEFz7kbJzUDlMwKbBVy
i+OaZbwOUGwNF9ReJjJUNbMcrb50/3MdHw3XGjob23JpA32otAb9Ko6oBEtvq6Yy
Qp0duvkTXhC87A1fpyEKFX2PG5Pxg2/fUmq6L10fwff/uzr0XLOed20t9WUXJTr0
JX9QjWIXj9faUddOn+0/Oi6oH2nkL6sFi2T1ds/7KIMiwkP9ZLjZXTnkQ0Y1BHYn
p5ej5E9t2reJKrwvEhvHFYQeM1kTFSrUiLSwajqUHsrFkQhLO6xwsU01jO/M5yzQ
l6Ua34i5SIW6a9c2N0YE2yyDSK4J2Zpaagqo+X6RPJoxR7tGkXQDIr4bfyEXJxBj
R6Wje54xZCtPFnaPPUYb9e/QS7jfLXoTFP6Zsg9QBQQR2MlYim746cCfzNRo8UZo
D4dmrPyHmta/8yvCs0BYEWx9K+QnbYjCEnBepP9WtPJRVGlqTPTxuU5KGLcBDYh9
zx5D0mvVLwn9vaVUSzc+axnHRLLI19N+z3LYnMDfXA7BWnguoF8/a6HiM+yzzUKH
JynF8hFIUjJPzjUONiUcwWDRq+RFYBdzaYFaJJWdLK9S1aiGeB+RPPX34G4mJyo+
hCGU7IaLFGxZxF02Qt+6G5hct3eX2K7Efy5Jx1eIng4POfz9eXb93N/mnjRhU4gn
KrzQfkFSDWOvHRSLfkBDhFMl4l9IfKOR7qP/KXZvPGFQB0x5ubiYW5aU19De/GIf
40MqFhqHPxlC2g1GGxuSsDgVWqiojnAc2ucu2vijmSpkNNn3zOCGDw90aZiz9e1a
V2W1obDdP6jocQc3/MK2LKLGwHngBGxfIw5GVTJj5zV8yuBuNW1ZRAkl6mLLickz
R4b0t3c21kgVYKNGAr1EUG+4UdKxaUaHxdkRPLk74nyZqw8OM6id/jrDFEOPy8f4
V619NlmM6xltNTj7e2LQA9WQRHdRj2EwjVKBcv47/l06lyAO5oDlFipLgO5YJTiT
kkOwabHrL66gZMuTNsa4vKNBtft7SzNUVmCfxtZF6Xx8w7Yn1JG9vezEGZtkxzGN
JxqjMBF2t9XIQvGDxKXQg4X6AHYEf5O+XFHXrjdy1fStHUcU3OMkVO0mgBfJrNjK
2Lf4+rpEiwKPF6MMCbCitodKJO0j1UuEe0mZMlV0tpYh3HvQ3lA6LTiO9apOWtxx
RTjzhnBY/xxbyTT7BgLRFlpZmMDqRjMxKPSYO4kLvHlwbZKAsCEiT+NAS+G2iPdZ
NX8rLRY3ESLJ6Vt0NzP/Ni7wcii96GUXbedu8F34I6wOoopfFdMKiOqOaaVJEMJL
7OSrU8knHyJxCit9Hx6km1iuZAkcA9F6Z5Zv0KmedLjNYzuFNUbf/6X1IQLIx1a0
4RixCidnGr3HTkWl4Nx0qwuxMCqzAfZW27sjBiKu0YL6SeozWTrho7D+KiXPsOu9
8XHbCSrK+dRHr3oMTuTGOrs5Cd6KxZngBhzxg6LeBTL3/GY1VcDV2yqJjxzvvhiS
D+c4FOqgHUrHvjM8OSzzBsAd8PKjh8/W7itBiNK2eUQ7zX//ZpAU7v9so0h3zxHe
wl9R9K5pI1/bJbyd3b7Ri/07YT7KI3pdFC2fgA8YASbFvTs2//nu+VDXi+QpwM26
vqyr1QptQdxCwLbR5/tkmLkdsxXXx0bOtyJM+m9GdWASpGlGECf73aBee+6PiQ1y
WySFL0fWdf/QN9pknRu65UgySrX7ktuueAVtb8rkgdzwHUnO8B1hPMnZr7lKsExD
KCjZPaVED19EOSAI0VehbeqavzlbVEvGllJejx+l++rInLzgp9OTEA/1O1p3afRX
Z1Y9mNuwkuMk5f0hRilmMjs6HmP2Octpfja34LbNgYDxUrUZFOJAA/fMBWnrBobl
+nEz8IMQ48TYTWjHcWCxPn8EYDqdDIVatS7/l4sF82M7FjtFE1Fg1KK2OWtTGqKU
QL8m8ua2IxyLrC+bj/Ztt4ovyZKhsxmKI3uqmTPQ1fQi3pv0PWQDH4eb6+/SnDZu
crxYLDXpHhw/OsZK/Kk/9VGPsHSumd2g34JDUUMFSzt2wGcKpDh4weXCP+dJAOEv
vrJO1hMsi5g85m8glD3glWhn6rh4nuNE7+Anmk9WsYo2zL6v+FFNRlQV74K/KbIl
T0j6bbKbq30Rl+8mTkxmH8HNzewaEUT2M0ZgF1Qhc6nFfyYPwUg7N47I2/Js5uQd
K6n38dOb1N62Q/hnVBtete5dsrKO55/cx2144gl6fJLPh2RcAEorbAiEC0E6L5si
3oDyUCEAGKyk5iot5pA/CPU2jdc6CKu16xwxzjnrPG1Nq8b1AKybnlbncsdmYm7V
gaSdpkWCVBvvJuYGpxbKMNbDVNM/JjYWvD2le25oDboGACSeYh9S4BnxaiVOMyNz
V8OlN5x98BupmEBDwLoKln/0VYlpPKNx4zmw2Le47hjFX/du1MTVXpYUBY1unlUU
NHHf/OyL/7K+o5WzOF8j0p1wF8gYf3I50BIuhbyDtmYO8cbiXlxELkjcJCHSc93V
J66vfEYgLcWK9TnomsU7OWpl3/y4yG7G1nLaRremmu8dWUlGYdfRNJe3aQCuG7Bx
mTuZ+JRcEoZ2j1GiBeIR/8U+pAvAX7jUCSzctueJpvrIZBdp80EmDG7X97oskPlW
F0qy9wk0VvtJJSW8wbTYqr0jcrxxRTvrzh0Cn9BJYVTg7aPGfFWP6UJZHalvD2IB
nD0UIbdACCQbRwIm1OAbcseYhzuj5ywL9QSwbuF2KdSLQHnz+STx+2LfcyqJmMYB
nT3v9GAyz6e3sL4IZHSvaBZn6Y+ze4KF8ln9bHXODlufduFIrgFOofuuRSBAR6Sp
t+/GGvIWRPbw85YRLaZyOwCD/57lVxPymkcZBzQbw6VFkYa5a22xiCNj/TLGirkG
km0X/GNSuFhfOwRV6QPWfKMOmfzxXujEkkS6JVWo4VXlL8+KFBjy9Z0lMDS7MR0h
85ndd2gRJzKOKOJbo9+8a5AKvJzH3yfskFfW5f3fRd/j8ssnEgwLOUTncBCGZOVa
L8P1MGA0KH3E+3Dtf/kGI4Fo5mHhLKg3VKeDpvNXklO2hSff2Lxgl0qJxNZNrDAA
ym8ieQP4z26mhSdTYwaKWeq8Oj/1YRd3IvcqSE6EZoXAkdGccech9IQjnnkru6Z4
Qn8xzKf8n11eY8LwVzWrqKHsCZKXLXni9hbbGgQXOKp+cfGPeovlGN6ngXcK8nBY
AO4PqqAYEF3LzZ+nFzDYOvo8c61C+UEKObhdzrs2xfynSj17zqBBQy8b3fiV8cVp
ewr6eKu5/6vPrkUEzj3SUzNtVJ/emIzAK/GUz/N3sfEqSylU7i+xYRdZ8HcRqwTy
CttuAS/56j45fOFzBarRkvAD+vuQSvmplSCpAJZJl6EFbGZIOhFW9v8NnBWRkhgT
BUG5UULhDExQyBsobdxzFnMNYp0/AIvCSiUC2ByfhHSebU+dZNqLfDnNKAnX5J+z
LL5fifmJd0Xf7wDAJ+zl8+BhLuzx3NLcZoQV1eiO53L8NbV5ewMseAxCCDNJpvoL
0LHgzWGC0LPMYt+PTZg56QwZWIoOkSu4Upxm7Yem+6wgpRxwSzMO2+tTwY55Hz9n
jGW7n4WyiZNxXRIRHt75iTHXMBY8AwlZbTIwnC2INPngELqJYJw4qJ868DfEkoKI
LvMKj0YmG2UKPYQypYU5Npddr0Pz625a+y4jCGOIgeQR24ls4LFpnKhWjnVCaEKF
dap1coaJUcob6ydcgCYL2fYrITyYUH1vlRTVO2yOnFUsMiapDLqADyVtPV56iYJG
90zDOp9p+YkHzDP/RbnCa+JsT2kVs2rI10xMNfy8cWqdz4CxsQ8ox+x1TxbSyaT3
+TGF4f0rPoLdyT8Os+l2VFiy8hCWSZCD48+Nl4w8n2efRerMn+hBo0Xoi+Qoqvt7
9aNDHo29V+RczA7ihJe6/T+AuzFB6jr1RGVAvhvHyBdstWIq+wgBLP9yQHU5qVee
WPxCTZqTTli+MhNjNBlngJGJK4uryJWTsvoCNYX4cb8eZ9pfU0+449AqG+2EF3EP
csttE/L8TwpPRoObAcPcJ+pLjgjs7R9ahRxJuC2+lM1mm4qtPjo7swUK9rZS6yie
Zz56QD0s6dkmUMWDC1ATuT032KF8vzuo1q/GuiX1fF3Jt7041Me8U6xGZQh3kd6i
VAeWCP+d+SKkWwOQBm8FmEHj0kM/H/WUBLuSwu/uHsHtNo9o+pvMqcjJCCkkFt5w
qv6mHYywiFzjN2W0A9NQY4+JsYbPR34RawHvuDFwXp0ut2fttbL3I+EX2HbcHzBm
PP3hIZAoCylHpv32KZ8QJzPzs8x7BDsktxUUcYWD92mKSQnHx3/FAShQLtB4T7ma
w+RwfD35T9AkF5ipF1wk9CubuuvI0GOX7kN6V4mN6UQwFLS5bajK5QOa+fVUtVMM
KLiQtARKujs4hS6NIRQoHST8EHw2rON+D9VP0SROo6/vSyx8uguKEpeAG+2mIkqB
b1MMeQibBbIQgxZqwyvhKcv/3yMXnd1a7XuRost6Y/JiLaGsqcQfdKt0DQ4f4l2t
PzmI1efHFBe2vLwLvDY/+fmHTOkJp/92BdkOEM7FNMN4U6ggOMAijYe3wr/dsgr9
D/OoV1VcsmJYjJQkY75B6n5aZvVGsb8OvFw9XN87MDz/CC2J0jrjKqY9wkA0JWXU
fuRne7qTgeRoSSvf/io+lEOaueU08ygnLBP3AJ3GVeKq+yBtd1FVWoDkB9Xur8ix
Yg/aQaJrcO3TVBPYSeakHKv4a6yJhnvhJzxstymdjX9bansAlfs/OvDxUhLD/Tdw
vsQ69HwJsR4pwDcrVZyQa0fD0YChTGMfJrgB9gJKxQ+UWgqU9jFiEfO9QtSzjhKO
cV0ZILMzxDzl12J6OLIBs/GfD5OlspO63DmBH25WvHshZtbHOaI+ji7/7+GncLua
vJ3KnCQp5ntqUx4pEcgSLJFYeSSP/rkeizAF377gMAKCQ1/Op7hEYfzqiGn9y6AO
/7rJmmhgv7OGDic5BSWoxlqjZd2Z2zMH1nmi2wBl9aNGMyefmtWYyzJqz4R2JPU3
QxLpiX+LC8lBoSpfnDwX9Ihdde2lMK0hTZHlyURq2SSFmGmjOHHk39BdcLdaEf4R
OJ9T2d7iGXBwTcyGkJ9B3Rg7VTfE12D+uVwE8Lb4HJbrelroU5wY85zMt6Je5de4
UpVaw0LeLAB26763OXXHUduIquTsb8nR1RaIB/oWDDbVoBEHC8Ny3u6u80+Lgg4d
Y2bl0gVOwYrQ0C4k28x6zpmei/VQOcBFRLheNHkHz4oeniVTWGa3h0mCmnRjRUaF
udy+lWvlIdKOUQxfvyPvCWuXDLgZNf6yz25PjIox/CRgq/qgwnBKRjCpJTrmXP19
U9Rdau9L5OFVD8iifxdQzQSsx4rqsykiTNA2MC+vdbfBGS4nnn+xfLYDFsBGDmNG
aP+xPmt0MXZ/AvObfZ7RawbsIwRwROoKqKPpxqq4lCc7AFtrjxm00uLHBlMyu0cs
MMf9FCM3z9zo3CJO8EPgCHjFrzgeSgHweL7yIPKQfI+0/zqZujxjb6QDBNGWffF0
4u3xtGXq5GMNFEKMc2JpZeQVoGaOZGJwFISsVHWlKRfjXdnjr+DCZfkVD1YJOk95
a3dE2ua+TXnnb9A/alqGtbMScJqclms7n4rTURWV0Rcwb12Flqun+eErU8GgMdIF
8E1JkFD86l05tI0OSEE+djFTANwEwX9ZE81YbSWlG+u4MdlFwaF6oWNEUKN6r6Ze
/Ae0l1OnVggRYaBpvi2EEqQHGmXdOiORMiikgG/MdiXsM+hYKhtOmDaIpLClaAbG
6LMBjHsgk+GLGT9nlCy+8O0f3U25/FhjPF2PSMv1SQNmbCiU7JzS4hPRpIyByYXO
WHQuu75+oEGmN4U5np1GNOfqYPpcYBPeaw/gEzaBQoN6+8ltlEJP93uoHbJCHwgu
mDTft4U+adjXWDy2cXnlBzQgbGwkF+zDv4VmAnY8mn0vp3jfozkpVzALagWTdDys
IEmmH2+eodCqW2nSbOZbOYRRkJ1XaOIPPB/wAFPlebv7iSdgrvgVmaSSrB6mwrOq
oW0rIXrgyRyl8CkXZNT5LC5AoIWXLSUESNaAO/ANvxxZ9/cUilXEKcBgN4JnY0z5
U33rP+JrQ3tT3AR3sM5D+wlyOZK+61AKli9bbqkEIwVerqoKP1jst2EfhCRq40vY
37rDswzuLki9MJMy2PRxgN1SmgLJZKF1CjicNJRWnvIZyFJFdjf7wpt36fH3UVHU
T1tiv5QXZH9uvsQU9ZlbipAH84awZrGtn8E3u7f0e/VPP0ohV0UvzfctQhJHnpjX
/cXV6aFRokVLCFJZRAizBMcKQq/fN656RRSTL/zE81pa+7ivnaCpxACR2EuE9QEq
COf6b2H6DvOQdNhvyHs83ugk6WGPI44VPXWgt4etxjiv5MlqWq01Uz0Ar1RhTJ6M
zwxE6tI96xeR+QD+T/arPeqMJgkuBVHHQJBMLP/g0LhyAPCOuXXO/YB013zSALLM
Q4bnJuyJ8Fv/7Ukgy4PYVJPM1RpeqRWiekYdGWIs2k419KUuIuSjXBeyFlzxDEsD
EhiqaZSl7s9X5cRbr+TCmgMejXjiYG/hWIlsIhnq0UGCtM95PKVQLdvlHH9TAJCM
3HScdjgt957L2Thlj54WeLuvf2HEwcn2jVNlwkm2e/MDShDfd17aTJHJubgpDeGb
BycZWjXuX1jhpQBpuEEjDD07Su720J/vrmLy7nvyYPB1LiB94khotOVDobWyZiV1
CmVY90aZUBT7q4o0F6nf35aGgm6r0Ovk3P0ObCQ5t0/tuT3R2tDNqhhIiN58kFEg
ah2j1tWNUHvJm0U07A9BbRIo6EhkfC78ydFdNvylepmk7z6k7VCqJi0ijojWt7pR
1iW+lOIaYN46exHYoht0cFAGVG2jXwyhQX6Lygv8lQa+hog1apnP4hVwV7AaFn41
reuC7A/Wc6tAeRKcjzbDI3tgbpGRrGGE8qbeWXoOT+AXfNpLMSrNe529j+2kEo8T
s4uBiSNrK895UQJ79PEbHlEKy31mtQMrCoRngjjkSr2Kyc2Xpr+85IQA2TZHIYVM
VN0b3Gi7BjWcI7KFnTWp+EzePpQ/8oZBhqIYbGg8Mw9eN9w2KXxD7mH9CNvpD7N3
6sZO3PfUS6cMGBy655QWZ1kCpYNpQumxPCDNjmtU0/n7HpIOwaxeqE1GKiGcIDw/
UY8oZy9gObQxxYvjB4qReEGFRlQHXmFzhmW2DRe/TBsYsdJriGcBJvHW106Uf529
pAg+Ks27WzVwjrKLMbQg3QdfgePNivLbbOuJdfn0nThCYMFzH4ODKW/AZQbIeagf
UtP8+sqoSKxSx1HedwkzBrLZFWcwx6xQ2kc2juqElLA2P4U+WgLW4XhQzetoH7DL
79fNXXUmHoE+55dVylYgHYQJywXXWUubTx63oOPENLVb89qITp4FvNNjrx+d/tb8
SJYHG0jg+2wftB7JfVLy9tVPrd1YtN14pfW2y/kV4XMiQiqfr7GltY7rnAU0OSWj
IdmWYxW/jIQ1ERoYLlRjrkEfUzxx2DkpeVsUHAfzlndSpVyEaofp3LsAAasgLYzY
9iyk/Mu68NTLrooG2buv8IFoUfouOsyBVxXq3rTERCtJRaEaRTZtYAbcuTYrmqfm
OkcccsBOpJco+KeeK8tUYwjYrmFg9DJ/1hc60T/UZWG038lhlulRo3Mr3vg5Wlyx
3Xu5ZuHn/z9eUfZq42DEi83LKmbmnVlFtuwER+QC2lucMkI3se1V15WeciK8pmiT
o6/2N+OXEYupSiLqqOWqyMJ5/zPm23XaAFnMv90mdDcPkG9DOi5AsNX2KH1/ApHK
YdKVUV5iy7+lwZQRjWu9ik5417pQKabQIAnE6OaN7FzoF34s+c5qQ7Dl4HZOjVWX
n3ioYe2TMW50Qvw2bNo26wOoGmozNE+iE9vlf1HQ/Gj0E69IXnbYkPME/1LY3Azi
l/3EfHQ7YxqgW9gl9pbaBK5Id3EYObCbF6gXTXrMn3uqgUfVhdlM7YcHU44mEJf0
kiVqGq1uv0gbngZ/LK5P7060dduV9yXV9qeCMb+zvLoAf+UdVaqr2lHqFcYv2KtH
6mAm7+Yk5KopSPAXq23JEq04vp4ngW4CXDqoBu9bax54H93xJlzSLC+cb1Q8c3H4
NaOuJxrpMSMMIGeje8tchsp+7ocftnFDFk2llVvvFL2DzOFHDTb3TsaiVe9efZev
G6M6pdKqalyal4dT8nCXv9sDINKoxgFfuGbR3XbKG9c+DfP30NTmb41hknfhVUat
TlzDxaum/b7LSkm3yNxwvSnNZkRHvtv0OHw+P1Koo0PuM9NYxqqWOx5jp3L0dBjO
LRcslagiPbISYBv5LKzOIe0F59sodLMduZH8npAp6IqF+IHleQ9uudhzhP5LkBYb
3EjM2R1S7GDePrmyMUHeD6drf3V2CgJilDsII4C9/gdzJ1fhaOgr5XvmAGqqfw+I
ANrkmzeTYh7rAlVpSBcpe7HdTGmb2lMcFnHEH5IMKHN3Yj3VJC56kFpXjdvbXOt0
8P7K45Gf6NCU30YLYoZjgsv5YB6dkEg3lJce3i+1Hvp8tF+j0x5sjCuLbju9h54/
/vrTBF+76jpCMQBZ0OXv99jit1zvE5zRtlgCs4yZRiPTd0JkTUp8KrIbft+W/nqB
f6T0FfIrnOQIQGpuJIYGKATOLWlz1MGvjtoR+gxLKjqbXv3j9/x35XGpWauz6Lo/
VVXzjyUCLNKsO4hPFXEX8hIwfkJbir9DESCqxBHy4vIZuCqhanMv2QtNDjZzBXE1
wWqe93NLc076pQeaFqcwpf/hNPpH7T0e/vANNVadog+BtWEWa2Z1W9HyklMXrrkM
iN95utSxtzXI+RrlUk0C6DHq0eSyfu1WLRztyu2pcoLsFEFC++uK/j00XttG/s+M
T3q5XiOhFMOBySMNiIpW+DPxIBR09NcG06njMJtNqsoI1k3rYLapK4JvaacIVK1h
LJXRUunFQXCXZvY3kB/nNY/AJhsDADQR7WpuX3ePpck47fL89NDeHpzNfv5prhmb
rOUIsL0/HBmB1bBjdwL3i4pNO6My3VZLSYiHN445sz1yNvlYrqLcoWHABzFyYfQZ
G9IcP4/SoU1JuJvYkCwlsIB/7jWDrJhlcqofoMh3l9ZAG0OLitBS9u8IU5ZdCcfT
VbvA0P8NKAgKIu46yC0tnVdm9xO/lwE76hPcu3W1euAfwRiWw+F4K8iHEh8Fd2OJ
uNz/ZHfjcdeGkRLDlK0StTZ8GBlMVVrQrGM0VkiQdGQNbQUhuIeiYei0jIm3H7Kp
MIykio6XU0thGOF8+qwgPHA3u5n+omHtCgHQto2i6Dmi+wFbkqtU5wfYYO45ujcR
wExS1w106e1INCkGnyF+zysadwL0P2cW5A9bKfZpPAw/65ZU5fxVWw3sC7vcUoAa
D0qPLcmpaaByosU+q8FORX98doiedK/98FTuuZLZITpLFx3a/4O2XNyJPOyDD5/R
tMA8wRiNDCAV+Xm32pmCBNrD6Gcm9gy5veoDkIv17ApqLwRGukX5HGTifa3quvH9
dzQklBRdjEkctLxAqoiq8lCnjj5f5oZQYuO/hTogwHP40YGZ5dj0aCD4I6UEUacM
CaQFjLHsWB/8MilYSF+osx50cr7RzFFMp9ZFJfVH8RfbiHcDC6nymbSpCj3HU/Hw
3yphbKiuB+2OL6mANfmYHzDR5tPrWb8CXCYgRtanoUjnm6OBvNZuHtnSWqt9UUBE
MGEk1GO/Rz4+1Yt8+nFeVBjQYY0aoJRcQz2Py/z2FHSpSqni5X7bjhuVzK6LQcEw
wCttrSWYV3PZ0nqNo+YbVHXKvHHiUMiQyzu9NWN5At4=
`protect END_PROTECTED
