`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK8c/ZhdP5lgY4y7MnRhVrNo1byLMmyeMsyyD7ujNsRV
SPWrVWu0i74EuIOg8LzYPJoRrO9FUz4EuoRdCL4uPN5WNpZE99/jka8vC1zL1KDy
uhyMvh/tb2fabMAWim8bOo224EFA6B0pZYCi56w49i+jWnrRpWf29VEEKzrnNos1
zLfpIdOciLR2IbmJhnnYC2Z4wcwvI6LqI26UpgvJcOpCi5AilHhaEacUjJPMuUE1
`protect END_PROTECTED
