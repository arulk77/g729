`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ab3t38y2wf5+qsH/48ktMDHnRSJisEOke6AT1Ol1HgOP7oAWSlo+VawtXQM31UJs
kd2HyG3w6hFSMA5WagfUEvXapPyjJwaGC4ffnS3fFxELYirw+G/qf4wWN4d0x1am
YS7AvGTKn18wZT031vF4sHrT3UiRVUIl9do/WUOkwLJw3HLjKMVUAlgja94zYqOc
wcZbtzXTb7SGPyHv0FFN5e/cMg/kJNgs3WEJnVDuERevuNk+RYF/4EFCEvNoKhjx
gwFTxrdo5zNSTZ5fsVKBfkuy9E45hSAbf/ZaQnY/qn42YEGcS/0eEDNV2KDsGvPd
MXLUWgCGzt7omUSRIQWxXOFAmF8Rdk6oES64j/DXsDrOT2sAKIBQy6j5qei0v2Ix
qjpjB8Go4HTmb70GY87/kNNgdV0NKKJRbH756nksYR0=
`protect END_PROTECTED
