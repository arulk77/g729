`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB2v2NEqdKykVYxGI26GVg2RAr0xWjiZmiQEHnyTnVOi
lH077IZrnOmnvIQF9i2xPIvTrHkg6G+cQfrAlRFBzPmQBpGqGPMmtGyoVRYOqP2E
b0Yf/H0BMsMRcAW+nnopk+oHpIc+Ai01LxNV53Xmk/WWOE3imFZWkKrRmJMu8gdo
uYaukN67Hr7HU+zVDB0h92K9GE/n+Xxwqq6F1GhEmjz0eV9KvLmqosduMArCJhU6
B8FQeonL1rVJtvcHwh1HIA==
`protect END_PROTECTED
