`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCKd48CKNIfcSlEQEHg4JkaN5O1Y7csPKuFhaUmwti+p
7MkFTI3NiYW6jgwcWI0QhHnbF5AP6mHn1WyTPa3Bbm5j5Qdu58molCCNwhwxRPgu
nqIJUB9cXcuMr/4/8ETxQLyvjpT6N5zGaAJ399rIUPRoyVT0B+bEG3HF6Owx023J
HXT8rykttgtcazq/V1sgdg==
`protect END_PROTECTED
