`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAuSELNAuQtBtxnNT+DiNdWKodXXaqyEycE5p3JZuOtP
mFzgH6Cd9fgpdCfaq1PuL3Ok1pQFwNBs1uLMjsqDuvFANBHLJSw+tpOjoKGKxK5Q
BZOThEgSOGQQGftqTJdJISnJrDLLIFzpCIA1beRMQr39fp+bJRdijSfk4NqMXIgc
1MlAsj5IlDt9p+P6n7Pk3w==
`protect END_PROTECTED
