`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJY5hjFnUC71lqaaGxHz3qDWzDGH9EStmWpdiJuVN0dC
0qIWf9iVIdO7BqFVz5DIFHZ+Eo2rB9BTBgA7Wce+jC/vKnu2o9IjihtfODu+qr6n
puQzj/+g015xdrWTMH3gCT8axpbZWaR+vG0tVrkn0O5CRIUjhH2czwGIYzoyHxMt
7G0ox2uqztKm2MGUjzJz5VYrzE3KUqyE/5m+Pe8+YQGlkrNu83xWMT/CZziS8/v8
SGjDP2ld5LOarPawipZJh8amYESd08P/AFQ0+rCHYkiD20goPXScvycpWbenc1qD
Nzu6ms0lb/ZjiUSGnqn/zvwPPz1UTOGDI3AWsYgkrpldnu5oHngt66LqAVAKzUj/
oRP9Q+wnJ2PTrf/Fz9C2cqm7rgZ24uCqJoywVta6YoQqNdfXEzRRIm25baCoeWoU
NKdMaPu0mWUWtbIwpMzGcqBLy3j5ypb7npdZ7RYEjqrUfJWyri/rTWcOzEWlZjwz
mg3G4MrHT0Hoz4gZr2vwNzX5OkpA2XfvWK3tP5d/ib+Wc98EUyGcVrGVtrNYx/1Q
D061nWjutp1+xBr2or6IkfNYdOmntXEhkpB8g4WUcnxReyEH28FN74DG3FXc/P7V
1dAXbgYC94B6Ek9/JrgLyWo2RS/pVCfsBYySZxC/TUR1B1xfpIXwNX8BtBMLmbf1
r7gIU8eMHEuqQytz8XxalOpy4uIK7VBwCsNlKU1eFmbPXlotn3ShN/ByYqmS+8iX
CmdxMr0bZF++3lM5H28LArGjEYNC2l9GRju7Ffhn278XE808Xa8Sc1YDqjT3Dl1N
SMo6U/gkeOZMO+dAKONpML+PUJQqNHsohDVSopZgAtduswJGu0UjFKgo464bBMmd
zUjSLN5ChgbEm7WbPAzG7y2jMPphX/DFgRFFqUB3OonjtIguXnVQVbxS51PKYtXr
UzMobTtbulM+xvDXNRf4kz+RT1xCw9tSO5t30EqEcCnfBiBdAcZ91Kp/WLBk6STB
2LGFFdLEL4Tzlm6r/9caFaWw4faX+q1ffCfHGBMhkQ3PAmRpZHNBeMBDquO8JtaZ
bAm91V1YDotzMKFyQvKQCko5G6lRD60AfaTw464d0ODUPgHWMfB9vDRwOsZ3ECai
+HDOk3CiGNSMZkwTpKmEgSqPXHhN0Ww02SO6q8M/hJZ7/blEHVYH5ioSZeO5gFYp
aRkHCTUsGIsd0s4CjfqO4nQZS3RAhmXEOj+MB1NS/Ru1Q2xZdLkOZ1ZcHcNCmyTS
86D1EwC3kEDTDLI6yFjkSGjLU6ElvQz3UtfVfQ3s4phen3F9ifVelWxSiluGvK/D
b+qMAd0DXU5ATRT9iPm95tyfL/tnwKDSHRA/QVXiGUtnidpIpUapQyllpDUCbARj
w7lrHDj/bM0pUMH1fs7A9E+4lzU3xLjsaVTfOUbkUsnhLGwOdnMY91IYvTtLv1LP
hmrnb6/6EeRj5dZhf/C8IQ3hqMpi6vJ/FJqGCpe4RwIb+doU6HBJKrSB4F/OkYm0
z7EWAnT9NeIKih1nUx8p4Sobr5B0P81ms2WlqNJlTlvYT1ASrQHJicLMT77m5a//
aBkSNh2dJ9WrHsXVltp7sAFOPP6BkoZh5ktbFd3Fn7JDKdYok0S1Qeb2XulTMhO3
B/lzCB3Wp5/frJ74X62hMg==
`protect END_PROTECTED
