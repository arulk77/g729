`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIUzkULtwJRUNuyV0hCChxwbKkUWRsmtqi5tj8npdf0x
vVaQ5vac2EGV1QFC1Seyw4+XUJjmGr+G4Ln3fSCLt8899MU5mhHCSdjNWQAGrBEd
aADwyUfNDrla9tv5xaPLhOs1D0ERRgnRxNdNHFIUoaRKWZSwl8oJMfVdceX3bmtR
44olG4sHiwbKWL+cA8CA09lkdhczUnkkcxB1qURdzBvxhixlyArDakrbZsO13FRh
vuCpi/ISmEeNyFpB1/uDfhBcdrrR4oBCNJWbZaR+YEDcp3/4/90SEjDiPTeIJUh3
DYgeTDOnbsIpoGBzQPueA6hNLMKgjZ+fB9zBLXhr+9VmV2OkHYFcRq2N+fmmHtXf
b9I2km2LLoJw8m7/ctfKTSHjidXJzDNNibFSLV9A7Dr41gNqbWUrNVVpMwQjwOt1
uWv1ct/WFA9IQLAsHmgy2ABowI9VprZLJ8Zsj0LsGafCnWJG5c9m06Ic9cymuITM
OufMYOgdCGUL4X2AV9tbCNyRjXHDUKrttNkBoXwXQMLB915I3JbW5DgLTIuEYMZY
EtCPJ1dk2alrR0JjZcedErVGdsA1bb6Km2rYczTUGGp8Ky/DJWkswrf2mheItN/1
cvCndfX04si1F9m5Eh9l3lnuj/EKz93c8sANWbQr4407XZ/ItZbUXs2bJBMvgvCe
`protect END_PROTECTED
