`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOVKbVx7tRt4eHfCz5JawEKIX2agqWHccESPlxsY/T+5
Lg2f3qYEN1Fz6Ck+ZX9NhZOqDzghhHDNYvvGIYOQlHUiT3YtM6slRvk6EAqimAh1
efOTw8R+nHkcbnPqddG6p8t0W8wfoUGeddw0igehZAtIaLHvS2lMref8ECH7yw5r
5GuFRJS0AQ6zfMfHJ0jNio46sfTIQPiFvj2hhwBwxQatByKS11u3WLydIVJrpZgs
aGo2CNMfwjiPS3hMVbqs0g==
`protect END_PROTECTED
