`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLDQaV9/eWoGkefZpkYvQGkCHGn8OpSjNd4JwaHU8SmN
FpDlEcq21cKIcNSmT6kHtWVFYefwZH/566+Wc9MftvBAS3LepXkQEZm149tLdSdy
JsyCYg3Iyz1UbG7WXqx3zsu4u/kVNPtu3L0N8VL1Bt07zyUIBEs/9zLWAGYh3mdL
7AK5QNfCyj4DsdpVBV4bg+BbLewlP6cX9JLpu8zNP0YB5VHt0wc1CgORBMieMK5Z
zSU8WOu040qlO5CS8GKwhSHcUgKgVfpMUHQeN+V4VxE0Am372vcbwNByJPnEECXS
NdM6zjqLdmMiXWMHejbLYNiNFRpvQ8zT4K+k86Yx/MD1CNB3JuC0rkSOFsHlFBLm
8uHyW5PXhksRpyxZpTgG10cdnf48cF20jHXJlp6j64kzP30Sc8j0G/OS75ZclAcx
HhmaqGCVE9EyQlxxBdwiqu7Q45JL4k2QsKubdoPvVLTn3hRSmtIRhgYdIpnCMm2Q
+BHOuof8FIPA8lNhjLw2GBdcwN6xIENJnq9BZfSgVIA24RpeZcM7CEbfkRZel7fI
trgY4cYZFzzfW6ZgPOnfGw==
`protect END_PROTECTED
