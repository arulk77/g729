`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
DBr92OAmfnUqwgPqX67nTWmVbgn1jBG7FIHC1yj5ZdwuDBx1f58Etop2/MWDuNBm
iLtYmSM0QoBbiQuC7o18wYMpFA+wCuOqdvE9c0B4Wy0RoAj54TwdAGxLHcnftiGO
xs9Ut3YrW8jWq0AJpi3bI7x2EzRftOLcLzR3ASC9uQsNPjbwfQhDvSHNbE4CF3h/
Y+Iereec4nJZUjiOlwwKmUEO8UqsVwEUoWQvXC6hIwvqYSubD+qFZQtNw74un+wh
lLK3q1v06ppUBLDGnwv0ssONt630exN7T0fYlbk5sAbadTwOw+EF5y7kF4OmSSmm
7yEo2OyrJmG9SFwj3HTzBO2P3PCc/LBYTzcoWHyfbrQ=
`protect END_PROTECTED
