`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNbLR8zOtf3P7I7jXaM+BnNgRK01eJr5jW4TZp46FiD4
FaOIB6TqQhyJTGIyNB26CxpaPHDd2jkmioKEXaFKOC+CelxEiKKBTvvn/FlJnA1X
c8Guwc2oCtwiHtzvArKyoSybVRXPc2ICPLhSLOhAZ4n9QNCfJ6pdl7YspFnV0zf6
`protect END_PROTECTED
