`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHzbJxMm+0dhVMy1l/kxMIU+MWVo7qdrnjxpv90aVGMF
SfTXVciwZDHtyI+ksueNvhkvDMqaIzduFdg/qepOwFSqcMjyTeqEsRXyI1SW+dww
DmljY3BejnMVcSYlkCiK6EGh2XwNQ3x9iwtvocwxQHDX3kzjOVsU5tcitqCnY2id
VcA4udwpI9LmdkCbFjn6ba8fv0lr3CYrum+uI3Pe/kiOp+tlZ/RJGteM7T0Rc5am
Howhn7iuWb76mkFX/MPvEnXQeK7iObhhNE6hzoV+CYLn97TOGKpZkIgV/XlMWMhW
uvSKFbd5Z9ueMH3wqDl7TnZ0IMKl9lKHfQx9s0SYICTww96AECCYAtHO4a1lFHiS
W32qWuI/IgbrV0AozrKkHcwjTo9eEQ9ywHgJvBJMb6/kKs54tDrHgBM74wT/OJma
Qhd5K+44EUtjTpbaprRKjxfCoXtkgPr0PD06VIy+rwNKd/2psYXBlNMNa207eURE
wWuFqFjJXtgf3vFwNSbS2THb4B4UfKxAxFYzzAmC7IRypRLGZvr4gZW8nwwC5XN3
`protect END_PROTECTED
