`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNy3DQm2dN8McPejn+c4BOyO6Anbp3N7oQVji7yr5lbgZ
6+yu1yPksBLWeOLu26czdqodE0BzIqyKYja6TboJq2Jpl0G9ouxdi3WGw3CiyWuP
BfRk4Sm5jAeCRZeJI9C7LjdtdDL+Z0ObLm9VkWOfWK78fdgCJnYRod9N52ZS2zVd
kb1VnMFne3EJYQtrTAvCvexmozh3l5seoVNYBHPKWoJQDKvR3T3bEon29TckcUD8
Ht+cOpMhELNFa/fdrKlyBiKhIZKeTiGYsTWhsdxjpKNNqboJ98isuIr+7xMdzliQ
pZ7PMqMhuva5+Qf/CUIDXfoVTZSay0w4R+CdpMhZjLQ4dJB+ih94Ba97gsUcettn
GIdL+maOpnOBSNxM8Cpt6iMEiBHLCC1hiJ8zEdU+cuVleV/2GylPK8Eel7YMue3M
I9A+Qp3nPQAQaWSstaIYhZEeHa0SAQITgBH9dBcnafXIB4MvcsZiOd9jvjZ/tg24
Z5PHtDbBWnXSTITYbLfpKxTwGBBfFbrQGu50Cdy1HJ9XrO8hnN3K+2Ewn1SSlTeP
BWCvZyObzadfkfmHrdglLZCz9arC7JUksFFIKZL8pr9+6KgMYuFyicbAvd2pnt6v
tKhJQa1egxTUtB9LkKrPehuBG496f8+p2kSM8HlIvr3LkctMSTGlV6KV+iAYcLbH
HNUViKtL6VkQNDC9/oM3qcF9XjbKYmlb2tVOTga5qdhNqEilF+7uYmzpYyVsbOzc
zGCGaWvtsAWJeVjpfuclu5Ic+Mu8lEHhqLiqapkKCd47HLBkTsvSpr6Gvl6sfEDK
FmSBPQDeYCzQAER+L+3OZkldf5W8cAQPXhudMR8nqAOiJtwZdYt04uxG/qYNVe7C
Ek/YW1rZTGvWnqzdRiIT9FaFAMRjN/StkDJUyWMSubcww4njxdUY7DmqF11vrtpL
HPUruJhChfH9Ut3YaikYHBNuHZF7tC7keSgeMa7BW7ikYZrU7l2xruUQ05qB97yB
W3wg97wdJRV6vz9+mugOmw0Mrf1h3CND68vLCXGNh7YiXLebuUZWwAhXOdBOBeA9
ZlbWBrIPZ0vxvoa3XrGKThZxmtAqnxaBqcN2fSLk7BuxCDdpZtJcZzUdYhBgh5qs
rzT9ztArV+C0OxHZ7eIRLq4bQ4rrohQJwxdJjdBs5Nt36NN7G0i/mXMYx8Rur5/B
4uh8tOjuKq1rdIALgW3KJ+cEhSLVxfFgCx36wLaoLhTNHDupfdjrp9CVGE1EpdLs
PGQQd/2loQ8+n5s2IlP4RwMQgYIgUjfvwTuHpuJpEgvBCqvdjBoZwzz90sJCwrhj
/m90XQ3t8GiySrijqb+j0FvTXuJ4LSvSUWvrGHtdCa6PzfPwfKStzL3p0dayX4kc
dNgplnkQFjNb7TyUyg19lwQkG2r1FnZIQrawfor+yqB+rZVPwbBZPPH45Q5aPczv
1Gkbk63J+sGw3k5dD85hB3SQ5xV3mYrpliTV0UN9byYyGHpf2yg9qX/7UyxM2Mh+
9VkQYafuV/CO58mOQ/I6TOYCcAed4HuKx/Kv33ugX5uL+F7dhixUap3tEpZibZ9r
t3vefAy5U2Rp9a1h5w0tBJqB45GYZx4wkpqV9nRSN6e+K51I6SYcLKP6sGBaSyFt
oQ3UM17+2EiTj2DBkzZr2ZvAQdpynw35ocg5kIkcA8ssdAPuE9MlcalZ9cQq+ptf
RGZQBlA4Xah/FRUJxgXJcKZxcvCXdA1MUBbNTkw3wEErGMrCijhTCi+7BJ2nC/GY
5R+HKPitcYvfmb5jqV2JQO3sgkEdaq1YlNjUpTkIpJAI73kaKt8xxDLqiNa9eyJz
vREpunzAy21FMSPLAehdRdbfGdxtQTnK27LmaHiiWNo6blO8Eglm+O/SgTBmPzH/
ijY+fyExsTdG/ma5vOouqABelrSqh0rY7cCCTRO+5TwU042uDj7hDELKenldVqJh
hBR9TmaA+XnNXnpQj5GdKY1nQGOazgFDvn2ssD4YRt+5P2e8y/FGSN9eo5xY/IV7
e8wk/DpZFHzfoReReOcb/Ky+BcYhFwZe/tlsh8pwoYCI8u+nvN/g6opt9hOC4/nV
PN8CQLd3bL0MVwrM2oNbiFiVmso61qdkjnNWkihddrhFgbEd0m2ncfomUOzRQpLa
ojJlRd0rze0P5AGPZnBETQWMEHOhhA/1y8ccULil0tNOqHKQHaNc5bL9YENXx/80
ilXhXz0TFtAGIM7YqJBOGgLYFLwQdGFOj0KXDh/CvuZvARPtVo2JZDiFUSAUJria
Hzzj2X8o0JmqSdeoLIzQT/81XBAMjZial0XXnKa2Epp1psMgDT1gPipIfzKWwsoM
4JaKv2WE/KtbhkZKVK5KBUJJI9Z6jTox/rQkpqg6RLEyZY32u8UYJfa9xPbzdA9h
S4R1PAmOWomNl3cGyrN73sbdq5XqgWZWODpHm3T7BOuUBIHeflHU6LPiir8CwzIr
uNVntRbxSfeSk0hPLe7Bg2kwRjaJRCMQ6qdox6nN5Kg9/mHLtxjt/2aIt+P3LAmB
Jg8jVuchgDmB24kWP4xnjxxBGme6oaQISrng0sJ9ER2MlXzneDMgv4dwvgwQl5TG
IbroDr20dVZCglL3Iht/9wZGeFG9RVmqR1RhP+t1qsxToyEhHwsqIUv4nJO8mvmV
anU03RCDJMOGSzkZZYzyeIPQ24qSAVX7YYm5g/8qYLetxyFbnJOJ7CW1PZHFAgUy
pON883QaJFF78SIq0RxzjUyhXwsOJOzAbnbxUNwJks/fk//WlqcgaZG671fNq1n7
S91c9U8nwC/W5SkcDEkS8kZ0z+jEi4l4xuXZ5qMVEciCFyn6SIyZbrExxeUVtCnd
eBujbaN+jHxLAUu5gDSC7jWORNTG8FFP8ZnwLXDwoxVKkW7xnn9qHOoXuV9i4g6C
1Ut7gIDsOE/E6scaskOUlKh9JORBbS1k7oznD/Jj9Askba+tVP9UnFYS8T3xjQyP
aFIjU198Y/yvFcraKHGtMAbS0sF1R0cmX+vXVJI77BI8pCN0Ug7RBeBKY28o6VN6
XcFQqGq5crRxSa6xLSijtslV7tUJdmQG28XPFszGnniYEGm6LyETuQgNWw16h2nD
QvnyAgNjPO7loXNO04UZZkKhKcfaWAKhw5EwIuoS4EIX2jH0x0UI1RQx0ZujSwJW
uVKCMKu81OGeNx62Tcd4zCGakj3N0qbQmvt1XAWIRy+LmpTSABzO/B+11v2ijuP4
w2GBpbNpQNiAkK49Xk0lieFTf9+zrpBhcQycvwTLeQwPuFkkd3ojo42EbJpbd5Ii
w7oj13krw3Qwi/5f6WyiFofO9gOjGB6jnhtK+Dkrv1w37vYxMOFFsB4CekpA2rUY
ITbVuC9O0R3hcMSE71a+z3ZSssfVyspOGHff+UiW2Q2h37fJIRhaEk0pD4/6Zjdb
kuKmqTPHyIrAX6KOWimLsx9GiMV7yAO3MjAxkTLZOeHFAo6/vWPEXJapuIef684c
DcCSZ+Z3J6PO5JNSl5YpXisy7R3DupxkKxlz0rKoP0XU9sfwyxCgZzpgU7G3QHPV
2L+ufxw2Fmvuvk3JwRv5HjbuuDCB1oyUMRIhLRxkBbJU81Ut8/FFw11z9fVsJN5t
tB3k8UzgPFaYXqmmAxmlg/AEtRn7kmlcuCiBGyTXbd6vL/IFKqICV1q8IVUfCW0Z
f5WylzhsF1Il9wOxscXkbbMkQuAX9218jHY79Hu9Q9af2klzf6LL99qkibSTYwqh
BIQzmyzj9m9/3emo6nXLinTxBSVuCYuPoRjiBAwsL03pSnJ9KJjLHa+AHqv17Z6n
ljCxKrcsGxNJHV5mBF7IOePVyEuBEpFknW0nKT4d723UspfG7eLtQ1luPOGEy4Qb
KZUVVKHqtDgtJ3SAJXZwCIHWtEsNW3o0Udz4h/Ub3lH+D7fvp8Q/hSxRiNY05Nxv
UsSQrWICk1ChkZyMNdprktfePiYUySAZT5wXae+ZQ0cxJAiIfbdDcSSnIjGLKHOg
i9tjC5eXAXtUddG6AHqgokFsRBUScXcndx/glcOrIXhMVU2aM3zK8XkGs4lyvsN3
tS8ygplOwDjKu9bSeAQQcIS4+T1MO6ORA6H4ywjAL5/0afVQQGd8k2k+vpb7EOZR
UQZguz6YrvVa/m0Tdo6jfA==
`protect END_PROTECTED
