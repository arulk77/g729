`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCe/fsSyuueHD+YDElgYVXqhoiYCZQWHjaQjHtXjhX92
aO08kK0gj78pYPZYTFuOnFLoLlzlCLCtHKqCWPnj/60INPO2NmViCiAB/d7gBJcg
L71Pz5zzbAnmlRZOUwB0nszkU4JlYE26NyKeaJpq9bGejvyEsXvyp9oPPce3FSuy
ewpnJ1TcR+Z+bD09Dd+aYsKgvtA7QctXAu9/dKxWch6DvPXDiUz2MPVfiTbaYol8
aFyRfdbLH2xWk7iJeBZMm3fjQwnbFRCBDJu2A3geoh6xR6Hk7k6GKhhrZUVpnpiO
o0izCZzhiQc1O80WDafafoc8TX9W3XpG+qssH+XiXqnzegSgAqmapXCcK1zI4hiC
HDQH3EpQSpEOYaHGG5PUqmGI5MAx22cyJg4RXWU91XZvsa1SDvP9J/njUiQ9nUCM
1VKoinX8TtRU6yF4PfgbgBCBXxxDp6IWeLAzaIX5ZuUcPdU+cxbbRfLJLbkdjFKK
EpzZDRAH2oOuDnSGFTyZF3fBKS9SZ+LVAGSTONstwg6IfaiwOfs0euIs7Q7vrDou
6F5zXfjbMtlPxHHUZqnyoIUcQknDldzJhQ50yAZgF2R2oPTKjL6ZhHFaaXDD7f+F
f413zehWAXmKsSlBAgPAn33fiHNXiG2LJJHI8tsRlpqcRpqYvCRbw85yLeGOMnMZ
LGllvMvUonudANEvkmN27pnOscuYJsmuk9LjBpaPJ9wUpNQHNG8bQ8PHbObgyQVp
w5e9EkmqBXUArYUUOp1ko+cYr+eZV0fKtFfYViIkx0+hsq4uVwkM5BJ3g4O013Ok
BicnQUqm5h75Ak+8vYFt9XsIJ/fZAKtnn1DF0SIiX94=
`protect END_PROTECTED
