`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOCladCLzoeLZ64kOxd6uCS9iUgYYVlXqm/s2hs/sVmc
2K72FkPmsBXebhHNF05733N1CNQN37xo06iXsuecwI8CjxD02WehCjlXK9at1CtY
MhB37QSOfgIKMn4i1Q5qlPsA7dxdtDoCRMjce+ABGALCXotRUUjF3HdrNSSuRPwO
pQy7Ft3G4I1/lXcqfRKWbPK3Cq3Yo9pPrdc8cy/V1fiYea9KmYJK9VleNuZPt1+Q
`protect END_PROTECTED
