`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePvF3yZxM1GojP6nzzX2IsJnKB7VVuVAOIuieZcaeiDN
IYV/Df5i7OJ4Qdm6K0xS137iWhrWqWKZv9/chol4fFdfDOX79l19yDigW3gWVRjh
AizDFNhgY7oCDkiumpnQtoQ/OW1R7ZvXIFYEpUEbG5JK3XY4wi90BTm5weqlHCK0
DlVVPVW+ogW38ZsRUyClGQSjfJv1OvUEN89pbcvlNfPUxFfOdvEwnyywBsAQE7vB
4Jj7lBU3qPtScZS2dT1DBPtu7T3SmV/b5/j6Fz2s2eTEI+dsL2vUnhCI9F4/O8+Y
zxgomFX3T8AszhRsRQuSHS/hs0EmHXJ7YvveZNXF9XdpOlbOFitDPo97ZQ9PbIya
LYwAknVlBtwkoFciF5L1l/Jc3NyWtiC1LM/hxudfF07FQAq9ndO25leuxDpyLOuG
cxJ71cIEKA9QmBgWiJ6zt5JOxPFG739DZLqBDcF+k4HSN/MYYADBkFwi2CgrAeJn
TLszfy/W4zMHJY7+zLQfrA==
`protect END_PROTECTED
