`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLsa3z/NqOsGc5MTuYbZE9DCf04DftWjYJBti/CeKgjr
9IyRYQ4OZycNL7f0xuNLNRn8PYam/Ic7mxz4qCbstGIepggNfKXUG+z6QorEiLh3
fdYCp+fPNqJjRYcBY8eRqnIBx1wQd1tYXEpqyOkvQ0FfpiE5Ujj1/AgFmT4Qrp7+
qQG4MUIIuCLBFZQYhQpnXIHp4qhh5PgYBM4hxDgZa+To+yD2wv5JsivlsWAUajux
dJdqYiBKFdbfclEW3UQkk2jIsHRnmStibyvIbpYf5A6/p+mhajV9eUOvjeQoIhtr
wdveXtS54LC0PAFEwtoUaSZi+8a+/Dw1VAmlqe+XsX16VCGKuHY1iFw2jp26+VEF
4mHlUKHZXJr5MmF4em5HWWECyMQACN1YUngUMY5K8wDD3i5PA+lHq2AE76gRKTrz
byxIo7fQfV2U5bSTAfQx+8qIhzVfi6jxrlSTkDP2gDpGOgypMuLWLSHiVmAuipKU
rS40+L/ovWyULs/A1hsX4fD1G3ddK817k+mY1nXWulv6fx39u0Fjv8PM5wmoBD5L
m/sb/70wW5QY3au+/Kw+PuV7oR8oE9F39VyTVdQOnFU=
`protect END_PROTECTED
