`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJQQtewkt2vuaQWneoT0FvZwIgVtTvTnQIgGpSzf9uaf
vyeZLir/EkhULgrORSfHOQHrfAXvwCc5i6qLlJaDX1Iec3Wb9TWo572TZNSsgyuG
8b05QFVBrwgXaGYg8ayb0PsVuphdASL7puDRs88P6nmEed4di/REBC6dr+xB9cOs
tyyTii30UUnX2vvNToCj/+AxgOkPKD8pKv2LhvUb7EGZEx4qqmpAHRbjR4frYo4v
imzZn2Q2U6Vx5/rsvE3N4pDnxF2DlZaZslaSe8+ucjU81hv6fhy/fYY7vH2PMamu
3yS0/XukoIoQAlQnmqDG/WDZK83ITiUpl17b0rRtRvzh00j1gzAYjPl3t8eDhHqW
ti3sKTIVOcb3GJuTTu3tSw==
`protect END_PROTECTED
