`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
76sFkWaWtW2g4TUTKwVVqmTLS/2OF/E6oycfb/RRWJnoPccFJyuTWFuZJ5yi3QjQ
NtSz5wbULbUGdyXNx7VuW7kdovTGp5DdtzF0hzumT14TZh6AfCKEMpJZUQfF452u
fKvDekX0GvkHpcWbbtuoHFcmRwLBu2fHdpdavLbnKoh/njlF8al1o7NKwX1Mzs+W
OT51RPLp+7l9MtpeLCH6BjPEJBRTIxoorB8KRsLfCQIlW8dPMkZz8t7VkWpFcbrl
ke1Myxi4DGoKGzztptmso26UtYTO3q2So/MNpJUn5gywduDrEIR+FZQojR9nWpkN
QkKipX/+eiehpX0qyWcNxYSDZSqFJeW6H4pRDIvYGjA=
`protect END_PROTECTED
