`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41Y9SdV6sLou9zhQkrC7rSkUI5tCG5okWwCnR7IY+Lda
3IhtcsUxEmS0NpRIEsk7lbcNQH3ZRpmLgCvKsXChrKD9G7svXk5nY8wAUVW4sDQ0
dAbrvk+w+J41Y/VAzFsYLxo8p7wgj8RBnDWt56dHKUvwlQnvbalf8pZMq1FQ6m7G
eRBK2cnUnOp+a5yFMUTte8U16w0PhLALlnxWRZZKvTJRlMxiyphQV4VgcjnIAuDt
DktsWcSPPWk5LoMXC3HTrEGv4K6XOyDepCJecgNeYqrwwJ/SKcHxacmgrQ5/evPO
P6IS0KWM50vNcpw3rjiWEYkDkhqN7IRo1+o/Xp9XtIs/seYnJdEbxNwwc2z6OodW
txaFQMW5WTZrQVPrqNOCyg==
`protect END_PROTECTED
