`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
nuo1Dq5xCUgXgKxC4YBeG1hhpTbfxxLy2r8wC/mUjcu2UX/y8IrZGSDPhoLN4Vr7
oHRy7jBSuBDJrv2mQQcbWIJOfGGw7wNlXF/D/doiu7cRnSdwEsP2Tge5rxsLzxBc
9JNzBn5nahH3d0vJXUXFqwcFZFWnZD8wkH0oicR4qzieQDaBAgGlTJw+xc1CgCef
Rl2zj3jdFlSXRLMPfFOcM7mpQv6OiUTwRaSYtMDANdbEOeAcYYqC/tOQRn/z0cX4
LOkvL7JMZD8zOXAcElg6CLIdHjCIQC+IgUkUtwO2DCy+7MmenLmiKVZop79376Ue
5fUrkNH5Me9G0uxAYJHfpQjI1yZ1iOzlBBNPpfRkZY0=
`protect END_PROTECTED
