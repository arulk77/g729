`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
t96EF3ID0kqLzm42bgx4ngwghtL0VN9tfq9LYkR+9Az0HMyEu9uNjQwEHSdDh/aH
u27ToWUcBo5I1NgFYPRBlRmcGRucAZOtVO1AGB3ucVND7Qt5rYlOIqh7Iv0ATRGb
mGxIBOwozkzWsg/SZMJQaEKMZxTL9QZkE/Gi5lN0CFSmQAqmz7KmtNIYRZSOViIa
mkiG41E7nIQ1XVXzh0zRqYkJIxsOP7M0eIvRm3bAg9BwUDIjIP1XHcnPnyEMpoPo
Z5JLDj0uIA690c37KE/sXTcflvg2vvk1q2rySvgS7RHvkPrgyheZfr6tJ2fDDMJ3
QEy1HO723wurVKkis/rOseejiygrgv4NGDrVoR0E/amziTTJhS3L1WrV753rRr4P
cSTGK3gkfc5RdKxAzcCBQhE++b3lj5ooKdkQVLXBPubNsReUUz/S97SN5CgYmp9N
xiQ33z+KDrMl4BIf3HkRG8jf4H9RP3aVA5pfkJuusOVSvQG43YoZVuuyZ46w4YKx
Zzx5wIqTsopPAmCUr+Z0oCb9y8Mt74aJItvmJjVElICvrwWNRre2OqZIsEBIpgsA
gTBml4gjjPa5lcuZUb7meRj3rhlZ4BfB5W05qnIpjxyChA6eJmwEg4D501MoZeNg
Y/3WXoQxTDFp+MZi0dsV4Tp2BVXsC2J0WLHBY8TvE/Rwf/PYOQhQ9HbMivI9pSGK
wdzLLt53sqYekXCCUD+uH8dSVP9cgXyKeagN1rc12rQIWkF9Ls2NRlH2pnYNpQNj
3z0IBMIoNnKG8qIcHAntPw==
`protect END_PROTECTED
