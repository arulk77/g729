`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SRsEpS0vnJ3JP33jdzM1ygULNgDESGl7+W5lGDhD6/sa
Kp7tww85IaZVrt60KVS9eCCKU3i9D9MtbOacK/o5tXr2jrovl0CG8RNimjUGRnWm
MAaztRTyWz71Mqu/gYsw7oAJbYvFXmivig3wFHq+6EuXunJMyYsKkefD/ld0kzE9
jNpxj8N60G88O1SqByc23xHbIJCee4Ee0FC05Lq/b2Gmo7O3YJYPsEhqPMdXEPF/
wtEpnJljXrSEa44QKm+gpOv2LsSCoMpwyDbbov2Kw5I++wIQsAjy0OtQhp9/f7re
G54J8krRQBANhb7VeJ3IcZzm1c+cI771qeTWovzzTklkyGiN1bEFs+9WwxDnh0ff
XgYDOf3S61kMxLLbofRg8ygc/7HAErweQagYpNxg0+ioxHTsUYkWpqy6ZDQ3QrbL
hZ9s9jh7INL/3Ggmt1syXOtOpZfbj9tvnFp7cJ/ikA0XE9cbV3pAfiJ6dm4JhEkx
BHMh3E2dUMlc1kDfqfmhGS6VfiqWsiRQaqiEqUgasFq7ep3OSN6MbqKrL0QEokbm
KOJWZlqj9/4s4WZH74IYOnzok1aJHXrLcFWy2RB6noKeFrjRafT9IFj/vbDrnn1w
7VnfZNz3OIrtd97F9x0DeCc/zZQKe9a8Pn7SOkN4CqLaBQ4Iaj4dV2Gn/9USGqn2
XnVyy/H6llIPqXKBq5AgcOyMZ+7JxsYwKRCV49AVIeq7HAs2DsyJc6lWbRHApE9M
G2+kiklvdaqRTYY4inmuykAOAqasHel2pUgzGQ7X9gBC5qy+JhApJdZKxrbDhzse
S8mHRY2wIyI0KQrSIToUPAzD3jmHSTCEO03mcuQCpYoYf4/mDQ+iUdJ0gVpmAceL
UvuZwYVPBCF/JhVCbKNxcucq5ZwPOdNnFT1kkcUMRazEwpANxH6H1vpE+P9PRwTh
5r7Gah6mh51IiyirMJH0AhzFoYx7s+/G5hm6WGxNQWJM4k6bZUBrdPTT/3huZnhi
T/EeHM6ttCU5+O/tkXDSiz1yIUeiKo7SVBDEreqooDPppsXed3NUhhafBtQHhRz+
U7UW3KTId0/SN7zMKb1aFpvU1/d+DovaDp307p4Yt9p16YjcgaaMUAQtwpjxrwWC
iwE0KjO76gpTqPbugYbvBinqS+ywnwMRdGhPx4/4usUMFvHc0Mrcor8NbwvLY7ba
SJLseDe2Hl02Al5o71LjiAhWgnVEiLaoXykxwEpF2zfjwkMMEb9HzJWiKMfJamU5
IRgQGjUDnpTyU+vJaZ4fLUgOL9JxJxdQ8Sy+Yy62rZk0d9zRITxgDZn6xjDCbgrD
1L9g44sQ799YScRliSdE5tSMTnbsYK0vKQ9prxFB6R6zEsLyqQOCQg7/9XiTOV1W
nrx3F2K4oHSkoNefD62wRgUP2Nliuej/W7Tk8lX+Fzmglot4SXTwlXRGHYuMBnWl
FZWljlYZ4ZOI1Kxglv8bkZJp3U+TutBbV4DzxOrbRbSbuU8DO53ZxUY3SKX/KqH8
I6B3jffPY7pNfOB66jI0D+vgR7TpyLOoUtcScVyG4yiqfNCypgTI8XChEIKP4sHH
CTeNhCtP2H6rLuPm/kRbwyi84c95CQrMm+4QILc8C+XTfOX2C9rzL17pa74g80f3
RAJqZUQqyB5ICAqvaj+HJCbfLKwlO/tXIQPhQY+uSRTtMaKnHtoNsQj1Xn134CAE
6p6J/DSQMospUjNPrj68tQJSfhdSq0t5k8APtjGal59WWukI73ZGla6abd/23bdV
OHatwwM0OgAJXTVnZo1v4ui+u1deyBkr7nxhmG0X/5hRO3PbYfyUqk/tajCxG6+q
/4dqmxq/78xZuF3Zh5nr+/kn3zBxKtcCVjVbYHL/AWTHLDXQfd538nGkwGCqkD2n
GhLSXdFkNmJSVRrwvgq95mer6y6/Kt80Jf9bJ9eS5BoUYvXlycn84T7B+3yszEKD
2Xkj6i9DKlby0iAwXMsQ0vYIvHDGGHQKzOR/01720+qIL8Q4pgktKfcCpLbFenab
F0ddk9SBAiK5VAjS7HKY9yOT0vGn6rfI98CoMZTLIefoqwKeR1ahCzxkJhqcgc3c
1foeeCDFBu4a5MOzU4bWvpnOpDLh1CWK/f8HZbuwE+Xnji9TWEEguMlIvZ2AYhOB
8uyyomCKiLJ9R1Rv/sEPS/C9o4PyQY5dYeqUtTgaJkUiviKKsnSeIPupwg49NaGh
d3YL2/GNgFjKhvoidEZVFTtr4q0vdxF/oCb1rCGP0CKSaqIKaVIqX7BN7IrVR7Fo
VzEhGs8QwazcJkh3yTLfqaJ/uajII8lWa64WEJ6BaEdb8hCJUxiw2gv5NlXwfSxg
jMVnpbFaqfNK/HkQb4cjm4zRMDILp/nNyrD0kZroafdt4nK7Cj1BmFnjHhYFFYMF
YSHhDHtbuCFPdu2y7CQ2N5Fws3O3HX4pSgV12Bx20TxuUSZYKzrmmlHfIkET64eb
OwsCqe3NjUth7CNSso99dAP8j4ChdKk+4prz+/rsm+oQwnGnJxjOdr/YyX5K/91f
IwZoFOaSRRbAW7RpHRWZwI5erRwMWtjQ7R24QiRAprW0eSUBc3nwUv8rv8h6Y5lZ
QzDbrLnX67OevwT34ez18t2XmFJqIkHPrl82+9Y/RL78pN7mAwjhmMWRUHgU1ZSS
pdqJXwedsPcAkqV+gpwUk4jD277nX9shvqoHOjH6tUmKpAfhaVKtdEE8cT0K9r80
dGDvy0DYebkny7N0SAELHDt/EQ+OvF1K8RyHsphivgyhVRB6/daN0QEUNJoh05gg
WTTDtDYy1Y5Xzh5/HDeVOPIv+/sVSjTc9JydWNt+3UtRaF8b+qHUGiwHPzAIc00E
KGTLygBYXE53G9sKxcEPaUCyyvdVONkISYfFLg/IgtNG6dAZWJgFRl7W6rjMbERL
JJVY+OTZ7yHLcIVyKxA+KkR+j5VD2s4Kzr+f+I618pdsQDFtmel3Lj1cUeSGT8G/
gjtwdO7/dxVcXB9+jta+pdHkGj8pIDOtIwVEJKH8HdC3KSl+UgadW9szFmxH6hwg
lp3kMaakOcDnd+6SEkLcDCK6CQbtl3ETRdK2/oI6wxL9NYHSVvZuh+5GKsseQ1el
fXd3HB7KH3/ukPJLG9zl5CDLDxB/ZdP9pEcvVzv8pB8j3EyQWwFNoKXNMwwniaoF
I8UmRzaaVkqpZYjpizKAMwY9t6ERweVvuVdfQ9a77HJNyYroQzesIi+oqZAGsFuU
da9Bz8mUmGatI8nv4dRctONbEnOBnf2abHzKkBpPLHhCnmO4IbVMmSv6ksGwcVxo
knndgfyATkeYgJWSVKJm/6Ic0VxHkgCYXSk42Ay/xvwBnkNcUcA2wTKlXfE4lEUX
oy/eKsr6kV929yDydgaQgpk6LeB7dIZxpEmqIzT7WXcpV4g94KHRajZzSeqZgsiU
jCeyyeoVw2kF5sURVtT98RnNXR1Ctk2KDA8WR67EEAGF/nRqfT6FQcRlTAAT3dot
ivgE/B+iYyHYnrFvIvspy2lxgqhhFhhRFH+3RI4B6TqyM4jlNKdKbOE/6qqUA35l
z8EELAoxzlXDCb68gCGPmga8MhpIGYXToLYHRqJopaxK5hXlz4kc2VxcYHYoGE14
dbmHZksmfYeF2fd1ve1k55y42X1IDYpBDTRtWoZkHCu6eL+i0fzLJdLG2EPBqnPT
quOUZ+VOR8iOh9eQrrkxtRCAjdksaiFDgl4gOmMa4wJsglasIMDUZrYOAhioGEDk
HRmelpPP2XEoOxI8yZ0DvEl94nBOk5NhAJCTU8TfIOk4rBVmuFVzidI7BzmnwTdU
gkBK/NI+WsKkvRy/Jv2MDau8YFLdLe+TUArZNOBiqi5q6SvSk8OOAqs38m81DM+M
3T0YHzIi66sPeHJmOeQGvMd6AgvbKOxG++7lYTI8HgVMDYJgOtxxL6IOfj0X+jHr
bGW6MoSEHZ07YkIK1MMbXPTxWl1FANzac8YRajUnzZzc9a2xSDU1toB+/32aLpBN
Rhp6PEMFJV2gr+vtrh/lprrsgde/E6GaDfNS+f/ytUBe7pYt16WQhtcUboZqRSRU
TCEMcip1KsDcDI7J/HJHJ/W1zW1LMOrCUyKLCKiyejEXzG6wUxVim4Sg2H1N5/B0
kCP+6wI0FH73zcXP4uLhp/l0DOe6bXCjXtajr/JUUsq3fFMCRsarLUkpOCKgfMTi
OMwaMjUIVC6ADxxhHRsCNkZHwR4mHoZe2kbgWpqEN8V8FytNfj2ywYA95V00tnE7
TlHRftKU6U8f3HEus88G69b+ZRNwg2CIlgBouM/I6Nei/2Q3GJc2XeDVqvXkFqbm
KL14EhwmjVRNZS6JVHKJwAa2WpgDJSDwwXTbCKc00b50vZ7o1ARqFuZ9UpsmHvZA
z9iCQVmzETZyiqxKrf8U0/uUujmWvM7pUgnMwgirbWJEFWNdDP5Gg1lXqhQbBA76
PzGVJEHF7E4JBAfqrGk9oiItw0U8E15VCvApSQeUUawmf86XraAbr8jCYOgDcsqE
9G7rhzGFOnlkYi//iZYWsztqjtoTHs2h9o57LzTI2ymU7vFyBZSWhzW/o4mq34d/
cFUyJ1rzGBTknzmGItl12wHr+0cTEt9IA8gtKAo0mnedoxCD3zgaabVMcEkdsnws
/5MI1ZaCD70vIqxVATeZjOkavZ7KJuZjQzT1XlKCei8MwgM85rbw7uHeFthcEYVd
UpXOfI0FqN9I4k7YFNoSgcQ+G9nHUDe51cwjSinM1kv6Ug/icbReJvQSBfeiaFnx
`protect END_PROTECTED
