`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SawgmAOwbeiNBlQn0qvFDngtZjg14b25FzT6hSwIHTe7
fMWvERNag84V+y025vmGAm1Rkwavk2PWgRpvJu6gQAX1wXmaNWJAtQ0rXwSTgXAr
ZZvlTIv4U+4OhR0GaZ869EDoo9/6Ys5u7tyEt9cnsVsqgCzBXD+QYikMHd8Fcn8t
C8elu10FD0YP12xBCnnG7R8nRaOnZGwx0+Btr3DvYKYNkbmiYRiJK8NN6QFqOkp5
biGo06FN+TDU05vN2zX1KXbBn0oawsgx/VzAQwLi94OD5Bx30Lrt1fQbqXrPDEml
zHuRsW418KZ/eN680VdE6a9gCpop0MzkJ4wgEAK9cqJ//+m7iGiSOa/AQ6CgJPVF
1tNapKgx/Aw8bBXmjpKIClaekoidNIjUnoKO7Depl4IdxCRB57L+OIdE/T6eD5/E
/j4FYK6JpPjTZwr5lF7CbmhCUSIIcr9k6GXcE+FYIwD3HMfOqKtm9GXHuEmmQu0a
0pqMOBrRmEhcKuRBASfG3VYiM7evxu/Ey1AgigAM5VZFum7+MM56rCZil181jUEX
EPmMDx+A1zOc5TobuCW90mNYQFXSWYsacHTZo2PHzKjaFaIkt+2QsNJKRrp8Fm6n
BJ6YEd1clJNq6PNGqX6Rg5RYTbMSHBu9hCgW10EUY84R7LbvK6tIVriA+KTu6IKt
oCwMXqZsnOmhA1s+UZpNlLYtyWGROxPQvqHpkJQEo9TAw9+pPsLPnapxT7HwE53Y
NyrkW7jm/G400YkNVOb+36bjshfA7ohMOHdg3x31BRG5d2oz49jXFgub0O24IaYj
RnfvXXg6PGmIhRoSfOLGMs74KeNflk3EXBOiNITnH7V7An11C0eUnB+iC33g1Bx7
ILuzyBtm3adlgGmdhfU4qNROT5ltfzTB3rcz+WUmkeaix3o0XzXFvVEWS5PbmsHF
YZiKoF6Aw0K21ZRyhLvCiR4gb96D+CYQLQFiOZWjZ6D2OLHdFEhXLaS5YdIUPJdU
MJAXwZrRCQpmUYJ7+if+Id9UzaWEg/Z7YFHTQ8GvOWkm/RFBQ6z8yTbUOLvr4lK9
mDJvaSRuofurBnOfrqbgqbUq8isfogfD4TzkZO/leD6/l51F+TCHBUKW+lj8Ci7c
CWDa8+1OHBSkzFfWMqAb5zBHt0NOeLuc4bnG74PqgQAwqszyW10OjwEYfyCO/lrz
u/kTs4REQnQbs7wwlLzHAZEw61C2t08W8OUqfbIIfs1XA3Vf1iU4rFXvV7AVLEdp
62UmLE64wwvWUdTMze4yhFMj6Nt+cMD8dkgDGOezu1bcK/sH2AooqojZt1d2Iuvt
W1uOEuRPszX3sKawkvbcunRcDx9I8fghWhfU99qvHiNwFjB/aLz5ad+hnNHnotxT
p4itG9qS5lZ8sj4FdJMQuEr59ZIz0+ifFQxi7EU8X3Y+onC8nJsRZfcpL4atD7nR
aE3kubgrYZPW97ITcRWSyPtXWbDfZxZHSBNIQDxkSn0ebvzAo2QIUeHgFf2vHBMo
nPm+UW8zu/vyFuBNPUl3wxqEaaK7C1hrivJBJndGX4Kq9sd3N/i8IpQ0iNeZ9BjE
diWdGBxO5rFgcnjTdpTqa7Wg121Lne2Os4ca2/08ICnyL9DOmVrpJY/iu2KYr79E
7ptxy1y0lNZpPisj68cucCW1ykrOSkS0V9LgKHt2FQCPb/YBDTH2tlDCOP6ZCepa
nR3uF0MhZXGr03Uk4X3mtHR1DZ2Y2u0D/nm2BYEEarMku0tZcgy3IxJgzzzW9yDb
S6sYeGX4RrL8/VSO4JureUFZ3RL5+E4ZQYK5WyohtcK4T6oeGl0oFDE3Ft2JJ/s1
8SeN7PYkz+j6S/G0mqXWB2pGwVhAzz3jAnydPn0u01txhp2wIs7bVgSRKFBhWQp/
VyYS8lnTBcJ341C+lU5B6gJKlez/hRMfoKuQ5pCDKNxAcfxACDIcjAeR7bcKkGtG
tZ20SJg+m9zg/YMN6+Uf0iCn1T1lH5WaHbem9Mr0JM5MM+rOwo+EPkPsGSpYKWpH
Cu/27Bsw/nAfMUs1MfYR17zO65f4B/z0qtXtOtVslGamsa0LqWVBB5YGBayUJ+nF
SDzM1gJTVPHcpUpDfuOCRpAzd97Uwt40LIR6h64ZJ6qpRS3KBAwm5cpyjmqAQx43
6UVCV/Q8jTr5CCab5BBBdkgrx9Jht/jSR1Eflb3V6oWzNFCBIM5JxBZ3fLiSl6Le
kzYWsFy5eVaz1ZOG/SZupVzV8dwAW6j8Xfn4WwPhHreGoLz2XUNIYYbiaEcwQa7L
GPARbkzkGCcaqkwwXEmnGoXuZCHDEOic4RqmZGt5fzu0RDW+uQYALMuxWqUhsMzH
YHhuTC7gxkal5dx61/3zpi52XFNZfqUXTB3RAkIMGbyJu3bqmsk6ChwrEbaxvP6B
easa+v5pAeVZ2Gahy5Dysdi8ifXYENabh3K8nDjPX0OR3opPKLq9QQqUV6QATyqs
aO3EWWekOVh5rxJYuYGBP+EuJOXWIE9Wttojuff7vsA6nriJkTkJg3Mk9R7DCiZ6
wCHHLpjHLr/5v2WTpSzaDh4XXHS3BtymbW6vUrbuMJEvgfwpn+Bjl44GTNZd7Rgh
KUM9pOE8vWQaehj5MfKzLa6f/O49dX4/lKtTXq3BHAFZFGkCkroab7fw02E02cK+
WDULlJOaNU82eA5k6u/Dn6XVA2sJO289FAFtGleYI8z8QAWXAXcwUnXffM7JVEyi
ddKQJbkWvLAagMqIoawxMqdf/d5jJ4nnFIMtnL1/2QuhdW8vPpNMQmfKFzomxBsV
/q42kzoEHaOYJonfCcmJwtWeejFpFtQ1tWEh7/6LN/4=
`protect END_PROTECTED
