`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C33AipHda4It1+TWZApoCZkXPrf9bydXt9GrgFLJP/b5
AKzzqRWx/BRs5UxPsS45nDHJSIQGpaqSwAy3G8W+VsKyCp6F1rQfHETqGfzRm1CH
wLKsA2Jcrgdzyppau9tDo5ppHSFyYLa+Re8jGlflNtC5xzRgvK5qXe39TD4RHCSR
r++dfNzCICup2zs6oTHesGK2ozkZL7K2orOG0OEOvgynE871EGD6RaE2zXNGXePc
D3o1r3gSgQuoO9YtvAIl+FoVKmprvwgovecUqwvVUeKxs6NDzQ0KCrTgh+qSRIA6
mMB1fV1Ee6CMou5RzDzO0yd4qRKT5knTh/Bc4soo5Oba8R6LDE79SyDfjEfHXYf1
CqGxrvUm6qwFnYXR0YhchYhx6nltl8U2UCYaufF6P76hUgQRVz22o7b3XL38QvfC
55PSFJShArH2NopL2l4wemaa8puKbu09/gp2PK+pDCWXxzQwGN4li1ZKEXeyVply
3uoZYjeU6zIbf89j33y8PNchglWO4jFYHiViWZkj5KNNe1aEXRwl/2ex4iEFOyE/
u7H7F/eS37zHNk8y7kIu//g9lQm0lGwS3/b5gtRGCCtyzBcx1AZzeoS3jEcG23FP
ZXT4zlZAtuCCMaY3cHq6k/oUmvHfmOOPKJMoZo/Bc9a7pBd4oI9cdA1pRx0lP5Af
IL8Rn9dQDEbYbOmbzIMqNns6Ug/mX6aJeOkihWQ9ZyX3KT5YCoznDGcFaDwtNUiz
WKHRHYCRSDHyRqNzkmuYUjHHizq5stZ2NnwODaw1OY1xSBvnEyZcfg80ZFApIanQ
4t9t75MOu81e088uPgDzihV5tWg5WLRuSAhMlGBpZR/tDMWosCWtBIubOfi3U7FV
QJTWJMSVrizucgJOaidIQc0NMnIR3abogG3VyCJP0zB6pzbH+2fNVwYYfrmmIlY+
kNv+CDThcJUcI92o/26uBjRF1A2NoiBSnesquPsvXlvTBHUjxJSjwy8BsjndlE2q
LTtX2PXOoLE7u7uz85gkHIuDk8wDTp3uqUseGBMyx7zZS/z6YSP0jeqJua+Fm2ce
nUiDQ+/CNLhJnHrKIeY4WRzEXKTeX8CC74gHLEPGcYho7iSIJ854An4pdxk6mfFL
FBx3v5DlG/SMXBYgc84pqFvNUNXFMBmcUhSTgrW7zANucBeGv+p6Rng3YlycEGX+
tYhKEZmu/Acb9PVHI3kUp+aW1jyzKBuDeV/r+3U8BjuMPqvR8mZ97BtBiT80ZDot
XZvFmiN/ydxYhOEwwm2FfE1uLyUQZhakuaBeoqYpDLtAXOGJlgOfdLI6uhoUR4t5
dHXgwgW/y4D7UevHrwSaJtfr9gZYt549h7x8dpKfhZPwQhiY5b4JZSbLkKyv0J8U
x7SeAKACk44v5yIo9QJBSmxOzyJOIGhH9lJH1jC0FEf3EObF0kA6ZrETSixsqbbU
bX9YfA4a0Y5SaZGvks1aiU61Iokhtg4rXYPnK8dB1dzS8RzCRUmvtqc9DX1D60Ua
ZPxHUqsKFWtLGPweXkgqTQMg8P/SXnSOq7LutcW0CEue3SLyrGP+2SFK8z16/uex
yuI0F8DGRpdX3u1rwenI/SvY6VR9NIgwJbh2MMmos0eAVYH8lInPdVGXY1VybLxP
2eFlRPAoFHRvErkCXGjoNFvUFTQc/PBhSffMJC7MGcNCxXhsfAhFQiZ/00sEUjJs
BvjtNuECGl1CW/MxLUGuPfrKwOTHn84kvFhZ78m/3NdFfXy6WWtWxyYmfixNzo0O
7i0+RCDzC8kHzMxYjek+E5tDI40yOg28rmp5U6ZNv9IvYXPAEIqQ3MuUFwnoAEqB
f1PV3OhE5XgZqzpoXc/hjRNt9V0RhemJ6sc32GFry+MkbHRP5dvuxXGWrXSI4VvO
ePAMneUYn467h4zv5AS55Gyyl2UdhGoUr4AiYcroykZov653MnVbSQKSf0MxW5qX
EPCWUpi4z9bLnMf11Dnj0cWdY5V/+zAYNviA2CLPtedYlZSmlIZ1k0MXROdoqejJ
`protect END_PROTECTED
