`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMO2lBbgXKqbtwJx1EvbhoDtpDM2n0KGxq/+JdbdfpPl
YVIKgdBq5iPPayr5uEffEkDqSDNsCcCZCgjQgjH1dmKt+QOqy+tKsRo+O50uEjKu
nrQ+KdQkcjhEKab2ANi8iPbfQEpu0WPJ9bKdQXGvgB/jD0h1mQFgFAlRlGBwOcnP
tG+TCYsCK7a/wFoAyad8536nXw2JsuvpiGG4TV0+7MU0vE4Eapenjj59zOMOJgie
kqsBE4gRCaHaeIbUGX8RhOzLlgZGnemrZF/AM7CBCNHHW0LPEjBpZ9qxjtcVghao
qR2xQbXnzxGPW8epFkR7dw==
`protect END_PROTECTED
