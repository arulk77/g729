`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGswdF6zg2m9UNR7NVarKlzKwconVFgwG5kYAyknKqPP
biB1vpq/atNVtIy0Scf9TBIjSi/LsDM3G4QkzrAz6E/vy22nJO0BG4AdzTOOgRi1
eNsb+XPZ4piea/uvPvftgXd7MSM0tR7PCBlToEDhnWN+3GaJB+nOm08aIEE+rvRz
Q/2wCkN/S9BJoOr8aNXEA/eamWITWIjvQ2yHTpYXTQg92+otFaPzFGAA8LkJ8i2+
`protect END_PROTECTED
