`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Xckf0xaaX3mV8wzRTcWX4HVorDkQ9TLecRTRh+E5VaiWXQMw0M0nXtkMVeMS4ffq
f4CtLg6eB3Of2JsY9uBCCrkazrwydxdfgRFNbpA6NU27efurenDy4f05zZLNLF0L
GntzSGN/9wIrtvBENVyZ0JhLrgopc+4Z5MXgk3NA0pwoB/mwWzKNdWK3N1/dzOVu
toHIRgvyxdGp0n/WfVJAVtgnzrd8gHRxW6uCpvE6k80UH5GG0MdfNaytKhs20n8L
067+WcIPCHiwi0gs8PTje8MHpvgZ6IxIRHwvTArjLiKmiVpD17G0hG/HfV7tS2PO
L8xdeVzx+Mf+2nPffQrgceoQU9dqYkaqplnbNr5beD4S/0b97nb2JugMIfdp/0/o
`protect END_PROTECTED
