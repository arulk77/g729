`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Qg1a/Vj5ld/i3S3U3woiPw7tRUvuKKKZ9TlAexr/eOqGy0e7Edpq4CULinTl7gxg
VvE/snYjnEAqF+tAamHp9RWTAq0OLbq4LnMU4XAXuf/U4JZuHFrClNAeW4422EPh
H5ha8PSH38dA2dRCdpvgnR9+gNLXDVZIGFktdMP2VcrnFcl1xEDgu2zZfRkBPHNS
x9I0OwPKVAvTlrlTW3HexgI7DiDWF0IoipTrUUxa9C/CZ0UIDbvAFqYiooPh3uB7
mxM4yDhKg62CTkq8gZd3zA+wQ3pClfIAYkbQZr6HsERTsS9OO3ge2h3pzjW9rgxp
mtvwGWuNMQqPlTEBVkw/Vp0zRPBK7FxzzlRnUUUd50GdUJzE4OLik4Jse0vO2OeC
9AkbxjOFNjKHgKZf04lSWdfU8gqk64Pi8p89uv1xlaE=
`protect END_PROTECTED
