`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAU1KhFHJ/qhFalnkaTGYCwE16SgptzcCyAfffW6T/6X6
Zapekp4UdgdDbxi8V1ex5uIHhxgTOkZ5D/NZ3N/RMQWsFVyZbGE8IrZaQ2Lb7kEf
pc5xLvFo/xurBJq3DTOkj8yxXY/4MvIBRyLz4uOZbjgRIt+z//wSMqfdetBMDwo7
YDwcCCG6ufcJ1pNRvY6fqmRRrNKkvOntfFI01GX31K0NGhLssrVDEeWzFdk+7/+S
3ZyGZlu3v+prqda3MyeLe4UGB+2wxu4KE0CcQyRh/VNBvYXxoUoOM8Z8JNdor53V
EoNgiQ+PeISYOriHiQu3Cjq0HpQPRy2HMtiYs7kRBTYSmyJwLmxXPxwCWA3ng1xZ
hU26EG+x6mPbkq93Gc9amfVgR04eKAcdey0Wvmqi0wadCW5A31HJwNooCvK5VpuY
S8nbpMbYRjIlyS3BK5n3p6hO+j3payNE5cf5F9ECjNv08rcoTmxg7fkAazE7le2M
X8Y4WdNuj+nfaj3kaLtok30z/s4K5om58pA0CO6a9Fm0l7g5jaFqmDwGaTpJW305
BfqBKqngOu051zerxpVXeZF1vKhiTkwo7b9Pp634W5eNyN2viBGmkZYeq3I8lIzN
K2UCJgBvEfX1/CaFM40/CzLbAN+TvPINtVgJkNxoXycASeduAeffNe6lMIeMlEzA
Y4KeUBBuLn7MjekNDEImaprymHaC30xCrJNC++0CE1TRe2qbu7QrqCptZ5EsyXzn
aDonjFu/XcQWPAAONTk/pbMQlVz/mVP7uF6NhKmcyd/bq2+ribrjtajOGOAdBT7l
Pchyh0w8DKLmCS2ood981ZYl9Ws1z/5CdymJF8WE9E2ROt/07W5fdC99Z69kttTG
L+n2N/TYUPVBbdIeexAfk7ScwVMcoOcYzDnoz/eNXKOaiNThP4VA9HjE69VuJYzX
vvuJSLh/TulI6oRkFEWpivnUUsEJLajiH9clvIRwURRv/wW80iyCVWaIUVpKjawU
KeCM+rLVR+J+9AbRs4qv6Z2rtpcrmywgYUCWEwGFTQ+8RozVvRG7ofUcxbYojPn6
GUW6dDn9HxCvrqvlsVD6ZgCVvaHreTM48UHth3XUzTJojw9x0cKZ81BLC3RkIqrc
SvmZoH5NeWf9zYF24BwqqbYJDjej3s1ImY3PUL4Y1ViDHxijfCfsmyysiMgln1NU
cMGnle/DZZMb6oTMBC5dwP1p4t/0C6RdlmCBOKTTZLC6hFtSGdn1gxu7BZBNh8GK
P+fvjxrbbenHar8PyUARnp7GAEeSkh1b9CMbYZEEMnIwT8FrWs7yzCYjsEgJ0xgs
Nj7ZMbrmICh7Auyq8dkHqvl3BGEUKfioji+CkudUIIuH6znQ1ZOboZh0+cZOrbWy
NrY5tzTYDqDz3lFXUExzQjZEgdG4LZ/n6mq9hHulXjoE7Zd6+bLkswQ96eDHb6TL
xkIL4Fd/Er3uCBrjc5TpVc38AjjkH5aKbGaZehcHJIdNpUzfSPJzh+6OdnD81dtw
IWoXtuUPOlJeKU3LlvhO7W27DHcszQv47263OIik/4z6YF8ZaT+uPrK2JfLRDbnI
ZdWpA5dGUc9NXxfqbeBmC7fdXMIyHJsDD8cY5ZusIQt6PgzYDKQ2enBOfqqQAHuU
ECq1pQ1mEgIxQuEKp7Gz2K08DV0ADRtJRBnImGW7fks3RlyDcQ2I//Luzx2krrdt
78+ugq4bmVWq02pilDBOQkQ7xyk1dzvvKM9CQR7sPMhBXcyp/4NTvBhiGFtFGtO1
6gZqQX0C/oZpzsizcUKH+D/9aMyhwvn9gStgHQLGfPSDmxIhJSxeU89KS/Zsl/MN
WFV+IQAtxvZ6lCBc7ORoHNo1wYaQTvDa1iCAyYVIQVuLoPxCG8HsloPOJb9QlL3i
smkogcjJjzljWfmAIQ2mnOCl0Lqj2HrgwMQYgvwe6MxTekduS8wqDIuYDdSziJmx
wU5Qab6VpSIrul4XnsnB/4wxak3Tfq3SkQvI19bUY6GjsFN9CPZ6CAFlTPeE4WO4
6AfU4LP8L5tOZOQ40x+zvSEyyFhQKRXGCWtTQL/IXlt0Ine8ubEa7w6hhl1dwkRg
SFy9QJjwB4eCSKW8p9r1OrzydRAndNPg92h/dSMAKSS5eO8hZYz0UVLjK6rl6saO
eOxJ3yPnRjhf8ucXOePs2khfXnYyMVINbAY/NHlHNPLPbE1gb18e4nhGxd4JqXQx
3GcyRJs+pGWcdmcQA9A8XQ==
`protect END_PROTECTED
