`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4WOzg57Aeu6zgB2ifW+nYnMAdlBc870wGoMLYTX346exw8sZ+MjxgYjQjpdQbCz/
AuxTYbPhlBs/2JA2+ebe25iOqXFi/psL6MCLxYXH5UGsN/10ixNFOuCcmC62Qmpb
xADmQuaAPlhqdcZUtt/d/YGQN0q3IEfJviIDkIxJ6qpgI2ja7K77zcEr4XxIa02b
x7eXTGriVJGMRM14YLcgS4U8/ujzDflgGmlg3RhA8BL/D8upXPOWxbR2FBX67DBL
7a+JnUTTJHGo/jaNCtx7xH2YfRhJtEyKQ2Z/cw4eWWgOyzKKSmbvvQqcYndagYEZ
c4wjjs/+hnd/iILAm12vaw9kXFhnW2LUi8FtsCvV2Gy/FCvNHQ/1FIpIyQpDFBV+
oKzXt/qz3GRwvaTtZFH9jQ==
`protect END_PROTECTED
