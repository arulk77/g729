`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4ztosfAsulrAay1BASmENzNHC7e+1+ATEMa4Y9wX5Pi3
Gew1BbgZnY1x1S4IjGasfLhbv1zLcSl3uQQVVDSOJCnfWpvQ5sKhZ94OW1s+C5Db
jsMyBVkY6eP427LZLO1xmkSdtqbR1xySZVqOwSvmtZgsuCVtaxnRjdLNOv6u+NZq
6jmRQ9N/4KExK4YchB91A+UEVNgp0Mm36sftYLyvaBgnLEqSWiol4yUA08NF35MU
B965TEMbVjw4qT3U5nvOpctgVU02eD7BHjQJEQyslWlB39ySqPn1QcnHewlTuvTA
bJ+tOzwZxc92ja2Uz9EQK7o3NGCekiFcGO4m/wUGu73s9mrARG6i1dJaGY2vPt1t
v+cQRlhWuoDpgO4d221eVA==
`protect END_PROTECTED
