`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ3fcglJLIp2NV/sROyQBR5VngigeE1t90V79+VMpfB1
vfYaPQBYa8UyOpKsJwldtGDzhM+8loS9VUXnmdNKoviI0DBBoXcm6M5Ofo0k81JR
rWDzgZyCaN32we+R3Vk3vjGACv/Qgf04zrG1h9QW14iYEJEFTMOOb9UzGKEAF6dw
6q6euTjGIFZa747s6G5QAjf0aaUGWrlHck2dGe+TUUj2Xil9UgpiC1lSj2VWJJ+I
LN2hFb4sHw2oyhLf28gC+XtvDypUegO/txSyRJxr3XN8cUCuW2n4nfe8np14Z3X7
FptQ+YHhO3pEYGMkjOWDuKwUdyZbk+wlisX47hHN/d5u2zuLkxXf1cZYl2zyjAN2
zFbzWDaio3wDWRCVitLmugfzQov1WJoqVUm5m7iimVB9ConlxO8ruQ26vb1sxiv1
/Abm1gveE57wBuFMjLn2kcJRzM0TEV5VQcAle5dulSs0rcQFMmECqwo5vNbAe7BE
meiMh+XYABc9fRFc0wuvQ6DZHqdqZN2TX+HcJrfZs5N5AIsXhR3BZiYF3jBA4zYq
3QqY0vVyVJ4x3/bKF7vGRkzIapXJZZHbf8Vav0HMSlqraPKqxtct6if66oh3JWad
w03y9UieqKpVFc+PPjWjGzG3n0u70i7bSPJt9AoDeAA+sO1+WLvf8O1benjLXpj+
dFUDQfC/lCgh5sKA8EoKmz38ZF+NN7NVydlmI4d87kdN2ZfSrv/CD2UROuO6fFbE
D5ayfzx+VdZ1hIYKsms4REQ5cryseQIsb7bSPb50BxEgc9xC82zOpQDWDlSztW62
qn86OJODdTwII4PTvvWxEVgCI/JEm+NSc2J6pUYwJ+U=
`protect END_PROTECTED
