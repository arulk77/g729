`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wmTAMJ28HJsHuT3Ca8eXzVNuCXOPiBS+f36a5v8swM4
bXbhu8tP4QjexuvVu33hBuw6AakEqTG8YwvDrLj6VICxdW/Snm5n+ND/hPrL0rfI
v/JXYhHIN2WK+rIsoeFYK0CzGDOKOaHULgnp5p45Qxm/zoAph1G/i5ucNchPffer
XoiTTBMSyomlHCHXmaTWGfuUplZXiXmAJYh2FyeTjZ4=
`protect END_PROTECTED
