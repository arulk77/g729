`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+wiU/N98DAGUUG9cwyAzeK1KhA2PARtlXyPdDDbzZhO
D6EQtLLUsG0r4dB2u8PHDhAcWd/eg2wv8mJHoNVqcjatbJyVcftmF/U+1WPnI+V0
+ni6feD9JmIwvu1sy+7S49QddyWsDcXOtUuX+5KyGH4dkaOEP4yuPj0xL0jfPM8U
1ag8sVj7M7sGLT2fpva0yqqVZRyzFq+IxryIXvM/rzgVk5Yx0J9nvZIKnEs1gzfm
yoHMET7TAcxBqeFdPBfppsk+4um0ZD5ujRIgNWR8hy0=
`protect END_PROTECTED
