`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bLBVtWGV22YgkAFiPhkCL9/gI9xJoDOXqFMEctXMDievSN87Hn+22SdrAB+RolBK
LDtwru7hEpoSwHKDNiGlZ42kR3afbckrEDiJdt7U6fSTo7ZGIxlaA2CpOEvBFemH
n5+fSwnZ0LABAupACtHjXCXmpavPdhjy/ESUjXjfM9vKVisrfx85rxnr28HgvpA1
MIyfscD4T75EbwwFGsU93GI3lwKF0IzbbQRPYXSuJh3o3L9udVl/3TB2qPTGkjMD
GDghSIwpDNie/v63fadkbkJV9FZi2/UAAbp55i5uugSuMD90nHgrc1df/uugv6xE
TTYrvjS9I4Y0EcV7coCbt78T1Xy5yLb4Nf1E2kw5S+BD2pShIh3/sCzVNbP6WuUJ
hFWp7d/a1gLmD34W/YHmNamJHCiFsDj7RiTIYIyRsBe/K01khi7PFlQfm/E3Q0Pm
RjYxqGjPoplGEg5GPIXvSg==
`protect END_PROTECTED
