`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41DSJzwBUQjA/ZmQ0xOjrvvLvqA2ExHQmNlr47zRKLCl
t2RoMMWa/AjJIYx8lLvyXL1/UD9DRK5Aof0pkLUs4Puek6j+r5maPCPppIM7TYRu
r1uHGCVuwp/+GudKYv7v4o7okixd4ClL/2KmcWXjMejg95n9Mr9dvPzRMUQOJhP3
FV/cKYwxEGU9l1GAYQo9wLoPf1CvQ2qeMUkhB69mCtg=
`protect END_PROTECTED
