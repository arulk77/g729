`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3ON6twM0bRyFDJLDX3TyevQhWWyPTk5ko+CfVDcGFDkYIZv0jwKGhXD4uGh1bjEJ
hDpsdMaZ82mC8I381wba4OX08whr+i+5yFMbfuZZ7VujbCtne8KtS3w/U5dHNxo0
aqZ4thGhhP60uKm0X8G5j6u5ii58LyvSQtIIFRLuGwt52G6VTD1WDuBN/eCVbPnS
oRkiF+qoBkIQjplGJzpVkg==
`protect END_PROTECTED
