`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM7JmmmKKxdGKuGx2yIJ6yX15DaKbNcjcEVr4NoAKwZ2
Hg8jXQX77Kyvz8cjsEEqWrUDf8JGrwejLlvWM37akHgfru7y+rKid91GBomZOQkP
fb41xavSuikGIi9BfkAEY6HLqO2NitkAor6cVyj4IxZK6ZWid//CeNazi8iQYTjB
8epTIwSTbSqJNBv5gKTUh50kXJpqe6j54NC4CEekty4c76Ioghk53tlGph6bZE8y
`protect END_PROTECTED
