`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDo2lXpdNyQay0+qgmPV76NU5Z7IdI7P6OmS+Jx+9uZq
FhhvzY2ljT9sfm3Af0MMCzFpZAKyCGUI2Igf6oOPxAIb/w63rYtMrt/WMJDCKjcm
v3qAiThppJ5MsnDTt8WgKjPGbBn2iShu8/LEmu9OiuTpilEqu5sgH2LeOtaWbT17
+Mosvb9Nq2lCWFTZ2awvudVhJ7lrmIbBpZ0rLjW4jBoNrDPUq0CpYaU7oPtu616u
sTUPJlBHrvwk2I+MH33WokMdFy9tUbtsaLOs/6JHNZNgEEuDZMuqLsDMEd6yrnZa
CiwlzsJKuPE8DDVMJ+UxpcK8BE6uiWDe7DLo7H/k6P7+8ANpS+ZTjooh0arJmaOX
l3Pgih6F9N/f4Y4s7BKigVcUGAvgOdpvyxcVTjHzrV6M28lnpv+RJIQHuwUY2QPL
skKpDa0LIoZPr+HJ17qBsZzeMoRK0PyUzwUzDFrB0DXgkCIYeYEWoWzvT3qRGCcB
/PQ7Sa2nxoLeMme8dHYgFeGHLdK/72RJ/08S8MpNwu1P15HzEk4ZIaglQ2PZ+1tW
S1m3aQImexLyZBHBLemOXwbOsLzk7vEk5Dn5ZmSy1G0RKUos41TvO10iKP/sb1lm
UpYpMWoywjV0arHh43PjE7Ooep4XynqYmtdoRESzXKBn42YUqGoJ56S8pr/dn7xV
+0VPsKcc790sIaguOt8Y5lAENl/fbcB9s1OvwXjf+Y4Gm+mu3QSpFnoUROh5mdc2
hZrH7Sgcw35vr8IECLkqlQ==
`protect END_PROTECTED
