`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C+TXfxSDkG5m0zjFL3ku+ufaetfvdw+Vj3PLYtlEsvsC
4xHvEzD9uKnOsnK14APX6L+XEk5bBwas6vxSU5bin7p+4daFwCM62rWDXela+DFF
xMsE9MFifaj7kJ2jq4krapZl+BOKQKl+dOZEpmkBF4rhDG5jVedKa+VPmhFgyzzv
KhPtQDgMCojO1tYZEto42bqXDhnrOkMK0CLHuxDyK9xY5AqUaS0IbUeCPIvXzSjV
4I1lgjHH9nVqM3CkZA7wr9VgHvpzF5e4Y+pF6PG7KqjnOArOysYs68VBys3mhfgZ
O1HmIkRiQ7mIiX8nZBdwxirR4JfE/7byAB67eL9zqod6s4xWMztztInfqgWssvM8
MQAewukFrEhlXeT0TSi93+9qHTVjw2pjvEixaJytv370TqdadyRD6wAzi581Cvbm
3ES4/4bkXZJgKbQBt1f1Li5GFt3pjtQL3j8PNWAD/SO/Jwo1GqYhD4YSdWgG/B3s
vxmJVCQc8kdbXOtanbGyW48bUa3DRJlfIJFExcxdhn863hIlpZfCHQXGEuNlSYkT
0FaoCEbjuWPtptt9Lc0QHh+wV6PommpyODpOp4vNIJYS/FBNC8WL5cty7ucRBdwH
CPvI+geWfOjd0kjwH+K9b6c6KWsirZ9m/B7XK32UDpNrVSRmsrs/eW6/LIUtztjJ
F68XVg+BbYQYt73RHZMPNErqR54U15Qv3gMk/rvkgnUbGeJhWhHqe1BYE++Rfc/x
tP+LicLn5F7+oeVFJP60lq8Xsb00FNEqKCfYCDZvf5c7u8D3q/v0ej484h2mTrTv
pj/FEcWnB/A7uXomn16jAwrmY0ktPJlnVTsKmgC2jpSBC7UhNUl4VzOuVNDgG5QS
6d/Uvc15s8cmgd3o9eXjTkmQLtR/Y69TlkMRnZVLXlyXatU3HyAQaCTY/G1KVfif
a8VNbQQD5GNbTVeEIsu3fD5BvMGlz0Aht7yWgXQ6B8WK41ASLyQ02wuhz/rFhOtK
y4bwyxI0WF57KvXNDb7csAmde757Xxrkrm1ER+OovYfTIgamDn0hEn1uYFXwU+vN
iQM2K+PTkGYj/JWJJfnIhftBdle8faCJwkebMwvu21YVGHWzaKrYwrbygD/TsiyH
VYhIW76FDXtc8R3ngOkQdXpS7F/ftu3ppNKY+MXAHyowoWeQu9JOEfChcxV5AiXQ
5R+k0vZ8UDKpRf4jEVXfzw7ICGqjBsPt4YXujmxaxttn7czeFzKSb3JUHv57twCq
+uUs8Wgd8lKzfGJSA7ltjqpVI+PWDGWs9jGfm0C+vTxI/PiOVLK9c+6aEhWgMD6G
STgsI0szC48Z3gjqnmw8KS/lpQXpRv9ZHqi4sOE305mFlGShX87r/uKyTTb+v5Yj
2mxYy84pURNJRKbKm7KSjAS46XiO9rRFQCGLmvomZqpWfOnxdygHic/5t7JMWU7t
jo8NlR7gj+25wc1uY304AQ==
`protect END_PROTECTED
