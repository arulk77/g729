`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3I+ZE63G0VvxgXdg5dn42fZ0UxDJQeWPGlB9aKAu1KoznNSczUCcLkrDpN/Cooyx
yS9xa/xAVBSBRCZ2EfNrOzjY7zpIfNOlZZ0pvO7o8+9Q6Swjd5M6z0AIAw3RwMt0
9jgQAr8/JMmEVG8IwtElBuK/3+8QMA8q/yll9pyJCy34p4vBaf/9/bdtMOgbsAvY
nyUY0lvgxqYKlDV21mbnwgQWuTz1JtVj3rqQ2wj1RhzKtK2H+b/hlDlM/e+z+TAA
ttqIeVJrwwfTViM4nInT1a+woVw8julUgVYdoEYv673OGkPJzUe2tkgM1D/Shjvi
4CYetc7VOboKfyO2EQpklHUE1iWi0Figlu2y4vnFvd5R+wdDwEln7wIMD6Nuzwv7
oSQ9sW12NwuFrmkMXe0eK+fIi2wPqaaFFEyq9nwCHPI=
`protect END_PROTECTED
