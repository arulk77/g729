`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
rDpeiCkLYPNRZHyXSXzLfrSXp3mibTedZLOrFhkLKA4vvqbPmJGAChvY/I0ORJJs
XT8cve5SxEbnGdixVdcFB9bwlkZQXEM6/lK55YMURbsD7rL/gAyFJlTdbqhnJBat
o0Aq/l87KCom1C5XIv9YfNF3tc/A8tPqhp+iE9CIWA2a3GJ7JJj5EuyL3q2UrRDF
6cF/QUY+5+4obgR5UmiW3ax6dX3Mtc12tkwzZmsp6mDO5MTGiK0xAiHUkLz/m/kK
43DV0TSae/ft7/6pEwxBG7CAtSZSekzEz//2+2kf7+takq1zpZv5ZFgxnB62z8zj
2eriaYqgCVxuHdx4q4g6vLigztX2uuDU1rIbrPElowc=
`protect END_PROTECTED
