`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKb1QiuQTBUrzNXy2GSqMM4OuLZj9anx3B+2iZnvbsvh
6zpMkiEqZqpSKmqcU/YlA2Q+HIV2fjbJASBbCxtFS4NMJ6ZRrxmdhzs01mRB9C43
uG1aS24z2vL7tcnSrLZH+lZ6E5vmA5XFncfA0im8RX+m1XVHcakEkSvS7RCx/pTK
Kafxbs/sY5Z0/6KYl+Un8Q==
`protect END_PROTECTED
