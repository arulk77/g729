`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveELEjhqcxUe+u2KACon8IYMeZBztx1m9GgjykoBJy9tI
Wigd7aDfAmurWpssuMF6vm5okp4t75gVuFkBOiGBO2ViFAQEA1M86rQ1orAb963b
LleuRiNCmLhd3GiHEZKnhT18sjTVTdLAGPM/6+puy/dkdAc62wHeaQmEp2I4VXqy
1LDIgZSG720OpS9F40/UwCTtb7zV2GCLol26MbXkjZwFlF6g9SmoAL2pk23j1m9k
LABHhSzOIiv46vciOsyHwikKBPOBEv3XSjYGIbnvefBaWBXMvT0bkyhSqm+7vY+2
n9j8LVjxVGJfmToEwgnPoJTyWyn/w0BLr8xUivBUaSbKe08veKnX52iP9KJJFVsz
d15KIXr8xQ1/GZD+e1Lzb3lyy59TEe3ehcwERXsRk1cXwUxWHLrK7s2f8MftzCrk
5qMQO5407A+6RH6WfGewN3jXlYsnlVoNFgDWbVUjzJx7MD1xZE4Cta8pKatLsxWK
UeRkdpjYBOec+9iFSXpG3c/wZCLLXpByLt7k6d0eUB3m80WGyRuSaXUaeOji8UYa
C2S2dwEcac867G9bAwFf0Q==
`protect END_PROTECTED
