`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
c70/bWEDmd2eu11w/UzPUyPQELvl3y0QBDIonhaVy8CDqB3n76rqBEst2urtJId5
9r+jNzKes8+QV3FL2DbGmJqDG9Q/yGjnP9ytBpdxAWscROZrmcdWLRsJefvpUVPE
F1q+OvP6Vn3ia8G9rKdTj6pdVTRwS7zaQ+H5r9Pmi4qI+EPaQqzckfM8ufu/YHFQ
vOGXukEuDyIIZ6Kgw5c+uf9V3rmfE3lu6vSkeEGiS6G5sgHOwyu6g3jiT4gbxWbN
RUkykuWvQd6db5wTeJ6p0Q92Xn75zh6QZO7QK1dRESJI9o8uhlypNJgoX8jd0ndY
pB2yhB16sngS1BNhe5z3PW97q2tSEPeS+Mv9QzReJqc=
`protect END_PROTECTED
