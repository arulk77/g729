`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN+gpfKFlBElZMwvoOZmalg+rpfS77lpmY2426rULmMEz
FfndCHT5QA5SJkwwgi69uKMC8h3zEBmJfW9/s+7GXJgvX7k5oTKsh0oX2folwnV4
/N1jFSlSuygsxzYfmbqhqj/Nii/5qbNLT1PTSOIqi9s4/GS2zwDR1K94LUhnRWBv
RMJ0BP3Z2CewSGU1SREfIk+Cr7XZO1bUt0L+vBMlu1aAWadtsc0p0al1fzRloDnH
MCp3BY5nnyP/k5zyOtvOTZdhqrrhcGeDZ1Dq/cSMHcOBRpmWtojchJs2C+aduMLO
fjD7B807BrP5zCrqCN2A/rhpcK9AqBpq+ZSQbjRxkz2rm2AHMgnq+EEApC+ARMMQ
uReCoLFAp+rmq8ZGDqfP3Qg6k/lzFpP4QhzrmZxMyb5cgU8lRzqxvH5H48ukIPZj
G+ba2BPeXE8mrvNsKQAIvFOgpg06CMXl7LgoqwUuJgB1VMrx4Ro6OvuCn8Dk12DX
azZPyAAqu9Aa0d2n+qJVzbamXaERQicZqJK6nYW0/e0f+Off0SCRVXo9kNojJmuL
Roxe+5plULG+gCquz4R3PKWBv5Ccszwfw+Ze32ZDPVIeuxRNJRV/n6GmDY6sD1W3
6qdFLjsJvFOWVEzrSPYA3B45lB11xsRxZJs19tdOf+Tcvnxin2IHQGkzAgxfJqwb
8zPB1mzwsK9WwKeeXZI3os+I+sWqeyaTx4+9DAMut4hMk9fFnEoB1QsuYnXv2MiH
wYsC68a+7ln5sgiyg2Aa35BToBj8Bci04of0cET9Y6+BrM/LeWeX+WTAkUOefugN
KGTTiWV/lPBJoGJ+acryYhpZc4X+DD3gwhOuxZ37evuUvEXOiSHckQwaFy4vM/Rw
I3kGaRUqPjmccsdZj0OhcWNc5AnWofdY6gu26STIM5swwvv/2c/YiR+fPtUFX/xT
th5g35dY5gU/dKsuYf6KZnvCY24ABu93iLOgB07HzkrkcL7tR2uwLlNy6GFg4/Iz
XcPYiyxI/2VNKSRG4w0E6baT0NY52OBbVFFPT/tDANcMF9SPxypypYm/bVVQJ/ra
LzaEg/MJG9aqBRKEyspsT0C9zv62yUROnBxziqUphoYB3qThpkUGJo1VYjFrt3rL
MSmeuMp2HW9JIdWgxcdQeXR4g0J4XYC5mYaZ5FcXTPNg+g3Y0PXmzR5hDxttCvM6
s1v6M589JFDvzaN1UaGvNlqS1ZhJgfZfOAY1zREUrms7Vtw4QSrAsQlQ2BUEftqg
/oNgULFeVb2iW2Elv1d5N6GPR7iIiw1vIlfmjTkU76dpMqK1MYmLBOrdXZZYxzO5
syD2vMymYH8CUk4Pw6johEbNJ50xjZVdfIo95ITVkJrs8j5fZAELl7BcufIIDdtb
b7ijrWu6p5XCBzt9RH6jqRYPZkBWm5cdnyNv/y3Yk/fP66UJDAkUSxpUv16eMbxr
JzJ1dE7kvXSrc2xrJs3lShsJ5WfHCjT3xjj5t8gaPQwDTQ/I+f2HxZAkkNILVC+y
hDVs6bFGJZ3M8xXKaB4F9g6ahBNk5a71zV+BiJ6dmx4a/vlXpjgRk2Dbz2PuBbHZ
2a3b99BmLbuJzeKJcY5Wuw5bSIfFVcOefm8eTf3GMLkvSYkEu7/Sr9E2b7GK36SA
esImp/nhy8pD3TmDJmm0FN0HK23SCV4SfbtnBhPwjHIqmxU9+EQuQuqw/xHqB9Gq
xtrUrFUuj7/ppcEMNluQqyN4Ynya8w3jEF/nqfWSc2Mqm5n/JbZde/TNIDNCh2x7
rhjov8xxo+Wqe8yFz4F2gcRzjNUoFoE1i1j+6EtxwzMBlLcruEJd4QmmzGDi1LX0
G5s7aHYLFDidI6SnPeHsQ6bTpjKXEztGZm+Z48YeJznvJQlQo79P3Ag8fpw19CUN
rXc4Dm6KzvSuFyAYZOYNnVJW33xQEAFLhLl+qVS1UWn4DMLwzHF5bw+pzEa+5U1P
GI1o13Jqk/raP7ADVR2jPkWNMdnGgath6CAAKGiCwdKa9RvqNa6jjV9JXEBZD7b7
QkZ/EL4KKNla3O3hlo2FEYpQ0UlY/W0Z8xmYFZM3nlGhQNeYuC0dDFbYwtMrT0+C
zv/q1yb89np0YDjKaHpDZGP14s9PHADzR6p2LBlODrHhqI5CHDa/SCwre2EYESVv
6LUi34yIhpNBalsvUMAIvTBGzZI9Eh52sF1cAKAuarR5HNNmwQqgnxEaW1LwU1YL
doxvy9+F0K6IwyHTLl2c1wZz3x3W77Ut+P5LQHUZM9wMOsd6QlbaoMHuqPSDCLPr
2kmJT7N+zc2k/a28OkqQxqgdDxkZ3Gv5j6hpJk99qo56qjOMzZOPBX3/KZPJkEGa
8Wy0hvs28T/o2AIXYpw862u4uNLY8pEHdEHbA5MFk0oOKPVnTEfr/GVdtjh6elCa
PhnIne3MgGA02WmOasArZF30yxfgIHxB/4xmj44zYrxwBuaqwbJ6qF/ypFRQcaDx
HqOM30FSZzs30ee57ARe2a8Sz5Vxux5eIQ/J2r1PKd0GuAsEjst4Nb299CLmJ6c2
9AxTf3/JqJqVgHzM/zd9JGDzP4dd8wOKlTqTh2ZQfSBMkDh4j6Qi7+ci8w+HgBEy
bTK7gDBXxgcLLuZtRWbbuQB4tKkivcUh75IU4c064GhXIy2UV/XQwDA5ZX4NP8pq
vAk5DTzV4RdtKQ4++W0FGfmjKR1BtNmy866d66QC/cAjMXzZRCvNRfPdiib+5xIF
2OSVsBv28+PX6XnxJ4xz+HcB4moQPwigmYASYhDwnb+QKFDUbcMmZ9lMf95Rvg7X
jVih6T4i7YFIGuGaSmaLLj9Zf180EoBq1h9WOuBu7UUL5J/Vy2WOpwfQoWn/9f2B
RQXgDu2Q5NaWTI/ww/QvtHczW4O/QxACIIw3T24TSc1FA8LFRcV8+iMHZLjCMveI
TAJHKuXsofOnrW+mnOyh2kPKns0F1YTuW1L7OpgeHmy57pATaFnDdTPynbKA5GTQ
biksKD7aNMQ6CDHOBFphVXFqrVjn+miSJJUrHkUghdMYdrTZd4lcdzQpbVob0Ea1
GEonVMwdUxPwIUC1RhVoSzDDfNDt/acfILtZJqU2OOAZfF+FMkEzL/4aysaMhfUG
bdMHwidb8qS1dYe0HYl1omn1FIyPAF+A+UhI7fHC/ApxeEzKbGVEyupEaRSdQ8Cc
0ddM/dB74ZE/BVV0rYQn2IgrqcWwtEVnEbK3r3KfEcSxbrOvrDuudZzJRsPxXOan
VD5hxYhb0pc7mDAxjZ5T9CceclsX4DH67110+HS+roTQyLXj/Wz4XUVQPmM4iYPF
4retgpqkBa1LxXCY58OzjL3I7lFfwqOig/4qAvlkyFu95yeEsZ2srjHhSrI4CA/y
q5R9P44veREa4cXOoAsuUfrOpBz2KVolNLDWPBgYxOhvR/skmuvUlRveiL2nCBqo
qzT/89irKw8F1PqsExXywavJ1Q7SVjU27wSW0A2YKDNKqCDgutyjY18Ttu2wkCDd
TB9yqSx2RyaJVjFsORahTK8pw98XzyHdWohMrePi0mOyFG+FqljyL4z9tUeWWtf3
6eHsSmIbpshd1S4wjXcacWZwxl/z7Kvny1lS7CtsObFK1+OPSKCDMUjTAEAJYe28
d7REq7C2bZbQ5hsAonpOyg==
`protect END_PROTECTED
