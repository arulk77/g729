`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAaH0o+NEO+FAAxAmMNmiQSEdx/OWuZkzGrT84+I/+7HT
LzHkLW0WAkpKpLe4LZ1JrjZKk2gjZpHX4PdmUVVISZTrBVOa1vfxnfXBwpuZlv7C
zfp62Q3gloahUnjFXWEXifj/Y6+v1bHUfBOySpBmNHbMX0h796EoAzJgEKNl4q9J
Hqba+z7zuwY4e73//irSvkbO26Whp8dCBjlcXtHS33NTf9rK/Pd62Zlyh/zcyCiV
xSK8GZi4F05LU+16DpJytpHdt7E7dv6NpwH6cjftlRGGsiakTpYbsYRx1WVu4ld2
CdwYQlZMW9qKVO7wzko1s1NxNaUY0fMg4NFIt0qVsUKGPXv6KCbrwTEPBx+kuTbz
pjtId1yryFlTP/EqyFuKV43AucEtfTIeod2p7H3/6b3KNbROIu1SsiT8VS13/nTR
ldl5SKQESgMTyKv/QzRuc44Jfu65W7tUYXVmh4LcHxcp9UZUhqltcGUvJGASOBGr
qIpvwvJH69QvmUR0VxD1Mxj3Ff/UpP433sY2Ci8NZC89mWli+8n/HEJvvFzeMQ6F
Guucafccxf0+JfYoQXpUvgYOOSliB7y+VmFs/vfhRFsYaZVdW38DEzvcmtvuN8WC
mZIVUwGQ4bbwXLdQuOjihFEyB62fU91+ZapbevlDRixDQOROSqda7RKkZFwde+Ae
zg8WBofhBUCZTK1r1qdgyiuHiXlAvvBUT8LNgA7vr74Xa+CuGXcshYz47cfiuo0X
khipqw+7FO86FbYwRMdpdg7xntyBpgOTqXJqOLg8mhL6A7VIFHLYdtUw5TAL3z7U
lSdpnXmYrzn3VYJlydyxovSfnAE79Bq8NlnEgOesN45xiANpvYurnJuXJDAhuakG
02wlusPjQokYlcnsFueW0to9f7DPGP1vLid/yJUj8Fle/oTd7NWPTOsg78/zyDGl
M7wEQhoXmdWFTRgCw4L9oM2HzoKQMM64oBG+xXUB5rhQnScUosWj+UhnTqq/6u5H
YJ/Nvn8+ZWf/BEyly2GFuh+EIE9W+l9s8ysJ7bnogxAO2hcRxmrdjHg09p/rusR4
DGmCm8bBn/KNyv178zsI8HsLZFwudNI2TPWVcJRQFTwA6vCLwauA6NseXtNiDhDq
04Aemxpj0iMHM6GiikSbS9mjmKItwiGbldYXAKxDtWB78y0eGiD+xx6kaZhmcDvx
S5vpfWE3AxCH/+0Jp1T+PZ/xR+0Ii+BwXMxnOkOLfg1zchxSkWFwPN5MnQCAYTP2
IZrZ7kZIZ6qhrJPmIunvV3Nqpv+rqtDVnxdB5kzuK4UdiRAqD7YdJ9H4TfHzGYzb
qNMqlMg+qXcLHXsTpsotDmc9aSZg3kzXkrvMWFersE2x8WVw4ZRp+XwlWUxyztEC
JTTZEuHT807uv3c7VK0PktrmJ5FGbxCBmWroFNjuadHWkfbQc2b8IGJh9cB9bPSs
9M8FJ4uytpKREaMGeh58VPH4X50sjXUQue764dTH2Mh7zTsxoMaER/gfJQvXC7S+
iFvllN9uAHebCIKaWEqwvQ==
`protect END_PROTECTED
