`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
lQfo6O4+OJfXZmeb5lsHiudXL0mNBP+fE0Cv7mNcZlFZmCD4qf3IBeO5OJTfKhin
tKxV4Z9BQ9bWbORNOYWUpNceq3rqkfUv/mZ705oO9XWJE+u53Vdve1/P6N24POWP
WNvFqttqFKGNW/hfa9p97b506GTYCaeUEUawEpkUXm4Yizs/Peqmq7BIcl16pCQJ
E21ka42By70Q7k1TzQwhgX8R2Y6lf7o3SK/nrJPuHQi0L+3DF+NgalkuvEX/pn1+
gsdHVqmujBB9dpNhAyj85Ur25UDmY7plvlRsgiIiQ5Thub6FsBdAhQBs/hfR6qJl
iiz0zXdrkIe7nWsT4bd3oPr+ALbVTpuF7gYaU6HeE+zQaBR5P8paAVh+Y7xGosXC
GPg/Uz0EHaYCy4wr/yGgeMd3DzSCsupiBchjMg8g5uuhS1jyaSm64KlFCBmDgCJ/
Vbgdx3/Xnh8ySfbYEyO22J1/Dh8FgvHsOzdI2NYEMPdeppBqyyI3r1oXjvdVmA3P
hQd2V99FE80+gMyucf8eiuLhTukT3CcC+5DoVYknuxXNTgUHqnl8Jx73cEZ47kbF
/DmxfNCYPvx+4AoLjmZ6q23f1VAyw1gOYzCsayk0zLrijeKq7qfuoE2yIXbVteTC
QexGmJanfgEyzLUdxBFbP/g3Y5OKQgGpgE8uYyDgIchG0Ju/U/qp7uCsHHoyBfXu
ZC2fk1QfmvQ7WkHIbPjdFG03Y2d7AgsrgT86EVYfBG5g0K9rM/O7HkSr9a+o/9yn
`protect END_PROTECTED
