`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46M/oZuduu8XtLBBz6TAdmCGXecc1bII4pVzw0+RV/VC
l09WMQ0FDbZZI8jr/7OlSjRrlaxCAdFI7bV3086U0mB7uCkXV6F7LBS6NkQhcrIX
8HxqoJXSYx+Wau7Z4ej+CECUqXesxLDB7Asr4zUk+JcSx7CyDrwPw108+BDGNiNg
9VdP3kS+AzyYnuPSKl4uIyh9iXDNunEQde229v30dDIWn1fLw+O4y4DzFoOQWdaT
nypPwt6ADx0tebvc5lkthP9DEUL/zCnebyLCg41Sy3udjjyYgnha1Y4JEkL4eISu
tnr8ZbVoCUlG5SD2/dGy8w==
`protect END_PROTECTED
