`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
vIL3Gjc/co6JGHf5UpOqW1XZ2wNiPYrBLQp0t7Y6UIJdECknGapKkQuexYdTq44P
ANYBInJ+Z2wRHJtGEuk1gSSGfVD7e2gAW30ZkobtLnMpFoEZNtIj2GOnDnYVFyTL
gpqovWZUtrO+F+hhTwjrjy0DdfUXWGKEmiSjTi3RxR1oSN0Vv1z2lR/hj5alGw83
T+yO/s4HoLhj0cDQajUX5YZosifcHz7mFZAdY8y/p5KPyX6O+W43QcMmPRE0xYir
01k3538Oq1A+zMgk22l7Upng6/cgPSB0ynOZ9Q/J0xdFAkjUCj//qctjrYM/VIns
j6OAXGFIuEk3fWTOIfwGqe/AQ1lDdUFgbkYOU4ViKJI=
`protect END_PROTECTED
