`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKRyz942uERF4gsVGi9hq78O9MtWUHxvDokWQTwWGPLL
wqhdkHs1BDEyhO3sbdrXMGoxefuFfCus9kBN24mP24VUZxx4vsWfbgWjBlUjGSto
05eL7J2/GqRDUuXsud20LvCm9tmiRGpFtk9txy+kVYwYRWabw1CfpUS+JPko+G2c
WINyM8cSNF3lkBREHCn/ELVb67hLRKt6u+VMn04TrTkp4BylKFgeXwZJtoUp1VjJ
ugdly5tWfWgIXJFX3hgs5pUZyWv02bMni4XZL45XE4U+J1xnQghlAM9oiE62is6t
zIo7eBnSST0F2d/kNCD3P6hMUQV1tBqkigO2CiC1BrmEbpJH19p9BQX6IBcEUuGO
4Ld1nAJ2eHmhqszMraIgvIL2hPfGyquWGaGzdSSAJa982bid0Yq7n1uInOSIkxvg
E8bYxWLa2+AmtXf8qMkhGv7SpOYdMem7kl3gzj0cnAhgN/0NdL39Gi+97wbNaHIP
hvjAnqstLWGtPiSv9IrmCvhsuYOrp+ZubI0f+uKMVAXou3wAIfn5NeiAluVA5Eik
y+Y6TZo9lfDsj/rE90pB8Z5CCN5sHVjlDjkkGnPRzpq/vBgQH8SVpxw5glfTW8JL
zG3V/E6pvwSzxFtwOf3keTSZFI0MKh+BCYPzTzMZY7+/6klEdgPyLYvRGJfv3zs5
vwUOUyyDfpV8yrzpp+P/skw34t31zyCyeMubNIvMeXvTl90ur8cvXftmayn21tZp
5/BIMgpXUBchup58VPboXt4FMGclfSboSfH90vCgZ+F0BgIt9dtiD1f5JnRoZOVh
5ZI1EBdLvVjTYjklDQEmSA4hPC5B2PpxfMUm2riVX86S5albpGf5bdIuQUvw8FQY
kgH96xaTicN+ad+/+5S02Cf324qnX2hNKCz8KbEzfHfcPL7g+x4/KfqQO9kIUnrC
pDLPKUM5Q6ScgZiC4WeYlCpOC0reLtMvuqFNCdyc60d/MBtsLKfnA7XRXVA+Fpq2
9hxvx1mKYmDvFX3qR0MLV9ZhP9t6DWTfKxTIQkbtuzOvPlkL6FMIx1Jybm3wCPDL
e+pIunGoRLQG68R3rTDSL0nQ5R/zPx+jAga69E5zqmIvEkWRgy9IFHC1myv7QwUC
CG2P3ZvLUuSnq7+Dsq0y+0miQEh4yNxrxdMU1lGTO+9Tfa0E7wkzaOaNWgNxRWZQ
`protect END_PROTECTED
