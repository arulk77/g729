`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C7deatfxPDwi4lIAYGLAhPw8PMs+5CgB9rRO2QSK1Dkz
UcqyAfJtOXsil3IKnvUJLE8j3fGwRZbncHKQY43yzadXtDPNsHhDj3Ba7NxzX5OO
tRMVF10XXB6uo1EP2meIJjdc2gpItNNcnoGRmrgukW6e733M386ZYQN76KJdTLSx
3ERokfzi7QoI4DNnBXHZ69w9TxeIQ239wlxSaubYrKUimUCmS9H1aZmptOxpCiYm
L1jNcLb2g3x+iq5EGq/6JiG9GoeXCEsIN+rAsKx/0uj1XjZmB1paa1hPR2m4Om7H
NxzTU0A5+48l9XggPm/NabqDebGouqTOn0/EMVcfd5YO5CgfnEJz4ictruX+uxEA
Bjwmlj7JPnYHCY+GWb3KI5OSnamyim1Qpix4b8WXXldu9EhJWR857A4dXPOOXAZn
MZ9QUUm+S3ixqZsBzqigl3X5tmDXbimQU80xHTyxLmU9yzscV3nqVcNzcTl1yRh4
NXxV5/SNWZfN78za8pNvx8WIM5oTSjSLStjl+QS250KKJTZ2VpEmVtsqsCMb6nnC
lHl5G1+bcD0JA4Ctjkx4ruUr9BzOZX5LCOs1vYy9bek+D2gDMaXqRsQuFR2bE6zr
OFsZW2V/z5WvHgANaFXaMtxJp2ba9zBnsTQsXdMF1cCzU2VsH8Fj2Zpf7vs57fEZ
azBtk66l7J1ROStDmS4FTHpEW1JPjxgBdwPyTxWCSM+LVD0dsVPtwXRYR/O0lya2
H4WL+5/BjrpusyAhMQVLj27n+HdTjJzPH7aLyfYpuKELfw4fmoRAjBQjWVNHKm/B
b5QgVAQkzMLgKI0nAS2qSLd3b6E9Kg2f1tzAtQcEPrKGj+48/jcGk0t5R2muKQ5B
`protect END_PROTECTED
