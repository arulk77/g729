`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN54qpffrnsYaQxLAHpa1sq9xWUishDUbcUWvqIypRoIF
ZVfiTaooYSEcee0DEeBmFKk/UkylvUkNZcqZRBBw/rW5Q5HO4TkvUHdrFCFZjh31
i/LIqih0dC5MB9UaqjT3U/GH9ghcvRJvjmGynd5D0Lp4LEndZBNhr3IrF9skV8lt
ieQVj5KFZtj0cE5qxRfUcaXP5LhxIjtdacNY+hD75Jx4u7ze3ADv104YrQRT1pVT
MVfvaJXrIPPEeyprFmnCbP+WCXm9ZifN/YwjlUbRPyoN/HOjFUrQth5mT9PYoAfy
tP5EvYv8zZF5hfvtqpFhztWB0f4IbOueZZLWyrxhJzjJKMIZiHAT19V/bAHd89sM
JGxChsb9dZcDm6pZ/ZBrohTxQscpuN17pT1GmICOv5Rxn65CmLBBDdwa+QoOleRf
dMJJTyF+aqlh7N12ONZVbvoJKXbeWZZzXUsxX1YVBA9xCrTVK/6jDv1m1S5fRWrK
OjvaVHSOe2I9DT3C7vRxP9EmxaBjNT1EGHfpLWqnrTiQveTfAYr0p4BD+rON/Mhw
DsPCmOeRnULxumSrP2W0QHLEJNOxxbeoN3NTND9c5DMd/g7PLL7+2Ae3k4GrJaqA
3ENi8W28ZzwqNumxn/UX9mrA2AyvXrnvwTiURPfBEl5S02DPlIwxtM1hlvaRt2pV
+wOyj2S6xX/kVgJoE1qz1LQ1+IVuAH6St2T8xgghfdSApXDSLLpBj2Sw5F2DfIBs
qklE2FjwGvkS0LUVvm/qX+0CE1++DRqnVLXqf0zDQpX4BWmYlAbTCNbvqX6xBmWX
UYAcgpg61nQKkPy9/1WgsA==
`protect END_PROTECTED
