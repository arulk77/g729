`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
5xW8y8SUhgOziwb/AUcNm1Mp49vbj2PH7mfqrvkj49nWO8Ds+XgZl9xklEoLtblO
b6agixKt8ajdVm11vTP0tgw2IuT1YBshwF4tDtgWPqgMJAY6HweaGHPy1HeyHkrB
u2oI4ePb1ncbKxABI2UM4JphfG73aObBc+AVjUD278d0DJJp6n6vCmSO9UqyE2Ep
qMrdgWQFepZAO5e46EDSwP48uYR+va9Pht88tlh2x1vcY8i8Kt96wG3zEhPkXWP4
nPNbK9fZP6T9pTya9MSpOC5yDPhLfwOrBug7paTuIJ1s04KXJt6nAAaZno8IfQL0
4i0lYtMpE/c3p7j+Geo3J+6m6vSKSJbPqSxXW92yBdnCSC5Py981tgby+cHEETE9
4WpIgqfUAMkU3f8s9BXIW/j2GZR//raveMmwdDWVGdg=
`protect END_PROTECTED
