`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCAh906EZPGsEqNfdEzN09SDeoYJHeIWztw8rbeWDUyc
4MXqbmiTFEp1LYiQTjFS0BXt7IDSD7xGhPci+2fD7n9IIto4WPMOzfm2baS6epzM
zua7fZB3zfK+dOuJ4RpO1mlAMwpkk8fGxr9oEXtS494zVdqtpf84aT+pY2BBk6K1
4PVrGO3nyPWGLTaqijlLBZ51iZj9NJd2Z/LyAMDI7xNEVaKtG9Q2ghcGps1zRQRI
8QXhDqxagETDxdMaWBrmvGfgaR9ygzNEUxWcoRPsitUavFSw2eo+f9s8HNrIvUJ8
YH4BMLlBv6lkk0Id1isCOhvfFTh2UckYNseTH8vq7Cr1pwzO6S8ds9vJuwXx6eSi
AB+CFLmjprMZkWdvXqyFWgCLZsVcrt1pqTuGkbFJlgN+M29rEwVHF6M3Z3xn5ZCu
iPnbIok3dIogf/dnNCxeug==
`protect END_PROTECTED
