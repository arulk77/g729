`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJgPAAdQQuUKgxtO7fumkvU3UiVs6aTKEIxs2K7oWrYB
KW0jIqQvG/06nRZ5V/Co69GM3YodQpdYDABTnFe0Mo30SRDhfXZGN+Jnx/tHLant
dyfpkcfPPjPGqiIF7EN/Gd+0GqLkyWryRcHCVXBtgDo+0XrdPYk2T8Qfu9vYkV6z
`protect END_PROTECTED
