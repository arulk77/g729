`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2EBoZu9tBf8wFLCnm6xiM6ULr4rfFis6wzGtaMtBHnBC0en3P5gZuCi/+bTVkpFo
6aB/XWurjC0N0mqsAKKBZJ8n5kqcLri92J93pE1mT25VQdgXLUCeqeKJ+eXBk48X
2uR4Epl4f1SA0aqqfmFuKz3Tru/w/Utpcmo63SxD3gxsU8Jx+PkMV5kIrpZarSXW
gDr3ZCu2Naf5F/s/wy1Pt2IgEJ/B6AxI35XvDqy7xKRb48y4k15vu9FDgnRErbj+
`protect END_PROTECTED
