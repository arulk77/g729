`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveASs8au7mI96az4nzBwX2K0RaEyGe8fvLg8S73ghOj0a
/D5zk6cLkqkgY6/5zPonPJcH4FNvQ4rhNXgOgyJzSyPX4O1Llj2EAfC9PIU+3pKm
D2H+5lQ283dx1Dr2cpqRTNj5npSeRkTcQjTmEVP9jjneiGwwKHWIa8uEnMlSRB09
smxkVfJCNMxLpE+h77Nl/7b1ybyy0pfyC/d8/a4nghqiilcux71I7XxANYbgYw15
Lw7+SB37YjbS+1UcBPK/K20c0MIsLZ+LU8tAU/60EbwGAP8WqCZk6kYVR71wuUAt
cRxN/0oA+fDCPZq8OUWzV66MSP0V7654kgN5ixzDStW3WxkQ/n2W+AXbYPsike/5
YYNFRNh4am0oIkctbYCo7A==
`protect END_PROTECTED
