`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMD8gNZojmpEZnDnqtKn86b8S9xznh2CcYM2Knm61Z+J
cKWNVlWppG91xvUS2+SAhUE0m+aeDNKjDvffnewsJpWD4YIPU0f7FVNlj4aQ0yIt
6Mxk5zAiYyJGKzR/ZFp84jGcYYivRGC7sP6r0rVWTemgvf+WRuogRq8zH0oFBUqS
q6yPNvfqeTQCnhnt31pU4lqIjK41z0HRyM0ufW6XxXim9YgAzsHTfoquMR0VZTQz
dqiASKuGL5sNFdy4hvsMJ/0O3AZ24o/7ljOD6boKoumsxldJCkcBRnIC3HIj0rpa
9mKQI0z9HWfbCPS2fpJUYF0XFGXOzaG49T2EkomE4IoUIOhLE4azc2e2xQCEo5VE
W31JKrZ9HR8pxk0nts6QiAVpQX3qiflIt2Trkj0zJkda6/dQ0WKr3brNMKc2bcty
`protect END_PROTECTED
