`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
dZ2xupVWvM84h40C/BcDUzkmwlfS0dh+yuTHOJb/vRknqi98+8oRjqyQH1wwRa9/
f91G2BAnU4lRyPR2TRnBTMBkI9rVbwTW/gftezJUl44CnjcXjEbqh+uem7dGL5dk
HyVvU1Y8oHQfs1yQy8eVRdF8icbRVPi4GEgkXHv4qrZTMqlCAxDiwxMDzUPxlD3z
urDmNLanArGHBdwAbetS/n676v8R6lTpCc0eaRE1anj9TdlBDLUIZslu3Pbc2amm
RKulrUtUS9NTPV0yP7j64y3daOY/KjI5nPvDLCpFhFFRhn1KaWcayBUiUa4A2nDZ
7cney5RsuVh09vI3DwO53G2uiQ3R1UH7VMSPu6IvjLk=
`protect END_PROTECTED
