`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKTp2I4f5G6bbt4DB+K5KyZnkvmwh/AhU56eAu3sFiaF
thci5ci2dY4qCZ1BVOcSdpBti7XrDt831vOLJSD0uxTcpg5AcrGxSoNYaAyCMcIC
jSHls/nyjar4wXndYUagx7MMNMHc/Ub2KZs/NWtxTM5C3caick76HbKD1FCWZPQi
POxVaA++4jy6WdSTvoD2XzT2QVOVEEGGD9hi8Sw+pKJ4zrZdbZOvVjw7iy2lvq/O
`protect END_PROTECTED
