`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2eX2438A4/xkTNxycD1OF8OAMpJgBlps9e0GLEr73Z72IaWKkBV5zAQzuzXecNGO
4CTLpDsMSZ1FgwAPqdvmMKWgr5f/G/ES5E3f2dLlc9ksBQ7CGCbEwai1HZ5cREe3
enuezsUXI+vVCme2MrxgGwSpuep40JfzXS3SQX5XBuC+C5V7U5UiTzhUYODEDniR
9GjxuFEjE58xZxjozdXZqgDpAKTkLkEcrrugHauoHPdLFl56z5kybc3zC3tq765D
mpG8SoJgCd/0u1sH5qpQOTHT5nfxblbyJyoGAYjZo7hTmLVaZRAn8GQJj3IS5KWf
T9j15aVEpXgt/SgvymhVflM8Rs3dZjLKgbtDkzIMdPjUP2Bh+mUOULW5NfVVUSGc
9EnHokZPhNju6d7Rw5gnOa17hJgC7z6NJbYK+NrV3riHUDKuJN3v9hcaFbEuQwNI
rJUW9IdcgNO/CAjE3BG15efagS0fsEFO22n9YAz7NES3ZmGN8I/IoSZooRhO6kQD
ULQupLC2zFZI6/AYhangz2GlT6fMz3LF2yoP9UzeOcI=
`protect END_PROTECTED
