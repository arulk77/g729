`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAVu+Fxu9F/hxx3I7Y0aNqit9Pwu4W1YNHzHjWmMJaaPJ
twaTAVmaqNh6+Oht/Mo+nN4igZRB9S5x6aGyu7DG0kALt0q8gEUfpRvDuwt1Vzd/
r9d/3DnKKLQ2o1EWFQoy3Ke9l4FFrBCmzrgBzqb1/KRVFnxU6lmncejaVIs5Od5f
7Pb9oLaNEsf4dgiUqbvO3JEXQ4RGb13FhirDqUuiMvoqOd/7tfqS09yEGkqwMu6d
NI6y9bFxIjEnLOWRlgjyNLwuk39zrjJhdjFYZDDrPsbkQkaO3G7oj+N5SIaPcvhJ
1hlLGe8KNUl3Cz6F+H0iHRUwju6l0iRE+gYGk0oRPGFlFTBJZsk3f1hw0N/hOnne
+9AxxCPK3/8cjbyWT1chryW3i3HIcfSHItqnK59ZyXYsupfbKqgJlxNeNS3cRpTl
qhzvwxcdzcHHmKaL+F1hQMm+Wj4kmYOAF+dB2x39cUKG93bEYDjLN9zJteJh08Qj
vXCftYjJqxTpfv1Ql9anaDLgvqDd2keSHmazfg0llXUP0eL8zWGfRXvJT4lAJDMJ
XaFfiS68wCtOb+RaOu21Ik6M1UAWVNHa1J6r3KgXUJhF62vVL172EYIVVHFG5h8G
cfhIEusyHlpCjdPAUT/T/J/7aZAFl1NNQjNLujwz5wgLW/DpIrFhZMcaMyaYUb6b
Q+6EirDpD40zMTh1NkYGeWmXoadn6ajQgIM4kbDY3DoCwV7q5y2Ak5gWo+VPzeUM
vaxRb3TqXIYs6+GVVe2PKgGldx/DVoK08+YpFnKOPR+v+F2A5rDKpCvVpOh1c28I
zk+yQ38jltdUoqTjwqRdB1kX3XK0MDPgjGPUDGhJljdBOL6UbX1mIiLiej6sD60z
6XmWUVCYaFWscOM6jy1LzKvYc+k7umXxSMrG8051fxwx3FmQuhPn9wttz3t+AHKT
/xYwEFC7Q0LADf4SaIA1f7AszvKtkdi4p1DCxl1nUTvRskWOKCBYpHEnG9J1AC4d
iHVQqoSPgLHtlPlNiS1xEv+ZBsWPvW/HDQVFSWGjnWr1KCMFEQa+YiwH6mULj8uP
kaXNX4Kl1qLk6sJdoIOnnATpTHxDLAro16wiuBwO92QuOBTVyks05pMf0jveB6GW
yBZOix0U04MHzbgaadaQ2mXOfHWtTquIDQNfcS8ZbsesbdN94/SL3UfTe5Z2I9Ub
p2TjalXhzf0NbOnRSYYXelTxeEad5pa9jacOSwqgFSxZ08fMi0WNysMWiUgQceaH
yZBXOZvFti1lUT5ajKYsbu4JT92zd1/ZHYASyQb2A6DyO8lQMQyds7Q87H4p/530
WqOXYl2bvtouT4V/SxxGcu38h7OiFv+XJ9ocYWFQ3QECRwnICqDmXLnKImX3UDTn
S2+BdI2Hd91U1sy8xXi67lctT/umQe1ICcgKAFWqAQulFTxiRdpd2RZzWzPTTRlF
eVyR7sV+k9nWtbr26XqEOjHqiKG79Uq8L26+3xY4SNC2uKEosM1fJUyVXZNRkwEh
gnBi7g6ZEtniyinEa1jx3tz5/LjCQE+QdSPw7KIK4OQwp34z3Dj+tGm9HW382Viy
IgK865AAINUeZcY0iSYTl0loswe8MG5CCvcepbX1zd7ppM2ydTW4Ao+3qoQrlqOM
Qla4huVmfJTNxTJD/As+4r8fGnw7pxiQUHfwMCD7yc4pbJ5CKmUnVfeL5A0dcDG+
/GwnY0YCb/b7LWR7+L2PB/90tEMFpawwg3GP4UXfW8yUGPB9JS35NaWCyft7GABa
GxezxZb/l1zLinfyVMgdiIJBvoDzYH7w5nzinqwhz1xzsSnpENByTiDEz0z3BbY2
I6MY8PYqvijyYXILM7Jsy8NQEdl+O3cITNT5BRtufuShf4gaH0jfmEvNlP9t5wz8
9iSg5qAyitDXC9tZNGsluFHnxUWOL+Pasa3+rPmNaMe1e7Whyy7/VyGwTvuvtVqe
xh6xk3AA/COpVMugZN/EgGdsEmwaDShqrU0AQ6NGMg1Juq80j+BAKFp1RW9UHVQF
TgshNpHzyrD3sHney3jfzQ4tXj5wn0/7ZkTZi7R0KQLaUzjTw4nqKqQUBQZNyxM+
XHybTG2bGPyAnIPdVdCLkXkXb7ZcCz2viXkoi2d6rLh4bDVLgkzP3D8vXNJm/Hve
/J6ZKYCnib4WEV1f20r3AbRFxTOZX7ZoKWRJ872r5e0t36n3EKTLOMcrk9er3vaj
oBuH2I78WlNRAPU7YWHCHpoWiJwsv24aBNfUlz4YRcujTOid+Pxt2FNMroZfwZ9R
Vt8pBdXFx12fQTrWmY71hgy8/0uR6SYWHcqj9Juy70/dnvID2hy6opnFUjMGCkCL
g7+D6iEbFmITUyCrNbRSsaABtFjhTF/F/USoqfvjZVu8zqT0GaQ9xJagOmgZILPp
RJ8YfV8+J0zCRPAxrb6p6YwWDBddfsdRhQsgJ0xiiVvf/Pf4GLyA+WBJ63bbgV6+
tgicHOaB5wyJ6U+FIJwMm4JYGR3lscWLFp3ht8+Yuk2LiT6UwO3cZ7RF63EhlYn4
BUjfI/o1n+kV97HOvGPnmxj4RsxWdJE1lEZS+hs5T+evNTZKZcucq2f+oBE/i4VI
xJklJQ68T3oHHuHOLiuAuYCFOdrWAoc9+IrxHDYK8135vBXqDpcTYGYk0dD91jZ9
fEYnFXFywxp8Ax8ji/Sw+s75JHSVsO9evCNtdKDA+8yEiCTbkrkBfvBqLOG3CJlL
86ED552K6TEDJG5Q6lyWzzOGE9IzQMIw8x2tsIIGJXitG9ckxduSxYJpDsNQ6BWV
i5FtFsD+CsgJJKX33ebAsPBQ4PO3j7DSJxjs10q/XfQpvbkVJya7+VzRemPJmqUa
t5JcWqo8M7BFk5jtQKWCS90+/wgCfSXO32aBP8wSfEWdAkTxQyZCjH2B7rCx8obU
5SBP1i+l3JY/1scpBoBPfOgFgtANyWa0EnEplmYGUubpK1+24DVmzBSQtY7YqwUA
qWD05W+i8a1q+rZRLdoXan8t9IeQrBEjDRXJwjAmVwhHVp4/Lfv9NMWUFsvmszYl
yeBI4AZY5CYvNCMUTj0TCP2KajdxbwZk7Rj3cindgQ7rL7Q9lHoXQ1tNc07V2Tyb
dlktfZaTrcNl1sySOR61ZTK56cnv0XaUySj5BvMxAh7cvS7SbpUG2udFKXPkmjGu
bZ+qYxPRrwYkOBICC0VorhXzPhEda2uhUwgL5d9MU5zQlS6NY7EQXLLw7Pos3fcg
ldiY1lCKuwjRTr11I78ZO/FUtAuEuCUIHTpVtAQCe3cb3dXRWb1zTaDo1qLok7bV
HokuMbAZLbwNqv262urPqR47gBcjgzxZ0HqzALqRPAVhziAeSAcZSYhc4D+5jnGi
+0Em2rpsrpgM9us5qWWfrrahAvL6q5pmYr7Tp6qvR9g0I6colLwn7pnnWJ+9eWkk
bUvd/iSgvs68YB2khAKlojYCRrB3JgYEWZUzAIWwA5yUrw7Hxxt+k4TK0z5ebLH1
3k7C/9z6UOUfO+ezIKZKVh4hj+mTDKJ5o/Y6VYq40e4aCRSKAD82cd3A01UmIom7
xMJhlBL4zFgqxEysLHaQpaEUcU/JhHPC2Tm0b10LDsOt1aaHTjzfkSUOwIeh+prt
0R6nrlAreoDHjE9NHY5AdZ796ZsaHxe9Sil7gpFIGJWlXf9xNA0z939lXEi/fvX0
Arcoq2H5nhWX73FETSDNpm7vq49UH30pyfcKUTHhJ+owpnQ3AfyguxD+F6Y3rNhw
GJEadIuo5nUwCWiv5FRO6sB6W4/MiAZa7hC5ejMD+b4QfiUjP7qJAQA2ogm8Nu+u
W6AJ5c7zgBM9L+bsAVySEv6Ur0FP1s9R8VrOvU8Yxnv1Ho3choTF9bUe29JZEMnP
Y0pq4fQXitc4viaFFc+Z0k0j12i79ZOdoY2kLxTmocsEh0AmzuAd1I+jh9xmWQmo
ZX17FDFBpE5W8OvUFIppyJ9gzSf21phwuy7CKe7pshhEFCMDXGbV0DnS8qjIaPTD
8BVi9WMWcqPNoRlFrlzcXTHJQNyjPOAgPVEWgjgsg8zB8NGR4da2//eem8T1iS05
RyaXjR6avK+UDQOrqr3knxSgJBQYajaIOWe7rOdOYnKAdf1LxcViImFTxoLkzn4F
ysUKstU9RkgIRxSvPlMd3aM+X1z0B5UKw5J1zsxHXSwqkJBBaIK45A5++pfhKASV
kMgfv+5dDU7tiEMLLEhVQj3/HDq8PZF6VVvr32iIdquMoRFcwLvhfLvZXl+ZKfK9
4ZcQPVRTt0AMK6/CY7BdmfL2PF1FZHc1QZ7ZmZ+s/fgUiVnZGUQ/jvKUVlaENDfx
0WiVXnAjzYiAC+Le+D0YFnW4i7DROf2ZueKLpi5An9e0mMz0fwFqrVq3ITQUkksv
c1dX/LDu6oVe4d9WjNxI85lCZc8wShFYjmy0ikrnuGZUsfJnMt6lNXHyWB2wNdRJ
IJKxgWennJ+TfxqfZIRqhZrjSXfvwgmVU7roGDUC9wrjUoBDYbzj0s0bF1KtgW+h
FyHSwKxngzfKsVWSXWiImsly9/zBhx20b98PeoEKNfRPc/rxAMdT+vOgNxt8T7aJ
5X3QGa5qR0irzzCkdAT6XF0yMlO22lhQ1Ijt1bGIwJGzlUUwMnA157vdWXAq2T5l
wBB8Ob5O+ssdJay8zfRTiTzWj/qZPeJjhCQYFWIepBzxnZ5ioi3xEA99Qf2yjWjp
pWGqcT7Vq0lRMQnaPWIfdzJ5B4ErOc6L4xKVVMDe/E8kARvGwJg1muMoyeNmeOGd
Q2sx9sorV3Fl3dC55/YYR3McPgqT+8fbdglpiscH3hxyzWx0qpnSWb3r7zTrWTKZ
IHb8ypE/b9vI835M39huWRPg4TvmSoC5A6paHMcbejYXsn5sykhdXVhtuXwzL2lR
05brqDM4JdRrTgw0QAM9J8iidDnUTfQ2sQg3JLCSSt1b8WSqADvURI23sYRq8yuh
jOFZ3iV9dThL5LK+T4yHuUSLG2MZqib4fJL55SdeXPhUklTI8kMDwFsxTRtCpGTN
hP9VW5l6mfVbvy2KcvE693zN4Di0yq1lqQWXnPiD3Jwqyv+S2yN16eezQyBluJPL
KUFYuXgE16VndeetNmwvI6pOFXQR+Uh48cdsCGFsAXzkbD3d4TDlgtYBqeQozGl0
LWT3Q0zYAjGP+fB4Wx9zJPIFkst21myOrw37i+EzqXfksstCuaUOuOyeEwUBMhGV
3NLAv2P7hEZ34cpz2LS6/txg+xAP78N1dofv9bl4mfoW4L0ZkPKkae9glkY2yoi3
t28moKTkvG25sLnt1VvSpztPbdg5BQyjc8vyDq0i0tRHBmErx0C6cb+sf10hfecC
/35KglszG+uC4ZHFTfAro9xZNX4zgBEvKzMiGO8W4k5bHfniUOYTNuQP2qDQ7equ
rWb+zHsutGOGam3vr20LEq4cBpr6tK60XIKMsMX1B3SyOIA4tN36xK25llJZouEf
W90WsEyUyGN6j08ivV3vT/8bsdUJfKzwj+o2jXIjAM/P72qX8Hb7ffCUSuvDZUKK
pBjgPb5/4032RjtP6CG7ks5s0EXuNfgGLR4b50fdROrHiHn25Bb+DOpNga5xTmop
GB11fc7RL+PRwldsfq84duQZsR9Ppl2hWidHODck8E+UrlOjluTjidRu9fndI+Lb
OskaKNZiNWO0DNuNQcxP1bSC0LRW4+5ubh/jScxmW0fUeNDSk8n0/RqQ5BfZgICE
ZbZ+KDhh9RY1eNekzhGQk1cTL+ox70cd7quzIAQ2r0WDRW+vWJ365YjJp/rTf+Nt
e99LaKNeWmgRF36eWrpnK3fy/gtMtWwvPq27fgrm47d4R8D8Gwnbo/BNVpK+DgZl
SNtWkXW2DV9O0XktRrcXuvGf3DeCJjUK5+378HZuRESNqbm7SLT5JDnxLP36RvFH
OJ+uZ/651O/JQQGbbddhmOfhZlnjgPG4dvRDqYl20FHwdjrG3Q9Yg1i1hXyJyucq
etK1m6dg+YAR+VAxu8OXQht+T8F45fb/oeK/8jAOCGlEyiyG9OA5fEZL/XAJBMqs
3bj3o0JqamiwMv6Y1G1YohJYWQmVDm4ZGlG5LmwFy4OJo2PAAQR2AbgGTfGSD+QP
WgvmNc5DUukWHD3TiNSaWsAfEcw1LMOXwJGvsmfxflUeijqw4dpb01WcEDVLKAi0
8LA4Y2v7il8hi+1ApY3n0WGcn0/aGwRHEcZDjoMM+U45VLThWf25w/mHk3v6CfM3
p/7v0YrFdzVSlpcqbhqDVWXy+zki7OVhCtt0+EKAPtdYpyifOi13Tv4YtiM+pE9R
fwkH67ZMUUSCeNr/TsBjiYhxMkm7x8YGgWIT2a8257LqgtSWGc5uTnzVsgP1KCMM
gCJb3d7y7NaZyql4Xze+cKdeOj7KwGCW9U10xI3ZjSnuwhib0agEBVJXpkbWCrCv
Cch8JIsUx5aY6HpYrxzMK9SZJ0UUiELMaY/MmJZN7JjqgDoQh5a41GRG973knBRB
Q49iLMu+kxag8mJYR+KAY8JX3+4ioB0gELznfdm8eUoz0B0AI2raUabw3Id/l6qO
jO15YtujZwMDwqnVbDfw+gYypdG3eKPwPDd40d9nXHtHfPj/tkPr0QCJIGm/RsAL
FbgFrGADW/cHeEXOp/HaDz9NFLYJG78hnv5FIF2X56PvDmCBIsIeDkYjiGagCrvs
z9l+gaOO9oNUBAdrygljZAN+qEK04PhJn3YBeVLAwazKmgJfjJcNs+xDfBvVmW++
lj1iRqxanEHwdJGAfpNvGK+DMissp4vtiOKOGlPoZGdx/iSZ64DEwukocFtPKSqp
+zUeFzNad2mjqoPPF3PRPpnRgLR83fl0MSfTlvLHG+NDnjj3xew+hpT5vfN7E5Ep
xl8dGXP9hBjpbAlBGChwzEv2UQm3S5Zb3HzS7uxqQynLpPIaTGQGnGk58Tok2Yrt
t1v6BPDUTKOWjCP+vMOQ7mjT8hHwspb/gBC8/fBv0MYvZQfpD+wemb+yojex0Ykg
rURqdXK0xBPS11i8SS7gEJsiv2oXB65zTZ371aFg4swLf/wy7Trp0Fq3bXKLNsly
6VWWBVhFDKIB/6R6GW+CPancqx+C6/+9JiC38vRrdhptH4Yw3GmSTiKLrd4FCtkO
16f3PTGv2N7fn88qzqAjxZKVGURH3rHe3iCVRlqzHc2JMk1/+Avim0h+TbdqTLat
2P6mHDoaaOAl3P68H68rdGQVcbob8xiWKiTr7EiOQ9DC2H6WL0foJY/n4SsmPXcR
3PQSbzqpiBdvXoeOvjPXZ4gERKJDEXI1KIUy8n2D5SonKLCAV9nLRyP1/QUpGj+z
pEFsnZ/YARYsbZkgKfOEvYsnAU5S0MsDBJ8tP2wTsiVXCtSr5xpJWqTCowc2LE8y
eAibfMMzhDTwcexQMu6/l6sEGvG7hpN3RT3j68/Fdw1PyOrr/OzX5T5BJMsWCK77
gzDdv7U9h3tDPwdwX0fkXCZIj18ubVp83GaDoehV1BZD3fyhk5BzoKA5fySPeDta
3ITvBsvXPqNXa5G4G6WEWD6CFCzly0irIShBWrechFEsVbqQeNW8C3+Omxx36ok1
zyc+o8kNUoRjyxmQjaZkNT6VFfC0u5uSsEuUIes/Pq8gkqZvxyz6IMmXiZ2ATvrp
mkbuQeUe6h1w8F8V5U4q5y9G+J27sbgi9yiFCmL7O+AY0d/nErBdO1Yb5TqTRBza
LELrvPHhYiWhOuEhryHODN8SksLXXnsi8i0lQN4NEUOrsewazMVyTm/KSF1MVU5L
fOCr2bWg4KR8mFtEhmqel85y5QjTcpE4cp7MXuzSnQBNq6ylbafpVZU+SFH71dgK
BdAscii2IBE62Uisvr+i28OQozFFHOoO5aqRwEYhXAx1afPhDJmFEBLwZ+ESpB40
+7iI6+QrP4CbHZyDcjufU7SWz7ZQgjOB5cgU2Z0pcxvLcs+130Yyuto4N322Nb0u
PfpFEbOYYbMwbVwkXBFaWTLoertmZ08AgDlNBlkFL5c74452DxGWtky/DXm5yn3i
xuuPJqMI59cU+nFCETuA2y3RyH4SfuNoJckHwIIuO5SrlZEiX5BFGfWgdUoxoeLz
jt8BdIay9TutVEY6JLJzIvPWFr2HMbfCExxYb3DYkNfDzNt+aO1hfcHRCgWS3AL3
aR/lim+Zxg+mhEJbVQVjUGbxQSrbVX6doXn1TEAJLwcRe9DHFLX5Xg9SRBufvTnu
xElJ0pHLY7ENfIxB2TpBi7dquR1gYEr5upNhyiF0rkFad+bZEeMG1kwv+s4kAjpm
D3oxnNunZ0CppLWUpynbWGv601r57Y0k20CAqDsqfw3vyTle/l4shyuFtgtkGvA2
tP26L5j8k1p3/e0zoM8cRNk+jSuybUZdGNg6NNSEPYC7fq/T/ELlruRYuuqoN+Un
wuHY/sxlBI1BWG9L/e/4cRZ/DRLn8bxzXVTrZcik8zftavx+avEGTMN5HpHSjwUo
OqDvEsgtIaCdk5Ya844T0hYe3P+bXT5leKb7XzqgshVmS8ttA2iz3g5oXWE6qOXc
Z9V7mIo2spZ2UJC3NNTYbWYO6cqFjXOuD6ywErTIH7TJRjheqoftyUQKQoeVJEnr
qjx1+m/deAOMAx8/qg8Mmyrd/Ti62CHsC5r5IF4FYH4A2wePuqu/tI9NtGSsFuBy
LWL1kTykPxIBta3jOZl5xDnD3wjQ73j6vgJNeFGVCiuhNF24tTFYY+pb2hJAKGLa
Ni/HtkzutJNJvXjyhqr2y5wqHLSEabk3xqS7/yFchLomZ0TNdZwRkOQvfP31Xe95
rKn8hyEUK+AN8+okRH5IPRun+B3zbQFVbURgMakSyQW6wASN7B9e+1a/N3Jw0MoU
dEUjbtqR0gG0cdCJ476bjzvggfXK2WTbsKxFNKCTI4TImHNsygW+GM00/mmmqq7i
xfNBH4CY4BXkeIm3/rrdaUaKiMBqoo3/m+7sPwaAKwbdfDi6yId3k4E6lHJvXIOp
ZxL2tM9+6WPnI1V+mbdONKFJtdV60aX0hxlpsNnrlv5x+Qvwclss6gpGMPiulqeI
8QcwZcwf1hPL6EKm3i0O+/d57E2lAa022jCoAgEvCjAcl+TtmCoZoZtlL5pJ5G+7
O8/oRnMQzUQ9WdR3TKl90s8IoOixmowEPD/uOXAgStS5pV3JgzLFxNFggBvzl5Pl
ZmCrGWMiPURNCuOK1kF4a4AOF26GF9zoCFlT2Inr4kCnFs08+b0USVqbYnWbjqXD
2ukrobuddeWohFvLBWmEjKPAIHQDYx4YuD5bssdVotFSUNKpkU/eLGEjGxExdv70
doCmT+oIXV3ev73AXftjU5wwL5J+Hy7gTuuhvuY2+mBGTFo0z1le1q1DsZ9y+Jcc
Zjw/8mMUHsC/nGmLyLB4qSwgem/cj8I4elpf9JC9AyRUGKzYB5zDhHZIYlWC4eQd
aCW8Pr1+nD4ikZ46xmYTAdtPIGpsyXFmE050ZfOkkDWQuD1WFXOL7G6tNZRScgKD
EsZW+8xPQ5sSYvb7fpnXP9Ly01F9wDa8qjrHVqgYLXjI/SWMkhF+JNHBIUTkHMCF
fxIqa5U+vP+JxnZ6LK4RCy7IFreaOFPkQbhQvaIfPs2gQSmZsc7uCcXwBkTL7JUU
SjYKMB/OiKfZrTI5hGYBfJxKewbLM/FAYLegeMOVqxzjQjtWu76wBn2F/dQjwrn7
mjVSTu0rQLelhRuYfrw/xwBj8l0SolHWfaMJksoMg50AKmpvut9I5wyGK19KyvdC
cW9JrSbZ1Vj1Gp1FBxk6c6wfdq9NYrSmGiUzkR/4ebDl6EtkmK+qIoM1QNCeVy10
XVKvjpn5+hs1P0e7vTuZ8KLsSse7FI1uqlZdFtgdAPP1k5qjnPoCOpSyl5MZibRe
q/A4z+wETB2uvWB1KyXQ7UhCHq4iYLc/4bzL3NCEex84HxsWgqzD8eUHGlje9gXe
ZliTcoIwdZ1RY8ToWzOYG+JbUVld7mTvXKFuSr24YMm9TpaY6ibv+TcSz8tPC5dX
UvZZrcUkaVCTKbjYxSbPlm1hWabUQUYORHxlQgtqyHrH7iY86fZq/xRJzSsmsQno
FXLLrkDth4VpWWanH7R60FgIf1j9jucSbLwdjv2QTaJBpTw0QHE0xVMZGdxyPvA7
vPGpm720mfVa2roeEZKcbHywd4IrC54rQuH+vNaJ8EC/Pw6MXiZ1zBCDfXPJzY9m
/OJaaMst/Wbd9EKxOik/6Q3MQIBtOo2c55akwb+NNDZW9F7+dl0wdcYVMgbzmb91
08ZFrhUDmoxYshkAdKl1NLgM3D05sp5fJB9Fcjpdrv3WAn8vBYhFwOAX5rXH3tgP
/rRXsYC3zGUIU+DUxdJ7XAnbXeDbnO/DXzmkc3kywEAWAogijTqYBkSbJwPTROi7
ImfAhABAcVU0FGc5wV167scOD4mGeX4bDEY4EmZjWeW0WEcQgen+KRpJp2ieBWC3
0A8pbFdkjMqOYxLk/0ycbETMi9StohSepDRw+bKTtz/g6HPDdd4yJDwTSQuzThvA
TBYcudNQe5FbfXg0ZUCXfy7epJS717f8P8iw5oB/VfhBeIJSXBjR/HzkByl13DO1
2vWRiboMImx0o/2MNSQjG4U7erPW2dyfS0kZZpEWAWbg8ivNwdxH5pmnd7kPfrHw
xQ/ptMH0Dsm7S7jjn4k8FwKvVXmOV39sq+ht0dRLPCDLt6d1HGs1EV0YDHMtNwcL
HpzkLgcj80lQrBCQNYJ73GCrE3NjtNB5l/3/MxDP10ZPC1jX5jQZKYW52hP9TLhI
eZP5OmniIp8GeKwDx3GGCKHzm7JxLN7gNTMYgFiPG51IvYTh9xoKExMyJTMHp+eA
ZgWuMpt32v1uDcxFlZ9swwQqXk3IHGtTXYoGFjKhPUauzatRnz9fsIFakzNDRsyX
EDsHuJszooHlgxREj8SdB3rWMpEPjaR2/233SoTRySBMYQ5GCWtXl9zbNK/hoLwE
TYdDX2XQU5RIUty9LzvalYw1OSC8ZF52ITA/q4hrCWgQC0NBpquGxFXMcuG2HXsb
1hAgGKIkpzUNEOhyjk5l/0GUfYNlZXG3a0Gp6B0UC4Mp09I56YkCeKfyNwKebKP5
2afabn5aEsezbl3sGI0eRRN2dysqO/uMUV32f/zBCtEapZgpbZnHPe8BRIN45WSN
LCQ0w8SfOlOQ3c3W+3LQWLzjlIddQ4kS9ZhutI+WaOV/DhmNy57+jbGoEAg5oLUJ
nEBBwNsIb8H+ZHTvRFGI2HvVoGMaeBY2xwHqw02UeAOYobHHN25yipW5aqqnZNdP
YawKUcuIpEs6f1x93EbB+XCLPZaFJROT63mtHOwNxosvLu93nDrh7tsx36ylo/LG
lmmLvWjzJNK+2M4tYaa0MJdQmSaT78zL3HwkrvyF/Fhzhp5rHFaVZwExgXW6IVVh
8DwrMVUOugKS0t6yv3fn2JjurYXyECEhFfyNIPouhfVeRj/SHp35Bn6k0a8iHh/F
QnKLNiunnN14p1kcILCLwK20JkyDrOzTa5ZFMmkubD77lc+MC83Qjq/vR3O1E5fX
lCm/w5nsI3x69JfwVWPA3LnCMMPowcqS5q0lexa+RIgS2ER086BqJ6cJuy7rgD8Z
eTQddVNzQnFqLcTqdaImUai7Bhns04s0ZSQu1nyELAk5t+dHJ7NtNFfyw9tzwrk8
TwitmTefWbTNYkrnFM7Nh2/qI1BimVbHEPeHuJUtvMXSFsupDmBeKvo0Ouo7eRdz
knXUOaG5mF6tSI4WPOXjkAAyxQts7FH7maMuZb+kZ18O4YWrywLKCiQfS+NuOR+Y
dfWKsYjuPwaHxu/+IoJhfw0v5EsW02Ar3uBSIU9V71uckFpUceF+onyG29/JOxzS
IvodNPhDsOxW5jH1g0PKl939YGp3SbxAdmvFJAu+at8Jd9qXC0aEIuJh/7/1ZvBw
WpM3zisK81xK3jL14w/VAm0LWxT2Af1uSksPyiEseilHfx678nFHfHevO+eCf+0R
wPW9+M8M+XS3weC6pZf6UMs9U7mDlweoVH1hQyL0Rp8OmaGdRC6e9PZyvV5dZnyE
NEj4gO5kAhv2HP0U1tCPW9LmYoD/bGc6T/IsAGRYUOGsg4TpHSL1LcKWrQiXA6wu
7CWYNj4bHB4rP81Gg+uXxo3di1pZeYk2lR0S5Lcm8Y/A0yWvEWQhuhWrxH9fEZfp
2B/PxMMsnXhN0S5+Uk1dRD6n3k3AC4ogc12oAmAi/NNPZcUqhhXU+XIN0vbHxRlt
D86h+s3ugYnlBW/drA2CruNqCki65Sg+IVifhyuGfK+fNHmbGqoUCT5f/4sfVBu1
WGDNQ/QL12EmMuOjrrEyMKRbC3dLmIq7HT+v+fsnp/DVA+HcQe0EtKw34AJ5A6vU
nlWaIDdlIH4S/tRMnfQe3Nkrv67hLTG9hU0ksDVnAsMIkoWAyA4l00/AjyxWDrfV
OekUJ4mBC1Z3EdNli5O47H5GwKYX5/BFpct0GsXNwBqbAbdzcMlbI3aj1HBDmfWs
lQqrDeHlE+mBLx0L77PmkWS/cS20p6cHm/DUjRu72k7GhqylPJGRVnxMmcEhRb6G
wu3s/BAMhSq3ze6sRZwpc7Vm88PhW2MbinAa6GDX6Ji6zTre8hYNyu/8GCenZhhb
5eA8ksN9pus19CWjILlsSL8KJw3Xn81B0q9CyVx9tV7oSGEZUUhPCK//u6A8k/0h
pgDu0RYR/RyVuEfpvulGxdhCJGssd37vbMrH1ENC9VEFRtsuu0Ne/OD7Q6TmGTaO
6nFEqK46+Qxe2HaOwn4iBfYqoRcUkZLH7IOIZs0hSediz4q83I7wd5aBFcqUEx07
zrDjyKJtyBXk6H/For1p0EvX3QfC7qisrg8wYiSmdSn66teeJzo1GI/8ETg/z143
L067O1PcyLKRBkQKK4v6xHovUvzR20oeGvgJAnIie0U5l56iECwijfyrhprJpmva
8My3Q+e4FGlE9MfAFkCUjZqB6FTYx2P147L5h4/ZddpTrsdTGSsQAdRGsT7CYuY6
RRz0szG3jPn8N98JpvJsuz0/6GtrIofO24dX8bcF9l4txfFlhBIV1e59HsA0UOcJ
Hob28NY+D6Y9Un2rDGpo+o1M+dRaOXmp2E+H/fwWi8UVcCPzhlWe+fvaOO0ZFoVr
/m2nNc7oNnw5sQz42xydTDIzIQQz1Ds1wORSdEYNesT9zJc1Ctz53o6tR54vOg4n
U87stMXLHhXd8QZC/ZrE/RHgEjThpJgpAoo8wYXrev2a6mN1GC+m04teIXVMw3NZ
AAvXlpqoWgnOaQ34Ef5P4dwz1EKVUAcMz4BvpkraMxhCTi+us4Tey4l2oeo5+bpx
jrjlX2naeGx0u8vSd8q+1ChfvjzQ4SqxqnYew/5WCBd2g5S1GPmG/1ih3puhjQb9
gETJ9TJcApFttLvLhIp0+t0RyTUFwPyNC90PXpWFAb2oeOmwyPOLCitCpG1gaG+C
jBPl0xrhuBc+c/QoOeySL97f6siV8ytfPlsQftuITp6KPblswLwvX37Xcb7bXXjc
eu7NIPAZF9C7X41y4wLwmfdSYMLgGnCR2mgSm1r0IR6Zeijx5HXCEGpCQdTjecJY
+Kel3XusKWnjy/XYfuhxrAEEIiya/CsLTNERL64wIJDMirz2KMelGT9sD+RkNsth
nJcyzldVHaPKEtZaHaXgH9EYwyUNECea57/r1BxTgee2b+2M2ejX6271dGqyeMP+
AF07uL1Whn9B9i5Tp4IL70dwsu0WD4kTlf3AS6O2P7DHO/IjS+4KHoYco/IFX0nb
XSJSCqJ3rRbNU81p1MyWCPlVaHGl971UXzdYWXTnJDuw3yqq/cAaKnThygIDfZgw
yxkkJ/BQ+7lK9zKWe833qWCDQpcOIgDyeTq2muIyZOjEWHisHDH6PAVWGifHNrAm
99iQ+Ccwd//cfLEZCq8r2ha9BY8VqtkhIZG81+wU+GowQu9PhIVKH7mS/YVBHHLW
JB5xJaHqWoTyWn/mS5oy0e5yNFseZe6qfSwRv3Lu9irgF1W5hT7lrYT7D2N/Wn+5
qVhFBKYoLucdpdN5hpxpQpNwAps1Ei1sSQcoRhmRTn9qVsqzKOCtJ3G9X6S0EGZN
Ceh+cee++qbjM9uE6j51L8eAIqK3Fp2/N3Il0aXz986dvW777NqfN8s7CiqxOQFw
PUZP8zJJgVEQTqyPpqoYqcKM40KGj1rBhlgLUOk0NmaB+2HayF95mKzFNfGCuE6r
Jo60jD6ov7CehoN94DfIZLqbAoqmj3xRutzycclsefihCkSqk5rq/zEYAHYrBUE+
FMGjvAI8DvbU/0FEqfc6y84EtM14sxWOUPxfTVx+Lqd8h8fYPXIxqliITuVka5gZ
QqRgd7DfEnbtf53MOyXiHuP3lAFrpI1QQS+AASclm7Jk/fpzgrwDMmoD9Cwq8/o2
KJcQO8x/BeRNBZi7udwwbBXSmAKRKSO/s/S3zXsqMM+oGWrhTN+zz406YhYTVR1j
WOZGVL7i+j+y85PjiS0zP4a5E4HqEgOo6ynWPR7lcTQuUU5A/ecTyYwY+bRZV2Zb
+5ofB5t+7fPpGpliWR11sBms/U7Gajcjtck/hzNYHKzcw2+xtzsi6/K3bn/baCz+
ROYTBEJdTqcpNvblr/fAcW6Ux0MLCff6YWgar9wnv1fZGNMs4zYyoyK77UYpxpqK
qZ5TKW72/yQ+HCLlwDpvH6gp20/78+S0o4bWOhHogAM7RJ1p37QIP1x7H+KA0gFF
bZAYnHOpok19YWLueUbmatR2OvEl4CH9u6Q1ht9OOVceppe0uRywAGIsP/AZcb0v
wD/Iu3QNlxPN0PhYU5AocrsxUvx/JU3+57+o63MuMGYcz94jLLmthoqOoASNWeAs
jDVekZYA8X1ECoch8/Y9XmVuSboPfRkAJjSS7sUPp3RDKQhOBIXU2OCas/3Qf6v7
Qwosg6CdOVS1wuXw3FNPP2L/3V0ODBzUGdeIXRTGKmuYAMy8l4qwmfF1gULJvX8n
vZ6S9sfYvws10uJfSzmWaPE9BjtFDNnqNEJyV9JICOJfi+ltYiE3udFd3mJhqmkT
9/Yh1u+EUtKNapik54VbeLXwoOPvVZNL7VZDTetURrg2PYL5zA0jjmhBsu9J4Vdz
Tw0419PPtHF7ZvJ6l3LTHtG8nb42SHtw3J+M+mjuAfH4U6z0r3hwK8SKgy0SSZ9k
Yij7d1fsdqGGxHLlxkR+XbYaJWMujVHMwAh1GoUY8Mlk5HJZDqe0AKzzCLdWfIgH
g3X3EEJYpDRKbvefFW2pUtVq+OQjAAxb8xZvxuYPGTepOZheJfUer494Yu6GKkNz
BmcGg29A2Epdc7UIucliJufCKSNIXPGu5Z1Dw4hdVQbfYi8hlEGnAG7I8e5WzNp/
aKhV3go5KG51dGp8DxIdDnBEZPYPXZ65cE9Yu1jhHJocltBYWW3ufs8we6VQ8neQ
SW9Bt72QLfciPL0AOK1vZOCaexx4eqK3dbWKWwZiZBKV5d5EBbzLAPdQtG+0DxO4
+jgVSe7qYXXUl7JJKE05S+sAAGW8dBA4cqDhJmfeKsF+rLyvklSngE85LLK1OUN/
39Fs2g8JJj5tKmSn6kkgcIzuIYLP09DOEPoX+DVd0OEqoQGOLePF1imCdloFy6Q/
24u/pFhVbOSIaMjabGRaq5DyYDzWC74gWFqPC7ePjFnUpdkXiNcSQ464E2mYtkU1
AfS1nBsjej8cG5t8qZlYg+BgZgU7BK4aMHAiAexikKlAqKuOmcHTMQCE7pHJ7zBs
tmO/K0BatufKn71+z9J2QUkInPJi16l/8vRdPmsGdSPGNOgQiIRGxE1eQYWhfL2g
gGmFusoXKwUsWKN6UsCwsihhCWpORMC9ktJlisVNbv2c++W8bFibrHhJum5J5vw+
NA4PhgOR4EtsbNahj2655ke2DyjdbMZrwPPtOMTT3wN+VY+nd1NPUlSsZ5iAlwbC
Hr0Frzx3+7IhbRzJ44W5dF+ZdeHLz8PcoXHOUFfQibD7oP/hSzouq0w3x0tqpUWq
ZbQlpEG27kS0wxXCZsR5JRqwdTyLyh59RijCw01nKdaSxYDwyZiwWRAXwKqSafv3
IxF+hUnWbIoAPtS0AC6GGDQA2lCJLnbKM5sNTe6j0FkxAjfCLsv202pv3k9wiTXI
Wob56Bs2kLaGz5XdJJWpTuyrS0MnPHJWBKX2B83r11AgRx0J49V7/xlxYaEqr1kP
NzRdFxcialWvGpzr6DGK+yFeWrhcaEIlUDJHurD2gTttS9WRmdQ4cE1PcqNuBWk5
9dRl4DohcAOzfox8rfbTRwJm53+Klv8ioY5ysDMDFr+oWyKq2DnuLaws5XDAarat
oQ2xOQsWLQU464VHoEV4ObYd9iij2z83APrmFmV8eYQIv6vVWSFq7qrfTnscV5cx
DHnyw6X7ClwJX8qY9+KAj98k/3/+22F74AQv1Yg6lwB6a2EEQaPbUKUufqlSEwDC
7GdeJk8FJle7YFQMCluOB/dTPysxf0ohNP1smaGjREOratxq7G6OXcM/z5UAftnA
a2fPgbrTWppLSHs3xzc2pmaDKzmYbVJAtRvHPL7CpH+NYl7V0nPVmoItcXzs3261
n70oJq2K7G+iGtzeH4aBRI9RS2aYQ5vNKweVePHpZWkIbZ36y9budHChgpHBfGhE
I8czLpy7SNQPif1y80ZPmfGeHo/ly4S4n+AP3F54t997oUuZkHpjeq9s2Gcpw+d5
ULCd1ZrbLtqkkYyWUPG/87PBhm9fThhRTt64SNAHtfvp1MafDuVMIHZg1Uk68nw+
19/ia4CqjB0z7/S/NAFLaJ1ZYDnmC3syxelNR/k30ZopuutBI0sKoytWx6Mwi02B
22z98R6s3/ozluTto93TNjH+L2fCjxPjcPmHsnXzm8jJ97sHVXUCSaDKDD589YiB
AgTuzrrQ47cxL6WETAynbnRtjgmpGroFNQb8BRUaQkAmDSf1YHceU2sdSQzeQSc9
kOQahTnuLhMqKlOLovpBlhVxcFwfvnB4bbdPtZy5Zuo3AVXXAfZbrDwSRpjNUCa/
fmle8SXQ5JV4vjH0Hs2f0DJG5YIfBOlNNLoxYZYvkLJw6GLK91ewFrz5CTQ61QD8
EhcXySVMlaDqd3eFmGdow8Hr1Bm2Q6Zb85xk7Hi1OMnun4yo1F3pZ9ZeRa6bFWtJ
FLLkHRdmQA8hS/Feg4DI/yG1e5sjPqfLM/msgxsbJIYphtywWb3uLPxewbqlqmaA
ZbbSRDg2V8KPxpOMnleV6GGG70GXgKa5tMvEVvhlAJiH0W/oYjl1+Eq2cxAblDr9
fa+jDKWqVOxj/kjugr70iITFG3gj+6yrQvU6YnNOHFNRJFQzg6T7AV2T+p5g8pvu
Ug5kGO6mjKiVQ4cvgUuXqgVFGwfAxqilRqX2rYZFRe4QH6efsryCL1/z+vdrtywv
sD29t77Z9sbgQYTEpNA8M/MX472pUEE0t9qTVwBUEIEMCp4iHVO65EpShlLjwUfA
m4WVAVSjq9+CEN7VoiyKokK+P/MxKb0CeAVmUNu6YTK5cSlg9I8wfyurMktZhe0B
xUUehSSClbq3Q+kuQbZra+XIf5fQO1+hf6CBWef2GKXSmQXWVGWLGOdDhn39RE7K
iUr2B0WTb9FQ/VSCkesCtDE5OYKFq35/um7dVEmkELrFlNoOlQuglpqZcKHJhi5A
BvdxrwLpXZTlLclHsHWjqOktd71MMA3CPPPVbq5+fMMS9Agcc+//jm+cmS7xlu3t
a2R2Ru43hdVzJlLkSAVLevj46lpn6GOkV7hp6QdZDA5nwRvq/4Id/dBqEJFVeY7y
gSHMecVVTgnjivbERzz0DVGAgChfO3ykpj3SfvlldXavHr29PemJ0jm87euHuYjW
3DhQ9mOKYt9b9RsHNNMWJZ/3FVMHyIP8VaJSrNdxX7wfsqHz7SmVXXqTO6kKpp4m
7Wv0AgHy2PgFqBcolA0n2gkt6Xe9e+RDylQuOqlLD/V21rVHKOKolYeYiQAnPs+k
iiNdj8c+nrao1Y0ggzpQAGhEqO+bLMKPiHL/h/LLo5T7aPgruNssIVbfvvuIuEAB
1GU00D9CGBBulI8SoqwQbhY8jgMoTjhgNU3JxHyIgPnQkEqyrb9K171T2UV1ZOUN
qhdQMYgc+PUGYwiS+UHVXp/HB9cP5xjDylBuOD+zqbeF6YwoVnd482K61PlqbAcu
AGFvqaqF+ZfpjSznf49Ka24k6MMooXqkei+zs57E6Wvgbgut/y3IixrzzQ0zISdf
It+6OsYXaJ6wfTeh85AEcRpv/Xna6ITG2PpddvK5eu+rF8nn7ceFXmj0Z/uSYJXC
mTTBV9bTqVQYDKtSH/Yw4A9YTkrYUr7cK6Iv5whNC9VKAVz5Cirf9E0h7aK4ppMa
SFSfIQAIuLuhOvbpWA/lsGlUUEoPH5m8Bz7X9XYsKu6exNOJIho8SLewsWVm6phy
7QrikqqrRgDAFVK072yQYss4p2zIg9RzR4q94d3RFcbneUBxobKFhrzWALEzokoQ
SGgsb2bJxNADiaMr7gs4Q7P5YfS1BLlY8Oh85DrXz1DeDMqHUKSyj5P8ZMbWq76+
qU0v7PKhLEYLR2iD3qirEtdWFloO/G9dFvas0a43iJw/o0o/xSk3VihSrs5NSukS
ohE/tllfb8mhTWeqCmzvYnspTddDDqxD2Z0ipp2OHf2B2LcJ9Fry3bvzIICbQfGp
UfburfZAgxya8rpfuuTYnEO1pKgY3kqtJPPiCbnMO5qhFBUG16oNoZvaXz4ULTrG
Ao6HPnJ6jCbo0EuxMWkbncnPgEojCku/GO31hk+Kc1u5LGnwMWy85DG5KClmMBn/
U5tPqyAcQD05GEmJEe78RtWznJHg+siEzwG31+90Ill0YXvZPUWU4f5FcwcPrnxJ
a0kogMCCrh7NpJX6VFadlJhiki5UsNZPuQQOaU5+Y1atkrKEwGmaGYXbr74/jWJq
PyF8SJ3h3SRAL0Oo89vrv1a20tvAWKkHdjJkx1PlEgu6sA/5ZQWLPKXStVxFQK7L
t6aIQ+wQWP1dSgBQwEN5qdUQzhD9hZMcYC2gTRe4qlqVeVBGRWHNrZHoq/W0Sbq4
C8lRpwtR+51cER3wehHsRdD31Jfa3ZT3B/QfyNQfTJnxSk9rLxuxRbO49GqlJNiD
H3tAqxasFkuF9sEYjtSEBB0ETJ5VHdCuoVQTPxoo/5BjIkB3tYd05KE/oPyor/Lb
JI+fD/2wMlsgpqL3fq3kvpzjNdHAMd3apIQMRVnkhgSx7mwMTCH2o4fdg9T72KC8
NqDDMWLwRAf4eXvjbok/SCToS57x/aRWaBngSij52p92UHlV/TsZq77OZdYCESGd
L7pYmUAaR3DGsOlSnYGIR/R6MbtLYSTWEXRHLVR6hzdd0q6Rke+1Zfk7wqxSXwnJ
7127SRoNXNxRDu11V+pzFEg4OSv8ifpq6wxhBqXwwwfAE9HGY0NK1Pu7kyaTaLqr
7ZWSsHtNjtFjz9iD9qWFOKAlh2dRMBprgnw+nlnxZS99uBYJclpL/U9dpIvGTUTZ
j/DP+5kU3ta6V+v8qix2wGE74pntFbKbU0n575U/BpuVnXPtRXUEFTUGM/cMX3dJ
/dPZI9OKVlvWpKCcEaCSqcc/OPNdsK086WBqr4zJTRN4YM8/vfvfgKvpan2uR5Tj
onbgf4rNJdSd+mR+1wxuAPVZWbSS9TpQqK7g4r2Vm+il0iMfowe9LAToTh4xgXRA
A1cY/pOHtbArEaY1Npqb2o2039FTv8a1DfciFBXexxLMp414yxGlSgvF7YfdYMNM
tlkvL2RTz4jG8qELIOt/WoTGZIMHCfKC9L9I3GA5PQpaEdGdPoJJO1l5BQQkvcIh
e0GxgfyDNcg4awG+m4GzOWxqVYuc0RGlSWQLBqqyLR/++kVtEtb9NldjtyIzdm1M
QtBevYT90CWDeAr3tYFZ1qnarwSI3pHlKHsGCUiPvVP/NOmOmg3lo84HY/gO7N09
+3rwDzqlPvGa+TT1NZoJLHnZKjfgRu0myyJNxd4EWzVQJntYD+WrLBEtDHwltw3I
wXwpGb0l8nUzyf2pXthfZh/8TzI4BIDgzoG2V5LxqWB7MRFhyKNn6/BaZxW3MSoc
b68mAFhXppLPDKCaGJwXzCW4rIpIUVl9S8XW/Jjon6uB53SzMYD/ee5qIifUTG05
Xs1gZFn0TdEiS86KyO35lT9bhpSTs44vqGqFP3HtNrW06z9sf0qh9/zu83/mRQRL
YVZKtjbUhBbjRazZoHvIvRBxU82nAcVFVu79dSZWB85INp8Sri8oAGuBlJBnW8gV
HsQqGkKFupaI2JX8Rq+6Xwe9eyjw+relzWLDXvCehFYTHPvaAQfVfAsKRmfM5rff
Keq73r3Kxs1n369cZgUjNM0wkeid/bmcT0kM+OVfGJDZ6JK2cYePiWGRbZzXEgPQ
uf6ZWxRxajCeMtiEV07Roo0OQiePjPVYueXSkY39JiZdPPL1PSk5bMoA1T8ZGfC8
LqOlpthlz879+bUOyLtyNGHYRsYyqyYBZoFwT6ql+pWnM8FKC5TI4Zk82PMQ6ybH
9oMxAyFo6ajLCsldibaj2lDKdvPy//8GbLRe5WoAEPZCPvbdtnBxFZ4xg6uU7PxG
mtjYjKcxmGgthr0qXqYMom6KjfqD8ANttWH1F6bxnRdrhCteBbKh2DkWb7sZiayx
lDtBpAkhY0TTpiF4h1MBTPbyHxoTyh8idxXetiMjrF8aZqq8Aq4Kt4d5pKiKJqRJ
MSqEe8p1D8QdYHJkIX9Jinmzm6WPbk7pLCZ4Z66L3aQ3tvjBYBIv2WxFNSrmJVHP
GHFdu7tY96DJGt0O1MbO2uil3ua2FJlbuNl8UKRvvxq8K/7t3i49Jc0/cHCdVjQy
J53E387qS1SMBQGbJ7cAWM1gFkIemKlFbZHlu74C8jCD75ArVDBKk+nv3tIUrc0T
ju9QKBKOADgcMqOK3Pd7Ontz5QRDkd5il4ppNBIer/0B5Dia6MbCSmqp7AdmZC0w
4uOpD0TPVJG1Q1xJLYYLBt6qI9NsMmSH67k73sZziEFvvETZ4+YhAjYLdwAh3JvM
+ZEfpfSjwJUTk9ljrcG14HDXwrj0nsKk17oIpXlpNltlLGejG9o6hl4lzQaptG1z
Ctm+4oSz5OmqWuZLZPte+YxWyx4Cup0TqNR3JY8d1FuzRX9EHGMY4mX38pv/8gcX
SIh5AYel9DEP7e37XbXOje/0zD/a5O0nizB720ClWSUSYw4xDyij6eXkUjj2ECWT
65w3ZAWTJCjKVd7GymAUPahLMrwzluXDJnktXMkKV1SxXlUw7zEDseAOpZoNk4Gg
xC93w29l91qGivHPvqA7X1PUP6c/OxhQ3GlzohQszt5FAd7nZC0Ojvzbyy/YPJsV
9uNkr/1RiLTFnCKvbD6uRAHtWRZzwoBxMkSeyRiCTi3jycuhzpWK3EoZwKvaqGI2
mjYlaOL+vjJdOgDLaRvB0rAIamytI9D5mcDlEEZgIed4dmBS4muIXEzUeTLsvs78
SZZkcyx1R1EqUrk5EfQlvxBHUVoIIsNAaLw+bthYSFM3CboX8qAWbu+MqPtlbfOM
VniVa6j08Q5DOntYIHWmWVyLAesqE/1XOdPjP6CW8Cin+usbO0dC3hFaUYvBFGPu
ch2JCfxjPq4KZq+4Q9c5yqBKJ6A7IU5Xdzko4QQ0apnnvn0G3EH4S8rjU/fTTi6K
OCpIcTQq2Qod+uk1nKvIBOYCemdd0XJq5JMREEAz1ncU3CQ60nFZPqkvr95HMFLJ
W2rkEZV/2OtI628tm8Tpq5dy1YVlVj5zN5GpdgyyMvhFP/yx/7hl+5SepC9d/wuR
43hBeuOR/9vTAS7RUgOXpbwPEaUPwqpr2+jhCnYeFcFbDeSxcjmY7ENKyhIZLZFq
cvyznSxbo0OCP9mTHgYg8dvqiNWZXjhYauc1xuwQz3T2BLAc8QHjJ5bV+nKyJZma
WTfLBIak01QW+toFEywGij3CX0qktPPzF5Zu+DISKhHwc9shtemwlcieGtyI87/D
Yq7m7HchGJiSCYai+S53gOBtRpsspa/oJJiIwpkK64PfhM6jjZqsQXduCL/Vo5to
wYRzyOXd3CgqUNsH9uQNYZLjfognzY49BrWbzzYQLi8F3HrZRWYHOhCOKNqBo84h
G+dmaufqm2aFRbZgunygACLE5UEjOM0mu0psWZ0p+ytoyVPYjxE+9NMaBGx1RDt/
icMAmnpCKiaxHPxB8HRu2gm0cPOOPdTLB3NxUiju7NwCHrOTtIgBc7kds+K/rdZC
NlMAuRXXFzWmDAQVcry3n+a1h13fMoylulJ1OTaGbSbNU3NlUc6w4bmXy0ZN0nB1
uovCfe5UFdJCpfv8zwIgsR4YOznytuPr1SDa5MWryLkn3uDJQti/YE9LZxDXi4m6
2Q6it7lxKcGG1ERupO7nptMxQNMLOyS7rN50QInyX/Fu/zwtCOOs1K33kRDmYLym
EE07497bwwn/PFTdt1JbT8GEFvMZMa/0H0r0z1gETMRcOkJVGdUIo0T2lWz7DKmX
U7VydoRrNBmruPCbZGBhgEsZiIFmHSjJd73p/xgyLj/TWWB1drCt/ZhFJJKthbdk
J4gHt0F/9kdXa9LQfgyeLMHFDyXSYoceeEozz/EZh6Idv1FdY5Kt2t5ks4ipGCAy
wg7XHNXL1kNX8QBocgwyHt3BE8WXFMXexnfx/PxoSlL3kgAvI3aBMgDLfI+feMcI
YXEN9HBa7imOI3/E84BqIl+Wzaij4/DOwOsEPTnb5X61m6D2/J0tpgjxV9G1BkjV
uH7EGBa3iUl0uDZVbWdG3ESn8btaD+LKURaHb81lTTpBdnOae2fSSq3JQxkfxYAr
AayJFznqowIbqSPAUM0Y99TS4T70zkEvT+eZTno0blFFdtAs8TJavmsGsoWovwxV
RKz9S75J/ECHqaX5ZfQSALtGJwHuhiriZuAtNt5Ics+gNnLuJ1JaJHA63j09qu6r
YvFys3oh2oa/787lHFSPY/5+2jI4MaSScubmjXA5dffNIKqSj1kIcagBALoYEQlj
uOy0K1XBVAMZDv1NPBWvX9mtn/cvku9ZwGT29rXESFjfLnMuSywyvIC6f+w9Z7Vv
BwZMzaLuBUPV+CG4vyQsx31rI1XBjJ/1C9TyVxpI/ZLfZdou1+hr1Um0eg+clZZ+
2VnKF+5jspcFA6E+9TzUzpPhtM6seAwlW5fdEhNg+M6hcCXSpT+yjMYGglK7P2yx
s1P1YSnoxkOR3yi0om42PAk4D1jSYBV0B+aS9e5vKYm/LSKrFBTYwjAw/sSlCcd9
tEv+4HOdt1nLJXTzRTtOYfKtTC3PKiXHqGFT9u7VpklpimKSS6YLamv7TU0QyqGg
3THvwbG5eyVZGqdsMFolH0IJgYd1SuopcFpKq3qqIIJbFAWPlWJT9h8fORCBJxdT
wHLCg/s18YhUseQZIGfEy8zuZFHdt+Umbgi/mK9GsDq6wh9aXrvHjrz61nquzlvL
LnzxUKWOfUzbd16F8U4An7HFZsW/buPmTgIxtXPLJ8Xawmal0ir5lZ12BMQPDmG7
QK+YYjVNIoJKUxkEx9brqNvpj+oudVX6wiH2xznYvkNwFaf9BLJtPV0UR/S86MX7
XfNjmJNtbj3bDK8JmTsP2j7Ap6sIWL4nrTCFKx5kHF0ES1N24XlDsGSEEyJJmvxq
KsXlfi+IQw7EgcocQB0GQtIpO0CGkZ36KRywE0s2MBozfjbe4i+W9VgKxIMHULWl
hquSllrs+yRaAq1gKZ9rV0dKgRtn7CPY+pgn5enMtzDn8Yg1sQK7DgTVs5btYpom
aKYPt008gSjIQMNUe3zCoyc8b6IWj+6xCWoWKA+lb6u7ZiP21DXJjgoZTnZ/o+Lb
v9tYNjywLOZ4ZJ9hqM49R+IVFrlZ9VAlWELjup2/XIGl6MdBIEqRTSuOQ/6itPek
8gzpJ0MVBuvO1ksU5uSvcC86xwB9Oysh4AKX/LyDgtce7JEF5UYnT9HxdgXdd/Hd
ffobPMO0O08JZQkMUVc68DpzCV6dMz2bpypX49XMRVHeYutsaA+ZKklrCILnoq6t
MUgvZYQZIHAgPT38V+bIDQUY+ZVlDPuHLo1qNEVHVT+Sw6DKfyUz9BGWqM6sLeJ4
f/uUJ9UIlyLqyL3UvrRvdLvpMpFV1s1gGzaSZi9oGGZY4Wp1pwUuRmQ4D1Opx6jd
mPq1pt1rDkxA94Ia/Uor1HdQnrIOYCXGGEzl/0va9wmuf7BKo2ZZJAVxnMU5EQ9L
f+7XnceXa1BmIOo5vOGf7rtOBsrKy6U8k3JfUJtIb5+9WD9GnI8wHQzB//VVYtGC
RJBumWKyPHu2KnfaK/m3RkF1wHfxH3Yj47fwhHn8YCEu/33KyRAij7kOpf249YWL
irqUfm08Uzp6y3tUyMYg6RjKLj0r9ysTuFt+ySq3mF9FQO6sWH2CU1VvSdw8TwQB
i4bWfLYHAQE5AIy7VaTgS1lNURVAtqHRDNdophKFrw/Xgq/4TpJxuDRRHPmwGuIA
9XzD7vRmQJnG1yP65RmKGgZzUpM3I0EGoIt5zLUXnZQgj+X8eKmizsZyDrPjiEW9
kvo5Z5He7zTDgjq8tvoRG48kf6GaIjm+kB0/EgJqzhb9mxe3ChLPTH0Ab2GVkr6B
ue5lnAqxlzc9i4dzHV1A/oEbD9RO5/tBsj79ImHSPq2b0/G7OekJnQD96hSVljbm
h+nqtg5QipOjoKKcemEEAdkBauwdYdbhlIH6hnHFgJFDeq0XUTr9oJaxHKI8gllP
MoieZNgqM2Dm5pkXW1clxHymKKFB1qW+DUIZGHJDdLa2lBFOrCbt6pEQH1cdTPb0
aHCMDw9QP+opUUDi3gjSzMjoG6NIZo0hyH74ymsPmp+MSQnCiuml4r2c+v1dBdIB
N6/OLK+KpFsNDBjdLSPtH6bWg98f2X4S86wfpJxbwJArpp1HGdV+Bn8bm24xR7ei
+8PTdlm3pMB0Ok5hWcWeCltWEE32fySsZHR2FAFO4gbzbt5mFrisWtubNmhWc2MU
4EtLmaW+8iTJzdTHFqzd3FQgx5A5nwsp6QN6NmCFea6s48e5zOJACOkRCNmuPscB
qaXy2UCjv3euMYWIwnr5byDzMES2jH0/s/zOxt7UEFUni3hxqB7GoeEAC9zy7vp5
bA5HhpgvstY9WFhNewDZA13DXwmCGOareWP5ptpAN2lB4N6xF0wjkWfP52YpiGNl
1m7gP8h+vHzXyl9h6PewWf546ZCZxBBb/oUUWJ0JHSNFmtUIX4JPPOXV8ukwQc0x
gB1s5kv3lSor0Z41Wqw4rSqqB+eecMhuMHpF2lepj3R2RcuogEQ/n1sjShoKthti
TyH96EI0CAi/1CDL9weYMlvvzuwmxQKBsc+IE2oq3zLT8HY8OhpzwDWCyFx06akh
0yPtLtCA4+L2nVREGTTCJbZbvgQnAYX4nlYl6wSVAbW6QaltuApu74hhEU3MADDL
dQ36/pG0BtV80vNuaQHNPNT9nBoNjY2+KICglBp6HhEoS/IjIYGa29bafQg8IXGe
LVdu2VmjI2l+6J6Ql29iw1FAMq33w4nKyFadCKFpgD3qbRwjyfiAnjBJzlz0OoFf
EP4KKcSrtZvq9Jj1svjRcyeVqHVo9AOZ3/sx9JolMelrlDzpE66AahGGb32GI0SQ
zjfeoA3xiuicGoAa4KLXJld4ZKYhhdoeIXqktdE4qEzP0JhpjMKXFJkBV7rD+xnI
v9H9p38iycj15umNkJQm/i4qoU0FGGDMgOoR2Da2lBVJGVq/xMWKzqhJy/6qAD5V
Dozd5LbsCyeqWsjSK9NC+ODjFFnVY3qxKSAL/UsvimCmd8MFBvwtI3bF1Yl60uH7
Z/3jodb0VTkxJxdy4g+aG6gLl701Gw3wS5uTTIs3YEb6f/+rxIkrRgfjzCKzk5dG
4kqOjmYGLvK/Vl4U0FtSX+8BDEUb7041IInzlYTuVxVOSsWqaBBOFmYx3Xxjp+3D
46obEh+WWCM1MXtav+bLReBgY71OQ/JYM026BLGzXVu8bnhhUTEEbkRZidBNYrR7
pF6kSQpNIAOkwp/J9U2bT3Z5ewIu8uOdtemuQwDQROwt/tQgvnAQ70BonpyZSzWu
Z9SIkbAZYMnTbOmP3HoTudrY9UrTd6COoeC+a9iyTKUGb/g+RlIePQItZ58zJQ3K
1PX/8ezpXNh7ZPZ+GHr5LXLWVTS1acOfpTycKfTjU2JmANGVS9rd5ncNcF7Z1toa
7hmLSpmNXvMynp08Kc3XSZ1w3+H/UkorbCzw0S1WS5B7LMiLOC3ekzlCM3lwgoTi
4+iASmdLkFtAJH5mTFwsq3rPmH0JMStO3WBJzp/V7YIcA4N1N/3ozllB91vrDd8W
N+T0Y9dkErxjG1t7igqnb+9bPMozSS/XR848CQdCNd6ac9SXh5DBwrW6X/BvHNvM
JrRseItPgz5SX573ki0gi1grUo05SJASy4t2vYCamjMhW9l4GihJv5OpW5D+od2/
wyg5LEcx9mUnqDIeez+EdeiJWmfYE46K6uYgnZbO9h5tLJsM7miESZdj6m2t+gZw
jZPkCe5m0aHol72UjhTU6mBpAQgy2G6B3k9ul0dgf06/NY5pERjElf1XJ5pq6Bp+
I3iAr1I2DtnugZQ0oqqodtkDEGLXWiBzkdPTEK0Aj2481C89gAO5jqi1+OKbyW+X
HETOmPeCV50hJUiUCPb6SQYbkZpJZQ3Kvf8GMOs6sjZiEr1Q/01e/9AcO22jxE/c
0cGZrIs6iFbh9WAJeErY5QL4mZNJKyJ4YkPvzvvnTs/tBUw1Yp08kUNF0decHuYL
N0Rcv4q4HCShjxd8HnzQ7CBpx81id4S6RNMMD8iltJ9qfTVrthPXq8be63v38XIK
CZTkmJrrmVj5Jm0lyfxnDq20biJPq1oOhgIP7aJR++lew6gSWMq8sBkX7q1znqLV
4zJk2MjIAzPkNasZpRhNWHHrMKmAInurJsJUFFcHnGwEJHlS4t0F9G4EzDmkQOWs
yoAYCRgtSDC0rtHY0Jb3qJafEVkFSAE7vN2RBVqDiKIMPoyFJ7b0tSbp3sS/eWY3
mOFKGEpdOgQnwyq5GZj8QrAZnViVUN4YEdOjwLAEj/ZykVbtvxiCWodWgFWGRwNH
Bn7oRtgLHFJsfs2XkxenbyQW+tJ/uge5j3leepLeNTuDB+ZCDKz6BwkI8NqAr1FX
tYmuMF2jcU4Db2OxeZ6Cf1+hF0KxQawmWtzJ92Mkgkq8Eo1U2n/6ghPRL+D+S2d1
8FF6PP6y4DmCKYamaQCsZ9WQmoXbTOXUl9FxkyHB0C3PrW8h8U2582x+/2ihQLb/
skeXy+k7NtXOTuN3vr4E7TFNWhs0Cq9biI/else4znRZmS0HlPOhm3rpOtKugbkK
MnLYW0XGOdzN3c/XQ8muMQbOXVRnjyT8dtKgIxnAo/XZECSFd9O1eWNADjKl8cGA
ZBRfc7d4V0RBzZvGx4tZVHMgDJzxGMP6srUHcn5zmHC3uEr+yp/osoeqYWyREHdZ
B/3tuvIqzKj2dtIN5QHFLJugnNquxBeBUdNE94FYNTITzFEDGZBBVNFsTgJ3Xc0n
FYMUUcEFiQ/XsnqibHy98NgjfBVmELX8OH1uZaAPbHnDs1KW0yXLpJ/qiiP3cUwX
tG+Lm5WxLyo4OvYshiG/tV/7DmsY/nU3qpderSrtuFBEirz9i0IASz3LBDnhO6Lo
+vuBz9ilhVLDlEhN4ahDRigPfolSGYkPXjTiN42Y2OL5IGpdOTLKfw79l8j8vP2X
efq2dFzm40/S3P3vN4DzSLbldaIpZMDcpdlMUYsx5DRLxEHV4yfT/YkGCNPGHTmY
5PIjN/qmpwTN0EQY+p3ZsMOv1TS8AqFxJ/42gRKguESLRo3ZAkMvu/D9+G4k4VWA
InwfJgd6i2d0BykRqpjCB6CheGvonmcOxM/uige6J+lAQv5ThlCGlck4LtzcbWvy
4dofgVCU+NAcUlfrMeyZ5RLPKuaLgic1v+WVL4ECaIhcMtZwULkV9OSoxAi3I3Q4
sJQBHwha1I5bQPl6C+Sa+DQLnmGJTjw9Ih3Mr+hqP9Qn6EpDMmwipxY84JSLWiSY
PBSF/mWEy9uKvuN7zpug6cg7ZLYTv3vHQU9+nuABpzedOsZvOZTsPve3JRRlh8VQ
/dHtcBUOSzbgHjO6p/HjGFfzyw5GEJL2751svmj16t74NUiWDw/lE8wr0/7TRLAu
A9NBDnHJfAyjmATSzXweaQjiaOGCqg8BsvTET4Sf/BhmR9Ox8TM+UiYGQuW/u1iz
gINR6lenvLwrXGk6Ckwa25Ebw8rw/txLH5kizTZBk0bQeXM1dZ4cpg8yi+vGzBIp
D4nrtpDbXhkysAbEQrzREGupfOeuBHP6rYekK0UXI9gzxhd+NFbBM4kWmC4/6gm7
suEvIF0CcnO1uwXLPnCchw7gjJKA0N7hPZlB0VZhULE2i2cAjBSUhNzJe4SklcbH
c0O3Onku/SoyIaiv8w28aL3zEweZ2tH/43YZOUpg4i/UCOF7g5j4HhXByKjqEsN1
pKMvQnwFFaWakxFqqkQois2EJHBYahGo+ZWOwcxtJa72c1cvjXCslQK1PFsGqxFC
Wh//OR7AAY/M8AfcBkEqwmnf+vqKzDo82knq4FLxiWAaqET+QjLhxfWtPh0VubFZ
UdSrrdpXE0D9XmKrOL0jFDN8vI+uAwH5/QXmxCXDWm2kXxIPxU+61QbtaIPq2T32
x+Jjxmu00QblmJjtqtmmcjtx3CjNh9jeneoqaSE1WRhjAawaVFil9NcCL86gF+y6
IqRdD6wva5nU0p25gv5c/LRIrqgkRY3g0kBQZRcx7obyWn1Unw9ytYmbLGRoT7Yp
hDImsk2Zj/4hgmuD0FfU89Vvla9Dku8YtEYxNBIkjU9C09doCdD+HDaY5mTrYhAy
e1TPVQ/KefpFdSk1A0t9+834dtb9GcQl0Z67rEgICmcIyQLqhtBFDFbywFLlB0N4
U57pXkZWPhMlB4rcF75h40rMS5ZPGXDwcchNiGD5ERSQZsVYh0RQJTu8o3wQue6S
Z4ZgcIWTa9WUl+7my5e6P0cEIZdn9cjYOkddH3o57AfJ7Jv0yISEo1vO3S/E2Emp
hX4/pSAyBmR4wYLM9xAbCHVRK511CoKo2gG6pO0OtO/xF7Pvh1lc5c3I6Obc9knO
iIry/a0gc4OBCPcbKiyzLnjoTRybGHScsDqIX6WtcwtiybHcnawov8fkiSU52Zvn
jUkYRoej92gML9j/dtPlsYDXVvliHdT6e/JYZgLSBw3jJZ8d5x7UBB48vRLvpPo5
aLYQ+qz1FkZKeQ8Z2oD00sd6UyrYzKye2ILHUNIVAicUnU75g+IkcTkoZx5IyQmV
hVBhc40ioK4ncNBReIwKDHy2LhF1IxDSOFF9alfKq4gBw3sEssICR/m9B9YUwT2h
THJjn7OETiGu8h7L1zN4gKniCDB69uaBa92uwaVUt31x01Y7Z+prLsr4R1mts+bF
xorBgKWmi/rGDUBn3LG277lCZ86zdviDWvdyBqzDQZ3ugDIuTXsB/qJL0lN6MoW6
9of3kNSsZPhc+nLUcii022cqZ9lWLDqfu8E2zOnAyHAdFS9npGCoT1bci7AKeMRJ
O4tIVILKxXGMurFroEB4KaFYNFyZq79fY43TbiGvhulcCfqNqcb0icCLYhQ/aZ6/
ROCTO0i/W/n5Z6ITomCSnoe8vERYH3ldb46drffVd+iFEjnJQqL0uv3JqMNbDzWh
blSDSF6DO8Gy5S2HHgoJi5qeHrUdjKlRU2aC+ATgdA9YrvNSZAe3JmBmoMigrDRR
VkXd/GrspGhjEsLyhmNl9smAUtLLZwqri+smPZ9VAQ46FF/t9F0f8PxIr9ZcrrEO
+YuMER/R7sIBQjlXrqUhQ7V9PvWX6gg7h0nQvwGj/ZWvOJ47y7nrtSt3ZAtA1Un2
Wz1qCoITI5svGMmxvzbUljKI7TBvQxkMpn0dRFgIH10PpYJ49PLp6kpRzTlNdqYJ
i8769KouEfCR5XpMgRZRbc+NlsaGGUo5npaDJhN9hCgp2K4bxQHmgmiocA+5x/jZ
YNzme1b4SnabSbTzIR1RDhatZRRc9tS0VJjULw3lj8AAI9URJM5HZOjdzv7p+txk
ekjpm1wThO2blPpa0ncjrO93A41DvZMawZFifpFMcwlmRAQWrGDZLWm1qmjJjaXJ
RcEIOiHbvtELNvFhH0iNzu6QtISL52OG+WwIJPWyx5IiJkjZzKadsgWGDmGQlLcH
Q4bMRoagbHUP/Wo12qJGnnsN/8kEngDPxQJUh7/sA5UB1ZDR4R7Pte1JRd41ioMa
TfbhBNRvjWWK0S9pLlVB8WgEiE+QBThjjC9nEUT9ERqqM0u/GFhlpEBsQg1um4gu
S5TVOXjHYcbCNVP4Hb96uI4P7sba7DU0dXfggqLn3XjvcjvcmnuHl7EXHSa1muN6
Sh/zBjwqoei5aeFfL3G9O2KjLOl+xv63TCSLa7o5uhCfRKaAgHFJ1iwhn94i5hi+
W+afav/FGrz0P1jeHPkopkPJPHUtyIc2XNTXIXXM8yg7Eis91cFqDIK4mhg2TEA1
GyLXa/xMtbNgn1OYFzForx1xvVecIjcOZQ9IqiP6kKdgskdEdYhZWJNdwhPiV079
whKbTG6My3i3bpnrAEnHY3C6pzqGkTPhp551df3MO+TChYETEva/V3sRSMLQ2o79
b/iR4ZVQ6YEbOYmxumF8KjMS4qDEjztx1zLasgWv/RtschKtNuVukgQY8+X0N3iy
1adJYK8vFlPGHogTwn1CdSBT5+W3zW+Hivrf18Nh+Omy9mOU/TR8vxj/KMsSQssl
2JK+xZqupNIH6e/pPQjYwH80qqQg70WF5arl4NkOkm7rVRiiHr7jG2KSaBWYdovi
mIXEkXvnRU1KmGSefOY6GF5SWqTaD5HWeuF1/8jo3L2vMwfxWy7HQfBOSri/HZgS
QaxRbRAWnKv+yoZMpX+0wYfiM4aQrvawsoVWXvfsE+OA//n2v6rWhnHfNuop6ByF
z7A+Gij+MlApnr7DusSQHTZEM1hvM3RfDNy/UZRgSaZXt+RO783NnzPhAPlpwajg
MQHyrH/dbjDcVySS2U/hb+LZBN4owBB0o7hZng5KoamnJ8MSJiTW4ODfOqIN3E4C
mgWa4lCHKLHpdWY8H91skeQp/nLyOqF+l0w5Vg2Ki9yR/M+BGDQcdQI4PgL9Bzzx
O8kr9QMWIX8pdIAtgQiwvLLPN7HHpfsc8jfhouBaieK5cjDL57GD4nsYOH3OdcUa
XuWIsldkEh2utJ4HBl8dmTL3fU2VOvmiyJwpZHTHJS0lj1qagtoFtTZiBoFDGCGE
qiYAEDckK73jAusqmdNIKy0z/Bi3sYMf9r6l7KQWUG4xiNpepfk9GPlxyv6F8Zd+
IIRIexsjt9WvfjpIisbbhC99TP2E80lR3E+K2hMCu5CUaXhL0lHiPdTGnUuANo+w
7qZa/rBsclRgP8WDuV9Arx4x85j+OT7V3l9eIHVBZfowxTGWP8qvw+XbZ63NlJT2
lSbdFcyPY5QObJN9OGqVZ2Oe4osc5+BloL2kXU3sJr+cOrgj8HGFB1ngppYSx2Qm
drJfcWxjazMyxYdnPVaNh77W7GqKxPYEq6faGCKninnZEQQzfEVnoFnKWHyYr2CB
abfuOfolMxVx1kIa5T6oTyNl79QvbeVLeTHpGwqrDQctoebKHoDoHH0dqTD4ES52
6I5V/rTWXCFE3S4JMosMZ6W+GHduUgTVJxQ2poT7e9IksemEwP+E6DFGZ9WS/fbw
oN+7tbpd0rr7sVpUmJdak1M+VI1y7mHSLO7FPMn4L4ZEVQXmwgf/0nFiLZQMlUdY
J4hJYxGgTLroKXIuKi1hPRESIGG5AdeM5lSq8f3NQpR2+31PiFocqI+PQrBDMU3y
GNZSbgynh+hjECgEi8F/xFEVhYak6hCp4pusOdVEr+4NcHd2VL2h+Hmhuie/hKZb
MqC0OUnAslxgJeeixnwFJfnR4wx+oQlmR2jHEk5q2PPJCLlf/sPGKK7pX+zlf7a3
UJ5JA5hUscGrsy1WLlM67GhVvoLedtMDtS/y8rnQ4vkyhGahcSPAnBEDAKdaz04i
PpOqAjaiRlFnORgS4EfysyiANC0crEr/W+KM/53plysQSqpIyMaZIXcPPK6M4Yub
E04hyhUTHQRwXWoxzgREMAZZ/5kL21jc0ES8DCoWShySX/NDYziFYs2ZO/Dpk9O/
/tIhLpDOieAtlCot6YcISXCJWGFrlhUJtNw/dGUwYFGwcDYnWLDWqc9zgp27cloe
lT1j3v8Njz1Miq4C56XtEZCrM6hlHe9JtJOkKdSqN7eNx0DqjbacH8f9lzraTL9h
GLy5a61EGtR19QBrfbYlEcANqBcRmig+feev7jt1QzgN58ELrYJ+z/cAJYX0dZ7P
/PGcjdAouhOLuLYyouUPlC+JX29d4HliiycfeHoM3t31m7l+RIc7R0p0MY9lLSa8
DaTgulYEdpdJ0raxtXTGLMT0gznddCWb9v7EXgpq5nOaOmSeDzRUb//JKB4RpjkA
M5WgoOJBraivJ1QA3huzNI3XHl3P/s8PHxgDX55rVB/xC8RWq1hrIRGDuq+uYZKn
xe5Xu5fo+eK+ipqRPNa4im8GC/LOudxkYNOPXVZxP5cotEAfUc81cnL1208ucHlM
7wX9m1kSCHjpPkPa4wJwlj01P+81aOVOq7l3jNPFJXacxraYi3C40c/ugGCyMsWB
UAc7MTpcLWz86v7igmlS25AhmVO1+3PkRAkhScLoZNaMEZwmo8vLkZ4DB4N61Ejl
8mVl1cvzNg+9HeFpx7ijaKWjeGJtYbH1uS02o6D90TIHfwUcUXHH7lPc8449PjiB
NM/X6oj3q2gd8ezOkHvSabRdtLY56nCj6MitHffevl2fiS4+/7OqDW+INi+F/0e4
62aXdShnUefrKCW7mmwt/Yq10fkAJKC66qxqHj+ssBk9m0eWqGYLTMYcNsBwP1XK
HA3Zfgn+BeeEOd5VOX+IXwsexbzj54n9Hn2SHrzAkKqvgYVkD157LEG8fGQYhfdj
tebD/hF14Rt4PnJsVIZsAObbsN8pNzsfF9btteqfKVrMMDOiCn66TwK5QhfrQUQ3
ymvdUp1ONY6FykoPv1X7eu5Lwr0cRPKiMemTKiJBwnMJa2gfCAD4N2r8rTD6DKtb
wntFTL8BvEaCkSfHgpkQox/KMXlxyJK9p17Q6bAvZ2Y=
`protect END_PROTECTED
