`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
0rHGBieYHd3nMrURlLU2kh1TrujcOxOk6AxeTYnBREIPsMls+UoKIFm9g61dN/BH
QyQaFv6jkkfzF+yY5zEJxZaRDkXiXD3NgN+GfYXbKWNnnG2rzI9A1oV88yncI+eS
yKqWWXy5D7nE2A3ln+Mz5hlbEhbUwPmiPvPyuE0RMtny7r3tA0tpQ2jAQkvwCKPt
itPbtTrvZJjDannQHh1MnevgXwyZK0Gugfjo6gi54X77mlKGDN+XfN7Me3oMDdiU
nkwfPmJCPuJTr0+zctlcg3TGQIIHz1jm1IK+ANKeykquRG+fKL3tQu7f+AGrnTEc
3dWe8SfLL8XKNov/VB/cmaxBFZ6jmzf3InMRXrlDz9o=
`protect END_PROTECTED
