`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveE499SEpJkrowE5HWbhJUrw+kbrQAC3tgBsIIwoB2LFA
jgU3ewiMBpm4m1Lpz33N/bMarrxAKaIsWAebgPG+Wtm1UV3z9UrGqhFOuxXC+5Vw
zmAGRWkAKfOIxDK6Eohdo8G0ypO9m3m5VVEo0GVjtW7haoxcKwEAQoHW+RoMF9br
KLzuEAAh8G+PNjXL0ocODn4RmTMizMPwXTN5CG1BYy7G8mSZXIJ570i9tsOLeNjB
RN6AZeifSE7Y0fA8hw2c3Rs8KIuak9pI1FBoYoa6z61WVUKpf53zJ70FQJ6Jmqni
dslQWkH7u3Q88bI+DvsgzyYD1gDEHrScYlWRVMK7LKkOYxvj4SVKnETN8P+S+JGb
oZWViPtOvVDAAoHYmZaLl5zw8oiwq8pC++OfkCLIO8upBpwrIpGUKPUMB3NwIzsy
aowXxmA68+C+7nlu8MugFWBXe+v6LAheiaJjolXt6lPNX9kyLbMWPO1txCpKytPi
OmSTQgA0aIVwgDYk/DeDwcevcDVj0McRjok921+m7Z5Zbfbv2kpIGNZLKaJEAcUb
1rzSavx32IUiHCwwClMQZ+NTQ8SecGNH7Jts8fVH45x2g/oSg4GIiTpzZJHZ359T
o7/pm1Ko8K3SJfpn61ehIFOZ07AEpLaquYyZUhSvxQfa0qpPmlL0ZSJ81G0DF4lk
`protect END_PROTECTED
