`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN3ycBa+j+9kMUhkN+7216kWPFkrbRgVFyGdxEttVPvPB
Ag3ad9EqnGTbmPc4muKWJ4hkFMN54cMNAq0MMlI7V5TgvqiRvOD0f5jqpgVccJx3
u3kWyZLcFeh7JX8ba15WNkF2U1zCHKb81Pa1bcdXx925baNAFIXK/jEqRYLoIpGJ
J5meKhfWJ6ITcV5PKLRAC2LzNnkj6/uoirXInHLpGUaQMk0HUZFoSz5FuIGsOQu4
MwiFjeKHvI4xAeo2BBLQCGOkZZjNdilpFHLW82ldt2pqmUv/fAkwJ4tjbAzX9gj3
htU3eIOfbt/B6scwFKS0TVaUs83Yw/4XDym2THQUGW7oh/vKWT8CsoCKe9FfiFus
2+/tADXf6tVi4dEu9hADKqD/ISMCVw8NMxN8PMWZC6KKPF7Wtzhp1rFsGt422la7
AMorUd1zFXBb2pjKut7ZUn9dz6AhPNvTvIJQin5jvjh3NtvKDDn2gf7+lJ3nmL/A
TGHlvilMcYJ+b5RXt/RrX4kLDaDfomOlyDWj5vsxmjodoHs7VXclLdgtb8UvSF2s
rjLEN7ypgOz7Pk3dA3HY5jbaOvKeYuYU3ZqhH4wZGBHdWfLeX9K3Bsr+TGON/USQ
g6yVu8Gcqp6N7xFD37Ijxw0aoQuuRP+M92mzJ9i3dd3h3nqu4WaLgao4I0V341kF
nf7WW129s00MArJp6JxEaA==
`protect END_PROTECTED
