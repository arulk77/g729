`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveADRdaOqBi85Kj587hPi+R7bbKpfPuvkt23m755sAsP9
ISO/BbclK5IsCY/DvHkaq/HGrsTCCpxQlZVJFhir3VCUN5UVB4mpvzVXfAWNRLux
OradKsM+g8t+Y2p+2r92wwUBgM/gQX1KMJRplPyzLoQ912uP0J1cj8Updg2XG9sG
7dcXayKUd9mO7gE1YsvzMA==
`protect END_PROTECTED
