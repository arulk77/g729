`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
SsAV4zHs9POVJQ5z5KMVWV5UP8K17gLiyI9CpQSWK0v6Ip4RKTiAhm4e+ZljE4dX
5bogFvii+ExuVa6JyikYM3YK4XgQmb6mS6Y6whv3N+Sj0PwXicCZCprLsLAxV3Po
OIo1il9EfUgr4jZpTM9LMDM4OXC6+6lpAvodbY1H59gScfq5+LbsSYkd3lwx+S9c
8KxnVJixvLWRE0mOxJYLrt9UgoqKQ1CciQ/bOPX8NCHx4qCs/eJzsfvwjws1gVL0
2RLr0Dhmvz3by+/L5BN7zOBBm0hyl5rdhwhjeVB884/WBtJ/ap+Wd+G3gWOntrht
LFaW3BgVzNRrdTf5t26E0AIvtRYRTX6VmNCUvZdkL8A=
`protect END_PROTECTED
