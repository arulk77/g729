`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
14+zjowRucobHTvwdQnAlhKZ5a2Wi0zXFdbLv7+LZpt8cx35LJYuHUYAfEHIf7CB
lHhEaGXmkudSlGSLjuV7NTG3jc/D0BHcIPrztQXgdLHORc8LsLky0R8UiAEOJNWk
8KNgNl0GZrsSV3K0kp8ejh65fZ8W9r0Tle5ADKdzdt1z0hwi1zhx7Gek6bzD52bT
ikc4NxSvPgmiSO9kc4HVOm/xR/GVRJeKfhoLHB4DY7GNLOJZ9UKzaSzFC5x4vy8G
QfXHfJpO62tMlcmj+4WOshu9t6SFEIy2lxdFsu3hsWA7uyJHNHuywsj58DsHIhsH
v/4Xp9Vf9yJxggm18K1gvZ3ROzgtNXE1WFxq8Si8YABLtx+hk8nmG8dH8XQIUZyq
Gpue0SwBLVsnNjE+CF/e+DKC3F5CAgb60oa/Ocl1DswMzl3bMdoU/vEXlt2gEyhf
7OmykHg3mZnfWdl4JQO+TPZC/hFccVCTNfgwWthGHtahyqPUr2LNID83gCLtSilG
oDxBsltGm6pggbL5iShhjrmWB0uIVuhBEGamOrDz9uGZIS3W/FBQtnu0GtQjmaQx
cP05JvpZvcKb4RzBZPcA1rQT4vAIH0tfQsjC2bne71Ge+QVRrAszjv+XD0kNMQVK
0SToYe6ukcf438XYuTmnbvzQQmRfgFx1V22WIAeEWe8OxJ1qN3EJ6DX8XraC4heh
NnXR08p7+a46y3OGzxKzZNuanzoQSX9+pFfJ4tChTmlRKXwm8ojLtwFlZ2cyPw+G
zGPAFSsyydB+HqPn9ho+Gs6xv0jv9IviQGl4/H8dJ0aF5I9hjBAiWlEW2gpzcDn2
Qg0E0A6h8GWPOhcbMcr4WfIvBDKtqA0bSBwrrbG6KY3GSMykqNydlvuBzaCJbNT8
OdYhwtMr5J7Vnf6AmPlR+ZR+3QeaeuB21w5nMIxytpplJzsgUeefmiHCgDrfP7Wv
kudkwW25VbsHwOwqK3Eos/BTglD1tErMHZroZvA8WkJks5TNXoRyH9eix/D3yOfX
1hbrP7AOoE6NEW1x4TMXdqCi2hiVbk/OIjcG8UDkAQHV9B43UDuAqRpGB+vvv68R
rWOaOuWkBNLu+3gT6OHzDeXk2f97JGj1Q/zbe+No0gNBnt0PY5VDcf4txKxhlm8w
d+6r0fYvsm+NXZ5IT8e2k3ltk3lNqIMkvSQTi/9eAYebaWEwJUO3nEWQOAjg83jJ
sIWVLSVA5Dg18s/yGXTpARvPXMPEIyNBNKkgUZgrkLpR4wpjfZkBCzwqF5HeehSy
yAh6ekwkf3BKx09x9PbQXz1ovb9rkbSOymcfnxPDttcY/1k3X+3H02t5LUp51Tw9
zQCO+CzLVZtz6Ku/5siZjQ==
`protect END_PROTECTED
