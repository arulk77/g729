`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHPcqsPJXsHNlho7ZSPCkoeb4cGA/6jdunYhqXmfhcbP
U59g3kchpF6GSkP729oB4tVkZ5M/Z5DWkHDUrqBY69rp8JGwfiLKM8jS1GSrWgso
l+xUofxuRROeSJDKAICBqgCr2o54NKpo816BxW3o4mcBORrJtrpqC4MToo283IQF
2MGjpLXzJtGWhx0Z/8c9o3tqLFjVhkr7nq41oMhG4p6m6QL9J7OjaE1+5hXJczuJ
hPqNndc8wCNLyAIDHGxTbcJ92+cZwqXRz0nC1DHIuM2HiUbGS0UdErIfP3Yudezs
bkSrU6xcADGWWeeRTEQcXLOj6D/O6qNKJ/jDqAYWC5pcaUUdwpAjiGiWwMkViaSK
lQxZnKbwYF98K0WwoUUMcdl1WFxOVFi24QnRb6H8a+zuDMaZ8DCGIfA2Z71ug6aX
SZg5KazBT5DXR5ZGnSTUONKMu89hXRqtkMrElqUxuNuYTeSM3oB6onmUNnckcj/N
2P7V2VBXl73fpv8I1P/clDsMD/1n5KHN/6wkcMfmLfaTsQPGx0NuSuFDr/SBJNht
`protect END_PROTECTED
