`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL+f+diE2wVi5K6UQu2HFnvRPqdId66ccnmbjLGFNpiH
6+4rgtxRGTDpQgJYsBlVAYbaHUXQn28if716+rehsJ4yVbrcXxaMHK5MBT6bqoDq
zkXv0CK3owSFHNtYZoM2NgwCyvSApJ7ruR2quN69dgYbGR6oz0om+VAvUiE/woBc
5VWefaeDoCSc7AJM6xVYVtBfS+weYf9vPKNZkxd+mBv0kL1P2t20J9dr0E+SiMUq
65wZv4AhY0P69kqW555wxTi4kQuQ3PCPOJE7pKqxd82LkJoYHXgqndIshmX3vYz5
H+VnAS2nhKIMm8bpj/OWUySSbu160/aE/coiQdxO6Xn5AS4oZCPShzhghL7j7/0n
MMT7m3uoqq+F1BIGpoSdeHR+ekidDb5Y3ZZpJdPnyI7Vsm2uZ/PWJUihgJxfh/v4
zV48oq+A1FuClPg9L1ZmxOA1hHcJjX89xmTQzWFUceFV17j0BcYXv0XWWH5bGQsk
`protect END_PROTECTED
