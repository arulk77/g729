`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43bepv8pHsjfUbZVnelyTZTEpXnd4GRiMgnzvTJTTZnU
LguT48Zdb/aHBqdlKh8m4EY8KbB7ZxozClWG4HzDzYR2UwPL3G9bCJxK8ST1LiWJ
Roz8CtVe1/FZaXaag+yBRYgho0C8wSfjmwoA+Xcx/AyduiMr0xTplmv1ZHPDL/3o
rKCqoiTUfysYxcWtaAxofZxL6dZiTX+0VUrBZFXUg/vHmL6SXF1JA3npuWlKPPkk
xIkn7ziVQLIrG69AhHWSrcVQV64c2B2kX35UhFXOLUW+L2v1PAxAObJB/FuNzAOi
XMwQcGefAYdMtF2KAqpcqg==
`protect END_PROTECTED
