`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46/lWG/c9006e3J2iktezUEM/Px78qmuERuUGp8M6bo0
eYQUvIoxx3H8c2r0/kvCsYNT4QW9ranK9gbbdzaRWA9acT3TngBYhgfUCcPd5tKh
0bmDvqSKJozYtqAakUExMc2DZMQ5HyrQfsZVDnTkLzMJDzL/7NVPaGycJiXU8Y5I
003kSTFbLR5xui8UeeFiJyjlgZXf0jcnBGZcBHQNRlbK8Qua+u8tSTAyrND+1vq7
RaL2p5kAxhnTq/hKk4tugMuB7uMRLFIqqbPKMiUvLxxC5QXg7+26uXHzptrLK3Pw
rVaAzWQv1U5WqjlJLoDJYg==
`protect END_PROTECTED
