`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu490ZOiLdQcKDT1QPoAe3GOyvmeF+4pvzdJ1rjUWsPK7b
uR6DgZ9chJx4SLC1gpEy/PHeNgmCdK8CKfa+t4LMLS1OrhRNv1FzbQ9iyAkeeo3M
0h7zLwvH31ddQpQkS3K9BVUTsHt4HyH7L9ZEfGqtL80uN15nGSp/B/XB04R0eyib
INAsNcBd7eP5jFUzFQTk1P+mI/rbtsZSZCE6qlOD6mcshi4snRwORjYr+qaNmXdX
Nh5+hXbHr2RSpJzKdnJDmGK6CzvcHh3F/J2DuZyQDjI9WK/yr74qC1LVm4sHtmoW
5ZhFCts4yLJPYpKsI9D6QKmLE8qWNom4pyM8pd5C/S/ncaC3S3h/4B2uuL7MDYxH
znCGaQHyEVfLJ9qYxfmTJw==
`protect END_PROTECTED
