`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHxWzRby1FqejyESYxcsCHgdfJDypfLfU+AhKt1UM9/H
Ngd6t6T6ltH22NPAvOR18k02XjhQf/nMG9hJ6Z7WbCB7N8kd1k+sRSYHpqDN0C8M
Qzvu3Ws1E9Hw4ohTlpTz9X+lVSuTQDHPbQbAtpF/39CqfSBLw7IahRN2Z4QdYtkz
max9zFO5/GcpQ71jkmXKaA==
`protect END_PROTECTED
