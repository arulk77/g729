`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNYTw9juRwZkCsXWMZcxRDu+/zW+6pVykY5TbH7DhgPP
mVd1OyJUqe6LgHMqNCHOec9kd9D1ml8vR7ggaDngMcsUvD4pJ89eG71Xuvq6wHhk
fc9Hx/IYtrgReiUC6DBvjs+Bm2uKw2VDKQ7Ot2lOkmhq0lyTTXYtHKzCZT8NqY1m
HIrh93DyD1OZe/2kXBxZilRZHpmT0Ks5env+Vi2akmpDo7vZDF+eLdWt70xnCuEx
`protect END_PROTECTED
