`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47Th9zisSo0wp0TAjT9C8CoHryEF1VULsQVuNJxFDpbu
5ja7lg6Zz5Iy9gCeelSpKlGFcLR3YQlZtQRCFM6b4hT/qdCSzgCdoiJgo2hjMohZ
vaGrw6/g8KGXM6S3V56myZo9V6+Lcd8sCvOJaIpN4C0igEVKIYCdGKBTnJCYqvGJ
YG2URIWYPTbiny2d9n0rQZxL3MW0Wj/V+9Y6eABBY+HzhNO+15EAWBhERIhHDSA+
8yj0vogrbIlLFd1mRxb7AlSXiuLhKTA0WN7DIp60EFu1RBJy4pNFW9nxyV7dSdms
ToQtzJYsM+uzPtUVMoKr1g==
`protect END_PROTECTED
