`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1abYeARBk82/yeNLmG0dZEFLH82pfjP28SzpctYP7JxQr
W2rGPpBJsBH57pwOu5m2JQILGeu4aYFz+6UBk8OChe6C4Xu3oAmEesgmo+6ymGik
wCM0w7JZGB3Kx/uvwHHqjRAhxe07Ugpc3L6dR4uXJxC/4+4rJ3YjXn/IG+zQiQP8
TgQKwP6KzwSSwnIR7wG625xA/IiPZR4QLJ8ZAO09jdb2aWdJVuQxeuZTouVbBiKo
PPDmg34z1A9VWBJ3sLRemTCBQfw1C8UN62893gHz9iszQ2cWm79jcI8kc24bza//
/eWxoMHfziimmbV3wPgCs3byZsKHohQXWZpZrfj6tngwBJWpR0IqVU4XMu7OjoRU
wlEsXRnjNcxBb/pxvpX7hnPriiJJvS0OEZjWl46qrDXyBbceBJ9dTqU7uV7aG9Z4
cmVdlQsqYUw3PLIaGensKXI8vet3K7BblGZIqAblrPBJNC+BU6ZFzIyKlzTfUzah
nKryVpeKzPU5uenSvKH+9bDPVZa1m8lrfIaRu/lTS6yQ1zeWkWPNtwNLiG5VU98v
2Z8031iCuBJO76QoHAm2VprmJF3+/ymfM98CCoQDT8eV6T16dGEL5EhZEr81dnVd
+6hylO2zdXIVuVvcRdudZG6fqYx8mjidOggWnh8CUfqwmBhEAHcgDnAYuIutyQZ4
dpCncEBGDtJ6PNZtcq8cbvFgwp1aOeTkuaS5YUZEcv7LhVqgmGxF7CQIs4pXa1Wp
qpgVCBSh1pBkBg7VWa5brL/Uevd7d7qFMl8X3b9RE8x6whLyqhTALkL5z/GkhnH9
V9jL2hJ5zvahqyyzDwLW9wU1F2DvGh5fqW4CBYfH8UdyDz20I6mgNMuJd2MfIEQm
t6j0N04zHMkwwJiSJD12QD1rmwTE/dV0y/iAsNR2V92RDZxkxvivqLlkLpulsico
jA4Nn8vYlGi05UjXym8zy8nsLm0jIvT4JEXftNf1uyrPsWpAUcGbKY2QyPldE4aQ
Tyv1ZdsUoaosWeIjVfLlkGibJ3Bfi1ZxkhoTd5ZALC20p1wkSm+6Rk1Vn3Vxn0kZ
2JLm0qNV/V9IL2Mh+dhruCZmBIkwEu9IFnlGm+QGvP/yQ9HHUM8F1LZE5T4VuoB+
8bZlnx0uE4HFHVq7GgT0nMFYGkFFmTxrTg6WWhQ0pApvYncTAjC/tZnosc5UjiBg
JRD/CXUFoVA6XwdFJHxKVUdTM1cWjO/cnJKDLuJcsfVsfBPwTJ6AQqhjQtim8kt9
zAW04eJJXh9D7uN/prSSsTOHvIfZiaY3SX0CLTDLesf+67iiRDSAPja1mpIWBtCV
Vu6RtAIrKE8F0JYtfjNnaupbq6QuRjwbpYHwjGFtzQTWz6DQji9vGTBfsWmumpmP
GENW28Skf2oYzfTrA63aypXRnAun6eVIO9iD2TsuCows0QrdnXD5OTHXt6ebh1it
h29rg4AzNe++iwo6INwGK6fmvHOc5D9uOksh6q5twPMTavaAucRLMRJhh47iYlIC
dlW7QZsHZUyBOybi2OLCF7Gl1plQyDoyU1Ew1fcHpmM+c0Mqk6Gt7sgwizrSwQmF
pIrtRaoCt665BHYjVfYQe7DBaIbopXP4nPCl/pGtWmk58WOWfjhg2iGIXRJgblP1
bdaiRNHJfnQSnr7e2xbeT36xtPDEYOFEtCZXLfPTmdSqQbUN40gnuJAI0C6hHaRX
SNEXgCdvH3DxhNF50eYZh3usXomwvHNwDWcnXSj9d22hAmlst+sRa+DpyIcl3GQG
LHIfz6PrIWanR/m+FtJQV+1JIyRPk0ZO5JsXInr91LEXrusrjNNPa3aAFZ9T5hA9
xSodLJ9gKVWLOjZ5r1iF5JQYft+aj2h8ODHBBT3WVUuAillRdiNUdo9J85OOK4UM
VpsMy+BWHWbB2upJB2M+JPpBTprT9QHPJBK6xBdW+Sf/u7RaU5ZpkwkERtr2UtJZ
PE0aurM/9R1t1astaFooSLGDNC7TKhW0uDjflXzlCpSFdiJU/s0as9DtUfqSpmBY
4YBOwtkKdbyifIXSAS3FZVSw3D9m8GumZbvqlIWmpaApo8aBfNmBxxHfZ/r2omvX
lG2TAg8Ya7FTG9uYpTERHDF/7P/srMlu+rddNDEDqUPSDbY+MGscjkZnrDeXxfS1
3W+lRwyE0bN5iNm0MQ7UA+1OrjA5s0Kp3+XUJz15G+6lB6Z3K3UxouCUK3Bi9vCl
7sdw862ws5F0ONAvqmZ0bs5f8FSZvoMpVhFNtYdk1DrZ0+gPcEnMV06YHhkaygUi
5RMyK1p+vXb/2xJb9XfGM+emWnd4tVBpEuxzlv/Yl7FBJ5sCITGMGCsQ1JZbMHj9
buoWZdaTPGpNmm7PEIFskpTWMmf/FG2JPiMksWoeYDqrkBXgr0OzcQsyN45LmM3a
Us+yzo/adZijeGTQh5yc9qRy2X/lPRn28fIDzlp4C8vwFNo/V80ZYVhA4uPPheXp
k0T4F5NI7fDS4ZC9dzT5+KmmtG6nq6Wii12yMbzbIl1RdQc0lA7D4p0GbvtNCpwW
b05h6fb0MlXf81e1QiiJhnUKum/CxxW0I2N9Zti0o7teB4b6roR+14gdJElZgaEL
Zffvkr9VDmFYXLFsIY5uk6IFcVyDb81SjqtOTzPFZyPdhht1dOIWh8G2aHSDGLj2
T8WZJ40rpfwIODVhNSDDWOc12Mr+M6BZddLtLlfPyx3F6Bsbu1RdyfHi5tHpYjVT
LzlGGqSYVnEZhgiyAsIPpLAA7r2P09niIeMPy8NcUmAgPQRSgPTurI0bZ3swm8i8
/WCQys38T+BH6Jic4n8sr4exHWICG6t4DYZngU1c5odObKUKTwlWsPSdNUU+q9X0
QmdHruJV4QDykSoYcxxt8kH4s29dqYrDB39u6rkcJ2QUNvrBBRuTSQo/v927Ccin
srKZBw9RwIR0x+rkVoFbD93KnXOaI6kF5fxCAxM45Q2ARnwVxrW0QAljXQMn5HRZ
ABR7ZdhUpg5gNZWISZB1pCFZhohBk+DPFKLMVYpADWfR32uVi6/rtTFypL1tbuSw
AKrwLODvyAYlFFqctOIssq8Lg84TlZuJse/qJuV0nsf2Gsj2dMEHyCu5UO7eDXif
EwjFObietUilAVWIZG9KIB+lVZ/TugojaXiDOmO1yMIZXCvom61dQA85W8UOWYFX
xROQo/mH9PuC5Ra0oXXeLtZsATkz5irf3HrT6wLPi7IXA1FDUbExI12AYSGk6JtK
ElD6c8/k40j2xiO8eCrrOwsYAWMDQz6Q1crDTGjXPr3beRom6hxo7dfojlYCFAEb
wavIv81vA7T33w8Scj701xGSp8YiidEXh61zviO3o16N9hl2R9OmYp8jcSY4GXjs
cCEStWEC5bRfPnVm0MkMAwDBhhHfn9vR7FqhD7WLiDK4XY9Ytbn3wgWZlkQK0VW/
pB0AtbFNiF5kZEo8jw1ezgATWQYROBv5nDXeFv0FyZZYLPYd1EdICh2wuDNA5Fv4
F8Hn+PyI6Ip06vJpYf1SKK8e0ewLjzMdIFtMlzbsqpXiPW6pF82dkRZbU5WPbLns
Ciuip/cujMPdmcFuLcMglDdAzgXPGDylBeFIP43HWLaiuVmBz2jRoGDTuTek5luC
Q75xnzDPYjqNOyqcL2MLlI/Vsle1RB26Bu4pDtWqdZFHjdPn105KHkUSOlarEyKA
65IKXJf7nyuSkOio2UqaEk1L9YWXMBvV7JnS7ug4vpisUjF6CVrpoi+l4CPzTNsl
59hDYcCl8PGdNpvrK1YPkLBoMxH4bDC1Adht9DbiArZ5CYNJLgdrli6V/umwh/9U
jWGitrdc1BJhri2jGs9Yqugbnx98uX+9kRv06vqURXyxmtwPyWrlyCB1hnftu/Bn
Gc0uvM/31vpS44Pnnf7ea8w3+KmXcEv2g0wJsMXIPy08ICUHTgY5YpOOhO4ISen+
hsVv0t3mGc7TbmhLyeg1TA==
`protect END_PROTECTED
