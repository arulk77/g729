`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aeWMSqAWdJBQSOBVeo5ydi2+8GPzzctoHfJCrbO0pGTo
sFCr6U7gYXsg/Q4TMlFONsp2oorTo4kzv+7l5Y9SWTsbCeVDhxV36R9SYEay2Sis
g25mXUFbRTif1hU2gCuXSLACbhuqUbDqyj0T+v/484+ibhl+UEyO4/uu7YHlCKso
jRay6XjhiKJnaJrCkyWxs+6qhSdb2+oVXJ0+k1gTpGLTDoCGf6f1W4gtUfh/1zC4
1jAX7V8VoEgU9/ofCWM8Fdaq7MsVIbaCOzfTXns4UEhC+jUW56V2YYJhjrkh+wph
wMEQQvNsoFAYjzCx9gJlqtoDpWE9PVSFZJS5hjl5S5Yg69v/PrlYHZe3wewMojwO
5oZvG5LA6cQlf9zG0CSpdeuqCgJoI2SZkK1hcNGWJvXmqV7PMiDzNtXdd3e5navN
3Wu1abaneduAfle3oueRYKdMV9trWzn6YZH2xLLjFJuBvvWgxVlJka64uuMmjy4+
jPInbTy3e3/SQfuWW8b/18GRF2AeHaZ2fRiDgzntnLpPi+S5tjv58NrXceuoiXZP
oIeoglv4/W+2Ez8QwSFoTqsRpziwKuZuaHhnJ769v5cYQBNieGs2Sey17FAKfFMq
ADnmiwUM7BORAGe4EV0gTH9TXMEVe65gpcAbqVeF7SSxV4XtcJ6HMIfhbu/UslH3
/3MqajFRd2tb14NT/ZxJdFzD0IbG3ff977MQEkJ6/9dzIeHfmHk8UzbkwsoiSK4r
7g+nn/F3774mLfoEjoWmehD12J71l/rcbk8dgKssgn3s1v0KcpCzvS0uNYUFfFwc
cV7CQJxvP0P2i5/g1oxK1ewXiE84gAKg82Vw4LCmUMFivmzdP1RpzRZ78d7Ombre
sfei+b0gEkse9ZT3cA1La0jauBIPNJDh36ntWM5F9ODKvotwtGf7YwUCwfyvD9+t
0wIfkQvZBhjl0LFmHHtF3T4r0FPqmw7Ah7TnNppPq0lsBxJiUWlv6T9yIt7jfmUv
Pi4rD1YAaCfmZ/CqG+VtWXCpQa2CTpUNru1o5GdbCUF9W1dpFmdKBblBlszJHto6
VuFvS1rxnLBC2Cn2OcKuxXAjtEGIpCkdQLsJudLfP7ZDYN4qA5EHdbLB1wihwIdW
om7U9mg4mIB5OArgF4sFcLvvuYIjnVwMblaQLoBnDPeMPDLTIWtF8cHAfnTrCORP
ydMnfrIK5Y1EkU1lb90oHsAUodRIe04ybonunxDjDEOB3pk1pQLQ5CTMvwpkI2TG
mmNHDCJXglEN5GVbdPLRL/q3QOVc88z/Q5k6GVOv3YUkVezQfwJ00aFgkyai7Zbn
st40MCIXeRRH17co5fWqrN17vAalypmeQJjgoX7gQRZo6Qw2gcUVeoje6Bxag3T/
TCYGEd6fL0TyqWJxLQQh+S76wWoz6fdXXnPxBDKq0C3NyogJS3CPzCSHbnF4LjJx
vQw9TzXzZXKEDF3+v7El8SwCTBA/jE7yapO+XWqCvAx992XOYqvkp+5F/+Z5RKpF
MB7h03J21qLsTv0g54tn/WL+3iPNIdHZkROPpJFy1+y/Nlh1dMkIlUX5N69zSooQ
6zJmKmIEiAsHCiXHIvG93GSOyZOGRFs+cz2CRI32bgK/CNwN4zxRtkmnUHl/WGj5
TQBh+8IYRfpf0wtJE/k41rO7XoRmdAz8ctjMNWQJPZMvO5NIfphkcOWhAeHfv1nY
lDawvYBu6G7JTnz8Bj57l2G3tbbZ9bi7G97Ku94Fm76I2mjRWQNaHhzZ2tMqtOmZ
cMApN3KUqOoJ+wOEFNk7uV/FUkrLKdPGcEp2iQDcyoWZqGr0iSPN2fvKV+RsyK9N
0Yvx6bkvhUQXwAImfUd0gl2ObXzF5RFlLrPYzkIpl7KY3vzWq7davmRhKQ89dBmZ
zLDUnHDI3Z1eSxIsoF1dMMEwgRqXS4QMY0735eM3m2FWnxUO6AQmXPwIqumCEMl7
57VPlxh5aB1H8Ig+fRR5dUMJYy3f7A//ELYgRdHBjSCUgU7cOy0oh5MHSUQ+xIGs
UBr4NcD1V4y1R489zuYyzxyrCPlBcwfH9Ka8/zaicdJ7OGDDt2H8sLfMbDfr3Pyh
J+GCEWTd1rFX/OEvw8qkZv8Jk+G/ZGlZU0Sz+zl199GIAxNVIBy+V0VYo6eIiWKh
nTiJazOTgyTm5XkSBBVp7RjWodJxiYvfdvwsJkncOtYRRl8IMcWEtgoBMF6raDCU
jmtpoiOWAtlCEHtPIRsPyyoPELDdy3mmvyl2mBxpJ8GDf5WtRY/0vNjAS5jaGvCx
/TvZNjWakOKbBra+5yx/Gm5J0ztEaAah3EFgHktZUW75SIZcgmpmxc/3ZkJV8n36
l+KTmM58rKFc+IELxow9DFAJZJx3pDxCP07OTjGDr+UmQpsYPvMVw67M2Pk2I6oX
Y6iLonylHILe/it/BdSBL7OjuUQD1XCZlrWjVGq24fNUE5kOZkdbBv528DCUw/uz
2yALdQBsFviyfW36OwRsxPotZVlp7FjzodNf10JcyjmiFOLwOBOw2xIm2YpO0nLX
jYLf7YGKfOii8Z8NMzAFNy5KTxctxV7mga/kicU3qrgzAT12ZyG7DLFFgR5utDgg
/8uSDI6XR8VV0eTSPHxrGJwIlACrk/qP7jRcslN61yZbE6AnzawM2H84RfoJyAfJ
J05snLw//K2AD7YE/DvkC6f4n22vpplg+V3DKrmRzMio7ykt5XkTsvMmbceulRyH
JBZM5yrjs79kXwRl+retK0XncJbOcxN3tyWqnu+xu7BNyWKEiQGUk8te9nQuxU8u
trgbiVP+pSXTj7rp63nrqkFmQp9pnoQegh+DDe+OmWsQZ9XLXswTeBHDi8/xNPjr
WVzaXJ6OxN1fl88DQO8xlYe+w4HsafYZ9JAwTsqZKlSAwDu7Pqd/WCCm7F7Sp1Np
E1AJ2FG0LOnWm7ILWlLVctD6hhfwjwIz3sIRIFFwNgh3QiOwJijNrpJqHzxNiDo1
dBckEXHItf11e2ImdwLqTTtkH7k5PnGn9IvZdE7jmDQmudNzC3KxqN11yFv5ZHRS
lrgoeGy7tPp4BhJudZ0eii7Ee+Bhb482GbONbolZ4p8n2PZXGBsEE3egYXJYIxur
5Ch74taHSJKOyhBpY/ykk8urrN6N9fIBt8u2ajkTw+5Dv+MBEszMdq1QTvO6fYj/
jsjHq6xKGPUoxIl8zVe3bRuw/Jhp5mZdG19U7m2k2wJxqi8Vsd+aXkLamJH0AzsZ
vr9qeN9t8cfbZzYsrwTkq6NIRxXPeBS3xdZPsMcgPOIUcjPkSw9BU13nwU/A0ZyM
CX0IU5bBhyBVarg6MH/1Jlmbwd9cGygaawDxxGYXUgUe8bf4KJhfuH5gn6QreXm7
F9QjggLTuSEH2CtOMU9ZXCc9s3aDQ44+uXfj4C1C3iFOAk66QZC9lebkrKPjTb/B
ZBSr0ZS634ONg9DWuoSN1frtGruxxVZRvHKdcSTCunsGNyRFrDF/gfgXG9ikaS6W
8dzH7aTi3MWmGSIcKmVdLBr7DDvxONm7RXRC/XQh09EKHvCh4laXZXqHWhSIGwAq
d8pQLvhRiE5YeYd7uq6Yc9kp5t6JrQoUYgVOZTegvZFWqORFTvxeznDZnCSzC628
7U05OD6WsBr7wDE3m5+gFhxXQsQVhAwWIbk6FKC/SsKf0Eu0r1joMASoSiLisfa7
xV6ITDQvwPUhMtDCRJL2lcuoC9wRs1HUfqVqVx+SCErEqHzqHA0bfSynInSuMKli
gqyIyRQrW6EuKLv9pXcwoZLPWCwkzn/x5aFSUwxX1fIPVsT/+Drq5zj+NLNOjvpd
deXGP9f2S1KExLHIEkZjXz5dVnj5Hv/RyUriip8Ly+VVpmKJi80Ifc1hPLaKKnjv
KM53a2vW1cu+/SZlQUT8rqtWrdUg47giVGS02dEyPra+m1CQ5uilc3W6PaAL01s4
Vxujp+8Adi4tUyyzHAtBsyl2x/ZCL+O2q47RrhSgwmt6pD9y+k1tbam/YLEQm8Az
Nt3Mj1OnpmkoXvPG6Sk83O0b6JrBnKfObmLOVlAQbMxMfoX/OwpLFf7msyeTl5Fd
bptL/m8ECKBh9Qm63sPmFQcDlQ1TENDBMJ63aCU87eSmbrPRQtJOT5cA/YG4K0Vj
nhOjMo4P0HflTnHpcaFDCyifOAjT4z2SV/MDlkYy4olefdMZgkbXTUPAQHszC/Tv
YH5jNWxSKYM+PnBjX6GFJMCXlvkZevUZiV0rTeTFi+ebhev+pCLfWiF0WHs9mbCS
gMo98jgaylrHrsfKxZagHcQTaBivREeXGS+lmjDe6I+QIhNoWZhifuodpWCdyL8J
KZX/hA/fxSQTAD8oGX2E9zci8AAZfhpTj1t7Ow5OcD0fqYnB6RY3DKF5mu/Dq1TL
wbYNebNr/HinIbgiTpq1w/tonNW+PHQFfSEJdmpzIroiDlaIOiFS7qe+r0O2hUJj
3nPlzK/jBua0lWAGVifam4RV1gaImWyzHFCw/XZvz9m55nJ8S7p4jDMFUKvbkWn3
58VSo05hRXQp7DdtOJnUVfjsXdUqY5a+WstA8s7eXd1nclCi6F/ePgAx9WND7sE4
HTskJct5IJPcVvQeX5uA5QhG1VOWyKCQJYikPxC2LmO/6ZlonSw1gpWekVafNZqP
4VjtQNLGblBLuWUTbWZv5/49AP5pOaagxfiv5EMBLA4ZaTeDznYmz+m0djtWeo7L
/qIqsnKDWr1EdysPv4LpxKOJSZI/OKPIse7QoByjI6iSR9Pfwb2P+KE8dR+KvJvc
hPZqyM/lxoDNNhefAX29Jj8+xbDnPG5ttf80LEvwfKrJyoTpA7UsJgic5+gKVnMX
w9E7NAGQeVr1Xo0ryDdK5t2SpDG2db8oZps9Fk1LEfHCLx8V/0Qsgchqhy1NAeD3
HT1sZ9UtdqfdxOLI+nOC6DtexNKwdMKK1wqcdFBkYZzMzYJ/xj+i4+riXOGjE8hQ
Taxr3DegZBfQIEoou/imvVGARrflu2UtUAGa/mOCZ5c=
`protect END_PROTECTED
