`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGEFsvQKXA+wXhtK/4PMRspJqEyefQd/WDBBTL5SQFjU
c9jWxCST4HKYTuhfmJT67isu0PvypxX/mUC4qrfKmGaVyWtB5eT5ajVgTFslOidA
LjhEuJM18V41RFHWn/ZD89jA0ufAOvKQr0vX/oCCzdB+9IzG7htK7RiTDRvfuFUI
u3T92SQEIZFg4ZjFTtyJrg==
`protect END_PROTECTED
