`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4ymunnioox7dob3wFIJsu2A8e9NZ4HuWE6ntgSrk+SDK
ksBNT+Ik+4uiaQaOpWduwtVGKFBF2EU2bKTH1H0snrmRo27QVd3Zy5VhN/vKzaRp
oakGPiILqhgjXU/w6glNvgzVPBEv46UyB0JmBGR272O88JZIf4ZJUi5jx61r/jVj
N4P4Liu4gdBV7YF+7z3DxpyYUcy+gLKcocvAalVSnIRafQoWsM2FdJFxY+oZB88F
k49/RF25ZpsRt5g1LIsHZwCTgix4luK4QEGQmwjJkEisYqmm5eno5tt2j4vWfx/B
bHmLb14D2TDBW4OCeFcUTCL2k5GJHxH0YIsDNs5oK67LNrZathUlnTINLD8yktwc
ehiGdnFE28jyQta5dlEn6w==
`protect END_PROTECTED
