`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGacdNeAJpNZDrYLRF1gG1IdbxfvNB2rZhZa+57C/hNK
xfuCljJ0TkxDeT0NuulRL2+c1Chw4gAg5RmzAjOQeA0bXu813VKIHgykc4Xs84nY
cfUWBz2eUjmzXIKq9kNp3xHsjvJcoQOg2gNvcI65ZSTtA1h/IvGpa/ESOKSAEP6g
2P0XO1+GYYmBAm2Gd8TQBMkGQqfaUxWj/y5tEvWzZwZQRYY1oQlAMVSS4uJ3hSrX
14BuTbh/4AR7gr2NKU/E3sX9y12TxjFi8D4GMUZLSKWeh9+7oqrJCHgWuErD6MUg
2zVyl65MOGYEeD6rG8TL+/YX+qLe355ncH2Q4BEj5dzKNzWmSfOHjeg+euILTkYF
E8DFBYYxT39MvWULd1ZzapM/5EuJvGkFJJZ1VhJ7K8/+5PzSsqHm2tu8U4HFybpl
V7CWwDsvTwnoHZ0JDQBHjmU4eUWHKy2NXSu40FVDolcfWdpjKRVM33X+kwi4lFrv
`protect END_PROTECTED
