`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHBUoCSgteF/1YK7sHLAjtEfhdKsT9JF3WdCfj4UCJek
j+sE51uOZsbDF2UnOkGt2VeEr8YUOgRXhAYc3QijTSVwS6Y8Bz5Q6svXSnuNEP0Z
Pph0EJuMaMUqRG0ErTL2+wCSYGApiOZvsn4/fvqI4qQzcl2hBSinZfDUS21797x3
XZKd16NgCQ4rF9K7SNoF8XlzokYW7JuXoOrljFGDGG2RNqDo6HNh16lQLNRpr7Ac
JuhJmPjRzpT2zeuSGNW1Npq660bCHqcILU9nq7kQV8TDN91NJnFG+nf9Tz5VEzKM
gkDxTNm660xvBlyLzzU6sK//2M3OdkF+7USGTmumyTMSUKqJu0qP551LOgy7Yyu7
Mq16pw7ctik1MRGUuRskZd5dwXqNfvPY/msIpAsjzpMs2/lvfEJd7Wvcarh4WDa4
C6hQ5jiKijwcYInEmTtmGsBgT3wuRaxO0VCFYfn5meTuvZyL1H34xEq+7wmvAk7e
6lWT9uEc8ApPblEvfbrs3BwYnsWmQGRhzrgdMNhf0AMZ4RBgofnwI4jmpBjxM+Hf
Gr2wAGRBubxTpzX5Ug9IpiDDSdZ21ofRDn/ve2gdNki19SwgscdMIJYUEk9jMjrT
IAUFJEspdVYYNblMRsqzHgosHCfdPGkLdIpfos1iiH2JWzSD37b72xA7Kxcdj63x
PhJPgC3YJnMgndqZEz4CqslDr9xl7N6tP0MUmnCGF85deayJ69DksvdI9VMUGq2o
DRdchCyB7vQ3i16cGOUiyos6jVaiR34W1BZQ5vTCNXJKVzH16y+pKXNU57OrhDAG
ZJVIKbswSMh4I8S4Av8e0p2cb1bFpCa6XXBlxQWquyg=
`protect END_PROTECTED
