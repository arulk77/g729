`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
iEBzYe0UL4UYD0k8vEPLRNAyFyYyYHZAy6V8Jcf+jbeZq64rTWYub8Re7EQg8A3x
UwqY1Lf8ye2KVpswXQ+YtauBqLdBn7h95wPybNvxu7mA8s6ynY1y8zNNvrjPbDTc
Ly3KkodfHVGsYwSBlwzvladR/HChUSdZpH8VJF/kytRwN6knlF9SPrG6q477kUnc
H9tSC/TlW6KLWgKM50oBupZAKFP+FgY/S4Sxzb6yBL37xssqiaBCS7d8eMHdWKuN
4thafjnJd9Cv/Z5aw4+MguMdWX41RYsa0+NkLDYG4mo=
`protect END_PROTECTED
