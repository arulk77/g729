`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
MhMFLUc/Ib2eizzQqvDtDsv0HExNxpCGreYs06MpH2//+KDqL0eDzaXZUHWbxXlZ
NDbJhEOFBUl3SaLQWHei4AKu9AnhB+DDGMcYqyP9pnQlXElUJgeeT0SkRpDZB1Xe
yHjRvTBnSuQwQX6wtpMhDeKNFlLgd2nmifylz6vZLtgu36Au5BeVDx1TCCPur9Rc
IUOvTENumgpyx1SiN6FjV0KIV+h6VMtNs1yk806tJX4=
`protect END_PROTECTED
