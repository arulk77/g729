`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK1qOr8UjsZ86mR1Dk3nlwJwVCwqJUrXQ++o2YO0IM4W
norf8bacEllmv3mUznyk6tBNoLdXDxsuD/MW0CZnVBuCQv1UFjbIDr8q3Ug4iG2Q
siGF4cL4BH6Vqxz80guVuCXIWbApUL/rHVCKE6BOyaU9zjzvvqVM/ud7sSzUeRIx
F8mR3Va0sNJEruEiP3Yj4uzXu9BdtK7/Iug5H3BnMXmWMGYtudS5o3F0mvA5dBG/
ZKCWyEt0SvMomQZXo82NjTbEjNyI8KZ88RvTrLStglZ/2iaQZbNmnCK+YddqOyg8
BpPk/niEwyg4+BLuHV/GrLZE9qPBUvkYPsCo+F58VuGAZxAD0d7j4jF7MsxHqr7T
oyVqmL3/PqOkj2iAx0cjl+sSqzWDCOetwdSp+HDvSqG8c6ZvZmJRI9SKCv5Z6VZQ
XtMUlaGc+8wyWHY1MEWvy+ngpGMcNANCGajiFDVwNEUIdAslpg9wYD+I9JJ/SY5E
vDLVhJlsPEnPlRMrmtLa66Z0YgfnF6jAdPjdo9jSYP5M4cYs7n+/ZtJ7dYHZ5K4+
`protect END_PROTECTED
