`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
z/MvhNsNEy8LRPKbHqjBJWPRLkSlfBlM00pKVAgftNBLf6SvlREs7Mprcoz0e9lk
tJg8GHtCRcLZFZfPkac/IW6/7FCOoh0nUJvZdj+UmBmX7kBqo58t5bPsAa04df5o
VxjGmJFBAXlvtxpeXHQcsG5S1jT8BAedIkLjCjrY0riTSFf+gyR/9tlMSXmSB/mS
rcHQabQokRGIKpm2AmCFkKHBmdE29p/5WoUETYvQJEogyG1ELE3ymCZlokvi65nJ
PqUcoZVCU3xhBmrE09zmDKBpT0JTzAuLbB8Ztar2je7L4R24shTSsB3TWi81Yk9Q
Ik/YRVfLEMws17KHs5z44BvjlwaYyXk0UkDi424+gPZ1fAqV56LHnEWIvusU0bOM
wdRnxzFaWBanu3WSCKZrSF1tSzNkayqtyk4T7BTB9nA=
`protect END_PROTECTED
