`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73CzMP8ImJ4ZSijuv3HzjYXPhKei+BsFMQ2RWruCAfhNrb
prZ4SHN4HoRrYiGtzBTYlOEYSKdfwBKJVcJ5hPwH2PPU/SfoEcAfBV/VooIRHP7P
SMp+kueKfEo9spJRCkAyDt25rABaDjlQDFVMH+LNBftKIC2S5nc2b8jPUfG+sJf2
yjRCiMR8oim47+M89fGC6N03IZpNl3dhxsA0kGwHxmtK52BLck94OrkB5xFvLtqu
n8e915bfULwlih5ePpkxAZrHQWwAP1aUf175JgxERcYwFxjD+ux16qwyPkjVqh5m
5aJ3sfNdl/CvVtlnNJ9H3XxM1VVnrdqH/ts6dgpR7BY=
`protect END_PROTECTED
