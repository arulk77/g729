`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zQnkP0DmtVqn87XDqbn77uM3dNrDmEiZxmkadQEdL0e
x4A2Rh/fEp8xAuB3vScPjrZm1ua7GXH80MGBQDaZ9NXNbhvqfD/6E8BXNS7qVe8g
OKeCs4+g5gw2UxcZkZ/NsK3IHWMXOaIgsbVW1dFO1My3yBTlrGrSEC9kg1MDXU9u
lJ6wHFfYiqvx3A+Q80glTOcM/WxlGFlVMwZ91QlbH1g3BBaOoZPsUL6VTQuvajZV
RFah+WhgLvjjl1hcoAXHfL2v9DELCapsSLEMNqJW3dTPOaz1gWntXGkG2F/hzXO1
ZccTai7raOfTBObs8wTI23Ylo6GYuUqXdIsdHIbzal73kNMz/B4nxPvwOvdS4lGA
8oHt9jboNOZ6PQcl5EN0RQ==
`protect END_PROTECTED
