`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Ynhg5esTbEMoXi7rBuHQ5NtiFZfAG1qACQ4zUjE1Rd327vC6fSyEObjycbfBNaLu
C8LoLnLepUCXmb+MWCbMJgCwtTDdkllMgzb7OBVmMN1gGhX6Vg4py6BpPb4qe41Q
Zmi5ZzYMj9mKqAFquVTvEC+bjhR+JzqSTAMGwYMmq8w28Cdx4D8PEceTt7udVgdr
`protect END_PROTECTED
