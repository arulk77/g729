`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
DieLZT3nBzluOzvcY+xOB3RdVM+YZ+NgJh1OHUNy4+roKBJTvuR3O0uok6t7Ivsj
oCZNipG5riGFBS1zODbm9sfAD8f5ZmVA4cjMkB7UnwB/Yo3rOadLvfM1YMxUmOfV
7HfG65gaHgaIQDx5dvq3sezJZ2eon604T2d0t5Wr5s2b1Si4MbZg1CjeoTtcxVAF
vph2cHOErfOcst3LUYAjtCaFipPatjRjgcZnPO3mAkqdh4+G2p7DxHWA5iirBDLP
QnDy6QMci9TD/tszZZG9z52yp1CT0vzoN/x5ueF/2dnSwBEvyglvJj1g0rDwqYbz
iYW3Teury2FfI9Fs8fhu59pvSnPwkx3xcLVy6L0S4N4o/ROFMXTHOLV/4ozAoAFI
XTLIn5xexFEkWLw1Z0IcqtwIt+gfKYQPwjN17eocoIbadawENx3YWtUwjzuhF+Ps
+EdQ7LiUrAWeiwXPVqhBWBD9NAjAeM8dCg+Kjzkpcbc/bBgpTvK5CIs918fp5SYJ
p2oo/L2VWJ2w0bEG+EmQ5G5vGtjXqste6nHA3NwLMRbfTjtPjM8y9e2z3dQOjv61
RppRWuqeowWklWlypuXG00mxGcJGLjk83W0IJogQbJSykqRL6UQ3M4JaeENrsm8U
6HBcXj2NNnRDjnX9rPIIddV/Eton/b/sP7tvpCphwIasO+KXkdlE4IlNjYaNs3xB
iSr74cBDJZ0e08qLyEeDky6lnVXRzCpTtS+6Hxr1De70EA+TEnCzKyCCHPWwGgT9
iUPL8fl31g5Zk50gGJIy+zbKH7fl/9hUtE/y7hYTzg67cl/EXVcXMNpDIgiqqYFP
GqoDn2V0id0fU+49IeNeJGBRMCepCbhz4bCUuV/2ZaoL2MNrn3P8+3QLQiWG5F7W
Q3QoMFXn8+eqwIHs/K8qKpBMOvSU4Pn9kLbh3pLYfpNVv7EiuhnHt2bmmwW+qrxV
KcrL5tc8+SQvENw9wFlXZg476EjQj7TxbZDHK8NIbDy6ebxHAv0s3dLtfkQLxYQI
pk9uG86e2PEXbjZ+gNjbPl0SjnCWA4/Sxy3FpU6B82j5gfO/cbcB8oGXHePmjERq
I1kOB9otyL2hqkEKNF+9Qpi2Plm5AFZ5SRYraj4MBxsT//0Ok0Z8wl0SW7+cSqre
hgOOmESqi85Pe2MTaZEeoTGbGTT9U77aWOj0SqdvJNdWzempf9bJS1aPetgJsyXN
Ipx94eKjXEwfYll4LSgOCNCWQiKDE90u8r1bRm25n1eK47/osY3aStzt9G4SEOtB
GksLNa6QBSpOOJut+0K0g3AEHbZhpxu30VHpDk84TgMHP9SAu3qGlhML3/gp4xj/
9580lElaxVEoT6pi6Tfx39CLjBJsX9WAjMznoPyc/TDtpWQO6HF9g8w7PJpeQuip
arcYxXO9M6OFRxw77VrESOtK5keBx3+K0CzGURLZahXqG9klyARnktX2zK84lpr3
FpxtFn2iUPJQtImgJW2PvD0ciQanmw+q/CyritLD/yDPXviao4V/Y5x0ze0Mci1N
v2H2X99Mw0gR/y5Od6gsMNTqePCcpBDSSGQSEvQTVyzYhtiOQdb1GEjuKVz+qVs8
v6WEzKWW46cxWHaa3VxsqAfDU7oZueSECqnbeI1YxAQe7V2YbhbMwP12K0TeQ2lX
I4ARsxPyroyLz8PdhjPNuojgTgaQ7oK9QCAc9mgRdDLITMU9wxmq9xtt/BB+8qau
J3eNudpZMf7fZCTjfnWRi2DQsUnyxnNAueIyLxjy7SpmkzMi07GvtIcHUbpnxU1R
6XKBiNsUTdw86pDB+AJK7ewEa30/x0rZZox4cqyWkN1OJovon0HjcgYRUqMtN8eP
hBFOpx7IOvKZ8+E7SOpOPDcY6wRf/RhuOMyfaleg2jeHQ5wfbZdNAsz8LodNWuTr
3a8EB13Kg3Y5MVTYfCFRkLbkPQvdCWtJKT+MfeivTol34a/ruFvQhNxhUw12Mv5Z
SWoV/L303OBr1j6ARCgpdQKGND+Dtk1bc7wdAvQy0yhAxbj23xS8nrL8nYXVJ61B
xqnrgZtnjzIxyLLo0h6fh6eJsyX+3EPs3ZyBzmo0bpS+8bc3zdDkxcPci8KQtJBb
kMf98wKxH/xY675oVWxfN3DKnSrMfBKxvV/jjoG9FgUB98l81GWNhpXvDmY4WnpX
CzkCU6Gpu7UOsrvpYv3V6EzgHftbcYO/hv1JHtH0SFzv+QPghaNUDB5s9+vHEcQ/
UZKY4Pr16PnJGuyGytUc569z4pTG3mTBTmq8feMk85bMRnq/Em2zUjwIC8kYpDxh
e74SZWIQLeEBOxPzk2weUPnRbwocVjPIZPyms/Mw7OgEqlnjDnG5Z6k1G/Ww+ili
hGiMmRiok4rpcZYLJOZ/6Kmj1NTA5o7xHNrCZjVot52/AI6s+xkey+pSzVTLXh4C
syTGL28JQ2r28foitr3Qz3JQk0Gs9Y4YCxTVom1I1GLXXYx3llQkxk8mk7VO2aw8
ERQZL+Ss2LRX6EC9fT83cvyD+G7ABy3nf/Y7nciw57AkmID7Zsh8xWeU6jI+9WS3
w6iWQrGwT+KmagEDjzKlIc2Sy/SPwgxGjTouG+1T6vF7sQi+whYci86mnlk83xVh
JQ41IGyOYxkua5IfMagl6Bmx+Wg9+oa5y8sprtWoDUC53WWvA/I3iWA/J9vJ1Ktc
MEi4fsZODT9XX4d/f+M4g4Jhgju+SKQwAfkif0kde+nAXSSYcO2S5e58qCt848yM
gjNTiVx3G+73e1YOwIFMwL4FkSxFDGMMZMubv++BS9IbgvXTvUlTqD8n9pN789U9
NNjnl/gx5yZSDnOQYniA3zjulm8pg4qWUZt9DE8XFiqnUeeQ9eGxXVEhrI+Xvjsn
DWaasndPUVoGSwZwlW+jOOcbtnIcg2Ke4DuX8dgRzmbo1QKHhSz5OAPigjgWc4pT
BKD5n6jvvKMJvBSWZ+QRN19CalJpVfH70IF1X1erYLsHxbfCQgPBbaBjfQ/l3oGn
Osnpzq5RibZpE42LPQyhCYgtYM2BQY1G9mciZ3dQuf3+kcS4wvhkcmwJ5V9BVe75
z4hR55srmWrmZnVDBv2XIfJgQLcqQGq0KD1/ktyup/ehbYTjIdIqgoG8PPzf/cH2
oj2ZG44kuvUcCFmznut5ly/rQ7JtpOe9eKcuDgRRI5Hu3QqAAtUyTJD8psOg4VLd
okEtDTMChS5LrspXYJpBSIc4NCrjwM/mou5RK155RKnUQxV4+MQWsKzfrvptXj4o
SzI+48yLaN4sMIzEEftllkeTvkeaqVCVVqzfZttsRV5TsYpCi3vhh2U1Bu46Yh1Q
Mhmj7CvaBEfKTu3885P4fUuASgarjLW7wJl0EPiKNFqXNpHXKo7guFrL1HBWc0yi
U5fQOPnsuhKLPJ+lprHvvjvVOtiDB0e+TX1Bh3PbfB6gh/EAElh+vOKUcjkARWgp
b9EHRKkBcpguUamfHbR/00a/KFj4eWPKlpehPMHsCNbBW1RShEuS8lplfxoRrBtO
xAGSAWIG+dnvNjpzYBUYxdB6MxGMLKr8qKajOOaHVT4MY+TQJMqmQPFNXMNAhhYb
IXo7jSmtgmteNISh60jczs6QimYPMH7p5Kge9ciObwxtuni26qCDGnmWks99cs+L
RhVHWpe1X1gS28zJEBTVBLWvlxIFHTW1qugwfCpmmCaxMrIv5NmXWAOXKbcFfK3w
q1qogrEvlj4KYsbWQJGflFb9vMF2FrfQtgastd+Z4jUCrE9QAHdhVFRuEru1rSmW
lxS9HJLaCCT32ReC7mWzDUh+hXWeHo2C85LJMr7NrL41wM8p5yz0tIq8X2upOClm
28N/zB+CqAQaLXDm+AO5KPQqZ7y9lBeIyGp/vRDrlQDMxZ5xqE8QphwA0h9SKAqO
iSz8pRguoF2Iy1mAzJhckMnBTOUQnr+JvmHoeIFiAzR5RBnHr1k0D1Xd8nz8+3vm
7gHroDMF0EhQAcyiHCXIxz3A2FSdSpQSe7HpZln/PDAS9+O6lZxQpEx/PhjXuQny
mVT8GxkjTpNpy6ypoWGl+aayfbns3EWWvL2D8dlav66rOlg0TO04XaA8CJoH/baE
J/TL3pB4ZtEtRC3U/PI9V97ey0PCqSOuRToNsHOq5Pq33vSQghLRuOayMynsxVlZ
Jq3fuZ7ptssIVqVEN8Ke5tU4jFeEcT9ZThCNdDBHLE7K/4ZeuNwC3/eZ15n8pytZ
jPs5Qf/tCl7a5Z0sr3PJHY/81r/CtRNbBKS9pyCfZb9YOzHkR3mfAKvb9A4Pq5go
mEFp0JA/4zvaPbqDdqq9vP3jbKwRYzMPwg9CpdDGEuij0dCEJCOBFRi3wuw+zarI
nQcDnWunto7WP6VMk8XSdy2XlIEG6eFNnOe4M1c9+em17YirDXUEtXT7J9nKEdir
YbBMUZ+C+62VPIh+69vHT9tH7IEaVK4G+YKZXB0WPBB9u/7+f1Z8JjDL5nW8ioXR
rww8F5S8rjgAArw+WY8d6oyxAIhmc86rlWaMGpATjUFEKmFoF28FkOSck4HrTOot
JZNwZp6JZP81MMxSpHgUW/K5qUsvq5g2lU8Ud+QwYGpZP2TTwGXl46jtwuN3aBli
zEK4J+/tPfSnUBVO8uIOJQn+3yTKWu1a99eSE7ogdiGMyWaIbSz27CyKhrwGeJX1
Odw5WJu1Ps0VcjkgKX4HtImQaoBsY+LqOCDRfDSlpCLV1O1OGBT3OV1el2psOrx8
QuwUPt/JHLW13RZLxz8iKXZuYfmqovJdm0MR/qoYn3SYBzq37GNTmiJ3bqP/wwV2
1wlzB5uWBzoSztdIMa8Kv0eO96IHlGlO+Yk2vkmgLKm6BUgxivKmr9AMoAhvdFq+
QXe8JnIjG0t6UuPWfP6aL9h0XiFo6kD+oBOPgwKqMcABewnZpNvwKZVZHV60NMGk
ksuCWn6JS6RkCzBy+IVouI6JV20WMSFrQFIM1SUzRqqEh/xEJIQEfU58q5UPlYBI
w38+k4uwoiA/uQT3NKLZRHy5tV7CGb9RKIR+X5Pa+4a/1bACmttcu4ZqO7ppU10g
u1UVt9vDEMHNCXVjS2ajxYutuACWaKPaXUU3xQQ+iVo4UJFnZhKJ95sD/hSkx4oJ
uCAirL8q+OU3Cg+k/cZmJVLN+0Ni7u7up6yA3uzQ40tL2Ony9NCxeHkNETlhPDVy
Sf82HzlY1frQyn8U3/V2Et8E0Va1GDmlx4+8x77J/hyZG1c/2KX4SWJNPWPPJmbd
DEveo1Pz+xjexEgvNQweIC76pLKgKfRf1XYyd4a2SaQMYWgbElezI+R3UOm757SP
V+GYt2rV/3DqDXr3nnPhFPXJdJSy1MXfiM7QRL4j+1L1o57iQtzzVH3OJB7AgtlE
xUzUrse90WW6s+BmPLHjQM5oJVbO96A/a3ff2PGk9TIEvSmHFFi9D54Qy+mWwHLJ
MwRRWaBCxDNhW7/VnzN7dk18dujtfHhI8iFctobW1CneAm4R9YAkus+lHDW1V7w2
hPUpPn2nFvj31itKJl2zb9jRr/fgjwgvr1DcvcrE6QCDsTqY/kfv1AKHQszg5OsG
PInr7zmjaEEwLZ36jvGtjqsu4Jj09m5CRG9xMq8pzskrz3dK54gGw2NrDdtb3yzA
chX9pCZ+7GQ/VHdHt6x62X1hmFth4YnxV+N3WMEpKWEjcKWI643zmBuGDREBFJHf
87Bof+fCmv5bwJ1Z9CYqSk9eLAWudeuJVG+JylkqaZUcxyO4sbgzIV6reYEamYAD
7yqLxYL5BmkA4kT5uxwv3BdcfsCwTyN0y2INb6qCAjfGaCQBc6Y6WUKv3dGdUa+0
NPL8J0Ztxfa1hiLTiPx/V5k9W7MCRiDLDLrS7TA2GbYf+ETieRPuZhuNXuT6wQpW
aDdAPxzQ+2/RdZCbXUv3hJ6OUfoBitvGrB5kt9cJj8wASsssz65DW4JIaRL83wEQ
D6JrmOs9ozohtIvg7zdALOS5Nf0ITOetyoH+6xTFZb0SH35VOv2jroDlSZ809iRb
6OSe29ZUr4JZ9PWEqQqBY9vTKdb5Fgeb+FUxvp8YpALE415ce3YKnAweCDGlpLu7
85iMXsejJ358A18dWpOBNFywfg0mUTajXUxyeLtl4L3L4iT0ToxkmrvdPIBv+yP2
aTnOs2C+rRxGddSPL9vIMFrcfbhiqS1Xv51q2a4NaIsQcf4Ro9zcy5yZUoWQG7yD
RTJCI7Odzwl4VoIiyn5VQHIJXZYNC2pcMQ5mCdH7dpal25Pq5tOa41Ebw0XXn3zT
dBn1ELuuQ9OLXwmzWWPFvf6Lt0vSb33oYVNOmJAHHQAlhxA/cwCIBumcKGeuOjL/
CQA+5IW8F+p7Mr3dvESCBcq2ikgAHiDaTw9k8liSqTMrIxgjbLd+wlv/ILUchQlj
QkuFbgMMSESQstG178ODVP5/OehoQFMSPSjsVXSAwmbgOI4wMTGNmZSeWMFwAbRW
5dtR8WqyLS1jXo7MdoOzZTCsdvxzjT5SkL0NsI/hmdV+9TcgEbNd4B8aN3hl+0cO
dMwMuKgnuNFepYY1U1/gL9nvhg+8FPKMUXrbOCVQ5FGUjZ04J3C6FuTq70neJcAb
bol/PNgC+e7J5Ys2YePNrvzsu6GdBKdvUx9saVCofNnQBZGnuji/jgTJ9UlH3/Mr
rJkgso57Nqb9QXDSC91sSA7R6DVE/x8l0M3ihEvW32v2yIt6fZgE3nUAYCjuaB6M
S8UjgSbJQiDbQN8bj6cU0CFfw15seaQQHSh6t/DuKNVaYlOOdorrm8aPo8eXwqkL
SuQRNu+Otk9iD1Ynl+IDFOV0qRfT7O3w5hiqG8PmEn/O3cdhFCEV1ClzIX1/8QZ+
2GqRBA+CinvnNCeY7zvIHGo7ILqiL4qjHR7cUDXcuQDDEZs70k5bjrcAShJCmtDH
JznWVR6XxM099hneO7PZe9eTlF7KIKgo/NQsOTd3oO3699w4LsAVhAccg7+8BQcW
iZd2TvSXGn4vVRvREttHDVaIhN0hcQU5jGGOcMZcAQ5anUV7EbUK81zsIKMKqSf+
HbLaugEbT2+4vJZqRqmR+bSoQaAAP+YWXcEdcumwMULjayFiepu8dBVYD7dXYMi9
OylBs8fJKbvPjFOpw6UsoF1+A2oK1ELKADjogp8IDeeaRvVc6mKyq2CtgM5OkQ8C
IoVsjBJMts0i5Xf5rLJtoJeM2UScXwEozwm82ul1XZjQbLxwIP2mEK9fXjVpVKJD
Q2Qo3rvBCRqvcWRvTYhjbAXvYmQXYLXXmj4LOlJNK/qMNQoT9q+jqSBSeXjJLg5S
rXtU+KdMzUMje+b6AkIOmBYOdDfoIR88SkomKKaJ+wQIR9KQg0GTN6u6vamu2NKf
OAN2Zg56mjEu4HNaEwMDyfIcHDA5CtzSgk/MHXTko6+NzP7PyhAUxtidkAgELqD0
oCzfFl6wyHXG1xWF5r7QhDtKDjOGQw9E2umW15f0za3yMX5rOFHiW9Ap+XY9q/5u
8GAmtITi+IyYt5FyJgdh7Vb72eAMppgYeBXJEgL5x/bYgN3HYplcmrEI9ggxBg1V
IcDjWxdmZ4cOOT96TUbMxl1ltOFBlBwI0rGcUa6/O+BRBaKxEbWatbZfgCrywg3C
LAXNalcuWF9rSsFp6TL8bjDmFGe/wuTYTCyy8HUcyGQ/djFY6yEU8lJkBXA+LBvZ
/DT7KgWxYfRptY7FgXeOEnFHfG1ueChq9MTCbLmRw6SROvZYIH++6tx8xRBPflYA
tU0Pd4yskWPDuhiYwNYo5717uaKI64Qg8j8uhgt4/xAbFQTLS3gwJZCYhngSGZMt
Pu4sqqz4rprHwTE6fsvR6HC/AZb6ktE114Ieg0gk6wpvqPK5FXalOMK1YTSvQfXJ
lJXEu9j/n0BuH+tPRZHCvzLy3uJ7Sn2SUNz2NYgnPlI+8Squu1jfoJ5IAe2ZrgyA
D2fCoDmZTNc7wH/a4vziWcs3Gu1qTfMttAyzOEITaUhgNiWSwJ01LxtcEGEGeQP7
yOGumHh0o7GLMJv/VyvRiq8+ihLPq/rkni7wZEmdyMbUD7X7Y4yPFrARNKugBUZa
LRaf5rH98VCfoXzMkdZlEXEZtlCuty1rOtQWhsUg1iPSYT5P4fa/DUcs4r2h3RN3
EJsdOOTTkSgGXmD1U0pvNYyS072DwCqAY1hLEBmLEiGEyIQr7LankWeWcB//CWWk
lAMPqh6W5hTC1nd73jaSeNijnIuORAZeUERxPqW0Zf3aivr9s0UmdiB2FcHMMdzb
+LKnPEDO35NfMkeMbReli4dX+CCSBWiGp8nVEnWiXsHmGA6wSzVqDsXUuYfFrEuc
EY8swY1wLLbM2jrELHlsAa+QSYpxvqgl8Gmux5so4UFyYqrtkiV5jr33xPZVtfIg
HMjlkh6wy6sBAvGqqh4b7rxzaQVOAXsnk8lHgTHBU3yN4aJzuQA+1Suvd76Xa+W0
+Q2QDCRi8DilnzZmtg5SQv9ewxPF6w0N8r16nQGsZF3Jb78rVaRSgyS+RFGW1Wnr
SZ0ghap0D2CRJD2ZhKlNfvJTxNijpIiM+rztrLvXCHT58KJNQLVa0LMFE//ONBdK
4SeikNMbOQpd8VXYG02gqa1AjjO+g6eGSD6jOLvv7moPPxwr0TtvOYCTnfaOUtCu
D0Q/QkbrWbx+w8SlT6oAdxLdgedeUDY4943hUpc9jQQ6gi0NfrGyUgAyd+u90sVN
rTR/qZvljWCjiqr48oizjioEF92/Jcp22u1ryqhGp1OS08+G1G/dWuhCzCYX8PlW
fCeAEder+fbSOI9i4964lLX/m8LKvSP8CtjVWGb5DujYkLV13xMfeipvIqJoknYW
7kz1+dokW8kl7aOlmlSG95EBaRCy9+6HvNCFFfjKJiPkm4yhVGCDbh8t6xPe/7cP
ke9z86V8hcZc7P+cdlRQU5d3c4IlCT7U66dOwrQ30sbMHYsE8asL/x9qdgj8+HB0
tOZL7owycZifMhcokuW/FlH3eSHu7BietYLO0JsjusG3l+kmu/REY2s4HXH63AFb
WQpONLDU8+C0qa4GT1qCTZ7WzFGRBLRbPeL4RFlM3A3aTrPbBwACImafQ9qDjde7
zwlZh72I12b9IN/qTlNZjY7lDIZmZjS0meZDTEGcDy0yXGBnkgMHoZyiLvI+qZQC
eB1oWUYY6tI8GCfm/Zdsk4eDXJBK5WYIbmVcT8w7waxpR5gSHL5/0RxBUHd/RzsM
Tt9jrvYpofNAMMx1TbXvs84yl/M40OX9A9MRxN6vn7cPYIQnHNr3O7SBd7mxghB+
hK6427aAr/fES0VLL5CCUuI5N+WT7HdNcyhfCTsBN/XADaFdqgtRxpgGWM/+zLku
bjOxwnPgzjabFbUUYliJu7LDR0T1FIZkAmqFSFeRWOVVlNyauQaHl5VSDXrlu51m
1ws9l6XG30peGUapyGXiP46aBzEHlT25YPpCowVqkfxGHS7+lTo+8YmzRKjh81v2
MVVQ3kjcBi0I4TcVDpHTe7Rpl5KjMJp02uSHrNLQ7Rs8cKHOqoLaJ2be2+xIyxGn
MbuPauh9U+YtxweqT6KDsTNFcHjxOWF7IP5QRQeMK3+yoz3OQ2dcS2QRQKAbunZs
/2EfE/Xis/XDteI0iZW3zaeqTWY/qnjyAI7y/KUbLLlAriVmAtkruIpq8zp7AlxI
3OWqhbcSyhTGZGtZn48jfS4ZJo7ODiilLBxE1yTaNT7ZQnU+GtqoQslL1A6ZTGvr
N7+94YtOvs9pxn7c4U1OhFnrha9FXaN5Z8IVvGbRCAPz77mmqfs6PhtbbxIUURp6
nCyjDqwdjyqtnzILW6StGKOHhFqYmxvQKhJovI7qadCW4gZiuKBvAXbRLeCZS3Xo
vJe0lBDipssf0SQy9NnP+v11MAJGs+AYHaNLoYr3ypj4Q5sB/vVCCLD3Ppt3i/Uj
x5PWs88ZAORQgxJTBrOQEUJAg0eMd0Rl+/R33PYTjnAhVMuhjCulbe9RXiiscNtf
I7BY4Kywkg2GhqNDtfirMWd7uTLLxIGdD6WndSnu/+5X+mE4Q2AztvoLfAjIqeHL
VGipll4/XndYcWDVHz2msW7xM2HCdhge8dW8NGlScoAP0TrU/15/ilOdZnDlo19G
3ngaeHSNJgs4PkOJtHenXbIRBctXjn/qnLVGiOSd6U8Ulug5EZdYG6xxPTxPQAyn
8aeKwln/kyB2CEuTMqcnXVZccKPuc7Ks6yyCKx7P9nkmUN6WvAgqXEAPR9UUK7Ok
SOtFyZNoaIMRTX2/oJHBa681eFxQOj5vRbBv1hCxqN/YwOOlwwKl9Xz7oSkN3rPN
pcrDSmuy+bCtwvzWriH0VaB3X6TWFz0lcfV5lUOCSTRBx3c5Vc8oLlRV2V0FtfJH
apYe6yWu6Ax0lRCpuy30GzDr3mvd3tux+3l+EronwXg6RIb25XQPatsf2uPVUaDz
V20lEujyIE7rtnkM/6E2k19Q7O7kgyo0KZkIDIKhvDElLSrdM2agncTORFrs1dta
ssISnQEdHZCsN6wtWs+aEGYpGvBg1uUAmiTd0XBeI7X5AmrBjD25MJ5VkTYT5yz4
o/ADuD9k2zaF+DnD5BfAVUUCA+zUcSiJVQGeTp4U0bm9vMWZe1vkGn44GjN8VHqm
rtBcfXQnCCwWlFaqQM2b0Syu4aZDWCLk0ilKsb0lW2ymLtCHR+0DxPNLIAMLjPKK
A96UOsBWxGsTWTe17NiwBeQa7vVrTG+KlCHI7pjqcgSeKvJWDqJttHvO9z9xqPB2
EkUjb+SlKp3HRoTmu9/dv6QEV8Fq6u2/b0+y4uW6sCkSY0ksVk5Q/F8kvDy8BFZz
GIkGcaM7JUeDnRtS5mRAsZ4VHKxawhqueauZHsGoIVMkvx3LY7mVzK9pPSTjaQ1n
ITKeB52oOPGFAzsc3ApCW4tpYr0Yfk00/R8iATGuSNtr3mL932O75BaGLxi5tJaN
Tgz8v/B1XuORS2rFUSeGi9PfE/hk+XIMepQydwS1EtrlGe3BYW0dPfqqBA2ifhbk
5e1CChtAZUCYE3J/mrLplg3nBc4uqx5+pJZ0TRDVGrYZIBKquxcEiNrXR5PDN2qc
tV0smBuMDDrFy9rFi5KQBpOA6BAsQeNqBHtKiZzX31Pa0mFISI+/stsI+06En0jJ
xOTX9EKWcxq/yFB8HkHB+7mcoi8sbyxs5YythBJlkpu0SHZXAqR6wr96t2o7/7RB
JZ10Fht1v5Snx26VkcrUM3QSB40jQod0HVEF/eaA2jvYb1/TqfD8XxXqbn191Dds
iLD0vN4SmJb2yDhVDCFG1h/qhyKIcEV5bq/6oHqXQe9Cm4wCseqp9AaftMMKeWia
T1Qvsra4mBAT7DFTtPo0xldT7f0Pj5l52FdaJDjirtdzyliOLMz6asVoeO4wcUQP
W4PGWuWrsytmr4A7c/LKManuNDF0Vh6QkqZnVnh28y1l6zHpxrqQwaJs2proylYl
p5mw4Y9bEnfuUcypNG3PQvrYGaBz2Wn8/HD4AJnycKKVo1lYaPvPcSdzXEKRtBaX
Or4/sEUVHECTbCfQo4WhMs7Ig5pFsOut2/run0RZbo1HpfAK93/g4OBXZwN5Wz6d
i58oPp5rDwTor6LIgdtOQVp/hLl4Gi5t77I4UF8NhGXjcJ7II1VqaeakqUiUyWwm
ZjMlubw6FMobPu2H+ArrBnXJCl/2jV8jzz5wJvaxjEpy398HNjwP/1XWz86BjorQ
o1scbDkQApwUI3AUdNqsVLtCw3Ybpx4JX9m4KijhpltFJQkP9HK3+4g0fdqx19ht
G37r25Zby1jCQBZx0HChFB5uJEwW+rTabr67Ww25SE0IAVeGqJvMonEusVYYnIHi
rhffU2BoL3tQePd+K0akBxlymVCH+u6+rXwl2DscRORNUhILhq/m1CZkRr27U6Aa
IoWpYi9lJCXiPO/gcC8RM9kGs/D5hXoDGvcGieqbfXzLjNy194Pa0Ec3OINt20Fc
5ZhQQlx3ZU0Ir5iqogZln11gruWUhmk/n5ll2FxNgyZNGFUnUKEi8s9yFNDLNd5q
FVWZd9WLnAJmpberWOse2w==
`protect END_PROTECTED
