`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Z1AqoG5fGgX2W2vLDALliobNDxnbTrbWOxJZ+LH7foVCjqPx3zgCY2p3A2atFwak
l/kV0r9kjLAhF1kmQUc9v218YK3JeHBu+thNDKe8hRVT11wOBsrvAVmI66I51Fez
aOEMpBZ/O9dwuhh4joUGMeZs613Xb6fGompCrybYmiV4HSJdv9HUTmJd8W60BrCu
bjHzjj0vK5IaRcf75llYqxUNZTDH90PE2fOx4L1toI6f7O8FD+GyRjqvLUzdYKGb
cUN1W4jVkqbl89KxyOzp8o0epRHW0GThtmugzJWKlmgdfjrNnGwmIg0hi3xTvnvB
zZIt3GpXyD13uxtX99q85zwPprXVkrr5zjEXonxohkz1VvEwal6nuGVjhFaXtvct
ol49gmyv/1CN335TDnA/C+UTCFNXTY1wJZPdsqArsg5sKrFWUTYR5S4AGkhBNCkA
D8qqaFAkfFQVvLg5GAn90VPILTzV7wD3RKZUeF26/VbKmHZ0aOwXhEkK4CvqJVI5
vjEmAA+FY/w6ETLsKzHCQqErLJFXft17CQLfXPM94QUHeMSm20OqmSgcozC/A+6+
Td+JzTo69rHVK/xoxj0/dtHudnFxxC0cAwSuxKwrQDBCavXGVW6J2o23fbEonXmK
JxXn9lqDQdULoDrBjR0zrOBsyFGN+wVbmQQvFPOJ7i1v08feHRW5QiWTRQGKG4hm
wnltHE9yG5D0YzWcOuQKOxy+xWqrHDFMvl+lS1jm5ZZjCLw7fK4lm6FICCA3GWFC
QKZV0EFduHvCpGBWwFTZDBemOWi6rezLCVPCJi50S9s=
`protect END_PROTECTED
