`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGEh5CLCZdSq6qvDP6ipbu2UsfXMuCv4ecH8l1N1k43q
R1bqfOtK1I8qSztZYCXY9lQBOFJyU/kOFHmCyMZCFkK7c/6UbjRQZBsaGdMbhKiH
3DXv82jj/BvHI/sWy+lfh86QJszqcP5fHAvxolnmKG2obUFzW4FEfMkVeS3QV7Ul
YzvJ6l5bnt59kh+AJtykywo1UttDZ+C19FVtpGNKSOc4E3OxK0s5kfsKf95rRTax
UTH+5GzmY44riXPn2ZkS9RDLcpKC4Nur7sBg9Oq7AFrEvKm7tRnp4Kj/3LaGVGwZ
xIvvsN6YafSVwJqd8vqg+g==
`protect END_PROTECTED
