`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN12Lpm/4a3bMfpwXRyS5oYcZXMNsIGiIa+BnYPalbwxb
7VBcwciM+CkdWMjm8/LibFWwD0AjrIYtMt1Ul5J10QIquO3u/wbNxBkUztTTLYek
nOBmfA210cw7wEYa+X8fj0fICVRmJVfmY3rwto1sI5Q1AacipNSBClZ/wZtqYWtE
q1OnpxjBaPqNyh35BM/V51wJeV6VLnfkB406AAmkSobh6k3bjInNQ19EfYEo+Zhe
`protect END_PROTECTED
