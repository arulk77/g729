`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aVTP3SEYDYemsscXnFS7rsjrvYov5tk67VNFKJDuecsH
O0I2HM0XE5jxxZt7jWaKt2knmsG+gdnrRksnQ8Z7olIOTeszPDqDsGRH9VeRT/42
yDPNfUciiYg3NHrMqJltmRGUPgpb/A3UQviRRCX3lBcOIc+HWKFRui92ukSjPghT
j4/t+pnoqeANCAzzM5wdOIT8z1woQ7PWhNqwtAMVdVQ/WMH1xvVcZB1G1zsZ+KU5
QrdXM/kRzc4S6qQAtvC+2Ctvj9cjaq0eumREZ34q3TWUVpsEATwqHTKl4fjPYcxo
FIhDJDCaFzx3IJ4R8rl01/A2gemyVky2ryDdGWQ94LBoV7F2aHBnYOWS6KSN1lIx
gtfmjsvG3x3ONNjDfJ52jebO0Yfw7pCJMINv98t/NUklpx1aB9exhqfIh0IegjhY
KKf6xKjstzl8V1GZ2XdEofjXapTZINgHN6EbXv5GLIAsl/moYE/3pcw4vPQ5OTOX
rOlQ5QmfT+/2eKHwPbAGWgQPn+pGFPpVRGbNtBa9MxrKO4iTXAy5Dpo+muWT2tj2
Mzg9geACg545lQD+XRopUK2J8wsrNTfG7q0W8OMO5Yxe5ewwKuZDD1lnM/a3cbZb
edZ/CoKe67RkAIm3FxcyRjm0bNxzXyktgD5ofUtP8j03U7ypV4zwsbOtM9V5CWvV
RkD5n5v5RmJxdt/nXgDnpcmg+RZdRLlGyWrj8DVQYLBEiAs4gmk0vzoLsS9C3fur
9PLtHzInyxtPj3swipSEDUAROb48JxJc0Ds4Ey88Sdl6ZzhnOtiOOQzdefbut4um
hWSwqKanYCdSA1bMjKYV/NF+TX1QX5c5HgIo8EMLYJ62PcjhrRQ/pd8auXSmoy/T
rLKNgXpmyGOD5fAdl+ldvMyGAMs9qAazfHEJVoBzMPL91eZuqc73Hj2N8YEV24hZ
gl5209/T/oP89hYgYxFCbkDt3qFn+gim4cIHORczpM3UJmKUedr2R62JHxtaPNKR
TGcuuJnASkbkIP7+4RffCNFYE4+85C2f9qme1OIkZijFlMGkQ0fm8gpVE6GKMRSj
Q3vcfhAOsAqBy2geARpSJwnbGi6iaxH9zF1K7otzm3ehJ0ucW01FF7B3Uv7l7r36
udfFZ5NWlvTKbBJ1hbUq4kMzxTW/4xTSuzEtyBFd8q5UsDC3ibPkGNZLA0Ryg/Ey
zKwPs88O9b/22diu1KCBaJ9e3GsmU0j4tF/xOfdBY7C5ed6/Fqsb7sewfa5P9lU/
N7vXH5cvua/dVm6QhlEstEyYxUc1Xm+AusW7AyjY4ob8Dzn8QwEz8hqury7gze1J
o+2yU0ngMDcoigj2NZ8sPSwf4kN9nrW77e6fL9XPXTQEqrbm5vdi9KWpc0/09Wqm
5k7mGHIlstZvTZZHw4zxVaDHJiPZ9bE4xWWDOlS9fBMXqvLBxFmUfMKz5ViRtYZr
iw6vNuXzmZmY8Pls6e02WlC0Nc9QmVY6xzAu0DyO5TLvnUpSByzORb6sZn2tF/+C
RRPccdT4rr+dCO/k/XN1EIXBrw9yxJ3ZITAtpxgm8IwpbkZ8+Jk2mcRMLCXEo1jW
39K4OD7NoDYZZPef7OP5JWZSFJUAxevw1URRRxjsO7A/g2AwZw3isVQ/SLEvGYx2
ZZtfC8cHhm8hGnB+WtNGYP+s6nwHDWbei2FWMQJDt2WPZcSxJmDMD0Yby7hfrIME
qF9l2UZqCCXtTKneyoZ1OdhKNMiyvfQzv59FsNzVD5vW504FfXsiCZRAcX1jeNsq
zeIhCwyHC3sMLoNtmonUKNTgt7pabgELoaTkKhaQhnZfPq7pNO5a4fOpSk0Bzini
mhXAJKQDtIXYLhlAzBFMBOX1YGpGrJFD4JfEoErpnAjB6PTWavlrGXuLV0bt8cWq
ETIOv54rSyEuSY4evTfgahEvDfMId/uB+/IIPzlc+LzJ0LmxVzge5CBzysl4zFtb
mTR9sSjP/YS0sh1OYoI0ES5ejnrertTW/OSAQLm9LRLjQHzXSZmQLCZ6hkOqAdWJ
f5VLbFJSuFsReUTUTaW7/BDcdQkEGkPfIisWC6EQSsa5+gvlV/VufR6M6rViwF1L
EqkrNLVM9XWK14gbf5zlwzPKpVRGfRaTl3pL2RIsKRMq7eabeA8XZy463/mA+g/z
+2/JSlUSNqIc/zyysD2rHZ7pApbvnDJRXPEImfA2cKI4e/hbpH12RVmW62z/j9NL
EFn1GOyf5S5RLiPKzS+0TQ4sldAQ2+pbWYO/QS5zcIfvtPlXVwUigkzU9v+B3gL/
7Q7GlN97wDX8VvngYva8yt5FYi6pn2k9r/Sbob/1aN63TnzduVlCHDvPtysPLn0p
39oULJTPkn6e2SWE6RX/eHgMcLHP5OIy1SwCjbs+tDOZDjpNBM59C+cnB5s4yelk
6e1YH575TtNjKoj9edhE2nt3AbIDVeaS6XLAENxDN4ja9Ki+L+Hc731w3rm7/3HK
1E9W4ZhE1oJ44Tf2OtRtvxz5Hazc2L2Ppaf5xfvA+Edrz+oxurKPFqk6dzkO1v4u
xmsheXriy54XILD34ywTkhFYF7jmN9n28pn1jSLOZTU/afRr9t0d1Fufplv2t+Cq
Gpmm9yWdtaw4P5Wzf0PRtlNjIuUQlGIStm/Jr9yfCKZYKMud55wsdry8qGcwktj+
69sqSL6vaAmlb40im3mTbBIn+w5bsfiFjhcbgtxkGJlbfcNSX9gzL61wKtEoZ11R
Bnd5ploeG/cOI6G7x18ZvKH+aRyhXdGeHoSF1ZVoghSutNoqI1dn2ajUyHZ0vTsT
NK9lSYNv6K/2kledLukrJ1JVKcN2WKSuV4vo+UGy0c/iHPo+QOjBYOCEN8GWd3Vu
CS+NdxLm4876wrDSIW25QUmazrs+rd4YqFC/dPTFEcL0Roxi0Rhmfbbs2803nmjs
/8NvRH9NiyTeRt5d+PfqsqXAXBpqIIdsQRfFneI2IKaSpFfSnf3QJU4bLrLqQCOw
wbVWwX/we9ZLzSl9ypKWAvA4UVsIopshHk4O3xWDCTNlk9hB4AaKMTlnbf3lBf5m
8bBAAC0iXpr4hE/WbTG/iEN17OcWdvS/ljWHyHUhRQ3pGKHlfJFTFbhsvgFz6pD/
RY3OcVIwoRPcNAzYEjDe1iwnmxJCykKH9IUScLN+suoFsfe/hq3EgIhDrgPVcHar
AckPucXWAjB0WhOzug3qTFiNCHT3X1WUzxH7r3vOJN7B7ki0KK6PluGkmqTKPzU3
v0Hjg2cj1cVPiTqZFeSMv9yuc4Had8kLBw+RTPUjmCBx9zEL1lmhRwglJ7A+ARoa
kTES3QEb7tSiMbPJq0HyquUDVH+oLGOoGQHENTzSCF1mLERDqTc+uK5fPquWw3rE
3vI7gaNpV7vHGFwWSUia6Rq9wQiQGrV5rJqFEgaq3rdUsDrW2i7mbTEgTVd867DP
XucfG57sSuo2VRIjzMaBhiGKq+a16/lxTsBIFRPh65xLQ0/QJR++ry8AC3vXsNuq
ZA7iiMgnJTj+vXG7iESNgFIxOZDA373rCv195BdTlcWc3UunTpGP7x1i2VqEmWhv
eLUXZHXZ2TI3oYs4KJki2KvKczq3YW5ZIEluMZ7zn2S9NamZa+sbUqZ+0V9iMvPu
fDO8qWj4lhfR2JlLNZfzoF43dQo6xPwM4nb7VQLNBxUEtiscqbcj8z3Ew0tKa199
uP3JMoptRnT5tf2WLbAMjv8P4ll/iiyzmdR2oegN4RZ+EvgUx0LUDgV5qp2EsazI
XIrLZQ5hYDAmvR6CBQ8Vsj/EFEy3xP8clJtISjCCz5LsYUAaiUp70sSIQDUac5md
Z064SwriwgjblIXLGrzze+FkdkQgoGkB7+0dkfVSYsF/6YcQJ+1w8TykmpHa9j5Q
+gaVkOa3V0oH2dC1DE/LZQQBWv9CQsCya3ERXlawIPuiDMKCyqoiNY8ah/wEBDlN
2nvYEWEps21Lztv/0CA2Oy15Yh/i8mAUCX5DJWslprU1aiWhasKVZPhdP2Ow+wWT
20PiN0F6gNVU+G3yL74G7xGDanQ+HV92jNGTFD5hKSl5dAl1I6K3rWwKkIAU4Ob6
7JMW8Fq9UrLM8OTgAC3pdVDPwn1QjO+nHfZjf056TlHHbEioaLximIQx6ckkvOjb
7pYS+DVMViQTTQ3G1Ls49rBOlS+RLambxZ+2+16ulqFvZ7gNveDXmqR0EqCxQ3AA
/rWkgfQ5c2IKsJtIXB80nDkBYMGxgPORcuOrkbcuL2+bme86IjkIk0NjFLp1hyb/
w7yZ1Us0TbWjwyOsytP2BBw19rVaJy1Re2sRdspblAF9NGQr20Q6ssHYOyDGZ7I/
dNuCXfx+1GCDBAJRcuqJqE0w2XVajDT5UFNyfNhlYyYSy/oaWvqQNQE3rmJ9NNK2
Rr0GTXFFd0tO1k79E2BEAu/7EeGM94m8KbRxbnxSshrXQCcZzX2Xl1y8va8uqPSE
Pj4Y4QINN9OIfwFf8XGac/fXIh8rFjY0SYIWpJ4ypRItJzj2hLm3SP5fm/2c70CC
cLMywuD+pyyQTXiFLoCgTCZji0Vqwz1S7sV8WB9lHELXXuhqOm8srKyjou87MCb0
YRQ8C8HDclGhBMyOE7++eGKV5fv/EknXaMeVmi1qJohv5EOqzqQsM3PP1dgJmRXi
nPWAeSokPdWxkGQEWlrkFtPuXL0py9/yJiSgnDMDGu2P4B2gY1K1A54bWJ2LFVLo
ihlm9gLYEKVvRxJYwklqtg6GhqoNLVEuX2e87uhMcm9HdQds8KyZhq29mOTkT36K
uew6blVfMknsPSkecxBJmh+R8bT1Y/jnbs8MTA3IoLS+kAAgcbFEdthHTRRpukrJ
8SESVAPnh9XYDmaChGwJnbBQbv4/ynWebjclF+EFp2Ca4KMlHIthGpqbJvPyrDkB
ROo993yVC5c7//cBxQHsdwo/ei+Rg1ragIx6N3dFL1a+sWgftqrY6iM7q2anJ+pV
lz4uir79UkxfigZT24aYXE/Lswl5NDYbcjA+MZBpiEu3FKb2psHrGuHR1sQtm2I/
+9uvKFdbus3jF1StRK8FaY2zkvH0y1sbY81B+Qd/8r7N9pVuxrA2mjk+J6BGeFZ+
AhnRYCmFvzZR7Y7rC46Se8imI5dpEEv0rFigicdjsjQbLUuEdGkKY4QlnmPgYziD
s88ZgzZXWzY57Pm7piXBj32C7/IkdH5BNFP5ztqXDgqqc8N5cWnJvdADySu3f8RY
dwG0P7gEF+jG2SkEHubRVgylNbux49vMVKHemi6m6Dd9vqPE9fRFiTG57UDtC7ss
23Bna9+TeFhT6SHdC/QZl7ORmKgQTJ2S5iOhSCdfCSc=
`protect END_PROTECTED
