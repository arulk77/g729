`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN3N8GovPyqNy94+cAhcYyJgqXDh6gaXvFFcbk1IaBboT
1YaZ+kHQ4hFIcJXOsv9hX7rpmwW9f+fQB1ZI5VSWZWKvJzkrRamfbNuWgza7YzG3
2dYu8qojP7AlMvQ045GF82iKpYSpbe0fxWWJMGIXSdCwCFqvane3tmfww83lG8xg
TptD56YXMEeYSf1JKyMyycsCL0HrmBuRMHEA0I1gBp17EovP7sas7WoSnHmiSk+M
uWGahJ8+YQrsbMAB1pSOnbW86RnoS5xOhChS+7t70uZx8V+KqgaoNO0BFH5oQSdj
7T9WV/0+a7pNlrKh2tRgTSeglBqc+waDhD7R3+wIPRmdYcKMyI6VpgKToyNfnhUh
54Uttm3GgKRmetH1ni4qeMmOCKUpcs0LQviZPJR1U3FH+43MktwUQQwPDOltusDD
iPrw08NyMM8KRkhN6Tn8xWf44JUI8l56J8ByozDyghon6gmjdwwQSLyxucCprveF
VfBn/fwmwfUo29NybLQojHWWM7Lh5EFBNnfzu3jXb7+HleJG/BAx3HYQz5aCzbeL
Z4IawFXCHliTuB5lSpxSps0jniQ98bleTVukEPICzv05zASrO0HPLuG4LHAYXkTM
2XnOmhuRdlSMiHvfKMCUbfvC7y3H/wqZ/dwmT0SwQszvln9qoyIFb66C9RRGyjNb
SccWhUHiUGNoNPaDAZzPWkyGOnR9RH4xtqlh3FMXNfa/PedIqeqQs3g/S53gpOOg
Yviz9/LsvXw/qLIPfDn8YMTDFIrkV4xwF2nXmuu7FCXaNyO35AkQ8Jy0Fk+y4hCH
sA7wTMoohx90PuhbD+PKQgJAWmAMDlDoyXcBCN3Tf/o5MAkhGBi3OqI7s5QcgBc4
5g+1fAYyZ0AFpGB1JHChfzUcjwcbfWXkuqvHGUA7PulehZYLILJ2tK1MUZxSFZir
SZx6bYbCxEptsZxbyqpEtAbnFbvsBu3TrhNuWI+gBGvjk6jwBi0nZ6l42DD1GR+E
nRaPI4oHaJEtEZvZMppljV+WGX/c3dhQRN8fjMxKHok/cqReM2Zhy4klVTNB3WtZ
fkSjdJUX6o75MgAZx3/gPzdOOlY+Gof2AuUxQu0N/EfyafGJFKsLX6XhNQsTwF3h
6TQde6QZyEl9gI5L8wKwgC72iSw3CsyJ37iUFz9ts3OOorHd47DaVKklhAXZoymi
GgRh5d2QUhjdLCMHcXjpFy4+dThuLN261aI/AcGD4m/yDacFqPbgw3e/UPnNvzfa
DF23E8rD11cvFe8dPRdtxHeblJ3tRLYl/toBWrt5Vs1szQQ9HNi2ZqvIIk1Ozntm
tPZxHWyPysTtGtWPghsw2pwDUCgkFsdqBN7cLGBMLUI4q1sVpyI/fUbTKy0JU7QO
M856anHqn1hy0Q0f2GvLTW8UhTr6pS/GjAkRDAoFvYR7bPj8SvFky2UbnU5BFfim
ExHHmelEuHufHS1j72tkjH0XXnziozX83v2tBZOy34K9lcRAveMQzzHMlFvjV3/w
/MXJjhDRfgDhSPKPge8HQXy0xaW01VxJCMlN4CvRDcLWmcKciJ1oCpwIryzlv9V3
YNg7CtgKxqoS/0h35cTsx/2BBQguSUAf5zdF6q1j9uc=
`protect END_PROTECTED
