`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
7bW5cGBP4dxRig5YuqL/ipux+afM1Qo8IJOn4Zz0G0upfpdAj+Ws2ji3z5nljCi2
6EMGB0M85WSwdjFYUdtxoAZenLFDowxv+vOaiaA2xDLpMDx8L+yC5Ddk1ROPaekC
Bsycf812oNcXf/y7VaLcVOJNGo09vQPbmo1kYMqhVqFjGtwocbPONGZvUye/qbso
jY+cYr/xrtFts/EvA6NZdWcurGo82QG9scytBo/DNb6bAq+/sW+sLsgVC6sJ/Bn6
OyTAl6Je4FxlEKh/QdrJIah/dFyM3ZbLgflh4aED4BGTdDHNdiDXgBrIEt/peX9o
qylrEvRFsC7x4WNJzRrB6Kod6nHClLN+/kUm0eItBjoSCYVWVz/JFMcnt0qp61bP
ov9GEpUC7U/45hCjivj4hsCOE81lkkGu45LNLIZEorb33PCeVJGnnuplpmudMiQS
GIAL/E1AnhtMajTrcaVX6YkhYB6WIqkEYIZfBVngMjKNFy3LvXcwJ0eN+TuNHmMn
NnZMEUAZbatxIhvdUebLaxDOjK4euQvrs+kQwx1vw/TJB/9T+PXEK7cPNBF0o2N1
3fA4NJfkKEGdxDFRehLQuxWNA84oLyJgx2bpzHZR6cE8YGytqtIEilGX5u5aT3ey
He0LctwKSb2OglKdprHuQ6Wte306Yi4vOTEbxzw9aRFttia27a2+IG8ZX8FyuYxD
hDfOTlrrqlmPDxUzYeMnFteL5shlP8+HPI1pE13JYqSZ7t0wkbHauyGmSInKCECz
sllyfkYfWAxoDbHA3aHMaCT5xscv3eQKIRgAwGOoW6WzISels+T615EF3q6P7hJZ
IebA8dRTE6BVC1Sq7wFJVumCUoMc1JKxtalh5xB99BLmM6C+8mPACfZB4+WzO32c
DcRj0IdkhJeKwz2fjS1gHclTAwFmeaa1+4HCXh8l19AQXWEYHsMRJzPVI7NYWJxH
429nXDm2zJ2lMvzgA/AtWg7U+XjBOcP0iZcHxtD2EFuHUKuqoZyQk3BlFv5TxZYT
XJRzwS7XzRQKpG1aB32MUHPOHdVhDcemK3R9WOCmEPoTu2uwHJWhMYjsxgC1r37F
il8jXuHvcXh4jrLIOE7c2s4xvPVLHeKkwmuMvHIEN8QRwFGU5OjvHgQQtR01QWey
thmsrh+Lp4FDxP5zkTA385lBBm9ivVkakmR2Uk6b7QEn1o43pH5b8DRkmPsq0PW7
JFOuxtlHeezXpf5RxpCgOld2mgKQ4k4W9v412CZ3yUCWoTlZdloMGyYB7NA5cQQU
Od6C2A1clwmH0li8ZQb78Grn3kbI/cDHwKg4fezouJ2UbQqbiJa8qpxTpfbzasQF
FFafrLu5Cn5oTTOiECFarJjTPsUfa/XCwQE6z+sAFlET5SMJJvEI2zstoYOgTxPW
bNB7QG+MA6WYgG98R2Z8rehXJ2kUBwcfpcdUjfWXy0KdZ9fwcYmpCXiz3ZQjrCBV
hwxZRlGv/ugnoCj94pj/td5XUAOA0KREp429pOwNmxZaERciGQ7zXIJtpmNLgnAa
RsBce8mXwFQmY/ZSrtuim27yRdV0TmGHDAMVecQ/C3yh0OB9FzYsJcpAw5lGVbxZ
AYqEs3Bhqrdr0aCERpCyR+a/EepDfRj1wamh4Hoh6N0CIxvril0viwSnI/3I0Vq/
DHF0Bhomd7Nl+mfaroukg7qItSluESTF5nvxC/feg6ENFDUCYQZRktdodjryAhSO
Hm0BaquJuye6RDDJV6Z5zIZsIJc7N9SvDAXbHDp9n0ffc1oZhElIBGOWJoX4eC64
AX440aNsTmZrDcAUl35opub7cHtxsQvmwrdK5BKKX7/xfpb5pPu7f7O5dPe5fOo8
cnKE0pkCsUctQhd/hhOP0wp3NWeV35qjXk0kXll/kZZ4a5MA0Ujj1xALesxHpN+I
mGkL6nT5Ty0Cs88LazrN2ssFxBpFa8mbIG7JVUpXqtYPOKM/G6N3dWzZNz4/5dBH
K9koP2A0WoUAbyih30fo4IoLi5cVHu/qBmDE3WJrBXPOVd3ZU8Ya1M8kIDPB3068
eoI6be7YVGdmc5puFYhEDMSboBk1fakgpviVEGHbloY5yob1VzXwoYv+dGRIsWE5
2ooqxB0WmjnJCWw21KOfvMS4V1qDK3OlwRJRcNVC6ikS7m+3QVWbr6EYJlYVpwHT
KUJy4BkRWhARGrxWBJ11YMJ38AAcfb+cbWNNi1h2Ghgkl7KnkRMHS61YbqAz32rR
6HPnyspNy0/ISMFH4yuwIj9RTDN8XZe8QuM1ZRWU04xON1C6SfCyfN2N2ofjxBEs
ElKvhbr5TcJ5ywr78X1XGiu525hit/HzHA5a7DrNm4xLNx2AKkjk6z/6tcsKCYyu
/TSjNhFlFCjMA6H6w4FGCiy0XdnBHmkVthb9XLqR91gxEHuzuXcCuljThGdZLKlY
bC/SBUKfY8QAzxLuL9iWh5YxcYwUgvcI/0N/4VQ92UUM5+0Xwo+ljfuF40PFr2sw
IUd74/VWhHSm4v+jJ61MgKL53KSlitPNaHlltpuJFeY=
`protect END_PROTECTED
