`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JS6Ee/OUguv3S0KjECptSJIj7CYNZHY8kcEf4UxLaem+8g1BYEUQimhPp8EISumL
LRqt6m5lJrZ8yif08jGRgR0KRJCcx1eiH6Apw690SyCg2WID+50Zs3oPhlEQHeie
YFOpJfDOOnzZi/whHecudeU24V/dizlz5XQPMJb/Y7RbkdmA88pe0sZ69yPSzpud
shTG9v4XxOGClNOzu2wVKek4Gb4mW5Z9m9D6F7sRlNjpCWPAQA1xJGKARqhXrrsh
SP1Twqz75A2co7yb3S42ZBLNfKUOvyy2Sf8BxSAKmNKR7rOQ6YCa6cItDZgNmO5h
srqntDUwZSVncXTACkGChfmU3wuuNPq++oS5QlaHPVcmYp3qsyA7kOMujaYsx/KX
fzsJ0GaXzKLh9kZ95Dog6qfHEJwb2s74yxvY6y401/M=
`protect END_PROTECTED
