`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40+HA1OlDyreHiPJP7D6M5JILAXZl8wYg9ugdVniCEbr
UMux4BVeWzLOdpJA9Mdvb55/Hov5sIfNxqeCGbs9I+TvCkubM6gR4znLcJ683XxV
X5r+gzqqcOsL/aDkaxnw/VzR9YmKk4OC8WjDy4FFdfb5WVuKupYwJl2wq8MrZOS+
ULTux4y3SDY/zikEsAm+Qf+zfMjQfG91z6uIyDFtAun+jPKvRhlqyD+uxB/C+9vJ
zLqEcSJKImdiA1p0SJQNzMOkf3/4TnO42YfQ0Tozf+M=
`protect END_PROTECTED
