`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePRP1O6mtBJw3ciDqdrTTlqONjsaIuo/rTVulEQnTauc
k7BkJOLKt8sm75pqaJrx5rAIndE1Os9ZtfIze/B5vR1YcJuL77yUV6SLtkaBL+2j
iKTiKlg2Ot32V51P7E3PNErJCwFUi74VlMPgv0V+bWFgbJgCilW0nZIDnrQuNW0l
rTgyM87E2YA3uKARVhOz2CniTQumW/cWGkReZFky+Rg0OdfT+NTrzo1mn5WxbnBr
tyonTpUPbO8x1f4CVn9xdUO4lKfjMTLh+tl2GNO6+PJIDFP7ZyTdCHAWGPAwQZkT
QeRaHQS4EOSLh3KP2TH3cNcEUzdR3qRRWxWT5u/5iCsTqkNKq926tnmCTyaZo1T5
+qG0U7617sHBagJC3p6mEa0XDSDZMPXEY0TJ3n6GRJcy/tq9gDpHP3uEmKDtfYd5
TN6mstgW9CW+DLG1wGM4WB0O/kPU3Bmak/kH9yuhCeQjGZ9l2MWhx92R1PSzJP/S
gKtAT/IRePVv1SmbKkkCID6EKmGVVKO7nJxAGE6OvTGOEUQuOThTiockk+AP7hFU
AStJS+71i3TODUIf9NvcdMSVAFmod49a5lwWXwNgQMqPvMD2oVdquKrZENcd6KT6
yvr6BH6tWPWZKBMOXg/Fo/TlFkTCYyXN9aWEmp8nXDYCNKoOduX5faFYcPz1vVwC
W56RLyQzR1ePNCC5DlpeVN90EQXwSBYkU9YLOqpU6h2AyoGDTIgGS8dUvBqUa6LZ
eyJXlGxl9fcbxxvusE1STUf3z86wi203D17INjk98ZRtJ6BbifnaDMsHCO6nBy1z
JNPWcBlc9e/XBzyf6TULR9n+ec0PG5ATtCd9EVmrvxOJFH3+bD7qtDnKvQvvRH+V
oT2MsjTHQhn+08Kyvc2P8keOBLr2BtudG+0lwTX8pDGeW9yFg06Q4iF2W+CkAw68
WL2grNhJC6hHRkQLUw1M7Q==
`protect END_PROTECTED
