`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFu+TbZTr9KGRMakUS7ZlasmGGo7vNlrFaXwpGBZ9C4V
tN1gVHXeW50zygLUfMnGlaJXpWDyTRIMygcVCBle4aPJFdigFGw+iHKK9wT8IU5Q
4I5X2sMQS7IBcvf9EBx1esd/qYzYHe/dziLS52O9nQPkntD7bXQE2VYc1WY+dpmL
GSXNwDJBcqoBqHT9deAGraq2f+m7pmW4uEuSOSKs+BFT7B7zmYcJrcgLoR4j0n+Z
0TFAYKcfIts/fWZnmx5jGzDlkLcjg/NMb+xkmQXYyDJeTLUjlJr/CQflFQQOFe+t
KaaHB4MDKLlakPXlOUwnmGrCrSetdbk4KKS19c/WiRf72XUbweq/MlfjmT9X05Eo
Cu2H2ZsRriZ7hxl+oO6RBDPLRIK9snXJL4lS8vor3O29JuzwYhNLFA2BVLByqBDm
hoIy/xmbddui16r0vrfWyLuhghmHEWTw6XJtyL6UAysssXC1ehErzMHpeTbcWuPV
7SwKip40GmjVhFCM71mRSl7Fw7sIkt1FsIL2xWDa7f4WAw+pgrzPb0vdd5TKKjrH
`protect END_PROTECTED
