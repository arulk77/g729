`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
F8S+AbaZCtWk0whsAcolA5W3djoDnel2qf8tOD5QXDq9r7Gcg/BljE7GPqU1Lj6Z
g3Jc4nKIsvj7rOxMcvu8tLUXX+pR5qysbGyMpiwF2/+ClxaFSwn6/Gz6icTb+wNg
fS+vJnCXjczcAfe1s1bzz2SnxmHBps7f6S5/buCoDlcVrXeia4kNNaEroqpnkAY2
XuOSqvItfKAqwYqmHukC59tjkUJ+zZ4KohqZHjhZAlIHnjGnMRc9dZIDyIJ7estb
QIgXP98cV3pl2O0sF0Kmz9mKO09I0UARxCyMyvfpQL4GJ5EeJI5scaban2CJAD9O
qH75i7sDHA1auocglENsBlNYw7fjfAYoydovYLsVxMTctcxxl3SbhF0s1hb8iHNz
zsK5kgnwewejWzTi05PDmPdcl+DxUYllm2IHWS0VHHrolkBKJkrDU/5XVkyFoKC7
2GaLGgji7xod2TFEev2VK7as71php6e9z6mWYDyWvR0=
`protect END_PROTECTED
