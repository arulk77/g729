`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOfZfMPJfI4IepA0boIhdJr8x1KZJRulfgPBTaLusDva
fZmf1uJKp3CapcUWu9W/8B2pJMYHEXqJ4SN1XnK9/MgVVxJRcE3YlbSpu+dFJktP
rc3ROgnfsr+p4NqowvG1iIM+VAtRrvLEZ6l/4usAuo85z+9IgEFZ7FWd2W4xqGca
tJ+asBtuZ3cWVIrNB9zIkRL8MxdsI8/nBQu/HMzSdR/IG9QUmNyoo1RvT9b/4OsF
`protect END_PROTECTED
