`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF6HxgoO2qppe2FKO26suJJ/8jkieqmf6DiTpHt7yEIG
50r3TwTZ9mYeGZOKeeBgZCvzAqi7MlZa1/dv7/InAGZs+XkLE51qQQSVGTgIKgSx
lfawt00Qda9WeOh3i5atU+RAkDNCNRlbiW7gOEy/a3ETVMo/2l9MUCRSoeqZ38IH
0owCYXXhhXpoGBhfbEY3h8JC4VfgjQTKxF6PMqYjE55goX2wbUPgKJ97dO3cDtYA
IRAALgv48pDD93SwHNcKfwMTvqLLOA2I4ye8H/6Qcdk4ivVRqfNjGshKQLpnw2VF
BsO8IXqKdBqfYpgOUdBZTLvzf9/6Br6nZ+y9ncXth9C4cZi+3oucKtsIu9I2rJPk
5ZFFNrEgUOVYCvlXqcHiVkCKtXsEMFtpt7K+OniezjB2qq2kbz0jBGy1fyILtW0X
o/3ME9h8uKazMFXyHmvP3hxhO/39k1MPcgYvz0wk9usf7NqYla1bh4VAETykkhER
SOGEUO2AXrRH6yrkRaf0OFHedRXrxWb1lpIsn0n/MJYyCG9gGkMQhHTmpV2i5CbR
`protect END_PROTECTED
