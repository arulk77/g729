`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBpnKnDvuxDKOyQFJ38VxDfGDJ2HID8uNsOd9kDh2vc6
0OoWSmvF8Rq45viTyLScPiTimJK8wuJ9lOTuAeYUNdohKf1hv3f+6QJ196w6OBsD
b00DsIlaoWfHJkBviFLeaVPH3EzpcVUfsqr1JQA9L/Krqd8pslqpNimxAPzLMiUq
pDs3X4YM5hDkI8TBUic018yl8zR8BPT3HTdte7Yv2gvAhYZbUzq/Lsifj06wA8jf
LaX2D4y3Y+RfkJ/32QT3rGEFSb7IH9zhRtweMHpwOA/Zxdtjx/WzOza8BY75y0wn
4r44wX3hSOfq8K/0j5GwQ0PmjimM8klFOwp8oqV/kkkE8dCBuMwjdNdrLfbxTD+K
zysh/1XCIGQqv1kIx9uyGhGXNgAO4SnceiQXuskj7J7qXAQVSyPf0Pzc2nc14kZ5
zJBaQTSnKNdtSYPfPRYTOfcVgbT86TWP/9cfZSuO8xiBzGM5CHNJbEMZP8OG2Pqg
LtlJ3Mt4+oa/gb0z3IOhqimS6W9XhUb7/TtSmeNGyBZd77flIm4JCqPzl5DqtkB3
ysNaDmoK04Y6M/nEh/5E94yCeQpgEN6iNMfW7NMM/AIPcUltT07Egf42+96nOfqa
AWwgO51KZgXZIwIPTukqM45Rtr5bKstrL3FpaONJF6WJMb/PUL0w5Hx8/RiGp2m2
nXeURl9I+AggLXfB0k7bmcIIyFH7R923IM1m2T5U9q5lTVwhQPpnwtFDeZ1xkvcn
3rj+/PAB9k/SZjDsEl2fG7KW3RGANQ3z9FfjnIAVMYy3gzWvx7AucrQh2cqj3SE+
p1mtVMacNNfhBrNuW9tdKlcqcBlAJKhYlwM/2ywgPgQ=
`protect END_PROTECTED
