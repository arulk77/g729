`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SUpo6xCdlQMUgK+32v0MkC8yXst/6810Pcntl0oTbfvc
YdHTDYpkmA8+Pvgr/2Ov0HIsKzcLrerTaat231rgn4kSPZL1pFUGH5XY+2afnDZ+
GBmuQwHBxQ6FO70NolM/touREWOhIqyZEVlMuDN28BiHNTdF4jGLtDC7ksgMaBrB
eSW0XY/92zVRYS2GH3F9C4fyS9/rBseP/lUjJp6EGNMk3jcaFeep5AURi9XVSNsd
cmm0Hb3AYhsH8j469Ub/01kdTsmOMzj0GVY2OtC7BMku7EhbON/JuFOXCC/VoqNv
4GK1sfBWYDP7j5vPTiH5YB4QlTZNjUgO1a+1tTYzBBwlRohNpEmnCVKtP1wR0rzm
IIgbwCJlE7q2Fxe4h5NVy6vpAJSmZ9ItIl8/T2K6UwNduG7LQk8LHQyCIe2NpWcd
hUEajl1SSXI7C54WER2nCQq/94BitbRZkoYaK6eiY9256zgHIt69RmjxPk6pzu5k
hVnOPK8bBymsftFjUHECnBizOdUeT9AyLJF3x1zC3dRfBa4mLW5L7uNoXa42KSfH
lVwfDsdBw3u+hbnWO271LLYKS6jC/So7EDQsPtH5zDoF+fkBn5yAJOXewHmwECdl
tETpztTdRkY1mOaRgZLL6XsFtWrTUb8KzRvo6O+5dFVjxvt1jfHqbCbhGvX7H/Yz
wNlO/mk0BsVeYO8ih5+g5fIDxt0yGASIm7KaJ2GDfr0FOKWkZFkzqw3rV+5wzcG4
/HPwENc2J8d7YQWaaIlnjTs9dyKRWzCEaxJxMBfWVISjK14fIcaLLDJ8Id5qmCNJ
rucuAaxsbK278SjdA+5vIBc39CYCejVaTBK0gyittLzB4LNmrWleOYibPLnm3eix
9JhoHYmPvfVjuhC2a8rWAY/owfHx9Rz5j0r4X89IEM2Qt2KAgim8XuCvI4GEpT4X
KGtxSt7xgAukmTQXiMXs7DDSJUWuBGJ0GvDsVlIEJyvKtal6HaeJ3oPZ6C0L6peL
hGpPbjLYqZR6fExpX9KdWHLJ73lsIRBXnm+UQ0o5B2fGlGQwWXvotp1wBqu4NfAJ
yNArXykn22QJTIROwuHnCoOO7knmJ9RvsTARsh1Hz8Q/ZgErX5TVNOlxgl8ZFIwT
4DodzQCR6XO6RPZmDrMAj6twem9oqgjjQYN+D8YY+qLNx25d+XWgW6XzbMOsWJW0
rw/HCL1SNQ7mV9DGTdMo0W1sV3CGzXdeCBGAzSsZZgmmH3iEgH/4qeHFjhwHXqbM
VffNzLEoljFY5DEQWJ/r2qaVyB/yCQlp9r5jisszEXlwj3GIBKLgMnzHiGt+JWOU
EbK0LCx/BTzJYGxj2dXbAjUauDwmeNMOo2TV348YeucZ9h6KaxtD/xuzscmr+XiZ
W3OCMk2mHv2DhsPM5uJ9HZMofrS+9l4YvgpfnllzbR6ehowV0e9zHHiMq0/YclCo
aZ87GpypFTXeBMjl1I314lPBnlGa4BYKKOlxgHO0AZJPjkv6/2FxQbsdI/GWbP+Y
4Wb+LSfbEYV2ushyxbrm6jEqD6YQhEq52dA46GqIsZ6vWbCD9W3caowGOrPjKh9B
QDJA3YZLtJ+HU0Q4Nf0sg4VkmU9XuP5330a790l7FNCh1E6siSSyxUfp43OF0wgK
Wr3PRqFcwPUh3kfp1pWe+KZm+rSRmDZt+TIxjvMzj541vHSD0DVwz6nDRClpM9H3
z1fBLEqu9J7WCdHkTEOiFwwXQCpTwJ/SAAYRWbLCSgIdZBZqSymwAgBArFb6S/Kp
k5Y53HaXQf0uvRzGgGHIpwgxitwZEh5GPFIT0h3zjlm/RZGQJaHK0mnBu8A0yXjI
us2EUEfE57LdpL330QLjGcT0NwxfwKfu+E8xWONXdo9rNOI6Q0Gk05flPZXrjatD
aDx/NRcy6dkX3QSviTN41w9KHgkRxiHo2vT+XU+wJKUd/+3aaq86B9iQOHf41F6i
gnk+x2Uej+sMFNovcWNEXaU/8iFssL8kWZEjrve6iSFn7g5/iw7nuLNllbXUb3Qu
1/aFoOsFpEc60aGC2MYsyO7IH04zQdlXFBeDvb9jOZUZgvd0IzORxmamu4n1OIHh
DGRLmVWUdTIgcohDBQZU1Usv+TbA+8nt+gKeWOZPrUqTCcSaSceninORjbkZwc4b
8i9fOZPlJwzp6qNjzDn812r7t7nbYc8vAlagfLEzfE3Km5l67dYGzmFlQYzAViTT
2lPKjBKIDRAtA2+Cx9lia3GXKMh66GOmQHeTrNRAvCVj+MhRz0cPzWIU5W81eegC
jHWQF+Bcsa/0p/mI1dUBHhIk0BwRPppjFasy+g5lhhtU7HguJkxQB+kRglL0/nys
LZ5WUs6h1qwZyrq5ey14Ww2veLtjqdr3fDJuPGLRo7+/TElzN6wer+2yzKe7sZNq
`protect END_PROTECTED
