`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48SDBqnzMm5RU0V0eOuN7IWmwi3RuAa18Q5RlC/FLb7w
mFEyKSYdxhdPw4DYKyl4RymOtNH+Z3FUub/cZ52n4w1MiFaqKOjIahEWhCeyYr/E
xmJNQnDIRkhLjH5m4GtXEhbDfafQCVXQtZe+oTeylw6mOTovLnnX4QMVK4rMQpXd
fz0CshCQADAWz8uTEMP3aw9fZQlHYVlaBgruVIobj/du9yubL7nMROF34axmRtE4
Im0yvbJg/4CarR8DdWNPMN5GMXEZlnTf6FQQhZKm3S32X9AzVBj/VWr6IFGkesHP
B4w+xWVKJ4faBHIhMxm/+w==
`protect END_PROTECTED
