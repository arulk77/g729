`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG/VOFwmZYnR1CecC4GQ50/arGr46UJF/Owt9jckDb87
YS0p9S5ZZFY1OnxvtVPlGzJMucvl4kYgp+eG5y8DoRmyLQCVT98gRmgaBfLa8Fdp
rDtnP0buFAY9bh7RGulwXl08ZEG4vb1a+LIq9MlWQLoeWjmOwEUWIAY1E8vSscUt
qU8EyL2W2MWZxkFu0oGzx9e/5Cu570fCDS/+Xi9tTUfYp6Tr9hLxNqDFW1jMw/L/
yiukyQ8whtX5SzpZDjNPQ7/ETWwOEDqZ8VN08xMDvc6q5a2pi/AGKPdQgw/+JtDO
vOPa6EZS3FWtWPpyXBT67WRnoIvfMwA6rwwTUjINIG9Mkyu8GPTpn7RbJoBICMbK
+mREav8ST1VVkACeVX6lQiZTAwrdX0NJS2b/cdlwiGdg+13G6xRhgxbFeSTOz2aV
bu3tB+WfEerR55D2QAZmeYC4vv2WHDL2/nXbYuxcD75Nnq18RSNkqgLOSbcIroTs
`protect END_PROTECTED
