`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3cIP9E1nepUubGBK9azHi+gOibH6QDZDA65qNn4qwOKjhlyoLQyHnIftT7FjAwR2
NMnkvHIrdss0aceQAcKDW0X7fgloroN+ygOfXJjK4LPgzAWqp2Wl51qup0MV0gtF
ozx2iIThpwbaYvznZsohstmfnAgE+VwCC/4GnrQZMt52+bqCHDKX/Q/udJAS5QTj
qNcC0R5vHkW58oI/JlOH+LnbW6GIMI/b/fLu86FVt9JoFPVncfikeWhvKbtWmiNd
DZY9Dg7crlxsHZl5u9RrApZ7Y6bMZwx87ag0viMJ0IvrRA2EPPP8uH35ufsLC7/G
qy7b2tiYM+V3RHJ2kHDq0KCdoW6w2qwiEYRbeRrHxlcJdGnwPsqIa79yavpKAd/Y
O+Hd57pcBC1QjchXR9bECrF2mB2GCuIcvfIo8rOTrErOVlWNaQbo8lTg8Wgl49E9
z1hB4NHQcU+bf2PlKMcqwOzIMIHUbCC3JueTnZz7TgSU9gkB5nSnUy52qntMbaJf
C2MmYkstJNDb5QO/z4DghYQ+qE6cSBitngzDj9q4I5F5q7krgMHAr/7SH5V7ndRv
KndV9y7hIdaoZGX4uhzeSrBTX7MOjxI9i20i6SJRnL69oflOq1C7/q3u6Z1BgiTW
x+14D1Qa5QkLMoVPYavudEYfQTK4ZNu8FCX1XZQSGPVoChsczg3bT7KKxDDIUhbP
AMfAHzyDEJiYFyK3OGJm+bYI0eWwl67aW+TTrE2pQN6/cjSq+CpN5SLiS2jvIc7c
qCFa3RjPLbwbI6rAApwKQVjabmqlVrDkRChjjnoNXjSjolaxcB75tbx2jypvKQJE
uG6NQPjteTGkepfuJOL6CLSRP0O8zWJmm4iB/YANPv/qNVMUT967tCjRjzes2EEx
bA9hXNFGvkyCsDeuDQjFpBwjjYctitGUEXyuYTtZQ1m6pkdRf+nw1EZB3oFcmIfz
+PUzpjql0cKr9NDTRWEVRRjkNqMj0MWFR5NaeKiszR417jbkHxaIpXmQcHvGfxZn
mtm4XWCA8x3OkmuIdOqyjmxSdRAhf1pmXbWUSmhmZDbsuATsvw0NDBOx4uw52Atz
IxU5RfZB2N35O85fJUK2wsuR2/X5H4wkqfkfXu9J1FiKeOyObMe0gNALfqeD57Am
I0Dyy8HU4FacNpdvBvi9vyvVkO4U7rmugAHhFx3+NPht5Iwn6/gP3sN/8ROk5OXh
eY+A62enluVzAsWPuP0GvTXcJiz3NR9pVvob5IBg17EzL0OjlTOuzdYZmZcEfCLo
LZMvZvxkXxB0Xi+jjqxkbiDlHRofJ0scw36DB8LLE5W9ix0gGGKcd575CS/PxhT8
iPC6fBufdUcFzcL8gesQHg2kwr1wALui5zMP4IDLWqpc6RxYeXsDDGi/6DTVEM9t
K8cFKmQyIs/ODre1j4K3FwWBmz1oEMcXr4UBJGb6x9v8HZE8Ajw/OrnglsrtK5tD
STkePh95AEj5da5ZbunYdTvINPLk2r2VNSATLvnPTqXu+EViNPX+dZPjwAXU5WUx
cn9WwWv2mpwZwlevynQWVdYoiR7ge7zcfwTuAevH06bfp3TBNFogx3Le+StDFNuf
TIofFesj/TUkg93vjqrxiSWZF8VsumkNNsCyhv+lJrEoCeQZDtC7xIlIQUAKLj1L
eEZk+Zsc0OxEPKV46zMSyQV1mR9Pr98vc43WYblomVumAY+mgRtdMfaGhg/XFhQ3
YUjClqZLLLPckLIB8IMIDaoJcxOBL+TthGGSvjyXgndDNfrHAJsRiVa9S7x/MRY1
2UwnX+uT88jYC0QbXj7s3l6vITuP0zce9NBRggLnQM/Jl7BGVUsFcrT3ZBTw3NkK
qfQ4vNt41CljCesMbQvfcI+g5/bCQOt4LBwBDrrj1HiTvpWm902zrpZf7rGmCUg7
sVBbUvszY3YwOKhy7S/W2DkBuV7ceVvCF1AOH+KpEZP7Gb75yKHfSzPSMxRVl38m
QQMabW1uCi+WT2HlvyP2rtnLhRomINkIufoC6y8RXvC1j8soR3Jwf7Bi9aWyo+Gz
16nI8p8Fr59/6Fp3nDkHmimhyV+2C8bI/6kn+27OJ8cdBEGhUqxUzOQFgzmfYm0+
QocamqRUHAyUS/7pCVeZ73fciXuzf1oLgeV1dmxvYETSQHpnYmYJGyUKNEqhZUW4
miQP8BkSsGk586WXkOwIFffmd4dSYNxQkUIVXc7WqsJF2D+R3QEfdxdJuR3OwKmO
8hgL70yKbgqUUI5ctgdHWRo8zR3fXxzrHT2VB5v/JoIeU0WV3SfEDNJfpY9FNOUa
uF71kvD86Y+sEn3TsI35OWEdYEhOj8GPkOMu8StspVpSbZRrgv+WBSVLe3N436E6
bTyKW2drbuzfe7mXGds9vIhxFthaGr0G8G9k0lIrHkM8LK6hITnF+euW0oNk/Sys
OiaZbOxXCeJG1QFvQuAkMyUgNieozFFMc0XWngq4HZ0H60dc/9cEVVrk5vcZLZL2
tIzO4tD988asEr2327ltOi5XyH3+c0wCILIYz9SR3ztvmL2MdPXKbbGgmUU5eawi
YpF8D9cGeGpBWVt2rmxUfvI/EXUzDrD6GdOvOTwdWvSqJ3Ef8K+clR1W5hzcibJq
SUuS4+JekNUv1uGYekLyIqdTgr7jJuGE9PuYylLPFTjuj78BbYVF6sYTMWKcms5B
EvDm4n4VgXKtFSNXOh+Hy/+ndTfxAlO2hgkzRNK1OQ2F8EoH66/h34digZm1AP3n
zG1NUyJQj5UXU1A5OUT1QhMMCTC1HwJrKfXmKpBU34GsK/f/ERjUTOWd5cSXAtTS
3pnzZYEVg576XyLp8OSDTGhJwqerKZWroNxwXNHeX2kI9KSYOSpuRCg/eIblvECU
UJ3zYDlIah65KXPK/vdS3iIrPrzHccBH46vl1xJXZaNm+7xAhU5U03JWpFAT7OTS
KuNAepv1U8b9Zihh5VMLpVJQ1prRU81Rf5IvA/6ARq6d901eADY7QHEwABpbHPfZ
SIILhpmZfpE/RB5+VEb7Z5kq5SD6Lr6w+koQw8Z2qK81Ua5ZjO9PalbaQybT8UPm
d93hf+kCvp9tM+s9IyD5eopdeLMG6sBxrYvYQHDwWgvwmu/O2E9blbZP7gLTro0N
0SlWp5bwntlLr6XueuP+SrNS7xAY6XHUKE4oUKCCmF4jpIVpJIGUJwDR4z/gEHIx
iaB6EFEqOcvtQJBh2LLDmKo1ukgmtbgeZocvO/cLneEruP+1FoRqgNoh0orLjlNk
1wqvrMcAv3ek5MAJouKnJrwX4QVxMkeuxYljnB80hki4iOLnrAKPswV3nxsoh9F8
88Yu/bx7jIfB3RJCJiT5GdduzKzwusEWME6GZz4OpoD6Xg12kgdENvkSLn4wh7J4
gdAyrva5GDgBXmWaEphcCXLVpz8unzy8NQFFM/lT0zhJA2BS/gwp9WZWNIsDgTOl
M93YC63REBvVrIQC0rvRh7gVn9TC+dysGLBjZy7B98NvIr0geQQ6tevSZ9+4LTq1
vf4F3u4nLYZw5WrzgKNiziGgF8UeUnoYH6wQiZq/6zA=
`protect END_PROTECTED
