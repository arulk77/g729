`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJm+BuNyir9YBcXFbenwxAhYJY/dt8yaaiN4sKULTAPF
Ms9e96UVMXTpbrSitSdordKMW28EWfMKUjjPOhExvL36J+dZIuCm3G7LJwbbTZij
fI/9dxEQ/WpTSIC4LbPUKIy28qUbZMXu3S5LSOXvcGKvr0hvjfFRNzdkmtPPeCbZ
VQ+ZR3qG8jw2ZSsvQ3ksFMpaua9ohr/PJ1hve8rJHLy5VYktPEUVUWUneLQJQnUn
Eg9GO2P4wx10K8FzMz89OlLiaTOPPg98jucNeeKAsQiSjl8K6R7cy3phKUYWwuyx
kunmJM5c2JaVhUmKDAefEdrbiBmex3neCt+ZXv1o/22NH8WHRf6Om/GDaaYU7NGG
YE9USz4aCdUR8tO35eT3cgMm/GLHFsBRmk8U8/PPDtP2efbdgK0TMCQAHmg+Zf/r
k2gSZP+fwKlv6DXyZBJCeJlZFgKoMhE71tkkx1NqRjVDo7C/HF9BrA3nOFy61zHe
Y1t889N0U/f5LcNFBzlPVfO4rp5noOaTkR7RKZkhMi5EkRKjM0Mt0mTFFn5l6bhy
jQLFkgAZ+SX/FvqtbEqpZMelA3Zwh86Of+p9V84wPonY1VMPGVGC3qePRmLGeY7m
`protect END_PROTECTED
