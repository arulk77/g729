`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
sZsoLj8clRS4b/ZwGuGEqjnGX3Yf3E7YHd4uLNkBbAW2JPa5WV7zpaGU+isi4wuX
UUF+YBd16XR+TPwTQsGdZwDG1BATnpJj8nZEsACQyzSSbLwDpLQ13xmAG6T1EfQM
RoePXL9f7w/0Qxp3+FVJ8fdJzFGIIeMP/6/EiymZh4J0ohAi3enjj9jXVSYpKNRG
eCrcNwCz119adK2UeVK/GyVS1HaA3tFipjH8wgYbMBEyZlOUX0udDkeMxCcZADQ3
xmhkF5gid20e/bFSKmw6ppaVHoVktUQ9sHP1zD2wap4=
`protect END_PROTECTED
