`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEe1kq8RtU/Riy7wv/L24gdUzpLhC6MdvNbay3h7vO42
r7XIp9vWS1/gcaoEPpdKU2iTFoyA2uf7BLIJyAzhKP6NRmszMESypOffJCiPvEPS
jU+25GFmtwPl5HHvWZYu4upZstK169qCf3/r1lM9A9GeUts869XKCtUAlb7ebBpt
qbaVLyI9KOL9PmRxH3NZowlCRYd1NdQikmLmRT6IpGTNupMObA6lNz3EfUkYRcIU
xFQZxxyesR7rU+IsqQnXJR3RsMc0wqqiD6W3jy1ZgN32GlAWqjdgnoTOGnrMUfPQ
bRO74C8x0B9dK+5zlaRaHJAr60cG54QrO+xVP3mLC797wayu9/rVTpGWd/nbJCzN
sitc0+deyuhK+4Lzwqob6Br7yghKXBUeachY8AnnCoOYkMCTdpTRZT07Mut460Dl
CNuVZXI86k2cdZHckZGbq29+jFIdDXf4sSFwuy6It4r8jbVxZ0ZtPAxRQZvCxnPy
PnYxIx0da5qkkZYM1mf8CNkczzHzz17fprI0zAYLWxU3ZTEUEd5pxOFt9WYpMkh/
`protect END_PROTECTED
