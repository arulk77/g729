`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHobwqFRLAXnd+QE+GsXe5nCSMrAkPPqna4zrgjhItEw
JLw18j12/3dDGhgeF/T1OVT1ixvrflaStOouFT/tAcqEoUxrvCEZqwv62/eYXi6D
sy6gVkHOe5bWAxS8ZlFKpJKh9cM5P0MbTl2Enl6etgAH3VBdJ3jK9xA3LXO+/rwd
wdNmBCH7EnxcQrB9Eb7IMlKE6RdjuVaV3ndHwZuPjus3flVUKlWOPmBsVe6UIBfD
Kh/7rFW2m6lQgYP8q+6FgSKX1l9Wyt/H1ZleiMsXxw51PwuvChoxygsY6z6tI7cv
otarJGukC0NTBk1AfQD2aZOr93Kbp8yDD1OSR+VBCWfHNLjbEDZpzvfbapN5Y9Sh
p+pYCCKEbQ2tuIunUljHAlUEM9kgDullpfAT17bt4tG2YeQYcsvYHlgq1owT6TRt
4GZX70nK3PBo8CkwAnkctPGDkIqKzwS5SI9t0ti0ro1peaSVbPQXx4N/DF5ghd/T
`protect END_PROTECTED
