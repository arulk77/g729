`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
r9N/jFx+TkSSDj9pOt+UIZ9j1LhyxvATs/Bo8DSoi5BFuixYmC6/ylvQdBDKg+EY
298PKNxqR2PS/6MVYnjP6DkVeAMd14XYyq7L2kJ3bifvk36OYE9dJO7cl5xufF4d
wwsDg9hw+4eHd6hJ4Wy2gU2A3czgRkvvOaD8OPO/9f+RpzRavYE+pU1xtYJxdcFN
LZtl2RCnVakyglumEr+tymfmRTreoNQhazwfpKZr9iJBUHjHOLfvjA2qVpXk3rAq
MsGbTkHspbarhPFxsn9xdqnu4Op8cVB93AuJ1hj4xZJFVvaKWl+OyvyxCXPCqMeG
J5BHyzGewraTjE89wdHiahcEwByLYiFHoug6+VWDHUezGV5j8LLBE3Kr+sBlZHGg
vq/s6hn8UE8+3FDeNWRGueNNVyvSL5rWYMsVop9+QH8=
`protect END_PROTECTED
