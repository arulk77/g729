`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveElhZ+wzc8CKdWZVT4jpklgsefS2eaHSqjX1QJvDMndV
W7xTOk1QFetdTmz59+eDVisbrgX66YMljKQVOrwPMA+sAe4AD6k0KtxDsfDvJLmR
mfymaRN73bLboVK/LfBZNjvA7nYU0fXZLQgg25wCRg02S0zRB306Zm6FYK/2TQSz
O/WkWDTyqL+q/JHl6Ry7fPdY6lezrkb+DCLOSbcJ8wfOeDjIROVFbIW3xtqxe9wx
nFj46o6ZRqxEXLT6wT5m46dagODNlnCtXVOlaH3ps1DsOXQVLjV0GhgNs6X0dUTL
C7z3P+ueXynlIGd4V7YJ94kWmn7WgxEyhfJbR/omlROYVtnzLg5CPjzYCmLwEZuB
3vRs5Il7mTeHOpIbNghF0KifpS1JEhWb32lP6svPQtxhUssIc9X0XCl81BCjuyDA
OBoMHWUyTonNzMfre1FQFF1ZNKIVk2kRmTZLH2hn12HlNcCrp91mzVCmXof1k52F
Zy3WRrk4q+VetbEqnQgq+1NToN538aIp+J/p9udLqWHgsOk25qU5zgx2Gw3rlL2W
`protect END_PROTECTED
