`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAXrGgL3XItWsd0ORruHDe+PyG95VhtN5RncD4NFgzayU
OF/f7VctaZ7tVFm3ZXF1tXTD4szwUBnHFFjc2DiuKpZUKRcNvFJDjPOe66dcCtiT
uaqvIod1pTsshP7dLzmeT8730SzUe3jSkUumXZgGVBvVdJaDMAAIQ3AF4gyQgoG5
saW0zzhvEn1OrPNxwEKHvtRGa1pLdARK1I6iKViG5hbeLGT04gTYXAvvtkS3s5UB
3jhKcwww8UtIWh4Gea1X5A+gJ2evOCSnCIkjVKW5YtTUaqesk808NKfNaUfoSN+0
KbikcYcptiNU7WFkUuOuXPWrZsx7L5K7DQP47iW/p6fUUuwkCnVQUpP81SYPc/HM
o+yzHs52ymTSQ8+AG62XD4H1EhPLYx8Vs2F8a4zqrbZ9xUCIPrMrZTvml34zqegW
++l9vaqiSvNwaLPm1UJTAn/I4C/scYnpkWINYClY8eAxKiEtxkCvg61u7XgjOGUX
9VzhFfoFiQLUEGYAOx/bRR+92SgndVgz7e0JyFzRHYgbU3Dqt4HQn+jKGSxWkdDv
P6VwhE/SQSo3y7u8JjOQair5bsmHUUePkGoqqoZY22J2cNY5oVw4un5hYnwmA8cX
QrpEA12gDalm/kDAZnnMVCoFKXz31XlLW47UE8zGk7rwqBBnta+L76IvynM28wdQ
H2HyQ1/zh2TaQytfNqxJoQ6SK0YwTYDMVuT37rjFdwdnbWtb4S3bVa1e6jZs4x5r
h7n4CwZdxzIT92+36jBS6Ty/hd4zaDqL6mJaFVK7wlioptO8+xZvJnu0uX6Pgu6Q
+SJurlydsSZDo8xecDxZPhsNeJJgw705tb8Z0If/PrBU4IELzuMGLuVdri+osCoj
3HxO6WvmwcOD2wJBLyqDPceSm+MsxvPre6dRok9vghYyvMxhKCsR7nFa0PXCr55h
bv/TWlWFGjkQsZLwSRJKT70w0zKSej9NdysVLK6wl3Ka21NoSBm6g3jUZ+ydpP/D
EnnX/kQ4J9wYSEPXfWKWNXBSntkI6UMOAyyl2GG5CYazfF27HU/mgs4LM+TTAMuu
4gsv6Gju9Gqx46F60NIZFzfg2MWk/U38NImZg8eN4xCcE/8tS9dtm/vGsN+nHgTd
rvPAl6r7uUiuApV9lAHhZlpQe0an5OrG2MhaudiVnApIDjh9DAOkG2Qiv2TtxHkU
8P12IfA1FJ1OvgzFttMRjtYeQ+a7rmhLqauofcPp0OkNskmxD2WSy7rf6lV+dAkh
hW38qYuO17HMGoSIKGOh0X9ho4q3Ff+FgRvm3JJIvAdZmkxHJD29L5UgC/TXGFqu
9+JeMsqAnvTKDSFbtKE7Tr2dqzgxd+YkvZI7oHdyznZGtvLn2eAU8egYCiyN9rou
k0wfrUBAFGijvcSxc3JuH66OsiN06XSc0LP38xjGDMB+t8BrMbUDvdamWByxYEhq
MocG5PnzKNYotIWfHz8azty93oYnd7FySwsqrmDKldvRq9lDeQsI8ZiohrvPPIWk
I197BD5pen5kv5xyIas1l5jg6wiGAJWGrRaL7vutkFkPwz0k5jhAA5D6iiQfWuSp
TDIWpbsiFmcNmrZD8mPYfOmET8jPXXCUQ7l/R9vYOaV7+iu/NU9tOGEHEj6RngE9
Sw3Z9voFk9yvVKOoHbl26hBWsBdjfTrPJ6HT0eUbd59jWrfD4kgiDDRM0GCfEBnN
tsXiwBmP1jK6WLUBN6XlF3mSAx6Fu6GGt+tj12oAdfZKmtXlPPxOHqAAwiRMtRfu
aAG0N126H179+p/wj3Xe66v0oJYVQ8Otq0eEuanq4fe+JsBChDno2mrGkD16JUqy
JKitigzgBmxHKzpe3pAxzdu9iooUZ2/Y8GqUcbCUpE9mP4RjCn85cxOPK/BqktDT
laXAvd0Q3K9+1f69DA9ibjC9AiKagP/NTgzB7ghiOkJRn8gDCtjo85JvMcYkXlMo
jafuMtKYZBgR5eDOZiSYXwvyQbPSSj9Jd/+dbrbAoiRRkHpGYmQli7sicPOMfXDy
RP4sbBmqCY7tNbZNEaFbvJT4wDJW2T8EO/z66DLT1PJ8HP9T5EHnBKf1WamHjosZ
SAk3m5K8/cZMUrCSPvsyCIOxUHUEkiL/g3/AS2y12Z2JvJ6DPOKF/psx8sr8vNMn
XHmkkoI4XEgo+42jeyGSA4jOVYZDgYSVGjNQ9DHViVAThR996p0FBCZRIIbHKuAb
1AQ30Y0XzKVF3Hy0tYK0g7BOfsLnRzFUSwpqJ4UT9xhyS3p8i8UDZSKnJlp8OJ+l
lUNi9IWNJ7xN1WUohDjYRF+DDZbvySsY+zSwTTqUdUCRISl3YHhj3IzdJs1nPBdC
erUr6DaB+/2t47sco7iJhCayXRpNdjM4szIUWDLBqCpF/ZyZwu17BRUA+yh0Jf4O
CvJGf6zPq37f8VrVhsTUIIHtJVfPSfZoVxBg5yzfvFOmsKzqR/jjGxrzcybtpt7Y
VyLVyXOBSdiJxno8YikPQI2FH/ZZogaCGJKslAykizeZ2lgXNOA5g9L7XgA8Ohws
LlYO9Zpv5exrNReFcuCWqp2zxEZ1LNXLBMshjphfZX3/8/vH3m+u+RacanwJmJOT
e0BYLPe/pvFWXdTuRBn6CpEsbs6/ActGBrsAJh0VomusOXgNirG0t3Vg+T22xW/y
PMMu5sx8YMCHv56L9Pub9U0SdO1rIbdSWjgRay7LihnbgtGnxq6hMHMyAd7QWV6A
1ujRuy7OmoRG9S62BQDqXP9N1wQ5eS1UF/v/g8amNI8rCX55zFbQelkCPifugtRJ
V3jWE12xQZ4RToDZG7YeQv/YOOBqYtR+Kd3gpbEt03b1qnpLDsa0gCtl95mAQhaf
N+G6b4pOeWPnp6YuOqrfDTfG6QfDgALesJ3JFpnssZcQ02ZWf3aMrjSOa1Lz8SEm
+wZ44xKZVPFaomW/hv2TzA7DHDHLtIQerP84K85Q8+zxxi8WiqWlQbX+NOB1gcLN
q4SIRIwi3+/v1ZNoc48oL2HiUipqpZBjJcHaw+mPbKKTWY1AII7yGvFn+b5p4I/W
KRIzpIxcTzkapnVADQNpNJ4AfC7DQ5waj9SPcYoRVrnUf5HiH+E2AP/k4QjegLJ8
JKw5qGG3FWfZeIMyvConz+gCO6E1q2oSOjjVbw9HJyKTTYjROrYqQq/tFtxTFbxW
xNgag2gsaL5rf3Ouhq1PvrOPkL37TzH4Z3eQ+YRoZCT9o+MuDaqjtsEm3rnYCyYc
fWI2IxSiI9aW6kdCLFXtgISUIXTXhplKuTYKfdr44IrbOm9krVQJdwXdqhJ1i3m5
aXAj1gX1vKVLy+r7/jGJj2SGRS3CWseCPy3vI87sSHyt4YfnRu/jlxnt5+GwzkQ/
5/StdHqIKcz4OwL5NAceG8nNqzVPEHsprtIgOj81UF4MV0cEiURVBB0F0N2BCqx5
P6DP60r7vjY+6iXG0/Ir8mMPk1a2xCAsI1qzOw4tKuqAEW1SoeLH75fk3ToEV+Nw
SwvjPyU3fUuassBY9U6ObhkUF9XsUgW+Lh2tRduvAWAHPzGjcxGheA1Vvapz/PKv
HY2G39jlndura6UBJqjTcRZipp67LEEcbqbiWvE8E0z8LitENW7XCdP/+o6/nO51
kzKIlpXpPubRVuFvF4X32XO8DiJw6FmDnX3+eb9EetLVBWulOPfchEAh3s2Rgx7u
5y6a89I/WrEtmL7n+wBFOo2kSu/URIzxP46D4ToUOO1ALPSxYyiXrCkirHOAR5L1
9be+TjnXzbAGN87QI4Y/GIIdkCQEhjeUnWJZPRdH7Fz6ciQ85zbWmF6ffFaZ6+QD
I+07GgmU6r01pGiHjzEoUE2fjAq5Bh7i2dEpnV21p8DWn0MfRxmESJBrA3UrsYqC
AX+9vK5aeC//RxPvHYDnITJUpBN6XdZ68kw72Hm9ib7nfg0HXn+KTgv/PG+dTPXN
qgsR5ejpSEcCIw6Iigwn9HN5LsPbhFgW2P3VBiYDziIX6VCUxDQIAM+KfuzqQI8b
ikEMRd6ENQs5LO395I1Y+uivLWoQnbrqtGfXaJFr48OPhKg9C5SYKpgzWcsZDVUQ
krTUsW3GRsw44nTZH53Y2gRz2dkYyT+sHFOlmjA04VeP7Rq4hGKfcocEAbElVB9j
n3GyjQWRoIPe6Ze7NHmhCrZ+iFLXsUaHaDz3AnSgOpg8FusILRsjDFivDGkIUFCd
vfCSMyJRyMSfnNbdfYYJO7YGPpwJjEA05FX2wVTlr1C1eqNJiWTOiSq26HdFUrFp
YYcz4hBAYo6UwFgR37SzEzLwgumVKMm0jWUKlz/RUqetEjzSp00R/txdim7ZEWJ+
9iykO28z88YspanipZTgfl22vmxefZcXNQ8RYztrY3n0OiE9TgGiQk0YinTcA6M0
UEd5Cf14NLgy4XpfkyHuFkQPlg8Y33Z4jl63vmx17nlLdwiBPjHIbU0D92zONBes
pgSXEqd4rBMqTbr7lQ0OAe3++kfykEMXZbt/jnu8M9tDJTvoHHJ2+WLRRlLYa7E1
CHeEyjAGEhH/mVtgbG8Dw9c0G25qZQcLOGadUawYFuTfaHazM7fIq5hvg0XoaNQz
CzqWDaajaA6xfU48lcvhK2YDAGsVLddHgpCoUINZEr4FkvwS4PRJpuY44a4cu2ZA
0og1tSEuv3SHQg9Qk7cP9QAGSvqByZ1ojwhkZYnv9WBaP3/q4nP1k9bMXZxM3gfS
xatzBmf/tvhdEGradNmKwVOvnmpgspb2tAUA9NRt8Tbrw1EE2eNMX9pHIL4ZnZjH
W5AjaSNbGJsd1Q/4OdZU4UcwgUG9tNbqYwvCi9OSXso9ZOm9yzltHqFSkkh6MSgX
zCS900RpXPsdhEKlrIboLhxVgFMHOZ3YKPyfknmsbqrcNd97AravfklhBRY3s11m
NkcJLo9Xy35fSoDlrNSkfAFVSMTzyvDt2CzmISvh6Bq8ZE2cRrcF+r9iAYBnhbpC
BAHJjUKvN6PCeNRk1Cb3JrRr+byONBdfZHrC0Msrojisd0KyDnxcyAMnkzGBiUj/
+P84CyGYq0vzOUYVJHRouYlVwBz6QoJ3oLH4doM1L2kZbZvhiXGeQzxrFlMCHSxU
naWEbgNwc3euZAky2as7opvbDphu4E5oXpTgj27vGZWXyCavlb5vMBtje0fZhKlu
hW9HTLRLqROYI5EBHRi08nC8bHyIZoxX/IQc4UvxeS6HKAmJvwsTkQby5ayKJO5w
ub0nC/iDmaO87VdMesNyTQgdOCbdCVZiv2XIcpKF7UflAq8FjjWgFZqDbZyDDfjI
O2xpnCEovEHBv/DqsD+OWxkKS0GT6nzERNIgmg+U9jKFJiOl2n3p2sKQTUS2kOTL
sOgDtMW7xgVdrdvGZDTaHUlV3SSr3mEbLYS56PKuP6N261SQp3cOERgY9JxJZMWI
9cs2HxP9iKzqavqZ5h7oEtIdaCIHU0v6mcoJuwMCDFrANASE9olPaYNYWoJOe6nx
x2sePpr0GEOweXyfj4itFUgJSIETpwSRvilucSoBtc8J+Bm2wVOwpU4BMWEMtAZ+
nsgn8Lz/zsDo7Fa2oNKe9etNoBCeKDnNTTEXYuInscm4X+VPUMPFw/L9kf1PO2Rp
ASfkm2LANBOAPuxzpj2ecPALN52jLzMYm2Q2LVsXAi3IhSW/BImZaA0PSve8fqYl
4hDqkM3TD6HTrSfrd5tEa5m+Dt4f/dwrMAoiuJRTUgPQseOYWPmaORmnIbFtY0m+
1xRy57yW9SMAVwpxWZ+pA6gwUPiljUqRGoE8HnSgieOnZcOZMToK7Mg/HDojWo16
CX7N1wcjXEoze5MNhxPSGA6JnKUZbbr427OEo2TA/maUrKBhE5rd2R9pP0hJQbD+
x+NgRVP3vToo/OcivstdUVv03/fjolGfaHNf0f/VJtEmh/Gh8edDVM3822tLfkId
XxNw7u/nQujDsmYDWt/7Ow==
`protect END_PROTECTED
