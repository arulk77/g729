`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49+N+iWwP8tRGwXIgPQzS4bjwwvNlGuuRsT02kR+m8Uk
HdMtOfi7DT1CW7IDDbGCSgK6JdoFPZKRN6z0Jp4rpsogFDbst7OyuQxR18VPdCLJ
feHzyR2AlS3uYRW1SekxW+eADbqRRcwgwCTivRffaFQf90h/dS8e8OsCx3fmuAN2
DxPtFtRmI+zddRyEnCUIpT7LVrnSDrH0BtfWsq9cGTE=
`protect END_PROTECTED
