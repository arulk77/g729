`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8Sdcv9CXLSF/cLUlY9zwB0PRjdXxucroHImmv7x1mO+O8
BXisjBJgQp3+Omlewzoem+foAaUqBVzgWZLAf7MOGU4SJArj5stGfR6LHJ7VBelO
9JcVg2Ve58wenRMGI33K4scQ6U4pLMhmGJka2TEAHtw60XKvaV93BeO42M4VVZNQ
XNE8L8YJ3Qn9HqF18fndzJg47R/q4bAOVWoFJ9mVFjyT+Z8XKmj4cXrhsTcnfOIY
htUvtCZRN5SvI9poKDWNY1txkWqQvHnkv9x2net6CmOuJEWoi88VC7JKB7+YzQdF
ZX0VjtwNldYFuqx32i3DY7CzdO1vZI584WHkq9ulaiAHLQwS3NelJXePjOH9RRPn
SPtt5SYHrSOoJNUyTZ1Uj4DuNEHs+OTvwXXGDqHoQmg6yPvw7W4e6+eNa34EHO0f
4bypiXEf5UY6ji73vHojgm+9Q4Bb26DR1VirRUV4R5+71rVRKjFlXKqII6uROEJY
l+Rnb1bgKJgV6KF/RbTVOyRi/w5qQO8s9Y7RIaz8ZTk=
`protect END_PROTECTED
