`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG6n17iw6EcA4zHfJmHZ4lPI8csrOdRi9Z5k2ayw3xsg
c/F9MaS+zEfCWE9oN9+p8mMm88kz7z90o33Nq/TRqFNWJWz/Tfn38EY9EIjRWKJf
UFBhcefh4ucdsSx8y3JFrw4QP0lCNuSniPbLAuWdrpNBZFlosQ9bulEGWfW8v9mD
3y3ybS7bm4rYkg5/UaSZlE+DvWZ/skRoMBoYuSITH2Us4zN+0JsGdq5ensDJw7Go
kjKmSTn5MHNpoaatHQ32v4hUY/p9NYNHb6+IzzMVGXgHfLS3/5nW+kSMJtv6U7xW
aD09DEep9mMgaOZxjBzXxyce9XJX6yfISrfDEIY23tee4WMaXe8PQJBmuzvzKOEW
m3cWRf0QKPvcU04Xj03s5WYUWbpe9oXFf3IQXG4MMKeq4E7ZX4CXsp/w475nB4PP
88cNS8UivvCE2TtzNVg1/tUo4L8lTarcpV0BpvO7Ep257KdQa8sgEt+at+ILFopm
X/pV4XR1bFuWkq0tCqOHhSWtnjn76Mx2+ic4adNKA8yveMStMAZ3JHCN1L/JDpjG
CktxVWuv7jYDML3I8ouKzg==
`protect END_PROTECTED
