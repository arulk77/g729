`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45l7RTAjFX6EEOYaO4S0pF0C+RfOLs+maUPNH/b0jkLl
Czl9Ef1+qlGMEJLjITdtzrhtJYw5JS3LOGWDC60bSIgHWfFKFcbpEHtdImpJMKK3
Vvb/7SgWoliVQGiacpEGvDgxW15fWRDSeiaF/3Spu3zZQZejfogl1pdQEFylSv13
b7Sb0vFyjuTaeDm6QFgvCau+axmX/LQHD6NDO9MSIxkwe8ppQo3fEyn0Sf6z7IsT
nxZaH/7rdEYatkjG67oKrCYxlW+oQoFy9X9wPPvZvfM=
`protect END_PROTECTED
