`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNxrVoI84jVut1qVc68V185NfYBP9GM8wsHRVNoEAYkV
kTGXq6iuz95aM7/XLamPuzpYID26jv+CRso1SwYs62Y4X+DPMdis7yDCYEGu7MEE
NKCDlP+Ggk14e3a7WuD1wMO83vyDhoioumpbYNPLAccfse2HBNrzvg40mEy57QUu
7aHcvCHj4kXogdof/JSSwp0a673wXFF/v6dMdLGOqQhE1XA6XXLksMiygMFEm7+o
d+O0e3pTp5KsabVt5hWp6zVUqtt+QXlHyXvgg2/l3o+7Y2lHp58gNaxcLuvxLJsH
PtUUpck1YdHjCG2yMBbb5qyNZvP1BT3EfHcMbeYRMxdhmEt+LGW04kd8wzqlUuob
2fEMu9QEsdxgJ/lziLY8KIaawy8z77pXRVLWgp8mBZ9ZkJbW65zBSpKG7NtD0tpU
mXJNzzk166YbZnmLZHdXVlZ5WCvuzb9UQIRc17w3flYY8KP6RycO5bSvaL1Kbhd4
FKgZfZMFV1eimwAI3xVcVw4a5T+y/+/ag1txsU0Si6gvYoUiH147fB10uQ21r4sc
W0L5MrH7GwrWiN8UwNjgDTp+ehhOditWrtfnLPvGTSyJcE6X2RRNGEZCnIcsQvXY
+GL4QVNkKrlqlsJ6K96XmGWsK4DwC/LXiJW8NmD+1p74vmbH8YpfcOoUubFc8nCq
QvFPdDyVxMZlbuFmxvS9u27G5vtMsxBYVAuUMaGUj3kDTrVzq0o3ZiCCwBmp72LL
Tuj9SnM6deBplQmwqzu5lsC6B9A77DL/hYSb/Y1CCM/g3+oIRU4vWsnqt/HA3uSU
yb3Bw5SinCmS5V3dofmXZElw9fvkSqOBvx/5vWqf4LYJ/SjvA5W4/IZu4tUD6Ag7
Dcb5ZCt3xmmog6xFVP5n+D387sTcWZGVYjbM2vVJVxbNA16YCqfRX/3HKZcZTBeL
RPJLrUM+K0ahtzLfezaTdUqEuZh+0Y+O0jGxhKqugUgPzuUUcFyEjVHuSRa4QnXq
N1k4GTFUPO0tZuCsgfaX2DU8VeXCFB8HDvPK0TDo0xb9BZlQDxI/cHgoOUzqwvmQ
60CiOOYGy8NLc/ljLqOVcfFHlV0v72EZNy40iU/J02eupjknX593piW8+cv6gAaV
JHJVpQ40mFkXkP7AevGgwgQX1fS2KgNeknesHExUjexWV+joJJGGyqLa2t/72cwd
NjbLP4lEXnwmji3ShPvchwXTgkvWVrOQZIuA1cO5apBFGKO/Ynqv7oG/BIF6j/y7
rsaevJBvgqySFcNmyVJObAF0aRXcm9A1S/wRClxoJ7mYcyaOODg24cD+kfv7qQW/
hOqKUKtZvi+8B5h2r2enS3RwvQd+2a1LVPVCuAFFMUssl6OWdhDaEtmHAV+cgi2z
cdH6p52xl2+saY7pdfwvplUzNe36Z3WWW2CEwn4dNLk2ExOrTi6Ef9h/rQtjQRXB
b+OzZFweu5qkqTp59sbzKAWb3RMdiXyZ7FwbYglkHMo2BQBGlVMK6RNjsIjRum4k
xp8IFGZSOsXYKyoB9UN5w7XGMCM6sp2NzVplsO1ZXYmPgh/viP3fB+JcYof5Wh8A
i8RJfMUa8g4G2HHQhJ4225W0vi06c/Q81A0HVDBxq9hUqlQ2vc01wKegkNM24Ogj
sWDX/f42d2vY+PmGMUhoS6qB9SBy7t5qa651ifKlyTre1cHIT8eu4P9XRmIaWCUq
LgeWkX7jzCoF336jocRykfr52ug+LRDabbAYC3AKq1b4aAvBwgd0i4LgHU6xnpWj
N7Etz+kto8Zt1xUtDg81OwbAhmomM3pPIKu1rDObGq60g79ihpALG2xQ9BmZ6onx
dv+7ssqEXvVdMIeaaW7phP0CkQrOy4DNyWRYIfpu6A16MxCU7gISVkMQz8K2Itrd
0Islz2TjquSifwmaCeFZ4ca5rtRhD4GKm+w3unr1oBHJyHLhxYju0lukvJy2HpjG
Bt/kWjT5bMN1w4J+id5iGsekDKsqBUMtERkDn25z9uOQ3UHa41uzfRLh/BO0qqlQ
8YLUbc2OZdZAW0f0/XMgUU57FlvNCdAeW0if2mFI//b5PW7rwlkRe76zHS0mfyJI
xdO9uzxD91w/pJLHC/34kXFWKrQKAOgD3ricnQxstOgfzd3ixH8cjULyOoMXd9e9
iHvB5rd6Q4ofxtyuflWsk43EdafvpSDFRORlI6hckRf6QZkue1Tt/F7rSbe78v3L
AI9OVK75nWGWnCABQ6Cbp6H3pQzzKkCII3sB9IrmWB+5X5IzVbUSvMki0pE/kIKz
Ksjpm1ZI0VNp1of5sf222a3kNAoTKEUOxeLRB+oKtmS91sbsBodY3u5yWVtFuX90
aW16QC+y04qmj/rpGjoG5eMInBLDBUUlmQwGtMqVMCeuZ8vuN0smhktDmjJYIhPW
zJFNgOIjO2UHNUd5IXP7VKTxLd6xF/XXkgdTCbUQPGGJU7ha4ihyE+M3N7UgwJAa
4VRACMi+mcOF1Rj2vuonKisvAfQb6D1G3L9E8nM3ubhkH1+sRPGuyNw9E6IkStj6
IbPC1GrRh3DCAnfaQ2WJ3KUBaRws5lx7+u1cKQZoHQDqcfRTc1qMSrJ5SYKUPhXb
w1xMey54T6JkZ/lJef2M2DjNZuOXV/N5uXhbaCp/ukO9s/5fqbUQTgjbSzLZdJfQ
Wv1x05bdS9TZbIlfMZhYkewZPGHt+JxtbNp0vPgNdMxmdXHep/S/QgTFG08ndeF6
By9nzyLsSjAkiho7AuV6I6JAZ2+arqzUURemmhm1cHCOTuEEDWqLO6J4BZkOwmvn
F1Ya7Cav618f4jg+Vfhi7B6UiohhN200F0TQ+VQlLMfELDehOJnjA5M5UUGLUPkH
zYDl8EvAEP0trcY7WXS/HYI9vzf2PQM8qSp8PVY1Y1IDOIPxVyB4xFsUYe14dKEI
+n7B6tBcvMYk504eYREUISX/+soBtxih9VGXzB0GKi99tYUz+6QH0FsqG3tpCRv9
38DgvU6KMCa5o7r4nvKBPrd8WlnDrTHFXIoUxHvUOqUwjZOZzkUVgPrLdj7H//Y6
lcZCfODpSPWUeSyquhF5ZtayfexZ8X4mr8g+UY0sckdnXgYIoeFBlvC5mY5bmIiP
UcDffJcnsfegck9KqFMl3jM3n7NU11Hnz9mnh6NRf5WhFg0cBLCPhHah0tRWJtbg
k40TytSonSK5SQQpeMpLtx6yvceY8y3LG6kcSwylHu8DYnLgI1imHV5IK3+h+qn/
3zXu2QllhWaorsSxJ3uEO4WT0/VMD6mNnAT1DHPauNEhK7tRJc5RV3NUsYoohwsa
ygrMcU3PQs0d6hNV5mcLCPe1j4xW5nDICLcux2o+0I18rxpKnGsna+RW7Yip8/VI
XgXw3urLq4WNP6TKR1bYUJs4f6gfjFPuM57dY6DMJl/mOvBNnkA7SfFNpkTWbcJy
dIM4PQqhCfjQl2ZZNemTYoWFcSeziA2lJYvO5ZSTEWZ8COTYoUHNAhnNcuIrno8v
ViTq2x6SQI7mpNs5UDEKk/CwtHP0pRGOzp5nAFf2kE+fzkagmb/SdCUdSSOjyRWN
LdCtMnMUwV3I7354OjP+R0dIk4yw+sqchG1ULcXWuZ83uTu6n3Z6Ih59sYaMM381
cOwiaJbbcAHj4CTsAp1y2xBJ5CSdsQ/E0D/3i0ZzNb9JuYabnd+68Z45QW+Yeyct
DNRuMlqkHs0+eHDZpxoaWs+/2QqmhDXePpwRrLYf+Z7KLso6TaznB7qWr6EZWi5A
Q7E4du1DJihPG/srwz9pEZ62WWN+2apHq5KMKVSJp2F0LrzbHSBSZWEOW/HB4id+
JM2OGoJy17kyrSbVPzDYIhWoWssX/QvnTpMf93fExqVv6jU7lekYjmm7iFSf5Dd6
45tB9Sqv4+Fp32V6A4xtfXqYYSpArbPh12VWHo8ZdDlstKKWDEzAK/n4Jvk+eu/Q
9p3OOyG0TSGMm/pY9P68OfL+anRIRVxC2X6tTErG/I4FSNQk867Bm+Sp49Wxb0JE
o0nWT3TlGSD0+tjojrRbs/+maPokS6U+rF1Czr2zyuKut7OxIbz3glsjUkTGNunE
AirZToCYYFxJw1LKtPr5GwFr7eJQ3Mm2ceOJYty9axUH3nbaqhxjauLjdGX9hFWr
8iRgWRB1mm6Ser2sj3T5Rh2Sk+/SRhBti74RLrBIBW7rgYW+I16W7cmPgw42410/
p7Qj0TRKALargUlvx7iI/xRkNJWo7m5xcII3ENVnbS35mwumaHLGw0jW0OndlHv1
6bhzPVj2+ujC8H4n+pVpobPkiVCPUF1KfX40Q/OC6n3wNj+L2qqWvgGv4pfVVCnK
MqW85w7Ta7iaN+kNgPF5cCC1QQ3fzq8/a6/jgJ3H4t477VT+EyRaoXlG3FqZg0e1
+QrAt1C4U+2cBkHIiV+VPyUSVhszyr2qX9+JCu/MATqA/iKkzaT4zjhzrfZVg4+a
or34iDnQ+13dQ4z5no+aBbciuaWDhDSuAhoo9fjBZwzEur9DdbM/RyQ4yb5sm8dg
/8vGJorEflI3RuR2HST0x7+9eynbIhnY5LtLuMUxsaPnT3VfIDtNQNMELR2SRsR+
ezshwbCVBSWsHXmbskCCpTezqFFkVhRAUIaevpsGMKpOUA1KrqiJDV7RHGDlQFib
WgEeFe/pL+4+dgXZMX4jhmkXLmLJn2tHDi5ExDBVUQP9fkQVXhhR5Rpntx9GEZ3b
dBusuqcbokWYNdx1mG33CcF2Yf2g3aOToigV7KV0XZzfnQnanDmB9V26+wzxfpZO
166DO6Tp9SE1vvVwKAGFI2+R8xarQjiWCLARkbHuQDTDwIB97d8FZAO3cRGG/VO7
FqwJY1gsAbYornE1VSdkr18zH53KKShtyOB1yUCrffAXCzCgGhaNKDuWFQ14EV5i
2YM35l1AFXZP5OxauetJpK2SRkr2xRBNM246X4TPQto5nb1Vwe5Xfdy7AsY7bkyS
hPmQa+bO2xbCA1YaQ75E0iPQc3LgMz4rLwfBad/OGGHjfxkZYzthJ3E6zWN6vuql
l9djxhRq+/AaA63I+yee9V60Q0pIP/b2C79jWBqHrh+Smr1Qgz2vM36xGb4cYpIu
idS4KNq2ey6uBl6jVEJYKfjJRWnOyoEOlXC3ijh4orTk9nKVJGgJv0+O0a2AveO/
xRG0XMGppPpDYIFTsSy1KVuGRrwGl8hvipoaETp4i5KYRK1Ehm9MjZZ2bHBeWaf6
GsBPGC28+CRktafbkn3yrZfC3jxqrJrM/2Kmy+iLDWlmsgYGJrEBDdosLWygPnzt
/1hdBi7uKLknGSwWbQLkWy9PedPLCh8gy9YC/8sbL3jBqjXNOh0AJqCDLY+CZ0bo
CNaH5mx0NfiKWAxGJaJzGju2uWokN72RqjZCtf27jOO0qs/+lzziFHp2mMeTZBo1
dft5UuAh5M2mOoL9gBV8uZp0dG98P88w7/CQ2mXjG2NhtieUN7+ONaOU1Tej8gf3
sani0+XddSjjWMN+vhMjeYkXJsMGpwYNqtyZedaSECE4rJ3NTlN3CQ/az57i3Omc
1n6Qq3pG64DWdWak6cXMwRrz/orF4uUzB5w7Gw/6faY88tpK9Ty/ONNjA9D8kIIj
fVOR9O+OSwqR7OgMCNeOSK/5DsU6NFLfjBcGSSYEoo5OjLp01x9TQzX2A6kH02xK
++744T1hJafiWkgE5GNI9EHQW9Q3cNH2fCZDZ4AoYfg50h9uHqsTOursJd1fixfu
bB5GEqRoK0kJZx7xGznMKbC4l0bM+/j0D88Zrv3Eq/1APgLoTK4idpatbPPD2voo
L+e1fwkUHkYa7iscXoReuKgAuXCOFdQq5FZnHTQt1ireu7CJnxeUYKUpzBu2+719
B0m4lhDO53iLNoGYXO3uJx94afX0DUjj+AZtGs+MlUHTenXZToQarFwd/5tTED3d
1YDH/1olPTsfFNzGFiPylZ62QeWmGVk5nFVWcRzAlNqc34n0M3xXJ56OMXThS6g2
AWgqmljaWKvT6cwRIGgkjDrJPq+sCUOSok4OUckbTpoGz/S+wV5aUozCph53QW5/
RIXXo+rMJp0Yv+HycqBX3AlWvDX6NEpE3913EuvvJJrq/2+Wpkz+S4VlPW54i/iu
E43QuDcBTrJAFzZdRB4swFM4Izl7nvsbo7XxnaIrrf9vBnscrg/xEjDUxdKwybgO
CzOQeYmjG/Fn5UrD5y42VovMxvAwVxbJompHJ2qwaSr4jd1700bsyrJZXlcmPdDQ
Vbb8eFs0B2FnEmhuF5gXFcgFWMpVRFonnjerpbOEsdcn3zMsIDX7TN/Bw7ka57JB
3vSt4QuFqy0DPXQ9scjFEBcpVJ5SWy3VHann/1S39ukVMeO98w9+FSOby4EGrUpI
3jrSdYPI7eOxcqk5p/tT+pZV82/0utegoxsrELRLEft10ysfTClQNZLEFxWfUojP
Wf+3uYnw9vwsfs0Iyel9sYczCstEdf/7oRdIjxw72doTMuQGMPp9abj3k/+5uqF/
ZF0V6+pT7GEe0vA2hBgQ+ClslvnYvAJkEzMZQIwsTHIviAVmTp5T+PLKFJRcfAUy
fk6xi1yYUAPAYIh7A3yvIIPiPZf55vSpNJY25JEer8zcI7pQ5UbiCFU224OvPNxy
SerxxQXuhH+eMpdfF1e9X79NKvyHEOKpTfT8wxn2WONIH0d/WuFBvKjSBY8K/C30
AourF1Kj+QP3W55Vn1d0gv/4uwORumoB8eaIvWMPgzqNnnbToBCZX92lMK8NT1Sn
7I7/TjueEa70RD4oTzMM+lv1i9b3EcRZfEo3lAR/cPK/qVJYpy3jC632FCikNKv/
mdF0BkGQfhcVZLFJvc4oMQX69oQqJecp0B4Qjmz4Pka7aAu/XkuaNdENnlSGHmRx
1YbQIYhPv3RY3iP1dRy/hPdTbwT10DAoRGLIYNTgQqbzo0x1RKHURC4a0alj9cue
Zx3ghpPSEul3z9PC+Pf9MU37TUXKMKZq8AWbtEdX3KXh+393d7Z6AZTd2h99D2Kk
4JcMq8nAUEYG8UoRUzXGa3o2wUA3m+lOHSYvBASGHyOnWvBASJRfExmKl0X09wbh
Qqhw376K69RvreFpqWrlYS8fZkztVcYyC7PbRlkx/WX5z7BHcHWN1d3aUuj2SXaM
37Ss+t/LyhxctCqLZgW2SfDfCztDqiePSvyNmnYUE6yj4LZuYmdCAwGlxtnomE9h
Pv3D8p8QzTxh4hNwJTPM//295vo7oYsUkLTFYuDUW3INSjuWQWWy1m3L8bgHKrv5
JJGP+Xz9FOG8iIKXUtZLUg+B29TU6HRO7ivsbZXHNwT95nj4hg4UVvKl4a7MSQG/
ux5yXB+PKiMDdOci2UnNPo9sq33yLdQo/xiS5RPEmebXzDNd7ewUU2vM0OBbLnkT
0J5z5qeunfKoRTMxwcwo0ybT4wYDNF9bluX1xTGcVkJYrIF0tIEaRAcysEkXNuqm
kxRQw0veujQisOx50n+xGM9n2nIRktaBNHUMKTqm795C9w9+8CKZbHkD7yPo6nuO
ChGp2xSxKMc16QywV/FPxZBF6BkD049XrFxWYDHJl+hKw76RUSITH+LqUGmPk0to
e9R/2NkTiJbVaT+E4tTT04ePdylgnG2F1eaEYTtLk4aR2WK+a6BdMstO1fIC9czf
kEorokFQcmU1ovx7t1uAKqsgtfEpm3RtZUrOZeGX+oiDazN7TwXZDUGL9LxfAITu
Kclq0ZXMC0xJE0es8shumungx8NY+HS/s9yZiHFa1HeaA0YQSfvQFDJC6ArG6TA4
ehw2U2UmyxOiQJQBrjYC0H5lGo9hO3aLIyhQ268oYC7UD1mHWl3GHJg/azyPZaQe
3XEgaoA/sEegEJh5QSvMSfu56Y1emG0UUOluCEuAlh524VpmlgSSXWm8Ik6dhm8/
q6iAz27fmVlj4puUdkUVM6QgsS+Zymc9Pfp2iBZ3l/serrvQMQZM+SqvY5/krkQw
7O+P0kZyjFeVyPhocGaf6OtxFn3gFrk4nh/LZOh3td2GWqaWgzprstwH3ZPTUS3B
cV7Y7mcZTAKlEODhIHekV8Qi5p67+KM1lZJtZX9voIPQW+5HHAJYzasn22MdJ44X
28MgIJ6zB5286j0sdnuLh2KIM8amJRH5Eq5sKvLUIisvYroskjv9u9GjWYg22hJP
hF4i1zA9UwTcivlK9ZrTpjub9RIXsJElN/+qyKgv4TTbxj+C1WvaiGd4Hb2GgTxY
mtldH3NMSDtuQQvNenuLHVPL8xhwWJZaybX1U4EYmfbvElHH4338QENyRH8+jxA2
Z9UQ7s7HOUX68j6M6pMq836kYnkuMfQmYRC6WnbTLQXTJIGFjFG9xaAzxey3as57
iWOEb+qWiTw6S7qgo0B9l6PD0fTRSmi5/DMeCQvwPv0MF9ueOOcJmWsJ51Kaewpz
tZMGT8Tx9byOZDTZIGB4ziWSyu2xYnlOwwhyvCHf9EYZmMzYDF1muQIBsBYqVmow
ZB3kln77PCpcOYLMM+gNI6FYB7yAmGS//sSify49ynKG8bA71xmAEIpz5iAicyJd
8Uk3ICZ8yGeKXZFZ9uJS/nH25EAZhQi3zfrPRlRXxG6d/2kTNOi6NB9BGXENAXco
ETud9cSpuW0eTzMqK0RIzHYHvxwVwg8+LJF+IHIVYbWeMfuKh/I4Bedl6TwiyYux
pupZVEqi55LYfb+Qdf0nkB52iKvIePN6pljcml17HYWwUPrwCtBWl93ORTWSWsHT
JCgadkcQetVW0aDPNcQfWboww5d40E5TFRVkUlKS0MH0nCpMH89dWqCeRZaSO1G3
QF2e1UjkKmjc9+nvqGFVPY2+KjCHNdzNT7Q8QX84rc9J/r5FmXkqhkV4y/86YBtB
BDgqwXTohj8XrdUvp4nGNhK6WPpHfIkp8rE5xB/lbLPhhTXfga9yS/v/SATnUcDD
nTIurTgxNy5PbbjNp0Afk38sbABApFY8IoX/lmsT0cp5ULmLOzE9Zhz+sfqYQjYS
TNO31FceG4ErDvXjdqF0TD+efyJoi1K//D+qpElXnJ/HV28rG+4hyieelccQoSKL
Bk3UuCIdQgINTOD1GXaOlwWYGBAKdzF9gR1yb13qslOH4F7wUD1rng8+gdUXcRst
7jE4Vw9Aqtf6txSBUaAk4Tzoj7CaJRLlA4P6TIFLtXvdXJyTT3uRSBNKtgxKq/PQ
k5jWnjEKfmNKrQ0rUidIhwMf/AL9rQrkGXqmWcg7uaLwV4fqyECvJDguRDUjMETz
4ILmuTG/JJa0/rdOwX7fii6leSrsiBl97F8+LZnlGLU+ljgqgW50GaK+tE4rGq90
/UIqGh0uaiHM2T3xvEnV95Vy/uUD7EFqrMSiVBUBHEgBZgEDeMoXnGlUG7ePp0eD
r4c3uopkB5LTeZHcAi7t5xgCWPm5CmdTBuic02ULjgGOhjUIAJjTmP8e7QT+Ct8b
j30H/a9ZWBqB/1E42NGBUM1sv0QfA/8B2J0m3HeXw117EfnHLg7+T+H1fRADGtHF
LhC0BuxS6ZNJOcHEwfjacDb5uTQenAnn0dvNn/BpTcMqctbDz6zP0yFWGIrPmGgK
Vq6VbUley3psNAR2ijEGKVa7EV4J5CF9WkqnJLbtMIdhDPBC/iECGRRw7Ydd4inl
O5LjSMrqUlOXa7FOjVfQc+F6wASVabSjK6ZINfTlCgElar2swOjkjqhSqDsC3mdI
Xd9IiGAnviITwsAhydFuJTklqVziBH7AMDbDc19N610wt/lum7strEs5y+1smEtb
UJyLdeFmcp9Ql0YmtSvQovJp2ywGug/dlHk2Ai9705jrOJkxZQuQH9RgmxKUTTZr
xmHTtcX+hp96fLWKk9MphoRHPURuV9Ag/adXYALY2JVcHxk7XFPnW2j4KXRURomm
kAqCZvoYufWuenrJWkkcUoNXB1IR2o76FdLFxQfmF25WFh01eAm54Bjb7ZByBbgI
qWnptPH1xMTUEHkzO9ZvhrW0fe6Ecf6jdvvTXlS3/uK/yRnQ5ok//p1F59EdNj4L
9tMlzqLPxxLS3OB+0T3IHkI5M0uRIpTfUa6kX4Fh7x4WyAPomgyA4V9nFmBDw71y
/ujItYuctq4pzW0hVrjEgujGpddFs16VWU6prZHJcqsPOlaUopgtRlDDvLI0DadP
OL213LdGoZFLSrggRB6ttch8B03vC7D7JuLDZssAdU0nLtaKOCEIJKPOYo+84F/x
lHXNdy33C8ghhvpkEs4touJHPYxxKxudd7Gua6q1PMkwJEgqxg0y3S3R3xHc80W/
nwdtEOIu10Wc9dRMxz+En6/yLe9/92Jg4QDr50GLmYd9T7sZwhYSXNRaAkiJnOu8
kD47DWNYJvRmhE25FTwtOMYkTM2UZ557Ta5mWFOZ6AJ9AkrUdBLm0omX5OQ7xJ/0
XFBss1DzqPl/OhLd1r6JbbjWH7bLoQuKgKiQRqNjFtlu8IgIU/OzPtjmxbEQqXF/
XnKgHQD+iDin5H1U2mb5PBWapOZghg3tDfaDJnLR3TjKPCvebCcy4GKp5GnaLFa4
yEwdWVPL9VQssQNwR+XCEbnBHMrPLscAlMSnaFyDdquLQ41uzcDQX8qwSp8UskD/
D+mGh4da+bZ6iRjrLvEtTZJFqYiKVD5moE4x9blzRVvfnX0WGPZW0vK2/wFV8GPv
Of00y3AEOykyD6TrKHQqcwOFf6C1kFYqXTWeWLVUgG9BMat5zJ7fOL0yQ5mq5GT/
zdUwiLMIunfY8MIQsGKmDqyK48mBsgvw4fZdfJ8uyLIhX8VQ98M8Hi+6zTPB61wF
mCkUXE6Iic411CObxQo7PufSAdvGxe0WmHgrHW8mJoEp1vYtI06GTvsjcr5RHuEa
9eYtOCEpKwrPHOY4W8Q/4rStl49fUtqiU9JHREQqoJkxP0CePKNmSbAJ7UQhWLvY
p2atn1yT3FDLsXsIt1vxmOvgU/LECbL/FH/dit0VyAvXuJ8Z9iY+BGojG67pK3mw
x0Qxzhlri6DntdKBoerMNkIRDgs1mC/M0dUEQ3UQZxRG/36cxckeuLBC+pwe9KNi
R5/dSN5g0tKtdeRIKp3n/UA9SDh2PzSVN/M/JEl2XV842nZlUIscaOnxfbWAk19D
TTOr13wF194DN+nR6a0ldN+XgaFJJoyVGD07Napc/p/CZeSowDdzUMHAOqiuaYDW
l/MI5tQaoAMApKOmsqslMPk7zyf5aJQaDxaCjd34X5dNGBuEWE2hWw1LesKQvGGz
+umTgvhCTL7yzSP5mfvtM9gYg9B2U9a88X3XqM5BapJH0pGMMurQJmqvqkOZVKqW
xEa1IShVKrNfyvvNeCKELHoe/gtnI4Xg/XEt/lkBOlz8W6WaUnyahwzYshLwFpG4
G//lqwZ4lgJSQGZYp24j68bp3L34yC9J9Xx6aZXCNK1pPKUHI2/qzR9/k/iw/7gT
cAkEW/gBA151BSRXRiAah3xUenwqv9d/VaHpi4aQ3rGEnG5PrLpcbUP+7LfLrOiT
W58IBI6EhG1RIA3yFvyC4H16rQXwweljLTm8ciEudSz28ZZiQGK2OwbL6S7Yij3k
QxcbXXy1l9sW1jKjC2qXHuGdSJSPB3fexNbiD6nKGZHbDJfqY27DuBzVm0l7Q9kc
TL54xHeYpi84uJBJRxhnlPtHFN070uaVDHV9CN5HPCRO34EjUHKcATDX8LGgidSu
PqM1WUAHeP2IWFkxS9B+RwbTVwL2v43BAKTAr3zc6OuaZQaR9THgTUXTrBLPW9yX
WotG1oqtq5y3fYrubbSDrii5j+alfbCweTPlZ67ZRBAbJ1AViYp9cyaURbgbWY7L
IN2xzrTIXj777gYK32veLo+0H4gzZ3++t6dhaauBCnLrljRJdPLAh2JRKxYXdoLd
OQiRYXI6rkrITOsL7lodk/KsCWX7+gx5KdZgOS48YQ2W/i2fy74F4/ExWeXpd2Jk
L5xoQYm7lGYb/QodPJ4jNQUi160A54cIah8xeOI2bbYxkjoxMZ/wQU4dEzDtojoY
2/axkfqmO40+zWC2Ty34Uq4RYufouD8zac0OjvpDvDwuMg6JjbGKhOh01nrL0HXj
UCUSdCI24DFzLpdkkNqgFjOVOxbEhd0YIj594KcwwNYH3WxlPoYan4YC62lIY+gr
3qf0eWsVNHBWAKsPzxHCJSIQmAbcRrHXR5lc7NQy/b5gcnYMrLkjQKN99Jz7IdoC
Xc91Yw/l1Ql6z5K3SyGH0JJDs/DKnnzSFuyVRr3l7pdNoorbz/smFBcKqA0FQW7y
sKOiv1FTtFTUxKdQ5uuGpHYlYVVCsj2eVHfSzY7AQLFTSdRFlCdZ+FuldNhpTJGp
wSUCaqaG7W7X4OMFYyv9h5qVg73gY1LCR+OZjHoKBLN4ZmJlJl+dHwgQa6kAEGw3
XqWXfQ/fGn9nD3jc4a5CUIhEOMVY4EESkkmYMpCvzvFG+CCJ/WtCHihJGjvz9uBW
mCnv+E4E6IABxTzEbZuxS3ae0Dqym2PtQpN7UQnTpkyWFAiu84ZkwAtgtiTY8wK7
CH+OhdWdqDleGOMYHiWVLy/F6uX9ssgYWmfpWBIKD+VE//yL2mPUQXaoirJjxGpS
6ECH5eT1BPMDOVVSFPmafMs96Q47G5VKG+tXr0sr/uPxOLExr/DlDEiD2+3Rz+tB
xUhpXYxicJQoYjguLJ7p1uVzHBpugLqihWBmWsFCFi4PN456v6narRJ/P+LNDPVT
PKMKIE0+udBZY/YDxdy0fLVCxI1UgRo9rH1e68G6ptAsdvz7BPKX+r6Qw20aAIEe
Lbe06iJlvxOMyPRYWQul4EOuaG/kctHbEvJbSU3kTjRa8RmPIs3lB6MU/lWuCAKZ
7eJ1j0Fu2lzSVZ4stSf0l+sOx4nQUumF9Kx6fwMM7XTluo0ZbhzBVc+JvfPZdA+C
lHNMS9BKrxIFiNya3ZEBuHGMryPac7ubuSOJilvxHTzC4/eC+7Y1y4DXzUGD7jz7
Pv7pf7WmR7OwSa3JDJ1T0ngD0UhLDMu8eY306pXRDS0qJ1T/kZxYz3ca3WEUENzW
mCkz7VpSj+/M6u5MJpD6uL9CAxvyEaTBLexDog70kw51R2TI/vgUVbLWBzMsTla7
IepVakq+tJxlz6EMh678joO8IX4kO+elWApa33y18p1/YpU2dBL3/s5UlXi8tAKJ
8MqOO/fB0nV02/74EMGUw9SBdncptXi3qG8QgdhqRJHnVcs6Epq9kbPO7lo2Im8z
TjwRaEBVbswMa1SNsVrxq23jZ4Zb2fiMB7uEk9GfNiSmd+CB9G4twHdAQgy0HO7L
puMnW084wmBrCFv5aHrs2tOg40R0iGE4cV0VzQMDlBls7fXPytOY86cl44JVB4kr
cFFmFcLDMQ+fOgoITNW9lvfwdKDfgtG2u3g5YaBBqy4qdpGo7OHJOLH12ndT6VUc
mPICrIepImxyBG2dqPak0B5NPAsO64aCZu874Qkwk7ZUZMXxURUIY4nR/9Y24nxX
W1u8oLhB5HPXjvBsMdhs0Uxf3Ms/JOzl/+bVhGqNud/S7fVJK4BF1cpeFh0JeIUY
x6rbCW30XMIDcYi5etBAay1OhoPxEqfXxd5cUfBXlHutxkQ9Y5s+/KtU8JzOtLD0
`protect END_PROTECTED
