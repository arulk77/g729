`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMnEMgt/0gnDSHEviessrNUsY47Oc480BnWm/JIBhcve
JT+njUOGqBKuIE1ZPDFBH7Ss7SkzbH2LqcrIELriOsmuMCQsUugbOcN15exh2sK1
cXg2Dpl7nA5SvuUFFROYPmfqCHqtwRz4fjse2m3eblkj/xnMBSo1IOry93kE1g88
sowe5e6k4gthxv6PyVuoC9pK6BQehpnHANGDSJQA7FVThUcRC+D71TmaZWqEzMuy
XptJNxeczleBAJ1VgQRoU5hn/doJwRiK9EeQo04rhz7EuTmhMC9koI4KlUrkYFUf
yjXqR8Y+kzWfDyNZMHRNkJn+xNaxnaOc5K6GH5mnyPF+Hmi1FOCoVO6f4yYqssoQ
Btw6sTB/CX5BBt+Qe9SJhSztzMJ9hdOartl5C8LvpTM497k7+ZjJ1mURdOGTOXcU
OifXZORYuJFmfYCsk36Xh/RnynKEjLMysk4QjzwrgZwgIWTHOFH0lOk6Q+NYU5UH
jOvgBNyhjZQwWQn+bsLbfIQFdn3bLYGykj3AovqH9TsqY3gF2SOaYaQnCAcjHxGL
zdTar7uJp+TavNG3S5upyw7eiEnky0SQm39fqkWW5uIkkuYnDBOmH7sL0qzcE2SP
U/ESsnfsixTTcNPY/9nf018CkH4VoJpq5danMupInT44iyxYRrugLRmWU8O0q0Yx
r6lrYj18LEFk5v0wx0L5BLQTuki7/OpZwzYnCtKBfBAwf1+mkptEhOjff9omkSRV
BVJrb1lYjLMo1ehOyCWOLsOWhQGafONWw3pe4hCUoqoqI88j7fAdccn0qSCnTbmW
N524UGVEakaq80/gm7UDhN+Iq7wxVgwzkC3FoVUT4GuczX8gVzmDw+5gTDmyQTec
OXxAanpMhlePe5DnKg+F26e45Ml7eD5SrkjxmDat88kx5bKjl6Oe6pbmoNyk56Jt
bqidj5MwKhdY8q08jGWoASuPAXEQn08ZVX62cqV8x/ILb/fB4uHPwvUa/vdS1/uC
`protect END_PROTECTED
