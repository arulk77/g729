`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK2QzVBF0tYzsJRZJBJYYABCma4SXOHxz9VnYGzLbMl4
5Cg58rxKd4nMqZccsJwfFnAef7u+Yr7UVGrq2OdNl2HIy0wHQFHwtQxkfXFA/2Fs
RkO6uetS4prNGKLsVNcRiOhHZeRWxlF5Wirl6DAHCZlXZ96kjecBCYnCYE3/JHwM
RxkWqwcxZ4GCOvcBom3Xl8GWUYzR/OCZ8v41W41x0z+MHRqFRSPYyPlNWUaAcrd3
ivXgoZGniNYiCg5ELN4EnTe2YZ9q2JuPl2dlp574sQx4u3tIQUdowUuOwnG/tPpA
Edn2g4NKVdynv3DjVLituy2oQUBAfgY1PN1Bg8spg9AWWLKXCT+DPXDe3ZxsWOR/
+MNY7wrfmRlmHnYaObLR0UW1OHsXGN+pjB7DnUu8ghL1SeUuZFq2YIra72R6moP8
V9SqN7a4HN8h/p3y/jYEzLWGNphBxKdB+fNGiZ58btP4Or/8U/VXY6qp6yittQXG
5547SdOWi1iLb0kuweAMrNr3edlqFK1TYR6HVjvU5raBxmisUFiQZc/MthHuIuRG
AMF4OR0pJflUchc0EOAgA5s70UndravojPhKF4/4E8ASNhFzkVkg4N3hOOCg6fjI
kJ0pchvfV9lwmHRRP1MsCyeyA3yHvYRm69CoPKkOTKzzI1R9t2kSgsADCf84JUi/
D1cWHYxeRJmrSjeDN7IxpubuckMVbg+QZIGm35NpwDgYwYW9eQdnD52XV5cmfa5O
091LVuSte78uGeSdYF8Kq4ssS7XY1V40OJtAkJF5F1HyXPkwSI+uKefb0qzJ7jeF
WbugnZPGA5yFTtHilfrTtLnQwwWV3RE1OUHyabLzmyE=
`protect END_PROTECTED
