`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
DDG7Q5MkehB1ZlrJkAb1Zn9NFpnYK3U5mT68s590Uq2HYhCi+W3HT2IiGXepuA8W
cYCmxDmXm9X4a7wdUHxcRA5q+z14LW4NdOJ/06sejlRlLWBiXCSIpAPHZF1cni2k
yFEnVKG0N935aYgaPFtEm0srbdnjbFaZpbCbqf6P1FlxtChDPVDB6HShK/SeqgKf
5tE5TCrn+/Xp6oAeyrsrE5YVlkwN8zgsDqS0nilQ8gWgbxYvgtHbmYpMi6WaGJXv
Xjg6LltZQxE5+VR14bmNnprVzkbNfpjs5dKLlbp5Riup7W4RBmHmQnKKdj+f0DQ4
`protect END_PROTECTED
