`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAZHh56qsDFONy5eDrCYWR+1IfPyN5h175Wk1g+dC5NLW
L0exFIWdTJornrmYqmfzOk9Kg3etFPYBVjd9cqhvyO4JuZ+XmZTPXfQQfLMoBJSb
uyvv85ikKCvMPDDXPLReRYctziE4/h7OUKL08epLf4RNVoN2r9aFy9xurCmJ4PY/
ZydOAOMta4oN8E089rJ/WhNCRCDpY/pjyHB2UmAFdQhtWLwNassrU+T8xK8hdO7A
nxBVB3GHKIbo1m5NMpbr1cdttsUvvR2GzSmvkvM7EDV1OtFAYbR6CY5f5MiQZeQN
j/lNroyAXEqXXgktBPiVWkbZRYYpVbTrs2nfwhX4ld5hyR8X+eEdkxoWgQsE9F0H
Izpo1FSzjtpi9T5DK/VZxkI7fFesfQrRhqx3ycnf9KvG2Dt/KB/aZUZ1fY9y4pWr
7qK4CtV9K4HjsjPFWAz8IbiEQGASaEgAovNGjb9olbepaRyG67biCCIa5foR+IM6
RvBpKzTN7BL6KUAzPhYpCeAB3SdsLCghgsel645MPbYcF9thjFdg1rqhlJTEfVbM
KY6E5o4g1bx04/H6iZnsrXAahv7imD5yFX9V2IwYVzQQvuC13O6lkgGYCJSAAe+Y
mScReMB+Wrf+r6EnXV+ssQKn0TUy68ea7Y3nl2Qsjn0oStgxqtxJ1WOw1ZXi8pa0
P16sNSYpM5tq9QNPO31DL6tfXQ/+lfgvGNRkd9v8Qw6uyIkI0W/tb37IjEZGTX7G
8nOouJIFNqleLYxorJkptoMhH/YxtSlEKWaMOxv3SphaAnpzc7v9lGHypFlT76rg
MUEGrn+2hyUiRTUvKV4j5EdM7YAAeYAqPEUSTq861+O/zxHmomWsnrwP5vjy7WKn
ewWO2kJ18ySSUmN+2Mx1GBFL22fnbDiJ3y3Z6+AeKl+kWE43Id9AXockKfAw4UWU
OAMzk25dfP34bNw7UQiB1bcBfjl/uIk0jJ0b4Pmc2IvPww13Ql1yCqvveRUsACvv
sAUGk5UCuqGZlcOEen+xxx6ef6zrvPvVForEZaknb70WPbqLv4441NNIvGvhGDsM
2BVoJKao/K8lfVp8lUO0cqLQAsUA/UxQDC4kIpe4woKQZnf8MisLj+Y/l8Pu0F3f
qBkiM6gZ6poEPGc1UswJpVRLBPeUUIK1WTBmKfE4tKrIYFtSTvwN4fftrp3VdoKR
f8HY5OqVhrwMu0evOlRJC8KSEpPzE5ovRQU/Kj/ciWDGoXdQoLLHWNzgxRAJNWnh
j9OfhUvvQF8WwJIbEw83KrXqExjKVirVKmijVFVg2gJHTSmIgzWvXW4/DnavKJsM
NfP1biLs+CCY9YizzumRUd7vf0RzcFGD64THb9QKtgqVggyvkxMfpsxUGgYMjNHX
kDT1lljmzbEcCm9SK+sMx52sL9z8kLzQggdRS6BZLnG6G2JJbqgWNewHrLR4E8WF
G9YANy3cmKxTpfUVLRARPWZjlXoPTdMYsJWbra49dUGo0mvyRXRj+Rbz76StHLUl
ewF52B1NTyBzXVJE2aimr+zrgdFkLWQOKUtFhqjGHWUzXHOad7xI1OBegxIYVp6J
RoR8dZDk9Ys/WBAkzQL0M/Jq/8zXUcZPSFwCnhKmV7zZQGOeKmkgH3PStoSP1tIc
MJzfPPO0wC0RoD4CJnxO6mcElA7SIo9zqPNyytEYqum7b1QuJaXR0IlDngxNzHr2
/pyuELpqIBXw5pDjr3vPSR8EGzVsy0OVZ7goKkpJCWKbCH4FD/hWgW9z/NbQRw4A
upk6GxuUpwizPkTUKLVVroekhBx7MARLxUDKWm261rx8xF/MFRfdsFCZmM/J8Sel
aA6w/TGICQujzk+Hhc4v1MiZ6CQLQGP7Utb4vEaz5cPwZrIltcdi4UOB3xrMXZza
VRPdTb1wflhUc57wO3O8xtoP9EA08wh7lVVBVi/+SGSaCQKUCz85fhB4K3nfuppR
lsZIzUHjRaWjxTUkO2J+N57hMccTQUe/J6ThA50C42xTJPRkzGbaJ5DYYqxL/5Nt
pW5QkdeROt9Dher3jAJBb5W9OC0oewNCKQYs3q/QmC7nyLjIdIdwljwHZXko33ZH
2Wv6AOPjWYsc/tXg+3OgHrqqGH2gaTX12lGNaqlUwN4GjrVCwj4aHqIYu58HnWiN
8BxRTyJfSoI3TP8o24MMWFXknvJSDVjhqa/AsFRcJdahnGthtx+WeYBwpxs42bTY
mq4C3w4l+eOQeS0N9ugWMljk+MtW8hgaJAJ8/WZQVKMA4H135oqZEP3Y+Yb8yoCq
SEflPqJ/+s9TeYk1l+HL0LQslOIlk9qb9ij8gAdbZvPm4bK+YOa0QQ3EWxWvTV6P
7ziDN+2ISlnlIzbGYGiu6gJlt0qTbEClP/5v57Ow9J/gPbaAfmNbVzMlnfkfmmCD
2+mCx4L5zWjICrG0sXeTdpiHXbr+wSMPKzy1iu3jZZAG+HQ41TQ1pAnJgwKdOwUh
uh+jkbjKwyr4PyFtXABFanbTQmBOKV1mJ5QQRcjpyrs7f7H68iY6P9DyyauTgGDL
Zw2OJxjrrXLWqem1rIa82WGiMHNlS1cqHBHdzw4SWSxmsfUGvM+kjeV6MZE9E1Cg
Pcx6xk+4OMphKPKE2xVfuXVn7Joq53BAr4HNVa2igacmV499KGzTa6ifpvW/hfI3
MRkbilA0aUY6eKWKlqHose/eKzDhcM+MKKxJPs8d86ra9ZsikQuM0oA24cMXIW99
rpjh0K0X4lcIR/asPt38A5YpfsAF53Yv4E+1e6dPcNvH0njAS8QFblSK3WgPRIj3
KcTUOHFjQOI6hXN+jN87QtrgpOvqX9x751YXn+T2BVvkBUOwPykUM1Z95MXQ3ph9
wu9IO1ca9jKuZvzkGQHwkR1JWuz0rylIPX+D4Qcwj0e9mmPlzPKUG6qE5Y5E5iGs
IcKV35FpZXHB/VPg9D1khR3UO5+XPNGUFKLDf+23czDE2/dT3FWGYVGOFpJYQJLX
S7B+uk+qnYjlCqjRiPJrFfujysZsEFS/ydiQDLVs9urMZpAo9NcGiH0aP8rgpfZG
6HI8d2M1jThwy5hGM0VdTUYFZ99s6UiyuoOVcd7L3xa6oQU7wMGPQtdfHp7giuVV
l5p+eol0P+LLFyb//GfWgld4yof1OTX2o7K6dgKltL2a9DbG8Sf/b7veprMaDoUU
WTsZAsbrtp/1U7BdLcNG2YWXgjU4CC1QnKZYgsX9SilaTf+vthAnK3H7FZLhSfjJ
qTz4UQQklol9ThK+N3EOhuLhKv2xPNFcpbchgw8x1b1lWlOI7DEcc3DlvulnTdM0
fVmPlHAC22+qRnpudSTxkRLOGmqBVQWh02X1AVly1LgovAyR2pdqQufBqJBPgLZq
Txna1SX0vEN549Qv4rNSO+yq5d2zBx5SiDvZaj85603DPA+UdNPibkY38zi9SxGy
F+KxfdpiPrpcln65jpjWv3okn+M/eCarHRe7UmBppO8MFqyCK6BPObzTkJuS3Oio
6W/VF2jW/Mgr6+7Z2fDO2l6fgwJ+i4EHsLQMRDNj+BcCND38roEp2LIr6YMeOGMr
l4tJDLqaeCLrHk0wVZa7WSrLV24pMAowIJA0V5/uXDVLiRCTRlJzIWa+0c9f29wA
humjDVT66lToiKxlM7NriWuYXBJp+fcbruUiZBbpFKI3yyLNcBAN0wJ72I2qoUow
2phn/MkDHA7/6wl5LqU9wYySH6Ovcye2mZYto9aAu7FdxRvRr5WEp4uLhxr1ZDrn
moMJ6U40lmZ//35i2Oxl72xkuL3O2IDPOUhjf509LMyAcmqgNc3Tog9ZH7mzbIzL
34IEvhIr2qEbzRvC76AlH++BnEB/xtGQsRoQOYBJoAHofWfOOIFQiJDghdbcpgSB
5teGKgs4PTBnJuXizBzj3MRkKugE1fq6FQzIw9dZf85Hl83JFpSfDFe1bbFgfdud
8oSr/J/XgSYNB8VZfUMW8aJJC9xu6hy1oXXfJZJPr1ml3WJWlnY1MdzVR4erS7MG
iSG57fbA+rNP/vejfSAplEDJxQL85lK22YwOd1KSiLa149GrZIxzCxJ/Di+Tjk0Y
SX1WSJqGUBZzHfnCVO/2guVb1o11KlVsXuE3t8aaVO6IOSnIuUrIUk64oFvLb0gQ
xIYhcHxHr+usAy4yX7riVJ9CIbgd4bpzLSDMQvDwIkL7YA4y9AK17Ohlcc7gK2Ia
1AtgFX4RNpi2O1/IUytyiyM6MYpom4sAtXxIVVjTMYFIxJYusr7g4bogYcxeq5l2
8PzGvU11xiF5qWVRq7mMcfD798q1QaZcYFw0MmsPwk5QnxpcvuwEUMjC4Wg2JpGe
y0+BFyJgv7ubURANG+ePBsoJDs1lIaH5mVF9bxmnKsr9LF6hiV0sNPIYYhsHX8FM
n6oSvqhMU7nKUhzd8uLe44q89LtibQcj6gnCZYSWepmetN3XLLSYB13ttMmt2kVo
GNT49QfJkcRL9hxBVEIHnpejoLcmQQ2zX0S+y9Wiwwji8DIcA9Nj/+RCFmld6elT
mw1mFrQtffopES/tZox5F3q4+8Yag5p0hmd8HSIZpGGFnt9q8Sp1E8NszxKpzIuv
HjKOKZg4Mb3X4f+wjlA1YXfxnks1wpSCD7UFtyfLLvw9Au8RT0Pm7oYoFphhPmVf
5sSwn4lyvRm13eUaa6EE5n3H5KK59C6qBu/vPbdGipOudvrgMq4g85Qxi6r7hgjs
DAJEAN4hWaDbMoFybBBhafHWK0EszviMOEhIuYt3LrW28Rwvt3TVeYEs5kh76Snx
5GQt9/LGkUuVQWDjhWy/I8azKxInRmrl1pCww/MTia2RD9IDKklYeuMmpJA6GM14
ZZmV1lXuDzfLllDEqd/StM8nWbDS0z1eMvzuuqf0VUguLo7DpyMxkgJ6s58sLKQV
/+9ccK3qW69btDRV55hWTcdMbHF2IknPjVVJS01bzTF14WPZUB1skzU8+FrbzRaB
tLMY/V031dzR0SLUOpm1IYRkNeG/32ddtrv74qdfAw4Gjoh5QUd36QDNxmPPdyIV
Tf/ymtGyCt+nSAfIzykPWfAj6bPOQ+NUdP0h/DApmKLmhkYKdHRrZFIA0lt6cuJr
yFlJvys7jXrT4in7dMLRgCivtiGgGD39KkhR7uuhXyWcMXsOD2z22nKoXyTHvz+o
hL+jW8j1iskdMGzsU/yJrKV7l4r/ZJs6HyT7J35ur3OfErCS1wslHrhssF6H6ito
3pj3W5F2Sw69+6rFqzgL/zCk7GqfgbpScnrLa0sLqvBUV5TfK1PRn480DVkKOVfa
GGCvzxYkd8w8jYgatooR/y6UUV3UVGSOvTC0wiAcZ0hE0ZXObVy7nETfq07FhHyY
ruY1fQZCJqLRXRSFt1ehmoAkN3lTgMUmrguSzi6tLMDghDlR55NBgEU1CufS96xo
aFodCLVfjHexhh2wax72W4EzWQChpwukkC1S2p9o8Pmy75bFlt0/bo8T2dU5PmLW
VsbkHK1B8BkLExfG4Rs1ml4uK1tisLEmmdJWH1dSARTOIYAM750fEz2QCGIhzUWC
gJSf1lX9JO71ZpWkFtt13GbebGXwWZjRlsxWulB6cFi8Hfmfd5zg1YUmhU9MozXI
rsH7E7oQqnkkB8rJvBK2bh236d19fvsnoFODYKklJMeGjxgSy301DsMsJMvvBkGY
2f7ut61b4kFRkQPOYcjPrtFX3He0JjxTMBre2QIMQVTIdcc8blBMUyF4Wc+nQo/6
ffTVR8okByhlNO5la5vcTcouXyml1RB8PuRLrdZLZnq3DDNMHdvX4i4tVdGFKFwn
isQLpNznewe3/vKV3svFr4lc2cbkA8oMmXAzrzxQcp/ncwT16i2ofWvOiKs8OAW9
FvgTswy0HgrWJQeewdVFXJVA9ahP2gO5Fg7btR0NRqD9WTgsMZFfdIE5jZ0hKolU
S695hxzMIK67ZX6aQO5NwYL67GaNhe1J2K5ndWnT5GKxM1T3r8bd7zTVrwnhfwxr
ffUVd6hGEDKnelDRMj2mXzK96AtWa8TDAkDFEACuS4i4CLrT8QB+OCOaVNroDubW
/gWrv7jjokVPMSho6ssPEsvJQk9gvtXc6GbzSoHo7tKRbt/fKOS18DP0PUKpd2lT
pWLKe6w6Gp38q8n4hYLn2/ciFZ3Jz3PMck8bX9Gxfw1QcUz0qb6iAYA/ZPiRNW9+
iFxKRjx+gwF/X5+gKPWbRPn6cxgBLJL/BlMaqz5f8YGSPrC1wyHJPnWNp6niq/Sv
Cj/vgd33n1796JfrMPOCPuAe8Bm/5BYAZKeXFPNtwyJkK95hMrhD9Cbv0kz3/M34
MVyR3b6OIQTWYlSgKLfV4cskszGLcNAk/kVmmg+YoZNmUQ7yTtn+unLYd4v0GMwH
n0mH0Eu/kyqHMRfLBoHPjkhj7wkphIJEno8Gq6KR0Vo32jxOaotlslUnJ6duDSsT
G0X/Hmeeu4D3/trHRW8OgBn9LaHHhBeTpDizDfu6I2lr8LYIKNGthaOGNEGBHiZv
Jmpu/wc8IBtWxC+Dx+J81yv6I/mHUxU1+8r8JCGAxtjS+IApiJ/+/CXdFffaI+oN
3nKtsepgo6Nsj+yRpjCNbxOw9mph0QKDt1/Y21dQFpXbaMhkiUltSeIEUkIaRGfi
Q7kFHMBju9W3r5cLVy7n47cfG+5sjR0g+2V+mKOOyr7sa332JJ4sILCpNJcRLTqs
Bk50RGte03jf13a3dKfLC2pQ0SnEDDQPo6L6L9gWD/6onpKcC1CvLf6ct3XvvwUT
ea5xbFoq5pOeegjr+C29WOu8MODlrim2Si/Sg9J+XFoLYIKXN4dVdQ2OjGOZyQNE
hkdm5Oiv8izhAyXpQp3uh2tOtoNTDmM+dUwiS+qb2yRlKs7nYhuNM1Qb1B6xeDrE
7RydIhwGf+IJJwIYXorsErZ5/qad4FFgBpkNbSQcmPesxjqOlVlCOjcmjrk5wDyp
fbsSv0VPEfpgCiFchqsb49zELWpT03BUO2Zcc0twu70EXibKjwlDZU+rOSchKsej
Jst7FH4YacTc2raXSD44lQKo5lKQzD5T+5XceiogaUCv4l1t4FsiV9kXjfWH+cFF
eI5IXKQWNiJuMUKzopzh4hH7fMeZP7Dge8hZbf/8V3FJKFNsVqGApq5tY7F/IxxR
J57R9sdLLIYugFhz9pE/wqziTwjLoAh73xEPm0qJbB7WxWFf3zwj4id0xjjbz3qM
dKrLuMHEST2InJZ9g0aDVlD4EW1CVglt3K46/h1fhVVSnn4ScDKej2XsuQixIlLF
uD+3/6wBqH8G5kbPfhIER+1Vk4Kxh9r6leoQUwHtjVVIq8r234HH2ZloGE05k+x/
wfR+DDAD4bGRGYME/VWKCaiv8U/8hvS5A4xCW/NP3YEXx7Uyhm0e2vukLcMcbGfz
UB05+POjVXwtyAQHke4gZ63tv1ZrohOiDBomrp/Xy1phSyceK7KV5WRblf9lG2IO
O7TqplFbGwaor/zxWnvO2QR9MVlCagIOQ6T/y3p55Bo=
`protect END_PROTECTED
