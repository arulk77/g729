`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
5SWNf39yNd9y00JkZE14QmxAxjDh1m3hJGt1wR3tDHHMHEh9LoeDcyTq2tOLYlTX
gdrHEi2S7XBF1zBDx3Ir0qcpw++ttaVJrTZZcT5PtFVu4SrrBS5Tg4qJAE9C9wKk
P3eSKW3rkppzKcg4LsfycL9fNVk6oBPDtkzP3yUdZNCed+UTAyRYMrqSox0YpDmI
Wo05ySH7P2Q1/3rTbcSyiJYvNz6nRu9ATNUcC1veOobBnroNVoVgOw8dkX5+vM2l
`protect END_PROTECTED
