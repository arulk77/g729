`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLrmhLmBW0KIN8p0TPa8C4R018Mai3oZ4Dc5kpPgbAKk
abcLOnOO4IxLx+Uj6oA+NeZgaPRYFs3ePbvNzdnJRoFZ0806v9NAvxpEa6OVP4s1
hu5InDZOijrW5LkQ7+W0dalziZru02bIJCgsDJjHo7r5AOMfpBpb4H9eUQXXyx+J
CoZjYBWMnAZ2H9qMf+qQJIL+/vlzvMkTPPS+rfCu4GEQbZ1JXi1Un36pNEsWkkgE
AgRq+7U1DJ3huJP+xjYqjcYP9BofFE0yibnV5kM1E1/h6yreNla/PrXoWLbtWZnQ
w0fC30b/RVzOsmxnxeA/uhakp3qNHI5hxvLd1U8iJ88sPsrTazpSJfrYHqzp0BfE
K4K9A/eMd6d4Q1pHH0NyAZ/7gOcC18KFlefQcJrdNizgj4Zpk41jc2eLcK9rYRJN
0Lc6ALpudem/9uF38kdZKgpjqDLtm3vHy0gt6j3k2aXkOKN3TSwaPIyOWTSalrwK
`protect END_PROTECTED
