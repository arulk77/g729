`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
72DKe5MEZSH9IT4s+0rFcImHc3Qcec0up4InvNz05mk/o7Wuw8AaNnZMixWugTqo
g7gtyzo6Az7cb1UO3F9vRzjk8/psy50Xy4IduqWvO7jUm5SJQqBavkA8JL+HOsqM
wy/9pHqZR1mAiTxNFD/xn3kY+nwULfL1cEhflkuqnPGZpdkqDyU2GAKZcN1eGvVb
a7FBdA15xXebZuGwFhjqcP9bv0npgWIR6oLieqc6zhlX8CPWEkNuPRUkKkOVARFe
5hd9tlh+BzX/06pazvNtQTPdlpQo+2MLNEPNJlko9jkv963CwLdGH30fpRQl/wam
DKVTXBl0r3ASpOjBLqtuwkAUOr5g1y4LtRnVO2FskbcGNRwb0M0AEgEwDs7/OLYS
`protect END_PROTECTED
