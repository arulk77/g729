`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHfAh9PLHnWoX503ltxwWzjCMl9k59ejF8DF+Mc42tHy
CSN2dZqNuFfqJpAIdKDFqXY/hzcwoc6mKyrFCFTMpS6fG4MtZI8uey5zdLLPMq+I
iSUJhIu754cgzLlYWhWRR7VSdQnQrEpq9mzfGmqFbUQ1FNFLh1ywBQl9M4z2/23V
`protect END_PROTECTED
