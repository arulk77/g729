`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8STBKHJtm/IipXAv0qTHY3EQqusvGJF5JfGuTiWLc5YcP
a72EkR8uDt0ZiEdxP1OJAnRxtgQ3PPuTT0bP0Pt5i6/+4ndua3Hqn0IYJGYBiNsa
65+lahoZFiMZHMMcllxXCnNK1SN2JmkDsyKvIqf0q1+OM5Foun5Mep58mTuV54GI
cxo+Wyjx4cGC1WxLTwtJwNfPJWq1uH73e6gsjDL0DoxX9UsDLCCMobQzu5WOVegx
XZgJ/neo21ViqxhqMjb9Btd4AW1hYV5/FTx8qA++Z3CWLJQSPRTa01OxiTIje2fR
qHFnEEfMuq74V2eKKRyB+8NL64Ei0AV4wuREkQjcXBuenInedJZWqtIeNFGetJtL
xJupdUNn4DuT6MjGRc5iV827iypCSvScuSqIYo1wL7/3yt2ksEE4uhCcHv6zZN8u
wZDbVpQHbLxOCh25eMwsffoTm9ylooFETT0wtsRvauOkZwYsrkNi0cEpVayfFfgK
y8vTCCCcPP9VSWUwn+KjqAMlQo+4wiOSR9NcbKnJJvDu5nqf+6TeHtzP8eLyxMzg
fxzFDIm5CEBxt7JiVTDzG/8O4CF6UWN2E3aO/HlQn/vnF4mERoajGr49Z75Ikddd
Sm/yz6vOD6X1uKaH3F82wjolrnEPMggzh1ee6qkXRvNEdomuLwSwSoC3tUMePoq/
ZJ+IJFA2SfadZXc/nHGWMC2nhOSC+dY0iyw8XxLf+ZMAiw3aIziLeJgUasmRDm8f
xxMKUsSHcugVg70Y0jv3CPmxPcpMkfygQS9TMr5eJcBBVkaMq4fwz0T39EDFDue2
deAlLKZp2zy/+4E/u491N/Vee4QfA3YjXNFY/kIZtNtG8mASyuUWGGIBfE5aJzhe
E1uNfKsn1JZ1fj2Y5U8Ne1rnZEiIYIKz58Thn+mw/Y39Ar+n+Y7W62de/a2x9E8n
/Oi5tDIUj4AJrX7Vepc9jdH3cCUsJSiLzpCbnx524bNVZytsLqHrJmDEPP3kPHdn
gNGC60K2x+SneIDl3U0QdfIVdDFtLK58gak+Yvn2r0fDU4+i6mJcRsxk5xKnX3NI
DSpUCa/BnInzdvoR6vup3IVgwxGUlh+x+X/G4016hh0046JwXYVn9VLUx86DQzSR
JabH1Gi3S7CaALONp8H4ZSKNV4FG2Imi0NCfrQ4RhmUGBexVD0JZiSqOInT8Fo1Y
AIwQ+2Nq+V9eaptXUQ2fbcAHK2nLsf2MhS0WP1YLVUwzSGQvD+U/Nx+CXEchyzrq
PMrdTs9wq9qmqdirnplnzEI6BqGvuAZlvxcue75SeWZEuSWsMDMdAIKSXrYNANab
kSqWmJsZYeEgCUatfW6y63JPx8hE3y3PJ3usMQ8k367sThSLcoS7rW5NNpL1cmsm
uPW5u/cD9BNwskwgu5UCupVyuZsPowAI5xiMPbPz3UcMuZK1QkbskfxwkgllPIWs
U85MqdaytVxZglFOR7/i+ZOXjBK5llzx8JAyKGzC3GTIVHWfk4ANXUhJSME5GyMX
KeP7QEH6EoZlu0q4eviohIqcRn5zCvwbMt0sOxk4tzzUtZisdmGNeiUkIt2sXTYA
sMeCwxwLdV0G3N9M6gT1fQ==
`protect END_PROTECTED
