`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB7jeP8OrW8NRl7D24KJ315YcvY8Ictm81vG4X4fujjo
4ljSwLM05pqypO0xlDsDX7ncrMIHMSW98/vYj1aZhwrgrRrRNXAoBTfu4bVU7/2h
86xAOy8yVE5olmBPwuQUynqN6lOeeUgCoou/wQc7MMGpQFn4hqZz3+VeXJ087Dqx
2WZ1Tyv3IjdxrBE9tCz9i8q7makos357Dlj8FDHpEEi/LzO8L/NOukyyvpJj1zVx
Aa4U+gottQOUySrJk832eLiPad3INyALyglUFQaXXCyq+e1Q4JeKLu+2xVLU+o/m
lkrI5EXxb68U2pLhZfc9XqikrmjGacP4Jf3YchgyARkxnXpq3T24dupVxFwtOsk0
MsYMic5sCJ77+oJMHr9Qmh61gH9Aje159+hDaQ9RYbvtJZYWinpfrTS/VwxaGUOy
KOAkCU+Q1AEG1+pD2kSKwLpPc+Vsv06gfh7lnlHqbxP/wb0KOTpbhFECnPL1rNKn
zG1bDafRxLRo3NT/Zw1GbqBEYWLPH6earbwDqK5MyR/itVc6BHuY+G9r8SmH9D+j
d6XFlymfRI+CBbu9TKwhk5q4Hdfjoh81NyVlIw1VV10CUqJA/UlPQkdg15MjVXQD
IKccuAb3AVG+ozFWlac5BdzwiXdLnhIZ99x/obwHJC31U/cPeIS2xHbDUDmynz+8
mAPgUwnGXOahEg6S9e4SylyuMHc9QMdui+WW6d0oQO5tooPxAITJBj3Js1gLrYEh
fZZgdZe3qPaKrh+cWWLvUZDSWy+ESCe3AkKdPJKrhVK6STU/GE6jkMEEfvpORvPU
E0jJLyZi5AjgwhlGNNYwhZxYqmGFQyJgKnGVGMFot0LovDdx88vStQepBzHQfOa/
rL1inSrI6hkM63UyOr87uf0ZUzV2AAl0qucPAehsn+w=
`protect END_PROTECTED
