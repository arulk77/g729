`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
dEqZFXTWEN8fUChU3amGpW2V3enJm1hfaztIHeomI3nqGbNhfLg4DyAxFwZ1615R
d7yWRrCcWpVXqoSksgRec1jl3mSytEHpPhaQd7D45U5GA2JNVy/E7+6DqDfJSiiX
m9cEYkK3XFd+NhczYdnqkF8dL3Hi6lgrQQjZZjUoL38G+T4UsMqkiArlHPfVj+/D
`protect END_PROTECTED
