`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44yE6HDdIjQ+8IZ9wdJ3fyfv4qrWVhU+pBEjZYBeyKwR
LHcGBD5RBFVf+DZ+ZDgepSvq4i5A8gNtpfV5+V9YC8ySEICy2gDCp9yppWcPlocd
ZWtEH6sNSN/Cbjja+DrceIIxDbZUUfKlh+jzBmkFtP9dlXHY981uiMhAby3zJLoN
J8kDxu52JlluRedlu3Z24ZWab4IfglqwdAANvjIKMr7bK7FLHjinfHd9W1vDwOrD
KZXjQvfS3MmjmqDTcPs11vwke7KT5kZo8AHazvPkqbpnvSAhD2GXXiWydKj7f2kk
AZGjheAc8zUUuwZX9HkrQA==
`protect END_PROTECTED
