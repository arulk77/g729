`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45MBhcsCpA8AiFz5TAHeN5OmDQsbjAGX6UtzEtDljZjI
D7o17aeySPN4UzEabQlrLyoJ8Gw25QofCWM91L84f70Bl1OzRmfXMDwxpEdcjpUq
I9QBNR+dze85CINJZfgtSZcQIhGEpQd5yRMpHZI6cdmq77XyMYavfv18I0tgmqk2
ZLN1E1tM9NnfVF1LPRE6uKYWJCTtZuuaJ7bt5/UrBRUKjFxIfjZyijOtSNvV+iUy
5eTNriuMra0skD58Br530OO3dq4fCYodoyeD6/GLY0kL4DmBkpKR1R2XMbFIli6X
JoPa19zuaxwseCA2V/h6CtGhUwHMHvJeHmnAts8QMOLm7V9z9CCkflgNImnzOP2w
BPM025yMIuzTfizRdASV8g==
`protect END_PROTECTED
