`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEoHckXXNnHb73O17Yu7cpalCsGZWGGXPDduprTbuefz
aXuvgmjxn0YPq37OLAxcscR1xKgqsWeG9zQ9r2x+3E7bE1jTC+59NE0HrLs77Ui+
EmuYLhA/55Yow2GB/qY5Tg1xlstq2r0zan5LsH7GhuqbglKPn2drZqPoU757gysc
cq6lutzla5XERSue29FiFNXDYph2onvOeosX2O2Ou80OJSmouRxFP7Yjqeti6SqN
B003LLKCYSS4boVqWEr8BTG/4l8RfZjAkkamikf0Wdaa+ThC6PPf5fQbw/VbnXhq
ya6OLubDpzNu8MiBTYkS0WEtT9ZYZSfQggrv9Kh3jppmL1S7RcS+EhvFly6RECrO
`protect END_PROTECTED
