`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ5C9xgcPmgeIta48VvGenmazlMb75NhUf1G8Gf5OkVX
/2lbuRucB7aaDa6N7i8XINC0rx3ycekb1j/akmDr3EVI+E45SJLOTdcpe6eIiai4
e3J7RraqMcFdBZOJwGdn/C3QAc/etGPcZe3+SyITKiBAY69qLjNmH+wfAIU4NxRa
mbkYgQmHVjdWKZptiAwiByFDqXMhrqneNSAcixNy0EMM8uy5wIX1x76a3JSYzAgc
`protect END_PROTECTED
