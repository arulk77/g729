`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
O+yElpGCnZgqqY4af2hepId6B2ApxSw6YF512oEPPQFwmCWzVFP8OvYPqvcdzaU5
9EEq+L+7CNAM+9mhfpn9OLtJcu+41Dr1WT4Y561+CdXkQ6B1nFj0g867qeENgY3T
3ubvKpZjsPHelU0n0k0CLZ5cSPhfP8beRNSistItQTWeJH0lgLygzCO3mPfIYb/F
Kr62pKMu32mswHky2y+iYjvBsY3aDflg3KwAILMfe49t0PBp721fBSgdSCTgsDBe
wqAjogIU+XscCrwMzpTNsYmVBXAObap9f/ljhOO0bog=
`protect END_PROTECTED
