`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
VVK7x26ylIQ265w91kLC/0msWybGrtyCEzEP2UGISZDkRH2kEVaeYWh4srb0Uncf
8L3D2Z173cNIM4T6ghOq1EF6PjLk7g9P+JGURcdH68SsJndszHK0d5FqMq0mHWSF
caGum0R1ZEpKNGDYPiVh0B0BuedtQBXOBIH2+ZQwdUJtYt8YklNJRsJyCqpg3P2l
75w8tCpVTpSLJv70hM9Pu04fj/xXhQJM0NDsxMR+qdDx1vAmnZTiMMaXoV9wvish
Y1C4aQdOSFBN6J+dgg9uE87eb9Jt5OW0x/Eo4IlhRnrwxcp0IN1WOPWhsy6IlcL4
jGebkMjk3ZWfv3VLZ6i3yFqThHGpJCkFpkOqA58txLf+0wsqF3SS5Ddd33Js1ptO
Bg8M0eIiuXurUtUSDICoBRKe6/S9zZR4fEpQkU9euDl3kV/xtOLyREw6tMzKjaxJ
VnEpjzzO+MIkMrODDhSh6YfhthvXttTsos25kmZbhgE4OmbzM2vTABYiMywE7XGw
2V5Fb9OugbBAorZsFvKbPugpWkgRLl6ejIicU/EGAXY7S70wbK8knQTKflIT7SdB
uAYC3/wJuaDQssUoQEjA2XSkaBDQzfV4kyl7SknJmsCXbGGmwiX5KXn5J0DJEbtX
yN1MnxBXi9MsB0ZxYrnT6PfRHKIceWBo8R+7yFJ9GJRETLCtbcnYSzTBeHAGa0wV
I+5sOeC6ijXPRG2eZkW5oUm7T3Ec+/2zdk59vB6MINYaCJVw+UNNKjAp5dqx/kVK
SJJb9l0GC0WuUHh5UdxnN/Hps99AfDhSwWDFyKkJg9ExEZXoOVEOLJMF1RsDoaSF
lMAEnANXoD7uTDAAkerWtwRu6/SZXCBNn0/EhGWAYbj9yj0tHD6hygMScbJxTKoX
gPMKiqDn1QE6KeuZWy4L1ZWwcmvdIdTmakJ42FLdYxfnIUayRXPqsf0HQpUAlJLM
Cu3XYHaCMrjrQGe6DExBNKFqynDBsXg0vrTt8Se6sISUYkAh4aIOq04Obs5Xea3j
7Q1ecu2e74Vdi0IaB6ufhIzSkBz9Ik4onLSIiVnk7oU8GsiRxMK7NUfCG0Ly72mp
v8f6NnQmrEOde33diYlgLIerRvJ05zfRdN+ON0KfIIG88Rcqnn/e9rmduzRM9m61
W7qKKWE1zqssQPdI01CY8fFCyMTba+SVOi5gYGiBJ8fPvzz89CZtcCF0XMPHxHZr
Wn7M0pIYZH3nxv+3JNMh4XNkb8EeEwNLZ1uqXMuvvvl4a8btwXmpF0fVHhTukhcu
lU8j7SVJrchgp9lUh4v13AlkWCcRmJsLsZLLoNau2rJkxBrVY+tUSFd2WJubVimm
XpIb4AZim4v7jwnCtnwPQahxMZPY8b33WS4oumV6IySpWxmp/YD2AwZTudw/fHHs
1Md98cnyNBPjQfCh8mfwO/KI9hlRwxARBdEj2Q+3WEiHzn2IzizS1XwDDkvhRr84
j2gkS5JUg3dxEBQeE/tcIHyIdUjw8euqkrhkN5YV4gUssUvm8jg/MEAcSi9UWuUf
MsRb50IcxiJhuHoVBc+SCtgl9rMg5gJGZGkysCCUYyTCm7ziSuLhNxNTXVSv0RPE
sVXS/LJAtQ5dBXXtO+0RvLiVTe1Z2vIwVJ2FJTTyCKIpDJ1wGfj0Mzbf23kmSAwU
lvpGKpH1OteEEx9ukUCOMmxmid0u+PwnEBV5Zxg+rMZgCTd7WhEdIWKQ/FjSPv29
zdIGDMMGD9UHIVPv9Wl9EXqnqpV3BdEHno+W3IGbBF80nMZMnHNj0asUxV70VOtg
o0mEntCZqEK4HocKDA9IqI2pfvMd/ndBA6lgB/HKYPfl9Y9EDJAOPlzfPiKx9Z4v
qAGW2rCq4updjcahgrIhFQ==
`protect END_PROTECTED
