`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
YDZ5yQEEavcD2s2NsElQ7bJrUxxPNYpUjJ48y/0Iw1zKkAD2iSlF+D32x/dP4ZM3
BCzM8AaoQhHurG1bl2YYQm1gUL3m2aUSAo5OlBsrCeIPKJXFiW2RskPMHPdb6Zjp
3sNgiYKCV4tXsnjLOerGOUxVZFRLuoMh1A1bOEml1QqQTe+Z7RfmTs5WCblx5tzo
WxkQGI9xyPIz6evcjzgkAmwlViMIosxyQz3y/MCHcD8/kmUzy+7KXwQq6bYqKBmu
OP7WUFmBOemW5mbiD77bhIdze65K1QAgKT+JhWVAwbY=
`protect END_PROTECTED
