`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C/qGi7vmvw74SynNB28Nc7QKshEqoLgUhoxTxE3TTPGW
vMEklTMI+XMbAKsyrWMcNTQkH9pcVsz/hSsRs6MS8Te6/a49Hy4+E2NQiz+j09pt
BDLbHXAIFi4kh3Cbn8NhIQCFKeJUjrqXsNGj9jtzxs6Hjft/2T9f2UAdcs9q1NuZ
Dt59lijLl/O9mbeB4z3rIRLHv1l7R8CTBtVtNUCLgXCQyJp9hKF+AY5seHtRSUiS
S+52xgObPzaF3Yj0NEy81UUVOoAHosL7VxF3lhcWuQ6p8aPtiO/+0Kx39pc0iWv9
D+aLqtB5MnpxLb40B+faHGpu4ipr+YhJdO3Gl6yLLsWtQd6MF0z66U8bX5f0N2+W
RjPADkXNfmg5g/b1oSQ2IjOZM9QWUgQX8YyKz4bcXzaQNIiYh6gUMtk+W21ZDAad
yFq4wEv17aJEp8HSiQ/Ho7lOCOp2L8tiqOyaUycyraIi+QJ7AQ48BlqpN/ATJFau
gWgURcQeyG5Y+VvcGq1mbnm0aKdoE0B7IzwPeBVqPrehOhqqvwZCk8IWPwQnleAG
MPnVFalwucxB/GcGzMxkthsRCsEdESIig/KRknAPWRWFPa301sGQmNmEjXJ77IpX
P5CWgPY6CO7WiCuhqcwsd9GJAeX/sOIvJkSsSzrtYh8VAkCVKfU05yN1w8tmOSff
h1Z8aOOEq04I8TNrr9P4cDpGfqXEL9Ub/hJHSB334oAXCNjOvsHpdTlts/2U+maX
AYQXRyghKjOkF6CquWlO19HU59+OmbM97tEQ9AOJd6/9XUUnAlrdfcfbk5LbxegH
C50Tp+GIsk73w03NEKt7IPGihaZFp073+syK/sH7eT67PResfXIjuoLKRat+8/04
gxBkWWVvEYQDpvC4U+3DrYRGWe/fC/lIJKPKNNeY7LAH7Fs0cRSvQj538iuRk62F
MV/JW8bj1aAITquTZjiGoDI/X9Xt517j9ERsxwujF1fhl6tCWLiBPGBoIL/DWa9r
EdvmX0CWJPtd982EJxMslwhg4SJZ+Tf4nLZasonsn4QXmciQdlv6wdxZq+P4TIO6
5iSDBAmcRDl6TDasFAC+AUbsnZ80s3j3vwhTL8pnZANiKiwys3dxDfkYqxrku+b/
GYAqyiwduy3UOce3f7I+Lpn1u1dg6E7rEuLW3q/ZVpZJj8BvN5ahDrmWiSO2tKeb
E0mTB4vBkfYQtdUFJwv2CqxmEqDYsRejmMNDemRNLH3GU0xWsQfOK/1tHX4FFsjn
sUwaDCG8UucdORh8A1HIex9V2PJ6dAbTGFN3zddqLkP18cahn3ExQ0dPkC572RxU
PpNrRGCU1ZIab0zLHTb7qy62QmVrPP8WIvRZBG3PzKRNYDjfTkcIlm6qGCGDasXl
RYjm34kXrd+fSAqX/4kQ7lGwoczt0EjnJVqK3z5DeVjoHrNmQa4bJgXku0Nwi4qX
mVOqI7+VvVSjhhaCggxEVeW3e9t96tvH5we+HNDDMKlB7jrspQcj1fIuToAKt4Qm
PPfewH955m9L6Np/149t9WrDZuf3AH+dpBdb2AN8Ui+WG2TT03/KN7VR1HamHGwB
dTu+0v+93iRPjBBZ7cP+1MRH0q2fOJXefYrfzIa/bkhHhvHL9DhlX3S+f+SJxqHB
D3RHtMQh4KvvBJEJ57ffp6W4nysh5l5uXeyiD/28wXCWpWDSpMHJFK3AafTU3I2w
ATi2JfqYJ6wclgT1d02LBCHp8RAnU3/jmHCUEQwlrUpfc83pz/IAQMWqDv1F0/u3
IuHZ2bJ62uJq7IAU6flfVHIa6u1sYKpjUpwx5tbVC7qGGVA5BxJPbxLU0Phc9nv9
IfL0y0yMzzBcD/c8tcd1twHCnqy1ty411E9QMRmHGMq0a3hrmOrLWPm7EEsJLMbB
N9LXq3cLQZFAIBqloa1XW9SLkfwQCD0WYXqUri4psPs=
`protect END_PROTECTED
