`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAWr9XS6nPV0rEYpmFszj2K4bXc3d3wWArAcDBL1w/Oi5
oAIUuQHsXUbl2LyXkt/KWx5Hww4MkKtzUmomBfdf+S0VvJcjLJsAHFzd1mAcsqC1
EdzOt4F/mtcIJx8jyKi4nIbfNOqeheVsbJj21nsPfB5Z9ihZyl1itZ2dOQLd1aC1
QuHR8T3pU9ZopySOwVAosgRaqMqzR88/gPSE6kC+M65HBDZENrTxSYyzM6P7ve06
QliORq25GMNdQjbwJIn5t0i2bpTgu2vmdBYGRgOT0olKgxRe/PZOl3y6zMQyFo7t
d5+E48e58hhpHb+NtOrTvw1opQz/EFWVOaXoFOVgL4NfwwaQGZN8GZrFU7y26mqc
EmDqRoJ/lpl19bx9BIqIEPcJjtzfSga8QCN7FW8YJaVuxwMmoBwQkjEqLPtVxeVW
ZYyFu+glKzOTxim9as+G/wC/g05YKjGhtM2vaWhT/FEpDQK+qazyXKW91z617QaX
RWmtyGC+mP+OOzXrGqxQDdQGJjz/fLnAUUNiHL66Uzj7smDGazejI1vZBT7K8suv
1GWcpW920cTo1Y4+rW/j48poGZJEXojkN9VqENc+JO9pl6ZzKXpYSoH91i4ybmjl
3rqkDp/uI37MVK+yp6OIATVP8jOh5Y7iKe+9g2oWpyHZibVLn7BCfDNLnn3a/SV+
j4jUDdgTyTtkqC0hPRyx48Z1O2VxiIvOBW1eO6dnIvWanHOtNsgVK4qS1aN5w5p3
oaGHi9Kb7/PJV/tAVXCSn+OCRMo/gWU+XeZY1VDNtqo5dxYWMl4+k1aoAZ+wCt6x
y99hzaNVzcwamBK5Fy7LBS1tpyG3mSD+PgEiF8N8HvuUArydOqo2MM2Udq2oA+cS
RBPUL3x2fx6Z8s78T0yq02lQdKxI6OsoZ3KaXNRR+PUk7WETV8G2WMPxwTCD4DVu
zTax68hB1ITankcGXu81NuBujgfxtJcIIH5XrrPhb+34vgVqRSC0XYhLBx282aNt
uCZwXPUMMIo4XXnR26n9qaB3ZIlaVOPgKgjiNzsvM9FFbmPgji7aDRVrXAKBlfCJ
5eAhy/R/Ki8AkaKLngge3r9KhQUcvY2ZteqQ+0tt6fqtu61yG/aWe/bebSEDwWV0
TXHwEQS1DNkJD8dWN4L2AIVflXXCSp2FFpgTT8qBM8Rlgxg0t+TfRu/C0rqxcooc
aN9Zi5D2XYvxtYL7KbXdXedIQ2i5rDSJibjXa6iuSrRSl1EvB1m/eNbDY9Nq1Zwq
WBkvBjckwBCZCdjz8Ejf/guZ35BQCo5kSo3k6HOet/VmQkJCOjO+BpR0vbK8036f
SLZU1O9Is5FTT8g0MnA006mzslskj9V1t5ZhyjZKjbWEcRxLtAq1ap56xNxUtXMc
wXo+5LMB4OK1m++IiAAnG651vSs0lN0vsdeaa42MpmHQcVVEbGqnX2PmkWY6+BBm
mLtLgx6iu1h03MB/KECjf7M7E9rSRfYSd0D2+NoMDGDg16T5nfF+Uofal3v9AZY/
YfBC6At8cV1U71GeFUPmC60xclx/9nTmNrf3B0wge2ORhUrzHp+kjIPA2A8SFF9I
7daW3m2wcbZD6FuJk2XDsSDynucngZQb3mWT3lqUb866sdyP+JNC+rOEYO+z1XZa
7ObSnRx0+nFH/6ZsShdrkWlayijeEdgDr/AFcLZY4I93MNAkEbwQ9zgYTTVuSidK
sBIWVF2xeVsNMK6489tX1gHoiXyOB/wUR53O+E9oWDXhLf7YsCV7C+0O5D117zkH
V7HoBesvyrMs5arFf+iQEXT/4MGvCIo9GwJnq8N9Wj4XHeGd7Y+K2U53jZl14cKA
JXx9OqSIRlYNYLfEqK1RZ3KU5+hy2nhcDWlSPu0baZkSt9cTst3LaNuMu7NawCEO
qV+YOI0Az6eqULDjMbfoJ1iSR7c2NrxRGE7g/T85YDI86LC8RQUaYlo+5lsDeh2F
Fwh/KjGDYlAz5v6tO/Wmem+mclFPoZSMhosoQUqM7Us=
`protect END_PROTECTED
