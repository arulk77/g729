`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44PPQRQEiZmRihZNX7NzYifkw9gCvgZZYzxHJidop6EF
F9mWInmgv1H4i40IuBGfO+E80KeTIM1CHuc+DEKPPPZNxkuFWQKLRqTSwEhYGbcR
Kc/fUkZ54sRzQSkm7jFm3XG02zPETMKgv4UFZDtTHZLszWjT8Y5IAjYhPW8zC6DJ
Bkaae/Kv4M5zO6qJ41Xz2O7kouf4sjhwwqBIIDdovvw=
`protect END_PROTECTED
