`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI+b1j8Dwwo7iZM9GSL/AtYAqGA4PIQd+T/fWwE4tVXJ
100GTSCjnME62zZEf2JSZ8R4qmfTGoAMac4KFbOIYKlkEYDjEnhdWOSl3Q9Pfwo6
0NYCsWTzS/xM27BLCKct0epPqyQ3GllI8BzIVJZA798WfFhPfvf6xMDTmWgcIV2/
MxbvIUgwPi5yohB1stkopSNqEKx94FuXbKJvzEfR39Z7vAbW3Ug1UoM1XK85e7kK
HVPFWRa6VN+k2vFjvUqUX4OadWrThOT4EK7ugEVHHwEKT1M2qfHaFHFjwITD2Eu+
KQ41urmOtuiyNHtLJYKATw==
`protect END_PROTECTED
