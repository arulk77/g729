`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aeG9AW6Qk/WSFK3HtMRY/RiMiL0r0duG6Yf758dvm4RFqwtNJxBUa4vLsDHLmYXW
GqrWu4ueGhBLW8GezE3xstGenceqS3EOIB09UwmHr5x02fHl0d3DW9E1Wc4TyYPx
8Kk0k60yzBUnEfFZRUkNGkHNnCVgnuvB5J0NgUYxSNk3fW4Z5uWA32ajMECgAgsA
1vm9ER06iWsFbXQy5RUS/UOt6DeX/lCvfk4CQY5W5+NMZ43025QXfL650Qt1vym4
kSeUyrHgA6Zst3yj4RdKcw7Gn0MSZM+1gt7beJMbQPIQAp+jPWhs+eTVxuEMXsD8
07JInOkLFYTXlboaEFZ52ROhHtlut5PK4au1VP2gF2SzMNE9U0fw0RE2vw5DmRFa
IwOULdm8xbXfLdZYPT79IGi4906g1zpK9fWJvXi+gNmyum3P71rNeifrFiJUDv+6
QV43NlbmY+9VvkZ9u9uGIg==
`protect END_PROTECTED
