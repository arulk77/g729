`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDBM3MCqxVFLdI6I2DnQQRoxzIHHjwUnN5t7EBnHoT9n
IKfvFi6OtDc5hTeU3qhBYMev+cONC3f+aD6ezbGwyCQ/wl68k78VpXSrFnLpAv9K
XRc7GYPTIDUbr3p6xl80XYo6xEYJYstyzYl0tpksMtrxh+QEJBvSHQKkzT4Mobxk
NziV08bXHrtFdyOrxk11t7oglWQmaNw1AM5vg7g7fphnL86Z4Mr0ZZOLMmXWNxZX
7lfPqbYqFQNRMU9+ph/0zvPsaYQIodqOumek9o90Nm0iiZpZUxJP7DGH3q/UTdr8
Y6liN8LcOwg3HVCdsFPAaw==
`protect END_PROTECTED
