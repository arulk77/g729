`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SUHV5vQftxbEoG/Salb4BEdQJiq8XnMqWC5c+6r5wXwr
FDCWUZRYOgqaHlUeoAwbHtqChOIDrJn2awwnAoYo1446IqOVQAc0+P6mE6FHMkP+
rNyV2xspgtJcgupTK8rrHrHAojHMlwFCAC5vdt//mye7Zx5FHZxuZqFOzNB2aY1N
m9n89tFf9D7xI2Wj8I75PGf5oIo5ZTwwN77PNSDO1cfOSonMhaKEiLq3QThFo6kn
UPxHbWEZbbkIlVJu9FvFNhb854kjQtpaI3vJtjbOS0BWlzcRC/x8aU9GuBlS1thq
o2TIiH2xgPoizW36mHGJicoc2+SJJ5jjwZct8qlklh5DrfNZHxIaJCKv2cs0+qBC
GTB58KhqsPXYsU59ciyjHeFPLfs2lu9pYUougbmiEeFrB1K+QPvaFFk7BdtlJJMv
NAu0JnGN9h7r5hxIvBBSnoD4Ef8O79B+mePPBlync6sbKx05azZruoOgG+KB3Ejv
f9kTB38QO+WCw9ifR9SW2o8O6MfrrnhOm0EoAFSdqPNGRw9ed0ZnHDLsUSing9h2
0tYdHSC0Tr6djMMjYBDCllCMxEAIFSnV+AdTPf23k7VGPDSaKMtgL8Yl9XZ9nqFl
cSewbkML8nqRQkVGDJvUEI2nUfyvYl4qqJdAkKJxb2TER4D9AlSDUyDVAnkne5CI
XdG+8xoj9sQK+ZkvBwy0e3NJlg76E6HGm8bOMT6gVApJn0gi5dnvO+Fbwb9siWvF
ZwcyWQmDSisbhZ8E9DeLkPStu53WPWTcfvYQU+90lZFfaYzWck2Vg655tGYVXtLz
ZT4GxAc5cudDVLUJxkWP9nqOlTqkMg4DCO6vegykvg3SauFvOnNW/HsQpCQu1e7v
ebC8GquOMGzfhVPl+xC4qZBGrWLwYN6YulEO48Ze1a+paOkfQIlC4XrsVv/4SszV
ZNUPXUtfav91ADSLOzzEH0iarnN1zCRd/1xOB+cJhYlV8Rek2aG3zQDlkGXCDth5
LOf7GOiElcghOyAFW8f92II8QpDqxEx+HtutxTJUNLB7Fb13+FeNuN9NWuWSB/+J
T2E9Pe4LIpclWDMjaHic0MhPdnrqfjHKUXjuuiZn8JblgM54CJA3akMTu0EVVIzc
I8uSygaTgYU2xFc62yNdwpmBzYI7beC/YDjp6JWPwMPWK45kZGPUVAwjlGFrDkUo
/2bNIzb3sKLd/5tKPsehi3pP/SMF5c1uZ/Z+xgozdhu8nMxuMYXYqbkpz6CAzShT
F9SOs7R778ElVZVKuEjKc9ylI/iYwvdY4hx3uMf4bxZXkSZ0vqmGFR4GSUvpv8HF
kwt+YweVlD3b1R9qCv5eXZGTr/OMa3+VO31fL/Lx8LNtckyovEqH2C5MRIUxlJLf
dUPnyEkTcPmMP08Xmvanwd5g0ABJiXTR2NsbtP2bbtNKQ/IIqTJzl5JVLAqLopYM
TP2+JJfETuiNbyRERBMJnz8r6whIq2b7id+Dmtv2hWeV8uj1k7WJ8EuF6sMwW8nZ
BXH91P0cTdTN6In43f78dCBGHb1u4ASQtrZjKlZlhXN7Z7esqVpUqhYYoS3LILmw
18dS7baASyZP5V2utHd3wNg6Ez7mmzeK1bcEL4C5kKl1p6MBwwiIwQh1ab2BPm1j
cZk0KsWTkuYY89ohPVhz08B8G4j5fpXSl5mKjJYUjXE=
`protect END_PROTECTED
