`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
uxqkUqUSjJgau4ensR5nmfJnLVxbSp2C1tsr624aN7Aeln6ebJPtuUKoERwYxHtd
LRxVB+qANW+k6KifoXjcFhLsSfq/WxNDNZo+ZkeKGaB2Xopzi06ovtKvC9VDZjjX
GC52KJeIzNlZp0s3yk1WcAPliEaChEsisfubJfUp+9OCA0k9kjCKsB4y4GKOxUt4
Lt1LlfBIHrRAATrjUf1Xj+ww0SvD/jQ/6uJIEP3EjMoP3xnU4VXsGCk/UQ8SFVel
qMifUnK4MlIBBHK873FxGtWiWqzrUAw2Z98Lj0JSL2g=
`protect END_PROTECTED
