`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
oInHZR+RfKworsitBWKNz9n3yJD66QCHZqi4wPdUTEyMbQSDOPGt7hU8g27E8bT1
1eXZf9E4gygsYcSxUFQxNV6H4yItPdL5WoPLLvf8WJiSJOEA6g6ioeTR1AeYlJ03
Lj2qhd+ihsk7NX9rJT4XHcywl4aJbQj6n5xU7k4ja8oR3E4tco9/wW4ZIOgbQOTi
x+X8p+OQwqgUHkZQLv0nQdI0W3N5011X/KvXRyv4vBxI/CFsImJ6dZSSILce3qjV
AFVUC75tOJMISFVFwNAHdnngM4GqjkE4+yNRhPBLEbb7MB1ZxiF4pLtYRfK/Dxyr
p3+oDXqEqIeNvuogxqvCpKs9Ubk9o9AtoWOU9neljTFbT5+LFzTZNxNo1In40pG+
PtEbs2DOLdljm5y0RImLd5RL80D4Honufrtqv6GJMQctyCyfYQo+6UGo2Ug3xOwg
8z6LUm1Jp4H7756Lzs5PqA==
`protect END_PROTECTED
