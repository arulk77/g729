`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN6qEAwfOrrez0FKPoal9XNRPGKdm+dMiz01lBtd6ix9h
I50z6Z1qNraEG3PSXm7VQstqBYcMqrqSq6pd2e/jgLuoHNh/E0iCkBn6bvbxCuBN
8Zw6Y2QzeNs3s65Z5pfaw6ihVAGcfT+xbOKKGaNih8y9MExGPx2ua0hBkiMKg5E4
VkR3BA8wKoWsORg+L1/8F6QSj5nO0fa7IcBpi8To1qcRvlc0WE9e/foEy/JAGFHj
NdQIDUHXURAHPtDOJtDYLrLCv8KWWFonlUDpt7jZSXVeIXfszMrcpU5pp7mKcQWn
bmfdH+fyprmeU8vjz00vxWimMg4uHC7BJI0Iv4vFIezSSwcE29Z6bvUSbfg2sboz
JyS6IovVAU0fYyDMwlloJMyqLovAU/Uu38cBzFEYMyRBb868YwcrSPiPoYtQ63fQ
r+SdRYalUuaAgw49p8SjJo9BQIt7FEVMCCHocYSjKmgHXAeUJJ/m+UZaGi8P8xM/
p+B73yHyA0NBS62aN76H+LWKqPfTGUoUbxSAzPKgzZBiJ50ZgS2yvRkZwSdcUdUy
4Uap2ST+JpoFO+1nm61xX+qUaXNXGOwH4dZJx327ROSuLDMmDf6xp7bRFgKO9w/a
LRAO2rEMZfO/X79UhzoNWYoGC1aFBNFlbrtTFrCEsCR04ZemrEotJAiTICzH+Z0O
xcVQQ6sKvjz8+ru1R80UA94sjc+2dLMPDp7Uwamfz+I5ct46456kPugiaDKCXdNJ
`protect END_PROTECTED
