`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
jGSxwPhLdDLT/sj7bYkebWRRFfvE8GGT0Dw4GfM7V+iZNbAaO3Ri9SDNcW8rYvZh
rtx+G9sghS3lnKdfurJR8UEAZfjHWcOMozEH3E8nJFF7rnKdqfNjQJPIGAzwYxmi
bBqwEO9kg67SqA1H1VME1XpCPPmNs4Fhqhzgqbj3fZMXjytbkt8K/QUm0I5atg82
wnTEt5LskW+9PfIbNN9UpCldJeV0f9VKXoNDF7Ea83pNZX5fKCk5lwdtAc43amB4
mTbUEtvRJDIUYGG4RJtwQ/DBIF031eNWGnW/OaVWmNg5PLZM+eITk8IwL2GPCOft
PYeZBgSvC3hP8vrdPgkbsBJRT8mVu50bzaMJT6G7nPA=
`protect END_PROTECTED
