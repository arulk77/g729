`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCIj+mJsftdo2yalNNFYhsbe5kJ5Lit62G0ALD4Kfs3B
vnfFmTfS4wOLCrmCGJ00o0ay6xYKAF++LJJLaTP9eBy/yIL4ltxuC+UifhhjYGub
A3Y2eXQzmM3ZcEv8WGFVjCN1aajY2gQfzD+6vanA9yzTWotnu8D5w8zp9SSqshTG
mlpTve69kgDteNXVrJdLOAvuKcpeGXJuvc0j2rZhlicpBv2A4ZagoMcnqMizI4MQ
j5ZVGRBg+UPB2Yx13PE8T+K0cU6Gm9+W6LPb0tICXV84Fvu26WRt7eA0moMq5Bui
9RnKVvdNtXZIR4NIznpswA==
`protect END_PROTECTED
