`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIMJSmjqDtDXxmMIj6sxYbXMbFXAAs03giiqNs8z+83s
6FBJvpdN4A6J0jCB/83BXq9eohBa1LAT4F4xV3UXXnQv31HRleiVzK7r1JX+AvEm
d6O3s8YMLYqSPMTc/G0tsGWlKN8dI9L7cd5P6eZ5C1be+Qqr3IidCje5mOEoQs2W
`protect END_PROTECTED
