`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAcyEg83Gvt1ipowubSP7ji7GOom2qacK1CNtUUxUydSr
bQ4o5BsHL8AcPOb+nXZ0PovUqi2pzXkVFOBgRSUrrLWrJm4vePyoN8FdFW5X6nwc
JMDjQpvi+/a7KzmO34k/OtCINYFgxl9c1ikYzeEPzV8DM1YVmGm8jU02aI5nBz4e
hVYAxZGh7YLasgIlnTMJKK6BBhOCDLbJRyIEJ2L7lOqFlHMikO1/hBqLd+WkQbkZ
lura4bgaoM8Fh2whuI2Vd9832TnYxYrZ+5KwJRvw+Bh0pzXcKHXeFFOynSfV8nhe
OD2NSOXSz7+BLiOED1xPQwpsnytgLEeJ6dcrPFAUCj9mECX/QhmBCdu1C0iR/olL
l1ykIoNsPiMLWIhwyJ9bqOOXOuLvzUNREBZlrkUzd3k1XKdsbu+05wCyeDOdwg9h
CxU88e6dLegYeDUihcNjqL51tZLDA6R8g+WNzveE1l0YDCKB8lWM/lVMpPPAJOJn
53wHcM1ZFzhWcWwQP7h+oRdWaqg9kvN8noqstXpi36bnuqBNoBcaULPSpdKdDxDl
B1nmtMNUdN1Mr0L9lq5X/dT9NnXJa3Uzn2+DEMq6quTSxXblHwKPJuPffr1tSidf
7douSjXZaAfUl5AjyGDdTUYKKsmzThMb0PeWY4s4b7cOz7yXRQYp7zHn+Ctnf0tF
GyDT7/jZJMOiXv5Ozwszcos48bvGCEQEj8GugdAphRssNoj9dTqZgfnq9iAzcKOR
64o4dqwoaqAYNeKg2YRnQ222TKPAumH0gqvbQYj64vM+bQM1GRugUienkJAKHO1V
RRQby/a484IweGh+qkvZs5YlG7fi5zDhW8ZkIqF1A28T8O9X2LnGmjEeX6QKnhvT
EZo8sMd5jbsYPGHKTv6ReBXOh/yZYFxgtsml3dQ+bbN2uPrPyIAcIF5smdUBUP+r
9IzATMqQiq8xmsV0kiMraQtw8O0NYfAzrsP9XbOiZm9ST7uD2CMXrMy3byPI+VMd
1RgJeo3/gM+gUFus3l5TGH5Xfur1vKFUzdwJJmgIN+NGPVfwq6ar8GzlYImg0lYF
ETA5x2tFWNWlo8SaVzNYYVA7Qv6SUK2EHzOD/YPyyTDI8HSYPPqe9PJZkJxZTIj9
oeqbBgaTq6mHLS4yYkF3RG1fQFGpjfXsZuccYlYIFELg0OCyXSmONzGm3Lfq57X1
4xhkN+fcz19a3xGWaunVZbK7B3euVyfNlJo1mpnfiW13mQSjXCgYWYeA/sHnlRS6
aAHKzVS46T/BZoBvPuXsNaBXbnhqkQbvcjvD/pXNuA2Wa7gJS/0GF8/nqAGrZg4g
E2NUefY3hw8RMjaJHLkUYDoRX8eoLRV4XPLqVF2HeOYjJ1GcvYdgaToqZVv4knLu
YiXeVUca96cI3rz8UL37weeMUzqaCAVk5QdSeWvEvM9sKT6eA+iD/ES4lex+JMCa
qr0I0/GO2y+WOC3hsnDv4iWXxsEyuEtObrNO0kbmgwAbT8oM2WHoe3EB5p6LAvcd
aXsm8YpMFrwMh0ntHN5Q+yQG+JdldBlwalaYAUwdO7zosz8vLXj9FPNW5SdgG2IO
jIFkfMIVysBZECuRjj/8uqhxGSLwe/f3LtOj4FRN4kbAdDYX8uDnWVt+/VdpUd/U
5H1Yp52+UEkzdOokwbyqoGKw9tfu0jSU44GDaBy5CldeIs1DcHJkMcRo0LOz65w+
5D3eu1JWzo5hlOypXHmStos3kbOhSbToWlnbwri/IjdZP1mfE7UGB6V+5avz5X2f
ansO2E72yo0nQeHmzb+U/cLYZ3c9TGCii9bC5DTB0VIlrGX6iQPKzOckUVlpKuaf
fGiNrZ6fgTzu4uFz6usf0j/zJVSf14AS0XSYfxFcQBL17DjYDAq7G1rlydIhOZVm
BW5rIzD6OYU2upLBDdoHA+sYnrFHzxvGuvVMfElxc2dKtIuZ+WPLoVhcTpyKDdK2
jhDABEQ5Mw+k3DnF4F1BoA==
`protect END_PROTECTED
