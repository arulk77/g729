`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
jM5/OLm3yhKobSc7vli9NdGs4UJy+fj+KFug4+4TBjKTRIGEVexxhRkWIRpuiUkK
KPYmX0emO1OMcCL+9PhU3s4zm1+hWoolEE1P652UwgiMiPLa6QorCWP4UOtpMyBK
W8mlByolV+5THXah8fEo4NO5wagRDr+PHzswkrkroxJS/wIsGLJmTRZltXd31pBI
RAM0FjeWPcuNeV1SIrxnE5lXwXmcAfhOAZB87nrvDtSj8lTLBtRMm+72+MfPuUsn
XyIMjZN+fVSieXiaAH30AlXjN3ep5YL1DGzUcSCg2XY=
`protect END_PROTECTED
