`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLhbNfOkOXIMoqmdfLrd+/9Hpgr1ysVd40KZ3w81mpnt
HbJwqD8nVvJ2VJFNpV9skwuIfUazxrcILccw2MvuR2Yu8T3dN4F0yuTlGaWXjLhc
NRIgtWbt81w91BEQ8fXieG2o08kfOFACk1otmNEJDGAJUm3a5JBW7N89o97zRzXA
d9vnX5rs3NpDTvbeoH+OhBzL2gQ6KN6tXwC/vlQGodVDM/YkibZxTkwlR812zYqR
6YEx4tQkjflyd4LQZQOUYyQEGrNDSlNC2aOITcT2z9nT8HEjZhZv/ZiOOMh6NZZU
97H3qKvjqurjgoG3F7m/mmykmbuKtJyoh+qi5j8ckWGPyC7t4WSR85O5RZm1Z2Es
s9ImLQ51h5naFrvGoK1HZA==
`protect END_PROTECTED
