`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAPKkHkyndDNT0F1Fe+jAN2Eji6bBN30A7TnBzrMbzsW
Z7GRDFbpPPUvGbf1Do3D6sbQ1MaT+NzlGImSYDwUUBHdpi9pj34VyPQWvoInAUVP
4FwsTLfXcUnZvOZCShn+voApOO8+fbLAREPjkAx6cACyAN+JeLghUoa6rx172GXH
BzyxybwmiJ0VnyUky/KosA==
`protect END_PROTECTED
