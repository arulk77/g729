`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
1u9KesXRNxHcA/V6oF/b3mzk85LmqEMrfBelbpku1NI6euV4zqsTt+DEtCaH4z77
SvDWOBwykimtxBSVPv4Cix3lHA3xmhAwRa9s5ZQHVDGi/3vYREcOHuKaOKd1kjMO
8VQzeThFA+KpeI4nCZN9ziol7u9Q1lUNU1mAaK+3Xa+ld1lSju9AqvtyR9HyBY5a
QXQb5RIbmyo6MSfgrX9O74furreTu3ZP4pDAsoMnjyhIGhgnsZqjZ6dS/v4S+SRu
qgJp8E4TGym0Pq0tCfJOE6RiWLLAKtqPv2MflWg5ReNV/FOOxyfOxHb35aKRIWmr
VkqYPFg9lyrp2ifNN/pRKpM21HJ5v5Mj6y9+HQqbLw4=
`protect END_PROTECTED
