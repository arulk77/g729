`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePCoqMfuqMS0fp8Xg/9+Sm99+s9AXwCiDY8/G6hut4vn
k3mtglsKxCd8tsjvz68YB7XCas7jAbVWKMw8VHqMKOCHFII3RMQs8C0Z9LPO7T92
yfhAN5pHnZhFQMWTs1plLaJC4T/xeflioQ8jXQDrR6PDvy3aCptM/6JVjQWA+ika
3IfGZzcHMbgJQjj5Xvq1b8bl51iJKvrFBvg+G++CECkLBEb8kmZ9rsu16WJNSDO7
wOprLwW29W0kEa8n2uiywfdbSfjdX7l4si34CfTpXWlhZaVtjSfh1A1jLvZFFBPT
izoOl5TcTuX3pl+s7c59PwapQfnP2J8t3Qqqm2s5Zzu9ZFHmRnlm8JNVlZsfLetr
pfIoBj1Oivt74mdrT0rKSEYbMKKDEWHeDxQX10NNLE+nxgZY/4LOo0nArETtrYik
`protect END_PROTECTED
