`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bh34MYDvuNg8L2FnQCtSDfHh+8/6zMd1BG/S2yFZiX+hv6Cr+H60KMKOe0q94Nii
W3apB0UpmrkWYpgxZ++PSPd9GtfGl2AvxcHMZAjWzjReGYmZtkwP1tcXQpDyIcm9
BLpBP2RrAgJ4xGEkLCh2GHayLK29E9rY2rnfVlBXsvnCxY72ZIT76EpFBNhsCxuc
cieH7+Me50zeBgg9MuWlh2K1taMTNLCJAufm/xcRwXlQwrHQFHpWR9HnQQClohRK
kTb4YwfmS+Zuv8wJR4ZIDEKaly7VSsADLx6lYMITIAgm7noItyp8AMRk1QsNNxFF
/0SmzIo2mnpHDxjOGKcmuR/7MzV89H8gfsx/lQtSfdc=
`protect END_PROTECTED
