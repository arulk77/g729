`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mlFBzCyNIVABC0bhYTMiK0vai+iO/XbjBVIeVpQa82j40G+y9xoZaVwx/eDuy2ei
BkG3b0+Szwq/bxG21cfbmuxyapxqheUO5AQfCxjYwkXz/VlIs7URb9DhVxoI03Bn
A83wo/3sqnJndy6HAKAHXhHSz/AUq5sZu8Uu87TXxNMogdMEpLMnW1k5eKpdBzq0
G2EdBGfkYG5Fdjg4Pan8FXtbhLIzb5oMyFREyGscg9BU7hi3AsgjSlBoLhP44yS6
`protect END_PROTECTED
