`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkTQVZws21HaWqi00rB014ioO8kMrW/pXT6qziptpFvlI
hf78fW+k+11Yz6Z8eorFdnqZi5V1saY6viZZ7DuzOxQ1qcVd+EX5AtNs6Vh+jh+P
w4GvgKoh/yxp5MoFE1IJdHbXTejAoWKO4fC9E5T1pgLr5KbuNomZWoCDueCFTHC+
uxkYoMK5u585an2op3lnG0GQkntrsn/5ie3frqg8NZ4cJ0g59/FqxmDccYXYck1u
DNmA3BpJEkuGdjSi13zfoooopUnMbuKLgtWXXpN1HgQkCdvdIl2KSiqUq/RIdR5a
bB1IL1qStwbEDKhwAteT4j+/951lF1/JOghXOnvUy9Ue9nNjKgQOUuZHD0+dHmfo
CacEAjf5kpBdIrTkBGWIi6GaHZOOHJyYfRUX1vOcV2ulqs0w6OcbkGLJq2uhRDR9
0x8SJbV3qGnSbHCp4bW2gg==
`protect END_PROTECTED
