`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42m6zLA91fhcqUpIZwK91tC6d4hlKvFNjse5Bxt+RYRV
TnKzn6FETApa0e0fDUw5iz3u54qRY4NyjjAd2lZneOZPUqAvqrERGi2AlKUF0iwP
pkmeW6FgxCE6xzd4JynMbtBanRQHY+J35lEI6AIeydZxQjMNP20yh5ElOoD6lf6p
U6Ev4ivKTunPVKbiyspuDbqdeHhOJ+XQ/fYJoQpN3b4NM8Wu6rfyhUg4ZGY1Y0qz
MgsPSBAMZDV23BuNysMncQqlDKqRSBemQGV+BnUbIu0=
`protect END_PROTECTED
