`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41ZXbX44ZGIvpOWKG8C68thunUITlWjwyBsR0/4V3/yw
UyrUNA+UbuqoMaIr10PmO57pBldD2mS6kZXANdt+ebdKympy0NCKP85P+E3sv9VM
JAMoFz9WAFTaKsqTsmqOpPRRM9QLT/zABrrdtNk0v2t4RZvtP0lpvJi+C59nOtIQ
pON5pof5kr71tq7Osgj3XnNcu/ovGw9iNVZdCV9cOFPC3cCDEcCzn0pOEgGzzypy
DnKMCAfgw0wk5IElGGgv0V/woBLrj3JX1u/BWwd7Ank=
`protect END_PROTECTED
