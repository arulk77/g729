`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42Kl+eUKqDmCe35dZd2aYBrf55Zx6Z01aMTUptVmXALD
OKlrt8JokQ+2P0k4I/CHl1ddLiq8R6u/nsF10MvsgecLs9kS4djekG9ZhRsYJLXq
mAwdI6tmw2sAC8SZvLLW+Q99jL9HDwP68gMs0ns1Rm0zA5VlvpiZiz5r0KQSAFZM
hKQUNPf85N8c85SOvITqqK8MNnqkc/8BFZ/B81cbernMhsOVd9lRoQtQi/JVG9Qh
K9++MUS8OOSJrG7ptZ6g6UQcQFGY5RVqVFmDwFiTa2G+sj49Yzr/TVStkBuzq8ry
ImsoBgo/lNXSzGKJJdIMIqHgrO4DdD5tzRxWEfmHVK0EuvTslSNrOmCyCmaK5Dtl
VgjGgR5ExS3lFVYjkNOoZg==
`protect END_PROTECTED
