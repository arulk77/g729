`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43zoUhnlctk55Hn1xsHgRDfouKaX2ZQ4ZPPLoO4kpY5A
S7fX3KtkcIl7m4lsskJ0iWhb8VHO2PMWp1/V0r5IV5DYOi1s0j8yWr690CAYVdTh
EdWk4SybKfgUGpsFkVLFMGFR+eEacMKfYgaqCmfoQQ5JjJpky9siwVTZIXVotKdT
G80+9pShSZXOatJoHKiqEtXIBERgh2AUn7QrYDHMm0sj+2AopCRC8H0TPskJxShq
1hpFhQ3S0A3z7SqM3noCD8h+EvmUsHtrz+XCshXEma4NlR//OdfNwf2BWi8fQsRl
Ml1kSyT6MTo8tVdogKVdPCbEXvPHwMtLbJruImhOPQyGI+0EjXgRdox7Qc/L2Q4v
ChgK02ENSW0JR21PPd7psf/8YLI8Qai1UBqXBlsmMsqNmCSTcko+VWoa9LsJS8SA
382T2jyIKOs3Cp8Or4xHYw==
`protect END_PROTECTED
