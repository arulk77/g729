`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4776XX90NugHrP6ciWnLKpoQaCq5MqpDRPSMxP26DzAX
8cA1QvVV50BHST8gQG1q0fKNkYNqofRVzSY4D5JtfSHvmtd7uSAdf8d6/dBgRDI3
a0uuM0rSO1dYPuCMcgLnCa4ZAjPGfTivN3FNAXFbw41JYLtmV39rmEX348VUARM9
hUeLuHxKG20wv4kyhilWneuIAAIQ5dBcRSOYtFq4wA1DXh60O4VtzWqz5igbQgTc
0FAC5z5HU8URpvANbJGT26XwHZfkNsbNmU0RBgdZoNblCHrPpRUHyySVFrok4LS3
sk++R5B2Ft834uZIablFc5BoHeMbimL5MVGTbZwf7phxk3J2U7O/ndmf3i59pVnA
eIJPVWEK71h5cLp9Um4gjA==
`protect END_PROTECTED
