`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEwAzvjBo9Y5lWlZInoaQmER8har8eE4d3N8cHJpvgnI
rDxJp0p5aKo2p40Qszyhd7fJRNhaurNawANUFsmGQdc69iTIR+RGke2YlNZNnZW/
A5THGpsdWcy6jXE4GUlURpJK8nEsAoMm20aQlYpCDTT5jbGvf1vxv86HWqsOzfmX
bTit8v0sda19WFr5LiMp2g==
`protect END_PROTECTED
