`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
VN3cZiJB9f6xREOOK65F2i99jSzsqlfzdmFj4/Vm5aDWrvoJFRBBaySeODl6RpU6
LLmdkq19558OrbgnMTbg9UgBe7FnIF/gNGCKwO5aiTJdzuisOOBRsBD+fSAz5C0Y
+1vA1QFajNMZ64UY3J15oAL/pw4MdW8fvoCX9RVeGHFDYkkVfqazio7ZrPSc4TMt
6fWSwmhZqaL6T50055sLPvA2/xuP1wQChCFZ6UyHtnQ=
`protect END_PROTECTED
