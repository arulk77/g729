`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN7TQzQVtogJ++aAnCp6HAnoOFa8DKvDNnqCe56mweAgS
batpoDHARmjPmkjHyYaZjO12tKcb/nPxxwNQ/8FUmIf6BF4VEqbYnYb+q2CQQ39u
hBrLt7xDGkGNIi5uuuB207lzRGAPAQ0NQ20NakHdHmu1c7tcceBHZtNzY6z5+tKc
Zv/PIKSfD57suF8yHWAop7Myi9t8z/u0kN+F2F/nnST6I/OJ29EbblZCaBaee+XO
EMnJb2qhqPceK0dv5I9aK2Ab/3NFCIqrx4GBSqEPQWws+//jP6hnSVviBKj4laD0
hkjrf3bSwtoQ/YgrAYuRfej2I8S1B9LU/hl08Yepz7M43GU3aC5mgdUq2jBGD1eW
hHdgFh91r40B0/zZCugKrUhGVOuyA+PgzU3BcBCrJI15AfSmSoghmfyvkrKH0F26
P8fgDNQS4eKiIvxUw49mG0nR/RuU/5phBA6yfjiay4n6A42KYgpo5uOxMYA/TgNP
YRyDc2Y9FJI8na/w5ov+NHtkQRb+LCki2R91mV4SwihREjaxfBCBugDDYvay4VIY
+ooq8JwctSPffKzjgBVJ3J4jNbmDZ4bD5HG+eIOf99Ovtmg4xuHfTctpQ8n2b5rA
/xjcZg0HDt0twmNRQBb7HWHimXW48hf307Qs970QiNL+ko0SJNWS07un6aKpN3cl
eW1qiYUm4EH6XK/MToyKshuz5QH1GeD+33StYTXUyMehPty9j20tlHkw1aOA4fCy
aEEoGttJunStTQGHVSBWEHLgOFdPEU/89UwajqSGilXZlJO47Xp/iAqY5o0WA1eV
Lo6ClD1o7D9RWWdzy33oHSLeenom+6pUIuuL/v9znr5VcIclfyy3SStC3CRA2G+a
YRO90/wYtsU9mXe2RDgHLTUUc00Dl5EMXc6TIY37iyEHthQj6IpbK+o8wCHxWZeC
DRACHKv2/5KpvLqihLuPnoo91wiO1+dnjBSvRvSKKCgGn/XqCq5TgQjwMHs6AeUg
IiPXYFuHXOduOAxzSQonA1J2LSPEep7Cx5f1SxTt+cDNSdK128zxflS/RFvrpC48
mqpob5EHVqwt2eUSXTBMIoLYTXz6hPrgH7bjYuAzHwP4Ux3oP88DcHuc/VzLMLFm
bCRUpAEI0JSzZuVWpQ4h0Sq7ctn8GolLTVryp7g3sg1bGwR7JJtpZzr/clGePi5G
hPYa5h0xzxp51P7eX8TI8UXmB0BjEcTBsEHe6MsLu9xhBFKybfu9cztt7A+sYLqq
Bm42CHdRBMFGQPYDhr8fyYxUnVdz9FkM8ipCakP4q2eKN7mjRMW/Dk0BbB+AjsdR
8uueLuHmmv1N/uYo/yIOQGBe/Xjg1obbfN4R8vd777JUrYjTt0R/KOB4zCJkMOGh
3lZ+WOzVdeLtfjYum3yDPqmUXluV7tijBrf9TWA1rCD9gZUG+e5VcaJ4mX5O3HVT
jo+k1/zvDrv4b1ZzJKnnQVoyW5aUYXFrjTDew6yte5sENj6gd+otJJ4CDwzQECYP
cSVzgV04D4ks+G5hl/BcxE8GPTwUrbkEIsGLBW+YbosMukexqLRKFhZSXDFFLFkX
sbwvTvjr+imE9Iw2reO6yacUe3hD86hsLImfLgxqz6PRvqCydKo1DeQUuvdCUl+M
UQvEvb4tFSVC6u5KQlEjZTFmgYPpj8oRrh7JMzx0KXUO7PNi1ITDlKzW+bgMdcYr
55nDvzSU94pYIHxySCxoxiJ/aOdslfYcpVJVBJrkZnyEkfUEyTxNr28/G9PyPUCs
PjIe01BoWvo1Egfh63bG6ZsNKQPucsfwVqY/e/Po5hf1C7FF8oN2bOLRnYkLy8zN
DjwvrcFGvpGUGtHI8UrDHELDABSO6a4v+avjEPKb3DiDyyVzhe5fRUDPZXQ006IP
sVVQ5ocmRNxa7P6WuWWfNZotUxbAuehylFzFY6efOUbM9yJRX0vdmtGOpSiQjVYF
fvzpvDhwtDe+reYbEU5XupQLYC/CSYvur0IfuUXWHwvUPz1jX0VXn+7WRr9jEoCv
3Pb8MMB143EU2LzM9kYdTBlgeMq98tmsdDNspHDAA79xK9zD6Cz0qiiKC1S/108D
N1clF2KgLSdeRMqVd69xz1qSfOwZmWcdBz4LNe6ZCRvsmohTggL3XxQxeEpoDbye
/dFkq/82vB18V9y+POF22XDlk0srQI7u3rUWB13jFP9wdzF2uJ2g2CZxPH0crLmu
q6tt1klORkcGjR0NfA4gLqFNPgpGBeKj9zF8icjAAbZGmTmRH0Hq7pelIWc8uU3S
0PKAER7ffXSyqtnj2qHuA/8PDHSYKcGLEcJcwXcupfZV33c7sLVS3cSaIfRcNCjh
Zb8VPZc8ngku8slI+iN26tSnx6CHlWikXrJB6/vf2dgQGCZeLjqEnCvSF4/1eEG7
ZxQ/JE/+S6ONZkVb8QGQh+dwX3u5b/RulsmD1ZN5tITPApD0Du5hvWC132vsk8sW
KJJta9Ed5gOc3BykCN9uykLpPZW2q11xf5/ECb7Ej9n3PYdmwwgzP3bAaGmMZL1g
6ihbmAogppEN6eILcXrxNyVbRy1HWbP1iiJamYazPQkaKI8qM4pN3jpma8zHM6ir
7BXXJo0kxKl4m3VwKOuvEE4U2jWS6ie6eYYDQixi3QqocuoZr111QK+N1QVjwES4
0pxqbNMImXHTdpYrmQx7IB7GybQGlkfIMl3wooarz2LEFkF/zkWdaEyRLwFouvih
mpsBWdrhjWycD04aJ9kdskQTKPmn6pA5bxGvltJijiA6VdpHVZy5+gOms2q4utoA
mxa9zWmy7nGoqg+Prup9RL0JELckR2O9vYeXPBZUeGRUC+umzR5zetnYQZieo38K
Wb83d0hxALNqJScJ/ORsh0W2E+hRsMIK4gZCeSECm8yP84fymnFuypoT00qye3Ay
Gc6250/eeiGrOzh7ijgDiXbjBNlO6l9uZZv48So6fcEV1KDZZmloayV8V1fKjrsi
O2CZcdeE8muIR66jiZpNKpdz3n21Pqfp2Il81/mkDfn5IY7Qp8DOoo7kDQCI7Q68
MHgEO8QqJhUKwShvJNZ6udok53FcRnbd1qkTofKsvtnRFcmamhseHEDjxzXAA2gB
lmEs7HwL08G+ML3qPlhQIuxY4nzfvKY2M6/gzVLWn4Hq0vz6SfA1pT+7bF2fcVPM
uDs1opX62ciBXoAOyhObE2Ts69Oq/6jzIBzut9kmMe29VRXsw6gKUCNyj1f102NW
Y3fFEZrhc8yGMSpLXunAr/K/TWd73tjvQvmzKJjKGUO5nlsWDFtOM6pCZYqkHrJ0
tP0mTxTqIImzpHf7dPKOwfmRmCV8Qyuaqr2gy2lp4vIa4AbE283MUgDCftIHeJsP
t4hMYjCsADyF3aPIdfnKailpKbQxpNimwTQtZ2E4J2dtRbLSIllUFAN8d+TuMzP0
0pjVF6ujFtB6tHeFMg18c3qc3MPvDKqLM6561pInB1/vGQZ3IpOVw9AP2IeWT8OZ
la9HZ/zPLMGKaknphh2rPhJ0Cvj/MvMIxtLRNsRx0ws9K0nY+5zXzBMfJo1kvDRq
XbDMLmpkB1bYKHe9B7vW2BWeTQ8YGtg45NtooKF+X7G9VoYIUzQ9GWKK5ypZVXan
QiZxQKzq4PB8QWRAA5rsxpR5N4qgY0Ft8va95HDfr4Ahf4wSY4Mypj5OcVC754DE
uARU19iZq0Mrmx4ATKG1dUdqj0fbUaERF46jQl1cMeDSQPKiscH0aC4PpZRLYlc8
hSs+rI0JMW8V+4binRPv0S3xgyk7ZWqBn9Qvmy5KoTLSeDKFeIhhCKqi0kre+pn4
3q8l8QLlFYRL9rAeXT1WTHWD5ytGXmvOGinOOukVxxcvgw3LRbd6VZbI5ulcb4/O
O2Crq6tbQ9bqzyVKSSaZ1C/LKVxLXgVj+xqWzSUiN0uRNKiiNPJ0lglytFH3U473
tP911Mz527dvfWrMZaS3QYiuzptIz7S649i8vgdMzNWK9dfwe3FAbq3Y9xKMp5Ha
yzBkMPgie4EZ9Cd05lZVDhPro1l9SMOqNSmURcrZFmbSKFN/zL31QigKdPczK19S
C1KQETph92IokEKAQ2YQDuD6VL21nu4oXE77VyGE3lxPfZpzArOQu5b8F8ffqQTw
jSAwsfYkyP//k9v+sshSCRqXGmitAn7BhJNl/juJ2K+ZvKpjFhhFHNJxDJx2nAb9
Af3FJe/5nO4OiRZvc61pbuOPPbB1u8TQevuKThUEQKL2I6t1Mn9l8U8l3ACgNMZ+
QiTDX6VVkE4GRJs2zNBB0C3+yngrMQ9soOOCTElkNtDgSD8SLL4egWdmx+qaVovw
JldL6Ph2y7nAIkL9IxU1Dtkk98hfx9KP6xWw2bcGQFTuo4FnQ20yADrdMLIPbUVp
yhZKoOQYkbTsdfxppgJ0OJy2B1qkA6x/0Be6COuLq4OGHZzVkdJ6QHYVTDeAs4Iw
F8rG/UyZs8hOi4wHz1Jqf97hubU6ETG4n3NID3OAITmzhNZUcGEMCE0yH7SbHdTU
6RHXfcs/CkFAC2eB53w2VBD4SXOWX2oaqx5/Gu6ElH2XDsPo8O/M0yob6oUt0SBt
Q5F5FK6fxVqdTLd9Go2NJJ/mlpdlOdpHvESG4ecXb5ksMSYO49iDJSoFEPluh+Zo
AUip2sJaBVO8MdDTXs4UgU9Fs0TIkreMks8j5H+XEO+WXFkE0HEv0BZZe4NMG+jl
/GfqruT1d0cMajiJk6/b6puP2mV24Eyyv7JNRq31bPlz398g1FsDaZb45FU722jS
iCXvrQPYMJwaE7P96Op3k9pNMontiyKcrdIttLeG702t/QqLwYoZVfby7ewAZiJZ
qZKWgP4+5xx6RnUyHOk4Xrv058uT7WZU8WJelAgPMpXY7c1BH2kRH9dqg2K0MXi5
SoxWQ/tU9s+E7WJQkL/PUl5uokimBiIjKdrcyQOUjdPABZUA58Oel0aeTA1TZ+kh
uKNGWceV/tMqe14ptHU3barZx1GZtp1OKgDH0zM7ouwm7sBmRDfa1JVSwsjBwjFH
t0TQht301eUpzDNdVQl2lrbqYHUFHuHav8jQXRK1ZgQvbB0vuAsXa5g2KraaPFFN
xmhyssqrjml7TdQbzQhy1tcP3bgi0PJ9R1SrEDM7swOzboiBBUoWmsbvmhbmy+Uk
`protect END_PROTECTED
