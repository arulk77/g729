`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
qjTGYIx4220HBtt/vUd5sFJKVVzikl0jw8I3hkpN86uFQD8K5MHeyhtjJMBL0xNz
Nh9Ju7gqZvrslXtDCyQKlD0Fd5yVEtNDO8T9ufrALiWmT1jP4DxM/E7mREymr8qo
IxOhJzm09KzF+LuazzaxhXB7WJSpymWf7UDUVJHA7voTziY43HW0taP+GDF3TaF6
54aXHPeuFZ8xCLhveTAvqhkAX3WDNijNHLLntr/C7Db7xs/ZgVdk1Y92uKHEjr+b
qkUdNcsIpR+3Jb2syrjLrZL+98bajHQguaxR8X0UidsWO0GYiepROEuDNelmQpSK
blHGsUGp4czxDl2AaQE3ED7nz6iZHaqycIm67ZTj9sEiw8f1MnaGkyHGzyjnXKGU
ERIdBEXS2YlkO4EQ3gF3W3yOtHNwjBpXAcHwqhqsCOWt7V9WYAAdMQiBSccn4/G1
OrbgNJnj+6r3Imvvic4r2s1qDF0NhwEVLuHpIK+0eJ+fGgsQIYGZ/X74Xukzorai
WioaI4lm41/a3rTDbo+1vWK8OxrOlHumhlt7CyZQ8ZdbAgsYYBplHRFwrsYk7gJA
14vDXObVDv217cAooCk+4flDRYcdLKuAglb7V2A1S0OoJRx0WvQ1gd8JD9ByCSJG
eDj/4oFItReKnvyEanIj3w9PpFmNKRNVAfcQYh/nEgqXIG9JCOMWDFyzKpvWO0rP
+58RCUYsksnHICM4s4ld29FMWVm7w/S2lCvBEsP42T0UJkYArQNNjQkmPKjvZOhg
RiIluAxzV+nmv6DK29VUUJMrVM+CBDhl01L6sa8jiF3utYDk6j7LDcIbSsh1ko8L
DpNlyMpr5IrGNCSR3ag5Xua+C0SF90DGjK4GOFAqNDcBkU525m0ZlQG062qvUCvy
8BQYhoAaJeom9+73kpFqfggMtPz4Ilo4WFXxiUNgxMkw873gV+iPPYUK2vqsLABR
S9Hc/t5pd4AytxNQ1rUSGjCcSBQ4uXK9o9LYP88kUIZRK8pEvsvkSLpnfPMgHx4s
kppjRVf6CCP+F1zjRj4mg6d0zdgeRxF1AyMhGNx7AzaHIeN3xm0PCqfPdyOYmn4r
tlGaBQ77JrO88Ed7AIqiL6uH3miQSyoKKGNFqs4Fi2aU4dtfM8OWVAusQ2mj86r3
oVPAW4W39jDlUpcCG5U1VnlOQ2x7Rs13t/n58PSoYixmcqpIh/Xwg+YF1KT0nqBj
QNAlVZMBCqXJaRYncCcNKaDQsCJ2A37EBXTj3azSzgqqa6IXZUUP5iN9MJPzhcTC
vHqj6PZLflsFioTd4KLhZxmgMGe1dwJNtuhASKWMUAVRRWyPZe/1GrwKPOHSq8MK
8m8mBfhKHpuLzXh3jZlH5Ix32TZAw/TzcOj/ndRFaxz8afFJNv3sad3eoQOuoWeL
qcb4EW0WFxvjfTlRp26NDJvEhARkVcIomG6PPGF9M9Mp/q7ukgXiDwFSRSL+q1sK
a8h0hED1WdO62jjWAC/GtXip/yRXMmg7X+ilTn4Nu5DYnUUbcfkPty8RivzSmJjW
E27chOtl51/VlEFuKxhS+KZ9yQbcmL9pQNr2mF5jQ1tdfZmSvXPkECWp8FU3FHmN
P9LLUrUo/Ku5gF6lUVH024PiDU/Yy4uBMOAwRjURCJNseuDzDkE/3z2KeT0V8be8
CTYi3cRDQfoOshbVrj5t01JEKl8NwYaU9XXGQV8nlZZQa+oyY4Bmt7zAx8IklFNS
ONCC+qAh2Q/FYhNHb3ELreMsiL5F8h+uBmzQbuXO+yint7s9iXO4lYm+FKZxDbPq
KpFBaxbrHM2GL61sKLKWjqj0y81BaATvTmGqlgbgomIZogmep3Mvu3xZ4LmTwnt7
EOy9aO9WmrXU1Ygw1yFj96v2HlhcRIWjGmzfEfk/r2r570D0XWv9SsWrVzdbjend
WJ8rjALeVeQScePckaPT32h8fkb3ubMWM773/HlZ5ZH7zYfvaqJYcvteC9YydIro
DDTjaW8iIcBi147GKK4uBn/6NXX8lLvrLvmcq62wIKSYsRhinYNZ902rs/XqNy+y
HfuLO4VnjGzO9OGTYbNUOb3PQxPD0dIswiDlUDZI7B9d0D5sAaWYdeqXfkvUPwNh
FBG8ULbWUkn0L4GvUOLeqgwR7sMlrUzpOxT/pwn8rpUHuq9ISrEndRzNluq7po3C
zDvQqKkry6o6NTnkfAN2QWT6p9+bJb6TYCfefn+gp5zkB1J2Pw5JX+94TXPGPSdI
8eNUIdY1MOgEsg3Zc92ShfwkIEiZM6/B0RUUgSzOWuMeCr9X22/hHEpZ7AIoASae
+leXv02stw4dMJfdDtI0bh5nU/8m1GJqkDF/cW1Qlxyx9tt7QUBlKgqtXEXqHO1j
3iau5Ao+WnWrmYDw02wpFXJk+vYkk5LQu7KdM1RruakV6pad0zK7bFLf1xrD+296
t6CfFfGov0GwwjOYW2zP4ML77P4Yz5ZPVFAcJt4imxIpxQR1z+62wJWdvuNybW0g
lV4Ju8q01bKi5kkiAaRs3kioGBO3+AJ5BZ+1ia5kT25uYYnnhTCQFP1YOYBkpCgN
Dgf6ZKob7WE++ZQFu/VuYOxR9V50kjTXnLgZwKzF/XhW92VPysc98Unh82tN93o+
l241HXHEvozSEidLZXRXag==
`protect END_PROTECTED
