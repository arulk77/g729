`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu476G+rgLifFK+kGNUpe48PkbQouta4w/owUrpHXcAyel
eU6GRqKEnu6HkJ21Ra6rcmCiMjm6P6Z6cDuKdZs7lKQKf+CuORQ3Zl6pU2SqPIW4
aZIjs/259nJ6knWjd0X1g+gFpjaSslRbcacI8PmvIJlAgCsoTyDvAbKqoVIwmjm5
jCl53BL2kejmO24ZzlTbVf/jRO+vKSeIl5BRHIboAWIyPJ7tk4/MVdBEbKBvqXpP
sUdzZRtVpLNpXcABDw9azt3FOD1DONpqvjugYszgiIF8jT3CKsvB0LpCRpnlnpMZ
Y3Ts0O9mEMA3m/Yds/Titv6dYl18c3VwmI3A8N6a/s3jjdZhzaS6qZ4Uvj0+W2Wx
i9IPUhoAFNwCLzgMfOPIAQ==
`protect END_PROTECTED
