`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
qKokBNu+8T9jxVu/jLhu7WxNd0Zvn2jlcsoNm9pylnqBb9hHb90IXSQp97hpjBcF
+Igwhu5WOw8tC+SCoqqtOqc5H0gbNPRQ0MFhFoKKMWxiRKda/VLYRv8eHCIhSofL
N0TfA2OeMGXpdwLni2MWHLXC0r331M+4KkMfW4d6hi7KOv0HpSboUaefJRHW/2oy
qo5EPME2bHZrrI+V9AsoGWVJngU3bxke3sI5/0nNPw32vURXnOkU5UV6pj9U4j/n
33P/uBBbmdjg1hGGRoDuE99Yb7nIXfaBkffzBZMabJLN6dbsuurzxmW1XUKidNTz
eHTr16XxK4rMdgY6DYqBGvLU9ggzQUjUQycGmUJaiU4=
`protect END_PROTECTED
