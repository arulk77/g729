`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFZv9iGb9Nwp1ONi9HkGOgD7Q51wn14qnYPmhq0+iEGD
GM4LSapXc/cYm9mxMGPQuWkLQVNDPD3LhwkUTZFGhCpjDA5KD+aYyfx1JuRFjydc
m+X1bmVnF76quh5iAH4D9qAtSFSup6mmfZ5vwhPx0Okd89qRTxQlhvuc6qPYou5H
QXrh7WG8lA4qfMSszYeJJd+zubM9SuZow5N2aQXULykkzXzSdDVc9xpsSD4M7i3u
EBj/rmhz9g7OE9ylib+BHuQ+A3UVRV0rzHGiBhW8IcmekZxnEJN2ewel7nCHWAWe
oUV7Mo2NWrOPLaJE7Q6qcYlhXXT34Cn02DBfnGh7Neuy6OpewomrekYL/OHBRsVi
S7uANmqJV5HEjNmb2SCmJyfk6aRMp7sFIB1256XZ4qM=
`protect END_PROTECTED
