`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46s/U/j56p/viqegbyXDz7qy3decCCeNWJjPA1CqkP9O
RqljS9hxA42uoiFyEd6W4DxaRggE1mV2bvf8j8SitHdRjMqeGxFIbJmwQafDltpO
PF1OTzTP+PS+xOvgZVBTAbmsTo+AqbKHlmNqMUF0MJK++wPu8tHNdq2wVpfEIUW7
Z5qUGHemaBtkZaK41KT7Nm1i9bhLEU+C5PJh7QmotgK2EierSf2QBU+xhyDrwwai
QSYW2ZVrpWN+yjbSQIKrKOycpGPff7EtqMMpnuLzjDieUkOyOvfSmvJxMazKglwj
yFiixOYqHyW2priop7AnOA==
`protect END_PROTECTED
