`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBfem+iZNo4oMyNzDTqN8tU0MYMEbdWBsTb4W9L+zZ3e
aNqjHlhwilnHmI0VYD+UA0qJZcTYlXWK5TwFpG21MVSAMRXPTGRKpins36NJoPCR
tHQNFIY3vPYl6OQqRnXh8EyMYn4nI/EArnv3sbziZvE9k/bRavNluiPW2JM8DKTj
Kpp3wnKxV2ckorM/rd6bD4aFJxi0jMedPeOkAGnxqNaKnMBoSCNYNHbDeX6oUN5e
ezKeguo6NfjTent81aXCLyfDvf78QjLnJiyt7j0Ta2MZH1VVp4MpUu8OLBPpGziT
`protect END_PROTECTED
