`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAXy3lTixT4P629dJVwJsvV6Ulhh8o6g8Yekzu+Z73Abt
oMujxJul4SiXJ/JyO4G1I+1o9EdNr/Y/oo5TFeeNOyhJlbgYa+GmUJ58NpPThEMz
ZK0If/46uE04FM9hXfANICmdvrMdNDVd+PdCD0Lu7+B9vyWD6ZZGEL5m0+SjQS0N
OAjr2KS83DNnLRz1mZoz3IgDwPvsjfS2xahw/HaFUsuM0HIOCNQthAIJDkd8Y6Q3
CZufsHIRXfl89PcNmQmt4tj/PKBusBbQ0LKlXYs33mQy5DDGrLWD4ygD3RH9x1GU
oQIwnIs9TROlMyU2GOY2gBJMIrs3kklndHv0XmvmQBilUW8s8a1BAOYlnsuCt8dM
BLRQRmkBho78HKV5HqTWC13jXBGsGr1FDws+9D0u//X12eQmIlnQYMiAhhvGsUO/
PupcCwOLMeA36vaO0ucGAUXumpBr1kGJSRB+59tofeAKSUv75VDWNXnqZstD/QYr
a/Zt443QL5Wwya/M01jVAms0H+ERir+6Yj1scwDXF8G3Qvg76wTSsnDGIUU6WGff
thgKQEDv6w5swMB7UALHM4iVSIMa3KpS9yna3R/F0aiqhFNSIOB4oV7N3yNT4nfc
F7yDVO8sh1J1A5zdofHfEi73QslVRIrLsJ/3EdIkWFBM/BCbU9KMpe6HApsChY0b
to5ZMOweNi2jNfEqx0N7LG1NK1pR7slnOqY7zYzj+n1XA5dfO8WoWxgYRqSFRRuv
pq2UMrgCFfEKv6afXWAxCUf2tdAtNhJMnw5NV1EhDXYN69ap46hkAp/Dt6ib8vJ9
4Zg5/a6pqJQU7pw8thv3Wr07a5OKTftC4S/70ao3NKAPigGfKZt5PAwhDF20gQdl
+zPB6Z5ALBgtYvqX5oWbjtTlEvY0Wv5qplveKCP7b9c0os8rx7rfJ5DVT/zuBkOy
JT2WFYH6d8fFnfk0jLD2Na1GGai5hFtLX5yc7cRykhjCOOfa1al39Mhh6YQ5x/ia
DlWcFl4QMI5aZQRW8axrdbX8X6Umsu6e63qD5tgxo4RhsGwjXA5fCX2NNhL49F0S
UCB12tGBMQa48GchMcC/4NKuW99WSAEx2KWtLqb3vfoepB9TVryS5ki7mgOauclV
dwV3lBfs6GeBBIdNTyFlvEsYPltejfK+ybjXMOGzsxyLj3xuRKuA3xOxGZjP2S3+
s7EAcCjeGsmS3BKzeUB9rtzF5kpwN46lRZEdhOxd0hMtbrZLaDie1znc5M/H4z9N
T/U15teP8CkMfsh2rGZlyKxDs0VWkAX+OZFXOx1LcAE8LqR5S6jhPZ5b+a3dkJfH
rM/DVngx0E9sh84EHkuwMNDFJ25ueMsvYJ8wJ40pDcsj/SxD3rS26pLoOtth4p8s
iJSk+Ghz2tXZqEXwb9sAAhkdhF5Jjd8IJ5CJM2y3WvlVxWDS3nyleUbe70Lrf4z2
qme4JuTm/MmiuaYhEpSxHGVFC6FjNHdNj/WV9K5bFGUmvOlFzLfbiv+IOUWNBkt3
A6+0PE3vztCxRVUgjh4b787wqIkBVqp30fc9yjs0KFZncJAGVWLUhSiT2PFdkgX/
b8UFl0mnQ7GLbsVXAJLxzq3Upc2EOYdztHYZkO/KHv6iP3sCL40kENfUrCQ70gii
a2vQvpM1sw+foKw7jNfIgHJ+GjMeAAHHguPu5GkRj91zMz3TZxNhZSUpy2SLVBGt
Ufxq7qiUR1D/izoN72FBXc+G+e399KgobLfa4U10hQrWYlqFRf39N068Tk8UJ+EG
rpVdcuyFkOjdZ72yoRUjWdonajZ+dmv2coyaP7mQTrtw36nCv7V9VwE/pQksAUFX
2wIQCbHKPkP/QhSEDu54hhL3kOk98MtWeCEbSNKaFM5pcf3DdJd7xwBI/oeznYgk
OrJ82QWU79goYe9g0Awa4U/QV/ylRpxUfht9WaUGtnD4+wVBApjyJLu4GkdApIao
Y1Zk5KtG4f7puux9bSFwNHG1s2D1jLsieGyR0qBqPrRKvkMwaFofEVjbLn+a6oro
X87M7cOk8snhb/bvUfVyiOeUbLMrVBkmGJBUC+YWbvAWxeSYqz7AlhbtSCXj6I5p
JQ62Uxl9DtWXTsI3HitjCkbupLrx50dhvrRCzYT/vnGnZkwJtIB61ZW2vAjVlESm
LK8fzLhOeAv48D3o9trXRuATZn0/UuuMkSoUneVNqyh2f113knFAAtF+41xrjOO/
PbxD51uuQ3S4IBu1/iQKhbk36khmsJRfnDMN1bMY+PsXk1bttbRjtdDuT8H88e4/
geVr/DDPfoDSb551YrLYoXF7JV/ugVnG+vu6WHCeLAiEFInwpwyVNLbVflc5KE3i
CKLPfRL2ufMNzoBO+yx7bS/Lg0xU96kzvfrDE/BtVMGbDcAJDk3uB1W9xaSQSfxd
MVZ58NIMRIxUJcuHS87/shiYQ4o22UOQPQvZdm+SrB7Fd/LDQMg9Dx/xAw9D7S+9
/DQmLFGTrpkefybdGjCZIht26GZ91zQ4JP78oQbSX7bbIV0ir/6+IRlpIfoGSi1D
habWNH3HrnY0KH62oSm+q5K5NAtK1Cm9eAF0G3sRg9Vy7OvhHSN39/ZT7Dmfk78e
GajfIfHUnlSbsdrxguPUCp76eN6yt7Yhx3ChrNC6HyiT3hRVULfxVPCRjlmp/GLC
7UuR4OlQbXMxXXN9BuW8PdvxayeazT/sV2L8wzXWj2a4ECpU6zvj8GRLi3P7jJFP
11QOArtC7EmCKvlHHXusZc8e/ETG5r5oTFxRQfaBmTyziYzqqCu5zxkhTbB8PLvN
kVV2qjGIo+Lwvsy4tYyTSX4Zx2uJ1mNf7HlA1AG7HhurLwue/vZr+pbr1H2QzFrZ
Gckk/tMTPVmPFZnfSJs0yJykt6KscpC4E614ZIFhDZxYitFaebCFZ8cBVVNHvRaB
M+T/VGku1gjQLU9wxLJfwRhEjVFAQVJTeX0S0R2749fltBdwCxW2lFNPEvyrbMdF
LDSHMEh4KbPmD18OwIluG0UnQ7X47FmGXhDeZJiu1ib7XglFb5yXOMBvKq6gGeCQ
nc8ZQC+ej8NT+jhAogpJ2I/5L96Lq0FMr2Va2Ibtk4qyDwqbB1nvvBKErQCo7oHj
oSiN6O+ukTPDMQQX3rfRVb0+XtPaXWtNIem2vDfiUgwwSjkNWc2E8Cqhg4S8VNTq
p8LFQFf9vaXFUNrHDShmS9XAMbMvblQT615RyiIpldGtG+BuCKug83nBmNIv8UQu
PHuRauxyyHwDFJLtMOceew==
`protect END_PROTECTED
