`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
E/5d8KzEiLiA4FadBGa6hKP2F9KcmnJdFNo5c67TER/YbgeAGYLbiVP80mVmzDKn
Ss7Iy3q3yQyW/kowJGd8W6GCrWQOmgimls2I3H3+IQZf6Y2tBSSeVWu8nCcdarH4
M+wfu9hsVu0mosE8Er5mN3XWzvh5Yc6Op5t2rqbALS9LmqHGj5x8mcxcfXBXo3l9
3AqVg7jeFFlxSOqmZNuU8xp3iWaVOeFwDryldq5s5EhCTpZQXMJFyYFgMecCyqf+
spXM9LBUo53cTxLQRKzzlX3uQmUhPGpMIaUDv3cYnyQ=
`protect END_PROTECTED
