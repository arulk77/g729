`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41qYOUiGdy4xmPgeZbUOSUO6oEnEo1jD5MpsR/mPxsTt
vDmJ4MOuoshD7b7BaOnEVv3+RXq8JdtTv1HoiBPwXG/CXD4gX4+VAiPlSXZCQYd3
XDAAl6YhSCkSftFZ57hXb6Tj3+XsBjLepSAW3/ENWlEGLgzSz0RxEza/fJan3A1h
MDucod3RkoBty6wlldiqsdVyRedRcMunRIUzwsY8kt89fMOaU4WboO+o2qoQ2sLh
5CrbNgl6CzTY+D2cUR6gXxNzppN+Jz/9bKzIRBMz/CtaBUIn65k+qXAD4DdtW+cn
uGTaory/WBXPqJoY8bUwiDpw6Tm5LFEqnXKvnu7WE2YN8v1l6Ly2F6ZSpcsuYihv
byMByJ6hgJgOwSCwkxAbwNDOuIJDwxOAuR7hBEQOqVDdfV6Qwf/kc/qOA1NrDw2A
w/JQ0aZxKtzxJRvaQZHg6A==
`protect END_PROTECTED
