`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveELATlp+JUhPe8bAyyDzG2kpJsa7LdRt6RXjTdrB+0/i
9n4Y5Wbl4xsL1UvbE/IxcOlm3SCVCpj1DJlF8cy63tUIMN5OavWL3ozAOLOlrG5A
LowiSz5SV+o9ltFiQE+SrP7RP96VhT61q7wdSiZrI32SZN4/qFDOsynMem0a0Adr
xsaFChjgyVmoK0cW8kbdLgtMdwvGpzDVCML+r4bdnjohvSk5ldeXUzJyjuOYAa3J
`protect END_PROTECTED
