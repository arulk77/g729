`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aXvg4zU62GkyIUbWr8UMnQdGlX2wU1+gQafOtXJYhazW
9hgrrFK0K9udiSAex27F65f0xXps5BT2Ge5SXofVSKkSH2zGKgYDOEWDSZ8dW7n9
986hWQ8CT5pMfSAL5CeunQ0jGo22DNXWcCiKG5NvI/qhoJkJTKcV+RiVY/tSeQh2
3UBVuUupzredXbNC+EP2PChD+K0Tl69MKpoogz/20BpB1ygoRxuZWAGDB2mIjdZn
yR2VtrvgLsVho20SiWNv//f+S484oXtEWB5qdufdxRlwyxjgWFo3gQtLpL0d1XNN
C/gyH+toFM7ndw+qFN3FHkmpLiUoUv+blM0JTwF3bqihT87cgYFU3eFWK1KJTfrm
EDJ1+DLYdApzD0+yJ63V77lSJSGeeZadFeVVE2eF/DEOsf39i/L/6EkZPtBqK9mN
29mbKvLIgSZ5nRACPUEqmBEVGcL6pU9Xs3TMEs0d44mJ+4WdiqtK2WCivuHM0Iw3
`protect END_PROTECTED
