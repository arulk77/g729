`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFyKTGOaPSbipWCx2mnnL+U41PZ9Z1GjPlJB97JKJDjR
2w2jSyMmuf6B014KTkn8j+1jCnOlvUPuZHQCHFs8G4TT9t7s86M1AqDwLzjqrPTz
jNREzqU+nuxSULbNX+9z3HErawl8oBNy6SlKLpboeYB3FKsU2uDpGipqt3qpcCn3
7qb0m5D9F3ywWyMu9GIftBPllN/sQKS/4ponmUk2AKkqeVfsmI+31whiulRuZ/kR
mu90Uwbb7TCxSG32VgjFyY6VlREknzCam05GoxSppu0wdzSPsKb4k0jhjAo8PinU
11CK0XXa9AP9uhKHr8SXnHA8k37d1nMh3LNMIJD4BJBYTUeWfv+EENaeLFYh0PJJ
QgFKNpoDD49PgvtMcIylp7xXx2VsEl/s1c6l2T8L8JnrZu1pK80H6Puk6A96rRJ6
uRZuNYsUWq2++4NfDRiPx8vhMlUzurUvKqD88fZe6T7/h8sYHuTJ61/4wZDBTkT0
hbCg0tzvqRcGTCyRs5z0va/c42tnrJ/rJH/FzvjhnShQGrmMEJQs67Q7wJRliWhd
`protect END_PROTECTED
