`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBBPZSpbxUxOhwwgqXG/WR8Dj3k0nzcglAAl3lVxTL+e
ZuayR3zWXChCh5dG3qhrXdTB33T3yvD5cUADz/impEMiUUkEPtZsDmQOimZgus1r
/gvqZBhhX+hmvZ6Ld1BryMJEh/kiRf40h3rat5cE0ayq963Vy2hcmJezL+1rIWUZ
cc1HYJSgWEpyKmTQxAO9J4ODsBmEYwyJNOr9rAyCgGl29+AZJE5bcj9V9hhBuKbk
`protect END_PROTECTED
