`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAbL4J/3MhrNDtz0LtSdoHJYEVVyV0baI05O8XXti0scV
S+7GZybwsLCQs81mQlx3PyQ8y6bMshKbPuquEysypm+VjswmGQ2KcXh+aWIfMCB1
ZJIf7lp6YUVrJxKRMkgw4WL2W1ghZwI/GKg2z/y+DVSAMA5Q8sLwQb036UXm4ion
LbGlx8rfBizhDixYjAYa5l2gcQoSgZIil4aljWSHXuAioQFk+IUczJhmZmR5gTMt
DFIz5v8ehf3hZ3TJ71goWTRzeLa7HEUvgCGQm8Uf1CFFJpUJ1pXJIjva5OpAIb6O
9HP0CBsovQYb/VCfIn9oHIYhRPKAX5ONzM9XYLRcVzFb+biV7KeKobE8dihJAfHu
p1WN8aIP3fHDXTjTpUlq/Wl1PppLL+h3JShD5ci1MnKczdJyCLNk18UnmlsMjEVx
t9OjomKXjlyG574R+lqOYRFdrhcy0UunFNr53Sc/9YtDoMDU6HaY/Qf4ugMENwqo
VUerRma7uc4mO9gw9PhHaMUZe82YG4JHiPDyQpCsUb5mwSiKj1Mv2GM91BMyHOt0
ffCn0Z75fCeExNRAUlf0drsuAJ1CTBOvF5hsnWXFSHZtK+Zrd6ULZYEW1NQzSFSt
smFXaNeNkAWekSBAqlDPK/Oy5TqKzevSh4vpf/UZ4/gUDH2/I7hE23MjQD3iQLAd
YMd0UIUm4Z8NEWIYZewNPQnevRqqiywJ9vBKIq40sPB92NgMm4RCKljX6B3hjyuA
gmWM7/BTyoQTIqob5OJVWTmHYqQQ1isBFRu4dZOcGB7SE9CYJ9L+8brmcJ6Zjhco
rx2bmJy2avoQrn6cR0gIaUAO2Xwk+gMMJYjCGro6AoFdZDAwl+Bulqtp0GqwWdQj
1uoFIzqcSuFNiZ2Ojc3Zw9Z9EpgRp6MC9Ly4fbgGQ55xno8Cs6h2NGNglRiuNViy
1QY5UyH89+XPk/vhX3QxCaICmAScu0frcU0xC2GU/LoXkGZwAMGfaZN69qjmqawh
mupsg9RTUPWtU2Yp4UgmS5L0LcCav+iZWnGhBv152PUpQaqTa8Z3tw3UIk9Ri2k8
8XOgu8u/b2Gq4GBB/Ut950Aux8zZCh/ltmVqXJllsxZXl89kDRYTwvTSh7n2F2iu
CtgToSRj9WIfVbCIqv3kBj+hec2L5fIi1FsIEIPUaBHNm44JT1E3q53NbYaXQKQD
jUcKxtm4j8ofUp6y9qYupRoFMnuxRhqk+zfkN0qzN5vcBfjDMft7CXsv/s5rPtZF
FRusHhU4w1sCREYmYjwLOCFBZZH0YQIk8hWS8t/qoCxMLy7eTqpnTaQAdp/8EmMG
F9S6zPpad2FT/KgMY7F65w6cngGRlF8SDWUYtZ1sIIJ1PO3B4ae6fDrXz4Ohvpxu
fy5a3OT+sT6kunUcT7PvyDfx3BSIgxsSktXxBnGPjEwOCPbUCPlVh26LESgR66ib
DP+h3stRn6dtGl6XAUsE6KVH5ge5o2RP5USaAlFRKu+X7xOVsg+dJeaHrUx6GqKK
4yemcurxo39PN4qSp6u00pwhQqjIWYjAB/+6l1RWCJ8pCvlaFuXUqE9uUiCDmQO7
5BhudfaXp0HVGVEq5v/Ol0YsFDCzT4eVB+IruG2QDVBcM718wCP0UGjPVO1ouNEl
jxiX0F/jgG9nBzLWPo0LO378JRN4FZb2zuFTY6WuNf+a3uiNc9GHTC6UgIegR1ou
L2yRPy14PVkBagi8jyEhmb07PQW/9cRbxKj0oA0CknyM+N409C7mpzskMMKdrc8c
PXKLLVokB98aWnjS7YTJ1ZTuMgfDSqTuE+NVBquZ+Mdvt+1DB9vfCNzexIbDsKoo
bPEcslI3g8vwHYwtB1rqyktGdy3p+tGitHH0vvy6UnxNjexlkJ/TjuRL9agu4Yh5
WPoK2OrP7Yq7yXUibzM6HQBzZSUsqFq4LkN6wwUc3QyXG71dk2NhjOuT/zLwkRhD
zXV/tr8fmJea4D+tuW9RDP7BQL8/d9AAfjJEO/an+KI9Jsgor4W/bs+NAzcosEMT
6YmHWX7Y4MMxiW4Rgndjgw0kgZuMfzZdwklxSXQdJGqSJkuydss04qWwXkeNmBTN
rD6EbQWZmXyGy7AkjPxekJyvNDOnuY1eaQqYV7WfYFmNS0iwQGQnMdLVJpVWsC6x
WyV+5Gqf4821k/JU/8euIpGYb944KuL73rIH+GxfNueZZMAOb5PdNiUuRMcmLfki
Eg4Cn+VqWFuy6IG0KP3+NakbKOwT0vxQ2frnh60RdkH5SKwLzasXFp74rBpfC7KO
nF/a6VxkjObhCoAe3ph4d8j+LbkeeXFN5XAn0JHsT7Kc/7ue/XjoQZs+/Hb2zhzJ
NChPog0u/vxv43YMjj/icpKFJAEK7xpTRaiavcRnyO/4u1+asxzWI4kpDfvbb1Kd
x19fRSqBm6THHa8EQSNPtR2xZAMDFoUly4aXNrXod/dSj7sxX1NNuJxGJh3bEFMh
Ad9aA/pZnYYvHkaMMRTs19AIduGr+erOcANiAuG18R91sCIGXN48FQU57YW4przV
fgqPWh6wV3Bl19/aIUBgsfVlWy1iYg14YjRi6JUDdbtzA8zoKCtwGU1llHw5rmQY
YXV2wUJLr3JOyoVMVnsx2Y3Au/w/vjVCAaDSbe8kGEIKw5GBBBV83HgVTm+JDASs
80jJMjC29DXA/mLuVVFPseCFxE6aqzZd/lh/r1L2qoEWjVKfDVhnCHa7punNTqwn
1jG64oEPpLN2yXU3jULNe8Du9J0sFSt0p5PLUBnD0HbC4RYp/faktVOzNpirgJpl
gqGGMYoajAFEBkUTBxEiDOWC6lJIEHTQ8/V3KPIUDROTup62hqus6QJDO9S9LmfG
R6h/ReZAIIFeaolGc/LxPR6m/Na4o2eoHh1FuIDOgRO0iZQ56hi71UpqEx8lkHBD
CJDuJiFGOnsRoAuOzDZgvylBPfVpHEOpe2v8cqT8YOfwn+/lOXN20d99MTt+81gh
ya/cXzy65LlIauWlh6uErqwIt6/eL1GJWalVCfXXg+OKheC+tZviM0kwEnk+8GjL
u65WIeqRUHHyxPXrN5Z4Fnm4srRuRhBKlpKz5R7IbW1k6y1+JZHGebGg3r2zCjkP
r7SnTyGs7144POq6OqXFD0+GK9UFHPL3PqG0SqaK3T2XMtp0FyfvoLxtANwkIvq2
jUhQLquN/2cyzobYnP4/tPSL8XRoA6zBCW52osx+orEpcDjDFjxh/J+BuUAO0C2e
XrwdaZ6+gfZCmJkLvVhW7Zzthlv+ILxwDqZzTImBetF/wQKbsof1XTV4OSSccnvU
jHCsUxKisrlRO58kgyM0uiPK18OTnWvJEqoDAMLOsAChBxPZ4QDrHPxRLK3VgWxT
fSQWrJ+ijsMQGgECK1/j9+q8L2AYaZW6lGTTiRNCsgi5zab43KgcRaCMxcp490RV
3rAX+w1PSXlVwHBVHkFVHbQ+zyVXNObZ3xyVYTZzSqr6rvcdTOUpFitKtx2p4968
niKLlHIXgJKaI+Iyd7E2hguuQ5FX8Ija+h0HUvf+P1rkhjqe4zDjyiSvROqAVk0l
m9g2JDqU+TYSAT948ZKYzE+wu2XFm0SkOsXm0eMB7Lq3o++pU0MWGrEg0vMVbn/Y
KdaJ5aDsuVp2kRNYeAjPztHY3Ixj35/KihaVWFnWA+mlbCaBNnx31no28XtirfTk
WCiCCi1rdUPs3QzZuHebx5cwwNEcZh8GgB6BNiN/SUIdTlp1cOvkYo3DCormNnhG
JBaGxo//YDbInxKTCx6Fu1ZSgF3+V0riwc8rYa0GAJbIvyaRzx5h+azZNkgCzsx1
b5LDqd0A5Y5uRPhuTbUcX5Y36FNqZ9it9PSwOTtAFbPgwYdBDJt7jFsC5ntQk5hi
fr8lnagJfXb5R19GlMJIObQMUxEt9jMgHsFUA1gx6sCe09R89/Qr5ek3fhyxpDLK
b1uRIhcmIYXGhlL5eR4WXRtngW6wKQLu//zDWFjRMIrkQ4u2KQ4lJxFluLI14uGx
tqTLdgT+dOSe3mWKLOWSHbncyamXG2cHx58ZE+diXfNRDMmwliBNcJ+n0suv8Xsc
ATjeo/MO6ECO7HNZ+9KNp4F14YDkP9c1e5hl7sYStuYk+gtdhp3fDp2cQlSAUM+4
7G1gkZh8WvL7+yL2bUECi2HHgsvlQ0Xx6PD5dEvZ11eBzyd1IFPbKk7PyzOca8b4
nDAKLpdyRfnGDHx0f+mfg0tFMi5wJVGNBZ6sJNJnlw4/SNKn51QcnZmXkiG0RAvp
JiQSTZKvyeycF2edhmqfvQ30ONfQMzCgYjuXy2A6s6NT6MOkjop8hhCpaqGVoa/w
dKUVQFVbY3cJmrTA72JoJe3tBt7Fl27SoknQWOKxWVRt0LYlmFe7M+DPyEWFq2Ok
266xkZu5eqdpRNArcAfnTXH3REuISjGjsgsZSFESFxNmiEvDE/KnnaTXBN9905qW
jRsY3RcWDqayGRSEAKz/epf7BhaassLgN+4Lj4jzkqZvoy20QrEY1aCjTOgni3R2
eb5unbSBPVgqT0qNpkm3Qq1m9jm0qDnb1wCVg4X2+1KAZzGW4NDLR2xoOq9QH0mo
rTP7pV6jVo7I3xic5VGjxCUeWZGeioJTzeNFWLjbFUO2+BngpohHnxjrxm5cScWj
IFTNwL/D69FhquIpMlwZOAzxetsn43zYVNupBxRQOTtWn16bU6Ik8dzUywhsiO1M
vhbCs9O2UEU7tdjKlCVvbYSR2tUUWo9IPge+j0puN6O22vy2tnxP13ZyZnkwnXQu
/3pFh81OEoiiJd7/XywUhglh3XXAznB/6LGja8zHvNIB4bv7TZDr/psJxSBOgZSy
PRn4rVe/20OlCLa2iJ5hjKm5ocmle9HlhUlaSXkU+yIYkU78FX+1w3M6YEbwu3E7
6pB7CH0vcvVkjDpu/7nhBkm2CNlBgamAcUOxRNtN5NzbU4G7UZt4KS1i353w/p+8
qq2XYeE6jLE7NziWUzuyimFf8Kua6wH+D2K0OxVeKSVHfeBlqgS3aBk+s63M71vl
We/rmZex8w6oT7KTvB4jMlQgkHVis+veu+cMHPiyZWB4LwifmLrcZtGFzizBcMuV
Z6BqeQD4B19ao4sai6cAuMg0addytCzjZLCRFtjMAvulVoC+fnNt8jBm5aYO+ivN
isgM0lxLmDuJxSLkctYZTXbRgRrjHkwhYPz9LvKNPArvIJ6914YJPEk3RK7/mZ9k
3riaIctFUFoH8KEhnNCJ1e7hGH/qHQ00Tr0EALGhu5Dy+0Rv1VockQHPEndzxwBr
lLn4Aic6s3KL0k60YjgR2axiJ2QnVpc3icmFvlX5p0Tl+lvVsT69xOj3HZ4MSeeU
NsAX2Ll6wysPPYt/+iDnatFpugQl+KbfPFG5SVJsTDQ0WeFY3L70lVjXc0ndepKb
fSrSg26dJCHjbQ50ZrabLI+ie9RawwjovC1Wek8gtJwDbD3+DfVN2jvQjtw8cvRH
dTwsG3S2V3oC6oVqBal7ZQXLKhYcdJrwBt9TPOq0+kHrERZfcy+WCM80W/SF/0s7
U1BWo+eGWeRQ8k7YquAwhsfGRWdP01DGflbSX6nhRuBuaIQjGEyCLIZh9DAtLYtn
Pv16RYY9+Wdh4AXWtw+JD86MO9j0/3tEA4MbO1GMWelPEk+zCKXE9ndrJOCHd0zI
qqtBbuoY8X2lvUu3WKeoGo3rdbVozxKsQw0ExlXLnmK1C0mNsoqgGvwosikAwEfu
LfzfOZIsiHLMZkQ3SIAAXCk8wedK7XIsLyo7dlvygM5ngV2SIyFpTGWHdSMEdnia
XXOpVlrooG6ITOiNrzxvVq7xz5c+eUnxUScU/Ah1vXBULEAaNhl0T5mZ+jTQyalV
gOwF+Pm+y13qRIhQmFDbl2drBss9YQLzyNOUMgYMxsHWHqyQa20LW9R6PtdobOog
8ig3BOr90wo+0skTmDKZqhiggHKq3RggUnTL9VJW/20hg7BSlHgauSzlDktZ1zlw
O7dkhIP/BFQ9BTMSYQc1dyq31FZ4AwCG6npwkXNeZ2P2iBAw/wRiGLVjuIA4jSkC
UsLBWCSx26pK1MRnqZaABVciWXNl0pCly8Kk5MsBncQVEB13Ct+h7CIiKikrJh5Z
EIMvOWL6OfEoFnO4I+PWwCT4zB7D7XlDiFSNjFGDGAtIc4JPJfo7blqzswU22Jnn
Xhnmsa52qPDZKhHObxbo56mvA2jMCN/kKA6eI0YdlErahLJZinafzzCwDaKS0aVF
KkphOBda5kJDC0F/rKDupzGwwtU7YcOSYJXqq9I15yILGykN4wvcwaW1rdc42kwI
7Zsrp5arMKz96SjuFkZZmXpPpRK2KWKB9Y3TaDd4D8N8Zaa6gDYth9evYtK4HSU1
cblZJzxJ+pkVgL2wX672aF/eV2YgH+K7oc9ZEha14eWUkQ7P0sUg7OY+Ixm158vt
9DTmFk1ar3GXzNhePhWGYaqxZ+IKpNItgt+nuTo03McdUEA50CECzwEMktyN0AEq
lH4O09s8JOADWWjXUDeQ6WXaW+T92H9BJ3YU7ghIn7nQXMMTRQUjn/Ty/miEueri
Mdai+/zmUslzViNrSELeX5L6XvRZcMt5/zZrRP/FHePJnkRrvV6iWhXiHNI+8Usy
E3LMpOCJzxFIfrw8mRvl8xqifwHcsQylURzyUTqkno201tSdz7BXBXC86WmaOWpj
1PjG/uKGPNdzJWLayVzcWIo/Ka1Pj2X59XQND5NNcBVpD6K/rBnlbIIL+E3y71qP
TmobOtU9pdnpGtTKEAh2XrystDEx4xGbeUkCpAZKk6848P4oL/Pkg2rn5Irfg6oF
9nZbiAaLZ0zt42bC3zP9oipZKxaYWugsoTL6Vz4FXJRiGyTm+vCqcBnwxyV6KG/Q
BbvHxfUq5JTRHzi5znPV1tGYEAVXhUTPu8xNHENBqiuJZcJIGHt0s7XV+oUdZhNQ
2T5E8fgE5+OlzxxEpfVtT0n6mqmMwc8ZkiUt5NHUV90ebWQHNkhnYllXl3p7Ms2e
ONFdeVG6mCvp6a8RMJ0dyxGNmg/USdj7YQTs3McXkOd93jnmALex+GrGQ80YYWOD
+W4BLVAkOtaAp+tAOYJOHKVzh/n0EBg/oDss+QHRix+awIEVmDDQ5/NyEIYTGF+4
VPvTWx1qh7ieErxKzcwVyTHXLMuHKpkZiiZwlv/9RCcNWFziFevWV4mPNFSUDuNa
a9ZRnoMo/fI5yck4tsi3gv1OEBmQ9YnVy5GqEftjQR9efefOX1yK+DsyriEANSmZ
Y3z8imIEXFiys0BgVmVxbUZjLN4e31CD3lEtkD3V9FRBc/8eg2NxboXJa6RMosRU
nYQ/6tfNg6T3qLd1AvwYvzvbB+TWRSsJJ30s2MI99Y/4OSa2aglJ2bEXDm2w2ms6
YULkYPkkG2KDzzmr5ULaCdcvyCkkIRgjE0Cui/j3/TacHY6ZnCmIlEruhxQxDYCJ
o/YLT+15iP362N1JTKqLmySbIdjy4xaZXPVDynezOxr+sHa8aZpYlIVhL3vJZscR
sQIT1lTAMTxmMzVXQH0a4PxMlyG9RDwV1E8TSJq4Fj4SE9hwLVmfwp9kC3RPMy+h
B+GWz/wo9fQbY1xyMDjMAPL5HMc2dWa9kSq/vZEvX5sEqSg0F0Keq/iRC9ZrCdit
blnC+OxebR8h8LBy9G/glyjhgZALZumDTAK4OMd0btDOegJLQqL0peiMt4wziX+m
Q1tHX8i0I6ywI3Q6MgV9DcQnB51TmHACOnuVJhEtg9G7tl9vWiJYFhON172Dky2C
/ti2suZwbuWyjBboCJRWU2MtzcoYDlu4VT0j345SG20BKKi+vEBiMSzVj+RRbdxc
zp2zEy6OmsYkE4yxP8TUY/Uqn4tgAY1qzy7aXampe9O8B1JEb9QkQqCN6h36sp0B
wR8ApUsxQkC9l+6+0hTagvKNWe78eCvPCCn9BO64sVZtTNXqEtDJ8J7+UT4D+A2f
po/DCbMbAZo+03byzApifyTdYAM4VE7yzN6LAr59SD6du2QGs4hnWclGTCwGXb5D
tfvd0jVqfBXnIw8P7D1z8mRMIvdCeUgeg/cfxJtDyxaK0uJS8LlrxmyS9BM/9fDI
f/s4ZRp0igruaAfgbk/Cplblyh1qRhAJwHgLMjbmk+s+JctElGWI6x6GzB+yatiC
lOkNguGoqprRDpKIGqnylyeS6wDCzTqcb3xfzTb0AzXKqZFcZxugErb+bG7aO3Ko
wFDNbKGQFUmrUYLeU4qlAh/4a7mOBqxJTbpLeXsO2vzugJpXywb05nJ9GGhl7o44
Bnudja9P58NgEQKGUXY3Ug0K6ktszi6tWcxzT9UiG7qnmYyi1Hxy3DmCaTB9ycMw
oBSZILW0K5ZfRGNkHxq6HSQ7F7DEt8jz7xDpvul0a5Ske6aTXNVwUuPsHmEj7R5K
DNWEM2jLzIBSIWkegsl/QJOWnyPjXB/fzXT7ed+LaR760Lv8BFJwN7dBUtuXYriV
2lzdNbL+sQ2w0HzvV2mdrms7NU7pkEmYB85CmW2QEjRKdKfs/LQVuEkp8HmC1+6l
JGg9mCFmmQxTy3FP4HIicJrUMi5fm0rjo/FY4fK20YHLxExj1PRWwqwd7j3rHdbb
8523pmqJ3P/fiKFUiuUCvce4ZNVpWFaavonCOY19CEDGWJfhay7YJ/cpRzr4oBR2
Fu7Q3uuQ4oP7Yrco5bsXpjDU1hYzJbTmZZOolBbFgxjkiFRo6xWSfFZcMfU6jUVJ
Zb+9vUvmizDDDolsLGT8hbahTee0FXv0/CQAU237aEQ=
`protect END_PROTECTED
