`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C0j3v8+AtcF5TJQ1dTy2XCQbdDzHLfuyxZSj6JuEwwHe
382hsXHS7Iq28kikGS0eg/whxe9aFf12EtSOigJeDwrAmlX05htEj6mm206vtHmK
So59ao/RM8s1qQYGINkxlhKJRigRkx9LsWlwTmV33brx4un40Kfww/mgIJp4V3vT
PoC3yievgKbaGqrhInJ2oTdRJmg6FwCAttMqBrsIShxN8PgBaIqNtmicEbaX1BUk
eMGnyfW15UmNrkwI55gS2FqUKN+LOSGCBHksHM/+BEUN//qsKY+Fg7+NsklSetF2
Tx6HgdNle8UYi2/KG1Mh5IQa9wLgQdJm0LHy5eVon4T1GhUKiD/roUTTeJvU/dMt
+BzNl9pNO/pCJhTR0+sOa4UfPnhvf8AX41OYcRwImWxBNllc3iDT32+2EMdj+/e1
HKeMhqsoggdOgktJPT6Fyx3Vz1f8qBqWP2HjYe4wf511Q+j57XRe0PIJ1q+ajdhe
27nxD/ppe7WdNR25Ikra8lQsbGCKE8USRVuvtCPNAtTjEPqvaoyxpwvrMyKdDLbt
+Vf89UfDBVkk62AdtRih0XqqpLp3/+7TFvKXfj8mFEAoXPYfOhf7gei9TMx3ry1o
eA8mZAPSCIUDT/1yCohCkYGUjnx19DEYpk5vf0y1t230v1OwzdRPsMDBsp1K9sbk
OBlhFDrijb3am1NurwzmGi/kJdPKtQSFKyeSRew8AJBNyT6yJABLns7cf7zQUKwb
Cb+kLgzcvmgqjASw2zW30hQgrHalR/kJGIhXL8/pq+S/OTC4LwEyo65T3XvHV12O
2OJAlAzPVsmdgi3wQm675SPxMt42w/otLQvGUnZsPwT0KVkE4/YOKZlhCE9PXe/y
jGpSJMUy5N0iN0xVjFViifc1rWidxtMoSlvkn3blBiEjRPJE++uPJjHE9gEFTe/+
sCTiTx9T3IK/H+nfXZSMi4wZK5C6NyIF8PmhHFcXaiOKMnJaPpK2lzTdJwUY3GMl
0dYYYw+rGT1jrOoG1GxNVPoWnioVcRzHJxv+epwC/WeJTXZaX8xtCantw7FGccZI
fAmKH5KVp/8yMZipP4N7rfevk2CjOj2CHMGl6s1/JITfKwGJ9rR4EXJ6KNkUYDvx
oL+r5GYIk7krRBHRuR5Geji2Wv47MDJMTLeExkVBjUS6rYOs7T6PVzR4P3ebmqc6
KIQAnDSYtTFRteInyj0bTJgdJxU692Qah1MQ3c1SEieA5AJmRi7ehPX9U0blPFJQ
5CIJa5jMsBhpYcdgHmnd7r6NNK6vAThnTPqA/uSjKXWauCY8TRBRXJK/p00x7W4Y
5aQKtO++oEYWfZa9D2gWY9uJhumx6stzzieQAt52jFF3UPYDK0c8PEIhUMDgAbZT
31L9GB9var3EwH45ovBadHh7HQhU34Jrq1Ynoee+MdxeXQRi641Upsi0QcL4sTNO
J0orsx8AXOFQAs07hpw5hmnAVBse3MKo7t/WgfZScsIUnwsu4lf6FTWzH7KD2If0
RZ/RRUvJyuREkUlN2KLJesyu5rYTQDXLxQl6dFu0HvBX+6fNLLxuI9oEam+6vXns
YC6Bo9lOJ2zb2t7tLPPQ9dJatZiSDnHXmqpC/4paQvJuXGOMtLjY4GsynhoGc8pn
gdNZe4z5PYP1oeChd4JfXQGjxvRNDg616DdovrTuxFTiemZS8SD4W4nqT8lXVW0b
Pvs6flRW4s9g8uIGvlf55lvxPzN7QQ4nparnkCwh0fg9IvkoE65gleXojaLTygLi
kGN3ocFm5dHauBscCgqGVbFDkVd6hjaRMIEkcyI6LnMU8tc+P2i31CSmDfu7AgV7
v9eruui1U0j6aFEat9L1nzSVVDG4atMUQwwd08uU7p+CT8YwHCaibBNHfwtO+Mz4
vdFQXOGMl1ezHhWVCO01nLDii+vD/md9tGj/aouQGU6XCBHbHfo6mLCMQwx3v+/I
yhdJrbEC3ZwLy8cXD6M0bVGtMbWjHrYQoXRJRz05GRiCu7gkpINBxQNhCGWJjDyV
h2yDkWYGZ/lNnCDzf/CljvBd0Z7kHtOAuebpPbYprSXZXFaWjIhzVudCxeioIFG+
35I9XYoNvLSp+xjJsp4TmtzkdswNYfcx8YIRFDchG6+z2/TTE9ZBfX3NrrSA6wuP
HSiTNwp2yxbYEHr/ukcSHt0T4ukJjdmGZRYmtOhycjB/DWMy8nVf5bcMArIyOgIE
i+eCmfDkvevsZlgv5xvdPKyoFJiu0hX5RxdrzTb71l5sJusF3weviQxhbkiWft7j
SMR4pnhDZLGasOgLmEpfyxg8aBmp7z7olnuTcdTmMnaf+tHU+5SKgHyZ6J0mg3F6
XrsWfkr1l//Fy+w4K+pnOMdWjVIHEITkhah5NK/oQggtlBjS86V/+n3Fm5F8DfQu
NtW2N82QeQc6HRjrXKgOangkuiFxgU3xBluo+RSLV2CJ3/uLu4UAYGgHgJ2Nog4B
FqyZ/zUoRDRyV9YlLVfCZpgEyBuGFtsh20dMhbqw7r7pbdJjkyPMxf5qU2GqAQx6
Qe6ewQFE07sNWpJUG6y4+r45YP7L7BgggW4flkDuilEqPDu+cqMmZ0XsJppsdVsU
TrrRzJBFSiMRlJwvodfFOamrE0GibjSMjjWbAkIefeNhmkG9ZpLPljjA7dIADxtB
Hrw7jCUyLmSQGnh14bVnfpiiReJ2x02t9Rlv51vfS/Sy2OT7f+VLfcywn1fjfHCb
/XW0awmCdMQBuNGhyqVa3DOD7NKsb9Czczd1grR3+pd0+hfb4IXRrC3b3pbIrsg+
xf77Vnqnyn2qWLkVA8t/Rjqp10qcEpOy9WVOCSjyyeJ4SxVRWBoz4mBZPZ2C21hs
pil7MSIq8EViqo6cLHuITp2oMPk8QYhusFo+dRak4HC8OOPGxzgnpolPZQsX5tBs
NA0sRxh3Y2HOmAw68Z4vg/Zop8M+lmS2yVhi0pEDjKrjL/zFD9pdBMRBCFIqXeuw
JFU9J+sds4gUrOkfJplj4BUSIASw9YJsDCGNAfhDNLkIc7Gh3kBGk0+yqBA851Fl
dnHmvmRmQ+uOJGmQLkKALPrKDmBLfckWET+gHqlyicEZo/B8lWR/c1pVcxBoGRlu
G9oupoX1PeSqP1O0cX/MsdYDWiQ4/4hSiDJbLznjTZHmlx6JlaL6VaCz7zUjuHlL
pHmJTLkq2rtJunH7x7rZh+G7H7uKDvXDhrO3VsIWU+katA/EEX8LplNWPe7BWqUn
oOK8bK1uDxtksVYshBjmjZDaiZ5YE/Vfjalg7DdNs9KxyvexKJTKiodhLvoYxhPg
+dfgAakgNhdi5dauPa1cF5ZO1N6tDX2XlK/CMfyLB+x8KKmwYLg7K7PqDxjPX5PP
WxU/OQqDtttW6APgFbAxrQj2U3J4gywhyNUa0vKsFjuortHprt8wHDxZlhGmJWq6
WwUKrVyW2TfVCBFPVLpMQkmSbZHNIqoZSP9g+HC08Ctamusokn8vadL2sTDJcbv0
hvImF+X87YBBFi3IihAjU1yJDCotEgS9BYPnxWBA77KOcW2zkJkhRqdz+Fg+Ah+V
5BsV2L62gpdWC5P7wcZFDhiddGGvuqSGOVQKWRd1w06JWcXBxEtCwLweuSkUL1Qb
spSIMGlfqvSyULSWVd7phGkfOD1NRcAupeBRK360ot1kBGRccHMO16fMEFMs/wCW
ebCvcgLe0nOfA9ptUmpb/rRHHTd+jcL8OYd/wxDg/RpyI18gcXrDBrJ35L043EB2
QdbZJwPvnF7B998pcV/ISidDCdT3vK+l8X5l4WzNagrjGsV9Lks4KVbjzn9h29BN
+ASJifjyFI6f4lWbDNNfta7d2q20B01RrznSP3Jmjq0sabcjrH5iZLs0uTEXwSGZ
WFt+f1A0TMCGZMo0ZS6VdZzjPna8LlJ4Z7CKWNgmCq2IBO1cHldyoKFExUzkx9vY
GvJqMpRXExWRM0sDg5tA8HjuSOlPwGfmlETytJ5dJ30N1u3RXftJ050/P/zU+Zm5
Kce3uLXFxxo08ep0YVIVgvEV9HN8Aer0OUETBNAFrdZKTNzRKfsHY72cEn8wod1o
cx4rtPbhzHWFDv6Tz1F8Tve7hUCxzfdqGmAPQLg4jI8qGfeH15TOK7DQMhAnKKuT
gECXP6s0HInPM50koJO5G0BqObcEJMxmUepdowt4fWRVQ72UwzahT3cee3BATURO
jbZtuevFagNNhVgaF1wSTnZsEQVvjbelGtSzpu5pMZ8KlNer07XcKq0Bdtist3ZH
XmdFzTLt/5AaxMxlsN/lsd6kiqByTs9cNaP5HCGX7SkwE0kpep0cDSo5/mvkZ7Zp
e+UucTLohlQqd1bIOQzft3YRJ2JWQVM2Z+TExrFFxPhCStDyydM57oJRB4mdhhT4
gML7GzU2dbzaApGzxzrpZYuxjWy1g1G7fSpYJGdq51FTFVtjN1SkrjUQCivFtvzS
y6RIP1HAi11AN0a75d9Dqr40j2l+id23IssdmfysiT1xFNHfbHkb09qGFsfVydLL
opacBPjr9P1qakOX/Uv7c2P1aij4wsdDe/22LZeh4ijF80nYHnA793pm+BBtc75m
CvYVaRv+kRqmwPT5euMkY2wo60EvJChzrjS5l7Z6jSpH1MySGwUBIt57LKB9QsBt
ilbW7g6xvrEBKJZn4P7FMW5Aq7UDMczUKlXwwvvVnToRWvboXQNTf3ol8EjtDx6K
s6bt20ISKUDReS00vNVH/dgg2SAb+2ABzoNkGM948/wHSJzYjz9BK09AgSbKrCk9
`protect END_PROTECTED
