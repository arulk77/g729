`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SdpGFj8DumNb8PR3wn//D7ORqAdo3hUCWah6dh125KWz
2DEe+xkAMnTHyaYmh2/yEoS59IFpyV2F4H1dX+VEUmuJZkPdq0zfWuJYmz0B07iM
mfnZgpVq2hGFR7SiJYxJyeH2YWzlYhgsSVzuX+I6+4a9fANDVFQ+dBTZ4SDNwu5z
5NVPCyLmhapB6HTpA0ei3vcNa1qot6ZG31+/DR1Yh1wbF3neKsB/UatMeOA+O1ul
Vm7cJw5oeE9JS7o26FJI6yR8CpFFZgZoziSArBdYjuWc04L/YSsgLavEJ/M1BMvp
1YjBB8Q8mSN/nLbqJv6BiR9Lv1nSfVW++U6CuCz3YIUgXDP+a0CyloufviMd0BBc
+0srewZWBpd7ujmlhRmHSdd6Mv9I+lLkpSkt43q6kG2evuWqgsU1kxd97QG6nXww
v2ycSvOgJ9qCaeCwY3/FEdsKyyhg1hn50Zwze81rQlJM4CG1DbBM+xhKnvn/O1Fh
Ck+rPp89w58GiJ8H2EY1orddqQ1cIC+aiZrccpD2d+Fca0/vsJhIAfJ4uEFQxunK
FPB+03lCIV/Dt7WXSs+4NuF/zF9x9yOJmexN668O9LD+xTqrtPjvhjsT3oethN4M
frdZ0zt4i619ssEXujO2fFOIRHQLK6fflRDsfN9XumRiOr381hLQZ2A260x+keQZ
lWejf4cWIyb+EsPV32AeatSK8W6I+jMQkzChn9Rtt9Zo1HwpJnUgA8R/nglaULmL
vRju7sGVyx+Gu8fEQmg/5qUpyhK3jGdrhYXlnKUYTO1tKmvPPLBKbiQh8wdq5f7w
xID59Wle10K8+owjIA0jSZoNJWC3tYRJcb7afmxZYHA9eP0zuKUouZX3kv11LBjX
bhfQeBZWCG30xZW1zXFvBaDTfDS22/T/r/KoqmPyxI+jUcMH3zkaWoSc/fiZjRQ5
hLWDr2YdplNZUmbEBSS+KlF/abDxghfo4J/dngfSTO8z4h2YGD3iEQ6GNEQXjX4l
wO8q6xSGNfL3SY+clBbKAf96yuXzNdIHAkH+hQCl2IPRyNgEgNOJjyha9FBREUmx
s+8mX9zxTSr0D6cmtI7jSA==
`protect END_PROTECTED
