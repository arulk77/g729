`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLH6lPwyRc+2qdcz7DnwYyn6yFvptDCEsAJDdSCo1lU4
1rRhlbssShVFa46AGhcGGHqWtqkCtp8rmKvxYBtskLTpBLeaSPxVyta6yUh3SK19
5kcc8ld8t/RJWdmhj//fn18qDwru9BmKhySph9Fh11UpTLiRJPkRw7r1/NjxY6K2
MfFHbtUVrveEvoKDlYoyvaQGitRhs7bj4Hg9QLUyNaxKH3jA7wBo3kXCjAVl41mu
AWeOXMzlnyuMRS8QOkDPigDaoPzMOJQrZMkfudxv/6gzvFcPbdUUkgV3vfLYV8Sg
/76KqvPgtc2UwCJ1F5nCHoDBaQXbizE7QXa9lCgI7pCsWuidcNtbQdB7U29TwPFa
EpqLMdIR5hd45hsmcky+axc6sPJBm2k5ABGvfzpZ3oeaMC6zmlBP7qMXi/LKZVy7
fWcfig/WFFi6KA4yPiad5FBhu/ZYtjGEmldRLrmEBiwFn4KU+0OlvBWfXXw+W1/n
0lbIAt6Pq3gL4gS7n5yi7Q==
`protect END_PROTECTED
