`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
p/mBZCaEdbb6urwLUFHjmBdGPnGT5LRSWlsR1L/qdsBdU+TRwYclxp6jmhofPKtz
Sbb+4/aySt+kUYP6pSmxGU7LjHx4hmyEpWm1RJGOB+e+U6mHNAYZcQfn6mj+doWZ
JEUuNnvlo9I77CMTv0aZTotJlzk3AUx2OXZCzoQn2RmV4MDazeWs+hJZNx9llAfa
`protect END_PROTECTED
