`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJKehe/l2XnW+cKvonnD0WpJuzsNYBIXKM46XDhs09Cs
CkEAObt3wVx3s28Ch7WbogCAXBDLwYDpzwloV7ICAhFkX6nV87ksCxZ9MRFZeSf+
4+804l9AnaHgKxRGG2mxNIHPBjZQ7ogOfZtQBjVr6vNrouw4TMcPNSwX3FyjEu4r
UKG64VPNyyAw7+oKz03uaHn03tmdciO2Xg1NougR84BsT3rildiEMJd8ALMIYmun
Jiw1AJ7xR58oRXQmeltRD+tsdqrqqYl2MWwuI3Iw1gKIrTuMAejad9TnrJh5Ovnv
hbYUtgXawHQGvc0D6pYjXgcFO4YW5yZ0phBvoABFWp95/DRg3MEybmpoizvt9i0R
xnAE0tSus5U/1qU68Up1hs/0+JdC7pUC7upQTwPxMHEArixpX3bvsneQcaH7+Cfd
7bQOb0qY2fwdutQiD/bk+HBT2h14MPLnkIabemYoz2D4USa1m7agoL0iKKLN9EhF
5DBFcb2RD21O7FbgYCR8tSzuCxIeYeSyGi/E60U/UzXREPdJ2AsqBkWJMU4+v/GD
mchJEuEIeT0EnkUfDOilbe2onJGDeMir0xKwFThAa5MoICWotUiRQAmSKqtpLMxE
mRPH6t2A4ee0OToj36k9nfoS+/RulXqqsl4Ms/phO+aMd1jqXg3X8kgg9rT+H5Yo
z36qbjaoaoSjgFXfGj7r/yGuN+OfHqv8W8P90jdCfeR+LaGNaT/aBgabRmKPBmIC
DYQ2U9LvJLcxP2CsD2kedydZ8SxYOPXebgd8gLqgzjA=
`protect END_PROTECTED
