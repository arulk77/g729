`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL/o+s+PYiqOlV7CqrYxYizjUozqXYCyAImHD8vU4IgM
ie3t6i0vc2axNedM9W70PGb5L8Qo5vsxEiVl8gu4VXLaEY/a3lsAa4SnJHUwEsKg
u0bc+AI2l5E9zXGQHbWmwTV9Nbhf8bgy4BJ0AZDNBcdVSx10m5LiP/fqraUemYVQ
5Ct2M/9y2wI9AbLuh7H/2tRc4cEfz89bu46xuZNbnzss9MzeiRXY0ziqF3JbXWr8
u39wwPfmAKKF8jVNzPtV4ZIflnSFtna2sEMyIjZZwUQUIsrU9ofrmMAY3AGH0b/3
GuZHPCEY0ulmD/JjmwJTwA2IuLVbGDT8JkJ2Ogwyhe0srCVAeiETRMP+bLF4HF3w
w0Qo2oVwhJPTpK3PlqqAAw0KczuV+V6OtKeVqP5/X9FgMo7Ek3jOw45F0kb9RjtG
lmjQ8jG0LxY1HZjAzVoFBBGNiofNDVYh2osGIAT0xZwvi9QHOLvyHAHmvi7TiOpa
NyNXBLalrh/rfGBsnGl8j/OaeifUho8M7JiKmvFnUqKurdgdc3+94xWaOE8nS6kb
GRIFxaWsYJ+oqKEZ+eptrvE6mW45bu3zTdxCE/eqkEjS+7R8+xL2CWJ0c2euJXr+
J9nLrrzajCOcL7DR2zrxsww2EeQrtaHV5cubgyRQlVb1CA+V/Cscae3AuHYosWTC
ikfMi9eozB5h2T7Y6Uj26FTdO4Q8i/m1chDwl7aQ0Bo/qp0skE4BGUYSO+eHpWDY
mBwYftJmZrlZfeZYBz34nNPXoxRgY5+cJtVt5oa8rxpw4XRWpWqpdFUx2FmGHuO/
039ozNFXJhi8XfIfz9xUl+QqZX3ACL3D0PwIDV5C9EMfckkvYE9AmriLNdrGstxb
tTC9IfjwUpXDcRT5dzKpoz1M6EzrfxBzaZrTvUX8hMmfX0v3yxdb3RaoJqmSlPjV
XpefeB+b0Pgr/hI2Iwv6EwZFYxK/WxjvDhcV5jC6JW/08wrxibnENdCOwoOQIikj
CCQtMiP7AMQCRCdQuMB5wR1lsjThXyKrV+WFRdy2dHaZC+DecwyW/7mcaBzcrrXZ
EFpEZyx24vD9iOMUVTYXYjOX+ike6iD4zZ5/NwaT8q3eWRQoRNBpqIDjAxSS95b5
Bs2iJrfLZEm2FT5SQUgn5pnBFO1blD6gYR7dzr4/ujd3V3dKB095CDQa6vcrd69I
oGla55H51Ix7HPQQ9clrw9FK2Xk5hWQE+zDMAr8akn4UqlXXNPUroAxBYI0MsM5h
AQ2DcXCKHBs+uIpzv6tbSNCLygY3V92aiPejelF3HsGSHJsfFkMmKjL0vSjC+4f4
YOW4X7dNehihK5Q9MOwMnZUvrh50GUO+XiwgKqdx2PC7qlzMmRln1jcdo+VnEX59
VQ0VWNCO6O9VJ12WE0Rsbi03Kuo2qFC4Z+NzMBIYxMd7Ay7UH7tGmDoRRjF4oOld
0YCtcQCWhVmTdpqWQWdm9Wd1zr5BaanrbHmwXBq2BcikEIWJCkZgThh+/l0nO/Y0
Bik9CmZ/lztP44x4WLg0HOBaqRkTjmYbSGrWTo+iO8QbnUK7CXXvBFZ2UIVEH9oa
jFBvr9nSv/vEBhCniApvLEIhU1B1fPwA/A+hM7flJsaelSJssEk8XBt3LHk4Hhnz
82FTxE1V7VwVv24jq5dmU9ksfncwlpsfSR9G3cJ0OJE++nFqqunfyZyjYANIs4Tm
aB1jc9kBEYsN+r1LFaL7bG/TCO7WAcL1nCxs+3o5nm0CcTSmY4B5CWgAYiql23+P
s2zLi+8qb4UQ8g0Ef1Quld4yzTeyjDfZPdWmwJyx11An4AsgwKcxQoQnnLDG5LSM
bs3Fna7U6+gZtXq1M+lC3hQlBn/jkBjx1lXSWNewUnbXE0MlRGPRZrqbZsg4UyNw
a56kbwoEb+RL599SrMy2E5lWAtAC4x//cDaAVcFJOJ5tOW56/9yk27M0+NKAZY5O
R8o1vVo2F4q4ztATJZgx82Z428dlihueHES7uBSoIJeRE8IPRnfvHkGBubg/kVxw
U0gkfr2UgokCVexNYdcjtexTIPd8SvHcXYbKbpKBtFzEXjmqJRYCuCT45cZCi3o7
l7jEk8YKODMeQvnjFRks4pxP3XgxIlnDScsdxuFnsY5cw0A57/Evrf4keLDQfswq
QHx98VkfsNlQ6MEOlkVLJEudNA/Mb23nW6RWl5y0FzIKch3r7E93h+6eyWQ6yn+G
w8c0sDANYmeJb0M3+IyVro37mHzjs9rybviCJHzJKCM6vOYF8pRZG1aWTtXjgK++
/iSgQFgzYCtZI4+r0BQxjMwJZWzSWz1i2e/zSS1GHXfFfcwZ4SYimNjJXPqW/iYh
Z++SR+EK1NyohprCTlzTBGqEbSCe8rZALaVH/Vw/COexWqjfCfUL7lVw7l+Ropmd
BmLzL2Z0Gkihi1RoyGgDs67ojLMAen09FSlrBfUm5rCW2fh8Ygt0FaU4+BW7vMBI
1DrDYb1why518UyQ4UHOBZ6wwHu9LKMA4ybPihu4LVH0xb/MXnzYODZ6852IgXuu
e8pvq4VSu1lx2RsmWmhWFJqb5PnV6tcCJpcppfxchcegmtRH7IW2wowDQa318Pg/
Bm/LvyXOndb0IeAZElZM94MVm2wEtXZIIQy8F3Y0rXWrU/QJN9gnRkVliYCTzxs4
/9JCalxn3L8ErbrD4m4ju6QenlYnwRO9pFXkD6NzComw0DMWxJMPxED52zphD8PN
lKLWwGRRPh1Ldcpk9p8QrsCv6T6EMUXqt2MUIkKwgPyUjR3dEnkJhaH6/g0ODKDP
sK29RfFqzOQ8aD/EvnsGXBI4iQA1BwsrOIEZtwOXGtcCQwGopMx9IFfqmFT2Sj04
o+BHbZZcVbkztabMOXbsmaekp9E5y42fvflyIxn00ZAuM66+kWucN6TH0tDTlTKX
bm0DGWtnmhKywF2VwuC458iSgEYjW7YcXLpEnYr8XiDYueZPG+34iz8TvcI9XKDp
mKuhH1BR2vEixCAS0yI4c+BhsUBaJ3Od5u9POcF92ipfvHQz46+3e06I/N27HCfW
+Pcz6PHcvFpHcjqdzABQvRFoU7hgWJnEfrX2s9pVIn8WQq/o+E9o9TZNQe1tm/So
lGFtZeQUrXLcmDdeCR/dlVyxazyY8MbrzhWZqL4mj2jS8l0bNHTFQr8JPp3ifZ/T
4ql315QMZNFXv0+YHGSlcKL2qvzykbtxG3oN+2c+eSunQpdoYUCDY/MXsRFY2gPN
n7W5AlCY6qdQPfKGQU3/EwTRW/QhYDBeXzzx8izqrLlH9q6gjZuLTzRLScl5Pwgt
K2yoEEJyosHJQbsMtZzQEtsgB6JR0mqvyxkvgT7zAYjHKmu5PhYRTPGOmNopWL5u
Eu+0f6kjT8Y+rbvgYLVJWW4M7f7r0NKNdHFnSA/u7ndT0JPe8yGD+edtKEh+wPM0
qwGuh3Mg30FIqgLlr3TUqg8jOqLuAmT5douGjNIBT6Jn6VcrtxbKRWBKk12WjNx2
fApV4uoSDC5Hhyqg7kzCzIlLWkiEP6ylfGtFLuFVY8twXQhWgJdQ/2Wu6tS6Wlb9
4NxbkkdObb2yvl2Cl+acTTHjB7kKyxRxmiheZCVcNyxqXIdRRb/RXXmJVJyeO4Hu
mvKM3oWToSnh9jCWIlUspc5bQg28j22av5CbWwGgd3AkGd/9uGzEulDXM/6n9lmD
KZjagX1+vx4VgGHe1q+tfEg5IIxfV0eOCI5MFjYicV5WSaRRFXoOlULRqee3+Nr9
t9JlWwozE/PLdJDgRQVhpx1UWwbBleNufDDl5H1v3EfuH5Gi3mDbA/cJLwN9XKvz
TU5zI2zhHL28rI++lOgRtoJak17k+TBw2SWr9i66blrIkFc5PXuZE0sAV2Egzxk3
xfL1oiRiuqME515r4w90o2NyXmwMbpszxc14JIzp/XiOLE/8FZQQYTtjIuQJ8Ysi
Sbt3cRteq5H+ehMSLv0us8o5Rdpl1C4+4Swi0S/u6jQKugmVOLc1aRsmvuSFWuRP
Jv/u5gTTgNRrwi3Fy68JOYkAA3aG0XZ9YHlvCQWFwiocAPkyJqpN7lLYOU5tU7I/
hmTI14qEzcykvJlxfVAmDOA75eqju4sdY/H90EwoASVXMMkAODvzAQH06sE66gnj
eeGkDoU8/Xl0wucUZ1aPZyiOCngKfTkT/dJxXIZpPd4PYHJr3yt+14jB9CyaXzQm
DXu2NDN1lv/ObcXcgqGVMja2PMWDUivcw5EK5vPvaMMQZLlBMy/09d59L3sZniN3
x6Lx7F2WA53rsefmPI3vz4ZVzM/jZgSk9KiEOAILdN0hGiR+/BG1B+CylLVKvpbI
SNNRv0cRZn+w6C8W6jo32TTE3YtUX+KY+qLM1IZwrxE84YoVlgQ4lXW8n4Tffv7J
42TCkfWFNhEnpm6w0jv5GLZvqor1LAbRPfLcND+EtQEKExUve0aQWeb7CBfSew12
jV4SRnpfnhKOsKNBaR4yHKnFd0LFy6BQ8F7N8d4Mr5gYuamQy99yrfBKesAA11SX
2/uTZc/c/Gl2NTv4Qzj+2R6lwQB/T9d0sGoXjLfLPNuncc4c6GCW/g3RaoTmwwil
9+UIutDn5ZGK1S9sT5SQoQ7UPTYs4yt5AYqBsmt3P0tWFmj/30lMoZkvEWrrewVv
a+B7JPZsNJrjvvBar5DzBTrQ/MA4devS94v8+rJ5HI36IEqvZgQKKPf8HIdmvnM4
vDbtikxzadxgZy8USd5XN5Wc0Jzy2YVT0HiUu+mCxMk1C/AJnICKzNNPH7zeQUyD
rdzMfjmQ1jhUHKJdqp8B3xH4v1xShAqJuQj/Y3V9Gf2U+gE4bPX9XC5LHcWJ7ux6
Qyv1OwXeWqnrO7B4V/dKw/CKsYuvcLH3KJm4jiveQLSiE7eMSpclDYwzkXQhOnWB
4DzNPBjQb/VWeiLYb+f5L5fUop6uCboGWYvts5eeFvJ1E/BDOcM9E+tsdR7Jx3Dt
wWcTSaP1aK1p0cE4oBarBL/0XORhBJOhvsuZwmhaw0kAcYeX12omYSgmemuudaK0
IBkcnDQABO614lImT4LaQIf1nscnbKJle4nQb3ZrmnlmOdJ+cSCmbe39mSS8URxK
fj+/D21xiuuuMeMiqn6mwxFiPnUg3RSGqiYrv68Qw7f6Yg911HEBPPO2esvQf3Bh
zXn9LjUtSCaQzGtWY5nXkiLPyUdXpy5nsdKX5xdffQoRqL9kqXcvpaktLQiO/F0k
RsTkCdBaXZrXAf3RJzw0PLDXuxcBSNKXacgtfs6ayJs1HW59m4HD/+RMVOzka+PU
/IMI0b3Smr5Yey8w2ssmI8B8Dc21W4bc9DFbIT0KidU6yf/ENbrlxTC3AIJ7SGIf
o9f0gLtZ4m7SVF2xcTCJnntwx+b1RcAXFsl4sbrI+1KbMuRgQ/w23PuQ8FcL9mMf
hIFDvWYO1RpcWrxrGBUcdeNIlvTRLSnOnyCqtwWloPZ9hGfQQ2QIpteZKCfkna9F
O44uMrbzq8KqT54cn/R41bYawIm2tpWn+HdhshQ6He67PMeqCZI2jAZ50uwVzhHO
MIf2Gv8Z8icBPIbMWu86FEFUA4qBS/R8/QlAQd+WMLnI1z7EWg4JNmAXl+M1OMRp
Px089p/BHemvw+zIsbTNP441NdBdbY6x/Pin+kbuDJ0JD3ivaYOqtfV/g5rM/r1t
OYMKNgTnTb4o1pn0hhDHnu9+F6AFvmNGo+0W+3j4cdG6i4ftyB7Azgqka4C8K0Vw
aycpqdDuryw2/KGJbpnmeSlXHUE4DbY3UW2+s5PfWWFzUDuCSuAAm0tH8P175usK
KkgspuhGK02/c2MjElxOtpYjIdThzv82/g7aWkoV9tD0jFGFQCBYnMgcd8qOI+UX
eAt+4YVuppR0miOzykZlL2HQs9n73R+um+N5AmMuCg1YCKviCcStJL1UvDYN/oCU
TpMugD0i8vvjorZtX/9iDO13MOjkFR6piGy0nwX2oYXuN5ssztHh2ZnOqMSx4Ryo
OVvlIh2PB1Z7efvfckoaLVRto1Oc7WvX/sHcgicr2AUlpz5n4NWDyfst6vEoFCp0
vIj2AEEa3jov+HFoPvyp+X3Wa3CCq6EA/54N98qy7QdlOq/7/msnu7SSWOgj4TCv
DJQVjCIO2Ii0km+f0JVxA3yzffNiUX3aaK1lHw+dZtJmK9fx7W4eCbTAH8tAE6x/
JmGh4uzn0eSgXlcUv3NOP+ewRzZWvrJv4yP3Do2nYCyUEjk614nEOPQBoTEh0KPW
m+PkgwKl25C963YKFSYxVu2+aKIzjamDXr8R49IRf7uhRypIhZFIUldjc4zgmoKi
/dCBI/rpcN9PZ+bCFrlTYmBHGvW5RYMvPFpaIz6Lp1YPM8Jq3HwdrVlKDKhh4ky4
A2ZQbLjYsQLGBms1y74Gqt85XVJA4yPgAtMf1eNuTzZgP1s5+aY9asz63xwav7Ze
qSHB5Tee19RXY1kOtRDRZsMr0Lbx34roiI1uyJz2BRgFhHB0ITGKv/eTs/QI+rK/
MiaKqwpY8JkQ789vG4Cpeks8/LY9LK7NR56l3PyH+x/DQYeE7Iicz+eBP7H3j5Mg
urdpj9sZGXK71DrEJ8lpHZSokjzfio5JwN/tqQk7wYYI/SSBpfFIHszXRakfKUNO
d8ybS4H2CD8chBkddF3I+mG5ilA8dmfhSjN9g+gDYVCftFjLzC2yHpfod3ZGjU1p
1E8peqHqCH9Q3qlTos97JE2s876qgxur/u59mUrzqvj5Fd7jGpvvJ5mmXBzAQagX
TMqF04g3LA4J4JAYNMhGf2VJFC93NpOMX2EODtB44OjHhMBY1JKesA46SHDRhtyS
AfeU6BMJSVOzFa23P2HRjBimgcrn0UycicDgmVD4QOh+lE+dxFSnsPB93C9o6dQH
VBeQ1KTN0RIJ3iyi3Z6RrQJ2VbzrG+wRk6RF/ItAH5xVTfIJWQnhnlf5+JlRk7ry
CAzaEYMsxqsPiVZzunJXXvv5neXZoo1QD9M6nZKqZxZ9H0x8QY6f7UIJz0RhSf7f
d+r/9N0C6XXnC7EOWNauPPXF0ejTNLcsho/7iGGe2//GLVV13PeLlYcjQb/TE6IF
59883lyb2cmmsDbEmkwcGvDk0408tUa32vwNTEkgEj3l1dg4Lnieng6ouIElEhPH
1KZMHGvGUVzxYwCreW52L865/hXaLl/DFv+0OTSzqnno7UOSl3LhHcLIgdjzFc14
k4/A3tgE3LMOjDclq6nZfpKUcy6Otpp+v0PvBLfOv/2Gw59voShSQQLb+bvZolkt
E4JVpwuZsGn6iDqxZJiup/6D/5Iz05USaXjFwSSi/Ac+zfCfQ/h+TJ7zb8xlxX0D
+koVGfBDA+Xt38szBdfiuh0fI2q2+rRLG/1t+tMqI4LHt36TziK4loYNwkDEjgy1
PKlSBLh36M+IGYnQ4pyCJC6RBHuxJrJaAvo5/Sb5MGQcBYRoUM2NjO9coxJQC0mW
RSJO5cDIldfO8BcX4cvRcVgHsmmzM3AlSlv0uO1FYRt80AjcZ/qRGV530trvCfoT
gsLNAdO/0BNLu+uP9VLX0wPp4u/fuHWk4fH+VJYl8zK/a9xB6QNllZil45WNcdeh
vZcmf1Cxxlng9TxVelWpeqOn7VxQw+YrDjMcZH6Y8EnyTeUa9WYmEK7sP+Bs5i5K
3FRXvk1jY2yxAf2lVXtKRIGMD9K/B4KrSm8rJCaBACVZ/+zS//7xJxgy/Q7Qfzoc
iAxpDXicjtxO1pLez9xkU2GAFvZ4hqLYwNeiHv5LxRROVnGOssDqOav/GuANWyBw
TNPW58Zzv9UXTeB3u/uyggp8NOvm6h6F0nlHYqSAPt0TNX/CGi2Yh/iRu6fHEFo6
8yMZu9546dJ2ArkIf4POp51FRvY5mOBgo0UwmNickhqL10yVs2Wz/YXc9KSU3oQM
Gh0j/8kLY5F1PfSVik6VVQqKm8RjPGee/HkJUYkZVm3Gy7dkQfkFpLE6dO82xPfM
DV3WgeKhwljBi+zIe8Eq10dqskwRq8wH2XvZviD0+jWxbH4a53gTWyi10hdqDCQe
2mrO8lapH8s6KZZyOa6xC+G/cTDrcc3eNYBGhbFi3Vx77mLRCH3G6l1wYdC+3tqb
2jywZq+ZkuJsTBEd0Qcb50AGYNbJpygJINcrYQeg0PijOTczD0WagpoY4D9fpCz4
ntpPtmMoiC1SYfL2Sxj3tikTmlS5EXDLxh8imPq6jcYBAVMAhHI2DO5FJan06CuE
LX+LxLzpAEI6pnPGD4VmrfvW3YRocdBQ8zX/n0glONKAQTsCeCXMP2Glo3miG94F
CRe8KCpZoXdbc+6tSq+OsgMS7W3N6b3poXpCxWZGMpVQGMjhsaUvSLSgqVtlFzBV
nrVA6j8yDFONmL7mUOIGGxY5TKANYtFJgu7oP23FMvIeiZGmxnyfsG2tDPrurFee
1uHPacsLdIht/hRNU6+fo462YH5dsFxTQbadb0Rvpvaa4CY5SAy8Wcvv58ijTARi
4y9rwFaB1oh1iiHp1VQwG6i1uVC4RjUBNZ4Pffh83Jy8Eo93aosmOFDbBL7XIGO3
El7y8e3D2ok/bBrTSIeYYZuaIQWY7O7vP/obKXqaK/Dt0l1smno8ITQgQDWhYPMx
mCD2qixBMb8hNidv0oKo6ittDvNL+GZkZqumjU1nsdUCv+hv0tgAtX9J4MhjwCzP
XPDpoTpYw3ji7aQIIVCJ5fvPd/eud9jt70eoT2IpBUgdooUP3KgArQ5sXB+txk/C
+tYFl+6w9vZZE4yBovLMnNuZ/Fyzu1Ao5DvOjOLcWzO4MbbCuVirF7ZIn5+XEQ3V
vhPPZvbe+tFP8pvM9KaLPEJ/5yfA648pzfzzGtcsVpkOjToDcTIBTcZEtdQF+cYe
Bh7P+8R2ar7uRXyFxYjq89t7aTMYCqPMS6t/STTXdzRNULy70GPsYawFYg1IgRH3
dxqWrIzDOlJ5xksPE/pBBXNjDMpRChwq01Mzp6Lc9tZk5ZwtaiuaKFdX6FXAX5BA
FCie2Kw4kpU7ivWPPjDNBwqUOGnCXWxOEGfLzEe0bjZt1yyk7y2JU11PV45CoNx2
XBkXjJTUYy6c03ODIuKogcXWeHO2gb8xF2npVSabciUe40prDF8K4gkneiSUz/AG
fg9YUboaunkA8pWXDh4tow7A+UbuS2PwHX8I21oka6KRLytTwiQoTCCu/XieWll7
N+xbx8SqAMLjJBPi1mL6T5xYhEK63OL6PbeMc79vdaXbbYEMK/o1BgeDCxUpMnKd
NTu6XOAMxs+Ja3IS0kcLlHYHLI1ccoCvetkJZpWExQ+uDn9/sVAW0QsIuOJDhk/O
YZcP86PfBYU8WWi0kRm2erNvS+Zw1/lc0iRNBFp6ZJKSc52wRqWKP1XM4cg9/2KF
dwaVc0fYZCXm9Z3qDd1UrJvOZ1aCCz4EaQwEVphZEaiBR1AyYetybgCV6wdSo+C3
f2UWrjnp1sKMuapBaZGVEtpUW3+HAZX2fR0liIdL2aQUNrQa8x79AuE5yoQmvWBN
UgcCggEE9I5OiN5C4JyMRqFIp1JBJAdfc3wjNPGKQ2r8xnbZQP5bPgPb+33wjb/B
Lj53hujC+7gv6p57tVDPhpk6V+zCuxst5n+z3utUxwCRzxnjtOHPUObGArxdZzYt
vr/NlcmafmJCWx0PHRjCciptCxH1Y4AOUmAAvXC2hDpkj5MXErEzevzZbqAG58IB
Q2sUXaZZ5X6jVc8ZgQ73N0qL9C9IOTCMUvPUzOkJ4RwhltaqVQACYr+bCrgK9ch6
i67IXKhe1UiRQRW0vbcaw+TspvFWWvcYf1WCaLEKWq1Qz5opWPqehF1lDXOM8Hi4
o9bVejHdMI4NnxMBOs2uGywyCBEidadVG5thTZZCN8//d43d1i+C6TyBOOQX+vyh
Rq+qwjuflsq5x+W6HbSUD9kleeN80+5EU52bG7jJGVlsLngyvT579QJJLMYE9CH6
9JQM8BkFcH+q3wdr5bz/RnaWZNGX7pdcO5GnaaBnCymDUXviE3rnCprxRwHSX6Eb
ebGiRCIB7TnPqC9HIQhq+E2g4cdkW49ed4kj3YucU9vnTuzJqSo5Xjdwt/QnD0NP
uoj0tlukYcIdCSFCByHd3FJKaYQGS++i69rFnaEX2c1PeRkVFKCsERmlaRBAsC8I
Aapv4m/PYLkLYa7QbAgs3a6shkKA0JX88D5Jm82yDqkqGuwQP4jOCdMhgFFQfZpx
bNI2LKT9lq+vFj3CMXsZiveJAIFbvADbwSOL91/iKcy7voJFJM7VkrSWsgesE0iI
xqZ6huwDNfenbGrQKCPqo6sNgqjhwGPXhR8qRMcnDOWHvKV5U4S6X6X80fZ6U/V3
x6R6WcCXPDI/jzukf04F7r5N4NfI6G/GKWZ12sIzVJK1NFSYL4wsD+c2kCnXbmy6
H9hUs/7pODJ3s8XkgeGYdxc0PqorXGhIg+YbDph6wg/+DR6XSjnzcN2udsg9baa6
kzZLEWWioNDp7HYpyWnbyivOh4NAmxsJXMXZ5QOIbjzq6MHl65EFTD9LYjL9uxeX
wCXwXfqa8BTSDP/HWSspY+pqObT7/ANc214OtUPKYMeLyxn6+vdRJOEaQ3Z1IX1M
P/TsSIRLeiJdFRmp6hArCn2c1rf0EtZPraV3Z5MuJH5O0e9b4Vm9Ynrfqk48R04o
Fd4lBfCOsn87pRrqmgyFgFaZ4JMowjWImBLBkGHbysSdaAMoOZSQTzLSYc/gerNq
b5i33j5Isc1av+frxhlsBA7HEo/jTVrcNtpglnM1a2+xupKyiCZEFXiOE8YOWfre
8p8vDJK0JJaA20FZsCfP2ECghPNtlf73/XxDR1liC8IMQUMSLmE5rDbf0rFwQ47X
Gbi9usq3l2a74LmRUHohx9b3xUrBMsRChwOyoflP+PdZhilRShjc+TzMDTDWNhF0
73y+3shBWSeptwGXOjJl2tbrhBSiTIZs0ainGzHshW6yi9sAr482T600bJEfTL19
P6ctPmNl5Qp4E5QreHHRoLttpvIixKO5p/ZTnb4O0uvsrWP1f/UAVjE/Sv8k5R6x
tyOK4xSL4WcZ5Nvl/wHzSRukME6nd0bwBKabOXckay5wOMUgYeGeXoSOqU9B5AKK
QsN21D12VoQqrKwukMFVYRBDdEh4LsM/3RkCGib0a+o+/b7CsJ8FIOBKMmcWyGUk
vgCj9jwGM27Z9/GbCKKo37bBMNijGFsEXUVDfsRZi2Q+0G4fuDffse4b1FEoQTHE
WFAFWJFTaqreW7lgONh0vzrH0lc+YAUroN4GBQPK+Ubwf4T1QuSWQF6iG5bsD7xk
+fXYoTP0k914i9x9BWoKPKXbg51bLVasmdMvK13u5NUu8+5RX6KaX4bS3qpjAEWX
8foaQobJT2vTE4Le6jxf8jpqBb4SKYrirKCQ6P2Srs5SfKZ9sLMzIADGXzeQrYQK
PAi2k2oH4Rz6/NiYCgcz0rGmMz195nKE14mcwgP7zAentI7WnkPpawiMsPyNKnO+
6xsAbNVN9I+YCkiXHgckOaXei+tvrJhglo3APDS4yCwj0MlH6vSM+MGq47/SaN2L
vF+QkD5sqENRa7+zd3Bp6sUm628Mwuu9eGocPc1rtNU1B2+aSSE5o6vfJpqLmUwk
ig3uuZQTYp8nFl54ftEpJlzz2ofF5h0poeq7T4eC8D+6yolM/o9LB0TrcJt8NUml
F6znlObV0fKqoL130omqLjdZms+7kKfUdMFRFnPo0S/gettseBhBOOlko1eCAcFm
CZbfimJze3ARdcH5g1U0Wutd02TYP2cyGiZpU71TJULImwBnnD6KjydlIzcIgTrq
QMdxpL7XE8Gd84osAWtUGTLiAArPPwJe3A5SbAqU0Xmvo1Lfsq4gaIQd/rBSJDMk
geUUcau16p0+s5Ri8jRWE7MOxlZz1MtM38plgsdfPqbwjTMGgdX5NHpDE5GagnaN
TGwC5eotZopOvO9IjNjXdVMdgcbgCjn8tnkr79PHmcXHrsPKUjDC4nKBqWDn1sRf
HwA+Bqrs538cKRnkcfR1NK3T9bwsLOvJECyMh+mAJThk33mfbc6UeqwCrDMj30BC
0ckvsUYcWP0SEuuBcfnmye6ZOqVX8pF52/bhyKbqYkMBsibGIJMuXoYPst0putXC
KB9FWp/6wExNl4V2zV0JCSKwSwrYdG0OCQj2ttEyrxZe7WmBOou2Cp2Nq/ZE84Ib
65s3mcvWdGdiBpmvZS44Q5GY6OOJrXrgQl2Ota6KWXD/UXoZozzEcbrwYBOrsK+e
5UuwiVKJUcWDnfo7v5125DoY6kua2DDk6puyvILZ75NIeps4ByHVzOYxoj6bBXFS
hxzZeJiLd44CV63Dccn2bMMtTxqxF+KWDFJfOG1hskrdECk4LAMw0z7oogpGZFaA
iDGoYxSa2FDQPi8KoObFmPBAsI04E6SNpf9BYGqre29ikiYtvgjcfdw+LQqmg6iC
fNbMOXsn0ztUMILSUdkAaeGkp6mKtw86CnPuZh2tzBQ69OBwBMHKKBVSgRzXPEvg
DVkhnF45Tm68D9p+wHMJOFzET7D9JytrM3NR7M5BQiirc7SpxyL/hBry+J0D0u9f
BreT0FbmZ9zTJi+TfBGwUE8FqhNfR79N/AOrcrIgznI5YHBKiF1UB8ZXmoBor+ES
+YoNrmiIluadkbGf4DQR0WJcPQOGG1M/aYUzCDii8n/+Cfoo+A91XyA340SVeRfM
kd747Y64YKwIFHcgg+gET4j5/yCpLTSwo2GA0AlUXqtJf2/5TGqoP41+kaNq89YL
1pe44vEmxjFng0ctOTYbGnWGv7RjSxLJtxqRnUWdLB/HP8vA1HnUnTXMnywz+jPF
iKXeeutG2xlUc1Kz8o3+RxHvy65XtlyJsh58Uqj0hIILKp30zkJncLY6Oh2Dv4fP
K2QDqkoL27nHQbMvitGjcicuOguAC9Inua6hitSmqXGYAQINMF2GTwLgZphXozdJ
/Fa2loUAuKfjco+A4aK8l9SEaZqjmXAjdsESDvgrmVZAVb/Rvnws/8FF7xsxQNO6
L8Dh1m78MKsiUIngQYEep5E7lsWC16PpEBGqj8fbgv9R+pNZATc4DlmUJBQfwTxM
SJ+MH9v7KUqJHqEwzIAmhuC3DrUPljkSb63bUkV5UwnPzXaQJrl6rMhvqqU2ZfEH
+FQcB0aNOMSIWcnISS4orBUgbaOPf+AiK07GZR9q1vgzkn0S9fHh1/0fKmgLmr11
IznA4Zcn7RadYj+0dnb7KOz2MU0UJvOo77oQGuLxaf8u+8uNJesdEI/cXSH6ZQnR
3evMc0un5Ml97RoW+JkVbNQDbeaJIgfgdiWUzQSRMqj7x+Nk8t0kjKXQHZsKIVd5
obV2FzYW+nysgcChvDdtZhF/tn4axW045R08Rhwq8ctZNzXIJ/zrkGv+JnCUfgKY
6pZcouxSX1qWhZpLvDYLWaxsH+IOnYVONhBMuDr9rUalyWFdb+F5czzJ1X1t7lqR
MiXEh3/is7vhGGst+dYBa98Bji3CsMV7nx5IhqmEdhFxWe7UWjuF3FOgwcg2iCIc
aRSzWp4EiO+XtgkoyF2djw==
`protect END_PROTECTED
