`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43Nr1zAtJ4ZN0Mo32KdsgYKbBQuFFiboFEigS2PYrZtn
bzjtg6ciptIHWv1S42iMEG631EvEmgKk8wOyR+uX4wTGRwu7d/0rEBBeIiTUzpfA
LBwpCgDyHPcqMQvuGr/kxKdtHcKesNledMEQYGGm0Vw5pTDxzr6qWq2coMR79IcD
PvChdLKzHsExn8eY1mX7oi6oc9JQ5U+fx/SUY8oUVkmUPdwwknzspwaReWAK39mG
1SA3hiKaAo2t1viLFpyD5QrYVhvosUvX3/3CgIZ/c/o=
`protect END_PROTECTED
