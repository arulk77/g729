`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHQUi4sofP1tLzt1MChHJuQyfbhnOqEgBu4JseQerfg1
qGUcbylfgD7kLhzjco3aDvdu2YYEJq97VHsZWMzG4nfimnVV8vr88bMB14FQTEt0
w+bTz9opwLGBU4dRvWTm8v0cde1qqciWd+5HHjawev7U1WD9j8GwYcSPB6ibBG1i
`protect END_PROTECTED
