`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAr+W7OvhTcqEQltWuKVQevyQbDsi4SwhjfpqBIvhXKg
DDU5snUeSYU6D8+aE/dX6/UQwOD6ettBCWUpUx6iS+UGZb0AsQplGI8/uk+p/a9o
UEOlP60bq4Om0EQBkssnPb3vYY1lF8GTNV0T/GmXV0tOVBMtTDYRRPqnOoHgu9of
pliZr5a5qDwrXimOBZRiercyXtxuyxyGc1sYUXhTYxYuKAIh7+tjskCfpYDxpqDl
`protect END_PROTECTED
