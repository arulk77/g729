`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ec6EFqNTOtehCYkUTRBJvuRNW1eZilSCvTWR+/KqwYiuRj4HNfYvXe/SaK49tBHn
9K+aqaDbdf9h28r9JeiNVdqo0oE5JVW6YUnpDuOZv1iScpvgwplcXQfaJ6m7SdS5
QfBeohzQ1xDDKsvTTkPoKoPPW7DQ5I5vNOKQoRR26BfsBPeY1DotLvpXUyDG0qMB
1uITFofKcgQocp1qwHJUImfpdE24TN1/k9Z4QKHAL09ZBFyerSAujF+Y1dTIGCy3
pO+DTwJZUtC/8q6esxPrQi6hZ5UXCurU8xz2dyEacZmv0BqHC3zQw2VyP9pB1hdX
/N0hrKQaw6mNFcmVyqVWMoFlkvL3YpKRWpTar56V1Den6yGup/QsNteCh/70Rb65
1FxLxyFcrwcsWg3OIotYdYCn4f8X+Lm1kPmPIwoLxv0Mhhggc+TCVCQbTXsLQcQH
wsBDzRoW8t/dZHDfkW5eirabnFyA7R1S24ywfOlot5dDs+o8TGSWQZqWkZOMhQz0
XVDsZt+HV3SEz9M5qYNijTyMXmqDUhwbkUxYLlUfecLUOmN0d4cw+iLRR7zRkzip
tYw8izIjPA0mt1e6GzWKOzQsfXp9ZijO6m6oX6kcohlY6L9ZeSRW/QQWqwaYkybI
0KGxgvfXVSvlAPgged3JeXdQ56DUCAVnTFsDIzPczqXCT5JoZoM0wfnjsQrVpotP
8EHncKLUHXTyiaAX09klyh3ut/TpbicnzMzTEfcd+InmNFo7oOI/GVlYXglXVLyv
VDBPTiSqvb+5vPif49l4saJz5CmtSwyWAVLUHqM1/X1asHizaOUHmRmvA8RrUrvi
ACugFmDOhzgCbN6PkQWOTRapEyPIKANw7qgJ2WmVTt+0AeDWIFiXA6Wu/6yOi4nh
OO8fAKd+loS0lgEb9UoJklIrZjxPhHzNbEH4WqPxligUss1ern/bnYqyz/gpYUrj
s0pOa7piiuIOfFM3YiSsHnykpdde7gaAUCCY1qL486lAKFJ1DbOFjXs5KstNljx5
BZAlZhINvuMlIGqa5MfyfbcmaCNFzTfllsewvoDnseqFVXwwiLpOeODNqktlcMZP
Zw6EArqhxjEnIX3hefgqtit99JHwsjtqpAlzkZEJgBS2FvmYpGVRTFNY1aaviwpk
Gdd2Oo7u46+i6dOdeS+hVkduybx0eS7D7xbaqh3TxLciOatNoiEvrDaXO6CPkf82
B7xL2Pgi2/4PrWl7tdMuWDoTGHbN74mSg59eVgvfAO2Ld4zrIMFvupqWqTZsa4DM
MbXdGRAh7I/+Y74/7I0R3mfwH6XauLwjhgDRanZDD+tYCPGlRVl72jLi4aUBhadM
yXMjqhQ8UWPASdONPq3WuHtsjBAAer9uIk68NBEHUXZq7Q/vTPVLwYpLcpUYykAo
6vLQBWpBp2NTPLXan6jtuw==
`protect END_PROTECTED
