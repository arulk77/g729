`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zMbI0Ayw3weV62f4QeJ4TyydFWpIoRocr44XhGRXEPP
wA2j9rztdcn1ummKnczSCX9tAdtMJEErAVRGyls/orqSUeeKpJFj2mTjOW8hRAmg
OycU2+eP6w5i6/wa5krMTHYDJgxpivZeRVuQxr4TXuqP2qTtay6QcLzJqEncxJMp
EOT1RqfnaYMYfJhzuZtR7CEcJt5GtT1qLoGPx8JjqEyVUYVCHm6bp9vwKiH27eBQ
p9VrtUN8uA10N17Z1/2l8hoT5C7McP6JijnIhF4GdRCdpaKaHay5gLLvcYjqwE9Q
e/Urn6pT8DBg/PiDjfygoA==
`protect END_PROTECTED
