`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMb5zKfNvkGxu/iRoJvMa52qLaY1WVwdeyrGZJlSBvKy
pGAkMNFHFqb6cNLbMp7+HRPLwouv5mBPmOupT1We8SERiaV0FcLq11zkYgZaVd+i
bJD9ZKhdgTUCIYOMUpMNtmKFsnu48HaraB2P6JjhXXcwQt7FOvJsIkPdWE1epmk2
fi6BRCwfj54N+nqihsG7Sw==
`protect END_PROTECTED
