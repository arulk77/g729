`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
l0OYwtmuOqZI83f41X5uz74hmaHAgEGOoJKRTt4TXwwBNIDtERn4cIJcldgvn6gK
pUmnT3NJleINNOLP6InJgygM+yazG15GZOpbAr5rg2acTSRoWS0kmSA8zdjEAeA4
MZItXU33pGfckQPj6E1YcFFE/RJkZusse1DtPdu8wd1Oi5hgW/S/gztrWCCqVZHo
DvNaLQ3epLDsXe1l8EIeY4LhV18rwJr3qAMLBoQk+1AvTOr8r9ODnMdrBNwgI3Bp
3tSPpKy5W71rDltqnbXS3bFeqOZHUVuYv6ihfpjkVPBdDby5MMlhu5C4M9teh9u0
HFgNoM0qd15kZkuX4vbgquFpvuxAkY0tiemYaDLyjus=
`protect END_PROTECTED
