`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SZP95gTw231jVTlAnEVm6f3arf0Zz8DnuqFe9PfUucyn
dK+XOfca0kFtJDpAe6vO2ZS6PLAK1rziejeu3jIKfMMrpizDf4r/mMEMJdK5fcyb
iAL5nQbLDb+B3+7v7nUuwjByxHDRDViytGzpOD85Rvm3iwfkDwnlUGw99A0ohEyt
v00sxUhvSWdAZI+S04M9fg2Hd7UZxNlR6e+4uZOxiUtQp+SG+gHKw55aeSYH/lig
E/PLR3tFywMsycXG8Y6iz/B3/0bgqBSdQ1Igvg7cYiSqJooBlOXfFLIz27Wxai6H
P864MSxNgboFmq08gIjDaNpnnp85DNsG6eoQqau7VEQEQ2tA3iRbvpytRRnATIuB
JQVAUywu8bN+2C6amE+VZI2fe6VWAsxnGjTPC8M9QbVmOdHOdeVkAOIDEMxwpBH/
/iGptP9uKpo/5T058pLxrWRsLRic7ZosRqfWAohC5be79Tvd+lz89qbLLpkJ30ru
Rbpkq9IQbgx1LA/0ub8wCILArHaQz4dEwUHmifeOxYYGHU3+Kyooxnj+bmnxB/G9
4OsjvbZ/Bn1cgoVF0gXcOrF5KvIDVjeI+17Gw95NbvFP7W4ViZ/s0Fe50x1fzqZx
Ra0gErzMrJ9fwoPOiwUdZifZuL1rSNJviDjCf0D3tb4GiDoXekrnFVo+QGhZ2EXJ
rdxj6QfxTBP9IC9EEO9zEw5wj/99gqYM3lD3x+XI8UHryMLHk9kDfWS5Ea4UfW+K
5ps1mCl1vrkkI2r2P3X00PWSNZh3P8PFHpTiXKhTO6rz1fpzRpZK1ZPWwOXO4WCP
z8mwXo3ypEccVapxtxtQ2eDsSyFldw8H6d7IoHBv0jrSmWUhyZPA3IGfL72hOcSl
f909/b9iqqIqjnYOn4Pb15i+Aw/QT0mRsYZL5TOpuK5er6NeZG8bGQhtpyi2v1fc
f97fUWJ9gljv1uwdfGKu6To6yXO1cbB3wo8NFS9yt/xA8MRdZKS4tLhdAzUujWBx
InhrQqS8BibBJJPs491HU9qqzHM8X/qvwIp+h8F40flYAGs5Hm/94L0q3k5XKkCz
vToScdyYdyVt+5QDZxHAu4Yp9gG+Bn+uKbjdddcVUeq5i/2XZ1eyA3vydnKEjwpI
ML18wnjFFQEk7LCXDhSRPcfua2Ew92DGIt5SUV1dLaLsU25l+4FIbXmvmKUYhr74
gAtgqgeOD2RiFktByWJ6SJTiwWYLzpAGD7Ddzf5MyREQZYA23oWVjWhxhbfS94X7
91+qBNJNf8/EWuY1EqZIEAP1pTOUY7dCNwTRSoIww/W43bE1aeMqZPmu6uprsu46
+YKXrJS5Cn7FollBqOyEZGm4ulLrYg9V6Cv4sKuJzj1XgGWh9LBb4HtKrLOzLywV
gJnG1HUBTRBFt9Pn2StFTYqe/CmssG1645kQN83SJB2IPYTCRKSrZg32Y9JzVDPx
UG0KywLD5bvJdMeDp07iSy9PeheAN47BtvZFsRY3KtWFea4pJ3EitnilYfj+d5vO
am41ilMCX0snOe9fP1kbyxLLDvurHBPlyr6Ng0fV6BCSkKWfXAxyTZVBiAXZ6I19
VqLq2FfiUfNWdMSN7mDFgXvYGoXNso3rzcIlW2OlGup92SRErVYe5ZTqCUWIMlBj
ioclFXP2uvDqBLUbwXB7Pw==
`protect END_PROTECTED
