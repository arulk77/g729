`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JOziqT6tO94csM1R/t51EV83Uf0nM0ORjJk6L+8znl/CmcpuHcFoxo9y7kWE+x23
X2kre2XJ8/Vgi8TFC3TwU1HhvabBhi6t8sVSdVp90bXW/xYYPboJmLz/vtiVn7yJ
wSmd0vtG08nYRdBxjTK38bumRbmOz1O0QQ2t0ZReISOfTaoZtusocZEbx7IyW69O
Z8SqDl72z3xyccjjOrhMIv3PwbPfcJZizNpmgoviEV0QKJ7Nwk5uTaYl7wNw06pq
RnW8FRb/1RJfz47/j6Iz2gcfBXXNj4l0DLBztUVh4gAMjZtO1JvCeN4lOqG3fUJ5
WnmG28uiSnYzSUdytO/Z05VPsMBgTd1OtDb8p1D0Ivvtmi44bl+s0jCXYeTfXZIC
mpZ9gQI6fYYjFHFmkzy9KSp6zKgcZRE+B0rwznS2i1fAHSe0ieOOqAPwmly0b7Ef
d3zGl9hSQytdcOZRHU/7nAymrOH6CeGKATHziGZiTPDRFoL25Peuy9ltHV/yR/Eu
xGjLxGTjcWNUdd68MJfSY5wUG4jIk2TW9x7l5fgzIrBN2z7A3odI7y9cAsTtzXRr
M5VkVTWcwLA/pFnNYoyEtQg/RzF0+FoxeDVDuQC+1pLv4A6HdFbTul7kBmbWvWEA
VjDy4c1CxvwHXtQqFJy/3SryLlH7DitI6hlc8vtdUdqvLdn3A2LDWebD3FATIfNE
Of5kcTPgjUcVrup9UmAiFDBbULOxJhOs2/NC23pyKBBemH9MyVjyrEqbA6qDe+sF
T/tjl6enOaaiDmD6sHkb3Yw0BN2txT2HBaDTGaNsb/0Rmut5L6fePO4nmjiHD1jb
zaw6Xy2g1A5aLv+lJ5nrz7IVcow2YG/cLw5pVWC5VBM=
`protect END_PROTECTED
