`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bh91kMm4V6rCItaAm8IytRV7ae0ViOwih7HaX5C9xGE1pnDVVWXe0L7fFn5fQrlM
9n1wZkFYLtUcznvakyksEBzvuWoh60mlt+O3QZo01+OJiWS00eg2r3uI7b9NKbF6
IZSIExHQvDqGkOAwS6aje9bunX2RPDh27DGVz2Gwx6j6PQX+kHaICUpnLwmpqkfq
+pCKo7z/vPsiWCDoPbE4a0ciWHayn69yw8CiFPFRmmHSdy1tNfYcZ8ckmnbprndo
sRMAvebkj/z9E3tOGDFM7zGAfW28SojsgUYkzKiVpo4ByBD5p+EqTfCrJanewnW0
1Z+H9ui4ImWZjantyCQb3sxQWrDfA9DSBfSr2O1V7SE=
`protect END_PROTECTED
