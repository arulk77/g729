`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOgJFIRUsT4X19K8zjOUDKupT/trflyfyvefsJh49IGl
EER3deYL+Paursz/lYAvhmXtNdi6H9QV2DWsxV5dz62+lrmovMVniy/vS+1fKyKM
yOcMCdDTWtUjuWtjJvYo0KV/5bQYNtiuiWVnZeUnoDoI44x/XzoOL26dW3hQQdMv
QuJkc+QphDlEjfOpPuf5r90punaZA5lRIWS/AF+hFxKdc2YTIufQWBjZKsB+7epJ
FekJX6/nrr/Uydg+JhIL3jPNGnYVFrw1NhjiGTB5Dte+eXRhJb4np8p9Z6eqKpR3
vEEZgQmuCjRjtTfFD5NsugkFTBg1U55CawLIiFNU/CJcUNECN99hwVZ4CdAlCwqE
D5sGRlgJ8kkzBeuys3HHJrnPIb9rFrJMHt/2JLEAMKzxTU0jRrf+PZi4ntPP0DPw
BInbyKwkAk0QL+OY4ViQXKWhBdhwUoXUDYDuMHSei6ubmGpcv/osnAEOiz1+9Lxn
XE2Wxqkmgpaoz94mSKOsvCxeeARw4G6OeMZ5iC6w8tsRV/6sMRrvxy7l+0/Oc/TY
`protect END_PROTECTED
