`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49TqDoY6eFrja0I/2fbdz5BV8+Q5X/4nnUI1bK8eqwb+
x8yjBAWMCGUup8NUFfLfL1YLHmaTiRWuY6P7qiOB9O66R79A8bPIvBUjJ3bbi3SW
IM2xXKCs63A97BbJKWaip8giRKSrDjzeCCtX5jsf5/UI3PZTHw03eLu56gQV1wiD
eftU0oKHbs9pSaoJeWzf4p2HxjRSX05UJsgw/q2iiC08A8Q30T0R0xgQ4UHEPpMc
olR+mZDjtlomZOBMZ98y65M9a18pbsZf14cI9yA2lr5xhVyBsHE3AJvhg9KMKAez
UhBckNZuqAqeWgDkK0jcCg==
`protect END_PROTECTED
