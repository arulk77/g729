`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBOn1/UTF+hAWBXNb2pWjHjaJEa/kAlSVJVgeUavtwIC
yHfkmFzSpphIgpumZEWCkgIkDXOuDUmqT5qQVJxngEArjap0kyF1hxLuriew1vms
inm755bHofIA+d55VgrZedKYAlOZQAveMMOgnLFKl6lJ1Wkw4wjFKK/HDbZx/M/h
wuxzlNZMtGc5P6Xyoi91L3iaXdO7tZ92FedKwHdEqoCgOe7oB9iDrOwAousgQt4r
f5qKFC55cs/zqchHq2Jf9Btz1I1nVC7tEQP3Js07PBn4ToFsHw4nYz0puIhdT7WE
aff1S2CwWVhtOR+9YpJWqgjOknga5n3Uf07MDGA3KlJqRZtcm+5TNTyJhPS2Bq4e
adWZ0Y+EO9HTlYHDfd+65Q==
`protect END_PROTECTED
