`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C2tjwm8Ox6p1Hyf3x4kOxiVTlw/AJyaQkTGdBimX44wX
h5ojrcaT8hqZK7dZ25Rq8A5ME+Ok+LAxZMYB1VezP9aKsIMVfhvabkMSc/087REe
JDFJ9iREI8bbbIiG+ETsxGJ2ZBLa9gzLgcbY4bmKbOgjX2aoo4AMCG/YAPsTbYDe
DdCvWsgvkm5WL6Bmtx/RMuKiqdERgt5ywvTFBysXbNEE9nzceIV0mTChuQ1v8kpn
Jr7buw8bK2NyHpiivIPQ3WStbrIgxvVeINmD9MBmnWc8jEsfTiVpHhbhXnlNHmRF
izr+T9QZqu2/E/cHeNHC9sVQ3fToWgeFA1ey8TvPNrTt5f4n//LUe1aPQAwZHTex
+VydiHWTsaxSzC96IGH69vl6tZyfUPtTSaZgx7hOQaLDaodMwGAzUEhpGLh7W3Gs
LOgBPDfdB990gbMLBGgPafuqG6c55SSfKQU9zfacTHlBJ6D55x7bOg7eyKq490Ej
al4A/8aE0Df2VtWbdQiWoZtC+O1pXQbQGdYYexcI78a2D2PspdljgFGMfWNh8tqM
h27QQjiJEhH8Ap6eU0vIB4APQL/c0pKbsQDvn8lvZWFW/sPDf+zwV2/4lmXgB/9v
Om6TESH3zf5JwqPReWThTSYdA1kTizoRVNNvzNvg4pGcmTo+REGMRQZTzWxNhGs8
ry0TkpbXbdF84m8UOm6yXYX3qZTjuBCfTCdWm3K5RuPHqpifpJnFHx3zCuGGXjXt
xf9X3E4FCTOiO9IqZmDlNVmYI9L2FU4GBEFXK9ONHeu7HhFW4omwS/TiBHX74M0F
ufcUxQds55ckLr7+ac1RFBpbDE++EfJlBaCeg1KupmJW9SEP3beTI27rJ/Si9Ut8
BVsYeyQRfSihxmMG6Vp0z57MeoXfwRPEFE825snySvx4rRP0IGdJVO4ElBCMNAf6
erC5jo9v8UDcx3lPMJc1lthlny1YrFgriDjmv6R6632Nem2gfa+TJM0SSbDdu9e7
8FR6SD30ru/9TxNvW81VHLXm0icLCp1dEZ3wVADBAcjnb5p5mH3pTR7qHgW9KjmE
RZVgQp0kAc98jJOG3TtcoMtljYzZ+DqPPTWAAAazB+lnWToNv4ziAaQnEk9EJ86P
6WLXoh7lUEfTxFJKRVndynpc6qQF1/cpAbkPjyZyJc7VcHcuTlXuoBaNR0pJSbDv
jjitpBXVafBZchKau5+f/tAHdWiAjpQ/CrdRKX660wUPb4cql5Ppi3O4zlezpUEE
mj0wSyvgZs+lil67X1FDMXg5zwzOGfmLsfnqHl32SvZwtb1rxl4LsSG4UZCWTaG1
Q3YlGbQaa+DfpcItnQe0S6s56iDjtAk/e28lWo+7h7/8YwKRGnhb13msgky26y9A
uPaKWqxM5odZWiYPYVhPyYik1A3ODXpl+CBLBbSYT331VvqizIPZTU4QcBwYfIK8
MpEMuWA2wg49n9v+iNLG3HIObZiVRdOWEjGj/9skEDYgp/QuImLAdFgh264Qk7z4
G6K5RTpc9t6h/JfVArud9DCP/yA/N64dbs01Koe3CqBXDXTqbIbP4uD+gyb8iVGo
aHsGGF0ULbPOCUQS/kkjoNL1Ves/1AIrh2wMtXqG1mUbGkp8VkG+k6OSzo2B6H2A
LKwmbQPmwpPw8e38RPsTxz0NsF3b0ly1GT9xRzcXeTsbpgHrwunauN0N98sQM+cR
gTYMbck/U8hCZWghCzuhvei9O6NDwMhGLWkEDcLBgrEIb3Cz0o5ilph/kjLrf6WT
ppZqQ4NUI9nybv6uMDWCo6hH2AJzw8Icv3ixfJvk2qBJEan/C0OIZWeCUHIJ6dpG
YfyJuBsVg0MWfQ43l2p4kwt0hCZI4jWhsEACo5GryWH4jmBcnxCBTsgLVRNJtas/
rUFj0dL4W7zKsFoZh6cHGUjxAM7qmg/oMJe/Jrl3Xk3j7R7ScoNYjtKxfZ/YorKH
DN/Up1BjSVBs+ZEIYsLuHxrU7R+GFWDKg0UeoX++0XNjJPXv1+vaTJdnO04iES+4
niL+IQV31LmC7NJugs646CUygB06yZb8GylCeG+l4uqmt+XzFD7Askne+wVX0Mu+
cJ7Eb9+6Hpn9jY3wacpuyqGIi8To1LEAHPtcur6HBeYWlbVWYaUHdYwoaZjKAGRA
qZOpp32gio4Q4+UyiLshSVJKN2kQqsuGqxD2IfC51X5zSJgtC89xNoiFwsEpu1VT
9I7CjPumyIgrv+iKghIDL9jsmr1UclKr+uyC5JuGYr0995tQHVSj8H3/netZnlf7
O/hYW82IwNzbY/wDYCmGWUQ4qjp4D6HrBpo6f+KKXUVVw30z2gkGWCMzC+vm4gp0
ef0uwo8ICWpb3k/ZM4gQCjmJbnGEIRUd0Vus7wYOARYqHXXkU1F7RuyKdaHKbrAH
0rZ/KF7jTtLUFbDiI4zDxV2p1tzwrRpfYS0WYjm2bTmGmn2Ls/bkP4Hrzmo8D2KX
FuQ/Vnits12FdAokXWil+W74R3lb/9saO01gBdoYZ1sdY3lPJpErK7HDYmK94/oT
HFdglzAARhIimSZFYT6bVlwlvZPLyqUjPDpSqEMSuuhuH8vUpXk52GWomxpzPOWP
X/O45Uk8z+tvaVvKCp8621TZCaC7tPuWrroQZQFeY7ULpDMGG3g6xKT0wS4IoqLs
ew4uH+LcuXe3R55dfkguKePNsEkDG+8mFa1XZTk+R1cteSpVuSY3nXx+rK6zBW6b
14BLKTP5hHU1cU8fro/f4cajoiswyO+MIOzJYdLEctqWkiq95RjQwSUgJkOLpvFN
gxoKwPyRT7nwDjg98/gLwdxTTxTxVePinl3YaV0JG1YqTnF0BtpjSstaTU61sgYW
CMlEeThopqE+FxXJ9axrW1dUm0+Dynu78mnQTZfHHfyp9G9BqZ8wYBL1OTi+oLMN
Fab6OO5zdhtMT+Kwl15mu7QzNC6YjQO+alEyQOue2Tv8QZJJIUcMS8L4sACwUr9f
3i19dpAHmIYFj61jKsVhoYSRnujCn6H4WwrQpCBg6hw/B89bjdARjdu8Hrckeqx4
kP3p58S7eOU/CyLtTUrvfsbPIddnnSbA5tOBS6B/MYE3wPVywIR3NmCCGwrDUXiB
XJA1yJ+nJa/ktcPwYeybcSH1chicIf0HetDJm0xGiYbbbzOaBNegW7go+Jzeq8fl
Qrccy2WqDPtw7OrL4SAQffxgNsAtgGIIuiax4nxP8e1NX37KBWVSo4ImzWxFapGz
jnxMuZhkCZuT4yn63RcD0Gj62Q7hLTCCf/wC1Lv6fnPqFmi7Q4yQ6/K07OlnXrGp
X0rbhNt7GaI+wvBt7NhWGtoXG4QYvRqZkLVOjEJCmI6PuUhoSqqaxTbmgpqmybbw
gsoZLMPGwBRo8nDBD2eOewYSsaduqbk4hVp9CuedJSH98xlcBPs9LR5mZRw0K8XI
1rcdFU07bqKsjJPVqV3VInZah8JyyobjK40VdLtLvgX8lrVjzrT0Jlc7hAbazEv2
6icpoyNYxH1crujC2TMZYJFP9UjJNvsYxCXZoeQWPjB1rVWfNG95QYC0iyyyUujE
MMr2oqbBAlgO6qptkg/Foe+LxcnFr1J8npQcZlhjE4dckuA3AC2PtU2wOaAMMCvH
pn1jt/oOY7lUgZjmbWQ9dlfHIezp1YdYR0vrKlLWyBck6fRAjLI0LIiThsxbxA1e
ZFxoO3qZpWGiPQV+bcvhKXVZPgHold+DlIaOaGgGJM4yuUGLg0/GlcMQ2MUE2Zku
O2Hn50qctjaQ2GmLxmTtq73xJHzddby4Lr5xXyl0vUXt7UJC3dHPvi8IM2cIr7Fy
ViVb1OesEjYE9+lzducI/9aYmH3ZCQ83CFuWWWxK77jBZ93at44SGFayKbVuHfFN
vt+QVOTXW7vIdBajeA0Mex6FHWPYWvbBDWXY2/+kloi6rX61ke3vOHX8D1O8PWMH
JMuBmO88evL5e694noepX/8oAbZgBANm+FTd/JBVuKjOUJaCbTqb4tbeUf4OoKaG
6OTB7tTzKirB17n8QobgJYiz/FsJV/TYMzaF8ew/VnXfsVYIJdQ2tuBBQtG/Yyp9
BFBl/Qg0dKnZXE4IEskVkNo/bLyG8zJvtzbFtvj00IHCqqjAwLdx5y+OrrE1iBi0
ZKZsDXu7pkqb+cYtZ6HMieYNqLFfD5FSFGLVX2cKyuNg0RlPZV6A703XaIN+qqYO
1BMIox18FRM41q5YMj1A99PHtQ4EopYPpR3cIFAQrPyfVmZoDQfqycpCib7TmMzC
pbTJWpc688Skn7ZnJzOXxV3tg4h0W/RDpnDHJE9b70jr9aAsvxFQ41Ltwa2JM3vJ
+TNjujyTZ3tfhezFUrH5GgugZBSX1OAdwxefBPdUtaBsztSTSq3hNWOg7jtPatul
1uXcW7M77vMXNfqMcN72adQUGzOktWZQht/MW3RyqTiUjHHU1E1fFfr+Pelclg6n
fnCwTfGy1d23rtWqGweEeCbbTf9P06B/6TG0e7t9wjs1g/D3V0oR05LcesfAdRcy
RKqZU81RUQ8ZoUOL2o/+jZ4ZhvBIvHeLFhqXXeaHfekaDJQWm4paa5JlJpH5HK8M
uV3dghGzF10IsNtPS13H7hc8cEftgQLNVOxsgpRuxw6s95UJ7/yy3d6MOkC/otqF
2F/B0ixhfkOUSbYo60LjDUr3qufE0vmZZJS2DJAW+xYHyYrNlklH1jJTF3r4UWNo
QAdAO9NmUhsClrxjofQ5CP+TBrZpmepN3lWi97QvGJrx0TEIUuABRMiLWcWxePO8
JkeY02F+pWmXxto3au8ZlP4IP1qu6rjO1TyrJn7Ut4eelo9eAX5+/Vy2+wUB2V7M
9YCKTjHUdXiUcmJwC8X++7uI66MAupNatStOn51NkNTn9bepKsw0KBYwRS99pR2l
cvX3qavRqAi54ml44I3D+9ZJaDMvNedzaZObnPzD3fNWW5JOyQQ2Cf4aNzbGET+1
L2nVAmtu7V8Cgj9mHXX8eKLXNJ6bFx9CPCIm8QFJTiqBN8Rf6y0VvLHQb5oxfIvp
OMMUSk0YEWOUUjZ5MHCOgoeD5u1lH+CNPI9bGqcrlNAZ1sR1PG/9nV6hvPI0PERP
PGkQ6QRvFAWbIIjqax2jig5aM3VV23RlbDHa1ufLvkpC9k0nmyVQUSqYxeH202Sv
XwuLTUy32nAtK5xdAwkZ4AArQQ4A2SyEy4odpCOTbXM6kl3WuASDQ4RsBYOeid+l
KedTX6TMlWh39gUuuPdoDPDkJy4/TVIlVh8OzsvvvDPCNfr9SpIAvbGl+86pR3yC
qYvWFc5VXMsBfkn0qggZMBm6/CDmRRfLVDQpYgegayFAxZqFIn9ih/lihV5mmdy6
CKbg0IhqzXLleULuBi+BJOvZcDdu+sdpnJdJRPNGzo1vnshyRZeGJAFpVkeNA8Kj
LX0Ys2OF5IjJggjZ705rJnHktDFipcxEpKXhi4aj/yFKc12vlIFkKghgeQ0YKl+l
1TaxX3loY+Jvi2Pk8kUGNUzKV+vK3TbuWEtWWMZyEZ52xSBo83ryMk+VHlVlsHGR
Ms/PblfFZcfs8XoRiEpTtCb3tJhb79rXuoIF+npaweipcPew9yNJ1SmRsZvQ04IV
J7lCDI9zr+Y22FUd1k6iVHfuBNZ/gzfoagxLYnEQIi8Ci+rzBD3mFTJahxX+5ws1
r1L6pOf4mGWrPd66OFjpkA==
`protect END_PROTECTED
