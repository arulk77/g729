`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
/QR5nO0+OpBTrEaBENH3A2iplK0428NUmLn1noiFCw9UaUDNOYB6CwLYRpgcJ2am
PwAtAEPBcnE9Mec1q7KKBtud5DnmLC+eNsuZ1/G4ggi61OLuURmjoGaQ6GNoGHj9
x4UlB8ETXK42osv7RVeCXK7v+s6iodlD+gdmw6mnj6/vicFI8cTdllA1DgGIfbRJ
luNKfEqxTJ1Wb76oEp44xhDQAuHn9yV18GEj4Cq3x/0AaKDClsLNzhMxJ/yVZRBa
xuvglGD340auU/+wpu9kAe5N9+ZOwbe2VQ6iQ8GR7Zo=
`protect END_PROTECTED
