`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkYG1WXT7OvUWBfLS2xcsjo0UNNqJlw1A0jM6M7DfgXaI
q/VkcI3XAcWQioqrg4Bvrtz3TUqQAxVycwJp4Yv8zSp8wTof/IIaPhQYroDRSr1D
26/8/+RNaSWaxVMqM2Ti+d0uHg7q6bFqbj/vc4kXmE/K5Z5BWhXLQT3tFqMTCI1I
bYwiUcSHWEyYd9ZP6CneoLhullccfykbP0AieAI12lWwJP05G3hUJnpWCZXHq/xv
fAvF9DOjsjEoHK8q55g9046ebkWCnH9PXYojiFvfp5ce9IP1aqyC9SygbXZa/nHF
qQ/03a9hRGbV6EHD1bclv6K1uxZvuQWEhRplEiZKYy///LvrdcU3TvuRNHVqhNLq
eEzah1cxcNguPZWT2IzEh+ITHN/c2NRiQffco9CIQxiKnganOb9eDtf2oLnuG6zW
w3KicdBYJlK+w7U7TtrAPIy4h3yN+lr2kA+yLrDOMFR2O8SLYl0qTCme3fGtQnTc
DNCoxmZ2Gi/EkCMXwygL/dgZjyCphbbk5Ija86P3ntJc21sJAANl8a6L54TpySCq
2FJ6v8wWn57/vO9oAWQt1wtbiq7p9XhiyXRDIs8oF6aCDZ79MCYAs6B+e4v3Bff8
y5uWrlmSHVHnWYhfREPuXhxBQLWAQvtvbWc9voImJsPwYwGFj8VScUFdQYHd1d+D
POY/pD9A7osXyH65R20zN4NMhT5OwGpoy3ThiOjs501rTZ+O++LYfQ5daZpNCCp6
HKBi/g6jzbHbkWkpiIdEKAF1JYT89EUck/HQX495L57Nr76cPeQVH9PqCGRI9NEo
fuBSSUI9nezuSud2ypXLYrcHPDHrLgsjclS1Q7xN1f3X7DURBZhD/JCwjgyxoXJK
fq/OwG+qR2KQE71l4i+6ZvPVKshegAR7gdQzNJjGBgBB8UQwHzVREbPM18aplPfh
9fP0MVhLAVENSB+Noo8V9x4i8qc07/qmJ+8vtiO77XJT/51DLuGu42OHVoc/XZMl
YB9xFeuTbKaTOSZO0579UBCQeC/hxroXWrQqrTSxp9cnnPg0cXmjqhK+/S535pLZ
mxI7tg5neciOg0MtPYApEUvl+5or+U+NZf/FExdG3SxwExSF7q/7oN6BHC8apO4e
LfsvoDC8xHphtRcu5quyOjKlDZhNAlvosiQHywcphFGiqfCFVQt2NOKCuntNmZfq
pYsuRv9t0ILFyszS8cZu1pWupMgf5EuyZRv/aH6BEmW5cuc7uoWKk++iRH+AoScz
eO7/oP9raRymH1WhL1l9tdjTI0Vdz78iBRdd0xPdQaf20s9h5yVbVEXHTP90ESzK
mbWVsdxE22AZzfFBvnUt3+6+rjK6HlVm8gddczuKyankhSW2bkU8Lzd9pIeq2Z+4
ap2/MpwqVDfg2z+AtlgYlnE+eH4h09BzeRZlF32aCN332GMU/PHskZuIs8vPVZMb
T+GBRa6OTBX1NVxI8oQPVm5kkJRfxSQunJ4z3DDhBrb8OqBDZpVKL4gFQWAfC5Mv
kV/I+pJkW8RRhT96FaNPQdqAZy5OXStOMPTPnu5FyBE3nM4Yf4ZinTIR9J0Lqtc6
d+hU6oKKKz7CL70ygv7OXg==
`protect END_PROTECTED
