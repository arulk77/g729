`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40iuT5Zo30QMoSf9ikdxZFOhpV8ihocfwmh3mw023U5A
vs19tApYIpZR6E6P6Nzq/1XEUapyh0jBcqE4QpmvtkZpDOdxj+Pn8Y9OWN4gB6TP
a2D6oaga/ENmi1U89WXpRjCdxQailq5/AkURM1D7+9cTc1G/Id9873vqTD2bHZ3W
JMkxuRra/iWGBivA9/N8JUbcFy3ZFowOP6fAexR7lxI=
`protect END_PROTECTED
