`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44WH0TqpSOEAqDJI9XGG9KyhrjeliVU2OP9QEhUSAX4B
b7tH5VS/aTeWpzHKSU4G74WFqNRuxlCDafxF1s12SfK6uH0cCWKhSVDAdh373XrR
hksw6zlnKklRj9Ds37dT27JKQlvZ5olco0WLpe+DU0PAqIcefUBf1CX2pF/TkcIy
637FalJUfGXzpQxXTyemXGFGqKyDgVmuowQ34pJr97wMCMqI1wldKZRYkuJGzQ5L
1frFkIq6R7/2KVNCwVH5TgwxeMcavR74Otk/pyjs9NeQILEpIiPFBqu+7G7cx0xU
iSwyE9TtBzlguArlZZ3xxU+CzZ3m7R3p8AxQ/kwwUq8hOkGxQL+ya/UfVoc6GHOE
izMfDBf3lCTLZltZ7kh+2Q==
`protect END_PROTECTED
