`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDxGpxm5rEuzPt+p8lYbTJXD43/DcDmKt/cCiJFEX99+
uiKxqCuHIzd9QeudOD/odIi7JWSPnGemkNzcwi1yg4oxe5xFD7SgVf8mqSB1K9YP
ir0ZoH0RXpOoPvzBkIj2daCZdLltPiWM74zsM71XMIKOgUQzhBU7Q3DAXExaYVXv
SiBUyFaxSTq8NgxZSE/7oQ+wfprFPAJ3Fif6GuiJg0E7cyPQ0BH8A4zul0Jtl6zQ
`protect END_PROTECTED
