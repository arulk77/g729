`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu498VreDeGV74UmgbUKF3khRve8bq+Gyq6LWFQPU2rmYh
hzxotJ7+GMqnib+MJpEBKD4fHxIQDjkh2KUkLaMqwk6jqasM316LwFtJtOy/Z6x8
yKkiORabykDCLisAaN/DXW11U3mpTRRCEia8qIHjZ16bIxZX6WLwzS4ZW+TRB6fb
tRbXlTbyqZwdkrnV41b18a1Y265WJd1hnGtEyDXVbVE0QZHGoYy7PY57VKEJVPMG
dLx8KAmtt3ZOl+isPfEboXLKqOOFGyyyhnljJFNvCq+bPifN7eLn5VugmmVeCaHy
u/mKqhZ//v+KQTV5FifJHQ==
`protect END_PROTECTED
