`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL8yrrsPPDhGGVQH5g93gi95SgXwRmjrbJlJzUSLWWHy0t
Ww4t7CpVdkEyxLj4AXTX/xuPlupfjmbZq0ixUQ9nqsdFSB20FwwQnXOHfjQOm3Rx
utbHYo7zzui76xN7TXqvRZMlniwW/uOj2sH82jROwM1SGeFB/Tag+THuJtk5sCqO
NMVZqE9Zryhn82gHz/U3M0wMVKuC/6bQqegv/fugM0lEmPDqoINGzmRlHOepCOOv
/BCik00UIepNrmkxtFuXbeXog2MiE4cev9bgo/+qfIqsEJ4aPT/RjO6k8Ir9CBKH
9pRawnyUbvVSFu4HFHJAr3j5rsErcwDt7sFIBKtFXFTSVs2NsaKCn+h6UNiAbmKn
JOZcA6coe5WJDgJ73mEBQ8AEN2z3Oeu5G9Lu+A8hKbuP5p1yijTJ2oNtF+hO4j3x
0bEYC3DJMXFOoyZE9BO1NQcCgE8OfnsUZdUkYke14pugARlZxkaNdegEV0uCG6H1
`protect END_PROTECTED
