`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
9UCKqHRMhYxdTsj2rSGozztJNLVQkXulv02S8qI0lY+6k/Uzfvtg0dW1FDY8slEO
g5tCyaKZe5jy2haU9uM7bCyoHx0v41sREA2IsQacJPAMHrfDB4s7qjs/R9+QUReQ
qOrx91ZctCrj7Mb08xsMTXQk1QBgqf0vbqfZWXSHAyi0Qt52F259ohpx0YIbEOMb
DHJHs+WzUHZVvkIFJzrbK57lLeyCoMNTD3tsvg+TznHOyeyrK5wlQuWxj5vlERXb
ounNMKdUNT6o4t2uk+fAte+dzvh7e074rucpcF2JepeTNqLEbuRqwNwbv61Ijyx9
qcajm8nOM2ZwdU8WaiN7e+2gewTz3BShJSInpyeH57QStVeubaYbxA7NeUrEUNIV
ehKRkYiX+8r+1SX2X3/1GA==
`protect END_PROTECTED
