`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Zn6daRSNzeenlx6kPPy8dH7jfi0pN6DsXw89NSBTJ5ESWYZcDo5nSSf/l4bq9kTm
X3lOFHnqbhStDEbfMz9Pk/ycovxVdJpBzMBJ/8xWZtCL+F6pAiBRSmvQ746LX71Y
mg7W/zEwWjpyyQ4Hoy6D9WwpGlvVDmI8/7pr3VlOCf9DvnyOoN90IyTUQ1+9SR8B
oMiIGnY3yL4ZmJeCyyPeAtOnVyCf/o6T+05QFWtXe9SVd0u2/dHWJ8x0A739175J
YWs/WqvTcaEkgU8LoSnht9EisMrh2ABkR1xKU77u8JkHoyXwh2MtT5aJgD8llsR6
aF5RpPEd7VdVHol26xw9u1OT6ketY8zoZMc44zQ0Mrk=
`protect END_PROTECTED
