`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN+JN+kb4X236aojy5Zw+Yqqgy0CU/VO7RB9vXTx4LdkH
VqppWbT+/hd+irRZkaHowTZWfv+Y04lI2YVbzzFenSfhX+LcW/lc4MU+/1QoRYzq
VyRDlw3kGrjjO55XOOujLVxPkIX+Z1DXbKZ8VCMOhKf6bB8lrnNZ7x3SPM5h4Nms
4fKe5HcRBFSyLBZ0n6iBsXcNLgrSP7zUCQ8ZtVP6OEWX5LsyKxhyBIZhx5oe+zvQ
qoBSmVORImF5fLY8C/+Uis4uEdB3fSauUdGvJvtCBLVeyC/fpM2reRjriRCQRh8o
AfjU9abB/K4EHYm768VsVZiFD7CpzTvYtAY/cEy8iC2340aPwdhn71wMYPTdh5Ks
gREbwnLmc7bX3QGxKktZ/vyhtMJZxx/+C1ATwRCIpLSVQX6K2/o7mTabsLbh9M7Z
UfR3Sv+7HtBbvAN4s0Or2il5QTVOMgaNOFetx7TMpPkQIwKEdYDRE3yVGfZlRIXH
+j2wOcv/QSLNOuBLwtUgm5YD0IY8R+DlPtoES7PGxHZq2EGgEmML4zABp8d3YXSw
XtfUdeQM9x+Uel2wKzD9kUsTEEntniR8nFk7XniG9yK5DhzQnxPXEeE4wtJFBtNV
iGBeyQwX0ELc90T5fRiBJuHmiqSS4tR2XcJ5ihXKYBch6mQWhxum9r4CMdotCXf9
rmqJ6pNNiWXiH4NDrRv6YTW6DO+FEzpwvFTvg6vzEMHMm39OTQj2e02Cg832z78w
s8FuOfO+nB8gS3tmvkTwGsiKO1C1WW+h0SR30DnJ6Q+z6U/5YN7Gq0M1506C3f+e
RYxbHMl+wONeJBzXef2DdKI4dGNWIRmGANCDsxeXKXypp0thGEvTa6BolvxmxL1p
y7tdaF3gzSHqNg8vs3PfkhgplaI79919ZkXcru+fH6fhKFBoJW5uFyhdthzXge8M
Qa/VF9NbXbgQkfnj+fzs2u48VPR7cqTAijZLSVq64x55t0O3lffSN6YepKsxhDGM
lk5ocvLCxSnL6kdLX5bxiqAL0QdvEIn3+boA0gDwXcJv1wbHBBanypZw8tR+cXb1
gd4dGQhMtVtgfGfk/ESOhlLvLVyZxAxO8GxuAHpxeootggrnlV2jbsJFDnVGsXnQ
fAz+zLZSkQ+sqyzgfoIDW/kZYYCY/WI46HL7C498xDW068zMIG703dN3JOQEgTM7
XEyhE5UYGQnxcT00a6m0g0rJlWCQ9KzUDSRsmOy3M+xvcuWNtn4Pfqel6pl1UFlL
KIT95NKBNHqfQF5PifZF0wDPnM1uxN7sJaOOK/H5PG1uZgl4vX/UCE0lVfcxfQ1h
R81nIlTqF3zRQkGtdYH3hpLR5k6iHr6qdGPA9dtcX11+ju/WxDbTWfepm7AiGMyw
oDb01cHl1nK2k1aec8e1VtwOSwxpxd9hgH4ASPDdSLptCzqGkEWulMtfNXxizKXn
1wzY8yNrFvCB5apsrNHrTeyk3esVBEU/Yr4AbUGRA4j0xKYco6T40V2SwA/nI90A
Yio2aft3zidf0lfFS2TaEk23o79T09Mm2giz2wPAcbhEibDtI8j3arO56NBvdGLv
VHj/7pbsRRQ2NBcvRDWH2kFFiffoo+PAjeAyQxr5ovHQjMmFkThjHhLZkmn881ZO
dCFJMcVlhfpGzMOkJ5sWLV45NhWhZbtp4K0RnzsiQmlW97X9irHWmYwFcBn3tV0h
RfwycIJaSm3W22y1YU08kWOqQRCUk5R+kkXXOyO4aMAwCDzB+NIoIOrKtFw2A2hl
XiWlnkmPoKs7y1IjvvgMbPBYg10ijRO+AX9Wr+nRYXM2JCqjn3R08dHCdGgeoDyC
goMEr4yVSb/Z5EJ9uWTAXEls8iWytt4dAxmx6zZRJ2z3hSbes2Eb6EbaaBgETMO8
6ezjIgEZim2LTO/QRBTpGjG2VD82FWuOAhzCTzpHdAJFDhX0YQ2Wrl3c/1wTp1qQ
w3owfK9LNnAVJB7UIP4wfmTAUgoKSDVN1T9yGtwxJwut6oXlUldRcWmbvbxEXWOe
o6s0S+HW1MuzIeU7yOO1AklM5SpTrQYEai2SoCBYPOJNiFjZeWAatl9dT1Izxsij
cm3mAhmIIruKwRzPaVYuWxXyOgnwl2FSPjTs2edX0iXY7r490YqHzKyI+l6XRayp
n1xR+/Bim0iqZE6IhC+kDg==
`protect END_PROTECTED
