`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wqkstJzaBDVGtvNKgnRSsdVT9l6KuIceIX1EHIIKrii
svlEL5J1/JRegHpQ0shhBhU4lUKF+RemuVAvm/INdCmKnYtBXxt+T3KcmkrWAQrl
CSjbMeuHT4OHCyxtnSe5cHMqz2/d71t4uxCnE/jXf403PnaeHd1rr83u5/9pjEFc
waaE2McQCCdgbGIRu7huTsVPpymQHTXTUt0HXrc7RcwlP8rfKdTstvsDaqkrB+dO
AcD1Cx8UZRk53e5qkY+yMC/kK+F8ynkgF22cgkVmQd8=
`protect END_PROTECTED
