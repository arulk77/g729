`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49fa7AE1FzYpr/9vss9F3R4oKY2s9TzT1/x/t2IhpQjp
NxYW5KznnWEj40agRtUVFAhUna+fuljYwVydrjrHWOVB90JOxFNZICkAPQmr95Kt
42TMMDwti4WdYoNHFXyjmcIdfS989gR06IuppXOl4hm01C6npTRdxjFEZaAannP7
icqxyn7Yz2DAFLHfG0zfmsIFrOHIBCzyY2qbqI9H1HPtSO2UyqSF/l1blM7/+zPu
O3WlOaCyutonH3uWwSUNCJ15all/NrMVXXBc6J15WsmQrIPox7MDFwP7BVJ94oSx
+AtcgiUyT1+a7eWtadaIsmRh6ZImoa1jIOhzgRCxOTcreWcl87qOq8hxN5720iKI
HO+9ezUQRrOsXpJV8zVvGtE805VsxiUxwYGk3EzAsSyYIrOoDaW5l5YnAcYzK7Fb
Oz7hr3EFGDKMUSHtXb3douiRlwvBmWbkC80bptRU6PlSF/+daEsdTNhUgmlBlh1E
`protect END_PROTECTED
