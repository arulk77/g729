`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJRk8FCFA6mOUDxxLb2itIGHyVWoyRSX2Wjq/vvUUirC
QHOrOv95OQO124sTz2S6sfY+iF1cxHyJdBvn15jcJEqrJAbzUv4YvcIXsv1Yq5jx
/u81PQHiRd5uWdUIYl2JCciBotqNYW5V+fJEasjmu8FatcvtCRnnslYltGgMltJK
khbpG2gVScpHm7NqYu285A==
`protect END_PROTECTED
