`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDHmxdFICtT5znqHi0MreK361AdKJEZLMFKkQ4hdrnlL
h5IfLZ3ZTkCZbGjFobsC1AeMc0LmPzH5Vc+OddcQAYbdIfzv+KU4Jl+a2cMLqytt
9ScCMvH4YuM1BxV0rP2OdIEHAl/2AJ1YxbWMTL8DcxqQZEwN6U/Wk1knbLeXGzS+
4qVmXeszzv3xZENuGOhNgA==
`protect END_PROTECTED
