`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDARaF1uaKQRtBjC4nFzrKGi235m84D99ayH162QIdd/pa
RQBLwP4rQ713S4Ht3PXPkKQ52afJki/f7f50IfrfR8cELfhEkblDQbuzYliAh37p
EHxHIGY1hUcDzD8wpypZZfM9UxcIqqkF7cIGlv6BHsaYVWQOG43sdDI+i65OpUxl
JFqKyALhvfG83xfKXcWla4dzd2z8wJbpGOMVGpGcWd3RYXkxYqH8jKvHy0mROiVj
eQCXqZYR7RSbnJK8FrL+Xj0CVs3S/AWl852xWF3oqjP2m76QYYype+bi3/aa4Idy
SIjYxreRgtqEXRP0PXibYr5UN9DXaEhXFbgC7vKr0+9QnrJTzpvHKWOywiACeXtH
Y9ZfXl498L+pYtrTKPTriMyRJclnFeiPU3AIOTGURwukGYASnvHLeXKUeAAmNVpt
F+Ozc1v4lWOFmGAVKCY7gxuODgPgoDkaAJb+H5v2MkVd4fy92H6qPx8aiJLozMAm
TVdYOHvOh7Gocukef6baE/xd6hp2RKseBhtJbz3Ke6Q2zSNGtDXhyG1UtitzE2F8
WOIXpW4H8cqVZcui7yo31YiAehfr6bVotgZZrLmwAowYHSe+ZtposIYN6iRieyDY
qrPA8hAqN13Py/Jcanv4f7lhl1mV9NN0eDlNUT8/T6rys5pj0No6lb0OCmGsYePf
6m93f3fTVbs1BBFM7zgq13sZYUQxEv2rPZOkjLjrPsgaHC7qeQgITjV9tQ8MY8j2
LExn/JcFJYC31GbSm75YtHaORoEreRL+DPCJn1r3AbnSKeuN2VdlJ+BgEauu0f4A
dtdVMmqzFfX0qqcWfjq6HsIAda1uUTjNI6YZ+xH4+5gViGyFjFbeHCuf/YjEhuws
OJmpK5fv5liu1TNKeU1aPDrNb9RGJGYvZUJKL8zeSitBbNWLOcqzPRsmmc5ix/kr
TvXM974jW51dJvDv5uJv1GW3pge/Sne+eSTkyWqwVLKIVkUES8H9GxXTzZuv5UwE
4EAf1oyQ35segTfw0oVoVS7AF+ffSo0sr37FfOmzecpGZJUdS7WUryASgvPMwuVH
YUqLOSdUPP3gZCtowzlvNpZr9+wSpHkGGn5/TIDT0ylVJHzS5tzetN4TqE01GtA2
MJyQAYvFULFSX1JumrRs5DL1bhK6p+kmuRjGpP/2Kh17+yVFiW3Ku/2+G8VZLvN5
BRF5VKFLm0nb67dpZ9suGkIlk5UYu1s4xagDjse1CW+4+pEmPLWAgYUQ4z+ENfXU
46FWlAHsyp4ijZWevZp5SFSzfCBfcL6rF8V9O/FhV3X3ObiaUXCOWHyiqjsjTXOY
ulWwSYBGEPPl/SKKaGdRky3g0EhPhBLgJMbRSW4KjpY6CegGjIWP5s3jmQFdudat
krU7sVQX+rIsv7H4LS4jFg1lblxLvf1o3vM7dKj4+/ALmQ4YrIaZ8yPKELzh8MRY
G1PIGTZaU/RJO7tVGOoGyWFkfCVMhOCGbL4u1yr661tl6kO7Abx0rxzYpFU1vz9E
r1LRlmG+UE340+/YcRDldvpE9tMXmZPzw0XSZslar/Klk/1FtqVn1e4rbQkZMsBy
+Bu+WaaZeizFCRBib5TCd/uT0quOpM5RxaPCZ/EvpubDfu9MFKFtrtvN0BdyhDt+
mSpwc6la0EIFFU59dQvKDTjNBsmCWuoiXE7a4399Pbbm7fj0hrn+/xIU/Niof5eP
TFcesvGdTr4bAg90LqISisLzMNFcezK6rdplXPmWcOXuUA07f0lDSBLjaqrv1S1t
u7rweVCnKEmOSgwhlvyEJxUWCeT75YIpyPh5vWRp9MYIQA0BWMG0cJM87k/u2hu1
nsG8IJdEjJknxb/8+tp/VEezsApyBjcGVejUmMdaj7XmttafVojA0b13ly43uIpq
tBb1t0BN5CYT02678AvOPMZgJbv0Mx5Jpdp0EmS6P3aLSxU45H10SXM8CKYSTtbi
T2fhLzi65R9JQkrfzBDho8uh6xm1ZsuaBqtvQzaBWt12mRYMQmxlJUVqcgZgbLVt
ruwy+nhJPrhkZupGzgtuSFopMd9bKNClDrbJTRUHTiBX/ONnDo9jaQDHfIjp35pH
1fBG62QdOndJRMqN9xgEYnhoNW8ZEpNbcoOdE2cXP1myr65UI7hLXeTJM/sfP61m
bVgtHznf0+IVY/55K80N/GrMmGsGpBM6Vx3Vx7mNInxzZ03lx6cRiHA0bNGtGeaG
LfFuCc5t5JPrNqZNVAURlanQDaGCY3tZnc/UjTL5B2kkWr/3ZwuK1EcRosiNCYnh
8UQHaO6oj+EtHqnPMPKVewAshYGCe3RILKRbtDyPnfb8yio9RdwowudUUzKp4C3y
qIZnMqfJCJW5DBcUHtVPAf9UHYV6gmzyJLK0bfZgaHNnOAlKbdr7ByHG0RpHev1X
KsrNJD6dB0m4m6jWLqCUkzG9XdW4FdKX+0Fa5Rpn50wI21Wq1Kx6dbAhpu0s0ZUo
D7v95KzhFHTueIUNd4gGwZa9+P6QldQlHsnVN0YiVCKfsky3QWUncxj0VABcyOnf
94dDCAobwa4/tb5c7LNU8jTzZ3VW0xnTyZmjJGUG6E9/lM7FhgC5gxSkCc5Ax0dg
ohTx2auMt/AgnyXmc+EVWO1pIakWKRCS1kPohX24DdIT+DQPKXySrkI0u267SJDR
493ZXt/lfOXT33Id/tIhmmZvwt962/kOsu4s0U4mKJeI+BqPj0vP4ZiR+KT3Q7ga
cwkUbgb5kA+DgrqXa1nkMk5jHKmSLrOrlLFCagRMc85wD0zU8NVaFXeiR36tARX3
hrKLgqOsqcbHCYS9iEPqg2iZddfvth7BVL3defqNhVzhUFpQMrlSbueGOjNfjcWn
JBLKjsMUqm32RZEJ3dDly6hVxx2ytf8zY7QB5dyYS5/w0zNX8Pc2wU5DujmyBj21
eXsY4oQBqyv2F2LhDBEvPBCIZPMCbNbypsSbcRyOfbgktI1WpitlULNdD2wMz20p
l0JX7jrzVBnArnEfjgrvOb9SakkRWFv4mYtv18AQY4TxOEGEAiY5nK5mft9XyZ8J
9V9Xt3z1FgvsDqjlURoQx9CyoxuOPM5Cru6OIZeYVZ3i7GrljfjOl9zPjje3YwZk
YbvYyl6WYwl7gp22z6BbQzGWTz9Dlkg3qWXxmS2FwC3WobOwJIjebY43PkofhE3K
R2nshvRrJPH2NqlykE0no9BgyHzbhBQiv18ZDp9UWAyEvrjWElMJBxMLr/Tt5t+Y
4VWzpaIrkQditzJPZUqICocrRrh+Q4kzPQTGLrSuBjV0IK43AHiid7FGIlZoOW9n
9O3hJrcLnW/6rJIpHMd78Fmh42DAfpS48BsxrjECRm8BoC3CDxnJUj0QHHvPiJMc
UHfUKtRTFoDfnjBhmoI1lw8J6HPrDUB2qEa76oQ76DPZkAcpyyuNztxcUYHFTffc
oWZxcregKhE2KN9NJnNF0cm7v4IyZGoFflLe8DBKPNvXK62DlMHexWO8CoNiyj6J
NURgnoRltX3AZt9wECMXlwRoB7E40K0llNFioVnP3jDhBmsmMA3FRqAbjHiNR+xL
ckmsXSqSwEyWydwE91mo1oVdLjDB9KVOSmX2QqaHPkbsac/56E0a3LutW7J7qB+r
yWT5UzOud4LEVpboolzMRgQTeH+cc5RqJ1NGP78ucLY0YdefJFB62D6+j7sOlw0b
T12a/R8tYtrvZGfUjnD/ykp2/KsHrKFvNmPqYRiw3gyXP/+6q8Zx010HuT+DZgZu
hapBXP4sisGmKCzdk3J34NFfpyxGWmvrA1s6xcuxT9zjNbfB6s3GpPkC+1YqAgbQ
IqIqiDiV3fhuM/zkurI0f0hrFEKBglildHaumB0LLh5t4rG1UQGGJdkM9a0OfiUl
IbHOtCz9zWxor3dOjAk3seKxvhQe2rOr0qSHRsr9QXuHYm3eeLIQ9swAq3Gj6Cgd
5XjwOC4zhU/XyrFIh0Rwk6kmXELmxY+qf09vDuGaJpLFc6bNf20xuGYqnL8uKBXA
c/IPFd3Q0EWuTS+a6T0zSR2MCerHVUxTUwLf40JhdIw2xDoLh5CJ8rxo4WBaWP0o
2paP/WgV7yIayIwRCHCs+446PTwcXq8mJXNKox1yPqJAr5i3xqCBfRjuL+eqZze7
B/ytlgR8qaWeC+cyiNnEhVeida0C/LkOCpLSuk6T76KLJ2r9wwb5On3dRCmZf8X9
8EKDfhegRnxs0IGO/gVxfTX0dZML5lVscTp/qBn8lfoMkHGYZs/xOm1UAJJncOQO
NUAAlo3efgFve+iTD1UhbKXHbe5TN8Op3nyWeekqVrg9TQV3bjJSaKJ54Y1133qs
EAHkaEeU5nuuBYVaYnintEIYreB7lcwR1d5fZwZyK1Dh1lsUSVVXRZPtU9BZ6JMo
dVqksxWeuZTpm7Vm6tiKjm766kYl1nR2ItMsZ687SNV8JrVf4CG9QGGScNUnTxdI
LB73olQg+S/9SWiMPWC8kvlpUzf4ZG/Pi3gd4jK86/p3e10JBIhXavoxtfb9D/w3
+E8GbV7mvYozLJtTmHasZFiS/hfoEU+8A/wvTSoonpCbkSibY272AhENi49YeBS0
LRpKhJ4NC11Puc4Uhf3XWXuIRBJsOjmUtA0lNcKsvcqUL5mvMi51fqFu2q8E0Wfc
07WkMJfgcSgWrwsWcMl3jPJXJLtbEQ8VV916lC0xcGq2yjdTNtUBUmROqHHOagKp
iRh/z0SGqmFSq3AZ6Fa28RV6wO4EuEirKx8+1B7wT8A2XXrqGe4a86dbc7u3JxKA
7WzfESawCT2mqzPmFyTq6ULF8CqrymCmDNsp9XQLNam4hCWV14XholJh4g8AU1Rx
JxWoDW2rXXFV4kjegF62sE6Oz4lTA4xhTpMhJn+CPqktFO6e3gh6KPVeUhlnpPxN
viNCXCiK5j6ui049IXKFS9P3YHDcY0h+9XAQIOuFDDH3GXTsK6ej/KBNZbzTP80/
/zkibbF00Xl+z0wTkfm4JFEEFcGN8i2WReIN7ZPNyOl9scwn5heitNvvzba9xj8M
mSRhkktLs2+5U/5roGCC8/f37HtliLtfgfi7oJElb7Bp1BQek7byJlb8YQYmx4wU
JT9i6Yjeu707Nl/77yPNk9N7sKj3gAEijE44+irNfVVw1E7Rl59jKcLrGSFiDyv6
pT+uUuOty49Okgwv6cW/JqcXCKE8AY0c9vuM1AHoP/9/cjw11A3CYBA9kK5OuMKO
wzW9nt2xZQ3HnsdUZ1qiRXUB+SCNegbSZ+IO0jNl/6cO5ezP1TcrZNgTvuXAc3B2
YdS/VvDGCJ0hP4bfOKjttiTGtvYj0D4cHH5okoJpVcxgGd0rf41B6Odfom9AtZZy
UvoGv2Bug4pdtU5Hv84yRcGm4D/vBpApPQpM03op8w2SG/PRyqowBx8+CZzh2bMU
DdeLx7/L/Ob5fo8TlnFvhGMfJwxBJ3vOm6YiaV0G5K8gQ40AS4lzeXNQ6O2VI0OO
7AaGcllR1m2Tgcf5lZxwgpknVF6Wtr539ZoUxCnMyNZvl+LSYUYP4Ijs6KDmD01R
Fjbjbu25HBhl9NUTnnG7Kqir3Pb7q8qsvSvdCAUZhAjv4YAH9l1obZAgEP6TMijx
HXluToFkk2oCFPO28mRwbZ0NhKDeik5IzB5bE2MwLDM7Nb800c9AqBx1NSsCl8B0
9TEE/3MclXN+fVKePqWaNPdLlDuleq0ccY1byIf5jQpDYJ5+zrb197LAgf01q/7S
s9pAUlvXgzEmwBR7b4S0FsGddbdZ8MCH2cLStQNl4JFyDedaDJy16dslIdmEbYgs
DDkxAEl2XgwsFXnZem2vECzvOuxRwQqwn51mRcBPkG+xxelCxdWawLvmJMb/0INZ
ZUvPSYP8r27Ge93fzfS6Ym4M5qlnc5x2H4Vf+oJ/5J8qI3mZM9bePNT8O6fje9g9
gNnsTUQ7KQ1eel+tT2sTTXIuTfyh8nBwRSQle4zdjxG3GOZAGxp3tVGWb/qwal/o
O0lDclnMGYWra2jc7ZsdqYZ/svzF50JTDwTve0aS7tGY4NfFsz6UdurU5RqJ9BtC
uzdg5lB0s9ZnoqcdrUADPH5OX6MK5OQ6wFMqs13LQ4b+PIhYXffYWyUBwDPZAP0X
IJJ5lHGwAwJCS54mhw+h7e7fzuAfErpuJ4QP2rOS3FmWPU07fgjKr2zEQdNYE6f8
U7X/hYSE9LxH+D0+dyCZD4rGHZQUTHmjCrXqlRcfao7nvFHTdG+qM7o0kMoVjTbu
wLi+cznVcyzD5zLRzySVp1NW3IixVWWcx0facb351lWY0QaQBAEdRlTsVoMmYcpj
HNsgwf2W612iNK4wmYYITwYO60iVJgz2rPGQGnegkt5TyY9KVKbfN4U5WjCl8lBV
U6g5ePer1nnWP59FaVa3oJpLpXpzYr5ibE2Vr+tUClZANuiwSzPRqgCcKk1XooEm
TV9pJK86Ixqmyldk0jSgIJqPHp9zK5GV3260KMbsORKbxAwUt+1VHV46PqLm/bCu
LsKGMTX7UiTPKd6akn4zizLmsRXZtPhdIWaoS9XJDSrihUBggiGFO1BChjb52gXk
e42m4MWTZaxQocXD+tJNH67HQgc3aa7ORqV+UacONiXm8GHDCaHWI1IYuLDon13x
f4i8rmVYpAept/GNFjQ/S2sJZvIiegxMYt5EdOYVcSfTfsWMQB/kHqo1Tu/A9zx1
Pwaup+X01OtytfOvoJWQOyAQxpT4Wq+9F/YPIrfPZog8x8md/bjN0ZsJc9p5tK7t
ml3DSjYYI9ymVVIWCzcw7y3ulx6f/1b0O+TdzNWzk/ZHGjpqsu3UKPJ/m+c8ATLs
FWM9ia5yvBuP3qEUinRoiyd+MDWnU8sEIxOVjje5W8DipzgjoavAR8W6WhWxF8VZ
OyNCmR6llFNhRr2lCm8INUcRzzm6qcbDeoSfYolpK+81UH/WCvktvFk9f2TTEtuP
gckznNF46iDvXg1ufdvjnhXvCrKDnghqdnLIHsuKSVOXsgLH/J4F62UYBeNstkxV
Pg5li030YwQvh1GNPVvR70tliV2uhQ1wnldO2HYtoQuICCf18npFdnaI23UKeuCJ
QgaOP53XhtqWTe9dEXFezGa6O/Tl8zgAIMN9Mvq8s2wM6Q3RyzwCCYEfJYAkUTti
HXWCIG7zz71Gzn40De1+bHBoWXlq4zHwW7WD1h5O4GgptAklZXx6XozeykNVWjgO
mSBtWRZLAEfjfv+jZhZvuU5uT2Ycx47oQUiIIpx0GWgbCNX2PIQm43gqh06ksH9v
uQKkGWRGGJbBXzUwXJbbFBIcqy73X8TEHYTELxMN2wnQWaFDeboF4RjHOgVDKMFZ
wgQ9UO1bQ+gtAOsskMpZRp9cka8QwhNwIFthxhMVZSZll/Muoh4GFw+vchnXGpWu
VlZxeqhp30Ls/PMBkxpArRsuorpJWg6d/zqntvNrQyruR2aK0VoBOzqnVV5iiQ9F
gIobI+eKysV6ybjUPpQrshMof5ad+Lf/b6sdOEnhjRz38HcelEwEpXUBQe5HnzR0
KU8qd34MdCf4IdzSogYS46wKk7UcC/z94W9AdN5YHFulwBuLxFqJMgeKUHOwNU9A
eL6LQ7KPOWwRGDe0bpwMSLS7hJ+hZdKHspaTg27qFio6SAGuC8E9BrpOW1g/peBj
9OCk4FvWXZtGASbzWm2HqgeLJeBR0v6TxQqrGLwOfZ/Tb7HakI5NzV4epl/wyc0e
c4gFxarU+38Va43Ezvydv1b7xZt94TesQwQF1u+gtXh2kiJp7NTZY7oOcplfX2dk
l5mMoa1ha+gDo6gqJnax62b+l638n18WnhE9HYNGTlOsWsudWPNYCH/yNzbUgCQ1
fB5LxCeyw1i2k/UI/8VNVUd8F+gh6VQ+DDWCXx/VXkKRldDk4jhMX4STFxhCCpA3
CJGCJkcfjpptwljJYncux42FgHOIQfbTSlKBtnVo+mOnN1fVRYmOOJr5qfUXhA6U
T40PMhll8CPQxaTBOKRNzmVW9mFPzladshP4A2BT5Lx5Ntbs5Baff0LTeFpLDt/h
twYes+fDKKR3m232rYBJoT072VHyasIAaPJt6s/TRDd3xtRTl/J//M1GwkjShimQ
dnj5xt0G4CIpxZAIBzD66BF+EQTFl/e1jMDIgnKkw40d/hPWbcfoNy3N6q7eeF7a
gKeq05PSLpKsl/jdmDuQcaW16hsw9K6wkIpA7znJdvNoO3/QG9KYbXet++vYzzNd
92fNONzpVuPY1x1ycsZKnp/QrMhLH84GEj84clTuSLViDWB9tg2v1QKVJHtYOsEV
8QXOsU9qSoPcjuyfOWxIPzqx26pGfTjZ/y+rbqV87uzEp3yu1RqkGEll80jgrtT/
Ab7blby37x6kh+Sx1HZVRp6Y1CSrkYraWHXjYx3QiKjLKUKzdvk3wCjbzI4ADLOH
nQ9EKDuKriqiP4GLT19Dr15Ep/VxvptOWPPr7J92GCjsa4WgsFIoKKcP9CkMmZxz
3tjBOXvc8E6x6RF23qfDQQvoYfh8WvEwN0XwejNIXaSxZtyouMvJwFa6J+wdZ+M1
CJFN78OQQ6/zsh6/DYtfqgQI5X3SgqVjjIefwErVzgrvXOqwX2uuvBPtumdYvD1B
/zFC9Cl9LYf9v4rB+4mvrSw5uffSHXp3IvRUHRTzZOjbgj4ZyxFuPilx/1RDOzQU
JTao5OVF12RAAs3v6jkVM8egUwSeLKqcqxmNyXxRtBHQrlg+qeSz4+UFFjQkzUtG
T77sjXM3bxNi0cT00kOzhqc61Y1gUyrGWXqvNs13LtDzpxFjJ4a+0uodJ9AE0QkB
6bn6co1vfMIVjvzQBfGNuimj+jIQ5oPExwdO81lbgYQj+iCcVHyihRDjb5Ml3456
Afd18uT/3H6fMXfTHafBLMzEGEzGBbbc81YDH1hawxvh3Oq6jjiGxI5ShezBFLBk
hkbMFDoGfVVMoc9k4Xjaz4Ucb3LOZPV8Yrbp9ae54SgLFU0ZtHD+OlLObQtlkb2W
0VWQVAtkjklL1KB2R5Mh/77x1z72YMAx5Ow1nyTRQrwqrQ4uKN8wcV9fPtQMBPaQ
/GlxfKeQreGFnIUyaLEp7ye2e9DlimI0UtO/V791k3zNHSkzu2p3rcHFjbKOV7Wj
9xJSD7tZBiGIZUL5iRzMldaJ4H6fF4UChT8zyd5hKFPm03m+XLwohzLhyzjO2UNb
VD07ijtaRypXQg8an8borkKYH6wkAdqPubgqX+fF6Vm0dm1y18pBrIr6FTaXidNj
7pSSQm0rqfEsSyXEJQ28kGWEKWcR+qRTWe7GzNuim9Zgocvon7QPJMZ29bseK33l
hMzDz191mSK3a7yzdKUsbuaA99768VPO2t+5eUo/XmU6HQWwPG2UA5t3E6CD/v2Z
uZ1x9K65XhgZls8aprBkeK0bPk4LRxCXAcSbKN85UFfEDpOI8OZz82GS/Aw6zz1r
VvJWEm7ZCOoG3nfIjv1vNfKgI8yRXTN1IYDd5s5yek5uDbJ7HoOk/XSmsvd6srb8
ZlrF0IMgpKuNDwnPJjBXsuJYjdPUH0iY74tbtBTdBSCvv18ah4fYRGJ6fudEGHsX
KjKrCEd5I0VEaRBsQv284nrPNOtKAzBKJTwDunJVZXyO5baMS0xKUnIBXKN+Fx2g
dR6dGJytsUKpgUXdQeMm+70YZZwEIe7Tuf5BB57e+FhTbgB3OEUljdkesjOIdPMU
zPF+FjXwxPjTUbWLW89ocaRns6KIWptN8CUUyNDfeC44gnEBt5mybAdGbT3i4Aaf
X3HEh39yEo2Vmznrf831yN8v8qCn/hEkoMkVlABmG++eQ+DZkw0pqEfE7MAnQlEu
FCIxEoZ48WXkDFPVrSXmmlFKScEeVxhN+fKx9U5Lyp2QQfNFgQeRQgadw41Woq2T
IlIPgyESNhQcB5Cfq3Kaw4NQHNgpnG3bhpn8usZV67GQmqYVUzy0sa/m+zOGGKxf
nKb4aHmw4o4Soj569CrGvm26xuX2z6Kn3n4EBV2jaqNabrwUcIQvHoFb5ovjxDWq
dQIQUAUiOyecodrI5TVAaTDOikbf7X0ABRYD80HzTvoHrq6nHUdCVhXWt4x/YkkD
DfzBq3zOsEv51oXU1XCrfhSqUc+dZBfdwJGil9TkaN1JD6GTI/3w0csRs18EoO3e
838bTKtQxw3/4E+gZN/L93C70nFShFH5aJxxgl8BnG693cdxW7qZzjJpw2Od0IGF
gaU2c8A6EvQpoPXuf21SjqnOobTq97y9GEET1syfRaLbvZF8hTZ7mClmO/OPs4W0
drl5J1mys5qjXok6WG2PTF5pr1n66Ir0zU9J58XQklq8iPHcmsj4riepBB1toz7J
E3fWdj5XLGv7zG3VZvGP1pFWRVwYu8la1wz8JhMk15MLo1ifENEPbrNvLDh54b/N
C/F04HUT9vBUTzvIUjFXH3ghclXhF7IJ+n0FxrOL/3X+QnQMUCi1l+N5KhwRy8Hd
K/IYvHHdwMjZGuKpDMBFYBF+O8U+0IRV8S0X9/iFG4NffMszJBrx3yuox5VB9zBN
Esv0nyYCO/vDkvUse5sST7k/xeG1rx17TUGKInKX6N3u+4t+I2Fge7TN83rR91y8
Pu2mVV0mZmyBvagO41ZIVR5tq8TeBVT8vy48WN3Qxy3z0uKy7NHBoeUO/0QMqoMR
KIojD4XKfivZxHV7X0yB/FUd2o43x06oIJYycnxzFaDuV2+dNau/z+Be5zv2RvA0
ycaq8XQTOcliduLSF7uJBgy6hgHt8M0cFGw0ERCnI3sv0yjRXWcdKcnUAUKTtZ6C
h+7ah+Cu1UH/LgD0Bz/qai8KxV9slr5gDzmmrmRTySu7uhx6L8gS+QProHGXefFA
ps/3glPznwGCSxGQSuKIzPEt+XfY6UfB/fC4EKBtD3dMwL3DKo7SOxkkQwees8v9
gYH+iLjDupgmFISoZsZO68EzQ0E/DvV2JZ0tljsFCwkWd1Adc3alwEfngCyjRSsO
fBoGFZU9YRTFwt4sP+4p+dF5tT/RVKlxjNWgRWit6etF1dXXg3bRyFfV5/XAkLiu
wyneeeEILBdLE4g0Xsm7liXV+L+h2Cm52o7A8Zz7cXwtTNbcmwsE9i5N5WOdWG4P
oNvjzl+jFfBLiEOIbBv7F7ekS9LLNBY4kVH01F2Ox6JHK8TkRe0OqyDsvZaugdfD
EniDC0aWhcT2EuwpAdXCIPLDDUHhiKSPDN7yabnj0v5gemiqf7bJAAA94cTuVI9X
WDByhxKxO8JzplCZt69qKrtOVIHJnn7LscBSK8WwAjb25Yg3+cVnzuXKxyxQ1DW2
YYUFnUO+L/QKNTf5h/JiUVD4u68pT3LLtUhMsBTj77HkHXalmmBw+A6k9VxZ40JR
mOZpqvIXjWEKTHn3Da3WlVwUWuEQaiQj9XOtZKWswLNHoynVYMx/cak7a3pEV+en
8gVdYqmpfjC0yIbAlN5oIl/8zzIIPUu+GptthpsQLARdN80+So2lkhHqOutp+ua9
eyib//Gw44LMwfdbGPZCxk8r/siLo8SXSrs1VRYnRE8HlDEsDoHvW3P+q11zHLFw
d5NzhuwFhrzdoTLSUJk0xkfeK3b2obQa5Mqv5S/YfweFV1ZkQelm+IiV5kx0EndL
7wXgVwQayVsrV4Rpt0Mxz+Xqh0qldxsd4LH/ao/sD54ky0y0uGQQjD5D7dueXTjq
bCijKVkEYTCiQJr1iELIa52nWnTpZ5mymy7/OAm3FXPXozjg62dVlNPZLbbyBf/Z
L81I1VhGyJfIYpyTOSQQTU6FMzuMv07tRqXjiJAMCeZJmOcsxs7w05LkAEGmwkqq
/EhFWqsK5Kh+vSoW0hnUqa4yPDiNVjw/t3e4mqkJZOz3kvOIWf/bWhWFqFev92Ub
87wYpl8oW2VRjoRukl8yackZpSrmAEheJ4CCob3FxnENqA8Z8FZQRnB063IgP9lQ
RlRyCEdPCB4uV6mAs91ONQJYbDupwcFeYOiq86ZMqhw/ymPXq7v148KPZHck/Osf
pxKWgAvS2D8+6ZgaOCEXkDNWsyyg1X94ulj76gWv3Bpb9fGoU5MX1nydaKyOnj5a
lnEImpDGjFfAeBuyW/yr2qbB9/OsaieXG2Lcqt0L8n2euqRxU0wzklBgC5Z1iIOx
oUvQV7P9tyagbEokGzqGYlqOvh2S45B4K7iAho2Qa5fq29ZOxhs3jx/NJCNdIrk3
SqZrGEaTP0fvzPyDyeL2Mh1eTJAtJZ2nn/4jGD58hYXVo1tsyA2YU/ydUVDzfIRu
zaQ1CLo2BbzQ9MvQ5QkCEydMVZClzG60jwdl6HrSBtk0Xd4EiRnTU3gKaiX8jt3Q
+nB/1bnTI+OezCymFy/ZrDVsKTZIZgpZ/WUxKdUpf8E8m2oRb98pq7nxmRS1RTxS
Tj1i3aOrjQkrx/cVj82nbbs3b1A6JD6VQvQocgpMo3XQEfOTQ5xaBFjKsdDW2jey
FLuxNclq1r3+JpASLeAJGg9nuGGudcVxC/NOOx0xd6xbXP+/sNvhTJy37nT1jTup
a2TDfJdTRL0H43svVuj8rQ5ERBHEXYnQNmVPZSFHGET8pigPcI7SQPjSw3ymRfTK
9CvFadmI6Sj9X8i47ybz6V9Tu57jTrx7su5nxRQQLVpcrKxN96D8XvAvtUWS3rYE
v/YgTpE8ktzOJr1sEZQ7Y0kthZgqn43Qfy6xN17R2CXEuueE3ROugG9UmpoGJewl
rqL/hUUb1YuSjBbX398TwIRln7wk+fkl69r8sVkwhbX3wcyusWhHX/AYNik0e6bh
hvpuDGlPwdHA/TxHpMYYGI7FU/3yGnHObt4fcNFWrcxiaEzkRcFe7oKQBeuqrDt8
MHf/ugPfqYf86dBVxkN7ww3tCDM3OiF6Gt9ilgwBXuTNpOlnpkI353Lr7vbrL7I/
VXHBploQ/1PGstv5y71UIlrtG9h/74SKO4pOqolTjgQhO0QXyolpRfjDgHB4ANFe
o/4jpU3z3Q7pO0tXlRb2JjwbrPZ7r8X8pF5hMoRoXJ/gdLrn0XWNbWMLWuZnkDdR
bC3cohOoqHO4mklPqcYEMMDRY7BEllRmpudJkslHOdRYiNRuX+k8Rb9vGqUPcbC+
mLS3t24b6gNla0ewUVeUI/XxZPFqE+FLMYXlGdXGqGR0RXO2foCG3P1HDBmLE7OD
/8eg09XTA7JZD5KWgXWvnN+tMkCI+jPtOl2TKe3ZyfK8DlTzoAJGPK7/r5tVNUrR
fzzrpzyALkvG/f7MMwDMG+ODbaEt58xBLc/AzPpOqYlT46kQ91bJ2P167gZCRH6B
QF5p5GkbsHcIcQoviRZhc7ur0zYP0JKPcXzUMKp3gvXkI5W0wR93lyuryh9m5qux
/htBn6tZQ4RIwqkllMpOD2uJutGvGOCkyxoU2uphi9bp3kAwaXIwqlKK9rDEgJG4
3MNrVRg40JgTDFlWcVm31awjy85iOT1ltyKUwO9zK6K3hzV32jV1QYVT/IFNthLn
4nF87brS7DwX2k0n8k7nb2LbsLN1uMiFOZXkrzVpnYY8+gQUCV3RuMZ9FAFW1hW4
U45JS48mFhcucMcfgNMPSqst7+gSNDygkiqDv+jf7NXg/QhNH0j/YIVQtnu+aAVT
s5RFW/HuhODzk5O/VY+uglFCg7ebqq49cOCNGhIXTbtp2tT9BRiObDQqSoDw3KIf
Q1fQtoDIARgLHBvHCYIkh/ozRFcMIIVVQPJwjssheqmBwjYe4spsE8fHFj2/irpv
mfhOMhY606pMYwoPVP4uPrvBKuYpaVK24KUByO7RuW4woXxtYACrb6+n7jRCY9Aa
1FRRFz6Sq6kiV/rr4LrVPQ/bin4FROCsQ3vtzyASXkG+u/sBz44qdk0zdXHXny8x
BAq4NdN+HAh2xnLCitqn+WVRM0HDFLvsPltHL4YyFQM0aBvUiXOaxKy/fiXXf7dI
6ZZoepIM/19P3iE5iT4zZRZhMMNSdMTMry7+sMGl+dJD40vpJjP3SA8KdLnUDphF
QAMMFGtogu8zNkEBOCzIIXg9GaU5xqoVP4oJR3+6ndtl8ZrAryoqC2JDxLzMOmlt
O7dgULRijgF1BjXF1AWoJJrZJ08MLXbKqsQstqJf+BaXNLQbHtluFwHCdLXoI1XO
H5pwqUJIzg2RvxCVD0joQjOTuavYccYxb+MDNqnhtLHgkbsZgMBQEpRmOhP6rpTt
KIAm97ew1il72ULFfupZsdTPrLQxYZLBgYkSXP+hhwN04JW9tuhByUPAK3QTNMfM
osFkYtbTRstoIwyYDDusA7WGj6eB3uonWabpvWTouQhTF4PJK/KyrxwnOPknp4Ib
/0m8bMYFPDHovJQ0RHCRZKiahys/ni6md9okjo/SLuWmEyhHtVfLEHhBnsMs4MZf
4lW5tING54dtKZurrKKWO+KDP6+lvmM/vjjP57CJvSFadq1O+EZEtopkpZ0TIJZz
399ZxH6tTMMoDc7Lr1T6jSZbawu5f7T0Q6mOw9Et8+ETkNJLJTZCYZLC1ECfdjAc
Jmmu8ZLL0QC7GZ4LhVuoguRxBEz6slXl0SKWsssokGLebyeci4tiocEoDkmN9Ebf
n7/OPo6yadWKYHBNP257UMSUfV3DlJMKaUjUU2n1c/TIM6lHzsxkseYULc2Ec9Ni
Exzc0iyPh8FdBKj0JVYAUL+DMmJWfUyySPw8GTvqUmlqerQG5h42KW7NfkcS0lP3
t8RileQii4pym1uNw0MD0xIbhy2dAHgIlq/euA2lHNjBfqB7La+s2gJb8U4n7Uru
JZtQuQ+aCwgT4Wl8iltJ0ic3LME2P5lB9ZTAXryU1jcVgC9eXKsKw14AnfIVidfi
w4DhTFwo4Qt6vB5IaXovuQiDP93ihGliwbVVU61WDVUqbLEAUejDBySiyLFuELGO
eMNDWB1iY3cnJMbrOOewuh+hqfewLokWcPtKoWKjl4L99E0ajC4qNyp00xsLrxbl
XIdv6N6++kRW7FgdwzPoXjmIyM4gzbvNQ5VUE+aF24MxGYu4YXgIOz2I9gSJDgLR
2EPTEVnKVMZEkHDGHivIilDEC8pgafqmhsgv8yg+N0KU2hGOfBXq4D2W6Nav0oFL
OhLc+SujkMaj5on+4n5Hrvqu8cro1DvDEjy5gNug0ZvoSz2BV6twBUakPe7ltCk4
PmbEjsA9xrA0kcMAXlZxiY5GMbhayxzF7I9i/L7HlRjGHHtSmQ5OXAKEDLzIBu6W
Kbe0ruaVUwmDqK0djmMC0xUDOHAV0YuvT4+desRG0WxqyKbn0fqoXsosaOcrOAqW
uW/ktzrAwlu2oypkMnSsHVsri9DYaDKCIOpUwbvALecfESlGOS81C6B3TjBmUBwr
yGZ4y9G4JAVLcNRK3PgSTI5iV/R2Gly8qyp42yZe12vIKlRIhldVFBLH2qsM915D
9x1xinLe+AcrIzDYjWE7EzKCVrxkm6u9KW7FGv6HHQQqrASkuwshcNc+xoSD0HkI
BgOntjZVqWAme/SU8BkktXfML+CkP7CnNJKiaMWhQWb07chJNOvbDED7yq/y6oDV
DuwcjLfy+1BpXO3pJT4p5ZRaoePzGShGQlYyqMcx20uDBVNB/MIU8YZ6Wv/ShyO4
MAwJoCAfE6QZH9SKh8p3uimogx22gsyzgYAy65rlGHoyw0nA5++LDTtXtM4RVcDm
pMHeypzUs8BXUUlPciq/BoXXfjlShqTYIrwRX0HRdUsYjtjtcWwv+xn2mn4M2b9F
Szr38UF9/jAsN4duNQPOFdfUkOfV9+4NI90ndB1wiUdCMby9MeznGzgmAIX2yktt
RKkOG2R7UmkoqOFY7nYPVLEOWvs1dVMnIfa4NI2z90BmyHtUe/JAGmqrMmNaUVMg
eivOpfoFtCmlVJjQMpH0LPydhG2JTXMjP40B9M7ayBzzITl58zpYM+l8CRxAynNb
HtqDeqnxPcTok0dRBHIMG7KCkCsT5MhSAzWAUaETMQEOZ1QSkykaQVYrd5uS0pDI
mFYKZUGqDFz3kXwCHXLxkhMAT2efSWnFxSCG3WH9qfGwxTHJ41QKR+IotBHKmAuv
7Q/XP3tgRRXMmiiKgj1MDZ2U2O5Y6Fh5Y58kHuP1aH/BTiMsUrfs5RgttEwBntDo
ry7iDpCF66n93S7QAYJRhUtWRQRrxp7mFcLzLlOPg670VrDyHYNzholaGcKs+qyk
T1BaNaan9sdSdbfETNOsxlBvno9nbnalT6x+YAgFwetBESRKUlNSfSoZ9sOyGdpD
pk2lfs2nVQYHqwoDUx9xczIzALPjCkCdPgVd2OfennfSicKGdsln6MAldIrpFxFW
e8ktW36tc7M7iMT4Ihvq2nv6Qe4llNzjKvG8/dmgYUSsbAfG8+7ssV8xL1Pql7UY
tmykrpRlH6qkUIIp7gTFruAnmsWeoVLfhOkUlm3N20Z12VQgi/57BAfXYl1/JJbp
mJpvnj94cx9Bg1/AsDBJHGX/mPpAYAOJMb2+pJSA6GCiDiirqW7oORlp/fw24jAc
LgA8ag5fSLP3wMA0C0QrpsFDbfo8OM/46DkLC5SL9wWzg8VgXCRE2dS/lPztURP4
AjakCyIsB2m7d5WjH9B1Qd0RJy+kJU+jjlDSCWeVTP0cN+y6Fi6mqWdeks86ZFts
bMYcqzFSJHHN3zbTDPgN3FGcbSrKgtyzFLOvvw56iy01WAzaFcP4ixCkkZK1EKIr
neKNQ4ALwT9pG2JE4og+4U84aHhwgoBHpquD7emdDPyX1WUfensKLYb1nxccyrIo
owIzs7zgZgcke/onqIXIJcgVXFB/8/D5AsqT8hveS+g271v2hicWGrMXxRtdMDs7
CDYupKmX0B5ghOj1nltbnK+R4ZvaIhPNG+zNlUVdIZPhca0SEo/hMYWGpDfYLjck
X9BXRx77QJb/SeITe7Y7alr0+1iyvWSPn72yrLTt6UBrwb/GCQmsug+vDcRDrdiV
5Q7AIChIyuPd7y6liX0TWHE0Og9kkqgFQkLUbGLlee9MIKzAiNMKbxqle/FTgnhQ
KD66scdV7RClSnq4/Briw57a42X+C9mN47Brj/bVKqhS0x9mBYb8u8h0ImdHQCqc
sH32anZ2EUM2igRP41xZ8ujMCXGbyAxq+jXtoPtvpJOVzHfFyeKKRlv8WeWYrp7r
LgFngT0f3TrNb0vEe0bBkNZYUgCQ3szoD6ylJgIKrYLh1L1rgpXC38+VT4NkTC4N
yCf7qqDs+u6Z9UKXiNJI2JenEiGtjalGqStyq4ogGktAI++0jl1KJJFKaokPmQ3U
aQGR5fQWo+TDPWpGXu4SrVL3HAH/PK3E+5oBRVJsbsUME4MjcCgPjBPZzueqR/RA
CZKHJNN8ekMAIi7jecP3ULTFXeNbM3Ingo1hjoLXvOrYL7fD4ysapvEV+ljAhim7
DZgt3lrTVx9Q8ElJMNcto2XTWn5PO+f+NiLVI7BYYaW0+FkqzQbvEPYoGFFCyQZa
XT/M4rKjZn1biZSfSYY+GL3F/LWZReY9rF9QklPxEhCI+UxDs0ThN22mJzaqKpiB
BNYInmzeaKYF3PpallR7/DubzASs0hrjURE6OmgCeShfcnUQ45Ue82KwC2BU1xpU
jmbxjzuX3ATFuyfUa0A5SDMTZeLtjnU3mJGZjbt+ScJyCM/y8fr1I065S97Y6a/B
/UN2HfhAPBYpOIZ5DBAXBfLsTc5ugv73aNOyBxplt9v0YnxlDSV1j37fmxGr1b8o
08ja7wD8jttFVaBY4uZhLYTBiXXeJKxdcoVHs4BvwcdKI3rHzKAawZYpBJjT3lUu
/98ffp7pRi8IR1b+HwPOLpTUpb4YVnAvKVqBfxMhmqTlwQ/18nuL1jY6TPR0i7s4
pJRboB7FWnbmd3xBxwLvLq/C7N/9cZalH9iNKr2CV7BIM4giGR8rzubGvw7Un1Qd
Y8iSYiMNpi/qvhaowkOFEZfRh+X0Aoqrih4YnPFVEe7Yw2tVsuuQ48vy4vnE8ews
sQf/GXoVz5Xn4w4xx7hhXL9sS72Bn7SqX+Uagag1SwIWb1SjHk74BxXBoeCmjoxs
iWd78aPuFZmkfqVt83SiWvhtmsulaweUex821z1jYsLpzuUlGhpz8m13/j0AnXsp
FG0l6zr6u5eISBTP8yg7T7+lLajXFTiM+/GodFP6EGC461o7KBG/QQIvlgyrB7li
wiZ0uLKHtD/0EX/6NH2TT+tzwmw48zc0mRPl6mEjck7rbsl/7/HBDe9fIcMKPpqk
3NViL9nu8cuNOt+qEsdDQpUUGvk91CbQ/9Fg1jh0S9JCBosGirZcyHWTDS9QGymW
EA1/kIPzwnErJJbcEPSKEanuG2IGe0AjalCHUhm79sZQCwjhQcfP+ceap+tFBRy5
xGFD3ebD+V8BSMIc9Nb0DgRuJdqI8WbKDrWs5SfxbE0PfqiqDSfIGK+9s0qgdfZS
SdpMaZJotURxIDqIKz6Agn3difqIUWP1LlO3w0ryfCrKHKwaWYvocgG0E9BulHXe
dTNKXbrf2mog4gAUKcJxld5gDUI6RlVXrZFxn7RKC6my79gy6bsA5iRVerLAx+YF
kqI6Ml8w1Ggc7jgZYH/U2cDUaQzvWMh9CajKlEEsodoFtA+TTt3fwcZKR8Kc/C9G
H8eZe7dxMTNzHx4/oMeufuuddfXV9apVblraDPEDQQRsREmaBRXDP6khtjOGtLwe
R6TiBOZuptiytTHJWNTBX6jaRqjhOOb+639toZhDn9t/Lv31nxP1EjqVM9nftStw
1k5MrI4LYxla+aVwzodrgmPo3pk/QmPq7o8/138+iDRKA5fK5PMkZnQ3tv39XrwP
UckHRtHWc2qF3R5XCp+Mlcp/K3muF3v7av716iXR18b+lJ0GIM1VLLVTg8qLzcfy
j8NmEfZLfbWXPqe8Ru4aQ9/ktzByzAPjffZJwVZSh+KWCGv12bLAb6lH1mklsBpE
z3WWxb7ZuD2HoLBioQ81IGy57f+d2PYf4ht3TL20TqtebCxX+nFLRgAsjxzLHhnR
CUF1vH3UqHpJt4HrbdOe9QY2my1PJmH3w2TOHfBKTNmAe80ZVDuZ+uCl2MDk3fJU
3t8ZBId5UFGDHbxSH6wmY7EDlNEmO7+Gg9U9Or/rkHa3VIzn4RjswcvJFHOU+stC
TtzkvII/ay7KPmZjtU0OXTzClAsO7tjrhQNJ5PsQpuCte/Un4FbdwB/JQbTRA/Xh
mJnQDdph3Mkdmfkb+ykuhiJkQEq7ZX1CAvUm4UGszCH4xoOOtRnn0Tl7IgM57Efy
RGz3G0equgFZEgWriAyDDK8f3h6NEz0K5wvsviivnmbWhmcCrGW659Y/9D8qRGpN
TFEnEOAGgNFxNxCTPzalggCYJQv5AMnXi6sEH+TDyVJ8xKvcMOcgVqWCrf4ZhLA/
m6Ni/4GAGzo3UaRhMKa87CW2gXt0ZOupKZc79NAxbrlI1MjtyCrzWLqowqL9Vpay
C/MJzAIH2dqo92k2CsVjlI39VaQ3QsqdCmhVrwwH42KvvNGmXZucW1sLDP7DnszP
W8oDc1SCW8jPhqAirXAXCJoBUcrn7rm9q8fjbzfD+4IYDVhOYN5PJEF683so3haE
72i7W03Zc3aZEdJilvHdWK2AXo7kvE/9S8QrJIa8ZhIauXsEIiO5qAjcFyk6deV2
`protect END_PROTECTED
