`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOyACt4PJiLCsmBkqVlZGgkOdDDH+WaGnxfqmizvAJV7
22nrE+NGbEXmfj3smcx+UMx6UYkkAZfHJV+o/jKupqx+1PlzQ3ksMqgttuwIhr4K
a+0jHIAqbK4/zDjceucY0ECzujau5c+3EtvmGDpElCX5ahz0Rf30xujLWGpoCrx9
fXllQ5EvaG/ONN2WllOU588JZYy+EfD3B9fa3RJvtzw0AO5Mg5SPUMngDjH6LZ8f
`protect END_PROTECTED
