`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
7wNuHkqssMBdmMBADDhjut0wAYpgNiYwcdVLzStLIlyx07ohIMAWHS2JvHKtmwI2
ylFMf6wdsv3y2jS7jOhIOeaZ87Ky90ZXVwPwpc9ZTVB7xBnllv4ynXMH03OypR+v
f60DY+GOWlHwBA2vQZ4BMeTZjGBhQlEP8oKHB723lWrkLoDuz61mwPplFmpFZL3C
H35yJI7oCylS0jAD2IAsqEuFq7jz8ZQz8q4IDkHRcl2vychZHYPNdSXlNSSOD2or
ZZQVF+I8FO/MflFJEoFQkxqPexXV7fg/Y2D97qBVVmSHL548RA9IHHQM5v+WDXer
fbzlic+rDxYwJKZ8X7UCq3cbTUD3F2pLPO0HCHs4/lxcw8eSlN9KVw5QNhTX5uBE
zoeTZ7HD/1c0XGHi73NxW663fa74ocy7rS3BOK8+Xa4AMqN+o2onijSjWxPKQsqx
d32pOrbtsMvmudtXFPoN0IrHouVA3P5lP6NW++zilDnkXN1Okj+dy6z4tgt7Aa7T
oLTqeGZtQlJO7hmq5ba9IXQslyiTOdIEqjBl5HOy9ACIgwU2gyo0Ku29RpuhZmUR
OWwWMiyvXe/43lnjSJeTdYp5HPeAXz9Veqnk6wc/YkQuM/duOEwWZ01XB5D1IgA5
2MMqaw6QPE5qKqKTgyZU4FCnscuq23RFOHB7N0ySnLMk+KwEfuvxM0ZkWq+rJ88K
3QXfXAtHgBPbaxe9eJ8q7zwy8wtfiY1mmoF9fTvjZKciPAg8bqZitRsGMZyZBk9t
nMMRnx6Uje4RKYrByA3iI+V870/HqL1XvVmQ+IZBkJU=
`protect END_PROTECTED
