`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePe4joGAr98o1ShZALEKlur1K6QZ6LTUaoGNxXPq340Q
lAePKpHoX/HLLkdyutLC7YneJOSd5fmYR2XMw/aG504rPdusIVALyWRRKHx0+GxM
svodqjqMm+z/pCDBaZW0SFYfMiIoirl9UhhcGoub1q+Y1xmY+kU6vyIalqwl2B9u
YUqhKzIX58zP9VCoNOyy7ViNm+Q98xD7grtC7QGLKzDIyc/BsgP7UYIkL4jiBasL
wqqF1KEojRqotfHUpK17OUK2aZwNeBRaGguELprRGQruC7egePMosnSMlums4rvi
U1MDV3aI6kZ+n0CDqb5YHKlk53KX5QwqBMejlCZSamUnKNHZS2DK1vLaUPbF1QGs
aI6AHoqo7dqmrFauV0bz2xHCPBc9CHMjIq27lg4hPD+ICOqsgF4cKQkhSD0w1QS1
hpNenisxMWAb7UiWEfdRnDV8KqGCaMnJrlN8IV01LUi1YmP57fWclelDr2RH8fzm
6wIhba+Iz3fo9rzGX0yz+c/cLuWW3I8zsLx/vTbhHEGRbzsAfSIIF1jidY5qYV+v
`protect END_PROTECTED
