`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB+XFG5TtK6ZHW7UP0SlXWSvutUmGPriGU0UZNhMDH47
pbpSMPMTA1BTG429tFHojl2jqChKeS4rv3D00qxukXeYd352yC4xVgGL/13Kv6hP
PnBDPZV1OmBF52nD8YjdbYexgEtw62XzxW8HnxL43jLMuUxRZFfPLI/siCErDQas
aAwEIdTowfNk/mnyucbyHKpdbauZ2A0t7ePbOBrPe9P6O1JKwCjGjEwvwrUXPNS9
Dcx9nPP17WWGJ1HPi02uV8hNJ4HuLsJx5H1Z97g6YPdUMhzblU79LG3ywmSbU5tE
FA5KeDNzac4NqqnbSL0EjX0o8/Vi7YaApocGLacpkyJ73QfEPgiqfJngjSaHUA+H
qYHR6VEshxxdIIt4BVRLoIGKkkCdd2ZvLiiGkcxtX0sRgqk9yjx7NyL1TPrqrOmD
lYZLvcsEnpkQIVThWBoeoTO5+9N7LGFWmaN8IoK1xqUWyiLCuhXl5z2ldKTHzJLm
`protect END_PROTECTED
