`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNttXZUilioKtwPRFfaZ/jstnpbk/Z0t/Yfssc4n5UXA
0FfdyjFKf+rRVNMioYgrBBAZN2BQjhkUaJtiLZwwvdnqUkzf+mB5e+ZoxGpZQpan
fO3Uj/It5i4zhTgIZFEtIpDO0HQJv0y4t50SLza4dasg/RzxUViEQBQH5axvLd53
22AFRIMcwpgmb1oFK2kR34jODt1e7z4xSsO8E3TV27Uc7R45WgVTWOIrKUufcOTH
S3klpG1OpGIhQO6fAyDSDZWAmG1ABVY83Nf92iFpXLadojEN8EZOaa6n+v1F7JP1
0b8UUGrJmMKXkOZlpW62og==
`protect END_PROTECTED
