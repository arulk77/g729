`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePZklTdELEupP5x0LZjqeJfpj2WEvHvZ/cw+JEUfMCRg
+sayUwGFn5NYgUmu/YpppvppQazCC6/9+UJXNZW+jlg7G0c4Yf2PG+ID1cK+l+Lm
6bRVlr8/oWRdGHfnph+nhpA+eWFmtsgWKXZq2Illp4M5NpQQAAg9vI5yysrevF0q
N3vFFQaqF8ZVm67fS0QDkTmD3C6BuSXyB9NAbRlYQIDgjQ0ilfSva4UeJ7bEs3bm
qYHoCwbRz9VEsHsbtxl2DpMcGH1GsKv47cNRzyRW07i6Z3xkpIi+4QmLi5oIlDca
PrcL31n1WYLP7xfQK1sq3YMONtrI38jSuxmQFZKCU/ns5C27pq/5MSKSLTMu2ONw
wWaHg5qwOOLaz8GzDTtf/zc+iJlglQcxpFHKgC9ldKU4b7jlf2SMQ5JQ2ZJxO2pi
0Niwiod17yxV5TUTJqPujJFS+0AffpMes9S2jfrh0UYQ7UWGlgiOuBq9em4CIktL
EgEpToatcEy8i86w20QKOOE3pychH2rHu0sSwEJ5b+4HEDMR8BCz31HmyPyOyQ+R
/dwq20vw3sb0hWmS2QPrQbExr0FO6V8f9CRKGxYGdIgWGYP6baCE2MZlRgsucIpl
`protect END_PROTECTED
