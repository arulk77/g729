`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu417U7KaiomzFuAchz20kO+OqdkvJqetgNDNPWLhbFOSd
FKuiyI2IyH9EyQGxiNDW8aKpXD3KQL9zAszkBRixxxrGwXyULpz/JIUEak8uMWDM
+TCehfQB7ceqD4a7X/qL9phrrXen+WmDwxVTMM9OFXfzeiSScfCowoOGN2E0JsTP
OMbaHGZ0rs5YNEvNBJhKoVSlNIF5zDk1k27Fg91u3Nh4MCH81BNNdYU4+b/kwLdC
TXmGzn2+NACUc6mq8+78QcBUFMd+EUnfM5XHnTdWP6MA6PEVi9v928afXL2+kO17
fPASJrJass/gR1f7DNtzojqZvQVhnIRGL2nZqnJ46DuCymLxGExdOixnwqzmtSWV
D1z88NoZc9KbTuYt3Meckw==
`protect END_PROTECTED
