`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNU1h9vOarYlkfHTACqHY7x9qvQVikQp9Zy0J9AVhwS9
Xjtu3qC5wPNNL1XRmxQ9vaKet1kLTyLT+7QtDaEtOrMUE3kiHuuUoXuGTwzs5781
4Gbe0Fej9rL06wt1jWoSYq2bPZ8VikOTZtU6pkGco9n3kkpbKTO+ROqK+O/WzpXS
4vsyZ5ytkKniLxFlVH81Jg==
`protect END_PROTECTED
