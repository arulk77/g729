`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xuXqEzOaOx6QFrr4GUMRhc66J+FBRdu+dvKZ95kQkyH
TTPWMoN26VxP85ezIom8Pyjan6a0hCx5TyvFIEQzS7osLyWTo/Lk5O4t1oOug7ea
5fAcugAapgmJ8lMLlx8oO8ZskSwvdl1NncwgDzDGd3dNd0oWHaV9a5C429f8T5E9
tQNhbg71M0a5mxQQLm34/tSZy+bjGkC6PSpV/ettw8MnqXMmW55NrZaniqXbOlLx
aBdPyjgsYKGXS3LZ3i5cmhNCqfcE2pOna5x+tovxVHCoe25YlotJQolanI7lrZiq
gLbRBhZ0XlaeNSs2Hcg+XzsMh8tWsBxNT7sg1Rnwpg5du7Yks+KNiglqI0KLUdf9
BFquj1XxYmsv0jxu71/Ureywq7R1JZRV76pjoyKJBxY1ZmEZW96Ldksx1ONLNWud
Kpy5pH0tnnPtWnmLcb2OJskUehephVIVZNArT8o7pgG1gSHXI7ICvmqmBtSVNqYG
`protect END_PROTECTED
