`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL1MrjN03HQf9alMYicrBCd9g2eVdpy+It/zcyWG/zQG
2RpUH62+MP/VPF4gesL4rAyZfl6HbzCXxk1iplVkkxJhJtg3haUAEEAeib37/Tdp
bL5ZmW6rsDIVV7Dj+cja1kC2lJVyRZzSn8lhkUq4L1C5hsD5Gc59A56X7A/z/ZKB
gOnZqNduDlxZBbb7783mW4GLVooE4DPE0aOo0KI8mAQMCQ36XfvS/yMD+b103vQV
`protect END_PROTECTED
