`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEBdBHzdAK7WNBnEKoXr4ApvVptTeF4CrI23k4/2GmNQ
C6izrO6C247lmNStCLnC1yEdVM9PzbWyulNrVI+a3sBXLoDTihES9RsluoUFAdR+
qKEX8E1Guaz9LXlXgUqP22X8eYIcJv9cHUmpgjIl+cn4YRF/30gYfaa77hwtlSQT
wfyey/ldgZxvznRipPZKMPwsUrKcCeIdUhmywrqrQcfMEbjvxo7xZdYE+hzCrFoP
pjAjwU7P7WFHANI+TeCrFW3CfKWgsslmzDR/VuFDyjL7myl8NqOaMUQ1I0aVTKRe
JjCXuqDWllHV7WxGlgfobHzvwxOMlmdNf8HCHcjX0LMN3+msRLDV2qF9RZ2dBp9X
tS3UmyfL6OAAVA4mW8SBJjIiYBqFinsnWP2iIhpQNogFF8WnzKlByMeIXK3cpu+f
7DKxRcyG5Jfn4avNH7a6vDtN54/JMlvrx05//E9KKAVCQV4ls5papgyoaqJ1LHY7
/GazrfK2BMrEBe1i9YdGMZMK+b4A+hTukvWOS4X6EtdX6SavDYLFA893Nax+IAWo
O30+V8q1FypKSU6E4oHrwTKloV2YwyDPi6QBQ6w0FQhbRCuYqRiGfWqhuWm2EcUX
3eKXyXWzcR9BmoTkPqhXb8bdZ6BSRMJ5kUsrhNntVPcShkUT7tTgH9S4rpcg1WIy
`protect END_PROTECTED
