`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
0ey6GqgavVAZYbeTDFfnhhRVsMACwhriONYJmwLMRAWCtUW9A329Uru0sXS8kqu2
qCOPETsVSpSK4VFqqpa/TpQCYu82V9JAYB/OZ92DNGUMxNXyS8PPgM+qYsPCC0kV
MP2OYbW9lCcXxGegInYCAuRmfZCClJUx60rh3PgDaZL2d/ECiXYX0gLNlOBKV2Sx
cWjh5EAaWzUCYcz/bMN+1IPjOI1H6b3uWg3KMZ/Gy0ghkE2n433L8y8z2atLMwf/
gnfwM1zx9t98wuy6mJ+R1YLRThryCW1Z4jDdQ1Z9l4o=
`protect END_PROTECTED
