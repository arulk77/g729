`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKG9DIxWH8m8aNTliS5M9Q10PpeWRnJpYbt4k6PvrctS
YkorqAcQKkauTiXkAGYFEhwfaH9ZJo2ahVdopXnT4aDNvGvc7Uutp523jvguOKwd
PqK7rHfZdnFnkA04lelbfYltrNtjYjreTgxAKsPQ2J38fRdtt1WGNo771zz31x/j
t7MgglOk4BaDllOhUp5bIsQk202TM35RsrFHTeL2bmc7lh0F2MQk6jbNj5r0JdXA
v1+zDvWxtkPed5COqVWvDcEIuVKT7wsS0pl8ntSPm/uroZE8b6WfqrGvn/4Nv7ha
ArMWBi3mHRBaFHHo63o8mw==
`protect END_PROTECTED
