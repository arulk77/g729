`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDGWVbH51jHRH5ldOD2vE1r9UvcOHUvp9Cm6kjMhxSEX
xweaSKUBuBa51zqZA6lAL7ScRk4DQtKHbp5piSHgNHeSI1KZrhnGm3CMLn8A0FaA
Rcq94UiYT0Q1f6YNEi0mRhJjjQFLv6ojy61/ggC0rScsb2Ed3Ri0jqRDWUTDK25Y
Lt1+PB7RhE9WXd/FYnTn4yCYJWMd4yPgXzVgf/wLydx0JxkxlcqfK1FeJTuWl1wk
odiQLwflpCSa0sKqEfb14aQtKwXg5yLD6wCG9hHZggJYEMaOSzcw28yIcWeCMuTC
hxpLILa1wDbQdLsml/REwr1uL4SyRtxqdIQKPvOGaFG9Oc8lvBW/mgBx+Tne5XOc
obT0GZEg2HkfFGsWSCEiVNRcgD6nJEE4VOhV/k6l2CzjKdwjzZJjQnctHjznykrt
3rabl/J6Jhfa24ECxab2gR/OXkH2cwryRVzlsa0b/0iC7FXbo6KgEfS4IVL+TQ8Y
QN1ASss4xmkQmRD5HEWzekYSh2Qqh3c95dLs2A2j5pyfeVQpxtIggEQnrzez/mWP
`protect END_PROTECTED
