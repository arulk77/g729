`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEukXWc6vQzfWMKQqnyES3YCf1swbepVFCAJOLdXTxox
XqmyPHE6fPUs6b5ChPzdDj2OGVEDaKzhkyIv/4p+bj1aR2kTeo1jyHPuIJSIh5j7
FrysntRa15fx20A5pRvS+IAM2e68dIBtyzeEt64ur/OWS3qVCgdBvyG6mrqK2M5/
YYbA0PAjiD69n18y/nRT3fqCxaeiCDANnfZJanWR9Ivc+p3f/osABYoTh4C678aK
nge//chVWtW1+DvBAmbUxD1kK4xLYv5ilLHIsxTniqiMrO6quEZaFAKUMOhdQIL1
weq/tIeHri4TS8mL0MNROVSRnPk4G7hRQrDpMqLd1m+l22HhOVKRJaDYps1+wiey
QeP0T83IYjhEiuFqjTtRrBamGtr2PNlNKFsS/u/CEa6zxDWtp4WdKca0u/Q9rQY/
Uaq0zEQF2DJOGASTbK29cw5oK1t85Qx54NMNV/odLmb7eN4//uc2UltCrRMoqXJ0
wA4jWiPNpUqE2FazIk7Xif602UGu3bubFt+8Xh5shHgNAC396kwYSjxcmgkciq1A
`protect END_PROTECTED
