`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKA9lgkGx4frN999/eQUX4IVVJhiiYkrU5oV/huH/WEE
kY2J5BP3Wlax95rYdu3+sZ4u5gSjPuGub09ho3MHddDDaU53Huovair+1c+JW8SA
rbum2qDi3Mq8uNUb7+4Djx4HEe9LhW/H/gbtdIqgyuO5UnZ5ZTuO9wJc+aI4t9iH
kUFZPP58q1w5gRfJYfiWb/UQ6KXqB0Qaw2qmsrId/Ohs4A1Mem7Upy5j3/kUep4G
QixIMFT47K355jo2hyfk11Ov8VkcDoVWzpA3D+2l0HE9bNDXwIA1+rdL4+MWA4qA
Gn16G4gN5eQBkCOPflXN/d/EnfdgcJXkcomlL8i3ToyMairGvELPiSAlgL7cJct1
A3mY2iicpo7hXTdOk+eoetsIVPGpx08f2kR5mYLEbz7O6Tc40oD4tVYzTCVNOwiM
9RSW2uqidTkKoCVh2pNgQB+RhNW9lhztw5SERZR6aw6cm2Ksqv92mnforJAyGW7G
Wq/1rXYydB1fiRaFHgf2P8zIVN4vNi9ULBH0KyO3dLqRoZgnEaE4UPLiz9+jTDRT
`protect END_PROTECTED
