`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHylVCmefoCnKIgTKcIDmBCVE7hFKkwTQMOKE+EWmliR
NhedoSI6rc2nHWvhwXX2L8AW/1IuPTDLGGhU26OALexBQ63GkRiBFqDAfCIsZqTW
NJceh5uIuiymkXVUbe1WO61LP4jlC0EOYrLs9nRtJ6LjKqR3E2KjpMPHSc5Jx8bh
jacDyk5AMmY/DzZ5qPHa+ZTuGQdXhRZISk6GOX51z7DpblWkgl7+F7QapJZ+eEgX
SAruoeuRTJSiTa/UiJNxdYWPwXKz5AHdTP++dxBjZQ/FHGoHag+LHzOc07Pf4xMi
CzbtqK1l7J5mfKPmKHuiLIM6KQ4xTe40EylU1IZxU23gvAPOijkeUgO1j2O74LJp
LLCNthQ0oGbMznySB48l34Rtgiq2e8jrVy8T5u7C5enKKfRLMu0qFvoazL0rkZNJ
PNXreIUbmnub4UphpQ1vERtmiHiCZmMyojPjI8803oIH9JMnI2Zbk+8VNvOAt0YU
gRH/ztgRldS6hJZ5/UYw4DhaTLtk/ZFwA8DbY5nsu7ux47yRKe+jhavWZAWHC7BU
wxYSz5u7XMiyASw21yOSuMWCSxbl532QyZ5f7NpYg0pqOA0DGxE3Q7/FO9PTjXW2
5zR2urvkMBsqPB5EPr8uhOpz7URTeMVOyY+HThhPEEbnrhyPoznnDM4pAoRmONee
`protect END_PROTECTED
