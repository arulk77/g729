`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49GUFS01ZMYj/INhOLRL13zJYJNchE1vUFmviPC9lKuQ
XKwyxP62SshQp9eB+4xzPM7WGHuDV+P7ODx1UQWGtRgCihRT3pp6VDsD96tOofl0
AagwCuZZ13aqvw1OQO4tz7xSBj3IBzhaj1RxkQke7XH+9+VhXZ07TU+CiPRD3UgK
MhmaxwCgFZa+hwWPOS0iFmGH1PdqsHdFZq+QIYHMgHY=
`protect END_PROTECTED
