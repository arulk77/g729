`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1accG9o1SXmCBMZvvt0WfJ5DmwGfVhmidvpa+Q+tkLtfE
HfEe8T6hfSMI5yR4l1957mLM+gBFZ+i9urz2Uixdb/WONN65ud93+I+KwtKxTAxJ
xzV86lX8Th2sR9LkTSdrfsu50FMk9g5/GPXRSZVzvMQayHcAcjGu97jKsgtQ4pF2
KTpObqRWAEuqRGy42nEwb5FBUSnCdykzChRAYGw07cwc5hKQniEHBl1xR6n1UCpG
gWSXX+MX3nsuSuD+wSoDChLpHxqAVlRT+Y0nqV7Ak3K+3wEY0hNZEY6txnWbxTV6
xe2SIhSGXhyp86LUzLhyUmnhZYGjegRYog7xZMKg54JiOdR/WU8tblLNwHc6+PMz
tBxazev2Lcb3rly8tuJMh9FWbN/fmcpVlbLtF3+1R40N9JAS6o11rZt5Gx7RnCOv
RAWIaWg7TR+oYq29QkP9Mp2suiXFJ/HOJkS/X7kDNCU12QOFnBsQbvdhX21R6WOm
uGAnuUiSka4wGNi5bYQkM7bUUUlVLDq+JWrUhh+39mrxGoPgEZ1BrmOJH3V+YVoH
hNH+azM1UV71HFJ1dxuCBVt0uJR9PPzKmyRSfJd35RbJNf9gzR2j4uEbk1B93t7E
HApBlDrnjJ0d6WLPmlg2u2tFBA2DAwvBR+HG45XfLssN2FBJ/5WY+wjIYfWfYTpc
qxmL1mqSU75WsM2rT/gLi0NgRkW9j47+dxtnwtC0DT1MlQluIyPsjBNdU9hK/xKl
rTtufvsTI7f/Uw3i2J2MWBE+pYWcb2nX3BTk7ClqociLEXvqPpWdf3bCi2DgKTCP
Jx1ayeB3TNK9T4ZdWb1pq03QuUw52LpHsBJu/MZqAWaQ/kjizyghkdb1PuTj0JGe
2cVNpTXSVQSIuKPUQeNyVKL3UlhLFSn34sQ8+8VsXgXvqWBzQYrFndxbryEYMQfK
zfjPxXnTuOt1XAeMVEX8bMF1b3MyDG0Fh7TjvGk7vBfdiUk/yrcaN9OofoaKxl4d
xWVhaqdjttlsLg9dVR+d/1MhCLVlKCIFdEUN3VlILVtdJ8b81CvCZcekQqW8P5Qg
erCHBeg8y02vsFpxm0EDbVk78ip/Avio9SLfm5tTrcNshgfK1ioXN97FDINtSYvi
PVAbDgi/qjiwvLQyWmwh9V7h2CuL3CzpxJ+xKnZ/XIrNuwnT+pP57OLFsko3cFSJ
FpZ17eZtG5xQAlhjV154gZ8kyyudvTJdB0VMh0rV8/1QmnmccXF6+0RurtWI/aif
1RB0I9LVKrlzedkhIrXMNab4qLxFUoUj0LI4fnZSMQJ58MqJuKwZtPhtUpCIS/z8
`protect END_PROTECTED
