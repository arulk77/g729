`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
klevsi5Up/DiMXdKlM5OWDQvk5qz7s70WqPgiKiafmX+nZWPkQHkDZBVZ0HpzcdA
UiE5Ko63DShq+fWSqj0JtVJN5Xad1W3lqqbqrjAqvQkhFAof3Uh9xawOcj2b8ONT
XyOU5I7LjvizVYLft8YTMq5LauhJvFC2noRzyeDBRsTxVxOZLxrn2P5nX54m9jkc
jfQY8b1owaryy/PAsW27GH3mM7fCZi2o1+m+3pWR9Z+v4o7wfCd/FdUNjzjkunHM
CopeYZowoReZ4eScZhV0WVVPu8/k+WmGFq01hnElmywH/kyCPxRlWFSoMo0usXt+
7M+7otoy074in2Db2bA1jg55AikGbARa+C9wil4Yn9tZ6uqB/wc3DH23uxVkd6Ia
HrV2e9tdepRrSfe3LIv631p9yfp4b/kX7xRJNJ5vCnvceBt9lPcbSLx+l7rqoqDJ
QmiMv7ZmjbitAeqzjzezm2yPLcmIuX8vtzRWurexJifW6/M9jq+M/E+55xgNAC4q
kMGJ95oMrsLdnoCAr/IrVR17k5c1gU4LWvDu4iLy6vwe00qcwLpcnDO5y7lKAsr0
sN3r7fudHKjRJ00Dl80jAQ==
`protect END_PROTECTED
