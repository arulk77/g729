`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHcAGZmHxpWZPV6teXF/XsbYar65TN1a16XJBlbo9Rwx
osZ9nc2Pz2ILwEjaA21LsWm56T+mTTeo+cUPFYTrObzqAnfFTcmKOr9yKiCJuLTN
rJJXNZu7kSJUo6Pwsj12dfDvE5IdLXXJXZC5ffWgyh3+BrYwBsaahUdlXu7c432u
HogfVAf/f97jyXBUczY4vQ==
`protect END_PROTECTED
