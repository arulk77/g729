`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zw6MsRVCcdtE+bqLGpIGb7mRF3NvmcQ7TEqm7O0YOaF
W2xoOI0+HOd8b65ML+cLf3akTDlaDQOnhPF2PZoVucgezzqPm/hd+Jt8S4jFRK57
0nd66hO0JgUOBLn9DqWWEDteA8GLgUCGMjMHPrag6qmHzraHbN6IY+HQWqwKASrd
1jO17bUPYRu/I38uMYRG63V3HFXO4tTw+dWVtFUkXpglbNUS4TOVt5h6QU1jAynd
jrbkPT8kKzZBNpY9VpBOcR3nA1+5jlqasbpWki9mfvdgVMPAMTZBOJiZIBtz7UjR
fqVAEEkEwr5K6fZjGJMxgA==
`protect END_PROTECTED
