`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNo6LBew1xG7uqsmRxg5nWg7HEyxhRtc8kS4Wfix50TZ
Fa/UnMUEpe8fuVcuu6vdUaixtb2KGLVEMmpLMpO24/MynCe5FLCaCC9YgVKSGEU5
JebuuJCpyOvB0N+IVELxfHjWzf+mjKA351bE8rhb4wuv0i8vi7g6fvtZt1+SDPA3
P1sS06tzzaHK/qr2FDhzGOWO4vhXIpCJR6apgSo9fLHZ+XML3RaJG7vVRTij2uBI
jLbp9d4RYVOu+2qa0K+QFIm9rlmoolQyHGiq2cXCW7c9s1mp1NHTQFEW9a5rdxzP
c0wIhB26EhccMFnnfW/d6NVn1w7cUGEXol4CAVFfndeB6PXjZmfliZjKGNk7NtTg
`protect END_PROTECTED
