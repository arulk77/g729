`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+DtLVidmqyA99DrwDtjuczYb68cVpGSJ2LksSbInC9V
cnTMxT6mbImWW5vWML+/8dH8eDWz0K9XZJLVKm8CDRDLA9LtjD1k6xMsRZTec4GE
evUFcQ3hzH+uSkIv1PgL7RCzBQ7QLy4MVlnbvec0DNyCZJcprILgcKXDH+9ZTqye
3FBUFuFMUPeHh3SpjOjf5zOMg3wbADbfInQNb9u7ZOdImbPvahUADJ9E9brYDnZh
053qF6NOd2JAWQeupXufgny3dCZFB8WLIcVG2AlvG6B87c7YGEInrtnBYKR2Fq65
YzEjh3ByyApgT4+3QogqPdXNWzifzUfcx93getrafnGCyA0mJ8RIVEwZiQfdkQ84
v6diEaT0Gpwr3aYbDEFo3/ikFUpExsLZ7zPITBBzmFinIZTbbboSqEg3giJdKFqA
tXsGJZdz6WMYxGA+kG46n2Da9qPGCSg053E7m+mXNkURWe0Zn8dnZ3mf4R2AS6gG
utZlE9NaivhraBMwx5Bg8VninnTXN80TbwtsziRQWg5Q0Z6sN8NIe6ihFd2OD9mH
uLhKjjRlVmvMsRz1Dz+kpmnERjCbXbc6bMyYkwiY7gVYzBCFCdz8f0WYeDlZGZHC
akQA2SVhPFa81DQtc1irKAZJLqYpCoLUUwt1M9lKRlTF27PkRbU9c/UbBK2aEfh1
`protect END_PROTECTED
