`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2EBoZu9tBf8wFLCnm6xiM9TEV3ui9TR6mG0WNXVJ0x6ft5wycXnJUMG7cr3VRBVd
cqKKI1tZB9oPRiD90MMDedRDacAJYSh0X+ik2CclHbJLtx8jrCW79Mypcl2HlcLa
ZAE0ycoGzayNIWqCJgOkCIgk612w8fSLVVQqGAQ9mSd5UhSEd2xc3HF/JPbH0aYJ
OYXvdofA8VvA2Eh/fXoqBA==
`protect END_PROTECTED
