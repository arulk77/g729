`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2D4LnyRJ5Vm5ZoX8N6+meBp7s+FGIwzlyZJRPNNWIQ/LugtoIv6odFxllTp2xzuO
a8AZ81PZUMH8Us5TeT7o+FaDz4lGRFYlbSFbAvilacyM7rR3AH2j8zndL8LERXvW
4/BbntQrjUE9arAuRYahRTBqJBYCJhmfWIYyEXA6fbprO5jb3dguqjyIos75tkZb
`protect END_PROTECTED
