`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
o82Uu3CDYqlkdaJdgdOZcUX4CuK87SeOdyy5DxQkb6ebE931+bp3KBeuty9CsLyu
P/aaDNj0akIAgV3kXp8BlF0jQb0vfakyKkQ5muAJCHmdolcTyATRc/1A7939HnBN
FojXJ0Vj/JEjyfMov2ZBkY7/yV9wL3bzTuUxtQDh+qxEtQjUF2vWOrwPXgnD2/fa
guy8RU9aRBfG+UcS0V6xVkf5mFTZIgIfpr4/CXMXQ+Qn/yZE3j40eEXg+IQUiIkR
NIDeSX2p8bDeazG+xha1zGAZADvuS9vJISUY4SSxjgM=
`protect END_PROTECTED
