`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHRS45iAjBCJAjSm2D/VdBj2uqFCG24rZy9WI95erZQD
rdeDGYquE59d3xiTOxcVfmaqIpcmT38HA/ZvXYi47eA5ZfzDGRTnUBtQuXi4CQKW
O+7ZhJHKEWww5NqzH0519JjORgWNmwzIdD+gygzyIdkfVbQt2Asdw4hXgpNr2vL6
MrkonjJXjKqxf0ksdrOctDGPlXLbr/cDVSzz3whDckea12RM++WTPEiND6H0u8F7
wIPCuFALt+W6OEj7FXICtf2W3LQ9UyODY1iN6PmVrXRtSrTs79s5MAptqUSSLBgH
bJ3+QIiWZh+Gp9gNTrlt1967Hi1seDXS1dtJaRvSJ66rknHiqYxQx2h0o3VNjguR
iOpqWleO/7+CPzWLqOD11sFTuyNvajep5QexCsT9Dq/h7o+bFcDWjrJmleJrBKxH
EJgwSWN+3uhHVt8fhB09DLJbZcG4GfOfxADwDzqIUSP1NXBSp3syKtO2Zg8TEEvH
+BTT4JzwTUhOW/Gw4Fh+96RqG0cc3kQnk747NicUpWCncUS12fcYUCRnpjnIY1/F
hI4bYNbUSneeHFWZxJ5zJ4KRz5Jsl/Sc5yiqtU2hlnpHFeiXI+JRwZ6TeGnJnGCt
w3BYGKlfmJBXrXpQjTNoHWe2rS503SYfXOVqFzaJGU86WTF7G1RbHsX8D2P1mCCh
B84iD6bELOloKv0A+SNSfmZYUTj3pImFmfd2HFfvdvphUezMFHpPQLr+I9W6KNut
M6+Yx2yeupgMJ3HA4BgIcSqWrb3dcus2i2UoShalRZlmhTEVfititOuIME+XJuLy
`protect END_PROTECTED
