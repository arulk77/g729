`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKAj5Jx3fc6S/9UUVrb/OtVZ08QQEAJ/kfqKxaX8GRhh
KXX/ofVDHDUZC18BkGw3+oHlr3b0BtpBBj2hu8FtXtRbOdHan5BqGTyq2Jr8TKkD
F9i/33zdGUwHtFo1Yqve9Vj4ihTW0v6ud6g1s2kMeWz/I/YAGGvXYf4gv2bm4fWg
wn/YLb8/TXWD+rDfVI0YtyXAuI2yfJgRbhd44Dqz8N68x047vMIeFnwgWpYDdpKd
BMMvGgyVnChBO9YkER5sNVJp0ojs9XvGpwEDjQefACCU8biWYBQFQSHWDHrISUUi
WWLHduAAzKRCduYEGTM8Waycq2WZt2YwoFRkQQ+YJYIWnRsLF1zIw/zhZTIZLwTD
`protect END_PROTECTED
