`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
76sFkWaWtW2g4TUTKwVVqvL9/Z6QX9BnlWoNoZWDE4pLqaPtttrg+KItwUNJYVpC
yGd4IbGryn4lM3/VVcFHBjsyHrncqTdHByp9oPixecPo+gL1Z1fPTDCB4GkVw6/4
G57tVYI1kd1oXNPmcgKOzS9fBggn1T40Jf1CV2bGXknMkxbOBaCnoA+VEhxlNYct
JwHqMbcwMQw1Kn0fzTN4m7A8CN6S38ehf9/50feKwUruaiLFw0FQPn7+z1KrD7ld
t1AqkVZ2DtRYGH2DN3aoKX/UGKA36DUg2U/g+kmerXbP4cNc8ZX7dv+cgi4/SocL
`protect END_PROTECTED
