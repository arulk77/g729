`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mNbLYbR9OPpDYhPuqsyWLy4Jy1HZjKOB6ljO7WarwCm9yAsgFOguaiXYZrEdJaXc
mmE9s0BYZDbLmM26AOD7ZrMVXov1OQn9JTRwJakngF7yMkqJFxO/3q0XJpaQjPID
xNhtFz3dD2kLVsiKqZcBYsx+Jdhg6RZsp62zEGyt90/itXKcQhFsVLNiKqJVNdrR
8Uk3zQgtKJRiLviBXcAu27hs5Qc1UExTbzk4wi3Ni5JoNTiM1dgcLAG4/K8ZFEC2
Xr6obLhYHNgYelgH3pXCaLsPNzvQbVvpy+nCTuqtwbc=
`protect END_PROTECTED
