`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKGkVa+tP8V8mjLYUFitjptCSBO5b1EZm47laGLQHqRO
W7wAkricRHHTJcgS5C8fm1dBFFjR3rGBbc5JeOS9C4ulY1C7aczAvX8Hvgfl3erH
UmchABk6ORv1px3grS0l/NqGq2yFfgyidErYqMzBdXMom1QEdXdWaVvjSVidkjIz
DXsnTg6Mn2WB7ny7MbRE4/4efxrfALVh8qxBG8bq1ple32EB3a4DpIxs2p00kual
EkPN513iQxi4+I5IsMJgTZRhTIpWc02D13+qUxdBJQfn7mA+y16UwAYteTd+B9XC
a31n2g0EGJA3U7Z0R0fjU6RJjHSSMBixzN78++Hw93mb09ZK+TIjJwhwBKMxBhhD
eq8Tc3PLeCq692HmuKw4Zk+22Z9abstlP0OP/SoyN1SBjJ7lOJ57RghhUzgDulzu
l+gqxilK1nE8G5GhP4zTwcFvZ5k6uj0YyLTrPF4N7ZHj3vCB01VQzaKUQLBKPQeN
BzLt+pSfLMM8h9P1xdlWWg==
`protect END_PROTECTED
