`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBzb7off0UFVhW+wEq0O/tQwvpnAq6l/3NuJs12Ziady
EiEspWgdHysb5QZGMS07jx6rx05EgC9nffOhIb/z4xQvpr4Mc1Jh5A2ThJPJbmLZ
FOghLvDi6OISZGkdH9wyTQUpGFHptyBHIpZL3tU5p0a8Msp0krYMrMHao7APVVp8
lkMFhq3AdxB3LhXeI/7t4g==
`protect END_PROTECTED
