`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAVRFnE/JbteffOI0q+WdjRq62ih177C87kPUxclt1uf
JkCiZPiHtJFYCixNxILEHfgc8yg9WClfPbsck7zvMufBREUSQPheMUSzkHpSdv1N
IpPLWE1pc5WFlrKDncu7/wHxBOPsANUaH6sMd4tfeEV8j27j6eM/KvvpiK2bf+Sx
tCzNqcwOyvQZDtHmkILDd4tPnn3NpM0SeiBWKUrz99ciBCsN98kFe6X2RrIVaNcs
OotV11asd/tr0+pz6vvBnvtkGMj4R6Y39IRbI9TEN76LfxgaS9zNkcz2zuknfaZT
BapBRV3yx3oktbX9mNkikkcG+H+nLf3xy8xku60hoHS2y/EKcJbaPoPmCIJJEvV7
`protect END_PROTECTED
