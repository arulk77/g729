`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNwK5Vms0A7QwzrL8LGheiMHPNwUH92zpJPul5uE5lS+O
1DVt8D/UGl56CP58DT9G7ghM4KtxZD0GTpw5vvuWP+BGXqBVAF5gO0AZNb4AGSrJ
UbLiISPy284dkn4ttKmBFZ7MMpmmSh67hY/ZHS9R6V8Qam6APyURBNtJJZ09FhMs
CtNu3DT0eBpUBmV1FYTvjt5H0KAE1BxgOyVlu+pe+nnRff5A/SYQ1wEo/wAbJNS/
eKBLyrZtDc/ia3SzQic5IxV1/Gw4vAqhnzxon+eRSp0O/2/xIxQaeCcUYMeajRoV
9tQ/u+kc4S6i6etDNSyCSGLjqF3IFp/eOQQlJllpsGu3P09754qszK2EK2P9WBuY
lyugX93O8y+GBGa5BpjVDv1ovEcmE4CVlNWmxcsx0N6fRrGs6F024MF8MhINrJzw
MoWazgsSIRhWSw4ZjP89Qdczy/l4jsMP/Ser2YLxuZoXdlxjt2onu9o24p84Rbqp
nCJehM82EOPUmB1wnlwhz8FJgEV9YzeqaamhmQJAjme+NeZHeJtsKtlv3V3tka20
E8ICXtJAo6H/KzfRVk6JeMr/GodqU61BWEVCxZwsr9NK3cR0HcTUJSua8o0KDtOR
BQaqdXGgG2o9+YtH5yWIprg3/gorGhR1M2B5QBZNcwUTFK169ROe7d2nAxdBNGRR
O/s20enTi9irq9Zzi4HFQPEIWcjO2czwCd9HS2Pw8CXyqO/NVcGr5IKfT0NR8YVd
joVTsb2DMHFxRHeFRt9IpT2Xzm2QUeh7OnqVXp6J+LSxC5hclZs6ARzQhTHWJAhq
gKYisTXGotQisk+mIOjUZ/IZ+yjibdyHbgPqCvxBR9bGxLWEiPH5R65tdCgC6jmF
xC+yVnFRBXzY4VmcpEQfTO+ud0guqKWzuekyD8uvf62w0J3iodptMfavh18VBZJD
VjPbb/8SqMBEbEbLXqoVMrkJc5Uhi2Y8G0ECLePSqS7ZWv2zG0q3T30TUWsfVLTZ
BvQ7gHPJ+ENHPeGD/WSUjMB4deR39uU6Lk/umRlaXCy1IrURCO/rG2UMYfbg2Djz
9uNq2nmzqktdKYFyXaioZxqSFU8CVB4f2sVGPZFPyrnJfQqyJ1OZlvZ4+pnVhE4i
Dt97qQcjQ70iVg5TNHJXLfInbMQlE6M6i7+BVwTpOpz8OZU6wQjCvxD9WdZaGXch
jcP4pcgyHNcVICTuTty4sYRV9EXwwJBx4Zl59wmloRpRKgie+cvjhQLrhT8XUWmg
zG+Sp4l2WN52tAr8QTM8mV0LGreV0NCcp0hKsmlolDEif3DP708RIEcXiY7wxsQ9
wGb9ISPaIDlbm9x3aICv8f9Uy9uNR9rWEaJBOiWHfmX+ewyIPVA36eLVlPDh8jte
+D2hFLhc1HzXf/+NXwA9P24smI4jioqC4PmtQJ5ZyaUYl4VruLq/aDuPc87/dKAi
lUcBlnqIz0Fp6BDXzmpKBxyNJqjg5MtpFrHePSKqDalJZPnNMHqRcwaHjyXP2KPd
WK2qudjK0tp1trt7ypKUq8XE+ykTwF0Ef+uc52t4v1BZCDSy+uFMsIGEw6RksFjz
JP27Gq46IOQTi0eknI10if2XR9C/3/nMtTqp82FT2h5uokiTpJnvi2629PP+lXWM
E/+WU3NUfCtVg9OtieW1oq85Oy/z2yFl0+uTmieV1LWpoviqJhl4ueQD8RhzQbo+
OM2SHkHkl5ioRtQro9fk5TamOa7pStqDfukhQU1ezVqpsFDONNECUIGl+MzDbqyf
eVmf8U1feGTg0+IjqFB43f7a6PTK5LdOrm5F3ef7bXDeevaJcT+R92+Sda1bgtPF
QsH5Bw+z88sjtrqFg4EwCgG091Xph3m8O04PdyLLjZnUEZmYpSbdeKWi3E+8eEN6
kplq2Mgqy0JXfJenro+ZiNrR0apcGrjy8WMOLm0/i3LIEj7Tod7ZDQN5uYvyP45H
+4mINk4wincl4F6y3+I3W4FaIx/qy9isEm+9xMS/uIV/Kf7t8Gv3cvmuketLLpRB
GSe/BIPqmUqy4Mli7klEn0RVMoRR7MSxZ1PjO3FqUUFR+gJu5nsv+Q+YHYrP0GYh
m6gZxq1IzxOipRmcFpGnT0iksT/3RO1m34JUoJXVyzJY1HP12OC/b8MJTxTkiiC6
r76AO886cJYn0phlxamWpwjMAiidlq69FhAVWVIKxdPF/nEsYwmxZ74XK/8Ug5yZ
RziuEShg5ZqOVGVJwQ/x+0fv+u9oWjIiZTt4FiOVu+kFerRDiKAMvXhrIJym9go0
Netb8zsVi0cuQYcm5F6kEYraTG6mG9SO1gbSB4b10ddlAi8vcBtG2cBbYwOzErW2
L34BZJVtazzCMskEoguvcMv7lnTje0g5iEQmxF+2cUbVGUfKSBvxzJRYJfuGY/GT
hTfZeDN+tIMhtTdLpdEZU57jhe7WgX67YjSyXe3GaUz/vwlrONH30XrezCZePjAb
z4+Y1yFg/ykUBGXh95szcD2tnUWAZYVApaDjBG+mwkE8dmLgA+9oKr02GBPSWBre
9eMDs2UGdBw7Um5CrFavSWshubobhCzlNSN0pNr2i2O+AJisRjsJ0H4XvnDnTAcs
`protect END_PROTECTED
