`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ClJJaVQDBugUzEDzyA5YFuBLlgDkDgz4s6cco53zqlxrLlpvovmgzXB/cJVtknPn
xuZ4QH6+9PSTXoLsdXI7nlazYf4+wSTnQPk6WGC5PP45BgNI37m1tDWtlCh8y+hU
3sQMGb7+5NdEjS/hkLNHfvesAMbx+uxjc9nAL9qAmaYa1uEmx+oZOl1fGmQGxMlw
3WkP4fEatZhT56cyac/PvW1C7s5u5kdggpJtisDbg5emzV79IVYFwq5QnEHVKqHw
uS+YIvnvCObm8vn3JVVy19JNz7hYwjQ+D4yEhrq4Gt+RrbCYc5mMeGxxi/5y4tiO
MsOhiLusDDBFjhIfiC67wEXFHb/KfavHcF59Klz5OkgsDiWKLOZEGs7mc/+h7gUp
Nw6y8uF7Zf/+B6JhD6sLYWXNYRH3ckseeQH2ZJFlV2WcPd/XaFetN6X1DIcqsuRA
gGAK0xg1GMCUAQqqE+/9L5glrNvdUdO7eKmrQ1ILZBhUuiO2m1KyHrXJSjJE4EK4
+Q/o9RFwbzYAQ4ywjcxRVg7mmETgvLK3tOD/npegDTrp/bh3/SR4bfl61ZSB85Gn
nPl57pAl8hPmTJkyTk6goqiyLKsgI0e+nizckxfuwwNLbWOQKEKONIoxoyMhSH0z
45Li+EJJkbBOJkXuzo2eS6e5xH2EH10BjQ0SK3/nYj1SU2c0vOlg+NUAcVWykgFH
Jioa9iuLmC1t6wiiMjVD9JbAsxti0Ly14gKyOaSxum29vVZRgcYKPUvvc/BXYwdE
o//AZT8GNGReSLUFsjG8zzSg5cHY7wXfcHqMVbCfWj1z3woLnCtQrH4C8DOU9fj0
D3r7ZxxK+Tm/Hjz3psZkCs7Q35LLbrOCG89iWJ7DjCpht+gLM9XCqtCDQUR5fonw
KjuHZSMv6O2vtwfBSeEvem8zCATysRclSSJv/MIgEZ1lLMpTLNdIRRUONvKrQuqK
gXGwQvaZrlwtr9Xn5mmO1EgOcm+mxH5je1PtvZCWDZl9JRnwK+QDH55ETZbyZbjs
h9s3JZOboLKnV25dzInvBqLlMfMVF9cF3VbWS9Sd0Ypt34rf/D8jj/3AJ+7go7pP
XG4/gjPHhDhO60Z11jy7zJlHKmKlhv9mMaPq7izMF4xeYl0nZsgJxEkMrj1Nqnon
MBl8vGdVxV+8B4SYnbbSJYIZTH5gnqirN9bM2Ew9vcfzzYCDEs8HMZwXavQUQ1Zn
wj++EmhgT98aLhjSqlpiwsYuAbRZ1KKMf2gBJ08ACxYwqOv4Cs0ODp7itwfmq1dX
aJ9JXw0nHFG6kudEFJM9uK03MtsqZK0x+qgZOLiXAqYZr+O+9OpR/U9xeLbHMJBL
gloKJckjNkxUKjB0NhnOKQfa5YbMRaLH5gGWN4wGBBAlhbjdgSa2hmplTmYEpix1
ECvPZndq0hyRkvdhwS/7++Fp6Nq5TjS+VrRZfg4HxhBLkXGVyHvy5LxmhEI3oxWx
FPSjjEtiqDBYoo/wfVWGmUNzmEM9E5Sbsw0usG6mtJlpoATxHMLvw8uC+1zP14Hb
Nl4N4ExJ0gxyWiNmRskDXKpmvmJkvlRBJ53EZ0K/gh8V1/JUSD4lmQIgdp62WT36
3dqKTGU0pYFar2FwAiMan++fUhuu07sCedR/cbQUU5nQj2j0i0vU6kx8YpYQRfYw
CEOVHvRtFiHwze7IbcYh/RclTLMyEFg0SXA2YeKD5Nuk+IWPCJfHH8S4eXXxbNBX
Kz4Tl6qwL6JYnwOWjs0s9XO6iUGBCFL+dVfWxkCbHaMZXshnafyFAhceVhqWI6SF
Dkb1VL4yBbid2xlOscPsiGMTAMDV8Hp4M375GByJUdaXd2+/uRexZ9p1p5v00+VA
EUwHroguAho1NqyipLrQZVlRRFz8yJZ9OyJOYZA2w60Y5reCsH6D4pqfOaD2ibli
GstKlKiAQpZ6IwQOA/B9ZMT+UcN8UrInM/NZkcv5pbDHtQ/KQlLAez/tWvwT6pO2
zhp8H2cmJEw2bYaJZMHvjn3W3mAk+rhIg0AxUc3shR5+r7MTVfS9Xdhvi7OuOeZS
rt/stAm8WAPYwDrExBa7jJkIqFo8EKgiaTuyIZSVE9Rr7QIhLVJhwOVY9ST2ih5c
3trHAYxzN+2DRYJDC61Zgrjg5990vP2HykA12ptf2nmLtYcNgDsioEhbGsTWba5S
H6lpUgPblJ8U2ZCmz7aKdSqLQUw5mkWxhG+KW9QDNW60yYN7J5EYeI5ZG9T5JCEm
ZfXHCzDOlVLzCMi6FO+RzmLRg9zLErLZog3ivHMMVOfzfXrzaHpcWKqXpXIOyFrP
/Wp7oglMwoH4BF+6BnpklHk6Uxz8erQ6oj5hvIYcds6j7zIqCQDONxhVTpYJXigL
JvPXZRihes4Qa5G52S5muZR7c2K0XLGx1+QhX2lNvRS3ONX9UtqVOuwdngvzpNjZ
SDdq7Ef4AJMwppHmqVA/WtlJE0FehtJnvGEmi7888afQkVTyHC4HKiJF2uXm0DKz
NW5XM1ks9KcS40Uhbj7TzPrZKDYyfHWUp0aW1fFZcQ7iCX55fm2ZNEzEmcvwom7O
xT3mtsDpmkvZpcOR4KR4fkU9nDfI5FQKt094GNuY8R6S94dODDWfqDQ1QQlYSM0i
xtxLO252idFybfUfHp6BCl4nBO5mfGCpvyop8424zgWRbraAKhnga3J4dLnEI/qR
fodnAVTAkK4A8X19ItCsGJOtGrkiZTLbrPtmXPOT3mUok3XNjmNnpe6XNyJdknom
dtX121sfZDJ5Kzb9CwqpgIdFsL+kKZRfeguhpnQ5UGTW73aR+te1Maya3Bc+pzOX
C19V7+/CMYV7umjGBgn0hCMBEvOLkuUe+Rv7WinaE8sYOpClz6/6rcF3ynRQD7EQ
606BwFepdsVEmRcZBqhCbFRyXzoA5R9P0xWo1PKX2Ja6NfBKAL/7QkfczMByFS6f
BhzaUefj68p0kpByJEBzA9wLClFisbxilH4ToZlUa+G2ugDwJ7BEtnThGfJIKd1F
dVi9KbxiddFMu/pMJ6RS3q3K1t58jEdzgI1HFh1YxQAMV/n2YBIf5mfiedl/0RuP
r0IYBNCCnOaBij1S+/9hYQ66kakWyPCUZT/QFqVDwXebucgqtZzNGtFS/bbeizrz
M9/SGaslq014+d6M6t4j9rj0CXRhGwCFTHiowNf63WCv03le83PUIwQOgXi3wHQv
0rS1i4l+5R060eA2KnPXocdstX7V/5O/SoncmNkRA70B/jZJrbVJo3nHp6KxgiJt
VrgR3cqWiHF+NPZSOZCbvOhV1G/wJ16lIwO567lUjzDg5m74gmSyVZz2qh2H/9Sk
MGgOsYMTUNu2vfuG/mUf7+ZTVoEs15LIjGRPNV5vIMz45JCBSjy7hCLf4u5zJdmZ
iAp/BiH/uMNKzNep33PQA0RDZ5ziC+vYbywLF9rFm9L16TEHFU8T7TyUKWZMEYbC
EczkEmt/ymFtT221bapTVNl5lfU20b5JnCx3GC2R2w0wkHRyLQCVNqQ5mBM/FKZ+
ixrRSaTif+j4BCr+zktM4cO0F4812fORI1l6apA5RH0JcXt9KR8xN5v1B9uWi5l9
mMgSphwxdDRHvLrkHxGAdoOLiupLHBjCboDfrWH7fmf1Z6tpg/DeYWByfS5PA6vn
DJ2T3D1/zJRjOHKi3bxjmfa+6+WuWoexsoTjSSeqCCCeRt2tgJGNizrMJsytX4AN
xipBsO/NhEjfOP6gD29E1BTLcPx+gKtmdb0dNs7AmqdptOPzJjp+EuUVcORfFN+a
hkMc4bwst9DNMZ989tgBTzDcwcj5L+5ZfxQPxwkIQTPvU8sY0ONVbp8pTg7W252l
btFpMxkFLD7WPTszkoxHT2mqcGKycDnkRZz5sr1u5RjmmW4Wyfmh+YSV3C0h68Gr
llsHtcqD4EUUT7Sg/qj7BZIg+1TBbeCm0z9dvy0xCbH1dSFQhy3deaB+aTYPjVWU
KbaGWeR+iCZ1VIW6PL6kmoVFrcK0oWqIkU/9ILiHSXfjqiiBV2uj9D456mIHULg1
Gi6nZCAanloCzi6jRzAcYBdbPERTm8SUijo+zKtyw5KCDAEYRhsZKUdDBJnazDs3
kBEManAm/foFYyQ/k9bv8fylVUFkt9WV6M6BeeZqCuF6W0nwbqnirM/KVaWaXhoo
wgHMqvYTzwoA7CAZAYQf2qSMXgwXYL+R6Wq00WnBzqKTjfMb1ld6FIrYzzK5/Cs5
Ya8H9/aM8SJ3X7ZhhU6W68ankFDgAeMAzgvT6HEzqyIEuxRdGnPKfEiXodvPMw0M
ulZ1VU0nW4y0yTruSAQMD9miFE/U4ojwkBAPSg8wl1B+uELC/HD5LUUBb72nfQWZ
e31pyyYAi4W9CP9IQNBFm3HHLKXse4NDQpjdBs3a8v/DDMHbUDH1e+SnLOGwZMLo
eZOHh9Qo1JE3l4T6kSZOckb18G6JcT+7VGR4l1dT9wiaDEssuy7No+xnYyjPsOrF
mHdpcx0XwqwORkUgGUBFYNnH5447FX/8kRTHEfourpeg4s/4J9+MyVhl7LsBvyvd
hcH0G1ClVJ0JL39LuizQN8Q6U7FFD/unMVE1VeHeljgXgdN/eyqYTRpsDHc6cmtI
vDnt6EW7bXCp8b8lmlrsXFE33rYnNfMmBAJ2wGE8FG/vy6OUBs0ZzFqUJ2nITXcr
ZTdKJ7Wlul3AuqDcSLVvhCiXdepNx024zzNkgvj/sBRj5/JFECc34e5COE3dT2Sr
P+aHKHrGWiG/dJl5ZWlUuAdw8R0pr4Ha6xXHAqJEMNWRzRsxecHCPzhDJmSavkUU
EGnLHpxeeDyJEVXOAxtbof8jXrNhOOnsP5tdAAKyUduqXNRFgP9yjQE5/YUBOlYd
GrTyAlkvxoHSYHvXIY2PDzZNDs1VT3e3l/eKLrGFsPRFy+UkbVY+O+tJQOc+bIrD
3UUQrhwMZ9qppAHDAA7JdbGpTkeLcuhyoJldKDnHcDCMXFmTI0eC3w4J/BueJjud
okdVtEKn6/4h7Ntk4KJ22yIbHZiLhk/1akqQZo0s/ShM36d4oEDgdNuviaJVgNyF
lJE+flm3iA7rxvUZ1YUcyFDl2oJZXboAh4DLSCySKTxnUC083iCeLiCq3Gvmc4E1
fY1RwlJtBVP4gwqB5w+7v1ejclrPcS99+1H2xaZTyFQeb4WC9vMIlGdORZoKhe05
w1ryQZGVtK/5KZeWE8Ffks6Y59bvCEZ1mZEV/LF6QYz3zM1J3sqI+c+UCIVn6OpX
uVcuFkrnUBs5K8pPorSzZAc+arOzHocriX9RfwTUyYxZgWRkiaRFS6pK84cWQtuV
fGydPzS9uhyW7XKLO/SHZFFFUTNgQznB404HbvorZozwIZT2LzcgXkQJfmNi0d70
iEK8VC4Tb7kVIv4tpw975pAqOU5UJLUK+SjcUhNPUtGJm3EkmpScA0pJp3taqqZ0
2gKB9HUgqTYwg9PxRgz0CPrBjtysRxMi0JYFXQUThrW+xPThLVuZxi4MX6FaUQBg
+MsBsrwIiLKa2PfABUOe6qUfmrJwaNlsch9McZ8ldHs1GvjNf1Gn15JVRSYnSsLa
UGWDn9J9g8xEa6gCHcrxVNCk/bwKPshKaVcxdQlN7KRn6HIhWFp456RvzY6tMMuC
FljTH4y3cu9mUFjh49Kfzq17QkashQ/ncl/SVIEgHxjQsKD+fYk+uYGg5UrlZRDm
Ct5ybz6dPXJODaaGbgUfJGMUp6+LbGFfpH5aY27FpQKv3THCkPhM24/vmtuuNTf5
Wj6PDY0FDhFLqu5oXHUfgbeJlTyGFmcpGrnsNFjEXibTu49SMwAbZ7v5YxBYdJHG
wQWkud/Ksw+2gfldMTwNZpJYh5Ws1I7IVBZCfKL/kfR81EtdC2eJlUlID1fCvGM9
UiArc4X0WQMSfcECMvgB+rIHH+T5L7bl+jSDsjHcdnh9fsrNIcThkwJXDNyJw+Dj
ebnLyPthv9MX1GHOmqXAuv8rG7dUoLamrJv6LdMQQSNmIiNsCfVYGgdP5EgQ2TUX
De/quRlYGoqq5SFg/gzTz8cN53Z84hzIzW1YOuyQjFyfdWa2mCmyAGVyKHsUZc2X
jK474wwmh6P0phEPqBFLaSADAz0Xy4e7dnOmb/ZHPwxSy6VIkxqkLfgSlYWqy+sF
k6kVFplOPZJptBLvpVmFVj8iTDr2X3EKF/dkUFvo6VftELgDVxYX6ow+KmKaVUFV
3IOzwTvMHhTsmmuYd4Gsqg9BRWkfV/BKyAJt54KRvnZhS5XFm1g1un/3i437ubIj
nTliQd0jyOloCQxKvrMg5RCYSQY/FmhNDPx93I/pwq3z23AdQCyYcWdLr/oQH9vG
Iduwqog4nahXG+uNLeQ1pxut6Pb7odM/FkYXMlAmmn27m8frhG3hcdAfo85t+KPN
BFKyebB0sGCi84ZPxTueXz+l58h5Lv+Z1LYw0nN2IjVRY5nc2+p9yBlZm36xVeIZ
WmimhdwLFgIs4q+gKAiuTj9neAqvgJPEHe64ibHiCABg6Q9J4ZhKp0I/WxZSgVj+
hw+k4HjXe1LcdPI0PjK8s9UTJZi75Bq3oiZHBv4VqqS5DktIjf8Z7YhhU5oFIWKK
4V2azYQnvk2JJNrdX1GY8cCOlEP7Ef4fn+dumh9uOwkmdsJ9//5FeZYobH075YI4
rCpE3nRANDc5CSC3efkNcv8kIYeOd/BV1xS/GsF5Om4h+1WOfskjiMRYOFMzVqNb
NTkOeVvNMlc8lb84OPpce8c0WattLQmp7PxGShzHKoiDYHOrN2a/Q4v9s8tq4BgE
q/ZsUV9S5RN1L8h9nQTw7vlJ5r2Jw2tfg6JBdqso3AmwXXSL6N44flYvyiVOKjzD
EVnFrk4C6JbTYWBbO5PjLByh6U0rTuZKw2RS52HQD2v4wEu333dr7urL08ivf3Ss
uOYpFLYP6jCPWjl7+GS/O6tA72X+RKG1IGpCo6D1mws0JEUzfXAcwVSIFJqGmiSX
E+lVjPvnyhFYIfxv9gGowA1coCTyryS2YV8RUGHawUximo29e2szl7rs9NH8xdCY
hpsiLhdYFFSroovl9Le/WYnIWbvru/erV0LwjzMCaLpE3LRDA0blIHOiXxPunCpE
gnVGgCEfEibnDIqaqATn1U13pXu7ACPX41j8A8eIGq5YhRR5Vgz7O+Om8a1VPeIz
H6opuFBKG2rrbX9Z71Qwws2cHoEwMHYlN9vEIPRh4bdfkxJn5OG+ZU4XTI3dnMym
w17f2ovz3f9TtDCZOfHDQxJLfb8AiI5KvMNG9Ve+djYZxOuDORf9dmhRxLPhE/ce
K4kHk0OtqygYAAhNqQhXZwHaxn/NUcBGo2g++B0symWCk8E3+Xdhnd/sEFCuOmXt
N3g2ISXxCWyIgbfyh3zgHfPwsUBdrbtTumO8niySXsKYibkn7qGhW1kC9kygkOnb
rO/jOM3VbdBDreKk1NiACc61vmdxEFHcnOzVFvoHwsiXaDZW4Z2MtwwFxmt1hEL4
3efDHDw2hc8GCM6JTaoji1HFPYP2TWRq5ofkzRT08umAajUmdOZYSFZPprx3P/GW
rXqc9nyx2MnyoBTTUK4th66FTwIh1Twb7mg3SwucbocHcxdtZRXVXEk72X3OWkNc
Mjdu5M2riuncTJqhoWWZfECSV/gDL1fXHpWHGpsDia6mjFWPied6lTZsixX2OZFX
mPOe8rfhAyhssUcyULsfZap3QJPe1+3+KeRnPga71LnWACmrcOvCWi7ON4OEJQQ0
rQ29p7hh/FVVfFlGPzNA/h8JA4IVbrhSgfQJD/x6wgLQo325fwBIIPCbU96PmQOE
2bQUZvEcGRV0RU9N/hdhJKmOUwovkqefVM7fUwSbJpVqu8Vd87Y/M7+OLt4v6sBf
h70/B9hRNsjJZCdvV8DPbzOl/3EkvjU1554L4Rj1iRjymelgeEHrlcauBOM+BlDF
FrWUBSQmpF7NZ8okJe8lzmS8WDK9+LfCBrxhrXDXLkF+yrsyMHp7ZhRB7kkIlUKq
XtB+mK7LStAy8shGJnbEpjbJguSOTMVO2h9nrhexJmSUwUNa1s7ihkfJTc8EeD51
1xQTkdt/aUfLMCH2hMA2+nnotbyfVP7I6J2mmedhZodI/PMO53g/y9IAmBHcLhys
L5VWEZMm4TN3xhEzF4I6gJKchPOpTSLKcySjtLYDx8JVtuFk0EGpB3ywVqegdwI5
SKzUp7XpbVadK38C3iC0OYwBYEwpkKUUi2daum01/qyN1Ji1qKlhv0OXhT6f/ewL
YWEz90+Zs4ruSytY2jYF/fEf4p2osODsqrARTLm3IQnGDj6x0zp3MZZ9R5TYHy2Y
FpJ7Nl7k0PbfOVTy6EmqhqUErQj2EpID33qVfP7aynBdZV2CC7pumB6sYRKvk5fU
uZ69pvMjo+JQVp6Jt5Jxvvs6n5kguWGRB+yDnT+L0iuPdmVntIT2kICsM5PpoMWo
goq/3HY64IQ2/UEvU3hhKLguLXB+vqglKIDb6adUNE/oULMEUGfc70jazxIVGKNY
AEXDshcS0ygJeipgl4UyqjsxgkmSmxpg+A4dQqtVwU51c78BfJAPOXdxHj8I0Yn+
/ylQo0wKIqg7q9wfT2TL9IHSDiZzPP6qDaBbdUAcbbfXNGid6zKzfZ8mbJHuBV5I
U3UQbdVwdJXYv/PRKAjxGrfdlopi6EK5BpRRobpDWN82MlcdXcl9byv9nu8w78iA
PFc40f1FeZvFVUhAzhZoRg8CxX8KnF3lTg6yT11j/O8JkOeT5XjmD+P+W7pokuxA
p/LH7QHQhTEKFKOfOy8f5uz1vHz+9nHdBoU5ERooS7DWFRGeBG/qEUJyWhD03DBH
AW6tw87ttdewLd6cMEwIfQICf5n6VDm4T6Th8OoPN6sKOoFcaMFE/K0dcQP4oVq2
u0UoAxA7T8H2aenScb6S5rjay6OrW41P/qFLCPHisBVRrYs99z1Vsu9INx+erapt
5RrZSiLhUK/5ckbGBAvEQ/8vXKd6aLWg78wT+7MEzAHUx9jxX2b57JgpJa+66IzU
CfoQvA+jwKe742SBqJDBia+iI/nP3W5XEcqlMKYoQC7Mr1ERFEUSRH92W98L+0Bq
uYQ75l8nrhRK/3z91nxPu735eCCq7hQIK37tUJXXy/oSclSNpAPCTKu8S4QtShVY
8I5v3sZNEdCjhBHmobbWveseFY00j+Jr8A+sqMCjMAXsJuEkXPSM91EVCWg7vZ8N
Vh7qiW52lRXd2kYZon468B+FMFYRNXvMupmV4xsRtXDcosFykIIVXzl/AJgdh/H6
OWkNmk5pKsk/2IEgIJ5TyH3Vh5Y7+V2xx5pe5TFHxnhlzHduefkNzdV8MlislgYx
1YOfa/8Y/Npgl4AZC7ZfODE4FaGURG9pXho/In00Vxzr7oSybXxpr9VL2t56phOX
ALK/l38W2YT/XZddjjex8nXIFyRwcm/4JeGmx8xXv0TCnmKJKEFBETlckhXr7b7f
gYn9YoZOni2GRep0PoH/2c6Yjcw8OlynfBCsb7fNOIWHZ1XmKl/l0WAiyUrPrNPN
PWKpOihh85GT/bvBOl4H+NUYBgH3sf/dxnjYms9cXJbJ5mVfSO82euzxVVq9NorG
IZhZ41tCX8YITB1At/dzELwl/l9eIss8QJt83UG2ucIpQ8hWVCRhZZ1AIfnC9t3e
Z22W7MtYGJY85dNn1Dk65ocIo1U5FGT5xAvqzwzD586jFEJUSbJ9BsP+Jimw5ifK
EY5YlX+0o63YfOTHF49Y/qW4R9W24ywTMfG3dSbniLsBPUw+QeKijB0PTM6VzAqw
kkXMGFYc+oaadWXnYt74NEIaZSEUIAXLku7tG2vvcvS3Ql4i6zJtKiptcp/vynxu
3W2Jw8HJILMLkv8mvK616x2joaIWdVODuVIOQB2Y0J4b7yRviaukNFLLE8/BVicF
eap0SYPxJLlyofk+xsvjKh8dEmzbYevg7o+lCyviOQ3BwYPpqSqT9iRXZMhyOURV
zjUiOiOD5as68cy78GCztm9j8lsdN6nJ3yNzaGCxfIfGZYzuLG78L4mi9XruuNek
`protect END_PROTECTED
