`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIY2rZipGhO+1sNOcmc4hbLQH1c+U+2xDsnph9t8UPHH
8SSkRxtpjA8cFTp711HeJELG1jTsT6Sil+B/ZEZpe8o7Q1UvfHPmYOpNXRN+6jHD
N8/G6/+b1zLNzaNBUiNT3+lsgCPsFRAT10ImiP8omJ31ZoCeVRom1wtosTrJZ6VY
Z+YGZzzpl6ovQnAS/Su7XrAWnFyOETof64hwWrYYarn4cg/wSOOPgIsm8nSXT8El
tDKShvl6uVX/3sx81CuI0rcZanm0hWpVLZoBWkmTLkMRgd/gB0moTHYrJ+4wn9Ev
KyIFr0+AqvDOoGEYii/xSL9FAeJ1i7aLQj5SGc21ckC46j1QOvlz82Z8OYep+I2t
48D8g8YwtW6XtOkI0UIMNGaXv5pqSq/+U/Xj86Hvq8ai7NVL6hJ93A6oPpof9Hq3
zffGlDzlo5kVqX7Y2O65UVX6W8l32Sn/Si59Bx+gf6SffFrvcXxG37t4bFD4MLpz
23lxsf/C/FWb/lhxGgN8y3nwksl4gbo2qrn2f1EtoyAMV/0AoD8HVGN0zfKTSYya
`protect END_PROTECTED
