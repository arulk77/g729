`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
TE8/el71YwffH4xJd9PBFuCbb4KhtwonTnfHpTb6mRtPJC2hDhD04Tttns+KZJ1T
x2v/2DL/ItsabRWgbEd8WOuG2lIN+qTkuhlDdB9DNxfX/fTVYixGY9qLybXszrOF
W/OuVdhYfIW7ApKY1vZg09etdPic5zuZGYeAMoJ9qOUpLdjsnWYGSk8XPmSx6j1U
lXuiCzxQGrWsF6Hy4z91jhZ07yXtpf0lZejUi832/uM=
`protect END_PROTECTED
