`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4woQTW0mQa/CY2o7pMi3mdht1g1HsAJ/KRA6S6YZKkkZeeXaMVUpn6bbSjv3dG6w
Fkh3Bv5vbR/+q038yLRrEHQ+0GpwN9Ai2tDdozZtcA0Km5/dl/3AdWoa83GX11Iv
x9PC3xrOOnV6NqLQmZGA24PvnLaxB9ZGbvusX6iTMDK7d0KWcwJhh8jbLUFxQqwX
HWXzxHooYiiuF9sr9ibGQ9twq+hui+dhP+EW7BWUJ+8rgdY0mg4cjelX7sYhV9rO
0dWIX9Zf0CWDkAf7NT7MfIH/a8ksi/0FDMTY9yiOKjQjLtpNVOXWq72QnMUWrZAW
OKEbeC1bRg/2bkxFtcQT1BbfP8RLFjZVYUuv4b1IoqN1pf86qAmHGVubeyEpEXTz
i3b11JzpP/duM4htPA0t/83jX+tvVS55aHWGF1dx1Jk2gHJqLg/3QuXHX/Ko3m10
MpvB0/c4fKwBxGp8sqoarPU+YwTqzv7F2LVih2fNeJsU2tDQV1gvdREGP0UUTQzh
hICIKxMLW22SLg6xpXw9FQ==
`protect END_PROTECTED
