`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOzxgDN+kahHkvrR2sqI5a9wmm6ZVPboX537JIPIIK6c
aphlzGNRuRWtL6OQE5TMd/V0DTJRDwfsfXnBJnfpjDWb2O7o77uLH+pH3AN/9ms0
k9/fyGTBMr65UvqYbokiN1fc8UmRn6UZdwASm+3FgV4DSAH4nIUUx2YTMyOiPZB5
VXAsEL28nx25VPYIHnImaDuc3rOxSQaOFgiW9+CyqlmRKXeUzfU0y5unHIA9X8Pn
7MP3UGMSVEaDRkA0TH9D0joBXLLNgNzOkSmOcav+iAzrQvI0mdbcYUdkkqpNEczl
qN96PpChIG0xi4WnQUvw/sB7IIOYKCymKVlph7NqsoLMChwm+NyoSDyHQ7z4zsUQ
PS3EpMAub4eVE5lGfDWXE4VbGxalQyt5slwrb+AjZ5pE+aCqn2iLNKsHhhriUHM5
CGs3qCpbHLgtImBLEJLlELqECqQE8UUi8rt7EkEEGfD/hfheZfKgFikWX47lOXy4
uz4BDgq/CEJI1yIuqNYdaLd5FaEckj8ORJhDkIXfx1zm7STw4lQX+KVKVkZ92zc8
`protect END_PROTECTED
