`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44Cfb0jO5fFR23lbHkqZClYtBbp4Kncvw6Ios3I5WHn7
oSdWal4jOUc3sdjd6nl9k5VQM3iIImQ52LrHGzZRH2E9Gg3R9lMzZ4m4MsNIK+pp
6qXrvVxW8xuPTBeyTDbRGos+kERbaoxh8M1F46F5ghV65Ev/RwtNbWVwb9uOc+LY
oc3GU64ARlv1i3L/37no5FooXYRI8s/mDamqBcSvr+r9qgNIyDNAmF9lqDqYIMIl
ySQfcJ18e5qUS5sI6myHXrsw+zsPw8jwlXCu/QDjz5GbbO2q55hMzzDQUS2RmQko
04+RTAwXykOi5cmQbhgu9Mtaq//SrixELsSJsyOFMS62j12xopCkNmvzBwELnAx2
cOopzDCZ9CNphDcWacM0iQ==
`protect END_PROTECTED
