`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOVC16uyrtHkt91USDaodBlC41f6lxrCsSfEjLRHPjtA
NJNPKuZ4Ye9tJ3cLv2NgsobA4Ma5QgK1n7uqOPmAdXUiXHKmH2hJvr+H+v4yFW8Z
U9WWAaF//gsswnDvDMVQk56Sll8bODLF+6f8DUbNdVTyRi4J+3f1SminVtn6vEG3
mmPw0K9AIA8o7uGd7xB6OXJiCaqbSlS6WwMNud5j4HlM5mH0TuqgiJwt4T9YPd8U
`protect END_PROTECTED
