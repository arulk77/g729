`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKsduavHuwmwLlMaqm2BKeMnL8YU08Sf7DgDZtl3/YeT
f+2O5ouWg+SBYmYRZramruLrMh78yU6X0ItRFBL5xKaDk9QJIixZfnaH1I4PdrTN
Cu1AIDKupfgW2BsDZp+geirDVQMvRqkTAYNLEfp8h+fvzdfaOBQpU5whqrnwOKRi
AKdbfOL8hV2kWAFXYjk6x5cDATjV8cE7MG9c6VqUG0gM5G8aUcFHq2Tksr/UfITE
NftpTPcm8aasGLK7C4KxqA==
`protect END_PROTECTED
