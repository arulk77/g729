`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41EJX5VnLRKMpyvJ5alqyBqGrUOCD9vRMhCjAIDSEhh0
Ft6oiVoGBN9JhS+E9+Az3TogYVsRoaEv7QKGs7zmIDtg9VNExeuUQholfE+dQ0RI
hnmm9XTyfpkqXFQPiYP3FpwN2EvlVUjzopOwtjTybwBX/5NK6Gy8UzGdxwjEozGi
nM7smQITBxZQqoXIk58AeThvgOKTv4LZ7jBhKhjiSg0=
`protect END_PROTECTED
