`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aQsDYiSRinHmL3q0IoPuVoEagG2oMVThuzCm+Bn1+hM/
ajUOL071mDr6VqnQbgOUpykJESB/icMXyt6C9xVaI+VddeP5KgSmJM1c38BMwggs
zGuusxTG6xv0xMILLxyIZD8FE1eh7QCdZhB8yUIThd2+SnxbI6w1nimwwuinataI
u5LfOb9KeNVTK8LbA+itRuv9x2Qg6W3r0MumuPIHCbep4QI4BgzJYSCC6vlSCKk8
+yt2HJSR0rvrDWZSkgqrJ6ninui8F0iljABUOFMKfS9fcKAkd2ZFxL2pOQEDBg+I
euChgE3rCs5mn59KdsDjwwdv03TP8Kq99fsoqSTdsihCspou6KB7CUX9GCPvHEth
ci7AN3Sj8okUiEMBKPjUp+II5niwPCRn/461FbaSyEuRK7rcwzG7ZI5AkYoilJk2
pu4xDXP5fJ8BDb40qhh53dl0DJ6c/VJ4wqNZXCpYELxqmnhEPy8BvhosiadTwx29
8G0fnf+Ip4ZrpMTZjFYO6z5NkB4X47U2vuNP7v7opWOINS/e45cZeDEnmRQl8q/G
1/rikEabwpmh/3Qboniw67qrHnqBCkZHaxI9a4OOitq0lEpLOwOhBSQr2F5gbEW1
tcvppUse/mV1NGb28il6iu+GxJqffYDDEOgTooRLDzqaSJiAvlQ9woLxBnjFjr5T
nDCzWYfGUSk+RdGisqPW+2WSArkF+U/EnspYg1KlNT19Xlq/IQ7EwMMxPF9+OHqZ
ZJNEHCm8fyeqQt2S4GRvP/U20zliL6xF/eJW9l/0FZd8jbmOutCyCFVleiJHkIIP
LkTvqadhLmMpBv9arfUYp1mt4+9FGV/+AYazt4afPL3glYDqeQGWT8eaqkdxmqv7
4QVxlbzCNtLKpuR8ni91ssIn2Q7JVGWn/25xAb2ozAJBEp6wphKY5LLkeHxzCh+Z
5DIrcmjPQ/w/m8+fhIZ8VQHoshXE7Wfpw0D21Fcd2SZqor8Z9fEJsKU+YpK7WVxm
DqU3jBaAqt/wWtLU0zmS4/hIxH9ljFKskUQL/6QAl7x6LlBehF5by0hr3BYhYGjP
D69a5bvJP0isVXUXufpoG6e+UoCX3Osblykrutd5cLHITq7rOelHF+ICzzmaP7ZB
K25ltrhzksyaIPRo5PmEiMUh+sXMykzbAoSzCskfmgqyPcTIjW9cvMYcLA02rbhV
8otE4YL/sxIECRrF9dhzTLivYjc9ccgT8TGgASoBAkP1UwBzCkBHVFy2lanox8b7
FE3ImyeMBNl0O1oVSNIWcVZ4IoESk1NrMloLNd7CTaRqiJeIBLN7AXW6+VDK2xRP
YDo3z/kNK4v6vXdXZrdPGOoqEPuKBd4lCBgWXQnWjFi5Icxb10/AmGAaDH8EdmqL
lEc/yNIxWJDg2KsrfnUV778Rc+gsHVwrgGyeOWWi6Styw6HsgYs0eWncjCj4I7gm
vXR40r/2u7Rr8PbFM2PPVlmUN2v+fkqpX00lyRYDl7Spr03YF04xRpg5GeG9/MY0
YGlHuwHP6n+hoNpakos2D4JdbxQOC+u07WHLOcIxyzd/yx8Z47/au1cUPxI1EMRM
S3YWjHekCgo4f5fbr1WYEK1qQFDae7IWzfwUqSK4RCytgNjDeS25iwyERZ0iJ/gW
JiiKfXEw9Gsnl7IlBbWp+VO9XHqOxo3L5bH5JRVTgmn8w+87vp++hi+RgoPNF5qd
l780dNILdlBz4us3qgeqBe4BaFfLBs15IWSrK/YGxb/gG4FyM9wlF4XMZGrOnopK
prD++rVOb+p8OEXaZ20PqNzbW7NPUHbGX3Xikq5Vz7vLSPhWoC1/e+oUWHTnYagX
6QVIHaEZ8quLR5syW98pqEuejcsIMvaspLo7mrmCcYKCfH3csdvnS7lU8vDKdi8q
j3rFJnl4LZfxQbaTBNcLtd4/Fs6zYmF3LwkalTFmVsf5J1Ca5JrVC3pudViqkHGO
SlyLaZQISvZl0W2YlO9MUvhBdVpWNBwMxVS9zPymXs9jr0beJbGpoLVJ9HxeITPP
HtmOfBtfrcrD7FbO+nvqziuruPeHxSIyXyCErQrBhU5BVsTvLgULrHt3ol4JJprv
ZCCUB4MQZzlKPq+WFWT9BErzWE6OVTy4G/Tq1wOlk/5OvuJbvTE+WCcYvoHd+EVB
4i5zfvbjqudL9Df749CTd/SJRggSvIuE+QvgMifwiUSVseJE0AhdsUY/DVufEeAv
F97bz+ZhqX11xF/vnTmc9wAFe5nd0LNuhZIZliIR1q7IX7/hfZzMRRDxW85fnXGE
Wa0nD+sGh+modH6KBT3BLh59cAq2i1Xq31S8CH1bHBFgzHcwdqenJg88qhq7dJcn
+mbjd5N1QdFRyG1S90SrmndaXK06d+OW4Sl+rs5GnnQMgM1WC/BPTmFP0WW3Rw9N
WbXQfogDkqdlT4Ng5DvtuqHkRAhas7PEdpXgUm/vWziflu1TeEV7vzlXQ8DikKrf
9bGm7UV3604LMUOvSynBRG9rnpmgClGYY2KiMgwEpzwepwpgqgljXwGhS0zo3Gsh
KBIXCgQho+fvZCdXUyoj+6UPEBsEuLRmybscSTDBwE8DzySGLpSJMfFJsBUSQmTf
jOwpREpie82Un0+CDda4GucOTmd0tyTnSfZKJIZPEnP2zfWtcZwmR6YysgEFlzkp
f5ryh56xKgNnbOtCT80E13pIfHIPudl1TBeUXOBtQtsN8+Rf0n853mKTz0FmVk6s
IedXF7A5zuOV11OHVTrPg4kvxuf2v5S7MQnhRABjSOsY+b4Z8QQ/gyESjlljVdKN
yqwQP1Ay4CJyuq2cSQsEufdSYuIfpB2f1d/ZHZIx/FV8t4rQWCcPDfJ45B8JH4+y
fQ670kIEZtaOxbmLbkbXl2hzXDpZe6+2tzPe6wE3O+Xyhm6HMz5pU6buhWtz9kMz
E4p70VDjZ+NA/CP5BFBBndCoaUcL0hchl7QSbx02Esd91PHKZ8febryVqeMjcQCe
tiriLflUGug378ZLDGq343kJfH9R2o0G1yGY2YCKTBZOGfousutMCpCFKFPK2LIW
8JwvDTHkw1IWr+YTTCwERvrV1IKOf9o0f9zMdyG1Phg4uBVjD3saafM8BePK0Pws
AYO+ktdtkRJBQ7yUUEnO1blmQWxpRtEddRmHUuUU58JlXlJgGenC9Y/X1TXqBgAv
GpJIB99AZL0VEOjVpSkkZqX/8QD5dtuYEWUukKu5IpmFSqkVr4A0imBKvfV/sM8O
3Bj6GCiaTLMnoga+jj0kRr30o5cl8etLC7beL3BXQHXAiYHmLP0vNzqMzv0Tk4Mb
5RzJyurAc1ZJCZT/GQx7qSTIZhw6Soarr3nLsSqpZqD/eOBr/PaXmXa5z9n8kFNk
jUszZpLsUjgVyL1CyZvBVBn335Xn5NXM9JPhecftKj9EVO6NCSrT4qvWVvibL5q6
NLna7jxDD3f2QJxLbSW9r6UYS6gugea+nBhvDDVs2fI9dHxiOJ+e3HgjYMl4+3Fn
6+EKITwFGk3jBobaIKxR32PED+kumPxQ7XOijGl+jdVWK42nretYMqT/h+G3Uajv
YtqHJlgdGDonfQPfbGMnwO4J8nRYj3bhOatZ6OvGV2cnVRL3bElYYyNx4aZ8jFaj
fBl3hzkFskjKjinxeAN0pb7Y4PFskWlu51V99MBlVOB9RkL+VNCJv0tyxzcqWjjb
lNc/HvtMeqsaZyVPH+rV6BXby1EtkizEwwZ8D4+E2OjsmQoPJhWk3BoQQwEYDHwz
qs0wGsJX4qCjhJfTX6CZwdmyMmSBEHXvLCI4SCYVAAF9Hlt7aoK2JmeknTb++k4k
qLf5QBTGeF4Tq3AN98J1P/G2hwM3WXGwdPGp5v3acIuah9jaT2RoMHbNsfRPUHtT
Ga84qHnsI77ZneByBSmWVl5D6P7HP8WJsmaItIxbJ5jLZVXYKIh2HfAUw4U3rgLt
vXbHKXBMdg6adcbUsrX6dM1BI7g/s0WoF1t7FTEOugDrobBl5ZWGjjEmiXDlMX3B
8GPBZ3eSur8L7kp0KcE6HaknO2r5OiSXNvqVncG6nAiYUDdPEPHEScpkoNWiY7TM
K3HN/DKzaSWkGqh/7RmiAUWwb4wM6uwGzYEvQcLlUy+i7smSt9k7tJ/6iFVb9uYW
Rll8FoeG1hqLYFycilHoEJhzbV14aT4p4X/FqtqXN6axyXk74vRYHmOG2hh6lIAb
u3lUN9tmbFE7UXsnuwqyvfOzDAbP82kTtHSij6Lw7wGIUwVHzMHAOu/Y3uNLtrgu
0FAm68OKhnZNCDxMDbpOyqOEoxejB5P4xwlUHzW7dwrIUzGw/w7vEyarh9EtymJx
v+iLnhswpwfKK9ChWvs2SuiH+3wjy2yHu4Ysyugk8EnaaPxKmUZPmavzuE6TsFsd
2bNFil5+hPlVmk9JdRT55RwAZ1XtwcoBsgvdZmeU1F1ZDF/VUNy0Hl1FyQp+QCEH
8kQk0NXnk22mZULfo8RYxVvdlMc3XXnTOAWKsRnf8kARgF9Usc4k6IHqNKUfd+Ly
eLvrPDUdV6M6y8lNFnbTiCNfKAVDCjlRsXlGOhavKV6vaV/es0zEzfrDogoeu9Te
snvNQMtTF6dRgaUTI+lMsPINHtOzhD21p76o6+fijp3DPKVzc2oSaIt+6825Zbnz
0SCZnw7/14NYwua+Aqxxtq2mGRmZeAEETTtxz3GajBageUHhgEcvqNuQkxql4eHl
sT+W2HgnB50t32J6wK0OZwFJcZtugPpntwbW1/q2h61Iwnjj91dbqYUe+Fk1S17H
+z9NBkuut/eeVMvfG3YtIGmN6J+NmY8Kt4hqkHzTEfcDEJr4wk3XNS8YTsKXwjog
lyxZtwRu0tGuSd7CoMzb+6laF9Dvh4c4u2ri179NNtK99zqvxmh1kj9l162iQnik
cxtAsxerh006PdmjcsdMxcVZw0sUApiLyhT88BHn7pVsNwoOWrWmyBxexpkHyvW+
zECoIdwtIRkL9SVN/kx3Lo+OiTyziYedPS8dgT/smJ+SRHXAVxBbN4s+t+fklKrK
H7A076c/R4gMGaP2KY/9TCfCOmY6CazQVQQmtdNuwlDTg1XXeUlWDR4jPcIuA3kd
Z1E2Toc4O5SIAXVRvUP1Q0AHgp96tgXkMYk3ghZ3N7P+CJ38m4NPN3926/WoT5mx
0JLjtxld8tjv3tfkiqrua7M2INoFnYCwK5hp7+Q8Q4N0fqmdPQ5Krq79hwIu/x7J
gZFBMEzulXibJRcqytPiykA7R/kayoE1gBfLVBIbXTcXKRgAmhjKqKo5z9s5vi0s
A+ir/RT07MDCPwLhvGCGaxgh1OkqLUP7R5OcVEkuBKTV2N8c7gMwfmhLna4uCuQV
+TxRuwpmPHU2/wnJIy+oFgDQYqzSrprfitpDMkY92bksFZiqMf2ThpuSzReB5TjX
Q1gY5a4i1TQl4Bt04UHtsJi+nQ+xtYMVHHixFaIaZl3dm7EgKHUUTvA3p+HKaeQW
L0OaYCTInf1GoEbvacXKqPmwCxCg0C2P/CcgEM0nyRgdx7UrDUCTzLjMrHCU4Vnr
mHQY/4B8Pynmqd3TD5YaEVusjGV3zoFtosWjFWciGFIbQOzuIkkb5OotobuxuCll
ksTgUkoNg6uuawEEZoGhe4O6BW8OY/2n18VmAmd8DFx6ynmLTWoIJBldukfBrSYi
Ip2PKfsASFqDRpbn14jL56oRCnBdfT21/zFwYbqQSWZh1KBnMUIRr6emmxkK/TRR
PP+MGkrju4G5Vhn+Xr/Dwrp/r+eFTw8tAZSuHyxuCvrXJvXzZFh/1+gyzqNrCqEB
+5KOFrezKPHSUROXPWTnbiQlluhY7YfNeyyefEa1+LBR9K1RmOEJJW69rXSIJLrx
FeX7fZJwvqlPdrYUVlX0hHJdAiqrSMNDU0Iq30x60voAcQb4BOPnKQub+5jn7KxC
b6LQNaRqTsu+rfBI40cWDNH1DYkHSMrIQ2YXlXb58rZchNkhW3EwwnAbkzd1y8GS
aDpQy4dfqrE44llTUZVTw5SYTo7zrSmQEfz5Lxw9JAFevbQTWy/Vwp6AbWUzTWRn
PklLADhWF3QjcUk75mCpLjnyUA+oA/3sXO2/kT1mMKmlN5QdzjJee95yHuamLaNc
z/aD36Ekggz6POVMdObnGIEeo+JzZIz5z+m/Im4qQq18S+bhIaKoZa81eS9hBt3V
BuvDOCoXLKpdL7a/Mte/4ytS4maxv2+ps85hvuF2fN3N68buSiMZPS7GdCHUPUM3
EZ5YIT63x49vkrBa+BaID0LgDNBTBqqv9BMLXzXvQIanPTQmvQWlvV6R65nUlyY3
/XbCmb5nNf/xATrPVjhbX6t3axUchtPiL4r0p1n2yqZTVzsmI7deBnGZXlt0KUVX
83RPt4G2TX/DzlXvY8gSkCwYgdapMDPMUO66JMRODU+7icpqOqBwIrwYztebjUdU
agYKwgOV6GtTMZNuQ5W5Z3z9VbNW4qYSCVwkhM22+PNolr8bOy1bNtNqZGOIcxuy
EU0CToy7BB39LvWQzKS7xd+B6J2gPtI4fHOUimv3bgY3HBhgGO0WN1O+5jsHn6Nv
aLpz4CZS7aY0yKmOhSZC7UqgPIKr2qCEC4ikPMgcX5pbCIfkCncwTOVyMZWU/4u1
VO4X2nFP/vUF+ySu7Hs8aC6HjPtUFIn6sgCiRfvKcdBMa56RT3RV/K+NRnfwWCcQ
cqFgPbNVaoPow4Z3Gug47cIehkW7l2SYnN1WV9uOjJGJq8mD5vjqsaGM3hS9iArr
2RGucZTXEOWngrmsD/HKwfEouJz8JyfXF1uyG9EbHuE=
`protect END_PROTECTED
