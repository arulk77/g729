`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47dkvCr4dzrR0pomsN+87QTCBnjcUGarzr3blKRsItTp
wkNuN1ucFLwj9jVIwlljwY9hxGhGEQvesjhOIWOq7FXrOiW6dpm03oBrAUkWsLtv
ic9OwcTGIUvYi/T9uoODjMJ0RtHo5IzR9ecoP1U4e7ipmdFJGbhjzZt/9AhFEVPw
S92gigW5YNx+Q7vSjzUc9CKOeV78lznNadHLablse0qpRDRq07L+gHEXcNGnVUad
w29bN7UZj6VJ+YhVza5qZw==
`protect END_PROTECTED
