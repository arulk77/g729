`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42biP17h6SCx+N3eGZ4IzLgHksykwQStxpd4FN70U5zk
DwEpKFsSRVIP9M+YIdTPq8QhvxxQUVgtlNcDwnlvHBZRyNllsnk2/1BBZxdWbKco
vZaEQ9Kwe7v3nPZvv6vXKjv/57d7a4gyz+uO3IoN9KWQ+l4nlcXnIQ+1vDdlsv8C
QAF/uKwpsiaYxbJ4wadc+DsECjzQLmDHjuEKE1xSBTIHCr4Q0IxgDCLfAXA3oUl/
y+04iQG2XabYuRlaOCWKVnH//1QuQQqpwyikTqh1S1noIFylBx7jMGq7KftAaOAL
PKB4wW3ebtFybdI4B8GoOG+pTN9KQuUv4YwGjPQtAUAFdAmpXhKtZ2dTW/gnXFYX
5w7R7En3wA4Lt7HYQxMP+Q==
`protect END_PROTECTED
