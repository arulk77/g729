`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDx1CDSsUYbtASVycbTym4p7iJjbBahwxQY8S1gBA8wH
bFGzBTb1ziYWP8eYGqhOMRIfOBQl5lQPWsobwerhCf894RhlpYN+8eDAUWg0KBdx
5MKVClIqlJ+AkGuY13ym8JnonY2EG0mbpgyyJX2qnhq2VNWdYzLiFtfIkAoZlxj5
9R+EEc8Fvz7xrrQkSrUop09h6095y1ATaUgI9QQGC8o/li0YijEqaW5MfmUTTj1e
MJ8u5/P91+9fxm0zyM2vpteEfFDmcjuXVmBihzswT2TA1wKbLuW9Hg2pa0dFCJXo
6G5PIXfvpZWpVV3ov1730Vs5i3C6Hvx4cL3ytEP8a8KFz3hWo16IyxMUuPkm8a97
OSUMnr+Jkn9A8zqMgr3Hgn6fEEtO14KPzExNDAPTtmfDuzynCHGeDJlAB/qm6eKV
7YDrhem+lVcYjRuHy29AVrWeI/Tcrhz1Dhiy+o0tGll9i8XUxUe4uX/x4hzrDO5J
E9ln/s1lJ4J2XFAFLJyj2CXOpbOborh+sIgzV1IHFYOsq9mk/ScWuEfnSMZbzRdC
UlXaywZhMx3IGaXbbko50eA913Fs8WsxDbdUq5gUPql9l2TTtF5emmTG/GjMkmnk
6ZA5xgQBq7fGLgpVSLoUH8UTRIdXTnp2PaCDqRYbtMLlSdCPJMW1kCLJ6vTPBdYF
fqxpCknSP+1ZllU09K3IsUoAiyNNHHfkenDwz0K60GKJirc3jCpP98EH0Su1PcYX
UJbTT7WVNDU80VKCFZ+jfSSAaRs+uIWANQ+Ls+W+sl5P6l5+m9U3OjTM4CecyGqy
xSNA5L9rtgjnc895AZZvrau6/m33IMf6hUe+PPyg5P/4kuZYb2nYXXoPgkQObw9A
QspkDCtrFPCUDXm9+aVV8EnRHkx1/mNV3dSopIbChnsGi67pqX9OIHCQ6GXh+XKt
MsXUeNiwmOQglLKQZH8RUBu+UdtVKpkNzcTqnhtaoa/M6DBIUewq6cJTpmrj/tPH
h/Ifbu6teMz0YOnwGaql7AMmzlAIxdJge6Gk/tgIJSt22F1gZjK5PT7+urqxMQoa
P3rStCp92jnG6Vcqvr7nxCc6xaqduPtlhGCFFMh/iGsaDsf0jlli9Mu2Y85PviEo
SMU+QQmBB2fQJYpO3clK8t61JNcwAJTgOoCAeTmbe7Nisw0lae8kDvNldWI664KD
hvCCpD0goNSjElvz3MUw8UKk2KMYHQ3GAG5GTt6hDgo75HICChUhpcrVCcC+bsPE
pdxmuB3xnAZi32sIoE0nDdVue3LC6hGRRuf0waZz0okfqaUeIa+DXPZnCzocuRjH
hqRd4bAMOQOeW81hjpwa+rqmmZ651hvQ3/9IHyORB7FA5ryKcNua8RLMCw9gebLc
u02UgzVooYJIdu4SnJ1K8afVf2RrP69OnYD3ek4x3L4UWw87ugdVfzfBumZOdNh4
Li2hcjZmBsBPQWkNfnu5J5PM9IHX2EKJ9Rp8CVuEt6ZvYV7zqobWWzmqxpRRB4hO
0jIs94ZUVWnhfz1Bg94SLRkmbNSJEh4VArcpamRIp78NKgm1Zy2+AiyhsbQeL8mH
wkw9yG1I52tgzgjOIAYm+VDw3x9kkoSXuMNAd8DpJEmBH3Xg3bnuoP5FbtcNJ0dA
OCkuQCXtcLyzD1OYHM0khBWjD7RY/uYXv+2+sg3PbxFCb00EU4T02qVvY3aAo0S6
A9RbzvlsqgaINJjnwFzW6G2LhnSLSaQUthgqcuaYNFqiAYMMs34Rn83TLa69WEY/
7hdtL0JPEUlzwJa/I1T6I8j+QP9tkcmQajG+8TfUAvGVS0swugSd2009fFfqQQCG
YDsC6T2e53Ff5OrYCsW1kb3R8coGt6JLKVxPzbyk7wnksCzmzN6c5DTa7fGYtWWa
btz7sgtqThC8r9brvfBtzejTF3PPk8iQkjGggfWTxv54RKzLkBuKB6sBCICLNs/3
sjwGzbcZRDAlzgtu1jr4/t7Vg4zGo0YiXH3y4zLFZjNRggzkrEVFgUCMmpXE58C8
s+p4U1/hiZCpGXQWtbwZPc0PpM48lhEl/6cfXX0E3CkUvtZ6TKXs7MKhIGQhVuow
6JlAPZHjJW9mBg9m8lRKmOlnQkwUVPWykDxN20ulhjXtPhLAQXIU1+lPxCmuKSn4
iUrYj2B4HR7F3OTJi0PSIOuByAgUHtg+eDEbsXNeZfM6IIktWfg2AHXjfTGYBQDo
kgNW0VamosER81n1t/Xh/br09Iavyduvh5tP9N1NVAmcoiBv+T7oQSl0mzJtkiGh
/D+AnzriUkiYXjWyxryYqy/4ENedKQ7PO06iiptoB7Ek1kP1+o50FTJDhsU56UXa
1x0KR88A3bBn01vUt6VpvUKL5UQOGAqf0cnJayAuLmyl7T4SLr78LIqDHdtF6TDT
iYUlfHJ49DpBHd+d5ZIyBWS4yMedGaudV94mG4w8xUGJ1ENo9KMqYgtgwG+tNtmc
zwoVb1TjHrUdpUCKoSdoJZRGGnFTzo1dkGVikzRm0h4mK7F0OXJJ2Pnxvpm3TDnI
qjqx7w1SgBWeb20nW4u8wG2ry7F7DD0qzzVuY7I3KvaUheiFH1laVLijAiaauGsJ
pnYvlHdCR0lVDhX9ri2QO7wVSzOCEOm0yTAM+wb4ePbQGXwMdJ9LrEmZ2rWH+aRn
I6phCy2k/nMVc7yq4/msIYbNi+0Xk+b92Xo0FZCZyCTOverVJ2xec6NE8z2Ihk/p
iFewQtO3XN2i+knDR9vpQJzrpZRrQVa7GfUbWsfn9gFS62yauOPIiLN0PXZqvXWE
/erSohCh/PgGXDrwMSsZRuBiZopmq31smy/t+R9LG6tENIkS5J3hOIZgfYalznyh
ih9FIscTPQSZTgzeB7F75d/bzNLNNR4HGrltdndMQf9f5FyUqZQF4uiYhFf68wej
V2QHUZZSt4yASxmgpwDqjWg8nskVpHd2LLO/6jSoEz/dsHku2x1Rik45KoUB5ctt
kGeVV2JfpbdfhNjVgrC+zA6KiO0PMLfXBBx3XwylYWgTeqoweUIHgmOGMkc3N+Vx
u/OWakAG9kQQj/xzNSULwzAVDrhjE6YFOCzd78pOMlIqAP3s9J32xfUd/oOVse0h
0aJBTYlFXNqd3/+sEqbebiThraEqWtUhv5PtLp14HOBxwhviNGew/ie7CDNr3IHr
hddie74SLBOU+OPjKJtAu0rg7jvkAQbE8dfBOCquistJbxrzeSUU926yDIS+OCBd
sXF3y4p2wbZE8p76lay8xlJp/UiLfWF5QLvwoyZ/nUHf6vXbgXANeAwd2ypOfRqo
WCqL2kxUqrme0/F4Ph28bVs04ab4sfAUc2uBHczN7+IYuwG2+NVWtQx1C2mh/TFE
3WHF3njVmYJhRXm+f5wBYCugpfqSrwiBDj6svqoGqo/Ef0JBJTBKvXZci37n8HPo
cyig7+muo1Eia38GnrvpAgne9AmE0d8LsFWS/NbOnNo0IL+kXoTaWen0mxZhBOK2
z3Lf2dpUYZAkmRzswCKFygVUfKxHyAxm5lM1jzjLgaBKOgsgtCYVxDREGvTkY71j
UibZB06jfmlP37Ai5U55sLhAaAE66bth10sAKhzm0MUOi1YpQDxKdkTOEYoA8FcI
rZId/vLbIF0uQEJnN4IxxN4Mq9uotogD+MZQcz9fFXRgKhnnqsWcZLQF4lswX/1G
IcomulwtFBNhmUk1tbzspKIAQMHtBu1zB9LG+tZENIZ4yWhHuOq1iUErI9ZQokA9
oS5Kd4KDoRWrLQTn2X15fh2tC52bACyRAKrspEjXBHBkvXdvzA+QEUZrrxIJm5iK
YBqCynv9xgzIC6kS17/u+47fRawZnYa513CDAyYdbGKrRZo1SXXZV004qz03g7DG
+O7ItjVfqzD9rujpAA708htoG098nY2BMwRT1utZx1Rzh+u1oGmbc6RRZTPCDEDR
u4nBudc1idEpbY6UCeAOHC7qHHMq6j8H547YKocEvmbJjasGUq1NLuAGjccWV0me
4h8I+s2bhylkueji856voBXl9e27m2VoT8EyTH9C4FQv/dX6W3UHFKgrsptOSLk8
XNqsknPglYWDwVEAmCPlkG+joyzCcorJCXRiOeRhI6ABKtp97mtXlaA0LJS8R/Ns
JYKLrPcgJ2tvWhcAzSJho5WFY4fhmNp6/xapo9iA84x5N15UqWlxlJIw0wK3gPyG
17y4osp0daGe+QBM4ym8UX38DOlXMvTDIsyGS8khZqijGCikpvfYFK2Tb3V7UbSP
b4uHk81VjtfWoXKNJ9zPn7VWCTiCTSVDm9kmYDJyy2z5GIc3heMjUwwen8aC0Hen
CXeWY/FDm8wWTI5gXTMN6UNEYrxZxgtjE+oXdCg7P33wEjxfB6I/QioMkAJKHvH2
aexZQcwnLleow7x6C7dI0dEpCSQQEjRFLtsePG0lx4SA5w01sniR5gm+keIqZVpt
RCRN5IHGHq4li9b7eWtqNmVbydc68wHKzusjj2KzeaM96guTV770BV7IWb3DOIlf
vm6AreiJxTA/wV1REKvwUvnBTGJ8FH+x+X2PMhvtIj8Z0R5o8JjcbdYvjyrw1Xno
5l9VvyXzp5RvUBXKsNLtb8sAtgbFDIHCy7GXdMTAp/f9plJm15wC/N4xhn7+2xlN
/JhmfIa5POe4yAzVugxM0tS7fjBWsOPTU25k6fDipHritFkMgJut8hWlu0RmWdNt
`protect END_PROTECTED
