`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43sW7BETxaTCGicgmMsfDoKHri7nVFGT01qscc9DRezY
VCM6VXJU2LQTtAqgPbgI51G8dNv+YcyDDdX5UNkcmx6bHC2iXIx5CsCeKEze0SNt
5XuTPcAx7Xvj/Tmm/nhRDtlUnoP73oCJ+2mOHXOQVc4keBHW3Tvvd7T8144p6xtG
lCjbVN5+Vq+4KGjMvcZmBqe6m3R+F5hkWsAlMbcTYAU4bwG/KnbgJIGnEPU7W3FD
luNk3NCpKjmn56qbYfL5KqxtIvNCjjUbRTS28hPzJBU=
`protect END_PROTECTED
