`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHpR8LwkWIWj0sK5+KJnkjtdQL+4tno4f3CzPjS+i35j
lg0/OBScoN3rrVOnTGWwvcmGKs15f8tSKos+xmIg+tzM9vnRPBQZtT9JP8jABy6K
FH+hGuS2rD3Vmw3ivpX7SWLHJT9S4izAU3hwxwHSzH8bCGq40REYSsrchifG90DS
VquLr3YqQclg+wXVs6nz3RvVo9lcYIlgF+a4PNIPuJOxIyKc6+RA4+ROsyPoviRu
CBPLelYWcBYOyXB7nSWusyFH08ZtuZHBIFm8Icqho5RPIBZMPv3pMK8LFrXUhgXA
KK3WBHEKJidKr3+Y9o6M2GNH551qtscc68vV7gAEgv/nOtuNQXVUMCnzKLLuwnSc
knGBYgxu95XkXJZLJ6FKLjwimr0eSX0y0WtJ7XueTHS/qgjWzLwq/oI4xF5RX5To
`protect END_PROTECTED
