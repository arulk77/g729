`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKVSfrMoQ7VPDC1pacFKL/n5UR46fv/D/8AGIPtpT8aO
BSovLqSFyEIPXUXRzi85fMgLowYcl/qLMEYMuVa+KxhKeQY8hQ3hJztt+sRtOzpz
hc+2A79+alRKKUTQnovr08fBAjCOTrZWcauiPMQ6XtJtJlc/oI7ht3ZIX6jG8Ang
FlrY1LnAvxi12E5kD1zydBnIKEoX0Q6BjeWcG3YlbnOd+FFFy1xiZliWVAyXYJ1l
ghK0uC7O+uXJCoyLbAfnPA==
`protect END_PROTECTED
