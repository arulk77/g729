`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wfz9/hy2WnQhgL5JSUsb39DNX2t3Fg9YmJp2My/W0Q9
ET4vZRpzwXTqQy58UhFJvRFPPvbmcrMjZr2AkOTomi2RwR7rvL/w/tFDRj6Gv+yY
g+zOZV418gMa2PCnm4dhLj7ccjMMt6LK9JHcZjp1Nv940UTeJbnO8TF3DpKQOE8i
P4LYOT7u2RdR1dgBLn+YuHoiR9WKJFSs9DGZ6PMn/ZA0OUq7x0P0SlsiyXyxijSp
EwoB8SmDwRQgUHLx02RCTqEmuq6O8sNF+zmuRq9b+sIRoCVjtEJeNukOlET/0L9w
CNMEwb2gP9j9lFSkz1wAIw==
`protect END_PROTECTED
