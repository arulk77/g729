`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDcuDgqC8ml0BAW4XC0/kFvpFsZCxks45+9wYzt67bCZ
Nbsz7jehQQz1He4jL4Ea35vBUUh30P4A/K9TmYfoZA07FE4TQIFrrPVFOAF/8lK5
1+PuIqv5DtI5JJ/oBTon+UBQ81Biw+9rd8XxDahCBZ2zBi+wPZPab9WCjWZL1Zgs
N4IANKW/5NNeeg5txf1t1zNTzSnjV1Jrhyf69+YSp/oECrRmy09t8U4OHCg9f6DW
oa1j/2E59Ck/dJV/9RMsKAn5UbdMR8ic/UPbS+CfhF5/xfTsq0tth14REe0Iv6iE
MYBC39G//TlLv73CC524V+4byPwPVxmSGLuQHjJdNSSH6afb6JTNhL4iD7zcqUKK
kGghAgVj8+H7f/PaIrZcjRG5iUcVGEIk3/KmugljUCX8O2XB1BXlKthy1i/QE1P+
fIQIRQlvRthfLQEJpxmOP9s9xDs1d9Qkh9wJr3jzJxK+eTmAIqx0Q7aTH8dDqMzv
2m3Zuvz2LzBpPNkiDp21hhjBzj2ws399TrVcEEYNfNHRKNatJBtCSC30QvjtcQyH
AlvTq52lJ0YuUdw2OmPWcqQrMIROAKclh6v8CtoBqVjVdBMA9cGKOzLycJiyxXbC
3Pj64G5r/nh/rxpI+WW4MK5X/fBTOs4sefCvIH4AocBDwIFJINjNPswLHJtbSEXL
mTyd/Ba0FgvtjHkUAnANTGx4NVkzoZXEs53qXCZAxifFRuYzC9MjCF3yQz0oSPqE
t3MtFlZ99WUdZ8nrLxqn6awmAXtrvsgEUVqRZ2UVOTY+KRG88kthsWzorO4NkRWR
`protect END_PROTECTED
