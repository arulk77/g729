`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43Nmp5FATg6/9HXvZeSKM01g25xdr2zsZeSwRv2pjk84
8NPcqazr8InlBREexfTRDmNpdA3+PZRtwwwJ3fFBESP+aQQ9NeNxKKgx+qHBoyLc
5UO8zPfkDgK7d74gJ3/amIUfX8zDFCfD0JZw8S0wymP0pPEej+DTTGddHnseqt7t
K92lqgt3cjJCkQ4qqrr4arh0NQXMoLo1zY2a6lm5Yh6Wk6fJLuB0ZAEofUWrDp6H
niAXQsi6ZCkR2zq+HHEFDG8tBOGzEOC8Ur/1l6Z70XYETOpvp8f3iAljhdpOHdlG
p0zuzTiLWBcuMEUhedFaqViUCRnTyDZjD7EZzTPveh/S14dSQNeP9xQEyS9k27JC
se6aAWtUTz1ed47HeJ4EtQ==
`protect END_PROTECTED
