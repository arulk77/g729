`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkTYujNL3NKn9eFqAPx54bjR9QnIcBbc6Uz5LvVX8WK8I
zrc7s+FH8i3siPqYpFGjkVEL5V5IqWIgrqPIfXv/WGQWSNttmxUbQnIKdcXDY2Y7
vpbVZG5O/JKmEcjNaEOMZ4C6j7Ts3TkwD3gCY+Xe/4L6oy4PNDx0m373Ior4saCY
J8hgESeDlP2uqPBn3an9KTkXKp4Oor7buxxy0itF3Aeov+P0IBYE06TuMMa52fCR
0QTV7jlTeQoNiq88TcH9UkL32kcV1ElqjxsHc3GZJkzm8H+/S3uEIQPBcDPqT1U0
+ESioxTUz4Ensw/6E3P+dn1DR0lxYBTxZVYjmqSWwZMAGTcvdDa3iW7VK+uVuWX6
j0qG6bn4CIt7FDaZGa9wdq/cmIumXF9JurlTre6o7Mu5lLg/74+3VeWuMhD9uXRV
+J7bQYqjdHoC9+SQcCNZpOVB9Yk0DCQDzu1ieaSQE9G6+ic6tFDLOrkb4wF6W3cO
Dym5AJyAaSLk6XdDibFtpLEl/JZmgFz3eFlapihfAbp39dlwkOvPyi8bOwFO9BC2
4tdJTmEGu8iWBdadzdxchDwufhC15i387VGxBIJBk+3DMACgBfV9pkJMfupLzRK7
IK+l74KgudluKWg4qCHkXD32cvnVhgh35daEsKnapa83OumhNbvvVAwWooQE/CJW
Wv3Buh0MkzGx8Q8C3mCnYwi+3eSoVwfGbUIXxGOe3osOisX8f2ANl3/FCMOL4abD
k8lHj9C611ZFiwa9uHdne7PMz/6KlNEVb0A7QMy/ODF8Ze59g37Lp42JLjy7DCSw
3J4GQppJYO6EmV2jbwIduA==
`protect END_PROTECTED
