`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47uORCVKUDMggx61qVAgHOe8WKvu/wNIeJHga1IKaB3r
aOmjstadl7mMkP35fjXeIiAEap8LhtbqpcwV1AJhqU17xeBXKp3lklufISrvcqHt
uanBiBvHdp3vaN6iKx6ouRFlmX5AQc6a9NB1+NFomXFLO6Iq34yR0tmnHXaWNpaZ
uTOgmuFIzag0FZ6oL0RlWWbs77coCUEUWLEH4Sn8pO+yq/UP+STDcBXa43dWK8nl
JJGrGaSJtwJdNo5BweIvyS3kKIdibxScA+YBTTwcX4Y=
`protect END_PROTECTED
