`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C3UOLnPVNyQiHfuYg48YIlqTr/J9rB2oW+1ybh+LVlah
zqyJ+AiLMwlHl26yMY6RKQ4jdglVRE6rnf98aU6AGFUITKETrNDtXWK44TGBCCuc
Va1Utzaxp99+BDOXAK43UEBc2Vus53RZ+z+465jqVIPUI3LklpbsDtpv3MonDp+D
NX12/i4G22BjH28QHQEfTaqlZz+vvPP5Bk5Nd3xEJX5VayzTC/+UrMuALaIzYQ/5
o7Z4VBi0UrM/wwLhACd0/rDoT6F8ZRhaadUDfQW5C+8XQCltUkSpu4cAVQD4vbYb
h5RR5+t9xrN4qGItjQUUsk4ID3jTvTzHdWdn8GOcpAErK02+25NUfLqi3qozKo5/
6MnBhaVt6YuQPR7MHKSohRHk78nXph8oyKYpEs6IER563js9Kh5KEs5YtCRh812N
fwP8TmI7b8/7Sqkk39RK8EJxBgwNBhoJgGy4UNvJcZZVGkHVFxfS5Vxp1bBdomg8
bMuJHtcMjNFvQ0JgeK8NNw==
`protect END_PROTECTED
