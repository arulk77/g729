`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAmAwDOw1GhDQK06RMaADWoAmKa3pDwdw1bQ8qxc6qbp
M6wbQa3G9riIz43nlzmw8rcgorc7GUcT/UopzHq7/JD1+aAQ+0f+vFedrCaIiEj/
Q5p3/gYCBR7SYtmjtAVsL2dwKwIENbFRI9djyUlnXIszXJzTZplQE0tTmVsQ1m9a
ReqloCtOXflwjX+fin8lMBiD4fkdTkPvx1XMQqEHYKrxywKyh/TA0MpDyeDdcb0k
l6rqd3H33Qj21Pgqn2/B/KQZBPCbfYmQXuOTfOPf5DMbH1m1mG1tMQfYIHHU+Dmj
+6NPRxHl1EyCc5jApYVLL/uYe2Du8xhYbtIUCsn8ow85D5Bstzr8K03AWPwwnQzP
C2OXOBdJzXUBcX/7bsTjjEmnSZrlNXtR4z0+iYMrtioDK4xGydVOXHxA7anv/TGP
WFUgb+Vxx9ZdK1i3tFpPO4XS9HHcSlR9Ngxpc6/4xdfWpDmLdDVtahgHyGHeSF1Z
6GmMzsXkttV8YEXdgLFOFu8t+JYVa744PhswTTnPIFQxbWsn4KU6KdmcMj0CEQ7i
l0RddeGGZYlFceCRHeJye09XOQJ4juIa6FS72D0gqmCmqBXR1fBmSa24ULpWu7bP
WFeQSDNbs6Orz+SU1lKJH4Zdy3xCoOXDo4VNwQcRJgQOYKIaVowBFHNK8EzNiMoP
ilb9YoIejKY6eEiSPRuR1no8zMB6FsGHVozol/DUy3kiGE21l0zmk/KzFeLnzWxE
gqhdYy5V/rXqUjt+x0I5FXPjhcLdwU8JHOQ8/4oPIfSIyzAXrrTSB42zBSJcMI5a
OhQr9kG+52LYtCBGBt9aqcPVEIU/XU1TCRyf0SDBec6wF94pSYRTdyJYCnp38UQj
meDqw3eoeQCSfQSnE3HUPORzmFlsqQlV2PaGaxpTHVY=
`protect END_PROTECTED
