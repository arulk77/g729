`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
BLgI0ySvvhf+Ugp4fjw7zUvuqs8JpSZCB/Ac5uDe3Z+gAJEc88BT0lRWKYXLwnso
FxukE3WpAQAKR4vhbYr1VaViJr+ssIRcFtAaQ27x6+GOtuMv9UsUQQ4IsxBv4+pb
dvaAhpQrDNwaoaTXLxQ2d53nhqayajU/8+HP/M8q3GzVEJvOOmeMkxd06D7sRgO1
`protect END_PROTECTED
