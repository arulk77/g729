`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu414j4/opKodtnu1Zf1XEVgnJHiZYp0Apwbhsj9Bw43JB
RXmW5lSGz6KSW5eFAGRlywUxu/1hMtUUeAsZgvMJMTpjEnZmX9m6O8KyX7CS6O5Z
a1zHueTtkw19YVQKvIeTuYghg0zlGa6JzcizCd5b0cswEDxQsjB9QuHafUrUYVpf
lreWjtXPZ1WM4w+YCWHxtN4sRRVf+WfiVlxavtCYI0cW0ijLf8C7Q6BHfe9+/w0t
dQ6ZHExAk8ZSGI7OQblWyt/2GjCDIwzpttlUQZQ+2yYcBnLH/q8RKD5Nu/VSvcZj
4fzp7iv5o5T274d3FImkRVJpfxZExAb2698ynjAcwilrtphzyYvrWzu3yQvcFzxS
AGC/wyRAgz2m1w/MyycalA==
`protect END_PROTECTED
