`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48h49rI4kXq/zQJEh/f2qsZxLrJQ4D0MCcqzF5z2JggR
9XVBsC3GrPptsqwSOqwpH12h/WmX/0qVSEqDBr28E/5vQvEAwJzMgJS+vRZ1sBNu
rVMzyGae6V+20/woV56qTYZpaFEMfnnM4HOmcV+2uuR1HClhEtIaSs7kBXsB2JR9
vlReGgbVgye066UDG/AaAPQVMfmi8MFEkXAKA1i8IXCq0zLUaYLSVVNdUt+rDa8k
xdboCHERt+7PTBWXns57FX6bcvUgb923EcTcqdPASUpYrMUZw4jUHJqzWF3jyEx5
SgqPJfPjeHu/5fq72rU+CQ==
`protect END_PROTECTED
