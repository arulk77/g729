`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKDtfdtXEB6GU7dZJDGW7Sn70azx+gYdEdYBcnhwVnf8
DTn60Mjc8samg4i28LCMylFbzAxae502MJdEJAtRrwlrIo6kHvXJXYmyroxG9beO
uZR6rxYXL+fpDZXq3dmXJEFLXA23vY0PsrOmauy/dCIT7xzP2szwzHXKRTWEeztX
cP6Fyw81qsKb0RZh6r4pkqWCRNm7Hiy7Nu10rg76SBupyqtrC/3811vE4L5QBoz+
i0COvv3vXae7kczwF/Mk7SniNVJ4RmczfQqUALl7VYTRwcsAb4NyS1rPUvwRXdDy
+3pU44jk3DXHKJPh/VY87uWqdZigadstlvvHzcfL2p0qfFNzK303MaDGO5QjCBzO
q5wL2e+W1k5CxIHoHj4FKDzrPxZcbYNzSkh/MuZjesPFl/SjeWJ/Pg9+uAA8ZSpo
OrtSEIXZ6dW1spQtQJm6iNh1K+cs6e0vb+wNz78mF0Cb39yU7wXAaQ3DuWWVBGsY
Q4CSaUxJwtppEUJGozf35RHpb6oTj0G+VOtX5CwiZoOWRt9lZaRmWOh2/PzXpOHq
`protect END_PROTECTED
