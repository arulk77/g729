`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Prgb+lMGK4ankHVaNnLDqxdcxP7ZuJ43FmpWx3YXsdftYQwV0loitHHFM59amAW6
HmDOedzHpDM/1Gky6bU/tJX/StI7riqYU3jevFupnlRpibZSSJ8CgU3YlGM9HGTm
7dt1sewPKkmjHAXGV8DvjuixQVOaWGm94qVxr8cwjWvtORLXA9m+tj3IgqYhPR1i
wvn8N7DKu75NKZvcNvfJnKS9gOyY2yLTr71pZvcQXrDzdo1UBelZKSi7K4A8l/Q1
62c2Z23i2JFqOPJaM5W+zp8/o2dgGgivN0j/1SCni1N/A43tbvO/WYZbidVWnHYd
`protect END_PROTECTED
