`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIj3fll3X/fLvvOrfRKBpskMPbrkOfa1kljyJ9byaHE2
+Pio9U/j0UMdnwqUxyXLdXBc4xTMfyH9t+emSUDzW3StaheAxpGPmkA9axsB4i3l
J4dgGsVpjNRPd981aCOFC5dnu3B+QQaTL/j99mgK9sbKBDEnMcfyfme5QRHXAc0L
k2WeO1FBqkS2YZpohHlkdKQGXN40CGDqm2Pt0VRVacy3pXcA7XTNI0Dq8OyFPFuo
uQDKGommumk+2JayTXBKehcmIAFsIpDseaYtmXk+kpPKPA4ZEdIyz1ESkT3TPzTY
+t5/o8PPbbWRz24Yqyr/LlRA2/mbJu+fEKd5fe8LOeoJLKbtl9GRsjB2skwMMD9k
+ttMkeq2tNm99IoQdHl5yyoWpzwCcmuyv47TKQ84MPA=
`protect END_PROTECTED
