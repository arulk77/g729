`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
RQ9GF9qSwauqeWuVIL00JyeYZUWDCfGpxhzZ2ZyeZhY/snhyw2AJmlibVgAd8Ogk
Y5G1gk9UBjvteAnTOkZ500gZkMLr4YKXbHaoypQpQwsXWbL8BW1d/tZcy0TLnjUp
DOqH42TS7Z0Kggc2Ehh7L9IJu03Y6TcSi+DH9i0HWLBNvQmTIhHNlCpOVnCzzRad
AhDogJSQWwCvqRWBysvWjca8kQEIOQrdG7EN7+uHogFmJsLPs6Dnl64rCOt7dokA
VXFYFXFwiaJwagtVeO+qgsIYs1P7nFGDKlyU8jVomQs=
`protect END_PROTECTED
