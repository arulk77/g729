`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
L39LfCw5obIW1IsmmD5gZprOv8s3DPQxWkRGrBakHUZopM1ekzkdHRYQ2K6Hi3rV
kCyebhCFYvhqkkXLVTTyjYPkYpfUB86P24zZGZSYCrEg+w7JKr7aNDZ1Y26EyS5v
6ZIl/ooWFaW06FKZWtJ9qGp+cWmZJMydFplmDrr7l+oG2XN35TcoCglsRDEzOrjN
Uf82CjRSPMjTw1818qYshB9eJtmjrGgsc7p2leuPA68KT6QzFmL0SiNyLcv4jqDk
jDKJN2WuX4oqPr+M/DS0rxo6iP1Kd03a5f790OmQj3FZXPIm4FdAgJE2WCFwZ7TZ
qbfBns/B5ljXh+x4Ay6APcBeFrKxzVTrzESgGTpEr3zNTs5dne20MUoF6ZGhdM7/
I4DaUCwk6TpptiWWw9mo/+gzvnZ6r6O4xKjJ9q+Vblw4DDU3KD5+pDXf5lac1xEU
PyOswSxTNQlQpYQzdSSnqc8vK/9Z0HXTwUd4t7YlTscJQCBwzH7QdoS5yaQ2yMUn
NN2LUS3fNfxfiSff8XhhjFp6E3IGk1ebPzhAM5nMBjz6fbVj2Ks7mXV4VMZ6KEcF
SI/xx8IFLwKHC65IRHwk42ApllpZJrZALiPUm9TuxnieQ2VVUTKoc+O05FdMzAMt
Dw9SMlMOHzsW0QIMv7OHPhqFnQFPtwNFngExRHMAxHlxD96zanmy2v8SgxSyX/ct
+rW7QivzoiNo8Y02yhHrxJ+KiPg02sKpGZ61Uo+0aeCbOEfQKDexetAmB1bgjOXV
s0YjPDkdejdLQ5d9SWJg79T9DZj1po7polD+GMkGp+/wLlZavMOe5rT5AHGTHSqo
`protect END_PROTECTED
