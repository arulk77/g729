`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/6DwMgxXAmRqg+BKZ3uEQ0CpNCyjBGxa43Hsgqi21JW
J957z6wGIidCJgS8kB6qfKMV+N5qiz3VAUXh8hkbmK4z0LKnpttnQg3Wm8TF4Mat
YFwzSuIskKgrT81hphYANMKNIYvKZLkUY0/C+BrTTj124xFoH3UIrABjqQomJoJ+
9p2c++Aq2iv+qYF3caTPeMboc2faYiFiKO21tZznPBasdJzOrGdLWcdNP6mhyVFl
XX40nSxrwRxa8ATxclkdqgBiAeZcdxSKK3JbGrKcYjQ0W23uV9I8pvyfEipy+LZZ
/AwQUx1Cd/PDu1DwDfFsSRZrl/Mv3WO7iUTsvGfm2kQtzuurrWl0Ms2jGJ/Y3IWZ
xTgYXQ+wUr1B6ahEc46hAWbRy9WaBxBEPxX2nTjzeMN2V/DiuyxTs8mXvtchu+ft
ITS4jT6ra/mFCxtvMNBEwlQQoezEVslSRi/IZ/2dNkCfNWyD17r9Sw4taM9zhlY9
tti291Z7W/WtDq+4krsAlO/WLkOp7yuJSwlNny2R80pXHHnJSRDIgIRf12L5yRQQ
yOGhZOoAj/emsJ9GO5crSLHaM1EaxBUXdEjvWSSaYR4WqGA1sdTxXCTXWMeVEF9r
xqdrlrha3xUgr6KsT/Hp2H/IoW5gjf0bqWX5pNWSWzt9z9nTVbOJacDmK3+pEipu
+F/KhNET8bdtWEXzB13sfrANTkMpSedzA7Av7aapbIZfp1oUb6qk91jYE1nvGHVC
vZ4lFdMksLGxj8pwoGEbKHTZmVfPww/aAmdSmHFZf0s69nWMkfneCaikFha26+b+
Qdrhavj6OLjK/5GqHfnexcDdN2WZRctpynolrcdPidvx9lNRvIBNBrktT5WoQ1oU
czVDFKEk168Uql1IgpzMqnFmZTmmrXgX38ZZdrSswECw/Owm71rJwPRaYMUnBAow
31hFvnj+pLnv90b6oGQbK8vFeqSn/plXkSjlGwQviOSkdLpVmdIuKPzz7GFpJvPR
csy2gwrHVVcWcirwYH6/ia06XqiCNf+FHAWr789+guE3b8b/RL9WGMvCEhVlWQLK
cz5/hKG/sKvlMW+t2KZp2JT1m9pqm1gbbhyjWjkvfN/zPCBWDSdDoD5cyIusdrlK
MvdvfNJZO/5jzTCxni7GT/HOnbpwDjLqpUYk2Gl11Aqckm60G0bHEUPQooRXU1Xk
CzcGxXvwH9nyyEpculS/dwAUxfR5vSRL9fyO37WeZgkmetgm4/eWfXNmh0u8wDjj
HYzgVwru01kQu+lLZ1PwCb6SqUdVgx2KePqELsJyq1CnHQumey4bA6bDE8HKlPST
t26jtg3rMS81B2xKpRURQLAa/wq9SOrZ3/8T+OjYDmE9we3C3jPFU3VaMCYF6GSs
5oZJJ/TknhPJh89NZ9gli0cYFmv84BmIx1Ft8WXls4Gvu/me0z/9LKz0XCf4UmUf
mFIkkWDuoDcVx+22UuZuxdWYa5UIWoADI8C4RiyS+0mN7FmPWlgWHr4uCmOig680
G9drhh7Gpq1mOWx5MdVk0DQ9rowOOKrP7KIlhl407yRYnLL0GpoDkXcEXKgn2/OG
TBpeoGVzANlUxDX+iTSbLdg940DqSfAAAgDHbrAEFDtR+21gYhslJeeg0tlPKHb2
RnBk6WlQDuN+63YYw9VK2BzkFtSeqCW6IMXIpjunBU4kN5QQVoxs/sDGNrdl934c
tcYjwaWKIpVQ6J6PYUeTWD/4r4U4xYIPcTzDQKysGGGb1urknk7pGGLM6cLOlndf
dXn2EkIZH4fwM2Yqy9XvlzOOrXV4WD9fgyrm3z9pdEyYgnJWoQk1b4V+p1yrndfL
YmmFzTtxh55IzTPJwPG7uaO3RyJKoGIJYA4Z8vwaX0wt5822JddcE8Rno1OJcjVj
Kat4qKJz20391tYgLwH4RWNsWVhLsHVPD90AqjeAmDmSOKZg58ugqvmjbg4LN7GX
dLB5wH2H9eMNz33ZtopHOk5aajVXrO6zUxPwnTr0m/LloErj1BHwlZ0o9MyHvMeK
QLA3vSP4GSq+pOfYbsCnhsWCrdChjQo3dMXPMCAu10SjbXEVaa88Ql4Il6q0GMRx
bCtww1wko0IP5UFv9C3ksvhhxo7CV9gkUjk+Jp8/GHiKzZ77qPCSq9oLHnyu2zjW
tckH6wthd0LKIfFwZO+6a7XBj/uNOhx8kr/N+XMeaeTJ2bp6GNn8mmrF4dBJdfeJ
u6mH4d3sTGwU5iRI84xZEg6/I6DfwQafrX/zQnevsxc2rNQWoZAKULoHmPU1e7M9
n+DyrkLXtYRHUptoqcsE/WeFwRjKWg/Rb6ZZLhRf1Kcr+XhQG9U6iQb0ZJhTc7B5
VHYqN+RigaRPPqXbD6+gPc9OW7EgQSU+SNYe8kH4/F1oALaTauPTMTp3jR3ijwPx
P1RGkAjbotW6oxipeY/G/SLmdFLVEUbyGvemccigE7Fdq0hIXpnAzb9ueaVwQZml
+qu6rnw1ccuR37vavCFSfA3IDUgwtR+9SgcEZYuVjNpVVPcDZ+Aede3j6GHmOfp4
8jLtuGoIw9Os+zdtDtKQZAZZ7LWGklLfOAYBZBXAP7O7cqZQXY+ZDwbo/sgEg0Nc
sFUCxK7377YiKOEqNu2PHkqj0bB3oYF3cFnD6HTa5JKAsog3hRmRv7a170Sb729m
zFmYWXr+nESzXRF+DG/Km/jOox0/XCoywm49K0PYuStfxXk6bRACuYqnMUvtsiFN
LxXBTtoUZjTMzJQ2p663pzPtsiMgIojukLS2gGqQtmMPcQswyqoNwgsE1ydnCV/M
2e1WOFwDvpABeBW1wCXZLgM4BOA2ZlJYg0f2sxlGhH4j5+GdVydCryTMh23ZYtJN
DxM3aYVgmuqzjTK5QSiHPs6QUI7JIoFQSOWFA0bn00xbGh4D0DeX5GbasaI4Z0WO
dmjIji7NE04QFeim8Tygaa2TQlqY8ZKq2OC/Lj+K+iDTihUoAc6FyhY4pKpTnUqD
+MPPE2jtaFtedKuWETOsDZ8kysNxAxEmvZcHs/4HldaDzxGnq4AqpdysZ9OmY1M0
IYxhDme/PtURxjGZ7DzREjkJJ0LhYap34m6mql0qO8osg3F4BeUjGKUiFgEFUzEU
EXE1tIr8yV/TYWkzWEIm2dXNGT/FotoSVKl8ucX+eqYzV8pTnxPfITKYgjCUss7m
GTFDTNf3uhs6c7WHyKVPoiI/lqZ+/W1FBYMD+ocgZWxPga+b5ZC2TK4wO3dSUWTs
q8ZeDtlGL891kF561bCyld7E+DLoJtZiizn1OKbytTFJ0DCm+muJ7m89/YzeqLnB
Kof62AHzvRIx1GgJ6yOXaIcLV0M70d0vWDN7VXojPbUmmrag+9dHfohtXcxGSGfK
M5Lb1WxM83T2qa+AMLDcoIw4XJaGCekFXvfIDJzLL3TEsCuzOr4Dm0BMOHlzchi3
YE20SFE//TqNPgpjDywGwg8B/yZ9g0dFtIbWTgso4zoRXfe1v5m73jE6z0e9nbvX
/bJujk8+afyXW5cIMSD9Fz4Y7CZrjOx8WtY8+on+CcFXmvfmc90H8R8tsk9BRx+L
PqA8GJDH8LTUchFEf4MD2RRv4L1+ZbyjEcp9UHqBGGwKL/PBQsi7Gvqcq40StfRT
WbZkHpnKrh4UhnAJxbrzanihAYffydhCVuDQhGjgWAzVcBoy1oFveCqDXFPbZP+h
gdGb+XQ4eNkuWX2jNSm0mztycVBYfOFeTAWDld2hgk/mE+GsaJ37LeG6HfFXsDIx
7fA3P8AE07dnEWXy61tYBd6R2O8y4y/be8dNIHCAUEy83gbYP3ptxtiBCw/elVD3
NVP2OeNK0NnwdqRGGOCjcygVHVwsT8b9+WEcKESL2AM+0x7z/rEcPXQrmWiJ2YqC
ywBQlTBcXx2xwnFRccuJh7O1bsXcSZLRHqbv3Ze8O16xJCSDbeMKMpfhfcdPrMuo
jfIG8fJ28x53HaFYt4OOP5Zcvo32GR25IQ9JAXBP8U9p+CdF7Jyy2azqcD5rbqcK
1TttbVNgM1bTsu7nY4cVBt7vnVX829Iie/XyrsJc4gYSzwWShvszM2HZ1Faxyo07
CvunB+4pl2ekSZBNPRt/6hBO8uv8qKWXvZT2Xm3DD5n4YFUPW0J3nAK1mBePCSl2
80TIxv8e4pqgCl4n/Su0cH1fCSagn0wIiGYQxZAjeQw3sJWvXcurJUAGF1Dt7RBd
RHFyTwZ3sSdXEqLtKsYWRc3I0A99MT6bXrFAbDc9+odx4e4s9GWX5WPaUqVRVHNf
IFODttroqDgRm8UHenOqs7AHxRSyK8u4QjZBA8XRjtLIoaeKIV9Lhu8RjrUIxpTZ
67WQUqDOOSRt1BSeeT+HTTCLMEms9Rh8WE9iIywyps7lFnJUyM2zKugDvDFFDKiY
vJNVtQYM8eJsgPLSdNU+D7zmH1uV1avtX0ZdfyEmXlfuvEn7CRPlJ8Pv6tdaUTL6
gBvlqGwWJg5UyXPH8AtvIP+TdogSCR3o+jHgH+UgJ15Avp9tBiRNE42+8D1Fh8+A
oNsVh2ixW0Ixz/qepQN/vsw1w2DdjP0UlbWPUoS9SOxjK/KqKZ7nexJ44FpUYTu7
9svd7vLkz9gVDisksPwpBSmW0Q18q8vvnqi3O+AJVzprttPRWAf+HgH0dMH7hWe6
33km368WKnsPmIyBvGFKP/jLlK33ni0o/o3CtHngRR6lCoT0zFYaOUchhsmdd08r
IJn5EKre9XEbkjh9xD4eKqfdb5KAKviQqvcEOR/06fZvgGiq5X+8fCWf56yRzfRo
ORs/gQonNKTpdCKni/F5VSHvOTL2ee74TF1RvibkUR5uNEHN4YtzkrH01Zlf9D6w
iOYKxqqp+fcWl+NYdukHRMpYzlaovH977uxN9dJVYWH8EPkqSEW+xPw+yUzDP5Kn
HMcvppPOu1mdDlMncOzhQEncyeExiRKCchUK1V2EdRoynEtQxPtNaVORUULSrWGa
Er4M8HcbR3QJNj+VuMpywiFI2of6EQT+yR/bGrUHJ/eQDysHPRMrA32gwXoRwEBS
7Vqco/S20Puikf5nTZNp+ti8GUHQknzO4WFAQsVOlnJDcFImJE7zoTzBOVMJAxJc
HnjKvWjUTDBN1Frsxnx5AAyK4tGqIG/L2qRgcxZLHEk/mODfSmS5jZBMvc144ECg
q0yXfwoPdRPrFjp5wN58wgmi1cRCPERJ9p4Fzj9ZK1GAtBENwFyguPEbpqG+A1Zp
K3TPJ5jEgLgeiryq77LiRuMMxu3GrMpKnwLzofs4dE8Gpb3SGXubHY/Qv5N49FYP
oA7oh+RhVQn4a/IaD0Xe5Zg8lB0u5+7fhBtvMuHaD/zMK1LVhbPLSH/25VRRzsIM
j7fn+0mEu5IxcijUgfETqWjc4c+ZrtzqFBg3gTq4lgiV+osU+/VRPrrazPb2gFlC
g55yUnGkW+apo7JrqDBUgS3t2d6y+tU8quOcdqKy1Liq4yHUa7ftwXASMltTa+1S
JLua9MAFiwL0OueU2I5YELqDWScbcrg5Pf3zLnqP10p2WpJh8ZDjQDVMjTGqN/Rp
VMHoy59osYB8PIYYDY+qNZLCup2BhZAYCNzjBASJv/Z5+KDxcksvfpB/wyD2Cc3u
ctvY47HHTEdax2HZ1fHMRGPAMjRqdnPWgZ9PD7j4ZwPdLTKfef3BllTgzK+c5t/C
kpedW+QrRE6qkc6UmKMGHbr6l8aPfEtlnXXk4PztlKtgvSQgdYyPEkx2LwBUnVEC
0obiEkWLrj5+cPvhpNnsWI4LTrOCSt6mJXPBCgBYDrd1s32AXHHXUd2vwlGjiOOY
ltapwtPX16oMl+lcADQPKpYsE/SXtYv+zSTcRaQ2DW2pfp/mFHTH0fnlQQJTJ8dn
GNgnvtCK8EIXRTvjWH+52A77fg4fJ+9JBE8q9CV3zlwcAQ0oXOmob5tIXXQ15eao
MnMTIvUEsNmv5IMFJyuPiDGZLVxpfnndEKRbtkhd1d46mrBkMJbFIC6FSjgaWK81
9u8Sro3o1Bg85Jj+9JnNmr69haxxIljwZ/60+lGUMA0FEYSBmLsXaoG56flJuyYS
wqkLfpSxDxHN762NgJel7+rDocC64QvjNnTwEcjZMDtKXBTjtv+rRsvIXm6lTj7z
iz6bjxaca1foRnDQzkpGojxgFJfpLNK+qDol1MLBRVlgy/JomD9aLDRR0lvO5JfD
GVMHVL99sNxu4P1DaSziZH6X9c0cgDhivVAwsw3+VR2vEYvI+9t3Cfa0djAYdOEF
Wod8ENLdWM3hqWgBAjpac0Qclfmd7gPmnkCs73uMWLHZZFMuCJOTkQUzQABniYCd
aeT33dnIo5JahaKo5RFxJnjIe+HgR6cl2HoKsTuViRwXaWf0HNU2TR/uCAe/Io9f
Vj+GFDB1RiPmqCIBjQVuJH3JoCr9cXThri1oEmDVTcsgrO0bh8jml13IWHX5DwJD
IoMEmZRykWnR8ugqiTY+5X2jIFG8LlMZxN7FeRnRGWi8fxWIDXGeiA0jnPehfP1F
YBie8CpZ1yZi6YbIfOqVJl0zTsrYBGWIzObffIRcx9XobFU5m5yWC9zCDlBVKEu+
XY+HSB9ZejVuBAC6hCHDnbeZghID5ruWd9JeVOr0THK/XTaSNySFpSRo2+mS9o1j
/F6Fw8DLiJSTaTVR9+o/jtDUzhom4jNWT2a5dnqy6UdnvNBa9A0WL14fshFAyvoY
xxNRif9oRzYDeOkq8yj4XVHviKUyGfRCXqplUr2ogenUg4Nn7A9BKlgMeBkJWbYl
54M07Q/aWgpTOFtXYltUuEbIrYfCHGc6MDs8xYVUeTXrvdoet4yBHAlfNzSu1MDC
e0cN5w78IY5piQM8M3LjKAPmhAksDDMUWLhCCK7g3BBGII/Ig4jcadAkxurXUfYE
ialgZ/PPqn26XKFAs2KWyZ8s/16+Z7axJopDf0eYhQ3BIGAprAhEzrLjzu00UdTG
rDMf6WOOtlvk8ZSfVSfrjWTt+v9RWulym5/xJXcdRcsNRYjh89WZM1itGg2WWk7G
OeR4FAkTsX+ikE/bWjStBnYfZsf6Ncwd5hD6QTL6ZjAURt3xkgc5+W2tKoPBuzYz
dyI1CPf9N1Ek6ydsZ2t/hzVYDeo1gi+MeOObgIvwlCh5gD0eDUgfmsU9EqiLdOgi
+XDiTZNvKykmtOMXxviOFvQPMwqH9kTEqfXDnorM95IUSBHSJQyc5Bz3SFxwHbdc
zv4TgVyxlUWw0s+o3XpwLvft3LaOPqaYhZf2Ex9tehPiKMWsAusWs7bcpQpujiWG
oDxPDEsLPQvLxKzsE6GimlvRlDAxcZeD4wqU+DCJAO5EE8rNE8hfMpuAuYDB6CiX
J8FGboyk3qv8chEwG48HPg9g2kQAwHAf+xpg+VMOxtA/QvehTeXg7z46X116Xecj
mpr8ia0UauFZnXhv3uLD2Fr62uj9O1VjnuQb6xkAdIPoukPSalnick7/z94CQWuS
g16vFBxP4PRnIwdL7pWMLNB/+PHfb7rhWXYRzedm8nN7jDrflAeDTmFgWDgl428y
4m8BthaRwxNLBvm78bsnLoiWtUVOjqT6uoIb+3YK9TOYZW6LxJ1SC3Bb8R7rJ7Yi
y/5lFzHeGz/BkK9YfRHx1kacBeo82lJx5GZDafSkudLJFoxlPWPcRpvEpNV+tJDN
NRnazdUIx+KHFGQ0+KwJk5qmoqdQoBIpMWpjOBSUKyvqLhdX8fffJZOuxlnaU6qt
hQox2u2eEmwof0JXhwFK59GMQU6reI9t3zdEcbN4qSCBZEfCJgFarDF1WNDr6rDO
Fpigw6sxSK2rMIZuXZ1YW6ij191kmOnXuzgkRQl1dkSbhXm82bS2AJfAelZ68G5d
M7OzlR5a0+r4Q4lDqI5WyN6S9Q7eIeyNBc0hLQWOwAT22MlNKBgt0cNQqJMGMA5D
lOfL37ppnOKspek9/IGXRZSLyOE+IEF6U6WM92zfd0e0hntljiUWYGTS/+6dueJN
iGZ5favp5293rcSSl5g8rrG86N3MOY6hC0RSnhAd0OMEmtz8ZvDTkrRcwb7AC9Fa
jBmrvQ29LY5ieFDryadNdt+yR0ot5PJvnkcEE+bPZcNPZyLMSuBd+yIoerPOUvlV
oapTWA+WEz6ASBKaQhriegUTqmcsnBW56kCgBXA92tHbFmQU9VeSNEJXt9NjllJl
1VUyowRhiUxi87mVv7dr341oXsmhnCZsRZsF026bh6vx/RxUwNU5oCxjjw+kO+ki
sZrNYC2pSVhxAGoZNYo2eg==
`protect END_PROTECTED
