`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SRv8Pj04gmsBlh5llkACc+sFXjA9pdx7QkNALCM3kWvM
jrjyGZD7iQ/4TiTd9QcOj4Jx6L/2k5C+znbJn1du1J4v7fPHjh7Y2NkOExGKALjd
+SUlybZSLsXkSjaS5YOwef7Tw+NxYR0C+cBJ4UBsUfo8jc2AlQ30mn1sp93nTTBj
yQfJhUPGX4YjAG2sz/l33C8HfhDbdNen/icwxWuCRpekivv6kBAJkeMHt97qJlAy
VGctqBQuaa/HrRqOpLo+s/SU4gQ7pewOHs5gvdZZe/vlxdbXOudL7oQ/CIeeXCCD
KRRz5OI8ZJ3lzK8/hXVDBBQi917WTyNuepa5Q+E/JD2o4AeRPU2T35Ij0QdQfAfF
`protect END_PROTECTED
