`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
VBAJKddLhiisED9ExTIkw0lS++dpDsHy2oB+y/5R5i1IaH7YXQFkYCfTwHskBk7J
ErNIj6ZzmUwnXwkQSgu7j+3zgN4KAsI3Qb6tb7CUG8kumpbSJIrRGZTxL+lqr895
a3a+fxDeT0X5ZrVi44HHjG5iLIXn6ElkwnleQ0x0ELPUhbSL6sT/ka1aZvuBHRNM
9dIg+B03sWpuFYXC//sf3NRoqtpqPcZEEhEyuV4A9g6ExHtMcpeIFWwpSdpzsv7t
JqB4q+QTmCAEDYj7KIWwuNb7GirB6K7WkH8tfsFZAN2vaxMgxdrYRS86M9vp7fwH
`protect END_PROTECTED
