`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNX0ypKmsg1JZVIKwFXo5+64wcTRUXKE9UtQcfLwQqQh
CN5dz1nmiPw9YwqXNXLofmG1tEyEJRNIv6JX9USpVJE8CnDfWVLqUDFSQR4sPPnf
9h77UT4h3qUvcXhEbGQw5wBG2IFzWco4sNju/gWTzjO+lkxgYHkH039wHSEJn6k0
ZmJgGbCvTUYuzieOMl+uBSS03ZRpKHwD8/OEZtfhvvb33YkjDOWKy89U8EjQGiKP
iM0N5n6EIOdlpv43vKBsNFh+c26QoHtX2IhykIxG++FvIs4Vhlc6zUnG3KerUf0S
tmjXNWwwzye84NZoxSpk1mKrHYjruxNTzy8TsxslO/YX54MFQtYaSOJGcKDxOs07
jMhg+zbwRxpQuJP9r1+v7wO5UehGM01YTF6maSjiLKFaPHzE5QpQN4NrcT0zdYZV
I0++gKco0f973IOxabQOUp1kLd+WwM4oHtaPZrIb/nLhhaUEguP8trvVC83cO06U
3ZfvQdsPkwDdAu466PnhYKpmgF3R6cQI5ZI1Wks2r8B3Ade0V/bNdUS536QMakW4
fzfsL7YqbFQ6KW26lwAs/a4qmdn6F0p5fbMjOUiMzzVOAqZspCSkKD8xZXDgLi9H
1ILBO3265rkIQ4Hlmjv9PDZizzwL7KFTE7PewiDll2AbEzGVZQ9fFFU2EPLGkw7k
DcmONM2OsHPVrVZcI3VOGy3om1Zeo0fJyI1ZV16xGm3Gycqui39ZfpILXWY2+cOV
ZhzTEWrhL83ZByUdpSIaBiOk9f11+YP5NuS4akG12bg=
`protect END_PROTECTED
