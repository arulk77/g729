`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
BOqNFHidh7FGngcmIunI1Gx3SMqt65zjJdhmDLzxQYTV8c5Lo4RTuiBC5fwktH2f
sCRSI21bY+Xmnt7M+pQASHM+mvgjbcl9T47QcFbsaH1vAMGhjxAyv0Pkgn9eUA+F
p4OzWrt53dJp/jCHUKr+9IpeyVIwta+133tfQsLq7cCPHlYPIvrUzu82n7FoZZYK
aBeDnfBXuF/NfjRStX6YHLDy+sayAb3aBAuFory8pP3U+J8Z3qzkBiKNDvEaLTe5
`protect END_PROTECTED
