`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Prgb+lMGK4ankHVaNnLDq9rn1TgS7t1OSsPkM/mjX1yqUu8Q04PjYHoRo6yNbAMC
9NUKTNrs+UQ4klWfcJNmP+hZbvTrD0ASb/DBINgz8lRwCXhNV6BHD6lojyvkVtnl
164hE+9eSn3ZYmO8q0QTCl7wlActZA+3fJYRUF0ZqlyWYSlHPwssNApb6DOb/xoN
fQeCXgy/Fsh5eQ7XA1fCyuxXwd9EO6jJocIlJVpNbqGwQjeM4qiy+B7Ix8unrffq
ZarjE7K1+gZl/9ElEDb6IxuHRsMXl0DuyVqUoQdwvSkXTFkLL9RJ0QARF8OdgXzG
pRYxIX46duo85w8GlQsQn1xtGrx5A+G6q/+Uro4GQJsA6k/2qDeJ8tI7Tf+M4d5R
KeAHsFg70lMi0Dt40CuT/4nzgHZhbaRZazDX4shVt5A=
`protect END_PROTECTED
