`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
if7OW3neLerq5QTb0GME98fz/Jw2t4nUfE4Tz/FMevN8ZPOEEAhB5tCOc4dKd8mg
Okm8xwopCzd6kQC5HYb+1ZlsdlLgAeKVOpNCnF0CvodWm5jb1PA8r/W6WopxdrP9
S15Kdx4am4SFTK0uUEpAj+Ii42y4w4L5hJ0Q02b4AfIS4gR26Pv9BwGpR4w6N0yq
6OIgAZdGfsOn9L7J77tmKnMUzEHB06qv+6rBKJzKbHFdodqdnc3SeuAJUu9k8wdB
P/Fhg8D3SkN73PLJvJkDJ/2c1eGVnwweRxRv1VOUgXQ4OQSOGioHV3wXIB9SbHci
`protect END_PROTECTED
