`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
rdGd5HHhlJAbkK7inYyh908ys5MXzCLrZptm3m//aJT+RsVlpCNVhVrbtxxSvdjJ
6ofFyTh/5E7QPJZfHPPIsvkE3+cdPdMDhXvo/JC/gGCwxkCqZvVlGzohDqHzUIi2
AwDaqZ4Xzv89wxGOJjFekq19yV/IgTM0urrP2Qrw+IoqPVLV81acjrFZNANTBP5W
+07iKX8ayb3dO93rZ/a1tj/7CFmQuDTwTjcZQjYaUEUL229coIVGPVC+jAT4RdTq
fWQR3YMwHPLq4Mntbq8/BZ0xItBbhykKwo5r2ulDsSTmS50FLhIcZE8TzTcPgWe2
ECzsl6IEuCbp4h2KSjKm50HZBVeX7yR1IbZDHoDYoqTI8EgwTXANeb3qjgnRrdhQ
t+4+Yo63pPbJaMr2B1+uuq/2TecF10OyiZuEK6oMQ5E=
`protect END_PROTECTED
