`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDj/rqtYZNi7Ql6P9i7f0dK3XNfOsBWD9M36eZDGErub
j44sQLpCRqLYQKiKn2+4f24LqFlsRYUPkMj7MTDNk6tnDb2nLfcx1F1m8Dy5ij84
utRnAuftusBkOIIZol//OBkuxUfNrVWyBG8S7vhcSc6uUjG/7xNNaO7HHd15QN+T
PVpxjvl6CwJilnkjoDJqFLvE11HYmZep6kgfECbD42xnrSRpvl0CXR55N8IfXgqS
8L5h5/1F6RjbdxWDOWdPcKzyo0CNdg7zp2P96arb/NgQNNQVOlukui0r6m20Ma0h
+fEUbSEGyK4nEk4bEZobACjiXr6ST2wRirsroERSDYlycymFpiTOdxYDwU6m7ph7
`protect END_PROTECTED
