`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveITLjAR/QBUJZ42U9Fz5hNgI5YqURzI0cvCOGxkf6FFw
r4CZj/PUPHGxpSx5jtiZBuyQc0bz38lr2Rt7I5vVfL9rrj4Mg3tZqXcgjqAhO/jx
S2j+cRfUWptMEIqg3Qm7tt8y89hkQvGfq8qWeHSxAOZy6Nxff+VaV9UvVhNeYTl7
bfmU2Z7Du211cV/8+dNlvR51ReUpqdvfRHfwa43NKrEcJ23KSoRP3SUU9ap4us3e
B62YOUmOF9EcDmwLLHbUIs/3Om/aNfhIb8AncJxD81P1+j8HmTLpV5XNxdWSkF0K
xYLZqDhMG2qxUZXTWnGtpV2nj3TRWejm7kFS6ot/YNOsrdwQJWjrRnB+wb2K1Las
XZJPJ1YArO/JOEaCsKQ2QvA3C247SwCqNXe35WhO/gtK/KvRNmOafBeCxRgIucdg
tCiwXoSB9kiePEWZWEhbikEOz840oqRuyvlC/TGRg2oJ5EE99TpAyoTj/lGZwAZ8
kfKrlg+J86zkYsDYnQ4ZE1e/yTyymkhRaaScRr+7MncHDM1Xla5DkvVUx6xr7HGc
QRqib/zCtjaAJ7iLCNJi/TsK5zs/zfomAQPhjGrR1nNxZD3yBW60xX2QscyUnsSw
0C2ypzJfH2HfLmyrwarpfpQmqOJI7RPf8RLztDmhR83xfiLThrS4cEPWBAzd01iY
`protect END_PROTECTED
