`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMUlAIikyRwsKWLroZi++IlcS/nxZgv2JGodcLA1mj4w
0lb1Jnvegvhtp8ZCapgy6KJw0FFfkanmrwd+XbX1JJRw7UoIPLh/Z+1vXrXwLu/u
CMGiOk6bH0Rmk2gayAUFFd2Q/hjzr+C4LHH6cvHrc++xhokCE0B2UCnRoQC9Q9vg
oi6YIUSjKCnsrMvh3JZkOR4GKafGwpaq1mfeeZKDJWCtwULBgrsMXYQwB3fzLFOG
Z9yW9pvhePZIT3VC4BrtuwOoc1dkY3UcUKPdDXbNLYEo6sh+ijPD8SuBq2bl2x2M
g4DeVJUPQyjiw+83GNDFnJMrlsYW0p3wMmQuzxvbpUTaynsBWo8y+075Mp9FLtSf
`protect END_PROTECTED
