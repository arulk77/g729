`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNKSg3t9AYoiRscYbIUU1c+FWH9cB8ktb9V4+OTrSe8o
rrOwFobUlqnvawTbR9iCGzW8B2zJhAIUhawgvcilZUGPJqDkzzo590NZrfR5fVeN
xGbMThN+dB8PBpqUGC/ZbdSPdXgoeeg1ev/QeNW2AVyNb0h+O3bZVdk1ZqdtCGqT
/aAhVkSrgiJQMgyruqowddWZY00IPuM1+1pWDkfyKm9/hBH4d9NnaqhWAL6uJJKT
H3BbWnx9qeTSlQuavnbbBMXYp8hrkoZZGIaLjBT6qKlpLIgNqaTUAXz1xpg7fP7s
bwt0LTVsVDANy3kgAWt0vXSSSBrnnJLlLHIzD4vrWPWysqjpS6B5htRGChthQWq0
EMrI2quJtNCVn2GDK/OCvW9ossZyTtB9R3C5kwOuynThNg1HcA2l5chBc9dxUqzi
Q/PalLrGH6l116ceiBzoibnA6KgSVQMoDS9SpEEiVAVMEq5VDv29TfpM/jbZo/Oe
BThdJ5LMpfbLrEywKw9Gqioto6b0HLEuTfAdp+eiQJxMphZPkr4+TX6mvf+SVhf8
INXIIYJNmRAM3H8VTmHQdw==
`protect END_PROTECTED
