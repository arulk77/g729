`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBTxhhZ+Tpx5I5m8j7ODNeSEDyKyZwxr8HnXGNTLLrWN
Ex3MzKzm409IY6ZH6eOGVoWFLV14f0R2idodsTcb0fT4g9PCaxVIWODHVAaWre3h
MADNSF5m8B1HEejA22aIUwp+4XBn/gKFDDxrgwgR1OFpf95/Mxi+dKBmy3Ipu1gm
pw0WzpbdHfT2FMNJ1SVfrtDtVLbFNRnwQTp+qiOxHMAe2+tcxjv8/zZsDmNxo4F5
GmLmD8N2D6VMRLxDofT5WZDVfpjalIEa3kWW4TGwFgloZRtcLxR5fZ2i2CjHTox7
/4WoejKU3+a+EZNxq2rGjDcQp1CcyvEm5sHkAWKBr/16cyJBv0N+X/k1W9FPK9N6
2jKzsg14mx73Q9f3QQKO8vNKOLNrrpVe+YmzFMh037K5Y2A76LbLEPbiy3Yw0uAv
2uwO/cJmucJdrZpsQ/yMh/2cKrc82qR12ghnyb0J0UjNW0nKIND6pkXF9aYif/fv
rSDK1R6cuCH4hrjdSawv2/EfVfAgL+SIGEepW2YW/wtq4WmF4wOFWwOMiTS6Suy1
`protect END_PROTECTED
