`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAfFjyaMm8AowJqrkmqFVIwfT2Tzz5RlFVE1rlsSgMaUq
zb65muFBz+GKuFwZl3ruwyDZDksSOjV4eA7QAFGBlt9VWxN3mPp4e5fExusbeZx0
HnE/7ohxg1nA7BGMlEqqdsYo/++VuUWcarHnKreFb2QFDJ5eC5sd+svnkv0KiWNX
/UwxBzuvzRJk+OV05utvVXWZe+CzDcC1FgLbquohQ025bMHvpRkgqxql4EMiRkAY
z+VrsykVZFD9QuhjGfgMd+/RmyuyvngWDmEcL9lA1RsrD2HWmL3d7+kvSFsDtrE0
6+TTbp/jMzqs93ouJ/bnjcN9LztGUw6o9H7yUZsjY23LimlQ+iFf3k9uWYdlBZ0j
bf2g9bpfzMFGEJb95Bl0MfriNs/VA/iCY3f5NpofKu9XyITc/OCG14ngf0LoQEzU
5pUOu38j+WZZr0ZZKHz+J+esZIlUw0OhYDbbZppjp3sl/SzICNt2nDvRLeUVK1LR
AdBDzkBcm/2ED/ihm838/RzPnjfncEjEdnWKaQbveFiBJJ802CZm7+RHnZGvvcNr
ik8488oHwtQ6AZzE9TjxVk6cIqlsInOU1p8eJdILhFtAKN0zqQoPNNzkJD56WgIw
mkM5P6sy1Z+6aUy8zaln6BrlmgjehjGcsi63Vqb+nnmcVImIHEyv7DcusuqxVK8t
ZKi3GlFnvV1ubOU7500p5VYuB5Ckkuf6232EssXn/T+Vhel9TElEAvi/xnFo68gY
veTV4m4XOoPkwzjXz3QdYUeTC5SVxXmde2Fh/1p2pKDqkN/k8TpjYNZDrjEFZW6g
Iq4mCsj+Gj94aCp5IpVfHfCVoFLqlCfHf+kACP20X7y3SLMM9BWEkDpz1PSxpZIH
55+3dGk+HE8UKYtpFl+SJMleMDG793uUZyGJNKF2eaYsG42f01h/oh/zrJYdssix
Ziugs0KOpYjLKmcYQLGHw6/46EkqIqCnSWn5uOjKZC54QScHS5rZLVVRxyziyF0m
KmbFDo4zVsc5kVlzpQz4U4817Jv15ubF8IRlC3XNFUO7y6l6L9xyUXpzpyPYCBbe
r62q6OUF4QZx1qs6uBbTmlDHWKLnVLjyuQBjyK1TMyVR+VklmRoCxnm0Wi0VMrgE
trFZmPCy9MxD5XCFbP4SQ0JnHhJRpo0yvY+/AOMARU3mOHYDfcgYNfRQ3zRtRalD
ahJryatSO/YtsW4AWMAjTOs1VzsfOk2xW26IWuPQ6XMieOHpLVPfDpkDCf26yuwh
lHYvfT7NT1s5U4lTuKNVs/UoPTJ8UB1G+KFlcn7lTE0Lw3wGbPF0O9L5IWKlgHlV
`protect END_PROTECTED
