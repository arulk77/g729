`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4ztD2HyPrWapqWgnpjFp4NKhFFn4j9Bc1kR/3nigQjeQ
PbkcCOWl0fAqYQI/pxHCsmSL9brJgL7IfhY6gHmrZl4gZUMsoIRLBhq9+oRQv8w4
6JxyxT+grqvu7u1XPTdPkwU9o6GBcG63zCttwGNYSsBtaUiS6YLdUbfaeimdvk5N
kKf8bNIhq8BL7HXbMHFgBv+ScgyVZ3PH61B1Qpxmykmn7Q47UOn6poKYVKu73Ys8
3rWlDtObB+kNcpzB95DYRTcCuhxMOCZsnZidTSb1qFw=
`protect END_PROTECTED
