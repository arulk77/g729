`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zWxu2ApZcYKf4wkn7bOf3yDL9vfDRjHvegzdOZ8AFt9
zicZxicyDusmt4SJBheubUhEHgijXw0hlK7nlD/wpS6Il8cLJybsxNfEGb5m1ijF
EmPyvbRKPnpsD6PO/JavNpdbhqzA7A53uGPgxPxzQTsAE6S2ifXCy6TmdQiE9nyY
SPT/8mFkCdu8MdWYhicSwt9Y6t4IHbOUfqscv8eD8MtV5/hf4D9hEUUnheeD5ni7
eUjKU16QeihmyaSDrmlu/Gp5i9YL4N+bul8K40DARqSyDZTJpjjZtV714XXyUWan
7jQnS3WMFyogqI/tKQlR7/XeQeYD96hzZA4KHMZlbjoC+2RSUimcPUj9KO0rOQw+
YbwFj7N/EaA3lj2golSwpNp10VFLTDrQtd9XXVY2OHNC3VJz8h038XjuOMWMpPdR
VIA20VueIJmktru0w7ZRVmp2XO7wjLZQ3l5kbGuiOaEJ+UnvhgQVRw2wx2MnhI6u
`protect END_PROTECTED
