`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOo+C7xHf7yhG0lxvlw9sHHd4lZJHoHB8eaM+7XyXATE
iO/OHq13xnkX60JKIBFyIPm9GSTJfxbE3tr8/9QAZK6UlEM1tVkUNWt/UWAzNYnw
HKTsyYBQfodMISK1oz8rrNYFwElNlwuRz8zo6Ws2EZeKW4CeNXXo9BdylXF5tobc
QEX0rBJ42yWrIFGk3FMGCmslMtHRx0HF9r5VPcVmiSxcgY3yFqgrAkfMTauacCTK
dEEPvWcVE5xsyt7AvUdnxWeipz5a+8E/5bnn5X190BjLWFrA7lyXWVD3qC1/Rs9h
+SKR0q8/haJTMLMCkZYwCo227tI1MmyH8LrcG9SYWhJW2/LzQSTMuwctoBA5Mqnm
jFhkmt7UUpRsk0xU+JFqoIl1oXBsHjIm4JTT/70dvxJrWZ5ZN0sF+dCEVpX6BrMV
TawhvzwFmk0Bc/IARv27jN6NirZ88bPyo2mEC0upRrMB6Z9fDzYJaqRghUmfxdkS
`protect END_PROTECTED
