`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
yvvxaAWRNptbE17J40JecPtQN/w6Y8H8H8JO0FWnNM59ISdd78rUak+UaD59gDPS
TK2Fb2aFbh93YOweXRnVaRyQonp4pv8dsQMdq8jJx8/GsO9+1xIqm/9gTd9alC/I
17vsd6EIDcDy3vcAXIzF+9YemrytCONm2d+EggL2+AWvJFXem8wGRwU4DbpiE/7z
/Wo+W2dQLlZEU/lpJ0vyChnVQKKmLcnWRdXXORXJagCK4EXD3watoxGjHgjgx6Dh
C/+fyCZWkxl2jZ/9+BmORzaopMOK2M/5jZCILWyDtbc=
`protect END_PROTECTED
