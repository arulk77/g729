`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
FUVq/jfLnDC6Jn/xKfOOK5Q0u6T2xctjaSCt/94/0c527sETnUe+Tjb597bwCpcb
+wNenrcui5ypuVp16KucKtKzqPt5OCwUjSp4A1M8gsH9xJHwZpE99LqiJBb+NAnr
z5TfPYIME0NpnWI1/vp1syDD48kfSozaAWW7kgOtt5mPRqKWb//LxM/m8JxE6H6j
jhGRwjrHRtxht3XMCUTo6Pbul4xdcTDoXcVmgztcbICubiv9gHwLod7WlQ4qikui
ePeNNle7VxHgjAyv6p0Is4pX6y7czBDsICy2m65117JafiIX60v+W+Ik97t+tpmg
Z04UsttsnHp5Qh5KAGuO7ddLMQcDco/ovf6GYCpyzc/NpfH04tRoPSLSgyQm9pQm
n+qndj3igrkxLRZHsBWqWt0ynABRxeppAKWNsyT3G04e+mvDuzk8U408ANxHEiz8
7RB5EluhJgu3rTe9WFXkz9XqcCBcgOcvuuEFwvmpZSPUjQBhCVGnNJGjiUJ9Qnlj
oV+3WogaCONejdJ7+VEJ4vN5CiUZYcjLCZx788u124m10n9sbnvfeTM+MY6Il2NX
L4ueTEsH/DmBejlLrl6SpA==
`protect END_PROTECTED
