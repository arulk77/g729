`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLc2g2n7cRNiSha16+tM8lJfRwb4djvF6UxGacPxvsWJ
92NFDrW+D/Zh4fXvI9B5v51VEQArCOGE+JhDqf/UXyVTKB9IP4UpIDC54HUanlaC
mQo/kVgG79kJHtHS12cMwWdsP2/7sY6mkoL0x74wldeErlpsFg7y8Nfo8emoUo9G
GkOizGge/09G4uzK7wE3mg3/EVrbLk8736zgj5lnveQ83FDjiyZTeqK0XX4wVhfG
zz5gsLTLcc1tRu34tlIDVN/b/bmJOLC4zhuNlQSjkmcxMJcqPIercVqYiQA0EzYX
x8hH0bG+BFI6gDEqDKhcMw==
`protect END_PROTECTED
