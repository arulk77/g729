`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJMNvdt3k3+nC62XGnHY1qSyVwqIKNpmc0KKcsmgECmy
8cpMaJlVh4HBzSgDNyKqCoFfDSVY/p7RFCtNlr3MVXTOSoZNzgFWWW1ER1Rl7ED2
QVYEbZqdUbWWJ2O9CyFD8ys2ji5CsgcrYkuUIQT979oFf5RhlOXpFeC1mqdtPbGT
zBBSKgreU37mMrv7Ner871IdGDJeuzzdjHN02TgIWgqyYTFV70OmKcpTWo9kIuxk
`protect END_PROTECTED
