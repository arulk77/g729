`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aSenHnro3Lxu7OCuh5VNCNrwaTXE7ZD6BpVv+eNwlERZ
YIsIU7pmqYgLkW6J6pFfP0vCn6oXp8ho1LWeFhxG/v8cPfFznOlgndL2v/7pORXM
ETYWkbi0aBQZEHRLH2S2dgY8jXYMs2jKxU10EcyiMiQSlhNdYdJ1oDVBrNhtmgf5
XgnrK9mih76KA8W/r3I/mSdsOFPOibrZpEKUdzR+sQLCc6/0MAvUPdntdp47Rl+q
RT7PE8vNKw0CdH0hfpHkNQ2+SLr9P+UaKksBOto1e3d/Fm/nD49G+FCKPpMQE7Gu
q+LxLuIcSvXzft6q1e5DUtxTdOylg0kXOEzCdP6GvasjJORJ5EdjTY5K1NpQs1zq
nbeZE65QfHl0SKyrpbfFihIRlSuXzkh6BbE5GP0emXwnADdDbhJMrhtsRn6AOAgh
9DmQoxKVPSjJ3htjKH0zbt5M4GYekShfgzRB1r2ze7XWHuTLd75B9b47YZ5cl+vW
BuCEYx7mSaLSUOsguwAIpg==
`protect END_PROTECTED
