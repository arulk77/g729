`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
/tOehzaSQ1twCIl/WUByAIp//JK/pRYbLXVWyAcmUrZB9E64KWSbXFzQPRpN/NKR
j68d6kfhVaS/RxDU8MaouXXdeNTbdHMmOJJe4K38vI9CdrwLFgjZ1T2VpLF176KX
z8y9i2d2oJH0ejJ+3WDpXTr8PcHmvSkqLJyRPcfYIeP6rbVeQ4mu8ZSn3eECevVK
WrVFKhi+RsDR0VHPcO9qzzUttoL8D9yuu/ZALnpTC2/Rk+IGigJYPAAkDXYGaabc
KGPp8bZDqg+93Xps/9m10HI2iuU9ixzVHPtAdwgxCwxGmemUYVHCLl++3Oxe9QMs
3mKp54ke9DaXtH6SomEPXID2N6Bb5DcCBtt5fm8ftXcnvZvJ3OrIy6X3BT8c77Pr
caidp4BnAqWHhqpKYUc1h3bOGhN1e/T7Oz+Ou6UMDdIhENvXVZpkT1NzSDuFgXqX
/+FlJEWgvOOkn902QNQSSbMA0MM99IZir7BBOSnC+iV1TgMOaSZ0q1wfFzyfP8vP
vswPNqoWa0PxuhaSIRh1Lxqw/1EOdcNXqtDiNWv6Zs52hP0FopCdCU03AJQ0/Q7j
UiSYbjl/G8odOIDssZ1ITvk7scpaK9LSHl5THrMuW8dPvj+GQNB4VvIfRVGyHbTm
CU2itGQa4DfhiAf3DDMV9qvwBlIwHl3mPaipfMSwfSupIy4Fm/Gp0cGJ54mrSkBy
yNCZJ50dZ+tOYL2RVsrNtcNv1GjaffZQgYQgWSP2cjqOlpRold8JpfgwEIiHOiou
MNd6JawYETtnOqTIRS0h0W+PZ9AOxoGBTdT5qE96GfdxEXOkgsOnrkiyzS8oLODK
XMMUopC5IB62ZHSeYscF5F3m0J3LDS3QDpGF/hyrFs66XFs72XZgS21YHtffnY+O
G3Ul5ctsO6rzI1F1BiVBJg==
`protect END_PROTECTED
