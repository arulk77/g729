`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAXM+hWVVK7WJ90o3mfLXacLMLiawIjXnSO/anZmH8WX1
X6tY8S+6gNliJqDEqwKheuzpY/ZEWko079/4RyMOwdAwmE+7oFYJd+mauLwTksYG
OjecBqYMRaaGSAb/CIU7qepheuAYkaA0/yITUgM1UVR6mIp9M4gxKk9q9gSIEkRj
o1DgCYDBgIRTPjhpdqKmE5hYa9Q/+hjFjm6dmq6iU1bY9nRIZHP4L/hhqzqTbCG9
iI0pyYcgphrHW8inVBmrWji24v4arl8LqC0QmV3NM8aihcfVttnXV/3NUOIWHpcQ
ymvXXgDygDwViQ8rsuXig5imQbMN50OEKReTG4Sj7p//GPAM5J+0OPJiNTAkJCoH
TEWk88mND5MuwVNtuKkSR8uKH6P1OlFSotDpcACkbiEsfS30Fn5v3+U3Z/cRHbgH
iPJqfpRpTsiVGWzKz27JctAgr2z/7CKdr8YEKKGYCoS8rH3RQQT4joCjRcorek6R
4jsysZq2BuV0ZK99hgVt3FpEgfezYE4nULsx5RK6FUS+uGdnyTecGqQdu0tuswAb
GEiR4byWS1Gas50qIfTiDg==
`protect END_PROTECTED
