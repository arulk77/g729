`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49wvdSWu3CZYi6ENSPOTZClpeNfy2KtKGN/1b/uc5eiT
W20+vnSPICUqOH7EbXQEGbJ6iqCVnpR+dmTOoUJqQKsetkXJQWvNW9byCVYgexGz
/nWoT8L8h/wkflh88P0Xq3JHyFgmlru7uxZY041NtkL/nJ8Ols7pEyWs+2t5sF+w
V8brLV13K3x+EM59hqh488d5WWoTTAWBYCdve8jg0yF1E/V5N21ul67HFkZprwi8
Gpuoenha5r0NqhzEOBTEQVzjJotp3LVHcEguMMTjP4A=
`protect END_PROTECTED
