`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu459N8DDGDvspV7RcLue7PVQvj8hgU0We7R+BpZVriJ6v
yfuzoMnB9CjEJ5CSTsN57esaZm7hC4ZdIAY7FFCiUCg0FpQrYYvtq49tWT2+NTL4
ZF/1g2VQYLh0e9F9dpPZZl/fFlA/ZTkudYHN3G4ok56uD5F514EUn8gRW+ksjsxe
laM+aiRSmr6ycyTGlilYDNooFTQ3DC3kkGugf1glX13K36ZQWjWiDseuZ2yT6Pz0
YkK9n8MgGD36XfdgDmKVVnSGSQRjPSTM7/w0u+3Z7gZ+HoqF8J+QrHNZb94TUVDb
zUz7Ke/UVPd84JZuv8HjXA==
`protect END_PROTECTED
