`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aSVx6uLpP+aGadwosuBQzQAyy/0F5AQcQdbKDE8UXOMg
h+GEe7clsyHRE7K4qewHc06jQtOOeiFNa4RXFkJHi+A1zWWAsDGmqeqXMa5jMBwi
aP03j9D5B45m6y85PUTyOUvWsMCIi79KJd7/SY9mHNDcVoRbT3ysSKbzKV+3skpS
/Ed+dFMdE7FrLKkfLWiWG5Wl4offwgStdBdFIdIZgHgOsKR+3EoUHat9uYA5YXh5
174OxKqfD/uxt+42ej6JjxU7VNkf8htfCyMtihzC+civD4ebJ9/2+VZ/NhQOOJwh
V0da2NtpRsLM3gI6fWUdfaGeKs4Q0jAMXthaurzJuHLJ5yeks+LTrctDLfdtIgYB
9mFs3C4/iZ45jL+HIhNs1wSJcQjI1+fFZ+EBLVpzO7+IGHTjwR2UzJMrixvqfDY7
bJJ5efEMXun4ktoIML+zWBpdLqtK/T+edI6vwfEKQroeBRtlf0T/dKhFl8k4nWvH
zASQgitavt8bEwyAmm2K9DkpM/3yEH7P5fJzUZ/mBK4Vy0yojbZ28YF2FiJHeD2q
ZtTrthlVL2ybIFOxccQDwBwyk1NJndtwi5QA0/pJnTTzCLJled8YHmgAXiJG/EhE
5Z7qgDpLeVYJ7C6DRkMf1pW5mstt8qOcP2j9PvjhubVIgyE3hIaoPnpp0i+PM6K5
NiLm+OzCuG76YR3mOzjixHOqsaJlT1Q8zEKN65sP+Cmy9Tx1HCKEoABsVvXi/Nqv
wTekPu+lmtuqZABmA9h2CcF2QatPO7lQc2Mc1UBfurS2ZLtsMhh2ZSw3bBtRE4zK
Gz8WFgM0JpVylzBo7b/C1hbotG7WUzEnm57BoBDXlyqeTIojqtklts4Jp7//pufc
S2dLZW5FfQeh7CuWr7pldqKx/5LVdc0rEY4vEKH/46K7C8D1a2ZD4gybB7ZHmIB7
Fb5GQ+5Bw6uG9SJ5vt/GOvNNifBnxOI5k8QApk+cjsUDlX70i1QrZkrt78vVz8RW
FxM75zfJSSKkGgGAjR5L9rANfuhRswqrKoVxRHcfcw5XkJlwQ4wskcch+RHggiWC
5+0W1e8vPCu4hwSKCTi3RXxNQynB3mGZv34aIltuUe4PvXrCjw+xtOnBgvNTLe7I
zeYr+5Onv1mvAIpwFpP12TvcW1BsdU0Tam7SVZn0TudoloUw2fvdN3meYNyDZjKY
W5hLoNcFOZtZ5BnwoXGaZqqJR/SbueeBwc3zKZMp1t4UJ08tDd36e3TypO7qF8Bm
DNJsoMYoMCD6dYiouo3R6FCwjW/4aev4yu3A/yXjhpGiO05iYegDt1AWyRwES131
XkzNbx0a7z7j/n8B/Lr1tpoNAcdsoE8QRLM956RXd8VyJSuyLymwmtuG8F5rtuCx
ymp7Obrt3ITxGLYaDUQOPSryrG2IU1Dtwcc6fMxYmjzR6mecfD91v8hzQ+pXvY6I
cvXFqWqBWvM3+4hPnk2hrABJnRMbImcWCpxRcg13MBsbKqjecaF8WUKbJVLKIPoB
fD6WilwbBM3Ua5mmNCsyKeZavRY4KKDFqUbCrIgvwdfdvZy7xb5NzxR46e7eCp88
rlvsq8YMKCHAmccOfZZ7DH+JbKRvhDcqHmIgpEkbpmmKSaa4c8bskxqYJTq76Av8
LlIAxyr7BK8Bk8KdjvdezUJr4k5LWKd+uopWAksrL4QeeyH4ga+Ogj7kJdbQ6ulP
GAs/lsISbUaCa7OYrwdWxqfBWtrRK5XEuSwBOCEIrmjtxmIEeus3+tJPEqn6UaEW
onC51rs+tx4NBQTWR4P/cJY6GXrEeYnutKJP4ZQPLp783Ywoyexcmd63KMGi1ouG
KV9V9Oo+TPNmZcMrrXsOSIwX3db1YzLKCgEibtx2PYbOy0mc9DN/HWaVnerXeKxa
fE+05mUxXVUloW6/CB+p2m5YaWv+Oo1cdt7UBmN3yfqrwabiCDfp9CoaXhKWq2wk
xSZOEz+sar6FJA7EiA51U5KGx886Py3DaDLCM+HMLoMqhG2vZNOx0SvDYnEGe68K
Zeh+lJWzRPdDC/abNIkNZ6R2WHiZ1yoelAHeLvmvqLChWYp9jeQbzdnJTIaHsmWd
aVx4EBUzTrCCnXPIriATcBIiwytd7qe13gXgIYEGCh3xdjaOuzQIw9L5B3uSIYSW
zRX3drpZ59PmY9Dtq5JGbEsU1XCTfBOeFHhLHaYSxRPjmWkar/2QuXhZkfWbszLX
hNQlPF48rcIVcrIYkBYmFeJR0nyv1/G/SINYUpUYymuMKRcr+bdRs/rb0zEow1ay
GhdlS49SdpZ9SoEb7yOO6/lu9Nk1V6sfHRJfEyU3terY5lAVI2spmQsN0Hwcel5Y
uSfZ508NKSN30hTwDZRQvb2Teg1JmzOr12zt3GL6Dc2N8JWK+T4vMgLBc2tCmRWU
3FT8V9wl1SJwk0Y8xE70wzIQC0OktVI2TRX+ckwXcuXQDCSGfXNU8/MqwN557e34
eLEIRMTw+Yzd0+lKvu6lGBIa4zPn7BDeQXUNHvZIpeJ1LSvqFP/JWJ3tDeEYqzqp
hbhJFQTGF7uoJJV3/qRuYFZ9tUQ1Z8m+chQSxMgDnXIoqfvpAFpThxbP94QHt58H
hkdVw8Ucy6eGryAsfpczY+0DyjzrF6beOqLaHFV2FD3/p0oYkYgCrg+Y7NquITtG
Mn5sGSaWtGVDAtZCm6uE3qwppTF8PNdRBB8Du/t7l+hu5ByrwSoivE6uOnjoU8ZO
eJGIFlJ1aKBwM119rMHEP10yfX1rsraX8NYVqANsXMcdTBHK7vG7/lX4fpOtAgqC
42yq3PJ1tS3YasyZ7lsAXigUShvzB5S7Feu8yJY4HpTbRim+0eSI5MCscpGdmZPf
ZhRPZmv++dG7gb6dMLH7rlbxRFGj/chKu1RWgHI2kn6NMx2WXczw1AxwFe985rwV
YMqNrQ199+ar2hwigjzyaCG6I4bPVHdrGBztH4ZgQwp3AkRxDesKQVap02RxV5uK
MRaIQ362wot/fn69Lfm+v+ggQ0DoAJc41OS4kUjkhab5y4w+KgfH33J4vNh3YlKD
r/NhxcaZxuJJZQGyGjeknQfzTw7A5TQZKjNYpj3JXCY9qYkxWwzxfMQF8iyaaX6q
BrGp7hCGYDjDwT0LtzgpV7FA0tVXQCLq7uxawJ+QI9xjHj32iqByGWRDwd9fc6rX
Z//ko/L31abLQ+6nlpE80PJPRQ5RsRj67j/uAXjgC8hxuPTfw2weWa136hzvKbVM
AwjFJJAIM63JIUcJEnlYAzT/KJbxCTJ2Tbro6QHRu2GGwXQsFcNU5FW9PzdAoG0f
EDZOAj3PwFVwtyNUZ7yynXkuN+OUd+H3JsFSbBuegkRhh0Bit6ZAqhQsF1AHBr6x
QU9W0w8FJUpbispOJoiKBmdJuxtx36qyjxgJAxGP8BE1fT+fKYwhjLhYSGKhjoaT
SIgrQkf+uJYSB4cgrjnpKCL8ixm1xuI53GvvmNcjKOVZixx24AuCA5KppbL7Pbyi
nzFvmgyY3WrR3s/VszFaRgt9bqNKNjUVbbOvWr9NtGEEZJeIoBOUhJffiyf9sOv1
qhOkeqEz0aCki50jxYdwQdp0DGU3geyjTrpHmztFXTtNXy0J6KImw/96IXVDsDaF
MNHvvaRV/n5vbZiOLtkr7XK5SnTOxBL8FfLZtqJ8yFi9m9qiOYCvh4FetLskq2R1
et2No5XBnT/xp2x2+4Clw3iKx2dIjrI28SriHnB8T40Gj5yiMihlw1Zmz0Lr0O4Z
2UPaVgx5iG4MlBxwOcPgDx2Xfxh2Wy6rFJnYG6KkqCDEBxS3tmNVbfIKESiVb4r0
j5yt8pF5jHF8LPtDvfMRpQUCd23nRLQ91NvmpeB7NtJhAcF0vVjf1jG6NeQU9hrs
U3IbwzeOyNsF8eZS6CvYHTfvLYRGoEh4YacTxtoOvpVoXYjANiJSE/UCotEbidnd
iDPh+YlljPMlxCMEuZY4HUbcAl1lVNbvKHgQv79LI9W+R4+KJBOTs3bsJPSZH2kQ
RxPNUaXlUff/1Gd6pHUFOlOQanf/EQMcwTEPoJVPrCtWocYEBmkBz8b9w9ksNuKS
6hkg21IPBpMLjK24P92W9pCRh/i6YYZw7uotrbkMOc6e3GiNv8VMNV4LCRRJ63Sd
M6iosEVMAmrQpf9uayZzbHaGoYLeQBGUAEQH3E8r2egOjrjVLvt5cfu2/FAA/71i
4zYCsq9MxWvjRYT0yCmOL8iy4eYVGupLi9asMmph3yVIOd3Jx9o94b+I/XYwxYBN
SCKepRWasHkmFR70Zq8uhdTWX/5PbvxekfRqf+fWzzwtm/FguETkR4/GL01aC+iS
Y+bXANaF4VRTrVyFTFpMFDl+cISv1kA8ZYKAT1xsfHKWGX+BNfa+/jwwxZLm18gg
oN8lzt+7fxIgbmMJEKCdWJnTBuVwW437XndFFJmsN/0eIVQfVhiR2aTelk6owbrt
IVoT7EOif/+Hb9Y7V3LIQjgYHNmKlx8P3kjh72751h9S1+8vpsFHm7LuEI59/iGe
4V9hj8kmfxPWVJIZn0S7OMx4pdr8W8XsTUrPKLIbEQZN+daZBSk/u/OzdYamwiwT
d2XPi9ho6CbKikipmMwoE+iKhBaKqgpzeZUrhgDenhwWeVqAZ22cFGhBV/IUFFhL
1SKal9gwzcCVGjBNGHvB5VnkbXhxUHjWbtdq1l34Wp8eW54X9uvBCN4KDftWiuD1
FvKTfb4G3gm5KQj+6Jk+fLqzb9MgKAS8xa6DYfxQr3KwS6XmDEb8FGQsF8HGdbUP
VKniUdALbhRHlzJBWmspWM39e+wUGctxKeReYMy+RTEzHvhCLBj6iTkHNbhxJiwY
jtIDEDc7uexjR7a4zWK0+BBWRmMdeUQVG4/WUtF+qiDK9t8505jlW7Pvk61OGs18
FlH5/F/UhGJK1tZQnmzJ7S9UQH1KFG+nYUccAlRjk9GPUU0xOt8ILrIjAoOv3+I3
/N5+Txxzto5RnjUopAGa+gLOPed2oIua1zsCJaTFLDuUECE2aYS9SEpaVYUy9f3Z
k/9fLcMYzvYBSMKh+D/WP/sigU1ndKSzSXDvBbjWaA+5oWNMqFKG/g7ekiy2NeJT
PHC+GPxMoK93ozbOKjXaHHBA2NHJR+L8HAC3o4RmVSZZDxU0uL756gNaZNfcvT/J
0fXVi/pizV9sDDEyhYJea9y86CDM24wXb7uHHc8rCoOc3iVh0qn/dgBy4zbXJqf9
LHJl4qqnHa2bphMXY96Xs7FG+JVNkpqlGROeOBaOCppCKkNNFNESzA4A91xsvpD5
ylRnr5VrLpXJKgzUgtYQ2gtLxHvdD75DrYFp+8+ODVUIJaVRIZETj530gfEk6Zib
BiuAcInDkEmLPYoW2vZrm6MrV/KL4Ll2E8fzrGFJ1QmQ8ShZYgMB3qzwFEbM/RDM
EazP4qxZRIU6iWOTQNJ7ddjQQhGssINOBbe6ty9acigFprIClS6p6IFVlP3HJ5A4
b9ouYlvo5s84BhBYkUo+/9w03jPVYg8WVYFKxxiWp2YktAtG5Sq4Y2oeSHv51XlO
jkKQuw6JbQMq2r7VAfS1auoqdnO9fO3WqjlPB4m9/6O0P95fY6VvBcR3OoLkzYT0
/cXRee2m33AJw4NaSedyV0KjU1LBnc6/oJgBqWgTqX64xgJkhverz0/mf3UAUmlr
lGd33C+8CLDW0rf0f4olUtyvIi9/l4dQiypAd8BIGXBqfX6BCcrQmv/N7WpmM36s
YZ1g56KW+2x3sIOmB8OuHcz5NHkU9D6CB9qZU6mWrt9+0exSzK1djPnRLG+yigha
7ZWCs3aUQVqUpJcOPFwEz991EHh9yoPeSVej5fAyW//Tt3aesUcoVfIQxntkv8fd
9heRYPVgUeGdPuLxF2B2YQcGbSQO/TAI4u0wBbXSPAuS4j9joZVCN4PbsAnbqvUE
HAgNTKdd5QlTpQ5/vWjyu9UX9mD2hBUgGzCILU3kBd0wNqxBsT/ttNlwsPz4Q1Zn
RTfm7p+NQs0VhdkC9cQCOp6B5bkd+ic/Xsd6nTQIIIKGZWzTlI7oSGP9LyOAq5fz
wz3QV+/rQVc9X0/eYdHzrUvD3TA/s/h0WzDnlg3IejY4Qtd3//cYDFh8Ht8kSM30
YDFEj9z8ZfIcEdZN/WrfOlp3ZZG5JJAKAfmT1F4WXgtr8SUGc45XBOp9gZJ0Z+qx
A5ScXTil4gyrnaiANPV6HYDAk4ZFBHUScf/dPmG4rueGSS9ILtvKK9jIgaexrjhj
evnawiqouv1z79Y0+ChIAsol1h7S8BdXn1onz+SOT3kONVZYUt3rgvayO5W4obsd
su9kCjmcYB1pJptz1Oe3g6r+MHkQHs/KELWBNjfKyc7Y550kokq8BBAXp/54BkTq
gqceGpf1YdL4fbkhwcewhFbAbmMkSygDpe4LlZSJFIVNWr1lj2ly/85As2UMHktm
HyCaGpUxyfymNjAWSZDUC71o6F0y767xIqCXWtY4AeKugDHSBULztVNYbV7L+JXK
cXcRRVQX/G8gseMRjsoaDARkJaeJ9F4D+CEOqc4h1kM+BKNmnk2NDZ4W5pBZyeM7
Jj3IC9jDBv3TZew7EKXcdaCaqpqu0KODJWYBZRou53UUI/pUCUkOJNFr4TX7723x
6p/f9YV/bjFmRLrLYdu2KpTe4K2/1kvvJBx58ofPUmM1f5dts+JlwTIfHZitFXUo
1GJR7GvdTxl8Br5Gks3Se1fQ6O3/EwVsigeOX0lg+Ryh2kprHkPbkcMMAAA/bjeG
7SnsvBHusQdjo2PjVGWSWhIqP3TGc1L9KmWw+KLkjGP9QjXuorogBOM0M/Qtg28y
zivNz+iDP+6RlRwjN33pl7EOoIl+RzIFXvqE3vQb7i773dCIIjPFtlXwGnVSFDHW
V9QyY4VDaICvaWWOwScd2w4Zi8RtqFj3qLyo+sakFV2ep59cxvcI4vTsX757+ggZ
Whdm4TnnNwUuDjWWoWRKQx3egK4cmteg5a2reEI1IGySFLo1ZSQhYSQLwQ3L9Jnb
HN8P8yDh0bjaCEmK0rvGPHpbW7vMXh/gZQphEW8AhMA223+EDHSjKLzmRD3HE8/x
Cg880LtyprsdlA653tOqOlrG1BC2Hx3VpV1Kx6kYyeGQDL2/uor/O8Ff6e4u2d8U
UcsS6gQhbJbCARgBCIF7LLsH7awzheZogRRtU5/LUMANNbijkrZTGxp5lRcKbkMz
3zVVzhh+yXFU8cEleY6V0VEDOmCML6aurTJAqAxFXGfcaDDuoIehIGbhqjfEtYfS
o/B1TV5Imdyw9dKUk9DAay3Kr3SeWNkO+pi9tvKGqmgI67+6mOrMdMIJjO5DW+Lm
F7cttIkUs+gvGi3R8HK3PWq/Vm98Ll2CK3UFt8aVzecE2+zTKBqzwTrUrandOwoQ
06F+44eoUwFZnb9nsaWnYyDeiyYpk57FVitrLUmfhPpujA8Ar95q24/tTzg5BKvR
lCF9auow8xQS7i8QehR6C048h7pLM24TfjgczPPQtS1ywVa6fXgo0SNUhUS0sarp
7KZW9JtbqKpuyNUF0T1jDA6HJQZgQfXLmNphQW5Zuu1YWCWS1fHGG1Ra9KNLgM6y
atTZj6DQBFLHD3pUVkopqg5Sgb7oJhCrHb0M6vIV7YvYQCkteof4fYPWA2V5bu1P
7p0hI+9BAjOwzjEnHNKmZOSNE3nGfQ8aleCAnHQlWWyDKKiFymGhDB2sXf/M7UAv
Pa1UZfZSzTbSeI3O/oEditLcder6mARrf7KjUFL/J8t4Z5db7lGHE5vT336zgDcy
rXovPGDUFVYPBOI4zuyMfdOroJmBBkfURQCN5UH6RbAdeFF9lkF3q1zHbWhUNyeO
rHWdfm3Nr5NTqvjjkGIpTt3WUhoWtFfFFKPM+J5pmTiNI/YyPE6ZbntTHCujXSUu
WHu7MwTtlaaRM0ysTeFtkxrufPk+LF8vMm4HlfP0tleGx3JHr3cvTPDzyrrw+VIx
sHpBvJFCtVWgOUaaN8z1NHgBsny7XnGPS7Ya90ZRKIn9F96GNZtVRBXFfV8FuXuL
RXv7r5gWPzrHBkDlk30lcPjEjbZ/5q8pE48s6osF7GI=
`protect END_PROTECTED
