`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ab3t38y2wf5+qsH/48ktMKsQ9mALFmLsnFHqkMAYEsgOpeaoh2nziFEJyaBgWaE0
ewbxTcjAh3C9UDDnLqer3b7sxBq1R2OcQc+GEY2FmGLXkbRo9wWRt5cdalXeLwSz
CCOm5BR/C4GtwmwcOyqN3Fc/AzwOrIkW9tgFXayhMEwI7zHzme3Y250cVf0F1hbv
MjhjYzqOr/D78lDfTO+e0cQLqRb1T9deZCyRLnX9Xt1KbrV//QPO0EXgoye0NBfj
nou5OBiA7ksCi5PF4wwyG+l9acj6Z3hjOk4innBbBsbqRWhzl9Ruq5XYVItm+0zI
TKLVzmZD0w+5lHD0lGyyyOZ2dJzTCg/tXf58+uWJB71baiv+D3qJi5V0iDXKvzKF
M6sPaTeLwXqRRohnTtrbM8OAyWZiWgBrSgbKj2x0hJg=
`protect END_PROTECTED
