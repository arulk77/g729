`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP6iPB24qA9KAIHLlKezrwhUkixzWAka0BkZQANnEiRA
u++yv8Ro0h/1m1G/OQ0f9ScoN9+dK6VN8ZnUBv0JPhQ+Gap4cLCji/OggMZ/GtLb
wuZi84OQbjgcWa/6n52L7+FGU0DBgcxRXhkY6UFuQQbPctnUzWcljT9Uj0DH+WWh
7jTd5I6uLh8qFpwzXKHGcH3SSDPIB+qi/BnJETxZcV3iisc5da5GvYP1AMJMBfeb
O9e0m8YXu3o7xsRE7cp4rv4Uzuf+iYrGRXSShbGWahfHIx2ymboowK7dqixHnB/P
q2MwCFG0XjwnriATxXSVrH5mGRvFibMmX6kFfpulrC3arUFQy2EYHKGg3N4j6WuE
8zSDxJqQcczWZ4D9YhW7YIo69m1vvOXbWRTrkhzqxh5Bm9rDauNN4Ht9xiN/Q5/3
nf4Fqnjm9xCwlPk3dy6PFbvsJmrcGqcEBJxJ2WxA/ESZWDJgRW0Fz5lmPW3MHqFN
6YLM1KGE+5baW/ZetQRCB3j4rsb/MOIoWe20QTbYOYQ+WWXx0EB86TPub+1rWU3e
E9q9rVxx0vKwOXwcG7MXWlPGaK1oa114yQQRS9PstnkR+YWz/wvPaJbTZ6d829Dp
9b3IVfr+3J4N2tHbzMFz3yqkBuh4bEpMLhP359YXXO5W/Xk6C64GwWWu6c5dEtx/
CO0Inb5qhr6y1lqUYlmBXQKZW15Dye9HMo2nXjC1aZkFBRprekIB3myCiyKNBx4+
qV0UsKnzofVkq+UleglYQ95pYC0Wq7qiPIRxO/oesVntRfzCBmytpr53OuJsoU79
OsWRGN/WfQNR9C/cDM1wmJcNS9xajzUJFLnPuFTKRNYj+ETwalu0EpVzHEg3dT/P
o48qnC6LAT7VXrGzVpUxXIwIUBhIdW5tlJKyTUks6K4XOfAbzguNtFrJKyIuN4PJ
nXUGfwRb0srAqsTedMiDHgx0YbV28z7J2ycPGdi8i/yTaV5FWW8Sr7jNtywv6aUa
kE3EbS8UDgcm/5bhFfF+DIqu8H3Qm6j0vtBgj4j4NeTiBoEFT3X8t3FxEylRfJVu
GEZQRuZbT3dtWKHmtIVGbG7UOiAXNNzRMaZvYOOUhDzxvBjSmFC3bRgDTlS5cqAS
7qOflwozVMBxjccNxLKRdGrL1d6ECn+nl43zaNKJy0UNvqjik6afo0l2+/nZHRFf
oqZqhMEKpdwB7NKx7J0zkDO8Pg7ZHEpACMaUn8BkU6dViWWzD+6ngAkuz4eR90RB
LtTHv1rq2pr0tKrs7ob5xPfXHhIOC++AC8dBc+GO4u1uJ5yfIzL53kdA2j9115uZ
WB0v360MH3/9vT6BeUV2LfXzWQVatNjufXHKxTQ+0gY4ubcfiDWOG8OLhKHwpc3Q
cZbFuwlZ2QctW17TF+PG+TGA+HGrA9eATBdSFbtHwncWSPrb5xYm5fNutXDI0UHy
sfeE7ZIC/wyAilSI/y67TpmKl+BMRAzF3H1vD7HZFh/oIMwR0/vtDDPidUeFItet
lU3XU6sQxNGxbPM4gkQLBpSHfb4RHuCr/KQEHGX8+gfL3SemzMMlDhsX/Zx6i12A
naB5R/U0BARNJvYxatrcG5iRnSGsHIipQ7jitS1Ef6SACSmJRrFovCmQmeg/og+8
w4UCGgBTPXwhyJk3PbJ7j1tXJNCCdI+KaGG31OParVfkH/VG5RAXI4gjp0PptQIt
CZokoBgNyL8nRTzdJ0wz1GRHjx0GSSXVyav2U60V9KyheHvP1F73F6/GHcDN3Xhi
sSAO8U/TwqVYuVZ6GsBclVsSa0lhffAX4RmmwB561WS+zf0C7KYmm1y3qlliJa/q
6A7mFqIIybpeykCDHzFYEAmvGNdgUjxDUPoz+DEWW7miUNeCee/6CmkbnpRWIeoN
L61YtuS3ZxPs9zY75y7lFE/zrwa+x+WY+82fm22KYzklMF0DD16HfUVlJMoBOb5H
KfD4LMRZacBjbshJJzWXBy+LRp1EfqwwXuOJJBOXJ+RpeRvDlSTuDonHfpQobyuJ
6eMTEV5625tCj+V4tRlEzSAfR2rYDQxqieg46PzOyPFyvB0OUf8UeYHDMLMxYLai
pqitJ/RbZ6dalU7EUW7ziR0QoZfN6xtI+HGN+k8v405iFKI1Jl3jIBbtELE9f5/n
3o4SSgy8tX/ysSaxhMfEuksJoRzYIEFAzLZq71FGsbhtTd6rhqrn2B8s8ahhzwLj
mkekWZCitChNBismzR/Le1CbiVdb9NezcXliNKd7yflx1N9al6tB5YuuMAy0hR1Q
p3Vf4kWwSxL9supro/52/G4k5x6DCcMJDD6g9SG2Ko6WEuXRAGP4Z4FjI55cxfXs
SUZXqDJY032muNM/8EtPF7B13FPln3ptaoorpkDZiNrin95iKn7/vUaZzlzs2u8c
BibkLiSlvxIC9KFxgXk0IFulqNzkS3Jg3oczTB1qCl5Nh4i/gBO9NikZQLqnU8QJ
3GwMcJsMG15q8bd/ewAHhUXery/jyUys9GTIegVXtP6BFHUYsTt9YFA6drx6gA6/
JxYu5+bVWzYljFQ2U3OKYH9tzIwKoVunQM6cqxCZ1g1oGELVl2NSjK9BFimPs1wn
LSYX651J+cniFqALaWW8wjtYVwFupIaoM5LfijHfNNegGCYVbYbqs7cEfEz2FMGh
l2MQEeQyHMK3XDWwtqkayA29Z+31Xj46VaFEjKWFMC9XGl29X0/OXh5/W15UfrOs
w/4jz6lRuh0aEQI/os6FbEmiOpd1RXKpkOyOCr+DDifaszvDrprvyRsXKSp8BWhm
J2MGVY2DI97dffi3OfgyEeco8jfo6f6pFyPNc6IkcLZXjIcalaTf2XE8AVT1D3JY
w9jtgVMD1ZqrV5k/cIFgiawKg7gfxjH7P/oP0SOkz2w1LRMuD19aA88QGJcxzv7b
kcdZnq0kwSGySelDTvPjOqHQyS4OgKjndIr/gs2ouaLbQfYf+sic2uN89dSDwEIC
BQ7DptX3AbZApdd74STG8cafm0rzkg0r6qvwDenA7roVye16B1SJmmGC+m7FeQAO
s5vABBEotQ3xt7yL8wAiIAj+vGLneMqjscis4XlL3camnmm5zJXPQ2hnU1q1BPG3
K/H9Thpw/W/CewM9fYXK+Ao9YaEfeOQAp4h+PevWbUHAHSFW5dvXn8xO4S800EaI
m8T2tVq4TuUnJPw5SeNMdKegFj9q8CWHl4BZDoyZIWQDOBrUld58n+TYtRnZ4gFn
1DjUJRdYNXf25L0iBnAK8+vuJ7CX4zaOCegRuEr0cIaCjouoBaS2Rrs9bL0Y2HmA
QUcBKRLeEKuL963skDJj9tgZvJdSUhCS/NaeTVYRrIPW5k0fgK/nwTDeep3zQjU3
UoLBLa0x7fIQY0vPU2JoYpNlvEtf1X+KuTQiOxmMcGipGnJXC7E+/QtAmKHp6NZd
tzm4I/vma6UDxDFiCGUosvDozihbnl7nbU+CAU9nt8KZLMlbgo8Pdm0mADpaytBc
8qg8I+EHwzT/ZB/VcJ1coxIlfoc9G9i8pDEXGdeuqPNpqvjTa2qslVTgHZFsWnSa
Qdfh4g1EKwZa5eunqBrARz2nVwRyc+SirLZkzmcO0UK18hciEY8K2UaGDzLN+avh
ks6mKaiDA8BvCoFM5TY8Qkb0sH6U7JRJthFuXPrC7n34ghplZab4Mk716r2tMHo4
CtKckchx55ecAqtjcmzO6HByQOfT6m7FlKw4rjO1FDQbBOhRYhf0kQfaHKnLD07I
h5XTunWB/18vUhfmHu4ulLoDjSILaxdfaaCmcM8qvxRIbyxE47aBvj1p/NjmKiMg
nJN1cR1qk+KHIPCDa+inYpO3U4beM/pfMADVdWCRMYI5AWH4g3yDDCE7knx7Ol8R
3rJ9J1ESNEEXWFvpS21/LgvW+prYjkizudPuFRgQn+odv10jOht0XQwgsIjNqIIc
jKYyeKZiwqWTiOL0DDovKq4i6M+TY45Mjr1Nf44yehclScqoaEt0qHqGvEH7xwve
8MAAuDDNeXDMdCKzDSXicTGwBSIBtxU4xHl6HcyLwLVk8gIFBanitMVWkqONnImh
bmqhYXOW/7EUraMCT2gTlh20vN7u9msc0VvChloI9J3wJc6zi9ut9dFScfi1iNVV
HlHvRNY+lA9AEY4OHXE43WRPtPGWOXNI44T8PEw/QnID/a4fcaneyQtdJMWzNZpJ
qVJsIXJ3+yvQgJ3A5884CQtFOgxjnoHHuZFN4ALxGEJxrXTedEfp5g0LFhaHM5Li
bT0QRGxNFzQqJUGSv0qxUyZkMpveupromgrXi3L92yxmgZ9D0uBVKlTS1zWzeqLB
QunFYeO+yIG/jG1GxOx+7A0LIy6PeBLkW0c+BT/IVR7cHeL1FysoocweQNu6iSjq
j8fyouRQpzd11rVqg8rE4ITPTkET0imuF+p2wTJ19krOBBepnrLcJJKE4QZjTfO7
EjTK+QWBgy9cUA/QBbZmrYeW1wnh2UTa/OaAl9jzTeRI+UvQuoC9btB1MgcqoSH9
sCWDboYQ1X0/2g2Tv9TwxxQFNlpnKzY1w5pjzAXCRt027CkFiyTzKGJkbqjK2la/
8QFwVz0AgwgDkIhT+8o51QLIDznFGh6psl5FETCjqP4U2Sp8qDBn/y+HQv921Z4N
b6YxBsw2qwqWij6/WESc0tcbFtvloWuJUenJrUyRzCfW8S/WA9nW5tKw8JNM6y7W
L5L+qpW6EZd9R96elN90JAArIjXjORLOUcIS637iv39Foa3P/0sad9Z65WxVRAza
Ii8WNz51KYfRuOSoV6oIqQ4v1xap4RnuhImC7ZlzvjGkM7LsXmDFtStzPAOXiaAq
zQrh7DfmrteKfIG9XG80b9VLiHkPIli/h8k3L+o7UA43Cj4018MZJlZvU9DhTM5G
LbOAS06kZqrpaaY4EvOKFpr9yV6gL9S/RzO3WSp2NFN8Z+39jr+3mOXjBx+5L0aP
1+epjpSBCKBV23Jal/SXHF9VcxiC1Z2iON3lto8a0DT+8VBofKsJmKqJAp1T9BK0
FEzBCj0H2hElWv/FP/65FD9brl+Bku2ohHBeGJYMzclStRxHaAS/oHq3JHLbxvVj
w1p5mCiDkyADEqXVFMNLXp9OWakxNXtgrJMyvm18ygAV8wiDJK8kRVsfZdNIJ8sA
Z5EBkg4b1jdap+T+rYXevXNH7gL3/+JC7iTiRu7/S8C5pn+rMaDghFz1SMLRbvl2
pX292QQ2OLA68tj0s6mQwSHx5CtZBygaX+NAibQBee82tt8P+duXajKlbp5Kw64Q
3YNeCrHratEXsP4upBJx85NoX1f0vSlZ+LYbUN47V2LB/50bIvE8My524uK+iiTv
8XmnBn+BWTQYKtEI/Frkbhf/N8pjsNRJNPW4F4QdszX3b/18FGLi3godBLU2JuJh
iQHUKP9hrouuFocHoW/kw9ZRViUKzKNn1jJBDjBwuAS+MuVBmyY7bcdY8e3hq021
FzRJd/VDQWPxIhkQod5v4CNSFngT+BOqMtEKjmGTQ45TtDjP5BEb3exGM6/iqvbJ
TLpT0DG69s4puH3mAf/Y2FcjTQM3BXvZUnmVbhMdqkuCzhZG9nmaBQM7WqqwJVqN
uASGm3iM+4iEH2nm3OQST42qOOhQ/WpNl2Sur9PE723aVn+VLMihOY5xj2Ntat27
gBSPRJTSfAoA7V45Ey5FiQ8/QzEmsD9ava0+PZjH+o8M4nsQQyN52CEwBzNMGJrw
qw2ZQqAd6Ir0+O3j1whuEM65idED4zYjLdCjSIeLOet6UftKpXodRBN6vG115NkO
+NAMTsrrduDpVY1JpSN5U/24H4XjH4Z4RAdTKQOdkR5uH/MO1MNoA8j/tvAO42VD
ryyYIx0gLXqpk9TGsMtPzOH1XMzqY8seJfP62BaB2kwKz1uA1G+azP5NBabZkBky
2fOHUMl21nUIMhbsWcATQfRNv8iUyL7rgQhS35ImiXmwmzx6DXlBD4toECbwuKvf
QAOL3eWdOkKB/783zHliEE647khCaeHWaNxIRs+RDfleNy9YdZ5/LjmIKPE4Z3zt
YjjMxhWUL/qtdcli/90FTiZPaGk9YNW25GvsUx4O46TtctpQl8ucoz9pCTMdIRzJ
UAdcjgD67DZTuAC7ed02udubSLU2FWwmdRQlh/b3TOkcAEndNHk6/bXLq2GghHtV
pq0uMLRrAvRD3a7+1I5BpVwtSTPEGgrA2bX4domyyb+jQnK5wdFlZZw09IhLXxDF
9rjFCQtNnrThF2dPWaHUka/DJe3D1UM7eXWoK1F130HaukxsPPkXjxiiZBTBoLKY
td2Ajfg4UICA+brJnZFyZb7J0+2yKGhkMYYMN1aNT4Jdb6jKSiq4dU2XoPUlhUGg
LTPoLwfse6QD5Fl8/eBS54rPZ5JHtM/doylngA/jt1Ma64bwkDPad3kil0XfNXyQ
sc/StS9CkykU2KPhxyQ3po14es7DRNWVgGAPZuT2KG1kYypw2ReiXmbyyivmaBWS
+8Nj2IHCh8XOTdqVjwjU9b69jB3IFS0Yzddokb+Vcs1ca5qoyYtNNGBdjXgjSTtR
9HawoDlSIVEwxAJClQ6h7fOBSqK70XpngyoaQsqlE/ssFUzKP3u3lxlWgVpYKMRi
M0+Daqt70JV8k8n3Gj+mkahBu+S5yOaF+RIJH82sSsxmZ3SbD7UCAg51jqJILq55
OAIjGKWkfF6RTFr0C35x7wzEN7xn410vM8qWcTTdLrgW4pRdYPlPaNTeL0dzDagY
bGlV2sjfIyBlAMOI3I9aKLTqHLBul2gmm/choouphgiPI+1Bo7Knwj/0V83VFtep
59fnkuxGp+1OXPR/IEuk89kTzsXsSoL6nwdh1F6TMNIflixVZMW3JiHksJZeZbzO
+/Tq7GpYWXB9iTyK4qZc6UsinK7eKonnp3zqqZELyhuuk4pD13vEh6bmPo3KjQ+C
YE8v9le4/OFjEpqLdj8Vrd8bll1Rkem1wE2cGagNBIIMFKQDZsiCQkwCvJTq3yyR
SuD8i3ZYY9nzcKDpqMRh9dq7758d8b49d71Lno9rQTGxm4m+BiR5Y5t1Fu+jVrAa
Ovrrhi3qres0teLrDG6nB9laz3SSPKrLq4M7cy9lu6xUlceF/9BHtI9k8k20fhTD
0uFmvObjnhR1r5u1TdEjUS3retP8qI9Fk5wne3zM7muIj5+ERvYizJN3RNqBjrki
3Z5MEPHyz7NyTft4zwYVM8Yz/d13wtW8q7CR0Zg+O8mmz3hFLK/eOxhuf4u5+pnB
Y1i5ms0R6R8MSRkMKXjaG4d7nZdLpEdzV6J7n1QliVYHoGg9RfOwjgCrjZM1tO85
B/SdNzP5XLnQuGRw7KmiVDc+9MLerajOfeLJ7Hbex7Etmq1L6OaUBgm+wFOwBdn5
A5pNprUGV5QsvT//3HxNU6VDL917h2l2UJAtFtijDzyypMphI/Y6wdI/SNHlinnt
nTt5bj2z+NZ0oVpkz2J/29YyVR9mON9p310a2jNr92LfOo3+78JUAvER++ja3XVv
S/ry3ya56Pj+H9IYR3xOBuyug/CfDS0WyefhYb0x5VGAz/SrEHt6p3cZl2Hj5phm
r95leCWVfIwxspO+rSPDt1/WZ4tQk0JerLHTtFNBIDzDOvJs25gO2GAJHazouoMp
oswlRpmppUtdW3nW61Xg+TEBd0TBDccaBBkrq5HNwS+OlGLffrwfoUvsVvcHOpeG
V3T20UvYX+N1Sq0cY09KCxqOG+Jd+YBMGxqo392jfx34H0ZxTuQBP20uUjs2R5/u
zskCkNBwktpHkTyHY7meY3cfMIGV/qrf3MJ/Xs0tAZj5/tanhpA/6TVarKwbHnbe
GItMIMIPZCSPL0hu2Oz2kli7QAbs2FHoLkD9qiwb0oG8ZEe1T42YXS/0ql5EwEH2
bJBeFgn0m7nZ63uQH/fVucrXTW1ZRhFI8lJdYIzevAK+y2IyALtZX2GxH/rGy+06
G8XKs0M/Y1YWD/BnhH2n02LIhJOTOa98rZ6CVxHZ7RaEFTkTITVPAdOoHraMu3DF
OmTPBilV//hmeTSNHX5Q6u9hus0F9qewhe8kQM5vz9Mu1hIAlw2GSI8WSkODd1D7
R4wR1huLPwYzgIqxX/i0ykNvjyK25ZY5sDVacZARtrx99nbBv06sQE7Qts+BHUMq
CczqM/F8rAQ8xtttSRzZCnfsqpz6ZCfrR3l6kE5buLvSZ8K3RS7RcP1d8NRqnwZS
EZqVL4Hyx56I1wRwyWDoMm30Z+bDz5T8rGG4n/+8scTA2rPaR6YqU0m9Zd4HF/ln
HnM+dyzua2lvXC8yjvUVXz/qeIfRbYpBVXea2vFmHJsf8lrYEFJQazxeugB2PuyO
SdfkgHlPyGmXiVrTjHf0zmoHkDNyDxc0673hhJBntIshjh7hE6XIjAyp5ZAIgC4u
joaH0RRdMXlHKRZsDxkZCrjjKkX6bIesgqmvL8bfYidjfvCWPFn1LznyjNh4g+hI
N+qKqW2DnCEBTGfRRbpa1SBja8YxP2DnbSC5hQn2+AW3Is2sceLK0trFMsZ1Pz7O
HfpitOBbGU6fKYZFiiPSqL4NOoSOgR+skBt5Z2AHk4KG+q1oGIsVD0l8CSaIyH/O
ZvYo1CMqCRrg5ppRH26pKmdKtWOF8jLsVycLVAZ/JkiwPTSmtc4ea4Fe9BYUwXyJ
TfnLL5oqS+Ce+THj451akvhvri4MhQ56tMueYSwlr7nE8KnZKAKl3DryKRItx7Ql
Qj9hKMq4vbPacrDjd3FpclEOhwuyHvb6Dgs2G0SowiFCgcBdeKha7g7b5PiLFhs7
xHZXBv1WMtMi8U+m2LN2fx490wqn3t4KrOINJyDTDrcK1/r8KtVZU00LoQ9aRZGQ
DkhCGExIxoJNcsM4YS2cuee4pDDiuZnjSskIDWlH3bKp3QvDDCUUpwA5sMfn0qG3
U+MZWZMsndMl6X7tKoJo9wGeFvsW0Id9l5kLhlpwTbm88d99g6iMvI7sGib6eIhU
cOT5F6u+leOHvvi2IwFFxqWXfwlyZymjP2r9Ic6AZXqfYPblmfGM3Ye5vXWQjEyZ
rualv5K/X6az2giIG23pzmPrGaBWvKYCrznNy0LVQhJqmi0uORhGGEfii9eJwI7I
z/51fXVVdzQL3bcFlYyrxOFb0kyhVaju6J5DgzRosRhbWin5d1p4C3Ai7N91YhMQ
jqnmgeqcQEKhwtM6xO8RBnb+wyDbEUrRimys8q7GDlxyvpb4q2pAhYGVoe713swQ
zcl56OmZbW6mn1DBQ8TNIY64zhI5SRJ4lDdV8MSjxhd1/b4EReQkVnthP0t1zsQj
ZeHJ//ZwTnFpq0zkSIbuoY/aSqGwayLGMEUjURVYcLwOWJe3R6rt9WV4N8hlugv+
D76pD6D7hXLdclwNwjvp5M8xmwH22ZPIfuQkRs9EIHoTvC7osVfARnybmI7P5J8z
HvPRAQ/Fty8ve2vZw3PvhD8gnPeMDTPFEtdlx8G1UIAQRA7qP2lWkCVyWMLYJK7n
Mg5HAGJZHnj4N/CrNreZFDPVBmI48LdTQ6WnXlWkBFT2bk8odhlhdQR58xld6es/
kwixz2U6vVhpdMCHhU4DXJGZmy2RZgqLlRLf1XT02gJ1RP1/UjxJ8IiR+hJHOK0F
DlYMtJy3Uh3Js16YeuFhEBayTXIckzIkXHkKijnLiht1LztsdMqreMFP1PxjLXnI
acKRPfd5rmyOlkmPISyBtmB6t5iLCChvnPzk00XbwvKPib9GShVEpowmoDGrD4ve
MClQxln9JUpLMZWxdqEsn8BYDsIuSVDEhzdEXfKvJOa0/QIeoflI3GmhA0hZLx9n
PT6jP/ElUBODxIjqI2ef3aUcrjCcLIATCbP1s3eBML9dISbDYQEdoUmMVvRn2QrZ
HP/WP4mfCo1wFPDPmaeGZRSY2l9nftWlJfXCprNjL2oKEWddLo/VN11vj1ANDzmF
O0e/8jPItSnnm9YIk1vx0ANRBtlbDE/qSVNYlkdvfqcZEMpYXjuGby8eJlo6BIqO
bqJ8hb334CDGoVPQbZNtsLCKvEHP0JZ4Ql1j0J1HhvPQh3TOeyse9fEzBiX5Y8HR
wyYUW9twklYWGhhN9PEHsT5X0riqCPZuhENZYPgoI0xBMX383DR2xDVgKKKc3tTD
97xB1vOgiyElgn93eZII05XDf/eN3181JNs1anoMmv335XoR3EvbY+SrB4qOkfRK
la0jDnMF9137OHlLiOecehOR6eliGXNLagjhK+YOC+b43EYzN50GvtsbggDRlWJo
WKW9e/dagZlO9v+HjXBHCzEW5Bnfi+RJl9q8Igpf7Hg4G+Ucpq4qymeMgsxAsGmX
u8FiLzlJl87UpV/jCPd8O1O9NoP2+/0F24htpc3j4/rVPzjfkhtOJOpOLSETba2a
oOeaSfaLTI00uVPFGBXKEMmCZJcJQ4MHPXu3O7ABOX0uetBk8/YkCEBwn3UOvC76
1Rb1P1rM35vacKK0uhLQn1VWrp5OXJzNeYGnFxWuptoi7dc9LNutA43NEbBhY4FY
nP0qdNN58PoK2ZafPeNCCSwC3eCHVeMmygx1xwgwbBoU0H+SoyVLE6ZkCivQEBI6
OiLaiNpoapn6qoB0zKDBwFeZHKnhIE2G5rMmC/w8q1cZPpeiGZhGTaPu/r0B/8lN
KBCWMbnX6gbKotpjRMee3EtEBhn+mALTrVKrjpkxuAmRwbsgXEPfi+a6HbydKGqW
y/jq+AbZuguect6FGzs7DUmuLNK44vWWm4e45L8DaTa0fndty3rGVlpKQbW67/9S
McbDRqzg1a2VgQHPsp2cXxp6IhkLi7hRWL8dzh3YvfuQ9vHcuAACrXDLWjIQgTow
4Y12Bv3od9atQgRmveKjjo8KlHzvgo1g7jVmVYgw5M5rYla3XPwpkAmK6Z15CXGv
q8KaxjQHCKN+qnbD/rRBu5VZsqE3uVE9SK0hrOpVQKlX5Gr8A+I5s0dgZfKYFNnR
lmuDq70JBvE3ftz8A9xpEA==
`protect END_PROTECTED
