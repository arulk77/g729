`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePyypztiGGU5xzcjGEk8IUoOCa61NDfI6X8KkLXwgOgR
xJ3JEfKlXUewRnxoLpxZ61iktoaMwFxWhsc5qylh1tsf/W7cvEkHed98BZx1Ff+X
AFzAUG9XLtoM9B0ZVfEh3TfFmcDK8A1iWSFrCjuHzPP7OJ2LzWE1WHCLunHIKYA1
bGekx3HgzO2NOdsE/OLxtXxtkVT0uHTfXVUOerM/0loSlpsLOdJq1FHWpMaK865E
lQOL/oAlWkPNnhjJvh7LfRlcG4olPmEAqPq+fCAbpEM0TkIJ8O7cX1bh3oyMcvsS
EQ+44M1zjqAJopgIm93p7N9ZU9GVUsW5IlURRT0aaMZVihgEv2mtKIezfXNW3NLc
o6RYHMR4wClV5i/UEtH7QNgZaWm4ewwh2i9MITW7YIjn9LEfOj4PMTnOm7e+nAJB
UVNjxt4u6QhKRudjmOoDBnoBGT7SQYToYruCwyes5BVHkpzIJtG/NqfiOPzIxW4k
MQoiW0E57Yxbuh0UMDq9CUTIfUbvEOpXPfiKh2mjXobyNctC9dAqlkXnFPAguJ59
JQJ0LCj2flLil8GMJh7gU2TrqzGDFSgOCNw+uh8KqWoCUVO1FIkNGSwmX6WfN+fB
XYxJySAzloQhi2BGXlsWN4oRjmUHI0j8UEY/zDw8Z8E6eByDtFlKVyxkY8l4YbJn
q7GABS9c2JOWPiBNLlqSFhiLePnYV8+ZKFxpxnEC1Usd5cSDh0eH4Ba/FdgIdn4A
c5qJsnnJa39FYeIhsVUIE3tdM7FhxcglRIaNdEvGPJuknHvVrrYMb3HMaQfDNDAL
eCv/zz8r1BQxFmiB5zFvqPbDpMcCW4oVDJZavijZZV06wPUSXs8YbgJvNOegEOBS
b/kmibVYhzsR2iz7n21VS8UQ7pHjHsq9mva2OqJNi+GG0ho29EkUqq7VTrTCxZe9
0vEFsJr8znwsQ3u1y6FHGi/ivwyfZ7NbuqQEq0a/msbhbnDea2OTxrXcSAikgFgM
QJ4el65xjpsfmkj02NavGNF1vrNQb/1fZrUp0B6Pwd0Tu1nrhqN8brYDcSziSCNv
TRyH51xqYutTpsfQnlk4w3eJ5kjY6ElAposZErADPIIb0BOah0hMLzFyoQTRWlxb
+I9+13jSHzvstxy/XUraUxYo/iT2S0JJldGUNBZbYQw=
`protect END_PROTECTED
