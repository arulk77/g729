`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFgE959UOG1tecjzi+sjhgOxNqWS+EXj8Oxjq+2iHLHD
xt3ADMLYh3iVF3S3zr2WWJuDHlVYDNbW2Hi27NaSzsyTV3tteB6EhjBFxo8iNdKl
84uATfuM1wZ1ptvbfKeSuH7HeRQNDFsHEKYBUpnMnLZDDaN9UHZTlwR3gWmuXctZ
9i8A5Vo51SrPQcmchI3kFg==
`protect END_PROTECTED
