`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFCgVo/sRqymlHo+L76vABBSuQ1TF8aOHqz0eufBmv3F
XN/omXa68HVHsy97VMbVsPU6x3lUTKjEZy/pUiPXTcfA31djIOqQleSitx/rSnFE
TT0DnydlsF1+CPMJ85aGEQlPx0uGu0Dj+MM3fGS7PHnQefdwdAqYEHFbQ3UnY7rJ
WuLhyIrefpC53rpBF/ULzg0g5mzc5TQ8R4ldQ0yjtTU9llngCZxo3kG8ClttjnFY
oYEdBKSDP5gOwCg+IfctjTaxw5udP8UxNifjN+OxUC7n+/nta1KYylC2AGnMIP8d
kV2YA/mD8OV9mqTuHGpf1n+VmyCX4DcLceuRfY+v1FrDL7jcJf6YmXathXgEtMQj
w4pg2j3zTifk1qNFmuG1CAzuaQZJp88NaXQcDlFyzt6qXgXtFPEyzYpZYpntke+w
q92qIqoAPAMpBFs7mjk7a0zJd9bLVGT/0GM5tTzszsVeV/feDiKwsM/KZIJcc0d9
mWH8phxndUX2PFdGhO9nICWkjPAhNHhIJ1Y+yB636KodsSL6qbuIaU2sSCRvQBg8
7A+8FE4FDhYhjzakHwM3/M9C6VWNckHc8lAee5myMXuteO3hSmHQwVIUk1ZmZCHK
vuFTj2HP8ghgGaGiqzh4lCV916NiT315IMv8lyMQ6l+WteQdpC7cG2yfO/X5BIzc
B+g1sAdERGmoCTJSg5AnDivp9nl56FK6bLUaLGhctlHEeA7wc9wuiW7R0uyz5NCi
TzuFZWSPvLdz1Fqg1NQD7dpc+YkzUvIu9qEGQLmTeNGRfUOmbELxSehObywxsVds
LMK5va0i0Vk9m5tblaa35icOND5UYO1GtZcZ3MHurpY=
`protect END_PROTECTED
