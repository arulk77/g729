`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47r2+LSjSbc3VMJ/+wGfBMOE7StIznhlI5PWdu/0bcm/
od0IWBU+2gwJ1yVLJKTFJYpe5203avWU+OyuU230SXgOg+rsIadkGoHTBmi0LS+v
/dCTsUQNqUTCZiWSAaKx0hB9rLOiSt3f9mZwfCdm6+bTYEVqwZVUxeVjutbEPIdY
ZAZJaExXEk4uV4Ul9zkA11JNmR4Bxrcv0hs5LUo/fG3bRaExwLTGzaEVN8N/Ciqx
mWDhpnLGhncc58YXBSuJ0WpoG1IvqmY2dGly5et68H+2yUPyc5LGAYve/5mJIs0S
SxL0YgV/0sMR64nh3FLkAUyd1n/bqEzeAIFrcaaD45c9yNCnEhXEPkCtuA08Zy8f
ab4gHBQrOZiKeTmPtg7vgQ==
`protect END_PROTECTED
