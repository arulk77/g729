`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveALx9TxWAHzdxUqUpDXFdnoACc9b1xNYC3EcjEnMdfka
oM4bw3mwL02pxYqooPg5GWgyeD2sd3PmTjKS/00RvvcPSO62syFhyNyMGXqt8qSl
9xFZWRw+wW3EcOC7xub4Cu7WmINjWUSaikr0Hp/lfPgblvEy13Evp1t+1KN+iB1y
UYALG/0A8fU+JBSvb9U1vFtOxipfE+mZICjyWvYbiYhMgV7zuIBfCynJuBUP3dAr
YFGLqPrnktcNdbxecVWRxt+vNRc0+ReIfxADMmsqcZwePxZcxKkzZv9ORYkRhu6k
1ywqiPO6sOiL005JukD/wfZao7sSqBUtXsTymC29yJnEeP3OSVkbENkEFHwk7x3q
j+XKBZQpZLMAsqEqCF61goEr6iNfFgqrOib6Zz3VnHwZRqbIe9uU5kOu8hdJdiDJ
MvKvrND9f/sKVrX63SZcGB2yRQM9Mviq+0mloGL4EODMkJwJofvKCIcVyd+/eBKf
gDeSn7ButUQtbjdufazNReRcsL+3n35eHCXcT3XK2lBLr/RQs0ScJwknm8DjXdI9
OlWK/qnUPHAVOt+Bskr3NIGtOMB6APyJvbwyAJZIqLS4A4E5WoVaLJHKYMlXBoQC
`protect END_PROTECTED
