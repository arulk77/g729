`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAeXaf6g/W6946lEE5F8VgQNBJXzslpMIBtOgLzQU0cwG
M8phpjIzayxDjASL0Vip1QRTOD4EeqarZuAoQKArzdjW52486C0W9Jtc7Qx83h3C
KnZ2xqV/ydJHa/LmMXUzuTl+gh/gBJ/PQOuQuBEyKYPT3IreB7h2u9ItIRu0Hn7V
7pSULqC46qGsUjUqg9zeaJRi9/Zt94/3ZSGfe8EIxc9JaH5alArVntZONpYIXl9d
FnLuHcZLXLlxXNcJkIz06wuTJWHK7DjzTZkHGTdXIkqnNRSomMyOSiCIuS2MNzIM
gYrYH+er+bBZG5JyJlkviO8fwsQ4ALyZrCL9KF8hKDwojCb/9FBdZR8yNB+GT25G
4ryD1K1vx5BYZGL9WSlI1gQkU5V594Vj6+ifmT1zR2eqecurNOuXZ5AH2CDbr/B3
M6TVqmkRg0VzwD4Tg3wkTosN9KwPFZZum882xcRpSEp5qav5WSdkdMLpR2M/qCN4
5WYJLpLNulG0Om8qhUcq5flBXF9FdAQmJY4DbmiS61mrOMKqoh3IzXpoDzw0lXmg
fU81mhRsTJqMv67mGFOwjhKKO4gFoj6cHQk3EYoJKwRdXhO3/rF1u6aG0q5i5T3c
NBupdwHXDFD7S0PodGi5VdF+R4uPOAy4oP1sdBk24FTWaCGmHpYEu061DDJqCNDP
KwbDfYF6jl00wX4Sf32fVPgwN2bdprCBxlAdE2xGlUPPH8flBuvNuuKXJRRQeP57
d44LndFvFDHah6PLcaDzbwiyZ1gMQdepkY2UU8f36KmO14tI6gXQfpGQTUIL7K/T
ph4pLVXL7Gi5Qj1RwP8Lmz11ymY+3TSTXTF3fzdUeudd9SaNbYuy0QGrNP3TNcyF
c4Pd7gAJ8LuGH4K04iRMpRxragWXHKSdQEcYjGHMlBLp4G3/sWCu+UL15zAY+fOI
yPOWJrGlJXmWWXpSgsBxS2eEv3YwMtfyhyuArjyZJL9tIisGYFOJcOcwBfp9USP6
DmYas6ipDfbO4DI7mEXE9lWuOIWT5A32yJvTyaIx8XSnseYSGA3YDRObZ4ljJie+
CzSmYRA93KbJ/oc6Gbv4ifGZwkb9oFvamKthQTMp2aYjdhDRPDFVeXJsfkBx6Yjf
9BwWOAGGAlmQUWYfLfBKcZspSnudxjJj06/eirWlFT+a3tEk0/PSMU+RXI5VmOtM
sdob8WopAY4FTWXoPEiTYAuJY0EScquahtHQfb3t/oOxIPqLxmFreozEKVMjPde3
JultDEUPuLug4KtOnDRktUMzrqTKQLzrx/dFf+lsAcjMPfAtQFQ9eQyZllVCl9rA
BqyY0xfJ3dlAL9m9UFWXNr1AD9DEhEh/LJn30nOfBNtMddYI63V5KeAFw3h3Y+j8
1hLUQVIS+7AjDcINytMy6iZGbSHR+PFOO2vw4XVX3qy5ijjbzVIqwTYXZdSgJqah
i80zf2TNS/Zr0559zFW82G4d1DclY+dN6e0rIFZBh8By/Zs+XQTPSpQQ31HRmKNR
MXwpCKD7sPIZqwLNTG7E27ZNngyOChkw7XQ+LOHOyUGqb04tWKi0sH34uqps8hRf
EvxBXZZ6nMOzEYMr9FtUM2zJcxSd8PQzciNDB+GF6B3n6Y61CiYqoU4nrA6Xtpmy
jz0p+tTKeqtitaKTnbj+/DNZUkwp6AZyLKR6z8mCVboCCcfULH2hcD82Vq71cZ8Y
RANY5jMl3CmluzfsrkIvX/SiwAOalIv5IAdYNdMnpfIgDFpTjIipkXeJELhK6q+Y
OCNfFHZoK5iyc1W/mVL+ClJIGyyhVd/jkVgQXQs+iiWF+S90tzw5s8KKNWTrecg6
a+u5MMEHLVSp50tTf5u2aKoRzEHx03T3dBiy5NNvA0ExxZb4gbSjfPqhL7zH3nci
Ku7rJuNe+FL9H/K5+K+zqup9gRoZmV6D7Zcxnc7gsq7BVLoAiLfRVxrQgZnvPoPU
mlslNqHmDHv9J97P1UsykiHSrB5ZOEHNyKPy4wUaB2zBZTan8Xm9A82SeRb5jY4/
ese8rV1t27Io9UDJ5FEC3sefo1J3nJGWVV9acveJgQZGMtft7RKtxQWouqLAHzO0
5EV91O9ttX6SPTktnd0VH0PByhEUOA+ke19z+cl0IwH971Jm7soM5GXvmsoseMBu
2iKH7C2YBekaB+1URgT6WhOyPNTtfiSLocbR8p1JiR3W1dojIdkEPz9eK7rZJ8RJ
y0WoRgAV3aEnXBRjchdOvwSP69DV5sLwgk6ouEMx/Dn1OGwViUfkbdO1ck24oKD2
mrE6viQ8faFzsu1Udk0ilms87rVoqQmMr16CzjHeyOI7CMt/BSm5clQ1tYDCrV8X
CDkv6pbycWgS5KFIs4fY8SR+7BYYLxoYAmEwPatkIwMus+lioUSjF5yqdu+3tCYu
i/Ay1XHL2ul2ZZEMWEfEuPNlJssTHxPMZH2pOqz14XYM1yvtMYMpNeTcVt3H6WhQ
eckXdmLpjjh39XObM1RLnb9PaDGRLJIo102AChp4c+Rk5YW9BiDFfjTKZOJQroa1
QVs9BQS73iIbLd6pZv47cHjOGqOc7wjyuRXNdW8sM9ptgLKXJLAeaalHZkKEoZaQ
8+pJRX9KD18mq3shlkQQrWXk8im9g8zfjCRQqDntcSiaMCaD4hrDPeVDLtO9DnyE
9Um11PlxQXdx+giKHLVnSf7WG1nKTYgzOA8eTRR5vbYw7fF+69slURfrEtXnF3H4
cyLel+j3mMs4av0IX5eBJpECySSl0jCE/J0o6RhEWheIkFXb0Tol3enABfh7bz3N
i/SH7ZBv4u8mNq5MeK8zWpzHvt4qNnD2HGHT5Cy0FEVQsh7xJpIGNudeAuU8sjG4
5sA2lCuIfZh6oIlrqJCh/q4k04jco6ia38xncQuPSOIoNr0PHDYhF1y1zihSWPY7
Yu2VNmc+6L1Q9O7jF3ew54rgPcoTQobTU9O4uTkV5IwPOwJWI4TYsVyA3uwar0ii
867HW9ZgtECATIe1dWe6jERt7g0UWAjFDHFLUCnGpXLl+Y4y7HMcSS+CwDAZv27c
Ck6kJjcjo/+MNrwJGp9WnzoMIDqtksZcddFFn9u+hVWH2GuAW2eJjxHG1BAD3iyE
+hoDZi7Ir+psMJDz9W+EI0jUPs1yK1iYYnZO03R9z5J1H5pDZEPSiMenaoZtj7HV
uKlxV9QakF2g7Qw/jasCdety9qqavuxNWLzuffKpUcnkooTkJw/gQKvo08rtc/fP
ICt1yrya3aNc+pD6636uf0Il5xgTbp58dnLDwiaLh0moy91rBBx6T31y8jZSMo6S
dIlAAOewnTAdQQP+MT3SX5ozrIBc3UYVmPZyBwgrQCwan4JmS1MJb693ZfjF2Dbq
9mK5QJRBAVTo+6Lo7/ByXvslj2qJyZ/CjPQhYybFVGJbiVq91mIJRcE8lsBADJdX
BOaA4IL8uHz81FS1r6g8JAZj7MjA7V9ZP4gGDdSO5gWjdHv3ddN5YTTm9rCznbkT
QLQ1vPlshovehQcOpuEdDBHTZCCj71zjkyenrma8ery6g/DWd91610NfBsFksWKN
JljhYI4B8YCaWSzQsXT2xnsF6D521P0aNxVXAGBCsXvUDm6Y2gJiBKE1UQFFoJfv
B6A2CVFBRMiyINnLC40IukBhv6RkksnJfIriXSPuqTlHXTsE1jp2y4yH094JhFkM
vuAy01xqojdTV+prvwAOVc+gFDSBbjBwYqw/l1YCi58TY6syjxo9R7QlhWD5xqW2
C0TdmvdfZeyi0a/9DdNDtFSRQgBgMaHkqE0gdJm/F59SSJK+yJ1FXWKd07OhaQ4Q
HM7gcWfxXNc2BVAFkiEGtomvZmjYie45RCGFMA2WctX5bFG3qLghTFRUH2AjY1dm
5RPV2bqC8kViD2RlDX9pux8IOv76FQH0hKGqJ4C9X+NaUL81vj3mxMTStAkQY90x
PtFGMVrVr3eOmx8pQ3V5j7Jk/uGMtrLrmEJQT/fwP/80soy6azsCwWhijxAEak0V
Cg9SdGKJkWVnVOBgb/nRAad/GXAbUBxodCEcHxAJNwHmYJaY6xDzc3EDi2m+s9vh
VVpVEKhZCuv2xdzN/NN/PqO+RGhT4sgAV9A8lHOzgfp1lMIaPm2qGL00vx4qRgs/
WoGxVDEYS+1ok4hpM0s4Dlb+Z032opJS2b4SH4VfR7cORzol+g1WrbwI62HpMNgS
3HjIx381zn4I+MdWajxM5NX+8mEYdgKgYR3Z6atxv2+JwCi2xOm+APAE1k9fuFps
MMmgh0XiZaaf4Y0X1RTOfr7P9+T+AIOWZVRzb0vlqhSwngM5BleWRpz56M7XASo2
R687PDDlBrQwVXF7YXx3D00SQF1gtpvEp79Bj6lH9hyIXpI4hezzoaOpjpHpB406
nzVMfa9031aifQJQbmKjEPx1mCPRZ0GYz+bIccGV0aMqe/MZ/HD7imAzyJ+Vpl/5
4NEsfaGaV08PzEQq+gS3+7NpVNRYQpiar7LLAIpQtLGReoRfjZN3WSY5W0VwI98E
9sE5wrjelUSYWR7dQEpKF6Hw7S1AV7kcCx9+20pws6kic6z4omjBdEBx7RA5naHv
oWI0a8HQmduu2ykNvMQEMtpfDO8NWoIdqSVyVA1pkO8wJ473cmMDaOT+QtXKEBoI
hbMig57DAzmIXNXlTjZhJRTvrNkb/1LucQf+Axstfx4=
`protect END_PROTECTED
