`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42PMtHRha98HsgTDPWTQN01tQpOKApgGGcoD6jHScN7L
CaYEMwnGYLgZ6yX9TfZMKq8iafGXphhsB51DuyyZ86hDuqrVlqNLSu6P3ATXbYio
6SZyoqjgJ8t7dSJzyCr+jGSGIvDqizS7COctWzPRey856mN/vmD4gaJ5KILuVsRS
MWVy2K2zg+Pg3egMLDpS+sRVtSt5G0RVbUJuoK0JE8R6oZZ9+KDQeZDFBav48MNE
s5jDVAYYhAu3kJtcd+eJfweYgL+zD3RZVY8jlYgAYEr7ZHRc7PnyYDSTakzYpTYK
ehokYNchKeAZXT4KGVTGWQ==
`protect END_PROTECTED
