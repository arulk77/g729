`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2IT501eZw0da45JlosBrm9BD4EWgHNJmLQ6cUP9SP+Rartn3pjFfCt+8EEA1uywn
7sstxFkIX01NmRApXE4mKDUccSzA+7vdFTLfwVR81/7jkOtaGkgNmaX4bg7zs5Mb
`protect END_PROTECTED
