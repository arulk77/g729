`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOgti+VD/fKNfwZzgsgKt3NoQmV0+ZqI2cBVboiolBzC
Duft9uJkYmrwzUVnhGtdfLBq41awdnbTQpoNpQuTHwkjNRXkCVUMvJu9U7yS+hew
N5oF0ZB6PNpz/PWK0Qz9QzAvH/Q9WHJreNl8rXC40AUvcar3Dww6GL9Qj56pJArX
Fm27HzUCZtrfNJzex9IMq77/jut9VD7mmgf+Hq3XxOEoWYES5p9FmDbi/tGZRZGg
BIQ70bWO9ZAbLs0qVLu849f4n0hi53ML+XZ7z+/eZ/5zW5hfxV8wz5kU4zDIpN32
HE7SMAV350HrwaeDKJ5wAw==
`protect END_PROTECTED
