`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48UNq4KoBL9g67L7fQlwiyT8eYb90b8fJCjmiJvu0pfE
C04T/2cALjP08z6L0qMK2cLRUlcI5bHs0VFOc4c4F1P6SQI9Lewa5pNMSbf+JrAy
sA9DIuebQ6rXXSArwB17czric1Jk/s37vkziIGuXbf0+7S1yqB09E4TngkblPf7V
g0dEeMA6Msdbn8RTkTG+k0XTRG3JutQTBK4l4W6oyMMNIuifBol9NAlN6SDcJxHc
UNYlggYw7bAkv9aZevIM2bIVKoXbSqbxh+Lf65IzGWukwpWmDUK4Ga95gfoNnNe8
muIE+Ms9zDRCGTH4JMGY7A==
`protect END_PROTECTED
