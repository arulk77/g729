`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
SqpYWMA3YqC57KZJfQIKQwB4w/5q+8EXDA8aXg51+dFKpVLzUj5240WT4A5MN1JP
GIs7dd6jXhoBp64jKRSZgyuBTYjkpxInF/7NN1yhJwFVSr0Cnh0I0JTfjXeLByW7
Cnh0H12xYN9E5mcZ4ZXmL1Si3X0RzM7lYLCwdyMmqlSOFhEh4zi3ZEddfvibwSYT
RwIo3dL8taIakMevrVaIlu/b0cujcx/5uyN0Ln5J3paiQTe60AN150B2Vvg/S6zt
JsggGZUUkUSQackL05vrosaAIfWtxFHiSi/40snIt4CVknluZr7Z20QwVywaa6U1
8e/9/ynLzEZLYbdXns/Q+3gdZrbDFtu2m3BayVcf4Xw=
`protect END_PROTECTED
