`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QNw40IqJrFvY2E8HYWz+j6+4wVYggVXEmKrz0iruARWQkUQAwbAJ9zc/fsdwlAt3
ki1vD9cEzJCUi4z+WJNtyI9FXFk3N+bimwRCBItMrTHT95rfrOFV7q3n1P6Xtpc0
px8J6tP57GZVLLrbQEC2tYHgorUKJpZ/8bpB3ACvnzkLAbNAK+iISRh9HT6zugB5
`protect END_PROTECTED
