`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEWiZPOfpWuHwrvDNdjlK0Gwtd5J2Pbj4x6badtf4hdA
GCAMFrVSpnJ/g3Pm6BxpeTD5WgzyG3+rzFZdABTuYuUkXvAN7FWTL69ajyd5MtUy
DRkpujliHpJO6tp12MZAxrmKTj+aMXbnn3YP9In88GZGTtme731164FoNmtRFVLe
BJ9dztwqP82dDz5VijqDNCf2VYYuvCzULCcMon/MT5UaAyahWpW9G5nElJ/tWJwA
Q9RCl9UEtmBlXbbUTdz3SFzlt2TNHNabdiFAW52QsEPIJj6dcK5deqsv6fnpX4ek
hHEOmPNdi6Uiid88UGXm87J9VE/DGGPiBZDYv2Fo+yMpMUsYmvsyVmihqaEx8Vwu
UPnKl6cgc2ku45lYwDR50acH9RqUymBandepO6d9z6fff+Myk9HLDOFnA/Kj16jq
1pStCsSj+/cMnDwN/G7D/VKImXsC/rYptYn9+BHOZwksC3AlHXjaxo+hALFX3Asr
qh4oJfWEKK+JLzOXe7d6djbahMDvZJJI86ZZw4DQwj2oNRNE59Qag+p2MEL/teut
YqIDtCObi0C4EpkawP3phfVBEWwzsiqNeopIu+MwrKI5oMaYS5EeqVDlUvVIOYYp
eXQAtJt5ULobz50/lkUCj+Kv29efu+rl7g4of+RcpBTTyav3KZFw9WFGTCjFcrOX
`protect END_PROTECTED
