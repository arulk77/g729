`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu476EVXfN9buM4i+pbd+PCNu6TEDY1/lIpZdbbES9gC5s
QYhE4SvR5wsUl3WHbzso7KraDjue5IHj5KCkBLchhoTc7xo8kCWbtWo95edDr5eW
zOojvFswMbsMEnpu36NIpxfvrBYpee0/gz99Q0gGnoVyxKMhBLm5ESV3xaa/51vS
Gk8kgAfxoqsbC4+wD8L8kg+AMReuQlyd/SHOiwOmgZ1990zbDA2d25XtTNJ+a0eI
F/YJ7KFQAVJaF0wD2nWU+NDvRdvEpmBB6lVxP0Eq+rg=
`protect END_PROTECTED
