`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL89c9yPvHLUIpmyvKc/FsQ/Bt3Ey8BXSoL3ZoqjyXGAHj
YUiRG3urSTMVrFyGUXTnXRjpzPkLI/717hCoCW4L7CiLmuMpwlEnGN+XJxYRTiP+
di6927KuVyrIBlCXXitWvIVhFG6Fn95ECIspMrgVLcv6/DTBZIQmBTpF2JSCsox5
ynEyVrUls1gQ0y+SBZynM2m8/JW6XcYembJtZ1DSXlSqz0OgUf47/D7bAh+hN7h7
+8F4vIwqecBLHbOEWzkOz9X/tD+3vVgu2NS+K7rhfICDNxJ+XnL1t9oY2XkR77IS
ynWEbpZcm7iwsqcdkH18W/Mo56/EESjqlXreiiFeulMjIQmg7diNP8adu8kcArqF
wBXZxJfkwM0ZfZx1liI1G5xz2woXdcBxUaeEXPE4orvg2/mzM8QFtS4SMslEWj2x
qF/fjz5q7COQMidC2M7GhHX8VNzabKKK6mWtA4QNtsyFx2/LqWhL/9t8pEIQnOu7
IdpUCcPXarDkTX+jX8KhjNEyB68p6hbCk8A4DFQ3yp8lIz8ckCQue+fKxvLAtpzo
n8TWWCIuL93oLMf5e2TTPygh02F18id730TFFDHSbRSdaCCd7Xn+lCVc33qS+BuT
`protect END_PROTECTED
