`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8STC5w8m1ZfNthXSgksfv7xNDAivAsp//7ddY5DpmgMw0
XoMc7lwPkQALLIyILZ4AUDfk3gCfpmwblYRvGEAZsBioWKW/EvqgAE8ZW1Odpwdr
mPkFMrDvHXuqlQQswkNA8B9Z3I9MgeoyxT53BF0lYrBmkgG5RE3FkQDicT9d9deJ
n9eftUrf+H2c6I/lG0W0yVbM3MR0Mx4YvqHnojyP9N7fJGjQCZRNS4cCPwgEqkTB
5Wy16KlDc1+bc+Fb2EZGXK8Crxo7Kb9bMraz+sfSu1TGEZSqaGFORF8qSc43jK5j
257MF2RJ8bWKO/TwE7/BVEzsdGqaOonTyvfHUSKkaiDby2oHHe5jryirzt8vncHO
F12MNVtsEoOly0WgtgsdqevLoTLW0Cw0CIcGKySh1oGkUaxqB5PiSO523cvxmUr7
CFBz9/98C5yt/RVta7KJ7M25T2UePhmAgUOKue1DIyqJWRPTPHVHzINvTL3oDlHq
Ue+kA9hK+QGeuax6w1YxSzPpXIK8xeOt8DD44slIQp2w/qtDBRU9kxUaBiZ59CJG
/rmVc8m2woK//9G65Xf5s/n+H2KLkMPecqCSnTN+axCJ+zMonhHkpk4PRmI2hnEf
8ckC47vNbb9YkhlzMWIpZQbLLwDuosLuY3v+/X/4MqZ4+s993WzEyWZhPXyc/u3a
qhoFyXnI7z4DodcKe0HyHU9G/U0zJkvcEi7ncmEbiDMuTHLIMpVIqnqsYbvTf7OA
PQzRL5axmYYC9DN5OJmtz+Bkyow2MXRw8QD8p+TuxlpcTbmBWHwhDEluTxiDkEly
33qpS7DCjPng1ZCNDvdGKRy9qGT8sDy1bLFRjiSkZ1ST86HiyBkphzwiQxhETzFP
Mr5JCSqkMgfzJFtgF9Q0XUyfYY9Rg++JN3EJFvqpUTRH93An4bqAUGETPYA63/5A
mlHXqPs0WCNM0Y9Z30sozfHOy5FTViRKP8tI4w3Rx49Ypz6F39SzlKHrIIlmdnEH
OjDMuppsxHGuGSs4W8VpkEnpAK9L8nnxI/wPsfOYvU492DWyJcTyd8pND+rFQGdM
JfvfPO3fK8MR4BYxI5usi8XHuTXqpuaRay9ryWmKZo7XCIDkIJ00Ic493VUUg0b5
gJ1qyx8X2cE7batiHY6uz05s1UinbUA/ieY2aVCEAS8WPl2UVlWJPjSY3tmF+Pkk
0L0n7QdEqGvy77AiVCNGVTGg7oKj4P/xw62dl6JgkMNuK+eG+xAldkSZ9jBKz3pS
`protect END_PROTECTED
