`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
me8ffYIZHdk30CHIQ/TOCDig6wmprxqxGS4Cnhz+28mpVPYrt01gkYt7STgr3Ok1
a28LCtMauOA4NZQxjJThEGHQjaannwdW3anZXhCWvcIWMGdzTo3n3YkLrE+GiT2U
aomntbeljaNZvSrie22ni4J1wfmgojg6QVH1PEwcVAnHEKWJh41VWB23n5yvJH13
RAlS7FdNTZRfnsMngX28Elw/MKal0XOJBmvIvmZxcepVHK4/octUPH3zm3WQrE50
`protect END_PROTECTED
