`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFOkoxo/l/4RWJwXmFJp5Ni7YEsWbv8WYdC/V60/wbcr
bXZbP4NRUwr+hI6zf/tCfgPbrA0FebkIYee/hkvDaVriznpV/ImxQU25IdGCo5LZ
03urJ0MVr9OpmOPH3m5FTnjM5JT44Ro458VZOVEhmzGL2wEenkf7z45ZkSAxy1dL
3pxM6aJF1J2MJ7pwlXAYze2QIS8jVl7FWR2URCFyYsF1sR3fJRiQBb+Fu+Jei3N2
Ez/GpLRFa2XzFMWgnLcgsOqVnvtgplDx9ny9wfgXDdSuM1qcoIz7feqfDgmr/bMF
f+yspd+AH9rXHSDUhFS/HMZ2WPNDIPr8hvz1L+rt0gQ2uSRHL7zd5aIDn6RONvQS
wD66i8TqBBOkdxU0OsUIGDIOXszxOD3HRR46gx1Id6ioRPa95TNih5aXZDqvkV8n
I0rRuPoV+JWXDzoo1FOaTDo5H40f8pE/IoLN9sZfEcEcPg0TDthN6A4q9rvIljaB
XqWx0TT/J6lPFYOymVNwiQnmb73aVvSdV6qNqiOjvx9kyKJtXJxBlOO0YkScOM4F
`protect END_PROTECTED
