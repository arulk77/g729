`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
CXDo269tkFVLssJhCUcbkf5MyUrKdR9Wql1FdXMdNbKpHX1FELpP22YgRie3rxzU
er92fkvXlUWn5ccGaUkK6DmpwAfd85HrzlvsPaOuQEE1IB5S6vXSNO2JvhMQgJIK
r82S6Cw3uUpqh5QZGjSNIIMveJ4c9a9NtaHKrnGz/qq+QZxPIPePeiI5rcPfwZur
4mfwqd0+M0PD0/Nzwv5Mfrjrpj40T2LbNM+wirxmIOSgpkBlWrmP9VCDD/BO4zaf
WX+Uxpw0m2aBZ7yjEXtNrw8DRrKzrBXMyjWOsHtzswN4OCPTM9UbFo5uiK3UQ65S
gEqmanCrb5yDj7P/tXxL26UPYx3Ubbm1XDgX/+g9/PQ=
`protect END_PROTECTED
