`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43EbTXpQgC9q0qRaLePtYoIwQJUtQDCqK+iqEQwQTGs+
TDWw16XDNZmex3iu+4On1xUsg7Y3zvv/RYSGMpy4aU89J+eJmLG+iteF//hESfRj
jQvTB0FJKrqWfBUI+Ao9x2mX/KwhrCfUe8yzf4W91D0=
`protect END_PROTECTED
