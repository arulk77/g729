`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCX8Yv/6mZjQarMOByMF92vXBww1N7f87fpLAYI1UvWG
O/94KkCmdUG/Y5htrI/iW9Hgx/QaZuhYchzouMIwx25ub5SaRp+AHNGZWKa7yGD3
U33WlTnoAg7RpQaYLjVUsoLxyx/MFX64E2XEMCO0Ai3kj9VDeLxC58gRBZ5Aj9UZ
0/Y0PK5xz/8XpgAGmiC+oZdzZJ/7khoH8Fj8Yt00CUb40yYQqVzaOsdLz5NWeT9X
l/pU97Me4cF6lh0sKi27glKxZQbXdUdXFt33QuYhGxK1IXgV/vtGVRCZc2/BI+WF
TBapp74C/vgXH2jh9dCNjPot08wjViSXz9dKu1dABUqCaBR96JivzPCPEkq5r4TQ
ThTnIlStVYxuNKG2+QkL9mZtLfwQ0nlFvgsA6UHwvo9CzAhjql1xjkDi7K9m0pG0
PdMLePqGWXfbMK9H677yOIW2+XA1vdKkEJHnzVi3KVD7A79p1ZKA16NvgwTPawU3
PqufDDhoBcdnirodxzCiiiiej/aWDUxYhN7sm89Kc466oT0tHDO+9dR6qeKx9O0U
PSNSA85Txbc59iRCSJQiz38mu3PfZq+NdJMIuuJkoKIDnlu47n7qE7X9DqhH2SS8
4YCLQs5F7KR/Dt0BkJWjEJMC7v92WiKjBdaEaq4lsrEh4/jrxAkn0mDsA78Bp3Ec
YtnkkswMvID7ycM0guYmuojZmAPjxTD6iID78rJdMUlAW7kSNtz5jxUUsYelb/e8
FFhskKajcymj9IglUGWIMp3gI6zmGMZXHKbt1kGm/LRQVE/Cj5CzI6WGFivUT1um
p70DAmazH2+c0nEXK/0BqyGx0yuHTOIGDTIIi4K9OcF/Y2kWyy68fit43dpci1Xl
EKXddDwuuGqN35d2XVsAa7Khs/U/oY1hOcUioqETZ3U9hBD3oKnO44HGQAvF9fDl
JYeT5Ox2sgKY52ToDZd69rzhYYi9tuo+mPirZYf8pbEOtPQDxsWyPeZ+gASGGWMy
X0VWD3sKJb9ToK0SVCX4N7c6+3Hmk4+REEUGtwdv7CjoYTSoYit/iRniT/XkXOUy
ySgXdGQPV+3CvrtHOg3GDqLhJRXT6Kkg3cnZHcVGPdItfqqBQp/6I0EkD0Mv5d3s
HCjxiSSz5kN3RzHtvCb+dUC4vHlS9XJMVfDsLM3OwnsMK3SMvvpbI99NG5jJ12RK
A6L/nMF7mXZOiomwDahN0SY55n52sBTBw9Mp2NeHmTZ/UvDol+pcLql0y3UJgzmI
0znS/hpFzMUsXa3rLDhcbbA5mZjRc5pMJWvvb357MzyVXlSbqXVGJeLmbKX8lorc
w1BjUvJr+4FQbuCGM8Oa2Zumn//ng9y4H74fhxFa16gRYZBGynq7dyNdtX1bcErp
EQXUnXvFJbFX4DXNC4G5A8vghuGEp7d1lWNX6U08mhcV1uOgKMzowifg7evR7XeL
9Lo5CKRIzzeCG3GVpok8jFxeYM4M0Bkl4s6dta9BDKgv9rtQNqxltMm1yJCHPMue
JW4bxNCWLDjD3sr5xeXi5NqT+LFCAOZWxWK0Vp6qVEfru5aECEwFsgcqdR5S3Eik
8mkiwG8huhyLU5vtBKlc5mHkzt2gH/oTKOgJyFblWWAiksmjSqcBSAHJMpOIbFGO
nDoPGFVQinu5n4MvRTH5JDuxr9TXfH//d1osAuDNRGACIIycH+1pddaTVl35TpcP
BUo0ibSe3m3u71ogxNjR8Qn7RhD26tHFhzzqKaFOmX5iXvZhUbmuAaEBjOcltPwo
wlophFOrFrQ7n18DNAeeANI/BinqrVDjfnGqxYFDDrB88sjNLGYWomeom3NlnSBI
KTCmdX4hBuvkCWP9jLNHTd9vm/JCWahNHNxY5CkFkuKzpQRHiYq3vesGKfRdKX51
dGrE19O5HGza/7g2mXzArm/rBUDu28yZwXX6X1hRBqh6g+4XW85PcESoR2rqlfgt
N8N1futIMsbRUteX8DnZqAhP8mZ7hgakNk0HUiE9gvt27f1yTedCFnG6JoIUYGKI
Ezl52dfkJsB5K8xeu489iIw8f6xwB2vg/3bjlK7d/VJZ4zQd7sSqMIteKMEQ7Wzf
VfYUsx068eSka0gmv1DmMVwSEFn+5IGVOIwf09is0suWuysgW/rsUljSb5fbaZd+
kR+Fyqr7Oh3gOHZuXML3OooiHHWeVP7u5pOc72Ni/N66oIRp9tCY7tRFrPOGPRu8
oMwb4mGwnCBTo/ZoDDPDl5nZvB2lPG6Jh//48eMlv+GHNRUTP8VuX+q5n1q+p64U
nxvDeKZWJZdnl3nhRB+ek2dGFEdSBPADe0haYrCxndLXF437Mhjvxo7CcC/cn9MG
YFkAazT/smbpEsu5EK/pBvRuybb9mvrxUklrA7kc/aWJBO2J8t4sgbu4tduQlqDO
hcBjU6fSJRNCPoUt+J7fSYTT+ccMN4wPqHi8zdTcZEy5zQsOlDfmJtCkbPoffDh4
9tAR6bl4gG0JUwdG2BstzSuZDBXzk5bvbO4CM2hcQj9ddla8N0epSL87+yWG5o9V
5aApVw2UitPSsg5PlJhmb9BW5wR+u0ypb3CGBZFty8wL/q4i6hxwBwpNQykFvkQq
vb2OHgKig96ZiWq7tmqumA7qItCpGUM+BAJhnXVPt7Ct8bUoPmcd1/YR9jLWdCzc
orBvhy7+3B1rEeqaf4QdAgh12LKq7n0iR9N2FkpDmzwU889nFEf1cp9LVl7jox2f
rqyOL+ynCVJ3hHscncA3C1IoHcYOQBPErxafEZ+i0BgcNjaJQLehpIjZY5ry7+Ka
1yRn2rfrfHIIDEThZl7R7PtuQXO5XX0ywZoLgI/fG4C2q3YN7RaY8C+gcSrySRm1
nAgPzNRxK07L+g2RwcNalQykB4+N4mPLfwktiOJXHoxVt7z2Mq5ebxJqnWP9QEgH
m2rv41Y+Xiv4QnyjA5+ZcuI7uRT7fzscliJVpLgb4On6ehhOQ+y7YgG+0xc4tY60
wONtu8A8P43rO47LkPq86vTbAWio02Hv8MT0iZIcQWd++TOKTORd5t6mEH7S81n/
Cp7wd5FYnZPpGMg1SFZ7teI8BkSB/9jcwuGjeOVYHTggJyuQjWR4rpl9zleH0A00
DKMIE8+sLRjxnOzslWSWtXkU8Sus830OiySAHWJwD457Oad7DZHT91qgBM7UOeJ+
mifZWRELN6RWLfATTTqCH/Jx74A/97FZxybJQvUk9BlmGao1OumkKH5kAn/vT2OU
VqPCj/mQhUImyLO5u2rop7dapXtbUZv4efn4evMb2b/oqy9V17p3pJAbNy7shiis
Dd9YU6lYwpkvmbgfsrVgxvqjKSYla9ogh4vIW7RiFD/Sqpvh7Giw2CWt0OO80nTc
v5Mv/HWWoQHsd2X30H2hpmCN2AcO5Fgb10GRSJULYg8kcVVtE1dM+L0JxY3+Idmh
2fYuo8eqoHuoOQgwHs8A+qhak6kpfZbg8GyqIAijG1huE+NZ5hs9RQ4gowaq3Etj
Sxvj6X+kdFBDrS+YSzj2ZQ==
`protect END_PROTECTED
