`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveECbcSQ+jHxWj9YVQw0bNlss4CkpSicaTcBQmLiIpmRq
9d7rySGKr5QU7mf0ZSsIVKMmCoJqHqlnLzjweqVpDhQwN9vwxI2DBSN+10eBZKE2
oJrPwUgWiPEn1DPYCCcoKmm34Zcp5S2qP/oFSEgx1LtAGYFO/4UXnSlQfG0nqxQM
E1F9OtsTWHFOqF7eP8/EEFxZDr5r8FCkf8d8H4IENQ7oW1W7PxZpyhkF8cXnDKNo
pFee8BmpyMJp6NgBo8H78rd0hYPzsVdgWOVVqSpln7e2XXdGFpD4DBEQDD0HIrXZ
tGt6hm9I3Sfi10GjB8YLbWL0I/wyvM8l59avxPD04vBip4m2WZ1YVBnc+Zb+NAhx
uSJD2ac/jIFvWDjqxeY4iPkna+/yIDWsniuI3L3LvqXiExYCnpRj/E4WXPOakhDi
oRnlxuklnVJdul5Wu5108w==
`protect END_PROTECTED
