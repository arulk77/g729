`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
feEC16L3KKtCQQb5jZNG2TdKGx5oGweB/Fm0weH0qSgyL1XyY7Fah67Zeua95yym
8Y8OqpIfbnx0kO3ulfYohTZRb58ScDjvIWPFjNFT4McDabul9e7JV7J9qc9olo9f
CsxHdef/ns4ihX/ZoF4aMNTqYp7YZkkWt5gAKBaGnl9cnw9f8EVLJieMIwRqYtbz
XDtr0lNGueRxVpfnvAQTfiK31X53v9HyQ0NlXQ49ZxYgqiQxC899y6xlq4NJm5ul
/PwILSW3c7wbv42MLdm8klcL5JanDWFzDTyXO28rKnh+lvj7UTiYQjZaby+pRs+D
mlZeH7D9QEWpFu6q7HS2lxb5MYXodin8YPog6xlhup4=
`protect END_PROTECTED
