`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j6JzCPNdlGrKqMBVAO1FAaVXC7ueY1WAOAzepc893i10HHOWIzk6PA8O0hbjtoZv
8JkwK0q7yMHUoPTRedklU191ZypwOTI39uWpgqkpUIBPM/0IuSBe+LMZ1MdRJ0oD
IRNVmhXYPGHj18yPCuw9tPlwW0x+lFizpGVrrqm6szSdyKG7TXF9LtYpO4cJOlWv
p6yFo38OP/BIvJ54ZAMqgUMEBftrkX0ctNkkrel2iYs=
`protect END_PROTECTED
