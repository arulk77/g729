`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
XZGW23JwSJliq/axJgycZAfJo+oXdFoFw8aNx0RYT4hSTreMh+TQ/MLp68c5CRj2
htwMpT224Pl2H1V1DrIcycd8r0+xQXtH5dbEFKCrWCMt9xi6NKMEyVxQsqgJ8Fqe
aVAh1zE6YNdtv3AuG5n7sv1/T7SUJX/gh0HLsbbEfoQZQFHYm25EK/+qKesE54e7
`protect END_PROTECTED
