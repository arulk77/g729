`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yKxDRjckmE8gyVqmaooxpYVnKf9y1ypeIFY4VVzii1H
EePCiGwszk5qKrr+o3W5d853jce0YyUmGVcHNoGkU0s0y/TNS2nIZQDh2vvtE9XJ
a8t+MQGuKyhKSHkVqESeriqJIwTLoGYVwZEBLQTLXsEla2uV5uQXdOPCsT17Oglw
Q5ABKzqf83jWGrM0nUL4csj/a0BR4/81DIppVMghUoHCO1ZtHnsrIIkBpfEyWuk+
oFJy4kkY29pckrQstwkTGO3qW95RMFHbFZZi6SoalcI=
`protect END_PROTECTED
