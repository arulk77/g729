`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKwa0pmQ3MiWKqss6PwMDN63nTj+61eCsOMFitCLLQ+A
WakywhVV2sf+hViUCckAIWkCvtmVl4jI9XblPE1q3TrSQZPiMTg+5nkIpXXX1hON
Yw7ovDLdZ5IfZyELV3P68mNS/Q3PQ4SHL6wSvgnJJ2N27v2SKKnh5G8q8DLSQ2yO
dowySif/nHbWu574xylyTo/hLqrbWL4uSpzgyZZ5/C8X76xyar0hFyV3Bqkmo2VZ
9hmoqstkIWBrNqOHTzFHLKAvW41Vq+C/vI/l2YC0Mec/1indUmXLaxP6OpWDmXkR
T7mHVvxzX3WDOu7K+xxmfbySqGyeGL53PVPIRK6ljS7l+diZ3gEV8ABmfbzYlccL
YGHo/Www19aK7s+lbxtxiI9GaWdb8+zOYUcWjw/X12p1uhDnIGnjV7NP1LsqPwbh
YMuf51w1Mg0d2jhxTu+KQkl+joisyPLDoAafJoOZcMSYpzaXCpnxliP2MzWbj16Y
`protect END_PROTECTED
