`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGt6uYOj9TLV5tY88c6nc1+EeOVvKgJHLS9T9dyR3JPD
KlMMAYknMhenVjrBQxv5zCvzTkra4C+5o8W8bfJwco2iS3EJYc8dypBF6KWKAJuJ
ww3JTQWj5fJoP3otKVk8i7fM80qIou/4kc3TD+XH/qQ55/JQbMPmbH1HgsvPVtWw
TyQ66+i6/p2HUPHhwrW6qZ2BkPEg5AxftiSYJ8Rh9HmrlowAzCCyjZaStVdpHmvB
Bb7w5QkPlKf+tLDyp7xF8w==
`protect END_PROTECTED
