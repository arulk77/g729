`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDqfaK1wl/M8PZTXpNIFrE5sHsw700sDNUaaW5HR9bIv
9KR4pie5dpgC50ybsCGMoRoixwLzT3zTHZYcwh3PhewPUdHWrQUS7BaEFQkuXWxQ
1kZGeFLAWwElkMTr7cZlcap1wXZ8O8K5+eFiB0Uu3w6yvQ3W5by8ueKeBUh0aZbG
Meg4jmgPIQPSxwNI6j1NsF0RslNUFbr95ycguAFD55EKQ+5vBw9H+kw1d7Rec2N7
3Nz/3ga+sVYw8CeLbGmTk4u75zORZxb7xunAuWGGIKEs6QXXhu6mQZp9z4+B8cP9
94HEKTRxFFHSMWWkepE2KR0b57xW10LVaVg0cdEfsjP51U1Fya0pOKQXHtXPb0nt
AYQdnomzGc/ucG1gBAneL8AdhCLw3eHIMuYJyp9Z8i5AAf3HcUt8xkthxalhQe6m
`protect END_PROTECTED
