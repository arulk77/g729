`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG8Bxr4Sf2L2KhghcmBfumKgP/rBBU2AeEABAcSJI0xf
DyKN/AnpkMJKPkm7v1D/6232YKLsaR8zeut2GKYgtdfOAwg6+cFFgliiZOzHmmcy
PPumSeGwWkqdDcAAWfZRLB5plSIgyHAucrJvHGUx1FsQneMGWs5arHPncasX0dkl
ADduczh+J87w5IeYTIM00CqyR9HolshrgYh52SF0lZXF+VetJirOVnD1qw01Z7c4
ct2YfJjUem0V6e2eW/7qSdqRtjYYHKN6Rgxc9mkAnPRCeqy37Bgqos/HnQSqChWd
fKqklWfALwy/lAxBeImLyUtBDNF3k/wKvhCWZg35J3yexosX3+hKkQKN2BMB8H1l
Z3tmfkozOj+RT71WRDI9u3TRZqk2G3jEO5GbRXNHjMJ5jWbuOZ92YaJl/6caog6D
Gaemqv5k+tkFllbHnT78DT2I8KhbngDJ8GG4wAdIH+IgZHoBsky5uFbS7MvR7Z4Q
L89NANCf5sAi/6QiLAHTjv2X5TpaUK3VYa7oef0Y3MXAyQShkgUmrfSwvMAU16qQ
llDOr7VMTNFapfz3Q7OoBvv2K2sFCmWYIS56bz6F640o1YK17XsZjQHeQEOEb1tm
`protect END_PROTECTED
