`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNwmmIN11ggJS9x5U1sDh86ahhN9vx/TSLQmSp9jGTIx
4SIr74D/FD/TjHyCosrVmUpQYy54dlHF3KOHXjQ0Ojy9pCijEZcVD9r06C1sgB8C
aIscK71gGv6Sm6xc91nBk/aLRG0vJYfVuRTIlSftKDXznIDjzGgpj1TM4sNhkRrq
bVBjYtrToYgH6Lc/BfZGMHRkb6HtQy3TM5qSd0qSXfXImkk/KPYaLsXi9LCR9NBU
3KTEUMrX84vFoqTwkma9vSQpqDoiloNvh87pktHs5W5GlcSBToqWBYqJ4Fo1Ieo2
MLYdbaA4whBThWji/dZY9w==
`protect END_PROTECTED
