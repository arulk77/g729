`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePMAUnsRxnkDeFUEManTqR9/28jtwGKNZLZIjB08Oode
eDAirwwy/0P7q/3MxpvKoTcznn2c7JszgoidAGImWAqo2PHdqGQzcjwn1y4qZ2Kr
KtIkP+tWslep2VMnE/g3G6sr7GMXD5SFN015BlXQvgqTJ0vO3o0HU2mezf/QNoko
7dlaOpO+KO8lhQ2TNIRv3iQU0v/pJS+zARnkGNhb7GMnArQItf7wthBkvMagVxCJ
`protect END_PROTECTED
