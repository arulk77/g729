`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM9e/rpVJ78Nx4Ss9dGifB3v/uYSYP3iMsU56GgnqVp+
x2C8mJZEjzA/SonuASfryAcozdgGPuE6FN5DMmoQRpxebiJUfl4n9XncQZiigWpz
pz2H8mSZLKkwM9YybUqHh0aJo4ZDnLaQBmCEWWC6WVMxIQGTIvhJgzZtTFNZveII
+lKArU3IKjRFmkLDk8AsTcy6FdvgM0KOXoMHDTNO7MuooJLp23B7i128NUqupQ6g
iPGVG3iKtbiYH+D5n7k2f01o44hc8x/Eh/WxUYO5Qki9QNAFq8fx6r0hMZRRSSEX
J0RrS1EJ3f8gHNw+tnAnEN1+ZDLWWIg95NpLSTA5gM8J1tf/YSFHK3iT+Q3z6M9I
1yWY0BGTgw6/6Bzw64hwinrPAZevuNMkpjQyeWlX3licD7JemZfA2P+xY+phOsM1
16A1UDwVx9jPPI6yOmPD/rEtyeApFhOEPKH/PCuKx24l3qgZd3lZ0gd9rmDnmuIi
fgSR2bSy9Oe4HtbWRqO6qfLYQnLfnRHAISVLjgioCqBgbycP7mof2VIERBsMoJYS
wxrQ7C+Q4KGLNSGJ+cgdCPHuyrkzv4af+nCydnBdfxUt4oyrxCpg8oOa9GzWYjwo
M4HYoJeKnGfGA44Rn/Qm5C8HrWSsPf7WyxqU3gRmRntjbWjW56kbazFgZPr+90He
kCOzQ+sRTL6aeOD+zQfclAhI6JJqcMI1LLs9kHp3q6eemHBvV5HMpgTP03EgAQzZ
i6vkRyJYPijwu86XW02lQ2rh/OE94Sa9nxteuTv3NsfYUXY+erWVkjKI6uMTAVpp
J4ph6639F3gcs4qzayjVh8P7z3cUTVWq/wZZ0r5HyJnp9ipM44lQwels7bSPnbBd
G8xoi8bIr6rounHqnRf3WFpxIB57FShlmKhzSbkMjVikE+OwX1K8oNZPUiDJ6FUf
c6xEkp2bIt2zzFcKz8XhNQfzPEzCWdKknc84GK4JU0V7uHXbPDuTJMmSA5N3MLOg
I1HyL8SYKpk7sq4/ZYjzjKYVzZexQ3tCORl+ulXCTLy0DLrIYDe2gQ8AEamWfqIf
2DGvOOQfLK8ujKStgSR8GDOAobUg/s5ud/2anG4FwluIIM98YL9BvCngwJswXRQ+
Sthii3PDGR3SpjqZOj1aimPnlsZgeoTet2FNrFD1r2VAW5BUjBK3DH4Hq0LmvIsD
57WC5GEMOxREkij6Yd4Z1HOaOM07+L/eckO7cX6/+nepCM3/J2ZColY22KRDwMGZ
bhRC2D0b6PjuvSce1v+SvxE4a9/942o7RiybwxhG30sTZiUbObxbLqsi9Z88D2xu
RitICRzUlLp8dQEPT2Kpq2IAk+omn3De8BNzVghk4fRE9e/hYbZuxT4YHFWKxFkE
zCKPLTr1QXUfoU+hbq0DHEXk5X6jTo6R9D7jw3pl5PJ+YQcCZHk/zPkgq2gH8UE0
Bt7yIxFpJH9QyOuREu6SVHqQb3jp1rBPQMB3rnsd/QxhNarFx1PshxBRhW9CoWeQ
Z72BEefPuf+V4Qt1sEJFpm5RedgmohDo2Yvf0lduOFJTaN42PRwmei7s+HNbzA/3
16aTOMdI0Pf/sV4brTbx7a153O84lsKrMywAAd1MNfiSV+KgkA402n5yj1+NPLi9
AK9hfY3Mn+AAHkO6CYQYA6GfyDLFJjlOiNcm2CXLxY6RCTRtHvInREVloJVWnwug
76Fxw832QVXcVPq3iihU8G+wHLvihFiWgF6MeThIuDi84OS5XQNfIZ9B1YIXqn5c
QBesiGcWH8YZPo22VBSs/zkzy3EsTZZ/j8IuEa1Vl0NxDIZYLBdNc84QlgUHxyZP
mrAGAcxG4Gkh++H0Gpo2r7DVUqWWdNMxgAInOO/O56abNd6FLTu8P5PeO1sA7vNd
3hLYeh4qdzV09e8+NfmLbhS/RJMn9zYj36sZzudQrpi3pQEiwsM76GbxFV7Gov94
r/uFBV6ziMSfjlqjBXZHRuzbpL+9CYBOCCsI8V6Lr0QkBohY8ptuAMi8bJkaG++s
cQ/nphB9F2re+YksJo1ZiDIk724gdULsuldzS23Hn3DBxcjX+RBt0/ttpEXumooa
IzAtufetpcabSrn0bfm/82+4kQ3VJNCnsS7qPdBe0AoJk4/cwhIPXQ+A2b99LHwm
OSLC//fsT3pBz1WGolUTX8LGQcoo3aHCQqcq7OnIVEhhBqVbNmLth+OEfjYPIIHO
tMLMdoyRGr+yS9by5zxgrRO8dSnn9OoDPmomQzoqH43xycaplOnnNWqxdpXjWuuL
E6FX/zYmAJXHUPGNrG27PWYSas9eZggh6VyqBldTYmxQAsiKXk1IpEku3x2GhYkx
pxKMmSuuhltHq9PGYOmeCaaXH5XL2qlwItVMOX39JZwTFyD4Vyx4yPsbqkmCSpUp
jiShDYvErtu7oWIOOigf7Gyoof3JHCm1YTzXr1nmPerkxq5XeYeC2arL+H64Kq1O
w9cg+3EfTTTtkO54sAz2s64gsCLiJ1M2alO0pVC45S/klXA4eOeJFkX4fDoBWLP2
QE0CyLCJDbuknpXCkrafvF3hjkLLgrWwji9CfLoJrmPx43QHG6VzIVG2/WDjIklA
OiaCLFvK8MQvHBMMGzUDHkgUp0LUzzADgiWERdXiY6+GiYKrJBWtHGbqLNPsRFMf
kr5+j1YPz81iL16b5mtfbZaOiRlnhZPYBNsG7v+mFCnYxEC0sn3A1WYVmJf0Kr44
Yd/P+lwep0/hauT0vrDCVwistQ8Vh5bN6rB2per6Wl1OFfmBbfPBD2XGqRyhw1ri
19TKMK+byhFCH/Gevt7sCHfAJzSRr8HkaeTPl7ZJG2YdcncU+i6+oyWyifa5DzuW
2sTdhzjG1vKaWznwdbiLF2jDRdIpVvBNcVeldHL5k4IiNfjO+2udeUbcRvsu2tjL
LuVKv6BrL7muNUk85lyfqpWfgmt+xjUjGijWJ3acIWO+iNqYzzPYXyD8UCaZcNEJ
J1/LaTJDDirbTQ3SKPeBuExp2Y9Pv+l908GoHF4rfGFucakTH1CGTuZ45gtFo8ij
s5DA5N9Mkcs9ro/s2wNMlGUJ9XzlCNG26tVaKMmNxWoRqz2oH2pdDK8X0npO8lG7
xV7dC1B3mY43gSzdQvRUQTc3av4t8Cxf4u39KHwWrb4LY1ewJ8Bq3tsD6+MUl1tU
LYfyXPhtVRalXULtXWpdPr+RzGc8DBbfZBhegNfEi51eMlyG2Sq7wcMgkBvSaJFC
buAlabWNbmtJsJ50YnyfIvMIyqL/GZgFlm4VgPsSw3OyP1g2ipD4fsBUTPpgXCk8
Th2Qrz8BB8mhPvBhfyQGDprmktrPggaOU3sn96FLocKjbbFjckWDKJiU+Vq6CRPG
FfFmbnowvJHsjyulDhLh95te/JoP03JLn4GCg7KUInycvvkpWHtBnRr3rt0TucBQ
GAGFnhuWIy06YQ71tPDxhT5Gx029bJQFuiEtDKnel6kb11CvVTWyfYGddapGHZPQ
QgVK0YUTcONpwR3t56E99t3TdK4hvtesIqdrC0pQ71+bGXGhlFcaaIPn8I7OkNLc
exX/AiBDX7JKyZqBy38BseBugUwN5g1mgqUBFB9nYezWzNXyD2N306JgUpj57x+M
f9cksOyliSR7GsQrJcplQTFmdXcGBEdYk7oxiiN8O88JZIZVwvuK730m+AKG+qH+
FgRvmB6osER5KRtakj6CjbFqJBwl/dm9HQd/gL6Uv+FUOpYaOwL4pF7i/expEDEB
AckLk38jZZL2dkZmKkMrQwosu0uMYrp7fTGsFLxU+lR/Cn50j7bJrGC9Be+Hmno/
DQSITLHBuTLo2SOQfeLIJQX2JhGY5li64FWySXnSOAlchElusQqvojjfgBGz4gb/
KiEvoIBQkcOhQMQoB64be9V37Qfd7N6Eqvy4aMKOH47cmu2WukOigec+0Bes/JVc
7t4zO+XJwbP1G304+n1BmGxszbzpRgQLMrLmYRcp7/ZmbCybLvfhpn4IJMGs+dJE
JYWARnF9GR7dslMCp7xAFHKjayruhqvltCmprwUwqDcrxsSDTBNU7rAd8LngsEXE
4PMlkQ6kvs7BejmuMMpc7DBXeByFYJZQ5NaAOYPKNTh7mOp6PUyLcg4BcA8rhj7Y
SwHEG1wCaEtJ4Eg25cz4vmQIawXYp6QeemYe2syV7+xpu4uhIZe/UqmW5GQ4dqvC
Y1A8MLvgMHsJQjHNzHSmMJ/GV5/OULvTrhPWELgoja1ZK7VsNhGaQzcYTOYd6Lf8
ak3LI/keAVUq5KugtCtVbkO5INeJU4oLHLLTVb7x8E8Boy9BB4BJL5D1yQwhjU1u
1pQ9e8zxFogoFiTzvCYXXQ+PkvSbi3afLj3bPxnZpToNIVlLfvcfXRTA7WJ0Uyas
CUj1bcWgGtdJUle9wD1wWqT7oYM3oBDUu+pxDSbGnYNeDI33du2OrJYjc4ehUfQK
ee9gp8xhxUSa5iaZPuA0DOhQsYSNKKQ12zrO6DaEh3TZ2DTpmYl6+w5goAtH2hvV
6zZPz5XovqCab9jFpxqf8rPcaxoqYf9Na5LtEqnwOQhUua0qaU9jtkqlM890Y6F6
NF6sxIe+JS5X+/mTyd7a21EF+80jMUVU6/Z55YS0PpByEwIsA12cVjGXETXCoAms
FEJMlQ/6D26LYppeToXmt+N550GV70l2soZn+6+M3xEI4pe8CvVVUdQyWcXK+rwq
XeI5ZcwR/9rPVgFeWFAG3LjHnWb1vpO7wzpK8hiB/CPRSCE/ZPNGw9CLdBz5H+fE
vLagE2CHjaAi5W65sArhaSUV341gNCYUbQRvX754wZApAj/niWCNIoaIALPhWUR4
cpNzWld3qP1B0hddmotW0HDOkvLqA9MUtkhRu27RBepv80kGhU22Xc10euVPuMje
dugOJDiS+Es9JaugyktQIS8rjZ3+C2SC9vtuwShN3it2fKDHnrL6asgjM6e1UFKD
H5SVTg2kdG376R9L/XTNdyv6w+JKJRQysygT52IUmR/F4dcLOhZOLdT39IkrhQyX
VGFqlCX/LwpaxsohYAviPPszMxbNNQiGTFYDhWWNhiN5tBQMHXBtdyqjB3mxHFy1
3gij8IiIZ2kNEEfKmlKzGjSrNZeUxvmu+TPI+xWJuSX68lB8hGmp/rlVPPTNte2q
lkM5TD7ZCto/G4vSIIePLgvf1r5vdJwRWTfhz6nyD/tNvp4Uz/ntE2f0hcLM22y6
rl7wCzCOv7gdgBCPaIx+Hw8CUnEgr3VDIamSHGC7FzNlSVvGJO7u7zVF/oaz65yN
PpHiKDPmh2xEbmvAzgkToYoOjOh2GIeFfZerxLrBPjt4o/L/8Wa4fkxFXsjKKuWl
FgdmYg/a3dq6YjsIic9DIz8aK98oqXJm/xendpnaNyL0cxFdzh0zT3zrAOmQrIWm
36rHoFjs8eoYCOBowssidnvFUomu+VSgTtQi+m0RGYVCEEr+fBNBUFc7POdUxMrT
J6pkrdWFt6RfRyv5UMI1Ea/WAsmuN3ZKM26EyzFq53NozDASmTJMFVw8TsO7/Z2u
czthxVyKvY7Wdu5AGyT9tam89Mz8n0H8IEuBc9I+Lrn4H4Vj4L4B+IkjLGJLxszf
IOXiAu8DXMNtRi71ZsdfAhTjbpH2bT/Dw3a47oWwk2HPhSivJY0VK/U2GMlbFzBN
5iR0UnJF3bKF0UTADsmKf6ecQQZiosb8bW5PJ3WYQZr3wQ505Qan1trH4HxF2xHY
QPIMbygX758q7sNrcQeTsqM3KQAJreDrwRDIKwr+p1KHl4yzKTU2LUfD308U4bfl
55e6BvmgeVknh5M5+YjlxQuj5dJqMd9q29EnXPxdEIN3tdmdeDe+wtBMWTStAN4P
UU+q7sh5Xt/LR8wFhcgpgbLmSbJZyl9EvCtugPVq18tjfalsRTCMUNGJ+By7oDxD
FjV6jIc2uN0zWLPS6VQ29uHJT2rb4YcABcnH7HZUZJuhI3zIXkyUaoxANCad5rap
aGNb6qUxXt93ULkeauw9vAZAQUTR7AeXi15U8HNLORJxrqooP+87V/EYzQBN5jK5
/hzGjCeOqRoFozfC34ibJTRSbk+1X9WFhHni+cdPThQBVWA48bI9C49l0V7DwaFP
xinJPNF83s/eE26W+L3eJb7ZyaggjhrDrko1T/Y5xC3FDQAJYLVYJKnxsqgoI5SD
/kZSpaJLHkeloQ7vf3HYV24lrQyuUbdETXwU6hUQ7lAXcyEyHpcAwW3ud+1G+vI3
mKlkuw11EgzSyNhU5bPBNJ2NWJQjdhVKYZo4bY3HQCHm/hY8eADP9cbCM7yR+24G
o/J9dj55INZKhCYHqcHGvybTAIp/Do7Dfj5iobWn6kf673zCVBy/7VIiAWfUXUcH
AQwGrCsV8rvbb8ZQwKdXzJxsOBF/hjRjlfwq1KBOWDDaWS61bNztgaEYLbnw30uB
r4tZXOD+xFO6mhFVPOnqdA==
`protect END_PROTECTED
