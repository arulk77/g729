`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDASbOQKne1dLEmlPs98aIaTHYJXKTpVsI5u8Ep8z8v0qL
S3ZP0vfIB+qQW1IyNaK+fl5IDLNKjRM/ZLGWqVdoQSKQVZOPJnMEpb7roXuAFI04
Q4i541Iu75OhdZfGkxl3gAZTtV+HdffRzUDtVuA11GgsG2IrBdruV1+wxlIRJVjw
U0o4tx75DilHyefdnfvVrjhf8glyI4E02xwrWk4WaqBYAkHVwTCL8s4NkPCKcjJW
GXrx1JoLCGaOPswU9buKRYK/l79eBvqmZlcPjnmZB4FRhfMd84Tsvco0/2AzsvL4
KSTU7n8+0YDzv/UjGMcyIEwJHLdwotgH1+NVLuKyGNJ53S/v3lCfdQeKlRNpn3OC
VfOLjijGC8LPBP0iSd72pS1e7UtXumdnfKBUmRoDKCJoOFoITyGjZ6jEt1K/LWfu
tU2HjuWpQKqjEKh4y43cATLhP3Xw4giJ/j1VdfYkzMG9UlV4wwft6Rd2YIt+jkFY
StIAkg+ON7khFo6ZkWgRMOwd0u4UktfCxdGxwQsvRBfnDCO/11kua4qLbikT5kia
VHpdSDvzImB4FmgLTJFzOrt9F6Ux8TlRM76pUJ5Vz170LxHVoAU2k06lDGMaFW4H
f2ZHnRVTDhS4qVGTpk7XBFI/QBJzWWhWAi1PbxYststjLFUXh/X3SniBi5g3OcE8
CgAfinnB9yjRP7Q8ixPUDUXwmgWs4vZObM48DORHhzOuxfQUJNbu8ik7OS3OtURk
Uv6B3goB5wwtWlRdRkJmjdm1/1G9n9YXTJwAATupt/6G14/UaVNnGxm6Vk5F8dAB
ZmJiFdpYfxK6XIfRofBECQpdAKY6y6oZToCXqR9TYq7LsHI1fXU5ThvFFFL2yOEA
lTVzzM8i0c9gDdPv/NCJ6XUZZqDpk80YfEK/d6/EufsrA9fQEJyHKPzUKNY5UTmm
Tbj51Rtw5/WDZ+JmjspTbYtsMPCVYGLHkvLsGRg5dlR9mh15FVN9ehSf5Jse1jD6
aipg6/wv2xiAny8uemYnvNqF/Z/HVU0eMUaAicd2FLw1yOrK3Nl/6/QwHh/NHR08
m85fYCuJNEGkT+uuO3zB98KQxPx5kkS6xbQBXZPhEEE=
`protect END_PROTECTED
