`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73CwxSCz+pr/QfkrYDpTis3cufwQJJGR6mpC4uz6WHth+k
KSzJTqihx3mxbqlzJ2V0ebw9WDda2+luk2WnGEH1ZaXvc94g//G+ptevM2Ehrg/c
7ujGj1zZhZaXxCSHm+TdsZs2EgWDunBgQYjwZFdZoUsc3Hnp0oK8KiebEvq3wWZe
EaSGmd9ZgJqD3rKLWsgp5NOrPUBqZLrjidetZ8m1CF8echIItuVYqGqXv6qmL7F4
RjUmk+ockwVzSekKKZNgVVGIfM81n7A7VYUPmjWJooC3EeuwzyqGw2mheva1a/DV
KAZkkWxrAuNMuEZJxLJPpoU+G8QZ3DXL2Xa79u5JeEVjcdbLlOGJ2GkxlRxseHiQ
wb+Ng+UJlGxOGTblN1yFq+e+3nv1Gmk+BKSl+Fg/RUW3fsI/c3byc8qyM1mfq8/A
e25e0UFu+iJculVlZHymEQjAWTvaHh21lQH12CPpaYE=
`protect END_PROTECTED
