`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFNQ2lkl/aVxkTJvHwKNKdc445149IVfcS13/ywFweBq
rhXOVHmiHV5OHKUOvws72LgX1dUwyLSK6ZQtSzKpk/s6Yu3oCFOgyO05XTNa0VeZ
5W/tIFO2wg7AqBUT2BcvBnr6ZdtfASqQm/GmskPKhzJkCfrjuHIva1h2RMZGJ4+d
80K6OZl1vdoYYafsNNUhxg==
`protect END_PROTECTED
