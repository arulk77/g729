`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3Igf+CkbYUgsJFxMMXt9Oxlx5xDmTqr1CM1efq3fpZVfRyQtYwWweFq9lWgXgRoM
Kq3+b7eONB6b61WqzZnp9neEgR+iYk6WiVR7E9y5BPaZJp0RfkJAmj/vf3lXNQ7x
GkihGncvojSQllnv35VqfvCk0XIiHRQn8mCLM8swnVJmvZFLTzK9zcz8Z/ZxcuoY
`protect END_PROTECTED
