`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SY6iNfkctd4ejYahCTqNPXsuKYwdYDnJ1znEh9n814gh
N/fRYMbcvuBpUmYsw0Sz+auaijLkOns2lmvT6xRB9k0+I0CSHAJiA2uuJftwtkRO
ipAUow1uAi4ErgWRSztP5OQpVYbG7RwwZo19cUQjpvWeWkuGm4jxQlEHHf5+8u4Q
r0jAGbYCnCLhNxVptlBfHWkkoFk+iS6UhM4NSWX9o3LXznC1YQhTeMmFcpLZoTeJ
tZamdyPHTXsg9WJtc0q2W5vR9ro4ONbSt5aWBfClPdeeqHMMY/lRGbPAhtZ7cX3V
LQOEs6o78m64RL2BBv5JJm4RartXkJMdvdH6eV0F9FCVqfT18A75lCVRDQIYGWvM
tAR8CPuFy2qbOkJHiDnOGp4MLdImXlw5qk/n5vbEARJk0iPqXgmgi58xd/442+mL
VPAjaXdlhKQZ9iL+652xtuHCDMsscd1/00TYW6UFwXyvqsU3wSL4gjMSLUAedUJ0
FEaMlxvpncHhBWBMDLXju/Uz27lC0Z5xFUZX3yoGPNi5VcSOuyvEtA+G3iYKfVZo
26MjKwl4NE+GbdKTN/7xpj5+fAP9NExI4gwXo4wNrVFBtDeum8osi8yQeY1WvibU
ofGJSLdUOS+uPeubTAV7NjAA0b2wczr1h6wqJIZReS8Bo1K/rgq6QHa8wLpPxmdT
gx5nCZfZncutuVNsqi+apWFiDJkbAdXAmesaZbD5MBozd3qHFK/fa26fxKOnpcTb
opvxdsO/OBCpFp9QbsaWkLkIdy6CTllWkJHKYd8DoQpV4fZRLOhGpDO3Z8aMULki
FfJQA5cT6nkRIZZwaPH5KaeIJ9S1tmQnyT8kuHo0J6jndY7wJ541FxJ4mA71utQI
`protect END_PROTECTED
