`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41Hb9FGNMT55lSmVGrmAMNZ4onnb9Cc9yPerQXRAuYYS
yV86UTvpp68kq2QgBm+c0ZKazQ25DGHB4FBMy9IiIaxbcL7V4J5FMX+L4RuRPwOE
bfibbD+N9XORhUmpAW83/5tRNYNLAf1NwtvHn6FCG73yqU6dxt5LbVRnD61na0ui
NKM2rTySqzHKj6WDHDsNCbJ7WwRZRd+c5dmaILpr2gvJsm2o534fOAD+6msv1B/y
77y0X/DYPHLYw/jH9VNbXKFvvRBPOvi5vKQXTUBvhF3BnpXeG/lqBiMQjGmVEO4E
veB/DSJcNg8GgC0RYLAqLg==
`protect END_PROTECTED
