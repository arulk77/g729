`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAaE4xZ4/icDbOSL7hcp7YaW0qksEvD9fBwuigdleLBOT
cQaOPAfOCkD6OGGqO31rcGehEYr8lV0Aj+xTbTZ+R3LTYM36OUwFbjUkdYfenH/q
RM6WaEugAmXSV20SFlUGHcHpHczFW96VJwMi+awhXxtcp9yDQ3JwuDQXARPmWTSx
Jj2NT6EcqNZ8eOoDvvwJ/72T3vTmlCac34A+qW2AXJ9Z/BDMbYF5nu8UV4VnmzGV
GI2pLdYFNUT507TjSMXAhl4W+Riq8CNmc9LvpMtxNofncbognZL1uSEmBg5Oz5Hy
rZ4Lni46athzkw1JF2aceckM1WYtnVACfoI/h3nVAOauiW0hX+Pz1e8BOoh+frYH
zqdI28y8/HQkCRkQ3lfIdxWctjJsH/QXMV2P1UyvD0dic+EIL36HZYROgcd8TS36
55ZmUbi0lLASz+LoWKcPN6R7hKgUPZGAc2GMrYe9fjghaS8zaR8jrWSIq8vBiLnb
jEjLeaoCf77DlV42ZJXwOjLCbvStTulWIyTpsbnaVs9a9qfACX2IVmthF2AZPdjj
XbHZCJhMNs2w+ZuMVHxNzbnU5VWZd2kp09U4v6sgdyAeW2XNnRNTOkjNvd6Sa6EX
3amkji96VBm8pLEkNRF/6jYVbkOEoGUHZiyv9oIROKLjHOV9dyEv7rqCG6xo3CPw
YJ4qABTMZpTRXoxZqGf/c6U6YncljAVEnL9WM2Bj/uiZibpDxCgJLeNR5jKaAhLf
wB2lCyaWcbPUisb072v7M3G5g9OqGnxVzmcYSyoiRlP0+FHpLTkldPy0vKoXO7sT
kky9AE0qAhIr4K0adTtwAsAqmz4yTKyP/DowKja1Kt6TItX/3gboTPENeEH8jDyr
rWUvgiHkELzhBfvpGIqwonjII7ncR06UByjx9MWhAmRvf295GlroeTQigmNYPQJB
syF68ujXF27DO3DwmL7PAM47NZxcGzx5B/9K9kKxpXVZkykBkrT3R7Y4Dfn2xTv+
kfzdOayMfptXPqqReuhKuyj78GVVX1NSH/8gTTJ7mJ7AvnUQ49qocHWT7GOm3dEX
GoMeiXSS+J7rXtohsTbqGvD6a5nBAhkfYwKIkkIdn1OiCLwHF6yJV69eS7vBLa/w
CxOfX8onauwY0/MIEgkCnKnvJ7QgmlRQoJzZyZp53H91ofJc+CGVk3wyFDYxRwV3
1Q9xs35b5ycQCG0/+cfmIS9p6BsZwwqYA7r5NyoaYWKqi2ae+SQwmwWTGd4dy6Yr
Nnj9H0nTZJEeKkPhx1A5w4s5qw4JEAkmapR3G9MBPzHj6jC0eDnQhlz4L03DkkiP
aD703SMzESUill1E+kTkqYw+r9xcMz+Xq5m1g1VtOJIlp741vxJhtso0MZIfbYTC
ZbO5DIemFNwe7HobhDJVmz7aRKtDKBEeNLM9fxV6kQEWaPl9tDU4ZCvc4c8Wv9ye
zAZsyNjvVYBlSXdpQ4V6M3p751zci1JdIoFfQ2p/izF8JcWZendQyqFJ7JMd7n9g
StdnE6z71egTi+gsHf9sPHoFXYGHKWR2Dn9ATZhHr3ngG1xgm1ousmsyvq8l0WVQ
2fEgDNvXzQk5VpwX/fjZ9Bciu7yL5xtEpWbDiBCvCGI61zIp0kx2XkIAEvuqYE8C
TsuwH/W76tN8pOBuwADPHvhxgs1dW+aOSMPzlP3nj9QfVioRiXeZqreTiIzW2tUC
L1aI2QAtqRuySkIsOmKF2XuAw/xH0S7echFYPZeRXuxvqOKF4jE6Aq2aqO2A43CR
DjeZQFnEKlz5uVrR76JL15PoQcfwZjM1iBDe4gDgnyXWTc+hjXQzGrI+idH9jOC1
RCmEmhzh1nUhTUJt3UtzNNXSe0oFgWmmS+3kBJsjIexBHhbDAoySs+83ceJDCqln
9fYkJ3Qr/4C7u0Ej9+X7elGOo98cGuK7oPwZNrV8m8BF9/Ud/g+n2gkA/ZiwTEAI
V1smwmZ9sehmken5vz5ccf4nWqmYNmhwB7Gc47HsGlVRtAz5czHfMZOOjNgTrupD
mTOhUDg9Dj+lVJnXtRga6kkX9DKNGoUn3SbC8mbYrd8Y5IWf87quSS1LnDeVmLWN
hlJLPhXxm4GOD5AbGMZLwkXF0AKFqZPB/0XNNLgN9MYEvvgZ4VZnCzhOgVkFC49e
WbUsgBcq8uBtIsQX/nx9gajiEwjTxjm8uuXHBPgE+q9adMy4+xRoja9M3PSYPK8J
VPhkvtsMowxr3NKAJdawatQaSE04eddJkqz1uSK1+K4WiSK4jMtA1eHFwOWk1Mjf
OcVUF/WGDq1dyspCOd3fTlIUXu6oPY4dSDKfqeLeCaqk7RV7DXFUJ11xIfY/cXEs
OEreGyLwTyvKj0/b9LS6YoQeUtpTifwlFzXuVzS1kj7UZnOxO1r1XD0dBCum8Cy0
37m7ph2FYso9PW+zjDx+5xX13Wtfe8DIl8suE3S2iFeffLZzuxRifVh9RZcsyOng
l67lf0I1VdgJHR0Kf40yOg5RmcNIx4JX0ZKv8fLhSIR+gPTtALRt/NF1reE/vWvK
ctSjqCZJvS6H0YxSFfPDmTEY18UYGq2aW+zuq3oci0aJvOE7USYMoKw+HcnFmm8V
C0Use/J+4loRbeicAJTl26BKXecvNWEwLphUDqiVnLQFiseejEYhmppHrHMpkSP3
wzBUhnoNZajfWt8x6VgT6PwFpQ8DJGf2zKl6yiqx9ETgmSlH5qs2Sg80HGZSRf7d
83EIXiaZtvc/UohPpM0CeNPpwIjVWPrcUWhG5RypWmV8mH4y4CXmu8vrWo4BJub0
xIkr2VIdXiIU4hXZyP3OYrVXOlNEnX3JUP8K6z7lll4+xowaciaxoSP5NJyTf92l
x1PMa2OoABWr8ZPWpaB1zZsb7Yh9oW9zh9DDl3gMJmR813ZbdrrOgR2jT1Wyu1LN
RKS1XZcyss6FlrgjvErxX5oTGDsmgMUyZQeOAiLFfN6F8DjKK9EBns4NBWYHrfIo
QvWdA90pKLyaBgP3f7fVrZv0xNj9rEicWF4Qm7LL3u/iOIca5f8Q2EHZ0wzJIO82
wEJPgwZzpT+sd0cw3veMV3kNhGgTpXp4QzautI7E1Uzhz8bppOPP6ssaOaIVzE0X
aAAqedn5NTjQSewfx+puDcr4AYjsa7dZGssZIJfbNGm/UoC2nNfpB64rp+ObJ/xF
8Rk0q315qsZorxoR2/QKKfPSlWcLc4vUqUKxY+cgBCGBAJIjIdKhRQWIbNSy68g4
rM9JoockH93caAlY77XcwnQiLCDlfm2U/YNBTreebskWfzaTpscBR770i8zpP2YO
KwQaAwuLZkE2OCwMvMMp4sOsUg+S6PhxoheDeYp0seDErnlDiyrQ2Sf28Aka9Gj5
fq0kC4J+MyE2Ou67yK/NIcof34L3uqL9k866YUlz32gxyxL/MldwjuxUORgRCYFV
Lnb/PmGi5io/uwz7a5RgSpaGbJJ4W2lUXeg/wNNDWASsvj99Dr55VCJ8W2BG/X6F
80sY+Qq4/FORxlG7gQ8S3PMxRjl3K3axbVy93N4z44JN7WW6Kmqj1LUiZyl2xT5o
5iFmSmG477WiwxWurszgA2Jp/DDpT9kYo/tCYMvFK7eWL4xKLqoDvBcTly1dnFpk
EMj4KOGfdXgYymaSNOwb9fDtRd8g8ZaCSBvatrTsF960qyywcerG4QXRJuSDyKKN
bDMs2PkGuC9fIB535aiBgmAHFXu5IwltJckpHKBc+XiekT6EWtS1NZqleBeU40Ki
GuY/5+EELNVg9dHzx7FYU3orCF5xmVUD5eAOPgGRbCiUIV5UHHQc1OmN1ZbEgxtL
KIRJaac8tO8OTMwbjYqVHpQRXcn3kLZiUymZy3otZ/Fc7OdIvwoXteditVFrQ0aG
oPDnwgeIV4RnesKoKMjGQODGlicYCculyi+jzS5hpglVGUqReZ7cfq/ovanAHluv
m1eYAfCqG80rItrZ4RI58Uv89PpTsQJ2xspmEo1U5tvFUFqfSJA26SvgW700a8tS
2/iFr96YkmNBCzV730bQy6Xea2NB4WjKmY0b6Cx9dbO+ARtw/ug2v2SIInOT0+s4
tzMev+jrcY7DiWjcC2DjW3NXnnWhXeywVoAZv41gvWLMm9ccvnopIZREnEbU0ucR
79cCMFFWA2qAa985yCRWO/4yrQb8bqC8a8MS9hd3ZwdxzzedNrKlxj/cKxbmMGC9
EZJpdeJyOwiiXCF0Q2y7cP/iKHokZmjJ74JSRSETcC0jCkL+CMI5h1P9Y0JDRHS/
7zSjmXipOd14ZKWbqQfD2TTdE6pW4MlfycYiuh2rcQ76r5nnZX1PCO+nm+uApUT6
s6TMEeVj92eayJhEkPqcA1WhVaY4rcq2avRJofSELvjvsXmZwl4ygSfNIpuYIBOu
BR0juDDxKKPHBFNhC/qmw5ZKunMBXnC96fKDSRFwnu6Y8Rbb2Tn5h4ZsZdx95J80
seQ8eo4W7zT+g6yE5knWqr7i9dXLFh+hDGmr3stLCpFjwBKCaKL7SkcGkO68f0wv
pRX53hPn3Il1qr+FVbNl6TnOA020+WbxQdn2iU7OFoL9XjyQNOKSmhBbB2TQiEVA
GNICurg3hS5sbfNCpg4SNPJZ7UzD9EUvisKZh40xFojUfOGFUM97wsKVkXnV95vl
jqXi9idz6aeA1Kj2G0fO5ufWNUxj3TwsTMgI+xuXi6QMKadxLoLbKcfkrAir9xkY
fnwirWTbOdzCSpEB/SLmJRG4JEqkTCO8NzRfgOerxYyw5hk/2PdQDCdoJidlQjYS
A69zU4zl0utk6iCo+Sa9kpfRdQhMD0LOSo44QwcjwHkfVbykAQOwEwQmftFKk7SI
VbZxJxQLd+HARv+SgrvLlP1s6OGnld0VHx1a6yIp8qXzY9zqha0bJTIh3F2NPbAQ
vN7QhTeFxBEnABHOUAqd2QRRqzTZ1W8WMz4K//Y/p3wBJ7L/PtEdzNBkJn0TnCCP
WtPyubzqcp9zm14FdnhtuFB1Nhg3doLKzcGHxVysU6o+5JDsLmBWa/HGj/y66I4R
PSZwVfM/qI/a5z218uw8RcxhJR5vNw/GONj4wA7y2MjLEOd7yPoh8BbXNBOU4men
osU6c4vbljYNnSKq1QaA8nk2OrOIOu9GXNULaLXQ8hryig2kjzLmCAxN6cAXIh7s
CHMbOACwbSHKIKSsqVEfruywLtVL1ke4hBOdqSKWy4zaRAP5prE8Aw+9klSByvOm
c07Fe3sdedU/Haxq37U3X2hGx9+9/oqOjRMKeZPz8KVBGwZU3eCauEN+F76tEH0x
nrpnqus+iqLegtMOrvpFIXNmC1splfBuHENo/MwvoXyK9QEZPunrJI3vbvUQPBbM
l63esG3jg5PvxLdGUlIV3mhEVAiwodu0smp4K0CEvYOzGsTgQoDVycogmN6gCfKF
5LCYqi36SggVp68GO7ioKon+2g+5tIR58gs1T0dSlgvQmUF25Zn5JScm055lQL+g
CUe4SGSNnAwc66Y9jaikp9e2wRjrUVHQtGUsryAPC0Ax8tsi9aRp7bqNHDGpR2tO
KaPwTnbGIJSC7opxBdpgaZzEG25owc9tBhyeYU5Xiuy6bqxXOmDG9B4ik7MzE8ad
d2nPlDpqn1TDsdMjGk7wqoXO7vIa6l5zvspYXgHJVtIYK0eYlfpiG+/nnwFh0Xi5
0W7cL7sZos+Ht2HEyAkbrfyUsDwppYFIdaRqJg9KI1+irbVXpw2W8Gx1F5dQYYxC
PNqYU20Mcn/22jBlYVZbIIODv+iUMcn4WGl5fvQJBBeWpOXGf3+FJeBYhGbEpk/L
ewtVKhS1vvi1LRqfCH931ek+kM1N39wDxKOh/8BEnI0rR4P6UrPSVqPHV4DO8IKV
vBnsZtxX/LCEb+CTkehRL5mpcNO1PcWgklSujHveWVk2YwfjVs+MHsZueZIlqeoQ
OffyMEBERJhwqTJ3dh4oxUdNMFpBMQ8qY5xjLTmuURYruNvNjnwBKhvNEtP+6E8h
75vEwupxq8i8tBy3lNm6a6cPoFOsAElNrXy/ywAKGy+CPYs91fwOX/dcfs17XeXs
WuIeRzl5q0Vk2eZmfqcenFtpqNMm4ZyomNOEzkEEhiltGWrj1oH971bgMIL2TFRS
xF4GvM/qMe9yZEJnMoFGBWGLODKtkfEwuk0VRmBll5dGwx36ifk11huO51+sbOdy
sYvZ2ea1VCy8MyjGj4YSjhrYLwAFDXP81W34NjL1cMa9BvxReZmPpQ36NGXnXgGA
9URLusdFnrRSxQY5com1HVy5eL9qtQ3tez1RCJ3sVdkoIsZBEyrxNUBWgLzH9yj0
zWDa/kY+GR1v3OyrlmJcm5WPbDl8fg2mTFrm/YtVVVz6L5d/KnZw3+0o7d1cYGF6
qcL637dY8dpLPD8oe+SrZKSe2LkKBa/Np3/JSK5Ramr7OsHCL6O+JWfnTpE+ZJBQ
u91DfUtHzQ6CW7cnjk9femmnFX/e6ZLzKjo+Y5Nb3KjDPWpLialLMNie9tJxlQU7
vFaT5y51/+RiQLI0loY2/YDddXW6V6sTg+cItHE/3QGgpXcxg4z7y8axcuUsbq4T
Q5MHyOVSLDGk//5QUT70YBDCMTlElMBK49j4nt3V33AXA5Dppxpm/3iPDCeIbuAd
H1Jw0NxoPXmE9Ez/rf0cwv/10QGMC/sIm8DVDbmAUXGfT6yaNNd+435Sv5nS6JKN
Frpnw/Y93h0/5m706okiKknjxGiW94gGQ9LZbH3pBpv9hWKv4dGvRejBe6BlWdhe
JSaCY+XIVGxFq238lrehgpkP+S9iLbvU48KshJIq/i1crChQCW5q+39qMle/6pd2
7/je9McBprIcQnXwwJSYQ+NuhhflTb2etAWitSuSbJTCw0jcLxw800hf7n72pPPj
GuRxSD6Pi8Rdf4BFGfOmYJ5pwDT0atB2LoydeRBVtJrOEnW6CCZHQVwbClsWRhNb
j8VuZn0JO+3MsE5f79vISxON0r4/cOUCFM7/ohyehuwplPkRRdZD5F2WywYez2TK
P6wXd133+3xyFFrfb8iDPYz2ZDaZR6bfylAqAMYIhjN6qBiZOR/l6huU46pXYNnP
jonm7fo8gE/E/WPxJOFlHKPcBVi5TUFQf2rYBaFz3vdoXL5MN9FRgyHHSU+n7KYO
PZ+LtiEoxxmqFJK9OlqH80X9zxzhXDEZ4HOgoOw1dfNAAtIXYuaXYdvlzm+oDZ3M
lSn5Grzd/KGI4rY7tmUXCouOED2Ro1MSMwIRnt7Tk2bRD+Ce1ucD0FEp926UkIUS
W+NcZyTvtjUE7bDnawViznQD2quKr/EtKHhP3RIfL6998tRtuxXq/vUBih075UQz
iG+jg3YHknctw77yMKjVNz0UFKIilsvZ6/qzFCpNMfBrqp6wtBSXMtpG6/D+Kolz
Jq2YvvYh2TnFgVY+MzZYRQX8T6cGpG0IXOPlHq3ved/BamV6YzgZr2w4iE+ka/e4
A479RUcvsfNgE6/+LlJXt3uMBC9rGc5DOT4d2REbUnzrHvck1Ah+BMdJI9dwriiE
dJ8hTOCPxE9TTebIjz5a4RBYLtlP5zQJfkIWAF5fb3EBtgDViRocf+8QOdF4e8N1
s0lNJgADv47A0QSdi5oEiIxgw3LIfp3JrqXTJRdBdQec0UnqaMpssU+ovfXVuVp3
/CZqoMtWSAp2BRed7A0W/LlWR8nkbXTXiaCItMnER6fD/HnrXUACnaLB6L5dYAMh
GlwTl95/2T/LL2E2J2JU/m7DIBoa2oV8lIP5q4R9E5RCTwjRoY6RfhtMh5yxrKKG
LeUTGpM3wIgCnkdR5hT3Eb/uDXv4OvQbIbpGDE3OtUG8eZ10UMWt6IOEKL3tFOuf
3MtFtzG1mqWHYXUcK26QQmh4YaJscFMmGk+H8chIpPPTefn1DcA8JSGEfpnNavQX
EkP+TahqnyEQ+1sHi/4WxO6rCzT3DQv7peiCE3m+tA+W4RQgbJ7OXfYy5IPwv98H
zsS8bFAeWcu8+3VDnh0VAiQtmvzjtkHGz6Tvv5Yvo1VH2iKyySMAm+fB5E7MVm/y
lZuSWUWobiHr0aKQ99MC0azM0u/CtIABbiW+xekgmRncSs+7KRoHiW39rmklp5DW
9ZqZxTQIjADQc+vpOmg+k3UUZvYcf2nFmu3moM4FlnXJpObgHrlI3qjSzW79H9GO
dh7LUUt/CaQwjFsiiKCi5WvlNxcial5Qa0BqeiqGmmIrDUNybbKnO8ldZwOdobGk
gfNOSsTxsYaSkxJ29WiO16LLYsmpIS1pB6cj6n3HIqcnLSE17KW7KoHhzzVsrT3Y
TyrCnGVxPUJbDZMPJ7cYHsxXkEeRkyOSCqx0+7ullIor+rICDrDdG079xNX5Sox5
X/DWHYES04lL1zIZjCR6VqQ6yyGAM3Ec6V1s2GxeUHmg+oIEAsb5W73/mmKGh0N8
JCcs1YHZZHt7Vn402cYDYrv4U1LBTpdyRvPl63wSnghN4OtlD8hGKxXXJ+1evdxc
oFOp2o7hJh32eTFYv+CbYOogtWmdM28AJkmnNV+KuljDHEzrlLimmJjsuEr7copy
d+npV3faX5b9Lyhz8F8OsI4SopZwRQ28WqSHoRM/TF8bZUPp/NAjbsQumN7PGgja
1H3PE+EEXgkyFv42/Hk4aUQJ6nmWe5mKkUXLVkcc7w4Q0Gn07lFPQNFcznv+1S1V
OWfQcyCarC0Wt+D+kZR5k9ieppcnyJhBg1vlxKmxJx3yBabPdHS/HI2kFGtDfG6h
LfpLzsSSaG6wQZVsDuxcJAzUmiWRLVitw5VwnzeUs79ycQ25qBD7tRsToYxcmPP6
qP2ER2Ksnwn8uHYJ2x5pR7PWP3HwI7vNxmB4f2SdTRXW7UdToidUvnGMb5lic/Jo
108x6AkB+AlKX59+nr4e4UFkqriVmKrtXnx8gahZpGqBUUJpyLi8ngLLViToV62l
rdJ6CWen8kF47HNrOaaKSy5489aoDWvQlq1gOg65+Ax0HWc16UMClKBqg8y5cnPr
z1llpIPcrIlGm3FEKvIos4voqz2r0/d6aT1fJXyBsWDCWYu6aTaX0QT3rUgge7V4
g8qbP3FpE/N6qniRWPeaJE/2Tg1e4+7DxCvilCOZk7Xx2aQB7p6UAvpDMrP0dWmo
zRhnCzlJGPjj1xa2moRuAide5q1d9aDCUo5Zk1KXodY88SxpIHFGl0xLhhYjIUom
fJP6sQDqGTt8qTDL1FG3cRIjmuQ0yRe6k/kSgp8UjIcnAm8tSiuwNK2udspth2t7
S1BibEAWG0kFa8gJY6HuoKJuMCIevQPF7IxMv0dO/nUf7HUFShxXAalMx+98msEK
XVA71vi4Kf51wrnH0G0bB01sphhCFWIieCyGBYmc6yBmPaPZugADIbH7M1aB68w6
8qTWosm2Um247EUGBYhD4RwFE2z480JkFx+HHLxhfHsfYQ1SO7Oejkjbe+mgb6O0
6fMXHMMCcbKODrhjpG+YxbD+dh+SiKehmbNW2AvKeiHCO/iwMOhoiV/cLjSxoJL+
qBiaAogX0hD6/1vRn9TPSRTOguM0HvLkhEX8xDMXgIe0Y8JDYxA8ETlt9ZgV7x1P
xIN2dZdOypYF9qbNOSpKW/k/Hr0Xd5yVtv+oljhNXDge+/d6XLYkBBh5bLwKAGnL
FE0OH2AC3vyqqhTZiCXOIyWuIfGqbC/aTq2jR16dY7+mpOqZWy/MmosP6I8MkWml
iEGijguEX6E9QHo4FpQOwdpsLNIw2a8az5oIbhYNeuMSDnbfu5gEYWTmQwJrwiCF
U4Pa3jW+VzTZehMfAihczaa4iT3nRBr9MtTeRsXsjGRUCG5bF2v5DXuQSdssOcxI
sZL+UlTGe/JTEMdgCXKEqWP8a75YJXyCPlyBZWnsIFKuKdoXiPBdvDAA/dbNJTov
tMMYHv6gfJDsoki1nfFfY2YUXgbECvcCVwvbhgiTwbqRyIdZe/BDuEr+hbEdZ64R
qHYf+YdvvIAXPSAjUuwmsusaszADpm0K1dcC8Ssw9mx1LtyR75btLECmrgsozp68
ruwhQPTQpN82c5cg7BJwLuq15M7hJKKxevO3bdgFChwhSQ+GCq5aFHszHTr3Xr9U
84aIzNijhlt/PkLthBscdQ/HZ7SVpYbsFhY9u5fkRRsM6BgI0qBT6w4uv0VcMBRe
UEWz9++B2VtvfGevQHsg59/9+sJkaNZts62ThI/Dv/VxIv1bC8zd8SC1y9Xy9xot
kKfJ/DlX2MgljzqwavKA94K0sU/yLEzElgPjyx6sGdgrm0QPOIh+EqDBDg7PYfma
e4O4004VyLCUCHgg9VuX9kfRnlMeKpAl777eGWNi8qpCoalrGk+D0eEu4fejRmIs
sI8D+zDKWrkfOoJGuodXUmJbw2zgLQKSbth90uAMyRQtGyHLZjn2tz3fT43n5n9x
WcctL4ffFh35kTnDVXzQu/+7m8Ssb1X7k/Fk8JuoC+5ZT1SnohwYcjszlO78CrOM
kVBYzq0jFqvJLD1YIMP6XfkcWPf004VweGKnxIND8JzID7t28HTsLFpW3fcEEQVy
qIhrO4qVmePWQDdmGe9POzlnormZNGuGSoINXq6JfWjj7gQVuDV4KmmP8CK10Hzg
/5+2jlee9lzoX/FKIByvfdLpIN8VjsubkUnI11MGm1NU0NZ0AmAhbwSNXsYgfb3p
jX+a5iSA1bggDDtD4/I924i9faXcious7hT3iil1zKJYxkUuslBsycRBmHxhOZCY
zaV1BvmM2oWqovoq0apgxr5/LOC49Zro4xr5E1oeOS6WFEDIACYN0lqtOYA6S968
JAuESdvEfcfah99gRa16aSlrmDjfjrnulj+IIH7QQLAHUCqtRzP2DU84U8CHqtDB
wI65jO+SpeusELLIcpA6WVUGAcca1sDGV1auFeKAVmjUNHp02A07kXqVlx3RoAJh
uehjSwAOkeDaEFMMIwlLi67ZWkJthVRBZJuLBUnFAZ44F666qHEhbIgQmN06vGkQ
bxOAzENS6P+26UMj2Kms+RS0jKiD0NCtLudvWUpuOi2xCJh8dXnOq2+71fJpPayN
cbzL9M5SWlthzBUH5MmMPPjoMU2oAimyMP9UpmeYwpp6StZbjVVAc/cSRSKn+OaE
z3b8CHzNktpJLExiX6gSYV6QiuNbibH1mqJdbmazIFDVT40sxQnJ+GgRxV7cYj0Z
6/NeAq35ycqCxih8ytemyUPUATRjexry+WWesvGi/kgPKuy8MUW43aQ3ldgaGAnR
RGpnRDS1oQzuGjiDlxI4gtZUeU4hqJjXTfagPtvy+6lbEs3XsJ/8S2P1tI7KUfeQ
v4E54RfFEF/CbpzM4f02CeiYJfW9iYivtYNFLw2XOjgKPmkr3IFuvHsbrWaYaW78
RVojMe2qEtR2cBT9CjC4wfoJwkoFMJfr/fm4LkjQ3BXNDyqmAwWyatV9+wj7h77w
X5TCFmMxZFD8Hq0bArnWe4Vu9blrdTQBQIwB4pduaTbzhD0V5t88x4TQ2Q8qf7OD
wTXTFZv/FjAxyxZzYlQkdY6tHrERvAl4AK9GIuFi8LLXDKHui7EY1G9OtNroYGyW
305w/7fzgVnKyN4rH+8VoEb0our5FhtcrK+nejzkIXR9qkQZ+EbfgHA9gRtHR9yo
ceMb/l2yqFc0dpzJcJv/OfConZuVMCFaltXoLjRot7hQhf8s/pZD5sglr7taFnoA
hGgc0Fpq1fgJZGLymIVOOaR7XPrYebNY8DmUQkvIdxNZ5AEq6iVG3HugMqXR392E
mJruNahoMI3DNJQbdMz0T0iG8ekFrWT11j8EMFgitv1W2Ph7Vt+vQwUcPqlwlAgM
tJrETkpQ1hRNeC09S5wPNLzdEXT+l22E/UlORkUKCEWb3mL/Z6aqqGorGnHJlLSr
9MKCTj9TFHXPL+S+DZSQjI3O4ds8LVHr8kv+iZ0xIBayVR70So+w5pRMrNrawKcG
xaHKgnLInTl8cXETdJkYwxCB5oKlGsdWwGwHcxcpxtnGvVg8jpP8qezCPYI/n7AI
Yw4yRqsxOHT+m8XAy6gjldeF2P2wLwqaUiLCl7Z5tPPVf+shcqHekWI0+fxpId3d
ziEndquhc9R2kQ09y0sOdx244EwubM227lQjzPxu9jblWeYWzCzVX7yVJRq86xnE
1PavR/HveoTW0X4QzoVbPbYZDHncBnNwMcZ4hqyBX91wWuM6WYcLIEjepy8RDJTM
Fk4W/QuP8PfSsiIRi+U6JGtDYPQqQbQkzWdrfCe4SnGZ1iyoqQXb+1U9nxYxKCt9
SQYIkV7is8tn6P02HA8U+koaddMYT9bLyI87EnouAN41+4MvhQ6TCsa4nnHbUnro
fjl4gy66xEq1XMSaAR5VhWvO96RuUe/EXUlXKrZduagsqD6RuHrn47P8EuJwCagg
Kehu6ioJcTxTL8bl9afSfyEH//d41vfe5LLbx11n/mFrxolxLe2jIWZnm3ciVmaA
bInRqMi8PrGqxeW+RrpDYOE3MQeuP/oX64+aOXnnXvu2JQCw+c7KQVJsiQmWd5D6
b1G6JorfwavVAhKHL1v0xw/S+qTholet4/v2QjnlKUm5sKxHAOC8Fdotmo3GWQUE
xmEnqoeKviPHTpMfRfh6r1ubCgQPR+9HQig/KF7T4PvnnBnDlT6Pmdg9apIW/42g
48wH2iKvC9rxxQaNOFPj9D8PdB8kHXrSkaUOZOPzcDKf9bHotINk2wLZ7NiLg9jb
JbciCQ+bzSpuHTKOLqdEdMnCbzbk37FuSwQZEN+pvySumcbFAuUJoCdhNFm74tU6
H8GiyKS9cyfKHTRepfHoUhBNQUc/u+nqQZjCgGguq+BbOdJ3sTPXgYOVv4APxenh
txZiU/zABrwxx01cxjw0fAJ71Y7/Dp2DkM5kvAjOll9yYe5pCrEi0zfIJg5yMZjd
NXCqRaMJRo/WtgsPAZpkvmzRDEqdCclUKg8/4MHBGyiykhKuEuWBeW7F0Jt9y+59
Syw+naUvsYYBJqaQGKIaTPDdKO6QWvkRN3k64fj4vaLvPBPnTuDD1qba0di8xE3b
vaS4sya/9gf0lN/FXE1ZXtdV1sJi17p4gC1D47loIL/g3lNnM6nDI+u2GqKUCYNe
YvJk2h1RQ2DDi7fy+OUuPuuS7zeNYpweplrxcttpQYOBnGaTSYi1+MabbxMnXipi
Dh9PiItNKor7hybFApVhLGlf4s/yZoMmVMbRS9Z6URcampOXK6Zgx2ndxE9kEBVd
dJEQalxb8A1Sqj2BI5/gcxxsnId32ndE9Q8iwJxKuNnybIgWyqXOsxTKJjSex+e4
GG1g6l7lrE5xClsbZecqEftrrtqanT8htg22kg3v8ZygcrFqOZd3JIHPbiKOMi3b
MA/0HIK/FT7/L3ZI5Ui+XYOXCcb/seNehLpf1agJtUSxMXpBIYANVujnNEPVA6f6
8ppvMMnFxHTtWGE7Fbr+jBOxOTyF8ICvPHZrhcs4sXClliyGT0UMhILILWcObpq/
RcaqqdbQ8Ej2Vjg/w9jcjKdsnXgA9sjSn2EAVr5iRLHXZbVXve4rEW8cUFXnD6eH
MtOaL6OOszLYxXSHFTws7hlJR3NjtOK4glEC91dwr2BCDcBtZwFxmUlhEqxQxrD2
V5OPgvkcK93ZikqnlZaLygqs9ebkN01C8x6GNLo+wy/yQa2q7V79G8sGvGXfBYRH
fiuoA4lpdA06R10Z0noUDn6dcPYzPtj6qjkDXiSHQAK3P3U9SAZnafMZvxlJT3tT
9kA2aYQoS7gooqsN9med87PkEyR0anYl4jyM7kKWiGwF12/zxQol4dWe7NyY0nS2
UdNr+/Gd38zK2tQSAQ9imR4GmXI5TjI1ShAV1K4cAT7VDQ8eGYPSHkEHm4lJp0/S
bjvjezuz5yO3EmfFFCziYH5A81udBHrAR8or8CZ7Zs4USUCRswzbGoS4JcBPAzAl
Lt96b9etfJcEfF9XnUXDrW9DmzDrb8sb7Iy64MLWTeE9uFJMsU/LEyZXDe8yH6r6
t2GeJ4vseg+0NRuBwHTEDvBp9u0Ttody6n6pnXjC1c7v/G0ZC4+591VT6idzM8vr
vm0sdtMTDRchCNcNv8+P+5MQTKmQEuw6gwVmq2EPwjKnvH8IIcUq4YXlRzhTkKqm
blroxGkN9wC2A7XIunM2D6FJgzxK/TXXN/rKifi/PlZlurgQtZp9/aYrN0KfHqj5
zgV2rJ3kn/KZyewBAkuHJklai2goL+Jp1M7ERKtPg7+m0zQT/d+m7r+BWW12Khve
J3kN7Xho8cfCtiM6IrcP/GHf80XBozI6LdJw4lo9rAuCD95w21xxMdJtp3WEX5Ja
Kaklc1khZmclFg/NccaZMwMUQul78/Xz/IUxQAF5eqkCiRtNG76v8OtRldK2/rgp
QwK80X0XnxsS3PrAgFtRPrE1sxvgWSKkqpTPm3Vwqt/tW2LFbps/qG/5RlZYfgkw
tBw4zlm+PSEowLfnVEtwp+YeOZU6sk/GHY/+UL7HRcfKtQKzsEhBvT/X4sKGBDgp
OnJySnWRJr445WwDbLxcaTKV6dqdDRwWGAeD9anl+BVurAKv6Qao1tObiEEbfHqw
A8SBEISe5V8FGJ614R0Jlf4mEiKl7e1wsSqf5R3WCWE8c0/EEoQz4LNFfppG0gcl
2e3I8274ZUC5LufchdXeQI6iuWQULhSxvXYUDvi/di9XpDwJGZRzHW76iy+iggkj
Yv/TOn9YbILvaBV8KILDYtmkEphm3zv+TVtnLlrochQSw/EkAJJCnj6lGWpNEp3J
i0aDRgmqGVmQED4P7fQQYNQxRCGJk9igW0r5lMCupQ5APNcbR0Uh1N5ZHouUXr9o
XEWbRvLWWzr3lBgfqHhswMpE7eBllbh658xuc9aXnl9QQ9lqcqHBTxiPSGbPeDI/
ravlRE3yHoKYLaDu++3qRZ8W3fNhsKk96BXMBE6rklwP4DX3k8lFsFwWeVJpeh2G
0Pnm2DozvqjKaHXY747NSeel//zTQcgh8yibk0ccVMB1nNWmU9KtRCRdE+dzRV6H
WRm9OPY2RtbnPs6CwssCQwFAsGXK9odFxxDo3LnALDMXS3H3CBvA++ckVkWizsvr
olAxb6TGDQ5LdZPUBbOtCb0ksAv5JfwY5N8WajYvYlA/hZC0v0VJSj705fLmB8Tn
n/BW7b09D34iw1NrkI5dL/meGSo4kREpUI6DPzc7JWwkYUotB7JxyBmvzXHaQk9w
0eCVHIBVFjaMAF+R24PssX8ceX6RN6H+ge/tbwQv707/IUUgpPzNsSRUe/0itgb6
kG2k+G0EZ6D46d3jALAiTemOpqXNaCKwKcyyerThDPVykRA0YV3bUN/FpWC+l+c/
VkiQpEFgwvYPABUMsT7FOR4HKCjfpZWJVuQHUu6X9MebeCcii0KI1NELDyoBY1ux
5chN7KS9H7RnehriVhm3m1DbnhL97B9MkGdLK8yt1mqPP1DjKHbBxc8Jf0QC5nBz
81kh6hYrD6VulU0Q+uE3xJ2TMUX6KWJoGtnvMo1MSPmRIPx5/UhikVrCX+HfGQ5j
GyhjDgPrgWWkOphN1kYSqBYZ28ID7qLp/xnA1PSbgTi09l+hoF4wczMQ9bOpgOHW
RgQsI9SBvJLdKTwzEI8vPOdKEqXt1kme6SYjpwH4l9m3hIUYlj2Vv5uWTng4H+1j
9XwlEVBK2Czls4xMJthWs0VhSI3GbifemfS02R83i8LRftrmKkYsTvv36hs0DfPa
xgYPdu2ih/vYtOFCmAmHRMuDKGfC+5hxY86B6oNmYwAcwUU68NSk4X8wnHmsBg7W
Pj4nrqeAT9QpHor1elx7B2gz7gmPqQA3JorSpLFJDuKczIM9T3JvN5dLpwCUZDmS
vvi6h7U8/hvhSj4dU6XYaHpy/HgmKvitUkj1fO4xpSeAPTrJ5Y7YbNOfHfB717XC
ag2q2i6tg/pVQhaEWeRhZcEs/ZehzVVvHQeFplSZSRnMo9e+bOmRualfR0PVBO/T
TjyBxTkXdkZTeJwKbfijbEl5++bIIYkOMgAJ+YePBD7h6GLRUoeyPOGINjNu38vW
J2DVGAScU5DbY+7zGpmh+vFFHfYhpDYa7rORU5bV/dmyG9gS4OCbiB7mxBOnhZTd
ERK6qLS8VukSmBrsIXZkSdA9kbbjSbihDUNSzV3+nuUQaqpGzelPebMWCsrdTcQP
bhqO8MJLZafq4LcOsGDbZ5D1nfW46Y8bLlDpH42LyDVEk38lmIQVEdeLmq4Qealo
IdWWf576Cq8tlgELOmqSlkCc2TUzGrOo3ON4rfhaOOlLGvfW1CrJap+0wpag0MbR
zT/bFOZyjG0mzhENI0zr6T5l9AI04MDUrFYvb1cXoESAB67iBfwkPxpa2be2oWPq
049+io7NdX20ytHf8llO8o7E45oxiMVHu6VK/W7ZeJiW60eWbBVYNps7o1fk5jj3
IPOEvOLeL5lTBAxxRxBjLmo8ty4stLo2emZ+APpxKAQ5+wEFyM7orpW8hhlDG0AF
dZLoQp2XLt7tfvx5iZVeSMSENVnxaur7ShAywSAEOHRJlZkLOCo1qMez+AmCi7Nq
/QNEYPRg1XWb6BynbcRXg6wsOBDB8KxpouPa255hE9tcyrAfVTeB4eY8skycfueB
wwomFWwaWnSL5vwURRaZi1irgkrcSna4vcw6GCsetoZYCLS9IXoN7gWWo6cevoUS
tk3pTw4msaB6uUKuU3Gi8HqPpr24RQFzsekiPoW+N5Vz6YL9yG2i7PT6WX6qLRHB
pBunkxOSIYGclXRXeFP49WqULmz6IhTUDsp5CT5x+WbTtvmQ+Rhdc6oD0mtCgoz7
IlnWStQIG16SZr7GbXwQy2kn5rMO5XMF3DGATR3XQv7VsWCDd7nHVHwxEXftB0Lt
Zs38bvOTGgkOF7ysrrNrl5LVByvECafmGjaq3N/QJFIB9UFfi3b149FnK5QXG+0C
xWShLmFwplRa3ythRgkABPYEd7X2sOeEylCcNHW9wnhfKHrkXeWBaat7/0VkAdzJ
2fYilIsfaDcvn1WWKhatAM6XV5YaLYbFpMlAKY6hDHCfOF0TchOOOaItZbuOPmGk
ii4ih3TSLlrwzvvTmYViNKnd2pSEeJEJucjXxSaBUfYtild+NrO3opL1UE2xdGYO
QkoOJACIQwnffoY2fjJ+lu3sn4GNMJDuyh2VeiXWm0qV1BsWZDr1uwQJ3JJ0zLqy
/pQKVVgx8uiyqe3urnBJW3ZiUEITZjxCildlDu9XhAaqv2Gvg5DLOOrLd6lcHo4s
leJOhx1WwD5SzLA/liB4YA6iCAiPthdPKCPuiHXLU46jWj+IZ/huLdBGoqQbyHSm
IzFN31aMOWkaLiY1DTKAz9+Iin8zN7pkz3H+EWh1wKENc/rz8ABTBbRljQUDdgeY
0HQPt0p521mTHzBSGS32040fXDK3l3lZlR3E7evddEc96uctzcnLmS0W77snFUD1
Sz0MMuKiOE9t+dgKYzQ3bHBVl228QzTcB8Ae+Abh9y0Ozw/TBqc6i7rC7Y/Ym34P
9YMLwFudi97z7Lc1kuAQJnDafZZ+6S32D9Tz7LfFAUL6SO2YjU/dmssN0ISzcpdS
wRYlRBpVaHFwpO6tvKk56ABrXi+G+1haH16XJXBCfOEMLXY7M7lx+JfBrmTwr5F+
AOnBnqE8NjtZGi+0fGVMEGP9v8oFLiTBLwyJViquh14SDJsTalNAVtJOG7r9P+KU
S8BhfCr2RtnV67rCHHlTj8BwW6ddK7LEIvF9xpEQ3lnqyfRn7WgFThk4hlUSa4Tz
9Yv/kt+csvcw9kXDmYk8Q+U84wgkhyZlRM9ARIYeQmuosj8oC7HDT60hC0XYVFVI
m5eqxbNyyH+sB+BjLbIYMFGJe1faIHjKQqaKmsB76zNIRCxY0/RDfB+fmWrg8TfZ
YuoKgppZ/LjPxBBU8iczqluGKmhaZkzhKNhyZ9CywVtQqFme4eNVvd1TVc1gWPN9
dOc4x+b1fiXa97maYQeezNRxDaTjZMWFf34nSgq397m9079igy7iK7M38FU9wGpy
FreieXeN50jfjnbzVfp1szZd2Mpr3YwmTfrblY4iG4vwCZsEClWyZUFfhMQu7438
Jl1Q282L3Df8xT5p0HPmQGm5vIx/6VxZZXvHR5Ttas/hV63WnKtSHbXe6babWwRg
MKfz1ELaX2KvoMYxAenk0Fd0I5rhlBxvzz20S8ao03VuMPyeKqQGJa48Ig/F2Ly9
KjUfDqfWsKp6lOJVdX6wclLGHi8+mtVkYbZlFyC5hIVtwn7OS3AToRoEvJDtKGCV
h5+w5ceSqt9fgfM2oD+BLRbYhJfBNLogspS+UOF5PABu7R3FPeLYZu/fVLOqjQ27
lQQpaoZ5qvJgXny/e71ozBmFksT5nVkj+yggWBqNZ14nPqeUeni5pDHEfTU2FDey
/VJJrBfPcnhhozFJT48NhMorpjBmOnnj7E72DytvF0d808qE/qihRNALN7HB31Xt
aBcwucbrIpyinmPzhzapDs6sO4nPczdKQcvq1zNfgg9Gw27xDcVLo/XP81n9LyCw
yEITzcs73PisNh6lVplaeXup6wiKFZW57DwaajvTHC3xcy3bdiIQwLJQF0KFk4y3
Ju9NfEX7Og12vSfu6JpTWj2plVVbCU+uK/cB6I6xZq6Vnt/IqIltMl4kZ1hp7ATN
CYhG0TkcelrFt4bbgYDY8U11W92hQ4wnRyH54zHG3y3M6X2Q742cyDRF24gv/aOT
qzKdEaDziKOb7s7SJz05ZTOXtH3r82+DgLWw/DHV0yVZup0ogadaVg3+lTwp7Six
hWtW7GDLLDmXZ76E8gXnj2FdLHGRB5A4sU9ZMHTj2poQtOppQzjmSu8XxyKQlLps
WbBlNBdvZIV2j3N5+3gJPGdhPYPJL0erO9elFfcUjEPv3uGjX4oNljEPkecduTbm
zQvvJqFsiPLmOVIwEeKrSLa7wREf4/NpUxkhk5Q467DH4CPKIJTIBPgf/hcLlJ8d
fNFthbrV1jkOYmi28cp+WP9nBgoj2CJR0LAB1fiSP/o4q6a1bu/5yCka00bak7j7
lWbRPDkSwmM2XE4mGgVd0/vIL/r/nYf2p3+U54P2dVm1KuyllyV6dLrDHXcz+XoU
Bp++fFe5FcCOuWI6eiTJyQgOl9ZNxdg1KkaTycqy3kVa2xoerS33FhvR4h/mDJeQ
nJWgUJdoc5LCiAfA9wCLcD7tBx9vh/LrM91OWKTfiGcXWI5CVn0InKFWV8Hebim4
gQ9fF7p3UU72b60ppTrYdVyWK0YplDSMW0nuo53AA73KZhdAkOvWQAaKIUdxGJK7
W3a+MctXLpHlLcI5YHyL2cWtFa3vY6dI/AnW3+hYil4Ay4yXWxeZ5hwSnTqKQrW8
FzG3m2B3zy3rNLvD8mLzw+Izn1k4Zs4vxgys3uL1khqJzQpIMMzi+WcbuxZY8kN1
hcaGtCK+c9NaLvNHP1DxEG/+Xaf6km/4iHCmfmIE3zk+Cb9Q0BcysfxEClkmS46m
pO4Zj/a/Wb8WS+Y9ss42V25SOokQyK++0fMHjf1RnMIFt+A3fCH2HWsplMEO1kI2
Gjwf4irqeIBhd3tNU1xTAgfixrTsSa8A/knMsHbZRGruUMckd6IsAZ7brs+plpRZ
R2JCv2mvtrQEKw55ukw5aLfjShP3WzzzLZW4nCxAVOgiLhju6NCJWV8/v10Z6GR3
Gay4mqKZQxzFj4+wNtkWx4SEWUqAS1EFr0OG2HKYXoUE+yxWLpbZq4IYyBXENURd
UIU4PLF5NoBgF4fak+VKsqGa8BPOPIm+c9XWwTi63ESo728xAN3gP0voBQ8aqO+x
SzwiDIs+ampXngh3LrFbtcfShvpkuahb69JbjH/Tw7NoaDYlSRcGWzSJSjL+NUtq
wjMEacguMAyHxlE0bguwdJllUErl0ffNO37Zrp54hc9RQwuG4LLS730F1r9RoIbJ
47cXCzB0bxND7byBHgTVuopjmc+NZyot7j3yG9doL2rah2utcQkBgL5BCUEHDS/M
xNfW8YfIoQHB9IEbaH6fhHMgP56+V0a+m1/GV8lAtiYKMgdGobyPL2sClPXqysfO
U1egCuvjZqtqkE8ScR/+JHNUDmVj4Nd/a1IaEv4nmWwtv6molvECl5wmUVQYsbnE
uTUkNmN4u3flICl5QlelwM1ODvIcUQNGj6Eb7x1itWIbP49yrj8+PSQ3izCARsUY
gLwEOG9e8kXXMOWvMHcgt+e6IA2Wdaz6MzB2e7kCDI9OQ1J7FGoEVT0j0fCyTilE
W4os5WfYmzGgFEJMjwxFAuUMATA2xvRRSMW806cXrdKN3nED1RA1o72BoLRRjJF7
Y5tFw0LW1oNn+A4tfCDE7knGH2baPpAQ2UxJasfLIoGO52AVVkRcRYB61NPfO0n2
WhWyQ0jEi+1vpC0jV3O1oyrHJaoOc9+02/46xsunvajvVW2BJdhkMfCfqoWYdl0D
s3HXtjWMqe+gMRH+cvP9pzx+PYj6aCOLuYJTYZl5TVVHDCDcdOjQ00rOec0QOEUB
oxgimW4hwmvNMQMJGnaP6C4AjMOmGuZwdQ/wWM6gQaG9Xqy4waMy788hR7DVDQBA
dUNpq3Hl0UkjTpL14M8DvZGUxT/UtpbQIHLN3DKAjBM4Hp2L1gZiWt8GUGei8V7A
D4fXdfwmaq3TgIViyVUa+5oqL4UzNctZuEHBUMQhGkqICQmdlHszza2AekPA/dP3
W8wz6d3N1cyY3E/8M/N2tNgLUcOoqDwSa+nawvcIBOXmv4NydnbK9fOEyetTD7/L
Nebn0TuSbPR6ZSCDjyZ3CN0P5VxRFk/m3eLk9uz9qwRoE30ZN+Aar+pHUo9S2Jy5
dDwpDv4biriyDkAcK2jylWrOOcDHnVJ9hh0kskx8H04WSCKfHA6e+/oDD+KdHe/p
WIyhw1qgnANF6tF/MZ6JX80YGFVA4escOfTsujtRJMQEJzS+uhH4xUkubC03KlIt
Pfr8uTvWQ7MTQmRntBQrJJHyyRSntiVF/qLgYmAIZaaCo6Kz0C4B5sVbWL+T6SM0
rBFYqIpTIiCSrsglYcga/vPrkYT0Orj54CiQho9jGtu8eELmuR0HCYb9Nj/kQGx2
nzYmxBmvQeAbEm4IYY+PsnVzuSbPVBRFWRGrFQLCwre6fXBTuOKuteLUDrz3SxW/
4PRZ2eO/LYSMxOcmL9eNvptmAqtD4Lsibqw9tk4oA30c9vnQrasp4ganRWAW4pKF
T+94adD842AC1tXTRlGBJ4cTKM83gFsW2V5ZSd75X+5Kc3WIwIroJhzlYFG3jvbs
SGmgVYCmoYE+TDLdLQ4O7+2h9swjwGCRqswDHkfNEho6s7mskOfJZa0Eb0w2WEVD
prlT4hGBgz6OS3ckvSb8+7GjiFyj7oP6SqYa90eJXqGRxrX47Ua4GT1OJJs0Fcsh
CeYV+kN5lVYWDfiIkHxUcXqg4cIJ9GZc5Lu+de7cN1zqErrEoQL+52sRaXcjEaM3
In17kZJ6j7GAvxf91JWjlQrcijII0+Xa48oej+FHs48s0li0im0qVUUgQvPgkqzZ
2KS8hxrl4KLDplNCHc9D8+i4Way3wE3+MHIq/GFSsOJrEMCX7q6bcMru6NztflFm
bRe/k06TIfc9uONlLaRt+E1nl00QU036CUjfT8BpMPtMwtJhVgr0nHRjqodOttlT
mA0wWRxvtRPhlPKLxkhnan7q425ejfHOooJfLVePokq3UN9sgYxLKwHsv0KV38Ql
J/l8MnDQulB5VE+WvrRYQJwso4xLbgQ+mQmxCC9Izk8lTrRqhBFblbMfNDgXEtmY
TW/KxC66M9tlC6+srcKB6tjBgKk2nVmTkcndt31tTDtQx5jJPDx25IsIEHxEUgKK
ejYpOwc1lNZGRjGAJ4EbZHsSZrWGGr08VfwwTKXP7+GjsG4mWQaMdW/B8OzWn8tO
VHsiOmEsDBHJDP4ki0kADVcO5VS7smE/YTme8p+mocpxAgtW6R7IWufAkh7JDsks
NiBi3YAITybMmghgwhhjy1hfcTglxLWN91s9Z4INaL0LPKalAC8Ez8U+nzQgV0cj
G4Z4zX8pjHd+qVRQGFroGzOpjFKbXrww4Go1Mc5ORnQrP/nqKkKWjsWgUtdWcNus
qun919bV0HUHQsk3RPr/6RmGAzaL4VcAfVaqARPf7AtXfFNzQw7sqp2eyzRpCWIy
89mwwtIybACt7/F8ox059jseXimESiJaptF7VJEuPz0Ffh5fN/cq14D4NwiOeReM
2DRrdXrhNY+KT3tjDbVOLICI+0bXLFvzgs8hzTbswgXrvpfcEGXgPyV1qPQ59aO9
qUR3gUTxDqDQT1rC8Z3Xde+aOV8m5HBjQMJ/s/nm1dL5UpTUKMT6B6ogBXAimfdp
jOiA4CsCtvI4/e+ljHlu+7wz9Dmq74PcwqoVwMfNfmO6ADwoCbUWTNNbrX0utmGB
MV+78aN682jtlrIRz80kUXRPlwxWqJF4XCBBOPSVRGdEqhRwZBf1dzJW/9qyZ/X9
WzBnQ/ty9Zeh8VpIzKclfJRTTC+XGRQny7s2AKpWFTtByr56SBlZEsruPCALtmXy
tc8cJ6/YJPxoITfMcm4FnDwTAlYGHMkxN19JYtRaRYENOn9UK1DpfxC7oRWG4sgA
0YBMuR0ONR1qA6dXfi06MNou76dUuW9z/YLRNEu872ChazKLSqSDzE1Z0Vagv+0R
i4lJamo7lVAJI1d7HOFGgOO9UUgjI0f4/uwzVHdYDM8HIRVeRYsjEhxMo/YT9X5g
DLFZ0pU6m0/JBmAHBTBxV+tbzh2nc5N3MEsRrclIkzCY+uDZOEpIbuKIH2MohPnI
prlAgpZL8M4z/V8L3Wv0l60ziZYTpzPqS/G/CTnMX2c5a1Lix7s6xEs/5y7ls09q
FxcSEo9tkIEElazMUQItp0hh0goxInl1Z0JXdkwhEx6bQZRTszCL8w/Ma6GYa5NP
rsun0Om17VibB04WXrK5d+JRZNiuXOFG6Zj5lHqaPH7IkumPE+ZeTK5TKfMedw/t
XiODHq6o9kcpRkRrWOTxP9sQB8EOtMUOcxW6n/+IFTQBWRJTv5xWJOaBEF50CeW1
RwJxTX0YovehbrNnv6i2rvmSMmKAnJzMPf21SVWnqzdkD46bxzslkJrlGwiP5SqF
wQY7RTA6EubyHRdUQpoXTm2RIu8t8RePPH9+YnKI5oOph0LMwnTla4GaxZ4odu5g
un9zVcrZSBqADb7Yb9mes2/FSuMbdE1d2wWXUCK1mWzLveBKsl0vgmA3mnYz0WaP
kJv0KtMjrpR3DDkK3eYpub4Edq5hN2w/S8yHUHTG6ZTd984DdaAlHy+D9SwUdjVx
FOK7XU9WBbkqnh1vMo63PozV53slPsTn2So1H7UaBWHwwc5uZ2AnGv8OaXHAbEmp
pRm0wRjMy4QbKv9NDkz54FE2BRGJRDhb5E11t/c4Mhcls6nqMi8B7T6wZTvHPpbt
dBTMRnceQGoCh6e6Agd73U4llfDXj7E0kFdjKEueZrrjVoftSSRz/QUBnUXBOxuq
nNx8g6l8gIGxfC9RHgDlhtG3+o4MYKZgRnr34gKUIs4RK30FTNMGv2ZDiacxlHf9
6yWH4bVcsc9L8bLvkdCp+F7VzLB5iSUfPC1XQSzHi51jov7rd8lHQJzi2xXo9cAh
hnG1757rA3ITA61merj+hukpg0eG1hLw5FHwTRuqLmcdt2K2tTR9TI4WBTSPQsIA
mk72sdUrFghVrJkMQvYd58UTU6TbfAvcCWbovO2D98uqdC4f3YCcInhfbt0wlyDY
q/qJXHCo4X2AfMN68dedbnQWKV+iOLh2XN5mWFvlXLX3+1D55mW+va4ssS5o6aab
T4FVPb/KJHNVFRBREMoVu/Bev0pYuqnru4A/iy7RFJ9te2FhciBllW9Vq6SjIrCq
WAsjyl/ymu3iIKR3BzRNM+a3QDrYQJ9dTOzgXRa+a78k0dyxJOeGRH37qDv6l9Il
VCaSlhXeuhQKPDKvivsHpLAfscg6InEB7q2+qk5NRukWusYDNOGiBUvuYx8p/0tF
Y4CJQjPnU0ulEtx1nBjlfNQBBmjfMI27zZPM/YpLkuBYWR/aBGjwk6HwbhbC+H/9
bXguOShu6UEoU7Mou7n9F54RECVs2loGvxt9+PkUALrToEsrHLui/PgVrB3lrCMu
KFVydsDNz3EEAQ41z3sCJvDcM/FIZtNecK+uzMys0MRYcNv23qA3jQaKqo6LdnGO
rTdttYBzf5WayKRGaI7wQBdTCcwtD9wYiy90xTJ0psbpC5mnxMJdNW03011sBwQz
qqiRyIlLJWYWQ5zzJd0k7v4hekpSK5Z/mwiTLN9XBaJJm/lbXHF2JNwTYghUu1VQ
hcGAcQ69YtE91oujd9o0Q48bSqO8s99J27DRwJ2X+sxkobKRHaCzAMz3snWxaIzt
lfmDc8O0I/MU6m0z9ekdqboty7r5ebD9r6LblOJ3yoGl1izpeaOdDDLshbwef+Ss
AemThGe4u2wkJ1RNcpu/W7NVRu1KVOIWUIVKZwSE8CyFMPb4SisG3N2jH1ytzrja
DTCKY0ZIE8SaNtMKftyufkhlK6TiUYO8ks2Rv1EOd18rVb0pjx5S27hjDzGz1uft
Zto65n9cbRR0i7OArsGbwTt0e7a0Ostu+hF75sqixFSThCX2w4F58GmbexSbnee5
stFNWoVFiUqt6gb993xD5GXhgtdPu2aWpFpI6/OOmqoDWVHzcyW0twYNvoLWo/D+
Szea/2eIbVrvT1LSYGh3QvjMfZWOkyYR6Om5wQqAETWoPo692najt4m0CSW8whE8
Gud7/VucuopzuhV+cScGWHUEi9liVRblR5K1YX3rRsuQv+XQYTtVUF3N4X31jlR7
vn2Ody1r1T3UiGyJLhPoZZ06EQ0TldT/gbJ34L/bocxKKSTOEf11suar/hKcv9TE
fxBuULFDUCk4h+d6X6fl6Q+ZN49HqtqAuQjdf7G4HIpvRf3M/hwWoCtxU/I8imwm
Y5/BYWEGjFZthaI2LxA0a9sT3xsUSapgkB8JsiEQtzxa+iFI+csg2uhMC9eAvD1e
BcjESDZHB00JHQZnG5Beklvggx5ccD7L9kXQ7agpTRPue1CEDWjFkVguyHLw6wME
3yzYdU/FUTJEJcOVRtpJPptkkW1OS3S9twRAVzPaFNbotrZg7zdtugcwbFkhiV4F
u1FSm9zMKkDpgDOdcyCbl11a9e8xezSD68e8OigZEPKpk5BzQhodlfKQstleeHfF
SwJyA3U3Aqand/tzdUBvpTeHY+PBvt2Yq/X+VcJi7BGSeWpp7soX7aF4McOxsEic
BqKzS50Qvv5HJj311qqF54I1EsdiGne2tBHAeFFedeZhK5rN2fpASRReiuvewKfX
PtOGMoEHOaxUUtgIKNoVLDso5uxoVI9J7jLrj3l7B/TdN8Ka4+Y5qWR09ahPvDNr
diTuFM2FBLWLFA3G3hJNki2wKrYBu9CE56+yUNhcQ2PIxJ1Jlo0OFJ+QIFqq6nbI
V0b5pZu/XS5KRnEuVIti7dj+yRxvG0D+IHjULlKTl9OWYhsHheq6g8TYcpgGOiid
sTfMCvNx0Kx9YfjBLMFEnvsXZWf1mEx2NHN9vzvA+I5YWhBXSIiIz6mS1bVkVrd7
t3wP6IiLB2xXwIFdVF+W8Z/o9GSkopUNzQeto4AotEeD/UcEk8TVNsUXdkOxYsWb
of+HrLeXCyP6MmR7pETBMIIkdo/qE6m37RNGdTqfretTzQdW0fvukfqi3A94np+E
Ge45j5l7ptJIQrr3VE5zvv0YLoK4IFIQOzxxcJUdvt+czMfDGsU2u0C3G2ucWQKw
hZDJZZPbRBWznvwkUy36yEExdb1I2keAgbECREQJ3o2x4qUdWVxVpb99V1MFFX0D
ej+A0nA44tuj9yviFZe8+EkrUiJmrFD3mVq4sJ0/CSfphaIr39vYFz6B89LbmINw
PSKKrjhiItLGPetD+3WBh3rQTY8UT9IHyinRL8b4nntpnIDuZbtXRw2ejXhMYOiW
E5fjYMn6FqZkwm+PhW56eapVeTdJFAnKDtAFhhuPdEZbOMKSPBck6gdNO8C2ICe9
4YODwuedSWkZBRD2//uy32umEoxAqV4lH9lfJD0EBoQTnBInmnUqnAnQ1rNKZf9B
UCjyQyzPLOpfHhumTNp4oiyfl3er7OYEqwWhcOKk7yZLN/RJuIDt18nuE8VDf6p0
TlzegqJyRq4VxUrwTGkplz2oPMyPMfBgXmIlx7inavPuDJ16MyO3chNDrOBmHIeS
CmmVaES8uL7BJfC2OZz89pXhAN6wBFSgiHZ8zWCSEzEVl/Lytw5Fx07r5W7y+lhL
2MsQgQ3nNb10blnwdBj15J9OLEISTxssaTc+g6Sq8m0u8LaqnUAFmogbPJ1DhYi/
nJ4kntlEHGwlaTVTitjr4VAF1lzuNx3dPt5mG5rM13Jp3I/rBjYJXuIHYVnS9G0k
rAbxJ+cNWwPkRO0E8qJVtYUPOVYht2G9wtKn1EmTr0eiBr4L0LfteqQMdZt+i/9K
rjqSZIg0l4kvsIbPIBqgp6WAjCzJ1WMVjyotqCMh8pYgf7hgXZ90FerwvOhatMhw
q6k6zoxSI0sS2fDEEHep4jtIYvBJfIbKhd7VgcxrwmZQF9mE018Jw75Ou0NFio1c
NI+eUv2pgl7/pn71d0IWnFL/ZV9R2yQxQ3FhWGho9Y9UzAT9fzxlL9JoTarS4qBu
782QKdrMOy3NJsNpwC1hM/kQKxi4ERA91Rtg431sK/1cKPT+RFnUvbJDTqR0QlJ5
yw6An8r9Sk+DvPmLgJOpud0Ezt6yh7+SRrOKT1BOVXMVAzkSFk4RqYpZ4NuAHEVr
hmHNbSC+Rr7S6uKK330Bmd08Hjt41PfY+/IP8w84R7MWVkBddlvifFH9Sq9NMyJ+
8U7wiwWlTJjcQjUIUc+zbLFf8prmg2CrnSPBLH7VLgT7IZXQetcOFIow2/BLEUck
2tUp28WljnzXvmr4rjE9MhC1th6tEgA5zV51RCRx+LQ7Iy+U0ZRLfaRKetlyfDFI
66h2VDm7VO41B3eQZySLF16pAy9y0+3eCs1wbn43dtib51AqL40dc+hsVOmR7/j7
Rf8G/3mb7nNL0qhhG6LPyQe1CRSqJhurvHKisAJ3qU6RnhODWpBUrYBdnAOcJq34
0tQnSpeKaTmZb8ok6TXCiuhhVagEH8gzoxJqPAXuoH/O8K7dH9o33wM1H+cejL0x
AGYPpqmzKSmKZpSG4lK8W2Wx3bQKDmN1ISftw2FB9U6NfL6MSLlFKYrUx4o5JHRs
Iq8hjlrDZykIUacAIGsVK/iejhbdFx6yUiXHgF1rdZ3SU7q9e1X5E2GbHfPGx7FT
/GJkhZCRFrnWMBDujPNrSgO1MXpxHm50T3ghMfIxfWrdjdxkBJsHpWw/gmqn/ctz
pt+120VV8FDvwR1XLApXWYgQhTqRjzNaGXi6266DNp5V9lmq4q4JhuytXYFD5FfL
663/Lp11XssntXYzJuEMI/fEUQAXPzJ6mrCNz+tAFnOMf390oBP9+w6Yg38tZkxq
4Hb/4SEqApgku6ktNguaBNeFtPpnk0ZXXStZgS5Ta9biXIQc7fD5h3mPLhhfYSYs
HmVHTv9YfP38igex9kEJYh7kUaIVZNCX3zccmOsVOKE24FYAWBrV4JJz9b2RL6cN
z0pTYzbJkkji1/I6kH6Gqwv6UPVK1tsHHjXze4tYO9CQtMxuLKnT8iNxztms0nt8
qMh4oUeeIXvt6CDG29sMIZGbQEamTPbLs7M+8Db8S1SpzkKu/yOMSUjthRAQk1/c
Kv77DWw73PzfNVa5yeNgvqU7OTrSssTvhO9334LHEl9H8Rb5gKvXc/DuD2MYrFCV
vuIxsK8ePrlXnPfPts1ZbGFuVkfFqPg/Fw8o8alyl1o9OzuXlQBNTBtSV1T1HhRn
oQnUqLFCMwTkwgFkQy55KxDdZjTGf5DeV/qsYBTadKMQKUhzj3hf6j/kqhuGOpZI
GWlmZUUBCUmX2MSWywHKyDTPx7Dh4WD028I+kjWrJDv6IUPnErATYlBDgsGqpxPr
D4HXgGkGsU1Lu/EEGQ+m1dXWH1UvLoyYLdAPuH4zKA2MGMUUVvm24gc6l9/UsBE1
3Qg9cJG3Ab1xzHJu+VMUU85kQlRpaWz1BVXxYGONIEvBHNKHD1+c1VAZLR5sQrZ5
VqZza3FbJ7a9hSMAoMU8pGpScK8RWoOT1dM52dFIRjB0IsN52l1VFL616gRgpXzN
3dT6fnsAHp4Nn1s847xMeHE6FF3JiYRWj3AvEL/y63gwWjDbfETIV8g75At1oV/Y
iHDdI3jhNI0wj3ebhtw17HaQLndc137RZlRT9kj2b68d+cNywaDmkNNM/gmmXK/e
iA+3SNrCDWbr6oFtjoPuIQfHoZZE5O1LFUthCtCraXHYTCj5H9d10c2uPPi06vZd
bSl0Kwh6kxecSsnwJfwEXR2BNrmXEHYioa2+xjaMgI6xMmF8CzZ1sAOngbhfI2Ak
VQ16fufO1n1AF1SDknUuMwwoKuSX4XTXFyWfTN//i1Y4tjYrJOZBtM98GcUmFavG
aQU5VuyD2jkEuVFEyPMqVr4onCtufC6+NKpYgGbYuQH4Yfa/gdXMcaTT8fcdJ9aV
VeIZUVs+IzTUav02DD26F4moGPRz1HbOEG/9KLAQ8kY1qs0J3WqNDPum4UBv/C+j
BihvwvknLGWuWsNpJJItGBLiNINfD44tYHxP3h85Av/ksbhbj0dJ5qlQIc/3K65P
d2AmCPGJm2gWxvNXOdQ/SYKwkNiRkPhs9XpLnv22qtQDw71xy1C4EWBMX0AnUdMK
uVGqkFnY8R3gcItMenSGRYD3kOTIs8z7pUMc2a4bOxU6N/octH7rR4s+TM33ryUK
u9qTj83I64SlB4G64mHGkLKhrfbJ/QxtOMFOlJmYASYUgO3Mq3N8Foc57UU1Znep
S9e+wTp+zdctPlTy24eMVDLbOCOETo31/nByXyDAl94AbkZvBA/2j+ZlsOdCD3JT
jHg+0v4ohepWGBRLzGtMuXWXS7H2RhUCVNahWlmPmTzBQwuVOuh1EyenWtxO2zfs
a40Nrcf/i/Erukxe/QpiFYIaVEUDkorbU2Ziqb27UTG9WyJPWlLN3Mm/ZuBN9VZ8
1EGEKYKaAtLls6FICNdh/mZddAbtG1/ZAEKP+RQfqzYgO+2m25fdQCMTiQbqy9UG
CzbPh/CEzii3dyg58RO6b6YZN6wrTDupNSc7RsXoyTzoLdQNs9afCCqGmusKH203
3LhGBJYttKKOw4sUjo2sXrq6O35VuYtWUP3e74T8paYV2X/Uuvef79wHwlB4nunM
9aZDw7dMLhtl/u11qI/gUCAKbYQKT9zRvGWS+IWIImq2jg9aJnbTtMUD2WB8TZwY
+E9ssD4FygEj5aHjxKAuIZcUVT6OHGlFumbTpoH/glSychTlNAO/N6D0scpPebo3
1BvIemVFQb22inoXZ7/NhNYmffrgz7mZZKLRj+E4tMR06q7tiDhaDl8bkFOk98Xq
1AZXNgoABmmfIMw+rud/cydRbAELKlBASHHfFGm/f8Ygo62oGFzCCWLTHRDicL5e
reGJD+2C6uG8AdEc8+PzJw3AXW/AUrJfk6EvQZRSFb9Z33nNWQSbG7lWcjEZLjcw
hTs3FPrQd6DGhteKitDLMuG1LIzggxX/JvbqrG0RsDYZp4wKA69NL/sJDvmmz13u
jCk6ZLJ/d8BfrtNMujSogtnUUbu7/uisv2e0RqMF+s7ZaYWA3NOBHPoX/3ZcRsWo
EkaSRon1FEJWsBVsmTPjA85pcct03I568YrX7s3Vpk2J0Z0Zesnv2O0AEST7U3PG
y+9HGmC7ECwkaJkB7OETzHV/mNZwvfD0xcXvhCh+qRQDfQy6euPh9N0sHHVbFZ18
JX1xtOMQLDI5Po+TmKOpV6Xi2axZKGvpkNFpagNFBbR9H+bfNQVmPg9KW9tdQRCY
OIYkyUqv1UepiESF7WFbVQzk+VBxGuP3nT0Jf20zwOvNBMbmJ0hqV5BRgHHC35ID
LtceszoRXvqHHnoNjW5ODnLZhmJZRpFCHKoHRmyNqFr3VSCO9xSHb3jbLqws5r+U
HkcJVaqdS1qaJ8Zv+ynfdUrR3Ya0NlRBRHDNAW+jTJf3TkUBv+AN7J0stWq6V2R9
n8khCjar4zDDo6IheyN1a38asuOzYUAOgqlbuoXmd3r4CNyFKnttr0iAAFa4bZyH
PROJawwzspRc/DPmyeXV+bV8BCbkC+iU0Wh6W5RNAbkMfNnqMt+oFreTLGd0ek8/
HhFEltSqCdX85faJhu7Vlhoe8ZzSHifiEYSCKyUre5O1EeYWbF6r1gRNyjFikUoR
fIfSECyGEjHY/E9w/KTbHku5MctMz+xgFDdLtCtS2j4yPeb68gWhGK0mOeZN9+RW
vM85+mEaD67Ap0sjAM3geXV5SecMIt8VITuKmcc+wv30w6gsh5vPTN3yb9JQ7f5K
x7bRagqCx/QszV3OjziGvCtBtr8sMhQ/XIIayASZiTE6Pjf4qli6QjGm1kjCK7WZ
oGG1wV72i/x7yP8ephPWMa1f27FA9We3m21N33q4WCprX0lOuy7q9VcZ/X9cxMZ3
Md0UwOn8qoe+baC+hdTs+Lc7UdrLYKkxtFDYcTuUEz/3KX3t3FFw3iURvwG1jwCJ
qwvyDR47NOGlpyN9jl63B4+sjJ4UgJmkIROnyt8pOjzT+g0EtFKd+yM/JopoG3KS
cfkpUvhW828Rm9ElGWVKakIVo+RnW7TpsLJ5UfnXcW5gQXjtaUjA33BIaGohhyC8
12q9RU2Ujc6Ny5BqdkFmPhqbgxrFmndZ9nAp/QNCBG3GCJpcJFV6wby3wZE2Gzpd
FrDVE0Vdopa06g4Ep39QKYRoh7WMQiu9q4Jaemmd+9ecD/wXuQzK1b2cR+bqG+5v
Rq+56uOgOEJj3RAFJb469kYd+DbozRKpxgcjMoaHO/39AnfLCl1cpquImb9Rzof/
RhTd3ZMkkK3jghgKMXttj5ix8ncqG/IlJMl6nIxEqd3BSA1GJ6dHU7a8ulYuGt/T
NRL90MtvrZWwjeyGxvjXyBi/1Lt6mPIyTyal1OoTxoh5pCqtleMSRUB5K1Pa1oDY
zQ0V/lY9UJYntaysSZHrF/AYJIZw8lev+N7/hiBLtAO9YAbU5Bzq7kf5V7zBf4bb
1oYT75zrcC9sXnXi4AT8JkqM/TglurJITK/dPWGS3tBBxHEwFCsWVCAEpZVkwR83
uYnMTlELJQrcfjfVfnKvIPVpMpoHRAmBEY05qm3Cjlk1eBybe9DKG3Sr6eoQP2EF
H2p+ruCnkGNfQ1ijHPOQMUrRXGqDvUxlo6B93IhhwiRHRic2eGa1wvrrGxu44uib
+WcpS8i728/nhkyzJYRADFOm1PXPPbYiBLTxzTZce75oXQ5UbfJj+6XefGIdNrmy
hKRlolgQkCLPHRtRDFi29V+x/eVqAbuJwf03Dy0r7J0+HIKQtZNmfC+YxLxBjapv
FqvNGXT6+XVAF/vNYFCBjCt51CStM237MMfXX2+xhPBnrLicAG2/yuHnkFupn7t5
7NBP+Yg/nO1V+G99fkavBS8QTcuXuNraxEkKy/yRhKklKC6HsZ7eqyMPrNo9oL42
gVZl9QFLTRKb2nsDay2+9lCuOkgY7Rts7VYB/dyRx9INm3qY0CvfrP2BedouEdrq
GjGUEF5IJwcZ+uLPMLeBxozqN2pb9vJEPqZ1JM03241/66dvtmQrp7tD0ihJ+t4h
j20zqRR5c3L001MGBOqlh644V4S8gUAy0gnB+7TI0R4p0UtbrE0dD4u/pTOcOcyR
QqAQ6sMd90WODCp7yeaZgg/CKSPFq+fB0MlXTiagfUm/Wx+64tdyFJhkAGzMczoZ
Qn6048RZjAIVzZhPgy1+WW4gIejVuIWxx5CneBiFMEYCeV5TX6KFycaeeq6uiFXk
9MrfptJSC01Bhl/DSDiqwzF+Q7DBLUZznkZ6I/C7crPHYISB13e/upbMb9+US7Yn
X2GziQpsMNXMW1RB2lKjyhnvrnYBc0o4jhBWLuHuZj5MO7GZL0la/GJs4Qjkqi8O
jUzDB8HdxdtiPWBcmXSW7ammtFXYstqP4JQMpsIBhliuLjS9meTuiUjApmq+Y1ML
bt4H+9NG3ZpVjgV00XSax/TCkUYxEYFa9zxMbnOyuNkaobR5Tt/r5z2ygOmEOTnf
xrV9oigHOlYFqNPscevDTQMg3AuKJAKXy2ZCyyz7QsXoxG2GEl6WScwlJm4KLEWa
eV7NG787tCYQ5aOURT9LTSy/Tm7VnVLOMD5TItM8NIl7GSgHtt6nDRT+D0MYfz16
5SDfh8eh6waOCNXuDvqgZFLVANTgM22asRoB33YkWF6LpubbnaDKcGJlaKnpVXfo
g6GpEYRpvYUXvaKZGWPEHU3Uaqk0LpvXD1xoAGyuGeBgG8uLFpXeiOp6E/v0jDu7
smGNOuJ8BY+tjSnDKjSAHX3WmV+x+wZ03vX66B1gi/4wmNvkGAZOD7SiptfZ0dd/
G7FcnoUe3Z1LcA5E3t7CKa6DQBVy8oxmpvBvt8TSN0in0uCQAiQoZ4GEpRD/45c9
p9/DSWw075Z8tSbhCf1lAOmVpUsK2XZ2dAt2HzSfpGeyXYXd94XS4ETZhMWDBIiH
u7gAJD16o2oepPwtjd8kS1C0ihUtWRtPaSbOe2VG6riMTfF1XbOjd/VIpS0bKWHZ
6A6k67feMBLa6Fv6qf7SBzwoYLr2oamSdfTuS3AiBoyGs0WrS8wnk9HPGh/Xp9rt
EnaZamZzeC6VCDafy0AvQ0a3LLxpRKdaiMTF+aXEnWVZzdfp7hCFH0ljx5HHqOE2
lnBpKB6bTyYyYq6/0VV766Ndu3K+ZSJ0/rTYSkdIo4kdzOjOjfDcRzePDY3K/Icf
HjIJXOlp5WHhOotgxXVWdeErilFtsBlBh2NhgKRVgV/3N9UbMjdA9ChuJQ2o/O36
IVsSWTtUTwj7+mxySE5jAc+1uUma36JKDvxTt9kOW1eNx8bvLjXVfN1Nci+qZuB3
yZ0HIujJdOs/0QaU4UJFBlZmo2NnOfLtgioCp3k2H5+02rYPRdNSqbaAt4iekVn2
mF7uhH0i2lXUxkoFbnkTp8ei9fn4mD0B7Pkr4R/IsOmx1o6PaqaBBwUmtXdCu9Tw
2+2gslZzWIp8SdyCuPMgLRdttXiT5s9h9tRvVIu1rNdblXWFUF8Kkk3LjfFCaFWi
mfuqqROcRh2+lqW5RSyVqV7jqrE4MBnLGVCJecqX6UEbIhqtuUdMDOgssMnHHv4M
7l4g+ie1uWOehLHQAPE+g4P8JJuSX+OY3mDWXiiARrsBcVbqTIFWnn+csJI+ClbO
7pm+z3PGKEvvrAtuLTkigAM0DRsUZrg/gT/gGf8n1QdUBt6swXEoYhNfPxNiiGX6
j73YY1QYdopePDoz2EDTffZLT91tQfXikcO7TQ5GVpfWbL8vUh7ziaLkj6I48fLF
H2pQmqqdGa3Kqc04og7z8auLZyRVwh/sWped2/KnJuTy549fIicI22WWP78gi4Ht
0Ji4XDDnqCrmCRF8+K7CL3YT6cWRceLBObMkRxgd5cZMpqFFjH+KjkNRYDJAqnAt
PPnHZfBLMm+br5G6Zq0j2hhvUmRAnqppUuFU446U7Sg+Q/3klzin4plbEcFUec56
WNNc66hMrm0RRvSL83y9isRIrlG5C2rSLAYACaTa7YXJqErVI/UCfJYLN85Wjz4G
+YLe+gcf2DywqwdBlWwVvAR138EL0aWmtmK4aWFUoEN+Emh+tqlU6oWyYprckr54
5unYsfdveXpFBWw85+1yYTmLedBsUDiLF363m+50cxiUCMtq5+YTPjl/GOfrYNMn
z8pRjW/LoY+C4TpYpSTrU80gO7b+XwoXsRctoF+bjqPrsVuFcfBEmNfJNoMLN6G+
lLnUZglWjG6gd43zJRgDaF5fE6VrZrjMkyCyu+TnBl+3RACy4vP8r6zLY7L87W6D
nWp7DaQuYJnam4vyehiwrb+oHw/XU3H9k9SZ5TSZnrmMq/FYkirKZ7cZnleYymMr
CyDXUMaW5db8daCecH1tk0eK0IQBXzKaD2EEIfpq0lfzM5idGbn5TvpLaYUyx1St
lpkfTY/V60SPkbGCl2IqaK4Rf+vY+BrBtK0cW1Emvb4OayxArEhSGKqPBKYsfkWl
Y+UgM3FPO0GZzFVFRyqtwUNv756ct9z9EDyI+KyjuZX8Y+x1cC4KifUf0xh3QVjj
btm/4x1tlva5c2tL1f1MPo2P2u6IQlbeeQAnTXuWhKUWeU0ExHEFF8XXw87WQt0T
vkp4VeK/CirqS57t5Qfv4rbVyIAfYWMcRQsNKRmlZ1+wAvTapj3d+/kmyw1rhIQV
NaRZowOFxBuKyDpEGHByI5YNzMiJQRiXQ4vJuGcUr5/nEBB+dJNOPKgKQPWwiUlD
54+037/lfjSxegOIhJbGq5Luutj3BGurz8ALtAnookTmKkD2ccGWRv69G3OJX83I
wgMz/0wwGlakZhQyzumTD+kltoa7G/XzeKcEJm2G2JBYkiNtMV+6b03CESDM+hpT
9l7bwJyzHEZkKsdIXL+u0RArkWwiTc+pJiwF4acV/wnYebiJbbE6zoo8XxeZKQKB
HThp+Ta6dTdODHrhsIcKLkhmKHQD8IISNlSvi1TOQQxXpYb+Ak6R5Dhj4WuRQrGr
FRMBGkKvDCepUdi1MLIWDR/H7nuSxFEup2KFpmh5Yu1dZ7kn9YZTDQn5LcAR+aUd
IL4AGQs4kWId2e0Ei8C3phTUyucxjtfR5eAsFzdFm/ZGwocJEI24us3ULCYyFkJx
jG7FUUjI82pu+CHyQ61VTFrBWbzsGNqL5YG+Ye6nTgnGZBl92zoE2wrMzHkJ7Ddx
gwTXzeWMtAbtUkHxIyglAQ3eZi3vpMeBoJ8rIZnxZ6+vK3om+XNv8Kzcd0LjYZUA
a4b0VGhz4iXUCDXBlSuD6g52xlwaQH4nOAYoWEtIupuW9dHQr0UUIEy7hL+qhthU
Q3MyhSF0XStW6IGO2OSIUu8P1pOFgsQN/8pC2QWKiRVEeuCxVCArDtLw+fhF9k5S
XsDB98AbANTQNHMdLlVW1ziyUKMoGr81TfzafVMRqo0TtFV1mcCzVg9Z7cr1C8on
90tmH3O013NZL6NZhkAEIny2mjJcE2FY1v2Pv/dK+EWY3gbcvhf1YcTQdcTBVngq
ctuooOaWj1n15s4iEeznOQkhZgxaIsh516exPYUc4LxX002EgUEqWjgYGeXcxcIo
j6QKVsGuPOPz8gjv8++pzgBmG7q9nt7Ty9Xnhc1MLoPpQLzKp8Fl5FENOcq0AFxP
v1LFOzeKpx8lozGbIn5zCKb16dw3chUn0B76akZhSTzf+zizasGObhBDTEXflr1n
qZ5i3tROSBbO+zv9uaDFvk/7yLtSL/Nj49K189LlmRvKES7HLQ0+k6g72KYg0LlU
F5on0ye85u/OxJAwwuPVlkTjXEKHm2eeibXPeA0Wgu8/inBJ+dJPSPPr+zcWQMgG
ksPxbp9ySYuhG09U0iFYLFUd2jZIu1seC8JM+y4toKvCFAuJQLyTnmEaHhTK7CCk
lHKA/uNTkynRM+4g1b/k2DrmNLoGbfbFICHIVJaNgumyoK3fct6ENGdu9P3EWPK0
lM2U1YUw2LEZHhiwaDI0GtOhVKLo9DWUm/iVfH6oNTTGI1+TIptzADkh4iGQNvTr
k3Yo5emcogyo7xvyu5V/IEZQaLblHbOjX/EFuyTabfB+svrgPsn+RyCm3SXM/gWc
iwoEfTw1MF9fjf9AIDRPkwBFpF5yT2CnkWPOHSwYbADdWyvLsteX3KETG2Kg6Ifg
Sb9g0Q8ZwZ+9D008/C7L4pVjn46EZEDdPkMvbcz/bod09u72JKOlWnyyHYa0jhRg
7PxXArcqBePRqaEGhHTJv1WzpODUBDMDE0VVKmcmzIvdnyDFsdvlo/uf3fq3chQX
vZqPnoueTAVETbXCCd8adkKNpvRy9XAdEYcpZUuVXIjIYp8YZfx8ggGNHUOjEUQI
X5moBNQh04hsZ1RfRcIY6SG5DcEV73us88kaj+wlVGrvnUTwlvrMRqaI18a9mSCm
WDoXf8SFFjic4fLTjzUH3xdB78fhltAFMO9HZhV9NzBt80V/MjqoXbUmRh6slh34
ZINexhkbaqC4TLErFuREANizR+Wx66OwHGKoiXMOh814BmY4pm+gxfj8tQVfPCSh
ezxEXm6o76Q2izL+vo6Ir0L/L9Tva6YwE8yj+A6pOYX5/88useOuxcSBBn80mjpr
NbX+kKzg7QpZ2Ps3Ul8NRxiVTbfNae3tKLQzv5SeO8O8MUAHcgP583DmmcJSrE2d
VOQE8LWV+b08bJ1bM8jFanc3l6ZqztsLw5Wvb72qjBxXg8Lsq4Mt2N2YgIV4a3a4
f6OaM4lN/V4nY8Uc3cpfvG7/x1Qi0WwZjXJQe7PhflkjaA7zJCTshHkU/04+2ngV
OAlyYQCTQFE9poS8XZuf+f3O3aQkHLIAuO60NLdxv1ev9AKIM81uL4VAR3uth2Hc
9xqoetnC+Zi9Pz7XG6d3WS/P5CqI8RypImH63IrGSL8rtzyWmi+hj3v/7xtwIhjB
tf9UEJZsvegxT0zzxRBybKTC7v2UtrLI/pP8D8Y2KdfTRzvfWal1eudWaVc6GVP2
CzqzG7W91J+WFZ3AfNyW0+tuKJNR1KJ8NUtsMzLhQlWYsM6OU83NlbY7NFJSqeCH
UPtfpkeX8k21KGfCOnBAiByXGNdJ8XpoC4Mwlqv/SOKVGPqhwGQFvq2hjeETuQ0O
RpHDu+9ZhGssnUePNxszu5coiuwvHW4V8qwYUZcnofqJryEcpmS3k3t0BZMOHZ1p
4SESyZ4fqjzbeXmBnBlSt8Q7y/iokLoNERFeDkuhlgM1BwxMuwdgOd0ZBLenFgUx
ZsSq+/oawXC9JuCU4K1xTUIRGwy//zi+QSAgtLXbqv4ixfK2IIgXccynFTL6+pYU
mApme/L3FwEcPTcaiuSplTIDuwuWNPiVdPJD/BBw53q5MqueO7rPrV+cUTjDKF4H
avS544b/YtbVCsVAZasfvNtorGIokdj+EZs1EYYitdqfJ+/ZjraMby+oZPqEwJzX
oRyotcCd0U2MZL8R/B5UhIGDLVhyPDFNZsFhW1XjXivXOiV5lulssqiYOFCMNF5s
NKHC9Qa9nVMHSK0J+ro0Y7aSSQggqpQQ44+Xqz3f/Y+GEEbykkHCeR4WhlXzxGDF
mkbl9PaLxBOSMSRaA1JB5/dgffuBoAFjSlYnu6+0FDJXVV3hd16+9nN7BQp198/h
6eyVtBOBXNopT3lUIBy7g0CnVwZ1Am3LjuyyH1dW/UlLLNm+Z1+Ow+CYbI8StStN
YDiUI4/jRifWrwiw/k9PhMenesyXJJZuNQaLFQ8qboC92s2CrjuyXzlQ4VcLaViK
LfwZCTucBugMd3saPqXrfdD0dcL4bX4PZgU2gFhZVOd9McKRIzxYsDmP/P6vuFtT
FjSDWL/4yDdIcnub3Hl0mi80vna8IskiEV7qWB9GFxnNYqnYE0xxH6pdzqzzI3FE
PjofDzaucxPSiGA6un+u3doVCdSfeW3+NeAhDhUvJrvzQ4THWgS+SB7gdyG2zJb2
dhp7oFQx3OsUGSfTPaNgX2FQgZl9xuj7UFl4KVz/aRQ7pihpNhG4kAiW8hYqHdAn
UyfwW2mHZ4rC+IN2T4s4IPe3m79ESgC8KcYOn9tLrQDtACC2UYdjEd37FiEDLJj9
eprb/U8CPw09AaT47exieD4UtRGS7pwlc31i/nBjF/RxdNa1PoAaBOLrrX+jFHQy
hNsOt3/IThZYTUAO60KKjKddhtQhdzCphdaisPmR6TU42AQuH3wa4Yr9V7pblOQx
xFKS+g33zRSqtpDKsCWD7SYP7xO4EeooA7Yox5/pnYQsJvxlYCtFSFQ/RYfH1Eru
Wpf2DoJSHKe58HwgnQWfEaQRvRs8WK7jUvOYeqdtyTt5rvBQQ6Xaqcsa19J71k5M
Q7FBD9o4vk4TMLAY7GW3ZIl+XEPon7UU7Sz35VUSkO6zJuB0ryadd5oCWfHeKTwQ
TNiGQqobqaZyqIsr35xxmb00iQOErE0qTTh7Fmic/KpwenTtG6CHJKO7Zw4ar9Zg
56VCtOro1c9SDveK1dLcZdzDaD4SRjjKg0LxJSrBZlf8bzc0FWMFqZYt2hyhpRnb
4SBL4pdcX4V9dGUS3BKicVMpidS7267YHWsVPa9ea/RrPrZTd5EnIz7pa6yZ1Ad8
eSvsH9Ar02XlutI8ecvTLXZ1k8dRPct9fvgYZi65ES/ENWUSfv9OZp9mciopxNHB
qd0EN/14EN0QwrNLcf5AoQZCJxFUpvn6C8T71sdfp2PHbVQ4gw5LVdG4LK1NQvQm
+jSrMgMSsVJKwaX3GqvIWLiGir5OqQHX4vBus2a5+KTdmL1x08cWke18AzlM7zZe
T83JX3VuNYyL3i4Bq3E9gQNe+NrxW6JPPftEtFCyDTS7v53TSk487EPf5wG8rtdj
DH7xBhpMKzN+LED4b18mRJQwnhz/wLhAMnmHRnFbjKtatf8sQ4F1pWR5IRuEHrhi
dmnX8w5FiCkyTUBwsSQtkbNrUBn8Wwt0hKSvN/K1kgvPxoXobIXJv2FjGISwpAw2
nhUXKEkOsqIyyfudewiOlKXMROUc6TkN0aVAupD+UWYd46QwF1eFLCj/fXGjyAtw
TAUcxNdPdI9sRMiSgbjlqsTO8zhno4YflKNqk9T2bm/yiAWUlGmPEf5DvpduSeGI
frmIQWSA3W/dk08ng1y3EFPP8iYEUCZXlGBOzjGbwI+Bkc0NecGZkeXHNS34QpJf
dlgu8dBKLW2bKZ6SL01HR3uyNKXHLpZW8TM8OBUZkMy02KP39gdbtqa1L2Tou7fR
1qxOp1MTHfK9bqShUKZBGrN2v5TKI2OeDh3tXqovkoXpdZTSF+lVEQGahDG29Oct
M54p5RxwENSHz5eJnpUoaxFyrJDuUcIQQdAhZZrsPB9SGhIUi4RzEHw9h0CY1+xY
WoyFsUpNLBNxkw470ue7gdAJ85wzabnTSw1XXGNCLwcRf4QDjLHi2YDsB3MN9x24
KdtMkkRe18Qev72ibomZODFoNO1xPPTl4qd4F9jECKywy5aIvOfhWyMMpsY7Fkjb
kb21N4tteCUJ/C1kt0nYY7Cn//F2WU8oFGg97YWtAtW5JJXwnH32J8y3lfTjHr6O
twYo7ubv04DCNKMIQ3DD13A7p/02zrnnOuBjWEIEUUTNWLn+m69qvzclbexaITQ3
fKo6ouUtuAlpY2QB7TXAWcKBGFHxZHqotb5SlsOIE3t4nys/fbhZ1y3Q7YN1SYy3
azVXLRN6xsf+LZNAM1XlGEoqlLdk4Y2iu6ziP5VDn1KGCOcqzG/9AiACpfkNHsZu
QHKDni+3rQpesA4BJDPBcM4XIqxSptAVagCHcsusRYUoUT4rAgK0HYNiLIGwJzvN
9X8OnqzNVcqC7wO/yTB9AfhaFKgLMq/6sci4QIffZPRg1XD3ESCXzaRzRDTSBhzD
cCjyXJsQ2O0rooNlhEDyqVW3WFImLWmSFZPNi+UEWVtfPP29UYEF8iiFPk82Q01T
ynJqGZTn+HF/3tgLBVpC2tfcAcSqazOpH7KcU5GyfjyKiIcj0bcUcmkVDBclJa7g
55lyaKYQeXghHgV5LnXSBOdSavETuD7YrkOzXRR0WMKZZZ7R4BbbF50oZcDmL/+y
d7K/Jnbh8fjQMjGkN3MqXS5KvDIawszXowwIa64S4KVgxePaz/mb1u69geOi9JrE
SHfeWO7Oj/6ePupvQFXDApaEhl01R9Wq7DPNcWRBytcnI6cq5xCs7lnOSykr1cic
s0oXLWaqgpEkjm6hYUVv+xPO6MsnCe7576HcVogX0BUddR3vhwr8eWWbgii4Qt5G
ZioJ+VM8FCyk23PVAQGHKbPerUPB8Mulm2OMiQSIqFDT19R4U+HpEjM9nv/sOZ2S
NUe3w1bfMmHTU9+/aKjs16stftif5XS/Pc8cAYTuEdfaNLtzZG/pwJlbdEUG6wvc
9NGyaB9KXMenFSgmzziw04RFuFKlzPqbm0DHGXWo2x/P1yFN1ZZxKBDQOa42o8kk
9ohDESbBao30tSJ2tFkhDi1JByyA53Bu6oiVtpSgM1Sj9Hgii3vGxFZ+VmpOok77
hcNDdbmOq6DT7rgf54gmmb9VK22DHteD+1eUe2RuO11liDmVhCjqw0gIP0HTtvwo
VNtKjNnq8C+k0K5CvdSdohaD5Bl5jkWJazORaD3hRaxeECJzURNipcVD/dz9FuA0
foakAuKSD5DaqdZHxaFDNi+DJR7TQKXqXzQqnP6oGjecfHqCfcdm8Ms/rExSzKCa
uYpm2ShRwt58/Rgjki1LJQUW3qzH1gWgF1oHBmFXrLNpfd7X18kyvmZOiJVBaQ+5
+y4aZenWecQGGzJvqOL+ke95/q7/EmRh+JN55wlBy/J67lUMceVKUvx0mw9iaUyC
AK2vlYZiehMgiMJP5MVIN59y/fmMSUXseE0ipomiWLxBQoJGAzSkmRNbXLUJfFOy
NBWSviU/zJLunn1d/eWvKvVxwtPSJrtb6IZ1MljXDX55X8Q1p639uwiAKbT+y2WN
vQ+CGk33wK+XRXR5k0maiWb4mobAVcf/Lz9bliR0m4hjBhbCDG96GEsigBZrlbxY
Cq3NhyVWSuzv/99fIaSbTnOZaENbyupC2NnyPxER2NcRNSjvLD4FB6q9uhBUjYHy
vGnUh8sqy11oGv6prhxBA9Gc4YZsKnXzAzoNjiu6qz5RlzpEM5QlXwnVTxQzngqX
z7dHMMpTd7dxuusGFbkZFfdA9fUNH0o9CGoOwXC0//tzDT+I53/xAarbapSNLsxY
GTtzsLuJCjmT0c8gOKNlOZhN4jbLo1ObIdMXUcI6gIJfIxYaWuFSRuCFDWS0aIYc
Zscqho4nwhT8HXcxTgsW2jwRh6fqswZZRsPB1oiEen8n7qMvxXxXetu+y5ZuFran
EES2NJF+c7bCyBmaAPDLGWhsodqrxmeU33ujp7iWNWanD7JGb8gdqZr9znWpuzfx
zgF9TZD2Wn4D/N2JOKkXOefgZ6TzR+GteWKmGlAFgq/qQYAmXKBRdvZqZn+mc8tQ
W9XiYrL8pVaqJ3+65tkCKgGo8ybQB5mlzmpAX//+IDATGjrZt0k25nthdZVwr81I
gXS6Ao8Fq1E5jl3ZcjzOzFpSIxiIpff8nuFFxzPMyAl5Km8MsJOJ8JEA6m5aNBJm
xG8Ybxsvz5v4GjHN2errCgotCH1z0Sz1DDXy1lYzeTdEWdU/FCbzFQ5NkAxY6bkY
Rds/Rm9eaMSqn3nMfx1ByaNyTLDtWNnyY5FvM7UBzW8QuPY7eoU8+0qUkS9CgQnI
M6RFFVE/aLY22Au9jmMlI9x3kthvcq2ZbS7EFUQ+LyZT6mlk+e2Vf0ocGOV5gp7Z
9y00SG6Gmt3h4LSPaaAEHzMiKl/tWGXwQZN8DBFxLr8kCPQEJKeSTHS16UWZDEYy
ysaAHFZX/bPX9SO7T+mU1UCEPnkVvNwIc77x65+KFEm4EcFwN0DRQWx0STX4txrZ
MFJg7YZ3IF+8I7QmdTfJtFe2VRD6sCPfoNRjBe0bnDjbU57SB4aLfVw767tpgrIB
lPomEecwiL9V/I4TYKxWGmxMQtqh59CNXgMku6hvVDRXbP4B4O4kdXXsH38BcYCT
md0M1HkuOJev0KoIZOvQ/YJABKRh1hf3LoWA7CQLgXRSmpXYRhI4Z6UelVzVMGnH
MyBZvfiEAD7EbgjzWIpXuonSJxPjBNmBMeSreNqWTWLdLf6ZB44hIUX5fKHLXpXf
EcwGE3ONh/cPfChHe2YXXbQWBK/oaKEwSBarthXGwJk05onC4o9syfyrswMRW6Hk
5oL09RHZoC3MQPUI08Rd6HsLKG5pNi+nHtzC+n9ObnD8PVlDecJAV1NiqFzx/N6V
HuLNgRnf2fdiT9RCTcHNK//MDdYbTUM0aNcjVsjbYcFigiTJE266AE7OEzgkHhT9
l8kxxLFnppiWqgSrRjUtK1EVHm287fGeK0nbpyp8DPxRYvwlrmVG2m1huUZ2iP/n
y5/fkc8yjBbNN9NYocBRo3XEaZXsYyt3bI7IOUrxlCSkC5BiLs0cP2bg76sXRiTd
r5N7ULuetHnmDA3EZKFP2tCWGtXElva5/uDwodmW6VfMkzI0nELUp4Y4VpxLFP3D
IVgwkXoN/QEEuPQ0A6fiulJ+gwXPOcslTolmKxQDkAyMSC3fHQsRvT6JArs6pVCu
QuymonISP1M/kYrINoz/Y0LmY7TypFT0Kfq8vnh1FzXdPtHmLv6X+El1F5uZXMa6
euAs9S/V2vx5sRKGjyXuu3K4sEtF+Q686OKl6G92LOCLeNB4wXBb9Ru9sSwr6TPP
kknKzXaCjJnq5yx4emmtEOI0/Xx9SBU2NvpBsAEnRUoYDxrpsAC7BVITODn13nIg
nL8ofXvZbJiqfk8ASBJM+cgLz/zDgZtl2T4JdoACb2VTamtkSyW7dqBLWfLZMo29
QZq9NHliN9WHR9klxzw8xUBQTBCuTGW0DjkbUHcQwufn65fiDU8e3H72H1FAZOYB
bLot/hWsuX53Tn+tL5H+Z51cU9AuetuThdHDSDvRWTMbwvtfNIFM0FvyRjkaVCww
o/aUWaPvhZLKIT+bZjoYx/untgyTg5FhCm0gN4Uk4MwA8GmSOlbSXoW4Ym+pWvcv
zlloQgBa8E4CuVPED0BYIv0wPyjTLPhplKcuV6y8JV2WO5WQikIemvtPPvEHC1dM
0iI5y8MaXA2ZTSXem+fVs/mkJz/pxYJFhU8c2oBbY5BnZ6doj2lXrkIrXFyEe9bt
0qopqiDvFkAYm6oiu3O5A9nmTtbFxzH7Z81WT8fQMmELwkbcpBmb1puY+RXfzxug
NurmVrDfSGwg4DjOx4/sBQ1A/ueCUj/BrvBnGlVOSButRsORnuZZ5bpUJBNessR7
iPL+rz3MisLSyzg1bbgMTi91qODo5Jymt6xN7qP+QcAQ1msFyICs3VbC9vi2ba1F
We0zNvFn/gsgUSPzSjC0n0wT+ZAqFBJKGY7bEuRY301fvQQCmPvBM+PmmO22uoeM
l/QPtQQQA+2j8CTGGw/qq+MRhFZRQSPuft99USCfH2SSakDTZErTdZ3ChVXZW37v
LgzRbrBkzt+E6yXFkXliV0ODLXeiqFiR6OPj9d+M9/MtHQm2rLu+2XWKMgEmjgaL
9kCoee3sh4vQCR5jnOzdF6l5kwHYKWJ1v6T5/gwaa5OaE1QIT/Gwr+wJaEyRWR2f
8YchPucAWSoKi1OGezBd5LqIGDu4j8O0OeVR0yQj+WqueEtJ+4Nlk0ucpVKV7Iwg
DF5vs8T6zJg4ZJuPWcwjDFby6IQc/JLBzbvMZUPBZI1ZOB7lymHkfPLCj4gkR5hr
qFZtYFTcEiyoKHiz7b3NOvWqjcrQyA2So2A2SvQby32x3RXOs2z/dG98mzATPO9W
NGbxkeGh/9ggKLaSRoDsClot94Zar3YZFmu1tu8WFIOBwHyeGSj80tx4/A4TgHqj
wsCaEWV3D7xWw7rGsfJnCRsMTB68nBGX/KYoVpxXRdBJSf3Qh9O7Am//GxlVpXDu
VVjj2ayyVDvoEI4PTgDjjDehC3g9h3xoUurrtsJNK/d9cX7g6XCA8OAmk5MpNDlJ
cM3gXR5nDuex9e+b9L8tm1GcMmhVCic6GkgwHoRysrjrc/vCpOc9t7zMn6hRqxFc
jvYekE0514ym5+VSD9TewLZQWO68+w6I1N1GnCyETF/dOwrcfwi9LxErwSqqTJZ4
IucQmFheQ+NObdl81hnotFmybX8c9euB28UBZ1ajp+9qZl+oY517f+InS5mS3ss3
geEfuVd+jgITjq3ZV+gbHhM1KaWW3nluUUJ5sX5+R8oT7cN2Tx4crt7as9hzU3NC
n/ajHwvON2LqN41pjlhDB0ygGoIyfkMGH/SRWzE6wTnUyxivvUwjiSCCshLnwDV8
0Ep8w/8i6QP7bhFAPmyNk9QklbmC/lBm0gh+HpJBHeis+AjqY9QgplVgVrD88KYe
Zn3YcCG6p706pP66fNP6SJRgs+fI8LBgHk82iTs/WwhSj6rAoju7q5teyZKaKYXE
4R9jfEmc+ESFCCEfAgFsoD5xlEo1yF7MIM+a69aVd6RssIPI+625t646L6gjquTx
Ty43cqBwd4wcLwOuPA9lXSM/XIcmzawDd+Ou34VskT38wZG8Q/MjYeSai6O0Fbvb
fCMvP3GEYoqUDMqR9UBHHGXhv6Wm7RkfwIoZ+yK03DXJFtrlXvL4K9i/b//uVzoI
+EUSAtEnD1Ih5y/Kp3YYBxCBJj0TTVdwelbk5/zHvjUgInhweaq4DxoLnxjQUcZb
LzFDFxys5/6M5dn9plw+V/3vmYOneXv45RzkUrMBvrqfjaPVlCPW96JRHv2IbAR8
XB9ootXARJ+PZ12mVWrwa7HvYDJ0idELRr/5nVxlGmVRihhy8z12pofxNmgB9Pfv
ZM17fbZN0p7e/MPqu5UpvapmMQ1yoMrIHth0fNdE1NRB/SkrKuDbDl9a/UY+1nE0
mLBTecccJ2MQ7RhpLS77E4UJw1Im9Siq3MlrjDOwdMNOrqx86Zd3SPXDuueuKMrV
QfklLgdk0w99/wmVkQU327KBNAyzr+1wdfLRy6MsEc1NazgJcOSWmPmJgLWz/Th6
+ufyYolpofdRfZGcqVwTTjXISaDuGwpQDPrn3xVURrf5OrLpaauNO16D6Xj0XwJw
omWUx7tZ7lpY5YbOncI0ME5nK9m0jiuISzb+Obfxnevmo7I99Lw0UAb45mMBK5Xd
oA0YZb+6JkQAF007B9tBeoyqQUxPTXlgRakZt1YErFeA0KfGjke+CUMSl3bTclR+
bZhuZ0PSWV3TvGUPa8yneaAskuDUQrycmBG5XXJDRTbZ8fTopGHtQZc/nWqsGa2T
BtoEKG2DQTvb7qY2xjeZOeNcviO/kkIdtg0oI9ddE8rc9+6/CU6C19PjCp4je7x+
5cjcjGvHx3Is4SrCQASiPSjViOSKxZIvInNYhOAWYte1NYVg07l/hJzJ/k5/pkFv
7xt7itKq+arlnxwLOARoDyp7a3DFvPJ+/UKgSDTHaP1dtvDbpXTKnbxOzuP9DJUS
8X752STQJNAlfe/Y5q6yUKq0XZbLimM9w4mD9AT0P6ImWhGTpxJJf0jqqH5AYWHV
94DkxOvhsKagrXzb0FBS07AagVg3F9y6cgKoyTqNYI+qqAK7yAgz06d9oIKE/plb
40CSXbs+X9djZgUAkoY82866gTEKHw7KImrcEZLd43qkb8B43KBE/52UudToXB5h
MP6q2snQMbOaByVFj9uviHVNGn5pQzIoeYSbYk8X5v0Vit3JlkVoD2+ypnyQBeRA
cv8rTAzk5Rrl+QriOZBuy/YHDFJllN42H2eh0e09dXzRcmxWh4fpk6FDYd0FIk0k
9B6W0WtNZBcFaTSEL5mGr1rUAbCR+lmr3uLQaRS4CqGtMcpq+4Thk+lawZHxx/m1
HVtCOOAoUS40m5TUW/Un0NixnTs3jbT1SQr7AzYX0A2Rw5wgrN04p/g/iQpkjLXY
ixunNHxgN3kI8ImpPcL6HIvaRYPAl18tfEgdIU2pqp5CH36b/J3nhHAyu5DGMwYM
m+OLsAvStDK8ksHbRf5kRx6b/OQi/zDvlBs8d/Pw/2AIXj3+dhL5gxam4x4Ft9Re
L0mKrm/JY3qvop6Dz+ST16aQzUExRkWq8fYHLMzATR2/pMC88xIxz+iRmqaH2XPQ
CS9fb0SKKZBBL802gId+eMhvDyq7oZJAC/IsHPxq7Q8pc0MmKCyE5+LrwvpaRBUo
XZmemm5r/4O+4xNfJz2thhM5DoVUjnBICwK0Ck8vlHVJiXHshAgJ9zarlUCraIsL
dcQfsnR6CFkN8HuuWmyxpI5F5vk2fbbJL0bvySo7zT9FrU3lQtvT+UapQbWlWIMD
obvoR9FUZa/Er8czPSA62eij1Uu7YX/lQyuRGX0PNe4WOXkaT/foRh/VCh+3N0I9
EF5bXfQhDPb8naGHPgn6j3kUV7k8DVHbPCj1OKl2Oeo2fbTZyDkxRqCuQrzsYmte
jnr/9+oDRfgief0K19StzK1MCCArk37pe3HpultVYi6CGFSn65Vj5FQ/BMy4azAh
SSsMcV7uzL5TsB0iS+ALAZGRKeMjptPwLCNCXMNADnct12478wyBjE7eKVcK9oVr
A+yAZvOYU32VlJy79h1wN+qWBYDf31STFHU4XqApTaYBK3rIJ6L5HeX9nMpu08c4
nsWxkET6MvfarirXY03MxaTnvIvUrd0ggGIddc5Cd/x8IeYWx3RwuTc5Y/gUKKow
o0n+lvw47do5g6aDTpsp7SsXeIsGvpHMPnySuUV85nEECbQtEMS9tQyyNFHvA3YJ
sgdZdQRtEi0SUxKHgxMQ2WBC6FdHOAIV/gFkx2owX7uZ0FLl4hi0WcBbBoHrQOl2
4HRR7GcWYE5gEG4S+G+dAcWUS4dtPuYU+nNA4jdoxmFQJU8BU/ginCX72dapMg5D
0ycIUrPHWMVc1Tdf9s+ssmFE7BqqWt0qG2syDAqmBcjk2BkWbyf1RNCjk6waH8fy
m3yyoWIM+jC4BTsbcqqwou8xUS1Ccdwc6Aq2M6xBzJ4tt0/nagvJBvorSIRPNwU4
se9pMshXWNGWcp/SdKyGNKLdHj0krEbaNwQO2ioHH1sZklCyj5CTvKNbMpi5ycgi
YkzcXsLsjgeMOIFszZfCjS8iINgzvBzWVFmeYxUPEi1Dm+dE9OsCoDJ1ei8GAdkp
bK5EDkNgIm/XXI+cDjBg4w9h6wmcwPwhFOvFyd7V/XtR2x3fIbrfzV+vezGqMDWG
AqaT0L0Q1IeRfv+V1uwbrg5+xx6Ghjw8aRSCsXzuTNh9fDvhiZn5dIfzZKd0CGpF
7eAZpBUXyLlBIeLyzQlRsFI1g3x8y9H8DQpF9vKN8yAEDligDMtp+FgD03Z6QOJb
SZDTO0RoYU/BAnxLGxyzCDNBA8SEGgPCF2Bz3+D6eIvfG3D+VjzD6adINuubY6Mf
A7nWX9Ak/B25pU2zi7WVHhTgkzv3m96AqUbaAj8v14vAp43wBWIHzR7xmbSzauMP
A35Mdr7x1M3OwYcmmfVK9FmBtRFsjKyGdLcNwy2/854JJGuoofXnLwL0wy2Qhvz8
P0EGj9D1MbjUokI9zvOVBTzAT+fiQw8lQ8q+gvrzLhPJOc+kGqU84RjwOZqpLw4d
tpJtfGt5740GEzYIFgz/AcjgCUXxPy2ZIwoFqIhXmeLbPfn4rB4dpYbZeVWREq0P
j69F/tCbJEgbZlXzbkeu2tF6rSGphalg9BEP33jNckVJFAvK+46KXLtu4ZRwOiwa
KHM8bP3oHZFqNNomPL88DdWuwl6cs1yn1CeSlrQcifoEf6rel7Deu3JtGMIXZRFS
aACniBHzz2fdCziFxNqHxNowwD1XSfqgXYxw2GMkEK93wZ+XYavL2DFdJNGD4qpI
o26CiPW1UMJy0aNSIhkzu19mn/7IeIMj/PCXhYmJSsMRTY79b5ZW1CXz3l5vd5id
PM2rMm1qcYLLNdFR3SwTBmrDA818P7VK2OV1hEwZacU5T+ggWcmp2/58U5SXSI7N
zCIv4FrvO585RNMB5AWWkekhuUv3J5NJbaiEIr5caB669W3evVD8SU+KeYZ5OMRq
Mn5GI5MFYUHizxZl0nbQNPpXjg1MowXoZQzAvS3JhkxenMzhESSDVzEz0nZVkYIB
r38pWPhxVt6FetP1dct9DkQUGJB57sPKVcD8js9H4MLuYW26ArnQRS/ttSnLz1kH
S7c+uUdabAHLO8SrFp7+IcSf/WGjp+Y/tO7ZeeERLmBvOceVTvjS9wb+k+J4z8hW
Z2TOhancMb5H02eUr+iIHdetDNCrcf8sf0AskxhtpNjMDEWGI7UHW3ntLXOkWFQN
jJJ/TguixIXNIEpj/O4cE+L4t8TDx8CwBk5hJJuITCnV23fZohRWD0/b0fyGasIY
wzD7j2bMdXcmCqcA/r7oFWlmNl9NcHAkYdOAzHLfpzXpeL4SbbJtDn7pyU/hwSUS
RUOfbnEomHuIsmfRYWNg1a/bRxQSQ5n3j4Z43cmf/thzBSTqIdfoyEiS6L8FxZWS
wYu9joWwmyysVP35kCIZOj95vv/+ytZwf4jJvxfgvPkCqy/apNxxFZVMTZUCIQxN
uWq0jiCafDWrtQOj2u2PzV+A9YVa9tvZKT0z6eGu/ep1eSGdL+VFOHyLTr15WbI7
OoX8OF0oQVjHJ3Dc8HsuQC7oAkkfktoUaS2dqb+7DDDZuQiM5rcUrR/P3Ck1Qp4E
qR9ckkzC2SFbKRYh6RVzq9w3VBPFzxXN99bvNFjsRXICpFCpY4vQnQTAXvVW4fGN
hq0gZPxKokJcvTdQvXZ0rNIbj77szutK+YHfGwG9vsynEBTJwjvFbG0OcPaQCe1s
uA+fttfHyWAs6Y4xZsJL+7Zj6CZYoJAkFvXDmWwcu0lHBuCYNY5fPUN5xNdnwxgx
8D7Jf+uKSnJnsrOGPvo1b+nXscZS81qpama9U6tbl9oUxjvXdo12Q80fPO+fB6vX
ysJP9OUlLxFr6F1PUxZGVxj1Sap0PY/TZ9OnMuPmNleJ5EZWUpdQw+dpFXkiFYnz
fjLkXHWiRWKWuTQF8BopNXOFj1Q6nIkNUrLN48OnLOUnQyDVGrZ4Xfn+0f5IDmmu
kKJldkJxAGaTsKMq5l/pssSFYHN/YKtRS0YJovzGp83SlgI3ax5jNAzYuS32xPWS
U3azPj2+0NQnyZ7OicsJVpCltOcFefv0/t1jwL62vB4gg2mcoAmbWKUzn7ljgIlV
TzzbBiCg+Spx/3zXzXByw1VDecbklkWY0uemyQKoHYNws4uGEIzp9CciMNLIqoFq
5UbWksDDe43w4j39RnLjOxZfd0acM9wdB8iilU+ym6XwnbnRsDRBvtPy7xygYN2G
wjA0L2LkdlYjn8+VZ1myVVseudxe71YAio0qQpJl0dtEBCQxSHy4zw5pvaaMddTi
jjEm+jYnB9Nqb24XATtEIr06DLbYAwnIciUPwsCFJV5NJnZ1sK2/mkAsnLG8NqBw
mZGjx+inhW8IOdlp+NWrSqtwamMrgoM4NQ+I2K6VBChVTIHahWgzngFEI7f9hf+2
qW5Ta3fJjg96RW5bM2Y6gsx9J8E77FGBfUs7uQImB0sdqHOsmCViedcKBbavxERt
Fi6a0Dv2POBvs4SmZUgfrIE/845SnDojeLwuzfAJ06JQrpAJFEcEFm1ce0DSLphR
OF8q7VGWE65pzWU+wdXhdXB8dnVqvnb/xP1YNKdcTRZESQgjFLekzTkjDAtKXdUn
4CDOOR/MQCADTQZ6hsxmEUOHGZ569d9gDdHEpcghOJUzQuBAGCehDEs+Pqlro5gJ
7AxDvkp6je6YCoMP2X7ZhOq/pAbHeluEZSEtmHvddLTpaC2Ac5z2KLZQOVbmVB6R
g9oepAKXUl/r4CkBRol9Kj53BTKcdVt/t7wuWER4SUaXXVATyeiMRQtPTyKgy20I
EbMgLrr1LFwHzi5ysA03bYd1vFfWvnF7ILzCLiptycqy+NvWUibuazFONjexcNbP
wF2ZF2VGuTKI71f0VVGDByc6qM+UQ3fxs1/bkjTjc31eVDvOdNSS+kATnMMeMr0e
qkVJHgZ8Yp0gQki7K0M9mXWr2wgdkmGVV0c8Go+mdvNdfzeEWOnUyrGXe1w+R4n4
uPLsrdwDP8ZMfA4m/bZ2oLOUtdJs67S9p1kYHJEL5rRlcOzqujlA2Jp1KmV3UrMm
4b3j4pD3Bok+FBOTYU5I+UyV9Shuax5q0Qs/XVftkg45+98YS4wbA8lrZ5lGp/LN
v9L5sPxBWSDQgo7JQ4liIGkXe5Rv7lSfVAZEuP/XOK8np/oWZVkKhc1k4aPO7Pgx
Eco+Zpg2jaOWixT0jf8AX0SIXWwYBNxok0eZGo77aKV63/PGqJqzWfZJQCIqDAPl
PCcYgEV4ku/Z61JJQqmJDSdakLXkLgX4bnwV1rWTBADQMMkI4zQRWnkeCsUT0enF
mr4vo59Bd6UdButB6KtCUBKXaM9Ewb1bOOeJOt9qFz/MutEPWlSICv8uNuTHmGiH
H7Xdo/Er9/ZxwN1AD+kdqGfhFXkB2JgGD7mi4sl6/wFWPH7TjRhsLmzpZzDMiQ66
GCoxACwo3LDLvtp9vLH26YaveAKBmR+JCtDlJ6izVB3prSkcAlSlQA3M+T6QS5sv
EOPLP57XF2ndXX0TBsrYL1yP2Wst4SGwOEXdtp4JvqTTM9Ms1vwzSUlDZRo8nbTA
MzKaeeLu+DsPqXaWLdvnWpJQk/zwV2AqmFGuQf40oZvE6BMP07OjKBWHNSgxC6fg
XsUPwD0SjVFDsxaSzN7OEN17k82vHQkCa4oQVWTJZWRz+XQzyqt/b5puMwxp288Y
2tEDjddIv6sj8XHI4Y7MfWSLEzk3CX6u/8NQFr6mw4P1UedaO+i5iMF4U7PC9w+G
l37owi+UH5c4OcSGqCMhvAyK5mjIWmiXKpwUDqPoQCkMjCHEKTAJu8xMff91fLO8
WE0P7xrpVWijly0yQS+MJ/6B0DeDWNydoeduBW/rm+DXyStcUTvGjoul6njQzAiW
EcYlLmLKVvxvTG9ghclorrNfmFDgyTB+3WDm2PK52jam3J76wnepHocD4kQQ2jM5
6JhK7R0f24HIAd2RTf4B8LmiXI8kr4Xj7lwWxPqJfLATfANEUuGFGOV2ZGgzW8+a
Xy6rGgE7UxP2IZZE8zKNU1nyT1DseIDaZ5XijK1LwL1rmSwJ/KU+T5o6JcHbGTNq
8d43x5E77em7VkkpLepNjQeREnMC2G9cWCPlM/n1B/3UveHgrVTE+bukvWa5hXge
u13RHENqa07PISdjfMOguIuJzKRyi+b6eNCY2BeokNa+CRbFftUCGTMjZVTF2Jb6
6KOhwEZiZAK4k4EEtTbSTOgE3Q/TOPzaeG8XXA/qsyB88kv2fs1lJxePpnvMA0Y0
YBBqTyUmPyEKkilAe+Fy04efCM6AvKD5WDkDhwRUqke6WkMHvrpwXq8y4gKhlkhm
ZeSKOYs3W2mmLAqmy1vlQpqydAtf1TYakebWlEjmolMOAm+78bfLOwPqVuOD2SU0
GBMF7f2S0NzQUHSA5+BEWTv/moznvbJ4Hu5WLWDX0mMsd3xloiZ07igKt4COg04j
3VCK2yqLRmxMipKdb/v6kiGOdhHWw2Wt2xoxEAKp7Zq7FpiX0J/kNtk30HLZGhK8
u2kUCcyb/DW5e2knPGlYkFwcEbgsGocsuYAHCoCmY9wDtW4o3pzyG6KlCHGxOl0u
by8HAoR01j2Vl9S5IpodMLO/+DphJE/u5YCDTHCR3YyNNgjW/fefdtrF5wNjvbOd
Hge0gH5xyGSbB4V8KmLyobIZbTnknen4r/rK/On6mHn3jXOK3vJdhauo/pxZ9pes
sq/oyk4S9tFFyXuqmvY46GENCchqTi1uZE76z6svWOtlEQvadrjNv2YS+TSqKlra
9MgIu6EZNFQ0571flOaMbbyktcTt/LyXXxtsNQf2SVjzxck7CSD+UvZD+Hlog6x1
Orc78gESuToMR8gYVEf2ccd/3xzDDomIFE6hYqcfuUSpVjKDYJTumS0dStFLPM9B
GwIE53DGwdEY0+rXNZk/Z29HP7MneKbrS240arKT+T/3Y4E8/Dp4DcNwGCsqxZRM
DF8HunPT0Dh0YeEEZVT5Nlct07+YNHmiaTvHuLKmIU8a4yXGltGrvV+WwUCrRsCX
UmwXUS6bHGORXp4+npZF3wpQqKcKE+YGpru3YINImDUwNA7txTq84cl2RI4WXLDo
9s5CnfJRpx9I5m/6WUjAW/7HtJe5QwBhydlt/acMboTilyf6Rr22Cz6TrYpcrHHh
eCD4LUL2q1Y+NnxvVBT9AKsEgvkZGZKXJyAbefjMQP6vBy0dgu+Ubkjyw6Xma/69
mA0wsVo5awslQGauFxPdSxV16gZICSxTQRcYbEC+uFylRHllyuyw/zP6mFx8Ethk
wAScH4Ip0di/teSWVyJi4jQp/iv3NJo+ZiSjfzG5aQXvJrEBgkeiA3T8WFmibysF
tEfFUUOxYXYNmFVIn26D0fJirZBaxtrJYCCjNgXomZ0c7Xm6jI3PBm9iBXNHXLt7
AB2B5lNw2qudHnQ6xMb47JS8kFpWEFiYnSEoTI9l9OfvlFmc4y/cksU5+upwpyH5
d4z6abRU1AmFV5I/jpZMSWersYgAwXhaWpiHFFsGC7SE0r78MoFBrewxFNRPg8aT
Zr7UknEN/whSUp42cPr+J60UeBHxx4cdjAdssegluRPwW637w0c9Q25aw3/sRYHD
JvkJPeyAXSbwA2Wie5zx/fuvYQnqXrqKZ3elRoWHu/zs0JxrdBcol2pc3Dse/YSy
Vh5R5svHiuchRURlDda5CQ3DcI/hkeaglKiqTP9usbskt39c0pf+tV9XQubreUSs
cq7o7zvb1VJgL214hWqQQfabd7bXLLvWi5pjJhzZq8VdVEjlYl+XWBznwR1mugpm
AtGpwVnRgvr06wyXMfT1Ekz8cCpL3NnRCf7OowG14hnycTaYu48lnayCfhH/ih+4
dk9Z8c5R174rO3BSLD69pfHaAvVMzyJUidqVDFnYzbZqLWqWR95aFLjYz/PDgPux
qEyMEAhBGwoKOtHk3DIzTom5ylYs0TnQOg/QhRM/ROyzXpdYI8Q/dSToWq4pRnt7
R9L+O/2UOSgSll9Y5ETUSzyTjOn2MUulqf2QZeYWhNys+60+a4FnVnIRYKNOZQrW
XrePlwZeoHSIQtVvp4XGg+MIK4FOkC5vQeIZ/E6szFHJwGz+oxNbtS+XauGe87DC
T0tzMLEZe8MjttVR0dIBjZstuqzwZQHzmVkM9JRuhBG3770cNn186kGVKMwTR9Cj
y53uZpNrG20nmFlYPM/+VGp/rvhTXwfMxuMwZ6dDcp9sP9RBBxkcFS180SJ9nCol
vBe1nm9HofDYxEE5W+SOaW9rymnsBzJFoMPJ0le4yW5qMfCujQunAmJ72q4vwdlY
dDRl/BjbMdZ/QoAmSTdi5kJRsdjLJO/+fJ3M+c6qKlulA5ulukQYodtVASSknzeA
Ui/A4dttRXJidQVYtMd7U2dOaHv1zsbSdGWBtFeteQOq/0jqkwhsCmhsdwvRY/fM
8COWFBv5GjG+3F8E14xYGFKAzDHfDYemieihoAbNGDr5ViaA1xglwYrW8iF8RpA5
5OfYbrOylCyEHQpOwDz/mVxmMTqc8gykbBo4RU747I1+ASdgBowwhtGf8mz3fm80
+bLdifNNRiDGKz8O9rglSUyM2fSmiyDUFsZoYoCBQMvsjsBLqqgOPznj8YV9meZZ
QfkhDjCoKTqfNxwx6LI/gcIRhp8hkw6STXAn6oiJcmZzANYIxjQEdWc+2gWwuIF2
K1ogKZfvgpJAG7M8CubeHItN7PJ0slqbswmYjibdTeeoUy0s+gVNA6V5Ra4Q8ZxI
kGARJpwIZ4YzvWKfMkrVZMZjTR9wfAqdTugvijnpj4jkrIf1bbSsBqboGBc0AcS0
y7Jqjo09v9qJtuEggyOsGNTgzR5IjfVmAew5lNbVRbJ5xOnUD6jc4doczSTME8Hp
21sTYlEAz6wRvcFtguB48rk6+3P3+tTEDCJvSDGUXNkQVuiHkl5POlUeZi7OvaqI
9tsgkheW+a8mJSo7dLmxJjhcl/aV2Ay5hzEz0E3mK8YGv22eOVCqtQo0cra6Z/tg
edjYyVAMhDhmGDdpce8USGSCjx5lZyXMrlMDR2fH7D/J3AY8WO9ypEtgtIBm1bRK
lqJan9IDAfmOUN0+SIOc/lPCjgJ28I8n2dMmbMMy+R5++r30luNj7984qA8nO14k
UGPIvvQD1R8z2ZgsSuSbuBj2HyqKTYhyRFLfu3Msu+aS92xN5XfGb+7YiGk1YmjK
QOmPGENbj8vF7D6UkYLVbCx6Y1DMCyD5DzIzee9MXJKvu7U5wmNkRZ4PPuNHmArz
e7BCC/EZUWYvjBQyIByqnvcGDi1mq20kSd0ho0LYgMQeoWUyV3g9RqZyQQrJpGD2
YahuAiiS8fcsZ3gE4xtsydb89fGFLv2pkd203EQbXEtSd0x5qhcldD6aGeIgmg7n
BLxIxjFhIV7kARxmNdV6btzrr8pK6LYrj4w7pxdLloUO405ACsqeZqOmh7Q29Rwj
BJuiB/uBfkKgOTVslcZPaaE422z+LKM4a38rrQl+wN2US7pfrvP8DVC76Vo7DTfR
nsS03rTowvOVSWf/W7NQ9fVUlws5g+XplmcY68E4FRgpKkNGUbPg+wUieYa9fmjG
1D0mqTfqGifOzH4vpESTJFaowFTbhvkB3FTIUHknN+DuG8Sl3p/ZIjIMVkcwER0A
XbV3YvvF16j2dTnnz82k35gPtXRGB1J71JAuqljVE4Fu1GMlHzkJsLJzaaDRy/Gn
POYz+Ab8M+6cosznLnJvo/NTQ+AtJoU1nj4of6tz7TILuynqV7KNzcs+jCTuLGzi
rxTir7lPJ/QIu/Iap8i3XzUpmjECdOpVvVlkg0vXaQ2J+3x7kHXOEuWp3hllmAWf
JFPQX368OCZQCwIzwV5afBLOOFOjFWPCuS8TDAF6tz+7tDZZeGU65HDaI5BbV59u
bW2RphljVX8RT4LFLx7H0fQyv1fjJCTpFJOJbSJKuwNj2PFT31Ycidef0YfgJyA9
e9yIFwnskYnVxRYI+c+zJy3kffqFnhEwbHR9rk1esU1H2NC80YDXuTME2+H5dN/H
fq84DVEQC3aHgoTPABDThGhzgJARtxzD8EiaBkHbTXVW7azAXX6lL0w7uhufRjvb
LE/6Ocvcz+Oqxj+b52DgnR75Cq4WclTsCvP47aLJ8s9avksH3zvpwaiEpjOTVe33
YOnUF1a/kzY3iPsJzdIHbnuC2LMqvrsDJzQnQmf/A7AEOQd9CzTL0ZSGfernPZxH
DwHvxWB31lHwXQ5wmbjPVzXgFdKaEf0wCUn+dCfB3bb+/I7rojH7YdtWoK8bza33
hnDIECRkMtqF2NKd51eOtKIK54blE2N/BzSFz4uKw+P1UVyqPEascn+CgtmajX9g
/uErifcl+8RsvVTFeqqQhXFW9NQUiQgz8AXgXWvY5ESdZ8ZiWER2H0JIymwc2UmU
Xug5XIcHQUJctP/bolsBtLfAtUKryYQAYki354+Vn6rS0SzYqIVXLcPmW9hudcRv
oA+NjRpOkrRHOs1yxCTcUd1cihySVReRhKIBeVvg1Zqj8rA8RXb58fo3H6nMr0VP
oxMjebeFaHhTyX3hBrDeuypECBnuRs5kzNMEPu4c1WQXFE6GZNGxfnHD7MlpLIZV
cP8tcOIxmhu40sWKZsQHtmeUl1BPAov+HT9Dne6YxjV9qwr8rVcE9+uMglQuNB7u
JC+2my68GNprLEWeWp6kdwDrOIiJcN5L7Ly/a2SorYM926zmfMX+2pmYqs9OUFPD
6qmWRcHjBT1hzFhncbEhFh/oc/E6PjaX22z2/w80OKkMB2nhR+htcrSztTgXEPl4
CcWKkM5Jyh3IbGx/DosXwSKELl09TrrNXFmFEzXRHSgqDCQ9grCU7eHmug7OVNNN
2FPJW343QfeoYYy3dJq8dJz9O/dXi2S2e3NNe4+xYgmmg8/uOOrS3kZA+sGz+w94
1XmO2PDoRe+dxngdW9Hb8sjXTqFNOPEIubOema5Zduyf4C/xsZqg+TQVQl3EX8m/
s+FMC6BpXfOmLLi0Ohj1Sinfk/HCLPOlJWui+Hw1N7Jhqwgv34/rwAs0ElJQlulh
FPOTLvz6xWfvF4C34SdRbV2janBNDJPw/0qjRnNEGFdlt9a7mhX2FUgrAyerivMu
7nPenIzDCc3u3m+CsuRBeQJz9PsTWMgWwaZn7xMLKTPQITW+NsT0s9Qeb4jDxI4A
okaajM5bLSQxgIjJ90Grr1z6RxUEIl1+3TK+b34TwbVtJbZT6ywcBwJhB/9is4n4
0jQuICHXBMr+50qgsNbKoX8kNQaotzvmOdhpw0vOgI/qDx51YZyKLN9q9CiH2C2S
6WSd/yBgvKXcFsF/N4dAICK74WluWRU4lfim1JBTCul8bWC/xWU7Hg20ormtXt3o
lk/yIaeCp/UezndqAwQO8CmBWcnnAv99Sv38XE3oVY3P9gFlTDhy+jNNCmifLWwx
zZZ0/TwDIfI+4jFsEIpvzpvxXQi35OKECGWe9hOZQiF0B3L1SwdRBfYbodEWRELb
AIaD+jmBrAY2A1B3GigGw6u3qse8SEoqx79u1VURf5NXsu9KQ6TQWTiTHY8KViav
a5XHGQLx/YD9YJRJO+1MJ8qyXgw1qYPoXktlE3Qry3BmrxPLyvWxu+PQM8om0+jf
R0XjOaVb27dUBk6NcIIiqFiIY024U9JFjJLUPxF6z7liCQ+zANmU1ZzBZXdLoznV
Aw2lom9QZtkSO/yOfDA4/vsF9kD2kGWQDVRyjAYxCq4QAvKBCVahYl3TwVyD43k7
QPidQDM0LN/LwcqlVEmGxThH+uQUXio8j+auyox79m+D3O2qmqDp220JQq1MYDCq
ia4rydVRq/xs5Dnq1TWyOx4nzdxjMWEdRV1fY3FzihcDSmh933SBDIT0YScugke2
tiaIEXh7v0vrPYCQiLtRcxgi8vZ3xHHViEYfMT9v1kr7ryH11p5dJkWO7jypmAQL
R9xedOsKTD0xwkw8PW+Ef6mhnYA03Lee444oJL8KKf2XdHbnQ60N1GXbeds28l93
tdItfq9GtbbEJf77s8i6uPAX0yU3miAOMtuDgBjad0/fLxzFyhwZsJCXmlmENqSQ
3qiqMKFbAKeopRwDUEXpFwO22trWX1Q7x91oSuVvib+Nf6cKRaEt76kPisZPJwx3
8l2nXlJRXQ7VADyLIhVhTSOblbiF6uRoUn5PyvkU2pgaDpczUMNxtTubGzCHscJe
XCzlFdew6quY/Txc52cdXGvDAjEBOBo8jn+P2A4DYSXIVTMbv6YU95AMuhMgWgZs
Y0vAPuyhlrKwQMwUbGH2Coz/Cfj62qFASsL79oJni6mSCLXa7hfJkTtW1VoSPzAj
W6FrKAS1csOjd5I+4vs98dk+j8piIU1kTmJ9YuhiTtcIShhndmVf40z1TlfaK4C7
NEu8o5rWOm4hhThHJpLGBuC69OaD4OUcTdWs8HhdGU+xbi9x8oA/pMCy9AXBFwRx
sVwEFTUv+z1jD0BqrXj16pQdGZAl88oONcFIXE9v12tnjjfxSSQeb/reCY5NJGFq
YijXAe+vCyoO0+qLxCq0gYgNs9BqDVtPOtRwlZ3v9jgdTydphHW5xOVxIR/eyQY8
jve/Y+szaX5MJFBnUI8EcsfAkTsray8LiLEv3jGjE6390pgGcD4U+ppAzp+GZZM1
qK7QsZHQXOv+XzDbXEbfnxH9j79JyCw4I4iArF/6nRvOL0nEKZ36gEvDCTgxRbNR
IU5nTfOQpMwEhyWerBVc7hYvO5OnRUUj0hyBRgjr1R6Vno0PwaGtlywwSPJTfIwE
2E9F5loTiEgcvPdHoHQJrSnoFsIiCem01j2NqJJYZ+Oo3ohTiASYy84Nc1A3yNlB
8wHJBy70QGjmOZ6crdkM4UFSFvrr1esM+XuJpGAfJ/Fa0oGdbEwYTGW5OWG89yAi
pl38ryv13ZleEoWks+0JgDYPiYEUZc3gVmxN+AR9nkZxZzhbmA/qn8/oD4huuS+V
U1KhD3BhlLYAzCChb4y4q6xkWByamsZC7OUv7Kv9J2mSKJUhwpZToYK6vIlPzYTI
mEMzwimaLAbs6+8DFYgz1a7hHnJKCZgTdcg0TVWUt9PXrsLnCn4eou9E0bb6+toj
zw4TpBVG6OZRUSqVmT8u4Or3rf9YcKlo3tqV3HISpEQInC5gVnTDc2qu1YXenLoo
iziGA9ItMIgoEvfzHqIQn8P6t2Q12cfwI6Gm64Qtcits2D6d6sM+2ZiLPft1gmf6
MLg5/OPNSEoEc2eIUk0fCN+A9bngIMmsOAHeAZnC4pgSCbdmbWlR8+kIXYviFBmi
u9oXXKnLeWs63/5BBNeNif+gCFU0wmVWzq0MEZ0/EX9v9wuB8Hn/wDhwS4uYfF2f
+sg10oOMsSfp24d9dlgfpxUg2cL/kxmzfivAITL4xDSlfK5Q260QnXl5SR78cXh7
+2AG0ySaGrBuyLVWndOHps94zm2ZG1pnXAJqrEBsUP9Hrts0ZXm1/7ieVmCZJQ+G
Wpg9tcH8yTu/1L1YAqsIXg7Btq9tTUXs4dJgh0CFPf6Jo0BzyEAG5EedhdZq/mVx
sS8CBFmwJQfuCdhU/HopUjFKkKCW29xvaoBw+V2SoLV3BehWM9mSeeLRIQmsGt3T
4K6njTOMfu7ZZqa2bXoJ0ElMGphg9W54xvChUHnvZcM9BHkGG+rq8fTpLH6rDgxN
KDZZJ3uvG1mWZj+wa0PEHVTID3TlzjdkXgjolgJfLpNBtdrIaD9xEIm9WcxxgDjb
MB0hnCglSdy94BSw7qj105YDtxbNRlnvHzRKPlSReYWNVv3RWN06P9mVXbiNovn8
+Kz2uj56s3n1T2EMiL6b1M3G4P3S+zKIsvjRzd4ekmVMTxDkkjCPnGXzER5jwuKM
2RlKqHxgWgd238vIoMCQ7LcyiUEB0mf8gZVj71C0hfWCdNOGV85vw33VjFaWoVzq
/GLzYhpEpTIGQPUMnz+mbaZC6YXWpPgIPmxe6zWPOgUPjLaXbNcllBEb2/h/Jp2j
5F7aVK+UgP1GWW/DrPHPZTCwR+eOjwioV87hFVck0GVQiPRI+0iW3PPDJ0QySnVX
kGCeHONo9VI6qaCLLbcZicjxHw3uO63hJPFJIgJHG3nFcsTCvcwELieDFgGdRhqq
H1i4ghRCHxgNEaU4V3MaRc+Sc4Crs2RGNf+dSLUSc7T2p0KztJgJBtSJkmFaaDGR
SLmifkyksMAv5urxqxmVeEZKK74XLubZpCQr+AevN5JVDNUDAFbIBvSQITdy5b+e
QUywS6PuG4TiN4uTrWkn6yimCGnylhZvh5g5JBqtLMsmdb71BNLSkfcIpvIiV4Yu
ZD0AWAyo17kql1Q/9itVNcTLbY5LKs/L4794I6t+zXoXmsLQ2UxeE9JNwk5y4zdi
FVng58MNH4SuUlm1qEvWMOH55FXe5p0jar0JX4uKfSHU9SRajaa6Jh0eLspNWw1Z
umEF/4QWQJO2slAT4ULHDlmsNTXY/1XjwZVDrI2PhdI1/6H3f4LGnK0jEPCDVByO
cmO5hPETc41XLewKCTySn3oaqpZej03eWN6rSyIlnce5svSkGyp6DNlHso8xS9/2
Y/gwJ5ZEn+7bwiQ5re+HnV4VS9dV4B4RDDCW4nEl9naX/jCkL5cfJY18V0anszXF
AppaJksvfLhPwdOqXBSgV19CtiOWG0YT6/eU4YnnCF84me5rnZoyNQ3a67Zl6Viu
yr+Rkse/TXYwsy6RoS5I3oo65ZeJf+rb+GGBYeB2goeQ2sXxIwx9QPkrp0pKE1oe
+aQ0v3wtIictgtJC8aNwZ0pqWsX5TPdxRZRjvMNyIYPYy2Rkq2AwJTV+taCA+1i3
d3m/CEE6XjfG8wlH3AOx6tzHwoHgUb7/V7PCv9E2ddoMyZeZSvpMqTOcXK/7FZ0P
bDonVvbrtPnjFl3eN4MqH2OI7DqcVjBiz90xxA3KSQq4xchWCsMJauNTfg6ANGh9
mnHcAy/tpyMu3uzth0e6Ub+rwj7noiOeyJnhKPofVKCrMbRYnkaPaaMtj+mQ8QEe
Dm6zf8TLFxpRNAXIoodybhjsRKFujyp76Smqeq2YBgCaWp7+m7Ja6jQUvGkERPQU
MuQ+Z73OEDBKsJ61DTEB13MGxR9ugmVCQo1yOLmy5rcJ894kFI50A5GXstCjZk1b
tRjwuCtXY2rBL95j2WgcThSNtw4jHxnAG5H1JbNQL+Vp0He8S3S6NIh0QONvAiDu
ce/pbsmFqqxWZvBmBtUj1+sZHYqMvwwMihcaPE8y4W9X01FBTo+MdfNMbyB3d7Ie
Nzrvt1zWM1SI0265QQWiRCGnfRPUM46fO8xpsKwdsP5862m0YWiCLPmiQxDC+LA2
/7UbHjOLq5o+gBrJYhmWplh1Q8mQscutUl/bmtGXQPNN4u9ouGTkMvDlkgiLYZDO
m7uTidPxHpPCU/EOon+apO1IK7vA6Hh02TqmW0EduNk0RLkkUcszdGfwJya+POdr
w/uWRtrbGugP+wnetplDoZA63j9jZXaDifgYDtISSeEXibVPXGXP6wpaV7Edjeud
TxvMlo4ONruMPpH1G3Ifjv5pjC7btGpAktPpLNaQzGyJRAa+monCYNKpUuxDyvad
cBL5C2a4Yz/i9U7P2X3KNOsYvviMUv7Fgp6T/daN/0dX4N+lfymgGFMIV7cv9RYs
W1yasrJxWSbLbFS2auuFCoXQkPTUfQbly3skj46px4Bg1WHjpzMPLoNN6E7uEE5Q
plKCbcUnQ+GUCZ8XoURIhGSfoob1W8q5zlMedLJB8sag9RMwdvgdQis6Pafbwfhp
703cwqug8174mkTrx4uMlVMY2pp6eV9lsdPCrLIOHj54DaGMt8fs0C9rC3z1gqxP
X5yyS3hhs7+lPfq4K1IJOSr/KUDAWz9eRHwd9qvdjSRjZLOSqKnUtARgj7uHCWVP
JndgC1JldSFz0agqT/cBhsvtCTxamawF/6YDMnDBHFe5QEC3LtlryL/tUUEDIxIs
iWdf4ceYF+YfZb/VfMkFUOA+dlc/tF3nOz2xS15c5rmRzLxr4esEZ5thieQ0dzTo
W5FBqEzHUDk3sqNQSbz3aaFn1lsklEBjvUxHCjUyZLocpTZqoVKE/zRtXXfxhZYX
mq6l4t5QZQnA7GwWfU0p0FNG8UCPLUWCwInyd/roAawjSOGFuBP3f6QNxd5LH4BJ
+DC0xlcI667/NW8N7T02inb2adMl9iWjYUZhQJUVktvhZhkUHwAU5b+QXRbtWgEi
IPA10RlZf+05bOHhURFyElNu0pOTHG47wJtSDC1NpZDuGCawkgqa/w1mQ1Y+ubVg
tYNp29gBlZXBJUh/HepAxA7YbCcMtN+e6u2BLb7jCtqvTSguAol/dZZdfBnAovdZ
HV0Zg/SeMZJKsIsr10TPrt05FM8uB3+2iTEqmoiW3Y8pff5ZwhrYRL3fQAeGh9LW
MI9K1i5UevhQV7Tj6PxFX1rLwM7W9i+zuY2YyfXYm0M0c/zklBaGMcHRnDaLxEpY
F3Krj5rY0+nJkdSNBDgOzwYF1BKWL4SkDifS56dLcRLzrX0EYBaxjvnS7aGNjS7l
yOcj8RYfZBlS9Pmgko1w5SiR3LkbJPOQuiXy279UqX11YRwKW04CyI3mYIR1wc54
IBJTOXWTzP+5VNod3LQF5l9oaxjW2DDWuiON37qAC6PXgFmHQEZG7yrWBdsOxzz1
12fsueIdVDEa8s9s9bO5rNQDIt+2ZuPoW6egZD/7nhgCmiXSvRsQMA6ADCnj6OL6
ezQQ0AJwsA/fpTImhJZSZquSSFKK5XgQzZcfOqUuvbxAl8+8UcMcrngTr2a1Ci88
Ey/xfAhyM6n5SSANvLF5pCI7OmJa1xOR8sQsVrMUsjG+7WO2qL47Kpqn1ONV9vuw
AvaFZhMpJS9JcUOi7876z/4Tl1ugaFrdHOy34OF5T5Gs3QiHPjdv+JWplhRBumll
JGOzO43ghRuaRdFYRyIil7llnrJ7uV7GsdFPOyzn5KoSahyEG5BbQCMleUg1cI0J
8AXy0CXT52RBG/7WqVKDFxSG9AJ0/eR9rC2zYR4SH2kjaSeXnzcuyZ19akvizmPe
Npv6eFMqhn/ioPdTaUeBaFijxY3ltZiH3eQASKRb4QaucBpoYeTDn8OWjrsAQg62
/InmRj2IF0FrQ+1BYEciKo2vnNMkhPNomoX/j1awp0Fs13We6PKfqrOSr0lP/7Qs
8QZige+E3qWgkPLntEhAduE5/KBW1VURi7UYR9qMq9sagpOn29U5SF5iAIUB9/JH
Nrse8m7emeuKM6w2KJ9HBYpcREeUX9VZaEgeVRG6Q49aHNYI8HexXaG4C1CIHydf
SSSIe0kP7JK4AI2FKb1Rm3b3EPY6F1c9P60ZNsPxCWpqsgtOWZrjq7kX2Y4zCEwJ
FvyqHLHl2YTnwnfFMkEtBeB7pn3DQkRcnLOeFzqfsmjhLRI+uRziuEf+0DxEx195
3JuEZ+eVn6rtBuSx5xDgOTIvoYkVMElJ4Zfl3TURwFSC66ARYcw5f+4EsVQxjNKq
BaIOLFP02AQrzx6gJtFBcJu22NPGJmrVDxrT5jjK274Kz9JaxhWx7s4hJ0dpISnV
OLVokK6+m+1zuPB+99qQ/7DwIJ+tDL+orj4htvbep3pLlM7gpMhZf6CCmWdQeaEX
YNpHr7NOl8WJ/muPtT0hTvrACRY2xmXUOqjTaQzvPpkkxGTZHQpw5zfZ7zfUTiyn
P9Sleq2tWVpixThcn5sVouvTlIir/Thj9Dmq6fkYbwTqcRRRzb6n851x44y+DW3A
PRi7sfuNU6EcHet0DBLIFPrUWF1pDc/RgzrQfOJzeWsD4oHHYVcVKTppT2pYFSLB
09nqs2taSNHphxCfJiPlNycGtY/ZjPjIUOCw563jF4igEqepwuMlh8Z+tZhy88U7
/+Mk4dC5Nmb0wpTASgW5r4m8ZkJkIrQ5DnHjEcjFfTRavVfGN74e2KMSCe8w0Bm5
XP8DU25G/FkMsSWpfRN/2RR5c3/icTT1Uvan8hViePkm0ixTM867Qlv/fI22Wk+T
QrTeJyoUwrKdvcUXS57eheB0dUkxwpwO1m3iv/Ihyufoppn2JSb6kn9Er0UvCFyA
iz/B2lHtRWkKqVO7d0epV98kCbgYOdffJKQo3Q4FfZ7I8lZh6F4vHRUblZDz7U1w
eayV+GBVYdj3K6nLyukokbWv4Bguev3NXeB7amNLRbvSG7oJ3cDL3aCZLBcewILg
Ol785+2uqEoZfqK7li8jjiExcpBhvwkdxxmTgimQsFSNdDeOVA1zmTRWD3BBGT32
py9OaxO2bnMQqBfhdCf5Hbi+oT6mabtS6QYDRL13LMa7jjZB/TVgcenp3xmweVdL
zljBHLAshi4kg6UrWgTCGmbCKIuNRBgJkVqXxB5T/wVWQaQQzDBta+Zr+Db2QfKT
TdsnxU65+sky07pPtiKEQ6a3mPQDXZ00fGMkWSWJFgv7WI/EO802JA0Q9pnvn1Hm
vAfpNnhkp/uGVSp23OWSsxJ5Y4zyiUk73yeIXj1UggZfc51KJDocWCwTyA0YMM/r
8sdJgN5Oy0faGgpVCQq4Q5sZ+g+g9teUY8/Qd75mbWDCUaaQDO6i76UvDbkKu4s8
39rHn7bhFZyYyzI9pGJEEMI9x+2A+kt0B5IMZdTRbwra3jEL1Gw5Z/z5TqGRCQlv
uLNd3/Xj0Zq1x+hZalJC0YPUNYf/W8iHTi3StI8A2zoT/YwaUX2mWRGEAJYkOTbd
ts5kSX3His4x9MP3BYPtlmxxDnG7bi7WVcU4ZLEVx/uaQYBLZK+uUSgfsco3wnkh
YyqRkz/wZfsGl8k/Nwkq/QZRIIw1UPSf8QkNbrxSI4szLI0WrXYcb5a6HqL0zOG2
48fbF2fi611j/HXR+pcORO30ZIRVaBMggckC3LhNByKXjLRAoQ40zJqDRpr+Q6l2
Pht2OwCyuC8BCRijCRp3/TNTly2pHmsQzjpWog+rN7lS68NtaDezwG0xxacClo9s
4EplEBkt+nO/chBf40XNZok79vB+Wq4CDx0MXI1NG/+pLbXNZJgkBFKIWBuKPOau
dC/1oRvulUGSMQsRXMWsO9OZM2910UI1lVpufhyKxMUygv0zsFXjzm2hocVaMEef
ACM4KNbdZMEVMAIzJ6wswezeFZXKtNUCdLsSS06+MdN/TfdYFwoVI9BFnwx+C/t/
uyAwQwn+KF8qrd0mjh9JBc3avQHDFedai3wfs54ehYHFR22lpw65luIMUEQtpOON
OYRC2zhJUHtidSgM8Akm/aJdJbTzSe0v+vVfngqiOgVgMnWlB9d1tKgL9HZJnrKm
+EcL9rzKPTsZ+fV6BLR6WjPNXlX7HmSBhKG48pDt+tHCEt3pJSvwQEjsy61dBybv
BU/4DKGyBLrlt7DpSMK9D/ZtSw2XnW0q5fmHJIpYqY86GF1q6dwsypPKuUuVf/oL
c3Ef+9wCEEXY+8+UkC9FAAzXTlmpr3eUhsY1Jk0yjxUFUIftmRHAN6jzllWrpCrp
QjN9vwJ3Ycf41LL8AJLr3IzL5FVQJJUv2VUXx//3Ms7kw7pA9uq75kzEZq7KHa8o
0EemR8enuvNUbT9lvl26CxO5qzWY3ZVwxFIxMhEujx9lA/CeEjYsn5YaVhMmn4Q2
Qt5tifMETY0tuyJj+JLDgQ8mIm2ME2e50Nk40ecmVsgc5bP4VYWyjyDP6mP1EkV5
ABZZcZq2fbzsF9ttyGX/M+/9tgQkE6t3PcFRUhPhw/xg5r5nYr8NmhxpT4FrzhFh
BScmntx3La0klvaAmT/HWcr6I0i5mieIyUdXdoAgrOCbPQPrbwqPRqzeA6i2NcqT
C1AIqp2DYf43TkjvFuje3L+W4y/7UnzyubxHen1A5MDENxI3QBLHykehQf1fP2NT
sgR+Xz1KobEDwBoKde70aCXXmRKpYSHk9Rllb9op42gCBZ7ZyNW11LIQ23pzkscw
s+Yds5uH5zLf13QHXorRIZwmALKPS2YB+BhjPcFHYcLgZky97ywHEHMwJ3AWiu4k
54HUb/cts+slEUABhZfzv/W3S+JMJABNk20XJh0Iwjj6dYjhK//y5nhpU7mohCWF
o7t9E7TbZiD39YpJ17P0PS3lHEm4xOdSH61kOIMoSZW72f6sNl4etm9LPOSdt3kK
nH/U6CqDf3zBIAWMR/Iwb+hsV8Sw8nH83xBQQeP6NiS8IDP0zt+RLuHjxnoQjx2L
9weHghmkzRQOYEBKccnrawc8YVeKTh+vQP70uZZqmAaIMGGpTDit8nxd/1mgDz66
T+yahXIhNgoMWZ70zHzBrw78Osc68l9XD8sm2RfrHd4jkIrgrQQX1TtqjTj5mD3F
s9qZYpNQkX3p1ivHXhs+CNIDwTzp4YZX8pq+SL+tRjIFgcVejtoCuuA4vw/2MGLE
dnW9hf4F9Ypu9mAgogyjEwqcJGjvblnvsMlcw2KQEtzLemLMH5aabU0LFSeMtLLh
vQdngVlRJGzFpnW7NOxRdrQmJ93btN0lP/BomGNULApI4zwtVAV0MTC9GOFYyWF/
rDyDu4EtVcySM6o/dhHuLNJyj6WkC9YTeWwo92QSByLbTIQA7OUGvpm+dj6vO9/7
WtrBHVyOSrEzzPjcfXvryOzF9JO2vmp1CwzztqHTnZiKxioXrN1QpOTROtMRPAHT
0NtR/MoJBMp4CH5fx/KoZ/TrNpw6jph+kJKBeEDcfOo5KEE6Wyg24T+8R/i1dz6x
nJGMeUdvtJJSXUGru9rGijVjzV2vCwpQv/DbrV4CK/SZ6eacqg6ObELNSAbYqL9J
WHPmLFFsDl6Xlre1GlWLpdBvMdsp0ExD6vNrec9ys8bqL5Y10Sj/8vpYqxELcNOk
i1wqYDLdv3/xbhGKGuvByBTul6ZYwVAyJxYe7yh0PxTeNSCW8CtDmtwj8RPULTTb
ijkQzyNcomfn3Sp8faL8xRQJgi09DJua4AIg/kheTsrff6AoN4pPMyz1uLRvP0FD
JFsMB9Ay2VIz3xeHnKpeczMu2Hs+TNUg+0QTNHNzMJHrrPT2D+nEhl7FwK/e+R43
d8hXilPpfFsbcVFKBARilCvOr/oynWVcCdHZ+VpcA2yiGPPZimGQKlLqXkMySkWW
4otso4DT7JsMmgkeN31PTfHgIGw7CIEYI5HYvQW3v4y6AbdUV1I+SHqZL5WqjiFi
zZaV+XJssi+7I3JpilNh5+GdfMKaYwWM592IBnaNGlSKWNrIYpHS//4YenWdQGWB
1IhWLcGXxFbDgpwsykQcLmOMUaOlJrC+tVA57Chc2c/lh3652qZDA7pXNHjj3d/j
akl1DGkITG+ZQdyzXmF3QbWSQ47K8StuGEbOoOM/gUA5TliKsnrIAYJ0mtksKgjV
5k9jXUxKIdZm5JCy1dWaJ+9SYKKDCkNbINpOjOCF2syhPyLYXmVuaMDPltCx/hNW
4jnuCQlUK68KsBCB9ZF1ONQSYm23z7Hdaj83PlNL+E2+8gHK09lp9tMEQEreR3Ub
GzWEPHKqhH5zICVnP4IYBENLuiDk0paumAU9wYj9Jq4z2jZc4QkYMupy4j5z43DO
kABBd/UP1TP/zIpX6Hkw3uxXCoTL79fvJwvaTwGkqVpOh7kGb1Leu4QHaZq1+Yv9
I+OkLvsjQdfhlWzJ9Wb290zoEV5UWqcF1+73zrMiroYHiQqTlw27MF8S+PBQIL0L
TOtgqDN0CkUABy0xVLTC2YHMxGD5EQrfZCRASgzpwF8MhoHvedIc/UWqx6Ccmxfw
fO6nHG5ZSBS+sHXx/OfZlc3w+7Z0f/69V0bro5vF9j+C9nXFjRmxQffw+Pb/BxZN
S3ceitUK0YyLeONFHgyfgFIkd7aCm1yDMw9/6MP0l7b13YWYVEVfvKIHqeMv0XM/
5MXYXWkZNbSlKEngXN3F0TRl+qAMVkWeNkC+AIWsUqaVzCmsuN1hcdRC05B7Inj4
4u1Z97/eBqfYXNCffmbHX7Sf/DC/7idaLd1URhELeunD2eHfmT4vB5qX1lnsS0gS
muVt3jFrgOvThJLKabusWja7+9kx82xMree4ffps4RUi3anuqy++s0Gcz+bbj82E
94us9+FoR0tWMXEtWkCLvC+QOt/dzddvVRIs6wE4OtZKEZCaDGfPfrvSCasUPyzR
6KuTonSYgLbnjCAMBS5W9ZvaYsqrJC9cLWbo4pcbfWACLH6ALks1/iKSuj6QJc7W
wvkalb8KDB5BtWBdU7lFlPN5yQrhlmC550U60NYV4Fkp9RdnpyRVfLhFf3vjivDi
VVxXQ/rMVEA8nIAdKRpAEwmmj4KjX4tZhkGO1ivQANeKpsO3g3PTSR62CHq7JpGB
3+F0vt7loxmw4759wa8eQhSKieq7oNxVQqLG3nG3AqeuOx+ujIMDeUo5sdE1wdIW
LPJe69H966RwXnX8Eh6GAhs6qXEApawJZMEiioEXJK8gDGEtrll/yNP2kLVgY9Pc
2dhiUoOjJfWS+fkP/tc9SalsYzOdeC6YVRdWouKkUbWXpNxITPn9AsC06FEdAmTe
t/71SYGnzGzfUx9VU8vIn5Saif3oArtzutmeCcgCuHxK9l+Y2kCCxqJzlaNFy6zO
AXJ7WbMtT07PisBk0WJjbJ5xUbCsNyjRbMb2EDafwgUu/ydZXnCdO/ir471IVsXP
p0PF6rnVhaOSvcmzBtQlBIeUshB15/9ofWiXAhyAd8ZwsQpWmnD4TVKdb1gfnk4K
sQwqHaJd4GBoDBSfzw+rAG7sBJ9M7Nf8qWYfD+SvgpIUWkbfYgKvJIprErxSSyLH
mbfQqLYaisIKJqQUQG3PKoBtkvgqEyBTmaPg3aoehw63PhX4eelpumgyHRHmYuBJ
j65uZjetkUawG4XqbVWAHvc+gQ5iqxouYYchVjB1a+0nObjzccEp6at1ff/Jm1ny
lek8mEev7bH8jeF9Q1618KzqgGLl+j+TcLBOPBRAY89vbykCt8LK7i/kEy1MUUvN
ubxPPB6WuNqUYHzXgJx65gzxkP8ImvAp9OupMRwrBrL01kYJuFbNPuiI/4Wd8XXm
04J5SjGJHWZjvDmqpj6slCdZ8tThBNruRkC3gi16EigTHwiib1CVicb687taIIZr
lCIPj3p2s1sb6OCrHhtK+l/ls5fylg7wLCRUlU4/pE//x3CSk40tW8wMMXgHEVuD
d9aHu1rsHs5oODtqCtsGZ3bwziVIC+LQd4b5NZVeFEXg+Rq8joZK5Kb39m4fZKhj
5xl7hqhAJ5v8de7E74e8SqcUK2qpkWig5/jsGSC570aGgwisNdHDsJnP5xocgKYm
rQ5V3kBRgGalt4G0PIFoGIEnFYSAjO2nZwzhPMlbbrL9YYZKuAK2QNzVucf1Qi9x
0rNIoZB5ZK5Hs/ai7KvtSdo2BktmG77IYfjHiFccmMufgDJ5VpGcsjAPuoN/hGjp
x3jKGCwsgJGGVbEVOPUMXEVrjVGH30M/12rZdtCC1rImpHqNPZtj4kvxDhlW7la6
1+H8+0ozXBVjP0y6Wf6B1K3Rz8upVpqFfH48I7mH7mUQv32En3qnRqANpog4zaML
b09lmgLErNyEELR2LjoPxhnGK4WH+enVdSSh7auJY6w47x/dKwXFjtw0RCnwZLvN
me6lBext4Yqibl+Z674mbuR/IghlY+yILaRdqQpM/Im2lEERZb3UtCktiYchbqwC
1I7AC0Iud/ObtUbhsEH5NpfJfoG0GOKXzvEk7lYmIbRTyW22Fyd8mviSYvEJhnOl
YexdmtNP8KDVDdY9Zi+R8j2W4C/ppyKkweaz/9dF4eiE0JbvwfLEpoFIHirS4xA1
q8AfWGqct30FysrAeCoOblUqSGAy0KiIPhLXOFAQIrRdiwztWGEw00QPVRxT3zeG
46vMt5ZZxQ1CIBChid7KJVU+JggWPws9ii42xyWGYMpDKwe6BbkT900tVp/JXya5
Hee7QdEc39lN6lEBClipIBunsv7ctX7ITs52IYzwlmthc6gDTb+3b3YXZCI0sPN5
D9f6oAQEyi2VhKP0U9rRl9lnlSyVOnh6oA0/sy90nsvDqviUWKgr7kN09d/SqpKa
Wga4lxBAPXIywaO5jY6lNwcraQk6HsRHjYAq+fgSZBmrDf3ADaVA4CxkLDRvcTC8
yNRet8UIjBwxSju0rBgtfJMmdrU7oQzGY/xrKumIeYRsAsYl6XQb4DCXF1U9lkh0
O5zmSUeGvCFEoDSzblEOXDk9ZaAxucjMMlpNV+9KyLyRj79EOctNgYwPVn6T6zJf
oQeD7R5LB82mKPVMVS/LGvQrpcGpFJWeNEUTOXV50+QE8E26fxiFVFnGYyLKTkGr
F0k+wpD3zsw3ZEAO0h0kT+PD0qNa0f9UDHyCsmk8znto0lTIxFox6oCgnV8gbUNi
I5s7JDqNL3l/7J0I6unCMtVn8+GTSmno525cISL1t6dlpkdVXIM/IM1PBbDbgfrQ
+zT7jdyPARY4mvx6jtN3yw+qbCbNUnkjymmu504D+8u633OvFAHPkDsGL5Jr6T34
3hbBBXqptKcZjjjEcA7zjG3Ft9OxJhaCc6hIqlvGQIc1L+1vvlsuHIOpPepNugLJ
rSLeXYs6rlUxYneCOJ/Ug+vSIBBTqTLIjngtODOy0Thdh1O2Z9A1ceFLXx1C3iYb
A6yWdA8qpWgYzXkSjlNfCxuGGGe8lQSCcxzmqHpsbhoj7tnYCS6UCG6cvJnzDAAL
YknuRsCg1G8KNbROLOLk7U5yVf8yzzsZnmKxq1WV3GQnIEOgcBfrx7uMsS25ePRJ
3uivzSb9ZlNCgiPnu6QZy+7qN1KRS4fqsJyEVnE4VqMvWy+d5cYM5m5vfZ32ECQr
O2qCUwIkA4Isc4wOC7F87uyepxlEFwTZyNHFOkJtWwI0vOr7ha5h1Jr6Tx3UIu34
rjVZGfPIpp2HgBXklt9OHkMIqbcZxaLd66rMluK5c/z3gzP7F04wN/wtMebqzeQ9
mABLeFTJCjCqC5aacGT7ijfpKyWzTC70tyoAXQoKfE954oZH22goYtWo3cJ+atd+
sLzaYxTSEyqpLtj4djmlBZStr3yAg22jqjXHrXwVaGW24bHpOpY+c4vbHUabXjhw
YVp8uKVudrXT3lhidY84zVPX0igQMikPFHJ7E4N5lAbaiccZyvDFHwRjoRwKSBM2
35nuj3QbPcbueq4mkApzZjuBfeusVdgvKu/ZGrvteeY0JHYqVDzQnGDHx7n9sKfn
r8FbW1RnZ5NI1hZId29wzI4A3ItRVFoaECkEDDMevSx7Th4//m5jTwhOahZ6oPyb
kK2K5UW/86kW9YoPZatSzvDz76hsOGDNgyQ137olcAemimTdV+Ik0QAwiSD6o2tG
R82VOxMVGXM592IlrggjhuCAJ1VdfqDBc11+RHNwh1NRT8pBRCvbYInmmWIkUmEW
JRR7giE0kFUqFD3d8nlsopIl4QtrmFihSWI739PZUud4mYx77+M3Zt73wD0Mbcm6
XYEOolNW+DG8E4dopQxKALdSIK5BJ+eSzQx8QKOzBJpQ5si+XuZC9v4g3AUzyVv3
b8BaI1E94wa/ViV0KnksVrtShNEU7q4OBAO3zsy6Mp1vja5lsors9eRhvtmZCxTv
TShtuY0OR5iB3AJyp4I3+bWCWDRkcYEOZG0KK/ceF67M6nqBOuXNKqXysf1ZoFbZ
KYcGlIHD9O9dpSZIxOCjI3rRG8/QRtZjsOdGOnqgoi9G9ejmAhtBeip56x6V9hL9
oPnwAHmnthAUpqk6nzJ+Q/LSC9EoMiyZzR/Us2/I0Xd4nMEtVspbJO8jt3ypM669
LwJftbQC4UdoM70YcSp7VQD3We41r0OZeE9Qgzy3p7lHzaP8cxXBYzMMsuroO2mC
ws5TVW591qITRcl1Nq5CbBwTk2RlzvYRr217jf9vbrm37H7Ut05qkPAfpW9oBJnA
AMRz6XDvY+Iwfq44ZZNyRdC3pNLlCcwnHXkDSQS3E0wyU2CwEoaMu5+pJ9YA+j3e
RqdfaeTgg0zbeSU/HuA+9vhXqi5zLQWwEXg8IvLri75HouODsfBoHOgs9L9uCdOX
3b5l8ijYywhvoMDyLZd0wIe91iGhI2/LFCRbLA95kBOEaVJfy7/8+Yd5rBZ+4Bn5
Ci1mWk/HE1DzkzUUlzGnBpbMEBWdQpKxDMKJk1TYwaPTzaDIxKRG92WC6W7+F/bS
1SwbbRg7JE+IB7ShjXC3wvmqoGITBDYVlfCJFmgx8a+MtQpH1Sg3W3etsHP/ztSS
1BpCSJj+McWfNm3iQfAQ8BWnSzzYnSMqJtlwNC64Wpsr0ZVVy52mYdEHtiipAqTD
pP6MOtXLx28UT+MnK8rvldHNAbT1G4Gq1gjdrWrhsk3aNcIFIw92TIYd2G+/79BV
9cGsbivkrd0qBjbenKoQQR3IprX8no3PAW0TenKTyVhh1otQglFjyT6MnMb1/LLJ
JfkChsz9k0TQ1H8oJR+QLra7vfqpWUMe+q8e6UH32ZqL1QQwkgnm9s9oQrnOHQ0F
2k+Scn9GOg6P3sZ3ZdHRYwRpTYWEJUau+Nv/O7tbPa++Yq8FcvNMrLUDTdv6clo3
mWLby7qNSnyy8PVY/19pJ1/y5b0aKSSaT0eD1ELkTI35EFjKR3F3HzFde1hg8Tpt
VXSPhrWoX3tvMktS6bcymkIOGpySat8/RdCreLboy+wHkpnobiiKN+rWppNGZ4uW
0dryx0Iyf89LKPbOxTUqHOC5Lagi7NwS160QdpvER2ob3MYsc6fZIaARjgnxApAq
LVi8PfSIn7jfl4nXQsJEUZONycU/99o7iGIRvdPMpFZPt2J5cr3YXdIh8vh3hSzE
JmZG6CP8bZLsbFL/33iXwIVErARswQPHBOJAF052/a91L4Q1cYm5EaPNU5i9im3m
ef4VDo9v9rxY1PUwnrqAG281eib7UTpid5s9cJgZUFjeeeoTdumvx4X7ADOWm86A
LEOp/HvNuX5JC9ZSyuq4rCKvwpuUDUscnYpQBVmOI6/uLhjIh9V8vJjrokd8ZP9k
aP5E/vTeKhc2EhuMujr0kWs6WMoors2rvg9pTKedunVzBj9xpN0vyED05N4FtyMd
Rps9CVAIipIEyZrpBvK5jsLL2zvdtVn7NlEzDD+a2278X+04DUcv04enMMdsSiAN
E8hYnsVE0E+8yWK7p1/S4VAvG7KJX7+LHZAqXEKiNHsEWOt5xNrWXPo9zS9rbphd
Iw6Ak9eiF6+yqwXQj68wYvbie3FRvZKj6GRdR7ngyzVVbnlTGz6OAOA0ZWtG/Q74
quQhECARnU9h4ov4Mf9pclKNLk6/rbtsrX9DyYNcAcUb4CCo7MkTtFUYbZTjezpN
Hyq6yvSQG0dwubYbmXBZeLBD+2TRvygbDEn4YhLQPFtNeOXhJqsFPJDCLJNT/4np
prt1DFf7oBqNJw1nEVF/Z6j8Frq41clLKKe+KCxUY2uPL1qXyZjeK3zjSNPl6hwK
KVDV2mqVlkEWysqruSl/U1oSlQKB09Xs/y9t9FmhqbfVOyrb2o4rPGp72xwBFjen
dh2xYeoYHLHrqdM6qHObSvXTZHnhpgHEr6HD9l/bYf0d9y1CddFV4vTcH9VUGtWT
ZWkWb6hysD5RWMjuhQjXh1olbJUFnfaiX9ACAoaf6O2Lvt+BsT0hMoKs7qT39cj6
Jx83cjvVnWfYYAyBQYSN7UnXFgPpdFroyFQxnm/MTbTNU7PygezlzGzT7E5r1kcr
G+FcwkEMF6at4pxELfBVcleUBeLz9PfcTPuIaTU+617ALiuFlBjGwcGnKywYJFqW
+hJpFPolTFr6bK54y4HlRXcwCkvHv5n/+6lE31/lnjHwZtYlXOoiVV/oj00HkGnq
qMN9Rbj02miV6alP6lfmiDpiv8CIhjrJyeGAC3LHqfohwR+EV79zaziB0RRHOFjF
DOfBWxcf4GJT46EEk3ML3MvFpWzLnvyJBzX2HlWM8dhQOwaP/TKLWz+eWyO3K9fR
Oo/G0jobGg6ROLuZHTbVKitaLS4BVqiu1zytnTyzG1/CmGSePJ7xVRMXBlKHfvTC
T2uhF1BPEArxn32Kk9DfqRqw3zbdRJkoAVXWKrV1R/2eqeOxJBgKJ7/xshCUp7Xw
XVp4ClOgupEpDJ4a3bYwGbs+UoI3TETvHlQsr6N6hKyLaGPHCROBYQYf80CxVrD4
esj3nI/IDOFbwFs2DxUUJkJM3FQMzoC9FA18V7GPSb0IC/TACwz+rtb9F2V4+LM5
jWV08nq1dO0F8JhJ6EPLGyqZMBIPiIyVSM+Q4LoUPiDGGPoQwtVmfRygKVy1PG7B
cmIoHEdsaSnJJGZllsumKicHdOk4Qr7E5llh08tHA9PiPhHKa+G4Zy1RJWaaZMNj
XL3UMHlrtTiUF2gYgwGoEtXL8k/Ij6DFyAhDleDICqPlBFgfIT9xQsrnZ2AuGD1X
m63Ty+5r/k0v9xpt1qXt6clEgmrtjg4R9UZ0XELmXrfSF3/mVjNImGvWXvQi9tPO
r7CW5WzxRsz8Yzzw+iALvVW/BUEQpx/WFXYaS5PUXmKFnZ7WliSVLxd1AfVW6vwA
uRMRiFdW2KYKfqlLRBAN+ol1viTO6hVQ8NVAf4X546xiHVxFw8zziXIJgRaFnQ15
4lAIdaOEcXmFIV1DecGZvyTTzJvSDjZqs2jquN2h+s4Ue6fAbFiCOlNvkq7xblgc
4us+QCf4mpTSnfd/OXWG3i5VFnWThi+GtRJarqUlqDqYKz/7HcJmBd1YEea+9SaX
SD09jxWR1088OTBz408pFqFC8fHGMNXysMPnUxeNGy9Dfb2pOjvfB0gh+1KfkUwo
lcNt75fMgjoGYgzfLtm6fPyNxdAGjYSSuV1xWaYIUhp9AVUXo6R/ertpR/jRtuWU
gTdtnlb+g0+6yi1XIlRjTN7Mo7OCtiY8frl34WVY4sltZrXZcvEvdMO2RxEF0wsj
e8GxJl2oF4MeoKIGwEc4+NVCIcJYPKp5QAYbMzzeFqyuV54oQ4VFZMLSkTqBSTNT
GQR35fX3w1attxacgSKrN2yxOWM/kGO+lXbuoQ5td5GEPdFq94SbHQidfqY7+85p
IfGUMJolNIE6XKelUTFAe7+XGffs8EGJ9nOKMAkzKDQhZJLCjy/JBD+IxGhgv5e2
cH+MVV8RXm3eldY1Yn918Dc6e1wbI7TxGPNbPel5lA9p/Vp+7bXnhPnGfl9O2H7m
PKLfoOlhlQ3tow8kNayAKZ/1m5wgrVZf/AbiUsyzMn+eKhbzYBcJYv6+pkxptxes
tH78Hvxc4ldRrbtpcHMvbmoqHqkYotZm/z8zwUK6xQvMMcVuAoN/OjXGy/7X5Zr+
CUR/MHZybbzAinIvOeY/DGJ6B6RKmck9AzjWFbnIoxB9mtyoJOAKtrH3sUpIvga0
UAot1FOB7WwwUhj1FnER2VPFR/X8t0beJknSmFZSX9ko26K9IH3dMqkmHnpHEd7i
U2Yq8k/JPjzT2eDWIO2DAVscriTovSY8cavShmuplUyi5O5S0Y1S0I7qKly1LRp6
ImDB0RcEz4HE6ZZrXIu17g3LgbouAJ8tiTnsqySu6I5asDWBFEPSb56Cwyb+AK/m
zWdheim86iKkmFEH5dgD1An0fr2B3heUJtko0u+0d5o2/JZ0n2buKgTqvF11D0Cr
ti560ZgjFPEFHGFUo/OzGRHGg4+/USf6mcHbW05EuUWyjr8RtaS3LYllsQ+zgvhZ
uwQBc7RK+MgHHSugWP6CIISyzgd411FrT8rwX6jvPLIU84haD/HA6gwD468jM31t
IpnjvsOxoLzqVUQNKqE74CvSxGIiWDKLngb1mNlyCkEakSoIxIpWTIumIQx7SzRe
PtyZAfk0UKTNMX88vsXNehSx7qAybfSaWR3cLXHd0qivt54tKmcBi/dojM3VMW0s
JTLLAVz95A6D34i7Liw7UDnSqFEwzW0ym32MoVBlUswozI7e8n9lYXZ3QsnY7qUW
Qqhql2nBKUD2XheYcaZEuyXAbCbo7wakmpde44RVu2USJh68z25uU16LgRPP7DnB
gsyI042xdqGCC6RfC9yMDiU5ZECagvThqZpx7cpVjXhZhIqhPNReIFsfJRxGO7YF
Bdgs3Ps3Rm+XYFDTk5DWmw==
`protect END_PROTECTED
