`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM9g59DZEQ39Kt860gi7gFD5SUJPxr3x+pZjNOwApWg9
k/b8/IrQGrUCro463zfOS1UbkHorpcrxLIwzWFLLdRkv7QIINbsJwqhTOsp8mZp8
Ebihe8L+AR/QnxtcErE+qelkITSH41IOhBDYqnovJDGd1vko5rWC9Wsvvi/0oxSt
y9N2E/6y2LThXb0+/jEu4nqcFncYxH/U/oP7gyf/x9DPHg9RrkGSvfiIF8Fxd8tZ
kv+x/LREnXJNYh5L9oe/1aXVObxeA3+vm1yFiyQn7U4wgzwYlIGr20m2R4pdzr03
LZDigrS6uPRw9z65Fto0xdS0+Nbu47LXXTioTxtZeY8LvAOtSiX2mC5/0w+62dQ1
Scooxhjy8hbfFdhws3lcafHAGiqaEJjmLnfM+BSxdbDulY4DZI2otbFg3ACNAxNn
`protect END_PROTECTED
