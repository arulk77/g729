`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
7LYDZYe0waC708W13y/9fYOc0YQOB0139aBFHMghlqi5lnqsPmBgZt3E6wjfbaxL
lV5i5n7xe+zUN5t85Qff6Miy0d0pJ5klW3xHbwrTkcSeT1f8g+Ssl4H0Ky0lQxQd
A5EkIDOMw0kGQx0NqsK+7kj2fqKnCF8W77YJADLnExvz61FiqeTPGfPHT2JoucBO
I6+8CnhlmA7cACddoAZL6RC+D7vMiIdSXK/QGyVu4Of/64wFOuc+CDXcoL4deHZ5
8+NnoRmNY+k0iV1eelhUcb9Q92QoLEUUkF1o2hUR2OxdFrlCWX33xUp7k+5IGeJq
BGmuojRpy/3T7XYgTo9QB/UflTJkaiYk5qZAjNqOD5G1YDlNcRrjwShaWIVUcy0x
YQeyWHthFLIZK0T3qpHndYc+nd9BKiD191j+CSSQLgzVG+pPsEPdqn2lIl0iWjgZ
V/d3dSz803rUBZDOVD+LeK2iJscW/pJ3s+/wkWCQ+5UjTicKW8V1yO1ocQ+PfRpL
eVC+R+ypphDRRmTA+eMX0kSR3paarOwANqSziyuI7C29YrBB6WmsSKVVsQxYLB++
HqNJAt6V/sgth8R2rH75fMC7PnU5tSHeq5e5E7Gcq3vFMv+7yqDy4cNqq6Tux0BW
l1IlRdFWrZ8SvzKGGI7r+PE7OM2mPYzQLn5RTylONHqXQADa2VPqvvQ7hQDTCMgh
Ear7xW2u5N5X00WA5/PDTc373dQUBGWbdyyruDBkPWEMhTV0A06wtvM5cfQvJati
aRQFesC6axp4LAX+PJXx2foWBifUHN/VYDuJhX3Qj3dK1Fcgm1vuTienj45b9BTY
OwvYOadjo8giBcdNqcrLqLJCxuxe4NY88/bimo8WF93v62K7jMGzdhjPfjY/cdHl
QSnlenuo1ZDaTjETQt/c1JfiptROLhO3zSXNGz6NQqr9dCeoBbX/wHkBAyKB+YuU
QEa0w0gjJQxqYyYRQ0ouv68tXLuHeVgMaurOH4rhDm1iUzUHAqG85bj1U1y7Hriv
omsCKg6JxwrHL0b3UeSdIYFoLGY38jsr2tCTiFk6S/vDRhJ2F9Q6cgr4AsFOmKU2
TdnAcSSL/kbnpieP+1C48IXS8f1YIbtCjkK83hWO5om00JE6YEH3IOqnpynCU2MI
L3J3LOJ7L3582RInsDZ4uhdJLGWrbT282ktT+ukkEeHFfEW3HiDSXj21sAcvmvYB
8QsoAPSR1cAzpRc7sdPjWWkLyity9jtCoTxIEl1j1ZPGYKbL8aT/VOds6oeynQzn
NADijJcdBVn6eNdAjNSVkNXnWjoxobLbIpzTyn2aSwHj2Db4WniQP6RPZsn+5v/n
FD+gPTmNtkv8Yt8g01vVvKHAZZI7Xz6nFIs2zFkNkFjOFqXiIymxuLQAB/b24sEZ
2eRN/g1bFmh11YGcEHUkgaARfW8Vz4AuEOpCL0+SSJ+c1cmCM/9WWne8wFOCAh+F
OthpnyOz/tvyOpYG6SpxK0ATts1SY0jLPg6NerXrVQ+tz7aVGF2AEI3gBF/fBoav
cL/W7fxCeTgkCaMYHNsDIdJMDVo8Uwbta1TjAt2Kn10r64ADLYm7z8+UJ89L2qC+
Gy4/MzHWsM4zP2vpdbUl3gkIYnQS/nhUTwHcxKXhefU9phn++q4NiQcAJrGqXS2+
FsdTtNT7DMQuu8iJwqFq9O7F8T40i1+7fDWgJkjkorjcjIpwgGnPyGX4gL15OsQG
t5cRr9EA/8400mNRvYUOCr6a0rQUHQHU2GANC3XD4PdjuWTwYjWCxrBWjuub7ZGs
UW4qf83Rm39BwX7qhrDMYqhUKAJuDTBEVqV35I0W2C6UqmlyCITDp9GJc+T9VRiD
KA7FJ0MNF5W/jfaEVIYr0nj8DiHocu7W1NEb4lnNMqjtbNmrkbH+l2IgY2bHZnN1
orv9i6jLMcumXM0c4jK81pMljWtI+E10gOgFLZq/sbzY9hd/eEhSEsLdDIst9PVf
2mL/DoRy3ut+M+7pVeu5Yp7cT4miuRRFUtqlw2QXm3NirlOL05gkAN7njZPNqxLQ
sqc9Clnr2d8iS+HsZ1p5pQT8zkE0rMy7ZLo7uXvUygM1us3gHIAtg3GiVvv8FEwk
oOrHgl766Stu0MFLDgiX2YN9aFQaXJRTfBILRW2wWm3Jlo8EYoOWULn5uDZO5GR8
/XxXJL1+vn/NiyoeKIuIlbkk6GknMTum2ieL2iqMMGRGXnay0qKc0CvwNPYsWlnF
JGR5sbbQcI/goIWq8G8Fo/MiucKr5cu6pruzrMLN6QQlk4mIYLje9yEWWyXNV7uc
`protect END_PROTECTED
