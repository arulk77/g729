`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
HXUqKiGzJzopEMbBLk8kmdEKYQ+Fr+Ssiyt23QXUqXrTlLYJ12EgaZMEsjOAeysw
2ML2I05MVPAusRklIfc4Qb9vCcE/HPGLz2ozvvKNZUn/MUpq1qFLzWlirVzCOF/u
C7URxG1aoD41ZHuJwEdzwL2AriOIY8XEVh0H1bwZ2/J6+zI57SVFVSc6eLnVOBQj
8qw6sciCnxfAQ4HYzHouLwVFB5IYEn3IF/VPSl43WCtDhqaakP+7b6NtRalkwWM7
uFOsGFuVVpD5WZwiP7iqfUWnXuSEFJcs9flgoAEiitD1LMOehQ6s/q0Nijx0zkGO
ZA60w2NVVAp22lQibqIWGG7Q4WrMEQh1718iqoyiS1Szmx4Z24L814BJIEJPIXYW
JGeBNTHyZUg2Dtuy0lKM4UXFFZu8IcVLTD6m5AhoWq0FWz/pq18+hH56SX7tWjSq
u1wu1MvBV2wtT78tLrK6A7P4KK4VzMANUt7yGxpwb2/RetB7N9rsnflGBomNTyTc
yBAQk9nHu2ofb1ZcFvCLyQ9MC4e/El9sl/+Sh2FBExlq13LmiuwFuIE46pc/kGtd
UYGt+owVzYB2AihKkL04BoemsH1nFThIhvbyn7ezKGlfnzcf5lOurKzbsSMtoGlc
ybLmjUrZRecUQ0RT8vBSnnK3on2h57DeJInqZgoQTpBPX/J3wWFzBF3a0Et9vsx0
qVIazKRUY1m78Q0hzODePN9i0Y1RlKLbLjm9QYxlDJMMZ8PIgEjVyBSErb1BMdY6
z/yOYao2P79C0SU5MzsK9SMI5yPe25EEI8NKPg4mXoon9ZxbN2hgSg3BRxsnKbzy
JzvcaNiSTryA7bsgS+FbyWhFd9i8tGNg0Wtz3BhSSOdj0JL5X4YiXauENQwefYzA
5kuCo7t4F3OFRYrF2svx0b6BP/D1PJlDYDI+FAxxiL9DLJg9P0DewyXvU1x2SzZv
J2WrUB/iyF17duRiETJZXtWMWHpIuXtUtsxDIvshAk5XKTjWg0tyLB2endaBYKz+
HbQV90E5MH3ktmXYMPm+aY9vSCOcziFOzmVDr7iNoghocKlUJK6UGF5nhCTB8T36
/D3+6+sKDPJks24oLyDBtuf279m3Rm9mb/G4AXhHGlqkJVoEkhBU679CkWi6nhIK
z5Hy20Tv3TNnsgDPC3veEfDznlqHTs2CUdRda8Xdp+MZVRrwZu6qSm1wEyjwxq5V
u8lg+lvKwh0a87hY3F9r0iW+v2ti+9/0oUqw/TtvGY6winnJ/ET/FOtqnCrdOzVV
puTtRh3P+kbHRwXGNCqE+5mE0i+L5hxp2lVSiM/dT6sW+sgGuz4pRoVib0PjrvlK
FGPn6rn+G1Dlb4WxH/E5QOM9Cx8uMAYve0EQUrwXFFxuke3sBAf7lxGxqPKsFnVT
PNyiYo9f/3PiSmNFOinh+Og8WOaEkrzUx1DjqCbcwnCd1TmChySwofenlwFpH7nr
DTC5LK2fFOYZIPs8lgb7NC1lVr6puqBnd2mP9fVlmBdKoNFuM2L4WH95wxZDjFRq
5LSY8CZ4YSj1Hfh78UTyfhzGrIFYEPpqBQJMyYetsdgxISC77r9ufiW9n6HHR4kn
K3nZctpMr8FT+u3qPkCV5j6TXIxRqKxuUxdbT0Qn08/WR74btSMKDV0Cvp7Y2WiX
y51FElXyC7sgb5s8zStJ5VE+E6WgNPceVeVWxKZ0fPp1B4G8REUPVTU1uDXh/eVZ
A5IPxLBVNf9y6tkMXF+kkAKPNHVK8TUY8diTE6drm4MpdM3AucgGX9wZzMCxeJC9
JhwujLxKB7DWicoWZASC+qyyuvFNgk3y3I1ird1pBK4JwCtHvxfu6TtEd71L8DPC
yOhuSfOimITuQTZToitlw9ucHdW4yMW/l5dW2XCnydpD6u+XcjkzGGp3Ue5hrvDa
RaUb/R0f6C4qnEWYSpWGTcscDK895Tc2urz159CS3zcxCYfxgrRJfs4MvASefqhT
is/r6hz8IM4d85RPRDBVC0Z7SVBey7YieOBFmhQii306czq8IxuIgz5N7dCNBHyN
aJ1zM4V2zcWmCb/AJ8hgm1Fd4gMyRyPdLJbcIk3dRIpWsfdyIMsdTf5odUVsDmUR
L4gQtYfoBZex3c9BlzsWRZrEkQ3cJnVGEF1BOat+To+0gRvSF/AhLazVyhelaeyZ
tpUyQhfSVWniD3KC3DS1ia95vF9LQgivi7nR6WMVemedPEchFlFeyZOFZBBmcF+6
NUlJjQNJ2m8E948hUJZi+faZbttowzjty7e1o0zhD8NjATwwcGKjEitelMOTwhbp
vkzLgHTo9dbWffGTJntpc8OQcBuQbpAGygK+zHCZITzMUpynkdbAJAvFdjMZpMyh
QgMwhb03TLdqy4CM9dzrSWnwOVkpcPpUbnOV0ajXRvyeOJTU/9FBSEiYim6DQE+A
hNYYRPV5TXjizEDU6XAH+NwXnWwBj4MOFlHmQvgzh4c/pbbLToM8m5g29uhpu/Mk
DBWmR22WCbdRtbwbQBUJ/l8l8j9/Ttpg6H+BkFLN7dnNCZ5vW+OTWpA0o1h5pXw7
e1BRjURxtl+ob836Z43ad05ZBG4L/6mzFqneXCfAHoDd+ByOqwFIL21/HFHvEt8n
pgVPU6mbbADfMxiZf/jbaGjZggbIHDVnPAaUkNfOTNeYsUobfjg5jM1kepYnyRNF
8aZyoYv36QpTn8DDR0qvux+FY5t6bpERh+1krG+pS3KUZ6b0wUKHX9Z0BmkxZolx
Gwy10lJAilBjsCTBYQDoKiHI1dWoFveRCB/bPwFzwvd7SScnaM92CM6XHoY+9xHF
WGYGOFBOfXXpO31fcRgxc8L0kxv0poPX4VEd3qcquAagR+VqI1kXwUrGh/kcD7zM
N9OCvgmsYXsYqtuE3zG+vIGqYXDxvdRQPL4bNBJoahxPFT1DbJRb1fJa5WGBcAZT
2Q2lB8G2XTSmbb/QnwTfxgYTFDLKTjPL8hHuwh7qWjaN44pjdWmYNGREiAXykutQ
dwJyg5GcpRbe4dFxPaX6mC4sUxrDmT4NppTB7jGBBtM=
`protect END_PROTECTED
