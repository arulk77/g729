`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
9OD1VINrRNU+cWz+vz2AcvX1jeX0KOgLhXus3M2bFh6MD7BdvwfoljO8lII4VTR1
/kL9DK612jyk2Y6F8PdNgbZ8gPDlbzuLVGJ2jFhexjnBAi4wWuK4zEdXgr4JzPDV
GZf+oiv+Fus4x8PD6M/PkwXNi0YwdXbWS0cm9H8+yFB2wcwL5VVoS5xbJyj4Qv6g
Iu3ywihu5FgjwoAcpuWkNX0RmNQPnIp8Xp8fjq4iaYrxvTe2TsdGmph1mxp5mcWD
16n0j0faFUsuyqero90n8JA1XGOZkfqZiApAN0+8fiI4KsZ036dSgd5zrJfvyBy8
MgdOQT6oRRtaWY/KPFGjU5liMJcwGRfXXohi1+ZWhnNvs8+YP5JTllg8PHiSkAQI
laraFUffrjhElN6OnKzbbHUqrf3hOlg+l6OvLK2YYvDA18lb70D5J3WvdVcFFdCA
OEYzjNluhvwKpqYFYjLbCqdG7xD5CD1Id645pCfjdlxdzX9qV2flDMhaokCe2MZv
P4mRti4QvTBiqhNf2X0Sbw==
`protect END_PROTECTED
