`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C2koylVHXsgstbzIJqYzp+ViAuRyh6jzmuH3V23Mo83Q
2bcDH9U2C4uWM1YtNs3ajfr/nneQYfRgUoyvhIbrnLpU2bi0Q64l/b/W2uUSTwve
AWWSHe6a7JB1YVWmeWcWYlal7m5BwrqQ6vQQeLgOitko7a4M+P2cpkSp90To6cam
5rUDDkGuMNCbJgRP0W4FTacatUzS3n2jN5iiaX3eTobQnpuWsqpssWuVA7zP7eT2
KT5lKUQPKLZHk0jTXgr32pEHzhetB8UJiwSyRLdFr0LFJbyleOWXoEn2qlQ0h+fW
l/Q/3KRdOmWvfNiK9uNrXe81f6HdvswV99A43GIAsZDRzgNBz5Xu6GTIh6lDpXZE
RvQ/Q1U+OkfbwQi1ZPJ4pEYyK9D+ltKj+cF3OImp+hNhRRTr++EyEb/J9e2GUd8+
ifcOVfyQ4wkZb4G7q/AuDfmqNsuq+P2ObvaNer7t2Hp+mF4NIpaEQU0r+QxaiKng
BrYU+79Vwfs+5HKcpA8n8/2Zflf9GQF1Uyq3eds/YhWu0YswJgqO9g+jRXK/Z+tc
Xw2WxUrKsLQ+2qAMMJINX8PSABjkio5F0xlin7TFdQ0=
`protect END_PROTECTED
