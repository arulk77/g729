`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEsjcUB+SxEIDeDY5r/kd33UWya9aku26Api5k1HrifO
rZm8YRJs+NMzUGx72nw8uKRLIFRPezIlRV6SvB2A88JWtDBYDpYhrjXdbvruu0Lp
rSqxrF719pUK8YUUTYaB5Ja2Kpt+DMluIB2pDbmUClrvxsKe7IW0+pW1RmOlVA+/
VFruWyfxXc/XrzQcQNc0BbiWugyU9YRuMXCat4AK38WCCesHVfllPllG0wOSrk3n
b4XrhL4k1XECQ15wMNRyfrsuB1Ndvsoj4gasbd+jcc4WWIFrkAKl4hlJT+ItLcg+
i1tznDEEruVEkrYTVPtQ2NxaXdpSerXSdN2o5EHXU7Sb4WmFUPvKfptwvd5VpO9l
eHLIt7C1SDGHfKjl7OpDcWKnklkrpRs9zzIVViB/npEzZbZV6SE2cMiXDSlif84a
IUZO53douo4bTQXO1XwN66RIT9tHGAqjabVXUeI4bP/82JrmcSLDaW6BzgwZZ32e
92vjwW7vOu0JywMKtdmh4VdgyaPjrRfVixTtz3cPxJHvshCLWHMi59kFCLV+D+fa
OJPpuTaskIOD4TfnT22cm3qEViPg32zhBF6fhd236S4/YMtquGvWGWPBZiU/EmS0
tMr0jt8jo+qwfamE4xGE4YywxG/Wggv6W/sA5n2ItnkNxtcxac50bGy5f+mMkUQV
T9xCT2vRw/KNF02mWhOguF46KR7Ef2DiNgdzUT7JGYUcaCMkH9rQYfLyqnYW10+B
py6Vb2CaBw099+mNB3+vYBzPEQSmqco8P2t5JF4k5TYEjY+1YuY7qikbW86o9Bej
BaJ+4ppcmq1q3MT7lzUjSXe1mw2EQ5EoGN4J6pVc0LY=
`protect END_PROTECTED
