`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pHzzam8aunU0yp3D3VXJ0qwlwHX4udqzvqGRo21rSuxp1p8opJpaOrupx5l858FT
RnU4zmAoucaTS2b62/KA+bX5q+xKniPiQ1s2ZPe/ecWHTpzxVY+2guUJnDfWd1p3
GSgqW+2NVDLywVOxL0Vbrop8fD+kPp2CqgE3wVzrZT6CY1sJHvWdl3YItxW0gyZA
Bx8RDPMyqXiIQgqmPXTHuLj5wlaoKWhdGiWJJNC3hZH9mC7ssgLHhu0pupLnNlQB
iRxUebS1H8JYDJtLXWSx0mevzLUgiPc+aFFtUbKr2XuFXCk5ClglhnaOxyoR7LEy
9byfzDwUoBjGTUBzELi6sB4QFlyAZXYuXm+8WQPkJlqWlalsvpWxJlJOL/JCdq52
oaAy0GCGuzDwnFSztYIyjWc+lEyWFfq26yfKt5Qjpbf+AVOtA6gxna59B5vSzVO6
hyiWY9qRFL+FZUoElZz/Ywhb/q7JZFKeYinzwXwi1PvJzfOK9+EmhhlvxBHqDETy
4dzlmG47H7VLuzeJmR4oDleptiRm9LNGjq+JYU7zvWS80bm6xwTPD94Qo0aubvzQ
8iiVc1HBFGtjWGtZ9Qquu7QJmF6XrZZRqlzBG7h5ZLxN65c0XdqPkUU7OqrMVo3T
TycNjFjTVsOlu895wigRwnJWY7n0/oiD6x9xxfKdA/C+xz4ucyOvdY1xKsWYBN+Z
L8Lb0cQeDyZyfuxPxjVb/0Mz8GvSoMEhFULfn7LYd/ukRWzmW4Lw/1gfgcR78qQq
4PDmK5Hn368sEgfTD2ZDqg==
`protect END_PROTECTED
