`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGO6tUup5KYi4JdWGL66OewIfqiQLFn+BVK+sMQUlzIc
GujIpjjctElO1bbuZO+a8ZvUyJNc+QMYOu6pFB2wk8Df6/a2ZeyQ98bG0wreRmVq
4GQ0KYHqh71axcaKlu33trTSrU3GkZsPm4VGQML/6x7HZyU/mXWl6fDLzEPKLvg0
jcbmMIpwUuHQdpYOFj94PQ==
`protect END_PROTECTED
