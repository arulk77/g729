`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAcUAHUx03gtlxHQxJp+m3180U1PpfWX5hmPmzEBOSy4B
5SQ0ti/V3Zqzz59EAXZ53Nbn2ROHlwfOvpbl5DMqkDFzELIr2lXPFqsFdPDqmxUE
4twtlLJsbclQgje4WA80sWow7xfA6H2XdUTUedRdZlVCtfjlIf1O1a6S/+CXb6O3
N19nziuTBugPydSEpoabTI9VyJbO09d9CHgLCL+ijpmWdPzMLBwHjxEcKdkFa1JK
MVzKH7yQFhOENk1QlGp5fdfHNly4/HoYBAxaEglz+BgfMOpmdpTrmR4iBYiUq4hz
kanej5Wn8tek1opvEIWFxste2lCkob1QwJgZyN80HLrRtIlaetF1kBzknnOaZp37
d8rHJ5VPs7pcOMvayicQ+hKXHdrwY5SN5rrFxr4O+M6iG7eRM9ywuPZjafiu6CmX
r8y1acN/msCTGaOzs3IAAgvbxDO7ATyZkWWjdFrtgvbtbxuHJQ3DS4X6HX3wpAvl
/eoxmvNkX9E1G8mYU0TggC2T0NSbanVepODEtrvYtgAYosObcuLtlk73x0DjTzRi
RD6+1EijsoxZMPgdwVRMAWVBSWsfD6aUMTkvWN92qv0LON9MR8/+t75IAaKvkvoO
kt3dKUePWlmIeKyZmkeO02Zxwj6eybgRLojBbnC3WT9W6DSyOxDkyLOuKAlx46wv
6KiM6w2whQPF4trQG6EgAv+AD44YRkdWb+ql1xsxJ2FtEk5mXHZgEm6Uhq/EfcgK
EWdKxHnlrUVzA3mDYDcgU5MHT/tCrNXuzhAfpwvAuhahPhSgA/0B9P8mBSSwd5Ym
SPYVQehedoe1fUUFV/0e5U8b6KR5KwCvI657T4iTaAU2HXq1ItQzXcGP1bCvFPBE
RXcIAj0f+YWe01Sb5cnrF/1OaenGC2rkfBxFe7zxec/A2TFc7UBANApOIZu8jj74
V6TvHLJ/oM8wUqA+4TW3dYTf+rZhwalCQdisDKGbWkS29bWgExx/0UbtwTmRSr5T
vEt4dZ07P83lSBcEILtA9eiaACXKpZ6WBLGPxG2pECnVsS7/EQQn9sf/RLmWYdNL
BCjUnO5Es4BofkYYImXSHjqba59zL9AVmYSfeG2m63J8z4zvZSfVrjAriUfzzwFH
TpUJ8gW9+eaztDAbxId/XLDY7eyC9XcR+mHGLb+dM4njnQf3aXg4on2fyLUfrK9B
w2JEmJW20ChhgK+SbaoNGqRTq16Fod9pHifxmnQJTXgkOg/HfabfumzH7CYeCPlD
pliZpp1MS+wC3hna7nEomDBzw03zgu7fY6dXygXRE/m3D9+Z4fJG/5BUu3pms+Pf
SLpHgXKtB3UOSDEpxL+ulujdM9+AtBlzXcLquQds1+eo2DEmhvZbxto4Ogg52B7r
pj+FRZK+MWkMFXnc4wlBQlSCreFWPXDeA+N1UCDDlir+hpRKxCCl/rJJ05OHHc4o
jUyQKLm0iHLUciNr5pvn8G/xohkBd13WJzB5zSyrbMAsDfjAuFUrk9n2Tz3tqevJ
+CHALnV7exgUwU0O3qtCOmZCY9yc2JhIiNF6VJ8Xszi606nvuaANiHN6pT1ndtt+
PurCI5l6ZUXY2bMaFiDBdfKWsuhxR3KaQlyG9Rizo5ZtCuQi2ho17eZuk7OVcMdT
3aOblj2g/YPcfZs4sI4ERn2v+8gwfkOhFoI/Kiw/N46zyc2sXG6CQBikG8eFZpUo
SVfyUAeRdfbb+5RqpASCb7Vh7Qhrn7dMDO4en3z7qP+tNYZu8Gb1Hnzv/y45UAe2
azDamcBEGOAs8CyZGvd5yJkjsLyrzjERR3GhYQO9eVnNJWHUbPb5mtAD4itairOK
mv7PPWBl96mNiBG/MeqxLExlXv+lHv30cmEA0XQk7+gOOPf9LSPDZbb6kyyk+BL2
uoCKvi9RBBOR4kN02ac5OfrpBjDewk69futfmvLtw29rarXjKLfMpiiYppXwOsoA
5iapBvq6L0+or6BegNqvLj+dwVGOB4ag25uiVn9P0CX3F72k81zHyerqfwoKAJic
e0FCLus/4r31I/BkPWj8WGOXw0k8KJwJic47E789Ofu/qS1wK++wa1dYbUIjpvYK
jCMvpsESqLXibYRlQi4reXHxZu9d1XZdf1mXdwYmGp8+yrAwR3J4XL41jtR+daQ9
ByyVfVx548JwEf9x05X4WeC5AwN9fp+iTwi/aMF4JaBzp22ESrCuSlQ4L4CO7Nqh
Do91XZmTRHreV8XpQ/dTNC6r/srEd4YcHwgDmyVwem3RloNxaXZ1zMExOwwymWNg
XA6FNgM2AuDW6i9IzOnZ7Xph5tQPiH/XWghHTBv/kZ3VwDqO8FaXn9KOEt5/Ff0r
fef0F+xX8gREBn/JP5REfSrGNayupMkX+iHccr2/EnG8uL3Lc86pRbiQq7moH9ls
zXlL8mmlICXAstgljTSJoDMn7vqM+5a9JidblzXyQzYkaTeUXzNdSwaesqwDjLlW
ETcKqR7i5AXAcDGe9s0Q5tU3KbKfVIBO+MPuODDYaprn1mI5NA96rLZIuyN+x5v1
MD6ifRC/oOCS+e+8+GR2llAEHR5bFVeKj39xe5EAHVayt/1oApvH4MX1kKWFqqFI
8r/REeK6h9UNwUai98gqzCOW4raL0/8shJbZVULJ7t1xVSL/2df2clLuyTYFXc07
rAafqbCxHZUpqR6xMz2/ZzS1OlDCe9FXbdDjuexbKVIybNQ8qqkKlvHKPhWUsofF
WhpX7Ka5DBjeHyv2YLmvYYqYDBiosU/AtRJw3Mn82I5k0T6w+tGbeHc2QmG6ZC4j
edCgiT1763/jMlSWBq1h/k2in3BGeIsxUvIWnhx+XBQBsuwiSlqm8DFISdaNnwq1
r/2ek2FkoCfEMJhB88oKUN7pzN8G77V1L/IgpkelPPc1do7liv7V7kIH5jTHb4y9
+3Ye/7DEDmoHKlxUABPL61WrjqdIIAVM8ILsuLx/xCXX4k/eqVs7Em1VkXBHpDzR
Tu2/4uLeYeWieT3lhxTOv5T7uFQkdULbws8rgn7JRROOIweHdHct6lfOC4tDI2wW
AncDdT/HmD51ifDDPXdgkLS38UNSzQ606jkfDf22XtCJ0viWKYXNRh4h6A4pbU1m
prdJOIN0x0O5upyOU60ttaNOb7hAjFDqM00f4oA69eozBSEyhGOsPKr+a68Tadaf
xoJGXduoQFeNMJMZ+YEVpELT+YUuU8gjUDErbWZxz9wo8OYnGxF7IrNu8STKKv8b
km0Ag8u8rCSQHhGJY7WhYW44dQbvxycEbFnEdVW+jSK/1npNktdf72UjYx6HllQT
EDBwFWBJ3XQAJDUC2sDGCapVXwXqlNOF8sVv3+8DJn0E/7fQmgZ7FhVAB2aldA+1
A2w0JirFP8QTlH/8qXlb8hqatePz+7Ub0ym6s2vsBgK2MEObw2DKonasKWTwye+i
Z67UKNhFEUSVggFEud5q5F12Pix7YHYNX4/4gLEIUQidEGvp34a/gt6vr/kQI75T
0cRcQJyOOrxKodpeoDsOlccEu+v8tn6TC8qgm0rSpBPCAqEdT3JFPz9Tq033u3Ns
h/sbwIyb8mEsZHFE1wpZtlswbJv2ZmQ91Ie26XP+vGJzp+gBpPbRk0Lpg1I3c3PU
K403/gyBv2B4m8vzHMTtCsOBjqIwwSKdKxv88CK2arTMCLkfxIU+EpSN/dyyVGg/
a9PZDb0v7H99ms+KSpzeFuIUPTk2lZ68GcRyPRTI6gq3XatvdR9da8OlqmCk8Loz
FN82EFnhCwzlXv51twoEA/dWfdpudpauEuykvLgQAaGwxf7g0xDSmEXKkJ+b9WOx
fylABKabTup93aHHRTSG7x0M1Rw+hdjcSVtnwPkWHjz2ZnyGMCDUzXACXNYlLnEb
rsFtcjDy7mPZ2wIE6wF8akf3eoF7Iuj7FavtOhLks44Q7+yk3JzsPUyzpnviyD8V
raTkK+LVWO2pMxZ7/FMRAPDSNXOcLueMa0goYOI7OvXlfwnQEyUrsUnDT6N2s1H9
GY08/T/cqHzkg1YB8Kpt0jupILDZ7uxmvcRvHIymfnYM9rQZ7yOWxX0PWJlnSxBz
13W3l7WsJAc+VDX9ESIXEPsxFbxtdjg+b529lIS3hAAwmQZ8gS4J0Ske+noHFooz
JPlW1UrsoCbnmORrLxBAI8orN6uyhkDEY7Op+tApaQBAI68N26BLZo9OoF7H6T7N
F3vHfH+FEdcNJzPfxuH/ZE4H4jkJ5XvYbxhZgZsC8pm8cdRjlKv3CvvsQ5j8dIFM
lCvA5JFhvlaqII1IepIpD8LGAUCwM2k+juC7CQMzYac66ZeVvryP7Lf6YBJGr2Bv
xwR7nSHSPAK7hxcwhAwZtidLjPO0XSbxVJ6UlV7DkwfSf1/R0wX9Ams+j8dvdUeL
uF++v/4Z1IvRydeAW9qx87UC9qiII2QRhOZYEQ27/4PHZ1k+qx0Gktft5FyBtN6h
UTKTQ99n8ZSYlAIgYIeLGPdpVTvZBcg0Gsd5X4rKCx4PUR4D42MHFC0ShNYdWEI4
+szC6YdFQR8wlBZevjXj+GOvkp6uZ79Wo0+96vEBjqkc4f6IJpc2Zr9Ywnk+1v9c
KvNQMaKmDMaD01F8ibLg1xsehV3CJO2vhwoHNqTCPa/+LcrB/fpuhEoHNjWZ62Q8
gnBJ6/2RPS27TPxduzwIY0hyD2nAu7EHuCSzGiDVTDTATbt+bKHbfGG65291KaGm
C4QLjkUAB5Md3T2FbNGxsEiPcOxIICsYh3z0sShllZLXwKfbI9zqqhOA/F0EyeR/
dQ3Ah+t9eJeggk4cfzMND/Elb+jF8TijBgPuhWTUZmNYuwlK3PMM0qWacPiWjH00
whaqwNafnzRYSleeaM5YQl7XbNEWk8828tU+WHSP4v91PccLkbcMsUab2A98R20M
my7/csWVVY2lzlulGthnVgrb79JyhxBo5mgo0Mkzpf4x95BcYanF7mlB2qdW7tU+
0nTkh+asgfVFEapbm1skGtF0duOB6QaZhod/UQNHxDO5RNluEpdoXLKkSymZ4Mvj
RkvMfBn+UHmvk+ShW3r8KE3gGerJ9s146J5OO37fk2oruB9W6G8Lmakvh1f3WxLP
Ic65iArY2P5a4itCxd+rbs02gMGwTgfOkn+7dnaNqxNEfs/LoJdNpodzTlhWudWL
BOzrwNpWdqCPpt2XgwlucvfTrgRQpo45qykvTYjMD4lQcLybCxds8Tmdx6VnQ9G0
nP7RuUdSk0wAH+W0WI4w0rSw0SokjOhypUJi37fM4tCMS5bjMSMUd4SgUh3Y/DrQ
xZdCOKEimIziAws5IDNEbfCFgkKdddYkylaxEHBVkt+c9tru5iiSpUttPBo48K9Q
CYLaJZzwb4Q0fGTdYae0TM6a7zLTf7VX8Rc2UlWiJbY6l9IvbydxNqtZ2emIlOgr
/r0yQHBYMWbrNsDNOYgVWboCi4REdbpp43mlxqaU9JFwoNSmB1qVz6f4GPprWJA0
DtDXS0xsfY43y4VwqEVXO0sCZ6s8goAKnWrqFrFTBMuuVI2WqFnHIoEdyS1cZo3p
MvgN4utgULU/8UNUlPScMC+c+IrsKl6HG7br0880OcQpiy6HMy+CpL304NMaPPdQ
AXuVL9y4m5LGwXo5FOvG4idUbgyQaV4GDWEvR1z4yoD17AB++OYUcCjCUU3adP99
tXXWB/9FSy9vyo3xUW4/KZqIy0DcuBRYpNubzwFtE418oJnEb1UfVExByzjBGIS4
j3OMSJWadkw3IsMy9iijNSnqvimdyzKLqd1E4lABNuJ3dwzQQkDbN8RkSyGddd0O
W+9oPdZ4oyWLS3Ohsrlt+0ff+N/o84evK97ucMyprbU1ATbh1Xkvs4Nxns9rq3g8
o7o832uqHA3kW41rpZp0+f9tgTwSLxtOmJa8GhcaUrCwT98Sqr7NFqkB2mwy0Uz3
i+ZmPr0xNe2/DW6H2pJQ+Xu+rmXDDWWQQAhNOxoIHhpEiLUFuGknJ43xkhd2Mc/j
uHc6e6Lqv9vSqt3WcW5Xa8xXrOLgGrI1Cw6PewGveNhlsGJeIGRoLWu7fsTa0/PV
NGTUgBLxY3EqNT3oSXYm+UO3g3HIrExaq+VmSM/xWPtlZFsyumGU50b4mbE7JE4s
p0KEFZiO53C5RfFRSOhf43OqBNA5D0ri0y9mmKs75b+scqi88FR8omc3cM/cDrJj
bj/AhON6BaVroBueBKGOe2L7wKi5H7Uilr0c/sYDeH8R4GDDIwHWPpCHQQaS9cpU
hIzWS+5QE0k2GnwGr7huIn/Oa64HUijKyRxByjHEjFuO8xfbub4oVJTd+VfhpSlN
VX4uzaDRJrSpre/abPLVsB4s3yuw4msOZiQIyfh2MK+DHLIJtCwL5BR0NMZQt72p
wMWEZqjj7fIA/vJYGyAEi6OChINxv5ktrizBN6MDONYt+ZI7/TucePN/XTzQYXcc
vusjZX6WSIIS0PGYzW5lOkyUCN+I/YkfEH+50cEav0sj/NKXZPR+qgxWcOhijJeP
BNa3vI0oDMg1P5yrrGi4MpXFH+PKZJvpJqyMO9rVFLQgQINSa6XF8ZYFi26UwcvA
RiNl3EjQPXHl0TQ0z5vggTOcBW2voTOA8vyp/ZE2fKs5qLAdMucc6CROf1AZIlKG
zPYN/6/i4VSteR+3Rc6cRGKtYxdKDWzZwrmTe/ceu8gMux6kdAHVIFM/oV3rlVwK
Gz++7czOxJv4CeAOXrAeK2IrZzfSY1oVSswJoAdxVVoIXbr6IBPiKvoT+0NM5pAm
Z/T6iTAS61lhkbb7KxTf2scBc6nfIbm4ce/bsXGgKAGNGJioSiBQdgbBq2CyngPj
UI2Px20keLKZTFnFfHdSMogw4QyrFKsLhavkA/AbBUZS538iPSSp0Eq9SlEi5hT2
PFYKVlhUNF1iCAM0LEIIF22V49YQw2c+/ab35+5YQah2lPMSAFcWMDlsXJGlDJ4g
4pg8zv1dMTwNKfTTaSJEa3JZMOAEOmbPNbo5XEykyG0=
`protect END_PROTECTED
