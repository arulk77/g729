`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
RPRXE9PT3aeNC96vwnbhYVGPcDMFeXii9RUHeWoXTrPi73Bn9oSWbU+j5eQP4ppT
J09Elc37LH2lpUOYAV3KDZXYY+XlRAp0xJ124kFEiDgFKQSdmIFvfxo58sR6CbpV
C0pVknQl7u85YSQ1OWwAFdKGGtTnyky1iOZTmDUlut57PWARZ0F5gWP3GYd57PON
Mq1D9y3zx7lRdORCE2sXTsACIQ/2axAsZAt8E3lju4aN9rNI/7OKj3VCDvApel5K
T7uRfKfdQxiz3UgwRK7b9Xm2Ca2d4yY/Fzv25wOS0qI+QxGpKriFz9kSFp1/FU9+
HgMQASX2stHPCnpS3m0bJ8MRBOdIa1ko+gejo1Z5Cakf70cuM4eqDsBk1kHZWyXM
/nxSdR8+85udZyMbgcfqcHY9JJ51cnVcR9EuBRvi8bLy8pPE/GBZAm/ujE1J/DlF
aqTMjNkdXVr8rQdziliNDac6DdLXKhTkU13gvUIrCT9GctqMnclZuIqTeJuxm2Ab
uaPHstXSSoWtwg9pF+fuDk02FVHWH9lHrOtPbAoeFwd3d/VqdzpwHTNg513TXPfW
khsvFixMvcJ2Eb8g7BZ/P+YyiaUh4qNEP66yd1KDzyeXHE4vOATwGyKcxnlx5ry4
Rfhl8ahP71Yw2DGXNgepZO8hEnXRwUEu2I0Y8Sz9Zq8ujSF66bSDeXiOXxNu0OKa
QM/xlgSFPe211rfoQYWedDqdDRtIlkO3N4ggQNwq8eXgY9X1WNERp+isZ+fqZTA+
0PLzmYAjrWNqg7tNivmku1DAz8ag6u7BgaKPE9qVKBXwp3WcXXOwO+Txx5WQYSgj
N6qC5dO5R658E5ejHMfQfpMw58Nt/pSpqOs0/Y2x/I6VCRH+tYbtJ/7FHl+UlXwD
BqP7NlbbR9v/d7S2pjvXkQpdctSwHTwoymKoMj76iU8OgrciSFv+ogorXiQZ+6Ik
lM09YSErnmbmnndShI58oDGyMHtAE3IDp/jIQuvSeUs=
`protect END_PROTECTED
