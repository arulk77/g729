`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
VN3cZiJB9f6xREOOK65F2lrlcHSb10efiABcFWR8kqCMFbnTBx/hOcp/vBUYcdyN
Z2SUcH5S+Etyj2R/pW5Nd3ephyORQEswPCVDdg0cZ+ioSDRnfAthyfD3y1IcSPIF
rXJ4u33FHNm30g18YqQdq5NUgtcbNtRe7awiD/0EWVHwmROlybWn0pdqhUuAcfag
Ms7mWb9yi3huMLBzRkUJ4w3XjLHJzZHJrq/jrJO+ZAcN+Kzf+IjIJJ6/a/r3WEHg
3Kt3UrXACVv76Jjlyo5urgoRlWmJ2icfLhJJzO6E4hyEyaIHMWNDzDoxNoKMADId
seqChPym+sg1zWStoVce/w==
`protect END_PROTECTED
