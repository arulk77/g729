`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOH1ImNto8QSBJSuwlF/f75BICSYMoNXJuAN+BHULmm7
1yxdk7YgiPAAHr1tz3cnfZANayiNm3XdiShv6SFrfke3dSmgLwuuxiuIl128IWr4
YnawS7YnSF84wj91z3Vm5WPVNgaKNGA58c397qdRHXSPeblPYMFCyh7eLKR9h2n4
x4TZmBKMHLNNfOj1I2OX2g==
`protect END_PROTECTED
