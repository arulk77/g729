`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLHfSEYpRwbI0N+6dKxfW2JNY4LisPMZEQkFOxLNRk5/
r5Jm7wDEIK7fxiBKuqgW/jT4Irs7fmGkMyY5OVfQ7FVxHLTnkJf9YPQPOZaliqAn
8Cx/HgghzffAzPmkfzL6d1JxYgzaej/eOlU6F8QsaGHjrx15Ok0yDIxRJt19WGKv
Xw1TW2DY1BjlyHs0pMarxEl1dJRLV+h9bKn53stclgwq5j2DgOUNiiCMmUWzKPgM
qXrw4Dij/TrY6AprqtxCRw==
`protect END_PROTECTED
