`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
xjzU7ifeNt1IFkxgZsaUfzZ3G6rx5nBEcLtOHb07gCra6pszSdR8NBiqpVwcek6w
CPfM0Ffq1f6f+EugkqGA8Al8wYq5zsTBwqFq7/EeBALiXT1HPOQhTq9MyqvJxKBw
oxHNzFMumXJeXg6tVmFXwZPpzfu7L7/1jqh0FHOqNKmTU+yWz21H/MdySaG45TMW
zibR4rEIVvUSS1Gg5ardUWP/QkMhA10sUTmiAMkdzEe8qc+RV/Z9ikCjPSypsf4o
UKl2c69q9y8WIpTvWwJATMc3y1INZSnQPxbEPlI3L+6ms80iC41f+JJsV5LadytP
Lgbf64qFdJbNSmEfSjBVMHqYqutPxOWPZ9rp8qYSe1A=
`protect END_PROTECTED
