`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
V2TAAKIG52j7kDjf9J4H+Jp0Hxz3mXbTtpZsIrCJxSBchKU7mDZl7uxvFfWqvVzu
1IL+nEzX7BJSFCWMn6RtylQkzzeb0TOYQBnON8+BJI/eBZ2VMpjMxm8lIRMQ+BgZ
y/0u6PAMijW1kY0Jp5Gw2U34PHo74z6lh2GxL2D0Ji2BdUqL3b3TfKiD2CjzPLDl
hCT6oDtwsvcSL0zfntFw41oWcXcWm8lM1djF/FMywjQ=
`protect END_PROTECTED
