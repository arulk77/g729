`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDASAnDUXU8kRuDEyAlrJpR9CSCCYxolmXmVtDBf/bUM6g
NzZijTd0ej4QD5vxv32XuI1DknH133HtLx27s8FHnWyMT2zzpWd2rpHLgJcBbP7d
Gesx6V1pG1XnAIXkM9Z7rzqkNEnyNeoP5d/pgI1D7jfihgpIAhhG11am2vJcSL3F
Dbz4oPQtshvh8EvRWEEO7oYHaBKxqkKorgJITRUZViziOk9IH2Mdwc/OeNXjiz8F
rkdYK903IFgQMwc0fmqrKQXU8L9wl2xyuv4MS1fO6Vr3IV2MzQrqUReTZQnCudrB
DTf/o84czTyq0eocpx/93yiiGJph09yG5h0fpD1xJifJcgzv60QEv5+3J5UhsQBt
Ew+7DXkvUf03dcUMlERy3wrlrCo81IJeqyaxL+BJF+5bup2VUo4aczcg+R5MVj0O
ZcFa1Wwqwxj5siAgqRYkT0ZNexQL82dDKqo3lkmIChnc7iLuJagPsG5I3LlMQ5vd
J8C4XDY+0bot7ITPVmYBlu+RGZ+L2qxxvbwOUmXW4pNk5ne9198BTSZ+nrxXOpqe
4BeCeaApPBTJkcJej+P/7Hx5n+rgfMxHGnyc1BP3uODDzFTg/kRcZ1NEvi7fwup0
ihEj8xErtYZeSuFXETL9q3U4JbGMZP+0B3VaOcZkS5t+wDbJCT+rXaDrxwzRIOC8
nq2EteKW2P/s+Ouetwk2wZNI3/PYoYYTIxAD6UtXQv60iQ+JYg2I2R+aNZ+0ZY//
Yk/XMAiSpzQrSdSMeeuSh8BkfTRVZnGx0Myqms1/Qd43r7GaeElbn70IKLAd+CJD
21AqwfIu146HPK07VnY0M3c+5ZJqM2owuDHlJqbhzqHvtKAOifSAR5rMXSZtJyon
p6wKgFTx/YOBNst2SiWgTtwfJiCexMapB2KN9/l79DHMv5QZBN0Vwv8XPtHNjXZI
+fGKToMgfukKPAys5DKUlNcQxuoW8QS21e31zuZOK/GP6xNqDJ67J7HcW9nqK+5u
oDE76Xs8kD6nZIWc53yEi+8mzXcj35KhAvOkUkLc0TM8kYMl941pytZzBdt3/kjN
zg1Sj8FMiiBr7uAGmqdyGJVbur/8xiiO/uwf6sUCFq23VC8NM2rS0UqyWkaJZrs4
vlN4GUWizpMoU5ROIB6T0EZg6MzmSAP5c5P2BgKsEUOBGS+uu8s6noovWVfIYMO2
Se0Aq3sVn7uCBYq1Vi+RyTpUd401Uq47+083X7U2JUBzaM0N82WXLsM4KApQ5RQt
TYuGw3je6+aHb9ctKhvYdVWv8UbNtqFHkdM4q6qBdDcPuzr3ix2qsDqz2Ecs6lKM
/Cytsy+lNbUyz1xolVzum4MxDiH8VFnglaMCeLxKgmFsqSktIGMRBqtSBxQFVbzV
SiiXmfBN95II+TFA1RspG70/FXJwR94Xc1eLb+bmS2MZQWgP3aeqImK3MZY2ibYx
1X2wpP4ekchrrpCoaFMmgRBN8uyd52dw+9SlGIFIlQGMMdA36hIlHJlDC4ZnVk8Z
02YNi0PjfDWSJ5rsX8Qpm1PmMSEvf/FmCue8DknSz6snSkdbwG72BRFU0eYDr5/o
cakrbhzY+FBuFXJ0KWpp7KdR5s6fAxcwuNLdAd6ctW5KxtPtV6+qHIRRATkyuhq9
DZev0qDwXNfbw2nhPphroA1R5SXH0tg90D+lhvX30gtJQ6rZWOu7JeZMNzMnsift
DMAbWvGbheWqVl73F4dD8+Yn4bH2i12zn/f3OwHXs8seIZh3jAdJqMKGdRk74NO2
GR3oOsJT+nxFqSt1I5v2C6rHTMGzV/8dAzP3xSLmRNlmOL25ZgJR48azzjPuAoQx
omCFmNhCWsWbnGfdiYdf8w==
`protect END_PROTECTED
