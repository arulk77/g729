`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
NfgAPjtD0CdBS6fMjvZdhaosaVqZDJBp6wCuTh9vCH4gf0oCmKFrxwYnAm8/pFs8
75Dg5P+TYZ5GthyIN+Nt1Qj3sKZXJwMH33KM8mRO1mN0uzwYeYy0BaT0mwnVdIGt
iyTaSN/5p85ET/lSP6xW+kwxsgZoMl+RIGiT5NhvgOW7wOWt16ipKdVl7vBiUOoj
oYEwTysKX5+w83DLpeQibuskx7fIGnlMH+z1p3yZYUNVzo9c9MwpqU/m5rcQkOQh
kQaSn3KydNspyOOYe6ejIM1WyNC2XqmPHOWb3sN1wuE7Pf34qmSiQI7c5+GVOEB0
d6g0z2iTKXctPbYVKDAeXDp0biOEHR+ZxW23i80sNwjK1ts6wPm4dHK7i35Fg012
MHsnLr0lqppiAdfvRmPbtaObZk4CbbelVJjRmZZgBtlorPKNjkv98A6y+iHw8s3a
TXsLV03nIz70LV+/Vdloxi2K7X3pblAxAZWPkhVFFK5/cJK9e0tWM0kKtJhZZ4T0
W80w/g9iRZUT4Jd0XRa8Czg4QGFxIEUxdIlk1L40BAEtuVc/L+l8kCkB48GYm5vn
8g5BbqLn9ytJ16HU6k0iJQ==
`protect END_PROTECTED
