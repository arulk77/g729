`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHLMLgMTZgwzR8LnPLqsbEUpSSEK84SylEGeyJvj3PIk
yA1q+DhhoE96VMom7AGf8XkHMb0b1r/avq8y9w4CSfInEu3y/THSyGXR6xJn8+Ko
9LkhMuLUKmd7ZhaseW4wi+tV+53MpMHp1TaWXGHozoM9GTfFLo6XU1iCJ9EkSXYM
9VQmbVDW7G+jJKZK/OT05f3oJvVjIw43rY7la3vbuk1q6EDt4CLVpHtilGr27JFa
`protect END_PROTECTED
