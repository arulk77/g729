library verilog;
use verilog.vl_types.all;
entity C_MUX_BUS_V4_0 is
    generic(
        C_AINIT_VAL     : string  := "";
        C_ENABLE_RLOCS  : integer := 1;
        C_HAS_ACLR      : integer := 0;
        C_HAS_AINIT     : integer := 0;
        C_HAS_ASET      : integer := 0;
        C_HAS_CE        : integer := 0;
        C_HAS_EN        : integer := 0;
        C_HAS_O         : integer := 0;
        C_HAS_Q         : integer := 1;
        C_HAS_SCLR      : integer := 1;
        C_HAS_SINIT     : integer := 0;
        C_HAS_SSET      : integer := 1;
        C_INPUTS        : integer := 2;
        C_LATENCY       : integer := 1;
        C_MUX_TYPE      : integer := 0;
        C_SEL_WIDTH     : integer := 1;
        C_SINIT_VAL     : string  := "";
        C_SYNC_ENABLE   : integer := 0;
        C_SYNC_PRIORITY : integer := 1;
        C_WIDTH         : integer := 2
    );
    port(
        MA              : in     vl_logic_vector;
        MB              : in     vl_logic_vector;
        MC              : in     vl_logic_vector;
        MD              : in     vl_logic_vector;
        ME              : in     vl_logic_vector;
        MF              : in     vl_logic_vector;
        MG              : in     vl_logic_vector;
        MH              : in     vl_logic_vector;
        MAA             : in     vl_logic_vector;
        MAB             : in     vl_logic_vector;
        MAC             : in     vl_logic_vector;
        MAD             : in     vl_logic_vector;
        MAE             : in     vl_logic_vector;
        MAF             : in     vl_logic_vector;
        MAG             : in     vl_logic_vector;
        MAH             : in     vl_logic_vector;
        MBA             : in     vl_logic_vector;
        MBB             : in     vl_logic_vector;
        MBC             : in     vl_logic_vector;
        MBD             : in     vl_logic_vector;
        MBE             : in     vl_logic_vector;
        MBF             : in     vl_logic_vector;
        MBG             : in     vl_logic_vector;
        MBH             : in     vl_logic_vector;
        MCA             : in     vl_logic_vector;
        MCB             : in     vl_logic_vector;
        MCC             : in     vl_logic_vector;
        MCD             : in     vl_logic_vector;
        MCE             : in     vl_logic_vector;
        MCF             : in     vl_logic_vector;
        MCG             : in     vl_logic_vector;
        MCH             : in     vl_logic_vector;
        S               : in     vl_logic_vector;
        CLK             : in     vl_logic;
        CE              : in     vl_logic;
        EN              : in     vl_logic;
        ACLR            : in     vl_logic;
        ASET            : in     vl_logic;
        AINIT           : in     vl_logic;
        SCLR            : in     vl_logic;
        SSET            : in     vl_logic;
        SINIT           : in     vl_logic;
        O               : out    vl_logic_vector;
        Q               : out    vl_logic_vector
    );
end C_MUX_BUS_V4_0;
