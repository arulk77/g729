`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Yu3rdfxH0sX9poQFeDMLDtc8YbTP6F0Pjut0pSOnhHDn5ltubBKEFEdezzEHC6KG
0oYI+7FHdSetGLkEULOMeeEB3PUZdMDpUeWHjUvgxZ9ychCdhtg82nIrBniEGmY3
iyJ6gXUz2y3RQXe9cgt3/HVq3UrAruMSzemVAAICTs5FljdI00gF7alfUIDgKukh
QUH/3747mwlERlWyAcqSuORLcWMKpslAvpSJlDZxkJhFcCmEaT/ZlcTKnXnnUfek
dq+qaZwe7bxaunrvMi/Kq2lltOdazJ2BCw2ReRxXbku1PZlFNnMt//zAlmC94pGb
kSVw1U0mBLl6KsafZjxrcG8YBYyLygg6+DJK+5hpEiyEIvytKqqMS7F1RwOCH7IN
+egYUYHBUGiPDhoCunaBw0rW/4F598uk9GdooWB5YjyLtTTj1iih1/UjgAwPLv2e
iO++0kdi6LVC3f9O3FjAcxfw9VBEI/O6MKUONQFiJ/QipJYAYe5jLJ5LwNK2xlBm
IIdvWCvnYHTIPeCs66TooIdxVnrKKsRuS2P+M0N2eGH7QkclXHiiga0M2c2pIDBI
hHnH2Fs9SfzsRl9tH51cu3C5ZBSL7mYiH6XY8+/ct10//BKLL72Ge320TwRw/wBK
H5NTZvYkeFWLuxY20QqvWcyvY2qAy5/iNDwQOrGpzVQg0q7Iw7T3HQlC+ArwmpDr
xxlG8WnCKobatz0i79dQGyy3wVIBMRLg/wwSal2XVamhWyL36yCErJLCIBXV0B0n
lrjRMGrSjnN1tIPmt7fIG+ILJgZYCLrxAhb9EcaE9APkUgNaCPkqjEHE7LrIBRSm
wxjmSKJcojvKVioQY2NontyuKNqrWfnONGMo61KPAqpvIt0xmdPZnR/p3KWcQQCh
/4DZaozhSHs3+DpJeA49MdXE1v2Druwg8dige/Ch4BUvlhrk+rH1cF904zdxkxp8
HQWlrhTt4FJ7A7x+KIhku/z8KZMsnQdZNW4i8RhhZDcF5hBEaU3Upbj6LZT/RsQ8
RTOtqxY1kAvHEnvcUU9dnTbvpoLiK+vewfNIpBpaPni5sdnrZSznhxYn/5U/i4dm
2c8LKgBzSUohZWWABDWePxM4upEvwQmyd++hr5yL4SeBsBt2SSYZuPW/UjyIFOq8
X7+KDVvFWmoL9u41c0+JhMOYOVMUj2o2A+w6vGOWOXEvjfQ/wNUwg3k1Nzoa1YtJ
rgw6KSuw06ghc3D0iwDLMK7/5Cx3XdxWyfxwiqIxf+/Kckfzes5ryvdYy5nkUMRe
kET4cuA/QXl0/fOZapqbtdMOB73ljOsDr5LYRerlYncJbgRqbQq4T43dNrZfzq8i
agK8dkJ6AnyFRZCYDEHb+o4O7FXbcHvbzzN8jsgxZm/KyvhqtthGa8M6TlSfQH3W
PWsOGnny9c2HJ2s0zhHmMhh3wml7GD3EtHSx6Z7gB8YViNCYZ+YDx4UXv6MgfPWZ
sUpJ7c9lSXeU7gv6Ylm+JgGEAoDk5bdNykElK9KyVOkMORI4yrXoGoFYlpKWhKg6
3wf7MY2eAE2zfr6Xilj933EOXrdlZTzvQdIpI5csRizblVGmLLEpV3I/xz6ZbKpj
TH40+dub82nzsHGB0rlJ3x8bXRC6t3Q5a28Hc8cftgf9nKwRLH7Jz6B7M4iNWbvK
ckar08D5RkRXLWFQo2/eAuPFcsHxyiZeUcpedIdRv94swXtqQPyNcbFv7WqU6DVq
D2pO/g1g4SuHBtUMz4cybX3mg1ZlloCfVHSsH2bLpM3rwIxEoZ31TOzLjXrmW5qA
CrG6wGLn7JG9reZXQQO2rPQwpgmhpETpBrjPX92m8gzBR5ENTX2iI6XH1oZlHfZi
0Sj+eDxYJMcT2TV/XKGnSqiT8asojsNR7IvEuZjFOXbZ1zPGOLCjbzo7F19Gv/8a
0YJP2AL/Ba6+JJT8ejh5gNBQTrsjMNuyGVcJlwGNC4Bh6nG5UOrJ+WCLLV99xvjb
0q2aAB7NH+iKULMajddr+MrLN7gZO6sVx5FU1iUxs5d8qj7sE1/kHLeSZ28A4bTr
UISdrCQUFrKSzCyqATZ6eIlLd3dXbNP3K8+mwXZa/mQcCONz5J4Y2giV4B8G7xGP
DFLBU4BgbrY+DOo1B3WtNhlChlyggm8rOgKNOMuiET5TTlICERg9XTP4Ae2QYIQK
KZzeUIkPPkUKGK/CTSURi5BfnG986mosHMPyqGNA96zUmcz0qv348WDLKsF9DyFS
sOUxdcNN1ba7su4i8u3MxkOF0F7LZEgaoqOvAJqjtiBm9O/egyVkcE6n4SHWNSPN
XV0cWyv8iWOL1I6CKWD/W7MmSdz8U2eCx0aOQtorYg8XQBrALMsyRZFL6ECgVH1K
LfTs6OgAnX/Gc5xLWHIKfjYT99WYIUEcmS7pKdm70726u772Xtcry2oyzhs8AK44
ruVyVr3eeNFeGwoLQsYKw1WuHvUsG+oGRBsDt/O3z3ZqEOF17+HYKKGbr4sf1UaJ
qGSPT3DmDUrY4c8Wm9KiTt0LBcMkcEPBpKPDPkFxmqxuAHwfJlkuIKa+UKkIyLAY
GKs5dZaJTkGkBEbDaQOPqDkzOUO39ei2iWDb8S8V9djw4nKxZKwV5LaqSdgZGRT3
WShCk5T2BZPIwXWQAc3+J73otoQ6jP2cq2a5hKfWqjrDYKGVNCAbm5eBZ57dmUjl
dc/oS35AEzdZBEnyn9/jic1ZHA0SeyI957leYVFEIT1lpu8xGPSjDnHi+pn4fxYn
QYWclIOWRhd3bDVlhO6MDOHahVfkZsmLZbuKaiU1jhgt7NoFOEFlxWwXtCrj8ye/
NzSlymajJaIhXAgbHKn5PXba5z7PB+Hk9we9SEgL1/j5iILP6i5uDOKNiIslPaM7
rY3+ZqrbbOHGo3ASUW75TEc/a/XtR5kd58S2faAk2qtFvyhZEqMBj5N1ovh0yifn
wY/q//SnCnlljI8TpON6c6SNh6Qgmdr88Pe5o+DWsGGasgmbcZpjHgZkUkzM9Eqe
8qFHuSaE83qVcfot2EMdcDLE0brUCDBqpz9IdLlfQWyspXmYUTT1UbRD2Mo2Q+FE
VqyPnVTnO7mAW3Tr+uYWUShrNkmHtnDj+DGe2n51EyojS/JaaGYWGwJ/ITDMwT5F
FCK356OfhomZon2zf9NoCgap8BzRakBYegkzeE6nUnV6Tahk3Wh4BhpJ7t7Dul44
WxIA5FIvKtoe46iaEgyiem3xwj2qXwrETnmN3n98C68HdQmuanXKzsgcYEBDgZGG
xDDK9VXIBnCx2W0sDlILvGUKKlUsWneUbHmr+m7326y75VaNIwIoA0srTmeGQs7j
KZJS/kVZX4taCD5De702MzLxm/3bL1SSNtrE1EnfzjEicIKR6B2/PiyHTIPVB4bu
VRhCnsg85+jaBaiKOwMctxBHefBWtn5qKBOpLvQkQLY2/uqNtz7i3QFao4WaXR7e
vfQZh9YUexLqj5Yb5iCeqD6eH+XTBfKRmmaYtO4t3b5uComEU0zUNV1a01LfYSVI
KJcptBSwnvnY05XvgofyhkRavw+Kb1L1XFpQZzy1FLCyP/JBo+csWkX3ylcc39Tb
E8FvuLh5Ff/4Ggy1rd+xn7HEy5Pm9bkdBIZbwlFRXDpwBWn3ssywL0I08AY1w1mc
MqOPfrMG3hlRy5jOPBq2+mu79eUAkRtlWea6s18DUTYdM5LrwJwokybXGGPGfgrC
/eepfwDrr8LXUylkTe4FJ4D4ZbR+l1Nil4B8iujs0Ozz2BKAOcXfFiNUZ7K1KXkY
lvaL/KIpfczN6yXCzt1UJBzsW8/I3msVTAesgynSDyw1GEML1Dbnwf6gHvAdpbsV
Y3bn3jOaBvW2dxwe0o/q5NIA9uZh2ETsgAkLVYaw0iEkJaiOs6iMKxaPL7xzoOzl
jDwHRIprwrWj9LaxPGEi4uS/BdUogSvuQsfV4qVUFBuNmKbRF/i8L0eMEJEUhydW
XHqAZJ0rVA/wU0GcE5APDb63GJB0obf2neDUEGZ4kLOFnCm0J8mtSDmt/lRwcPiN
FoQJhcowtKTyILyhh7g3trzs4D5GDhTlPmMKvrIfugdcK48/dr05rR3ofTGikHRt
nxPEhnR4phTJXGAyQkmBrbBTF2H7DTlVqfCBMtYEQ1xLyksapsJfEcT8ptaPMMMj
o+jEMXR1H9cAz2ZAm/22geJxYGDBGPihGtUJGRgDsULIgQb0M0Y75/YIfJrkyvgp
V9FZTKD1oHR6PMWvN7/283Fec1Kst1VDssSqVESq4/SWk1A2slZk248+sQ4c+jyP
DPwiqMTsAAFB7o4ti4qyrmUfHHtAAsmgOBvzldHWu/b5IWDqOs5C6XmIqf03Syto
S4wQaAVgWwyW9ij9WHzdic/aXDECS1OHBxrVn7tnBwrCr93I8q7nA64OSP1MaeHv
Ny/expyUjAjxPHbi0P6cURfiC3Q9CO0Cyscpz0Hq75jTGl+/gBE+/98ciE5MMFMs
9TaaeVGPUHWE7ec717qKdraZedbQEf7QmNDxkWgGnnSgJLsWPZM27j5Mgr2R4rPn
mio1xlcdJweuBZzP9z7Cx+Ni0LRAutXRm9HqzwEaQB7QI1fQTR1O2aDI7K2xsuC/
jEXQWubwdUAJBEe3h6tm6t0X08q1nXSOO5DJ6npktK0T6BYOug4JYqu10XV+N55C
Myu/SvWoBJz3J4CDFOIhcTQpLwMBa5PnNOV4cIzY0narQPuoxYGkr4ZbX34wUpTv
/dwMQNKafKFBklD2+PI8HWeyQPksJMUpgakYSOFPfROZ4tl+l03fglOm7qiAel62
bpwFbYHCgH50hz4Df6jJvQtUNljkIaV/BFs+m29A22jEOU1qY8mtB5xXUKJgRS2f
Inr3R6nYiUTskF7k5CAI/KGCVtlF9ZhKjrC2MuTwCoztDu3OalAXhYVGBeQ46HOD
fH78oYDq12D2oHsu94v6wbELBVQDdI7DLgcHX0LChKfGTGDwU3VJMEAQpJpg96no
2HLqYfRGK3xMWLadw24/LMYDhm+kKfnziNM/wAawiIwZToGDIzSYLzHK8928fkp4
LxWfxhWoBHKbvxyhyVqAT7NjQ6H+jh1E8PBUJ1htGkfyIwFKCakHgHoOmhOwvMLa
KAOaCZYWDQyLR573M1ngADV7l9nng9Og5tA15Isfov29P+R63cm3fzTNCmW/2WKb
W6U5nzmRc0F3goCqqh/Ke7mWwLAd+AVWfBm0s86GsAtLV8HGoiVxlVG4fKmNXzh0
iN8XCSFlv82Bkbxhm22cSWODZTxmFPTU6mIY7A66DiCpn0s1G633R5zebzwqQPK6
r3qsNG/QqeKMlNwBCznMNF9CSm5b2z938Z/MBHEIXMAGprzt+Ng5BM342HtZnWP4
a05zxfhmY3QfJBFgPEcZ5WlkO2GSz5BpZOrr/bbuKs6N0AeoBARcKkvfonSVYktH
gChJ3QB2HZwb408p/Sx+OVhBKWpH0U0yhAM4CedVOyJJWDku6IxKItQiPrZzAzG5
bUqGG4USkRd3+oXKhRPVXFrEEJo7Z4pKKDwglQylITPeT+ooXZqKqqytVdvsVSMH
uldiAqpgE01V4/yRMCvn4dWZ6/bOtTWDntR+H4+MYQV8GzK+P1ROAfkRm0+yJUq9
JxbtEuNiyyLJmIxJVFzqGtAyoPCwLmsqXkNgDaqOXT5cFA5a5DuKiKAxSroWWa+R
SWOpd9R4hpVg1XOc0IHvxps6K/kFArE1Po90t9d/aJN7/fmze7l7JoElRGnrUwwt
Ly1XDNrIXSHQfnAnWnHg1zBkIG39pw3jkkbG0tfiNj3JJRQsSXk+UKrAIWns/ewC
kv/nK3ALUwGMsQql6erUkLlC3RXLfn7jncHL7YOgD8cA33tV+5CUMcMNM9sCQ/60
B/1PygYYGGsRJ57fqrV1xIvGiNtonOr3VzRkHmHhpkc/nBEm6NdZQAItL/I/Ep8j
QyzlXKFr1lps0wIvaScT4EZei/sE7KYp/0kEiYr8uM3c9niB6Nnikj5FmNh87lAx
gNZFO+PzT8NGy/HkO5ldROCC3gQkcG+DD1GnOYSf47YYWhlMwZBty1d65tZPOaIt
0KjXkm0xBYWfUEXBJM672Gr60nJRK1fkErK/PW0JQ0oBVN1EP2KbSlOPCa/VzQ3G
VXYooNSqVWFnTnwA2c777m17psujcvcNxxPkwzOLxraHbc0hy9Xfg1C0nVF27Kva
VNZQdhSvMz7jEfYR9u7rGFpoAcs+yx3QvJnkFBrtx5veW8+0bblfi0CmBCIh9NgL
mlDU4ycs+UfmxD7+jCMAynbYXPwJPO7K2JeUnKNwkfFZ4fIfYPIE01D1PN4KhLtp
PfzqNt4sEwyBlSufyLKM8+Fkc/JBMdlX4B0Cd7Mucq0xMywyoCuqVuVHXmeBEo6I
S7CE9XH4B68DmDJ+PAhlENBQB5VlvZ+gWbXn3vTpvaqjS/Lq5WN8SFJL2tlgFoz3
111xeVOSP2qsY9eyLDgsYvgNVnlBLZ+2pUiu4YPioBlUOMdZ+HgcXyPx0uTNMhdL
VXHyQPZ6GFO6mUiRPHi6uW9483bdbN4Hpr86yQ95X1y+l79yIvosfcRrMDyiXPDS
5BpVQVO1Lp1LLuaVFbtpd7sopvIpb0YZV1sCwZAmvBFchxmBEti89u4FfPi2UP/o
RklT2aIxN0wJEw0f4awjQQC0CDCrbs4OWBDmHSF33EcuFSrs8UWM67Tq3i7rU6/X
OvUOrSiy34vhGuYVUXj94wrynVEu4R8cOgU33fPGrZO+NvQt+H43VpkzyO8+A/WM
kJnyxTaknNxEJfvB9SE9cmbOHR1S6dVD6SD8PUD0B9qrfJjAamDz/ysOrSJ1wc6/
H27yfvSVgVn5XJ6w9vWZ9IUeymuLOdacaN0U1vQLDPBJNKMRfmlZSdJzXIJlSLtp
EnTusBhZGGOtYHSJU0fUEo3nmQZSSqdJ1uAyg40tLXrBJF7P0/Ux2z/in1iLqV6U
7e9LpixVIrJrf5G+H5C9BXYf8HU2MIyNhq5J4JNdW86WRJAChBCJO0KxT/oATr7F
U9m0yhxD98Y2G/zYadvp8iaFOpoPYscEUIP55PXjAlro1QP/DFWOFUjYK3R1cPSY
GVrEo8Ma0TxQzr2PCA9CMlwsDO+aEjOLCJzPqwqOhwbwxBDgCWhiYAcXOGtNYSax
MkXY3CUn+WWidMEkh+iPexBmfU3z78SYu0X/kf1Mk+q53pbrg3zovEgTiewyH6fA
HKYMLHIOOwuMJxdaqDAh6sCCSmHGGPP/Xipi0aPQaRvJsW1jHmPZCuJd7OQ2cdW6
Cdq+Yq4J+gxHXH5QQUXotv3geKYrch+S1WFz19J9jjsNpD7YlaxqQjyHqFCav0MI
Uxi5X+VrOhnP1sU9sgtit6H0ImydzHB0BETiZgtyIpfmKbdOm9PHet/RNwnryrqj
bDM2trvC8NLsv0EIg8KhPR6hVFYNiigFGya6wpf0lqxCfznjbg+C4u//r7xyG412
UbRN+d+kv83FY0SF31BeLiMT6xZ3t5SMjmHDOiwex/x2sDhG1cNB9398Okv0f81+
BPwa0GS45KhsUNqGiHjRj7N6QxWE1FLCGXRsUeLCNHnT2cuTxGgrkyDRGexK/QIb
KEzzC7RriGU7slX/Fj1iB8W3j2+fvNC5MUz3IwCYBxMXeN5H8yjykn3H/J3g25l2
zY9zjrzT4OIhExax31JAfJFbN9DMudTyzEYYHwq6znrtWa5lWXSRAzLqygsAgV5g
FQyq985GRtr0ouQKIMFSRFqi/QVSb8JPG6D3j9m/UldYgeX6uSPx8L+F4qwFhett
ghIeOLKydM80ZognNSEPh5qIlpkZgFP3goxK1ITnz5P4tOxpkzVXapeh5GPIjSJe
zI+6zu/NZ/ELeRxd/s/CjH2+4NjXpm7l9lnGdKXyi+VXjdiw+fSc+GNfROaWO1lW
fr09J+lXleC4lYqFGvJJeG7e8r8M/VqKrGFABQfCkugcHPQI1883QSKsLwnI8A5y
NNPK6k+IwT8PW+JWuMmUZ9laWgMTvgJCUpx+LGI87K9zAaPdGciOo1SsKPqQkHra
QkRO7A+Uh2QgkfeF5FNDp2b2kcEoQ1/szdZyevcBDIcRY4Ihw2Bw2G390nL0slPY
LdeK2A5kTPvYvS4gUaAcH8vzsPvJGunKLhSQfgMSjpA4DElhxM4kw2CUoPMnx+Hd
LPURCiNE0B7dU/sCUU7WmsG/qjXDTqtHmFtBaw9feYqs8e1tOdunZ23ohhIog6Pa
Ys6XvC4q0mpeRs6x2mo6LKjzTKgeN9tcHXU1lF5RNYSLUIC7NrKRBpLrjA937eEM
ZlMEg9grJm7YajwlUhp5+9Rm3yfvYBmsYECUxnzlPv2sYPygg+V92jXr8KTlh/kS
ezV6Kb5ufDTx+RK1/IKKtxq/oFOYROlcMkUZVQd/KF/T81fIqDx4M24GvtK+mhSX
qF5qQ2OOoE0IMyNz9+8ja7rWKtXhzTPEPbSLSmHToXx92nwjFfvrXtB+FjlMy3Jr
OCSlQFlu+/zeNIHho1BNrrXVr3PCjD8kWzSqAE6lzLxtBbUv9ktnbJoNqREanCzt
QPEt9Pk30urrEtA9Q8jvJtl7mM8G/9YFfNMi0IK1YUujn3949D8yOZVhV1itLpkF
G4zRQdHNO8Q1iNT0mE6wjgijfFf7j/D95IU8mzYU940=
`protect END_PROTECTED
