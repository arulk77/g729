`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C8Y4H3FM/WJRTl+wtPNE0qMzkdWEsdSLca02yc6ykhRm
VK7F6vLBec4w3UR9QeOHSaKI7wMqB87M+ujx1ATB2yUSzkk5MuE3zn4m09VE8q3Z
3W3Iyp+lVdsN2hbx9W3F+T5n/vy0fCyJYvo8V8ZdtMiXQJYuLcHwK882LXzZlqgn
ur+ZTplDvsUi2+FdeVHGRYiLpTMGp9yEKo4/Ldayqxk1k34P0pT7DWTYSStraBeT
g+TnLZcdF13Bx66z9Efm2QiBC0dLwwdeDL513lfZDSTIURJ5nldAJkGzQ0AdCg1B
zKqBoFFrLbt7+Wb30/dfBYvc9iv4W53Ugr0XfVWr1APPD0ks0MXbx3mHM08RfGT2
3MWQzwdxDw5cUcJ1CiCxcjIWR13ZROI0D4vYDAMyo5tGnpb40jBJ9QH0RHou1sUf
ny2YqS8q/M68QnvVBhAFT0vYqdmpZL1+Esczksqw/einEhX6mLhetLRw6BxYNdfe
NWO5iordyIalNC8HlOgEkzWy5odNwXPngehwP1T58HupQc8RGkAGBP6bCL7atUbg
wOe+tiZv9hGXDNbGwXDtRI9I3r5662b3L3XOrckOcDBHOYgQ/U86l89wkw5s/llF
8tkLLzvWNXOLfhre5CP8sOfeVtUSK0WpVLDZYFrg/pkEJsbdNx2fr7DBAnvYLl9d
KD3kI9BhgaQn/do/A6zZmXahSl+M0PFFzYWcheNQLsOEx4yptQJDyyDs3PKYnclO
4SiC7TcKk6YwXZpcRR96zPi9I9YBZt6PW3rIz2eSraEgeIfbveV+RaWC0Y47ldWP
5M00ktPHDzQel0VktaaYW3+m+UapYKN3VaoTayBZvUMNELdx8Babgi9vd97X3Fb/
tDBRlYm9lyPgWJlAMLZyys/j4bVw9qjMhAaOIOMJ55O0HcObXO0PHBa/7UJPpffO
5zoJZrO1SjVIodP5FTbi750ZSin9y+zpVpCzj1ULNJxCXbJhTUrKHE/zxx5MHGuB
08ZXTupXqYqwSAhm8Sb5u6ViwUGRTT7NGCrDvqima8q2YIbYKqbKck+KH/bDf4dR
PxU1kL3VNSMeqfJil6SU2SCwEiML5nuSNo5Yt44QFc/PwtvwYJojA4Sjz3el1Iue
n093NB4iS9c6IDKuX2YIigMr6N8qavqUBqbhGpNtBKLy9Qqr8MppXmsJfx+KaPqF
gbIe03lXzRwh8UmfbEx8xwgbiD0G5NUs/H8KcJCF6iRwgb2wS7YEnUHi9VvrD1sU
GCPmj4PGHEzAlQJPJzDlxRzEpHeSDuCzmJVhVrAptiTqjyBlXTMcAJSC+Nd29l1k
U8BcpiwLPqqdM8vWAQhompXQxehw2+vJTqSO1SFG2egcecOA9FKN+N9M4cahE+N1
Q/iobRUehOsIJRNhP3JBz8mUhqIW5Jy95jIV1I4F1H/aLlST2soR4eVg6CsnZscM
Dh/0wyRPFArEDk4z2FSGBlImJ64IGa8m7EyO8t/6NDzPfrWqhduHyHry0l5dZAOZ
yRyItdytkndyhZQsD8dQk4P4E9TCEh4oEg7DdGdto8VFUbjqRHApIvbsprYHFo5i
QBKjuwiNC+cL36iUWgKr1/I5YQ6H1Lbil7eMWlJV1bHGck9en1qrjklgkDawD6M6
a35E4VYXZPRxXgWoLTTozebM83oovc/8VyIpzc5eEXW8TeEPWwTYVHKZlZ7ZCl7j
aH1B/SUG0PRl3rAFQYCtlm26zyjsW/XkdAiRQ+uog3+iP/MH458X7qxGym7EprL6
4Hd14QR1LJ1TcdFXtXr0DvwbQ4I+OlaA4VlxlnwABPRH70yuAQ+AtDS5lmoznk32
BgsiUcGBFqLpxs/BK6ngvepLwjbTNsLgWvVEyw7ySFMln2ix375vmxZ3CjdlDRG5
McDbNHzazfcve1sjDKWtD3p/qpF1mxWYp2NrKg0Eyz45YlwNu2qxDBV0bC2UrDmw
gnT28JZ9v1N9IB6jkYdJtYc7hUcJqTe8O3v94QPwOjS2LoQAGsuwhlggCxO2C03n
09v7YK4zwarJjcfFj95JYZsEfHHnA9UztPLHQS5yIGFdanlhmtV8xhG+O1DblaPy
CzzCsQyJRXRLurHlznWCQW6PlUSsvSlAXp1y22mVBGfVlhFHvASgYIuA5s+Tia3f
j2av4yCsDU9AvkDquqX6T/EEWXfoi7vrNBFvatuV7MxrVoybO+HHYG7hwhvj3g/p
F9AGTn8zZ4hABby0fIxg8VHsBdUF2Wsucl5tm/8/rZqlsleoyJWL2Zs8yumlUZiU
KOkjhLuB4p2/xhhwrGJG+WR5VuS6Y+/LVTOV+OOmYzV/ghYZrRwM75iiQ2L7tUsZ
VwmlJDLdypdhXBMf4r1mirQsc7aBbzCrfEtx2V8oe28JW89fD7IvEPHj/0gxfkKZ
iVrKSdTGUdAY5T0hiEBOHM7JAcsSSy76z188hNiVZE3s+C2R1TZ2W1XYk+86fxWa
VnZ/4r4Y/kBSUBnnE+2iRqi5/0lA6L9kmQc/BaTc3WYvVGvVMDDUfsdIzBTpO428
RpNiGgn/SG+sRUUJiCkx+QUmEibXBZEpPgo62DMwM/sSY9Lzg8bA2DS2G5R67f9J
dzM2sJ5EiSysf05J+HR+8LN+BBQxv2m663laNmsSrDo1qzTYbdRjvOKvWxfcAb0w
GilOBJzu4yX8eMvBvyI90xvcDgLECcRj7tQ+PTIZav794O1LICLZrBbGKyWvsQK9
C6UngVymS8QxJfl7Qp6Q/pcegIeNxtZWqVau0V2YAEi8FSJNDE8pro4GA2qv2m4I
XNQ7PRgq1n+qLbfY0FJKvpLRcImoaXpbmFH4F6vGqXxnkGNu036BnRz7xWUIYh32
kKhkoXEBaaSD3tf4o5gvEMcnkXgaVrNCoXzSZGlCQ4YRgzEJ9gjg/PyPwBbRLC0C
zw6+BQSlLPds5fhCso2A7PxV1HCmtK/XEmA2NxainTEGlWmV0yY+FdwyWiyoeitB
vbTZLy/HxLs1C44zE6fX+sHnkI5J05av081cbIWKqjy+Z1gHZlBtlyf8CoRM1bnt
MdhxFuTPkKuDzt14G2B9qsYUeVHAWBV3sGwUfFiF0xDSoojCJLnN2hjDypxW71qq
W1rjwxXwi55hz2QDCTzc0B+GNmufGFq/o70zD7vn7coKpywkR7GZEFC2cWqL1BA+
LkNmWcqhnpAL7mBp1qM7ax2BNYRwzCTY6+vQ1FjTjMGOXtXiOqoUb2qCyoCYKK6n
ElbsfQZmo7p+5ym4aNNNKAJkmfY8PJJT0E2d7LNgMvKpyvis5jaYEMOJeVHLWAsg
qunN8uZr6mW6iBIoBrT2qrm4/OjWJZkd7SEfETxSyotuFwn1tilBBxTMKxaIslxV
3GnICANEAefL+nj4ZtuGkyVjlOYuLsC1Qcr0S/5rVZIp1OmO/xaXtAXqjUbymhLH
5sjxuIxzZCwzkVRjxYRee2yyAdUUTcwRHVDIXhowpOhsMS/V24+c5ypxyp3oGD4/
HkBMeylcNzxFUrUhe0JvSWu5lHABTAz9cW6Kpi8T4+BOyGe2SB5QqtYBdCl6U8d2
A5QSv8v5TThOERYL7khVzBKNQDTGqZXt+nHm7Wp6VXyQrIT4wlb2G6Z3RjfZYr/M
mA/AnLYcnCryGIz5XpgmVy0U571u3OiX0+b+POOsixcOuUfh0rsDXK9uUxjgZA7B
gQ+5fKqGe7cEASCAMN0asK1sBbST+Iuo/JAqRWb8J/218PDJmRPRoeDujJdZ5yif
lL06mwErCqJ3QTjzWikOVhm4Ru/UuRzuMNHRmHmD0MAIHhaHx1kj67Xh9CldTxoy
u3UA7Rur+mOW4gHfjpSNihC55Rj4JkDcQB978pmUO334qRNKIROEhjPNW8vVBfj4
vonsI39V5UC+cjY/8PZtyIySUOLedUF0LHURW5a67nwANPWjiWBhr10ZaJ28rYRa
TWcLVG3SNj3HSDPVWu7I3uRL76WNBga+eYf0teZh6K5Qsxcp2LrgeSD2ZxNgiCmT
9Qvj7rwQlyZ3yCII22aS2PLqXrL9I8UtCs8EV161P2b5EDHOrg0MM+EewVyCRlHv
Kx+hllBtP/xDXRK/HXpPvRuryGZUe2stCUGO9VTPPJZJD4tkCC4aRs8ZUHLUFzF4
MkKx1I2NHsRyg2Fp/3jVyzS7MFt3FaQkFvk4Ukjq9sj8gFAtM5aPmMC0gSOP+F25
kIB+0zklVZMHls2QnO2Ex1s+8QBCFzRFDSWc7yF5qK6DTjtmT9h9S12jmYdIK8Ze
NsVhlugCEPBtFNUfb48ODIiEQyMS5fJRyT9+wyZJTqUN/kQF/jMsJMYWqA18ZfzQ
anezyusHYzE+7tFOlVTZjeG2Qk1iaUwUKygn2vlCO8ULxPlomBD9GKaLQiivlp8x
/nxl+BHi/j5o0m7sXCMao+8cTx3mvvaQPyLuWLYRumlq9Hcixj/F6sqzmoqqQpyF
WVcOBPauNMW5L7YIRd8l2n6n5emg9Rtzjp2akQdYEKCgQJfr3t5zXrLJccyM4Nw4
VX7SxSdN6Nk0DndClB656smnDWkdtKoaJUEIzkbkOUHqQGBDOV3FCVoUimq8Aciw
Y2rSHQfjByIayf6jddresFGCBlAxRlnKXB495FxReAlhdMVxPrVgoiN28FnnNRoH
SqiVHAExYFuCT+JpAisYR46IIR408zs4Kx5fPvjkzuYq8qGyDNF2yvEhf2FB1x8C
TSbyeJFTmAiO1PbSaq8iw0EZ480QMtRkv3ZGtLKzmX5LPIShACXD7KgEOyFp2M4u
L6AoekvWAJ9BC6FmYc7/ZowDgFbMualw2JUMbcDmYBUYwJzRHaTebXRkXW8t5OSi
qoUhjYZ/guSUK+HnhaRwk7sLH2rG4MSaol4iwuiY4s8tiYF2vgIudk2n/DiTD6xJ
s1xFyLfF2OcEz2Ij4Pf09hxqgA0fZKaJUZNgtF80z9ucqWBktJ8DapusKfQ0Oxpr
zacQ+fDROJOINvSw/06oQNsLBhfGW7UZLNJcXdcmP5arp5t//UgoA75RJPa7TEld
/EiI3FXSLHAjHCQ8P6AtNWp9jmwidCqy+jkmaAMNcsOViqE5FvbQovyzHuJ2qvY/
JEpA/ag+HWtCO0v6dJ5XzSnCchbfrWcR1jQtRcmR7c96ZKGx4QN3bCMQ0VTMCH0e
eBu9hXewZfU7FUEM3keNPjmYqrEHL/PiR8rKsHa8B6cCxfII/m3hqW5b68ZXwLBf
+4XDymkfQeaMR5UKTtvDDQ5FnZQkFCLaliTGM/AApLoDj3Yjo5YR3EmyqfSsWsHq
g75RVqALI7RXu7W5fpwT7HGBCirkjTUlK8wA2i1fjzOgJKLqOM2GYXJvteXBmskB
o24O6jbyHDd9Jie7JpWfboLIZtgOA4hJGSadvBF9X7Yel9NPclh4SU1nesCTg+n1
7oSZB92OvQVpzdEKftK2jEnKnxbYYuoUDlIz6B+xLxdFnt0qHdgRaFIxgvBcIMFJ
zMLsyE+Jrxs5UWX1FGU3Ck68638gVLZtrb9X4BYV3hgv+96wK96c7UBNRU1yK4yP
0eeKvRYfcO4TO3cbhZuX1LEhXV6NsmV2OYayn3ACRSGYZho0jYS+k4pUk5dxwYuu
UTj+c5U1j3f7VFFsD0I/y1gKCIIAy5LdS/xrzVc59us=
`protect END_PROTECTED
