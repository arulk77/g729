`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zBrJrsXYKJl19lVhw1hsEIn77qP2gUnjsl/fisO4/sm
o+rSmpTdkYbH6sUGdUuZRW/r13S6NpReCH4GZgf/JP2lDKxr7AbOOrkJYZ5KGnHF
VIy/As5x0boz8QUeRQBIYUG2J2Il8YSfccd4T02B7qIVmlBPDAnzCQK6IQ8avWab
T+2MKhFXJbYFnIIjxF0wg1ZiBgfVSZviev1HyTMcmotDd4arFrj5yGyVUeBn4Kby
8mQG2JUG9XxouTUWMMJcRlV3fc9G1kXQZ8skozNC4dfp0XQP7L7F2qb3HI69rtcR
e0OXnF6QVrf60EnBdh19NPw1CwpOHnIBBmgw5qPVYr8pGzOQGAt/yqEISmSa2QPe
eJDr4DJoQV4PHv6ZMb3DHA==
`protect END_PROTECTED
