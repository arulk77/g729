`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu419DOnrKpm3FUUnQlSu+4s1Kd+kDr9BLNzX+2tw2ei99
gxXjR8+hGg0nkdnA5dsKxgFSVqVMo8lev+c3aOd/PZjFpmjdLuq3cR2R8kC0FIQg
GGyeZ1R6lvmtECThHwyfuWG6Ufj5U0XP20Bt9Hiiv+li2mp1LoP3KyZgwFBXTV7l
LqOkzWXPd//Ml38ncHibrc+ppfL+E0OQ4Duf2bfJYL7QmqW7zPVrbQby5jRdiMz1
PI5zF+HnVh4/waruQQt9Z8MRfEumCKdIT85+YByRcYHc6BjdVNNiqVh9XO4t94YK
JVhjYMal6ulWvr8mlnZ4nhxIAbTIOdT/UFQgKH9Z+AO/gv0P1gJBoH6A5yV5jE51
N2HE4Lil+OiAZ2LXkWxYUQ==
`protect END_PROTECTED
