`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePbK9wtUIvbyDhGvH1UKhggI6coCsJcjvFjYfIN6zGiT
Ul46yvzDzSSnDkqmUET/GpkC8q4QWGF1AY/Nx+efqjAL+s3uegtV0ERBEfOdO6Vr
AmfPpXKjCt5KDu/SCc/RNSw56dCOk/RTz1EkV5kaR6RSSP1SWxfpUPG+QeUOxZeO
ZkwCtkoj+cxzGEflhPOSDVtNZxWfAdpkDE67cPeeykuEi0IMgJ5fJQzrz5uukNEq
QpTgw0plffg4Wgla86C2bmCwBnX+xjEFOWNgAxWrbD6O181qwGLX91RFsj6Dy7dD
rafe6iEMlOk1vS3ux0ZL1Hk88qs6C5G1HzYzvVXJ3ZW0jenWYZq4q5uHFXkKwRZI
dLAgNVL0f8a52oF6FQqq7I9fD7SPvfFhPeOtgA+13Uq8p1vlW5QF16SQu9u4uVHO
INfOPx4EK497XxBFjD7GheHh7dvkYgWhC3do6t27702bAtXv5rr1ybgjncrgNclh
`protect END_PROTECTED
