`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aSAjh4RJhUf7VEEdVwhCU88PIJHE0ostRSGf2X8Wywjs
9Lbhmlna1ZVRJU8W7eiTMNBa5TnktmGfiAfi7StC+nFvwJvxgHmtHe4SFP1AK0Ba
KGDHMUTdnvaoKGFx6sdRK62bHGceDCvafRUkIh4Hl7xOdkWhvaFlWEuWdGFz5oaA
Jvp/wUYm/Qu0yjJOAq0z1DerQPK8+1pB0dnv/vYrI6SrgK3oPfGLSRQ6o1CjbyGu
`protect END_PROTECTED
