`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN3e1taIKEQPk0KqcDiElfrdmyIQ7xlVYD6n7d+OLyb7
XMCHWEI+5SOiUCOk+gj26e639Dx4ZlLqLx0kdpKqQSa5QttS41isMzKVH06LvpqC
IuZBWcgOGZBf0give/2qMIUAHQFwjmqnUU3e8BiB7RpT//KJM112mdftDyiG+fO0
SmC1a5V0whRekOUTtn9zI3WC/8F6o6IJsXz8FkKaHbH+uiJyY95ws3Cl8uGPzTB3
fkxsJVrsDOPbCHVLNu57aTEUuaF3XEC8VmagAcxxYKPrBc2+Fc6Rxa2zbwRYgfJT
X+MCe6QYFaFKOMuMzLnKJw==
`protect END_PROTECTED
