`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLu7q/IjgQnWuAbYzk83811W/f+AOQI5tfBD3rF/QZVB
hN/LPz75JNGWm+S+ITen3GIDFjhCXPTjDgrauouSmJxE8ZoiChQmp1lndrguEh40
EwI+60YLP2MoUpuJBAK19Sr1nraEQWoCgr1iz13DS2mrZ59of/m4Ur7JtdulOU7H
gnb/ZLi0phSdhFmR8jF+CG3YkkcgJhkxeAUrV43yv5WKnGIorCUH9a2+gwC/xSaz
`protect END_PROTECTED
