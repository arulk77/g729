`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40U0cD3w8T3fFjXtSAEl3khEbe3oHNMUyRglqSqYbQUy
oSg0zpASm4kocanWlYAN2lNBIO0LKEd/Y/1qLXztGfoKI13sY/KP76S5/84F5Uom
5nMwA5cQK+BY+m14yJJa0rYv4CsVDrkRHEgIzkpytWL1uMOIMaS9c0DwpA4Vc7OK
gkplNokZZhpf9PEPsGKcEgvuqZecN39DQr0BGuupjK2yQWqgC+POE0rJ5HaqV7nU
cxzka/OhwfSbrIR7zoifAuUzrQljKFm/OPAWfEGAB4+JSukNcABxNvYMblLhAXff
f1HfAc2BqIymCx6Y0igllcTuyu7UrNPV6OqtOsMd6T2vFBgGGekmKYaaR3wkt7i8
dXsDgtYfsFGxPfFkQqM+ow==
`protect END_PROTECTED
