`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMr0MXQ+qVMKEEQFGwtKI1jIF4u7Qwepj47y8171vfQC
mP2s9RnO0nvyJYkdaHFdTIZtm/xGnxdT2dDPG2ux49OXqUO62aAFwgrmg1br8EKe
PbYUImaVe9yNBNKUbksYsi2w8zfCX36vPcLv7MiIIcig/8k5YqsPstSWIxBjMq39
HlEqAogKxSPRgwnp4VdYCQ==
`protect END_PROTECTED
