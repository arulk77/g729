`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
yZyd7WBz5DCoW+EVveXdLgd9/XyulOOjeBju08tS55Cq+gSapY1eSwdXb/dvtHEc
suiMUGFNedQ7YJtSmOzTh3i4Vj8QB+CF9zZ10zYqr5X/9qYxHZfyNaNdHZCv/QU/
A88LWjdEecyWld24wdTsRaHRqMC4RQlj1JA8n5ZiRV5wefCHT0oECMZeVfz5XnKu
SmLEv5Zd7bVd5OUVDTt2tQ83ce75nD2YWLzAz6TfMEwQc5cR1kKCXDFgh44cPx9Z
CjkVYV8CwDGJsZrhe174n9t2eQzEguR7wsfW/X7QG/xiUAfdDKX5jh2WSgV2lYjH
wV8j4H7mL+xLLyM9bGIbrjN7eZ2n2tr/2k5dRA2D2yhOVfNmwvAaHqJkNcTFBDQQ
L6OT01xUW+NGhh2bkl48FTnTWs+SwrZgvRICOIMeHkeN5WpQkvS3a5XCl/X2dMVP
gn0+9psE2/ilgYazE5KYLSAXSum12lxpmB7rW4Cojcte4iikVHAX2z0qvwvyMKT2
pLCTEucWdTOKCw7e4rFcQi4BHalBot9ENN5x9ppPPStWanBnCKn5zawm8utagiKI
0vG2+Y1NadoxgPFA9bLMt1u2EqlaRptBLnfkysFEygfV6an6L41plEsjOoCd0MDG
p+qHOfZsGzkHv7oPIbU+eq58XVB368LmJwXOs5+2ax0=
`protect END_PROTECTED
