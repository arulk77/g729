`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOQUgvdE7rejK2TVNId4i/r7m552UIWLMg/noJ2Ajb/X
vhwvbNhjfv5r1UQ9lDprq4K2CKzLTIPHvxKTl5mThL1lMCUVqPtrnzShCXoyw/mo
ZF1TGPXHIkJO5unSBlmMoUrW3H0ONc+z00Zlk4TL0xmnuCvv+N8e9xBL2+BwSFlX
NFtg3pV+yv8KMI+LfCL8Y9VkTFN0f5SDjc2qlZ++e6j5v06b6X4UxYRvt0PMMhgi
0yT+YeGDmoLtq4DIzJgpNZh3GTzaMDGSJDr2O+OKQX2RUfKBs2iHS3ry1tcwbA93
QnuYh7xjVol7zpQb2rB0gw8IuB4N7WKO1rQGMrcgSQAEV0DanaH+cEbQ/E2fiofL
ePviMp7ZKI4MDemyvkNRH1jXvBwkfoVnDh7u5m7Sbn6Yifv9VELR8NmsKtQ0vGsV
R++rT8omZOjKHUPYq7S41CTmf61n2FErwsXHO0UgstkXSEJC0tzH+6x16GLWn9a8
o5uykfXmpdXFAIQqCpWsXNlBgJDNO8bUf3zZQbBs8O4nEBVIfgG3AzRBtFOliz8q
8LCD2zoN+RtruFC1MkaRPCBWod2mMaBszrmQqWrvIU3zNS4Q/oDagpk69nZAGjWt
0dIr5FchdNlMOlI50LqZOMQx5jNEy+g1FathsEIf1oE1dofNlhXbEwEFFJNdIdE/
Hv/2rrmoIGSYne9ANXM3f0mobQCvJxRkAJO6T962PQ++NRuKzDc8zI3DaIWOs7q8
`protect END_PROTECTED
