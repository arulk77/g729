`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLTw3KNGs1/xkBzY6bqyJ2FAKpclVg0NoLB3HaPqMOh7
QYFnLlHPCUyRQNtHqXUvKTPcGRNhGHCMVhxlqB6+H+mPnMcM++LKR6uttSSkwJA3
11p/6L808QQKmGGn1pcfNQF6iOB310cuZToAGgvIa5c2Z+8aAWr2knupbdfvX7ya
ymhACMG49pyQVp0lN9asusmPCBYf+h2w8h3uywa0BQN532/ut1eLUOWR/jcJr6hR
Nr+vizxzLgmQgYJuozlGrPnqCJaJIR4+7KzUqYYSJYUD/0EIpKGw3pQ4BLtDsomP
YWywwjbrM3ny1C88qFYuapzexvdt4hOZRDoNCkyLBbWax+aJvG00GxNh/FQWitpT
/qox18Zp74ps5dfRApNEp5x7g941u0zK5yOJKsTXAiH/0bghf1vT916Q+8u4XOj5
l9i0yxTGuHc0AgUZrkZIjGWo8IzCO1AEnTgqD1DcF7hzCp6vwe+ApjdFgyTye9pI
U5W1GLkDDU2m8bqvKqGJT8hGYWwF2z/BXo5rKVv+6nInm5IALxB+tgpNkp7xdR38
nSrmIQTcOLRB42gJebjmqjmTb4t6XGDQzfaYpEytXKHoDNm/oehnDNYwHlExjJqt
dP0FPudRbd2eaQvfbLGYlp830fNbacPCAXeLJNM848JRNOR38A+ovsq037pO4RbZ
lZ0KRAE1+cxS+7PgFDKsCiBMcnkxuTKhZIsvMVDblU0QCWv9+a3Gt9N7J0Z3rYr8
MJiC3vMIz3o+pbSHehlKauSS18ynCGc83eKiWEmPwnP6Y1UqDBYcyEb7DO4F0bnN
uc1iqpyR5AD6qbMQT0SwnIavb3DJZx4FbVi0qM8eUZo=
`protect END_PROTECTED
