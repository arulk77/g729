`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAAvf80nZIv+k7PErTMzZFn5VRTqyZz8WCJYDz4pyPvE
2xvrO9zj7Iv/FV3FCrzh9fxZW1wuxLzVi2d02asDCKK9+mujvsZy+y93M5bcgLxq
74r6hYbz1/hh+xsf5So+0S3VAnOgs1biShkl7hG+4bF7+1q5Rj0XQ7Wkgd0Bmpht
/aQGc5T+j3+AwIIwUTzXUATnaFHyEPj8a3YxAUGMSm7tFbxDMtbzingV5PeIXYSg
pARZMypub8n8IXPKGCAohYwwyqJYyz4lVxN9EvtWLvIVx3lbrrfjtUBlAEyQKkkX
derZ5WpnrcAkMNzHxfixe4AXxi8jKX7SHIHq4su3mrR0+bUAHyc+s4tKysDV2zIv
duhMkYED/hc4ObEZ7voLxXCqvea7kvkBrJ7O0XusgZJV9ztEf0m6oLwiMLjELDAk
LTVGCeyxKVsmVkDgot9FlPZOp/2phAcZRkaTHf/sJmU=
`protect END_PROTECTED
