`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
5ofDvMbxglgRLDysNpBhAhS4ThK8za6ZrqBxGltv2B7kUDSqbD7XJamCg1dg9pDe
amCqX3zqjHnXkHCjwwivUtfw6nZIKzk53mCNlBnFI5b/cJ3fOMRYAbOKnYmUuEI2
z32fcCwYoZiRE4cW9qBENDCy70MxWOtV11CPrUhg4KggbOEH4iUUDpP4Lzi3Trdb
vZ8NnMKLeihl1S7zrUQA19t50fKDb1W5IQjvtJ6fyKTNDkQVGNCwdcZIZaARi1Y9
EhkOIvhc0UTnWk/CueyL3WDeDpY0niX0FnDHm1fiqhZaA9LNYbqSMbLxD6T5vdhD
fTjPLKAUp34xDDjBjQcX25PG0FzAWm942NFY6pqV5SA=
`protect END_PROTECTED
