`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveO+JQ0wZCxGdjqLhKIHKnU3FAavt7k6K7T3w+9MBpXKt
g8czs5rqrpl0QNXsdrkGs1PgwwxOMFYLbtvc+NlIRZKfOw+Mguj7MKrHzu0rTc/o
JheVr3FmJUc04Jrq7VS6VTuMccBz40fcGaCWJGL5xUjenOASRSu2xcn+EoM36cco
NZElv9p8q/w/Q5xsXRF6knQiSmQUnFULIw3x5s4zGhyIhQeUikFxitzNdNxSHzHM
PFOwVEg2qHEpmx6HQ0vzlf1xCZkqsOKxZBJqmBoiWW/iHNRvv5h5RnqJK3wyB/oo
be4fBVgEOkfdhIHmHrYv0Au544axNUc8eFWAyUwq2QjmJc8PDYNdaKYsSTXtP5jT
fJPvQA3qYplzAg+GKzIm8TH3DU8noNTreVIpCCywSh6xu4TuMOUpj9kt2p73WFrV
Ea8YmG2V0BTp1T58dB2I6ovsDq6O25UxjHe8vK8aoE9mMeEv/axcxsVgolRIalB1
m5rjPrb39redwqLKILBIQ46WbBE19ERnLfpGvX1IlXq6QczdXLoJKZnA2Q8RGkt2
7fiWariKBoOw//J2WBaZm24NoiJPH/cIKrEDAaAXQ4y3d5ThI8q8JIc/cHCx3rhG
b94YlMjEpsHnavsQ0HmkXOpNMbA6ImcM6PP6As7hQTiT7IJMREBcUgeA2qOVbdcU
`protect END_PROTECTED
