`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveA8QlO9hJ4V2dOOhmOVv0x7d+YELaBz+QUnNaS/APeIJ
TUeywO0sH9cWt981QsdcVdAhwkjmU8RRIu7e+iFEhim/JouOpL+SDoUtM5M3ZU/J
b6P7VRZO3c3yYJClNmAYAXlc5k/XUX7eE62xc6CQLJ9a3/fCBULBdWVOfXc+kGNL
bVT8/hSLPc5g2gYPQjOamw==
`protect END_PROTECTED
