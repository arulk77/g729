`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLalvN2GxqJrLDQF41smSHQLyygv0tCyTthAYAwEePFb
YIi3mkDHF0Qc8h6Xnuydfxm29md7GccMD+sfm+LVkLO4r/BTVjd36sQmAahEtbJG
eDxkBeMtlseDRmLWQzX9a3l9dfr19jxy2/aWiVMU6TKlE+egQIkdmRhYPogiwc3L
Nm3k4UPCt3gFGbEO8fHtDA0qmRt2u8DTloyj82D/MTeZFODece6oEw4YkzSG8bpD
+0FjuLyOOa0kI1uVJT1s4mG4tRsOW292K0IOBKdv25LxgmzBTdiUR6eCsBaUnQmF
xelBdhPnpD9eJcgOscILChPdmnjZlncZtCXpk0MX6NEjYJMzZxpN6pyrclSXcO39
YR8f7ZWfqUOoh12vsehLtCXBYBPDCncoc0KdUK1dLUbk/qplM0wOpezNW+kJeLvt
QmFZC2Dodg735HV2JcQa+nVIKNU/utWgmUWWc+OhoiM45Wk8iQzNnvJl9h1FrllV
Gcsb35r/yLSW8o2oGlZNhQ==
`protect END_PROTECTED
