`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
9xJL8kBl6IDt1Bw6vRNbaoLze34K/G4htL3lDvzU1tu0GUz4oerW5piTfAjtn8Yo
YnA2NdbDZCvZ+EGpGpwMKc/eU2mifDDr6oORiqLzoDaSQ61nz9LtrtamVWAnMydT
Xi4Co9b3DPd6H3v9KxiTliv1wZotIyp/tpcOht8WFGJsuydb5IMlak8BZ/hnwVP5
rhOU3EFfHarXDBwAPfA4bheVNyQfXwMymf6/RZp53oXliDW2lcF3ipzsJXITVg88
`protect END_PROTECTED
