`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN5Gpk3ETORYm9eMB/MT4VxzNTKlJ1A4ZTmGFuIU/f51O
r7/pTRnTou9nPv4xKoRqCLdLplY+eGCpBqzL9HU3VgGgyNCwG9fLQPypSsxlCQ9l
o4uIlPQFGSajgCKiWKlk/q43uiDenbBmZMjCdGWQ+WuuFQWCW/d6yhXr5fo/ld/E
6s7+OTkAc8fnEHaBmpgjhCzys6YCKD+NSfhliXQXL6md14ha1q50kLtfNKum7GfX
xLwneKJMFGTUG4DAir4V6S28ffmcVVc26/N5X30T24Ieflns02Lb2fvRM8GYV5L9
EwMXMicJqWju+iqb/ftZeLF37D+AVD8P2jApTPylLvzNDzdhxW2qiCPg0nTNBo2k
W/ZZhF3kFow6H3W2tUowPl+wvl+MivaWKTDfGfCsJzkMZJwdADB1mn2xv+TNEG6e
6BQoB/9dajnWSHuAnJuml12IxKzeYNj0gmss+AhZl0NsbMznQ3TEpAwE0jGP8ryi
h5Noq25Uxn3//ewmaULZkDyKSxL+WOGFiEIz1TMqWSDNh6XwnsBJagoC065Lstao
L4Yiyw1/5EYvVyiOJHytFe7KocyMBGTXymsg2NWQUJMrObTU2SjQdLPlYmEJA9s4
rrQlL3V93Z7zAcO2h1VKFbCuVb/b+X+14JaiSnKVUKTbkWa41XBd0J15ngU78vxl
P7uApI8DnENdZP6HOrXGRuS+BUpwxh1b6kpe7ub7DrE=
`protect END_PROTECTED
