`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJxKeDrNBqH1PgbEcF6rLrP7R7Wn2EBwRQ3VKiuVFvfj
gxAb/K2mooyJigQQN2/ABXhloJvnnpOfyp6PLVQjQiQqtwLdIw3km75mjEeDUk1m
+c+rNLF+c8ehjFEpRSahd8IsJvfCubWKDKODKWv+o9Nf3nGhuaSNg9w9fR7R6Jo4
GOKwyRL5VW2Ppj/VBP+hg4TmtNFbuEdYTEoe2SssEQ0xxClvG1mwXcNOwwsaD3Rp
yzu1WX64r2bg0aackTNN7g==
`protect END_PROTECTED
