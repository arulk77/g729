`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/IFjDDQENj33FoFZCHoezwTx4UuubAUQlrv4cTacyb0
w54qIuXqsY8OMl4PLBg13npb4VAIy12d8QgZEAyh9u3CzdQHs8L+i8hJNbUJg46U
JuoDuha7tf1zKiRTj75uuHIWLxQsEEc9AyEaJ4AyN8r+1ZtUM2Ii34sgYBelp4Vd
PGztlzP7WJJKrd8YJ4wi1cEGAbwlHo7M12bn+4/mJ/4jVI1G0LrbqltQjhx1BvMt
ryVnJAsGVkHy7y8jd+AcPRXTKpiA93sVnBgoRXKof6pkcX23Brk3S5TXTFIwAj7P
6zxcflZ9Kj8+4sPwDrkjWGXphe9eNAS0x99STY9i9i9z7HmWQHFiCt/tzSn26ZOU
U5h1sY6rwsyzRegKwcrCgg==
`protect END_PROTECTED
