`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4jahNb0brbuV/RfqVptNMcfoOp7zM0O02uwkcXuRp3e77jdCgtiYSORvBts0BRq6
xrRf+5U6ZFbqsyE9T69OpHMplidMoJ/qroK1B9+A2ekPHprtt+2qeXVq86/pcD9r
RDMFc7Vuy2huDIOHLSdpx4fHmeOnKIxw51yTRINs5zLBkBbFerFg4sKsyx8bpNIy
L0aoKrDKjNqybhk8GHW+/W8wD7u1f5WwgNTFijGIzjcox4lnp2ixyRIc7xO65dnY
9GXBzCjW3MNp7/WeRvuEdXytSypTw46zo8NbwEEAxOZLxRszDgQDFfFE+ATFY0bm
eSPwwLt7IH0jp40sDftyIgw7AHEifUtsU5OCm9AELEg=
`protect END_PROTECTED
