`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCtBqnAzKI7w2upBbFlu+wpt93DvjRkFhKP1iEhAt+qT
fa4/5j5XxDff+DejNhlFxhAN+9Zv2rar2VoPZKniYPwUhdH8qYLzX6AbozI1n2va
bBJdw2ivCsfYmkRSJx1f/UCSc0TUa6UKGBBFJeFTv9yh9gkh+5Z/drZoVJCziOrl
P2XO72HoHqGs1skS63fyJR6n9/VsT1JuNJO5duTCtrHG5+WIrBOn+RGfYLBjY675
Rd3DIngWDLh74h/3VZrD1dsC0rnEWlqtYZShY9BWbsJoJtFEBLverX+jNRg97Z2J
NJ5r2NesW43eViDetMm2vW6Q9OWv0dGJFMGzduaoSct9rkoRzh5HoyxRSVf/38uz
kyEM97Lxh7UKEr9KERg5XglyOgjMkOPMCT8JqXVeJZe/WOIQONvBBEGbC8bN6AE4
4yhOb0Ajx6hFOcpJxrXRW1lAYnUT/JoR20OBgAjTf+UN5c+qwEAd9mT+EyhEwrHV
58eubGptzn1O2diys9nNdL2ViMG8IBAQTFMLi31varCZEv643vpfQKRo2vkhPzhW
lO6DokjWAxW1Ry8yuXEfLvwNeM1L9Imc3rHENGGjb9zD0hthiVJANcz7O+SCy7Oa
tTWvyM/cyNtDeifHL1glwvUZzofFgr9jEVQP+L6uCv/RRGU1Rx1ocu5GFDrc2oqv
`protect END_PROTECTED
