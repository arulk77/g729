`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
zSi1rF9cyJ8dSjFTxZwm/SDthdOb56ayiSO/N4XUEFvSseZFpi+vZ6kJEFv1/KOs
k+Z+xR4OjsQGV0s3TwdztM9Eh9y69NGdDGY5vFZN2AYNX0S3+AantmwMdB+7D/lI
85LnEu2pj3QBEo46TZ6rBkuVzUwZZDV7fpHWEWcQezhIsEFhe+JhK/mqximbu5Df
ef/NbqqEkmIFqCa/KZrV8Dtr8IGWtZFgU+RghkPANyPT2cRhAdQexxIlhU4hWvJr
`protect END_PROTECTED
