`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveETXzWQCo/h/TBYXjmDX9SO0hAxHuQFwPq6J/CLKZ0p+
D0CYb0pzlynGZwDFAy9SqRE6dw5rctEW+nyYZbPt3aZRS704vD/6IGgqqaSb3yRN
6GuJnEdUAGC+cRsDEKXF+xvjSdkGbey4Mfb9JYYoxB1ClnHJiC98QLhhJ2fXUpeN
R+pjM7AjGAyOAM3rhAiq5Z04RdS7ed517Vkre8IYWsxO8dl9MaS2SQNNf8wXZb+q
U0F+IQVoGcWgEUNkfSjjAfgJ753Ar/bsa/FQMrZFvEtQfWD4aDiVb6MBTbnjED1q
SFlT43626EUxWhPeX46713y4JQsz6/WHs6CDBccTevk2vMNYFYzGPr7geOeWCTsm
AaIwREP+Ngw13Sj7J3mtYe8L2dFp/RoMfr3LkClRP609W6s2IMZ7pg6DFwo2MzTi
8cIz/HIBjDBwOH+IBUccYWGIkudLL8wUaFiGBDyV+VurO1azFuIk6HXIE/jaGzg6
sS1N9XFVT4q8bsZoFgQj1g==
`protect END_PROTECTED
