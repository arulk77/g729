`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIYXQrN+oerf6OzyvcyXjbcl6YooSPMFW27g8KdIjh0/
2d9BbGcdWmG9cM/leEYnJ1fdwRZok8nOSI1XHFeAC0TYz5T/VMrNXULg3DNVojU9
vkr+NATRJenBIXac+g8RJVRw4laISvE3aCGuUgq45HgmZ4kKHWHjDXfezXhs86P0
9/BFKmbWa0rsKFEI1uQXzA==
`protect END_PROTECTED
