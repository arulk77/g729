`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
W52by5FksJUdhgHLv4Ym9GsJPJkPb298G/KrE+AWJZc3vr22DcL12OrSQFmJrOLu
aitA3X+xz2/2M/fccNZCFH+WFbxXmYdQJE/oHFZeWUYBkNAdN8Ft9Dcv0mDL1uU9
SD/hnqrd6N6EjciVs2HRTRnP4uRQFq+r0BV1vCBk3+Inf8fv1vuEGNMx4w/JezOF
VCq7kP+DZ9yLc5fFv4qS4BvEw971hti1IGPWczEpX89flUMSO+wz2i/7t11QVXWd
2JDDVWm1fUYHVjR7e0k3PTvJd05lAC7xOdISfNYQ+8Am5/CMBetKbEYWCYCKI54T
jpFkzgMGDW7apNAMYkue6oPIspjFjgj0TeLuLxotbYbcChkep2fu1wVfGcZPxJzL
AbfrNeQ85iyT3QAmmhNxMDpgmFbMQM5wTCcRLd1pLII=
`protect END_PROTECTED
