`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
jPVr2hMI/b6dL3J35U5J0Ua810HarEMrj4ykfne4KKUU5yXlEQ834D1i+7vNTmWm
M7LMnF+JHSWJJ/EcrSBL+PUkfWwPikJV7vMok0h0hUTs76xqyWNGZXghejbeksMV
0+9BJdRgEWevwvKq3W1f2HmjdR9GK62nZYBuMnxEHdeJfRVRcb4LtI2w1ImpIxYH
8VNDG5ZMbMiCEHJNXrLYgqhCOjHliJ0ZAaVu4GTuzwBpf71TyaC+Rh1oYTRp9r3Z
caUrnWxi2LC/OnE5qAtU+rBmYKGE2woD8jSlerAIrdY=
`protect END_PROTECTED
