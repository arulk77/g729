`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN1HWBFmtyVMr5R5eCl5v5XH4VlEYjMmmi3MfnFtvnw3
aKVuG5FVsjdgPxmz663CqxIt2laNxYQ0AcZIDyq6SVUJwl7LrXW/Bv4fH3YQb6L7
GB2qryESL5i8bRxwz95pbQK7h3166/J5gAEKQ+NpZj7DATzPJ1PppeAfelBPihSI
U+12tcLBf9aVaEFupBBgpw==
`protect END_PROTECTED
