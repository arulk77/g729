`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCKXIDAutzcq4C0miVVizxQwyyaTJNUN7NhqoaJHiw9l
/9EDzWsDIbvrA3PK9dG+XCcoct7ZgA69AhxaabZcvsbGXUbBOUSSSDUqjPQ/rMRC
v8Eyd3zbE0qpPtmZ3ExFQB+cJGZovpxZIekNp65FSzmmtjlAtWUM6Vqxii1atSQ3
`protect END_PROTECTED
