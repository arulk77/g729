`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JS6Ee/OUguv3S0KjECptSNrwgCCh+A9IOedOp2MlUku/PsgHBfG0c66mfkzBQXnh
MbiZ6OqzpUSsQxxh9OW8RqBf+qSLiS0hW734np6VM81L+5v5BCULC6uMNdPZaZKp
uUCG4XRvJakVJnPJhnAKLK9SmlIfNNS/l6yk6GMRhFE5Y7gmWfS0tRxiNxzXJECO
oSjJ3GgrzjopJnL2PUZU5dAEz/3xupsU/DSsSUJb/hi9b17cjDypm1ibqtntCjH3
`protect END_PROTECTED
