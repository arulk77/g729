`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
N1C3GKhX5DPT8Chj+mgrLFIauuoa5/g7zoQ/xOdl4luKpShNyLGFk6Gv2EzOaXRo
Ij7lFNl1EJIqltLFlsKQvuS75aSmeaZxoPdvd1Y0QBdEZC572q2S+JsfAcyf3qwj
UnuZRkt2FwRpIxvKKR1TdopwXWB7V31FkzwieWdfyaT53MkSsaHaFWe6NJ0t6SM8
de/+PKRV1miDcdnfEaLC3X9pw1IciB50MFAojUP9FIxO1D6/kRpFgACtpJSA6kl3
cnIPUCulMzn1bGEFWYGTul3sIZu1hjlgVlipTUNkg24=
`protect END_PROTECTED
