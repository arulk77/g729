`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yl+HPJkvdeGIBduwDvFcIxYpe8Qoa2FJsCcJ6BJvGPj
cLf3gR1cQjrTdV7eRJ0HYfLpULX+nBBGW1bvTBvzEQLBV2WIL8QYlX36J9PtbtWC
cF7bOzV0/SDVi3tqyk5dsxVdgxddur13c/TkuT/hpTgLVoqd5P8DkjuvC2z5crNI
uHSjFo8SVEZpOjB9y1dZf1AW9Yllrg/jw4BZy+0GdmGIVUysBaWlD2jk1WOjHVbf
+/xhJRLpPlhkxDf2uhSmOt8MgatuRBSvz8MwxZTQmHfsENCog7zTXcJTWIlk5ARz
B9om9rKqPkntzI7VyI74/mS04g3pdsF2QQfd5089EwejG6L7GXgAPlgbptYlYz6j
qLcJhiCPNslOapDqrsDg8y/DlQoTkqyZ85sh+c4fMT/PTZwW57YoBROcY0RFsfXJ
P1s9g5NdvZW3gJbUvUV9sw==
`protect END_PROTECTED
