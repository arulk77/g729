`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42HOkRYrQEtW6eUhT+vpTDzY9tgVxFO/WGbrnf9+rxNt
x/jLCm5okBb91FxzlInsoF5Ol83hh4B9vJxgjeENqK3n8vv5oDcjgbX8cVAt0efm
bVOVsMIBZhDywoXKkv8fQfF9cqXhcFs+N70zbPOPcyuzdJkSsArLZBEmdFGY9ire
H2ffR2nSvcG8s8nyL8cw+g0qlBRbJWB9t1JYJMtE4WduD6dKB7oB4Hg9hxhwMl9E
p2+cJDvX63YCbBq3zs1buNJRBbrBYG/sEiJUDMRcdgBAu7quusMHmTmnbRvfIM96
C52xyiF9odLBTwmb9oPy1g==
`protect END_PROTECTED
