`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveArPQqkgAlCeeuusdqftUIf3GfeP0aPdpGaENcaGeYIL
hSurK9rkCE/i99rHx2kCE5dRa48dGQLzyPnq9C5Ns+z74qtwJFIPOhmbqD3ovLuP
QNjvlqurTS798y0X4s3zuWwUCevEN7sJbjWYtXQuDtGdpyKXXc49YvtEYEqjE3ok
uPxI4jw8F1YjVpZTyzRcAhHtITZC7FYrZ5bFhGfE8R4OZSZq1NTzu6RLuxZwVwRi
krM/vDfgHnPKZANjGcA8kA==
`protect END_PROTECTED
