`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveO5NLvBG0JAlYANr8R2H8UobfUWFF4+VHoXGAXHF0R4w
s1uugI/UoUNtz/3a1q3GN1AOcONqpA8pp1+Yc61wzLyRQ0ivlM9k4PTZj+CrKaL0
nYkwEIpqJCyj0U7qB1nyzu5UMt7k/SnI+IhllGjoHFpkvDE+iGLk6+k8RaNJ825o
m/ySJv/PpVQSucJprZ8uQrhG4OAFOY3d4sBmeqEp96wxDVKtSneDeDUgH6FZ4ZvW
`protect END_PROTECTED
