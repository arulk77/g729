`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QltYdGPWBScWdGVTC0DjLak2PnEnrEUuYX1w7gzgiYTp41EEl+HhC8BgPUKYdZ7u
ygo7Uwm0oOI0t2dsTc3Aip3Xr78Vun9GhLuGo3Xt2xDnEghpfdIg6IYhGtzZ5YEe
`protect END_PROTECTED
