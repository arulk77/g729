`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
n8a8fEgwVsk4XE3MbucQy6+244Kf21XJJNel0pEttjH/UDZGOoMDSWu58MqJScBW
VyTi473CSeb4obTkmNafwovh0zJFvayw0SEdRWhmje4va7kiFhf9zKO7mTbrsTok
Wc1okhgpacTRBIVx16wG9qGPsHsyaMJgt0jVL1BE4YWNnN6UV13zZrrLw5rd+GON
9hFjt7wH9QYctbmzQNjnJYqNSmjXWPTbdPWx4g3IFadGeP4I8UyKL7sE1Lcv5VLw
2YTe8xn4rJ9wZz/vYXz1c7M2JBaHEKVjapX72rACiAXZb5Xll3M+iYRl/yIpqgkO
xaCPJExkuRTRnqQF8gqxVPzfNkOODfInTpl9tXq7Atg=
`protect END_PROTECTED
