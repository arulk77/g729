`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNal8yDHyUINs3S9Gfk2+NwD4gJQIXbMR3R7mV3AacWo
LFYQGg8Z5OEBwqfrxh1T1TWMAKnwxF87mNffoxcQjM16P2RrYdygWHLu8Jr4n4ja
A3FTSIivuFMpOge5ua3Fx4Zdbel4THg9Z/2rW5T8zE25VXLUr8TrpSXLSOL0CB8g
7ZQTiYYGT1mHseNpltF4QxXqTHpXODsT+8NBg2IKg0WJj7WLAs2m6FJghEtUiSgO
H4TFFoxw1QX9/02CiagY2j9MP54DNuqvaMVToxr9y0++bUgi308cSFyk0C7ffenK
tdEDly3gqC78UUACBCIvTNX4xOYRe0rJW+vRq1D+QaEoKpmcWTOtnC5rwbodxaHq
2a5aDdTBOUFJYjZzB5si87gkcqdLXcxW3KU2aN8AFK9OO0zsq+jvlIuDcSzx5L0+
wUcmlZtiumxnCDelOW2+wJMrCgrMFrPDI9eRI2SzNcYGpVK/sP1GCITvZeYYa+M7
`protect END_PROTECTED
