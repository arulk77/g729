`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44uUYLKOkK3qjK31dnlDyqFAi3rT1qF6JfpDP7FWSJ4a
F4srLtZ9oVhvM1sFCb1ZPZBioZTVYfh/922CH9dN4B6Ah2slQHM77kZ1kYaaU9CH
4ka+/2yfaFFolWRY6/XvQyxK47ubBnuFiHAADVp5fAUGiHub+BOQChu2/YcW6kfJ
i8W6O239e+YhqkOZGSIc374+/+9/sXQfMNP9qXb/QsdDU3ZbI93DKKQSHRQHu2Cm
PnHANmDmVVOOpjEbkNnu/au4YyWGvJsHTe2/EBPE3gKzMm+7btaaj48JqZxIbvqO
c4E+4N0EBUUW8OIWhtT3KyvG/MT4WzGIRuHnXuDRbqdQOGp1CS+9ep0l637cLbYI
DtpYntXjewklBqOWhOXEfQ==
`protect END_PROTECTED
