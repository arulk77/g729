`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDlwBrlijcHAqaP9w3fdWYpVEN1oM7clGI94ueYCe1HP
iDusNL+mlEK+A0fy48XoU3J3c03sjDkYEc9+twVhJUywGYrFu9fHUfhZvZjHFKsw
cH0dT1Y+b4m63pfs9aY5SxAal7ADKZ5DcBmP8CGpexp+cS5EQoje5OAxm9Qbnv7q
+84afzUmay5ejPBjWFkFi51G427atzp0qvP5Y2kboJH6dNql9Qeatg8Qca21nrSF
`protect END_PROTECTED
