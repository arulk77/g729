`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
9u8w5HBbAvrKq8z1du7XGgJ5ZG4+wLBJBTkedO0dy9MPPUINulLuOG6O0hHrsezB
1I5mydxhU5joVCpyMsNPZOjeVj5rDEpTsI07s0bpFGNzdlsC+c2h7xUx7ziIt809
bkWNPSgk+5vHmg1Eb/soo0zseXCkpjrbe+2VmDIYAwJuG9RKQixvohnLXCvHbxvD
RmbjqoPowhaMehaRLkA1WUAusT66id/E+z5Q21KfhgmO0lV+1W02wlbyjVkhEIvj
h0tVO9n2CTo8bPIZniATZ6RbeNVXaPlSN+cAPR2ZkTcQ8quyopkerB7O9ZFqwpy0
2UgIhOhXkI9oNuC0B0LylNyOhUthmIifv0k94hppxnB/4AhVdGKEGeGN5CptPQev
QNsqyQ6X3bUuJd3s3VWIAqGOjC9a/dSwKT2i6MQ22P+bTIHFT6bFfI8jtw8F68h0
/nmmsqno1vTT5hrS/Tsti+cvqcHkuuZJejHA9ZanvUQdcSZCrYIRriaiQ5b8Qd7y
fz9TmNkq7cNMLOTagumeIT0DbQmVzNtQKm6/C3Ee+a9ciCg9bfhrw9n53+WN18O2
k7d5pflPmJaaAFlXcFxRRDcaHDcia55UwL0h/Q+XbvmEBVwLqlO2OuRm9pX3yjeL
BO9tHmDI3DitZPxJ1ssnDYYRgMvbRWoSuUMmO8N7eURzak7UhiZnuviSgH6tRp9T
Y/ec+70EBvgcMbSKQHqqVv/rcaGyr3TLOrXuS1UxKLKyhAuP9yYa6cq+ccYlvuC5
T2c79JpCyfRRwuyXFtpvzlmRzn8YT2U3eYW6uQny51Qj7gQo4Og8LsT6s2LNA3s2
GPP3+OnD+d7htlNeXXTDJjvwITi8bRyTuYsZNKXlUdSk8hKzpgcwoAn4W6sFwhYU
Sj1FgGmuhtQVq+zzA4wQWGKbXjQNOOHBebscO8/rQdckXca2pIx8VIUUCYDaGh9g
e226YFPbeK5gZQ7a7k6BaF3LvpqlhfCgU5APLoC17/MqLDpDFpelfjMAg+v2Azm/
4kmj7SzmgDYffcAI2u22u9o1BLQwklZIG06ORyZdjhyf76w2AccBPFpgVHEbfLtc
6+58YCK9DJoVwqFxQ2RHfRWCNWI7IOfGAV8Yxv2gj0w8Dw3l68oJYxnZ6A0Ig09g
yk9be33cQSC08pgLpJTLM7/nO0A95QZQ4cbw3ZEHYgyC03Pvsl+pbJ6PSr36+jZB
eEzK2jeD571q0TZUoLNBakRW4ijvZEBUGbTd/9EsUbqhEYpxK+vAKsQFFtcnD3j1
kq0MPKmE6sgSxp3wZ4ERunpSjtWPm8CS6eEymap3Q9o=
`protect END_PROTECTED
