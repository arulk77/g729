`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCPB65RNUkN+TSGYX5/nbkjFmvS70kX4G6VNAc3JK3TB
l6XB2aKdAJMpHGAmpPbg3iNTT+rBQOQ6QB0AoX9CDaOXEss+/71oOWAktGDNAAH/
k820xiuP6YabqN5UmAa82RWeLNq5kUMcU0pwGw2HBzLX8OV401AQk2BiyuDOcJ69
2XlondPAgW/Ln3nJBv1sebqujrHWN1LioOqfH/bF1Llas/qXpgcL4Ex85+2RxF4O
npyJx74JoXrC9dsCBvXcKg==
`protect END_PROTECTED
