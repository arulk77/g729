`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
EdNWefDLeXTw5H1cWAhu6FUd3uZpEiz08hnvXbyQ2QsBdX9oR3IU8tDCxeCUOzft
Bi8lxVJ5k+50uemAy6qLrj+14BFeqWO9dxzNlhL26lGcO5CIYm4KzuvssdzCkBqF
6jfkFFIocTQlnuNxU6KIDJm0iPSso3DPtITkU9+Els0ILna4u4hoQXs7c4DTtiZ6
`protect END_PROTECTED
