`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCEoEqSGb0sxRudja0EiLxRLu60ehKtB6aY+xcJOEE/j
YE0ih06xee67TqH5h7/yM6mn1SumbjHpndhxszUqvOq46risV7cx0cqAsApblmW+
TAFEbFnxmV5t/drhXvfbhpoglVpGbKWiue4uTgN6tojGnZgxVcjngV/GDPm5hgkg
V7AY3BfMX14BtrBO+TMNQl6qapi2XoX6nYcv+elgH/1jqmipEQPrxVdf+Kbo0rhl
GjiOi9u/lpIYlWDZY+ThuUQhGhaKRltgi7evoy2dp+aZ+gwb5hMdpDs2/VG5q21u
MwDsMCnjphzJND12ZCmAYWXjMLxDplUAFc6mpEs+FZ0GkPUBGYxojhyRpXQqTrSJ
0ivL7lLMT1ho4XOn5jvxlok60m5FkN7vLwV91pnp0KF3F/RBEyXePdpNctGJlRcX
ukPiPKwFY1wzmw+40cDWbd0s78gTXtYwTY9CvqOtdqfPP5UAtoHWOAuhlykwRART
cvlqdUTwNahiC64EYK6fdA==
`protect END_PROTECTED
