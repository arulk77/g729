`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
YJvkTYeBBOorCvXw4oRLUtpqL8/+sSjp9d3PwO6G41U0Qj9MvJPc3Ne3kscjTkiw
K+bJf06RH1iRGqCsSAnOcqDJy9NczckoauMlZNhPdZvmDR0og4cHhBa5iJYQjXgJ
O01HGXPkGy4abdWa2vRHasvWvbxJKiKZC8u42AFRD0Ny/+K10U7f/O198cbVX0As
t9xOH0TunoQsTZEW3YD9VL+8qPr+yL9sO0xMdmClk+UDdaCUx4sQ1nveyeciih3X
fCrnw13M+JAQqEXspGkzwbHYTmdsMJS380n0O8Eava+pT+nw+xR0f+z+aNOvK9Wu
+sKmCga4ZLPDhb5UQ7y2x1WhK8mf1KQ4RZc2xvrfaYw=
`protect END_PROTECTED
