`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEoirQQ6uZvcM5g1L39jjNL0OzCngph7KXTLB/Vw0FH/
e78wNcdQuQkZucLMqmDkg/jP6lCRtuaLf6wrPSPZs+pNG6cDf5SF3fWU6cJopdD/
b2rCaoMhpfHuilaGgnPS5odvYktOMuddX8G6r0YiFCbuJ5cDP1pjV+YEGh4usQwR
T6IAUGuW4Shjqq54QGp5CTUuyaV+ztNr3IwgdbN24E+XHhWGraqh9iN5w7udI36h
NbSDkqExP/4I417SQBrOjqoFUKcW+4loPLp5H/JcSdiDNxTik6NjGxl5HclfDRyn
Ii0i2Hw0LtdB+edMSlXIsIDIUtSCuR1a/z6PlWHhoI4uUNn7zFPjj+wknMPuyaCu
Op09DQp5539nxa1diIE1QeqFgmK+cGMJv+Jgv+y/NUwoTyQZUMOtrmkrwrkZUnW3
RnocMZ7xDIS4kr0vaS7zJQ9zUCtCKj2xIuZ9KXUbWFKqOtDTRcCDRhG8QzMBlD8C
cu5a2ikQruDOEeapWlnrDRKIMZiFOpenSnEMpJ1ihu09+Q7uohNejSjDc1PKUSTk
HpvZ2PArWjZ5wr2HzVco3AiJN9jb3P50CKOm7hPrPVf2pZFQpFfdwBRfCkNcIcah
/yrnSRLS3sNiyJUP4Gx7M/jc7dTUMjHTgHYJP248kY9lFyZjNXjwFfx76hlWKijS
`protect END_PROTECTED
