`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOW83pk4E+vQxyK0QVRh993ZQKX72L1awnUzAEd9Ulzr
WcpNJbjDF3CKrpk1UZhtBQo1A11qSw1Ch+UYUCIjy2/QfMZlFkA7UwIZ/xf0UlSC
rRsGrHhJHRnksgxKP6ParI86H3hgNzSwcjSSoVDDSSfiZVPxQDwZRWq0lQSNMFO9
pAlnHNCkcp/E4nJDQBXkvA==
`protect END_PROTECTED
