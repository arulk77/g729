`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKyO44ZSZvjZLpFIJ0t3EJIOjeM5H7ptZWTotBfgOvnC
ko5t00LatrR1MHOgQXQOd10il/Yip+tHH3DovhyTCG8s8j+iU5C28J6aX53eQ3GO
XYlE4S1h0xEsMNYvBCJaLgLCl7DDZb14rBM7hX3U3nNlEv+39C8+TqBLiVzrxn3N
NufGTFooe9epXe2PYArNWZ3gSwkFG1RvYSXYMUc83W/AiPsmUVvpYNqvwdw4UJMd
uHHRm8WAWjv9xdeiaBEyXbp1CbAPDsQfHzUD34SSsuxcoZhIWcaNw4MhXaY2h2rQ
sbTBtxwkfR7G/indHkQuZhzXqNuibL31pBCoO9wLh/gHmWRbCYsbvXFr39SaXCWW
dbNTKaMRkAKySA4oRJms/2Knemkf2vuj5T+M01wOyp1ctyLNnc8svtzWLzMh7pW+
QAFhllOEvKw6R1c9U4YGQC+QYfHjZavUEJo/fqTF7qIjHjbjJGhJjEx6/mGyTGT8
aiRLvvvIbPkyc/ftG0gid8W6roxO0Ky4dReZwYfVVFkBQOkQ31b/CTw17cXMaTPk
`protect END_PROTECTED
