`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAWyI6fKd3pC90GeUztBiGjQOIJQJqkc6bFwGX4o82enX
8TYOQ9g7C5k4X8QuR1e1DXKx+yot/iEwqNhXnKPxMS/jh+TLORZDbP2eaIJt15J+
nu8abPU7C6XUXKzYnYTW6FCz0Vt1bx3+q/hgQ8BvBdiHqOimuIk0VyyeIf2miNjv
ZKPH+rfxkD8xJUQpd7kCYV7AJv+dGlR1Z5wsNY+AxXaM46P2mWIMk7Rv59evKDFh
XhGgiWQ7leAVnGLwIY0XfOAJO9tXtnDIj3FWX5am+2zUBJoMRr+s3n6rWzKjFRxc
C/AX7vtQIOUkz979Qd9uvjiEy+ijN5nbfaXrYI4xYySSEr5ss7z55ySNJGZSynKE
WS00NbD0DJMxadMrS2IW+heY7QCoL3Yq7f9x7NLnVFubLfUmTAROwVy3IgAbDn6V
knhRxwTK29kSnPxkFo0w9gxeeus1+09T1gh2wNcl23zrCFTlH2f7kmyF8BmVFvsh
p6h+A0Buyj69JfkEpEtpbHbvNBaIwUl+Se37CXfeF5xOzUfJmXYqMC1hWtOkBkvK
drYjUbFWdjmFYNUYQDVltdMfS0kJajow5eGTJHnqsdd7R8Tj3VggiyTA0Kze8R9P
DSvnz3PHKLEfqZCrJxanVF1LUWPyFSyl0TccqQrpFcYJTfQ85oZhzQW2DNiXn0P5
hmUC6Ady+Kt+ulQZzYEdVP5+K8NiBVrxPqrLq/x6p4HRMfB7u41giQ7AxMtpQY7J
ekteHmtLCMEK/UK0PxILYMCde7D1gzAOxMvzGzc8ymRqjWEugddr/OSL1NANn0Hn
9cVveUohu3WjvKDbZH6wWXwUuWZ2lQgMINwBjUqx3IeQ9abUyInbVlVBYMVVsdQQ
GXg0NeujR0RdXr3Ao+AW1GtF/2ZDWTD0MwBC3NEK4lntpB6XUKdK4ReGMNelNZgE
Gzf1rf3pya1yxSdd19dy6Nr9CgasWkTU5Vpcby9jNC/kK/k0vRISGrPN9S4xm8r5
iVnJXBZQAZJ/SINjB4ke+K/r9uuS/Zf6nlzB6bWtPu+O20TgQUrJVunDbnDdaZ+s
h0P2A2cNa4WWutCoZ5+0BcG893JMz2LCrEUhShbxrjeHaVCoflVBWb6fLH7crvYl
42uQEjbWt1y6o2CCgVVTppp2JdEU5VyBu3urXRTZAQlEwfn0MD4BQdYDYke0zZGe
9ttf4nRqtYatgZbIETvf4no3pLDzmSZQzLZSeiJMZWkVH6pIe6c7rTA1UX7k0Phm
`protect END_PROTECTED
