`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAf1h+qDE+KlqWN0atAd6xjZfbn20IYrr3T56x5wGKh8
C9oBsrCaCj/KNBHY5buSd+uYDMT7Vazl1wVLXIBeMFmNFHBrJVzzXKdOJuQLZylD
eS8KpLx5xr3LWLvurJDKTnYNa8pICnPA/ERfAymJ3WPOIhnl8K6EHb45xy+LkrtZ
f6YKNEv2DkAEyYQJ6j0BoUH+fcdpdNDS28YzPNls1gq8Jnvj9E6xfQBWANqP59CQ
tSmbIjp3q6apKvNEW8NaUP61SyLFlP2XzIvXZ/aO08u9MHeKGXkDq/m7nFVSwZfa
dz3HSonWpgNvyv/D0RbCTT8w2KcuiVDnSY6w600qNP1JerHKouX4CMAIgsMJYuD6
rAQQ/jMc5GKRZoN8RjuSw/2bC39nnpiM7I8j9y+xJYB3hQzlBySUDAKXsfu/kIwc
Ouq75TWXrNGPuRc9cX5L5GIX1EQ17aTH8sMbytQCbLGdaQsHbO8MVkir3TKpCVyG
`protect END_PROTECTED
