`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOVOAyiyifpc3u9tTIYGogoVpzJSKW1dWzPFlZ01JsDo
YY/P0QNlQMvYoo/AXEOEpp5qUNAkEWn6cOiCvOtOROrRBdEymPZVgt0pNsrDl3IZ
pS5FNz6F/sJJWkIDYNh3MjlTR5RDdQWEdJAN5XaXeTEitHQHgoscGtzrwzdqZKVU
`protect END_PROTECTED
