`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePIx1oVLXDX646PdgRMiyMQQlU8XjxRAWCBJx4GdLfuR
2T/2OnftaPFpIbUCOa7S17z6UzEH/kocpXnyyMmMnvgb1EJsdK/qTU1yyZdYPZOl
sfGhuV6uDNrw4h7G9l9RjzGgCdQ5xuCKoT4AO307Drybj78Al+T79Z+QfhAo5UGF
WUvo/OMhdkmmLW31C+oE7rFXFV52HfBamkjfQcyXhJ8ZW737XAl6JigGbFMasvaB
n7DrBtrFdQ0kVXzxVYfZ/TqUUsSvoPBKMg7zpq52ZaW4rx/rG3OP+Sw11gcISQJw
5JIsk/HDuZinnvxsAJakRg==
`protect END_PROTECTED
