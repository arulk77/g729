`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
arfyX+yB0wDqAvlehZmq55tWwjC6rz8dr4ycegnyiLeVEOq6JvitS1yU5HP9F4Kj
f7TipuaiqSWV0lhEDXvvc8+4KadGiF4jxpsjyYlcQVM9g9rNLXu60yd8FmpxGTp/
yR3VHxcPE/p7Nq0f/OyhWU4atm4FZXUMzlZ/zigVw4PeNwp4xoN/G8MyXlKGYi+w
`protect END_PROTECTED
