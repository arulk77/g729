`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49MmpTRUUg0xDs/sRwOpksF970C927mzZhA6KStFyGo/
5sGP2lJsxwAf+9OrewQ2d0MM9W2RUtYiv896+pV7LbG8RB6uklcRUCOVSSUo+K+7
fGWixwewV+XBH9ChbrHa0tKb6PEYoivB3YKTvAu4IAekHb+RavlwmMs55T0xJWhO
saqVWgsfYe7yTJoaKKEu91jMaokPjKtLfRFbSLkMg16YIeff0OpaiXJ511f0yjc4
2vbsuGashYDQqd00thGA1jTT2I6K9/Q/ggGX/dGLWjgjYRgblFkRdZaSDeYAD1Xy
w7GuCJYuMlZu6H4SV64mZnU19CJWWnoNiPY5b/laDaR8wQw3QCo9E0ieDi0geThm
KyxBgxNVgyQBbt4OUJMvsTbals4W3sMvYDe+mSbxzOtxnwDRCqUfL9hWl6FgwpPd
8PreKOSmtumLHC19DCwtrQ==
`protect END_PROTECTED
