`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aWKAALRfc1U3O9cKRdlB5AY4RsWWXn85dvuBYaBqu36R
7WH0nflk4uI0cojfDQPaJTR6Bmsfbzy4jC60h+4HVLQSL77YNC/7pDOYFwjDaS9b
/gl/IZNekD7mKOGTT+PWK+yMtT+BnTFw5HVmTAJW5PawC4QAjXqD4NZbKi/5Af7h
RGwBwczPDvgv9bbCqnILZhuOd61jYwjszN3OAvOqJWDxiBRmFWicdK7tIeVPq38I
3TrffwsFZz3X+qDDaibdQDh8q0d7ZpzJXsGUy4u+aasVkRizCMtIWCUs1ydRJjaR
OwMRIc8Jua1lgyw+dGgjo+h3u1QsSnJn7g4MJm34/+cS6sYR/1Eb8mgQJX9/+sml
BveQ15NaUSWF4fHAdzC2Q5quEkA0AluulV6Mfr4cI0tWZS2F2RKy4Mm2Gnc3l4M+
jJfAu96P8ssbUPZyhQvhECCU7EMFk0EArwFRC+nUTklsx9uwR3fag7nKqlNP9phz
38v4En8Zj58NrBOaZOhUHvuWbDLmuxyjEvdVhEGgWzOXGv1p5SAZdcZOlmXwhZYB
/YIRdI1gyGWmD+63dGFKP3iP6l3O2dwed2B8cE7vMI9sihVEbuYovVRaSWMpKSsb
luJDhLrzECe8dxGcbz+8SfWAKQHA/pViv4cLNcioNfMpcyzpQOWjneCApo9jbeMw
t6Qmew/Uaf8dVDlFZA0+eZxrhNGhqRlIc3oWeFmdpkUiOBzXHIq4o/ojGCTYydgi
lI5K58tYhou266xyuwohx790jb8dBzNUsib5ek2/2aJHyJ/2Qw5KJkbfHNTbABBv
GOzqbtmNVmP6Jmx7AyeNo9PaPEOE8rxwql4M0QGeHG4HAOFKt8Y1YupqsMiBC//z
AzLEwOd97BmDmSP0pp3nbcaNp8qqYa5BAKYwHnxJbPY=
`protect END_PROTECTED
