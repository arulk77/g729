`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFO+CwYXhMa9+LnKhIMGnxfYd7lwQGO19tqxo8yGdWBR
zeE0KFB2cVQEPsPtXm9fLosQ4ZV8u9X7wv8DmKaJsSFGaK0y1fC8BHhGdM2SXlz+
ORE1KEmtQxVjOARr+CqtiXqieDftcbIoPhS9XiDqJuZZjfYolj7bRWGOF2NBMuzb
vmzSKrQQdr7Cn0NgjZOe+xzpUZy8yMYxLFyfGmkkCaaAaSN469ovB9BjqykAo8va
`protect END_PROTECTED
