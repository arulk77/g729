`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCXBZP58BIsi/cBvpiDOZJ7t8APDczSnEKGv4EeiQjnu
2ZA/Y0a/iQuO99YXVyjkPh8D0Aq0l3taB4adUFEXG9ogkE51/jTEHqet87FcvNzM
kv5l5d7Y9Lt/hxkrsNDOwKcBXhbGZ9JTPd9C2PqdooirKyfWIpp2BHZMsPpDxuzx
`protect END_PROTECTED
