`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAgMKvi2jPiV+1hvcTvwY1eWxJAErL19OxbtwllpG4QL
34QV7Uq+f2cCCOP4F1SuZxm8evucH6Zg1swhIieD5WZEWLAUkZrzAFLhg/feQqKh
NpPO6tG+TUfNAVY8cK0wzMp/Q3bGgSC83uKGq0d44+QZgHwCOIaFFTtr4pe8sDt/
ru4aPYednFypi+QPAa+Q8R8a1FuC4UthlUfxyDURw9EEVcqXCsVgZyNwlw3oxj27
gxiSeDcDF6APFskm1TJxIGeLzCnZt4eIJxup1TBSqXZOgSVOdtx7EFO78ay9VMUQ
nXMrld9Tz71KLg9iZ8hQcsNCvlOVcbeE73/It6cm7x6ySlRgypMe3IpHb7Jvd6u1
X9ZpEi7S/42TBeoIpDk2tw==
`protect END_PROTECTED
