`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN7aDyTnZHhoAbUTrntCDzMkynzaTzejlH0/c7plxm6ls
VmjIgCmS3Go/N1opJdIJnESPU4iryLSG6bQ2e9ENukVeFiy6kJGpK15++mtpDWpt
mnnB2X7qGpYPUrwwmk2Ry2Z1fq6bGZ6rcM4KynHLkcn6/fMy2DKTHklY5n9t/T2G
VFN2rXUYvbaGrgMN1tuoVowxKyfQx1Ll17X1XZWjgd4iC5DvgcE8WOcBp+49j5Aa
O4IOasICEY7eBWwre/kJVdU6t9tGj5+xxh6GqunzFx244tWRMoblFK5rcZVN6wvH
i3lRu5QQxU6X8dXihV/+cZcCLyoLfonjcWGt09XO0FmVem9rIDlpQAfDma82V5p2
v/xWcnARov1wiwG64EL1myfRRgZzhXwYlbGWWtn46HU=
`protect END_PROTECTED
