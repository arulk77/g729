`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
A2927ATXC6eBL+C2SHz9p+cxBuer4WHQlJCqPZNO9PYXPII3E79R3JwJVnmqOvHa
UQ1zQf/KUEE8XBvk/fqg0Xqo7Kl6I3JGpHYxq1koI6evo/2boAo9p2ZEOSaOZWJH
gxgFGX9b10wZ6DRxgoBWGLf3v5d2yEI4+ZsxY98pPVL9oW4Gx/RfrTHoa84pSHV2
kCOz07XtvYcXixkibs0E7F90Ty1m+exWKOpknZRz//5ibJUsvNHdIxyKgX2FnVgY
ztMLQMig9D+h+zRiFB/67ilqyozFQDuQ85LzcBEPe9QBYRBxHaZB2Is9R3tdPtdX
3vSh3Wxcs5X9qmJNU4EgwjwfJyNbnujh2rRM8X0DvxvbUP1wdFTdIstq0HgSqi2i
7/BsmFhkLz0ItrZnp1sguEwpHJHTuwioI8+/XCv0Acqygw8OZDGsvHzNwf2pDva1
ptmdjLilP9vL5uMritObRZVN0Mmg1Jpg8wyNCF8dyjl8Ilve404Ckxhx6/G/khz0
XUhTQFMIjeoJDBZkpwI7Nff9+8yeWxDtlFtGncWaaZvuPJF3/tJ1V5/5FK52OCn5
JkZ5vKKgJJ9QkSUxc7OiuMS4fzVdN2uA4ADt/h6epLSWS8O/z4kw7fBZXuTym7br
M/pmqWeMbkoEkw1DTbUKhjJiK3RpDD9X99FQ2R9if0mtXDz+sefRFT6b9+VolStJ
ji88SIHDcEGZKSHmd0b3yQTWZ1sAfVvA7SkoEHAZjA2cqSvVj8vuJuNHqW6oMrRj
YDA2Ol5IrpV1kXM0qyksPoPtmhLFEQrlpRCzszGXcaUlIaX3R2vXzGPBtvx+8psz
`protect END_PROTECTED
