`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xogxZiyDyKJ17bKN3B1Gzoy2gS4pwckJe9V+3urxB8n
reL8BIIcydBAG+VaAi5dz9m3N9yHWGHS6YDqheDCoXvebXcLDlu4doUWfxv4YpfQ
bhm/V9jz4AWV9Y41kXA/v3I1rPN3K4fkJ0m9fNam6xNlyvoSXVMWptEyTDFN8JJH
e9w8fHQ4Kr5Ib5pNPgc76+Ck5aE7YBKvQA5XrYCUtbBXcVr4ISK/EYjyWLXPU1+S
8KVptp5IUjzUXbppUGF22wJtODkF3zuBYtFUHg9O9g6pBQcitkp0yBhrOrp2q1DR
L2ZPSO9KY7gCu4FGzEIR0wIWzDSrOsYaR8Qp7JBLbYWgcIR5vu+cPnkMwFpbtpas
tSerEDNOgEZiWZxEUiJHs0nXK+UNLTfbvrPab53tgC5KJYoNOhF3YiBlHNhg2ndQ
ydshvQGyfiDffNLS2JnZ4g==
`protect END_PROTECTED
