`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SRGjiillTjZQydpO/XMzPELwhmXwR7dd3fd0sBxjWVmH
28biyrKBZcRA+8DXF0tTeEZbA4E5Tg+VdQEedvBmKIH5Ydy0/AwycKW+UgLP4uUv
YWOTiJx4WeB11nczDGS+CzIO+12qKeKOR30yyZ2xb5lnV8Ey/GoggRS85qgB+D1O
kmsQOR+xp4lvXzjtny+RrpU1al1d48gFQ/WYKGoVeLl2nqFfVg2ocmYxftu4+67s
KHvkRFA5vW/SElBCplyHjqhmKq0uEwMv3qEfO/yTUE1kmq8VoDTDGa0BDXE5wVJ7
HluCWsnBFRwJTnJAVcFo5yivZ3HXk2iGVXl+hWgWIuwSOQcH1siSf7mjoYTVB0FK
V6iFFeaR1AvqhX2H2F6klPbvWRNbYJa3GMbE+zyDuLXf5sd/rTbescmMFsfdmpN8
MRFVYqc5LXrft03GWB4ObEUWAX8Fof+INRusCh/kbUez8Y42F+OpxepbCJmTwagc
8v7jlTEt+LceGv89LYhvIjKGCwr6WeIppoFV/HCx/2QBfV9IpSd2b6Fp1554YodS
5KqIrHh4i/is6IuyFAOQL/3zXjPHPHMHQeLtLAWVyqwEkiY+4ZEqdNLNWRzq2T7C
wCKGFos8YpWPjVMdWTBeK/+HPNsHjV3UHz1v408lVWDLVaU+NsgObfrefr9lMPR1
mIhf8rFRkXtN/L71l1Eb+5o6qK5ljveTDMqszNPZ6qKUOAtnKHuNPrzo9zWu2jn9
+x2mTDx1m8wpki6zvoG/9oLfmFLOZBVOijUxMXRXtHCNmm+LSip64bb4xkoomNbf
6C0BSIcnc4SseIz7IWF31GGjoWv3F13vFOTTfde/IF/KOt7xcpRRovJiLe+BB7VA
Z9sZ5291J1ID0tiBtKuIoWqH7OUgJrxr71glljWX0d3THp4TTadJ2PhrDvrbxx1w
U5tRkFIGGCdB8kKerPkTa/zxxzBgrw8EuYYBJTpXUt2ganGcS7drp6UmBPVrHLCz
FkRY1MIvxiLbAHOl4cV/ZWtaYSrIyZDUGor51qvz/NrtQY2J7Ljqo/vSnlc8PEQa
ltKyLvkFuXMbhVfshdBBSKRV48MyaPnQgDnL+BfNXoMhNR5Jt8ejrn0oNm3t8PBE
DxHsD7ZSkR9NlnrAd+cIdIHboVh5Az7i+nOnVmOsmpz1oq9/ZwQhuNc+DgXzAoVZ
TnDxigwVoEc2wLpwpArth+jRsmccnOp7mBk3Lx+qe7HeWsQZrI+ZGCRr1jcYry0l
RPNIM3LnwTvVjnTZ0GeNBdrwp6t2V9WsjywLfsfMPGFfMxoFj6nEungU2TGDbm7g
fZiZwxE+zxzciIsoDzQSlHbkVFJAsnoBYeKczvdOLcoYFbWRpSnt/a9qE4K/upnY
CPwNahwiF6DezwiK8pzzm4j19JHZ8uwzPCg/ale78X8VbFzBHIFA15KoJINoV0mA
g3ch/vfvU6b5jEcmI2h29RYGtkQfwDrysSJo+jRGS4rC5zGbB59WS8TmIJYVYGbg
AL6HJH+QpCl/YQHUxfg6ksmXF39xJ493IWXI3gb8E9z4pD//oriRx0a57VTsccn2
D3c32R43M6DBj+8sFbHY5W321ObtIh8yHOUOcGPFkiQ=
`protect END_PROTECTED
