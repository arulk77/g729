`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePzk+R+HB1O0e+qnOoZ+DD+lYRSuG3/oFhszFPB8a5MT
b7OGbMnRQMJXg6MHrvSyzCkCaHuOPC1ADmSBUWg3HBIjezLbuibSmsh9zbDK3QvU
iw9muNWicvWf0zbL9tGvzIClo3sxo3pWI/hn8s905KYvEEH8udBhqQ8117TnMUKd
IvvWqotJJAqTWlIByn+CPQ==
`protect END_PROTECTED
