`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
5Aas82WX+NZU50I3ANwz/rs7VBAd/MxTkFW3QqBMMp2SBCcl8HeedyogHNFYxgQm
MmF1TCNxs9dYGa+cIcIKuG06FOvE13EfynndN7xxiYNvo9Jxou3XtMpZEBeH+KNo
8J86KYqxwMpY8kyF2pQ+Atf31myV+uRMDOXR6pLpY83Y7BzCZ4QC2cz1cXUOvDCO
L/sjW78AxaDmuPY42Yi54ud8dutuTokioSP94iFthjl2puW008nOkdY8HybWThaF
AMjGkky9oRqQS52I6OSRMDTz7AOAQUuSxnUfESNc2QiPUyaoD4aiCB9mAUibapkh
Fh6o0nUUwYveYiQNDjdPIBHr+4ayK5irxLv1Jj6c9YU=
`protect END_PROTECTED
