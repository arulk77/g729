`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu438qMASl28RCPSCzXGYfNRZUoaOykPZNiTSYpkcvx5I0
XDGb4wJyceGtSMYJ3n2ZE996MZSt3ulZmxGiIZ2rKC/34h1CokiGk5HU0z/SiCk4
rmg+k9HptXi5BkbQHzVASgR5z/Cl5i1NjeyF10mRe2o7dqrcjTEDz6x74EL3hXqA
UQ96wR0twDCWKKKovlj0JFclb4zQ2kdPxiDfXRKX+6LNXuVah3bysUIr/uV/JYPq
YmLI4LBhErl4xVCSZOD7YhyzyAMpoPgTWTlQjesm2clRwAmKWyzQKuZ6is0IcvVZ
f+iY7wEVlcJpqgNSpWugoQ==
`protect END_PROTECTED
