`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73Cw1vzWhPTAGEneUmalUggn6VHrOoB9I1XGKgjChyFO8/
TX0MxEQjYBuaAytw+xRdeKPZ1/ardICa/NQbh8siUrPR38cG+8T7W9BPZlGO5wIu
aFs+lv5b73PR6Equ1insbJprjygyHGYneFIviWgokNH6OmfFw1ynhyW4/kzm5Jsa
ngi4BlXiQRY5MGpeq/qraPfduklhafeYIg87Q6yHb4VL5o+dUoneAbTE7tPnjB/f
k55Tdu3NvW1xn3URcOnY0S8utWCBeWJPwRWn4cRrUqmjutqajsF/p5St6DgwxwjW
5ggbp3p0jWYgeX5fsHSdHuQ2bP6TB4jynYfuU5s6G/eNTpCYenBTc+avyj9SNxId
57nsFzEeU5hIwdMCoVhcJHgGwlpP6DjB7QtF/W3aguKQUasKcMKsjcFS68X9Ujtb
vuvCA7ZOxGoNCtlYv69OpuEAPpBo4CPQoWTS1eFL4TY3vcpK1JaXu6VFUiaYfdgj
LC+mjb7QWXA3aNT8VvaA1ml0iCGPkz136rsmqZrsowvVFp7ygx/Y19Ko0p+ImEbu
UzSOxBeyQZLpOtZRrvW1DAxTp9u4G9DcDCyMP8Z8IT/Sv6ULv6NkD+UnJ6sszFS9
rKa+l6BGQImKvnmB1TbXNiWVgT1JYm/GK6mDuNdfPS9MOCaOnqckGm3ZOCUGYCFg
`protect END_PROTECTED
