`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI6ZdiP55JhDWRzezf/jU6GBShuUMu5aiV6g/6+huN1p
og6lkd80Wgd0EXOmE0ZCZEmg4VGryCu3+HYsMJxToYs9tuqSFZXrjG00sWO5diK0
8QMX0xCjkNbw/2ae52XYBtVDH7lT0nWs2BipZBhi9yC4//MZ65qvWgeeYu8/NTMz
`protect END_PROTECTED
