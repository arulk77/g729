`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SR+RIE0vAxt36XiC+/ZBJaLUCQM3ILmwI7i+Q/vtSsEK
hMMLUZA3QajOtwcPSByblD5//338vWOpQkJUKiFFlHgCElY7+6QyC/Lyu0hmPPf3
DKaJYpKqwOCgwtvDgUPNfikQ0Si/z0tW0fz+0/rarFccEQS+puAK9ypU1Z8SPBRH
M2MJIuwa6BOXRP2G1oIgZNWciDz6LmJ9P7HSbrQHh99HONet5KR21ixD7hmH7+zN
eUUmfjrE1QrIJRNLuGbZHIfwN1qn4MJw6qmp38OIP/jha2hOSJqnEiMAKkqNgwCh
`protect END_PROTECTED
