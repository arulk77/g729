`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
36A/U5tO69wVl401zVMLLWGRHPY884BFZQErSsOZVLMSwcai82KBcTELNBTSBEZv
MfYWG/KmbUXpjwU0up2VIIG3yU5yT+ljePT2oWJSDSRXiM0rEfFbKd9VUUDtmXNM
jNkX7KyOLV+AYpCogxFp42MOImOW+et1Lp27gm5P76/KvxZLi10fezVZFN5SSGyr
a8Xwk0W56vvSTgy/I7Imcq9Ql2cGESyMkRFA59RjTdhZv/9qMRrKWV6IFsGjGeor
2Y2WojUu5av3B/pOynp4FTdXTMCB6RALr/x3QPaIrwGr/DX0yJc5yRNPWHq3cLYY
TC1+sUMm+Sza65QCWEDJ0+D5yqt54xsWfsOt7YK1bj9toGq6bKgIpWO9Oq7xUdxF
`protect END_PROTECTED
