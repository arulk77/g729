`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDGSdFx2pWWvzgygk8BrEtLuVkB6iV5z1fU3fsRkQ5Vx
xS+A37hwz+WOhXT5bKafs3owXgJKltAm38+eHxJL5ie5W6YyI09AtdHxi+jmWKMb
DjhBX3GuqQstTBeej8MYLH0kgJChsWZbAbHZ2M/KGWqcmOhRXfb9rVO7iFQZxJE9
/2m0zzFjGa2ilogCMFU/DR2MRWhMmUOiMgYIfeGCNrpT64Qtx5flTq/YI+YnV08X
D3OImiH2szWuNWFw69VTkc8AXYWrWr16cWKJofbnS78EJGHfQderz0Qq++tk/xoT
l4XPSVFfpzvnGR+HZYlxppQaxOOyj0UxAuuktN5R9ryDYMCiPP0M+2U73g8UebM5
yia6mMsYtNZktqUSnnYYsiiT5sk+ccqtYKJiFRm1LjBsJYxJyBRDgSyy1ib+8SrF
TeUsjQG8/ORlLAPtMigf2B4/4F/7McktHTUXxLI6V0NRMM3Iij9ZWdvNK5Mu6+li
aAgCNPw6+XNS5n0m0SB0I/QndtXki5P7c1E1unhT1rdTkX3+Nx9NPN6bhdENHCY6
NNyLcz6cnVfAa925/pYV6wQoAh5U+2hjZvUt2HK3+/k=
`protect END_PROTECTED
