`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEKgHD5tfQ6XGWRxT0ccsJ5XbTm/qkhDQbC1UcPszFaD
zVfUmIt/lwdRLtgY95n9OMpRh6uA2VggO9bEdxsskOCo4PjC6fo+Ac/i4Tiz/k+1
rt7g+GDgTXVCcs+3e64am77I2Psu+U2YbwTi5V8YBcdKSHfSV5PGCZzCydBShUu0
qtHEM1wJeYlrt+lxF764PDA+9Tt0dw9BzvJO0Ygsi7DxH6yhuFu4bWRbaZlgq3Mx
BoCfch2li6C3AUUeUR7oSaF0WgKlivvOS/7Z8r4RCE2bmBUf8U2vRtMEDaTUFT3D
XYq7gifFN6BHEx4LctrKWcknyYTl86uczYpQ7XE+4z8fs9VI6qYOZNjtCXGUql/V
kIYiDQElcXHSQt/jzhp3WYyIJs27Y7h1sXA+ZGbGLrvCzuGpQ5W7rsPnHJAKc95f
Bd+6nQtAxcd7PZWMUJ7KtvIsoNaoQVTku2aSIw6MsRN8cGcxVF7iJuzCAqw36Eo4
gQFveTGidl06nZr8kRCXFZz8MXpNinVNvsGOA2ckeabIWMiPtZ2XyjARv4f9cGn8
`protect END_PROTECTED
