`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFUTozwTYa2Kcx9uo1xhmn0hrbn242J9qaRU42j6uYg2
DlJIM/8FELD1JcbrH2QrAU1Zt2P0VCsFKx98KzjFVatOjl6GUGq0gS1nAKcZrDr5
j/+xln+vXJZ9cAkyEF8Qwr2pb5DCCVMjltj/YPQb2zS/DRShHBHFiUFZXplYHlsx
cGdtfoCpthQU7BOQL51x0QZhOZcEWVwjtA5rTP5wtW1g4nFAmnTqGiIMM5gygbjD
`protect END_PROTECTED
