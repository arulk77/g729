`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xDDyRBgljOmyzMBSpAVodmFJVf28ldM19RCF6Re+Mqu
RQWiD98+9D6QfvR1XMFKiVZGe8g0TEP4Ol1SFGFjFKFI2ESzeBSlP3ajy60KCChc
FlRVPmTzcXiiW2z3eXWJO3HpLc8brK4FW2/w6fQsTS50aUNzSWYH10CQ2soz3/pc
2uFj5SQeGxaugWtP5sC/QFuEd1FZYKcGWFM2uZ6vKmPzQg/SnwztfUwWiIBlj5d/
it2raDYfALgpXdjWw5no/q6hHz/XO5/HFbCOymUqKpU=
`protect END_PROTECTED
