`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
84AZayied4u/d2eNPxMP9hRgIAsZiBaFFxpwTHvScqlbFkge41ShH0aQ6rSX2HAG
Bz7HFjZaP0BC4Z+anhKoySSL1+IxRZSldpdpKTK9YGkrF6yo+zjgJP5iH9z7DV13
62D+/QiyiTWYd7tk/zAS8FURL3v9aDHxBX2a0+cIXfKq9Ios+CxiLLIyYKUF0I6+
PoVrwZ1eziTuTxkNQlNycNgAquvQ8vSLlQlGCb51ezWcl1xdkMEbYy2Nxv32qAI+
fn09JhsqGoOSu9RYSAA7XyZ01TkVHdUAiuFFXrL2eoRDmgJmJR1tBv7blgD+1oOl
Gmw/rxnORF6sJoXxOVit0G+5X5u/HOFmz2nYffEQ4Dc=
`protect END_PROTECTED
