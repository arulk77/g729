`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/L8KYQWnMBQQ8SFV+o0O7LjnMMQV2STXlp3cqZ+bPZG
pkREz1PhW/YsvxhZpO676KtSfy13V/1+y1CyxjoVTqGSm6Ev4RBrxr+zF9A12duY
ENMHyTj65ReYeyWvzOveVlDtRNBBwt4bYh7bvyN3O1HsJfVvanht1bubs9HXifvT
SS0YwqLbZ8RviI/2JvSToDU87Cnvdlp1ZFUbt7M9IS5CyR7+b8MXHm/EP9eWV+Wm
FlGZV1GDJ2Zu7MClEf31DBokZAGrLuPrQDC3Sp9KYtjGkJz9JY6jchzcELszMGDy
VnvFTH2/S3c1NI2iIS1HYQLEXRpxuQNhbFHHPa/h5wPnslDGgCIaG5yRXsaOr9Uq
s6ehBvgjRYi6MieSy7YEVRQPkYnkvCodxB+UnzCxmdLZVqEVX4oy7GnU3lIOj4B/
U3ieoVCiIobuxbaDIgTm7z+gFqN5bXClXcE3SMDCHxFI8jXWYvwfStro4jDVjFHb
3DqZB4KdJuw+gEkAEHjyKQXxiL/flx1EFKgwV1v9GbjsHHTYFBKnYsrpyWKB1NIy
ydY8XPV7Q6RMT/v1mE3ngfFvnnPQ+nebJE7Hi7VJcDx5hlnfAUBQvYsobiz+KG6w
uPPsVG3JPZkfS89c9ZbqhR3GspCnTngYvwj6yybZz9inKTvcy3h0iFijPyFJkY4W
`protect END_PROTECTED
