`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMVUZ3+XpF82WRMHb2wbPBjP5OimTnKLi/2aqP1UTega
mqHLph8pdIyALBq29hRza6p8WUxTRr85kN238fT1GciUhFZ9lCSn0ikhWJfTL5lX
S+Oa15T+xkz3myMPt0lyMLu1QTs/e6XGkxcaxcG7g4B3j9FwKQKUq7+8s4nH23HC
HzXBlrSxV8xpl14F19Gw/TD7/o0TddlvhB56UVR5DEyj1buuRL8huihEuq0aKawk
5R6kuwicjGe6iJswJkaM4xUFlODAkvk2ShCEUwEYLUPrVy2AKQciApevN9bjyVcF
ZJwp+JfNl1p3o5sTJ8aEdPYV4mFyQAH2fPlQY4vvQZt0+rxPKSKs1j5EhU2kpM3a
ONU+OOJxNo15NKdETM7F+Q==
`protect END_PROTECTED
