`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEqglhKKK2QBxMQB1X+aH/oXW892PdAjqiHmVn9quUGc
cgQKkNext870uxY3R6hxLgGbRi407dGCxiTR+Qz8lh9LvgeJixzk+byiF1LpvB3d
tqewIQ/lz+ApRUWoj5IFuPJ7yd1pX3APHIz39pmVqUEJEh4pwMBLe/LmQdd/oG79
zvuGjqbugjQuvxjJDYDrXw==
`protect END_PROTECTED
