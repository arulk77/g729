`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOSuTXthE4w/DGFfZombWQWepk2YbOkNljZVsFV5Iw5j
WxdXze+EAk9/yrDeYLyuc5Q1tDMGBRYomlmDtDGmU0anzHs0ddkgZHy65Vpb1rSv
S9ek+NsZzgOQssqpgAxU1+phXW2AQMpOvwNkFcVda9pCNCbVh6i8agnrrU6vJYj7
sbu3PsKUIetFHZYTVgR6DA==
`protect END_PROTECTED
