`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDASoq/j3VcMQucrH2H8bgMtCms7NeWnGwL0LpJLA4xdfa
hcmdy3PHIyb6fYAX70bAP6vaIhpta9Q9ja9GVOaIxEu5ReJCe6DFDMh3hDcn+pw+
ZhfM2lUJg5A1kAkdgkz32mynLSD2BvIcauefwn0irJeFL0CpCcrwGIBEBHAPJ/zB
L5IuXIyFkaSVxQTggRSuhTIgMqUd5BgZoompNbUiE2WNCmzwDsFzVZh85Qp2s+k+
G5SRlC2nUojPkFHsJfPkjWbGaEvRFmxbBxv0uh4KmnUjBPFB1Bv36PNcuozBbJ38
xSwrkORgr4+fglnkIfU7SSf9yMkaHD4mxfr+LS4EyhCADnCSjLx/p4wZIcNsHfHp
yJLCJwqN2otkqLLm6R9NW4RGt7YWI9B0WucRBCQlmyqMpdKsKFAUb+eD6HGANL5i
SD+DzYncTavBVSo8qv3bOamDg8c3k1U+WY0gPVVc7jDK9xVPDmfeSTzUwffJOUDG
t2UZpntXcsPG0FuDPxI7vv4rQuiT3+b2YaL3a+FAHbfOHo6h1IPw/iTgslr3/csl
cyC2+0H6vcktSvMKaYTIVPE/qog5snZ5tsWHxjyfjrF4ShnhJ7TMeYPmpxL/pbq5
QzkE8VnWG/8NyjLvs4WUkD0Ur91vzMWp8RlErRt+Q0MmPyPdb1ZUdmZH4KkiGbx1
yjJUOmVKGlhPJHjlAZgnBblw4Hfe+SSDXicX/Ro/A53qODkc+W9XbJlyol7spO7J
bV0QfGcGEIdCHxd2ezoMVl1sNbnJ3JWKY2WPLpMrH1SHnb7RBqKqokdai4uapew7
3spF6TPkQ8IUk+kGCo3sA0Nzj1AHUhabwxj/2VOHpQ+YP4+du6ImackTuEgY4tYn
ZmbBvQaXEuQEAXER20mIbt7S+AkFhhcvUDZinYTojNzzVGcq3Kr2c+Z7UxUHg5JG
iBQHkwhUALOUuH0mAj01RHrFeFb01siw5+TVDFK04hPMb2X97Ib7pg9r6eNjsmYT
bce9YiaSH0GTAHq9notj9bpe+VEKSd/IROrk4mOmKbe2o3HYbvWY+IAMOOQWzY4C
S5HntZ2j9Q+HL8Z+EyMue4oel/Xk6LixIhaSWpPw5sA7rZiLTqyfYGzi476nBWhS
yaDq7QVmRYxwhMXXVezUlSjjnmnstzGFn8t7g4PfbFImYEaOtl/2/mBSPSHBeCwx
IfDWBoW4QR4Sw37e+ffU2vTmyjOee4yK4rnCr7ukmffeSg4KobxGDJn9hj6IW/L8
nYaTgytnj0LMWu5YQwx51MHROgEpuJXQbsvSo+MZ7KwVccjtrht+xrpDc3PU9khL
knF3tuuRtBvxAGKlArbczl9WWGRpY+c9ksfceM7DHNPon4ippccOjgUHU1faVLCl
sBkNuK2DO/Qcnlpc7/0+dn6gsR8wRlYVnTMD9IBfg4dlfDDR0hlAVekvCieWjRhH
qmN26PrK/k+8RjBK3v+MUMtgWWPD1mreuU0plf7HTsneJhsj4b0IezFqQDKPary/
iuDpeSP0AKIwkH+HE34KEaAdIaIRMhuhV5Si4GfPPZTIzBg9GVp0yOFv2adjjbo3
QmiHkIp91oI3Q9WueINSBHh5jv3ghMFCUH2TRhbY5Y0KTZ04EQOIbOWyWmhvCjB5
rNx/CwvvtmjLmKzVaRdUx3v2DvZWsd8BJvh+ytDBNFZqVRAQ1sUOCm7cduHuIv/j
k2tUG4lVx8QSrmQL8T+4pK7kM6m91h+opo18D/2Y/j0FTIHcPP2lPpdQvNM9Q0RM
i0NYSLu1/mrhwUk8kSskuUDBX3QbmZXmcHL6Yo3xGac2QXXuD9MeNUuy78/83lcX
9gUJepu0HZtlyH5XYKaru/Lmu7ibgm4L2CCToqBwvDFH5t8o5KLYaeGzHwLX2Izt
`protect END_PROTECTED
