`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAAJO/ynHU9SQ2mwT2akIl8LKSkm0ZCGRMmZII/jMROP
r4CZvHww2YgVkEZ1O21OSmAs+1L3BRlXmnnhxHiwd48PIKcxV48sDOvaO73DUpah
4NhD/4rtV1X0/yBeNKXxX7wQEfKKQSxWu67wRckp7EshEJ41BFQ+TClPUOqg3Slu
`protect END_PROTECTED
