`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFgMheL2dXK3Y62yMQOJlXS7EgTSUx98TThdA/rG0cfa
U7cr8qmKtwFrwFoV+ozhc6IEJKAL9xANXOcdqBzZ1tY4RXkpN1fObATFIbpx2Ydb
z8deYOiasv72eENSQ//0FnXg989BDuIUeQJaguI5q8WCWU7/iEecgC8Tslh/Dmav
tGPHWC/nOpY22ei5BZJJETvpyjRJCFE0eLua18pi/uB70Cac7vLN2dPqfKLVuTJe
TaS3+NAPI8LrRqZXcoimcxMGCKyxh+SWrblug7TyQC+4WB8ux16CTMbKcKQJKRbg
oS342X9nJwGg5Dt9aMc1SLc2aA3/SLJso2eKdyBKy3znYi8Itw6rs6zfQOJbiPca
WCFnQVd5V7Vl4dpSuQab75C8DeAWiH1zS1cHo+DwkDEJ+5sfUYlDsDJ6ScEKWz6Q
r8/5vd3ng96QcL1V15z4Eygirh5sx059Y9fTvRhH2oI6DkVIdp08zeJfEWsG1Tx9
1D9lg6TRFBHc5xhTcPaY0AM8M2I2zfGy1sXRPj+SICVTQMGc5lti5ZmE2w5nwv4i
3i8Hl3Ry1t1+RdIjO8VyfflrowtPrLyWZ5t2QWZiL2oVHALeOAZDh3mw5tI2WW0M
X4yfsHSMzPOeNYS6KdLuoU0rvfxJTrWP/1PQcqaHT7AcIdUhYwMneZpqMS5sh7KY
mnktW7K9bpkKf2nhnYfbrT0CR3v0uRVHO085mPq3AX8TP2vP4oMIm6DzrSdcV3WV
6wUbQJ6gn7uRldEoPXhir5EybIy/nW8ZyyknGHF0FHFOhKm6/drL4g1pp05iwzmK
a2y5FhnS1uvxNI262ilGdPNMWl3sVCWMp0hDRO3lPnM=
`protect END_PROTECTED
