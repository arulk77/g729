`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLaWrOV/KyWpso8SjKZloufwNq3ZnIf08UFjxFtLh+5J
j6KCDlhUMsROiEzSC1tCeEM3qO5VyU+VY8yk0i96GXVVbHSMzpgKoUsq/mOJILJI
/lX1Gj78G20GPpV6bK66cJlQRAayFHKeeyUccHS9YRccVdSgpaWgZtXzik4v2uHy
d87upEDOOLi7m3BuNOYWzQnYBCDcskMZol8nKPxuYxsAj3Te4R7Tn5EI9sYpOtbc
mQfRR748MKtM8x08POZI1q5NglUKJ3/0VX5X75GMjxUo48lQDW5w1wqcrZBsZs4C
bQWm2iU572fOuf7wbKfI2Cw04QhXv0Ou2Of31lnPVCRNYtSFHzANiOeKQ22HZLKj
9UF6RC0mjDjJQYIjyInVyCjWcd0IeEc0t7p9q9k+VNwD1fbQvfU+M84EYne+N7j5
VzCuhdAPwi/fAEru3+7D9fm6SNKoxTGtyuf2NK2nzpBno69lW95+Ae6DiphAuIz/
4Nj9bo3ggNXWjWtfRDogXGhdVWuwg9qSqw+HhoOAIhRS9JqexTMit6ZyXiF4HYVl
`protect END_PROTECTED
