`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIlvimlFD2la225q9erFTUN2BPhbY8kxcYD0xQX/Jr3Q
oKeKc2XVJ2JiK6IhiNG8zSb+ODXNB7B3kGq4d8vKHO8qZ1/7Dstvl757ta0lawGE
Vq7m1swfqHoCxrm9rTDUE/2yzBDVLmyyEo6i0NjTUKukaQ7faEseConI+O+OM+6l
BeYH7YU8oUPhCYI/aE2kZwi/DRytkpdnCMuLdFJNdlN9ZJkB41PtFEJhUa98OFHC
2OaT5kUPF3M9GkmWMyevBMDEqgbGPYJiHRTvoKzyH3tZS16amMJs/aRTQMxz5pOi
6S7EcD7mtx+OU7GLYyJjm83lPdzGk/UuhgJIrHllGKvYAK1NdnZe7yrC3TXjUMLD
6Uxvds/y631YAhW9PlnMceL6qYvMM+wBXBeb0Xy2wgfmlqUIwYiArfrLxb0/BRI3
QkQR4ePf1yi1rfBX2V6nK8FmrypPY/cfK7A4P0LRI6j0ueRcEOxSLZq35FAJqunD
zzsAN5/2+JtN/AxcC19Rt6570hIMXRjgLQm58VMB5P1bVDMXyxHEIVuLkAmXroLY
`protect END_PROTECTED
