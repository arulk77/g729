`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pnyY3jxGyCgnwWklYcFi/bXMFnJwA+inHWmKmO8gIGK2NIqF8BubakBLiNT6hvsk
wpolh+hq30r6tL73WJxJL2ooPD5jKNXe1XyrSP/KLhnfBJjUP6WPCqs+yAt/wdF4
y7GvmplbI4GJlBi+sLOIqDIBgO65S3L2BHVq471BuBKTT3/01wbs+ssDt1IhWwHY
C70tT2ZCrK7DTNzv0jU1G4Y44opchJb820tYIfi1k1x451yvkmlTjQ7mJrJi01R0
9PfyeBYjtikM+HaazYL2jTw8C+Tmagmo57xXMajwpoRrIfA0HpN5L8EkdFI0plqC
MbMl+4k+Tawnkg01Sb8xV4Xv0FVZo6sHnljsO8fDQ5gqRBuvZd0vt/44/GWj83S0
n08WJn82StEgkZZc4fIq2udfiz3GvB+yhSikVGpC0fo=
`protect END_PROTECTED
