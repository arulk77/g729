`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42utCncO1ceRBledwx2zfixlLdzcsnv607gApzae3dAp
erQRKfU+Q7oQrfavL+l2AtxzoJVrTZfpzNglJuXrVP+4sCUIDIJLUPD0dmRGr6yi
NGDIapDUiueLjaLxKS84Ud2UoNsHvTkqgMcbBIMz9J+UWs7iL/yT0EVWHGGBUH+o
yifvdYH1edLF9qHe2cyHhNqjz1d6JrE+2G4nX1DagyT6sanBQju3eI/sGRCZRUOQ
h6caHGKTX0FPu3WM75IYyxAybApfXpSLEANBs/qsNtvP75ThwfKn4b/MzgW2J5WL
0/bv6YVYqAAZzgwACdTZw32vm/Vy+uSMaBQ4sFQMQ9eIGPXRVRXAlSLuiMSfGtdy
hLrpiVPRWYLk3fY4u1q8aGfTMVOLdNxxUT+zR2Ac0MKyzxf81q5qmsDs9rFPR02X
jU1dKxJyDrV8HT9P/5c/cA==
`protect END_PROTECTED
