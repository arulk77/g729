`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
lnpf4ModKYOuaIeqPeKH6cJANUkbUQeZ8ig8f8/TIv6oIZ9c4ojJDCph/nwiF2bf
6pCkpKC4sK2tEE+B84/tu/Avv8AkvN22rMpNImYwSju7NxJNNstlTGssdfw4qoWt
A9AjjEjC7TsNgqN1cBrMi0L/K9dtqu2/Ux7OT5SUqXKaF6y+WYe6H8kxqS0fEgvX
`protect END_PROTECTED
