`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkahNUdF+NPEQ+GRJjq43XneE4S2e+S5iJFvXYvJ1iEkx
pbu5yaLhoKtRIUsYwQL7lLSCksoFKlWL5oTK8Dps3S7tBCxp5eneb55g5rvQmVn2
cRieYoI1ir+I/TCTl4l3VLPusWdMCx98J3cATFbygBiq/8XT7Z5l2Q/1IVPDh7o6
zuMAhB5nMt669KZ7yc/CZuZV0tdjZPEAB9erJCube6EZuxECYbV20SL4HvSWM2Zr
dH5bzb/Lg4IE/ZOPkESHpPy5ZQ6nLAMqJNpXDIYDFrLSevsn5A65KjPSaE8FCviw
pD6NiGgsSo7Oy9r6KfXGaAGnWynQcf8jERFphvMp5fWWmIChdn2KN/NWD58d7xti
JjynwEx5P+6e/RzPaY1I4QghgWdCx/q0kmC/PzZJmWeCvJUAlc/j7vgXEyFUV1p3
1FK80v5O3w/Hi5Ezil/e977k+73JGcO+lkXOvs+6ytUAxjsRZL2qejeZWEWc4K5v
dR1TgUY0iJmPim0a1sImJIJg5p4PxioDFGiRxI8W7tNiDqA3J1PdsmFxE4HXWvQF
Lrfbo2yAOrYi5q/BF447YysNTIGwxsIUNJdb4xlUbrqtGWzPx6BBhaIbiX1aQEJA
LY56J0ryzHGGpHH1dPCZN+vyQO/OiDizqEDGMsMjov9g+YepsffTEUOGbLNwGs+2
cbKxO8TLk9RBl88k0tEB8hPi5b3Z2i6nWZYAAyN7JFiUJX+AxvXILOXZMpuLME2l
wHBshn47YVqLzpB4MO24bOo5wlzExIEVO8tYlpYdVp2T2ErDkHbjYNJpF+zYCaTC
gao1XV/u7o2evTtQcsm4MWzRN7xqCdQh24FMQjndYnVEEwA/M3ok3nOCKe+1IzPe
gHVvv8TpTi+q7famMU/ziBTdvla2mESYRQHq8VMFXYju80+6b5d7kjfv5Wyg/i8r
E7/o2MykKE15x4f4yX8Q3UJEX5uJqA2HQAo4SkSc/XBhKaDpXHg7EV/IPeIR/JvQ
EYS4upjicR/r+MCq0z7tYwsu+BytS/b5s0pFSUHASA12PP842qkEA5yJtGLzUVoP
Jfcl4bW5HKI4rtm42uhBsF+W3oPok/cZCA5cTQjTP7cMUUsHvg+hOJFfEt1WJUCA
KQmULSmHtxIHFp6X+s/zaIsYU+7AqPZakmtPOaP1r3joBPv2eMSUXCweree4TgKC
WdO/QQqJ2qyiekBjiLwASeOVcO1LK9fU53bHCrk9SgXBjNrcE0QeDEOHQtYSPu2z
WIGNJ69gAWf6aM0stsbWvR26cdtxc5JzpDHrNzE9uZihoM5IJsNr/f1Z3MZ3mNh/
vilXOQajz8A3tyZ4Sncl//REUB0G0FIiCbVBCS0eEL85W4mUm9WnJ1Xk3aeQMAv3
eik8hlJqJY+uA81tYvX3aGVI0mL8Lc3ixpFvnNurjZR2ZBS9nIF1asxjvPSJ+4Jl
3ItLyCbS1/Z+qSgwzVe5LcQTOp01WurUy5kC4y3mk1LqOUavZHNJ/C6a01pYcJ1g
bwH7CqYD5qCfm+ICFv/IBbTNbt+8LV/oOlO8x/eWh92BJ9n02R3OBXHUwXNE7kq5
Ujb3Kf2Wrcjp+1KnaluYX/pJ9wMxEY3sM2Tv/yqeqe42dvzRAeQJBfWfrosvzH1u
tet4Gt1K1U+75i1lyG/FfDRFoszokNW0yB0DJKUgnulvQOCQNDkxXqlZFAj4SgBD
S6foj2pv9pO41brfbaY1qlBeT0zXCJzENdS6XIge4WO9RMw/omAq+aZO6ANI+VrZ
sMentlvmDX3aP0XdGoPA8PISpWBsW70WAZmoIrGl7u7U95KrwuNnotEXVk5kx9vE
GpsbxosUi6drTagZ7fX3BAlzrK2CUAfYtWN/tAgHcMDJtSVTaNPWR9TQBcLTdhxE
RnTXhZnNKZy2jE0ynLslMrYXrhEKD7lhnLmg7oy7rgYLBTmo8sCZzyebBvdI42ys
KZbPlhGcRxek92PQCsoZPBnbZdlGG0oEN7HeWTiuUgIx7s3wSgN+QW1NWFHyuoFU
hz2n+yE4SqADmlTl0wP0GB7JA8RM4srIi7Hqbw7MzuSez99ZB/A++PH0oq8pSgmT
gdBLNKo9t44vXGb8hFOTrT5Ws+Kd1pVoTU3QOCQud5SnDrpn2icmO5TCdt84fjMA
FaCefudoCb/J9pLsnXBs1tqu+bDQjiS0JgejBa9VwhmDWDth4OywZh+g6j1KemCk
KFwrEplJn68hxAD9cm5Xp0ZBOE377LWbbUOoFtuBTrXku5mjRbJYPJ36tthbBGoD
6sNnntsmihNDTcyxhdo4eO0iOjZrVULiYZnb83cVDuJkuXN8+LbGeBMTrJWLwIdA
nKBo61YTiUQxcAaMFxzwzU5vcZ4NLry+xZezl6Qik0NaH1S0E2QIN8GS43sIOsYL
nH5r4SrIIPR5xrzafwCGxB4BSbBHmRFmIr5KdrkhCVs=
`protect END_PROTECTED
