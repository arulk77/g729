`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49D9sXF2TjCEhh3UV42YYsaepAmxJ28YkUN4Y9KDFpjg
1Ok3lc94WiKQtGhXRiLEBXqXMYLtkhczYJFQbVPCQBL0EEp5pP18AyhQuvWhlq1U
eauZnT6vyZySM2awnHXZYH9zEW3i8YVhV0DEnLfY6EhWmqkH8cgABvV1y0CGMP0g
BC0G99q8efLeCrnV5+/slJsDurSNV2Hvx3bOSPQMUA1mAh9wImPy3v3DUfkVGgup
7tX/hxGs1mxbfId8fuSjMGzIxtP0N3Rh/VZoQUEvs6jNXCnn5dnQ3nUHFQmCMz1q
HBtDH7OZ3wHJlZkWvmmKww==
`protect END_PROTECTED
