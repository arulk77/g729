`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SRlvatpfSA35o1P/KlrKO7FsEY+y1Az1IEob1XuWcWUQ
PmPFCKJWxJRLfHfuz9WKgj+5gaZJphPamW7uT265vFkA51yvc7tqjOWC1jyo4vrN
MT1EgThjRJAneFHxhuWG3hNjHaiwWEhnkYeGCvFUd8DSeJMOxDwCPMqiQTO2HrSa
/p+KgGygODigi3wAQ2GOyUeEQYlRk0/eu7hesufl8szm435wWFX4mmyvYjVRIoQm
PJ4WM0s5F6OYQw2cMOEftDQThs/J6SV/DTOdmKYGRMCqz5XjrU49fFO5ZSXuig6H
c7sTbVfKl4ats/CMsrwKcYlBW5JT6xe3Zmoh4lwwE8W8K7o5T0ADsytqby/Ff5Nb
NAjlczLQm2JVkqV659orwUHjK4HN38ytsQlOZ8zg+cWzuDRntM112lSVUBR9lmw3
eAZ8AY7hiDE41V7TqdXiQadKrYJkN3gd7aCq5E/wtCpJP+u2q8aTGyVMAz37z3zu
j+B4Ak3bcNHDq/aYtqzqGB6/lBFRAy9bRjyvWq7oou58K3x2ErVo8Fyj2RRA+968
pqlZkvgy4VAyQx2VkH0G+P+ADbSPpcEZL7JapSAvxxKRKpFTjTDGjfctL38OjZEK
Cq/V0OXJABKFv1cLHGfMisQbB2PQ0W4Q53scz0JSjcxr82wWhWDxJ+cpOc9BiwPt
cIy6aFC+lpeqvcbWD7SZQwmPtYVTSV6Q7Jr709sONwh2lOEzoT0BlDouADidlkcq
dLBtTktADuM0to2vXSA5RtdlpaYNPahBVklLkAt6Nqt28MRXOZjyQdh/K3oMWVVa
Zy3lQf9eKGla8LhfmQFylaU0q6Mp1ZKD8RXO9jbNoCyz+9X7okLW7DnW9AjDCiWG
+sTOhwNwqoUZwxtzeBt2hiPxvewZmXdF8pyJA/MvRgcJwixvuK3OhZzeoEEGlhM6
TDrGHT2I3FFfiEqX74QphtwyS9jgv3de8ioC92LkZ4fTdN7GPW8fwnSMy37+7OOL
Wd6ORkLeWCZNdx9zMWGkDE9x6YEbnOv8kE8UBcZOC9CDMfb1NfW10b0zTniT+DRs
31xrflRW5ucZ2SxMtQXpcd5Y4s08EKK3iXUBk2KVl996SD5FcPLF4et3mlkjv4ac
HbdmRDHdL/Et804tIbJMZ4kM06fQOIWNal7ilwvWTQEheu6wdLZx0BGTUnAjOLVf
DBTx/lOH4a+IAOWKGE9NeQ==
`protect END_PROTECTED
