`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIGl+U5CtmoSifXIZCcEpRQkj7sgwbdea1i/oQTm8gA/
WMVsueNy66V7z+WCmJ0m+ev9peWPLZn4IXMUnOplc1MnEJfQIFzecYVsnOvxdG6s
/pQKCE41MCaWqeaGSE+jm7616R3Q852kPv9EfSGoiwR/nV3pn/3/C1Xa9tPKGoNT
doLqlXKkUACVRjsCvCPQiYWhVjJs3jXwJtcRb9tXYG5JA6pnVS6lzMf7kb+wCigx
VejbzPh9BsqTdKq8EfKi8OZNCyzbv9j9515RYegVixwyCWr3iscWhk1LVtDuutsC
7yw1jdBKARkIoSsfonUm91oV75bkNdhs26p0ehRj6W5ioUU+BhdXAjC3YVzJXycj
cV+ZsBwsvb1JGc5KSbsG+2kEKfsAdnJioeWtXS7FEZXRJ37BzMz6e4ofsEDGerZt
XV9JGXEPdK8BAuCANjH34NjDcD6x5VDPqPGQ/Uz1ITQ=
`protect END_PROTECTED
