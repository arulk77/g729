`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL83TFqqM5JZf1WEt2arccWJdI9w0QBB5XCVSdJ1reUdAR
ZBMVVuWDqPOjEHvJ9eChVc86mt09QCXJclsS8ND/lVd9//2KQetSVgZTg5+A1wH2
J1Z8rEPuHwCxBOeIGgtWSa0Ag+ZHNmvns6snWLPt3C/T3z+W5/kx3ZjH4cIRwGZa
iMl5Yx43AeOcX0mDjhr2AJp6XukXyUF83/YIz5HDx+35+eJmT9NXluZSJn/E2Gug
GTEIM2fo7cZxhltADtroWgpx/wXC80Z8hAO7o0oKxl3UsmWvEb37i0WWo2ZF6CzU
fL3Ik62lGVWenHTAieE3sk3iOeYNscrkyDsvieezU4i3A4Oesjf+pPSt84/oxRr5
Qbiv/tRKxP3qTTTCHCdNFUwU1g5i7PRBYdVF4p02zu3c/L6dW3qZ4mCxKqooFt3S
nq3lsbbdJaeqTRPj3t7ch5TPlALSxpW53LvKhHimL+M7SWBe9d+woh8C9MIuM7Tu
6N6W1qIYSscVqFuLMawwEHnQnvwcYaZEo4OQofgg6zmuwfRQzawWtFmAftLNSAid
48h4+pZbfIzmlZMNqnUB5XQ5WxFjK/eGrK7pqi4L5kF4d9i1V26ZGC4nHPd7kMXH
9+dOofyeyjt0BWrdrXfc09Oty6byk4KrJeyJMhLActvKCRy7xFqGx2BSVsa1a2DI
sYN7EyB33k7tuPorxXXvOPniYgMhbsgeUbqxqcmys0SOHyKBty65vmwELmLcKWte
BANzfW7sa9D1ZwYL35AcHrRPeuqbZGby6Fo6iV0lZmiXausYPTsusMQORlxc6Oxf
22ERs9YoGrcJdxa235DBaHagrRmhWU35hKUPm1GhGNNJFCRrbXG25T8Dhn9SWSLO
wRiQGIFmYPFjznr2VBtOTK0I4pMCyWfKVQwBpkOMvbEwofY2aF5cvDiVoV8dPfkB
pOhsecAgUIdQvJCiCjz4QqgezwOBacoXTsnu4wPhxNUJczS8WcGDxVdsVY1HDKAd
a3slPDGr00gvzF31Ev9Xx6kbaaNQekYe6Fh7F6xZwiDuBeP8cq1NzXfIPStzlsWP
vCMeq+npnQoBNwuFnmoST3tXCrHeowXXl5LlziBK4Me1JPvakIANyO5/h0el4aHu
yw0Mg7vuU5gZ280RcPxKE/HY1io4ef42vUl6gfO4MfnSaGzPD0a3NE1G4+0Ti1lk
3lvh5E0TDthmi2ytqDFaEu4Lf9Mwb/JaIHy7/gcCODoVXU2IvtOfj+Ue7w9MJpL8
1L7JqIm8UNKRRTvXuMYTWYLBnWxs6CUjBPJU3BHWeRL3pxY5ezLaWuCaZHYgdZDl
suBqT870wRYmwL12FRJ6X5yW+fVscHISzuUp2kiqmAH9ZH0E2uKjChvM7+UuKe7m
JiiXbM0oAK/EfxzfdgEGZZFtKLLLzFL7sW8F2LsfB7G/RT507xy+W6A0LWBJtmuw
uwUh+pw127dWRInGBhvNWyMG94hqI9aFIJmNi+PHCyuOLBKvDJi+WJ/ZTQLrH1hY
ljvkbzADfnUDvGhclzJqnoKb9jkm7wIB/kTEb9slfKLWf7zxpUIR0pu+03AZ4bX5
4hEPs3wV1xvvsZ1M9PRfxENPLkgQt/dKRdtKC2wjZLKRdz/gdwzn9MtiOiqLT3Xa
96woRhs3rXXM4FsdeHuQW0qMj1wCBPlprVuRMYVjoRvvaJJ5AYXA1bkcrSzWwCDu
OdtHDYjDIMdEPqxGvE+qZ4m+56hOZlaTMeLLR/tguiN/RHjyCowtojfRWJRp3AZx
f/ZHOnPbsr7npHEB3tHtKg==
`protect END_PROTECTED
