`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBbziyzzzQb5gVL+RLkWohGc/jfxjmSZQALipU2hxWAR
0BCFiuFWwYglqM2St5/SA2xSRm7KFALzhBA39/5a3y0p2HTREYSxBdnt517JHHnF
XBC4NnF4qAdamKv/3a7dUMW2ZHfyAZHIuppMv8gf4/GMkUq2NUc8381am0GADR6M
c9Pq1If9RgxzYaCi7v8U0g==
`protect END_PROTECTED
