`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNmUhaqfAbyl+2CnbLPkSwCsBWp6shcPpIIcYGNRt+vd
v8g+3sxHcyq4QUyQaZ3a4rfI9YuA5gol5A5+zn01orbGoOyj4n0wfOVtmX6jpBpV
jB0EFKecgiEIvliY+duMX5wWcQ30PYP7EXiklzXoDi49eX4RU/gTacZCKNPk821v
ExEX6H+vO0keyLS0qI7oyZk2v4MQ9L2eKFAxo7nTFtnWq/3F0qv5tf+pl6i0fEyK
Av9mG6UEk/HXYwezmh/dW3MYTu2QmCGybEliOUM6iQbhkPXksrAjQ8x1W09P7fRP
5KBUCxKAbZalYWdXYDl52/NephSiP+rimIUa2jK1yJaYNuQJpOE/v/L74CfHGZtx
REmg1ao3LJSXHzEsBt7fHXOF/AqgiddLsfFcDvTQtIiLWC1EwTeYoOjUoRJoKxJh
0LOpaz0rKJ9I8ojJeP6F6IkDyRZHBa7rIn1GRxKhXE7eaHfsXqO4rzfHb/FTk34R
EvroZgHg6wXU9wqPbLuWmM8GvUXzKcfBv4PZizlhB+NvN8EipoqOgpvIU8s/wPjh
8UMnp7s479PymGV3aQD5RX6t0lhi2lx4HNnUc8nMYkZLfiTYuPCPxXqLzoaoWDBR
JVpaiLRO6aEsY+hdAqDvaCEgBgs6YwOlw7Z8stqxRlXV7qKUeS4Jm+v4cttfoPUv
PVgpNM328vcyM0PJ4x9HjdK4XijzIIGcJE3mfuWd9Y/MBDRlR35vjzAKMsE7bpnK
3lgePf5uo9NJI88ClzzYGNdbMcu7+FC25YT/c/cWs6MLNxxAxaBFedXumiQPkzfN
qn5jGrlMiZjYePOZMpSfsTDCAPR7bcu39gP0eeQcTjw=
`protect END_PROTECTED
