`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNzBxBPDJWR7F3BWXZ0SXh3slcibZOJWwQzRZwVOXgHb
QnltWIun/E07hwxt0pVop/5P9DtcQQHF3Cp1b03nC2bH6FlrTl3uEsgKvvAVXyKj
PFUqj07t8qItkovUrY11gQyIypOGp07pCyVMRGrBMxt+A73qcNmWdF6iag+VFXhl
/pfUrILy5EIUpYybbWhQjA==
`protect END_PROTECTED
