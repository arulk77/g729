`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGcUyqylSpOpJ4gO1BnOvvqkNqkYT4vtkvKRGHgmCsSu
4ELsa5W2SknLdB1VZVnV1bPobE7/pVCYXLufYuIl1ZCIZYsOzGf9xmfyVODVnkgx
cY9dbNJGJLBps4jM+GfrzRpdB1p/SSjgrqT+ki0PN71C5vDK5m6E+H3bnzlfBL/n
LLM/tj8rdmcA3mXfqBlnytobiz16j+jEOeynxHvXAT659tJ1SFfi58qTbZXOPxZ0
hmY+O0tKDEsor/wLNeOZ2WF2UxF4fCuKAEJGiqySAt4moTEZU4EuNCV0mEESimkx
7h2EM/L6Sp7lYPxVoBZyV4GP/DTNLEL51CBvEpXfOut3BEQQMk61cBf7cvD0mVV3
lQEY4Q+20ab/yVX0Vd6HI9HyKt/pxDbRLpxMxsLRk84gsWWAxyE4zowKqMf8wQEy
i9/RObwdJv6pcj7CYDeCs3zAiIN4kay6kwnwK++a5HWS5RUBh7rYfStXpCgViOAF
A4TCUopKq5+ySI7nmmzgsXvSpzYpIrLRcEIFLV2k/uwvS0R+nVa71brJ3L2q57nf
fzcoHYSV+Vhcx8n+5QcQEH7ombmnsLFclIP9MsuzZ0Wud0ucURTE+Mtpu4/O4RBQ
9X6XYIQo2ekF8Tt+BEeoDrkyBGPhUrilL9D+xlpdCzHw074lEe/inFK/Kg6QKtCe
`protect END_PROTECTED
