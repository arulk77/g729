`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47bfB5EBFomkbagNTKmKEQsUUQE2MFLVpR1dmkM52uUu
tKaQVpD24H5DzKFCwwgHt+jz9KNAvLjC53FRqJxS/sicvPfgr0THjJ9xuT0TnRvA
NP1U5y/0e888IsIrUn7k3+TukcKVbTZORQ+AbirLUbkynr3ZTsylm/88IpBORyHw
Lf7sHgRcJdTi/B3qsGWy4wd0YwslVpx4zDxOEAPNV7KeHJu+C47gP7CzXmK7GJbS
QMuFSJqtiWCT/SH17K+fUV50LykC8CazPozUeGlEw2InZBFGhSo0tI6yXxs4BsbR
OssXCO3uBtTbS+gnE2KquOvRtqNAo7ALogOhYr+EzunLmfTMP0vCDgTZE9uyz7hi
uyvsBLOPdcl4U1yZsHcuRA==
`protect END_PROTECTED
