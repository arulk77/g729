`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEHYNkG+eJLMnibie3rsLcNFVOE3Sb/b8ldhKqWQWVT4
DeX1lOl59m6dK0SGXiSzxWlidXQF3iu78BzLstpKY5XuFQjEGkgyppvreXRVm8I2
Tysj0z2+s8zzBmSZGlDlMuv/5kP2RPYATwBYTnU808gsWQz4NHZPfjL+SmKev+MT
CCrx5vGrKGLDKbPdsctKyrPhHkWN73lEcvs4uHfRYYRHdjUGS/o+7l3O0g0czH8F
8rGYuhlpQp0C+ddOrCFWHZMHT0amAt+F7tnnmQULaNz0d6IQWQ0gvPIaBD+yM3pC
B51DldAaIiq2MN6zcScOaFr6c04CIn0YHMNQvgIy3sdMDHz4ZZvwemBlKgMtwxYS
19agp+L7hEhM7LiPmHHj7XQtCU7R9tCXvdTzvlifGu9jNnZWOYEv7xI+b4ZWzJML
fDDc7gqqK6/xWA5EK2ebWA5IDVolEs8ZrrXywzSfB41P2ypseqp1vcvQPtMBfITQ
`protect END_PROTECTED
