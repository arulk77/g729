`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEtp7yA08rOb6VevIqIs2vDKhHiP5jiHB/XEvDal1h7b
01rswk5/ve2+UxpnQlW+/ec9EjeXw3AIB7rBFtO97dZH4GBDYk6tQFCwN2//gKgd
H2/Z57S/8//XzMU3QLYcrQ5Ge+Dt3lq/AaKkRdh5VoSLrC8BuRtRmJmE8R7pHC8i
Cgg7VS0pbVX4R4Qvws5QDCeYbWgqDyOqCU9EAAYpSyOC45j9XXMkf87iBVXLy4s5
mgntPgML5kCVcvAG58j8m6Qti59J13mslLG7PjjdhJo4S9WpLRPRhqfkP0z4TlHH
mhMUyGLZQE8wB9TWAOtqsKmRSbqZ9j1lE9V/QjJXUtAms2A3czV2J1q1+GKvMpls
l+YFK9NcXlxA/T5fzwAkFw==
`protect END_PROTECTED
