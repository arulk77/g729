`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
b1jTVD5Pt/SRdmnwbHuSsNUO7XS+YKleoMfeVtlbxEPKFXZZWCdFcWsIHszBYNNj
DFrt+o92H1R7Yt5frWb3MKvjQQmMwl9rwdY0k0qCvjAHDnqEG1wccHSTphdx5lNA
dQrDnuVPAXzKciTAbdknoPy5mmWzKJYecq9dw2pJokiPpcsgOVSm9oOIhXSDB0AV
H7GV+IGE5uTNJXGTHovc0Te4fjbA4UHq+PZG+ZbdJsFIV2HNrWF13tOtFr4Ev1mB
mBU8k6qO+ue2P/hCommht48yEGaaCgoufPtN8niWUmqAQR9YkXhD/9yzcyePOwoH
tFrWaCgdzw3EMQ+9teQU4LkTh8DkEOAMZCZ11DEZgG1kXh0q7ZGlAFE22AL2/DeE
T+1fMIGRXo9mHS883iYzQEOhBhH0haFyYAdaVp+YAgCRvEahwF5btKP/FsuDyQhn
xDzl/bfQqt3zvHsUMi6mioKZvsp9Z3CrPWpJpW+a7G7y5JEiyBElOiUcWLJ1Ot7o
3nvh8F5xS4xFkwUyDovlBd9gryE7w4ZuZ/f4Rig3rAHX3EsRzXTilK2jOjiKxL67
qBabgLqgNpoA9TzwYC7zjrYDOCkfq4TbR63z/yBjOqwUc1P1848LhPiLmmx257Zf
/FHxPGu5SEEAyO5qbL0J9WsDd4/Fz2tkkIu0CBXvdaqOkLdIRNky2gb0/nfXtiKw
hIQWyrAJI/PCXW63TcChIRh8AgvCJiHcb5P1jdOyMVU1HA6EVimyTbI65yGTsdcl
GCjVxiKyVPO1qxIp4L+wCZ+qAVSxHwdcU5ObGw+rbyai2TyxgKx/Dzyi48+DBUhB
NzY5M4CoCrrKVWpKFoxYSQ/LjqhXHoVQtUMPK9A0H1VspoUk3NAoM6JQ+UcZqKXB
UQGTf/pXyiPlhRo2yxKhBVCopfVTiazh0WxhLhPrjwevKEOQ8N79a7cPr7zCrlns
EerSNQ3dBtv1+/tVCSmrcdd5WVuuqz2ZI5L/Oc4XP1IcR1RYVXarMu0gtO+QwQDL
/KbckmjAm+7kPmLXTP2Dp55Dp1QjFZUqhxQWLQHZcJNo7q1dBSosdw+lXjWwz/Hf
RDD6fzHbJ7bCxgbdQ5Ua/eCyz8GZeDGu7K8NeyDvL4N+/7QfXw9ilf7NrQtjwhiO
sbFfTO5I9l4XwotYhn7flfiXC2L2DB9+fZG2ufOhMP1iWW0i8nldltEkD1Y0o1ec
GxUXY7qvFyQiMEu7Gef4vu+FUX1gJL4Rh/pDbsKaAGeAbnDSFa0GkeEa/9uvh01E
Vw6+uLrTJgw9+QbL83AvMJ6PAx6alcGc7gwi5R2BquDGTFu3vbmpfg3KSgOevYXJ
7QbVru7yWxa8rNcTcv8h7pm3lDzCMeDeEjHCWxkR9T6+rhhbd0PyAY987GjfNuaj
VEDt5oqrgFzhCR+/JkglTt4BtQ9J74G+XwvynBYNZvLTgmhGcjnCxklNGSsPX2uf
j/ZB9uy38OuFuVDe6ERclSqYqpPUeZaSNKYLuCKTe87cacfqK1Jj9YuosV9kqWtA
W7l1fKbHfVzFmK2jDc3HZiqy9Pg63aRTtYUiLinj8cZcWnP+xPLbtsmkpjPlsPiF
Br05W1LbEscEw+CNKSnyZvGPW5q2kwwvIaP8xREqO6KatqtCHYSJAK3vI19S6San
NdFZASyLNAypysb97IOuGCViZJnYPxItNKVxdWkBaUCV4l4KH+EzvUWpequyV5qW
O+VL/S551N3f8Vnu/72/9o/WkTnTW5voo+Ptqk0naMDP5tUZJKYTDPe0K/0clv6B
bn8uMSsm7KpKruDfdW3enbC/zaxdDNFVhoZsxL2ovRaHA7phB3dvktYZyr7J/66C
6zHCtQ+4P7TW+750qS3NO4v0PmORRHPvvpZtpmnTMln5Xv9c9mvvmEezOS7BbCfv
KBbKz9KRQNq+JFcMaLpnarsBVP/QgGsn9Wnn4G759qdluh5OnTmTAtXQ5q9pM7Ag
ryWhCb4RvZtdeEqJydCu93HpeeamqYA52CBkbzUV5CPe2ReU9YKWH8dnGcAKWsk9
4NkDo9b44TZXp3YLDzOufWObptb9gTLRw4HZcV4wOqD01/V01e1BlB0dEOA7sX7f
KwtFihpcx8aEACjXQPTWmvTBPmX1vTNTCRBy83L7XMC0GvvzsRDlUJkyJ5Emv0+A
eo9BzoxvwBUPxm8KK+uCK80Me4PCaZ4YCTAhhsWeqNvtMTDFeRgIHzzZxI+Bz0+8
ofrZ0S+ubnJml4SiVc1gfuVnZuIR4l2LW5afXztSioPlKeM99pYfcNxC5P8bOFSa
8CUWCa16bQMmf+1LnuyUvmd72r6yiMTx8C/KLTLHVYoQxwnB6adZiEfgNM69Vxo7
RGJ46PHOZcJDOUNWlp9J3awJbcwioiCUaCc5dIDTF1nMQ1VCVdtdwPNCqsHjqIHq
9RKWf8x14PY9ms0c71KFXJVG7ksvqEu6IkclnnYXxEG8TGMem6kmfFaNFu6swiAA
TR69+mxO3mzzqUBv+3CuiqJLGMR220lIOg+CNum3hOJcvJCdFJJhJ2GyraqOM3ZO
Tpt+m2ztsaAC0cCn6vqOi9nzmaPy0NdMHONCb1IAS95lyncHBmA5vDl7fcz0Zs2d
Ks8KCmtRyPyIQ5DTQHXvZDZLhwpfkxM8r1P4MqtoXOhB6d4dh16Tcy4SVG/dKRw6
5miwhY/iMDiBoWC34T+T+rmV9Hmg0FunRHQ1UNuc2lNQkxy65pwsK0zwLiXBj7Un
N5mdasmlK9xMvSwvTG1tnzGvdGSxozzcppr442bIQKMbBFhIYtezkJDBliXzrvWx
If30lBIBDLelgKnPClUgJWUhtkGM8v4a4s0vfzsuHFg7s7Fic3hzt0evfkX+kRgZ
TVMh6DUyNuK8mqehakdKsqvxIhJGG8LJ5AI/yT0NdfASGZUQcokhL4i9EaYXLs94
Eoikz6Oaz8bgw3fFaZ4wIbNEFXuNJKTtqua18knAidYDoSdibFFv4nc5YejH0EOV
btNtgRpwH9x4cR0SwbthAGiPLt1YW6OuysckBFFRlFQ=
`protect END_PROTECTED
