`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMec158l4G+dXVEHmHb8gH1O6KKa1/diKlVzr8aWj2A2
Tuy0fXR3W1K3ymNz4LuP3QN7hGHUzrkVde9Ojjr/ISxk2zyxix4X6OAEy6+SZbnF
d5RbuB5hsr+fBhLXwKbsd+7w5+lHQrKpPBqLSk8GoaMGOAT+/7ryo6igsAapn5tf
gPzoSVB8OIH8SUfh0a4Bjzx7OD6aRJSP8/uWTiwOyeU083ibRVts9KDEm98vvIw/
`protect END_PROTECTED
