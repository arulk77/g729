`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
YhWfva1tu17a6Ifbs48u1iSizIUv2JxdGvntulELC/kKaJ0nCzYU2sTCrOBls8v6
L8evE0TK3I9lFS5K8tcVhfrzACiNju9KCHhE8ahA/jBvJvKPAn9fWsaJa+bus1+3
jsiS4Gue6HjekHJTQlS0JVXtxCBIr4NY52yuSbWEMJoGdJUYzlyrAbemk2+uOD1f
LbMvk6AgtupcV47hLaZGMJsgI5U8G58wIH+4kvPhajOlzpXmBqKrpnpnUZ8ACL01
gSec5yqEUQgU8XZfivDOO2Vvq2ufWKx2tCvevmud5WXcIDs7eyaai6ISWUVhK1zi
39Kl+n9MZU3tJDyquwWvWGV8ACCR52xYtNp9AukBeHGBk387TbP+Uh0GWg2ayMx1
sWdpVa6VPf6kPCrKOcxpbODMY7xqEKeY/eRDfIMiSa0=
`protect END_PROTECTED
