`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLElF75GBUyPtHvQoOZoJG5dijRYVmFLAv+tjB6QTM9C
Z3xPHx7GYHdD77Drxwoq6YnYcBVzQaI79CVYb1v6k55mP1eSHndHvxgE4yCXZQh/
OmXyMZ4NY9YtxnzkQ1mi+0X6X7Rl1zyK2Z7nfX66IhNDJFPXfmdmN/An8gep4/RH
/a6zb5wetf7bk32yyj1EEDEpFquJoGAc5ljct6Ptiv4VDVXp7H4+gkAoThfjTf/U
Mw1BmDLykmjX1iCO0B4K/BwG7IDbZTH4b/FEmB68KiH2i/UTp7Jtsw32r1d50kEe
GUBlI3aYd7V9sW+j0uJflQ==
`protect END_PROTECTED
