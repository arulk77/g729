`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHYedUbdATv5my6q5Z73Alo7pEIuF7U7bxXNloxYux1z
oWXmBUtx+/bs/h4kj/mka6I2TDsTaTlNACjEh3t3fV1vKQoMHvMST4TudKSZCSOR
shfLlX0dWM8kX0THOtZX7hFJKiemoDTF0OYMdFkfiMvRjmvgNVFwv7GfoOgzbRDf
WmHWBKlhZUsdvkKAUUb+AKtFKEPp5FZJjOpytkiZO1VD9wXZLMzRcfyzvTEkPiof
vuzqcFixH1bqZtn7UVh5Dkm0+ONn/Q0S24OqEUv5f54uAUGWz8Smo7cGSAnzpBMW
2BGJ89iHT/r798leC7eDBpMeA+SXtRiW3LceXOTxeFpFiUI6KR5Ng06GHLv97Utb
dne/Y7lPsqteYOG3m2eedbJMKjzp7bW6QBq1np3TGEVMLv8YqdCznCh+wJ8YCGqk
ZYukpUnL3UTGgmMMhjANaGxhpWLhbnMRcxg1R1Qev7X7lnXYS6xYPOhy8DNY8Bgp
LZG7t+C3i2aiYGDSnL/MdNuxhzAcCTOpJk5x0KY9AMxqAZnhYgJIP8+psn4Wtzs5
1yaZg8U3pvWxn6iXdBW+LA==
`protect END_PROTECTED
