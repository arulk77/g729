`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAm2wQIjkEXAmr57Qs8QO2Aas9w4i7aG5DDwhLzQq3SH
Guvj2OC+bBXQOatS00PUsbN/heHYAIEfDQ4HNA5WpM/+Jo28ivgRWXsXtuAc7E59
ippbtV59uRmweGmBn+vgYbOUklqw2r9tuS++KmMowTmTxWLwW74TaJo+riVLSDvA
f057C+Qrb5MW86BDMU06zO/xAuvDtgUrPmHXVs59Y9R7WUt9Ti2lt7JmE/UwZMkk
OTb6hybOn2D9TxAY1J0FkS5QMofF3l066IvDTAxSmbT4d52I4Im/XzlQqkKccwFQ
xMv2yA1yAMJ9NB8siG9De1Eh0AOIhVDx+5DHiXD8BeRI2VuDme1RpAJorU723U/c
fExcO753a5bGGvps/mEhCREZjOA8DylvbsOxwONTre9uyDRz1Weftpm5ZT4X10NV
JYBBNM+rnhuslWgIjRQAozxQyZ4Rvuvo3T8mMweHXJdQlGpHcdj7I1XBGzRQG6Xj
ruCZtJrQDgAWzaSV76uTfQ==
`protect END_PROTECTED
