`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveA2VNvIXtx/YfjFAZJ1vdHTISZnYGjSQ5wb//O9W0+aZ
7zxXGYr3EZQ4c84fUkEAV/emy0M4e7p0sYnXuf+3EZNH8HBy/SyeEsuS5jvyW6Yu
eP+9V+WwfX5vW6Nzz+FRRGSJcedhBFP813qMfrUuKpg5INiUCGgSU1dP49QZ/Ro/
ZMO4VH+8IHnUxInzXWb+VzFb/kc9bGnW/SYhPdZsIGIL4Fmx0zo0d+lFLwUXL42F
ztfPXWbiJh7NNVWbvCNXvhY1KNm8uAmE77ib6n0b2GJtuyo+bESqifpkoxxrXAZg
/OlLcN8Te5DXqNvZDn7Z2WUqKwSEdinwo1fAkJro0mYR/+39nlYB/VeNz4GeEgxK
MfXv3MR7nkxEwZBCkkNnXbY4nraOSU74CTGXKd02chwRIo7ppDkND3vid3Gn2f+k
7ZJF7DSec5/pmQe+RzYn9kHeCXgAt3aGwd/xgqhS3MGw97MR0v1oX5dZmeCHuREt
AhNadn9klEru3ymeWI28fCDUGUpGceYP9E2uX2YLR/cLSo6va5m6WEFgazk6gSzg
`protect END_PROTECTED
