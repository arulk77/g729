`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ah+6FtI4W/upaVgdQjOyNbXQcbdHlUcCsy4squzSQ7FaN8aVEQ8Z6JpmmPhbQIuh
wTC/wUC9GlHXdWsmSwWNdqHd0RCBFjwxDRP3rxbh5VzPzC29a9gsRBHTYXvaVQNT
ZTU8HjftsZ3/ihOp/asE3sZ2xbWA+PwFCKM+1eK0VCy0ifcAvkBiimhrV5FIWfY3
3JoqRhjqfeG1poLeIaM/pLl6OOkcEYO6R9hxN7ruF0vebjDCO8agSe+F/OTOI4/X
67A/wE+iaQVD2ptv6ndVi6wHlb+Zm1ko+U6cu8UjdbNHKeFmUNstdZZvV9vOVo5Q
yO2+4mLWFn9y4EvPNa9ZFgrkjH3SCovY7Zua1HesuZ0=
`protect END_PROTECTED
