`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C0w215wiXUKK0oAye3asD1QYrSNcM3Oue/nb5q/FusSn
f4TOy9My517na9ZBa7TY/R5lDNow/o5UoZL3GY/QcXiNoEHQ2D7nLGy2CCY8GGdo
oMVfYrKRYlUmvmWwaPKgzsjoU67eeVwRxdPJoRz3+LlbrvaRKDvb7Z9LZ9NDmdB1
LZk9gbOiIQS89HLSmOrIxNr+TxQsc+jvgA8RDAWT1wLnaOLwiUs21Z7kZ9J5Q5/a
2VNFyn3yENO4DAs9ZkfxkMYznrGqwy8kvSf4yFF3HjMf64WY+5pSnE+Q/LRUqqs0
W98xfN4/Zhlr/xL+Q7Nefg4jgl6Rr2pyk1SRLsUkiZ8Hz5inoTdD71Lo5CHbHomD
3hY2hHw/9I6GezlVdC+1qfYDKEHVvUycyVJ5UHhspFu8bBhk0d8sNvu1Cyylzzap
lMNf/26SY4NhM19lqFVjrdAZulZhyyEoBlb3HAW+gIjHqNamXThOGtOXNKY0gGo4
KLSpaJ77gt6RtJIK/pO2bTxMyfdqS3KYbsRDzZZsgSgV/32MxWRpOLFy6v3vQJgL
vjJG4J3Oncl2n0PSSRwq7EVJI/aiCPKkdtQcFz8yb4F90Li1tl0zmkAa5FOS+z7a
p7pRe/nsyiuUw+8UnILan5ZQ8EVZ2eGLqe/uE5pQ3v61OvjtobrYzxHa7IAWznoE
NG2l7tX7n/HWSR417o3QUZ/Rr++lE1pA9IiY+8D0xlLLi6Kx8X/J1ojYAAFnaVTp
8km7i2REBldKzHAjY+tV7A==
`protect END_PROTECTED
