`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveO5FktSxuX/ogXDINav2lav1yOj1z4rJzJGgbxeRGksr
lTaTcIAMLULT7n+Uz/Ote1gqsuSZo3Zftth93aWOD95p5aGDrtH5X3iVLp9+cjIW
xrLypWH4NUIel0tEBhWWMSmGxaiGZDij+FTt5m26fO3HKTYc/KbPQBuSWQ2zoKhC
prEvtZohEZoPB1yz3f4ZrmbWlMSEy/DIFGNRr/ROm1YDtwo15OPRs8wD+9EGv1x+
CFeuC3B4kcqRh7hj/9YHv3x7mP1Ai1liqRhyY8Imk5cM8/x7psN7HNl2NPTtuAes
CN7h1AClQxq+X2tvhipxRcfZ6xwY7snzaN/yNqG0/0Q+E045WL050Rt9YqCoGafb
83aKPxu6KB5+F3Dji9r8r2hrETHqRZQe3UhhPYGCWwnCHgIQKNW/OW0F0T4lIV86
YYDmDQvkhFHcTBsH/FGiFdEwS3LDzFdo8qcLOKlPvuQ4uXs52Aiyt/DG6bXQkhYN
Wj6aEPXONtsqZU/0MeMSGGY42HesFLDzlgeHQ1XOf8dqpzB/capspTCtqmLFt1bb
xh67h1JuDF0OFkKeb/M7IZICyqfY8Naz4xJL720Dysf16SSkFs+DXnWy4Kk2CmHs
OVIFvXXw/7n3K1SOD2O7FJiq2RogvcZXP7frCEeHyoA+V6ZxBhqRFweDrxgA2mCm
bqjwU8fekgll/mbbbnXAmCu5ZLSo9HaPK/h2kJfOo2DzC0gcSJN89IrYCxF/X+84
0ApK5ahRK4hFJU7lPWa/EVzhxkAXLy3x+TLYNLYu4FR98KxzhYSLwqpbP9WR46Yo
`protect END_PROTECTED
