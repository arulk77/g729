`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bXesNfN1spFtsQWh11R6TNXh7Zt4rLMflJ+D/KOBgxOyRtibRXremQx9OPOd1H/v
tdRDzN7aWD0NfNrX8qg1vFJszPcvLqr26JO1x0rwN0blhKmsgq651YBFtsuxa8nH
t6poGpoFgRMs5zN7JcUZI/AsCkcz36Rp+Glwp/rnovRidjMtyTWa8Q/jB88eSGSe
pt3fDGPD15YpUWosiPqlpUCEJFnf2T8W6BtSWhq6G4bLTeEbypuKXSGsDp7rj6K6
1EYCWAVMTirAsiLt5kD8pJ5asBBAPcToDKiHZxEzOJSS9uNpSHBEKbl2Zwm9lBPi
nKnX4/8B3LeeOBkLEG33AOJboFMc5Zoi7lzZAWIsBlcvcbLzs5u8sXQTbH/a7Ptk
6cH+R0GbJEtQQIU4D5R3BZnuS7q3pkyU0HibxzWZAj9hgoEEUk22Y1M3JvwGvt1S
QBjhVJlYhNhblaparwbHsziyks4ql904/tZozOpuZS/5hx5brCNp7K3w8DGip0ea
cBxThQmCp4oSUfSVrKReDgu84Fn+WqFgTEcXMgufNxq6001csOszkvfkSt5mkvG7
yFjYCBikCahJeoraysTeolaCJCAv2EpY4XqxdrSamWDQ8Vg6pT8Z5WTNg/lipI1z
40BXSJk8X/+sVz8p9/i5cT5SWDkZjrOlWqhBDL1+5wzP3+YZjgPxb2s83XLsWwvX
pHiHMByZzOKAIJGeG+PDanxq7OAc1Bij3jWt3vWYYfxcSiFQHbipuyP6i6uVUdCL
ossYI/70qqtit6LCzbAnnOzrOfDkh9dd1NPzBLvHYaLuYVsb0dQMzg0Nr6vxM7JD
wv2EZEAB1HcWaQP0mvJ5HJVbzZzZke+dcesCMHs3RCf/C9Nj7XBgQsuM+DyqlhHk
xHyfGTI8epylnmS4QG0FhGudihFW4bOxEFON8+WS0OuLMILPguWQioep8j8wp7Wy
syveBTp2FTCueiOkIP8UUwv2CFQ8SKqHnX4y9txVAZ/b+t4ANbs72HzjS2pN6H4l
Yfqcf7ueUj1F8+SbPlAfvd4uBnrMCrWBSkhbzC+HlEMqN79lyu8gi7pCyjHuZpGY
AL7DZxhgt1YFONdDP6qp4z5MNIjSkeU8Rm/OE17WkxeQXJEkkENxp7RGCBE/CfKJ
D1IcxIiMfWsGcNjQpj5Io7djJjNNYzQ1AEo4mH41Fxve6ddWOwtM5n90C4rVuaV6
GXdPdIiMuCqbuQXpGjwR8BhawUIJw8kW9cAWlkQniepKk7fG6u9Ko4azEg3c9gPj
BO/QTXB044BQhsAVypwjwpnWv8yxO60cniv7mPtIQ4VD/EbrW9+P44GVIHXP5tpn
b7aktedpoW2+18upk7TuqCWIjqi9PlwUvN9hnJAmNHwvokFZW/P5DMXaB1EsWxm7
fi3EbxBXh/zKfc8tY9WeU6DlZN7dEW74iIZzp/n1RG5h5+bIlfPAHifgdNoRnLqI
WSrtEVvwtYj9Qs07qZC/qj/TgnIY3z1fdhEwNJyuWLXXZ+Cs0RW+h3YqzGfSHT6R
t1fgRCqABla+BH97icD53jDR42MYjZfrY42/Qnv94HdsbVEzusSGw1/aA1cbOvdX
aAN9Jb9eO/pK6M/z3Sx9Qq33eKD5p977cMBMQ3lVMNChSBkNmr9aNB9luMKVHLSA
F6qs9JnRwmVYtS/zMWaAu7AnLDdZQ94Na/EIFLZup1E7/y9UE/Jm5WtY6zN+qCkY
LfksLurM1O0nGhaoIYn+NNkfB52vMDZYYhEsOh7qtNZXAKms8a7CKS7cARfWyJh6
j7R9IzXds/dJvvCysACXBPYcdwu0VG1bWzYSK8rf7TFwceTiYaZ5BWj+ss806jN0
3Jn774QSGDPB2mKxususI3rAHKmGUmTu1S/gCA1Yt2dbyvWPPrsF7Mf0U73OyM04
ZC4PqdlDwozbRDJtDdE9uC33qVgGbHRZvHRn6uPlo3GLrwkhC8UmgvMDyTWv4PRD
xkrnjtpAmA0tztdOaed8gliLeBk7aIX0UgTtBHXlo8MKL6K7Nk1sM5BQrargRqLR
4gDPIKeTWnuTHZUnfyFaxBs88/BjPDLRTiJdGgpMgtpAF9calrEciQG+qd/2UM47
d0GiDny6O3aVm63AkjiET7RuJUI443whXsEo7iH1nsfDze6xCfAZgImOXIfJDHPb
6UmIg8l6mfZeBsk2bZKv5FNmCONpN4jMnUtWNiSEMHE=
`protect END_PROTECTED
