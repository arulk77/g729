`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePc5HEI6KtdtpviJD2E2nhGxF+DhwTXJZSCqTDGdG8za
v08PAN04bgCrle3LELysaZZSdQV+Ex65zoxeDLexQF4JfgQL0/EhSLfs1/6gR1uI
1C/5d8+rLL/r+mSO2qXfkmmcxaUHG5vdgE1LKcnIO5OkML1P5MkT6ZiGGKIEXK1x
2Wd37rLdCAfqY7cT7UEaVpRrmrl7jd0RP1obXtX4VzI=
`protect END_PROTECTED
