`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEUylwHEYJBminR3P0bocX03o3BSnzSKBMwSw4NrDsnE
sV0mZqVVEl8XNTUx0EAvqTTi7AblV1BX9+QOYzGlHpPvbBNpL/NYZyd74QxosrMe
ZHOtLm24qw9etZUtntR7k1xXinMuLmmwwdWDNxWV5rHvft4EQLkRvzUpOQf8GECS
C97ZVe9rlqWI5rEHzplKgs1hL9zUmnwmffxsFYUZvid2ZPwCCUp8xFEWUF1d6zzK
xo/nGKRlXFeHrm6zOVqwV5GKdzBu6cuj2ltjL+jahmgGbboXfnn0cK1D/59QRMZY
iT/L5tCgm9vsyo2ql27ajVCt4KkDyZNAJ33Uqayt2oYYugZ0BgcK8dR+yOB5Ca9g
`protect END_PROTECTED
