`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
8q1blhW8VUksv8joichTQtjhbE5hhNk2A3ilEHzDMjvSRzLm6MuNqjsY/jiILrQh
8NjoD6kOepSRBbvToD9FUp0RIv6P7IagKfAhbYKC3vb0b3WRijdpaLiBAT9VmFJY
G3v4pAJUqve/tgrqUca5Ts2X/Qtojq9lQjJdI3mvGfdB6ioAiWhKqHCpY7FQgIw8
HQMgM3GG4OVCSYyFqXHFjk6WEiidAzZGL5mQAKTCSeFkUCzVipgFC46+lMj3nX/s
uV9J+adgxpP2qh0ft9N+W6OHhStgb8oO43vb8lxpulfvrWzG7FKbZAPbntDY6LRT
KxmsEjU8zpJR/ZF3wi0twYXXNUuM9voh6HcwOr8zwW8=
`protect END_PROTECTED
