`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI15o89y291yBScdJl4vIloD4qRRlZ+/gpne4m+rj60+
QBFrgsUJLLXhPx/yjBMVS7m3VxU26Kn3wYjRxX8MjYcQMsY4GYoiCkCX77gBl3Ei
01jc4r9rusyPxxz387bNjb9+1SRY/HbyZqDJDw8Hl7aXiGHo6HB3LFNsgSLFUcRd
DZfNg1Ik/G1J0wIll35SaeNAU0jYh5oVgbydkTxRge9YS+bWgIJ/kQ/QFhei2cty
TElMvyK/MpBL/RRwMTW7GnAWVVeHAYiffL1a7K7HYCNFsWHhbo2yAGeKb7VtyRxg
qd7Kfyod9wZfHEThUde76nC4jTFvA0N+LS6Dpou0uBGRfDnV0lK0Yjb8zOKZHiV5
dt+2LfN8FXjSOTSrIiwfamT5AQ5mI3tlKk6l6heAITw2KUuu5BRBD3e5r/c2Bvki
vA5GZmMQdJRHml5L7HEA7ZBAqlzIBrLj9wmT5xdT6X7D2cDdE74nfR/sxnglTU3x
qM9VLkfVX8n27ZlZqrY/1oLESmx4rcEeJGFlZeMdSfR+2EwoEwYEfwnV8awH5jGl
`protect END_PROTECTED
