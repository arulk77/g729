`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aTzbBYleSnnq4aHszMf7erlWNtbt2kiY8lrkqsxorFUS
xVLfEddhWb1H6QQgD8WrEj/KgGDziAU/8TXs8ToIss6DcqxoE+zDvp4IyygVR9uG
xs3l6dZ0+EYKgy9VtInwIUQ/YAoHzppbkSjygsRtb81Ee+iEHriusXuVvUoOsbN5
m6MdFEyxsmEs6FGWe0bSfM8ADIG6JlZFqIol8XRWQ63bYqam0f+CEREFyun6br12
JFFX93TlKnveLvJJZtQs9kzUzaHxCQFOaYLUoGObKrI0pvukqiMFc6v+56Dw+wzg
vIi59Z85QXec8ptTA/mp4rsJcEZKr+aceEgOuDqSUIy+xt1FVM0DU+Ru4SVn6umJ
REsapnHsWuoXBL4bcI/YnsB7QEN8yDowRa3rw3UXDhPp58lL2dgTHbuwkfrdoE8S
t7K/K1Mpbw1mfoNIZMVg4GWQy+C3puE2tuUfGoRFv7qJMS+b1xncp2EZ+Rfjmsrk
WI5cONbz7SD92YxLRSq6/ZOGx+r7peadagfbE1Hk5ybEORfAbdpZ3/o08ey77CJu
9x6ffWzsnqlFtp4sypzOwCxLKYLx7onnEDsj6Vmv92p3Zl0dylNU04Y8dUX/COE7
X8ETsKkpUxtxrtS9lr5hzCf/hY3Fll1hi4YpWZWSvlAlEbFZsVIU3gBMswUMNmZ7
IPfIgbDT8HitkDFIa3g5M63zFHZ0GVMuWQo49S5wBw1l1CiPgiS2l4tnMftUZlSR
H9XnFlwdxvf8/fyw2Kn3o47Z1pBQ4r2nzeXPs95FMYDGfLvEUcllWu2zW9LdmHGa
XbG+0Fc8seW/woS3mCi2mLvoVaqH0M6nd06aNA0CpO/Aoa86Mz1y/8m2Cr25fZtT
DkpYg69IeZgOxaCIz3EH6aFi8kS1ZC7llH7WHVM2Prqz6ZMloVEP23aBNPW5GmGD
`protect END_PROTECTED
