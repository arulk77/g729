`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFBze0A5orb1KMfZzwYMCZUY5hErvElHIS4tnKBdYz2c
vVpd8OSeXRB4pIRllZE2tVgqGnTNO+ZwcqNpLUPdCsUFzd0PHSuXqLPWkMd3GUl1
dhbAvx4q2rFexajGY2+VGFdkz5Up/JUgPGHcZoyo/w7TcMuv7e+wsLw6NRzEMFtr
PRW5g86mdWOG+ulOgYtza5KGtbDOeXSulAQq+jocN7TT1GYPj167RXrvuTSA1UrN
o+19T1wYqyFhctrCG0TzhBzK5AU4zKPDfDOO6mbR/JFtMGxITcZldCqIjMweN9lp
dJOjoA/lLj+mX4pBsSEi6IE4s1EBMknJhWWbBUfWYxCRpIoozb1ELmZ/21uCGFY8
yxDTLvZmPGtWovFSLh7fg87ZudW+TY4FbfznFMbdEPhxZ1/u3VI1FguLYVmocb9p
vlVqSS09NQW3668F2maOQNmeW7SnprdyFktZ+8sZg2w7pc4YooHuulQl0QEwlb+d
SfbFSfT3kpXiC4kNROrBo7+WM69IzTSpPIeEye8oWmDlbkYfzWaZGbjC0EnZeUxm
Z3fy1J6g4KtQ/Ykcb3PRooqeS7auKzIz5KDuWPfFNv+zlxfvxecQtFv5OIyKmNvC
niqfvuXmkOAM9I6g6O6/XJOpogE5teXZkjl5CL8yLR72HBh/VtTByrfqJ/5GJBcW
`protect END_PROTECTED
