`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNwwoXeuGjgLIOv4SkvZ1nhKhITeLJ3V/8yWeNt+Iiwdk
h8AI7bacIDBOoOdVrU/XQNWteJeXujRpXGYmxshVZOErlRRIg0LyjGd/aaIjR20I
J84axzsSYmxR5JUi0xDtWH5mvaZvgGgZ8ijrHzdCLO3jQ+rWxLLBbUgPPc5YvqUO
aUv81wlRYkn5E1cbh5mytcecixhdeqj2cawborOGRVtHW7OElP4K6xFm/dBCxhD5
XnAdxLSIccC4GZBl7Oi+rUUxqu+XdXYgIns7vsR19BOpvstrii8+8worXdgH+kz/
b14Tt7RsTCU3a/ibbRMFyU9/8n0pBj4hiCs+Dy2lQMk0iEQeisgJaGg76pegz8xY
bIjdy2f/PSyNZq1h01/VDK50VcmXcCLJAMHTECJYWyrf4HpkZ/d+IMCBfLiv3vp2
dwbAfzeNe+1QwlGmqjhrV0zjFeDtN6SjekoRmxnnNaR65nZnBCruWiduPMqjlAqa
XHQqYn7GoUu8DYRDoEseIYBdI0br/yzeViI/WGEbSw3sGEWpBsq7cRlu4mGYGkBs
Er5Lz7I9DO3HNCUl6zRsyQ//i8Mbc7GVHJlptERfIyUohX4oTTXifni8XjJ9R0Un
MiVg1IyREgHap037BzzjPXIb7u3mCUPJCZW0g5F9CNmQmqPBnQzQbimxVpuDxsge
EYJJmYjSNYxXgqiYYZkv9BBt0MGAf05GjXjJRf2jHkex9QddbXdID6X7qZ9E6GAl
lfYHa67IWehvOoBMr5AYbVDdLpJ1FuHF7mLA7wXJk0/AxjYyWOHPUdY3lovIuODd
7K3iFfnmgrO0ueZLMrNvff7rm2FWzli58KOOMTann60FxuwWMhemENJN6XnGwxIf
s/AwiZTZidDta/T2M/kGH+0spGXduGe8X9o/mX6h0c1qiFlk/s/3OB/jhmoc2lpw
ewfsICAkisrJmkzz4Crb7Hv/ZivyKkKG5sdaVnJu8uMwhqp1+99g4sOT1rMZTQnM
UC/VheLFhiBqiJZObojbV6+TukYWr4C7oOUjFNNgpvj6IDlGxXkC8bVnHRTH3095
Lg5kD9nVrOuTHAuzt2NYjbosGm4zNHyxPBNQC/DizQZnsn6o4oM97UxCoKEhtfL/
KH5K23FYru/Sk6VW7FHDG26bUeHsQHKENW98Fw7k6liQ5y7arYhEMc9ORFJzwTie
u9fFiWqtDa3BbnP4m4V0tjep5CdpgmgmMnvizXElKnMM8k/Cp7EE2SgCJFVEet8l
GUXWOYxwce/HZS8KjlEUjkMsrYV5LsCZGIMnMXEOByRqcZVJVcOphdXRQBS1vb58
vmRlkgloItks71FPdYFS0See0eq1lExacmWj542HqWsF2loWO+0onm96EpWrdOXL
G4yymILf6gWCbVGS7url7Ue4qbl/CX1WJMyW1A2XcJWrjL3hQF0Xt2NDr5FYyzz7
SHUbxAltpjHUvpZStgglvKR1obPytLQ7Rwq3BkCbUo0A/UbET6eZPU6X43QOSwgH
bhIYjIAOCidgKbOXotsy5N0jXSz6QpkQOg4NUWlNHDhJy4vcs+KlQtq+JqcWeCFf
RVE4iIbHHUOzmrp1lNb0tMF9X0Bx4EabNy1pfy4Or6YSoZU2438GZ6sdN5JC1ufg
vMvK2q712yuGjmrD+fT5UxnoXbAJpQBxU1MOn9LR0a32KQOjjEDaJMpoGl46q20x
7gHcclbYvzzpCGhsb3Um5q8aZzfAWOwXUYWbZAZPgiM9lKI/lzBdBL+Fb2/GBBgd
SRJphzYdV1oR0xZMyU6CVtDN4z/+NRZbhLzymWpOyeXHNW2lLRXag4CVWw9NX7jk
Mdt3Mvnl72I3R4xgj1rIP8SH93sB0OfO2Cr/mGJRGnrIlQuqKogERXAaP8nHUzuf
+gzHOVhb+eJ3KxJ+Bh6/6vLEAhKTMPfNxEkeMT/14UiMMrLKWUVVrHNsrEcTcN9U
qM8wJiOKSM8662ZX4t0R16Td/qeB/jBzgwqSZwpc+F2NUb8KCAcW6W0+KnoTpqqE
mo4THQM0jec5nxD0CafsIwbpNE8QI3OdE6WPhklVyZJ4SYeH+2TEDgJPrBz5GX1h
1wNBhAQNj5evWcxJIHUOzo1J9Cle7zZQkKLSVL8CEWrFy2i4L73AO5PWGLxwahzc
YkuTQQjvcnSFCd5tjzmwiwldBDmwjiNT5VbU1spCENymtxqLb6FAGMYnwIDvacEr
Lr9P77PeJHtmvtfYQqPIyptxFcVl3bNQtOSHTzisUdk7rYMtwZWqcC43xv8D3aYP
yglvltOph4dHPp6X8c+cpZOvvUukRGLdwS5ObzOCU+2VsebTSLMRyYhAa33XOHWl
tfVT349KcY5JQPchYFk2+DFWwesZms1YkIFw9JHAbKe4Ywu4bdKILYVJWXnuTEmC
c4j9zj7xbBmNjNASlq8OlZ+nsRkgaElZHvy6yxvr+npKGtKLx/Wgb+PeSIKURrdW
myv54VUhxJdINAL0B8MnOoliASU44oSdF0HxcZuhjKsuulmUj/JMd2JEdF7ds142
CNSYxDIDVMU/L4s1OuKtLnj9majWvN19cPtm0R+RdcR+a/euDMuzsyArvzMGbT8P
Hl9FPGyFJKo+dbMRtbGHuLLUHpcTBI4IucqQ5yn3lb9vVZrcLKRQlvoO4aoa0ZNe
Prlyj7TDj6QNDn22p2QAnaufpRHKx52gaUN97NdhyxKYPYGQ+MZSSFjufQvpjPo2
Vh0xYDHedTBiN9y2N5o3o9IA7LIyO0H3KR4h3M3H8ia8I13gWUEyj4z00ShqGOT1
U6+ImfqzW6TIhRGwergejuDyFiMQnhwcj6uT+QiAUC+0/JlImmyoWgVIDo3m6XJJ
CijfYvuus270o3MNYvWJJTfc61pSTHf3pJPb1vCyGJs5AWTKY6URM81IMA1J9CBR
Wwvc+4x7b05YHjbaKwXliWcFoUCTZWPTLBZQt1aEOZRnTn2brVWyfvyTJZyhZY9o
rLtYsXxvL9aOqJrAUAzjV5tKv2S8B8UrsizEsVR8oo2uAcabPBrPxLBgDdqgp0be
YMn1j7qKoP0EWN7RO8t7dGQP5zZ76bHtmVP9uSDG1mbZMyBnnp4IF+0KjyxVd4su
OSmVqWqDiUwY79m+JCxmiLk+sicUY1uuRd9OQturw/97N7vm+dlSNl5xvMZ0KJCo
icIxWfT3tZZbJJK0/poEH9jz8DiSSsfJ7RfWRFd+ARnKUYehtEacgfDuQCCPJnA3
FT4Crtv4ioz/jPov7Jlc8NGJByiSmfpEO/sbz/KaYgEUM2FVXlkhy9FpguhnDaYQ
hR4FaraZCFO6vu1dqAMgPselQPByvJW/rjma+tQn/tImqRTpDRKpqftTCXqQLMMc
hQlQ/cM9wVqbrkI5N+HbAvF50OqCHfEUN1emBueMI2gPqot4VS66ySkIfewjrx2n
USyOCZzZa5yANT4K2BmOCOLc/7FlSvnbw1Qq09oe7IGhbXzqQsVmuF9jBkbD74z8
tIO3wSsAJYIGF4Wnj/VgyENfyVy3TPb7QFd/wrTsgfXTnvBq8859JyPcqNiXmH8S
naIWnLxU1X1yOwpmebkKNMi5NoqQ2sO+VHDu5RV95kCWwVJjxD/BU+VVNrNax3r0
jtIOVVgmxC2wbZp0PQQlvaHUECTwQZKu+6zgztvpoqsnrZHoscZJCy7h1n00oy7g
VIgvHBARA5QRB8sPWpr9RgEYdCqCaBXsoDpQbsQQKZxMotL3xNPY1zRMUyzQINsY
OCy52STDU3pKodI5+/0uGH7ShO5l1JbiE1mhLXtcVQgxU5WkBqwf55oFpvFIgm+C
7qiMkjueKU6By7EvGWHOsolrbHe1KOizsUsZ9ea8gnTRPlixMSTthEKIlhPIs6zr
is/75SdWPyRH+AhFjhKwBrCLsS1FN32AVQOEmJS40g0MCrsUR5w8DytPoKxsNdfr
+e1POrpS9jno2sZnXCglx0HP/4SydvaOPx9xLWrDsKE9Wj+3SwryPwTomWDQP24p
1h3MWALjLGd9PbdUP/aYNZfFj6nofrF1iAJ37wZygXqYEtBjzV4jrpw/m2cw7dnX
g/KgSZl/ktorh4Ng4mI+74u6x+nk2RfUdgrHtDSa3uLZy1E5X+sUw5JikFJx8OM/
f/B8vzWiNBLxYlXS3V2x/R11lj4KOpiWddzWgHTGBRL2+TyWIuFFJhrvWzSioK2l
OP8yrOrMJQ4ybieC/Ut53ToHhXaAtoZ+A6GHw1wGUzrmn3zbocMaaU9pU/YqBm+9
vQxgbVQKPTuYpdHol8Di039UJ96wcCovD6Elvbmm0Oie3rH8NTtUBKrkNUkW10te
B9pDZsp87rxI/Dc9BjDU5F3XRlwT/lbxaqrhqJmVJr3HDBma/UBJ7Dj4zTpUZiK0
Oi2rhaTaxAdpjZ6SI2ydrK9uIgU4aJRXSf8Pk4qc31AcemmB4n50GORmvzR5QSBK
nE1BKtO1PEXS9+mRXnpZevYwv7VUG75UNzJxGph6UGwiENusrZ1ja09LowozzhEG
3srBmCYeZZGBWO2acq/dBp8oTAzbLrZbLFqHVDmIgHd6h+nHTE8KDwJsNYjE6vur
kliQbXXoWodu5Qp3kR0qlzi6HZAuUR1R1aUKZ/fhDdaxGM2Uo0gKOBinoV9CZcSy
QMal761Ig8BaN48E7KNfI/wdzpN863BPQWjKMCpyuD4wAMz3/W6uU+XGVNzmpL4V
i9u+nnf2X3W7V3uWGoY53xq+fOpzsUuNoDbDK+31FDKoeKj//7j90V58k2NAM97K
DKQP7y+GfD/hXx5hpTyqvHHpyoFwfCylNonHC/DYesGZcoG8u5FO86LzUAPAaem/
MHTeEPxYhfYUQwEchRrcmCp3vmAfqW/PqjnlfcshZScFpMfXRBAFUx0Oc4cl4Smg
zfS2jJgJ+1GeHHHExZvMTH0yXxTfZ4lqLfLK3PFDQ1f6wajLjqtxYRcg2hQbbEMW
TM4NmL/fsDwyfM7Kgpn+D+jdVOhXNZXj94XvrgHJirHu0M2ATqc4eU5F8R+PUUK2
zA/SMMEeRZEVJdNAD+z/IUj6hZ0o1SGuK6fjz6m4xbaIG+KOyxZ4YBReXnfOB9Q1
tVJTzCV25uPTcB8OOTyukkKPmfTd9vXiYNUZ6C+1VZaelGGE2RoPFzjraOAF1VA+
3Df03vhLj4DRwc+ScXHFgq9LgiRHLdWHdjRD7HE10OCYAskNbLwHFLDXNmTUuiAc
tuauaupvXXA9+4L/yWykHefkCmX1lREh61aC9h0nScbVsPPsAcv2gtN66BFX1YuG
6IGiI4l1FscLs5by+qBsC4q1EISxpLRNwbjUS+cMazGX/SSAYIIAg77V0E6ngjZ4
LkQC985oqKyUqu0RW0kr7DzL5+OQfF7FwtdtlrTDiR5mhWXtQGYACpjPWG649N1K
wyJREjfJqoYQcC06BfmRlksQ3ROJ+CyIScZCcb2Vp3neCd2bYW0+aokM02EHRPNA
VRxHN+suPl9o92vT5bSRXo5BkFyG+Fiw2nYTKNN7ogMurRTv0k0GcZWJTdxS/v1R
qnRp7wNVo1LZN1fhiKvFj5eOIMfcq55uOx135bZcnL+z5HgwixE6cX8JdyiS7ct4
bQrpmr/F+NmoZLks9XfdeE+sT/aVNVjdbEtoPwSazOtBioJYIHVAsivu8sjqcWe0
20NmlsO2zmRlSUuyJQ6rBNPC9iTPgVpgTHK57sQIXDjkpATwQN6+q+C3laOeL6nc
/mZMD3SDQUTTFsT1JiJgRpCn4SRwfJvk52gbd+gaLppWH6EhSLwyiwMQ6LYfMo9r
9XdbsHyx/pc6jUm+JsPXoQOidF6NvpSI8jEySFrW3f28zvLnNb+IpfYEnKgrMs/6
sk/4J3fYxObH69rSTecia/rjZux0IeYktBe5uiHnXyAmuC2gRHSqMrEWJzdJeZf6
GYMAHbVcjyUiXwCY3q5mT0nMrYh+hj3qj5365ymIkoMlytgZLlHbNlqkQ1vXDLtm
51hKstJgVD9yhKLpsmhgGGMiRBb1v2mW+JGKo0sMrXlMO4/q8Mq6tEeY4Lh3BF+d
tg+1HcgZwZ3t3mnAAOuDvfn4MvYkUpubMFIs5UMz9g5E13CTh4EavshQF9CMnvmJ
KB9pCScqn1Bsp0tVLL4unLVZ42EbYENBc6oPJxcIkyQGNNxQQyyeh9pSDQAmd1eB
veyxTclF+vzEtn+07YI1cIsQjV6OJUf1AebH/RoEy7RCHo7+YkBpy3I0jPW4ipCV
V5Ii3PhOXBGmZfNsN8ePdwVmaYWGvb494wqX0tFO1437w4ozflMceuyaVoxYwH1p
90pYdD8CujMs6Feu6oARz3/3C5qfItZ5s0E2xjM9oVHTY7ArcM+wZQoVsfIIzU2D
TPg/3LkZC3ADhRnWX5V73qkFJRD/V9L/o0AgRRAygiy9pf17N+llOv1ZkP5EqtNz
zy0kYyPJpT142zmcKp10Hng7uQGv1DhYbH+QUzCte8hz8PoJs1XnYd2x7ipz/CMI
Okbp/Jdxn/hvVHu2FjypBsovQXGzOm8LMVVOt/8QMqJ6h8sFoqs39aJ1YS1z3GMl
F4ik02mXgSD2JQaESfuehoCGT9Gjp760kZxTQ8zrZu5gZ2+KfbFpdfIpbU1Pc8J3
J59q6YB10R/5k4438GarGHMkvJElbLYtwa5mjy9HItCl+tsVSsCuFUQe3O8/CZD0
nd2Yv7kfC+RORgtQr4iH+550QnJRqRdx9aUmZtef67+k37X87U1XeSb/TF9YbBNo
SbBaqi1PoghkPwlyYjf7/vzCgwkVV/cZLmh9xXn9TlcI59GhfbKGIH1mPGA+w59u
/PaWziN+FRStsJlwPLXdUJ6jeQeYjtEdrn2M8gDxtWnYC96P50DjuG/iWiXO0mFn
kXVYbXj/o3cbZOJvyiUU8L9J1GBxpbYnvOJszEwyhA0wqUSSlR9u5+b+/hzDIzVn
sZOjtCjjVI+gjJ46w9zTaJ8+8/JD8ZhnzUemQU87tBPvU8OdssQVrmGkqRq43yRy
Po417n7HtcxO8KQkLWwW7XMl1VEgRVQrTgrMhlMr+OMlBhyF/SfIDMAVcqbdwZ+t
uXbxdaJ5ZT3aF/fEcQhyYEZE+SLobGhriQKoMLI8wUFumPOaLLuz2NcR4hJblFXG
AOKZUvMnpVutIgggbfwpWmv+woI5G9dgsi8RvcFp1ZzfnK/y9AFEuAE12/hpVRAV
jvmXVpeMKHSkMDxAyW6QY7g/JHyQtutCTDPDNLvWMbCBxHNXHNmC/vwKRn/Dxnwd
D4DFmHLEz9t0Lkg2ZBt9xcGG9zRQhghhLULhk/hSm4jMTiF3BrCqvk+7iV6tAfq7
zOfA6d1ZB+WY6TN91AFCVCk9thaLUTro2RcNaQhQPQyHJ2eGzx1L9hCH+mcK/Dud
U4ueyP0EfpjKU0o18hhEEV+v62UXVhWMsr10+ngt8R3K6wYL+sFIwIX0+KiWBYbT
r/+MdFB6zQ2CLunuKo5Bqh79cVzbCn3ZdyZRPf6SVWVh1XY+nJAVkmoHyXv19+Zz
mwp61EAAzgofVcOqEmgWB5a997UUut+dVSjgRgB5dqqlFOsn3U7tZwCoPitw7PEi
8zrdSjvaze23kZIUEsDzrTpq8uxd0o2C+YwY4WOwWSDLyof9ypxEqNJBGh7NFGyV
h/wegYZDuWwYh1zn4yJmd1PW0niz6Txn4G8A5PhCr2fY9TyDqszI2JC94GcWHNrh
QSA2CCEqL+qmRB1b/RzYVgCwpLXrmBaQU5Y0k1jdMhJJMZa8lIYgntF0EIHfVVfL
D6/cbeXNpLDzR3iqXRPdoMZOBlHTIucNI0fjSvXDg8EhyHwu5oBw2XqpZzbqU17k
tmNoMsANjJqV60rbmrvX+A7jqxt5ea+bkgaaXaqjxpuJQoTETaWr9DamOdq8y22y
HYeh4mWRwBxxcYTpypb61nGfoK1sPM0NmI7GM0ysK/nEmUBE5e6MnWz2YjsO88bu
UxPtqluG5HzIosgMkfRPj3oLMiZp6zw+bfpJmpCdp1qtPfBdPZ7FheTcaiTaJnEI
z/4Q6EtfQhOGY73XCHgHeW25kTWqlaxI4MsjQeKLWjw54kRi7LuniOqmpuXmZj3a
U/d/psTTGUQkJ1Btd8OMXKdsj8V6coTA3SmTHje6MwbMqjE6ILBIUdt2zKOPSK/m
NxBYfNTmxLBHxqVjBLf++fMyk8+VllCGrAOx/9DqRrOwxWH2nckwfU+GU8T84x+1
yTm7yFBLwZphgSK0MipWF8oIUpOnxPfCYMl+UCeEVRckIFynI4R2HFU0mI9JSpNg
6afLcZfurPXqWJ7neDvH8UHczzAUtCwQ302hYUjT+udI1CGTQKX5wcJAUvEh6xkN
mxQ3ML3MB9f3DaA33ewFI51pKD9HAP6eDGCu7XDOyi7vTYjoXxh1FHZWyRWH/Siz
w+Xv5fwtX7KPcfCOL01eaWMwDujlofPtEAqZNqCNRewL+/ga87RK3+crL5f7ZH5B
26qYG+tv3dX627jIDkooaD15cddrJ/XQV0AMHDTeNT4j1GOB6ZcTsbCjRG19gBGQ
ErTKnsKmYsnn6G81rWKylHbFCn5h+d5h0jT3ExscHw459Q1DmqZrruB4OJP9SzWP
jZdKYdQ9PP2pDdwHZ/5sV4DL+hlPXcq4EUZ6thK+qGOsnbSE5GbedEar7yd89h8Y
YMEsrGh13PMuuidhq3tfUkkAgXIJkXcJwFZGB0leePsOKTgq/Fd4X6XuAcuJW8n3
sSNMGpNWDMIoeKH/v8Byjhin4Wo92Qu93PdDXrD5Hkp47G4MoQDm1MTPPHLypTcE
oN4J2LbA0gNtDVa1n0dtzSKnuy8Q7zr7pM3mc/2pg5dNI3OsrtEoAUk0YbYIUeoC
rjtTiVei/lohM6Y720B2cHLC4zjIXXhzjM9l3dG2MBjcwBZwAX+FpJx6DI+xKggQ
peeZ5lExQYuctyqrvoP2i1onquan7itKOdU0PunJ7UD2W2CANcuLfor82Dnh1g6e
r2LLZDs3WrmIlN+A+HD9VHYO6TGcselwGSvB30FDOVmFP3Aik5uUufFSJSkGXFxV
PjCWx3zvqzJq680nDoSoyK1OYPfDvV1Cz9+n2b4DtKwpREUoTxeiAqJtAb43oZI7
3BrQl1CfrhuKgngFJg1f5yHcUs10Mt2Ue61OybsBHjwRW4Uenrzm32R4lrtoUs+u
1iDLSnVZpf9R4MNph8WGUw6FGJgMRaCJwOzDp1jpM9tjgT3F28rF+GS3/HapCTCJ
rEBFnptsagBYVUkH0WNVLszSs+iHeyporuK8LM7z5h7Cuz7XK18MSRwoCO/ehbrZ
22Vf0KncrJgc/iKu3kd8BRNmV9MFGu3nnX2Lfu/6P15B664CmINnFcggFSWHmCMG
Ymqto8xiWgYjE5J8ESDC2/puDjeJA7r01Q5tvY4ArvKAUAu95+HOHt8qTEdD0V80
5DuRxGZTHyclmAc64/Py2rtxORSNGjeL4jQmaSo2xtCW0t/Z7JD8Uh7Ic2mVoGgs
/3Ab2XAT5e4ZEZSW1qM7qU6bBydp/jp65gMaFPNCQFjFscV9gqDx1GYjq2Ei10Lk
dizXI+meGRw5NJqe2DzXGEcEUkkWko9bXlJIqZ01TN2cugMpcfQQN866M8oPff0o
wooJruATCrAacCbtdQE2R2ZZ+SPg78oV7TVUCQUdM2P0IKitcD6HSIrIO7vQnn1l
lGAsJx5NUmVPuwWUZALrBjwW6OEl4lERZcFL0ksR8whMk8xC5Rzlyu1JPaL7TpM8
jMcBjm4z0WYUCMvGfxerGG5N48mfQ5J96KHDf0FOmI3QMstB9BwGRcbJQ0oga1VL
W4Xjf2WwghWs0SDVTXWJcpiv3bUU+mfz2fCMa6PrHp2UmGBlquzt/qRaomOFKN1E
kjTdB21ljMOAKo2TZspv/zCRj1t31ttxTU+u00OKwlWrqakqIPl2hcXobjROOPEm
wbUQJn6sTPwrPt1C2LLgY8tTEGJiejjjlppm3ySeentNy8iaRcfJSEfAJRwgoZ22
jmBbioJQfgagq8yQ7V4aN6anmjhBmMvkgRIRMhedI6KCv3W3+jq+ZOYYaGHRpYUj
2cpzLj3iM59l/xk3zkr1EdlE5mnISOY3CAuwlL6uREgcCQvpA+xy51fIwbCVUTVD
4VJ30LMcP9jkdW1ZMGDa1LH7LKLEkBo4Em+BnWKS8SgennHGH+3eU77CgSma/R/a
Vr0mY9ULdLmsUQcr8OXEP9YvmSBOs0Z0Gm7wYezQqTHLYtrhcAY7prp2aYouqvYC
683oprt0Bn7X2Vilqpx/NYCRK/Kh2iOkAjpq+jBO/JZJBWeFBAyje04pNSQK4CgS
iE1ud6/wDwxf+Za2f6LzUW3p+WKdngmSvtM7cgjHdc3/MRTW9LRxl9gPkUu1TjzS
008879fWgmFdb2c9drECBPtATvGixY8mOR+XtARvwPtLY8O7CdbfnFjCVOpv5XK4
CnV5KvEHx0odufn8DfryU97e4KzhBHaAae7AciLuzSxJ96iE9TI3mfNFfRRpE/KV
nAcFQVmQMm+16OyKVVd83d6nrOSCi2cBDDoGOksSkP1YavF0bFVjWne8dyRRDqMG
hb5aWGKzSLyJBIXR6J1ROInOPVPTi3f7P6i/u9EVT8jSrIgEyG2GmXACeXnJ3MdA
rq1vUsPaZVe9TeoExGapw/t6GzUzRzp180u0YB/q9Yydruj/ifzXSDMq1RtIDC/y
OCgWznOMb065krL/ECIqbUa0tBuT5BZSM13ryo9NhsP9wzmICP2kRC9Ph2k2TASh
zKEww1k7xWytdsYj081tQ+Ay1RXUePCzLW52QnwNaGTHTAW7EYFG8dp0Q59Vff2n
enGnjRCSCENRdbram2SoAE86P3hZRZ8lc/pxeRVzc6oBUnIKGhdnIO9uAEnzamKw
Uuav+oafOCom1DB1KpbY6il4wLhI0G8uuAWJAHXj5vjyB5hAYfkYP/CRi3RuM6aU
nOudd/HMUfH43UA9TASFokSF87lmiJ5Pu4Qwkrowdaf3GrXci1i7PEAH/b742Zfm
EBf7hTeDaXxs9jkePQ6V0/fD4xEUKvCOM3ybV2IKXfaCB+c5wA/LEn3i8CKTsYSC
bbkXb/fDtlDLQl517pXMomUyQ4xv9yCAd9T+3CbxZwuBBLxAy5MBH9uatJb9SCUo
B9nbfBffoUQR9DUhJ38eMUJRx5sbeEU7LawI0DvXEpEWFHaHlTuBw9KNrZSfWfHi
VUwy2PC7Jp51Qkb4foe1hWWWomVB8EGeje0+BqR8+c2rTHmcq9RvVHIi2a91tute
x7H73UUHVl2hu676a36P6eeDvfrRNXT6kabdezS5bp2Ag1q2dzsYXY9IDAvpZjuK
O3CugxmXly7kcIOkAQbvCk20mgEAfqoCxE2dFnw+ZoDPPn7+N13XZjZ/rgfadoAr
7WnFQTPvgrpBMHXGQl1aPSfL0/3RaLWGVVa3esQvpNM6OiJCibADZ11KtVm6DSgf
G5HxIcgB7a2QykU6bwA2xtkRUct1vIm7029JBL/4lCXXXH6eRJ55lFsP1zgG2reG
w/e10a62DkmPPumszqUDGEAjjP7DxBt9TO5BYtaq9k2HaIXiCJGtpIXyVSupe1k1
xl+3ZvBFx93wSMOyJ7hyzXUbF+RfYFJsVt6ROyhQCKB5Sja2KY77dtuOD7d4cLQk
fyokNBbNT1gHWxqulZZO21IbolRcjhYT0YhGHNu3TcH/3JNLsLmldTQm3/4o5mbO
HZcR3vh+mBsn8+E0XEVTm+TXRtkQ3eiRHiyf3B9JyBeeXPS+S1h6N39h2ow+2aNQ
xZ3d9BjcG4TtKOYw/6joZTtdLt7NENaAb1MxYAGJ0SefQ+ILs0UNDHmVWNGT7PVv
mO6IB33JdzCjaBMRnnyV2ei4vpeN8MHE9lr8yczsTfhCk5X16cD80iCvK5fmvF5/
oXgdtlYeXjtYwoECPjWyBFyDQlnmYQIf+3NhiytZ4H3emIY5/35FcWgRy1KFVXF9
qrk9Zx3u0v4nX6FGPbhV6SxddoWXaqhMegq5Bp1aMeBbBNE1DfPhBywqizqOi5iO
4KD7EcptgdurfA4v3SJmFHBEgaQf6bhlEftuzKxDj3RYrf9E2qlWAXf6ccQ7JM2N
F1tGZVCp6FpAnvyQ7exK1LE+B00qr95JbYlRwenSiGtvmNIqaIUDgUc4D/G9y1RT
IL11W5HsgmqEP+WJAXjqIW/q8En/U5zdV2tIuT7Et/VBFehCw4Gf+OdFH43E7Jdv
rAe2n5ZsAJNcXkVEPMtVF6PLxZw0S+/1fqZw2frOaJmgZspA3OgikdMMeF8OYb5X
ivUv/uhlrJM/e6Iao9IwSJgCOd4QLmQll6UG1MzN5F5b4JtUIq2xOQjIuRawb8DI
SZbOhj2uM8W+KBtnUB2lpd4hoN9PLJOM6LcYwsV5LXlLDhL0KlEZXR5FaaDEeEQS
JRw/V2kMfJRR5M/7iBf2Vh/1te8cHXL1Qg0m+BcKI8Gmrdsf+4/gw2yxFN0j8mfv
C2kSNvAA/y5gSBMteX0sZHHyjpgQ8tQ22XpJ0ovJwNYNIJe4UMbXK6RDxu2bYoBw
cufj8KcxStOXoAvU7AoDURtaJKujHHUOlynSuTT3lkPQN4C/bWQ7MwdSkFn3NF4A
F4Km8y9MAOazq1nPq9Iah0trRIJ6MMgSTFh60j2l9Hg+tlx0Mg6g3/J+Hre1AJHe
fNyAPMGRz5+t3Lay4AZ0iibml9uhlHtFomka5o0veuYH1T26cwX6hnN/BxWQ+RtN
WxHELcnrUGsNeXSoKcN961nOyGjtc7LJcIqP7t1cGQhimKmqXKCNbv7DoG0EDO55
yB2VLV9SWzgGE4AOCCi/cwdvfkX/sfhxSoiWbGsrDrmEsI5pCnxgY6cVetzz5jb7
2soRYalevvMQiy1mJjvEJ5MW3NnwPAS1mvnTnOF+kV69pJBJjUVgWSigMebHiwuT
LOu8ApO2tN2qgCSrnqsh9dtejTuUM9j2D9lrrF+i2NkBxXYXEmvZW2pnWuL4ZfIe
MDdME6vf1UiHdpB/TfG9qZx05lJy23UPNFlm9LQcA+yN/Fw3/MPqbw4CbZ9NsisF
MfxmSfUNqQu6J9CEHasXORSJYYm8uLqtNBdXzhZct3dMTZUq90AQY9L9KuwFByw6
OVtnsEly90PC5b1xBMmx4DVXVia1tLG/wHZoC5cqNmGETjlI2Hb4YCrru2wTVZvL
wwJAt3yNZBOw+HqDseaNFeCaX2yN1muUHt8EAptW6hXmkj5sNPcsI1RfsvgfGs27
8SgekogQWkxiXinVEzD75Wq55Yo8yPqgtJe9+CYbHiURNVmMRj709J8s/AEdbqm6
Tjxr7cifS/SEEl3xUzujlifruGNRRE/gyw7NQWK5VwwE/xcdhyX1eNIdCff8eT5X
BzPEFDEFyS3wnniHPvrQs9D6VnIGa8S4lqk/rgSQJ9GqI2H3KtdejaHCUCVxDbum
il9/vR1shc9wQgxlSXpYhCEjyQWvW11pXhn0sSdnFTe+RAQ4tRJzO3Tj8BZCEfC5
4L3PTMTmvEXdr4DBcVfFMEzIKZkUod+LFKg05INaOXHS1P2Im7A3ah+9BxnjOHTy
GtkrYi3YPGOvNO/WJURnKJcJLJw5aVNcaZzer/g4G0nQq2XLFrSg/v1j5taiMerb
2Reuolr6AjU7pB3HvH4JiDoWaeKsQ4Q9cWNKTZLTQA/y2cHHP9C870V0TAKqrviD
Hue7ANkbVXQLNgWGYdNr/k8WOd+RBP9OnjObNfTyDzm+1rQ0gmcOsAnDMdxxpR7W
Oh8VysSyMWyPQdaHWIzazQmPlssB4LKBJfeRKuLAZxopbNsNYun+/qPfhwovA157
c5RBIP4vWc0RG9T8dHrWI9Vumyl+NqFaPATxegEaYrGvQOwAsi4F6UARWGLy8hq3
dkKU/VVwRfdPsou+yMXU0kfpnotXKULJPNQyzJdIrA+lVRk/xcDjGDJbApqjuoy4
bHz0tT7u6DCcEzQR9heAbPWiLF8bfo/JNQKTMmf5gJivx4Ps12mzKF8p+hn+y0Fy
kmMTUAOnfms7p65KOoYsNv4B2dPDYSQSQN5c5VvnXKLGvAn/Eoyh99Hdpdi03wtI
CFOr5ViKV1LNnldLy3vSYDmtFqJRktUdFYMmyiTwweuoqAIhRiMikX/k4Pfio2Xw
gUOnfidUVx2apMSWYOyEIkhCf9EZKfRhHc9QhelBnPZOT9QHa6VO+J+9rB16LrXu
n2hlqJ7XVb7FDT4TbjnGy6L+5I6wlo2dgxoYx0yI6jf4HF6XLm0+wSWhF8qr4T21
FtD2BP47FmSDQTz05Xv34SZDE2Ect52sAlkfuk1TKnHyQqHjm8LTJB6n9YsJnrT+
qNCMpQQz6tHYs0uAhefgQIDW8fHfZQeh1KRt31ouUn9pYiPhwfXK83+HgxTFhERZ
S5bU+4JSekX7ooSlZ+zLvitgxQ4d1yVwZolWJI0PCv/muUpHACVMSO4DF1EUTaBi
hCFtyHdQW1NPGHMs88zTrIpkx56zRp/ywPRifuqp/8R9w14lCOEzr/r1Lb9mhC8f
62yprFkLX/rLXWZDDFhjE5qOM6EgGQWINar4ZxCQCMGmsdU/QGQqrOJly32P4hVv
iTgX9V3d7rEYVsxjXfW1Dh6yrYs6LhyycZ4J3qdK0f1uJY1REMin7s5CIFUw30Ip
RJbF1vKXnaO/BCjCr/p0AwLqE0ln64ulAKVLBMZtWzDNt59BMYc0ugZKTIhIfP5B
N2IoW6z9BvQ11SLTtlYhiAQTn80DqpvAr8gTSBFknSukfepT9vU4MohguTk0t+45
tzoZ5UocA3KjD5FC3AJZqonesNJc7sG5mT9eVwZQjXPq1dpYb9UW1KApdMAyLYXt
IWnatP2JlfB48arc2qSHzVjvS2qzwO8UEv3bAKlxaduBe4jp0256lG5ALxS+mLNa
x6g4tdpBEVZoBnG460RF+74f35aL705tjkh2iYEsKpa36X95njULEpKGzvGCmPm2
b+xDtsFs0WV3WAZ2oX8JoSV+a5jTBayU7ouXKSExH4fA6R8/CIkKZVFqessqxb0C
Sugxvv3qtFTO2hWLtxD5mHoygProCkx9+6Q6VTSoX9tRiu7QTJeKj9KBaYLL4uSL
K5zQ85vWAOSzJJZlXmmxAw3A3jHmPQ5YHL0wXZhpI0D/bl9I/dMHQsTe0KKmS92k
/bz7iOglBchYxHiGzg8xGLMj9KeBqk4haqkKx3yyGSgPcNHGXVgnoytiBRSFq4zM
kWhv3ffW74F2/Hg5nZ48IqBI2jbOagnbN78RT+X8If7er/Thfx4Aus9r1PQgT5eN
OfGFKPD5krJf14yirMIRGU6tE910aS5CqR7gjljfj/QGETdp/yyKkVB8O1u/zwmF
89EBdCJ74bX8hRN+lS+r/Mn22E1q2kTAw8DS4dRybQGVf/XNHCxo3gfCN+cNsA5V
/Sg8Ng4dFk/BT0TsAlo4JYooIoQdWLO3UFSrQi8NFY/GyWhDXAD7MbMe82amf0TW
yhFAPSoE4htVkl3gR/yju3inMhwvavPmeO7M2k9oXRDEbk+JVR5AzHURRzUwv5OJ
WNemPQuTLWZojL5AeO6rRnSPJ3YxXCjtgiFOGoLVbTC/+5hCqgOo/wY3oydPUNU8
gM2a7MtyzOSswB6SHCr5QFhmnmvcJ37JncFGhum6g8JuehpnA/skCRgpc+p5/8ua
ugkJ6QjIt3lUzDXMx+rOqc84NmFqzYG+RXUfW4hNEHyXunh/MQ0vG0n4zKkGDx3k
bLWvsOv5hLs91lEa5ZmiACco3NM4c1ZS1tW2B7qtsJyqYmsMDMJmZtp2Y8ImVkiE
WwO4+4pZ6WmVkwIUQpetft895Gmal/0ROOmBZdLZNFzPjnwcVMuePoC/7a4qZ179
4dkfRcqdMiw1s0uuwLD3XoxYuBCWGLwtf+A+fEbrDeULJcgLhYNPmkmJnDMssN8g
GntiWfuyV0e69bkmUzPi6P4h1K91uBMaLCC7xXZ/9dHu1DJdIuobt/a6rrLXvvja
TobYErOo1qsw/MgaPQkBxMyqiE2gH0sAR61KmuZkM2vrivmlbf1RhVhCpoBPKhAA
DhiyO5+rdeUYDGLGX4oh7nB1J9WHOZBPIu0i6ptFobjHDHh7cS3r080sAQuJpbXQ
SFTi34jjpN19fDMmyFPOJqKkZXg/6V2berf5W5fp0FQb295dUWFJe8IJYVCEsTC+
pqS7loaZHKLnCHRmNa7LqJpF7FgTb0pM378Y7jF82WMKhVDEQFb6JYqjnnmi89s9
w1C75+Bs3iCQhC14RnIQNUT3dz6/VA6rpaejKVEoq2sycxbQH9EMoKYZ5x2dooKi
nqKHXn0ahxIEmhBFy0BRMNJrJ+q5h3kt5McvowcBtpZ5NrGMpzz0pmFMNL2yt+G0
c0lZNU9Mchx/E+L92Vdt6QXaovtmBfZihEchQoMd2uZbAo/tLYCTXZJYbBDoZPUG
v4l/t2apusZFRiwjykyjRZ1Qms9r4z1h+GpKbwxINm2X5g9zXn71uTE/2ueYiLdb
7luM/BbfwfSy8IS3U13PUI7GOKMfJbnYO6HwYO/G87IUKx8MmWfu+MIR364bSBaw
tEyLagtapzoGGT6Gq7SgA1NEfPFHcAObJupOeXNmFgc3LaDGaxpl1dsC3OKt6Tdb
D8g4XKtyIx6xpHx+8uPpdE0cMY6NKiPHjVggH7f+FSVjyPawU2vFoqwiabe8pV/z
84aXcAjK8sh6x4KX5/wF0yNCdyBhaogebSaLqY8JEZfzVLj4lAfuHdkAmaNBwuS7
v9Ccxcd1QjnogziOdh6CHAxtmlYTXUuW70ksmTT2REJYHB/3x/iIXcHxwnAqTSKA
e9w7gausOMMQoiIOwI3OWSR3q/HOn5drJmbJ6KirD67M/+Nbo5r3CeC1G9ppOxQl
GHDlopU6D3J+MXEHL36CgKuxVVkjqH9HqRYNNd/L0RrAOrbS2Shat8xg3Y21lH+t
aAqkKnAqP4eSBn5pSPECYu0exQmk31W7Mm5UHSYd+hbq2oAh0DAoIh7MlL5y3Zh1
80NI2GHI1nvaJNT5z7G4DnpXWzWs7f/YohNmUAd33xmvn9dtqziFSm1toRwLppL3
0gjnSSs3rwJ4+GRAD/dp+TmXo17PwN6g0I8Q4JAuQo+oOG9fzLf49gVqg7uPv6UR
MOWy/JHPICU8QS1tK0dlpJjJTcjTJwoMC4AEyle1Bq2hqa87U90WGGvWtB8j+GML
pYW+SEz0IJb9A/JZEZOcl3SqsZ4yjDfs2J9DlaUVu1YzknEdnyyWaHgGfwyTIwaj
p2P9qfG7IxzowsEBeZPtRuqOjyCgF715Onry6X9sh9/FOZldpmHclKAmNnsAucU1
YGNrENJsZHAjOrOh6iJ+1PmAWHvWJESW+IzBYLeTMCvTQjhu95CQwbbBH7NOVtjW
oqDoH0UVjyXUlYfsveoa+WSHaA3FQ8o9pQHnyfjI4x28wbIITmB7XUCov/mi9bf2
CT6ARqAzQIDyrgpTqrgsXO1FObgpmUY0eIUM3xFfpc0BGkJ9ElaK0ncaAb8FWdGX
NsVVPg+7YnoUrSyRfdgTe5OfqQYndGddDDked88Rn9d3eRcamXH7UdFFOuWOpL1C
zxgmQyQSb/Uf0zGyoN+VyY+8JGJtMoTLhf4lj+fQfWfooWoi4DtGyYynRIPy+4tr
Mi7tdo4cdh1GotC26sWPTACh7VmJ1KNi06SCUNQgh8qk8+hChY1yN+MtiSMO/7Dv
xG8SSXAURKTQobdjWPZF815hAqOotcWJ+oEPzZt6+cFV5skQl0A61DgHZYCZq9ym
2IFBB3/mG5Hl9SHmWQ0PIee118ILpzJNjRPx1jwZHU6N6Bfg4d8juIdDi+iLWp12
lBffeisVQJJCbUc9Du7i9PM75VmgXUCyJqmQob1QUTXAT0vCArOVyHmrWnhlSLtT
ohNqhcgmghTwayez2BbnA5mzOeNpAhnhZuK7MDfti75yTM0UjUOvRz6X76UeQio9
1zbSviz4ayCCogQLt/edg2UwalWKb16e5xx5T1YZeg89vKn0kcdvy9ggM2Oeg9ct
aRrGNPWGUg+nsTiueYmQ5BiERoqiO3E47JGsklU5I5JWI43WSZFqYmQ/NEYe7HfZ
JVUFhSd0xhNYtIlXjg7k7GuWDKhV+43E/Mp2aFgAbluHnpsHSbQEmLc6GergtBpw
q4C9J2ZUahdVtzvpDemoqO5dUge6cACJAbC12i7AuCdjAld5OCeKFybFIJmxpWgr
mYJSraSKMeUaCCeuacImi++JIZHpaFD/tWlP1ctGcY4Ypfw43miV4IjvdPyxnjce
xhio5gPU3cEnEnz+ZC8yoiTyVcvBJB8VNaKiasHVMDSjMeGBb/0CQ4cUZ0824u5S
kD+EAkP5gZvrHbreTn8W3AA6T4QCjKOA9X/INJ1zgeCwafpxnPdr6EG8WQf+/24Z
HbLYKWMvIUYq2lPyBqxuGnpwIZEuEYx57K0p1hH8l7XIM5xQaIKrmTbqv5p+suGS
tTntRkUqoL30gqZw9rf6XrsI0OGYaOYid7+sefgyCRlFy+x8Fi1+HZ0WDV4/OGDK
wH6oIEsNHHkYuK2gtpUH98N279QhuW030DQ9Ux8JF+GC7eyA+/BKOfSBvCBiNOlP
olDGVGJph7zdOOHlk/QShCO3+VdH7LIz3fEzGYcopD5UrxzPGl9F1gtFZmdho6yt
i5xoBkZ210Wxm3/WChIXZ/3kQL8dQ7NuSEZPa+AOwa98BaDqjQsbk9S4ASQBF+Vc
lZ9sIKiCkQnkd/2qlOtdwUdJIUOBijkhtXAX1h8XKVHsjiebNbWFfhWt4IgnT6BY
6VlctD9xuMjEQjfXtNthJ7X+IPg+mLSMrjKiV+Gm/JcE5Af9fgz+sB97H4VjO8Xd
S362h0jbhAUGEuxOqR6/bkWY4ZqKHkoGw2FMMvX8FSaRcv7i/KVTHf6TIIC8McJH
wqREAoTDXCH1FNpZ7PO/8e9AOeMH9xZ/m3qlZ/Mn94NaNalcGtkI+rQHIpHX0K5x
W0P1DEj0FZ/IeA95XWnBrowr0ORCCq32YlveS2kvAMmkxMmB6Kik5+PTiqhupv7C
1KTYsaLmq2J7fF7lPFOwNXKP/SzzZyEDfUuaPnkfC8KrsMeFEhWST0yY9+reuvqG
V+a+gfKDOB8TCG8/jijOtKZnZPESOZf6yQpbOoprCb5VYeHoTB10W1rpDt75XUHU
MxeQAfzIClRxw5UrwUNBaA+sL15BtAEV3XSqK1Nxp6ZXiN+eOb+gg7+Pn1XBDM9V
YZWU6cxhDEQ6R5Sj6GQKcBA/l6o/mxF3ztEyXI4oqmyJLZm40Oh0wZjlaGlaJsO5
F1R9Zhvp1ywAAIHR6oIuL2HsMNmdDxQRit5rYPO7sSX1KlxAhMOkIDnN6SO4KFV0
LrXQxh6iCeNzmeQIZC8P9yX3hSE2oB5etrGo2Qouv+0Cze7P9eh45VMlFmgv8wIx
PNcR5B4wTjeacuVgpY1KxdoEmfE+EqcwvDntcdmsam6/Xn52etoJskbl3jCBslIi
aYUpB/eb9DCKDvKbsvC27nMBmcxDoLXC3DFnhA9z+/e6LosLNaW8npVqwVK3U0fH
FLYSiYmyMmniyOumDwcAFJAM9qZ4WwKonuGhLpDM2lv813HGxTFJgXZr2ex46Jy+
9da8ZJO33oYozRWPhvjMfDGSIQoeFz9bbiL2+qy8D+J0RbABjo7GnuYUbs2G58ij
wj9Wue4kV2Z2HW1wpHlrRHg/lbpMKthdLHgAYPSrzTB1DCBs6p53ivWPWZ4wg6ee
lUxspiB/lAaqMywpTRnaXxEe/p+RByWrqOvqUqlgoIL3D8w+ynNT3W4b1sL4Dnlo
bvuVEILlo4e1Oerpd+SUCtkyufgG6mYH/Y1GcHeaMSJE+Wuzm0fTP7fLgyrYFbwq
/XhGIoTWfamb4XXsMDMcN3Mw77TmnclP45Na8Ar6/WEtI23Qe8fujP0KP/23YKPS
L5z9pZzKcB/BAYLrghsd1/b+QRgGS2Xmo1DLxzXtv0EKX21H/d+QVPqE05CSa9A1
11U2ppxEKB7lipPo4Gdz9gTnCZfNLNDkgNKvAMM8d2Rsg9Mn0q67Q8v49whOrC6R
aO0u5NLgOmzz/EV0TVwPiCwphxklrb5HE4DphePcHxaBooTerqMLAFxB9dIx0gcc
arPyhPLDXnQxf2pmsKKqVqeRt4q/pSGf+fpV8IGtdDPGR/xW8tOU8XOutDH93zbJ
Zmd6zGntMt9QKqjDO5PP0io5mDBjaOPqVx0CGsOg/UTMq+rNYam53DQNAL13LmG6
pADJWuh6JPiaCbVbVbE6pKJ/2f9pc71LbPQ2F0ljnUF0D8bxuPAgHIe3Ec62h1cr
1pSmmsTZrLTTNDT3YpUvgArR5R5yDjxuQ75xDP0zPHe6sBjKxYxCw3oSiIrdkmSi
8gmOvejGf8yi4dmS11HEB9Xq05F+8hD7mvIYCyaRB5TEFjoSPlrWOpYXvbZpN74f
6O5dWi5cvSeV0HoCmup41fjNYlGSR3rZ6yYxayZlBKT4bAeJu8OhU0SjOVPmpCHH
Wd4mWziuP2MJV5tBF6RhdTC13UprMb08Slak/q0zOKLiPeajjMc+fljF23mZSlrD
jX3f7WUg9wVDlGMFTD1xzURUzJZqfrA8eOR4RuGt1C0hNhQs0gs3e588uR3aIwnt
pdz+1UMUulmiX1WHOJHsSB3rhlUh4aMBhnxpI5XHa6XXHpI8ef1myrzMWo2QLRKa
HpGN3/xpop5gYKEn3mO35EssDoVNcyrjQoIUL06sgP4nCQJ1VUsTbC+d67zE+PjI
08NMqej0/+aXFzEOjkaY19YrTk0Qv9Z/uvGGxhsdINxO7R6xU/UC0eF7Q/HP5VhU
yXe8DX3re5x2FlSuSRaha/bgj//YlZ7eG+etqquOsOZoLvxml7wiSn3ObwPt+M6y
DjFnVPc1dmV4SG4mR+NT5TDmJZa8rtIocTCpgg6MCmkF9oiBTHqb144NhRxywT3q
STC/IbKk2Roca9Iy9e7JIBfUMM8Pbzuq5f8bQ4CEzGJIhTBd0+1LlP4Oe+5rKzO9
FtrE/IxB+tlGkLzM9yV8/gv26qaAq8Ru7YZY3Gf5tBBAfy1roceUqTEW3Bo9StfQ
CAujcDol96UAcRvIie3jFAx2CjFwQnIki/LwSl2o8M3SSxua3Jjc8ZJTTtZj8pZy
yCEKBjlveaznBcHw3q2XyatGJorY+mySo1YCGjuwLumZKr1LmCn5s4BSx0m1wClp
uuKU74VlAZdibbXusCZGvYeLgmKSZGFpkUF55enI9ACw54Cl9EBSGP2qGqsjSn0W
MnrymbnCTI8+BIq0AQLE8txRQ+hoqvn3vQvEjNW11DmEniVb01UaXR2lk3xQpuhf
yUjcYMSZsG55hY3YM6gfINI7PdG6ru3vsCkEM6KoOCMNf51xuXxg9+Nr71rNHpMu
smvUPe8nIn8rRspCPTq5LxC5CX/X04v5k/C5XDVjKeN3YMgT66oFGiJhulJn/bHa
E3bOg6ttZEej4BJ/y+fJDBhgEDHiBE+CxApfPNu3LklwDRrRPcxC2ZyG8CiDZDTs
FTo/38ZjhXK7IngXaTA84ckf6RX5o8Xz9LqeLEA5ZGFWRBDylPlUbJXxB44w725A
RJe5uGyVcyDh6eIRnVh5EbIA0dDGWj+DRKIGlFdi1wP38HWSU5W21HJpBUNp6IsM
7sWHXcD89wZe/U9TdoAVWR2Bk2TXH20CAjDkI8hGB8cCQSWL4tRYwptCZwf5n/rb
X3N7epbrdaGuOfzRx+IQcQ0W3SliQDH7+gxnLV7kUz5QfdkyQUUKhuU7OPWcdn/E
IoBrhjf5pgeObidDQf3C2Ybaip2/zkdOKC0+jRO+0ns9HV6WQJazJ6gEQKTXdQtp
69t58yaZF5Xo08+pEZRyWr+paSjnbr2860fe/VEPtFENq6UHooOH7R0IDTL7D3em
Unrra0FnFzu2FeDntKtlxiLavJ1GEKssCitFwfei3AsgHEFH5zp9V56tB9haYb67
h6J6mwLzK83j/FDMaUoKo27fmFQmgSmPrMTYoV3iQ5CZX1kYNJrNaoEcpsJhYAoV
eE4t/J0LtYdCwBMN683Y7MWZ/3w7XZb3obtizeBGP1OpBzeuT7ssoO8nHUwceD0Y
3j1HX4hnwp1svoesXMQ+82lW+XISz//1aeYXEGh/Gs/ZzF/kCY5euwXPAnwr0Sm4
xDKtfd2NB2rEuSnL0XXD0d0fz5PPPaMm9lzuIojO4c85mxfShwNE+4AMr9oKgcvP
Vk3tcuaNJ8CWCLTD39KuIfFhTjPJ3XLhXi45+oLEuRznDwEl8T0ugKWtmvL53hlL
xONmgd2idE7yPxOvR4FEwa3v6qZUuT0iw9eR+aVtfoNHI0iyoAPAYE85m63zr7sR
UABxietzyXawOcqVdmQZBZEayat2ebUWwNlb9OeVG1a1cqkVYCjUI1Eu3UGXG+y4
43kS9AvmVP4I2vkEIzPs0CpqF6AD0/kgZchp8eU/H1j95WxdaTTuWo1Txl4cIJic
4dcffPbwAgkZBcBV3umk6fPb9/6qhxgj2fGgMXre+oOxksD3NuhgV02Bd9B/u3Ll
cmYpwfVoiMR6+RNUBTol40Y7l8W/iplXhRe/WxTLBbD4z1P8pV0Y4OT2WJ79t5aK
600w3QoorBBglRVd+Qu34Of7AgyjQY4qn9TnSNTDDs+10lBbKN7a1d6d1M6NIr1h
pKLTSJdmtHEPX7iRAf95tF3GVPaafnAElxWhMjr/RgZ0Q1s/D6/THLs18ZvcgcNE
jjvkUICJu9xBmc5RCizFIUYuxOBnFk9Osj2c+2JDbChMxa/EDHnDyjXJBIpd5uMT
XJaiQrI6cJrYHsnjoc5dMcs2nA0+9pEweXUPX3s40SL+j84Ks+dTkol/D4hDsdGp
6BGytHjh6EYkDaDCYtt9oiSnImT3nZ5pxZejT3dHux+k7T+y2st2GlNBpvTkbc4+
nw/ms3LHXf7Z3LCJtKCTQms6oRSZq0NVUbvzo8IoeiVVmSrznt1poDPU6MvBbK+6
wj6IBomENpDizrVK32qDPEJrmU2hNhDkNXLFUXOazuhrCGbEiieU3XEuvxyQo0fP
WeUIue52NZKGYDm2MYiU2ETt2r5Nu+3BrCPfkgCm9hMudbyKibLN8kOCcFgJueSb
ofO5ous3JOe1chWtgtGVouPUCzaBdRx08n0wY1msmHv9np4l+xt2iYjP0G8bd9m9
HrNVsk1S3tkrR/9CCUqRRDbawP0icxZv1F0icz/EDL7d51KS2Rt++XjNaE6PyxZ3
JK7jGYqE3Ghn04U6asMXdEKG+qlMqe6O7y1vUJMJNCsU3Fo1g/94Fk44ROVggwUO
Zb5qFjzDz8a/9SMV1kRx7/d0B2sB2RPSFksncs1mXlzPizvJWOkI3SXG1YzvwRhF
DRBb4Q7Q++AiXY99pbqNGR6conmrSJ4EnX//NSawNUOjevgjhXx51gcAa9yjnc38
RlGX49/muQOJ16FPMquEMnw6GaZY6yU/F4FJi85zQXVneyq56i5sllAKawo6evA0
/etUolO23LKING6TSzHzZTYaTRTmqGHt2YIUNsgnH+2/mPqQ+PUvCQrfhjl99C6Z
pKddXC0l3eBlL+/lBx+VrEJxnRjV36mw25Fxji3dY2ar46rFXLdfyZepLkHdOQM6
EnTORoMGfeGmzOOGjC7fNPRKUZ25ss1IGNeRvlIl/vEAI9Vhv3Joa2bEGqMom8Wk
gdr4gEQ4IapklqfeAwu9auKpz5TRaxQ6J6Fnvh9WtfGraID1CkIeTJTin6VKelmc
T5D5H3DLBbdCqpGbC9miYMjd6JJh9y5XK3DSR12AH39Aq5ovptIWwIyP2CXAoUib
NYbA8CHN7dGJnkGu7swGGnKk+JWA0Ah5cNMWS6sjY03++c5J3Z43iaKBfH0m2RYV
hYS/n03FKcuqKuXjN5J6o9UnowdwTqzjbGTl+teeAHuwLPdcK+mFXqIKRofCpBFk
+qcbBJEasxW9Ek8hI13lWc0fDB5ZUQT04gFcdtwqBjDjURgzZPU5XyaN2Rg7RiEq
/+LVW+3US0BR6gkNaLcC7HFsulRYLgeVrS5SrBERK4wYvWuXLOv3ZLZrMA72hCLZ
z6W/Ic3+mEoswiXbCdtzCbbVYktmPrBY8wfSdBGQuZlEjv4Mzzz6487fhlIf5lHd
GkixjpAO9DX+JtYPmpPCloMJTmzDNMP5DEr4WMvWj0mUITvqv/+acRgJEYVK+xRK
7NjC1xOd8jIVYVsWNtAmfnn+WUNnKFkHerZ1Vc/jualodJxEETEps5OUVkeRJchE
hXBxZBHgZXwm7UbROuy765dk9XgdSezL/Lx6C6XP5wmLU07PcmAQPxluiTmjHNis
FWOtAspm5o2n/Gdj2veod1sXwI2c8Xr62Cx/ASfIt88TEjuZPS7YCT9e7oqcvZ6Q
kHttFMOt247tHzlxvqcm31U70ClPmeQbjn+0wZZB2EAg1ax/BZoOl5R6RTrtiXN3
p5hyE5E4t3/sgC37W7RoEcTPXwPLSkZz9NibNzCT2ikUKWhh4MkgBWS8ya/Kh0ZG
pAlH7kBLiChk8p6RssFglJSZdRPFunehHRwJF6QdxZgFK6KJRHp3YOQgrfhF0vQN
qAUOLPsO3iEmP8PneuGH8N/H8GVybxNKlXdhFLRzfL5sQxXio/CNvS8oOZjOtLEC
ZUddIWsjzbmW9aXNuf/CRThCDADgESHzHtk5C4eR0KPPeSC1jQpJMB+cVt4vm5u3
uz2R53SshS7oSW4+h6KJ2IkLM8DYIn974xW1p1gKV90/7wYhU4nyUBmiLqiFelCo
v4xvnEPd4UJq04/akdp+Cgq5hyysufhwwSVyw4LFA5AYlDFP2vWCpzmHRIZiSkfl
kuSlHWxx/RebuYJrtdZ02xq+VqFVLjdas/qC71A8jYqoOKQVUdMV2kUfB+f3zU4N
8ml/1asi8luJrYg2Eqijfht3plk4Ar55ptSUP2FIu5P+HlP0s+839kp3YLFHCSs8
4Lv5DsdbBld+vyC3vGumxP+Cp9BYF0KhZoJF8fzuChfkM6lGvdojMmTKliMTYDjP
7ODwGlY8kwjMRZHtBU2dngU29dFxI5L1un6UZNIZ99a4GZ8jXFdTPPBaKRjj8Lt6
KsDtgy9YPQBBIKGIwdAduW6GHrVUqAo0mGe/9dG0w3nCD72XigAqAMziB3xHmmo6
uEa99NuoOM/e/+SqsikEyT0ixksthxUdpuEsDcS9aTw0Ljykpty6pcC2t6FX5MGT
b85yR9JiL9eZtEoRapLPRzvv1P1mNu1fECkMkGhYoIZY7j1MG9oPZTborpzmNDxI
FbL55BQMZVwzWLGVawZdCHvxD9m5vuNBhpKZmUIuIFZVibe9iWbilZ09psVn0h7l
4+ZUNl8T4AILqPbGh7OMYip0ZFdQyE+SylSuhir/iUd1cxBD3ZU0hZRW7ffsQwO0
TNEdRQdjeOc7FULOy/iL7/NxrZTvjlm9ZNiQSPIR/36P9Pp27a6Jzp5fFJRAWxj4
N8/acVclmZ6Ghkkl9fZcTt8VaQMinozXcU94UuFad/C07B3N7jhsIOTyAHkg4T23
k2HKnFshFHH+p6l0dzpFnhyHk2YL7GkS2BzCRO7sdFkrwgkqEqU+fq45e4ryKLLm
vl7UBS91fGO1oi4tRl0u95PiClqDBg2zjRwWYPH4A3DpkAlcHEnjzjWTUXnE0+fP
KdfTTiIm5nMmmBRjX/YjMdqHTJkMpgdGQPBKyMiGYxrld2EXW9/gu8USuE22DB/E
ImS1xJ624gGZjk82Hn57T7quqDdfmLGGWws6iUlcujobgrAh8oRJaYU5oBhV3nxD
/NUm11XWDfnw4UrXZs3sNLwfXMTsLv8hB4VZ9C6LnH4gLMBimgkLhkyDgKW8JIFz
KBAMve0PaMcTxsTo8PyQHqwjE6dpR1U3WXWCgNzpdokTrNpfopa+Ttc0r4S9jgAd
ihlTgWZd7wgXZimvJwqQ7A1d7JZ8ZfyrTR5aauD1TEA5jZc0KUZYHosc8IwgDuZ9
XtUkzo8vPiSH+QyJ3F/Ese08HTshu9+cdIiKKTS6wAbMrm9CLm3Iu7sucgSNY8cK
vOBvgASBeZ5avv54k8iCQdbzfpjFCEo3w4cL6r3zJJljk5SrQ1qqpjt7e8pmSXse
htJwvlIRjYs8bPMCQQ/IVTc2lLgYI1nIy8nTHNa7gMiKLyJeLCrtwRjAuooB0Trj
uwFC/HVQikjskPy3UKyEbIUOAcUfwsRZ2QfVMdvq/QsfGQ56YAiPWgxD1zi+U4zB
LJPHYEpgS6/oCW0dYGkmCNgk6HDwHrQLm6enZVcxy46dci7o3BJEP3c46bnaCE0H
cf02rSM7eD7rRVr3IXfXEKyTtgMVCjcOeQdpX+cqeh+2mUETuCCBGxwTpmInT0YD
A2I/x7JARcgvq/y0rIk7Dl1rnvtOYMs/U00k2uXuDjWJeGnUZ0ycbaYQyHjHF3O+
cXx3DU0DdI0wQBnDUNecuYc6ub7ZK9pg73xkKZl/xZumCB+lCZAk/xIK41ug2aUj
2z929ex52Lxydpw2IIlB90PEv/o+URDN5dZBryKd/YvcTZByMpXH69NEh09oJpjG
M/7liQHWdJOznFBD1FCWMUwsb/ewi48gvHaBCjyotobGqcBZdIgsp67vxOAeQs+u
BbZE3aJOHpL+KSEZGhFPQOrsMFoln0a1yHH5jr6n0hQnOue6eLlzkFsNB0aKBY0/
c9tzyH6ECC7PDPzcsLHfs3ZGlYSClF5SJxS1RTVdyHjlxuSFnzORbs3mNDbfNFMN
Oia2XN8p+RvC5pSCFvZ7lWo4FKC8WN74E+kgk7f2SnPxIlm/0vusILcOsffvhzug
0394JoEu+TfAPAStzLj6aH2ZPC0UTUvNdP6SkxbHwMBVTTHKpoP/z6R7OyLLbipm
uq09i+c9VNKqL7WG96Zk1LK5jp4/mZn/md3ZujIOzMQSCne6VK7A39T69GISpouy
IwBroUW+1rofW9A2MH/vNng/rzNHiZjOaR3kBBocshd9A0vYAvkjC6jz8sSbABAP
+DLCSZrRupxLa9YNl/dCRrDguA1gGKU86X5wsYwyVSNF7cdr3e8SZnMHi4NM171n
+cAL+95Nv2OQhfy3tBBIfee5AfRNvRtJfqU59wgaqTruxvJPFpCW2z8gcisgnOC9
J2S72NZbzzXhcnAgQNCocR0VJ2A9cHrFstAxVChWtyC7FqsjmLydq/ECDLXSEYAE
imAl7Kw5MK63t3FrReAwipEq0y98sE2hOBPamXzRuFF4agWfDkSRqg8aWK2OusBI
G1N2jgfEu5zfED5eiPY1Z//HGtjpe3Rrvc3tfx6U/krfcuAmhdBlPTCUPP38l3od
miRVA/iyP2OuOfx9CdTLudVPUH0q68eWhs3ia43OEceBnwfX+/2oVdVTQLhX9hWN
FcEGg8tbcDr9FJlpO5YDyTeedueJzgnmJdeyZh0VWI1ylcnvITXDCtk4E+iiEQ4g
c9yqzy/onYMbh+gRi1id+Ko58GmczQ7Aex8NLvkVPnxdwkMDu6xVf8iapSEP1R2s
tIZyB13xxdjnR9X/icJMaMEQ5tp61LFwxvGIpCak8lW+vo+ciUj//N3GCCEFTb2O
/tlEeqswyuraZBzChoTZm9R4OjgAr3xExWR6b8Hui9Bu/Hosc6cdF4rqhSXO+Z5H
ib+PXs+nlXio3TC6wY5nk/gv+yqAXK3BMgOuehBwz/vweqljxkPhBR0RrdZK/olq
bZagHMqgdcdlfh//QQKsjYcobmC2XNu1lvnMAu/NPMlVzVCOFTRo1AN69zJ5Ll9i
ATp+nE7rZ8PTFYpzJI1vdR/TtEDi4HvFSIzU1AH4q5cj+1joo7oM7x8++PLT5N66
6EYMghhFGYSM2Kh+ffyzgwSyBiOH+HxI2n73Dh3RyvNCMA6Ch4RpQhh30yo+0fgj
MsXDtqp36TEfSjbJNanV5c3sIq4K0u1BsfR9kfxVL0CzNt4LOJHuefadXr3yB/n3
ve0mgrVZHw2xHkVwbXn9D25IlKEHy9UEL+WUFtL3KkL4H+OON5YORNylJBR8Yjjn
yUpgE00QvYitxgAPyAQUfKHGB07piNigtseqO/58i1Me5NARjSf4GQg6AmBwf9f0
S8r1OW7uUkha5k6skkmM490wMEeOCFP1IzGCbSiUuew62PnODXMA7y4CGHDaTomw
/sVcSEoEWLoB/MtxUw3vhiNMUyscMN0mbD/93hhxi9jPNCG0CXoy1C28jVzCty2G
Hc9r2lXrAADW1U/WDuxwIVjqSdnJE7WHL/ZpmFT3QcNpL/OQ1bC7Rg9Rzo+4Sm5Q
dqqivqfde8w6TYvKcIWn62t4HQvonDFtnR1ay4SIrJoqCFPvYxWhXG95TJHeuz03
20lj1NUiVy5wVFmkeDWKKICxu8Fr7DfZXRodZiSUqdDM725M9jzWl7SqcdBHADeE
kOmQkXseded8C6GUJBLawrU/l/27fNi36jSFFfSSQ8oVBE3fe3Ze9Clw1OoXaDL9
RZMcgdHZkZK4ABaYCcJNncYdVDNJ3ucGuDRbxGxaZWGxPYQixTuNHiA8js1UKkmX
3zTpq8bemeiRZqb8V7gjeao0dMUey8Iq9axaKI/KMq/X4NcxzRsMrXy8wgPHZoK2
DsD+7N1oBW5awVW+QflMgGRwhWJRnc0/79KcmrD+1eGpSbGqx3YgdCGMh1ePF/Gs
S7NBvXzarllTDjbK7eUs/MurzJXPG89NhoqkspY63y3xcO/nh53J6F66YU08u23Y
3KsGmNTNCYCFf0d1gxbw/wQgQGuAFRJB2YeF2ts+SHp/7zhq+FRAhAe09d39LXLn
Yz18GpQH4nX8VbLG4exXQcIyhdE9MmOjjEFVZurOqok7bfIaZbcf1eIxq6DHQguF
uWTyoAEyTIpLVGdqV/8//fjxMWOGGDmq+Dgico/RSV18NC1Wk5cctVgYm+L20xDF
IdSeakiGZd1Ug4u57xBTcfDi77tmIjTqG2GUQAJvJGImHhIqzaUTjF1rLWwujKak
aa9qJRB/TAYOTv3udIOzpXuCN8q/Ghax8gS541w9AL2/vugh+bxvwyb6PNvYG8ZS
OidjchojChnSxSQI21kc1rlf1USUPzY1pOtOocTIvu7bEoayIdrxyfKxFpVS8ffc
b8E4tCNZOMLxwxZIIotf+xWDOqU7LP5p+hVkCzpp/WnrSa/FSAzhLaCD/6sQEmX1
AtdF1+IWc8v3JXgm4HlR7Q/GAD/vS2DabWhDuHtlQL+jo17isrg5d5gg10vGPwol
8ramf9AxjmJKLR87VDtwx+fTiDaJ0ERHZySyZ8NPUhPcdIM7OtzpLfr8wisxjp1J
1EdkBHUyJjHZBEOoEjjaOuDWOTXOGOANACdTlOEbcfSMo+owL3KYti3H2J+eUXju
t31HdaDIW+P0rwmtDdKM/RAy2g5Mq77F/hznv0GfA8U+zK6Bhyf9z+tC4vymUjPD
wpURpYmFY+M5wRPmWwM3h5/X+5Mjp9bNbeVapRQ48YvIShClAj3HjPV+nK7LY0TI
irsYdu1xDev6en2XPrkmQfxWewJmwENMVqJotZGQ+tst/Y/kpf/7PsqjrivJheHw
iWzQ18ZkwNkzDe62bgjRQS/wBEyO7yqgvCz6FndkEtt9girT+I8HwnQMyo3wNdaf
usEiI24ImVhOCuPVqoS7OuvYeaufqiZZ77P8p5s4CYD+ITc5OejRy7pX+J1bPDZQ
nVc/IGDOErpsToHS2iZE01fnh5zYfagIshmLVzhV2Du3CS+WrZUDozzvFKVzfnZw
p9MSFe3Afzaj+iwKjRIkaQ5DOUu7x9A6w0Z5899NAh+tFgDqkUjuFvtUsEIc1zoF
vMOIltOY20ho4SVj29Y7P4RxS2IAxdAfNy8IDb8qvQPuB8/Q3TSHJr69h0vao7Qx
LQk/TbEAWOHszbA9NUBGlGg/mO+dZwPUCKq5I7fWTpEo/3ORHQWhEZaJnmBBc8EV
5QdwEK55szxQ5gpuUnq0T5AxMhQ79uqIn+F9MsmPY6BRjQHCXIFHyVqkybuQug8/
CTXYquoumGm/+U5pvp8yKIHqRafcwWBzNjAMPA6pWAf/pu44XOueh/soJ9dzeIMa
iq+k0TV7AarfMnWNN9/3G8eVWCBTnaoExWsvRx2WV5Olt6j64lpbw221pWf9W8hw
r+EYRahOxOSGj5VH9Tb0kdsspMKjA4dcFqeILbsem7TowQTqUzJxoVvkFUTnycj9
zfCtBF+xmpcc1kiq+HMmYG+xPE/HjeXvi60OsNOfD2Hnqji2Obd6ASCw/keCO/cI
uDtTsUK6B5/9/SIHfC6iz2mJdPjx9JtwB+LcdCX1iinEyq7KVHdPvamYjgC0wAQC
IPU0RaxGLpQENiLF0SqoGHZcnf/sazEsUo6lB8RKl8sU56ln1c3lUQT3G0/+Wgj8
J2IjWK2DYHb/3vSMsCjbuaKFKdir1naoiHwvtXkFyyvdwJ1DZEqtYru92wmFl8dB
vf7Y6htHPofUIADXtPgYjMmUzktkwBduwnqijBfBuNhfaAth35xPtjZjCIZ0h7XD
2PRtO6tfAbPo6stiLDKaxsJLssCNv5H5dwb4bs8RKLZ6W/YZkbK3AU3FpoFareRi
9qIMZVQoc24xcrsQI9q9wnmUsayxehoRLxLwChFMXjzHQazPCnkmjP+lzkffoPvY
uO0b13X/FimvqW8m1S6YT9oyFcu06FjGrnQ9AOScDnS+oeKqoAH63KWh4+2qVAw8
udZGG8X4p/Y44YTibfJ8wBebn0BZRze7X+cwAwufQqlazimPLaLmwcyNl195kPBv
fxOv36sHsfrmxJXMdLeSMZDVq7xpHPlbpFixlHYXAGEtWyczYXE6u5vxMid7ndMZ
46H7TZH3OegfSdQ801sA/cMUsT/ZecAZ/t4SCeEvJlZAYukR/BHcLWFHfV536KWY
qo58T5IMS1yGPD2MvyRswYu6+sLbdjwlP7kAYfgBzDZ0I+iHGS06VI/U19VMq/z5
x7wdQ5pU/KaTs3+oYXuJvumxZFfEgFTUp+E79RKWO7lnDW3SJZo2L1bVAZH8Wmwn
p9pftPqdl5vVG+YRPl0Pqga8JofOkzT2ElG3wR43EMvv1DorPz3WLnbtmvt4v4+a
dK3DuXmLgc8KiiY41fujkGGgDObGl9xrL07phvTEpK0OjPKh7gVMwJIerJ8L/Wzq
GpKr2yF3gB8burNdkxig/Ra6N9BFzT5oJo161tobbJv9NMC1EwzVOzBEUCgVaSPf
SugXUC2C2g+r9bi/7JY3JBW6MnVs+1Pernv/EmOKtQVnXHNk3LoU/5ARxGA981Uo
Y23jm1ILPdOjE8t8wty3njlmVRXvd//iQJaFgQ6AimUAK1NYeYhXoMuo6IW6dyVb
i8ffhOvJPjR1JGLXb69RMKoNvrea50KUpn5UcVrntvZ7ZGDFvcRSQaJZVBmf3S5D
xPQ2J9jUICyNt8Hq58RHfUy4W/bSTqFkqo/uKAL7IecYQRLlX/u8/mCAMwapqKv7
Ny4j08ADuuJBPx6UscGbNb9OWfRwqcTU/mLxggCgoDu8zlgcKmZ5UwauvwkBHSCQ
3M1XNhPtiPOe7FLv6HUnj6qYFvsgwIaghLWVcIYKSyXq++PxazxJom/iWSPNgRCA
xpu8NMdN1jY3+eTHbT3seLPx9t0g/G+mHLCjngP7d6WbMfEJtP7Uh1C4kAqyqRVZ
uXKZN3aR29N7lK/yiE6HKisINdxMMRLQJT4quEtfUQjf7EZiVWBiCGpbMuWF+MkA
ifmZKfHcheniVYy+gdX3LP5gSbFwrWr3B+bmEvoQohZq81ryz8HZ+MojyumhWT/7
UtlJeXLbTyaewPqlm3nXdfhhVT2iMes+w2y5w0Gv1WS8D+dDEpA66qrRulQXlsjd
+HY/9MpmBG/v1QQhwMoyZd/6BWmmHC0ypzmP3UYoCFIOEPAPr7h77g26vnKsmDnn
2T8u0iloMh/e+aCadtZNxARXvm3EDTxSAi8OU3ncB0pIWZ5EvWHwNuEiSUWYhLEX
w67ytDHkTjJy3aZQbB3OL5SnRP0GSFw8F71cKl/u2eD2NkYVYukHnMrzVSXCXthI
ollSeEVV7zIFjc4zH0NFTs2pdhHS+Dz34TU8LaOkSth+AgGjYSkMrHec9v2OpY7p
/iYlZ6p7WsJ2GjLn53rjWatgl1pKdxmv/5ZlJk2lB79rLHGJLvRhtFj1sNSqKuwL
fhisw9dUhvSzooY7RKsO8UFSMsu2YXskTI+zUypsXALXDhnjkO5Na+yPmf6/Nf2Q
LbVX6EaFlWqv1k3i+cQzXi0sx9m1qZZEtx40ZVg5BU3RDlikOHqwSf/zcLNOXSyy
X69C0tMUjfbs4T9OTvWdvuWdKG/bM1aXZt6QD8Ig0op3ju40vpHiN3qLgL/6W7x0
Gjjk7rm3Z5iQqrjCot0DdLszbUz+PgQoWFM3pil2BE+4BZxCq8g9+YSuM8i1dWmX
uWvjOwryirHCxvs0ikaFNogJJDXu49zm35o45CUv9+8RAlVSDIm/0QcCJH+4bbGl
73CW3GMBHgoeClhCOEOCPwZe/9Xwte8xiTqCxhysjifpWBVgmtloKQ+114ydJ2Hu
azTpdIs0QtYnRJDvHhvpF848cPx21q5qJn/yyt/bhM+yJWUtvvIWOh8+MlFfXz3F
4tocIHOf6CvjPAlzZhwjAIAqX3hVk9gS+gDAG3riv2aSO5Hf1Hi4VGJqlhgpeQwb
IqnCeCk4NsZQh/n2KDoS4l29uVnGeNf+g1CuyCaIgM1kVUtL213Lik4f5UsEIoQl
lvoqpI18x3m1/Kk8IYqxK5maNvpawKznVpHrlylWBgDo+5XwNtakwFsuxGenn76x
SlrML6sD2fLweLYJWbuYxNI+mIkGhacrmM0K+iCysQhGbXRJ3Dy/Pt07A+TD59yi
d84JPIBHbrFmQ4Hs2q1RNgKwA3pQ84DC4pM/jEicI3cD2HBGcoThY26XUjof0Nj5
0MvDZiBcAuBYCu3KFYyJ0EcUIXmyvwq0t5xJZm2T+iRf9D3mRSsttd69MExUpiUE
4EQ5lMRNASq0xOnKajiQue59KFTgwiJgCxG0v0lM2jFA6N6Kb9hrTi1UCoXbPZXh
h9ZA3z8HwzomKSo/pmql4BzNFvjILR9XsvVKI5rzGSxvhIzx4sAXsvTqFRKdjwPs
kTWbGunnYnUZvj1rMuoCmmqtOyQNQ9f3KSYUCffGfrAVFwXbcCznkx8uuhevrIIo
Lh7kpgVyyBskb5B6frjTp9ovvlpQ0QIa+KEXnz6zftMhaK4wyJx1GVEQyrZoGflz
KRGMy7uBET1gim+szrtk55ybb7wKw7DONFR8VlyQoH5NWMnuwBKMQ9rjAXW8R8mo
j8X0tlp8yxkw+VfMnrfvU1EGir+GGFuhn+y5fHkpshHTJzgoA2O64FGNB8EauGah
uvDapCTeAbkOa6IPc+qHNP+1rgURosfQDzMiCebfhdudlCZfc36ZG6ie9FgzWjry
gREm2uWoikVER7kbvVMUTt19+m1fcWW1gKxFCxMo9kjWuTnwFLDvVMKGptjZlHeh
3n1afk/4VQuiB+C9DtkJd9rKgqENX8XhAq8NiiHktZbjzTjCL4QyfhlKpSVRzlb9
HfUS1lYZb8Zv1hKfs2UFBgIpfYcDyQGMxvVFY/oV92ZrylSqknY3loDhcNtOXjJT
vrgW9L/h4ZAYQBSr3sgYAh4MtzgYW0OG2vsWB/qks/Zj7gLkhbDpDgQomuwIQjoA
Hj5PX05THI3AAtN9K4MMY2PTItIICL4EYvTWE0cAojm6DnQLUFaFPoc54qyvzW7m
jTTCgFLFBHhrp29hitJDnM7v8hdhk6JKKLnYoZNb8XfIIRLRuNBtwp047Il7RfqQ
mfobbNUvUXvD/SQaIKzStSycmzCFUREfjgyziJUoLhkw1daqJ2chNRHsJVqhwvvv
TfX9lNjuTZiMUzCekhi5EkpSiFOK5oUHLm2iIvT9exjbo7ncpGNeJsXJ96oJ/p9m
7qOXalXgRy/yc5Oy2WvSwHVeldrgG6ixIZ0B3KErfXXFxDWjdXo1/GRDWIGaZyIU
Er3n0FPeT5sv1WRgEUgDx+Sslbc8z5y4JUyzOXEwQclLhknP084k1GVYRJ0X0HO4
uJqRdyjA7WiLbn/t10IYwbQ20QHeCU8JVfE0xC5ItAtm4QjtC4LutSLunQJi2Smv
OxT4aQeD1FILWlqP+f+xkj1OKrp8W1ra10lorVqdDe4Q2JhvALctcEjWHtseIFc/
s0UP8q0BrkLl5lYnTCi5drHu1VhGtPXo63+0L0yTeR+RYaJJi1Cc4zicx0wyRO6y
13IqgmWb4PaGVLy/yMIdAVy5HRTCVXvbK+8G6B1gRsyePkjbz/AlWZVMSvVL8vFs
IRTvwo2VEA/hRcpLZwQD+FYlF7whXnoCGYrqzwuJonP5f4IN83N30OW98DY05G1u
qE0DEmopmDMYqN9XClmIvk+rrtlmuVDFE12unzHQdwpLs8lbOb2U+WNaO+3+fKJP
HT4BuuCD70hmlP6iL+9IuPb2hu54jY8qfWp+p3DjnqbaBTR8pNB3N8+rBAgiuWtK
PLRMLudjl7opTdvoKbKV2gO9wUoWTJ86K5rkw4pzb2K6gI/WIM3aG6mhYpOebtER
3gEdfvgajbgqqprCAEsTEO6L8seLDAA+G71u8bCXgAzk/oC1v4D9pHh/9DFeTZgP
rOagsHbewofxUqUa+5MMKnFABp5kUTw+Xqdpwno4BDGXXCUhCtf/zV6959l5rvWW
XtCLkhlWopMsnnH8eoAqriJ8CqQbqCMgiyLpmRfO49oTtevBdrlkU2v9R5zN2eTJ
u0YJIOx9eUxKnnu5Bj+ZFDtDRCMcregAq8mAxu9dvs7X+u2PYJUDt/TmXBRjauzK
lsD4tIk6tQl4gnvlXc4fZeMsfA9dRvtfyzvc5LdDm1TLROVJ+KKrHEL8v1xRpg8p
kKYSs8FF5kcXVW2cElcU3F5nBMb6t1wKZZxeXZpvnvX9ZcZl1abHzcvnl+4098ZJ
brTDMheyjcIzHSY8a6Ai5fxl+04TEpN/T3nBXnwwAtlLNs92a+LtwCkWGiCJ1uvg
mVpMARvvZKMKmT5OT39m1St6Ol5wakrP9U8JaHaiuTx19uABjkT0sn9Fu1WpH+vy
fhGxCZ0XXxazf9H5tl/NaFOSFlCJuXhFJD1xM0xuuvNuYyP6+3XMsSPCp5c8fMtn
WckLB44Ffvf4+im4d/ueOIr5LdpPXJpidHTN08EDdouTioei83d8BOLjwtQTDde7
sopKcN+a5wckzAWn4mWGpR8LkrYne9FDOHlhSxXM/4oQno4STtQ7NWyHoI8WieU0
HQFqSzCNkfhY5e6YBrSWMdQIZIn5b1JNleEtdNocJa6PhHCGp1wSLwg4h+vrP47O
aeMLZv2g6fn1akX/MHLV9M1oSHgsYrwFRSuJrETADaQsud+R6wO/X3hNY6jtKxRy
Hm4pGK1sYnJbtv2K2F2QNjUbk3sw7BjrWkHKMSsVabd/hdoO/HCfBbJ337zEoDBo
VI6k6OFZKGlcVyGnXBQkWXq8QIJnqLpn9jd8pHyLKk1foIlkxmS+7UYlGxTTnmP1
6fpCRRQJanW38j3v5h6zrK8WIZNnuXdkwgRZVgac7olAP5LSxZNR0RkcgYsVgnQR
n0fyiGN1GFvznFOOlR9BYuPaYgiU+CAu4C1e99DhOlcdvj709G8cK2chreDyOOKd
SKuO2qIXutXf+i0fyHDNhtstHhwwAEfeiHZ11DvhgF8VFH8XUEugJ7ZPAhI/B+lH
kSb5FicEHg80Yho2fI0dE4EhVAZndOVLtTxbkFoqAy8SVGAjPQduc7Qa9BgWTzpf
MCillUF0QODXoWNgVE8mUyo5n3uv2qvksxUJXrvUXemSNdgQreDKaSWy73lMCNV7
KPBG1bNegYMULkufjjl3UEv4vHRbmZVf1RpEO1Vqp7tZplD8wFDpbNvbe/Q7296C
xUSuG2gG9J8+Azu0uHS+jdtU+xzuKspZZykEL4M5u7DJgIifpgOsQJ/JOs9kqcow
I9ZKjfbE6ofi9njcM81kWMk+ytp2YGUY5DAr8hROKbw35bs+aK+Y2YvfR5UhVJ9A
x81NRWtoxPcQVtKK/XcGuFSCswI/0ZgBtcnHOJN1og5Z9Ct7LxU29AU76ztxhwY4
PG+aYJWlMkMw9zhS+ZrVE4W3FggM02UB4TwaRsnPNFyRoHlhzSVKoo0XdW8OsPik
ZVItmlvKgu3EhXyDjlj+OGWfBqhVtPk6oijs9ZmT7iblHFgVQnV/1dYNFPFmopKE
tz5BpN+kKxKV21YOLiF1an6k41nDwD96RGdoYfg/+XT8571O1LX6XINYXZAoefXf
1aoB9JhaorFrLpQ6vHE8kS32ikweQG09GksXMvO2OeD/nZVYHYn0GVq2Cv5JZ1Zb
HYm1i3joMORQ4vEfVFnVhoQ/llmlJ5gEnbL/RfanBHBF9E/ihVET3jiypDj9gZGT
x1J28VINIucvhUHumiBVTuQQm7Rv59osPSih0USVMXKQ6lZlznSDG8NALd5G5gPG
6NjcdS0wUwdQAyDCXUWI4XweTM/Fl7HkcIap4r3s/g3LSFCgA+JJKn/vJtoGPvRO
EMrHBa4PKSQ2TOgnLOFAEic1KWtQS8HyI7+iMHmxyqZRvQDHjP0yMuDBhWYuFJ4v
f4ul3Qs13PHGhlKdMP7pWd7OlRfGY7ncDttHn/UP8F1A1phUHwv+/kLnhG+RSxAr
hwwUFnvgHiZ/bx96zermggO+fkYcN6fc4Yf2XspKFBvBnMHg5kQbUspBFO9Ps9Wp
ghuEkVDqAqGSf430lykn2SHhJx7x6LUXghnjjpMvbX0Qc/j/YZxLkScJeq76/YXV
zOHHXUKEEZM5DlzoP4kfMb7Nu+E/SnOHmLgPc9la+5mLGZRla361xjuUy7AmpMWT
dT4qn4A8lJ0JR54Km81n6HOlQMvR8MJg7yXzz8J5QBG2m6fDwwfSaFaVnZPRs3m2
6z0UZ0ydoO7sWot45yA48rSOHpo7wBbT1jqY6UumaPqtoBibdV+JpvJmPXC+dhpp
kA5ixGU0z6HHuT3hHB5XW4GcC0/WlyTj3PLd+KnsZWaHEs8PCzcLDrRQbiJIQyCi
wRisTjJIChEODqSQFuGRq3DaqFQIPOwU8oZv8sUls1sbdzPeVdsibJZqC29zcJli
fXgOKB//wr4c4OVINH3IigZYjAagZ2DEm8iu8NpERCeWo/FbD0TFezQERr/IRCnL
b/HUzAZvLWWp4xp2dIVKaHVhjR44MtcMcefzp9Crp5h7SP6wiwJYIT37d33ffuXN
9EQwo3JsSZBKMwyYVy/cOKXuQ3f84BgDpzgexkcP53kO9jcj7PABz/IHHSuKR9CT
GJ6ESjS7QaHYBa+gUyg/H82i45hdW7pf7EcZ3cRkunzniJcfNFFbm0e0mYPxmXOj
iEVVy2Rok5ukks6WgvK8E0pqowpdFbhUZrdlKY4WLc+Wty+fTHj8UNRu+3VvQuSK
u5zTGO36SxZToiLJ/S5bcRGA/kXeJ5ATJqvP8cX/a0X89yQuZRti09EwgEdMMUyB
l2OYS2cake58VFtcWJUhllXMHC9XE00qLEQ+L44gJ833jSHP6MFqxhEThbeYfMuz
q9RZghi+4nxAkvN6MWQ1e3Emc4sRsb6B1/V9y/3YdrNDnxXMcF6zzcRP2RFTWHlt
hJ4fbKFa64RG/pIn+ZctRq/1es0XIszSDB+VpL2p2FkT9v2sjyFFvrHUEg+0zXzk
7t2kgJHN79uWivMaAOVZNsptlZX7YycIth2PPobY7lyBNqvngyuXVGE/TfB0CclX
URwi76CL26sKAqnIs8S/0jVdAVoorlwAnm5uG5WWjZifOi8bJSY1N4eKrFpScqQZ
QMPlRbgPJ9sy8YiTpWCPvTHr+Tidgw4FEAEvdxYnUq1YYwq9H9yszHzh5zmAt6vd
FdP7AGoV1VMiObDxZWfldzAT1PPTs37T4cJhER0Q7bqoRk6DWbQARlhI1jGqGH0T
hCUp4VkYljWi+B3BJwzA0+fkez0cK5snwruXjl05Iqt4y45xC6FbD7eBzKjzR6au
ZZbDBhmI+iYozxV/XrUUrNzMf22J8erLUJT9AssRQ5EHypCaj6RX+IDkSFt0Wh2F
4OT1yoq5X2CJqsSaoBw0FV3PYCZ9lid2XqzoKsx2oUwfWzmstyqeMSfGF/WpGWzw
1LtC+79UkaCYA2xKCd8e+WqVLK7nHV7wXeWGpVrXKZJpKqirV5mYr+BkBrhrb0N1
ytftroUJ1SfhpP4AhrKumB+b4n33xsmjlvcKLR6vmGfxB6uLVKk0zX0XkQDetwJW
mp2cFsQpWMnUOEpQF/Ct67eXlsvg31HKCB/NI99z4Gnk6REweBcEOJc9ndT1UfXl
i7YjMpyVs+GR4Dz3YZ/ku/oV7DeRJDajh6vuQO6IRqf5nl7Auy3Z/7Xt6eDgep62
l3dlkgRgX10lvZVPn8F0ztFdHn1u4OgciiEzBu4a7hoPnR2PYj4HOSVvY5AFANPp
NAhpp54GYoUI4+Nn7/c8Hk3Pq5zp04llfmK+xarRL14iA7y8ItxC5FOXHZujs0tq
+6zpBy6Yz6ZcWzun/3YEYcf3UVr4s2LNLLC/fqOwzfVDqYGAq7SM2FxMTtfonfxN
EszP8HEW3DNpUPRtunFBPFl/BMmTJrBhTLs5d60QZP8wHkyEPsnneHR1ofpzPWH9
Uis8gv6dUo/F00rtMDE6EfUpGIQmsoOsSVJFV9AWNCqnz9XD7AO8uxHXumUI/vpB
ZGCztwhdAVIch5xFyGUokjUYFe1GfMqGhRMw2CPVN52D3UVyHNapJHbEoYS+cceN
zYBVp6CLfhhqFF90Lk9gvX2Y9Yh2b2TEz31rf7slSkVMr6IlGho4/vcGiM9BeNtg
M0nXoM3Ihd9YqtJVLsgwSocLmY3b3VT9KpaXeV9EFEpms2CerybxxfQS4ktzi/JG
h2Q2ItcXr/u3ZlsbY6NvaGLzS2Gr7/4aJQ2b3nHPuW88goUJpg6Xzb02otT/2XN8
M6HsfyR6XmCQj6YPfYVugx7Ep2xIYekbOH+34p1nW8rieg5FNXr2TLygxL3tWOUY
k7az5wqfMFa6R1ZqcALJYdGVMN/3xXtpOTAixYb+CQGAFDGo2p3N6FlwDBpK4smp
knAj46kaOtGUdnPq5zvh5e96mPtuRcu57Q2ISh4hJ7oc/qEJ2kcORv59PLF94kYe
wECmeoV6gp8G0ZGDhCyD+qcHVnOBAxMHfsHd36kMz35WT8waPg7FvBgq42w7qfG8
euMeAPhHKgLViC8wJ/Bd/C0/vdiQMzsoYrHyucyDbvlA/xWL972A6VX1a6brS+aX
BwSAEQJC6eSv51zKTg5G5vGGoT+ek5Lw7qzBtd/ZyQSd4+0ph4VwoHmMootMxvp3
se3h0VM3ITFEkviWrJlx+zTuEUeca7R1N7NrzFvxXrQJHFLQd2RJsc1xe5H7B2hL
y/8izksAFIu8DucwLoBShtvL8/iwX7TsGXop0TbpLgJGfUngGp0gSWeG/dVRNq5F
IugkqQIeOS0UBxc6scMan98tKCnINUcmZwTL6X8+xpK5nueIRCMLEnnB4JMH8kkn
zkQtglgAGfNoonUN4yecP58IPG91QvA7kHT/Qr9soaDjG6e6jfpg3ZzGmhut7YU0
JnolMC1YjgPHwxvU9tWu/D4DI1KsMWFKO6+mpG2hPAhAkNNyruswu7jhp63PX3rp
BxlK8XOboDCm8Irb8GN7ueAuKMF6lUCpkfoAnQNpSuofL2UI6IkbRgo8wOSH1ami
BSYCc7qudzTqXJGLrN1nyY9oGSyrsoOR8gv4eCa0bR2B7ZibIZrhwOX46m5rP8jN
0M5eXn992mljLIhb+b4mLk0tPPp6PVjNWU+2KLU+BXq9xk06Nv0v14RcFolHrg7r
6HJEFGN3phhCCF/KbzDmROdqNFV3XLUmdzkavCLewWPAwPd3UyA7T2BhtqYtnvtb
1D9r9BMBWJHb+VWcGkJAxAET36lnyCYmK49UBpd9e+ejvVhpLhifXtcAEJyKYkAx
PG31v1sbQUGSzU9WJOLNXTGw7AzS2MezWr6RtqDH4+jtfwErI0D0EPLX51Fgv3kX
m/aqN0cPfyrGfKYuBDC4Siet/whG8EGnp/Ak5BbQcX8P4qcquk/HNOk1NCuopcyq
medxXw8/7f9Q1uaiu9adI75pMd1bgQwLEHHv8onTYnJFn3NfMSudokI7zh2LZ37W
CtFR92uKHybSW/Ms6kYsT7ZHEU5manHQkNwP3CfPTSBVYnTKAtkGOWt8rYUVrzNy
XXRD8gU3AIm7GK846nejCBu+6OBTxoqEZ2Metk3Fnj9yC274HWFd3JKjZ8lfIqu9
EzEr5MewvDtTWELK/XmvIrDV3NFRjID3fOXtRQWGfXaYNPVBYJOWWSiTP6rgUBbz
fK4KudxOL7M6cmXMvcUi7omKaWuYVilOQgTxCq6TSHL2/Yo3ABE32VxxlCs1+M1o
RTncbkwhxMQljYwJS++Gau92h4kU4sRJLkwP6vN05/27OVEcHsY6QXM0whsdTv61
zKvX5qq1XrxSLQUihyzXZLYmfIsBY6fA0V0zOn40/pCakNxYlNwy+MN3A0HrCFSn
zH6lDtixjS0O5GXIcVpsj8xQ7/MlJAye6pDs2yBdsiUdK76haIxDBfZNNvjuRBDk
GzptDAoZs+OrnjcsdsW9nSheDtWkpSRqcUlEPq8sX3LUtdpkNClPoRw0aAr4N+LH
d4+wBQ2tomE/pBi8ybKq+hgvBFn/e0igFVZ7Nxcw3bCKKBMnIl1zGfyKXH3zJxhH
b1Q9QGP4QofmU8ibPRi0L1O32JZVfP0jhQhsp3LzBfRaKfCMXs3dOLc5kB8OH9Ng
OG8/qDBatxtztEjksph5xnwN4iFrrFeSlrRaG3HNRQGogNOOK6sJcB3fittIsYyb
Xh4eD/NUL6TAGlOccWQAF/9FRtKYbq/sggcFHApPfSF/y/oD+H72pZuAfB10/mCk
BeooFJkqnomoNF0eyBpIuvwDL+m+D1i0wY9l9Uge7T8kkXsC1QOdr84GqUpNjZvO
oq2FlxOKEG0D554BrZ/bo0ZeTwmfO5GKL5xz5uVzOciS1oenDLnPicdME9hj2x5r
Vq07DzRMz9QqzDGuqfzI19fuO/r462H/lEBBGPuhMoawS5+DvQOkn0uprkZEY+mh
wd6C2Lp8QQboO2t9bLrTG2+V0kMNtOjMocBqaMt0Plo3/EPaEUHNM9zuC9PFKYJy
6GrX7DOkrxgVaiUSFIWMAUOxIiAQC4m0BJpGMwiR1zZTNTJqlfSDSJoVEdQW4paZ
ww3YNQiu2yb8pfm7lRirfxjrx5bV7MQF54iwJSjYKsgrO3kz//wWcbXNNV4Ju9fK
tzOheRFv8mVrLDA9OMMgh63aRo+EcWZLrRsLQdmO3tbQ5lN5rONldhOmZy6GHzBE
OxTNvYS00/RLltXy99yl2QOimWkkiuk9d5ClQT8oXY70SVQsDuATuQWN6rciLdhx
2JKCsIadBHe3nvU7G0gzxcHM0EB5lj7fJLXyAeIMxJYlsj9InyofEA/qGzPpPYEG
SE6NJvXk1A4O7zWnEYhCTh+u1R+jYVIYcKBscPZdo9Ko7qWSelYVsiVv6m/UkUDz
zQpUZ86MAJEtg5l/2KVfFz2YfT68ZZHF/KVjp+XNWVvT0gzzOn4XTH+evOFyUUVV
7XUhsCc69RudH1/8ZAaUmLw4wk0Cod2HFcNWzxUyy222nZgXjmoEPtCQQ2JYXE4p
nqry87j+z50RqHuHveW6PSS4i3J5GvXO0ke5GkIj0R66ZUsri9pXp8OWs14z+N2y
Dks44yYm8kdeJ0Neg6pF+X3IewaUhuCdBZrjE6UBrEo0zk4iX3+QaB6/W7o74nMU
l8N54dHcB+BNU2uqrSnubeyGfdFLW5IrFtZ4qA1eXTT4z/ARD5drItsu9SDhuQfT
YDSbiaam6f70lpzUhdOj7kqBfn8c4DcXxuConWQFhRMNhUjLhtSLdUQVg+RmTg30
WlqC4yaCrTnUmhzKvAoPcL+yxINwf16PFBL5bJIa6cW2GmImPB9m/YLl//F9wvwl
G/CSu1emOh3ot/kIHgVQcR7PehmOybxQGidKdvD5OfmXWNEXKi9H5YDRkapyNczO
M/goHN+ABzAlsa5jwth2nCxIVWWwEx07lyR1j1y2Oj0G9Iufs+PHPdq3uMgesqTM
MM8eeN7lDSlM+CV4ny69O7n+yvpv5YUNDdpqfCVAz0zjYppJ6Ol+gyzBTTSxr8Rm
ESt3gbSK19n8ob8u5moHshGiZhrgOaVCQHiIuVEdiSVhOG4dvHPbrNfYau6V0ErS
oA0z3aDBSGM8qSKhCSgz2GkEZrMINwLYADquVnyRBWHPtBIZQjzIrXsfL7vQu7DI
MDSOO4NcNx1hGTNlPS7gYlK1yTg7T/mjbzX1agmNi5MuOgvQyCEvikIyBEF4J2QC
gQTO5uh3QANCZ7umyD6m0slvO5rQwf4I6HdMea2g1sV0dVIZRrw3YxW3vL8lM5uZ
fu3pReGEI6WZn2ullSZDkjaW6dJH+kRRS0XpyVmB0ojjLVWpeHpBwOEkzsHPC1RX
ujdrJUpbXdcnr0DOnYpQrfQTHT+eyz8uRn/kO6YkMQ7VIRAbrkvZ7aNtSNOsr0ZW
NxAzGRE+lo0SyzhW3jIOi22Sx0GlU+iH07gU0zrATD/FZXsBlc1OZ0uRxiTrtBd+
sbW0FlWveWUd3FUA6d2IffS2Vg9b3+k7Mv79IBa5n4g+aDNbIVJP50AbSYMPkMW5
F33I9pA1UYQU0/+F1G0Nul1XQiLaZP6LQpEO2ERlMzxCbA2u/ujjTzFA/3M7il6M
IltEyd0PPxe+V9M7+7Tg2pZEOC8nev0JqbDtzTNb/sgOvPboUN9UcaecCcsh2Msz
EPlkzarfKi0vFuE/KTZL75aVE4xQnfcWSuDqIAenEGvNHpOf1XDaovB1rpDo666e
eO0UwhXImgSFhJdQRrK/XFXhqIr5XdzXr3kVNC0Ku36Eo2kPMIYO1jOAKRjwSx1M
xkyk+b5eeFzeoG4SgeJDicx6bRiltrzX86Iy87rMc/oKFJKlgzExQlLJOPUwF3Md
I1vX85JVuTUhU3qxWL5zdnEECamViJdir7xbjhp54z6BgmjGp5ToQTG/Uzbt/FHZ
GOnRK0u6h6ogFPrTk20+wCgjsQdPnEuYOxEpjt89VkPfu5Uca5++9DLnlvTXc+Tw
RUuUOOIioa7tOiy7BmMlDxZaZ3Mlm6gU9dJ9tOrPl+MIANGePWoK829+oMNmUHTL
O/ps8d7BcImsrIAyRYDzlUuoSW3J9pB9l72uBRe56GqGL36DEhwD9I+KAUy3/E7Y
pgq44ngoVVXZiOLLRRAvud7klCta4xU8ko4Vjd7vCb/jJ5eKCy6rQtwmNOrd0Kkz
7mo5qrrXNpxYYcjzl+cHVbqMqhIx633FKvn87oEQbGUVSFGRQrm2X0eiuVHFzcJV
4znaHfUhbT2rwBKwYZTloADlkXm60pV79McqTu9eqcJABERT01eLrctLSQzqHICK
aY0ok3QadIc2YE6Cm/z0G5toqBRNCO+yrkK+qy+ws2GF/rDh2dn4X7xgNLc9/v+N
LhvPKEuW35tiG+vHRSdiPHKK0HU1e1KQXk/M6x6biadc9wO5s/U3/xeZuoYvQDzu
s9qo9qwsy2q9+LT9LVf4xcX/P+ijMCxqYVJ63u3wq4kXwJvRKjirxPOyduKS/mID
W8K0wAppo4n+zFT3Et6R3Q1U9VennleMoYkOckVwCEKaZS4d49T8s6JMDLjKK7a6
rwo1v2XoQ8l28X3arfJYQJz9WeuM+l/Phe8qOHTVfDVqx6ZqfxEDqe35OXfUIrkl
2HtPV8Z4yBj8gmG2YIsTqTYo6FBTV9f/kj3ROg4mDdKfPk+ZY8Qr7ZNdsbgHU+ze
D5Eqf6jTNPxOuHYaZE5CzfPY/gFSm4o8D/lsqJV2gixrbAx8E4NZCS7+Y5QmiOdW
MHgxQNwY5bsfcScbFslnUZVaiWiT0ZD8KkdKl4Hplf9OiBcX5EtPpRay8xs/CJEZ
R0FskNAQVxsISksf7Nqic/qdFb+05wFI3AlCrsW5gwjXuHxLkyzj0jjk8ipOtzaK
5+jsetrlrV7NMYRovy4myrOZCa+LMOpiJqdw2+1aXSimz/Sx2u5yMPMthIZVB3R7
a6xONSO03OWY1ddJGm42athZ1urgRESCx43obvMhZgqw5SAZlkDXufn57qH4nuGL
2oVFQgZLonV+z7sWthNP+LOg25DAD2h+uSAMvmNQFmd2zqURxD8FrIlHurRsYTvL
KIQpbeA16wmIwLA1a3qSsNcyP3mqrqZT3+98VXO4ZrXXQHoD6yALLI3iEpr22stf
5k2opE/yDaDMnO1DjNcQbE+if6uxS0L3lPXf+bLKX4ZfOVeSPnQBLzRvLDKNtIBz
//nWco5OdDuGR9Nq+J1KejGqEc4ejp+4m/+rOvJWzf31QIcP4E9VLOZPbQHA5CO8
6Zd9kktfE7oE/+Bp0laMFicRkYndWA8CmqmTX8TYSKIuPKKMiZbqOJmTMiBPkx1/
ANB9hXJZMNhBUYePvLjMKED/4PTqR4sicQqsKxjQppptEYbgsn213ZhXDOe1G269
04eV76VE9L/t5kxpWHlva7anVp2YKCisaB8FulJiN1QuF/ePL0c6Dvx075WqL/Bv
AkZ13r1JRolx9pBHyO3UiHNWq7cZWK+p3IE+qX1sRoUFzkA2Hiajziqk/xy98FVx
V0ZVspC2QyBzFtXzVYZzYIX7Wd83U3eTFwB09PDKS/qLFpLWcSu706xaX7MtTDfD
8nT45v1mspUQwfCYNy2r4CFC5rxiXbu+2U1JsnHlWaqofgY+CS0bZziDo/MdO41M
Vo6E+wxYfSSoXxRdPMwp1ijAlCFUwM2mmEmqiUJMMrRlYZP/x0aYaQzs8MRrhngs
oIvW1he+xvDSQNiJW8vXsL5zzoquYy8eykDo+FOEEKhnOQn/anOPugMqTLKinZIp
uy1Mxc7cW2wrMlILp2EBFOm9lgRTV0xL2BymkoQjk7XuGfHldoR16pmXJdCSb8sD
qdHTtDGS1O1QW6VxNh7BT4O3laFt89Ak60v5Iat60k7jjgoDZE+GSwIzpeUi2URy
ccADFu0EPwq7kI6X5RYFoz1WkiMYipKywc58kFM7P0CDk8CKouMxgcB80MxCoH9L
edhGXPJhm8ADAyda7WXzzBUp9mpHM9SKDRvsewa7P7JqTCckJnOEW7gkxlk000gS
1i3gGlip4kRDVuA8b2XtFusfk7DDjUeF15vK8wglnllxjM2EWuDez+e9YzBwtSlt
aEXVcIfaHKB2uGL1XSw2H9exsQ5C7J3SMZ+MaTBeuwOanx2mZA1LObybq443sB4r
S15hAI6gyGLq8hQ6gohftFC1hwjxAd9E9gVZLZ3b1QeyKOoV/6ex24Pt2+Z5L7RO
WR2Jerz6FmPHKqN3VuhxNOithQl7en89H1/nvh5hhswL1Baw/uXenaXpGpfKnYG0
rvvrSY0JBruz+IqoD5KTYEIu3vlH81LKo3M6ixzMjrGqOOIrUq4hW/r7R1mVRySO
Zsu8rrL5j3uoaOkAQpK9IWcDrG1bZ1gGPpBeTnLU0tJjc+/FLf88RcuTQ51nd13t
2DqyBtdGO1XsQXuUS68UoUC7goZ0c1wTtNIBgHzmV3pbtm3A9pZeHgXlNlOal9rW
KBaTqFLHOAvt+XSW9ypC+nAMADBHv8lc7qCtQZVfv5elYRTzr7+JTPJ6XwmqZI0m
ucz5sClJTz94LohR9DYX3rFzzss0WAEmo/akUCVmGSH7duNIMn1Quslh/h6mEKhp
wUMubKJbKw9JVwaXFoxi23JoRievzCQjHjZiH2vtFuWBRdz+SjLDiPUiWeuo+Gtu
jXcfeey2vSoAjwSw4JoiH/uM9Rw6eSlUUoVa6wRfBJhOiMdH6azSVGzRT6Bi3sNk
HDnidzte6g/cctoCVVzUmeFUROvL67GkdPxa4mbS6zFcPwifPfL+ERAZgRplKL7X
pGPQ8KFS5q34y71PEq+Ml6xDL3ZA6fw0VT6wH7x3HW+PWeMRDF24Cs25KVg+WyWw
LvIf67vpvAkmXTkuRzxov9LQtwI/gF0Mkw7OZxVvTgYtP3Oi/5ct/RcuGO7o8PKp
FW9U1oFZovtd4dqTKHuy2m7P1sZritbNWFltggiJjbk1JmN5fo1yrw8Xs6Kcf26P
lYq1G1Q5NoWaaFhYzLVw3MhBPQ+GAMaRupy0LmUTee2z04Y4c8l5cmUg4DwukDgF
3Upi9zWe0qjpyWcfcKjZGhofc6DzeSz/y54hEkp0BRM3m8XjPnpqDL7FS4aIcV00
v7sIgeu+e6t+ylNyy3B6m7dqXqFmeTQqWVzYKlcALx62g/sjQXME0q41tVfERVLq
YdclOLXzKsnOC88J4ebxPneMEbKR/6um3crqDMOvUl3nZpEMFfOY0n40fDyKe7zw
4pO82Yua6ncggKmMHD/VO8KoA/RcYLi/x+EsDe7dKvN4xyS2OmGxjnjixQeqfjen
OG4MVWCs7uhbtv+CfAWFxQaYq09AygMzJcwcSFPNAySaylPlv9A6Onab8SNap80/
svosrcRPXMIDsU/Qv+l1MGfUepasOKjC04xZ0vFllY85unxPZ3YJ1uul6qPvnQqJ
3ybn7E0ts2oRcuqf3Nj/k+RWUydANPBHJPLqcJwm35/YwrcyQLdOEG8ZGU7XDVKy
4aPnX3c3GgOgRIa6qQIJ+jet/qHvc90GllHnuVXiWyJGqX0XgtwtXtOjnF3Xm0qd
gAZgStaXwRQWMCG9fYNbzcisVH5i+0MMJUp9vFN7os/EWOqSlUNMgBcdtippLQvS
kSh6+AbSaa9fbZT/qyA5Lon7PhLTQ/D62B1ojGcFpa88wmvUGgqqyLMH33VRlvdg
KN5CB6BJGy9C2Zx7/ilaRnz40xyGIHuG0JZMNiUk4plQLs3dYr9nr1ikToCJNuux
yu9HpEx6rTl/R0+4/XEGh+My89TF2E6umdiAOui4egzqA72KlQ7Ja993SQ3Pmpcf
D66T07gdumm29P/EzZQvolV646LuUUIJIXYlTq5u4jXhtLLE4ZisemcaNgemYMfr
3QUDbTXrHwlwfj7/j1669zh9pr79BaBK9VRUXKArDQ/AqYdWcsnBe78ahFiNOQbv
wGVP3GwU7JIeSVHuM0935A0VxDs6Q2Vl3xgQarR74RruYf75UJcMmTFUVzvIZAXr
4zaNv0Gc61rmIuvTgtQ2Ve/UXwbTjxX8duGPlvDPgP+JXpiayiB3Tztsgc5rjnw9
bEcMwdnxN2Gk9JWpkPyKrvldu0fsK9mVLKnCWj+lNLdbwHLl46FCROUbrbhT5hq+
9GLd9dNv4hlfjuAbtD7xDeoD5ItjWmy9MZ1aIQ4p+d9ljGyT5Oxu3WUkeOpbeqi5
IyvpG6TkMvUf/bqY6TjuylZsYnvdqvEDc5ViGukwtbqrz+3yG4Nwwv4qBozIaPyd
Y+/11XuovNtktqYlHDLYj9bOn8M1mM0QnWiJLaXHm96Q1FWv3h5eTgYPrqZN7c4V
+U7/h49k8bSTxD5aQgK7wt+jiUdw7LHqmKI4Jta1vcA9VTnhnyuMHpLC5HH04CWR
XE9KZ+G3hMRn+e+xBse9HjX93OLya7b8pIo4LQwyRcblTAevCjiKoL7gM0/aXFfi
i0hPaWyyLcXIiuW0ZSoq8QqOSCE45nr9tEGkW05f0/8Qf89Bc+W1t2PrPcOBMnbA
04jrHctmg0LODxd7+7RnYjNx4QLY38tUvOY/9uB6SUCgeHbRE/PGwP0BJjyBwQZe
xEJGetnrtFaKKTjaOET38aniW+VzXKRxCA4ljT8HMjtiw9s0IAaouPAr1up5yUOb
9jLFpZShHh5zgZZFsGsDnBch73JSdm0AbmtlnVP9xESwQEqNdFXYGH7cRqdErU2b
cf84pFERQ+/n9wVwyJnVgGZCUki7JPyfQR0P2T8I+b3hVD3GLMHblroYca61a6Hs
eF1Ntuk/xgldLVKpYh6u4bFXsxlVj/ltaZ/QHgy+nDBpaoDWtc8SqNchL70427wm
RBxK8DgE5OAbYMPt8n3iJukxvMIx9MmnrziVlg4EwiV2PjbY5BFOtd0xC/+1pzk0
+POztQ8O9ky0h8sLNwJN2nogTmj8vky34TX+YZxguXg4oeI7fEP0g6dzflrSsAMI
cN2UDRaQyoOWmZlITUgJzIB0YeZa1jlpTc2+bNOGIhJNUXkhSG44Ly25MLabYGM2
L2ODx5LjC6r2Xz4a44u5yzphb/6dDjoK6vdU+d2Ds89C/HJ24VkPbkQ2ylBDwQJd
Y1XHkqK7BcnElC3KTygbGvnk0hGnJso1XqRJAheVlJdill7cTYvxWdwSUoGcmlvH
yxO9ngucLwpGQJ2leU1aalahzH81N3HRf6TlAi7BdhNqv2UueMVB1mdB1fkyARe3
k8/DLIIjbtZKZDNP5sGaJIxIwMqF/iDlY0oz/qLeqLbK7YFtu0PxAm3rqx8gcWu1
6SnJOPDBaJMNZahEzjslcYtQi4vqURuK8A+AjQbNxqXrHMSmZaM8pvk552eiyFxL
bYKe22z4AvH24/M5Uv5M4F9O2Rt+0UEKgonDV58B8w2H7oCdNqsbjjARAEl50eDp
zb6nlYWIc9Y4sDjWNGyx5DWHuynD8qmyosZC0xr8lmO3VLYEptl/T1UOsMOT61Dr
HFwduqZIFn88U9yKtrrV+WJ52vbT+c6LwpTPsjDyoNiaFH7m77LWCuPbOXoR+MXF
10VU3TG+AOVpmoGwaUgSU3Bl9g0u3OtqcCJPXaT+FQXzoVaU6yzDkr3bnnamBNRJ
GvPQkS1ib1Ctioj9KIBB/FS5d6Vgr6wwSV0pAzgb5u50IMgtiNwlh/whQplT76BM
ZWyDSHXp4/5O6PPgvVOVJHLSP+wdEGO7v2gcBaxEA3mrh2RysnibxPATrVpAbFQp
nNf7ThNgXEvbDxyUKDACoa5PTHo3BWzjN4HTaBUBhaklkVd3rURUNOmLczze6AxQ
tiH/qz16W7s/uW9hgvdyGJciCfVhyLSdV/h5+TLm5qH9YeQjtCBk3da3Vm8ZrGxX
0xDnmh3PhGe8V0LjhFGb3tIt3TvMlU8An8T17hiUJP6QkV6Kl3/srgY/LsIsmFkX
Zh8aMzaLJXIVnvzCS4SJrDRfrZtxO+4N2CBL2m/VkqsYiOY+gqXkihgxPQU8ZIlY
EPGMBPt0n3uCwRh5+ufaCDoZIbE3vIkUH3MRx+SNBfpGNFvO0YKUY8kOmuL3U/ly
g/DS5LWXj4qOc3Ehq4jXR8YhdGlBZvalF3S6lc2/jJpl80aefMMU6arHuhUbt+CB
jx4fsA0Zh1pQ7comG9hGd4q+sarImMrLL78bKQDuJ+LMwHPC3R7h5tFiEyJcufYa
Xb9Bvj5GL2lg4UvHJM5vC6x8ymBNQPSYVO+JH3LW1F/ra9SNlxiWhqWG1kKQE42b
nBMnlIK18T5hbViKlmK/8Yj1hCgkB/KZMTkTZ3/NX84vmPsPNxZflCyp+jYVbYDb
kFnN85XaYqJt1OtZq/Lhh2epoxjhXbC4QrNUMFl59o3D1czep+V/jXN5a+3LFN2B
AadLmMhbRUW20ivYW0qce8Em3uaeHuIR3tP5yS0nst4zQY+uMdZGfTZTcVgrt/9W
DwUvk9Zw6mMiXU7rzr5IZJ3YTVWUCwq0+1An16wPduP3CmTWy+koglkfN+xdDaIB
hlpv6I3vPShSMys7Nu6YGxDkHzBN3eG1qwdWN6sodl/lDR4ZlCmYicK0JGpB3C5D
1wE20z0eiSMp02mfKIDqHcDrbvPliawGEbQWyjRbOtg5NFgbd8wEewJkoVEsBkm9
GaISaSY36at39CIcAA97l8PdIHiAep3QsQNy2n8jsHCIby5k8PgDr1SuOGydWPlf
jOMJrPeuQzWu1ICIw6aLy0l4WxbmtsOtTAXegmXCf6zd/aAF07BBcdxMv2tHVIvp
agmUi0krz1sx4zYhlPd0hqhAZKEAmwCI8xNDHLcAT5NG24Wwfa3TyzVrThy95saf
mrmS3tvPBOBIxUcxFqeXg27oSnr/3e343pI6AtxT3gDVA/yGUUkokDcwgEMIfxTQ
jXAx3H5a+QOgM1mBvnQDGM4XzDel/Xbz4TBJ4dgZi7R31FKUthrHiNO2DmotwfH+
VG7bYa+ikcpBE1JTxKUylxii4cogeBL31BYmSKltMlz3rK7bqsBHx76O+Z9aYvMz
WYHZC6o7zDBtrOxwwzwHKA8UIkd0UWW3W8lPLBEOPCg3ArWRrEHSm0q/q+i2Ws4O
SHQsfQkwiDEkBmxCvMb8LarzwfDZubNwPpQQyUjSjzF4uuwWzyb15OP+5dwvG3sr
48LEaWIvWnOJxYhqSchCtv8OW+isp7LTqbUEUD1KfheYIIfxFbLgYRWByp4We6BM
BgFKDYAihrJ7S0xe3VgeLtu+eleSg6mEYyP2XiGCePAV3N+Nvrepx5lT/vTwCUsO
Mo3t02Fsl6oM1JSM5qBCgUcpu1D4DXQrlYslgBaazj3q11iv7/MD4louBgKKSqow
PPhBVNckjYYhNq+UirFWvD49QExCXMUyBLrysb6OG1d6H8Vq7OVvPMucoFb2I5QA
YDgpkwZsSfZRqj92GEFxo81AfxkkVIHdV7sALV5iZvpb54jzkecDFZ5rUI62a+1B
cb8cQ9XIJ/E1g2tKZoRSRq9Dlj0Qs270Z7UMUiSlrHXvYEUfjX4iO+/txphBKs5G
w/V+IwuMb4776Qys8mWZ5cfgIF1kLSSBdIggfRxIJJQQ2wNAEbaYjqCOT2CA9meV
6NVLVoD3dDgTpWjpMfGDjZ6k+f/zxG+twHFAlEbkC/1Q5oMEZMp97TSCK1dihj92
SAxJ06jCqSMCuGxyvjrxz3MFKjatfzeyGLhVyXTx5L6p6wqQMrkTA+NUgEBQ0Sqx
181/V0NTnDdsi4XwmTD0ccYxw2oWqq29gPfYoeu/yIguEH5HZ7H1yweQt/34Ls5K
2KpwkvUm5jCRZ8iWptwyo58esey4nS8VwQ9TYv4RhbF7TMAYYFHqV25jqjiXrRr/
sE5bDn2KcQwQCkUsOI8lxH9S8UItZ1DilfSGr+VOKv7G9N3v6NmhVISXnl6b+jfs
X/MZMxNOSvrGe5kF3bQf2ZnFD68FXgG2M2RL9oo3szjH6Fz31l8OpQPF3n+bi6M8
mFZfAW5odls8UhNKf19sgeq5brX+8Bp/4gkrh11s6jvQm7ogYL8S7vE8WdH5BPun
jPo+O7DIWRCKta3DEMvnR0ID35BzKdiqRoVYG7peWNXtAU/zsY9e1779X4Q6djFX
woLfSFmyWicwIoS1di1jAvpKzkftaY4bGG2U9tfYb4S6Z9xnvvmzX+JY5JQ6jf/Z
REYeY6dnJJe6tfS6Auh28Rvs/IDqBBPT7OKXP5QqjeBne8qzMyKtCyKABDWXPbST
a9Cb6WH7L93rviMahm68YnjjNgTcFIMNybRWD5LVOaBogzU1Dk+43x83DXZh6esJ
OQ/FbvrpWKH/pC9gX4WPrvsZdA+OSgiOpAuVALewWqM0Yw//IMz6aVS575xMF/1x
W+AkjIckr7r3ZafGPMx1fksqfQZxcHfa0JP7VJAcyls6xH60SG2TWtopW5HgQyGt
a8cAifVLedpTzNp1DAcC1Hl64JjzQ1MNfiytmlkcEOjIp0neR4bYRn5rqPp08R+3
Nyv+tVL8Kf6wbnjzAwqHvZJlEAxmNJtzGLDmBIoxXMtM+jPsLVNiCO9f/P5bnocw
XsrrXSSouA1vTZfk2q8CJi0xkt2p+mNo54NtvyGxVOKQMTRbBX01B0vLwGVIOaOF
DKbQoc9GNPg8H14pBnXEkwRFHW5yY67O3D+c9fKiXgSWF3a0ca1Al0gv7KbPXkzJ
s44IsnRX8SKRf5oHZZdLG81EqZrUFnlq3a1o3C6/l0zXypwUh6CfanJn7I6giJ+S
/85Om4epCReGDDc0KH8lbRdDp8wijDbMKPr9pqvPh6IZGyF7GDi6YU+5NCWggnSC
2KlvFwwfqW7+C3DbMlgsZZrL9mhhiP/nv2eflZG6B5dsqrEQ5jnRKK69so3x1ZNJ
jgDUoCvDoMyabUyOD2fs97OnsAxO/dZnZFhjl8/rCTYDAt3Cqruey/DK6JQrrBGq
hMk/eIOy7rkxUFzBUtJcnOav6QzPBW5CChl9zQWA5nhX5D9ajMXNkbrdFX0rUVtM
FJ2oHM2bxCsq65g5yM0O7x5azCAkJqkvBMoWqO4tNXKN8UFEQRM/Db0dmFZChleO
RrkMAS1RWdvMbQoJVQboVsR43bYYyfgpiQ3CdNCi8czC20zzqOZTfB8PKBaygFeQ
prRhfDnWH7sWCEm1Ae/l899W8W94CkHljI092BsudXNOlnY3x615xIHDiaVtSf5m
VRIzQVVsJqN14DunKMUqB81NpkqqMwli43P1D9jd/Ue01s+vT+/uDrYvMeMtijtC
xqcoWGPQDz9Ca5c7Mp+nq/CXbHQyIG13Wz4P3mFIDCC32yDJwlJ5+UToMr4kyZGq
U612U4C1hdc5ddbEF4OpSkKLH3Bdnfel/zjZXAhDUGdAxPVPVTyLHrmotdwLABcA
zVVHdKvnckbDk65PRtLcLK32MmIDfa7OZsjjSRewgZnP8vsh7DFvMWjKT59kQSUK
QE1z8sldUpRDMM3kuKJqCcmgcrGOfRA0YNQ3af6wuQA98emI0oE8cFCGJIEHvmbE
q1yNU56hvmmE+sgq2RmidO3ag78aH0W1EltOhSXyTXZrFLI87olS4dPemQNMu/w2
oInZ8Xab1C2qrjatHdxbK7C8qA9rTtRLSDBOOC3fxOmId7aaNyj5SqD4vKaXJs3J
541Ir7IGQxNledwRZf6fUTWUSyC4NmhsdeMnLKx+4SChnbGBA95ohfpDNAGnQJkT
UHBMDNLVxswb8GegWRJhPEdmRlhcsDG2jtPIrLNr2sHeB3tVNyEuvlMxFEMjaHD4
sENUc4/TXrPeTX5ff2fLzLM35pkZwwDki1YYZASVmqeKe2P6h9oU2IxGskmE+Xsi
+KRt3TUHcVnnobEaApSI4LK2OAoOBDRG0tKShP1hRmdTWIZ4/5dZGkKuGl79D4Mf
aJvaKne7tFtuIQSbEF9nHrhuVw8mWvsrkaIwHdCS8Qg+NdItLuytCICfNS1El0nl
RuOc4gowp2iCCjcWX4A+1A5hG6lFZ0wc1EksjRlliv6brw0kPexTHBoaOJObB+IU
ggVIP9Mw6Iu/e12ZxasrtswoQ6jql4RgpFZSq9byZ0dOAFPgZTVAvtgwJ3xG1QbL
M06tt+R+oA9KWNSInZsim7WB2Cf+shyTI4rLMirrHnFbYHash33hRW6hqJAXHqSR
b+IDyMz4Bl2+336W40s2/xkX6GiiryHhhIPBgnjFAuyo5yjkRvl6mOiLrdSuSlYJ
tboMNuYP7VnC/v+hZjz2UNwpZ4DjUN8WR16C1cdjqv2RXp9i0mshAQJCU0NGnwse
6na0BZoFkUqlLn8N35FPI6s9SENaHBA2k2XmtoVCs3Qy2kbAAStmCJ9PvjvkpCxi
G1oWfQpN+cntu0ivlu849XrjMGk3Lyr9zcYCU8271760J0nH4lrsEC4Xt86eqORE
yaf4qIe9D6LDygIlHDE7FmRdMfNmhaGhT5rxXWkcaNgPQgB6P3a0KGl0MHEvf+pa
GHlZ8sUO2HUlLHBC9hEi611bgYJKBLhqxM7IbeL6+fEPkWRA6oHlzNcNb1UdC962
KIT49OGKclz4t4EeAHfbfzLoeF8o4TxjFjbN/xb+6NFIPRwdl9TU/XC9/U8To4Pm
g0PjItXH7Hp7OCLfVyplwzlhMuMVByMR1goBallic9jhvAYdUch3R4OBV0gmJ/Z2
1hP/iE+R8pA/3biJG9iMe6D82LcllMeuEDv7xloOEk91ey5nNPe877pEBedHB7vs
lBK13vYQvwAAS43Doi2LXQfhR7JAE5aFrr6baZhXnQ2v5awtidmrCkIrXH4Yt4BX
7oUtvAEThXBw1aVsWNoy2GHDwXQvLu8JN7Bj280EtOyr4u7M5/yafXpakysPrI+c
8y7ruH2rgzRkpBbaJh845kslJvHuN/G6iUdKxAjmAkJ5E7FjDq6Xx4v/P8Xu30r4
f3C2hLImEK2v4PJ9Bj7hJPvVVJpXDPB7JEBVUdEngt9qBDuWsX10zT0wjA5eoaYo
uPEkH8plIQm6s01tQR+tJ9O3YTZnoUkhI3ZfECJroK4JxdCvJPLoli/I4SbYUJjV
dFbJqngeRH0V+n0F7uPnlj8y8PBvYwqhDUwLrTmtSwrJ4DwIIIqT4uxUa0+MyXbh
ck18q2dukxseqZMeupIU2bBlUYlGxPsPQMC+FNPk881dxPlEbm6pvEyHL0a1kk93
ZuTBYJV9EUVzmLIB0bC+NPeolEnzJdcZwzoUZKhd/y9UsLobzulUIW9sZbgFj9XC
ky/TYmOKjtwl7ju/Q2TTMO4L65gfdvND/e5Vf5cKcK2+FGnAx/rFJnq2s45JDQ3z
5x9o1QW7OLcjfBkPpcCU4b5KGA4ZkuSsrMiC+a6Bz7CHoPGcnDpolq69VTf0epMi
qkI4DZ6wXlFwx7KcOVz68rNZVdrhKu+nvThsrBwxtPVdYKvPWDxgyKKYw+x05ox5
/7Aikz2hRqiVaGcp24nXgZC3vqHJ9T56AUK95RLjkVanxGEdWs6XHbvtXF2Kq0HA
mCnbO+962dr5O6ypQM6ziGUkzCeyfjJArilLu2alSdaYyq3qwebpzGw1623rOE98
OIg6O3Q/z9/uUSG0OOMT0FxehcKsrhUm2IozE60O9YFg+G85Om0r15y26xhlO16I
RmSoufGG4uqXWnlWSKWOzz52JketzOo05m0II3gAcr8gSV2RmwiZV6b1no9KktIm
2CcgOxiMp0LVV1I8LuX5ozFP+ZLfdTVeJpZNJCOriP5DRqWOXc+gg/9kQmf4VMvR
7e2Yn4y5N3xZ/YO2Tzl/2X3zLa4CPR8najMZzRnILSVajCkFxGjoE5s4jHwG5ypG
s8DyEX13BhL246wZlF1Q/WzBGuIbeL2p2+aF3a0JA8IhwdiiosHYJuFqmDhLlMF0
xnRo2nUGJJc2DIeHd98qWICmFLSMGPzMJJtQpZUoAqyUpnnCYN8ppm65WYDOI8aX
HsTJNLdjYs7QWDCgNBOmYdJd9PXQxCa/iaanL0j0VFfMnPVjrY020i6gDeOmED7i
PXjhNr33bRF7m5Kjr2kPb4k0BIdQytYfnHNbZfzM9lrq/MjMXI3AWJYd+ExWOc5i
iw5Tn6gAPSMagsBFzr0+GcQdxJIMPphlR6aC8YLXdYJ+apwn8GTkoC1qvAPWZWls
QWhTbJXxwVH94S/pVD7bCm1S7HAzESIL2PgjhZMpB9vaQteFyiYi9OcLT85gEmS/
NhuEB1gJm/ny/S/JTBXbEsQrgukjSG0BIZHi5cIkIs7Kvv3GZyiKG4rhqqSCS3oB
/iSn0Oh2lgEeH7KVW3TDILpXWz0pzMz8k97NfSYzRY1Q6o7UCROdEaM9qqYQ413M
e27xI/0pnLR9yiPMlyAwM2ljkb3bZXj3D1JRQad6uHtUMVjwlkdQTjoKr64CESSy
cU9nZKSupuzl+eHk2+QAU60E2aoYKMz5oy0JzKtRdJwEH/nQEqVJmetwuKAel1E7
hvgGJja+yEWVmpTJNpVAo4eUiuZzlEDpLbUimUH/Pu1Rg7SQHCG/DgvA1516X90x
6Ge6acbbVzcJsW4b1bKOWUye5f2PPv9r6iVEOJXJMUxeYNoRyVSkhla+aTM5wZ4P
U2cyX5DZTEErC7pgbP2gMkuy02Di7K7duaR/V7YECAYt0FDgV7Ibb2J1xgfQ0i1X
TLGpWxFcfIWvfIQy6MgIqxjOALXRG8eUGgCkySOIgjpDqOjwFkxK1NVjdAzm9OP4
s8V8TnZ51W4RreFw3tM9HrOrVrSvrbAkQQsTSG6/p7sjBCCXsZnjyib/VqiL6y4t
jtTJHsmCq0tKfmkVXifeKz+Yu4UDKHeHHynyvfc03TCoM/+WqLA0hT7sTCLjLuBC
yyijdDfxI3EiofZVJ2xAj3fOjzxUB+9kvkHwgC8+EvTubPunNhY6CFBtLd/NOZyp
aShd+R3FdVy+eE/CxZFY8lJfGgdiUxZEaVsTrlrURKZmiwC8cvbEnVKCh1jl21y5
Mmbq6QURNOr8m4Ukeb5Ovkaw8QuK68LN/kWzMIhihkuqN/N9pRJ/g6NZxtICh+Z3
odkziY3CLKwJKgtSwRy9KNJUmvaWcKTtH5mQv3OoB/hMS4ntIhH1CRYWwl9RcQ44
HEuCfkK13Edo19UznkOM4oNoF2nvykzMgq7ghX3Zk1099wsbl6wRe5ydRDfOt01M
JpzL9sxjTL15PofrmcAFaEehU9XqTKQLo+JZrerH01gkN1Dc+0/6OqNr2Ac3IxMm
RVSszbxFx8IZXrw7++uSbnGuMJ256IOv4t8DG/zg8HpPSuNCtRERefxMhdZZ6KJK
FRFyh7FlDp0TObaKd2yZJpzM5pqv6vmFikhrCrt5rkjv5hzL+++JB5EQXZi6zUCT
rgnAgLEfhN5NQIzK2Y74o3EFmF+JROqhESZh4a6A+qypHUgY1fqRoRC3nW492jdR
+GEcJ+RyUWU+60WUCZ+/cjMoRf1zZ4Slcee7Tu8YTjpw+RQsLCIc9eD4PSwHqe4W
vrcH33bnxcLhe/wvISO4E6+dOAYOCiBXyqhc7Y8Og58bywyK4KwqXuR70GXd5gqz
1IVpgHztCpcI+OLlKfRZfv0kJ/+DgikPOayYIjB2e9u60h8tBIbq7ZMEu9xvKTwN
+aVCK757j1bDdjmJ+KjnclRiLK530DcsfXonWxopXm8zmnr2K1mkfZ/Q4r9WdLYa
pRR7SL9Yn1Q8vluGES9gLUQkdo2mxobow5W+QU8J0ZnwCrlFTtGuqYyT2bxQuIXc
MpQdCXosKQ4ccs9Ow7RzQwQ9WexJefYjL9JmSxcl2pIn9ioCxItxznhWMryCy+Q0
QCDPtk0/xtu1m9GoaKC079G5FBRcZQdJbBC7yxxqSaVt/1AJXcXiyOKd0pczYbcf
jmitf/PkGFHZfA8tdwSEd/IxN6q3O7+Zu7YSSQmWR/oB5CIbZqAq47JkV3krAVUW
IoFqxQRO/Hn24Q8pKDeF/YwnGkpQJ5BY241WFnBzRjjOJ5k6mlVxpXZP5yE7DtWl
W4UC9F6/GzGJLQW6IKBIR7mhnhjmvn4KFEZlvwKOuX43h9JjfIUM4f85Vrsuz9SG
vtlbmnIIAVf1O/tA/QjFMmYAa+Jrjbd6Xd0LcgeRdnMC7CI3WEf6tGPtXC/YDp4b
vdW/XeZwqb5/W3VrU2Ey7ayWgl669TqqiDscowLwa0N01vbvPtW1A5iZ9YvBmw4r
36EhKY2BvdIoClgF7/CKFy5XDuBO+ibUetXJsIkknYHtKOLhxnbWcQJ+Gm14M8+s
o/t3C1ySHVC4NufLwg3wFH0t0AQlUZO9lDjgOEq7o6/641vaiC6BPAEZ8lyL9C+6
m1i+3xx4QlNE67GVjTrWknJK+lHfQmE6rYKjusAnjiREPshZcTloMRNypOqQcNNc
PouoKAB1PStdTFo/PFlv6Grz856aeWwO3p/11zClyl9OWWi4smLDVKnBXTlgAT0k
bD2wZyfP638IVdHJ3acFHj3PLg5eReveCTXHx04ExiEbhgYuX539KHUPNLF8qqal
GPU/HjxtnbBHODDKos/a1bt3RJOQIqGELBpDgCFe7HWUIoCLXFQkB3myIPnd9PZI
OqKx7vRxV87KpKTpbCUPHWps7hTOII5ybjLO48a/DVU+AxnIX+F8TgLoFtsMAYN1
wj7jr3SQwHmKNlc8YE0MydXprG3H5M/KdNSDAurwizEU/7SjEBokKS7NKa5oKR65
bl4LAydp8+MpLYq7w8fEc7tYPwrnDNygLnColFSRtJqmVkpZTTvuQjzH7NUIlY9T
yP70Al8VnoWQmtEK8AEH58ACQMR3FkIIH7o5jaGMwNlv6HWuTfYu5tBDj46erzpA
yV7RfryWVK41J5txSnZcSjHNUebQRCiPpIlUR3sZ16FMsnFj3oU70fGlvP8sWbep
GuzhKKNmJuMacgRL+CffBCN5muNwlEiE05iWEwKKQe8RjczBIfQsvHcdlk7fg/Zs
0YY7RhaKMjuxkmBea9XO3xKTFbhPSXrG9TNSSbSFrdxK6qCJdkU04cjkMKl8sx4b
x4oHZ/gtWp+lNWtLyoyGvcIrdSbh/4EVehjKsENXpjNlSqd8d964Wygk6nKm94YZ
NliSh6G5etY5pobSW8GGV+AoQR9jUDdmVlD77gBKc3Gm/G+h+qzIPf5AD31l7I52
x5Lau3d5eARGq7OHy9uA4rFyMa6mEspaGglW+kr3OgqvbBoO0cWQzGeKEjO1UoYP
QVOi6gNhvVAviQyx81gQplTkA8BgmwhoLzSpL5h+a1JFugNkjRnGYsxhcXUhCoxy
6CqcL+sPnzhW4lwMpjck0hIkd3OLolUuvdf5WDb0HGECC2Oako4uHnCSQZO0Lf4C
Y8XmqhlBtRPM+6C0OOjWUVSl0NWln3glefkAPEKy5dNt0uL7n37hOvPOqSZYvcI2
UmihFCoikd+x9g5fvg4KR6CLGZN3FXvImileMs1wrK/WRGeDLue42EmjD7MMEu7T
hmZBPVnJnkr5QzMvOpucAffAxWmqW+8SHigJ/ayseCQwMDV4rkg2hSsLiI7aA/Vj
wvCOYhJLhiI/t5nVRdLRFa5DVDwMCUJRdnefLzfba77ethBKZmsZNxUel26HqGeA
YqOZfxQXNNsMMRgOLYqKcrYVskqMMMDWpF/1suMx404hO9K73poZagMzQzr+fT5Z
F2etHmaMjgmW7plRJppi0AXkAS75aOlVyVQEBrHwYjWM3I8PRlBtKix6CtozIcwo
Hb6DquRUrGf5FqZP2vMfUwu2RxW36k5iEIb8/Sy6bAiAccQH0eJec3seuSeZbxzN
EsW/8GyksErgAVIPn3H/hHipEeIpda6maiKAM8B7zQN0zlHEDo2o9vwinL8Qrvzd
Kl3Wa++/8FfX97/oPXhnxn1EvJaFx5FexrKFIfGJfQFKmn/7AzgWJ5TjY5a52zkV
KDEquEwUTmiQKvfhsoKByN/VlxT0vpvtbibSnoPUYqkpLnO4a6vLfWwI04+MijNa
wXeBwwlzIs/DTvXF16leIuvtaUeekEapV5QjtcgyrXByKuznw1LGlS4V6xEZocma
f7+Ss+dWLmVyCjX57W6qF6gZZ1yGHUf5VqzLLU1eGL5Tbvg/Lsfhqn8jV3XiJs1S
Tdm+3TZRjuvnFyHmrYg4kCCHrVjkPpn69Xv4FpbVbS4dNppj+B0DZF2ObW21gj9G
ELP3mjCBSgbTOdwJ/R4c+JxD7By+o21q9xWPPCrWwAScIznaKpuyQvZUsY3hrHKp
3H1Dk/+/rDjk1HzTvN9C+0OP6CN5biVSeoFPQbqKZmIzhDfVLQi9rOl5Nx/htPJ0
b0zr5eX26shvdq+vTFISWhFieA0YPe7tEFX76xqho5GQtvbHg8KgXdZwYs3wYsO2
ruiCGBH7Ph3UjTnUQ9zmZK88+cDMrwrpDq1J6FWZJK/saRApAiQLGPpB98JeGwJ9
oPWtdMYEs3toliCec8ucef2kdRWvxuWoAh/ZKXh7GshusLIEpbSnRk9eiuWwa1pW
3uI3T1MwMVdUDvwKh0xYUjq7nKii5b0yDEJpFUrcydRvNhWhVe6Xrn6ZVp8h0poi
oJh0mcEjvIx+C78zUZ8K3qh/FbRdAZ9Ci3JVENpHGLkBVDo6EAc0Deii5hv+5oJT
dJ5JyNWsQGiM1xU/X5cwvQfTyt8COfQD7DjdG6UPA+E2ibBcpP+JUq4o0EYrYeyS
F4d9Yr/Z+fnzyE0OGHtlOVEHUvMQDGetXACJHFBpZ7wuYt1GF5fgloQgbHDRlO6B
X8Fg7OuY3/01EGCCp1hzMWwF+s4Qi/Bnrfvdzy8eljYoX02IJECxdMKLdhT/raDw
rC8kgcIdzT29ewSyB2vEakIyO9o3WQ2WCEfy+FI1NO/Ml81stgiZAJX8hmHbH0ow
nDD6n/LyEgOXBkE6PjSiU35lqmFDXBDyUTRr0POfWMMzIy6r2ymWlTcGBUnEEMX7
vpcowfTdaYjwZEMcSb9/aRgen2feoqIheJt2jZkDlgdFQLGNG892237V/Ug1ne5X
VLbg/22RExgKhDXPvY2akcd93LpXmZYv/4ZNNk3RQocCIszvKlYcGNj8Cy3YPbMo
kStWZkOxIU4u3oQ+5e8EiFzFjyb9FsC9FLdz31VxB4tFZLhP+TlqFTyVKONu1Cbc
9Kj5Z9Vj0MVpL+kN50hqHDM9CQ4H0KmVXmfdhH6YgKKdS/fuzEt1T8W2LWeAz5qc
jNLWpD2gfrUCbsRgFd9a1i5MCWjvRR+or6o4yMzZe6l5EGSIj4v2xxXO+ecGi75/
RBAkjNpFA5iu4I1R7UDR2OrAhkU7P1GzJ7UtA5H1hW8AYhdZFflVHNdz17Wcv8r5
YPioYn5wBAK/AGjv4tWAbNbO63ylmgQgeseToclJ0BieRpqbZ8Fejna1yjhNeEtB
TwnO9tY7g5zeyXMd6h56vYDtKDhcyNSez9XalJZldzQUreM2qIo0Ibd8UVTXYcgR
naXd3qwFv6ywqv9WOjy1dd2yW/tPsXDv8+CgoXFFkyXVhy+sakXELJwbamONkfj4
JVCA/rK0a4/PwLK291vEzISW3McIEd1tPAsIwqCBgE6vPytNxHvpVnV0AmBULB1s
U0Ljo+RkIG9if0zUIPhOhbPA8YuJAFMdbTfVnCX5l8YXiYBzuvBstCgKXILDIm3Z
T4CWjcDkpFbczlKjsEXPvPUV9/3MzBl0bzrjKwm5GZC51B/ygi7Kt4wkWh/o/Ll7
sFFwGNce8d8A9eqAfE8F/i5z2eC4Otyu845I7QpFOI4XhiDJuuGEeiS5qrB1CQdJ
Kik6HTRmedtUnaCFja2tGb4unE6IINxEEQfJBTj7cwJgI+ERMt+9mJRin98R6tAs
yukngHqugjKUXtG1MXAFOZbbYsoLpDV6PBL0iNjNwOhIFudzB6M6DIT3Wyn9Toej
pgFgtJ8GLKjVXW71wv+FhZ8Z2DTxzzpLFeCt4A7i6UX7wwv5VfEzTMR9TfEFJRIC
kn2YqNmU7IYtNEnN1PTYdOABXjFeymxf+Vo84kVvMrtAwFmXF7Vj79EkzVjgDIHo
qnqmrl+QOa7Ummqib4EpX/tuUzh6SXu4GIlNWfd3nKGq0R4hzfFfurNs6yEAoqN3
NmmATv15EyJT7syssoCFbWsMa81ngVBWefxbk1DzaCswBtXfaCT+6YnUBpkv+AJb
VWc1Gt89kGGtvvZXkRhDNQwV5dC1si4pL546t9OTsPjnVSMo4KoiuN51ihmvIe3p
1C+IetebOGQaYhP1nBiOShOtsgtC6u+9wEvi16CEVBEIhO+tfd+KAL71Ikr8wQbW
DI7OAeRiCOU8rvncB9oolif5eUwc0SCjK3PH1ggxnQDrhNIosufWdQxGVaYGcSsM
YB/sQ+L3SlXRjAHZ7buhsFkv28Fc/bNXBIpNJHH0EwpHCe1fvYxBTGKoEErFSEyh
flQz+ru09/aM33KYIyNoWR/wMLkjJ96vgKtskT0fObQ2FbVsuvZfI7/VbV/K29lD
7KJA5/PIS4JeHY55KamC4ixyjj6lHV/SIiXNpTkI2+WZB3nyT/N9fUjtlueYCDKQ
GrVbJK+X5Ass4GiBDOmQ3iG/CVAZ6IfzARU8MXxmFMzmhOlfvF/iF5SGotOgZBfe
77Ww2DsNvL4IiQC9AGqgt5CN7kWHvQ+FOfyzEt5eldq1OL9mS/VJLC5RAUP6xcZl
20enqzTQhkjnrQmyLQ43d61Hk6qdQrAjeqE/oz4v9xYJHKGlS8PEKu/nzEoqym5c
1gB/wZegs9lenYLYAvJhlYKmaocHZklPSXlHP/7xDSzIMckNLq8ychFzD9+CEi2W
KI7w94Z4QKLWxArFHTy7gxnQPcoZLmNcpuLwrjlNdu8IOY3wTL6iBsYcobH6lnYK
CNOH9Vs9bNvQEd/CzIWV2VACTIYBubAZDqpmij532vz6BOQUJuurEMxT5wgJtIva
InBGglDF6MjoQt380tnCzF3PNt6/bCLjCCa0IXbfpTNjVWHDOfJnDVj6RwHqdBZj
X4ibWu/I4u6E0XF9pxxpEQcKyc+SCEiIyUBBG5wjOWkijBW/f7hAm4s+dGEIKAId
nom5WyUrEdsWaTWXKUP6cc3R7ZGBnHZMzemfnT5sUxv+7DftfLB9qgXVFUdF80b8
ICpil2qr3OmX7Y30tugT36/RdEurJO65k+w4eb4DH+SXMfbehhgba1f77T4b0cR+
CHwipevJzCNnBQs3x2YwRvFLthLjUGXlBLbT8kofmP8e2UPxphg8wpYnZOh2UZOw
LKSkBNTamaSzON/qfwXXVPyQB+/HrtkOezwkhfb0yAj+cq7GqTBz4hQw9TjRvGgE
es4jys+gMhFyU4siLveGgRcnZt2J5Zm2+cYmLIhig/VUMRcbpz9Yh+Emy6Q/3aci
93uRpgn0xmydcXlO46OihNSJ2CSc2glWuTzlW7jpW3xliBpEbZux5XWitQfXWfs5
TROuhW4LyYZcqP1mb0XchUapPAC+jSBmOXvRjNh19MYV+Wa36B8eCudS++Ol+xzP
3FRkGD6Mpy6WFqsg076IcwWrgKqH6JOS2Bpl0td8n1YXvfsm5/PFky254O3Pw/V/
LouAj5Wl7vw3pHb7NGfMofDhjbq8C+/U+xv20ZNO/2ocWV2kXqMggde0EbeHp/lW
8p8BVv4Byp6TC/AvK0BrwIumT73D+u5a/PG9Q0Xph+8M+FeJrBtuh38JV+lNb1M2
A0NrwRdRLVZAimY0CgHnfAx8xYsjyaLIlT/SRB0zvr9VEt7gbx0slhobvK/ZFtHy
xhKJe6jxuWAG8MPAKqlyDL5Ui0SEcDxZS/VfIa8KUIz+f1fnUXnKypMwimyyF2Uq
b4oIDQBXOzxKk58Pi4E6pLY9jGecBPePsTNNEyKeYROKc106H1do3g9U8dMZtNMx
JJ/HF16+RKcvB17fOezqEq64MwuQlCho84dIkbeFwvI/1dTZqQfkzfkPtrHKCUgn
sMBInSVCnyGL9jIMmVD8GahISsSc07L2U5QfX9R9QpyEcc1M2CEZPoz2BOlALjlm
XwYwliRyUTPA3UevnxQhKJ4Pllh1xqya7osDLtwRto0RgCY05fLaEMmOUftLsTkN
yxW7UnvP9IWyPKz2Xxk80qdfVsjjcNQkBaDtD/Djc8KWZlS6fvMfkGz3XPKUBImO
uXRlyAFTRHWIzSi9lfEtH7t7B55Zk6N9Nz3lwZlcgPNzjZt6MPAThI3wphrbr48E
MeQcxh6l8PKAW349W/svZ5fSdS1Waqh6knB/GIiE3LqzSHSSqyQ74SacUpsClPS1
arv+9ZHlO+bTdEyJGI7ZbsVl5UvwyuIXnjFUeMEuIK+U+TxcD8PXlalRjs1J4SJu
TGCfWBh6b//zy+FUkZQZsu+LGrhbM7aYloE76TjRqx23Rqj2R7sLFvp8Q7zsPS88
MoEE2JBY6DPe7tWqUfKev9hoaxay1cq5EB68i+1lo4xw0lC07YBPQ0n30rQidWqI
Dep3kYNmSFKI29oUb60o0mbpFxRaD0LEX9i4zDzL/sRht5Cwxt/G5TliG0zJnekE
XYWQfGOgib62AcnYV6RXh2c0OnS78Yq+sR8XJzASnqHNKO0eDzEu9yZlSiSRGhf3
5tGOMWVoCLF7SjUDgZB5XBg73Zt9mz8bx+P7E3FeqcPdXItbroHnvyTarIuRVCuQ
YRNgSvJMWuWsqqLyO5RC29taLxel2OzBLQXjyMerpr9g81nCoY3hPYCFIGLo/k+S
YXJnBD0YLq0DT651QBHvQybRjJwJZkcpSyPq5dGYHYE/4XUCS4sdSa/e7Le1ICKi
h98xnkOy23SvFEsObNtWu+6SJkxHV+alig4qxMeOKud8ENXkcs66XhEv7zTJMfy7
1oW9qJyVxpNG1zMghRGezKaoC+BMhmcmQBbYYHKsYApxssA/jgYWz9oKq3GsEPdg
GQNzR7GCtFvX60/QoLhS/R2hxWginq1wbEntWe1SFE0uDrOo3k4DaonYbk8bzpT4
r9mtBhzM74q59EDMp/ql5Vh9cZUOxE/gniCJMdAPFLKareCJfUg9C/UQQHvI9X6C
LsQlX3//POeL05aR81sNOeIE0Rhp48Sdh/EVdYnzbR4r3QIgtsBotHLnkcliFKqS
UwBZ1pmkVuVeL5jdEwHaQSbmnLGYF44dmbj4M7gelSpC6sEaN63yxf0BMDTC5ist
5KXNpJo1R5EHE09cE8OnTIYXsREZZF4IFeqvc0WABOVOxt8jJnM0OsBL4eGbk7wi
EfodjPKuxx7Y6tzMq73Ang72VAS7CgdpHA4DhwMPgaCX5FnqZPieh3zPS3oJOUAq
90TxPRNv6dbVJdzOzytjTXt5ml20UWF3EofLfJNfRTt8KFglVZBPs2m1v3aca28R
jVuHUansDOh25d5Mhtuc1Il38eQ1cUb47Pb+JjTSKsltKjkAIBbI/7hMZPOxloAV
HcwMvy4qiYZ9Awq1t9XOJywBvadM0U5pP+YQJrAolRInXtHRXHf5F1cLZFBh4d3D
Q3w8ukoJOxUcZjq2sLHe4KsrAchmBNbkuiuhGMyqBZQUTlionPRPGqmoYbCs3a14
oGVXdYL+YJTYZV8LCvYWFk3jbwpes5zPmYUOHgjLeCkMdA7bc8S6zY/P3jyfm5/6
7/SJekiL28L/yZ6L2lTkb6GF65C6E1WsKSKPKXITA1PcMjIeva/1UVo8t4XxL475
kjVTuGPkeDZeo6u1nUCdUHzl4f/IYCAFvGfLgqk6FaOFnLE8TCHBCeCcZXrPsjiS
h7u9ZFE6hJmgvLT4lR6CYhmJOf0LdwRGbGXnKQMiQl8s6MbRs2H/ShSE7VLgo6qf
SDexu8PqnnwZmcrIB/ZrgJt4WqxeisK0nQiD0Id7LIhHijALNt+U9F1cvl4c8M2b
TV+vGc551t4Cxz2gCvqOkR37Xx6Q+HNoxegkCN1ntepOpH51RSyrlUAUHjPJdjyq
/Ij2kqvRYna/46R/wgk3NZmoL0C+vUwIDtd6nS67LwL1crD0RiK4ZTqgB7gUdQD7
Pro+EHdBF9fHs9dqtPEjTycTDqXmZC6c6Ct5L7rtxfn0F9rQK50fWUMr87ZaLBdr
xShcwx+mGMtDPK4rzFyZQDG91zP4Jcn5IFmKc9t1327kQnx+dlDckVca11JwzDu8
Y8vy5WFa/fuSStEYIqXDXpF9w29l9ePkQCWluy66zqAxHBSbD+9ne+HtqCsWhGLv
Pv9VqNZDU/6UGKHuA3U+BkurkKpkdWyqx7Anym25v/QRrNCd6XJXvms/AOKibHd4
/lJk0ziQ+ZINp4sSWp0UkRSQrBYgnPSOsahUBxjfWT+rdTGyl0M9a23JUc2pyVJb
cw4KrOQt58nB0mC+kbXqA2KGNt+GO7W+5/AGcPZaEAj5GKIK5ti+zkcKQ4gpDzLP
8OmPDOFiyvyorYjlhCc0VOt3Bsb/BZdvI1gzFAXy0ypa2uZoCKAKf4NLzOxbtaB4
uBGARUumhmW/JZbY78LJHWJbjTDOETyofMlkkHsiK7s0/TiUHs1Re9wZ6w82MZ1z
/c00jgY/QlPe4/7whphVQixxzJCi92thTziPEcxMtoEq1DqH2mJFyNCxb2k893bj
bN7AxISfdHq5hBCb+w4OHmyLR9AxKxL0LFSTh4fKSJjQ0hiEZGKTNBRzq9PViQfr
6AaF4ndWDQDfJGl9oUMCbJBUA7RF02j2VkloJWN8crKzZLTDLyC7cawvFklmm8Z/
GlvXfLt6RingjXppugUfnknuXKerFlCKjztKzs7RfoVSdrGL4Wm4vkz7+clxOgi7
gtq31d+F8Zwo6wdbcU6l7DH9GOHg4U2SF490QmYt5yrohoTKVyh80QgFjIAEHaNP
xx589PM24YHTZYQS/369ljfa5+BPHJ03ufrmW+bQPiUsDLujzc4g5hzUbiISikSd
VAww6jjqr5pP+QxkCXid/PrhDcbWugvYpLW55u+JLqEylh4NBA/LvKaftpECWuSa
M1zzKrd+GevmJyjiANfRWfsjoGXaitIQMjz/ReM4S4v2NP0WAiU1dbJBSv2GraGm
GcGvGmE9eLwvkCJC2h0ATZIkDQJ8wNWolWQpOrmztWs3fw44qLuQX8QIfMnRoamv
+pxtNOWhk4oOqOYhT9uuv8ZMCbEkId+agziuJUXL59MfMZUF/shWMi3XmouyxPQV
ILbf0durVH8NDOrbhTFydwH1d6raX3FrC9Dcu0ubrhviL66SY6LMjUx6B/su1eLP
UqSHwJiz75aWey5l5v3IDBLf3lxJBziF7lGh8ZoQWv4sS4lcdxsFI/SRBE8zbUYI
xxnaMpjWSJuhEg8qaSyELkh6Q/bgsghsFIACV+2APH/obwCuEcx8HdV17G8xKg7d
6rAQa0azexbDBLxdrA/37m5yYPtfyi0lxDtVM3fyATOjuqkYSGGuMx+mnuW3oLZK
l9jieq/7IKsJwmgLd8RL3eiQ0Z/EsKbqJ80RjFcK6jiVObINMLhqNvcN/xqjlJjs
yODs8eFVsx8hchdXyCaA+Gxb6igK+JkqWWJGZPujBvl6D6F4ll8O8N61h7vVyVvb
Zy+QniyP4F3RGcblA5DVaQHMyMeB+2VSL/WDbuPqXv7XJ7JBD8xSJNS3w1p7edkA
SxW8hn7HL9vbdvxSMQ1C+8ar9tBEyvbFAQVPyiRydalBE88T4vVmSKeQw6i3Hxr5
iNzkVeK0agK2RSRORJCVThogYkittp1nyVPhkaXNKUYowWnpnhYM8lR0BiBILbKP
0Kk9So+dyDCziJA+rVxKddDoWrFBroji8K2G6rjRvrbzt4x2ZpxzmIA//AK5RF0K
SyKmSTWuYa4cz03Jxdo/ET9CBcwnYtHi4UOaTMFfoDaxGpE/jOVy0ZfYMoXArJJS
rc5P9lffpZCtfhHL1SKtWhHjP04YPjQ6vCOU/Vh/vyXQQyQoaHPpXvdv4hSCbAtz
+5Yws0uYKIcPEZXOH6nqIhZP9C/akgFT+aq5ULqXJvKw4rfu3/I5XAS09dv/Cz80
uSZWjyuha6LlcQZJH2+G25DcCGiL17edC2hGmq4zj1tq0jsvEJ5Sine8Wdrvtgwc
M6iUq12NzXlNZVkl5G7YjEOBprsXpJceLjBd6ZlsRUlBWVfv4U74ezmjrSEmYd3Y
KMNhAbjITEDADDwlDkLVpMFgJFfGwZyg3Yc1OV29KnMy3aiiTR3h/jH5Sw92aVCM
fu5f/YaOvHaNVdfI92YYz9tXScpnSAIaVhFbVlsAfmHbcQgZx8OuTexwu0He7NoG
PYQsb7anGpWbwoIaoiwq6MfS+pfDzy2rQpmxxUCv2DtmkKTUlib08dnWxtuKnbxM
LACDOQw28ZPPqyL4PsSfZUOghvRqqLwOlfyNNCKbSuTdLj44FXC/obOecboU6WpR
ZqZRSIWf7sW+RCF82NQr3Zxua60UwH0Uf5riWFyzkAIW/+8xHo+5lXlHUYlJcdJI
ibFjU7PANwbAyhIVjDG87VCyYlvpa+Reg2rbNqvtcKamngMyac9wzckJkOMdLHUj
6BeG57cEdkvslF55U6k/6FYtiClwo9sqHFHVHFkc/iLTSWgw1YgVQR3K0J+a71mt
rAvsUTg9eD/FVzWxL1CEF4svA1cZE3BLkN24gX+GnLW+XtE1Uilyp25yv9OiG+zK
CD0B2TyrSlsMqBp8qEIJG+f5fIfMRnolSX5YLQm6lKFphETm8uWQPS/7wPRr//sv
BqprkasNVTY+zCcStmIleTo8+3PLrZTHC8UNKiuITNtd3fqVZ+Wb3obTOKBGmf30
sZFE8Z7wWnu8/YZml5+9FGWMbVPGaKaFFx8q4ipYJm7sFPvR0T9VXkXPbYk5sYp5
Ll9krqa/bOvV3kCpULgDFyMvN44HRZ9KQavnpHSJSIHfby8S6ZNVtV+YELWJAaPc
1sSycjQyPrC0nH+amDU8guhGHOxz8C+TQfTjeYdoRExTOy4xBapYlGRw0bH/XPrX
tK2VuOFVPQ1nVbwTmAMPFTlwXtgF8YvNByEQl3JBTtqrPXtOBOrvKRZcLb8KcxdW
dj93cfHmpUAEJKmeulQt8w==
`protect END_PROTECTED
