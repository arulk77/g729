`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLkr4vnrV/9ptoqvlf09W0puuNhH0czrwvbKsJ+R+CcD
h4JK8BywkcU9LGBVfW4QSV9iaiEnbQHSrN+gdBPnj9omgjNYzqnQL3JNQdnpAHDP
xYOPI27xKWDlOSMHojilJBL7Cz3mINplrCkEVPLbraM=
`protect END_PROTECTED
