`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIZucvwjaBZ4y42O9Df34gGToXFstYxjtN8iOjdo4mgg
dL2V3UJBB+XTd9PIId8zX+syDc4dkfXUpz/xLzbQCdW8m8H3NGS6o9blZVC5C5lg
xd60f3TXFv88mdt4QQmn2bxQp8NcblDsQWaLXQ+UlDJbksyf3k1rMUiqQMxr0yx6
Qtga07htr6vaOWTLqEJ74cmu38YMZ1seT9zjrrdtux2Z8och1WtPxiW+BcPg0P5W
ul7IM7E3XC6LoQ5yWSq44s+pn6EQGxBUytHtdaCx3hMqMRKwJOTPaQE0EJiW6HGp
Gg41+RXe2bBOQudDr23QNtI71XsW1GpCNxkBK1aIuvQsf2lM35a8gJAVKQ6ftJ+X
bs38JlG+p7iyCrxoVrcNJDRAdDwyVPrM2rnVv5rxz9zuoxhtusdbF93gh5Ab+9Lw
8fTU7Cs9PrLW2x6rXbFr0zWMyDbY1Hw6EoD0BbWQqEA=
`protect END_PROTECTED
