`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJxBS/1UqXvyl3hTNIr7XARuw3+F95vglSuOSkkTSKnP
1RO/Lyt2RY4ObXSh4xqPSHffuv2B/A82IzrnwdfvsHZQzTt7srPRLB+G5wi14WTT
2jfTqnsIKGdmPF/40Hc5b8rNhARiJCItVvwUFooC9KILNocL6HNMRIPVT8duyGt4
wRcm4+R9azzu2CaDn5uxx/qlYnuWnYqTFG/TEpHz+YHaIjo+xSFgy/QP/Ju4ZDMj
oXytlABg1aM2G+L4UNjRPS6a33ar43su3ZCMooT9XXQd4dsUNmo4JXB1GRexiNs1
z9ax1ppL+W53rFH0nY7N8saPbiFqsyk0WIoFOlfzyqahE2/6GdmabOKCy83EGusA
x9OBQH0TrVoPVOm29IWBZyGE9kiTBfqfsWtA/gWkWAl6Wc8pHBOKgJWctTJZK/v7
`protect END_PROTECTED
