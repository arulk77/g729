`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+XUfISc+9VVl/a2eqfoUVFjBjcQ+QG4ZvDcIG0nkzXm
Gxdy8oPd1M2acLnY1Ed6qYXkrJtVgIeHU9GGuFxWxiB5d0AoONmtRffggFBpY195
SEFJw9wYQDTYsxr0QNhGsgmT/xdqqM/ZECyMEa83Ff/1VpvoS0bNuYtivB8mTodA
O9T4oHFtHZ9tbn2gnOoCfh0AW+wEojII7nw26QFq6jbJ7kyxIpmk1wSQJJoG3iub
GrniXedk5aA9hD3RS6mr1R0dip46UcKf6xkF206VocqyWrSXNIaPshEPrG14C/DF
RPUgHFLTngqAT4nvQpRZDy7Pm1fCzNntR7R7D84udF8dmUkwz7d4OHBusrBHvT59
l6CnwuoKysUzHTTaD2Zz17TZB5NGjp1bfZ8XolnRyGNMLpVqWJbcJPnUQB/RqiIq
q8La4M8AZMYGj7XKxire8DKsH9hYSI+Wfp7/cnpK2ZRfjtzgZwxZAbXak/oC8cqm
`protect END_PROTECTED
