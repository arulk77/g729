`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
W52by5FksJUdhgHLv4Ym9PrTrSkhdNy6DC7eK24hzAQyvNPu4x40LNQ2GZQTXAGX
Az0mmbry1uHXYy+ENEqfM3eego02uhchzRZx/qMk9sqGYnXK2pB6g+W2B8VScaCN
rkG2f2+LOg+cao5UBwTcwHnjtpEYlY9xy1FfiaUlJO3eh7V1t/BPZq6z9qZGso66
QNAq4AG1p+Gt/WHt+6VyBIMGNX1y8Lof7G9jMlLwFja2/aSxQB3Qsxf1GIXSHEtx
inPSn7GUr2nNvgMjWoWeT0XkRAYp0wrYdNAHTHrVvjSZ05hpZ9Rh76UBsiSk+6Th
ZZKlkRKogvUV66/1ABo/mYp480PJHIS5B39TTAO2v7ZqQE/wDWtD3oPqlG9fAh++
`protect END_PROTECTED
