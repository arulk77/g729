`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4jUYkdt5VjR8oFbu7ZiLkinpqVdbhuQ+85rpO6YawYhUgeCkQdUfGau1iAC7Yurh
BkV7/MFTtVDXWIa8KZbmtkzk1Umzu0hVisiRBNk69y4JgEnMZlP6/iWm3ASkl3Vy
e+p00p1iEIMnBdTdzOToWSyrThI2y+NtflIy8ZTlYclG22P/ZoQf5rHB/+B4jQWw
CSoPvckWxr4pxifXZRKNSaBB2drQ6UhFZv7QabO4EFExVOOx+TJkM6E/NImMAQyF
`protect END_PROTECTED
