`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOzBEoYPXSZvaApgQyCQKHW/dTTE5NCxTbOYOjEncdtz
A3qBDWJc1zEeajhYonqCDAWJki6IhS8XfdCS6SHkIni9rzzmMlVCqgpGxI8CHB+l
JfJ+E6xVhngdYGnzBlFzRMGfiIhDDw/qryh3Ui7K7PjPWjmfo+pmQGYAZ23MVTju
LCS9ZWawroRnudV3Jwgmrw==
`protect END_PROTECTED
