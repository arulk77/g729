`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHUh2h1AI5nvKrHI2/9Uc527GUIEV+oLxGDBpi54m9YL
AXYPVNT9SGHPOHLoyxrhWcMpgWQy0BUhGC2V8JWZMPe9XUKCMmWvK18F8GErJORg
2/o2S0G+Dk8pyKn3SmRff+/pnnlKlWMfoWF68/YM1M7s8IZ/Bx6qN8VuP8IWJN4Q
cF4L7DNkjBjd0aWmlpzwOQ==
`protect END_PROTECTED
