`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
i+OsWkvvDmrHSB20uQ3Eo1j/MPvcU5P7SoMVzd9bHOuG4OiErPcXZg1ghHkGAltl
h+cAR4QLw8E4GGPcUQjfCxwh05agZnfUbAQFTwdPYGD9EoI5FVoSRRDcG81SaYQq
7PRrR57cIo5YQIX085/VciRlmR+9Fhsaupuls1HXEjIuC3SNbPj38d0A43DhfK2M
NpT2YrIiPkOgfAiI1QotjITIvIHWmBba39SPZupyZqlL43ncOuvxp5LkrVYBNy6b
EBBJ6SGBB70J02Sm7NLh7sdxLeQuanjDkq7SVWe/3ngQVTL5ksmntbl61HbO7QmW
Um4+MjRv+xnOtbhh0mjyjzCDuo73U69XA0GiG42gFBQ=
`protect END_PROTECTED
