`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+7qg1di5b0hlJbTdaROAxmUnOK3tCdUPzkInyq9QZsb
bBHlqOBbEArF4SOM2rZFR7VqxZqdn6h+Jmp3A+T2gFVAsEIEOmSCcO5HngJpO6ni
MzJcYIWCysSMcYIRuFvYDGi5l/t56KtXzmOBL8GzfupLQQW33NZYNRG8RBvyRKJs
pnpWIwNL1s6zFI1yqKpis0YMfCPTlH2nnPIPbEJHpcez7HLJ5JWfLMYhPJcw4042
Dpcirhjoye7WchKaFPV6aTwy1UcYHHU970kDkVQsCDrXeitdWmnkdtL3VOndAd5U
3u983qLtJmSoSZnBjmBl64DeXv99fyyG1ctvEIyVZu6pbcmfTRu4vaYGNViRRVOk
//Q1jtXYk4LL3wnyftOGMw==
`protect END_PROTECTED
