`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
z1WzEOmjde7I+wamwJ7Z+vuuNFoiYSOsuuPy+Z/Q+wwxrD4d79wQR0dJktwAERkl
pD6/n74/+bRJq9NsUflvNndB4fJXh5uI9NFyWG6CAi90RIOAcDfRi7eKr1hngIfv
JiQrhj3Vzpp0HK+6MvMixFtUX3pqTXQDfhtM/QmLhjrivWLpZmkTUYKhk96wILKA
Ea7Ca0HgSZGtbW92T9ibXf9vEebSLsrPfmohNIfQvKENWiRYavSrciXXvwUUQNFf
DLFtFd49ki0ClfrVEWRAqkowU3gQnhpg4VB2JUruB07ZZy9QXUBmoYONfrjqBKvc
9rY8bY0kW26atMVoIfxhcxiE89W0rbFzb/jqDTOZ/gPulBRIOnqrJjHmMqbra48m
JanA8KnwaU5jwJKo+d9y6JgsRMnIrbrzmA+BLl5vWNwPzvl0og4QgoENSRgLkY3y
Xh0QdTCi3xkS8ezVQ5ckVuK2KQYA+/EWPIMw57z/czD17U28OURJSu4uhI/bLunb
2/wdcD998VyzTd3jCEqQKOQM8MvhacrObj5yseJMqJUDfvJh6BcZlu8qolKzIuM/
Du/Uw2xZwv2gzShe+drpEWu1IlisQC8G0HIy67tNyiFmoVg6F7EdCTqPXrD/P8bM
cth88J9XPryFtKLt1Z2xXCNv5edzLOkG9km2Uk9bAXHSzGZ622xeD2e6KEQ0hKXP
pDL+UVBOFPm8bm7ZiNPiWwoanV678/IZ4TR43nPJDqnrf5kvi94defYsoAln4feJ
pBlXfjfI3c+EUnX81C1kzL09aE/k3UD9rWQ6VW2skly88SxDOZ3LTni47t8i4ZmH
0ZeLJXQxNBm5Se7gaKqnro/NPWzjd9jOhgGTiYtWcADIv2UdRjQvcjzo5YBAW3iz
ypc0fjnEZ09YOBHj4odJMEwJf5EkvrEA1MZDTHxh/yLQJkbCKnH8X6zGogG5qCKz
ndulduaWw4VKFlHO0sVA1AFidFXQpXFhRNfu5fRzIC23CrlIb36pJvLtmiCn5UvT
kaGYGTutsm3RL9qY9RP2WBDM7KydTR2UyigWQ1szwCTNVlcuoE3mtaRcs7S3FyPL
Wcd4Hhqkvpr/4X/MRf+xMXZzU/6L1VEt7o7KaC3z0BjrDLE1pZcEl/mnJAE1KIX+
wSDsvaBabCayH1rXVY5KMPfiLlkuGelUWS9Z6H3HuRri30dW/Q/Oms5iVZhCNX76
5BO93zat2KHFzRrzVwbIUF6qQGIq0Kun0dEMckJqhzMjophhFWwE76t0zi5DT+HA
XyvTH64MHoWm3jU/7qivyZ31wAfCv6O8lcwYZNVZyvvFetlwu4KaPpZVxuovSZjF
1vrHnXzpTzCe3fC6Mp6pEei4a9qbvddv/qqiomLgKS4sYJV5b/pyRh4CBtiCRxHf
Kd7CW9XpGjYiZ1HtwHqJGZADsUgwHgboK9gcIUaZdBtb9bu79CKZCSaP7uYViUtm
ET6OMYLpuP4xEyoXvG5V3Q5HA07kflZilYEltGwf32pLgCn6JPyBmxKX7zwp9rge
wLTtayvZ7WDe+D0+r1Sd5LPxBJnBi+wxtPX1OfzMWheTQ8XaEaY/6SziTlQY4zVK
lLdeK5EuuUyE1cZQgiJL3Z4gYH4PsYlNevLcItLsDUJXIPjp8Yvb4c6ZaZClHmES
Db5itlm0SvWi/nCDlu4DzrgNg5Bo4sydvC7/1UdsdMTLQxJPZ9dmQZujrbdYWC9g
0z2IuVX2neeP1zVNFRwMGn35pSmEbqY1t8mGntuCS2dVckzPA4aTwQ9nH3C+RGqS
cQcGe6s1fBAWipBMsBdiKhsKfTryy/SoY32S40dxucuWQjuXZYjwWze7r7VcSbeg
WsNBrOfssUH/WZBYoEoDoFoOXhh3Odj8Ph9RI0HRPeVepJeC51RN3sspOHZNgFHQ
hXU6J2ZOyZ9iPI4r07mFTnuTzLgW8lbElI6FFUXR6yAWpaQUB/rducRRsRpIV2HO
BAQZn5XJEz9b7EanKlBCyThZkRXLXtvhjeMTKrALauqayvD/W10CXzpHHNSoLdCS
f5jtKExw6U7X59yZhp1jkw8j+bD3t/qjFmVEDPrYpF6WbIwVlhRnmzl1ioxK4cMh
h0CT3Dn2sHn1R8+V7hh3XLhwb5c4G5JePvy2gD+T0uEQ5KcdNqhzjsze1OPDWZgT
SrQ7cnGm1+6q47H+lTHwF+NrWK666dzXqBpeDb5m7yT+JCVAQgP0xpYQbs6E8JG5
RXbEFa8jAW4N8amnUWKEYLpCoqtY8FbGqcDDowxL2pPEbVfUylLhv7xQcKp4WXO4
9F+Pr9+w+md5XvEG2j9VaNs7KMNIj2z9xFfiGQ+89D9dQo/bLpbQ4gCY7zwyrBn1
7TgesOhkyMJ7xwBqpFslWD99jDKX+fY7P/ATfyEGim9MHk1qdjj62X54ESU44ipP
x/FWWOLqrRRa6uyy+kAp2/EC+/8FzCQiH02uMxYu4JINulbw6EmGQ7TQzqN2+Bbb
5YYWHSi6jD0MBkkXrjsOu28aZ9gTygGLbzql8Lg5841orRNvQ7AzXMoOzZiRdSAv
lixaLiKkeLfltNDj7c2eP3xM+ZlqIlgJGZEV4ErjjDVs/esVm2vBUlFEVG/pTyCE
jHPW/R2pIMfpqYCiLDPreVVaaYwrB+244xZhiH6n7vSYnmaVQGI2uVvNAt0ahK8P
BzuyoqGHCK36BMf0WTl20zGakP3BMHbLzyYAkLVLYlFWM7ppsVAstNqBQKdP1z7q
7hg0hLAJ+3XG6LE9F5Ho+1BZa/YR2jilmC/uihgMnZfNrk8txIm49eb62xw01PMn
KqeWX44l9xZPJTI69aVq5cLouj9dmdaqZfNkg9LNXCc1yX+zurmg4uypGvyu1bXb
rEpipcrlma1VScu92bf9gjX7ygDR8X7vp/QBsF7oWIBiXQXc1GccATtdAl6bIJ1z
bypbllj5rwXms4tqvcGZZfxDt7sXYl9kBd7zP0LaZi4mwPL9Vw7deFaouNS8idE/
iWQz00mZ29Yk2x/Q4Wh5fPFTjT84o6akOY/eoAEUughXMWHQwrjycmUqrnNh2oOB
K76+pSND/CNFJPK/qn4B4DstvDIo5EwqbRJ7eA01rnndLvHCfLmIXcfcTnOPg0/r
ejTOHyFUVprVqcb6NvSMqV9tPAHEaPDEIoqe1rAbc8CcZAADU9FX8NoIWXeiGgoZ
hS8dz5txS4iJf6G2KQlxFfeLumN+rWUjJ/bs0uc7fntvTkNPF92mrCbVf/zLa8W/
sjCvrem04+HbrGAXeUM5C2z+/10xYqLdRC5qfEZ1rbyfi5nY1cLfcxTBlVNtM6Tm
fh+KuWo+KkAwKcIatVC/j0cBC3NPRB6Z/CMvNIyTP5c+p8NOc5AkfQytPI/C0MgC
R+zSTYlzPvCLRJigJrpy6uQD2BB+POkA0dZvawGIirTRxSThT7ESGaidzkRrw+Vm
r2lc1NDl6htKwiJVBl8GAKuz7IakIYk+meIxN6HULFnXEeDZoF5KDwqFYRCz4WAk
8Nh7gNELaQKucmjDECf7+wff9aGulTiKsFcHcHeky3yjxNolwxP2Ojkb6By3qKJz
VuMpBcM56azHfNrkb19Kaf8LQbHrGUWYmut/5SITxDoL2paO7U8HFpHGsnfdFxJx
pRQW5zSY4EWyaZbBZKwf6HOEE+N1aDEQyxthUW7B0MQsFCSOuHqDBPKOdPuZc91d
ZHvaz/iWcZmajXJq4kNvLedCa+QK4MbJdCyJIhDYxaUbOtMZJoI3aiCDJpRIE/J0
i/E3Dbh97v/7ojVBcvVxRL5PsuaLqZ8hRNSh46ZoxYreDMyUp7rsEpR6fzxhPVvV
wuRCNRebdyzQYo3slO775cELCmcslKpVAJHj+DvTdca/pKbTQDxQ0oY0znL6HWs0
GiUNCFM+ZFsmoC5zaTD5f5GP+HFPEs/pn98QG29sTzQ29hHGOjJE4eYJ31HiYxpS
o5slhZMy0qNlCNX6xMPHQCezOMQm5pFv+0SxGBcQia3q/8OrvqW+dghbtK2tfQqI
C0EuqsN+gcudFCYpu1SY/qdg1/okExEUIFan1bA+xDvw1zhP46ckNL03EKIPY0ZC
xF7XVj/gJ+nf6vhju5eiR6Hlw3dg+d1JrjK/VojMbnNfFSPDRurQI3+J8s8cc0Sf
mij4IYQgtS/+3MDcbS7brJSIE7Tq+JRYnngyRMBhS35qzPIpwUX5ge17VjqcLwdw
iEVSiziuoFNIQNVTUsR6DIojFyrKISayHei0w6xD0O+KsNkU1UIzgzFj858Xn2p5
n5xvMWKo8h1ul3l6jngwLgBxNvmpWMRGYOT8+MByJLdwmYxzYsxzi9Ms6QE0OQ/K
N3gEIukwWLDl3aaDx14ILYk9ulvbiqm5GyM6+a4iAodFRWa5oJks4IwjoSvDiVYI
2f6GiNjI3eVUnJFYWX4VOv6aviG3CCsoMhmNXbt+fC9sdCrm6IqWeBXHy9rWJFRV
DdX32zjNHDnBmFz0II9AAX7Bdw0saqX1eROxlR9Cid7AE4RHAvhlFbDB3dQCRsJ3
IbyR65tTUMv99TiZWaxXG7TudA+/wA9VxvzP3osjweBr4EWxNbgPFz/AGYNoJrZ8
0Dnrv/1hfxJeU79fEuagbQi9SL/WfzLxOBAL7AReJxuWosiAhtw0akq1XSsEoV5N
uunxqzsr791JQ1AzEM/Bvt1Nhe3GG7g1ljSjm4hO+XTqCj9Y7hfh3f3+ljVKbMC2
0LOWckGjU2V9h/lpet5NRH/tTZ6+wcp/Dpoi4DXA5hJu6DOHCeZff0EcCSpf6LnY
WZfHuB2MB1YFGm8kMt1OSWiB1e13NykbZynUtPZcmXqeteplpNPc81uFtPXWpVTw
xIAiGDud53FHeY/Mx2Lt+0Tjfm0+WeG4M6bnf40J9emOg8TnW28AY/6Us9izA2aS
C0lpboFHS0CEhSP8/sJewnEQpmKMsTJpIwJpgZNEFSpj1TemxqH5z/TTcIDsxDuz
MG3FFMZBAlZ2+g8kUY0+vYeCeVo3VJo5S6AiK2z0cVuNwi02VNnGXlDmg5qW9tIo
f+b849GpAzPEdE56fQuCNZootiot2JXBwr1wZoSbBmkDxzZwCajVH+OYlfry3U7T
uTmRX4F+PADy4kY8IjeBrWhedNj/l40gSrvjvhX3sYIw10tRnjQVK3ShyBuPcGi/
UHcZ80UQLvLWypVz9HLS0ZIcA0HSzGW5YPK8uL3TaEOKV5ZqiAd9hZb1TUUCz1gy
oJVKUZW9+GRry3IHGHeQO55FOdnOjgNJ8I9D7viSXh3Iuix0fMbTANx8XabSoB/A
M/QxpUUmzm0jWAZs1CgYSRbVROU/u+hJE5BEddZAyvGRtFLD4JyosBMgBNW6tKdH
XrU7GVGcUlu68y9JYl+uQMTiKwYFN3KA/O/PvsMy1qXHQU6OCFwDZ5vH8QD9l4Vv
UulFxX3QU0CueZGrR69hyl0iIlB0miDIVV4IvTRL6lLynaESmJWUFUAgqHWT6Hh9
Tm9tqb5JKJPXbxDgqXrXodUsj1y2G4KAY7dj6ZTK/5lL2KbLAXKNndYrTBfOWmSB
s2PCdofDYSYmYSHFK2jDgtS4VPFTiHjSPdCMSQWMVznvhaBvY/gJmenN1b+m5A3N
DIpsdo1oTRm+qWfNwuJF6kytYu1zA07DIHzpoLzBO0BpK9o0QC+gtS48GJY/QbYo
D611TZMK7PbaxzmbNL4owUbe6ZRJsKOBWalHdDFrBD8Tlm81UER05Td87p9i+GqI
NsY4TZDZkPJKiG/MxP9aMMh5O+pTLI7W7+7TR5FkT1SaOAi/rsZhmTd31YyNvQYx
W83u7rEZUGu/jjinnGb7yR3z/U5pIjnMX5ZKtQu1JfOneFtRtQhy+hNUd5MCGY0E
jnDX7jSSf4PRJeHDvIx8YZIOkVnwkWy+h09An9rGjzWY7F1WhzjKdWLeJFzhnZmn
ibF68YbMWe8XMX4AIm82+2up1iVu17kL0BgDE3sVY5/WEN4Fp5iKs6SpqKNXpcqf
/AgY7AHFw9+DcN+GI9lP8CUgDf6S9YO1KiYafmYFOPHovQIlxsh5T+SHPllX6Cx2
2D2ttgPWiRb1UJfkG1r/fp0zCrhn/3K9p4AX0iAqWpFmn1uZMffsBKcdGi6mu6eY
2EqdCJDjqH0rhB/gc70cr0CIusOcNo+f32p9KiAym+NVKMAYhAIekj7zwcwuUS1K
vP9ytSZV66puHV+rTBzwPCVmEz9ZsbDH19R1ztrKXWIwQONutDRn7ZO7n300RmE1
WdTxKQh9R9LzTSSDarJ0+Y4KSN5pswi/ebvaT6Vd7jbe/lFS2+UPCUsxrF20qVk4
MWc2utGxUD4CRNum005/WCJww6PS5+59Z1gZegsycLRTdaVl3zgdcAq8QrBQMr5J
+use1Z2jb+BsNps1Z7s0trSlZNdb4b8ZlMMgwyeKp3C/MQgAjLxmrY4Hc78KW/Ye
3rJMJ7R/sJrNzt+/IupiucLzWhbEVw63kezSsP/xLzbhvMK9kp3WjKXT3yDYbInR
0gfM2WcpCziIe8H5R1zC1k4WhLJ90olDptNv+pyM1Leap2UL7/75La8f8n7nDZ+s
8qepSYfeWQE+b/oeI7UuWThw+6eQFIL0Q6J38cMVllupRZC8mcSvRmZB1eIVk+rn
8UGvR/sXtcuVe+pfImpcROwFBLgJH2PGFFpr2jArD4aeB0R6vj498YM8MoZW1GJ5
BvYBMjwkUzyUVIkDUoBxkDp9tC8woKU21dMzZzt7hYeNO/C5GDugmxBnEXc95vi8
YDBTHI9qq4/0agSVLp4Sbsusp5y+DHdOdv+QlWJX9Zho0Bt4JGvx510WwPThWLD8
122SY6Jkt0aYDDOBv//ml0a9jneI7TQ17WEXyYp4BCd7kDY8/VATjDqH74kqK1Re
5EPzKRTXYYzX4OkseYwzULjBRaDQzzgqRQfsGb/RFib7Z+QPO4U0FZ9Zq6/gsUvy
eYqOO/iENbvrztkHrAPEjIJQlfPj/JODjX9Ln0PhZl+pmT3AmtHOoPLytqFI22bw
9g9qElvBurxpw+v9oeba2gCNjDsHCgKhZ/bHpsz0MSbSOWKpBDeVzfWyHYyuR2Xx
NZl5M7s4hKRCgYHWRNPeXksJ/kKVgk9mm6araCWdUJWthPvnlVTDLfI4GFNZPrcC
cWISKQ040WpvmqhvI14Po4vT6jmd0nXeZCV70LTca+Zojd8k6CKL/CfxGCj9V0yz
BQzn97pr4ZdufVEhMKkSvIr+ny++b/Z6pMIAVLo/EDGAbTpXwO6g5GaA/qlw++UU
dsCnTls5T/HKtUtYn6xhN+59fwxuaHEuWlpfFuQh/ghJhLSet5XFnAwAI51I8W+9
sAOFIbQ3pMtyUEje7yDoURXDPs1lDzV7JKCX22ugCTfBp5J+f9jOmVEJy/Qf8+Df
6IqRr6jMHcScqQqmRZINI2LCedvs47a0EBkR2SVLWrtXaG88jNYRl5OtAIKZn9wX
q17xVDGn2Oye9yEjEM1xNFbQdOLrqLCuergl0fuJpQjXvparHn3pSiirUkAJAEzk
cTQc9IXY5YQeXyGwIsS3X33SELGXupW23/4j2hK4xAE5mtUmSdmiFFDvhfCdair5
qd8Cg++plgOAhkzXyIwP+jdQ+toN2X4MNi9087GJEvageMRtAievkpuAib0rV8US
ymABupy707hUbtv0s3Eal1HBSDS4M9e4pZIiIx/OuG3PPiPUXB+SxuWY/Und9JVi
+iCo6lziwZtjiXcIYxnvq15m/shTupPnO3HtFOpslbuf5FFun9hELxe7t7eBDSYG
/R4RCLDT15ln7aXe4i0KrPsTXDnpovfNcIZ5E3xhUsN9sMxoOgE4WbVIlK6Pr3wH
CoUMF5nmEDeE54JOpKmN09hnO0ew6O3+VPxX9VdFyxTOwQesegu6I935prEOU74Z
APnDoLVFNBOYlYvKCJgCl72QJ/wTofBIKoMtBswhJ1WbxUaQlBYiSprfNPvVKxt9
1TFgygqOq7pxg6MQPsc+1U+RTlUtOm76nJb6hpT2XjcT+fr0P8ew4k+o7LhAIJY6
D/7UpvhtIU8wSfF42jPyNgwcMtIkCHamgK7PTUvaN3ZQHxD3oNB6EDbiaxD88JX0
PPtlzRV6630jQTpvC44IOx8E1lHbKhK6wkA5pqJEl8CGftgo44JB/4D0bP5ji/Db
dgwoo4wRA21IbS9UYcg4Bceq/iEtljBRM6gc143GLNsZ/efSTV+bgvQ4tZJQWKrV
xh7zIL/SaCyzOW0VdERwkRB/BFBgQf/Se5AOjByS2ZUpdLQLadVpvHmvCNMpKmxa
Edmyei/s7seSjw6A1L0/o5RqsvfukrbsW6wT/Gf+VRQtewy/8gLd/91gD0W2a8lB
Mwia5oiJmxx7o1xgvcCukw2WCVGiC7NEpScxpYqFPDJtdz/jpqyn80l69W1Znruw
6nueATQPGjw8Djtpi3j0IaaxNS5B5gX18QODo5802qxVDVYz1ZX+ZoJEJ2rUkYRf
OqJ4s263g4r4lHU/9aniWlFDjjksC7Gg13NuYOq53D04sZ5Vsrk9Y9PiUP9Ln4m7
isUYzHY44s6+rsoagKGEVm5jZSlJ/G9mx12WKZzfCmZHj/dX8Jpy+gUZN9s4o2fb
pRJNhqmplcD3Mx7LcXHkbmrXrcKAwIqZsUTS6VYVsHFJxaCpGN7uL37/lXfG7R9Y
rZbz616ExcK7PK6UWt8FwUBr/EoRvUsKmsQ9wxQuBS53uwFb36kJHu3b0DhcF2Ol
tg9CWUERsldi+HORML47SDUX2EtXorYE6ssJej6/hUw3BjtCHW2aqUAKs1YVBE3b
q7wfXOFASxNV7amiGRZ8UtP7l7Q/D9TGVbu+2vzn/vqSwX39yfotZR78R9jEp/nQ
SRBpCUlX6jgn0nhxClI2OHS4oV49ouDAK9jFFrkrD4nP2m/1HRh3KTC00zr2wrYB
wjHNaCzqJC6YbffUZKaw6T4C6bfnC041JXAz2Fqyhp4UFrqgXzhRPemWdfK8RSTo
LRiqT5FhxqJeHkieZEdweFDKjp6QIpbqdYSCNtHx/JTnrK7UfrN+obd8Yzua4lso
i3RsWo/J1QCfH3p9jWvKtGpBCHrVpnOpSJ6zYVOKJdHaUa1lfZOxIZcpcLwoCVh1
X49sqtnrvvy4hY37P++W0RdxxNDgCg1AKUuRf/1jgVNxWl8P8LgVhgEc5rQRh+5O
R2r3VvGh2D9bQVfkkRP2yBXYFrLcDaH1E9OImaiMZv5ZhrA96inMIuadm6LjUHH3
gFVTQ/8Iao2rQ9XSbN4AkDGlq2+1j/9xAOprnZIiMvlDa1HnjLoxngb1DKfBBP77
/f6VrTqrjF0adRJOa6c2YNpkgkOChNaRaFfODZuoMKE1reBdk0mONcnydiu1qIC3
pD2tNN9BSsq7U0KWD43nFQ4Qlgow83UvCfChc/WqQm5JMgBkhhYTCtoJxAc5y+Vf
LEpZSuwvKdki4q6qO8K/tHfft3UygWIE1nHIW5DSkwZ7hcggVzd3/cJe8v6bvFSj
sP+oOZdbyaPQpzEJ8AHnwAXKufQWPeI5H2WXtNrbplasUflZ+5IJN3InAOtUkruo
LXBxPT89uqjvAPGFw5Ewtjq3F6OlxpIssl4ofyCVaU8sfBMiUORTGvPqLBOjZaUa
sqgQ6KvG0eN9cM5s8RGzEGAZZineDEilTaF7YlVn1ucXwr5XJHY1fu/8M4D+cM3S
w/lMyBLgv9ReifdMowWH+0erCkfBgqTEGHe5RStvgeEnqrEPcOt/ylV5STg4JoRH
EV7GWKaZnFy6hqtt4u1S10Oi/qXbCZpq5yITGlPtvMnb7fX5Jh6amGK9gBRoQyZ+
4ab9PilTGWGl7CSDu2ZP/7ySWSZUEUe2HfJqV46XO6KPK9tB+cbyu+NH2rilTRTr
jrzdDcSzFl5gGbO6r6m2QtVqBXYFzzBkgY9fjE+eY4cGvazdX7/rWnb+PpMH+or6
+xp2k1/W9wO/KxysYMftvYVgoXh+hSudq1vL1qw9EeLkmXVN26ZjUULqQBRxX+Qx
xP47V66FQE5y83DPjkkm0ZoTx5uhlhV7Up4lV8WUJ39z0VES9qHuNJH5fZwFU9ow
41im0rJQsTSCOo4AmRpZ/+zQt0hjd3y/TG52l6sTemp408LGFywi+CGu61hMrQc9
hxnUi+UZuigdnFigIzs3/saTErbyxbXS1P3ni8CzNigXOJ0o6bnzbIrxto/ZBnLh
TKagrSgZ5qlYx7B+CctaL4lZ0qkWLOvPbBEMed99/fheJC4vkp9e4RyLwg65NNnv
my6gy7XAZbJ0VDEqhtQc2SY/7dalkdsHAtz+5P2K3DQGqFWzo8+5RAjIZ18nGVwl
JXVvp1/DTnmi+r93t0Oo9QG2jTw+2cD7Rd1m1BSZW4QOl4CUJmYnvUHTLqwS/cPB
y5wg50WpxJBuw18QBkO+iD5ethsEHDqTNjUMP+BkRixgobG/bLARKwRMmIQ4ZSwj
ob2jglepcIJac5hqgPq8/1Wm/e1UNoyLGiscXeoFLtQvNzMsWV/pNJ+UjEukFheL
HN3DFcHZHVJj6jDdVgOK1Br1FDXbN4gq2DylbcUbSddqs+DwPx6tyw50ypP/BzVn
wdnSrBh8C/oHS3xVvw4xaxRsZ2PSDRxAcdNIGUh1qomrHPAUD8zjNaZ6Tg4axF0I
g5bktB/hN/kAZzKvK8Bj+oCyOJPjf4vozgBMk816QslQmKfObDAl0d1KdghL3lO8
HwufX1H2TSEKeIq0ZWja0k8uUphpq+g+2eOtW2qec1DySShhx2w7RZwPS+5apPOZ
uLH0j6ioz/p+ogryh/QF5NxASE5EYdclbrrWZb+37HF44rkrhDPIlVtqissDt0x/
7DbosyCWfE/jvo6AqsSpg5wBpwmVZJqzZ/zznB8S0DGUVByXLblC2s8nbWsRA/wG
V2yML3bKEZyNiX8bQTQI9UHlUflVnrJm1I3w1qRToe2qkdl+dY2sl8Z1CzitJByt
HT2c/NlJexvFer4q6LKnQghjuog4FZyHOA2G6G/LK1tqplg3H85p1JIhaljhKiAk
Fjrxl0JjzQxCjbYPNdFT8KsucnVQXQ4XMJenJhP+egKcZgTbsEZcFWk0YOjZQvMj
XHbI7e0+aDJC56S8r2qKTnsACCd23HbjQBUo0WAOWfwyp2FeqIrFuG7asqEVEr8N
soJjzwBU0fEL/ZnPRXTdkDJ4jEfXaavBQ6vLfoMCsWPmIVId1ULMyfT/RSGE3+QR
E9tnsVlA5p7tQ/UTX/LuMVbLno8tEJgoaYBt/Fi1JRSAMAgO61ZRygtbmJvEFaO3
pFu1DGX00qnFbQ58Lxy5u34ylfkdm2hPf2D5Jy7mWHEXvc2+x7STLqLUcKZN97zo
eAIZFT8X+U2OW5mT8O4xhnTP1Tid3Gm8Nbi9NW+o/hlYdt2JpavdLZTv5fj7EMeV
32en+An+CUkp5GOOor6dtZ6Y5rmepM3e9asysWwuedcb0kfWhVA3ys21B+6a3uNB
1i6g3jEvtFfHPCiSWuXfavozp11L7mNaMFeGkZBlNWC7zVzekNpUQjRPTQBYtW0K
KJ8BwVE9JRSF6wRV3WSvVRubBv7pj+hS6GALZbS9jTeI5QPtIoYZH+IZdS5wPLz7
QoB2WCEm1w0vxoehdKWV8gyx0GP25Axq97XgG/fvVXApH8Dkt18yvXg0oEwwcUAa
h5Af85nWQGTyPls30DWQd51aKxqIhj3JIKQyslpz6XgN388cLhSG/IMzDohOX6Yc
Y8kpY8mm7VDU5i3/A56CFoqPDGTcp03rK4pfHdueyZbXbUp0LTgxr8H0hohn8cBw
Sn0IdZEuXQlOqSc3Ritf4LfOwSMI5RwSHs8TTiiqFGBj9UnzmJ4H5uWv4GmzaDU3
82LjEaPUaaOo4a6ZNvyK/zTimyEGaZMrtPRLx/1dN85xpQllBLD0voa06M4ZB0+v
1WraIkq3v7Aj/QocsDt2b47cyuma+Eiophe7POlO/m0nFkzJM3/5ilmXyddpa9nq
8/nTcCRWG/hRvAM4ff2goKkVgnlU19Y7Jp2gSh5F4/KvHvoTLgq2SiM8XtWIXf3B
ojOPtsL+3HNGVwcDQH5synd8O+kGozveSCcArDMDBrql4WHoZRUaNaw3cLrTWYn7
S39iVS6CXvrrz2YgCCggxXUFgLvXm+ZmavvPeZUkm83AMSBmKTrM8lVxr7+tIM7a
udFE8G+0EJUtkTuY/5bQd4rIvEL8E0R8pmjjpwTyjXiZ1AOLdjiw55MK3wUyS0Gi
eJL2x8uSNDYrfSRRCfV1dn+gXbXj7lS7hx33x2TlDyc4BFwddeyMw01ieoxwQOPD
poI3pWlN7RQjqEpXv3O8iUt7Qe+imGoLRRLYtCoVM9cfu0PTCdavuWr23m25jrP1
ci+L3zO92blSjVF5Y7fMVPR2md9ul9vV8tj0UoTKKvIznjtMUGxEhNn38mPXHr8o
1kTw9B9nQ3k9Pl6vJc8mSpxIY9//BXHnwzDGLl2wWN2dcMCg5X8zUQTAVAusCG3/
o5dRHtX6bjCwzTAAe6Xaqg7u2lcst1fWrnwR38EZX+fYrVTHv61FWb0nQKo0zmFq
ICJ+J4jZgjaSLsexQy5X+DSFi5nY6AXodhs5WD0WgPiSZYUy9yjrm48iJk3w6TiK
ur+2WZWiebdCLDi5HdeQsysBF+kR+f+vkFMv8PMg9pR+23SWSYcqxwCADoZJ4sFl
swJ6TIbCcPpt5WL4Emk20dquI0fZH2B5KY0VTOscUuspFJ5ZU3+Lt8diN4TnaiFc
dXuHZvIFDSaMz18hbl0DRqnZeWPybYK3tcPp0r+mBYY3xAHQ6eUoJ12v2pbyzgdA
TxlX9bKXsBaHydmHMIcq32SFyW/394ctUSIy4RZLC0tzmfueZiPsSlDOtJf/Ma2d
K45MkvYO1YCt1hDIqfr0ZH4IjXmY5lZVHFdJlMgvEviPtJr79XDBCTgjG0GOkcGk
9Tt8MTXQ1ejotS4gYhPu73CHKxNSE9tF1s/ZVB5RGHsKHGOnqdo/H1JfOLT47NM9
dQL6BJrPzgqjS0AIJVRCMSri8Dl7amJuJ+2wuUBvzSztLBxnyYtelwKnbM2+UckW
sPdFqnmTaY6Gm5xAqDKwbL54LVaHgutFKjnqRNCIjBJZVgW2sYKlQKyLAYJQRFUq
EZpCetnf1YwSXC3Uuu2fj/asuiodfGPcbvmFq4i1Yjp/AbuyiXU7PGcKYgbm4cEm
jW9/Yb90bcP3cBK3y4STZ5aQAFsCdD6S5TTkDquwvl5r9T/A1eaprBhYpKwmbzNP
d6pxP62dGGdu9Ic8Jncp6oIz7JDUJw2CYVSNnhcLyPKjmXgKu86oLdqpBuooT50n
fn2km/kA4nMGWctpgCX46s9OSwwPH24huo9izaXJmxLywy1EEZ7qdQeVcsx/vtpC
UGu1ULOqJRWpVxRxAbU/8ztAFOizsRyGNyyRjS+ujLE1xH50ZBdJ9gdqTEryU9Op
12aNgpM8llwbs4T8XXv+I82A8mK+RpWup3dLM9kOQVT7EkkzLoBimJJ1aciBf7rD
h/6PMTRvx3AHoXxYEgEj7UhVHa+J1kA81+aFQat7NSxuWxbjc80SITdlqWqDcrCS
dMqGGp3QLUj4IGcmd9z6207DeBOSz6yZF2Y9ZwL/F2d7rD+4lpl35WwNRiB4l/0Y
ZQYPmGun3wU2UO06FPhM0A0LBDv+cVTgyF6K6CdHTmrjqGM3nLlXi6TJP5Ip3rye
+BJLuj4nxYMoZtH2KP1pr5vOz02zlHJCYI7dqB1oCx3h511sFYbg9C6Nmj/ZESBA
fVyIreUtUkobwM2syFK0HpvZvDsevtwUSXe3xTUVr6NDLRVFulJGcjheBu6SbNgH
Uq/3OkdBHbwakR8G7c8YWo81988fs+DjThc4yPAHJz2vtueOzRzkVxNZqwBkSlT8
sPAaKlbSutGNPI/fDOvUG/23zzhzgAP28+zy7DVOvGxabiGiCF0SsWwGtOAWJ1si
lxHJOMDbJc/O/K0+IHBV27k85M7iFEjIyuIdNbV6wer7CbPNmjIpeEUe8m7VKFfB
Fc0qx2k6QMARycL6f1EMLPBQkJI/ef15xPQYqFp4+7iDemJuDxwy1NP8+l3TqGoK
oIIuZfOg6OjI7NSL+DZ2cE06PcMU20fQSAE6pblWngWS3yLMwPzfiZsDrsosqpV7
8lA2oH3mVaWw8Baj+C8VjwOFQuasKF3qcUBm44pZQ0I27ehpnexfVESoP9Y/BTpB
nCsjm33szNytCgZV3oy1mkfDfE6cmtrRbvqh4fpXR3oBoRk31BxWOFY4dXfny0jz
obmI1OnkNhvGp4aS4OT77924gFIfhe2XvECCTguc1bLG8xx5oyXaxXWUFwTnXuZy
5JJVZw7TsUlS7SbRqo4omeEwxWazLGbSUh1QO60OLULy1DcEsi0v4OrPGLNN2twb
2NX8QWczDTu2GGkMq5gubk0VKZJiErFnsXOUJZVbn8hUkdqTETOcIZVB2zu8UbHw
BYpWaiy9tPzkeFd1ZMfDxi1rbhkkPzfqgBhDoP2z/1KyRlOd6xBPx0/MLH3yvr2h
JjOAyyuVD5/SkxMGCrP58GA+zeK3QQIBrKpfGADhHDUmA84AV1aHNOzM85wXWX4U
kjm9fIv9FO3ICVki8jF2IZNphBcbMCYuE6cryuma1odpMmzN6gHTkPoQxjXYTroO
Bb114/NBWIAW9Pyc4unbnoW2KoBTcqCZCrwa+YPbgsLl0dZeO5rpZRpgrSEMsa8z
eJI+iofLPc4gozoElWhboY5Ah6gyxI2mvtag6LHl+C8+f/ggoZ5lNXU7OxPwSSvL
XfEebOaytaCY5Kr2++ZpeFPUqqheT5D7jtf74Oa96JIEL1gfyPSPJkpXlPyW2NFd
i/azWcK5jHGvTDiuqmXdGvg2HIlM0y6pThoWOt7Gb5UrIMSBaOSmftqN3ymw30dP
B3BkjrNq6JRx8VGOb1CGy4oD4Xa4QzmMBJ9lGS8U9NIrVvnxJddmc/C5SNR+0EOX
SO26bydqwsVq59Cl0cOI87mvq+tJRu4Qu94TCDLt0rIGvvIJAVzvZTJ0Sbz0LufV
kkdU7BIizEvOi90XChVUd7XJa9xpch0mMWkkEpn3W/Wc82EHYTqSeeXyNj3n76SB
6/jT0MuAZ/MlE93R9su4OXVD+TOqa2mb0YG/Jus33l5VBmeSEsP6RgDCnx3w0YtY
167VdCirNRU6cBEX4H37vTUXAJil7pk09/nHXyUwlBbOy6jDEKMcYFzJEzjrJfa/
PRRoZiyIC2sGuEjRMaIJUVHwXePI0GulBnsM8/tqvOGwPJr5U5OGa/5oo/zS/1UB
lgk1Nh4YQQwYmqaaByPhU8H52tHlM7gAzSXFI4t59LtqH0QePiqdy3ctBqW/BV/z
nwqB7ceafQMEE9AnJedD/t3Ln6YKGG7XHfyAvaLDE2C0i/JBdE5f7De+GENsMN18
3PU7Xngp93wBF9LkKXrGsdsxCvx00cQkpCg5axlLOYTEBLsilhgRWR9rSpUvcfib
AHRp+r3ToPs8LY+Oed5z33r6ykzBwFVb5FTNaXOSIqNeLl0m0jtT+oviVYUiDmQ2
R89it6g+GjcMc6fiI+L+oGRdS3sXRr31qBctoSTYTwdgTHL5DHIVIvwyl1+9PR2Q
8qDjnHIbEQeRQJFtDlqEboan+PAbAERorxC6WKW2MLVWaaQjOVJ9Jp5WNe1W3V7d
mGyaYilll8E3M+4vAkMQPi/mTw3rzvtVjSPd1L4mLTHoQUQGoIvu0wj9LNm1E1At
KD8fbdaMDF8uPT8F+AZOPGFgOJ2ZaC7PAc3+NbyTez2OnWQMjF/kan+5nA0oIxWz
vy+D4p9wQbWoU3R7V8hX1UoksfRCff9Dx00LYoGIjiNgS3XiA4PEhS4FsPIdUTfF
rtnRhSdp9ExAaUmsSlCAhDtqq1wPOs8Ywj+8AIKrhB5naZPSj84jz8v2YS9pJwL+
BZwTx/UmbWtOHZJ7i6Y5xM0LHkCP8TzkGThPAgTTjyOhLme9QjjZW/5QLffutaq0
oX58oo4FfyD2qvW2f1820xhQD/e9R7X+qo02miSwPgmgMmq0q34LlTf4mXObNBTE
C0mDncHwpASiXGmEOsId9X0rDF2FtNE8XfpKN4wAJp7LMwZXWtqdp1AmWWI4MxWn
`protect END_PROTECTED
