`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveO8HjrrlYvqL0yoD1zuxNVLwXivKQLiqJbhXS0xM9R5M
RIn9pRKr+jT9OZHrh/EGImcDrI5bbRn6ZejvS23d41HvfHbUExfxkn742pvrbUoc
6PaXGNi/yO3PWPVVIH4EakwpatgSEoJmfkhtJVBZlcr1ySDA0Pi/5xb9oIbdZfmj
hJ6CVWe5JdyTN352q8WIwkLnL22b6kQxbksBzrjFR/wB1YJHkZDQTrVNSGRkJggR
MwqW/TVS8QRzdzLpc9F4n8d0yx/wcaRkn5stW/B7vDINhx2/a3KBgG1si1zsd5Oc
YNBJ7snLLWwTcbgv06cIzTLXN3foOp1JNTD6KoVoTzIW/0OVERtO+ZVKK/2IreBW
`protect END_PROTECTED
