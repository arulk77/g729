`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
OakNWG3rsVFqSFFlnFzW+Yk3Wql/X5nF4Mlu8bfsIc4Bx05Cf280gDrOGfCH/MV7
0iLIjx7X+MK9IHfXvTjFVOpKF0GOwLR0WZtZEgHstiNXZIqQjtwMBVXc7bsTRF3P
rOPrNNzy5xgBbfD1bvs9kjTiZT0ZfMhRAZoDgqKMMLgofIv+k+EWL473XkIw8pYV
1yK4UpbK3FF2+2xBv0v4JMNe0RQ5vXnhPrLMtsk+27RptUBW2l+Icz7tdL2cZPkL
zlUm32dPIGlf/yGEg9ICfjF5EZGh+4fjIJqx4mrgp8/INYDEKtAkH5FDUFwYuCiM
5yxEZCBJ6uzYdpsARxcPM9BO/gvsJEK6YLnvODd2A1NuxB9wCZ1LNIj2kZoCemml
oIe0Z8ymuL3uQdihfkjOLr2UJKKj8nZCft2TORcFLspoahnXyELn+gnsBse2vzuw
YT2XaqOzB5BjHn9e0D2930B1NAiJoXs+mRjQhFNufTE7s08ExiuQhM9Z5gkMkeNb
EhwRTi4UGE8kC+odT1aNvO80tbZldY5rdNYBdCQxJs1LH+CVynIhPg/fpXDSLNNR
h5jrXz6gsxDrqTUql1bYhg4w2Kye99ZfFrFiqDDWSRY2XnMm7rInzpPw9IBLnL0f
`protect END_PROTECTED
