`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJRMbmgrtPIlHNu98UAY/bDay+cDRmjswsrBttwq9W9x
Uj99XsKRjUE4dIylXjObplGkXwEkjzb9GuCKFUHMvXRsP7OBXVW3l5csVGFkb1+2
qa7bOo9nEnOucC1uCgLddWplZ8ajZItz8gP+4D0+zM8bsiJU2fATyTdjoK7tV0n+
O3LkCGv7J/jOYLK2/8umkcbwW/ZTNncjVx/Rd5QbNL3MQfp9pO8brnxji3veivKE
fToiqchoGh1SlitN0QVhoESlq4nphHGwo81myVdFCm5WYOOTde3RhzsD7yRdukYs
cCdm4kJqOxXbGdHiXjY72Ht33SosXjGcAobQX0V7X4rpx52cFuyjd9ABJcSlFjig
ggo5yTCFLchdcccoyoIxdTad2e7OGjkEM92tv6e77vW7VEIyuHHvT1sRDkw+ldSj
DpkEI6P+BVesBHZVToL0I7424REwq5XlooO9KcLjhN6hMlyGJEMjJvllQ/+X8iLo
9nbC/KeO2RvIkiy5QCJKNLNqn2xtQvwFDEkINVVW6Ysxh6z5rH1QJBA0xr6TUzfg
uPDV7Fbr/xXm1M8EhyAQpowV58x67NqfRIHabMFgUwCs6freMAkDxUakryrhSldw
eg1oQ0EMDLejRSYw1YwbMkUr0DqIKXXdjJ+G7NAhfAqomYNnu39I4blLmMI/dlsi
MriXGBe1lk6/k6+e8HMqknRf10389gNRitH5UzMHkxXffjlHoRAK3h9ejXXyy56F
UT7SftxtGFAQDE5av8ckrT6LXbVCPg/QJ1KqebhhGO4=
`protect END_PROTECTED
