`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIlYj2IHPB9rEnpCvqKz/rAHo7pRzVYvka315FO4Gv4o
i1107lHSmFnVTN4Xh+aIbDjMgHlEx2Grmrfi3kmqMsmWP8npC74NxqB56gZlJlXo
UGmwaDo6MNUrz+hGh21ERn3hKAhmjvepVCX2A0n4/2c+98zmqezoX6fRYIpCLkH9
OEzGjE/JfPaIDDC1Q9yBBw==
`protect END_PROTECTED
