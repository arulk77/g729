`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNey+k5J2AKS7J6PsQQSPUsV28w8GA6pMgWeBJJcjXur
MCTeNMGREM0mItFpSFlhXfFn8cSJXe3hey+LqJE4tHeEjkxiq272/KWUfnU4HkWE
P0cnKNtIjF4elFhfQNaXB/8YPas0mzpRGY9cIR2mCht2gyUwzYo+INIVYYm1jiHQ
0ZVlZIlJtftFXgNoUlvVKvvtBVr5FDCVfXcFsHBmVzEs9EzhG9B9mFiuzuwJ15KJ
8eGPcxTtFDAuYQye2TACWDsRVvtHZmjbSTgw/cGlkDN1kni122XD8o0RCRiHMlSA
vgmITz3KYM6gbNlnxLT7izS2rGpUHaBDxyuckdeaa/2x8UGteZUiTAh6hdcsrN1v
D6XcIpqiunuv+XE4z90+X4tiBhwILYZLthWn/XZs5MEozsXvO1o4bheu+/LzVyos
atJK1ywciEFyajwwQm5lnh4QqsW/MB8qIHepTkdMppR8iKkfsUSt2XI1uXESAerA
AK91kyR9Zbf2x+XsGve20BE4jDV2U85k2/tUHFHk3A83l1FR7FdDdy2TqatjQkhS
GYiEywqJcpuFX1ZkaxvuG/xvfJjAjCF3Ru4w1Gj6gOe2ABDYnNwnGieoEOp6ySll
DSdMtxLZ5l14kJd+WBFVb83q55djVCoePopJv1jiafdWhbAmDaFnqAfEWFma1/B/
`protect END_PROTECTED
