`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL80PCpsrXNiNYqXt6ehhEH4rcP9prFAyI8+pSCb3xdd
LfNE7+u/vsMno4xyL6SXbz17CAFryp5YGDkcESnhAR8h6hCd2yA8yFFvZuhiBEXE
ssiRWp2vL1swmHfufzgVNW1oVa7DxuuD8q1ilDgS9AD/i03Rc8T/hBJgXlvEH8Qh
KUupgptTc9ixIb7eDV4hsA==
`protect END_PROTECTED
