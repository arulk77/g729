`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAQE2SyCpJggxmltBQneNQoiaFjpBX3GTkXnveYKyJ6F5
GAhSfDSapT+Zj1rUg8Fij879RugMBe33j/jJCn893IovxGPk6N2OCyFAX3/6zVUD
dhTE9+6Ez9b+UgE42z1gNeEyZew0x2PIEJ6+FRDALXsbmCPPeBjh4tnncMosoVCt
uS0sqbdStEhUD1fB0BqidLgi4TZZKjmB+yXONPR0EM5Q7pLK0ytC0nPI/JAjC0VD
JpTXZdcZOjXWpLh2c+6rYz8AoxBa0aYrbW4UaB3NaIUSZbnWNp/YIjZKa5xzk7hk
xLB34K36phRiaA7KphGv6mAfZofhjbXd+CtQL7j8rNTwL+Piyx8tMt7mimkr4XDa
nG5gAjseEU1uDW8In1NfBCsQbIK7labYvcXaJRUT1Ou/xD/WiIPiRahfyPNCnmzP
S8HiqEskYTcAKwEaHV/0IRYKstnIKFcKaFYq/dXA8MSaT880ps+UrKngUHYBuN+9
ysXbW+PysI75120AiYY/kr9ciiTht5XqT7O/F79yqb4NwHLRn9QT/qG1qtVnIwtK
aKn5U+dMlvCo0JDx8NnRrl3QJFQF2HvdNuIXhzq5lXDV6/iT4441WCLWrglun3OH
TFH/V5qbAGP2I/Af6c2QCOyGI0tsrRuJn3OEQxeMnKowa0iXwhfmkCZCjo6LjOuO
SRTK21YtMoJyUweU0LBX0O5l4yfca4rFqjsxVZkSJfNtcpVk2/Orwiv3mFG3gYHe
m0jy31uKzblQAykxs9o4GyQhA9vBfGVUO9o1afc7rzYjnTh1zeLC/f5hcdJSSccg
FbJTV+eK76GYNJrQ8+kXLfx7IZW76y7eNHzFk8L4KBmxS7NrlZiA5yn5PJTL4wqf
tF/ZDevv9w2qhsUKAieOD//o0IBEvUrf4sYxoIw8odwLCtPAWhZEIyhcqJMDwdc9
FXxrhazEAWynsrUGSQafZngyfpFF4vvk+IC5KXCywy7siDKdAaiTgSK2NgSIwIOh
nk7v1KFvj4bkJX7xC/bOSf3BZOZoexr4VJGe5pkfC2rclSOO2zOqJmSbYoPw3ZZb
OKINWg9wn54Qqg77wwJQrSD9TsrQf3CBIk7Kdn6TmzGcLpTDxZBzcrhFCDN+cfsk
M+kRNMMYjAFEFwCO79IGYcgjXJTNiTd7HhRKimtRK+rmGM7qOQ4T4+a7IXSd1cQN
akhHmgc4yvDZFjjSezpzW88lWF8leQ1btrwITHphmUXA3eAFxc8pdGQvxU9tMsYi
QT/gPCUmKJyQNFwUTyhOYDAl98M2Lp/Ygp48Q4nt8+s1x1QHKlKeBspP0BGpHCHV
VpbhmL4Y2PNBIw/qLebStj/iq68Duo+HNzvV2jR3pE/QErFUmlrsZ5wY6eoAoIU1
uaRyZsmbO/KeWFI1mRzeFLA34WJbf8Q/jzFAvZ4Qv2vf3yvgKPZxOD3+akCbKmA9
naC9G5dlA+fUID5ZTiriXWG2uEAi3eaci0g0gS00ScLBblKJUmGKc8XtkTZlrIOC
1ocNy+5dG5q7SYuXzz9I0pREDpF8kczjGXRTpDdDQew=
`protect END_PROTECTED
