`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKI7ONUBzv8PFWuRXya4NrhU/W1HkdeURnB+/CIIUDBW
cxHmbBcZ9aBoACMMdKsYSQ4hSPnRgPyHxT/O41TSmhZJ1BE8+WhxR5KIORpPBEa1
IRgv24Tz4UrhNSV/TJxajQ+OpMSc2zIga+5/ajD/g0iDcn4Dkv76BaVra1VcWf06
JtYvYnMzzSVpZQtYAmUb66Yy9sHS4J22jYIFoJSVUi6gbRpEwvuagXdh0ConGLe8
ohEr3MxINyhPdW8GYH+h4txlWFZmN3pcp66g/VtPM53hDS5JrPmRSSVjxwYVL0sK
4ZSo0ZkPJE5BevsdLEYC7w==
`protect END_PROTECTED
