`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIaq7IlYJqhnjQubtW0lfvz7BBjxhxr7nloTI9TQh0HP
aC8PojVi5abdKNwMe6d5lk+F8n9HtrP8Xxlbhi5OR8+zaophB1+Egjx1zhIogjL+
VxK/zasBmKM97ohDvGtgbTfBfnJZIlNDYigwNjntFiP4IpCFp3HErwbNoxvnjtwQ
ScpfwLbm+6EtNj1PcQuNSDDWlQlFroyravr0Xrfe+7vuw54qMtFJfjlqNPJD4rO5
GftqvLLdR2N7ewMNbaL+ZOCvuO+kKLCcqJzez/9j5K6rYSTV6re0Nge/lrSj1VKc
qhuPJoTLB+n3ZCxXQ3KLNuRhMynbSsN4xOvV69fSg8Uad27txm4a2L3XKmtBIZ//
0PAxMt5d4gUddie7awA8BXUUHgwIj13y68GrlBJJufiKS42+k3KLbIz3chgxquB0
DuMZvpSLVrryR4XEvHXqXvuNQEyuwq3iaF8bqBfokEwTONZ4po6aZAzfpkah2sLe
rJzP8y4QMcmFlNPLJwajmoNZrNAqKhdyYK2JJ3uV3ZHGaG9GeOqHD2UiEADaGSxU
eYzrQ0HWMktlfuNIBxoakA==
`protect END_PROTECTED
