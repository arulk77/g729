`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49StAEY6pxq010jS7jcUmUB9g0wUBPZzjqVCKmwExqrb
0UDCAxsHyRvKF7dY8UIStRuXXJCYF8jlULXa9PFad7XOb0XsTMkS2w3+SHXglWoh
NnMoKnVvhZSYiLVRZJxNrgMBXw9QeSgRbb2y5yOHeZ+tYD9DH6oJ+Y0nUo/YvmHI
UWSOa7ilVmbd3LnWtwxJ1IrFiczduqPnrM13hzLt5tXVTdUasyjEpcuI+PZXml/I
4aoZk78TMKh2z/+kY92CwecrGjCDE+2YvcRxAuOu+CAy/tX2dZnDdJce31T7q4l7
EgForhYiw+KWQpfdbNyx8uzz9qU8USefST3Iwxu6bGIBuU/PkNgnjpcoMtaSWn78
f14AfGyFPIzMBEnuFyTdUtaNJuK0mB/c5T53tO42WcQ6HZ4fSQe62HRQ3iW/E5sg
t56DCCE+joroJb9qBF0IFotdRJwUKF/7yElr5YZd2LXu9T+UoZ8ObhFiWxcItU8Q
`protect END_PROTECTED
