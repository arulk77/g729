`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIhyVUqhH4fpQ+/RUYMGI+03MhxzvMs8Z3gSIwhcxzMu
0TK/7d5u977blcEePtS0KyuyBUKShToUzUdZH8DcqtHsgV3kA7eD4ZEGPJEkFCNl
B+W9t6WQgpUr5armZplJPpejBoE7vsaoXnBrr0UqOfgraAzL6pXVrA3AOrLZB8FN
FOoldtKK3hki74VceqcTU+PBncdyivfdHWQrTrM/XBzngWH7TYA7qLrE5RPx1Yyb
qJnOB3sjOEtwaPSJePkVtqAxqS7u2+v69HNKfkHvTzsJbnUZ/I8BCZjHeDbdpcuy
YY0kuqcTgdhEFssid35GLM/XlnlCXk2ub53pHWnNIuu/vmTbNbrnDWCEqUSj0hVy
GY3y2+oYFbGt4Z0LZzbM2g==
`protect END_PROTECTED
