`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGjcDlgioLvNNpQYk6P69htQLCWQjoQoCCJuTQqalxxj
Gi7l42LiANkj65nf7hucYxK4FuOxjaftQGoy508GKP8C/6MuOD5d0gDNc360ZXFr
1h5S3pJguDdn4Bwd/efwNWKVBignELC37k4OBmJpfOBXwjKSBjg6W9TdWT+2nYms
nnr1lGZwSPj/hNJ71ZfzKkiTZ25RzNhhatrp1pVV6s1cwHcLeIoocGKMEcX4ltyK
`protect END_PROTECTED
