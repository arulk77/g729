`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
36A/U5tO69wVl401zVMLLShKh5c08ynbctNtEGBvLv/100B9t/m7ZU3RlfgTMgtx
i99ZjzTcBWixEG0PkDMHt6OQXTMPe+0wOwFg9EzZnKy9YRMixLZZgBCTmvO5qD4u
JlMJ3Rh8ATE6bmxAw1STgqoKYd5u/5DJokbx+zqgufiCGwmqqOm7x4xmEmvrSODz
akIgUsuSNyq7q54YaI0qNjQc09Lz0wUDtg4Ma5TNrnhmdz1PUInBWu1SfNCdhkmu
5FqvzSoFEIc0rveRhek9+blp1P0cbcT9xeryZUAVP9wKlKKmS1ATTAz48p87RnfT
KS4AfeqelZgjkx78bmKbufkqQUcyi/yca1SE1WsO1bfOB4J59MxHuog7erTkyhmh
`protect END_PROTECTED
