`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xEP4ysk9HqDpr0Dsp/lKRqBEdNPao81jHFbhobX8HeD
3NS5/qTrO/yk1QvETpYz4tAAJXAR4HHD7/oDLXHQEJ/Zxy8JnR77YouHmu6Kxo3J
HuRR/wm+I6QWa7cL//eNAO98fYEqBiROlnPPySxQNYPxtXn24iY3q0cQW1114y68
ItiKuXMuzo+r6swEZjPIa3349o2IFnsDSshjF2k+X19S5QlViuwSxN+b0sJcuWUG
XopktSbKX+8m5O/+4xHaD5XaiyPb8azoLv7Z7asJaz8=
`protect END_PROTECTED
