`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFgKYr8eIdlla5Ir4g2k1yuszLDODsVj+z9aLvlZ3dba
tT1ebrzjG3yOH1Bw6Z2PyjAgMBLi4U5wIll0nBXE3QXMQkxHfuYm/lSjQat1/Jnv
QB6btNjKHarhfGtNqnO7JrFY8Et/zbww7j2vxcS8+XI3ji8IwWIBI705jvPFjkxY
rfrb9cx2Aid/ppGToIRDlg==
`protect END_PROTECTED
