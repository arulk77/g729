`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEx9gQoErkA+kOa/7cgcX95Fh0R7rQr3F9PdbnNGnu2i
ZaGuZzJxb6ZoYIRheTPmettejjUtUsUuKgBn8/CB/TcHMWIDAvUQTqVQzCo9mnBr
jNt81AUpaAji//gwLSqKX5RQaVvv3TGC/PcDpbxVTiPW8+gQ2CQmMBSue1nmvhxB
rnRd4kT3OvL9iL9bsGkhK1GhhYQ8Uq0txTNeVF0QmpVWWq+Re16EhHVjmmpTXq5/
1UXND39AXdGbN79aPjnngzXiMXuu7XyJ8+2LBDfUIH7veN0uIDMluorzLNkPJXum
xvwWKh0AARlN5f7+Q547eUhMvtQvGqdYbS9KiV6EzEJnPyVvwiOIUfc8DvILjxFP
jEM0NLzubonnrx37/6IbhHc4b5X032hEK3RV2e39RA9waKkp1SEpLS61R2etk/fL
9mMS4Qoz5YHqWYnZq14/QfRy53Q8rU2V5nOGiqIVQuXws/KeIKxH/bCn46p1yMnR
8qOcaae0oZnW8gzxLMMp9AMRtcNtmc1yEBJAP8sMMWBcIjnQnShvxzW4gkWtMdVb
`protect END_PROTECTED
