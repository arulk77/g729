`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDxWp8EUZOvC0+Pj4L+w2kOq1EYqbv51joN7ilgDbXTW
tbJrfnL0zeZGwOVPcxYVTWImTKnGPhcBdxA+A4xgRFYxyehfnnyzJBXkJteMurlJ
JboiEoZk6tDksXzNN7+ll2PefKYKxe3qNypHFFDmMaDKwzVl/X7Sssoo/J3gy7Dy
GB0HxvSmMzvWny4WsP8dOSce+kvBG5YVRmnLrahSgz5Xgh1//RwXilZdKWaEO9Ik
PjHrZn0U5bLp9eS+Ht2xU8RvfTJ0kt9suxdkR0vCJ2RdJEYptxtVz9kdbh07zz5s
`protect END_PROTECTED
