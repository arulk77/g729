`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCe90E0V5knUUKbn9JVmRBv8mi4YVWPEBhNR2O1P3IG7
8iALw2MQSKnbQv4tYvmgitPGsn8RSd2OBlU9Rswu7Ybzy2No9+zAnzl9Yo3UgfJV
uNAyyxLLXZZE5OiQdNLix3MxknA1qeQ5cOfQPtiIjZvunYguPTBIhreyIC8Jh3Gx
SUAkhLJSX5gi2/9jNIbx6Z+yREbZicggng3beBizvBe9xh5fKvzW9sHqfx0ffFaP
NS02l/LIs+HOkvzP/P6iAxQhim4ZzaRJuIyYoqUX0D2N7y3+J7TYkc7eQR/N/m3t
JteA68twOE8U/M+B+M8dzl+r/KMm8kFCNSx9yEtg1x/S2GenizQFh5N4+ZcMMMTO
7GzQCbUF9FOkTXSUq7yHlw==
`protect END_PROTECTED
