`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHwZQ5YAIVXUkAnOCx42fCCAvGmMGD0Br4i6S8GldLWy
tPLTdldkKDjXN04JUzlOEIRlB58oYohyTgPj1e8RHyE769s4M4wZkSZR7nzlgf6e
4ZPPDe/6ZcZXQRl6ou8+I4l+8ya7xWBReP8KkzrVB3srevcO0IL9SNR3GyEVntW9
JKgo+hdNe1Z9ptx7WK1IttaHLe7ToYC5/siBDqGqeO185qowPbtzbggAy/SNhhu4
`protect END_PROTECTED
