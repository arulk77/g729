`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAFbYAf+vJUDOxsWlXzhCWPQvAg56uxw0Nluy3zbjBF9
ycxzGh0hNMNItVONrdxpYcy2RYJhCVJqoRZgFe51zYTW1IdmyF9Fg6O99Sq6Y52t
yNAFKqjQr2AitYRfhj7M+ILK0Rc07lfaJ43ODp0B9PcAqd25gzwya0iDRGHqnOzz
fngSeGOIINE10DUN/59mMA==
`protect END_PROTECTED
