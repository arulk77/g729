`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44GTJcvaHNPHgfDPGnc9q32Xtm9kZ0QVlz58K2DDQCaG
3l4/nyXdIamAwwD5E0yLD9hOuZt6eCG+9DmchRVy1CAww60iQBxtNo0/HJ1Zb3OT
4lxem55Gz+HV6DiWg2dS+1e8InGBhckE6tjDMojhH3kk2jQ9BKH+DxSLDRdw40Gv
ubNd4HZp2H+W93R9PA5lObJs4wzMMozpF2hNM8CK9/sVTQgeLzR/kyex6WpfXdO0
lIlHQ3F2bSmuRsJW2n2Ibho0eco1D9J1b1PdjB++ClwYNdK4Pru98SkpUvGRTN6e
sFCqNOYdBjs+iTLIZIRGgw==
`protect END_PROTECTED
