`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEA/ffYjZY/T85FvHvAouyfxv88TkfyYrqckP7N8+1n/
MsFK4josRlKpwKaSevQzaPC2P4xb4HAoPNC24SRjhtd2hbiBi+sbu6JBZljV6CeK
6D/LAZ847pC8cDy6nh6tuWd/74A4z/OIyW/Kzmf/J6q7DoLiwOHP7ySNcV75kbgy
Uq0mww6N4JBcGJ9cD/KWKcKo7vTyRVY2ciFhLtyyH8QM6VEgUMTZ2CleIMNghz8O
PkavuLvxfrBW2eBWDdmNpPB0gk5kn2E8G4CTwKtP5ihJWdZ7ZPM6RgyMp0qWiaej
ABg2yXYTEWy98nlYYmOb3eIyw+M8QC7DQQF5bWdUhzqcxksTu2NGzvJK8IKnZMv2
GOrPLmOq+JLy0hrPChhphg==
`protect END_PROTECTED
