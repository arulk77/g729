`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOZjAeID/RTAvnJ1qVnICenMGlBbXZWsmyMXUnWgtLlJ
wJoOIJQGQXb2Mdz1PtUFx3g/XdRuYODA1QDI5zVuBLDaNoxghKZuG+EEwwZEk9/D
IlzRLixJXGoqtaMJ+lzjEJzTQNnX2lswg96K20ewUhCz3kjoVv+lIODT/APOITum
iqCRSMoWq+/+KWWQz1Zk49TFQ7x+jv6RJXZ32nJMAvCbBONTCD5xwyDbWxjhJUK3
`protect END_PROTECTED
