`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
gy7HdhRacIemSFionrLM4e+dMxHj2h/o6qWaopnf+CA/J5Cm4iSWPXJptmVYrDQn
djYfotjxrYJaRQz+Br8OwvuJhyhC5s824yj5jUN+wGDUXEve2iDu3wsvmDt5Yymk
Z+UP7SmvgEV3drt9474ryVIvh8nr1M5L1mlDy4FVKvBd3lOswu1n9VwKs3CNKm6+
71SQpT9JRUNX+nECT/658BWkJRnBlsr703KKq/JIU8FG0sdP9UYJD75y/4ipNaJ9
OsBsdfxc6ieNnqmfqjK/TZOgWoQuu/+W12AiEdk20+w=
`protect END_PROTECTED
