`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
xTgi/qkZVQx/vAaTq443pSOFJ1koeHQTWb5Iw83dEUtC1A31OmdNwxbwKHX+sVk0
Qqz1qTlWO1Kb3aR12jD0vEeAhFvcRgqrcpp7/5w3En7/9o8RWvgI+MeZfj7gCK20
hOhE2uhWZGEpiiOl01+bGVPBAwYTHkN8HZpx13rMpBZ8KfTRiAfLvzfuM76bVICV
i4eiK4jo35ZNtbmi5tPA3TpiHqfdRzGPHjkyuaOcKf6Rbf7G2fTwLJSZJCYzUwzW
uUll7njLivitUbCbynFNE8eqEQozM1MxllsrKrTQPOyRU9ohreuOIjmcDsrBRbmv
JPM3gTDuzTejvoU8Kivlkg==
`protect END_PROTECTED
