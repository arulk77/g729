`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
76sFkWaWtW2g4TUTKwVVqoZyLN7GvTWjWeTsC+/zBo/kCgchzKsuMOleFjdKf9rj
X9Dt4EumWxZlM6HwWVKJtcndo25pWdPerOcvdgaP8fq6ahJzC+D01pxI6NNMgmcn
8vgfDlS8Dha5tv+aSZQav9DoVPgqlltT1+ncDLgiwwvNR99/sDPW735S0v4U4aKN
GmSF17tTKVtmifmwIpyAAxjT021Cuwn5MY71hZhfqr1StYWZcLCa7HzW6cSfUjDF
ad6MGHlip/7itZEq7e1GQjz0vWlaiROgIEfqUz1IyZO48NERq29SS/wd3ko5Gy5H
m4h08bSIStmaLakjgG94IlUMyus9bZPhuc6MuPSQQcw+8dfKsw2qfMmN/jax1oGy
XaRfvhQoZ0E6HgcbP6FydGUW+nGk2JQOI0yQCU3FU6AAcDbBiYEn5/vWHm6fT36V
2sottAMzV5E30hkhLlYo//nbsMP0rqua6y7WLVyBarQ=
`protect END_PROTECTED
