`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
cGNdncqj3qygDGZyEZ0wFr397m50DKsXulKY3jrsyuGx0WElOROLka4u3R+5hZ1F
Z77WQ45mL402Vf2CnHT5j2TKFqkCTob9gF5D0cgiK5Rc4J6aNHEXskTGdlBUjFyV
7dDsctfVkdRgNwRwYdzwPNdv42CVZEKm3zRnunpiMFz5lC/i+boUFFyHiBM8wOgV
+Eba5QOviTTK/oQTVe3nVaTEyIhceSPMFq6uLUKD7J/tuKtjZbzQ4Nb4kpAZmJ/H
E4nGMpg9b1KUJeL6vX2itRs9txxne8hjTpHCIpyDTic=
`protect END_PROTECTED
