`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJzABYeb2BwENKNYZbicFbdxXrTRuIwANCogEq/RvZG5
Hoiaj6s7+LMXH5am3pSb7a1L7e1x15CBcKRD8Ara6OnSvlsXXotMSpNjwWJH0KhK
WiVqvBPGjCtSWizXuFeaYIn2jZ2RWIfJAcAUko0Zxy2eicZEmJATd2FXe+VVeXxS
HVT9SQE/ZvJHsH/3C71BBDydrHLo045aCECUI4IW5tMBEeAjvMmvSzbbqKtqKZmb
zfhCWByEl2zGtoaS2yShe0MbFso7cOEhl4EevjXuPD5vjFBkWQcgSf8B7hX5jXwM
y20CyoV/u/K00FSOaEKbq5Fdxmx+GhMVdxTQeI+FYczZzhNuJOX1041qAutL7dn3
`protect END_PROTECTED
