`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMy3Xm1Kp3faMD6+jB+0nKbXbajQMQpeX1edcm8HIc33
GuLk5fXi6e7v8V9+ohIJFWD8O1JEYMZaKQk0/PPp6lHI/7BojUZ+eVjISlOlvFG5
YS192WmGlHQuOd8u9HL498bC5hJ/iEEOA9qGhpC/1UJ1ekEBqpypvVPOPpIh+csi
DReljGDVuvqtaaKV2w35EM4yT9v3kGyuxWNphAK569EX5bvchgj1YO+BkH43eECM
EnQB6zCXNtR23w1P9wKr+TKnDyLi7FzHxPHFaHdd1V2lO36wB4WhjOJxIa1rBC69
0u/A3DIh/Htu7BvPRpxO8Q==
`protect END_PROTECTED
