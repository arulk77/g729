`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEFyrhwYWYS97GuDd8PqS7IPp9yDqODwIQeoHdE95IBd
gzjuf5ih3lstEVHCR/BoqBQO3HjhZC0fViRPbCwqU2JvRCg7OKSC9axdKIf7oDj3
VLIlgeBF0CG1BIb3lrhaEuF8WEuyIH9lcOdfGthZMnlPnzGbgkmVTve8xxNFKjbX
Lhlr42Tf0CwfgrkKEoXLamoMpK4zLZNj6mFdlNVItNLXqfPQjHWTIoFy0NKSLMZ3
fNZ4oiY/5BII1NdIT3kp/FZWSrUoUApyf2k/0KanBOG3IVt2eAjk6c5tn2r8hZpd
hg5zJDdgpOx7218tPdc9JuLPbpKr8Oe+rg9KpjbzCU3qeXcX4lLw/PStVDEQUI+j
S9rpwLO/w3ml0h1JI6eaA0CtPntYhq/Ss/V8+se0gx4bv2n/RFE89yAEpsNhAN0B
NwNwBWrRiZOGTeqUzwf19KmMGAhdyky3pN7jr3LdvjoJznbpIhuUzfpfuIWXv3kz
A+JBskcqGwmgjiodSwL23XqDp9P3WMvOICs56luCUgL07QZ7ay9sWw0xR9oiLl0h
`protect END_PROTECTED
