`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4y5hZaiiexCDH81mVUtQl58u2bcQrMz6ZuCUy54GiJcl
yXijIVxjbVSHh+2xoL2JciTkV4r+LFKsyaUOCqRZUXan2b4L6q8G/4h9MeoPIwZH
ZCsIKanzgr4uEqthhDQsC6rMSOhN4AQ8glCBh/74/dUz8yfkB/dozoE3jb2J0CK7
moOtImXwg2If1/5Hj604LtLvhzYlgqrD/D1yurX6hLI=
`protect END_PROTECTED
