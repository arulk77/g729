`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN6vQLbgcxatbsg7H8FfzuuzyNt/MLE+aIlE1TxOM4go
egEGCvl8BbdT1hbdZbRnVf+Td8gZ6JlnPiA/H9S1BZ1hiDxQkn9mWY3nGXxtKYky
/o5Hn2I6b4oezAktU6c810s12xNMIJlecp6QTRETtkvUfpwqahOlZFe9PNaKRRdN
HsE+7SMEWtu/IPhzwvSAXrhV6hN2a7JVTW44+/T7aR5gfT6t1JzqZD7DXish1Z42
b8O0k6pR1KWq08uIZrVRUOx3JJz/5djlFu4uU8uw2Rb0ZutXiE5O9RoyKiN1V8CA
Y6F+17/3L+HaMfx72j68nNXxMXhc9jqE9hTjgYmAKG16aHN34XZHiiJDfBwRYr+i
qjiRilPgX3Ldlpkrx3RkEUAoJYSdObQhJevXmJTlLPG0so5myXXDoWEq5J1AtMiI
aIo5chHOaDWm5r8ODn8l9Ow38m5XjAZNJ3sgTyqEMK0VkJrCVmoJdo4058p5v7yn
9c/hUbEWBt2EV9aZ2+Al4wwRlnJ58Vqmw3QGU0Bifqu3Naf8tTYg/rJeKG3HNGXV
zcnfUAx8GWIwwd3RN+rlFQ==
`protect END_PROTECTED
