`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
sJ1Xie3bhD4eTkc9Vjah1hVUsamEx6ZKVVTMzsdBXDUuAXSD/y6MIyk1rLnxijX/
4oub0Ipq0NgvPhuOhKOIsExlXqa8Zpu9Bp5aUkPjgYIpN4ApviIpWzh9bVVhxCS+
MLt4VGilpITHc+FPmS2KodvV8TPU8NsliFjr3u6xH+b5mLZfqK9n0klWvekvJw2m
NGpEJ9E6rcQAachf++m3sxqUbhw8XgK3Y4TP93lrbZX2MyMD/POAvXTOlgtTCsuQ
Dq4J/0sguTzQbfggBIPqiksH5Im0GWovSk3Er6Vd89H3F/DBjgZjBaMdMlnQ9kFq
GhtK/id5neeDJLfX0vxraZlhB0+qLNn6NTJKr2OOkODi6b9FkhaZaJIsH+gjJ98R
MiBPbeuMiAOOEwsKs+LI/LoFBrY56uhQYIjwfTmgLZe14Y4bWVXRaRo3hTxdDcJr
0cT6NQyEXtfaUJmZr5uE6IT5AIllpKfB74jrssp0MT0pK3c+SGIpVfFyza14pCKl
bUO2MNxlt+JKcuguzuBSU1pJKPYqaB0DW++UTfj3P2nsWMcVv9XD9qgEP6sW6Ef+
KAhNZuJ6S2w3Dt/MbOiMKngALqnc+7dMq8IfTjtUydQ=
`protect END_PROTECTED
