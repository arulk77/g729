`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
nT/SH/82Lra+X4Jy/BV0DifVDVg2f4qA0lGJ1jSa8FPzJ6pCDWDwtDaERenq6e1N
UG1oXwWXl5t/sZtE9BehSBSjU6Y47K/Y5GDFo02bRoX3a2KURzM6Y6UthMnXJk+z
LgRJQdoRabMzoo2A47OFNTS3A8tb3Q9bxfaLjfyOUiOe7+UjAga3kzjxAhxwI+Di
dsrYyRRfoFKQfHDs+pIoxxJQ1CwVVMnXZK+0axZj+yuJ5m2Ieu0AwiUIowGREUQE
ZwrKvM842cHVvnY5oNoefq078LxXAUxcgX+HBlabsVo=
`protect END_PROTECTED
