`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4ww7XN5yzDz0mht6J5Tj3rv1/r5ffuIChLWciKUeuBsG
i2kjmmxcKDUTKu3jGl0OgtgMi2Eb3CvYSfPCZihM/IynZSo/gGVhAI89brNZSg0q
4owrXgybIaJphER3SLPeQUIYHe9CZ/DjH67TiZMM4nw=
`protect END_PROTECTED
