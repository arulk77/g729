`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+/Jy4TwlOtoMndl4OvxqWx1y46cpcB0jSDxFmuSfnFb
6i44IwHbNkn9FwrjLpEvwfYU2ZOeZ0I6fGq+Of54VD9zlQeYmkNuGtk/Km7IpOvs
m1pGZ9fIbIVgrj/3qYuR4yUXQDA1SchbdM0HQOmXwzj5IE/UaOOwkZrQoMCWzzIw
i/yYHEc9NOU7ENnzZ3RbkhCwRZg9YZjQZOVx+yiYWlGBSyNsb5rz4YEHSu6RHBn9
OJtSnc1juVAaRTLDtCrz4ekmxbzyq21pGA/FZfKRUklRyEi7RLabU5fKFl5VnF6U
dD0p4fY8CTSomtzKMcrahxXXlEr3j8P074DXy7ifD++WzDaV8Xxum6UrboIkI94U
4DlZptHgw8yf6QGnHfEvbDLV6N7eZt9KbAPhZ8zmNiikqkKwGf2yC+6rI81SjAyX
buVCOgG0k4BYYGN9ldOmt0Pe4/7+iSL6DM/pkM9PcJg9FqMFtD/VFn6p83TmGv7S
`protect END_PROTECTED
