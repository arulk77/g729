`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
XrTlrloF3cVJXvKrO9HUCZbpe6K5tItQpQA7DpojUqadSY+9K+hRxHpxzm/3mHH4
MxC6+Kj+iuJbIdi/jtswnRHCuuyZ3E0QCAS4ENH5ctoRt3vXZMHy6mlLXKkcnuxY
pOYNpWG9NSndPIXa3crYpjeTrb5dLVeC/dwWcpOL94NLHFQqN50QDT8d4etpG4bc
8oCYaSaDIfFKZpXL7wF/ktgrjwYXykRMK/LdvmoXfDNcdpDwNekUI81IJP3z1K3r
xPLd5J3ajxqOnUTXqwjrrup4tmIdeVEMhSUf7va0or3azp6fyq2yuiB9rA3XfG7o
PuWMh1kryujBI3uiT4QqN20UVJ1d1jNLVvLDUHl8hitvBHEzV1PIpoX2E3XG1L5w
OxEsN8J9sTjB0D7f/Bla1aKh3fPXCwb9n2VbEtqWLwknmZWuKFsph8H4klSG5cdv
Ld0jqwCe15YZHx2j6tDXkIglgV7mfaxOVC06C2416E+1VX9lKTlHHppUiDVVTP4n
IDa2wpQwonsVmvKdnJ9RucoGdxTCpDvkXD8RzrnKEKvOhQ8G3JOTQ3WaqxqwXb83
cKGziW/ZBgYuKjF66bew/g==
`protect END_PROTECTED
