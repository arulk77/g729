`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
eX7eXjdMg2n8zf+K9Hhsc25SEMm6T/mUrZu6k+gOHj+GCleg5ps5f34TccOgA0pl
6ZllfQGYmE45fgfLKY67VLkiSDWFYvVKQzbKalRmapnjMPQcm/tDfCVo41MfzzFT
qLcEn5HiwZ2rN4Wys/0JOKr9EZ4koKICruheyUik6Bk2BABqsan85XCwTt+lISVM
q1MMnlSZjLV5713yw2Y4pPf7t6c5HRZBLM/MMAJ6B0FgpET8OqHmWxy6jC5Ztu+V
fgzQyGauF3/5MGFi+vUeWT6Vy61Jn0mBj9qJIBXEYSMjIvGFO65J77vYdwMNZE8o
5TJcetu2/47CUe4pngrxb7oE7mvDRg511+vH238IB/2lw34O1cIPdnVeqpXOR6I0
6cYFODE2TjbVFoducsp6lpqoO9vV9ne8Y4D4uvet09zmnul4HjbwTrLC2ek2Ey4E
JAM07B8xSdjPaiYD9TKIPYoMwXhvTSf3YpOiBCP39FgF5cxff6fftA4c3eDUddAJ
`protect END_PROTECTED
