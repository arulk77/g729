`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGHQ8j5zpBV00pctMbRMmRmp1V2audk7x+4UUSfGFP4d
v/V1iuWEVBUTXmfx2/f90KJN199staA2EMuWqE3hOJIoWzM+QOEAlMkQeuq6C66Z
8geDWbj9QNCkaSbUhM3vCR6INmx9vxpGqcn7nI0hd9SP+nUstBo/7xdVAmQaUOgE
g943XPHzKcAxTZvoheeDL3IxagtJ2hG2wBUFJlqzk5kIVkS3bTPPK8OuoCUnpuP6
yGRo9eOWf4adHukQS3FOhHW06McNQtgEZqSI9PL+WUKMw51wiuOqG81cUSdSdu/T
fjZjMfMcCD8YXOrSG8HAOHlPKwQRPWkfMweBSpMGngVb5z9bqQIFCzkJwVZ9a6gD
liRm/bTHnjsi3uWv6CCFy06ggUsHfOdHSTQjENfohlJiokF2liAATJv/2M9M4bOF
`protect END_PROTECTED
