`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIjiBmhEUVYlNqrt58f7gdHm+y7yRmaP2tNLVPSl0K3z
rmFdXdWwppkfNDPgspdhhYE6639JbdDh/lsuvW7UaNfV6yzoCE/0oOEtEvsehIQg
RFgzVlXF0Zy2xEsmbvJwLNa/d3bH6TnryUgapgwMIHS4+TPOeYyPvt4l2J4zykph
0hTl7CjUBB6hxlE514lKDqMhzCpJ4LfGTEnhGd7Jmm62EH6RLcedf6X8657f4Img
`protect END_PROTECTED
