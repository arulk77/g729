`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C8x2eiWqm2vW6MjY6483rY4RrZg0ceFtWHQI4Jc4a2pa
nfCYHFMV8yAG5IrS4x4bTyCpt77xkbYHL4K7I5Wzt0YjYF2gRCeTyNjI36Dffr5M
ezq6IX3XM+Qpg4AcT1Wa5W7EBXdVDpceg/hZrvFWcAI9a/Gs03/Pevl4HOnvVynx
YaPaK6ACFEgoZUAT4+z2r813XLvCuyFx5FCPwVBDZuQR2Z9ZUlWPIZC5bINuoB1x
sJSVower5tFEezxk5QXey77YBkP8hDHJtlApfroBbFlItJXgUSXqC5Eh3B+Qgi3P
jYjHqCyn8nfUfK9uYi6p8D3vBYqK4YVzOn73ZGhBFyE2Cgt+57UIN1vtsdUo+XIo
cVf0DaIZ2Lnp6pwjGDtVcw8vpYe5IK9pWYuRMZDYZINh1yjewnkiX+0lFIfGizRl
sThQ43h6JOw/y1/4390XB42ps2Jn/F1IT250UGMALDrPi7YOboSXh3Am9nHjG7dC
n73HgFRo/IMyJ/ghDwYkHXyJCta86Lm3Sc8UGUV7yFSDDYdWj8xjTb9CCwjvXLzU
pu7cnpj/zLVikEG3Oz/0KBKkyyrqcOYi3MdDLdQ1Vc02tRATilOnIF6V3lONuNhI
gvQO/HeocZde5pVHw+HLKa9qDPRE8EuGPkJPJ3hr/1lIdPMgVokZgSXEHCd+2rxp
9nGTPhINloO9WOvb/s4z60F6tnFNTi/iMsfcnpjtG1vS/YFQDIXoAPJaZYy/sMCs
STqmVk7y1flLk6i7oEZgZiUanY23xnX65//Fk9l4wxzwVi//s9E7zmZmaj7WWCj7
hCZuUukoBBfDY0qil4qS0CB+M4N7HyGp/EUWzxXU9rNHhFcUC/WlzQ5ICtBmbYov
rR93PSNaDf9aHozhha2uYr54gCd3xywS5X+BkZquZLlhT/rUbdgzk47r349Itacs
t5eUKHrvWZPHcM88FE4j/KUhyC7rwgyB2m3Fn/M91B/aQ+IpCEpPk2OYhhWGrg0d
/MmB8MDUBTBeLMDmzgJ6D2g/Hh4cC6vApRKb4fYkQgX35LvRICag8tR2THJHqQOW
Ltjh2/I5v+/vHcCE9zQDgUYQqgCBRGDVIjCsybne/KjBtMqxdoVEaOFQSYEmZcPz
4f8EzFptRYPTN1LHos9n9zwVVqzdvqFVmB9ICXQ3wMVmVDQUqbJkn+bYaivRKzEv
WimgTqQ0FokHGIPUb5NO2LkPIvEVjWku4QvMvTBDSIF817ZAtiu/HYaokvnYABcS
lZNOmXLjrnDyqDutIBSu4TkTPAyGMZ8DLryFYBfAWrdC+R3s0xNQ+BAzAdqFNHfU
f8x267rKwdyUaqVOKfKyVNtkNRDtAs6gYx8Pf511FQsjEY+1n7qv2y5IQWnidgUT
AaHtw+IypYnfzy37VAvmAIDgiNY/T5yki3IImRmQ1zCO3HEyl7djqBEDNiKBonks
aiJE/AEjj9WqQ9eGYnsU9W5BiFFaIy3HQXVk8GgJxIn3NBCipr9JW6fLN3rpjdwO
lB3Z1M58g70yJv5gHv0QSo7ZwVGDmj9ttyYgr6ErOiSrM33TN/tHrnCg3p44Hlyp
7X3y4/glHmRLSNSjsx+MPr67xlFF2u2QyjUE6q+JF2IrrSe5b0mON2NlG3ELXa6J
lRzGYnBA/iKwiU6mblzYCYpS4Cju6sYyI6oSQiWu4QInSTyWFH+KAVw7gpX6mf9y
ubA/8cjn/hxaHkqazd4SOKcWww1/SJjDtr4KAUt3DISlKzscKIJ+fYpro2pKuxIR
LBI3d0FxTwSYAwwrobz4z02BCofgzeFM958Fp3U/YWM9AuOANy3IMlTYjLLub7es
FBGKQQXFm9/+ThRL7lgUnL0DA+Frz+gLdwFu3NiCZOcE7CuNcT8faQeyIvslVKO5
YouXaGekNRBXXea4a52bchzfSZg+wGvKbj4OrNWnqkb12lRt7yS7HBiqy1JpcesC
JwnLd4DRRBVZ/ASTIcOqVCDoF+jQ7ldVA9U6lwodBNDhRQqtoeLAUipl266qSx4q
rzU/1igomUrp2gKiFx8wDfqHGZFugO0CA2vzEp5m6tUVul1lAvu81wdrVoRaY7Xl
/3OnTtV5FNmH8RC+lsPS2fMAVbWCRTi7y0eRpq5U7s1Mb+Q25M9ngG9EoDtmZC3w
hMQR2VCZGcWRB/8KYWu8aCMznDenMVsYAJDKUE/IG8MXNz9YpmBAk07ixeMLglcW
VGBveDKzxz59Amo2arrxanUyGjPQv2krS3qkyaS+co+6dy3xhHD7hqQ13bgOZMMB
sjzIgzvueFEpjrhOmKt5Z3D9VMwnJmKHxxW1iUvo2tyCE9eAbhaXPB/FCe9LotO+
R8gHg7+hji57eDIrhlSxglH+3bKb4vA1BivulgJCtddnLVSGBCH4/pATsi1QfOHh
PM3a9TivdFMSHYUK3Wgw/ezRgOOmdJuupI8WFj439b5fG3ePPRRjmwdXCQToM4Ml
mOAT66oDNCGMlKEinid6d7dYuFrWLK9G66w/s8TqtdkkC6JMlu/wz3kRJlu4C2cB
cUiNzyOqmzDAfwB9r5k+sMzRWREmCKrqi0gF0xqRP/hvO8Qeuze68WQeB+Xx7R5K
KWv+1a0mdmkMbUuiZNc9zBy7YvXJDz3kpemyfMz9Z1jE4FPQrbzURhQ3L4rLPDPr
TC0Japw6j6A+/2bb/r5ZlAs/kqmXso9f/kb5CcA0BAtB1nLZI1OuoPa9GdR5kv+k
6SJvmAJgS9BQkauT1nIzRSP5THnfx7ocCVqSI2Ou55iGM+/1/dYDu9rkIFNmLrvF
3Hj8rf6lSHZr742QsJy4RvH4DFKoMxBtTi6Fz3O2u2+Q1xsUb2zp4acajUkwiIwE
KBNW2PJZ/cFSViBmhKGVbsXRv/2KsGmjWpXFTMR1R1tR8ILzuQ1CKFA+bKVLAbNh
DVnhR5+ZgcTLphSV++KHtvpmi8GM6M97u9Msoo4ujDIhIhOWzaO+VzaY54iVYw8Z
oMycNhGNpxRUmT5UFkzi6YKtHafPcUYJddmGRbBLCkcYjlwh6FxQX8m6fDDdCP8l
HCJoHmZnXBqK59SOjBEjYWBzxvsgIb+TH4hbIvvL2jD7FiGNbc0lUMFz+SXx71X+
+XR3Y3rVNTz8xfY+kKUIQH4mJj2gkLjpphzknKZTKCvkzBxn7XVz3FqiMX9gmUnh
D7diUC0eYGno9T6VVyRy7B/gxmvSMY2ib23mJpvs0Pf90ogOVe0tcDx5qjTVNGG3
cUBEWWuxbq6nTZb8eTXQGWx8zFFnUidiIUhxD34fzEUnLYBxddWvyYv1DHP88IcS
5i1GiiFl4C8NcyyaGqzp5jUcSYo0MIKa779mHJvnL8Ii2BRRFoeiW9PqA9W/ZpPL
KCXyao3Tl3UYWuqS+eKXxBgsDFQUBSapfde/KEddyRphX57dv3tQCd3x29j3XQey
c+3itlbyM9aZ/FpOYuH2V64vi9khlk/20Ao3qVxbSEmZAjaRe5wKq2QrbXCpyJj6
m6gk613Uc1y4vdrxegY1S7o5edKxty1wVPbOiT8WnH34j9eMMNfbvJDNboFfMrU0
H3t8SyiJAtAgXrxzgxxksHZIIw45Bg1umnBHmE3LtbJ6G6MYKQ4pU10sSCIsObCg
PwFQiLwB/WGYS3dChe0G2DVEDjWk9ceWlIYokUfj4rGGBK4LGyulm6M1RWEAdvTq
YksDJWUd++uFQVd4l+whAoLIjvHEUvaevyqpuYYw2fGth48n1eIQEp8fB4yYBqGL
ILkWgEctvLaiO6007an+pSBp+lj2djO2n2QFuZvFA+IQXNfo6MM3r5n5Epnmn1+8
tigdmOKxGndSQthn2UBZ6v1Cvvr6NIAUI4GeV/VZw9kTuOTVGb+4a8qu0A+vqDL7
+mFQbuHt+55CVX7Sb4jobhwap0W/LD+RVI4mvIlZnT38BoHpRjQw1FpdixYgIByz
qVGcjokcrMSzf4v6UskK6cmhEQv8lQiIg9Iint4dVfP5LuCxgtBRn0o04JyHAOnc
/+jswXzgBmw8roQBg0XyHUlqux/xhrgfe1uVm83StjlCfqc+Lt1CigNR8Ra9Qxsc
HouXS2Tx1F35Qs+pwQATIHCBHMITH98hPvpUqU36Xo6koc6nsv1QmPtkOC/h8LXf
29TtMYia56MsedtljwuGhGhbYG2kHVJuDjER/f3PsED8jY41Jmd1vpzgMbcW18vC
w9uDGTTWTF8w4eUd7Wl9OY5L6Va1QD72eOaDQleDeFxjAvh7dDQrj5ALO2Y1YGAI
JgGb+yeeulo8dr/5Da0rZmsJH79JVRxZjZZ0ALBKCLcslYGtymnxubF4dE02Lw4V
QvYhHCfXPU7s2/Dc2e43Ri5eSW0uuJCPycTzzaIWvVPzqxQcAQvXQVePZ/P9uXgP
h/uzxiHmZUamnI2d3SLyOMlTie0mBbjkAcv6nCt7eEuHgdYzAZ/LJv5AV+CDOFV3
iNhl+zoICsRookonYfXTvltR4H8/DViWkBqMqVH+f1cIutP74BmYxBS6Yjy3TsYO
N7umivZKN+y2AVq39x88i3NuvoJWeh0hDdb+aejr3U9scHCogloXPjQNDQ5C+JjO
k9ckDQ1/0B4uH+f+Z4i2cKbZ6ViM4dVGd0nXXznQ+PaZ1VErL1V+yyzDvJ/PmR2/
U1v+mwTRM0u2/p+t0wquhgZlXXMV0PP83rLktdSwjRlFKAE1IvdIUcFwN0Aizp/h
bKXgPXfiPQ/4jRPXCGUJCGvpmNHA1hLGYyuyV9r4aGXmCQAq4eiiNyfC3o2Eujsa
V3gsAmtRwK3Ayxsa2+uBXcoYKklCzMCb/zHwYo5G9AbslE97uKM9xN75Q8JPaMAs
p1fGqZVfmgYfbDslsCEc6oaZWqZRIehy6/LgAHL8S1GbBjFctVSCIKjvDLVKNoIQ
aGHjP8oeFwbeD7OWsnKDJoN893EtDz6Fs/5dtd0ch6VbojfmupG+sW69M6q/rL5x
jyatYYn/p1o4V1G0KmqmB9/AA+fV8Y8idnBTqzV2FZsFaRNXEJVbptyZqz2tMF5B
Rfj14GdgddaAlQkLY1hZYBlZd+UzPHxkG+MJcAkdt6t8BssAcBQjV7TrElCOfV2j
TFC8ZSzlTKkJX+SRw+otk5jX7hUxjzDidhLM60esG4/G2YuuUiFyl55bV13/EU63
1bjP6xNQUcGC2gymYjkGN8r7wK7Cn+DAJ891ASW5EDLxWKxWtVjxp/lkFIJcp0BU
lJipdcyVgEmpSbziCXo0VOtST8zM9sC6HKi8jBNm2BZeOkZps/uXZagLCgucOioz
9zcsWD9E0cHsaIcSlD+u0tPTgX2xRQ8fW52hLSc9POdFLhnc69aa2WIYi03dcEA/
GQoI1hhqtxkbo+DbKnWN7izVsfN8R7CNQLEXfw6poCMR7XQ15nWyHDc7+th6Kjju
7n7zIb9L+ApR+r9+hP2zmeVb+Awr2nmHG/LnaJT5pMp/PlnpDR911rvxhagZvfXL
UeH3mR3YqMaQS6i72lvGRcsG5uLBEvT1wAzfvK/suxMBuf+ozd2X2AvR63gRzaeN
9kUL/dWOOiAzvndAQo1w49mZGc/gJBZihSEKhgOCu4K6g4gwaIJFrrgO4zqq73HJ
C9NaeQVE++03qZeBfwJEiQWffrFgqPxAFq18DD0xiytoLEv3WL938NSO1C/JmDLD
ZSKEzp8oA3H3WH6CqOs/VysAr2aNstXj1zhad+8gO7kZ4tc/YC/60xi8jKpcRkHb
+RGADgR9TC2WRacqKM5dlKwSm45lSR0KEdlzsm7YHykcZVkuyLTnbtPlg6ejsIWM
Hg8+MrPzNB3yS6lLakGwaZjfj8h+FKCduFaxG9BV8RfKp/KkRZhrH1ZyLxhCIhFf
x2QqhNFDYxhoV7yLE7hxp44nS2VBtRr5YCCMMbqtwl2XFaLPopjtZYWB2CvQGnJ+
ocbgzxCgXzP7TRaNA4Dz+avrJExkycp9yTeIFveEFALjrd2lmutbJMA2kT3nKjQU
Ed4v8OdfamD2bWtpU6b4wFIgIKpo0uOvc4NtF5SOFxfT7gZcH8is0/WThwEZkCcu
n6iXjIcIk2lNNGKM2nj6KNiqSp7uUbj+mrTKoaiHnp3Zq5ESZaDTyVwCDWDX8aHw
m6PAHKmwQaYkzK6qHVVG9wYnr23s2yYZI36atOBFpLhN2j/KsRh3qv+/QVorXLhg
gyxsAHTC+vGdngobi647dt0N0EbuYzhOJVIEjOPZ5Sp3N2z5G4gsn07A2pz2iTFI
u9FdnRIWKFPj7gmGqgEgz6JRMwFok8D5fJoM5vWxk/2w75K9OSGHN04/4rTJm+Il
PjDOTBmxTLpGQ+Ynozs5/+iwfeUMtzrRDOSXCnyjbm6+32SNgz8/ikaftItfJlPk
3UBA6Nin8c6ALtJy4WgpZXpTqvQiCnb9FsAKDuxg9hez6Rne29VX2JKHEirAU5XN
oRmTKpESR0sZ/3N4ZFITO9YZHMCeysENkf18acunInPY40e8LcByKvCkzCVGUiTB
MTbLfuT3we0L1SE67nEuQVeqQLBVK9SMXFdf8EXJPM9DHhNkwoeTmGjKykZ9qa98
YFtKlXfnyRMAvvdnhX1Kp+KXZFjPrXRQDMuSF092fQ0YQ+eGoUCG6Z8w32ZhGEqX
u+gYAtnEVrBj7kwO/hDM5pjSNzrqz0eYyNMTNMItcXoB3TNMKpHspfH2yrLB/fJm
YeZfnYAHmtP1h3IvWTHsNgcPidx6g10LnSFnboX1wlBAHg7hgfdCYfve7+BylBsI
IpiF2S9+S+AmwfXckUqFyj8EMv+ESi/4yJD70ZZzh6c3/iKnvGGQvHU3/zJEKPK6
OZbHIRgviE4LN4YxQblr9KtLwlhi2T3zaNnDBvctFGOPbNLTznVrmzMgnsRRIkug
xWa5Al4c5p8wFzRxKn2YiDTHOzzh1BsuFRAfJRgdMx0okm4NvUFG3qb+x6EqckDx
EfFmn2E/JWUvbWe9YgOP9lDSIidK52syDQX6NOEWRtMvkVBNwDPt2RSTxbukm/8i
CKB62+fxdcDwMWMzaAUlFXSUdZnysb17oNd4Y/koVU0bS2OsLxax5Qzc4cG1uiVx
L4WKb2PvPQsafm4WfvbqKQ8EamFvBXFfauZXhIH1DQ/DbpwkIdkWTRTrKz1yEZEe
QG1kBVYxNRuNLBCDARmzPGj573ojDuBxx1xOgws4JCRMq0pnPiReYY4RNfnOnnvO
loAajlErY70QZ+0obLTyENmX/8jhU0S+UFG3/8mSjlIY7Rc1hwZErWul2JkRuIFF
hU/w7tOgUR5Nl+8LaPVAJE50xVqLoc502fZZHFi4Klm/uVH2bR5IhOT4l82HBKjP
ltCzja+PgGw6CnbCYD/0HG8XGDf+vC3Z5gMbULOLyfCOrB3907N2DPKIz44ukF9m
Ujbf/prPU9j5asifxA31v0MNvNttN+LEmcTWkvE/e62HyQTXB8eeWBb+b5zyFkPU
B86LC4wSRfrGJ0XP0o3tn0bfe1JWZW0vMKrnsr596sib9fYpXKXu0UvVtxREvc0/
QHfqqCzxj3jYA33mQiu0f2RQt255dcyCjKLhoS06JDa+polAziR6WBJgTphr7uKd
EsMQp2WhSN/rQCES4GSU5AckLDe4XaJnKzIq5/DrtmV4kdekpC6C5+sNL/kiXRMq
jzsPAvICshfeL75LW796ZstsRGJa8oGdtu0jZQpBB0uJrhcOi/tO62A0mAZYZ5oG
ZlfJGr/+TOHr2ZuZKERakz/oX82iPwCZhS1isRYDhlMdNXCwEHTjXgaAcpmFxahV
KjTupMX0ON1guOBWtLQb0z7ikQ8gCKcLTCOwDVenDATUbRBqSLyRuLrGwxpfU06L
wl5W9ndsUYwxuXs+JMLS4mhohHlJU6bnwZeOrSENP6ukd8eKIIf9/Sv0Rwolfdnl
g3BKf1IED0IH2P2WffIKu2ZV2QMAeqwdUIINsfA7fg8SxkNid2u8oDo8dsFCczhD
w7sN3QRsbQ96X5rGkP94zIIjOOQnXjbMgRA43NC6ErymBbkMOx3BdCiFfyQ/Tse/
oKz3R1QGRZX50fYndw6lAguTbqogC7prGKf3PQ/mpuMGQRz0YNixQLHNguL0AmhA
5LwDxX/yqB4yRx/EWY9hubPdz05FEi31FdQR9LWua9Sjy2UWb3J87tn2vvxhgm8F
ucmLyUxKlZTmqVS5VDQP2Rknj5A9som8nRPtXXnsTPZLasnixJ3bcBLmAH+U6Muj
MHaB8GCEdPEJjX5oO9qyCRmoL3H+08q9PoLz4QYO9OgivDIDNyeN8kdgJwmQaJRP
eZ5UbXU3vqvWJWonOS8SLF4jJrCXzOc3FYo9uRuk1Ip7Y0IjEdjDIpU7qyfrjwt9
yNWVVYt/Z8WfCgSipOi4HnljC/M/RHh73/Kj/zWrMPYyRkHqWJ/PlJTkGWGl9ULq
pvmkmB7EkU1/CtIZ7xx480Cg4QhYawR9bUnExear3u4rHEHlwM2gyVHQCK/XsOmu
Nbp9pf/M34ZiB/OYuLvPf1ooQpwOd06tU+ipSY/l0nQusA9Iukspno6FFaIHOmrw
jLuLt1GYf7oLyIkAVtKDXXYhLLpenKuTMJv4qsAxYFJbSyw8zlKhV0rZFM95JY4F
yp4E8FZ8UI9hnLbSheFheSh1sN9fMERz1/ZKVd3JisRRIkIhcMphbSmM4WT1oYLS
IL7VuUNlFMM1AG/QM6iqZRMwvnAZ/JSbDxZBvlLDTPS1AwraS7a9UkKIn96YBgvM
i7rIb1gLWC7gwA7fbCzFuPc3GynYXVFqjsCycsrfvaL3pCqUwlPsFOigcurntV2+
zbhuvmoiwJs5phclSIIe+xl6P7Qlj3yhJjdkckgZF7+JsJHSc6SFo4kP25WeeLFB
n/55+MJ7dHlKQQT/sbiQSoKYXsRB6/6BFpDyqP8swnghNNmUwW/3mMdOAN8tavcX
WFWbLUpkigx6Pm0TmgDu2R67SO+p0ZAxROHvKqLNcEvozcZ1KyGHEkaDegQDbMPM
xFyiyhkTJqIMxh+AhaDVfPMvLARll6FonHz/3mtzpWz7Pe0eOTlGiEoL5ZSyTyNe
twltgEBAQwkNUXXrAEuSgZKg7uyb1wvsUrHOSzfhCvuz/1KRLK66kn3h3c0a9/S0
yZjJ6gb25dZzyPIgi/vGtoJG3u+DaPU+d9yBu2zalEr2gLF6aKpUuerlSXIWdHc4
x78j8yHJKnwDT4uEUetgFA==
`protect END_PROTECTED
