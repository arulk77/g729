`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
jTFYUNQAxofeeLqJtKeEJ/U5juaqdXvA/B1wIQ7DRwWFYBSTIJ/4eHZPSOf+8t5Z
60pXtHem7+aZDvnAetZrSPF3KX40gqIpmq/EJY42Q1c7rmDfTCjXtRonII5RNKcw
XKhKlaxOZF3K+sodopBvI36GHgjdND2L+Jl8rCd8Vb6ItvH2Zq7VofAfo15E1sD+
P/8W6UU/gXG3ofrHvp9pHb9EG9Gg4AqDGLjgF9nx9ipAmcroL6Y5fRbWTwJf0sru
Ep52nsHLeG0mte9tv5IKfFlUpg8TS5ADiJStJK3i7rETSHqpVsrKwZfeK2BB3Axj
voFl6ceJzjva0Avxxt+nEhRoYq8VuGJSNJzgREs7/Sg3t3V3r0uZ2IMIqqqwy4qL
PWTo9iCkL+aKUL+LFHKXW4jyBXXKylWSVEUZf7PQA2I=
`protect END_PROTECTED
