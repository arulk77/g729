`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44rXkfoJCqfCbkuFAd8vRBQ3NQi2HltmmLXSKw7bWuof
qJE4wG0nKZCLAx7o1mNP51RoyKICLRAKrQJuuQZdBqumbkS0zC6Wy//vLxvs6gBs
4ysfNlqgvBqzhldgECHNEnL2cA7/QlKjgjFRMRcpe/yGqr4q8O4WWh3aAylNu1HP
w2s/dCbaPDwo5H3aPbDCbWy3zrQQrg12bkEP83h24c7loAJcAzmklSysp3ZCodjI
IuY08we3s/KKEJHg6TXjUZlD+0PAZUlYp8c+F8FpAfTbDI0W4q4bkb0VBQbCD+7t
ZUxydABtZfuJjwVyokhxLzeSK47BFrFjRbSgDNp3JQQv0mdezpt1MB3lV54kYd8o
Q6B4wSMgH0qL2rPwXMv+Kg==
`protect END_PROTECTED
