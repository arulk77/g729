`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/k2AvPfi35SuxCF348AIGlOr919a0j1AnLkyqrhQ0Mo
0UCkvoJf05bJvcs4pU4SNd/LdxVDQGhUsEWRmhxyIPS75/XBp1J7qmlyEm0O3Bgq
HVFCFbU6eK+XtsBjfUAkfBsRdoHWZ81eOUyDisfsembznULWb+tDqhhyAYnq9p23
6Cx0fQbam9FEffNx86vOZh/IA93Ygmjpy9lq1G4ynUV7KPjzhS3kBsAMvFTy21EZ
/weMWZj9X8pO+A6Vp7eAUqI/aM1eTZiBefP3XKSCe+QYcFoe19bkNrrUFt4Q5z9r
4gLdMnGk1eDvdseYke74c1YPL9bOYtUKjeKIaG5PtPEcMNd6PhjAt0/eLewSt+6v
bIDoZq8mXbmWKtTFovZ4Ngc+Og5Tw7IM0PtXS4WEEWxecSFs04QtBbgn5IFJCoQ7
QxU+wtV1QT59kubQ6vaYw4QtgEetjnBCbGLRkCinQhcKW9w6kR5ea+KIWPyE7EO0
aeceV7W1urttEoGTfa8yAc009btHCqN+nzzkFRmZtcNZ/x5MpOSaD4Jqbqj/ES9R
wo205cW129g+a2evk54DEncf4k3+MhYPc5rkYunNG8IiJdz8Mf/W/bPYagpVCaYN
IIouavf26EcYtFwlxQO85SLetxshyQFHcFx3gDaHvGnfDDPxEJbz1uxI0TaVdHLf
80F+BRPweVR2aJyjQazzRwkmLGBrK82E28nGV8JGQUJBGPV8+jDwlGOu/tZsAFca
NT0tfPRLSrw2qml89hSXB8ZLib8c0lYHm7XqDghKAVxLRVcwl5MO9hajCupxdfXz
FUwIQA43qzN2/4fnwxjgK2kJZ6X/2rmjUX/Fiuw5KcvjWXH51mYxvgQSMIWtPi53
8NM5KDjieDCtQUvjAxAuWPqK5XZEQOgLad0hqb0oLgLnjgaVFpQjIyHOdYwOPH5l
xLgPK37Gs07WCNnQmkWs2hoGYvhDLqj5vlvgXY6bR2lT/bGS9OCNBEpT0rXpm8g5
ubIacSzoIXKtriQPTkJd2w==
`protect END_PROTECTED
