`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDARdGJOKnZZWZo53ME0LG03I4xHS++pIvP4Ocv+c2l2U7
siBuEYsYQR4Wf7Oa6uEZ4Y/5wdR2M6vOvtvktaf6522+ia5DPbDqOl04Hw/DXAKY
4PN1NkIjex1wvQL4fDvkcWWvTQ+ro8A4Q9+M1CSPAy2/8Ba1e6i9CyEGtwDCEklL
npIBjI6SnxsdmJKACIB5QsrOsPutRVx9fHIWO+RTWPnOx1DAjjWZ7Y9xFz4sw1jY
tvKi39VGn7AgT60cZABP/GYpJAJfxrohb/pIznj+tRKpGCNFQ5BT3+OwBXNP7TjL
CN/k/cmN/Cv9R4MJ786qAVHwZH5qUNRYaBrGNsIL6TOEkvCvVX0jXoh1aU6Cdgx3
2ES7BiD0vh9JT8YARGw9xXx9BpV3gjM/E78xLe0E1unGtK6STn6b2c91n4hlpGjp
XGqTvZ/5IjStFuPh4taSVKqn/jz05tlNGnzz+nJ/YUsG5rfdxRuAXfjAp+ezqmeC
aJGHKYWNbPj+Mcnl3ORDtJE7zlNFLJprVygU+geJYvs3qIwHIBVsf7Q0W3AYN+i+
e0+GM4AMsZ9cJyVvJ8tBZbCMcfwHp7xkkCCwEw/gJATZeOvt/9IopjkbYRLsNSM7
ryhrIkymgvfheZPp6SXtsoRLALTusbdhLWlp259eCeVh+04u9R7FsFQFjerU4hs7
Rvg1XXvemrNbj/OFMxFZRTt51xJ/RgKXtUhCwza9ibwcAwilTBLYro+HO7a6wqQD
Ikxzm8+F07Q366vou9DpSoGfwVs/WHMhu8JrTP28NDWdJtPYmgNJ++lg0As4H+IM
`protect END_PROTECTED
