`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xBbfU1psfzKlqbcIbQDvN91G9FIwdaOhrprHyjVtx/d
8qPSizhIqPsbqW6gZZ+jMfGiNn5pb9b0C41j3NpQxDqDLumvfDwnAySV+OGAEyra
CYFQaMGeYAcT+tFYeUnk48VXJna4wjUmxCCqv74WqC1G7zr/jAz38kzNLFWPIo0U
D/ErnqBWcDoAKAyuYR6ePw8R37LN5s2sfgDyB2z68EXVy5i+bITKFnWuvqbKs9Zu
byheSAtEgOg0O4rTj/QKLU63jqpOzSaAx9HGh+4xPLqcP8A/1tekQFXp0Tmukh4V
p2TRODj7qWypY2/CQztHLA==
`protect END_PROTECTED
