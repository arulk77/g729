`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
rPDUSYcLsRKcM2LZ4zppzEFRw36u+UwWPmDc6TPjnvwYV5Tl0P+bmYt3gluWrUCD
z4OcnQnqALB9di/gj66Y/vJGLt3jJI+AP0lD/+YUX+ISslO2kJUuPGdOlOjs9l6y
jJGbp0Xz+r5R4YMWJoK2SOKqTrhwjQwD4X24annJD6oAaSPl6GDe+eWaC8png6RC
TzI9kqKtcPok8LBBFST9BU5dGQ9yfTlnUFNjcGFzYOC0gmWAFCx/Q9EhUG91QJWu
jhfRk2S9FLtHdU0nBT04ZPxPJydoBWQaGCi8iQY5TJxGGH3osuB/e5QPDe+aE20Z
SZLI0AkbODtJJyWVHSjhn2iUgLH+203ct7dwp3Ak9Lo=
`protect END_PROTECTED
