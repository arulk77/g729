`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAR9KAalHJasoAwkVdKkHY5C/AGHkh6LNFOCmEqtroYO
Feg5nFCXWhPmDNwuZYllONO7yxY6kV5hqGph9gbOmQVCxCYsriL1F5hzOnH1/Xn+
c1aE5/BzgZC4R8rLX80MkU9YqeYoDkmTO+NKVHwT7aqt1JMgD8LdEIxWCcJeXw2b
8d5lK7SBe7C44yJmCgsVRg==
`protect END_PROTECTED
