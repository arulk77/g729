`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43v5mjpEbCV+KAMqKHBu4ACK81jc+SVdocvtDIwU2x9G
Lz+mrbKa8RipJaRIC3SXxatSUe16zWPUrQN6rMnYpOgvc6wAkaRETjk4FcmyyN2I
1SpmmN/FT5LjvpjOtu8tlO/8LmTNdBATzk0I5fp5TPmAqZ3lHMzVLSs7tq/iobzW
4C3BiCH3x9Ixvt0ya/zFr6bs8KPTyBBjFpxvj03FfhC7R56vxR768amsHSVW4YWM
0iJiercEA6wM5AB2nc0oDSdKCuknHqyS/dROhltgZh8v/kotoRDrraEIp3vKFIr/
YxCSiC1i6XsEPhqerkJtvA==
`protect END_PROTECTED
