`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
nyxv8b+fltrvVZJtnas+i7/3ZFIzmbfugbjm737atiFnIaxlbfx5nmxFiaq85qqm
+mjaK2Ci2iH3qDCTascfF+fUr93H7sHDPrff0ZaZd21XK9/xgF+wg3FzJwM5hxiB
jhO2lc2xwkmn0l5id5IFWSkJ2UyOuZ8SZoFjS8KziHsnurF+k9hwDPkmCnqHWAr7
v8PrF74XN1pPUifFvpvQdLJ+LPspJE7bXunEijWvUZuQma7T78EbpxXpctifUlJj
s6uIeXf/XXi8aTIgHrtFi0WKKc4HsihoRlzQePNhCq0AetYZ270wN8pGU5EcqRf0
7hycYSmbGow4BXScK9skt1clw0znDuJNf5dP8ip3S/4=
`protect END_PROTECTED
