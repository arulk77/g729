`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41lvD2VRLnhF8I7nn5/39B+6NRWnAN6hHVi2rYh7I4Xp
qQc1wzyv0Xo9Qr3U513zPcVxKaMNW3m83kfBg/2n5KXUfHHrHh7YEyre8B/OEnj8
YaZcuX60KcIdDTLyGMpaDdxx3CoTYqWLQUfJjMJ35ex9525p0aD0iQQjhJEJ+NR3
yXn1NeTTdz0nS4wN18RcdlbLZcui1NyiP5V9TGzc6OV5YarLdgPn1XvHvhzRjSyZ
KRpBwUwuKLcE3+LFlLNUGA==
`protect END_PROTECTED
