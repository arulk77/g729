`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
jm1bV7+s3SVsv5ZbLSw2usDziAgbFuJDBiikI/KTc4/wYMeN8xifp+AQX7VUtgeJ
GXS6fsgShF4W5cQ6Hu5uH2qGLg3lVdNGODjaepe3NfRQR6sGe/bXTcR7SijiPum8
QuuTIBEmue5t/iYxoQHZKOi7BjArioRvI4c4iarwcBFMv2w+z/INhE+OQgTCSn4C
NO5zwdcQH4xr3cyVPTDgvLwI6lRENAkoOFdZ2eL6RwTtgwXe8/Uvn5/i7CXa8mQi
ZcmgZuOw2ccEm0UiVL0cGDbn7QzFXC79OwoZjsRNW7gkGOFQYXKksDz3yrJ2lBgJ
84H8gunIxgf5KlZBYHUrcUTFq32y4/DbUAP6lCyNOEaKLhTwx0FGJNCTcPsertPd
trDB2dA8g6GKlBPxwPlAU7k62gbS4A3Zkni4AyFd4rwmpu+Sb0aPntGnWg8CbBTW
0Shxjr4m97epiOaCoRe3byo4ndbs2DF0NJqsDxOLMvT0Xj10Si4Y/hEXIHgPB49w
e5BbGmEGuiYvWMkiEmAaUzRD0kTSJCyWQqXxUTVmkxOxTU6mYN2pY4Qy6w2lwLFX
UqbKZY8i36HMyo75S+qh4Q==
`protect END_PROTECTED
