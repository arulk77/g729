`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
gXbLCjWpNqtBtbjs6YCZ+jnQlMcltQ+6S1nEti8q+D0jM/TLFL8xCAwncoHzRPKQ
xnRbnGTIpVL0pXJnpld5GyQRz4c8MTbeBBIJ/83k3MemfC40nXk3xgBArCYUl8cZ
I7e31sDOj9MwgdwzQncZiOoM7o86BNIqx1ncIy+uH0yU5dSQ8dMrYm2yKD9idXl0
`protect END_PROTECTED
