`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41Kzp33PolVOtvTqFc1ND+TD6Xb9efSUDTTVfbAYdIzT
ZOXTJo7t/kSYcvhNrLBOScUHdoKfKZe1J0g1W4aKY+z1h+QZCDPpgXz06zZw9emv
W5K/bZCqb5DHLZLoLbmmUC/uXj107Tm2gvPBdqh6UJ7tVVP2je5VeVk8xzW9ULOZ
e9kXAc3ZevJagRhk+DSSnVQJHvJQ+JTTTsHgtkEPW0jTxiqEjOorXc3F4aIKrLsi
yXpKzEV309akzdLyPQTVHYPUx+oWo2y9Zk/cFanhy9+GAW1XUrGX2SRJIbmKArnQ
vGlskWFtq1g37v/htAJYPgco9VSXFisGMLMcZkYAKafs0qok1/tC9iHITskG0AXr
UqOTnjmKjm5MZPKVAohdGw==
`protect END_PROTECTED
