`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
L74RQn/I/rqW7QuuI5+873Z0bbeXI85sGMES5r52DGMz34uUI2wv1TExxn4YjPxx
J3HyxwFgzPrMbNR9K1WKwQAWUXMIWp12KVv77GGgAw/Bas6SUsqshU45VTEY0oEM
f7fIrexXvzHFsQbxsm5yshQDHcIiiOBIeGPoYTa0WWJHga9RAXJStei+ITfrm5Wd
Xv2JYHAzdvSDWUDxEHKD9Ebqww9IXeuWPkXDFI03xz71Bwd+Sshm4+JqQyhu1y5X
8bunDejgECU7WSHmWCrbpvinU4giwcLlso/3pGuH45lyaPOEAOmfGp8pbuHobynF
lJSiE5ozSK52WBAvYTD35R3dOMIEnUpXwOmrz7UuI+4=
`protect END_PROTECTED
