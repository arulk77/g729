`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMIsnpuBBmRSWU6h1iB/BUz9smCkIab2KsHnxXH4F2/C
vlUpwmmSBQKh4vl0iL2lKwpsfbhwc/1tkdR9hv/5Aj8EXEKsHGO0sY2KR/HJaXLh
nWRtNNBYr6YLK9I7I7NPeQ/qyPDh6+i9HpRDRZI4Xh9MugnBIGo/Xb8JPFaya4hx
eG2K+dJDnJviuKJ90K2oBegKr4D1cOFT6lIky+HleLiM5xlYEimGTXNUyLsTy7DQ
mz1CrN2hI15HJ9LFuqKegBH4hQgGhL3o1wUArigRsL8EZUU/bSffC8Atvm+EluZO
AohrBHjj0ro9bNMnXHG0U73yb+11J5WepgT6S1AAU/Yn4r+pRBQCyytw98PXJFY1
PsKJOlE7dHKlGR+99/V6GfeUpLYBiDfy4Eu1QdZBkQyvEIET7BtPLS0wqz1OlYfm
t6k5q7srwLlLCgJAF8zxUOtsJPrMCackahb1/yYJ8e70ueK6yvT6JfdVNdzzCQul
BkPGZ3QbbieO75w5rXXaBvIHaKrcxfKis1Ujf4haP2atO3UlYUSjKk1W7PpN8K9i
N+B1ICGijSma5qAa5mrKEw==
`protect END_PROTECTED
