`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM7Y053y2L336ggONvRYBHVxGsiBzrPR6FXvAXNtbEEM
54WcThftUg9hXlwZ8EG02RfnyvnmJuEw0SG2gWHaih4IZqwDf2327soOP6ChbibO
S7r+x7JHAX7Dna2acWaLiCickeuYsbZTFVU/FwsTvliYhohNk46h4M/lIRcycMeg
hLhGObzFjSSh5TpNxtDj6u90MhIbTEfeP9hUk+d+q2QcDcAAzWd1J+H1XrAouzIn
`protect END_PROTECTED
