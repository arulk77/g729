`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN5sKuGErwqkWE509ZQ60hQ8tpNHHjfrWBVGITUu1MlDr
Ji/eagn8QNn31AdAjejc+Sq9Pn9WIOhaqpHp38ImIs7U5d8xUh52yB+shZiBAv1K
YnfZpaAoa8gBbwxD6lrP80eNg5PjUaSk3QKtKQSVf+88SiOIztKdYDOBpfjsWJaf
do3fj/SgVbA1wOfEMGbqSM/sQ8xftTM8jQKZHAIAqbFTtaqf9++LYiH2GHXnHPU9
uw8lgBzOxDw7lX+ujp3DcHK3SGTWTCM/8m+qMLeGrgQWY6HTDx+kzlLkJgSRRia3
PCUP2vfvivPimorND5oJCpkYuyGdk/7Dl7g1SQpIorzZXd8txW/VojZn/B7ItHv9
eMixmcNOwqVByG35fTW0NQYso/Nu9gyE0QAY+mbdtTYUiY+a9u+VQZrdxx2kRAWa
MrTcbNDQgqgaEL6WcTztIYmF+hgVVw548gydct3E8UDMGpNb1sbF+Nn0O+zxhexZ
1xGHfVhz8dqrXd3hFAFd96Ta9DKNytqLcRRS2rl537g5Ff3/ppazX1dkuQb8nBsZ
+zO9y6JFh5Z9auWPm9lRDQ6h9S/fUIAwupt2ocrWIb7v8lDzf+eqMaVVZ4vZv5/M
B5sCoKDQB64hsTiFiYiqPRZ72UuNqE/xgh8SfDyA0TA91popNRs42MJuYyefbuUw
3iPzim1iQ/caWbnqwkCrGAViI/ql/kEAA1OKd1eD07z3FqaRzAh3XzuiF+8yVmJk
74EvSjabnFafys73spNIPWu6NuAn58CS75u60zMhLw3vbGGAW4rx+SYuDDNgBFAr
1qtVwvbcmGkmUUKG2M18ltDLZTQq0W6ah8aecd3Q5E0nXZQmoCxMSlrutJsBGcQm
tTqJpX2peGiscHA97cpI7ax+9NjqiWEJ6KaTEwvCWIbqA9DbbZgqEwEGeXANquU6
riI5ukbo6/ulreffAghDtKMzKzJxKzZsQQ6lzY7xMuzwpAl4yX5K1l89k02NLL4P
rrA4rz8ZUw+QqIhb/uNNToCn9o3w3mg4vXuw+LHxKOX2XWnh5omNbzNFdKeOcVac
AlypBCiJi8RITsvrdUizBH5OIByMTS+S8j+WXB8KZFxKD6bFeG5FkEaNVVHRk9KO
rM9FR9vknN6UM/Dg7QRerYMcFI+psd9T//tUXUotkLyfSXPuE9Dx1QPQwSmCdOfe
F19ITl3dZDGZWwvnhFSpruF8oCZ6pdLVJ8oA6xdRhuPFnjh6atxTXDgbptBkqdX7
X/Kdhg/WaK3uZYAsMwTjz2kgj6chU1eYezXqY08z7zpewFqKhPeJcNLyVJF3qe/i
o6LDLhPCIEdZ/n6zlQIDbHSSD8Zu4GxbnwWfSYCaJv6BCB8r+62yd9TCnV+gps5D
rqNKV2hdEawdnb7WPJ3wfxwJU0CTFsFR0Eantw3v009hNdUdMnGxutb2yC94vc4O
I00s+0YjWBRyYgdbOn24RqSkWEBrgQkaPf8nnREMQn4MctIgu4zVC2M9JCqiaQeY
XTleEe6uHRrsRA24Qn6N7RBCaEQQAx8IDREAELlFPGFvfQn027HNOOHOvdY5an8M
aYSXQlxa35/Rr+0IPSDkgmjR/d9No2eeFZ5vY0t4qx5AdOKCTx7YnftNBRKeV3h0
csJHRyYqIeshI0o5z3KSw82J7rt9sA79zdWQh8JsxKxGzpQF9eenXvDoECx05rH/
PfVAWAWH2fNEChfJl6U8fikcY5WV5ARZytXPWKhVX9EISfEH5PYrxtviSCvzYo7y
Qs0D5RJxjPOSdMVXlOxJ++eymKEnbvmkvs8+wdzk89Gk0uXf6xZrCOU8I3boq61f
iCb46jMS8adNFl120IFGlkNPwfXaPe/guVBfpOnojx4kYZnCjwXZuEEUOuwR23SP
kElso82mNMnD151DTGTN8ZNuLLFzIRFpfxIRb3yrhnWoDKdCz26orNmdn0N0mSo9
pwVGSdqJsnOQ8HIeQ9AA0pL57YHLpTv0RdxzJ0eN1HfcJnMcLWT3MknpE280vXwU
r3Z9dFzSsIJ/+nXn8eA6+RyjnwYa5gwDkEjKNpUTJ5uivDwwuOKhxJquAUOsE7Ws
LzEvDZGDDFS41IwQE/GUTTnPiqx5daywFj8TZkSicoX757LUR1wqH4G4ZekHCUsl
2wztzqB1KSr94upTnNod3hoKzWaqBJdmpalcQIKDuewBZV3yRKvJ+wDAAj1bkn6z
eOqwpLGSlx/+EFOzkfmwYfDZQVTxVEoI9ttZ5ypFWZldHIzbhgKCKdJE/gjEMEG7
ihYESDyEvXyiBBRKQJvLlAo46vNklZbSswYPeS3qGtB26HMtQ5kXL2FPYk0fghh0
BZBx/cRAqaB3O1X1o2HJ+Z5lf2zRE2BiuphIgrQhtKqknyJu7347yh70a170+CMQ
CqTkrx2wWFPRAgg/kNSNpOrGFb8Ud/YsNWFnFvkNLXkB0h0PXpHY/cr+DJZN2JMD
hQbUASsbEKg1ZR50WNj2FSOTVQIMLWcb/tEkpWIFcwpMFRMIBMb8m6ii9KyyhOwD
kJH4UtDfesx9VkK+o27cQ1Z+vhQsatZ2aySj1jE/35/PKXR/Hk4V+zetL8G4juTK
ipbI7Yh8Aqv3EdzL+IP3MnZJXcqQ/XtVLf9/IgtXj5MMhseuBK9e7XIMwnGoHal/
nFyT6EvqcZN8ugrQDS5kujKaafBswUPQOVciJphpSVCNu6PrKj0P8J/0nTqB59+V
ZmB1C7o+JUNZ/NIaxX9cNdT5UE75yzbONAmLag8mcdB4mBDR9tVt10wjLxeAbtWH
tLPSt0S+moVPMKqON51dM/bCNgK6ZBXYf9+anikh190RXH1nqCzVadneyWMWEX8q
o/TJrIKQfM+vN8zrlVpAV+SToz8nkFroHpNKB8RZzuVQWFAyPHfZU+DRvd5BTfRT
xYLzuVCf/DqfhourGXUNSF/qyF/0HV2SUwEWqCtoUtrh8nCQ/QUUkpE95ZEbmm8N
pKuZuGbnjOyQRnjyz2VtWGsJr9gG/7ulX1pdSy/nKRVyA9octFmDEjbLk5tXlmIq
XLwOXZueXe7olYK4GJKjJT+cUZ6TQbz7F9kbjEcxkwSXlir+RIEkn+b0Bn280AFI
dTX8/d5ox2PG//zKEVB8/f44/MoApauLb3drbZjJjTtrs2R5MJ+KovtF+vmKZ3lD
lntc9MKe1k4SWC3bNuuNsUn5WvNJ3FD6UfmDqaoDFWZs2PCj7ztvGzxwxBBTewQS
gu9XrEyz0j+naQa1PMnhrclUAflKvLLtdBU5Fzpwevg1lFrFiZ+gTTlj1OvoWUc1
txNrd9K+dv9S/IwvjwxqwFd7PwEn398wu/nwwneJH+2nqlNpbF1uhuwBqVIm2YAi
tGFJtEVsRhNlqO4yJikPzacXoH5PAfVpm2QyqUaTyJc8xxCxoX4/6fFWNNtK/3BA
6pN65SWW7B1Ry4i1vW7cCa8QcWBaP7OeYDZUUdMxsMJ+umrSa+FDkALe+j3RHirP
k3KpWnyatlxMkNIeCBarLmeZBS+H736WrLh66XexV07WpEF3ybOr/fYPnIncV9x9
WmN4rhhNh5K7X1WQV9h5Py/7moag1uAiLUwgjEJ1/devBcXKc0rM/j7TOozzHA1k
jkZ77qVQiotBABU5PEdk+kzJe/lhDc8m1a7qnPQTKOy5wYyPz89TN/oZaN37fSN9
V76tc1aYj6cjswOgULHtwASAGDFgD2z3kTJvPx365fpNFbLMkhI9ScPZkTzepLSn
vM/NJiveElSRVDCTUE5qNxp/D89qYVkodlXutLLhrraPlWikpaS/kb/iVwHe5vj6
fncSXsN0JdzgLg4WTaAJ1XryvIWqvlkPMg1cTfT7ClwcMGoeDbZXUorCeCbfSjUs
4Q26id+Nh+CMEc6iqmdN/G2+Zth6w+lQUi5gvDp0FpMTwpXirlk+3eP4tq+qEcAp
InXGRKETYTzchH/AdVgGySusRyzaaa7isDfeDbYl9dx7/VAKxeUrtLaFwVNC/+uF
QXljDNdVtal3WIXzN4LNfM1XwbSykh20PAifhtzAQBeIuG9lsAZ9uNvLuGcvnYyu
/L6GerN5bRhelO6o5PCyshRvmOmlYu5KXg7Xmc+r9B9MCvCTLi1rfB81rYhZv0WX
iOp/KviEyrDVu43WemZGniW9+vwEHIPkNn2aENFsoTocY7qmUh15C8k5SvB5LCDy
m4G6w3Quj/g8IXWmOBEO+AurBmyFs+eDjA4p5PNunZdK/M7ci8CngFr0VW1j508t
Yw9JYKBFfHvT4yFUIOAhprwY12JEOtlrO/q1jAD8jSxJmdOFHBzojbG9562XulRR
Sm0zdgDez8PpS9imqdAK4PUIc4N3GXZVff1qf8hVugXoJAz8RNilcnEhraEGr8G0
OHDniKx8/DzGUG/9vjKvWx7z/TwnLehglj0aLlSHZjA46yCYCGYxxF18c74LSiwO
1pt/cBcdX1jt6sVFDVN3GCz7aOyHgDh48pGLq8BQI+sHZWZ+cHa6l7pBc3Frk1JV
3hcccUhAXiwkEieE7w1PV43Z2nbsHAK65riCgPzx7F27c1Db9/kjddIeLCTqiDKU
SSxqLIJ157gJQdwx9taQI0EqpWCyPkVn90CxMjqtHLruwFP10WIurMnGz5YI5gPR
tXQJsxi5KfPDofr2re/Tz9MvE29DnLheM9si9OFZOjQ7NJsvzcDrRgANMbdVWaBv
vk7DKga7jBbNI//Ny4NevfQP9QjR7+BgyDSUB8DpyQUbI8y6wA8Bks6PGEUF6RvY
plZhl+5cw/runBDDq5q5N9M/HirtXqmfmwl4+bp9bLv4k0b2xcG9YRDWddBwS6Cx
vf0m3f4qygQN8JKAMpKvuI3/BRPIZvGAN12ftdcDHRVZe+/iHTR1YK0d97Z81FnW
OYQNhamyuAeODtxXhZMggrG9PPGG2SpPxp7yvfbj+j2V8dXE5iwKowvnq2w+3UDO
x6qfBL6RKfTS3GRqaN1BBiQFV/j1Qurmb1PcNyfGq24P6pY1paNyiMW4iFwyLnlH
n9+Qb00AGA1R09u9o0fMzDo0Q30Pw4cJwhmlrYTwEbqtsf3WxRSRp5LJE6MwgcP3
zDqfzgFczXGsl8cyS8Wl0lSH30zLrWFqV8JVqRpCCmZ6DrdQ0rRbpw0ZoVjFUNCQ
cgFDpIiWC7TCleEb7bWlmJ8oNPY3eROazQ5RkvjHWIHN8rll/oNObwuX+qPlMXq8
26LkBQm2wRIxUIWUhXA8JX/KK4hMvuqlW2ILlNL6gAROjTG30FBed4xC++FrfqKb
4oL2e923OKwYhrMEpulTEF46tnUzTu/kODijhsVNR67iArYAL4NXfgxSYI1ZWELr
imjeCk7bzDMNzwdfP4ThUgqCNmcupZaqi3A4S/FFzuXwnqP2X9fwbn7bb7LwtqrM
hTkr7FD3sl59KYYPJOv92cF2VAGT3hBn2RkRl1w+VAH4Kn88X7H9p/MvtMNCdlsv
f0NXF8XTBqx5KPv/8j136RB+lPnwboBtK5YWoqalUDDWZAZfyoxUKFLAKbh5vbop
RWWf1AoipetIKHz3I/aSZCIUWewqQe9sT+pY2+xH4oAPwiojB6eSTXlQiUE1/Xxr
jX13I90WqUWEJ21pk0bhpRZX+K4y7VSmZUFYeyd/0LLcAukD9fru6k60raaL1ywr
zslP7czIfS30eLGGylbbTy6YuJYoIN1CKSFAl1F40EVJYa6pUySWKICIRORGR38O
XRge0f0oQeBWWzpGR2GyxSonrkvuyQRMnzq8gem+HuULfHrJ2YM5jXRlE0aG+S2R
8aqcV6HGivzAhTgdbDHS/K66hXPx1pBD7cQYa3Eo9CJd2j9TBbpqRsEXpD1uQQp1
OV5ZSp1sS2ATr8ObsJ+qFcKLYtDDg39xWSjTrQda5NTcBbtdumQXohgTJEbM+Pp/
Os0Ey+MPxrP5zpHKKX2xTy5MzKj6uk4aOmFgLQ0JxbQVKiXnA4BMa0qAQdczg4IR
xQ+y6wR0C5x7oFEfaa3GH+hoILpfrxojPXR8vWPvTnAc7EOuxeN+008Wrh+4q5Kk
GVKFrArUmbiZOtWh28y7nR19CRv27efFTfLCReZll3HiMOvVtf0ijpGhyyJsUxU2
eyCKnIioBCEm+GY8uICqdtMhXGIE12/J7jGtVDeo05Vquu8FJ7nLrEmRYuorw1p3
Z9z5UWzwHyHtzo6xi+MJI5YOU03Uk+gkP24S2NLN0IXPirNM6SDQWfuTn8uaUve0
MtkbyJH6goX1hJFLctRWug0ozNT/HeAlAIDrM4ayQveXx0QyG7YQnGtIPYd6FxlB
5dyV3KVd7JrXNzDnWO3Aa/36mWK8mKE/BHx+OhLbEjFsOmjBGlYlinzUdO5BloRb
pIf6bzHLZvYBl2CL52F2Gruk6yLrf3KE98ROIY/ou2cNeBmus/GKxsJ4dy2om7yh
meSdJbyPr+7WOm5Yl4kxvLr9+4riMXDVO53piFz7c5NfISCjXYMo1hpiMJd6Wndn
4b5VqYVhCCq12bC+Pc9GhemYswAF8Xh4N2GJY7R6GNgFzB26pmXzbsAmO3CJxhnD
G+2rs5cOxzn5rV7AZ+80ZDK9aqDxLEr/23crAbIPqDynyEWApsA8arXBRxnbjKzQ
ejT1Oo9+pvk3XJiQseOyUFfc5Qq5IBYTnSGs93zlYLOe+T2ALLXNeKhIppi4mHY4
0g97o5rPVvyqDI4+DzDLIvC2Q0Wtok8w+2l0/lVr4lMjQCfngQCtUH6FkzM781Uf
ZFqu8kI42n/Y9tKcebX0tao8vQmE0k6koHGzpWsexTUJaUv3+NqkiEDKiZ4T7ZwY
iCjXzUL+E5dufMlTqg+xnw==
`protect END_PROTECTED
