`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAXvhBZCxZEBBFhud2uQugBIYYzViWKUXynNW+OajtvbA
6rduIs9GvJGo/JgVIVDVQQr9bEXFhrUGWjYYpbSZah0FCdKuLBvni01wrj+0x6iQ
4qeibeWN+ts5phEcw9ZBgWt0rSlAhiiGl6IDlTopV6HN6MiMVkxzvrwLCuE9NIsL
uUd3ItpTutlLQ+WtCE93s+X8NFGo5dDg/pwT2w/gl3yGyrulLyHxuU/auyoq2UdL
jcqmdkQTAcrwYFoRtUkfL95fr/27v3XVkuH504n9a+NcmJl3ghfGec+xncCgi/yj
xWPe8WGHtc4DtqNz02kqzTyJu1w6FK8gIR+Lmjx1CxM/G742kT5rCk/cw8eVOCP8
dw3WchZOcDpmzf+TuntCwRxGFqr0tS6/q6IfyM9JMYAMaKyJhGyAOjrprdgox19I
oihZ03oFRNtgeCMjTbiXNM+QDMUQwvcVC4i2T7J09tNUMRyZ1nnqFb/j+x01z6jv
JYTyWV9W5XjqMLdZnLvEEZ4jzQblt1/i9+Wuj4Y8OonbNxUvxDG5OG00M6JL+hxo
EfXhV3crZXilHpcKthJwO7b9UBx0+9yK58X+YvIPgCJkAtST7XIXgIQLewEscisd
B7LB3tb+MVj1X56ACrXQe41o0HBtw8LmTtR5af2KH9cmi3TNu9HK2Mvkug4jO/S4
3sTsbbAmcXoOQj0gVRPKaHmDeg8wsMVV9X3CS1t8N3NB+rdzdnpLmJSRwccywILl
eLHpxju7Ht9Kj5ACDMZoxqB/7phzozLkICwHxukIr7Eis7M+QVYpXPxZ/ZoQCBHn
lQl4uOBqg+eNm65eJ0sVP2aOkufsi9CJqG4YxFyrsLqV/Tl8xLKTsaS9CfhliFoP
2M2gHUFGSGU+hVZBu3yaa2LHPAzOV63ZNxOCDaVHH12pNhHNAtT2kvk+DVakkvO6
r30i0wb+cuk3LnGgfLwe9rULZz875YxChfH0z9yvodifiZm8GwgKf59D9ZxtH2bZ
pd9ZjOn1BCbzKFaOQ4/xvLwscvUeX+iI+B3HSQyTbhhdH1WqXncleXay1+I6kVfw
WVUiOWieV7G5kyjmCju5p3SRb/PfclZy0BexJq2gsm776CD3mngKWyOHIK5X0WMF
H5s9ZSuaEk438bF6mdKpYVbdh6aQQxtjzvW/l8uADVH1tM7gtV2aBuleghuL8Jhy
QCVPR9xTWs2PO7QrFuXa0QnUrRhFkO3j5gayZi5lArkOph0S8Z8qU5AOzfgF7cqW
oSyZt+aHpQH42pBqXiM1Ee7NERCJoua+SD2LX+RRex+75wbtQj1Q36A8SJny4Bx4
nwb0iStWk9mvCkKzbIGrj8ti1B8JTfGbI38ClF9PZ97FKQBbxUyQWXRV6SR2Zdo4
QgpLmFFrG8KGbcidiruj8Q0K19ncFnM8HpySnSOlx184Ma8sE5micmjinOmg2cr+
lj8HVLEkrQB9m+m47BbqNlkT06h0d5We4cDzXuDGV3OrpgopiKohCJ3QUzRIKxyR
Ej0t1AfQVHjR99L52Za54wXtSQYwwlN88XrVXVibSr3duKyQk22XltA0x4BFftB0
EuvPTEVyft+Dxd66MSS+VRJhFiLliD4LWo69vkxtExV4d0JaBDmtHaLrbO9ZALsR
EWPbkNYuREuUJhwRwCKX2XNI+5KI14pT58tfn65fME4vTAzwqqYcxyXO52+IhvFo
C94pQgd/Vzj5/X4BvqOVxXYqpvOPSSZhkhy+IfskWtlXB8oE7aSNkW4WBoxNR0Lp
UvP/W6f/rOPGYSQ/3zTSQ2QoyVgfOh4NCsEXD4+jDP+DqhuobC9K/u1nEqWtEPmQ
D4xO0n6kS2lDG+G0uEDNdewoI+xaU9+VQDw2GM46fe0FcoVKKBt12UFyQLfkyP5C
FwUly77LvYYrstvGFowmcywSv9pUBVq/6Ppx6w4tg0oHucRLgdVvDf14Y6em+xK0
H/BwTOVb2ncCL0to+fIHLKTJsmOGl4R44drx7oRyBaMBV+PgFMD7BtHiJ1DpOGzZ
g1keJUMK0GDiFiPph7/70BymN12NLuLrWGhWKFBE34W+fuYLckmQpglUDFsUnS11
43eAoGRtgx7ywInd+3o2/NSqt4OFxtTd7oUbJ28tRJJNGBfpVVurGqoVZI5GQ866
s0c1AEQTkVpCHXIH5bItVh/R8wjY3SlAmGkEtFXzL0D1GsIdznGvfSz+x33q/Yqu
41IGxdbtlGjx7BxqNT/kU/9Plw1K3iVjJXUZqUrm/dV3gvcJJomfKRhEUk+ZhAks
LL/u6HRmwitI6ErkAecMlbjoUh7rd9sy3UqXr9MIsQ41+hZMQ3+54yLdByCXjM8X
w+myhbulcosjONiQ2xvyzP0Zfl6GzqOF7aVKMr9jY/od5w/eThDwNa0CgQ29YlBl
5d4Qj9dtYKIKOVv+ZI/6CrfNj1kEQcXRkLU+d0YrZraHuPH2LiK4/3ASLQHa98+r
gmDmrqkpntXGy4gjOmBAjDhzoMdrV3m5p3pcJ+hA7ALCUfUa3wzYDEVx8ztK7l7H
t2kZgMs4U82QQtWBMhSmqvtzWnMfP0rY56wIq427oVlMi65+v/UTgMi5zjlS/VRZ
ZbFTzo7q9+/b5bcHjNu4DHGZWSWq31E526bVoHbX21MKbF3uJh3C7i9nA1gfH0nv
jjiSXIe6M8D6vhliTUn9fvKNyW7kaStErvqWU7I1H5j6SRZt1Kb1xrgBM3yg+NGs
cC46ngjlOTDFmlsFmo2OUr76nb70pqZqxD6xFRnA5tkvU5eCCx9vajwDfSaALw9f
nQYIqwdunnH21H/ABvzttLmvBBqzA+ptAmN5FathwJz1AtVwYZ2EcNosq0mV1Ejf
vdgL8UFfyxCuBQy0heKTLzJE0n4ThpYHHmuRYNOCBZ/EpPlHp4SycrYCyVa7BYqt
iKr97hraIWugluYE6QaHD4KcDG/bm3gMlePCgeIUvHLcf0PRgC8Eakfs0NLD39IK
s/mlip61+DMyNyCarlVwviA/gFhzdTlE2rhB/5angHRpaT7O4MVPCqjImDoLT4HE
MPZdkw2+LjFATd5T7Fy9WaKzcNnF/pH3UgUBwHu9AMVQ28ekpGN9tON3ZJo22Vf3
RfLonQJGpolr8QFzoQdHspiG9imSY/5hBm/qLGugb8EPAM4oanhjJnXbnDNIpo0m
l2HN8z1a34T4abNaMtd1QeW9OX3cFrAYLnaRe3vRRaE4jMu05O9BM7tg6UxVxSfh
+W222QzofNMh1JzTdjl8fPLacVuDGB/d7qw0rijWO17ZRb0Xk4LkSZssdogf0z0N
m3ihziZq10T7Q1ph+0n8XKj2K75ezqJ43dnxXX0RZnPSDMA88nQ8UXKwt8jhQqzP
wSi1tHBPCNo3rf9LPeqPC+jpkT/+6UpYjT29LTGdxvKKf0+ApgJ7PePM2pWNSVk4
dfKGoMUPRs51QdZ+KZjEGcnKF2zeCYhUdt8oEpn68IN/3ol+/rWW/5EPf+sRuQUV
vo7wNBAnl/egP+83NE6TqRaXWZ2PN4DUNRGuUnFzS0x1QNmXOelWbMEOgLhwVyTJ
yoqdtb0uhCRpmpxF6pG26iAvNnZnAEwz1Nx5RN9JIyBazEkAAwl2QySmfcVqVsND
dlPWKGVncfcH4fy+VkFpiKMiW4qQONg6ptIaF0cHQba6BbzBmTllPeZsGzypsNo0
9s6KgETmzD9gsgvX8FTUqPpD+/0WwEY2vXMyEPNXIwlGPeEyKtK1p6MGxK+cG1C6
/z/ctff63L/HosyvfvDaTiP6IBr8S4lgZrZA3sA3EZD0abjxrF9j5EYu8Te+k6Cy
DJ/4hd4wnJzm3Sox0uVcuebApIMj4hvDe26cosnEQORuKRSRiE7c5V3IrQC4IwHL
ljdhdhcvxMl3fnR69+clreR9c+PROR20nkZZ4iLwfZiIM8UMQk/76IPUX765IDpd
fzettrH4f8pnX5+/SRW9bRLDxiPrVGBRf8D/SYqJI9HaDHDD1No02j/ksbM3zt7B
cuOt2/kuES80WoQ2AWgDsZzI2nHViosHKE5+AbRozMOYEx3ypDoAnJ0LJkOZba5z
eJLdI1v/7uN4c6COD00wYPMcJsF+ra4ePLEoyrzR8zmJUbf3ydDOvV/Mh6hWJY85
vNKshadgQBRP+fa8ETLaS+RQj3sIIUEXy9Xn+YDwGjj57Fc4uGiJqVb8qDYE1U6V
UkoD9Xy0HSFU0CJ0SJvpCFXxuf9CmKgREu7vtGW4f4iyaSA79fES/njrcjIQl20+
D03f1HAPBp4u4mc1T2Byd4HvQgIS6HUr06DExB0unlM89lnYZdzqCtdysQ5x/MXx
wrm+/tgkDoV/P6dlGl3tAFukANl13FAj1Xvht+thTK0CQ/6R4kFoX1kft5Veepba
3nM6ZqUOdEB8SrSQ+aFuxcmWjWvgotkoL/26JxTqtb3mn4qW59LT6UPYpj1Q/wIF
+bQ2loNhxtF82A9yTSSsiZ9xXwSF/SB8iOvd+sT2Fcm2EWh6Nm8aUrRzdzpLGAMl
Kv6lndu0M/OL22b1agF7MFX6fc5WmK8xiq//xnZ62JLxl1Ai2BgocSBtzXs10D7S
0ytzppId5dqdGcvZJbRgEhcdhgNESJIA8T8F+YmE7QDMNOtvkvLqGSUFy0OOUfZ5
fKFmBZLhBonrkHv1Ntqbzd42cfcN6Lf22o58fUCmtGZjH7wkC3mDeTrJhtZ5S8h7
fu8vr01I2QDp2I23oRWkvbXy9zqmGHrC0lnZAHxlz10c7R6KCPmZqbB2eyBpHGUf
m8MnZbbZf9Kwu48Id0xXn7PdAtcBu5Fj8u4kaiZHjdTGjrAqmw64+pOcr98E8SXP
TL7FvfeiKlkJ1HysGrYdLyJqFSQjSNZ9M3brWhhRSjtHUP5NjqFBv3IhSRAGl20I
f/UTsnpVtNo7IxDbvIee0TP4cYRPFtPP+027PQnQK/bw561ENtS61+UsO5mCl+SX
ytcnMK9ZcCVD91Am7r/8P4C2Oq+NWZpSUKZeeajcGtQqSuZPL+6zEivlVQzAKc38
/NJnbLesLnCTmhFjuicsuFnk5HkGoj1avw3PImP/eaBFD1f+oIvMWzr/y9hvAHBe
FKWkHvkhLhkv20caTdq/5VdLnjVPfkNAvj9sb38CDsdj5J/kF1qVsrDk7HystrgK
Aoj321VzyiimcGODs/NoXKaDGTGTmHkfqBPjhpyLCawjLPTBnrjCCO3QUmJ8znwt
iDJ7H3GNY7z2I/+lXVaP29fynvBPwSttFAYFMbND0Q7m5IuDZf8ew04eqSFkzUWN
22MhtXZJ0fia5B+wATLox7ptERlo8esDpo5wqIp3mCNrXUx8yj3h2YP1no5CJmeb
aToS5zJC34mKEyuuW2pbCNzAC/cghVidZL72vSJKGV47Zqco9rHX9E9yX1iJXqid
hjgCx25X2ccopZhJSulkS18wqP5sM+T27QxDZVWe8CKnxws2RBpr5t7YvR0YReyz
W73aensbzIRtv+vdo/pYn6flG5UhRCB1begIxV3wWiCYfNdU4dj14OrRtRNqSygY
2iZIeR9Ry2g3B38n8ZnxVgrqLXdva4Kxg9Ijp5wVl22yCdLJb1Q64+14V1Of46wk
6olEs7SyEJZmVm0DmXNdyzWEq4luyH94uMHOZxptB1/f4ZryEmM9Syzx/sPMc/B6
9quZea8GEEpUUqkYZ9iUzuh2wfXqBhyfMzi/cNmakC4zvFrR1ki02Y6Ka0pfUthO
THBj/z1GrK4Z68EEgHiYhrDQLVzlyvaJ0cVrBbWNa0ORrkUWZKh8h300ED0y1Cs+
hDZiN7Kasw34QtXsFc99/6PmokJJrAinlEfLhq41kdbLvtQscFYNTBBU+eampmUS
RnQxGTa2ZLtc9E1zRR40R7egEDH5GKLJCvPrQJLHqNI35+ygM1Wc9NoFGnPyoE96
RlGjTT995CgCFUIgTwlCL6QHZid8kInxlixbmclyC0Yum7cSU7i0cBqswKQEWMoB
+hUreLj7N/W9njG44nz0c8PLXSPXl6fd23UGWNhX2gAgGqHzDqKRUvhTDS7+QAGW
4WVbqTDEuYfNZE3VYwOGagJV2jq4l0AM4YX7f2UlnSj/IoC2NfJylslkGG14zPjq
AbCBgI7zs7XOIbj1f9z+1OtGE8+WU4EXcf9BD81WoTJVgRAO1eeqbBrlu8Qjag0z
TT6sfozBevx4KH56zz6UNaEQEsV6zgx1PQMuBH00cQKthgVBEtxryam9dX7B2c3S
iZ84WTjMOdlI2NQeEBcuI2AiriGbQoS3fhpDS2AgiBc75XBtSHdCtlMqvcPB3lsS
0NngxMVK9XJSP7+RaU2uIUuPQLfDF8kV2CwubwElrU4TEq1bzuFvm82YpyjLuRh8
Z8dG7R02vo5cVzvjPgAKN0ka9tn3NoD5cKD5APip2vcEMKSfXJdJv7aF0J/O3PdY
xITYITv4efllXsSZnJFdLrTcKnlH9zAPf4wcpr3XQtz+4kQqZnV3yuNrocq4RKp1
CU7KUEeM58/nZGf32TQE5Ke7iQBoC47KZzcMkLWtDk6YB7qOHynZ2qn2HVA/XAV7
0nRAKAZZWQ6RySbA6kX7NCnXlfADzbkziOGxi/+QFZleyg0Q9HKCt6hBuyLwtuW0
t5Xi61GIm6F6WrTTOYJqH7yy6gA0R3+n2bgND364E2J6FC2WEHjnJnfz8d8k7+Bx
/ThZ6TJUEy9d/7kfPxO7WLPJU3nhH83fEi32uA4GFVImwYuK4OV/8PxWcqCPOFrt
ZccYJQqyAA6LynzvLc+fWMBrbBeBi00Ez4ED8C2hz/TnmFPYYQyDfHwWgHr5PKXn
IXYSqk22SfCk2UTjWUGhXOf3gpRVeWW+nggxwBREwH5dXSMnN8jmAVnqzg4zUkEu
A46XNosN2TInroi+q6F+n0DLrU7WNcrqyW3wfl7XIWNLRNSLmWmqvUX7F/b2F1Js
d/rv8yDX0YpZFeuqrzaUJgj1ICpXxAWh7jElwGM9TideedX/fi3iUWJOOEj65krZ
2k22jj7fG694IL92G5DIYkUZziuaWGaz2hcPPT1DgEmUMi6TUG9UbU6OPaJJ+qbN
ldzrYtGEeVeatigw2yprvsJuGXIJCfK5FxE6seCkm0r7LVuO382Dc5UsfzHQxZJC
vjvAZGC1bC8nCPTvE+uB69ZdWcEpK40SLWBBldFcRpqz5RE4WMhfz9LOiWIVOgES
gZ36Q63l9mop42iTKptsFQglVSjLDkiSwkgyUW7/4x79VhZPBPTR6oQNEJNDv07f
tJAtPdlKhEU6Qlqt2yKKonkSc4vYRx33kEPO1eLjCiwUOq7vCYIQg6TPG/4ALcrG
r8dsJs3uf3gPD4fS4s/5ZgUUROU+2PdONMG7LdSBzm5QITvhSIQwfFATiGCOugPU
nb0MwWqHuIaWYougOqwrpJz5BPLRwus7yFG5xsT/6hm/0j6MHN8Pu0wb52LC+fnU
t/eU/vQ6J9sI96bPNAYGm3ZhtA/HgTFV9eVSpkvrH+BYnwS4SMsKj+3dAtaXTrMl
/dVljlifN+DHqAmdOXUpofw0sr/eZdEv1gRiQgOytelcrJMjkgp47xQXE8jLoAXV
pQ7vVAZxIAchOqoc67KMJSBHZ5D0K1gFEIXZ2dujUN/AIccGhEW9qRa8ErfSXH3n
ABgHKm3VHYM5zpFgAOYz7o0kX1fNIIAHsSAoyqRY/JFjW36jsovSNBec6Q79E/dy
RXM/Dsff+As2jhSgnAFWzXuemjWHsFeka5qCf8R4EEuPctrPavh7199yeqmLk8WS
TLGXseRqYEEke4FS+8tZq5zZC7oix0FlWYmWUK7Zt8QkP9qTIIpp1HkGcNwqMqIN
En62TAVKb6FBYeOHjh410Pdx8LWQNV4bOXA9fHUcE7WORmkb9Dh+B3nq+bFGikYW
9NhaHb+iTpN7Airp8sUQc6pLV3NFsSxBv8+G68Te6tSEVLPAGP6blFpJ5ndnjZsP
PLfoC69lGQ7EAzZe4zKRSIg9TL4xLTHoTAHosOcvbBbSWTYDdW0XAjTEs4VNIthh
N3wSpu16B2ZbUTYcAotevEtvWkUmck66FkS8CuHhISLmF6wBO3HPkvKnfIpNtGHv
Y9K56SH/W9BG2FeSKs9TVeFkJYQTqMuGzHtDJjCf0KZrfovf7b3nspauAvL2ctj3
PL0KunBK23dXbci2BsA86zPiZzAdc0MYr0woUvqCd69xzInSBPoKABy/53xpg5fF
OP6aP+htwF/eTnRybKNBo+1GHk4tVeWv9DPye0bCwUvpZBRIIbRgpf8QIKnG59qy
c/ULqfiYv5oWgv1YwusOTV10src81VEcddxBxlgDDbCwgqqRcH6Wz3L9jEy6LyXb
Cnzn2gK+rFyZYXXe439Lj4C7cPLD9V8ZHdM/+645GCbjGiwb2fY8LoFfZwKcjiGb
d0+e9Kz/V1dddcu+jABEKbQuuHodpj0fAZM3oQmHq3YRX8nky8EO7oLyYoai4efQ
R4/VON8bdzckPwi/ZHhTaYMDEixyfulD6TV3+CkBzJL5Q3So5SZniGoCqyRtl7UF
7Ouf5lLpXqU24JhoWnu9NbTaa+3t54AHPK89NBCvJAlihbqA05KRUYVvLvkudWUd
yjPuQbNdNCfY9UomK3FumEntvqLUFLRvIfTkCyYoOiChU1++4Cx6N/FXxKyx3lJz
ArjKN0U56D1uVCei8fubjRcWxTzbz0rOIqUFQEagDb8oMDzaORW02C14WfLjDK1d
rpSawaZdJVFmkCFqzmQrnKYy9xJvY3jtTEZydFe+sO/sDcVl84Gz2X4pt0v/47l2
4bCV6fUUnq+lIYduZufUrfgAxBpp+fi10D/UDTOj48GUttBYVQykAJDEP3pngO7I
DcYiV5/BNJj1/kcsgsJb/G2Q4tud97u5+5qfWc3A7YVX2oslSAgiYlkTfoxJu4Jt
jq6JzdUsuU3TmIdQlJU1vNCfS5PxDDIRLfHLI0MFRcm4U9dWXKMCtvHnpYXEMMNN
mbg/tbsXcyLfoMrdD//9qoc/MWwyWWpf1ekxNzHOeEKAS12k3V6xmbWDhs+GS+3L
X1r14uGWf+LFEeh33NocwIIImQaEG64/RJfFPxSKCu438u3vlwlnZKmMUZ3YL+86
JQkqFW3SD6HVuKapBPgWKTlPHNlvhcUYeuQMozcwD396DzL4g711naWVF8aKRqFI
vbMSpDAf46FR0AoE3+5YpqHtW+C4dGt7XFLuDOJffr6o9KC5ydAf7Im1LCc3Cive
mFVJyCL2W1GEZVwtONgIPsd1Bhkl5d/dYrSyKAYjihbu/egcGg5XJcWp5sfhqgoc
E1nMeJA1niOAhuoZDeBr3v2KKv0CL5kguWB+0QFPqvUFbXs4szShINvIweBmxn+5
9grCldgUVCHX/CEDPLJnPD87fuQXC6INQ5uSK6YgGSgm5M3Hdmq6BwDi4w7LkkRx
+Wpgmgp4uCQo2JUjKqhoBikUJPXafzTheS1os17KGSODAfiYZoQMlGNY1ABjplW5
qSWw3NFsQAJmYzp5WabtnYWYF8ZLpgKGud2GX+6cH3QJCGF41EmptX1eLzNj6Vsq
4PLkABFOmullTZscIZQ94h/Ly2r8F03/HKVuaA4mPdIHjBZZvWx133tZn1UYgfNB
XEvEaTxOzt6MZiFw4Y3JvooW8BoNqYwXr/7W8mMkbuqAY8z859c4RBbFp6Pig8ZT
PhlJf4Mf0qhkjhVojf2RojFI4bC+vdoqmVoT5/mJWU1Ud1idT0PncMl45J/CE8rW
KOs7SdmBIy98MMiRQvDDTdfPRp+7v08RvzOQppWBIIfpxHTcGBq+tmrQeb1Cax2R
eONH0gTWqctBZcGYRjZVJJ042SNEfKvnlgBcralR9H/AkmA6k15FPlhpbaU2hx3u
Gv+/YHGSw20iIsiTKkURhI3P1K8hQb7ysa0PvqZgSiiXvrcRF4/81tPVf1/NX56d
cLdDEGzbwhZLDQSNDFRGzQNtBaw1lX7Izr2ZBfmjN38zjfwLQSnTJQHRGYqxwYnf
p9aFdPmEv7qs/uJRVcuEwMfh95KaxAvhxxYbIafI7G4gb2kR9svPHF3yXEWljiwj
LGDKPy5VBkPZnYoF66xuVaia6dUoF/h0TxlAz76PvQhQLi1GG+fzeU5YeecPPpzl
xBgN7OmAsXbVFLhylRhJPXML3oreMTOBF1a0ebapA1/tcwdI23mOwlZfLlwFcJKW
jU8adcUyOdlW834YX3UHJuBiE8AvKutNoo8RmuIdW6hpeDFZYobpL5Twza8UVqEc
C3QSf/0mzJcItx5RHsJfZAIwLRmfYdOsQ59KHnNPq34yszKnNZXu5yTs+4h0xgaD
UZB1cenxhnPyWs0+dZQdFszWlTl6SFiMUBWu0Au7PrSBAjrFn+5OPt8jpr8GLo3d
TF4CA3g3rKe9WbOpVzZcjVVFr4XlV2gCgQG6HdRkUFY0QQIhMPA4j/1ZLce6sQ4y
I0WWkrJZY9aoMKnGIw3z+7mBoeHwcO1aTLuAti2nE5V2Begl0GZFVct/bLk6O7Ao
zhp68+OqQByv5WXLy3IhwT7lZ9S8Quf2KLz7vaQmCcRgmlZbOGWG9ItXhDe1ucBC
S9u8Sdmj0amof8jcSyw8kwujQ+gqAlZu80Z3iVSR5YBasZvZ1rjs0nml5/oKtLMP
4vypYnqlO5fEBcoEWPw467slnKCs6s9uIr6paWn8jtPSlRKjKVK/3UK6SJpyapat
A4DH0AqYf17nylwFQNdqNX2S+D8dtuzNUk7onfADLIUlbph4DO6Bg4/yf/wJjoDM
EEZ3QvqxB0/hGHMh9MsQQyn+700akl9XRL1X14bTZOXxmFJOI/yQp621Q/b90nL0
Bplne2KoUtPOGAnGgdYF4eumHojYkn6jdNQBPHKDViH7Szh9+AHE+3TsVYCS838A
5pEZ7cfqurb0cw+HYb1uYzcgvBloE1CUIITXB725W9fUORFxefAW8GJI9fgrt4WW
Vuh70wHfw99rq+pb//Ex8ESmdPIGenpbn84zB6Z8SOTyAbdcDM/ExCis6hcWN52N
U2Op3BgrAgxgYHOCgmiitcRxRfWNyONM6ET7OriXqaOgLqhCptntwlaS47wCjLcz
0bvv+VqI9YcUBiGOxXEDZmxVE2B6WWgLNU5mu5Or67R2/JQ90RGWgPAo5+seJtDz
iqtw3zhmpwDGJQIkiG0DEtvbd23H4nzpnE2ytFQJXQF0ZOT4rcb5N9jYN+tH9rB1
6dC05yUghLVlnNcAJmmRL5NJrZ2dmG6fentue87UjwqlU+AwNmNdO3WOFoPxQNU2
WGpH5Af1JDjGqki36hrWTygZvcbnRgcEKhD4DFKwaE9HbkVGyqVDFrjrEaAXLiaQ
L+VaCumRCjrt8HHgw3hrPHuy2pce5htsmvHKlQtxs/cNiogAwFLj10uTDtYllY3D
4Jnjf0uHHK7Jm0k8dpRIDKbxQF9xctGA82KDrJxnwUoVmKZV2jP323hPYlTNrJsx
kOrF/PAdPtTBtKwCqVUM3aor2U8gYOVGYHmmlmi/UW2vaM13J5ZH7oqIkcEadqlc
A6wqtWpoARGiY3atS9PKOSPw24rUx1IJ+ktJugbSxjrY2rnNbry4e1TLQMnpUd9A
u/TE866d6M01oUC+QvXdxQ5ItHTYs46apUOZ+UwS5/XNy76YNZNo9WQiaUHLXYvJ
PL7ybRT8dJASDGhd2eTcucAhVdul7I38OdW5CengtUOcokzWqO7MAPXRwoZEsEmB
a0ZPHudKRE2mnRgKrBdrlA3II5c/Qlu4aEgNHmouX4IcQY96+FE/0SSLACgWgRt2
z72jxf2Lz9DxOvqRw93xUJN6lVVGJ8tUmPlfFcsJEd6uq5jOg6d4qe/lOhC2M3XE
7DWImoSOhoxpzDw2bFhsgGxzfMz4iG7sXMfZyiVKPYGfGs2n5e8DWo5enbLtT2CU
mn48D56fCy5+mzr8jey1bMOvO5YcmxiWcXPZUT9Z7QPcFRY6Unf1LhSM6/GEOCOX
FxhXRKGpXXBviEwHy3WfIR/E0bPdU1SOyIwHq2P7edQfLqOteqGQcEk5RfhO4XTh
smlYZ0zZg04oYcQNfXeeO7s4m7Mt1FTw4CNqwdtMeyfTajdZ0kPQcQkyDoKza9/G
jEobDE0VK0V3rnU92/Gg09BYib3hL79RsjiCU/SRgPKOtDm7eGMjOkc3LMEb6MqH
G/kHyesv+ZAAdnO4UeXewSE1UuRdfk8n5byHAp4UqsyIU61B+JQ+a68bYuONguD3
m+ZBZcloRRyUa+DwSWDeMeOsYSv0KwQV5y5snc1f+McZLQ4MVds0xlEPZqHghAy4
CcNiHoxKwv35Tm2U5bzaQx3Nq43KqOGf5lblSTMjWaQPyowPTejrcX58cJ8RNA52
xOPWcIdUcqhdkClEPit6oYM+iMgXiPmYApJhTby1aCHheP8k5W0fMbLgbzLYZM9A
GeJoh5YWgkn22esRzQ8WaJ2zcqD04FEtTbXTV24XmacO6veuNyFesz8SLgpEAui3
m3vuXwzDEPXRd7c2KDW7Am7r5NmRA0+Fch1maUzONVNaa70Oc42DUqLslBQWGH+v
2TraOdgPDS95dR7DFgJe27wB3Ak9fmXcXU8z3TTVnLXQqsnJA3sUHNvtgQcf+B5N
0ciuxbsDvcJQXO7IaSyNielEDUa3iavdxW0dxUz98eaTrP6GGwthT/dQj5Jy3+ED
Gl8XCwOKk0L86zjMmuiTRfj/ScFXcPWHvrFkrEEYG4YIVtF/nB1tFtLL5/sA3fLp
l/bgbw70BrmgdLrHvfy0utXvXy6a+uRamW1mEzEh1103hhx+Zb1U5p8zGdMQlW34
rrpqEaYji8HpKd2ywpaAa7GMqRnS5l2Eyj8L2L/RBbiiD5wlQO/wp9cgtevFjuVq
6FrdKPq3L8yO/PXGjdtipkDgaGDw5OqyL3g+h3uv8TVMCJ222VOqf3BvcuEK68Zv
+P3+0AIJ414p00yEt2kIqxJHyGr/Nf/O47lfPFm+FIJxM80buG0zfQotbLKtl3GV
VR3yMEabLVBxbxcRHVBmuJi56HZBiIn3y9eMY82v9sNA+nR76rF+b8ke/LTqxabu
1XP2fiXOPaI/31Xd5XDvWDqKwG+rHiVoeX53FQMNGY3ll0mpajA/SQK+1g6JZe8V
ckGaa53kAjiAnfLvSV/gBJjBJNWZ1mX1oN4X0OGG0Qw40lEAj76Dv8jAK6nFxftI
EDWDIGh3xYyd6AzV2FK7zEMgqJiUjw4zVtlouVpKVK9ybi9RIMEtKQ7R5nI2cXb7
ddFjKYXk9yFbm/qLgqkM2veb0XxtSwUxd/EcNv+LWD/JfogY9N0BYCMqJLCWyxrj
FMFqbVPo1NdkgnvXVmk3eECe6LOmJmyKn8eHAUD5CQPLsm5AcCSZMYGdJatNsRfo
OcSJ6OMth39yIrtHphfutOP2ypSp6K8MStcyNR+Pjd6zJBV9YaE6HzOrp2jfL90W
bIUIDUDkcPK70r+DPcalqXgLiOexSRdBtT+DvSiJ25LUcyAkaX3w868afkmiWJ09
7vgTLXPNPBM0/WQJG9caSrl6zV/t/fWxuc+27+dzKih7KynSjEP6dpDYUT29ZxKu
WpQb3ZAJeSw1I0TozzWeCC3Jqa4k7H6ax0z9lL5N0OhWcaZrkFHqT+kve/01eKAi
yF8ka/ZcWkpHXQoMp4pANuftCWaNZAjd0iZ1LgVG1hIwnqPmt4WfiXWqdJ87uI6L
0ZCGJccMvEUuzUV4nS+lO98cvzpLIOTZjsOZU2GZOjP2MjYYTBEiYjy4pFKflSAa
6S7t52Hpc8684ozme7S58tIRf2MMPWvRZpr3+GuMvpGPwboF4afQVIHcMTlR7ocf
ZnkndS1iAiOLdAvdblF7r9nOeGrQe8Atd+I4O65+pW0HaAzw8MfL1vh1oBjKZl7a
zvyJrYwowWl5Jf5FH6K5RpoCVf+/mE7qjwChk2xr6g4LBHSe96jz9hb6icOMfUaf
G4vJzjCi8q7qqjOSASyz8ODbnI7MEFoyxspXHLtZuUGocmHXzKtWMvNIKvDcg4zS
cntZZToFsEb23pgbNl1yMqyQO1IFDSkbJIk4ZcqUY6ZHKbFocTBcwWR8yiwg5+cO
lRGsRy89+LvgM+WluAoCvkm0TulQxEeUgrXAX0sAgkUxjoEWU5cQ8jCgX/PKw+/7
R7haOc/Ig0nQgTRfAYzxewgofz3S0TXAI4SzoEAvK3PQX1V4Mn44ekvxdUid15/D
4SIbKWW5evEX1tMdS8XS5vsHw1vieH+oaXpVJpciN6KY76D59e21Me3qNl32QG4W
BLlZeloFaxQ5iFnaifUy4U6V8Ho86n4vA7e8bAiskwg4DuUKucg3AzPDLpFRLsDy
8s0qnck7ByMhwvknljxEDN6IIJgdUlUe9tKX3CmCeMHhznUoqC0tDUxKVzyue3Ib
ZH7K8mOPrR3D6MSNtvLBdAszX2/niVIOZHtIP31sCIP33tFa5oOUU6iK3IEfcMuf
sOb3TEAFR1PogTLeSaPyBQP8n0W+4fF+kVKI7SIFjBUlqiEiaP6J1udS7E8IRU1d
MXB6DVmizEWivkptpG+MVu2lk4oIZf30mLMW0vqsWS+TWG6FRGX2VWJglSPYtYdR
5OdVTDe1IVPfnMZhVk31yYfilMonWQljR1QOkJu3ujNpUHyitb367RT/HpmLKJva
57x/NR/Lg5tBY+qtbMyQT2Eem7b5On2YqEH9oLuLHH/3kPJMkqyrEkZK2hvowH9n
n2He4FeZmdyn2HDU/18LKD8RJ7r81Q7SE2a9tOpL25K6QsWx7qfEfsdb9Io2JZwf
qYvdqgHdsvba53BFgIS9bdzxf4vipVaQgRS4TcLa2uTdNykUkE8zUrYmvXWH4Pum
MThHV/ldvelCZ2Hppp72psld82N8piMoMzcvZGG1Fz8F9OSRb/isgHV/uzIWcG3d
fHvTIoWoOpyVtGYwVKRn7WPV2hxccjNnFZ0RgAi/I0ZMC9Wgco578rMkU7FOVrBg
U5qZdtsZkD8/8MPix3LENeDCRJQHLSkVTO0dheYjGcnZRXXL4k/F6tyzC6nvkYAb
deR0khmGfqm28Fs0RraCu2A49Omy9aM2cSfKICqrGzu8NqMLxC09G2sx7k0zE2aO
bMXSSbIb7W5wnXiKZmzTElGCC9V9d9ashvhPtVwkQXZfIL17to9S4uhAkBDNrYok
pA03X/DSu3rYlwybmsdtNgx24G+EFC3JCpQky9NudubhCK/PjxiD0lA6lxxyYqaz
CnA+/0nu6oiO7CtlDqfxF7x9zQjX2ZWvh8OyLvSdDCGgbmpNPhhiEdCXG1A8DMdx
dy3huEj9JKxf/AWOc2w055mTXhhVDHgq6Cwhrgx9xKRh8UTmkqJuvCuxgiEnqaKU
lmhNd4Jq2riQceJezeb+nSP2rojC4JJ91uUWPsEnas18bF4OttXSiBcmTkAO608y
phOuTbMdLCXd7UPPdjRm/MsWghsm/b5NYjOxyibc2OxUktslqVouUMz0pUzBOU4n
/MMtPxh5b9xC0lWNO4ZikZ6Bki+OKiIAyl5suMEHA/ZHYFNnuwjEOvJkFkobP4eT
20fn7N+tzH6z5sqFTf/8hBsdXMk7RHqELfYuV4iv4maGMf1mp6iwnjzPIABzQnHB
4UmKze3O1T7yjiDG7Eh+Q6SQLJZbnuF7CL+n7yPZjMBA4Pgis2NdylWiIPdmtiHq
OXH2uV5py84uYnT3dNjEDKjEfjo4xQlHRbxUI9YyvMDe9AT0C5TPrdNXW+CatAe3
fq47v2hp/Dy4QlKTTfWZkZjcPfqcMtzMKOOWMUieJl1hfLH+ZYntrOYqnf/hq28A
15nn53wT86kT+qj1jJkQcZceyFsuL5mx7QnuXPrmBLIOy98vxT4aGeMwAKBGgDdT
GBVqTjjy4pBKj94SOw889pSAovbEgslsHmIWuUBUcTt0eUDL9pgxCiVXiEzxNmH+
oPvCfwknFbddfCknzFcLunwZN10+k32adXwUa5VtmgMb+Vjv1V88/P16HG2Tm8Md
8oNDR9Pll6mKlAAzKonbu8YeEQ+2Z/533YA11KOvnQDU7alx1g1JjqmTZaOyk8aB
OHF9taGj5wSBsoYw5PA67fLLFrgz4/CVwbMlpeQzmEuPgpFDHrsVd3ct2+tlyqjF
P1AEzTgfBUoY2+D3iUpoPdQJtJ7wSHy+MGbpBvvWcWezk3te50nsRKfA6xf0XtiK
JHCV7+KXzlGN8W5DoynVs+5RHU5qrixZlIkDKNpPn4idqSLsAOXJ8FT8L7KI96Rc
XLvHeyER+6tb1fJLG2ARUEk3oJcD0L1tbfgM+K+l0L5WFCcUtyWuBKQ6OCmYTr7j
LNxaueoZ+sAj0YOFv3jkQjiqYqfTMgHVFuMeTZjwxXTXrXerIsNavCuPxlLAeCxk
Egm5ULaJ52ArOMkh550q3Q7o2EXh0EYaIEA6W2Y73a3D/BDMwJbM5f6eSEwiHPhR
DgRI0DcvM8IW7Gd97cCbkQcmJBolepzraS78W1hxKqyfeDrWK9hUg2b55vYdDXwb
2CHec1M8w94Q8uS38YTIZGLtpDmy9LlxqULAmAjDeqCLraV8xw7decZk2ws2ipcL
7VLdS4QCLo7K6N/EBvO3FAyxMSFFJKgtU0GJmamEbNSmPq8GdJFhpsyJtsByftfJ
cjCLaQ5y/75BJ6TT4iDulwKhzBL1tNblesorHvvJjZlfce8bITlurNGjVDDz2SsR
SO7zvQFdExUz8F+OtQUz7+roEYoyS9k87y/ELksvm5A/v6V5orLFX3Bc0F9fmtXS
J0T4dU6oNSMzHP2MzRQgGCR4rGCxCMZmxcptuJTlPz/YNYeQ+xhwfNlQIYGcgzUQ
kiPGh995qrXSGzD56dQssSEig2DWlBf0NK9eQn5sfAmm1PrL0Lq4Rq3UFZLoc95U
oUWqOyVa0m2FqhPxYuqj32Y6bzqZSKeYLCIzEHcTB8rok8JUrQU+dqPCPSylGxl6
ime2vXAqBg62E0Z7DYo40g9kw2cnV+yuI5CxSj7BnKFM7zLvk1t5jsrnruBJuYD+
Rwp8StePCKINcRVMi18Gi8S3Pc2vYtlF6pJ/HLSR0aFIqtwfcOZhcwAe0KG3wajP
toWRYD0i9NsKP4wc5zMMfiLPiaScwrcVMGHfymaD44XAbJDLGFpOanV8B8/2KVSm
5mO0q35/K/RgUWWUCOHyb7bKhGZxrPKocDX7Oq4oNc7uyRSS83cntCmFDW1oL6GY
umd4wTLEkVDRkU4wPBIpT+yF6IiZvi640XXXtYC1RaDAWMhog/jfRRtM+YYs7piU
xUYWzr/4kL4G2ybPvt4g1rT8P8vXJ6FvddJxY/DC//iexTvhqqFyc2vJ2T+226BU
aIu/wG2Ev9xwe1SOWsJAOi+WealyPyrOH02WLnGrRr6goweeDbrOpcmkHtQtAwcP
QWl/XxyF9giz1yCoo7QGpCuXDKuy82ukaLOYRwrdyRKmXxzeZJb1wXxI0fz+BTyM
J78bo6CtsGUC2FPVsy+OYMsWNjyaOovkOiZj3gZbMhpBFB+QzHC7xvZfOEbJcnjV
P6wsZt2rfzC7zWOef2PCZQFFbMphjUvwDvN/cqrsYMcocoCiAawbCCEhvDADELJC
kznZwxtJS2mZSs/BxME+tTiCBsn2PmcP84ShGSwx5RG4cfaEe0bNST0CZMOC190u
jYCCHXbyCE5s+SFnwsQc+dHgpcPMDAcRadMMTJIb7xzT0vIX6pqn8lzFdj0tzslJ
IGDBNscwG41Tbom8xusg3ZzGjfmX2w76XJUpWgkaHPRmL19oj2OlJHlhhatlJ+o8
vjf9bVHAQx1pG60WfvXJnyTho8yieMp8aK/u19glbjHq51a8oeLYf7SJBoGgZmJF
xswfpoGSx4ebnS/U+Xe3Onyz5X3hgiCFCL2iC4AIksUunEAw5lsrTVdlYnb7TdR5
KZJqphAGvtkS4Z/oMj/H7s7Bqf83fmLgvKS1q2cB8gDoT+Doo8r2JRGsim5cFnuw
eKjxtsv/81qXrlHWH5U93Li8Tb0VMc0Z/Cuwolg/738DIqMVboqmqytMN+SnFFv7
n9Lse6o+h/YAUyj7MF1MiccftI1s5VjGWm/Q5zmKa7ZRX4ppiU8zq7JGP57K+TiK
iySguspMYP1vLZphhXTqDkQLiT6aEioMaKXiTGBpUj66w9ro5WRnhNSRfVLgWOal
ylFN6qwEHif/gE5jvWasOsvAoFgGI9OSaGsdu/gKzuN6sEbjGboVEds8U4+ghtOR
x+6mYFxkYIDDSNDN+pYBOerrInLOQXgUy6FOflysGSSIbJXprJgtPmFYu5aaMiNk
uYqUjBc7hzcXpE+xLV9dIoCdWW/XZELtFxVjuYit0c8u7mQEXE7Y4/Q5NjdHvp1j
3g4wKbi/azf5fCf8Xxjj0PW/LopR4UifNoOJ4SNde1a6eAQA4G4E1Qgm0fTkyGeR
aTSzdy7LHzqAwVQEduSGi4OLg4J0q91ivbdNcjpYKkY8W4YFqGmpckQxiX92ATat
/8X3M3w4rtDnkMABEvdw/j0I+dto2mmu1x9IyLZd8PS4kSumyf89EgRirN8eMNPz
cYAl3HZFGJ+ooSPNJydmqXhkYZLyu9EDRyeLT0qiwIhgcPoFc1hm2NXfCbSQSSnl
FZIouOi+8m388xUSVBbzO8/XDhRmIVuX7o2MGugrLnqqsJfqs7svZ29uVqR8N4G4
vK/w+lYQiP08acPAXN6FyOEYpKC6XjeHN87bSaEHWoPK0Aip71XBIhmjg7rhQ2p7
G9HtUChaPavqA/ZmPE95/EKENPK4zTPPSbvZEygfitjq4DZpEcGFpfYXjEsshHc7
tnej77UEeu5pNuhnKX3xZwFl7dGbq6qXyGb8PRusQ5Umwwo4cI+iHnZcG2Buv7T0
UcPbpNwEHkL0NVMtqLNqqB2hRmAgTtesLlAvmsTruJLbJRensJdk1RfFV36cRJlE
l+ZuLzDoneSe7bNFjA60t/VmlBsNf8vQ++dfjyQAGvvyVbovyYvzTk4RGZDZq3sS
FO3zDvdXM6vWQt03ScIWMaYhBN/1tm8ubfPf95PEUedfytEOgxfP+KtThZV28D9g
DZgLSF+J99Lf4B2AiHfXuzLqzOya1Y0DC3AM31WMU9KPQH9zqhLo8XOKvB+5WbCL
J1SSk2GDMy3S+hyXTDB03J4B7nsZEVC482zeAaP7KT3rFuueLMGgEV/FTsP/RFEA
QKg3Khc/rIpV/wbD0g9i3Nr6rIEeXnRZnfdX1cJCE/f+bVqMdN0s3DQGWAsid4TO
3GwWJjxvPh842t8Fq+1fIVyiN9zcZWW53IXC22bVNmRFF8bebJHMo7QRQb0gdAhQ
X4NXJQWnAzQJMQ2JCTuDPI8AHJcJKLQFMkl22xEgXqLV4c62/+2T1Yey1bYml3NI
8ZGqEQ3F5cMI6fSYGNezaWVISGPrRVrBoRM1LTpN4CqGcmorRKmfLHdpMsh1gA9S
fd+uzh6eix0DoKIev52A1TNfYFkU9ky6mpxWGDzj8ifRu2tTQ3kpgqcaRkUSK7x1
8sXf01ItS2RLaZHsyj/bK8cRVhogkQ+0x0YPPlSCWeMyQ8lytGWwWZE9sRlrix2Y
ZAXJofFoIOE8FMManzSRFjpHP4uLFLhoQp42Ml2+KBv9l5bF3myaAZ+d2nf+9HsK
xt9D1MUPr0GzgH48GaYnVfHkOQDiDx2XqyWFqKzFrtv0JDfx1g/GxhtMYFBY7xrV
T8sZfl0ylSjUuvB4jhyc2dlKjiszmIOKB3YuNlPVJNW7r10PDYH/S6e5HkYx1G/K
6tCHFGBzCOWPdn7qnA2/ILDRsYsFszS7P1AQuLXjXj0LZKcP0+Ccu2PaITZlQNhT
OuYpmE4hUrhmZQ3j2ZaVpm//lh0lItAQWhhGc/HSZu4YzHUAbNMHF+xRAKToAUMY
psO9yvPnNWCdN4iw5M5nZ3d7DWcEBT9EZfrqe2zRURK+qmVVUZXEHosrXeThBoVs
TwedoPmsj5RhtClWxi9nXc72TofuedQC6TNia5pxZWQKsEdjk3Nv8Vc0yuuAY1Q4
ejwolYuLqoL/Tmp7fbxEgQFP1iQsMckEIf3xAfhRDdTJaS16SBUxg1z3HDtkU6Zw
gaRbDfDWAqHiJ1bk+zJHyrStgOq1pcLCS2/w9ELYmDaZsKnfW6KzTzypmoCPM9ZX
Vf9X4yCX4OnEO3a9l8Rf11oABszF3inNIrinbl/8xkrq7wQ5uAt8H2cA1tEaFEzL
vN4V8Q1ynSh6QtH2J6F7ocx85VVSCAKhroO/W417ZkX72xY+gC0JDkhgl3xASiEP
SoH7bdcy+BcAmtn2iNiTri2mRsayvLjBEER3IdJsxINJ8rUy2cWNxyDVqOEPrJku
MH3yiAeQ/GzYy9pijc731JDOp8ebjOtIuMFeWIpJ7n0+6fjc/tdTF9Q1qXzNRGUn
qA3u+aPZ3G72WrzKg7keT9l7Bt5Ut5q7pP50qcCi1dJurGis4ajiqvHXjeidgiwl
z1SISUx1Tp8BArQ1vl8EaP5aX+yqxz9hKRComq58lp9xDg8myuTTnA/Kk0VodrLu
TpAoIMgTnr2tza6n6yBpcFtUWaVx4sscM4MUBlWj3idtaO9Vsop3nYAuu9vlWH0A
Ym7PZ85yDpKvtWS7zsBuPyjfDd0XXj74/hz+2HF1Yizhkvr1qrIsb0qmb3kyzc/h
nJXQi0TlU0z4ER9jEvTlBsXA2g2KNmyVie7q7nLGeizA+BfGv9rMDha5ef6i2IiY
pC5oe1x5SpZotHGT6zaV3yLvYalq2ugTJGA8U2gipsA6S3Z3Q2htBJGklVuTz3Hg
pgmjwM1ynTzONKLgRi22fFnQj2OUVvm6IX/iu5Xcn1mIVrrdeyFxEwizXcmEs492
TjnhiYs9Z7Eqf8IGUPMG5x4aDyahQD2PJ6YVMScDCrHmPFf1FsRA8vNI5Ej9sBHQ
YW8zelVRBSD4UuqneQvPJ4lF4/o7NZbGwmwS4rGopvM+H19lu7+wAA0muYimuQUy
BrxdESAgcqPylYF+790PwztXA6/2HuB6KTw4nQkEKfGL90P7zuredYD/mRHdxpb0
h/wnidkcKjp872suiVnhWvDMnOf0hYSXgK5t8wUj67LCfaR5/dtdGqwdXlAIdu8O
/iAoZvOi+floRMIe3GrBLAMlDSBN67hNWocYAS6GFCsUZgxEfyRdbRsdZmodPBVW
dlM6HzZs/vpqjbJm8zRh31831f+FlPGv3PmDiK/KI09RDq6WIdmlax/k7xIH2tKX
SXQc+LSpes0CgUF1GQkpqSIT57HKUBWPim77V1XHQgsdgHNbGu5CLX5r1Nm5I7dm
xhiaFgRXjaOK6aMXms4yq3WBBYqAEp0Pd2qD96HyCAtB9+tf0J3yG2VA4311CGFl
JD7S6Q9inBkhylZhlrHJ5k4UCB/yJsjt4CEOFC1md6Ql4JCR89Eb69VTyn+eV7oR
rPByqYQhHJDOuytufn8CXTb7Mg0NdVXLvSQyz5jjsEF1GmEVLw5js/PScW/8G8TA
19WNxn2Stvit8XWO6pymU9Qeg/I2OaOhjSiDpv7IUnYABD5lFedqdu0aOKT1fX8M
qfTeN+3opJW3d0NK+vKSdHVnAhHqXXJtZLndzLx1FO/al9ZUnlgztd48d/eBJ1AM
JE6edPVkKkwvJU+5ntQAL1k+ypNwV4bxLMjSxC+4s+n0Zo0wjIpCrssKw5kHyy29
ucDUzyOH1YSWPMlrwrinhpmyQpcCXsRVJM+d/1bwg93v59kjJS+hTv8e9IrhKCGQ
FBXDha3o5Zjvg0Xsg5ZynllVLOHkcgy9XIeqfDPFM2EW2DusCfYcuMrzCCEfY5ZQ
Z2hbk5zniWpV2lyFNVdNkdu7umjEykKRXs2xNMVlWd1TmcUwusZGs29vnkVPhpYV
VFSGOBjPNSfdZLdfyUltIZ7OVKPJuTKtjDv9Y9OVaKLSRppouDulbIDHD2z9002I
Ucd3MjezIasW4z7samQPfmRjSShANsklB1EpwdZ4rijwgklc4H2rDKSgmZfu0ktx
hoz1qFbLOHm8m5GJ54/XHu/mASwIH9CW1V/yKQcTOiJ9+ZNPd1Psnqzs8n/C08PO
ICrI/7nLoThepTu3aIVoIx05c/uCygJi+mLMrr8j1QQhhWNLrqR0xaFe79ettGxp
tMlBm5XyTeFavQPYCcuE5MIseE4Xw8wskHyCuuBgqQIxqmQ/0OaVsrBARwfvoBNs
mkGdD0R3bSZG7//GsMU7HB5016AUFivf+vMOiReWbXz61obztByhiUN4cw7+5Ukq
67PBvTcGCCY4/8LucmwvRKcq0lDG9Bv0B+Q4kjjYWMpN1k1MaKmqdCQ1aO41yy2F
1n/24/PPii+AgBfcLiUDPkZPKD8Aq5UA5yWBf63iD5/pwpnIc1k8iY38LrjMlCGo
Bg9VGy/nqDUY+ujdix0GqlXDFk0NkRFumvf7bPxmRVejyAq4rrCHhk4/qyrOt8dV
qQT4wBAAnrwr5MYz7Cizx+rgiRTnHqkfcdAcVweuknyl4/FH7+F7mfpQniDu5g9Z
LwD2u2uun3wo9qlgrIMS4L/ZZbQC+HX9wswx0yo9j7hCoNnBpZiTEz3vQc3C/6fP
ZGQw1ChuuTN1LpzEUTZdvdXau4csxDnsI/e0SlsoPmmr9OBGQLWGasQCjau7JXLb
qRP3uuY04hAEy7RyJykfHppbXxjKyLW6C9hb0lTeCyHipLiq7j5z9x6wktwh+4V+
94BkEdAfcnfFjiTYFAgj5JEweWtY9kISBPKIn6jMSnRJgAUXEqqQNVutl4yEOAfa
yGrN3yuibg6vSAc1shmiCA9DKn6rl/Av7mRiPwH2NRflebGOxro7fJM3dwv8A7bD
majxgq29Iif7/fTnF1doH2uNqxw0cdwSeIWXI0Zm6gYqO9Q1yFSmWEIK+rbFau5h
c31eezfs3XmBcA1+Njm3ZUD2FIUvl236osCn60v86bS/weeBw6JAy9pUTdeUmJHp
URhrBPLzVjZiIb4sTtGAIU4IocRpVS6Fk6ec5V8ecMxPkqX+OJt2/hoksEENqU4j
aGM/t8CIAGDB8BcTboBuby0ty3t6hJ1h4zqGCm8UPkirBBAOQ/e819cc09p6WAnj
dlybHJ2nxybRzdC/RTgcP0/rPLh8DoeGL2yjv20LOMi5EJzcF2sDT7WjTdPZKOJP
Y5G0AeBt1uCvUpGK0UfjGvvcSmUeO/9oTI4CyoYh2H+6U2FKqi2E4oVdBzN02u7n
8Q25hy5kP7/XlgfuzmQCizIikohFFpRzDKLj2eXM2CrUpMfc2ONl7+19CR+PKPhF
ll+bK+NFh/W2IkvLAPGqi/QiIRNVgMj2GEKsCp73Tr8ZTKo+nw+8NSUZpr6sK+Dw
crxqUPGdH3AeuwZLDRTVcjRIWPGRYmnicj+Et7XF8ArSc6qeFOCl6IAa40oHDsC3
03h6XOIlRLoLLYDhT4XysL0CJbWbIrBvEcSZWKGEJowL6Wi5hXQUUdo1srxLntio
q6Fdloqe/H42QP+VTzftoKF0Y7HaH6rWliTYEX+1Et0+DFx/FtwGwgagHdisxklg
r/ly5DCadzPTRdlUvPlc0fs0XYUiJwkeAqzfqqVeGvTMLDasAVIsTE7MSYnXwtdi
ondHX9V3KthkM1qkp/c+ZdOK+tT97Soc1TUU4IB4HIEn4saE7Q7tRTw9xqkidxmI
6uFVVp5gJ1sW7KMnx593IOBFTNPd9KYpzPTwQPn/vHSWtib7di7GLs9p4OOFljqJ
oPfKC21ydn0BNNHTXbxswWFL+oOos0fXV9LzToAMC3bbC/EDVBEkBtQxxSUTuk2G
t7sqFLn3QKCXoUUCC53fF8krVGKdOtd/3J8A4AvCgc6tCNX7CHs2Kk140XC5HcHF
GzrAlZgw18e9IODNlVDhRFIZC/RzBur29k4+reytjC/QD2yecfJ09WQlfTBMngOm
TK8t344lKacYzrY1NgByHnXLgNm+jzLjCZoKACFF2ZrAhgTvC/Dn4KwGvFM4OUv9
wkby17UMKyYUJcHaAQP5T8Qj+bSAUkb1BXhcIuxtUhd8zuoNl9TuivXQX58I+eij
iPzRKCMpuEF/Nwk2Uo8bsDxRY2YRr3K8SMPoJgnc6mZxY0EwoMZPH/jJEVuxMP4K
AVCE+4ZZuee8fcuSrd+nvOubJKI3URbF7Cro9XJAauvHk/yKb7r09j3vbZ5mL/7c
i/W9LZDF2plcLGiIsCvQEDJExcedTqXTSE6e0vBkt8o+AVgVVBMpCHFj3LRj8MJ2
73iC6VgDEq8XGo4d7ZLjG2C2Dr/C8Yd/zUyvzVoKBVSyz6I+MZsEIhNybcflUUUJ
CZiO150YEGwsmMl7Pupj0MfbpADJIcic6qiP4Xnem5H+tBbOe+A8AzQQ84X5ih+4
8lcnArbSLrHaDfC5OBaPL3R2A7KKnKt3UlZcaQDo3x+F40wwiP8JYjygBS7MnMan
5Er8JjVa7o6NBUmRXlL7Sd+U/jHs1EBmKVG00VXUC6WSPgIyIgYMe7X/BBJi+8mS
ukSFSwPZHnEhuXkTHWy+4h4v/5DxzsYzG18IeViJEUF0vKJ0nc8m6K2wgFMZ2b5l
nJeFfmMm5QRsYi2MJkmCSomFbzlarQTLWbHH2sCFYIXhXB2HU1nJnqnFVv+tDq+V
W51m1hys8LTfY56PBqYHjZ3cE9V+p2qebU/ZcDAmEdDqUNml7ub1Q0x9lbtYT0bi
ljGq3+M5XBrfefJ1m2yXhsyYNNWvOkPxVOes7Fy6m9cxOmKy5zftD07PU5wHmert
LAL2o4TEY+ECdOoSHKtBZqlThR0t8fPZuT+E3/fne3tWI9yzdHmJ8e57DbloOGWr
hMIQbNFJj1eWQax1DdhfvvOMMfAGx9Pu0GnN0TEajT8uA8/oLA1K/CGqyoOpIZO0
XzCgnxGIBvJ6solUvw2+FqPWQ+oXwi9iBh/wv3QjvKf1Jw/4JZT5hkxLUAyJIsZB
5J8y3LlBdjnACEMrOEGaaQ6LYGCwb7dRYo8qtSUaEGeIF9e9HeCsOTc8YFfinRAY
TNBNB1jtWSl0yocdgU6S1sG7ZOVEUsCTXtQFH7HI3GMRAuK50KwYGXNWWeQt3qcJ
Q376tJfubpndAVz0GUfOwmsM5gWhl+NtcldlvfWF3uIV0mqbAn1dlm8rgrwY0iBZ
QSVn4+xex9COK16HSIjvLEPiiSQeGQWwVfWvBYvuGWvmlVSZCbeg0jxRX4HwBMVo
sZABSxg1hz64+53ypexJrRris+JpBAxlEe7zFBiwHUStsbpLcuYWxxj5wsvjFqgX
cNK2IuxJ7jQn4hp7mbBW2/XzSCv04Ul9vMeeQCcUGr6W9QWvn8kQj75FcsGLX+2d
/dyZ6HNWCmbOj32uI6hsFkaZxT6FE3zxGGhRmQ7Wmwx9RFDYqjDbmhIzmSjjvw38
4XSHkpRUWbZTh6hBl1164vt2e6u6hiaH7EOPmaYO2Q3UBvdtN7WI38p/fmS+cJnF
hWsQpLKQhiKyUlP7Og1Vp2TEKqf/rAMfsKNKFvbuwKdfbFYL5BsM0w2FFtX2ABI6
cxCGdw89IfH6fSKF6bjWYjwyQEu4USVdCYenYYIuf8iPFPW3BfsL+eExzSwiEr0y
MiSRUHoTcCYLBrSTap6eB1ycQu2qxhsPfbjm1ScfX1PIRejF+LrWoCj5HbYZvCSg
v0UaBeOVYExQH4mMyTY/tzDUlvt/rFBk+hBihcyHffSm2MYpIOkCq0xuOGdK9stM
dVDKy4JUBkk3RpeQtH6lib3qLfl96LDMku5hFf7udgVkpr6SnG3U/kGgg2sDyyr2
cP7LWw6xsTpM0i7TGD/uLxiSpVEn9O9z8+P00ylR6bweCsTqmx36UJV988E54kil
d8g3++zD0KbtrYNtPWPpI0EOQKwX94XPl1jYNauThLx05avfpF8fDle0KfwymbID
Rb7CX5/5CXsBdz5Qggb3lfZeX569yH+T/wUHfqy2AaBeAAuQiHNt5DZjdMu24VVz
JmKCrLeZE0O0oTHfm+YQSKxuREmfeg+TwO3x4sNTq9YjKX0y0FZ3embY211CeQMi
VvN28DebTG1/HrsqDI8GGfnAhJeoT8lCXSw6HEg4aMPihjEoYH4hKNct9tOsY1lA
RIf4h8XPLYKAMII5YvqsbEsf9nvFDTKfSj9y4JHYjhBf3mahWJbAPenrPcezShTL
llVKC8ola/+vrbHWJegp+04ehxt6ByjjNyLavoPyHI3lJvgyr7+P9EgQoBwcWMIG
j0bdCIcRWpM5g6Yh1e46Kdpxwi4gBez10546PgpF3XJTy9h8JwqL8juqG7wxrbF1
D3+lwiY1DkVmucR97o2Vaf2SIW4n92EMn988LTdkydAHCWRazBQTfZ1SUcOFCy54
8vCeC8md9gLJwAaFELjz7WNfvq6INI25GmTR+kxba8W304mt0R7GgL7T2W/2kb/L
c/lbH961aRiKLvcNkiVv0VZza1KhPJ4ZUdU7I3pu0bW8vlMKEO0BQlVBlJY/aMJy
oyhrq1BOV+RNZV9YAKSbOtAqmx49Nrz2pOOJTt5qukQ6LpEKVy4iwzkGNebKIqyL
/W5bklQgh4+R1UgXui9nHK5hoYuUI64TMsrYlyhYSLgtcQcKIlySnQuvGPnynBM1
5YzfN5AEXwNALyIQKncJf6acv/jNN9AIk5tyd2I2tobdP/zbFFoqlQUL4hEGUR/K
uZf+66IZczDHaHkybTtk/2bNcaAtQJKRJsie9rLtlcXeFndcOtCkGGBaXYccSe8a
JIYksaRvA79XaL8YEj7WvdaVw5zClXU/vgbjnUPiB4ps6Wae+IuY3MnbKSvcpV7w
SANTlZ0m21+ltKHQPw67+8wrt59qfz0hHQmSAf/FV844MHbv4ZgO20ND/KZB4bjU
WtEjXY6Oda44aAKlx5tHxGsQueYDH0j01k14oaHQaKJ2+eE/5XQ5qTxhqASR3YNz
U3R/qFVYktwdZhJSJkr3bFaxl4ZzJoZJHLdlsuGTN9x9nL0BzLDFscUrGC6n6uwG
j4OPxuZGLqXcRrQMLNe1CK6ri3jxhq61nTuc4TUVWzi/XwKO2eKSn/Li0TMihBGG
jhfvvAdpjQMiGe9aaDHnySlG2ZfqVtRDmDfIhDrwsjSim3eUxwAM73oB/Cb22ZhS
LR4KbNC7jDK2EHnkBSbppFGj/Jq36JGCYzt37QJP8OaKi6CFg/eC71iqJ4ON/dih
G52EZtpYiMhYbl2BeIgwCphPHT0RBFw0J36lRHQeL30hepDZa0muFTa2pwTSPlaj
AFlN0qvi77XYS1ZJezuBqe0Yh3AqHFv/2VlpMMChd4eyPNjXOp09qUdgSLT7K5UR
qqtdrwjnw90bUNqNl7ipOilEyGOZ48pFCTc5LUpwrWGxZWGpurpoZEBE/mo/nOJt
9WYyF/GFrkzrPN9El9WCidedh1Dtwa+pd4Gl5zeIoE0gVXEmv5yzBWkwLvBVkXYu
yoHiSazG+wVDx3y+aNxfgU7FgnaclSHuaieIDPwb3nT2/kOx8/PthLrD6Lk5dVRY
YW1WGJuFTvdFLlw6CpCsIWHe2U6GUV56+3IR8S/rfWUP444Tt4TwhsX2M/fQGqjg
6fHAYxYu4ZqCv7sqt8cq6K7WQvnbLqIMO/J6tjfvm5x2F95dC0jGmJ+gohgozMlM
rMhiDojwtgajKgu6pEGsBVkYPY7ZwQ2OgsVjjcMFXJLQ70wk2Rl0ATi/wQRTVGdb
q0NFcQ+x6rZhKUaqXl5XQJLwwai1fTD9KiWTFpURm4gROr6KBYEcLmih5UOcdTw2
t7Kri+QCeJ9EbCGkdtUgNVDWO99WBszSWMhxYrqX/ZDwS3ZJZcTmNK79JWznfb/a
As5DkbV4sPZjS7bd8GAzqhH5mAzave9BCKBidBlL9S8shlT7b1/1lV0WgBnB7riJ
gehzT4x8NminB1RNEUtE+tUVOXF+UhxPI6DRBu7vxhSOXguVIp62/QJNPy2TokDO
0CqGHxc8scbgubTN0fMWSu+6okIouWmUMIVh1TQEAO+1UdultlLEDGI/rJmZSVXE
rH5Q/9lw3KhYVFXkDtz5q5nC8F9COyr+S4QbiOVwwfI0H6uPPLMoGkgTPCYPGrWM
V8TBPCqEMXNgu6sXIBs1fqVb5LLVCaEsYjReQklkKBJAZIH5iWLuVoykX7JOgAxT
u/0aFqNWHnc5BylW6zMNbAxNog/TUVzB9ml3baSNldCdpz0eg++7qPCMtcR1t3i0
yiAZ7wPrd56uA/iEaPAQwwZIiFdOhfLubuDljOZjVxG8575Tc3ln+od5ARJF2yXD
hDTyBYmdb84zNcQsMKR13y/T084bPzqKl7CDoFdtLy1vRJady7uMSDM+TJo8YV2E
C9fKPKFqAHD/sRmrKIecoim+AtIs1Cdh+ZKiTUpW2p0EjY4AVpZjdqEOLfMqn/j7
ahI4+8mfZTWinrg7JbO2JdFgvHg+POlgMTvoRaxqQJfetvSl++0Vn7fWWKm7A+BN
ogELFDahTDt8c4F8yiyNF8RuyoFY/oCKLpJNKMhM7Cq9e88febs7Gedf0iJHnPam
G4wvgUTn/QeM88uDruU9YnAEN+kiFHe71t6CVeKNtLJNGmgarkrvBuO0ODIc3y6/
EbJF+INxPkxBw0y1kbibjshAHh84KCgnPAI7wbl1DcmxLm7XR3qVG7E6NMXU+td7
50iaItMjNAaKkmnG1X/Pjr3cudFgg+VIqRSUwyYfff3AbL6zpTAV0vcMOrdq0ep4
dSU/6vAInxukzlQ06+P+cG41gbGduR56FkJ/GSkmxd16kwvj9iwhN389p3ICwJIf
ZxfS2bPm/6gOVdMS3Km1UtcePS65K2jNsrbBkGVhcYieNFooFSRtlC2qZbvc2tuh
85uoIFqgx64LkQ59LnVStKConSBywJ8i0+zNbkBE97jtx5Nk/IoqLWmdoDf6MEm3
UEyBgofozUmkfhi5IsnmzfM4SW/8KlZTTpSxUPVSxOfzHeYcxBTevSx/86DRg9Cd
ColiFRX4yWBNY1j97YXsltcJAremsy8xXOlGakjXoP2zH9bREeFW47cei9xNcM1/
62etVYSlRzIlAFFLW7yTs3rX/0/mdfR9lEi2btQXgGIUY92Y4GtWeQ+ZB6ftiQkb
oOJ7wyEC1FVE7t6vgGkD7CguzNQGrK8NdqcbQ/bo19917Wzen102WhA4eTB/yEOn
plDKLu4YJc7KVVAcQ0RXA/DknzBCXTVM0yy2VHTBuN8FJ2XeRwURbU6N0GUOHv5O
TUM/yY/k36AOsM2RMvnG6khGBB9/m1RV87lvaC2wGzqXxxcYTkwytS70F6ZayIMX
hliKiGGIX0TIdCeoR2dw9LkKoMHRNM8maN+kgIgq+L+ZOy9NG41VOQkBlpn32lHP
IeVmlyQAxZ4pQVrnHM12tNxuhlS6bn3bOf72cQ2m9+h7QxLJe6gN/1bMMNoY0w4f
OPpXYDVp5Q64Q1OswvdNmA6driJeiYrYN5vyQXdjvkStOKK8EOseUAGDQJk7pbpw
hM+s7xCjUaIG86GhAQSkTid+jpQgvObWFmiSUFlN6kDlRFSpI+JMkB60J196m0p7
iCg/zzSA/bgbL/vhZHCFo0rLu5e+rHvQ80/43eFV8DomwiDGpPoQno4QKlayJj/C
tahR0R7TWku/H3P91qqHpCtE7IfQx4iljojx5N1S/4Cm8zEAYmw9CnkPVLhyrkmz
9HjRTRRG0AeFeQk+UkHikzRH5V8yi59cF1pUzOJZWqBi8CtUE1eb+HQJabKWfJlO
pNxuHa5CnKilSGo3HwoV8bqtIft30KDWL2b8Sv3btOHTJbgwiqhKptVQCq67DAZ1
DkoNR/GtqDw6pO61eCcF0vRbI3DpSmwqfpcny4/lbAcWynMPxV83tGE1r6bgCBcS
XIVI6gS2Tk0pUXFuJCs5QjrnsZp+zuNwVD7pgVWRFfK7bMUDQdFRmD0s7P+zdFYg
4mpWkG8++AaW7231fm51hiv2c4AOiD3InSe5JfVK2ThcprWCry7/V16latQcqxU/
ORI5m1SNo49JfrnP499fXWvIRUzcxDECPhliJqkCVco1kpWgXhqFS866pOfG5/kH
/uGh4+61qlvY4d6JUIadztgT0d5xz4E84Tjg4/I7jX5MSP2Ve+njYTgHn1Ordf1m
5Li/FAVncRXXS5lDbItgvfDpImfZI5nMLsKtLXzWWw42DrlZEE16O3B7cULi0Bpm
3240O2TdQgRv+7wnWkbzVZN2PxF7VrhQ3xntMl/XAkTdIlLtbJlwHPGDuAmo6khA
FjrFTa5fx31MhqIINPDa9kWSs1DDByeCOs2CvGnREUskzd0mOH4+5y62p8x9t2kw
tYRFpKzZKLfBQLeKuszqYOKltHoCPwqPsq1K1lEd9hG5WHm85dEaIxbm6dy0krff
gRPsO4W0/biU7RxPGbRwJQCSYEML4sOXkf3s0NZn/o5bTLRng11a3gkaAL4YQ2wD
a/UlX6rAtFDBIRhEnzbcuIx55bR49/OiViBD5Bq7fspm8KHvNWAEbuEM7oxLUEoM
A8jdy84dfiJOFjIKkh7D7ZgePN4RnI/C0ZjQn/dNbD/3LXv0/s25RYn+oAXhlnzG
Za1Tgt6/SqAtoqFNCL5UEr8Jze5xnFM+vZZyMQaNhU9w+D7aFhZqPEjd1/IiXeh+
MrHXXwJD39OHixflgi43yGZueD34YtlbhG+C7Gx4BsY1ZoDzXB2nVb+/PkoYFWpV
JNnifXn78b3O6W7ajygN8edt2xIKZh6bRR1OL4uVx4KtA6ZIsRQGGHaeUm/kJk6B
+CosYk0sUEiQgK9+6J4sJemgd2HCrZpULYBpSAx8jyC7LDyqcRfXz42/3g8neh9U
9YVuKz/9aJIy2f4X7lrYq47PY63TVfi9/gTEwuiUTI4wN9btVZ6lYMx8P3QJb6ii
n5YbTsh4o8JrW68GLLuIzbNF9Ry7OJ6ApLTEdfprj+vaZsLBW8HjJ1r+Iiwy9jEL
5OLMvIgeM3UasawOS1XXUBxOD86Bq6nz0dICYzGQiye69fJ0/p30HEi6A4Xo/wnd
JIwpwjRPNMhHMhZBXeLhnkiM+uLO1TOVt5HK9tODfCIPbOmpg+OxC6gKREKH14vu
LwMwZqr/eTe76pXvFO07+M+aRospQaQtAu+SbBJzZ54sSw5Be3wFifXEhAdao3VW
X7Aj9lryn92Vy8vcHtJssqwXI8N/Ca+YWMON7a1PTZFFckho/1+Br5bWZg6vZus4
sNqmYw0HBJvarbFcRslpYcZHYdisi9PLif+WyRXsEHfRAzx8q3xXP7i9LOwXMqET
U1bye+pTmVa9euCISeIDAlEU7EdCNJ5ksxA5Si0Abz8KLYwDqrYOG3PLr+hXYPmK
GNco5miFIBhOl4DBhtKoUed6H8AlJYnuQJY4E4xf4w7mjDX7/cQ99RafOGCrDCRV
QQurfETneHugrN1I6VW/ixPibDiuuD0ycVQfnvvux191xcOg3R2OSu2EksEysvn/
FM7lS6+TLnqxzQGJn0pS6+bFAcQZC4Det3A++CALuAGm+cceZMHAE5k78KI8Bjfb
tUwKG2XFeyRHR3u3r+2VsMwns08ZlMP991Rl7AQ4ruUagYPL/wfDtmBvSGxT6Gr2
nvNCx62xVvrw0df1oByme1Pm5X/MpifgXYrWkRkWTWng99hg0BAu/VP4aa6Xo3Zc
uFPuZaDHQvXD8nGCxu97hddDReZfzV4H4AhJuI5TqfCXkY9YYAVTkgmFSmtzjjuh
PmDpazhZfJrhiDcgAHvx8gjjpy7venSA0FEnbUvbcrT7j/c7pcm3/OxJEcig1IhX
y8G2hDYWjZ3NKgWXJejtlBY/xB16BOqH47oncC+tNuIkJBtfZ6u/KpQJui7ojN9H
y9itnFptf++q4jzRuyenmwsnbdU65sikDTKXQ3KmQrYCEQY4PXbdqS0q5nij9tM5
KLKT0IaRqzY9eX4EgcIKp1AcWKAp0HyKaOBnVy7r+kwSy9pN7xN4w7v5fsmPSV9L
tEUlizjAKsL8YZKuzH1iWnvtRChXTWGo+gRWZB4PNv705KuB1OiV6IedNvKZMKMZ
FcyNclTyU3AbH6wLieXGkEzsqGIzirveGmkF3LSzoGuKvVMWosWHQoLz7NLX9tAG
BW5Yl61TPLts5JJmwVGpjSUsTA3UNRpZUi55LtV/FXHxJ4KZJ4HPmTPOYpD0LGaj
TXEG1ijba4p0uM8DBk8sl1naOKrsiIjSezT3+60gf85W5cSzWnBqcEOSibCvgI+F
8l62SYnFBvswVnGC706OYkXpCJmGzLw/cHJSXdkSWRR/qFbl+3Rc8I7jRIlcugV2
FN5+gI0qHETExCENKmVfdavGoXdfEzRA+hY6uC5elE8p8zyK8F6tbSsJ8ZWHCSvr
5/miD/gcj/HEZCHRhS/ymB6HVjMoXQuMpgvQQAjRoZ3O1A1fBj9oam5QYMG44gBX
+kMWAOG9FIwm0aRSp/4gzw5QMHvKoO/429zXpDta6i2cuBdOo8hZY4Wc9K/ZBghe
ITNi5tEvJsT/Qxuk225hvNYQXGcJf5CTjE4f6hAy9qwEi/8lHwpIvzON3ghok2XH
GZNiZ9uYBb/s+UgLw9UyrnYsSKZ9f76+j/MoUi8XxtNiU9PyVEtEZ3eET9NSfO2T
3WiiCWHphhi5IheQN/1Vef2hnnNrtcQzBwrzIymBgB/7lHtwOfM6xdFBs0zMYa8O
uNDFH3kl+4TWL5XizZqbbx8CgKcx9s38H4WuApGE+Cad8na//bxeOg4ZgJPr1Thd
O7SRcRRKgDyeE93GisbujIHvTdAVpNQ4uheJne830g3x2NrFFWjw0UK2pR/Ui2ov
HJu2Pi4CPtwQGNKc3Pi8+NxKzNR+134ea2VzpsLrmOMK63uJYIrChVqOt/NA21ph
PegYeoZWXOsMwwN0erEISWWZw1IrOGRdg5FmT9sgk1ySjY3l+lvzfWAMiGi/yV77
sN0EDdw+lruh67S/4xY1A5hk6STbKtFQGH1E+uvRw1aWqSdOncc5Dm7YozAs4U8b
kKLzcoVLqSN6Jvqj/1cCV9kKa9sPDUezTUR90zNg0JGACb5kMGYRGBwHvAi0bRmF
cvclSLdcoS9irUCvYK9BlEk5nVMuHIzz4n0C9L8WWk00ssuEKlcemKTGOVRa3dsW
ZQqSdOaSCOAi/tptZHz3MaX3CBHn9O3S/R8f2e5oLZyUVaMVk0JOpzQnTNyhv+UE
rPb56YOm+InY+BQ+19FLV+hgb0LikvEpA07Xr2hmrVsMRbhuhCIKF/oksu+I94VX
TWrT8GPUSsZxlU20hj6y8/PAcsx1sFHeS05c7JiiW5u+Z4z20bk9+TvQdz1S0O+y
kvi2wj5xtmf6ide1pWOmWEKNluA4hGtHEps3aWpVNbN7Pyi1geV3eWciGCTTsU+A
OhJlEIZ0ZSQXc//G8kIYRad3vcsS9wz8MzNU7tQDOp/P9MPLAfN7qSLEyAeWl/cC
C6Nhx30QWny4hlo8klASglMjX01ATMGIzGveRItb6fy2GEmvFa7AEroLDQOdUwue
ettF6dQY5mHfKlkGyiRKwe1tx4xW4+C0eRuIZ4SmehYQLdfuAC5jc7t8U4xW1xOs
RQzUx3HAw0t/+agMAMjem+kftYbTzAbcpp73g0xxvfW+h7lRxoGrD8O6170nokgU
f4A/CbxE/EqC8rUjCdi7xJLAluBmPNkyioc1Ji/QkUxFeA0siAJA0ob/BNIsGZHP
6HaxE3TcqwsQWUdtODr0s1fRB0VHiF4WguPE9imx+CVvNSfLfALZCcOhNdhebQXW
eZeZYpGaXLum4k8qu4N/xZSc5AR+HLSjDfBUxATjnalzX4oItmkUaI0rcE32PDEY
c+VMR+MD/dwc+PFKt7SDsCdLPSd9JhYtZ7BgDm7lSZEKhxxNMbC1JYXwxIlt9Ico
gDwReS0ZqCj8Yj6wk2LRSWYJPFWu/Ieu9F/bybtY19WbiTzat1A88Gc2VR4hYS9W
UcxvMPEoy9A09KuYWpojP0vmZUHbTAm970XTmQEh2Seqf+VR+2dDWKFFQVpa52hz
5yf7lmdLgB7Ydoz3hDSdopeEWxGPheUdrhd2BAfpdmBDMYO65VI5f2Pzy4XOM8dw
4SRi0kzeqbGwlrp//nRzLkT5BdIJCaEH71zpmLZ0QEfVltYnJfFcsADqXB9kUTTb
hASEWFgotjLR0n8h7/mlQDLLLrliLTMlDayrgd+W4MVTeNcgGcfEjqp0yLALvFj9
E/yWPXrcmy8iCKA308eauXOx4RNYJdXG1KBhTcNbejK2Gnxy1ck1LAXVPsVeO1dM
pUw2SqskHgwQm/ugnpvxMsgSkJsq43cHDs7sJdjT8X6zLM9QSKS24xu4qm97rQIl
VVX+vz2LHm+nBIOo1N9CBizCYbJCWywXi+g4+wnfIk0iyDsJOfhCVEfh0avyZmv4
O/WWWh1XpJsWB0yt70L6emUNCkQg+1p0gpw1rp6F3AzQ88XJSDKgT1NPckYqMAjO
TkTOB2Ity9ufHbleDnPbmTSVHmecK68tmfO93vHV8UU8aimg7C9WRW+vEHiHywKx
cfpJFkgeN2tnTJe9TNEjFUcG1jc6V6IYa6MfN0BvceJrtYFQLHCFHmyW5wLlV3Mx
2bMdGCrOQemdtIgiThSY2ek/mGn2tqa4EePShc5cBvLxKm4tdTZ4fZ18LUoUUdGE
GM659dB1R40HpSpi5j/ly3S7EGW5IHlCBmGdKrh4boBqTBCPpXIBf2hg1aIOFXeY
uZGE9ClyulOB1GQ1MPuMWI5v8dwG3o4SUx2+L60ENbjM5wnYiApHY9DEHYmFAXQJ
TIsIb7NLGkB5+FLd8k0K3JDsrv8CnkM4QxGhFXCoVJjYfl73dnqR6sfOaW29U9fg
srPwkPVqVZTu4yNf48ijn+spIxbWjmeHBNyJePnl3+fP4uRIZxebwT/QkjkXKJgP
DZL5an6TXJYaZjj1HqfC5vkI62aGby9EynEN/AOu+P1sqw3ZHRhw8VbRHxBKj8jQ
jJMv+aYl4VY+5lr4xTdE3GtR6KoPBoy0oPAj9chKQMatRb85hslV3BnMHCreEs3Y
PmxiPmHglUG6LNWwFOCoPiv63ZQXBmzGqcKDoexQ7QxLOTkVoX4AUui7tgcVZEK3
32Z/OkoqJ5BDncRPPLSrJrSiQQwmk5aZg3YKI0B1k3CAO5vjPAwKz5osB2Kj+2tW
9vjlAL591rDG0H29XM5rst1bGe8JzPAHv3ZHT7zbI7Y/PgoRQuaM0mNVxgNPRzkz
FCAIGqZFzEsQz6BbOdX0CEBURoIVR8RNoLB759588+4iB9M2WjFO/cHrcNti3H/s
A8+g5dS1wIVsGNOsw5G/52NHNKkBA6gB1bO7t1VHbaC3dFCdSC2MdZLKdFZHGCjn
KnId1+5nSdTQTgjlFos3h4eGKcBDvCep9XE9hvWlGea4jfeZhTI76mfGAgal8m+8
Nqj2tzuflodYbbNXyFOrd/cglkYJGwCBe88T/YXLL2w2n7XQmPzD56LIVZLe26Fl
S5OYZIE7P2BIQ1gmhmApYt9+M3qD3xZqKP1tTmwas1fqTSg1Fu/6AyV7OamhJ6nG
FLWkAUUXM8DtwN/1k8RsmSVNYU6NDRJE1oC2Y5CELNKBpmVOaLaG0qp+lWw5iOgj
ThuYnqs2SPBHtzDrN7Z/e7/263Pzu7Ou1lZCj0u3xZUaIfMIba/xPGEjsjisRWG/
zspMsNBu+f2TIsJCuIjoMSxfX1+K4fnLa0onIgIBlEHgyo8Z2yn4pnIARYyZBw1M
3ZdZbtVncdgVACmq0pk4BglJrnRZrLcqh4C7HF0MCmpx7DaZR2D3oIGsc/YFnx6i
KOkZLuU1A33hH6YyIr6JbhpMKkwzFx/VXn5u0SLD9M29x3noKADXDei+1XS8F++j
M27m+wMhwfW4nrnbPLJbp4uvjaoLnTnVSQ51kkmDZnXnfpeo6Q5gWPRN53T90CwL
5s6ZQCfppHorSt6Dtw6cGrNQhfIxfg5+LZ3eFugSEDv6icO5HUOv0CXVVcv+mk1j
WgjR/qPRYldrQA/IUHcACqIOg9ew+drV3lrXeqOuq56dq3d0GOpHCtHBMOGcMRgw
jTf+Kz7FKRPuq320LugsN8p+xiVIUwl13AeYuqgZWX32E4ltetaRAr+c19tZIiLH
to8nCfA/pq3flWLDiTIYhZeJ+T4VhHqmjeYsqK0CKlY+xCb0NQln161XXLDM4IUV
9L6xFW4kkbctDNuSIXho8iFg7Ng90ZUAru+AesKo8oRBfG2UIgFNWpFlRydl77XN
aEizSbzP+ceiO23kTP29ngK6DJg+QC0aBJibTKzRF7LGm/YYSwXkg1InRNHth8ua
/Q4G6Ptwn5kPhKRF+H3+RsBIqjIuL7ziCxndGDpRuH1HuAVv1CC0rPA3XN/LSBrM
RT88UZzTv9hp2Br6zSsk6Rq7CB7bZRydWNSzf65uJQmt83ZlXGXhseDD7jFlMDyZ
cS/0H5ZgPzvwZ6qWscMLFe8flTKM988zoGP1J5MfbHNSIB/xoikd8ckRcSmWUpbF
gKAN7p5t/1lIWp77crBySBBl+9e63i/F+vmtT0kjvG3LUf0PfASTjijjqd8RlAFH
gBoAmJqPAGNv4DqoRMB/rw1YUlDGRhIpIeYNjzmskGddcAA5Uzk1VzV1mIR1XbuB
NmpuW55Yi2fZMiNNwf7+/TXvGTMFfZS//cULXknzDKtk47Jcm9LrhyjTWGZpsc6u
jW/UNfMaNum7zhE/USwt1mOCGtc4t2UhRd+fOMjF+GVLYpeb0xnmucXmu7KfWqXr
Ok6p1K45mSUsIa8Nj04Yu4GHH22d1i3xLfAQLEc4vnufSm8wyD2tLqSoJ8zLkEPp
xZtj9yB4y+y2UnXHxUSTufqDswkZi5QuyjhZksU5/ByrJmoMHWw+mPyRFFCa9/CA
jXExYSu5vjZyRUUzYB3crJPdA6KZoPzT8yWQ8vsY0eW1bgn7GXkyUyQv8kUdUn0Y
vMJsWat0Xk1f0lgoOJxhoc5ZIbX6n1n7hJOqSGZEg/ljT3zRo5QECXBrHtkEq67y
/ZytMerPTR2jpsQ9IamO84Hcy5aJdMVcDtlJgKRjJl1RSfAPTIOlnCoclh51y+Yn
cD57S2l7vlmSKQgH2RIb2zDmEFVhVStEBllG77tCiHA5tNhGWiqfagKxjykPClIV
2ijjbSBVIY8s7R1CrIWrA0QEgU8bRdyonfuBCL2ooXj6W2E7Y9E8lMf2RIf+xbnj
rfDr0krXedMcR9Bkm+jaZySTeeT33k4treUhL70/EsowzY2tZZyR8C34Qaenly15
+wwtyTldY8Nl5q4zJSCIqmNCJyUJ0PaxlqqhjFMCqQV6moxJSZb5GIKYLneVX5Jp
Y8vPeUUeeoUwimkXDLFKXlv1U0pTz+jT1GjduSVbQjWpEZ2OMAhqnG9Qj2YphyDs
OPymo4Ga7XGPjKRhSsviSaDqDBGBKbV3MQI1dHrZpUomkIb6CyirW1p0W93MWXUM
nRvpyvGvNECE7sjbe003Dqfi0T1tNv3zW/TAve6i1kuNYd7ej6FkUJVWoFaZExJ5
zdGt9ycbYYocxpGL4x9gdVXmon7ioVAff/n311zAmR4nrwosprxPfZ1PE4ivnb7c
bSgG/Aunoa5N0Bc5cMvMDS/sc8iTq7crNHt90PqS0OPRLHUwu9Bvkz9rjGD1llbf
0e9iWxPDMXpZRulwp+TuKvZvxZcQlZYrJbLR0GvPqHl+SEOIMWbHQrr67/ZzcydI
D7NaxPQGafbPGdte7sdlQLhQ6PGH9zizvjGUAA0UvqNQUk2EetveEt3J/pL1f+2Y
hoDORu5xKHhiGoAI0jfHIkSETRR9yoGoFUklzYAchvS07FIHTJvXf8CS9Nmn2wZ8
VWOEM+H4Uxdh7gLBA8wykF+vfpGulogD93+tO9ytfghW0HrkqdOolH2gKEu02xMe
VuM/8rp1pqCo2qxRzRFG1sTBONfbFlpNN7jqpMUkQsL5dnmTCwcTt+85ATQ0Da9H
fRUMohn4sIGesO4CywpglfqInumkoU9EY8ZdYc9jYy72d2Q2N1cGEYO9HtL7wGn1
1GPZpF/NFV+xLRDRTcS1qzArwv/ZdGlnjCoHTD3abvCYHpwS7Dvt8gkbk02bvigw
CPT7dhWICUTDwybVq0AifWRSJ/yjkoLdj89HlB/2zpw6ntpMzD709UXZYGFn9YbW
MetlXUgg0lQfuiNc4IBK2akeJeEbTQBDu4trJ1s+iu4kAdNXKhwnmJ2qBVkrD5AS
XNrGbHg13DsLfRvm7tEtYX7zFm1DD0CX9Zt1RzYQsugocDP66VUw6M3uOfTgn9Jf
fKjx3xFSOIyGtOJLu1AGh1UOsUUbDAd9PThWys7pjxX0Vg6hC9vMvBh8pV1oLypD
+VFyqKO3i2gTQUof8VvHf4I2ptwsZhJFhXMBX0OvqUlWPlfRZ0tLaejqbOi87GQu
Ar//PFBoOOb6aktQJeacz5v2+77SuwqzGSs3OwnrbYNRzKfnEnFi2e3kc5rZtCIi
XxhXjI8F1dtK4aKlxUXMVh8bhUiKr0t2BqQZRM1Wr/k9gvBMw4kDXACjHkY3PSSp
2ga7PU5tnuOjwhvfTqVExJ+oav/2wv6YUdSEHdMfJU8ymQt77jSm/uwPVFlMkaxz
igGRJYbL7hwWzfB0+faB/3i+5NV/2Gc7S6uHVj8eTQINhoAzJYh0jzFGbeuIdwf9
6LD4RWcF8fNUfzLWHrSg+l+gIGYxZcUTs/5ZJcdaYugFoOmVPcBsEGB0mp6QTdHy
e3LP9d4kbBDC+4Cs9RHXeY+TTyqgr/4OcCLgNI21aiII2NPxeQ4X/nUU7f1uXcg/
V1eWy92iiLw9jIahaPPnw95W6x/ShatITUDzZ9rj89TMUw7rqt7Xzsm3TRvsu8+Q
onRtO7v+QwDHrN5Afu+8mXnaysnGiNnDiWTEBlt9oB1Cu5SPRBZ/Rg4vww8RU7+G
zZjUeWLSzHTzC2rgKlz1dD2EJy6rEnVp6Bd+uUvWlRrqQHsrDwBgII8LurkySnpN
8NkTRyiANwmpjLcfRQ9akGyQgb7fBQC7n4cIBgYIqH44HEGJvX3AioEMCUg7ZVI8
MPIM8DNWFhl06Rw71AzdWsw48FH6ZdLHd+oWX+AR7XxHkMhrBQNTg9S/Bv8ZDVvm
ny/cJIAZHwD+96k4Z22sP0Jzn8VDZiycieErHxHeWiSYewQHUB/LHeZ0gBBMg7jY
qhgNcw7CtTuCYdXffZd8DX7XXSXZu/BNIFwf6qua6qzrgG20O9Uk4vZivujN2k4j
20oA4mkAaoM592UvEEclUxPslwvrcz0EHNqr//+vlFvyu1Xbq8BHQGeXXK6xtF6x
LrKybRItF3Jkf/b2Gy9JvGVnn2Sny6+tCo02P3DzCQTcIVOP3gSNa/C8z4v0EZET
DC+sf/lswLlE9t+0UnmZqmxOEdE2vYy4lcHj9+b0bXhNmHCwRb+Qjinl/UNooHoP
jIY5It0RolyuiS2QlfqH3NvZpN8pyq+5z++oCHhQt8XP5fWmwUwrb+5ajbD2E6lV
uJtQ62hJ53AEFiEo95pm1kz1WRG/cTVYtcSb7TYnj5NIAjMUGFcpG99AgGiprXso
rpbhjGb+XhDVhh3vyyZip6qNGKNQ1nZVnUqGDknNESrvhvhZ1GA+1cqnr+qoFQU1
Bie9TOve6RTGgdUkDfdkR+I8lJ4lLw2+lx0pw/AOgWMa8R8hVLcUPzqTBkHT6sTC
zrrbzywls2YDNsGDxellm0C8VUmktO3IbVnZff3rKD/kRlSR8QeN+s/oFknrfdel
8Vcko/tj3p8IabBFdp2ALaDEjSe7ZliuJfZVfGAxNhMfaVyQIKgkzUuNvi7rQVfZ
jlC61GSU3TScXw4KaP4gTbEXcwwyl/5GeefjmZqcIdCjr67fQnAMWoRhaHXNGG3X
BKRZ8J9sujUHtYe7mivJBjASX7xFBaQEx0qnmEKbO+7251E28wyJtplq59wzukbJ
qIOBdP4GvNbNl649WhUyi8O7p+cmmSJfKPzCjIO1G7/9rRt8BsSV5pf2kwNc9N32
nDvmtHMsgNqDzPRauufRRcZ0+nwUTs5ftlqlMlaB8xaMj8V5H1Nf5hSgRLxrvSCZ
dh/7oK/WDfFmMTbydA03t70nNkKG+IWXRWbqbEhnC+aVdMMg6s/glKsRFPkZOSpk
OTDfy45+BrCT6JXF8pufWLcczrM5KlpHemlBzc1J/b2Ld/pBGUYphvxiN/VzjReV
ZP7KE41kUY14SMG17R2Q4ITl36l2leNMcb7IrfmFHEmdWtaiOSSStp3X/lmaKF4Q
qwndtakF2Zgr+nwps+NNxXXRvgQ+PhI+pKXgPPHTISWKzz+rVKyqbppBVIEtaTDI
fgqRhOQxoKqKV9kku0nV5LH2beLsbgZvMTdCdzbzLCzakkuaD2eiwuHs9iqiAcjF
O6xRhhSDqSPXsibzYEoDALVxBIXl91lj/JzqouSwfiYDOtXGeYXExiRck75pCwqU
Wm9GAmnCANjw4JNNP/dcgVphyupw6WJM++QnSq0vYVY3n2q/ao2C1WX7l1RvQAia
IFZ2hLeU9Tw7qooT4oHs235KoSHcAulFE0ClvhXt2/uesaRW3hPkmlC7BiEh7TCx
WWh/DPrX+9BvFSfRPy2X5tNBvR9I3m8+ucdf6zz5u75vkXwXAYQz0Dh9H4NOvrVJ
m8LLaCr9XNTlBeVegzswBe5PHL9JHbZ1s3zbpo5D4LNCZaYTQLXozUyKgyXIwPUI
+xapeKJVNdJSbrvXkQWbR7LwjVdIpsbgoEAhAaBITT4Sy4XdGABm7btQMy/fa0Q1
2l5LMP6Cgfqn2fjq6R5PzYN6UIBcbepPQ7xsDw5ihzsUfPY1AKhPeLyTgpsZwzNG
5Ig3Mkk4qLUGPVbX24Xk+tY3FK89C56+HXBSy+RXPsTlvq8fphnpblXIbY6NetpN
cYZuaCtiCOG0Ua6jyb92FIlN20JDiTbp0tzQ/95miusHjD1Kfq0HUZRTrzx43Agp
qqGgtDk3nE6mJvxFtAD6+Ygd8zVUMGxP87dsYYlQS1d5HzURcXwKVcESgSoX6P3a
w8PIP/iJo3pX8zIdn07DRCylQeHDFJJ2O+/khIho7b4wL+fGxWUK/gzj8kHW+8mU
ceEnwDCAIcm3wUNgBy1dd5PkRWg0ZXthSE3W3Gsvz8GFQpRLpkv50NF0LzVE4TuH
12MdShodfJMAMl3vubbSRCX7hlm8ak2ltbIqd7rDHAnkC8D49aT5VZ67K53Mc8uN
iKHm32h0hUxMX33VQsMe1hGT2WaGjCu6Eo0RYtY0gJouMB6cHLUwv4P0NnfAF//h
dXlOnfnOfhBF3loUoCzevd25G/XsifvenmH68HBtANGA3N6Dqvzf0j6z7NluqjUj
0R9GlRD8y8VjfABOpDm+PFbKky9AgCDm2LECq8H2ipMIvIm9yBr1+S6XmtC+B/wv
hug3i5lHsWiLxsnmiMAeH0hHc1qiISAdqQY0nB3vgUZ04lpRHdwzOiacpN/4Ux69
jyhkLvYOfqaggYABfHRyAieiBTQ3+BjV/A3O16mZ5y3uWiPp+W8LMvkkNHa9aq/D
IZGubqmnhoflQjezpuIHFc1J4DNzX1bhC0oZSSomiTfX7XdfLkJU7Zt/wSTp4wd6
1vbh1Iu9VwK1yy5nIuUI9neczjwk0ls0X0nRKW3DHCsNy2qBTLmdpsNLkR15UVMM
nMhjcNNUEveCCK9xGjlF66Po2HRCBOQKUgRyP+q4zLU5Y8uF4hn9Z5YcABHNhTdB
3xVLKa6ECZLkwohFRP+por21UJd0mWDg4wsYBi6gHrpHNTTo6WgCYukEWwDyYoSq
vzA3b3oPappUOUoS7EAiZfOhdKk/rmqN8nhrLf+vRBw66rOUabk4y8GDP5OsF0dT
ooqMGndsxL7hLWNoP0x1B7JmGLBU0uOdaLcBFZIAjWdfAmV1nKo/+Y/+5L+snTG4
PUZHNXg6yJnt416Nk67yGTvEhQW+Vp9SC0XUf9pUV/5mF0LFlCwP8EyTrh++0B3o
S5DpdXq3J24aIcH1WQ6ZsALJokk7OiLrhkM0NMY13BOCP0eGXf+2XazvJB0/IexQ
x22DH3UfjgHB+XMQv69JfIKv57b90c7OlAcYD7Crfn76VTX4w3T7sOI819mbvI60
LWBzpiqwg3WNghTW4/U1Pphc1BilG5CBWtmSaJmEAkMd0DtHf38uW4JN0L/d+6gF
+X/rd0RtO1lqFul5gNbfecgZFsKW+D2PrYJLqdhbD2nIZVxtLF1fKeUb7EWXqzGB
nwni5HB8Nb/Vo8LmJWCrE0+OlHmPKCa6Ojyg1Z9UKMhBmFyltzqx7sPF9RY9GZvd
wJ2RJl1gKRcQhEEqdKCg1ojxLZxZFc6I6wAc2m4bcE+kkkPGG+3JmEphLsfjXfIy
B7D8qAM3qujy04B6R6DkUa/fdEd/X7lYnUDjlNgj6n/XBidrn39sAj0YN+ZpDQSR
8Q+TbZ3bYcKhB6vaWYbAuEY5prG/LdbF6t/KlKG8GSG4+fDDv9sRXYNm/EdfTFab
xuIDr9sYNPem+fuWeEyeev1L0oWILwOuuZ7yLTV7cAcakDHjpU6AJwLnAQwGu3fF
L28+kaU37/05kUE/RszUxQzewJa34lXpHqXDT+y3fObK0GHst5kd/Al80/oHSqI3
vJqsXhno3NhHM+PYueVKf2k4umZjsQ0AYu8xlwuZ4RvxoFmP2LvJ82bv6v0aZvBD
IF/7W+Ahzn8oRl+AXFqnFH6i+T6etZ8tJ7nOIgh0XRaevmFS9g0QAscSWXUH2p4a
QvhB1bjRc/H0gYYx/VHmm1ox5D14SV6417ZrOnBsaGD5sJZqptWsnu0uukc3C9Zn
LU8RVIPY2YENg8Gua1gEPtAZG0gZXf5OKcG6/0Uu7cck0tsln7LRmP3yKNNzDhSb
GHQXX/rZ/OEWMG2vx+ArFL9FnU8Cv6UxJSs0g9VpqGOJUBTKjHnnsJybclcMasJq
24lxi4OkJQIBtA8fkmjIezgD+JnLY3RtA7OGu7tQq7RJSw2qXaiIPGHWMM5QTlpQ
JsqJ5wC25uaEGN2qLP8UM5srzcUkisjfuUTK2/aR8bUyy4mvdYDFy3MOc+YGozJS
HZxgoW7D6/4eM3AO8tO7qW9rf23fspTxDkZTAPoTv0SEi1Hn2KE/rsbgn2Q+lX9N
u8pmx/YCcEVSvDbax/9z//hmGbMDx04wYN4gx9jCWiZt+Z0Mf2BaxI5IzqAhIWY5
SgCgVJnzb5G/lSqF9CtJuKJV6jNi40XNqF76oY9NT7RPvfreBnrBz95BPAkSlTjJ
AU5Y1L8aQC8wGWJwxx0SgduZpkHvlbXVbF9n38E9GVabXLWUlVbjCwcpokIJvanx
tvYGWoQYty5dy1HCiTWotrnMoGSdorc31FrRY4XLrPSNDhLlarlhXv4c9qUuTLrk
AicLuNk5HRHmo9HD6FlGuh5MQEHHoIy/tatQB0VaIXxfHyipi+O1vTuClo8+vu5/
7Cr6lQNS5rDMjYZWOWj0lMho7IuqUpYtpytR3AGGJn/LoDoeSqzeSDoQUiaoJtHZ
g/qDw4i1j4iDJHA0ivvpGVGyTvY8ELbOAdcPJFMzKKi6frEoRbYRavImBh+EHZm9
Vay2mRXH4gvapIP6ODYWDVGrvrVWlf0d79MNqxjMtoU/kJMr4MVFWFejItP4MgpN
ZaoIT/yvg99agpcNBw0nHejYyyqk+2CqJ6AuCWIT/H5TNWq8aaUmhITkblQN9I+z
9N1Dbz2Y/Ingxv9m8BgNRvLyyneno6lQxOyBx7/EBQB7CmfMSyqL0QlmM6VvB8oU
uZXcPnJFAP8EYZrCVuxnmngJXIHe+oUA0Pp7jVIWp0FrbDA3ClD8JVVcL4MYby/V
EzX6NHpnRaAVfuxL1PwrEST2kq+2GO9Wn8H+cKf05sufKf/eHnMx2KHxWcAOds78
wxjPcxFRgoFD+1KLPVgZzf/bOd+UqEt51VDRogBvCAmMJeydEX1Ezd0dryTcfpWb
NKlCpxfO3GFdKPbPr06a1IXUyL1Hx76GQmZ5bI9C+kpW67068ZGC0Gv3Fx6B5kq4
N4t7oELXoO/kGk2IEtq4tp6FKK/j5OGcGph9e17s1sqHSXGX+n3eIarzulSwDiB1
t93eCjNIXnSdj9WGraLtvhu0eyK0vHPRL/NqbFP/OLVfIAOa6IaAkbbv2AP4lCej
o2Lq86S79VbDfShdEgVWef+cNiactCwaZBpJ/0lUiVsl6rNY1EKuoA75qCV//eaP
GtdoON5PD8mdlXMLb9OnBoE0B1WhvwdmFuyynuiMWx379ob6Wdv2d9VutWI/Qp6P
SIvCZxbMVh/hUv178UqzJgSgJSinKXOytIDKhpr70dRXxYa3gzu6wFjLRl5doWs8
z+kSOZp40yizgVqwEEjyIzZzS/PjkDi3D+UbZnz2aRsK021f+eQJjIsbHw0weVma
Y6BVOXprw3eLfhRjzcJ12rwrZq2v+sogym37Rl2sj7MPQdMn8y/hfgjjVo92GVl5
bZD7tzM18OTSwArUIm4xlg+G8KUtnr4+qu2GMM3gkgbnO7dj2/zXdItPsoDZCa7Q
+P69q+SxsmVDr+M0BalDkx7nc1H9/6aYH5mLljiLg4fZgaWuBtocMi+jTvEhbU0E
LiqWw0ES8QgTmv+hQQsZBgpufcw1z2GPINxqt8RX7v7aNlFdNbqHmCnmkogovJP2
UMFWh6+UQ8XkAYExXRkdIrLiD5GedBjsnyZjIJsYfuebCe0LDl+67NOBrvli857Q
iGUHIOhFHbhOmFmtqK4ANzpEwo7f8QHZKUM0wc+NYuNAl/8qU+ajPjMLrzER1maA
tRHWuVUWDe67XoqeTi2i16Lne4YHFoIC3uHnSKKHZHYgfpHPCWVM7muEtI88ZDrR
7F+3WD57E7inYTcqkJzP5/RYxulm6fED0lukqMqq4l9f/4Qfsx/KgtP/F/ctC1OV
kt9mIxvYkA8TCX/cC1T+K/8eDU1Hyj5HRLVQvZQVVkoAwcnSaj9tWGN1vb7S8LOL
IdYHf2cx9q5mYBxZN36s200j0lvGSzP6FOIKuCTz5NeRrtxxFMO1q3yI/9qihz96
NRpNRjxVhGTyNz0tYCPJHB5k8sMhryAN9U9Dj9gTlpTlg8ZYnvJ9TN1pZGpsYLtw
X/ruKyRM6y5zj/34h5KpzN4WqAMVK40OoIaXigBb9BM92In1MTdugS2CFKR5gOxR
BTETDjHy0ecJj6rMdGqaZpSjnpDwqg/sn0eyFNEjNAgOus6IPEwT+ljBBtG2I6Dx
gkHzW/d1yMmDsLO1lu812ybiUiKnPwBcY40/fd9pP7ON8QbkYwZ6syvMyaL7O3Xg
+Yh6WziPy1UJuEj8PEsKrrAmMSZj0/5CkxnkVBDgzs58VCVhQ/tplTsrasx0bqH/
/kqbfxfCjw94J6+5ojOIF5OHCA3VxtP5f1MtK4Lxo6A+1OfVFjIlKtOB+V/XBtgv
gqddvl5eCjQaVvT8a0usYtxCkkkdO3f/Kawv+1kV1nRLLMtzMQYrb4Y9MCzPgU2D
94SznGrOaBsptYw2PwVmaiAxoSJUKcLPALl7WYeIzrCAqS295/bb6MoKPjn0xuWU
YLdZNwST4+9UfvdkLGmYU6jngjyLXd5eWWlsUveLJ6jir5Dzp6qTVtB0hvsx8nGh
WH1hwNW0zdLm3PTsqAMHXyb+moHuv4F0aBznMWosZmX6OfthNZ/zzu9E/AKvJP8b
h4f3aDpqeXl9xsz2zwf0e8xLVpDjaJapkZPyjYIrA41+H9dwEHSQXvR2pLyeMqvh
8WazBHOiFchVw6inVVidhXb8MHF74xJQ6vy5IwqCXrlXdALBIb3p/YvKMRUmZhuE
bFqrzbOV6N5dlAQD8OSfI61T2vRrX38rx6bvLtngT9q26Roi6OxRCiWddBPp2nWD
rGT5TqHDRaOKsh55lBajNqss9r8FxsYrnd2ru7C/kQJ3B8GTEsZzyrKfWUih7tZ7
iokTMre1+xn5wIfSHc4joQU7DPiIehxFDC5m+LR+h5UTjcU4dWiDZZGgKoQG2XGW
uRQbfmzhxX34fJqzhuuS7HN9BcBsVTVt1g9wyPqAaOz17uCtWBDDAC4yhtOjnEnC
XiAR733il25kQjKwBiDSmO4VLwkq9ygh1F6mFw5FTKBYIyveNf8IxNu+QDvofMUu
PC3KWyco4gbBjRUepJo0uR5p5/fL7LcFsjrquWpBv6m6Oz1PD1ichD3O5gkNFccj
MypagsQi/mEl+VryU09wo9/xkSRErje9lY7vG81mHntWY9UymOEqs++OuX7zPm5e
vIgOBjjyxbpfM4doYmV7HDA5Po5rQSpO4HQ7dOTuLA+kCojQoUHOd9h7v/Pr6xMB
wBsc7phmyo8r3CAzwOu/c3uDkkE96xidum88IoSZJ2dYNlIVoBryUf8Kin6EgqoZ
b/wPjnsQ7UUL+7dXd9RBiGlrJJrRL1mUdtQlkqsr2GIAqFKqgAbbTxDPzQi0xeFJ
H9uPb1bIMIcUC8UPtFUlgWMu2XKc7ahQ7RV5DJ8OoP3VXveKsBgdqi++UdZTb0ua
w2YqFMsTeyZWW4jp9DiGTEoqVOxU36pC7D6Ex5MLWanKZEHu7cHSlI4vNlMCiXbz
DGznP1E756IxvP+YM50YfwuJRLzD1e6owuobmPdx7M3rZsjUkqRCawZVKWJcmuu3
BhSBgzkue9uzcUBYomPKw7WnMI3/g2lsmIz1c47A1IiLp4KCAtUzEirm9an0+iUl
lhGemskQHZoXtOFkpNZn0nu0o28YVdIyJdTTlzvW8yXBh4yzC5a0HecEPgSiyajG
+1xqQTXVbcaIe6yw6xvqJu1umPo4qgogh+vZ4NcexqxM6mGCEoAUBO5tUQ5IqNgj
d8KeK1tErM1XlfX5C/bgQf+rPObQuQ7Mu0iCdoLFYaDwzcsXAk5Ja8Um0uKWuB0y
haM9/4nAlCIb+SNOUiWDIYRZSCHgpZoG29CYMTqBPVjaLKbvhfFZzWdcL2GhTaOw
I45IOTz0osedFkq+AOfdLF4G0hf+FQHvm6ZOpuODBweUGzxQJWoNWHEFUEKD/1B3
lvBm+srau1DUSNZa+jVUU8Wc1ETx4shRbFMa/R56wGgwmrnxiIpmOFeMvdJj20/A
U+qvaXOH/BDpMwJrAV6vyflXdAA+Z7Z3VDl/av4/4z2JwHN1+/Lpl2ah+iIVZ2hE
V+cLwcqH4rkc3PxHFCYpf1RznezlpwgheVbFzgmAiOfhRKtVoIIh9Ixmcl3ijmT/
LoXbnrHhoW/cEGnU5xJ/CT+F1b1KLbyXd8p1U8dMr1ACQCIyRFrJsNjXYWVdEy9c
kiHrL+UECd8q8dYpnJuF3xs8uVGx2XG/bnSPSHriLAN4lh+46DaLTF0tB+z5bmkK
Gs+OQT7+oWlTkU+f3Jv99qXfhEI00ws1/UHotqTLlEael4py33vs6PrxQYX5tb9l
meO+mvBJ97t7xboeE6TpZZrDJUKy/rQdkEa6+BtkVh3CfSpmt0ynmiVhrd+7Ro5l
O9rkt/PtPmAeYfa4MEdEMukasi7lecr/9xl3HiZXYkjQF/QRLvZDB6wWBGApRLiL
ZMwSMDMeysHnsJAKTZTojmTcSeRe8psstVEN9ZAh7/IiSkwoJCGbEbl7HoJtdC6Z
CLuvegfSU1MkNqM4k/t0Yg7gSUR7Uz25678aQAzlVaHyvW7KYl/g3+wSYTl17/5D
scAW7FKWSMdPp2s2jaQc8+YWeYx6B6FQkAd8pn75iMA66Vay13i88X7VulN3EQN0
ta6VeeyWFTKl7ncK6eIW38CcJYgBvCvC/hZe1yMtSd/VW5nr88W4kCIGdshCc+tB
tPzONvCdToSDV6xonLpOCzYzJg4FZs/2KmbRm0BhZ6z7hwUqfoFtE2y4wijOy6LH
lba9GonE2KohmRygp0m/jrwT9Its2PuW9ENwoeTtTwoUWeHYrbz/IVLSPeBF7apB
IQSYPkViBNdAfDuzcsd9vaIWup+0q+1+GkYhltXXKs0lJAgvoPCfOx50pmXlB2bF
64JGvjYy1EFj5/hjPc5HRCHN/dNItVMTNH4nLDpXRDQEFc5Ee6K3ob4SFkvNcX+I
orw4ppsfrgZEbUrLBe2hitV6KhFRiClBCYjkpzlCkzNtuk2ZV+hOien75hTNDUNa
2HlHLZdcYd5BlT9d0n6oyurDBzYhS7lo0IWnVqsNEnrqkyugndNAhhXg4ms/QuSA
ovj3Bpjpqt70LwDyVofNGOjyJgccGMsyTqz6Fsi5bzSucjTJfUgIxOQVvQto6cqw
WrjngjT6EJwwm2kISVdhHz5qgH1oPlNAr3R6O19RqNeN4Wku8+m00VJdBVS+gtRf
pxP8gz+PCcoPaHrp7P7ImX6kwwiizFBqs1Ra6ckMTTKVE8FLWP2Uh48nRypVikdP
gTjgpP1buJmz0Ik4vLS15czSsGZIQmxONebsvj8cni0+TyurTroCzcdFBF8Cf9xJ
1ACL5vQSekC64Kbpac88gg9b83QRKfgIkctnqA/FvbxHd/6F5zmPHi9rbVuJth37
Ana/s6PgusoVSWXEMGPdSTrxYksFh2gW7udA6B9DXnSUvCMskUqnLFUah6TEJGPs
Kx9JOiBRVLDaIqEDqkqwh0AD5xDQiXulKlVcKIS1UXLc3yTQg4IlF6Faz/Ft0Wk5
+Av7utz3sjoTo/cP8ZR7q220E3oOTLmbD+m9FRQe7g5rm1xeSlJwLJu8aSX3QSJt
J72ciiv9bbS9aXT+93NXzJwdUwoTudPEykuXhqwblkqjHnm6J30UOy5woICK3Q0D
u252m4gdsS1qekYkw2VgSd63ej94QbO8KLkQLk0euLuAB2uXQV/oyZyQOw35ccVB
tIo6bwQIc8PkWKV+MsA+dL3vlCzO7sz8hfvVwszFKs0SCLaYXSg5JfNGs884hROT
i4DRIcmo7p3udT8nhmLazEP9q95hqbq7gOCNuJk68uThMGOo2aA3GPcZVikZR0oM
+/qmxyAh+AhMuu8pLU9p4FvD0g1q/BwhmPBIcC/FD0X3AkgJbrbY92400uLYCMW3
aWOGeUcWzxksmYBqCEpqve8EAbPiEwVSC8NipekUoHTHMVj30EjTh6Hg9Mv8qmpF
PkigBkkLkuhP8XYABwnZqkomCJmyEyEUdBn/mWVJlO+6H3qNTwORJo8YJCvSA1Ak
2v6xFWwPvMWXNng6rhNSLIGri3sJAAqVVVqBMJS17sdmO9HKgb5yQfxQjBerwzUD
ZDRZ+vRNtAdMXXUypoLvF7tlGCVNPYct4J0wryapSltPwwuYUfAtwlEPIRmHQOX1
i7Dzl5eGMHlgZU7Ntl8Mfqq73L4QxnGTc7DDfPgefOYcq4zyc5bwqPdk+LeXjta6
q/ISf5o+rILRx70FpAq1FLjSS79Z9PmFhiZbKHCot0uKKNwkwMA1Vm1KZPwrpX+N
rOfKIomFhIjpbqxyTJm69DPaIpfPSR+rLFeOCOZtl95hY/QaeCeT66jCh4M5lMLk
KH1v0CedrLL9VnLIOpV7A3hEIfOSWUnuavuBmZZ2g2sGnZr4+ZEpy2tut254vSpi
LxheOoSCNjDv/ggcEJLfpYJrahE0yEZkS+IB9oQnsXR6vF5sm8B1+rJFM/7Wgtr4
k4gIbcum3ZuD+RmXXQIRTg1CwwIdQUErhob/oCh368ebYBMnkBmVb7Cb6c6WfV0z
areoABHsLfx5COM0jn5oRB4RMgNE6URFefRm+PmVnk49vXNEE0UBOICpGV6ZH+Cq
46T74ep4F9iPaKGNi3juNaWsiwEnCPAKpKsfLo29YbUF8Jkckw941Q/ITZ4/aytz
hTexa7A0/DnoNq4FdHIgc6K6syWD/8orqQtQEcjOqS6z5Ylt8SYTqJq/q52/HpSj
DbqJ3TuCAoxNAs15kvY0nVRmHyyaj3barxIlLSQbRfSLhtV3OHdB44GaxGOIQ0Jk
OYCkhdu84uunEPfLeHPYI5sL/JoeKQvCwhVWZDpsGehItuORKv1Pbq0g34mdwk7O
NVqjdQ8aV5+qG1VVrNF57M+N+4Odb+GpVbyzt4q6ZLQ65iRuHq7AmpHpcn61xCYD
0TiPwJ2gT6HQzQLLviieMh4eUcsyCK6uUNzSZbnI6SXqzg3Z5sXfehV3SS5IEJ65
iucZwwqJBY7vX8HmvY90lHPOyXpBqLc2daEu9pcXlMvmvDu2GwZ4QndpnEu+JbPC
wCJDS5eufZcOcjNZ7QpRE7DYH56bDDqVfbYjgUToOqru+uKGT9YMj9yX7YbR8M9i
oN8j5biGqD6bkNnLws561yvdaAuWze1TI9xTTr+G6iXfoIXmacaAbpgy33rdevBp
siPizNFtIHbDNQ10JdFqmluK2BC5gc/SbLxbrfKiSvPy+DKRyWnaPwOQLB8Yq79V
tvRa4fXuujedkHYPghrbpNmBaJx8/n+Gyu+U6xYZE1gfosHgllXMl3Y8BFfl/0+1
2ZCkYCYKNM8Z7Tpx+YdDF/1skBm5B+CTfMuVvdggPsUeMr2LGnGdqHMyikMUNuvV
IphZUh3H1ZX76Gj3F7Tn3cVOWzy11aafbO4qdQkDB/V7qX+JEGCcoXMOm1q4OpcZ
LE0kTmMT7iPZrHTAiltIiO+yIC5BKCcaJMHlIZs+LUfgVRFOqNv3zYbuY9Rx/p6B
bziigYnZhe0SZvCb51ZKjiP1037F5kyC5IiSyDFKOHvdeCSF+jSgxB8CTa0h8NW5
JMh2bqxXofjpfNheCEqq3JhJrM2cgrbqlPmEAga8UCWY7nImQEQOeZlLm3foFD+s
32RnNNb/78r+GLnRRBxxP+x29nc2m+UDpWmTq6pNJ2FCwqpb6P2Y9URvAw6b/h0e
3WQbR51BCdDOLpWRb+vr+7fGmvEPCPdgv3YyAcHkTRNe2jhMAqmMWJar32PI6jC5
NbI9vo8RFQWy3lNechKnGoRsJyF8U9jHIjGF9hRG/6SazZsuX5zqa881hOX4vQ38
Y2V5wqfjlA8LsaGeotUfYVbtxxLyFl5XAWJ3jrNjv4vqR6xwzrnuAPERJ3GMkZt5
yms5vN57dDtW8xDxfNOuH+CwadSfS3zOVc5MQeEAAY/8Efw6/B7pezboYp/V76T1
Yp/ur+XgTj/PSP3MCvjLAoRq2nkXxEsa4pgQcglBJXrfuPmPtm/b+2jyPftAfDxJ
7T4kUKbMroAJXNNc06F3WNiIM2/j+Y1roNWFlS2IVG2bX0vKNjyD43VL9TpvEAgF
PsFtNsgDqEu8T2THYy+yNOhDVJxUr1iK9ZjQhnICieZdnsOjPPh9sjYRu2xVY+Hs
WEC2DmmNy4zWGTq2QiByzkkHwYGTmgPSvCnSfgwD8t4XWt6T5z15u363UsDGSuUG
886DS+Mm7m3nJD8T9zJC4uNd1tefjlOnoWu2y3FDWeD3Yv4TxheYdPgAlI2ZRuTo
L6eWDc2DBOzE27USBjuftnSMQcWQehNsk2o9JKU+iEkzUsjdL/svtnF6VUWyb3Ft
9Qayk+NR1N1GbsLAe1sikKk7O32Ss6m728d5L0fujAFWJWRkgw24b1Ai9nnxRaBz
YPNGnqZ0O6y96V6h+LkT669r38abYTEh7ShIyb+5II+h8cwag/CO//g1w9LSFjxp
6DNnmbP+1H0ngKWQCeNLPAbVxCZVU2l24KH8qxALrw/XD0nJaB97MPwZpLbe2Lv9
bT5dbMGYlAvyrhv+PQ9Cpz1t21d2+NUgzU1W7mn8PVqQSKvrEE3vCOQzQ8idHYbG
U5k418hAKL4EsElnyJIHACYiwE6clD5lmtYRm5ZGf5gCRpOfU61Fd2T0HFfN1ub4
tHXIl5zXxfgmoZe8fC0NiT/NH9lEsTFNODY41tj1v9uzTAMaJjpIFU69pdBoSAVs
d/5cI1WaN1MBRZcN8Fpbs/5ayTArkj1i22zZigGEzWF6u6KDwh7bzgZthxLNlHuh
1YsMftFS/8gSpfODWt4lpTpjQFS0sBopW7kvWz0Hu1WoKm8JqfBkM/rtyRsRNTiE
NBUiyYVolwpQlUlnbhuqc1LN0i/nkX9gs0iv3iMQ/0mn6NriIYYJ7QYR6rSl+r9e
9w7qvWreIhaf5leAzBxAxIs2flSi2JTQfeOUUrnBvkPr6cE19E4U8AcWxsY3kjaR
VWqFnxxV+MP0W3a24jaVlyIcEr+Jt75TUEYeIptzafYBgq5gUNSx3KgSbAlpwvnY
YzJ9MQUC4xBpKycCZTYiJ/J6mHFHlAYFiq7HEAQIkyEjFBi4PlaRCQcKNFag5pIN
85XM36DktYRLjgYNW7dIXtFHR8rQIxC1pxbKmZ5d6ToYGqBCuoA4weypr9w530FT
ksm1RGbOQUGdP1xcGPsI9jMhy+BvIOgYYlehTwzcMGKJg/j2rziGGkR9X2/9Pe3+
2ZBcTsWGkf0d4p1VZ//4qcw0VTNXnIf6+SpMGfrUQ+dOAQqcL8yMLRYOPeqpaVa/
4KVHqgHBbALzcy7Ov4L9BU8OOfdkor7fR/w0h5xcG/8gTsrxfbUa0tTohXfk6HMn
T5yGcp5NBpe5PAo8J2GZ+ZkucjlkBhirHjIMr6+GKLH7ATuMm5ZidjdRc7ofxJkP
q+FFdaf4dlkWBMGvTWiG6LQOAIysG/47V6f05oX57xBUhZ+OBBI+l40oumygVbSN
FA3wMc5BU0CJQXC0axplcixeXgLiViQqC6eXZynOEJJomfypxM1N/BV6GqE4Rchq
gFucw7GtY6Bb159PQJ+i/ShoP1a4pjtPklMuh+c1PqDCh3LB/Xlm0LyVL1GcKGth
/YzQ6iFA0hCdOZEbI5MEYowcZjz6Eb5oQsZ/ZSUwudxxvaKzDwAenbh2yB4Fs8cR
oMGSs8loDA0qbiM/X92T1MWFYZpqaF0i6yMD3QSbPbuFFFqlcd7yt8P/ZJqmFJR2
noUFqfYFawfpu0B4+i1d1oAJq8rcBy4L5t/aRv8Suxr+vpXS939dJZXAPyRUscbr
3SoUBno7Nw6vj4inR7r0MoGv5Txw0sWemS4z826tjMzDKY/I7Tu+9nnN327kamlH
DUrr9RQbuyRc90OvMK8H3MyBUosYpRj//Lcv/X7M9Kxwxf7zjSVOZV8jp0vWaEev
HCiJ3+GQ8LYDuJSBPcKcxEBmFG8ed1tWMemM65EsGOUcSKccV8Iner6qG2SmRnPN
PJzcjeqzzSxbzeDbehMzzoc2p2lNZ7ReFmT2YOSC1g7CHI8g49/7eGf6V9EOb3Z+
WoaJ7wmauAfGNuwQ+yC2hD2dzn/C5+CyANdtnLHA0E5YKlWT2st0vzCIGNYo7D3H
lpNImgcLt8ZlzGin2ciCdUVEnBQkQQs3afdLlwRbfFQ1UQF8jOk0IWrs46509yJ7
8T1KiSESTUQajsc6jBuO/urHkFm6Q5LcUhG5EwNR/3BVenxuojOtIJawf5hmQV1W
HEwS/kPAuW1OJuhJ0TSdfP9tlv2qRE7U3b898RN/3mByz+KjWKl/8tcszYp+xhi4
b69detQa4rVVimpoRlp72NC5upninpxbeF1bIrOAePmmaW89BRmxgTE2zfT+t/SG
ebgOhbKat0nGMQCyhGQygAxDlKpHb/7diWRFihufJs3HUc59OkvxT9ZyUqyPnq5k
RXxdiJ/xH8qAzi3Xa8G3Ohwy1lTBYsPShk0yDqpmI7J2Z20vXA+cCKzRtdasszDi
HhX9PuU0W6mc+2Robi5EpLsGN+xDShchr0m5wPHY4Sur6KXMdHGBw5AHVwV0GrCq
uoyjV0rRsnK2yIKV3rU+0mT/hhch0ia3fzrgxlZVzliVz1VgsWRhu2rkFarVDlJx
L85caZCcmxyvPgiNjf+C8FkkfnKQhHGIh8QorGlbA4GTMY3w55rbzObeERt4YDbf
9isW0aUdLWdWfUaE7q2geINiWiWjeasV6OoXcZOKXeEjPBJVb6qfutxz1lhPO5kt
H0ZlEwYlSCU/9q/OepudPf8EKtRIIgJNflmnf6rY7tJRqedzt+bGax13ucwx6rqk
VB7u3BtfcONr5RGxv/Y5j2cx20j2dB+Z/whAAv2WkT4dK8krzOP9ZQgNXKeRCuIf
n9TIAXv3XpQT7KqsFCromyLGy/xtN99UQlpKMEF9BvwOL1QyPSqgyVUm2wbJCGHh
HkRKjBQ14d3DRx5gSlaKuiZGpsEIEVQX6zJR9KQVWHrEiqNvJz7MSgmTqmooS3QU
fIZNm/Xzp9CEGWZXZArHcfT7hpZ3CYvHIgvND0sF78tU2upK3O6odhSr3GIO4ius
Fthxna2DbCTfunyq9R8e8QBAwxkxFVD+vZmtIipULSQBZdaq6iF71M3swszvnMhL
WovALpKMbCf42PH0shQdKLhPi85t2Yz4odtxGf4LlGOir1N58N2/5UTdLPLiKf2G
bfJNK2pNSn9jzfPPjx+mkuvuT7AIEY4JHy3UB/ova7537e46uoQYM7eXSWwUrtqC
ZS3G/s24NdZEZkBceXcj7qM1xebGXuBQVYiuO6JLdxeK+VJBnEVZA15MnxUSh2M9
2ziaf1N+S73IbliWF8rJQzHgFMlnPlSSlhasRfswBQEdh3+1BJn6+s/e5Z2MO03+
5aj54y5FaJAG1GdsanAEMynBi5xKl44soxCykzbgo77DQiMbW7OUCRH7GG/+rFmQ
ccuLxwnalfSFyTC5neH2A431rbvCeW9FqOQEBjyXvqVRbwZEl/wDlo//ewZZbvkn
jpZOau46o1bNSr/fFLBORMCnJaYSpEokQQX/Ahr5Jq6bIKORfiy3UGB+Vl+kVzqT
Twcd4pY4xUi45v76rkS44FeaqEDHNL6T3+zzTMCLwaG5kabsMV6vvCG6sKw3HRjl
WGvrS8XVZlDYLAmNnDUniKVnnmLyiuNOx6Ya5UclMSlzFlLJ4ciz+FWgoyOYqhjp
0EYvQyEHYCWFKQoZYEGTkChhxrffD9kE5GiBapHnZRkPxU7AP4/5XXmpE3+M3AUS
9kkN7vAZORwBk3ANU5Kw52K7NtqGjNooxiMqRYQAI02Kdem5N+4S+9EAd9saCzeA
cEM8zPddSZ3MbDZyfVKggzNUO1HusT60E1fMppm0kTRdPT0Kzd+MwDTrLcan1gBh
BNoljD9NKFUzl276vhbaBtAw8WjoOVyJm98PiB9PYEbxRISX0QvGYIX2zwUWvY/L
i+7auEbTDHaIUB3U1U//tdWIsP/jLuJcEpuV3bVY38cwMwxXFRum4whsHjeW7s0M
Emy7Bu/x2BeWuOC9tQMwkgPh8aJeOD57dfBMYnBPRcN18bEMkyhP4Q1pTKQveMy6
gkFiS+5nI1OVuZ4DGqFYLAOMnwzXPZG2tcQ7gF6TG7hkh6pmSqAaRbmov8e96ZSW
z3vjKj7ZjvtSBl8uHQf/j+ZYqaCfO7rLowLMkSHF3bRFbNxy9vsPU2p8gKAlZYpu
sqmLJjB3HeGwoS+KJcP/7T9uG6Auzr7qoNyZ18xSdPsUn1Ma9WjUhX5/McAks5+2
EmQ2XkIoKUtTGQ3IVp7D+KyQ0Fx1uCGDVoENAefCBtBOcz/b6N7LtV2XDtI+fl6K
qGH3OkZcF4It+Dr5LydhgXbw30PiiKPvDVj9+3sc+0mS+npk4vydkCtQXCaqiZH5
6DX9QrO6jdc2Qo/4coy6YVV5HcXlg67Cb9LGPZLq5jTo5zstpY3a3I1aPI6Lki6c
cNIku5AT8G3ml9lzZHo2kY0OytK75HqmiNXaVRm7Ymb0EHVOtmoEb+eKtgb8ZcO2
1EtKQxZKi3pvq0EJrodvgBI7+ixfBNxihu9IrVLs8RVPhW+GvWPp0rrAnRshYl7t
KZZYkHqG8jUxqCTlzHv1KdmKGLtBrqAEzsaTZOdwzN+N+XYizBpQ7TIj0zSPBl16
xZlIF0jiVj4mQU1MRRXdbI2Uc441zvMvOBGCzwjM3GQLQzKIhMJ4Yea7BaatIgoC
7v+8XSypHC9P+ClQOJ/E1D0iZApjdtkeWT5cYBjew9le/ymZoFkU4DI7rfrB87d5
+6/0sTQjfhm7iTrhyZkr35ZMNZX2kiD9cMwake/+ykaa52Eutr+uq+Gw3jwIwk2y
S/DyZvka3jzvC45woEH3RIFvpKzxwWw368/gJhWrZ/tdBcgQlxReia5R4KsLpcLm
5q4mtT+sg550Wi9meCIhWOU8f88qB4Cv1ejpHr/7QmrQuYnFFGUp6pGIHG/OIsHN
JidDsKVz+zzXnT9j/2z64gPLoYWjLgTFMRN5OORGKCgaMgeAgG+9LQjgrxndIzqH
4eNlPF6rjbKFlsqyoQJqELPDvpAOMYJYcxvd9CHbURk+13+XsCkVkmprXrUZYIFq
8mo0TpKXDKRYxuEoTGLZborcm5yr3IVWSJlLMsLWRd7anjD6xliktZJlTSMGGtLe
Om96vvTmEqRQ4gBDoK/dvLMYEzZ0jZ9lKTbPJ+qT0WdLYUvUjtB8s6VXztkGXi1V
sB4uwXWGh4amfeo1nIa8yAF8gC00LEebDIbZjDMqMYR7RT2yxb1FUzBDgdRLgemV
jSBph/yNcqvqYdKLnXt4farnzmzvwIBhnywBMgv2VuXcHDzThFP7nfWCjUWymHk7
uG6W3Ni/TTgp4NhAUhwHWDsmR6kxLsQzuP92qWpn2XvoJn9wygr+Oth/IMn66sjB
vIgGvmCZL6T7Z4Gih1A/FtT363Qav9gXBCF9oPSAbby/xBcJ264bk676Cn343fAY
bM8Zo/VjbRH5VAE9e4Nu0ddv3U0ErQp8ZDSlYmXNatBOz5xrIv3N2iuvv8zsxEb7
U85YZ7qby8YEqXC0LsSnrvxt4I+pv2VoOj+MJdu7qbPBp1LWMJ+fOjkOLWevKoit
FG0yKp623NRnTV9mGiiU1tBlKHWE8EU0JyjoDqpa8lrTfp2F+ZuXpx9YKTrcTdhY
pFzU5k0qjlgCw8gr/tQlhtLA8Etx5vEPcoLo33CmRdZmvMhpF8/Huvjyt1oKoywO
exHLLkLhhBZj/qUP7ko+/M0RMmgQIw9MMbiATTH/ZCUkmPZFq9Ku7Y/iXqAE55Ui
diLAGLwZbLYCqBaxzRt9sM7CKAoTADiQyPjlZVY3BxD0A3vC8ettuF4wTfcsQ2CW
LxSdX8QsUqQvyd3cCYyTxjfAGKKQha3XtCr3KpOHFarm7C/5t820fjvumgRMmnPs
Yvl/44VFH/YIQzvBC2iJEGLO+yc1Hm98qpoKpnHAUYfDYL0b58Hzbpyilq59xCkY
3mDEp0MjpQAEBdvAnLulKpbchyvGEpBkLzmHPmouAos0FJgtgnvFz1D/UYsEDGeB
8fVfZieBnAVhFy3M6lJlJ9Ysb72k4JPCY7yEXc/IGQyWgW8k0m57TAflU02Viz2J
eeo281eM8hR8QYgNwIoDIG0EmTQbuxQ7ArqjLi92LAJthC4/yt96KPlHyPo2Vofl
5qFGtckdBBJfCSJifjAN8Z23GfX0mJjqAGHfDkR7JLsOe5nFRhMrPof5j6qJ5z6f
Gy7MRiDQtywLcYUoCDEU/IU58LLMnZTfPPZfA7AXfqMWEwW142hJd8NVPonBECYN
ATl1rmpdZxztLQtU4foeth8usipC5PJ+cNXwNaQCgIlAXxLYIVS15cVxZhKWHeF0
/4ESFdnQey6ewL8/JbpNGFPDNp5C54D2mFXDFZRyvKbGJMK4buzGyjlWQ+OpH2hb
RKPUuu7B1mTtxJAITmNwOOWbWP+ptAjDrQq+sXaWye18/0802cqIy50YjDOA8StX
F/lfUG2CM/Wf7AcC+7MB6/lRrPsYwzTm+bbclUN4/8x5fGG84bhzgMohepW1LDhK
ry/ajNAoFhGF+Xo77fNypwZesgNpkOGnjiO2o+V0mp+b0kNY0bLXQJ7Jf74q+Kd/
WuMFKZEgYyUHcXV09bmzpS9cRqbTjSGLtx3SmxsUGESSNrEDzFNAJzwsjWsg8vVV
KRvh+f1FzrMdnVqADm9Yc3lpcqJHBAVBqwMEDGxHlUwsrXLLi7Ae1W82hLJp2noy
xhIegsbfzSqn62gFsXC5BhN0OIrXDaCavEZzPg40B4R05PFnfGhUZEdJZO8EEHQ2
6GCPSNDic+MGSvK/1b8eSVic4nrSbdWXOfJAfFvITvBPRmHKdCpUheSLK7XRgqiD
F3c9xaUb5q9BusNrAhlXWPimycTbT3jZqABJ0kwJrwP0tXxvTWUfj1KydbqQ7o8Y
mc7WsPuj/HVtlBfOrEMcgLom1la57b/mR4jmg75MxqoDt6O433m0qypahdAqZCOk
gHLnqPuZW958gIEgiQXi7vnibnxhS/4JIXflifISpshGETyYNqWJlB0U+j8mlYK6
OWrALvdXQcnTAFc6iZ8yiuRymCp5LX5jOun67D0JVT19p0OQWM5MmSBIWZRcU/Pl
ibZjt7Gx947kLVPb6GlyfiFyUhUlPMWZGufwoLtrIVK41eATP9PiMzgT3OAHgny4
HbPhjfGyIae7tFJgL68eQRfyGST5dg6NjRjfRQ1jpb1P/o87BdrJQVIl3MS1uZwX
Fma3JLXwUaGqEFWTlnZASRzHnxgAWj9TWNp57gFUSfIKFYRKI/U02AhCLvkY4XFq
Fbo5Jy0CMQbvytpvsvaEhuFrYXpEacn8GASWXrjjP98nkrJxKZ+ShJmA+ofigtKg
Cz/DLc47FdFRe2U+LoiuOrgTaAGaCRmWn3vaCRi3gcPejoqQLeirBBtyQdRkeHb/
5HxnJr2EavmwzTfVbNtUEvKrOBn50yeaS7eEdVamJyUrKaKm6F1kPH7ZLUmPutUP
slSc4bHThf9NF2Eb6Dp0JyiUoGl2dQWJNd/FPRg+r2rfcz+VuLqf/EV/uZJ9XiyF
hqq4gfu6mq66pd4iKik3DyTDlPpXKK1ZsEcQtU1s7jZUmbLM4+ZAxncvI0lhjYyq
OhHX/esJfFJVhO3UE7a5AhRlufWUJyq2SNsglNSd1r6cZf+RiahkdgURAhF8pIYp
ZFhWnptrUKUTVu2diggDWicRBXXaWoJaPiaix0vZEJ2J9CKiZirfpzHz2ZBU5seE
yHMzkrQbcVKYUAPGygoSGE77/hxKQabylu2c7p0ykqPW0mKeZtbmrzLwXDGXtMYR
/YXXwkJKDrFbOFfCHJfJaLr7XGumCk0j/83HP9dfFCIgWchWsTmntPb6bObFWPgj
6KDsUjIOVqx0gXto+NMylWBApzCVR2Zig46ZGqi3MrGKRyQNKCBZdcdS6QXgmO0K
OPdS5Vyet2jQ+UptqIOrK69HvVCIvRSrF+GBxaVg+HZRwPOaLcS/vad5O4vfb/Wl
3JkDAdYnOnL79WcEe4NCyKbDaN1IHKp0erw0gnIErX+C+UamE0CfCbV5a1b6y9QO
5srRynxBJrHLxi5XW9JQf7xTul9te5Ah2uBCO9FSIDq5n82DgH8rK1tWRGHMlg42
dliQeAq2K9d5js0ex7C6uAmI5+mGSsZzpngH0m8fywFCKAaLxxt3pzrfNIptzjZ9
ltpHczC5mVuXuWpdx4WI0mqsuronFEeY8xs+fKCDtXmyDuUaNO2ppAqaGIm4lmG0
iHSNZ6WGBh1DYxae40CWMALUWGcLfzWFOJj22V0iF14WNHTe2CkEsg0wcqG38zM/
EIL3Oo8BH9+yQdr0t2VnL7BexnzlfCHOO4ql538wAnGCoiRFL0aWQwKTPAbfGUeb
NDUnLVtRXLkRZa02QtYHmRItiT3pBQdR66ulnL+C7KNZZGNLjWhJ+RgHV0J1GKi6
DQjUnYudrG2wKs1eEBzmOks8vKRpw+Hafn8DMxAuhi2kcqE9GAAVPZiheoYIV8Y0
PNTWsk8F1eJ5UpABL3d4GuQRHnbADAwHgBDj0wVX/S6RwfrNV3IgBWe1Qv1nULxK
PPOodGw426yW5zxbCIp3ZzSSoliyd99OsKv20KXP1HXzikPdVCRldbEzvAiqvcYi
RTBNYoUrJNKKfbbLSjMni79ADHTzMMI/ElzuYwgjuoaO9HfpkKe3Mk7iSH41CdDg
kt3a8IDYwZyY/tzIUfZIBbwnT3q9p3oFMpAf/ciwhrZEbintkC5UPI0ACu2GDbi7
MxOL804+qRBWl0IcMtzT1tHzl0TmnHplTCRi2YvmR0lkAKBxJpUjmXpYlede2lzk
wniWVxNfQ0Y3fuYlX5F9brbdMvos832WVIdSlmXJtkAMsYzAP3UkECnDXOhTsPLB
YiGgBwlhJwIfNzrL7lI5g/kpMVjQwHvx1MrkF0RYePlptF6/EYdjnxpTRgakUMtl
B4JDiJgi+HzBcLu9TmPijLbAFUMeVRI5zs0AS+NAaOHRTExdazrrtgig18M2s8qr
a2tM1mtBHZxi78ntiX4URK/QVRKkrlBdK6RFNoXLDOigLaf8E5nDrhbzPJAEho/W
xGo8nC3kZU4gLgXD65TBFmNid2wyQlw+4aaS/9WtyiPBOs78oz3Jc9iwd0j2w6gU
UKAxviVNvpqoWB6g88uTVWlLp1BgwR6KlCUrUgzQp1ZJAXDcIXundMtGltpNH+8h
qEYJPsky/3fLX9q8owlg6zXLCHZVKKwaKR2uvNYC+xAYm7+64bj7SB+YeOGAvlJd
r2adwaTtEAvyev/HZSZXfddGMG5KM4AmQra5TD4Qo0tfTBwdIiQHXpX05+Y1W/R4
FP7OlHqEHfoW2FUIkv4iR8NeXaqpL42pjMbEtrwrIpAbUyYWOhfedtzfXQUSMXiz
nbM49M3SZW0yASif5cTQL+uCg738DXl0RSSg/cj2RmDuYmxIRgW04W6Rx2kvZJSD
3LqbWdxxAEKq4GujMfOODEPjIwl4XE3TMxhsu2wcAaeUxHZBq6DfxX278M+wFX0p
SI83tGvisIuFBwNwn1bAoHlIA1WrjNm3jFFfM2caBB2WJ3394cMcoQ5Zbp8hVwzN
SX1Po+ma8mTRbut3wlx8WAtYch4+XRymLGQ4Z6Vb3oUjbJHz1XF+TrUAHkGigs5z
aASJzipGYRbqsdyh2H5x4Au4j4TI9Lb7ymklKHJ0kTmoDaINUHL+Zf5VoI2MGNUE
YkKVniotnhLOIjUvF5LwLoCQo6UUu5Zg8njHicMqe/6hM840W/5EuvhYpG703tjC
qu0is1FWrgeeiuaafHa17XspRw09CdTT85aTu/HEgDjj9lv5r6LGgXD9ZAx9ArrH
WBZhUwSsytOYkg8LOhI/gedM57pMRYobLKWbZrh1TofRropMbHwTk070fMk9ancj
Eoy9NTZJYO0KruyuV6bJlnbuobPKos3lanumAnESlkIekjfvxQsjGblAYKIBKu6b
t6pgPa/Qs1oXzc1bpPfMvQs2zdbCBWz52IgTNhdVFze9eMTOl4D1DlUcolRTIZCJ
0fjX7KK4CjUQqBwWGNx94kHQgeKYbqUwjqcxPwg3y/4OPI2pbBFTtdPjivEaP1Wl
qP2j4JS1tihI1CMXFR6uwIl8nPAQatLLTV2MHBf/xRnbAXL1LdXck3p5jIksGeiU
sXWfKfzq6R2RGtmee+Tgocv3cUc3VnHFGwEh7xnNCbn32s+9y8SSVJYtVrCMvanx
icp/MRi27iPdLv4BzdrfW8+roQKEDWJbq6WeFF1siupqi9PwGvqzVz5PegQe+A6B
Mb5NmM17sgpuL28OMX2C+zpMePTM/CWPKwiiK/fzRPf9QNmPbRnpgU8iAijHSkBh
waMaF5hDlhL9AgaXwclY1wtQeVHxPcc6CY0rWNH2bHXi16zmttA/FXTU2crideKv
dEzN7kH5QGtfC/Qt7ZKXm5A/S5Moi6xoAWoI/zBDyS0QO5/a2xqgtl6E4UaGVZ7N
6WhCe5mWQrQW9F0Z5SeQrAZSZh15YNStsoMa6ClOgQDg4wxc4zQCUrP4ot6HMfZP
a2VjuTLBFgdCk3hx6MEFjgCJ4J2q3wSbgnPfZgelMrz6diqf+d8xPwFsz3and1Hh
1Wh6oOiXl0BckqV4uZ7phfGZlUtMa7pJUzXvFLc6xeT3fTmzQH4s6P2kZT8Zp9tr
FNx1CGqzlWQ+ZhOX1ZVUI8CWtFLNTtCJ9cKe2Zs1Mr7zce8C0t3GtNfk46JIjbCV
hrrlytu81D/2MLdI/4mlwxheyZNGvMD27clDWPYxqt4UCAtGTF6IqBXPlXwwkBAh
kxN2XjvyeofKDQiSmC2eFtCYjZAR+AgCFUgt9oX1JSCUxpP5vui/nDB6WlcXnYqS
hAUM/QUjM4VJWBQHJuXeZii9mn/KpTCNBjOBFJf9ieJzwYtyObClm5u5hzeysrOt
wsv1V8Z74E/mm64BYIrTWvEggmF2JYUNRB0GwXx868rS+0jrVs8/4J2q39SevFkD
QfgyFMth2L8PDI6iSXVrhpgdcImFWlKlenbri3fqYEAgUMoaCFMzdiJdjHmmfpzO
vJdpxpfshnqzq1a3S1hY9sF2nd0RB9rAlQq78dkxg9x9kkQSonSonC4Uoo/j+9p7
ruESkVRiujqHYkTJSQLpcJV6YNHXRJLN2WQvb68CaTpIfikOiOeB+86lwt9YgU3l
cQ9o6+t+unQuXswKxPWqh9Yw7fLaZ4bouEe08GPbkt3xTllba9aKIAO5QeJQXoWX
B2XVY9tl+UGhLqUGRolBQyCzUINxbFSvQAJWqTBCEmFo6MMZA/R/MokqHWAe92+V
R5MjT3h30q07QDucn8US20TXOQEUlT6zefzzwQWcV9HnGGcEjyiKyUR6yO4aL0Lh
fFEbif6FUBYyuyoeJhPPY/t8eWVXH8KGAsnXl6VBzEc2gRMV181ln0XsVUm08MPU
BS+gijavuLRf3gs6zZdcn9F/6JIXpPGBiczz/hGyYqMwIiAe2Hh9+O1TtmhH1H0d
/kVcExgPUgaY+SJA8tta15/P3ZG3KdCgEh/hHn+R/rnJSA2CJWUNfVd0j1VuZOIW
Ch3DEtmHIXtkudiglQnEpqI11GZTOjNqS9noCsIvC1j++npTL3NCZrp4omdIKVOe
AiQKgR91phBmQi/vdSskHqw5w/2V9ikXvDjJRj1do6E+7QO9/XUKp1GHH6vUQPRN
yKvNckpb9XajJxWCJprKAUX4XfNjlX2bPBadaccxjsnlZrBgpbuv0rpuwUOKd690
2FRXTtGikW9gIYcbuahqseKodLRHTeDfFsuH+AlVeuqmot3D/Mgczfs//KxcaEdQ
ByP5KocjKAtciKqb/u10EeOJ5UumcXpEFx6FoMHluTawApG18KuY4QU0uZfZqNyl
GHpf23GnqAZgVh1XbGfALMoOB59pEV2FiesnHy8EXtjkdPYeK5AX5zYvfBDmlYda
1w57iGfIMaMfsXIXhPpoVb8RsQvK27hfA/rA+SyIfJXHCfpB4wU6PhHO+8VrAREQ
ozBi66uYgNxuEp9q7kJd+UYpUrWUlcLBOh6tc50p+OXTFG7rZrjw7qaF/7nuP6tv
22iPVICGaBO7tkF9lhXuqCN57jbbbxmz6OWBpwJOM62Sw2ZoUI77y6kRx2+e72Hg
O3sDsASEU+a70TTbA/ABtA3zaNVflmhsN3ZxQgGF4BJmZmTY0qIJXjD28Qb10yi7
X55eqHKFllV8Cn7WwmLMopJ4ize9gSkuPLreWR2DfjMhnzrHG+8ww9eWGnbP7KU4
m/6mHqyVOc4h/lEw3lWgbby5U5WsRfrAVDV9mxZiYk8gZv4yqz2D2TU80oNEBr1u
p/evHghn+2/G8kSMCgW3eoscvoj1gGS1TRq+hvGgncCBDZ8EyGiCpWa3ngC8/hqV
BcbxKjHgi87c5A+fL7LUAVfBdT8dTOWdcaueVLUHZ6aNQUR6N5e4cBewPchYPRd9
kBj+c4JkpV3b15CKbyp9N1HdiZ6AX3IdX4ysHfkdhDS3BXYykAdB113NJDEjx5jK
umhWc8YJ9rA5c5/e1tVtL3EV5LD8a/j/HolUmCt2+HQxKHOQIlqB5zDvJJNyixeN
3LNc7FiEJ8qcZycFummr4j2ebzchxeQ1XRbWEzLcLFMSB6DJkI/wc4PakZuWNale
jYSs0d3+Pp89fiZUUG1rSjSTClRPyheGTyW+0PsHkNSTp9mmCxdihHSS8bvAZfPR
M95QxXCFCCG8p4sSxq2OwvAVb/9xyoESgL+AzpPun6jM+/+89vrHwMR1vSRFLZq4
0y7nDUo0HaFz62KPwMcLNVt2AQBZyKnfgbaew98G+cBEwsNRIHkulcSXaIhRrbtA
lMhJRf28LUGCq5bs2Tr5nf0HfGzJfgKgx5ZgPeKV+sSdk41oY2SsmWafpjAcmcEv
6UI6+MIOvFbJeq0tAnUL4yLeeDdoe47ZTIIY9slcz48hsXiMPgjXnSBTtAMRlCIo
l+957cuittpyMeCYNhdVhLDIBG/b3NMRrmhg/onfaMYuuXbJ/nD+BE6a2eyKrPhu
wJ9zTxqoR7hk7KHLkxa55waNuSMJNCWPWAHGW9Skq3Fjpp0pBYV7Uh83lC/qO0j6
uAlGHTwKQv8S3GaflTKq//LRkgAXEPQa9fOVps/dewwuLE1xrBOYByX8ZeYhXagL
L/cqT5tlN2gLHLQWQx60BnFA696QkvZb2hKeAe2pbPtKcPpqTKlm3YCzLuOp4bc+
eTZ3uuis8XM942Ryk4WN68sVG56K/HkwmADfvzqadnin3qoSHX4jNyrb02QqRRpZ
pSONVTc8HU6uRILC+Los7osiRKHv9uueQ9yiYDPO0GF9z0cfwcdIH/mNrFO/BEVE
iMKc4ZmQBG/E++4GARTr6qhqPoahznqgmfEDc4NrIdhtTFB7rneR+ChDjG0Sg7Kg
fw40df4hoybEpHKSEHuHxSvLyVN1aeruYkKTfnF1ADxIf9zkMseYA7NzXizx5Rak
Tib7RNbTc4Yx9Yu0qqxGiF9keQC3eJwOa5GECVCAjtvShUWolCvqxQ0c08Ynjej4
6YxEROB3yNfRRF54XClR/KdJ/DmyqoOXKrt/DnwGJJGT7UeRTF9aPckVJ9NUf7wu
n2e4MlW1qpVzHTnp6xRkwybjLMgn3DCeAESzrqD2qB96gbkQfepoBA77dMXtrzfL
l+xmYg7v8RR31vEfWlbvasy7KUSmH9935nXDT7sly4bT2WPFi4gVJDSgsPn90tQB
dugCVlh5uvTMNwOK74CZQHJ3qwrSIJBoWnBm/COyRhGSwlRNvmEmVPKp3pjPQkJ3
F4W8aT22PJzgIw5mDGfEz+s3pxqAslGc4oAFY1VkXTjLtMZIihYzB+Eqc5ah1PLR
bsC21uCMtI/H3E48VInLKBXlQpOcQ0xeXSiP9uO6PQU7WTe/GSZVV0QYoM/WSqZI
HdThFweOKKc7gjEEqjE8inAFm8+vEmq7YpApcR4Wgal6RfZQWNAuRrTyUaLbCFfp
kG66a4kg8A4v7f4XF91gGNPInNNHT/xWEpWaE2Qgntx0pAUUgJKd8BwY8lLWXTEX
StjJ5+oHwryyw0vZydmy17RGIWjQqaB9hvhhmUJgNtYoNAmLcIFpX4fn/WHwyG8r
JAyrbavlQUZfsd1EXr8OOvgWIs31i3oCd+RZ3XtY1GEeah4jcY2W8T7Po+llyYiO
Y1gbUW6uYop9av57s/V7wlRzwRR30b3Z5X5rU3CbJWk7LSZnIliIvwjrQKgH7sYs
nFXO037IU+HeeYctIzMsNwN50pBJ+ao7Aw3IrB7t6J1gE05kNCqbkWz8JwECe09r
FNhj+p88l3Sb8z9GrSLGhTmFgfSx0lnx215g38cnOYevonD+47zOPRFsep5sE8Wz
u9v4ggc+scu+QU0amhi8TBPee92NGvFzw7cFsYXvpmQpbKnf+VHVCPg2BkLp1BZ5
DS9u+IEsi6PC8EcL6EKTtu3oGW3paetFA8XQGWyZWcyWwnkICTHO0LUR61vElPs/
H0qFTl42Z8lu5N+SDokM8WJh0H5iry39Tg75sj4ycgiC/MU5KCWVW4XeoG52r78L
ZiylH+hMJLLlGU7cuXiqJS4N6hAjD7u/gmNvbw3LSUfLkXZXpked6l25ONMUENA0
62Ni06q/xB5X7B7k//iUAgH5gtZgarKsuKaBbxliFW4JUjVJWhnU2lEjSiCQFlAk
U0tT4EVJGIhmMej33Rar3paBv7gsB3uCEaugpdiAdnW54KqbaBIdviBtQa9ECtvF
M0IsPCDF+WbTNM4faaOKb/eMRbFXsblKTt3cSAcszUstLlOrhLZO/sJsZzm21o2u
gb+tBNuj6MeIzxPJTahaCndEbfOmvoFzcZ+/+HstFJq1MuRcvWzBbZnr8ofuAUZr
fUH0aAobifUt4Vcrbd1zIfwcyzTWmRW3n7yd4+D4YQXMKJ5j33eY4o5agZULR7D8
WwIgsVm+CyoJok+ljYhv4rYJ701zxuZ4LQ3q721gLwa1iOic5nyxeIdq3c1cJ5HE
5+BCLVRpocTGBpRXc5dCLoH6J4UjDQ6Mffnbzy+jBsyf1ZfMfnzrdHch0Hvxn9q3
Vv0k1/HvTFV9APWaiFYj1smDTThDejWr8Sdmh9d8Rr0RkmuiCw1IMmTpvmUnipnK
mbJK7lZNc6Uyfj+Q4BsttAz4DlVI0oliP3a4laVXauKLlEnGYjFQMCBxG/ALssyP
7sIUFN6tDiXT2eftK+vn1Uj7PnKdeyd9iK6odq7+kzQvQBKe1tWpbGPSfIoazxeO
VO35AEDoaI91XIF/A6bllsGTUBJe6FRJsf4yyYapDVYOfHAthv/fZrNr5rEP1pWH
F/+uEd+SYRwCh5pl2AA4iU+v3hmt4VONZkL60Lv8oCck/2WtoLgPlLN6wXVn/Nlm
pKAaKYJXwhdyy4kPSi3hEBowN+euve1fFIFtuMOhJpQIs0q65hGHa2qr7XetmDy1
dFdhuV5tHSfg8qWNaWbhiKqcZ2BIZ3+H4+SoZPlghi/4yz4djHqVob6VsNqJHZyS
/gVaY+Rfc1KWP75k6fwE8mZxUYq727RJHfHPUfCWoel0vJ89kEgcM8lIuAMLa5o4
Mtq4euEcS7CNJsrz5wX5TNhYiKxVt7SFs5s7+ZkfpumeW3XcbO1PS8ob3gxCAkcN
QryUborPlxviYl5LvQWAIRiATP8dCwvniapD5Q/ZOmeiCrYiV2kW6JqDxGpLJpRW
0MtR/j4rALAVCdTeuLwZSg6pRaD6PGKG+5CUWvG3PLATZKKn3U+PpswE5ZQNuZjY
DjRu6xtSjtIMSC31ZvBpfu99xcwQVXRMTTY/4LPy9XbuEvSbcCtityEnbFAnwG55
Io32px6xCNHn6/NZd/rwTlpWmg1weUkcebMGyhohy3RnpFSlPhGl2Dgl4bdIyjml
1VDhd4NcKaa4mSOCO9rTca5mqZS468sQXWzxHUeQKQpDj1kkyPJi55l5mlJOBX74
esTkKgXCQE24Ozau14MSYbCNgyHPiB7qScxq1WtMZ9vSd/DZGfkWZ6b5aEIwG4Sx
70knXdY72Ue+IQr5n0KdOHzXOOksFh8rv0H7k+cpVe/bi/+PDXr5yGJ30ObIQN+L
ZeeLk68YGjDUp6tMLgfY7hoqPJgChqbfZ8GmAx11CTj5QYN+Io4HleR5/g3YY8RH
UAVj5VSAAeK3YwRNvQxMiwb5Xn6Hzosnx37l109PacFyS6EPHt7YeS8GdmD9ZwnR
HrT4WXznoDiWp58lXmp21y2wd5ruZLsgdKlKdikr/hL8gKH3yHy6LJSqC5zvHrCw
lNFhkmmVxLfDWIA1tK8A6y1gN8xL02UucyAELq+UsarWEw6fGNeufrSUNfWuW7Nf
MnDXxZO/O7kag02G9lbli3HA/DvRKHxBLtdsUuQ+OoEGiXnwdxnc763eBUGwTLnD
5mFh0eJgwFjpDs7cR6RfiZLS9kYFYRezyi2w4lut41ACg5/7y+XULjiA491K++6c
KS7l5R6d7DqLizKxikPJitPubeWpgr7MVrI6no3hEiS4wRs3f28RXj5KrZlojjI0
dmMKBqBUOxWfA1OX643/SRf9qn0T2BYaYyjBlRREKneAms5py5+npkRw7cffB41H
24EVPAVU5h44YZ+yy8mNlih/wU6QXQofe2aL519GsEM7AUcWZNWy7nqfkE8dc+v1
9vnUbhMWQiQY4znFZTexHqjJA1hasRpF58igaZUCyLjptTjEg+jaYAUB+39kxf7q
fD+ouVTfvBuoKSCsKbV5Z8xwGePgnmWRsg4i5MTeryQH63uXAisG7T/Z1dLNxodS
z9XLFKufhcgG5aOeWGBGEQF0kvYP6hwFncd2kmJCsxR39RU8gojoA0/qXQ56cLAN
c30MGfXUd5KvfboVxSrRPCzsSeHE8avj7AXO3DX6vKGxw72dXZ5eoGRXX4X2E7Ke
YsGsrWec2KTzR1vhSO5ao66WT6sIkhcw9fwb3JSttBnd4y9atCiwdt/8LRtxuoT7
wmIfPm3ZP5iO9uqd1M0GqzLeGsY2WJZ0QAImjJO4fZrBEfMT9BU73lQWwuaC6JZp
KjiC83RLSfJMPOPi83Nzy9ze9YF4f9SNe2oLMQ3I7hhIq2Fsa7vlN2uaUduwuIAx
3RqwKymfLTC16WnxDD1+I5Fism7OX/dY70hBVucuTXHThC73n27yjLnYskUaYtzg
XiJYortfmwOPvfv0CYXmk4HyCLso4L8OpRjLX3SuucHIrjLnqOQ7Q7gZ/1sCgOYp
LZifGiZzz3wcKbVfC9r1D71rMxpBugSeMylTP/xy7QAPAUCabmoznQYXIGQ2cPFB
wrzSNazPlVFF9AREn0MuB9yee1fkrIGI3DVN9wIesPWbJiC/GgE5bk1ugAAPiHJb
kAc8gLWI+COvCDV0SYu3bSLL+oZEvcUsYG4erzkjEpy2/6MhaN5ifPVbt0rmLQ2n
WOiQ9zozQ3q7Ihu25AoieI2zWgefCnwEu6aOl9VOwFtwhKZnUO9cNj33JJ40EYdQ
EERwtErPcs+zQ9d1wiuhnlB1KAAKQpNOimi3QqePCcX/oZJr4ej6BGSs8fNPr9lB
DFQjys6ATaryQQAYGLKs09JQPUectY7Tww6HgYzKN2zra+21sJLIZTQdIYr5/pS7
CxvH5vHwtYqOcKcU8O943ZnO8ul1soeSYHvXZPfaVCN49Vb6H+Gh79Lij71qsskq
HEn449wyKOf6jvdXKaXIxC+TbcJ7G3BWAeEYy48Y4Px7a6NMra8Ym8TMZCeqoXIZ
in9luWyk3XvUIoZ5dKIHhhZJ5tJCTYeRHQn7v2zRRtHlvHCVlDq4bIivfl9MtyPI
kGv6KnNZCv/5qx1cPUn5kyfQp5MwKljF1ln2S40aMooFsUWalh04ujkIUSMHSicV
k3H3ORpr4Qo3URxJvKjyVtJb6lTfyrPAtH+YC4x5iRYL5Pi2ZRqhIydrrrx0L1M0
RoenWki4RoLcYqW9FaARtUk0SteZV34ci+LvZPWXTNqhfnYJD7KeWl5PvWnf0O5f
ES1KIpmYoZ1FOeP0mYUZ6N/peaJUmHj0PN6XSc6u0yhiMt4YLP8XkTOlbslv6+nq
JXsO487h4qs14lCAgd3w9zsvt7i9EPh2o+5ru3AXKm/5x4Fm8mRtub6VlsZOFKBH
w4BXm0/sEvhkqRtLIhgOd3q8yzHZlSLS9mo7nq/VZMVyYEpAStG7Gn0gwYqb7dmc
a8xBRns423pamMLngHqU6FfFcRW4ofBAL8+nivUD0vEJU1Qsz2eXYJxrmIdjX0OQ
9+r06+BQ3jl5P5wsCLa3mZN7+RNvLOwZEyQPfpnASR8PNIqU9EvDOEhfjaICiQX3
f5cl8vKijY14qboc/7pSKv4bg3bPIaoHX6B5JJBhymG6YzUM0LTFgku1AMVYO46S
x1G0U/Ni6MNHqopVxtyMfO76cpnMrwJps22i4NHw5WEzBvMjiTZySAHx7vVchp1Z
XsR3ipIuEP4WLF2UzIpcpY3tBtBB1ERUDTzdV99SWIoFRmoZV1pcbdhW1HUrOIjf
wn4pBzaN8sQ7/BSKxa+x2mTSyvlmEDKLnO1nwcbbmGBbRy4IbLRCmKrvW4KZg9Ot
ZOX9Z3s3IKBnkRcj9CjHHUGDXXPVTs26XfhdZ/vVi5IcuNEKyEl+dvN1+g5iEgdm
10Epi+sHZeJPA21AeMXVkvsclOkjFZ5UZte001AKY//1/CJnA1YYmAKOv9qk5wYC
TJfvwFo6bTQQtGty4t3JcmNnMJ9SFiryaikueXXjcyMocvheoOJ69tTVpS33r4oA
QPPVyRxcQtMN71g1UcV6O46gL63Qco5donNxycbj3m+2BTmH/bHqnryMFDITn0Xd
xjyevMkCW7UifxRjtHZnhMLBh+K+zuDXsNPqhFTpd1Qf+w+z8emXlaSClbVxFNQT
46ktVcXprD768pl4DRaSpsBqrehAR+JbGhtEjFYLpLSCWJvBniqVT7yq9FFCde7Z
5WfdNU5VGKwMxQvAFeD8cPrHNNFy4C44D20xT/8vxjdiyZB7f+2IwfXO5MvEzyr7
eZcG8YhXqQXG9FiPmUC5/eQkFIkahhbIG8UVCIPgyK4KFghOs6MSYcviowIUZRxt
opTdr1TWsTGVZZqdMarktX1iddz+ZlttGTCopVEvRXMB0BbTf+6biVfL+fe5FgJg
S0CqOVR8R8Tcg+ZoXVpwVQWaT1zqN5syplt0IoHOvcleAkXxVmUffFHlllJ0/AQp
QUAapyPCGV9jGHqOCf67wjDX2GQpjHsw45sQuDu8Xl7X0WcPhzjnvklDkmTsEzT/
Pwo8GqbjzDidljfL1KzgN2QHFXT6XaoNbfEfKfZIDH7B/PXgqlFMAVEZoRkoryb9
jrKW8PJ6esCexFvxQAf8/ak0fRTgB+TQWXB7f02iEOhwI5b99pm5nvnITVVOSGnG
91Zf9wh72lwBoBXw+enwRfbANzjhHAgTVbEbahAaJVzGPNNtGOi/KzVn7TTLtVvH
ciRtoBfnx1/IVW4LhMtWC1rlFgvSVP/9y4sq5hgoaDfFArDNfDooNqAH9dx6A/X/
vz0b7nHRTv7XzhQ8NCcoB3sJhMMUSVdXUCsqE6qgcYov39E2oNdkEXPFnEc05W9P
W6pDqxGfq4yQIBZBLEY1MUZYPAlyX5dwzsAk56SzzpSnhL9VL2bt4vCVuo/GG7oH
GfbCHBzOyiHDsNItr/+e6SQKTfMqtnoXZgeYvlSAzakSW2wBr96w3nHRE+WG/UXx
VHp3Nb4nGQRnWl0U01g3TTMqa0zlhXzlUH5BjhiX3fQOWGzrawwdMsKVsbtNC0xh
cDRj9PQcFbnVWz9tT09Opt6xmnx9yfcGBytRVIwgQgd2N6PAoe3vTQa4Acoy4TOn
DHaLt9X0t94mHkYdfu7Sj/sIUh69HcMdkKeF+Vw+CNkH3/yewkf3G8uBrKnHCsOR
Ele1qk7v7PR90+Ys2329UD1mtdDhMVYYQTafYr5KQS0XtQlJDNaHz9OcYwiDNoh5
Dy1UICRW9AeiDpuoYIOqZngkEYjgO2X0Cz0HEIU6jA2bNOeU7kqhSwIZf1YeOsS7
72ASBIWvFv25IVbKj4kG9fm5WvYOS421advqCIzkc+VA/Wc9ZFFz22a0P/o0iOsH
jo5fdEw8bQefeICHSxTr4kQeTfO8DT6d6TQgYEN7wZ8Q5rPfap4TpPlWV+3dxBkI
nqVUVsNfJNltsjOnlScUCiQzpu5+qa7NDHiRuoTEPVtzclDVRh05iqaolpNs7dj8
gNeQHUpd6B2szgU0UY+wQcX/KRBiCkdUpUVLpnOQFClofPgT34Nm1kSUc3xb8wjY
WO9aZZhL3wVnfIls9HXH3R1WjcDqzqq5j8iRjXWL7esDyLL4llgnYHaivr0ngN70
UF5tJI5SgcCD6IN4XfQ8VXiT2cUBJA0MnEJymuq92N5ehssdPhpfDAR7ctx4hyMg
2qnmpys41UrrZIuaTAoOi/o5ycHEOonNAdxJP6tD2NEZZG/eStUptEbaiSTKYe8L
ai8pnURf78T7nt97bkaRrmWVEH9GjP+TSSjgGF1F+EEGms7+3DrHipm3uEzUKDEU
XI3Z1CMJakOr1H8/uMSXnSOknmpJmL7r65X73O7qiDfjBcavNocPF0hpAsLWp43d
h6acqv4dIaExUEEePcJ/qGh1aKGa7sPI6+qSBfBTD0fTmckL+fJYemU0rR+Dw8sZ
Err0xgADcOJK/BLnD0Uf4cC/ledQrBxerHKEHLEM7set7g0D3YxJnioHq+BtFXPj
yDtEY3jqRXaTPXuhcBdBAb4FhbhIVc2oIrcAhhLPpUtuqwTN2S9eHrM9tG+u/br+
ApEEZExeOt8BgncTeoKdxTHokZXklFQssi6pgorZoQHBJpJAsiyw+/vVbq2zdEmi
RW6Wy/91Tb/xr3uE0Q5uDJL5bsnODofGNVE97w30r/yru7Okl/pN5GekF/iqgu6f
jjh+fGnlTmWwwRpTUz4BCZuSEfqxIDxkesxkwrE/uNeNybzHb9WeGqMwCljQTknT
yjQc1tWQnul6aUZh03fu7TUhiAYl9646Twb+lCsQYc9Ou+CZHut+Wwec+mySLLs9
B7xLuDFORgMtYDY+nvrR+e/IPJ7GPTEAj5KAl8qP51pTvCdK6LPWdXQKmpcw69MD
S2nIBVSRJvkctnS6dAAu83q3AFSRWCbGUuH/QqiScJh5wqlln8ASNwzAvq1drW97
CnTa+bPXROCobGv0CMqF9qZqAwGDR8anRnoNGC2kudnqnqio3IroT1hvnmxzFJ0n
YzwnJtBG8KHzGVhMz3UKbxuKyN0W5uuDAe11vRw3eysvA5pQFGfHQcWzpS5C9DL7
oZ+i8k9P5h0l5/otLoS0M93xyeyQdFjl7tkbxpNtEGcyTjMRFTr1jFL3yR0RaxNV
h1O3VgGt6IJK9fw8odslP6mCBMQWj2xiaDJZgbZo23WpRhyhaKJ4x+6WlMtXUweg
VXwy9rKFJO7a/H3qqqXlvJ8gx5gorWZ2QQig+ghDC3vTFbR6M8v/QVBYQREvoC+v
wcAZP1IipejHtJUpWJ3CRApJfRTTblbp2V7c269eykIG5nCnjAXJhgnb/kMeU1XN
yvMwTTgRFddMP099zKtziANDrtugoy2bv/Sxj3D/p5FoRC9yJEKQ/KjJg7TvSiku
rLa2ZWRlU7ZFqoRatGIVS/wQSwxfMEHL62AikukykS96shFeY5LFy5dQUbsanJE2
o2LIeAjWxYn4DF31YB/CGPACEjPLt7ChrGQBKdWaiZAa1aBv4rrjDqFZ19gQI/Qa
Ml0s47mZqn/OPLmwltd6ddCge1API5vao8OGuG28+dwlgkXw+Q9iyM1aF2hUNNpM
4rDfqC2AknTDsAXee3dLIQ6xpD+UZ/Nno+4iDq8aOIooqG9sbdbDq3UParw7s9Lu
ZAx4LQZQNgZ65dKVvbNXh9JHHD0w+VH94E1QdEAwLT9lr5Yzzhn1cW1Wjeo0oGaL
y/rtlx480+vbMVtAOb5zredKyyapQsFk5K4wvZPpRqlRiVOxgtD2WJleJigjbYgV
nckvfKMZrXqbGZZx9hvMy099LVe3M92scgXYSZMTRf4Di6GkmoOBTNcUv2wzhVG6
wzGpzZKCmuLBddfJ7P+bW202a7WzI5+nBKurJWFZudXH6SvZ8e/4B8GeNk/zUYuc
dGVnWiQXJmZct+5J1onVBJ37EDQr7J+QxQRUcyUIyNKPcB19sxSE4Z50Lno1gpE8
P4SDC2fLZItm/dcjn56ClB1oNXpFNkSifQnMISPabOQY4VoJ0d9sjkXB6Pwy8YXA
wy9uT+xjGrhwCWxb8RzoI6D9n0n+wV55fVeII8pBvef4tjfT4obuy+Xr1VcQGvkl
CWeR7+KLyp2HUNCN9ifR3TQVlSlYfeLNPhIeei++hlebWmafERBF1WD/VMtNgG/P
oHUV6i48uKvXHlMzE6hFYi9w52w0j81Tas4hENLBFj+qcCU/jZasH5yoQBX7hEtm
wMvYaOF51Vj21vnmgibPpXJ/hWQv0WJLu6q7jZWvbJdMnQB09vkh3+O20lI7jYe4
a5pp89Bu6pph4+BAN0ZXSAk3FW6vexYwu+gx34zB/yillh9Owxzlb+3nxoCZp/NW
/pJtFYikhMdvrRfG/s+KTYI4nruigUXLb1sDwM/Drgb4bKWYgvVI9q1ukIdiic2d
0HuHWrdugavHuexi72ZgT9NYSl3mxhFeSyTvwPPExB/HD29j6uexvp9dA957kipy
1Vyj4BdyYS88i0uTiMSKZTqFLauJN9NxOrSU62V/z65r/i26Bwsvfm/bntXSqu9W
mQs2gMPh8gamfh8AQJ3sSZANQ9q6+NGdYTxmAWczhYcu8XZYx/wKpHRRGI1HWgWQ
nsmdaNCI+WrFB0ODwWw4uKEj8eMzh0yTE+DLoguqdv+LmLrapbZFgrAGE9TRoUxh
RLUrNYnxDkJTpkCqk11/bhT6QJ2/XWfLH27V5bgM97X3igAMbXZ/gyLfZDHdS7P7
iDHQubhD228lw1IVuud1jlt6CrZGZQx2iVZoRkScFs9PPPOD2AqCHWnaufy6kUqi
F3fc1iFMHjEDtdolFvAHSVvLR36BU/ltUua7RqwT0bYvHO5ST4EMOG/HVSFPJOTB
M0pmI4V+NYzvYg82wKW5BAVdXDmV4jT34254mSWtY6QZ+Ag0h+BI7bJhYYgtZWMU
K3WDMFVhwxnQHMB8YcV2+CWeyXNrb74tEPnguE10reL2akU+iYbfGvODM14+wlGe
70sk+eFwq9OdzV5XqCptfaFyWrM7ZXpCwOZEqfQwcm8Ub2wx/+wNotfQ0dE9sic0
2ZanP9qlZTEbMa2dlTENOc2U4eY14oHLZ22pJwT4rfC3eoUUMXl3KDzEhHRvS8fH
ehkb23hDWXTFm0uAQNyJok2AdjyrXs2qKAxEUXiQWhVemNaDIPQkSFQle24rpCDK
navBxD18YbZpjFTRRdSRzC0gmr7VlKzr8mJeBVzPNgAOk2oklu7L/2EX2eNUV5kH
kZLJSTbheZdY5ibPDPk2zRFGR0/O+Oh1bWWzry4ODSYRYtHrLcw7l2UFdqoDM5tl
xtqDtF7wMtkAZZAw9iFsmPUoGPVqaHqJWWlK7wxlIA8PyO/5dEdaJ0Kn02/88Yj6
ph3PqJuUn7m1502AVIBv22twcqyR4jAHjzKdA3mWuIa9SUJpJ/5S2slxj8KjT/j1
ugIB1xqvRKIh+9biP5gv2LWzqyrMgKj1C3ggSyrzYktEWw/4nA/k+MaVp76JgCVM
qD3y7eVHzGyC9Hb83jlTBGyCWlTPaeL8IkV0LZlAU2fUpd0lfgXnT3fPfRrfjQQZ
P1VpJGgvlZSwOQoi4+wb30ouPTbq7JocaemYaMLi37yrMK05iP+ftvVFqpx7Jbsy
8eMCRAjC6SjvZKvuMLPOkoAo8/sbCSfntUIBg5T/BLGaNqOqO3GkcoPJkYH/fmVF
aZLhjHEIXKLVvkoQPGR6okSbaI+cFhwjtW9OheTxzBlng2YUsOjgTSCXJtOQovvV
ua9JEzVlC4DHh9BFUImmrHUC71Qd6raL1CO0dXdxNWOKCdFIPT4ULr3OZueKtXeG
oxrEaUQ2hXZ6MALeMKQfmJChKOrYjXcUJKNYjIFW/2oj4FqRKw3rplwIxMYQou1N
fAG5Td0nnLlBXnn3rPOcIbTffMR/hkxobzB0LTtFzZZWyfRUrjozZF29v+bu3VJA
6ep0Cr+hvKPPh0SMXDhzKsMhE9dvKh7t5obtJfnWjQg8XrWFlwHpOQOiie5Acbey
6Pppu+fShIih70cnutjolWy2aRzsVZ9luJv5cJTkr8oEKlTThD1nMEqFrD3wLdSv
rpGUOUZZC3EJzuDOMjt0pJBV4FdIgwsBpty0i3BH7zRyhMNxucWQ9rFEJHme/3hm
RSYtKeRX+IfAbUtcRGvx/ycwKUXstPEPLvDoPDuo4mPnDkfEAMQK4olPYUwalv61
l+9a4oLWIINJXsMzfKSHLZq/ZtlLKf3EWKkfV2sxb35kiFACxtp4Q0M6gVzfw1dL
pRRQ+aGZRg/u71rdSAbLyLT6nsLGkrpcGpNtd0/bkf7U6RqoJcI9A9mJNEjgQwXl
tnCKEwPOfKLoz2SmUZg5K3OnHPtG8im6d861cU70kOiIfRFIXNAwEdSbuqaKGYr3
mKhEgt/tvWOeFKVPw1PVln7LLKE/adUmTrj1YQNCQlrrS5tuQSnZk97YOwdRBO2M
2SB8v84D4QVxDNgFUADLn6n3mIMPWx5v857rqYiQu56sTdXIfNAQXbLcxFNtqphS
GxNcP1wVqYrjTAFoQj98VDZEPycbkJU0GKrPZ7Ldpy4waO+mLFrAUN35CcYMpkSO
rmB3++SZcA6id8K4jWZ/K6Ko5nuHjIXF7xY4aRYM6xp2y82PwBXmJsj2dV/td7Xt
5afuwuuIvYMknoE7QzssWL4vf+hN6ap+8lqJzJWspuEkkpb4vwlWdLWph7lpgvyl
5EpXTcopPRu2cT0zBJE9U4Ih+x/HLRu9Fz5ivx/49wIvCgaOqTpDC6BIlkfMqZeO
eVV1oby1UmulraPGdWjbvpwjjQLV84eezZIeKwimKsRhkS1prydYWh3DVxovWrBq
NbC0kvlPasKYNzZSzt5IDKtJfrZQqJYkaWFXxunnw+GY2e6in0nAlv81Q/w/8g0J
wxvq/Of75Vn6W0kbdewmHvz+Za2VoeOJtPtXyJI8a/UE+pqZBkdq4I/E9SCpFwY5
Q/UKIr1aDDWtS7146vBalvkuMUtDuAj7s9PWBMXZ0g0YHD/lvndtKE4ZKURUBUHe
/Isgr096+2oTxfIuS1bWJSLkZHMIIExqZlGg1cMcRZuBaU6rcp96Bm12i2N2en2a
poBAqeOxb+VA625lMj8k/2RyJiS3DFqjnGtK2BTMLJs/octuvhUdc2jF7U0P1+KP
ZanPdTaTaBDnV9kEREUiUiXRYnsPUYkbf1/B+kL4Y+W8tBp+3OeX4b+rLCxqKWcl
nbiqegNi/gaupcwo/dR7V46Hi7PMTxTNafxqxlW5bLJopwMiH8ArptNli+z17SW9
x7ThP7vj71PweTs1WxEtlCNWIhLzs4TO+UHq1L4HDunUl/ymA9rK5UM4Up3VggSp
lq1qmUmilKcpNLCIPX9vOl7miVNQZ4QQiyuMTLXqtWMJeBrmEt5Tfkg2c+1hUfHP
TxQcf+0HIi77ckEJMfiMfrrySlYyZPtFWS+wnoClJwMdLv70kYM5BC/jnhl9GQsp
07u1lUxmp6vYqZkneYtRWvo46VJttgaeXnmIO+sH9jrTh46Oe6NtQmgYS+pkIba3
GuasCcf5lx7g61n6UUmkaAbBKKLPFg537MispV+LlGKCVaopWC8yNEK3p1nue0s1
O4fynLSrQnkbpSTLHBjsmBa8Jcs9Ays0Kyte9usQN5euO/EX8iIfaw9d0LpGmJIL
Y/Th9nLYx3pw8HUbWvF5fj4oJXnk6hHrtVMlIpl96qpoptiAbkkiebtg0x/99HMj
fxRPphqDfmKAWX8gg03uhz3lhtHCYm4GR+6R+NfAtkngIR65CCeQn8tl+442K64D
ZO8lLUv6ZnKZpONCre6xJjb77R/FfJkeatMS02npKFKldNo1O4S2UtQ0KgHKOUWR
Sjw+mRM3ohmQInBbnOAL799uWGOXJc3fTnXlfzd3jxxyWqyczg1ssDHq5Ebl85Ib
U1Y3ctNr7Z6do8QUnueUWsRKOd2mcLMrgDIJijCO/O0EQHETXvcasQCYOwLhPeYb
/O110ed58N1Jnd6bxsUIi1SeTZYHmrEl66kpfULk7ofoNca8PmqLIQ1RX3F0NMXD
FBdz38jLG6lZb4ntCgNqGs77qfTMcMyRYObv/E0U+SVUpmyW29r8+2OiM4BrVCfR
sc6d6AsxRx3AsjiyZP+Zwf7Nh1DzP3EVzdXYD9d1DRcVGei0/03qUj62aQoqj3lJ
LzQXNmml+bEMJO7iWLe1kH2txfFQuw9SthsKSIpo+iJXjA8Ga7oX7FYBDgEkuusH
lQiLL5bDR2GzxRV4xwtxqxePe3aUXptK0IBP6yR/YKgydyaRL/ss8cOt2XKXuAkc
W6QdUtpak7xE02f7P+3TloS/yOUkuqygxWJE+oQ/XsB2YaQwN+w/2JJoXtudMSAe
vJf1IJ3iyT4WWZhKMO1I5+7OqnTAPBfDdJ41o6dM4abzoK24jV677H7lVBKYRziG
XetquzMjn8+Svzx5lnXUHMOlYWojedteBUesc1SW8NjS3y0icJTW7RzApN/FdMla
SO/fzl+VlZNAElOz/P7aA7BRND+I6FXlyOV4DLZv9PBYXI+bsM5UJbYglRDmv4yw
DBFkJCadqOzrNZ7fwuYOAp4I1sngJyoMzTvGUhmH2d/iiRoyQ88Tof5msdK6pduZ
hCnfo73thE1Cq5GnZRV6YSqaRcwSgXNIKoocLli/D/fQbRxLdQxMqpY6UvyD+BeZ
ZBdby5sZo5y4Zu9kU8ta84gexl5QQq3dkuEyEFQcpBzlxe/mioO0+myM/bJF2PwF
YMQATXhvQ13E/o3DePnFumr+jBmwda0NP9uqVU8cv+wV7v4cvX6B6PQz9zkx11Ss
0J9gittrev3opUXQNvf0JhWQMWAI7rTA8yyMp9n/fImVyj1PTPGog2ncu0qX2nDw
0ZTstopRZ++Wz98rKsjBMO43fJY9teWYhyMYdraO5iL+vrUu6Q0A9uolrC/gmv+a
JBxmS5myet+Qa2oClXets6fBtLYsKVpnz6jjAjZYDUTJXrJXF3BeQmHXHU/MOBS+
hq0RvFj6kKHJ9VGad8NOKsYVC1dYu8QF4+9TcSGnlW3w9Bp6auoIgowPOMkhG9jA
IBW/p+2r3ynvouJMboqVxfUR7QzadEEgGellMX9RUTlcxeeL60tVaRPtf6grB1Af
IMjqa8dNdIBWPDB7G/IQU90syrhHoFz0UKjjq9HtIcYPlgXFPRkC5cNbI0iJx7q/
qUQW7uMbQkQkQ4wpK8MJvf0IQ/Q9+w8L0OHSFMs3SWVaNPp3BkORFoL0e5FlyCMX
Q6g4t2dC/svn03oIP6k6yYsFiS4UW61mOLCHB1tyMdHQQlbFqDERV3A47P0AiW0T
qpnThkMWVoq5s/v8aXR131yY9MGYTaLBM/YnkzAOrikFzRg00d+bLkqm6CeA3ZHW
yf7WgdPgpOkF06daVcd+1oICA7/45pU9tRt7cLAtLWT5hLU854zBrk+v5DMgV/Sd
eE054mKcnS7MkQyLznZx3wm7tXlEeta3oPaxCUg7UT7/PuCLVIn8upeSKsqWyacy
hwNwtta/NEYN7CB4dL8kGAXKC05y+Gphv3qva+v01i7QrBSJUHU9BgNiW02+TdiR
NPzySmU/0K050Fcz49aFAUIaD8tcAdkqJI9271H6Re1akXQHU+qAHR/qv0M45Lj2
0675pZDHq3XfwW9JLbOJKNRMZvnbiLPiT6oA28Xr27pCo+T00IydA/gOEr8ZPj3d
u2Az/b43WuMbVeX7GfEhXop5+1wQn2RCTQ5zGqiu3eHJYQ7tcgZsZDD4KMOcLH++
EOpijkxFhpD98LQS6aiU+LDLFEnxVted9Mpqc5/2eKqXwS/t9wTBhfZoFRa8AYxu
PwtJPaZNrCFjtm3zJKAuJGJleyIDasw8QP2+oSOhZClWmiSg8uGa0piiBHt9Fp3s
nwWgIvS8bYXAMSTHg0lej0bhmyiD+IuA2l1rRXb9q8acC9zkghdtvSjvKlF50oVl
IXW0wK3NKjHI4hkV07lyJeGPaYjUwrwDSpCLHcUNXcLR1Q2ishzLuGRdxeE4cYcd
UuISX3NvbjcqMqZ2lnm+KeyFTs+YcfPLE5+/YLwCYyFa60l8r2UAqdpL4FUlfSLd
dDAf1fepu7oeT+ZUaqKkGr1LL3sN1oJZ+zNpCyZHi34J6qN1XmbYOaZLEXyKwRUI
MdwFVlYDCJLcas8mmgw0CIbwRn9BNmBplAsnCX4h60Y0h18kZBQmydpnLtY7SLRX
1Z9yFB5yz33hEn2snJtY93aqaeVv81fMgSGBgQfbMc3tYsUs91pVVPagZW0uNQfi
HCdpLmqy9jexLV82ht6d4hRkH45m5WppBAA5ZB7KtrLgDSNBxJ0OdNcoc1nVW7iB
1eJrWD/t614qS9ju6hZJL9FXTvkFyICyX+R8LZy8Wi4niyW/f459UMqitvaDjVvr
RYpXk9VW96dWx8RT4bP4qzHl1Pd7l6Tq1hAI5vLzBw91Ao6aBZJj2/8rpCdo6Sr9
bOgeer8PQor6PpdoHtyBx8dHoJ+CNq61PWbVUrXEUY7dDKYhetqhLqXBmVkX1Ijp
smqEObhbGB5yBpyvfCLvX4wP4L8S2CLtpu+BQvDw4XceW/Z67Cp7p5qQku67SouE
ztCV8eASBmo+8QOOLxU2oDS5ISdKTMNEVJhzjSO1EHxLCynJYlPNZ9A1ZN3xr+D1
v4U0UTk6UAGydevtBJ2iaacndzRFR1Rd045dnk0HD02Kxq32M55bRZ54vZWUhwGu
R2DRq/s3G7/sjZ+W8bBogQOBgZCZBTamSAScpu6Gkk8yvo86/jHkXNLYlzrHh2LG
kEm6nu1BwdvMbswm2ff50hJ10SK6Ua9Zz+00DSHXviYNWyPOu6PNSe3htqOT2nSn
9xYzFHCMEdOrw+8R3yVJmySjYOsXMNOnQOHeYv8XeYJt/wKtzslyyxfvqhbWrkFz
TgTd5QMooENfIdbp1kUZshzc9i0/HLTA+U+4w3a/AzTMPAgazSnVHUE/LDXKXZfX
MXiQJYcwfrto4VV4HHjSjFXlZUBL7nmDk5PsTGLLX+/VCO8XpfjXMng3gpt0YrBs
xMEimyREl28948VPobuwRnmHQv81yc3QTQhdq7Xc7tCkwxmpJzDCKQ1jplQABSk/
N0HxtdIPdpANU8Q7YYdZ1mj3rkTXO98WaSVvzTGjR8KcAxd3e+/OAPcGfxgJSoIi
yy1II+NzG/fgtr2E8nsWFKOUlSHWW8mxXlq109Mv4oVSPoIDXGQXIqPP8stbUG7C
r+kRIZOJBS5rlZQTg0QDCRqHRCuiYAoq5kSI3CjVuKQbXcp4jcWW4D3fssEHnVIF
5asdCkYWMeHRAt6TH2mmQpI2UmJZNzpqBQqSiXXZ3xsaCLyy1YneYgS2kVryHQvo
ssdOPOSLUQ8S4mHPy+f4Ulctla4vdtjy1oLmHUTg5b/FTe3Jis00Nq3PWgWPGCa5
YhA6jptHYKLGZHBrh0dIn7GHug3qhOsweeUi/zcZZB5RL9g6Nuyh99RPI3Yicpuo
002wZr02KwYK0xTnbrDK5MUeSFrVTrSc9dm2n7lgNkPC+QwID7GifQ7cBii2q4Mf
6KcVHN86a+JwGAqQ4BMaSFJJV/x0fxUes5V0Cn41pkrdJhxrPOgUcrbtuNmkmNBn
gbY8f/7ru6U8KAjqXJtmm8iCIGi3j4dq4BVf4UzZCcNLFrIueeGGpJy4ETWtMpWh
+4X4s4F8bmdcUn+uKovw1+ZFAGeicrbNycBwSI5egR+ISPdM55sPwNxACkRdT4iX
7WrVRFTw3uYKqVlHjWcQWd3luf9nOi2rkwtzNHPWLtiOL4d+CF0OtXRRepr8yznw
gdsmBYycvVY2yKRQXHkLlEOcOg/iInYbh53xQO6uZFjoCTWUd7no5uljTLaRQDWi
LXOMjQrUvIgiWZ6iNj3PUlYOz8D0uYWkXxXS7AH9fhUog3aRgWM3sO/h/fVuqKx1
Xz0QcvSjEI8P2yI2lzudFI4TlZkHaUinkkzfTPj686PyusbjGviDVBU882EDF6vE
Rq/gJ5hhx6ljlLZMYscdDPzw1odPfy5esqK1KKxsQw7LNZvmoak+VItIyRHImrqI
eT+u2079XvBktFw64aWUBubv4RlYj7dNc4E3VPQ9M6mqlctvgYu8F5x4V4cqkS6B
Epbf0YQgu3C2dTXXEycTg4Ow5en98wHN4YUCeQJwcSP4hN0KD0OSN0rxBHWU1QV4
2WiK+aql9HMuMaLYhQJBb+SLZd/3jmMTWsBB2GK6HlPARLdC7ArAgi+BSJ79X2+U
n3zS2Ngz5A6LoJlKySOzLUvAX5O3JX/qKvcd2p1ukmo4pfbidhv7vgLuQ5VYAoZi
OJQv3LgI5RvejPDtgHdthS1n1yNqbCTYEOoKzgxWC5++pVtQvDE2jr2uwAuuHktZ
TH41QGGMHGIXfD60SKAg50xn3PBtGqihY8BfFzjNCYn5yx2MgpylSa4WeNuXePOB
TKPIeM62EmPCMYp3sf4W981S4ea/d61VK/V5sQtgi12StEm1c50sDU4SsBF0i/JD
yKuC0z1+zP1QpokBKxPo4CxEIy9X9PeWrpcEy7UYlpFXsvqs+VHKl9+d7+EURNf1
jgln64nwsciQtLdn8yvO32R7zZvxv6RJJk1ut+V3NlL2MptZzErZ5hJU+21JfdUR
RbhiZzQ4NIj+JDeEnzJL3ArodTg+TjVTkxMlA6p/r43crpb+SGZ2Dv/9V+Knwn0Q
z8q5J7S2QwwqnrL6yOfbH4XAYQIsapxIU1NLfJo2H0Yf0ZmSJPhu0qImfe4WjLk3
4+zy2SDBVmQGPKSU1axs83xgQZYPQUr5rPhnkrbEFe9RCBvVuE6U/8vYxH4z11jf
XM6xRVittAfOq1AiBqVwrug+Yy/QfsLRFpgyKyjS2cO3uFyU8hklS1VzenzcA+0F
lAOxnMe/RnMyY4z7QibcC/YzAID/1lNtEOjZKHE1mZWsKZLj2tsQP+eQNjQbQN5H
H7M7DXPIfI3BTfh9WnhqZVXiWcrHtqFX8XojCSTK073+Mc6Xt2IVeJdG8YKem0ih
hj4bAw6K//CciqWY+LPEcpvLQv2GEhJuDFm9YwTz332iKODn1F8/ohcXR56Hofq1
FClELOu/trCjwF8zS4VY1yK6QdUHvNV35H1hTRV6mFKTooYnd7KMtQVcHrnK5k44
dTxoI3IDWwV1o4zVt7eUomy+yQRha++7sBOMWrtLyFfKvSI+LjaSvDTVd8yqtX7q
QyVZbC6Rb6iyGiR8QgsfDH4wmF+PyPsinLQR8+0JN1OLwQN8zvhZT/kVTVtFYoNg
Z+te13HA3agyacM8BOiQvwnvPfX9v/172pAxnSzcgBr5nlyDJjpyqtzRWIAwG5tD
YZto+rLM1joGeKPvxDL7pr4GDqSp6ihSE25slq4y3pAbGvzCshoaH4gIboFOssfb
PIlYHwpx2+6V6gZS3qvjEvBmN09iTnFh7HeIu4XffepRCNhayf3szH1agmoRuCrF
cjbFy7u4gCJb3EGi98tvXzx3tp09GGWpoVpDhNThk9Qn2yuMxV3/eGduKmZuZgix
+l4boZDGZ0MuztSb38d6IP2TXy6AaeyHLh9ymgDMihAqZ3kmq6QOxvL/68YqztSa
brbrKqnRY1afsdNYgbEUPPu67TbN5Wda0kIOoo53XSR6HnBuUqPTRFMc4gO1bk+8
cRdACAsJnBdri5G7sKohgXLakvwawGL7JyR08NepNEgBuBNECKq0rvMhCpLBmgUy
mSQBz9qUUVYtRXo5Y1pel8pRtot9BHOaX1HPuFLMMVxstKQjFiXYdPNu5r68VNtf
Sc9i0g5CiPk00g+MaNKzO0oR8uabPbDs98rVfBgxcfOfjnBtmmHWX70JGjuoKRVt
csUMIZSQ55c/BlKkLXlgMqWnctXqwJZkVHvtVUJ0XeSKlDUvHhldKmZyqEFgFn6l
x6998YVPOfNH2MkLzjn+OYIfPLj0NskSoCmw4IIPH3DDEFbrR7CJHPh9+25wNCm6
C7JzG8fSDyuv2pzUiFvt1rNb5gUr+q6MccmCY5C6ZKsId39dGT+myEMFIk74DJDI
Q9FBx9JKpLCZ+So6XoMP1qjmS1aaZ/khtgBoCqJMnoYznkKVR75wVCDrjfRUy0BO
ddWqym4ONtIXVzImQszTidUj7ljtVXmz1TwqydDp25+ZlBh5qDrdXpuFo3zrAaPr
T+NaWYZvGN6Rbbec7KJN6NJ7vWT4KmN9kt9ttCRxLeYrV2Y156K+GADCUFym0q/d
req8NI51jcu8cw87ZR4IKxW2xr5hAAd6jhhVRIo5RvcndTUSv5KZ7N/rvg8C6gGK
+Q1AuXiTAn8BeDvEbQv7Xr5ow/w1LX6S3h72LyTQycGm+VwK35zH2pRKsqr75zko
4e6xLO9GEnF+pMny2HM11arL7TvKt5gCUXSr+nPZx6xqL5VzHWBpaQJvu/joqY1L
zOIOUo3cHsDJd86CvAuhYIj3blt5B0M4tdoV91T3A1JgWfSaDH6YS9ie0U4y8IFz
6gk0kzvFef+nQ9h1aFwIiAa98fPd4c3o+qLgBUtoauCu+bK5txVVX9SweQHahQ3p
lANUogjMXV6T28qGOT5h20bveBOagpxuPPdJ+b8xant1Wg0thTKjhEAq9npH4AC3
LGy2s+CdmGmeBr25wSJMCVZzJJiBeEyfdDUFwN7Tlu7QmkuCss80joAjCZnFamS/
MdQfSEVrTrjmiGeaIN4lOaUgEBlFCzj7GQXC7VweqR6jq3+N3TShnoydA0knFBV5
ekvugsHP3mDQay9nSd4DFVSbKsq6OxLLgSTn6ITY/Bq3bHmWZy7e2NIX/7WT+93j
3isbk1HySdhnLaYitL9jzaO5okoykkfA6QrLXdjb46SHYZhDZhBgy/X/3uJbX6ae
2oLl7ud+tCIZCtKuoJEYSfqPZ0Zw6VI4S6xfmkhJroMIhpB1CEl1eKtxKYzsxLQH
/R7F3FwFIOzUKMwqurBm7FUyKuzdbK4l8IMybzU85pbILgjWvIXypd3C3tDMJB4U
W1tYgBNePz339wqLFKwNMw8G0TMXOc/zvuMiT51ni4K/hpvd86nq0RbMeG4hpUxt
2nWhX/PLU6KiKWNBy3zhDF43efSfqc3RNW9cdBqXFUHo91mykcgmWkkU8WvQeAYG
6JzY9deN7GO792C92UykEZEhbdDY0SS0qQ5IPeegeYcfx3PNlQ52sXfzJ8kRKj0s
WLfrkIjqTeVDkoDbi5BDx3n7d2IxYXcgtLsB2JrQ+UKZIH7t6QqPp5zgJ1nesezh
5swMEHU5zslN+snkBdSCpraWoYx9xfSnGjDZDl4RgRJM3o7PuoMEt1zZzleBZM2D
wHbKaoLgTyNqaxmt1bhZIg8f4b3XdVQ+ka6frULPzyRyP2/ElsscDlscjD+pHs/5
eHvuPx4u+AWX9Ho0SZQ+kipLsXTXZS6dsOo6X/ixoPRk8OtEXHxve7A/tijxHyw9
hac4N+8xuIs9MmwBVHXr7jZdJ+r9OE80xxBIRxE/BkHeDAfsfQT7avZpLfW0XVvV
HQRPcgTgjSpNnq004c7PMYiLSy7kKL7PBEHwlEBDNMxkSpb5yOKtb35lLBnNc83Q
+GR8MnQVItmYVWEcrSqN2rxHDD75cIfs5PoOqGdHSQc5n7aF7hk38ifjhPW+DO8J
AFUeYB03WbXiw9m8DcjYLF14vCUjM8iWZE7UTEdYh+1SIbQOZNmfg0P3ve/4hXmK
hGQQvni5xRNTLOvl65YLQDR51Lh3HyCJQcjVcKQyk02+88mvbgtt1xFpC9uzUdGN
ByLAbA9bE8zHpsvge+DrwxTStLmQ7E5f5/Q2+MqgUD84NAxfP4jFs4+HeYO3kExy
qmatWnjaamNCpaEz8UstMwLYlz0bKewCESqKUP2k8xp21Z0wV+l+7WLgSFdvVqIt
uNZkoOr56Mwe6hMo0OU9zm9H097J9DPVTbx2rmXbntOobRQCxquHBoJvAei+7XhJ
j2vmLMkQ47P/JqFVc0kBlb3F9O0SZlvBVL9Jv6jtgsRmbUGpakvf/OxRCepEwn7B
WpUI3qmMnuY1XT9OhlT3FGbRyVb3zRSmkpW8SbY1EaAMpYkH1LQK6fUTLV2duLf3
ENIbv9ViP7ZD8pSspSmvgjA6DXMK4stFC9krix6u4BVmuDBoxSn4aLRyBSpHhoPe
C7zG+VTIrYPFUkQIqcdZxbt9IjBQUiMUmtqadS/izJO1Ke+qF0+N9x99tch56La2
XmMjWU2gPEbwhMQIpLfg/3h9xdmrsROj1wGu0/ditrUglWwa37NEHup63jBavGO/
lrf7wpkLKgjcLlNpRFH04K1UTlYZiIPeY2mGlz5vJh+i656cmbetn0J20tZD6RT/
Oj2rD863Hzj3lJco8RomIzJMa8/eUh9+DgSZA6/dUJ7/b45C9jAWXJzRpTAb1V8W
HkMKA7We2hwKJVuylPMg28z5dOW4R7q++4yZiM51YhfEX4hANTxH8wfoW1pptD8W
zK9JIwyb6LAj5L9ddVLf/nqosqpOnDwe/n4etUuHA/gm6/Ov6/Ap3J0U+j2dVwW0
YggBwGeQP4sPexSYOGrppLcTkzUvzfueVYi6IHiv/yad5z/OBaEKHQv6/AU0XZgw
SC5MMMxdXj13hweH2C/b0198nfDcs4y5LIwxM6BOGsZDi8qXBOFrw0qk/tlMlaLZ
3xb+1WN0CI8c6SZI/AZjChLfE/oCktjxgZ1/OORz2V/HfvR2uX1yiF73biWLtYKX
oTTpr9VVZDK6czhUcerTJWLEykMmbGDmsh1nGoLB3bt083q1G9qWk8zCPxTQvDME
iqAh7ti4Dw9nm7lZMGSlGLhEaAIEzenYDeP4hPzoMu2KsQdDCuXTu61UfPjpYDbO
1nJubc9Dx5w7r8HDKoLqXTIBR8hvXLb503g8wg84jJNkEQsGLUQjqNjh2oIXW8Ui
pb/EF0QcS9BsiABtWZmGp/M8aiY/D6wu0lTGrMypU8lO6Cb+2uuHOkr/FBZSsXDB
5NLQguI8BBhuNy7cSsMuOBGIySq503G3lnxc7M8SDrUa5cyIsWJ/14t5z3AgD0aL
KM5ntWnNutxbN7lxHxexN/oEqzrJw3Cb//qM9s3nhoIIkQA30FIiyu58D2ZdTIGw
T9qIENmVm/N4m/2OUPQmh5lZZCTp5GyWQa9ccFj1djwFC0SgHhwiTaFT3WelynVM
f51DF66xP+BqmumR2ClEoR8E3hgqpct3qoI3SMcxUsX20i2QnQA/vyx06NBEPd0/
nc9UyfMXwY7YBnwSfFZTJwCoOZYn3PidDdkju2r6yFqXTcvvxdJbWwOC5vy7Y/vH
16mLhEuTBL/UlqA9NeNe1B/gD1B0sJP0r/o+V15jqXeG8fzj2QcVi8JNVZUT/JXw
70O+PLBF6rWcegLytEEZHmZYV019Y8kO6N6hVjarH83aIYI6HoMkLSBAfKWJ1s+b
F0vO+ILGyKxg93rpXuoo3+qm8SZLIl598ameQgEQM6VD5mpimhFjp3oRqwrVZCyC
Ly3nDKAI2jValTfPrr1rkUXczt0+JRvs9mDm1bGzxnI2j0OaYzl1rybADUEgz6lh
+vMPnNwKFx1VIMWLu/GQrcwC7PaxZeMNwdeodA0PDg3cdWFOqfmIYGdS04ZYHr0i
8grcLqBwSVCoyGTBkvtLVgDmgV/PpEWXV3g+tpbY8ps2w/IoP8CilEVNnYAr4ZqH
Rx+JsqJqiVEE64JN2K/BGqWCmKoyorGTYJM9lpofLaEDZizwjEOEgRQ8LUW8BLAk
hdeJiT31mNwDHl2B3mL7lobaDzpDejcAoD/e0nKPTVBQ7WtIx1G8jAPLFfSipLbj
1yWBxOhiv+2AeZgJL7E+5J5WHbqaCLYVHfSM79LLKDvasqg8Kl2Vn80AbunIpPcF
wfPJiTUk5z6IzGDuWfywKCYeVTZj30h9xfFpNZfx1mKMhH73mUr/gQfLcVO28BZw
NOZ/ChxJGePBuCmc5TO7cjjqkRns9BWlDB78UpOtfIi6GSctP5LlWvIGM5OzgpTm
ycq4KgQAeVsuU8DoOiAfKUT7xC52Gkh/DQ6UU1kJwX3RyRWoqYn4wmMFXdvlbVGg
SOS3dUUAPqajaco2Vu6YXsU1xvWRXEi0Do4LicI8BFx8Qe9KucyJrsBRDtZlwiN3
EmPv927uB9W4Ou13BtYfO1adv2R9dCGwVT18cCuKqxvGBRjel2nfegnYUrQPnSdt
f1rTb/cAymDhXN+IBDTc12sMftEpF0SB7B8KLA7yMwNG8aQbG+242mmEuJltkiIE
AL6MRYIrmSIq9zJ60hzSf1RWX2XbrUOxrTzZPcC7zvovwKReZH0MA25hHEZtz2ac
b0OlsLEpYrb4Vi+0fBf0l/tux+F7If5jYMfzdBTyZh7fMg90VR6Q4Jqgr1TqWmQT
v3ZF5ZaHq3ivdFnHWBJdy44jwwyuZNdjx70c3qvvwaXYk95vT0ZWqTvt9mAh2NbC
SepcFu33qcS9WdEUKIjLSGWaKwPTs/qZKTqYprBUwSK1jRHRN7yu9bb1ZYgckw6T
mIIGQLoX3dGuGVik61n7OFjL6znlANKXJIg+MmevXz2jd34PivgbBWaPoQCGSXUK
YmMJ7DztF67z5viAPOIWe3scOXZszhI4DO0UGZAPVyLyLGX5FJm6Xl7YW8gSmr5p
knaCLg4ta3FZsN9D4ce6sjEReV22eZRY5O7+BUAxZt6GQRK5VfK77cGMn+TnJxxc
D8L7Ed4SDnsczZObmAD3SG5YDEKxLyz7wAVr6qgwGVgw+lUlvfPMPZbwN1m9dUcu
Gg/JsWhuR+6hl6Ahd+vR1NoX0FCXaJIj0z4jyPvLw1AIqhYQCJAWwvWCwpAVUbmt
jpo4dflVDnfelPecIndaF1WUUDo6rhM249M/P7UpZGCe4Cytq/hUchMMaJG6Jk1d
5JYFWrtTUZuvhd1s6Rbi/PryPYF96xHHN0QhvgGBNqaaYN8A5fS+TJ7QTCVhXsDx
V0gOYprTykbJwZHUWIbNpngarVBVYCse19tcp3BxDtZuNhuIiUGLB3jvwDORQWki
TTqCfq3hIPaoXsAJz7kce5DE7k2M6F8G35dWhV+rPgyin3gPLYUqALwCl/3Vnqno
QKNJoF889aBQGzmQpMPrGAMQ/YNjS+T2oh0ZjuWY0CB/+dMrYCpACGqmLsSBKLGK
oqwwpcdJ/w3ThEL/mEsJnbQpihx2vifYoqOtfwdM+U8NpE2hPln4XYO0kb4mj69a
bkDAXrUcsVQzfUYMM+gHz78bVeVNv1snDwZumnTJopsbZZiOGR63j4NncOKv5zcq
sjbjiJPetaha99m7gB8KLqE8vm+qj2zQE+47v6NQagLN1kIX6TwVVgbnT21iQqq1
Zgepp8Av4XmP5my4DV9lAOym/Xi1ypzgI3Vr3DVQiheaGyTySJkxL0W7D6rJdQdI
56Vv/SUCZX5wCz5yOA7ApiTTqpXDuGJMjOqG7COXkLttE1RRRncp6W3GyIQx72nr
u8fCtHpjFVVCGVbSxmZPMdMJx+1xx0OXjTkVGRe9VxA9H/tg08i8Liiupv22lrsc
zp/E7YWRGOB8XKoZ/+BFlsZXvgMT7fiTbdGnLBj4imCyQJwpV/6zLLCO0FJ6zFeA
3Ca5c3CU/evTm90Kr+9MY8PhXnRgPv1NDiV5ydE+PmlNlzq3P4DSXU6+yO+gn0Sy
qfPyW83cYwnFWzrM7RfvtpqKSvy1Xj80yj5skHpwTIl61ZOOXYnoOsrnII71nnjc
JJE2BEjUwfMbWQn6Sq2BVCuPfZqdLLkZh+VLRcC251L+r714GeXYnQECsoJArqmY
Sh/W0MFNtA1RQdzsSNq5LoDJlRoM1ZyQiW9MJLA5PQmdonEYSTZSsVKnyJ7X7rPz
B1WePZM7Ohruhz7cCHU8YhzhRjHAUnJAxcMHjoNgZSkuVFn/id+fgqYWoswPRkUF
O6Nq8JQsa7frpXetr7/GyeSDe2pXVYV9gFZUH06tn9+lKbMvkbLGlC2x1PEMePTe
WUak1bZjri7Bd1uc4KpqnCC6Bkp9RXYZFCMuFTxklD5lF49KC7xXz6d5q28SVtg1
GI53upu+VY8ZNo58T+1hPVFMDqSdEQzPfNRQLBjDNu1MPbSfJ/gJ0hUbfFJA55dd
e9I+HeMR6aE86eQUuOzqMi5AxomO+JohSxHViyIBiZeVGpulYdhGSLHR7/TI0qr+
PqAeFlViEm+zv2qATSDbbfHSBabJisMsBcR1ZRz+ua//5XGjhPmvgpO4Ni0c6frw
lQdYueLEE8lzN3AD8m9nHncYW4acT0w8pXRukxKJIaHXcf0H9SQuzTuGTDC0RZDw
SOaTn/yFxNcgXUs6SdHyF+ccA6BxJt1ebArrPYzvYBUd+mG0pt5aQorPSS62Y/pO
8uqVjE1bNEwfFkAuS8LY3xDxpBAdcG5rXCTpSbd98vJ31Sm1SMhxF1Fcs8E92P5c
5xsLvwrRrETwT916x2lG+sdtenb52YuE8K4Ik/jK1UAbOGJ+GJIj2y7DblNny9Q6
51nqeT8O1q1pC4LkwpqTp9hw7HZzeBjvhkINjzKZrYXMG8HPXW1W2vgHRNOQhWsN
x3gflofWfwVtEIlrx/GyWmYNb9eo8e54JpSanIlDrO38NBZ1FxcP1PHh+rjRXBpY
KcvtBOqw+qc7ChTQQYGZ60VMXi4a6aw5LLnezpHqIIxqxwR7/b3KTNSmjwIj5WS4
K53MPwr/ZTByw6rBp6Rirdq+k6QCo8Fo3FL+wL4UXzym8yodsB4fA1EXjH43PXTx
d1gLap8Bxa1DS7UyiTTh0RelaD38SX0ai55hagngVT0bVMWP6kgMR+DGFINpNSkN
Yc7p25sK4Xy0LEc9M4PeOVooPsIBM6s+vhqQxlA9r/bJ6ok8653VWkUay8WF9kIs
Ea5fHoI24sIUs2dxKkRoHZmh7Kq6Xfx7lZABMMGpt3jvoAFLVB3gHT6LuweIrsKd
kUyW8YXQ35m5LYgJnH+xoJBoI4jN3QXndT8+G/rb9SChvN8cfEgZ/fhsRq/wE2tS
FwqsWyBidOU2bB42Z5jssFiNQ+le4EAEAFGgSZ+UBXJbEXgMygSFuYNPcPL0TZCW
DuYuaxzw0bUbCQEax1kZk1kkstlRuS3ZQNhXjZUWCzEW9CYP3fQVtzoaLdZC5ZDy
imhP2p+TgTrVbPhb49/V/AhBPbY4eLKkMuLuhkJDyurmaRr3por63AZlsk75xvLV
tlIyiDjJVDOSnEcnkf1Mr9hdvEpDfGOy6g8rY5HHOtaoz4m/jdyUbt6/p8TgA1d+
86efs7Ec60Uni0l9IJXT1R23Q+KQO5xjCrtgQi598fzaR5PDhZAfUB3YgXDHV7rY
0r+IMWSYX2hWTm4UKwaAUQV4O9Gc5QYLPvBjGzfeHs+8pn7PvIInkxl1ISTco9l6
yhQl9ntEPE8fSCqQjiz5Iu4aqX7PKNs0PnhRwFHaP+aJHupvyUxs6ZW1xn3WZjiq
mR2m+Yc4mnPX23J+gtfj+b5dU9dWShfPUzeRpXJqRaS79MxTAmqGaFVnr7HACeIO
RsC25rpXrrtgejIR9B40Z9tH3w4sf+LoBeVwdGeqCYmro+q9vnt9tkpn5HjCiEMv
da+3oZz/MVmyV7MsauL79U/M76ljVcoWEmwuuyQ7RfywPEfKdeNWqgEsBlvWlZc3
7AAgYG4k89CTxM95eG6ecJqg+WHeuj6Ypu44WErWMJftci/B/43JHLNn808ZtT4B
erZpkZOHZSRXID/vMUvFyACVsrrX/jAVOahHoUh+c4mb6mKZNgUeFzxUveOg61bq
i0xj0bZq67s8lwZeslPuX4tzUdkP93sA9n6bD+1wuV8f8dRIT1x/MjWk8NkN4DmH
UTsZejF1YfKepr4o06RIMwvq7Ef3ft2wiaxFCwcu6HLqm5etBMBhWUTjYJxNkyK0
r+bBmkYaoD7cnXYXCt/aRu4U4X545NDAnR49LkZDDI5cqSCQbbZWw9e8mzkWZIT4
0lyEw/7kc5iIuiNHsetwVoTbCoiJdAbiQhHASCnb7NRdPIOCf0VC4VU2cyyp+eZS
T+Tli4Aed/3nmQOakyx/dzmqBPMu/qqF0EE6ucdRVqBNKPSUIg1FA/sCfx2clMbH
oNARAnJx6PPlJ+VmfHV9Joa0X+xePQZZDQCU8CYG8wFt/2oX8IK9gej/L4UoBuC5
/uYKzfavN0hVMTj3cDCTntVHiCt/6BuBbT+WBc+kXZW7A6zs3u5EptV/Ehr9ieUR
rJ02oiHI5vROu7AAgREvWMpfVaWF5EzYzpAqUS3Hy+lANsf0S+Vu9HCrRCsCQdOV
mjZ7Z1syd7zWpu3o4+ia1+9R1gDxasPwFDDzEkTWJyFOMPlNomIOuBO4Qc6J0jSi
Bf7eUKcHNCY2B0+eG9xJaePiERNZsMFe/jNVFZWELcJ7VZbcOwXV0HdCxai0Xi/z
IWBiLtU+CMyJGX6hd/cmJS9i9qMcN6/0cKBkXjuNLSA+DlCobPmRxZsNKr2mKzV+
RqgnMNVWEg++eNK953RulC7T3eJpKBnwoCg5AG66rVVPXg1OZw0qD/kODWRSu3PO
o6aHnxqxDPioiMgUO36vDW6Z+Ed5cFtJ2XQYR42JFlbGg/F7mmlLH9wEOauiVndL
trl/fG6AMW5kaCNGTuleUoaujVcZSD0w3uDUgt+dxtC6l1uDH9eHTMeZvcEVvgQF
MuCxPCGWWvQi7DK0PWwP3dGD0h4pW8jOhKvibTQMu32oZM/03/NhViHW+XgnoPed
j2TD1Vf46K/OfUm6WVzRHWjHgvJ5ObfdJS4SALfrnfrk7TQEC0LTDS0rftFtxmH/
kWv6PHGw2mzua0VdcyFzhI/eXmEsOeCIto0qm0eGhE+gmYHlJd7YLCxmgT3yfBfm
BE4JS79bIpgsVfZQamBg3B0WgQ4PqEw21fiSZL5ewbQQ1zDB4gBkZ/cZshc99bNv
kYF7OuWL3BgLUbQCwFL4nx/j/jr3fHx6OYo4yS+IB3+RlGmBnyArPv9LRP1N2sV2
9fo+qDAFVhxO6GvmtKbJztvDxD8JSdbR3bp9qlU5qFiAws3dAkbgn0qih06gKwux
2NBpFO1UatbBJMc1bzwv+sfuZG8InWEjVbadoemTMqD4r6eo31MwwPLU4VHuJCuk
gzqbca4MkONQR+J48o18OXGNtwgM0ApmR/mSPrpCSy1MTdKNL3Pv410Y3Xkg/hJ2
+gF6GOL6ZbPPVQUpX4vR2LEE8wLyRNCxgxAXRnPg3Bc2ZUgC120Kkok43hmaU0RE
GSHnu6bLVOc4bYI9/HiJfF/QKbcL8/VOjqwCAxUmY9Qcn7b6wvyPiZJQ3gLOLDxc
ijHYdeU17Qz8ecKZc/zPlh0IN4Bh6O7yfRWJ1rHzwsA+1Cq+QddQMqQZSCVIlMRa
tizBwf0AerfMrcJajrkThBCD2ClkytM6zHMfGt1CoAaKgXF1HVc4CR/w5A8Xr7ki
7UbW9SvRt2YS7pe9UDO9vaD0NDEGjVae9ouJyJavTROBgJixQmGigQUSYCzZQchh
ANZuPGwcuKzsOSs4nEq40W0D+5GtOxSqEkftt7vnyZ7hINrpEs/c1EQKsjhX1DN8
zvs1+CJOMBjMtqBkAzC/rasjyIOKS5YCOlcxBtxEQXeD5b9qkwMrpq4Pzj/ri0G0
QAn1VWwdLUZ9iMHcpFe2GaiIC+7ri8eMfaK0pMokc8u/Dirasw6XtJO9Bz8tMTpQ
JsXZKr0OsfcRT6kVyIrp4VWPPRrukloCmnKphbCTa2MdzoaFU88Effldr4VWIDp1
iKtqrB+IubG+WOj0JwxUOrSnnGBtKkITJxPxV2ujNp1YrKpyIoEwpc7iWDbu3UDx
lsAoa2ANGIWiC/4Qcfe6wLOlm81R768MleFjPLMWpvDwCNxXZYbmkvG2G4wAsIHw
tA9ukcnOpLQkhj2QAeSzltXbaWbE/q3gJY8M2Gk5/jK85fKKZWIF6neJyKvZZLqS
RrTPrxIDQ/lWqZ6bZTpf8TaoOOrIZZk35eL5NJUwHvBnUYizMchT+IoFV8FjiK/u
9KQiBpbsknjhiRgVVY8LaykqBhKoyTY8u+D5MUKSLGZAk2uT5VZbdoUpXCUpTWgE
D2NysGgXCSxWmFN9StO8I/Gd5A92d8jQan/iUNH3FqTfwlEqlNixVXiYmlraa/5S
mY9tLWDzqi4yqgWtGGasbeZWwUxWT5S7EGHlpCSxqF1LpsGb+j/inDI7TGqqfyvS
ce431/NNZjwzaRa/2eHNEcJCFCr+s2S7tvthAbvDl6Ca93HjFgwjaOFJ+k+n5VWF
Lif+GSVgme+nrPijAiwdI0L6YAp3CxJmYoVJTo5r8ZoZsrnAtJBY5K8/cjtBRML3
+ngYtreY4qlCzpoHs1N/N/MKBic5WLI/C4G+L19opBkmysQVW6mqKaVSossWMcU5
kiBmcjj3Yxg83RgaKafHAZI3KxBNXXSWm7vPDT16416o6L5d3KS/v4ilsu0O5TJ6
5l/LQjehqd39yhJJXA3XPf3N947e9kwMaQ3+WWMO7+mvFbhHWGT/pikv/BI+ax+z
Yuaj+c9LrYoP7YhiXFDkLnlHC/sb3Q4uea8YeU5lJdu61FUtgb216KU5+vCuUMc4
20Bevf7acmE6VmK2wxTyq/mTIIEDgtP3ImU5NbSNYz6zw4YhIEdQ5lvyUDFlIC7n
GONgcx4r+Y8Wqg4MagKDfPxDGTu8rTXCBo+oaK+8OtT3I0nTflYLmtGw+yLLyK0/
Swer5PKwYmZg8Q1F7wFX1fGBUIGDj4F2cif8Lsd/ac78d3P/kupgjooJcfy+RKkw
HIQeaZbfi5PDm3JAEBJAbRj7zNyww5kNxDv7Sc3Lrvazp448D9U/9pe3FnNl5aEW
VBVjBuPnNcCrkxSheQoORKStO9vr+ROxl83YLWmCKKkDmAVtpLdAB441m01ccd/t
JQ++UAvkXASGMRzQq/q1D+SrwnmT7lSfpoX+kayNxgtOF4qzutTPjfx1Vfesj3e7
7MhgAZMlpJvp/LzWBKxTuarrejXm4FlUrrQvIVpTTnGeLpBt/ovEWH+4Y8d+mrBx
w/lJKpS2F8O+iQCcpRTgKA6/Nz2eVy37RkQFPAqAP5x1H/N7tQneLQdl3gz6aOuV
69TspS8OWV5dhprjgukUqiE5183DwdOkmqSQuqr7vb/S5Helv4FnbSORxTBAh6X8
d0z9FI6jDUYxbQFPR5lg3+C3FotYKKTuixa+a388wbsULbpeaCC4sOpZWLxGppER
av76f09gPb8h3zd6MG7NAwM8AUjcmmsS4CdBc0bT3Two8dOl7hjDBLCO8Fq5i7Nd
eJ8qOUFscyeuNGLUNY+igrZnkf8wK3fREcEsfXjMHeuBD5sFYiTLZFx3HqJLW+UE
9IZyhiDBpFh4vart8c8hkp5Lcjt9w1k72f+yk4y7cXubQVPdkQIO9nSmw5wq3tFw
mEUtBwGzJM7vrvVpG/jfYyr9UTrbDK1nz/NuTacRCj857DKY7H2uM6BaEXPVC4E7
8qiL2agbG0JMeqAqJZJzG0ZmFazlELIkH3f7LEZujy3wTmeKc8D6WLviCn7CZ6OD
dkugNpFVNUpIQJQn81yGAgwr/XJrdaHhe8IbMGkqHErYQ8FclwZvttXqKePsLTyp
JamzwYgq9bKu7fItQKPMFSl3tJBw7RITO2u6DL/tCLu/1DRMo74rBqSOT8DYdvF/
Butjv8vPysbU+ZC4puKixGNTv4DhZLT5oqHwAQlXQtHdObApkwm0c714vSuIvoVr
AfIpg0jETYG295vmF/FZ8D4PoxSCBEkW1JjGNPlQpVjZmbgEkxCPdrEsff3WIj8i
CQyY0bSBCo5wFYGKd8sxhPJuYLK939qL5sUqqu79O2Y4/fcnTjNEjSGX/XDbhsZ9
N8lTfP2n708IrvLTsSNlW6Sf85k0yd3h+Ngd6q7AuKakQYVZPBudAnyrXwngOHw4
fm4lp00SthTc8+t6eOOQux4furyrD6U+z6RV6u2D05L21Av1uYqVxmx4qh4nX1Co
0tDKhU9fXJMnhVPJVdkK5X02SnANmLAuezzFzWOQpxhgqF8RQRfdAB6qLAFhqrxV
4VocTK9yq0z9bb3jEGpav6sghT34PSZ87ocwJBNhpbaUbPNAC/N8lPQ9UMk3xT81
OYTTWJgqQ50Y0ehFEvMA8HLW9NVMgj7Ga02uP7rwJhz/50ZKZ/L6q6RSMEOjaB0S
h/aqsWqAfwpYZi0OF7Lehd2cVgxdgPYDTzmLF0faFyyZvENK0ylvA7IG4Vu1LQEz
e1EeJGo0BU7icZMQoF8BkaO7bvlCn4kRUaTFkP/VH0mqwn39HRKEILx9xQm3PkvD
n58hpZ0CtsBnCHIMX+KBgVVelmsH7hjkjqtS8SVH8lIKtNyVFrd5Ko01xqeJnnAp
bAlWJoMHOW+swZpH/LhJ62aP9YBDKgrQSt6eHyaagSGjaFQXF53n4+lV+R3r66BH
41x/LHBhzCyCgFXEDqlrk1ZfSqhskwNh9/f28tuVB4ai7v+xOzH4nqBlVxeWaEsJ
VPkhipKUBBZQcjDoV0NgeCTZQGEEAVEtIS0QUFoIIQg2pDoc/sjYOl6QGNyaprXr
nktCsBYThuulAhCOJSLCNwqegeR7fJgNeaYntbRVrXudQRr0FujMhpZ+jCNrqkop
S4cuU8lS3bAwaWdDMX4D7FbkRhq6WkLIfruVVSojRM+fqIP1L/hXbUEKPG4AvMpB
+dl/FXWBwWxbAlzbtyEcuF7SMQERndgNTO0uhgbCSXEi2kQWaIzL46/nnlipjyb/
/3ENTWINY+TU+mAQ1sLRpJCPa4Gcta5HJpToxj+sX9OswhNANAfWeUESyMCGGVtm
ufBZ56Bgw/eBKpanzGo5++Jot+2l2CQCEe4KQtstncynZcQm8rGvHmd5QCxUyLm7
s82n6VxGJ4IlXAJ2ZcYHyaKrqtWvwkX2nZEgFPxm9bZUZuDd5nkLpp+pc2j81hYI
qXGasaHvzKOx4e84/lkgcPKVn2QXxrsPDhwQL4dgA6VqlzecE/aIQfkUKfpjQhwr
5EQhuKi7q8zRShhjjwNUdUbIRCMa0oQaB7fNR16a6hh0i1mjiCXn8WBCKYC4pPDG
HOYK7M2BycYmjYQDvQm19z/ysIMapqrofQ/spkOXNHJJqiIIgrr6/lk/47LglyAS
FzKk4g+GfmACXajDBwtj7y16PSpA+QHnForJRzWHkCc+nV0QE52GAdXWDeYukNqI
jrEozkPsMZ7eGuSh4tEi5lZstQ6Svgzc55fV/KZRpEDhQVJT3nRDzjIfi+uLCJ7z
50qLWnKios+LWu6OLq10u1FnHVK8piHGavO2mgY/CCEolJ67YvPs0dPc3PBsoHcX
3jx+UoeVRMmurAklNhSvqjH3WHZ46CDV+rs6IE6aVuy2ZhkQLFvk/v0g+F8ZZmOY
WWRtGeSyIa44UzMI2yW1m4oJYNCV8GZ5vNfiXVc7MZI4tkeW2TMGobOw3x7meDxz
zB/gpA7nTt5vXgHt8sjGUFdmoPArTxEaIx/rW5HU/XveuGB/TA6113ATYxHAF5qp
nDaGA/Ch6o/I9DK76lV+jUl9hs+KT8/JOIcHJHvZGB+JD9iobKcDDxZKSoLUsA2K
hxhw7a53euIAvu27jtX80oTnB5X6mjt3+4IrmT//OUrwSS/P74avNjIzNhlpRT7J
tU1g1N9qg0fyPysQYkPTMClSw1eujK3QC++DBPeYUzNX2eMflLHWDb7w5VIgd2KF
EqHx3Ci9ZoS9/E8LRiO9XtEHbiZ/r51amrAFWQRKOXvpoSwGerzxfuaRPj0tNRh6
9OgWvtUl3p13/Ht/djaCDBvvVgsQnpEBal34HkpRvGvr0PfcGqlYoj5KUqqaibBu
Yx1TqMe30GCODU64jDyhsRgF1AE4lcXOJRASzl4QuT+6yNPNVvQaSVeLDlBFIKe5
Y0zGT1LwYOrenh+4uBy327YdxvRAsTcQdNrNAQB1Vh5ecfAu4uNsiwsbmOYI17y6
HJobdsaAiVXDQD4xzPX+abOVqe2LSF1PMInbRc+NqOPDeaaf+1ktfiMFv/n6OB9R
F/VQDoUayNyymIvQWZpFhB39oTbWuTkIsNDwhyA2lgSMUNu/ocMiTohWZHKwJew4
DLKb65h3nCCiwYV54IMVRf+z2EzJrcRXOYGlaxgl1oOlRBcwqEXedoHkyhp/vPh7
rRVtxcVZBjhA8QPNn+YMej4ZC8/+cb/veUELrnOcnRXekFYqvABiMmcC5K19GM20
IE+VURUSUE6gydH5X05tHGvSjx616BA7t9Z8Fz9sTmG+7zFrmAogRRmQ+MpD626f
MeZo5S6DEXYWsQoi6w1kyaVOuD56M6xKd9/oKPDLaip+6ZLZbzV3AhjynD0kAc9O
TnMqHPpNst4DcVuL1YQ+6DZbRowmiwQyeWOQoOGnh6JP+AqOYgt9cvWPYHruZw++
4RXIwq4ifuRy8iY1OVW6CdPgGDttsvE8dFcZ91ZwwvRRwarHM83XXTyQdNlZYpE3
3UiDc2oWyK6vIMorRKOs5zcgxR+0xvCT5XXd/jlu92E4+OvKCTKPh31kPpJw6sJC
X3WXwxy5yBjovdvRRAHa3J4kQqH096XlXLBRhPSQjmPk2yQk2koBvdpp8ixvrrAJ
8tcUKYMDsgd2mMIUV5Iem/HRFh2B7Oz88iWwcLjcO1OEXc7nsn4CiY/OuH6URKKM
N2596twqoefufzAW2GlTd3Cm66fgu7lycQ6Qg5dulXn7RQSLVnR9Zc3jh2Lvbhz2
pF72uKkupKAtnBwUIIaVvAJrkS54VbKQ9C1K5lQvRT8WN6J1os+jBs7UtUgw/E+o
B7jOkbOM/jhZm/zmuZM+UMugSmZ2/doapCvZMGkh0F+d5AUpIBWXkx6jbiTZD5Ag
P8//COMNaZdvvqbQdLXhGxE2YJiM6vHHAIUCa4Mf/WjoOU7VhlTc0O0OZnqIOV1j
g8WZi/iQJRgk8ThkU0LvT2nvStAROsBeKpi/SN06cw33ZFyBCK0WUEZZh3aI3wQU
qrkH6tf/6HY4C+JYcV3EtzyRo+6jTsWsnCrH5jijcZvmJQqyfOCHgyhNhLM9hVQy
tzHvzPkskkS3/QtxDVEe73ygbGuARIebkjyvpck3GBmSwluMMceKhB/VnZnBR7fE
GOOjrhckMfehVYbzlJfUNDIl+POfYqe7H2AGkb25v1H36xg9SA/lZ4yWVzVoAbYK
4L7C+eiy0ytQzhJ/jxocjain+gMnZO1BMW5Ht1ewu4CkzXMdZVxQW3QTLOZkl3o3
uYdyXohbkG2C0SdmryUdlJ3ZNiY56UCCj8FMMidOz8xN4JBKICD6VZ6UrRXtgqFe
Y8vWs3cC11amXMPC8K4fgWNEJtXu/ZIEOQWsxztUQ1RDAJVXgfM/WfkN0AaRnea8
igVbLO6J2UA0tex3TBNInw/FzVOmuMFdrT1JiYe0q9coyrPmZjFqeqS8R0gJpCll
9s+FPPMeBhZSxJQoQGSfArLjMTx8qA0AlagJMjLk1+cVkva1OsVQyvNSoc/ZXe7T
URHPUSG3FbnxIr0RWYq8Ab4SXfaWRoCNUTNEJb3rfbXdIuIQUkFTGfS4wkMr7gEx
aOsy6dY2UQD5ul26J02QecbhGf6SlnzYTPRmpd+uTlGVKy4BqLB4HsPgl42JGW6N
hvq2g8DARGiJ2JoLtaAOjM80sVo+4ml9kodOOImyGGJACPst83jRdoExCQHhhglh
2phe41BOtfHLMQEpPQiwKxJlqJBaXm0c8TYiK0zUnZu/pPWBjFZfqSGCGaei6wwa
zqQ5jmhG2dUD4eopaQtgE7XVB/NMkA+1U1abaZIl7Vdxlaa+VHyQvG6wfxusdwgT
2axKAwkcm3GiErKtojEL8weH1QUNFOFm4Q6PHQPt1tvXZ9KSQPySwy5vlhnrGwTA
+u3Y+qrswLkB20BCo0bMva+9QIEAfEK/pq+tssEKH5afAIIHzQlMcwwR7U/a08x0
uAzh4zPSQEJhVFaQCiaZ2hFmJD5+giKXt4xPz3Y320UqbsKbWBr9hqtwSovC/6vZ
vSM7N/8gxye6QRQXKP625syHHoyWdUHkwAWBL1oRM//QmOJEhh1X1nN2k9lpixy0
vwbHvaAOZ9VTuuwuI+gecZSTbVbBIotinm/3/m9y+JO9MCUkdOsgio5ua2FKWxho
0y9o+2qOpRJOyYgkd9+tRX7m7F0aYJQA7yG/biZQRHnwQ5E6L4vrrT32CIPGAdie
pXg3AkvQ7ftSRdqMLesZPCGffCbTXnpCAWQFzYccMcj6VeoYXIhHs12l/oHOLfJv
m3Wvmih978VcaBRKGXZhEdJ5q91xd5Yb91tCUv21xJglQb9nllLJ82Du2p0RnFpn
IiwRffgN0QEGjZ/1X0GvgX6l9tw76SjGDA5EugGp3Cl/U2Q6DWnwlGAzOmre11G2
triUMjDeqFeJSm9ExUG7CwDzvOWPfnxxHZhVXzXrV08IMgy7d3JvrJS1LYT3kAZS
gSS7EOBbNkj7AM1dtHuW5GuVXWBPFAukzrQlzb8TcbGlLuG4g/didHGk6N6pZrgS
h19936jxsHOV6fkYxYTxDPfLQpUn7BCQ2Pxs34ygvBb4LXjZtAINTNzFscwkrPNn
u9lUbstLjAB0YhsCtl+xY/0ctYQmmzcQjLMkCZLjqN2OyeVYSm33YsZiP0/TQ1qw
uyCfyXHKXTzbhR37TFO9U3llMt80zkPPor5eRo7nVbaj4hSPHYoilzW6hoYIUaVW
Jn775ablqtvDKm66VKmJGwtthmtxE8yanba/my3slrUk4K8XvGyC5Kbwv6nLc/De
TlPV+AWDvj5nagHXcV9d3qiewJTJudjBY4HiDXWW9sCVwd54YKzNGwawUDuqc2S0
KeKrh/prlU9TG6/gG5sYcbNqhJuij+XDywbyxKBmBF0TRZWp5Rz7gBVCkteo/61/
hCUyOdVcchYPXP784qkdHWKKAdgPkQ7SSU4VPu6T1fkKMZ/UEoiPOTCBN5R+33HY
E5IWH7QyGEyrQFwjfT9w+jHCOUEOFtLwT7FwqdheWH1MlCxZdYF64ZVtGfvbMhWQ
JKAZ3oXUINo1V8AX9PDtiBNEc4gokZfwqVOmfGbiD+4Zb0RzuDPFVZXXB5b0P+h6
ou51MLNXNuHqwUEnVzuwWT9MDQuxwkEDlLrjFm6xACpJ6MqUof2lk7VSWwcYaD5Y
9JeSE8DC6HTRJHT+AbtjlxNWdu+VGQ4+fW6inYW8WwAp2CFwu58CVT0oDZTLv+Pz
3aTWIrG3aG29YOynIHGKemShFwa2xa+KBx36Fq64E7Pxj8ogW5wLFaG4jccIdvNc
eV5FGmXDIePmHP3aMlWsE7YWqDZMDVYZpbrAllVDGnv1l7pmTOViPyBxdDr6wgLU
9tbmWTG0zdqLZp6fNcQxZ+OJO2NQLl2+KHksebJ8pE50vT3W408C0EoibUn+IXiJ
XzVuB/kYmfFZJWfB/+Z1BG9YrOV/fF1xIaho3ID8eh/WfUqyyrD9OFRWic7DNqKn
limZ6NodU0kSTbV0FmhmONCiQZdKGx9YVo4CUPD8hjVr3t5taGWCXVDr/DslmPx9
NvJ7jVX4LR7xuEFahOg/blPwPlBqghZANRtTpHAcneb2fKRRyjYV/lEhJVkE63vO
1i4UcUSTF1l3cFjYKKUUuezJYHAmYnZquhXJXNCYv1/rulV6oDm9dWd7eRZ9FJQx
bAp0yD0CTbRNcTd6REi0LHYb8kIj7JUnf0CaK76PH0bThwfqp1W+a07n7Co1NxtM
muGvJmEpmqQ1T4safmBkWHQ/fdsDVEkZxcIfV+2LmxoyTNhx6t96z6g2pxqxclIF
v4AIPOZJ4DRvSxUfKml3LCkSnYSJB3i6xg9STkgs54o1l8p9nk0SVNAq4onTtneg
05v4RhLtVBewhVS9k2kefnEArfhXJ0k7HUf2jnfxUsRwDfWVOPGlJPe9Aj2U5XIn
j+7YRey9YJv3JpWr/HmJ19TbfQ9o/bXZSxU1V0eHQpD/ECtb+aSD0XtPp/TDTNjz
JlGoGkG+jq8iXVONwwrBx89afAPreCBofLyuEnt3GlD9W1SpdNbExr8Hpr5mxeAZ
zoWNo+OkwAnXeMyuLbfWV6jrmQKBX3GV6YN8yolhD89QCjhDXqsiEe/wjYWAShb0
o0xzK+SaaCA2cRQjbqcEDRAQxDGkLphKu0/60CWCpH7G3bRyWLOAogf008MhCwWw
XALDi7KcBQtm2hUIuy/hO9Wco+nEwd77TEege0ISl23PORubu8AldmQlaFpomAac
szke8c2w39f2szyTbFz5C6e8wicRNDiS9tKf21QmVt8nIWhwmJ3/fG7AB+Uwqkcm
GT98WiVZ3anBiEhGmK3RcRSm86Md0hmncgrTl3zvoXnQMgFl4Bt81yFQVkqFJq3S
jLWarCJGUV3rj411JlykG8uaKmUkuzDZvO42OPaEQPdraLmUqMEXCpEmV9jkBzsf
+02mtoEbhWrrMebHmXTl7YxhspFsAOCzB5rJb/AiV8SFgeU4/ti/toqSwvOySCy+
InuxUSdp8xJDtddGNHpuFJqtQAcMJ69aC144x7sPDy0IEdRAriknipGPG3BPHe69
TmF85FNP5ANuy7tNDj8jKERMyDwkc7ClS/JzVKGWNJN3BOaSda36c3ZxhKOpPk1d
fm9Kur+ZWxiPvSkoYHTJ+2fYWXhT/DEUBgDGoPhNF5hcVZ3o3Dz8zh/kXXILS0tF
wHSaU2Skf9qq5vel/D50xM1z0X9lAMoh8HI/I+Q3HdnoMXSLwPCXALtI+kCpcjjV
O2UVd6B+C3lLFMF6cS09ZRQ/qrBl5n5FCq75qRIiJleZCFcTQmcQdypowekP7DwF
7nZN5h/UAGpdh/K3kKuiK0bIN76rgRfBC/W74lME16wx1Q9pw5Ax9MIJm4Pa9K12
yIXtP4LJfqR/RtPzmgIJtTPEIKQSw43OHTeTxvvRReq7Fdu3bsUZ6JQE4IWBN4k5
2KFrVVeQ3My5DeudOMNx6YSfiM4Olfhs7sPLLXHWxXDI/OuPbPjkG+vdbQcqrB/q
R4OoVsZNgbZTOp4dlHGGmi+J4ltn06Ld83u0GCfCEuC8Fmh20asjdSplizwyQEbt
x/nm6qvdoGmLtLR7EGZyA1iDMaWBNbRLaz5818tr4omMOb+pVHUqBNPImzCsyXaX
ToVFYNuHjnYyCFOqRajIWR/rHECGePewaAA9o8/tReZaZ8uKbzJFwYLbf4d7wgxt
4UW0N5Ihfqf9BSxvcoAgGLnHmRtCTlQWox0VWCztGasA0wmOUr32onWuT9RTgtgy
OY7z8jHza5xqEJl3IwozH6cjI8+zPwAHD4X8qYuYGP2PWJ3kB5ApKwde6kNrM3JO
ulzyDh1LI6l04MjkErG9TX878UBsHlsG2/nAt/LR2IhWDqYtcXLznEZUKlV6fJ+C
ezVCboVRwRE9nCpsHaifwphrjyvfK+YT+Bx0yAgrNEa+/M3zmDObCUdVYSQ6ozzy
Q3Zm5pU2ja78otqCGvIMg8d254IQysdsptq/1/1IvBWBGQHFj4gTu4LSjB+c/6/G
mMog9D1rgxjEFBCDkbHOoveCz/tRDyC/FyK0QZZ8zmXAHRiiAfnjTN7/zeXkTDHp
v6xMkofqWCenAIm6K6vTKZRR3NEd3117GZB6oH8vCjombrxb1zFyN9YwVDfMtEik
nIl0KDvz86jSR2ZENvpz9VFTGa4FePoL6Yxcqg8FyszYhH0gBPop8Fbrz9JRjFEU
X9RB7Qh9g/D2Y5C9qsArTlEiD3pnTBbS8txHSnUZRjozF4YEkZwp6kfu96JEs681
BuFx2vXIo01ucK0PDN5eb4CxUuIVLNnedmnSHZAvFqS7f5tihnFxQ2cNbpSlJDOY
mqtK0Lh76bTaEQotCuYboW5f3x24Dbd2eV/HbwhQV2t7EreV8T4m0615Ioo3c4jH
T/7izu1fEywpE3XCTA15AW88+EC1qn22n9uvqTyReusLtPKIfGWQJxj4+gEcN1Wt
dEzk+BstgnMuqWVLw9W26OxjvkMkhUgFF3JQA/DNIewcW7YjkVv7Xq4kor84GqXA
iwOYrxFsFYyrqaTtPF+39JidRSbfjwsUrdmT1m6Vv8nfAUQoGG2MTxaQR1/48y2h
FgQtujCp1DExiU6X6uCtFoL4oAflkc0LJeXAXOS3LgXr/V20RCjJXpryVKrKut6s
zGqBT4fYlQEsW2ji1yy0vnrnyyaU136v9VhisbqH5JMEbOtefS1Vk0buL8vZK0/m
xHWJuSyf6/tZv/gp83qtZMTHBDIbXp0ebVzg2Z2vFpZfhbGYqHLUCI2yDEs5J6CL
3vn5uYwBAsVEJ/q0eBxmZVlAFzJ3J4ea7UPumxNaHhuQ+35jH8bSPzj/K3QhahlS
oIQItz8eU1Xqm8xEgpWttiRKhiwqGJRJ03iv8C+1eo9CCbTdfX4MNIfrat388rkZ
P6Nk/RvayOk3D7Zyb7pUhw99fcJbPlNsJGdXjvzar17cd26rT6km/7YC3/AREo5I
MR8i09Sj5sxlHjhR3pmHgmzQ9b7TEIexjgxN7FThSTuRc+23igNPXzB4KrYEmM1I
39p1iyKYVDjSTiOCR3YbxgZF9wVcJRAEJ15zkczXEACJMTBHH57YM+/2Ce6yWkDO
FluHKVe08XwRQ5URMPGFsgld038S1O3TWSmCaW4Ee3ldssDX+ZXUlp00ml5QuMFx
dl5QY8ylfnZ3oto0h1kE7DzQumDiYnXkP11s7WSIX8zRJfZb26dkc9y/1ctW2gYP
+vcm5NqwaDcHgcwUK60CBXOEcuYH0aX0rVxeKUCjW5EUOdKx+HuvaNWcZE5I9BnP
mb/P/4tvtYDUFaVmuGUAHvq1beXXI9+oF5Cz86Wkjwp2rdY+PvvBZhTeTSVb5H1G
2XL4EPFreri72qEv2o6rZwKEkwQI8jnnYHA03DPX0ahmDhZxEwKgy0Hn5LVKk424
EhgAE0qFzwzmtUDDpvK2b2x+gnr8oMpP7BhOPycN916X5h8t7EmEF8s+9+PHHfn+
HP2CA8wX1+I+/kRxzFAdeNrIkbBLWqHimFYNc3BiOuMaFGFoFOrXdvfJLcgM86M/
4SeJ+89bGOtNWKS4049jt/G5fI7HqKePq/CJRcDpKHDTyHjU4UyFC3OyZLpCfIR1
/gTEh/YylgDemfJzkcLk+5F78CAf3R1hY4g2YAIYHV090KjJN8AURBe5kOzS96Sk
LdI7J8NoObd1+ZYMd38QZTGt8firNsx2zlusiuxG/fIqECai+7dSsyI5zLY8DGVW
FKZzwpK4yjD+3zEkSZlGT6HpOMZFJQInBueIliXfW5wrj+NMtgXeO9c9/JSOTSJs
kXTHjiHgWCr802uUIJrQutkOEKd6hmV6ioJMgv1gweq+DhYr/fbJKDMFq15yIqUD
bewErN3hUo7PzphNDZbWfJCzA6lDQNRSPD4i8SvipKQazsxS2+iW2ND5QEtVFANi
kItN0it/x7ntQUZVyunrKaVDdqMXqhVPg4Qcv19pD8oV7UJRElbNkgeIS0oitoEn
v5guoUFnrkQ3XDyBkBkJKC1FdLelSXjVSj01Ko+VFkEqi0sRuqQ0NSFncKHwkedv
vtDAxLHyPXntoetjUENMPrEd/vdlIpDH9Ngjaiej7zcoOofkcFSW366c7wynMgqs
57ccrRYsB/+5wq+D+0gYleUzoWh7rxaOkxxRZF1EEOS3uJJMZS4PyzF/0SDEJ3Pz
biAQeRktJ6jFv8aE/0Mx7mkMS+GvPTLnMKLPhvGkhaawBZD/Hva7CIGcqjqZSTIV
dxVC94O3CVwYKmIrZLJVIz9++yyUnqv/Gl3fGj8+4qmouJ3H7FksTWvxGr4Alqzo
k/Qn0I8lXUiOqEXAvIhmaAXl7mVyHQtWfib007VgitdzXhrcQlcLTRYsCpSqGoUW
9eFsC01BcIulCNDyQkaAryFdHrz0ykwojGCN9V0356DfmjsggUTlQ3oG3KqKyjas
KbBQDoGlQk2TSqMGVE/UfIwaY067TTQM20zEf4M1JFgttYi5KjZz8AWL+zTwlwLu
71LPdisRz1b0z4sBqzwxal7YrQ3mlVThGzMiAZsM+tbwjU0pRlmshJ+N9BNm+qqV
SV7emd96Z7esPRTqTkGBjaW6iQunKhCu+ZkOS9gLWXeCzc7ymPo5e/JY2tlt8/rn
QnHX7Yp0aOSbR6E2ROoTi4m3FteUakSUP9vdOiOR+k00zAl832NBpOSy8Z5NToJb
QxTYZErh/POFDKTAU8o28MtHjKeBvhLMJXYwLRW1nR9RYwbLlTbStFZQbzzcpWdJ
0JLleyKc6DFUUsAla5/kKWDo5vyiytf673htnLsYJr0e4NOtQFIXkdtIcDPhLErB
vDaNGYJ7JUqUcwFJ7BnBgX8OWBpzIutIYRIgWN+awCrjxtxYp0qCR306YpZMDsvN
hfFp/imTavhbgLuqUgKRYvh5C/vpDkVem3yg0d2Q6Awd3PSiflZJ6WVT3IpOQMfG
pSHJeVooIfqlkgK5A7km75gDhyLH7tj/4NMBd54oeJa1LVFLVtwVqoP95KSV8P7X
wifDerC0/f9EkSjYzp8mCS7bzvn0Y7bh8VrRinvJZNVjfERQkZ+b3U9RE6CfP7T4
Tu1tfkhQyb9jbw+6ijMmRFAXJTxosT9PvUFzZ6reYR1vR4I1J4aZiFKz7m6M56y+
BuCY5yKQEiZqi4g8xS/R9C6PeT8/D5WIXawciceEufAr8dXuzQ8ZzyRbnAVelY4O
mHWMnI/AgivJYsS5gErXFJi9yM8z7t1FSdnPH2LAgbrXpVlBgaFcwgEwxNERMDps
zygkGzkxkVsqcYnu1O9RpBtEh458TQTHlJoG3KFLV/UYM5X0cwp5hMJpLcnO+P+h
PvO7aGGj6wtoMsvaOvmTRzcXxXGnwUma6HpocLQEkGb++lbLBs76LUfO9kBhpHHI
cYUf6IxyqMK9R9xZJhgln4yC/XOa+Y1M4myA0Cx4aesmiCcOKNGDEKn1FdXyMo3G
mtU2JXbX28mC/I5oyPdu7pMCtb4OpFAMhUtdKoKsKoIf+ngkeFDKCnscG3JKjf3S
9HUeHt6hdiEf9OpmKtNA1Kij3EdnCayDGxQZWfB+52VQne0wsGWyIhhAHpSWFl/F
M/FlOYmYkA+6iVsn5BCCHMZAo3hMfZXSxxE/PIvy2+FvrXmaxPGuRLJzpiSSq3Xe
N4R8imIalKL1LlG5iY0DMgEnhUoEWTza7NyWuc9g+J0K4Jk52Zj+4QUJYrvq0YR1
ZX8Rx/UoPUdJP+98WVNvRT6C30oNWVHZSYalspI5yu65KJglfgfTIaqWhTHGvCMZ
RaxI1iZedL9Kd2ROEBAFKAH/H900TbVxyJfD94f0eH9i1FAu7F+TcKSApiHY3Ztg
t0Yowpd/9kH38MRtxcMREYprmyGdmOPgQdAiwsGBhUzGVg5z36ERM/D8GHQ/NWqY
e+V5gMJj7P/PrDqSL4Y2FVEVkmeWaRPMXrYT4VhM8bNe/cIt5xMPS7ZF26YCY7Sn
92MVnRfWACEjI0AKpOQ7q9IgErju3NZ6q/To6QeRkvCFJu9cjpXUc8QzN6TQXV+U
DwUkNhTSu07+nODO1oqQp+GDw5kP7E4aNqPP5GtdpfrCA//xQRnAdjVy/Ey/Ub/J
7WgoLtLrxg73lGQYvEZA1iNWPNoYyjc2qXJWZPmqZ2ezLuYzlmPVLfm5W11ULTa+
BNzmx05n4V9+cdY9kghqhPikF8E2y3FegSSpuNx9aEWg5q8JltDGMMMDn6O+1dpL
xhZYFmEFrTs5ipWGtIQHiE7WGc70pyEo7kzQvlhg8moqCP7WUY9+L7YJ0QeT6toa
3EjobwvJ6r6skv5vLW6s0lyYymSnwjUbrp6UFtD21tqYEdz1WVipP8V/cNA+8Xf+
iYRlZbwZC61s+ogM1x/xbjachYl2JGB7iqSQMS/bqTF5co4mYsGHe62M2/G+02/5
yzvLruzjvFg5s7JBit+Dm1bPsVkcVZje/ejadvi9NnlJO0jiVf3lnucQ2SUIifX/
mZ8qj1c7DDD+mHXuqUVV3StYfgxYG0dj9zzjxIBKIf/AD7riAa7zmn6PM5xQgXOw
vm7YEoN+f/Mkh3AOycMdc3ECMB6LiFZOGZ/I8twARv07w/RIZpyVmUz3nrS3x7ev
AW3ubu9o4w4jZQtRwA2rG7c1o9vyindY74DWIK3O10Y1Usdwozu3kFiLwibJIdrY
INlP+giEKicp8BIkLvmaiu+U+fdHMoXq7RhRhuyJMb/obhoy2DWGkwaTms8017bv
wCp5vPl9FMGnMZbOIyfrOufIZhdbMnbyOqnjtPvsPx95x19G33C/OkcTr9XTVYXE
HN3LxqL5R6ndnenDre6N3B4z24zyZ1Sih8QmCd2S9+icgHabVYEWtWqva48BCqXc
MyBBdvR63v40+vWfFx9lZsm23clD3cnLur6mfprt5KeaoT7Kd6QKeObIh25HYm+U
coc7zQOQ7l/bzSQb9QUqEVy4YdXLmSy1i8jki4ikPc3/gp4LIK4OXruh30pDf2Q0
uKPuBGA+8vqm9GQV6jrLl9TjdnEsGGWCxNLJHtSML+NjZDyDAi2URUj4orObAaKu
R8BhdppD2tLtUmyTkUpYokympAV9/MxkHAXgtnbIcZlcqzhpOBGZ10NrmpWkgtHr
Q+CFLL0+zveP2jz+2M+YTnU/kj/GM+itcM6oylCUt3jRJfTMXB+6JwA+exo/Mm9G
Ane5ldCUbrn3W8arwZUDtOy+s1Qc2ESHbdCv3gVevHIk7mKg59VVyG9Rfq7ute7O
h/XOpY4ny2nTjznjn2DiHJO5w0V21/pv58ZlHYs9p9RPZ3Hl93dr9YhkDPyzbYh4
muEArh+Qp8hTceySRsEwrEdjHqM1RaxqTHWHVPsEpSTmq23WiTWwKnMulThJycEP
M5F84Y0JWxjQI0zAnVvauAJQJmreJ0+bu54aEM4qegaNocbAp9qm8VfyyzoJ5NJS
IPAt6biz1flCtdvTyppJBrSVCARfjZ+1q7LX91UC/KPwmKyx72V0vKAJK72LQQ++
M2kCTpKcuuiVmmhHaq5v7t9e5ZaljavYBJCzSzzopdF4PTW/CT0N5YZGywRaAwc0
vX8nvrY0BHaKELy4kAFB8ZNwm14fP+6MEQ3ZXTKEe+2VbT2ZbfucdTqoPZ+8o1Mp
NOhxw9eF7JuzkjGSjo1ZATBDbQrAAameANeU3BWa2Rp/omPcd0RTniTV+eM8l3+I
SoHy1n6L1ruxLQYVMTF30l3D7S3Qeh9FGdcAacwNDGSQukUKe2ey99MMzQLQYsbn
z5ixSPJ/YV//lSMIRayajOcsADU1OoSU4sXIG15R1z0t2xynu7IVmwOzeATcp1jV
cOw0/lpHMiqE+7+oc8alZIRyBLASr/THGy/5KKvvd8D56ATX1VeJkJqNTs4d9OhS
ZtuhQ95hiiim6z7VlD+WUWds31P8zRhsBOM9t10PQUCKlwkBhMF1FsUvaws2ouDD
YASwBQm5APNxrEZDBnzseAGqr/QSE0OTWjtanTNkWhXFHpi3egH3bci7Z0YSW2Ly
B4gHUohWjcX8ca+6KIX/86JGl+DGEOpqxoBgNxqdCgK5JtwIVaFL1yag05UOkEG0
IuhkqIi+BB60kTvlWi6ss1hfvPgy8cpmzCvF+/OeYIuEyZs6LgmpVA23D6bC/7iS
GVoXSR30tY+StNJcUhVeEkFqvdgNOomx/ByRofdOvhy9ngtj/yXlFCLeJpvhDTXO
Rg7Esu8eUXFq6wRL7abCJP8r2tZcMf7qGj1tm8NZ92pNFwWf6ik0HVwm5wluw734
kEbLnw5sfXZCqnouZ9sH6MwYI2xZP5CwIJhKC3w7tdSUV7W6pp8bcFevGyMCim5b
17zhZyMg0iQZWpHmKWXvywTK7SE7GEYIiSAc3EcNKv8+CV8172ssme5PoVShEODR
gIKWmAWM9bUVKmOVYjGmb//zD6QzVBgW4DzVY5j1lkaNT/drrIfuhWlPeRequ0eP
iTsVWl804x9BtBe5muoJyOQTg5SUG8fHHpGHh0xucLF7bOlzrj3+fHCOP0v+3+9k
/k5FwlWqgYFfW2zVx2lihicjiFN/GtE/srcC46UasTxnMOU1/dLNJGxZoFz0oeEL
Eka2CwHOeRhfaWy4Kl+fRyUpAymCNP5R+2o/tfPCVdoZ2SXZV8GmIu+dEvqAzEHJ
eyo/DJvNApUS6IEUgaFEGVX5+ldSTPmSq4xv2l67b0inJpUbYl8QbT8cARuXeKHQ
Czy0RhUaS369MYUGiv4vOhvHu4Tk2nRiR4WzLLAXITralY9xc4B57m1w+LkS5yuV
RmVgtN9G61G+Vpa1QeJFMjWW9zijwTSm+OXS/+ScfpLFA/zzxhkCVFulDsAfMUYI
nv35GUMkJrgvUcVKQ//5eB8GlZVmgSPRqC9ez+wwGNMJw14bKjdnYVsOwspjhGDv
A7R7l32K+Y+t4vWncTUHNE6Rh/gaHy3iETwLy8WtCMyAu9nsrxHoMOoW1JnO8Uo7
7uyrHwUBT6SCh3JqMYpefhCgJI0/WEnIts+nuR5lYxsKFsRhA+m/Fh6P1tzUhheO
zlJihh+o+/+ia096qmXfOdYDMBClQvt+yaHX0hPDbJehylH18l9AAUH+cYdeyRR/
b6pEXyS5h0YueK2BTVv8h4mCKrJQnbi7HM9tqeRd19TufsRVMtNgWlWeKY2EnfmZ
KY1N3WzfHFJDiqafaWg1v1U5DbSwbju6FWTOMkGmtl4rhPNjmNlmil6QmFveTiga
lGHLu5E1339EDtYyjkqjHvrZy5cNIIq+vZW1SK4U4gMEqLOlkiicmzzBuPHRijtz
cwwOsreh0acxBOCg3apnekY1WPf083kuqHxKQEmBg8zdvFk3O5NGH3WCnBE0YsOW
DSjOJmQNfgIKVmjCOzZhPFUzKUIh0uaxNjGPtbo3ZlrTicFw2In8XFsxl7hG+NhE
S+YQN1KMFwJ5KQnACRf8972/q50v4NQss0k0jIUXjuaSdM4hkQSMlCiP8lv7AFpQ
W62wZSk5/DHJl3vE5VcZ8iLkG1v7qe3G9RXL3+ewXu3kTXTjPhwQkNJEDpY+Ea25
QEIfb0Tgn1tofXaVGVWrqvZoEMtjHUiWOtMRa2285KeCE0fg0oTVzvEdZePQ7bBo
bNy2u8SShDKEKkPMhsizcDkD+AftTmun0XHAHHji/ZkcCJ9LZq+U4xR0MgHgIho8
I4ZVxL2m4tcyCn+9gUWEl4phA7IXkVBQ98+n/yVH3rcInozYh6VcuLvVG/4xNzE+
mGKVVWKfJrxxjBQvSWjkojylLsfN9+l0P0K0uit+TiVm6/L7VU5sQksfwNvU2HO2
vWB8Ryb1UvCyzyvwbWu8g/nFz/P3CTkQGEVYLbAuzB7kea2b2U44id6tUU23kYuu
9aqoHtzSmRHW4nlzlUyr3HAa7dbS57/4DP3O1uA5gkhtnBPFF8FXQiRZfOom62je
+ZIFo8vHSif6FrhnvS0tZTGb1ainLNTkkNAbNrr1xp0TQiphTsXNZ1gW63RYn3n8
Xazhd6BhvSR4DcnJymQ11daRP037riMd76yuatuWY5n4lxAWGS8UtDkQwx1/++1n
PgfMCc2QMOK3QO4pxGfRjZAvtCPNRdJmPMkyPeLroW+jChJd1jXMdblEcxWYEPbb
GKD9XlrUIaKPaLCOhc1xcHliQlppN2p3eSJOlZcMfrQ6BWLIYQy7SmN8EK66i0nL
OL7BbCS4PZvb18iIuewoM112LTRyVRIjTeR3RKUnbfIIlPp1JB7RfxH6TSp/hKl5
KjRoDAqYPn8oRv2qOCLsZxlEnKCLr4Cq+C7Yo4MVaI0Bv8kOFwcmUQIuB2+lc1UG
G0qCeo2kANp0hD7iuhMA730eNDwGohJYe9dEtRSTTot1JENbbereSAlHEf+BcLlM
NXbDmr9o67tl/OnwgGlC//ZgV2WnbSCYr/bl6iN8hdhYDNxdIXCBZMBerPWpCwa1
A61ov0jdR34X5BFipqjPFiYnC0iaxPPc92suCPGyg4EDKV3PwN5eBcYd+U3jaw27
w0jKI4gCNsut0WE0Hod0vbC/unDMFu3Th3Mha1Wr1UMutNjq9Ry++F5JMmzZkEvO
TC2seyns053LQy2h22amMj9hcdyIXPk66mE5ufHaqcnFg6p6s6Ch5ag+u35mHVXd
vd8NRJSBaQSf4XaHqWXJIO1SkPBHdCffpntFUjyHwV5h5IqjUq8tWGrHTy8H/2xL
2tiuT4p5UNzeaGRHBJiXNKg9OayAElIA/SRw5HV4HIwl/f94vkcA6wpv2SZEQ9zm
GrI+pMhXw2m6Evxl1/WKtJwffOpf4Arde3WtdYmXL+r0obk+vpArYFV8S8bszRmA
xmySNGaLt0bujJYi6g7amorwvF3ESbHdnumVFqKodEpUzvAAcFgBrC7HsZ/DBAOC
L9bCrj/gvfLLtrYJixV0zmuLG9SRqj7IfnnKI4oj0tBMrBAP1qWkeyIqwfsC7TwY
JP8ob+BIYRi22Wle0THQNeBuWchZlyx/qWfvdMhyccII5DMtSpAmM+kgGVZI+1gl
N1Q52hCoDzy2otKArC1PKMqBgGojVa+sB2mRNfCEQZRODX6NsZdOJub++V8mI3ZB
0R5GKWjUdLUmDqp14D/8H5m0x+pRcnURLh3yCjEvai+J236/wXnSsTSkjldjXFwD
ksrbiVfnQiKUbo9p33EzLvO3mGujbYam97q/4KN26YBKFkSlJ3cQIwKGty6sTBL3
maRMb/8MkGq9srrC+CEoykPJKg0U98GsRnOY3gxTgCI9rYDhr/O7/V3PjuTE/tqv
K1HwAmbBnvgI8qX+m6/kCIQ/HwccMXN9rQl4ZOriHsUbQPblSZr7K8QEOa3+htdc
4rg/+3Ijm6g6GnUiWJwF/KOlTY70OBQ4tZBQGzRF6Tqhg754mdI04CNOAYXTHmhn
txEvI22zRrAL+z6PlnPIlbPbTmFezoiR6Gyt0DtICGgmzGQ6DVQBtkqrG6+8Hs4g
NkeUlY5P4EF2mS8666hnPyseGvNcx7LaR/N/6TLxUvOsZbexDQVqlAJOdMjGz53F
uu7U3hOVIiNjgGNAondt51uAPgqUc/jj772MK5TDnZhcLVB0V4hIogOFMyoL9eJx
W7iTt/adHvfuXCeknw+BcxjX/Iyqz4QCkEDcZGjGJAKXs3U8OnpPJCDSx4ZNcp9k
Dkr/cYHaIu2LAGWDjzSqfEVXagQsTZw0wPQQdqJ/1nJT0KcGkgM0oLlOBC5I9R+v
v/8RXBM42fiRD9ku51Dj3zjzZy3uPmjGILlhFZIZFvTIFGDailmFVWygbEWlmmux
c8NRtK/AED1PFM7fNx1K5zShS/iFs37QwIhx7LHCvJMzViVWI+9pGe+3hPTta4mf
bUz9VpKIeabhZ89P4LhVNPC656yo41rp0ngGaO0UTU+kTFVnNrNG87HLpo+ARRTZ
nCTtvKejTv1oBiCXhousILG+gKdq2kj9lsxbKBsMHNaWhr/fAddU6xAVfjYqykzy
QpGTOOAOoIUMBPXNBLsCfFD4qtFJyy9i4GQaVnyqNAtJXyrOFiNvVbbqyBKRLCVr
DZp1Mb+77DzRgQ5NICxBH6FNMDg3lUuSRUcWVeC3Tgwb0JNTukiv46Epwce3AzuP
SF5mb38NrcGUn6yShwvCskjbkg7QM1o+jMJWHC3lj5xLjzV6i9ANvikziH31qEzC
5YecAJJqiGRvhO2BrL0SV4CyJMyKwVOvBneXgmm+QXeAHvDiaUC0zJEXAyr5F3XE
31nrdbm3PpPkq5FJ4jIiy3GCT/JVS9oLmj0OcFtw+dWGcd7rs3n8RNfKbeNwhvnv
qrfGW+saaBBAJXB7hdWiy2dkyKUDYmn19eP2W9FO5GfP3Y0YK3QqHCga5+9dQXMM
eE9UA6uE46TA0DV8ve5Rc4zop+IdNbG3lcuYdu76wKDGoxPIMt3n7nHdjaFvpDwd
UZd1unLhAyET6RJKxpWbhLUQb0kg1DF0jDuI9NOzgyfu+68ggGufA8ZdYr8+5U8R
F1t7CB0Az/Q9DiGe575Tdf4H2PTJb26iHyT7zZPpK12gW9aW6+aZaLLe9+AsANTg
FpmdMCivAkC88VtKEYCJRbguBY0Le59SaqaYMrviKDyaB/rX9qHlJGu2CF/XZT3W
f3UVA9C8KLalaNLgqwlui1oInB6HJvEqeIcBBkrgoB+8JT5TfxwN7xYCr0Y7VgtZ
nbK9eWUnEmK7lqYJXukLBLgTZBiU9UfhB6m0PIuQZ1fJvwae01+DzoDaaD5xUhcZ
C3D8OgFy81VvnTpPmJqER97SjhvHBDby94n9YDrFrEn9jU0ITXbpPZr3fsYjXDg9
4w3bDGEUEwuWPVV8OhPlqLMWFTu25SbZNB9ofdVKe1ioA9elFP93FQ9tZeahtqUe
niVuZX5peaZaEu8z9L1lDjSO6WxTpNNo3kGhg6mZLKgyNOEmESA9y0ZgWUneRos8
yY906AGlS/pIBFM684VMXJx8EAVPwxYq9HRz7zAW/xWbctPlpL/Le9DdoA8M+rCE
HJtpUflSz96gfVGjLaPYQeG2y+NbcC+8caNTerVeq2fqmQbA/RgEJO+6rhJGtnaP
SnsYEP/GZ8GclrTAJCrR5R51V3H8MKGUgGqBMx68kRv3r2v1B2GVNVE+52Fv6CpD
WGKM0d45xxczCfHQMOyeCishZoMPRJoKUk2n4j+2yZbAWxCkakYOWNXRM1W42zKu
Kwqxj9FKRPO5oG48C+1bmSiozJ1ixKpFSkHYR/iGHnjAeN+XQwDOzhhoZeiKLHbP
waoBnuvx9dB9CzO0S56GqYbzXZmW/tFvLQRzgcuU0sfN+/C5lifG/15Jvp/QL1IS
4tqasroIEOGTJlPrT4DlDgudPxDB/j8CLuvNOOyKjsU0KyMvmIxkaqJ7o2N1TdcW
wlGASKK4Nqo6Ch6de0t9aPiEtPS+VHyWm+3rpsy3Ot5FIuUOSUrI/8kSLzbk9kl2
rNOCuh4pXXeIAA4CoVh348COkKa3p8ijGUL9jfvT0EwSb7fRl8ZsMUnCulH0VXZp
RMIEDAv91HjeD/rCKplJcRiowutBem5IPf43AmTwKPkZ/zD2Dxvdm59voqZ/oeT0
3BlD9bthjRSLkD7Uhp31lqm/QSLolIffq2y/OgK9vNOefNSzASXzcvKNToXnYALZ
iiyWaGgcUKt8Di5Klx2I1WCtZ19nzTaa0ZJQw5M0vX2p0ot0N72G642M/Cw+aASL
L2faLYtz039CV68EnuQxexSuwMwQ0/toYx8Sex/YOy6ggfoVDZq0Y1rBFli/f5ef
p+IHSfNz0YL8mF0nM6BBvG/hOcQK88Yz4OY/+bv9v+/MamQnxAwsBCcbXXlLD+Iz
IPmIwcTz8OjFH6IFHH7ZvRrLBSJXz7qAsf2OpzJTaBN2cDc+Ix75dIQXCj25RKcP
bc9hBFz0A4fcqkGTF+Yea74MvdTqcY2R0N1VloBq38aIDlSuZxk3sO8mgURQAwpP
B1uHehbE+Ix44KahoUqp0XKz/iGuur5JTE7JvooR/6jgSIgIFxO9NR7lZwNCk9P/
er745aGm5whCebm9+GLvw+Qi4WzavHEjiA8dOuKo0FGEl1hr3ln0yDr9skR8TBqe
oqmj6KnyIR3xC2piwBXaYCqwTNFdRmfPH5fyOrmvxGDyueeyKXeSJfCnc9yhAJp4
JjH+ZkGwyylBmbjYq9QlI3DXOMO3l8FlSODzvGBaswb/0WeyzHWnV0Rmy2wq5avM
XZNUHF1tM/9sJVIvj73+pe/oeqIs3jMquUbCmh98Bp6ZdH1iR3UYekDZLrSuEBXD
jTR0e8ygxmmXMJPUlHx6dl3AkTIagfUyw2rGRGjQk17CY/F10CsqdD9+At7RhfEf
bcO/j182c6VxUgCJf8w4fhRm5QkTf/KcoJiUJxB8/0h8GmVQ4eW+7GiZOCaiCwKe
nfOsFiHIQnX1r+jLkoFAIq4bLW9l6XTM8eU2mZuwK0c4p/1pUSc9K//cL2z11OoL
YxZF52+8kCf+FAce3dL88g6hF6Ngakpq/4e2oVF5a3SSUmTVZlMhjphJ8qZRRhSO
XiDkO2DTi6rwf4JR1K5gmnMMmv9HHNkh5cybrypNkCkYbnQVRHkelr+ovVy1s7dY
VXL8t5x9OaFC3Aa+Q8ST5B7bG9iQ+YePt7l2s7WWfwknsDR+5wefUj+oFFX77EKb
flhBSOuRBKd+Ir2Bd0MDpDGf8S1vgvQ0bEMlfeaWwsV2zT/YCBngHVGv2MYyCHoE
3tbD6l9vP9+jRAkRmy/tLtTtt6vDmRji6V6Ta7wY/Z/TlbpYEBcay8dstkh4D3bs
7VjE/D78FrcxzlCv1UHRXgYiOt5kCbKyXkVTVVi2puVysZ+BzRZOxBIUMzqYIRi9
k8ufg66axSycN1kJkkR5lROD5Afmv4XVTFQtM1Byo1h1wxr2UO1ksrXzEs2rKlKK
D+SdyTdwuxqK8dbWtN1iIRiES9O1fcQGfdpdHjm2BxHJR2NHDempeMFkB0VP7Bdj
uSIue6ntP0Kq8wvgWG9s86yfNk0VsUKPsndtt3bmDVBb7ojl7EWBc8/x7DY55bw3
2qKbYrxLsbYtzs5I7TaBKtczR73WgaFL+G0pd14fdG+eU7LkB6Mof/hz9CUoGBwR
HXlKk23aKe+HkThKCLnm6sXFN3kQkCWAWQKkUbLSGGSqtFgIzGSuhSyomZIPLjPv
WK0m8AoRlxrXl9UkYvNPsxDWFcprzxT2v8G4A8j1K2dNdzgawjfYVp4mExFZmbCw
zw+fEgeFrMg+MOOjWxXJBstb431ifoCvM8bpgk3J8iioBwW3T3VZ3IyLRGNuZ9oe
a3TJa3d7bbeQD5hYzIQ5TtoZ/ZRyIfvZ+U+XbieyDBeAXQNraZ6ibCAtTZFMjg5W
dQ+cj+pGzkVnyiJ+Pz4gtt+SRBGNmjdule1GyKVfUVNO8/JcObInZQwenwePGk1n
GU1W6QqBFuCcFJdZk6BDM1x1pMaMXBYOj8/Efg1nPYb/UhdANI9JzYTcrlEgxE/z
dhWNE1SoeH6Y2r/CPtpzcrHk+XY265splFpSRmOGWI9HMQYd7Ena9HT5v7/Y873+
+h7MTpcHV2uBKsucouEJxOkr0i2Acf1Cbq0Wsnjcz0I+NLtXHN1BvIL5EKdJt/92
pxvocxjiDQEpHSf7JmcbYpLMfD2wCMvvrdhapM17MoUtFi9lgC6guNRRUwMPqen6
vyb7JsVc3oLN0O4oQeVVTDPiTEGuwfK05kOFX4YAv1sHOYyx0MeOXXqRVEXbVwrw
e4d4YCNprTafsKA7/sqT44cYBvkHxXXtlgs9nuOrnAZAXQvZPpl+lHtmRjATcVJP
LL+wS7Y5jNwZy1xjtzm1ukNteUaver28J/DfMO+JrJ/vvLXTlNFpOiJ8pAGwwtll
d/Js1x+w2QW21JsBxhn+INBexvyNKWdasQ80wHk9gc+vnptLUZ8djaIa8fnf6q7+
w1/xPnvT5MqCsjpO2CyBYK2Otw9zchGrFY+zF2+1LE2wLIC0c0/G4JYP/NNFKVWz
LxNjEMpElevWyasEamt5qFt6yAzJzdNENHy2DFjUQcZd3oCX9s9ZbFc+cqfeMlKU
npYJJHE7+FOAO3nXvIIYMAHqB2ATpXVHDIPamY6SXIjZIn2tSkJUJkL/cpbuSH3z
G/5On28SOyi7YvUrqqW+Zfk0VUN23UHfhbmZcDq4CuZpvs+l/QydktwVkx4zpJXd
RN6z6303/Ugeg03U2emB5zuip5MEltYMn/xY3DGZK+EyMd/kpBin95NkyTT99SBl
YpTIHj9ETibAeSbySqR1nSsxDb3Tj1cYbz5sgCVDRw4gQTBsDO0SgwZh2MQpJB3L
PlnRpEeixKcne+1MQT+UmOHafr5E1bX2ZGaYkc1HHa5+gfgFK7zhvJXCS9u/tPos
bAPLAdfE/Mx3oAznoi4cQJK7eAARcmduaRFKBq2FBH2ucZQOyyQcXSDXmUey7AVq
n8BTox5XSN1T72Aeb8Ayc8ffOix2ol2JLuub7nShqf2GiTPSve94G0w5g/+Of+G7
L74oS5SPV4ZqKcTOKCq4Bcjp8RAgZ0cAJ2S9BeYGO7R+clz+wl0ECC2kVNJCCiFt
WJDXR2VVoaCPbT5UWMWJ06glP5NeBNkc3fr7zHpZU6RtZ3Wfx5uZ+DTsnvG9p9FO
5WSxSbxPudmKyw0/Z4riVCFnHvqwz9uJxxJk7j3B/FhqJyRtwQyz+fJYs8LZ41S3
JU9YZP8nfFNxr87Zm+x9UY1vaIAc8+jImTFMd3qi0WmOjSaR09qZkD+qEePoho6n
2NutII/Cm1eJwtyjv9HuMZt52vi1rAh6iy1vObd4Kok2S+YoJo+79lRHels2by5K
nPHOSPDnmsSOOcFrR5Lp+BA8xRx5PTXi9NB8x3FVMmz5DBTEduGNZBIL/4h6wEmn
oEmt6cYLCJsaPucpLSrOn5nAwoAL8lpSe+IxZzbbG9sO3cSVoeWK+9xc0VhyJ/w1
bx+6efpTA7QGAw4Ui7OIlYiJWwot/boSZVM4ZHy8ot5AE7Wcmz1ngjGAN2qHrDv3
tAf5Mq7r4ZAQ4EIMB7BNnz585clXeqDKGhUVqxok5VkjaHmSdBv8luSMuYccXZ9Y
hs/QCJXJeo3ngFSGI3eLF9uGWY4LC1ibAH6tyKOjMuDbBN/jSRtCs/48mcZlHFKV
vw1GQqFvMu/DyVOlj+tO6daaHAuSPn4sT99RIZAQ4rzF72bs1bBzFwzg593aJhAN
eBx2lcuwB35uFyCDfZnhg56sU/molQKJ0C0WwexKhrA1qBVeZA67v8Ovav8M/rdL
8mJXp/Vzuv2l021rAcx0wVZswSX1ggNnUV6JldOX80Ke61F1+SP6XTw+M+99uGKv
83jc0SKEeM4JoQUPJHj5iKhKRAxEH5J2BAapzhzk/NaiLzaZnwCZhQl3SwXOxM0O
wMMU4F8V+ZiZPx222SRC22/ghgToy7TXfI2IsWzj2BuzBXvyC5cS5AntiE2kXTYh
G8zJ5Mp3dQII93J+sAu556nb//dOyUMx/45qtyDN5djh7k+FRoMUTKiQ0O20/HUA
JkRFR9rzQx+Czy7TicydG6mtVkRqCKiZD7c0tQjzCKnX6ri4I7sAOCqREL+93/x1
VwQ80vZC2lWE7/kwtQcjzpRPMq3GKXOmtlCPEtwwKyXfb4o5fe+rDczwymtbLf4y
BfO1NE4jbTylTCJDHtA6ickKoOxnwVnv9UuDUUU2BF8ajA0TcKQSE8F6OkrsEJmG
lSjDf8rs8skf3YHMU24BLWHV/ZjPBR7M2GNS3FgSd2Ru45ZQ3Gu84sdhrSMFGbAr
c1DtCxHiRQaxdHoVnh2mSHJZIRHs/L7dOD7W9r7xSeXynPUqi8xNZ16OzFTHb75w
4SNQaL5AVsRAdNSltuNtVFjC/Aw3ZvBfygoYPNj5rgmhBEnzp6TVp/u5rigIRXt3
eiLDC0mneBh6gQoFNenJbhysJhzn1Fa1MDJfEr6kziYV+oiNW0seSe1G3swZ+b4C
izzvJw6ueddKPbHkHvjYVrQKPWbK3F9fah+jgr00o5RiC90KFgFq1RSTF+Eb5T9x
Uewm1mKxojgeO1mANPDQUU0xGplz+6KqDw0dlnPxXTHxBRrzZx4ZYgeAy6UYhem8
pjXFL18zEa08vtQiwPkaBXcg/8wbCRhMsGlEfOZyEsKMszSrMCQsOZ8CJG9a60Vw
FL9ENOxHWK8uWoeOQlmvW4F0K83qljSKBZKsbUJK+0shwm4+DQENwaUKfpv5Taf6
xyChq/fK5GxO6Flbnqa4qUn8fwBbLvKE0xfWH4dAtF4q9NKxitDAXFKmWGz0V9jh
0VLGkFkWHciOESyQqrE+qMyY8ZH2/RvlReu+EfnE09+kDsXCYEbos7OLx/KKAYeG
AXAxm6bArZwOREYToOk4P9kJ3kvSafak2wbgACxU3Wz4nA6GfoMqYY1zcKW+/F2O
q6JIxVKnsZ9EludzvYa+0kYUR4PaC0NSvKdX/ugC09VoSDMQxvj7TLTy7P6uiKN+
fjo92idwR9Ag6DvHzAcGf6jnO6uNde+vfxkVW2GJ9Bm5BEXL1Ebo/owKf2ZTla7i
I8rGu9pDTAEQsAl/5jK/ClCIBVs4eKUDoxJB1qGEHmmwch2cVzQxcHEn1UPKBQ/q
KXCSHg8NQaigoLK7soeWZzqh0ybK80pwlMkVT/fkrR9kg39pD0Xg9QhOVmm5z0Zy
wl4H4R817zMfXHRy6PoYr6XSEP/N0BDQUSE5tcGe6GQ6nXvwtqDSGQokDcE/MHWl
Wcbz9aCQife/Jq5Pbyn4Hhw9IRKOQEXqGG4ZyvJePqr+k30h7hgDP5ZMs8NkZZec
rbWLNp/i5F+uUyyYU7CcH8kNS50BmOGlu5IYnEzXQ9jOpwtDV7RSRreE23LD5n8j
sZeAUbVQWEBpXg1JZJfUHdJYtzij94DGCryFqAzeeSAu5lT33tz4+h2TszCqoLcT
uk6+P8UWw70tEevSmuacuK0phtgfmL455UWxSFS1x3glmHQ4Iprv/BRQxn4O7CXB
7e1P2hOdoxXiOLLuNVanV9Co94wWyE5q1YKIXJe97u1SwYm7Gy2DmzM9IN5WHsA/
H037Y9g9mOHPHDT3XYBMgSuH0qyvJ2EAq2oQ+Wevxe+tTnqaa9u+xo25noVJOJyE
WDffNTGIfNOP6sghgCirkhC8Rvy4uhyHB/qNDQa81fPCqzocc34yJ1p9N8Cy649c
ZpcpnAOTRIoYjlDwWIRP6+o8HI+al9+FGtlrYC/fT/OObNzwNVeZeoFUGaL4iknz
4IUCbE3tH+R6vTektCCh32HUnEJ9L7XJWu7BM1kakyvBf22Ighn42FjTHvqUrYuo
Zq1Q8p7G98RnmDkCvw36Uyu8xRBfFIPyqOXjHfKIP5gjK+k+MQMTYZbHHAJpCwL3
1wwZLjjHTn9N8dibkY9dGYJTmXLcCw/BvlGlZCY1E0EtZ0G6wqWZrFFiY76qP0yn
PkmL3HhZRJCirhNmJd8CWISw99zF+fCfmK9mkWRS/uQEI4bWHdMAb2vxSELJEEpk
E5A/nYHgzT5Kxi7Mpn1xVQAK4koRFETiVcL0F+yDgKdumIgi1/hhJ/hj/sVE9McT
zpIpFzjBx7GBmx6R8UloU2fSKQE2Ve102lJryKImPvoqVafsFaYc/uJawXsGDHpN
xjTXRBvhoxKxvJcTYbcytvbqOP1zX5rF+gYDipSCvWKYsvwP9ivp9j++XGnuFwLx
bwEqJ0Z65uGIfP1yrKQopxYZhzvsE/eOZBi0MePqgrFG7Sg2eHTLbayfV98CicCK
mGgEiPYgYTCISqbaGS9WSXmlQp3KfE1OrutFUlLvBBoJDVeIGhAAAKifru5CaCkZ
4UAm24vL01LfqnzwHC+2U6tZIpPnjDxHPOoGO6i0ooBqoeYl0jO990FYBfy7ZpSn
wkNgjQLKp2j4iMP7h+VzmCNy+VkbYFw3nbvK3QwToxg8k+Ew/UF3FDXSnH4Rq76T
HdAXa/61RUroN2y8fUad7M/mMIcmxgIazPM9KtxbODlyi6okUZcMrNvugx1V+v2X
Qslr65uUqFyx3WThGbApFIFp5F7GfWhn8uKJYjPIFdt+4ynpyEPqJsdaiIaX26Ni
Ps0Td40ircfHGSuDMcTnj790e+8pHH1XQ5VgyH2yM8Bc9kGQxyVSiXZgzexpNjs0
kbRehoUCR3DJiplzWeG6/ylLnRjgnHOidxoBTm/lU5mD0+0X6cmOjEnxj3oxrpN0
PZICtaDm0CeY6f9Cg5T/VtgFZ1GHLoysrgdzPWmOs2k3jPCzkYqmTNgHqNEcZHNj
j8QvQQihmxnvuYPJzB1v96NRJAidTHTIZJKs4eerJBf3369DeVjN63onrfo/W8us
qW6+mVwdaAv3LelABo4PBV63zYBtVm0id7dfUqCOiwSkfycgLeGysGy5wJDo77Jt
mhGa2UeMYUABUdCpyzqQKB1J6cvrlulgghO+EfqTFFPtE0wiboT3mJBIpK1bvrpf
/yChG12xMisNdj4ipf5K24W+Gr7tVpfXDDsMQ0GJk8yLEWcxycA0OIAGTg6LozY5
zV+xuLi/5PA1OYv/8q7PqwxQwK1o02f7HQLK2ST2oJkGy9wYl0TZi6go81i57iAD
SJVQ3SgMj4rcgB4CvYog4ezssuCnnsQ+ZChH9L1Q7T6X2tY95hU1/IvhFmvW6RQJ
X0j/Dnf8IuBHC58KSiie090UM7LtYDhVMmY/HL+z+yUGNtSd9rNtTFMms1ABLSW1
+jroSJ7OXUqzMHYuCAsv7nRRAVd3u5kqvkvqLOB46d1TQfiaTbnnP9sGMKPp1p55
Ly+8u83j2v87TpLUEzX5VfkD0zc/Ucxz+Uso9xxHyWs7swaTLeg25iOtOf/LK/ve
wQwfHl40L5bWOftunDxRa4rR2lUnuJpfVEN5PPvdA6XZm6V9DtTuqT0JtPl/kyVC
UFp6InjDhKT/2dxENnYpYZAdYxBFBK2gR2U8VQ/OhKk5rLIv2mdfGtDtbWJ47uW6
mie2SwMrrfigUIwICrPsgWGUREH6TbSRmffCAm3/jqLfOAeOxdsTbYoxpSWAL4BQ
pAoCyLS6Jv+HZLrE2Gv/aVYKjbbuaubbk1FlKnshWz/Uhf1iScSZVKYib9D/BZSF
kh4gwSKDMG0j0Rr+vYMkdQTK/dgDw9AN5JnLFcxDgt8j3MQWoRQve3H2B43hwxBT
c8bulhJn2PasWlOkow/cg535PfTD/M7vlj8E/ymOqonMWJ4QhIcZ7ZZUtpiq/mT+
eCZYUBdpGgTR8htdhxVkp/+UbqjEQ0jdau4TZ6ry6fDx+Jva3SZ4Smc80KpnZfX2
C5//jOsrtHYwjz+ndz25qmb6ofeJMEs6eBY+hts3Blr1+baCYTkaoFJkOUbhfZYi
CrYSsMNzcvYFmZYG/e3oOlICoj4Bo2FMtKYd/h2QEMgUiRLnMv7NmCKoJ2vIfdkp
zU/sUvBCVkRosZvojhF8Bfl3VRG9E56ofz2X4B5Vvr/c029SbP60M0dXr82kVBaK
iFgg9CcgeFfKICO1i/JEMDa/A131rEyPBtKuBvHWxn1H4a+FD5ewHsdtoTx/k0/j
QKxU6Xl/u6hCObOwy5noswCriJJTI3Wb3AWcFv2YcSWmFnbjrdItjpUEMWHCv4us
tncdIhOXmZsfAN+NOWyWEP0W6y8n+/BkBMe+osfWts0O9Jc2mAjJjcAE1dgIO5yj
+7JrGQlQr4M39jwvUdwnSr53cj6Nq9w0xIta/cUF5JPp7fdTtyT4bLpvIpAasZeb
JlvN9Q/y3nnUeyHMH59s+cF4EASiGsVlvL1u6wL1WNbUaemELrX9jnej7lluGIna
46atv2sHxp/t0bw1ggJY65nTUQ5Rn+9XSu78wLBvePmYM+qoYGNwLW5aCsWviITE
Z+QFFOpUNuOhngG4TQGSg2WgNZFuc5Kkq+WdVFRvkdkeWCSbCu7mo4ot9KOvNPch
1qgUOPSjswXFbJs24hoQSXOe2mziuQE4luP8vwXyXCucL4laHxizwxAkLY1/eYWO
Yj0bfsP9kr6uPiox+CUtt/pLX78ovemAfwlURSl2oVHgyT9YfyET3LDXWgxRubg6
RKcjp9ndVU2NaL17jCEsarQgn8jyD/djgHhbSxh1vn2RCMoxS251xBDZ8b3bWApK
aqB8agAPY5cAUAHD4AB6UBt4xBsdiXsLpOPqTbLGHtehOzElXTD3yW34fn6FIlCj
Ll6Bh9KpxjMBfQ1NcQ9GE7+Y8NEJf2C841HBYpj3YU5BC3ALoGxhjr0Yi/6C5ZPe
NjpPbTeFsbLOOrlaFmIBbMWV77+ndLbceT06qkIKKkNxgMUNXNOh2lkXV7fdE/pE
dpQYys1k8U2BQm3BFCqG4T0jx8AajzxNgbZz6zwBhE8dtnS8z1eb77CX7dcoq9NM
4KePeyULASvnvue6zrU39SSXKdxfqDfZVoUtBZ/AFNatOMPIv/1qGB0GvQnx6+Y5
EsIqykvXA3+tmU2OUeEc1hJFGU0VS8DmNUmXAV7xpy3CGO9TfdiMT7rVIo252bVg
CSxO7B/9/Rqs7oLCQGZvF8FGuVhEJSXdOckeaph3XFAQkLemT9t/XjQkRlL/0v4P
spnxlmkoHEwUtRl3wFQHnIWG6CWVET8hup9ZQEjwyd9SZTmbhYJFuFJMlseHI+C0
WnIbbQOEHN2EpElE7PGQHTL2jvBBYAoJUQKyFR/+dJ18rGq2/INUlIy1iUzo876W
6NmqN5VwMMtJP6mVcYk6EO4B4NPA1EHRyxOfUOWu5u9z8TvStkhdN46osgs+aj91
LBGeCWSqj4cyS/QM/Wn4kQJbTlsqbJZuQofmsodRKMkV8RmU5ToNEAa2TWdZMWq9
++Co3n3PDfov0t4mvteSwJDeyh/TwF4otdegXRjm6L5k7MnWUlSQ/0AXxb2Rd4V5
0z1Js8oFBsVjg0J6l0oso+C1SGlmMwSIJ3JvNfYNz6sufLLVeYxpatwJPklIH599
wLvzqrBKSMLReJ1OwEAUlrQMPiY9vrbUhBaGNVmJxJB00gc7Uzd0ttrXi2760K6+
jcrIvqmcJNjcCLStgJ9JS9GP3lpM7gmFQtduhwwjeU7pMC7YuYSmGGffty0S/J1E
OzGercYpxkw/BMlFaYJKmx07nZIvuNi0afsZqmcvWrSgCzGnhsAZBLkN8TREnjTi
h7nZvzH2yJHGCEVSGv+qnAnHJmPRkh1SVh258LMiKkzxjNrvlYaDaW3A4qszgphZ
Xi6BlzrWqdF5ceIUlQPL2vaiTGol0Z06ckKDhPf2qR8Xp1SDBMxd9VXFeXbtT6eO
ys6Vxg+s4fRnYQlIcgKpJ3BUS9BZkyVbYqZ2NfUKNO9JnsElcKn+ARYmAhHCbQk9
yYiVEsqhpYcSdyuph3n2udRdH/isb2nGSPGklL98dLAadkwU3n7/QqBh87ju08Vm
hftavI9lg6SMwHVux1yGoXkcm8IElDxkATI6Xaq2+wL0ozmsUNWYgAfAfxWd9tSo
pHQ0KpqVD7uPOFDaUaP6V/KcE0DVBiTVnHFeH79BNo9s6NOssbe5iq69gu4ARkjX
3aWEMxkBh3oY2Bo75z1+vefRBQ3FBPTYF8H9S4FFpqe9XpOq1SsEGr/dRcTkx4m5
Cjz7FQL/WgIHqYScvlefc+VSyyloz3Tgb/mUYcBZkfUHtsS+b2I9l1IZMUJz7q5y
Skskoa1lnymg6BshuwIe/ejMus8TSRdpyGlFw9y5WE6i0OQhUec83e8y0Isgom3L
GHHA+Mg4yuQrjc6KBZSlum8LTawHcZuL6uELK5A9QB2/29kcnkBMn0ajfHOVkNxY
VmkfpJyr8dB+QlEbCeXkWXuMCP383+6SW37QKS3YMfUEH0hvblKgU4EsGOsSbLtv
oU9BwPtMpTsCIGTjBhhRvb0JCaUFccnI5sPCql9ni82XDoJO3URQiHGN+GN3YwUr
tuo+fHowNUUtr5EPU5izWaBiwd/TP/ICCqIx+ZtHMN6kfbPEzJcpUUIEJHfpJuh8
GvkEoCmYYFuCSdjLj7c44aq+GZweWC5Rq4W6tndVBTmZ0pAU5YJPGUUHniClAcwQ
SH/SylOIGvYY8JiY0CFa16Lj5kie6ySe+Hc1qwXRieI56g9TtmkXNWMYlrUggtLC
t/07RkrybNr9R8g6JY2amxataKCBLbWE3/L+BXhenI3kBoyBIhapPs2ZcqCnE9Op
jjRnYdJga7NXqYzxJ6gQmA9qy00MgpuEU/nbJgti5mE20aMWPeJqWE317KerGmT5
JmY7Rvu4PjnApPa+E88hGxhsvzr/eGNe49x9z3QK6D7mQL2DJpekEanUj5Zq8qt5
bqRB/fTUAHanZZlxPuGYex8HC8ZgWYCeNFUGYUMqOkcRDreaClFSCZ08aPmKQpiI
6cWazGEP9ApcNQLhbY75fNK5oh5fx+a37+gw+Okgkg4arUbzRuLcZZ0IjIREqoxt
9zpj2tUD9JIIj9jnYW7oMXMN/bdmLtw+He/7ooIg9vgIiZk+HlkBIRyoHAPo3fyL
WdU52UavrUzi2Wgv80DbQWXUdQ/wgUZhTZH9ZCljy+s+PTax8Uq8we1X2O+iLZf6
puJel62ZPMHdWkA++RPNzhncnAyP4eIlF5GtA0yuDqzkdI2BpZecM8L+tmefixpX
umAbYfZxApsR1WmficcO6Pf3TxqOi923Dh79420GGOascLuP8bOM4OabBPP/6Sew
TWagXpwaSDz88UBIbGuEtqkWaPDWp29XT4tX2NqjfM6H60CJuiEICkg3JkfSq25T
fWWTiSxvTqP8/g8/S7NORgU/H0AadfXQqIX2lEGBDRSUnjn39xFZimvApQMUdCqh
dFnzWmyE4Fdt/FWxAnJf+XboTiwWaKvRnvPVKFWLlvEKL6dGR43w/pXxsYPVudqO
TyQUHcdey1UD0AS2ztsmcuZe2NX93roXZV3rNPh180sBH1HptGE/moIhagwFz3df
c3Ad7zhW5e2hGbTccnkSGfH4GeRKhiyDls9YIYScJDQ06yv1dKOV8qSUVd6EWCUe
fhlCNCDdR/j1838d+kYoW0ZllQSHKLhOrw/at66NNFRg3Fh3gUWFYnZRYd3/407c
/NB9BEJXA7K2ykuSPeNT142yYnanbi8g0ix5qaauJkI+wZZbDOzkA81X4QxVrvlv
Qw6EutuheqLFnF7ueO6Tgtr2+vNnIGNkOevA4Gx//O0XS/g1qzA3z20eSD20zona
VK2eMtIhBbuArnw26uNVuiOdjdAr6MgREQ/cnw6F9Zdu/T85Owoy4LJu5GTaKT+/
dz6sdAeTwNAgJOcWNIXT9BOlos4GVyM0oRK/aq1PilMHf/u9/WkENb/hRKjU/4yz
EbmFCHmS523R/SoYHaHP+PLTCsjmncgsisZlcX9yMWqkNxL0VScOp4KEaWWmgXnl
xSvB/XZiQcZ0ApXecNqrtr8G+K5omhKeSrKI+KlnzrVptTMMGzSNHvyeeM3G731y
5Bmit1ujtRmvqryP+4eW+w3bCPzcD00Mh6swI+0zQ6q/4vBrSUkspqDpcLhCOkiv
5QsTOPEWWMNuXSUC/D1HzZsDbJwcvEmyVhy8PFNrnLtBwp0llrDjv6/eq14rixOU
M57h5ZrwnLpKhkNpwdjfeNh+LU75TWR8v1vyeS2Ism58/TKArM0pda/NewJWY47p
9e9j1nkOmRTaxNHIh8FnszPw7NOcaJgctidWIZkVOGvGsytt2W1ch90AJAjzyEaf
YFz7nLhb9VEnJVO0m9D4OrEayTWEBlGH91/kyo2DvnmPfMg/PQENGl9MZhSbTjeE
035u1KGQmbn++VJTGt6NxhTjs62V2E1FaU0HN4mxczMnduLB5ASy7qPssxWvgoRE
h7mfuzIJ+5WZFXfRjX03yX+4sru/G45vn2s++4zowONdvLjBjDOwZrc1tmWx6NBG
PwEzi7q6oWPf3h68Y0goy/3Y2heuKYo0tnwQ0KWYz2cSAq3FpQPcF0oG1OVzl3SY
kYiAMpw2A+vDR0mFzMVtlwM3ijmfR1YApi9Yq42nxl1m/fLS02cXZxV2LTyXFRh/
QSaj3xKsGHOOMWNQh0de9l8HKar1XdziNKTnur//CeMI+VizTosAG/woGq4+4Chq
Ha28mV6gnuOBsCEC5nBIIb3wu5SE8iX8gC3GhSM7TlAsOkodq4/go+22knrDwmk+
+0HcsSrL9Z8dtjLGtnslmzcHdOceChSsCM54fI3QHNGtLHlmmf07YwUqhd46caYW
TQldtSiVhVP0I2S+ywLHtLvEhMV3R/W4fIwiknFp/HfdWV5chub0NFVFhjH/HBpb
5V2xFPgmnFZK/Up1APWlieejmL2vUEux7whDcklPASphADvzXJL3i/1pWWYHsbg8
b2kuDfzvRFh0z3KlkWtL6hPmdLXuAYLGANZIwZkt2FswJ9TpqTTEtzD9bTb96X7m
rejuJEm/y4dvat24fVna2WeJMUBm3vNFUlVlsDrlquxukamJxLPbFiZgihMk9eIG
f61mehIqZkaGB+ioR0nyETsBK6UXb4klbwH7a4yj48jlZ+zQYfkahyxv/TYj+TYE
dYQ0v+YfS1ZQXcfQ8LrmJMmiVT560NKtNMJt8x04XDai6plZ2vHPn0bl4n6NJwdv
8WqsqaWSMEuaCSx7c+RH0nULykl/66z0R6sxg2xu9G4xaNXJPfVWA/0JJlpBfMWO
nbISuJLeYAb/K1T3WpZWlKx5GYJ99QNAFLZePpTU0Q32h2Cxhv1KWSn9utOL2Jmh
qoUPG92aotTBCL/c938czJ8ZRJN8aFK1stkXM0Tqq5SBiH5WTvtlXlbV0rfu87t+
n5gjd7wkUl7Eiu036zmx2c61lfIUOKdbc/cXdjcvxk9O6VCtU4nu77yRcW8PSULF
Rjl6CeKOmMyBpYypKOMa4DGzsH9/3ABpYwdAxVddHy9PNzs7ZI5ddjvBNkBjqkzJ
yThREfGlvw7qhgii7XrqBhzcvLkZvMdtrk3APQNL4h3zdM5h0kep0Rm/lkQT1Vkx
MGOHfGrvVdynnK9shwwpNoR7TdtahbVpCPxp0IFJPrbxX/8tYE3iMvuTjt432CYh
zNydhGkx1MBaNTYbbmtLBCyS2JFBHJvO62aKsADIBLnAoDIpO3SoGU8CW+xcT3tB
Vs/LjIWDIT6DmgHFa7d13vSrSPpOJd10s2T4OjuanRSo7WWncVIEqfh/LM+TVfo/
GwtwM9MRAbGY+xZBcHXU9FrIuH4SWli68wvIxAj0EyCPP7SXF2USNOJIuiN2Ooac
j3gG4TOO6WlWi1xqZJSa5mAG/U+VjyxNNQtesLCs2IU8fpTxcSBjF7127Ps00j2x
kPJlIdAJHIFhPJuAqibA1+BinWFoUGVvzalxJOd96KiHrsTaqrnlIZcuYifPHqgx
yNunIIdT5jOynirlvnkQEyPRnfyxLo21AgtGx9cQ+1NcmYNbEO1LP5KJ40IEIJph
W4em2tt61BwoFmeVvvQmcXnj5vE8Ok6iHLdbIOTgTjy3Um+kYVHBfLr4wPc5Pb3c
PNNoktt3NLS/+5VnpP/yOKpcUmaiv+ozfmTPWUEFlrE0lhDb4EP9CpnIjn9sS866
QTQtHVt7LkrYkTvz/RK4hPdWmaSpPVxcRahxdt6C1BXWgFjpzP1CfaBJ6FxP091d
17k8k6okcupXR1uFC1kTmm27s+FbvfgSPwwwz+4o2H0ZVSn9QHTcpu43jYbqtZcx
BNU+YKkCQ5JMua50vHuquXh58+acpOhm2YzYqHRH6k7SNhtnBM9KnszY1+NZWUWV
uq63zEdYzWlnNw7tcukk5KSZ81fYN1nsCJ0VhuksZmZOwcxkN3TMGTve6Zo0WENE
38ijApB21B0b8AmqbdIKvm5IcZuw0Ll/lYDIDHArDNmH1QEd0NuBeiAP8d58haTq
1S6mef/P6K8muGMS7UBV3yUqjU6Ze2HcvedgCGH7Cc8DqMsOJjix7RwtWRiKv1vO
+EUHlFH7gYaIIkXeDq9PURN+vzNcjv42QydAgPBTOcXxJALamy9YeVI9s0qg87gO
MAyrmY1mgzvn0m6koolT4Gcg87ZY0dEa4QM45D+BBqLsf8+NejqcK7jvpys8D4uB
sQHAP2Z+xpbEOWePX1gxR5OLH4qCwE4WJOkmRgSzSkGLmKCajR4VbMdP1YahBTXX
dBBoJRQ5jN/wdWDjcLBTaulMB9gT+MVakBPmTb6dT7VjlNMRIpcyClbqqpCkUkV9
kMZDgSLSmN8V+vAZI2p0zlWbJa3+wwbXMQLnjk6tMAyhu67TQ4uk2Y+J/y7OdPpN
kyw/YkipN1pAHD/IpTjxzIbNESpO/8P6dMU4l7aHmtCz3gdQPtt+0xs+DvVddL5q
KgdzRUV7VBdqRbJPD2Z7UuKNH3zOCFPhSMXBCfHryjfeYxgYwfNfUoCvf5t7CBWV
UEr5fN6QxeH7mwmKHUnLCt484nLtcISZgvrC75WrrnFbwXWkpAEwHdy9IM4wBVSA
rG3qMesLTLua8Gz5QA1gQnzb8Vcp97On5uxHXX0+b09htL507LRPFRImUPfDr9J2
qCy7ud8zGWt5y/URecTUOwf0eBz178eRNHxfihOWHH5CyFBTrV8tftzXPlTmEzh7
sOc0A09F2SUZNBKMYF5BoeQ5Qrt6GKEJTc4jAFl1W5v2Ww3e5WPB0C7ZymfVlK5N
2OpkcbqKGWjEomGlLASsNBj/UZpfyeO9dmNwaHdPoagzlL7S19sl9lRIKt6y4cdn
Bg1VTmHskpVAuiACnSvT+rMi/NX0m4gvz1FvFiajAAkVCE+i73X3DF4VnDhgWnVZ
8hzt3okq1oPL+bQ9Tqe1pKa0NqPC/kBL2HC/FtIeEkaWAZnDcoEJu7hKjo69fn0g
9J7TCmF0zdrfRINYwav5THB4DbEmefwbZExYmbSNTyBQUcaMcs5+f0fv8tSPudML
i+g1DuMldc17B7bjFazCPxI+g7rsPKFT6jHEex/qdqBQgTcSeY8OnShbbUQxnJmd
azlgK9XVxhrMoqS17AL1ZhFpUWOlop4OQY07yc9vmgS2YU2umgEMjd5IoHa25/Zo
8FNh41kG4kRzJhjLsoUQBbO985DCPasL3uBTtf17OQnrtJsGF3Hy9kTKBzP3y1VI
A1Cwxm13aPvlnClVYcyLjTNU1HP2MHiinB6UjqUFdC8ShOGrYS7QlJpvUZ/FY/J6
NAZtiLlFu9EEp00YWf8gpcVlrzj2H9SAB36ebhB25a7mi/Evz8FcjPhHoJh0PZw9
0/MR2KvOBebmBPAd6Bb2x+IV85S6LuJXpRbIej6OQ8flKzlMWQtkN4aWl1yGJf6C
f+OGPP8+ZhOd1NwfIMa6qWdOftueKljhkAExIsqHGiQhB57m+ZA3VkzP1qEToPvc
rUcotJz4KwOvPqpqdlUGHohVEmD183dWdUWNZNiGNNnoEjSlZvjvEk4WE8VRXl5E
9NcvT2Bif+JhWjKBXfWFDpuhwpPLMX9LYQPx7bFqsFSucdyL5/GvChrH3Vu45zHF
BH/Pognw3MWface38saR3tRbJNay1baZ50gEe7sPpXCug2Z5MsRUC6GpnjFBvbuw
PTL9xGgLuw002T80gQp4xZLD6ARccKkM5+rhDEpEe3eynQf6PaGIrmAgPgyo76Rr
MJkcK6HYBQvtir/x7H6A/fu/Sr4NV5tSW2I8BtKEkLuwBfKm/phF0opmiKtP2vrz
ASi59Nig7bMbXX6tQbabPgrVNf7cODMuuGzzHtWr+y6wqhfrxsw7CN8l8EVYziUq
BAZHOdHj8DCAdj861WcghA0fukLXj+wr9O8DiWwex3PaAKjsoPDTmA1cFugPBow3
om8wib+jNCGpNTOpGbBTALtsgY72NZDvTcZ930lPICS4bFsDhm2NEriEWScreff8
LLSCPgB1u49Ofui3AUVVgMOy4ItB6TYAoTECHX8sV5FhRah7tkJTjrEdTSszWhHf
5W3JGJ5myaKZm0vm91ztPuMECXBCUduhc476wLu/UU7cxmDg2UPZ38X1y8sMVxyx
3Tln/62FaDoMjjNLSERfXfUQHCpu+hfTYVqJX4UyOy/N6vwc9TJHNCTTPzBIbAHK
ZImWSuTxTyvaxwAQb6BOH4zI/NE6XOJcV1yEo3U8EKw4FpMHXWNpZx9lJSEwqQ1B
mQP6Se643R827/PgxzZj5puK2qq6Vzl8RmfD4nWk1KAEUVndG5/xrqTnC2Duz9AM
PU9qekAtzsXFwJLA22KC03neP3V/f91kZlQAbd7P9fK2OjCBG0HdyENX1SZCy59B
HD+5pHQZw7ro4JsiXLeEKHX/krhkP9gI31+DhfOoIY7GuSPLTnl312Zf9jEwbhfx
1GdOXxHLQyUMWjVt2lIHeJrlKMvfjEpBnw8ltM+t3xf8qlEolivl8pEOTsbEYo7o
9V5AQq+wNZ9qokD9LfcIUjhFV04jjLgGNK16OjmI2K2YbkLL4GCys8GZNMVHc91s
1Nt0jEgsCdf1Da2RGhkk5WF+XEDFEpB1b1Xv8v8Po70ObthzuxlLm0JeJrQOQbvl
eUcMJFUDEeOa0Bc/1Fn+DqhwwCweZQgd1+QHm5MSCe9OWitivLR79jO285nBNxN0
eO4Pe1JryoNgKMZtbt23+U1yXg2REqRxvcx0zUXsVRifQjy0SU27Q7NkZr+TFOlD
mWRf+xH0LIN3RblBKvmcRW3fomiKrOKMtGIElVmgSrnKdbkrm2P9WsSQDOXW1c2O
HFf6ny/iI5Y2rnvqlRNV2OrQXBa+HQO/VNM8Aru5Z/5C/qp53EpEKpDXGBDruPX/
gMVEwD37ktRKR+KFkYuiwLWGldWh4IbKcf9BGIomMq7MMhv/YC7Y4Odia+NG3Ydq
zpVRRWCI7tpdnokOTM5c715SmYddGQLLiSkQF3NisWnih6VOvQddb/mZODHeRkid
vBW5NlLATciGTUH8JjPyQu7zKjCKYpidHfa29O1bRPVjKDel/DHt9bqx51X4rND4
bjQUrzoxLujNKt4xYMyBlFvzRxKGQPsbic5S/xIhjeZJlikUv3L51gbsQojusdqJ
4l61wgVbSvoQkn+HzoOGAYh+Y6vqnOrfiZxTblLvJkKxpQUS/yy0C4GA7vNBddUj
oHz4mPCqNEIk644EWAFbwJS/nP1g0HZLTytYDL2AkqFASJ0Nj8KqHBHnAyeEmMuQ
R48LsG9wax+BCAny6StbC10+GPevnjK82QNEEeo6cPgplGQv2WVuF0QeMpYsze9S
rjHneaL80y3OyBrirRoXv92jrzGDJSc5ulj8Poy8tRzF/t9Dej2WgDoZZ8yFVIjg
dJPfo0Sy3DsQO6g2x7c9OQ3m16763/6N+dHZyN4rs3Y42WvnRc9Nxx4IoKSBdhFO
fJGCCX0dKE49+0F+aIgZY3gVxniNhUHVlTJvfkXnKYjsTINRWuAhzbzb4ciJOPW7
HGuFMWtyRhOpgx4CkRFw0i3J1AL/WlvqLkRJpMyfpE5xF6d5Kskz60MC/jlXg0QA
zqzKlM/ZQj7EupeIdD0tkUEF9HjaVF3GdoPOyIG9idUJ8wOeNIJt+o1bCSe3m1Zd
N47ljhwbC6ejryszczI4MpMM4JTMKbD9tfVurvaevHmENvKO19nzdPjoxhCfHuxP
38JOlDP4e1lWeR2jdzajAX3iDT27Mq8sxxRHuV6aA1F4uZzbzTGlwV07qiffeunT
jHrT4MYir9nWkY6J3v5V/+ZDVD06dmV/OyLZbumlUM0zUcCCssdSLYRxDVz8A4+4
jeaClQ031q+gYnMVBF+hVQqYDClZhq0Q3AlxPSRU1LIDIyBM1DF0CutEL8/+fosT
cjevfqhLIs8koWofG+AQsPkmZlZ0l3FNmCerPQZmG/5cHjfLirRFQmuKOOjx1BHP
CCJOwZQ0IhzxCt4KXlPG6R8qWKhJO5TWJab08mMUMY1zZkOMT2E06Jw3zQsOUsU2
+Ru6Fy/e+/SEl5r5ch5kuNkYfxn36gpU6xTlnC0aoCUVnuvbqkBHQk5PVXOaDNx9
pbGu9BqIsU3yNtzAssd8obqfIoJH6NtaybVPBKWaaE8D9CYCv62HbyVi57bYBWwd
4nnof45FO+md0EC5/IXEpSQMG4zAkLP09bJjGOrL+Wjmj3ZmuftXy4OJjmUP9iId
dSjzJtn9EBROrseZ2MpY6zvtquaTT40y2B/cxlXmdMTwnAC79aEeiXGTw5ea6e4m
CcSjdPrWpYkFKgtddFJ0q9m4RetiXBOWBWirs4RlNt7EOWTdvOT2gGgoTTKG5HZ1
1V3zk8YPMNwQtVjjat4MtwtFHEFzZ2DJ76izaCRJ8vgAy4b5G6e6AlFmwtrytbCY
dok/1YJxv47tnIIV+gTRGMW/j4lbmjMgrPD9EVXwPA21mvk3qWGxTvp6pn7xiV9J
z4sN403aBpdJVB8HK5qQh0CBjnC3rKIIVoPto5bKS0CPPMvUi4CHe6yk4Xhnfifq
bxo2s7WbZBkHPbxJUo/EmRUv24B5fshkYr45IXclGcXNLV+9cXqNZ8OP+56wZ8ip
jouZTs+ZIF2Mgi5kR5oKhVLsvk3GO3+QLO0M9B/SD7/hypu2G2B4LkgS/jF3zv1X
nMZKq7aKd63NjtugQa3OD2cBWiLalf/wOvt/FTT3O6Tb6TfL08QSZme6brjNAzn6
+sfrVn1jFQ+uTIktKN7n7Hb3vFJx844+Xxjyaksqh3xLpuZTMasrIhaHzTrSlGPn
aYjY23/TYRt6Jc+ptzLS6sSaEecaruGUBixoNIvVgF4Pu/Mq2LudlXdGqbJEEvvn
N2+pJ7ac2K0VIkPvalXC0dPJqLerpdnlAQFIUUeKXxVUfJpsvFkeWnl+zj6Y+7Zr
zUbnezsqNopscNwYijcyBr7fuFgjq5lKs3JAbrPzcy0j/6WMlCmfjSLS/DwPgurU
Nb8CUWxe2FeswyX7weLbjdzBDBhpHxs1Q+Y6gP5Sh3WmWZHDE03t5aRimsaLP0MG
OilvM+mIIV7J8Nla//dHMp+12GEVQgOp9Ug+/h6Unos876gDbWBBrMBpGFirGtRX
bdZNiejwYDUzRmWDLAQrUS1UdesieG4Dj43lDAv76qQb6Cyr6uj4JZckkaFBgwAO
YjU7MMU9GTBMe+OSHpkWtaCbYJlAMJLxUZo2wo8a5HBQmwZR2JT7VGfiB9SwTWAf
r2aNbzEf5IUcmif4R40Fxf9gur7ZRIbJDSPA+y14AKEtWsi1/gHWn6MdlcwHUXBa
AbKS+CioJrBSavKauNYftS7c8M5VVUKLPaEC0MCpDoJj8WE1fVMpyvH2h9iS+iYY
AqMKbykuP1y1Ub0Y4iWNvqEPpjvdSi1vRdIrj59WpS0U7FeX61tfb4IokinPixoU
JlZ9ZWhw/09IXFVx0goQ+b3FPO4kNIuD3ISFsbgmBqSKb0HWmaL8cgzEMTTtLS6E
Qtp3vmNTEgRrd9ZJDCvGc+n/IDGD8kCQZ8gDM18ffAZDRPg5CGy7sf54sAtn8pXk
6w/EneQw/dScqRX2B3hMC0khch06WU0sbV6zZ4aCRLV4ujEyacD/iqQ84ckHl5Jc
daYq0cujy7AFpu4MynS8rm+luAgwatOU04kICZBMgavhzJrE8VN2FXWF7DL5iGCn
brf3iDcQUbuz5C2ByXW6mhHZj+2KEbiIkGLED9jfCogiM1ZPcfq0XSeFy/Llv84a
hpGUmJ7HAEOt9Ow/8r5GnbyByT5mk6cmceFo9AIrMpdfH7ptLmHp2j+QOWV0e8m9
fime78x7A4uqI9SC0n3aq3UtKCgIOB9lwWsb3XA2L2JNs6Ps6fgQ9i2pAkwAcUWd
DNOoL50N+EZEFp4wqas28S53CfYllT1NQC98kaSAiD+iQHtfyRqcavK4qbNrUBd7
c7ibpM4wZN9/Z/zubrOszVZ132aFO26aqqRVfzthu21dBInW51c3vO3iJttjnkbG
KzkzwHajT6JVB9h9elPKCjcAT4J3T7sUoqJWz4mljxCN1Apd+nuiCD8gjTjqPWYm
GHwxGzHGs5woYkWi57v4iX6/y3RRiA3bDg5/Yfnj2J1n+4KM6IlfLRko3brYfLcx
Ctckuo1O7XI4bM8IA1hmS/GGs6zt84L9eeFHW1CuXXeq+zo/GoWgIP/dHrxVt0m3
hnq/SeJQdvB/D0QjuiVcONOftwg/S9XKuEmpcuDb6nqilwoQjXW/U865zIL8U6z3
JMKmpUGD3C3+nv5gyBgKfETA/1Zg3r6JENDPdJQONRwmONlDN+TPnhQAU45D2AeX
Ifqff4Ef/tlwXHOQ4XvHJUIos/grGmLNNwMAvqJwE1TyIM0zZnfHAuOpTJda4W9Z
uO1gdej2cJHZR/IwP5BzZkm7ooKDuN+WxNSWvdn9zN8y20XVFzU0q80di4MMhzek
vyCcMuvobpEKO/whmlVp48N4/Xh5DRtFxXm9Etp5n7Pt0SNBRzeRbwX0oVlc7MMh
LuWVBV5jBkB+oKBtigIGiLdD4Q/UbLesL0fQVCZ2WVLrco3qY5A8rYEMwkUBdoa+
vu6E4Ii+uiIeZAiS15lsjAw+T9udSul6UB/qbAZ62a6AxoQI2nO+4ZUXGWbu7weB
skmxT8lbeuPyq81dxfpQkSElimEWuvkGov+55gFv2hSS8JKIbKHNrZFJNf6U0gig
lbg29roJOaAuktn+YLWm9ZfuPsy+CyAmfDBPLH2hK/xrDMR7FVI0Sg0BnvPvyxEO
IeS0ZnY5wpX27UlFdM44uAHrQGAI1j/9fditsD+wxfFnLBHMqZhKchBBed0w0smk
eTxELiQKu7Ec6lq2Gr7SQWuV/xQZFc5ZfWu2U8Scc65GfyiZJO5DzfAIMH1FrsgI
XG+supKV9oO4SNR0EE3nLlUMi9xx0/Ob1Sv+7l7NINfioJyjmGmdiGvzt7i9gm14
ajNPPmeLOay/X6T4R76E0cztuzZBcVsCBCUSyZR8U6zA89Tm3WnuqUVuvb2WEq5c
VrwBAcsVag12dkWNdCLqR7AwGkC8yxVTAs9pptmthpxaabqRvpHm5ajPWHSr+UfM
YWPtkI4JnLQkP5qemwctdA9KD5fcgVq7TuuSUWPJrHzf0MhgXfxqjoyN4C3DnlZQ
DE5yZ2GKX02YNuQLn08MrsZGTseBf6ITfx9CbL6GgflZe+WnQNMGutvFKeIV9JhL
M8dPdEaIrfl5rqYiIzGsb/mtMRwlyvcl/WluQt4AMOLtx3BxIp9Vrc7i9G4+s4lQ
30iMa953wjnZ1e8s0+0mhIuEOdgaKjxCFGSLcgwlLXc1Ft2rH5ehgEo5BRuunNZL
9hB+RxIcqQYHSLv2aU4aKllKpxWe/6atdkuf2t1UtTI3EyBLdZT+hmL9d3lqq0f8
GZqYc8oM00fAH7Z9/Vuv5lx9H65NZb3CW0dwAPb9VNdnr+nmctjE54JmaJxk9shZ
hI3d8AGXWwGqeh1leX8Ep7H0ncvOEgFt+oDdvdi4Zd6qAfyJ5+xiDlXShSjuzWi4
4eZtZNT0WUIl7wWIaa80vqh/r43xmNWIiTWWL99PeeErE969tqCAkE7qocLgNCGc
jgmIzjOrYRmp0Xrow8x8uY7WRTNTiXOqFiriUDA8I9PgQnSLDSaBw++jeZyGE3R5
Yg3JfA+QR1m1DPTLcoo4CYveUuq6soiV6IYsr51uYGc0vki9424m998z/vK3KS0J
6TSrxYVbWxh0YgUVpQo/RtpCCfxV5ebim4pc7p0TgH3WlM0wEa8o8ND3Im8bohj7
3QSfetWvxdvVvIOZb3B2IsNAegxb/lLMHlDwfWpOvmh1eMckRKHF8B1Cqg0TcCNT
nQ7UsnbN0gRW9aZ1rb5GuNvk+Mhoss+33J6723G8AoQI8O/Fh3JoNodpoJ9e1gNI
p0qbOzOav2lEBiEj92l/tq0pyTJgGBEljeeUsE9foJe+1SyylIdag1xa9JB99BE1
1Ow003/UZ/EHTxMW/+hzeDNgVuelhUqPex0HuRewCJ745nMF5cAOmgN0d2P16185
hhUhCriLtyqcNEy7W0+QSF8trvwPdYV5g1BgoEnu6V8au8epkT3AN4AvWACraX9E
2LUD76p/DeN/5SzxqyxrjcLwqQ18gKPEb8FrodsllI7UqneHWsuew+m7GF00cWri
OCYE9SbavYi4Z9DQGNoeyUA1Jcs8SCZ9q0vpF6HzEcsHAHP5Dnj4yfMrnLmwiiEp
VZgcIDOw7QKBPkB2GkRilpCfdKdjiZDn8+ELzad67/RDs/kjvBnbR+pstFfkh1iK
3lWAmdFKDEhToVdigPGS652ZGTOhKTh7l1g/EEscktbd4wA30Qel7v8BVFvjvgOK
5WuZJKVBeaZcfI5AkE1VMKHCBzODkvvwsgNJpMAYK77aB17bxVtVJz+5pYllWj7N
YM4SxwYOgoI7PsKd60GSPiHI94TeQDoE41FHnFSqUhGZtpnvmPkVSx8WKyRXkGjD
oEjK6/AARJi8dKUewE+IgCzaVINCmNs79b5f9iTF7D+aY4zGmxpH7cf5U3YWC+Yj
rlNhunLVSgj4DquFrF0CD9I5b2+BLtf9a1uHEkk+W1CeSFBrOO5vrPywSn0Yragi
16ikUtjtx7YPnym+vNWXSUOWHrt+P99JkYA0gCw45AlSWoJ958/ByQ9CXLTFAQK2
cgRElsRIyw/ZizJhU/bAMIyY9ofn187+FoUqtMBvR1t/MX7kyFcr3BP/8LTD858t
GDjY5balbxW4OD95ryeQ471k0TzrUM4Vl3cjUvhIi7K0H+Ni5Js02wgZUyDXwEI5
jPM6+ahiojQEbq2euUcGEvYRRjUvmwYwkJVU9QjyyhifW16+i0lVKTp7DYdaAaPQ
ZhhhiZ7MT8MjGL8J3vA8/FbJrGQxWonvsxXa/FqoUeBnZwa7LTkAtCTxi4a1RZv3
heRPSnjCoxW6n8bA4B8OQdVHc3EB1OK2cefP5sYaw+QKiIOq2BUpvBzcujx7h6w0
pXmoNLB6/xHkhdtGohfdaER0SUsGBo+5PR936wybsmafqtV+lhzBzn00nWFbx+Tj
ABqZGN7cqWz2FtDf95oHdA+Ulnr/8M/GOHcDO0IEmPVy6SieM60gvbtnkDtUUA5F
bK1XOZXn/EeDgtrE3xsELiXCQWpKuJ+7Mff/fjn2UjKPhnlvhOR8DuIDb3Brp4oA
riQ5COhbm3ZOd+LMWhjdoMb/m6/CL0JvpiTYUNv8hak1m5uYO80lk434uTBiYF7J
GZv7Rn3/8xV9dtQZJVuU5u2VgLALv3CgrK7zNbUZhnGPfJa39oqq5/7xX5uNfbgJ
P62B+CRy3tbqzQ1y1ADFyDBE0jp9Pz+ilNT6cWRC6pDMk8KxxWs/3WXgeuwl92fh
D5aJ8dtcbZbI1i/Im7893t8rlSsz20zBmR3Pq0b4VqSWheapgepnL2/SSFTB8s00
jUHrikeZhJv5l450UoDhsWBCT1/rW+X/hhqXIlu9C5izVxAGyka6xlmX7nmTscs0
Pzwlpo/zQinWjRMKG9mOaRiBCfpm/mNzCeEOOsAjo5ki20lcq+WLWXJ1GvEOWGe8
D7z4lUTs4YhygZxTHDoEdI1rztT+g9XiGa/ucGh+5x/i7puzTFXY5YK0fLAtuXQA
FWoY+xtNqud69HknN/9ueX1lQaJ8beh4xRydRIADbwIuKCc2jarr++cTM2dvl5kH
Z4a0EvDtKtHbCGL6iCKjklXGfuUNnn7WulvsogsWHT7jguvGdYQCgTPc5/r1iD/q
VX4VG1/ZgxvrsdE1pQxM15zbmsw9tSTBSqPhPrsHaIeNGQbFNZdXhl1z6aEGE28r
YLpdlBxi/58H2DNPyhFKsXmw7VS2nIqZ8/ASIWhwUYZ4Z8EpjGadinmEu/rMGqx7
UvU0e+AfPt9PnbPPf5nYTrk6SVr1ZrlJLJMRS9JdnZsVphjaFmVsM/ODARvu+w+3
WhPrdOe1JdA5oQcxv9zQ5hliuuhzcW69Zk6sm6e3bAOUmIncPAblCQykkfHJzpSb
ROLh/9R/WrrQjWvklxFQFQcMRpNrmbMTrRPBy72cW78W45J/pxxTk5JDza/QkTJ2
h9w49l9bUBG7Tee0JQFJtjYLoXWw2d4UWX62av22XhKS4ecwBYRCZwAu6+0mVNVM
acQ2+K8yrZvqJbqo1ZBsKWtdzZKA+IPeYfa080oYt6aVMNhbiMbByG3TOLyf6Pej
fdiHAHbarYzuLNFXMZ37XQ0sjemcZncosP6jT65lOmDCtTYYUc0T3xDrDvX6dbkW
nvM+75V6mqymzqGubJESrWxUgLdN1WfZ5uSrCix6kIQ9X+nx6Y+7xklrU3yxXvxM
XGxZl9jR3LxR2AirnIh5EJUdHBBXvwdKBIMLfZD8JXL/kZ0EpuTuXLUG9JCdCFWD
XvWUbAeR01DdntCuVtSFfPc10QxxOByzaa6rnhgkZw9MYl+e0R9Fmm0x6QHJq63/
niFzhtplMqJgW8Zl8vugBbQXZGrwl43c+i+fuGJ8OMns0sGp4pUR0fLJVZsStzNb
GbdcgP257IQ62zErPeXBn9K5ilP/l0rrXjEncZc5dF9L80VcPYSIzIx9D670HLGm
Hvw8s5LrXwddbiLI9Ix9vI3vlQTkxYMrQvJeAzRspbFT+7/9Zkto5G7ewo5u+cnL
VPtRSqPmyF/jc5BNX63ZcrG/ZbciwMwcqmco8LCZDBFxxrGE1adDFOZkjoGKe2A8
zmJcCW/182+34TpNoHSymI89rj6aYEd9kf5yxjelb/DP6/qwOlcQnidA/6UV/oFz
caEGI43nqH64OFDoM3QS+YWwzVTkcThZMuAq6ywsP09c9UOM61cvIJcLxELu2TrL
EWC7oFHuouxwx3uIw1E056oD/iHDWzMSNO7rM0ny+MXtW31XHC4o/QQYhLL6ixuR
3biZ+LhySUiECQaHgqo57NYjFBYrSK3MzODZFkCFQXrR4Fc7ZvjUrpUgPCmQAE43
HHy4rmhDkb+UX6wSAD2Q2NTqF3qW2BEv6wrz3QCUi0yDtaV87hF+7VfLGMg+sxcp
pwyRcxa2N0NfPwW7y2Jb3ifqw3CuyiUltouibVAeefVUxanb5jWTL2L5MM4c9kqa
Nm9rlqvTk2uZNYGu5vzkXV/jDOzgcAlDedVy+viQKtMmo5rI9+lD1uE1FOaEoU5F
dScMDzOapj9+8wlKiEiNpqN8Rg3yhIH2WAIHROhaM8EgACbBu1ChHjrJm1L3nvGy
KN27DmohCUXULyDB+FqBAwUyIyNP+FJjz+V2+35HYYeHtSl+E00DUnJsecPPslOK
TWIvRdVcARDRaCXZZCbEdUe3RmmE8YqPxP8fnHCfV1UIADaoLYkWba3fra77Eu9H
R5JRIiPzTEtu+mLWZw/ncz7mCJTsiXyNPGELE9gSl4fZmUIBLLxq0oLM+ujjJ6nc
TCBZrxN4NkvCETNIULieZ751dd0y2aqSFySY/KDE/CUwyg3xXx9oGn/gIvjAdvz5
FtrT2HH53FBe3pmwi5tHTA/4PLMWAGt4Cc4Psn74o29gRamSrHQVSaozQOsGOYOx
pPuZEuyTUXmBcaSLVfIR+WwMFLhQoGjYKfFAqTZ3MIrz/wHx9ZyxnMqlpzt6Bj43
FZK3N6J0vkiTuFZtBLQOudPcjLkyvMqlgQidlXX45yW8SQdFjPPOWyejiK1tuIWn
U5WSCuRZMY1xl1E/W0h5SIvVM3TML3C2lIjVS0ZIrwQ24EiEp7dQ9mGoi9ofYevo
58RN3jD8eI6CNBf4/N7s6k7SOnzgA1uFX/jVGihKmnQ0V++JPWr+UuU7sxttWV1U
a1wPc0xnaX7pbrcyVbu7WEUgEbsM9aB3ouIbbRl/tck2yIk66Hun0DrMv1pCz7GN
VIzzE6K27OhtPkUcm4Vnag/gMh9IcdCb6PL2z/FfvuJ7g4JR5ozpuVNOy2Gf01Oa
xQSy8/E8iZshcvoyf5DTrK9HzytAJWrrUpOg7sj9qXXLbMEhrxhNPmL01eNv7LWN
7fDbRC97uzOY4sHaELXZVyUVwYD8+AImvbGfGBr1S5azZvMy0juOac9QHLl6WIBC
UVE6QW+8M2bNGTyBGb/FN3SdqycXzGdnewov/FYNyG25FTWq4MonC09yql4tzFde
sW5GfOFzY5fmYZ667iukORuRYmQGFIWoHH+OaswpP3/kHkp2wtpym3ReZy3B0INY
2Qzcwr8uOU+Lfysx0ldMRZRSbtULFF8+xaErBgfMmqZR+U/zqO3ZKqH5Y4ztHZrg
t8RgUn3LZI85wKT6Z7qgCBaABLtTDhYCh5d5FlGo9vNcc3Mdv4hX6EVEiBrnti+f
pToLWaWe7bWRoDByq9nrDlanQ6Gc0BevcXF+VtrGL7jPyrX6Fh/mP3LawIOk0cgK
r0P813Z2hHNRdvJiYiGZp4XrpdgKzswj9IvyM8Sh1MKPcYc5GyHcRwLldE7bKTZo
+OgaWt7BVtySyg2JelDT7QXUqR5qK7bzXJSljUXpH9lLSuUFqPSzQNMzE1YGKGCo
GGnjAuldosG3+g6MMG1WSLBUXdL56shRbE9LVYlyPGOF8O+wVYQZeq9kaR2OC6+J
OHBQk6wWaX8RBVvYic0Pa0/aPSszFJvQJX7lW6s3ZUspRTnGG/59kTT1geYs3W1R
9eGAQ2kZe1k8S6LZBWkFNi6f23q0W2Ik4auLwOGKjEfcRbylWb4gh4z9Rq/0PQgy
d53i1M+keYa0gl/hLR/4EsZ+jKXWzefrorRHUJmgPaQbpME8EzOQByDv7MIwdw+s
b1Z5SKMZKIGZ+FUFRA/i9+kSIRbE27GxHn67TJeVAPtI4ytobjA97MMhhVSvNBMh
r2eQy0hXtfwLgO8OuSgqYXt9S/ZqbiNfd8s8t6I0SdMojoBRX/+gKDAEFnlFSGRh
xXDDwVKqC1IQv/kig8b1pDS7JlO8D8k/TAgBZ1DBr1qb17ITsTa9bBbn3ucttBR9
mbvwpVZL65ymkCTV7ZD3DyJiGwm/8pFmo0Ze/lA2pSO75Ci/NZBUtkdPXhc8ZA3Z
NY0CnLSGiktpdh8uixmCJLilu2RTbPMTZPU3XCUeFtGQYaGe+xw4fRgVbyp9VJb7
KUdmupTTYaSFiyzkWmi8dFA3XEHByu0geBSuOXGIDOh7IdBUXptzIao1G/OnoEal
DEWN3LB6gpNAKvAA8CLe1lgV8cZn6h0WFutKexVnf9UjB9+rBrTqtpRbw7FDUxSN
vCUYxiT+aadFaNr3Le1lQPLwZoO2u7+llCcb8qgoNTv5IfvBfC6VarG8IJtjsw9h
ag64ptAw2+qpeMz6Mnxz/I+yuy1jMtDfGJqSYLdf1dbpc2z5dRNWDtalJ9En0MFT
RX8EaXAJAmXHs0YK9ykADaLAhk3k7qNyYiJPYlskBdqCw1XquN3EUzkL+KGCdSnn
F4OTyW2CcnnHrm5axw8hWye+6zg4xqqSqh48E4LuQRPNvKECn7tpUHZwatqbkFDy
KlEQI9Ox652hj17PXMtF+o+5rqG5RAmu5KuK7MFD3Fd3E0T17Svlu5m1ZaWA4S51
fYbtRC+95O2UO7wS7IWXvb0mn5Werwd2poWAIM9xpSaLxJQlw4vLyvHuVIZjxHMB
kCvvJJpImAvknZscNXCbGncaK1iEGlH0TTdjOSJZLIg3dtxOBOsMbKpdKopOzvrp
jvk4oDpi2bH7UkMOSq4+F0FEShHPFXVtGFTUgAJmKR8PKm6/js0FI6Iv6ewMamDv
KuGF2fVv+New0B7l64hTUCN0o3tyIXx/qJmCZ0LWkoDmmNO9yknMfCXiRIcEFWc6
9d8rhWU2LQqKUwR9xWT4YOo5soNj1r4MDuNB6ecMDKYUutx9unyfYm3MiYmWWowX
MnexqkAH6J4U+WVCbP9YVuZ1inLK9Ie8geVu53Do8S9KSLGLsc/6FXZXDCYSJuvB
0E3Dp8qOfGYDVmxv6Oa/I0yXejgqhj7Ac8o+GP/6C6HYfQz2g67Bo+ggjUotZPXd
TRIJ+u1Bl83c2Jc0xCuhLTbCrgNzO3yNXf81WOjcp4dYTAbZhHBOpXdVnxictjGe
x/ox2Qt2TcUhPpL2mLcm8osqKhqVknrcGj2ct7YNocPzSXgluMVbr/9oDDVND/fq
VQoRXmIiCftlMkGhbWr2j/1ScoXPHdq/eB7L8m0z3xkHJf7r5XgxAWL8jcYFvWn3
I5VGUwR5InSacoVrUBf90Jx0vWOqszrqOc/WfdIWaiyoLgRB+022vhqSaVyapAqt
Zb8TgCDua9gjSz0VMtZjpw6x+VUEWBcPMIs48pVRmfcG2y89BxkbHYoDjol99GCz
/qSdA218CLb2d7vXxsYO7GABfiJ89/iOZNPIHrzVxFcIh5CqbcYiw8Ml02L26a8B
0WY+7Hb6YmHTdtiocdrX2O2K1Y+5CiE1XSlyLtpJbXl+2Q2pc2nwd5GCSuOu7gfg
nkdmczoOceteVCiz2t/+9YhM3TJCNTKmDyrW5iJ1KLX+GBNX+YhkEWd+5FvettyA
tOgb4s9mCgnNIAf0MHtZzPDZHnDzAuPctRRJ9Lle0k1OZ0Rb3L+M6icy1/uAegTd
rGmBT5hNaNtULKmpBP1CoIGmgNRD6LQ3vNMluRqwX6pS7TZf0jb3xWwJGvSDcXNo
0CK3hnilXRa6OK58rPpg6h3W+1bqKKUZjCUfSyRdOMKZk73bwO8L+7rA1R0QGzaG
JOsna/oqBljLh72osWWPTZQkkClKkyIZXngf6ljbic5lId9MQhF8ZVqe2eiWZV2q
b5vCy9BD7nO3zYsboilh5UXhQOhqrhlT+hEQ+u/mBzkk6gGhkDHVpIygyWK3EOCp
aTA7UOFwykUmOkqa7unaYUkGzFSWFCOJ0T9HjTp+UQrCB70CFL6SJtopWyreOhVR
COhWK/miOFogcjYm1t0YMXtYm7d+QpX1VG+SE+u1HnyEZFKPrLf0eXBtIA43eQOG
H3TgZJNKLIArqa5cskQEMyySatfah+XqBHjpM+6/oIHs1WSbswdHqmx4y0nuwHHK
Q0/xPFJyWF557d57WS2lxFQqoVQ2VaD/n8yE7tZQYHopzddSN9mwXrbPIJ2AlO4G
B5OU4aOA35PmT+Srfv2SeAgEmjUKrLNQSJXt69iKzMj1D3Lb3RXK06+faJJ77uxm
dreBkkgDEgpQKnHG8I89gDWdBWS3pqWrd9H12UYYuw6Q+vpf/wwcFWOd6tPlZ25p
c50ZBnX00RSBtVoJt2PcZo8mMyZ5Zaavr5g1td0Unn0LwyAf6ZerC+s2Mh6fxQu5
jVPY7MmkJ88OrS6alhP0aqB47m4/0UEXFdIC04IfUp3xzTEJeTlkCxiUwV2fELSu
IL6N3unrxZ0ND4ejs52gX7pnpjG18bqjArR2b1E6VSRmWThM44WyqCEAC5Aie+kG
lx1ydQr2kLHrcaWAN12GHw/0DmVmCEFxv6JkRfTURqp0CVrzNHoEZqnDXMnKATCK
2obmsSZuK8XT0SEHZrAREuejGF531rkwdGS/+Y7v7F3l7KMMjQgZNWZl7/TpORyP
I8sNpHfaqgikR+qfoXZ1Xlc7zB+EEUtmmB2njHAfLgV6n7Drq54C/rIOlMFMob8H
MU5ZWkFPIt8kRRarJsqDKtBK0+ccJLVs6fF91HZcO21ljxAmZ+A8ug42N5QfdrZI
zTheOHBIH/r7PQsQS/KNoVd8VCJtBt32bawoSlXGnEbnrKPIbVgX3gLeGYoTDVr3
MRfVOBSZ+OAm0Jfmof9MCg/VykaT0UiqCkZTuj52+ct6OXmDeezLJmosRme3hhKd
7AUzF4bTcOEluwFERfVSALxQjjTac0bJdgikpXriy4tdIztOR8BYQxjrmJEOIo/o
S5O7CyKSlWd65jeK3Qlb4BjbfVXtopnUUmH0S3QluAKWTeQ4ruHzkOFjpFH5KEK4
9EiZEKP1L7yAIORvw/QdQKqAlp2tPm0I4vQQHQ0EMST1GHk3ULFzfYVIctZ5vmqX
FfAulAED+pTrG4XhB8LdtctViKIQOYRadnO6D8gdCvvDv83L3OwvJ15WFwPGcU3S
7YzX/TpCmHt0Etm6Xjnv181UdhSPqS9Axzg17mFSx1o3fBU1R+n8aLwkoVFgFiDi
hiIB8RJQZ2HRfYipePZ0+/SdWRNimsfHdeYx6NTGv9DXCZLonAb42ibNDpuBCMCe
49C+pCrSrFEihlW+SkdIl1LFqa76qh0cPoT3JbZC1wgjacXDVirGKrL6TE3f6BYh
ht8pT8Q/lEUeK9kPVGuEGfi/87DTmSL099DaH+fF8Hd8Q1NTd8DpjgSGLQtMmAoE
pkXdj82jiTm/BntCL13lzMq4MOZoylUghc7pAabmAORPismL0l44CsidBdJD8EMw
ekWngqfPOzMXVYGHhGK/YZBpv6xngs/p7QXL4Tlh7d970ovFboFtgKIKg2MQ/mGm
+o6stjG7IaLnjcaUuSCBioKLD2WWKsCo8dxUPmL0tBgDEmTX8/3Zls7K2Q74veM1
ZfnKVkVUXFe5nYyJRAm41/4n7pCZhr/IzJChCysDyL1a4oB2ogzbjJvd7hZYFDL5
0AJBDgS7i8lCvcg4sUDi3H013eC9wwPFNHhoBSHTtYbSe3crvXfr+YZfOWtvMrj+
3U4bqTTQUdCNEYyheRcZPBEhbt+kFjlhsWg+bNOhXTRKZfg7ba5bbIh+dLdyFYNw
J0t4kP3NWiad2QBlb5Gb5VBG9bABirvNn9Dh8RIUWPnxJSO5hQ+qu0FOyTawnFlK
lRbpoDwONYRHLxVvHlFY5ZoSD7qsZt+HM7g2vevTICPVZhKbMOwiYXogYHR4uCT2
w1WJYtb+RpCvX0Nuh3y9epE08t725Mct7R6LOYcLU4VkC35rCqOOtlAU4enR3/i6
1ChJqH0tnZwrpFA3pzXxFcHQhpkehUjuk36uLVY20u5DdbQaSJteJJ5tZyUUpkxG
H0Itl0BnU1jogRCergPryvpSRBH9YlRFvPQhjfjyVilVfkoUCo6Wpofu2WeILk+G
ePxxOZahwOQ3JatUv3HJSwx774gblouQKlBAfygCcvucnmjq59ejjze7sUOCRCTs
MtwW3msNoY47PsIA4VAyNpEeqUsZ6GsSRrBo5eXvZQo4T4ozukkPQ9oBgmOouzIS
MOjxk/60txU4e6+yAPKX8P5Ip/jvPRzBt+olCx0l8tY1PyIoI608/0XT/wrD+dPy
/+OT5m+oYVwLS4C+P58PMwhjANfpMU3zXbpjTYbltfgx0nCQrcWzU5mzvChxa8VP
rRx7sXSc/WJkWAgEULRaf/HVgl3EweyFJhsEw9SfhkRpnTJ2oY6ys1hOkBMJpnVT
GgidSJIpSow6aXX1d+taz4gTnXmTQAgPGuKsGbUDZuDpCcutoiUuxHa8snPvrCyf
CIAlZNKiYe6kYRHwXJD6uWfDwD2qnznhVqcBn1pua0FEVNlp4+40COrReWzEox37
ujGDmKLvgOncXUuQ+/kBmnCwgQIfs0UbLTdyols5MooRQoXQUqieolE0L0pZ2tAc
4SA38zRr4a/oelBLqa/GpsRQY1BnLnhMzpQn9Uirj1ItiRR2kEPV6IAcd6JfqyAc
eTNknP3/nmSawTOsKO2F0YP3wqIkR7aefJTQrWUVmv66xfOgqbGIMe4tFRzw/D3O
A7FJwL9sujpHcueo/8YNFdLio6Sihi54eEQolkKUnvXzO7VPVtez4bTJAPah6sCb
YKtmqJLFHv0CfwKoHNzPILY9/k2ifNjWZaCbHJPFJ5T2e697E8zL/8weR1C98ELh
5o9YE7CWbIsY9erVLCKONXBsWlCGRI2vKvmO+Wgr92wA3ymSu4WBGI8q/yG8gpra
/+egzhNHpmob0ULA6lxnM3cSZ/P/p0h0tS7m/v3MUu3EB4BWL7zFlP2J6wM0lHnb
9Q/LLNenNQ1P+sGJNfAzZybP5FuPTB4sEqgBhJOzOWBl3lKRIwsRIIWpelFL8hp9
VEov0jzz/4rNoTb/m3IwRkiWKTCOjmVVZ1S7sqtByPVElY7zIH4sVKBWt0PuPXhR
Klq6e2RIuVgMw11W2M2HbgxLpDnQuoWFv1Ap7Uu2n/rb7yx3It65jJUtI+WJZuVk
leDeWnT0l6A9+SiLgy/+jVHdLrV3zje8EAyvrZId01SapTmV7kQ8rwirbASIlvX0
oHDRiP45zW/bflW/7PIrHTJBhkGsEu698QB6BC9X8SNx594oa22NgewRqwq1JudM
xw6fG3nxGStFNweoCIWfiIaKIqKBRhtc5Qrt4aoe8CL5iCOZ/ncVBsVq2YVFE3E9
7tYIgvvqdqI+NYDkIQTAtJoWUK5ScgN+awAmMbxr04RxnbrkUc6a3hzAV1siY+8K
Txe4zz7o6tBtvC5uiLt6F6hbsFqUeWPRWi0Dkm5q30AcWHEVrhFSNmS9dD+H0fAx
4J2ATaQTZ0je2d97akuBtL7mSnOF1yODaZRjWVv6Y7TkKn/Qcw5wieOnoMkPi7UQ
XC2A+4uWvQbio13UuzzoOCy4c+Q54bf/BHaYmZOQYqwto8l2FYveQnGbbzAcAkDd
hPifNhZMtzfsVAg7CYsRc5chb8zB5ptCyKuYiH/un9hc8XN+De0U/1Uj46KHKmtC
0b4PH1Nj3muUPDu7ViBmEloWVWKSHIa7mVLjaqMK7VKcuo+goFEz8CW9bewePS0f
M2R8nGk8r+xYHZQiRGDln0UVHHzQRRYhr9E7DrMspMooaZgW/jvxcdPw2BGBW2CR
VU43xd1dF0By2A6mLHI7AQBdGLJCkC2NHGnEmH/uhLxQ+H/dRqroRT8UNUDH5Mgk
4wW7h28b+X4kVNTPii7d5z7UQ1Bwbj59YS1v+1KWso/LX91WOfBYMzLPoRQTt4uQ
tCwARLLS2q713jxUagSRj9/yJjSLIgh4sZP7E4tTVIVB38GYSvqNR5gxiI7EiloN
IYPMaPfBtJtBB4h/bt98ZjXleMP/HoQ/zXEa3NpqhnfgVzKQ/uK223OeHM5uauKg
c2ayXBnbk4y6BrYqWZ57Hf94qjyCiWjK6YJ1MosvnvVeG9n78675zV/JFLpc3eCR
lZ9oNqu+VkgxzrPVfm/8z234TsoyjzwwuIzfbptjVQbqnBLmYwtlr16O3uPlECTB
w01Iz7ghgQbCTpjL9Ljulomcrd6c0mY3XBCIY7gwtiHMVTf9DXQN0x85UvpqwVpX
WoJ/xrsgG6XYjUmrBmo0UMbElFLalD6MBve1uaRgFJfKbBrh31IEGcuaWw46g6Hn
4RXRyoKOpRiTFB+KhCebgGQl5rnMDGxLG6pVanDh7piei7bZ0+SYILiRnvMV5vc0
xcS/jg/MWrU0kbiDOffipEuEF6QKn3FVyMfHi+Szqdfz1bA/5DUq/i7B0t7PO+rW
4gkjEnCKfe9IHJEg1G2XEMYV07bHZsKDzurjOM1nrzJHbhrzp5ZXaFHk3lK2BYJn
r+BuuPFCbCKvGbM5YWEhuDe3q1NtqMmfEGKzBr2XNnWmsoPGiXWrdURN1R370y2C
eMG33TU5kDm7rdEzWXEXKPY9IEvhBaU439sHH0azGJBfsHLB7prl4DtJrVqiY/w4
4BoHgNFChaeMyjCYT+7R7iIutUEqyAq5aeceGqv5NvsKcPHZ0zJFOWSoFg4YA28s
DuwtcoFUSrPta2KjZvO58kv0EVVxRv2cG3CNrVMHmfE1vEDhrTdEM7VoB0ccePvu
Xj3WKauduoFqtzEnlBxGrN9nhPE/KwcYc43IRUcuN+M0Uve+lwMvHDOUfQWE+SME
X3cx7GEByq7LZF5DGmljcXFaEHTJVcxstLOgnUhUA3WQRPeFijJXicTG62UY3G0n
nzzltsrilgxUuN3ywF8DW722DQNOPwqGAec87JVHGZQRCC64K1SIPY4GgE/PL/XA
G0X7PdwQFsmhnHz5Z6k//f/Ypw0fUngZhMmhCLjLjyJom/W6Joia+ZZyEpJghzKY
l905LQGNfsChtdIJyvAl1Ee8sRBH6ZlRWSCW8ZAZQxvObu1g+US+NNjmQVLQmaGi
Afq73IfV8dMoGWGGRnbUfSETbN3RCvfOYXPXCRg+hSdq18kK9dYPgnxgFvZWfNBM
+i6hAlp7VhRu6Yit4rXgtPjTVQbUA7aB0LonU0wXz3zkwijwg5Ec7tG4rnY0pG9Q
yWc5t1HItcyilg1YPLZwqjswgIWeFINt3TRcgGEtZ5ycvxiLjhaVFFP0tq99qZMQ
xnXa52KskfHPFt44lvZrDYnQ7wqFwbu0vwYF8uuPpf8Xe5s9OTQ46RbsUaPxXeC8
YGYCQ6PE6oMdXRSyTFPsY/SoOkRSUNHeoomX/tXLUyIZ78JFtbTr3TfUzcO0l0aY
OfqIzq0t3p2++JFJ26BpJ/cUZqt/nhbbK7ri5h56YLvfvMW+KvDHOQ3g6tdTf4OE
CkJXDHK5vFn8LR6No3G8nGQLQdZ/ns9GT4OOlH2mnrtAveMlQuU8HFQWHBzZrzjA
/cvm5nqxGcnsppzzGjoR80j6Kfcl4d60X4dOR8vnV2+GbvaFqGckpMEDnW1zTB77
dFNXha26gdWCom21rsDS4/JmJ8QVM39XOhYVKI2vZwTnMuoIt06i5P48qS1hL2Qf
EuXeftkGlrti+jnXXx54LMiTSR38aXQC5pxId9XOhNlN9ZBp1pQIPIJ+DMYb1EC8
X6YvM7boUFMEa5yLE0yXottxbKozR0ixw0DMY66/5WY+WCCuOPe9+8aRw2vGvAQd
eR+ZQdy+7kuqu6QuOJPJmP9H8X08RH79CY19MvJt/eVGKA6hgA+sE3fAAh66/42I
4bkX1EY8lkCRDLqZ4IQdU8Hx/f5GeeZH/uP5wBkkDloWYjWUA497h7PUncsN1FSD
sSBVmQIMiSRwJ638sZKauSDpdnTbbFU+2rA4R6qd7FDh1dL2MUpjnPvSZ+WOmUM+
fj/hoOuyOI8TLRUfl1Q3eBiowwKaFHF2yA5A92btBmdscitJxjH14JH2a236o1cA
UUiZ74pXc42wgaTQ8LZ5Pi5quqil1w17vuhKkOSHC20iyLwyNnWKTbvNNFXYZ7xp
biRonYNSY/5IxoxKJKh4LAcfZeBiR1eG0qn4jeol95BaiBxJTAul6peb205f8stS
q57K91bcFQ94zteZ21TagtgmkKlOiUsyLdmNjGxVMDTOKzVf7Zq7igoOPzen2Bpa
TZ/raHjZM4kz1qRXZRNJFEGQwbQTdhFzRtnNV7kl3NTCrOoannZr1oxGyiRqnmBA
jwc6JDpQlCV7Dk8IB2xQtrBUvkjEqx+bDBxvjKkUEfnM82aGbg7OBm2QLU795901
JR1fbDhhtuM3aF0PebFo+KtUano4J4EoedhaeEog1vWeRFEzBAVGzNyvVkhH16Ia
Klop9FHw75LOgn3tr1PW2UKqJRyjSAXjL1T/8GASRz6WsY/Ca3F5F0vr/MVSmQ4l
LrmLtoH8oXzqcCItyWOUCkf4on7QEZBo7ABPgtQVJjGBpvtkig8J5/2Vr6wYz5GB
R/E+VhKEURxeXfTeFV73MMvbE7qe0Tq1UXAe146TmjRpICKhm9TgmdotUyjD3XuN
d8AWz7FzeJDDloUoNK4irhO4NkmSkGTtiMVwAX2mK+IdaNd6yegDeHYWipfBXTo/
d7l4bTmgD49mhlWlmO1k8KXd5LEMnEQw/cgGOP0ayk6Tzaffy5en4Yfnzl9glEAB
PyctrH1Y9ywF99vdORkqtiTWBYCCkRt99JC2LhIIXvuH+foUdeiaGkrfVD+vpe8/
wrq7eONEDbks0i2XONSvL+3K7/JgvL09U5/RGc3sbcvUBMKzrEU3caBJngEG2qSw
ZJV4oQNDq13wIzAfI6D7/53LIGLel3EtWlb9NSl7wf4jZeQwelXGD9JVzIw25z2t
wtQgsvoZSaq2JCyTpnApC+RGDG8FcmK1PVI673QDZJOfhWiGXIFuGepM28UmUZgH
X7Xza59omjTvkQuSJKD3EvFteEYjKbdmdBtH4kbdrm6cKaVmdYcV513gv7lxusyn
OWW77LD0Fp/t9yeUXrj8zrvxBfcDstrPJcfjoakbOqTSp/TOsAmUj6wxuz0iNHhP
vTXeclBBG/agQl7sgIxBm6672fjBlC55KHaBKCUIM1uSyqrLPMsRb6eIDnvn7zCr
BnHQKLo42wYAASqCsQCbtuUNOw44sMuHaM1LR7iyahMJpm6fisWgGIsZWQXKzBGA
fX1GdvzsX2YmWZBf61xg0if1ZumNIBXiw+W12jV/d6gOjmWC2StmFhTwc+lsO7Xl
Rf6lH0AMsghaoMrpmSmZxsSM2s9k2C7/7+87Nx3NVp4fWExV7SCLsmXjVNmo1JJM
vObD6h1ntHer4A28y6mPTi2Ty3LJENBxGFJMHI7MUpAamOWyHryDCDJ14sLjExpK
ZzK0Cp5Pqhr17W+UmGNCbu3a0uLYTIflaH330c8t9w/b7p0aAIYXqGDjLiHQYOqt
Ut4OxY8XQ4tXS/4RTJK9Qg0j86S35MLSOPOKkYlfmyqJ6sL0obUC2rbsoQsjPU4o
yMEwAyXwj2jsYR0XLhUi4cSclVlzSDuHbtc1PjUqUdX3Os4aW0uOwtWHuHgmyoCu
k353WNvlmq99egkaPvQdpb+VzrHp0rTGJAVU9FwDRtGbYid8AqGEdtbARaWeHCEk
XouiIcrBSfveegaKI3ZSQblEmZm6fn1Jx60BlwvSbMBiRrRFAUnpM+V360vfXOH2
On93kd0FcU28rFGp3Y0JOR+MNZ6tYvbDT00xgNkU/wkAyrq8WWsr4sEcWgG6J1yp
uSkBrohYvGvWYB0nw2zdJsNCsPU17jd8sBqVgYfQoyaVRah+u1xgEn4LIR2m6O1i
Z0gTGYZc7fiUo5gbDMgx6osyxIBuuCnTNkvWuu7ZhTCmXstX9ALW8TVaow4LLTFo
67S/0kdjQaHyAuVHvnNfdH0xlc9ve2frQFbpNPJXpEglRevh+YOr2z5ViwiWOQ8I
CVHwAsBx0pFeq4bVK81RIYwSTMJBaNr/JjctlCarNPcBEMzwpe7YG6bd/QXLlpMu
UvRkEKQSAVuSvzf+YSMd8iXY8MiCjA5cDgX9VQFsnR9MSEiItOp0P2iFrPr13eZg
pTG8XmkO5eBHDom0AonytqAKCHtqUc0Jy+yENQJd8kzevSfTIVbFwPwf2EMY2V25
Gon0I6jAlOt/xknAbTqmiXrrX92Q19CpypPI2GDPQyUgIF6ANw/0ooeLrhnkzgZx
+/nKWeWrRWrSmX4GvGi2NvqYdvBY4ntNPfyHEZIadF45wpAJJQBQZWyaaHLcd2Md
BizZcWvpp22gQ3YUMcZzx1cKnQ7ZHIIf8Qwq54e5t7DmTs1JdwsmAD6Uf01Djdqg
PHWAB3nkNT7sbOZmSsZnD7/hveoUnciRYHi1a1ABsu0V7OyzVCZC1RKdNQ+YtJIC
Zzcc+OaeP8CPKth3I25TAfKolbodnPezbIA4CJHxNubl//5eWnuhXYGcbXCIBLcM
cWrNF58/QXPikhFYh9Ct7yvHs1AVQYYfZrC7+mbgCzzFJjoobVimICwkZBhNQOSc
EVZhKHfu4qmnUz6aeYLDAIhULKNpXyxjz2gvUbsn03e/qsdgCa8ZpVR+BWAPxu/7
jeVwVsq/PBuXOlKYn8IuISGbe/tuIp1pWedrGB5Dta3BIMD0VqeSKyiCTElxxvJ4
9Ns6Ws6q+q2rdYW3iNr9TBkfaLaA9YSWBapmI23dITiH3ELn7CYij3o5dJuPrqcl
BnKoXCy0Ck/znVBl0zh/PXvCEQlKAI7wFd62sJxqEAIpk4XSi2eviDK9n8qDhyq/
d2D06M1dttzCBZM338jH1V8c8a538uuR8H5ChoktVlBAcB5HWYetmyMbvTFsIlvd
+9I57RQ7jYJvMtiOB8+h2mqkKadWemWidGJ9thDVDBmelaIGNd9oUoSXUc8SN9u4
I2GspWvQBEHU1TV3BBQiITvE13789OCoTnUnZP/+5RCena/gxWvz/AjuAo9etv3W
JaHzHLigSsZ1KMBiK4LPXKEEpFe/pr83lQEz4SlAkv03gxRy65u3Lw0ozXJCZhbr
s95tt7JKouz4JwX1x55ClPxas0vRmLzMM7rbgUcIyM1dDyfWv1M2S3FB//3AmRcp
mLFfBjMEdrPs+FsxBEeB10jKAd2qN7SG3TFoekLlwctNGjbp3k+CQAnSxniGfMYs
kVkpe9WaZs/plqC5vs0ACLGkHdFJMrMWol15+iq0npVBM6hc1DYq1x0+n5BK59uC
aKAtjEhRUeZ6wm35FluogXYmvH0HVpvNMPpywA+Cp6+r0RyZ3uGc14NtnAirMQX8
k1JmGQhZQJDzEUphxA9JsG09y3v+SnKx73zB9/q0H+s6HDoz//19aBAgPUGRmyGv
S3fuGWq5uLXfgw5KxWrwIdmQIypw+GAD/kcnDa+O9ZDqyePzybVxJvYcNKDMUAc5
YprN/lQnXy8IAGUJLecsZVOsHnIoo54FcYXP5ImwonooLBwIx2RJNUPx3WWKPfDA
BzrG31QZ9WvbN5yX8+1Z7defx7qgX4FHGmJ0MCL6WYTL4f8LrrZn5PKcgoM9bUuF
kGRllNueAnMNQZrdy+eGTVOqZQB3ZZ829r6OrPejOXpHYdQ2fl9r7sQLHNuzPwIx
57wfOcgqiHxkzjSxgUHJB2G8ttBxSV6h65hlpTHxFLWwctw+5fcBWLsKmUwnlumV
NplzYHeQdfjtsSqUa1tSVFMz7YejSkEEzz8pVkcs6X1i4TnRCBzhGA2JZcdsgqOb
zGN4wrpSwVRpJndrEZbYmpihrWdAvutsPFLI4Y3OJKn901NbTdq/sAyt5PmiEFjG
ps75+YER5tBKQiDGD9uDfB+SCmQhjOljkXRlI9Tm4IJvBzJ+4sTUmSFtRCspbEfu
qK76AW/5XnEYKn1mqSwliy+v8PwBKmIdypFTShCI/xixXPQIcJ5RmRwR07cWg3Qn
5JeeGAKqjHxLwAUZD81JOUJ0bOLZriNEfeMbukWAd+QPRXQ2yeoiScBl43TVQ2aa
YzQZvNX3EgLWSeF6shCzbIe1J4jw7/qb3dPurZwqHuHUoc/n3urT+6jt+DhbEVSV
WAmvKB4B3RBaaK5BSlq5j9UhS/HtOUpBuJ6QtKyQ5jJLT/1IB9NtMd79jYmCFAbb
11CR8Qd3JYYXDgClmSqcA3bReKvS5d+J4NMTf32bL/uiJXF8G8bd1Hav98CnAR8m
h2tXeqvWCTQPpC3w9e87eLOR8NCVhpWuy/S/V0V/vLN0sj4B+LUXXbEly+2sIz3F
buKz9yBFDunwvCVoCz/tdK8ZAAOYVfG7ct5EyW/Bie3AMAdn6jNoKPwoKmvWnRgi
sJgspNAUyCeIQIFAUnVJptHrQvVvOKqhpeResw9GsoHs8HbZP3LzTav9IsP89bnK
oit5gUsdiIT6itednCtHkpp7HJ28JYq2rQj+3kx95jYCTJBRG92Wx9HWH7SnbEkF
D79RjGnzyZL3rsv6NmyXTjdhVNXD/0u9Fko9KLeJ36YmX12xBjxjULs2kMlEjcDZ
By1gISYxwkUeljW0p0wVuXPB8SiUytTWk3rzvhsqmuwT/T+7Tgdv89S2fj4Wlt2N
bcnl3dPPS3nmsaARD9bca7DfSD5c135Udd335UPuzXZ2qNiFGhvBKUSig7Et0L+0
C/m0q1EiAcy2KaCSRBsUjE3kfU7Z/JxBkJ8zuHgzi49ewaZDyPxcRSLhGA8jlJRv
3PensdXh4hv/XUVktUpz4RDyxDy3VKeAwnadcsYoEGo14/LBtmMJTUT8lolkX0VL
6JzgBQ368W/8dbTSi/i4f4cGomY39p7Oe2TNWz5pwU50Ec4j9KWLWsCWg/z4hgTC
WAg2LLIGJ3qoaQ5N8eO0E+3Rl2PvlcEtZ0oHCVEXFrwW8sKDL73dyjJ5lhVyWQVh
5h6q1hWMWmRN7OGxJC2pHCjg0OVLvobPNk9a0x/HRMaDfQwUApumrTnqeOMcZAN/
NlnpMUw9Un1mMq3nCRYoLmUV8151haO2Si9v2uG+yVi1QEv7s9gLa+Jd1wkm8C22
d6nSnNFnDCP2aHDp1BfEcPhuBSdr8N6tFn2KMsLiw+d6/D2Yz3inrzEWEYEuJVue
p2XrBvUIfcYnlEhnr3iAB3upXFmzxMT+XgOu+0F0GCQp8zc0dhY2q9b3xCGn1BPo
bv620HEtBEQ40uoTDc05omHd/aq1GrbEcxv+oWi/nYWN8oXFbIZcNBFvUCd1EDSw
yHp/Y2GNYEosmYSfstjv+/TbXiYhtMzPWBjOhlIcuyei9tx7TEWavKcI7VH6ZhYD
OLRbIioBkjkMSZLVZq87z7eRXYPRasG09vFKojyxOuafo1TYX5LHNDEu7ZVtfLYg
8lm4JBC8SGi0u/9z58tSZJkSuGPuTsrWRQ45HrIy5YPvzk2fZVumZ4Wm2x/On9yj
NxwHIEIETtPIw628bQnCj1LVOEfAiQU1yxzXu19p2aq3ksRqZpuKCfxk02YLV4G/
fB6TPr7at5t9SlnLBywyyq9guPzk4ywatu+x5/Cb8cEpDpT2SYNeI3rf5CBqr15E
VzQFiLmGe7gam9N013ldPm744HVUbbD+oYCNNkUOj5BCDWqz2m3jF8T7qKIGPZ39
kAQ3ylQBcL5U5Eur47JBr04vJnV5AKdsprlQPRBEylf7XeDK6RPio9gm9Den2dAV
yOUmRCwIy0aZkWAfocOHzf7DzmUl1bVgE+gh7DzkB877bq8wEl8wvI6NIoWPc+rf
zUpXVJx4dhyZgVMbyVbYVRO1amX5ETPBcDqvgvNYXFcmoXYxLlgUZPVb6mpwb6xR
xBjXLvsyeT/InXIteOEmoyPDLlM6V6nTnXcEsr+SCg1lGPmDEW3danxVdSJJ8Q1x
H7YzA2/WkfjRBgevmYHMJMoRrxGQtDzPQjD/WrIqQNyodZJUpefWc03yUGn75b3V
rJJOIMsgjm1PzkKqim5sR+xionTHE8zerOTdKH77SkIfvFJUx/UkqY/IVDQ23DxV
KxWbTjrIyXuf/ZoZR2J7eifOJ/KxBA/OOtv3783EyPQwlIZgkUrOd2+kjrd4Fi2E
HVhWtFJW/ggaR5KBuoSjqP8yByu32WfRhULjxHM9N/Bj8jab2bK2NuPE6tUtiBk9
1RKrrR1NuYbwGwIw6lqH1Dy3Y4nA++zDpYqBIfICG163iucJdA4oFUhkeMyvKUul
DLulUer9hJGcO60M+d9Br4oRQjSeE2v2zikdHa6fa2U+EvLLp69LrCxkylTBN88k
1haOEy7T2mjkvOSgHry9/L7V8OwJVRYjjSt/imumM+BYLnbVeRRS3nyM8GZxQNn9
fD6WweJqD6xg2CdU4u/Ov614BaD35GknTi9Zk+0cH4WTKPwVKtknNTKOJUs4F6Mv
8foHbDuZ/zZFTc6S6NAnF+NtJVwQs3Hrpq481YeYZMdj5C12VxDqg3y/8ud6y82I
ODkbS0fQuYQAsD08o955JONeJcDToN0ovq7AYYXJiuspy0cHWAGjuafebHoHGmcq
hhuVlgaUGwJI8htW8iSn31iXhcq0us/J7FtSlWf5EOqCS+h/2uWhVUIVtuCjN2t9
oZ1AB793xgncfc4u2rk+7KFxUPOEg5Y992EVpdfkob4jsFFOIJa+3rzFMxdCSPYA
p8YE+mDSQYL9lzUgF6UmpEEa/UqOWj0JCsIkvRecTKV9emCYOYhH5JFm140fH+j/
GhvcPijdfRuLIH+SY0GGItgHoc8G9NVLhvEWlFdJ7Q1qCauQoTaYzYKPS30XNeRW
GqxQTmJXtREWa90WmsyGfnPPjnvpexmIwJYOwuabq4Z5DaBd7jwSe3M+V6W3GO5r
GR1VuWFP6gnsqd2LqO+/7DBktf2Zw+KXOITYXsO8im6H2xNlmp9jgZQZwAvbr7m/
MsgL14xsAM4Z8AAY9e3y70yquymCwUF7Lsub6Ccb232mfXT4fuLdV2gYm9OWlZ81
ovXROYPisLlbKAYc/5+npvf9zFk30NyX6sVcHxxSUtC2lealKPgVJRUH7II+T3zi
5ucvv9pIiAosZizYnISgpzEEbG6Aqvu/wE2O9bosR4L+6ca/jQrkto7RZKv6BqAP
zEBB327vKk7i4dy1NC44MbTtgApcf/rNDevoIiNgWSxIgTGA7DBVt9QQ2hk74hZM
lvy82yZOPSucbDDVOVI+KwpbjTzfghHuOrODnieT+o92C6caPghES9GUxsvT9aJW
Hdzw7FVkcUK0oojTtw4czloUBqg2LrglXGW6ly/4bUyI+3sqlDT4PY5+0/30l27h
q0644pyp2qQRaDtFwtgKF5JVbBfa0Mf4c9Ex58hhcYSRymjdyy5/EhwyJbMvO5eb
duHw2qGYW3SEnuoidetyv8mAYyGo+PdPuk79K7pnIo65GRQQrJP6+CeYmMut+GOT
dVlehihefDbl/ZCVnC5NIh1AxLt44bdSSO5d/1+HGYkCxK7b4KE8D6AQ3YfYY2ll
NlGJyKUoOaPVkhyQ5zviucIk6kbEVo2Q5dN4Wh8D7nGaBkq+eUPCE2Ew0DJGO5Dc
IB1WSsoAI62mcffmCaDlnfhP0AywmMWHva2mZ40kRe1BCZ34II1Mmv0ODOdxw42A
JXnPHV9e2oAfgSq5gB9gpIW6wQJZkVihrM9KMvI3/7x04g840jQp0tInuqQj65Qw
Ch0QuGUjUVnKk1ncu1Khjkgd3n0n4D6hcE3krM2NNdF5+2zM3iyw976AEhLKs5e6
h0j/fQ5oOOIuTFJNatNUJyA7r8cqWposCKBbqZiGJWwUWExLj7jCuvJvmFHR+TmL
ABJSOL/QQulXBiD37laflzdqWxRBEOQU9lVkxaZ8dqldmunPHFeCIkpGaI2Sqpd9
w1LBrvvg+KIYy+32ZgOeVOQCQk0MlS8ldhrgZz4XN668b4Perkae2M01ZX08KWER
Nh6+OMi72jgPg/R9cSg68a2ZZAyvXQG4n1hpCofzQ5SHML59pYLWS5b+2q3WeOEO
5DfjXWk/0IorUOgwPTVBk2YQAJaQZhdTilm9OY+XJ6P0bU4wqGQaKmLqDljrrXPG
2XfR2u23apu6oeZVMZFUuNSmjtjABAETF81jmuYakX+xy5sQzrq3Bx4oOnkeUDov
A7mnHtwbWtreQlVQqE6da27BKfr47YF66xJ/ffVIMWMz9JivYieBmWzoGQ6S8SJ+
yqqPtuKuo8eJ0APJG7evj+1F3/thbFqoE7hF76idea2k4NqSmj6Pi1eSLvMD8bLo
IaCZxYDzOj1RUHnktfqBaUDj9aYpK79fRMlpmOi37bN5xskrtHB2/6p6cngk5CTD
tMyADWZQL1EteGDAKFQjQHKEqz2AdLLWB8ec6cctvc2v41nml83bLaPDlH/rDXg1
rx97cMZjIC7+N/iIlKxsycVYzPLnoXDr6890HUYQyuCoVqLsL4Xv9AXWkwFIjVdX
pJ/zpk8/9xSEStFdek2JiuIlasj/gjOVGdnLh/E4pqkYQI43Loly4CmCGE94atCr
CSG0QPznjp4/p003kQ4v203NNawMu+aSVXaiGDfBJfDW+BRgiHnsQKY96j1OW7od
PCcPFJLqUJ4fbDA+ZYv08dzpIfZ9gYEXYhncfs2nveMs2X+yiCa1UqdIHnr8zDuf
2xbYqWNzZAO/9yT8v5cerFNg7eB0/8Em4VUHxY7L0lkhb5dS0Vxn8AuFFyWzj65q
5EEtRDEAmDoKZR0n428bHtGc6ElhPa3qmNfoN4Jvsnv2wmOlKXnYT0KcmCPHtwdO
kZOVKUkwmZSQ6tljG1UI8jbc+XppvrioieW7pBw0kl61mBByiwVnEtXvRTSfAHAc
tKUVqVmEU6e/FivYeOjm4pJbCT/q+9A1Rr1RIRomKUdOR3lEG5o0YCHqXsKKJ689
+kFEqB2X4sNd6C4QHPtIz/5jfjTkYPNb0HeXDIl5JK3+sNPVWl9kXIG22Y9Tqy6t
xBOOIXWvBmb5CfuDV/J/hJvuJJdSfTHQfEwNI7xvpcgGL7nfySd9uqBKzyKZHmRD
YovWmuZ/oSa/rDxyF0RlMWoYjb8hxU6rx/E0Gt9CcPHPTu5lCBylpkDZuJNy9a90
TVviFvPRz8KaYnWjUnH5cVNj3y/xErhlKMNlh2nWHCEZWIfmoVSBGXvEjETuRmxB
F4BfGNdzoFEHxZKZrWwXdLMt2VFJuzMOwY9yYV1HudXjlwTxUUYDefvTUxfPqyqL
On1aY0SIibexrOCvv6pVQH5NbbnHncAAQpBzxFqTWVaTbpRMMzBgYD3a/qOHZVsj
8XMNZGez/c2n5CKmZDUGdHtOqIgDE8z95MqpdDiRHmQTYJxuMa7IClQemdf6Q8Nj
6RwqToT/vBvcqUNsiFk3Do2u2EKiu0wd8d0NvX78/clsV3D2Ypy8S1R8frYb2ElD
LHgeD1qdIKOoxDlVIWVALny007zXaStIZi3TPMc8u2Z18cIVdjMypBDwRVlbZ2eQ
nnk5NsXmWeKSpUv1TbDMwqVZL4A295dcNIxheWSivO3QNqMzPoG5KOcP0IhYXNwS
1Y1+phszOMX03nAGcd2ZAp97sv7HWuUHlhZMmix3MUYnUt7Nqr1LTy4bdvckk27A
HJTl59puN0tZxQz2hk57Gf79J7plwmnyQQPFnIfBr/Pz7P80OLqIogJwf+Cu7SGV
SfXj9beaxdIqtNVbIOw66vkUT6Y13eAEz74cUR1BCqrOSxFmCmn0NKjTb96wu0I3
HsjJTmlHytfhSYTlJLd3wLqfjg51pf+MP6NcxeetWheA+IA+xMNT0hEOS5rsicez
XiqKFMIcy2qOGW7NAPbvtoh4yINWJX8bvUbWtIiqBD8R8p3VymHGPgobjX6l8oQ2
5dgVFE69qNson4YwN9WawL8DdpjwaiPUySl/e0K8jJ4ytLXdTdnKD0VmObsRFRvT
AQmuMA7on+G2aDNBCuiXEt6dx+UxVgCasFcGNwpZxGLQXnciIkDik490xa7p0BDz
P4yXFuNKpeD0T1Xkt8P01PffH0bP+LS6rrIub3WZEDSOjGpRDkXb9N4/+nIGkTo5
38M3huNvSvjSGzexp/8PtLlPLzMvWg5qrxwCYg3aCXhdrSfXbizqxb3FEQcqrxZj
WJXS6zayksHwS38H8LTRSBazwjG976vFwEJ2wpk4FymyrLQmqkGXED1PD/xC5jzn
hDHpdc+2swDCm1BrKJm8AzV95rs0zlKbO4w0MKu40anaBVhqDWgmDbdbmVSfiR0l
NgLAaz0nr3mg1zBvTHCQ/ipCDE5rGH06jjtNAcpk1E8jk2UtqTOJ5EIo72niSLZ2
XzLU51Kn58EFzEffnTqPz77rpaWkade5Ky+Pg7Z3P0hLp3PkawaJ6Y/aFiiRMFYC
uFDpG3XiKajQrOfYJEscEX6bqRZ+dqe3n10COPYVY3H0mkifjhmmTW9Xdk3BSLmq
jSRImQpaWGlCBuPaGH2dqdKHzSc9EfmK8fIdgKRC1mWpWKYnsn0ChmEJ1S6+xmi6
pMBuqY7SAKEisI/Ameo2zgbpdEqXfTkwoFhasuwyx19EwCimyirNJfU8TmWSKkSb
izyDcTkZXKyz4Lyvb42tPA+icaoqMVDOKyyEzoksfPRQnd1z3NdJNLAYNAu+qmtq
tMxJoShGmH5GsBJap17KfneygETOUuD+bGGir6hH0UwqoQA4Jn6SzjnHlNveuGEG
8yzIQwqGmLaL51WIA+sesaIjvsKPgNOqSMIP4MQYEFvFoI+F1t8hU6UIUPRaxxPh
coP/VryvDjTtUF0kr/UddFZHxVCRysocil6oHJKgyvaan3kaWNp9mHVyJoOQigoV
Vz9sUaLIDZl+LqprlJen4c4IUEZlWjMqCV+pHZ7A3//CTQQptorxplxCnvT08FhR
B97Dvz3u58mnMpLBfsbSxxtqW+WRFEPInSVmDeA95EdSZWP6VhUWKLWxtJjfJme9
mbhSiCNqdjC74gKGTyZwU9uS8C6ACkINf5dhfOySyiJQZ88Sn8te7iSBcCEun6hm
4XpQOyAnbxlnNWEM6Nvky2/u0qzt4nJ3QPGr008/DGyA7fKVEPKHoFDIUnkI+KSj
yiV2IEhwBATZKR5V68ahEzBGqv+mmRwU1APFtA+SCHO4P7BLhJlhEeHnvTksL/c0
WMN2/w0nllLME/9gjH/Skun2PZMqqkfK/z05eaJDxqiW5RPbVMAOag3tTYUYDpiG
NkGpT/TO3R3hVEzINYjuBuJsESO0MGoNV43zauRBFCT0Z/SDxjWSuLPEnatHJBRV
+QlH7z7FQEa+zmL0WJ41clyw8ROk2AZxqxpDjAMk3kxtdvbEsNUfQyCUNtyo8KLe
NQALt6KnqMmiEtPrwtydB8dtw8PJAOtrbq+I0GDXQ2P8bWHVCT4gq0jYxcsJHWHb
1S3de3Gl5lWFPIzUiakVsnuHmQs5TOFAJ5yZc0VZR5hXgrh6obnDVQGp450EHcv0
0KBhdyuk5/RfNjjklcFtu8rzH5J0MOID504X6LC2OYOAuwj2kTzhzv7/VYe86nXJ
22BA6Q8NgpI4YWjgcLr98US5BjtWkVAD92C0YMfWXTVSUgfsItsPbVX+fl8j+nKS
7cKFQyNYW/DhoaY/fqjWavi//bPr6vbOt5l5J36iaj1vEdoruUwRBJzg88BxTKTC
XmoPMN1mC2EpOWfdBXAf3dewkHuU6A0MvQIlOj6s/L2hjfpRwp/grElf0tsrk8tZ
c7U9nMRGWrG9lJu29oZTn9CyE3kLHcyhaIIWMN0clN53ywf3ATwcusk1froT8Weg
3+Lr2Ge7KM1LsdjisosOIz1kl3avUg/4ksYWarwfYIysiH0XDxxSiOa0ASE1BzAG
K7psD0citjaWjevCbnYfZEbSAP553PUO4SKqkPtL1nNyrVIoqklRdckAeVHuev1O
WWZdXtrdO3sgRdyIDjre6E0q2r1H/9p/0RX+P5KnRt7X8Knh1w8cQFhdD12ItiB9
oztHTPYAMRBgHMC3bDPEhkO71CUT8XryWGluARBGwdMQqmiPfeWGFIbY/ufqGA2H
r+uMS9kkq8OFHl8Y0w0isMMFFkAd4vbeJtP7n2EwlzJjZo3Erp0qHnjStEjY1rWD
QByJ/3YEki43O+GyIj/MTc8MaeSAkLN2By5VmZe/6TnE8IVGqBaNdsLt/gD/Oqvf
DNOu0RKfJDsY5YAxxEMrlrEmrdM1w+69OUIB3DYGhLX4FpLQFOmg8NLzXfBOhrNM
Fj12Fvo5WfEyp+DN7UHjZzEmcpKjmrsun0tT+UK94ZbwHO12BXOovZ5QxENJ+VEa
5mFCj3OlRAaAgboURRdEmcJTREUbxT/Tza+P1A0ayDJaoUfL69mAvInk0xy/6yku
DJNjKbF6HLUbvAyV1+FWUwryq0WW1Zrp1XjnRmP7KPtKNsoCAGBTO1Dp/zPGoOqo
uGRzxeEOczKWo2pQvvgSHtiwUupZha2Fv+GOI68vKFUFI8lFGFz4ervDOx9Gwbm4
AZwFzfM6W23M2v6qbmm85xHcnCjKAlC18j7xD/43X82ItmPRuKcYbh1x5uIC4qvA
Zh+BAnDBQimMqbgPM9OLiE+iogek3VjwTzWy6QkcyAC3sIBM0Zn4wBa5M5AqvBFM
S72jWSWePwX9EB8f3nc/JR7i3rJrESqGTAKuHvHusNxZXmpZkBscKfWPjNwMJ7KT
lG6R1DeCrYMzkQKHojdFfBG40pp11vtaHf8TT9v1MNxrwIwhl4dvtpftjn7s2sfy
wGMFXvlpG9d9xkbtB4hcWYmHnXMsCrRZfHJ5+VEwjfbcmKRk5e0KtXh1rVsbpj+7
ENQOhXyoyzUkwgmPMUjS3A7W63TJm/ImVTUIt0dMJf4lxwmLYC6D4G9YR8tk99/z
ygauYLckSq9C/fEGH+S1grvNL4GFbn11vFahIFsOGdAJSS+Wit5jGeAaU4tSfjBQ
0+3CCMqMTZQzJTQHwNNO4YYmlaL2AvxKHo2bfVwjdntcGQFupTqdGAz54KhfE0My
8m+Lq2X4wZGwwpP7R29VzkJKbFl8YKtFmFHI2uz4xKZDDfpAmyJLpAZDE0zPR6o1
/pP5e4F6vgOHNik28niEmDaczHdEsDcsdEAtrqZb9eT526LeFjIfi0EVGCdl37m4
rNwRBiUmGAmj9AVIpCb97ilrnxhJpBl6onjwbPeu4F7C+pSDejRVzUeR7DTRLncz
eFE0JCNp16+UmSkASjE1fMc94dc7n+HEw+uvrolWSzAIYkDFFBL9KwvnmRhg8Rtw
YYcmqaJ/cP1/PzV93C3rQ8+zwOmmUYut8QtITAUqb+cyYHKqe4dnZmo10IdtW9ed
vU56wPRq2fsFx6yMVVKCH3keTU/LcjU8FBHXO/hTRsSJW7F9XOwdFh5o1ZMC2Gn8
6aCfpRj8ZO49TNNrV5qi8FpPjBak+orvVRNC6/Rl3Z9dc2aBFEcHimld6nmDicE4
BUDznvvdK/XkMOfEekPmYdsBdcdS6uJvmGZqyN4+jqDKqEuasHy8tK8sogvWXSu2
DEl3tAzXsrOYgzcVJjCbJC+s68P8oEUI4vwa9o5tDKUDGdiAnUESZE2o+akj4yV3
8lkG6G2H5Q4QRC6lIX9OlWfhcZpwn1ZSFolwfWjxtztE9+NgzHkMa6wuNMIBIUj6
QwlQPJmwvbXIa7dZ12KqhT/62oDx70JY53/cjSd4qd4NZJjZHPryv7Q+xJk5coH3
f23/br8mImMgNjfR60+fv48I1FGTTeI4U10M/B7vsFGG7Skfk33vM+/m5Jv9NCnG
mB+sOUnJ4sKrWOZSODtmyAJsHBtCkMeRV1s12TZ5c6IH1TjL1ulfi02lNxR9Fu2d
y49D+8dfOJKbHcbuFpSl97wQ3m8G1fsrph6dyrwFeX7UQYCvNv9GdrreekSZ27al
uxl7tvHbFI24159izz8oPAyLyS0FDIxUf8Ob3SX7MEsr0kSTQxSo6hKUlHFXsuo8
JSHCWyDb7TegmZkaXNMJbdWwYYrgbtuy/EZ3uMdDnzkZ1xq49Mb0oALXtrUHRDcL
irFdcKb+t8y6Ef2rXe6QqVE1Er/+KPls4kUG/nlAiyL6xoP9xziKECU1HUzqpTYG
UsL344nO/ZlBQdNnpYxr+A/5i3Uldabk0jXtKJtx+T4/hB8UOjl8/Mp1K98Poizb
4Imss930f17da/4pYR4PGgUHbrY4/y0DU6UJFPsNIayZGU5n+3d8RxpG3K0kSf9x
PafuEZuBj8gZd0t+ZFJrzPnHDhPszN9WgLP8ofYFPJMRim+7+AM5l8w0sTS6+cMo
97kD0TJFA2hhfevVNu7cOIHEueTjiAJR1VgVTa6Jm6+CHtxVCtfNGJ5HTIqQsCMV
TgQivRGPz6HpnZ4QzLQH380znA2gaKp96i5LhAyO6ZrWaDO8ER7Q8oCxgkM/3qtF
H1tkTlYZf3G5OO7lI92aXp3YPEHntQEpHpU4ef+kc2brKQ2Cps7qXQhT8CHzhMT8
Oz3AyNJaiOQ1kYEZYtEoeFP4VEbyz7jn3e9j7TizBKJI24AwbmYk0qaKYggS3Ydy
d0m55eqCPqbAqObKp17KMza6oHXyjLfo4BxuSDQk9TOkfiVtc4vS3bea5ZorXHe1
/umrVe27oggKIdS4yIa7kHk/OhP2lW+KPz/ercDQGIaSh1yOXsxlu5McDLbjdM5n
ebJ2KOhe+dvi78T6baFrPeOhA/IVH98faAsuHLY5CFvoSIRFFvD17K/AsYm/DLfB
ZBPFzuQOKe7DOen1YwdutphhOT1C2oe7nHpJjx+gl2CF93TAa+nM3JELyJQwy9Tt
wAnZ+74MOi7Uiwd/njU7PjyLTIiiSv6dLJVCMi/Wb8YPizfbII+W65OtTx4X/2BB
fJnkMyLcctiTJEteSc5PSHSDedBzkL0+tdYufOc5KkE5fLWh9zaQ0fWcVihAJljp
cpilPeBNtb5sgrshk9Orb1ZyUn3RGAE5MTQ9hZAb9cSZL4yI/TTXo0Wv+SHGhNiD
76RyIgyL2WcnkR2I1hCCw2zhKlJU5S4BKOy6ShAI6D/6XfPpDs5smN5kP+1pQCsn
+VKFkQMU1AM3qAs4jT6in3xuwotxh9clIANCLISYt16doVZ3VTfGuoJYL6fKEtuA
iOar6RptjthKB3UeDbCuwU8yEaDuPYBPJfnszx7lXNAa0bUobdw/QSwcziWuMSLt
6aMTFx5OTbt/4o1CryS51OxCvyRDeNv3P168s8ccoPmtDtwwQ8R9yUGkX7PwSho9
ZXyqVPzKQKba3aI5LnQkjkb5tbeBLikFSbYCpuBCWZ3wKuGWR/pk+r2mk+Wob/g8
Rfho6SZNCd43ND714d545FzbWFYE/u7AkoRvtIsU8SgjEGYbgr5Pqo1x24yR9lzt
mZXDwMpnCq/qfK9q1SgEEdfuBvklin5XaonvYZARWnZiOBKipEoxyLAuRWFnp932
9311Pzyjp+FpZElxrIqpWavaHJinxWQwv5YDZgIeEP5rk+vGcM2mdx4oT/0FvyTf
Ri84lr8P4GXMq6TY0VTszbkym5r085mkoSIzAkk7q67doVnIc1UqJTcG2RixyiPd
AzdHS6LBdwCPp8+zQw6LeY6a7qIO7brMEpDrrVCaTpyh81MC01gTEDg1GS15PeoQ
OcwAW5zdaNU+y4sRLjPuQCk6GxRAl/ulx7l95bJnoYnGfU/Zaui8xj4Hw5B92E/y
KzAMaTj4voXZPcNMRdp/oyo4Efhxtotz4QsafZH5nC4pWNupoZHs1mWkJo10/IPX
mBuEVIL7WQM92Q0MrFYgYDnSZz3nia5vJLA7T0UWvXU4//z3Bs3UTikTgOwf3XuJ
r6yR1uFMPrRatkBVA44lML8Lza/ZiYQ59hd1HLjQGQpgmsO4fDRRMbOL/Xa/XvXr
k+PiUIrbRcmmPl3HySEp6IrwVHXrJvfa5pWqdq6brpg1AvndO46WAU+fclrCOI+B
fJkyiEB/293gb29JYat4p1f0lmuedC9ooWWJHqvYUnNubT8G/HQnKOjrFUspQMjy
0WDQ/oexbNfEEPxZ6fQZTSvpSHNBKLtgTIS3yrTAU168ndy2Z2qqJEujAv8lfUWx
HlixMTbkiEOsMm8vPlPSFItUViDnqYyokuXecPgDNiHxjIdNo7pAC/uz7nNdNj3r
K65PTGRcA8TEwaoZqTk517KNfAjgeleVu4QGGoYtpcC398I3AQ4Q1pt30hCFqY59
ChhEiT6bHURC/Wqbux9vcC+QtMk/3IGBen4OQHYNInkY+9HtNfmgPUMEZREMbSvF
bqeqXAywnKbxXSpwKcbwZVpKtVA2PpvcuhtuMrdfI6AgUtpqM5mtD/IF88FfTKN8
WiZJYCsUzQ/WequTWZZaBraPH9YMvRaSrJU4W6cPJcjZsHzMG/u6wnaiH+q9lVA+
aS4ioG4L5AcOaashXBH9AsgAoUtBCFq5AVLqyBZ3EsEbnI4vNipkrE8RSJLiELq3
k5zkRwuhFXNwUyEI525WXYOA6WsucdcLBD9wgvo2YZA8FkRGzmdvRxKdI37NksTe
Q7cxkAuHjnXfqWgM/OPPfHOJgefigtk+4G2jYCGE18EK70L0kaED/mgj+6q8lHzs
lRjgvgrsv2vDHeZlxwBDQr8WHoAX+sOnOum8npA7Ies0sps6bHseIWGBPqmIw3OU
05eSye35m6BDaS8cualnaclJvhOdH+t7+XkTF6qmv53YGWIxs7PTF1M+7XNaQzHz
WQ/6aEhtzn1L67LmD8x0c/kFjww1fr+lCimveDDEZTfkOvYNFQadqoWAHvbbosuT
Skg4fH6MR4WB/fMZb7dksU8zS2GzlUHn0OQ4j09PhbSQQnPPzMBrT6b/qjsXmBNl
bnOcqq7+jJMPBFJRsDUArgy8St8/c8f10mtOk2jiR2372AiTk3XzTbBcpKIkGULW
3vEojlhIOqx3vxhgqoK+wApR9EimEAO0/7K3kydCupMlsgJkJJbRXEB70BhOnfjO
LYexGQCw/TSPEfEoeHhnfWoBj8BcRWX80O/NuhFcGfXn7fbbod4ywyj+5rGl7tCA
XotiiQq8DL1eJd2XYZZVBoTXVVfkblneAIJQDJQuEbKMmBoW4BgHs4wbHqJ2mM8p
HkaOb2+VmyiBsjSYTcdEx16Z3kxYVpatUBCsV3mmXbQdaNgMtr0Pd4weNZInT3XJ
gKYZSDkWNmksDyvfuFcyVd0GkxmBrHkTIM3J8CoW47QWa1sSE1VIxPEqS4yRemlm
UrVAK0EZLcV99iJ28XDVWufGwVnmwQ7eyYi3ACiSscCR+pQTio8LiVv3yV/ly34y
fKsLlvBsBYG0uPOUARrrPzuzmb351lWBN8DCtJuQkcDYPnjSGBfrqsZrVHmrj7Nu
R/PZ/pbHeNcv14K3ImSfP0JNYOI8Ez+Fy7pcVUxXgDCqS08JDr/JCwYTyrTpxprZ
/Cp2uvuJZDQi4SnoFn0+R5Gw0ADSHZHjDlk+1r8ifrDHiiQreuMw7DMPjbPYnIpc
p5QPGGfqkYfhAjQbn8mKOSpT67JJwNLxEKVbERoCwJ/BOs1JP1UXK3IyP8vzWA6j
M1b9ZrTRGBITwBMlHWhZnKIP1Ys7RjatMNeyubL7I1ZNXv7CyVA2L62+BAVZUTli
2HKwJw3O++HzW9csVAqWy2xnKlxsiwmOCfkRlkObq/aGkPVyhu1E5/wGc4uno1jg
M7RKtqXJKYZUkpyuBzFxVLl0rDBaG+jlJNaEfw5/R3ZEtmlW0oZHJQDkBCKmMFXr
NCD+1cOEPyT1btKpJ2e4b1fuUgE135lJMnxYhNGvTshMi1/SroL89+moQHGbsKbZ
Ml8e7q63QtWPOslQlKQR+VLZDaSCZDluNPIV2R7u0iu5yIcl6WAgIPszMFsSL54W
mqpD6Yb0LZHWy8LerOtt0UfbqxDG36hEsV8K7JVQ9w00FyDFeINzvlshiheNb/Qe
7sqk/x4ltrA49VLHHENxKunR8+kyVcjiyBw/bYtBilxT9KZ7FgqeTcCI3tLfaLEq
BqWifv/bapSZVI4V3Fyc2Wd5818ArIZ5VFrJWQAOYqKpiLxSz85hoOnakZQJhv1q
IDsbC1QJAmWGMXOQAtS0GNW4WbpibsSWWYQ3P1Y+7kIr4x9Ck7ROOm/myNFmUNWE
n4JSZgxfamQ7LkfkpWJ4j8ESpburkdT/SNNCFjienHux3vQ9olOAHesQByzfBYN8
llsUIYy4NGcA8m9LU9xDcGeQrgWQSmIsPqYJh3bguAl67cBKqPUoTCmYPuECjL67
ik/aKKUMWXvOrvCPeIGbEQXzhS/IgofeAdE92JEkBn2jY5q64lYJMXgqwPBALopT
35proA5hRFNRkOUCI9KjUhvLiUSTINBlK1AxnUJ0VXTArxLrdZ0ui8H8ScLWEwvw
X5JZgAskZAyxD9JOckQNXJVTUS+BhLzM0qJNLi9pokJIiABPBbZe7r0FsNPParFp
bKXIJ8O8dtv52P2CaCg0NpfEliQGmdFvihHYmNja15y/8tRPEz5hNpjAgJKwckOk
r7wy697fwvQFJ8RbPGvjhXOuurT4kke+3EAtRFOxNKmS8yOg0KBJ6tNl96RPL7Yj
NT0gTuBdTi+g8xucEEDEUYtExkJ6Ymamp5N/wMmomPQyXtljxrZq9mNqDEdRY128
Lrq7wP8GKBvYW7ajAlfLBvTc/JjEDlV42nV4XbzVM1EF7RaLVh5UTkCVjp5Ye1Ra
2ExQiUHRxJE0BjQnYSDr0g4zHUaJ/RWHtli/GyhuX4PUZsHM3xfOqzYbgs8kJiIc
qE+eQLfgtiud/8L8rCgraP7ma2htDQmZOXSOFv8OAfU36uYf/73oKx4U1kJiIbF6
wE2Pvf8tRYxhDZFvyhwoZEZDOvojJ9LPGERtctYrzLG5+oEILeQ9GTwNnGzobo2T
P75WbBGHZbmUrvoWBdYQ8SYPsudYlNYDcQA17H7DQ/TQ3OD05JCVWqyfDtONrywi
wAxYAUC8t5QAA17ItbE2oDFC31SK7of7XXp9uuFqV5+VOfNxadei+aZAXMzcfQ0c
XwDqbBNo17kUMRsFEbx0nS2jf0LUsHZBG43bpfbDQoEIhgnTplEbyNyIjLepVtQh
hpDDa3K7Y5CNuik01ulCAxflz8OH9HtHe0pWsDA3RYqz+DuWdLZ00C9NtWGun12q
VmgC4swuSDDTVbK6gWZ1gnngu+psfRWUqvuEpqvzceT+Me6wSrdgmfDP27lewf83
PGmDv2OPdk6exl9wIpHFsFGArzerCt3uVhkc/ij+nTP5nBUUPErmKxigEbE8XUUt
koYlpf9HPndz3QscOglyZj4jzluB2vkh1C948oMMOdXK0u2/EvQ7ab0H3gGUl8Yo
oKdqaGHaDbbd3347bXKWNZtyBYdZQV3XhXErmtFBHcdhPiPjUsGApQmFDlJNwRvU
Z6HXr/0OK6W9d+VCB8rUAAN2xBpG4GpbS08w6dMksLmX+R/YwdfwBJoiOBjRMoT1
NWrvYKQnefk9mAH+1g6dk5qsXDr4xhNzE3rhWEIex3tTUWt7GEmuN9VF/BFIpxsq
rCw52iedd9amMgyqk9utVpZwimxQ0WDCAPgkKLNfyrUMtXux0kaeUnCuK9IQlpbD
3yXzle87etTGrAOuVqYuBleOP4zbVlKG6o0jsu5lD7LCoUKCiJkgKeS+cCpA7vio
U4Q3NsJ3IFr5DPNzkZeUy+e+7DRBgxo4TiRs0WxKFU/xQS/23YVEnJ5+VZdj6/71
5qz5mtEBjlNeb8ZENefQO3RQ+26VjMb8zyOXEBp/nUPPqJexUYzBf3ktvjDI/AoY
v6ICMoaFP01h2gJc0YUaX8ArCOn4PZd+8rFnO6tbHKaFFid8IQ0WioL+2Q2FSrfH
8bVMC2PwllLwqaJxHR2QD/FUWWKS9e1s/Tz7v9Uk1+BvjMOgL8jKGmRxU4KqqGMH
oZYFycHWPPrExe3MBe9UvCBvd00OQb8Q2OOx4lygQD7687bWrUgxuQ7bNT4j4Tlf
RkqvtKdtjdox7ReF9PEYDkRyJIGEwqAuq3f3yCdM8uLRkLGxLQh6uxfbBxiTBOtO
UiRv7rGhXS3sgj/fNpW3zvBGLrvZKpGmAFirdpfbF6/Yxn9n0kips5Cvw/2Utb6P
8RDtkhKAHfNGmCGRQ60yP12xjXvgGsS7hkifrH+eDitbx/6JZg6NoiLyGiscLIsc
IaSJZPJUqGHSL0lUNqxxwz3yR+Y+/LeJVAKbsAPSsjsP7s2gexKR0Ea5HZ1HzzKY
zbBsRKHUHx5BsJzL9BCC7ktHcy62w7yQM2ZyuTQZKYL4UGcUiPi8kvrQV9hU00yF
kZ3mHHz2YWxmZaElcB6OR1uNsuTRENvUE3NzJzCyRG5XNLzYQ8953+Pu8pSdiQgV
sarwOekrkHxvt0CSHwiLevR4NWsdj7wUTEA6H66mOGY9cpV3yV1bmtQjMdq4ExtC
xjU3qx4CYPCAdtpMpvbIMsS6hcPtoYnbt9mlD4qtiAEsKPrkjyUyTGXsbqjI49O4
o1uv7VL5S1GPXPvPA1GygW5hkrhe0BSYXpjlrsqRAjSaKnyNRLRgveC0Izc8E59Y
qwiXewV1YhGZIt/CRfFz4MUF55YNwI35FAu0L6Bk5u378pP+NIVNNSOjLnvduFlo
cRCQCONowxdRGDsHHCzhol6wEkJDowoB6mC2X4z/ci0+oGZ1j3k4zzoz6D+SRcQ0
4bMVu9ioyQQBGcrnY6VXoOC/8lo2b2r9DxlGDbcXYCByPVgFVmrffgoOGsKpsskh
q6/6nZbQgTf84rKclAF8/euit+e2SrRYW7anRbBRWsrMrNrnv+Eky0ACABnRQNd/
I/KyyBLG2GCOZ1NHf0MGGpekOp5ZyaDvkgs45GDlEH2Dz5mKUpL8sUjqqPmzEA6B
ZEM479kxlQteEOrfc49+Rnzmo2w1fIY/1L8v7FCZ1uSdfGkp4Taf8z3RzHB6qlpm
lY705TgiX74Ouzdel/BcHVtPmM7fIC1MnMJuYkkOaZA3po0EGg4zAiniibgYSrJh
Gsk9MWy9XuU0g4LDunPlHG5rCRJoCTG7ohdijUCjZzRf9lmta6RKxCiA2shkfgAg
byMf+wS0HhVbpWMx/COd5sDhcEAnLcVsW2t6uLY4+J82/NIkEGGE8K6qcETvFI1U
WjbWDvO3A0lsmcwVtCY8yZORiFDouP6VUXaJ9smiwN4x+2+OJ4cJe825SWw2LYQB
Mr15CQkKrCAaz5JyH6mYR/LdyHur7tNuMOc7geVRWuVhqNjhUru5+FqrSxHO1TMr
v8WHrRNjpL9y9N+0fp0bAut9yqHeF2diftvof/aVU5wZ2demShggFqxeNAJSqg98
kVqDwcaWogprYuHL78kJWuqBzZy/ETvKqfgLTc1QpH0mFLHK2HtEBkYBRHLnPhOP
2zanZcGJsIbpIAcfcqduI/AB85uvysqyp5gjeA9Bf4Kjs1TbZ/4ZwFpcNrEWe1h8
TU5EVX2GnunksSwKyB6hJ1lkp5zEAvkUW3MViJePokKhZfpz3RhbV3yyt6/wqrTi
WKTdTqyTbkrVq9BJcAk73iP8AViJ0lgotdNuRsvA/bxofa4JQZIPrqKHL1C6YmmE
fShG9e75cZZJ/5/2wL/MTXe7DF+6aYJA4QTCS0fJmOGPEYQNiBuLITlPH7OEIDRa
1FS5kJ+tHvdOr5+d/l23ie7luovgCVzgVJ5PSst47eLfj1R4k6gE47g2uV26E+yq
ClNjNCaYE1C11up6l0xbYsJylp9BExHqm0keK8yxcc7Tu9Erm352R8Q9DZudt7U1
Tqvq4pwWsbJWID1wAbn3JIpgon+w1Y3Siu1bIOq2LTeVQuO6ogzVuJ96j9DvvQuw
eRxcbZZck8562bKmgXI8rN6C3KCWVUfpyauFMJygxBCjcH3OPGZU0hh4kxNOShV/
J5oXeQhivoKy69izsXf9wITORnZMugKDnEFPWX6AmrNXc+08BLMNYx4fnKkPFTEj
dJB2mTS3pIHgSFLrOEhv5a6pkVjvhBQGI4KypD0FgeVlBIRYMcuhy3YEHyTBNdQC
kx6tk3M92WpRfLSSO2Ir8MG52e7RvfkzTCAiQo7V97AnPCi/8usNhC9jAz3d+3p6
+W0sRga7B9arcwL4zp9Js5lMJ26pyvO1l7aflPBGWpW18btRn8nlgj7tZFPwNSb+
2X8pYrKeeHZ4TRXlvPaDZsEXzOQrdq/YyxgLOfrDUYXlku8+uNj8BHbKkatNaueh
waQ+qkzQ/dq2BZTJaoGKTMT2Z5fT5Vd0NYIpee4CjVWcRTty+Tqjnj3qkbY+kVix
IZWhtoTBKkF0ez3cSfzJDl99NiOTN2JGIlKuVsc3NMhXZjqKrlZCCX/LMIZ7fEcA
X/ExCkBI3uq/3xBMd5hB0Lj75kypNsr3vs144MBOqlanIJ6vkH90WVRyw1eU0Rpq
tNKt8sSlE5g0jzVoufb0cEoZw/AJ1w2QGhasoVMhr1WpP4GHclJklma9mecM2tOo
CddyBZZfYY5313O+gNfqAmfJaBc9N00v7QREzy546mO3EqtC+FugqW9FwwCGIxcW
oSbk3uZPWizXqydrbBjID1OxElJMBl3+YSGxyhjxNljSCK33BPfU2H7XP7jwjTzx
p7pPFwMghnZchL+ZM0z5fXxRxbQGlF+LIscCJaUi5jcuoBmqeGANyoeijG0QrH4C
z7h8ol4U7mRHewLC7p3SrsAh7j/eghson8mpPrFBZfddSvpD78+lrgArDTEDaGA0
E94PSDyJsiy3lnj3hECT5ieeRnBC1cCACI/d5wR8H+mOI/A9kWhXNeE5zdEm/gQZ
KFqZEIqdbA3wD4STw2igsZ4gFHX2miaqoAiXXStUjaaNv7bsIQRAn3BQd5HHnrrZ
QCxU5nSImiiqGlBZm+pvE4v0iDUY6+q53NIWXIMxI8jf7MyGwGRzqr1roPQBBciI
C+UBDZcGJPNpT0AXur3z0lBLg8sMdnX5d0IISZo/n9ilPaCzbQZe7tNGbI9WpKgy
27/MyWY0JlsoqtwTnKblosfY5HDhfz531c4xePkifa5KdJKpjU6hFJDBF4fqRUD2
fBSB6WxoVoAee6clpGG7EB8ricp0KRLL6NaG6rzIdrmSYUu8QLGlotI05lIFc3h8
mHhJ22w2zso4Matnv0qbzgG2mf6bsnP6C356cPV8BZrMZ4l4fd0YKyX0pin0Kh0y
i7OhNMflx0tryNmOCSWcvrz0sNyc9yaVoYywI2XlOtjfW72AC4dxJf97iSiSELxB
RlQ/C2aPDx2Mgh1nr1BSGPz8DB6drqK8f1wTRCGQE1heW45EUiRWIoagP393eSNT
tHVaFMT9RLBRaFqYOVUV/rY76IwLoUxAd6HHDtwJNWIR1FflypV7WwtOHfU0RZSV
qKk7/Plqu/JCPFIWgsV654+y3A2QlKYyvMdt2LLAI0S1IwB9VEO7aBUAF0tkURBO
p4CHTus59QhAHqjnp/yAVI9KtLNGC8R5xmCzuUFCqB4HyvkJvdwUvM9OiflqMTaq
K2pcMZwIQjs+Xs8On8A7Y2MiM212drbHLzXvacfmDejd3p6Y7oSlN5Qak5jAx6L2
aMRH4U1O46EpqedX/yDgVK3XhxbODtbo3dFcS9Te9ynCRP61H1kVglACRA/5KtJ2
7JjZTH53LZ95frGKU4amp0hgcu/SCCQ8b5DUqK2StmR8KcCGGzo+Cd95q5FX1wTL
6uEQsZHaZBimn7VF9RxlzuaSCiZ5NY5ZGxLzdsG9S59FU1KN7gB3a2goHkvgllIi
P/F3yJjdZbaQ03mbDwn7CtnfaBTM32PiIfjyTv+fVnH5Ob8hafZxwJW9BWkVL3J/
ZuEh6BZ72s/lgrXNC4OoRMGR4/UpxBFmfsoh//ETI6kuwije5xDn2p5iqCZA+LuF
QA+vYXZF6AdNM9ClTjWrvuqUYjgEVJAe7as0Zj43i8EjB8AYEJnps1t7sw35pZci
Vmv8Sy/T981h91maPhCaupMsV/3XPYcJmyLNtg98zzhkO0DzDnHD/LgBw7IvhXzL
5/leSbCZw+Bb4PR1Y9Zg0sp/yri39zo/L/F/9MQtke7rE1ytzdqHT795YnbyiSP0
4bNhj+oKFv2Nu8w+eYVlZnxvq9Vx5D17xqS62DlFgagBoDSGOQ49iAiCPBoQ5Zjy
REGf9RipGa0fykktHkYS+zFEl51SuIP8nQ9L/ZeZhpiwp4TcLokSld6e25l3bpWf
NEZewiN2GhurwRHQT3QQ/x1D/5fu7lAey5Gh3dNT+kZn3pB6mxV9m3rUd8zUzWU8
WZTA1LfPZUSCnchzoVCkd4IqN41Gw+f7e8fshOgaVogghyx8elx+9xsvCfQgJt5c
3yhkzUhNeBzTwgHM9TQfpUkfxZePx0Kx1DEpXeR9CZ7PudTAZyTTZ60Naor4ZTC3
zsP7Wg9B/WUISV0ruJyEo2WjDlWNPfk1BdVuzAhpzbB7MSmS3hsVjIN4fZQFrGR8
EJmIX0gltqCourx3jB8ocUjX0xYfT5dPkdm9MSki8wF+BlBs8UqYB/46vwwuIfCL
CprI+HBvAL8X5PN7BYak1BlAI5IUmWsTLgNEQJoT/hsiwO0WEa5XEuIoS2ytCiD5
xzZo9PNaMvAnJPoito3ANIQAQhJjSzbnpqA/7g5mqUV0shcYXjWwk0ZUvLjUAR14
sRVQ7TWe2VMp6851jNCyXa2kMhUqWXRYczXBue/OYIgSh4h+EzhQrQeYTjbhLJlH
Kx6RcNWKy4gW+nTUGA4mmS647G8DoVxZ1rvTl7NVtoJnLE56/eOc8mcEIlvzuVbM
c5qrbd8/bTSkVZhgcC5BxZJofJlbBMAp/VXhDmLmB0oedBBJb34XRlQWziTino3X
I9W3KyHkzk4/mT2paXfkcTO1AhPWTomwi4VVDd09e1zzWlFUFXoyyursNcxXnovj
0oCIZL1xZSf9OFFCV/6hntcO1u08LoPoroOcqTmoL+oXZDqWiNkFwIXI8F0YQGN7
c8g8HeOdQDB1fD0U7loEq+zBkdVCJU5U6VvsVaj5cupIF1qBaMPXi+8XD6xjdD01
43ta1sXG7hM6I8MRbljIVlsAAQ9xZ9XV+3M6x3UKxLWgKwxMVYlIf4wT6FvEwScC
uW3+ViQZAW3ndela8h0xmMwAKtSM/i172dhLpLKK2fcGwTok7nM97RERVEtuPN3E
eGymEXVzVTk0DUe/7HN1pEfHF/S2k5VgfIta27dafOXRgn1rx6LF5nH9TBMWiVS+
UO/WKK7PWjOXXp9QMOGHxyiJGOCiCP/qyiPHvgd1Qg6YVnmN40ix+oppp6iYc1Yb
Q8r3XDma5m8q06gw6M0Jy3d4wZQvBuJwBw8+RqoM6KEvOKb/dQ/sQoWJyMFPswhu
pR3BRXuN188A/OFhhjgopbbxxGXOIE30VlSVpq+83I+V8wxQ/MGgVkoPlZpdutU5
CL0QvNnkmOMTWjS06VAyWTCOw2s2/GA8XopweOv1lZCHEa06U1CnknGG9gpjgKYd
JO22ZATxuS8A6YSr0/xGeMOl+Pt0LzK+DmDvi/xG9DhixYDvacPgXI2JCe+iQaaf
BC0mVyXVDoGwTbVOzOD8AsluBZo1+QFfswUHacsvXleLA70qCXp4WmZJ4hrX8fix
d+r3gLzRr3gLqv83bCAxn5DV3zBFNHYoBXPyaLND1sshU6teY/oBYEJ0e2rC50Jv
Ugitzuqa+/s2DBL26N9nqIbDjomFqE3yOzSL9KC8LlTMCqhy2N7PTwmiaKri7i50
F8p6j8evAPieezWxDs5LG+annWXCKWv98CCUz2CLCoI0wklkvWX+ijEgmespsz8V
A4SZCpBgah65SFmVNn6hO5pH4AXfZJPYmCK0e3fFv0sZGXDXjjV33CFfdxND4BuV
KPXFOe2QAc7VqiKAxN6XAqSfH/IqtrcwN7cArw2Oy+66EyKzdDK7+SZPDsg1W4J7
Z38XCVfjazOoOG6Bx+tTAqM1YLP33rJ7zhTMxCQ992YSsIICWLbHcVEIoqop1NNV
U/NC471jKSfi0pe98GBBEZY+iRP/Ejwr6RBS19aSgDR7OVZN0BbvHSbT9wYu7ajj
SbdfassADfH4xS8t43yH7XnRpalV4sqqQmIosm7jEOTaSmEmhSpKc3EwD+9SmSeF
0HsX80kUCbYMUprR440m2heOxTHquuFDbRUjFbtT1h8paCnpN58GF/FEd1tY0vEd
/GlQT9AoCcZz0EN/AQpLrWvBY2nyQGqKKwyPh6FQwStjMierEUa14pkU+bdsb0rJ
GisVExyNUkj2oxuAfuEAcXrpdeCFWJWtbpIfbhhvHRtW2CRUIvkf1W6edPKPESVh
F3XPCm/YJ5ZzXlUqHh4AdM2XYKx7cgv5uevti6ZIH3+ElDOtT3Revlvs5wREgE6p
yC2eTfqcz85XfuMLFhyrijXV/kMDGgj5R80LgJOI6AZcvJP+CbdQkoTiz57TrolM
nSqn46q091iFrV/4nMHsCxI5vSfbFLbc8ZlFxAyTAqWd4ECf8fgyYgaiUx6bQX1B
3DLuB7zUPk0dO1CI/+rG3nl1gG8hvrO8hjA7pkqmDwka0ON0NZEMdASPjoDy1xQz
sz5Mvlh4p+TD/ta1deLHe1/MfoLznb3d+zKkNsmq+l22JeJFN70Q/0QbjuTooC6C
m1V9YZBtnuT20hQDkRBm9VGm5PLf/pYqdZNN7Sc+fRbeiZLq82E+DOa192Xhv5an
0abPypuUjb8OnF8FI+uNhUMHaDUXovy08fKD8GlnAmvN73dNnCJhLv9PGwyer3XY
QanEBC5WEjAyjipn7HSPIRRmuYN3arlOMvxrmPK4Gh2EU0X3TzKs+eFC9zhfbfF9
cM07RlyTtKCBcGayzZ98yisbRJx9eCgDkmm7BT61IpfZPgL8zhi49mKHZ8SiSYov
oUdw9ntP1fG8RzMX5LAvbnMzVweWSeHpVI2hlMv25gU4qjjy2IOSkmSKvt0kjDaK
1QE3rN//WLP3pyJYGBT9IqOPF2K3wTGViPtZ3uodKYK0A3OyiC69pCZM3939oaAU
4tHoUGRsgQPoxuBaAh/+Ugu6UaTTyX4nmVGrvVCGLj8RW3CfXH+sGRisgCm1EPXJ
Jvv0QzgCnRcNyMKW942chbHHYm2nmj8cVzRBTFvIqp6azta1nblWZnhJyg62llWA
qW+yQQSlD3GNnJ8MQA1Tl6uzCXshBXi6/kmNAoTlYev7umyNFdObnyf4XmmXHdSl
qPoINJ6lFO/BL8pRCv/6bhnCieNKaxr2auoYS6AQkMNbMMnIP6jR+oyYMfuHVL7J
qq535xWokrjG/oQZrb1YeCMx3HC1/FjgSqky+XI5a3LshZecwqs+RgaJ78rQSuFh
ddwWZP3o4YExLAMJZLT+umG1v97KlKXKiwST/12DkhHrf9/fPvLjNBGMuPX3e3En
9dWv5/MksbeiRL31DpC41w+AHkws4WCuR+K60Xp2Ed+eDYCnnTyM5ToU+LbskBdK
fNufEQimILCIXTxu+St5jTtJJYpCkVCBJW0DchFo8AOf4NTb3WUbJA5rP2Pznd/o
jW/0KTV2L4eApqa2xyyfD8vW8RxA69UdFBt40oNb7Xak4Oo+b4RIACMV3jelwuqH
mZ9dpNKlTSKs4kdZcmjm2g86MrU9mHxN1QhavcrS3x/WDlB3/qKvCJd2fJ2osRI6
/apK39JiwLugmdtpcYQTMwzyH9HQdIItIvAop+Y0ySP/QNYydWjha41fKVkIrPfH
jHT18z8WyqGdorpMfraoI+DmoP0G6RaxYu7jyvMgG0tU5f3H9Cn5uynY88ECiRzs
bd2gv6GDV+KbjZMNtjhAavNDfW2Z2orcADejSdJXDehDGlwY0EoSiD633NoZ4TPD
ewAZdBmCPVtH/EW+Iboz7RQo1Cf04xU2ZKA+XdQNZeGNrzLhs8bLDRKDC9/NgtOA
w7gasa1jlTZbqYsDUNnw9VvnVbJdhmakQtZLd8hFNrGYqTyT1hkgSsQWgLm5/oET
vjLasIIGW8AXWbQT0so1R+U8yQA5Ft/75Z0LEOAk6w86MsAmoI/LIOIylvXrIKkb
1eBBrE2BXL8pRzoTKyG43i8AgvLycLYjKvtxkt9M0E9FDWvR/S8cYissOra4hg0z
6uG4u6qhJQ/NTjz7Nd1UwLaZb27BkBB8rayfAK70TaTCw4NJ110AkvXYbw1Ae75S
masR+5OmSzFo690Qnm8NGJFjIxP9vP2ZU4uiAh7OOpGJv7JLq8vTDuUbNXYUzPIn
AyR0qdNBSw1yfbP9fo8itc0pZnpqh8Efbf39wQagDsuWFuWMzIHeqJ/NKB6a2BT3
0GJG4LjqOxD9QKxBaDRK00KVo7Kjaegvjz4yjGLCyXB/+q13p/Aao8Xoq/iDUJFW
07PYgYDdclr6XHVnUWGjlqauZ4ri5jEGA+sW42gH0X440SMvTo5XSEiRvjJQMfa6
KAlXEHoM5BE5Duxq9c0nxhBdvbfsXd1DqSnuEtOkDjrzdWS10OHA6k8WsS8X/qQy
b4s046XwJICZbRCekt6CzY0T5bvGfCFAS/BDTfsDoDpPmxzH3vawFQC+olxIwfRz
qUfwOYxY1tGt6JDuR+PVTMoHddMgC9Vvfr8oDW9ao7q1HvqCeqROqM3a45NNjpkJ
znCjkMC0WPUlkzJ+WVm60eKWPHj+WkGTb9mNWFFRJkcdLDUEUFa0AYWf/S4ATO9T
qw8cTpO+giNX3wSMKN6EUqKh/LPv9jI5asY3SfTfT7FT3rifSTc42Xt8HNh7XaZo
oie/vz2+i9A9G1ABVU/ZYBsHOG62D/t1v/OJV9K5Ff0sOCa3eZXbh24AeOtqxUXz
i6Pg+CLCe8WfgLrTJ7dO5k/FGUrU7fnEgIrUu/LhTHiVvLhZ4LIOkZVgIkcf0zrn
dy/OKP/uq7K0wIoQZty8pBbqiy5xTb9kDC6nwQBosCxLQq8hnbmiMcvVTz31hXqR
LRYL5ZwGRzSa9hthrS+4LMkVYD456zdEHo1VpoNh3z50cj/S14H0NKDwWC7NbzaY
BmFCwpbXM+crZSu1pYXwNAPgWy62xwbcNLgZ5bVTFA7D+UUIjFvBuAqsOMMAkQN3
oVXMBAOhxVN8/jthfJgMqCqqf4qmYVtB7GClW6pO6pHd1wdeWjOsalRQW1qtt6gn
KX+DQnYLFty5QweNoRhMFuH+4xS7W7qZwW3y9/8RKyDx9+ZkS+KktyuItc9PbcxE
i+ZbUzy19qsRTUNBYrV+pQkAc5I+utHTW3HTQH2N/OUdN3U7F9NyyUotkt1+OzsK
z6FSTsMDvRYrd9rMQQEQFEVcRc4lHTv+VFhH5pF896MuU/wA9Xdb0XpwQdFjIUK0
FlvFqNHWadAOI+7K50wNIUNjfTrTZDBWY2aHPMMfmtz8BE3LCrxrzVjAULfQXdfa
OT1FtmhesMSH+dwZoyXkSARW0cRMdX22cruvktz5eEnwySzjj0xFqMpx5C3F1PFu
/iNYskvw29pkI+JnCFcXr5jetPaJJEtj47pN/MFwHQlunpLjENRfh4Q/jSkEc1zj
BnjBGxWaOZknsxxRvWge6FJEoR2Y1xjkSv6nz3biWZlgIWuYLwOeca4dOkDSrGbK
0A1JCfytyMNEjKsKYr/RnD2L/aGsxMl3nBudFC5+5hXQ0MYLhOBJGSGEZO0k/nID
Hs/DB+sKFeF1+QuTNmgnoKBQkolqaQZGvBcVadIpsYnTBJcWkmTMLwfk4Tdlzng9
2DEb7tFfwBWd4uYwugfJne5Tfi2/cRiwNJavgbaHsNDt1iVHGC6CbCYRk29VhUSX
OkUWB6nFXoUKkPNZnZvyF5tYRexH0vgfX6JU1gCl+QLXdqUo3aaGZqAYFAovzBOU
KSg+i0LaA7SO7mKMkDSYeXOIZ3b6pghZ8uPse/MSvBYl2EpwXZehOUXunwTdBaiW
XWNdI17gXhE8JYbn0XUZtkpuJ+9uHKnr98GjWYMM3/Xgvq+dPGVSFw4nU5qYd6Fp
9fAv3Y3S/0NrW6givRaYg/o2ZTjwcVJRzkOImYxMRh3odHkPPwcv2rwXPNOwn6+e
foqgJXH2/PPcDVj/rndd9Sp5GwJAhxOXITr/30iKj1FYLh5ZZ9BqmPFPrAe+QAx+
z3ZP+2JlAHJ/9B9YY4GCY8D5fMH1TCe73Vu0GVt9qEyPV0SqOtn2EQRPNqP67+XV
0JoM9VYUx15a4TUgLpUzr0EqnhjjeVaJa8+CNoSA/kPA/TmFsbdUG5Lx5M0wqLXa
RJaKDMdeogpFzqkr34c0NjSTd6pLox86lhGCsLUOqerofWk6trkiAkx69tnl/8mg
CwJ2up1mPjFDjtdKnZvo8bhKcu5/BYOlLyTJVOks9E4P0alNOrvyoQyHHvFjlKe+
vk631R5K00yomgoboKGYidyRKMVvuZQ/lzMSScWW4pNfLG9u1PdCQ6K8zG4hvKia
WT3Qz0FjXar3ZGXaD4qE3H5eLkpVbZvbYgjk8utzoBme7s+hdYFpUnLtbww5z69L
Z1agSUXPoEBpy0g4k7FuDEz0xzcMGYZia4unZ1JBQdSPHP+tZqiCRByyHFPNXB6Y
KmIlNq+ZMwHqXDlz8gINAfwrcl8QSR++A1VtXdK62wmP+6vc2FY1epfcuJlS/pNh
XDMH0l+nN/Os60xrlxHQ5rtIMC2HZaBvBtCZob6OkGuGX5N1e7ThpmejWz/mG9jn
V474wNa3VsVe4+EcapLmOZ6Iapx8MUzzyuv5Ft/iebQ/EFsP1LNxQ6RME7e4y8Qy
/m3gQK5/VGrTZRzskrVeHI8P3oogXsoDJs3G+ShcuWgOxKVrcIB21o8jzk72VirC
jwwWi4FbFXA7yH0HW9TANsy6VGkBA0XIFHsBUtw3+JbAy+JPkNOOuozTgBZZ2tsm
xRYBTHwq6oQ5Fi3tF83V51uW3h2OvQ9fkTnIW+ycx8l6COz0CmJjQHCJNf0N5qcA
ZsZD9rHZIyVnndnZ23OwTorOsLUxVOw7gk79EkVFyUGrSVvu49pnx/BcYMGIc+N6
Id1fMvN5UYhn4tDh0oDnTvYSzj5r2bKxYKSzhE8KlquA/WfxgZAwaUcbI6Ukd6Iz
AjMUffH4l5bE0Ma5pTuDbLAv+NyPXsHatKIF6I+Gk+PcPcHKwMvxn0fmVvahYvxB
UkxuwcPJlAWRWM8kbH44uC3KIEfulT/xk/MAwiNq9HkTpfFLSUJ2ZSZyRpHvD2VJ
nC8cKzovdVmHMuHzzykb3z7XgFe5kQLc3mMLezAJlwa7DGQc+wQwkggUdyDS4Y7K
xPkYK3L7TpHp1YWrUL+jkZjo53wiT/pB/ZXnNxBXmHmkO70T4cCVKCGqyU7DZPOR
2KY15ll2ZO0+Q0DB6XXUZ+M+dhXdjM56UzmNxekZ1IhZfILzvXpV1nQGMx5ues49
+Gc/HrP2C2ynmZ8HU6mPB5jsdEN49dNrP6OOqxiEaDxH1womP1xEEBEOyiB3Ectq
XeFYGgQTAgAGgGUXwp6AP5EkxNquV4Jii0cRKXDZEicVmtysqgFmqRPICoT5IP8h
40k7yzComsZaq7QSeLff5qL1AajyPvP5e30EBcfQ+6g2DlmqVzmxtr8CNOPcusck
MqWkQzmkB8Hz9Dz0v1YRV/yYR581QqCamV4QMem+9bgqV5xRP8zG/1UaBxYo/t7R
0jN9GMgR6JXjMhxCitJus6hLKRqA460Y0uj9DUdtRg2MKXItBwZ96AAz27u0WjZg
BlN7EmxxsZ/vDkeoPiltmDNDAPWFKdJyJjWlGDf7yZ//UgOdVWKWeYiFIEpm4Dq4
JA/MDawzWyBoVCvT2PDgiQSV8k48iSoC/JnyfKRF9Ks994883MTDX4CHWT+bTU5l
HnQk5AvheIWiRZfJ0kJSFcZezTK4dRrZI81t90cdKWJnTlJp9Icd6pzU7HT0tq5Q
92Bur2JwX8P6S/6cOH8ycCkF86/B/L9150uZCcPPW9iOi/Yq8oE6nUdxdZuAccbw
JhmxcbrTRyYYQZ3OH624r3SGu3qpFWUwvU8U8+OTsC2w1IznIMkPO7rlWRmw1Nou
DFVU504LbbcYqW3FERHuIyRB6PNKNhaDDttxffMmBobVBCepj1JPgiJp2RuZdi3V
j17mMpROjd+CbVpuphFUuHqrFvIIU6f++ctvFA2LFfkC/KLKU/JdhiB4TNuhYkvW
4tsN6feeCJr4NFyZaKVj6Xy5wBBda/1oxUHbhwlv8AmVmhWmKqIE1LD03KKBpP6x
8FjSerO1Y3mi+ljc3KsdTUa7UMPAoGXMb32XweR5/dr7fYVRyILbnFAJN7yj0lql
3Z/CHiD4bko+2gwCxEZEo5s5k2bnnxMlBVFMmA4sXEtMkyCHSj33CIhi5Kgpzm66
P107rbIrN3/1wWzLsxq7jH5xydTuSmBoHEO46H/ej88EAIZJaHKZz28ESAxm2U5G
XH8LgFhVeAUQvVwy4pjQphia2dUOE3RLe04L/bpnoMt3xqPqlDRi+n3NoIvr5Ppn
k6iYSBGE7mkl62YtdFwh/a3gQLCGfnyGVdwt8xwS5VbZgedg2EVak4jEr9hPx/eW
VFLXNO0LMi9F1yZQ1jG2zw7dJX95fzeMm8VZomZgLkg+IaXJYvAYPQDhB1zZhkDP
bI0UUgHslDVv3uF6qSiJVxdR3u+GvLAKdesRLoYPKmVytWBUYgQTukkjwSkJSRrU
0DvRG21W5UOb+KXDuv1nREmqgy+mgiCui74F81LSHM0iV54ft5Wq9h9PpE0qS0pY
HYiipibnRn6cDy14ybw+nbsI/0L6uTxA6PK0MXDNSYaZOjThAtKV3dSwsnTIxBtF
ZjTq52592GameF4sYqQzhgfsL080VyQt+OBtjfBt5w1gd67ROhnUfrbwPKFcxqj3
hu+bZMRDQIiW/q6jO3m0JSyUjUEt3UsL6JD19CwI/cTa07NTQh/UkTgGn3VgGU8d
XDTPXmMH1UGzjEg3Rx0hq1307qv8y7npOZKhkSodeOC5fHctiQOl1YCtxcPoTJnC
cgPEFEcwgaS1y0Yflxv8tsahI4Lc+hPx/9yfsgSPkjjzl3tHFOsjWYrZAi2Jpaup
jxnjlAxcsLMwuCMVDgcbMHqEJy2aZVZiE3X3uVog39TtfRjJH3NnUYjbg92c5wuB
8d0zyZTNU87HOAZV8ndnK56tVedxpozwGKTGNpFlV1KtetgW2VbkvQzZmek/ndP1
JKxEkh259PGf3CBu9HP26Bk1tNDyzdvZko0cR+UfhUaci0Bq9R9mFzVMYJUwVZem
hEJP0RDei7mtzQeK37rvfMxaR3Ubs9dD/BEcUwK5ribSLpJzaLO4UP2Duh5PsJ7H
bc6OfWl6GcwTILL6mTob3PMi9c6giDvJGPs/yS/MlkfMhwFW+bf/YCD5vBanp9wa
DyOsq1CThDsWLF/hYKOLV+c8qxjl5bxtSZyzC/OHvLgx8jqZMAem2H6OfAi155Al
z3ModjOivtWdvrsF8tVHge8OXehNpM6AlpI/9YYhtyUYhajuNuHtbXE9yICzb7Ym
8HMaFi9xMNZexWTjzFhgrJDZ0TIXK+/6OVyEshbAq6LWYgXfmxF5OFAN8n/8R6UA
Wv+KAO6/eHEiMx9T0shjcV6AeD+06VjsbQR3lVuQRANofBQYM4sFc82xFc6eZBvi
hGVo2VjXsako6RUecl69pKmFZAushYQN4KGpx/B3J8g2938tULsyRQSbphtb8Vqv
yAiyGNsB+qMjkS+x4WxQ+lyyiPvliP0Tgl94ddrQ/6PovAPWyzvTgzrxZzSN+9Tp
Cb6FMaDVQcWkwTAJZOp0rYxCdjsxWVedrtFXsQkDTb7OWMNBMlC8JVxpi1ByUaNo
6KTYerStRzR59K1jm/ZEF4vxNcumDvyrD5oiM4eHUzXq4tGyYwOqzkwMDDpUrmwP
yMQ8UrNIYYTssSFg/OorVJllWv2aerIiU+/qQQ87XuAVAhUIJ8tfnNDEpA//aQxp
BKRg10rWbtvcBZfQc/NEVYinHsFWdoGErzF68dqBRJ+m0rls5CAaZD25U+BOj6dm
G2XxyfAH6371IPkgrE2vcl/teK5TuMp9qD2EtG8FlvEF/gONZyS+Fkl5SAT4+mvj
DhBSU6dAn0sCDjanw1dWMiUR7jkYWHjpk1O/EnOYYuFlSjktbRkjJsnqqFhvaY6d
b+/2hOzAMyv0TgGZ2PzX1O4HVYGB9/qL++kuV9JQe4rNRJJL6OgcTFS8/exsvrkN
MNxewh7ix4s84i9PPtu7E2pnyL9tRUjHi41x5xwuVReSmnkp1O+ILZTmNs0/9DQq
xVM/53Q50zjjg3hrrUC2V2WFYfQSW2BIoOsl9Ku6VfBbBke64HFDU6d6wR1tDftq
JIF6uC2vEL7XZC4R9iihD7g9+r8sn4q1ouEeA34UvV/lFO5IAi3SzJQeLOWlStIj
VwuOxjewCCWcx5n5P6SSfNv/3i/GGQ7XJYb92weUXkPBGsyMA+tSyuTTrqdsQ8Hu
BoLbLUmsqgyTy8+GhL9JOTel7kNIUpKY1cOo6c0MBQqmEaYy5PKY4mrgnZ7yhnwc
I95tDXkDSBQJBjVSrTq0QBI/jcXsmFgOJlbc5/q0+2xWE9u5cjZA3GsarPpH3ltM
iB1tyXBIow48XIo+o4zENLINr9p3XtDpk+0iP72yQ6aFn+NGiSmyb8uJl4qoWL3g
pjHRKDHg+aRS54CjxJdNWaq/TVcOZdQlE70Fk0PqhP+8uKfTMz6STmJxZNPFJZUB
wCpwruuu1orssRjjNFPFkIyYD+hQZ/dAVwhaAHtGb0XK33M3keZmNZE81dFzJv9k
Z04COMeW6Mntjb7Y7/wGv4sN+2EbLplpIcq00MjNcujAe2Dzkv1ffhFEixgdbsd9
mAFQD8E2Q1+DI5xGnbfu7TO9P5k1PB5xYSqRpSD5k9/iltZPxqI3LnMAjD7gjtYK
1u0DkGoJmTmPLGh4O3Ok+CTdDYi1YL+f/RDsD61gQzX8RFGbbPKe9s4yclPTkaHk
JMxHzti8kKBwSFwdWPmDCNmhc4iLhNR5a1qJhWRT6UBGjV1Doq0XMWcwmZWOTmJc
EMBh07JxhtceJjrdqekl6yGu6OW86yhd4Q9RufF/Ew4Cf81+ztNWpOs+5246AZt0
+Vx5uH2MCamtLlbKYko1npwA0pQWCUYHvk0W0pKGnxtTtmODBSLH3h91T2U0rp71
lXHEp7ZlpRYgwYysRopX5lLl0agl+WNj3iv78+VScHWqOl6wM39DVxAMVwl4TFZ/
kpf8ikJhZzTxs8YPEgwL/oadEg45zUxWSPYTc3c1yYfe5QFCaW70J87BePopXvWw
PRVCJ7DiDnTMNxXBJv8SbSLuAKzvea3gwXOW9uxoo/l1rqKlf9HLN+DSx6i26g/U
5AANmOBzQC2ou7mF+SM+LO1UNt5OZW1XuxLnCG8SjcAPG2tQUKc4Ov6mQsW/EHse
gSDHX7Y+rUR0dRAs3aV5BBa/ilr2pEFZTNmjUbRFN5u/jP+GPXKwqkDgymsa0vQh
UANyqcuSvphNFZY91FAoIATOzBv9ve6P4pM+f/7sIRvPgeQ3q3pMfkcBYnjdLPxK
1R06Ee9cFLMqTA5xVZmqOYwyuOleE7Z80Up61UqjCAQ3WAtK46VE1ICHR58BPrtD
jXM/chgv1RB1hxTM7zcz/aqY4StE2P/+ulaIab/eGqRn8tcna9GCDaEr8hbRuCzV
S3+TBczFNcQ7UaJx7tflj1lbWq5Um5gQc3n+ATQCsJne3YJj62aNKM4yaorqI4OX
6mzhZRVVKAGeMoAnxSTMgiBPIs+GI7Mc1HjXVjSpaVQpvQC4/yLweF86gti6zum7
7GmYexFvI1Vs7M3LQUF9ecHLvGTmUzzI9vUxCgZD+1jxfk1rCbibMVnqfgz+VQXu
z1nMVC00Dp6TSxcVadS2gbIvZohmznnznsjXu9aIRb1El6mQP/+xhaBgJfZc828o
QebzQY1sGShCkm2bc0UD0CiW1vR+4XnowaFrOE1nwtqQ4nqQkycpOu6eUPdvNAky
r3ZZ/Ym6iLk4YlKSQ2t+UX4loyj267VHtiTUBvNrrHurVskb7P7Hfa6vyO8saDOK
w4sIbKHyG5q6w41JUqWv+gJtw0sWx4HVbT0EmOwDdus6YyLBIHgbT3a4p59KjYbL
iaQGx79IqnHFu2c278q+wacuXagJXGUhoJLh0gtDT7qkmbFvbgBcJU1uK7JIQvDD
/G+RMfrUwiY3rbH1VtHxMIsYNopDyjtyRa3f8ZHFOfjwnpAYN07V9r3CQehiWQeF
nuvPMpLgZTpgjrseEbUUl1iAppz9B5H2e/oQk0+p063GqvRMuPKYAHyZ4jpjxz9j
Wxw8G2enIqhwYuvhpgVkz6mCrfocjStaw7mslSCOqbpySciMHOX9KOnq15dvPkna
SlSZFHZjTT7JNhT/1EG1Z9+S0Zj4ZncOwHhC7P1biPoyNCBtQpXa3ZAmzupqbVl+
71MMDPLADXkpVkS9cgDSV+F/ULjGdx1yqhC9NMjdhgBEdH/BebzujzJuYJLwbxqs
KfE9MnAMTqFZFLZYvN7/QRQEftFsIvT1+8raxVexDs9UaApCeRfdbtyZnTgzEsqu
z/7itw02w7P3BQdwQxy4tOfRuWOqxml8BEbzMtHrRPud6AcGOPzBZhB61tNF0HfM
2ydFbX81Velv91jfKCU4nNXvuqfdqvuCbhOR5BmfJMsg2J47ADR1+OgDbRSpipIO
1MOosrEUyTWPi90xviHm5xray6mTRNStooDshi+gdA6/jkTZNH7oPmiJue4pljBh
j1rF+NLAoy+VFe/SHOwaRTFS02OodkaQQbvYBENUTI2oFZdPJijQ2jjDqpzSFo3W
2QWDXm3hWmxza5lJiqWzby1fHsZYYaSnlQ6FJ6KL4s4ffcsD5hyouC7MANJEENFm
mIL0Jy421WrJVH71Z5ssP4gXHSCtxBm39OMnlLg11wPdpG/ISCVp69e3N8C4kB8L
6bp4eguS54l4xW0aNbhJeGvSkMCrZkHX650yk4woXxAUzq0t+k7SYBa9et6bDXgD
gBcVKUj0C31c6OZr271umDD0NO4kCMov0znai/r0A5nKEAaFKpymRzqwC8RQW58H
7bhdVTf1plQBlMKnp6+4UTZoz3AJKCowkd4WF2mhm8KBrSc7fGogq1skyleOw/la
hX/WYZi963Pmtd/iepCq0rWLtB1KIP5GxEMih5SCDxXcf3HOACRt7C8Qx9jusnbZ
wG0kDiPBPeYYFkjHkvmF+wm9u7h7W9R1VAY5LzsZexhh8mhnHl4KU/3PUPwxou1x
zHrx3WB82LYDQ95E8uDO3nxtAdgPb7yhizSazk0/WjZ+8GR4F7kE1BXkhlHcE2r3
3s066UAD5rxro9XO7jgVqX1IMUXWm6dIHrVpUAswlym6P6opuaKXiohQ2HHMv/WH
kX9aEDYh5EI2wC0ysn+Q1+7JUTqmz5ril0Nn1K+05aFlOPoeFLODxIt8/L5GqKEf
rKCkyBtWy074OoVOLHiPkTU1TQWovwQX+zgLrdiYn223vHyk8pP5uYLGECjgtRMf
ReECOK2Ap69iM8Kz/vbA8iuOQ5tpYNjXK6amS8Eosu8gECvy+dJcfcD0coZRitpY
W2p8+d+VIPy8ggSNtndhojV9eMQ4efOTRBVGkkJ5XVeezIyossgRnsq8pQvxMFU2
whVbcqpsjN1J1u6+TouMMVb3PU15q41gcOcUrYsQ4cBduiPoKsXy/U0QybuRhs1V
z/Sr6liXtTwmiToYFPRXQLqqolEy0+Z74d1KRgivEQHu3/P/GBl8KYucp4+wT9av
S31JH/smcw9INCZkSo4/7T32OapZBpFLxg1Gu/hpWjwirubwu9uSBg6Az8Pkb6bd
cLH7+6BI0yULnt1dQqaMpDSTgu+kdG1O42+7VdEktR3HIhdRrbRKoBFmwnpFg1dk
OTORPYzCGaO3271ASMSbkQ4NBiOaEK8ry/Tj0qasvMxcVYQArNEaalywXjnS3A0H
HYXFGOKg7V/nxfjZKWbaWJBIKoYMclJ0O60DBX1KRmLs4/irTPfxwyHr09AZJSUR
25Z+huFWIHfnLz3beQSaN2iU6SPTsRCR+qGrWjfLX8FBOCcuO2/DO8edP3mIlVQK
b4ajJV5t1Q0LMaA2C6NhzcDcW6Zou3jPHmZA4gbSQvbrgyD8wl3Irghrwzb2KbEx
r3zQNDAJEyjqFtL0WssLsb4eK2MIob7SJUy21lauGxzNOP3tM7Dhn8YGPGYfVVjw
9J1TJ3urlK+aIF3/PYOhDZVc365B4cWv8K4kGYu/WiUjzozniHPMTv+9C80MKaeQ
b0xhs0ujOycw+HruachzFFk2ks1QuxgUjFP7Fz/UHnDTqywt15u384bFa//fN0WO
sfDsFXDO2g1cDpT++8SKNFYfBcg0SBYng5nEGr5japKeHNKoyzjHNZT/29ZuE1E8
/dY/LQORZYr63ZXlbSEB8J9xvp6N3yaFXzahg4+uJvWL82otZFK6OjhJTBoqmKak
ykeupwo6K4pNobMMLggCVGksobuMY7XuPk4ZwBBCxi+sRbKNMk1NU9VeS693LgUH
c3Wtwku3s23J3lKy+Qd0xYoivd10CnGI20mrNvYPNYuoE9RcP/6G5+z1qh6Ivjc8
yPuruOqTcPDFxrP7OV+8dIMnJCidvCgysZEWO95X3L2WkG0sfitZS/PV9TKwf8ZN
0WXSt5YQnz/fZALbEF+VkaGiWWohrDrmHeRHYGjLuxLg/G2MPAX2MoarEG1AtKEr
GfDCxY5LeBkOZgTyr6BFXSQ0cOgjAuOb3KV29y+FFSw/7Wv1a7l6tJBxf19G+KII
ZXpP/51UHTX8fa0WnkSNSrhG0BYzd1FAENGZn1dprsytcoUJ1xztxPWcge7A3O+I
K/cPW03d6KAyld1uKTO+fVbzAHjWEK0C7c3ZaJ9hNitHJfYexA3ZrynLc1K2O5Vc
o2lXd1+yKB3hVZ7aCyrFzcXlhg3kmwzaTYExn3/vT3kKGDhQ7AT2LkgxcLKNz22V
yr+pCt5WfBcchFkN4HfCND6m7kWN3a+QDpH/Je60a5ByYprI22Z2x2bhvyJ1c94S
6hZ7L+eUuvKAbqvprwkXna9sLJwqPWy3Ze+fisvkkSKe/UKhHwExMWszZIlcWWQf
VFPrxWMzJ0N+k3OT/bF22/OatPTnrDGBHbzhK7l1U2KZDXkcZkDmMybQ/IbAA7gm
XwaAgy7qLH1WI/7ou5FXhuIxADD2oQ/+hEh93rwVTpLeB+n5vzT3wKu74rt6/OvG
1X5fxu63OktmEn3BRYznLATgW3q8NhUpn7swOc0wA0Ei1ZMKflMr3NvJOSKBwhZ2
MEH3RfGPHP52UJvvBs12KVjEsB3Orto2GtyULekXwoTTKhZ1P+Ea9Zzl8slypQND
49gyMn/Yg9VPSnv0XjwMWNJzdx6XGioPhhEcozPkhjJWPLrCZWwEnz3+MFKLowQd
Usm38VnUbA07n65N3Y0+uDbSiBD6jq5L7X6gl3kSn6LrnkCFKkmOEu0sHmpF0HgG
ZtRIhZHPskJbYEaNS7A+dqZmAVo9tv7T/qU2oDGnxzZVHBbNiZy8bcC8rW676emC
OCvLatxRbef3+Vz8LGmijgp4CA7eQykSqobZ67z452dOtCq/gLn8v78cy8Y7GXE4
BPzks7pOYhUeSbt8NkhKAt+LBtFQ+jczX5GxwD4KbU7uJAHhiJmjBkRwFi5bAvY3
0Xe/a7K//YhFYG/8gh+9B9VKU2wjelFATtSnm5NHEyplVUM0U5APpuz0f7P92Zs9
ee2zv3TqZKHbCqrAZrV/AeoNAzzzYTu1GjBdu8aYHYRVETcFC6toEQYatqwIvVGf
GaSiuNBhtDj7YckxKvDJrK9hU7mbIZ081WTW/TjAIULIrsPcvBVycWhOXMRGhNqP
whMA9e7HX0wAmbJObjybixVLOH6VXxiW4+3fjqNuXzkbcoPeZSN0GCrZFTUbk5Ys
hfVkyxPQQN7+Atj3DmVXl98m0t78uXki2IUDdz/I/tfaTn/LpZzGT5Yd6ff03fGx
EiJpBj0PR5lCOp2tWwkO3ExDSPHxvidUh6Sae8ujH4WP9WeV47rkZe+MW+nTY2iJ
Gp56p16R2ljibERwP1UU0ZTqKf9Y68IGdFARe/Yh5Rz6FbUDYuL9A8a84Vsp3rPh
VjNWXPvLWeto/ANC89SFf2ZWXt0A2fEqWkdk3ut4VmBFbKu6TMx48ottGkIoLAMZ
5PXjJJSLuRCewo52PXtLjr2gna14Ti7QH34D6EFHoTAzONQff3QSxLFYz6X8DT2X
IVd5AXEdSYu+7MZXQjerXcND4Rlw55bZm3umbwd8sCq/6Hn3V6zGOIPnS2KG+5wH
6p5yAGuJiFLsaVws7laMNgSN+XHCE6UBefknqmegP5ugydH1pelBkGPridsF0HAS
UsINxOjTdEzj1sCU+ZE68UdSqxEFtmr1zro4+r1mxiNOsVlm0mjOLg3lgjpIrvvy
Uck5GSVCQ2cY45CMm3JPCZmtJiXPFvbcvdAcWnr5ij8V07GEtakRrh0F5nD6MiUi
QbDeOJFKsC04L1cb752bL6kFFXIIzL3CFmDDP+RUHzwP6n9E5j9p0m7thtHwXQH5
/tHHpcC7q10lhqSoYGjPysrkQN5KiRq5ulVYDS2VP0O/BdSTWDFwwikEnIp8h/6w
0p9V/YfCkPreB0AO9Qt+vzKjj0TSIinY0rizJKREjeov6mGnbnpRL+39rXhE5UyZ
3sQ+UHM967vJnRYm6Nok0TEVLS1xTr3ikLjDCdcEosUBzTGl+Hr6mMBOjvliQk6c
mTQ5VTDsgXUwXzPj8Bga1YTQ5+IqFSMlRPTwo9eXqlrJ5XuI2lpjnfTwtyMKR3qA
0+K1ng0MXSy+1458+Xa8Tsic0w+G0GEhCjwkiM+bwy5pHhETO6xTVjtKJFsojh1E
LqxLpoKfZMNtbxi9rQHr0dBV7A+lEWWd7VMsx4jRgp9MZVELl0o6NwSav5le+4QE
PV586vwNkpbyDXmwTdl1eZylYhZCxQi0/BMcLNVTNUPiQLcX/r5pq7c5vI4ZvhJr
85LeYxGzDcnH0E06pVDjhSvZHcn+10UOAKSjdIaeauwNUrhw5lx9A4dYT8JWMdcm
MTfkf2HfU89MaEzTEO0jpmeiTgE93Sq4BRd/7gkNwh3L+0og/kzpvKJzGkpWDOnL
erR8ff4KrsMscfKSo/GiWmYFKTLFsTrFdTooN5Lg47NP5NA6UVBldgkqt+TvoQ8k
SsfeZjBaQoUWZ7SZTMcvZoEu/bOkkH01ewfvi6hFnyk7BUGLZszTm7TbRLXBz/fN
xwfXb0cQUcU3dU+bEnWYksUsjptjj3lF/yftrXWdisEUjXoZXSe3QaAgRA6oCns/
53Q7DZ+uygnFk6OJVFI7evXehW8TLUxMaMmqYG+dIwyG2qdnUGUrZzGBxMr+lkfP
u33v9WhYvrwWSymAzFtz2iEdVMjSu9CtwkBAYEsxRZ/Y5HpJ5w1UWhWPQLLbXQTj
v2O3J7A+KjRPv571w5njYSBeH6mb0k7gS7K5A2c/BQAwt+ZAsM74InulYhlo6N6U
nOKerzwVPhN6Zu7Ijb2fW+2a125I2PuCqyvVAmqqhHH8K92olMeSdfLdkyg3+fa1
1Zz4NBqc5rkVavoZu7qZd+WU1CGKwwJ1E4ucEEGX2qx6AONqcMkUHjCix6JHBdwe
9MxvilhMCzBBrNQECFNroAHpojxVBPR5YEJE9tQ+yTWjuTXGSb45zygySoQ7KB4r
gw9RniLM8fBh8gn9hyuErQC4jjI1Wf1GGu2zcak6cO04QpYP5sOuctVqdIr88qc+
w+aI4/RXqCurt4zw7wkFF5peGGL9pcnML9TzUwc2KZMbEeIMKd3zt10AJEzha+8W
EnYCORBanPK9vdz83xwRh2bOGQuFPV/+i/AFbabqNrg03wFbjCDFFWJvqipBgPAu
OC8GWXY+X3KpofeCxfu+XdPj3jGi9yr4qGSzxfGbMWmaszVvUO8GbfDMPxoizQMW
yVugBcl3lGU29U3Ka50Gj+58opT6sgmBWD/hXzFt96iS4tH3bSSvYfubEZBiaBYB
lQrUpaEmffKuc9bZkwjJRXYdsYCFJCegcBZWoVe+WKUkl4Vco+rnGm73sCmLsgrk
nXBMWFp8zR/T8olN8HOxLiN28VHFI2KBA5a3CCERzg3PVo1jcTqAJHd4CVzk0REq
b4wMsMdjAKuY5eXrAG7Be6wKG5RflS2FlcPF+3EkRyXXZyfgUJg+OQMU9f/vqUw0
WxmDJ/1RwMbL2yNJBBbZVv6al2vvD5U12++p8bjQDPlA+4DRp2/1G2d+oOattMQ3
6Es3+2Ho2fzf2U3wSWzbj3rrca2FOQg/Tv5j4I6AhVcRI5hSKyNx2PRkrlQEZoJi
9UkU7vOmQnMgoryn4/eKCVhhBTkJl3/TeoI0DrhAwAS6D8fIKRm0dzUvDcqpArTV
QcqHn42MXKxRND9z2rjp7V+6j1j1wbfOJSqK0HEkdlv44Bsh4PHGhav8XHzP0aAH
j8gp+GPJOok0533j73wl6L4Uva158pTSCUgiixi3zk9yUNSSFwZ9cS7XiB7vACIR
y2UlbroqKTl2Zs/c/ImbhI5NvVl4hZy2jqTPceOEQcLvu2zDuwdCQYd6qjlfDkeX
E1RfQfYhy/KfHi/rsmW037wZuoEdsA8ixd4ieaS1R7GXOuOOBfF9hmaLs65mWVCg
moIoCXwHjC2sS1WAtY+DQtrKa/2+JQl6SG+f3s1VloSNHT4h4FYQEq3UV3zVw49Z
cUSp7H0oXxPhcI+BajlbtwLq9/JTVTTWlriJGh2zXz2IK7bgEuiQg2bPbZtf87gp
4Iolp8qmsIeqe28sfvqWsqHxjfWJPU7xQYvOOdnf3yFyVIdzH1Sob+1pyTFZKCAE
3Egm3OPTct8xerwd4sgafkq9pHbzFsvdTk1z60byPJsJ/pF/YDdAauB8meGEUWxy
lAlA4bZhITilIqECC1l8M3k10U0YXvwzw05rdKhogsx9dHC+oRsR5nkv1EOBoGME
AIyvOvwFVwMCdFjQ4Ik8cW1uZthPnDmULu+Z5rc/10yNRjQuPyKPIAZ4N+evusWF
lhC5NV1k37PPTjkR8CnIbIBKxr/AWfnsFik3QaWFoYBuMyUwveUP+OBteXUQsNdX
4E8I8Z906cm3NZfqTIgfT6x03FNBzM38AhbWGnOX3FyrOJnY+NpMLKQrksuFiaGz
dcX1SdqB51WpfakNJvd2vL9fNg+z/lWtcHyX3MhaHbU3Sir5Qt5ItpH57osZzfco
3wEXXCNuHS6ejhrgaPTukcwvIHdIzTHbHAhx8Q1YD7Y2EjRc4frvRP7Cv3Zt837S
JZ6cRaXqT4wFeuZGF8yV6S8szy5WYOXPL7uQmjlTG9tCRKUEG4Gg5XF3wl0BXHkV
TDwxB0mFYgjRfYd3IBnZP8PZJaVBY28AhDp+hxPVl8jdmRupoURLckV+GfH/dG74
0SF4jBm2AhyFp+VLasl6tOo4q3ILZc7EinWtNOtZFBThOhqFv+jH9zgXXwvDIg06
KV3x0yoVSJfjQIsT3zyfVh6/Ksk6B2jKAPDkj+tgFDPYYs7H5wl+/AR3fdKoIdo2
phJldfTKr68o91NVObk0vbzGaW9vwZufkdcSRhYT0gsKeO147zEsD2bdw3fB9YgH
Q9GNZTGLRzkBumYQ8oZtwXbvcS6VOBrfUYkobKngmOCrhqA2bmeLatLzzrVx05x/
AlPJfTy15fHmvMy5lprrGkciC7/781VBcXS9YOmEr7bFUSLiS72MuXKAwI0OyHde
Pj+tZ6FBUp3qZJoDGz0BCP7l/OSNcYs3u6B95i3YVuD40VPbquCfhdbaRthY74cS
sifTdh/rGrBRB7xG14sYFP5FG0lfz3X05PaL33JsBDbV8v57yqNiunZQLoe2Ib3m
VHoGqjME4FBDZNSgaEGGIGB3f7AO0ezvgm+lDH/MsT8uvzfqy/d4R7VT51hAkIZH
bppUabbXEcwSDSQryE6ndPAur/UPUFeCALydo5pGFyjHUAAsykrFCosTLCXk+tJ+
Jqpqc66ttItvcuY4SwCN2SGdi6jlllHOlcu1gDgRFb7XXAn40QtU3rZ/T9uFgZwm
17mQ66fQi67HU0V8UlldE0nOqNY1ZNorZPSLXqkNZnX5D0EBGxe8VqgF4fQvJTj4
fd6G187vP5bAbxSn4PsoPkSUNyLbq95c1pvYJOeKDHnUEAFrklDgZu0LjwBk5FVy
cyORmBb152wrOD2FDVciJ+a9CkZzlJhV7KEK85Z639KHFpI2F4daWY25AXGRNSLf
vvU2YDtLTW8oJTDWTvdvDs/YjQEllgN6u2gJ2zmC5nF6c+QnR4Q94E4t4vUA82Fm
xM6iv3NxUCckIDrH/Ye5fLGOqvlb1+ZrUE9/Cc7HSGdoKiLbQ9SXv53Kl/b9WtZU
4zywMKIGDeC7bx9SttvdU39DIPy6SmpJpQIsHVgaiJt48+OK2qh3hykR2VE08+qe
HpZVbAPtEJwYP3oVBBwWMzlcYQAQ91hR2OdMwRv1CkaKV0xw5CA/vuJiHxpuPBS8
/SHExXeOx+DQI8biEKb9+AiSrt7irKw9Z6FtqXDD6+N3QjCPHHqg9HO4mfmmmAXD
GTpL4f4R7cycZSRwC3gSCp0LU7TCsioNOo/VuBeoftQeEMkJv5uJasek8p7Whn4S
zIGwO36wOFkYdlQ+qvUjAZjtI9f5WstMvp5lRpADOh5OevALTB0BLnsYq794O9M6
IlSeRHRp7LygC/6FlP9kLb9NPpOZ0VemTwp5K7xHKBrdgM7hobPTIjLCxUrj5qOJ
G7U7QMLjnqYFcf36SNO0XYghhYfmw/jRMDofSI2xKI+K6rGHOL41zjp5Ypoe2J7D
i2sU6bIk7VjFt5k2DA4qCJLk2hz+r3S8YOqK4O6l12MGxg337d8O6yD3sD9Xhizl
pp7CknZgyEphWwg2l92RTd/mzXfTOOlLDeDxysovYxazt1ZLojWflmD9Yj2jeqS1
4A+9WRclVOO1M/Rv4+nng/CHtTaa5wa11qnOFdB+q1aCU0NmgexGgqWY9o9jigYm
G5w7+eSamjZvP9usp9d2DgyVKuupKqxg/QYGyhIyIbWVaexsYtwo5VBpk3rqTeNO
U6y4bzP7/+T5iV0hTKdfZWnhceVPhtJdl3NzCdBYSnbbL2XGB5UUoANCX6IaDcvi
PEaqt8yuAqdmOZusqau/rELmNbrn7joLUikm9hbl2r1M0hzdNW6bjZJ/ileDsT8x
7ZOVh+Htf/NjEWv/eOuxGuYDJ+oB4rMtLt5jpWslY4Pwt0f6MfH6Wbn4Ny5DUTlc
ILMyRsRtZHTG1sfCHJp7RbP9VrJqv84+kMBa5R/wRSYHpTVwhcehsicMrdTZaU92
ibVSeaotp3JFAQJpGSr83N3vYqewd5rFDNgLSVDJRgmhoevomvu9uB3JfxymCtYf
LG/59eeGPRvbnlrU8LfiwlwSM5/IdooF5FgLWpK70HNfa9HXf5V5vNKfiCdK9nxQ
WPcd68O8HkGtUrmeWc1wsJmb9cEtz0ESDRE99gfqgwNSNwzZ1tmE0RDgzdJksNpu
Ruvb5gx8wndMVzEpvEY1wroB6uRWhoLOch0LrcZgg4xWvmWVHq6/2UspaT2RCB06
i8SR+H2WoEdZR+E9iK8OZdcwmzSxJEP9YzOGw7HIBvE7gc/kqzf/wkI0ZMpjsj9b
cPDbfcxieeHuRb+q4645Pi6DplniM/+JKz8lxLOCII2zZGzo5cPKa2G4R7lEfzw8
DwfAkROcOsG2hbwchgmiHuXdf0CWqTU04/gjHZYxFgS74x/ZQL9HPHMftBjr3sJq
MvwW2m/KyZlIupeeC4UWDtSS6HLHWBJrs0X9xOQ0Bl35iV3NI7rGk7NY/pXP7W0b
gaoE9r9NbxaFNVC8OOB8mYxfT1298ztXNTA3sqhCcg6yv/vwS88atgHL/7TxgvzJ
fjSsqRx1SRROSF4/NKJYFXR2u1qr/zfARULo1k62hLmyj46waBfso6uALxULloUO
zO/tuG4hCT4MK3/Tk0SotnV+yrOsmrINMftRV9t8xvQQoBlxBZP52gwYLH6FIB8y
FAnuzDa+AgBj482j4Pk9W3zRdRXQJvhypHqoPzfV2NWlIlcF6oN0EBLhTOpJub8t
fh3BRGuRdgNsG2dWtRTJPqebrtWmrbCl7o13sLiVEorGC64QxMdRL3KZ8Su8eJ/m
sAY11zR/iULjq+54j9EiEQC5rkLz3QTF/3ZNauMff2QoiioPQCg/Z0QCAtj2mFlp
9IfTdLhTO3gq88kT6D/+98KNRwRV6fPotik9Xb6+Z7XSob6Fukfl+ENcPFisABeA
Q+HB00WV4MgBa0RBejeckihcolzw3iP/MDp7FelqM8iuFNBt6bMq9rR7qGITXrKL
RGvObCOuNm6RlS2IFuS/EN2NSw5tpJ092oa781v3iyhzXNpGY/Ysxral1GIempQE
UC3fRDGInuuOBWWyVnpdYLrsCaMcQhSz1GDGE6AGMXS41oH8ZaNXisnCW0/ElLHe
g3yhOaPrckyWx9aWygiNHLfnwCQRPwhgO51ZIZbXu1JC9AhdFxJ3WIxSM/hZch1V
PhMN9rwH7ymdxUKDZRHFcIApgTSXTUH1dl8qSNFRkCjedy1LjMCUK89fSLSJRzDX
37gnBmIOLJCyRYc8FvOxG2zYEd6GaQpAHS68fRNIVslDlEmTQoig/nvRiWRkozeg
ORacgEd/VBP3JfxMj/Ba9OOaHZsPgmdEB1h8W7mzJqgVFY7+rN8TJffmWiAtec6/
6LoBWX1hbd8pWY3YMKepAaEnfUbQO1iupw+yc4t2KENcgt8jGcs6teoLoN7cpe9l
a3oMS186z/Db1os8xII95NIDafOWNmt5QG201oq0rJwPoisXvQ4sO1r5qcy3qunv
YAPIoOFauL+YcQsV8BmaRvxc1EpIoFXONsy4ZZvHOv4tgrt7zbPgaH5+46Wu4tLO
nd2H6ZWr+PreLXCq9kQtLe0///buo9nkeRSfwXsh45lkr875HAGK+4Jm1XMKnyAh
v8q0XIBfKLPsu4s3eobDVtWYBnz7oErCCTxdrNnHVK9f7C/EMf+6YjSK3zlr63hx
sID78C/zCEkeK2wwMQkwBvGoUGEFEH7WXsKzYg0P+dZ9xKVE3ML5qbdmcoOu2bLd
xw+vLIsp2jhxjti6uBsXf8vfHweDtmhdwjncwBcij37kgjFmnutRZj+S9hWaWR+b
wABb1QCMBXZ994B6cUz9wdPAaPqowKNP5VVb08cXNxnF1lsyJwT2OwmAtuO1d+pW
X/N9liAf7HA1+oraA6ZeLooy/ZAChc0ZySBG0rSgmZ/C7HnoDbOrsUXMkxrnVy/Y
OZsdUyjVQtkCfVfilxM8XIWtnT0nCtE73pAwBCCWg/tz4iHwIPyFNzwi9edsyoLN
CyHr+QjXO9mHYj+878XLUjVhUe45e5n2fo9bT+UbObslpBvWBRVPoNibVwigdFWK
ydF1ISsCLpR4m35K7C/PnpWpOcB6NU2FNr0BO0G7z5a0lR9M9cB1+LAPTm00xNX8
UY4cxpASgcd1A/lQH4r0YRIIY5X0hk6pz1GNCn3tUzKcEXMZrI+N77Wr+449z9Z+
FmdsE9NdRdJdGYOR+aQ3xoNWyQfi1bZ3Xjf2xXtyJi8kOz6GMxreUfoxxJRo+Hhe
iItwHQW8e5ec+GS7lV1u5z8OSDd/+jne+3S/CCBy3DOJh52JBV3t2/X8laBBX+JR
IMd2C2Q2uD2OCCJTGvY6QtV+6SFq2fKZ9Bi9TdkmaSzlLuUwjcvwI7KjZwMswhhy
xCvkDvesJ3UIRhM/EdLo1fftwBmzWS5+2p+8V4CsnWYFfqtp/vMttLW9LVcGokv5
Zh73THkXvTSTdiTPW/vv01kPlxsTztNi4G+/CzOA81bDlBiA9D26oM5uHNvJPHFE
TfqMf5yOFawTZTJmSdKNNXxUWOMiMyWsUkYYBzl235eNNyP+vsJ8+bLSTLHyfdPn
q3knOEw082T2/3JXkLZPcHR5e46/nQ2X3Q+YbosDz73BLVXMkumIr/D7lecg/UCJ
AnYa1zyCnNwsxgadbrDTJ5tG90MAYGDgaKPjGlERI26C6IB1nEzYH4h4DpAdL8Ix
HVcBNyqMUeT8Tt61zH1LFHKkhTapRKLz7Cy7qc5QMWVyn1C7duz+T38ncK/T8AGJ
ke3FiAWr9q6ujNDYsRqsviMMlpo4G7itUCtRkw/XtR5diGLqBaYi5EFmwJZpBtkL
AnEavDYPBWsQeFW24rajCMo/KH+y9g7SsPDZwCubEPk3MarhJdsQN+cLKLMlnrlf
d0f02o6yfutJwCGSSYiThyJNgSSzpc5m8lvLqXRhCl1yI5oupio+Ao3CliKw2JS2
lMkraHW9PyLqvD70WsD0/JwgnxEW4K1CqMPtTxxjcZNzqGvSZSrm4+BSSob50zDT
Wdik+2JoAq3zwFflTBd2E+8yAuH0AewImA/P2frT80ZyF+j4rWPbyvfv8rbxxAsW
TTSSmkqGqZANCdxypOLo/6JeoJ1KmRhTFaaD9+n3ecZQ10vcb/4PUQm0nHsm6ycu
p0yQtMUNVSZU6woMW8wJdmy1s5+UrCat3GhIrs8eiEFvsMeLCv5u60BJZHrte1CR
voJoDB9vSC87Op/CxY1HCZfkTNpz+jJqD44UTET16jxqikP9i4JbOGLHjTtMN1Cn
velxA4l9fziWHOWrfTgXuI/6oSHNmIIjw3jEL77qev9B8ElA+WS4bYz07pTeYLTg
BAuMcFA91ETSf4wkrxdGd5J+UlNTKQXiceIQrF++NH8rFQw+j2QXG0ZsIrO+UiTp
BEJApxQu/hnXe0LpILkJgDtsWaBWG/cBMaMsuYzZV9UoZ1CfXj5dnr4Bbb9TV0bh
+mi78scRrhjbwCUQ1hQWxNN9esY1D6XJnlbE8oQNGLyWhgyvv2Bi9MYMbz/N2By7
TqO3dAjioR9rkvIInFovUUUBs6xNR1rZuZmQP2k0D0m/MjUak9ky2jGR0mGpoyck
Jb/9x8M++TQWBQOwkNoo6Fo4IX54Nht7CxrDdGzMTX92MYwEbHOMLgB9eM7zK4qB
2eyihqGVBVj/fs4uOlvPJ7RydOYbpmOHBiS35HQRIJp+mXrTWgrdJHfMaMm8k3vK
mRaTMO7I0Jnjdrwkmfo/ZCueqox1PRADSsSiT60BJgvXo+d1BwRjIgroJJm3W+hq
TT7NCoRBWb+obgPNj8xjmit/a3QSmydsG1Gb2+PVi0aw32PTnvg42ugBhiWOb/c2
ZxjfVXKpBOF9C4zjL8WEIL/qRE60QA6oHCqynfu9qcFcRMtNX8BvTuP59ZELUmrj
Gv03FF1VYusSTZVC8W0J3rcf2FiiNOTDd1y6kxfPYieqOaxfPvL866FfpAFI8Cv5
4t0ZoXF9cQ6huhwv8XLprV6fZWBRUgbcDRgSBOp5IRl2QxAJuqqxphHKsbhVrTfq
ozjSeYvJrWFUjDGDJCuLk9HjU1yHpQCs0vQSBzK9AQHckGe1/SoO2/fIJ5vaYy1s
4ybN3qbvF7AAuBJxO09A+zhdjCrXlvw85DFFuQKVZHz4I9jRUUiXSzk/J4KL/ez6
NBDxa86ay+/BytHmvkH6Wx/8yePh1DIdBc0NFvjcm+7heyfd9F+aesI+g4JREHGF
8aUrZmNpGflnLe7wcvlVpiQ3/TIkhGcYsn6igL6d3iJXgJZBog1/eMXh3Kz8TOuS
svW84NIGUTIwksCFmwe+Pao7uv8jhSeKVWjeNboMXXie+Mumda7oqazAHQOy1Ra+
PJ6+jkQmPephgU0cSrYbzb80f3mFSkwwpfA3aWGApKZ9kiS5ORN4DyNQAtubgFu8
7HK0hCUTBLgGWAbYCQtT4eLOlQXJFQKmQMQHYVTtFXsWZjP4rp18V+lFfC4pQqpF
hr9V8+QkGdufV9FU7WlA4bZKYI6njXHer7pvZ9VEdYGI0WgcP5Q6yLFmdAORa141
/H37W8KOOlbaJ+x1SVggQ3nEF+Gg1yl9KFVV3i0kdWit0w13dqUlbSYOkH45oYmg
VvgIPS+szJvfqwTHTx0k9QGDCFr1uIlSH914OfhdYi8CH1+/ziQjJvRuOOUNeanM
wdNgYkpJxC2SB3dyYOoSyl6QcKLt+wsTAihXuGV6J90QZr0gvKnMJfg4SxdBxUa6
wC/SFJwO1KssRsUrYVHHlJ7eAoH2rQpRjk7ZGI0iqUkYSYePiKHCDcidN6hz+PUX
7ZJZcPQw27Jqy/6dT/GU+eC1fOp/pJ70R48lwWmjYfmC5FMiQWm/3T0Pe60extlf
vbDiQHPjnmKemaX2O6flOLtOiV0PqqcA6ssROGQ6FOIJHdhGPJlK3rSBuwbBJPck
4mhzsjfeAjgEp/FczSiIq+cc7JZhyeDRkO8Bech6YUv2yssClBsRsBo2z/0aaQNY
USEDqiBhXvLxQZb6gvcDTbTOZXLqyiG7j/Ldy6aPvcIhkH1XeY9lsiIfqEagNwlc
n73yrll8l6ji7BdkQxyuXN53NZQfBOQcsfJZ3x5vH7cm2bFywSLKTvCY1AdVv99I
1KPHosepJUVAKQPgibJQ4MEKzYJul3eVm3ThXmxQdoVk1w9zNhbcZp2zIpsobR2d
6DlnZY9orPn1krgvxrSMMCsavWDPObr8vxzgnxYujtmf6r97IDRrB2Wu7GsZZVIy
Iy8RQaVMoeTv4WPT0lHc5AjumaAp/p5DPc2nMX7QzsVZIDhPQOijOBogB+iKCb1E
PjFMBKAEvAaBOMyhA3XKQwpPGAvIsOxjU2Tx9ic2WPrX6+wh2oKqEX2O7EVhEoMi
DA9bOuRIMP+NUIuFP4hdqLkc9zoODCRZdHqSMUMWketsnn1xAAzvZiV2ysnJYe8s
ZTACJL9/EN/bWOIacHoJ2R/1AB+ciCqb5G/gTTFQmLGF/WOycOzy5fWsUYAqVBvE
HKJK7RtVb0NWq8TNwRgPRcQLAClcIB8oyRffQHLOSAb018YZJGX2JJ20TVC1hilk
0oDFlAhp1OUVsIF3T1U/+IMXYTVJAj6vNhZPG8QXavAq/fL9xwYx39jM/KvGVIDi
XC2eZvjtHv7+ZEhhN6f/GkmGQmVwCdzHiifTmCADIR01v/VeaX1QSf0bce8fMmjn
cPTjitwwwdJKe32KkqqEn3Ynl1ns3tEfNrBqQnCmeC8hpEBKFy/1cYnE6hNXk8B6
M3s4yHJoOs2zNXgjXcUdbA1Gz3CtL+J9Yg9Me1441yhJSTwpG3WnQnOy1TRzlHn4
1YxHN0j+F55SV3XqJe2LCViM7Dw/W0hUgauMs+GTd0jEFdTtbMFDTEHSeQh0EX+E
u5ozsJ+BvGykaZ/vNlew07lmvwwXvrDRBibW227gLt41hH2LzcfqUU5V26FtWj8k
I7QdxOV5Fz8UjdjOtSBMvTqq/J4zRyEX7MIt1v92A5EkKtnh4qC1eJCrHoWedIv7
FnPJEcQkMH37BQGkOmgn6C2LTlpoT/I7aNTmk7Ij6eN+Bpx9bySnSPc6Q7fAEORb
fk9o6c7wGPZyjwQBdzBYNbp8ONUMnaTcE64jk7ChtdaF/HH2gimpThztAYcFyJaC
nVvi084f0raldIK/YLfShK1emh1MyL0yYvjwXMczfCoXbxIn2ho1VVzw8TXVPPUS
jqTAtIIzcLoXCubZGgtzEmT1GpGoTbt2ciS15avHbopQIvlPvpt+2ST90RyRXC8r
xB8+6AQ6QKE7OlQsJiXcKX5Ssi7FVCyu6sGNkUD8vWrIjSld/gXlQrpagwbgbiYa
UrMtOL5ErRfiXHAWogaqNxhYQyr80asa1Kuka0nm/CwQDmD2bs0oV8LmAg4KagNF
ZKYpNKtULVT9JzmOcSJJX0iDHG6gnLUySwUrJ8wFadg+TQT8mH8cCxU/4lo6YQuO
8k2iPozHo2aLKeNDyQyuRUTvNGeA6G6X5n5p5B3Kpa0wm8Lyso6HO2ELcafKE/Zs
wHj8IAC0Jci5aNlqxeX4iHaxKKctOYy9XSM+68L3BS/bKWRVlpP7EM0Tt5U5VoC1
cbnArUyarmhDf34ouWsQqm8imx5wY4LN8ptRf01aaVAiAJ4jOBKFt40v6t+qa1u6
CHDUK2dftK/+/9+MFc9x7dn8k7M5YLpYwEktGDo3Gg1Bg1w29d4DiMQjHbPi35Gr
qxIA6rbmJEqTTC4zyXrfNUiM+I/mBrezOGXYcRIZkSHdNRznKY+rVlFUqRdLwK4y
R4wJxeB7+iRk6BGk8Ay5pho7YqQqeMpkJsyR8TDn60StAmws07w/DkivpyOWWKei
BoV+n5KT6o64z716DoHHQPfA3brSG62WDWH423mtUbIGLtNq+jB0MeSCZxCBAEsn
mGe0hZWxWsjMgOfNeu5mj5utlNpkz0GVkj5/ue+hTFCiHVERshom0QtwRsSLu41d
cpJ3jrQGmo0ENqWF5nJGQvsslKxWIeFmbRI8KOmmZ/+BhaAJkECy1erbHLsS+BNm
MTkLlXRlKYcy0k1itO/MbbRtVsb6T0xLt9Zqxp3OSBEijWU0GQe+V5XUbY5dxTBq
r0Gw4TiRABtXZLKvwLMPAB3g8Z2bxAdpUNa2DViyy1tKtCpE5J3/krJYkvcgEzkm
vSoVveAtPL37WnmJ30LEZb566zPGBVG9vKvm+OH9W9F23KVci5YZZHn4ISyDS+DA
yCmrIpGw4WmVNlZUOBl2N7kEzGHEVbA4lCj26IAIjt7TMh8A6cUK603HSIgJoWgK
iZskcOQNs5S4dyJOUSISdmLrPda6MQV/fF+RNrvl4bQnhi85hOymkJCvne0u2t6+
S81armBYLrTpjz4XdGpKXL6PVmAZHmng/Z8FXPQB9p1k3B8hVKjnmCzLk4VolJE1
j3oL48n0vJKYCpKqSjT1YXg/fYK8NtSb8Qk0Dx0wCAw0obBjyCup9VrFSrxdI5nQ
1B0zYgKWp8dy5fJ+zsGPukESm5PGi3FhczbKaAOCSbbhe6BcmBzyv975w7HY2pNd
OQhWeeJoUrLMGIsWdHuZfs9hgswUgaNmtfPMSxi0IMW4C9jyYjfVOMoVpvxhpzkL
BCcuRfMRqbII8u4ILiRqBtyGwHb8yfcyKofnbUAHdWWl7jFFQ7Jd0ZyeWMLAvuct
E+q73gLjd6Mmfm3mukCpeCi6R0krl8xxdAbG1uOz7BUJVOhkwgrwOdinqLqoyvfY
syuTRDe143+dHu0aBy0A7aJDEVdvFHcGKcXDO8WmrQfUk1C4FSF/D3ACXYZUOfme
24+nj9jXCl9ly2QRr20hxdUMHwc7iAqnhKVNb8gei7wsscT2Ate5Et9ZzLK1BqwN
XPQovKMTcykSsovyENhfg9wsC+HXRc7LRhFJ11ZeYO8mfEYu4oo/g7wEg+u+Hkj/
3eRoWlDVtnDggL3PGOQdPqinoC7fMe8w9Jf03xbv3YY0ohOrVsMLY40Dv4Dx3+QD
euph8b0WVjeKgvPZEbE6ay5yrMpGZPpFB1TN+8gxAXMiyMbfVtUevhJyGxVFj/U1
BT1cAoyqgOA5IqSGtlEv6Y7ufdrwl6cKSdLigl/ixNtZIbpxZQDzgjiP7QwSKdqt
oPn7Rx9hqZMrNc+LV6mAMPel/r30rKQsieOg7B2hv5wadruBrjKQNj70PkxJ+9kC
RiN3ASqFoebq9G1hs4rrtbwzuSm3o9BA8ygQZGAxmNV+l5v5eKsfvi+1xwMR8iaM
d0QU/CGzdTC1KQMsysGXYKCDYUC/en+sUNiUge7a42zyE2ri85mNwaGX1TlV5hKH
syLSDe75CTqIzYiFDGkwjdJ8mV8P9cM+8VNEa3AGD+WzYOx+Xhn/qzEhJUwN7Agw
GXNJn3duPbnbRCR9yclzbCU90hgER2yt9KJz0fH09YN8ZmoPZxIcXcl5QGHLUaP0
EowKDKbvL9207pg0lwiddoexUswuZ9JTglE7pCHZPufDd8cT3Z5xlG9WdOMc7VzW
O8KyThJCzawh08buyC3kzXLEscqxnyF3sJHBzN84x8cfEr0DuM0Rrgyzf17TgLvK
sfzTnQvMbfz1A2z5knlYFCXZHOJwKV/koR6xwFka5K6mTjdsTyn3915LaXyr0UmL
b6w3otuUTBVfREfqG1Ou2hd0STRgQ9XiJo2jR8CaITn22h+g+jGbyKIKo/iU77sY
dIRA7Q1X5TRBeCKfiqnim8vwRv5BMK8K7NGLNhjPlnhPrb6eyzKP9hiZe4Lt3iiH
15+iX10N/jSiEcXW7Y/Q/JDX384k/5i4HAjWagMldPyU+2j+CXOciK7yLK+PcHOq
dcaKHakSgT1QbFRZkOyTOo+LhHcfLTFOLqs2/li5koN+08Ew2Bn4PqhIqHf9OZGM
Vo/HeUxvQb0oSQSurUJwiz0iGWemhzmMYqlZWRK3waeIB9bvApGOjW7C2dURvQ8M
kxyYzvjK36+7pYc60bv47/C4mXMSh15nQc5BMb7e8XYelmGIa3J29ne+3eMqE2Cf
yxVCqdtLmyURS0ZzwvfPr/6ZDVR1vAyK80mn9Ic1EOl1oUSC5+P5KX7+G+98QS7a
4BkhZtfvazXdjqyOz9ZSyZYZELgRD/E6uOGSA330PXyrAsVvoy0Wya6eVO8nfGdU
So1jWVmSNW/Nx6HuYfsiz6K+LmyFM0sAxoV2pXuuvBP+MnaJbtyZ8jy8rbKU0g10
4Loc+OlgOv01xS1ETiu7M6ClS4VHHy4OnsAk1VTPs9WEZy3ZfZlmOOMZLuOuJPnO
SESc8V7oIvg7kV3Barkm1nY2jTNj3vEaWxX3VIDlQSENewf+VIsn7p4kvM9U9aRd
MeOF/yVFLbzCXH1FPPFEavOjr7uOZkkDr8jtolkm+Z+5EdlFc+pePL+7hdiWP3PI
q2rx7fFBkfMGhPjERcvxQc1Ouk+QFP38A0CYi1VEuY0DsOIMZ4R9D50hoNCKJHOH
d5QnyytWcl8MM2vKyUgvV2ovekkR4dDy5xJ2HR35Vk6pOzo708h0p4qLwkoqZ6m5
sRLkx8rX49aSdvi7EoDppjcrTAI4oBH890i5rjZIVsj6cojD22s1DWt1617JaW6Q
f3Edjl4rFZjylCpI3yCxLiPs/2hNbcqoQ7Be/5HTqC3ZV+nNSwD7bGcdkcee9RpI
FDB6OhM+lfn4u+4PqBw9g3O4hUOpTbC2XeGAd8cOgesT2ueR0ocqvL0sbY6Vf+lm
7i8b99V/tZ0wJX8FFLs73oOc4Eqcczhdo8Jf5jZk6rk4OW1PCQHqAd1S4rENHRv3
pYJgh9ni4ntC0xZ0BKVS3V0aY1PZwabzcattQA/eU4BpMEsRrGzL7Uam+gLjhlnh
jLEDSDxiNYSy1+dj0FvCbjVpENQvG2/3kkkcYx4XKhGe+vcvZNKk+XKDeRrXxwuy
VZW4xvvAG8h3U+82CCK5Bz6CPHnL+2BTm4Y3jCe4ExxhESN7d1yIhS4VwNsvQ5/O
Vquz0N4GoYGY+pblEztDVlfMPrU8Q05+BaTOGCWbPBSb+ltf9MaS6Q0dib8pUZ1W
neqZ7fIPM9gcsC1+iANsMIZJcASlqFJ4enz5jIvGyPwI5ux26KwgDFUv714Fdw8U
+98F6h39VUpil0eBDvzCqbkadNJ2V57Eq8NkWiDTHn0ociFaoPvGbiJyaTOwVasV
KACUH+L+EZp/1dkTGctT9tgvaOhIqOl8FsuofZZ4NXT5CC6u3mAiZ7UE6AgumGER
4dOlKQltI4Esxpp/iZoLV7AJ6pcXmcLJWtmVOVSHF0wnJaL1K0pte3elVnVJiKQm
ak2f4ifbM6q1sMMKC7M0fjGEzYEWoVuXyPUNMHdIfY2/uiJdbgpXN6xOUjXwhXQ+
k25UTmd+BRnkHHx8HZDhddAWlFWY9Mx/Fyj7vp2ZmgG7BChyfQ/YDT3pilp6EZLJ
nIJDoCjtA/uJ+QyjpH0SOThV2hC+hjlhF/AJBAueGjKzbScuKvPtXIP6iEVWtAmF
pD2cQ+nh0Sez4sw0kw9h6NriEvn/8Np82xFrUz7WyJQ8IJC5leq6Ez17g2xCU/r4
KUGLjWiQrJRnCfeGaU8jSqLmRsk/gsw8cvoAz6CC0+Zh+fxEKV5O0l40PehEPRJA
IL6aXjgH/jr4vvk0L9l0gyLb2xnyKTOvwJeySkPGP8ZXh7XlH+FciSzHdzcCgf0d
iY2ZEzwwgqhkvrCu5+LBL5GxzWoQuJpsnKC6wctisVdklZlspamUFBF9BPCvQ1b3
0hBrlpYWqb/fbkIBarB69T2Yrl/gqAiESaUvMqquFZyMcwedlY9O7ii+wy2LLqdD
DvuVadRhKvw5/ChJ7XieFb+setqqoq6Na+uXXX9I6ZzltbinvjxRNF6wiCT8NsAC
vs0RL16cf7j4qDUlwGlo22AnJ5KTH0/G8xyhaiAL7ZxjT2v7qR68NNP+Si10NStr
bFLr78A4MR8RCBN5A5ZAF1savf2sv/agMbi+f4BUPGCoC/8OStCsW/geiicoUAMc
OH4RZZTiFj9W7grda1N1fFBYBe08a96+XLQYz7L/fp6MW/IUi4mUPYBq4Jy895Mg
7SbWWSJiSF0LG0cmYGJQWJrU1ck0X1fklsDwC0GhcKH5MwdQI5jyIudhfhlshb3b
x41fCZVIjiMRf055rYg9CTJNViNsQg9oFvWADv70Kz+e9hHuawBwgETltRqyXwMH
5mHeNAyxF+b3JLPRYOX4D8uLNe0+GEkOC+C2RLK4tHui809BD9yH7fI56fAYje7B
M4LhqgrwrxqESQIjAz+HVjXbPD7IrgM/Ct4qE+TlLhu/mbdCQWCBiC+tS9LjWWnS
lQsSdgFsO8YhqOV2xSbrmFjdRSBGBXQ0wRzbI8QD7XLm2tK3i1+nD6FB5r79ZXqL
tUV13YYs9UDky1+ZcsGOG/xCKl9na34MvQ7KrPIVvspYJoMMups91b4XATxA/14s
RYwzxid7GpsqQKfshTF8kG/zcS58GElGjsny5ZiEWUxkOunVkRkuqNAxnKCnsBIP
dYG98CkWXzvN+gDaaGqWmi5QDUXUft2a3JXytj3jYUmQHlKw61s35nDNaxO+8Jm+
kocpoABeYrbT7haaHoOSf9tNRFy7NVI2XVd/W/FD5Y5OtBXxZG5rSJYaIeFNmBkc
cEe5oThRuueFBfvxYIDYQqL3sZaDuuddWtqvWS3CcR7W4VW1xPkZZKO5dT61+iX0
UOQZDFZivrZXjcqtGd8iFiU35AS73tAuYwdhCow9i6NiotvWMBiY7Mv2se7pHb/D
TT3KAH9ZKTtOkGUp5GbFCfQ61EBn7Vhu5ezLfcPCSIzDZ0oHGVPOVcAwd3IrMeIG
IAgG/vQtZ76xJO+ZOPWonBEa0519guEJl8YMByBAdkAaf7TG8h5S8oQpPCsTKWAr
EtF/sQF1xVXZ7dtYuGnpi/HjrahfZl9paoXwz/dRbvIb0FXZd3sOh09GVS/AgnoK
sjgezrUKjnGVgHLjd2ZnU6kNXU4gQ52L5b/pM8qMNNiZc4/r7hWNM0byUBlVFvtO
POL4iXUhcKPCBK53EhphnpccROzQ47ksVy2wbwcavAr1pGw9fSkHfjM2tBOQ9PIu
dc9hdv7g08V4ncr4H0smJ/Ysd4JJZYcdRBuQh7CXyHimtkhTJOSk8KFSqHJ2dlqA
77YiP10YEbBLJJe7IGHQn7vzeIY/jguI6uMQgZgaPIJE6rVSeOWgvibduRr4pqsC
ynix9ovE/WSyTZ6kuC5FH0cBMwVmfRf2T0BtpXK6l+KFJp+Yl2G4rt+8NJb7rwbw
s8hAh7bXbeI+q1oPaDnDJ/0ZVYJZ4L1Z+svBWLdCUy1NBw6tPGBZXQaZCDY2gDsQ
D1o3Y7EZqfvc80cgYbr/fT6Z7nU10WdhRI9W5Ks2RBfZwsDIY2ZVHj0hWMHeDFD6
QHw4K9CjXeJWWr6SARFiOB9wDePrvUFk5l9cA3KBdHeHM4X2gsk8xGKsAXj7Rsm+
ONBNeswDV/Gds37hoyMOM/4AskU9usAx/PbJ1SdwoVxcEmukz9/e30MZE10CiNAB
DMnvKts1F9IRN+aFKwnaLETZe1De5A/Tf9/HlKnNjPBiZBjdg178imYlF1O9cFHq
xhF0Eaq1xluQwj/AWV9nNQqSsje9gndV1HKKAS95tTPLSPbQy2x2c7a7OU0kbfo8
jbZLI+iyHV0SRCXH3oBVDWZNbCHsuWiLDGMNy/CunPnOhHVgPOmBp0quoni5unqQ
+vP7qL58wKwavxDk9lOVHssSCiGXk9e21Z2tVexnskwwEFS3ht2IfXycIlhb+8GZ
96j4IffdtDhoonvDClV0jxi/xwYe35OZ7eJFmN637GZ+MyIoXDz3RrxqNZRDD1Cu
cL5eY4tXGdyjkipx0QM6RQ9y8sak8jE8NMz9R1yaqAXnDkCdu73fGNqzmGeGpyum
Q9xQ4XhU1Kl7ZuUKEV/o7kGnIPA7ot873RihAho2owVNXTq+dlTYROXySTQi7PUn
dYvYbelIaiHT28uKTqfPMrStjoiP+4EEKjk4BSefbXRMssCnvctIIktIMNaqbd6K
NPlvpXuzWP8Vc6hhCJKj4B0jdQauqAhb3lZuj2QnX6hhsZ/E9O0fM+VpNwVcL3P3
J6Wjj8QjSfS0ptSYWUKYYbd/2AsNla/CN0mQBUT0eHsqmgUzG7Xt1LZU04BpOr23
lohqKl5EcgTMEyEQFU4TfPqMN/Up+pOwckiCQJZqokBIAKy4rmePq5RHAuTiB/D6
WqkwBmH5nNfP/AngX0jk33oCiWMP2tU3beHn+cntJ7BC9Gcj4A/AMPc4poNKqBiJ
lZY1VreUw3CQubJt9+7GARRMpnkD8prUcKjYqnJmMAZ5M9NELsDk497Hx6z5rU+P
bIFonfnLtRMBnUxmXi2x/71pxSiMpoJiUHX+8O0r0l1khtvfU3h+0aYpSRYhgstd
KzCnIqzZQN9/9JfFMV6b/ejjtkj0Jhb/Rgx+6GotEBJ7cXGDP0fYl75PZjWR3Uqz
AqHAhhPRAYE/D8zc0OSIIZm020x6MWnMByzfAiCvj0EGv8C9kydJ57I4QKHPJcbE
tw+swZ5Jg39xOX/Cf2GG5dVSY71Foht484FTVCmQga5Q6Xec4hegbvHJjttbf50/
6pJGKMgH0hFwJcUREMvF1yGmkt3fxdAEvHv/9DK4oi2ffSB61nPIguN0WLJBbcpI
dRBZkXqaQomPpsD/vnpBJIZ1G3+hMxuwD08PjvHZud5E1S2XEIgRju+ZsA4HJK/7
qXkZRGQWTaHhRE25lBb8Lyo05ifUT6Vlox+r9GK6xtFrhDtCUUm2IB62HmJiSp7b
eWW1dHWBtxSDnGNx0Pv0pRDt/mNCRdsqczjqMXr9BrEqb0usg20Mcms5ey3anxgp
g8VOiNBVwl+gHS8pPMoRXzMpx8bZW9GpOyJgnY2ZbtF4PYTihQRSne137iKHHf4G
dDO3JC94umZzMSZa2Q1UYSntGbXlhgkX27K9CX6Vj7DcFr02K6GwhnIU7Fqf4BZ4
nP+tA3evLTuwmb+ge/r/qsukCVWwugeAyhfLoqarVT4ncSN35nS1UqayiZYq7Lzf
XuORjdQps0+sPxh5PRVqjlM8sCEQclHdmoVTmMyMkDUq+PL1WWiR7FQ/lsV/2vqw
0pirj2XGn/fBOOkvJcz84r8QNikDFBZJ9DXpLzsYgjMhQ/9VgHsuZY4ht+IERZ75
xHbO8h4qzTIbwocdOmWGpur/fKHvTL4oP4ipdNqhd5B9MA3nuxjJ/IUB5PekgwDN
zcFSNmFGUENeVzNpEgc3c7W7Q1d0RrqxFAMak0p+flWJZyBaYEvs7TjXrYm7tQY3
PmB6siBZVvk6ILjOETPJ2fHxUdSZbJCHjI0va/3wHW++smVcHkCo/6GEZCjIKKgV
qwgizu5HuJrKcDFI9uROWNOf/o0bczeNobhP/IsYqQiPX0Vq/Bz13obb17E/vyS1
rKa01Pr+VKEgeLiWdf1+nUTaNA+VxmlOrT+Gi6afre9Njj82PXcSa8vkBvSLqfCn
P98kdUQEv/h+xhv9PRiAr3D+z03PCLoMsFbsNUFPC0PKsjsVqs76I/VmzWhKiy8k
JDqpJ10z9TvYD6ruX2TeZv2Ef8OcRYqqyV9+La2R1gSLLaiypflnvQ1CpShy2BmW
KolB9a7kntQveJCLN7b1+sVtV78Qdp0QYVs+v+GBXZgTyQA4WWcvcjryu0g5m4th
3so9HP3Xh8+VJtH+wBEFfk09Oq6Izbty/HjJizugFAI9BgBG5AW4ScRSd2DfEd1T
jFuhJ2qAUzcr9nIngupRkuOlgLmyvmOFFdoc/FAm8dCkcPNE7DecGJZDVbxY4Wwq
ZelLBwtpUJTy8Ld7iGUaclwFfzTWO1B7c1paQax0WyVCeN2tCs0cpXY35v7wW25D
fMPH+Cg31AWZv7MCgcoelPKrcwkjPjjauCKYYDwEz5YV3SVwfak7fKzY5fa5kxi7
2pIamP8Lpu2coYtJ3/+byEPCvR/0cFi8I8Q0IAAl/vI82QqQWMOpHMQKoEfNcrqs
YqqW2tAalM4qDrMhchtXH03HI3MHUOaj3+gFaHwczR8FDS5jDKg0Ic2AQCW8jfXf
cvgNRLSNmFyFDDZHq6UJWJIITuv0F/85XO97bzcGVqE0skm1Pq61jRiK3/J03ppw
HQfSWSMWD0ZhNNFInXjkyAR1fkcz02JvfrTO8BbBAmc1/zYaAs2KY7BIZb8DMmqs
Atu/H/03DQQ/6ARi6AQq+hJ4MUCiGswdcSINiQ95qt9QbZV0DjHmfelY/p9eT2sL
ZXf+bYQovvtk0L3ec2X2hGMZ1m5XIUOk/0/XZH0QKcF+iItpxVCX9U98Re9slXKL
1bXNz8YYXZkiPzYaqoBbIm5Nd/4tPPM7trDCJNTiTmWh3Yks9BRZ1FC/lAxZOJEe
h6zguh8MiG+w7tue+xQV/jsgm1uXde6z/8F+fQMYXysWZi3VvRvHeHV7/mAKhRxu
8ih3ktfqoeRv/t+fMF9GiBaUdS5v2Y85F/gxVHd+j0M1Ie2wl6oya+pvCT4zzZMW
+o7k7sVmhqt3zkoflQFxLkKABRlo54DkmLHrH9ZcIrqpkLMmapdH04LRoZn9BT4U
VeS+Ys4wcXbdLmjpAV5uDv4pgYeD1fYPlVW8O6cmasRvA22zuyboptVmEucmM503
9cbdzRQaKaYzcqgYUdH2ao975BDn6MMjTtHIPPk21RfSliBoOgSBiNcHH1u8HNW7
LicAZ+LH+dGJYCAAOwK8ZCBOhPFQdcN8rt27BLr+l5pCedcl/4NoM8ddn0SItJus
XH1Ma+a+7QnMLr3XFPcbGyUoue4Mr7jlZC2T6HJj+Yidlth0tXNf5JAf2TiQkt+5
AS8ZqEWvQTKcRjutg33WpplNRLwSYj2YpZISIiVAtKc7BflXj2qtsQhraj+8IoT+
vFTGiUhmpKH7MhL+o224uSJsQDvlWRtKnJ836tjO0CH8Uq3o2rWPMq9O8d3a2xZ1
GhxvKT188VMlmUMadF50pZSrfkhvG0nIfDQI82JSrKCvl5vDplgaTQ+aau/XpMXE
gADs2UiMZdPdidZMU/hpuzYN3PxqkzW23tVSO5Iv7+K1b6Wo/7jpJ/OPvM0pS4dT
0obF04VF42ViNj2eHSbWmM3C5iG7V7cL6jNZqGaKAIlAw2mPRTVw6peVb9QYo6gt
FeVA4G3Xt/1lsiubapvoq1fZleLl9X3CskVxp9+dVRoTB2GdTHZ302rbjWqtx8hU
4XsgwkYgCRmWJhj/GZMy9JbU19NsNhYfhAVC6ooxx4cd+TW9RhOyFn0QVqIv89uE
GeebRm+zDC19N/fUW7nPx+RLozYuUjewcSX3B98sBXDC/10lxCZH5yA1JjJofuSb
9TTOE7cMmfHj0HRjUOXdYohqaBjnOy4yt2pQ+rPJeZKQQRHJqjQOZ6XxOhQi/x16
tjjPC3IR6f/AkkZ0+YVC10Nz8Ysi1DbMdYrXtM9ph3sjYqwwJ1+LXtQD9HNwHntE
HmmyI5Za6HBZptGsu0awg4veBqWnE7Obro47vZwohKkTzcXrcu2G2kTMv/xXJNNi
w47iwqq2fhO5W5wzfJc+fIqDUjg7e7iAugr89cktnNE3+T6p4cCGORgTFG00CKF4
nehyJ00gUuEUKtTnIIUi/U+Eo7sPglZs7e7dnY/Ib0Gk9ym8rWi+hsgD7WMvlM2F
lpniZFZcmlo5imzskMJQ7DY5NY2M/CLSiMYrfCfZvGQTrpJE5Fw98vjWbAwKyq8y
DINN3AkfoEqzDu3DUYaG9Cym+DGPTXHXg2CvATT5ZTD30D4yAZI5SD2gdMskGxHp
ug6Tl9GkEEIIT1sOUw+7s3eUcrDJzKUjwkTWduE+I4XWLzSzVsXDVQHa4k0YCZIc
V9lq9/XxZ1nCvUg9dH65Vjj/FuWwM8ASnl98+QEN8FbfLBmLvL/a+e4UBA9k6cJA
wUKh9SLoAPcJm9hpCRNvVVqh07MIYmliKIbSyFQ6FyNdQtzVC8oKTQ75f3QRMgYs
GRY68noGgO12bjcupcNeSyugPP9ANOtm5o7mZGzXN1rdGFDYt+ZKzbrWeddAvOwB
9zHz1lZ4BqGsI/171eH5B6hKNP56LgV1Cm/KmturH57pTauyuhlKGMG5f3em/eSV
zXaCYbSaQVVCS3L4S0mben+nyUNhkgGHmJsKgSrmKLe43lmbg2emzVd4ujih+K62
QPBg0xAt/3iRWcybO9Tj3dw/QsyUdGSbzcXRV/Q4Mqa5dmSze0Kr16RXMWvPiJ0n
VvoAzJX9Yeg2itw6mHcDbGSB9W7Uix8DrUy6cIq+B7unKG5AuPbOm+z/dbPMjw1Z
TvmXMtExO9r+M57L06H+JgHUselz+cVodJYRSGwS36LJ6NXn61q7m2vL5jzUWl9B
juu83OFwxG6wRr4yiIqja7w2ds/LGlZVH1VpJizUVVsp2EOHGjQKRtwjc/VrUvrq
qZPXhAu5YZUEwmHyX3nAA+d3qKzimeN76JSyb+5mRtCxSAqYnhUB8PTlLw4jm6ep
8a8tb9j2ImWz18pSAXFA+LOye4R0Mz6fPm9h77ujyLWrtgavpyuIafYWqyVqEE3g
23HqOF9mjll4dl8aPjUjbx3jcO5z2Mr2+L2bl08nNH7Y64TPcpS9YBKGXF/zABf9
+Waq09+F7v3Zl/957k40a1c3318QFrkOTipvqTW08e8wOlffFGqHhjnuLWDKaKq4
LlPsXm0U3mMMkS7Dz9VFmie/7VIDnHoSZef+ZfrNcl6qY6QOfZw7QBHVOhwr3oCD
Iygdw6DVqT27/bwLEdZIxPMyG4RWmUDF4TqzPja81NknJd5Uf9waIcUCU98aIw0e
x0odTCYxDUoTKEn0vfhflQ5b7YwX7rlL65VA26tnj+pPNtnLh/Cl/hQpcifal0yC
tV6BZ7SQtDXryg2DdsCmS4LyPFd2qKBvdV/xo7Q0XP5brhSSzprEyB94sg2Z1z0k
J9w8np1qeohku3UmWylssDE9cbMgDd3uq6EynrBnm69KWkD5hCaiftN8/71ay7uO
nryk+bCZ+iy1Ijmno8YeSLgeRyQMsjmwDNBG0SNK5N0SW06qtpI/GSwbeOcgWdZq
ncxHaU37P3dcEIjzHXWS37XccLyj+MUawR7WnSfxjkCOoua6jncS+Qlo4e53cuZZ
jH1x8FkZX0Vqa1Z9ZtARaBqkq/aOQE2BQOJEc5po6FswP3IbDdbsEiUOGvQQd5zl
1KCgr34ckSsLtnvIcidJNG8B35yuZf6b7Kit5MhGFizCqAXpIISmTd/OkGqcsRdj
z9FPQe2ggviPuGQ22a3jM3WWhXWxaKIHSEnog1cw9emWc9FtZPUNp/kurinMOhM7
pmgx5ZAjTHgOQTcArWwS4KhPWJMLZNRMlWOXm6fXHMXcwRqZBkxhVFIIkpO1r84p
xkfqMdebQmA3Tvc5KJNurYTBzfMuIqa3GNeUZcL8xDX8oZf1/fGy0L85EK1LzNjI
glNcboNrmUPbhiD4LARVlXFDWJEKZ6LbjNvuuIZG6Onyq+x37PbBcs7ZC2Ir04Te
1QFZc18YX/zQC4Vi27t+bGN6cNY66MLL9RhW1Yz8vRBNdbIrhhy0FXzqhn4yBUIW
JE1VV9WWEP+rBSf9mpyZvCTxGSJ6vSggTWWG4xnh6eDm+/o2mVLHfrtMJuZbjMsU
7civjK5XblsXqJLMQMcQ/5mQO7/928TovJjKDRZ2YcXc8NjVEr1BuTEvhBlJzClL
tYwCq8xBkjvscjjrPjVuPNTxFAqbkBNTO9acZ21rea1yr8fo65EKy53RzTTPa80A
nOeHtmGEj99ZQeTJK8yYDtku+BNYgc7pqWXRxyGch1S5j3sIcPXmNrycUSfLftrm
1LPJjw+qjWGJ3Sw/bB6RuYBoaTcoTQwPaFxyW/mWxCJE/d6HrO2LZ/i53JjaA6su
yYMHSiuRS85KzlK1N8E2RcaJbPQ224l52LUxP/FdX/es15p6UT0ty22G8mBvNjGZ
Rkxe5hXgnfc3nUhFAobSogMWLamX+jEGY4qhq/LdUA8Ya1RCcxHp0m8nSChpkJ/u
4DwHv6RrnM2DDE0TjVifqHT3wcvLgcopuzmR+RKNsnJcdxDToZEQWI0tCvfj4nhI
HWqjXwrGPqYfaWRTtU9crcNMOqojHM7B7AXLMC4KMy2HjkQ4eDcmdeHnRadLx1fd
Sii3ZlUexyTddHyQV0ETeB98qFH8aDq54WD7YETryQMqDUVr2G/Az/8gXBJhgwAO
2w5dcbUaNuVvgwdMBiGnevwNHfW1TbjSF+9veYkhHBtULOmmvyY3Q5V14OGobCAe
Pj9l5yV6h8R3gT4OYR1kbEHoGH4GMcM/Wur4YjTdFzdcIpMwNh+cwN61CwEF9YJz
Gx/Qs04SkJMedub8a9wuPdvtg2pRPKPfeyY2kOyMerXHXIWrQCFZW+yCV3JnsdD7
lXOs5x1DhQr9IMNQ0C+ISJ06WcstKOXNZG/uzy2ggr0LZAG585FzcCD3y9z7HOuW
lQ9OjDnX5tK64vxjcMAes9GtU4FiCvTyrbRmPaMW2rZz8W7MQdVb1EwbRWpEf1Je
dp7bYniY1zCKe/53L7dmJwtWjT8jrLuF1KTLYDJHNXLcGTap7scsdBcAkc2iTWn+
w+McKuESTsucDTdxYWAVrl5DvIs2b9FTXUf2L7p7YvZen1ZPd8aR3Ix5KzsnuAil
tl+VUMOglfLXmE56v3UrvQIWTLLUXXtdhENCmUICDqvlkmIAtii5FInJdAtZ0LWl
5OA52jL4xtoHLj9Nu+Gh/tgiAPusB0HLocNyPh9kXNTZUbDQrvdFKM3OoxITc+3i
Y/fdU8VQaV9wsiDeJNcasocvkc7x3qCLPKblkjfJ3rXTlx7NskehoCKQPqek4cdc
PqZyQeFV3ZNhlLIiOJcTHarpFCmTSm0E7wMzlez3sEuoKQXIJ/InWg1wWP5pmNe0
7BheOkS683Mu9EV2Hkq+X60eBaDIXoIUVtOsxlXKxks0wtiGoUSSyuZFU5RoWYga
g+QAY+rZTYcU5NySFMFIagm4fGzlj8LzgeccEJ0NvcoWPKMzyxnnEJKyFYGzIr0u
AkYDUqKhDagrJ7n3L5ZshNit/dB4drkujounCxjgSAI4LrsoHCaeg+LQxLdV+hcn
2YdEwOEJCiA+3MbAFaHwSj+gIeWabbXuVHBdhN+CtjD610G+1JcYsvU3S5Ki5Wt1
lm+dm+pgKtiHDEjGK2ttF0OUVAGB8LN4xuRO4GKd4I2+ApdztSXSfqPhNdhdm3zd
Q4S0ehb2Dcd/zPSgbqFqb8mJRTqCB5s39nMZd/PtzeaDIqDJu/2DWOXg71v4+sF/
FV12onNZYVrxo7jGl5JHouOPeETBcZS0vLtrzy5FsulF3dZIszNp16DjnLm3iFel
DqP0MGgyoRijvIzGO5xXdHwB/M71q707cFqKswT3wSBr1icoq0JWOiVr1MuGCg/C
Kes4JMw3rua4OpSmeuJwHurZW7Mmj9oPGcCqXR0Atdlxfh8ov7us46DBe2VM2I3a
jsGxOmBu+Z8aK3nse2+4Y4NTgg0HgjQzfDd7qY4hu2pTWMPao2Ddl63A/Njbyt/X
BMyS1+karXGKa6k0am4kGJXIOhkZxC/K+Qt4ES+QUt6aBWHcZBYeMEiV99WhFhUy
patb7ZHEfzXyKlrhwrFOeRnAPv57EWbqrqhs+eEtsT1lbF98REbiWFeAt006eFc9
V1vH94zkLEtltvNfzwTVir6iL25J5ILlBtklvas/WbSDkqnxnxBKDv98L6EbwFif
YwaJttLQ3kWk33CU5W2zDi4IucBG2U5dqrtt3ZtjERe2TRUUqabFqeqwNhQFiIFl
mvk1DijrBsPxZ0uN+d+8ZTz4n9mc1mvQcvidUIB2NwOUEI84A5u32qBhfCvMgjpS
TKtR7If822VWKFMY2qCQ4PweiEROtqH76Bonxc4/RhcB5ls5Iyt+wrGf9fuHkn0Q
bKFcuoqauCnXkABVI0ZOkmsTiVTWIx9qNrDPSVHuqV82ZzKmnyXDtf0wp6/ty1MO
4n1l5HUb/qjYmjoMsKfcrvmeyC4a6k8NGStVgWBNVp/TKF+ismF70TM7Xn+0B9pk
SrWJGnspDZr0z64smDdYCuGMpV/jIlRek9wQljNcYXaknYxxACuNPUSa2e4HnLAE
RjWwCpOJNeHm1fxCDcGdSbqOxC2UftwhNNdK7VxlMQsvZUJ+CRi1f21lj36TVoZO
nrb1iwjhcL2IFQnCPvAI4f2mZA2ybnikiRyFN0BSwOSlAlMReIPSJ74w+r4XSPow
au8jf6AYl/aQCWYpqEESvk8InbgYq4ceeWQ5+aqnqishwEq1nNSbrHtjmfAK10Eq
c0+k7F380raSzubxZysaWY4nat8Gl1XQ+ahLU4YM/o6E/I2ysoGhrBSATlGrDKb1
sGzaJAebTU7iBgL9KppwwBtwIsIa1im9de70LmHkQ26kuAyudCEWas+d6gtJBIx5
D9X9mGWrGD3F0B7qB3RY7R379w2fcoVT31c07cOzF1yWJk/SuHRVwc0TjKe2YKZg
3TObmWu9CwInLSLIp/XiE4Ap/AjzkIXE0E2OoFb94Jl8MOHX5FPoocWPFVeaVKfk
uVol/BXEnI7KARpCXnebKbct+i6iBgO0vGvib+66trK+jhngzTBwgXsAIPUrj+ds
haTArojizAeDuOm85vWxKuOzwL0RRYlaHXLKdrDVxUfU1x9wXn1bnsZdFvYsb88b
+Vtl1Np7+LIhDTDQrfO6bi0gMvgbT5xNldmwR2gpWfGJronkL45hfpTX67pSqcoX
t7S4bciCXeC67o/i50ijTHCVdThDaaeaKnCpKqdLLdrBgGaQB367ByXkZqWxfq6N
JDlTuWthqh/ntuCfyELZpXyUR7f102wMp6axnAOcGkdRutneyv0VZTAOusZ3KPLT
JkR3dRofbVkprE2Qj2dCI6rkOTqhPfcevuLWrlVerw1D1Wa/h5x8fNj2GQ+v9xYJ
1iZYnbAts/iqf2pxd0xbOlcgljomoORILnCJNs5PNwD0CaCzf2Vl3Rm56KcOFPU3
J2wMvJKB2Xy8Dzmb3UppaJRvNYdzUOk1gQa/MZG5RwWWZMgUXZurh49t+5pQhNe/
COrweSNho4ttzzqhwwgLH3lDSpfjj3XyQwaOBIPBh+TzfBKxDfhLtCWX5ubw07eI
ADfqgiHW9rNI+NWEv/q1wPld8vdesRCQWCTgv9bP5rWZJhSImpL7CYipSq04uvgr
Y2CP7Fz1mI1MUwhtTRDQJT+dnR1FnFrA49ntRfkZTSjI+69K8r5ZY275Y/DNBcGk
r7qcZK9MSNnF9vozi6wHAYFRgeTbTdhgxddxoLoAM6KmvQaFoWUm3oA9boHAYUAz
n9vHRCqZq43lK8CiGYdVxVNhzHWqdMG+8GTBp6vEmFTKw7fIXcOEknNOgCnj/nOB
9S2MmqObfUimHS0QNVSQRtNghg2YL6nkEmQdfSIRMVAeYaIa8bGKvi/kkH7wlDaI
59NweIDCnuvDYODE6nTMQsxP3yeeUgT2jJ8Cj9j7InGhuILzh9slEVVlvJ1in7+s
uZcg4NC/NUPAeHjJCNws7L4q1MxR7TliUocK4lL+cCQnsA7H6OYi36RmWFRCREAP
KrF0X4TB08rr9myYFLPoPcIwV0BwDkBJer2Lxz3284uq758RALxQ4Ly/LDy6wbD3
dXHGtJZ9E/lej/lgAle4yXiOiYJz/bMe7WYrPQLdR3NmHO/I3DObw2PQlkdCPGl0
5IfMcSgIAzhNI1QpeUnMQw8SYKdweBaOkMX8feJJXedCikr9MtJ/79xgeemjONel
Qy1UxB/Ths81L5VWHQhGxVONRPgeRvxcuMA4Cl0FK7g87GGSSon/1tP3Oiusrwdo
4sdNrO1xnFKPt/ACN2WSbBR4mDSeFh5c65lv82bidnLx76ylqBC1F6jEHR0fmteP
vACtKVfkK4oi9xhFVn2zcEplaqoMTUwlmUW0I8BbiYTN3BzEoSWW9EVJjcBcMQzM
3VYENMqR/svNFWoHksdCK7tDu2aSJEhskFcpQDypzM172oCc3l+BFMLlm0R4pUHa
k4dOEt7/4fYgdky181vPlQrb1N82CNQcf69zAEzs7m8YFp+U7ArNdGKnXRV1Lrrj
k2K2YbHbHez86UlKDhhnKixfKmLaJ7JpszJnloHn1kp3srsIju/8YcyrYuI0iHOs
Zw+AlplEJqe+GcrIvCAwIoaDB9NIn98HjI4rsG+4LO5u4roU1o0/8bINnATr5pYS
jk0c5Tqixl0bS5VxVY3Dy3ZjSQr3bWzILsqWUV4sYB4DHfwf+TKICtJAbWUOwjfU
hEA5c/fAXGkXddfO2Ez2IrV0vsfvSB1PM0CVQufr6CtM/NqNLldPE/EnGOdoD4CF
gLt5Hek49oxnEC59D9PbCM44T7gsa9/iTJ0VMXMke0ITKlN09uWym7TMtSETKE9J
Ap88LgaYZTn32RWalvqek5x2y7qZDoxuWivIctgev9oY4uJl4tTXNi6UQe99tgWn
2A4VvEWs/Yib5XX4mnOz06D5XW+FNDn82yn/5h4NXIQluMalgnGX1EuV3x1vbSD0
130UHy8ykXUjZ3OFBgUHXcedq32oWT9YND6tsA3UYiwucn4g+Uba9v7xoYrzAwtH
uYcTqsNjfnUNspHPtSUrNwElWuHRLrtHp1YeEr8wXO2Q26MvU+TAP0pr1GofoR6h
S8f6N/GhNmQ2jA78jZDT/9bSNKNPwex3rv3bLax1FYfa1H70Ymzlk6drMrQUSRG4
TK7eDGUHS+BD86o3H8cpJ9DOo2RiFaRqeGC+76XOH1K+pv5OLIXTf8g+IMaQ8di5
szUaHHW6mWlLDoBcZ7OUL3MnR04+/PY39rwwsXR5rro3NSJS7sWMOaUXrc1w7Ks7
bX2wVYpr9r2Fpwm92H2pGcIW2uoi7BTJEeC4RIRP8MRhv/pvylozoj5XoWk7KyV2
40exDSV9/wo7uwSllzL7ahlR0agr3fOtRY2Z+vNVJl7fZ8VVK+4ReYCW90fdSvhS
AApRME80lQUNLSgJKBTL7lTId5g/tXXIzhKYjjK6houYzJFs7DMTU7xphkqbEjIQ
uhg51gVgJO52heTWAhT25ue67xMYidMJ1ivJFRKTVPXt/b5NpHdC2EItt1bClSDq
bpzzWYXWbG73dFPIaTNPemZz/N9vQnxHXWpEEZTFkUD+ulkQPhEsY2asvuFqBbRB
hU5IXy/w8eNHiI3APEHFuZ3BKVwDRutFNL+ea1pVddGuyKEZTv4CSDz8+J16w0kr
KeO0lj7XkelgVOg6h9UQdDV6smhYDCP+FY6BUW0Hc83270OQ9yt3+yq7OoXZgo0D
cgFLXTBgMRiY5ZHknjtfzINM62/Qjpxc3+HCaBnrQ+InrJDqwSK45QhpEj13liLg
6Cq2AzBGf125ohbM7uBrFraruTuABXLiqCU6p4e0vX/CpRrh/GoT8mpfsgU3RWMv
WKvrNP0ZtHUJkYl7LNq0hKsYNS7j8iim/MbHYVcRFzRk5mCm7ozGxJ8s8OFDo+5+
rOMvS0QnFhzjsPGbRpVDMtvxljAIITtm9g8WHszfmzi2YL3W2qMUqa05OxsH1H3T
XQEQfVrilRnG7V6M6olYicW+ZqEldVRXJZjeSZ7wTaSIIyG/BVglgaXQcBNwT+cQ
9NRa1vx7ia1TWaV7XL2hbWroDdXi/s3/QD+yjyp1d9eQIvuxBtK41964h7OUIaKc
K1rGxgDeMNTzS6FEheWcQwDN2Hce0Yklv99SryYdXbZErIRr7KOGDG9CzqpeaAf1
Dy6mdCEHgPLppyO1NepsRESK7sxvj3UoHkxbyFFMeqhL91N6U3pANRMasnM3pbde
kpIJ3pbE3BBVYT9lj+a/dNZtyvkS7ym5DxhRZXvFbLdmTjEUNxbla4oWFdd/l/oE
mopdjnqWh7QERDpcv7frfbXB+LSQB/X9Mo/wZNgAMUn/YbsXHguC5kUm+Tc60Xe5
liTL/0QLiNyIfciItmhC8Bpu5sMEET199iOxYGhmQU5NQPqPaWMJZS0KmLtp22Iy
NSZbU/pg+sHVRJ3uML/HV6skNIga6iyB0FxY0blPxdeABo7SOOmzQ2TaCehuASR6
/lXRSFUcCdS4WQ8RKzDVQm+pKav+PaSyNh3NKyU4ZZI8ict/KQh+Oh/fsEvtu3EN
ErsX3hSVBH0UDUl/4onymwuTC+gDoQUiblf0PkQBETLwjR7PPDfWxVzOHZComYkm
QpFhc6adFLGDSO8NG4pfLel0v+64uf9w1CRuiK1LUMtGvHJQOYa4awSLT/nmQpdb
5hyKbtLuhDfiLPzTplq8zC5eR7YKAGxymXSAh1SqHdxYCEr5+6mPu6MTUVUHT+lp
RgXppErsS2bV0jC2d4YuiHCTwswQImHyNhfuE48iT2kUugmin3THRbp0PUrUznCZ
u5M6gXAcd1mBD2DnR5IIUIqAG0Ipb/lLFAzwoIadsVwJpcHd//htmsJL7kv6bS21
VShqKFu2jVR8RGg0uVmZHIylu6TASPk+U06dDEM6RxRHGbycmAiP9ozTxLtf6Pw7
Fzb8M8H9RfX7sH8Y4CCGpUvqPe7oah1wFHv8hN17u4Cc1uFlFZHiaD5U+JaI9Z6Z
eO8UegCDMOM4a5bmoEAZ0Ea02YEyxTgfUYwr4SpBkEbZ+JTtyZhOfG6kI2pnWtvU
dYU2KE0Kbj//CefJ/6lF2QjMtXe7CH5+zXzgCp/nUUCUbRtuB317iHXT3ZoLW07N
6v31bZIy6+m+YIYv0Z129RLlGR0b0Qal2TfJX7kzHDenyONgTOBkui3FLMm4Tz9R
EXYjc53cg0HUNS2mfIRik0hdQt8Si6hAKf+UITSTMivhB26Y0Bq3v76E/6DrxejJ
CQRd+f0g3UXviFuRb0P4zkbSc2uLAd8DJe7F1mrhdXsnhcwxSB6ETZ091YVJ6UIx
V1cgCO4zhF+nCLALmBbky4IlK4mZepqMjHTKoesdTLZ8cN1Z7sjVa/J0c0BMQF4C
Yc9K6+T71r9IrqPKBqgA/7WaORur5X9GhQtKfr0hjfpgJ5dfIbQ50bbAtQf43Vf1
NFZ3QMw6DLBGCZO0XdxRFqPz2dPntgL6BklpmgxC+ruhwedCBWWPMJETs9TC2yZc
1R3hLDMMKB2Y5g9mxf1AqBMt5MPD4n8NLDjbtC7Hpp0wCfYTI+gtrWEo57xEQnip
gjbkRXaTfHacrXwYqFYikmpQIAkNxEwWBPDkt4tKd4Zvmlz8NqUimlMdrhtmt3IO
0RqvdK3vogshEpd8E3lfng1gC/+u91RBX9ElsnyAni8LzI+YnZwhDKf9zwDVZSeE
1tHZe3SxLpF7yVwL1sRVNPNdhBbyPFkhoZGMm0VPjeMtMxpwn2tyLECsVy+KQzlj
IisO2SvXxzstrh7EY2qZVUGsXDHVUyMy+GtuEF7Pr8wSO3PQ257AtsPw2oVpe7jD
g72yNyWQTx/zyOQgA7+yoFp30Rs1YIRQUtwpZULzdYrKva7jSxpo6XyoEq/ewBHM
WOFN2bizq9vReKjpky8swrXsvF7LiQffJUSegbS3FkKfFsGECLaPUuVwo8HzszoG
JqgYGmA9M2TV3BouT6GRYl7vr0gIvcre2szGuTWgl1BR49C9gE+y7QQRqkoAgQRJ
m6qXEir0Nxl/YfdZSy7J1LiuSoxjs4k31Exm9LA4nfd3ZqWxR9Mlt4A3jZMYFMF/
khkAMvpwMmumZe6fQNDRx25KVLU4L5rrEDSiayf3Vv18hnAiS32J+Q5TvSdCw4Zz
/T5t1bnxRCSNpcV0X/bT+u0hRq4AS0izSnL54mMQc0i8auRJCZ1gCOT6vJ1D247c
6iJKriazK8pSQD2G7/lLuxpsDW9Us+AUwX09ZA3j8Ie3Cud30y+K4uCb1+Dy/Z1N
03XRJL29k455V+IXsoflrh9F4wo6SQzhfQnZaVLApQfkg25BCi51vUtAi4cVhl26
OReiWDDXJn/1d9Hqh0nKSE1WZNbgnS/mN8W4JRE7sx0ONGgYsIMblmAukDT0pcCu
BiBFL7rKiGTbmfd309t/8Izs/gTtKDQhytE7W6HVCQaMy8+9j5AYBDs22PQtXkf+
tFLdV330EYwYwsV4y1Q8+CWXyjv2LOron9ZasdHM9QSb1lXD9UTlAKciwKou0B5f
wG4d1Z01rlExaBivTy1nCy1v1DbY9nj+9CkOqu8eTUUzXxBDAtqoZylHgDfN6v3l
A1D2+5QGgyUcmgZJGFps+dcSgrCHL96Q4fs+vwjWLBhiqkovhu+omKkhsh69/cNX
P9/s+WStjY6fTtUOCDLfkNMzOz4UsTLBe+u99ONdsoYIqlWa0m7aSb8Fkjo4zj1D
ye+oo+vbieVxT+S0wV56TH7y/IK+mHwqN26gMM3DxBGFSoisGtOVONy4DCC8udYP
EDKvmhVisQYvz72iiaTH1pGBHVE4yP9ALbUam8ZBMaixtX4tkcC+lnAgwn72R5DT
9eK8DXt0zwP0irt5+8RQ6zbB5jq4UGb0WrA+ZJux9IM4eB5qBJLUTwfZkZSYN80X
B2DLx/GMYE0B5AWr83eAyMAnBy7XP7MdHftHNJ4VogAliTtWnoYEgo+TuGFnkVp8
xaKmxp0j8oWmGJ9wLCEeZcHSSjhoOIqdOfGN80FvN9kMbi+5Yb+bBAlK7qbxnMUc
LLlb/M2z5kRdcwQHCpjhpGJ5CCjR2jSwsFh3q3UIuv5Eex0HyhqXitBc90MvoTeD
qkq75cW5/UK4rxJSdj8RtzS0aspI2EzrDTJXrBe2eEGMNLFwS//jZywzN2x80zQ3
jubIt2IBNWVMdXcdtCm0ubUn2g0pgQ11VPpGGsiucjUpCOXK9BAUdQJ4EHNzh+hE
kipAvd5NRYC6xYTkoNuZdgbrRzNNCwrZRA0CrnUCyPJHjX7bteas4VkHYTHSM0J5
giM9VUngua4pGlEIKRVUD5CZKClAgXeGqHopmHjkf2Ad80iA/ZLFYicdxmN3BmSX
2PD5LpJmwYA56F6eDWfag74C1WOnffwrn94efVWf7pLvQjCrMz/yuYGaur+90Dil
LCUOlZFkZUqCjksqFSVhVditvZNP47Uocz1hp74UrqUEYhyP5tdmh+Q66V7s1Oae
Ic89c9aREGKxSsB2bzNqlTexNfEU47SX6RhKodvw55c0XN6ZNXKAe1S2UhoqP7On
nNi7DKFSE3X1DmUngQbQGsZN2BzhJnKJY/UE/eZyPXZqh2n5d1R8C7XUiIUZngof
yJPm1/wIYDaJrSaQLivXzDUHBc291QlW3FZm5KASarVN/ENrZDMLzJ8TCmzxyKqh
w9bChUG2PQfDFWPQIDxTQP00vs0RKoxLnzKjf8SlRp1t+fiS2nty8SayUcJAE58J
eSvy88tdbVz9gyByB83yCx6Lltf0GU2S6lXnwxxq7D3kmlcuYasPYCwT83SiVL3H
s+wZK9DhM54yWe7Qg1U3diRHs+AetgCew6VbCVrQjylwY86KWP6+WFse7G0qYuhe
j18Ho6glFJKKA1v1Xwv2TEXg+A25awPSXiCq01JrgpgZct9xN4Py7E0nw3xSRlg+
dEVwbaCCnQe5Tn/6uc6n4JzIKdBqfZai6hkxk41bAUjR6/j9X8teZrOZT4O8tIgg
7AqVG+WEyjJFVK/DmMsTcifvnxVPqPopLjOL+reqcBG2kbMnebGJkb54iyhw0KPy
ftdZoKXBdR0vR+5aoMc++E041wep+L/ng9Vz32UoesQ5upr5qfGDkxSfKLgRr784
wa2/wpikWT7N5EuV0gBRp6+6iYvGwccqqcAr80drTr0MOsF1jvb4KjO2hSA0Rxx3
DoTYnsRvZBtu5oWWjABw6jkTcuEH+4XMn6Qt9KVSBZOvKZ8lM935RSsPSCPssBO0
00prhjWzQe8PteXYjH4NucMuCicfs6Qj5KwFopzPny4cJPOdkhrayrwwiuVRJk/n
N7TR+FFJKjl1Xfcp5vNC9+8KaWyCk9RllVyrgyA7Pj/5k6tcOegi4Yg5ia23vlk4
38SyiZ3TXkLclsmPSXPQE1USUZQJ1EK0GXjBML1Xpx5Yr9OoWVbsKitt3G2rwmTW
JWezI9TeVAOU+1ThqUE2gikJVsGKv8WkJkZVl/X9VXxSgkozTM2mWQ4PQb2kicJ5
sV81PYk1o53irFVfhymRjizGojStpMk9hWxmAFyTztsadsarQrWhPmHnYzatuEHR
b19vuQ2JO8wVDQrx06JBgD5yvU1EXaO1MsFmwyHHA2db7LcSpQF1KDW7gpQ225Oa
Z+TXrwwy1kmnPs5sYuZOTCFiD74qC2qJ9+kg2zC+7Q8TaTZScW/2S/RdGGlvOt1o
fCMpiIcq3skTHJnwaYwWhnFkWtiDR6YZ/uZvYszSRLDSh6wZmLbl1YAHlvvVfIgb
dtwGlebShcwz+ZedEGosIz4gM7X1NgN2z69Kyfhqxoo835CdhIhnFswges9NRr49
1s+W8TcNNr2jfuyz+8JLaoodoHedfrTNpw1kxFX3lrEFmXkvlYA3hL+O4q4+M6x/
jmqiQFWstxs7foawKOkAnSh4t/4vAYc1V+wO7JY4MixQ3sCWEjSoSRj+J4cjRcgH
W39Fi/q4HeWvvoZErIAe1Q7dpgOcQ0mQ73/PjvkINrmmKv5DI1NyA+YGqvAqRPpa
aA/IqjwB6A+M7YPpggC8BK0czVeK9dtjeJ726BswNOtVtWkfAIoO0w4bB9n1Wo37
cCqwKkGmahxaTaZw0/pWO12dzhwCBLEsZ0Lbqx63UIAEOuV+ww7vlD1JDwQWDc6I
+FA3LevMxqkANtTd+zvxKn4GM2OLuMy/bISQHIDjBPT6ecxbGsy6lNHCRuONa+mO
vb2PoocVrMbAmPFMJEze2hZULeAg9NGZJLHRDlLgFemuTynmSKAubssb3ILFEPAQ
iy03fQ8nsJoMgNLxjXCNf0SlkDlg19knNL7mZoyawXxKiUyQpKfkiqEI+i3yFIE3
A7pmXBpUqVvmv4Wg+ur8p1M8cq+14jhbNdN2E5ljZXnjI5vRInH+iYFNfsBxff6b
AlQjVH5+cGm+tv+nOCZ8j9jT2rYNKb/d2HRvrE49puxp59/H2KbIVd/5kRPLl2ob
Gfgn5UwTV+wuumsZhg7Rhtg6qtfinqEisfALjD38cyCWFxn8VG+1b3Sb6dXu4MnP
WnuCuEUv1Dbkn0CvAaO3qCCb3k/LXnQqUYeet3oXu2u6sLKYIiQ+OIwH5JbUCH/0
WoCmhp2jqKkWum3SmpW7zIK6Whc5j9luQM9C91Fr6U0hxYbZAfDCD0Hpya51FJGu
0NrT+/TK1Z1uH1PtP4rgE1ZPSXb/ogeFSIr/fElFu/IO/tCWDGFOWZYs5qXFqEfb
O4S4jrBPPoCYvvhyI85VMWb6Xe0+yCaP5uwjtFBSljq7OPXFkV1n8FOpIazwVMlA
pBhcQfh/A1WeuvR6Hapeh6MCK97ZlK2pjFyB3l6oAwAzFIZ+AAgK7AelBodqH/yp
iJD7YhfXM8Leangq8ItmkWJ8/xRI8AFO0jENhT9T3qEqulLY3GHq/7yKBDZV2c1a
UcmZj/gnlBX6M6kGZ+FUwBmQvK9t0nrZgFx1aQoi7yaQj2FqXOc5UOau33GUB2Mc
tRRo2Akxb8HZBCxW9qTl3bx+Xblm2Nj/sy3jHTUDt52qJyFlUfCHhVh/LktWEXiZ
FII/xKy0bG+0/2dn/alVb9vQKxg18Dy3gg4htB2E620AnSI9Z/L3wNVia0QeIjyH
zIDi2wdlzqC5q1YmEfu+STQQkhpUzWBw6f2xYzu1GeebYPH911m7OgGaAdsJuzfT
+uxUB6DT254wmepn0XWZVKhhyQCDq7Z0fZas5bbOjKsCpCdxuRmRBmjYRULSoVZc
sZ9xRqRWrBPWl2zoGjuN61ZXGFPnysbqkwzz/H8vwID6RaoDYlNVtSoJw+ty7FEg
+iwoxoMDycYAYHHqGEVKgwOqhhXZNp+Kn2KCvM1pP3abcmHAKqxIeBFGbkEaMFiu
HbcskFtIdn2WFql4rzaAQ+KOpmnq6QlnQVwEFV1jKNI5RTz6kK0vCNe4SrAdlavy
pGE3LgBUn4qhe5eDT5SL4KrB3SYKFycxmfGZwmokCZm2HslSBTa1fJFYOb6oUGnZ
hguYxtRiDJ6CnIUYE31Mqn4NS0pwfdqjVOgKh9LB5nWyUuo/7xRLU0Qqmnx2Y90v
0XuNyUjCMntZ7HXhUIb4xXU+mXeZUKXzvwtIeVyllndXJipifo/jeWx8MVFqeGk5
o+AHoTIuoaNMzjQXdML+YfoKgDITlokanq25XwEM3DiarMOlvVAtgPCseIVMh5iH
5Y6YvtFyhVIOY6NaZcvqTIyVDKGO5ynfS2eiG2EFMswLPpUhZ0ZiWGNauLevEzt9
d2f7hVsK4NhMKahb9a8vqMQxl4b1070tcqV20vLbRk6zSMTtYpUn34fAd225MK4P
oiiuIN1XcoE8qsL4pFty8ChMlf7hM2uqbTXtPqmg+pcdUZnxfunCpr6J0g6uHJl/
IYZ0rigX+9Fc++Js0KbXJmOcZ93m9pKSkQQr19EkHGB40VpSIAMe0dBbb8qUwuKD
mfEMeGLnu7VzTEMZV2qxNoP/vBZfiA6h1IiImrVVtrLSMrklblQi4upP/TFLP/F0
/JJdhehZHF9/Nx+wntp8OYEkTuPpZ/789nmW/S5/KrxK2alIvuT6bFoalJFlZUZk
gCejHSqJkrLnrBjQZOZcUYrlnqsLOSuwhGlqx1mqq+l7jFJf5+zBNdFKWUgm7A34
QYJnppRKItgF3m5Sr24XQcmw1h0W1AUU1z11Pl2qBql+KjOjaXZthiclBYmVYbwM
sNbZEhNVBujLfz85k97fkvllyDAoS69ayTW3yG3W10TBuByIQqD9zBK1cxAXmXkQ
UCOy5aR2NwDZTgVK5ph/uX7Hiqi96sMpBKcF15VtnkyI0ldSLbFXpntjUiI8gqw+
gle32jC/fF1F0oVofJkUcLC6mbY12jHQvp1nak9rN5fT0tRE9WG8XjAeBj4FYEu0
jwHCNYWbPKRV/92/Gzv6WJM9Gm/meirM2jE7aunBcXQzWcZk0u7ch8L6ZajDEmsI
6PYuUWHKD+dFRj1fImrnU8Y3T0v3WRBsQ1c84nteTdyQdpE6mC2a80QnhuHTinEV
xu4XvVYXbXU8vtbq0X/t53vxJL5UOa2WwQVTpRhdlmGytLmV4XOqV4YJqPxFBBxm
fANlx+VJF2ZkOwI8nLfFlo1pGoZZaRCFEgPOm9jsFHMfgc6RAX80cgtELerBR7qb
gVNYLLShHpr2aDPKxth1zCVwqadvqfKSQ1LOE7KO9gG895O/v1blfMLiUYL+eaVs
fM6mcG6Hukk7MRZGZXbBi/sK6KYnf+C5kClEdfB6uagGrpNCx1oAg07qbvDAX1TO
g2CjEqy9xOXosFHkSgqgjjM3m9coC5umKiQOxe2w2Eh2ssFKRzCIh8hniemPAxp4
AcKIJx7M9vQ4dT9fhluRgyTBpM7aLCMmnRvM1ZS/qDZxdZy8OPN1/0TelAE3zIV0
UiWvYc7rTvAHVxH8rQUd3dZL2dvBPSavHO6v5J3PuomGW8rXtlvC0wgEfUcTymOn
WHskok7HlJE0aPur2e6deCgNnOGIElZhvLtmI1edIWpcLH0C/TAVOwTIJ+d2LBtc
9Q0lAZgLzO87fhOywwlmHZTchqg+Ema5tKe/bv/PE9eOerMH4fABaeryGMEABVs5
JCkI/nckhTCsOxn6UsTNcMcncBZH/J5vt5K8tHXMcBgfvAaHqyUMpwqprq3p3Hh2
/WH8uAWG8QhJXsoIcZJOgaHJPhnH3wxqQ3ASLrsXyKujSpZi2ySQf00oHOpQNOYu
Nm5uPsPLZszU1h5GSb2LRsJ1doCv0YoHzX/heAK4211jlCceWx5wqU5fY4E2FrZn
2NDOhpGOUX3G+w+sF3djcyA/wcA/felLC5lYiArKSUYX9uEwCiV4fDyKVaP6lmT8
98SjGh1E2HEy/1c2nEbUWnxqLd17Qp5k4SqejAQpnZfbjf0Xfi7lEhqhfsj+8vGb
sVI6dS8WBerpZQdM9kHpA04dJTerzXU5Aw4qydewUAZ6e1THghJcQEvvOspxqon4
3+fq5zYhbt5upolhc6LO7YkR+VxhNk3I6qpagbat2t7MvTQiNtJYzcmiXaRFhquW
fveLXuSKiMnXUQFx6KSyafjKu3V0tZhqYGxbEDF4KBxyWYwH+9CiGZPnHYNl1cZV
5sDX+OthnbDO0GLP1NCB9KFWAqzYtssMsQEtCHFh4b4z7RkvDpxFoD7uSsTCLWwz
zd2NYDs9lTL19yAZ4WhILqGdHRsJ1g1xsIxlOCcUTnHGXx9li+vDbFGzr2l2kseX
M+2q0di+RHbwQ5qNPGTY61UsNppsWb41vILWRyqfWqLUwQ3QT9+j1PUAgZ1rP6A7
7CuqDYolMQ1s/va6KT8EQy3qNrGwg5WduwD7uBT+9RGW1IHhqjiERMiH4rnnmt77
8ZImNhLfH9zjmMu5uF4PUhPKUqUd7CshoNIx5rrQYZsqFxoUJ+dCGxz9Z97IH6jf
SBhEEfMEIankiU/VXiFz4gzTvq3CcNTuT2d743tTGzTWFXpHXC6usNAnqPb40y4+
lxCxRN3JZw8o4jkGsb+L77AaHnAr+TB+6IHJ8j9q6wtQYe72TSy9vQ6YoN8vvrBn
plqwKXDAWd8LaFmXhAWEZAsC2ioyoCeuBLUQlVcspEffoyTdL+WTi1fHIv0HKJWS
BlXcw3uYOkDUfGM9teEGIPR/1FHG/y4SnqXnsrqq3tw079fWj6r2NnHXBJuSL1gJ
Iq5AM9Fb6JLEIAyUtLSmu0+9/1EnHcuBLie6b/TQmlTfHfhvrhb6oup9OaDSoz+e
ZW76+X7QDi3xkxzOFFVAW2S7PHa5tDSI/zRjwkLFKHyORRRnbCJsJK3Xs5Ceu/ms
nf4i1x+qPGS9PKG91F3Q3xJbynxRvx4ZML86LcLJst061agequBgFJLi6M90N7iy
/xuWXS57cWuArz3tIop4tMbKLC3QGn+P+KYQB1rfzvMJvz4Gb+a+hd7W7ANpBJXv
ZSpEP+802sjQYXnmqy9YQMtDWwWRrItaCkmvNiqfGJ8a8HIDfHS+Jg2YClGwg/aG
c4vmlN/2k6yAs14Beb/vzChWVazgzA9RKFDwyfQlEyQ4qr2VXJMr4cglxll34UF/
DmRumjiSSsGJLjqiTHdDdPiVmOnN9giY/JmLPM+DtLOrfesMzzlmGsmaytFUL5Xt
3tNSidSdCjtMA94fQ0B2Pog1xW5tAuFON3Pj2mSSZ5R5pc5965DVej4rYDsGI1kI
ldDxNeRDk7u+OaYVN9Q7/jx1VTCyyI1n324waGN2wekhDMGtnNiAHgRY6tR0uFCm
NJiu7wY+aoN9Ce5mAk2ydrND8oaHCKr/KXyCuKwiXezaLX6KpaGfSqT+stU2ziaw
VUXQB/8ebMD4ZL/+ypaOr60Q7ceGftIjgHkxkDdJOk849igsJ48jJFzd+Nl3jhGX
PmlTisGXc6qryMxkXipM8Q2Sf41NmwvLxETrvbfaKocvtrI9Bf9bfUEU6/BE43U8
zYQMzyrnrsPSLiadnpDP3CpAN8CtE8af5otQfUF9HLE31Qq0ymnNHpKOn7fHRM0g
sElwI/IwUkY0zA8iczK3NJx45Ie8Mma303/PPrdy0/4jI7XVMW1/83KwNA17KZsi
vY4KpEFVqEVap5SeA5WQLpwAob1YWesjDTyet5pVtlpkr/T5hxToPcQUSMYL4fTx
Ff4c4tiE+a0db2/Xi3cebXpfQULiUUhy2Cx/90jdABwHxwMjRLc/pPrJKzomRR7o
UVk5z9HKvNRpKFl24LFENYnrxIkUjykJ945J6XSF0D7FmTs+qt4Qt8qSyi9oqD6E
u3zBxyA7xUHGI7jpAFl0OP7gAWcdNuM4z9Mvi6TT17iSZhwCW1OflAvssdX2/xHN
SUBEAxQv74DDsgePMFb/JWr1v8Xz7eIbc3fxLRQrirf0ZZP6h/7Y0QP3hwVK1u+X
vay4OxoxTWixwYmnV8QBBWGBlYJmzNx9JBDwtVyIE7LQd1DSh4GHnIGXM9ouHY0S
GrVVXfo8GV6ZowXHke+4QCszLUYbhx7eMYVY0pfVvwbbBOqgKmVNbZfbZzWFeoIw
YL1MkWYwjG7X/kw23nal3ejD1213SWv/tBoToXdITyM1p2SHTPprEzYmgWEud0Pj
rT2t7g9T74o/3GF50K+aK68f4PXNBue30jcMW7hwAfZ47K1muAvXoDU/PIMJODRa
k0I0y7BRS+UMWMVSKAFP++kkblUjGgWdPy6yPHE+AboLLoWeZOtQfGVqPRPzWuYp
Yc8psIleA0Zl9nGMftNFhESHh+MuU/FbpFFGuzes5kTYPompzh0bbcS9aTy2mD2B
7TwP5jApQa9029LGeEar5f/rKcF4c7GDb00XVVlHQljCPZofK8MV2m4sCWJN7FF8
Tbay92notyx7cmjx6g6NZtBWOKyPUkocDYChSzmWN4RN41t+Rci5TxeKCk3oFXcz
vbYTwlu9tW33dbj5JZ8daRxbsiQNojjZJinSwoH9pRVWShGvdVSVtElniTQVeECI
wlRGRZkl4xFBoVRp1Yqa2nwsyvLQvEDRY3jLkjdix6622naHAWh5LyACyJEkIKzk
iLkycBtuSprlYP2/zdQDsreDGjrKrCyAF0dACo5eD0o7Cs90QV4948zuEjp+j6lY
HtYoTmltluun5B4az7Y8gok19BNrkx6xVHG3aucVbju8XvpFZoTaUdzWU+IwPtm2
nRKbxDR0j3aeamp8HwXzhETvlvWDUBzgYiyZ6W+B1SfjDRB1dsyiVyo/4PpZqeZt
Em+lA4znkhw5HdleY7EO+ZtW5SZ2B5gJqpG7tN3v/U6p6OrKuSbIwykJ3rR1yOhT
KhsQC1+3jDvYLuvRAeutsiKx8YQe8+Q/xUobkMNKqDzdtGjiy3r2//nWkDLEZKhJ
KDaIjIZ9Ijx/HZVClNKBcPjqzXuWtvPC1i3q+fyM2hLs48yKoxwneZvgeBekGyHR
dPBS82TemkE1yeXHzFPAMx8f5QRkyKtn3+KpQERaYaCdW5DQtBhwDCegqd4kIKhx
T+4Jeog1fsjDWZoJ+LUeqE79r2fpjcVYUHHNIYD+ywc4DoCBrqGwwXnaLtxYLXMf
TTpsEsPihGCp9rr2VOu3I4fbKp/4dlClAGjnjaDAWtELDzGyScgHiWKT2c3yzJi4
OzkAjiWw9TRDIrqxZhpPITMCo54CPh+/nmQvIqeBe/0n770wgOpnQR57xCoKjBA7
mRLuONK1+FkKZXsD1pjQ5TqrjXRsVvm9TFW1mjbLKkiz4amAHX7jdKH33ekml4f2
yqJ4e3Z+vWdD2pxRAgD3Mdoer3XAmSdGNHS6KraqpfhgSMbYcHDDOb5LN/ymsvSS
+R34uCDj9x6vhk9vi2d3jzVO8sCh70stXe/4k7KtdbpnLVhzzeQLqRD0L8QyEMVE
9EH3Rsi/kSIVgGUxxXPdKXAdS+ZHIE/9dZ3O9yxi2brAmT2HGvHp3nmTFbM4xKRV
TEREAGlYzGlwTXfBLq4VZM4CCgARIEYmM6NNvpbloeGlDN+ebpYhrgOrSsysWRw5
9v6ciAObdlSOqH5XTRqykj0Wo9ayqKwYu3/KtHtV1OeOQ62vgQIiTI9ng0CKGhYM
B+jmhADi3Ch7pte3hT7W8OdV1RWDwAGTYptF3SG3DZlnIo3Su3ME8c6J715FVqJQ
S5NFN1jQ17rQDgqk4zmsiqlk7mVC627M/2AhHyAVmE9WJQe0MsknprrxPqH4R6m9
1lC71Nhp3jkEoT+gbsfcfuTZbx+QahFNFUs6iGPY/Hai3zj/lYJASYAx4Ue2K+7G
PiuWPNEW3XQZS5NsyW4tZZX358DKjpIHFbtmF82oBt+nMKHS3A4n98Dvhv/HcUe4
weuRLEfKisISQcttTGMzwDrsndlqNCpa1SVpCnssXDn6k6k5yF/uv6zIIMZcjfmS
h5qEV7J1hiIfN3fao86BpSlaqsb8/nMMIsxoBhSkIEJUwYqelSnfNyybpt1BxoN4
CwqIPJ7n9/lFrzehaBeQmmzkWlXft5di3Tyl5CcbNSrLulwmGdGuStjzljn8s5j3
PfE46JeqW76rNe6LPmBVhDOp2IGhZakBlYxonLDnf9jJjE0RAi7AcFKUZgZS1XHb
kOizWc9fnslQ49OO8QWM83AUIb+Rb4mgUeaWxCs/6QQxuuaC0rGn0bb1QexL0iLj
HoU4suPRWjJljxWC5XlY6Qqu2moOE0SKPRsck+PK2gfcmXA/TWnKgQHfFW15q6HV
QHNZ+CJjE6js8Cxm1RbSL9jnVXI1WiRNvQpWh94Yd4JlRACGMRZYA7nY8+PVeJGQ
WGFYoId70yLlY5S+EcS+iMRlZ1Hz/k2FA7rvu1QJ6oSkoa9YBuSqA0LPwnX7TWja
hUx1fEc4IMjEdTra4sfK1PRrhMxmKaompmV3+OH0DxH10+HwoZ7SRtCYNHjbH+q+
oRLTmOxATttKEAHeZ5EHGUCsAX2DQxKiCJsDyLep3Dpcms0zTMPIFg7Lgh9stkA4
vZ2OzuemjO5YIscGVIF7m+TXHeAKfcdqKjBdFg1yBZ1dkvce0+N3tM5aGXUX6oku
Cm5zGOkLhSiNVrwjxdq7GDhaY5gud4E413U63tluC6VoS/J58vMcggp8rXYiygNO
5uIUnwl0K70hRgXszYVkbMag0B7tHtbbxSGMZ9Iob5u+TgwGV+my2puoCOel7S1R
k5TX9SS91lKLCl0rQy/s29xlpBTg70ls3EQwCF3Mb94YdDoDO0a3xyN8ofd97Lv3
o0tCsjizMrpccMf24AUjClQPtaY2X7Ze7JnzAjNj7/VsYo8yS0Hj9ovTG3x/hiPb
7SB1Kk8vTAkX8fKvfBwjQjaRGxNSH0lscF/e8tPoMpGJUWVihtPjR/75n+/Y1UT/
Vu3Sx4mYUVjZRGKGqxGv5x1ztxaSH4V6LBVQOL+V9D93h7wsK7tgtCrAXEOkG6ca
A3pOoUr2ZpXSxGH0Ypm4U+r/19VCjSprfqcAVC0sZd2sofuU83PGmHa916+dqR+0
wGq9LscemaYnCdIAuf7vpXN9d0Z+q+f4d6SDqsty5h0F5sixANIRojszWYiMrBxQ
BBW6x3+psP9ZChuEkpMsIop19Z4JlONSIQydw2+xjUs+OVsODHK05Q2U/aq6vs/O
3n9NiVpuVhAZqrNhIygoxpS6h24zVokmK/FJCM0CIa+7e8uaQozlt/ANAglRLfC4
1kdFaS78dWBgt6KGRZLEt6g6VWbJJFvhox2U7M7aX6gimLrs0YnyXCNbnY6S/qkf
7r3Loct4tLBFczVMunL/z2Y5mPkZx8r+23jbt+vPPp8MUDUYhpbkKk1YXQVHYoMm
XC/dBGzWJmvJs1KlD4zPp11J6DJSd+zQ/4FRi7BBPvIUSThioOwQ+hShFERg7fFk
J9wcTQ7JqCV2KqqMiatIKSoNMXCX3JTYh6gWbi5lJ3Nkgv+/yOYDBNpudbaiJOU5
J8rKCaM1k4BCCWHQjgYHQfmzCVrIYC7a2c51uacDCB026Jpbiq1u/8if9MTs/srI
MYche2WQ+fo5hTzN4Y6rEVcGYnXyTJ72Hh5B145a0cStGGxPB0u7SaKke2kp7DCF
GV0hnkp+gQ4hDgzA1Xzf67JMvVXBCZqensF2UopME3iz632vGKP7wC+d9SsP490F
zCk5vzjV0QBHM3o3cTmZdSwNKpk0mMWDxiKsvgbFRC50O6SJhS9wVB+30xAlV588
VY9vRHOjl1UuTLFe+bWkZwdh1wMa9Tm1HXbXQ88AMn3ZcU3yieAFvMqT4SFH3noz
gtsj9AzywBJvawqeBNwzl5EbbzK4xFDmBCrtoWLQQvVMfshF4ajIvMzyWtTZDVjt
G9POed8uUJfiZuNvOr4XtrmuAQqX5f4d6JSLjtrFHXf23jZJWU6009uWbSB6OJHY
HCbSrJVrzCzU9JQEa+8FWVK8qpB4/n/APAnVm2CLFyrPFxjGbnCnNZoTPq26jLg/
b3enrh7NnRAceG9BWPcdUaYIO2z3224u85NbSIPMPVZzuxwS903gU+0tptk0vQ89
/l70V0AFtrTEqVRI1xHTY6oZ0xJlGnQPTVYzJkloS7aL5zGJKvNwiJRdkDntQ1yc
ARAl6EIjBXxLHGLHGWL0A05cZUKAoAOm6smZAr0pv9o8LlPhMxkp131yEdy57iq8
WlB+m/eOow1C/20WGuhp8VNTtx+VRkwLs8t8SXrBzBPEbM2zYykhw+6OvATkdejV
KNfSlnRsAAwzXqXvmjODsy3Tqr9giVe/PBSBLZ1X/6Qcd5PuVa2mZE4iJ3JjstHd
+DfLhtNdtbDNSSIG7ia6PobSGKYZG/L9+Trr9jovtT2dEijesyVsN5lOoxgQzanI
qLy22Vy+H7lylMXuqQjQ/m2ErL5NJWhS6psH8PNMiCg4E/eENXL8oHfq5N4AlwyG
dkiyBd8PhVsYQgcF2lxssme/b08JBmjMz2YjfrNJIGOTJnt7QvOpsMTcqLVzf9ve
/lR5bvCMWPOAPf8KVlJLpiQPONOrvFVXv3j9mbnYglKSDZrmLUuYhEthdJPCfPmx
HgkJYcyGYGP31HQpwBBkWjljQ+Pz8e6MpJmj5UUA4B6K76zAdOgTPH29NlT3NPxs
TPa4QwqitvTWU3udPk3LaRhECL5Eff5c+aFfVtFwA51RcKX070UNyCEEpYx1nYTQ
usqolPnCjJuE31T7zCXl00ECmiYFwZZaTSCULik24WIlN8g87qYSuYbuagXodLRw
yo5y9OjfW/0rfIL7H0t0NP/bfyMpzx0/jfdBWqLivG5fKvvUHRQ8n/0ktAclEBGJ
NhPwvKYT+4kdRjT5A8RWHk8nIBLDPiaZok4ko0bo+MgPVMiuoq26iqDtkYGPig60
90rPmn38nn6on4y5FdInDG8WKkpQsjsQfHrS62qFRgOr/pVcE6CadmgwnkKwBx04
X+FO3eq6Pj2ERGHLt/16e46yp7gCi1rIa1NlEk5jN4ef4j7wZGV1NwXJpGJMFU4W
IZ2FXAqtTzRz4z7qb+aCMgP8A1w1L8/uxh3gAqrMgHHReV+PIsXnSQs65pH8QszR
hw5T7867Gp0hXO9trpk/KMQFBUkUcMKzWtfFkNHxB/1SPPR24N/NKZW7ix8h2YoJ
1iDXwW/yW1R5IYCY5Ifo1XxGIvCbzP05b9my0LFbGZwYozYEvAhNBDvijylRbne8
34NfP8DtpZn8CFymWzSLVB/bvZ9KV/SJDf88qej+ddw7dOJZ4ujNIH9F2wptL4Gc
+p0bXbHqWaPA5PS6DsigltO9QdsmN7HuhH0IXVp94m/9zTsZbjBSyw/GZlzqXHYm
9Fn6mnNyb9NnnXI3tSW8KHAz6Cm4+3nz4Vye4zUGTlBklhsAy4t8KwwkEmCoEGJa
voCqkdwZmhHwPtE+DkcEWbdHsH52mOl62ptwf2PpfMSedjARdMLLkgVaMjB9G4nV
DF/Y61XFUlv2wo+Eh/HC/WgMSthNQJniuLzQ6aZ1SeX4OFv86xsBJsIfvzVfiW4r
a3GvgGwS0EoRjFPcLdwJ30xjgr7Md8ZWaqv0nBCJOxUIZhoBAWifXgOD6takWhn6
BGC+2LUT1QJplVZJZPi0SElwJFKHzZqQ1SDy+EJUqprI8yLW4WvKFhuN/Q0Z7Tcy
q3uHE/o77BJkN/Wz5FS4K42+4bSJspfxAx1D011hs1T2mIeY6rI4KtcFL9sCZ4N5
ubZn+YqNaqCaZvYDrV1ZNhy0tXKSCq70bIiUlNF4kifYpykfONpbdqmspxAkcH1K
qu8+X+nXvex0D+2bIrrWVn4NgT50N4Js4XQ2IWDhL/0wp959jm+IZEOeKsabnqE0
Ao/WDWn2Mwb2VMy1btN6EecyM1N+nBB5Ycbc8VSQxcEr6mqZRsf/ti3+U5n0VEvX
l7yHNNRrGQz7Y/mrRXGibnLx8LNCUVWdU4rMjk/2aWJi3+4aBszNL3esLW88MZER
xEIEuya+sGSMBfSSzC6r4rmKj+93sgLjlM63MBbYJFotFNmGjuP7v37HhIavIz0R
vSCOoR2GqJQi15hLImqVf44kDV7Xn/BzYoi4EHVZq2Cz/46AoGXr4BnxKvqdAjhk
Z3RDn5H9xDyoW8x/luMTesHkIUFPQo/z6jqMbhlSh4VrlsjOtaz4MC3AMxQ9VBoC
uy3XmZT5j/Xyq5LuLOrJvAUopXV4hLgnYmOJQi/0h3xTXNsvD/Wb2gevvs5M24MQ
ZhLxHynoK1rrJ2tCSq6DFfKHHAvlmarA4wCvXoujnGeiyjRPks0qCoQ1MTOoj5GI
FsE/RBaCXvb3aUMaiqCCU/qcLzyHyLgJ0ZDopjxtJ7TRtSC0eORnB9jaDqjSp9gt
X/iP/eC33054pl1u2RxypLEraAx7HT9vSH4z3d4BRgACGzCIW5A0mKSL64FLsmyL
12qiLFREbF4S/jpv4pSPbtUrQE2G8AeQiIGsSwtb/CsZzCo4QqDcbESGIKXc1/cC
eaZ5SXf3XjT9qCnQ91wxRP+hjJP11n5g5tPvCggn0sBxZpTgAjo6hv5QUZj/jXNu
c2z/cKVGCERy9sEKdyIlppGF2wnI9IiGVNNo7Xko+S5diN/Q//eQU+6ykOItnYS2
hF9CpsCL03oFsrKAik0iWrVAQdQfW2WobP6luOtcee4MoW5EWLDDbeZuM+ZGaFBZ
8TO6JQ2ZVts/4d7E484Nx1XVMrbAZfdUCrJJ933IgE+ahIB9LcK+fr/fn09OoA46
6agb3xDDzbvrPpTo2lIrdupQcj/ik79dmsbamPo27Y9Bj3ulu7mKwgYgveMLAxZm
q2srB4OB6nYBwUy/UroLt4cks3j2ZrFHzaIzewsGWSVm9XKJvQQgFsozHccYhQLj
i3SA3GoClLG43GwMgHpb1AVcVeSa0wwG5I0O3yJSdDRPIN8E+9ERy64mIofMEZBg
kkwMwt68Sdz2MN6RaIq/emIshQjUEq62vgD/wXx4O609IZFpj2wFm/YAZqiJtuWK
4w1P7Od/k89B7p79fxVXCtaDssKoxph49Udpd6RHAe7eNu3lIg71N2BqBAcEH82T
aFwLyhehXMHARKFIWOWNweqs+9q1IaQbOZi3Tu/3agm4hmT6f6YrSiyjknlTA4EF
0yMAyMTspCAgZagynve8YqNYda+QeosAYcys9d7N9Ohlxsg+JXdKxawbL4A0ofMC
ewp2WXXksVSc7/DCRi4PjRqO3OEZNwichG+3jhYclQ6b0kX+VS9YAYjpYqGxKevn
qgFBZHwJotWlj2txwUHLGUQJtBANEOZXIfFPbPw4VnjlvB0Oc09XpXCJCcCL70F0
8+J3NhYREOm19aOvFtzWraaBRmaNAv/eCNBrK+O6DF36zrxgkeBuOvjNH1/N8tgz
dAgL2T4frX0yHO/l/AVYWguDBJ+1ONXAyikzs7XCTE+26GtsvPANUmXD6jWVOC11
40GFSMumTCrmfsD+1b7a6phxLhjtoqPFiSkEuIqiEHWeSVAXhe/q96dfRhs3V0UW
J4lgvRqTSEC82XOxJcRJL6BjDJk3qSCyAP3ssSDffkxKMk76i4Kz80XJ6aEO9OiX
il0lL0IIcxkU4bi/FfbRUa7ZF00yV+ouA6kDkRVUdNdn7AD9zvFHBEvgrH35Q38A
/EaL063FBwdKzfv+8m2NN8hQmUVYzJ/15Vu3+OuA3yP2pj/3QgUxjucvTmlqd/sD
LmAnTHNs0qfrwSO6DnOKfIJRRGQT1ysj4ADoN7sSlYFhYgJ9jE3ASiDNhQoLemn0
VvrTLHJ57tmsvqCuI56ivaLw4Ve21R58wyHKOhB22ciRRqmhqfXWI9FlUluf+CCj
Mw6INaYPfC/IWgR4GQwX/LGx1qeflfItHNqHEQeKQByjKjcd/wEEob28kgzlbexu
eAOlSDzs27ZrJPHgIEk735VtsnyncbXsgbfpZvUtDZqvtSql+sW0DpX05V+G9Sfj
q1Yp/TmBwEgRKqO6Zf+IAYun/Yo5zmgc7F6MwVhdnqgs/vJ1gnTxtSuhjRHYXfQh
sxsaBRifivJKlj9HvWazxvv6u6HXzF+QxOYirBDYkyUkL0FrD7ZwZJU3GOKVEFax
/FyJlV0t/en8B+EHbAy53VovXqqO9pIZEig1dw9vMOoZRjs7e1OAf0mKPfG5olHD
W9uKSIL1lTppVaDG3dY00PEk1GmTjbIeWstmL6J7AOKsk/Bwf0M/TIxyHlF/Le+J
Yq6ulRFU5kYmp3gtFYkRefpA5e/t2bVixQSbLucdqNL19d552lPzIKYOXsEUokbW
gBsUY5gOTiKd5Z2omB3NcO0z5xFI0S9yhzToPOrfgFOMF2jjR79r2KM51BDijgMJ
fIdp8Qa/bvKP4wrZN82GWYIXe8++g4Hn0+WWa2DLKnZBTzpnNZLt4S5tFiWyRmpB
nIq5QLTOdHsqIpGn9cJIq9HpftxjxXEo2Z16G6SCu4l1IxA4CG+/quT+9QFPYs5j
zXtVaZIEekbGolc1CGjqmPSTjX9rfwk7h/eOCzUDuC+QP9/n45Y+MSk2ejph32kg
5THrgNJyK9Ky+EIdZAgoNDfm8/mZtp85EL8wkijvQqzZW1t3o60+UvbxCL3hIDpF
v2dIo1JPnzg6IfodSlfg61bLI2UdrrEVf0JQaCyN3K7In2LHhEncrvZ+9q0lfLTw
SWofpxT6wCBK1mx8jdAXTDK8NMk/uXVXYMXpK8YbP4f0xfjhejivZgMOpsivCrSv
l2PWj7KpmVGyWUPUdJw3lIE5fNtt2oglRzYnM4aRE79hqWdRzqPgyGGbieyn8ipr
ylbe+xlctTij5oE1ggbYPa4/e041nD98C+9CT4GxRb4YneHSFBg8+sHPkIogkvgn
Pgv8kJ5b7F/gaX4mT0KSp0uPryvnJCfEkpsVm/oHrcl55LpR93tTMSuT9KB5mqdV
JB33EpZ1xarV5p/NWHGewH35LoMhA+vWptYCdBaFOR4FV43o9DfGbcU4hioQXDPO
vUoCLLxKl1/re8ANsKZIPmQEYBhRKZRiFW9F8BEdNxOWuuziUNFvNQrPD6N7imoX
lzHpROXg8ansVwNUocelHSy2ebvrhq8HUxHCr4Bj3PaEL13MV5OJImEKAt7ozVQa
Tt/qJP9Aqbgq9wf7HGB3JcQeLWo/W9lHVO9anP9DMy6UmWvSMbO4XTdv0W4kgOEF
Okt2aVQMYzxKWifZ+FB2Qtc1y7tkanFHmaOw6oc3MNXlWAmKW4mwYSCqJMTfplvC
onFSulrWzPDK7X/DN4e2FNXeDnt0GHKOqszLWVUX7TXhXn9WTNFweHiyqnE7d2GD
eHSNV8M9VbgcshBTA8amR8+/qH0/nhWOlZA4PmRbGBTlCdlhcqXdfC95XNaGic2j
OU9hoAIOwgMdKtUc+gV7AAitrQKmsvnyrS3NanpctQcOEbruF0rpieiSFmN2hQSp
dZdUb68frPAWmjGcH1C80oFRANeTU3ZoTemGjEe+hN55+GMYaZM2lU8YKXNPW5/D
wpdhRcy/eoOG7KS8nPQibSeauOv81zaU/+VTI7cNq1W94VilLoxiPp8c9S6G6+TK
i6HC1+pFs3cKgDVESTVj92+ojAdvtpUy9c/kK5R2wRpSSujmv0ivJGOeSCpLKw2K
W+zRLAhhD+i/qmPDBDWeKeQf2oPDP0yTv06IXbA0K6NApjIZwIuUvZXBIx8kEjVb
rLBUZLFI07qhkrjztB3ymnk7JBHwLyCJ6h6S1VLdN/aXxwSQLYPyqo9qKMnHKSUo
jbgjhE2YcWV9irdb7tGZPgHZxaRz3HG+aCAeSLe0iK5Votwe12pxZJ9mc5vU/c/h
rRMHprZoKawd0teiTzJgSCjqlvl5FjlNwJa46KN7OKuCBA9PYxcs2OEsKkSSublX
x/jp0orVpDzH9uXnHv4/CVaAeQOvgEilorMjyzsPkekyzLjpg2EWq0hZ7R31Rsiu
+0wvqVQhfka7OwO2ZVth+BnYvmaNIZ0XnTyVmJt1h9Urmd1HViutjyjrQdwb0PcH
7GCHzW/mDilFWWrGCLkFEyzaq3kzPpuo0fBdyXxiVZt1ZpNT2CKUoFGaisuze25z
bc6YTiz2RqyZ4nTxWYTRdfytvjW+8M8l65CFbt/3U0irddxyQFJkos1Uw0Sh4RKv
Kfb8jcgfDvgZO1fBAEkb7jeNfin7FitPlt1w0XFzRzxK+brUKGKUG0mmbFLzsoAg
/dJuvKXjWrsGf8F68AkbaPYxOxcwv6Q1nIGtaAUjyEK071gDo7vj6pZc3nOpJjBo
sUjOiZ9HUisFd8VFVETwp6RUyDFxHcP5LoQt4wwlYkCif5hVOvV8vwEc6Nb4oUjM
K1a51Q0gP8XRcz6RTgh7xeWIJ7UBTgSZwqxW9ZxC1pP2a2jNND1EDPtmnosk1zd6
e24cyHMvxlkdXvKrHkbgVNaIuGGd5/WZbzQYfnQl+alikPaEN2MqHRarlAoJW3nR
nOguJ2deylB+A2vJXIGTL//YlfUKzz5XXcy6g8pm9grfIuoE9hED08/PsaQF23mB
qGYSqavjNIhZy9oGx+hqoBSjuhbFFa1M1HQtpzO3lgG+UCe7Uyk+fE25K1v+02bj
+wSFquaStAQ0EBGLIBFhMkDOk2QgZDMZ90enYIGpTIJQbjn9HBJgmVGPTaGSg3en
URvFtwawo9QM2wO97hZqWPgnYKvvaqnrvkdq0TbcTKGWf0AMBB/32p5YW/GgB8ud
8JqCpoH6c9YKx55s6WkUen55G75EX/3BOgE5Xfd6tE6/+o69Bl75nRh60gfMWPs/
0I4Fl0cbRYzDdo5vq6lMefhM423puaBIC4bUv+w8vSVe8ml0GCdRbj/333P9hHM3
izzPdkcRNg3K4Tbv+rEEBT2AIgHJ2PS80JUgnDyUhkKWeXxFpViSkGNSWLN/YxOg
w9WlBvROZ9sv1KvInH7a3V01MoC3qG5+65YQrhysIjhBlue9OYZWMn1zoKzuCAkr
L8qIKTonNZUj9zq8R50/u1wyV5dLI6/4+JNTl4Sb1T8J5EA5Bus/aZbipqeS2s3Y
vCIpxR037InPC9p3mrmmFGNnPcH5lXDsjTBGV1hzZaudnPxr0Uv64MQmhBAqqcQQ
j2yKzdvJE6NDoEEWP/9b6LM4LJ0TrOFKtHBxX0lyA1JLXhs7Y0k1R36SNFpKemw5
203urwKdXRltUtm5OxqK0knlwzeCHhY0BYylXWjcueQk8Os934xuI4HV4UcPH2VR
ZyxNn8Pq71Ca/RsdD0m0Z+xXngxShLe7gR+BIoW9yFDtyZyKx1bnC9oT2RwuMQ/U
S7mO/eo9Fae8l3NSzccCcurpfQW5Xec9xI7YKM6At50qzhNI9FEter82ySnQiWcG
VaXegv4ZXSDwar4BZ87euQb98UgHUXE30HNMlouhiDUkUtrX1cvxTxC53he7sd3c
FylIusweIov8L3mS45AgVpJINP0kImRazGVLfzBMxQruJ4AnETZnQ+u+MMOYgJwq
3LjEyib4OJNat5/pUH0CR21jafinNuOKiLjRa4KB1pR+BNkA7eZ7SDn4ij7zvbjU
0JRL9ZGeFUp/UeBsSSnOZiPBwnityoJkaSECKx6ZtNPQoa2KKQaHf2NUz9DH+WnS
NVLGCqIgSBodMrl4/9ljV1M51ymd2hdSHzNFPDjVDp/T8ZK1hCCi7M0W3ax1yaid
A+lAKAbIcp15rEcAaFmPck7qprgXmOwYWKJ0aiykC9VNC8o8Z1ZG674OAkZmbCVP
3exCutg3U/FtuBHD/2AddWEJq91v5d3bCfqUh3ZcpdHmWplk+JYWYl3zVyytMWO+
wMVAfr0dOYubQIAy6tMlkow6LPUica4VGqRKAS8tVMz59eMw5sYnIi43BYYkD/zE
MPlmB4SsJzy5hPV1f0c4VGEGxUqL0UXbjq2PimsUxLiQxs0B8JbzADgR64rbH21E
ad7cvk5qh4AXy7tW25RT3gJ+2hXbwCMQJOxPt/DhvDeM0R+EvLgSgc5LTXJHtwGq
7f1vt5HhepKt0Bq207BmFeA0LEhGyJzpJFShPsBUcQaOOUe/jys4N6rC7/SoTeg0
NaE1CTUvHGiPfSrW+S9Ig/yH0BX7LuCgr1FCmJe1TC4j4Osi6lAM5bi5HWbeoLVR
gavcDfN4ep28g1fbX7gPs6NjSRb5h+fI1WQUXwazNppHvyiwFisA154grmJ1Kjkj
xpOipy3jDFs2pwGT1OdZK38lIeE971RIbxKPOxBrTypqsbIO1C0MzpDdu9MDHciz
WBL6mrIEFgwDP1GIZjidar2vPCp4bC0K5EwAPX/ZucZZSyWKuJbpVVhv3S/SBQXX
0k5zJDidxoDqGzXPdfkUXnVC/6E8IBqRY1SF+NLF9HX//CWBijG15LI2WF/pgnav
U4iwHraES6BTNoWliJ/sZr0qaF8IAqOFimQ0KPqWFvgVY6U0gx2b0eTdWh2vySi4
5xYwkXrFZyjFnDtEmwovsVXy2kehEOzOUDvgVFAIkSGg8xor0Nnik31AXcRVHXSp
SNzdyCKXEfYElD++HPK34Ml6ns6k8EmML6zBOgEVJe2lZtptcoeyWZIa7Bw4l0vp
IoinbcESyfwJScv8UKzB43GgXS8UMZG6gkByA0hPEbPCk65zj0XxmGIdVWyVWNQz
5xyFW3t90n4z/26Bg5QLitnX5YjQc79TEaWmZK1uNKWcf1CnpTSMcnQBHFCpNq5h
vs9Q0ocMzIXyqHhuz1wt2cOlNdXICWp70ZrXKDb7LOttEze32YYmHnYmdenAJWhE
Q/yjhHRon3dnkGiDmH+e7LQOqaU8d0upXekZLczYPyB1+CdOt+opaU5UgUhKX4WL
W9uUSz7Xmip56qrDHJXfYR46HSiztoWaUYukmFoxhk5L2S6AprGljOnYxd4/R3O0
cPTJ8irtAWFcJx3mfM4OPySUt2KFie+82+NOUPHKo//aGZ4iGZaYCvUZYU+3I72U
NZVlhV3cUUXRnKfLNLcnatPQfDyr8l74JZL8e4AdT4VDlZ9XvtovTvotk46FpYnB
khJzjGYdRpqtwizE7Nfp4NyQPUwwfXq6Kq3iiABkhVIRl+gDwWYIb4tU7DjEvpd+
fLd29k6P8uF7JcSbmjcHODATtOMR+oLAsZgd/Nwz+swDVr4hevEKacSfVcK2Z8ET
Ze3FuS2Z5U+lgWN+dZ1vyxFqC/qdaw2iXsTOxszLLNmhlWwU1MZu4leC8+d9c5Jl
z6y7Fv408QV+vDti5C0ovHlKUd+3mAvLSpCZY5enIqOOHpxy7sqRnotxjS7mZtE3
jKwnOJgnlK7YXNj5dxdrvVMFVTPqSOBXBjby+82zg/lUKM94gXGz9t5WLaZGmkQf
J88Yjyc/idwZFeD6dmCFSwKoZdC4lTDzcyvvTxEvDFNJgbqUEl8v1X3ftk286GFk
xQwutwSCwjMIT//fbZaT+lcuHHetl76xxKpGm4271ZQPyEJ0RzwaU7tfJcrMyFuX
UnBKNeySv7VLea2xM4wN0UhMz9xiBY+pLncwWnZ86LhqhqVelNm0WhmXRs9HYWgn
5+bss+M7zDx3fu86B2IDIMvEVrszztfsVWmSUdTxaaw48ljHbGFvrTw6x7wNd+/J
F7OJsTLsHNV7jPdYzcd+pgvtEtdnkl2xjVxFnE068ah6u91rTTzMQBZhU1sP44uy
F3TO7KzPAJjsP11TazkDjKKqNAmAWET/j3z2RIUSHHUG1XIBjj62lLEsiFSxaJkF
D55Wbs8J2ujQSwKZ4U9AT9p/waxmMb58/ayo08kaeeE1OyAt5KTki9p1xFVMwAhL
TNbQPOxF/5kwK5nXLMJwMgCimLVwZPjEgsztPUjqFzADTAw63nnnPhN2qyTvFeGL
iiQ5j43JlIR7V3EYibUB8WqBWNnbwZ7BXNoZkel9c/HIHSn7wxtEM3xaDPmE+KxD
5AQ0XPS+csUxGH7icqM2hpKfnI/qu2GNEyUlLcEECP9tXk60HxeEq0DA5mp1nOGl
ewLVCWSU/Ug6BWTBqkp5zgMPS9vTAL4V0DMVBEk6ByQCNBfMsjgRffVmQOqd/d4T
xnUrwBDaXX3dzTjcHxTZTIlYowMi2utGClVvq+fExt5s7LZ9smp55I3NitP4RbPO
uv8GiUN2P86n7s/c5ETVN2X71Co5B+cDfGIajXH79e7e94GwjwAixQTAn/ygVgK+
1eQPgPvfX+541LD4kpjF7420rOyR2txbyHRjk1Y7MiotobjbI7HAkIgGRT1t5yUm
bCp+tbd+GCBxE7FELZJpH0TLOK1lTYCwE/t4rulxCzPKSzc9cYfehnuEK/xz8Ba4
EQQmdSEzQbo4eypxDVSXJPzXrvgJ9d96H+xXmEWKv5w8fA2uqjXZX7/0X/fJOP6m
M6pFf/QuwEJkuOraeOQjpaq///4XtKF2tlAy01oE/43DUykG2+dd5Xccn3pQa3qe
nHvtFAgeU+EaRCgyvpoFUp+2PGyQGE8ngvVC6LGgglvbGCS0dVWWGay5PtKAueZn
UgLQt5+IX1Qe+U7samw57UrF/x5KgXPyJnjUuhzpkK7ESYIZAKY/pC3UameqVpv6
9cn7CR6k4v++sHL5rNSsiUqQri2wqwYdL8vq3O4L45e3VOQtrEs7II+Cy4h09taP
lDieB/o+xfo+WjUyQxVrzSJrhliRPELr82FWo19iWK7Af5wtsAOTkELpneXRSVEE
XQrH/0nRY5h/Lh3ompWarWLwHPJbJX+Sn20SNUz6nsOv3nrs6KLCkB8azVStSRop
pA+wiC/gutTsIj1Tm70fe69JPM2TmV33w//AvKZTGitDJkFYgj2S1KsX4iGaACn4
L20jHWb5rwoPwVKy1CHmLIbXj3GTO3FKwcQ77ui/aIogxtVAoKHUWdtbKYSgqV/W
fbdBCL97sYC21sLBMfHOnLXX1bJ4WqMsyRgvhV0yN+YkdiH+CCabTKByDsempl74
q2pTNUy0sJDnARz6FZLCuLpbqoGGd7Nt4kYz1heHjBjZOYcws2po0SSKa1f5etdG
Cga85ttj1BiTRRUd2ymdumnNPp9NR5w6PTdGBRbKipUX2VMBlK37WTQRnaond+aH
OvyZr6yRmkNQLWEo7zXjVvmHeHu+vLSFPutDjoHu89Dm596ZPCg5ZQUy/+6P0hj4
okn42mysqOIDHQAHZbMLRI4C3tZxnTIAl+NdZiQdD40ZAl5tWXhkaoT5rfm9MtNJ
A5cukrfzZmzyQR5Gp6kXZu+5T8fVn41tN1Fl83FvV5VSFEicW3RVVmPmgJoiQqed
FVR5pt9CxlDnXuaFo+1mz0tC1LDnfC52knCmNzOzyt+kwZm7HuPBhnigEa5sOPfm
kuZ8HFi5bSGgPjBHl5QGC7TrPfvWut0i7FPlKwqTpK+Lw7JD7Zs2o7Pr2Mliikky
y3qrGjf4ePu0HVts+F/pTA9KBaQSMB2pMuzE5gMzuHITarpNKOOsYf1Z1UxOqm3n
Pu4By9l48Hz3FiPccvo6PsQaJlu7Xr1YMVvAR79CFqo4UVXWyICyXUoTZJfSYfnA
kxeMQcQfg2NeM0ECryl4sAM70nZHGkwTdY2TNiLDOOA83xzaiz//XGN8wQLsrPZE
npifUSegSt0aV8BcF2Co1DRAcDxz55obnZtCgeYGYKl+OaZugXK6NUnncFJ7Padt
Z22KLvWn3kYX2vVmy/d/dk/XzLZTJLh2qiCtNiBNNnZ6QgiqU0BWI3/14w/ItF+A
14dr170pOze4RydGVT6orK4nOEhbTDzpVSNXdNE+AJNqHzBQJVMpKUIrsxZVlGgy
BkN2kIugzXVEhlCdAR3F/RUStk31E8zHIi2cILinvPWlxHxGh285lFrMEesdlRQ7
ENOUJTEOtCDr6wiT8nv3q46EoQMt6HMOmEkMJYga9HQGqmT0KS1wvmdh2DmsTcIB
eNBOq9cbW9/9JKJSU+ouvVogaFcKXP+wnNLfD4up/0ag2zSD38/SiDlcKOomb0UH
n19I0CIJLOJqdCAP2dnmYQGUeXZJ1XkalID9E9rJz9WSYJNaEjSLwRb53lS64xma
fQ5toQ7s6SJ903JpZ4HRQqWxe4Y96Sa+cn78TCSCOCtUX2djNBMhZ3Av7/Wyaa24
x27Fqq3Y0H6F1mv3xXWHBGKZZNsKr5iU5aW560zox5gbsFQvOGDFBej3FrNgwVQu
r8lbq0/Hblc/8H6GsfF0EBEBwIZtdEeAXYg/gEmiJ20gBcnMm+GgJkFzMg8uGjlB
YmS5Z+CtGBY/oMhlnGbTFwBcQ9qUD8tjgv/UuaGL2lSLrb1d5Zq83Ac5zisbf5rh
YxWopVnv4PUCLYTLUNpJ+ijr0P4/tY/N0EpPOMPvBdpsqOp10BSRKC7fc1MLdD88
T41QgQwl7OBYo235hc8fxyllWfp3Wsvx+tSmRQiBzrutfmkzJS9eNAwiZbT9Eqlj
120hSAdWonG3ZwcJFh6+SWfNVE1PIJe1KGftkaP1DUeNGD8olzkk0Rjp9dVCiCR8
s42mq8zUoyyUElKb5FI52ja8V1CV7nAXl5aoQhyIuuYZ4JFmqc/AlM6U9N0cuFTk
WultAQ42jWgIpHS1Voe+nUMM0NiLskGaVPKFfxQWfYYkAwo4lNxd3WPtGuUXOoX7
3ipiicHqqIwzr5g0Z9BG41LzVrbqNcy3A+/GRaQy6MMU28qlW7HSBzQYmg25wONg
GhSVPwBareMZhcbb2eLCtdRVpBFAOASfhL/BUbQQU43abDuN0tWt9tlzt2f4QR2s
Gqmqmm6asJtQnIjkE4jw0NdIpTURd2Ff92Dj5Z2bZ1DjbngBQ+aQ8GMbOFRAbMEx
++XnRvhhHVACyApr1M4zL/EYjZZIVzgRqoth4anb1UppY6egPESNhF2yirYa3ajH
Y3BSSCrO+hPD/mqom77IGSPzcLXvyQoq/+GL55iOfRBE73YwtqSG6DtCgDV4znbB
r/r+dufqT4v9sqvbgNPVDx6Ry2p9M3FB8POK1FQI3adglVyKO8B/6kP4RClsths4
8wH9x1YEbEnw/AsyLnGPMWi/54AtvTw1eDQU1jiUS1CkoO5dwEqk/Rs8pFbj3QjI
h2QtCcMu1sXx8cK9GC8W3bCM3FQNeGFQCqx2hyAT15nRs8k4PV9xgOD/Fok1ofFu
7Bhwh0op8PGk2dZqjo0kSrMdhHA3oIHQYKdgtVNTEiALOZM+SJZ7096+4mo444Ut
WoyusMvVOzOT5i7EFX4asrrZKArwWE+D7NwI9XigXFZQNi+YcfB5mPiqOTlWPqWw
yJZho/9Hf/9BVtVNXG22VP5Rqg/OoTKbR4xphSNJ6nHlTG9GeTZQhQrVdG7KmYKK
oLrbjwE/bYiqxNG3DcRDPUi5i7Bno/3i0js5ITI9BnjxO03G1n46vaVwgwuMIy0P
zNxDgvcIBhmhSP8pmuPHCOKtblUaJulUBhJP/dTfQoObkiPKdQDL3qOVTbWPZsQW
d/pZVtNM0ZJZlouDXKfNQWrWGXBlwVCOwe5F12u0awgiQeZLIHUokKmM8rsCMxJx
tDWJu3iqWYrQTnmtiNLghdibIOnXkJ6lH//obgw0aTsDNiXYFoZwIJdAiEiPqHbO
ENakA3atvLECmbARuklpstwITZ9IeYbWbPTOD6qlRCUy6N55EV02Xmk4bnLz3wTT
y6RhSrKBdrUMv2+7gn6y++ZfWnOgQDjTaemHYzPAbS6C7fJdDN5ifX6tdC/NAupT
3YBkwUKfI5aU74VDWb06LytXKUO1108Nktd1QCmx5V81V162mQZ1CaN5hdl+7LxP
+kYd1CbGcEl/Ta0Q77GO3/Qk4gE1vaewuJBioXGAQbeTPbXt/Dcf08njauVA09ZD
ElvD+ZTUHmjJ1jaog4/gPgKUB/F5eAJZO8TinW7mDjxlxQ4R6UMDr+yaH4Ir4K30
LnHBztQvZjIFfrMHcE9L6Z2BveM8E/wvMUQkImoBfQBxccoKhS1vD1/OulbbWm02
3VBiQUlkJko8oT7KfwBPVMHWHQvNc42B99t+6XyiSIpv1XjmP9o5mAOCwaNHSMiI
XVgvEQ64POibQAqQoZp8sregef6nBPctEnFGw59nxxbDSLXB8oXwIlljp4CDxZ7h
oZm9kZ3qxrLNGp1QyUlQRSCXBZg+K/7p4MNb8KZfqxBDET2yDSCdlexnR9jT9cWe
CBHk83Nha7quy4njVsZyoP1WtyykGz3Amyc2rcjyUYSvEIK3ZGeYXuLai8O+EhGq
8jFxkTszwOAQND6mfGnTsi3i004U4prZ91zGGoNcexkYDzfnubEh8tZLSxfWWRCf
0DGWGgZxDLu9rm5Vnwn6q6ZCZttEVYuVEYuNUSle0EWnHRlbBqKIMXXz0BDWvERb
+ltvu0mQqd0EOr0vmELQwtXkPoEVUATYlrTJyxeOGPBIwcdLGl8FiCpHJuCqJN0s
8kAbT+uMc9l9sNgRAQCvVnk5nZnW1wGkDpOuFdWbCrLyfXmwM87qw6YbS5BKo1Zr
LYbqyyTO0YzA5FVgFgHPL4VSbMuNI7sthIGndI/jNcnUsh3lJPfHdWYf5REFgl1G
/ShbLeXk1CQDA2J2GnZ5XtzVMUx4OFHUCiYBvU/MvXrRxUxxLgoEVLea1k8cirfZ
HZONorM2twaqvHbx7o3yK4rU9SjSFUOO2IZ+D91eO0C9NP5bOdnWwAo9Mme0BhY7
AUkNdun/AjoE8ozZdUnWbvF8uiE9rviTLr49EIHUEfnm+H68pyJeTLur7S9mY1Me
dsoF4JBbtSB84i386hX5TzmTR2qIS/c1n+irRyEkX8S2JHZyYhcR0vvkblDxRTXz
FvGj8joEAkKlUqY8jk3JxBTjRxxxDAolol1AIhMiH4HEui3MFbgUDTN7uJ1B3/Ug
yIXvEDxUGkcDrzH47+DXPEIRFI9/X+7Fkm2wPUN5t7QiOTmO/0qUrxZ+BHsZlGi8
yNPNlVqORpW1M5FDtUPPI4OQu0w7xfzRfdcQsXwOaJy1uEhVqi0hjXjzua9TYWM0
Zv2y1rG8T+CJdXTiFp5H7vba/8ASqp9i/02OXctMBkWJr+dy+M4SD3DUk/VKbnV8
rHKKwQVffySZbvl78blGDekHa9LvBwmqk7j/fU+mRG0M1JpDTnMdFKNOvbg7pp7E
onqZtv823sGoYxg571lZJ8kTjQuevVzB85jsEwJKayS3eacrozneVgJr7UvxmMc9
qR5t+iyZ0adx9Og9lfPv8gOrArcUSnI2KVZ32qHiIPCK55lUYFt/fuJ84sM7Ppwx
zvckX+k1Ja+dq2IoYgPW08q6QMCH3+3vtnjC0XbyumHLUIxp64RO4zhtSAi8SOGh
iIH6NfPYoAUV8C7vYt4rLcZrbOXes2Py6H/6tAFQcKnwetZX8U1tf0/PwTaVtGL7
4W163DFseABzEw/83btGD3QZAufD1GioQakhJ67yWvHF3j95Rc7lUBVkRFaLscWX
qKGlD96l/316EknEQrwnnQHhiSObdPvxHWENtfMcJSHHi1bnPN13qfpDDhZ4aeRn
9jIgS7BHPF6Cyt6U0BwWZMRblx47d86Fi7+d+hDYTO5BqY9mwuU2uZilLQO/7Uqb
PRBgsxEVpsmCLao9C0kaVIOyjPUjuqtWNhhQ+fQrgXz9spKCtgLLgbktb2IhSKpm
WHxa14Ds4dfzGJRmHhVVZbphReYAKG+1SCgeAYmaUfMBBR2LgHpbqU6XSF9KDQ8C
nmmcjfpaa/EFF1VDjDBy8I28L4YkZa21mBOtQKElUTvvvrpAn/IB+5DJc9GxaCYD
6yQb91AJmwt9/vpMCohTbL3MDGhyZd/9yDkkb2CQmuiB9Xay1GTOiaGpreoD+TPe
7m8rjIzN0Es6b3MDgw+w/rm4ryaVqCyMN0rD2qTjWDYMXNzidg49F8JRSu4HMY2r
zQZJwnR31PMoM6pLD/X5TQBjC6JEClc0cNm2pTxuApsKgfa94HNBhmZ69/ZcaCHP
ZIBm/Zt4Z2Zx7kJbEEjlH6D8/adyB6XlPaOzjk16qZZDUHT8qV+fh3nHiyLWcd9m
DGWu+thJ9yONjqbLcuvRYdz8su3lA12Z7Hfnavv+csVnCsIJh3N1GsUxEK14M62g
GH+O3r+udNG0NrvRzSpWIPFWsk8rhL98e6JMinJJyiy9jkrMUzHMr+nwmrlyICyi
oQJtV0+hXZz/UGn3tZNOQiFvQvPOqcBMTqsBnB153IVCpiL0dSXSGq/+dnWY7zDQ
oIP8t/gn/DL734p2eAv6W6cqAZisIhJ6nE6IHDLlSiwCtnED3Kc44gCz4ydk6Vff
u0stFwGu+S3TPFwwkpY5+y77hIFzRtt79FjsRjYhrXDXOZagst1v2DnjhJnQZf3l
MQQkumPZWJsATPbGx6PxdWjywgHM4ukcID1z2rDtu9y2CRYyMqK9b5CExa+Rsy/b
C9Tv5sV42sDJI5TX6UC3SYfKx+qU49rSXvEROMBZw2M6gQs16s6wrYFw4YtsYBCI
n5AwfM5Qz1nz2bcN+2qdBSfVXN4nsS2sP1lmyL+r5WSg0y6pCz7OrJKS1C+F99PK
mCnJvNfXhCa+jIkhGzm7U0jJCTSEoYl9I6mFvoaIgwnBXwPYbgQIfcUk09gwwSAK
QhdGGWeGn94ijP/xd7LPSRyCCPRQyAPtV8fam4dsCb0hGthgOZAQ3JFTtU9kDgLf
0ohsvmhRT37Pag0lpXzt5BK+6DeQtB9Em8IW5hO0f7pZsGmvxRd/4AO+if9EUvhu
9mlYykTw+EidRGsf+OQNRm2/ADPqW+EpJrgzZA9Ae6iWxbsrRbHmXVA4iQFPJJqc
n7GDN7Uy2phKed144kEgSFz8iAihL+n6FibAQNIIchB7GDIIsK43MPtcx37ncgHQ
8u57ZAOrZ83Hj63KU7JmRLINOb6e7QGEJ7c0b4v57qujG3H0LALWBYeSANn+1P32
7HMkU+AhrJs9RiZROv8YvVBthderUto73BRd8/VRXpzmYRVQm5V/mZgz7LOzMkmT
Bme/v11y2fTA9IQphgHWq/sA+zJ5oLWRsqEN4WwKFsjzGtOmFpzmflspHLDtNIRf
j3D1Go7RQDOEHybdGUrodpee5L+dxf4Lnuw0QUthMWa8ycLfbr2L7FRnL5K7n2Bo
ktGOpq55R42nORxOf7uq5t3r/aqtuTyUyD51BCw1jrz/Dy/6DZjmautNKQD441tc
5Dbgaee8lr3RX85zy0OjDtyI1JYxGp2o3ockvPOoQ5EsoQK/VZirX+23XvZ7x1Lx
kFk7vKe43aeY0p6hDZ+dCqytZkrzr4+GLoyrGds8uZX/UgTw6dZwL5MZclLRHcXw
Tuorha6w4erOL7kKmkRhXcOQkO+nmvuvT0THg55VnM9Yd/z0SArkOLumAmyNfsgr
3v4AH3bt9armsc9wVmDcA64vyvjJJebVQCDm1wkN/u839wXmiXXm7pzSM9QzwnkA
NCmn+DymJRW6CQwNB1jZQPsOzpsIZLIBONoKJsqAU5K/ukHCkSppcvVUc7qrrUO7
jRaeJoshfh2lVV4w3bPQXXCypZ0BnpFVQisPRUZ8xbcb4v2TPdnu3AdnbUpEBVpy
b+bBrl/vi4RcB7DMYOzZTbDPK4kCKSZSE1kxsUYrqQkplHb30/UQeQForLk56GXX
jGEL474WvFZsxJ56Twx/w0w0u3kMaCLNCBjzDN/W2KTIvWFr4MrSHMNS7aGOHLGT
8kw+JSeQz47XK5awBFBk8YtgVJvCVoAoRrlZQ8Eqxk2wRIH5iVrN7hIcEfgJ/Jp4
WXyds5CYzZOwz9s3rmiawit005DwVUMNXmtGPBPYrhRHiX3MQQI5KEG6IdMnsm5Q
Ss5xYyhYM8Iv9k6eDtrOf+Wfa2J7TUl5VkqhCYE/KSyodHr4YB7caspCQ/Ys0pou
WAGznHIi+giLADTFQAUzWAOoXyaZJuRvXCD27EPv8V360DFiMaxWsCxQ/L76q4OG
5bchKRbT8UUuTggNn8o5ahDaSiymufk/aCR6G8IwApExNV9jlchHL+V2uRpl20WN
UDCVavmSnLQ1q+NLR+hiK+U3IiT1FSmHfoPyvW8Vcy88ci501kO/n8esCTI6YbHW
D7ic3Uh1tJNpWa+Q5uYbe06YL1i2oqxfnViJO/ruaT3uFwidNUX3r2a/hgMXLSKV
d/2c37lgFO22R4Fs4Jv9TNfZpyNFQq8Q8DAGsE1bd3FCgFmIds9LcyUkf8++azdP
kHl2tZNWbxCeSvakOpOH0qr1nIvvz0JK1C4u18bObBEbV55X7kn93qFaAkuU9UBa
EUNuTnKxxyT1lNahKWBGi1YzxuhUbIeYjY0uxKYhhZqvbPnfSdtnuEbYKEz4Cwp6
4U9/BYF8Z0D+HDJYgTz9pRHBTwjujO7N/rxo57x+r4WQh6KNFoU07koyuceJuL8f
ViRIeS9ayP2aJRT8azLL4eflka90PInQmvD3/Y5hcdm6r97u/3r2lVfU2+rPVGnj
G6DUT6VzO1G3i8s2HONHSBpAKBz8GZKK+apkHwwf3k1kQcupe1+7wMxT5bLHKzEF
m7ttP4JNxzJ3gZtSt07QpDt2uVnjhoVZehg7tUay7drcmkVo6smN1wbyz3yAfBNJ
yJxQvminx1EiiQdNLWGHUGo10sdAgtryN0Ezv1/nqAvsQhlf3Y1oewEUhbz+mlsQ
9i5LL6ZWu6NzTHBdywt6z8NyJ99jvfUyGouK8GIprYHGvZWBoLQOYfbxAw4bYzB2
L+Rw1btW5szT0uZ4EyaUcRvEzuLwEhd7HOYEQ1KNlGUrvxOek6BkviynVkXyO/dY
e4GK+KnwGOTuO6B1gPfIPhLcZUFSRtYS2TZ37uHF25Vfow4MHgbdwO126zmmagEy
IUXRtq5utY6ZqnrzgilGRasFKFDv8oZt/9zvTmC0gQDE75kuTobt0pYYiERPhjjB
wXPr2XtnsKaUOrIp2kB7dRa85gPA1bv5QCQUIjc5FNIWObr9gyn2Afp5GtUPGZq/
59xiUvu3X18KDZNprg2lZwuCUnDdp/LITZrHAyOcgg3gP4V63g7YEDI36bjrQ4oU
EteYjQ/z0mVqgA3Az/ZzSo3D2va4//mpFxeVOQPYe8MazMd6SCFggY73ZH3rnZ15
Rdgfh0ll59TWlDSZGWCkI72IweaU1mBYaSKyVTmw7KqAUDZ6f9IA/wDB4YCltBxc
oouL9dOJ/2jp93AnmTJ9G80lUQgBaDgvmTSVsbqE2eR/PrMUn/5f+soXFlj9+4ub
g3TQS+Rt7iQlxmWIE7irF7a10h1b8tHARCYVl9uNRqV9N7HU/PJNIksqIXDkKQ7o
/I7Wf/nrdne/L6MGSWXW/tJZwqxXuko5jLS1KW0gQCTcJEfzFpJ/qftUXrgqGICj
Mgsk+iqMUP4BlHZZUwDxVw9gnSTf1tFiBfvkek61lida3wNQLupL0aLh/cecvHOJ
dPJ825gMQZvM5bkev+GAvBWaCFRJYst4AyK1anZ3AApi6lzIsfhOI4wyK4H8pgjG
jkCc33M5nuVkovKmj+WoH/ODBvqgu53eYB0ahrBunLxpz+2Oo6fdxWScvCDprpix
9xt684cWT0mHpb1wF2cC3H3rorLBGJhGDbwWLRR3yYgPE47+vyUfVnkXfmdkIQXa
dnxAKYdCNE7YVv3zlxQpArpzhwgQT4pw7906886X0iSh6Dc5bww5bHVR+pmSoa/J
bx92A5bpBx7mnDum60DkFJBavP7yQW/JXneET8DTH5pukNNuvsmgaoZCpIkINvvu
BNGP0QtJP+LLmF1LzdpB6iNcMKAmtmPCkEXxfh3x0Q4aVMo+R76H3ZXIoJfMDjaf
42ExvdCGwpP67zJhKmeI/uefHsP+2+sq+2WFl5QpRcNxTDleVVQBA1wwcGizqkyW
KTdu0xgnGqx3KMsag9EaVQMuxYbtWQ2tsOpdSINPQXonQL5k0Ex9+VBBRXSd8WEn
SB8/0Tq6QTDgBSjywKbCWy+uv5+LPbqkCh83qNyn/LKogWBPXvCtHHAuchIs5KPq
TtWX6kOiLJOigi0KSO1V4Ne0OfjaUD8oO3vHPeDRWtE/HIm7cP2wV9BIet+DYmBQ
MvIBwYCJOZn8toKoHoRjIooeVa8coWZ4uHIj7eU9t2Umpw8ynN6Z9u9H+QCufbfY
ScbrMF977BQyFzX4J4Y5jtbeepsWlN8uH74A4rzEF7kjS/DrTEw9RP2qeyFcMqUv
mMdgCJIQdBW6ma6yi+rZlloEXUEVVgMjhFIBNJ6iUhvxEKDVa1RjpjpJYHdAu6bL
hEFjPQ2ks9g6SHkSEPcYIubQM/uyFr05AZFmgp0vCXg0KcB30XwrWtuacBTNMfok
+ddluqzI3R9nGyY5Vuv5mqvA/mggU8WqRoRX+WJWRjs1coCMNCRj2tT7EkmbEn9Y
fMEGyqZWXlnpyfK0GHVAYf7hLTf0ozOa3Zy82i6ohaKUdBXdwNHG2rx9veO2VfwZ
jH5sg1Km9OfXe2i60PIUCDlcaq2NR7F/WlTH8Al4wFFTYAl/jhY9BqDGHwiINh2/
LuQlqX1fABsbi4oOBs5iTWfbXsfeIidV4YPcsiQabB5Jplm4r3YdyR3jynAQopTF
Wj5VjJfs0w0fN3wvMSSvFQyLyJlnWbDUdGN5xQq0hDxl9+16/p3vfuStQie+fwpb
g39fH6EBCO/0nmRGXees7oKGAV9y5l5/bULZD3QD8VcQzsrlmcxzeY2h+EwGMxWB
mmWi4ejBHaMRv+v7OihrHEVRQhwmoyPcMDEr0nq34qw8mfAxCOvQYAaqVMTjtJId
Oqm45QvaBFV4Rj3n5r9uvm7eUkuJMU23QTumRptD6yD+aSzhMs/0IXMf5SUpZEFe
Plk+RTY/SIjIb7dl6xWFr00cDT8SO2yCnKl3Zabsj/HuCF1XhDIeQcWdgGIffEHg
4jQs3ACyvk+O/IG7LyA9PT3Gv549EhfziI4rxZaLIDbdAqDPDArwzAqjFKiZDtzT
TlqCQyGSvTnn0U1uUCVN/lUeBi4VNRTW0USacXJEPMToDw30kY/P0QoBYAudOAXh
b3YV073qKiBL36/ltbQ8WfJZcBqEIQy7a8g8zM6V+Npq+wLLJDWiLTFXGv5hL/jl
OnjrSgeSbGOWKB5Mu+nxztT5JRljTBl8yZAxMVQnYFG+Az7pciYzA8uIYC61IfCk
y+OzgDc11CBXCtY+v1/NPSDbNP21XYOehpB7b5aM6djNnR28JG5dqp+f4TelS8H2
mzQnfDVF62wrr0Np/EjvrVbqcDYe+il2VnjhHZw9x6r1jWpXz0TP5xC03NSzzuFa
ExSdGueWjavMy0Q2GS1mtpH4g/+oe/qDUcsQJ6lHj5+6T2SqD+6QcaM8X3mM4phN
VITvaOUPD3lu9jAHOXFeYoA3SI+bhzLgHDEy5inOuByr3JIgSu4tGkGAqsNjRa90
09FRHTrR+G37DHmNFe6bU5LDK5qGzKhMPRYXPQ7db/+3WoqHNqy/eYlAu+tH8FKD
4fK7gVfclkg+RaFqF/R4SWVCRIk8CXqNDDkGQ8u7nH9glsDkWLoIl0mcJEMOqWL0
AiXDTwXWSX5b9K44e1HC7Tpp9tOG90O724X0MyPEwOg4l6hUZ1l15Ay5jw/ce2bI
wlfRqpIRgE4fP+OgJMcItNNo7/pTxli+bolRQ0borYtOin+a6ZF3J7LC0odIyWZR
75iFCkisY+PsFBjaGbB6lfV9l163DBnpVrvGSGkCiUtv8/qOT7V2OmIsHOCO0XtS
fwAA3JzXmLKIcnJhVZtMFlLzSHQk7qNdelavD81GGz9QJswkOcgc0CB/qe5+PkuJ
oTDcrFse9nw/Ab/+p8h0CF7lTxTYTSC6oKJYhwgqjcBWT91JMXD2hyi6YKEwe5Z9
D7hhUvAUyEUhzPUJlcS0N3Kbhxn6r1XfVnSk7Ly2hw7ItU6HVbR70vLSb714zvNc
2Nd+nlGjw/iLo+UM9maN9MjpF/TVQDzIGaAZP2+4E3e31rSCyyM2qNFiyhdRqKwd
llLLMHPvPSiTxEMqu/UVR4U3h+Qg4Fz8aBYbKVqyyeWM78MhEOKU4Fw4NovCsVqj
6movRLTB3MQOZ8/wW3+J0h4cwgmr+8/EtKe17G79VFyKxr88mCu3UM1MVW/LRArm
hSRuZDkV9E000y/dAm2fOlicBPliET4HExRhCBh09J4m0RdB2osaQjdOUM3iJe5k
Q4eBjv0+FYU/yuqevjKk5tWHZb4D/eCSUpt0GVsz1FjAnGH+VlUpamRJshk1VEH8
4KwMIy9mSNuz9ei6sGaz4k6YETIktsMS/cRyu9JlDKmjSY1sAyUYlqFMUxRWybre
kHzX4JiKoWAuI55qCcKTU1p6D70EnBuf+2oPAv1teCuczsb+IQsDDa29TM4LdqMI
Q3kyQUX3/0engfodRSv3yfyaaIZ0L8NDvaaTJsfYA0prtXb+0AbYZbeiVD0+ecMG
2qLwD0I9qRtUd2inGnYjwNBbFAG9mixq/4vBiFqetjPH6MnTTWQ5N+vtCsucOTp9
WlJLq8Y2uG4o3Ue5WSc5icNxRkKVc3i5oRL1bPE3ej2aXhBBWz99OkXynvmOf/W9
hAbie/dbtEsP40bEIJSyOj1f/i4bGgZ2FEzKtq03b5D3EEMdOuTuWWSffB5wv8Im
WqWJqKMdffADJ5Z5qw30kWkvUVB4fv4Kcuxos37i1r5ORfwRnnO+YonV+BhCITBt
Zl0FXO/WqKHMHLRQ/EltWvYHD0j1z/Bit4EL8QyhJcyD93XpwabGGfQvryA1y6Fq
1IAzonN74TBgSVrxx/PinL25gandL2vYiq/vVEmT5qiWcBePeXGO2de+MZJB3d7U
S/+mCbrpV0ZsnAJvuEl4Gpsd549syGUi49AlgmT+im3Dumv+Ku9mIz2AyEQIUJZh
IuNzQhJ7CCpCXOA2Y0nryk69lmIULX4edqKO3aGFEylmApmIZOnQoPURbh2JclOz
JNWV3IJeyjcCUU/IcfJ2KF4VG6vRCHDa/pkMk0w9PesLv8a1MoyZ3fokx7mZ80/C
vGWeDJCA1U46R8xhdHKIdHwDE7umr3e1thd9akyGMlNtUpECyS9fKKObnBj0nFhc
SFyJ02aP7uFMmNKPXLbQlRYxinpqRg3BV3hLchPm1KwIWQPpRiNaOlkuUR0kL4SF
ZMb1VApWbw377iEZLaAjARRKdhnIXaL6cAyi7LE2GSiJtTT0ioic+L0XhFbvz9T5
ZmjXNHqo7H50Uwe3atUUw9Zlr4Er7FfI9EeU1t/wqKTdsMlnfTkOQ7TmbnUtIvCT
t6w5QSa4edoegs7cnsX7KRCtlgv3KABmwZiFprn/NYE2aMskZTS9scgB1iGsmiEq
qGqy2YElgt3PVZAI6l5se1fTpqTxEQ1UnlW4L4OMZH8DYHpqUPVh6V/7qvL3pkBQ
0m9lPN/dnQPUm9SCeLUCUh9GdEQFEQI7UtjZ4Z3ChWEsUTjvKxEdH+imNftBrkz9
KY33DgWccpCN/33f54PcH4qhhbNFPmmI2DRfAwiyGdafITVYEXYTGNwSbpIpeC5U
ffziQFXRGe27owt/VMl8Zkpn8CQd50hdyBINwksZPTUUU5k7HTUfWjUEsbb8+9Uv
GbKEhD96m0a7Vi8wRevQ/g8trYWxHMuTblL7nAJ7XekMLOha5h8jbGaPfSf9U3Wk
qWu0K8BLZomu7WhxQkShj4zFRATnrDrKZ0dEJmR9V/u8Yfbvoyk4pnPvLOeStFG9
LrnswFjLkPc71suCcISSikCaVxsCVqut4m0XLkKnLHhjuPntcHZus1dYFE9CPZHF
N38EvtlMGHtwQh53i3X8yZVojXD+JGOwHZuKNl6+lv9+ahfmw9JXqz7D4R/S7FAH
tNMAmp7ecdYmkomeBD5oEH1nzUPDYpveVpA5JK8kTp+y6fOt4ZYNUAWDprS+e8kM
k9x7IY70aa+RkBH6U7KvEM1q1yZV/tcMpvzjF894u9AMvC+QYfnTgevj6waBNRfZ
niQ8VRfqNmd1mgaz7jTShscEHMB0ThyMajZ6zy4jBjF4OJkMvZfwhQYF1FINuWyd
/TOHH+Usqi4f2hilbOfgTZSluYUoqnigAESRuFj8fo/W25xch+lXPdThy4ZPi4B6
fC0YHOEU7szTey0Q9niDd7CLvv+pAaQqlxb1wp74Mn1BS1ht/6GGiMmA1BFFrpqA
+JtWj8cWPrYj/oysnK0Y1MqZpDt1a4pNWCrcq5yILB3BmX98eCfcmY6CD+2IEMDw
KNTUpT8w72Pfp3aCtmE7+6Wl5FghCWbfCUVVriP4UspdtYCLS9FeEya56cgfpREy
+TOYlma62QgDGwv7qYhRLSLcK58Go5jbejaR0hvyUfAcXUje+bUSzsBwJ420QjPL
X0JrHueMS/6HTgIkoeH4rSA+so2M+Okg448yGuEaRZrTOmu6LueQKIdVk3nmiM6F
gbGp3m00fSSolMnuY34T0YM1cbDT0Cka+KsjilbdF3Vk7YIUJK5gBgcrqQP2523X
1Nd5maLSP2Qg4mipGRYJ02gMJXURv1IsGkex6K+8aasrcoO2c3bAVppIsONBMn5J
mW6ll7Jg5tK8r/E3ABxe6H0KZY6VULl3hiesSrHBHCU6i+Eb6KkPzQT8hx6OxhVK
yUId0HVzHdPQ8OOeCNpfa5R/PAitnSs6tZbdYDcL+TfvnZ0HBSmCJVJgNG/rE7Ri
nuFxGCryhphM+uFXPqtnGMNGd3/YTC4boRQ+msX5HTa4PtjxjDHJKCMifIdyD+01
7sZsnOsJgYRUvfkC3Eemv15UtP4x4rqRAWOXNEzBVoVS3RvjIA9N4h2QZqSGrtYd
ekGCdUbWSA81HYcD2WQ+qzito6uxd2RYiZCtXOLhRGuk+qVRdelCjxbBXoUbt0Ll
CLrc4PnO0kMQgHcdQhbEOEYmmb0PK7Z8NlaN7rwjOZHIQXjEtvRPR/Ny1UtBmWwv
v/KANI6hlK09o9v4NaAONDpQyG7Os86Vmn2d6DxFz1KPnwQ7H6zdZ1c/o0FJUmb6
hv/4lAViW4qyqaQ6HPWPccbTIBBktgWciI71S74Ml0SNOLzU+MMU7NoC5oo0sKYr
Zn6gzFgaHhI9yXZsCxXGs8/3vadWzK/n7aGQBgoHyw1ckN8XRGUOauy3Gv6/Kwyx
2pmO8zSmE0L9l+6+GxdDosK1xcrjCABLwGo/LXgglgPCrxX41e8qkUbZ8Y/ohkrH
IRNyh+iQ37v3wpFM3/hp5++tVIuO2sJ+oM9jfIMQzroQFTfe5Go90ywwNRTrVT/L
YscVOvUgzPkz8ykdAmT8EbTdcBuwSyiMwUK0fSfEfraa/uzzEty5xlFY1wohswNN
a842QNI/QCzBlGoTXCAlviZwc5Q0zaHrvOkDtDANnjBwmGYESlwDoF6gkd+YSyP6
/hBSmX19VxFUBCgS/hQTnmdRY+l7Prdnz1zELislrwxsOkJ7xE9IyNqawFZwMZ8p
tZdJpWnZxzj36tXJ5Cz1YOyza+Oc7Cw5TJsAM/AJttg/7cKS8t7nXQXMK1y3q1Mz
5fIs58i2l/2j/lJTx5yD63NQOHQKKpHVYn9qjzi0TJahj+DmHp/cFgmwyPoDE5d1
QnSJIem6jqdFXeKeGZ4t8sbprDvuSclc+ICyTq1g6tVEbfxQY1DpVHKRt/Lm0Nn/
W7VUOTSv3oBu7oPyJ2izhs9n7Lt1KjQhqUOzTiqU6igHjBEO+B5QXT1YASBckKnI
1QHgpWHSHM78aWKee/xkxs5szHsGT9eZ8FbuO+pQIowneIZQNs3+rDW8nfXkIKV7
sipH+W7VoqBBIqt3q9JIsYKCyGrNgxEcNFCA3pUBsVElpDkw9HOsLZ+kyuJDag6b
Sw2HNh0EGgX0sNE6HrjaP0mhohlNMoJGmcXtg9OTrOUPKsvsmNTQLtgvFZAadzqm
A3gKLWwuntHOJH/dCXogMJcl8FIul/iPimJChgojwKS3KxUcB5VM4Q8Ef9WFJxMh
rgjfa3tmsxttmpRCME3Wp6xSSIUKu/FuaUkobAiL3PB/PbCDtKcU3MP9Zx3ui7Tv
6fzFVmAa/YWHExXnKlaZBs3X99t+1ZKJ8hyYCBLFDG+XQ9RaprH5IVO5t4W6MvtU
kJAHbjHTM2ZELFhsKAFIOtWjvhijjxl2XOdTvbdamNH6MRFCQxUGq8AzKJTGMUUI
fW01SuwXZUAYheqQ1tpt6cpehR4hNEUNtDBZNPYwDBCGwslZ+ncFPoPd+7VrSSk5
3puLvC6HB+6dPYe8CHrIn5wEa+rCA3fWYgBgHTTSrAFWEbbgm13le04N12+aKj4p
XpYE7ENOS0U+BSojCYOhIQ62IQIqxvC5L9cgIKNbcY9oRSLApwc5hWJkc78G/Z0P
A/HFzizwVat+as8yJtCji8k3IQSNG6JJfTiVdgoNBc19C7CZzMEeJJyU3ZiZCCoZ
dJXXktos4uNJd09e9MIRlKuXdxg67mItSQnbF6gVTXTE70maqMMdBf2iI3Bh4E8Z
y3ZbL0upk9eBE5b+509/rEbAJRRxoDpkzI82q4+c+rjt8v47IEA9sgy4F1u08uE3
Q0apwri1AFn+A/rSqcAVnIz131GNEguWGV5dqLLs0oww6k4TasEqTnzOS4aCwXBe
3MdJrYt4MnrBiu70Ps4LZZn1/0kfrNT2ua+EHCaBoYKI0zW1xO2TqAZVkiFVemjP
2dkhsZWIEVkN97Y6DRlr0nHvkX0RuY5Ut4FL8AsxcpK3jwQFaK3NQI0WiX5Lmavb
XGQ3HrIEBdJvTXZ3CoEmCwDQekvSe2lL2CfRiF1tfr5JEVcx0hVcEX3WSzM5Rycr
R6AaufI3WkwyPcfSD2APvGMqCd/gBssNv7TUuh+3tZhCTHmMwjCeCMGHKpDhr6/B
tFZ7NaCVluzs3he1VYhEWjaqKLqxjRv4JFlMZnFL/sdvS608CqYlarzmNAqy509d
5AXnUdfi3ZvJFUlEl4hPBPRq8YVx63fwl04zSOyB5ysM+5vTW2p3eBlSgEyUvQwZ
Be6wHcpzEUyuxRt1ua2DdlEMuaLNfXdkhliskmLHokNqF+/dKnK90QIOSTodXO04
Kl9JReVRyd73o9B5j9Wm0hjU7pgzfRZXqV6LAlz33GjSqC8T+UUHjaK4tNDd0IKq
Xv6ZSEb0BlIPekt7uA3GduuNKY5yOP9GteUPKmIuYtbqiFXgHmJuMgUCG4zgBPwM
nJNmKZuvbU+vxEQ3Og00yuyNkYXfKIG4dGdiPqP5pxtIwo5CoxhE/bfmhtbOplaU
vcr8kVfnHcVWl/aKGCBDBLmItPT4P55ErA3zqARdwrSBf7k6FMUvyAPG7mJjfnJM
28K5ANRuO+Jy2YIvwcI4z2zl8gdz639+2qHMQ6a33jI9y0E/EOy9HgYzF4HPQ5/+
3vfhO3lyR3aIQ8gXddpREebsr5a1GUwm1lsTw8xaykimpg9bkb1l4DFKYgvM32na
wiVw5F4dPLxUCURUoOTBO8gIIETag/MnylEtkLtRyjUpTMoFGHKe22wVGrVnvEp9
Wkh9TZz86x9aTsI0/qgzY00ZtYW3XsVHDILeXsx9PydsNFa6lqbwL1M9Kfu9aUxi
M7gLS/04wRUgYfq/RctElrrRrzAFitxJoa8tmP7OoZSLn0spsibyF1mEL+h2PMKr
CO+A0b+PLCnpm5U9chhOGYcaVZJP+gfPVCFK0gvUQ70X+pb/rnZy0ZtbC5r55La1
ThOpucGzK3JUX3pE3TqCs9pZ/lo1/ojgQh50kYPf9q1loJKF8e784cuRABU7/65U
qV+T1tOiGvzxfkDo4VNsZeOx23Apq8WNVraPDVKChU4j7JCOGLydv36AZNKt0t6D
nFXlA+TEYzwoIPGjJPYbQoB2CHxFUh4sBlb+ngcvOTJnj2+Maib8ptNV/+AXCeaZ
4ok5XeooP4c4NFbTtHCXpHwsmPSHT+MZUjgBb7Aqezt+wKOZDfY/DuoWk5vVkHuU
2hqKqJ9gAWioSsdSJj7ouITZOR2gueTMNsxuxbIdefNNhAtxIJ5ySU4LWYyyVYLm
5xJZ5TJLfuyWnk4hpbCTThgmkOg1VLTxO4JHRswCJl/NfIJaR3lfqxytjxxi5pc5
9NC8MwD7bkTlKWeDdHk99/Ng4Lf/DX7i3WKPmGWYXClDQ68PGHr8yY3k9PCPy+4O
nqjHYTZK3REA8d3IpxJnQC7592pYz5XduMdQ7OqCy0DTt3qK8GKRC4H2MX7DRNPX
sjxMgIqbN1TISiC67LeY5ddfYQ/VlnYlGcQCbM5FqUqKvDcFe7zazBnTjbKNLLoL
RRzX8/hZClnA/ZFqWPUc9r00KtBPxh43N7RgIy/rEYQhXNPr0C0kK3B8IFcDPX5A
TL48IiEs3KQQmEgvTZzKTGR1Xa7gm+B4tM0ns+GfPXtSUlxBmIDahpBwdfxKbyRk
sEssKdxniqi9ebRB+AzIJTulIIYvO7jvJsBzChBa8kQ/huGNDWvAV8AgtUsRSJIW
e72kYJN0Zen/0UoLwtwAWnaBvLImbqCEo9s9c7EWWTmRh7iyOxzcCSY6fj37AVHf
DwZMsx8CGRLjZ2K729uSvF3o40RqldZn16LNYTlSmLTFNI6IEjUCXjtc0JAklnxl
U3PyGH523z/1tv9GnMOxv3m6SfebEq91m949dCYwDHLqJpTkXOozx8Ps18SkvBSG
00fRkzPZcuFg4hDIIOszzasmgMJpaqFUYUo8dVgSzJawR5aPxF/HGDc/LRA4jB6g
8pjLgWU1fPyusZGpEFh+vAT0YrzLkbI5SMhPdDZKuU3yEceZ+wR/NVJkbpROJkVA
GJd1xPD2OW7PxucHmix8ANR6UgtEE0kPqstlZCE9L6Av2Mq+U4GjSiJ3RDvMIM+4
8jL6NmwLoxIN55z7PUuUVXOv+qr/00QQmvOKl3qOlWoBIZY2tjVFB+XYS8vkOpEY
eG5SLAnR3FK+a7aEm+p2DkZhz3Qd3d9tFXofzGFwWCmIb79fRzj4grwAI8Ppl1lC
Q3vGnd3I92KzgaG6+kgicxeOP1OcQ702SjyY69mjdtdazZWniSITwAP9GlBcNd5W
9zGHRVqQ3v9VaGpAZG4LweiO67DaPuLWO2FAaEnOXUO5t1a5ToNt7MLZiMuyilcW
E9ju1PFY3JVEPxt7/dlyKnVZ83bAE9zOhry/Vtc71c8vB7WofjHl4bbfhoc2e1as
6p68Jv0eobiQ0Jj4pWyYzbqEnNUF4DEKPxDtQTpkBQHrpJ0wUb0Hj+c8hx4UiuU9
G1a8XhDHzuNBCY16vV7R42S1RHohnp/Lny/NOp1YAf22cqj9X7Xyj1qRWsJPnKYA
D6NPFDxlY9UyPGR587VprX0ECrPpHWW4iVJnibRTJwVizZBSHjZUlKuk2vj/2zlj
nmWnNYU1oRoEIaI6+FfKqkanZxn9++N6mm7y+i/2Hb70ywmkmD7K8VkGK+z9LNag
24/h7ej8v2qztj4XZ9gPQNt8tiIPY9Qn3Cn6NTVyQxau+HXO5g/api63puWdpBuO
33UdHpst9umNJhfwBoA8RQDZeoZZZOdX5wWMibkJBUj4giMmm2/dauOSHMiPXMhT
5YJRafvX7CnRKPGN5WyLdDDAbejl9v0dcJ+qeX48/YdA6OqJaMRmV4e0rW2lTwML
XpKy36eMZpuT5WYqe2hdtA6JqOOlCbmqTjD61IRH6wLyacxc6F55Kv6m/KsREne6
FrHno7hKmU7CNy/biwthvI5nD74S19zmZosEem4hijH0WrcNilpRS4bLiH0IdTi3
zLmpRZfk+URRpftxP6VFziutSAZgZrPBsfpywdw1iWSSf7pzTpYm0r/eWaJypXac
1614ifqhOC7A5WUxdxzOaOTTWYSG5PPEoXs/r0/ty5fk1A2tFEhvua8/D5o65ThD
fwYSQI+GVaXRyhhS8MnizoleQ5YFlySJ14TEr7e3q7qhF2Erwirb/aDFtd8V0EQS
j2Qv/+AXebxwIPL0l6AjPlBa3d+gUQUALnxHeOQKG93qd60P4zHbwgMLn/hXteCP
LkZw8BPfch/EzSshWRjZMVhAL68svb6pVTBRuERgPgbOCe1RpBHvPk87OrnXInQ4
LoWiLqZVywHB+/bW7wegzZ0WOaRgHJmXakbRa6sdBG15qe9hjc5v14gbiEQr+YMb
2e4UpHsUEXq+u0HmFQtzG7JAMb8YmUfa3jcph7+IteRwKKaxrQ7tr/RjKQmc+QDV
bTmznT62obdyBYm1itpRaf6B6AL8o8iTLclLau5YyQVbyY8CWYHgnPzkocYnBgxI
0r5SWLto+25w45hJcOmsp1JSzZyxYYMK3jcybN3ErNKN5v49kZVQ4w8I/Y9wcsaI
zBj4mwXKBSjAgE9/eVWnHsJKBg9QwUDxcWM/Rd2LQRlH8GGm3CX3FDCH65nR9zEv
OLpfxJcPdqLrbq7zFzegQFoB4SsTSh7eNSl7LNzJXN5lKfcNa2cO3hXNsz2bdFrQ
eHLHwUE9ZRzPQpBGo/Jk5VYFLWAjEgwbrdsrdY6De8BtmnF2TVWbRrCNGzQ54Fax
mhI7O5/EVsNN2JOL8vX45fg7kZ1p8YurOyYFiBvbXFv9Is49XV0UqRpLBgagrX8z
fDmniM3age1zLsZvecz4WE3r0rJDvLof9rY+7M3ZUs9ol6A6Pt8jKzexjTK4SMQH
UJHccfafoCUBm+x3xKwjwgHl4unWze4Cc89/QjjR8RvzsKrcLAFiTh2FXuQFMRky
NYeDfGh7BB9Utt6dZ6uddUU9fB2h3Jf+6Z0eNQRUQwjc7GAsU/9pLwbL/IaW4afl
brst6ZXB9TYB3XONbRgJd3jQb5W+aMjsxgSUuJKt/qTa8oQpc8F7Ljym1IbUnwY+
/KpT4G4ZQL31J6iXSrZhVTq5guDocOOjz30bBHXzhbmLwvHhSxwWE75quUX5I7CE
QmA+bt4Rt4LwoT0SX2G6+YDuQ5lJvV+iwc8HpdFRTewAyKh0oA8G/nGJYiIoYYPA
BYjkpHyZLH9OygcMRwwvSHFhJq5mHS6XDtfnp3S/BjPvt5czZVrrs9c0IThyKlcJ
wf/KsbtfXUjN5R5Ive+TF54Rmh6gRlhfdJLmWuAhwoXcPnx7CAORcwHWtvXUVZQi
CvlV9mGCpeIClPhGwHAyKSvXyS7qLOQJyK4RzWEvpDOrzDnptm9ymH2UYOyAkExb
Rf62jKTUGY7QjKoa+q3bGpkqaPcLw1faoJlLHK07OBBazsXoWbFMPwQ5AxYrCGoT
xQQQeqgfnSYoiG5pCOf+Se+LsJblfRQlcAdcgbaTsIonndc2p8GI2DVK5nhmgank
TKcNF/44ihyDt9T1RsycyWYgjpG8IzEBrA1xDY7jWsxcrMUFZ6Rd9bF0GHa0E+gv
Nf4M9cjMxqUks5TpXSveiXrr3w7ME/8ljF1JMVny2dMyZF3WWkPlXC7qjbvxcsVh
ebKes3wgwlOoG5LaQ0QvTOrkfkvFWjX8TsRG2um5D+jkqKsfrw8HMJ0aqYvRLPSr
ektojT3x1rBeaYRvZcgPIzB5DaW9UQVB4WXZ7EtP4z0HZ4Mk/CIMFOd4n8J6RpBF
Tsd/SYb0xRgjlU4TEzSJ7wrlB6y7CcXpSMvIEnSMRjnDVaOmb/SXsZ8yKMts6v+M
3L/1Pu+tRDL6Gfgb8tyDrUrfje/eP2WEZ6xdf4uYQRJvncVfIM1JFpqJCXKCCkrZ
GmKyDMLdlMlfmnvhk3VXf7yTkX6+FGdnb/koovcOnIZYTxiHnZkYiLtAKbWxgNz/
jKLfFHzdDBfSozSRLqKWKPUI/pEn8KgkEFyWivc717SlaJNrDJgopb4swVvDEvjw
wNszXIe2xouhjX/vYDIQduH9fJXAxp7DO6YQNXyNIfE2lsfX0AnHJm0MRqsI3Kxu
3RMAjUKs0zCtT0eYk4cSk3d7wuiNmFu9RDzSSfbMuu7M+Hb87XJn122PrHTpMm61
aSb/2kYr9T5zJ0lrzho46CxErVgk+ZaT4Vvltc7Qjxqq/hicgaAF4rvItYRl+Pv+
52tBZ/n/hRkYo/Pn+0z9wgilzXI+Ctf5yYQ9NmWlsTZCv9LZZN2FuKv3plkPIH9Z
dXYCyuTrqrb5h2IHtnPKBofR5OsqvH7mthDBaLdhxv/wbS8nZdnLKWFB236Fznwu
8GYroQnV93fpoW+ty7eyHzNTYDXvbtdX+ggvVTup7Em4gGBE9WqbXPdC9iCRhmmW
sZ6Gj0B8bzMuM6VcyYKcsp+ETuOdd6uCpsnApMW6czoNWGbvC8ONC6YkeTtlf9SM
B399Gi5E92FhQJ5SDh8EowK4+XMJnLBbQldqMkUgenQ8tzt+2/Au0uv1su8nM4hb
p+KpYb/SGyBgRxTLkxEjW2SDcveYk/VaadpsFe/isxOB8Eojjic3V/Sjn0up3uTC
4BKYIu+rliCotglcBkNnPeEXGL3gbH1jIaTcLsKoN29O/5UPDub7e76A0QZiCZue
j8QSb5pZIbzcHfizT3C0AXBLU5runr7WJiMVDrzXlRJj5mF6PqseZy1k1roX8DZp
z2BcroS6VFo2ah3sLsEl4aAqbC7hl6QSBcrWl83MXN5dQXOFEX7ubXj+m+EUdZl1
r7xYtP7YN1WU+0M9TTfTR79XcD852qLetxs2WFBPQatuvYrVPsq2xoewEs952gDj
IVslRMOfSToNE4SrwBSpXUCLFJd9kZoY0F/NGCO/3bupG9tgo5EDNniY/83DZ4Zq
NaHLnc4GESwNqDbRQi/f6pRHWwhhwt0Hh0YyDBtHXyM3YnSONXBikAjlBlqftI7O
7HoUYIZJVRNMqTWCExPE9cCYuwWEgq97MUPjqCEKKsC9lDmuiRZWS4Ww3C9M3LKN
12OvZe2n51TBCbZDapN3wY19RbOogVEp2uBH4MxRzPUpqSal8eH+1El57DwSv0QI
LcfbWbsq6AF7VUCFSYNpl8VABre8L00YIaBm1nOBCgxKSUgsaYhs5SEqfp7FDrVp
eyXOEDI2gpFauNHMDAqzGU3qAVG0XyPp9SKiq7rtUnukP3d5KFWtC/m0ARGzB2Zd
vMfOjDQqLVfEDUCF2Lk4RmkQUM9eFNC9U3Pj1qENnoJ6VaJ7jG0aMPpFx+VjY/Mf
canuaaSsn3v1pCY5HTVaBftjHRH3oidPgAbtpoa8I3JL6JftUk6puFg7fJ+EhdTx
NVGrzYVh9UOspamgatc785oTFW4qOLzPt7GOdGN3VVZOmMi6TT8V7Ih9tVDqIPe/
BQbhjxU0dA6zY6syqqMqO+mxT5NlRIDvhe3xX/D7iLA1BsCX6ocbiO3d2bCoEGBR
JtFbupK3TCZX3QDUzJ7/axqg952TFGq/nTXqeO8q37oIZ6qEAQtlqS7Mb0hiSrae
mGIZ3pRCEZydwEzmP+7FN8i9fxRmTDzginKWIR5krgrJN3M9RHc5KJuWKFYbT34n
lJw+0TZN0b2IddVhw9hIhgyviaaPa7TUYZsVPjIywjtlkmgyRNrKefDZh3Uy//9T
irC2GcF1AglqNRUslW12Y2ArO213kzcv2+qLyqmu1ZTl/AovHzVPGcmXRQVhsIcc
qSB8m3eI+0+0HPowQTfiS7RwTp3JfQ5JmRQ2FALlgvDS5s/RhkZ9xwRQ80Z34f7s
zMykkHb25zJxWJcGj0c5+2CRZOEPsJdScQ7VxaWVS/H2DQed7/TvyqavHHk1Tk4e
S3YuSqi+NgPK/lyJGWAMRqSM+gfF7MkuHf94Z2pL4khcdXfkR8IZZqGmfeXBU+zD
ynVvAibYXKNA8A7b4VeBAIH7inD9PHDADSsmPTN03/oNxF0TWp9EfxdPExwY0/FS
EsZtE1rlD3R5UoGQOmEEfIiW4ck4NZtrkv2ZDVXt/5PuSkXBBxIptyhIg+Dcq/hG
UxdMwZmg5tuOLoSZ17IcYBxgnX7FCKr18ghlyQlzyBayyoUmNbcI2NtJ1D3BBQgl
82W1nuW5sbUCmiR+OX0qVnFF4DyGFw98PM31/1py6u16o5eSV0PeDPnWOgzZ2I3r
zVlPeKHjvKvtm8R/DTWbFsvgEzQMJxrRwv4yMpInwRiSYDvIVcd/xTX56Fm7rXi4
YP+Mz1Fx71bafDpWcg1q31enPAYY6URWk7St70362Ts5+Uku3BJL+3vvgi7uo93I
1CzFwKkj6XDFoeLAI7XddqaYmPb0ILoxpypKImzBc24pUXIelaoY9bmu40OqGzf3
fKFKGzM33Kmaf1DQNgEfEXfIhAwHVVmbhGeSA+FHczvGVjcdEf7L/S2dYXCzBFbW
ppbj0Th18UCA2AGjJXeqv7VsMii/dYm/2IiG6ncbe+TGe2lzUfuI0ixd8XOhkQiM
pyDfiKVmt78CE+dA3wv+t6ZlXRnI1qhY73FHl6u+FqKL1/+7Dhi/R3Zp3/eRFB0p
Eb9k7/h3UzW2ZsUx+1S2e52DMgso/1VyHWxRdGIvs5bYg1DqqMpvDEviUbc99tnw
a+stO65GmjobrRtW92edtekVBwDTEiopqk0XOMfipxxk9qztH2vXvlm9E+gSTZ4H
e8F8C+mT31Cm7mW5csfV6EfLQwN4/pCoGYLhedM1uWkdF39C3+uOR4LWSwy8G+QT
+/yIDWRqJOL2cTMN3XRJoULIGuAv40d7iCQrml6Z9ThdSFYL6Hb7u5pO/FF5j/uE
OX5bwBO28cMLOb7nHSM0vbKOsgIxspC/ba/E4/csqetUv1TdXl3cDsGEtZy1S/tF
EdfZoSWkppKJiY9rAXLM60HwWH/ExS/N6fmdk9t9QtBf+rG4Dxbm3K4amPLc7MSN
riSqwbaBtn+ohPpusgGXXvrNSfNbp6Ox0n6QvXqoQX5tT3M6STa3oB2QQhQJzs01
67zgFfHaKRngz+k3+eSMMZNCaxf1EjJtC6JV8bB+UV0nzdvhytT97yIPG8TY7p8q
Ab/yGsHG0RLXM7Qn+LSra9U/QkS+07zsDE9U0Ji/LHm3i/vkYKdX8y7mU7zrEC6R
kBtG3p5YkCxiC+ppdFcLMESIeasSZ9nlvWwMr5bHN4h6vsImc5YUab62aI7+27iv
xq7jwH4qgRsJfVbCW+qCONXuF2fxIgbZCSKe1igPZLjBgWA+C4NsDzfbCm9etpRL
bui6az6wMgs5xRrCAoQ6cfkXPc70YdIGc3MGf+Br1TE4UNxBxt2JSgb47lmQf1ud
A8R7csZurGK9i0MQNjaiwhXZP4JPk6BmmXhYdBzuvREVA/UWF9Su8hxSM0JMjM/E
47FCBvhAmJd9IVi0HjvX9aPzXOoEAGPK1VPijaXjwVkPzHLbgnCrFkIU5CfG4WFH
feVSc3QvgEkDaknULbeMERVQGVwEPs+dJ8WggFw38Fu2WVQzndygWBgtPFgqI76Z
mu+Dl2rS+MEGPuBDJPnw1SopCQjy5I/34//ltayK3lily8xr+n6CQmaXBk82gIe+
VxWJ8CMb5YVp8a9aM9YhuSxpHYIuC8nwgCBEypjw/VDsPYlN5xAfSzD89VrB4xed
YIusF56mlqhbnBp6ZvPlOnj+tNiJIg9/C6+qauILpzgn7W2oeReIQ5UHwibt9Cnz
T2fFJxozhnVrkkOTcYqWW6IHRirn+49gPJVQsj2iRceQOMU3sW27QssP7NBy86Q/
ExqQHZIeArdD/KaRFwE0HbzBeKJ+A1Z81TaxClvlgQk6+pQJRCcFgPkiWYFqdMxI
FTtdJrRsAC21qRHooz1Q43l1Yl/R0vGrL4mJ2w74YVl8cJWeJBMHYdZFoQtz/4LQ
Vva1IGH7/HQaVcU4ynJaVl8CAhjhRpNW5t8w4xiqlf2grOIX+3oIRURqE4FM6cH1
w4gKSZmSzK1qEUwx4es6V+oHHh06F3L7xnhibhv7LRYfx3bzSFIBVBXAS1B8xdvh
vWr9tu5wSiq4kLmwAH21qc0+5m3r+WaeFvOFTH6GmISHnWduODIKq2VdopZ7RTLt
RPQAD+Zmp7Zgohcloc9LyiDrT6Hpx/zFm30OrWSSMfP9IpLgIopqssLKmS8YUkAp
VvPWsz5hA9nsFg7umbS+0LKw10zd/fw0BU7ip+ETwwaUYrUogWE9Xq0GWChDspjJ
+YfblemzsFTaqfWlZOsArc3+HdFE19wtJDlmZ/TD59OMvwm7eH+cEEUW4G4UeXQp
hvX81iVDjutBkaZ17sP8ibrwn3O9IvHMb45fyoruDck2/xXP56XNJCHPwnSNulaQ
p5qEvo+P135AKH2nZEXRl08RBshXjrNuhB18iZqpVZHdEikLLMPRSWMhx8dWgssR
kTAerYKPDpcav41UYQGveAoS5XiobX9IiReKP36hpHtq5f5WcxwnuEc/4TBfK5PI
OkdF7q4W2rNTXXBxYssvIAwgC/GS/dk1r7y43kJyZ2DSJADj7caAGcgwtF1LKFh4
+a0+DYJhzikEZ7T2cyr2UBhG8UWZOfFrTeo2rMlA3IisteozXrt9P/R9UKNky7JZ
JzfwHvTFCA/lVXoXLoOFEG3ddFOxznNRae5GVv/9haFYWKOpifiRpdf4K5uTdggw
0GnAuXfqenVNZGYTTFnO9udmB0cjfz3Pt9262KDPr2RAVvefsA9/Q2Th7yykEe6Z
ccl+l1GDSoTf+kalfRSF48jrCOkICYkwiTG8NOEgv+esXsMN1BBnEphy2xGUIWon
v3YVQrcdJT/NvWiZTROa/h6AeKB/i4HYwDNVgYKk0hTPViwsXZP63TnGgbLaTsCI
7U09ljJ9tqQUPgyfvJIJQJ9egpI+uxePmriPNH4NlwsenT4JByOi1ZGMdX84GDDD
XZBr16NtbFmHdP5F6fbccCM3KNVrAgnshMYpp1MRW3rE3JRTcEpJbk/Kwv88T96h
6wCF4WKrzIPYjJ9CHCIxqPYGs8qhezaAAlL+QMca21eZXcXHybXCNq4Ff54orZJG
LkbfhBuIbQ2rTyRZRHgXDY70zHaQNEiP+L6sJRVatjExOvDtRxlJcUP1kniJihnY
qxoEmEIYegfI4FTvQXbujiHcrWHdp3OkJ8QSGBC16+7bJG6Jz9Gaf9sRVBSC0V88
E9DAULGCz4T3XegBNM6GA0vtpFr4TyIDeG1L0kQOkrAxt/S1og9Lb97IpiGTXt7w
Paf82RjorcjkQC2kAN2xwxf7W7qtsHXsXBTCczfS9JtfH+YasTKfsWnCKJyPEoS8
HB25Dd+NcBNp25RgpvFFLw8XRFljPfuw8DjOxg+QvojmX0nhXWHRwCgek3uD9h0Z
ACmwAy9szaSwtKILcGA9hfSNRTuqjlPBaf5frWLuQey7fKq3sOTk5cXgMpYevUej
qqcslA2sXPyrhD5s9NKCd1kCDLBvsQQj0KKZvEO02bZHYP5nlAdI7A+6cTrrC7JA
UxGiZF/fetBckI81tXiwi5GB73WwPFlxogMI/J8B1v2YjI18+okTvoOfalk98vQb
zFBXeIxNQBB4EwVNh0FwMGfHZG2y2kqeUiowli7chDU+TYuGT/T2VPo+jiGTayLo
XFEvsDbhDYhwW59etVV4nKy8vFZIYbpjd8dAmGpUuWRPrQRXvaS3Dvr0hg9oVniF
sVfTeb2Ez51sT2YVfK2YGSo5uOpd0sX19+O3+P9C5d4d5Gv+GMOpJ9Ahhty/prNm
OAF/SvmJrZ72AwcZWUHeUmZhqkUGmexrc4KhITAWAWCw0nOZrKqwMdWfS/avMdQs
O3FDy69UeCu4P0T5632W//H6tCIgk3V6/8/fP9PScpScyGZhaufmop893mdIKf4t
/pF3P0upozrrRtCL7kuqyIaD6UXqmmRKTnKb1FhHPpQhjU1iV1tKzHevH2x41E9Z
9fTOVbNOtTKM5wTeXDkBkZFtkbEP15INv/s7UvZ5udZfuSTxr3jr9wOaiDg0d5/I
u3X7AFXkWcvblC85OZUTo+3ppGp8TxTOgfpu2JU8jV2QLYiawlrv2WeyvxMfo7Y0
IoGBT7BXoeIK5o6KIPF4SRSziyeJZ3nOFzxRWJeTTUKfSJucvBIWHZOdidpPhoX0
viQBGeMs6bbx7nQ//6coQu8D5IxKmrNCwZEKlfCEBNSfQrz9OefRt9bkTJuGP6Xj
0RP8SbiX8tBrHFBgLBLyMMDTITb8seQJWhcilH+IbvjBzRuu1p7yDblB/K4Y49kc
ie1UKDOTlQsSBXlknQx70eiFWMQV+08nlVaZ7eNVOwZWSXB5AzQ+8b0wZ3ll3u5a
RT2dame18BIO7glD1n0W2pILVI92yAWJkio+w/8JgUrC17pG5cL5gN323xVL17Nq
OWqlSBgAU8zhNgXghPCNydpescLzKXUnOz2Hmf5jEJhfbpN0HHqyMBK/JlpRUh4v
eCdgZWQIwW0iKfJe8NsuaKfGl7q2jDtOmh7Zc5D6VO22BvGJJDEGsAo5Tg/SegUU
kHAZQz9Dsmt+gglEs1Oi720v6TLqkJoB8JStTGW6dttN6rv+D6pWq1wioFCOO/mL
9kN9iWGoWd4+mLJColwxtXWzQuVE0SzH6hjgx+du2oRD+VAvDimSvSk9dyNfVPmA
u5xvpjRwDuBYj/VjqyT6UTbv+sRuenAGJCb001kBQg697Bbcy9Y61Nc+6lBN0D2v
+bz0TDSyc8eVMY1yTzzHQ5O3FgStDKVfHDJX8ApdDc2NDnTJ/Wc7v25mDMOO7mgl
ZHkYVcSAS/6uiQ2avgILjjoVHsl4gIDmd44Gb4ogLe6ToMo899FHoann9OyWwumY
TIULCyizq2vNfEPa4Q8Ox4xaYvuGVkBCFsa5ZBxIA8N5CVW1oLaG2HrPf3OkAGil
8iFB37pk3IKtKhXreeq7Itf32xDNX0w9d2Uu7pFd9FoXxRPLPMqq/zhqU9k4FP5r
MgLeJQGg3dgh7ZmAG/vjAtJ0iVtVOnUwzpSeMBhsWKoa2lelsDYq7KllEmlTr+4+
JsksK3vzHhFoTAYZm+tkZHQ2M2+q2gZUkf3ADfvhpyn5A0CbNabrAxJGJq3D4Q45
lZp1YfV1ut0JJnlnkGpyuayhGN2+jqiMyTeBHP8llOthOj5hPzcJTQc+CWuwr68d
bLFqRKSdpOhzT3iixGeqZ1L6U1g7bknSw0q9i0MXCeKlTOIzgHBOsSzb6FKNAs/m
dZdkjcZn5GsbfYkmWyuYyyQyMJk0kTvh9e3Wn6O22+oRy10f0tAr8sy7i40CLAvo
SxFTVQFP3NbJ+JneA0etmGwgJeOfdHrvLgQDpd5Xsdya3koe7nSupk1vz33DBmep
XYdgncF++55XJ33Bbylh5gubTakEsyI2c7fTrufGe5R8NxIQdRucaok7xu786UCP
IPiGbUVXKMhmHHw++LF5vKr+RH9NEKBn8LbmAjYhRh9xBZPjk1+YXHcSIYzfMKgz
eVsDRb7yG13KgwDNbRTxQLkTZsFh0uuGOdYZtvD/kuIxwNOuEfZJDmXgsU3cwMq+
p7vPWHuj+Htmc52TLL/xrjRih7+HsLulnHhSaO4GTABVdxaex5MBROFVlHSfAKhu
ZT4uSfykhKwMryms5esDSc5SP7+OfjmoKFMaUPo+er5B5/0tIUOnZqGTZR7r2ILo
0azAU0z+remVS7VDqcbLyPcUIDI+RNEA/JNppr5ie61sFeCvm1GKWLopu4a9dlHu
Fow0tA6Y622mRLz3bCYk1vKQfyK2fkmw90MFcoFKW07t77f1pLgepBA5ITmYnX9L
X1XYCJihAmN8JrFY9oc92U8UnP8sIiCRq0PfYpQlY+TuqOgzmgMYx/usigPItreh
A78gj8BD0tOtp/LfUan9XKHrRFyLpDJbzaFfd9BbEW59G2c8+AG7Ua8nWideLF9+
QwLnLGPxamCwV+82TczJICNLoHlDFOruf92YDSYaP6ixa0Hx5YW+m3ktEJ+TCvbU
UPGcUo3A+zpjrvVxNxIVa29xHjkkijXHF2+RqrsTYQvdlAuo1ymxFijjFi4u+DAQ
XyqKa+splGcYlXKVio5WFmjoRTz/z75sse1t4nDK+LfmRgGTTvoW13sD4Em9T0Nh
CIOIXczOxbbqGTwISXa0w8T82cTWWgZQVxmko+BeKDLaoA5mUtbiWzZVDUHG6U9y
BAJtXjDbeOIBlTqIvFqRBEiv8+HTSkAmXS84FdqPl1zAQpauf0le4ZssfNoOlnUv
9w9c7eGy9H+xpffKA31TcJp1uvgAALltlSC4zVRc+YD332x84Rqu7cvnFzu5B8/X
fh9cqnnt8QO9UeECSPulwFulZR/eVdcFuYPuYnufxe7O0+EkAgIjpqLshmyukPxm
6UkMPjHwXJWHo62A3s++P0wLes36VXKrwS37czZoNctxhQA147F6SvaHXJBQ9RuP
zZ5ES+4Vu5qT/dWnR7DmvX1EHIF7m1YdiP6PvisfSngf3lMUXWvPjPMxF3/jDK2i
9V+jGs1njf66rHw9sXTBwkO5Iw9qLZSZ8/T1vojwwehwlLSqNkg8S5IX7RckQz5i
rzwTqk0zekTcNj77ZHb1WwUYRZpo7h7m3hsk+pQJS7gsy66Lgj3CGzlvNhzcskWz
JGK7r3+U0hm4Jko+7tkLej2Kf1iV2h0Cl834geZ8CTLT6XQTaIUyqIgHRRUPGi6B
/l3ZHdjRPrBm0YpsPAvIHR1UoXo9pAMzsKg7FYvGmPFhI9RY1TzqPuvPJBknzZyY
cNwf+NOcRtvQysEgfJQDzhX2qafILRsJJCvFxHQHNzB2yA4PrCuNfCskpf25APvx
saAw8Dmhv5htRinJUGLgSoXIHIqnZ2WGiExUQOFPxu6R9xSYD7eEbCLfjf9MwQXN
1AIW9AIt5MwEePB5OHgvQvX0L55Y8bmgnVnLtY6E6j260OYVwc6lCiXlFJYwTJrb
S7ZdMvIuXlr54KeC/cLJrz4fhAg5KGhpWHFoCamhMUiFCpxbrXObZPE6rRqM3ftM
j/nvHMX0l5CCJ4rieZU4LYqAAH9KA+XSTcGcIsVR2VvPgW+O1ksTEdX0BJ8wcKCI
VnEdjCoLoCjKDGSQunqHMwx4Cm2J2ARCY4fREVTlL5rSASJ5S75V9w5HnToDJwL+
709Nfs0z5Gi9fdVBeGoSw4BXRYMSnzMWGimQi8MgMgkLGT8DNNPbsuUlP0gcR/bq
DXnSDWGtprLCZItMZeM8dE0Ni90PqFXUkpIHWWFmUirkckc49PLH5DPemyHAP6pb
GjioNFWjFu5BlVjH+KuxOuhjtMprH97OCoYjo+oXgq4aUxEPdrKg8O8r02jIB/tK
hQOGZ/J5IlhNVJJc+6UX4E7qxmAto3wvBt7yES5dbNwaXYLGnpxZwpeIxbGkw5Zk
f6SpOef0Tloj5P23uyGo3MaZzyS+CEhryUaHzGbQgKm28M5e0T+EivJ5P6L3mvBu
ta1aAwziRH0ra3bbDsGOkLbrxtXpuaa9bWbYwfHzk5LqXjkkTYgWAAraZpa6Ut5k
j++gMYoSZ/o0G0FyAllEYD4yuZ+Lkhismb2zmGgloZsD6K9y0cNoYIIBNNETLliX
G1oelXokt+1ay4FFjKEtqGX6L0nD5YaUboEa43xl2UWI/uVcrabwd9vCuK57Xso1
n/sqTJR5R1KKkqcooGixTgvu8xI2w8Lg4RXsE0CEVsvMaeg23GFkQjyXHu5Kh8f7
hG1uKIbttQypWxfxsqd0ocet1Uw3KbmxvnN39mnt1dqzzvWB/dvpfBt01skN3kHh
Onx2dBhLYpq+kw8/IRv7tMIgbRQMAaskbmk6LgcTQQam4ahMf3yuekctsQDl3bUU
Puz6fYz+ohUlC6TXJU86GmieVc6B4pmgZdfthm5pcWe2anR7n/HWtq8z2YpnsYMa
1wFw6UmKTlA1HzPgPL1u10VONX09AzHEDxvJlGhmAb9p9KHWJ+JPHU31uWSMVG6L
0lq29SsxtyPQyfqGjChNKVu7EJBnFJK08myenV6Xa6VpHx3zfvKRJgvFl+jDHola
uJz7JqZ/WVR5jxDJAvcGeaxQ4ZUjt/M3MfCFy1/gIpcFXLg11yCilFM9TCGOKdM+
9h1v7m5msmuOKaTHWHvLNT+Kfk2j6QMTNWSgVMm2e3ELfqfrWmuGWocefq3DGIt5
jkiBaLnWJaNgIsbVqD6AEkZ10o0wOwGoWmehPeF+3WPmgCkfD0jrkrWwJpPgBwM5
wdV14ysutwk02Db3LdDLIsdDxnvftNS39Qg34AZ1znjlv8Y8ygfPrtaDSxCVz2l/
50gpHi2d7AO3tN/HLqc1L1PAF7hzzpMQODLEx+tmlbBl5ZTZJdujEpqoJQdLp6Hl
xDDMks+K0/NMPv4hrx9K4OdYA+I83ChF1zDzGoQnZUMjgMOWu0/wylGKBkhGYU4Q
yT98pEsz1ImFZRy4LukgjI3HzpauKy3sciQp4jEUOy4LUXa9MS/DGJWP1RawxGzm
Hjq88vN4AVS/I56hxXhHdSKd2fg2hYDCwM9k+2bU2PSRgzb5stgUl3coCJ+RbxWq
8o0BqMsrZ5VXot5gXRSTWf1y3ZqYZK179tHTREfeF03240i6N5h9MsMLXiprg1zC
726zo2vnq8UyyTqylnw0oqlMkcFzQVXakgANnr6QujEHlCFmDRXfRDjfXz3CNaAk
BtfUtsF9jRlvg6VXW1ThflYSqN0Uitlv/XWlGFGrOitkm+bfYqqky5ys2Tw9k9M+
VCzAx+nOZaljeeTLwuPQ/tI8eJYOj1h/t3ThGxvu3Rvio5oj+q7fJCAYfaP98k0C
zEA2Wc0EuGXSiSq8BdDLH3zOxcj6JM56ATSfHQaY/6do3jjbdlE3ygm2SAw1wsXh
eNdMiWz/lMEG9cDzu6IsqqfScnr6ATXSI+IUmccu6DgMTfN71iwgmu+RLA8WyrV2
TvGheponRamBZ0qUsQfdoRGj6S/CzO0BXw1YrZJgw+1en3OHGSNKBqxKAyIRNon7
UUA8jB/FReOHb4V8UAH89AowhXEzN2tvmaU4i9nwM6dFdeVNSApcGGB00VsjfXD8
5rWTMvK+HS1AtbSS1KfCkZFagrq1W09yn6B78duGVuVz3pTpMDGnWoDmHSpcov3M
Mibg3mciO4UWdgwNov/lItbvPfYvmbffrNQr07UDZlNd0bTIzHHzQ9BdBdKi+UwS
7orwP6XiNiaMj5JZqHjT/AMd02WvQZXN9Pe9MoB/Vv9rj8pCJGr5UTBR53Q8bpca
0Xgb6N+ZVEyyFDFWFGYmRFN0iDQTfRpSVc0EzcIGBJKe7WRGnS5pY7ErPSEpipzu
cLtK5E9m2ozcgdoVSNSxFVERy+g8S4eetvPRg1Gsq+pbE+uEGmVL48NkZvkBa1Y8
7SvQLk7K3LL9O+ql1z2WSLQiCulvVxQaRJv3YUHIzefmo1A6kEzRBuja0AUutGZz
hQm37RdpyGjjihLpxMqgXJV1N7D3dWlfvjLYbW3HbwpMHCupPljk6x+R6hpzxHU8
SUEDFoLHi89kBLvrjuZWGBrZQAAkymIeQnKMPFb51mxZCAm0gHw4SLXKyxYO8H4y
c/IkfvkWCNh+lAdcfNc7zVDqtVutI+ZPTQa5xjqpN0l7uYtyyTLsWCyB8VW237PI
k06nf1KLuri3/Wx3a4MQnpwukt90Fv6eNZOZiBarCG7nrFTzR81v8c4R77FOPRIG
/pGqC+lesuYpoywaRhKp1l5y0UEjaVk0g5fLhJqM5c5jTpSian82qjUHeNpPKHq1
fO1OeCXEZbwzfmeSoZ/2FfenVseX/P4eCgnATZTYNdvFjZb5v85YPljmjUAmwUip
oxBicPc1BK14G7dIaq1h2vAyi76V3h+ZsOCd9mYHKONClmG28ajfyyQLw4QUebBi
DyqR037r+kkobleaDr3DBocOSLKh6uwKiHBztWetIgxbHXyt2Cs5ForXCz/mtUlD
ZzY8CGdMs+21bX6fNLb45KTn5/Yiig1/oGhO41ykt6yoGqCsBpOAiekJrWYMtvhq
/i490Fvxf3NQ1trUdIeuXgPbUPnXYbz+omeRAIktbov0nUNcaLFACK840SfZ5Lrl
u2PXz7ajTklde8yfuZThXle9pMYqerL7z3Bbx5TqfRw+iHOr4+R3BOn+jh/Y84Q9
rO+rwUnqDaFAMNgSUwohC5ECzJFag50+chq/1IeEzcxTrUOEqkQkjU6dkcCTZXv7
guh/KmFC7pZGG+qvAG5Qb51KDUA01/YdKJGcLrpchtpIkD34p3pNhQKNPFEfP2/N
9d5CqWUvyHsK/+hYbHWs+muleU7Mp+AdLmg5MNvsZpBbNAwpsHxotTDFLXSbfCGI
CBofbZGn/kcFKiqU55bgn5vMIqvX4BOgbk2uYOLn766xt4Esx0MLxAJlu88kbWjO
0sqqKjnQlCqdvUIN+Wvz2L57mJ2pI5NH0EUIEDCwTItEBuh9M8GH7+yWl6ku7xyc
Oj7YGe8fyHj2O6IJ8yZKxb7lLxQSfX5LhKvC/k4KeBYpAOc17WfaujfGG4CY5+4g
EnCGLS2q7X5118BZcuH56F+oS2ksrlXE5f0RJ3bovtERY0Z/xbweiYtBbQXMJunL
vnN0C0NcvU5bz8gujI9NG8qyFmwQdfW8T6IJU/Q/L28F4Qr78ijk1eLEDtU1OtC+
CZ1OebEAL5o3cB3mWgrqzec2g35zWxLfFlU0ySyLYICeUVdmH0dkFRjEaFNHbQnB
ZAs/b0vI9gdJhPlUQaQ5ofpuiNPrXmo+h0LZ5KJwl/kZ1W4tFoxSW4HwZV8W7v9l
VPyTDPPrfdXH/LtB7C6yl2tqykv88wJFr7w+cfk14cgLn+oaB+LGMzHvTdV05bDk
bjX6GJ5GWhxuYcY4XpZscP9fKYBykbO7DcpfgW3x5ezqUxE2qx6ctbQW3uyBAG7C
lgwMwTMtecAA+7eEOaodePTs+ddK8aMS/aOTkcnIDbb7Q4YHoh9AqL8vJitWjP+8
kChhPWSn3euwQYftbagteGOf89RLzOXrBF0awe1CR/IeLJfcx213ewdqKax/hRf5
LEznE71WzlTNC7H5Uim2ncawtLriadpbEBsvpwO/IvrV/BdbOCzHkmr7RrZ3FzoW
2qsEAyAG1p6GuQSGXKqcKpyIQQ9WWVKf2VcF8Z3uuSOoIj0//hbghRo44MwxDVdx
7YCFMPXupZJw5RVxmg4XG35jb4CwRzP8jFuMKGn9d+6q9ZIzdsi10v+1BV4L++n0
D44M9uUeHleF8dWl3RnXFEngVUHL3Jggq/zVpYEpxVfAiRNfj9rChgit/nc0r+jX
/xjSfz1Szki3Q5aRcsuzsr85VQhBYVHOlwOm9KHrEDFGI/OFTkrGgb/LNXBrMhXV
mc7LbLl3nmqVRxUhr22LPyRsUjTocrL1wYbWY9hAiLRt6/o0I7w1gy4FnWT+kTjn
rceb1Y1TC20pAXWuON7mK51CioCqlxnVfY8ZCHM6sG0cC4HK+DK9bORzZXH7bMaw
zcogcEYukYBBoObC2Ride0DYpEmU4F5dSSQeuauN9QMLyR9tLnso+YPMS4l3Q1cR
A7V5oQNBPTXMN38ZeuwLulmGwuvJCW/NXsWjKjTJQFR33YzCpQcHIIAS2yRpWfV0
GC7evSnI0HJssqXG8TIljiigUuh3ZmeKaYjNa9lNg9F1JfMXtGk2YH6815Tur40O
ZPmjjNZvO/7uc2NBeGjgr6p1uKQLgwAQFC7AlOsKQza8Bzx45mIIWPJaVTxRYwun
07UrpT2AZ2eYa+azMcX0jvnrqVYhYhxho5gWn1aQwsxdkemEwSsD0dVqhjg8X0JE
A/G/z2zrYfnSk9lO6l+PV2Vf4ofppIyEKjCS4F/2JBXIkwyUquOTA6yO0RdC3yLo
/X8+Z3oaX7IDSHcStDZRpNiRSuVEVXqdhC+k8t14Xfa5RvUKStRhRm18tIXG9V5o
jWpfJOD2cSJ3ml0ly9b+5WAyOE0EKXCVHr17VE1SaSfKHdh4vInmpQagMN+19OpG
OfNapncEMGjEzIqD/4O2PgI1TJe/3ur4a2oXr1xi2VX3SQLTPe2RpJohaS5OzLwy
3YjyHr6EJ8ryS2tfNqKGAW9Mp7Zg+qaJFeyIwdkH9YQe24dRcbu2dyG8tG7oNcm/
K/4E8k+99m9C9GveXN6/aJ6yg+fxQlQqUnnju2AZY+mmJ59vmGGvfyZlk3M1zgb2
TbqrsUbM5y+H5b0XyZn5GKYDmSF3WBwYFsOtFpqVNbRmh3zInWn+SD1l2mm+8xz5
3POSQZIM+GXHn6F7EHIMYsF4wPj+TXJnYI46Rx4nXEXrDEB9kdEyv1IvM3kzgJni
WNCA3LxEDqQShHxQX34F8tj3jX0Jbl/0vg5LW74w4qRfpAjcIq0s4OL9OTGwFrbk
S+wM9GUqp9mCCOCFo79tGmXumByWIwaowId+FSPm8BKYLbrdtUaEyFILf86HoEyr
ydOR3e6RRVnrGy5LKdHuO+Lnw9LIcVkpQ70a5C1wVXkDV4mHRW1Gark8u/CtXCWE
3AyoHOYCVdKHZBwuV6SWlOYlHz4rl7LnZr6m8KrpZw7+84XP/T8RpHqYULbrKV8p
f1ylXCdxBb9yxudYjNlUiIPrr5AO4Z9+L5XPE0zY+qPsJvHb3+2OmulXrjDnPJ5H
SpiQVZELVmina9wtq6MmFWFhJ/NltPZyAml1vaG23X2MvfVEBFRrm4Asbq9qEATN
VKJRNy55xKF8IlMJg6BcdJ4U+rScEErszbqn9oDDxo1kdrElsuHYHrxt/eSQkTvN
CPusOqZ7Tk2nGSu4RbaCcZhwMtEeJbdYCfzxa9HI6GtMGK9BD/klNxjg9zQTnEVb
XiY6QrWQLBVEl3sFeMH1belXujxroI3K8HLAfs9t6PkETYX6/DXSYZcVez1YlPqb
LsqlAeZ/J0r7RnDFfOFyCuRBKOACRTs75t4LqJ346AZ3TFJ8X3ByvpzbxNBISHT+
iwYPEQGjiVOGu0FlC1+olD1yXzaZxNf1sAno4zPVfku9HgCX+odl96EnnpBSfj7P
EuTWqAfieErq2QXDgH7BqXqg1y4ek2aprEMQZYIsfxEUAnoPWt8UGvnmFN3awiOM
0EZtP3aLo4IoBqLrCnj61yxRhYjfp6w5av60N4A2q/z4X9/IEqBmlOSk3GqTamdn
/oVROj9kfjh7UeJDCNINLvyJWNwtapq9D4k3MaTwI8RL5v0rgvTA25YUmJw/O0Qw
JLlw5CAp3Rm2saF6Pdvh78tI5lJ8WXZR7OnUw/7PWZq65NwmFMsG8AKM0KJcBVAL
kGiY2x2cM8PIybJls+WUUnq01dNKVGdfUv9D+hfsCHUJI2l8M2btLQ6jd2FiTrot
OpkzY00eQIpfYqaOri1i+VDZGGq33z/AN8PfoPqjQ5tKMR5PNpJpoXzTofs5tt7J
J4vZ3IbjIEBm/a06t5x5i/nlSW26nD42De45R0PjA5y1ql1EbklfriECQSHj04TF
g4A8DQz6UlqDTdXmWc34QtCMMTRcgz+lMhGNG0zjTrJl1n4UV/SsLH783hwFarur
5JggkRw1XJbsiI8RtM9RYZA8LAWx7c/sJCAlcAGr1Zif88tDKpjhF37T5QN3Ww7v
EcuLK3vlvYfuRAhl4lNBcrMf/JACFzzC6nz1VBgoVsHyVJCuhh/51PJzuZ6260tl
5Oe+bA9TYOPGnZuiZZzpZ1WL4kZaJoKizC2aBMu+vnnHf77gNwaJTFmZ4Y+1tlEZ
3xxYdJ3juxzMCXs7aUDOMgTyLfFU7t55kHgiWbDu4SL8MDgyqX3vq4+LoQG2jzCi
87vSj/pPM6iaorr8ajCjF5d6bvTsSJLiVsBqvRKi9eAYaifLollql4vH4sFNrItS
TenI34vq836jicLo2a6ztMBdGIuNZbvm1Mk+2+t9oxNFBqJt7LqSZedgbso/GlFn
RxsTi+VCQKStbEAdip23QBSZuBoUUpritzm3MS7V/KIhoPv0k5KAZ7OnhKWbEg4c
ivxoy5WNlwflf63eKg7T2P/VClKY5vBVjkqQgpGwy0KZXwyYQtFA5wAqAzP1GcnX
l20uHntsoXPnYggV17vsuffvoOAm50gecTufrgVzd2VoThHJ9pnSQAqE0k+fccKH
TQ3bzbzcYJgjiSKFwrold6D0hkmx7ClIyKKaj68UfkdHSxkhqJroOilMnBTObCxc
ArSBbgfeuFi0rYDQ5qatptwLqCgHPfLKrLupaicAd/2ewcap1FL4ISzOypWlqisz
AGjCnz95K9AkAMlYWqZuieRadc2szFfLv90fPFHE3xaMW+2b9rGaykkhtHkmb/Tq
o88wRkKK4E4bV/Xf/TZip4i+7avsEjX1l8uVB10uKQHruuWsrrXaIWzDYBDPOqtM
jvtLgAU5RLnFPBArFd11/Xnh3oSzLMHuYTJglwC3KyDNnV7YonNFJuEcAEZj5Z5p
8kVFgTEd2RuL8c8kA7y4CUOpHWJfHeHylLIFges7oWlH/UwZxoAUOkNG84k3W29R
jmo3Y2jBhSckfLLsqnmwLnArvGBWzJFzyyIepFUzYviZv79bMV1jaVV1QrATMXSz
RSURHkC4+bDFhC8dtoaGCMa0HiMYYL/Z5LE0bzdEdeebsCnOJGAIY4W/oy8QcNgz
PEgE0EXwXPP0k1CopZC0U2EaodYNbZ9LXSV+/69s8PjYoPu8KInOINIPFyiE9Ern
+7C0/eev5vUUiw2KvGELFQH4Mj9vzHAtpzkc/eWvXxRFR89O1M3mZQSYLqtVJ2Ky
vgttriGbeI3j9EaZNx6idVtStZCCcOj/ZhHN5JI6EYuBfLfDOM2Uwa0IPRLoKhMf
gCa1e2ErmYi5c2mAouN+yL7clpt5aNxxYLCubUTL8BKvJ4u1v2kakFBIg38s4xGj
mib9clhwFbGF7Rpss8OlNLziijRsD26QBG7GtMkRLSkZK1Ithh9shYTlwEjla18s
eFBFP9xemptarmPNLQG7BnitLgnx3NILWO9mOgrx+0/+ynwks7ciplvLypaE4lRf
JSzgBsfDvTWtYC8YUnadVYALBmT+avx/b3txS53tQTbG+mcPVS+At5wVbShGrXbh
ZxbI+W+QmhjscKUmD+1JOkYF5f6PZKPlF2jEh+HXkPlVaQJNaXXlTzgPn9ZSilQX
n8z/yOPPhnA5e+TJR48k67bmC+TF5l+NP2B51mJfszoglVO/fA/C9FjoXPli5KlC
BAzEH7ZqXCETmk6/F23DG/Ak6dOOdi8SReWD3duByavvg9At6unzDKy0oncStALy
/+z7aMzgXZBO3UMgodlJRP3JPqTbq4An55ll5Jc0/do6h6zyJ4jYl5HDDJmNzikL
azcPksMMoAhJNfxY9W58jVuEll61EvClW3avKDDCFaadNguj6ysjIniBXXyipNR1
fkAMYWlzRJcX/W8YxIQL1mcis2UaZE2PXSKmPM+jLkWXxAae0THLVTTmh2ouCAYL
oxxmknQFHZhZjz38Wjs8clzpSyNq0+llWjj9Gi5DHnE8OylvgPjAsQmIijqyxwbW
WZ6G7beDSl6cf3Qc9XhaSEY+g0xYkDkFrl5rbv84yPBy/o1WwlkF154if+xQuEUS
QEyKUIBEq3LxaU27Z4UlYIXCy/3xgw719go0PRacsQj3roGKmYBI7QI6LLtGPZBW
L1wrdCA37w8/pL4CWb4rjtN8yVb0UxAj1wbHJbhA5x3pI5SYEgNethBHGORr+GWY
o2olf3UHT+h9QfTFtiZ+NQt/ZVoYzuu9jXZXfDzLC5j1peaSeMz89Ytm7hlyZUDi
mufMtQG2mXI41hZuG+Hp/8Hw/EnT2BYXIyYuQYSl89CobMy9zjwZ1AmJ40CNSj1w
8plOIwawcdjcphQG8A50SmhV/1CyumxCUzvuJraetRXQoW4AVdNQn8Bagb6MOMvq
+oDAhVB76Tt6N2daNt/9Dc9J6NGZgjPEgv17gGe4UQUTHitkMSPpctE7W3f2tbXQ
nlE7CXNwTSZ0PtDIHl2JxiKpvJb9L3ovin6LItmp8r0WHm0gKka9RcSlVOHFajks
eEgJLE11FDEmFj1dgtiS8858Db8FsR76+revljwSr4RDkDOwzs83wXMcXa+mR+yR
InAJIOx/HugGabPhgCEKcxi9L+8K1gf0Kuf/QTs+btSuef0wHJcqxyfWs0KfwsxN
7ZO7QLGY/7lhHvaWagTMXtz5NdRAS/RPX/dzvcqEEmN/xege3hX/L6Y7/zaKvbF6
geRGkYwHHFXqEr36Lebj+ZHiYka/M2z0OMVt+fP+GxH1XBFtoFeNg4rZjYCIKjG/
MEPbQbCFkUwyCeGWy/MULN3oPuPJ1IIKZ+rWg7vUlxdtvihQUsxhtMl5yD2tJu8N
lYfqKiQM39r7LDlkw3B+8ojkMfbegjRoqYPO6Ji8EMRVpd0t9rnHV9prKPt1t68z
RV0/XjBnhY8/MJ+TEDNgfPX4EgrmflLCHb60iw/P/yDBwvL/4glubn0SN2jeFXqZ
CK7qj5+oJi5U5E33cToh3x2xtkHsqoKOI4MkYET5EuWBRczyyP0nwqXLAN9mAyR7
X1iUuCjFya0Y0T8yREbPxJs5f65eKz5dAQFXpGXrG8h8QC3q7XaBTVgiQQwsEGJY
Drghbd0PW1GgOMy18B8KxCz2U3E1oFaZ9Ec4MbtvhescOXsUQWNJcmDBfaHApj3O
oCbkVzfyOssWaCMJqzMG71ycQhKRLb1ew+LJO1bK9ePoOp1L8VH93z5ityDlU8Rl
ZonNq2+EJ832qpIi7Ixz2RlXB0kHuY4xbXsJdq3FHakAAVZ+MzK47ZdsdxHczswl
0Wt4cCe4MYnUm4VOzKLlS1AibB4jw5u8AHsgCVObdB5aLuDfvIFvnQWvEHevzRVT
eyD1dGO/vkn1T7nNVT0GNefRC7y6B4J8q/sjJhTXv3YEKde0fwIhGxGSbeGsrmGW
7EFhyMRKsxFoa0Ds6q4AUGYrX5DHiL4Y4kGeVZGgUwl5cCYgQCTNkhzCJXA5tZGs
lmbIxH57hlAsx+IAn0BMw25Jm5SPyDQs7bC42GvCk8YMOIz45lgnU5PcE9XJ6mt4
4g2YVvc6tA0L7N3KwQvVQvBz5wExuQO03t+ln/MOhu6MJf9fsqAke/+VWAeMpRkM
2B+p7nagbVhNzpoOdS9yVUQin7Brb1AUOGBj5eiGvXE0YXVipYwvJthQw10SmaIY
82YLa6FtS139ERloKas+fsnJeVyrn+RyzGzmT8teF4t9vMFcR35XrQtxurj3Bs7s
PvkpFfM5/aeC1XO5xbT2kj27Le+1q28QnEn8BZA/iRWsR4fdeO+3XaAovssewLby
Iywot9tmBDHfpWaoBd9kTR61RYz3r9+VPBZdJD60BB52YjgZR/Yso7ukl4Pb2uU5
D6s5LdSLXZtJlWTuJCSi+rWVipxHcWgSViHWgEMLRd/mrgWQJnjq+gP0SYgOeGu2
wZ9/MELlXxQZIezgJWVcHXoTkdpeH97inhBfEn3OMFCtQ8Sbvmf7BtE3UoI3ZacC
gcYHJXeTIWGc/4n5Kg3Ul4rGQKSe0+u0Q4CCEueIa90564nYd/qJGGTRHUuYycvF
E05tlLz56Pe5F45wgco4EmPcC39jhYhlYlZNlQrOzbJPc9PkCYRGngtuKWzNAJQP
0iRqq17jdNeqvvMK8Vl+hrCVxHsdJGNbNOyBF+0xLWeVGJvAmouPZ+Pumjd8ukxB
9nJNYd/CkJz2AUgLjSeY7gurUw6Bxns2AFxfSnYi3SJZFOPkbOpHvmK8ECzBgMXF
AV48nv6H0bB2cO+XWHMyxBCtCyrZqvCDNrMvemhYnPST5Hrsk3L9ecVr+MvHmQ+u
9levdwUt3N3QW8bOIGQ9o0Zcxa6DTAoCGwezRujVbesC+TffiLlcjwey/WUojQKe
IRUenm/reekQUo5joFKJT/rVCIetz9OZOzALgYaFQetAnUtSZE5YP4j6H08ZzIDG
FkjLHF9up8VXPQXubwK8uaszAztQvLm+l4vXCJcSQZhxRG/iR10S7sY3Ux2WFHMQ
e4pzoclkF8qr3QITcVE/PM1Xey1kNgxNYswqvgCyBZXWzYOKErC7nYVaREU6dX3L
FeTQPwKbVM2v71PZBOwFHp2mO3Vh+5nQLX62GbzmTX7cXzySyp/JrrqwfyV06psn
Eq3sn1AXukHvBkmohenKyhEND45ZnNHHinXcKTfrhZt0yWk3esoBsT8WLCto/k0n
gFnT05GwdSXW14Y8bwkGvJ8httWrH2zd6ZmLy5HyOX9/B4x8mRRpNnkc8gLk42tO
/MJC3H6yXtaAbIfh6M8RsDwHxR4EgdiFSDU/H1jhyd2cy9WTr+ihv3yvp4Qej1V0
d1sDY2Xmj6UkC7+n1kOMPJg36zrerwjB51UbFUA1Zh2xJA/NNh8dy1tENNbWKraK
clxj8iySK/lMXlYBa0GDhvGG6jka2P0Z8XL4JFINgr+zV4cEJeaLkpToyGcZl5nb
xe2gzao4GsHhNMomELsB6jIgP/iaHu0w1gnfexTLCRJvOf7mA1oUzyyPSsINdwtY
7UTNRSfUU+cC2U0q7P0reWVz6w2h7/T4+B251pNSeh/a53VlZF6yMmN1aowyooqe
BxCCEgugiqzuaZSvWG1LkY7fm4EdhMNWbnDUMQ5QRtKu0GMydVInwXrPZS6Lu7aQ
KfkGmlpsBMrakky9sPM6CpLOq5srvVxOCvl8akG9zO4WeSXeJ5Rb8/lcEN8bvLU5
1AQWsIk7Tl6g0IK6kElyq0hjh5kDnN96Ywdeq9w50hAmWVUcZ1D9SWti2q1AEINC
ymHJbgjf2hgKg1+6DbhDsW1x66YeGGFsplWtowzjkvhLmEuMo0FFx+R9NCYZd/4A
R/nI/X+AYBqGZP2DnsheG/9gQpCBc0jEFl3Ib3w3bY7fyhKRbfkbbQlEOBFR6FFc
G1bok78xDg1iehOKMVx9nCNtPK/s5CZi5halm8xq5IseIAi+1y2v/FC4wtCt4Mux
C/Ktr/Iz7OWwQCHEX+zt49EdUhiOqMXChwP5qaWNYZ4W89aMmtNv12r1iyElLFTM
83584KtGGUSc6B3fJ3MN/EJ+SMJIIUAA6Waht+4WifmDILe1TXEqhkbzHxA2xWiq
ZtnqTxfu+RyxC6a78JtbCnFk4/YW9zUZYAI9kdxD3xsL+1wDaijKd0V1OzUirkoP
IhpBZqZNK49J9kau8X6FZJffoTm5C4IBhKVSmw9AKewwddiioLoVKS9g1OMt/IZ9
j+ocNWb99BvNX9iKmsjD/NdKQuxRLEb5Y12gZLwhDYe30Obv1QvF5P8ZHMaISq8Q
Eppu9LKBwQiWgDjxh7TNa2UZXOHPAq+ZX7GI4R5msbBiw9nfBa8O/MDNJeC8d/gL
+ggLPY5WjA/bx/tbgs02pzJM0DNZtYTS0QlMlFp3RqK6mQmm696mxYr4C+0Cpi4a
7ekVYOKFcDqAvfXV79yCG7T+Gyl05nBWQ3Ql9TNITgmktDEoTqZy5sSN+M3jXqoU
JzfCz27F0RRVCuwXTlhGuRkfQR4tsVejrt96iEHo4NL242nkrrcICTPhzKEir8wZ
4f09LpYsrWSA9Kv/mHm9noYLQ5zMuvEnmW41xSZ33lqk+QX6jBgPNuvw4OFtV1yr
6PXVVjUqPPegXYgnij66ygJwQWOK4C8etGAJSv02coeDDEQRYEtEF02AqwgImCQS
5M0Cw33GeB5vLIedvsJTlUxSfPbr4c6fD8UD94qnWDtPCmDu0D0SvOFpSwj52zDc
F7rvxaA1bEcIDcF3PqY8tuGXHU17xZDsUCADE+5FDHcw2YMRFg/zaQAxZugfgpCP
2KNP+UvcUnI+c0He7i4vFfSPV+f3FSRrW9S7sQFUoGdtx8+bZLY/PPVD0tKZqgJh
vbIIgSmKij9ZIow/vR9O+nw+5PZfweL3Nv3xEZVEnExyj4MrtkgGyPvrqLZAO9M3
xHD47JxocgZEQgAXXXF7vbMhlmrQg3DpTw2s0LidjoOp4p4aeIKFnNnq4YQSq0LG
QLkvKdDnBenTtCWt7furQkxLX9auc80yb+3fX3x9s3XlgKsOR9SrAv4WrwdbL7+Z
+SWf90jt3ahtmcTri9WWoxVBrDNnnkhQr8Jlb4iwR4QBohEQH3/oVo9mTuekxlI3
jiHCD3ZMxTLEl2Kb3YmXLoi8vdru2ZlJ2pSfL5kHkQ/1kLB2RttlUfJN9OeZT/Va
q+IGNjgDjeG/HxK9XwrEML+6wSQlPHB/GVdAwWaxdSjd5Zc5tEJsx9Ytivk7g68K
a6UGUtMVp2tMDbHS+PdlogI9IQVgkJiwkInSi3oELFh/qUxrp1uobAsUYRpOYXZF
IgwRDJcebFhaDfEh8JycDlqaOZTnNf4ii7jyz++OumfaMmUEheRqU00BlzBFRPTd
VtaSaJ8PQ2nmkUqNb05CAxeC5h9bk0jfoYNzy6vFa4+S1rCWUbfv6LfrzBysLmKG
DS4XE2NW2FZZadB5/3g+iLviH5lj/z78gApTZtT8zmMBFHyJnp10cxvbJfRnX2Un
6le9Tv8HwW65pwN/g+40SMEwlBVUUGyi+R+5t1ip2Zli9C2ijrRRYxOW+qVPaffk
tAT5VDgCK9F95Z2Ac0BOXsbCg5tednPMX8Frat4OvCQwDPDfD8S32dBw9ydK2+ub
n/Ym2O5BMpnApUCw5Z/yDQteeRghPrkbNRELc2IQovIbQjf38ddzTfvOCuV0G2OH
qxd/7zWj/J+sT7d6mSEY1WTlNqnHAfMBzIDk/AOjJ/GZGDsathOhvpkb0cucMNJY
gIO98rTtz8/ufuczJ6xV942ozHEjTaevjxrYrbzeP5rR3UGAT97F/vyELByRwm0r
kUZOMdF0hfnU4+FAlZet4Jy4FOAjbEe+0f+8XrSxp8SbGY+fRpkWwfrtV4wUmXtY
axJhQGNw/S7a/6UtzAED3Mj5r7eiCm4Cg/7r0J9LT9rYnEBWVyMqdU+um7zEFg7m
lT0rkq3N+scWsJMCC6/xk9+Xq8YHZ3IfZXHv75/lyjU0YpFSHd/9853XZS/SIZpd
NcNfVeH4cGC65z6u2HMM8oR2rvQvczKZrDygAsL1LAAQQkzOjUA51EiNz4xfxdBH
3oAEpSZi7iYEzgcAvO2/PiBPajQVVqisFPSBiL1IxsXkgOMaA/AI0gTR1mNO9Nsi
5nwosJSbDiyIrFHOGq4lSJaV0it41ohaq1hiI+xYLi7FmwEuY0PR2ujcRKla0Sq0
gkPOZWHVfIiQAURzNOET+3HRe6DOwTjQ3f0ac+libszFmmy/kVGn7MSlounCMMwu
vwzYoCN5BK3QAlWIN5ULKENFfU2Lw7kzPx+l46w7u5y7IABXPldKOxMU8dwu616X
wOl0Tq8eVc1IJuQPBkjUX7S8ZJue/zmZWU4MnUH9lo+sCXv+h1xG/BWGHcH8wx/n
P5cXXvq+oF7vhAVSvZct7zdOODaTvOgzXUl6ca2XKTDki7iWWpWFZ7IUGI3DRCSD
ZzVIufrJw2O/PAdYVbMFFEMuBNoH/p2aXldsgd/bjlEcW6faLFUBlu9geSLohhFM
v1QNucGvP6iY5yo1qUMH4bhIt7s8Z4Ot2E91yZpp0iXVNwuLNByy9U8y/ewDaADl
QBFtCGko7DAtnEcbFOxZnaJIYN7aIAmL3NzQPkm74+AnLBcLuQaSjejntOZC13wp
l3UpXGeGdOg58RasQhjF39fe3VG0L+AoQOByzHIeUWML53a6Rt7yx0YTtwURKAux
yLXdRmjRC47aLMKfNy6ZRi7UyW3YDGCxAS7twBmDDV6RYIqEyXt/Ao2s9gvN72Ij
UCeU2NJe+GzMDj+zQea47d0ZC6MSY7KxNtf5c1ySwvcW43yYEYttWAeKOCvzZPH2
CcPo9i45v6lDNakqBm7SM0y+zDskp9ljoyOz1cFYH04lX1Z09XlDr8jk79wq2H5x
+l7DMDZguXunYyKEgFBSGvA7EOEnQuJSVyHmQsFqRad26MwyZuJRmHDv+0NcJbbt
cif3zD0zjs+rCi/I8nvtbXFeQdicMJxo+Zs71ZQNy4FTYHLIbXxZbbBGZxMLuy3b
/+Pve4Y4Q6r2Oh4MHGiH6K9V/Q+KgMrLaepTRTkRKqfNWQTBZiyeZCkvkP8TeZzH
9oeeiNYsIduszAi6RO6eD1vqLKsn554jDRD5DeU0HQyaJF26QXt7tCwfmyrZlngk
tZquhWxIpKC/mlWH/alMNhghrSjc9JzzFIrTJi4tVAWRJOEcZAidgJCy5uEid8I7
tKq7KW5VFrH2eg1W5nOk4PoW33btkYrOggsbJtQktUz+Jbc+thbkyhdNU/Qb5mjP
rud7WqlcE/FE89BLT3pM5XB7hfvC5Y+vfXLHEWkpA8tqF6JK4WE5JYimzdNW6Y8X
i4J1imepVeI2CFDslaRIxTllMktxdRc+8lxsol95SoV7f71k2Tfgri6abzmZNAQ3
twS6lejosvTyro5lgEo5rL3ZVSqpVKTwH77cGeEWRefwVwh5Ov6E3maSv21X7qCQ
5JvGROBN9sflC0ppLWy86/dKWwpRYH21HUCzMA+FvA9FS7HqlHeviFwFtNQECoyI
QwETrxOlvIuAhhalZSZo/j4V3BqVgG6c8QinQohX2Wa/qTJDd7xGBjvftLaEC6iT
P3GoF+y8gSURH+gMn5o4LFbZ8PPKvoY/g9LGariL2td/4N8GxKbJywYI6csQ+Tpb
7FKhjLpotqVBin5gtwM6RXfBXcc+PO32+TngeGwXoVV6L5xgLF4hJsgeyvw8SYZR
3gvEehs3OUUF1GvWd7sr9QhnYJ9o6g7mnhYJkrzqqXISMXTXWnYwk+O4+412dI7N
pPsq3s7JH82RxEseYxKVom+GMS8xgVsKPx0Yqn6uXSwemqumkHS1XleKamN8h1dZ
TeODe/QUoAUzi9oBpBpqJrWxuB/boM7itZp+Wrq1VOn2crdgu3mM/bhFmPNc3G8g
PB/gxCVOuSJtpyKpxmVDaErRNCZ+pEtQM+JtjcjJUPO5ndrU2AP5P9tENprQ7raP
4Qa6FiUFecNN+Vm1mcrZrnWjbisVMFE3GLHvxHllAsKCdIdxRSe2TeX64X2foajS
auWLnFcf/DYCTFnB7SI5PL0yiyExDqzquvdexhxDtqCva6R4ndCZIGQ/hSpl6pQe
geCPOtCkmuVY3NtIqPRVQ6Hm37TSBCKOJNxebCcOtrBHzIGVKxbFIJmTq5RS3c0q
6i413sziXqkdKWc7Jxc2IUgo03+MzL8CUhrtm6WQV6/tS4xuU4TSbQIh89x77Gmn
sZGY+SEZrvOLihiHj8Twxj8SbhpCjHz/QbsbTe4uQ5caq+UruqL6gnkD6VG8Q0lr
3g0LSUldwH8ewci1xqP13ntUh0gpccBJCQajcGV0NyEwmb9XB48KW9DqPtCfX0oG
+S2tYzmUBl1B30/HvlFp0znEphduVD9zsZtMwW3T4i2KouKkECV8gDSkHMDjrcod
4B+M29ApJwDvB7iKee7KJrq0BuLHJB/IrTnhiT3QiFAIrNmAf4KN+a9VSLlsNO+1
eM8hMH7OGUpusWxsXJGZImEt10Olk3Ado+QUJoU5jPl2dgV37uueHPRP8Ii5xLTP
YpO3cf84RqoItUyYcVrZrtfFAPyJr1cw32p3HzVtXKQJ79TT7sI7RSEJVVTgPoPp
PpJeq6tADh5vhhvemPTyX9uo/tX7MVQjqYY/4lzcyw3YqIuBMtICYaA4GisO2lwp
sOdBgU/lT9STmFwoh6g4WN9+QDiJPDgHe64WZR/zm6j61HuwSMIvCycXKaBkY+L7
cDGvQebL07wNvAMjb8LIL0eHL/FjAxpyK371c4t0d55w92tOOBnwc8UGi/aOT3bB
Hg3fZ2R7YChfw2YIvzMesfxC6+87Uutzf2qCmE9VVSRzLx7LpVxKtC+0Keei2Mwh
b8Gm3G9QagJENqVZh2pJeGkDMCKF4eMpeS7QBBdDG/oVuJey3C4VqF9xqWrjuIn6
ec9CGGk/vx474R6eUOWUtUZYWn5umbVFK1z+uEHCvWsPAM2BeNEZr53BP3HryR7t
XH3HocPadXz5DyfPG44MuMI+rJO/rPdnxe+yxbMGNsTOqOuv4ahbtkiOqAXRTBCJ
1Rx189l268vnwt57AHGx4oc26/38jv/qfJDUk6Y0ThBKBmvT0J48sKwUbge/GPvZ
K3Vi8ExJnu1NB+gmEbft390L8p/49Hi1aqB2CBYvK4DtZifixnILiBZh7mNghEqO
T+/bvp2ZOcrtsVdBlhr8Wq9YCMIRGSafmtpkeujyUfkZnAWMX3jPKQupItgrG8ba
kQgBqBW7wswTQzUL3e9CwSSrW4ymx7+VTFnOpgTry8SvCTmOBK4uDyUsiWgXS6F6
5LjNuySdCv0q2X8W4lcueOM9IrDr/PZlwMQo42bufKqE+6LSP6LmU6Z5P0CQDkS4
qR9ScSPx/1ZNtx+jCGOfXmrX3MNGfEx8Bw9/HpppXm70OIWzvpnBkhl4Ibg/xkYa
JbmcxoXxoaFlrZxs7GXxCFeRVX6Dg8loM+smPUiPfZHCa784oceB+k0Torkr15Bt
ihfiwjpcRRbNbmtrrUJSLIcmOmmPgRmOoHEOsfQ5Sqmt4ePODmZSK7qE8b2p2rbn
uY0gqJDpY8bWt6pdgfD2RIhLlLkrihSg80vIGHETyU88A0+v3qAzBm9RTviD95ux
fVp0L7rbFvHHWKefTWes3osZjBbLQSw1Cer7dBHJi+osAVtK8m99wGw0NUlIqqVr
96jUEgtS6FpcO0B6rPbnWNmgRGy4MhXQTyLP96kymLVh+6n9h+jjwalJYzrVx6Q4
sN+JNzDiROXo579efRz9iZ/Q5Z/hUy8yLWsgvGcK4n6IwvN49Y1hz/QELCy9XyKU
cEVen6w+xS1WasxwPBeDXlfg5+RKlsZy9NzanVzlTwd94tMOP2pzTBo5BihMzYsp
C7h2fYouMIp9Jl0+IAlTdTX7dbl/SFoMGoCb7NaKd2m8rDUKVJDw66lZvFQUdNt+
g3YK4ugATHZxJZLptgLQL6j03NvpX+IReSp+O2aDRqZv6lhkI7PAYEO5bVTERql6
BSZKBN7N+rlLDIVMhCDnClTH8jjLtHp1fD0gwkxZ/FX4dEboE/g/kMchW2qKhAlT
mTJPoo1qqSuqLLGg8bks21bOg7eEY6wYv2PnStAfwQO6wyyWoBHFty/IgpWvzoW6
biKK2xIDIkjrY8+t5QQt/SgpmS9Gfc3bVWZso2lLZtQyvmHFdcuMAIB4ySLgzwdQ
+IWdBZqm1lfAQVSR+VvM3wHvSNTBpmXtJ7MLTUcxHglwhyhH7oP+bdP+gvCe14QK
G03Lm64mOhAYhcFkHukWAh1wIaDbzgRMeumW61V+QHXj2rWk7CLy1+hAFdRCpzlH
FRn2WpUCigs2ig3rffxdB0rxe0zyr/Sm/grcQpKMYiSzhGVAS+DDJmfDcspotOfD
Ou90sVglG2RHIb6pm9t0Yq5vH/XbwVgKUFTu+9iRChiHhZpMI19JlXgJCFiNBhRy
i3QV+T/4bZyeN0OEThNRrwwlAh5/ShBqoQysiv4oMSSBiFYNJJw33Lnxl3Q4WgOL
bttcHB8rkr8XsFws10F7eebo3U0ga74hqc2NxL38C+7IenapP3RfWAh2ARZPcH/r
lz903EBbC4jRgKBe4aRz0gchqPYjPLGtlt7wfhptMweZIDqdKgL//i7aG0fz9av2
/310b63R72qPWK2xOIq8rbR9An+OVgMjOklXaIZXZ9dsuNSBCGJmr3Wcm0kk4gG4
pA7rbO4/oCrhf+weOarct+f7Zy5xr2Nb/5S/xJotlbV+DmwcNP9ZlPoygwep3h/W
gZRdtRLn66PAzS8dRkECAat5MAGPR0z8LJ7X0muBcQjKkH4x59oZuyTb/9XQKUcZ
`protect END_PROTECTED
