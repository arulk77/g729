`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4ywnhUpJAl9LoJ8pmRX3Rsag7Bfek+QRDonlC/wg2905
cY58j1PYdFUCmNXMItUxQFYsK0D4dAVJpz9vSKgELitC9dbayyNlRX5PLsfAaEU1
4VR1Lfu/Z0lodtdT+EfAaOnOPukMGMTmIJFxzesKtQawUpz/mBul487kYAyLBuAI
6icIzs2pmUftf5u4K0vlRHPEdM17xHhwo7KAvGercBNr5l7WMt2YlY4l134Fg1JV
7D0RWncNLfnXHxNy9y/+wmJOegUbGaBDAkZwWMgNuyK19zR2ypUdNBkeVNGhR3Ww
rsIEMm6DRLKqFrshhX5D7NzBFFCjkqm6OSMofqtEKv2q+AZ7dCduXfIT36YORMcY
T/lqPYzjb90LNXNOwbr+Hg==
`protect END_PROTECTED
