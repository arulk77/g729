`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL83E4tVlEFHzYgzrk7bgVOOzkS/2heu3QyiE+3PwolF3a
tvKnGAsAnTMh7siLoTW3m/RxHtLbur+UCXosVOAjURNn9zlwCCHhLYT4VuA4qYQ7
DVh9ooEaDfFoAysbVevG1Ieo4QdNnoCpVWyaVZxDODNI04f2dWN5KiQzexG4pQ4I
BVUBLvBEvQD4hwuIzO5H5QzFHcRaP134X9nyHER/VayAVGXWXeZAK+gY3yj8PYCp
Ir3qd19avZKQQ8fdgbSeWmlAGkR/uEGjQtlivgnCX4wGqaYH5FXjqoN9uAdpbOer
Wygn2i8PDJoTAluM0pCs5hH1Pqswf7y06MIhED3lU6NHQsjwRSUQOYLxa0MqQs06
ppBQKLx5zbo+DIk5SXULbiQAucGjyTuRdHw/w103BwP6VfsCBH8L21BSoZKwi62K
1xJtI1IzVEcJSZvn7r7Sesq58dl1uYxq02iqZjg8oOKuHbgJUAih+giafPlHGsv3
`protect END_PROTECTED
