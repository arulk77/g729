`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45BKd3I+J00tLo8xXjvL1byjdVEYsF98hi0rc70WiLcQ
2Ko8GaQJNx82278ED2lqGK2r0QYRHEMr8xEWHwW90wvyFh6Q22DBogot9mpfqLwK
ymAqgm1UTwDozl+xKYFsngCn5JEsOy+I+tzB72IeEJwjQsd3XcIRArZQ7TYDfAzq
GvfeKgKTrkSdDa97DJDERD7Mqaq6TOVhyeYv7oAxcZJyelMm2UjjoWqerN/rZ1RG
ziXbAmMX6i0h9iiIA4skkCeMx640f2kzsjT/YPAZdI0=
`protect END_PROTECTED
