`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IVAQEutWJ+Rem04HAd7sbWG986Q7hbPaaqdH1WbVc4aiqgR/LkJXJ/fkh6H+4StG
lUysrsONPj8X6uaJSWdVpyX+He3dC7PkEx09tfyOTL4TidtSUysKuErCtuIukrgt
3xVs8iybAx+h4GZVH1AlAtDQCPPDbnydjnzK63w1RJlnqu7xT4e040wiXuGEVEmI
IWMFKiO/znTK9ujvVhL0VDJZJCTDquhdPiZlBXLfH7d/fAZ7qh35AfVq8gpkO0B+
hAiigUSohY6IgFwpvIs6EkvLt2Cny19f10Iry0jRZ+WlGRixDwRiLaTaNGaxM7s8
3FHFgfLrM3Tupnm0L+mmp8QplvvX8NDYC9TdS/lJTFng4t90AMMjZKbu7RzU9GyE
FE8H+6+6R9wT9Bz7Ww+wApdCxv684UbNZNAh7E45R96HdGf41psR3h8q1DrFplzO
EtmdOYUEdYmyIwIQuPP2haM5MFrcnBcr1/8DOr4qjg3Uf7oqxTRIriyV3IAnhKxE
yXnbDAcr5lL9tihs23x1OoBprSWIkIctb7Nov7+dJ9LXzXeBdiS6mgP6C0+S9NVe
IfiM8Bw6RQwxhzKXeFTi7wuecZyX0vXbBAaneCh1uJDXWhVCzrsTzvdSHWTRvTMu
KQ1vEAQzemuv2JcziWqaHQkT4IKkLAYsC9HeFy2q2Gx3xa1IQqVOyPPyKEtNh0H6
B2NWlegmP6ehJo3DTZECviqwa+p/Ap9qgPXbmgYeBW8cww9XyFBkepFnEV/ux/2+
4Uiw0LndbGy+0FaPrbP9V2/WYMPIOkQlMUTmWORkrsC2Gkfnfcxr3kUdiEY6p7Gl
ZudYFvp5eOJilUEMT7c0eZHrRfah0cgCr9a0J8xLJV8DXLWDRhxkBxfEEoS9+GAJ
TbnhFgJUhQug7waqeSLlkgRBWtOtbR/UJiybea4MSY6A9YncvwqmFfLedfcRmskR
InLmyOT2kHJDNeaJxqYnsMpGcQ8E4zYdirL9Lobq6Qqg3KytndNjm+AZW68mY3CR
0a7Wnv2Ip+INwsQf7EuPlYkrEMIIXnzb8Jn3yHZSsC110DIg3qJ7g7wPm8ZJZeIe
Hpq4LZD/METadkUOq1H/mELL6YFNOyf150Y3QKNbgNPMNds4McaCjWcRcES9gJya
dtheBEyKY0sVeeWsYzQWYMTX6gOlkSmNOYUjWZeGQkWCck0zS3JTuutD1TX0pZFr
ALjq//30AAL9xUm4mmYnOt4ilDqEKJY8mmcx9tOPW/p9W2PM7kR8MP7NKv7k5jNk
FmREQoHre2rKCMm8fHPAB/b0Jwz/H3LDfURr49CaeAyuwpD6yd2e2Y1jpPF8PQPi
MX1cCNk7i7QLkqNCJPVxHt4chlfQh7fI6SHUjNLjTghELDwElJbdkpsbhQY9dW6T
+wgjO1qReROFxiykM/VZ7I8HdJxchqr/9dxRTeHXTuviE5cJqx4IARr5gdX1WIG4
vtToz/YI9AmTg8gaPV/9pVUu9W1FaCekuWjWqVjwZ+z4Bzr2MV0D3AqOIbxTxOqZ
LLVOgzyzKsyw++2izvvuUwmpe1rN7XFZiNmj2cGXHrpfXP9ti9Cc2YMtmFfuHkUX
MYaAUFz3ZiJOaZ6ZO1bFkU+RDNVwy4wSNuDDyvZdE3/HFWW4V1sFqZrV+rdYttjJ
AOOabXFEBZ9zdu6ryAoCEjn44v2xCDfX8YtjY9NGL8SDJdS01DMs1RyzftEbHYB7
xrEaslwpTuNm9EaAYpmJTWa/lAaPCN+lhDKKdn2nljG9xnTm8ORMGORoqTKf3+hC
fitSR/auTMUB+mRds2D+t6xHlD5o/Oj7Myi2PyBUt3SygrKV7s2mJRt7u9wNPfB0
Rluj4OihhSGLUXFND4fSiYPo1UP1/5W3iAN/pWWBd+9754kek18BlxxTTIiq0Kpr
rM0xyrNH2AmObSuSAaMPhYShwrRlKhJVP7/vUQibPOBi7xKDVE8DMI0OJ9G5uqBu
tyXS6l9D/mNgm3dYdJsLGVyl4jr1vw0GRjPVucyUfy457OCMDg/MK3aTd+aFdaoO
RYKG6FagwJd0iNq8XPIn03iIE9FB3RAYTzGv+gy6RRVFwJZ2hYyed/In3jfr5DIx
LnEypNCrtKgqLKIQ8EEoP3iFVXdN1VHJQobq2TsyaAd0Dzn+IDePwBuLkTsqb3tX
j0aC116x89jZZUwMFtY8xPcu58R1Mi557JWKhU1KFZsNzVFn39QBP+bKMq6Nva0w
Nq2SMXVJ/dpOG6aL5eOPfNnndR15AIFukDOOmW8nGctfiQ3uqJxKXLx8ndmr7FSw
jsLJys63dUjTd/ocNYJH9u/ufx2E7dvZlPZHLO7KoUOBN/GBLCzddX9LSVsBtRr6
trUcq2zOOsyub0vq6QQkyoWl6AEynk39A+ztTekezEgl3KUP705TJ1jnkRAyxBHI
`protect END_PROTECTED
