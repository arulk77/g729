`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKCrE/P0GfnrejokTqWN1T5yThb+8fGfevfud0uHzSIA
8yYm2nRc7JaFt6DsNwEkMZoayDBnkMnp+LmzI3ERjNe5GwvLqRdOBeSlYQuHuA3h
3Q2n7BUyzQY43PoIGjNmO61QBNimqTf5CRviEJuv8qpVoC6T+P52V8Bhin6ojgVu
+ysCC6ssqa7gooRK3jGm+W4ee0/Wo61ptjhxoOAURmKmajMnBgHvd7qukvtibLz3
fyNP/ItOmVdPy+C2Ge73NGOk+HUBgjMsqBtYyCpYhEGtohXdUEs8OqH68uapSbU/
ZQfTdigBdAiuMPGXFaB9vyd2lyoDOJzu170+iXrqH0vPmDqJY6MILokanHLCrIIA
QbVq6Kll6JO5fKOEVTMRpcBLWs8oheyi8/ytbASx+oEoGJ2bvmSR63A0Nstq3zN9
I16egs1iR8j26L51ol1SBqWOlSXYCf75k1lRmiHjvVTxr5C1a1SiVxfaM+awR/d8
Ez/Is24vocyzlRdeTfg6GptnMqoY0iQSbLFKR+1ViLK0rkEnRBYzTOutJXjL5tGJ
NB1fQukHyp917g4SOQxnZVS/KMcaqqcGWwMhgejFtX6AaF9pFwpmOL3Y7PnoIm7l
sDmJlbbrO6D9wbV3Lus7vTL8aRf8IvfLZh/86gQ7EdBNHVHNEfzgndnqKuJsGe/E
/mdOmxFNFTkgRs3al0mHQrP5tOkE8e31tYLuUEjne97m/xHyocNQGKH1EnkaYwAI
xGYCC76WMblZS7NfL8UYZbJTQMFXikwaJOMzGyHcF63ejYpOkCdXyxdGG1oeK8uX
T92UHu7UP3LSqkgX3N+ItCnZiKOEYqGYdYTo2ptmhUf1oz8+btPqApEmguIFkwnk
5UmB13CVznLiFacLxqjrWXQ5dZ0zwuo/PD17nvgNipH3ssHqd+mjoniETP+aexSa
R/7BaIDhFsxSsPlxZXr/t4eVUHb5TdTjkIrLvD92tfRKdyOtCDTX18hJGgZPQ6x3
NhTa3pQAI8VFQK2+5vNM2Xfqhrkg09sUcyDCeR3+BdXEGagRJPRC1HNKY7B49Muj
N9q6KTYf97oeFDTTen44Fk8C5q43oF5PLw+HuXujY3FUbOoq6jZe/iUj8wTiwpGP
mNPPprOXpPJ5cu52M7486JtWFqyUCV4sFNoBhaeOrlrw8BUcN8OqjZ7bt8RIrnFg
qTaAJscZ+OouWZ35jnAYa8mZ4KX6CnL6s3dDCgjcwRWDsPEcNRf5+ctMcU/ceQ6X
wloNri/zytArnnJG3NEMcFyyLXR7+LFweD4jjBVRF5fg746PCGfAy5pkmrhRmmAv
FVE4K8vSIgcIebOUe2+XiEDB2tofwTvWhcbxbEhGMAeV6DtHaBvnNV/CP7ASQ5cF
znPzaQa6c1VRTeOrqppUFuTfewBZeJcGhHpjW9NSBAR/M6f3gocFbXSmlHfztpp5
5ZVLzaYCxW3f9HmwkWgrRRzZQxy3qE6PcIvI9afOS2TszDCMBgdnAHijjzTaTNbK
FwEvEda0xU6ZMsem731m7V5LamxT4bTRyC7QD7cXy9kmSiWR5l9VIR55TiT38edj
EAwn04wu3GZeLC9rMdcGeC0nWafQND5RgSEYarGx/rlUNOKCcsRF7Vx5NKCHxS2J
BbSrZ95hNyzxOaDWa7Ho959yCQows0rA7+NJYQjtZT+tNdRUg9VpI9AKOHlJfN+F
+IE+w7nxfNhtIH19HkvU2JZMYS1HIhMSxZVHYzUgufK7vFfz6Orpx5woorQ4nT15
nMKtfV/Ggyjroqxwu9g/1Fyv/8Av1P1ZJVuYSwYq+oUGcGpyuQau5in2XSks9rI/
YoQa8Nmra3qVJ0ExghlBzYbebYeBGfb4sSd5YUbjahHsvsYayZQOw9BPbTw62LhT
ib7FlmEMCR9hXypf66nD93HcTSoT/E/gdbnrF8kgbyUBWT7FSOKgPb3+1B9eeXnI
/osSI0BcGiYQSlU9nQ7iHV4sSSQcoDr/dUbAGmpI9kYzZWSv2QYOm3etV38omxSr
B4tLCcfe0mwesGIAhNEd38gkhzc+TyOTe/iAR9gnO8e8hTcQmPdMbvwiaJSWCpyI
se1BbOni5lvDfLw5VZ0XHmLASmf7MtCgeldxoOCDq/raSL6MffqlZMI8B4KFfsJw
XVysJAuiUNq4vK5MTkdAjb6xRgCgPazGbfZID4S6NDIRKGtsuSPLyfikePkqW+qV
PdlBV8MfwlqJF31GQgGDqPc7UlYD1LBK8nf7VdzC5otwSPJG67RKw+rzqiOu9HXM
Gr0TXxmXWvZRx9Kq1OD99+GySJeStF2IIQv/ulDobBKZ2q/9FlcnIPPy3V56K4tH
L/WBlm1c6Nh6qeU1mDgiHYHQGf1LCtYKHxijVKIv1zkrBYHZNzgX+ItUei1rIT9p
wd0hm6UxcaMyuu2t/z3usxExV38yskXOWXLtji3r4sOyGFJdI9i32OjdoJq9Zbbt
MoVzV8U5IdH1GIpP3nLqEHXl0iynnvXb7aWXnZYndDPv2jOmsa0GXY9YMqjbA2+h
OIhYRSixyeVowdpwKUEZoicTH1MEsjTMxsbGEN1ZZ4fNF/iyZ4qHJGHZiNu8ZOpp
ee6Kgejc+2L9c2pU0QW2JFgHU7NO0YmxcXGacUEIP4F6X7LjBwsALJglHLe3ylYy
WUJMjgdawd/89SAs8BG8kByS9eCpKgPoPEu8iGnuGGMpFDFySuLM9FTlzrZ6mPBA
932RBBds0rCZPF5E0CsuYfbDwRLO9ZPY4uZ4kS3MhZLAKDNOeaafFq3YF6fNCCs0
6YNmL1bgwfIXDM6MAJf4TmW5kl0WpNVRQGzNDTvi3sqzW6lZfIKZi4MJwcDC3XS6
ihQAzG/lvbk6jfCus/B98f1uJBMgAqHxpiNYufjGjNC1NYcxMgRdG61+BTwJ/2do
H2rzvEIVh3lbuV5K+nTDUfDOC7M+e3Ii7MtJkoFwPNEVjqFkU9eqhxp3qD79l7JP
78nWASjEI3Bx7sSqYyVi4Fqs9lJjOr6LYDxpAm2nnu4z1IfGM3tycmVNAYy5Viez
4wVBPbuGWJ8CUFCFYEqTTwDh+yNFnsZ7x1US0UqQGL8f/zcsppW2o9fBTbi+wltE
C3REaQ+UxCljUwhTOEBPxNcKCrdcvEuKuUin/2qkjwTNzxFPYrHr9hhyMnKGzClG
d1lKA0aiTljIt4PJEpr3hSgXaYCW/UxcK2uHPVCNBS+BtnrRPsnn9IsiedyHy5yi
2p0BlIXcHARUq2NV04MVtt/YyhA5+ndIGHFEsQTmD8o9+bhbuL2+Cmh5/ud714K4
jEm3/Yscz/wCZfkfKPaM92HVsW3WgCFbcD2cctGUPIXNDoIchChVqRy8bck8wj55
VCuqFlhpUxrUOQgYyDC9/yD0PJNegDYa1NwVfcQCaVPJoz0L+jcbQEStG9o6tpB+
v1W31egSovdpMxg7gvVyxWr5hKoVoEoGxOR5tdMnTj2QtTphrJIia/0wXj4hLpjN
Epo9lebhJMj45rW/bJYH/kEfyjEql75UO+aYzkS7hpX0aZd2b7UR2sTb4u23Yu8V
MufW4CgXnJXeZPzA24cu86xR/I/NBtx9uwCLo+6hlJrkOZEvzmfWWZQ2sS4TaF02
T8KoWKxFlfE4XeFHBqUNEgeUWFDAeOexOnD/CdPm3fnYhUXLb3Lv555TpMwFV+N5
Clp/yNfvRIyK9g4nY4Pzxpy4pld0wg9Qj/8b5UaGG7mmHZu06r1E2RQt0jDp7nmy
8w0qWuYq4UZTAZES4azW46nUhPbHxp9y1/iG2wAuSfpgIrIOCXpZC7ElhpRnPh5P
ePbM/kIvwAgPzl98I9MEGdsgBaOLlvW8Wa1ybgUAI/g=
`protect END_PROTECTED
