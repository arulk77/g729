`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
K9zYCpDtkaFUb4AJM8PDsA+xG8R55/LljkMRxZ0qvT+uTNI8iwgHbIBXgcQko4AQ
IPtMh/vkysa2R/zkPt/O2aU6kZYGMq4yzRbGLYUWH3HeEY0K1pgEyZh0nfG3mV7P
1Kgly+g25g+zYd+VmA0gT5tEIdzEfeMC7rmNhdy2jOXcNDaK7iW4N4cAmfFYzhjO
amHrCe2Tn1LlQTO+7vq+exGON3T/KXvL0DLjwijncejw6fXzwaeBPIGd81cK9Cb9
clQ+KNIQBNioUG7K/aHuGLjjVhOp7lRVTSCfmBQzI4ZGl7hYbT1QhA37J6y3AiUm
m8l71cvZKupBWsuRjc81mVE10tLKEhfC0+pxfxiHWmhfC4isVtrbVTid+ldoU+qB
DtU3sizXPSW5IB4m95mj5EeNxy4NB554ZfGp3qwSD+mhYD5bTBE95W33mhM7MpgA
xLQrZ9XBD3BOuucTdqHm4y3o3d6PKITIvVKFFIni51FKq8gysUC0vkul1CXKDz/T
WqOzrOLLGmPB5SH1tKkCgJc4foJgBldjt32osElwOa1kiMXDfVO8tnNHFYV+e/rQ
dNht6b6t6TRVIBbN3/rJhAWEDguBDIw5dtui5RNZyp2ouwtmOB3eP/pNszwmp+8U
7k5bkl34c2kM9bCWuRInZZFfo2fIu5VcteJF1/ZoFoRGHibi4Wt43iqr8QGHwUvs
`protect END_PROTECTED
