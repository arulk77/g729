`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCkrbF476OEpyobjQA90wDpFHLBS+Gk7DvytUanJaf+f
8dnF/IVQ8TNYciXGLZfyKhxOCaRuHMO7kxF1L0wYa3pHI8S9yc9g77GoN1jFRJAG
BQjJV5Iv0/A2l9LfqM51hiR9l3NfWPUqcibvwKiNUvCn+es5X/vxYKFPn5t4pRpS
icUkNdMC+0tk6yUuq3S2prz/nmMyxOR7uIw764uTUEcj3wWg+9J8SxpngfdZXq1S
AqPVXqrFXCwMeSPbiHiqazdc0gKHhGb2DjbgboRUmNHW4uzjhf5arjmcan+B/ouA
`protect END_PROTECTED
