`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCS/dLocTFJX3SknaMOj2bZEgRViXwxU6/gvm8hGS88g
APboh4QkUhb8xRe3k+JSKP6QxeD0egpXmNexYp6xdvj8+IdpN3tGaulxrzQjhL8I
PAbwK0NzyqXMKAxfo0KAw5goLKGN2RnMUOnXG5hxrxSH24Cy+bgAr4mSCiHgo9MS
`protect END_PROTECTED
