`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
11n63OtjxU/o+S4VrKJcaVZhh98cJHfGY1Vny8Efu6liWlKXGEx4I0LZCClhKN5t
nk76Z5ans1p4Q+XhgYNLbM4dopAf8diOq70YJm6BFhmon0ZWef8ePaAp6sRgEUY1
uhvFgl/Eut27WnTn+i9WbcaTVJSSmpiP0uLCvx3rbUFUlVA9SdedxNkOOVsvAnMV
QUc5rhpmc1ZVxDCujiDapPXrm17cZn75zMk7HdB1UsQkDWwNlmOUt0rf1vHlvDf8
sVOHF+Fk5YqgmSSSVieCdDxSmOxKr6Ce0a+gNp4mUxUcmlkJxUsTt0PJu68HUyPH
XbMJejhTUrPbyvn3JUVoDUBcxaT/dRfHmWUuXL3kQAo=
`protect END_PROTECTED
