`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF6kyTfsZe9tAd1LSQabye1MR8VKtvSw/l5AaATAlgo2
HgxWG6C8GySvEweVSMH2HNVLWbptB1bx7AlxoVVKLLWNHhRwvnQHd/AyNLcNtDat
uJnG2q1LTzYYqZEp6c76phf5NvSDp4rtnBmYii3VeRqBZPiistkjFnSYq+FnDpx7
S7QznjkmPjHWUsxOB3itnES6UIh7k2YUn0pU3MCJuEpXvzcFodqxh3YxJhfLK5PA
WGB3XMIQOmVI9IsTLgogH7Uo+Oiw0z9c90SFxDF90aIJrKlbzoO7ZjprC2putHlX
uWEzWCbQYEz3Cer7w/YPvHJvbrnRWeb1XcR8gBwm/Sw35XogWoskVEA9FawUlwoX
vSyA6668NUOHn1l+kbgsP4XeMWvh7MDOx9CMu53hay/6hx9TsJPf7A0CwRYQHmEh
SL2EqUYf5nr8X3udHNadDcFpBvn7bj90PwIyvQAXrhxbKJA6ylkMhj0mntgx7wT3
6G5JWtmuETQY+WI0UC+L62zZ2fhMjRsjge216BY9Mq1SqGT86tNWUmeuU6LFpTqG
pBseetAGdGLTGDogAkNrz69QqSieaI7Jr1w3GTeL8e/8dwzYITGHPdlVn67oQv2e
Lj3pjj6+fKdZ/9n19jqpHs4PbW5zFtg6idbwrksBhQMmV4nBlDdEqStfdkfUy1na
ok9AZbR5XZ8BQ7NGDF4Pk7sf6tzzZoJEx5oZwKdGokf9jeVwjQUk0JbNvns5LM4N
ViMIhecBgFVWa5+4qIHnqRA4G8X8r3prsHtDipD3+I8veoO0c/nHRvDCdvAbNTB4
wmFkMk+nmdQ0i52BCbUrF9SnLHHzsikA5aPOipzXD5FIdybFKYmvXchie1C0UFdN
c0yQgCi6mbe+UUDUcD1VLzIPyhnqsbyADhGcQEma5hcuDQRZAB1x4bw4JWw9sBVA
UIeDSbz8MJ6lo8DL8D11ZAu67mG9cGv62xKixtFYvVoyy/QUzlUDbqwR2Fbykw60
A0UKyxHuxfTqI6oxPtfhfaIR0pb9a4wEafvMOuZK+YYtBE++KfovRdRMicvLaYC5
1lI6NFjVHG1gIk55Zju108PNGjvM1Q/LUJH9RBSOLJ3twdTp0wNspqXzH5RLDW5e
58pgpmzu8EADjlVHGbu79abuORDi0WeWFXkV0INBP9wEokcswBWNSeT1TpIA1ZyR
g/wv63MZ5fWqcLvb/wLeWKyE19HCP7CsjumpOAsUImMMNgNcARobBpyhYijVPSMX
YXw6ZAGi+ZnyUCROj6+1lwTjyQYkXD9EfrFSlTCk9qtC4ew9gukQy+kxTvX8D4W3
eoUkseNooPcMay2vY9XJlDbV5KFKX85wBPeW55XWobM4S/V7QuR+QYasoGPUcI6w
DCk29IBAurc4wYl+h8VeU+q8FXbTc43gfzukoH42+Ha3i+B8mnVI272DUFDFMPnR
BIW7yevtfdAH/Lqvnm6OVHV79Et3xWbzcz5oFf9+YH30v6FcK23eSJs9UW4wIzXe
oofnfbg2ysd9RALoskRzLWwsGFnsa5CLomiTx/SIGAag9VITLQ0zdCB07UciYRPb
xDQdlVBp8hWmctXuNelqD7HGsdwYjs1//imGGXe9/EDk4NxW8lAMTGret2MQPcvC
IRiVO2Va8zYBhp+pwrrhDfjRUNXtbgozdsAk8Cbq9ovQ+WSpoYKvLrhwE5IIZhRx
FGH148u/t+eB5fkCbG+NEi4eCux3s3GFhyKv4Q1NPQKBOXka9n5bvdEz/Q1HFgc3
LRe3ATRMqsvLaNtFisdzxpkfbMj+S22ixnfiLxrP2Z+5cGxz0rUG3xPQhGzgzc/B
u6LVqFvLaNP67rvS7NJwK6UPRj5gsUk5YCGDQGRSpFKDxK0ZE2cLv5ZDgoLUxsrK
LX9rnjXeimKFXoM8bwBNqIE7HlucARD+QwSQnpqmf2Ix9A1tbHRC+RGEjgFflaAH
o+suzYpy1q+ivmbcxSpA3CH2pXvH4S2B3I4A05zT1wo6rzNTF/iPe4rYHrXIh6cb
WC06HdBJK86r+hFuH0xBaFN0T2zdL1L56Gd76WaQ7j3JLNlk8ne0it7SltxRgLIS
WVryg+BNlSf7mTCkv9AspA9sfoUJ83Le4Jx/ZW95aJJ0ORbyhS2pzD9UgTtJpqpD
C0pmJxdCOKXBevUAwHoHm3v4OPtvAcIZDWdkpAcPz9i6gP/r5OCPV4rny6SEm91a
e8O7s9fEUr1VEgC+w+WXHVtObByGvPNeW2Lnc4U2A0M70hv9sfZAkdffqFjkzcwy
QZl8Q9wfrF8qPTTTxg5yMCAd7vSmInnQL5RAUYtGtsq0DziqGxs/JvwCfZHbm84e
TCecAquUIW0FY7zxsVhY/tE/XYG2MpcKBesBCx9B0T/SNbGWmymWHqAKuwGX8ise
JFZeYyOs1RdM1sJH42Etty4Yh1CTuQ22pljSDVF+0VzODWZTWB9C2QO44JtnU4yF
gbPLqaKvYnM/YC5mZBRhDuapyTQg1sxRaQY9FJE3tOf5YSH4L1ft4lA3i/uEMn9v
/X9MkI6m601lXhYW8uvdV2OnnS+a20RikVOzlVDBrDf0iunf4PbALwsD8RhhuzlA
g3qDmFrSP9kox9gKFZbM7NhgauIyNuRUCDPo1ax2D12s5UaP6wENPT7KgJR5DFZO
DQqTvuzhTt+9z3Py6Jl7oyHwc/ir7Oi2n6KJiguiVeGY1pOdqqAqh/3N+0l1nuuv
PRZt3lVXt9VIvP0Wcp/lhw==
`protect END_PROTECTED
