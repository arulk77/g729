`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zowsZiPFFs3QdkRGFITpCMQLij2QaZShybZN7NQFs/f
YRK5WUTZM3a8xbZUAEOqfVTCUgAk6E4TFvMtIyCJa0aO8SxpZkx1YXP+CU+XKvWP
6Nuq6TowUlSq0KeGomWd7wFJRJ6sr12YB+IAiJiaShRuEbBFVNNGHvxLXKeZuSfH
DBDWREwQNur7X31zUW2ZhxsUpvLY4dOoEFc+wpRSWDy50FA7S2XbugMdVWU5UQlu
d8XdIhRLwAxqai4KMZQBeaMxf0e5/rdxXxWb+UhFAeaMvPwR3c9kjYmoD8qAZt/P
cj57psmnD3xSr76uQYX9PalnhuxCCXz42/oH2jqsHipviwO6FR2pDdlsNMOlP/bA
L1FcuKik54wEjQOMAnLLSg==
`protect END_PROTECTED
