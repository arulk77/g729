`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C65/FhcKiLeevd1o8qWvYqMvNTRKKZXeU2tVuukaLph5
zgQINpVgLJVEc6wEiTmIaQQdLUipajCuB64MoSvFNH8Svt8gRK+1qD7tY0vIl1ha
hQqf2n/xrK/c7o4TJv4VTm6+8tdwHoqrPB/qk3YrGtJIdqMAlYG7wTbqE1t6bsuz
vmqCtV6n4xE0bO7CdKNtq6jdkKNqySwygEfIWPDmDepYc48TNAdl5trt23Ajwzil
DQZQJyKvK8NoGISxQZjaD01Cpk2SpLang6whk7Tih4YlMh+BfIrAO8UUR1bGPQxw
VtRKllIBPd4+wbqYd5K6sT9aj6C3EpRAVXRgiJa5xybCtQ/VVQCWAJrFkN3WyQnf
0Zrcy0h13MY/PIR1Q7orVW1DMOiCreb1czwaqkX/N5KDsqoFf/yFsE1WKrqg8zFv
zdYFNZw7ps0CoonSYdE01FXOfGqjdXExZfs2Dc60nUy4rOw7WS5wnDKpK108zzx+
PA5tP24sIdq/zemQqfCGfuQBmjfnwuNqZGAWsPxiTSanGNl1AdXdLfVpfixfNXgh
EyWlcAMtpjBFpK3RnkR6mJRIpioeCxUplrM6NDEGdBRPCifk3/PyPJv3uXTemfjW
f8ue7a6CrORH4UIhlwXi/0BD1xbCL9JpGUtbX+MBSJTv3fMJJYDegZfceK4SbJCU
Qy5XZE6quNl8fgIGMXtehs65bI4v1WfvPpzmMAURoawrRl4Fz3fFNk69XpYWXoNw
a3m45+c7n7ADYrhIhpCZS/aN6/EfVB4OFGX3Pix+iR1FwAJL3CpgTeF77QwprO7I
MtIMzLawI8S3inVqBAJ0qGuw7VbGhMRw+B/9ppQq2JH0GT3EzgdFQD42mg9JYYk1
Z5avyr+FjKwfF3bbqLluQsN9Tclp3k0zBaxpnK0PEaRn/+9CStJmzyOaLmbW6M0H
bfvwsbUPCFyG/pUtV6nkpP7zkzuBOwUY0380LAw7fMc2th4IQotZ2tD4LXb+gSOx
Dp1p0+GsDE/c5uFK6qGdaTT2ybNwxsBKpKln7aMTsTIBTMtqX5QXbRgf+39sOa2s
5K2SLT+soTcJi8cL3cD169ez6GTqs+JyxMdcJ6EZr2B7sUJJ+yQ9TKW2aeKe1OTp
q93B+WT6dtbdJtxHnAqGEBwecMhBmv9fbzBRjOgeqvxb68u4DtnaMQSnVZ2yKgk3
iC2nZ1M1saNUz4Qh6R60JsYkQPpfsBHoIz0z/EF4cYlaKgRvgRX5CAtBmwVU69IF
c/BIsltuaJNSCUTCK7Py4yJ/j3okKBZmLI9ZsQl66FXOUxsQksSqzMxc4AC0pVHc
O+sfqI0F3ArRMY2tNkaBVt6G3rx2qghkGqraf6jJRjoLVBIIbvnO9ZjiK7G8SkSg
UnkzV9xLPn6Cy5GmZe5SesV1Z+k4ob844zRmSOvwLyq+A/BOQyYvmCWzIRE9HbWL
9lK+vowj8LOJxzmnBIzmVTUthqTnmcm4IqsCNsSxe/COYmiBClfG+0y9i6LXbhvh
dWe4KNKc3kuECPUHqsSuZLBPCm4FdB9SlQjxcIrVTwGY31wA7PMdNsI2FPXBmYUR
C5wBu/OR5v0P4VYhqSb9WxIWouPEZB4A1txT+5koIMHQlOk33ose22EZAT6b2G9m
6/2VFNd4qtZb2JjhewFABz0jNbPFkf+E5TvFyJp/wJ/l6lIdfu6dOW0Wp2Q/lHI0
ANOoAANx+s5aiJwQsPN6gK9Y9Z8Unsdnv79mhYDyx6EfAN60NrBtC1NDu8BKczGD
uuwBl7fzDE/2D4qQimT2LCcjq4oh7DYJtu3x/6b/y3nCP+v8dYfFeg97oUyYLLqA
y43T0D2dJqojKyYeYhsWjRzPY2INzWLH8lZ8p8g7eefXf3+q/DzF5NOZzdMXcrjA
beSoUpYxRJbXGZD0KRr6hjLBR1DgkZJTVpDKslr/wk3ZrnS4/KeI2r2rIkTJbd9l
P2UwJ+/kRCNuqg155cqhEUJyw6G4Yf/TEM50SekRXBKD5Ig7wtIUfnikm84GBVAb
YTNRVdGsR2qzhpx2RWhxDwOK3RKmiZ73miY7Wo48zS9X0LQOBmSrGqf4XIXjSihh
C2t62TWUmQA8FE3i6GJZMW5VI7Ii7+qaBfNxlrPOBJiWqoZD0ZomL4UFUSP0+AqW
dQkOaet3lorK4GI0kYqP+Tr9VD0N8yBbAe28+asohaIV+8CVczs2WPCy1phsvdIP
88iHxBoDHT+77NNjx5dTcC2Rsc6kf52CuPog8m/jJFnNaP3ljxhLdq3axIkq+VDo
fTyHYUaN4GH7RbAjNCHJWSW9x1BC8uMLvdaVoaaPgiD8UgTIUD6Ekrnv2HV7aYYF
nw59I7pFUWjjIV4lLhLNJ00bOWm+fd07t5kt6kCCIH8up8fAP6/mliTmW9lReVWT
763WJOy97M7WrIJ/t47M4y+t/ILJY8TZ0yIEl2+6iQkReA4KhivGFahzoOlnn9sV
NvnUuF7h/ZBy/NIL8KN98l+X3v0i/zOmoKA1sDJA8TxRiWDXen0vWOrUoLwEuBYu
sYh1qqua0F/l7RrjAwtJp+lp+7lSDSTWJlTQCFSyl4wvtWcGWkgieAwlGsTAMR2w
cmJgIfjTZMvvoBSxzEz/iX8uHrsqyUvNQPviZ1OZHO4nLSQU6LtZe0R7lOnaYNyX
BZzmgq5/zrI3w2rqeVUNziNS22sRYDOMfbihe8Ppm5TLP9sIvb5ldcVES9sQnSUd
G5lXZlGFNyNTf5zJqckUwb5n4Z7MawEYtmUztvjtP9pa6IE9XW5h6lL4eodUpjYW
DQM0A3t77n1MTM35zU2FDb5opkxFWhXc67SeDdNAbxIBcHhtjpwT4zRO4+SxFHht
yFrkVe+Aw8uJh6WVmbnKnSpIHaU1A1Oq3dpbXgg2XayurF0rtUqvpKlaHmmXm91B
6H57Lmv52eacTSf/Ha5zcsvUYoaxc98f0/h/u9MD76JMOnURlD6ZOVUUxjZKMz3w
J+Xp3GeiYBCb1OTJZtl/J9pvoiXtBeAjJIQ3bDRYmewNF9dN7AyNnuTvCJ1HMH2m
90rqZeS9tLoLsFIdMW9TRM8bFr3aRqc+7QLazOjTc5e6b+PkJD/92aLylG1fhPtK
ajELorFClqd/iQa77QVeU42Kn/uOR8yyVDAF660O55lpHflmsFl7f+gVjwxkssi6
Hqgv0MB/DlVEEYPM9Zmyn+MtAhIY8I/rcmXo5VVyvUUSQxFGZ7kbvnamB0i3yFjN
1TTnlMossW0k1oliTubJjJyHaVA2MEz5obsWyjqkarB47P9oCmnAo/KonP6CcjFo
QwgeTfjt2qN05dRAlnh2BdEiUWJRfjosu0Xs6NLZ79BaKP9FsW+eF5Xlmi8PLUS1
7C5vKpCzhIUWgrnG6ER79FqR9e2I2f/0mv+7xHVY4v2xW5p5naDV6DHiZFEbuY9X
oPU3bj3NLXKWbZt+tufLK46WG062Lxtt9lW2aRnOgPR8NxQ3g3ItmZMA5I0oUQRB
0X6IemApT9mWuckVUFBasKYdu6gs30fMabZiq8soFUuv3/4cutyzdJSf/zHYJSKG
DwcC6UUWoiOBjUtvcIUxK6DHlHL2QgOvnZlIklxfqgd7qkJv6sRuGZ9fdMI3H193
OxL7l6bFjK4s8T/W/TcG532qQxs7XxkURcHRUfkI/wlAOkfzo3euDUOp1R5xTcba
WEEMF1sDjBtdkkSiJ76cIZSxZ8rGhTTgc3xpTD+AsPR1sB3woi28k2VHGtMy/hBQ
Vs96PQEIMQuJ/byQ0k4AOh9LxJYPZgSDoxYgim6jaSfBJrE9Hc24eDVzgZkTP4zI
aGX1MHVgvIF79r2jdiitfXR2I+vQT2S2F2DCfk8pKbaFWSKaEVlpXWlK8c8jFfoq
RlC/mFW7of2DiHPOUmolU1oVFnwlWw4xjpRcg+Fh0QILfIDzm50kPKOvRG+3WJsv
Y58/HlFmhJjV8/m3odOtpbpILeIwdIGcU6YK2sKp6DSrtaaJEyRKvAgN9Hug8T4K
zQpI3rrHZPin7NO78ddk8RAeoGsYd2O5gY2IijA5RMB1MDb0dNUEWlsJkhiURP5g
fZ5g+KAJkQBQE80wJCcgR8R4hlgsRWDV4rpb7qv6n2aTZpAL+fVRv87kjKmEIDJb
tR2Zbre9zx3STrA8jUWnulUFU6FjAj2ZBlMTklgbgkBCMg5wZYT8ZTI0eRrk2YVK
UZE4j2hu96d3auBAzFw7/ZFT0Nu4UsvEmUgHwEqdmc5/zypzESdjDkjVdcLgw7wd
2QgopbGu6Y2wz0sE3GLzzLUvTiSDMYfpFyDQ6PR333SvY7WMYCDBf6HpIO3Msu8m
Y4insOYfAyqJjBO6N0kkww5dRcNkF5dtj/fWY6J0oCjnqMb57C1kPw++YSzblj/X
0j0d/eYF03Y9zpHsBWlR6WwMoeyDeLwWjKnMRmhycEvYdMC2ivzs7mDg8HcmJblG
JKsHoO6O5P+ogL5thorbafqYG3EgUQoMR0e59lqLR4p57xlJZEFPlDzppV60TY23
LJaqEKEwpuhkYHAMqf8I+MPGTYNZQf/ExjI2Qlyq3ZXBMJXkaU1EKlhGoRRT8vs8
bqyHVVlGSxQtlC1nHKesbY3nKQs5KolWFfPN3yUymxNlsQ9WWcmVxZ9ugZjj4jR2
IA2QxdVjjCnHyjiv/m8ZX4xLqQckGbb+IFpm64ePMjUk3OIZrPvDsp792AbjULiP
1hPDqUMcZujJiWNs1Jt/F5IgbFVPw1DqQIbE0onneXoS3CtzWB6OolILo6o/caEK
Yfn6t0MRv/6oIfdSEWDV7NLidaAmSECiErIotWDASnSkpDaLxurrdbOF6LpclaTU
d7B3pQ56lR5LxwEh+ABIwGSicAm/kEUHJLEEtqLm/B9458FDPgyLNpPrYGfPNPuM
zmr/INfMWySEuRSGPedZ/1326rIcyXmx1jmN97xutyf7tmqmKGXL4iCfjYF53qlI
gE0kfcUWmZDpd6cTF1ru7+fBrYuC72yj/wjo/tesLBGs/RDIGsyuIs5SHWRVQhxT
kdtzhyiNmrLxwngi1VKd9AK8RAsymK2ghC+/nCP6NnuLCpXca4IYeQhw5fXoUzBX
XdvMRY63WVer1X+nJMdlUkaqw0qCJ3c5kGG3u2lacXzjUk7J5W5KfKjvs3CMqFsn
ik0CguyHSBphbFwjk7y/OzSX6jeCB3YDHvYY7/qzSi95Li4vcYKKZKStVYq/O76q
BFiNZ9yYQA57dpbdL3/WnHptv0OUz24hDvEWO8zjdTYEWoZh2VCEKMhQO/q15t5B
LLxD823xKb8LM2bkNU4q22zNZit4G6ymSdYg+pKu1J9DIfpSE60NGUjgSa1C+XQF
YkYYm54w+ypEEd1FZteebTWgSNpn3NVO+SQfrF546TvMjpdhyAxJNhJGxTMgqhyc
622oYeB+5RS1/o2hUL/Wt6CCARgy3iTwDnS6blkk8QUA2lxqq6VBPmcwu7l2AK4y
5ezPGFW/R8YOtdcprFKRRytaArrKNttH9J9j+CoovxrzI02nhQOXqPe963f7xXvs
45ilf//guA40uRZH0GHYfg5KtUa2RZh+8aMhQxlc/vqIuU3a/Ulv/qWR+eBf1fJJ
k3ZxV4A0AadF1v9bI/KSQdFbzpyMyZJNKuASlovHWGH9446d9WqhWWT4AjbNDX/C
91/3zAYlEVhAjyKoVXruU9ltbDtqtOC107npaXu/rRebBW/Ly6P3jHB7RdUgr8Tw
r+KtBIcvXB0UT9zif6+0+B3j52dC1Mrwt1Sg3qHj9xC5ANIcy/GfmFmaZs+T+j1/
giUsX3F+LLdyZVaE2Y0rSq8iwvSt/ZaIHl0BjF9iYxsMOQHVscxtXhIuk4gBROAV
cb0XzIpnA/eiXEARhqS6H67O/CE7o+4NPbNd3X9Qrx/N9bpmYyELTuRPpEBtazvM
bAfnvmUC4K4mq7bZ/QSbnc0QouB9xkELY1isxDcozGGpS32KegaenyFlHom3G3bS
oCqWKJHLQXwP/LCLMJxdOs9BZw+w0HeX7VzlgZWhptg8n8aEVO3gIF4TdNvFKutN
CrVhmBJCt6zypAch/GZG0FQRqs4iOyqK/dzuRZvMHQBcTuk/YIhTZNn1wMn1fvDG
HDz7gPnTFnQAiRDecTDaYYITOkNTCZe9zjT5cTs/oK7/vvO0mR3pUjCefm6EnWMQ
2vfAlnlb2Ktg0AVn0pcydBtPn31VV23dDm2GMHOSmPpX22R0opRW3HlvR3fGRGx0
1PqyWrNf4EiefeXmCd/GV6vjU8OcQkGB/IIHm3JRn2myU4u7phs0IT8kLkXajE/K
s3GOBcYiUlhtZmpZ5IVJBL2LRe4gDchgDXVWY5fEPXrd4v2SCOD8uTPBYcG/2Q/3
DtJWvtc32x+BhzSmv+2ZKKpkCoZE50Tar1JN4k13oQHZM+WzkEp3XETHhR7QgZ3Q
q6lujtBt6RU3ZV3wy+6bMcvUrNdfaiFW878YfuBZ9PNLNjf+HM1GTN9zzSpiLMlD
uREJQxKk//9qz1odD1UymeZ1oLiYOnLTncVqGr3C4rcYW/bZBZU5wDhX6czUMpb3
Mu278RMizWyKr//LMjIUg161LO3sPO1oDRes1960xMtHqxCMS2T6tUT761myLx7H
2TIcVcxOryF02BQ6LWKnrum8diBLiudMfgUsq9IU3F+F1rEO9+DlaoklAjP0L+e8
rP85X661433HKtvw+5QiKNZjEN91uIlq7EK2rm+vtnZ0/xl9SeTd84xDEwPl6VIu
Dqk2IQsVRrYeti/2U64gdEcb64NWycRJHwMLSY9CGxhP2kYW6V3hgLRIm5nb49D+
tzoOjN2Xe0Wwxtfd93PcKNpjgo5HndPJ5x5HwYMwvOkrtvlg3GxCImKcMZf9d3mC
bsgrc4NrI18uTpzQfRdg/oEHvBCKZs8lHxtN0uVcjzTHeI0uocj506y5E9FjoTn6
QKmSy2oncW6Fj8fJRWCJ/qHx0M9IFG9VgzzBNPOF0MbvcJrWfv6lHvZiLQZ5IzyE
C/s+OpXzSQnEBHkLTD9p5aMgavfym6mVAfEuEoQMt1BmTU+3ootbgyzSJy+9sgTi
beGoaizfEkolUOWf5kjQ1Jk5KCABJ6Nt1jOQb34OZnHc0r40iDqRMH0t/mL+6c+8
Ju5nIAaYRWUH88OIjsgYHpJbPe/IBLvH35w9cVdgzJx88GEUFdiuXZbUw74bQC96
kT8o0QOcn/rHazk5xp51g6hznmG60kLZqDig4sWhpVL6RCJh9Hi1+f0rQcuSF9pr
QuVdrIdOGBtQRXPLi4g95lq/hC/2BSEpbOtZhZ/c/GGODEklRBWWUsVLdqVWCZJ8
vb8FvOIxarUrK3B/Eul8MiFpT7n6GV3klTkhL/mjfAvjfLP2Ow82bdDEeaQw8uXm
NSuza+4aYkDp0TB2ZFNxEmI+fESZ4XwiRtvaxw1Ly1NBnnXkjZozcGP+n8w6vIgz
MxHPalGnG9dYxkfR0hF3WN9fe3AdvFD0awBKBqw/LUc1lRym7vqodx4/Ho5S6kBC
qSxdS2DtnjVmea+iVhU2DrxupYlw76Gz1ijLCr2WaxKOIgkiHo325JYe7IcgXhvR
DQQKrf6gU3UDERrcF68hzpBMKhgWylOuzd2EGbtztw1OOvSUgVmt4EgnEEIW2vch
6DxN4eksW2yF8MC1lJ/q3vXPikzzbZtVOTCpZLE2x0e+Jt7zVeaz7iEo+V562+5h
SXnLTTBP81zduS5kRH1pofVJYNSb9Mus6rLX8vYiXLGe6goOB98EGHg8xaP2NAKe
LOdu1IUTc0BkNG2w+uzIKuHw9uqXwvg2i2N5Z5B5B1p00QaR4C2W1l/LgePcBQkI
oTgwkA2Ly2rpI5ne8zmKp91DDm+dZaFFBliNkEjKJ4XCemERgiRy3ZtkFQFlbN8E
S4pSN90VeQL0XBrmYOVmwOcG7seUv8eso6umrj9j/D3yP7inFG/4ULDYcwpTWrOG
UcdKZw0QqC1fF1Hb1P9GWLivOW+U75YHw0GZjCEUcabcrwNk+jwo4lex10jbXD9/
oQx7QqwyVfLDVdI37zQvm3R7pJVBz64bJ07WkiKKkW1ig/GrPk62pv6Y71Kwcim9
EQdO4/PcN9viTdCAvOi6r9wveUVCHCTzRRlzcMIFquTT6LNO4YVLci56L0xw+1Gx
jy/KgtCPh5TUysK9FmdPJ4zlASp6EKX89vyAFqshv1jJS/oocxFU291PGEh66E9z
BB9OXVK+8DjdpLpDgzpgWM723zciIY5SyD9dx5C1v1wRLZtXhVLfhAuQUDzXsgTP
FV5VF7QqT0yyfepN4gg9mGZ9gH5LaySHGmya3/GA+9buAnp50PVswPgML2LZI8K2
WrnHT6JR+Tva62b0JGR9CjF1BzZ3b7oRETl1lVaPG7ScNDWUvVSvX/iS9bqJpHBZ
uSib27JnIcoFJv+vpekdhV3GTO246+jpDfgX+l+2EKDc1E5pnbnx0pos0y6m1Jko
RW92n/TxbTZ71nxywC8WIWSpjqJ70ciR5lvKaifshB5cVNudAlWKC8SFDaaIpytF
uJHDRcd/I1r+uagVb7bEiHobIonzg94zIyJsy4Hw38aAzs7avMSrfgrpqAg9j0td
UWxTqg7oniLJd6z4eNYjMFOhKh3qkxKlDZM60CoHFlwvt/lXqNte8jMpxRL/u/jR
4M/jEnmNLIyUqggBGklAmefll46o1qJ+1IL6YhCPqZVbU79VyzRORhj6KUo1o2u/
m1NcZ8x/Y16vONy+jkNu/l2/mcK64J95us/SSvlve1ilo99SeUz0XYahWMrycaTx
RKFNG6NPHsukJZUtasesf3ifOi7GyeIw9kKg8opwJSGzC3vopXz/6at21D0NV4xQ
2HX4iRKTApDigD39ry14aJ5JLA9QTaD3l5aDTZRs0w8ZbvDcDw4BCSuRHHNdnJm0
dFO8dEflYK/Rrqbnz/wQmesh4R349a9LnJWrZkO7/jXps5CjfTK0dkj+jKCMJIAS
abazNViRumrjvOtM+GMY8QFMz5nqmyizWvy3tCkUdQWGrj2CmMIc8Q6YbxPgb0O5
JHLyohrI5jkOjqLMhOBzKbkfgQks/VO9RIZaZ1jfk8/IXT3JgzZSz8c3aQB50ElP
Yb4ikK781R9Ot+De0dYOWL4rHSs7krr1Ii/ZlTAamFXsM87USEC445o0o5cpOk+S
xoERmleX+5JaYSryk5SqeBpnaeaG29wkR/T0OJVAoswdyQpSVplet7LbJEQLtty2
RLI9GJTrk/wfXQI43D8xiqW12syWP5q+Q4PlYZ7/YG1MBs4sfmPOM72aPXAfYP/M
sczYE7OQUnxFFe1eRy3fG05pdjK3Vw/ZlOZ0b2fwavqetVAKdfR/IjuS2v3uMXHs
ueZaiVAc5jNBGqykLtg54gl4Tcu1juneNvgtQt7I6PWRH828QIS3HYTdx9rnPvwo
PScISfJqKOJTl4H/vgmuSl/CRdCGoehaGcUDD6Zl3W9GGlBNqHCie+2WzDkTWg28
BQrtFqH30Rrfmub9k4NWHszvUwcdsmDG6hg6h/QKbUYw2Gwd5qePagpCgn6mloI7
TOc3MQxkxwTFKq3zXOwLANMCo8T1cwa+igq4AEQBpZTsCZXgiWc3ajS4N4EDBiJL
ZpwLoZNJnmqKDppK0f92hrQ5GWDNPN9paTuJL7vuEpIgCH0NJXv1rJONNEbz880/
Una88XBhE0opjnmmLFBImlVjyUJm/DSFWKWYj8rsh/Dp5+hqxq1lWBaH6WezXPwm
N5I5JDCrDu0dS26VS0FkZnojDuwjys+maOhZxiaIb+LhZlsa+OZ5+aCTP+5GJXrP
dlcB+Nl7UjP9IfKT3jonQuWebnajcmSl+LXVTwwnm4eiZJXl5qTtAYeJoyRgsQmo
+3OwRGNc/HIKjYOtm001xPNwwcM6K3B5TnhyT/WPmTVPVkCakbsCUiL8fU/YyboL
aHnOS8GFESo2EVJbaZT9QTVTa0i8i/Rmq9m/8UwwHU2x1MK2O7vW9/HvY/Rm99iK
r9l2O4OFUZNGnP+mW5X3v0YbGxMl5rHSsVyPqALH5CwGkBXpV0+z2CawPHQz8v+g
0xrquRVk8+s9k67TeLIykJVi7VfQkltD379pWZhE5Mt8hsByACKEZ1VVY+z0ire2
W/iAPETDwmgbEmPf8DTa+UNuQYvg3MQZTcaVKi6YDAmvEw0x8LTvDWhZFyFZMIOO
gBJLajXC1/C/d4K3mJVOkHrjM3OatscdCQpLmbn+JyPDc35Y0SUEHQrysgwn7cV6
S2ShDiCM/QMBp75YUdeWK1Ksv6ncSGTfLM8+7ze/ayt6Q0VEVsQecj6yOshyEqKx
pxwofzmQlGN27/8qr6XVLll4YVUtP+N//slPVEDdQ+NweVfvgxAzQVXyXmCmvyOa
AKxOINmCInhqE/hQ3Awp6i3pUmsUajQ7FRgKv1y9MyvcJP66VgftimAbuPdNBBZQ
7bEZj6kVospNM1Hn33Vw7TIHQWxitD8dajmvPGCzu+DZvNTAspxSeaqVR5c/apO0
naCIxAcBeupZ/3/Qf9+ReWk3j2o+YMBOJb6ED1bi8YbK9Eb130SNlNluT1bb/f1k
CUdn7pPEIjAg2JPHVwqe5tDy6ZwPMensCPAnKmjXCRL+dlQBmLCy8wellfX5Wqz6
7rDAt3wu+ENMvWxJgh/+XYtf7s0OPIZQkH2W3NLiKzlIM29Rng+ylMKAdYgPyKAG
Eou168tzf4kHsupUpFJyBatixxAuuydxqxdw1WvzdZNlsWGw7uFYEUVxVa4/mhPM
ywcGptdnn2nGTeNNNYZUpM0RH3xOMFy7JGBhOrNU246IsQyDWyRicZPM2kHYk39l
SxfWRrKyhx3lyTWRzi4b1njcO9YwhL0688IHFiU4OOv8wxAdV6ru7jmK1ENal+FH
jLMXYZqOOJ0jzNHH1F5BCMCzzFHsJTQSLlUcBfNie/kJTrmxqED23XqiHZjJlI+r
U6gYQkzp86Sq1PPEY3v8HJTrd9buUPNbh2lcWXc94JQt2qXVW44fPPGBAnnt/Vm9
Aei+itFadwiKvTXHUit8WBn71QNqDVP188snihSG3xzOWff9Uk3XCcE1XD5oZ0of
Te6m+utaoVjJ9TLSG3OR0c/+Xo3kB/ze1oWi03nC02XF/9EC674TNFFRKJ3tLhrJ
rz8jhz3OxWdwl5THRj2mBwTJKUMfHUkUkhZjnp/MmL/D5HkKUaNXVmHft4t2SFzJ
ZqynxCEWMba4DKgFFSUnMSrgVK1IoP+XKjwWcvN2uT7wIkFaTzSNqC1fjtnMxDST
1E4vHgJcV8LkxHzrhIQPhAAR1jGcGpXmIBzH7Pp1sFAZlZaNjCZurhGSEgs5nEnY
XznzMYpNc9D7ZllKGtDv2wnXvmFQVwU0WAhu00G/shCG4EvtKXFhIyM2IPkn7pE8
3nZ5QafHu94NONRQMwsbw08N7uqN9uic8XzDevBYRUoeNd3C422HjZ8KP/xoIZ34
zwS+ZzQAtfgigRydNtoDJP4wj4ELrlhZH5Dkp4J3XQuBi7GKEEQvmrLU2BCHbu1U
NiaWgereWXKBG4zyOY5VWgXccbUn3+XHr1oTzioUOxO2UFFK9Ng96dwhm+KoOxhW
+VrJDiYow6G7p35bSVRO3CCFERt3cz7nowDLssw9lqwqRKls5i0stUPMpxWSkC5b
eXLJYrhAKMAvzBGWLEemoMrENP7JOkXYrgvf2gHMaefrgtHux5lBDVgw57r5Vvq2
XtybmK4G6hU1uXlZ9P7T0ZcAvT95ycPOVuxnKjQDY0+lk/XstfGxZN8DrUlWjRGn
0MSOT2XJhr9PtAVouDEk0Gf3KrGA/LrrVYfoZLjGMCpvyKuQyOV0St8tvl0PrRG+
oX8tMDqYlsCvGxjEIAbtER0KV0AOLolAvGiDkBtTg10Dfs78hwje5yYgmI+1qmGl
jz+3p7HFXFPkRkAAYhUfG3xBlaQbZ2M1aREWX4pZITShdxzZCJ2S1pmz54MEexY6
XksGtiviwMTrdx7Bx8tfxJ40VkQz7y+1W3ipYQVdEMaFbYfOusjtXVB+wadTnSm4
oY5mrMa/h97fzis5L5GRyv7Gr8jr5xOFdbxaZXgGjv2eS5s0mHKSq6vUTzSgunDr
bV34GvUAXTiYJtogeDCo0OdiQpIqvBSZjBcP9PhvW8bCofxjRg+ujpXocwsAuB8h
P/5BLueklXd08sVNBOfAQXZfeCGtUcuNSIoK5HVh8GufswMP/TxeeR2keC+yEII5
UMBvYNEJSyhcE5NrahnX1oXvQFsH1jR8hBnIq+X6BJfTnm6NTnDhKVl3UrLlB9Gt
XHkz5WQHflWUU4sy2U+qKCKYxg/V2GJBB7pB5ZOgayE+rRFHosakliUFdyL0GCHL
tHqWTiC8jGpijEmiWOfwDqL/iB4cJZUzodlRjnaaqPP6qVC9+64vMO4BkPaqn/LZ
wCBSEfUeMvgPig02nVKrdyJDn4y0TLddl1RG17kSe2ZF572nX6kKx5ccodw/x6ZD
QeF1yKQHejrp2YcpIaz7JLij05KSa2tlzAEdbOqGiHtSxKvihcXexGR/gdESxlkX
Ric/BasZaOnmpAzMhJ9X6rAem3okRWkkCqfOpDLqgCybCim9Fy75UOYwiS5jgqeF
5waO0Wy0SEarxisepCuRpIeS4WW3LO7tVBk66AXFRXQ0eov09KS1vpTucoze3lIt
NuuDUePIepo05ZNNfBFld11UckeDPmDBlTna33U6mLjlkqfrUzWh8bZx03chd3re
tVs/H0tGh8Ms6y8uMNm4hOfE7ZW1tEBcv23N8uN73/tZRTEtMdfFuAPYAYk0T59Y
Pgf5WRU6FS+cOOs8BV8i1YN3rbzGUZuzLUACKeVZtCk6k//jZYTZbKUczz5E7LLj
Qta13l3qvVz2bDrSAzkMb0hJ+ISk1D686gwfR/FmdV9vHze+2gP3xrhLyiIi3YPO
N9MXuijnVMfC8grNdRkaZqQ2ntSNehS+s40FjznEFM7X6Qf1ucJP/+1y+yBCbQOH
/1UL0dYsa+4XCnAWTSFXl9zkM6IT43aeNurHB3z6Rs9GAKx7c5MHBtzwk5Cv5l7x
Bv/Zb62X51qjmZW+cNPeSHEsV4T/Eew81qmhcvy8QczXzbWZYVMlKvF3U2y2Tncm
7MfAXzS/fkZ/gPJxXXc5S+fJQyyVBvJqNpvaP/5chyHrTSo2z0duWIaMCFcjPPzs
1YySNOFsekszQNd+7YhyugfFcMBKdbFZVpJ8zRi2Bq6WggGnhJP5k52ZcOHEn+AR
/GfdCTJaM2fNhMTTW0Q6HYrLTU5XtbNfyCgj5kAYRrpG/cHzzMj/m29jXuYQYg2K
iXRHtGvvt1WrwajXsfP/V5ZcHeugrsU20+cjeaeDsEe0HyQyo2R3xeQo5i1SUXU9
i7jZWpI8EGrJ+lSAsxOSTxHa4DHsfNpZcj6/KLvCUZM1BBkNzyBxJTE+X9eJPd3n
5vKwqM+AkzErBBCGwTxEoHSVu/6Kjn36SMnankips+8w+w2Q3/j94CBwy4FNvMSU
dN+xf0QFiPc1hPrBMoxSuWH2BhcDKK9Yo+BsmiphtGHGiMQ2nCjz8mTHoJ6Nqvix
FT9PBBtNfmfhnTs5Q2JLrYYnZA0bR5lo9t+WdKfDdEBeEHbMHuuJIsLqy+urdmj2
cOFWST3Uxhh/sS9oXzYKa+1AqZyg805lPzFHnZVIOmEQH9gHerR9UuGyhe2p+Z2Z
Fzd66kBYMdko3vQeEMjNI3GFGD9MFTTOomZr3dU9GmGVKGoZGHNslCjHqUcw1zn/
w9QxVwm1+Zhlk97DWDPmKpoigMpmo+12oyhWw6O5ZJKToajmk7QPCz7T5cHSd6VH
5LQ4PGsncxfw2ZoEosl/9MlJdQcZhqpdn0xfgJdIQ3I3nOmBi1fOPF29XBHBqcgk
I+Ryf6oheG+vCLQmRearmPrg3bXUYXpDi4MkkToMWhEfquh+iaDRYTrRvGBz2/rt
8flFnG50xropWQOefVGDbg5dgEsX+6SGsDhF42iHyp7evstsNqHkevsUq8T5pq8G
x5nXA1xx1MyEzHCTA113hrrAxlq+U+k2AfcMN9sNq6VXlXmYVl4BoH9oWqEif5PK
ShVzjCWYxnCPn/qHpnWgtIiN06rBZ8h4wgzcC7JNjMwJknq2Tuj/j9/Qy8TzxmfQ
lTuJxu9A4dxPQsozWOX4bBNY+hWxfBEPBUgwHHBhW98V6HuePvw+QNE/x1/S0lGg
AUL6hi7qZ8rXhUzhncFMRAMNA3yKJYO9RkQa5SHK2edKIY6Xjh9hFHgugRueosqd
qyMugxsqYgh4I26rkqda3Q4Oo9L8yddYFB3y6N5jkkEa8oevx0nirVZLez1xgJUg
LxQoUCwKYxbJsbGmtJeakDwl38RFklEKjPuHLbU4CUviWwtpDPuKnwNIpr9Wu1uw
TMyOdI1V+kDfH2ugEPqCPWvbQn9nmCrynHL6gYRxlrMmRqJHUowDnBWWnvxb5hN8
zNw1JvAFLwMnkKmpxYBeuEYljsfSVcmgB746vwmu2Hc7jADNjH9tiADx8Ufnsg93
+tkBq5RHi88Uga2D52M2kRy4R8s2+1mvh28BWHegWwurHfrXK9lcw2nUf3ud2Gr3
tLfD1K3dJzcwcr4NPz0UEQ5WrkFoQo8+lmXrG+PW8Sv77/DFxnJ2yBB5fvhyfHC9
DOUaNzvnobZUPfSqJCgXYDNFPcEt+DbmPccP78uywI9ro6rHGqvoZDcR7OqhurWA
/3JFp7u7Dvf1dvMK9TCEa6T4TAB7Bj4dU1qxo0kyAIwgpn6jIUlhJvmEzdswP3F5
dGrA8kS6RGE+D7Kbn6LZ2KvggFRKylUhbodKs4cz+9O0V3t1RtXhinofEoRTg7P/
uM/9nE7kV9DqJTKLa9KDiYt7LZZMgjNsb1QBlUkTidifGwUBXpcb41d8CJzqhwOq
j9J20mdIrGVRj6GktHHf3hjH8c0Yqq+jMa6dveX97UGp82M4cyZFRdmCp214HOff
NnT6OnJq31f25cjT7cmAtbH9oooczZuIiF8+SJ/lOibHWjFCd2oKIem6wdh7uYQL
Eh0O/VZh6CBXhUEfzBDVhvFXGvIT1LsBZUbJGiftHaJnkr4cn9n4yNIyGaySR7UF
9vxWK9JzuJhe2xPO865L2Qo4IyzKnG7zvm2sJfaClVcYSDxwk0TjLFGNaXgP3zPZ
+NUo+q0nDGii2jLkGxGeOwQojFP8AeSepwKB8HSpUPTLmhol3JZv8p2wxwwMlgIx
Sfr45Ldt0xdEbW3KzIUJtQsIZOBwp+5VPuB8aGS0zDEaJdf6lMlBMBMaQhVFrjDj
ZDq4Ynfnm7FlFiwrvCJOwUjuKo4BfTPakxI9MmTuQpj2NGHHzsVvCsHEgYv4LuxP
FdKWe1X1lmYyq6MuV6JpK6LSGqBo/UHfP3vRBpjhjJvaQkZtf3LMUI7jRvCOrzGw
Tv4XlOxSqr/u6s+NjetjMKYNsDPeO5V96CtLJXPEgI0uHDVWMMaliDGrJH0gOgQq
dkRDQMohyKyr+H5jzqiuXmUOHsJE2+5HRxPmEohXyhtpmX0jqBLYjiNfqQw9ZzGO
XEwL7wpT3eP3a78o4PhhsPTqgEpAL8aikGNgaM67z9Jy6BwaPPOV5iho+lPkDwm4
/Y0kx3nF+ZP6iU0UTFaOPJN72Nkf6D23OXWEcyjn1x/uvah651UGANeaMQpOrTn+
1k3Uiloj45oK97jNkNRg/wHVSQJYyws1H0Z8OYaBgfzhQJJnLKbPTeWoXy7SeRcD
imbm8MSDh2K75maSid4/Qo/pIdAbALs7x5+Bucm/oDMRmLxCzrhvZkJw8A+ukYbZ
gn29FiYjp5AeYeo7f4GFJu0RB4o65Oaifv2TOGynpJgxU+anNOgmi7YD3WFhmx3i
9STMkpqUFJHgZa9PwIvI/4ZY1JOuR15kCiOihN6/2vaDz0+kS5QRFniQYsTHwBNt
ombrM3p/LdxsV7r/8td0/SqlolnkH0riZjgRaugu4muZOwGp+6MFWI8yaRsDiB+V
FRkHiAZV2x2Bnt70tOe17N3Ap9nPoAyepdZ6Fex9nK6VspWpmL889+FHkeuCdn7R
f1kUsPLyxLJQQNO0YoHLX4w11DOdb8wtOl6fWZty8Qgj5A2O6/Q3Qa/LdAnUKeLC
yZ42A+eM0zAm71ZrqDlMAVFHnCJgV1Amn0cIHdaMfhRwqL+UANUN8oCZOQy1UXWn
lEoSVHyS/iZb2UQ9ZkwxWfMuc4SKF8irl+2lzuRWopLwO0sMKZHucRbeS0Pn31T8
fP/CSaBdufThP0+irKMqTrCfrnOVuhxW7kReuUCh5B/VyFRDJ3GvZx5KLd05t+3I
Y2BDRZwVh0b7XF0zPvwtE082qyElOuhT49ciE3LNRW3rVkkCftaYeUX8fvohkO5s
AoXvSFufq6Krgl+SuQe0HbWNqs0u11Bv+eoqaU0iMiN+JGJKaByO0O1/ZhrIL3Vf
Gl8R0/EEp3cRub2deH3hz1rv1E/KMbHsGNJNaFtH61FCO18FcWL1sKkMcaX1U2ec
/57AcurNW8D0J1kxuhP4rd+CXbog263MSghn3ScZK5xq/6HdAOleSLySNyfbwo8Y
/zbsm3ruTlKZqX0jkoqYPcjirn5yNT7FJ9WjmxHe16linT6DSPMjE2hneLs+HzmE
R353MZBoB9QasLw8/6Odbe70oiAcbdmspuxx8Gva0zsWRzvZ0Dw7lEvB+BbGl8rm
BWBEzQ6V629JVXzKG28IyN02iPQbfKNGQ67VM/PchrUPoIAt15QH7NRWeCMWqzxB
`protect END_PROTECTED
