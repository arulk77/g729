`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAQ9EFWbSR59S5JyhrBMoftxtlfm4QlNRz2d0kRemLW0
4916ZXddvdp1vQR1lsyAspyk1hUuHOQruYdxzNWFNbVUkUpPbbkutYa3KfJhJ0sz
A7ctELJi1K4ZjsTdzcOoCJEm+AO4p8X2qrfCAyl2TCEBIhtKdopLo1UN4Ethl5qp
dh/QPjQz9UpPqzZAcdKU1Q==
`protect END_PROTECTED
