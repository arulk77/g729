`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
VTjQtIy+tbvP3hGU077+tED3P05PYZMKSFcI/9F9jag+WgqK8xqYNxEDQjMFeUab
FlzQqrcoXc3vHWbs2iMXJ8ggQ5F9rnCksmz/3b5OSDOvtH4Qer4jKXrMAXfQzQ4O
FRW2SS+PTsFl4EzRlkDRl5k4CKkw0g/gztEsoPIbeJ9W9+5ocIfAPSEE0waZFIRj
wvieOGG+pFrzjVgxU70rtpaSBeN1XLc+IiFlCSIg/wVuC2BEGhZJUn4qxRk0PI0W
zRLEWMGgPHXNz6j/nNYHfZ50JYSYDHCW8vpp7yTDXuxs+MCqm0XoWgz3aWRiLq8B
BCOPJBArW4d8Zj/ASnanpVhNYRl5rXCtn9WZDKiAzT43tuoU+zQWnQCL9dkF5EgU
ZfSrrYwXbtF70+/CrObQPmCFDZJUFxZ/YkLzmABJaIDiLw4RDs7aG7cRYib1nRnM
fknQ19no1c+vCnDz2bUV3PghEp5SUURWs4Fh1J6wSnnI279xadqb+HCRJiOvajpy
z/IU/MmgcLvQrlwKQVp/pCYyZD8ViIqMAI/vFf/rxBGGUz+UcpnvAqeBV16KcavU
gTPh2SEJ4G6rHc4KmNkaMIS0/UM2/+CDDGz6qmm58TRcapmnQuMKyyW8CtNC5xH1
08MiTaTDCSt6hE39arpwyvEShRXAMwUO59iT3Z1YSOQkBO2u5OT8nBimwfT18ZyV
zBJpTysc9CNw6EwOTugKFcq5tsOQnFpjOA0IUS3pECmWuNWXJbr15ODcz58JVD68
f6nmsBphDKd28m4rFpzwDrN6puB0UfdRELI1jb8H3/pjw3ajrsxeDB24+TcwdI38
wpGtfPeKulu10j4BO9tCEUo3NLhFtwJydMjAKOKfPWGu8y1808Zd6BcyclY8fd2l
7D8oOO8U5zr7h6w93vEQm3efPMntfRK6rmwjLg8ffVglpaEx1yPPn8uBKIfjkrve
BaP33WQww8nkNMqSolSGslSrzKsAmR9T/fIDvvnn7+OEgDVcmOcz9TEf+68mbQYS
/x2SOVf8oNNSSOo80pEzqwjzk7iFmZL7EHs1Nb08l/xCpsn/IaWYO7P5ugM3uf0u
ggbR3ohx9QaVhoWT2oxKbBdskhbM5Zksw2tjN8jTdwD7a1sCjBeJs4iRUdpgFa9W
fAdTQ2usl079UWg4nwsMavVx/0sUjpfFWruASigMSg7hOQlisG2UN8bxGkbY4aAv
sZDA4QalWW0L6e0JCeHOpSG1wwLEfY1F81nse9zAsZLhfNwg7Uj57JhffVBG1Jjg
OF1/KtaLBes2h+CSf8rT+wYNrDKFOvgxDE6eDDtcfaXq86hd794f4Do88TnUej4r
7CzXKSB83v40+zQPOf426jyJEiJ9IxRZ8VxorjEBG/gydzx5G0u9Ir4mJBdvxdH2
Gi2oaO1Qpx8UzBrKxCDYfXTGxst9bKD+Ht8P5cZYy3G5lJYabCkD+tqL32ypdPc7
Q8sWHkI6IiLU8f61h4pEv3hbAmBIdeTy02uAmM1jpfpV0Ds4ZG3iHAAs7Zh2SlBP
LJVdwI8mOKMwaQmvbsc5H2i6WKKK6szL4jLVS+603TsD30hR0l/YUWFa6XxPUzII
zDGJM6dpnpTi0Re1hr56mQbe8rcTJ+G7IW31squ4HZzioVRX/XzzdhVr9R3y0bno
Az9ThdfLTZREhIpKmb0VNCGqz0LkPm69ZuLvj8b+3NWI8O0XoO9Z4rExN3GND6Y4
tj5unGFLmca8S4ie5tPGpUunNR2WYS+mwpgvPWFFPJLRDwdA+xkhr2An6+6R9UfF
X+n/8bom3x346LJZKs34ISILFu8elut3SfjJtyFDtAkHNGl6NChIGGh/2mV9Bww4
eFMWCCMCaIVT5P+BuTHwYz/fcAPqvOSl5o3cftJrd9nh+fyoieceAIuA9/nYA0jx
ZdarRzt71jDk0pajqguSCifHXMg2WPXKnMxkcxU2GUpGp2KjLCAGzRZcqyMOgKEO
gr8is1jjPe9D1jDf0z//W0Bw6yUbWE6udCKS2KklowKRqkBG878X0R2//yOG/SX0
PbI4slm5ncwu5T9A/16MhCpjGNmP6YpewUESlQFVPGZwajTFXsVtT/5CNDc0/jxM
deg7tkBH1oFL4ENr8TXqW35b4nFYV8pvNbAOsy1cFZ80G9qy1hApUFz0so1KiW93
G1LpGVsyTL+arKc9LOkLuY5F6V4iclsQrpOdLhzuxG7uqnuB0ko98NxRDYrOAWEb
JWexI9ZLz6gSZjEsD43v1uezjJSxPIpECxS8ZA66DhhfnJo1aLzc8AJTuU8aPwU+
RE7BuIvWF++CYiBf0Z0oOpqyWjlMfRjsKBvRp1oyoGt6WHitrIidRf0P12lAT2hd
F3sYVGduO+aYctxsXFbXfSl8M+Lu7yC1fbs/c6wZxmCDbUY1eIKJOiWbCrJyoA2a
gKTuQskx4iOceyVgg4oORV1axYxqS01NBQYv3T7R+ZHm9JqIT58a9slJRlF1CIQt
DR9aF/pm2t0DCVox0824O8s2baf0WvnJmQHWplri1in5uFOY2gwSZudKMDLz5ur0
DloH9Zdj8REYuwHfvZskcV57HflysDWgXbEJY/gE4TJwA6Ss3pBm4pIYBOozq0PG
ZAJhoy9kstuoY1FiddKRowWjJUva0nU9WBme7uaKkQNL206eEBX2LM60WJiAFW1k
kbaPQekZjN9FMN59g4NBzek8HkZhffvDYXvtjknrO3P/ad2ujF+nJ5fMJHf+jXnd
6QeoLeyBbr31z9X+Qy7UWj+htkCrR8PT/c557eIPp40n0EHcu6KaAQPeYEkv/phu
yio2HsE+kb+3HTnu17FxtuJro2FcbnOce1N3uYXrju3YQYJKv3+bOVh7CXVPKBqy
ELwoUKNzxnjrpMoZR6KBviPMTqFJmQalCEhk6YBYwnVstfoFowSaVUkmxCXNQbwt
O1be3/xih5l4hn2SALiiQwSAg3sEcJw5rdlOe2iRNVILZUnm+7qJ39QxI8ZUhrCD
/FDRS/ajxYm1vYgK4kEfwvENdvCCEP8nWw3XLqHzT01yeBXpwFH/sgGyih/zdeKf
BndzuyL9y0Er8ewXE44/dk5ZwY8NqQwYIBYQx4OC0GSePHbg53q+3OxeAAyRnwGD
2R1tRYXymc/332TzzfjSU3K8luRneoNxbk5HusPqZV8d/1SleFyHjGxdPMb3E85L
N24GziDatvBiK7UVgmUTCXzSfuViBrOB1FwCS/2JPNCt757KiZCj50DOiA0sbUgp
axXZX6T0l5+QVMgePQ59IyVewnQI5TaT+V27tqRyvIdVmTuqW3D/Hv4xUdfSzlKb
UZhEA/NkhN1YTsSGYpgCpFQZ/Pc7g+NHKXSyvPZWDQba3CIQSRv48vB6aJG/+jZ5
vQ1hA+9X9GT4vi7Xmb/vWOs+o8EZ+zrM4SOHtN1sDtjri55TxKuJKNqDuyWDU0fC
2ZeEBApbfddI+GBXPOkEmV81ogMqdmwIySPg2wuXlMxZOXXkM8dkUXkAW3gg9F3f
CoKD1/6b9K0/CgqYF5j63mWeJ6tBIG0hwV8awQzYlb0+VYwMkpUnAZEMpJvzTunz
zk72PPBF6PxbBE1sovLBzhVsoy2vOJrHGycETYdoNRCeEna3YATbA/w43P5hcPb4
zBoADuP1o21TIxVL10oHEFRxvj2yB+ThcNccrm2a2DpEyR8akOnEi0D/gGDLTeS3
Dp2tCPeVH5I2g+Cu6EYpznY38Y3Dj1VSA6nhEtSPXCvacnH2ZtsTX6MpPzXqDCxB
cMyJKNAA+B9fr98fNAS5T89myL4JcRbhzuooG1m6IiVRnceMkY/VihpiIpiEr/sy
fJ769yWcyWbIHvBpi54/Fq4LLyA3kOZbRgaHGgd40FnZcVw4LxpXSXRqa0NEvdwd
FqFlfGJ/ZWd+RJ8C/7MPQkJShW1pSfYlbhNiu7k2YruYlHeAuH4WzJi4lS2JjoTe
ktxgigGsq9bhVUGCetVKAytSO+Vsm6IGudDZNgD7vLHkHkS9z8fK3YkjOL9F+Got
kiIelJurWVmKjYVi4IKWanc3LUVY/+wZTTfyR6tqiqkikYTm8gffVs8trLece7UE
kFSS5FBXdqwECLkM3NSpY+Uyn2ZYhDPOdj5fu8uPBzZrZkkxCM4fSCFRB4Kwm+Fk
QnhsTTXlHfUHCkFA53M7n+DfdgIGtmpIz7elTk8jLdo7nIf7DgsbsLwBZYu27dXh
hZbP63kOzf2Kr53idg2liHvDtxKikbKixlvFF+jjfx7r3hvFQTCsEaRKn46bL2gZ
WTW+09zKoy22vAzYkzVIhpN3kyW1hM/YVlMRd9J1CPlA62xc7piWoH9M9oPFTy9N
DqfMEzjvHb5nb2aNm01hPbLmshwQFUtU0FdQzXjYmQyNZLfH5XK91deEHUih/OG/
EczRQJS3nMvl/M+b8XjYVh0B8MYQj03P6tsOZSS9+kTST794+ItetYaIkc3/I6f4
iInyzpuNEwdNx99da5Bnra5p5+3QfVJWQq9nnNUxQrunSVjiuvUcd972yvBor5cW
Ohk14PoKQJV/WwbLmf5i8ZsSxaA9mXVA721B9QO5fU7js67NXDStVixAL4HHQV6/
8KvcIXy9jvuPHuHN2aR0mnTZ3fgsHj68ZGuvU1JL8KZNUs7ie3/4d9pCwEkYQPno
Sa0oKaWpFfkxN8DAmLpRSpWbSzdqLHD4WbQOp6KG3lCZiP22N6JjDLuExaCwAnks
gQIfISovnQLyf2pCuQkQn6pqlfwkaWMYHEewF7iFzSi8/NRsf2X/XAfp7rtIbKA7
YzSTD/z2KIV7loDo2b+iQGeDxeucdVAp0izB+9um42wgF/hpsyPssTZAUG+HJi8a
LfSaLWHIp9ofh2ZxRScHiLqB30+s4T+iBAQUoTrGq1A0njfYE3ogmVkgGthARPdh
lyR3rRwslm2AL5qr3PhHS9I3+yIa0Ik06pSSe4G7W+LNTkFZUarzlYEytQKP3X5j
iwaA2MfxqEdAftWnanV+Ok6saEN1T0D2g+JtMDCtq7Yi5zMfAyQGdcCwsEX4f+56
+LbqMH0Q6yHHPkK4lX1gPZJtjsLmTTSsYoqJaAZ0C1USOXKntnOpQMQ/4RigiY0C
9A1QbUcHEccTOUtT8ZaV2yemQg+NH7Mqb/p/y6eoCwKOYYV2Q1K/CDF2uSt7mU4Y
Q2SQj9I/C19EKsNohQjFEKk7s9k+xBN5zW1lirotTdBhcYwk//fyDhmBgQYvfFp8
NP6kjHxMPBe1/HTg8BACP8ltuLHIdX3JWFeodoXF60dGu80/1hKyi7QC/+X1EF8u
XQedEoYtvxdB4gWW5dE/FU5EGUiKehHeAdYA7HEtycq5wD31siaBJX70Fg9v/KhD
cA8n8H6/St3/7KKXQvzErrJV9YiMR0ZMXyTZS7Nmbs2rMliSc0nbZL/O4KzfMIWB
PtVDfT5QgKAYzIbVF9W3BVbrRrxxJjNyR30JyHUCa3JFeZXW9nUEGb2MFrGPq3x9
NzWdRe837H25u8tK6KzWm5YyB+md2SDGSZHjLaqNu3FiEJCigYl2dIR9U4Fr8hsi
xhL0uDqbI1PeOPVW8xXsAb9rBnjSyMtk7enuQMhP4oBtfU28nqYSFnsfpuRxobJc
QppMM7P5CsBhZ0j4arKORTTURciGfZtRQBrS06RMULR17kEa81d2c5CyQl+v/aIT
pphNaPSTQDmcxxg3wQX6g3/sbVaRnaCThtLicMzh9hiPEeUneJc0f+axoe8iWzk4
XqnD0qdF+EQ+I7qcoTqagh9rUOrf7NCOymjXhNQ0W0PvnkpNThyvhfFmoKSkNJCj
qPtlL340NQvmVmmNh9l2dFe6rE6jKJWMBcJ0Q5UqTcDnJSzRfbtSWroyzO9FRNNH
J0+omQ/umPHqh9OgbW8TQlPVXAuNJnSegR/c1afBm+FoXMPHxS4lohmaP+eJjhfP
jxBv2fUwG5udZNP0V7gUFKbkii/MmqcZ+NzAN4UfCw39txBwIcdQNWGmP5nVJm26
52Sp8Vvk+cDIMKGdMBmgfpBndjDbM/8DNPFYVHXzrJ1mTrTEwUIljab/CPWV9+oi
y3B1oFus3EZBtnKzrXsiIWAmyn+20mSAZph6mQIfXnS9nD6TcEnqA32+PXFyvnN5
9WNkg67bwRtRCm8v3pOl0oTIwR0xbomDh53pQz6KSYmQDswSprDC2WHY/8N7DOL0
u6rAitcGPTJgjfLarBTOwNrEvEIMGa2eS1bQ42kBI/CUJ9tCOv5NaDxMv6ec5fNT
7LprCeaMuTa7jG5vrlElzh+mTiXrkCnUkjMYqK9z8rmwAe71S33jTSwaLSHGNSwP
3qXU3UcLKxwybg25srz4eFPoRMIoi0lnqb0UcTCBI0fNB7I+vualAmfUEvfjmnbs
KVZQcmaXV7q0r3jwjFRWdUTUbbXnWTEZjZsMOqTA0fEgufu/ebMqH5vnMMHu4+Nr
TFzagfxTFpeacsyRCrnu3pDIykUH9Dy3A4YCDsZxoj7EG18VtIMp2bDfG6AmmDVs
jfhPR3xIMKdZzSF/f5Npq8PA2AvJY/CRo8eAsXaaIaW+Sh9eaBrc+zefW0y7hf2D
/TcDaPH6LkeMFLBsZj1Ah8RWE1jH7dec89jpGqRLW5Svb6jo/UQ3bodDucPwJ2MJ
1OMnEgW+yGt0NVFkG6d2FgnvYsgtmlZFRCkD9zrj4Me/iex0Jane2AglkaIp1tzP
r/h0kMNvLGdz4RFSk/dVUBCXqMBlsNnSQhYxck7kSzAu7op2gBCa9QYZMJRCUuno
YCypQ1dkyotvCVmVYZiniijFAowkhFw4CLUoWdOy3+6iDU1FkOmKCQEjxsONscKp
ZJgLRMFBoaVfQa8VbOpoCX9RVb3XXB4831p10wyg1ibuIh+GiaHVaTBqtVZXkLSH
D2TVYNuqq0jhcdb2Kbo/hP/DHslc5EIawAat0xzL6sodJ+ESzTrX1fry0dcLM3HJ
sKlU9kTtdc0ExoGyuUI6+BsGG3jAq8Q8hIfsjXjO0yAdx1TG14BxhTqTmB6bGUlC
peezsDStDUu+xvb1BFtCdUqot/GMmfgo37PiZfECBSaET8mvPKlW9EJaAjk+0Zy/
4svxETSoksrLDu4kvn8Z9qE9WLlXXew4wKqXDKZNuzlKhN6J8kJC7D9tsAIuKfFE
ebHDyt0k1ubYf0XhG0hnbxv0iY4FNiOyou6GWANcxft0WyCBn20PZj0yVuot2fRD
kf4ZsCP7xL7bcksyfuh4TjNjCdTasgrLwaLRCWik9eN/IN6Y9+sYwvGA2ghANKFc
7x/lZ3LXQGnem1EWQQbIB1W052NqADao7iJBH1u4JXHRrCureKtPT3Zy/4JYKhnL
QxfESEhGhf0Stoap2zPVDLFCtABjHIKsNU3tMZmMGLczfO30nbMM3rvQK73Vw+fO
eeI2aQ0PzcH5LaMWM76XALx1JzWHB4JJoLoj7GVbzdMqaY1YarCQmZafFKYoU0Fe
9PoSIK7xHGC11YPnUr/33oHaM4Vt0C/WzMcux0jHDdzF9XIg9F/sppks3Gvpoi9j
4g1aLpdpERkZDWpEHQJi50ewqWeFZgqjwVO1X1oCYGiE99UOaAeMv9ZwpfzhxU2/
Tsij+j4vNIWXSmoAiq3838KKpSCO0MJDpAvRW+Pa6SeRay+mZMDdoDxIPAef+EL+
89r5Mm1BAYN24jD2DXa+CHO+h9Ggo9cJvEaayoohQRnT/45sOXvv7RsuPtFJVU2r
RPGwwHWamlpmWLooPf44PBU6/ug/IelMlSl6jf11tqjef6QanS2YrFq34rx5Ke59
9VvxiJa8AAGJRvRyUfFAaj7dXfQOke9EJSehvrtq3knnRvvegnbsM509QmMvaigo
HfPn4TLEXJwseKalfHvk/7WniQf0nNGuLPgonYlFIPYcjGAAQQ2DJga1cP8AbdxJ
EUxBsv56cFAtUcp1YcgzQbp0UQ0As423AadGkAIAUeC4Pqmb1waEoya/Xrjs2L7x
JnXaIQ4pEIdY8c0s5jZ16SBYiRkkyz8Un36JLB1bDdZhiRhaguHZd3E2xvSKawTA
Y/maSOh5xGwEb06/eyQLYNM9aorP+Mv7YxQ8EztNf9TD//wVJAnCsJbkMUH6HX0u
Ag0SPzIVLuRYJC93EIea8LP59pp4IjMyyzoE5kAUC8kto0N0AxxSI/tssRUBX5+x
rssJti4McJjE5QMsPrCAUhLTbMbe71AqpM09hulZJYWVExef+xLRRq50liqRANB7
jSmi2GfweCjPll0z5IsoKjA/1qZGeru8FhPjL6wOTqC53O+JiT0H223dDGbBmJng
tBx0ejJELO8ZJPiB5De5mbZHTjEaBSbyP6YiY+ceCaFEPngbVsG4uzZUVz3nFXl4
H9GR3UnWSo3KB9eK3v176NLrbQsBAlIfTbRVsyUpUgzBlXPeqqoVLm7rS51GEyDU
SxshZQ4NijG0jriDGSpWHpLIvqYJk9vJBE28PTA/n4NwjLs9ixJiHVXabKYBH73T
kn0birsbu2mEVpp+jQlW7X1i+G7sequ0BM9GPPH2kpbvEJ0sM2alQfRcvyhCqXFR
dqLdo/7BJ2n64FUZP50X2qzb4wW9by/uxtUKpm2urXNXaWU+Mklsn+cFZI+sdZXg
BPt0xFFkUTJ/qJMXbMav+BkioI/ibZTsVXS9oj2p4JX7gXv8ekZuduRJuZZYyj03
p21S7egj3GzirILvaPFXGHa9BqgDIzSyDM1NmnJATTcucp4FNT8Uj/TNypWF/NzC
9O1mKY3hVXbn8v22QfkdOLuLwxjUiYLKhMCUbBlv8K3StQvnHH1fE48e9IvAdF4a
UfbVrYcsroedInsq9TbZp3KiNYV7XV/9AOQG/5gmD00ie5UCdfUItoS7j4sdea0y
CROKO6WdnigOeSosXcsf/IBwmGP5W1XNkDwHOT264z2FfBRFMXZAOwWAM9jEFkzz
X2yxOQc1sICaPMv2gHC53UdEBqNgJA778hRlOQMgJlZVGAbGpv/UeaiO8fQpEMN6
98ucj/Y81rvHiprUXrn0pzmOfdppMeLmAL0jNYqoxAfPiC74yACSZ2pAGDEsr5M4
IkJjvEZxYIsuVPfrxXbWcZHZxOH8JGdKX+Jpe9zEABsyXEQ76ZGRuQzMclSwQclH
TYBx5F1Vxc5IZ8V420OxKh0IK3WtIP7xyayTOQkeVedcvwuYql6iCXP28GfpkMYo
uvSqCzbjR+E1UXK2vNqjjMw0UHxsnlxBzUGYUxbhaDkttigy6gw/tdyNqVRTwBGR
fAlwn3EvMlyTqv+hrx4iKItPgEmGlDNN1/HZCXBxDZdDt/D4SFPGMlfBiQRh1otB
j8SAX0FZ85k011OR0eIPnp4rCzbSWoW29KNbUfRcZj5iaf8Tox8un9lhyFDJ+6bR
6bzRJ8cTH+02Lx1NPENwLt5+y127BO6pcKhCLJgIj0CY6pGhu4fAPvzO8w0gPc0S
DfzumV/3OSTFwdcHAdsoej5uKqpb8HNbv8LffGofYT6P9QGwdz99NR6SVyyug0K6
QeP3FDTWy6u6ZHUy6hedBc7D2jOARNbKDzzpVbTmR07q6RNKHea9n28usoRtVKBp
RzYDQAYGDSrKS7yN+UjDMGc5l/0ljzwUeTyPgxM9q8oWYpLbg5TtExUTr0NsP2zv
k4sv3kuk1aZY8Pgm+B5kZ6xOhmwERRY9skR+dldBmqZvSweyqGnah1iw+XlU6Bql
5kX4BBd3QETtGkA169e5iess4MsAz6WQ5JbsYZ7vwYEM0UVJcnhTOxKYQihMC7dO
r7Ql9eqSRgx4/3uYqxSFvz0gRxUNnOdsYpRamR0PcbtpKrXGK+AoAIH+dAml5zpi
ffBVL5amb/bc2kG7CHLDZ5PIfT7OUWlq+6xcrORGVnFj27XsMwUWsLd29srfJwXR
gXuCZ+sSqbB7LtlCUI6KMuTiJ42CEFLMIAZ/+Bw0jH3YP5JdO2+Umd2p8NDUmR4U
OkSlWWNQnBrMAjMBGqZMVRbzAfMETgGJ6ao84CYMgtYFEMz+GkcYJe78O6NSjbEN
7PXMMCqhJ9M0jx6xUD2kMiZtuJ7VH8d4HimZl6QTnifyjtAZUj25nwZr5gj6ICTr
BcxbySAhL73FUkqU80q3cPxnf6ZbPGinR3kjZBslfmN9KBfhw77f6Pf4Lj+g0asX
Rsc/uJouSl648P/Ct5UC3Q3I5tMs28+lfcnK/L73jat+lqLx3oYVSZjbgE5SC0/u
9GewEARzsvqQRbtpYGrdVbdtl0xzENcc9+czfgCSZfe2hrAVi6JTbwXDJtsso4kh
Cd/aJoWTZDXWlzZE2gRB89AXwMJs2o8VTYITGKiJ99P1VmyLJz5K1C8fdlXb5Plg
Ckok7JGaW1967eA6+S9o+VHssmky8F6oVouUwKCTKuTchVKaEMTTi5viDA0CcsTL
xIZ9K+vM0Ta7mbqXGjNRJm4I0DUP62nLw19M8K3EUt5zSKHoAcKlKGZ3PPeYF/xT
9w4DZqOexH3LAbsRxStS7ZtusO4SAt9L8UWjPVTDS1JX6sCNx7OEVPDorwAnJ2fd
brnxerEeWGvpF1+UxqT+2SHeDIojNnDhix2MH90lWOHGsoW5uuJKmmFJbxiXVwgV
AAVxClQw+5Q9wrOhmZMo+aqgBZXM1scxV4Qj/Tvrxrer2FAiUUDjZZ6AkH1jQSwk
La+6+EgOp/98DpVCJJcQz73BO8mwoHFMn1s4kVY4GwrBfk5GQKBE8bMreIfDaBn1
C3iV3iLUz4mmrbpcZagJeZ/mCWq1FlweQNtbCS6Cn0/A0AcW22nANrnXKno3RLp+
/VQICzzB9Tm27Qh/iFTLP45duD9U/IK4eHIwgR0cVKberuC7rg/V4BMNdrmDt+TN
ryqRHFjbn0hgyFLt9RqMv1tTR5QhAV/dCcYx6qCtFA49mF+pVvIDsbPmzXLWshtz
FS20bxS0y4f/yyu5uluj3zA/fp+Zx0RtncyGXSjkXGoWVKoLKH3lRx1W7cL2o0dO
8B8rYwg7zO6IlMXVAhhFLgSxvNXpZ9h0MkO6/tSPwo7W9mPMMZcIfRyVzi6YOllD
4RpnzJgh4SxrgBSJsXV1MNNUYB0HztiiF20UvMK0Im7dTmePYPCHv2f3TJmJqAVH
XYtAn0tsUtUvi3r3Ax3cmtn0w8ASkjPIdB+1B1K7DjyI6LmI13c4S2idaMy0jbGg
u3FJvYsB7vW6c0kwgWN7befZDDs6aU2zyrDdi1ABg0obHAxooWDSw8E/7HlRSE72
9m3d/PqRpER2J0kUOuyY9o/+g8YCRtM988SUDZUzpWUPNjdFLIIYnPd5ZaeQ2wQp
JKJ+5sTN+jdMJq7FZeN3sWv9dkZxWaAYVE50g40vYMwlT2eTuUniVHcsrfzR/iS+
KiBGrW25hVrcdUoleSGNrNIizLkDtApvX3SqxqoBSz3F68VskKdq+tYNA5OpyLEn
lozenpbcHcHw5XNpkBJh4s6mTqMYQpecb2L/DYi+vLoSWXS7svWj23yMqy58CuYM
d/wuHvWm86wiEVSvej8u8YqAVnmlexqlCFSPJ9AgrO4GO4+3VkB/blIqLGvamLIO
LUi2JivQicIOr8ua3zjxNMxO1wQHTQ8ir9e1+CqpYOtM4lNEGGsv8NFIH3oVB5O0
9723oT6pknZnJ9SokeNcteUxk3916TMtEgxDHbGW5+7O85L0fuOurRWVk0YsBq/I
8YSDvYewbZjxRps4Xi2D9ZnREHczW5Otzu2Qt9r6wDDxdc3JbXjzImK4Mia+IHYk
SRRg/8SIZfmAxMRuioL96YP3BrJMYiaGgf/LcX8wKLXRjML8vYmaIvpeQdWlBGuM
ZNrxd+DU0vPJFC2KhmItSmxuIAaBfcHbTNg9PWDGQWjQV/DoSyPkqUqWR+yugDXV
z55yhhoI4TIPHV1TUNZ0pz3NasO7s/4vJXruistjvM+0MHwJmiPWctgmeDGHCr4F
q3Nw3PBETFuMs6oj5+bB9haJp/FVtRPNGoxv8eK9H8zzqZLkO3oJgS4UiBpTxBb9
BvOvhhgQEo5dk1hcqh9i6dVob8IYofc3S0rWviytbQbOhVrVJwDKZZzrbdrG+29V
Sdj684B7O5u+SJDnQ+5A5t4W4XHRThbPbUXuajauSaZzoZo/bKY60/NUNfu/eEyp
PLNOLhP0RhtyMJquXeIWXX9NXutg1FAN8fCBBPjUVw3lnqMlalBdh0lOqPpjvTpg
yDo4vxa2g4dMbfwI58bQMCno40Y+DbPSgt22farKwxgh8ppu/SkB1UJX5fkzpDT4
RPZFP8jUl7M2yvjgnEVn5BXdiK+Lk3s1IsQfcjtqUiUMKfI49Sf6TBz7DqC/SU00
5pmWo8YmGvDlS6KVWa7C/aYw3l0tgfZKAP0xjmRuZsINfM2iFX5BCQTLG9fa9XG7
tcXBmc4nZONWI/Z36NVo7eXlg9t4yxG+MaBnC8y8JxpWdR19gKRlEdjP64ExlDwo
922mLosaUfnbUwS3mmAewBitbquyvfpj+owDkEu9IV9ZSupGyyP5D084Y95xnGaS
aYUmbNDR+Oo28FzFyJnvYpERWW7/uAF6jJnUzj3URADtZY+DD0ZXUHqi8uWpeJHN
Unf1A4Z4vdWVTNfmgZVtSpmOyYFLxUsEGxTJOzgLPj+5uAzC7+innIM9Suf9vEKx
KPnc1XrtX0l4x5SF2ttnsKtLcbmCD6MZ5KJgTllsWtHBEzI0W97yVieMzx7SH9Ex
Sky1FkoxEUG560KsD7ugbQ30cAZrZu1hVEfVnzturqo74x2CA3ykuC8r7Dx/JwYz
o/ZpZuRVziNG5IsRx3pY3BiTgu1b+yo5LCen9YNrAAmy/Dss6tOdlJIbQVC61ocZ
vGHiC+2gSv/WkH6R++feFkL8VppwL4Cr+ZfjNHh5mxsJUujqg0wuGhAOX6QPO8g3
JlQvay6i8M3vyXclRftx9ImbgnuFFsZpHIh57/mV00hEjrvrOGKLcqqYbIj7fRE9
PeQFL7Ps4e5qdIlrYikbmIQWbFREV+HqU6Gill+eP/r+hRNOEs02ep2+pR8tAcLu
1QWpFRNkxabwItF6bV/yRgQGbEFMtgSd+Fz7DPSpV9oQFMGQwbAJN/oMIXDjyW3k
VUGq3Zwbx5EN5Dzj/uj0euV5pVJj4G8+7IH+mGyYFkOvmK3KB5B3Bsu0LVzvqaqj
bD29kjNNaqm42gZTakrCh23d5UwmcCJnpC7aKzr3nRmZ+02cC9FR2IRURSAzJQUd
sK43nWBvToXWrlxqhF9AdQ==
`protect END_PROTECTED
