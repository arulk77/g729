`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
jWrOEt12/3WGVXqNeuatBM8L9HCYo2NP1yCHodeBIiRj5PEhgkL62tgsMlq2Ow4y
enyMbAzLqXCYHLdmCxZ/SVWsO7tfUcIul4z4JKktJ2TtaYptAZwv2GQgJ8uKNMdU
RoDMZlg3jnl7xJBNQx0ovuQzu4YRzJ0dnFUXNyxCCnenYBXfp+f5HTHPVmph3zin
blu57hBWwNsiO+/++qzvAumPqBCRuXk2M87rv+akrn7y2Bw3cZKoSsMFpfvPgsyC
Bcf+b77h2CWXj75Dt7n9wHr8/WcnlgP1kZjCiEdWEyDDKhFUBPR1Y5rXgMsr0BGC
vnjTP2QARyngxkvw9UNtJLgbUQCIA+ndJ1lvH7gfpPKCRp0Kn6hNTio7zjIBRiKO
XrhJwPGzwOkOONzDyu8dUi6gbGFS1WQJvL9/tl3W7IzABl4OhCQw4S9tee3iug4l
duBluDZQ019zoFfFBPy0gfOtN9s4nvH1/6F8wqoO604urAq/AhnMmkO3AS7/i369
btuYB7ZbY3vy2Yrc4vATAUhnAVLXLyAqmMRnmcjcyJiuVg8Xg34Ajtp0l8kR42aC
Ik0oT3LzA1bP1A5UE/cOKVzMsw5RGY4udkKNNe0Y/isx96B2OJw6Mcjxe5kZX/KQ
OIBY2P464TCX7onNafrR8ExaG2nFkNF+U41XXtQHfOYpSBoTyc1KBo0PYid5f10u
nayVmMdb4rNxQxm9bmD3zNNbFPvI/GHqeghFgYVJzqd0DbCvphm7tGWu+GiHVTKV
zZLfkLpXZVRWkaro8l5Xdc6qJswTULz5PP2eXFJRokPS2jgCoGeaEFYRne4HAiIA
fPx0tKC+5sh4RTv+aOZ1Xw/NDc6LtbF57Qlfwf9+35ZkLWiHjnL+aq8lXuTTeRcU
c1GFF0L5GeCPfbu8ObtyI90wjxxaBQGKI9CnIoxtLMnAcnOqVVKUbQ2NMsMjHOpX
xNyt9eVOw1AKlBd7xlh1yVMa4oATai4byH/3dSz9F4F/mrSBhwUf6728tU3LJRQI
cl0WMnfZJ9LT6Ezpc2leGx3rsGS9a+vi4nIbquaCTBM2LZOy5tZdExZ0zFoCoZ5c
qB/pClUD7+uNW7jc8VHkeB02vZdq5LGGmU7rvcK8wt2xb3Ftc1EqrZvxMqsfLDFz
htEWh+d0qSArTsFuAddwdcFR76ny4XYGXxpaelyt7pSsSLF7BzgXkvksosd7aGZ6
MDY1ElOh//urP+0RGnk5gH0q0PbWRfmGBzl8DjcUHwyPqRM0RVC/bzuAsHHFUIaq
UchA1dei45YjEORV14KHEVWL8okkxZ6VwFkLqRAh9irJK7Z1uo5lIhXGYg0JNGvM
K67VQl5rQJBAmzZiSwlOAEShRvKg9iilJ+YVpiXk5YxjhSb4KBBTCwWhd7YwKx1d
4AD+nyB/Vgyu4NphMBU9SApCndxoBD1YjBS8M0crH6O8rLtftZbdXrD9qYAQoW3h
Xh8BcoMPrTQxnAOd+jRn/aQ3zOqt9m2QQakvV7fDbyKY3WzUARLxGx9EunTrkH1E
PnTdgcFjQK22xoF66PlsoheedWN19jKOg/ESYonbI7XC5vFHTFnps3HR7o4hUnBf
2gYfGjEUgH9XtUW0K6sSYmQFQZR6lvc6RUrYUNMRw1Lx+ydUfTEKeVSkpa/xaSC+
1OvQEyfjiJLssxFywVBUj/xpFjBCadEhPiAqfYcrhHayCyKeKYC+6lMGJP44di4w
Na3EavuoSK1JGUzg7R+rddBAaE2fopybUuR/C2TX/XjUAUrgHYpMlnV/SKnA5TK+
3Cvout1sA2aw1y5eCXEz5b9dmgwXN/ql6TVQBsF1WMYa6LfW0NO+k73SFxt8EOd1
Woq+gvmUHqV51QbshWuBSZ89mEel8NIroS+hRYcYj4oNP6aXqlCYx6WfTfeOWMT+
Pzz0BbzAdIDd3SRzzITMA+p5LOycXVkTUeLaJBLsqaMkS8WDzz6W0/lGUIIoCpv1
Z/3r8qJxOy/GfJ4VtDJ9dOh2fezuf+tpMNM7dkxVQCsl1yOFT5I28P2HNXc/bOvX
MMvV+y/3LUmLZURuj8pD1O8eh2EGqMQElHt8dwVLws/xq/4jkKXTbB3qkXWcAKCq
Wa51z39FPNYp3e5onU3gOdzWSN+WNnSpt53fAf72jS7si1vnAEKWq/F2f0nh0PgK
`protect END_PROTECTED
