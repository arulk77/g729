`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAdTde9D7tILS8XUmqX8D/Le2bS11KEgYETW+uCWu/q2s
72eeXGtPcgOaAe6wCFQkkyGNwWtO6CopPYI+A+mg9xqgKutTwchb4sIP6As2dahR
IvnTUeX70nkz/pAR3DooRUFdrrLFsBmTM6F6JuZSwmaYzmc33p7J6Fj+8OflNGiV
+kBUPYmkz6OLLgjMgaEm/DxNJYQXOLB0gx1y1RhCwgJid/gDrILl+fv1PZ0AElEY
zhxJgCa/3xn264MjcCFSiysjBtn0t/n3Qrj/Qwc5wOgnaXpEiA3z4iCQn7lSohJ7
1sevuG5i/4s/NnNeQEf/ouKjhJNe/s+uYnEZDUZnPOp5Dh4Ej5gQScYzZAR5hgvq
eNlPgxUwRmHaQ+p+gVwNKu5dx24dub5278EP57tjWOBbASnCA/I4N5n7ddNQMxMr
a35s9G3uPfg2o4Y/sW3PTtKaLPfqOPOGL2zcuMUKGH5GjIUsYpA96H5q8vVI1J1D
XCMUlNtmtIfd2TnVoOU843o8VDmZ8r/cTxumfpL3wjtv4+us4a21bg2F530AmLMt
NG7JWHFAKPRsd6SXZInzHFq/U1R/3z/SW7SbXNTOZ43wn9zxmTODC5SvqtIdJjBB
XDPFvv6HHWOPIn2quBXzFjEZCg1E7cMCD54BW13slTrthxMg7PibnqzyHKMXPpDZ
V+3qmMsjb23CfFXeZ1vvTc63ta0ULgJAf89MHNd5WFyv/tFyZ3mtmGG8vApHSc85
CV+5KrI5KLrlBYaf07dMv0Qs+nxUHfym2uXpOraJ+z8K/IQJal0cNOUzMSE0/Cdp
E4JFc5q0MPTX5bg6w01tHci1y+rFylQiHeureh5u4vhxC0dGc9zuWnaDr74RPtKc
aSNsUcpFyjMFsBtymE34MOZZanrvbafyKvOJ+Lv0ZRkRzZ/yL3NfBTy4Kz/G3utj
q0rEr2144BmSUhJnLmnKjWedEdzihF+gZqVTH/RT2C/aucg2r1RLy2QQrJRARkPu
cQFxvNT+iK0jicnUbP7dNfJxcw6j65Sf8JIaRR74sUD1+bob4Uuhb+X9wYuKe5VU
7ecR36u5GBqrAcelPnj8TebNawM+MyiGjB02y3M/cT7PbLl6r4+4SvrQuA4Sr776
P3xiwuOgm6Ene/eb4NRd2EiIHbIUCd/4xR2JTQH+kkgILhTOvpSaQ+sNt8MAYnkM
kic6JM95lVRuRKZBY/PM2p83GW/Umh0K8QNso2ZHfo0fJnS6wqdtZFSKiU7vVUtx
yOEHBwFyhlfQWqX9mbel6b1LqGCJ/w6144+HoZ/jWa83l1SHK+7y+AQHXGYQl7hf
RI52GlWAiV3/I3MhoML/hCQjk9Vhi/jZSvblkIhFzJ3QEWi2uHrMJjjoSUmI2HPQ
FMghcm1K0/k44ZXVoUiq3mkZSNhXHcpVgln0JhOeKSFx5QsKncUtN1zbBLe0de2X
R4PwCoPYP7PWqf2CF/KmTN8Je6bOH55oNvIMe1QaiPJHZBt9CA5BhYx0B3+ag6uV
aaS5klirebohI/3jNhpewWT+gQGz3Mn+qmwASCRnuWXNwmQg/is4V9m+ZZUj311C
f07tXsFL8nr907G3m9jSlW+aYihs0zKf5PnWcYPDApao+MOsM3IcI3aY37wLbPJl
kVAJxRG1NAFA0QLV2Py/mWt+Zpy7CJbQiucQmqPW8ScVDREFVvRSX5pbl57zTktW
Tro44AtkFI96vBiWkpkktGLgKy1MhAcRd27Hc9fAOi3OzPST5UG9rTudlMeHAUrc
SepCVrygao+XLp3pgFoWvVYq83Jj5J9ONZ+MRTNIt1kqCO6sekJu63dyGVVPss5k
8SUg3YyrNC1y3Kz6qVw6pwVIN9z1P0nU8mqQSbU62y09WFiYiY/1RAmgBJrLOnIc
lfco+IuLFaIkDNe9zYD9o6mbKUBpZVKHgOholoWnJj/+Z7znZ9fKe2aXBFmXC6l3
g0yfvKAZhu1u1mm7zSAU/pF6RgGFayxgBjUg8tHrQPuk584DgVBAfj46GVMvQyvY
OXUAqDYNb2Xk7LHN4DgHlxvikX0eI8MaT7A5e9bGHvI2gIsVyzgFLjRoauImrmhL
gHUlcByPrYKcjiiH08L+fxyXxIpMcDVvwZlJ7+4FS67CVoff6bodoOcKHd79mL/W
Y+grG2kMrrcC/6BPlyJDIbCD4ev1snYYiESHqh3CUUStZ2kB2yR6giUHywbnZb0L
bZRz2LP8iTzlCElc7jQ3wHxtddIyPKbq8RQzIdE+aELOxa9c/egQUnezrKnZUXJx
U0f3qRt8BhrAPPIBtFzhQbP+iRS3Mu3ZLtnwlaynelRbHueg0VDsUktLqsffdqF8
bWlSdH9bh1yrwspX39bqZ3dzCJu5AP1zpu+0xPLBdLOUgZkQpSpxOA27iv0i9rpQ
Y58GM1jtaAixFGD6j1oEgpFbm7J615BnXCAn4K94E59dB+6L6jqFFgz3S2BkzHa1
gcCSM4P1ByAI1nZj1y0l/GAF8+An5Z4EJgxisQp03AEGWEvqWP4wAcZDsTBRLZds
mTtPUZmZYgeDMvMb3SW8n3FmQi7E+qOrsI21BWj9Rajkk7Z5f0iiWnwsTqbdoVjn
Vd9TcnMvsUf+8AZXXhRlrWgFePNDifDThogCr4Rl/69qkdeBBXllUrC7ZrfM0EyU
87/E/KPR2AZTM9WKTDZQ+2Fd/4/qB6oCuaWYV/vS6Q+w2YYvilLFD8cqEiEtgNzp
PHbJ6e7y114pwg0wbS3CXuiDa7R1Ua5OZDpI5G+mIomllDQr5hvUFMT9CyROtHQF
EI1f7ofeC2acD5FVtgEPwF1ywnGQnFOScp+n31o8d83+ekf4nTGZPPjXeEpv+DVl
ahXnmaqWK5XvEOdJlET4adDaSnIaN2vZyFeACnzFeqf0kYf2MRsRCo1P5EGsFVNy
z7jPJXO2WSngUhLLQ6aMK2nn5VbreFqMP0N/h1xhF+T0CDLlFEKFHfR8Sew+jYD2
2SWB2lZYdoVu38h9T2+ZyzsjsmTovwtiWALm7K2PPqh9MGNFfPU9hzRuhTiqcG9Z
f+WuGkAtZ81eGx1T3eSFesHCjh8Xc3gwH8Yb/pM/NACHKDSt5NSCxBqSEwoihn1U
g+utZURX104IKFRXZMxSnCsEZD+aS/66aopssfdp3LJBMIXTT6c4Dxev356PVTwd
YrwZfnQoKMUS60Cf4BvX8cGF293zX8cCvhsMElvmTxfbyQmRp1LijpMXScy+T9P9
+E4On5txmtB4tWOpdP4NT5WAbNWuHduf3Xex96TsNXtT8shzRPGupnUSEXT6a0gt
/bGuH027rDA6Sx/toY0QMX4wj4ml408/PGAgjjFR35gYcsJ/V6+ghbRIsQz/KxPj
f3YgJQRv2js65GUgOsnd5Mzk1cgJRMP0zouq+UUJtPp3Ts6U1hFTTBemgM4d4ucs
EL956Lsjpyc9KNY5eslajGowap9zqLQFii3JRsVClFa+k5ZDW81QOlmgn5ctJfyv
DC/Yc++ScLhTnfutRYLInDScA8kz9tLR5QumkChRH6nuXmhF3nDIRjiV2Xh28zT0
JntMZkAvmtL7YBVLs5G8knrcMUM7ENByqIQQXxYkKvyt2odH9m2kVpc+0XTncQdl
V3Opdm3zOrjvto7+vd50WCVNgVDKLhl4nrK7+NmImRqoIzA0ktfFcJ8qtP9DMIJa
hOHi3J59LPx8y+ACfxaLNHzFja3RK1iKNn3qh0YFlTQQ586u2Czg+Ey2huzSBkBG
jNrMFernqSgy6chrZ1HbwsbjlJLk9G/KOKlwldfp0A6LEArsf/vAtCFZnYdCZW/C
452iq5FSaXW0/nQ0RI/UzarvCFQ2fyhu6/NdsAHGoJF9CwYSHlGXoSDuPcvB71ab
bd0hY1MCj5IOTI6uT27LI0eaawpOFmc6A8ZpYtow+WtNxmKWnFRy5oBVw1IYhzzK
sOjUzBLItyoPe5u495mkJwRcCfUfzaIHUwsPJ2XgG/L86YoLhk/6eK0fDruFy+df
o15saUpOwj1hrfJbWj0huyQ0ycyjzNxA+coK/oUAlpEUnkR4IuMDqY4ZXwy6O5o5
hn6KliR2BxdNcxw0pdadaPVol/XY2bZCtFsR+o0V8gdihsFGLJSW9nlTuMWmVUaE
hoMpe+lmyy5m5rSAUDfxqU4R3PohYO+39PGZLK6426HPzp+lXkEWl9SYdT9Pqhhf
HCepyarerp9jgWuWRQ3LaX0bhghhR0BmXSmrDzMIBmgs8C2EI5ZcE8vkOUDkOpGb
vOROyxyhzBdf/JYz6HHV1L9gkhVb7euTbCGXGIjBxOAMiZc5lvy2e3j6ZX2nnrLc
q1ulHh1yKURaw+nI0uNb8/WLGW8lF8qeUhdYbJCn/Wz8apDn11B40V/EZwVbntGX
m8Rm6fCpZqmh7CofGTl2MCY7974X7PArQ0K4AKYc6zVF/z3zY3xmikkQ4pPEgAtL
74+Nk9NW8AkaSf8LirN5rTAUiuw9cG8xq6lrI7fRt9Q/6qGqqmK76MUmWCsOmiLW
KGdfExPYVB4GZC2+fGJvPVP9VwC2gJxF27UG2I1ZHtHqug6/+RQTxKmQkHdgLkJx
FEquE1Dyy9SDoVx+4QwCA4Gd2wZhpo3seNc21YQ92XpeKV+9tWI8sBEwaNUYiTBD
FNyCbxeB79kL1s0LRSApcuft745OW13QrzZTbI9X78kU/usMNb6YV5DQeTykrHOR
KVRYLZ1LBUrPVovMjrf2rVFh0GE6BExpoI93NEUKqRkHeIPUvzwyvwTzjxm3c3eF
S1gXP2Wwl2uTYq95gjTdylA5zSM1FKNT6YPL5IrX1IHlrGSoAsSJHu8yEPLhTqgX
1xTUWFr8dz2O1+nwS6gUmywThCc7ANa4JBUe9Hr8V274dVbx80HDVdbQ9s4TcK3T
S29noShDgr0VWxpaepBC8U+GmvT4t+wbAm6uHEGP3QUhS8Y/roIvAZbQ53+8wsRp
8bgiefUtDZIgKPItkl8ej9feZhcg55FwN4QVGMsXG0EOBeKsqlvXEwhrcvM0iigJ
tD7VhJrLcXMmkc9/Tb3HebnYAJc0aYCUZFyJ1M8+N/CcbPOgE6dHr1WvFv+ndzTp
+H2hLjRoc3wp5yKpNJbEI4rYO0m7aoZ9t43L+QqUjF980WvIt31RvIpC9wwLSnA+
cZzQI88VvfMnEm36+v/XhEgsp3d0VQWCbXHsN/zYjh3cJETIFfwtrF702ixxO4yG
ylxqlZQlka8/9vbfs85bF5RlUrwtShxe3cVsUo9sYvuDAodNYoIrP9xQ8X83q1eX
HOOGnCeVr+QdW754jq6MHBDN7iwNJrefIwhgdXi1+lEWgH9MYyAJsZZDbq8ytZ0Z
LO9DovHT7ueilhckiBWe+RoCfigJgCewHHqQ+XhqRMnCpSbGLM5Yc7IFLhGMGs63
wxE+vsbl157cb1KzsmTP22bmINAzwPkKuM2y+pvHeI/uY3nXO0DKiK+GnWYKxqAE
KAE7B48u8hzXahQ1YG3Yz95DSrin8tosvLAOMCNHOXHg55QvLLImVloKjxHjiEND
1e8TTGowj1hhUrTsOGTaT/GAbd6NYx+pvEVSa5CFBFHQvzxcfGJLt6FIOpxiAUGy
HuHqFoqf5WQOdMimrmiYRrSi4LEvqgAe4aCVZX7wAezJVdK3WOvGPrm2LVR9buwM
BzUwxfuafP+WndaSFAst5KuauCAfcZeZP+jOPKGdD6GANa5BYxwOdCFTrN2AyDmh
zD7AIEKiNQDAYju9y5PhBX2aqspAM7vuXo8B7T59ZLoiJYyndbYdkEGwuDypSlq0
XJeGIVhTKofNcgJl71V6VXsW20A0MqKGSovs22tukRJlel/ntQMKnwKrN76qfQVa
7QUcyPCrIYoILmH8lmhHSPZ8qOQDeOdWUmSPAvLSlmE+sOiMh1ZIRC5iehF5ffGy
Pkz6b7bTT0GwKI5XxEAD7mnF48yiSjA0gfC0bZxyRtYKQHYGNQgHqouobCoVOfpg
vR/XsaaGBIiBNyF7tyHEbusVf7VZk+TplSOgYeVgDJfW8BsuEWaZydgEazhhAtJs
j8qCntjV4Lfn5Umo1BXvHHfdAbG9L09YSw/Q6hhACqni7Pg7evx2F+NzgGAbcAq0
w0WnN1nOFEFUmF6vZNPBla0QCea6vV9ylRIvNiZVIDCk8HR+CAEfc+lgTt6c/vU+
Q1uH0g8WLCMGPdH8tOk9qMgma6H/jwjbUjzAAG7xSdF08nW6+jZvBpMOEFI+kvmQ
NIDjkQ365Hn4ZvO0Mgf5TwOP8BgloaRLqC8gCl+4MWk=
`protect END_PROTECTED
