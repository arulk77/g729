`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN8lpX/HYfkdptE9//pJTZMlxy1Vxdeu+ElebqbcQKnRj
hM/L2fVECt75UHwIUaTLGIYvpYqXWSRIBGQlQ+Djynd87n9cCiLSqFLzVdPWgNJc
Sk0+R2nGQ/K5wQ14Ce+wOVWvbEuox2C2rxrwOxttJH1m5keye6XoR8hz5fZG+pG1
WJuW7YvCVTBIiw6YLNMhM0YR96+E4SEsrCXC4LIZ2/2Ech/yWrMOQiviSDKbPOra
qwiiNLNAfcBElSL5X34FObI+AcH/eoUo3R2WfiS2IvZjrmwFZdCDTPizdraW9/R2
LOIRtKM2wRixXW+/vyDEKl0lGbaZVcAmbg7vgNReqKcvj9EfwKSq6q6xbXGJxxp1
+G0hDeiibgxqQEJcgVor15X5YdvqXKrVDgOxHsXznm51ST5dwgAubRbp7hkCQp6P
LcQpW3AGbhDDjCSi2xmtyStRcHDc9p/0UUi8WBTQrQCPx6eR8Rb0FZKkKnag5JbK
v73iFn5HWM82uo7o1iaOBQV5YYQ+9qd4QcNuwPmb9fLMrkMbo0Js9DDY09Vvri24
ynGh2tmkHSxMouxn9kC9LnuPOH15p1pKxzLaSdfcBX6Art2YkPULBoq0HbNj0UNm
9IbQ5H2BXAIQSnxs2eCpd3h2o8Zfew3s7liH7a2ldQI=
`protect END_PROTECTED
