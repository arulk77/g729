`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ6ePP5lKnYlw0gAsiEFYwXThPA2zdTp+HxNk/KIP8ks
mS3lh1orgLcjuwu8jwIDnfRyYY5dU2qsTyPQtPNAU1m1w0mL16ssFH8Ao7ljhEyx
gBV5GfBqAsG++37MqltMAXaTkUclcV1QWjm+ikVQIZZ3Q8PcivFvaQTb393vVU0E
nQGvxw+pNbc9/ODVAz6UXJPNmAPsQiz+BkZ/523hAHuhAp8+VHm8tdo76x64DqSX
XwhJIhH3TaYfnK0zhdYiYwBTywi4O2FlGycIqg7BE8sprbbkyKq5aCc0kCefr+24
55iPVPxUfYQKf6hRlRqqp/hqm+WEcmtx6RFkfvfFNuBdKr421pzrEMPYD1qFHdv/
njZGkxD6eRpFxVFYyv9VQhAz9jELkLCb/oa6r4UA2lN0brPVO0A+LEC8+PJ8Qz7/
VyqcnvH5ytFOggUoYalmsCeO5YIITSh6t9reT2BYTs3+7EGFoIWjwCMiGzi2AVkX
aZLVsC8D/SFz0RneZCex1+95FhkvOGMgMAPFAmqUsXvAvz7dEqqRO3FuskL8fdJM
`protect END_PROTECTED
