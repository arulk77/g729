`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
TBdzT+sNg2k7RcYE964ME1+D/g0aMgCK0eEM9d+IZmIgNLJYlAaRymvr0FncZdQh
cWZNfdQ2XOlhBRmsG2NPx8j6DN4bnRXgmG1efKfARFQGSoW8sHBJrNTp51XWuRDg
/W3zvAty3OehJatlvQf3CPTMcFSEIb4JCqhw5Rf7aSaofjgwnBW2ZKN+AVIKG9Wx
gntG4aBLTm1Oi57ARXpc7BZpl2KsKXTzpkXP946pr/MY8PVYuKdCm8ByG2PKdGoJ
9cuK2HrtnOJ6iv6SsgV3jq3PPhmWVhCeKoDyoY6pMCBob2MFoYQLEcPWLtzRPPfV
jQkhUWJqd8O+dh7O7G6zoaNJkeKw9C2cyAF/h6jnEtG8bMKM4cPANSnXUrB8DhKT
RbjBUtiVwFo7IUG0KPqCMATI7mZYi+cEeL/vVKxVn8c=
`protect END_PROTECTED
