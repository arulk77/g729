`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAHfaOtudEyaA3sKGiXO/UIoT+FdxlVscUQHdNmUDYGs
SsKTakA7q5oTNj3QlNS/P6ius2u7OgBXJY3hEwqC8Ipg9U9F0d9tfmWcsZ6A78vI
+DSlceX2RdzY3q3kSKm9ghujs4ZEL3ibyjFI4m7xTuHcrO/UGg1VOujlmUZ7yIU3
/i428LScb/4YeIWr+KJ0G//BaRaTyqPO0ucHHrXG0rY2kit+00xuJ87N806LCvpP
Di2o+DpLncAfoMju/MwPr52Op3h7aHG24krc8KvbRxM34K83wGOmm9ATtyze9ScC
7Y6uqPVX76HJYg05gD9qNvAFeWcGhmaRhgvVn0YM31LqQoth8nTL9PYJNmTdTB3Q
P99456trckoDm++sjupzAQw5KJgIpw3+51zspESA6bJZ7FoWyr+vvsE/8U389mnE
A+xrpxTB7z7Mg5G4/xnXxXwv2XEHO6XyxnD21Jp4c3S5xM6YLTxHhrC0empAXI+y
QYODXoNL9LwhjgQcZzXNjm/ZYAzeciUQ9RbBpzG2XR6xE7PjQ1GPUCgxq/LGZwCK
sNJ9jGzfuR/ANs7vbsWZFuhjv1lGRJo8rxGOAJMvVTeeiILA79DM3rYAr+d6UQ/e
mgTkFYx27dosG0++RLGF3KPSGcr/rrkGMb11XPz4In/GyrGl1/5466o1Gt1hh0kh
9IYcdznJ7vDKB0H/eVY2Sa6rPkwgcCGZmUd1tGz2AXhRakrkTBGzYAIe6wPfB+L8
U/qxhT48Wxx04523527GxS6wMrSLBBiVYhGhkU0ReQq5tyFOYP0ZH6+E+lShfdEd
rZW6re2oILMTUxmq2Ck6ozMzAaXSwq/swHVFpS2peEiitDtUKcow8eZ4t6R41CdE
Ek2A49PGVC/YoEz7b8icjQYy3jpf+8CDYc6/dE7L17R7Ui2V6XiZ/js4EKZte1HI
v/PzFkfm0xI0ltp6hrTisrYH2L4jR9vtiLJVHEHtSdT5sPH2ZW6eFpOVpDokcat9
6QIcqrk7iJ2YRy7FfuOMoP387MctzOPIJYnmnbWr1R8ZHzeoxyypVsueA4G/mmwe
K1AGX2ohNNb3u+FJbuhHUF3Q1i9S3T3d84u+U7F7usPvHYoD4EN/EZq5dpnRUlCU
Qmrr/9I6yPystyLJOsx8Zp84df7UtPx7YCRGWRBSW4CoDInUtrmMyxJtIxqJlE+L
MYGzn647Jc+NLqFTMiubLk/WRKDOen5ek10/oLqzbKuG1/X9E9ofwIg1H+uEFQBY
bkjwETvwLHLdlnSWyHH3uMPo4R9yvX29cd3TjAwpT50f/IloZHPfrFvHLMGdYJkx
ImUJf5u3R8JjXyeL99/4pEVp1Q2sxoqdD6oboanGwzhSuGSU/S7Mw4g27wvJry4g
V+UE65aNPLj9wNPAH3u9M65gwIufJfQYZYQiKMO+eWJomSQ9OyUZdhAIkseWG8Fl
cIaDIBc6V6KGt3FRsehQIouzfhZbuzEX4q+cpsC5bCy/z6v6qTTYhwsIwTWMSh0j
blbtDYov5WwD6jHdbT6CRd9EaiJrA0T2ZiECKSYrLXyVf0VEm9gobeu66Od6Oncv
C0D5Fal321NRgHwbJIqD0BghvFuhWYPiXSeHYDuMZu1DajRAgSakcoRzxYGGQKNK
/7q/kibxEzr3qN4VJJ0zW/DbxVnGnaj95WES70iuS1UH2agFwjfgzXxolhGt1hjO
l7bzxBtc0Xodr9PW6/WFhOiPCYfFdCev0FxU/+kpdaxGh4JkzDs8m8f5D6z3Xoij
MekpXjmsNNTQqFnu6wApznPtcP6NAGCXvepOWrzoAD6AOxBkloYqTp8zdgaBfLaV
gOdjRTn5hRA6lVyOKsYST2jEUhANqzCYbtkxYecOMnTPH3KPO5aWbUWTKjqRCJa4
Psq+8g7+ct3GgJB+FB+DQ9OxDmV+z69lewYdFF/7uhotut1ZBnOi8ui/og+3pTzW
r6ECggw0rX0lYTcqjQ338ZvnlBY9tOCRBwz0xhmo4vWA5QuyrKGWPem+e73kH1dJ
8rLXWG7X6jgeWyDKoz3qvA41e7j5HqtUCEOyCndOlZUYn6UWDkvyOmrk8o0gzJgr
UpHojwhnytr2yyrmGBaBgWef0jXFiIig0v5PX7wm/H/eYW2pXYnfCgKu+jZ8kGDC
XhvYru1/NXWh6nD4AbrGbGPJugQpPr9W3g6XhSDFkTRcs4O8XDCMtKAHCpIdHI44
HFPMau9LQEZAmahGh8vcMTlw+ZELLpfoagUHtSycqF0XmhYS60J387YpZjMk41VN
pD6rB50pRRZRsuqaIJIqR0Dhea4ao+fHNIPVkRr5uIq/Yd1K/7KZWQ9jCsM2JOUJ
nWZ+301A7mEclrv9nOArZR1tkYHoK9hU0tXwgOaFuWdOSRupYxjHE/McYPWuOT5I
zRPp6hBgzIVDaj6DDkq3XajDuBS26Dj00OY4oqmYGIrEK9GDtmkq//zUjxeEfAyj
UKJaInSC9D0bDzxVP0RsnyE9d0FQi7afoHKa51LpJ/ahz/K/HmPA6faeCnDaueSm
4Bd+Wgg+gSz2/e7c0e/9fNZ6vZFmCQl7qR7mgC7PqChCjFdBISzCtbHYrEsrxzaG
5ofuAN5wBDIZvlzs2++DlgZcQJ56gAi+D0grRUNf10somDUysIjrAVWddLsi1Nyt
F8zDjtzVUYLjjHqDApROtBmT3rbMSzq7vEIuzQbzD6mMXovE/IKGS5D2iFi4r2lW
XLPOnwBesbAcvHFYYd2q6MQknXF8ovgjA0+R2jDhymprQDkTrsUaogm49JH1beZj
lIhn9B3yyBaydAhdFW7qqvU36GdM/rTfxhVc0UiGWWemDM5poxw7WyE3R3mb5D4j
GCE1G7+2G9DQ4s8ZhVXdVdeiseQQOIrE9pMJW4QhyNuIJrHbXAGL7ur7KFo/2MFg
jAclSQ6NA2B+2IuQ+sq4uYC7ahP2APAcubZg8uNJbznGDxejP9VNgC8UfBzLPZpn
V86VLbD1yxt4DYvKdVg6S9JEgCfdUz2ehrcAANJrX6YF4EnCo6AYVf4p7SpODT04
rgQLyEfkVcMyd8ykaFkH0nOdnyg4ImXP1AzWe6XEnFA8bisK1zLYYqgwPGJQ6Trv
cK7sthtkLFcqinKKSBGtYCuyArFumj/3ZSp0IlMzkBtoz0s3cxCDd69B1Fn3X89z
y5MG076HCTCjZnNaxzgEt7WR2cTvO1e2j7FmK7a7wYg0Vni47J3bGMvewFWH1wo+
3muFsZdowB0DLliGcJ3MN5wKQW5D8tJw2bm/QyzccIBlzE0pr5HNTbBohDrxbybV
Bf55Smdp+QuMWEJMmzxFO8BijMiN51OPlu9ogs7gncFtDLDh+DM6VNxBAou+gt5z
42Js7iTXN40nAZwK7L5H833kKg482V8hdZJQWTrTHH6WUEiGXaYqpR1SlA9TJ1Cq
j4z8cZdDxmlPnHOPDlLZPld0Sj52hNtDo/ZfpBf8FGcEb8wK4nNxLUUTsyNWIfVH
Ebddh0UPK7AgqyIhtozNFbPuHjXa7GZWkCWpDJqFC//iCjf4QSOzwcncMu2NPUI9
ZIszfgHuMHIiD5xxZSn88F0z5sViTWh06qro5HdzFWMDfmavHK07DIpj19REZBLV
OHXoN4EK5Ch2JX/fvdvz5PD3KlGEjDT/WOiygzFSzKQki+eBO+r1diMNLObnkM0g
juj92bV530BTuOYP03a6z7y2WYd/qdfqHOHb6qCrhSVktLErtp+ccSxvbsQvjlhv
W2G+nmitdRrrS5SCwo//gYvMWrt8Hk/UVdpagESzTmlC7Z9l4htAAbOhC/Zo/BaA
xLiyptMcO55hoj9+27zSFMOg8ItAT5HVsps0VeNqx/7A++fO6tF6S8/B+7CJ3MQq
6ZsFSzOi88jCGZ1mOLkg44Xoho6DTpgN8UfQTeLBEI/ssdG0lIFSiXuYruIcQ2Ar
Lmog+mYvHmf0qmqIENiPX2HeVMj3zXP8ENEee8maAVd8ijXncDMjhDEaPNBHePHQ
hn2xhyc9VSsLCldbkgud77Ktw5pXzIe7wp1yBYK5VgSPSdE3ztxH6CZEwvzG0Dnk
9I7sf3lHVW1V34f4PkWSBhwJ9CYV0sTmUtoPjNP9OvYG5j8+1aNidEeCqNa2ojtS
7SwshYOXVTB01fnF/PGGbg1dATZJfdQoEoORvq7D64bdWJrBbFHxovz7Y1sUvYnJ
6QMOd3dx8A+nPYPbNL1EmCpk5Di2XCC3ytStVkh+5UmGxuIDfIKCA0FYTKbFstMw
w34D7v3k9Csbdp1gek8bGJ1kI20mCgIe6ILZgO63rDbAhD9n2qtokt1kM7Obdndy
h3CZ6Jtx+ZrkX7QgxQLWZLYBuD3mDzC4vLwOeZh04EsAfDCmQvQ5raR4b3xXt+2M
aA/PdVjRF+c4C0kha4rMC5oYPaArp6nK8AJr56p883c3JPSP3AP4uy5W3cmVayru
YnbFZTjb3ypd3GU5LKpWPVw7rcJBbLB3ckfMY0YO+KeFsSomF8gvLthH9yeqhaKN
`protect END_PROTECTED
