`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48/dofoXGnH0nJj57Jof5mJsDbviWZWzBDJW37SyELUz
tFoPl+/yQQuv8M6+stVSkpZk3f3b08PYjgAdyOUZJ8CxmAxq0vKSqCw6Evyw4r1q
XSZTZQckmUfnP+0Q261gvMqkv7VAZWqm61YL2yhIwZxrfAmP+5q43Va5/T6mL89E
+i/C7ybP0eVQfPUMayX1pB2pAmkhrD+OJXjDsZ5V4mu/g3C/PiCGkt1S2IV7NgcH
V1UWUKN7OZlvnpm6IPATkmkA6DtGxHXTzpc2WO7qSyx6ZLIm5lB0kuMUsG6bsUpO
k2WCzSsyxqWB9/Yhy9NK9+NvQvE/XllPZLX3Vz/9lILsUB1twIi1/YFRvUWoKqZD
22X1jfxUZtofsktDEP3Sntjaqwk9GpuVFvH6G9cMH6Qy//grIo/bnsccuELNUn1K
ycpU7fyB2JgbIYdSMW5Ygg==
`protect END_PROTECTED
