`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aYJTFtt3gNkfmoUWbxz06q4tAldvg6UUxXukbKobhHA6
asPipUv+jzhmVeZpSkR/fre8KEd37XM0MZD35ur96ZdKEmcwahYCNk5K7Irapd16
jA7/+Lr9zZcOwF1QfS34qHTsBYPkGsqlM3ZoFccMRyzr2QpKeso+SsH/UBu2nOuS
Quh5bQO7VVGd8RpSu98IU3YqiJxEP2FgWaLK402JqH7XfkgLbKFwW2NdWci4Wo+E
PixO7KD4Ti76a0ji9RlwuSqitIktet8w08ZOzxML/QLhasa+ie0fdLNNH+mKa2kd
U7+Si7gYhdb5ink6Zr/ljUl/tkwcVENbIBjjL0QTFQQ6TmMiE3Mm5SZZzGa2Lbub
iXy//8ilGWezLQhEvLXzoD7yutKWSwz1OA0jLzQ3hlnpVW9RieEesmS/aqBdCrDF
idA5EXOlVLRuYcVupvG66+nahAsxwPtZUSB3ip/haAVopcDatT49/3A94rcGkkIu
mTsADRdb2uTEU9MuTW7irw1UQlCVcPJXgao7rHqSJi8+Ys3ZuRVcn1lyAoamGtcd
oAUHq2hG27W2RI5BtLyDw0tJtrQ0OiAp070HOQPbxbkZc3NjGhJFy/5IrK2eHSAP
B51QwdjJ+/doTlP7Oz0I4xLsthU916XAMbdGDbbNUYs2Tzh5RBlcnpymAJ7rLgZV
Ll2TkXg2/T82eE16aUZpq6fqsf0KFH5d1uSUF0tJhzde4Yixdz/bNyHrRoyck+xH
JhsN5kHDWtlwxlPgs9yE78OUzDOfZrlZY+hx7gxyoP/St1Q5P8sfvJvpiC1okSXO
dVVU+Sy9Z1fbgHY7GDsJRFySpJ0evIp2j9d0aN5K5qKy1rLHkNx0VmyipvyPCIgb
WO0euJAqexYxL5ceXhMx+s/h40HSXuk8tkf8bpEidSFS8zSRaJpO7+Lc+LbVdugW
hmIFOF/An68tC3Wdw8aoROOcpZdYfj7JDZpsg2UJJoCrJc5G0TJ+QCp4NguisbJI
3F6CXzg+ZfOztEJbO8hj0RKZwj9bseSYlAU8zgk9Ki3wVih/W45hoWHX4W51xGrB
Qb3LnL7JfXLUptSXMSwJ3aByGCWmQfJBFxHxBGZrAumNkuyZAUZOUj94em9hBIl2
fv5P4eRPfHqCLat7ege9g2WoTsMXSSPlOzI803EcxyPAhJsAF7wEHgjNgS9OsLmh
rlBXfp8uIFzWvr8o/Jl2gH7PY97Sdc2bJ2O4RVEFVWrpnO+Tgge2E3UIM1aTUxd0
pW4qJpA6BiXZpQ3nrCZGnjv5km6p9aDCva/NE7Xp30yIs9Zcpb8+MMe4CmyoIlj8
bchwydZZ1J/pHyc/ju8ELMOwTzmxo2mt7CILWaZJZ25CwDpNOZuTTw7uJ6EYyL7w
iQGXFfohDV5K1noTNer3cy64ao2x86OuJLlsbh9wMoGwA4t6uReSTknq30Pn4xX2
VjocExyMOzq4V8rsNWiL031OdfIq69mHwVoeGn5iHxzfknGeDvHLc39NHdur1hw9
qmeiGuWXh8SfpeWGT1bz7JfIrBYGZteLpTPhNMGpDzOmGW9yVcBQ7aR9lawOIhI7
IO801CzLnN64qAgvUJKVX5ETUjUXqrLYjux3OOxLC+jag66juK1eVwy5kD4zVDwG
d+FW//YhaAJiD+Ku8N+USxeTKPc1fYb0y7W+TSURH8zW0L0/03y1ftpqwJcAoyMi
HhmrSiEfUMctWcZqyVuipFP6VklBlrp7CTSQPsNgjLok2EIcNU9p7KvnBTfYxbQK
Fvamu/odh6bc+98s4cZxXScZM4gOl6CjvdmdCQ/cDeJ3WX/VrX3XgckFO/x+BUS+
P1JgoZWBUOx1Vi08dqH/QTT4qc+zb7CVIWltPw0VO2P37aPdp0lbT1XSYnhxHu4i
Hj9NnMSWurq5ciZS0MwIx+glAOWiSYm2JYg8/rqwldHD2gQRyeyOOR03UxsDLkCZ
d4boOyov0bsvK6QEZUE0003J7WRDqwNuvyPWYVl0ONY2FnqH/v4g8s2MS6D1kwuX
jB1OPPtTSMIU5GVj/+u71yi0ke6RO5o3XuKsGRnjhZCiC5VH4SmtLi2bR8UiZWTo
0bV+Ru389BDxxjaFaF/EdugXoZLVfm1auAx+VIVHx8RA59REEzjX0pHKswCe1V59
wlWxlX9HMlNFgCfuvW49woOrMMKwba7gOqk+w4XdRrIpyOabXN9F2okMMNaJPKYe
jrfYf1zCm6NtPyWttOBv3THYJLg1kJzP+4b3XgXbJ0N7vs54cFTT5VEt5E0j2QuK
zypjBtHACLCQRowdS9zesNBmmu6NqLvuTMsBNLsa1RI96EdrDovmihlRqvBh5vxy
jCya+hNvpyZwGkxPeCdv9lGSAtmDdU671bmej0r9HZ1B0r909aeL+ejJICqLkqjA
CyUtrDpddAYKj8gw2867A6ZwaGMl/3rVZgOuy0oRifjM4CY+d2rtHV/O9iIBUgnn
dprOO4JCqJyWumWharfnMQomW66oZtgG/8an1CCTnkotkNvkZ28QRrl1GKiH1CUc
hj6Qy0tszxWZBIi9ArvlfuAhGgYf14eBjUk63xccT9fsaTvl5/7KnKY2trdiVEgN
juXcXDFIYcKm0Arv7ZNA2WHyp/eIC7F4VB/AwKrX4LPa44GAEH/sx6vp7O5yGwR8
xqEpbN0Y5xMkq1tWQvAotbNBHGdd6+pw2FPxdCG7JOpCTubCvAi8F8h1K77DMHso
`protect END_PROTECTED
