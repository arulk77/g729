`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL9RndQsa5znTxp3gPS67fdds69mg7678KCxiC00gEcI
+YJpQMm48pbm6MPC9sAvXbC8ficOXtdZd5Kp/d/3NlZR8fu5JKDxYH6w8vTtUFKo
ZS4O5FD16SZLNHUupzrr7DZC7dZlCPL1CxrvRS0nXRmuzaxjOZUSFIOxsGHdkRKl
78fZPtGhz0Zo+ugm4UZ5b25XZJleWYd4t5fdtIG6DaraGYlpQQvnhmLBcMwFKNvS
`protect END_PROTECTED
