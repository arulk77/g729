`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48AdjkRjeEQ+ZQ1gA56GfWgt50K2to81Au31H2YRfZyP
CXeHVixFEQqfylq6Fcsodg2ThYr3yIqu9EP6Y5Ggh/QBg6KR6u91bjeZ2btwOPEK
VP97exxcupIYioX3/fVF9HIllC+YlxMLLL8lMF4AGfp0K5EjphCSAbtv/Qcevs5D
vtQ2GnZBHHFaUah5r3wsW71UgQJgNvMxR1oPZWMrdmo34zO79/LETfGKk2VPuh7C
JPoGBIq7Z5L2wBKj/mw1FK2epIlzLbZsJkOoICkfsjA=
`protect END_PROTECTED
