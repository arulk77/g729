`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKerXs0sSFERooxSkvW8lnZTzZDtOzmxLsC4BbWl1OHr
TS9xfcgi36PCUqqJEwo9TDW8iShoeIIANNI/WzzlhrBHBl2WF4HQhiU/NQbDSRuu
Ft8X1/8eTs8cJX1v3wGnZfunHLgIlomiHFyZLowd9T5V1WvArrGjZFZKsQbOtuUR
J7LnMYT5xlcwcS/HoUDIsut0uoRHMrnvkDnzkg+S/b34bMXv8/G7pH3PLP+Vk6pD
T7We0Abv0P2z+zx9V7qqT/jx6Vk0YDIuV5jaXlAyiRDIkZXfG4pVvlGOpG4IxBw5
3rx9qrETbQb5V8R88E4NWQIfUIeKdVKetskPnXXWRh50pc2dWKp4rcv84EL7egXN
L2tUFFyClVVAlk3mt7/NvN4CBYy3my4lxCrwCzFYXQCdUCAeiWk8/v/Glgf3j6QL
DPHwuIZOoTJvVEZFbRr/pPILu0z/zJjYqtOpem+l/1dpAHlkYZCSEq0laDRF4Qxj
UvRnAyYVV5JJZ3Mu24dj0M1wloUeiyOHeHCTtYA9LyP6y5+D8TQDz3aSJFDrsc7K
2+xQeS9ZIYUEFxwB2ak8IBDHZX1ULcWiHAZUcwH31vMX79TTjj1lJVSo8AIh/HAu
3cPehfVipo5JP6w6QzIxuSs1Xe1NJkuaOguN22DB4NWbYK1iEWol7WRKXH5zPkCL
/kTQUD06wXQMebzAEZ0cDtK8B6U1uQdu2BcOMvwI3PMLjSQPCTk9Yc1YW0Gt5ClF
OLXzX7f19fcZ+NwAA8WxNrJqAVIBKXtz5xez6dregYKcE2BGCK9DbuZRRHeUQ50j
sDrCZDy+c/7vkEWPI5h0WlmnjGGTf+FbSWQOdQJce8NRWj6t9Gjsi2v3mTlzkdij
mIp9lV9OBJcQA3y+iNVKdCPhwUvidk1n3NgcNcD7CqKGTsQ+E/t/5N69bzyJhaHx
0ESWcVRtxfxscf6Qt+9qwtETiujRHyPE+oL0QJlAAfr2DyxUmVECXvW8BEhcSQ3s
usC9V78GETQIEVRPRgFMuibkKBWpE908lrK0o2YTeTjUqbq7qGizFhUqf61yb7mR
mMZnsyq3Ol7DomM1YyMIkF8lq0gQVJ3GrFE17F0HlL6ECLP5TRX4EwDGQC3iuiGm
YPkSUoAL+MX1180uP9tWZjc17JE3LLNOJzocZFtS06CMaNhYLlpVIRDXbnZvO30A
1HT7A0Ty3hVcfFCk3IDyIcUMNUBk7lheNRVpA43tB7koc5w50ezTxgDEUy7TW+eB
S44QEOXzwBopfu2c2ViYDmf/3FpB7Q7x5QAgePINkWrx40BBKK/HcB+iEzIqNylX
GR39jqb9ITzCNtdh4kcJ9JW1vWbcL/nNo5OKZyI4+s6ztYpYo6DBDYzpF0PokdP5
`protect END_PROTECTED
