`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJRM9LvXhzpAj5Xxoov5mbCfTra4jL4ZevXr8na5Luu+
L/d2nsqJ6CG4nTdoIybwDpzHQ0t5+ySK9Lb/AtDuMuhbiAG7V/S3956CsoUpsgZt
tkAy1Wuc2FRL2PIZnHa6MylX/9oIHx0J8Z5QQZLY27yTtQRVUjC9jgeU/0nEQc3/
weQ4qOCIVsACHKBpdYXXZfek/4fuoXXH2TFPoKsppx7u9dp4u/IvYVm3BPzjxch2
s4SbwIHWJdf5zaQ3V811VzdCQo1QeDs1oT+h6mHrhDxVyBYPVvcuAxZeX4Tpc/+A
Hh3l4wMDgBhZm0HWvGEin8GEEvQtZiX5yA2+YwB0rxmSdrKj3quFARJGj2ZwqfBF
UT39QemYL1V/ui3hTm4zK9KVtR/wt4R4D7aqYR6hQgghtI1MGAxMNkqaehOEeIfB
X89I989kt3rIY8ZJ7afwPNOcP2EZmA2eWbitTj7GgIvWl/w9aREn1tYHz7vP5hr6
K4WXi1w9HqTbRoOrCo2j6Scxl5i0P+IT/P83OCFx/mWCJ5lZpG0gCEjMYzkqACcJ
0+74hncCF6Y7uSH8UiJg4A==
`protect END_PROTECTED
