`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMTbj3yCSw9nOmX1AiIsogwAMymNmlyhxVfeTDq7FV9+
pre4vdebyG1Ax+Hx99r4OlNGAmsNT0ATvANS+cb2uUP7WTuB724mnS2Sx9XKAAdN
/141cEp3EcGsEtIYhEb2FgvTOFZvsfVqmKktH5Wg04cRvTI+iEIuZMXDtTYXLZz7
m7Mc2D3NUNfI0aw43GHfuKN5l5aerONIcEAMtr0u9anxssPVg4GCovrIX++vri2K
lch6C6d6FiTfKgBrpllSA7GR2IP4favAFZ0GL10GDjfq2YGNHe3xo4d2/nlEEOwA
Mqg2P/xH72hi/rqssGFKifs+C8pEjxP7MDEqjVtUKn55Xm2M8fmkCOlZOsT1NP+I
kH/V/I+j+ZfthwLvbqM6TYOuaetvbVq/GqSjwTP960T1ZTbUO1OnirYeqoeNp8Xw
pRhyefloBz2ihUwJJUYZ6dCRMpBAceJ5iW+SO20OeGvDvsF2q+tNqe8SNFlsC8Hx
gKtiymkI9V9Ef8YrPP/rphazZVu4InUNKdJsDCONH41G5bk5vLtK+HnPkmpw8TqG
`protect END_PROTECTED
