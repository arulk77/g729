`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD89BI25at2yy5IJNTKKHh8J4UJT0FZBusA41tCJbRaq
jDKCPyzg1FbOjNq6PIE+HS/O+LFau3QvflKbuVqhIrlndO3+KepRNoCtZ7RY7T3j
dM7Djjdf6asC/uaP8tWDJ4RW+cG9/l9kQe7QpjpSMA3otTy4oHriatW0UpLZpGmW
Ziku2wqVbQ9JcuEILeuYIO1btLDSEq/XL8tfIRs5PeNOPsaEHQG5L3Jcf42amfs6
YBYZ2J3Onh2zBV23lTV+37E2P4Ugnnqu9TQCxKc/j7uyD+u3dQasV6eCeBoK/WyJ
g7FnVWVCs5tk03uqSdR7B4XbjPhA2QWoycyFH1ikBsSbTfU+xw4XVRxuElUMueUK
3BD6HES/PXLa1drMNvd1YoqUPVJ0d2vTfeeWoMYRONszJpydXpi14reDOGoDzRIE
ff2VaG1h31MWmYJfRWIDlxB9od7RN2x3PXdqg7BSHzOrQSmaxbINbZoVJozQwpeV
Yd6O34NzdwUSF7lfKmPdwhew+q32bLk71j8NsN8lsMMC3qaofDfBpCcV1fJxpaJO
9EbZTQPA+3Sjy2c6cKFrrJuEkV90NSgqdrbR57LX9Jc7l0GBk/GPFzTyfeieCdKO
lOW5/LTk9OAwzX5S4UxcDks4m4MKyMoEAzB0mtoh2NB81vEH8QaqRzo8ttRawe9l
`protect END_PROTECTED
