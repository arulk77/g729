`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL82qsigvvlH+rKqBlT7ksoM2dujnWGiRTgQTucACN8Q0H
HmxWLHxudjb7/gBIZzhwTI9nCj+AesnDUl7RKjHsIEcB9EFvt3pZumYnaZrnNRVs
qrgRNu5hBO4Onx/tGW1PLueDc2OUkSfAIxBnyQt1K+46tEkRQ/B+QUNJCT5WlqK1
Jk2di52QOTUD/hj+n8Cwy05XdtnOZQ5ItdbquRlOyUQs61J60/W7MxkjDCKNsrxL
26vWxYfSO2zFJ4qN4nhPy1JeZMWLPz279mYmTE96ODCQJAeUUJh7shO0xAFfownW
phtAG1LLB32JZhWHjm8R6hjahJHxt4B8eDJyrJuG889SnglJ7e+zv4aOYeFOwcQK
4cIWskXHDyRSZtedtXRhMVJTiYWZlPXWKDoUJiHUmJZKBOV++jxUNDNJG3NztErp
NG6A0/4X46aqEotj75KSFZ8KzM6rzY/eCm/nTq7Cz/wWVGnC756Tvm+kcwH8npM0
vDbC0A+QVrlHgqQ+Xc067VmLE+d9tXwvDyKp6t16eAV891Up/3H6WpZsVn5suRVm
ikfy4+m/3o2zqy5vq6pDSabmeU9u5xwUFcV/HASVNpuowVzsrFlIFdlJkaGnneid
hobUEsFfubRcGZEHQ2Gxbc+WupRCaBGLwQnFGPsLtiQvwpon2QaAQ2krvynjRcKG
IAOEvTr+PSxsfVX37tmkDT41plA21KL+6f67yK75D3WBxmc2d/Ooi7zWCiFGIJIL
I7Exjj6hh5shR7d8jC0MYz8bbIqvRRsBiA25NCNZQmICj3xey9xmisWR79bt142S
BRiCy2LUCncHO5xBo6ABhsLiBdv16cJ3EOkf2CMnupZKETro2fdyQwX1/x+t1wZn
2JND5HyNh5+/P4ax9kQNYUWyv+rEQVAdG7/naC6tjMfNDGFw8Hf9gJ6PHFB8q8qp
8tDXIRLTXBF6yLquS5F+lVgK/s5SclCQ7yIooM/ng//TgMzcR16XS3emkoeFR6ra
v2YJjxe7RvFxOX/0+69JNlBayiCaHcb8bhTTIOJVs5vIxjYdu/j15dyazp14hhEY
ZbB2bZ/Hws9V6Vc7Wqsy9ST2NNnz3mM7iInFNzaLHXIqNdjNT3bOY7iw1AGzthdc
lk7hMnff7clBLcEpO46NcNtRxrVqGQo0RekHPX8+MaZAJrlffMN8+qH6IXDBEsuw
1IVuZorBGQF9El0QW//xyBdFiIki3xKhAWo9d9nsoOxEM114Ri0veDRK12i8twrv
OafhCbKmNq2o2nKtH1IWdkwTRznQou1mgpicRiWcsx+RO+wt7Q8PwMxf+UIwTtwj
XPGoTaPBwP7dYUN1WmOnsYS6exSxkJR7V+UmEe+AtPwNSpYxV7bQxHBgtSYjBdkc
e4BW57e18W0Y3TsHOzJN/XGFCQ1NYwKgP2Z0NzlQbATFYqpDBRmnR3e7K8LKSnGc
L3QE0DJgluFG6L+Rnh3K1Cy4iREoZTas5wDU2guua/xUARLFHPTTzQ+QaPEPScKk
6Xyd6jTPJYpdaLFXD17I1PDZgYvr0D7f6bGOq934+5Cmw36RvVkYNHiAzz5QNB0s
AbmDonL/ZiPqK+Lj3rEcJFGV3NVQ/NGMcqxYYQj7HDMD1yNKDPfzCMn9uzQsmEVb
hiSmuTVNvxYRRt4ZKWYyXYIYvhUSASNKrNpLkcjAPmuEkzTTomXkbnKuWaCrM1KQ
NFrmURChJ8KwMCCkYV0+MxqAP3aocunnV4ft3pmFlQcAlGtyPY2ltL81vzHLrCFd
SfuERuSYCAkNZ1s9e97OGj+7wvgjvVYb8z+1skmyAd9ZAYgB9iF6Hy42V/brPDIY
l0rbmv8ko6y2ST7ZCyDl5asBl7Ko8nWMZnkyNG2skM/TxyJGpG5HPoABPo5dEd8J
Cf8mVYUzTVwzVV7rOzYg+YqSFl9v2I20/9rb2atTGEaK8Gr/HRjy67rfmUHA3x/U
`protect END_PROTECTED
