`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNO2ChH3GxbAKElWdFBeZ9FT4DPqqPi2r44zRNV2ggIi
U3nm+FzuiOPGT0Yz294EyszA8oQny0p9JYUpRJ2VETQopGYaClb5maRzTIi4gTqg
GW9Jfdr4boxwGBZ9+96lSlEfDC1L4JASRER90COv/b+Dy6WHOKNtpBCBOwjVJAS4
/QT6Av7ACzTNjgaFZHFECBmpGpi6fA5NL2k2JLlVUqXY1xc4qLY88xiOzpRkWjPX
`protect END_PROTECTED
