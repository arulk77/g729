`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yrZ6qxFehaiChxIAmMu3G6+vFVvasbFHn5g7CfZADlA
Ssgr7N9ygtWfdvPOUTmf3tNG7yBHyrS+Vt/17ZG78RWMN4Oh+Lht33L6mVZjdzyO
mMgulSwo6Y1gEq3RYrqUfl1SQOaStL5krPRqaW7dbcSgZ/c9It/8FaS+HmPTVube
Xk6GSHBvR6CwHF/Y7QPsIZOGRjEAxzkLSbuhRC5ac6g=
`protect END_PROTECTED
