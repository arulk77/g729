`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOmOUH7w+X5uMJSm68RMPAm3l8zJ3Oqt+0y+3xfSHVl5
ylsUETVmgMOMjddUrdY+FLOirCf33mp6nNS0rNNAzWp0Emw5ZkSs/gMgCf/E/IYj
XY1p8OYB0ArNajhPq0NMpOu2dA/QsBIv36/Wl++49/p1Vt8gHslvKXGq/m5T8pSY
zK1iA77mr8QLRgGy6eF+Jw==
`protect END_PROTECTED
