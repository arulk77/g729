`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
hHmtdHCJzKZombVd6eH2IHYNzlIBNvY7lAdvYmHOJ4zuTXAiD4RMzPL7rW0zQMQM
IK2toPwnTrw/JOWLpEe/CmJCz8O2/XQo558HrpaWPrdVeH+nvyydvirwVZsxvZ1M
irAUff5pE3BNQKRw6NeyByMuFu/AaeBwhzcc/GfzPJDDOHD79ikBmPYbz/+y9euG
q1DY3RQ5lpJ6fDHiRGlmE2W6r9psFkLx19utUQXUF90gXVyZCXtaOoUlkp+nzPs1
9f4sgyQrh57GA8N3Lyco4yqANRd90R2N/ZtxW5l9iNY=
`protect END_PROTECTED
