`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SW3vL+KD/HaS+7kLGP75TCYTK2pfOu8H2OJ0kYq5mi3d
tVb9PnepQ+Gpx6S3s0eOV0yRG5c9yom5LXN2INxRO7J9I2Ilp/IWxe48j+e6/PKN
9bG7+nbj1NokFxYBcvBe1L2IWHgf8VD/juluLz55xSBtzPUSvrphF1UgFcz39syT
gg8XcHrmNfQ8VOXVaAjsMJ2KmRgNmX8gVZDbg6dxJAF3uSOMuVh3m06LWSC31skT
s5VYAbad5nwo4CdUd2zG9ONgeVDwQw7ENZ4d+44JM83Hp5PGLo8hFfyXbu7THoUf
qLm9dhAGp/AuBFtZ1IZWloim6CnPQj9bo42flT4TMkYcWfJb4h2pOqxTV442ze3I
bT9CPg8c81JFJkIfgTjbTvcd49hhcB5UrVNZPYA3j7Is+jz4/xDwalRKTfH18x1U
n7xO8XB4ib/qH4qwaDV4otF0YttPtakh1V2np1A4JIL8P5h6YrL1sFeCwMUYu/f/
HjzkhWzpGnXzgzfbFmkVDx7FjgBgrmj2N09/LDhJhHhwr1EGMDd9/BchQWtZVQhA
01A+x50bYsApfMpVblInAu7qIo6jXwZtsbDsS9AF7zN4xQO+RLz44aLhKRpoC8lu
rpqVGOTgLpdI7S0k/ipTWm1odHkhQXe77l4JGMb9CrWh92d6KDrFqcSJSfTF7HXU
0o9PyZBYh3xY3KTItVZDiZIbHF4PxsEjO4rLjTOnoYvJA9G0vnGW4PittFHxMmNR
7d1h0ImTBVHaMO4KDBymPDJaYKqhBFcGhs7CmxMWyouuz19jKQ+c//EM9AGxIeth
Ruqrikr7ZdDcq6GoVMnn8QHAZwTFUtWpdaGX0CAhSqNpRktIAsSuiEASGjwMw4Nx
/OWt73kkQ3XFjzK3BZMdc9V6uE2f8OY0I9HRbiRIHZHA2fYxarpDxlCN8ef8KY+9
aaiaO36bwYop1pea3bDr3kwsx73QgIM0uCVmnEU4O7rh+zPEDIl0HcaOzMz2C3ck
bvqvupPGZQ6TGGavJzmU6mzOpty1jQy/JmltCC9L99wMpRpg5Ba4uiFxtuXgcLUd
DINfdnJ83FUbKFAy4snVGhXPOV0SDcOPUlxIMl/6ureM0Lcx94WbHEmZ1GnJJnij
eq9LkHY5hlOd7o1c664L8NX5xhOiZSaAIRWzJ3CGPjFjBHQfMc+dTxlqCy9cdAO5
EFXTcmi/hsU3sEv7Xt+PLN3hIcCJlZr6snNptGldh40WR3PDC08qFXJZ0jeMTM+i
v9aqTU6rWXz6YD8UjH0jEJx0zT1moj2MLaztrytrw0EYTduIqUJkrRX6Ps79VPKR
5OScR8uD8w3BUH8cJ9qNQoGCJjWiNKsWzsUV53P8lKRs9upZCJli4kD98HlxTruj
8I0DFibk2v/G68tTR1auO2m5mJEZ3YK/Ngbd+I48iTYt8KPyan2ZlhU2w4aA2lk8
hPTlklujdKZ0HRAiM2gML9gzBjl7ObwrYDODVI/8cxyC1fTVfPVv02qap7VuTfsl
feFb4hd0q4R/rqS+J6YJolGMBPxTO8l10ULqW+4lJgR3Mpnp7BmPQunA1gWVlENw
mjM1Cz8n7lCuSxCXgNJKNSwkPwSbX2wffIpy6B2qY4k=
`protect END_PROTECTED
