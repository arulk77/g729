`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ1BB8cQ8qJZonCkShZlKu4Kym73CGgHixKGkWukFvH3
ziwSSM619T+IIYYnfRecxUHZnHKK84VnKfxFWupZZFWDU4vJTziuxInxfOFg5srK
u5CQYy7ydriJBUffJWhuIFHL3eJi/l9+FHsRiUHuAES6mLOvcSv0RA9djf7b3Mw/
clsAaiRX5lP0BuuM17e7Wpg2vElGE3vSPwgGqtCYBrBjec7o7we/3x8ZdgJRHfUf
pArI1qNwutZaXVwYUoTAeHjv3B6+/gp3OgAMuIEQXT9XXBtb3XS7a1RtaZg+FMKO
lDdQhq/2J5xrgmW4cFGRVe5860eevGUL0Wwj0Q/SlQBjSem6BEioiJS3BNJRmxX2
ADzlb1YVL97H6SxOjKzdBuSgfajbdlzQTWO3KqmsUpJLvk8aRkzADcM6XKH3Neok
/RhsRtqmWUAew/+KiBrWF/KydM+DRN3TGScTyBkfLR17MUg3zMXeIWONgQBAJwyg
1f8HA1PkjZbhsHf5IkB4KgIeSVhDm55egdWMLxd+qGBr0KFNf4SYweaeGh6uCSkm
6hkJ+X7rkFB3L9RXR19c1vcaGXFUX8AO4RbUBDgepqlEvwKoKn65aTBVEoGNnbZS
Vonf89GDoXQCeCY3R+lQCx3EookhCxx2bBglEDOzgS8AEvQpe5J3CeuffSNG08+q
MiTLOpCy7tMJLKDVETwKN31z64E59/EqKm51OS6Iyy7IimInCpIk7/THmGc56iv3
cr7eGSF2WwTnb8Zi0aDcVMQPLpA3pGoYT6O9UUL0pVHPuDduEzx24C6SBop30y+z
`protect END_PROTECTED
