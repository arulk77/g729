`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zM5W9+TQndD7Src3uxP72ExriQyvuBLFcdIcy1xftmz
h41nsDtAkuKf6Nbeq8fslPGXWntiMiUA6NMwc2q62mromZxBPLAL/96jFnJa7Ehd
aoELp0l2Qwa7IF5BKuwh7JhYLIo/EbXu4rwJoZPmCw/Ns/dFUG9G8gaADeT64W9Q
r8PyvJQQGxhYvdtnk/r4GkM327hVLvYQPdemYStZgEeayMRUwqVwjvYCGx3RzKai
HyV4J0QWifbEXj2gigXcm/33x+KELCgKDvFf41c5q9eL03MB+0vsG8FeE5BzA7Wq
fPnwJuEXnGw0B8gSEARfWg==
`protect END_PROTECTED
