`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveELCqyebf0dxcgpf7k+szjRGp1mYW5cvjZKd5GFFHK35
lNyjDdwg7ISLzGTGeNuS4C00G4H/YhpMl9HeKF1y1hUJwXLjNTztHUwoaKhokq8A
7ZEAIA/HxD4sot68j4zroPLyGhBtGVKd2+AruJ7vRQun15vSz+F36BUl03X2WV/T
jHOv5fUYlLPHxVMs/sW3GPhYDjrajKx2HQMI9Ywkbapz0lIF4fxfdrEoyjqG98rn
IWVoSxwkxtaNrSHcUmaQNw9Y2RDEULPOrCVto/c1IW66fLMmqzBit1g80wl/o/Cq
p+N/yl6oqAO1RyJCrOzPEq2R835J21sRQEYHpWU9FPAo8YwMVTH9gQkGYS7U+y1/
`protect END_PROTECTED
