`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkRUCijt1erXuU1aKr1RnYicH7nasiVo7wQ1+/0PpGFEU
R2jFPbu0KLh4z/4F3FLfawuPo9PBEdM+9orUpHgr+PLmBy24OW2OFXEtKacNlLMy
la4HETy1HO/Wip8EdOn6ojzbVltqHcUXKLjQxrmPQw6LSgUtbcVEv8fvvIR8Gz0x
MXepiYOSQgLkxMcNHNi9wGfBaxsw1JDdKf/nwYd1PUFTaHlx1vkkNvgjFOu6MoQ8
DUq0Vpa5fXacrvJPdIc2rLvQOfMFvaj4au58Vsd7L9XOjMZNRjLlBgZyXQYICwFI
PrFUiR5OPcVC3uTiEOhxyJp2kuMD2abQFb4M8D18+fAgQ4/OpGrSWLXQWX3qeNo6
f1+peOuRg1EadG88eykzhdl3q8DkJWUKM0Bo+AiKGCA6tJuqQ4I9OQFiNqcj7ZFz
bnZ9YX6n5dGQ/NdbNSJz/6zKMjUb6+GwAaHdl1vajYdCOIopo3zoMo1gDRz5ARnb
6KHs1MxItoXietmChP4Qzp3XbO0IlGT9O6IdRy8NhCiFtFxKRQAzj1hx9LZhicoP
g5pnk1FASyrD0metRnQ3Fkwx4bKAMnhcJ6/ztG2UGCdjZoMPvHp4p6BMLtoSMQsO
Co/fMCPfnm9vVmGLp313C/71dEo4SMX+FyzaH6P+oRZNtBl16H+nud7A88TUyC4p
J23EMbPUwqgE/U0k6PLvufGG1KLeE+Abbrk7CJ1XfOdtj2qn51JuBa056YwH45zl
oUOQZcyVGV85lNzV1XaZV5OuffSGhvAZ/l0ol0inXuk9irCgHufnoRbbCTXIDEii
vT+r1HgI3tjCrtuSrVVpYSt7HxiuKGu8itxMz1WFCLAeUliOHr7JfqRVLnd8rtIt
TBl4U3sFniH84L5HJzCnMLATUsh4Nitv7hGWyx4ZakR26dNfvOuYONuV89Q/ZADc
bSH0GcO3As9YYA4+capc3yxREAtnWbZxPMUIhY5GJtOv/dloHEF9SM1UCs1ikoiZ
T4Lxm7rpWoV5vTWe8UpaQQhLy0ICNcAQ3acrinGt17+0KvXAVB4Qje2B4N9dnGdu
Jg9RsTQ7oW0lx6IxWn8jTG8djl1p7CoAT4eqfuSiUalSYBXmuhiyez/mADXLIwcC
sYXuw9WL2A4d6n3x5eBAbdX2M51M7LhhkbGqSVv1dYxGePWBn7BL2khl7GTMgwle
nRM7bP/qyhAobpVR1VO2/IGLWo2FcgCSJBizK18kTsKKs+vkhbGH3LTAS/kb1AVS
U33ClALpbecvF2EhY/IugZkU1Da0MZtLPGQzx6HLYEn6aOppinRlaILCcOlaRyi5
D1saLicIJjTBxdnJz8ckx5wheKMM0o74FFdeollz6VOli859r7Va9hxIpgku+O41
Rn+do5xaRI3dPFZvHy0NU+R4HL0BT7xcA7kiHtyJDcKH6Y5o+6W1ElCuNkwNfWZi
Z8KKjlmQQ+x59X/wxyAq8c4P+hG3OdZuYSeQLkxkVp1cBTjjigUVxnDrDQWcYTQe
7e7Qhyg+3nAvltz4QDS89xTq5MNY28RJtOuUdVHEqbH0pINaeq9seRuVUI6Ntcb9
`protect END_PROTECTED
