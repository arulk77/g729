`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveO8uRoeTsfIFsV28jjh19y3nq6vZXwPllHENh9L5RdZE
p4NbcvcCa+rRW1mIqmsrdJVkLn9jFTBIbu94dHIkvbycttSApi4VQ+Mqs7xyzI1Z
UQtFx8nxgNz6IkXa6mn07h41hKHjgnWN8tAE+BXvBB+F6ifgaGlqxfu4Hs9nXAFZ
9llM8Rlcly9iigIRp8xHKR4w+IcFKOC9eeDZlhhQopTTm+DEY6zjcTozFGBnNjeu
cIBjqzZLI/2DojZOkllTO/5eNoMh1X8pnBAQ8R9BuYgvepJVny55QbuI/QTqSz9f
IsMqO+WULwksDPyt9cneUEzj5K90ORyPcNvoZSFqVmOXEwa5mtbYrNcubB2JcRpI
Q5LdaQhUfre5b4BTVVRBpjeqrUWE4Vz3qR61R0p66BgukzpyNsbggHChtaswsCYQ
kE2yBIakRkWKrCm6T7EyVOOvbKwNXCgoMxfRzqFOPyAznO+ZiPGMm4u4UHKglzWG
VIz20OE06eI7k/ExizEMQCeG6wI/hE0yBiEcKJdmElwvaXFeHNP4NtY8A4Q8j7pI
b8eEE4uEDBIJea6oXkEWxQ==
`protect END_PROTECTED
