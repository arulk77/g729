`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDZAAmBrKO5sxb1Tsg+9fZC/Sm6KGA/Juc2GWEZMzl92
m6zk8AQ5ReqfLkBoIGYMcf4j+qhITE9sGDRaGgwM0mKJifOi6PA0MULJ+Oz0KQl6
s3blK+kw4ZW1HNmH6XCKhM9F8vNd/CDFSohZAcq+EhW1CSZDTA7mVJzmoZDj+cv3
/T/qorZjdS/xrS6e7lMoZE1oqHAjTN0tE4QosDZlBdTwUiPW2Y/P64U3QFY9Eid9
JvQK4uL8T3tzPnljjBFQA33o3t6Ir7PLFVdCNXJo4VnuJdP0AJV5WDBBmDJTIgP3
8FIVOxwWxtJ3qa8zGPdEVW7rxji2TQcL9F2NUzFuS4wpl/4rCHXRpOLqJb46gIcB
ALFl5Kh77FPit0eOIXehGOSr4eakX11xvHnZ93eT6uwWDo3GiYAoKp632QF5VVhp
EEr7JtjG6J0JA6QSb4Nr2Zw/OiC5ra3dq9VkpcKYa3T6PnE6bZTB2MV5dlraFvza
l25thI9keuc78/bihzUVansf9Hk+PYDhPs6BOcegWFw3tQETWk76c5nfbKfmOF2r
sHOZWCdKvLjk94j4UpQ0re6UyjW5sCYUFK0FCdMiMH8kdRzvPEp5hdi2jQ7ivmA7
CQHAO2r3VYReWLNa+CrywZ2rzTuCHdeMD3OoD23SuVXeJKlT22A1pRS5MklBC24m
`protect END_PROTECTED
