`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
kyUKPC20xrxU7IL/BnPLlbZcVWgDMN/6fb6G8UyOLIeF6scSGpgsl1artN+00wq6
3sJV/RCgDNMQ2AzSA9L//q7sEsBiI6TgChlg1G4sMREoHvuC2fPRFoOA5KRwGzEU
kt11lM9MXJ6FSUjZFGf32F44VFGxcI7WJ2AKkKD+YFnmjgrcgFujT2b9Ou6a3RET
PJXWxp6Mcuzu1k/p2mqjqu19Q0vPki9G66TYLJpBFYgVWoCl7MftLFtMzBgjcJzD
Ol1grb/ffyb1UQP0C0Eep3gt1QOQ7Dk7rlhUsGy6BmYqua11fnozKlv5X4SVXdcL
g8i9+d903WSfRsPP0xZP0diypwoyp1maOJ+1C4DjA+SDZCd8orJyRGSPc66BnuDF
5gdQn6aqVLpitL0neJ3ukfNe1j4JxifJK2HeBYp7BpE=
`protect END_PROTECTED
