`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK8c/rhYW01LzLULXLABUROAEB477i6CFCF32NHYdo1d
Awy1vkdkza5GvTheU4fAL6tYg3QJJyNZiXB3ckM4XzK/6Jj02he+NZG18oTPCW3d
f/QLZkKg/bzB9N8WseuX0oe2ZguJ1Yg8BsKpqmniDeq/hnlE2UufaBrMliZRUQ9X
vd8N+VAyQSSjIAxfSfMsBDx6I5+PO8Gg3q2fzjX8qxJsBIHPuwkYe39rBXQzqizR
1uIDSKm5okxkuQdJ34MNESSiTLRgGwi51riO8lyKhMg+eqKuBMJip84Oq5dKo0VM
jq/Ud1skl7WaXEbN0zGfRAFixtMKT890sh2Kj4hUrvxY86Ib9NsKSnouxrvHNFmY
OWVe8GbtCRsnTqEWrxnBWUgIezd392x+0JcbAD5P+jooYcf17VvZhNgqS/HNzeyn
SgXAWhD7zcFNsFhB8HzIGFbpDjNfWSD7lp7Y4V49VcNDT3Vk7o4ziQDJcIOkytaZ
/GpQBvwnTfof9RvFxN7VvrkEcWqiikw2S3poIOtsvGfIm4jj4T9CVpqvyJ51JT/I
K/xtVlcCaP8vGKI1tZZhkYrX/eiqmHDpflILdBxGMQk0t3WGPwwd6LcWQWltYPfC
zbXbgoZF6B9+YcuEdAPhZQ==
`protect END_PROTECTED
