`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1adUT9qWdD0lF25zH/aAWDrp1oYYKNQFNXb9oEYWWLhil
g4Lx1S76mrLwrRwhmbd1SPF79XMq9OyLzuIBlmBbVsObLdknA4bGOKhiruuNJeY7
HzIvFxvmZ0ONqc5dJ5rfWc1oPHaQpKgMLjjIWymL8fO9cwGOrtIur9Z0g2xBZMBw
+G0q7fC5OghwdssUgfb52Djn7+t8ZhhVsRVeLgsakAau+1Rz8d1aXYwUFhqZqNKT
BGVnZhGoQy9X2IhAAY5xTZDxjpzMM6Utb02NxQOrEbY/yz7qBSc5QqnWm0QStPYV
ShtuzBY+TmEqu+5iwhH6L41cmn0IEYw59gGmlIhVhJKeV0WjYj15DN0Ow9Aa5j4P
FeslrjSrYfmCp9hkW+1UEZGaJIUqWbuvGY/rS3Zz8TbWYTKgOQViHI1m2/7R5bsI
xc2VLbJ5urwBhgsRJspMLZyPQdmRgG+rVPic1531nrz9Kq+yzTafYk3tEQaW+Zsr
fXOg6HrCoGQuanv6sgLdmLHJokKMLE3pT0y7VUEFvtbRi1TDg41A4ObEGvoLnbIg
7qaxLV+SiS615BZyTm+UmJPGsx5xFVCyRj1gp/9CgNFCCpYAFEBE70Y/9RB6wn/M
UmN8fRwVECsCpPdFxIR+SFm/nOD9q6BPWI4E5TjTYqWmViF2bO/chzcgLZ1KpJL6
ifv/m2LN7tIqnjgzoSjOR3C+3OTl/0+QdZaSHpji8+i0xodKtSKdHiaaIexK3Qa0
GMVBs3ymCeMr6Vz86ncQnfou8PAW/+D/AAqasWLBcfMw7xjcd75QqlASuC1NBTyp
qzSg1bKpNu3xxqtZfi1mGGgvitfig1BFmN/5Yz+IRzNngjoMHrYmpURdXIcVn4o9
wKylP72CtxCkTyBEcc+dJnC/TiN1vxiWvYNl3aM1qruuAQnTtgZ+1xN97gegKv5V
RaG/jEpd1RdanpJOBds6udnfOyRQuNK0EUvR5mDLgUZ48IwryI9LpqIztyjQIPjV
bTNdi6KNWISBmSC82OEjk/1PlwU39O/muXRKwJnIwN86t86VsudRBof9Wrpe6bnq
m2gME1uB5fQaVgbuPb6NI9tyqx69Pf3HIbXSfwWsHc41AWiJ1LTh1JLC74rWS+jR
CMHeQwri/B0rnEjZZKXvhHqLjqQTjoXnEvhoIjpgvq/Zg/yR1JpHrt0EoNmItyHX
sRmOQx51CkiiVfJvV6/cMHTjtmP8AreLuR0qHCSqJ4QF0a7OWY8oemj/pfZBtnr0
3mDekEWFpt0Bb2phIHXtDAYQFwJ+lco4FxB6KK322Cf5XWmRGNruSjSfrNGZBmkU
oX+tRqy33XY6vnYRbtmPgm5hUvMvEw3qmdX6feFDYQKmEprwJLnoXTyg1ZHUYYU/
xW2nH4qsO+iiaVbQ4rqXzyb5WZEzhO6Vat7mU82zTps45CfMbm5qmLP/Axw5ls77
fw7e2gewLI3kupYO7x2EGe3npF0fiViXi+56p4IGmp51C+H5/c2fuVq524AIna2C
tbXqxZlTYr9u8Mh1iJhiGWmfIXmO5yhe1b6lAO508CrbGJQrsf1pr3GMtNd3qRR1
Gs2Gug+ZsSuIOBRIw0oh2uJMVHijdhJ7Cg4pZRTNdO8MXUsRG4WGZEp5jOtQAJsl
EvLkORBaQvDcWrYsJN4Qxc63j7rOP499RhXSKUodeME+YwfDpAv7At2GgODhjbmd
yfS8K2a11AVPfQWvDcG4xrO03/3OKZnUzNAGLjWFFhMx9untaPrOzIcLDqzS2NhI
pFdBBUAXji+BgZbIET9gR87F4VjHgfwz2PKA/8JBoqZ8yCXcSr5tIUMYk+pjXvqv
xju/beQlHPuFntAyADBeB23AWGp1r2Fge9AUj/Fnxco2WRdFXRwAGnXrOqWjNIqv
z6B4K6iPScB8GWJMB6bpdMKE+qX9ogBmP0WHPTbKQ/3H/5UThw7g3rhzaeSkM9cA
Mhv1FYAXbBGB7FfneFFhfI/Yeem8eW+04wAD3xyfxAJejT4TvhIUe538CV1BHwKz
sSpvZeh59hyC2vAJHuYpGH2f+zibDXQzIlTZ0TG79XRs/KK8gNVq/4qx2HZ+pA+i
ZHKxJEyIpsl5pCOpNTBjOyPizyQ0GtlHa/GOFLovoKgRDeojwmlXRRa2ifusRBk9
Jno0BQkanHcIPyidy8QIQnEkGcYLVc1W6xPDzqVZW8GDCyufoWC6W1yeovLSrrIe
oeWmFWpuH8vp0cKDrZ73HvndVMwa7T8Ty1GyHzBwLxvJapQhtCalgNZ4CWZsNHqU
mt8sstRcsYsPFtwVSNKeCL6arp9nfNvCKgqwW7Z3ZR/rm4FQQ3atup8X5W6Lyb1N
oe2Wr61V+jtgSF1YhnzhlyJJjJRgDHDebKTo7A7A0nh1GBn0rGaI0I7XGrWF1dEj
kNvitHfyT5ZGQta912Fdns9yqrawO4/pIxUa4pQkLZElnZ0nttYTwFyU+iVEGqeN
1xBLsLwL5K4bQaewDiy+djdnFrVUyKHAC7vPwkxo395mnaH8bw57WROM+5TjSUvy
w0+THubvd7jT8AmzxNhiP08yHmY1RgV0JewLO2p3oNqIRi6WGuPWOoqLBYEAEFu/
nq/fPogWq1AQPjZ5EWEPYo5t6jWKWm0WF4ZYwrfbxbx4rLYs1blMPj6qjWqiaH4J
bOHCDgd9/CI0tJaCfxjJV5DPgO+yofcq+Ta7rFS8HfefZNDtYI3dHjyCy/l6LWUV
GdCjQTff+6cr7jRR6kPz+a9oHoqVCS6mnj7IvocWXjVPPNSc1jKcT3+SP2VX3cUa
v28yJf4mfUQrClcTXaCzpbDWYyozz8Zdao0Uv/wBDQgfRypCk72oVOqrYMMk3duB
95gnUDw8ph0cLgwA9iEbMkC03OGqiNo8kR0CjLFs5LEPhMae/XacEvm1B4/IiSZ5
3ew6ygiIzboM2o0zexpD4oa28oE9eahi7nL1KDnJKqJ2tkwJx4xxXc2aFQbwmpM2
H54hwqQbg8jFpUZK9GK0Mllv67FGoDhGnQaYy6DOgQ5XsGs6gncl/U0URUyobpz4
4b8pB1b6JUhhKny/Ux+h2uNNugrbsB06Nf6cBnNuvAu1oeQCnL59pA8SC2QQnUc1
6UrU2IryfNvnDZr+S73jlZMfSCY38dyKrHyEfwNP4La23Q9/K8jvwvBdHYiA7NyO
hiZiVVj0s+GDN60bsmV6I1madISiqsFyl8HXdaW5MRYcs3HZqXCbMeoWevg0n1cF
G7GInMW+ceuo0rxG1qgOodAgit0uhQRNrG/61v4oNUcfiFXzQpNs1o25cUbIC154
8kdlPbvbq6pmjDS5SPq75ADCfUJOTErd3r/9RIAR13x7eTP7/HwUYXbyWt0B3Y6A
UoxoxM0ug6HCuUDcgHetMxKX30A5G/q+5u3x/gZMj9zNDPEUfwB4zzXVx9SjvlOd
EylXH035yitd/vlXAF80bcbVi543EvMAu0RqxeGH2fq2GrAPgfDtVmd6960NaMuQ
kd2FJe0ZKq9EF4SUYSA5IMYAm84bCSLYXUF1qHsOEmnJ393mDdgiGsiUubD0/sZ/
mEXsCfmI7+htUTp0JU04QLhwZT3XVrgb8q8GuhJ0dFLLbr55Dyea5CC5CsyCeDLb
sstyeF2hoVrdwDZznZNk3lYHOUFwDjhWMtr5vU1JnQqgX6GCnPE87CWQfvG3CiPt
PHHz4bn3tmpHzoRFOM0y9RddIR8c6r6LRVNITcIfmoThmhcnqBoAN0z//EU5SbUn
2S0PaEf8jnaS1BSFszno1eC1Xm7qB2EBzPspNd3882BLyv4gj2Vx21V8FsHKVGbQ
dtXPaY0k2RbkzhWbxjbr1H/HxvBEr2cRuKM1HJ25NCdGb8rtudO88z0/FgJkrjip
QQW1aE8EotPCMuQhZw8jEfUCEfsG1un6VFCE+op8audS8t8fqrXv4F9xOV3Mr+zM
m4MOVgYdtbruGIOOYTquhsJytIDEIph+d7msKMRMLUl2mUhBJwcfi+KL1tlJ1BAT
vCXxjjOZGaMoXGUrdsSfcKt6UQjvkYM201JWBAiMy2Ab40mcsFTQmCV+Erz0OaT8
COb1C3veArEbk7NPL2Jqp7lbOSvKgXOBRP1CldLBvRkMLxuurfJYWsVujgVxE5cr
t6Wrdf3ay7v62KFIrzhahsF93iGIwOmO07+h2s47hdZVLL1a6V2Csdph75DmFWcB
vf1y/fkVehxP+UdDOdINwcPsT0VkzeKu6Cl23+dc5Z1g1iAE0K5q5RA9vZQjNyTa
3qRfjDoVKPphBPOjko8cqVO3tbN3FQ8kZDn5sudW8LKfR0CNM58W7E1PA6o1uFJL
5jAyuHBJUoCe+SNhYQ4PNO+kR8Dve/CpH+KhR+ZLi1wlBfM+i9po+2QMOLzILWXO
Fsz0w340X7jneg4MNnMr9oBeB5Ha2XLVll9nkOHnCxamFA7htoJ7VsjyXqwMdbgt
+TVLSec1/O1Od+sQqIH6DjjZRXZlftC2YRuNs9a/8mQyPNZgcg2lfAr36am2Y0Jj
Fhj2VlULdlWn4UoQmFwzaaGdSzY4FklPHeRwu2uMoGZAHdX5cVjH92ZKIRr5LkJA
cAwrbFyhPmVkxGwA0DTU9GLD/6t8WjEqE51bhLzVHMLb2ZGwHxwqk8ZeGtviJC+b
cs107SrqaAOdylZmtTTp5skFwS32wFjDRCWMrvYRwO8CcQCd/+PXIjLrCYfJg5Ch
Uji7UbW6C1n62RuPVQjjiDuPuztYttFuLY/zpIO6JP6wTsVbvst2jWyz4hMKPKtP
E6KckcQNOPWuSLMnMiOD88NXg2xVx/IZrLtMlzqrxzBC7vd4AQVqfiedFyFIigX5
JDZOZ46AQsoLPlssv2uI9rJmiynuboqqWT6YyAvLPt8RUgDlt1BJ6PtJL8EeZ3XQ
nnIWYQDPBXEJoTf5WZFx2TiViQzACSC0VD3+vBQN3RoQa+PNvRprDpiJgQyxNNsv
FpCn/FURJvmyqgn8Tz9mmZ3n+R1FX7Q2ulDtPGP5HkIJWLcxLj89cu+t+bxBOzi1
hIGHvTmhzZp9pvFxI0eZc3Hn55TOY+Oc9Wi0Ojqu5oUdSUMjEdQr9wmi0SQ1vg6s
xUpikyb6/48eut+A6god4A1m+abnRX0ADvXIWT9aNmFjeTTpqVAfMI7Be5xliZor
sUMAIu6Wt3hL4sRsQK98jxiNoS2Yk/pmaILfFN8yFcesSyF9XtPhbaP/Esqiv3ls
X2IVvj9u3mMwHHYzil301jMy70aaCO3jIVlH2jI1+w9aXiaKyNjJ+D2EGbrzt+gm
wbt2Q/mcWX+SMZ1W+bLNMzHGizYY2S0TOiUpoDKLe1WYqZ/kxV3dZxZ/bYFP2JD2
nkq18babvUO0sC9Ukb5rfOmc8bELN2KpKQyL3INhMQhEm3HNrxBgIsKWtsR3DzcL
19JssFrYxOvHFSTv96U1KwnZgnYGRxRZlK9iZWmahxI9r2xUMDpeWMREYroPfLTu
hmLo+BM3CHIf0HoeiDf0ZTJP7XUeQHVRmNO2n2CkS/gArxCT2VzHnQJXVfXTJ017
Drj0e0btkDGM6ecz5m1hFNvSEWE184sxi3Oapx1FjwkIoy5K7wByT/4aCwncYDcK
5hAx6umBVg6FaTvjo89w+eFknJMsYaTwdpQltjk5+8VkOooU3oep5KbRsRoxeonW
X2dWeMqnmybJiatar+8wojoeugYO3IziEv8p1y4w0Prs/HEgzJhxYZHLWANvnP+I
2hfnn3ydlShnm5IwBwtqTdH5hnRn4tfoTMMeHxyIqb/z2BRV9pJ9MOFhD66i1eV5
CtUtXt4OoMNsolPgsbKV7cs04+HXaUb/+LbG+Mt6KrO7oyY0A+3FMLtkBz6076SU
/V1GNqwfxFoebWkhoYsf9DqeS85VimMa1G2EBMBae1rXAQviK0ExMDmy3CxM2Tpx
qwO1VYvZPm2E1aLfS9K2krzzTBeMJzcg58VImScui1zH+KzNCK3uxOTzfPVKnbFm
JU5vMHaQY1kMi5kjtOH151rMBjV4zgqGWBce0SoryJgzjQ2nZ/7sz9awlW0w8x69
BZuPk1MaNLDufwYXdmjtblBuy2YO83o/k08Ytf8jdSd17Pys4PEwIo1c79rtYl3J
/RGTTLuJCbRBk9mNdHnvM1H7wBEj4OcMVxSZPPpHEj+7G5EZx8nu0WyH90PG9co9
w+leLFbtAohz/0IItj29v8fvscMgbIH0Zfsb62RxKQOWSBrAyNAf5QV98h+UKzJd
NNFRim10K2tmt5ni1MAoIyy5aKRPGLA27na1dfw+nwK9LBqShBPLA13qAu5D6Hte
zZ6O/JaP+fme0EqsTxViI3TpUvGdgzurWLEh+Mjtcsuu8xlDMOhFR5tZDqFFlAsK
UkuROJ1qtv0KPl/pEF7bg62F6xY+SELAs31Cxn5yO+c0HaIcJFNthb/9HEmIHvF+
d+iCL6HAIyx9v5AmiI06OmfNZx49g2j+aWSACYcA+fXH2JX0aXaqdlTlMoDcEXIa
8wcOJO6VGRmqpIWrKwUtKsn3km6ScFMJHWauqt5dq2xQSD7eIkT7lSpGggUcfpbh
ayO2UKG69hYzmf7mHQJ+zoIqehGetAwTyrQbPo9RxntJUgwumNwJRrlcrn1/3dVK
6Z33NrNFm9g+bE77RWPk11TAwmiFY5iAQeMFeY8c03FJm7Ydq+07XBbLskX3woa4
Zmhe2tdYkUR3ZDtWv7WAXT8VBpKNjYRJl8vzteC/XiUWcWJdI5D2UcvVWPrjR+MH
zX9RM/ZweS+iSsQrg2FDvbR0TJXqMBbO3j6GY5oHfjI3LObbCsXdMhtzT78d1pvA
2kYnbJdfCvrNskDm2iv4QagRObqeEw40blCVEDJPcqvdKmpP2woCNIXValfOmXIA
nCPFJguA3scyfDjNyER6uki+uo9ks7tfSjVtVxu3Q3EybVc5J6FOYoZPrerUBZOk
h6IcCpUI2rQPv3q+wNNl1M7Y0jp/a2bLwk9JLfJH/Z9pfaacU3PXAgc6IAaoLPjX
yQC1pQIWVWUxnbRvVHuMETOZWTITrjHb9qePv1QvpiVDYPhbwH4fD9m8niXNdnCf
uvGFNIOo5vtMss7+thnMlao120+Ck1v5QklhLjvgHD5ZqQkirMMnIr53mZEjoCwH
GnPoaFzqFY5hfCLb5sZZptvQbvLy8ddLziJucThiyACjiNofmeUuYtMWuT2mCdyM
xxjy0x+vvUTfBdY3V56Omvo/TbicLF1aVjsaBq3tXlSq/DJ7AagDcTfzOLfrSmDs
FbgL8v2nqRKb0hkGJtGhsFPruGVw3YlMQLJIP0Z1D9qbQ7P0B6UszhfweetdNshA
+aoc6nF8jsB3x2ruj/+jt2kmcwA1HfVQoC2LsG+dy6FCFR69dH4b5Ct+PtJLEX43
jB20d5q8muPdCJZM9MbU5E9tVcbRG6P9nAcM81Yak5X4PIKIrq9rIPL5frGIFk7W
vHySQZJ2d2+PQ2XuZlU0eowxc7f48oM7s/TUCmgcpD8wOktK21PZQjkyerdeboe6
CpK2HdSkgZ0AYSggALgTBH8GemDMwZo3Avd0QLjVpDWxRMyYFFeBb8MIuwAcqkUQ
z+Yd8Xd7JjyoinbvzdkcfzxaRd45gkvGkLHmF1PjqQLWCWI9hJfjO0TZLntTIyNr
3XdgKj8X6RW8i73taAtsniGyToXMZIWfp5i1hGG6WQHHpFulqJB2iZzTjSR1knBi
L8L/MTZaY7TcX8e4u/amw9mg0vdcfPd24xhSag71Ly8TdmJ4Y3j/1yWNeB+VoNrP
WLbXCvZ/w2RFECFWd6cNbIlawmqBHarYA6IZ09V++hotTYONcsRxiiE8wSqIbHTO
EW2KFlsLR+aaLTBsiIEw8br1Vk8VGwzUx1afAD1SqPq11F0f6ZLwrRP8xtpIUlZ0
4Nvjd2SJmJ2G65Dsk3idt3Nden2pRXOlaTnUpGChhClhFXIJBikOz0a1C+eOx2IP
o+qsqevKEDQz4V1bvE2714RUswfFry26haBWS5FotaM+hYYFisPvauxxWqRPBrAm
IXhyK1GuRbJ7e/KhyUKAVLtCExGz8m5gQn/iEdiOgiMQdt5A7GW1BV7Aeis5R0oc
A4HSvcCVBAEbCQ+Zs49KxUmfXXBWAwx/6cSY9q7aRqtaVYpInbzD3VwM+nQh6xh2
LfS2IGcDR6cYkjJ9pM7ZyMmgkE5sBXgmUmfgVXoFLgzIgHy6MSDTE3dsOuKUiPz5
Ar3tM0r29p+R/v/DoaE4QZRI/L+fuIG3nHvTfEzavpP+wiOxL0INH62ddxpEmu69
dwVj+u0h7ix1xt8Fd7TMlCAV5l23r4RClFGTzcJokKU+2QmO0+dWqwSQ62RaLtiL
iL4temW/ZiktgRkGr39Lod06Xz6dDOR6YPTvqhvR/QgEAHfxm1LteJA4llbb6UEP
PwhAa7EjHnU9eYGJe95bEyC2YG++x5gqUXo88LjM/Z0WFFmUbg2sMQUKbTDlfj8f
wA3xFl1IxtK4Bz+51i16eNrtUAlffWyA3DGLnns8V6pvguRbBqOcQvTACRC92m/H
M8ezhFG+ZnspfjJbfd+gUYODI6qvwiET6DaFYtyF19S9UhbBPU89NCTdYsqPzQRU
Y1InP9gEe1xEnpMDwoJ9GgywopPvyrdC1nkApNv+oVjWwbFrZIenk479w9mCcn3n
9EzF0eTn5RTDPvk1X6LjZB5srFcRjwxTjDJmdOuiPlt/Qk39FGDtoer6MKIfvRJ9
xr3wr78b8g5fdfWbFOs2mUBOnWzSoto5BqiUV3FxIf0DrD/S3gQFntFD9XYE1285
HlcPTY4yWZ0/HvM9beeh7Mr7b8StGvv5iwvdEYeyfE71K9mhAM2vDLyMpRdpWB/8
SzBE0cxGaMg3P3GIfA5FU5pSSNdeIlyEUpJRGSNA8BE1iSkpGiKL0wma34P/JXzC
Xdxlc1ohoyYsS3W1oUm8MwdztslDclrZIFRsUsCTG6iAY26UWuztetxdkGQafJDY
H9hZMtUlTDuSYJEdjFp2iLLjTQ1ghTNfs10cLspiysdsQ6LjVS7p24J+qQB9zzaL
FZ6LRO21UFb0/V1NFww9Dgh1mtG+v0lklBBsZDD4nW+G293Ovyjyy/in+tvVTEeb
Nty4xXuDKa3uxd0l92dwluxcI+raji6nTBDuQxZ0FX1T7uyDiMTsoGWZbFJBIIM4
WcMRgSPD05kYbpDa8YLq9MFAbLeKwr5wmF6F0vh3eSOxXXfEGjr7/dUj7KniF9S2
iBNi1Ql90AIOoW1MJB8r9rg97s7erBoV2nbsSptT67R6NymIRccMP+C13hQHjyNG
l/3acDTMuF16kZ8Me9Q9ek76NZBUiA2aL3QXaUoUrECC8qBMDrxxh9c2f85UB3zf
BV1xvHOVqrQD5q8Lr4fA4PeylwPuKvbrEKuWUDuGQntrOZ3eRNrgM++okYh8EmFz
8wcy+1suIr4Mc9M89jx6E4ehQRZY4nbbKHNf1A+FkxUmtnFzUZQUdrnwwWsJ8x0Q
0KgTd2gC1ALHxafSFj/6YV7m+t2nYiEyfnNTs+JW1NW3ZmFMHdSm6jP9E75I/lw/
xsFd5Gp1nN5+S0J4RsObeS9wl9pCo0b19os9n/b+QMmi53e7hxC6nbtLFD5/7d9y
SBeLdO3guERTnHJMlCDnA+Pw/yhQvFRysToCjDabNWBMyaqHe9YbgnKCTYKeDlEJ
YIzIZezH/sfEgvQYzUCxi3ZaCdhV1Pn6JINkoPjjwQcoYRBHba8j2K2mX3eU2gOQ
njdsfp5yECo+u7AdX5nJT92KtrBndsx/91QNnypIBUrLDLENIzLdTTRg78TZwk1X
zCsSb9tKsqpugNOjv+PCFIrw1b0qgpbEqy0kTxZomGiJL9q4+Gy4sI7b701H53Wu
DI3EFR9G/azOcHlk7nySaHNh8Cyq8iAqUakCwQMeRo5WfITp0iRTJSXZ5CSZHqDu
ZyZxiTJGr1yarbJvK8/rxhWGWTtSruqyhe8dP/UB1xPN+FWQYGFx2XnLdmEnl3Wt
wJrALTl8VADemznU2RLdjhyrOikHm87p6M+kvGTpQBGTZOH/J0I3wsiBn8ndqZKN
1FgYvCBYE08EVrp/AMjcvn/dF81zMZmA+l8cHaNxfGo0XdFIapqwAnAJvEPNuW0+
XH+U9Xl71KGiNRBm1f3KyeyWpzcL1m2pyu9u0T0ciNyjaT2u9jXj5fdU3XX4c2BC
Gag1fOR1p4Umcrhvrjca6Omu2A3p1dRvSuMBGxdHokuHeuHhzVtAy5t+VNqH/7KU
DlsSwdW3hPmT+G8gfhPCTzymaSV/39Yeyednwmn1q3ifhiz5Egic2bU+GezPUXxG
B30tjLmWn0iLTLbTTKE+hkp0jrLXTVPaYufv82rvE8d7TCniEbN6TnpaDzoFXSmC
5K7y1S+926Xfio9XUYpZU3QHJNjFkiYl55vD0S4ER9yVQKnSxj/vXW5gXfBdjqs2
4hbLP99K7rTlR4XUvKwsxvMXEq+qrzJ01SlSZaIk6wUIIB29ILSn6nKruHdOvTo3
s+IQlT89tY6YOT7z+EAVNilSYB1VNYbouyzrI+MnszlXXeaavn9UH0uEb/8Syqsj
JhbnjCqkuTju7NHksl5e+lV4aYgd1WtvjZUb70ZVl9u16MI79QvPXbIeaD61RWke
ceVRfGkFADdS7ABaklEebJPMqXvmGDw7CKoqiMBc1lYunuMSswYw8gFZdma30xIO
9xdpYEgo5U5s8w4ZFpWJgMoJvx0dK4BXYLIkHoYrgpu0YP52HJzexzGmN/IbCIjc
xmU1MKNB8N9YI0Zljg17ERwKDZReved7LmuNqE7wgBsi0r0b9OMDDYxYQfuujMoD
8GbNB6ENjhwIGU8aUsme7GXi3SRQ7GPH/7MMAgRVn4GzPbq43KjKcxTB77ogWHim
jWeH8vy5JGaIqdIqEedCnPKWMbH30sLnwGnIE8lGvLrDOpP/kc53vkdlSsNawqzF
VgIp7TbMVREyBUbDGo7T5KcQsWkG2kLUpWtyDbnllmtmRsXs3ECuPTuguQWzDtw8
+7OGYMJmYfqe3riQ1odiHqNJ7caczpgHHBdOCQu56DLKIz1bhPXjEfr7dXb+KK5v
qpL7RLaZdlFJi4jkeUG6wLowmqLiZ9HvbpIzm4N7ivpaOfYvlDPE+nP/RDiJvNKB
ivqpWA6Se5VMa9PBHkBRFI7O3IJrqxCCSP3c1RVSf1/8xK+M9UbesEoQbB0Fflkr
+5ygU4YJuabdUQ50wzDSFG/kImxtRogFSNaOl7tlnyWifMr1+wJ2Dt4lIV5Of8Bp
HzEflZpgHwQQ6Ir3an5bU2jku7CgSiu/FUm8BJIUEuNFH9CYlenQxxHF6hjKQKFw
pUjepab5L5311K+MPhOlC0OuQvyNJEzk1Z15uJmbizyinzRIFpV/zq7+HviplvyL
6vm+47hgw+vU3e67/GW1LNYHwOTh/2pHE6vP0DBaDEEi6JcKQM49kIt2OaDf9WIJ
Te+ENicJU5h8jQACqVaj6/gb1NOZ9tBB7WoaROdxINNT0hMHTbA8A1rohjxvW3Wi
6KdQH96CjcZv/xafJGiNfQ5kriFEXl0dJgbaB4+iW+uWWuSG2b54p3E1dd++kL3M
00o0OoIpvnPKEjctUoiK91EWO4KQoA9UC0M5eQ7M1DVZaGli9xK2CD4aBHOtHuvZ
U3PJ6JovA0EekkohQAkpiOb8gg5fUwHDEBn4bcItwLRhdwGQcC7ncjOzptmm0h58
F8Qw6u+GSmFnkisbcvoNw+XOdP6GRj6tajunPBogUrNXqgOjYO4MZvKe8GQdGhrT
fPgsQ89HkQRbzsSXPLDHomX/E7hfQ8PN7/RWhNXHqLwkI8pGJPx3Oy69fPQwrm8O
MuNLZj+/VFZVIKZ98lwJpv12FEGwoGqAeZv1oMbB4TxvrtpovL+pfYVerRii4IWA
j6rCoD8oxsvA8zT0t48LrhBOwdU2G6xa3hZkwUeYzfPQ6pmg1B3oG6tDLnU/m7YO
AREVh4qDsd4UE+3MmQQPaQ==
`protect END_PROTECTED
