`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
L6ZeoqlE/mFaHHey9tXu4065KpqNoAwhpwkPcl+RXHf1Z1EZID7nD4qKhHBFQnd7
4QbCv7y2G8tpLX2KfBARhQrBWrY3GUe7UkMy2tlTGVcaZB9VJ4+nCP6Tp5ky6kV1
4Pv4rcYPfq+1SpQn8s10GvpB7OhY0hUPkwduZ/ANvT1BuabNF5OeAUpaXHRb4Ftg
psHYCFDe6rGE3in2AJk9UjpDib2Ay8XqEvqx372TCzErLxfsDBnJvwoRev5sDIlx
FQdXBkBWvvw/WsWlLT6GznveqyMX4MIyGBhgsDd6TgzmuvKzkdNQ24vlwBNBzUz3
nv+/3VR7m0xQ8zzfqLQdfuNBHdSWaGfCHUY9+vwGefNZVUPxIUKY6cKRrpEnAS99
Rikau8cal20qfB7cqcxhHcwF3FrGd4hju8MVJWN0GMeIKDEirNaI2SoKHPrXixXw
njpkgSEKf2EY1DoAMAon/4LNVfH06pzh/mE1rpBgsCvjFWR7g8A3dsOxORARkruo
`protect END_PROTECTED
