`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFsxZwSsjDscn8TBoFPHVGIOoo4Y6ZXjC2KY1CjdtEVc
IkzUVMqrHLCFVfcMabtTv13avJzweS8DkwlhCOYuGHr4r0iOzXe984buqF/EpE6N
vHXH6k5cqexeFL3DZw28tO88ZV+K+uYwJnYj1v5UBzyFA2Tx0SzJcE5O4GKZVPX5
yPuoxUZbkw56UyyKDIyQ9bVh5eCare3G6v4GDs9sXEwImTSlbaN2sw/LuDmTAQVZ
iScEGNPIrivjAbYYYLTWtN3f4ro0QkOQYctLg2JtxrCL9T3STUvBzL99NLgZBC+L
mTXEG/f27zvoCkIOhcQp0po9adNo3MwqA9Pl1Ny6vsaCZaamG9X9Jo0ql6vVi0B0
m81Gtnl9fMNlUs3VFk4sjlONGuL49CCxQqgo8jcgroY/w7BSNj4ldsUv+sLnC0oY
sEvNaefuYqzLmK8MjVSEux4dJ2z1jn6crbFR0Gs7JZqcvPoVq3UVN24e+dPSuI/u
zVicz2pJmo9Y9plsx1YfQoILNgwRa4OHkoRZt2gqfqGgNcrL5KzxqiaxY3hJH1C6
`protect END_PROTECTED
