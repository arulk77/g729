`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLqck1sDNFOuZiv/ahfGl9M3AkXfd5PNHOpG9Llcsd2r
8tHql8P8LhV0jKXYn4Q099K1Up4+wM9Sm5CBcy1KzdDe93BCb65UdHzKSVYuvORc
ZRiN/KxbAASnFOw0pGeX0UbMbnc1f3mdIBAgu47Xa6fcY0gkcORcfGNHo9vKtOK/
VoW2r8wydzs3TuM88v3vrM+rJvka8gNvGgbTtGXtGAUjs1mObiMIFb5JjuWPD3bL
U0YZbc7Yzsz3q4srJsWL6rn9tcV8DBiwZSLX9TKUACDSdga54dpY37xANY6G3kSG
XrAmVLcWCA+5ByUEq2yY+kE+Yi04hS557eYFh8b3oSvGnMxnXnl3Qv2vtP7j1HlV
p+RC3e7BRCUepoB5SmjdhsmzzLh5ATVY6ZkzgiX8Xd50Vm23CxSK0kCU333cF9ok
w8BlbxKntWw0NJWMp/BV1iprFM3/a4hOeI2SrzzJ7IPiOvfzivIjRoPVq65W5/Aq
yXsvlV84hSc9NdRerWkvXEk+uwLaHcUO3dfwo7GfjMoHa6Ao8QKIQRsdHGgcRsdU
`protect END_PROTECTED
