`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkZ34dauIhPeKRSRNurzcPyGcryclIE3YL8vh5yqlOPrn
QFH+f28wYtPbNW/YaNUE58dih0Y6q4QCATOMnoIhCLElFRWrKwtLG/8HmPZaFcYw
NJDng/HVQvzeb8+ZmEk6Rw82RKfToFdti6CRjWf3AnIl2bWMfXWfZokOaBARJ1/E
b3FB1FIHH8aYtKiJMPdbqYyl+sc3ghjo3sqTXhJF4v/xtGPgc+f7437qqMhchUgX
jQyA0QSSynZvJlKIn3urLpD//gFYrh0Pd0CGtLogwSyZ2S+ttvTiU7kTGF+iBnNh
tqmxdeho4/SfVjoG6EdfTOnxuOPlh+bRZy6ox+HK2cBMph/gTNzle2vj65xMeFLt
ttQpRlD9aJabd59xxeh/k3/P0vTx/HFt0pzYxBtuTGqd6DuZXD61XtbgED3TkM+D
GdhOyt8RyBUCzfMCMMkGHgTdmI8JZWtMYg0nse4NI5m4vSj9uHLUQLOyQEOpJ7S3
`protect END_PROTECTED
