`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1adI0QowcdpONOjOtcA7GgAOcFzvnce4EQo6Ed+FiQs5b
DNFC+Q1WaEyJ4Io34KfRfkqcsceEA/KKHFpCXTd5F0vGzNcEkIYUZcrwU0ikVV1p
35UhBhykIzSrhmlURRC066nAO8J6RdlJ4MjEIWy9T8cIQGMiX+1e5ZlMmc96xkti
vUfmlmMGlxp6RuEjruCKpO289ik/C6No3ywADYDsuE489C40b5mLR9SvxMy3TIav
70wiI23EzT9uFDOsq0U6xUIFz/Bzh/z5E451bKCevtQryxss21tIx0nOEzDtD0iq
YIXXXsnOvox+VePCV17NbvBlj0C/LzKKvV7YMsv/vkts5JCmJb6cSfAj9tR6UuTd
3jwMOs6godDVj6l+deNaIh54zefkF5vV3y/e5gcaoiRBpROtwZO5xYztSWM3ZIwQ
jekDRflmpsMolk10qRRI4vpRvPWnMoh7hs9pQnpvyXC+vUSRBs7yyWca5pbRZRoX
wI2njTG/lFtAMZ0fXPkC9qrwoCLuymopzkuSiOY1dY0281e+uatacu3s4CQKBvLS
9p/plxHiz7QCHYgcJ20+8loYES+GnuTiDhzGrbxffckCFAeRXscbpp/MFdrqR95B
oZGgeUihcGDBzJKkk5fiWqN5iMHSkm88U6oLYjlydiHc/YC38aiUpnxoh6o9WHNK
U/akLV+2ggrUfpSxxy2Vb1ON3Uu9EhI+WJxXVFKDbxaCaTohIbbwcjxJIjoWL35a
eTX2q+5+dznFOASjwLB+fKngwOaz3ovlcCmat9t1OmCcA5vKtswhTuYEuLwSJjJ7
si785Y/aMLv3Y1wahKV+ptH7f3onjHL5gMgM2qsK7Glkzwg5lnB3dnkzdcMwg27q
47NgN3uI+lyBR8HVIhhoXvsYe43EaTPjyw9x+AHhcgRIZKxxyl9pnWf188uF4pcs
L1wgOn6naJSmGbUOV4lJacvS7hJs91fEtjsmuaqAuccnw7W9KaSgpSPgOmVoEoXb
iwtZ/kU/DD1yHImCvSNa1qdlpka4an68DfzhEROcF6MShtwfyZtFxDrCv+D5RNxp
it7KG0erifEzlQ/veJAO8k5urj84jg+gDnHjuH8DI7TyB0XkAAZ16nocFk0zRwPV
RkEFPvnKShjh4WCAtG3tqJkIDGdC9BPa/uXua0nfIBBkrh+OsBPHTiC/fmxO0MR+
zNB0Xd+yF/Ro9BuXW2GX88hTse3PcJHuant6EUJksn6i93DwmByaTwmcNS/uycR6
xHND8Zn5bnGE6zGS3axfu4CHDJZ1a4SmO5tzXq5X7FJNv//d1zOLfwUljFkoGSS1
N56EVl52U7jWIrKUTZzI/p3XRTyiYmYkX7izeUBVLRA3Ylb6Xyr8YYydz4niN4dw
imtN2SZ4gPclKKF5EVsFozjNwF0YJOgvfRRa6DtFHInsMEtZcGBnt3gZjsiGIFJD
mbLT4712+i0KHvjjcSOTgIPZONfxztX9QTH48ODCIe4hpJ2I7t0AHnHZX4FiPUS3
q4+9B5xjuP1MPox6USE4v2vpy8Oz7xozuQPjCEy3CLkyWgJznuskR2CkwdLTAj/z
XhwuM4dbwFBdFQs3VK7wYoNPD+UIJRB6n6kwSuFTKL4V4uGdqf9o27hnGurTaTH1
TKAWQiAnEdpKUGLaGkYv8HCqgjTl1gzRJRkfgRS9e3Q/+c9AvZJsIU3NU7O4/dEw
oROeJo5Gsi2s+dxfAtfbGdN0LYw81sz93XK33UiyPBBaW8z4wKabkccCmqoQDxzE
4ABKm7GITNXlmLxQv3zqhUOKsfDVNWbkE+68Lcpj5bNHXC3PAnSnOzn0Xgwb0yfB
JrwAfekgmxGvZH3pYm6FmRUd3SCIRarVldDAKx6T8H5cB3qvGfrInH7o4DPiuXGv
GxESW0/Neq4bd4P+oox/0VCsIwuFTh7AAX3TiWXLuvxFFioMJsK0dDg9Ugy36FQD
5qV2hz3Bmp8nvsYxWxgUwwhH7zhORdeIN0GNnZcB6o69ZEId81ekFP+mcHp/4Lao
k6VBKmsx/wCWUJMr4rgGDgTy14iPpWUxgGZZ1oIc2lRsJgrp5azoBH9Zzuh464K/
RzaFuVAflU5Uzu46+O7LBtInJGjaVkIfNj1QWEQqVuXeX0fI20TWu1aPnDpekbW9
rutVAEKVFuANMZ+4SuqBnjFC87mhguKq+P8WPGZ/TF+99ZNH9x5+V7L7aFcvZ1+L
Sv5NEdjCsmTB2wA6fW1aQ1FBWHHaWkUe7YxyBcce6qKjIyA8JiylyQG+ZQyPR8iA
oxJsNOnytGG/lD1H2di8dVUiRyW4KPD9J3j3ZyG7yzE3gokuvX4A7MTrV3M6GWYA
45WuNcgFGgfd9IuEy/1tg+B57FocquECdlR5gxLHOjipsjAZU9WLCsG6lT2Q4UGP
nYBOWAMzrEBloog5hDgLj/xGEWWeKTotKzOKMnNi0B24+jV/0+vdOvtxz9xBjNO6
2UcxNmi0mJXrKVvRiooSnGz4fEGXRybGHamChasT+UnbWwXOQ+eRqtcV1HFmGwDU
jYRe0x3u12zMOPLlLhJSO+o6Ck5RPdaqf24XncQPU/NLN59qBHLLwxLhEbRjuVFE
v5vjsa3Ju+TzE2KhDswEW9Tp0ofAJzQcjhp13AMnu0jdZGcFZ38Cez+BO/DXfWfQ
IyGYZf7v80ay0dV5GMN9DgkdUaUuoSA60eD6245HdaCXQioyB6g1+AQHgco4Snc2
Sw5uClN4bUfqORPd1hwz+d6fhvNNa+zy7YOUVZmYFk8uUQKSdgzAM9GPr+oIUChS
yRYqIpCxCzQDtgVN1aJaf8jC/kQKwePp8Bj7NimPUM2YmNf8qr5FXG4V6aXR5Uuu
wikWggEkvCS/uEJCjyahDSxgAlaMGGA8kM8vwl48KJVKy8tIXafYF+VT16iyt9xO
eFIjZP/qRnjxocKi1t456x8OeLLfN7xh1dtALTnu4XtHgYHNGlPdRbTU5PMsfI66
7sD9FyVucnHFWlafZ/3tngZlIaV/EOdqYgMBeLr7ebQOdN6nVfglPvXCKmUL8Gu+
dfJoTehkdh+suYIHSZijHF3kzM2/QOX2MWvO8Rz+oluCk44veWjFv3ZfUdZQ2J9Z
wNgmAKW3eO8/Hsz+YWdkYZ6cKb9zLGgO/Dz3DDaVSeRYIvTC6pqD1WiWK5C+hMrB
EseqgySfuWXR7VZc+Xm96Q==
`protect END_PROTECTED
