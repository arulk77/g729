`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGyq4oGhy6ftb4JfrtljL+M80J7wk4YN0IzuUa7R/VMR
zcSthL4xAi2qttvnlyhQa6kF8+Idfdn18Sm3i+cUPLCXX53gy0rgGDf50KcmxT+Z
oAMrj8tsF+inERPdzpMZvKJV1G7q1o7GjQCoTqXF3vZDL2ZxTN7l5S/PfBmGtwVG
YgY8l8Aop2xHw/uQ1czMWds3Z1msew+24NDLBILLx1RWI0Dou3t7tMkdDRZKf/HT
gqInyU/zG7HvdnS+8Q+xR9uAc12IPgxXlKLC86bfB91fITPGdoTPhPLuKlMb+uZ5
wj8oXzC3cmldgYws35LiGURg/2IO3AzaN25ce2vWFP6Fncx4oT6vgaecxRgTxlGk
Cp/+PPdF+DtvO83HIV6JtjIerEihJ535PitFDm/cxp5yVLgp5C7XjBg1zEfXckve
SEt1S6iOzhqQe6GvSwIuAkUJZz7OEIY50elg5zMeH2EfcoughZNFLXVH3FC1j05x
ks5Ithb3NQf7S9NzyjJSneBeE7hdMrviIGG6i3W2BBiQBXJ4M+Okt7mfUdlf20rD
nFyqFbkwH+pXDVhAKnrOnX51R4lKQ3gNQsttyQ59ViKdyLWz1U5hVPs8eaEqMdw4
Gpr4g7UNkNgXTTa9CSYhxET4iwV2h162G96ncchHMJI8aeRN5shAcjkfJmG6kmyt
LoW1WYoJ/W4cWNt+/CTubU3Gl4EUyq/X0JY3+PRdJOWmRvZDcjk4s1yAsIGlbsh4
7mkg9+a8j7/bYjKXPnYg8cm9dbKeEOQobFDQkSWVpcZZkt9qMfCYrW6O320oa17d
xMVJAUs2jiELA8e1Vb+CSiuMQ8CFucVNAzyS4iTKMmFCt3UntiAC/WhUirzzDe+2
/rgYFe7SqjUIkKutT6cTM23AWGv42stxfVVRHtl/V/oG74cx2CBZJyVQIFiIq52x
9IlsQRWDHccKRnHWzPWanMVXLnbUs1U5cziPy2oRIn/ogIx4ht2d76K9tD1DMxRm
JGXMbcyf4JfB/NAPQx+V5yDYcSuZlg59gAiiGA0ceMdfVOXYsBNSs5Md9/MpaA71
SFZaNPqxgx9dIZm/eLrbHpQHVZVnhupiy+TZkBcNV9gi9Ni7SB3WA+oFNTlotMRD
7QH4tPifKRyfdUplhykHFA5c7XwE2xG4eYiHcK3+jrKRoGPYFMtUVXJReT0BAjmE
usBVDGKeRFDo/4bK7rIZqUIEBo9aexoPvSDMjjHOYr1xqEt6JZBFBcJxKikgjKOj
i5gqEy2ObmyRgFwvEChl3BYYZ7wf+85KSbVOhhhby9Y388SZ3DFovot3ydquTEFW
vLG2oMuTOJsDlW3+4o+F8Egwc3T+1FcNdoDxi2ttteYt2ykeGJkgJeOa1QOhPQdl
V5SxYMrPvb7C1F71Vh/UFx9lU6tOPADSR7Tjn2GG7neCEmNDxlMM/RgTQOkJpMq6
6iMJh3F55vsDkIug57UVAgVwV2+kSpckqZ5ZxE49UODTr6T7POsMLwe5RWEAIEQi
mT49ggykxs3l0MkQCK0gVfigCH5C4rQ/S9Ek9phWBtZW3o/YJAThxTrFqSWoa3uV
tdemonCACBIv/xBaVlUPbpS+AvmFhoqLA2VsDnCTdenROnx0GELHWyfoGXJprg1A
7mtVN6DGSKM8RvFnOXSEoOmcs06QZH15OK40woj6e5uJwUZA/mRK7+x1OjByHQPP
vGG9rdS8R9ZHZkcs+cy28UMaWYipiEoQ+xFJf/Q6gThKCPKhkgaimzkeUI8PIBkY
rz9vQnDR0fjChAn0DxItdj1pfegbzgq4qLIV15g4ZjTUYne5evBJjVKlBepeMFjU
xDXi96WB+iinlEiyIVmq6JWtPL7RlX1S0jwBKd5H9rBs0swTRj2Iztvnqsn6Ns/W
tdGmLRGh6oUBd9d8GO0IVAu5lKBwHsBXk8gtRRLJzarvVr2X9f+AjU4qwjIt5Pp3
Ss+gz0smmjm1Yjtxs83ZIHSgfT2yurShPWMDwsFipC7HcFz6RfVeE7A0LMMqxqXn
yp1JF/KSGX1q+VZotJJE9eCfyxu9YeAg1KgInKy+3zOYAL4QqyX8BPcl6rJ9rhXs
4cZGgYuPKoz2Qmr4O9TAn9MKK7y9iJDoPdVpt4fRYJn8pBGVvZO/n59SadUxyBfp
nDjpn2+9JEP1US2iVcY0zFlvm0rrF1oqqInck893pZFSecnvWnd91pmIZ/03SEpu
PScZWMux+bZfwQL1L33vUyEkKiiEwGSYrOaGQNI2RjOHZMpLTwV1NXpAL1Bdiqh4
kpTEY2xvbKX8cF2zH3WY0ojG6U25VkQi/eKK0p5k2bmKXEGxCQ4tlr7q7JTKAIod
ch4eqFEEndfj8EgKIfAE7y4vT2lWqz3LA7zR+pkPYU8j8WsGcWoQYFgsJZLu3YG5
hDqfkiAtw991XuLsK3awprotP0Ef/XS3gE10oTX/gXA9bMa6K8q5eT+lFi814q5e
WtJVdA10YVgjSMoHCVxvQqMD7P2IufHn+1qfKrqhVyFsyQbYz8mGKDO9j4AO9DAU
uMXdUqxZPkNCSEc1pGUhdaOVdrbVilapbgLWcw3GIjJEbNrXfG4eshz7AvwlhkgF
vAo4raa8bE53J5R97MTs7bHWz3/uDwa3Y6K34ulO7C5woE9mcg0aDRs75Ka0v2Sc
xE8qC7gkh9KdBYfC7OPDAWbvIOh6a/npq6HI4aDMhk+2oqtKhsIDaCxKC1Lg9EYQ
7oW1Ai0XSpRK3M2jcBl5pwX6ZL6BDSGdBCWph8LllL+8TUqP0Yb4UaiCaTkrbFn3
GcWxZSDZRZ92chPU6mgfgLGkNM5UOccJFdFjY2CWUcuiATxGCI3VWUP+E+j8GKrt
YpctDE7dTQZnNGzLdB31w/Q5YAx6En5ljRFg99jtm4dsnvDzvByBbXwtPjzqHGKG
LvzB8G2OlQ+XJxOiZmBQnoCwJ9dBO1rd9yWAlYkAa/3Bhld/8tyoyXSsHz+P60bi
WcjST9rq7O5BE+eC+2+buhhFnK7Ekt09jRLw7hzrmsockleKDR4behvlF16dA3Eq
aRNKdlwET1/eZ6DhYmV49xVVffc6Qq1QyaLQk03VvUQnPSbUZFK0WJWP0eB+W8hF
8PXS6wn8jlyeWbjJqf3b7yYu96aQDw8QeujWF3vgHdShIR7bh2iePwy/SRch0IzF
MVn3mxhCbyn8xdanTICzQZGNj1ytH3mTxdxT8dSW1jkuDAJNmZvvH3oDgikLLGW1
eIlVEJ5Vzr4q6bm+EngLAxUea5F9SYvXKq+PnInhDVDfJNKVpA0S7eNH/SNuoIp1
nr1/nnBZIfhE0mgGsP+JkuagHE0fYHH4WstnWBAVbaJCBATspGLjMqYy699z/2dJ
XaSdStb+5248iMIqZrKAWYzHaS7XAfYdJAb9rWhaVFTcG7A4Vz2+Qke+TfJAzPfD
Bbq6vMXO5riQWrcCqGr/MHQIzG+93mf9tStWFrCXM2h5O3Gpvoj/+I/SClcKeQ+6
9dkrdunw6u1d7tLnTQ7d2TiSB5OGxDRhRJ3/a4FUAQF78Y3FiRWGgrzV7aQ+cQFq
ru1eU1C/wHctblHucDjeVfx65Zyz4GHp6hFITxHavPtNwBaF4p4aAGOOsbncmbRi
WuYIpYjeYOVXOQeO4cokJy45jCIFQXtvh7H+y1QSTNsDN0t0dVcJa92TYh5Us0Nb
BDd059rlBrclcPaCGPkrYGUbUoRM4JKpGO5eIBgAKJJnMZeJJKI28snMJTLg/7fk
69VDm+w18FtAm0RExdW6uz0bbqRDGXhEGCOtQHsOId9ZmVwZL2TaMZ1WNg1Jb00r
Hn0IxMxz7EtK2Foj4RTwJSJI5/jy0umnz9dKAMjtdMaOKBJQdrs2+BzBHRmC7IiB
zEgaz4cTQzQQIK30CIpMAYrW/F1u6gd1GuDWPXza5oJSN1TPl6Fj0csOF5pSL+1K
eiaMBNNS55B54vTcYTL9fFcsnI+GAaY6E8ZPdWCqBNlNgCTyQgO7/smOS1COlP+J
xkUxL4KLvpiC2HEtTNN1P+x/yqsNzSB+aUka1ZOxcHsoXb5Dd3chrmoBlQJI/3g+
JAxg5OUH4Ja5lhTgQ+5758c3/Ts8bnhX49Y7DPX6VhB4CRd1ltJQC3AF4XwJ215G
egaTlvtokj1tQzAohH0WsbwN2cm7PZAwPhwuuWB3BEDEgSMcoQTKawzjlhp5a7Nn
aHTOMurb4CnfQZtJ3r2lXBmx91av0R7R7V5TYVTpPFcqb4MuopfolI+P5ULPtPy4
LqGpiWU8X6ddCh+iDyeZvkBK1VRQXFTONivpstgNe7mRPfUsoCch3L9zvy/7kirC
LPlQT6fXL2Huz4iJ9+/CjJcR+F8FDw7takwPr1xv1esogHM7FMyYJhsOhh5ScYRM
/CruOQymnKZm8tCBzarlTcyAic9Hz8iFwmMakiqOGtCjRs3UpF1q7USWB+82om0C
ErPyU5LKnf/CbG63HZwwMVX5bFvsrqe4yidNdvgumESEhZVxxH+v0j+Oql73c8S8
yMtqUkbKHSxH71crZ6ED7BP+JGfzz+RBC8lDZeAMcx1O1geao41iAd67mkV1CpGr
6evdO3D9vJZz3cvJ7JJGr4dy+jONQmo6zAL11TDbdQEg1Yjq5hd48Fpav6XvLMHn
ichc/n+7PlltxvzculAQbfKJFJskc3+SeEpGm9PD5KCZh5oXCK7MVm3s2Pq0Tail
ml9ReEQrshl2RWxd2kV+epKWve21QK0RszKZIGEaGa8A6d6zs+ymROz2vuYWwJK0
mTQsWCuy0imSvasMBUDjAnncLD+4sZJxXGXxmmkbVBBJez1EhJ0NHyeM7W6bdvm2
mkWht+iaeb3/WAM4fbQiAfMeUYULWYNWlcG2krjVhUZGh02Db7GAyVfgwYpkDwgm
72oCg8wtaIIJM513y6J5e0FRqKOzUlAMtJhlRMihWeo09k0cE3/4zv76zfEEvKp6
6GuQQKFwERuEcAMeue+wH34N5yfmQgntaV9zueR94cPYzYTWgeXrI8LN2BlxBWat
7JrVSHKUEQK5f6N0sxjLaPu9vIgR0AYnl1Siz6gsOEBYWufuDuJ8yYSe2g4TyXo+
MhGpHQqQUC78RfCiY782382xHCwEz6IBG4+yQ1CAubTQVVA0WpIgR3yh+hHEhTJP
zucVmeci0olWVZmZCY7hY5wzvOaxG6Z5GaogDsPPRcxP7PFJTZgIh0VBv+Pd1LQr
CC2L800pcB/AIw4KxJD5ZR2wRZTIAu2KhrNe9+j0yKPxW0YGX5elDtV2xi4j7OnX
/GHvPet/5cTYhx1NwvP6LVP6rQIdafEP88l+1QaXgd1TANUH5he/lwdvlwDRlGqH
bUwLTt2KGe3mfy963+SoNJ4+XDxNtgs4/1capiIeitKQRxukxKdQyUCsTyVgbEy1
sxfM9JVt0ZSHj2JDg9McLttZTZ5br6UODA/jpi1KJQbNHkA9l9j28+mtoXhUYDi3
HGooHiYLp5TlNOGvi+bl229VSvsPnzCL+Y72wTTCSnpdqYg8COMMylHgVQVzsdD6
4piFSm+Ff0P0pWfN/mrs/JRt+KCQf+UJcLthUm5kgIep+n+1RS4e/fjWV8+OgWef
HybWeuQ/y6njbhGZXa1tPjgaTHePEK2twjMXlvxm9mBZV8qy5X/YgMNCMqgGOFy0
UullEr5P9760Noj01dt31pW01EbaYAS5vM+Y+aCYrb1O0jTP1jYx7ADhH78qdwV6
8GPX0tc2Xim+iFNY9IivXxc0tpMFxnR6+RmdkhL8gAT3sz8/ghK8u9kLFTmbW70e
opFyKNMiXi0xkH0yLKL9wIru+RpkKYQMSLcD9Ez0+iI8M1ABwkcQLmMKrydKfDQd
neWrm5CplzZpUg5V3wgpWz2ajskHj2wZah8mCxAEpD2liaIZSuK8KDIeitClBYmq
imsBCVbMV/w+AgQCxAc6inZ1wy07zs5rWTlGPLlCpkk8Dh4Mi3gd+ZaZYeTMQsCq
RAv8W0B4zuulV1CtOgCKXimu/uEXW4fm024joJKu3oqAA9raV1JEzAU878bdmwM3
gWEzJGGwEsqvPYtdZscxpgh+3TYfQhC+2zMUPZnUCpOUio8zVQBlZPe+l3kZWnSy
z55fpMiNDUWua4CbnmPuGrXqMPMI1u3/BQH+5WsA/Xl9J677WHBznTDFjWRydMfJ
KZZmmB4wJ/AbutytmwqOQCOg9y39EkDHdmryj2m4UEcndAJ9sLma8CRuB/Y9upqE
OnuypdNBWquLHqs0PlLK0iwTNKbzsa+hN4Q1TZmNE8hCyi9sdiUR+qthp3Ij+Y5O
z0H23/WsWygFCk6S84+rUMumi3YsEiWkTaHuC/qZJUXSyU0tOeQ+z37NMVP4Owx1
Curufql9esWSBsaFduwzKoAWDnRirD1rER9uYTIIWn7/AX79t1jQu9+MvWDzHRNZ
YXwtcvnyzSaxe1MpU0v4CsGSWg87v71CcROMLGyPdnm5LH5RiQ3B5+rrG1/rZHJh
6PlvENT+NixmHD947OWwmwzApSPqx3ylGsM/95HDHUWLQBkj+hAybrOkUiHUDfZT
qOK1tnGIydKiO7YBRG7UqtvMMynL549f72Ui1CvDhT4nmYXJS8nUQDIJbdXPMUmO
GpSoyyfOgWCyEmNnt1MlqzYdYR2TSukoiOMN+ioQYg2kbMZnygWYyDnWGIE4c9Nv
7ODWESgv8KqOMZMiio1ax4UFVUUVcjR24HnU1jnFGdIaQkwlm3ufcLnMIopBRrQi
osuyd7Ys4VrBqnOs3vG9jShm2EofLZ/OOUi/g8sjQMD4TaBHFdsot8OejU3ja815
6gPuTVSuY8d0QK8mdJgpnZbZSfhRzMFKp4XeI9FGSzWxJQEw+cRxWlga9vTpxaf6
v9KdjGXr8xu+32v4Wz1AbyvHa/kj3OY6/ieLe7Qlf6bsHoD6/z7evchdY7jPLaZv
XwVjHaWP6j1FH/5sE8nN0126G8Cj20YrvAMvetTjKca5Z7R0O61i8vR8JsbfvNQZ
Lp6PfqZZKGrW/DsU8YkNKsjiZWUxwjVuv2W4VmXi2guhMLHfxd6wu1mWNCCwN7yh
R0zWoYEJtQzHoHqwnpfx8TXDDlPjNDezhWtm8CTDfXxMPOzX4iipOdps6rGb2JRL
aS9L7ezBBUgSZVdMcS1IOxxoEkIhwpbfMMuzF2uN08YZtlmGCJtZBsCxoMOUDtYP
t/VBDg7E7JJopHxbTdJy5z8FfgcavLnye0DAorI+BxkpS0pnTruFHe9EH60XZssb
iQv5Z74Bh6h8+L2dFDOBQ8KgpWwUQZ9IzhxK+aWcSn9P8xxO1BdpRX61zI/vWetx
PYT9dooFcHdBVz+rPQKDdsuc23clguHeyiEO246m67J+rr8am5G9C2ORzSB7EsB2
thCiJvc7rVQ5HvxkJUWZ0bKsdFUBC6EjSiMydiFwcv4WATKrDUURd0WebIFmO+Dx
nJuR1ScjmKX3sU+5fzDSirY27qN6SvjSj6dR6yxCFP+1wXtauUUfVpApCYcabHKy
etQesHIRGer7qB5PBOLNujqwtdn/3v90jUUiTX+o5go7fkA9vF26d4MUkamgmUia
366MX14pILrB6JYeM/qjT0D1I713cwRAj1dDixPiatNtpImBg0y6lpcmeZxPqViP
bou3+XQpR9kNwreddgXtIzJiHIPYqSYgbXmwn9gBTzyzv6I2kVgeIQRVhyBmuCeu
GLenmJJZDmmoQC22JoBN4E94qU2E+V++VFeAMxiy5/tmHtj4KtQyz5k00ka+TOvD
sdNPNx47cVBsdCpCrZWhqSNb+ZTxZbQqCYDaiB2P5vho1Xwed8QXsWOv88tOriPE
+0WeQL1STcCvcudk7Pfd8xHSxjjRRX4r2+gMxVG5vGpwM3tBaOUM7hQWb7idbH71
pdF6QZo4nrTv4XOHZ6mBO5orqf7zqHdGM0XfAw8vAOAxVADCrvao8eJgenmzP0hM
g+MjEQ9zHI8BUO1Zd12T48OkbCxdhRHXSl6HzHg86PPsZ3/ZrTLKHv/6Nhiwy2IQ
g8rIRyOX/D5QT0AYL+E0le8Z4yp93ZbLTXXdc6nC/hwngUJsMSsqrgHt61QZfFjd
/LocpTEBtY8kuGfnPKQPX34B7bZsLUyiqZPAqWqaDZ5u0NZV0DKSTLXQdaTg8RWn
OZ/on7URjm9uDnLIw2E4WvNpRsws1l1gqvK/yohymT93OxbKbO12otQ7/l5h7HXr
z4NNGYm4d8KgUe6v1LxyiL01boMEjJpO/PmFEMXK0wRBHSdXZZtm/TJWFyDL7qju
5ejHSA6S/9CJ+QVt0ETPgS572j03jdHfJz+PtKZ8rnD7IfAEV3itaDhrwreyekoJ
V2U/2htYphF0ZkI5nWc/hQLNkHmY4t8CaJUDsrBpp+ENrEQvKOPcir5Ajs4JJv0n
blzgq7D49IjlPIW2umtJ3nq9fXdLWcj632vsc4ksKO1s2fIKSMhOl79EVsFYmS/5
Z6gY95d9oMA7UUGL3+JR7r2Zj+yqa/+VtYCkaIzgrHqWBWNSnh4uHOmlBTfoxCnp
2MsBaD0UJADLjfw65xp05dkhzxbgltNSsaSgjI1MH3NYlpTkaMC6SpSWOpKY6JUN
hk6R/4KO+tOPQGQb6QbOYFLqfGlbvsmR3zYjz9eA8di3DL3/28BAnv6enXxtFVgS
WWF1OUE5a2kqZ4BhUmmUQq2kAD/X4qQufJavrOH/FptyREbgUw+PHBUM/2RK9jPo
QN6x6Mst1GgJ6b5kLQtHtym5ZciXiPN8iCc9saQ0dxnqm79aeVFB8IOX3mHvK6bw
YG9/O2MQ7dEfQVA7pYAcgouWF8F1nyGdKEODm3deSxwMIhqQ2JXiT45VLNb8bGOu
3x89JmC+Q/n3kxFCEfZH1/e+Yrk09EyJ6AEN3rqX4nlc4rnOnEMV8cEoQYVqctjS
bdzNbhnQ1TFcrYOPSQB1tTGZsp4BfsU7RwQCNK9LLBDK196YrYCyeujSiaTEa5eL
BSd4QjiMrg0WmACIaSEtNM+UWgfq/PTSci3315yNCecZfnbMN2JIeuasul8IfkFt
VQU53S6BWty2Mev5bniQBeptUSc7Li7CwGerFm8UOz2OYtXG1Lk2BH5hYGQwzbP8
gxAf44iSX5uO+jTrCg4soXqgVcTxxEsJ9+6OTAdvfnNQSuSPafZifhEzDJvPORvP
j+IMxyX8d+ER/deDozzDX6b9UYxoYqIv/T4X0F+GZdVXhNxmzTlxmzwwJfF7m6og
ZFlC1OmCY3hYs+rVUeLQsjb4HG8pxgle91d+fSh3oMeaXM66PQgbg0gvdHSRwJFj
yiLVYzjuPDV+pYj4q845xEjm+E7LZQ0n5Sxuk6pD2yBV6BxHRbnO/QPOGrXaeZe+
R8U1WgHvrxKkNH14iEzvXL12dHToahT9bOiPMQEd9A5RFzj0wPodaazN5tXlbZK+
M9byO/8dSU6OCMJPQXIDyF1OtCsue8kw5ekBax2wHQlzy/oDAuxj8nPCVD4Cd59a
PElCOHECV9DOyGKzRBPM7t8NW0Skbxehxh6/8Y3SUMqAjdgftxn3SGX2dUVD8T5A
bq8jp1hSKubKa2WClt1+qJ32XKdFlVegawSTvjcv8KkZ6qd4R7v8GZfTd+3HOVJq
RcRCrL66BVwEe57DYoOJu2FkTEuZVOwuAvtwB868wCCYTuohx7VB8mBZYFSMuwk9
DsOHTm96SmgRgbfySumum/vAaOTOTw7v+JvtAyCxfGO21Q5TQ6tdcCdxFooyGFnH
QeYUPHcT8nq4dco7zVYEAxPWHKHo4ij8c6RxB8YrvvB+mcbbbpakHnTqeTIyWsKV
REOMUD2jkdcRPi5TIlXjI2AOcytL46mDHmDN6IMNYn1usjePXPJcW6tlkHPUDrPI
TmpsYY4EQCwZXkzoFAH/hoeWLVxZc73JM56ULAbKdpK48iE2MSt5P8ZkUb5F0DBH
8Xbd1mxjajxSTrPY+MfWHPF8cDYkWECn56rBEHwqVilWk93SZ/1RfE0ujX3JqIMx
pIVaHqwOAwHQ3JXtttVQR8+kqWLjgwQo/nr9lbj5lD5lK49hkjEGrAuzoTSnVqwY
7DC2rgZg2tGvI4QpqT2sYsfRPex0MO6slzJyV2oXTJkZyVOCgwD77/jructziEra
hemsrU12pCK06v+KqWEVCJtY4/65GJUtJHrHauSFd30kgCvcsC88mTCvYLqbGfGl
KSLQxoEA2qLo56iIsymawRgsRAqD2flGD9Ds4PM5m2i8FV0eUECM2DyFPIiOhbvY
z0/e7nO4r7JlXo7jXjwW+PlyuFID1j0DH8HSRPteb8VwlKycJS7JqB7RiaXyVNz9
5hhfyr6zx9wK/79oJHz0wrusYhTBbaUYEOQguhIC6J5pM9gVAykPK/0iZfhPODg3
6u23fRL7Pu5PccN1YJCnsJJQw5sZVrTSF194X9oRDJ3K2j3RSUBoFUvGVK0ZB2pS
E4eyNwUMadXnKudR4BAxSZyHZ4jgh2sX01516L9Qy0tIcQr0OZFbCAadzumQdjKK
Mowx7XzPrbZHPwVC1HjOc1n6JLyOd+qxuOSROWNzZADztcf9UXxAc7vU7rtXYCvg
QiRvvF00vHf033+X6V0kLI2UROL9AM9MhwBndNK39nTN140l42hhLBICE2i9osvq
axM6NjZv0nfje9fs3pkws1vvy5Y+smb1i2PBcmV/0ldWdbTSRasTHHLp5292BXqe
o00Uoo0PUuZelOO7mdjpbQHwcXSjo+3C2HL5NralkouBvIkJ1xSxkuvb4YS4RepQ
i5FTkbJCRghMt3TsKhbKEkzz/p/1c1uYK5rPV0ltlbVhMOl3Fcgsz57h5bsZQfsx
t6ZGv0HyEovmbU7VIeXunGErilKimI1AADvGlORGFQMc/tcGwCEaDBY79R3CI3P4
4mPbnXpGAisvNxrSp7KI1g==
`protect END_PROTECTED
