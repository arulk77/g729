`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
agDLpqK+mpMBQOMkRj+xSv+9D72sdrY2PDGOR7GmyxBBU1FCuWvFsNEyFs3ortI4
X79CY7vklZPPDmLgjOeQvoELYFdsuANo9a+yLGodbvvBdPaRP1QPwsVpA2l6fHo7
Ht9pwhYOvIqUYLfm33Wk6eMG4bC2nH2T3hPrfrWlcsxFJowr+sRZUM/Hqwcz330c
RdQ3csxXSKxlzng5lLYscu+wmIU+zJ+UuTUnnAk28qsOBN4fGUqbR/1rLCupYs+k
LRhy6TSFmfhM4ePOJTUVQMM/8N6yf1R3uN0K8iKZHQsfvcHqBZ268/YB8nIrN+af
0yX7MVJMgUuL8DmHxDc/4O+RvxZOEW27nMWaXk9MFGS8JXc7U2dpHs/t5B2A5SEp
eGQAGnaU6B/Ui6z1YmAGPNgENcd3+3N1xMZrAoK45vc=
`protect END_PROTECTED
