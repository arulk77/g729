`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
hoS0/Dp5EsEZGco+qBTnD7NtsqF8/Ln9D72m7QhsjBUmhvpb9FB5ENOdeJtxPmAB
BJNZ4wEdyTWNNKRymO1ySqxWHkeUf+dJhgI+he/J/2tneI+IHu1odw7KP5Beoo7U
1vzELX3+BxPmEwKq75E0H5Y9SgYP7UWS4j0ZD9RAhd/EyNASSVSEQKSPI9eKUP0s
FloFnkO9MFgBmb5jZa7tLOAgdnBR3f0c/wHVHMydTAN27r19ShrrhElcHiKp5x7y
dOATvQOH83cXthHrItLkTb+dnrjL7a3xtpIwKuwOsBeBULBCg+9nfREHAKwIuArn
esaCmRyEC2hSUnOKdU6+G+pzBgatEgSdmaGA3SbEwv4C8SxiVIlfwsQz7EmEsNa8
Bj8r3UXmquKS9hZe9b3YOLQxRsiWade8dxnhoUYPxO8RJR30+WxfCyE+/uvubC2v
XVQAXvu0o9Zoe3CsC+b7kvkqDXBIkAiypgFE1DyTU+m3kWWeI1h+kPKdZDNexDaH
6+HvemsQoAw9Db5pMbebUWpglJwtWxecNsCpoNsNXO8Rt0ezQSy/T9tFh9pl2wvX
WVM+oxb1NOCqMwSjddUCCP4+0aisDc5+3wOfnybU5lPmUiCxgfXPsT1qvlTndBp7
/ANFGo7h/wJVe0sMCztUYJdyOL4g7zW2NMxXscQnDkqYBqoktEfPeRDeTfH6s+wl
7tQucYMwvh/fdJwrJcamQOItHlH5GkdNNicl0iDhcd68Zqj4gO4OEFs33fK8dWMk
wFkbjqzrOasHsvEvBVYJ83NRXQ/muJKGom9wKCqzSUo+oAGnQiUxSh4cvVN/4Olv
cZ5pHfUJcpAvlkFOzjTkRuNgwD0IWtvxW59st8Q/03OwmW0VBbllouO0WRY3eC5u
3D4AYES+UoxJ0GkukHt+5hW+YW7DjNCNVgnhz5c2g7PEmovL3IL9iJIANp1HMglt
IRW32K/7+w7MRpxhrdpdJPeXQPVPWfQi352iWYD0Wfy7/jL1IlDrLNCutmo9OmIn
T00WcQaLu80YRafLMcYTFzZuu8y56bFncaRNo75IFWYSInh11l7ZE6KV5uVm7VzC
6ftz7GeBnSYkdxaM4Bc7c7Tq7xId/6fXaDxEaMqZIDa70xYf1jKsHfaMVAENTMtY
hQo0rFw3OzT+SFJjbj9+9nhqxqC+ifpg6XcagGAc6C8=
`protect END_PROTECTED
