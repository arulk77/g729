`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xM0yy4mSno2xON8cN+0820n+9Qmtwg5ShthEAIm/sSb
RKrs22oBdsHEAGNSOwEndGYBZAQPK3hL336Mmu4FOm1haBDspQghL76KtxYgS/41
91URuHcP90q19O+gN1Rea46Js5DaSVR4UrE0UnwncEzoiKlptzyn4aso8CQSEwds
iqkbUYYV7bKpmiEVwFDiHO6Hmk0ssgfo6WjEg9wkZK3pC8X3OCIDJCJkAIrYEj/k
5/Nx99zms1cOHrElHapT8qU2ik2MUBflG1fzg9TPmvFXhsvYCStg78YdC5c/OYWF
Nsjelm38eyCaGMRxCHBnvA==
`protect END_PROTECTED
