`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveO618TzBxjI9+gdji0Zg9xDJhXEElMRM2ypX8SJe6Dhl
hlIeUttuJYt2lRfz/tTwe1Ty5igHJ6q5GXx5TUpzZvWv95+P5Zajx/VD4REttPWu
dtyT7xQtl9D8O+6DUEZwj/eWmGCjpwdXI5kUIhf0fzFg9lsylhWT8o2bwTu8LN1W
`protect END_PROTECTED
