`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePhrQJXMxBskCpiHCwqyVNQFzpw6dnPdwwxXgNqdtCy1
iyX4d1p4XP+/lwR5jYxgTAW6Tl4RdwfQ8NuWXeEaJV287xINHDUuPmDGPysRKBJC
T2TVzGSGyfRGRRF2KPRJWaujEHGGB3Oht9XZ/3WbtkxNhCMcensjlIuR2+Gco5Fw
ZjZN7ie06uq6gFi1wHPeLb0fuvlw0Vp+eq0KWZ1xKPun0Y6YbMj4TIQkf6aEivSA
`protect END_PROTECTED
