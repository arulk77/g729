`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGC78jRwDA1cH45TtnCw1eIvN2qJuOLK8QA1xuRoKlNc
5w4ixHa6tZiyNCcVZ1rqHFAYdjzvGltfTRxPPDBxmqWbJHGOis3ijp21Ft1uNHWB
6S3joHvxpddOCsY+Azbt8uMQlGcyRlqSGKO86+ptZtX6KiAEuQL7gMcIrspryGk6
i2PvNy+Euz273Ym/Gx9KxFW1Scx+/xkNpj1/PnfFwAd5J5RGPUAi1LpSve4u0mBb
O44I6hcG2bIoUG6M1A13dPHmsS1LmJNgzqBGtjY6rdfhK12qvcXnUYDtlszqpDnu
TlX3hWvZeqGQ84/CZ7b8ddOMhrMErYR6FesgXzuBSWPk5A8W/tfJpPbMYZvfCcXG
0+bok+Db3nX/eGxeqOnQq+zxFnrwwqfUAstYKvqrB7FkM+j4ao3UowhuVpLAmRrw
1G6pXARzgDQMG2FMGvLq1W/0ElbgWArgHU2UW687us++n2HrTkL+JiLuWfmEV9tt
2WB6T9DLzsxiUaoibU8M7jljHJTaZNC4ZC335m6t09IPn/ABXX9cyABL/LxzoH8e
CXYtfAdQOyCyx2zBwSp31dN9suqaVj4VkBWkJYIAmxXBK6FTbPz7PHsiVKCoyukZ
pf+OaK+XlXo1zvCKK5UB973KPa0OUWWXc1EcOw3yqEhRTmn5u0KEuVaKaDP89gcn
`protect END_PROTECTED
