`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOtZYM9fdjvmXGdaRcHBZ8o0I80G7bUJJoiKbMPb2vj+
ze5KEYlt988lOIJ4UYmZWrPpz6wppK1R0wiq8+/sz5Vda6xnbr9JEgTsx3cwXzG9
bU/4Eo0U88A6RM5c4E5okDw9V78LFVvmXuAM0GQTJlLJOe+lndSzAfOFWTh+cksG
xMbqcwvvXoAK/76w9liGGnAus6JqBhh81bORMk4+gnD81phGxh12PXX1rq0MvsYC
fCwKMHJjvxzGEk6NYPgkiaoT+QFGbUyp3Djyx+QeS+i9xbSGawPP3xkhmBOjfNsU
6Gcj75NUnY7Sm9OD1/UIm4tYp/gWYkAq68jytxRaDHYl56SmJfh9p7aKo+H2P1fn
uAHJQa2dVKsV7/qCtbtnjvZW+faV2sDBlcpCAOXa9b5TJg1rN+c6lN0dmQHvYE3Q
ilGBDZ93pixSqht/aKmBukFATnRbQA3mWkYC6ZjSktm30BgOJOmlpFAiY1CKkv3I
XwpRmJUhWv3M/pPhDvqC8j2CBvWRSeY2S83ZRRwvnPxi/UaI+KF89IGS35HI/MAb
Vh2KLLDULZCQKBGXClzV//09/zmcEPG0TrUbzMD4W41Sx7HQ3Mlu6xEORXaX5xTu
Cdc1VMfbTWOh3dXpqcnxBJHZLsJZ8IBfapTQGqwA2ajiCgfTCiJgpp0IvrDm260s
TmNma8MdP9r4SyAsGQU4/n/EorPgDetsKhY4at64XxjmIKrUGYchrYiJhLVD0lek
uatDp0F2EWVlqF06b5vy9hg1S4L+6CJIJ3nH8Fu/QaI=
`protect END_PROTECTED
