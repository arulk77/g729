`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFfOyBlVX9LZbHoWD0Ovpv5TUm8LiIFaOJTHTjTpqnHo
pLlc90AL+qLfmrBnLLeAO0zGUgJWD9Gu2XP+a1PyN9H8bmwH7XkP7r9pm9L8+Ztx
aXaFAHk4oNw0VufT8iWCcaAgCh15x5VswNztuxChco01k9mEDvNaxjlJSbdxt7ra
z1BxNc9pwcT7S8MzTpH25xxZkjA2Nhi/HLDGLf/FnntFpmtqyXFL32WohNXi45u2
l03fHteBFIzG43whS/EZwzUwYXQi0KQaPIzkrnPaNu+U/UJEXjugJ6VzCKDW86ty
6aC/ed+ne04LWkNXCa2JAQ==
`protect END_PROTECTED
