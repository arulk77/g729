library verilog;
use verilog.vl_types.all;
entity GT11_CUSTOM is
    generic(
        BANDGAPSEL      : string  := "FALSE";
        BIASRESSEL      : string  := "FALSE";
        CCCB_ARBITRATOR_DISABLE: string  := "FALSE";
        CHAN_BOND_MODE  : string  := "NONE";
        CHAN_BOND_ONE_SHOT: string  := "FALSE";
        CHAN_BOND_SEQ_1_1: integer := 0;
        CHAN_BOND_SEQ_1_2: integer := 0;
        CHAN_BOND_SEQ_1_3: integer := 0;
        CHAN_BOND_SEQ_1_4: integer := 0;
        CHAN_BOND_SEQ_1_MASK: integer := 14;
        CHAN_BOND_SEQ_2_1: integer := 0;
        CHAN_BOND_SEQ_2_2: integer := 0;
        CHAN_BOND_SEQ_2_3: integer := 0;
        CHAN_BOND_SEQ_2_4: integer := 0;
        CHAN_BOND_SEQ_2_MASK: integer := 14;
        CHAN_BOND_SEQ_2_USE: string  := "FALSE";
        CLK_CORRECT_USE : string  := "FALSE";
        CLK_COR_8B10B_DE: string  := "FALSE";
        CLK_COR_SEQ_1_1 : integer := 0;
        CLK_COR_SEQ_1_2 : integer := 0;
        CLK_COR_SEQ_1_3 : integer := 0;
        CLK_COR_SEQ_1_4 : integer := 0;
        CLK_COR_SEQ_1_MASK: integer := 14;
        CLK_COR_SEQ_2_1 : integer := 0;
        CLK_COR_SEQ_2_2 : integer := 0;
        CLK_COR_SEQ_2_3 : integer := 0;
        CLK_COR_SEQ_2_4 : integer := 0;
        CLK_COR_SEQ_2_MASK: integer := 14;
        CLK_COR_SEQ_2_USE: string  := "FALSE";
        CLK_COR_SEQ_DROP: string  := "FALSE";
        COMMA32         : string  := "FALSE";
        COMMA_10B_MASK  : integer := 1023;
        CYCLE_LIMIT_SEL : integer := 0;
        DCDR_FILTER     : integer := 2;
        DEC_MCOMMA_DETECT: string  := "TRUE";
        DEC_PCOMMA_DETECT: string  := "TRUE";
        DEC_VALID_COMMA_ONLY: string  := "TRUE";
        DIGRX_FWDCLK    : integer := 0;
        DIGRX_SYNC_MODE : string  := "FALSE";
        ENABLE_DCDR     : string  := "FALSE";
        FDET_HYS_CAL    : integer := 2;
        FDET_HYS_SEL    : integer := 4;
        FDET_LCK_CAL    : integer := 4;
        FDET_LCK_SEL    : integer := 1;
        IREFBIASMODE    : integer := 3;
        LOOPCAL_WAIT    : integer := 0;
        MCOMMA_32B_VALUE: integer := 0;
        MCOMMA_DETECT   : string  := "TRUE";
        OPPOSITE_SELECT : string  := "FALSE";
        PCOMMA_32B_VALUE: integer := 0;
        PCOMMA_DETECT   : string  := "TRUE";
        PCS_BIT_SLIP    : string  := "FALSE";
        PMACLKENABLE    : string  := "TRUE";
        PMACOREPWRENABLE: string  := "TRUE";
        PMAIREFTRIM     : integer := 7;
        PMAVBGCTRL      : integer := 0;
        PMAVREFTRIM     : integer := 7;
        PMA_BIT_SLIP    : string  := "FALSE";
        POWER_ENABLE    : string  := "TRUE";
        REPEATER        : string  := "FALSE";
        RXACTST         : string  := "FALSE";
        RXAFEEQ         : integer := 0;
        RXAFEPD         : string  := "FALSE";
        RXAFETST        : string  := "FALSE";
        RXAPD           : string  := "FALSE";
        RXAREGCTRL      : integer := 0;
        RXASYNCDIVIDE   : integer := 3;
        RXBY_32         : string  := "FALSE";
        RXCDRLOS        : integer := 0;
        RXCLK0_FORCE_PMACLK: string  := "FALSE";
        RXCLKMODE       : integer := 49;
        RXCLMODE        : integer := 0;
        RXCMADJ         : integer := 1;
        RXCPSEL         : string  := "TRUE";
        RXCPTST         : string  := "FALSE";
        RXCRCCLOCKDOUBLE: string  := "FALSE";
        RXCRCENABLE     : string  := "FALSE";
        RXCRCINITVAL    : integer := 0;
        RXCRCINVERTGEN  : string  := "FALSE";
        RXCRCSAMECLOCK  : string  := "FALSE";
        RXCTRL1         : integer := 512;
        RXCYCLE_LIMIT_SEL: integer := 0;
        RXDATA_SEL      : integer := 0;
        RXDCCOUPLE      : string  := "FALSE";
        RXDIGRESET      : string  := "FALSE";
        RXDIGRX         : string  := "FALSE";
      --RXEQ            : integer type with unrepresentable value!
        RXFDCAL_CLOCK_DIVIDE: string  := "NONE";
        RXFDET_HYS_CAL  : integer := 2;
        RXFDET_HYS_SEL  : integer := 4;
        RXFDET_LCK_CAL  : integer := 4;
        RXFDET_LCK_SEL  : integer := 1;
        RXFECONTROL1    : integer := 0;
        RXFECONTROL2    : integer := 0;
        RXFETUNE        : integer := 1;
        RXLB            : string  := "FALSE";
        RXLKADJ         : integer := 0;
        RXLKAPD         : string  := "FALSE";
        RXLOOPCAL_WAIT  : integer := 0;
        RXLOOPFILT      : integer := 7;
        RXMODE          : integer := 0;
        RXPD            : string  := "FALSE";
        RXPDDTST        : string  := "TRUE";
        RXPMACLKSEL     : string  := "REFCLK1";
        RXRCPADJ        : integer := 3;
        RXRCPPD         : string  := "FALSE";
        RXRECCLK1_USE_SYNC: string  := "FALSE";
        RXRIBADJ        : integer := 3;
        RXRPDPD         : string  := "FALSE";
        RXRSDPD         : string  := "FALSE";
        RXSLOWDOWN_CAL  : integer := 0;
        RXTUNE          : integer := 0;
        RXVCODAC_INIT   : integer := 640;
        RXVCO_CTRL_ENABLE: string  := "FALSE";
        RX_BUFFER_USE   : string  := "TRUE";
        RX_CLOCK_DIVIDER: integer := 0;
        SAMPLE_8X       : string  := "FALSE";
        SLOWDOWN_CAL    : integer := 0;
        TXABPMACLKSEL   : string  := "REFCLK1";
        TXAPD           : string  := "FALSE";
        TXAREFBIASSEL   : string  := "TRUE";
        TXASYNCDIVIDE   : integer := 3;
        TXCLK0_FORCE_PMACLK: string  := "FALSE";
        TXCLKMODE       : integer := 9;
        TXCLMODE        : integer := 0;
        TXCPSEL         : string  := "TRUE";
        TXCRCCLOCKDOUBLE: string  := "FALSE";
        TXCRCENABLE     : string  := "FALSE";
        TXCRCINITVAL    : integer := 0;
        TXCRCINVERTGEN  : string  := "FALSE";
        TXCRCSAMECLOCK  : string  := "FALSE";
        TXCTRL1         : integer := 512;
        TXDATA_SEL      : integer := 0;
        TXDAT_PRDRV_DAC : integer := 7;
        TXDAT_TAP_DAC   : integer := 22;
        TXDIGPD         : string  := "FALSE";
        TXFDCAL_CLOCK_DIVIDE: string  := "NONE";
        TXHIGHSIGNALEN  : string  := "TRUE";
        TXLOOPFILT      : integer := 7;
        TXLVLSHFTPD     : string  := "FALSE";
        TXOUTCLK1_USE_SYNC: string  := "FALSE";
        TXPD            : string  := "FALSE";
        TXPHASESEL      : string  := "FALSE";
        TXPOST_PRDRV_DAC: integer := 7;
        TXPOST_TAP_DAC  : integer := 14;
        TXPOST_TAP_PD   : string  := "TRUE";
        TXPRE_PRDRV_DAC : integer := 7;
        TXPRE_TAP_DAC   : integer := 0;
        TXPRE_TAP_PD    : string  := "TRUE";
        TXSLEWRATE      : string  := "FALSE";
        TXTERMTRIM      : integer := 12;
        TXTUNE          : integer := 0;
        TX_BUFFER_USE   : string  := "TRUE";
        TX_CLOCK_DIVIDER: integer := 0;
        VCODAC_INIT     : integer := 640;
        VCO_CTRL_ENABLE : string  := "FALSE";
        VREFBIASMODE    : integer := 3;
        ALIGN_COMMA_WORD: integer := 4;
        CHAN_BOND_LIMIT : integer := 16;
        CHAN_BOND_SEQ_LEN: integer := 1;
        CLK_COR_MAX_LAT : integer := 48;
        CLK_COR_MIN_LAT : integer := 36;
        CLK_COR_SEQ_LEN : integer := 1;
        RXOUTDIV2SEL    : integer := 1;
        RXPLLNDIVSEL    : integer := 8;
        RXUSRDIVISOR    : integer := 1;
        SH_CNT_MAX      : integer := 64;
        SH_INVALID_CNT_MAX: integer := 16;
        TXOUTDIV2SEL    : integer := 1;
        TXPLLNDIVSEL    : integer := 8
    );
    port(
        CHBONDO         : out    vl_logic_vector(4 downto 0);
        DO              : out    vl_logic_vector(15 downto 0);
        DRDY            : out    vl_logic;
        RXBUFERR        : out    vl_logic;
        RXCALFAIL       : out    vl_logic;
        RXCHARISCOMMA   : out    vl_logic_vector(7 downto 0);
        RXCHARISK       : out    vl_logic_vector(7 downto 0);
        RXCOMMADET      : out    vl_logic;
        RXCRCOUT        : out    vl_logic_vector(31 downto 0);
        RXCYCLELIMIT    : out    vl_logic;
        RXDATA          : out    vl_logic_vector(63 downto 0);
        RXDISPERR       : out    vl_logic_vector(7 downto 0);
        RXLOCK          : out    vl_logic;
        RXLOSSOFSYNC    : out    vl_logic_vector(1 downto 0);
        RXMCLK          : out    vl_logic;
        RXNOTINTABLE    : out    vl_logic_vector(7 downto 0);
        RXPCSHCLKOUT    : out    vl_logic;
        RXREALIGN       : out    vl_logic;
        RXRECCLK1       : out    vl_logic;
        RXRECCLK2       : out    vl_logic;
        RXRUNDISP       : out    vl_logic_vector(7 downto 0);
        RXSIGDET        : out    vl_logic;
        RXSTATUS        : out    vl_logic_vector(5 downto 0);
        TX1N            : out    vl_logic;
        TX1P            : out    vl_logic;
        TXBUFERR        : out    vl_logic;
        TXCALFAIL       : out    vl_logic;
        TXCRCOUT        : out    vl_logic_vector(31 downto 0);
        TXCYCLELIMIT    : out    vl_logic;
        TXKERR          : out    vl_logic_vector(7 downto 0);
        TXLOCK          : out    vl_logic;
        TXOUTCLK1       : out    vl_logic;
        TXOUTCLK2       : out    vl_logic;
        TXPCSHCLKOUT    : out    vl_logic;
        TXRUNDISP       : out    vl_logic_vector(7 downto 0);
        CHBONDI         : in     vl_logic_vector(4 downto 0);
        DADDR           : in     vl_logic_vector(7 downto 0);
        DCLK            : in     vl_logic;
        DEN             : in     vl_logic;
        DI              : in     vl_logic_vector(15 downto 0);
        DWE             : in     vl_logic;
        ENCHANSYNC      : in     vl_logic;
        ENMCOMMAALIGN   : in     vl_logic;
        ENPCOMMAALIGN   : in     vl_logic;
        GREFCLK         : in     vl_logic;
        LOOPBACK        : in     vl_logic_vector(1 downto 0);
        POWERDOWN       : in     vl_logic;
        REFCLK1         : in     vl_logic;
        REFCLK2         : in     vl_logic;
        RX1N            : in     vl_logic;
        RX1P            : in     vl_logic;
        RXBLOCKSYNC64B66BUSE: in     vl_logic;
        RXCLKSTABLE     : in     vl_logic;
        RXCOMMADETUSE   : in     vl_logic;
        RXCRCCLK        : in     vl_logic;
        RXCRCDATAVALID  : in     vl_logic;
        RXCRCDATAWIDTH  : in     vl_logic_vector(2 downto 0);
        RXCRCIN         : in     vl_logic_vector(63 downto 0);
        RXCRCINIT       : in     vl_logic;
        RXCRCINTCLK     : in     vl_logic;
        RXCRCPD         : in     vl_logic;
        RXCRCRESET      : in     vl_logic;
        RXDATAWIDTH     : in     vl_logic_vector(1 downto 0);
        RXDEC64B66BUSE  : in     vl_logic;
        RXDEC8B10BUSE   : in     vl_logic;
        RXDESCRAM64B66BUSE: in     vl_logic;
        RXIGNOREBTF     : in     vl_logic;
        RXINTDATAWIDTH  : in     vl_logic_vector(1 downto 0);
        RXPMARESET      : in     vl_logic;
        RXPOLARITY      : in     vl_logic;
        RXRESET         : in     vl_logic;
        RXSLIDE         : in     vl_logic;
        RXSYNC          : in     vl_logic;
        RXUSRCLK        : in     vl_logic;
        RXUSRCLK2       : in     vl_logic;
        TXBYPASS8B10B   : in     vl_logic_vector(7 downto 0);
        TXCHARDISPMODE  : in     vl_logic_vector(7 downto 0);
        TXCHARDISPVAL   : in     vl_logic_vector(7 downto 0);
        TXCHARISK       : in     vl_logic_vector(7 downto 0);
        TXCLKSTABLE     : in     vl_logic;
        TXCRCCLK        : in     vl_logic;
        TXCRCDATAVALID  : in     vl_logic;
        TXCRCDATAWIDTH  : in     vl_logic_vector(2 downto 0);
        TXCRCIN         : in     vl_logic_vector(63 downto 0);
        TXCRCINIT       : in     vl_logic;
        TXCRCINTCLK     : in     vl_logic;
        TXCRCPD         : in     vl_logic;
        TXCRCRESET      : in     vl_logic;
        TXDATA          : in     vl_logic_vector(63 downto 0);
        TXDATAWIDTH     : in     vl_logic_vector(1 downto 0);
        TXENC64B66BUSE  : in     vl_logic;
        TXENC8B10BUSE   : in     vl_logic;
        TXENOOB         : in     vl_logic;
        TXGEARBOX64B66BUSE: in     vl_logic;
        TXINHIBIT       : in     vl_logic;
        TXINTDATAWIDTH  : in     vl_logic_vector(1 downto 0);
        TXPMARESET      : in     vl_logic;
        TXPOLARITY      : in     vl_logic;
        TXRESET         : in     vl_logic;
        TXSCRAM64B66BUSE: in     vl_logic;
        TXSYNC          : in     vl_logic;
        TXUSRCLK        : in     vl_logic;
        TXUSRCLK2       : in     vl_logic
    );
end GT11_CUSTOM;
