`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD9I3EMdJ9+y8UfKfxRf0ceCnKU4IKo5QsATSJerpYqE
KCGH5ada+hdP9IvgyV1ZEmX5UXmTgUnRtQO8pCibUXtEOJWhOf7crF+oRkMLLKiR
HZQYyaHr/tDPQXVh25zlk05HK2n6ajmo3UgvreqKAwYXiwX4bnGOnW2F7xoW4iiO
q0X2lmrd2M8CL+7H+EmXPzBtdcJghhJJdtwWGudR1ygmLiQgVuGSUKVDApADKy6m
qQzpiXbcCAFMYyaL9d9oZsXQDV9xO4JCztB62gKJ6aji8U2H3B67rI/kTVDYTqSt
xJmvPInSv/ptJbJ8Ofq8OWgBwtO7XzVELfjiYPLhGVAc6twYxbTpddqELwH0Oihv
`protect END_PROTECTED
