`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47MhCdTnaddBDnrTIVaxztTwbMXpMbrLcYi90KGkZajv
o24wKxuI0EmLPGXmHblIiGXjKsfl+aKBiEqXDT29jFYiffJrYajXZt9pNJWHRJRX
t/Ghi0mVPrVbWFRBj0HnZwpAcbvk3jCWahbC3p5wTHo6PUOsTDNlmDI3XPxeZxpD
pK+5/RnMr2Nbgaw35B2hqwEnsNeD7Vv+8v/8lVGVcd+9xBf4Bedcb6dfD8XWVN9S
NFxYoYb5lSPj0kJlvJUsx8eeYsLsLYlM07GSeT899hMFqthoV5ttwNpvEZNa8B1O
jkbQQJNdGHeoFwBzjiJpv7X5RCDeUrGV50YVbK282DS8le57JPHn13XFlttd1S+o
Ay3V8qBL7fAh6BwU56xAhA==
`protect END_PROTECTED
