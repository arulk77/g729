`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
FQ3Qcmh9uMITco7neeTVUzfLvqJscWLOc5ga4YXG0ZZYBrSn8GjPY8AgXNd1/WO+
1/KEidpXERfT2wa7iHh+F3QwnxY3wCg6/WRLt1JN1OOdKxi4z0A2fV/hvjqaJbra
U7Mxw3mBVS1vj/YX/GcsYFxmxl2sa+qzyyajjHJ+SS/wfhi3igUtoaWcHkO2+is8
5GNz8TaLZVGsrfl9U35ItpSKqJU///X2xeOoCe8jlHE=
`protect END_PROTECTED
