`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKSJ6dprDjIKFzR9efOy2wfZROuvT6GyksWszYf1/C1M
luKww5B+LvEr6AAdlCVmStLRupyUMmv9oknNIf5o4qh9hriNDV5vzSgMpIM29I6I
BBfOhRTV4HipSTWphwUUspoowku0dzotDm/02jB7xxn2KdTndNQvKYg7g2gBVMbG
jvCqzmTG/lPwTY6bhQcCzb9Nry8A1KQGtFujo5Ina2z3j1cv6pkjNPCeKRlR2+c5
dAIwrCXl27eJiPlMD8g2bMxfQ7JTgjrTkc5DLRAVRTeawVy3vOjiqxrXfW9Y9HV7
BpenDFb4gf3kHVeBcUndSA==
`protect END_PROTECTED
