`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAQWwP1S+Y+IKW2BedNSjy0qSVV6UA0pD2S58j1RvgyQW
l71x+xnEwYAaHeZN/SoPlOU7XgXUmE8vb6LeaZpVuhVLEQCEyN9AYFTUo/hoI/Vr
dJTX4V2uw7yrPqIJOyRoEfOmXC6U0Mtx7LFGUh3jl2FDfPOFRZ1+1OFzpdL0u8RO
OiNNRBXe1CtAj+f/WIBj5K/KDgvfQFD50YMGW7KqkA5N48LnUMNIUyyadmcXbvIn
iTAtcPAnd2YtN8iu0CYVBTHrSa6IKJXZkOH9ZWueqbluKGgO4Q8FRHFWf2sOUf54
JiB2BckpGz+Q4y+gYaWv8uif3InCBGUV/3B52HQGefG/0gBYvFqg3eWsvyUM8Els
BaV0kp3ScqJF6NO3plJcPO0HyI/qFgQ0vqn41PhApMSF0eovRnCxGrXQF820hCHB
J91bEhk0HsVcJkDGTYftVJJP2bt/EtZhjpWtfkglAldQKbKmgFWh989ACxjEvtT7
RiOz7SLmLkxRmSLHnxvsi8pxcnAo63KYaA/64encxjUzfEcXZTL1CCE0aUMztN3G
vF67hpqWVVxakXCnhdwpjw6LFNOoAZBwTzm02mqrWNHtzJmEjrCsxUwYGkWso0fH
G0Y1i7n4JZ9pCzi6ULooP9pHOLFTzgbwcB2fEnHYUA9GkdyVYEiU/A0hOM8XgSJr
a70x2im0IAyJtsvEIOLf7myHwc8qLiVAaHan92KPTX1t2jeO+a+GTIDeXMdgjj0H
gFfjOv6Wf7BPp4dx52OPZLZLdskfiZ0BCVGWZqYEyDgT+jbgzziLDaBy5hrVsiF3
a/AFOP+M2Aot6iRVCNsB3wr/ZOA1+oKB1GtgPupi3TnAU7HpjnCojHSr8YPC2At3
TeG7Q01EVdJRURqgEUsCxOi5aKQ7jShCIqmeMLPQPNOm7y3Zew8E/kil/TyhIZF+
ldimpyghbU8H24T66Pkn6fiaX3AzTVXw512XyG1y4jq2g/cjaI3F2diyQPzPpU5G
Z3HpwJ13LW8z6eYtVXzeiakXmDcJsVstxpiz8gxKyTT+1Z6RFCeD4ICEnatA1ofM
JYinYYhBODr9g0AawE/h43lpEO92VT73hzOzjn05mfepBwtsI2ymw+R3ABMbV3Uw
PP78P/W2jrYttBnHluFeNkQHypkk7Ug/y8xRXk1ntIAU5hrASRSHUB1itb44gFGm
5HlR/YRuA8mT1nVJmhju8AsPFOeoG/E+paE1cPpzEoytgnHfA995yz462GoAVQw3
lAQeuV9CCi0C0blEe3u6Qj6Qy320E/omti1T6YCMnE73u4OTG1Zpri16i8lNKzrB
Chdcu89cacM4v0miQYXQbEaieV69blVWZ84xBeUVYqyAiV5oASb/WxwLoSMsHo2T
d8rtHaTPWlAaWE1Uhf2FMlQeXbWU/rwbLjo0EEPwA1HJSNAmM7pKoJPU0R/EDGtZ
IvsTsaBvbKorcNIKm2g7OpO53nuULAXTkPM40yXVfAz7zfNcp0a3n3KuBrZKHu41
kxW2nB7bQ9i9iE0EMO8F5ZpLCCu49moWyDs44UCHDJC9hzmCx/v5sloko5kKflvS
Fz+14dAYabWLRy0+jkZ1Q0kRB1r2IB3uZxJKQJUKkxiGfMP6zM4a+7wMKrJQfPbd
7EFMAkNmV/4cPUcBY6Lbpx0UOHfgqw47tMLCBO7XBtUX40j5rJYsfHZuYp6tMCCc
bEUbhsMhn4Fw1yjhLKMghblqvEtjBirsHUzt+F429DpGHx8WUktEkE+EsueAapEc
U7RQS+V9hmxKJmYMepr9HLjTGz9wCdNt+AjCwBx3TXWVq/Tt1PRNJXPlGTq1sE/y
4qKuuq7UfwLhJuriqMNkqedk/NLczJt0N6ScF61O0wKx6DSby1QULRndTCGk/SUm
nk2iIY4Ii7Ebglxde1VrGGkIpKZle4HLgz77jqtX/XQ+mc4uU3KMYDuceQYv3QiI
K+ltJcLe3tBeUkt+mE+Kv7oTlfaovSeUGNouziCkZ5HFayBbh/hXVo+gE9mcCABe
v18PRN+0aWPe0MPH/ezfUr65ZkhyFSgSuV7wb6i/CsyhjOMSAu2Tz41ncWBT/X+J
`protect END_PROTECTED
