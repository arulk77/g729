`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46e1vsqubSKhanBzucQGr2qp20IeptGQBgA18Zg5KvAh
KwaRlgSVQIFt2EHPxQMVqsLs7/aRlAWvw3OjMr0iBbl9ZvBvcmNHkEjWPV8AppI1
7DzoH/EQfsyqYCCpvis6kpJ4/6FCVEEBidiKwxjg8GANs2SodV+QsIZo7dcAjaWL
OTDNt5KnMCCuJ6aCm3+hf2MjZc/FuHLPEnpeuQ6icibeJulir4S/sSocJ7g8DBVG
z3G+y/DqqsfYs1zyfYLOlqbpMRfukr6n5OJBSBJeVn+YDblSHjwr1kzCTJWoXyOi
lRS0OIGrs0Jds00e5ImcF0w+RyjhhK/vgiztCVUnL2ZYejCrGZc4NojNyL1VCoiT
e/5ZRQAvA+xtLBZnpDPPm/0ET1Rpduwh9emo+yoEbAicgGV1WNtFlzPOE+H4/Fl0
TklgmXmCgZyzsuMq2s0xd1c3RZN3RwX4xJ/GfGRhYPKzwoF1q5x9ryTk4IVDMOU+
`protect END_PROTECTED
