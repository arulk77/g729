`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4z0Q1oZBeA6+8sqclHqkwDX8HajOO6M5+W2wsX57KI6G
04baKP6TFCLRnaTR/kEW621ibqikdi7aYpJ7aGKSO5XCVznJjI2yDtKQ1kLjfFmV
DVgyQX2XeEQZ6kdCaZN1bXF2nG6vISjXToG9Wua5Zub+BQ+cLi0//Ne0MkXXwfeM
avEY5ou9rh6sug8ZFDB7F3rtLq8ueIIJRB2R4LTaKOWDz27TDKvn4vExYgIUKAxD
o5xIYpQnbIe9IsNZLRbsdeTBVIirAPDn+wjdV4u1DVu5V5wowyTpQ3QC3na7fsZr
sMeTolp2lT4YFZxpiIfjO2bjd24XCDeTOM5JpFV6gyzfUhnG1/ubY8MOhTJYB2FI
CT0TBy4nk/1obTqSOsvINw==
`protect END_PROTECTED
