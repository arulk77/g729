`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNav7so+7hVE/zhPxv5EQmhZnybhl89bAkUXXmpvE6/d
wj3Z/9+SxYRCokvIvkRrP+eof/uqbvkBPvL9RVJYzS2jFfbKtc1RXaLKxLoRyOtw
rzmkJkj2AZYL4C813X+GWWYNO5CA9k3DinGEzC9vC2Zbrq+cckvyjaNz9ue0hPns
x2X3i2o5wJR+C11HAUklxER4rQwan0mZsGz2ob99LHlKXK0dNju1ECZfS6c3yNJ/
rpT4M8Cf/iG8h+RiDJtYhbl2lp0NcLQE0wXjM30c4OCVJaiu2SM7wWgLxxewMDl6
7d4zSWUklny+5Jd2tKpm8rIzypyVTQGijbXzX9m3TaS2h/NWOm2ohKfJHkSgRPkc
tQjIcs7T4Bo5GqbK+uafv/5EzucvVOUQwwmD0WlNM0IxMMCcH6lHGg+MMTky8Kkt
IrhuwLKw9lQy7SmLUYJfetwF3PBQVW9urGjnW04BvqQt/m+BzIkQT83tm73rHH4X
fUrOTR5p2ChVLAdRvtW1tt9hrodrV2GBl3gv2UOMkBeGfA1u66AoNjWrTu1/7prm
`protect END_PROTECTED
