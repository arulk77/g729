`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
fqIX4MpAYT/OD5N3OSEnXSeIY0x8fff1oWHOILgY9vf9ziU3Ikn3DZb6VWhO/pCQ
sKAM6MN6HEh5U6CoOt0YBL4g+2v/QUW1sflLUrhRbr84qgvvSkRlhcaH1gi1liHk
vXNrLCk93ELtNzcN5ERx/rZy1nkMxt5oyk1+Fk0as3PS/FFrVv8VerXSTGwN5aOa
PSYiwEqZox9TqFj+pqs6VQIaUhUsV9mmV9BDgqzwdqG38o0L3cEI/hl6g1uPe1h5
78/Vyx06uxT5OWRhTFqDC9miXL9pzRI3PAJqync6FKzwvCI9HImFU9vh+aE/23A4
tazOscg27mK+ssr+JqQeNIqoHP3GQF9GuJoi27BPkRfVIAMHUyQrzY2Ohc+kgwAw
RVUVO8a9iUJtpfPFzexwr4nRxqo0njIVyDsH1nQCtT0=
`protect END_PROTECTED
