`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1afyPjK79v5qM34Epa13CfWBQJmh+ttHaadUAsRJl+TnH
+2RSZ5TvpVDDZzrRw1cINm6PDnYc6ZKgF5RLK5hgg2WSXmZ18j2NfbXc2qNbcDR4
0VB53qc6jeA/cAvB6tZBhhr5KXQ8OQAbdfQEBsSIPUNKkAABik/pB8D9rkvAfkyu
tcQZ+RvGeOCe/fKmazIZlPFn9/wU29/48x8RXxOW4owdGltfHyEwHWiVcFUp5wS4
/lDvV1yQiF6bqQr3oqouHmHOpo11YFMx2x0d5wTS3JmG1ynGrTdi5w+gsOTPUrL+
`protect END_PROTECTED
