`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Cf/a//tFpkW+5T6Wvk436qU+svz1hZkbYZ6pm0E9QVVlIGxeYJGbluIWsvEtStYx
YNDBCYkyFGoHH1VqZaqqn1qeUjXkU1008Sxgm9Uw237jrhvmQxq9wU4v3HnUltii
B9dVEdKkCkGRXWU5oB5PPtnUpU1Ikx6hRIvMBkhm6PyKj3cUbpLA9dRh3WOUxsn3
/eJx2lQf/9ebtTe4EUJg8d7KA/f4BQX6nop5ez+UXAu9gPKE+jaaazy0b2mARM8M
zHaHVtbKsvppUiOPWMq2ool2Q7r13y6qcq6Hgo2SK1g=
`protect END_PROTECTED
