`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEXhybw7tobY+yEKiCrzefAiEeagFJtUHfJ2aXHEcqpO
WywbepeR7ZCon/wU+Q+K2GQbDlzDNrPW6Gue+1AJ45SG3ndf1KWixNHIeitxe3py
1B6vTaCNdcz8u1glwzX4TVRClAh5awyJvOz3sBP6mc5dgI4L3vri7ZOU4B2rejiQ
7TiHoAYAFW/mSFgSegimmoPGKCPrxGB6n1Hxxaj9BIqmTcyGi+mL9p6kOmymN/K3
l6+4DgTXZ6+tbMr8TnC20xjkacIyR7ZuukiP8yqnxvmH6GrT6QN5bwQdHMlKOq9j
jV2ppKFxSxGvQsPigTLDGQT+keeaKuu6SP1hTzNtqrk4QFVZSV5Dv/Okr5BxZBGM
INfq0Sro1eYXlweTURme8m67rCB27EeRAd9bB5B0cWXxhFabv5ALMatBgJ1KOItz
TuQLofeQC1OMXvHo0puwcc8MYMqgRIUxWCRWLc7V0jVB9a9NuugmqeRXojTGSOAv
cEL658gzQ5Q4JpYT5LKJ7R77Zgy+2dW0NaZT/dF6f59nvNwQUDKY7npd3k9BCcTw
wv8rGLG3L22bgFketXmwEtWEN8J2WSLuNggGbEgvrVHLerObddOsrVFFOiOhXvUk
6LafPIKPmJhVH2x152gbmuoFfBtk15U8BRrAls3+PyjOsAJYZo7+7XTnUnNSdUw/
ym16buAf993uz8IsIYIOChpvR8DfoEGeU6y5QoCdKaHs7EAvs3icGYD2lhqYKxxf
Ad14tDaTsIscKLb9wxJvUTbeXrYe80qYBDOY2Offtst6xZLJlOoXzQXhR+5KIEy6
0cGk51m0DAM8sKajIKphHm/tJSgt3qrCaInBvBDVqCU=
`protect END_PROTECTED
