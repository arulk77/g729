`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aXMOwsZheStigqQcTmI/BS70ZzGR+VAZViF1kW+/Z/gu
KqdhRkyYSuzq02JU2wYnUaIIk480ogSfBm+Y833fuRHtg2LjrmXtP0/d6gtDXViM
m4YoeaXXG/lAylu+Fb22f2KAm1c4bsb1CD3BjZiU+OysALIhdHAd1Y6CbfjicQA+
rS2ejzAM+AbYRTLE+fHH+YiH+daYTk+/Gy7HzvEpG2U4io1+SRdHjPmUSlC7XP9j
jZgQy4wdYdf7Y8i+gMQBFEL6efMt5ChQ5wraa7skMjXFVFgupaIDPGkT+OwkiRQN
oUk3o1oVElu15MXp8QhZHU2qLK84I6oqTRqnuzZWXryvHyA8wb0/8H7+PukwrGql
kggPVILMa2TB6LNk7ee7+SXC9hLXKVRd0Mouk1K3nz838t6HJ9t/L1soUmxFECiZ
li8Mgnj28kfnhtwCrIBngnySoxokfdWTighCMtwyump9zX4H7J6xus+GBuWi/P1y
e/v4xQg0VjiLAKu66TOE4/zt4mnr8HAnMRFkFC5Ov/qzEDRE6ZWLFTrokgcgY/A/
kNEzG3qTR+ORAySfjzz0CWcVbWkU8snOFozHZ/7YEREHinoWiOJQXef3z8PXVwUb
9vqaW5K+Y987YvFsgUqnea4aGW0v8t6dlFIxpT/idO5lt5BwirFMb3j/ks6Ibt6X
3HaLjmacN16UXV9p+uku/v1bbetIP0X/34ONEqIFkEWN/nn8mrPTYOh3lzjfMuT5
6aG1UGw3GGebm8fvtiVgltkUWoejyfLmqc6KRVz7lipgleo2UX/mvF5gClTgYszO
/YIvbt+OqM/8cF3OB65EiYetuavVJql9x+znxCzggA//HHVz3nqcxN2uKcvhzzpI
SpNhJEGgBGGMqrWK6/xVhV1Py4NnvboWPYlcepvIDo0Vk49AgNuREfn43qv0uj6N
Vi8qKgf96mRLgcbeIFiTPILnuUDzmCe9qTcMnlyqwoHED3R/BxZzlWsO5krvkpj8
8hMNQ32VdNaqlOyYQrTeug==
`protect END_PROTECTED
