`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49nOhZTjKCfi9wwe5cruJvpEg973SgQDU8BWR8/RneRX
3xikaDN3PB16dVh1Q1jikVhF5IAAOmssFPC46OB7uIcWsTWiAhU1Ib8cdaavAA/5
ORZEozG8QTk5IQ0DvKwrZOAXwmSCc3QlQ77glUa8JHqcH6ZRf7LpPgXbVq93Y6z6
vCV90ucBR5AG/vnwypnYX4Jv6l/VPXqgF5xKrHuwCO8x73uvh/E9pxDtwxaUgZij
ZSrmKZ7jdcy4xPHNyvLTY8BwiojPwWoBLpl0RSURECCe+r2sdYvqKLHYB+V9irGI
YtW4YnQAUwECbxxbK1N/NsMpoJT3YEIrtSgNSZUsVBXnhFv2him+KsIhvOyZndyi
6K9F2fPc7dSmVXvAvaI1vpAzX+vfFBG8OOeMUYbL42i67r+Z4OeHfkHMxL2ZcdqM
IDT0y1NiuaqqS3wNUBvO+30cRi8/smoa1UZREbYNeVOYE8AeD4EmJxV+wMnW3yO4
`protect END_PROTECTED
