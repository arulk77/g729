`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGph6p055Rwfn/LdwcAMboboF1lAOKWeDilugzBUAam9
MKJTeEIxXSEeQNr7Ym/SNM4NxkcHwplWCrz2iqq02RyBJBWdf0R2Fks1grpkVQF7
2Joj0vQ4hl8mCOVCrHl3bqFUKmjc8hIf8tdH5rlZMBgKTf4wHdyB1CKjoN55IiK2
xmCDpSCb+WS0si24T91MOp63nHAXHRGyWilMcYY1d/jDjLFu6UEjOJlpOIL6tgEH
mOc/x3ssHL4rIzDgyjxxwpIuHFQHnzl9718JUtZYlF/KEJ/D7YGrOmtdt7AgjOkg
rItSlkuzX5E8nDrtGU2xGgMotmjm5HwTs+dZf/IVRtz6t/hKq5FSJxmMwvXaZEcq
2VF1WjCiJ1Fp4rwgy7xWDYPTgFOxznRApUcr2YD7G1Z9X88Ubf5xiJPebcusEGxl
pNKBHw8InqrEBWsCrlWmUp8qaB53IrRHh5+3J4cKNlKW24QUMpr2vumFBQubCcP8
RKD+ukLiTh7m2D9LqBUrQQ==
`protect END_PROTECTED
