`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xspKX+NlnkcIWhy6pA9sdBuRJm8wSUFaxZXyY5GydFN
6aetx/4cmLsBt4/5+sC7+AGzhG5oan1WHoKutQibbagLHFmKsDFWtSJi+fHhQWyH
Bq6x+VCc5sfhb7g6Z3BFkoqwL40Q45RXBSjxrRJPKj0wcvoBlD5pHmANfgAKYCxZ
gBkwkViaXQC9ZK0h6Lz6wg/+4mR3OfI4Xunp5KbVKczbWbQVPREDrymkaSzB3Ok/
vWe93JQHpk7p6+zUT19xMjdA2O3VXUq6oAMewlFQ+kg4HT/s9oko/ZaCNS1FAApA
tn55M0Hi+c3JzVxG+qna533VWLyJx5kNnTHJXlFgi9OyGiiCNx0EMINTuTLdzQCB
7pc5ycHVR5TUbNKl9XgXIg==
`protect END_PROTECTED
