`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCC82/rlWUkwbW0sujJoE4sjTij7QB7MTjDjmJ729Xkg
2W9nwszTzWSv07e9dqj2VXEZLMC8O8lSnHe1oeuUJZKSJg5MlH/Eh53YEZ6crn2C
AAJoGIRAec0aYTIvWFQyihRapIc47Fkm7NKIPPfT1b5xyEn8fYxRvKRLDnoV6rgQ
BqRRTgh8Ams1su5a4zN9rZzTh5yIbsnKmBZdCtDSJxlCKsc23wcQnUmOhzMZHDZM
PoxvBsLK0cfzhOd9B93RHldRIDacX6LIunnM4VK7VtoizC+U0QlXAjH2Q72eOqFR
maWoUFWZG9d/PrS0yqAZMUTHHBzWt1UqEmugCO0JO7AMwssPud6URsd3qWk+IBqC
`protect END_PROTECTED
