`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
n77ai9c6udZrVNg6RpvXYFhLLCsHGE0Ow4kJev5luYVGwLFCeDxooUL+hik/gCGK
vg+6R+SMqly4Np+W1CvmeharxlodiP9jPweRddpzi6nL1baufBQiq4LcHK3l1Mya
qevSUDrNoc6n9U4maMFrhCB9YD+1f3/vkgD+UDCAlIh++AFDXG5irn/brPUMC/r0
b4nrj+CCwcIP6rUOajLluz1PWAElNLVaTjpTtVuYZSPfYlc1rxIJXNH9sZVNADLb
5wQ0ucIju7zy8cqr0AA7vUNy3HUOTtORg6MXC/aXe64=
`protect END_PROTECTED
