`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40SrBvT+6EUa/xd8HozWoGe+la4ZUFY8EQhtiO38jWie
MdVzkdGnmth3wwsHQDmCWH+6LVwCdG9KivF6sZ/7sDsEBJEotFBaXqX8C417pks2
7fkjj0Kf5zsC7DYyS6siWEDaekfkR197eF/EO8daYzTJ8wiMg092VQLTYKexCVQA
WnBoIyXX9eyYQgIn70Wxub/En8NcqoQPbLY/Tg7BVk2/0b4z9vesoAfKgeivFN1m
AnqrHPeGie68gtNOdl5bQEdiFnZlLnGfI1oXlkg6IGs=
`protect END_PROTECTED
