`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePl/gXZnPR7Z6RoJNzrx87EtUDqT8mplwV2qakt1x4Hk
2L7W4k8vGTS6aQQYpTG6+gDsS5hxEK9kSz+VYpfU+0Z3nGMeaslLJfZu7jeqg2Se
tTU1fuPZ227VuCXTgw8cpMQxQJZzeO7zTAL34+txDWCQHAHIrYkPbaC19nnanent
BmhP+P2cqvTrxxe9YxZIXm25Z1BMu09JJRcmAlQ2jETG+lgchPWFN+u1hg3unN5G
uNLgh2auq5lmI4LEWxDSYICjWA60y+AC18RlSFP1taB1Hn1f2UK/7JewRgrnTP7v
KODfroN6tpubou9UTNokBh9iMepVnt0SfJhcmpLfGlWzgJBMLqJz/1IK8OmL8DSU
T6EIgJjieeGMuOCA6QzDMUNP0mlbak9IFi4iTnp36Lq4/EOKDjAFaz3M2jsfBMkQ
GT06RwycIriIHGp6mdmEnF5CKycnxXDSVVBjjFYjaUoxNDetUGKc6bS68AKy6Oee
pM+r3KVgj8HdTLavrF6FvUeQ+sxtzKqziMCT3aDHfZmm7Gbrw3frIT2c7sPkQC56
`protect END_PROTECTED
