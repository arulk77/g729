`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
O1gqIn10a4g3oWmqRZe7DaUzQusMLQ8zAdPY/iWLPpMNvsuO1uvW3HhCGxkYgsvQ
qcAckvMau62jb+DV0tXcgjLWjuBFcGAYpTaMy+whnS6Kk0JGt9+ZqPrN7ULtUqul
JBBJy8Bc4h/uKfzuTkuWH88+ZZ+Td+//JbhTS8eVjB0JrZpIg1J9WZAtJ2w+99d7
qFvN7vPbV1XTB9WuXvxa2g64cX7FVfyXnQE+5idqXO6iDkdEVNpAqcAqnurjT+ka
`protect END_PROTECTED
