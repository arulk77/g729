`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3NStK26vEPehLkUBWdWtyBSmYWWlGb/TE5hdIyL1bxyP9zM1qmNeE+DaVIma9JuJ
7ElOjv6Z8af2IkbZL/XaFaQpFZd1guwFPAI+RDPDwiaYBI1h+SMYx10OJV5e8hgs
Zn9HcCq4if9CXa52amkhAXBCKFT6F+dJ1K3/jxUfjea+HhOLafMJeiYKr+b3HFaW
EYTPvRWOB2cT2j/56bWek8c7rDzC7XYsq3STscv2/yDks3XnZkSotpHIcaNF1qf2
XnE2Wlgkor3EPcqyDNv12t+7rXig1K1ZGKMHyzptLitVw0gyzxF9rsslu1sRK1+W
h/QLIZVPwh/X7ZVO/vA9dCeODq9NjeWWyVL/ti4/Bm6vPFt+EzLXZbvXA4xdUNEp
9C06+5IVCSnamPDh2VXCziK3ggJmaHzPNVuk977mslZPvTjnPBmob4ODlBaEerXV
EHl22g58xh5SERwC01WaktiZ/77E5hY8MPJrBRZadj4yP9hlcFASilc7MAbAjjt/
FYjJv/vcLVBcsM3Hqjj1hlw5KjKsj/2gGdgFXzy4L5eYMiRtOjGl5qipzYFnrLgc
7R7cDBe+S2tU3EFiLDv9qi0o8+dqDBHq3av1CK+vAwuhQnS9MN6m0DTu5QMPDr9f
`protect END_PROTECTED
