`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHl99oNqLGR/ykUtTx+NhPRagWzeUaP/C1oHv9PUgZFC
pgkmROocS9G6N4eovidqhgRHog+4GqGASr2yJK2xXBi8Jn/oSh9Odpv+SJjO4kdu
h7l+kk9FECCqBNcPYAuQ/UQ50SKdEOlfaL/hmR09nxQURQ5llAtbBDpaZ14f3aZy
aP/wNYRRIbfYBw8bAguAbQ==
`protect END_PROTECTED
