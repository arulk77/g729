`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI9hK9Le0j2E89gC+q9TSGgXc755CrFsCfmh0RMA/+IU
aDJk4K1oP3qOhFfw+7c9ninJ937099HL9WxRKh+uIJuNUyLdp2QXQ6gi57W28n1b
RJNB1qLteGjnpaul35kBi11c10Qvp0v3d/DftjdvsVXOzFjJmHtqrBfh9ig9BDQQ
IGBPRIQfihacsiRRMreG2uIaL+Xry13CAvI2T7zm7/rcvNUk8m+UG/+g0fuJ+8oJ
fj8ddbNXMaKbQv2wQEEUSDfTgkhR9LzCrQGhjcxFbWxiLzUlzqh+5ywbpKxy1TgY
12vEAq8dLLpBXYIkCqQuh58NWZEHTeipuM4yX3knVCtUH9+tFQLU6JstZpNmype0
chKI2/y35fzWzaME9UQqQ0hnepCAbBVsYteb79cHiAbbatxJher7biq2btMpB72l
9bhNcEAZfjTb1qJW80f9sWbyiy2DoJ34j+nq6O5D/AZkt4UdCeDAH5ka6LXZu/Rh
rbB523f3qJApIFFIUIQ273M03mCL9d09+79gbIAQ91Dh6ebTZrFp+MFSgaORBKZ7
L6oQXO265UEWsYnA+MxRGAWR5rgAaqn5Y6N3ZRb5nuQqNWBj3YutDevKAMjtk/0g
vHwNU92GpI++mE5RA0KSjnMj02z675DhLOidviCy32F1VAGd0JEf5uklcDtdQLSp
`protect END_PROTECTED
