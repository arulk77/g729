`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
o1LvEcHTTqXWu/IIzT7EH0knuKg33kOPfyQ9WNGue3TZZn10fHKNM9E1AfVMeebS
LABygUkqon7QebnWw4v+N4FP6lPkN8NIMb4OAMznySM5pHn6viTx1MjxwHS4xItP
cZjbUtwrmHIjlWUkLzNH+O3EAXzdj1SUC6sLAUwOqngNPIr9z0j/T5sxoABhAjSh
VJnqDm/xPBGGnssM1Y9oXe3SMS6VDyQzRhsYPLUB4zblO/B9w3jRPnWLxOkaS7fV
YGgeCYxVfH0tD5YSWGPrkOYVgaap/XZjaGNbSkYrm4s=
`protect END_PROTECTED
