`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHFPPW94Rg4iluWrnitH5MorsG0Qclh+WH6NnHZCSuPv
90Xvg6EfrMHQaqQXuRpiOpsWDZ9oFGDclcQR7iTH5DeEfKpdaD5oLL0iEZU509+L
8bR26znY7Gvp6S4PYzjRTzlRiG2TuebacdGhlSOoNELYV/2vFYCDXakUoR44jRZ6
ad8IQP8nuYgp5T9VzrydwQ4XYFQS1yvHzxnBPJkamIvwg67ZiOlqnrkDAlIo6GGh
4W3uR/JjLu0vzh/avUMeriCJDkn3VVcb4EZUo/eVeubLLBb/rW7ktwJIWa+GuZ5+
fumvKnUBfZntZnCWAq7w5bqvj8puxDQcHklaDtcp0BXRxZkOSptxqNX1F3RzPR6V
W9FFNLYPHmldk9ZMBDnOz97IqKkJaRovYELvBLG/9agh9msCnURFp96Hicf8pPja
zFbAdeOr7az7nKq7rsHyQ7MrAgxP3JD0ktQg+c8H3mZSAEn36ZctbxkJ5bZiABjW
3oGA0ULyy5zEKtTW86Vg//++X6VybnDDLq6euUy45KRmOg1LIVRmmvytTj/sRu3A
`protect END_PROTECTED
