`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAWxaiI+8/vNI4E2+UgLnQ7H9yS5GsXIUfm2YDmM9MTz1
M6BE21xhaNqJkUeSMIel7lam8l0c/VuAX4jtNZ+4Tq0e1hLoz4oZzd3ldDCK9ZeK
d1NUIl4zRAtaDJ4/HTEiULPmfVgZnRmiN+ZvDw0uBdfNHD+N0C2H8+rHPfC4JJMO
QoaROHFVMWDDuqm1jSOzhV1oNvrFlpr+ypUEH6sfW4a888exgMvEpRyaxR0Apb0l
6G1as0wT3WRdixNEz9GMGySwxhmCIhU64lTlCXIf21oKFv1SP4YdnpzLOmHJp5iU
RV1aVJQYR/ZApHl57GzGMZ91sWs6sqzrdmSqJ25k/As7lyTkM721cvqL08Jrg9Wr
QmZZM6T4c7ABdlyRIy79y3B8opEWJBaVQnEsS0jX7YVTGLtl9HMfX2Toys/X1v6o
JUToTqCf8XdVjbglEodMPeVLJWcVgHmQQHdxT1mjSMMBDa4ikgKed0AnHAhPbHSN
b3DhBlSfjWNJohvPvhgU/JSWmQlVrISSx+8CRHo+C1Vi0cEUuaw+9eNLl1oB7fM/
iZaRw6XlLaKWXXdYW8YFCp0oyGpI1QXfHIRiJZa5G2hLahOcvil5Sm6Z/HSfsYE9
fXr9MqlyWmfi1PftqCo5JC4efTHnQcskUdf83nlE1kEO1STjs+ST+bwFzvL2ButK
hRR2GHHlYcrUcbztdD7Bk98Zb52QyTZTxYLr2QubKkteZwoTwvK6p4z/ipAzdj7Y
l6q/w5V9Dt9hFUOiYZQwVA==
`protect END_PROTECTED
