`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDNcCrkr5oQMG7GCpVZFk4xG7oCBrvSqvIVPKCcG4J6A
XkOSC8rGgPIHCBe1itf9fXKFRc/3eAe7hYv5lB0ITZ3pBVhf4MviAwy4N3DqSJIG
BEuoau3uSSWekc8AulgesFyGzlMoVpIgBXzeSLWVsot0q+26sR9ZU/OvLj8VSkH3
wEHaY8h8bpRHRYmKIG9q56dqE6phRLqSF1el+Tye39yQdhgQ9PxoBmXFe51YYpwq
BzkFNB4bimSrDs3eaSgC7MZ4QD5ytdoGYKd5EfG2jzeIZdAcV6lhkLVjjO/rBrvZ
s/rvre9QJxXtlNCqjLHFDdBS18efKxFFF9lTPlqbTKoYYNqBaspqkftgpjhqUFEE
tAIuTdW5m19ZKzmB9t7e2EQ+/2+KPeoiBxo+OxoR+I+IC85NKRoFZ/FU1j6/8n5w
UCYccBy3LHHMs3Dj0ELnkw==
`protect END_PROTECTED
