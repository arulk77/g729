`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C9K8DfkjZIPUL1E8Vi/f/kGLKD+KRwCiuYjHpxdQIQuo
Qfcs0qvBv2qC2U1OzaC7W+Wl9fvXQRm4JgwiGcntb7CR15wXm2sJlHviQA1KS5gw
+a+IExtrXZi0sIdS5lpFqw4jetbxQkKmVVAdndfjQz2IqzYotjHvs9amaU3mUYWw
zg/Hv5MdpD1DzJTblM3HypyzYd4Yaxv5LDx+aMgbf/BAnbflzHUfLCjJhtVRUaGW
ncOvj3oWCbTJUP8WQrb+Sd44oUQvW+x/1p8i9wrS4fYNPKnqE1ieS8aPJ3sVYxeI
/tOgiAG6EUYJfORDB3CZROfhzE52BxWXWpCBq6NuNGkfqRwj4JT4ssty1RuU5n/x
HidYVRpl3wsoiDFlYfBboR/HOtfioe5zJ9r2W0zA+iDZX1xD4UW9k1P21Y8CFnmX
honexn6ZOedTBs4qj269/nIk7tkP4s2vHDtj8wY+5zRI+I3OoSAolUGsushRNDJ8
yLopbTYpw/RcfCkV5Rn3egbqS+dk6JcdkWGzc8kLP5YQfbwMp4xm0H7Ghr53JxUj
gNyY6Kl6hXMR+bj+9LC1GcZ8aZ2tLrNN9Sj0Jo8bS4pfmRVuxxn0TfnDJ+I96DL9
9uTXSif9MJT4ecW3Yb/oQRsZmuBB79buUEIkyEtPSP7EdgEoAWKntXJ8tkP19OhN
m9MjjhVv0uk+PiXrkr5zYG8ncSJbUCDuPP1JFYpxXQ66Ai1lk/r69Z1rUGpZdJzu
gq4ifMutyr7lOy2Y9AHseAZYSFwRuEkya5bLMODAgtFXmhFuTL9BIEqFtEUwARrK
9n+BkdZ7umVzdjrcfRVRH+Lfqz/PILacSTuoCXJGl9aV5nJIzgDA/YcwbsyhDclg
hRdncwBowIKZCNT3xRv/YvwAGlVHQOU6xici+dPIJlvm3+ukVNHeB+CBb/6UnsiJ
OpxDQzXk6v4JG/42ucbyhmNRSHiaRrwsfSdVx84mxhYhx6v53VKwWiPrTDqYvVhi
jCuTneCTaz8XtXNyDsaJXdjT7fPDIvIhQ2UWOgELZulcf4gKEE+hedGdGQ3qOU8X
UWCCexknz3dJ5rD7vQ41uA8HGX3SSdyXbBlR5cFIj+f8dlHWbpMUeScYkP7obBaT
N1MvspGTVmnLl+5EFGkuedmxd3mXYPLoQpdG0fKvPrV4uXq/BIrVPVRjsGejTmig
AUTfPu0Uf2uaPZgwznKSmkIaOEDTJym96o7nTEb0eyoRXpltExnEfhHCrcYKJEJx
ojxrEisRtT/6kvkArKjhj49YiZ2N5P6TEXm/KjJpXrRZxW8tW4WeHVkpUsqACdEw
vfUeZ7fNd5hkwf7wsDHIVkoUUsNEDQGZBagCsOi0bhWn9dB/K9WDbi1/G05V4Nrk
028LrXxNSitNNtvX56jmizM+hBK5xQ6UsplA7locI88rVBA/quk+kMp7oOm8QrM8
WK1UZSYOU788NWRr383isf4SI9sPjF001SPcARvng3+Oy4xIGwKsIbfbKKIgKTrf
0XzjSyK0GGIpebzLiJo13EnUM6e64CgHRqK7E+UOwlvPl8lehWMkHy5sKwJr5Fiz
tuESWA79XSik8Cmmrn6H3TffjDaGks1kyd8R03qWo1T6n7SNp0em+SHlxWd73sBA
600gbLNNHawXoArz0whtoiGMNWnATNrhIut7ENLjIxY76nntrIqnU1slhdLE43Ne
5qkhn16n9vff7DWhMgusJ/F2WhF1uKtJXH/CKOYwcp2s2MieeCIhjzKO1n9bIHLj
nEYg0Yz+NxN7GMBG2LpBzlZxo+a2gvY68HG+y42NXQZlcDBdc2wDG1OGk8F3isyB
BNIDIbJ3tWm6J81SmScBkjfnG7NoudKVh5uf+7EqeTwM4k/vQqOtscA8m3SUI08K
2obMCMdJNlZUY3P8F5ZAxkQWimRiM3PGpHgfgNSO+YxRj0WlyI9EoQmpCMxAL/h4
N1DhvxmAqsi2LXxwy7wTx7q6mZ+tuGPLqsg5rjnBgF7C8RKHp+RJINqPg7hLx5I7
Ty8eSssri33gJqujvO3JOYTf0hZWDO8kRvOlzna/MID9UglN3mwiBln6xNi18S6k
ceVPzPWTfi0NJOl94+DhcVDO4OdqdonETwnhEYNNJ/RoWfU7kS8A3fGCr2Aw/qpC
f8WTuG0qnb0GXBCAjfWtGKasMJtuQkXJALTpPBo6DxHMDfsF6/W2XlUAa737TgLP
3E9+pLsf9nTmU9/c8asT3DuZafdj01GmdkFUd0pWtCCS/mynvhOcHVn0uRRqIf4G
e43QfR3GcxUHKs0MHiXzb1G0ZKyKvINXOkEqlr3KIqnL7RKgsBBmdE9HI7j9vJ1o
ToT2r71mvySXaguWiFOa0RW2Pm4wKicjbCbHV6/dczEV7+HDWvRJTRnV6FVOQl0k
sn1o1ORS7vgwiC2Iw9SsAcvl5UAHS7GseqcAeePLczqlFVMPblaDY2lalxCAKxdM
mdXTRtnfGR08WzVUgF54zIEfmizf39IY+ue7P6CpgrcKnsSLSOTSwY1wp+uX3Wqe
ckfzjH+c9hogd1olfak1kpInGSAU1q1iK0XZofc5r3rzxYKMTzO6UI6juy4wtfyv
/yWXTQqtTmv1WlM79HlEWvZs8J5Dir7qLOcD3aCb/sXtD+pu0nYZUL8cwbyi9ZBv
t1Tvt/F8sIqNLFSd91BfxzK4naqz17zE5ZtLtHylLPhnNYakwFa6ygXz07lxrlfk
9rzjKJ7cPf+/4N8q0Tx1BNDJB9VFKzOwJOOCEpHgHDxx7X0/PkdNQcNdUiUh2eKp
06SIzc6V0o/LR7iMBVFWn/snRgKMctgVNLDg4WXx0UCZ9p7W0Mk9AMVYiP7RPdAQ
DepWLqalcm/EtSB0MdH08FiKlkwpYusXzOOxiMv31uSJuSnoZLd98ARhDD2RiNyy
8ENSFrKPjOF5sNgZ1Lnnv/dljf4kZKF13FG87ga5k5z35tKUCkqsVvvID7Ud/j+z
6ZScD85tH/+yt/2lVarUXzVUCKv22aAd4qyY/fEEMvMnIoHFsDcm/r//ibZtfXm1
3RsNrDZilOmswjKNHH9JvRfMFlkSALknAXzP/qydoTlEZ0b7PppVMtSRmn4QaF25
MSWSFn/eTWRaa89N2yDW/qChnCyVi8iN3C2FwEJPd2wkm4F1e1E76yL65Me+DWlD
orHvJRcn+oWMoB8JjuamVVu/DBZEB0m+lst+wxnvW+5ZMQMQV3EVDdRPkTz9lnZO
Zok6rEAYy0+1QgUr+LBCkauDiYRU1Ok5rmD4V6t8Q+ttxIJU8bZYAPyaqbYg6y8m
+VuIe4jOkYdwCKd1Qupy/3mXxh7ERi/lwy+0R+e+KlKtI9oXN6b1gfqco3f2GL/h
OJ2hQAuyoaInuRx87LI0+G6ONS2/HiXp4vo5a4kmwFSlXJVJGy+szmTIIZIOqf6P
MD6GFwQUEhw5CHkL79FhSI6hDqzBPI8zIxOfBEByXpQ=
`protect END_PROTECTED
