`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
7h/KVNwzj5r9TpExoaMnMMDhNR/92azD0WG3s5nPsz1OMLDTo1q0rQzczWRuqbGY
T0N55vl3ng/8TRnsHt8vhCoaDP85ogbudjWP9MlYJ5E6GgHETqt64uEiFYOMqcQJ
icAHRfacbNSNeZemIM0NadrHqFV2eaRCy3SgcTs9o0tK1OQTCoveM/Mxjn5d/iyH
lVaYV3BDHlXWSviy8AQ7z/nQzl2cMmx4jBVxhacJHhP5iIkG3Wnk5CBiWtaiapco
ePgJkCoZ5nUuUZpnzb00Hv4jKFpTzU9F+L8L1qnV5QTNsQlY0CsXVgWrhcBeWTI4
NWgI963t7oMfA+nB79hfma3OXWy9sL2pbBRLV0TRvzc=
`protect END_PROTECTED
