`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAYceqQxz5WT4hTUSzOf/XwFc3ZGW/YJ4QjxlXhjLkqrt
O7gV6m0U4bT4UmQP2mpXkK1TCPm+k3HClyzBbB8Qh9WZPjN0jaDwGNiML5FixnEU
m/asmmvOem0/Z0nhy5m9hJGZNWrMKhfkXk1bI8hE9UBSc7ffWkJLRzyRiPObMonu
jpuc62hwHkUY+ujGjisteNptHyQjAikj727FRmLtPsxD+hL+rjwO6cWTT47+W48j
jDmQ4ac/qQmZ4LKdR7LPcQlhlFG22C71L0vkC7UF/PJ+M6yQWlo0g+7aoxX1G2+I
GJzfrv2um8silR7w0QfJHoCTgPfM6N/L/R/NWPG9StHL5/K6q4KypkA/8IW1zet/
lf4vfEhXvfA9wfEFqJmx2iIIv3qwi8dK5qGio+Nb5YTObSoRBG3QlGY1zyKwWSeW
o0Grtjmzi0vVITu62aohNmm2QUf588N8oOogZEG0JicoQhkNrTCW5+ntXgPw9o59
2FUKx9LwRg/JYP5PmZRkwlo4apXG7UgeVdkKksOWQxgERxU7r+ZqNZDG9bD5cXME
ekC06E8U70dj4NNDYAikuQFW9eZVhqCRIl6RK3uHRf3vtwLpA6O/6Vzx+wI8h855
C4RQole4kk8VNNJssDGXw1asFAGwrSkvopHcnLyQNkFCGgSWh5Md4th14egBPW3m
sauryhP1zL1dkB6DA5ijGbXFWE9YAsxmtevX4bE41R1bCyfQ4oww5Gqbu2yuhuxg
aW/uVBkv19qrXF1gw1xF/Ya1FosP3fqehWa+kWiITSJG34hrx2GKll70ywfmYcc8
gP/RWS9kn/L404mQwIvCuHuCapqqlUBMOzESCeQNOksfbEUiUGo1R8aaS2yNauw6
i6XK11KzDb2srYMij8B+AtGlfdrihEH52pTE7kvl9hIdK2BiO2wK8e/UhkEfHc0E
8OPvUVYrlcOskyhNpnz17v7KG/Qxa+YOJBGE3wteftKZt5eyiXkueGxZUVabxgT5
bFddooyr8FHWcT/exnRa4ZG+F0LrQspRROVnpnk2u/+zV/dDyhBqQowL+FoKc0bu
CaB7dTgELqjHFJcZCQxRcqFnM7LC1S5xASwf24drlpJ1CtdMWlOh2gE06p9FuPq1
/nfrw4+6tuiMmIlkKUUsXWinYqvM2qM18b12Ai8ZMaXScxIDoTB84C6wfkWReRHJ
dvL+E7hqsQYs727hcL6f47CHeBAcg9SrRcCao3yJ/EHmEEyKkIbdZqXmAY1XuqS6
akpmCypJQsINpfzV8LjYm9Jc7MNYEruK+l+KN8QhBLSyWdcZAqJ6Usp2WZ0web8K
zuxsfytB2190V+0rBjoLtFvGbUTYQRqHdkYyn+QHeBZzkb+ulT7jK72elsxeOnjG
nBhuJdbUc5kCEm0GTwf6cdwHvhb6HAMUfQxw0x7ytD1nHRJFo8mbmnde934afoYW
7/+l1PB5fgdKIi50mTo1H/cmn1l4wSOJlco77wkVyV20LAw/wbaQ/Q0uAfDulPVg
1z9XnH1mR8MHSzkXZ3AHi0+JM9FnUgxfwY02Etj6HB2UDj7gdOIp8/xq2HifxyHX
dBc8Dvphx1EsxcZxtD66S9kDF7XrMYV5PJHhQyxwS+qvpdq3DwUgW5uMLYRD48fH
TpKiN1QS2TmfGIw0roK7yQId7Y3CY/hEGDGQDGX3LLtBPJ0292qivtwB7FfMLotJ
+i2YipE+Zf0VQt1noFCJ8w6C7Inqqi7f2fINlmcXgk0QdcFJqbFt6WB8P0pZDtqL
DOV0wO6Ih7TEjst2xcL3XAIggH6xvDNhB7JoLyNc365NZgPBbATyLIn4SBzS7tjl
JlfMS0JYApskmCGlrRo65WByj02Ma15U1HR7iu2GLPZNvnFVD1FvnadC3Szm39pi
aRpgpThZgCAua9IdqhCzaHksMoSGp74yH+ayh27PuY8qPCoUg7IyxiFr57/y8QBG
TNw7pa66A6pwxkx02bkKr7bihanyWGHjp2t6as9W2WmkU23tfX0oSqJuEwsdLuuq
qCTVd90Tt8fgKi++SvdSkuFAPjfZIG9NJZNKnTE9E8+7Zn1VQ+gcw4+o1bfYALI5
sp0vgrbFBETLbF6WkKkVZ+GA6ir8yeSWVcFYWZWXOUq0YAGoLChIP1GveRpOVhB0
2vM6JuTQrtHfLLwSmLokKNwGYBYnCYeq/u834Roq6SkAKl48KcLdYJl+KY/RZXsD
MwV7am9GTHmE2VROrdCtLDzIVGFjNqLIHDZET+7HtYShH49+JQKWRyIDs6a2Xaad
sZOrW+Jh3PbTTsYV7X7l+AEYJ2xElOP2jSsXMhS/ufayDt6kl56sb5HWl7y5ECkm
oRi7o6yaDOl9l323hsEW29R0iJZuHsOKEM1YK4CYe1Vp5fhWg5sk+lStHwSKGHUh
UMrL1wOq72KiaEZfk9dwa0winWkpgB4vhGm9UPHEoQp+HIHEwIjobMeJPQK8geOJ
AOH2gxj0rTxpJFvG6xElMbeBKIIz3ASzqPOMfGYNJkMfAiQEPLQsknIsWXc0k1T+
NBBfwQaEyJ8LAzSrKAejmGegqw5SMGovngIhuhGA0D65DwZMcVj/4g71a76WxD1w
NHfW8qFAAtVFVdbxQ4n1gmEG4vVfntrjEw81Utzx0JnPi+Za66uMbk6HQvZti2NN
ST2wBwQA/GPJv56UbFy7fG4gHcYlBa3IRfcS+hL4O/4ojgjVcnAyQi291NZWCWp6
BP2i5L/6cDac2+dT6jrgspQY/WLuRxXoZQVFzTRr7XP1y4E6Wx9FdPfJtH2ML8L0
lzIfJCFbirVJovhKnW/8FyIEQbMbPP22/JgdlowoZFQJWFJkJgzdoi2wan5iZt1e
x5WbCZYze/a17GBMbkhPUIsBim0SE6ssAaOplrZAh/xoQ+mLpCMDr3o1+w10JddZ
nnrm8jNF4yKKGzgMqzrwUGE5zCOYDehuxuR1ValU81F7P53RWNRUaffy7evX8I9E
+Uk+T8F/5XWjoEdER0WxC9nRR8RYQDzJoUDr8TRDaivAM4fyXdWwMmP4KI74PbDJ
G7YDAyOjYpk4tyzqlpnHce7GU6EP/kpYb0n/RCxTatr2yh2E7k1JvnCejHkL4M/P
0BNCc/JG/V/ZqlWhuLOI0DSu0AEAGp8lMtalXhUSPhjOgS6uxG5DeTnkHFBNha6S
Mfx8m3HdtWS+Zc7H494El5DdoG8otpdo5rYOhhg2ZZaPOs4WL1ym78XoXBb31gvg
`protect END_PROTECTED
