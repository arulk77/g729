`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
62G0NV65ZmCHkB8DVWXUFiJmdWvYCzPQSk1bNtymFPvNDT0FaXbiTI847nay6om2
rZhvrVbNXBR3M/qpHOnx3OGn7Bv/2r1CirQURH32UN7omKIZx7WKBpyl7ZnEpiGj
4c1iJ1fdJjZkvDH/UqZFSBWMFKwssqwKEb9U1BffEP6y4S0/JQLNIkMl1L0VMQYX
2NEqj5FvXZJ+r9c+k2LxIXTgcWqbUGw1+05g8nTNi4LQtuXYZIxVl5ptGlaV+qKa
vC1r5ahii5ORIalbnkUgueTlSBwsFrdBMIJRQVcRir0=
`protect END_PROTECTED
