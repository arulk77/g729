`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IE06gK9b/8WreQmxwg00ZDcDP1m58n2DeQSR+ADhtMOoXA1OjKvZld4GoLgL8SVQ
cLS8Ms/x8eQZRXP9nhp3TwKjwEMK6bc8d6hpGwV0KoEru1+hqyakKQHXdtGdQ8J7
/14jR00RhdrUlhp3F86G1wlGXer1eXRDXZflcS+5VQ/RFeUcBHWrgIOtG3xuyzIf
u3pjfdeeMZcVgUcawt8BM3gleFR7/f6/UDnvuRiheAfw0ToK6dpF80TJogjPNjVy
8YZmH3emo7VMB6Q06oF7HsdedOhTlucdttc04H3gekty1KzazgjNhrDUXlHyGlq6
Mj/xNMSWOM5w6z2cDgHvLJTwbN2VTNHq95YReZ+Ih3YXcOc/SM7beMWV6w+zVVET
aCMyZjUei3V7nJPnB6ibLt+cjvptcEC/fHrWcpqdMq3F7lqBJsjSWeld+ELMYbX1
hIDVNd1sR1vuwCGTFs7bPw==
`protect END_PROTECTED
