`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFokW9hVofVlxrNiPbVhxadv/X1UD4HX3jmojAre/Chi
o134NgncaZv8MTIluHkFWA9MV1SCbSrqX9nzeJLrGFzLSCFwzOBNTo7y7bhEmhVG
rQAnVt3//d3Jo6r+aQ8WqbFf66nJojeMWBU16rKq7utCz6d3v0cKa4NpQLn2pfqe
BEKMjr3bxoCbq9tWtMfGhWbjaVnwVbfcucmLnNRAtjVE5XjNfbJ0tdsjsG7KXYiA
947LaveOWmUSxqVoxv2/hmOC8ZuwTxidCjRmj4Iat6CDUdbR5lOB21ChgaNYXfXZ
mt4Hau84TjEk8j8x9RJOxZVYRHRPm2ClzhD2f3WWIB2B9pcYWjlC54fG6y3O4ACP
`protect END_PROTECTED
