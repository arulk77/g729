`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C0sKWXTqxiOmAewiNnGZ1zrENzI9jYUuXV5mVdvfSBjf
rnUEL2f436jNj10NlA2tUh/HVDoCGaQMYAKTRmPl15opA3MzHxLt7QZUQuxqXCFR
CoOCcpNFJ0lsamfKQAMZlxbCt+0pMGZ8HuJGQF5ci3OlxBmfus/2GWMWLUBY9aCl
jU4gqxqVtIccNi0LhgydyummfAt5YT8C17+vSDx3QBMEg9gwL4j2igGKt5vgy5P8
PNsG4hMt9Hi7Gib6OYOcT9gceHzD57A6ZqcSGGkYxQTrA/3CcYzoUJdQhfTY94xl
OV45Tq40cTeFYdD8RFneQU2D20B0ks/L7v/+MyfSMwI0Kaf78InqI92fYXgGR6ew
6wJ4kMAB9k/gqw93/QHPCZzNLjKpCsXe30gWVxayV5i88s0JOL8RaKUFaiDb94q8
sJ0j7LX60eQEIqNR4XXyL9DqcVCUV1hsVexElf3/tkOfg8Smp7h09XN3N1H4Jr7Y
xtGtwhDOQyazvP8e8y3AXz+ZnNtCKHIjDvpBhM5BXnGyHdvlDPUFHiiEBWnTMgzd
n+GAUP4XtvlN1WhaOQ9fwwiiokWuhkdfErnC2U1iOdzTMjW7tPN7D5JUsFcrya7y
FzlOnZWjJJpRNxOSVzOogVq3eHHR+rAT041mLoohOAp+4wI/8uk0ciN9CyPsE+x+
bYyzUTlMdgLMqxX0LGInzkW5vGrlZx/tlcerbou67Ha0ixUKajZKkn3NMElXizYm
TNQWSjBIBdbRdRsLpqB76peXIr6OhqbjZpe6ID9KuSZuljyXI8RVC6V26wnYaCuk
iZx4kbcRiJrnQ8SuzDzD9j4/o3WalfnQ3JduidfWyv6R688Za1upUnjlTfaXQ0q4
V22BO0IrifvzVe6TjHjLWRHihrQCqlz6Z4z8o4LmqoqHXABNdUE6YlbEG7GaXUTK
h8sriP/tjUa50f8IE73q7xcVNzRKMbUPVnWvWZKaNYAhDDWs163reU1MkoIiMThJ
M7jaU9DJO6KEYXw1qm6TGHEtkmJBkwuFpZ/tO16H0Q6yE5PE9UP5/Wrx2yEd+7Pk
FTppqCNltvGCE+kPt9Cr6V+iiAyljg7KfaB8Gx1sZLHes4MbMCJG2Gu7fFowBvXT
hhwQo/6tkvpA4Gj9dcLq69mO4u/8sqsCozBXKrBGfa9I6I0GLhapFwvQ5dnEYrXg
75o9kRk9MpATTTeDwPGo6zg9+xIA64uPkGGtnyHE7wY=
`protect END_PROTECTED
