`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL83TFqqM5JZf1WEt2arccWJd9UImitxThJ0YmsY8ZXn3C
6FqOhOy/f1BI6xzhl3TvkPU4S68ER70Dq2IDH8l+2pfY685bYZh04VBlsvZziqM9
VZD6ah8sT3SuoL7qSgCIrEJSmWebXeRbR7WwQ2Ga0Md6gcZ51PnPhUhrZW51ZpbH
0+wbAqO3MwY61LeLgzDyt1qs2ZU1UWnRPiLEpoVgtAcMZDDm+roveSqBdguMBMQk
V/I7mi0DnJwHj0xYisbGT+2pJFKWiu0JQG10CsMRHY2Dho1qZcLMtr9yBdke8oL2
M0lyUs1AEjzPzaNSKfHYRsnmNPv9mxR1KAsMCAjPnsslJF6pnoQeNwmF8EYOnZwc
teij41UpMXPBhiKi/p4t+aBONcV+nXLMc/Ewsz0DRq0l+YoBV7YBTfWrXYFPc/Sl
6lsGoWinh0nO+MxRtNLnrTPL5hMbnFfBRMGiayyA3XgQaXd2zKcsrDwSKhkmi1Bo
PWa3sJajKx1WL4nP5X8veR4vSrVpIrS7JBsg+SHQlWqPQwjmW22ypu0OMV11/cZ6
N0U4rHt+a/HWPqmaY3V9CPefHSCGX1/8KPJZ3L2WpWVGD6qVl3FGO8FH6ESDjDFC
b+GLMv17gAbh4H00lNP1wAFvtbbMimFOMqky2ChAM7oGKoG25GzLMRyLD5cwGVNr
TC3k/Y9Z0swJZtCRMvEYd8K2IPWrbhLDJzRriVGNCdFLf0DeFHY6NW9HzLylROcb
9upIREiRUx4mA/IWjxeghROy7oIS0iAcrmjL2y0vKE1i9nskbtsXaxjoF0atRZiM
GI1wdFbFqTs0Sx/C2FeRzU9i8zikpBNFEiOuY/rqB9/3AfApIuR6B3aP6LIu7gfG
le5EpZ9EkkYlT9t3OKsDe5q8XUyoWPzdvl5cACK1txmiaYe4KQR/u1p8U/+vsdrf
6uRWK7dc9JZ8yr/R5S406dqUj21Z+dmu5h0evnKL8E0ABEhSm5yEGHxF//W3/+/9
Ay77pByo1/A2zLQg48lJRf0tf2h7elP4R7zE/hEmQLLv/3SB21gDfv48vbcPRz5w
QJDwQnCnoRUkx7nGbZN9+/y7tNlfWbJVMWaRYdTpW3ghaHcVXGYuFbutBtUsQ3Vr
aGqLIwsqATZIi2uoAdiOQNbQKX3fS9FOn8+E1dOYeKLmZO3ZlGZrUIC3EmC69QdJ
os4dAfJ01AW/HkniBb0gBxj7Cmlekfk7EHORTTt4pxixNeJPfNIigualCX/s7Kjk
mJD7lCpnSLVjnTIneJKi2u/kYi7LL1Ai4fQuO2IB4caZh2X6/mRuxXr1yxYhEeNs
lNsYXS+enMIpQF2a1tghREMd6kRhv/qEgi2lK3tt/Yg=
`protect END_PROTECTED
