`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1afJoxWfeiOxlXNMk/DalSmYzsp6UzsQTIbKN/U6Z9lJ8
1sV9y5fyu5s9VtdluQ++MtxVB28ymYzf7zY7YOCEUlhCDIGXN37UE+8L5DfqpCOf
MLKh8KI3m/gVguc0ubffgVrAH6UOxGfnw84/4EYhSGZONkje2KCc7bZjmJrIlg4T
ENDqwUTScW1fiCbF/7YjWN0QZYbRsHjZg6bA0oJ1BCu8G1pzC8M5/qHgfhrD4bJL
N9YnxJ+qVMiruGUYj5QI5b5ko/dpymJkHRgm2oOJ5y1ukrZab7ZtS6Kl07+1VeJ4
`protect END_PROTECTED
