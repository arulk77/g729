`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu492Sd7plX/v1G78nQXsFFIWZ1Ph67ZIgd4d3E4dW2JiI
GY8y2IU4hJQESB/SHzHRifkqAcL1w3y4+UTsNKfgeI9BBcacGGzs/6CX3zhgoFIV
SXCf+iPODLWidi2mxU8tn9Q5QFto6gIE35wIxQXADCQ70cy3RC+V1DnaDwwWR/mo
Qr9sAy6/U8UjC5AQztAgTt0By/kSROOciRrkyBn7uPh2LkBbNfRtnSuXPSncUDp+
MhwHZzz+xdoPdfWGIId6lWSE2h0uqidUoA8Z6m8swuE=
`protect END_PROTECTED
