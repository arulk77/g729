`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aTf1RbK6AzUC2OSVAR2POftiRAPHbv7yXWmrsZsMHLw9
oP4J1LLphFRSMudWrlxkwM+n5sHD7FI3f00vui6KeRe3uGl8zz0U9hjRO6EKRXuK
Z2WL/Dgdvnh9BecNa6Z9jONE5yX7NyIqz5QInnUvbY/jd9LYME7YplywwkDROU1D
j8N0Es55476HnHS9+yXS9Riv6XPs8R3eXmD/UQ6CLLaW2iE/OKW6ZOmc/V3HbTXO
ZYlJPr2E3x/eCs3c1CZczZAWLSw6Fu8tXPrjKOOSXWpuXjumyiFBniQrnguw8UD8
m0ivsAzzWXlP4NJYuPVCADzfqXFvKgLEz9Vf2tfkpmC/hP1n68s8nNIxyYM46XVj
8pey7vbhdSod5Gvcqfo0Qe5ohhVFqEdI/+ONjPM9CoIUinr0KtWemYtZD/3qhMQb
j21CriEJYxykR1IDLmU+18XK3I1RIG6bx973Ij7iolywYNAFLVv6/tmmUwM4ju/r
IXSsYZ/n2GVMHBj7zzvGMoS4yf5uj9l8gIWN2OpjJE0xUygCBfrK0r7wpxspBasD
A/XAXrgdGU4bmjMssUQ1RSnCtjmRRyP3zLelugUwSvUEjuLLLwvJ/Mx0SOV2TiHx
kaIDmEp96JEDnrXFphj2N8+mHFqvg3CRu+u2H92vD/P7qq/OFcwVX+mmnZeLSpjv
jTaKcrbASqq6cLfCBArzJHyGNRXni6MP5b6ySmQ9KDocrLDPPz2uGjZWwTBDIhHm
Ceyo35eRx8OMePLJaApqUNrKMvKVvXrCGRs07GcCOq+ZwxikfHCnJ0K9sAAKuxqe
WDYgmof1w43ub7suMspdPxf67nqjMA+CdM3vDoK3/DA=
`protect END_PROTECTED
