`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLL50bWk4gKmJOWQTil7z5cE+aaLKhqseUWkOvmp2j3w
y7HMMOJxi71Wq/XH5YbfcxS/RBdr5oMmG/rAo4Hh0znNAyr/UnJCHKueRv4RiZoA
EtgQQVYdjY1hm6QUz22HDZpZ2ifgo2u7xTwceGltHV2dlXTE+TtEko8aSEd1oys3
76y5SYWMiHYTpozfj+Y7TRtN87MVFrkRnbW9D1Ab9kiYgXGj7H3o5XxuSfhc9guu
cseYeshEl4oE9mNLJNQkxx04ukap5nqEb0I1/js5eKHyP90VIsOPNFE7F5oTLBYZ
d6xTUQEZ4MfB+gxKac3/Ui2/wwb5lAbLVMJz8/5aqZtz0PuNiBAsrRSKzXR7AS2J
MC/FoTUdXjSZZFU1mUmh87MoG+1Z6B+rlQ/iFS7kqmRjcRVEcs4fPgHsHg9Ub9Yd
u+MhpqzjT4SwRPby8o6FupfwOozphb8NuCjbjpCp2cIv4FPqrSTxTD+UL+g0PKHh
Rbzz+QKsFKUC8d64u5Mg6EBJN00jt6xtwyFKW+JQra134FI9L82TjcxJxRkYbZro
`protect END_PROTECTED
