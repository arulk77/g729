`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePeyGJoW2FoqV14yhnbj+mQfbskQLYzRW7FcGrf0hh2k
yomkDMr7bmKosAb4VQOF2BQa+LZMHON+FDLaJKAGNqxJQx4B4OnpNAab7S6rJhr5
2hSHme2js5eUhuNrRsgTDNhuVfbyaWtGoWE/ED8JgHqT36VjHq1GayKcJsEesEIE
M7J4/xA/V6oa/PJvUUD5zA==
`protect END_PROTECTED
