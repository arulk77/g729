`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM1nC45mio6Ixv21CfdK+Q7jz4gxRNlb19MYjOWUxWr6
Oobn0fJDvblSFdDlKV9GndXMMmZMLcfpOQVoArL5Fr8xW0fqa/l48oLn7MhSRzHF
4OXP0FaKEVyhaARgCwI6u/Z1bz+9HkcShsxdDvBfTzhTCAnDkWqb4NdrHlaPxRjg
IBEMqM3Dg5+iWdg/+4l2E4243eYIiAAwArTQ6IVXkj5nLOIzoiOL1xYsU+58Vdbg
`protect END_PROTECTED
