`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD1uzgAXUxKkx+5VK2KVheqRG7KgP/RgueflmRgJ40Qa
OSdlK4yxdbAqIxnLu63tpEn8SLN25AFVyraygO11eKoMN9fXHsoiFrb2+2UGCZjl
hCi4nAeZoMi58g+/oo8tuBsdKaw15BOIyJOGmRDhWWQqiyuXhavQYdmGCxJNALtZ
xNm6cOsS3em64qHP3xydVIeOUtfXrq+zroe/GaOA5jk9KDQHjg1yY1X6x3eOquPW
8U+N6HZAH8P4Toa3AkKPFlaZUfqV706GxbypNdH7w5KM7Gb5SDv7Rx0wItYoUMoH
I6w5P10Ny27HrwNaGZBydoXRPL7ArvqEN89lNesSSuI50yYx0yj19sdL2hS6WNzv
lBJDLVPJm29uFyarwivnXVEua8Bzezxc0icOgKtH+WKpuBm6ajjCT0YBtaD6rsir
JXoej3pbayxH9wGZUsdz28nZCnGjbOTZsG/lxehYFYv5Gtlk94g5nc40GX6/U7w4
/Hh3fTJuIqNc8Od/HrdwHghANur+gEoEERiSzbldOnSIs3YO6i5Qtyz2/J+eag4t
wngM3znWNcI/TdEmLuex0Zwqzbrhg4aHHrJqr5CRvvNbpuWF2YXM9vjb7ylZUAU7
0b27pSKTvNKBCOUY1ptbybbjUl8EJ3UY8WQLLWv4u5EkGpI7M/021Ex0wml9/iLu
`protect END_PROTECTED
