`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
e8HmnbwR+dxiXeZDDc5BVAgrTWPZ7NhPjZ/TJyFF5IjxdcO1Tsp92qi/eadTGoIJ
m77wfj0IwqFuoQiCegz/ebhdFOadLFM911Hvld8w0o8u0e2e+32onty4nC40Wm23
McB9mvXIcb+yoCYLl69Bjp0LvtH850sXgrPNibXOWqiSkLwNCJFGxiddYmzyU52t
tW1QrW5IVF8NKt94QCkDiy00epjjIYMqwl/HGV68UoJSIc1Q0TlV6TmBIjVwI/Ny
eE3FBwa7luW7Hett30BipSlRaWP6BzBJjrg4Z9NvPPj8jt4uGbwu+tasTI0Uavb3
wZdlW0Y9I2LByqqyq9rxsehB/obTinCBHKny6Xtupcg=
`protect END_PROTECTED
