`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL7OUCox6GcN/UTG8Qd5oS9OzcRk8CB6vP+hfUYklHua
1YAaFhfQ2VOEZ8d62QIw2f8y/aH679Xg8+W7rLyGNw988hngTPEtgxo61Vht+uWH
U6DdYdcoPgnrr++GGMvhP+s7ALnuz1ak+wW2rsrRhjVLD7bKYjYl1e9tXj+JoTxP
Lqe7W6FJG0uBc8wSDUPR2p5qYjtVCLUSqiCf2YgB7/N7dcRkOn6jm1soEk3bFGVr
DfXStq2Zo3/nRlPPYqRfEkagK7+lNKcZzZlMexcv1DM7K1cmlTIU1FyXVqYqa0Ow
PTQEuFVubP/L4nwuQtOzJ/yyK1bE1u3jSxtDgU3k141bK3Z0f6lltJMnM/LTw1dj
nVWL7SaNxUrvlB6vd6rgog==
`protect END_PROTECTED
