`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
oN0Fynnnb1iLfl61QfX/X27AIX3zQ6kRGFSOcS3WZYzDkRj1LKVqObxZJiAGlnrY
Me2tEBVPcmwsrJq4xXoh96aCzyHzrRPoMPFWu3W/NJtZBKCvKClpuPsVdsD+vxTl
h+l1z3QEEVxY0QIMceNpioH7BXYudwagNyS4QUPuR+6mfI/dJWlCQ7ybxsVxw9wT
OEB6aBWOdt6DOlVkf5FKX39i0/0RJdEXHWEryy5b1THfn68UCeJBtqflkIN/EZED
hV4gEhHIr0KFOZAlZ8lydjLtdB1suOTjPyWv7Z+zc8liLRs3MVrS6jhniHlsG1ru
V8eBxPrPGeVSdCbhIM8Mtw==
`protect END_PROTECTED
