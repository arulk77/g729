`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAt9VPSGH7K64ouxWuIUxXcxtveJHGh2a5BTP7rbyPbM
tA17pN9xvXqx0FE3c4KPiaLqG/ep5Jv7+FtWENlnxLrCOUfNZJ6QLHn9GhIvIuZy
nS8fYGtDOk3VevT1Gv/F0Mb5MDra1cRdJj4+Fzlf3C/J3CI33IjoyuxzlTGQaLQm
1xwQ2pbZO9FG700CxiU9KBdGwt6AGn37c1SQJ1mMs8jhnqfv5b4woDPLE4lfZN7f
hHCngklEW+hQN469OtgXiAJ3mEdNBKmD0D/Ecx6KEqeBQ6bkJP3Ty9h/eeir8Jn1
fSV3KiMlI9oQmqC/DuWdo0f97XY3qMr1qcAcYB3CQntFL7doDXkjivw0kNPwYOmr
nZlbU9l8s92xNInw0mH8/7+wv53B7LaQlz6GhXcBsEIzyTkUulbWQFxh7MDGIVZO
8V4psbqp86q02+Ot+6b4mP7r+w+465lNf7zG7wcBepwB1a1lDhuc0zG76epC5DjG
/i+YLhrtw/atVBgd3/0qM3Ft9Yqb/B7DqHLjeNkpTqXUoDdH+WV2RYu+I47QZXaB
CskN95APT8vWY255nH/UmLSsonALzbOtVr1kb4BgVPYw0Ek8moyWKJCJtH0S/Q/q
Z+WipfoWqu2jzOw9MlY8d/r1e4KL/f5YjmPD08tmCZnJ55hcKK44hnIsa6CR0mn5
SVP/glw6kbd+M0693qxlECWBukJh05j0HcSOYhn5tiT1zZeSBNKTLdeAPgPRKq01
fU7mXd5piEsUdkK6YUCKe9etva3ouQbiH/2BhL97bDzh3PD57PrWMKqWTdDbFvEG
rE7H+j/mOhS3LAuaKAW9gWtbzEIsHNhoHMDueKA5WRA=
`protect END_PROTECTED
