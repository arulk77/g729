`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46RuMQNnbnmdRYVYod5CvyUofJBM7WfJ7U6P7as0bRPe
fZ/JVlSv32q2TMlTNMLOM0GgMCtVmCVojv6lQSvUW51yoPgI2kXEwqfB2NYcUpWG
1JiLNRaFKf8m64h9AnVLja+0Icb8BFGmbvsDomssLx12TI+lgPvs5366L8d3O+0W
Rx2aEu9XFOiEezifsmtnpkdHQrxeSKXxRvoGhH9mKfW4VuZ0dN1zI5nN991cbNI9
ClEnNVYpuu25DY2SygP7GNMnig7s/+WKUGfIKpG9MyzDQXsdvKyx5IEre6+c8r83
EWvj+4NBN7+zkDhwJkRiZQ==
`protect END_PROTECTED
