`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDdykl2HcKOnTdoULDb6F1M1T4B9sTjfwbB1Y9nDVZhL
6QlbA3QGAVvt/eSdHfxGNfTYReRbqy9lig8aPMnVpm4YXRF5P55O0grLUc0V3Qr8
anrIpQ6XFgfjVs1ZFA2PFunKlLifXD3uXTH9N8dBPeYPZWLX2UKxYP3e++0pQ6ES
P4Q34GU3NRMEJk/24U3sBf6BWwgrnO4oh0jU57ZJ3sOnWfKGSO3tSsY8uLpJCf9s
jDJrsKdhQ23t/fHN8JsiaWFF0vh7kmZje3QfrD0VFdmkPnYu8CBClNKaf2slU+sA
cXWyU+6+bgf6jdXQ73amubBBkkFZ4H2i1vc56P22daiTmRMajon3JXjRuQlxq0XO
zeBbYoN2MaP3swsRDSYcuw==
`protect END_PROTECTED
