`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
FyKNwvt3XVnoLNvlyKajFMjQC57d0lycs4/it12hWMv8Fdo+Y9y27ftbaCUKnQuL
Sl5uXjFRkCWIyKoMnSH3lT390KV2Ad0/riQ8Ploh54VqQb7fajTg2WTIVwR4bpVR
cLOYXRcD9fwDTTjsdp1FjR5MdA34k1oIUP0bork2eaLqH1VTCY0LP0BbsfCP7k9Y
mCL3YmutlyxjVeT9mUs9SJ/R+Mzqvb1OfggiACp9NxumrA9YBPTaJV7YLXwNyyYd
xUa9vr24xHCLLiKaHbMTYG8lP/NnE9pFgTor5xPDcNQq1wAvOST/fCBvg0yIirx3
9DAZea4IV7U2yzrChhF09rhh4C+uBI5bzNoMfLoCUXngdEsup+0kv6Zndwtq88eo
p8Mp3NqEYb87SJAos6/1RZVKYH1cdSFIHY7A7ePbSZg7MbaPc9GNaOq5N9FDWe2e
jW7VaU6SzgqPgHKY5wRYc5vIA/JyJTkR7PaxLvFpV2GnbEODJwjDXsNZ4/mHw7SM
xo7wZ+VwTz5mBSIjLrr0gm6ZiITl/NlbKqAxXhF3zEk7zxrOAX0pK22PPvjmVkBl
BKmQpRNq/PEMXu9+2P8eYFNSxWczMkBeCkTTJ5hIYiPOsQxvf8ollDm+4HRmSl+M
w+S/sIqaAXP7sRZzzo6qrJHaRveIjCwBjDllAhN7HybxtIIgUXmPHautmj4Guw+n
keIbuWCd1d6YyDPg9nWbX78tJh8EPcPRWwvcjgyUli8I5hkH2cSjXksz0b45cSv1
3y/6osjtSIV4DFD4rABm4cpPfDMdkSp3HRhs6pL1tinqO5ztclZ6V2nPlWbdYROz
BqJTznDfjnHXFrPWFII78O6tD7AcLbqCXlBfWdnIv7/FkZSrkpj30wJDQrO9vKxh
bsUCJCtslScLyVGfugv5dwzJSu+5b3kewkH32is9t/xVLcG+6alKxqTs3NrL7nkG
GEwyQsKKDXghNnr+7ohsCr9AV4NhPDlyTTP0BlqEJUigLBE7DZ+0sKRF+6Oc8XMy
VF8g88offsSPi6hpWBgrG2c8YLuLsVZ1PjxmyTgC/1+gLm8V+BvUqv1F/DELMRVA
HhN3ULjEq5f3b6nSRYNSO/uS/vqlJhuz9ypJ4dqVA0Lgh5aH8CZGayaA+jxaYfYH
liqyt8VN8isofI8I/pkxnd9r9IyWg3iIMey9QNZQ36BPJFWH0/w8eFO3ZLpl+rws
clrKgB8Tj0vXYWd8io8KXe6Xzqz4pbRWgddEfJ/wPXUvLaVFI4Ld2fib4g189QyX
kMk3LBSFeACd1+FC8JAbdGaTXm7MiR4/ZVgNGDdb4CHcbOm11FzWfdmrWaNv77fj
28ldDlS39mhMafwEz3ir1YecpEO5TxCmRLEn699VMu5zaO8WrLpE8PZjrq3umpmD
1S1T6zv2OKt9iZqdcVXEO2Fl5rzG1GvqM4GTLx9h5bwS2aOv/tye6zBAfIWIwEFb
1N8mtvbUuq92MFmYrn5ebCs/8aL20U8aE8i5LJsc3B9rdko6nBLv+1aBc6PvXAdD
sAh2psv1x7dOcS/YW87LYJBPDbjA4uWl0wbOckoNgByM2HpJUTGMlPvXf6MwpAJs
ZY9knEnsSSy/5Wvm0xY0x29ZJj1MKHctww/+fUawpUjKYYPrjXeOHbQmBE7+BwcU
unlQkBtf/OPcJbd+RnVzoYVE7Ef14uzcXH8F0jVbefm59eCbTGg+JJCOqWdeAYty
JaEGYVBXtkl3kqjZ2DOVSoh/5sesegjUkYMxgnTlbVclv0OeFdF3noWrJ0sC2C3b
YlJ6D9YqV22TVYwlPcL1Ti2k+Zr6la44nqmvIJUj8OditA52PVwxkQ2cI7JLJTf5
rk5Ygrtv/I7OBY+fRI7DuU6cTrjMT4ibM0Fk0l/W8uhlkvAYjlCoeOWyynbW3NsG
`protect END_PROTECTED
