`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN5VSZmJ33InzuCy1Ud2sRGwTPxJI0pvyxjvPKBezcp7R
xF65PjqJZoT0M/GbenL5DM8q1zuHmi0vuJ8zFkHdzsfksco7o4/RVSrx0HSnEL7j
gFp61SAl7yiRrT8AeceiMKRNquzbggGioCpMgVjTPdmRBkTX8gfvctHS9smElMg/
/1VkWWWgzXEEIzk/0twQZogV54NHV7q0X+el7m/YjAdu/GMMYlSX7m6oGAXj8jx7
+9uPAzOkSkqcM8ImH2+hyuZ5FFtbMMUOQ3ZzX9wEexjQrMRsQUg3jf+PNQmiJikB
7r+pJ/Ri9PLbbPpwtxWQJMOZmln0fFJf3FeffkbthTSwDjTazmOOmsxIBnyqxBUB
inOdurTEW4VYU0NSvgGEOg73pZBK7JkShcyfxWmniPqCTHmlgvdwyz7DD7KNZNDe
wAuIuW5BR9psHDpbPwhVHlEUSlCazXe+4bjsZ5vb1MESrweYYEXpYofUWv1DJ6zB
Y/BF9mv3pYymlURajHJeqY2Szz5xhdfEApJbcIc0qUJmF/m6ijpnmztb/DaG9zda
FvDL0wWtudUt30gz0L/eUwC49ir2wt/uiJMCLulLcfnWZwyBV9rNwAjGVB3q7zXD
fhN6nNppXBTitGXKEDicduG5ONmbXXK7PVjgcdja8E29Mu/rShHkdG7BDsZiduEE
xwT3UV35VEbbH6tbKJ1jCjf8ePruyvMhKmrW/umboJW6ApDHRrPLryryFGQc8pMn
9rRYytFkzUbQwHV5DoRemInOp/r4Q7lxT/8dQXU8LMgmhWo2/HBgxX2iEUFDMoDi
eKbXR5s2Ag1ecsSMm5QHHDL72TLSZDgoZKbv8mhhPObKs7ZhBmc99rUC1+M264wa
8nE4mCtg2i6/Uo5jH+5uF+cX7z3jYHORLFDksfIHrKVp+1eFU3piwLgefJTSc/U4
fm3i0ZHt3cznEb2axL3NDOLu7gE6xt7WY3CSUOwwiPpj59LQ6PUtTVGeOdYDeoqd
EGjX5rPN7iR4dH143UC96Sh0MF/jkhcPEpc3nZcJwkSIC9xwhwLE7uMRPqzQORWl
6ZaHq52gJV0gRCfBHKYX3sE8PYYSU5C2VhN9w3n2jlIwTCL5AUoolzTn4cfhAu+m
Ifi44lBL64KWFk6522CC9DN4/WBDnDIHVWNkByd283h8uEGZEIISCW+DcFH1+kSt
Yry1CPoghpOddnv+25JtRmbtY8f+sGYjh0WflBWEQYQop4hlyBG7/fEgbEsONUox
DtH8s3uymLP8649yKPSzgzENjk5Os1fv+lQkrAOeHYAhR75p3dMbtyLlKC0Fui09
SZhmCReV18kQzntCu2IpWmicGKBzgNvcoNbpM/u3mgIUPw3VkZUnUOyIQ/mdusZV
4Db5rqDHqNuqChFpBzKuYziBzDnq7BFJPLTAlrUNctsM8KMSe8BiJ7ZprjPS2Uqm
qSJsFy0bOUd3IQ54Ut4bOSqsFqzU2QcmFNi8Jzc4EyZoUk5fgpjzs+H2OwKRI8Dq
oqSwiILYzMGg3mOEPUjzmw==
`protect END_PROTECTED
