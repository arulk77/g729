`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB93DQ5Pytfqb0ZmmrRnyf3EEGHruoOljBk73otdSzY6
QLEw1xTZ0YFwYJzWttAGFjVV/pdsKqig2+npiMSsmM3QNcMrkx83B90XGuM24EE+
VVZWgw9yVDSWaY2cqKjyCzBiOmqKPQvbF0ICdFSfgDeOnLEf0N8j8MnfIZK1xM3H
`protect END_PROTECTED
