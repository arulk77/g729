`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHrRcyrQCI0DsBmsLYn5JUGg+srparjrrswGPI6kbfZz
9UZJ/Os3zGKNvsztcwTCGoI1uyLbLEDVnCSl7jIvlv/SSR8u9fcx9HdiSyWbKx/E
PipjVXBQMd1TF3iMYZLAYJZKjIVtyxPK1PP61rtbEE1IChLGueFXUp2QqPLSd7Hp
TSQUYw5KAqGpVQICibmTwvmkE026dncIgwrllxLiyDA2M9aI0Tl2UJwv+WdXFD6i
mo2Ux6uc+CREzCAvIokOmXjYnJlZnMO6Zs1csWYJreXEiWi0LmY6oEn7jezx88VM
zjjUhuxHYqgYK4PEwifKjKD89K2VmzMZi+MWNgx8aM5dua4oUkD6sz2MJarLyTLQ
otZs7H0bAurd1up5tZYJHOewsTpWjtwUGNErziXPCf+QN2kxJcrVS9kd5Qb8F0IN
hlKbmTPX7uMuBRp0FPByuzQjT+dl5Px/DunbFkPh8fGSPRsq5cIoakqc6tckL7nm
b47UkvzHc+u8hGtTdw4hNYRN6LAGPjwjKcxmVWjtohH9dVAin7AB0ToasPzIEDRV
`protect END_PROTECTED
