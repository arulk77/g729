`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveENDutkDJESkI78gjU9UfFqtlfI8iu65brlxBA/xLrRB
8AwgSMqwRG8oOVeJngGBfGk6CNrYvrVC/W5zh0YbHfpqU6wX/5x3trv77OQqTXo7
VPrgTYt+ZKMkvllk8QhtOfe34P72L4Mp+DPkomVZv5qQlWcylCRgWRENUaAd9Duq
B2P0V4m7hkr6q+md5iDoxZ8yKg1LasMEpLfb/HabL/TfRZtq3KsGGEbmWOKVmEEE
ihIxsIpwG2TeJCgupH9pEWVRtyS5ovQgHnsF8QVBZxvnDivVr63xRPqS9ISXjeMx
/fOn/0XAs2XOVJsNpLrrhtp6HViOf6iLNW+SKDlWOOvMwXoKUMrcuHbsBrbQIe3+
8IhISMX6igr52bMo4epdDG9PuGPeMUuZIEmUesjSNYN3vj14rvskxFeK0N+MYxxA
58S/WNal/tDL9l88q8CGRVa2JYiP1+62x9VtkvmGUvR7e1YFVSSQwm4KsqfCtAXZ
owKnMIz1lAYOJI1cTEsI4GNePFK+Esme2aBuhp+1qjnvHHg4AC5U6LhkIld3zLDq
HllYushui8yZBVUt7W1xcw==
`protect END_PROTECTED
