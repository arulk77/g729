`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDYj95ipBimnJrDczBynr9yflIb4ruma7IRSolkk7ZlT
tZdtrvKCdxemNWTN3n/rxP+Q2WFbboavRWsBjZYK9ByIFVm3sBg9LZdRTufZ9I1n
3oW9gGEv4swQw1HTYUu6vhjecbGTUmA1E72bLgPNVpBuKoY21j3I7cLqEbITFfS6
5qQsb5nPI83vkxoYMn/dodyReXBCeQvJE2LN4ua8fdPGH5KzuQUxDkapAdi2qSH/
r1JSjUTXXaidgIgRrIl0GyZVXKiqpzMX3BLt5+JPVnfxmkJOFttbEauSU5uV3bv8
dsdaFq3cKy0HwTAsRWRWITtHgcy+IVcOpaMGKisAS38UG8gWUONfSLSCJYOW2yER
l42XRTqOLHwVGrrpql4bw9jzILyOFujK5jB54xGD/5ZfsylMJj9U54S2hBvj53cQ
vemsn9vV3Z0RMqM/HKVEH/JDuuZYNZK3MNUliUevJ0zsSERLUI+ixQ6F9yrC2SFx
mfXAj4UOeq2Vjb8LU8j/S8UBAP6v7s9zoT+Ag8wYzKxwqzdb5EHKGu7+4FeznK0x
rNPnYuBaYqKBwdc3L0+akZPKBZ6Hh2QbNIKKcsump04j1jgEejAMo53ee/Q5cwC9
UZ97QRY4NC34Zp5ailTV4FIg+qH3fm2wUUHVuyLVfCOoMmv4whD65JvcYSwquHXi
`protect END_PROTECTED
