`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47J1bXcO3ydOASQ/YF5WxdeHI+HkrdPKEFgIXfWerObM
zkaTfA1LlSCb4+kpf8ANWlP4fYuB5f+xLAz69r2pV+8JjBGj/0XOu/6Udmw2t3A6
t3G2h75POVaYXqVYzFhmv5ktkynpcXFK2Q7kfsLaWet8LJJkePfo9DbmS5jI5PSH
hjjIW7IrTJVHvmkcWOSJAEfegGYYorBWVQK3XB/MYyotcKaeO0Z3fJWrZc0VV2yY
L+3iR3+5r3LJrAqKV8whlqIt/DuHivOsFDdWLWr7lAk60+am3hJgeofsMmNObsi6
tvAj8xeK884yfDLuwAeVHM24S9hHx+LP4Pm+hdA78hNsusjnBy5DkcegOPe7i4QZ
kRKzR94aKlYADvcfAanQ1MypOwF0l5bPLLmivK7ZfN6/DhH76ATsK4t9MD+A+k76
XMHhc1KcSl/fBpLTXY9/vg==
`protect END_PROTECTED
