`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP/iKqeTedReyRZMC9iuG9nvKI/rKsgl07ueU1qyNSjA
JJCD7IFOsvbtBCskTIObOE++5rzuge3rE57ola7fCeZE+qe0/uDx5eDHCGiyKYog
aoZmMyOCH8POEQuv7ftJwPeXgFdkD7sPaQqN8cYotBwCmaffWJ/+J7X6jhxO5bas
0H3h3YNspSwVDnBdGdrTRTq613UHEqFWEUi3syFbBA7WsAffE/M/v1kKBogGE5s4
fBMrInp2FrH2jihw43PfKobdQyP7XKHx/Al9PID5zB9N9gp+pX9jOWJrCiercTgl
bJ2p4PZ6+8j9dZtOgrf6A7hI0qKVhvCeYlbTc3QMCOFj46w0lZoL3runcNSOUhI5
0q6S947GCzWnegU12KnNxPy3xQpl1qju6jx/5XahYLViVOPvZ1n4LqOrMgsINWoE
WIzO2LCSbVdQejW9yMERs0CUkVakUKp+rT5EVKuJV/KICrPWLLsyzqhd4h24Vo3u
VTUK5ogNxh3CYsADk5+tCNB9tq+dXfbrrbSIf30ymDrLfE6qQbj0BUAjjVEu1SP9
bINGIN+dGD+oWOWkSHrh1x73yII0w8GYfZtBBxc0yAsCyHLQsTM8EqqWD9cFBydd
kdc3mlcnOUMnC0sTg0jwyl/SL99lQTqHPWqaiJkE6Mmza7IJRxh7RNoF6/5GdeKs
+FlSf9DLlmUmEXqUngRxShpdQDSGRzTBdmPchVudz1s4hjxjqcD1ttO0rLa9Mpbt
8vVnbj4hDvIaM8koiV8MudPi8LeVvSTFFfOI6xCtr4ZLStX2sauQPXamriYhFLH2
LrPZV7IrD1i8SAWnuI+++osYtjidXqIdFNkDciwn1hBFLtQoytrN4icujM6jCOaf
HCjorSP+k5pnfK3SVo6eYOA5gRTGZhxw5wdk7fT57GGzUHHMyIZdzCGZ/Ew39WFe
UVNECtzLEJg9uM8f/ybqLEA7hdN8yuG4S6U+kuul1pCNIqcKY4wGUnc4APBTZ/tn
CfaS7tizkk8+iLUT2XeH2AsmyQ2z/jUBltvMPViXuA0qtjr3Wey0UdydJefW95dN
LKDTdfiFh2ACk3gmBI5IozqUrR0i+K3XwT7r7BOLYyg6c9aT7ly4d+cmrpRHnAvT
G2vxY21DzFkS8+LmhoPj7SS6Bb/kDoQgNUoU/pSLNSaR1zb9VqDwloK2041zqWQf
cT3iXiKgtGD91ChbMPp18iMEEeVqjpbttO3WaRfCwF8c7kohAF0C0T0mvqxtXC9n
9Z8MalUAxDeCptSXtxlgQbP0gXspUKuL0rBTUx8wSAsBEKdONHilc4pMjsTKdv4q
1Pzhn9ne0vn/5Eaja0xmJXXPf9wrmNiqVV0zOMJXLtqpDtVo7BgH7c/n21ezAu2W
z8CiRme65MmR68zjHpVWAHVVs642SXLX51yZeWE/roDlQ14/S75ac6tZKZ+qp4xk
hsoLSaf19VyEdCjN+QCnk2f0D7Cr5dZOZHIgbgIFxW3/ZubRI4aE3XBIwGvuQjt5
j6hvhbS+lTqCcrDfMLVnJ/M78SFmLEgmAJd2jT+sTTUlYrvY1rwNdS/dPb+zP9kH
50ElNVkX1PgYf/e5z4LlPA==
`protect END_PROTECTED
