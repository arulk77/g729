`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pbi+4Du0rxd0+meswZiy9iubolyxudDCWhY+kqOen3SK7KpcQYDeRQSA4tHQbKR1
OqjjnRIjFF/HxB6xJ8csCFjyuJKp1piNzBzxFFxYejd169cqwzAer6N3lzqD5Lm6
2Yd8Fn4RXwsezb9RKiC1iRX/dr+CzKqW39R+tvw/sDFWEZfsGBCQLd4LHN6xfuSd
r9cURN1W1OHz9akiNkZph4nncYHLrh32gIKk5ydRoK3cvaTvIkWIt1G0kn5mhNBk
mKwcDkx6Apv+ETTv6P1PsDz28+p0BmsSupg9yM5u7Uc=
`protect END_PROTECTED
