`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAOPCj7el1PCbvRDTEeUOgJcU3nQOJgAZMa2nZkFUsO8
DK+xGlhSaa/IPINQVYdg6pIrTkrNEzTEK6KzrAeIptvrTOeIDcsdOWCIEeeetNuA
YTi8JjRl1cx7nGNpD9mA3A/gkLMK9W0G5ApsAxj+Jv1TyapB3BDKsjyrSqRWGAt5
MFDf4hVN1crx31//7nKJAWAiRo/N4+hSuJXTiTnQs93LZLt0PAI3qJeNi3rda/pO
DIW3Y8bHo+9dYdj42YJEvuyuLbydaR9ItU8bHpmVolbbgbJeJqdIgS/AZAWjZx7g
NS0Fw0NGF8EFHE7J0KZwjEJw8sbpoC0WWv7EB9qRvIqJJS9fo4ulEpBYTr2a1D8P
lBNRRP9U7ZTnfM3MbRMlujxJ317YWmnFq0w6E1GC0cpAJU6S1vKiNkG2V2R9gZt6
Muoc6FCNoUzIcdtid8C7Bg==
`protect END_PROTECTED
