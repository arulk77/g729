`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGb2cZNcCjcumKJT46gKTnHjGWkNRdDXkOJ/twHgbyIe
8Q1dwhgsfLOj+n+U6I0/S2OgRjQwo//je1egkwVea4hR0HxATCg16EOs/8SEBc63
OFZC8z0eULvBgzzX7oPU/pZk8FExx1+n74IxorFvDyPg3j4ebRKQ7KhS8gtnW5rI
HoJzk+LfYSmk8cNhUK+Q6g==
`protect END_PROTECTED
