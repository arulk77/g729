`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMsCgKBdYd4KNrqydKZ+cuwAbKNm0SpJfCdL4x6zUNvH
suUsedawqn9IGkDKFa1FUwZAlRe5M5MQ6iVtO649RrCckBxe4SYPQg9Ly+X+24NN
SaOuSlBiXhLahVbCvwJju4sk+L9STNQOxWS0ERxDljvp0ysrgKlvMfLhJ8UMnWCd
QIdWoOLnfth0fNfzZyJ6tM9vr7VD13F+ErlnybsfWuacF7sbihLIprMT4vUC6osr
`protect END_PROTECTED
