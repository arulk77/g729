`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1adgJ2Qtw/DUzdHhenTZH7EqTUaZG0pEwv1ebqcePALUL
d8XVEX60Dqu+Xa/Uv2eOLKd6uvE951NuGrpNjvxGbX0mNDzbsdddMXdmBdnsGeoz
C7sqb4x5gARc1rkmwD90LlVk+FnBNFM6bTrDUXM4b2MSWwPgvcmvaKDvNYMVcNGb
lbESQzJUb3hZABt1vx3QrPLASpCXMsT0MxLxr5aj3hMIceJMKzHkTZQEaQXEYUzZ
LmEDyAAeTNGIgiQuRmf4lrj58IwQ/QdSKWWl3i+rckgDvdU/6o3bSO2q0GsEK+5k
BOwFwfMkIZhNk8lMQBZiXNQsq0EAibjhWYcFxcMhbssbgS7uRpQx7tvXktc2qk3n
8zgEpJueyIsP11l1oazgFMDtqwv9ydY1R3kreUQfTgt6gEYLbk7GxJQpbc+HKuLo
gbkO2va0UTP4XAkOPFdt/PtEcH47jcGMXBQYnGxIAkrm43X4geDdwEcrIq1gz2Sn
3KXXVkb7/G6yLzV/m86v9Qiy3QZkK2/MhNzJ5kGYPTwOeICu6bg+FeEAkfCug/Va
iZYPQljOCOQ3H6xuNodvsQBuFjcAdkYvd9782z87A0mKVFZKOiUdgqG3BqxcFI7G
wx6Zlb7DnsDHHcdj31kueA9QBPFnk/vTAEij2khflPsYPvWdQRU5kQyrLR+3iOl6
ioS1tIP9WkMQfI364ddtlNEufs+CClRRKuGMqy4++jQ5F4uVGjVMBQFZamNercTC
+qrB8pIWnCZyso9OTtdmqz9p3G2p0dJ/s2wcZYdkMlpuTudGXvSAJJIvpbtoGVg0
vLkJrwB30lp9ZbNxy3Df0ZUdv+gS1ud5+jk1ARpnzXwiyvTnV0ODpcjedpRk7ONb
eiSd6W/CurGQUPVV2mCXdx/dS/qbf3yCKFZgYk5ZwqMFL+2l8EtGggNVNf3fIg5W
JyReDRregHiLaXBfdrrjenfkvfAdKDCRGw6potROj1ThyhWPiPJQzUka41b3Ufsw
0ISl6lcJztEwFPEVsZWIiMgjh4x4gp4UkbO+0lsn2fLGLT09LEB5eNTPXjLCNN8V
gaBDdazI7HlBPrimrvYe6JfozpljMEznBimXjUNlR7OI/vX3cPHixDt1tH/zCIzl
Jm3h4rckpt5AAcIA2SfUr62fauiD7vpam+0VM6O+i0IB14+Ax1yi+rh9U1Kx/GgC
Fr83u73j9qDMIwSUt/QQH718WbbpJPY7zp5dY1z/IPKysQ41ynUOOg7c7WC4NAoG
xYX04QS9g3HQ8ZLV4W0t7fz4NG5ypUM/efwM3yjHOcaQ312ChLKKDx1y8IDWv8V3
6llnMgT7uXaE9z2CVWkKqP6+yODP35RRtICyKQgGtjR5HjYZWO0m9x5cBnHJXImW
2TNfu9EpOIjgI1VjhGeuDDcbp8M8VpizIYfwuevIOIzZRRyKo7dHxWdzbbOPAkmQ
72scpkrlMZ93h3I0sUMqgnz0M4sFHzBHr0f5NNwBgZexLyKboypDQdam5hstnBgc
G8qWGbnipl2nQW+aUKbzBE4qJK5JIQExvIyxjLWcKc4KCJXHohbKwjPAJJzmgvvY
MBDcpYG6IwLzlROXh7QOPSbCdcnHN31GeJ7gW99Bo3T/O0KLTmI4Tj3YHC//Syxa
NHFoH3j4bswRftmyD6e7sVlOwzm52zqlUAywzBZ28DTvC8R0a9TGPL2GX5RJ4qbY
dmk71yQO2RvOwzvs8lmvgt3ofzjxZqeR9ZgFmcygG9m+YjMtUfPJVecuMxhL/tIR
nUVwDV9nVHDbWDxxv0L6yt5JTOuA1FWuF+oXlxHeGRJABHAOKhGkUqYQxrOHTG0W
JbB5FsUH4eG/pvIodxBkOOmAhwcx+BE/Atg9C95LhKEf+Ks3qa18Gyxby2sorr+7
MUPu+LIZ6B/90AW60imv5PSXuOdb5AS3Hbo3owYQJAA7J2DmzOkpk4M/AAOuE7XQ
WbGHATJwOELvoeRm3xWRwNqklSpdCXGCtIXvr93zeHBULIMCM/fX/tWHx1Je7R3A
QHWu0cNWjBVzx3bXUZRQnFFcenEnII0tVTSlpE5mFlVQcukDbxfyUaySglWvuGBm
eEOMH45azlq4mL/dBiYLmqb2o8FY4nKAUrzspCCuKKEv2Ma2DbM8p8gChQ+TJ7fb
PhWQHy9GP1NSfJ0Y0qPavV1kizikKj1R4HUa3VaoK1DSvrHTuvNHbs6WwR4wK0yP
ofMqyoSspkUaImKiHzz40HOIw5n+FC+EfkpgvkwYPlvYRkBtVIw1KxXltE7EdYgx
Y6P09+SNtaTse3Q9GoCY3ukZG/ByhnX8GgT650+9RYUARRD/J0M72O69mLFbAMwS
CZxbcs3vFHA7UNUQWPHdHvMakzuWS9NcJhYAxf2UKJFgxys0o6x3GKzXnTGU3Jhu
GqQPPyHya3g4F1kGjOZjKSlISnarZE8cu+sBHT/4MQme2rmu0ay2QQXtlLtUXK1o
O6vH8bduH5QD3kHbwsIyQ3Y5pajq14LZoXsEK22lHECFxf+Iy+oliuO0KQbCXGm7
5AyfxjVcyt3S5fIuHIAhkAYvdI6q5BGF1Be2dXN5qtISclzyK7ZktHFJMF2sTQxI
cB11r+D7PrFJPmPdCBAodoSX4gjwr1cILv3SPpDU3jE24cy5Cj9oLpPi9thfFnys
9+kU885+tNPw5Rj0sGKqmiPbTHEkGBH37YVMDSrTjzDDyL/WVxIwF2ixXYDJ3nK7
9LJ/5IZhbYszgxitLyESHf6NOTomfGFhCWfCUM8qiXRG23cntcuLBK4cYCQJWbaG
vvXclNn8au82/hD+daqhKkjKz40GiPyQC6ZNTSeTwYfBxhyHchXR7ULm4tPiZrMD
wyGn1yx74T5XugRGkXNXlkWfeJcFRxxV2gawxE1syk7HbiCcME0KhsFttQBQn/iM
0ZKxgwM3WEl9gNd4dkxNZDMhsxYs5/JIGQ9qWj43c0zZkLNF4K9tz4+bmdo4ygPY
gmWdMq3c5rnfLssPFw/HL6Ka10orLJThZ6APVYZJh4ojE78EMTh8wfvNTom8lUN9
+qhm2XCwHjcQhYsZF8Qf0cnqCe3/iEhKTGnJ4XsJEaFHLoGV2tv4OhZIFJfJ+zGQ
oD9ZTCuyxKOFDCeBOrVK99A/dDDsKuAWPz0Tw2gSBNPkaTzLp/sFUR4dPbQPrUou
a3QvgnrVQGJRI71KkhhcDfD5SPWJJnL7PLs/ssE48zii/C4SLFJm3+Fag3ehN4F5
woeC3x3SdfvoEV8gLfA9NnM5c2Zv6IyM/dC9phu14Y5tODijB6LcDOyPPmnupEjq
4juQMDqANW7hs5hZaJHSM3Jz6/AXX1etI3erq8PZxh7TeaEtAyjEUHaeEhrT7MJ0
68AsSkT8KyxKWz+UI/5V0Vp+R39xyOKlJv605soaYO+PVu7NDj7hj0BtZVUED2GH
5zwkTHdb55MtbOvVHIYQWMEak4baXBDa3axC56hiFQEFTMv88itv9yTi8D/b/dOu
GWvm3aPTdfrzB+hFS6uuBeyh4IwMqmj+aekfmoayx2g+HR080ZjE7dBYMISuQf3v
ODo1Rj2VnpaZACjuA+eLmKTHaExM8W+Lzt4fRtuuERhGl2onaiJi4nqTzjcSDqCd
9QFKWkm65ZZB1NBzxqTRULQmI8MZhJMloxHW8bBJdD2NTVCGN/ngtvnlRqE2BQND
W1/FLVMP9OWmfbWTAxl5urpUht28cHNzcGBKG+xnENwWhrRY0ybmUbK5qqvhrV0V
9TOuNaSyFw1MOd+Q4jrG/axcTr3ek5hkwYP78Hs9U6t+V2eugw+2sXvlwO9r/RdO
TlB1D5kvnevtEcnpw/6QaqZFmh0Eb92i+AW3EAGT/XqHqWy9OYfPUGJVEVn/wesZ
XgfXB2MZl/2Ir+J4L1uUJZmkfJVybXSucHk/xTJcA/Sg/anso6LmzZf36jDO1HNj
5PylL2WfkY2JJ79j1F0+ICYLBbzXoWz5vIROKMjXvkHhe3jPfNlD2p/ELUbsUvQM
OZFjumHhgWcDyq5G7rqUFi51iZtksMrR+CDhRC8UDQpva+3aF1gx6h7LcI3ZwIO1
cyhvGouNhTLGjlqEkKAJBY4FZ/W3QHYAqUnMs6+FYySV5lpRAGKzcn+eWH9zlYxW
UmnwB92PDkIe2KqGHcNLgV0l64Q65BuVSdrecQOepCkCl35NpevsR3awjFbMdHMg
PNcqc1hye662/MdXhnt/ssrO11NddxWLoJocn7ofuObPqimmTEcYtKf0YjukFgNL
bdRZtRnilcaCquSN/NU70QQDGIG4V+OqYI+1ja503RXpNTfBQU3wNkuEDOWqLMbB
v99jswABgd8RwJL27e2hItcLjiSH6+KsdXv/NnEne6oYH1dUPNLwlt5QCL2AYLF3
r7SmB5zIC3NtgHlHIFpefQDj8nc2M0m/niVWjD+3wP1JwIubcymu2QAYE/mfhWC7
7OBgeyh46skRYV6amGRpIboozgbwG7uEOgbfe0Vtml/0MSoXfBLCyUj7i4tJIPA1
MPrl7/JHR0doqBWvNDvHpkz4wqUAgm+pcwUa+ViEk+PAdj9x9gqPKwJSaheN8gcD
931ahKGQ7sdgPSNwJ+5e0ok07b7e7kkakke2PPZjTnt0L8zO0rymCXla0brWZyOp
DgKykPJUPZ5N0hS9mqZp7a5DGTXCbqEZqtGf3T40mvX7/l1URTqvtT6mHq5TC7KS
9l0jhq7G+Q4/ex9jtj248rS9/rsBxYMVBiQ21qx9t+fc3byiy5EQrV+ps5YE00NK
VXaCcFVqRMKeRGAil1kOV35xJ2lkQQNAW20PZSuKXmu2Ffq3bxEEU5LAeIB5oGre
kJuXtoJFg71EtMGGxW413cp2SQtYkGZv0m6ThHaizzHn3d5j4PmHiCzN8LN7jW4+
Z/m1N7j3e5bI+LXl8aLyndpYSagXo/cctA3uJ+5HUi7wpHcF1LG7f6EiDcTN572k
STqT9Xi2OgnLMwo/BPmUsTC3QrQRSW785w2kb7fG275H9Dm2p+Vjx9op2kvaOGDb
0+SjUZZq/3lRXNAQV/VjTwA244pZJjXccYMcIa62G4wpmvwKV6uUcJXLjQBe84yV
Z/Bql0iUVSMs1ynJDqzbTpRihVxfxpLMmNdsoreaGibTk1KpAmwrMTmYQWUguNh4
X7CKiv0a0N8IfVHlZYgowICx+dfq17rKanVRlaPnOkQAjpVXQrrFEBgjo7Y346z3
6o8Vvcn2to3UPnA8xCtEZNargYz7Rf3KvNZ+sm5S1INIc+KD6HFD7G3gt1yiUz1K
jH3iEwrlgUm9pc9NXtFXI7EiM3iFjUUGflhydiJ5UcYs+uz9ifiCW31NdsDvN0Ly
jCZwbVjj8pywDMn4WsTnz0KcU2p9comEVIZdkgoa+OKssFgsUYbWwZhceOixvdBX
NCZPhCBP1CfAVLZoHVwcB6c2wx4Rg9H1EaXGwEJyaaMHiuTbcEcQfl5SxOdhbQfk
FuXZW52gIq5dSra1tbKu4v4qKtQCfK6euxBX/6meZ/67M2T7x/w6yaKAkbSRa6eg
b2+n9K2nKUAtVXXnPcJZqKLOHehvS7bWnayAN4v3ofmaO3ZUD2TrQJZIfntCvWr1
SDlKHqRnob5H7crUEjwn6jJ9u8KpV+i9a1r8Dh/Uk2DIIa+3+hwEbST7Afqk4vje
MOqy6wTyLTxYriObafDftVjhjdTOtqSYd7QHEyvWj2aMSJNybhl/9FN+uQ95NG1i
gW7mCZeYjGbcOwQ6mrFrhgCfhMpHYoZwfhJEL2UdreA0HsdHvEbUkg1XEakpdQto
6xE3FnXeCz1nTfsWs2PD3whb+GEDQJRh16cg/um0L4aobDPQ4UX9T44HAHxI1mnp
GJ2K5oPCPu8gZNF7gAixSb1924iya1h85I7bcBfhbfhh9tzXb8lKJuHBslYFi+nf
urS+z1EcwaX3onHqHiPiwX1j/4kZqyz6UbAUcp/HGTT9P/JtzSZ0mFhBgEr7DDBb
vIEh4XI29EGj5Ra42dJOCRWRCKK2xn9VubD71pDJ2kMjSv1u6/yoNdcKX9W+EsS/
pwMQroDqRkOrGKT64qhxhOhov8OKxf5QYiJFEOwgIHBwv1UlfHqfBqdYZv0Kfjgy
+21LfgmxscmLH/R1zvW7nnX+5zfaJkReB22td95r/qdtTeuboAu5wxCPMX6OhkaC
`protect END_PROTECTED
