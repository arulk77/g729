`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOC/WxiKNqacMtuL6aRhjItLM9LbHRbJLNUGjuGdIhq8
YcH7ZM7g4MAH6OFXgQJltq8h5z2oCg5tw0lTp2mbd4oEagaAIyFbLsnlyfdZkjX9
YC0P2pHXAfHGmFwpZc+8p9hfXZFtmuKo6GaEwlm++70fiyR+ALcKpK21Gul+c0yx
MYJ6x/ZUIwmTEqFyTIyLfAoDAcIx7OQdIHY+dLvXxtyODjH1DK7L1uCoXgdgYJk0
UmzQ6uv4a9FbFwMz49bqPYtbr8Cpyq5eAOX8DkK9iVZydcxjDEWGGMC8LOl4El0w
qnxuZXPo44dcUngFoxecJ+Pt7LUVLPjR3eWOxxc8oDEFTeA158xVaBO4ejoV5qPd
azHGKjXxa4k9Uo2BHQ50S7CD3ZU8HJ78M9L69qjm26m/E2jrskl/InmG9o1F/aTw
QW6WE89dgYHqRyEdY/n4Jj6qnJKeKf5WOxavnkxo8AwNK51FZkm6dy46xepdOzPQ
Lwa9L32Oo1FJE+YHt5jtPkOkGWJa2Kd240VHmf34rsoMH1oNzpDOKkM5WdYMUcIX
5ncJtw+FszyqeAFRgBR9zF1kghAkjKsNGFQcQPjEO/kqrP7k/+h6y6gGkLTOepju
vt8lF2/ovElcH4gCQpZISXOuqzdyfi8q7iQuLQUkVd7HzFd/LGZwc0VbgeU1EkQJ
lqd1JVo97qudE+lLzlEheWQOfi5iwwpaNW6/EuJATYkqPcr2JUFZvS3xUvncB9KA
gYdZDxJcfRQ7nbJEVCb3BJvCoyTIGsm51qF9nYaTzzsGK4O3OhynGw8uq2Uh8uIM
Yqsijbxsou3yEqMuQDdU5pGeHQjTCYlGsoWf0doZQjX06aH62DHYnWpiw+aY7JnO
G8gKneUQsE3yW4sslK/BPA4T5uJdzdjCdIlOcekyejXDqJvCVqGI2ptG2gjyNZJ9
Y38oeggj4b1G9lcjCCw+BjZROYqVRyZ9IoB5mR7tZiZIAT55mNt8V8iZS2PsifU/
MZo6EZiU/HUGxUIuLSDZQQ0JNXGYtsTrjTwJH/wbhO72KAcOQZcczKV95lJoopP6
0BbbflC6obGLycAFp66NdlNnEF/NCO0rNmYeHVvGhVs=
`protect END_PROTECTED
