`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41P1o1ODNckhAsMQCNUqu4F0guJStq31jvUgOKHEjNKu
Ew1jrlOTjDGYX80cXSikatLw56jDMcNb6Hn5hKgKweT/gpsmU4q654PY2pYC3MWd
510mwT+GZDUCjA7CERhhXu7ET9nJrb8bh5ZMW4kUxBpTCvOxERPr5oTa2yBnNKtK
lkDwwB3GVpPFsyqWLfYrk1k52BYCWrzz+r1E7PKCoMtpunCi1aFHqZY+RQ0yOepl
5/VDlT1uvNtO1V/fHEPtE0LblnuB8Uuqvgy24j99qrrmXbznJuttpmHcMJuG8u0Z
7Xneu1rY+IenYZWpVb/fCQ==
`protect END_PROTECTED
