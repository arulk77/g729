`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mco5pq8lDAVaY9tDwlnxHwoTxcDXHDKLeQRo502q62i2PLuVsvJe2lCvsE5WJLlh
MWT1bYBo3jaKVZPAM1/hYl9Wg09A11ER4boI9ASM/Xcor1L0lR6Rxw9ZN6qP2pZ1
RZ3T5fXP2mI71U9qQ4okmNB8uQOyvvmwUKPSn609fWFoGH8HbvF4eLe3rVyeuF3w
HcOdHJFHnOmVZde5Uh+fqxiT12zDjRfCFLUv/axc2Dr6j4XRLkY4WAT75rIPnnSX
n7CciiQz/LL4eE18ca0sTarZgBeJfl6u//AvEHIjRJ6v/nW/Ly3wS75LWTNQr4M8
DQJPZOoZCR1Ey6b7lFzOWCQet9WrtfGbW0Pqe0fNOqk=
`protect END_PROTECTED
