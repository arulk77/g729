`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu470+oJMBnMbLil8/2wbQAYs83egURdUTo4b94kBiqAoD
m4TDvlhjXOIPh0sYqWw8eKoMrl8O588mCthiPjdjhRQ4BLWWyWEE5QOeGlT+N+Sz
Mjtth0IY+LdpjcoW4mL4nsdgOOqTN20RSXAxzQslmAbDhLRFHja01Ah/K7E6V6CF
OPpOL6PZwljnIdvKfsgqLWKvXHlM/PSx8W1r6lLzWkeWyq4ysdOEshcpIydWUWGV
vytO0YSQzFsWXU4IzNN1tS4Wuxqw5H6hgzzqfHGJW8m6ru8Xcsrp6utesMPI+mUa
s+2SuDN+CwV9EBtmUHMU840RQre6R98mlV5yFfcTYspZmk/dikSSsRE6TkWKntae
To6Vhd6tC6HvCpruX6fm3/sqUwqZWcHxYuNUaJXyyNOhzGfJBKmfdt4RheRL5Sxw
BqcJGmRKEzkLtsSI0jvfyINd++Z5xRdwTZyYe4nsRTKxSLdJHShxchRdn5749PKg
`protect END_PROTECTED
