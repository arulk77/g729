`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C0H3Q2bw5AKc0S6Z8HZ/nGPbc6nkuxvRP/+4ZbsdxUOM
8LTzofOOmir2IwfXr46rXH2YaxG5AotpqbcX4SL5x51lmu4UqwuNrtsBiKIqKVdT
1dZB62XGk1jL3x3KoOrH7rwg/gcSV6vhmCJRkV4AGJ4B7ffyT2h2DwbMBIt80fKE
kmFTBwudIygX8IRqHIy41oi82mS5HFwEDgSc7o8gyM3hAwUsZ/IkLv8dEJQuAUzy
qG4uJL2HWepxb/nA8t7aE7+W+kIWHFzUTyqQJ8oYW5WCrgpTvl8C9u1cdX+nxn7L
b5R9nKg+HmiIH4rXYVTCcKcsX0Xzb6H4c6jMMfI5EFNC5f7iHcyRgrZEnR1J19o0
pgNTiM8vKArj91O/HKDUBkRfSDJ/eoKYs8HBcT6pCSFyumZ+m4U+ZIs7XL88Cu5s
RkGEUigtke2JqU7tTYARayHEVLGxFu7z64REMXmU9Pb9iY5woP7YCXeS7KYQn8ES
t95hRAFwed40UhA0NTA/8h5M29zbBjcbHpb9w3aFhOjHGATIHtft7wD1uQ3hltNs
dnLvQuMbt6Gf6uVYHhOYaCQd91RuMqiw4nZozvArnE9MMp4cvrqMlOtnFdDmEydL
r5k3CEHDymMEW+aBA0zvM7paXyQnKIk+Kj7j29//OP60YpR3Frl6w+20OqiWKL1M
7LrY1gX1qSaZ/3wfBbi4so30gwZJAwCLRTnu7qPoueBFe9WJZHPWyYISwmvsZ3IP
4cPNc0qk4StPq/uDNYUpZXRX61GROmC6Lx4CCF4x9tKgPik/nO5V5bZ2MV2QbG7+
vb00t6fZPFGP7aqhQPAmCNN2xbsZg4S28PaaoeIruWXgN1QG6Q7P7bW44ourW+X8
9i7Yn+/+mCLBmIXpAn1hQphr1xfNV9QGp5rjOLetaVI=
`protect END_PROTECTED
