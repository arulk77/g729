`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAOdj0FT8xSWOWbMfG3k6j9BHiCfKrvTWeXHz3laBEYE
1Oaq5VYMfpSQET9i1WHpSLM5IZwIADvgYT0MQHmEYkRvZmtfXqqp4EwN9MbrGn4C
nBz1Iv1UfcGr+jxjodxQiiUkd9KfUO/DPLmlqMT0G8rTQ6pwzBv6ShzatpF++Kue
St0uzUJPiwyrYcre7hE5Rwkfmkyeke+YX0+qfcEEE7ZwekCE+kt1qb2dY5Yl5T2h
/B+DofPQp8n5s/j53hIZ5WzMJzltEQG+El2hr6qd9Fzu7VsIXwC3S/9kI2NEXTCD
or5fr1KOpe7NNA/JbnV4FYfhWuG/BM5bK7mRuMV977oJESUBWtDffl7tdfIq5tTZ
l5wxz+6L+warftiL56m07dQtP+EU+0LyF6k9NQjy1kI5PBMeR29oKbUYfQi2bwiO
9pV6/3puQ5bkORinKSXt0PWUqfDukJhPmzKR96euvGDyMkKNFHoY/YbhefOIX+DM
EBRhq5vbx/FMN2gIPO+GpncpeHyXMxaG2HFXpkwCHEtE25D7EByNQVplABikLAc4
hZ3Xrk3QMZnN2aw6BssF2ECfOGFvr+YF7z7y0ZmtiZhv9ioGGQbbjq1fEyNNZguW
mRjUboJ0HujAOfz2DVVa7NgjswM16HvlhzeuluHjDsRZY+kFjIwQliU31t6WfwQ8
j/7/S6SDyNQjir5OdEOwfxGCBaN+0Owa6NxsH01uODoJwlEO/uQ+nZbNFA9ecYI4
xUqRwxsi0TmhtciLQ+j/tWgIycS4nOhU0L2exwl/7syWoC2Vb7dddZAtx1wmJdye
jNf4xksQ+tOU8sRyBWH1O7oc5KkTWPwv/NFLbmL+Sfj8Kkt+RL07ueUbJPWD7oAX
9nEerpwr0zw+YEsAinvMUjlTinmffg/MN/aO8HY3i8np7S+0Zs+9zim0Jk6CjDuv
Kxr+kRoZ1QVtNs7u5C0tz7fb2igm0dNFlLG5q2kpXKZ4gz3fUcD/zFI1ym45Fcym
hK0aPBUgYti6f3Yxll9pa2t0PLeJXQl2NUsbmJAjcjAINZmGBGmqqPDQfho8LqB4
dmw8+MHIH7dJ/IKcYsBju/mA5iZY/9idaDv4xWJ+KRualC7x/xZ7iWXGoyt58WRv
aPLUWnFiiYSoRMm0vPomy0EKZgJoeUlEXcxwLZVRDzl6keMbMzm+iVbOVahyy5vs
G5fGSLU3Ctt6hzctGzAB+rAnjELOy2WQrT8FwlgIzNyrpaOOFNTLLKWvOKh2sJKR
4VVJOMwQTooQ9imh2xonepnSRrhjkVwxSnMyQ1QUB//t/ZNa0MQHvnMQlDozPLDn
JNh3UVBGkRghXAuYdaKueFr5mgQK1Npq6j6RbplV8wLqlP/3LAxQAtF3o5a6c+GT
Sv9JU25JkkZCE/kJowX/HCR6H6/GXqQpqj8p1DiNEcbUJhpnX4udPR+VTPRGn5EM
7Cw1KCKbJ/NfZ5VcAbyZA4XVxXONAeEuhm5ifNkQAijJQ6oSGaMPyEf+ULfcysP+
7n8evSpJlF0YkKu4Sw8uG+48vAE192I1yPN0M7gmFLb30in1ISSVrPhOLp4QQm6E
CrHZtYrgMfNzLw9URl8dw/dApQTL0wQ4FE+0LLaU+cg=
`protect END_PROTECTED
