`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47PPqZExuxJaDTY/srQl6jNy8XOjtIFBRVssL6amhH54
41skVB00MxgC99PEhxgW2/terHl6s79EXXCwsFXfWqj9iG3mwsLUalUEcSaHmOlr
XLdSsXxm0mOoS98nXV+/BPdtX7jMb8WGP4gLL56936ljOfu1zWe6flaztPyf7m/t
md3UgA1CKjrOxpZK+V4Zf3n/uJJAKoJBDeGtu5yawSE+FB+X9YeUXnD2GL3yqYdK
zCKITe8A6gXUSF39SkBKc81mp/biuK4vjXX8ckq9avJWvbAtfNpVWXRTnqKN+9W8
MWAB6gp51s3Va2kBpGXb9B44nvsMN7qitZIIB5Xz852AC0eZ8IsGGM0SF7z5QZU6
LYcPK/fOS5EiTfdMKZAJFw==
`protect END_PROTECTED
