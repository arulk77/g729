`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8Scl3LRJTdKM3ev+tzGyxZNiYGdWYqsAZlNtKT0uOv8H3
+edhnZRxEu28gAYw3NNU4YnQ4DVjykghBc+nNg8r/yH7Acps1d6W8HNLMPIp5dye
auXE+s03/40b7eebBWf8+51wHfBPQ5B89fdvdu/ks62O2GctZAay5P5loA0j8lHE
z6ix70r4YvzMfliU+913Kg==
`protect END_PROTECTED
