`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
o/gmXDD7Xixjnpr2OL/fpIO3zsruq5Ta1njTjGf7bGzLrAbQXs32VnogsB7t3kGH
R84GOeTQRvEnHEhhzDSRxJaJi5XJk0xdk2HBz98cf1473ov5K0R4WDq20ZQauBQA
ZTZn0tuSlwGJ35rUmPODpONklZjKLptEawJNMdQANqHY+jNEZAg5JrJv+a8QQk7q
rJ/qV/KiIP/e/sjUvhAPdnO7g+EO1HR8ddJRfQm0qsrDsYvt24hOIFRp/qhSkOMu
f6VSrVivXW+ww2XaQgy/v30xuXOQ8EgzlKnXnpYTWB4Fju1RWoXSeshlsNdykFeh
VNC0t5NWuhY0d/dKg9TYwdU7P5nLC2jN56ENOg+3v0g=
`protect END_PROTECTED
