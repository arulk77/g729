`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIDRY81ttYMZURku9qOmQZKrI8FtZ6kTebsmCMj+gKxE
jKB+dtWCushN5twW6z9tblkq9mqHSzxDvcGaeIrNDOV5ooxXKtkxjInSF+q0C0j2
wAHsxC8vXb/yjZGViQMWOcoAmYZv4BjF6ip/dybT+l0kJnaB4O9pGrWx7aXVPIIj
0OCSxvrINa7oY8TjJhynOQOT0Zd9KxKA2gArdF0ycjiPXxuFjY+HnbYFXCJ3DHvs
YNGb5MpDNOSa9i64wVurwQ==
`protect END_PROTECTED
