`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkWMKTOd+JIxGkt+cLzQl2XlC8qfXywZFO8pDLbt9mDgr
eBnBxW5MjbqH2hV5EOmT1LIZRfCVY16sWqwwax3PCgnZUGaRP/EYHYC3I06QcejW
6y/5A5XaCXm1GEsJf6GI+H+cCRa8MkzRDgbmtipLOv7QX6CVukwmQzX+FdAK0r6C
nR/yWkyyxvmiJ2fQFqRF09n95neQQHVCp38LzH5faemb1XY44kOqsiCPwaVzYhk6
O2jmpXfIye39lqUqXV2HIH4RkyLzfOCbEQt/Baajrbnuh+l6zGaBLgZZ58Dp+aJF
BLZmEG72OrgBzFnX7HOpji4IN+InLhRN/Xqvx9IdFXk=
`protect END_PROTECTED
