`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ2QNrVkq2dm2S9u7XVsKVAptbkZWcrMv9kaxQYyD4H/
Jdav+7Q83v2DiLDD84QFjgf6D8pixDT6r9fgpyc73x7ztdptKrt5coKOVWUV28BB
lp5k8Xz8vi60hziwNqPggx0HARuZEnYhqdsS3+GqEhvOBl78I31y0GtpGgmiWIe0
PI6cfP4KUemGkSIok9w+zk2f0h/D/lFivUAvn5ffPLWlkrz2g5uEhToWna4DjuyV
guRct583WW2fgrUNT8JQnEFskCDicZipnTaCpLbsmQBNTQnJpD242NO0Tp8iC0iC
6t1RXw7Asvfkx5wN304pxd8fJa4DJ7EhmUlEJfrv4xLr5BWCHTbsBnUQ4pamzl79
MEO0HgLdC93HrR+SmgljVLFf+Ybk49L/oJNUUfi3wU3z7TCmpqXzgMWpt04xjq4P
xCx3Ce2fqyXcCSrQETGuZVldRue8dR6TjH4pLWMsxJEXpzsZG+EfVmER2iuT1uf1
7IDoZg3hwJqXBtLXh3iFJAo1IEn4XgObLbOdHZH3Y+DqX8UANUkQoR4CmYyiAIRa
fhdA1yX2uFSqASQhz1wea16aCZPNqV3I6M+r6PM+ZWdEeTnNIWjGlYF6ahfFcOIH
I6FVipZqk7HOBhDfxscYcxy+oQtEzcpLFNN4UpoCfgnWZ6yI3atS4li6mYD+BMDw
eYFxkR/AqFAlwnOKWo28ybcfnoVrMld+pTzeMsv48FO1CfR4Ra10UiKqux6VfoZ1
zxFAehoPA/x/w2o52s/2siR661mMP5MWYF44ooja9RiCgmgxhaqsxSGITYB5fFEq
Gm05TZI8FnKzxBg4ik/cONtNyFeHgZ2xAGB63z8tLKI=
`protect END_PROTECTED
