`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDl922nfcESRSDVA4aBLkWfdyfkUDrCucyV+w+/eEV63
OVMVVhogxYsJzCx+ND6FH7vsYq1xFMJyW494JqDPqEQpPZX7XjBiAAa8fKBGFU3m
qpk9H/YnouZHT/pZ0xwHqL4ZunFPexTdsl0LxoTbfpb+cnWe3wFvH4kOZ4DTl8Vf
pZO21zbU8pxXfmwTr4Clknyh/UFD2p5XUVo0T+I5uZFXPUNwWRgngCiYcf/sQxyn
FXZBHZ/4zmtQS3yybVrn9GLifjeqorKJBAw5U7oDX92306fzi7hHJolEMwd7HwML
cVYhNvlUZa+oJW1/73r79w==
`protect END_PROTECTED
