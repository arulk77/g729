`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C8abnO6cGkEqNie7vPKoRf8VlUUyNwntgGxz8zrheryo
cni20TDK1BGKjdxb28DNw3cc+Z4MLdzS5LI3yRZoz2p3rZc8BkiHVsAgH4k2a4s7
jncNyKU0NGYWc9n7HHciYfa6y+evx6b73XdYQWfBAuHGYpGu/03AhYegfsO+iWQR
8HwGpyVktD8fqo3ywgP0DaSd2jTDFx6U2oOUbyi+m+8bdwhntkVHtrHoCRAy6DFH
Fyrp+/DZxyUaEjMhhr49kV2vFyf9zAeMUNIkPcem3DSPqQe3F93BV0mnTSMZ4Ja2
/Te/4EoLqrJa7VJWX93bCe+K1LllEvRbDCkLfcQM/oGLSl/lDMjnkiHuDt4cOILa
rQi3htKN4iiGL4SSKL9cOPYrKLGbsYIFWNBxIF4OuCv0n6hYtjC3xReU0e9S2UHz
mm0Q0UyRQaXnZgLNvOu/wo+80BwPCCkwzv/FKARcxpoUmoyLphSAG2zlHUSL7d0R
taExE4UpLWlNtKYrbgQmUWTden5goJNoFdE0zloBPYDb0wyOYl+U0pVZibNHQrsy
mjjjwjadi/UkBdTt3coIrhiUDbz7vL+cZ509w+vBbUIfeRbUvM7y+919GogGQbRx
2Gh3iGpD5JeCuZCHMClTZlLwWXTftaFFpaM1DnwJabpaV12Feiv4Rzo1T5sxjPEL
Sd2zZVTMzymDHqZUqnNVvcpG6ihyl9SleseOcVC+ZMwyKXX/CV8eVcfcsgRz0kad
b+wU1vWd9NAgP9lf0BmGeryJEXMU13Oxd1iwKIEFVD8oshNwsUUOUOWNidCchxcD
Gwc/7Yg9HJIz87fS5SdE2evl1ZAVK5uIocq44jMfXj9kmU2Z/0GL/ul3oWpCT5Nn
hjf682ZaeeamaGDbY0W5dpEYjTrxTJB/EjSZMdG2ZMjXgUjoP8z5ALVQCqDspX7N
NvZpiIdf/qmroiOMGkk6WVQyqTxC83NHT2kbbjDiCxvNaLZ1JCVHcdizv2Hr+ECO
SffHt7kzoh+pb2szjdjjU4dE0fHnz9DbS0/ElHlg2LbfkSsdEtFQekWw+9bJVq2D
mEZdRjcd1ELmMFjGiYA27uhWLhuxPP1ISeiC2jUaq8lIf//R19W9zDQb4o5beG60
ST4kqbhgd7lGZfD1eAr1dZgxOb0/f707Qx0mpgolHVbpHa191RLLx82tGv/Djiv4
/Ww6jrnDdQt8Pc2PMfmjauykghnKNa5bQkSJJW9DIglibciGzBFfd5OB87R+FwqP
BN7pHaKUzmtW/rMDuhfMoTHXz71vqQpRayIt8P2oWLaj+qUN83ZjWKnb7XiVeQRW
mVN35RViU+0aaDmZD904U39o9jIUuoqoeSRipdzVIVAjptdnyKQKndwsvIFs+sHk
KDOVZ9MnNFh0UJiOw9MQivzHbDZnrgr7sMNKiM4lgUph3/BCRLII1F5x+pWJh+Vm
rOpVhkyvyAjlgg1B+p0sD8gHC70aTnvEhEOonj+4Sy9qR+HbsjBYx0m9CtPNmHGp
jUyLdmJ75sCpGekp7XnWYNhDBkNQfhJc3V6UFu0RfOCFZkYuqKz1kg4HpmlJZtA2
E25ImyWbJ7xQsGPFbpwiH7i9xTgQWQiHpbkembeW8bpERsZzPX6R3FgBdoc1mkBQ
0WYP/Xr91io/vlOhHav5jnBqYYKpZfxOAoxITBnB8ccBal/9ereLsHShqm6e+W+n
EYFGmiB22/2prJ72VNDYQfbs+/OCbUtXGQZA9Vd6fD912PJ3eDW6h5eG2yzHH8aF
nJsdWMUA6T6JLeLv9iHPTf9x7RJRiudqzsWzoDeuYReVPO46kjU91ZY9+XcgaVAl
XCt20nszvWH7cjOCyko218xx6MPffy4+c55M2Bh3XKlrJhWANgVp5ch6+MfrI/wJ
pItaqNl7dvoBQtysrhCCmECfPmviSs//RUaoKsjqbdOrKZtGzZH141SrG7Oo4kz6
j3uxgrMbFfxSUOfZgywfLbYde2MsnHRNU/AjnXxWmI9Oh0sJ4UTVc3zo3LOjUOxr
WoYr3hHQH15rAgEMQFF8betmlv5Rquhe472888SR0WQmZbpur0e0jt2lN8e7qcx9
SoGQAs4yVZfPovkahe69tNzftaCApKjB7MxvmO24nnisgHOmbdGGgPPED/a+jBJY
QERPXRNKlWStSrkysy0iZVutbjrbmHUuT9KEAb7seW6GnBSq8gPg9jiLupZnQnzi
e9/Mza6Sk9Nq+p0+FqWYVedWvIwwUd8mAI0foHycfyCUbqNmESxcSZ6Prkyd2pqx
vyElj9vry76JNWRbCzvJ900mjMHuYC1euTRy6mx8cqR2bfTnpQLLcrnCHAk1hRq6
iALCcAzkTqChP7EyZ6THQsP+zlgKPzZdo8uMFjEz8/gb8vAu1uoYttyhbjA6d8w8
yId+YM5l7lXBHd+RljFoBh2qRR+wYPuo3lPrHDUKaP5norgPELZcfufAo0JnE44B
lakv1ogl5BKHp9GM+GBGVAjpOrabWdPXD7hv870ze5Se3c/+Rk7iOFi6hyhbsEIb
UUFnilsBA6oKRDtxulQLrbsBh36i3yKpWq9CIZYY21PUalyXpitNm8sySECsPAVk
WCJjngojw01etNcCsb4q03H4rz2ids2AgJksdmiSv7kPnlXtSz4XQ7i8+7MmWoIm
lFuvKLZZHyu4MqQhAkmEXWPsFevN75YXdyJcfwrm41l4zDqrsAg3j3CmQe+emqFf
FqcX/He5RWucOibfJ5nLNh35bRTx0YvKLmnNl10DIJ/gYy0qg8Vs/ovyCATctb+V
ltBeM1TjZfAc4kfT66/V+POr7moBOwuIMGq1b683L26qx/MLkv5DlJqHAzpMhR54
0LmbQeXNxUxKCClElc04py8fWLZMe2Yw694vmGs76XlNfwYSYWZ9J6dzAtLO5RMb
05SOyUwd22kB4cJ0ng0wUGobZhIN1I6wNxNHdrkxJb07zVPD20LuQR09URAbJeY7
IY8e/bHzjqaAzvXFcKpG53tV0JSCFlUZCuG/PInTEl1xMlMs1wjcRdxft1Y5THwp
`protect END_PROTECTED
