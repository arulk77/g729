`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
7I2w73FRJoVhn2QFRnasgp639uctA7yRaTwVFFae51esvNRvYnDGsSKcED6fz0Ks
ZKeaWnD1L+E/JMSmLdX0l7p0oxIbGg+nlehss/J+MG/qrUVlxu+522RmCuGkyB1Y
4VKerYfJH8hdeYih86qxv0++llWwR4o8LlkpR6XHsxOWg9n+K5fUh4D2WK7KZ+Pp
rZUWp/UWNfXW+Y7L7zZmIvjAKnIHStjC3D+nuIE0t9kvLadVOcj7oGKXzav0571B
Grc0bnvfDE7rl1ZUW/xbofL9oj/LOgCcmjOr05haoD8fwHN4S7I/KAI/eh+bGmCo
IVmW3OdHKvDiXgLr9d1HSRD7ywvwcjqz3Ar38uuBEZkE0n0MfGGSaTHpFtOyc1UV
IdN0edjS/DHBgrGpot/yTWntTEldT7dqi9K5yHpT1QE=
`protect END_PROTECTED
