`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/ELPyuJD6alYWa4ZhP3mMZR1jIz4Fism6GE7xI7lqzC
QmcdxviqRQf4FDwlqDWwLGl0Vq3tv7NLMlRXd45OtwZeaWx90JvOBQO8G4Ce0sg3
fcxNn628QPCybVOSE/Mcc2fAtLylZ3PojBRzBuqfg6ZhXLsMFscXFlmT+/bH1C5b
NhNyuSjfERRpx4l0qJANIqMaLihOrQjsZZqNvKV8XOkqzE2IAPD7MaqgbcbqZ8If
SWRZxNcyeD/BcrqKTkjKC5uBoILvt5IC4koWbX52gy4ZFfZhUrV2oKCxsPEorgqm
rDG0RSyVptzkBcNpriQj6w==
`protect END_PROTECTED
