`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2niYLszMe+KIskCEvZuwzhxOSOceLfbgPeBnOouVdh3xmjXgqQr/jxdLxSbLM6ct
Y0dtIJzNcQyiceoiRWB98Khp15cxu7YrOomXy0ul7SGwf+7r8MJ8CceJMiAG6ytl
jM25zflsr63BF86PqyqDDIrZWlEr0bJmt6z3FOVr4qwjVi9fkqmewMVyIhbCFoOx
fV/sZhGnE78iGF6HyoTVXIBJwWVKiZEncHCLqa8GPbq+HI1W0LWY36N5x85YUUcB
Sjsl0X7h8NeJq1S3CbML97sDGZapMr6Kf2XueeWyDvxn/uMfpMNrgdZRakdQkqfz
ejdLYx/xdRdrGoufnk5WWYJaW0Z1ihq3N4fYN2yKslNEfqMkDYEGU1yXh3uVGvtJ
cQ7xmQwFTDdalwe1Cv/OUZDbMmTG+Vg4I2gh3NpFEuQtSFQnN0ELnFYRq6j5VEbZ
8DvG/7SjdR1a5GoQhK/1plXI/sbDNB9AwFXRSQG4j6gzxkhM7rfK51AUCfKyOyzL
wGl2zYYyByKshdI3RCXBsr9OR/BLYfNOVafF6ghsSTC/0ja2dgF1nZUbAnpntFOW
cDEnbKeIUVrsl4a9vF9yKQ==
`protect END_PROTECTED
