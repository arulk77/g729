`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNrfcDZ/z24GKC1jCdGsUO+LHIXJS3pB3lPbE+JV1qXy
gbExNfKU2WtzOdfjsbrbIBIl4GtCTCAL1UKYZ4ENnpCNBPQItFtLKXDec12v8Axg
98V9OvhY5uzR/ow0kd9asCNW4qlC1RXK5s6N87oRhrxB+DIGG6JpVWEna7bOEF5Q
abCJ0AuBlQyYjNyFoDdkqQ==
`protect END_PROTECTED
