`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLONpqI7uv5hfhwYaz8TvKHXWeKr9enf76pVJBba4nHc
WqLTuopUfUxr+ckUIH+VBgxCgEkad5EOAmspW5NsyqA967F08LMi+50VLfJvl3a7
BICd1OYNhYgq7wyV5eJMQWUSXDfr/lpRrblaKhX5Z1PXvgdMubh5qHoM4LW3ztJA
KnuSPvYG5gTo/YomzFANcLEGOG5wz5CBXm57JL6QRZmBf1xS4L5vPyTzdjfj2Gzm
x+DDPAPOyZebZ42UYk+8L3n6+XJ3caXqojAhOj/TjyaQ0AXmIedhTCTUGeYNdOUo
KkusKekdRi6gBmURu8O7dYSKHXPD1LjASRr/63zofGftxTGA2numfJudpK3x7QTX
FByywQmUAupzICoqTe4pWzk9BgqUL7sf6wP9jUdxeDb2pnn34ZMO/Tu762sNZmtx
KSjzSfrXN0qYAgQ43UCfNdhgf3RWQpe+U23GdyRsx3wUmf4mZESKH+BBCZI0Za+t
e5Cmwc7pFlO8s7fvzRz31YcNYMUFC1Wn6XyMrzsP5iKIDTPnJBvk5DMXiim/MAk9
`protect END_PROTECTED
