`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
92tiggQQJggUlcv9SQy5B8AuzRoKmzBviyHT9dXZSFJr3WRbsp4Acewfi7sDXlBI
Qlzr0NwKPux4cEfMqcHtMygyhBENat2zVHQWOi8sFzvo54A//AWQXOOSzD5o8Lht
FFG7JQ04SeQWFGT2pCtLyACwwBhFQl8oCzaqAgKBiSVcvdiAGek1L2Wq+bIH5VaO
07dsTKbGd3VH9UMAhjMOQ/wioVFPeWQv2f3c3+yO2b80N7c3+eiSMJFzt+skGlqj
FEu88hEiJxhIxO++JZEKphrHL5t/H0l2PkHNbdtIILxIpP+7MRYhMCcx68oLilyi
js8so9tweOLtrr4sDVe55q1xeFWbbo7VSz51NCLX37gyT2q9WTZyWjX9b3AYm5Be
zKXhS9OGVhnSgBMy3d8fk6sWkruX05FbDLf8deQxivVsj0GrezxBG2Fnkno0L9my
g4248dWxXcH/nOja9yHW60p2Y1JgQoa/C+dCvEZjYyAdDw+lPZMtO4wkyNc5MbXi
XizXOA5EeOrwFkrji9+qHzkhHjuwviOkEsVmyJKVC25ZWDz/FCikfDB6JPvZJGGX
HZ6VCzlCR2aZOC/OdrN93sJWnrrbclT8HmR4gdvvFQQRtzxTNTTh7VjmtILjhfU+
cxe9366rEw4K4J9sdjDtU/4E5gkGyqWRWKkYouTk0DfFCGAi2XzpWFCzIOPVWmwB
l00kQDPRHgnsGQEjtqSMiZqwX8Y8LQnf5s0eEsKRKoXB7Mn8TJAjB3ixvpY6gZH7
QL77sTPSC4223FQ4oW86Gv80LgnMGxwBJxYScah6py0IfWa/5o5R6hpji62vvZHS
qZhR8LaeyOKjxe0G5QKuawvrMVLI9zScbysBHEQhHrojRPN2QBPCL6ZkaHAsikuV
OyM62jI6kpLNrLMoir7qHJ5S5E3cmIJr0EizmA1deUbb+RayhKARGSAlgq/q8sTf
xGP4wVdSdolfgqyxfxwppQ/2cRtV0DzL68E1zyIziqh2gzo2mZQFIoGxS9ln34e/
BGOoTMSFNz2yyb4oDWkWDNeNnfAfuNx8q/yL34Rf8CIBTMp25QXvbUe2Odlnekgh
Q4pUyTXhZfFRAsq/ls5SCccwD16U8uJjUU/72i9BK61fo6oAX+TdxQAvlaVTO632
PCw3fzQg+oq/irvgFJ37iGa6jhocvT/5+DVl1bARJFg=
`protect END_PROTECTED
