`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SWwtd05sOLA654/h98hOj9CZlqJs1X18pteiq+G+Y0Kt
4FvpN1rkYIiGL7rWRj4YcPkcxf8jPjyEKuUpMdIosl2E82kYG6odufiaGi2PrS/r
TKbFB49RDCiLfz1B8/FjOzAgm72GB4hMBhr9RJgcZGpigV8JaBUYaoWBV2vDvnNt
FT6rVuc9XwIbN+Jxwkl2E7vc9KDe+Z2B0aUu/RJjA0aQTuPv5mEc/xkeLvCf45N6
5P9GT2G3IRl8OGxJ7zn+aiYwto1JQYXhKuyMou9pBU6DV+81hs6L32BShEKCJXnB
b4qN4xr/MAkOXNgm7KZjqYjy+w80StSOQovki/3MdMGGJz7rEGzEEaI6XzLsjuxc
FTVxyfJZIAq1tTxcxFfZWqQfyb0wsOtvCa0llWYZ4c7r4ao3/d9x7hSBUKfAgxXq
PAiNzMivEgI+0+b3h5Kp/IyZEore3xNebth/sKc0Cs98pMfBY++W2FBPvQntvk7P
tIaEv1+ckbT4eh1k26AmG38PlffIaqq19M+Tg25vk3QhuH1JXYooYwPZiIhW/w4F
kKBOk7mOqsRxoxb6XtXgB4zFBkSQENisoH8PP0/t622bvkthzZK531hVOryBkvWr
0p5vQDVFCnLHMmN9R8n5/HtaL+98iy38NAZCVRMEcJRdvHReTh5kENL8tGA9eMg2
6YKQJPT6TvIJKheGwwVgSGhaGV+ngEk1GfmIf+1QuJzj4I/oOyer4rslfRW9fTeG
/K2g80GzOB8TB/h1hOpNfIjqiZ9EwEnPNITkdHcuyUXOishjgQ35Wn1uRSHcCVZC
fH9c8hzmzK7LFyoQlVbYPaRxKKkb2h14KlMmpKzUhDZWJ7ZIofxwWBZ9zVtC1brU
j/pcic+elE3QHzOR5Y5k/TgMz9hMAiqVIofDvBF8TIWaJLHspeoHIt/sGpw6icDV
PqPj2EDQUogq8+TWGMIM3gh0m5MZXcFddKGU61qWRHyOorDYEIOa+hSb1w6Lz6YX
+isF2rLa8pkt2ZtLJK+F1ewFris0b3C+MRIT87lqNvbQOUrQyWnizMz0JmZziRi1
Ohq2ztvcrxtP9nRuzy4S3srPL1UvbYjsb9c6/95EUTn9WvH3QIcolCeDmi6yzQBh
A3nTyacGmn5glsuW9rr42cdLF65mvj+l7c2HB37N06ZtrR2IgNnlT2vC2P/EgAKk
AQ8rnKT8Y5QDzc+f7smr9waCz1cnrXtLm3kPEIshZba90CjxY/GynRhCqVg120uX
ns4z15OfbRuc8SFQQq+dCR96USN0pBb0GZ+Yn0SM4XvAK/x3wLThRI5+13BBeIKK
XXdPBV3MBXH1eljoIg3ayuVhdBuGc4X0Oxii1ABJCvfciBQkoIKYuZFsIm1YkBMJ
fszubkFou6O4jm7C8RLKCv9u+uZbCqtRqgC/klBfOHHu5QToGar3+RwsolMYOwtn
07FFLfn1QoBXVPQiDKJdPF/4KzRc7LjTr99o4vVdl1twRr7lqP7XTp3n4mNLFOP9
dNxsNbXtbtOwak2GkJklHim54KhwmmFrOlFrDTI2Dy2zcIpmesIKqwOTy3Ye4IN1
uxHqBgf8PdboEMvKPe2N1q7bFjaNOFn34OSQuq20bn4+i+22jELGHi33v/BZe7VM
ZPppIKIeenkaPIp30++WSBht7k4cCgoSSLhDG8scHIBjNPl6IqF/+2LLYCwOx6gA
nKDAkYi3wul7RJS1SHWR4DoE9NxZrvTIJJTlWhEHkkes8C+nsMrHWLPZTMaD/7Gq
mHUPELXg2mZtRuXK7YOwyXmnwWf6/hECKU/29w7UJtADVlk7YHyiJ9cKLcmGVM6L
jrhZV/2LbCbffNVDU0pCtu+YhR4TygD8yqGmX7pqvTxky512ZWCmGMOiKsOS7wD2
jcnRENv3Mw5Ua4WHADN6wmOg+tTEKAOEJ30gl3SkRz+BFOHx/cG5AB+Wi4ckxSHE
ZZ/OnW4fROYo0f0vvcYIAx8evYKka+hiTLki3uctplUiWWKft/QRQ8QvVB+Y9Nb9
TW6/kMFoFfH1/PLgqjraV4O/Cjt4rwpH3ITxlN2kHnaPbyJxyx/jnus7Sweb97Xa
NzpRoEjduZKRgsyIzMry+1y+EZX5vt1KI1ZZJ37BNY5JEQO1ACcVfvFSYrHUnFib
W0Qfmu+5o0Te6eA8YFDFaZFGZfQL0RcqDSbN/lF0acAhg6GzpXTN5hXghfIKyqwZ
WJFaTu3JY4sp4DXbKnS++eZMS7eO6sIgXxe0pL3PosOfLb3376WNJtGpb17BqYV4
E+h+u0RGpkPZkxdJG7mFmQ==
`protect END_PROTECTED
