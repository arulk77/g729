`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
m0HxSBTcMrv7Jg7XTCLIdPRgETwXGD4wOORL+iqccMDLPehi84+20JdOSj//mFx9
Z2ydwPMWScwyXJ2xSiS8+K2ZXY051uWW1N2DjZaCwiwepSjY3XFc6m+8bKMrhZ/d
ABnu4y+QMafxbwbKqikw5iB/3AXgPzccRSFk9Ex81F+hMgLaw6QM4L9W3gzHO0SW
Fq+Wip+qd2hzGZJWMicAninc2FpWDMfpv99KV7M6TUOs3u2YLLTW6ZSP9gZzY1P6
dWI4csuXOBJfiFXknQd/UTUM+KtwhtONDo1x0p6DBz31BvH4WS+SRk/nTCybwjN9
5czAkriGKI1YfW1sYaBeCb+pET3otnJiIzyJXGlGqGJSMca5pCmvVgMrDLkna/rA
XuJS7DqhO2CHZqG/pEkt5eFbFhgWzBT5MGI0XX8yRY1P2wi8/FHT8RCXKweAQtww
tLDHRPo9BxUatKtjVhWWYQT8xGEiOcMGgeLgNIMV9uC0PBxt+91hl3vTexYuyCCX
5KHrYljOfcUMnxDHPy5+ri3l+Y2Jg0GBx21IJvHXLuSLSONl6Z7rJyhpp/XZbMNi
FRltJ3ZDKtkl+TIA2cg/IOcA4PMnbuILAuFcGStXkRpqsUyHRlw57YBoyCQDVcBM
rIJpXdt+VkD8cZ1HNa7gcmMCYKFwt4NE6/XKS7xDpmvTpbw2cCO2qki54ANPxahI
fULL8VzgWOGLz4vg6+L1HxkmuOKNvc7y5Mpgh0jGyEQxlX1V1xvN3DoyHH3Yk0yC
61rQDJTjKz5NzSRm9iXjvgvHGVDt3EJRVF2A0wEK1QZjJ9LiWs7QN4DfJ5LA//05
/j3iqnoT8n9i2Gz3uiq8xU6Kc0SPfFpcRZfY5nIMnyyKJ3qImt4Hvyd8DAgRvN5c
uo8xeW2W+sk/Qb6Nro1wrD1f2UNCOAF+kwlposGaZ8ccj5xNoBsfFLDWScksjEsp
ZS5uV3Nf0jKbJ2EHvmMMkLQ9jxSSB4ogbekrBVxRMp8739aexu3Hpx9iC1gky1Jc
XvvVTiv3LHL/QYyBsmb0Rl92JzV1fmrb1PWOL2LYpQ5eDTdDf9T6MQDqbpuigvuy
ZzuzO2vbrzqXH27+u9xRlLiUgLbIz1Giqvkfj/w6221lBMxl7N7rwHFL9v7JHj3+
OG6hSBGy8H2RjxQ0rpGJQ7/KM5dHvU179HIlDQwKQ1v4PcbLhVMqKNzEA/S2g3OS
NGA+5cgPNYyUvnaObc78oJv9g+eo5yZNgYrcLMqttQ81NKHixTZp9w2HCnjysilp
mBfBrqmEjoLoaPlgTsFF0sGTj59IpMOCoB9ZL8UhyRcZ1K+WkOsX7BpPKGsjK7Xs
TjAAtf189yY5PZtYR4sKj5I9+MXUmJmPHVZ/2Zww55NQJGJfOOwvjfQCHzpAybm0
Bqy66sRz0HRjq4lwma/WM39F36uOmkF0iwn23rOAagNErJ6wspXENeljtY5VztHS
Q4X0Rfd5y6rnsOpPjMnKTrskahgZ73XiVkCnaMcPXNTnkg3b6gQILnPg84F/gjbA
+tTLyhRHnOkPsdT98YBqJy05FGXiwEpYMrnaHetmNDdCPESQzhqKN62ECpbOPdga
uJyOpEToZev/JyRpQazl1kzXwREhbt8nB9flz+7lh9zYOCLoH70Tal2YLNXJ2fow
45WOj1nsnTKTRvQZvOTU8Mq1Be2E1/QVayTOR/KIK3MqxkqWx1lalnIHXOtW7bhn
qBg+frChQbWb+rje9cGY3tMJUJEJPEu3ouCMlYkJobVl5sXNPTOl++KOrhf5Qxz0
zgCfZ2ECta+0ptr7pjRAvT/jn0xaUDPVyXHGK2NO0Njd1EEdn5eFC8SRPnxBlPrU
A6GeYW0bM9dXLoi2bg5DVhKSkOIqQ/aB4iZ99fGeS4xuS8XQIsoaL8eCfjRsEOXk
CVfn5wzv8S7RtENQT6cWD7Uht5bIRX7GLLg4XgmtLXkvLjJ8674i/VSJW7t6c7/m
m1NMwyorXTjbvbysh4AXLw==
`protect END_PROTECTED
