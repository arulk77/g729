`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEUpBobEyooRDb4z0MKQOuCYa6wRaf/s8O8vROM1FNPm
WWiVNARBb5F49v2rkjkyjCynOzZxLSzZ6n2emUma2VLaNxTS4Nj0nInCTqvsSPdZ
Z+9xPeMyblGIth0hlz4peuwEUBXTmBgV99k4JLXuyoA8MI/j89/jd4VE9+Z7W/QX
wA+KDU4+XqOOwadrAfbALcaOIg5c81pR2DLUwJiXuDRdlcGMivuYWYRrkpwiyH8n
qyHrg7UruD77Q31jIgjNsOUN28hN9p74xiwkZZi4HQrWMT7iGTXD2iHcDJk+v9jI
hidzfThops+utz7YTD3fjbIrTbbvJR2aRfkep8k0udma15NDQRxt5j+Owu09lfsB
sicaz9R1lFrRQauQhq/Y1IsjGWH62krrabEiKsjmr1sKSIhrQge+bF/GDuienM9c
Y8YsLv7+4Y9t01I4VQImeKMKhHXF0k/p0VGGvoaEeO/WLAWImLquFSFBH3saeHIO
mX8N0Hp55wqthHq6M9XT7oCdUVMn8zW7KVdSMPa7w9/gEZXbFULsxU/f4qpnDfNh
`protect END_PROTECTED
