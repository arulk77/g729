`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEgzHXZK40WDzlnTH2J1jQ1QeUPKKeX7KQ5Iv8cPoM+H
03N82aoKoPN4n0fflU7XYLVkfXuYNQrRp++Osk876f2Ny0xwz1Fteza3Z6GjEsz0
wTWIGgdyoycXchja/UMwoiXUYXBAZDs8lzSDSVvOn1JgDTWtkBMdbB8e6vdYN2ls
zl8o06tHPmqhBJzHXst26OH8RD7VNAVV0k3Fq9CKGU7dkzWYBP17oAwxINsgbtfg
nAyo0zHM7Qogu6RcCoUIJTz8/CxqU502iTKh48UQkEV6rItD/pvM4fzhXcPINbF6
WilKUXfd4pqtr1qQK2e56C+2f+dYCjjsMIV6pjHSo8QLh4domju3hRdlGrfg55bC
24Yij0zpQhFCdPAz37uuG/rDcrFrsWJZVemqtt91aHv1Fyim38oCZ/aslnSuVvsj
PfaeDbcJ99MkSI9PkJNBzVQzBftPN/95dQOPLi1yMv9UUZqapJYhBIR54reAxuhR
YPgGJmbFb96cFMXK3qnD/Zqu7m4EIc8vQk9Y0XOLn/p0WlQeHzGL5gL9QpD5F1vF
dtSXYl4CxWo7iOXTcUlYYhUh/m3GKHWnmVKcuCc0CEyozvuK6POcyvEG7kXEZsl+
QQ1RZ4uiexII4EqPssUmrnTr5ZzrOP3E+5yG/1Hb76VmDuJqSJ0KVfblXsYAAo+w
+svk6CxCR8fbiANhWO6b7BizsqNeomCEi38RmA3evbjXJYJvhFlNWBMYhTdfl3gz
9DvKp0HZxnsovfdyPWxCPiZxZ0XIZErqDuVEHa0fkKJuYxyqcKeWgL5fspMLYsT+
P6zS2/XQvRRep4ppjZGdEK0PxQSx1w1F3Vso+aUISGNsP3qcXDdlVpHCp4FzJVME
PDTQ9SpDnxN4LEWsw+AJDc9oEmpaoBrf/2sZ5YL/cNXaa/yYaN3BAOOLrLdG9uJZ
x0H1VB0sFR45/UM1WhsghZbd3FJgHYP0CiQ79mTpeK3QgVHFKVU2l9A/OYXb1Plg
4zo9nQ+alSc9xdT2gpUZKjG2chbSKQSd9FvL0EzEP9NYoRqYY5/wVGjBeRy8eM+R
UfpAWmSHzZxrezVoKcdiGgf3/W8W7eDlFD7pa1KAxE95WCdU4NDOfdvc52VzT3Vw
JL28eBLJhv5V2MfEG4SXtCkD+zTOnL6zM62jXAdiBJAeSZm9XTSTfnWSsXMXb41A
OCGDhx5f8Lwk32sVdRiD7gr0i6O/Nreoqx6muQ4Cq0qcVB7CyiljAx9pnb/V5Twb
oix9IH24L8tVSJN94gnjDn4YpFENQHrQibC3bEomt9DUDOtEjINPZlpDWs/qyNPi
SOcDS7HFhXaSPxrIp4scp1GSpgMnJEppJ0zEAhsaFZyVZm/b029aiw3sd++8Kv0C
aZX6QZ4+n6m53yNx+gun4YIGB710DODfr0yabTOaEkVADgxY9aKjhjeMeOik+gDl
OWKAR1rh649+mQ3s7iDsbEI+d3EIWewU56mj+TxKYzzcG2G0Z1lqyzcHYZ4xQ572
NgbIDJNyL/3vSDDbTDXSAd423iXsIBN42ARdCw8fFhMtgX5TWyq2Sn07hEtob4G7
DGEbqRlr4S5vlz/g5CJ/dWpZY3Sd63JYUzXW3eFwg5Qvd+uL8N6jCcTdRW3Npdd2
n2xiVGGBtq3xs3CN2K1XJ79Y4BjR+crS1GFwQynuu8fH637Ky6JtEap0HgelODof
BKvfF7fk+scPn0omHY7qyGnuSDK5zyVYBZqqR12lPLgxEnbAH/ox27WQ5axp5qZk
kAcZnNiQ4EthWEJo9hHQk97XmBx65qwJ1lKz1nFw27/aMUcQA4ApdCs/XiOfaYav
ClRK0Vre9CPrPeda8naMe1bTiLQUwjU2qx5qWAl9tPdWpxpk3+dUyJLbItWzVZoq
2pE8GVDCaX8FzHpNJKChji1V7eSzflmxx6z3S6TiJq1caGj1pfnQ3x7X6eXIpfkt
+1GRIMz+ZUTdfwMgfHsiszjAMgCMyL2uDnWArqg6zfACCeqBVOAMRN62HTs64tVq
zZa5Jkm9nEze4AwUvZfWPI20Ff19FoYGRO5sqrQDc1CGniusmOSY90rBWOAwtl+r
ManXpDA/sDEvKBqUw2xJwsVFs1ywrqeLMOmqRpCnov88A8DtZqwcSBNXH5c/WRKu
7+s/hvwg5D69rItumYMGmcWMyGOoHB3kusfuThvG3jBfPAy2O2Nr4e6C6mqnZRlS
pdXkLR11A0qQhjIEqelPqW3E3/1W28ZIwPK7VRiDbCNfTiAwoyv+7uPZR84hXZ8T
uznmQKEvTMmgeGj0FM7C8f7CTbOdqlVCBdqALrbBW8uGJojNM507wyol6P9LHp1C
OBX+0Fn2Xe4ktVIovdZmrwwhw7Npt51FPdaJ6ttFIa5w0lqaIMqwUweTqzAk1nwA
oSEzx41UIfi2A3f/hD7LyPUGTfZgKMvwyDeTliecyZ5iJ02noT99JNCz/+fTUQUb
P3Fhs/EsSeixWKbSzHKVUIGRlPDKaFhuyYX6whj3zGvSgLOIWXmvfbqoVtRSHDXo
9M74sfXlYxsWuQBt59yEI3VtFoSiKjDOBBBJqjLaBukwfFI4OwGW09flCtzfikQl
JhS0niv57Pi3fd8Xu0Vzx0mWIvxy+OUjapc7s3lNNXj/W/0RbRLvT6A+ps+p0mpf
2ovP1Ugf+WKU6kwXzjvtiv8dWOmttyofx6QxjOxPysTxuh2ohYbikL8s9wAuvLLS
0X90UQat7WX/O0kxrLmic0nkO1kleYK9Eq1zR436kyPLqqDW8iII1xxyKZy4s7uO
OILjgzOFJ0fW8e3RoqzW7xXUGrCPNJcbuwXS0bu0Am55pXKsxoORknhboOBpn/KM
DUWdkRVHqiQ2qFLTILrTUgRnJInKXQeQtaVOARLeOd/J3KhyFnkpNJUg2PVXnSDh
YicyvMzhITbQ/ii8x+uh4Ywb/IrBsRU+VIWNErAJl043XormeZ6wedrjtU2TnxyF
14WfUqlSby8JB/3U3OFBsbinIc+AY0KoUezEptU13VRj3v3x3VpX06t8hH9UGAxR
pv/uFpdpP0kydc/rvsq6WX1VF6uO1PXbOXjca2x3Lu/1oT11ApoVTukNtukBQcSl
9YUV8KkYgblPMGSupDDqZIBjDHZjqSIE2++cYu3buBvqQxcA/jVIX80iI8qhzIlY
emcQEH48zST6itJsAZEWOqp14HB89JeQJQw7mDhhWwPGYbR6lcwvYD/Op/JAbcb7
gbwCh/vxu2fcO5pKnOjv589kbyiwwHBJpuOBvVLUgqw7wZKCSOPGtOxHXHSH+fc4
zCxiyaHPSN1OknFrN+uUe/E3Zbo64PmRMtT7JmEyJbbaHeQU2TbtI/j1hevVe+37
427etJVhW2gVvJqfZPhzubeVflyAdmgy0vaxDBZXcvfTksCMJU48ZDihFMMuadyI
67zlWBCUDW3raFtIAnNukklT8AFrV9y1bqXgaQKtKie5tLtDj1gSB1Vqebz0JGtN
8uPGpHMK7lLs69IhhRYuRu8aq5sHo8T7srieMGTYcA4=
`protect END_PROTECTED
