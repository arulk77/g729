`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDigDUG6QxXiV/Q9Kre3r5cl0zdepHHk+tpS2UQGRYYO
R1hyvxGDrvTEKinO6mj2grXrBCvfJNcGf33WjyaqvwkxopjgURLe99lfpeHOzLdy
dUzUAzeQac0m3UmMPYCRex5NkOqfR8h4IExnPc6re5qJxXUrt7c37fKCyl+C4GJh
GdP5gfb6uPN83XY8lYWKPnCdBptrLgkNGDZF5r5nlEPcOpeoNVdgW/T85f37xVJd
`protect END_PROTECTED
