`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
J0WDZSprj3/CqrYAEfVPMfAB4Hj8VwS+PTW4fjRjVneKIOqH+QYjkyR+KLhiQZ0L
sA4zk/o8zE9RmQWWRKk6rqlR9X2fr68cGeEVWgjiEaL1TFDzb/ywfywvMhpV5OTU
WoW9D7y/cw9wjnwe5iHZbfwDIGQdIS4crC/BJJGUiakag/s6ZZDBC6iHNfOYZv1S
1FWyQW8hi922REst+xf1MNyWLbCeOABh37T/QpDNSM0=
`protect END_PROTECTED
