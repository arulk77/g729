`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHQFaEA28dIFoqUWkIwZMJ1saSiWM4vsgnjMuUoeo+bS
532Pnb1HJGjbho9snQ6eKCrdQUxDfYu+r5fu7voeWa1I8KgawHnwp0Ttvy5Mhw3U
QZPoUW4gL0NkPGUk0hD5Zq5aCczPxbaS1Nd8oH1egMMEUl4hXT0dqfqwYFt1m3KK
qWjip6pe+BiM4A9ySkoV8nvwbQbiExEanldoKARbA3qzMd/dbjDmr/7+msYgDjFM
5dPM/GMn/xIE1WeZiovLWhLxJij58R/ENGhD1LLtZXy0YGlcg+2Szm0JrLABQPJ9
dxiq8roE0mHa3CRPl3h/nsajROYvf+YR+NDHE141nCX95F7Lk+qaArZ37rCyfB3F
6cwa4cHDiX6rUPjlJ2TCASY6z4TDYPoVKhPsznQeAdE2H8vD+wB8/rhDOYhGNCkr
o/cnJCtfx0qGv3lBHDOUZmMe+B++6YRjn8KGVRcUxit5oayCk0Hb6Ce7z9dYbiMb
L7j41hKD8VLqe96KpDO88aUq2wTC6sRpmvkLf2y8kNaWkL2u8zaNC/aWJnRqKtBr
7kDYijL0HXHQsfcOjUb2o8d5rhvi8ZPtLzcbGkHgZBys/SG0BJ4xMOpdbpJ2kf0O
B9C75ow6z3wBrzFrw+K465194GuEWbzWl+g9Pnw7+MOZJsYWvigMoeYX84l8EC2C
BA/Zh5/6MAY2UOhvrMXO0GDb8zxvbQ0JaUpFlzynde4uZ9U7ovpohsZZRs2mV4t7
ilSAJgiN3zJLMgVDqWWAGeikxol+4lirRf2jYD4ckcN9hTtPWLYktZV/yvFM6axU
UB8OCNRaGxYKrE6f/lNHcgSfRMXeCfN6iOPIv2GHcAovANHl0jwzs2jM1QJkNKHf
YGEzlEJHdBaq2mWF70Sx43oKDM20h8Pgd+NmzgvFx/m+YFY2hYrBO7WnJsfEhseT
jvm+NEycqJ+2hDFWYmEegjlswI1wEzljmGuuN5e0Zwd/XQrfB2FB1Td31Gri7zVm
PX/Goz0rwZY3nsDzmEQrvcCOkOChHq6my+OgIzCSstqkLcPKg907+W4wTsk+tKRw
hiDcEkb0Jjc4Noy6SwOeuD0UEnlBSvZ99VyBrdTcyVFXxTmcm06HZnklvubICUd+
YsNQG3vSxbXyrwU29DJbCVHTuIkvKr9IVZ5S7NE8rQEqZeTmdvkjpa1juxkR3csk
YFAtReqYOwDt9VhgqnhNXFO0jDp1idhlYLVn+Tj2MrlwRx66jRGvMoR5EARZthH+
ioMeXGdxL3b1wMmKYjb4S4oVoAuHhDZZhGJY6tKxoFpgBgpRfLzBRuvpVq9uMCMz
ICPoLuM00mPfWXjHYNNE5W3T0pswht//GQp+mxsfM52mMM44mLHxtYu4tu2aLC38
LiZcTOAu8ck7SqvN4rAQHLD6ByqfruOYNcIUu+AORPvZdmOQ5tkheIP6fY2NUp+c
3AkdN6d/Orkd3pJA43e72rKdnQoIQV9/cp10dzB90I9LHKjxdTxysRIVhlVUGo/A
D8+4ZO5DAGGEfS5r4593MLLNSsOSkabwIXAg5whQqbqJoLXGmHpQEdm5Xonn+XTx
tnCsaSX6AG1I7PFr6RBaqnJ1cadvbl1SLI9l+3EYB6crWusQv4eBeO8eC8MuUbSw
nA3BkBVrZCdUtSgs9RzGOw==
`protect END_PROTECTED
