`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
wPIHdWMoq4uhQ6ksjQ+UEQTf5Dda4hsLJFereSEGOpXea7TUrUd5CZPKOne39lia
j7F2E/PHtpjPSDkaHUy9jpT+G9zaBijCr2UEemfr7IFSscAyVX48Ta72mPM/+zIg
GglM0VKcHRdFmh1L4zja4q9Vk72DdtGV0MR9xD/TmTKoV9JuULDd7v0iQmrGMlef
ZHRli3pgx2hncMgvgEBUryD6z2WODLr42n7l3OpqoTuaxO5KS/qM9/sEjOcr7abJ
70Ych46BXny7lkGJ9acGBayQJlQ2onPr81gtzCDQ+9MUxlc244D+R9iJBmBny/4P
iD0GPnbS558joohIyp6dUxzxCMo9V4niFmARmrg+88Iw3eBn9ACghFrmbR0gAqHN
rcLJJhRVWu1LguBytU0wqBh6SI9/QcqLuOO2l72ktHTiG875cPslwi8qzjkmjDPY
JR7mx7LCBqiyg74wlZ0n75tdvugLXIl5JbmFeYqQpEnLZvIKmTPzx+sAK10hrGwq
LNYe1GtgE+SJBuDWT6K03AFLRmv6tZe5xpBDyHtZlvFpdTPwdV0rgYTAdm/lvALc
bdNb9XvCOuncE/lp6pVYVQ==
`protect END_PROTECTED
