`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveISskmXPYF9e+RJU+xBFAL2BTLSh/4I9705HiVX7QTVX
bsr4eK4O9BPaL3bdbFtgypcYFcTyhuwdiB545grNZxW8+Zhh+nxiLykwL2ei0gPA
pGBOveNTD81PVkAphuKNr16EP2geFdv2g5Iv6n9+jvwbWd6M+SjgdeFyDEWOWVwC
NbuxJdnYFjowHNeBs2mjKu6YFK5PZlxEjVye3BhIdrq2L7LHbn0hrIeVX+UsjZWJ
B1MFLQ7EiJ/xEx8ele+K69UtdJKyrpjpVIW6Ycr8mAkZxUze82Y8KTv09XksnOxa
Aj1AFm4gBcGvJ++WOLRlxMKu4ENAo2k16opdyIgnoN17/HfqNwG+uWDkAYkBnglp
yFLdjRX8oZSVuuZ6PnVp6xrYJ8/Ru1sUSPZfun37JbRPAhD6dinLkHojf5Jn42eY
z8rWqEyD0Dx2GAhCoCRqMeLf6RUWDQ2o5qn+aVRrMmk9aYdyQAsA+hv97qKy+5GR
`protect END_PROTECTED
