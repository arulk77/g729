`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCZu2W91JGJm6svvmF1LoIjb7K3qz/HZ5Fy5C4Enywmi
H+GHhK77q70cFPirDda1lKFWchu1f+YSpKSHZJXe3IYm9uaGQkJQAJAPQcCjoXyb
MZ1X4/UrR8ME0Xu2RRjrziQ5IcpG5V/POEASJuYnpW+rR5Qm963wSbo3XLo+cJD7
ihUjenLj3+TfXjDMUui+2oqmey6FHk6ztgL/sQHwi39kvpWGcWa13RXm887p9LWn
YDuDdi+cX0rjKuJ1MF2l4a1LidqlD8AVkf2L/riz0QIis6zEX/gVzcZo450swnGu
F3Zu+OiMxKrovWdhPBhyueBFDLuU+tpwZwdj1NBKcIfA8Qq3VNNUR7y5+iACRu5j
DMJRl0Lc5xodi3zQNNJF1O1G0xSFgKnCFhXQp7lTIE57Kw1j0q2um8WeMVApChRf
LgEJT8nw1fZx8jxwmQEAOBMHf8b6weE6UG4sbNuuEOFBkXXK0a440Rme5SjxjOQa
sIR6gOKdGKyy0ozHWtsaG849bqF32WDKfz1a9QiK/ab/s6UsUxAZbkb5ugulPk1P
EdrDjQW7KX/I77oM5Rl+fq4eFnrE9jcA+XHRt1alQryBdBED2XmVU4DUaDa5v9qM
HVIEeRn6s56YM6COvKuxc7UDetlUEWAG0JHjwweNKlZ2eFryUFPyqa4RjOFmL2Ds
4kpxf27AprQ1LRfXrIC5mIqe7wBFodCKt9KFvmsfYKm8msyTDi69hQNTip/jXjOh
M+V/pqf7GtnczvqxCAkslFe3wQ6G8b9IwXoGLQaMaCEipaL7xuBvC1hneZx/52iD
c0J9p5/E3GL+1FqLosiQMrUzikEAFG4jG7Fi2POx7As=
`protect END_PROTECTED
