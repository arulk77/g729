`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2RtTiaLwZbJSuPbraFO4dpTn/cz2Ty+EuESUabcZD48EDuQf61wzqIfu3xC7fDM0
XM674yO6dVEl6n9F0kqTLCMszoE1JRUSnAg+6VGElQZTifIuVccH+PKoCt3a2kKR
8HlgUobjVe6qjZe999PJHqDqcH1/qUFcrL4UIfdqNUw40PONcFy0TVpErVky5TUa
`protect END_PROTECTED
