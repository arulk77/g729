`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4733sYi5EwsXQP+Mc9SlBmfL8v5T89lzSWdiab51p9in
wVaHscYwurS69aeoJDRN8b8SJZo/DK5G1CVTx5pRXaf1dJroZf3Mm2kjC0gYMu4h
2SXvdOIgIuXXWN+VxXpT3HqSR8HCDa3qjlj37KEtzWN6dlk0EYF6LfVAUJoZhBlu
XSx9AIou1LAQLQyf2ReNdI2UFb3kIwm2Cen7z9DRg9alZKWt889XHKxvLsU918+e
EkCqjjUbxmj3zgQjqA0cCu0RgshuSxog3IL7h9DMkzK5Qhtyn1frI3ig7iKKE9cd
MhpvgbEy/Yq9D2FVTI3lRw==
`protect END_PROTECTED
