`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHUSDbv0MjEPd/Kl37NLGYz8jws+EzAPZkqroqBgM9ND
/0VGlUi9iXnJSEiCy+7cMCNOtEBnlL0opurKrCBlW33RGCwIOnproGHzwwYnqxz3
P8UFevlgavWHYwS91muMVhNa7RIHq5iySi+s3nzN9f1N2wZubCzuMvriwR/y3OkW
redu3C3MGfs3vPxgO7Y9cegdJBMS9SLNvDVd5BVYY8ycMJP/bovwMbaoESo35meM
fy3fjtF7L8a9sQk83fMw+DwaQyjdoZI6SuTnlRQtEh3JEQRQ15zG93xvLsBPD8b6
p2npeZfKoeyeUt6fU1mAvxunzEbQZ6o6GXgUfjmtBscLRtoSdub+3LkuI+VPORd9
ZBTpmVZJTuK6BdRgeoD7+4DN3SxmIIQdRt0943/ai00fsBfjCPK0HNNo6W+8RPL9
SH04kZVcDfF769j8nEjaAu6111C0WK9I/yQJeIvcn+Q9KJEuPdaAOWhXO54rkx7a
7PjNBsbH6cuuavbJM0uiX9qOF/uqgNbXU0dUk7MXvrINIH7djTaE+ReFXghbbL/1
`protect END_PROTECTED
