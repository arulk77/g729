`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48jD9YeRtezd/M2tv7rDq2W3sTtNnIBqBv/74OCg+TYy
6CEKxEwQW/ZPRYfkJcwzYipdtqzw5Mk4bO0+7E9nRaa+hOyVvTX1XlkHYpFwzMwk
92GTKbkFjksDA/kGtzVgOhqKLxsqP/lQM8UQQ/RVPYRLnn2oGAefahGzj1wPrJnL
VXqxr8hlBZ6c+NBNFDy6GNkECZ8jkIJT7qPvGdHxu+L/tcMyv5jkXBhXq4Bc9fZu
TuNEzw8aIPq0FlDYR8xDzpvppHRqfra+ACOMC6LRSsdnZ5d8eET0R8R5I07KK07Z
9gD9PA2qyh9dHromKwR3qw==
`protect END_PROTECTED
