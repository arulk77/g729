`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP7rN/bnh+d4qjJdWx5Jhtbgk9Bb41DKc/Ng0+yywuId
fk/mNNvnTnHx0HstyvDbr+17xI7a+QoYTyDH9WWPxvk0eptGxLVuYSoSTQJx+187
HywrSXr2BcRyLPVMsa8WyLMURw/UV2IKTGqgJx4nxPtpmGupg5WapAycdRDJyD2D
70Mg/aiKLJme0nsOJHb9XA8P+FxrGIxEhfEVaxToEybnSl2zrjeUVlr6C32/w0Bf
jzUhvxCUcRvVFme3KALJCftSy0MLp+NgMdd/TFW5poLLtDE4d/1N+auezHQNYzTG
SdFmrot1FpRt/9EMJ1B4QAYAf+p/G7ZpkqpVWs2zjQs8yYBWUEov4w60nzNkJmEX
`protect END_PROTECTED
