`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48W9APDauU495ry/tcqQWLocKSgamD85g+JPLZV713ZN
Bo6fOy1jsYTD5SQotXfuQRd9tudCSjuz/flZRhkRTHKZNV0/fAmiv7yuL3ozCsXp
x3RLpPvW0eDS1Ly9VkVUzT7jMM3VYkR6+vbji8Guk4Ru2E/TbL4jAYsv+6L/dYPR
XhadQIMs3rnia5sh186JTJMpZa6Py3n91eRPqUm9NkA=
`protect END_PROTECTED
