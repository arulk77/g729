`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IdOQsFb7YcSDo7CJTtAWrQv6DAZmJeCmdByJZV0vnJwxrbBJJeMeqnOIJ1XkWIxs
sULYTkCjAZWrxihg8rHzYPdv/2t7to0mZr/erhQWRLXAmf/Yf3DCktbBqW0u+jDs
PfErn0tR96WGsBx6Qulxb3BvHkEn+MeRzfDWLvheV0eBq0Mr5LepRiPjiSE68aSr
bE8DiIN6PeeldsgHs9lp346dImSCytrafNIlsb4uwBqbMkKoq7pkVKH8n2kka+ol
ay03CsyMFc7j6KMAiJKrH5UFWneAE5yJuSi3cLDL0gdcF2YLULLyWe53Fe0YAcjv
LNqE5+luEEiq2pZDYaURKgYnAadxzHSlgd1V6FK7/Ns2rwVahoftM2S5Kvb7x4ql
ROyWVyntY0OC8XDGQGpfOH4PqDTKC5kolOfINtTZoEnA9fv6ChI4qnkFmUDw8HBg
fKN4jTPnHOnSGLmW6RnxVjIkp7TlOmIETrlU44oE6CZxyzg2kxX5fw50jDch8wCU
F3EHwF37HyliNUlT2c0P6zag8jqS3UPf9iprTe8YGFCyZ34363bk16dv85C3M7rU
zg+0dxJAWh7HEy5FsClcc5yZQjs1EIsMhu/jcs92p3PKUqyRlcecpskfcUsP7/V5
EcHx7GRWh4tqWygnWoFQK3IBOKQuHqPLhCyIF9w8IrLxPOxt9smMDD27hABYz4jP
mOtHe4fMOxvC87Hqw655xKCXU/VPucV43VyfvkJ3/w6VDh/0fsMwlbpl5P+9gC45
uuzO+Mvl54aTGkBglC7+3ar1jYA0oAhneh8XGsFNmsDIBzeZmfRHAucJTX567S+e
9W8/pk2fDw0crK/cjsH/b0MGNzpKpu8qyZzHaKX3uWI=
`protect END_PROTECTED
