`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJVrYun+bYi07QEDNYfUbUM37iIaPfuwjWxwAj7PTxKm
hCZ0sthlMiw9IhY9FrMw3dBLCup7TE/xtDGhasErympaRRQlVQWblnMcvXkBUZmB
podfqrS9mVmxg017cHo+R7Cbc5BDghw3lU0uECv9DRHLzuGvzpvSRTf1cXtkpFsh
tNkvHQa8pyuFNGIVhDs36NZJ+I/GuArTXyxU+yjLo0z8D2G07UFBpH6I/sgj3EIb
wbnreVnX+bo88YY+dHk/XyNYR+HPP5LDNrtqJgqfIEzCSf3L5111nNSbZWowKiD2
yb21b2y8LKB73Ma3HWGzYA==
`protect END_PROTECTED
