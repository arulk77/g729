`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMW78ixTzMBBWeDY75A8ZlGScw0RKiLWHP0H1Nms/rsG
IQdRfKtHX/WHbnLx/YWhbvhIzA083AzkiBfNKVhuvQZVn62ljJAkfFASeyB7EIlv
1eNRyyhzj+xWkv0aHCsj5HA/ncmIu01NLvu/uNiCTzbwHMsrDAjvRNrGU0NK1CGu
OGXIZPu6TZRCFFdEVuY2ctdxb2DSAOTqOLvONlh9FmeHJHkbblgVnxyPB+OFTPUW
16zhZQTk175wMEV0mgjbyJyoU6mnDbNIivClqhL/AJPPqNJ9Q9tOS/TEirEIlM7+
DICgne1O5viQCwBS352Oeh8JPWIuOVsLzZR9LCKpXE//oz3AsqFoqIzQncLeqjEd
Qlt84EQ102z4huxu8eT9Um4IhvHeFozE5dmj4bqXhXKZE4K9kczIGDXJHj69ADnm
LBfSDE9jvT3TqS9X9XNpfg/WT9dbb696IzxvS9Mzk7sKFQSI2lplWRFvbiknyBmK
GDiAzpaMpGsZjeVSrsLuLevSQRvHkbVDF4h+uQYFbwWJsIYadZlGvtaIZehhqtDB
`protect END_PROTECTED
