`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJgcFFN4ZCJKXqSa/fQMsjv8PUNlokFAnAOJI+y5zIrt
hxdWWiCgqUZJEwZot88hvi2EbopQVu0wVHPRytyhSrSxKJQhJu6mUkUzzXYiT8gy
80hpXtJlrlD4r09clwZNb22BP7gv0zlUdXE5rAJ++9D1e5LSB+GykOBPzZX1awX1
41kVYR3TWgjFjJSZisStzg==
`protect END_PROTECTED
