`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN9SwytAu6MsrX0W23tYez6jceeci1aMizsqsRVWdKrHn
qHCyo7QbW9gLiQrb1gqdnN6Ff8rLAXVoDfxLnt55ccmPtyG0/CV3ochh5e9lJtI6
M8DRDJfLTrZtq1wPPnAlz/BY2u5KrQEbS8fgIlJiIC+LfK4xnt43Jc/J4qrchHlb
p1NuGaP4F8GLLkWWX523OPvfaDVGDpLlN3MKhMLkG9i4z9FZ/V77khy++K+W6Mwo
2BEvgdgfrbGy9Dx7ugYhTos1oA1dFtE9Go3mGtxYNpP4a+CxODcFd+O0d4nJL15t
90GJMZIsL8q5XzsExMVt0hHQ1Kp3IC5bb/Z0LtsyEkeI8nI/Sw2ig/jQK7/drc15
i3ANaAGrkkW58XVUoxtDhA==
`protect END_PROTECTED
