`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAqcUjFakwoS9fEzTOU5/LimxmmJUOQvRdoF1JAy0C7q
9EM/EkpZwAkrDwerfy+wHrwwPQqM07d6iakmsUdokOmprZDSF4Kjba4N9zoI01ix
VLyrcwUZHJ2PxNyhSPsBvuU1VbiaCM6wCNqgXOSg6VtzmY1sCJ90XSuNPRSCcuCl
hAOjX7A4kdL87+TkXGTlYfrQH/eOpPeu31KxsgKOg1+btASkr7+5NoWPSjadBBS4
FkUrlFd63ybFUE+ZGTwXgl5i5RNlOL8C5wMFTsz6+ZO1RORaswpib8izoEZEaTKh
kLRMmtOszFQB8JKc5vkWzeptp9CmSzlXykLep5VUvZWn3WXKy3IOpE/jjTcGaoty
FuKQFFsEl7q8l4AS3VDBRMAZwS8Wxb0vdwaIJoMCnqFDGfY7JeSrCZVNpWcf5I0i
`protect END_PROTECTED
