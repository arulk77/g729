`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAl6xt7oQ0f6oKBrCqw2GZGtPiNBPZll8U8PlMKrLkGA
ujNO8QVOyLCPIcnlWKTybNxJVkj/uXjUtNZ0lqRYUmrw6wYJKKTfr/XFyRcUBrW0
KdPQpCpUoububofxYnLbEYhbVMCpEODqNtN8KkoTTwJCFacjzYr73iXwYRdaop58
UEiOUNNSaMMV10j5BljfaRJHFn/JqBNGRTSYKlLDrOr8Gz2pnTKS2D+3XsSIol3m
4EntE3oM3rJF29DeHvHmXKUR78cktisXxaVMIMIlPI/agDgAbsYRICsBFjFJUNLb
`protect END_PROTECTED
