`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKn1F6IRbMZnchhQbuqlDkuS2VZzJQb0fO2XFpcZZs6f
Qv6VpvBPt7/CrVaNhIMaezJ+andOA19tg/TsSwBm8Q5oyz4Q4OqSvI8oTs3e3IFV
eFwmnGQ75QiPc+I+uziZbgoa2nbhAj3p7exSlAyPGpQViBd4/n5NIwLLe9XiftgY
`protect END_PROTECTED
