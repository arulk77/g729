`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAXjiWn6vfU2WR8mU9YgXJHvLGpva8yvLWBRNpOODJXQK
Q00WwJ5N4qW6fn2n5mqsSYPCjqPStvNWKNHcDXRG3Cd/wq+g37B1DZsZCJaoz74W
ZsNtQuK5hyD9RHZSMekT5f4f9j49u9RYBfQ9YaHFfMa7U7NvzX9i7alJ1vVo2YYh
LJYUJjDhj7jczTe1+4SWFjwOYfABznNAVRdA4NAoS5oqmuVskgPvRldn0x74QavS
+i0UJim63ID+qODKJANuz8+hPTDAoJeOqPQkX7bOEVcb58Vx34VubQpDKxFT1MPY
99IZQVSnMKWlU5treEWl/zolJfxbFbpnXz92DlkQsEuyI9Y2sYWPAYAlX3LndPsN
zlNwkOYTWFD+J7pHthaGq5uF1UyNrK6dpm7bb+cXbdYTgc6NG82Hf61ZOD9E4vJi
Tmq1e4EVnwTa4GYTjUGw2LSRHYzRRMmH+Oiqj+Fs3go83WtE8Y6kchckOFHLNFgv
Eef8zoTKoV/oYCG1tQksSKt908Psy1BpbV/iMYzl7j6tS3C336fdvQRvNJDQwXpm
/EpGGbZhjYPZ1L/Z4j+sYNr7liD1nvu+dCIimva/+87REVyn7ApCFL7pLsHZWzDL
WXLtseImHfBZ0hwMiSdYapZoHJQh0DtaakSy1C+53yp2Isan6PJA+Rkf/lbJCRGz
zbi7dudZpAX0AK4cFmgd814eG9e9MhHWyKLBSbM/bF+Aj7Z7sbcnsg7W8ymukkkL
kepG5tOO+nVj2TM4qwrUcfK8MLXgL+CP35+LMahOXGRjBttAOdwEbHOU9VbPsjj5
NqNdGHl575tNNSC2DcH8UEr8kY/XE8pfFuIi2PrAo18aep4w9Cb81NkqQNirIwXM
9KbuhmSdoWBjZVh/+7EadWTpuaEzGcNf9bsWjuL6X4na2wkq2uMtamLwVqkjUzXT
KhldDecWV0fKKt6g87wGNpCJIzvIhHyJmbPCY7o7iTO3jXzcxCj6q26P/VjJ89cm
HhCiwSMCUMNDX0hLIMJAGQJTwOgsRV/nmT/1t0RZgDn8dCFAYvbJV+9pyPZnuX/e
7wdFM82QSYsxEpFjSYM8fxT39ybXT8scv2oKo0Y3AU/Hd/7OpiWyAMWDgQG8bMkc
k4YOvQJA1wio2fjk2EXOwoec31B2Vk3ckRTaFAwyQUc0h+QPavwqCW5zGNPiCXx+
eY5BMvl0BHnsTQryxYnQ+58NMpFroD5YPjlJXTG8kueWpVy1VW/S/xUbuKG0X72n
98ADRMpElrittftrrR+QxCEr0snWmSd/b4eV2+5n8zjm4I93Th5YXjV7f7DW65sx
Dh/gXkyAn1AZu3QDOUwIfJ14k/NvjGF8mZImU1zECZ5zjeXvLGt/1o5vobctplkZ
8Qmeeskk2sE1HRUghjZI93TE/LwiVA3jYjwCWuUcK9hywifW9VsEYo4iPZRq9hz/
c4FSO5YupDjsMUTejMMrnl69Ctj3yt4Ez8DzGTMEcLCy4YzTsOMJ1Xc3DgDZT3XY
/W57KydDjqEkuQiSKGNW5hJ+X6zl0RlQwTNDTC2NOiL3ZYk1gp8N0pparvqwcLqf
ton6YeAb60Fi6byIeFIVb1PvBR1s7jwkxg6LEuJrruwecM9kgExnW3YYIbo4cfBv
4gSqrImOK7dLVY0OtTLiOg==
`protect END_PROTECTED
