`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNw3JbmCjBUsnCZMAh3OodqItV3/lxqTXWT7jpdB4j4sP
xPma4F6+oVMlAvZ3CHom5TyRm8Wb4j10eeP4effe1QXEm5hHXXY/L1zQUU7P83yY
UJ3OBJLwKUQYUaMavhvXoGfzVRXdQRiMJZ1BwLnRFJtM+Ohv9XeLpeNZFc+l6QlW
vp4FKNxkU8uGHYvErCO0Ib3twAnqi3MNk6ImRKQqMerYLCMF9qePvZoNfBjX3gHQ
SYw0oW4JW6rrxrDefsDENPvdqsVMNMl2ADEDMx21Od9r8vIi/r7HP+djhJQSEYRL
ivzkMvZc5IqT5kSXxYvfB0ZKQ1PdvIjC87djEzyBh7SnUbOlx1QNPa4xFxwm+E9J
qeBYa5es2Ot+hrSywkBZRyejxV+74Oql6Q5o66Lm7lj/f9U++EJNhSredTHHuW0W
H4RU2F3PbLc8DKyy5Ky5EqNshgjuPbxBjrS4xfw76rTG1z5oSyHF6rcZWlF2a7jh
u8YjCQMpqcT/Zgu6JJdhxI3FhaohzZsviuw/wMRZnU0lExTXMJ7VRrzQwsdtMYGj
oKe22Pc4I7jxlp75MT4cO6t1K/ZQeXPulXRNHOHbImNZBShPwqKyR41VtdU7Vwmm
VXW+4JikpZY7Fxa4uFOUbM+RCYcopPH7CgDFyYzAvvMlSq1UXPxmLzwZ3EUfGquv
SDjO95sHbXz4yjBZ+meSFUNrSjY4PD4pEg4QkLpZjkTbkoObBAOxy0OqvtBJINgH
Raw5FIzMZzd2XLcZIb4OammDZH7VZdrrl99p/NiDGqn9BQ74ODb98jis6JfOgdc3
uNHqcPgEY7Z+P1M655GpBTLV+iu4GYyTucXLc7AWxeiaTt8k4K2SyF2Qo/Erh0MR
ISFuaDRvpN+oiNmwSsBKnIdiVu51MehTI6W9/mBjrHuoKgBsM7AEVkDq/sdG1l6A
NPo6N25e0hzDYXEr4Lmva3+hKwELRqwBd0N6uakQZNEDdiYgw8UnuL7Yo7BREAQF
HTUiouCVWLok0BoIiapo3rdI4Rbnv9mqGATlipYY9FE9C40tfM9j20dPs902oYaJ
UGIFyU37CkObhr7obwO0Hd0mEg6pBAwx3D2oVCD6R7mUqatUM8nVOQaEGkQCTCL1
8QqHMFHUU43NDxkPpzyizscYHS5ZoO3Lxto4BW3XNI6rOtKr08N0aUJotkIdyUri
RVWSSO4V7WzAPm5dIfC2yw+oEDna3qndWqI/5Fq9kMSxLEmB4rO3BPS8cm2o5HhG
k30OgeRFBzSDmv9YpmpIxFqvpd5COnLBt4Q4wI7tbUlRPS8sjD9rHUdwx94csNq3
J0A5OZdcVbny9EG4pLWh2nxIagqjUFBEPQq4rK5Xzjh8om1r01MpdHdqH6DMj+V2
sIP+XsNwNDJ6OESIIYjdypcijWkXp6wHJEU+Lgx5ULohrCCyUXOtcks3v2QUYxFp
WZZ/cblEGAC4d6VEBX0fLNoaJAv4hIq1JmRk3ox085UCzIpn+9huEz2Ipivyd73M
5wrePz9sN4HvwXuFimuyORFhFWoMc1jeOg79/78VKnTeh0F+1u5D0cM40IsSBCFB
QKdXet9ZAZta25iJg4tLambdjSK1Zb/uyPmr6invdSgtKDpID9sfVQhXxq6jjkyX
Gni2Aw8ldWWUDDAsKtsicbx+eUuZa2sD2aycwfWvD6xTcPIrD4fRugX9j68Mj3lM
MtlNK+0+uYD2iQq2LSrNw0SAq2mXb96bWS4CIZgeZV+vgJ40obw4MHFyFwtSlLvp
+700El1b7DS3fsB9Nj51+oNerIW0xwHLKSjVseVpid2cCvXKx7/4f55SIfyLpdwP
J47hJcMScf04rFXcJhNBVEvmbXLVm5U3hxPwIo0+0EbDsDOs5kUVuY2rcW5XRzdU
6pbt/DTB7rumXVXH6XJKHSxpXxmRL0TfkqjeUQEfMed8kSQEOiPi66WY69fRzcPK
btxz12SSkqS9D6qiXl0MBNK+cKwZliD2qkS4IesT2HwqdU0rFFPjGQ/TnssmcAzY
32Mo/JBFVjCRazAJq933mr8KN8/KCSShqzaEADPebVoRfdXNJTdAtmi8KoAvqeXW
AZd+o3RivUT1RUI0k/uYoX6vzPxr83wcAijKwtKVKJwzNWRBxPVt3bAY24Y4ViZU
+6oLmGS/KlrKbiuc4oG+kSXld94qIE4dHPSpHgRc5x+STjxfpSafZ45OLdq/4kng
6GZ2JCwJr2Tv/NuM5djnL7htTnop03gXva+HlziVtRPBZrUqBKqAL9yByH6b0/d1
Aec6a8bNFTdKSqwoV0ca45EveLAaPb8pePqwsZDK1H0duuVCxR1DDUSiLqT6Q+Dv
b9b1HoyxKCqBYB3g7rBVEr1WZCsIzHoJ23MALpzcv+0TAMZQKuE8ZKjJjuWWuQoY
Rv1A2Q+2awS/qzpiXvfGgbxnx5YZBu3ThbWp9tBUjOOwMsnKOAIokhh6yzoYw59I
LI3fP96cykQfXslK3EZaCXpUr4v0IUp3LTvV2CZtUogF/DzQFNaUnf+wGP0oKoKg
AWrWdS5gVVYb07vhbABH1rNrFoDEEYVTwZcx71L2DwsmYy7BT112AUCdg1x6iPXC
bYE+M33/vcQfH3mp1r2MbFGCkQWiBDkCBHxVOlt3YIbmKS+MUTu3VhPrThdVy7A/
aO/mBXceVfGTY/glSiLN3khG4VrKNqntAoHrNTKw1Rn2weYfEvI/aJiEZ9pCZQqj
6yhGRGkAiNii6t8Yd2T2JYFfQeDDGq74IEXf3ukaPz4qN9CjzPDU0T1HFMUfJq1g
P11/xOqJK2BRzCO3XD/YwZ3/W56xTce/aVj7xbGL+U+XhnIi+vVWzfwvsed6qTqd
PwyWE4M50C2K6/+TgMjVOIGbW2MSCoFMktBYllO+YzhWM/e4zjYP4xWEOc7gk+me
Mdupdi2p49j/F5fxJZiwUD/SBaf/K5wQ7Y7fD/MKm4qzq3DDNjUzzzY5Hs+WCRqu
gFKLzQp6yhtAM0zCDr+FeqmUNJwy6LAe12y+WcaHKaAJbh8K+k7YUPEQCImeHzfx
Yi4sNRGFT2nGoqj3c1XagZ1MFoKF53TlJD+z5Xp4qZbVUTn847QxFClupjXKl/N1
gTC3tuGwcZvMhyBsJBTQ0D694S0653MVnFm5vyXL4pKtsN53NdY0Os6Ol1DKTRZB
g43CcJTyj1RpgAS0mP+/HpX0fwL1zPFmYqaMZNfrsAQ5rQ0CN0H78KYM8SoCfnjv
WnlGaLQu2FrgzMHQ9/zJ4L/bJp+WJFAUE31f+upQ0Q5E1M8Q5wcMaAQsFLgVdl1m
yA/rH1CjVewWcnA5x6QGkM4lE8To39bATtyw/qrEZC0G4VDEgwzWHs0CIOYkBWNT
9DHDsq19OBpIa1N8luykc46cFQsPeqGv6OEueZWMStRoVJCOFIsmCuGc85sHRCS3
NExyIabRI08HBUVuqznhx3j1IW3JSk/qy4qr7YP4aiOpL67VG1DunxFAHYpehS2z
IMKI1SWTkkQyg7upCjGITvrHVnVv/PM5dX4ojDuGdUqN12sZWqF25Wn09LEtp+kd
yyMbntCrjl/8XlH7Wi0XrWOIdNIN4bSpPEENU1r64pAox13uUpdgkRzu3r5UENOM
lZk7r+y/82VpQ/7xrJqro12bEoE5nSzfpj/eStsW8wdcjUUp1CwP8OOh3+qOk4Mz
kiXkiZX91dck+yFF7vr5jWWyVGLV4TOyPq1B8srgWSi/DyTbFHFUv9Oj4KqznxXW
hNYZu5V7+jLGl74pCu9QaABF3J1wQxIhWeVC7yZOUTpzTBDC7zwnw4zDJcd94xtJ
Ddzi8d9aID3Uy6ZSUXK7u4pR/h67SXl1afPRqo26srn1aqVyApwfdxsld6wt9VfZ
hPkTjLaC+9YAR+Jqq1dozJRAFp4DyZuSRovViRQUplRinZCvt5jow9+PNe8l9hFN
sBN0xm610ZDBHcYNJxMbpqMRTOtXVQ53+ge4jLsp1bz1+5tYmW2iufX/3oR10MtO
Vz6Gw5hTYbeL50/XUxHXjGkQMrm5N/xR9M124pLRP30moU1UYuPnUbwiSrO6OXFY
vgQg48GzZ1OAiK/vs2DkitM3bOZti9rqu6P/AfNIEQXVGmpSyvJBvrOUUGBWROFw
wcf2sjAIw08tSCpB5K1oW4d/xG/f5oPDn0aqjT5qSZ0tQbLYOy+xuVpFI8ECG3KD
8wGCQC9v6mAz+ejywqCpSE0PSviMD/PDJKsuHHKCXPR97skoOul8EMgbPDGnEiFH
Odb63UUeeC/se8MfxCCxHaQFJLiipQsQoUNxzashQfsLvS9YIhrHpQqeXNwrx004
+le7yfU/mZ+tWDzVa+6bfVab8STjxe1PN4ayl1DWbYen4clSlBcqoBU3v8CabxK6
5/SJ+GpgYMpzejgLR2qie6Jc8acJu/3KkGZaWsqKkI8CsQnaTNG9WqX6C46/ngTj
iWVi6VG5kWnN7avr4GoolcqDmhH676w8lirvjlmTd7k7FsRfK0eqW7dEHR+Q7/jm
ckTy72Us8+Yui5kh82iiV0/BCH60no9MCG5gFqtis/qalNyACYjqv9PPeVLxDijH
yDOi2rsUD+TjJCflZEQUMS5fYIeAQyJd9mnEds8v8uLUeL/bgFmE4Zz9y8tMq+3S
UcYGZII/5EH4Vh2Srrx1U4u9ZDbSA6Bv/LFK/MlLyXPYe0CGqQkOZmW6oeuprljp
NxWclYyDEKUVN8ajsqVnphs5bD3dFm9LEtHPTR9vplaOiFw5bJVDNEPhGsVefR8w
UDh4WNRKhdaBNMvA7/FLZOkGGf7LJD88D9jvtmhL38e682Eu2KK+gWRegzAjM/S3
qLDdQ807KjMsCg+H6fe/ymxifDFX3y+S3dUJcisHEOpSACyTGNqqnJgoHGZBPyB4
KaPy1Vj7OlrcBLg1TUN8u11qKrZrIoN+y/OQjfS5iihCaiI4Eo4GJq9z7BAwH8fb
Z7bNuBVvhTkjOfBVzXBJebIh1UA2JMmFuYP1YKEKfYs27VYOx59NR/W6smV5vY0U
AqDZ9l94M8qyjFl8DVDOJT+/2PYYFG9CdD1eGg/doht8pEFLPE96XbOIy1wetSUk
Cb0UCQS4TmrYLvtFzGC8wnAqPEV1GLA3zY5X1cTtXTAiqfo9NxnyZ9BRccW4Y00I
UU5Zg6cNvLSDPIzNb6tylwpzk4vIE9+mCZ93vcpdSy0uAIsA7yN/3YNnrtQU4t6l
+3N/KYFqTT2yx6+blS/5hNF4FW3OZwGoq3BOG3k47wcDxl9fnVz+5WkZ02svY+fh
H3sEx/TOeIc05IOZMgdIE5XbFk2iDAc873FVcR3oJe3hiWPr0S1nDRlZnHx4JyRI
X5ptuYxvxhlwWH+sRGHDu1shb+CSffacB8MfufJ9bh5JbgMh2s7CbckTKARPBRwN
Im5Me7wCo3FMjw89tUp3yJThlxHjM8p+BZXK1mhCcXoiDOVcQQUR7L/P27kpLx3/
KzAkeCkR23VQhsx5sOM4gFaQ9BPvCeenOlpATZ13BxngLIQ7RN84kxr9oCHxGP0w
4qbFa3CIixiqrAV9Ec+UlML9CoFwjFZxBKKIsnnT+QDNEDDDxQhsomabmyLWlwPS
CD2gBZIy8R8eyOyvYimlE6kP3Dtl/GEKmusrQ80mP9BlqLwgUFS4aifbL21icWLD
9CMPZuZwb+YBDXTVJ4VYNQPInh9lsAfFNglBAjvX6+CESPQZPIr6sh8+v/2s63tg
Wf0JJnH6E2sON2XMMZBH8GrSnCETMP8Dgwdyh6YEjgik9JVbLp6piKwqQzsXHRNc
fvOPJQ1SwgFXemXC0C6BOb8lBYu78P8P0MTRlcnDetnh6jlQQ7e2NbG6Y4brir80
vag9+oxWgFfkSQeGyXMl6W3aNtOH56VtNxcRscinIrXyKOQNc3fOD6lJrIVDA1Sx
PElg9DObSVYgddlZpEmJoA4mHx3Z8vNoqcwRyXJo2GMCflsU+mCHl++saKcLVCzX
jTBtm1Q32z3JBTWEjk9patMvsR0qdiQtB9oxCXR43rpF3onWE4qWcGfNMjfzPXDe
vG2w5H9XO66a90xvMpkpAuSSp6s4QfvTxxCmoIO5nSaey+T3JDcVIZwC9wqoQsbL
+VJYWdccU72Rh8KBtGI4+7/F7gzREF6FgsvWbRx2SKDId0gD5LM1DBCAQOaIeNsA
kthGX5o7fsOdJaRo+IsMqyrCccUY4UvltYk3McVV/SLx1rzxeAwf+gxv6QCAlpOD
amzybwUAVmKrrcaJoyLRjdAsVet1cMdh4L9m6OC0rWomBCdtkg8foA5DOdHG5x4T
icCX/Eh31RZaaUwEr1T6IChinBpi+6ZkxnAp+ey8wsMFfGhpY5ncTkvH9pUS+ISW
dCQEgUYJ1G+Y7wwHqxR2ziid4ujVORcTiLoJvy8N7u+jQlVgpV25iIRenm/wrcHF
`protect END_PROTECTED
