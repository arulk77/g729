`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
1W8HHO00qTRh2SwH9iLXXq9INAK8cCKQyMazZ5TYA9PBIHqlTIE/Xhj5PM2m/OuK
UKYS5I5kPuvX5fOJ1VfyyQNtb7kloHFSwtx/cZE+1/FJde6LGsGEVpZ76fyZO2rX
4RelWaXG16CnpXySx+jmWzFwHArWtq2GKhOctt6xFK9Avj6SErEvZydQJFNeojNK
iKtSGA3Au69ybgTIJszdedf7rRm0A3z1rDFAwuSQ/LGrhLjeWXSoXcJUcX8vaF5j
XxdjPQIkQQk60iTcj0unv06sO5kqoYUfIIIs1++mkeMZOFAEbstJwtZWRfH1kCav
ZEAw+NhcKu5hsXn9Wbn3PEkKH+kQzOw2DY95PZ+kVPsVOClrq/GtlyR/tFu+RY5Y
zQfoRA5LdUpiShVp6QdWLnWKreVmdh/DVCTZI86A2ck=
`protect END_PROTECTED
