`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QNw40IqJrFvY2E8HYWz+j9KKfYW3D4EiBf0BqBNnGeG3C/K1Diyw9oBLijsdfdVF
LBLK0T8jSf4Vmt6WTx0KG7bRkuSGHjCocGrn7G++i/NcDvdxv8Rzhl3cK2qP1G0h
YEOUZrtHAA2Gqu2Wea0HKOaK93KnXdXll/1ZDU8Kyap73sApB3lozvP3WbA86FXv
`protect END_PROTECTED
