`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
whfZdEhQhIVICrvn0VMg7m7ClPWP0AgeFZnv6jRLYTDlgMXkZJU5i1K4zchauxyI
CNY0QvbZv5cnlliC1PScRWoOIUnJoYn98tpAMvbJoEByZrZEB47Z99kV7pM3o8n2
gnfESzxo7lf4nsZTE1vBjnfLRJlfIqRIY17Qv6HCYg09KbHXhS7NQD+AK99TyUuR
EkOC4yUfOj7nOj6ryBQxR67lJeEOZbi2mdZIbV3f4bMUmL3NIOiyK+RSxLmIL18Q
Wklch9BOq5isG8VdRZyuW70CVBSChOZT+8YtklAeHKAujufcgBj89xLALA4S9ffy
levFRCoGzvxJ6rY9MulyfwjDbjdZAfDSBayj8d/LTKJyJ94CIDOwhdnT3mRaYxc8
`protect END_PROTECTED
