`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
OZmTVedTtmYGy7jVk7bqJrGnVz5DtzQAMy8SWcJAwrhYz1u/1CK3wc9vT548Gt0I
gVxJzye60FiSM1Q8OE+p/QrKAPzCizkI3eKdMP55buNSbNjqgd9OGBEQnr90wx+6
y8QlevkK9pkGsoHKUR4x1w05ifwlZqtMlFbvzC/7wixGFr3W4+iFz56MJXtjB5DX
bEs7WUAvPHUzV1SZvyA9hRmjIEvnEyPxCk4y/O7zPPlfFEqQ+ACXiKim4FIXp5ZO
SnSONpTD7FiA8TazTEXyjdE+HjQoPF7rcVyUU2S8PmDyH92jMGi1Mxo/5j0TNjdq
VzCEGRLyPGESiMhM9fIE7IIDqAkoBmTNO2nyTdafxE27G4tjaKGfWmNL6t4iNTIN
RLQu7IvFY81JUk2+LTLQ8n02sTUKMd8KI6LpPfdS7EfXgjh4OcuVS1VD1ST16XuS
IPIXAJgdUxOzDoEKFp/w3A==
`protect END_PROTECTED
