`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKAJAlTd1b6ZBeWFqB4J+BCA4jWN27zcOV0ZXrA2FRac
Pi4r3SkVh6P0GKA+IJhwUaLKuFF4RnYFNhljuuytalZQYjdqAB5z6Te+cMJ42btZ
MWHeexbmEU5X7l4FUlaiGOKrKgR6ankLtI81+BWJ4kUuQ9Z5FuL4zQDMWzMOPClP
pUv+9s9KkIiEQJgwNnFQPPHgzSo+1mZUQzsE5aBJWpHtRGjMbR2fExU08pXtshDt
pFjB+s3XU/Xs2HuSzAGVS35glqoR01bya2m0tUhaMPETVNZGoayJ0KKz0tviZB+Y
2riJRks1hyJaIpPYAe4XRxCUqQyZVKhxjhjsptdggIL5BvNqPXQqrFvtxAhpbAKB
iJW/EJCNfHxd3OTHoXWYhWVM0RGFA9EONVyJXHCFsVP6W73TQ3zi4gM3VlJd2QKn
dKWhDRp5D4CeGvO6Xpd8FPLNJG61WQ8MgCPKV1+41oI7PLLpWlJl6tbM5xH7PPx9
nRCeERbK+FySUh1KldELhnGCyYjT8se4paw9C0rStLJOzb3sJbneiJg7pBVPsi3H
IZDYeuv2f0ROcpjgecvutPnERe08duFluxhAfHvW+u6cE8GTwYbcX2uQh6W/nbYx
fUy9Z7ezAwz/wZqhnHHCMK7//oALyhOd26zKhiejTX+dCVSenCaOQ+q3kfLa1gzd
sK4W9wuUIYs4qfG+N4T12yrGijAvi4qjc9cV7zj6PvlaXPeTdwheE0JmT3SKG45i
4NQN0X7ug1SJFplnI1sL9RsaB+4/y0g/h5YaTujiWOjW4969EP8aL4hQfthrKlUW
lABRC0NrzbdBofBBucIXbUetT6MzDujpEQ3VID05ZEhOtnmVq26xx/s8yaY9UVCB
nuDrCWfwntekf1ddgEJPrS3wM0lL98N3VOTq2S5dfB0bh5DV8ipYrTjDG8k7kWWd
YHueq+iapnt5CI0GgWRCogP7yj+89HBcP9NSWLHlgbciH2LHgREjA5OCTX/gJsly
ZkR6S8e6Fq+F5pV6OLcOsnz32cBiJyEfr1eIBDqYvQ/l4yc1bee9pp9VLEgtlIzj
eSZcoyvfAHDJeHn+XtkI9DY6KTqPmVhMqj8Gzm0UqI4BB9ZLHgLqpUtotg/FM23b
kGnOlB4tuzTTvZRSSxFtjWWAI8Lh42TnysSVpbsWvNyLYnTP5B4ejLkHHxuWGxCI
mBVuRTnf7OJ9IvvqrKyyq8GecO5FSW5gOlY5YvXq5BQwdNHd0PLsyOiomEkRKkpn
1mbXVf2WxRPtgf+ITg+ci3FDbP0KBGMK7Oomp6Gxhda6j0GdWntmZZJ7RMYGm2vA
IsErsFyumMk0MuJ0Tzyp+ftdarPXIaC3+v4+NVul+6yZD+ErGg1Nd5eDlCtcK5sD
GMwxKiWMlNqo+83cKzryMh++ZWZW8nVTETpryKWY8B1AKn45cUc4OmaQUz9a41dp
eX/Vdu4P8lKYS4T/jhygY5BPHM1kHcJbTj+kqmYYkHGooDMKyFfu2bfolp418Zo9
mrKCncpbfrPuDCM1/RN40r1zEctS19XWycSo4waNf17X/a+OhydlCrSaeyvIx9zV
Z5ET1XNG/gZZ4LZA1ZA2tcEX86CEiKmCUqylGrJHUYbYHWFbObCri8rb9n56iQk9
eTHGhqdZPo57ZG7u3oETcTUwuYk2LUc96Wu1DdmgUsPPgfx9O0yBPSJCBM/I6XZX
UO5CAQL1SVH3tABTm+/asdCauamMhuDhZ39YlkpNqJeoMl4+PVayeBYtCNl6GPg8
6wdwUbv1k/jNfGUCbCywBJRlGTwLa/OCX2Rv4Cz7cymkzgrgoG/02wDmvK1PxaNz
QiMOOQa9rQ06FiujoVq/Tv725kc1vZfnJEcsfUE0r2D5aBdWkYIZZgYT4bDLS/p1
U/FVSGDwGNTNp7+9658B4kjx2Nn/xpEJ+u0h09G0esXBE4w/mzr83MbmYrwlBcSX
+wr3bpav9O3DhTsYNZUt6K9Ipj20Qee7DQBCm6x16kZn3Iz6iyU+c4+z+hD54hXZ
/iS/dzV5h84b5uUZ3+rPXYvRhYgFKLtJ/kyTKKqsxf5BnrDgisPgbgPijjLdBG6G
oArC8zZDzLFGtzK0NsuxKlzIstaygKYsThh6PMfuUv/nI87IvivQtMM7GeyLh9zO
Vl/mjcbnaSNpFyIHqPp8fbhr/wBt2EUeqb0yFTLg9A1vzGbE6KU1Y6EeiKX2xA5+
b2u+sTP63ueKuD33N8j6CIEvbR+ezkZBxL1f07PoevMqhT2QjBnoL8WIDT8M0A7P
okHiatZiBIKyo3Lbc5bGs/GVjvA4vH5KXc+p9TvYApxMeYXeYYLUyStSaBfcxbxU
Vsz9F9JrUWNwaaTDx36qBBFFPolOO+B3rbnxGkPk1iv+Ogd/oiVVTYV1wwRWJxDa
taAXLseIPzT50SeVPN/ovNZo4XhsgpVsbsEH4nMVX/0XDUchOz9yfshkTXVYDKtS
+iksxrLHk5JO2huuTtolms66Zx/qbggRgLhMN68Z8toSLfSyAQC3XlfUbWmkI99K
cAC7ADi8HsWGsMAAE226VQLv2jh6E2FcHHIdXFfVd0i0H1P0kuUGbOKmN5iTqdqK
i1yxQXpQY+9EptGYQvYqzzPkBYry5fUzuIyBIo061M9dGtHazHC0xd9Ni/+p7lQu
gQ8SQD9LIZhymohOx/zUacKnCyNd3RZfhQ8Jj4KPugwUAHUl2b0PozGxTP/G407u
m1rVl7IqmsZH0BSITXi7USkHDFwHmQZ9lOnuLYkkHIZLVxItqiP3v0fz5DkS1OE+
hej/vthwLWK/4HCLQFUQqFClVTucoIjP6YX1kFQWxaxGtPeVPVxvKgwWSAu1RjdY
2sdrFuZOXn5N/C/9G03UtgAgvTmjtV0P6S7UHZVBUfyoHjMxKpVVLzkKW7wO8pqQ
5R0AH40e9p7/1AuMwekZGc6XcUf8U8ZR8Dv37ecj4bpqlR95/0C92LPEZfTOYW6+
UYDNWCMFyYOoB+xKdGKDT5KURHmLTnU/2PZNYmyn/PrKSmAGtiIy29gSZcu9XnUJ
KEctfRTEh2wKRD7RGRsWS1ttmdSVVLe/6kQ4XBLGYQDbJjSLf2AlF/fzfxt6aOA2
iaFuHDLKmgBrIgBxG8k2q2p2r2C5z2OO4ECmd5TheuQI2lFX3H3cKiiuOu1/2/yd
ys7rZef84vTw4EUuL9ofI2soEmICqqF9max8hJ0XF660xzCkUPtAIbd+2Z6Tw7ho
lFHke6WFrdLJk10CxmoJlEiXhCNluQ1nl0jdAOexonCCFlDYAdufUCSLl3msdq7b
BO32hx/qvEJH9DeiPVneqJ1VTrZxx46Yq/5M8qapBZlvd2AftkADd5SzqWyHJvSK
TvY+s/wSoXSPIfOTb0MKNdXmkTW9XuWyCqomCczHnVdatdf+8C4nGS1piddZgYqe
Lk0P3Z9NyE37LcpHRCtjSsmdC/LQMUMhTXIQ749FLQ+7gPg7TDjgmPt+POQAxAP9
62y8bynWB4Zg/gM39r4fAcYedDyLVOdD1wk/6NMPZDuRrLX2OzNkEL/ED1NYbpUS
gqSMbZF1bn6lVov73Pc1jd8M4uY0fHi27vebCrHSeJTa5EorbvMJmnRcdriVsMoT
cZWea49bP1xTUXb4lG2SW/mPGZMqKkblfF9OdYCeIgy2ocU97QatD1n3c5IHbe2q
tlSXLcw1g39Vfp3RXcaAVZxJUqY2coJzB8/xrpgsVgp/9cRedXOVDmhdYJmYAFKb
vrtyKfNC+3N353z4roIGFoHNgQkMAcH5pUkhWdTi1c/5Vr2KK+2PG3hpl2j0hmbP
`protect END_PROTECTED
