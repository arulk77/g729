`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFRFbkFj8QhNoIzYNTmA+2XgirAzjkkr1aXblpp5li0Q
Ldzgw3pRzIRc7IMFzGIV0rQ5PfMWupjOk2+TTBcOOmfyCSXYIqEA7ObbUSt6B98a
qezW5wB5mFQkh2LCXSKGnsuh0DP1oVmtmk6YiprWA7PiRKfEInvN/DNNI3J7M+rR
q6fVSIiSLVZnb2hl764dY2rupFovTQIYVnYl0Ena13UOkdIJs+d1C8eaDcb8HIW7
69hFM5jyHI+MYSFcy9v0L0YHNhn99142MrkXJe5wxfdEIAQI95d+6eCaLswkwqyT
2T23TQujrR6MnYGMbIcnjxlCtgHgE/Udbf3YBxXYEpXirV0a1MmbUl+AT/ZQ0uN8
42hIG7bKDao90U3QK2PSMvQbyR0+sDLJ9/fmX8EASF4=
`protect END_PROTECTED
