`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB8fvobOExnNxFce+kCOu6wZwPUq8HnlIItF8tVCkYLy
V5xTXoGu1sQF+iPlE47x3hTZ+kMXLgQcD1aB4Uz6neEUV+eDBv8ATS9kCzSNSWj7
Vh8K/MoMdaL+Qdxjnn+pCtDZRVIytqoBH5FRTc9avtyMtywaasZ6oKbOFd+Ptwae
pKuEeiDg00dXPQjJb0BCS0++TZIFZB4lO+C1nwlrg5Us9Qm5/Kky5x7mbV9w4eMr
7QGjfzlsMj1myUz9AagvVRr+hkyLo2S8TBvmdpmx1vaUkmhgJerWc/ZIBfYRNinP
qTdxvMT69TOWDIFSG2Cm4vCWmo4NoRngJY9yJgpVUJO7wjsxtkIqLopIe3YH2pug
`protect END_PROTECTED
