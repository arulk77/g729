`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCQWdqDa3qME6aqg1scuoD7kMJXdSpXNz/nW7LGlWu6K
q441GcC2kUL/7ZhhagudDZtiBEv+YWRxfwPP1buTmMZlpUsIxdnDOTxN6RGlKipi
mQQoWN6cj2DwFI5/QeIZTkqd2bz6rW5rzXAGeirbiilKwE78M7gP3LqvA+NPOU78
fCMryhqpmlwYR8AYi8iE5/eAn/ze/R4PKVKwrAFJMw43fCxX+Xs//wbfwtN49c9Q
zmDTkiGZ+OOPi/yVY0XJ28zrKe48dQjlX44acK7HknZ7+BU2WedoC4hciUAI+FJZ
haZ7k9oXvlforpJ430OpMuD2ssD8TUUvaMTroj1CZ0qtu4VOqpKRmEM0rfyM0MYe
q4e2CCaO36l0Ykl7hKcftUP7TjvIELy3P5ZK0o2EBq2THau6vkqyM7AI9BPId0Xa
xKj21s+yJeFitOHuMHEs2MOc4fUJCj1sv8sljdQFS1bBQeDtdf3XwTkPxDvzGzSk
CoDFOucQ6bFjCrZ0H/0Y3sX5EbDCH2GsL6lz1wrY7ANQmkZnZ9s8aenHHzsT8kPI
zz65Y0If8/A4inILZV0UEzWXTmtXkIHwSuf2CxjL5sNKLTlWLAw1zWXggfHHogGt
IKmpKjXGVcfgB8GPxC+5rA7NgDLFc4Qpulx/tDOqqmit/wt8wtsa73eOAt5GFU6I
VSxJB7/a8HmeUfkTRqK+KOfhtHUVTp6kCjPnSRUSExtORr+T3U9O5VxSWhKqzDxi
KwuaTUPEVaW4m4YC2nQbH/ZCnN91uwK65oyB9Lze3I2K7aE7RyqqyTMrQ5XqM5ea
Cc4nYKcXNuLlJybhfyhD+gnsExoL44xFuOUXTGn57es=
`protect END_PROTECTED
