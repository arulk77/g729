`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu44PvLSy/6zmxFBg+R3m6WnrcJXQua1hx3Y9Y0oarfmMR
9sAV5JwNqB/2fCb/OYj2BV2cZXP4gsPu0ETiEAhBBgv1UnR178ePQAp+25wvnLzf
7JP+BnBXqN3myOb1WD0Cu3zse/TGhZ7nyuKWMXgesJCtWujRVWQq+t3LkvO9MZtS
+gQivpADeKUgiSwihoI1nqffVyzfYDeEbRIIRwHrmJUz7sFWt7Jcepygm/tVhFLt
kMjmuQdgQUFJTSd3UUsIv4Q9Tc8LVqHK7TTnlk3YUm/t3N1bZ3QdHytpksY340JB
k30cDgmDphQnzrywHLw2rQ==
`protect END_PROTECTED
