`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAWwPI6pAvy/h9h5Nw4itVm6AIjKiz7fVlY655yshw3M6
Tl+J6hW0OcJPh1H9umNLLIPw3iVgJ82vOG+tRGCEG7fWfnqPII0ebyK3XGwPxrG1
mBgRWraMfke8DvqWFvedFHu7MK0sEydN2zEfUNa0LPMzXUVSLzf+eX11nbC3iyXg
w0X/cop8agksCRG1Re0vzBNtMxogSN2285yY45oaCTFnD+dtu4lWaAljBa+UoLgQ
ScWstIZ826hxA5lM+j1YW9kr9geZEKu0O8HU+DxCgPzdaCtVSY7cExgFtyWbbm2a
EKOYGJtkOVWv+1XUTxuBNGkNSfUZk11GJqYH7/beMm+Vex12+aWCzz7egVu4tWqU
hapcwimZo6qRhGVi077merPmdulH/+MyOQ6Er5Gk0EWDHtfO5G6DMrqqlGwz9GGi
jECvdAvG9Po950CBwLKrrzNQBTgUchdnW3d9yyUenIRhL6KomrpwScZSVJ7mjiEd
A5veEBdWq8GjTR95nB24B2PmKGUtjJX4pIL7/4d7DjsqUSiYupPE8TDHMFCiHAhs
Brug8GiasZpO2uo+uMvzAhcBT9zpspSZNqrFjjoPLbSz6j3wiM6et13QMHgKJ6da
Os4OEFwJ+F1jBGGyLFtNu1e1JTsPpeKRsZXMtH42frrnVAs/IKeK7U18weM8XXo5
czG8Ga2aqLDEGkkwiVQk7UWZRg7dpRkHMKQ+ghsS+GjZmBOhHkCoT3M8mUgfVEPO
5hY3tFNc2AOUtvvIrnJG1ZUWZbf0iXlqg6GEA0vGWJukLtTsi8MdPtw/+Qe6frN0
Xc5lY2xbUPXYyk2hAZk3/6f7v8tnm3MtFdkiVhxI4fLx9VR2uwTQ6TS4ISilgS3l
JeVL2ZrQo0JuygZZxfQom6j8MWxO1qKREz5Rz+SQRf/3Z/FAuWh0CKU0aeYCVp1n
10ZElptQYyrqVnwVpNu6cqA6ZN5/IMu6UVSIVu3OxeD1MBg6JBczAv2xS1OFZB5U
rcaOXy/4X17VvKqia8Sig39/9ufTcXZyOVuHFIC0V1bfGpuELKJlqfQ6DeRSPxQ6
zL1FuMkZxG6eQ1vBgfxWruTZj5FThWUWo3Y8SftdIICDjazCI0u4lR9Oj6ENwgeU
iXwqJJ5Z/k9q3ItH/tig7vElm+ukl5ZS8oKy+GUsGU/PYf/wY29jd9Oy91Nx1emS
+5me718egFVmsWqSJL1xCoEMyQfwobmzuJ+ALC4YC87Br7us1Hw+HBCOMEhBLSzC
SYZY7465AaO5LMGSUmgB6iR8aZi1SPR+E7pRivOm2MPjVAFD1jxmEBpF6KmBYR4l
UNIqsag9YJqMOgETsSRtPYyKXSCnK+QyiURrcr4cX1MT3ogMjAXxFI68FxOm3xvG
4apj9NYMsW70zaFp47WxXLapirt5uwjATZsICytY9FpWtqN4EdqL64f1lye7Qy62
9NBZt9QeEmHUY+CHjaurf4L1Xen9YhvTKyT6rAg72rTqsxMh0bSXe0ZoD9qb4OAn
crtFA0M5uIYWKp6YWI4tMAy2zFwz110urmeXyEohWNxDq478BJiSi3Usq6o9/MbR
8+VpM+0X2BO+4srj7RscH79lAdou2wka7cFzsAXRCSjmVxlzWpQFEsv2/Qnt6oTa
5lo7NF+m7EaCkiaaOYTuSzczi5N5GrSdiaNVe0QMeUBIU009NJlXLGGwHGZbYsDz
0bzfQO9MRs0ZxPMP2svJmG8E1/T/KHoYOjZmhwVTax8aTEbG/X9a505khtx6WsPF
lFtiMxi28jAkbzkmKfjq9r9qIuBMWIkc/94tBboGBF0YgDV2IzCuMhZQ+tbNT+SK
h3KB+CxZCV0PENU0JKL6dfmboLURsFazalCXzOgPtQojsWJmRi08rzYkdVqs0nuk
yEGrJRXhigzrF7S3LKa2TajXc16Hv/+HNa6ARkdgKTmoUmgvu6CKwGvhIseS5T+L
kkIu/7mgpxKJCmBJt8cqNf+8xQ83UbSvqGp7XVLkFVgA+ZtBexvzZ84VGNFLJ/V6
whk+a1WrNQjCtZCihyDxWkbE8a76Tug0YMy/ZG5oJJ4cUvXc791E7GZacV4BKAKF
3Gbqq8AkBCyg8dv4um6Ouiv+2QN6VFzB95kPJ9nJsdDjtLmboYnn4aRfUKTLrr26
jQ4BuU4JQ3cuK2AQRTn+QlWkwiPLRxnwWy85nwlqmBS+3rjmzQYo3c6ioX199HPg
4M30/6YVKMx+7tDBn1ZZ1sWSHE8zS6mWhWQnjJoLYJk1wB/NieqUgJk6MLKjR5Vr
/Aq80ZRiCMb/4/+X6GMH4sGct4jjeJR1o8pnietz8I7hHBJj61cHCm2Ow8u1dQIO
doEyWfie23SF70qIy8rct2JQan0GZCRrUTjiRV8P8SffqPlbb1T2x6mWbu1kjgYw
NcqfU8+7ALDsQRsyCAiKXWKcuKhZoH7S/fSt8/f9nTGWzWpBxKqgZxh+WWerrUMu
Ijtnpl4EM9YX2yqEZ1sUkaydaXMzwEzImXb5nruJpw8nymZ3peB2dKqiXO5Wgnj8
siJ5IQK3P+zeq6rIip4RhLCaW/vOap85GlwPlLIt6C2lZmyVtmHBg7nyAE3Zg9QK
MJ5W5RSd/V4gVYwM8IzrEz5cEwDJ/sC4m37KsI3DSkhkKIyEUObh0gcRZL1TRWBG
eQOA+ybB5rJe+3HUTSqQ+tgCDFxT+4y0YZfnWXHMd2+L15xRDuRBcauvEktaUr+M
YA5htdL3kOazDnzBIkW7RHmK3SCtLAQoQlopMVqIkw4B2DyafrnwF9UyMH9Cc1Gy
XxksijJagTHtYsozVab5hk/GkBFknOwy1kiJvSNgkq17px0J4jPMA2O7shn9etNe
CIZMRkM9eSftYITyUwvlyyNs9Zef6usb9SwkatQ5oWSu+99tEoaqJ2eBPiSeCLyk
yQloHFUuXRyNtTWybXnQJpSsmfCkeovxywqS0juioNKvayxY1ZZUkFKNNmXZq32b
BzOp6m6bZ/eUtZLx8Kc3ZE3C/VdXON/iYF5hs+m8xmwAkJpf1N93IehBQcdBMgW4
MmBHPDFZCoLkCe4AFlD3kcAeNsF8Qe6y9G3//v8rSCk=
`protect END_PROTECTED
