`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkfxmExcpZTgpiA5Vo13QPN9gKwrZnBoMMV1bJIGAr1Sf
PKVAjfArjYzHmR8klWqsIfjHKmHXyx/YGDxWKSSwN5/2OZHq3O8Ua9hjJJboAd0f
m95dHItwiaVAWOX1+itSKp1Gt6bBY1jM8SU1CXH+aDyqhxNYmxZS9LG1x7kAMwDX
mFsUw0hESrBDhZ6sY16UMHFCB8fJ9tw9C9C/a0BkPNbdYrT7duovCxjf714wVsx9
TnV25zfPxgbblHJaABrPzOk93017d7nl02AxPim0k8v1KVJl6QHux7xhDYm0OjJN
0KfZ00Ce8qUXWoIylHoY6XdVEFhAYoml7bgqeVzZodA=
`protect END_PROTECTED
