`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
vwNbtE6ylh3CX60OkOIhF1ou5YCwbiXZ1lUSxNIPawb5xtMPCI5k4ZXwfYfh990Q
wyB7/LNF1gfCkVuoBAKefGEy5L5T7AcNQQju9x9wWsJ2ESyNGRA739w8w6Fh9Dlc
Zpqi192OBbGwsZMiK0XQHM55n4Rfn8OQW/JKp8zs+FQ=
`protect END_PROTECTED
