`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEm7yj/0oLkQoZ/MQxEi9LvCvnYhGXJqEfHBiUWWxQK4
FGRTfedgUh1JZ39xLbLPKWKWNTo/dkL4GX+KBc5RSZV5P2u/TyeGNVQ3VEyr/kC1
9ltjsoNtO+aMMV031a4+eoS9UdxweTSX4jFixaygyYJLpx0qRGNqxA5XM131ukTi
pn/6i02wqBnxWyYqKYzcmNm6Pa6/KNRtQJpMxB0Vv7tKCMu0Vq1pVuP9jiLhktIm
yK931TqKawJkWn4RBG99jAREYa0B68kud0eu3f7uikrSfTVnwHyfOzEtD8FkIwDT
ewsPqXwRKQoDt2j5goAaVQhOMxWkJMqhAsOa4Km5POOJ0fjsParUQu1Gv1EFI0+H
8M0bZNubdPQQV+mRSUdgTv7g/VX5JQN+7GahLnjWPMdFjjx7146wQruTMTZoUfml
vxYpRAirMsIcI+E29f63wIGZMclV69FI4AcOOtuT9c4Wxt8uohCzbkTYwvzLjPa0
M1I5G19QQrp1nCg71q3BG+2rIo4HJJtVi0yZy7iadF5bNHK2rXA476Tgeb4n+K+k
8GPQL7Sl/9l1AMJRqZTpQ4DNIh4rnQNUGw/19fQ/cove1PpwbmRYreBnWSl9s3kW
`protect END_PROTECTED
