`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLayf+4xVYOkrOalMDh7v9lREDzs4J/A5X0b5nPH2U3K
9vgrqSR8pwy+iZ20jtEpL/5pK/dY5g1slzdWId28keM9GTwcZuFpbogXsVmpvThK
dhv8ct0lPD6ssWiYGW2Aw16CnNGec7bsB8i+f6maPzrxEd3kF4bUj9ym7/1VvqDp
KiWCyESoNKzswfAn5NjlyOnhGsiaWeywTTVMI8fQofoMrQUEbNx8aIPrF24V7NAq
boSMOcs75Dn3smSr0mgXNM4aty+OZ+7V1D321veZ8JLxNvcQICBuEK/hvTmJ0zMF
pxwKINaA39WlHhClZdTQRA==
`protect END_PROTECTED
