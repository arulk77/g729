`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49W0JskvLT4QyJH7PJ+JWXadNeL+UEPZiYNPkAfeJTxo
Df2BHKjkSRHjyEN63pAiDNprIXinybmGpquBJLDuJGgndy0/EEvjltGsxrZjGOUB
0uU2tknyHuOeH+EPqz8dSGIZh4Kv/NkIbZn7J9YViXls0QKkHl8+E9R8tZXBSIVL
LPa1yLUPBOPaq8wlEl83slCRYzl5XLy6OVlOxr63EiO5ZlXzAEH+5wh6l+ukN35f
mwfhHSx41qvEt/ZZlSRthdFdgY5mWjdYwh89olofqUO2nEynUHe9OrwII/Q2dMcx
jKvpmshEOc7bJbOikKePKqA88VxzJZsr9IrMmbohjF3uSk/3x8up2ZwE4BkMyGna
n9+JLDuROdk1f0VW7GlKhA==
`protect END_PROTECTED
