`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHtG1AaSI0YMrvAiwuddejae8RviP+qSWW8KMqjh94a5
EsARMsshJG1HjsGeZcheei77FLii07FbD01Ntqnh9kFWvnKMfo7f/JOFUeNHuw6Z
GkHSW5DOLR8CnYkCqbhxPLSJq4ftWZaV0XEZUAnPQrKGTNh/+Otl9HtnJox3DWsr
coYQjNhH0GP1MdWfPRmw83Ov37HukkOUtX5yzWKCcLBH0ACa21/5RRzS3nwoUe/y
zMJNa1G5RoJ/Qb/Hp3GC4TxkK1dV0twhTTLGREc+Kt8TKGVcJ/XQBbWyY9T91S8J
brY9go0mZ2R0ppdOeoDIOMAIBuYm0D7gSAvz5Scx4T8WeOHEKyLjRnV5EuCcWfFL
5P2wSETS3vdqBLBByUzohEyFHbQgZhCeq2qWLPSImlaZdV9j797QvGfjfIq4tNdp
`protect END_PROTECTED
