`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45QzTmOLYC8HQDx81TXDoQMzfwWR1cVHajiOfiRlthTh
ET62dmjoBNzAzNKnFjMdBKhniOpGODGXnhyNKT4r1HXWReL2AGh5OPFwn5VhVOL4
rwyW8GLNnvDYDOgnjIhHROyWpSNkkIv3LRk2UzOhbLwSW6HmzR4sPlFwUZFCklz+
pSNdouIJE5GzhjBJfDJghJVySe6lf1k9chpwA3xjCmrxCdRoNT9xE8YHDpfBLUQV
wIdRuoteOdBvf6qMH/xM2Md0u73b0NM5Fja08d3bZ9sjQekNYUsIKmzPv4VHdzzi
uKAuSCMPPkiNtsnmQxYVXQ==
`protect END_PROTECTED
