`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
EyPZQug7Dj6ZZOpTpHyGfijLDEVoaoFKIGR/Emn2aqh1iwdfmMYyWoUin+HwzvJy
tYuL3wcMuBXmrvX4sZXMkQ8TDAYG72dCd+KXWWtgYmVIIwvqTH96fwgdZmeVxSfj
OSxmreiv8gUtJ7bL3JbouQQ8bXbfdcFJnYqWVf6/H9SmLtCWpN/QJisPs1Fa6U32
IN6a80kf/1199swdUE9//dmhlQ0VC0bmFt8LIAg5O+4XQEZnwqqYViQ9TkymIv9u
MVbeUTfnOTp/boaMwKFq3nde2RSjdgMFsgGY5Ah5VVKiOdexqCa2Xps7U91d4bCv
tPcIUfo5CXz/FK8Qeza4WvtkkBO3eU3vklHwrRN5LFs=
`protect END_PROTECTED
