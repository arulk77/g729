`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
jnh3tNoF83pwuVQMfI/BYsLGapprzJsT33YHWZFIC8w9CKErQGWK6YlCJPO6VrcX
1etiHXfvg8tUAYvFT/Bujzf1orAbrXlRTdpSutcnS2GnS5CnyCvRQmhmaReYWMhJ
0QuFzANFSfdNx4KM9HPLSggZNoJtcyBvGTDd//sUGv7IzXuhalWy8P3RxbxFyW9F
8wgmOa1Q0LNlfctYZhtfq31YWcsMWrKPyPeImJWWsfKRvfr3dFNiwhkBFfFOz/96
gKzzeSlcQzsdumhwYEvWQIWbbVYfY31leIQjc0v5F5QaFvaVoMx2TI3HHwsBcQOM
onDNwJwoo/oCVuUG3YZHrMDC6xB3JxV+oKL7t4NFvCyrQ/lyJcp/1/rdYHQZE8S/
tO4NI/c5CN6hNElGOXfrRq5lrq3CUarOuHhdPTfQ78vxFNJxKFc1T8qyVO+pCJw8
BSEoLOP6PUKDOILAWOGXMzYMnB1ce7ozcmPg6/thUQJ3L7Gk77FNxpu9woO+opQu
mYXV4qr3+Pi6bSMFyx8As64B8eCZmp1XCjMZTVXsEw3dTzJwMMsxTLy3CsT77aF8
FM+okjWybZ5MM8pj17nke1KFM/RudkaX6mhW8171gHozBBzGfa/Z0B5+UWiKOLmd
WzTZw95W/7LZeZY1pJxaSp36NAPRiEypPXCnor73jp5TPEXIKl0Krh9AzN12/bZR
YDFg5ymyunUiaYGGQIDOvz5WF4oe30ieuFqo+szRDdyoDthBLMIoEZ5MM3m86khs
3u8URRjn4eWCvm7ghaICRngCMCTaDHeSbkLqI47S10cxxlBprK0H3oiZ5dOSjjS9
RM5rqmYkSroyXHMtD+9ePsMUVn6CmjwkBqy3tQrRkUrK4mYe+jyhXL2xIXxQyRXP
4jwFR3yaC8hGeCaT+1vyKxItwYWkOYsnnxSkjJUOYOfT2l1GKyPgUaS7ThBB3+Ag
z53Ppkpb2bEtzRs0LPfRseMd0hGqZ34MEG230S5ZiWDF9L2AJbsjokkm27xcozrw
uJnVsydgWX1klp+pW8sM/1BOQ3O++C8j+e641qW0+zccaeWM1+fN5MOjJYUgIGel
Nz8rWk/KnnHZBDHp5UjCkEr2sNmr4V7iK59Z0ArSw8JxapWCFxU7aCTh1qWtPvAS
6Aj9h04tHz4/CyJ9+K8zSJ1TWBA4IMpC7v6bGaMARXVMgRKoMfLsVdJeTMBUEHqK
rQjHmL5nUL/AXUbV9SMhCsXoWPh0HcaIJG1hslGehJheO2r1XfJP/JKdnZKAquYq
y63DrIz/z1U8vpZ6L6sk1GRBw5ZJQp8L6TJrqdC9DbkOvcaF4YdtOtRIpeNKL1da
reoxqnQSNE93irOPIMW40wlIyfXWyVEN4KUx2IKw7GVKB5lymwU+kehZEXBrunwf
f5ydg7LmSKEU5pTvdCeIqdJ0ANwX8TJWfA4IgqCja/buaPAuphxJW8YEw70CtdvI
6W+hH0LdDD7jXqaHAdHgZBBxWRPAa3EiNJK26G/o+2+6elscT8uNOgytsLJPckzf
Od11dza+7zZfZYo9XkCCujIcxuo9pGErpEVDYngHimx7XXvyV2A1IwZFhaWE444s
HFq+FhSlrUOVOTSF0k+7me2tmRFJyTb0c/xaNB3J/qyj2yoC7Cs8Q0b8c2opIuCk
eKSdhW+vM/ygKPeucxjIILwRyWEVXKIehBjN1IrVU6ppiSNDyVtDlVZAw8VQ2V1u
0lNwSFZcE4rsSb/aVNIx9/+7oBfjMAQElXDP3kPsFw8FoNqwyh06Mw1swW1Wdmkj
KPxWRSO4fCVGaUoxvNAN8bMUUBTbSNTzNC2d2R4/t7JTOSJA+ZhsbsIHtNw/UwwP
nZHWgnBLTEwQisDnX/J0SLBjHF/wRcuU2InzNa1bpoApzebJDB/rLt98Pu8i1Lrq
cHgy/ZIYhhgGxoHoiBC3o1dE5EE5OR6FpTItQfOzEAShBgZZSt4mjPTEYUnBwxiE
TGtB4r+eNQ0hFHFwSbNRx26IMUFpnsEEJ9SkXZJ8sC1mZeaaSVHA2qLOoOjiGpPv
HjmfoyK1AvL2oC3e0AsQNvTVX7Q3saOB39CxOTeI5chIsSK5hH96vx8iFngL0dAK
5ZV69/SzrwYll8WFU2X4ie0+dT7jiLZozQJy8dxIxEMu/lqVoAIq8wQl6hteAg/5
N4NfphyxMsEmq1ZME14gpVbGEZYPbF/7+aSJUwP60oPsRhozxR6rqM2IA3l1amvG
9N8erwnjVbQIlEa2+o1OYD+zZq/v33pJ8X6JfiTnqUUv7n4KXoEMKnUbdt1/zuzT
RExZG62DJ0TSMnnqMNoPdLStPqM+4F2Dw1I/111x8E+jZCQrPL+IPxLRMvQDPYAl
G/5ubGmESlmWnGGafXY3C3S+AHa4kExUIZXnndALXFFvQw1Qdn0YZp7gp9FUG6D9
`protect END_PROTECTED
