`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
KEyilwfJAC/DYCM+BmbmGFPuItf6UPbQQ7o9CWKaQfHjzuFW/zLPZDgu/+YrbwOB
anxx3uIV8w3F6MPlmVMqATti0K5ybx2a5/QE2Z6D5kepwwp7Zim7kDCNWK4AKVFP
jtPqKh0E/qa2BhG2FiNdnggm4YCwGoPIGd8pe1v1CDfbmBiCNNbVKmtw2YHGLj9K
N1bYJGbVbeZ7U6b6iYC/92PHj8ML8ob7ceaYwoZSN6eGFJcrhr1GnBJi7TwiZuG+
4BPmhHBzyXMq5kiXRom44WWILl7BBDFDwLXq2Ng7+trlpC+1+SOiv9PVaLE2MuCj
sAVZj+SpVLlW5mWCsp5x1hvSTF4ArZJXWL5STan3sm8=
`protect END_PROTECTED
