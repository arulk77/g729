`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Mu8H3B1HOKUkhEbf0nZXIbvdsqYJ5Kki+COsPLuhrswk4Fyw38sKfWHNVNAlh/Gb
L+DEVSN/4sfM5oLLF55jhV2z2LZ391zmxGwBHLF4MW/h5Pb128vqgD8NcmPBuRZ/
A08ct7qdspZCX6A+pXe1ryiWFqLqq+6jbmJrmleXyryU/aFI0wRIMBcJ7IAq6728
fB6wZHMOFa+AlJCQAyCc8DUdcA27e8qAeJG96zukmVQLakERR4PI7R41yCrODQOx
oiqyXhdHKwWBMO12Le6rt2ZBQ8VCRq+qbtUTcnyN6JE=
`protect END_PROTECTED
