`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMxGdebrSOm4iXSv2RACdh+JYhOl4BgQyger1Zgl0LYD
1yS08522qid3zPSM1PT7dXl4wowlaZ+QO3vuXOgF+b3gYbX4bUyVXoSSPaWFomx8
rn4ekXD/Z86uyisiTg4Y1Vn/lSC/4Z965TverCpxVfDKRf7bVRPhMwD7VbsxfFjL
P1quWcnXdJ/k8ksP/UF409ZJDHKTP1/dCchr766CpuX85hXsmo2RnSeRxk9Lg03O
`protect END_PROTECTED
