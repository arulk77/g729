`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLORW4tKTDUI2mchUQnoK3IDRNUPUNF42+/bHkUpAeNF
e/gzCJw/6O9ksdUcCQBd0zRcK/YZprLo8yGlOx/fLEMeET9cMiOWAFpbyQ2MKYa8
1zAWU17FcwFDg2f3uoZLZPWYdHedaOEoMksdRbOpARGFNLqUb5XV7j6m2MpEjnLF
`protect END_PROTECTED
