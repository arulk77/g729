`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
uPqSyrWgefpEQvcKB81tTxthXVKl8iaO+5eSXd1/VeVf9te70vbW6EM+oMyqv8Kw
ptRjbMjDq3Y6XwaFxRFk4va788ZlzbSrBz03bxeRbAhNAJGHTtbJ1ki0Pm90qmRd
gF0sgRycSyVGlb0bIAYBGzSf2rSGvCCFcWeEgGRQchnoHTp3n+SPZUgDlwP1aXGM
0UxpR3PhZBNzQmOMlPuf+D6dWNFWsRQKyzkW4T+Xqvg3zrBnRsguoMcUvNq+oRJ3
5BujjU1s+sF+mr7k8I66HC9Wh3MqotP3ku6Od6SJ7uo=
`protect END_PROTECTED
