`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF6K+ubwj1D5Q+t0DXyWrUeB9fdUiC/rSgJV+4Fkufav
u9TUBDfXS7D7aspdyVJHGTJ0+RWctJVqHDBLt96PuRuPWOehlnBS6b2vHBOgK3dJ
bz2vyIoq4QlD1gY7x+U2mvCqgWgjO4wZG+8OYKO3siZStV5sMpxZIzxWG1Nc0Jyl
de3ptLKWIUNh/Kd80mLnx2/0O/fGbENd4dXwKjlvp7IHYMiDBAUyQdLVPQT0GVXd
`protect END_PROTECTED
