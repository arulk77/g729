`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCvnBKA9hRFqiR2yMOYEt0CqlDtTjxmCEZ+NAR0071jv
fKAIyBOEE+yi2/qPLr789GfinTdJgbIamW15jwJG79AQiG8a2glgMawgxL4mqHUN
EzMPn3Eap4WtGFL+BQOZ+y2XJIZseBCnG/kezpbdKwgkxA2E6pKJZ5vvyqYknJex
4cLv1kJ+ZuBnH8JY8d3mNtNU6VMiMR+04oBWUjlgMEHvGtyyoeRnr2vvlA98XDU3
FJ9mnRI9aQ4RM7uJiCjL3VPwiOVwxr+O/uXMAQZ5SgQ+I5MyFUWDcfPmG5xN25g0
uaGhUu0wsYFDX7VWv3WQtNzi63wocK5dcnJJqHScuorYYl1eZLxm+5bn3jvhrT9F
aJ3HP8rcx0zKkzHsxcxETt6zPExZ/CkPdFW3gi25/sR7iL7TwpIBdw5vCXh9h+wU
kWf4SaATyKpEAj9K0FsUqzeY7aLjvjC/Z4jNZdoHphEHsFWP+vaNMkTH3WkYa4xE
Y/rJINz2dnxNDvI8Hqh6KSwneYluZpLWxnB/v2PVhbHIjYvlbhldvS+TzfHKIDmS
`protect END_PROTECTED
