`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mkkYvnTv1R4Ho8ntydXMxq99Fu3PIE0Xaqctat92ljO3oVJAZPs9s9EQ48w7Zke9
eWOvwLHDfogH2KsQ4hq8+Z0YzBbsdmJCCCqgn1fhV57Ai1a5CGHcXZOobelzBF5p
VsmCf3mRrKERqFm9pJTfsRNDYh0OjJA3OrhkLw8fDyxX7TCRscW1n9lyiX/oM3pC
HoRjkB6jJacM7Zlk+Af4A0PWYrsFu3UjHi+bkJh1qUx/arYI/vfy8t39PdXXjw3U
Dmmnl9Td/DjGO2s2tIvRr9mxq1jPKGCTfc2ay3Ti05Saqbl0FoubLeIjOaShkjPl
5j4U2FTquGd9FqV5CvFnKUdUqIkhZqE+/aRrp+NxDcFDL/gQS5bLorOyZiXGXF8l
pFz/X58+7ncotciTy9w/lGXIy9RkU8Nfvlng2i2cOxs=
`protect END_PROTECTED
