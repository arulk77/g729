`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ldo5tR1TIlFkHjabU/imcRjCx34KjG4p+y+q+D/ALdE0QKHe62H0Z8Me8HM3/KVt
gtAxRhZTPI9suusFaYTFbsiKiiQhawZ2W7Z9DKQOPiBFa0P6/hXgkEYyLPhe9qAe
OxN3+/n0fsW4etHs4Li0RYU9Evf4V5dc1/hddtOthdfw9kNooidChgNwXykcbkl+
rJGPAnek0UXkzecaS89mP1lx9Ouk49oUYlTgeVEK1umn3Epgo/vW2wl6E7oXhZXe
KiuPY1Tpe868+1q5S0ZYmOT0mICeCzh2qbXZulTS4dIq26pKv2+RkQ4BVBHNP6/+
ZV4PEm+RHhivyb1iETe4WzBEga7Z7IbNp8UOTNPc19OCVanrxIuHFmfMAUztn6y9
HmZPtYKd4XpFGSkxEW0UhzVl1U2Dc3xZYeKLjGR7LuQ=
`protect END_PROTECTED
