`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEKwXZaKoC9vMd6Qr8vuIRBlK3w2FVihsA9H/eVZfzrk
a2PQrRVsmwCtrSsH9K4kiYJjpuekJ63udbCM8Sdw8812H5iXmNF7H1gP+SI9nbvJ
oZWOkxIbqYQ2NHTyxGUfTj+O7ukfRVru7dTkHpSBxMvDUeZPal1lg/s7TD3SpYba
lctUpXwJdJy2xC/CcfCQmx2OZh0Nkq9O9JvpkyxjPlnCHSi4Jehbo0KL+FCq6n01
qKvj65Vn/6XEi2gvoMlnMdy139XFHWZPJqszA2eksyu/+nm2sLgXfNUf01x7Mnig
D2WsZF/MXCydawra5VB/7yu2wdPnxbGjIbkVi+TcQnwBUdjmsZhy0pd+NykcMTVN
ejQB6HfzHDosxU/GSyVH96wBnNyOQv2RCcP8SkS5uGEOe8CKqhT60OVxUOREoN8K
ICaY899Ish7e5pekotrpno0vlQSk/B4A8DdEVMs23RfBNkDpzSRo/K2PzyeR+Wcn
KG3Wtz9ae8oILHjZnUFFtE1xEO0nK/eg6CUEXwtfGrGGS8YJ/yJZmzEd8vxZrhT6
P3UztPO1fPHnIIVZAUHSH5epvf97QKh1+h8YumzGXxWlJzGnhDEsLsf+E9GDKkEi
`protect END_PROTECTED
