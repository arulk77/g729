`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
g2Y1IHGqrshzeCCayy1dz8W33EHQspKlbV0WG1maOE1wejiUncTjtPpxe4jphgwx
GH21BtlhTEsAoa/JEn4twwmWJSPTsIApB81aogjyPqD/JygEuASbOc8JJfWCpKjz
jjQjf+DOSjjtRQEPKZMu0eJNARNhJ3jWViZm+WNTqvIqE9pUAugscZOIX9t8jjuN
M5W+d9J+mHTYBFjRhuXF8D14ePYMR49Nc0VTN/GnhwxY4koNUiqh+OqRPBBqjQVj
wXpyzpQF4l96PQQNnc2O5ISjv+mbK3IXH6PQPMDsKsA=
`protect END_PROTECTED
