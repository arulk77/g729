`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
DbDGhJIvsuXPlM3LD6bseBKw99u88mXeV2S4GajPUTIntgD2Ak00o9qPGQpu48Ys
Pyy4ZX+inFsnGIriqGbYTF/a1IMc04wcM17Vdi7M1yAXBf8u7PsHVafwP3R4llqg
tvUyqYC1OPXFilUMCZpk25ATIQm8Y4+xN6Y1zidtsBrRPYde9rFf26sJsAL1TS0C
EfON7bBPQobcquQ8HIHjyutWxKzG3F54c6PSPXVvpdGEIDJ04ECEfPrIQuHNMLiS
8Hpff3p8xs34O7jzxfwQD4hUxnPmJOxUSpqH8TVhntKIyZ6kBwl5Ni2ddjLnJDFo
BZegnc+FQzP9Zq0GeEImhM4ZHweCOaKHXET4lO4mrizPj2ABvGnbY/aR6rTfPogU
RSU/Pba72swfpmpjGbcmBixyy8j12a+khYQ4dAbz0EQ=
`protect END_PROTECTED
