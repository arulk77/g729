`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCtlqtjPUZYBzJEsDjNAT8aT8MkCWB6Zu5TqZDdKECfR
oCpiWy3kl5naYwzGaRcY59Mp+kn96xu7DCD0abz8moXduvumCPYFqK5mWkKKDgDr
vE41s8gjgUpINo1TgTv/VmWcfj6G4PNlzoctzYOy+2mOuHnY1XRxj83hx5Xlj7Ip
dtf4mut1QAUW0VHGwvkf5FWkWPSnebjVdymOujOrDFGgSfEphkSPxHK7IWzevVTh
Zl8YF4+qNRdZ43cs4145tg==
`protect END_PROTECTED
