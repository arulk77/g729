`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIgqFTyGoFoN/8DSv4ya0lE7pgVYOxkd1A9Xv8jzMmPZ
bORyl0SFgEiVRjElvN15et2XVvhzxhoAHGLiqeN6LIKVcLuy6E4p15yUkrEVhT9g
wNZe62Royo9m9LaMAdYWooLlm9hu/8QB7HDNgW0wg64HG+TmL37Ux5eepOgAxrFk
W31k0f6VHCrV3q1dWiKBQo7Vw4KQMXTqCaFlmFxnMetJv1bu455bgGALyh8rW6ff
H6q1yxqCisVIQjmh5eShMx9D93nOQidzVg4wg8C+ZbgeJVe1uhAalSiQS3Qhqya5
Lng9aRJEpz3buaC3kSa0A46uLKcj6XFr3Uvbl8WmnoWdVzv0XVm5P9B0zBV/8nDP
WD7R81TWI23nAisy0h9a9A==
`protect END_PROTECTED
