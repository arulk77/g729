`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Wnec8np5wbF+4zwQNycFkIjWYpOVfgE9d3PXHdO7ru++egwVW499+QGdV55Qg40g
kh7m9FrGrdzeR60MVhHSYU+Rgr/nlz4lcyWb5wHFNZXP0GDfRtz3/w7LQ1lV0ToU
Bwb8R2ldJMWd0cv+tsRMgQAxhyE3AYhu5QrnK9olWcWq0bCMyH9s6Hx5q/I4XfOw
eNPmt+dkSzfxlXKzbSA8yNPu+DwX0GcL9R5xo4q/up4qOIb8GkoCSxCYonGuPBTT
sP4jU88Thq7PTVSvo7Fnzis3YXnN6Dx126vP/hgTcuI=
`protect END_PROTECTED
