`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNxRg0Wx9RPhyTj2eH4avUCMfHvmxOOJ0GWcBENOI9w3p
QQ1TkOV+jFt3y1NA38bQWvFlxFGyoqOvrhz0yXgNE183iamQdFosd26lGreTVUUs
COBRIWmkZ2MlqfIpRNTCvRygMFfAS3ulPq8Uco9EHyloaivboLN2Qn1/prh9qiVm
IKc41LapZxnvOhZT1DQ8XgiN36qlTceOHrqmSF7bsJfR5vUD6Qg048oF7jTSH+/7
JV2GT4BRfeDoC/tZpSqYE48TfrqA/SOvGDYefwvyKrIjrbln6YDkaFAGwjgCvvDg
9zHSuQtBNigxygIo8az+OQ==
`protect END_PROTECTED
