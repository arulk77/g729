`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLl5U55vURzwuT+8vJnE5/1/+uJP3pXAHLapRrEQkXk+
UbumVuldesgYwerS2gUHl0I1gZMWLsdb2ZKNVkrar/KhNge5+xcqHKyI6ZS2QQzN
3PeJftxTZKmSsQeHzk8UHQsM/JRQmHaib4AkC1NkOyEX6xbRskgrFFk344SxZNPw
eflWrH/itqNRHKaNt8F6LYzZOe+Z2hTg988q8iTiumopNL7tDO6oVJrg76iRlkfA
N+ga54pjcXOCD9hTEbkdB339mUo1N+Eb8JPMEXEw9pWW3b1U+sqIP5T8sTcqq71C
Roeq7gRfPX+tpdCPqVUY4Ae/mGrv3W6Yw54WdVn3pXW+NIv5FurJX4jE1IDM3k+8
6TzbiVwM9JhGpJJbSmelxj/GH1S+JJV2UO5d8e8J4eIvvkLWVkL7xfVFgLWLRo9j
GCxEeTMJmucjpSfDqZE1hF0lmGQyvyAxLpwQxuSZ2daOVmydejm1GlbR9KIAd9Su
/89CkT0BzBYdu0TI+2+nh1GEkR8ABPpBf41diOvHDpVTk7WGXxl+5VRCI21KQfsF
`protect END_PROTECTED
