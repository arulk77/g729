`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDASVYgW6kVbq8/TzE7W5yRtsZUQ6dgzgYzz7xYMBLVtF/
vyEzzRHGEoi1Tb30VvuO4yNR9DbxxADM+fsagoMbvB09f+PzhhTgdx8WJCmlEHQx
fYY/45HIdjATKZiJfGxsi/7M40X1eZ+c6Q+BFsoMnq+xS/6d7DG2rgMHDLf+JhB5
R75MgFBsOwcFnQA1/ekuKh4vefWL6zjfePhxE7aPHs9X7JHWvEk6egvnmoHoUaD7
y+sbayYSl/oJcI5omD2SDJx20bxDF+0yX3Luz3YUNKIgAHBr1AEwIET2U8WEgG8F
j5J9y1pzI5DmLksIdQJZZeQ+QwxK7jxFnBNFLeog97xCNLy1VcTJfrEyBUfLH10L
Gh//E3Ob/3hKzkFcpKoHMzkV6cEKNQA2iYhtXxUaHxOS79iEXuoM1NOmcFcRIa17
N8sXmD+JO1Kii6PtUwP55jXl7GvE6sYJ9qcVy+JJb/WC9Lf/w8JVj1CC3ghM/5xE
Z+SD0kjf69WVj/wJN4U5+bpMXXj8ND+WEWunQB302uF1MattNvFkKnDCmnoAs1nH
eWB7vPZkguCIYckcaDdPrD/mMXFigfjMvvI0Zt8INNaqztopLEScc+ShuWUK8bnn
1h7vknXYjXyOFh7MzODgYmAnpxTXv/2AHdv6cE7MLMEfkPM6LveeniWEFdSkkRdW
iFHuO72tJUZx69YT/7M9eCH60qalvSqYWvJjxBrw/FtFKVe77/1Osx39XvO0/9jQ
HmMWdqSCDXlz2qDXZbkK4JudDJI1hfgYkp1S/4/+wEAgo/KAiszAh+lbigqu1rUD
/s41tmvSJa1hSW4dsgeWXecMlWzZpvLKgpM4lhhXXp/6Y0vHqOYx6iyAlHaRJMXp
O2w2bfSc1CuC0g/bp/WQyYSnW+5je3l4QgPt2XA0682yZs4hf2ohJEE/fvYzpam2
xiXxDHpHdsFdm1ExPLb7B1xpmFUlNg+zl9yJ5pzJlAkxys5Feb0nSdut5/K3ygvN
j6d71NLKehWUSjpKfdz6HKm0R44Z39aLBe9jnPKQ/wMyoY0Q3JhQ3mo7N4VaRQ/W
VjOGMzzoJF5yiZknwbiiM4xJ21UIagCoFiGt/iG83ZxtjvbGWGAml0SnVVww4nCO
IaP4gaVvFjQzRWOVJBb6qR0OY7V51GMhWci1AExiTX3KdLF8Ba7eRiBVRf7D3PdB
74+p1ETmGVjNOtAPRBlKzmKtHqGm+MqbYK0cyVnBKQVdoajxQVSEgZoauj+UiZY1
Pu0LrKXWNHep5d55L9p+wBCwJJGI3b4JNLyqBTl47fEravzeyFZ4fTWOZTlG28la
MgEQlIO47qIDgnjd6pr0/vmXRqUo8KivSkO49bDLhj5VL2ZMfWzPW9pJ0V6pJdiB
kXup3BpcoDjzlT5Sh9QGKlLeQKTl0KL7cBrM0CXqJ8EkkTl/f1xKRhpokHMEaaB1
ZUfvnp9XOutqkY0TwkazppPeOUq5PlJ0Q9kQ7XIdGT1vbwxJV4UCUvD7Kfan0XH4
y6GdtrGzNcuwReLHOLzK67cnZ4sSnlk/cbqljYh59ClJcQb+pTzW+OuO8HIpa9+i
rm4ilAI0JYXICX4Nefj8N+Qj5OjqiMQ9VcYp3xLGg3r5LX0oO7FPrbpULvDRgP+R
nHqeUxsukxASd78X4I4S++asq8IQLWEBXvU5LSSGe55fzLTmjZ6gJU3tEQeRJeeB
gpTq5UXTwR/D0IPYlIo0n3gh8AeDG5tsGn6FGgb1MxjT4l0Iv1dPZ7gmTSK4tIL3
x+U9EehZJxZPSbsHQK4u1ZeJR4CUC8HBUqEwdEnnj1EFN0m9FE5A40qO99UYXo0C
aQUV4y/IpL6hhb8NkdJvQwpiq4WnkmlXgrFSSCoQIGFtx7zTEX21Nmp6KX//CD6Y
zxK91E0pLPE4FWYZZh2i+FmRGHl60Uk82F084VBMdk91XF1NOqcw9NihkWMLv7XC
VdpgqROY9gn559Dy3e7g+R557UZ1xqSz6z9lDzktW37nw6YXufClRTIarl0VqUi3
5q359NV1vwG93TSJ91UvASpPvUEt6i9B7Ip6RjjBKvnVRVJa7rWO6rSIdBjBQnwF
Ho84o2138WBoFDF/UF0HT+P9Jkdoef1lxCHf3MO6UjnSlEsDfMZrxP5+/iSQKOyh
hVwzKxogw2MS8q4uZ3I0O/cyyZD6vCJdHI5SysshSTRnvDZJh44dZlGhZqSh4hoZ
fff1Pl2/UMSW1KuS8dALk5kEjxbbp4v37l6BhG+OC/9NXgRJZnkkFvKbJpYJ4RA0
ggUXW7DkmjHAAqjN/wUuonA6lvRaiGlqSMCiIELTmSgtq02ywAVvlt2JtGES42dv
20VEJ0GOdcbkHP9V4zZYSv5tc6yQvoUozZbd2cjkSTXOdeJ1X689qC4Kz3VFTZhf
dnlRMCBq0Vwg0rt/VpON5fG0MG1Ou7Z2VndEE6JJPZ3n2O2psdXIjw8lRlIYw7Gw
xMNB71rCQJrT8VsneKHGWOG8kpLX8RRlxdnIh8Ri0H4K0QRmTnDggJc/qFNC+mPa
7tsUbYQVIySALnsHa4BLQvMJYvSfNfGpowNCq8mWPN6968EsCMk7Ce4xYb5wMvJz
/kgSG5imVeP9nW0s6aM5bHlKc7unOC3/VXxc7vOv6LGfY2xyEZ/734GNSwBrsM0q
2S9+4sSubaYv44kRqQayoHjSMx28MdY7L4V7p8CdDFRIMMBnb1XzLMVLXRXis2Hw
pXmvw9UqXvi04BV8D/oib4WZcaWgl+zitvwXfxQIU21G+gAmcWvA/9tO70KOurOs
Up52xFvpopGyp+XT02u/L9eY5BUSyw76g/mCDusAqq/8MIqlOpaJJB9WGy12+u6O
KW9vcfuOM/rWoVWHe51oBggc2M990Cg4eVhmDwf+nXlxdE0Ang0faiyitwGr2ILs
KDCIEgzYTOeTQaWmDwqcJ0NJHEQ6fO/GafvfIx1IgDBVU6ToEE7QosWKO9avW/tW
uICQLGNz+tKOd/avqlJpxaqMRGJ3tWis3ufusd++btXB5ms8Kb9lUGSkqlsIkwzb
Fiup+5yTjTGLDwwc1szR1Mz2CRbofHG6QqOmqhzEwsJsaLy+E7TjPpECFVz97ptN
BzQVy/WkqpYWKWSRvYMnTjFksaEFwVNRFo7cUdAw7rq1tbHZ+2u87S0jlEesbzJ6
5dIzdcOqXECQgeadFpwmhDVLs5KXjwWUCzy12KxTi6NiYGcSCvH9n85qK2szwAAg
DZ0p13IiOah8Qm8YKp3DHP8vt9731MBnWmkVb+UW61j296e9Xow4OZg83VWRc6h9
5pzGvhDebgdI+4TrxAOv3SMMRWJ3HmA6PiUS4qkXzI+LhIMRdlMxx9JJdmb/DSqK
Lm9Nw/3gCfJX4Llk9nc9OtSiyhF77tINH3/FfQ90xyFKZ04+HkeY2rnseCyEQVRU
JWEqPJ52xxp/hQBshBDo7XLWEMImQOzQI8V1piR8g3qhwsnNr/s8blx2fYi4XeEt
C1leD60s4O+9hT2ECmeSvweSkA/7Twnjc68qrSkoruEGvL6jYZQznHf0pUj/dTOG
TjRVfIRr7O/ueV8RWEq22Z+FVg7ch04w+Cz9cbu3R6F+IiNCNKsYRL3D258FFRTo
0sngtmXDkFxzj3ENzF4Bi5qH/61AcNEiAGr8CdHDonluaNabZwJNcDlw06x77ZGO
Njs+BmL2FHemjgms2uMy/uF749FzNf3SnVsr+3BrVaSiP61LbkKshLndytmJXh7M
6j1wCHmelm/UEzpS/6ru+ZLQps2TDmQzk4NEytJrcuHQAZyTBAssqcGbU5UAzekv
B7D3j8L+g8fmb2LlRcRuRIpqkuroU8z16o3cHNoCmLsJaNtV9RPPEl1c+qGrIuKE
WLNWys4wMdXKswzSZpZln0mehFylUpRorXexNTaK0jb20ghywO/xFWw0j934pLj0
2nYnI1Rkw88FAzfSKR6MnbkuhCdpcJRSiLFQH7LwY4KDq4b/J4ns1QTIZ7ivwm5o
Bj6Mb/MvwvTHhYhpUgEReL0wvyEAkibFHPBsWIhldgQm3yozPB0vph4zCINy+pmd
GujF9LgMHTkmbSiamIUN/cxvTU5K0Cim1M0x2R9gtoKgg30JJTHuwOsXax5rTRW9
mKy+8QZnKrQ3+HPL2Cy5zp8ehlyQ1DIQaLzaM+fJ+QXbgiUcuz8rnhLH+mxFToIx
Ree1/NDpVCTkgRWrDgPZnbrVU8Q84RAohyIXHn/TBReRdsJifdnw4EQPMSf6e8eb
cLyyv10RhlXGzg4gRqU9eR4HZ7n/OKNITQiZN3ikQCRnOlXDaL7jEj850oRXYkvI
418EUJi/Xlw5PSMLjr8x5PxOJowZjhbKTdb2okH0sarcCwTSwhGbuYAdyFOUgVpt
LtD1t0hsT2hMwP0I2Dnjr4/LQD2meYw7bVPnPSkLD7gW0zcviZU7W5/uiKM5N+ua
l7hAD5fQgR29aBhq6tCxMn/1kGI/42hJh5IQ9NQGTNr6cH6v2W9S/JOiw3jSLn6U
84jMqaFWuVhqJYCwaUN7pC76qmX+A8j1SIYaNukSCVTpAx8uLpHTlF5BsZfxCzoi
DYQxmL+lDbOPQdzDg4LzavVxP4ha+4XZccMMGe+VpKcp7PUQaZVbbSHu51PYiRe4
9bxus9RNdpUJ2jN8XDOIJUaJoRwdUibL63VGUfCVr2/s5SbD0/yLJkIUmfBWueK0
wubq66e3djXkNhLG2vVg18A79WetnhSl9JRLDeWh6FN1HLmTvuiGp2bG2UgQncLc
aeSQnGYc7Fz2b/rNylRF6VjQ8J7HSz7WI7qkcYOr0WrX6cv6Ulwxbt8xWVIou3tj
PxxpxxZXzMwGZkT99sZTdmlAB88A33KtmPN/du+BeHry8X6Pzqy/Sc8STn0nBJby
WX+RaaSRBiK0epv04N2UdLg3+E1JqiaeiabBVnYQE8MvTtzmO9ka2JkbewMWcv5H
do4WmJ3VAnvvi8p5eDQN6xKuFa7QOn7H6K6YAtGH0iO13+JIJdGTttpJnIdYFqlH
iPym/vYUetPHMJpQ99wvGoKo+WQyMC25W3MPfElAqObPgagK2tkwyTpcEOL8ZQU5
LD379bh8f84Of38BJ03ESz01uldKknMYFgWjVAtbThOLOzlJM30+Uxr4pVUn02gb
0CN9iXmR0kZB0WBORLvTuDG4Ey06ll6qROTJvtzJYvX+BR0of4bug92fCmZ1LyRK
/Baw+wytJu4t7LXygonuHmf5lB+Su+JZw9PS06ahRI/3KBXC/RDpFXJQ03pOV/jY
jQVGG93/All990EgMasBoeioLS6LRjY+3L+MSX4fSSzj89FF4Zx1h8oL+8aYFpmw
CXpyHCSfeY29/agm7vFxWR84xerICH3ISR8Agmq8z1J7U6WrRSChcLS0cxEwy2od
sttnBKBYpTJD3WyPwlW0S3nnbZ9PzqLGHsHPTv6wLnfLVD48VEgqzq3IEaGfC0Rx
QBlCYC5w4ejyoZcLfambMdn02HmBZOpjx34hZk003MIHwIwyZbjyIVdXM95f61fk
Yue5BQD87OkzpCShKY3Kl0Kjj95ZxBEh+AeaX7zYEng84pV8oNNU/pTwlZvaeMFg
xJeHL83kPxxe3K0Ni5PCVgxEauNOvj3IziMQbZEMPagS2rlPOLuKorUuIFex53EZ
BoHrtgQ9pHTad1vnepXlHRF/JMNaHMRjxh1dKx3HYUUKrQiujoO6dsmmlcRUiSla
qbvSsjbiZzHnFFfOAqJrK8syOk6aUIuXXXDOmv04xSb1YM3cbaaYz0Q2aS1kR2N4
F3ix8Ye1ZyAydyN8P+RubVL6j+rp2WzNwHqStex4k2lh6WCAAqZV9jrhfLBwDkXI
OqbrX2MWxgkaQoNCVSyKTCVsuknod0GNN1xKCfXGHT/aUtIvT5foBF0DPEqO0o40
QvisbSdLfqHaLkhKLKuOkdtPqlv7n6ZXPZAK4YjVRn/Zfcp6V8gB09vOuUN5YFSi
UuN/96HijhykDj9A7+i8PyY5o3WvlF7BDlChgMm9kxoxPTBY/e2IuBd9fdTpHza9
bZLf3qodM0VNmDBMEwcVbbT+psmt103Yef0ZL2lKoydBE+6/kO7FFnQe5HZazZdl
FxrCLTJ9CeTcnaEuUf5scIWzKiRY+ZTrwpPDsSBe1Ejc6yeGOTxcYLuHu3CKwoiI
MQqdhbSRqUAEWYVLg27cWG6EmbMTVdtMZYamATiuoAfxxuHheysuWXSrRZLhF6CL
VC4h6dYGnXuPuL6YF4/Dlow0MFpCrdqfh7xXqGgHD6K0JvnhppFfvt3Qw4OepXaz
pBmPur60XJ4hEzjuSjGKaW+8rSBfk3ZozoZrmXm+4RWvryRoYGZl/FYkg4Hf+Pnp
brbVSujN/LBJn78oLPHsbdhBgPIJL3anbOeRB8AOcAi5ZIMVTCldPhASzoAH0GMb
vyHPAYx3gzLAhJArqsvemZtlP0wpB2I1jfv93Jcka18N+b6Tr/hXWB5MZRdN8muu
QkucJeH41xWQWQvTMalDVqAc+Q5XyeiX86+3NI15q+ea99/dGqI2R6nJmCrhS4av
pvGy0SP9S9jsXKzMrQOsW/ZL97IwkngZXP8CYaddyPX+4zx1LEAaVoxPnb5DtxPh
2PAfopInlTjubBZ+IrZ5tedma0bAlVGAB2T85/vxGJ1vCcM+fmyk8Kw7TzPQOIvh
Ixad1ewWvEK7EFNtOE2SAr5UADGO5fipK7ttNcoLc8XxwAGawTwO1glQP/+hiUYg
KBJPs5EgtsZA+Nve2tcswLK2XrxOJH38sOGR6PaBm/gErOxB6pp/ML0ZMUFZAqqQ
jZ67tBxtKJwdwNKq/pZhAt1kPEGV3W3yBfqyxzv0X12/KXmbRdgJOWiNfiwMKO/S
yGmwFkXq0/rALU/Ws753cHMauyCdvgFY3PE8odhoEP8JtsdGS/PeBe039DWBgn7e
nYzlHRq5ozdrQPom4PFGSU4Mx1epcY9l2/XJ8FgMWgstc4DHI0vUl2gYaLYTjjKb
vOkq5+dgftsQ/8EShQpBgdsa2KHszVfRXHFvHtP4WvxVDbku5xfV4/yRaoHn8RSh
CrfcO3H8RfMNKyhHymg6cnoHDS1gJY5qMFahLZuSkKgp3ECh4L8ulRmZwlld4Gk7
gL5iizOO8tca1GSsSEh1EmlWs+Xe4ASNxNdWy1QQxIItv5XOE2aZGiijkO0yOhKN
zZFZ5g1rQ6KPkBEN7zmErA5nF1VUflot7nMfQPbACSlJ24aFJACsJBFUBh7fzOTt
LJN+8WAU14d9GLWGfJL4jLobZ6lZ7eBIi4SZK3GhrWDWHA362GlhWAxEZgouvmv7
M17BLjw7vnzi6iFe6OdE0C/YA2c7L4H7DFmGIPh+0zca5YenFg+0CnnH1xDu9D8v
rm9PIqF+h1JKCwqn3/MWEyu+XiHXzqXYQl2dVGpsFH38PcR8H3OUl30psTk9zIdE
lBZVZlcsAt9RfHTEthSTFbPCiYNwiqjw51FI+CBZao+f7/NaklYmxeCo3tEKjhIB
LkrDp5NmETJOk4yuLT6yrkQUrsP4lcDSEOgrotr2tSWjUjcTCYREZRwTNH1TwgTY
8xvNEflbCfuFxCuurO1X1P7lNp2fKrAHor3+afHrky98FvLjhAxDULtnVc/dG52k
MJJe5907+lTlU4IbgDbfDGIXSdoZzk4dtqCT5+jFOiqP483UgykYJL9im4zYRbTG
cDu+FOqgkWOAIGZnQY8YpgO3m2bqQIPN9Ohy06rJpn2Pt7wYN1FQthAXt8H0bruJ
cVyuphvAUQ1eJeBlm0P/1RcJJnHGAFgp50r1DR2xLoMa+pSg3tXY9mSOBsGCQn09
6vWYX+dXPKEU2oujCTunnHEWtI3eNAfMtKtN4oWmBj8XGshTnPI6PxeAAiKeZHBR
PmwxPnV7j0QvDKgw4P+92e1y63za2/gH96unk/2oplETbD84uZa2IucghC+ER8a+
JpfT4tgJRPZelkCkMVuLPKpEaJAwNRJhfrCBKMoFC3iimo6d5Re/wHn9b3rkS7ke
BC1mzB82H4gzAm9dT7qYgVilW60Xl3rjxcf2UBFpiIDljAuqar151MruGMagZn+c
qZGhu4fXPDodSmFpMgOZpsjlnH7q33HUXwAB6TD7cJxPGSxYFeYbSv/n6jzghWxC
3gwojPavaIFj4lg2AgBxAhfTjGJ4cK9OqYfYHa59F4Jsa4rY7YwYa48dAg9x3cKo
DIT/1Sopvz41hRSr7rv0vvEv5G7cGzp3SLcRvkFBaHnDdKjJHPqgYlv61w7oj/6Z
jm/F32jjBYF9T3HJQur5lKcdntpKuLICNQW1DaqmTxXx9lEMDPgJlS26yWaMqipr
zyafrbtZWIyZ+eAOwSwPP0A0sPC2vSkTWG36o0CAIYdRSSIOYgCun03Cbvcd+PQh
gk8lsOd2hSSASa9VnNj0LWYots/I/Zlsg1gookFjx1nLx1cQVWGF/dZJU0HkRCpM
dwS9VjNVknQRol2QE1juCxTsrs5YT9Gx8vCtGYBczeX+XZbSpAjjzgvBvJwXiZVA
7MHxaoF6Qs59ZB9caWzl/dFq4J6SssULKZ2EfjM2taZ3Ms0mrfjYm0Fgf/Z6YsXB
EXfoYQs/SooxViTgCIG2iUoAH6P1BMDSYwszLh5oWbZBdEVWHwC0a+2RA1ToKUYV
Zlns0WyVi94ZKQpXwlltr+pSt6m/FZ3G+8EH9jyzU4zWnv+kB/yxUVd19KPddtVA
SFb0RAcqW9gsrhgB7+DLNs5vsaUtV9yDlarsKGsRd64/vc3zU7lSDb78qYK0dyqv
1hqqti9I4aIs8rtyUwh/LkVGJ9hA8JEGHFuSZh0l0b2IO+ZNnXOVnDXf+Ir8cxz5
zJ+lmgxb3Q0WwKMgzWhZoijV6kc3QjjPAy4na09W/nXw1Z7YFUrwgHn2V9hj9Zc2
R5kZIPwE9Abryl/r7pb1KZfmmWOAQJyR2WxzsJPpxbXoLYn83ix4FQSXVcoZnhG7
NVIb73VOOcFmtpE274DE7ywYNt/cYt411pBYpgrBn3aYu8VXf/XVVawpOMANdKiy
0KQXfW9o4+8XMX8MW3LF6IQRYQPEkEo+vzo/jUEvF3wnEqLSpY+ANLkO7PvL86Au
uLz971eclt9ltuCiQIunnT5Eqd61pCZQm2lCQPz/E9MuRd6pGr28dzdwtH0nvvXF
CxIQx82tSpdekmeBsgngM0rBcSKh9zEP4pO6995hJs9NELDU9M2HxCkyx7x90Y/L
HDM49FI9AYj7jDYOnPErnxOO47uaAwrEyYNr4z2gl1Oq8E33Vk7Bl3M2qHeK5nAv
+kVRGR0C6Q2cBV1SV4a+Y4t1lZd52HBQvBNUBctNgt4KRzSJAYjCLt5RVz6g+yqj
8+QhQtS4gzhScG2RnM7+LoVFe6P4eLngSAamVqJgFvB61F8VpfTmypSYRJe63Gg1
3rRd+/+lgnWzQEVp7sCPxG8y2ZYFOdHg0DMKmO4OLEGMZxqojdGT5leMzLztRuiE
xK9l2O9VQAgGCohlH78f43KhS9dsqD0nfjmBmlEQ1mlMll46hZb51ghXnPY+UI45
Bfl/BCRVo/vDwWMGIn4F3qOhwncc99Bg8C5YlB+tnJ4olGhmhCutRmXQtGdvI+GI
9vgK+Ds09NhcCKt41ns+XHGEHitGzshYgFLkQhJ5KnZMEcXOQfvrncHY0o3aButG
Bxkl7xtQj0FVK4OKh0YUVQi2ZRfDYaFxypOGCCWwN+tFDloLzieLcSVC3Rxb2IP9
vJ6IWHoRksSmE9dzvq2qd2ZANZCzRlZrjO1aKDmu3Lm1PyhYmxXaXqJaNVg4ySc1
xeXj0VG0z4VnvpLxHUYNVfmeEDuXH8Xm4F2Nneu2NUv3mf7JK0JHa7qavvYX/fdp
y44f2VpSz21Z9zHy3TgZdAdlUzFHRD1hXWroM9Oq3lDoAcJFysq1xr7WniX8P5K9
hBl/FIxNWMlZ0ki9GBDIv49gZn7txyGXNmgZW1CZocs82WxCSzNvutOxf5UmP3N9
148rTrdBvKhzuDZgA3zvuNOhrBq0qJUbBtDO0l3sFa5qXsfP1AFUWY8d3h8TuU+q
D6uZBXbMyu9Fpf4aS9F5W8fvT1ycpBVMj8xbQCTjv9yFCVb/ExnbKS00t12Ex31l
UDg1gejFJvgeGktinQ/pjnhA6J19lmhITAR7Fw0Vwv+XSAXoUoBTYFGyparVYgHL
AkM+NeZsxbiCkvu0D0kyx8xvnTTYCB6GL6cu7/VgDrEYJpuozOz9PMmpfdtxrTsM
Dl4femeqZhmBNSMqe+9NzkPA5I565x+AzFU53D6TqUlKHgO6csKEYjZsKh+3XQg5
QYL3zgzBqWxn1LyFWFeHqFk4VpCEsAOI68VEH2HopLZInYNlR5ccG/o115144+oQ
grShWEc9udW5rkzPwGDoua+sBLzJFsrV4+qYDGL43C/RcpCmYWN51VHOSpgAIBdX
XMP0fPjti17LnFAcMpx/8YAAHRAOo5KFtGFzN8jtyzYcg/pg4yfXRkJhNQAYLJB+
Oag8ShQf2eQtgETR+LHbl6ybaonFZIbyAbFRXjdCw+iaS9sZ9Gh0MWDlbGLFP4WR
Sw60H3tDWeOexgm6sax2WY35x8XTQF7TUYZTvJJNpiBDAqvCxYUzmphbnIRr3Nzr
gtiC9zTn78YmwLUTKCy2ZnVwdigiW/d9qfVpd9sGhrD6LMaz6+fF2IlVOYh5/FMm
pxlwXtpcJIkZl2LjBLgqNre00ZSCzi8Z8UQFx6zaDM3V38a2aDwqLEU2Q7qKnS2n
f9BZN6zhWpGDUPbhkWNxjgEpjyqGsP9oC7D2vtiqA7oeLd6oiijZCnAefym32QhH
OzeXJfuoE64gz8s/c1X78KaGvCJACKBTN4U4bc93+dtIdYnsNAm6XR9FAjU35HLI
uCWIgVp+jfhzX9n99O+dpgsCPpBPxDQqhAv5JQrNc4uDvVa59vWG0VQ1uf9mhDon
IfNGZGg9RnRBxiiGerKiaSt0QcC4SHp788R2kK/tyrutLwbL0Wc80tXixiwspVyA
jz8jvvrGa09JQXU28xvyikOE0cQ6K8iR4x3ULApZ1hwskX2s4Mx6ckjmjPRlSTVl
t1nSXWkCaL640NwXOhHcU5974EQawVZzBCc+yywjAE4L52voPAI3XMGawsJWe0XT
h8cIQqJaYDpv8krwmOHErueqh96eE+Wcn/kOaorWCHxKvmzyan0bwRrcNbJIUInF
6HAYxNm+AV+X76gkSHRVbwEsLKTD+B1taSznWilRfSaHpIM3+Thcm8+Kg0vFxyLz
z76Rm0emtfdWhPcfMWIZEI8HzBDtKdQTg71sgGV3Vu5jnlE/1O0QWMyvCCkVwXlT
VFzbhufi0aE2w7R0ZI5eGkUDtExHcjXjX/z0gPIYT+uK8dHs0bCUpSP7lTM++0BF
O1WbL5X0UVXNDe0eGGYfsy5DwuWgM0qkuOd8XBz6Q8wT1r5kjMm6aK+NZW5og7xD
I9jvh0lDel6bAqdhAzsVtiht6pOMZ1EKXM9hIZj5O6UprvBOhDiocWJ9hEUfHnDN
QwUHgrv3OPeTOPUGwBR6tJtUUeZ0HWxX2SgoRantwWt3lcPw2QRG29ktCCoCQ7lB
Dvi4FNUfeTX1velr+Yr0lgma4GT4gVrMp6wwAfFp0Mid8AIQP8ZTi60m3HE2v/MW
J+5Oj25lVL16se24ObhyGAY2/FshxGrcFVYFjMWeu5PXfQpuKLrXn3WqtVVvA/KY
ZAVYAetVuzuXYqNKRSmWU5JDls8VX0fGrQtvI3Y/tz0WE9Nl4Eh9zxetT+eKlRy5
c6iYIFuXoUuoueGwqbZWErXSgEJAQwFvr9yrtli2nyrySqwuzVrrXEdOs9aEWu+w
+V4aJjxt0pMN9DYa8tths99JuhW1yMegw3C+2f7IlgwsWQgx8fbH5ualmFtBNxZ5
B/xE5QGZr7plGCYQiqkuBaDE9zzsCLYyFilnUO8+9IanIpRhhW4cVQun8OzZOpyA
C5z7H4jukESbNmpzoWY9/+Ai3iCUL4krsUh6glyyB1bkYhQFvggkq4xmz6cmEZVG
vsezEeF/eauqWVZ4GzurZ2i84twiDLJerveMp/gd2wHCp8kOI1AwhQPkIf7fKZsL
VReiKG0GGV5JwNqWpYcChExMWQFxpHKtmJ+ABtgAKVMKSl/F1eMNTOuxh35RdbGn
5oIOpNfdSq4tnJeI8szlgi/WN/baSJL1gaW6PT7FTlZuja9KRD+qMZFMDIdl0A4d
nJxQvoo8oJVWSM4fdiJz9guqpz7/hjsscLQLdcf4xW1skwH6nIUlzUjytlwV1hQW
s0T4Zr3VITUN21eQkdXibtOYqx/c5/yy9/v4d5C3OggOm3SBIuUgL4+wyVVu9iml
8BNE8+M/EyEmUZZeLoi4wcvMlm6MgrM+RBmVynsosa63SKUNOGd59ckPl1iOQ3PC
j/nuaCdVF5DW5vjCvdW9UOBthYIkL4TR4YLLFLDl6v3SKaVf16Tu+isOhURaI1iW
ouWVZ9RkUxP6EGamypT4Uxx/sg4XPz+lRzchYzTHHBGRdi2BewmFsbpDJUseLzED
+rLniZ70ock6yIwl+NUGz3Be7DIcSr1hRxFnQZTChIwDt93sKr9tj9xl7ajnrYJs
uZuOIuEddpY5mh4NwFUzr19p3jzr1EQV4H00SfOq6JbuqJfpDn2jDAtNqqYxAQcc
Fset4ORfzyG4YmxcZUeWQad8psZ1z9G9fqCHBbbsQI5Q+WnolcxMJqa3GBI7SVX2
mBbqsqksXbVegThe9PxXDxkEx7eQXApP+RxKDmECHatjPe7ysZmYJjeZ5xKDOszc
14OxZBLltNNNSSs2XMWrrRB7r5I+cB5HMiq4tmh8fM3aM4hPzzfto+z9XLY2nl1N
XF5/Go9gYOF8GlQGrRXLDeKTzmul3JCEiDEEK9oNCONqOa4pAbqRK9b33cwrpDwr
0a5qiJ5K505CBzwpL2oR8n8Ha6Pw63T/kZo89WSaAkVcQ4hZgbEeW4ww+1RlT91C
l2Uth+75xx9yYntPB+8hTfNCVTn6bQ2jjDnpuvt2V+pvf7U77oLMn5WFsjxxKQtD
zCxPqk8NxJ77oedxug78g9/t9XQ82hBVtEInyl6oV5PFw3WaHcEoTB7Oy7Mkxd73
h4yt/+AS6wGbP+fQiScKGHkraAkMvlm+kyj23T/X+JB4jNHAysPUtjzk/Y89MgZd
L0TAB7PawAa+wEuYvivQ8w+UsegWKfZh3slX/5U/2XPdf8TL157ahtrym9p+4a8V
E1Sso0O2EBLGSN/hPhQ+oOMhOJKqOx9J/9L7qbI1NA/o+GyvCg0CnJupH5LAPBjN
2LA8rbREDdviIFQQ7PAKoELphOlMiCJLy3wVOGC6fAk87x8kydy8rYZ1x8/9l0I1
QkYG+gP8k1GBeT5CKF+WlOK1M8uGuUpiCnXl089/5Phy+DO5XTvrizZf9ufjURDL
McqhiWnC0lQIuW+gohJUVnKaRC0ZmteJPVpu6XfdLB28W3zVjjNn/zXq/pSKsbS/
I6JihhfGctV2MYqikh8ILGbL+0I7pjqEUsmJ7aM6v7odmrZ+J1FuozHdnEpiVdcD
WaLEfecvk0Y56bDHDlkMD+To2ec98Q8lEWfzzD/FdQV/HvkjISVQw7ijy+Myo20l
jeAgEX4A9LuXvSHJ6lRf2OJ0XoZhnCOZ5pxK2EPgX/5cPoLT4g+gL8ba9nHaVh+S
79Jhc+j/T5RCWVPfsLC2Wjnx0Ly5z190iFrEgZD+sIHVgwpEede/cT+DqQ/MZpDt
3zDMR5HnKYtr71ssDQYJiGYsAJe/1Z9c082CV60MxTf+6bUyi2uC+nOpmsObwfPF
UxhGfE2f9nm8PdPX4ohSuI8Q/66SliJvk3Q5r0QOJerA69ICsDdtisq4DRxHDifu
qHUE9d/0PeIRUoJx5EYzHLk3Psmoo1PuOz2cClL/GdlDZ5F6reTTrmPB4ju8Okzv
hWjOodiE2bCXBLMfnyfks4eYNMExz/5oxJ1nTtoELRlRjeVEdjEXfxOaaFaPPycj
BsCWfH+ap9oLKDM76Pp3XhRmeAQsicoG1TMc33OGKLhLixGyEhcJyknLVxc1716N
4Ze1YbHwXgrpCMfRIdAFkysuLSSXT7wo1pRtSbwXYulLJmHHXLn+TwRsorzhKM79
v4O8+LBz836itHFxvmr7I1QW2IShSJI+2yNlOLlmhp1tN6qwrMtCtXi3E1AyEJVi
w9VNcyXFFNNtQtISDV14//icYancaYOFK1IwQLmS4VQgfhRXh4WwHuON7NLxQ13q
kaG4c6ZM//mk8QbdB+dwQPwTlhbxZUZihfOIyWW8AYjFH4l/bKxTdbJZfGtMwxTt
rvTYam6Wg2H6QLiQbumAGju2oYmHGJ1uMGrP0McECIw21JTgluv1YSGnnqj3trgk
vlPD4U4SLLiN6c6ni67ATXrh399f73n+W/XM24be5qMHVbMOoiuuedTV0V+58puM
1f9aWzMu8NieMvNazAwlBhmpiY5u0qOhPMZJw/m4qMtv5p72bgZT2j6MNzWgUbnh
gijwt1e9bul7W/7+NR4BslO6gXJNcqcjB1L+A02ZWTmHAokh0DYkj/PKZFoB1KjR
f9Rm1ILmzEe7AsCppJ9Q3BvWJmCwdePOlSjvvv9p7L3gC4zGrz26bVGa5nTZv0Ik
gZsNCflw9vIYmHT/HiZeKeucAovgClYLoKU4nZZXNsdtq3++nglfwJoC7BH+M0xa
FjbgXjpcdk/1ekGg7AVQ8hk/rP3ZCIWn4GnPhbF/TFJB+bwN9+ce+rSd237v3gST
1db0XV2JPuQ4021/QIdczp+X80kvQkWjGtMxmUJkF/fITFqhL7BP8HyEtYUuM+KR
CFkxfknul5OEUFMImriF6OMAsqlqRRASyNkyiNgjY/3UPsrtJ0rynYSYwHSt1IOf
EqJq9lru3bmeMUDRPkPk0OKIcJyAX+LMWduUeNZXtmn/4XPhNLQVHdvyfEJij4zS
zh6cnkH0AqYRzJvul8/NXPza0PqFZlcUhqeX7XzlfQNMxsI+tzHgsGkFraUpqo+D
fZb+bdUkOCuqSjLU55nhb1Qmk+KGFI9O25rKmZLzDIvTcB1zNopDxQmZOC+fLmg/
ZOYjexq3VjT4Ha5UqJU6H2EzE656gWDyfGlKxEzzsrjbiLZOQTUuk9veip2sQd0y
4c5jhpgzoYI2S1ZRrrMigkOhUJu6penunvBa9XhgYlenVdKWZEY5dj/r45oXnC9w
5EpWcQCvmv64uNQDRsj+1v95kY1bYrxaHqpe1UACrk63SqQzcvkTpKZZvgzijBva
sdtgOl4h4ZVFxNhk2tH1Zla0e7MLrEJfq+0ei27CCdLipudojK77mdDhQ6bFh6Qq
fcjvNvs7XjerOxRYMm9d0nA8waKgciIRUVDqodKIfcdmnk8xUfyC2aa5DZrp/sSW
Yq7GPd7qtlR0000DyVvuPlK17MRhBw0MoeELtWLvDTJhWTthxBESILikM3Koc8ai
WDOhhQXf6mfyFWsnyJGE1np/CBNPzTmoksh0jHhDCa540BxZvRDpWZJAbhM8o/h6
7ytkPfGdkzTdClRS6J/wyoj52tGw86IlDZ329CLuf/FxL0rxVj0bUqxroIn/XaWs
EoqpOw6gIaKd73xJK/RH9ynAljU0fLZEEMEYcPjEizHZZTyEiqltL0heE1JsNL3f
2bwDk6sI391HbqCLONG2VsQcFHpk5wQ0143ojWnaBx9aKsTKjo7TdKqHn8GfzZau
4ya8BUTkV36N+fcMW8h6dU3eiEXGWrc1CC+rtRJN7QF6gweWLkYdNbqPaO3HHuSI
mKhbtoGZXzYYfuKOk65UIAi5bwDgJmRL9ElDkTugGrOXlLwfbyXPzDTHQXkinti8
WIbVTxhDWbMRmytXOFRVokIyG7nDr/Gbvdig9ryQtUutRnrMBMTIgWZdbvr0fXOw
+NZ4SFpcutzsZ20e8n6zaO9Jd1sNMc4udhPObjKIONL6Gx9+cmiD23GmR/7nyMVT
Wohn/MVJm5Wvq0+PuaF2I5PT1CY+xSa5DIFU0vjSEsKMGGxdUXea53jn31QES/D2
JctpjYMrTwC5nLQW0+Ho4N3dUMwA41TIXKXELOD0tXEQ2HjjZsxTR8+Qk6yV1/h8
Kpnisci4KmtnWOOmC5Ubr58SsBaqaUHbICbjsw0E7p1SaLbcd6Ja6pci9xzBr9eY
gXTbpznLazvQNi1sPozbUjny3iLWRo1nNaW7Sib4y61+O0yGDBjHGpGsS+2yiU1l
iMuo0pv4VFryWwcHKY66B9Q1I0RBsRwi8Bb3k97fJjDXj6PR7ye9aBwZXmNHg3fd
4/vqUnCbKB5GKglwSYqtopkqTr0Ijy2VLrbDPQef/GK+ezTW3Lwx60DIu5xHcgRw
UH41QxVsbSIeb4jAHiGcaIOXL5GWrZAEHbFMTpLPMRrByqLe/n94o/e87vW215On
Vpaff0glqLsNf9R6DKsAvyOmUTSRptivuryJXQw92QdSnDPSbAYxpDchydv6nFd/
47omjTH+fC8VPs/YaEGslVQdwNqIh2+CIV3qvT4nDypQw5fEKReAiI96FuZq1pew
flp5/QgZk3y3LsHTylaV4cQ7kJOwhD7f3JesSNQsKlblZm2qAafnwTIYChJcYhEm
d2dRuPN9Q8EH2oRxa8XG9Z579qwUJXmQnCB6qyB0ANTPXHV28WMssNM3nQa71CwD
XajUptLna+kSnMs7omMjzOZhNnV/nIbl68fqtoj0IAy52IauytNZcIH5Ph5U9kln
SkKhXHN0oBaiOKel0rUFslF4QWaA3ny1db0JjpNIHDAJTWqd2/O+cdUC8Ow3QTLx
8qFbtGEyEQpp4GS7bPeJpGjn8WWM7NdQqHFR9i/R4rLd8IlIR8y2Yt+zwZM0Md9A
ozmurUH5Ah7JE9tesDCsuAd3VW9UcRnaXEchzoFtcJmP7F5n5O69gZW3AeMi7ti4
Mb4CJ7QcBYYg7KBahO+3eoksY0Rvn89hBz95t8vq2DnUs/bp+8u3tFrSMlQ37m7J
Nf0O2iqTLbrX7mHY31yNUPqXfLyzY19QlVUJh/vr/ev0SD7cuTdrW86KV+XW/XPl
JKw8AG0FZz/LalBtfpxWRorTnbGVOCXUH/J8MaiOX5DQRtbCBJO/2goZGxanMzI1
8iXGrXbPRBLCOsMd84EmgL/7RGfVod/8GlG/KCGWPtLtZa7e0ymoScHoOQiOSxm3
dpukODDLCZBfxXcSdhl9yOHHyDYDcpmpIH7tClgJPHl5uXlPGXrgQ2OKMH/mraRp
HXJ7UCpVLP2/l0sQtkiARhQ+SY61Qtq6OSWWuC2kCAvH8zuj4UFqHcZgSyqVNWoj
ROmguE7AkOpHtQhDhawnAfy7cuLOWEN5FJJecYejztJ0fUtGGlY7FNXhIRlTJtPY
nAMFd3VcweuE//fd0HbCd/SHKYvVS4ocQ8Rwp0ZqnrxQY49m1wntJ+NoMh+lO4U0
8KxBr3k9mhVWZ192KtNnYGngDJDmkE4FK0lN3FZJV6HOhKEZVu5Tjsi0Jkj2EMQM
5L7P6krCWmnp8la9qqpDTQcwGDJqvkK+F9OJ/pSB4WEZJRBlfvnCaQRXlttxhqjS
aEgLeDahlZlKgf0kM+/HaqPgpuHePGV40fV7kdo3Ahnmv+JUsVBWOvDBKk+KdY/V
P9qlZ66whgGDDzcjcy7bSZTRb/6d3ATvbffE1i5Ywv8Tb34l3AZAOpYUPEvqk4Zl
9OfEIO/5/0yhfhZ+uFnH3vZC29lhCTTewvwODqLDIHNRJIsrDo60R44GbL6gJQBE
d7DS/a3BVL3BeXTF8PogPZFzVKnznhgP4aLfpO6EgkSMP8Q8U7X/21fxIyvO1Org
lH4Qkg3p/vDf7eJnXHyucQ6oAulO1BVL1sSgWNSKkuMV8sXnPSPT9VUcrKEUk1+B
cQJrxiXIaduRTh+lIBK3xslg2neiPJzGz1g6UsRCF93iTGwbR/irc+BZMsT1T1VP
X+fBhs/Gvb3iWcl7rDylxPa36wpImgX9N6mkd/d87eYawqdxl87pxv9OrqzoXg1q
eAW4xdzpHF74lp4OdhyvW4dWKNNHLlW8KFZY/tv88PrgsBxtCKbapyat2/QEyuRN
unfYGowCxbF5a5dR1VazruwkbuzhLAKUzBt5Z3UP+q1/dRIwBx+zjSHc9Z/hVJoH
EbWDboYh8u6njapVfqbcH36223CwjUrbsAHoV4FD6RDJJl0MKDNdheLycy2ox8xV
ncgWfByY0S7Sq/obbMaUvxUcUm54TEJRT7KcMJjoLRPurvgKXADPBbB/n8mEOBH8
pO8Jh1dN1FpFHrI6p8YVHUG7PeogWDjrKC3bQ96oAr//RMATGbIMvDIea0iGokxP
hlxsrLZ+0HajHP0JV8xtvyiIOF8nLq5pxSw6Dk5M+fZMgYmK5nY5f/p79Xpi3nex
lVy6CN70eiEbeVudNRuc+bN8zG6xznFtRKPXlnyP32jS+u4DELD69CAAn0DAOcAj
wha0IwBiStIMmzSa58bcq+LQtZL6TdMS9rEfX3h6zlywn4ff/zKrV07nHNZ0z0nJ
XdNijIFpoeRUr/8I3a4mjknvummWUgfHUSnubRo14GP6Y/4/fBDJblqC/oUkh2hf
nlydPOZUOI785rEpvkxmPKbxO3b4HjrRKpJ4zcQSIPr+2IWKHYRG9UepKkzfCijz
E4lo0jHRyz9A++GVjd1cf1VmbknJmeGgxhZs8FuRjoxg5mYg5wwbEQtYwAJtie9T
UyIpML285I6EV4+PoovG1Zzc7Z9W8iFmo6Edyt1NM4S7hd5ro0dpeL+v+SZtEEdx
x2Xd6xXumF2M9cl1w/SUMA7EfDXRu3qwIOJLwINx3OKlzZ/60n07H0rulb2o2IL+
UQpjKHhX7I7U94P+XSMQ4gXFR3nzxtDQfCtq0kJ89sxo9VVN/R3UW71e+Gnmo6n0
Zhhl1OlHNzLtEVEUi6p+3Q7ApPr423eOyHFUgX7l56tdWwiU3fRt4EOE/BPWQxl/
qtnl1KgFkro1bvkHqhplTf7PKkC9EK69UVsygrS37KyK7gxHVzjlfwf+XBqZnBpX
31pdtmMJfXek9N+QvncbEl8OT1eJmXPbsYy1FcfLJJLXIzl+katb5p0Vu7KjsxYi
kLgdX5sMW9rMSfPKKpF47t9dO9cntRRQXNCxUS94ZtCP8Nyjpi73hsYMQl2tf6bE
t8YwZxP98nfkGkkDit0ZwPnlPSODW7H1mSF9G6SHLsR6JElOXXlNUKec4Cn+1xjQ
RP03IcXM9URDa6ykzLatXVyghQVBX7tgXTlhXWojlypt9TGu7Bv/lbraLGzNXFoZ
h5+AgK7m5C1VPoAc9CAGN7+et/A+8urq6nyi8oqFgDT+hIColIvr0iRRvTFVxOV9
ozmtfkVkkPMBDylywiQCSAVfG6itF4j6OfU1NGHqHYDiIxXPBTR+VYutgw6rtyLe
z+XpnzvPOAz6GVMSI3GiGx8K0DInYE5ryXyjTFz6QvV0akK6wXcnvs/MDXqyg/fy
IpffUt5GucBafUdbWDelbq4amCvjk/9QeuMTLdpMyNK2khW9x8UqbPG6ColnzpS3
7qKt5LdYKer1XQsko0fwQ1rwcFbbyOMALaE6/dgq8kVl2WQxevy+rrCk/jzpMGkU
e2meGA7n5NA9/lUe1FJaMBRvkVQ/2j//AZ8ogSBqPKxpiPGBl/SSRy353tZEZqGx
rT8qup7GjscfYDQLNBB4Nr8lxoRd0T7cN5ZYBXGX7G7heZRsQgAyOZ/IzYHGbQmD
xn16FOOjs7NtfUQe5JSVcTfjTEfnJP10o6+EF983CmoPON3ylJVv2SuEC4yVdCKj
5uq/wP0tOa156GilkEisFmWLmBSbLW69ZqWcgSX/GPhda5E3b6PqhzQjNuJEr8uG
ircEBOr0c7W9fYoMaho2B46KQj9zLBXC+6850OMg/he05N4VjuYkoaBJ5H8Brsuc
rY3ngGpXsCLSbod88YcNskhukm0pJ7P9uGHVk2SQFotsFSaYu45DmSaXpSMUBBk0
p/PNed/7ge6/ZaTmOgvJVNAHWU2TxyBJoz0J4lU/DRp81SYP2pUWYc1hnvUroYPS
kqE/V3s7Zp8CHAd9ZUpXgpluXfXg2xO/EYeHfolRPU9zj+Z4zc6JPAh1ggt0gAgQ
GqYYfqr5Tkh+WYYywuo5cH5ezper8GnzkN9IUDHTH/ht+a72g3HLaz6rm9nk3PNH
zQWzsZEQkdt91aW/Tncqbv5t4WB/Xrg88Q1whVG6nu699seDhvzIG6yX9il90MPj
p5rRLD0gPb32PcPbmH3vancvvf/bHXNvifyQfDtZGebe0To1QnY5/0vwhiJ+vuHl
LWaNuHloi7XajZUAtWd30TheNdbG1LBr0rC2uc6s6jOaZSsx6nKH+Ptyza/1Sakt
NY4aYqjuB/qY+LfT82LvQnt5e2do/q9+vl0RZCQJfKfHF6mKHsN9h5FHQi9TyF3C
FKN51HzMEUCe5jo9lrW2kwDzKOn5ObxZI3AmwwVmp0FfbyTzLdB4Pfk6aUyULZ6x
Ccj4yfXYLVpWqWtCo2x4F9cOuf4nSBp/PDGIIfSPsHR4uhCCY3sfGdnzd6Zu4YIK
z5Eazoii5kGwIcUiJ3aej85iGEndZrfjSBLJZ8NHLY1JwikM1g3FM8v5irxOI+Qc
muMUzjcSICwNwBo5/lbtl3Ewt6YWNTILUX4PMySAWMc8G/jBeLWb38rxbNYTWP6K
PPTBJCkCQjptZHHvWUyTlS+KSCH6uSaglH8fODbZXdz/QsqsrP32FO6C9JsqeFvD
DPUZOmuxL2vx1k34cGcRLMLSGOYhWjTCw8bv2puxQOwu//y60ElAd0L2owVwJE90
/kCNXj95WGMiRHNHClKobSdnJB50H0YLWhTRYHh884hcFMAz3nLf/p+8DFBSGjtR
w+2YPDy9Y8vBRyqHLo0EhtzgJGMY8t/ZHIwqKRvlvd15MDE2jIghC+QI9ilxk02p
t5QGcClAWC8Bd4Xruw9cdxCqQ9eXFKUV7MdCY9N1SuYhw210KUPu7jtjtQyIP4Y6
kv1imT8lMEy5GADWn6o1cvN+IBRl349DbugRZZeYYDInS3Z0LmZam5mO0L5zp9Xe
llbu1e+rAY90bjlnoLaACg9+guPC6zWzY+DtzqY6ZkwEPAx1RV0noTXDMfoazsoF
Udiqbg6iVpLmMO1wNdC8YV4DlPFJNb4aRSp64lxF6ao3obdHdoVHFvyGkQMG44t6
U9FJV7YgjNBc/o7FVG95jGivNZjIn4NWxIWIwYgKkE9SigBvWptGnoXQHFtBBfFY
kDaoJmH8X6PQosvBSqahXNhxMRFhFXTVZsIfulNicPlmFUWu367ikG32UwYrFbuL
OiDS0Fgfa48MC4vsfLQwOJT6PHa9v7HNQEJFg3AzBLg7UUNuUtpVlY1OXb70ji++
VOTxoFIu8bh+WyHgxPe1lxYQRlplqGKdmHeEgaOl5e8C+E5rGirpq2EGR255jf87
1ydCADPjUlAk7h47PWyfC3NpXkt+ScWFTPay22ObNwNrHqYttHArokZ3BtLnOaMu
2/IxZrkNc/p/TTRoRR7Lln3ARV5htbZGm2rsCHQNet9YAJiqb2mgNSlSBXLeOmT3
6sdzHEnnrapAAKTU9jVHSDxhULTvJ3ZIMudzdqV90VtbDGjnj5k893kpvMHW/O8U
xetBIbbruCfB4O7A/NwkkkfYmvSj0aENEhNmCg0eybycjnA+uBd6SgK5NtLnf1HZ
sxiHGHpQDUjChn3iFrKQRM8EJexfq/9CQRGcXN9y5j8TetfncqQAQtWkcOwCMz6C
GumCZNgb+c3mfARMydervUAXhOR96jPlspw/ATufByW3DZ+RYWo0uE6t0ZhUTL+M
Nv1j9o6dJoJdqOe7oMU29JARJPv7t1rdnIXChqmZKZVM8IWJ39b3Lj3/cXtlAqJN
ZH1I+Ens0CCzFGYxWZExW94EAIUPCOcKwfBWvOf+M0ZDCxlXI7bVW7/nLsuCcQs1
MD7m7Afjt8L+SEyY8kZ4Z7x0m4Ajq9XIVnNs+8JOEuSioh4wJNol/Tze1ckru+4t
OjoOK8ramb6cEf/98uGO/zd21mstyNMTvqvWr1B6mXzXXsiNA9jPEg2ksHS5r6Dg
w4KCLCHUNElCUHTUenREabfWXrda53IaTIlhXEailYlhbDPfqLMzMPwHmT7YJnye
gseDGaYK0xYzpFuesX3I2Sq/D8l7unIyUdZ3jFQ7F3SiQNIki9UOqsLpHlM2xfae
5WT3ArRaZ+GwEOK5blsa/cUDkACT7c4BCwQXPBNTMqdA2yeBnfDsXTn8e6zO+gEf
RyD94Hep/kgcUnnTRa+syHaHCigEvIcFhS5Baxel3rcdSJcGo49q6aXLKDZVlZQr
nwIeyjNYt5uFZkm6ty5qyvKY445VkMH3jbAnkGhMP5ooT2S6RSnJPdABOVXJ+j3a
4T9yzL/83Ysz+8tGnslR9mgVsOV5yCajfUvnS99rsHpc/k7ytYYBqnkq0DVy+pQF
Yvr3UdGA18iobyqG3bgaZgRKJ2XYgGkAuc3lbf+703+vxIhtZrYRHr/t7iYdRjNy
0NeZNs+0OumqQ8stFXGtja86HYvi/kibSzjTnVLJyH/X8DJcg8x1XNU3n03AtvVh
3b8Yy/3TUXLjyW/NxQUq0oe+WTMbLq/UFPZeYIHc/ImjsrNyKeFQl28Anj5xlwKf
nVLr0jSy2rlf5YtmtM2MW02n8+9wV6HAWcuAzJTsIkyVoKZs/FRUbN+k6rZqFYeT
DW2oIZxz0t4S9OJ1NieoRp8b7kQEcXs3J8juFEj9sSOhULTLWAqdkzi5VScrv6am
OIo91R7R2zR0yxD/62KUSE2wQf6HlQIWhyWwrWtvhNedBu1nfjOHGYp32wTaIKq/
TxEssJLsqiPcJTyw6xQnN1TOWoCz5dzTxUTx2vDsxQUotUnHcjggmAPnt4W4q2x7
0564sj7RkAekIAiD+8UeiacigsEFapJzeDcL9gBJNdZg4qdJg2Pe0bdsOjPOX9s5
fcIw9uvzoZCBjxM56xaVAif83j/M9QFOTqv8AFBw7nUR7frVfdgNPF6+OkRFxG/z
eyofzoh4aPbTY/sUpeK+PZzOSI06AQdRrF2b/k6QV4S7JyxP1ZmUBTlpIBdk3mTQ
2/jgMjWc2z+NME/fa3JnPH6Z9ercCqe3y66NSlWBfGkQwcULAXyAcXLQPzjKnKcl
bRReR+ruCkTnc6pYKqATiOgmQaIJ1lhd7yPS7YriLJKBVa7BCSmoMFZpFdtk+ZFs
FxD4SbF51D7pK61vIDr8KJth9nGedxGhdVjpWG8POMtPMSBwuQm7P0F1bIZHJjBo
FJm2cEMzzWhZ4eB1TXIRAXHgbL4sZ0+qGJX2ML9MMbAc+qYp4Bf1KaQxM7DC2U7k
Sa7e81pyILleqtgdBwCTvu0KFtj/qDB3suB3OCb+fKR15oi9SucSBiMsymkDMjz9
YDY7Cge8UN7ViFPeThS/3bjwbPrRNRRD+YxQTPDZHfSBKpQ80NzEHgZG/OhTmLU8
RU4sWtYFn4qIpG4exxuCqRRJ+EYhQWCOsbOPWJ9iMrs69rA+DCyjRjlumafFKG1j
x9xXBBlNh9y0SFGqwBjYUgNmrg+yoEDpArFDA76xPIqQADHKmU9aXyfc7tRdXMLC
4fdSLBCmBBbUfSqQ1CGJFjgDCJQq5zXDZaBjkuITO2eK7tD0A1D1S+wv/yxArZ7A
fo081jaBu3lyVZoz3pGSUAGORzoZ1BPRoVfltm/RUOlel8Zl/6QfgtwABamuxlIX
YusIBu9a1qqzzbVgImUFKuuWoFvqBoQ7GAU/snyamduVUqQxV0jaw7Z2bCcnPoD6
fT1E56cA/Bj6DFzy/jY+ywmgFlZhuhPS6xKhY/UpTSB4OpPV04J16gYnnEQbIFg/
I1UZRhRj1MeP33dZ7VcRbLhDt5jMjUdnJbgJ9zo/cf0k0cFjM9U1v65h5D9bwPuy
2aLprRDSVHtpvEyyMUQQhjdpPOap0bDzU2f7hPl5yVX2QsOwYV+SNBU3Mez6SO6S
WI5oUhzxIkhmLh985hAkQr+XipWM/Gtd6cQjhAXBpZ7KHAqypVR3cS9pDXjgBV9w
TQSF+gZXS+MxVpZVZlOK2XLN6W2l9yfkKIgLVjEqVCL9xrXDBzQSrXSeyxu9/Bfs
SOitb8E5HV2pcFpMXRqDW04GG5sp+VBxvmMDecNf+SOgfeweN52/zof/EI4sqeim
qdtVRhGnG3jIRuMea4ozWmSn8rxfxHY+pOmO/6ZMmMAX+p3c41Pdxql+cTcx0IdH
mjW6xglllBu2kyQ8fKe9da+3Yw6tmi2qHjY2Cus7OaPsco9DrGkjA87BAMWKHHj7
Xjx0dVBjGNWv00j93mcn3cQ+n3vquycruLl0tqkIyy0Dkp3ey2CdMkVDHZP9D915
/rUUNdWXNH6MAUJdhF3WvmT+LTzDlKkhjjQdTnfbfogPaKbCuSXRTb8nwCVjOvLq
0hJoZXHBSIj+3kF3nyL/vdKORb2Vqg0gisZ92Am4wUt/U8xGgXqbHOtQgkID03W0
UPXI7zFGFXJz5VrA9VtWERRYjwQerwp7p3yuh9hTG/NHVolt0k/wmXFIGmawfJaN
1lgoGOYlUGItqIqWkrK2vjKNLbpkI4gMSzK4SQZwq47CCpA3Axr/0c5KnXCAdrtr
yG7MdIJzJSRDA6BwlDuhKBh0Tsf7U3i01P5I3Tkt50K681rBcxAQiuCOgPyk6Vx5
H9Xl6Zq9YO+SPmz0ixZnvbUwWA23pyG4wHlWr7VJxBy/s+QnHR+xt0R5PVbqB4aE
Fw9fTwMTlgZr9XqUBxRgeBg2jGjkUYhk86WQZlStWNFrkIGKkFOm98AGXFM4R7Xg
ZaK1X09X3Rgbp8EaLCWUHDse04bc/SvNU5WyM4CbBoqZ3I60XKUJTb/kYh43xn2n
+xnIMy/Sp5GKb3RVhi50BCgGxIze5xIUXsaKU3O97d+btAgYEIJp1LQ+xvakGNwV
ArUlffhC/ZMlIp3gqplkQSc+hWEaGMMB2wWIyb3uFR++XHuH1chG4G1jzDxPq7SK
B+7oEHzHg9TOGXpnnUCjvDRyT7OgSiEHkxivbP7bz6uKvJmA9VfmlUiJB6cb0QG7
0lFUPfOR+FUObntnRw5UKNWCV5zmzqlSnR+CHfXAoAMdHrPKtxD9JGWXlU3YZvVF
BYwALTKekc9UUsw3q1dstf/uz550hsBmAQttr9/NtrlB/078SRgvI2jd7INhZQrO
qSA8rZ05GHYkKjcfSIc1gcsxCOMzZv0NqogmJ1zwexRDCHg9y2L+EISaM8MOY9xl
28ljjcfoBmF4Mz5j5I6e8fQoIkLnAMc+uUXWCJYtRVjjaTqTClmqrTtjRNvnvvSo
vqJgEgSeahX3gu/i/8QBlLq0n2Bg6cb3XsNJn0l9acQidgbbPwBOHJaVmuQ0Cujn
RiG7+Vij/BCewAZZK1X9ys10IzaTHBLIUTekkvvpDYSlDcLW6E0gzacX8nGeud0Y
oRCZ6nA2/snaBsZ6JtuKREVMlofcjmiiWhZdbFJ6DI1MKI6XfNKXBvEBxrb+2pfe
pwS4q0wPligENA4i+kbcaFezx+ZcmM9WhWlNHHlQjQD8KWT8o+exTpQeQEh9PdXR
IKOu5/tFzRr/cdjxdSzwMNCipCwRUkrC2I6WnaEz4WYpzgYARwEwmA+07x2Pdqq8
Tsh+oF71JPbqU066NjKteTT+vJ2Q0mdICXY3NDeq3tg1ErZt8xvSRDCYIiGKGEqv
kb+2mOn6lXu1nAKFTspzgaah56RuR+uPIgmE6pouVKylOF63UgXKPZPCfSCD0Lm8
oASyvJOXoIxdLf61gXTFjqWUGer171O7z2Cs77sgTrKu5VLn3Iu3h6wjDp1dZGtu
4dELeKcOSWtLn68gGEZgqw/EugjyR4X2A08ByZLUJxak24Z6MWlSZiviq1cKhRlb
q9FqJeeqPZhVISW9y0rGI3CDFWd3wy0IirjvZGtv5J+Z48IPr6f4qvNRx/OuNtXA
IqP8M1fFoiYzTLIR63bVYnSe6GD1VG3i5RBW8Nyst0Ueu2oYnG9AoDvAnjR/tZyG
pqoUrcSnaGQ6ssFs6P7GN+rp9XZWuahPcj2Qn4JtXaIh0e2N1Fl8AYNjd4tMi+EE
wFMEygEdpsBAc0JFEF9hdoETumilnXqj9elQv353PuY+yjVR03UJLOJybLsx8FWM
PRZelRQUt0PZqal/zU46rkMxlwNZJLB1VTsafNvBPQvSkrtvbNsgAUPGQPjagaLF
eEF0ODoQjRxuRBLqYL5hrgJ9G3f5H5NWVCVV2CPLaLyIIrxHb20dm2t0/HC698xL
xYwaFIhrhZlSQerdzsaUaxA/s6JHS45IbVp6ZEijI+o9wlUCFddtMwmp5lkRdieg
+AhxngNxtPT95dWbXCRsRRPeAe+qGWda0v0rVJp7XyMUhSNaAvvAYR+7kgVOwT1A
QJaVp1gzFBehfFDIG3HfwepH/l4XKNdmJ5NhMj7oLPrNfGDriIoMzG2ZJeJ68c8L
sZF10JYwYJfWmY/lVuw8fIzXmLKxxzeih7Upscza7cHRc8n9ZVvshhZRQ9i4IWzZ
FuJhwlkAKvpxGI1sn0Lj95w8FTJmeNOCw1py9WE0RFQ7Tbpavpr8JmYTttX9KlyM
ah7J2RXp8ikjyRNnUfm6T533EReLaGihGAje4bUavyjWuPg1OYHBpUqdTgMWfZoc
W5cSc71pOJSqjO2WrifjwihSSBNfZNHCV4EQgd61zhJaIHsAITohYzjcx/IBDm3f
/OZGa3ZmWVogjO90+LxUS7dtA5Zh8v+LKUGU44qj/pWxUb0JEPTvEIhHWGxzC0EH
gXUz5IqA8yZvkMhRM1qUJh+0MvNwq72j5vxNcWDATbI/Fk4ycDqZzw/eTlI+tuMo
GXmVyif9oQQL+8uYlYZ2RRLcxo1tLMgSeLE/UIaMT0f1BD3h5sbrZgKF/OKTkoUF
myA365G6ApxjGkw4O02GW/qFG31dNW+Ph8W6sB6Q6sDSfLaIPsmEBkxTeA5oPvZ5
wb3PNe97TP6VhpGxArwxCPNkZR7Lye0EOzT3IcZe9veo/OEMPCAYvAPvKYCVx7Cf
4YERRhH3jNCsO3/ah7Sx/rvnrjuV+WmksNdACrPNkRfOPwJP/3/8GtpiejQ9zLjD
J9ytUJ+BN3X0MI46K5MZVOL1LS/w0GfyE2aDxF3WfeW1/d3gRptXghCv50NhkyEu
A2wJ1489qWe5+nxrGHzQhysfTLkrgEAymV0G3w/6+QcK+CPf+PnAey8YfdfyL8EI
vk8KRqgYNXxuXF99ky4crpf7gZPlG9F8/hi7O2PsU7+FO+nMQ8M+dPMgsHEtRXRt
u49+7OAH14jA2zdKLIYS00xrBqsStFjRzcXrMlZruKMZVi9lLaioGQZ7hdHBDSEe
DBOWiZofOz9wWnLvGPSFj01Jy8sjaTL58ku2RkliOJRVhFE2QiCq4Uan/kdT5lCr
wZAO+8LaEmsvSe3IJnpnzV/9xhCAgRneEXeKGKC+5FMDA0UX/DvnlmsHfYDgZNbk
oFBFVys1wyodS0x2ZnjeQYNMZhhUsHvirbOre0vmqbGnLkrRMMdZniD01QYnDFRW
hUgw9FhLR1ZsvhwzNcHADZvDkNBaZkZ1EruVtRIDU/rWo6ZqFsx7qPGNTpiUkN1c
HPbwqwCkbOeKKOSV20CiZhc/J6FqYsI+YEFe2vxDpHfchZtwe7TdZVSLT/9exYVB
4zopjMaHRtktfulMXDIYF0eDZOfzjJiXFyXSi0Pz9Lhx7whPQcZN1awLDzpklLpt
0E65WY3cWwdzrEUpok8FQ3Fjb9zKeOo1FBB3mpYqHAD2sZgY6ZAs9XCZ4VHeu3h1
hH1sqbr7JzpyvAG4/RliVXIMH/eny90NJYFVVHH9CJrHM2dzsoZAHN4bOB9YOif9
kwfmLaq+9Pcx6giiPq9FivvQy3k/CxHg7Xrpgsll9Htd3M2prk4Oh1rKPVGlHiOV
fBwCCbt5UoAshp8QgZ4parZFbzBMzGjM8k+nffNCK/fZ3+566tHVMe4pkYVSwI7E
d1GS5YYAxnRsJXEP1RyrcaPTyYyBobIjAOMI0OBKcuSPwiXqZApejEyvdovXy2uJ
F9r2J013FG3GTZMBm6g2vaUZ6u/UEZaZcR8Mgb8pxrfzdGSE9hjq1ypaFjWnW5ZX
SDzfA7XJ6R0ijg4u+FnPWSYxLX3vwjM1IFhN1PsTMRDNrEvX7ufVicTbQQrYazwq
OoNgn8hRzpeFQJWbhHvywUEhSZFY1vUvenNHK6zWhMqWz/UrCE+Ra0ulkjNFw/hA
Kwb3CHD6Fb+SBVM6EM/j5qpgGay2xoF4euw2YvzZ8wPpG2+Z5UKu78ilB6e97zoA
y4ktCDnlonxLdYt9QhSXVRrNZXS0Cuhg69kwDANzyfhjkhiNXHNKTaw4ACLOmURD
/41kYPEcSwiPyGijC87qisBQm8hD+tJhswsdUefsK5yC1DrLKL3eDGX7zMkaQIh1
kBClwWmE1c/Fp8relwjlFXITodkpTI9opIXtSwR/p864QMhm2f7a50kjOXnRmFfQ
XQkY2M68CKn6hyjUhlpTa+w0Qaafeh/WwyKwvQVbJVQ0ca3DVkXgPl8KV4H3Xpo/
IqXl7X9GDj05u9xn6XLGPGonGNxXz8hEXNl9guHNoRAENDNUxI2sHhVB1mQVpPmq
XfZtN0xB5bXybVtq+7j0uagv981xuGpvgAT8q/f+diEOr9RmNRoSTKsUAN9HDciR
SGTY3a30UZtzRAmSRmuv+i/1wmWxKSLvcjOnj6zZxVgd3AuMlPaa0ImhS2TFz8x+
eks65CWEHi0QcOuwVx4xVl8eNhtuoXvqY32LeYcSyCh+Q/RFXH0g1xtfaXDNV4wS
laDQ9IEwu71rYW2HccLGO1soTJL3px9EuivuQabQ7D2PhHWx8ffm+8XvmYFtP89p
6gFjg3wzdlaGmUNYzjioCDzdlAykYCbWBj37KW5T2HxI6/Sh61O40P/EKqSzcv8+
W7xWyDdNC40s0r21TKCCUf6CGCx5ImdjPPEjyVJzgMoGCq0S7i/Kac/0mYU4OcxO
cWR0NCTkuXaPUAaVTitOy1T7ioPzNmADdKek5OMuSB2nVkRpVsoqxZISFB+7/MiI
JFjAzdgNFjMVItn1nXQV3m9H6PBdCBjvK2SSVtARgNXdrq/N5/vLznYxRX7BaQHL
NV4KkCMPFn721qBs7Ll0FrB79GWKkqKlL0MhnbclBCgx/d44JNjYoWsnJyq7+sO7
ZlPVGloZggsFVg9BheVnVENXMmNNqcC3MSScqT7n0eRXbI1hcX6a6/sTT8u+Hr+n
2neOhDsT82ZGvBwV8AcdD3DGxlCeHxTh65CwCUfo6jfXHqpUBu+/+cBZldZke6j4
9CzLGY2f5CrWefhtaFSQJYc+iOYvq0Xk4nRrpRIMMH6ZzZ8bMg30lABCS9VzUwoP
REP3tgDaGzT7SgdVN1emSG2Rc61fG3hDujBYJc9JElOOjY5wQD6J3EWhxXbk5HnI
mzcg+m2C99rPkWHpsdUM0qz6r12YjQTHLmj5tm5RqgwOsVcM/mCuxkvO1+XzJ/46
SUCYdcBWeD6f2TxBnYpT1zngpe4sYeVEV9tdsnuVxCtz8pD5TKxHKOAhdGPipVqI
dnSCn8KVDKLisJD2e3KQ/Ju0sVOuR+zA15cMfk9cg0ZbTKuj1SfqlVCDKDf/yhkX
AfNXAP4W9Pg/Ldx3JSzLdhcg2jjixuBai5C69T78gA1+//mM8ZAWKQ8evdEcJ1yl
5zwIwVxOatNkZQrUJqXbx7hqmlumYERSeFWWF3vUdQYEZl+e+Tb1EBpNGh9xqcer
QqYx/LPgG151VuigBqL9eJZ7i3aBIJHUleCzg/lx5SaF85/TL2jM96ib2OZBWFVj
0/jRwh5RQJteLyDZcr0vsh/WC1YC/FXUWcChqavCNVo/wk+BAcV2ic+5ILHCyYk0
xF7emgjyNVJ2a6z3TlRs5x+v5Bzt4HThW6exsPUhil0031ZhXOwgILWRBhIaZkhl
ThPfsPg79bdrmglKcl9uuRXv1mjcbjZ8/+Ygu5sS+Pi16f36xHkSP/NETznqDhdL
e52D+IfPiTWWrn3es/oixFzK4KXulEoDIRiXe/3Yo5chZDyHATfHZj4aY2Xggyd5
pDf/hdSRCgmlC7R96+9PcU+G4Y2Srwz1xEils8mcbZgJBzmVkH8g4+br0dSpKGpR
NMhVw3oeyG/6hlbnSJix3AmkZr8EZ9XxLN+LxZLo8VG2L75AGPzGVQXQEyGFway6
NHa5+IEcF/EUDwMPUFN8nvp/gRn9tsR3ZEhOkLioF/84QMHopKRqw9Ro51tQoYso
ZHLp2sNqYWJtEa3Hx+u4vtBPAAK2l2AYrXdGbmycp0qSAYQgnYPr1lFZK/Ahaz5q
JtzrulV6poWQZMva0Krs55Q0ecru8mDN/FS1GZtoDsazt/pRDGsvpx4q36noXL2U
B22DpVusvuWqkJxY5URf9pNCfgRdG+RW83y9ZVxHiDkIIU6rdVre85sD5KQVoe9Y
kr/hdQulHMh7ODGMHu3eV7/KVIKY3yJhG0h1rTiF1v/L1/kf/dXPO9YHioBaWKRg
TyBCIBW+GMyyG87egrc14AZaHKNwDAODSlSulykkV6waKYCj8N0ilQlNYhtNPjhG
cYAsk/8O5RJ5nZALWtqkFHh6blYEbcL5izXquFhe7FJ4ElTHssEy866Qt4XgRAmz
snp+YnNJKiMCb89cv08/wPd8n/69yF8AsNIZ5nWe/jzJtZao5jDpClxJvl0Xypwk
82LheR7zoxgIv05WL6mdvfnJ9YuPB7uKv5d5OjEOwLWsTDsLgAMXdTY93gnoCHp+
Pxv9evy0whdj70EbxnPgL7HUOJ3ewvcoTHwCx5zAjr66SIPb5rVRlypt5al/yXDV
tZ/YWlA2OL3LF1/o/jLT9yOAokW9VAxcPt/FIUOm5ZXmQS3ExwsI/a2alwvAGSUE
HOUOxsuXRijrE/PZBkvrePmG/DSIPfauVQkDSDABDVVGFrHic9lnsZ4dkwxpwi38
apQJCiZX0Rd/tLr+vILjHzb7WQNXtPT/VvtKpLReG6Aq9Y4a78suCyMEvxIswrEB
WLs+GxRDf7aRPWyNXpb8SQo82nDqkBU6lxX2vW2KtbehPLa3V43UdSTCmiuUbRkV
zY6Q4JUIFo/OaOWBqnC43i8nOjGuelxLPv5P0A9pqZIHXU73Pti4QUMar7v0aDtC
PTgnBU5R12JmKCVlPNIhLD5iCmjCQZ+DUNwx3COHM5Yh4FBM26zViPQUXPT0iyxe
ysZLar6W3uujFzhugUxdiGQXH6BXX+3jomH5KHZoUty/JD9yi7wT292MTOtiTYU6
JLEjYKv5h5OGxOd6bnoS/ukOjhjEvNGAej2+PrMD2Ub8znCAGgbllA5xO1G6+fXR
nJK3UFpMDUf/gvaQfWEgPsYMI/J8o7jYwDliRNDtDcq0semngvcg8UxO2o0BYzeC
GS6UDXskL931rz7V4e3Jy6CBdMCNzRV6ZEcjCiMOy62G5BL9e7gv6+vNmnQDHU3b
iJygvlzZlXZuacO8Ant6ZPT+wD9xSsQXtXaK4zLuWbfKULz+yawvRW3O5bBFT3Vs
jNlqPFX4ZZvW7emitCQW5B0CT9nzGQq4CiiX2kzlWOvGJdVx/k7GAoZHtu2P7eY6
ZbAL4JHHdPVWhJfnbSyXEl15B/Chiu57BETYFVbURjUk+9iS4RyKewVWMIX+Jt5d
63A28PoRTmZaEvjrkKez9ceMBJudX6r9iPJ+VJe+GUbssUHYq81HygF+Zs9csm4m
eJcxpTRP3jYxEzQ3Ix37DJX/Pv1TFneZZ5RpD96MtsAj3oajXcqslbHe3jpkAQLw
Vikvks1P9nO4L4yhlk0uLoup2s07WEv9JD60Cz88fgqIw5T+OnXsr04DHL+2aNOk
1PY3n2lFfm7PAPv1jy/pp9J2BKV6HQA0IhQllvl0RpKVXNrkAGZ84Gvi62wnvUx0
cZkncEo5Fwn6FwKS6BJEjKF1jAConXVSzvDq2U18Y1ZlS7VQHOZY5O7QLP4u7Esa
CbUH7/uObjf5ml7WscG88/fZ3luBhtRsh1MHweSWf0u7/lXCFgC3a36q2SJhXkUt
737I8pdYR1RX1FVQZz4j8n1GzrE66xDx+zeDE1VtXicgmaiJARluEMGZaodiq3Y1
OBF564imH5GxRZuIVesJ6x2i1VRBsXuNtA/iQ1DZGRK7dMfGbNZdBYhR3ngkJBnd
JYIEaZwSJJscis5ncvRo67wyDcwH/mfeTAjLFhNeKOnLW80LHtJMDpaSm+mGTIuW
nbx5HPHpmCqvrFGwnS4nSx/B+Tg0cp2oz3evcjMdZyIrO6w35Kjqluu/Mcx6o1NH
9wEpnj4+YiSVKaWBKuUopy62ZLEy8SV98wV2F3Q07MihXMjAG1HTqSPRJsseYJr9
8OsAFaP8qxw9lSZX/snhFGvp69f1/+Kxf2O7Qv9z27cd0tyDvZQzDwaTaqtYlSi5
CXP3NirP791Z+ixnwqoMci1d3r5PE2xkUCgQlvXZvmzzUYabNdw/l0No+BVqtq4/
URzutyeEPJ/i6NjDJwh0Q1XsgnmRPM2H5AUACS73ZyuvZJPeq0lOgMHqURKHoWRW
m9GjxneYBp0gOyLyTmgLPhqf8lIQ8qOQ5r79dra766HzNu6/Q+q5nSTlUonIntCM
Tcr5G8iOcPP07A8Id8msn6r1bKn0XLrFDgqZclHezok7LtlPLiHlCT5ZRiaHvWyg
C9hMBkBKFhnvK8Tcq/0ELrkIIntiHJULUn0SgnaNKu91y8APUjVz3ywnpAWeIdYE
nr3lmz58KO6iHUSw/BCvwG0g/E88flIX77sImwF9YoyTiiFjpNZEtAEIhlGy551l
JAZM8UMIGv7vIyrEpTD8/1y7r2FekEAy2/gmwEgGgDbWNOXpu+Oi68jiwJwJ+nK8
mAgHgOijsgoO9AW/JfKZupJGWG11DHfuXew5IOQrby1OCpCi5WyKxwPw1Dwj+XK0
gwLlNWUTB5mdzQTr9uyOMwKFhZxFetRRDOL8QS1w/PjmNadEFCzaszo0+OUVoStm
ft7fWaL1ezwZwxjfsFhyK8CxUhShBkprymA+w36QdSVSpXTl8tvPhUDwVAhtezds
UewQPH90Zte07GoZd/XxT5Nxt62WzbvS68oODkITA/vSmJxD/a06oKCRfeRGY8z8
TZMTLTZM2PLYmQyPSs95d1vzFd8IQIjhtuXOrVFKqqIUZ37yqMsoNDgg5VW8z62l
4lxQP5BIJRI7J/YSTGIFePg+DoMKX6tl9WPSTy8DqKO9r7M+Aehnd/ojlpU0gmbZ
/gHD7krdwsXiPEmhLshX5f5yXnFjfDc1qlx8b/0gB7xLtjzf3S1GZ+Mz7T9UN5zH
0JBpQBdqU2WvtC59flY+iDqn/bZyjRSUdIeNcSRbdJBsMcODd3cjAQrs0qr4iORv
HUC+Mp9K+UKIdj0BFbkOcmfE12EsI7zwgXxTFzykD4kpZXELwUysAZ9gmoGHqJab
ZHbUFurp65DlP6DB0sSJiLGCuq17jFESfwKKxDUSD3CXyF81u9qGo5iM/lDvp5oB
myN5YV9j7zwdjITkxWWq4XQPVSZwJCIn/rVJfHP8zbS1TRllcv5VIFb29Lgll4dz
lgWxFT8YmWPIEWAtLWHv0f+0pHl55Nl5TWejcUqUtljbU+mUK7GbywEZdFuH910y
b4CZXZIkk+ZbM4qs1eNdHDfZ6mtec3r3kO1IwyqjK1wFhLr/DzzmlzGk4r7m/vHu
NGy3Z1rzz1HJpXhdJ3ced5I8pYfW/RpT9toh8GodFHNGKSyaXHRPZqOrYznkdIOc
zrIpAcL0y497/fTsPP8lm88Wk2qKrLhllLyZrO79JXJer7n4XzTTwAvlx+2EzDcr
hPWfYIz4gpMLwpQzxNeWqxq8C3UXNavRq/FCPLZx8S09lLuFxfAfLzjWVi+uCMDb
0c0XkZrO2r0JEK4wQeX6Bu5xE5QRr5qe6wZwuiyxfAI240OeQvjE5wtcNdj48Zkq
J7AYlKbeoJASK6vBysY5W26VoNJ1vsWTLc/4h39kv4HuA4w/UIVUEJjyWExLl97i
m729Kv/NvgO1WwA9lTYH68mFne9xrvnjeqYmGZSAP5t0frEMhGXcc2fcJNykQSGi
wxJrzhJub5WQnyM78JVnBa5aJj1DqB6X2HZKVNCuWpbuwHYPrvnJPIKdPBb/1+C+
DtjNoiyszbxoN4QCPo0I2zSl6+gSKA9vox4keWGpva2l7YbeVm/itwhYFJl6zPi7
AwtKjDHOlPrd27PamlfFMzeK4+mLJaTvPos01RJ5Vwnmh/2oO29WKgl4ZGjeIt0D
/i8FnsufFqdKE5EszIJ0igoLXUNgGyAtaJRhfkTdibOLv12TEKfO16ugVP3qcpZ8
kDmMdLH4E8r/UA22DYBEntXOwD8lxJSIgikDOkSDQUBHREaTYkigsOIvD2GBtRj2
12Z/OBPZVJshY+qt6/Lra1U9Q6PlXhKrJQOXG6uYqgmw4CInJ1mucrSkizcd3aAW
FwEW3wIWzUMrgrFd3DFulPJ0+T84MmwuHznM0ZYXMg0tYEOYF9MzxGGE01N+D+vn
3AZg30Gm8cv0y5IdTwKG5tjgVQ/F5V7Y58JOTZFB8fyQC60mppKHuYY4FQEWZlA2
fOxsZGOJy7dOrnky0ddHFsAGWK24DlCGSHjNCN+C7cOqXasgJfO/HwMQS2DFgDuy
XdQ0IXUpTdf2TNF/sHr9kl54PYVaHZFjKGTkVY525EGR+K0EL2ovjtvTbVW4/Xzf
mzt8WQf8bi4IfAx/3RUHllhs9zh2v+gRYCskj2q7gsZmWtty08XgOAAdmTJ5DqQ0
r3EnCo+S+X4WVHLCukg5lB6u0YyuDPcYEhKkWjts+h8crbg478QnD5dfOXG9AKSN
LmetCxg6J3VF2BTYjQRK7XDEn+PWExCalnB90tB2iG8/ChOC1MsyYqG4Z0XjusTN
IT34k3FR0Ti45KvPFiOly95Ie2H7wx081/FHTIvUndgVEK9dsxIv/4wm9K6/ec6D
5zu19BSfXTilotua9HQw6LsC6pZgSn4ApWy9Ye+hIsojwyo2ouTyIWFiE0u2Q11O
Swr1a+s4m9y/w+LIc3yT6QGp37Jhokw9IuHgUzJpVxvSEvpbbcGbO+8aY3DMffHT
qnCvpVnD9u8llYaJosJtN3KJOD+rrf3J/bYE9+OT81qbB2G8bASgUgOImQdMH8uM
V0D1U/O22nh2EsrZob/XBSFTRM+nJsuSqjxE+fl9jY2HR5u0eBnFOh3zMy2neqzP
AaBUTM+Ri88oAQH/uGWF/vL1gt2LQG08lCtoknruDSxwsfb7FRjJ3vBhgG9qoZdY
sh1mC9RSq4ZKuas8BkyPz5i8mGSyUN6ZVtieO+C1mdHWMwd1Z0ApeAMhYbljjfkc
DGDw9fBpTgu9P6481UF/f+rBBnR4etRxY/lcHvkqvyBF0qa60V0UTQrovwJljKE5
TAMRTFf0XkZjk4KQ5aR52Fl9M0/dFxAp+ooBsqQSwqOPCbvzRJTzByeJxmkA3OVG
bnfKWD6rcM1+h5mIl/yPGYLG8a8No79TsSo/3X9QxSd9rpT9tIfz3l6w+n5YQ3Tz
/Zf0SOOt2VoVTZSgWa604p5E5t6hGvMQVOXg31ngg148rdWqIHr94wt5jLoBLLNI
723MbST2Bk9KyAtcXDQiVSrqXrKqwXzkD/xUS9IqIbzBXeoEZR+nAfq4PUDmz79S
iZokW3VKdyWMgsUJYIenGtRCSOo9+FBPbTW495pUEDmJYiDL1hOHdMTxu6P5xWCQ
VvFFvs4q9Isp96HwDWPuUsWFv9v9gMzmkKAbvNuOQC06vbz57txhLSHq9VLSiA3R
RCLCcWU8z8Kt5SzU7k/cuKia0ZK8JURictf8SHM3O2dlK7QAGDl21ccPDdHY6oTu
K1ZtRfEV9MZAz2pDkfe8A+3bOhLJeY5NlGQMbQVmhrWYXe7Upbw5lZIc9b61FzV+
tt6JahD0lbSS4LV4V2lZ/lYOhgjxjCQV9IBpq9AmydD06N+yNL2wNYPZsoYVnhf4
3Uzqh85Xt+pxts+bOBbDF7zCcPOPBiJWEteXEgMj6eRvIZ84esQYHMj3RMSvOarr
MjSm9crIoP2eMRnreL47YJGcbyZhfam8rjuefEUpzz6U+NVqBNYiAjgJqA89oRvk
qxFxr6bhxLvgdkTicNxskmn+QDjkVoy4e+yRmuK3ZgctFr4n8xGfGKfQ7N2Z18+1
lOwByMflEl4J7yosCOqGVlrQ07HorHlcEFqTStRkAC3+WMvcHEG1EEH+rrcUDf5v
k28tysWVVt0tkjNKsHz0bDxkH/0jAXRPeYFMl+86R75+cwZX/GFXhZLbdoEt2nt4
RjcREJixPGbTCOiEnJDPvZhXoGVp6P9OBldY9tdZLfdiOr8rjTLz4bf2ygOfZSsz
/OibmnlI5Afb1oUvln5iU//jiTr/Rp5TDvtwEED+mhQbuGL8bgTmIqKyn+RTdn4K
XE5+U6q7Iz9T4leF1N/50pXz1Ed9jHUSntbl56HXYpDDq36rW9uhLTJNMWAF/m3H
sF8oRolwj30szJGQ5vQqHIqxxf31N21IDz39yxSIcvaNeT1vnoneAGWGJA5cNqGD
boZvvf+PFzhu63CTI4MqnqHOVguAcbjleu20tw0SzquuBUAaXMkJZd0MbhpaxQSt
vQJzy3dRYULGE84Ixw7keZAJtPWfYpsWjJu+WREtIZr9zq540eccNHAMGhXCx5HT
J6bweiEBHS7Bqw0oZWU9z6/r1hq6WQBxbDJkglNglDgLb8Dr2ZY1zLHi70n39jgO
0ZjxSSVe8Es20KUalaX3CnQ7WLp/a1RC7N/pqVWr+SCWrHbBVG1wUg4R196MuRdT
qQAoNhnFnprdFMaBk3Os2JGYAxxUcMtop/SzC7mkdobs11ZU/ZGU6T4uoR6SGgLS
9QdVr+MhEXTx9Yt40syTzJNCz0JmZUY4Y6TUGo1DA8p3kZZJV8PJrHwLN6m2/0mw
F+G3RYylyvBKdVALeelooR+flwl6kOEhkHX714/zj4HBqVA+9NoQa1LOfLeuv8dY
nDS5Dm7+GgMiXvGj7j1QmWVJQRRAyaorDmflc4M94WTcSUrZ8LbkEBaBbE8x4NB6
iDblVmSZRO2rwy5ylz5VOO2mM51QXbfZHTiNOpfxji7Zh9415dUND8UZuLq2t+un
DxRlUi8dB6VcaRpVCust1ydLZrSE3spATLQSnLszsP0K+X68/8uzBUAlKVhyR8x0
W/0vYUsvvKZ4U1IZKJwVYz65kFXFO1cgVKPC1Fo920/wbqrHpVYBBLOTCtYNagp0
zmQnmwwVFusPlAEQaZYv/Ywqg52xm+JcCiPE8w/b2zMiod0bGhMHRSqjbzI1RVUE
JZ59zAxXumKzXHT9OtqLE5lQg5Hj3QroSJZ3M8Bf0NxC/EyZ5i/FRvmf05RQuMUC
iaK5Ttr5gwsTB5AX7uR0tJqQ60SWDdiPz6k2amAyxf+8rxD9EBuGSmgbABtcUQVx
IA0S/nQXntljdZ3jhcyRC9M29wxiCclqpStA7LPKP1MmpqvL1v15YkTuxlfgJiq4
+yYYoUnCCRNTtPT4ID79C7MwvDGDtgbM/asHGX8qOULC9PuvkmbZCxiRYcmKNBYh
237p8cfT3BMYfKxaBET2L5ya5u0BPG8joj0vAL7XSatPc/crWPFUVl0WGFBBQNKw
iVmM+Xx/R8AsbnBbOs4XYi/ETkYfiwtkgGJ+9451tzqajIwYsgtANkhkK08hfL/i
6wzTxZbFnED1p31jZD2hFBN9RctknweG2ellvgI6Tqw6iKzYMBK9S8ounRhRFptN
y147A5RsPQwkU4HiZ3XHoHOxy9yHCOzbZuWTb3IM2x4knsrPc4nP+6EwY4e23qBr
W7BaMRlW5uDQixmvVdMZeLuNxO5PQKGPfKMoZEUFjWod9EL9b9Ex55xIJuNeWJ9O
RYFptBdSko9l74dtKdxHzYlvxYY1IGNNxkMWjItjV0q5ggPaSEy1xDRWWccZ6Jq+
w2PpexQT4a2RLOuFmQm0peV+zv1LnZ7u1x4QwL5bOwZGSCWdb4Bkupb1d5OfMP4E
O9iqM6NgoQjIC8SjtqzX+qdDLVrRvrvGwq+u8j1ulfTMrUcgQe27sP7NT1j13fJv
2MEfhFnszrEtBDPhIMikhn3FEKF9yzNo3pZCB/l0QMvclVppYJLM2dtCYRPMIRnR
vKmIO4fwiJPARrFSV6dcNs6Gp6q5Wn6tdyijKYnvl5uNYetXvxsqElyNiP9lOVPu
34QjUCY54MoWvFJqznYDjaIADFDyvdxjG8X4gTqTMP/VhzA3SEf3oxMOEwYFF8MR
IepifDQI+dFYGFFq4zK1Xg7BUAxf6MeoVoeqs5jZQKef3Fl615nzetwc/mgscDkk
td9O6QdcN3XpjQDqYAd0f8TD4Vhi2pB6rknFeno+flsxKFjeBBIytXbVgVtdAi45
3MJcQsdIP2KnlLfb9PGECLAPi8FEE8RfOL3WmSYo3Wmw9vNW6fU0jp0seFen/ZdX
aBmYsisP7WZ8yyg3jS7cxRpKjEas6CMPTsiZUDZxgUHDfFJPX8/YvSxPPELVLeW9
s0HqCVJaXBzIehbjHgXvwMeM2yXzHqiuRTh6hPg8YKEDEUi0e60fMq3NB7umU3QW
6HzGGfPNFuCSfVteNyaPzOB6RdvSWczsXQQ/+Evv6y+0Oy/Nyx6Z29i+ox2PjuAs
RXrflHfpzZq46lHQbAhzzqYfE1zzPGMicFXVK735BBaaylKZ1UscfdDh9Jf28bNA
Rqs0lFNVxDtJ6AfyEcMC1mqj859O4FuVuZt3cFSq6+j8zKduuoBPSXBGMRBaV/aK
/qErSYYcih7cYJCaWZo4g60foJvrlW5ktg80IfpbXYxujMsvNEPvT/ee6A4x2svF
kiekNPy4url/yBTZoDum7zHqiaC2wEgu3dEfhTtRrxqz8EGj8m/cbJSQR41bPf3M
UCTZ6l0aXdkoiSmGagSV0Z/nh+kosrzQB7QILXhlPbxH9Fy2naKc74o2lowGcAkc
IyG5LA+M3nvyBlFr5+63Urx3ygaiuN0pgaXL0fRZC059mT268+zKMUC/lSxH3NZ3
S1XCThzz+6pzBkyTPfy46CdR3+aqpJz5iBgJPmy5yOafSner5wQM610+qdMZNXmj
rr2+j7WwclQJO6UaXE0clhq4hxJfB5ixniLI8i1ykN7BZV2BH9Ru9QuPK60jo/aj
MsbJEU0fhJGVcWf/hXX9AcwLzBpHzKwHNiVvpKiPLd+q+bzo5wsbMfs8a4rcM2xR
cIk2Fu2U0e+PeBVKVCbkyxy+QVZxBuK6BkWHBOB1okCQuyv40la3NRtQQBtLFMWV
nPo1/SEeqRFhCO7WXsURZ4WF/REzFUPmewtBEUR46/HwuaeetJjxWQbm5DrZ0v0A
KG9zGQzo1i7vlqr9wJgZOadEzaW45pRRVdoR0aj5x8EX1AdXmQ8/gd3PQm0PN4jw
STrk+I226cEkuKeL+GU1GxhavdyDhbIUu+vnP43+XwLGc177btrpBtIaE5elWuZ9
XuPWQzLp/WPP2QQmX6QbUbS+zj2c7oUhy9dAZFKM2NHHXex2YQeS9NGLMRA3CnCz
18WllSpuKQLNEjlov6KUHsEQf0afCnjOxEq6J7mrWpYb4zEAFoU1NM0ZPX/58OOF
kS2ljuNa5qDPPorC/59Ud46Z6CAwSe+GCj0lDRXxJAMw+R0JHdLHX8BRX0F0cNeR
M+C4ePyT3NWWvQKCWla3iJ8HSl2ue32nwQX52hJnt8sUfpb6zx+xiDSJmf/G1sh3
V896IZt6gFTAwD/WjbH0OJWGup2ZImzhxBbSnOhII2xDprl0eliY/BjQY5Qe5Ekt
jcnR9hHGYgnPw+fJuAJr4BZZELoWv5sTEFTUMyHGATtUiNbGlkzJMLg/7wR+NH5C
w9gD3Y3iXq9v1pyN7vg/59ltXd4XZakv+e7yY8bnai2Ub3RW863zFkGsSqVEGN1a
TnzSBv50pJaIrYvzjOOejaOMAyrSXzYA4yA3+xfeWYxlJ41v1RdAnjodQLoPDeEL
x3RJef/mlHE90zJ6f1hFRYDh79Fbbtcyehgj3pIatHVGGGpUfXvYzpkNQdb35LTo
nV8KD5gre1e8PNtZecvCB8KmBgU4j/N01pSJ87ahyuxTPsHIWHmtP6bl4gOkRrXG
SrDLLAY77je4uI2FgZA5wnYK9FGBT/OQBV2ELJ1SMeh9JKf1cw44KuVztvW01F4e
1dkOmzOxf6uDSCPVXULFGgZBXh8COsEb6aoUMwbzdfMdsd/hi7XrRrpBzkJs8+yx
zhMPFc+MsQvNzcfsNSurM2F3rJJshvJjHpK3li98kWInnsBkth9Ae4AS5vE0FPPM
84gKNHoiPZX0udaldt2/fQauWH2nqZyHpfrEbjY4TmxG8ScQN0E9LWeUly+VG01J
aMWnUwyKsoB/jYgyj9f3xQbNW2kVX89vppfQZOd3c1MKDRJOFui3Z5hdew7K1Hdk
S4G/zaCUvTZAylShTsxaEp4YdMnqCiMUh+7AGcJQQJw877o+lqKPOR1v7clyeD+l
nsbSjGZpLcdrLeEk8qLF5TWnou4wTf49QUDE3Y1No1MF1ofigWlXYvR3NHrEhLIc
AsZ9DI5W0na/4aFhDWsyjpkizzi7zAZW9H5wKFC1FkA3og7uuBXOt5BbGKVv4KvD
zfGS1LFhXZTxgdFXQGN/iiZY01GueeBhx3SJMMbqfh1VDM/FbZ52FsQ65ogG6qsk
FcCLXAeHHhVRwqqoizHlOkVelASAJQ9ca5uEIwoy0WhOJPEcPLUJF20bpLzGHNuX
DSCWWfcHZ5jEJGO1+9O+ZxSGNfvr3nYp0Ni/zAfoM52i+xSYA8CJcBzFt2JM9hLz
HMV/kSvZPPewhrt9ff7CnbFEfKd7RiVOxUCwMGeBZgf2ECegdINO8fRFxD+NVO9A
tjj+g/qeK2loNnC6r2TdmpU1BqjoidtSNItrl/x+jjmr5swWfQydfyvWi98M7sCD
m3Wnk3HPsaqTZ+wRp7Z25OH1wmPD80wXCyYB5FJAOs1dG8i0k6Gpp7uHDyCI95SL
zpp1e32W75ZWx9BjXty2q62ZtZoDsgBOeGX5+0UZ+ljaIjT7LGE6Gl8KY/GOeKQF
vz36rFC+Gl8asXpKZUvgnL9TcNxceFabon0h7iuaFuWT5+E2hyX3K6TdW12KVyFl
5WJQE+U0RBnSdhn2hkJb16pjTozDkBclhAhViQlGQR4uAUyPdoTyZVfeSMLE4gCt
tR+Nhv29Y1p+iOf2ZgyuzjfmcdzIz3IcAgkbGcwI4ftwkhvhPsiNIwjxalW0Q9Bt
R1Rt797W6iwGZB2bc8AzKaDSXA3nSjOFLKJrRoRhK2hQad/CdiP5HN/vI2DYmYzc
S/7lXGXuZsw9l2XOkjPnCKq293IiZMPOd3CdgJOZ6b+e2Q6+Y9EiQfcYz38oPtQd
RHWOwNUXiXT5O0NghAsA++Om87OC+4BLaljUhiSASypi8FTpF0nU3KetgLSghJLb
nRcS2J+71jZs4P3VFdBrJqAeD+754RtE8HA9TNqiTn2ZKcsVTFtS98j6ROrkTMwC
BKLau8tAUJp7P22s9KME1B3ievuzT4vkLobVRZTui++O3ljR88D25p1YR2Qbm8NJ
3HvH8VZSUpmi3e844vRLMFkBpCd2K2M70WXmwH5APq9jMJ/WE1yV3V4WH1QJphxE
tzA9PnoTkoV5k/E8punPqcm8QTaFgwuxpimMe5auecEjO+D+XeO0mgdNzxy7jIVY
L5FSGRYGkzAuk2rCYw7XQlLjeO1E6vcQyFREl2TR+IshGH/oAhnWUuBtMbTcibNB
GESSMzOmtX//Fkf5bhrLD8MhMQyTMnzqxFp8SgXPDn2G0SYLjuSVhsusUrO91rwq
YYWoPWmRgHVlg04f+OTUTd4cim8bSIzPXdyuQHedqy99rq59TMzfDrImyEmXHXPF
DE+w/vbJ3u2F2IVAPspR1saL3Ymdwjn1HLKid+m96kUQ8tjvomEmwgyV7aHm0UTF
dnjtuWDmzoDJwoxJxsabxeY7dpKXZ/L6TJ3b7ovL29xcH4T8wm0Uw7bXJALxgrEP
dg39nKHxKij616fAPUAayJAe8s8hdo3UhF9sp6d08bnMY9CABGGjSG1xq4v8Rmd4
YMXYmca9d+AytroSKj2HF5XExxxDVqdQWLJ47Xawo33Ub+FIDkBrG/46tyBKjW8g
YTs5La9SpqKWTm0MsuzlzljDHxYJ2MokM28zdrxuQeeKoBfYX/tgGQWIbo5A2E3D
3TyLb7b2afIssk0vL7nIMxT5uj7AkcWtZXrqr1RtO94ASrFFiihrAk9XYZjfKB5W
AtQYcthdwpt8faDeVaNFivtcAP7LtdZKoNaKNXeTOe7+/1l6bQiMLOH5lu9bRHaH
Q6KtDG+HS0JE/b1tQNkrsB4yeL4MGvbDSIv9j+fYOOHTWmilI8nTnxRf+Mcy3llE
IgZ0X6xjJWXJVQcbFGjcsB7VQ5FoqaAyPn9r1+ZONvBMIqsXeGilY/qQxCCd1bEy
OXLwcEfkZQRD7xAuXYi50FFglKP2aESVfU/GWEym4bFxhyg8W+9XiKmcavd1g0K8
PiklvN9SMLCodb+VlatOpfM/LBb8JkC1S8TKtfDR5fNe32qlpuQW5UBGo285gQ0n
62j/vkUvBf3z7D7uA0SoqBTcaeguKpp+Tds4I7HLXM3hefa+FS3ztgM6D8kO0kT7
CikTu4l8ZSTVBra03R6VOzBeyeMyk0u8RZFYst5SUvo64pANLTPd0Hp19MIG+K4q
CCh3Dc9GwZJoN4XvLE6YF+t+3VWSsPjNvIwQM4dBVyQ+ZknCf8UNBzp+syRw9asJ
P0sYfGN6o/HrAJgmumCAaxisZPW2w5TmBU9wKxdBd+1TTxj9SP2nWPAC3QhVETnY
7tO5WjQemAZVi6Mv5seHnIFog3v+GLOSOFmhTh7OVq2IHpPgWhnyGe24Qtm8FZJ5
dMTEkMEC23wg4/lCfyzofleWVuvHJG1bFK+gsgZCWcksSmopRG9UT+Blf3B7RsAh
w++cJnYgkc+tN9I6Ank4WUj90fKfoiKXbz8bDrTMBRGIzHWY+0MKiXMMtMM8fsXU
FZwslre+vEjuK7lKdJPj7bAO5oZes3/KiqLa5sSWc66QxMsvom4FcPecAgqNJA7M
59V54r5nlGXTBZF0G4z7Ii78CwWhRbupaZd3l47UG+iyRhaphvIQQuP57sc+REB6
eZRdNZsWt2jXx441k13gH7SsqwLvuVhhZvSKP58a9XAZg8vWrMjR1xsH+TQ7czNS
2WzdkpjBrgOW5ak6SJjNbk6lGEjiY9xyq6mOcfbRuIK3cVqPcjTXoepp/i9dzI2f
3t+J82wU3qjtwr5tWUkIJ2eSaTpyc+RU9czYkJ7ZFP/lvkbOOgL4qVnyzp6c6LPx
sNN8goBV4JNyTnDaaTJVIsBAdsXlL3L9CDUKJTyMZiu0NUt0RRQ/uWnpZ4pCtDJL
3hhl449cCMwcww7mWsDlQXB5GWAd+NYMbhPZTtrorkEvVqGeNQZTOtu0EUhwhsGb
vSGw72haF+F7Gc4ksA59NoGYPYA+H+BpXOkkSfKgT9lBSPuahXvzRHKvDEgwY5hC
FfEhzn7qNG06xBGTnZLDODSWJxBdLQ+uewOi0BAZj9AAdW+IWiBI3S2lld1wD1Ne
S5ObKAWcCYwiXqak17T92hw/2By6FxenFf6lZlHZb88nPDGmmsn75x70PQM8XLsl
zyTCmAD8qrbM+NRO1hvX7bS7dZdpSPVZbGLZyG/d4eOpIcdkQojuWqatbi52ZleU
zFi30DGG0XG378fqb6d+YXFFrJvbgLMpUxC5S88LYegIAr7itBflzB/OeMpoDg4a
B+Eb1/ALX3omJLxd7cbDG+31RlbxLqCUKzK0shjRTAVmyn6yILef+SrVLwdwshJ6
IG9pbEpToVM0IaWuiW3G4cSi5MVlFn3dVWX7tUERpqlj3P6nhIOdaC4R1Ex7tdjJ
i1+Q8rPuyuei6rDofCZqWFVdBR8y466lLkHr+GXI+ybvXyOneqI062sHvwcSD7yt
WT52qD/LiSk+kjBM/1su+2ULtDJlnPqcPxWiTwkSPPYAxu536thEaJMrthxbH/7S
NhY2iZC5TSJGe6kcF98NyCryDmvIvDOWI9r9syWLKKKeQ4fM2vi0NlsuIOSKTkVm
YsQa9Rl66lYVEJDTw4zAXDublBgaPFlMeIWnv9LRYYV+K6B/wSaK+lxPJVgFsh1Y
gqIyQYNqtH8T7hexAMXCop2LXw3Zy6YT2iZp6cVGuY5EeUi9tnfNI2E3JN4nlofq
1rW5PKPjS797hstZ4/Iu6B+oA9TDhmNV5+ObmHyH6f6W4Jnx5tkqrj+Uv4Sur/fD
Ygtqp83wJoJJ1t9jJhb6n9QVxlvzgl9yn65U6jmTmuR2wm/Oiu+dEt042RhEfljP
FKm9dieGN92inVmEnsj3oL24gOPl9lduOfwGSIOFttFye6jsw01YO/YwP7fV1j+5
GuC6G8TqDfzbZ2/nZdglouLwQaShgY5diAt3HbTaaLXmZmAAwsf5u1jQliVZz487
TUY1XEMU0RQelMyeapVqG9qyH7toEiWoozWMIEIux2KhDmRiKhV9nucVlT8NSD9X
g/cch2Vt9xMYit9/kwFZikL7cs5t4fsIbsENBXsXBLWce9ug0fgQ7aA+5Sup+PLV
9erL5Zih8AqIa4uUIwK+iXJRIET++pgyLiBijCDz2iYD33QE6PMO4K6V7KuJJZC4
RmE77rL+rx5DJdTo2KY9ecX5aYAODu7WmZ8MFbo8h7t8xSS0+Bwkp6qf/9plgYO/
s3h0Im+6Hp5vVe35Jn/+Z4Dc6vBWfOJYB9xnO6fY/kCZWIPIanL6EwbIUSwNCez3
WYMLQ+kQz7g7JyHxyAdLsNahqg4qbNKgMWCm26Bl2QSe3+y62uEp9C4GYynRbK5u
0m/6WVYkRlzGZCNAXtuXkbhGoY0QhKBYNAgLhMY9RjRrVMDER9ie6ZTX1UeRlbXm
FymYtjdzf8aAFxdyNbC5q+cz1V5WByCOnI2PEft7IZ41YbTs1nLK1XRduwK1nyHk
F9UO3ZD9CFVyulu4AkUv2477Lf9N7t5jSrcHsCjiFuxJakAlVG99kVmTGTbwq4/p
wHUammhpbH1R7WXwWm8LKOw+HerSLtVjmdmZNpKklgmHeeuf1OkqzcWOuw7VRSPd
CIvvKlrRuPdMPkK6VhOLYeV08rxx9XDbCRdxBdCvQVqMpLqv7Lsk/oSygjshcRCh
ZYz9XutgLr9NBl7NEND1tcYIcP+BAgMM2nUat8cT3yPzAityAzWZ+4XLBJhcDZFg
ov66ds1PzEv3bbLvaZFANHkM+kMJnjtNqFfmT2FeNUrvvPENHpNP17x8hpjm6wnE
DDhG0ETRH4nQANykxJRHoI9JLAaJkxEOWrRjE+QPo0Qg+VW7faPo+UwHpr5ZQdWg
75DaulQGT5XCZA+d0y5KHquGwL0FRGIz80oXI8s9irjMwiwL4+4tya01iqHc/qB9
NLiDH4GVAGVLbEuarNfrPS4lpUOp9Iip2OFtcLM5Jhy+O/loXxMdxvMTdVfTwkg6
KFZoneU2Qcyxv1Itg01MyjikS0/SSTuLV8rNmYv5zhgAjGgDTE42QYh8rjGUds/a
9INe25iq67j0Siy41Ro2UovUB2dpjXtRVA+tdDSvw2Gv8gmC4F5raWgIKjaU5ZfW
nHZuaCqhjKN5+atHyagV1aZnM6Xz6enZUHE3VRmFDNteBdj/DHbLPYAZeZHyxox1
nq5phNvDJG4HfrQ5dPRk2R5OMWUoqvFK/1pG8rMmYtx3bk8ojYEw9k+GDTT1qXRg
H6NzwQVsciKHjsOaW7REF8yEWc3P1EJyCAafBXc1gTVpnRQ/ZQp2RMEESPigfs9p
Rpv/NsN3BNUl5GNdQXTkyxLixCcHN5vB34qmcbRcALBhs6dk0sg95nzjEIwz1OC9
8+eX8VHM+4OKFqnh1kiRjcj5jr+mliXJTgxgV9ELNmW7FxVddzCZuHRyiK/INVGj
nCjZivMicY7aGhPqTSCMVvJwzn2EQJGOaSM6G9vVopzc7TldCEtuyIo1Pn210zMm
Gde+UFcWmMY3TZqWeTOjvx+b+XwBHf2F9OdSFTWPsP0pfjdwRIXaXPrs3765Q3X0
5VZP9VHPAyznTrBXWBmpaKKmthATeCSy48XOM7mtkcF946gE2tfnT+wAMltLBoDM
ceWK/bo0x3n7+YDYuHdOc1YEhPTFPqTsEncUBuuYU+uA3OY9l1d7/fSg36U5HfF7
D3+mHbZq+jP7BUvTS3G28SJvdvTQMA1G4p6lVtgkbLUAhx+XSKJ0O4mwqzBuz76Z
jE4q+/o1r9v6wE59C+9TfumFUKqMnsmGIlVhZQLzB7v+9yMKGMgAxURFqDEvI8x5
tchLgN/v2UgHrLFBpqxnS1wf8tiISaQADgYeyOWdOEeR1xyNkcVDyIJj41wY/XKu
XIbqDHhILu/CUlmnnGgQuZSooWoXWmvFueC8HQLw1hX5vKfrne4tRbDcQI26E5vz
VdHsspuGapKG2oh4ClT5Z0HxD10Ozvq5Cj1Bmi07npZYzRUjFDFiPXwxUzUzmIO2
aWgWeNJlSR/PZjLI4nol0X4rBxii2DM91ztCBbvuMuyXfWndkw66FqyRDURsZyBZ
M+oN4Gxqy5QECyYyhBIXHbyzoyhBmiacxJFn5Obl6ZOqXGnuKCjQYdrsCSD3mQQO
h42JZZpJRbeIZnqqFZ+rpNi6QwQ5O6osnRepzyQyx8AkIJ4EqrdkgtykRWalisZr
LUttz7ihS6dnv+FKMj68SN/mLQB6y3VApH7z/KCBqcWsSCYd3Rj+nraM9RB3FCnD
59/4ih0IVsvibu3GnaMEwxV0PSUrCLuDhg+WLuiNKfoLIhMB/7Hq7sOQLTGgsCFq
peB/3jN8aZW7YRVz47j4ylu8yCZSEkfTyqm/Fw6K6rMLIcXaO4ZFVt+4ayeRiixd
AC8YE03KznJHRTRdQExk5GGET6+CC6lD6YIeR2+o8TCF+EJZ+gfZ7B8oQ/GQlHop
lte+ogELJ3T7WLX5LHuEbWdDml0W1+SvErMzUMXPhljkMeLLrXR8qoQFCOIxstN/
6SDlKyAxOp7HQ2dSEikb34ndDNLv8Vo1+Xixv5GXyBAndwqFIAApb7rUG8NZv/LT
In9+QBPHsIy2fFraoDi272iG0krdbdqXmc8KFza3aG+dLK8eMT3Y61RGSPUSPPgl
5Bq5CmjGvRO5yC4D60O/f4dkDcX811f3yMoqwmsyBL4RFp4UbsCWMEkhkbApQ0va
G6GIXa/Zgy1/PFpKwvw9CeWynWIkXLEteNGx26ysvtH8VE+DI4COWRTaFvLkfFiH
gx/But6YN4WIpl26TSudei+1ECxOWsdYU2YlFUP/fvxm3YdDs88b/4Qf+NFi7J67
E7kPhrCue4eYJKEM3raaRimYvLCPXC38taaTyRlSJ1GWmwU9qpn5Fk0PIM9iZoH4
THN2HGm/qEE2pXPpUTXS3SKEFzVKtO94444AImpK2sXqAeX4xU6OcNy3rO5ApP4e
q90BHmoNH8Dltt6GXLCeI84Qt7ztmuSeiDb0/whBWrCx4hGjUFzNnh37uPCVCZQR
vtCU3hEiriAzaEnVSt/KZzIW7U5wUj2P5BgSANymeO8Uuj856xtE00KR4Xqh4LGJ
E0RZoZZ0gDBXMyHQD7GZiwQX2dJfQxBDA0mcjdyKP3Ccm5cB8g3LoWA2xCRQTn+8
snypTwY7kxC2jkm5HIVLlit3jzBFVmK05QlS45qOZ28MKPl3CGV+Qv/cicW7lv+B
xmzW5NAHqI/Nbo+TynKP9hXFLNxaXzZfGcLNrsua5zZqZwCjHjPlPdsMyc/4iJ4i
grq7XSIsOdxEKroqq0sNsy4pMDBE8eDZydx9/4dMpGz+pQZjspuru/Xb3FXyR0ZC
RrmCNbNr63dHJcWoyZ1jvGFaBRrLyBGqPnF4rABcmMazf/o+x3FZwZqIJwwbYli7
INxiJDeLjgjoTanZKPgYfWsvj0FADJ2l1AFMXNkT5IeyGRdpC5dRXD6ew11AfW47
tYGzT/TKaHZjmXS7QO8wKBEcPBYSntWkQKeocMO3bhGNGmQwrvB7e3iZk7jES112
3FrqTRWGhDw5chHCbE1SGnnbSD9SS5ZuhSEeuq3JEuBloW/7qBJ6jl+237D6jYgY
yYzig2uF1E/yUcDfBdxcEOULyJcRZmmERrHhCBNOUJz2M4beQrG4k+4R7SP7w/BA
hvGWtPZfLvsN1lwWzI7mdVyUc2ejxz4Qnrb4un8uzXG6zRoaN3073T96ySF0Ndu3
5nizM3kCO9LMP/t0H1XoeHpp4Q+/YlqL6E6ae5NJPC34IFxRxUj8UC3nbZAWa5z7
nsnBnbPFkQ3koU4OSPzrTQu2oFcoE5Qioh+8kodaO9FfzffYx8EBqnxC26qKZ5lF
TeUM9EGkD549lTSVawZkk7gR1bHAwW5hLah21tVi1YiCTY4Q8Mqx7eU4Mo0XMPtl
JD5aS0fDwO2EcH2l0dbFQtKzMRGozTJ2L6N2gBzmDEpk+6T9dP/EeH3mrHEo5a1E
stLSirnxTceFub+D/gJiRp2FPl+AN84fz1Sa1lGwwTUV+g1IGZ+vvhsXcLTfSRDW
w8tiA9z6TDdOljTEIgq/5C6I9L+HfdZVvdotXDddxD6oRQHb9HPlj9xirh0xH2bH
OzK9xIXA0HnOvrnzZOuCnuDDexXeRxlGDLBWbs4SxRu1f+I8jqsRt/CMzwisb2p6
SOezuHkztxDc0Fuv4EtP/1/rnKiaua5tTmim+9H09sVYnzye0CjymWTyzZX+y9OV
BpEt6YRcJ5JEgfOddcMDxcn0FCarsHBjL9fSfvjUE1eB4m8AkEzCQIWWB7IyDit6
eOaSqg163L38h17CehDyjGPIvco5W2ho69WepKSGIfas/RpP9hds5dWY9FyMBEhk
lotLd1AZ+oInWLNYRsn2dTfZEie//tgUcd47im4LwTXjRRZSs6P/GIQlvC/lcLbA
o4DBaoyCCPiST2JlZBnzWmpLB/cFdiqPWRgRwxjf0vTdZ64MIBWSEvga2RaEXd+T
mgCWBBleGqoEqcCkWoNtD7sOIJhsBSmGXAbdk+hS3gKNm07VNlD2wWggWBd4tnLN
bQJQnOBZSxkC5oK6Y7k2btmf3o8y19OO0p7PekwEW1n/GXUgCvTKzepkdiPdNuz5
TZ64ZICg//4IbWkEfAdqaJhp5bgXk9oL6yHezeATnyafxlSiwIPoJKAL0yK4fGCl
sP9yB/Qg7z6eYMSUTiKlTB0eHRRa4VErjSWl1GrB1KN/BQIFvc4aI+78U200RHP1
9cZOv0jyLXDAoktUWcyUImCMbDgWWOmY35BXRdvOSjVsMYFxn2F8Pp2C81X3oFGY
wkqY/JxfaE5+Y4UBNR0dYK675X5CBlV/qArKZL4JZnI9oMUzrNvKPpFheEZNCILy
kFfQuLtRPoCnBKzTWuf1tRf2rOfSiusnQ+UKDSt0hMCm1ZhduurH3x0xumk5lMDk
RLwVVTyoljAS8r746K1GRAAreA6xzezLEhw8vgB1YVQ5aDYUsVulzF74tMMrp0Y5
TEkeJt5Vp3+HRPigJ5weBKVf9694um1NW07Q+5D3BtInI7WUbheGGMlGaKFjt/PI
hjathwn0maXysdHfVcBpiwn8068opmkkFQiN5aPYvxzSwSaHrYJ+CpjjLqonMkm6
6ZrSNiaYktcuX32vJSNzfAvd9MarLIiZ+yXAgJ9EAOLADOtBtbSv949PpT2YeCu4
7vSZAPbO73p9LMddmlP3ADSitU6s1jtZXmrGGvOCCHVp1rQwPPA8CoJphEA1VBqp
pChL3bisVCD9Tvcirtizr65nMyIyHbipfwlHClRd7U/eGcE40A2yBA6qolnyWkrY
Y43B2bcIfbMM9fEEtowupwuPkbgcdxfiDHlxGDWd4wJ6EkbpdxPQFFjN/iPK0kdM
yGT3CQPT6bo9paLyKkwg+ZcStu+Yomdb6azj8EUYWT3AzMAVqSNzaA7o5fH17vKc
vlOD9wAmexf3NJ+KEVQMWlbGm649bUJw150GknTflHRF9qa3ozpRwtNmiR3ikEOX
uXATc6m4Z6DkDllxXyYIxFyU4jdUDDLXlL4Mv380WV2fM0qdF/F2ET0O4AK8vq15
HFvc+ALH/BLcB71cqqzT52jOBw+w/NzX2c61Uz/ROfxqk3G24qRqidHkW4XHdPOa
tTpESKlBbDwRRr/GDs93FKqtpPXMBE4qZESk3PcSAWNGuxmUAqrp2HS+vTGnFr1G
FR9b9K+ca2ynLK07D8jV0YbYKwHRuY2dA3KF5Y2MeaK4tKQW0i8/XDCV+JjKJ9QC
2L19vdwwMGaUMHBtTxKe2jRBdE7gjINfXqts+78aYeVdv6QSGJgo4c3zUzubfnCo
J4Zh8Vu0EUwJWmMRd2s2x+sEA9OyqfUzrRaDiDPl1O3yaHHHAHlSmbJM8I0LSNDt
PDidy6a1aHFIiJXDBgfaxstj0R8CvBBit98bG/Jo8Zkeokuz9lQgwt9SZjzu0xMl
2bYGNoGRH3iHAIZEq8Vq8B0FTjmKtnf5efhndoemeTWY46aA8onOtkFe85zfOnbx
rR2CmTTTadssAhIdEoI2NxxBrGviXfdDGR/waYklvPSDnsRpnT6ENiYbgy1yDG89
5v6vwpf8vLZMSFyfFyKhCt/3dekzsjj0M5DTaiCeUbUSINf9e1R6TYu+FiY+7oN8
poCJXj50UEvegHtTKzqEqD2WXVHHpA5+7LexxhLYtIo0N2vxTLqqCwSvTVJF66ms
/Vd/mgVIOYg67gy0zExPB7qoTwam3WUOXZmNXA/ogRsAE5nTE2Dhyz7RPFGOXFyp
qAkbLMymIyZxuoGSJXQaaNz6othKc4l9HNGySvyBcYUAT8UJ5FWAaTWFRC4lXojT
3ktNgFxZvhecgHEEtGtKObUFUcWsuc6fruIbVKED0J5CvOijpjjMl+/JMtczo+71
3G6HY5CbqZGtuKdrJtLVL3H8ZAXuRpKM+/PNOuzdAvkqQq6qD915G6j7zpyHMMoD
ifKRFuGDe/E2h8Fz9JZxFSXrrZPLj5VuAbrgSUw7u1LH4BbdpqAcwQNE9mFjfjwP
0TMkOV7J2iXTik06Ub7j3Jvtv1WVIP9S/9jI28djQxXeb0c4ZkkAuR47UUp9NruD
ni3N9CfBveNNWaDF+xm3YL7esbaa/N4kdYAhOhjNQYde9V8T/5nWEJ/6U32LPD9I
HBoCyJ8JSSVsl1LeAxvh44SNuGYYpn7+efhol9/qdG9+XZH8n52CeZuqvD3G8snb
xLKTIbqwHa3lHRr3blsNt445zXnTl+15QmsbWgVy1wNK2rH8jwortuu6rE6q63hy
YvbNo409O97gQ2pvfpiGTweirOGytLUiNag45t1PxEhw0Hu7v+BsrsA7cdCpDU5y
iqGI9WR0c9tOcKw4KWRpAJzlSsWxVYgra4J/eRKJKhh+vuGxLfYh45fISMtDBWOD
j04HGwWLBMoWMtBJP2EHpJoSBcItmkKVH+mo22KINkEUeZZYP1Tf83FbXH7onese
u4v14osIbE2Ht6Jwk/h5HUIQe3hFQloo4sIifA00J+aS6dYhTeKl9N54IN4l9Fq2
VhZ1SaqzSq170Aelwu8t6/S4/tWgcvbmxP9Cq64746FkbFdeWXScSx3pOE0wrGsb
qvDZ7bFZURnb1+n87deP3P+XpMsBgQVUaRu7oLUpIOce9dKMMgRdBBKKtf2iAKUl
uT8HMfbXYRx8YPxnC+vVPPPYdtkXBWAa7DrOB5gRcdvxA2Lxag9kQM5O/BVvI2nc
tvT4MCPkv1QD+RB7IB5ggpJ9CFJH1MBJwcsialUS0KyzTI6GqTyBgZs5sQG+bdQl
sDKkYGcKd4xQ7R8/I6L8l7YMdjgtkh2CqzRLZg8NDqVnuy+OfaxZW2Q/5FlNdwG6
EFT0FPOXz+4CyKFPczBFJrHuL+05Mqw3TMwfiqd5N7Yo5kjLBvW2YXQQNEB299tU
X75a1dl5VMwjnwJrIgLIFnNth4cmZGguM/vZEaKX0icxmGIpv+yFOjMLTdPKaSGF
sSEXQ7zR6CwQaXwvsNDILqgikSufpi0iimgH0qCdSw88rfiYeiXZCUst7y5x/huX
v//2QWodUaJsNkcsfkkTYak1197zd/BXMhr9kwJbi0AvVPf0BvIRXFzVXZrw8HO2
b7G64pQOKCgUxPB0a4sz1FVHr60zVXzWRFajURl7MtkIY0rPCzF16a5ubsjHRa2P
xgGfShIv+ozRRfk3brD6LzVPj85Rc80S+QfavbrkcinsLDeRFS1wuLW3I9OwnBOt
OSWio6tnaDziM3mIUhCdBZH+OuD4fkVOEOuk0Wf3O/mNPROhSW5MmHN1XXXHzTLZ
aGFCQJEPGjCurAdGcQsdazIEdrH301Sk+u5fVokXsrEfAaE5PHJMFKCY+y3Il2IC
N8mf3NF/tUEA0jUxIGUbkXRGwuiHay9pDUhD35rHtFsFIMM5Llb9zHFzHXAZX9xV
JZUmA3RGmCrVtsHQykDgQ7ydosCPo4PPmYxsCoECG40hDIem8rJqLXo/mLVTqTgT
av2VA07UMTn/UjEc1sLyasyV7OXQdeDwYzimc/V0bQR047yBbEsmA7yrcQIBoPgE
etg6ofGoafvuQK2FNpPs9pjlhrqgFTszIDwN1cFcsaKY7kkQnpWB+GbnabIBO7+G
hVSA6SXjMbSmbpcwv81zQg+UIQcOrXVHPI0TU/4oK/BVxGa5qVl4NgeKbyqRchEW
2U1uAXY6ZC45ssBdmLxcuUcFzl9u8ImrH6F1g1ZBpEMe6GxxmvURMjPy2PiQiA+Q
gDqELjqfjLc/5A5Od4mnVVSlXOq0VssKxG9pS1OZGM/5lEOsgsz1AaWkD7HtWFce
pNPOsOT50dLULuLUL9ZEZVShtpyMnp+66Qu0wGJBfSkL5dkA4p74ljJMuZZAJ4Ms
mK1GiYNGxDNfHIV05ZZ15PIpDl388e22YWs1H5Rboh9APl1cKgDl/TRtL8Vy/4q2
yZYUEhb6rzogQHqf5j4huk3bfUBkezsKze9Vvaldp35Id4HaGt+YZsAyPuAujqg7
DBMRryfdZWjceciaLqgwRVk2nd5U4/6RilFVdbAjyNoba7d5H0nTZashrzV6C+/U
TJnmX9Weuo442OJZybKtuNSHDUasr69NoFpNuRUoCeo4sSu66Dj7+23WsDIc58/P
fXe7TTLvMG8q6t1uDDgweb6fO5H0OQP3CYoB2loXXup+a4uqySD2oFEr+aWQRnTm
onN7utLBXf1BHNUJnxDuedIcKk70OiwrSmZcVOWNW8m0W+ta7osSnbI230Hnvut7
0FDy7QA/C646u/2M6cXHkw306BUXnBcSHOg+27Vux+uhdDD+xFyHXzwc3CiFPvdI
OtQmbzAb1tMTLabJxjtotsPg3Wp7sOmLbDuYefpfpYOvib7mbz+dFgWRLPf3pRjZ
3fhhbTxhECtF33nWPjYOAGf1WRtlDYLNlBRy/GyMDLMEgtvo2CgUvVXehbKtQkaP
dRuE8peCBZOlkn+RJuyOx9kESoj5TnOOBKV01v9LUyln2yaL9Q/mjT085gLBvmk2
az5wgtH0YgAy3qXwzjC6eKlw0oC/enLEotot5N/58zE56fZJJ9qtSVJh7dB3Bq38
Y7IEb9ZaQvMqdesylC/o7lKY9R/8OCwo2ioBy1oEBaZHp3tWGQD/r6pPDWeHhCBR
ArjSPzOozrSfai/uc2YxOx55d29vDIRtQjW7rCLZM53z5snoJx2uADb+/9uSG2wG
bjqu4hdF8kTQT9KUueLpatFc3s29BCmslB4g7uof2nk1v1a46O2FgKIa0jAETkTx
dggDbk2+qSVt01Xh9lGsRYj+uwYrjNl1wGMf5Ih2kcVJmjdXZHn1Oh3hoJNB5M+U
/CCqFSDamM3JewLfnKa3e7yuoZaRNf0PvCznsTlVP4lUhnyNsbBC3uq8Q4i+J1WO
iffy+0W5tlWVnjpGnHS5ugySPF91Ck2AtsKRvudtK6nNeV1wKjjLLRxXpvwd/kc0
WeGpZ8NAcJa/mZHU/e2DxGmfiwpCIPkIL7eX8cJ9qi3hKjQS3kQI+jWosIGjXVP+
27wE5gUDYw8FGRd6JJF0DN+oeUqSuclLN8s4pk7RgNNvylji9y7FPE8l8Ge8wvPb
tODau3r5E/X79UzN4B1Q3XMuc2hKvxwymmnC/kcNeJqwx4wDxRedbpyVcmkvSEuD
yTJ9nW2BH2rsE2kQ/aRMEOyAjcgWCl3Kz5iwM6aAibfbSHIENdgrAdNtC25pgPQb
0uKY/pmmjfgXsF3KP3OSjXMySooXtnWtyMlZXvDyxIxE5tfJNN4pMMh0q6oP5fhm
VCUBUE/DoGt+FLLYyDAAMlzwNLjHgK4pRwgD1476hHKFnGAHN3/Que+ECZqt+ggj
32oB7UQKaKlqyMi93Ip4WI9h7/R9wAy/GCmpl/9QZApXxdeoGrPzfpCSYhRy4tgA
jO+3Uocog5vMNIl6k0KTfF4cKHRvi1EU0BTPRnbqWARJeKEugBgjGO/UzogZbkua
fOQX21xqQB1htYb+QZk0qrl2QMF/qg8nJWDEyqMXC/zWMJpYcDz7JrmSqRS8DE7B
pMF+Ehgs2XYo9Gm5oF6Q6zGJwFRwv/wvgSXWSDip4tZ6uTb88s0ctjIzqDo/1Qhg
zE1JRRW7S2VPWwh09E+nGpPK4OSXix+cFeJ6X+xZBjX7HS5sRr7Wc2K4l/IEQ1no
eBOTbMFBjyKIKf06IcY4U3cHbmz/kP+bV0N3sSnN+7189gLVWCcFyMsmUWRZdqij
lmtJVOTNeTf01K97d38yU/Z25vCY9jrsY41YyK8sBLM1O/FlEB+eojvLcvXWYanG
fTdvkiayBUFW0nGThtwxfG3XrOlUGMbSDXfQ9tchRGYiPmYbB234ym+2ME+BHGjk
Nv6BLwn/ROQRX3ya7q+p63Ull0UqXla29fkPFV0n/ZE/QcTlkCzXHBd1hnnWCBnM
4ZNa5k9FgOU6wPn2UN6Dh0vm91dazRBEHJ+Tca1/noL5K/FGt35cuFme+iEfjwMf
CjSphFX1lAHcRuC9e7lDDx3zXxVPQA2anjfX/4c1Dv6YyH01jg6cSn+TWf2zSbi3
QdZahna2du5g9cxN9xNZtj7wUzGihfRtjr1Y7rAwr2L9zyLWECflcBcK+wSrEo08
KmyKSYxb50YrvYDwnqZJaXdQwUs9HhY3Ahi4I2RYo97y6QzeGm2S72kZ2nAO546b
4YDf9rNJakBYq8kLM15y/uwFoOQIlQGJVE/fDLfkhcTjThVQYHoVwe01kxqyLWAK
L9ozrwdHc9tarDtLgvcENEPaK8K/h+7bYCfbzjS9hd366lD6EiTY+ypfETGugmeP
0VZ4NnHRnC9IZeRJipnunIWK4QAgO9alNMbu3v2BRAwX4xnPpCgVxw0fEsS/tWYS
ngIvefUFTV36J+S0UqE+tEMtfqTEDBbi9Zii0EbNE93vDB8jPLre1gns733yYKS8
bhf4BCe+bMTXyMkSwFOXFMBjAKbIwmLDf0C4HtU5x9RYaVemo4by3DGsx8/jU5c+
jnBjU1sx++0pr74NVoOc3rJjZiAYwEz5u1lLtGGqrPXXm73dfM11H+Y+4H7yn2k3
TJfJattV+loIEV+HmzSM2H+N4swfggJ76bvuG/OUR6v5IA5SXSQImcRS3/sjyIre
GWjo3FsZBMY1GHYqnAoXOj2Oj//5iOmDL+b3/7czgzmiXV0OEy7i9Ljxc+kQDRiO
KY+ezwQpVJGykFnnRB1Rp5VoFZqkkq9kiaFZ05bpYZVrMhxlNTw4Vlm58BC+FaVt
YQOmJajTKyq8uZ5ROD6canrBKD2Ds+cAqBqFLjpsKZEP7nB2D8VLXstuMBS86a97
+micMBT8AWgK0BbFebqV1YCL3M1UjMk2JhVSW/nhnMUj5/W0YYDLobRYvrFhLxLW
0460xLo3Stz+Inge2yTaanMQ3nQqLBkbYm/O4BrCYTGyS7j/f+XFAv7Rn81MbzDu
WjyzIoSOrO7g0Mre5C7LQwOOWnzci69ws7JLSSUs0FtSykshm1VNK0c3OycwpSfK
SgKkRcO14Ro9ryPXc3KWn+L4BtZFWkPIv2eMjcBL1VgZhO+UA6bRfyW1DyLDadRH
p9JECeN3OVDxvHwm4t+nIz2NvGlHAhQtg7/wrH0jWk2mzmeRgFz8eE9QeM5CldnQ
GA30ddFYQDpNRFn2rZK36t2+5fgzqv/yqjOk8W+WsKTcMf7zA3QucHkKF4qVQJbZ
N2nsDzacitvYgdKimQkKbPRPqTJnvgCNb5mx9vvoSLHhV9c6WLYtn4mxVQbYazmm
WL6RTOH6PIBwnwekNi8GO6frk1xqmKnQrKmaBBzoAqrMkcLNuhgk3B8UIDkRASJP
AxI6t5QVDQiEv8M3cLfcrYjToRHr1IZ2F4riNHxLHwxaJwq46rL8JNV2P7frEtzl
pIPQLcE9855N8KiA3+u3ADjrU4iS1H7grD1QpjjDrskpqhZxuKZH+lkhDQ0L98KY
aC7ZIkkHQETX1CUF26S4z3cU47AYSf0ao6DDxMCRY6No/Jk6/nzaM3sHYx00dMPg
03OGMnSXlvEjDq0ZUEVB0/vmPRZAim1PmJf2LcAE/cM38OLIzTLpoUrBZMrsG6fb
a/CtxzeyRHgYFjcD07LeI0FOGs0lMzId+gYfXxwsHJR5vUCajXJkVOQut7TnNFwS
Jl12Nv9oMu0vEdA8dHfEx63bdfXnzzzYRL9tUkDSHss0yxX4QjBJXh7qUSlOYmsC
DBWvn08FDrg95/LFgAFkYlT+po1j2aMGDFcipaoKFyY7HO2J2BNpyBDvXtfwJVwa
B5sGcPsFmoALsODIsFmYGBTWajhvCkNrYxyjL5+lavRLtYqJHF33KhndVV5W4xAv
RwJCfak0KYJSq172kY2cgeKT+ZcEcQzUD56rfLAge+zocri/Tk+b0d8hFOHbAobe
fI0Y89gHZWAgCJBSdY7YNBk3wfyCWwqbDyBcLOJXnnaZeadUs1w4gMHZs/hSkMkX
Z+Qd/R1U0v8fACWz/p1pMFEzLuz4P+BOUmw+Dwx9CqQ3m+JiGAUszIRqTmKwDRzN
lLd8OLYoICJaD8xHgkyK5spd8xpkjMZHCyVcPLfqBW0YPS7tJoRL2td5LDOG1NZS
5ldvG2fC5qeWJ7FAk+kRw40PR64XW+rhXRY1EWdpIIvcP6RqHmv2KGAl9C0bjSCi
hP6XF7I+lmtovXrw6QmBG8VSn5bJGGH79HOzciIMOmQ6tD/TzDdYrdtwf1Dgq5NU
ZuJ8JwGUpGcXSrkFxSke4gdofafqEcj9I1n7KcexqvBw7cMs4PC1kXzpXJ5PP+yh
bEgSiV+b7a67N+O3+1mpMZqUMVoXBt2eIyl7qD3mqqsst0by8voZ5UwFDjksyo66
jWCrKWAoyzSF9lnpuKlqthY+mP2Z4/6HMzixILt8POjJEQGe5+DKX46DORJFeayZ
Xi0X5BPbfXJsh4Vy7DXMu0TgVHF4M5P47V0hysfjglPgEfpdx6zpYnTJgbjpbsOB
ImllOFj5RyIdF15OleC28J81VYqwbbDMDMZRbLt7z0Ka6xMO/UCF2gcwiFsLXTud
caBnN/KAw68GlPUR33jGApTnF/OZaFtUnCVU3BfbL8rlLBsrb7g9e0wR0VfNtLgb
Xcu0iI8Jg5RgXWkdLroD86HJnxP7XXBRLyd5b55JD/ybZUrx4oJdGcyxPIDGkZid
04uRVLUfYu4D7u+HKIzTkzNeDHtKnZxMd14o33KFzsx709NoKvi76DSlu1pl/u7w
3ENlvXUmwiZygH5n8QkOzNBHzwYjE1CIvRNXQhPZ5/3cXNd38Z80Pr9sM5x+fsXX
ss2ofarFYHKCFVXbcOpCAMQ23n94DHGGarl8cTD5mtz0HVvXg7A+Vok5EcvSm3sd
3eFe86eLiEZxYz6RwxTEGPkEuFC1/F2hB0dkiVfKCp/mFuMXyEIY1UzURkOAsZ05
fblvkCLlOG6OYXDjbh/uzop3LgAgNBmo9hAvvjkBy6UR1OQRVzXeFkLvP2+lyt1s
8vnvLWJoTg1++xq41oTVFUpQ2IiYhhJyoNom7m5v6SHZBYuhotafeoieazA+e3nu
NdnMeMQ5gpgbj0aUbjXR3m4y8P4D0U5FlS9E/LpiMq+GokyJZLffR00pviboj+ku
fWe77TBInM/0sl66noSONczZp/WZklQvO1fT8WUaycWjICOl1nzvfdR7o/5iXc9K
mL/chs6YXmQZK5XrslhUUGluuPeyQBqm8jduqm1VIVHTe8IkOPQc0+2jMeCHnCtD
PROvtCyPC7rQru1Cev7vhhr/KZwtUJTnlpUv+E6DHGtvWxHDTQVlNvIwK8cNEze0
z72zA20b8fddVejuJptLTd/7DLMJF1tZW2UY7VA3Uc3E1lVrFOFmX0k+U2kQjxUa
19miSEO6SVqJGMm5GEeI+glP/T+uRoHnFUwEUS3w8bo0k9tA/glNSBBu7jIh4IiU
biMSCdDDEklKK4zV4eRDeDZn7K8ppSv8wjJeJU4ut4/2yv3j7vZjfF5d0EfMU7x2
Qtj3IIPuGlkef7z5mzsRP3kQMrDyi52W3/S5vfIouCle9dg7LL1QW0xBzy9dCG2O
TGX/wpqP/K0m+Xv+o2z105dR3XQSPzTgDicC+DYI2g7lH1Ks9tQFhrd3WqYp2vqB
W7l441hxJ15ooAff58LVcv4QvIFgmOgCYD10oW5lmuRyMmPLBoZNoohWkNcQd8Qc
wMYMX+C8CYF7sOVhT+/j+U1FvxESomfpeZ23GTfI/3Iypu+CORJx8rH4S47qoyXR
LOvgr9iHZ+sDHkHDRHsVx2nBsolI+tun9/yRysq/3/IZ2gLkHT0JuIiCJKvPcGdV
PXgeai663UaUQj0dmb92cAzO3Quxtg3ulwPhSvCkSd9CPp/+gxEd/0BYIwb7Tx0F
br6+vpx0aej0AKbZciQnOoEZ0YfxKy/8oYCrFxy5vjZ+J7CYe/I00tAz3Xhk2FbQ
F8pnVTsRw0PjJZi1nQ2tX06cHxUXTw05qFclcKNyZvqeXB/27iKy7VT8LsQaVRvx
UYv3XQTBYl0H0jiOSAGq86HpxP/FMwB+TcZmGrlzTPr2hF1b4bBgiKOqq1ba2k1b
rh4JdCP1aow3Jqm4SCgVEdiN5xvkcz3o1RpVnCaLUNHlUasMj7nLX3P+h3euJ4P6
+h34bDWGoAshx4sqrYY3JCcQXtE+L/y6hvpg2loAmo8FxAqmzEisHCV4COMZWGOC
LpOW+9yqlToefSBTlxu84FxlDlMKezoK20EVie0AgyYApP2g0QyQwsBP1e1VjU1F
XH8iPird26jhBGT1vWXZOhNJjI8HcYPuyheaxSrNc0z3h49YDSdDUbMJ40v0+Z9/
73Jivv+fTGHJLInYbF4K2HqAO4zxVT+tXPXQKtIMZptnXYd5Si9FXlALTdtTLz3B
JykQDqv8lhGs/hNI8XwUZnldH9PuvITYVVYtAMqsCRXYUSN8MGROa4KdzjBJClEA
mJtuOW+tbOcidHMEBuRnR9FXrRa+cc0QxJ8gqlDmdlxhynYUViLHXPxUzrXILIIE
WbFMoCyHy2Sbnzl2GXuZgTiZi0eo1r2UK9AYBYQBZZM337ZRID5T0vgjs5Gl+a+7
U43X4FTUL+kPP2E8f94mwuff+lWsX84/gZKQTBonqzyVz3VyjoIJON0JhBDFppW/
Uw2gm7DwZ1KvorFMP+ROV7b2YFS3PT/hiv8yYpyqWquc4wtpKKPDD/tzlOQFR4FZ
JkrnZlomgqJABIPyZYbMd5tzH1+R6KNGk+fi6gL0XQ5bXqOVuL3KgXqvvTZWwVHj
LEb9IMb9JXDyex0An5VwY1uywQcdh+tSIpnjX+wLQNi0EkDyId9KMMezJj/rv5wV
MlA9Gb/7vyk9fNN6ur98yV8QCfksU0n8XyEFKL5ARYQYhXUMzRh+i98PW4YJkkrf
CZEta34otXdsK3/ju4WKIgB6FTh/umDPqdq9Gu8cePr+R+zDXdTBPnUidaqDgU83
xB6GeYXGgIjCuDyrEm2m7EIqDwpIhZGHGKeF+zjvcYCXqB2sCzsBe08rEQkFcxF0
aGGD10IQq6krLsCfyK2mYc/nhETIqzWvcg0xFFepAdLgvzEwl+1I5UQBBhUFOhQY
YONAUMUJnlirVXdBm1+x3sWB9rWSbcSZ5a47J2Phzev7gwo/bIMaVvm25+0X0i2t
2r0JXlE5xoylvmomxha4O6GE38kQgAH0DMqX3mqQ0oAR4W4Ndw4M1VmHZgaMT7lc
EuHyGlwJCim/pojauF7TMS0TnyTaSkihL6+5y2xZJteNvLuIE5UP9dHtA7qi4Sdk
/kxZlnF5a3QunDDAFCSQ3ZwzZbTJa+Lbz8G/oPINxYUnUtgBFidlkSNM+sHdJO8f
MwWm1c9vmI8CT7Wc4h4YOYjra4aMQ8tosFyYp7UGpkNFFtfKByivjHZ9dwmq/t9c
XfgdG9EgR14nan97NUqIU9I06Dkzu65KlhZxQIhQgVOfI1cSv8c4CgKztSMrIKOa
QguZk9S40vf8eaeBysI0O6Sy3q4ptZR5ER4qMdA5HIE4DwjyLMQZUNQlHuJyih5Z
8ZS4KY2rULnaFPg6Xl6CH99VwM1cgL/MT7bk65CsmYvGhgek0k7hd+3PtzWHir9a
Jr7JlStrywyr5z7hqSNjSS2ov9/4v2VNLB6QKojgSCHTmGpm19wkEIYAupZxJKGp
2DXwUGSHqVtkt28ufb4rHZwqMgycg20GTa2mrSnDlhPItue3wqYE/WgQtLfExpHR
KeNVNX5WJMWWtQoRO99MjJ3+r7Qkj4PffgbmG8KtJU5x6799cOyObGTCh3QmN0l0
A1Zt156Gog3zmdeDjzjVioawb0+EWDkj121qWizbBilxD+c+jBcu8UMpScsZupZO
TOkL/l/C5Rt5K1J5OGOw6aeMQutj8nOStFjs2b1UXueridygzC/Xio3PEMpJw637
nU04huyAj2RAj5FhaSWBHzKI6FImNKZZEl3TqX3QIrwANMxrJFdIOLl+D0ECY2LD
w3qKssPjozzBD5CMJUmv46WIc1FBXslm/epYyryEqRNQb49CgImlEZDzYVkVQejk
1pPPmERWkdMxSJ32qNjWpWSV/qlwYqK4NHqWRMflpmnhCxEUHU1nKdz30exvUgLH
zdYOAneOTs4hLILlwGiAqfldBvYt8yGJDpbtaiOMZsPQRbPRy1mSL7J5iRKxGPH+
M1QOxm4VkCnzK1LK7W4GBeNp2jeeTx9JGykYMWvTKtkltEDUMimC5Ly8HuiYBgjx
q09ZSpSBOrf1kEsdNv9Xxf350veyDv1w/r0coKL9s0G6VbAtSJ6j+rPo1SGiOZQl
5M8V4k0bu46Gq5O4FLiR+B//GDJRLPOQVcLLuYDZ19rTJn2Q2NA9KnExa+oxBuOb
RXh0asbZrmF7OSuvU2Cvl6DGWDE0l1/9yw0YQ7DP5Ulw2DoV7z5VxXbHPDxxxV0K
p7DqVUdByO/SAF+U66mqkfWwlbPJ9TPhY++J6y3xsO41nxzFlgygiYVWuSnZ+WW0
YbM948sl6YfpNEvfQQmn3+y5dC8pl46fFLkbuFQlexaUq72I7xhZSg7RxFy0uHen
uGx2ufuwouiNnLLDhk/eBJAw5X8838+GqBin76M1BeNe+u0rfVpbfvwX8FKKIdiI
A1qXaLoK1N/9ImCjRinjs0SyU48WUyjZffKy1XbvJ97GE5Xpja5gXvTa44pxqtqD
rBKTMPtdIEieH3JEtvbv+KGyCHuqyftWZtccW2TS/PccCUBUmkie2qhHUScp+crd
48KQzIwrcUg9D7GaXLWdKgKTUca68nmDmaSKJBRzUQLVWKXTl+FIidyNCD+nRKq4
1CdV/ut/5kOn00TP5DDSgyc8qh06W86AlUz3NGM3JJVCKE8TjhIjA+AtN/CASuHY
3gNSQTHNxET0cO92+Gh3dnfJYy3Xa95ma9muKCyp7e+9Ph42VFLKa0ivzd6Dq0SY
qcnsjSGtWQAIQhyT6186uwNwVwzD2lV31AkNSs0+jwBSWb79ZWQ9bd34ZMJigi8w
Qawo9NBnewVLthiMO5J9HQSdyVg8lDhgNoPzqQxIsFyf6RWgrTEJvTrlDjx78S/y
LaJhkubLYL0Cgn6cjt/jPrht4jPZmxHY32A4F4xpNIAA11oTOzD18HO5G9sekDJI
F8xh/3FP/M+dhqdDLzysmp6fphisCmGB5mhHCqUibXHVeDQddEEMDQEgWHH+mZxi
MFN5j/C9nbwfCiaVJd9AqQq/DKT8sJ/Fa0EZn1nWnswgrMzEoI8oB99yQOxpsz6O
Ry/u2vGY8+3LznU+GMRZNYeOWc5JN1luFN9mj4J5K01sdJvEcjs6/kC8MBBdxce9
54hM6okj9IrrP04NeCWB+hu3/4k5/Xr+k43a6WrQvCxPFCTSqXg10d3IT6oEIuRi
lWKyCpkYDFT6VNVZZawf/0Vv0E0ljPV9+EtQkNxwXFarE62tDzTMZvj4vr/WHtjm
BtNg0ieqc0/nkzpcYRw6b+3PmdUIqKQ+GjQF0DOGKiYm+naEB+uzXZUAuXCO1NWI
aSaOTtm9y2uYCHFofE7EAMY2EGKF/52VY6JjRb98ImwKV2fcHwqs9nCkJfyz+y7+
OSSXcDTUgdXoThOPHQcZVxlwzkz0PiHGGuaBIVPb77IfqB1DAxKdMiEzoSr/sQ3y
V5BpL5XMpl02TLbpqG2uz+NkHHRiPU48gihNRAV3CsimM+fmDITM2+s+JjjDBc33
NUz9/gQyNEj0466FgYjuC+J4JWTKsbhhDiSUMvgX0WWu/bRMT8tS8e67X5hDPVCS
Rm4dWhJBWeeVXsOLD7DHLxoTWNa8sxc/u+Oz0C3dg5q9ViX0qYRtZFRwsM0r2ceV
VFvNCvZTquxrSjnjf7Yj0aYjY6iGtcYQwplnWkiD/HOyumEmzs6YS+I3izGcLaoq
zypP6G3Qqewvst9KdEkilqSS9ZEA3ZJpNP0qHvkyMZ5nHLm+Oyp57eOJ73MRNgg0
uujDO2wNYQWNuFDn1Qakiof9y2AEqvw+g7YzlD9u+o0hUAspOpnLMzuO13Z0SFAR
`protect END_PROTECTED
