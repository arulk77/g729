`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFdN/qJOeYX8OHo4ueHv5Ccins6zUIW+LVmCM2Hl93vY
FqtM96D97WCVKeU4tsRtRp5CfVi708SdV5LmXwRy7NUOHdXYe1SJ1SbkQ3yj44wI
ilYXP7jDXmD24oQ6D/2PrFmOKvkn0Dh1ujvKSGp7k4Rv/KLYvD77ZVBm/Wye/6v3
uOmBkIfgBI5hW9rN9c+59z1NcZzYhKg+G/A2xuFqU7W7eaUuD3kgF5Z8Aa8StuxC
7GHsCGd2tEHZskC5cmZX6ThANWo6o8GKD6q1OmjDcKdWaCHrSHFYZ8m8yk2e9IsF
0i4JH5z1NZeF7oRkWtEEIFPft6t3/YEYVqOIBPov7K6s7XgTTAZ58Nspi3W9x01d
V7Xl1ZL6NFUUl21EOWj2kg==
`protect END_PROTECTED
