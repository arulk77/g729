`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
z4x32w4b7PcnK+DaPPqEgsfkRxDs6pTPn+FeWZviVeqmDFFXmJeK5kGnF5kuZZTd
TuZpLKrjfg+5FUDwGbN5kPEpnO8XPGeLXp1JBXm/ZALZei/aRED4g5hA0Ly0QO2w
7Uja4O091Kvjc1LFwp6v50M26OTXDMpGUDY9zLEfFR0=
`protect END_PROTECTED
