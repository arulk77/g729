`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKYwgEwRHxmd6epJ0Zi1pXaDW1lUtVmOrO5Dz9yAuSWl
KMKqEIPh43KGcUZYyJuViAyxHDgaTAl3NmQERNPQ4gHhf2CdHtz58Yr4UCdehUo7
tpBEZM2CAb39ODsmT38PBarLTYtK7y2wbxIoowWpc7AveHFO/DnJRZyWLDqN9oII
BY2GBlbT2Lc8dU9euPHjIaIxidF9bGuZ0DR7WYgRlFdr5kuA8nFWbAku/9lTcDYg
vQAx/VsC7+fkEavrFMvqXiIEuGRvrxIPnQlK3irBIC4egG2crT2QzneqXHEQ1iLM
J1xKJ9Ho6cPcSapJ0UXUSZJYFiJFHiXYEJJ4fMPq6OfhE8RKYHMa4tH3eqmBrm20
s2irDLjdTTk/fBzj7/KTwbB43YDLYe1QN5hY6abuKwaUJ4LIWl4ETfLccSXKLiQR
XMoBWTlFMlG25fYtZRZPsVuFJCaR1oGtHEeFAwyRQEh6Cgub2Fd9NvRTqwVDAlWi
fuut7CBoZpKWXfWhY7blFcFmszF4oPD+ZytB4NHSt+D63HbfPRAsByxJXjYwxHeI
zNpF605ovbLRGjRRsAztgz7h1QLRWY4BrpDdsxB/0A8=
`protect END_PROTECTED
