`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wzl4WPwHt829TMa2TQIxxADTl114fpD4twFuYfhQiJt
VUxtsST8V6Pubi4xCknGYkQ22qIzLz/gJqLTN+wVBGOKYIr3wID9vroGDjTRnVwi
pCqkMrrcMbGhrJLlpfp7y8wQ8BQKOwz5HqBj7hnPqk2MGbzfilyAf5J4w3XWer/V
pFRNBY2JIbvea6IoMXa9gq9ExHSK8ZzpannjetyMA2s=
`protect END_PROTECTED
