`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDYvzvxL+nHQhwLK77PbwSuCo4jmMM2raaZPe9QMCmyO
OpUBA+dVETrKOWucaMLdB2DyF8bj9KeIstfWcbXyKIHdUf/bs4hyZDw+sZvec6UE
WH5G6/Id7rmhbSzes087O9bqhrDQ06r3qkEc72fzJCaMOlCFM1t5Bl7UG0TFEJ1J
PorZxqojVZjXjMLgxCmU0bow0UDC1FcHxur50ZQj9K38W0s9LedQmMURW82V/cjK
IwKbgT88k2pTpeb3YnKAdB54A5hQSMo7DipKPJ85//HASFyB9sU1nHzPOY8KdQZZ
ftMFRiy+5NIUtsEHY2ZPkYs83tEnAl2DsezT93r6GyH9rwtcs1yvOTWyOwvUHuSt
MbmcGH8+/eljs72IAAaLExbDLBbQRLnVsaIvVZBr7tPNrK/NDmKSvgT8SCf1X0SF
yP/kkXOjFOVPIj3Ybxszw7vTcdLYHejFTVG9lFz8UuTX906MORMl1T//dvFCr3/7
If8pKIQOqTy1rdzrZAYYovugRqHCGVHOqePHBOTtsGzxMdKh+5pLB1CyR1SFX736
vm6Nj9pgtIKjTr+igSvBXuyVYkpxtp0TPyo8qOGu6kzBYrKobi4lKhfbK03Rij8X
TR9L5Y0m/FagSh8eF3ddIIDloUTdLZ1yp2sfKSLbfpbvfTCcIH2ONLWf/7GbGlrh
HjGUfPOYMtVz8AdLYUC1394hyhdDZAnEGqXYhfinVyZ1kdjAkrNzzZ6x984g68vN
fJ7ILyo7H0mRGL1j0CK9qE5BENJQGfJn+nFFvASy2iub59spayIQbDw1fvRseFBv
2ZZTMSrImNEn0YAOncu4fYmnguR3HnEP2k//gZcROn8=
`protect END_PROTECTED
