`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDTKjUKfjh+mCT8xf5Zf+mG16k7GAEG8UhEbNrJtmUEm
J2W9xHo4M18YDx/sNSsECXf6PlwK6Xkv0utAWBh+O12YawPx4zPkgOgIGcjau+ao
Nq+aSX+2ZwADDkkFRpplWtI5OLahcX08kow4GyWqTEKxMUmnTvcYQP3xuMYIO8Qp
7ws84OTax/UEWXRVq4YgVA==
`protect END_PROTECTED
