`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+OK4H3goSz/TEm9miAbMHaxOHF1BQHqe+hlg9DMbecp
B81aSq/QKbWH89qZm+2P8HaOMS1QMpJMS6tXPFzAfUplJB/68oreeGhmQ3rDaPw3
kFUu8IXFP/tLOWGy/8INBQp9bROTJn/XwEyGmzVnKMhz9GaHm58W2Zss1cVdEygC
LhoYgCLnmCHHiTP0LbC8dV/m/vObTWfqXB9Sq2zgQLXGbD0PYkd6kSxFIRsZkV7l
8HrkhzDhY8JmWzAHLcZBWFl2a//CXhSmdymzNPlayd9Y3mDd31/pZqMXXNa504rI
1Y6Z3GD/Ie7Z1sfQZGftvQ==
`protect END_PROTECTED
