`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42IVmOkTdPjraSPolFPe/kcveLjWssoCkwgDMwJ/HnB5
WfkgtuD1Aftfk+6zMBD1Gg8AKgiYtKUC7FaO1TGB5oaL8tctkOKZmf/sZ6AdVgGG
7nzHR6jXFMqdMPjqBo6Zd4mgQG1C/AzdVw8kT0xTxiFdj+JuF1IYMDvUwgE7NebY
DEeG97fHyZj9yOOVruQu12jdmE8vjDQV4fMlyh8+vcZ4fvd9jftrApArzZ/WowUP
XWgNNuqfbnGVTfsqfS1/JkWQbLJ6vXUjfClzFIenpogkajeVN/YZyJ/17Jh0pQbc
PkzMpvTI7mehA4kPbj9pVw==
`protect END_PROTECTED
