`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBxi/oJ24Jx1S9CkVPiRUmwD3JWuB4QnXt8JYXP6/CxJ
j6phI8XHkgE13lSugFGmNEthoKBQi7eTaWjbTQ/BWN4swNxYrwf4KpBPJ52tW2Tx
JKJgCnj6ut1ACrwbfe3+QihcYPHRwfVvKhpwZos7xtrOM3PHc2ydVjuKFT3FvCAu
UsYHg1wydgpECmxu27ZRKd8Gq6jR1CmJ/lHoV3a5qmr6Dw40UvzuV3R77xwq/A4A
KeepuFQB6wmtXqRfFgtbW1ROu+PSaOCnc0mO041s4pbM60ItmauF48soonugfgAI
fFJb+fk4a3EYyJF2j09VpXMgaHmFJ/d5SMSgUAO1CKoGvvyu/36MqU03yyCL9wID
4JujDkSEWfXWGW4PdusXEsDA+hcsxl/JIiaTetvHs4qQdJW5IJ+qr1dpOUlduo00
5w5a9E+MoD/744kNPUsD/g==
`protect END_PROTECTED
