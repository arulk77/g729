`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFE2O2VqNHL9Sa7bcNcpoHX7AcyZ4ANXOqFvr0V6EW+K
aHO78Ux3UVT3Gbd3teJ79Zvp4+J3CynWnSbxu1P1XF3eR8FRb1ATl1BUoFzAj07b
yC6PGgzgtcvnGGIfntubdmcet1eFA7qyGmlWgJSwiu3MRcABYxmjZ9NMRXhl/ibW
q+SDyG00BUWJMuvd1q007U0Yr+YRHB96CLV6alfSo0nKHFqx0JwBkrezM/RZK1gr
FIfDV+JrbCkbNoHskc13espO6kvp761dfP1QM5GdR0iUYD1OcS4smCAgzkFJRQyU
`protect END_PROTECTED
