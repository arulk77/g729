`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGzQS2B8wBMt+E1sdXFyyByMhV5+0T/rnegSC1hQ/z1k
VQj53PZTpofJVtV2rBhC2UiFAd/6QVqzcAUzkmf2m+EKBY5sq6dLFFgrmW7KyjUj
0PwFj0Av0QLYyZcqpGdZ4dkOyQM1sAuvaFdQlKGGm1/e61uCtxpU72lcrjlUwlRu
hweqz3oB3Aaam8TDzAUSv/nicgtY3QD5okTqgxQ0Br3FBmlbtqKewUmbskJNqQJJ
`protect END_PROTECTED
