`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG5A/eiWh3zAUloR1HZD3RPHPIEWLsXNXnldX/MmB5OF
CHNDok3CvvEln6mL4tBnEUbmwts/Ky69H2MXbXT9cdHyb4SVR169YTWl+XO6vtbA
UOKekYYkBNxQ6ns9k8Oe29xRNpxeWy4L6BZwJ+IVn8VZV2EPrbHcKVUg6RywP1qf
OEkqKdBGWWdXungeURcixrBXgNc/5NW1kQdKDXJRYD+B9eC6THkzy9ZDhpge0AOg
FRPJ4CiflTBnojE4lGJzoKkJU9SAgWm0nSsk4gIo/K5XCE1gxgZgUEqM0SoLGfnP
Clo5VNv/DlW1u9aJhDGeqS8bjFBm+Jwku0ajp4irHY2C3LiQDy5w6SIgdf/bkfif
5c1Kb6FULxDCv2T/pFtf7Rj6N8/W9OMtdPOUtUOSsOI=
`protect END_PROTECTED
