`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aTuI7xfZFAVemXRoc4iPSnCc4eZk/7Kmjl75j99LndoN
2tZ8Cl8YCeormcpgIYdN2gykg0SIty0LzMhDhLSfxGx35RUcuFAgDe4kcrsrSEJV
Ss2GbovpuMkgVPm0lQbfVeTKHLH+GjXgg4POkW0bkUNwT2yj/58fLCLggUquwBfJ
tG+BPMYVxrvMgtEnsjjj9e4PY/CGF2gA3zEAZlxqGZu83Q05kv+bBWtkeoofp0OH
gO0/jQO9qf9GlFM9xubr8bDWRZytxFITQKp+YNe8wPYlp9SA8Sd7FDKZTy3FJ/Cb
Ku0/+NxIU2yUln7oJdf7/tgcJvGTlPxDS98AHzNSS/OSPOEeD4fZPYpI3fUKkVdF
SqbRareKVh8O/xx8bvMM+w==
`protect END_PROTECTED
