`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCTNC6oxkdw90s6asdS/Zghvp8OYinjsFc9eLthy9p8G
xncjfWpT7eIlkdpacT2J5ZXEwiZ0EQ0XVQbXjftnxvOExLJ2VaAw9nruPkG6BzCA
EYtl8CMgqR/1jruo/0cpkBjE9wmIeInQFJqq5FQq7ZPJAO+sj7O2bfx5HUp15wmQ
8ZcZ6hjOCRmbzG89CHLMsNj6fGo13vCh59HQ6wgXet0mXaPXNYF99xCac+bkMVLY
5JCFdfj3g96cZYsAchLTi/YApGozqh6ryJi6Z8Y8Jn8dEhS1bGaV777MMMfdClIN
7qcu4u/TQ28zT+jSd14JBTUzKgiDbjFWY6Vs0N+Y0yFgDR6coo+OauOk1e9epZVD
ijSw49AJYZrPgWu4VZdWFlM6KtC1xFB4CPo538Fii/jO8y3a0mIgSHf2+cXSPt4n
B2BQ6VgFXAm2ubGjMklOoCDHN7svbQAQNsj2cM/whru1Wl29H402QRvU8GuhiYd/
RQy8IP0kf9Vig8qB/9rJp1GOP5y04kw5wdlfF5HC6oBje3WgCzyhW2Jg3AFxzyF5
`protect END_PROTECTED
