`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOqObh3ZdnHGBxJLMWxSLPZhtJw/JkYuq3iQVBD7+ng3
t+voOBjz+Y9CcdA6ViathXMmLI8fqOYK+yJ4eP9MF3fTP1YMbqg7l4WGQLYUpBm7
LxhhwuzkMkgTSFfjPRyuHida3njO6C8z1oR/TTg5iF3tmEmHxF7X3sXTQjwvhe6F
`protect END_PROTECTED
