`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAfnvlzl0e2OdenB7lQ6EYb5LZKDuRfVq+OWA2WPAqt8
rfpo5U1fbz+irOzEipVvx3yGCuk1jWW85vEyBWUAKiNyVvkDuD15pyZLT/Rak8Eg
+9W1xj6mlgzjObPkKanPizGPHvqHCbOboxLZcwWfv+BMUofNzEsbaGBLDH3QQALk
nrb+BsqRJro3rypz/DcBmwKCxom9rOW660DwxqpS5KT88QNpJfnvas4zE/2yfTp/
`protect END_PROTECTED
