`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB+pcC6DEb2hCYVQ49J+OdC7J0Eg8JyQ6pa57qMN91hX
lP3ftrC5HAjXmVWxAZiJFjSVzCgV69pbWdEMu/puFHeh1WPyTjj4HCq2lX+o3VGt
xSbTPjpJcdSHnSyfaRSgqEDi2hsSwPI5EBFBCUt0qxg8MN06fC5o616oJY420Ju+
P6CgEZtVq5GKIHzr9uP4ym9qQ4XUz0xy3PTa633xEK5ZcciGCkPSCWogk9tXfXra
jiJDpS0i+61h5TNYgP8mm36pK5yeNOxhw6XDwtrVOxvYwwsm3Q9tKmX5LGLQiNYm
iS+GK50z7jYbo3FbGDWEWsG5zlMfX1t7mSvNfvebJEEGZUIGYscTBA9qKmkOW0OP
gUL+UtzrlK82/cmDGzgwJg==
`protect END_PROTECTED
