`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFqUllcqJ7Pmfk0zCriOgaWCZyL/MBISvH8Gt+9/b2wc
yGOog8R5EL6V46F7sXBDRGpXIGAzw1Kb1tQJ0Pa0mYfvAvUANO2mT8wtyIDPYZQM
dI8I2GsramrWLHwS8ns9PhwatCOeUwoKYMBW457GftMQKi4t+0D6NP7rZyPKBwRB
/EcDNBDS6rPZfLBV3on2VfbDXn4msEJeccztocK7ueLavzCNvodwooJ9jlcr2pdq
qSRvNeKFjYnrBQD4GYkL9srtUbxcxSJEUoij4hhZ1luXrNe5o+7PFZm6DumF43G1
g4kmQWoFe3mxAwjGFk1hIr48uUR6xz3wC56WjOyWyJ8xPiuBm+tcwt8JcAxmXz1/
v9eROgeA8frDQihSV9YxEk9l6f7+hiNaNfybY6rxSckqGwX05k9FfBCvFbp1Kp/f
CErYi62wgUIZVwlDy1Iy4hnGr00sC3q1KM7WyZlyjF//psGwa61zk/3nQJXZTROL
tFAROT44uBCzVsCPVWdto6vCVns3E5M6Lqrqqz6aSLibreDJy17tCivVNmKQ/2Pd
`protect END_PROTECTED
