`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveELtKFo0pBZq8379ADP7buA5edKWqvd73tRgnGBAw4p7
dXkxBWzVHgTMhxSx4BGhk6xtOnMqyLRonud5R9TuM1MEJx5ko7cPD3fFCb64G8v9
coY0QkhdXaAUTKFnh9tnVcPl2i5Yr8vfhGRLCq5WupBHzgBS2Jc2lou2iaLfqefU
aiMZ89tuH9wUvKYrt1JQZR8xfklKzlbOcTlbsKGLzuOUO6icT2jbU/TGelMAjX/R
F9Lx0Xbt4bAulvgFMC4fs/jmH0zLuJFKNIR/m5/uWKwR+1vGKMaKo7MBs9BGsUr9
N5eb+NaYtvuj+3Y+2PxgEEga+hC38BR7QMPhht6wfBwiORY6VzutbB7d0K07MTV6
Z94ZTxRuke6YTzfc2GUWy4/Ds0euhsH3BuP96UO2K+jYh6aPKLneOFA2GieoKvAf
`protect END_PROTECTED
