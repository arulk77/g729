`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCOPEkcCzibXfdPA5F94KzRrYiirva9JHKBWTYj12ZZx
EVyI6zJw1YGWCtYvAjrKZ0cDjJpy8JQ60fxWZ1mLJIjF7dRLcrE8DRFHgy9nZFSe
bnQy2LMhACtNAv+yJPVJM3UAp4CzXbxYTDntc66Zg0M7NglOCy0PzbaNbyVo8HoJ
fKKT9gYZnVXkpooQR4267IC3hdbhAtwlQhZmllsT6N/+oca7CWs5kJMv2mNCTk33
+YdKxDBzJCHmSiypbpgK4CdVqxZTYuAz7hlziNNIid8ogsmwpVIOkSDqTWQVcaXq
nObCs5n5s3mQAGDlcUiSHU+nH7qzfw+uZJIIuKH/yml2FoLWlFdtrTZsxnFQOCFS
fV4t6s/GG7aML6GifD1CZ/bVLCz3wbflXFUcJHdlNErwhNKMDCEgWJZOpZ/rQ6QF
wIegpie6T1PQWvGGhTeueHO1wIMX6p7JINXsIfHbfm3iGXHx6PPJ2YYylSCMI1Vx
`protect END_PROTECTED
