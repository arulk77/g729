`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
vs+MpH0RaJikKxVYQOIYt2HZvnH88NSH3chq9MQqAF5jwwgao/TwL9nyI8Y0Y6YX
VDEf05StzogM4KdLU18fXdHBOfGSf8oYKjtk6HpP27mRtVfyph/LFLErn8pj2Tfd
E9q+2WcDPLqCV3qnoTq0xbzhptl8uK8Vfl8SI+HPuW/brClEvhjoKxrMXpjzwUoG
EwvLSncgq2rbCChAYUD4SN85pdmxu7f1UtY42mO+FNzxIUgzpkqi8GKfRSJhz4vh
zYVdkoVpP0qFNOno3knJhGm6DhPR9i8plTZwK9ZJKSFwM+zKpXtGjdfJi3gwuVnw
ujf4VamdruCXVwij3sZuXg9dZlb8zEuZBxbaiqGPppE=
`protect END_PROTECTED
