`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePRwEpJr5OaDX9l6eY0bH3TRN5t/L6eBssddX4jNV+Qb
bu8FxdD/hihY70cCPKTTvRe8FQFnEYgQvmEsKbxz1S5KL2ZYYJBypH30QpztUKEK
SoYIlTn+OVpZgwWcBOPgxj486iuYrvp4v2EdEIhUSWBs/YpMW+YvO5pltPdeHUgk
swQVYr6b4RbONnQ9lBVrEb55CaeRu4xqwdsR4d7+1eLUeI3kTUJ5lSjzeKrwdlDk
efMO1GTnXNoLC582Y5cr9I90yilUXO+XMedkdtGU8GohQIaUxIl8fGoR3zK6sbp8
ATYE+mb/q4iyNQZ6cttF+9spopmv5yWfszfTPHfZ21iwvloH1d62D0zEMwX9TYEa
x2HgLHPQy2A9/8GpvDgpZQiA/+p8lguyezlUygqnlRUoA1yoPC/gILiAYAV1DARG
2MkbMQZqUfKKMqhsF0fDDgrGanXvmvhN6lwXs5UXBzGnfrIByATaopRrmhvXcclt
jYeRcPvECIodg3LRW2D98gevAoJUWWpYRr4PREEh3RP1EGWmYpmC7wA+6QDvgpx2
46kdbAb6grKHb0JLO4d9uc/b1w/ZEgcufnliBcaW/vMWO7ARiqwPXnGouL8kBIuO
KDGELh/w+wSSo+OpAL+TVxq8fnrZmxoCrGiemg0cmfun+n/4n5jHJKtTWuKTAQZy
`protect END_PROTECTED
