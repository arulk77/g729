`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73CxxDCmzkJJY2/KXqDLFf72rUnxLxpSS2LXcur03+mcES
VzuajXHvEJCeAuyr57MzG+qJKhPH0UXStrkoLnzi9LwUO8FF2PYiw8ZzCUSi4PK3
onUpKjionvk49TArPn5W+Z8AuCKfJ2j4XVcbTwoKWBwGuT9helmqdFNOuIsj+POw
KE7iAXDrbiwcV34QfOSnPEYFrbxoZzM2lhFy1H7G1WJP0ZrW3qUf98xtLic9Nwpu
XBzefxUV1QP+RCjaQbloQ6ncZIq0pyPGoyRdkt8DFtPu7r4kmdpxiqnUQTMQvDmA
1P2C8c+CLdYZ4ZKygzXWZJ5x5tJ4oTmoz+sjdcnABwSq7g9UbqRaHszeV6hMUC/R
Czq3YlWzGK61xYVMOOeq82KvQI0hxBxlzdPcvsjpoGLAR2o69c9OA56CSbhM8Dxb
4ndysIZhGizDkQJOGrFaRNPVoeNQS/+MOJfc0kvKNYS7u8q2Pp9WJGDI0Z+fbARe
h4qyKiEiN1cs1FRRpYcQLaeGyqXFsKwNx26i4AF7ZLWrZ9YfHzRJhVFs1tiefgDi
u4Rv5HxeN2V7oKmsXpS9JwKvb1RHIlSubnKz/j1epjk6uPeEBFwUnqC0C8jVxEUj
sWYeahIh5JEFMEwapAUdJhz3EX7G9qpn+WacdRwGfSOYkvn/lQZ1jwkw94lZlEaP
OzTSxnDeGwIUXlbF+o7R69Whz5Wgk7MUBy6UP2CsrIw=
`protect END_PROTECTED
