`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
D2fAHLLwAfYKa16/FBOU7c1ZcefuYhxSuV4nKW/Fa/HO6reZviqRPePv1BR3iwvP
c71WlXJNIbkzMIgTMPP+m8U2vqhr+aL/f8x5+WO925Z4w3P+SJWkv1pgwNEqym4w
JFFMNnGbXmdSsnsiHA9WNZcoDyHqeS67We25SBDq2hAJOhL95lT2RHC/9pQZE66J
gqac1YwlXDWe9I27yztZDQ82m4Oh20ORcpN3PzJKTaHEjBfMFmTvQlGyTVrmv4t8
Cor90nApXxgsiDn5ETFlgHgvj5kRavZjk+09K1O14jZ7FBH6oDdCNyrdEeskh8e9
RdfSJr2KM3NQ0fc0vD1TpOTUBQiIzcQ1tdszn2doHAbk4d8gpxVpOLHAHngZn2GD
afSSlmRUlNItg5KdzkfrAKmA7pVRzG7AlJo1Z705lKNpX35aCZfI1qDRL84Dl5dm
/hPZFSsEVzpgYbnuGDDpoA==
`protect END_PROTECTED
