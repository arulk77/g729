`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+Sa4HsrZu6z0R6wUNrrTsGZZPIkcvcxh2URsdUA+/2L
buOiu80o5SgGT8TWdc0JK0yi12ky0HFoUKInpEfU+Dmq3+/qLk8Ltcw/Xy1YadCs
2Sq4Q/oyPgm9r1hsZiJa3JtxTO/SqJnJ2MI4Q/B+rPWfLwOI+KF9Jd/9vBj8zswp
+gUeQCsxt5InDePPsKzGu27wff6+FpYNJHlRF5USr0s9rVvIIhM6FWRrf1DeSJhn
91PYRN0e8SXN3IMKbbhgRM23zWIxu7gpmNP6ZuFj4D0J9iwqagSGd7B2x/9T7eWA
8j+ADeKXvt27Z6tegUjYXH9oNKpnLTHQxEcNc70PtSFeSGHYV4n78eNZePxsvXqM
WSDfpz4JGviaFLkSVxtLlQ==
`protect END_PROTECTED
