`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHc3SFv9Is8fsr91FtF5XfO16VzbE8jrLoovvA+9Xja8
PXjYOvSqC5ePFFVBgFSd059llnGu8qeU8a98Rze0YWsU8H/gvekFqAJm7CImsHtj
HuwntTtfvPW6m57+VoIE3K/MNyXkbJ5YEDv6RUQk/r40ZT3KAuRH/AV4rQbCaZ16
b5tQKK4kH71v/14mP69Pwz8saEV13ft1GtnVFHOAy2dEXJHinX2ozlMHRgGyxUhA
PvPf+ngJSdd42m43f0oZWyIW+/0Qk6k+hAyh8EToKbZamFyyTG8XDLI2ON4n32kR
qXApoMQIr8HnZybbEDfqZw==
`protect END_PROTECTED
