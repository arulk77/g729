`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/vVZUZFiDSkK+0Zd4taGRVYQG5+vJCyWLUbYc99czQn
tFGdEvqzW0gimsCtfgk2ZLF6QVsJn5alzR0Ku3FwsrTmCPRNfNNI+3MP3KTOo6fh
avVPVJUrdhThg6EfwFxlIBmxlSXFAE6wx2cDvBkPW8deL6RxzO75TIzk6I1Ts7/d
S6ESoS8rXno1lZ05aoWHM4uJ/WpwDwFOOw9tWgJpiHDWjMmJTSJLgM/soxCp4oCn
digPiqfvDo7XcnSHoWdecwXTjqeYWlThAJU1h3zqWLjl32KoTpPyvBeJXj4wuV/t
UgC67cR69fWcqnJiObO8yKP8aQDPnEabqkiHeyPe1uqSyBVNEtJ7B0aLbtP/dwto
VMSBwdeo1uHXAbzHEvYCXQ==
`protect END_PROTECTED
