`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
J5r+pj642aQGWEqoaMf3I6I7Ui7JZB8w4tTL7Qh2bppyCIVFgEFuVg5A8UNavUGO
lUJ6Ph8craMPj3g44YTbQm1fhZT/Dt88SXsUBS3bP/GmX4IRknJCXJd35fOWUx/2
u3WJ75NQGiaOdWz/AKGYAxrBxOJaX5qNPqSgYEDwaknbISDAeSAIaBn/9w0E+8zx
gF8WvftlOZ+Tnt9CtbPu7h0jVzTHoJ+a5Wu3pZeR9SqrDY+T/EXX6XmddhTAEyM7
aAwqC1VGt9R8VZ2BiIpc6AJBO4a7FjD+EXRzPHT4TLZwdkaB+OOKw/E0LGWhsbrM
toNTruFhjbbpYgQioliXaA1XoGwBMGci0f7REdBW+vQX9e+q0vIjO8EA32ThwHmG
rIWcxmI8ZFPHrd0ZAyZ974nGbtKD6FBI/Tkt79vFO+IK7YzJ7CtSrsiY9Gn9Ou2o
ul5v15pFoCMV0Z54mOfWUyAQgL9e96b1G+cF4C7NRVh+mp20SW7gtEDZ8FPCr+xi
KyPDr0S6Aif7hU4noxj3nXxPkOk6gITdDR2wwH3kNnfUBVwF1vxgys4gTITbTv3M
nqbcb7ZZFAScjeULSVfW1hvZ+/DxPmPCBuvmCZ/e018YijqHi/AT/3rmU+zjZfGd
gOTPwBp6wZW0EPjN7wdBQw==
`protect END_PROTECTED
