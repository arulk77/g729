`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveH/Wj27nVN2+yRmOu1XjXLk3E2YkgGGDjbpNOsRz9Brc
dCB+MWiEmXOtWgcuuJb1x94KHkjYu/uHz0OtoaMgWtETEJKUMuEtYad7SXataf39
KZflSQ736IjEoT0K05OQSJadrKZHPKxj/1uvu056WDkGYgg9nmWfiOTy2vFEAWn+
J1tAOjUJaIyRJzQU6A6xDwojzd7vp0hjYSG3YWrTuOaCL79hKCrMZ4QzoQyDoj0J
bFxzjXUNyjQ2z7/KswT4iFBCZDybI34KhJqdQXZ8b7u/7C+mcS17evYgE1vYXpl0
tnYtRPQXYkd4UlzpWMSNlFKUkmNPCl7a/+CCUdZcSuRWH/ejjUYhRmHZq3kCbOmv
vWH0HHi3xtuhBTSHUTsb2Q==
`protect END_PROTECTED
