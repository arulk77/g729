`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOh3MKQ9xolbZUl/ywq1aw3Kl9N/X+y0EGoX709ohidI
YF0Nq0by77E4HzPoZqIY7KIHpxRZA0uIpkmhQRzRM15gH8rp8LN/t4SB2THdbXzO
dmiKmqoNfphR4ARCJcAotaXXGAjs+S1zahxUdBA0Sb++qGAJ7GUfnVzVIABGFNNx
`protect END_PROTECTED
