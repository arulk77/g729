`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
lPT04+PXCcdoNKXAu754/stpQIg/GD5v9/HumdzQeMT91YkeTeCXTZnuH+Ty/vZ/
+220bHbDupa8nS6ytEiETIrQA99L+D8uuhgIz+VUgne1nKYqCS9HuGZwUaXAe2Iy
iIWxS6QCKdkELfFKcI6Jbo5ZAZgpUf+PvPdreSwYZMJ5760dhPZi6EVwPK+Ktgoy
01kp1UCmi8VhDpMLv4O6eLrURISreVkZ/p3HuXIyhea8Hhsj40p81ooaV3PZfSQG
YnHOMVwBv5YG7aIlZSCGnea6yaTkjh5XBVHhS4awjK5Q3mOON+g9CXbwyi/Dryvu
+b3P+Y3080zjU+7wJD7K5yQne2HhMeMVsHvuROBIWxEwXswiPnXdb4VRjmKy+O9b
PYC00SA8IWD6B7EOfH8pIaiVTDXUelnxtKq9pPzD8F0=
`protect END_PROTECTED
