`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4w5dy3m+pO2WHGny3sUyFIPb2qmKvobzbDHjJsw/3/Sn
8HFtJPmttO3Hcbp/1NH0wMhDROqZJJ4fxlLNT5Wc7DLP8va0Cv2WsNJdiZAEvCmM
n73huPYg5R1+NSAB3JaefhN90Ag+fwpFXIlMOO8zs/g=
`protect END_PROTECTED
