`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu498q8ms8VmZz/tZxs3buse/G2f7ksXLGGy0UId5v7vIu
eNKxiouzLYRZYiI6GxQKaBCVJJNrwtVlp42kraT/r70VZGXIi+moxDJLZ1+JgC5E
6PGG44yNc6kW5rYrq55taKvuDRv3Dz5Yji12iclCTBcAKhtoF1oCU7Ys+UxO9hl0
d980uDpq4ZjhbpJWPPmTBubchZ6y0VDSyDzNq2Zw/OEfWP0/8jbidEnReE5IUDJg
BkCnKOeuFec/EvuusAZvSnIzKFSpa/xCQFs3U2SgZhD7uz5C36KeXiDWhuRvY/ZV
lo5i5MwMn/nsZKQTtABrkQ==
`protect END_PROTECTED
