`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
UqI4p19hkPSUNl2hbQffZoDDAng9ANzOoMAgNiWEC1BlFJgi3/RMp7QTCkgRlh3P
ywIjb1I0UH8l3checa1DQ9sNYwF5ngXomRmeBzHTsQQW7AtTbqEIE+Twd9wZMiuA
sWa9hNsTMr74aPqskAKSLpqA6sx8jIXZ8s5jMSxe+agfeks3t+Zd2tub/6nxprc3
QQEHqauJDWKbcoSMGwPGWrH8pv5tS5mAbeRz7Q2D5hrACW/uskYh36epT0nhlh8O
cpgW+EqNEwuC/Sz+e26IeiOr605X7sPY4NS+m8hFo1Y=
`protect END_PROTECTED
