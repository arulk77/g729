`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG/y3mGOXwY/swp2SWXqw1PcCzKY2Gf07fm0r382gP3m
bAulBhu3uBEzw+3TYmEvWerYN5LGwavcyvH+C+Tfnvfw6y6x8ogivf5gqBgBciTq
2rQT9HZtUNHJ40ZY6B/tMkwX3OPvncHqVfb+4xDjOnWR/oz4hlFLvO9Pl/o9Yj2e
+UFp734Bs3CJOARKTpaqCKt7K1jA33WEaWOyGxnXZrSMgp+IXAvn+RTHQVtqPYFQ
0Z5yqN0QdvQqlvC/mBo1diAwZVY+3mrPKk4AUYZGevwbHmAstRVSaJMDlVh2Fhlf
QdlkZTwPXmGJ6gvGJqn3gpXxQfJlZAAoNmjDl9uVWh/gMimI2CBQxUD4ANmqvNw9
i0my2ZAmHK8E2W4KAjMTAg==
`protect END_PROTECTED
