`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNkMmj4EMFBW6hbgzk8a+2bPQ6UE6oBaztmZfrzwwmM8
NpcFyzgLlwA+yhZ2ODT4QJYI8LKi830vMnKr/s9mqxBgLlaPPvlGCNCl2Y7H1k/y
FJR7cBibdDzXTzB8JN4mhyLqidAaItvsP2bMQRMkwdaqKDuT/XGpBGVl4Nzxyxjq
ul4ezfUlI+TTrQOtqkZuqZJnVCgCCgf+XiDNCo5o6lLYXle/PQYgrTyB3li2UP5i
jw0rA1rvocbQPSzNDwyGgcYVT6SsVjQhEBzOvV9mq6ZWnc4L4TeeP2xzd00pPFrt
GK3d/hM8nrHv5ozQceYqCj5PY1PJx09k4xfDdQwnfrWzxgIh6nIL7qybV5XDPavh
pKUtmtPnMWmTal0qSXogMGlcZpwRneAE5iInXrg/PzRGkpLU0dud17vBlRvEWm9H
ndQ7iPVfmg+LIDF0XOv5ormUGX0H7GB9n0/sV29e+0pSlMMkSFQzk/yv17EAjuzb
HTJK1Q/d0cD4z5gumOxb6fZv3A4b4+UW2shX9MYwXge7ZfoYcPTAb7CwhNMiOqQM
4CJnqAAt33askVnjLSddpxQdqe0EQ4S1iNxIxfz46zP5wZDn2josZxBHMGnggegz
`protect END_PROTECTED
