`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN/dhgTFFmq3hiNKNbz8h8DRzeBT7ANJiKfnaFZZiQIK0
SFOdunRlvC9Fzlpc35BZzurnkI5Dz6vnSST/JVg7nV+JIM14xviGmX6zPAwrzOFZ
MfucAkPz9dhbbS+DySLdN/QfpiSyajBKblo8kZ/PUPDXaGdOfcZr78KWuZeOM0YA
UmdOFbI2iMTnt6t5eX/Vb4P/7tStsAlUoKn78DQs5IfUpobTOcA6lz0YMpQZuHGf
zLIrKw/UjMB0QTLBXjoxNsHQ3dOGayai5prrCudZawfXdieTV40hFEueqJ58WiW3
Y2oyXnYz7D4cskI8hOY/hbDweVz9O3BXHsRmp5/FHhPOZIBVC3f9i8lbEH7EYNTT
gAXQTXP22COZdUg42hbo1Fbgv4hsNx0Gln8X0oADqvmMkQTlXjVa0mDc3bGzUHKg
OtPNb5YzOFF7SdOeXnB+VtA7EEqfgYJs688FWe+EOADW22vBsrRxGpQ/Z2VnU7By
2lHuGMBI9/kzrCWilHNuDw==
`protect END_PROTECTED
