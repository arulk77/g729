`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePWtPP9Vio1hIGFHEIqP05QO9BGSV560dDZ3MgQp1Lv8
Zuz9QWjIL1woTZQJZ96sMaNdQzPpoSva+Z91U3eNYlte7qd8m6tIfN/DYMjZ/wSv
5J+Rx6bv8CKniQFMZFHslajzmJrWotSKLOaTbY5ubue8rYUiS3CYDxLwMC7Ld8nQ
Uo1eATAnzA+TKDum7fkujKaSb+NuK72B4mmjsgds0SJB/Sq4Y2bVMXC+FyvZhl47
PgGu1knCMKvy680S4PALgSmM9tfS/zQwbDSfTuUmPOEkNZiumfXg8Tp20i3LgBYi
bCbYidzVEW79CCtN3k/CJaqUf3uQtq1UW3v2KbNEBwBfWP4J07pGEXP0FoAcr8lE
aXPp2RDxRxbDL03IzrGeLQnnnKoOEtZS8lp7ffZLNHzBNB13tYYicpJhnXLygWqZ
IqB7N/bCzFm5Ul98r5vVlaPHVRg69cre7xgoOe1J+F39WCDg9NucTx9oVEtMSw5W
TrvZjgDN5V9T7ezENEMJaVHnCobjYf8U+OJZm6OCkYMelqtTjj8bcvaUURz5MeGf
A2F671TvIL1e8i1ZCbgp3m31RG5LSWN4oVl311kUx1In9JrhKmY+134Fq24Aa2vS
MC62kcKEWnp/ee5iTg/FMDHYFxRSmhNlDSUo5ne6v4jRW8J1ENr2ijnXXP/f75Dn
9gUQ1G/qudtQgZDoc+wzRrPybS0ZJeeInmx/IiqtEMqqsYck5mOjONyYkA4lfCpr
kpWbGtdzMyiMhwHtLa64vZMOH4Ykm9DSusgrhU7vkwi/2R8dHBnn+QzYgfKD6rIX
93kpTsQG3KQPgJ46dFitnKec6B5CsW3WDo+ydKBIdEo=
`protect END_PROTECTED
