`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAunoRqLAdOQ4kwDyl1SyY7YRkt9Dd0uHccG5fWk9R69
OAyeTtJ7V1O5kWI3vQEQoxjmro1911EywmYE6l67u04Tx30UNY4rFD9/xjU2JXZc
gJvJr72hW6OQCe9pTsNBwIyFk+NPuqEcPyghxxf+DEbO1LWwy/F0V2pbmE6Ryxdx
rCJLDlU2X6DcVR9e7KZZnyvVlZO66d11XTYCmElIlFIaK+nrJ0OQyjQ0yyr7+gHR
SYWSxO11zFp6eD0mHtfeWQ==
`protect END_PROTECTED
