`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8STM+hSPon29iqe81idVX51kJ6AmablcMgbP7Z+wEF6oy
gS/HD59upg7WfueYypLMLZRi3HDdMnExhefYMDLGgkwU3Sj2yvqF8hH16feBDgW+
si5e6NL+0X/uVInHgk8gFDbyp4wxuRXSgUnlSNZO4/tbauCIzLFp9ugzEYGPrhYc
Uk6mO+4S0lZdAiuvcZgz/y1j31vuetupfVHNCYWOL1yXQgTMgiVuP5CmecQjxsCh
VPDeySNqN9ezyxbqI/L0GAiFsqVR+vhrcmc/GlngT641RKezKlxGhLmPLQYKuJJ1
TBRGr+JV/7uIfuPxq/Y85wEv4bF0bZ9W13QLTT5H0gUTvG/XZGW7KlJVX+RgjPMb
cAdmZWUypLapIvBBx62ovSUmjgjp8hMV7LclKBUqdPVUkHb19ZrM1FxJIqO+Lr6r
erW6s0jE+Xyg4+6c/w5CN4P6LPw89yRSrOZ3seIBRZjKeBjKZ3Ht6AP+nqhtYqtb
6uLhomQbwjKiscx90tYFFUKrprxHOqnAylmgL3KXpu87tOpMMFnmQ0CS+bwAtHBG
SkpOYMpwprFXSyKdk8+mpzstIqSKzKWDiFsK8f/8t4OqHMOrLJb2hfBKJ2e83UHd
eHW1BCsxjnu4gRwZSuN/U8cFlSwrZdjAX9iDlqI4Im5Pv4RwvXak+TJSkqDP1qCv
UDGzhAYVYQxJ/lWRn0Eb+NvOF4xbhKo4w6vpz8ZFwTm3GNmD9NpCUzCjOdLRoji0
atVdwIFnG4o2WdgWZIuro+tDZBpwFfF0ghsuxsP/RiW8h7j+Zx0OnlCvmUY2/Ld9
q7jM9L+A6JFiZ16JvRf7ewigH8XC2eeQL8JhsZPEZsBh0bulB1UFfrrMRCEULJwB
RVLFQ87ZOOCj8IWRu5L4jWIowWjstFHkn9wrZjHPp8oubTNMzy/YOUorW0ciok5B
Z/88WEi3JHpbllAfNhRaVDj57ENJS5VZTnxS8GcJPaCpzHCmI671U5BKTo3w/uuy
abHV+n5nhSWVvSipji61vw7/exWi9W0lf4JJarBJTXDhnVznuJ6TbuyEJTwp6fK9
0zkOLjgINaPwb/uHQ945mhlSOvDZJl71xzNtgq/PVg6CXzHWANxIqwdFnf65iZux
rSN6FxY9/BVMP0Jk5ttoHRKUu/WOJSf/OZ0uRHOAsCF4ht2YWiVaetIoOPSRKdwQ
mwSe+oeawoQ60xHj+/CuqN65LwkEcWroBoslIK87wNZRc3sYRIWEzEAS0X4HHmh5
ZDLj8sXAmqR0VpjxSoJ2wIhCO/BGULEUuJgTdt+8xRdIGxdcOjdSnyBlwGLMGEYx
yauSqLSZ7TN1tzhnRMC2vv+5vqxBqlqsZncs+kntpifCDGcbqgBR0Y2prpeHh7lr
TZt5E+DhH2r4KZ4WBsUtCVghQl1YX+F/YmhpzEZH3ebGL9r0Ai890pYQaJly5lnM
s8xaH6Ln0gQGVgvAe5UVQ76aqqbqBVd3q13n5rfLwFiwMPQUkAHyu38Vci+nOvQK
+BoEPLCQODrO64TfHDa4bfLVcN/LZj1xZKaUhfZPMJ2qRKSMuWFGSZ67tBicjYSn
k5QtvANaQXvH4019lACFEY7Uk/ZXghfSv83D7JXDXrOqNz8dQJA7Mg8uiGXlhQde
D0uBN2um8XYq6RSPS7nI31eAmvhPMlRUZ3a3FSaOihc=
`protect END_PROTECTED
