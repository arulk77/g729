`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48u5dxJJabs9aSNscM4cgBObZA6lxrC1C4n+e41CKRTS
HUyf5mg4er0jqbnrVFSFIquLtimoUGkkBRKTqmbxj3Iko8bNL1XoxNf6UXv2uBEa
ZHN42P/vi1HpNvu3Y+bHmBkngw9A/MQKD4eth7RndG9pNo/rc7KHmOdoriDKUk5+
BYD6VFE2bJZbOVcKrtWQyGChKp0zUpMTg/PzkGjwUdvLRrGYQQ1gHIh+MRYsf9N6
DyWOZBDhFOSn6BIIQ6MUq1ukm01CeONcJBSp7ss/2hEsx/8wAhwnXYawpyt6wAxO
ZHBUFMcJs6+ER5MiqeUpevuIzV5zNPLB5PLr11VerRWoqsgIAun2zRxDV9XaXeGS
Rkh5yBZjxVs3YFaJlM+eHw==
`protect END_PROTECTED
