`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBISXg4/jSwLxKfwjmwZXrXDYs2QMTVa3RonTUYUADyN
CUWnLuGPpwDi+eShzTZShmleimC4efYvMzsYskldvGgJf4zKp1SBLH94H0RByhcf
lySNbBa+1qcOq7qAISJFQ9HOEV8mGT+68v4uRCFCfNlu7fGVQU0a5kSfMP3s16r5
+KJO0F13AieJz0++I7xqIFe064plf8zB9s1DyWMW3Fo2M5bWc+xeQPmNa/A4yJrV
VtZvC62bUcA4y6I2jRP9TUmTJtIFwABUtEtvKQwF0TAEbFLi7DtFtBW6atkWUPUt
jv5NKUhwyfjbu88MUL6D+g6nEKfZrSvP61bqpALl2go5+nKlwcAShpUwSAObG5eQ
`protect END_PROTECTED
