`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aVz6i9238PQAXXPgG8oNAAiT5YCc99fG9uqmoyvi/I1Y
k/5cz+lWmWv5pERL6iJKCIgjjGk4w895muJQwv1/MJJiSCaXGvQGtYE5QPAhNt9k
shPW6AYeVyx5cJ0BVinsvnP4nRDM/k8MV0s8owiH13ZEMZQX992f7lM3u4BL+AKn
hD6Oqr6jNjrkkWkUabPdcG9x9Z7vhyaLZ6tShqe0UZUUNYLe04s8AsXODRwrwlNI
CDKfHE/fZlfoFbHYAHJWlWOzmeYLSONTpFwIckwq9qfkHzEOzmN517U2pTP+xENv
L3NPYntOGOmhoSR9bS7ZhrPNjCyQqTeuugJ0Qm5JKVdst0pv9K7cgZKjocgZp+qC
`protect END_PROTECTED
