`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAcxThDATvHUHuqzN0fI7QckjKDhRtED+n77ZAetFfus
8TwnJuVZfHiY9VDOcn6Km+CGlivPs5MwwNjlAtxnO7e+ZNA1crAtp7yorTyWVuGo
ZaQSJ12nJnj6WGKgJyWutiVvweKl0V5zkvr0Eig5r8wsOfopFEkKlu1BqizS4F28
ntEqN7or1jXPypAOVlOKD6b7WVRtMYB0Kt28QVIpcTqLNOd+F/Bo/yKRTsXaLnjp
Id1fEDHNGBK/Ihv2VQ2ghpW07OTs2K1P3HsipTUDiVocFmfpH8QDgUeqrZzdugxZ
uK4f6tFT4ssAaQFnQvCFZqDhxp7whV+jdSKlo7V4lNVdN9BV+eZlHUIy0ZToc5zn
f0P1MenjTY8pc59qdTb8LsAkMVynj9alLjSKgPQ0959eevZU+4gR64IHRJdrYo8d
3ekDpr51ceyUTLXreoHpa5art5H8WQgMIvX2xwkb3yiNvblvpUGoHZ4FwyBBynt9
PjJVeTc8yR5EqCn2mtgWa33laGDKIi/f/V1TK4Jwj2jkEgeRO/VL5CC6kQiWsnmD
26HUueQUiWnz0nkSVKjr7eEzXxjL3v8AuyfBuMTGUK1J2KdrQJvuGP63g5Y19bf1
fVOc0BSRxu4rZbvlNZLt/NUj+TKs9PvynAgMM5yDBCm3PwuVImKVeDE8MnD+mYJC
H66vR5vUhiy5iMJ0SPKOcuv4VVTMDTpBnbH9oeCdwKGbOafnCTz6fHGAVKloHXdL
VLjy/ey2IjM+LTlUR8WNtK8aRrOZ3kVCGW0gEAInYvjsC6XFcSkGPr6UGkpqmbtb
wdg3ontERdGIkuqmPHg77+Ep34osvn5lePbfsr2aKn2yK1wTGNaPvguM2nlMrrYy
uQvdZo6RNB8Zaq9DrX3KTxAHfot8xoQxhzKaWvUD81R1RzYWsIED8gnrxRtZfxKp
CKS5Zg3P3jidY+o7zO/rGSXk64cdRHbFjpcEs0iuERNrpavKHrlhsqZsuiy9qL7G
P3lsaHtHkTw7Eneud5qXtq1gwpZP0eaOEUTOmigGei91tWaRaXEW6+l0wwyTkuiF
FNaztaKbtBEzpH4JprgvZOZ7iSFO9zCVaQAwN1lWDBGi7uHkTqiukM2ZyUvyZOjD
VeUCUQ+uqZ1dWrqaRF0ZTIIsuVl629RYMBkhkSgSgBFKSdmFVJbgB/MfUnWAZIVi
kpn248cO1P5zC2vs0JI7+ic6aGulNFos82AEVNu8QaU7wMeIYext/dw1ZlkGswyL
ZPkFbqiuudO7HwhwytT6uXDMlIweK2GPkkEL4wTZQzelPdxl9sHUcKSO8gFNAwUX
3MkdS3fXkOUWCDp690fzIzU2MfAHIwsfVozbFhUCTlgb8sLI2DW2cKyNPYPnMl/X
MGcd5kaLUPOnlzcocRk4CosBBkstz/Zz89sL9xwlj2AZMhjUHFqW8Ea+qBbiafa3
ThR+8EdGlFW6sO/YDvKjAT6Q4HPaY3YYYO128IHAUrSr4NUIuhTRYVnxFqtg5pAT
wiiPwFa63UTWwCPO0PB/BrSyUJfizf1aNJOYpI7FrCKVVequFRCrxrfTmqtYs5nh
ergl65VaoksXrIwsQyn+0aLr35uRC9U/UfXXWwVlePSmZrWqK0tFJjXhcOZm/RNw
G7NKddr1lABQaAmQ+umcs1EdTWhjMGtLCZKw/JgkY4uCT0Qwq+eI35djVrsLhoqu
nCpOFpqIgJtb/HP+GY7zVq9IcdRifF852f5pR7WP4zVz2Ss5L6txEwE9QWku/2Yj
C5uecwiINllZF8Jg+dfghSD0cYaIXaTFRFc/yMWkn2jEco5jN5xE313bj/O+kJYP
9hV/rK95SMjFl6F9xs44S9XrqwGDUoPAqht4VgJ7pDOqDAKWBnowM7miWMek/GsM
v2KiOct4UzTTpJzS8majZNoHws0SmWU23OiYtdSGCZvU65LmE4yWf4+0u+Kfeuwe
MBGuc0Xp/t3DNC+wr3QMSv/YUOb0EuobyHv1kQegh7eD2E+8n7QXdEU7pev1Qpx6
ED+f8fFu0x8X35/yAzUk05M/FO5eatoBNFJeJX5D9tOmqEwqXbxIqKPblQyjsO3D
4uUmRxsT5FCm9+JYZKP/j4f1uKevdDsvuNQRonyUYWbKnImSVA16YnarP8qlsyrM
JuVDG5hm/XLz2/XHb/UfB/i5zRepi5u4E45zMdcS3YcG/dj86c76sl9kdKCr84co
HJIUSOk1j5B+F/M4ZF1eKbMGykr3q4ok9FwNd7iULX92Us2juWX8xrqKfIoGFQ/N
PUeDocv4w5IJ02v9DcOzJK83wmk6n1bJ4psWNsnwB7oTP5nC0SHqEMgj6Hy3NG5F
`protect END_PROTECTED
