`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49JraxTDFNbNWrQrDhykrmBvzXhHCY74PQmR9Yxrq4xA
hNQwssyaAjOD6Vs5P2X3xoCZEwAlAMBrsCEkCvdLgJ6ZB24pJVLHmxmV2D9V/+vc
Rn+xXyfQsw0jxePHu6sWTEgi0ZbuNB58dOzLVn3fJ/LuOE5EVS64AgwXqu7wMxa9
pfG5AIlMHq4doI7bO7hPq1dwUZhwOSYpbpkCF/x8qliiYPUJQPYx6z8C/FoFHp0/
+smmPxBw1y0ZoWTonn15ETVczygwlUOJTpVH4NOxJkLAzvlYjAuVMWIqRkRQBM5p
pKqqQPRBWlDqjvpcRa2zGOlK7vwmD408VBmuRpZZp7oGOIS1H2XNV8spq0Ibs3UZ
MsXRHUy83e0l5MidWR2tLPYjTMwrP/FAdCVZ35lv25ZdyIS34kw3v+xUVRGrVhnB
ovkSqVuGyoj5+E/xZpOdSb/E24Fejq+ZxRKuuUdopfpmXZJBnuFw3AcQuemSuZLU
`protect END_PROTECTED
