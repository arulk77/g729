`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
92HhI7KAyfBKb8hRGx6GfvcVNgQ2pqbwBmDRQgsb4iuZcxJwzZkiOqbUV3wbKmN5
cefSY8WgnTpbupTOltqOCBHHL0FkUZj8j05/irjjnUbFxcyW+1g6/6uy9/uuGddQ
F+cazktVCGwbCK/wjl5ByBq0YsfVYUzZaajEp5erH9i62ixxw9NTn9jUI1EyhKGg
sEOOb32mNH638LYQD837M+dgYKqt3SXs+ruAC+3OONN1uZ22/dJ74OYT6ZfKL2ke
kxlx4SOn7KM/QvUFg1DGig5fk9nkW9QVvKUz6dvwjG4=
`protect END_PROTECTED
