`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIbVFldiEPVaQkF85Low6SFTK9mNjlhaAj//6qowlHjG
F85NAzSW29axGIVj6hBfB+tLc8YqKGIF8XWEgxlAtiF3lDpM/b6nA00yyzR4RwRp
iyjaJb2l5rSjpQiQBUjk0lCmRB4Li1Wiq74SI4FYluFRe5K/vMAmXFUJPfzas6UN
h8TQcTx2Vup9cms678+m9g==
`protect END_PROTECTED
