`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJmicbl12FgIGPJaU0ku4AkW6Rn8AOkukO+j1M/HU8Hv
7zraZiPIfPwRS0MT9YRRsWndZqqxYVmrhmIUhGS8pEWVjtrAT5vGFfnsVpnjh91d
pYE5UNFir1Y92DO32haLdWX8/t2pOzwwF46ZawPVPHdGVkpGJj85qqwZhlFxGUUE
7VqjthG/DBPT9ZtLxvWHhg==
`protect END_PROTECTED
