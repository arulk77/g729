`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKGHurkDN/FWq46wMUOVb6NOSZAQZ9NOn6nHTf3vdHiJ
d7S0a4FAJs68qVTCdKG5wlL8DSfBZGIek7xhUFYbFSt8tMfeR7l9LusMUotTqKd/
qT5q6r8EtqET5eq/LK4Toj81tenChNPXJVsB32tI7IQA4+OHHkar/c+aQQL8xoAO
8xc8vPk0WpjGdDIVc4idgw==
`protect END_PROTECTED
