`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
LAlJs5qdnYnVEc+NFIJFRmF0KrksHUHyESYfnNP7LMl4yuttcC7oliO2fykX4PPL
p+G3IywwT96za0mEU57xxhuD1IS+H0qhAQF5HMOLOEzqou9TsWCkDsZ4q2TGsC/H
gNz+OELq1lB0mMN6LsSEaqketiYDmFXJu+8sO6+gaDrxieZx/1M1de/1dF/XnovJ
p+9lWT1BiYNQ0K/Ld2YLt0NF2rMP+6co9Gh4Tt4Uz3dTCpzD+MlDoPA8u7rNLLhM
YGbsowsGJhMYuGF2Dx6eZ18N9o1D8gaO/+QhospvmLaC/CiLZVk96olDVKivHc53
NOilxIKrNJo1zcupiN6aoy52UkposmjnMPa93b9J4IRFFKYVQAR72RQ7xPIR536/
NpWgPCVRdQmdOljbFATopyXI3S33pdSm15Qr7VGzV2ULZOZFGmyz7gTWteBcmRm+
8Ry1Lxn12Ie5y2UA5z7+pf/sDiVmjeYHO2d2BZvIgtg=
`protect END_PROTECTED
