`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePZbQyDZ85yX4z2h7/Q11ZKdmVn5PZ48RucgUpSbJX32
0QEgOP9z4NA+GQH+X2PwIssmKYFGAMeCU3I+Krpd2KvUyDay4oFua/UA3s/GUeag
SP9zYec8PSlQorwRNOgtpbmqjKQEL+KEnt2HEYy8s49kLDCJ3ScNXg6L55tigSe2
CAL6lfwTE3Uj8Pjb+FNJoQ==
`protect END_PROTECTED
