`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB/12SKz1FWUuUJos23gbF15FjOkkDUQwQaxkwMHGjVP
d0PgWsJFSDXrKiizvSvY206AYuH7ia4T0RGwLMHn/eHeN/iw+qdMN980zTI56Bg3
weQ8ZKjXK1igA6VSlpOhRT97B8FfA+RHM4UCAzojdyd+X/FxhBZ7AdJz+QbojSLU
6pzVm5Uhl9HzFaoowkk1pQ==
`protect END_PROTECTED
