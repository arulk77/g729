`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBqConBJweKmSI98MUbPFNtF3a4vJiVZ29+8xgYZVgej
NmLt+OBwu9O4zg5BYGKq2UkZFftpiuocAXbZSfkBOxVKgAsSmUsLdTS5tWHIu7dd
Nfi1W8GJjKMW4e/frU5U5vtSL05vLuaE8vgnbKbBLaF2j8wrcFW9LWpYO6V6j2FM
oehHXXpYHUqHrEWOySeqJZwrf/2uW/sxotTIxgEQLK3mIFBjQbXCxD+g9SJswPSe
emi9SklfNGpbWkWlyLEaT3UPlI2lvhGzkBjDl3tzpzj4rA+MiDLv38D54JwEXXoy
AAdXHghU3jvGpPdizhp8tg==
`protect END_PROTECTED
