`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI2cPEj00dBBbr/e4+Bjox/7uqjHMZnLqDybEBNzubS0
8zQxfkrNhctC3CavCcKKU9RrxVBg/4JPeo2QGkuwXZRvUTNj5B3fIJDQT6b90Fv7
i804ntSDlY3dRHUzcgChRXtuFi7GMaqCYotGCHa710fq38/E3DsaPlZ5dYN4VEiP
ntLHbYSjlL9qqqBhHEuQI0POBPxBY0Nn96GdF6Yaw00B7Ozv8ekiA7z9NsiazClf
VXT0vQ9C+DRobAW//E9uHdX94/cmzwdGVfAEeTDYADDFQt584heo6xkcdhlfODlG
B6XPXg2kFUq8INoYTg5gIt7j+oJ/JsmL/XDekUP5jqHURAZrZdTIbPKaJ9q/mPzi
ZZTRqjkr7FMtA/GUF0FMIQeHMnISWmK3OpCk87vZdwf6kWZOFjUTegQMHGRgugCt
`protect END_PROTECTED
