`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMZKpDAjpLgzZgO1+FNBm7wZiJvWo6x5Ayk8diTDXRrV
Jb+f/O8gn+KPOp7BV1ZYSbJgL/1KhNKjwjLuXAlFYHlus1qZwNXTd7CKTCbWdYF5
i27aGoSkf3mr82FOtFgVZFMaxfEe7FzfAf/F2F9cDNimVwfInFh7AzOZ3+ofro+f
uKciYYYxAOeVfb73s/qklXAStG2XfC7V3R4jUm0TmHT/KFvDY9GXmTQlyABZo5E0
9cCv463RKckxkQJiezbuomv5QFPrga0wyj6W0jg0T06pdUxV7LA7AZjGHEQKJKJz
tYYyVDddKICqUE2xqFA7XHvXHLG3teiDiQ7cy10FN40u6aS6D36uwdcB6TrkYB4A
S/Gy1V8iPk+au25c4xcDgp+2JVX6kd7u0mtQyITPRCw4XAcWaN+54Vj0wPRbXs6R
28CfpQLVPBYj18Q1lsdgvv/Z7rv4zUccYGfcIOqvwU0j4zaHvDsKddsoktZh+bvY
eR8pZcProKBNrxU/qXDUQuWl0yn9mHg4wqHflQdHkpyNmm2E4/jnnqqjKS/PHaNc
`protect END_PROTECTED
