`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNwnWQRkkf5CCX9ykzQerGzTGCvjq63Nw+qfljOYO4OUe
2BW3nIwpSNhmXJ+qxWH0tOM3aOiLac5yBkWaDUAu2nY5gK1weznosY+FcAWxrnwZ
s1WvIEVJZBjnpSgsRJb5zSFr9AxdZiKknUOKYN++buLv6XJrjfeHlYqHZ5BKDxcQ
WW0bxscUUVVttFCXsjWqEI1b2MRW6LEu99q2p30BLT6BllyYNplyzL3KBWkVJsCs
trZnd41w8JpLhwheg49g79qra9kmhzeSlhUWCguYJTxNbzTUTJD+uYG96Oo6Lahn
+fILncFdDGySktBpRxp6Ajl1sMkC9MROfaPs5vUUorQtgYedRXkVwzF3/PMh98ln
+3kz7EEHhand8OKGsik7CXesNh060opAMMJViKkqTXedITfYu4s+Z9tcPRY2Tyb9
lmheA5+VLMNDVIWXW0BeD1aXJPJpTU0q0R96+VJ70IuqZCMeRUU64N8xXQj+5qRP
hMBJs7eelPNu+VNv+uHHWdS5VvzHquK7wUAWUs0nPrntE7mGY6eI3UNDYrwyxyy6
DHQ8CJkde3BjLp5avRvlCXxz0veI7oClkqW6jieXC5+YKoZqoxYohSe5EOV4PkHC
XXkgK0PYn03N1rq3BxfQrRW3L91VrnO+Np+KWAIlqqqe2YTObwAb84KTxz/R7rf6
5axrs0CR2tnmdMf/3lFPR6T4ZpYdROd3TEdZlxIma1OvegvN0aLiw2ySAN0JGqw1
mhH35zof0VHKB24X0MnkbR4+zHCfBzmkK+6QDBJ3PqqCgdLpu4C6e+iBEWy2iEGn
1DxRtw6RW7b4qnZr+hg12HWoI6htH+NQuYkwLixzIK76Ut88emL96dLDmPejIqkJ
sAfopHo1equbXfkbA5TLbTZ//PlHkRC8SBiE3CQqkUabOkVz5HspvVSHLoUyI0eo
TlWde8I7IYeAsAIuFv4euj8gu7jV83bTbt0S/YShY7ZbOyKLALJYCwo8JYqjqp4Y
uTYKAnqvjQur0bSl651cjX3+P5BemXWYnG/Zg+LM3jJdjhYBGVpPAil5jnYx5lMN
Wg4SnTy2WX5QLh+hJoVzTeZjGaZpYrPDF4w+ecB7wgnNnwP8qzcRaDsIQgBW2sT5
oONfdVpfE4JBZGECDTQwytUKQHDZaZuqMcESkBMf1FVpnxmx8EWu0dJn7SZge6Cs
mZ1Egtme1G0cuFADgmopQh6HPntUMygk7Z1m5r4QknwE5A2V+LHrwYLchLnVPITK
9hgGKKX07YKf9S84QN6drW39eInI5/PkmpEzVmYSG2pmOZfaUn1KCr3n+tXK/cx2
ktQJoKwDXfzJ+TmjffG85DKl+OGyOzJ1FN6NO/vNZSdeJYBm4f06FCbtq2BIO3w6
fUc4EqVYlQXZCly3CYxyu+racwkZwf/4WLb8a6hdDnUoB7LhvqLTd6NNkKGgS0rr
Y9kJgY3Vj4c1yOxXUF5s8QuTrHlg8SrFV7Zr9cRanCcXCa0ULu07iFSz5xVjBJod
Nehhqu9/GWYOis5yt+K5/ghbmr/rspgh2CAP8qhhgF/zkAShnd2k8BDjRLHYEPMT
Y5iDkmwfKyevwnc/LWLik6gxhVbUT3WdwlolsW+odtyAU16U+8hCFbZUNgOQJZ0v
Gcq+BSCrGj9WEdaQylOFNRC6YYZkPRo4+aw8LVXJLHPLoYBoxsUXZ3Q6Tp2/8BAi
LyfELPHFVuzbNyOSh3jDjY/pmS4Duf9a59cQjqTgbkHZ/AUK7r7IyGEvf5Ln18e5
wm4EcDyujQWMerRzR6CUQY7hfMWVwjSoDaSQTx3Kq6BHMu9wpCpFkXyIUiTb8+Pi
BFR50P66HmZ4/N5MoWmnkM9p8ZIXxpbP5BkXbqQa62WWWzrZCHFz1pVN338lr/fk
5QZduwmSEEI8shNO2cpVuLfmPNcgNRaXXfjJoX5a0CGgOR3fzbfGuSU4NMvlbZjF
iC1RWQ5vDSIy/2UdAnjmtSxjZv3Y1yjpCDwddX0RtTpiG9ySPXy2ofGljpgZpQfV
jmGKiXX6k2iynaZfdfRiZsT5ScnIjWkpYDaEf+ki6rj3YFz6qPy2WjhQT0nxrtkm
qv9Eqz1wTF7HpVrb4stbn7aEkL0K2Vtgv8lFkOOmxusF5cWDN9fhyfHlyUn4ljxt
um1pDbZ1obwR9kcjJvssZtd0+TxwUU93Uo+Iy1JQCMNGnzxuL/du+p++C72HVs3j
uDMJ/ib0Knxm4rXas/70w3DWDFTiGa6BsCuMIMQH0VdJl/vjD/AvVtpu0k73w8mY
tKzIptpRxzgpRVb9jGXpGH7vY2WSaFyPyuA4v2FPe8Pg1mZlxKlXvCRINwPqQOhr
5aCzyKbmARrZSmMG3QgGES7KIRPkoM7OfS+80XBj/k0AUf9s5N45aqt/k6ZmTR50
PCpKRYXXjaQErA/2DFxHFcCR0JOqtQckccsYazmjaoxS9Yw3mBdK1IeB+aDhcAKB
jh+BqojfjUu78gdZMzEmQB4xX2JcIWpzuMRGKnMRzq6vN7vwU9+emeGrxHfm16RL
witIosQa3VA6t2blZ+dOa+HxQPEHBsJ+zG6qMt31RjN1xuG+aYgn5eLA9sp1uwXr
my1IYFmDvG5o5ZrHzsIAz2wNgBZpFsWStAY9rF6jnJyWmeT50X42QAFFWnlvAach
SY2TCOgmQLoS5iGpjRrru1HOSdmJGGdzjVhXG9EVvgPravHgV+9FwfrbYnI1917D
tZSjjD68FPTzwg8vCWphfUGwVnOf72TTnlj1YfjmeAYRvMfTpoEzjdM/YslJ9Mlf
NjvMJihKK5VfEDEf023smxokb6QziXZ8E6rPQBGpLVUi5DZF9+Ad0XDX6SudaCya
Cki9Y90IPH1thqxj5VI+OaToD6ObtletuTsRmurDdga9RkyqHxHNG3GDM2gmCJEt
ex1/NepQvPYGjT7AsYbHfTH42IvR5aQZXqedenRaCrH6MY7ploHD7B9kJ5vO4Onx
hBIo3Zr6Rk29Mw5hyr5XzbtaXxybiBcgHuoeOME0RsAKHPr8p3LKgcsPdm3Fo9rV
fo2bKg27k42c5Z0uagy8TVUHDa519+2jlVitBziUXsXBhZdsZokMuqLdrLeBAgSY
3eJtkJp/k6t65czxei0ZlObFT7s7VkBs5wgjsPObBmxfLadDwtf/PZnfxVFnY5y3
Cw/G2tkCPjoWDWLyLhER/O5sIRhImCD2YDbxndPKU6DF00kwavb+6QQgKm7SeMdD
bpWyltbejyvPkJQRqsFoELkFG5ULUrU25rjmKuz8ClUg65MdB7IuuM/7/P1PmjD6
i8spR57Khw/P+LezNrInPUZHsnEpynZNm248fA4gwPaETAA4mPRBjP+p4N4MAAlk
ECby6zs8ZUEQl9OlvkgEyP5I0kp4n2N5bSmKPCk7lj2uEyJKQZIqweVnp17KJbYH
4gCR1mySfYmcb0tyg8nmdu6ahEmnW62juosqGj8iNsvN1ECU+NYtwS51YenZuqmN
W0Fj4cH14mDRhVfxuIeVeiRLacmoov0iNJQw/5MS425wRCfNOXiRXY19aLNByidJ
isZkxqbp7Yh9NQF3zjW46468KK5i+4Xi7n9zfkA+dhPjVt72gv58YuOJZNF+GhmU
GxiNKOu28X2c6zfkrovs6IWeOqaKku2YCPLRNcsoty6bgfAwmaUzNpt6BzTte5pY
Xh7XZhWoUOt5BZp9I15FcPXC7a71eUUW7OC785UdyZk0WJySl5fLJgpi82L4Dgd0
bMbUVu9m3Vutd0U3ZxHe+KjkcyDotcGu2WfRB0p+1yfYGAjZF6GUL0ML28V8kn7q
Um5ca642xa2dXKqA2u1RXi4fbi19H04cBvyE3Hh5mKYzTfXgDayNs8tUIWfyU/09
6WRalj+Wf8SzQEbABr0yJ5HQaF5lKAXkhpinppG+YpRv4bLV43er85iL05AW/lvv
cq8paq/+T+bYuom5TRhM46UESIW/ciDB4I3KIE6Kcx7ckkkQ8sCgiuRcHHl+Nida
GgGpnFcJcYlJtXQACERiKq07RAJqGDnijPaYoC8xMcpVWdeO5kUW2iWqs9aADPxu
N9BMGXE7dOp6Lnxp1v6ReK/Zhm6rW/hvGpY15/kz9ZDTbBWsUASkH2c2ILpCuT62
3N9z4CY4UENOYzT6+jHit4SSxhpvQDVmaE539KPKNvSSwrtSlkhWA3vU8Jw/n64j
+DhbLRjAPjfFht5Apw/EOnZD38IlLi1WEbjAV/HEX1sNFCf2wNrGPWInfJvqBPz+
G4ORmhIXrBIEWcAxVmH5fdGjPnXN1yH1Wci7AxM+rZybpS5lzFtINQbAdzQfyms9
gWCyWO38gAcNGA8wWRwEqXAzvBP48RztUr2tA2i+N1V6rMD4a/pRSnriQWvsSZZh
gGEM2qWkykUKckDkbWoLXSFCPRTNDrIM8cdeX4rD0DvTpLBkEwp4qVBn9n+YdNms
tCbjdyj3UVQdUVvytg7wrsXw4HYSj9beHeQjhudjqfKFANzdeH2uCYEDhjfY3Agr
SdzdoWO+o7fnqabQVR9KrbnU4EhJgniBahAVCtCcdFYVgLivzCN611jtqLJJnLty
PZmczHGl/rrC7XxhTb7aF6DyjglPsgvplevfXfqKtY3QtfYkeNLa1N5pPgH3X+h2
g2WqmsY83g4AkZ7kVmx9qonPZXAxJsyQXpMZBVmmvnZ6Tgv3s+NYppv1knGPAgWL
ionKVxpePdsQsG1m3X7zEvVoGVTXDL5uxgLZzd+M7gUZvxFi6WnswqB7kUy1pE8q
0edeCvrrXSNQqoZLQxORznfEVF2Bh5OOcIowGxpTjm/BzUGViByKclDZmXSgmwNL
rsDdBVlve/XRHcbTZ82cDQ+YZhD6OlVlhPIj6t/SjECK0D9sVQRwMECxHYa383TE
nLpYjAKmLCU5DQ36URvzBJrWA0HSItep75MgdglXtWovGiWe1G2IbRnZaPtOngkN
C6bv2V8JSrKSnN91aiV4Ki61JceZjxXp0lOY9Esu0iIeu9wqZjIauz35Rh64nXvF
f4xZWop4yJle+N3zOZhxUMm4y9ITCvd9GbF1kHFL2+4//b1L8qtABQoD+IC0nnxL
XiMGROn3fuAHSAluJosCjbw9SBXxgyV3YxgZVhFXUUv0QE8dt6rMP2bE+fTROA7+
zQcfh2nOeeNO/IXjSesF7mFqV9WheYkkjPkplkNBs9y7Hf87uX9flnDyJpQAHtWZ
r9qh3s/oG+jvH9eW0+tdNlL2LGUYJq1LQxHm1X8VLTlaDNXGJZnKNH1Uo93kLzw4
Z09q/3TP/6sBWt7n5iJ4b8DPFVpsPM+sudjP0goXdtZJwobQPNn7dkCrZ/4FvTJF
NpJCc5b8QF+v6a8O/Zmc/9t6cDydZGY9gPDUMfOQ8OYkCJCsHmjm9K+jjhAq1xPM
I/pez3+R7tZzgws2v1tT9z2ld6yKbOR0518IAXbkfyOE71nwvQFbU/qEQQsDAaKY
OgmlART5QQh6YFXzDVyuzibha3USB91ouEjhmOfaG0I5yG/fpte/KaCtIppXqWik
ebEWo1wyxTavXrrRg8lwtjOtNwuImXFyorckz2Ydb+VjATaQ8tBPPxqppMwzGpKM
t0yYy5146vhngtjMfoa3Q2b+4Gb4kRUdcSBciPPhrn58z25pcXSpkwY92CNuCAia
KqvSUuGLZiQfcHUyBrxujpAXhD2xtn+GcS5wDl7PTbzJB8PXp/EHqoOiMztKepOj
vlo43L+9OQKrGTvZO+vxiPVlT5Sig8ARWJUS/ULsLpTDn1o8zRVA9L8JrupL1R65
ddu2lPtRxvai3CUN2vKpzTjEa94AG7agSm0axhSsdpHKs/mUOxLudnuOQseeVKX/
63xtnS+MPKgbRqFAla7ohszh5JUhGh1ZC9RKtMNkiH9GqwpMvBoKp6B8tclYkQKm
yQBd0BHPDSY5uXekEib6qaBxXvok8jj9sPQkCfbolIbrnmB396ccgOOHTgP3XcPk
iuIH0vAup4wECXWVabE2wIuMjjxFTWUTnNR5b3shB4usu1boMgSMBJrHhSO51CNA
AVXQ0lb+LM5Rw6GPlwMMZJXWBgbVmcQYLkkh1LwjQt/7FZqFk385JsXfOFIxLpkM
r1su9i/FCEkd06eKwL+TRIHHFU8F0W+QtrEmtq7w4OVZQdm5DlCFHLYUybyOQXG4
u5towMdkYwl80CrRaQUyNpUnGDHLV+k020LGQEoUZsyFcgYGDMKgbqoGrw0gQgJf
lEAI/cZ33Xe4/qjh/E4wNnbFo1dzboiTXGAIlbjxNdcwpfB5fafjzh5m53BNjv+L
p2Bh8w2Gdac29Li/7dnFoIpEuUIfl/+2BMGas9YLF7jxKr+EMs/hpK4caTEbERIb
KH9wX2N8oi3+DAYXBWiAULDwrjHijeuahesfQEpDWpUoezFnDMFlG4LTalxIcVuo
t6bDwuYO5qvUHYY874zFXa+XSGvLormcuncRqyavTpfbpPJa9c7m9XFHAQZnqHNy
ztw0zv2HxcWwAVLxXffvrUQrzBLg8vm4smkynwx9Zfjym+zfNF/yYhCBNjOHQNXM
YEL9Nir8AdcPhdAgoqQiPyS9MT/WQndF6+tekWts/h0DsupcxRTlSe6xpFu8XCps
uNm6bTlp7ikPq/dze8nHtThylEAlfWPnxvXbCCYJhqV7iG9tjwA5/D/pgFxbBfuR
kff4q4L1X/fW98f1lERufvDF0rfpqkRoSQp5KXt3zYuTgmtpUZjAUR+RT83biMPP
fCMaQ7VNRTFbzYBKBtG4CMuVxSDV1Z3w4gljNtZ0qRYbpgGkSkyoIj7W6X52bF0y
ti0Z/PuurLVWkt+KsjjkhU33BN+5FONhJ8n/rhBA9nXM7G9NbtiTcvPWtdTKGNuk
x4wFm5gJcb8Wz5Gk9Zj6BF92dUGRQI+5JLaJKwYWdH05mly+llHpJ27EYoQZVH8c
vrInZZXH2twfTwPUHvps5zsuKcsFQGWzE+wDyc4fYtIYsdezU7ji2B2lXn9deKJm
9vZ0Dw7xF+gCTPYYVnHW4Wrpt0riXbcBx09bzY5/IixISwoAOQjIkUbaLADshIy6
nShg+cnEl/WedYhUGqppFxhSG//c9x1qNmzDmeqr51MwoESVWQOvCk62w1rPskgQ
pMZjXDJJvIgVyUQ4iUnWq8bJ6bASrSoxZRvqKkNNU9AZZone3ErHLMS35u/+zE4S
GdeLgX9zHhuiNTvqzrvtjAeSp5XFIBGt3i3WSKO4xYU7jz1X6iA56RLVPt7cNdTq
LtlXVT6ygHFbwLxMnrIPSLymzXCCc7YjB4hp563EvSz0QiJOKpJNm8GRZnH//pAt
Ars3t1scH2Tgwul9y1gzzZ1N/L+Q7HpxZ0IcaLgufu5U5Fzd0czOQZhuIUISKTS8
sALV0v5MkoZ3jp/MQQp6aRqXL1CGeArFK5B90gfyeQxAk6brPK8uvQ2FXWVkam2B
tcASibT4LjnlY9nbCEx8PIvFriR63m5anYt+/eC+SGvO8FgTtIROjE5XajzBcrka
hM05UU6Hd3dtBvlvL2M9Jg+WfOEoc2gGyoi/TyPwgQjBYeIlK+qsJrMPmkV1cPQY
P7MupwC7CoIHfZc4LxgpX2DhhC2kQyM2dL8AQFT+8BW6j+I5bcUnkXcQM+lc6HiW
79qav0lo13i7bB9t2ai2q5qQ4LvUwkra1LSp67hXmsK61pBeEhivM9xVq3GlEGEb
DfS54f72UDMXO9zaXsnebgKD6RUsUXE9wCxnix3hGWc2WrqvormczEBh0HeHJLIt
co6vZXsPbAcfGK459MJxkYU4WeNcUw946SjQnaAOBAlWPRyGUwzi9BfF7xuZ2RUT
o8Y+ZCbMBp65g9gB+W2QrJbXnjcfKaWnVM3Haa27l0cuvACj9/Ky+VCYy2AZRlWE
L44aa1lc2yY/DsqaeR1k/UAWdRXJi5cC0GbV1I9JjgGK0hIc6/UZeqFHMoVgv+8w
glEOQKcs0IacgZEfkZT/io+Fd1/k8kfPooqkHGDWcQVmJBhos7PLqQkkdIokCM6G
TxpDlFkGq6GEiRiIkr15UN8hEx8JFw8KBKTkidCy9XcPZmVctkziUV1grTgAA8MQ
NP323N2RZPWTZps+a30f56h621/xF6CAzUim/Z7xfRYwZF5Raq3S5iqqUsz6QklT
sJ1YLpPTPnRXaZEB2RUL+FPChfGPHKFrV0jCt1as11KHYeHND+DBMr9MVmO4RIGo
BeL9NR13Doap0qht44/fkkwPd+ASVQso4e9GkvRm5mnfJmMMX2MqQRu2zG06tm1r
CSbdIMxilB2vTo82G6nELrugN4l/Y2KAveC1JPMfKjo/2y5gTtbrj89dsgESjY8m
oXsk511XTo+UyyU5m/jOnBaDJSptSpacafG9rWOhghi41vAnbgGiUL/oPPDuHbha
e3s5EV2XHmBNNAtG1bKRtOkmGD/FZrVVnEEkglecakZGpHgmpsEHbNGEqioqRB+W
n/uVCCbDLBzPpohCKE/cdu6icSk/stG/SrmtOpL3PbMZ+5+CC1/NIHoKxUQp14w6
ftw/WXFbISlmolQ9c6RnuwLR95L6Du51JYz2lzf4KhPjlfiFrTpIcNaIOmEGEcS+
3m4N65kX6hVznI2zC8ZZEQ==
`protect END_PROTECTED
