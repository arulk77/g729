`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
sXdsNIO2llRMG67ACFG60WS8gGBdo4y4bh+tg49o8n4VbFi0TyKEd+LWi/KgqZTd
43OmHulFLr2Wy2HdGWtdDfY1uk3AN/Ll5tDslClwSwmgO2LhWltdN81QI5jUqHhE
2bKjleVm+U/NLrbQIL8zIWmn8mWAOAQtnkOOxJTmQQFkt2G3EAGtJlxL0rkJ9t4Q
AmydZ+IQ5Zp4i/OsRPlOcFGUHgpatLyZJfEWnZp3d88=
`protect END_PROTECTED
