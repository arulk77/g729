`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLa/RFKHoq8/B53olANCFyOnULV2NSYVRo6zEd9GrFpI
J9SjA+qDPuKNZMpFIP/L04WinDNrwP+J03HR3ldZ0luojiAAlf8xq/fO2H0jKSbp
ztyJK626HYNa3gpGDQaU0MuMvg0TO/xe1pmJYVEHDjYbbmMbOAMCzNrjQY5i5aqr
te6dp3TbDjp2aD0iuHtxwN1UIvuF0RumZmDSYVAeuvN19Oi1aNN5GOsGLNhJr/lD
ZmITd2fdaZTNeXLXbizwpw==
`protect END_PROTECTED
