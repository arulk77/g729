`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHI4oL6PeYm1JKSNOFVtcwqgfXaa2vXTCX7rdOxaHOYJ
MvaBX4d1O+wk4pci0DO0Ta0IxgQJVzG15YQ6QZEyjMBEGuH6Im0zwvUG02hYsjY/
FBxxyuETuQ9ShXOgsLdzDafms2DkAh/lpA7ysJjTmepkAG8wGG3TG7qOJ7fW3hg9
Voo+vVrFibWBY13zEYc2TAxduDkv5YICYWJdwhx+f5lBfYAjD29QxSeoIE98kH7l
uq8ksdAbCiZCVh4gllGlsr79nSykyRx+IICqOfzY9ol1RetYGj6xpD/rnkLGypCR
5urD479EQww6UAbXZYj3DZBcRmGa7LZhu7+hN+1hLUUVkj+6JJRIxU6xFFn9REuP
hTopA0gKluaSIeGDOef2GzjbvyPfkrdw7r5RpxbOd1BQM/DVGtlis8W7gEiUS97W
+Susyzu2nZJwp1RBovgvfE2CYMtUtqyTMqNxn7o7DgouUw9IdHyctAKyLOpvwuQv
Bu6fTW7N7sMfZka4sED6VqORX0LZRU6sMXUF3teJ09pPXKcAWdQXEuyRJ9pRpqbz
kgJTyy4M/ZEDEvMBOJuaOY5WKdnakT8fgeFdMG0y3lf7GZaeWchtcQ7MuXyPK/p2
PQWL+wWN3bhsk7DV7mzS/owRsxWeKbqs8Hfv5fd9j6S0tR4dBsL0yewcMtNnbyBu
`protect END_PROTECTED
