`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42ekC/r2NDXT7XPG31d6bSPXQm04+8CQBUaen0YaoVXI
K6pp/tdXxM0Sq9npGv9canpp+HwFFUgwOZdWSnAyCpyX1lZEGk9n8RyzJqtyFg4U
x390dPmWC0XBzyvDbiRiUuJKpZXRDk45VF/LEOGAoW68mWOHO9pNyPfxrPT7byAv
Y1QniXM4DBmjSYs/u0w3IKdnbUkPueVHJPHh/RPXZsc8mSJOvSMwFYEvUDcNn4HW
ucN/aTEbMkskCaiP2WC5FBnGpvmDytyMRitp6WzKlNQ=
`protect END_PROTECTED
