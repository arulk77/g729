`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDsmt6Am58sPgjHprq5+R43XmhuIsrg7ZsMEnSLbreA/
ZPOyP5OFQqGiJetSXxbhS0DroUwl6cZMjvRRhUdS9VJmogln7Ll2XYmvTZWqgPOl
8IuNt2K+61hMSOr4FguVK4HgJ2dMwsSQqWVYzF+9N08yv89p/VC3AhTXzoZFqF46
Mu00iiTBwzolrOEIYgvYaSa3A0jwjEvOZdT3T5epl8spPxCQk4/K+sJeOOiHRSux
Dvs4YgEN8ag0e1sEf251mYnsMxs49SwnVb9PvpsAZXiV1umwDh1moIkDHt0wo8+X
/SvN8A+7ifhE7vfPGXxTSDCK3GfLy8wPVmuNXZFrBxmeMDerCx3H3bbxVSXtxhtN
3zDN7tRSscfmNXzJfjS6MPiMw+laEc1b2TbZ9tkiHR0fHYumlEnj7CIsbLq378Ik
Fpd5mIdRkXhXU+ufHe/+G7GzZDLBPlRUk6JjwEgPrJciT3grr8YeNyzShMFZZfx8
Xs4h0165ag2uN+NpNSoZ7kyG9SSaX8eK/otwAUTTWVIqTJQwwjPasqXsm81nq5jy
+BL3TH1CqDRGLE1vdUT5RiYcXRAcq1tP2HlVFaWa7CttLyZwQMCs/++0wTvYYeYH
`protect END_PROTECTED
