`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCu58P3Nm/LON4ARnKBV3XEQoYqtm8TSlS2gG4BwDXoW
ZOJfPrPdgosdsRkJD789laHl8DFJQYsJRO6q5JfsHRTK/Qbx3IvenackRMDrVB9n
dD/A2Qf9xmK8gplGUnLPAWSDD+cVr1uUocf8ZjzhI5gmhoihD4Ccx9PbS02G7QOy
RL/2dnmC1shHJVSBDflLW0WOewZa907B53M5jq1yV+MPzxhijkraglJ7LJmXAq/C
eyzCcTxI7wPJSqIbYLzfqiICqR67SUpeNkzT+8ej9/T8HR/7Ax6KeNG+gNNC5AMY
ctLCL/Lu8wV6Z7Ij+8iJO/47KU5ZCzYxvte7ztMLGzDDoxYT3DoGSjbvYEQrAgYl
YjPIopNr4PDRngXNFxIC8A==
`protect END_PROTECTED
