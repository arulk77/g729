`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/7djOBBk/nYkk8gCmDLb+QwpiB7ls4WshUFOReOiSMk
TJ+kiBIzqyPcQJCw+umUzIsRQ1/SD3XesM8j9R37akI7I/Oq6M/dg3FApr8d2SyK
b9mFftLa4We0KAq9nAtkNadbpMmIpeQbEdT99B3lXIPDdl33vAYE976iaEoEs3Yi
lqyGny/omrhk9Bj2+TzglmMMW6Se39J1hhusdkOqi3M=
`protect END_PROTECTED
