`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JZPjqvXPgH4BLbrGrTT2XLVu/3PlYvmwZoseXgWKc/1xJpijP8UxTTvEsAy2uL19
7gU3E0KAi8HPIA1Gkiu3V/htSDJgJ/G7XV/IVoFL93NG0jRS/tHjivsQIjunXxS8
k6UGE7mKZc7rJkwPRQ3pLFWGlFaoDRIuIUPwh3Sl3j7DRi8ySCeHbCwK2YQX/0Vy
xmHavs5vT9s8799IG+Su3BXBt+QSY+BDL0/ou6vovjSsnJNJP3srUwM7TMMHznmz
ZWMH3cg2yv0DTtrSdQZJKxGBjrbr6Omil5I0vkXYANaXVTkKKjq85kqser4K3/HY
kE0C+0CkeA5cPT9e7BKDL9YVcc+cE1pqx1DUajK6JOXtEjmCADR514UWczhkkTfX
kofAiu10yggJ74EJA6NIB00tsk3P6NYb8BUj42GvLGosOJz2NGzUunCUdnhFzLuW
WRH6botot21V3/m5L76zfdGkRnsppnbnm6hR5riR1wPnHQ4It1RSFy3XSN/HwJyG
GURDFVLvaO+dyLV1kn5cKAW3ohUm1eV7vzpqv9YoaZYPIy3W2Tb4PsvG+JdhVtS/
3/UCRaZAQRbk78SC6zma/2/yDVMg9MWJC8n7eKGIuuwNo9ngdn7lGLfP97CW1Ib3
VPT5HE08+r73LWwHsboQBF+pMMi81TgUfE1ugOwCnEr5sLS+uangTdmF+OZxAYmB
uqw6wMz8kNOA3E/bLcFpOVnMpXtME6GKoKVZKNFPqBNrdV8oops4ztLV3xLoV3Wf
m+wTcU614E5J6TU7ilOdDu+3I6XJwFU/XrQlqDFs6yAx3OBsTlH2zOxM+INnvA13
kzp/o8m6jWKK6Glu3XLu+N1G2ksPDi5cOheXOd4AZeokTLrIzUzaHwwRiXgYUR46
99m83NVoEinmdOnzTCbdI14yFPS70e1n04/TuUE+7M1lWMBgCa+NafhyOSwAQr0n
NVCasBM/TvRxcCeAMQve6cItSeSnmCesGHgu9NeqiIhS+/LupGV8Ln//K1SQSJ5c
q0w24mpYvFkgit2vE4zfLbnP1QubTrJrUlh4YjibnGGNrjlnIQcPaydWR4JI2ixc
xBkP49ytKvB67xiDjG7wkJjQ3b26lIY5MwVTm8h6Zs4v2g6d2wNSf+RvH9xIxC9d
xwVUSbr25j77FWPjf2KajNbe3mIYw9t95ZMcazktlCpIz51WCEbOPj/e/bVgY7mL
kde25NfvLs7hkM7Dga0wtpWmz/hdG/SZAZ9f3a5cS9Rs8tLcoZBo/sjDchmbH4uC
EIgDx2fJIC7cVLCYGVAfK9GQu0oD3VppvxzxdbpURC8q02dPfppa8adJPPVWpqbE
EQU+yM/cupE1FqEIg2euYK+ruflv4Z5mbutMDgTgfV2Iqvdv9Boeutb2opotnddr
ziKYD2PB146SM9RKKD2mrHvF5k3Cqw6XOtUM4rMynvrZ003k5a5Zlm+sRTUYIr43
Jvtao3hBgSAPcE5AiaaP8zse7PgZGWIe5Qnv/nl3aF3P3mvOFaBlA9ZZAc8SfryQ
ySrcJEChDrQbEW+ZSaua7tvr9MHOLnWzupGwAJ/9fOYFfRUS2XmIml17Z/jiSSqM
LFmQHR9QHcrNhaIOEvyVembCFD6Cy8JuSRGVS0Bz6q3VLXGDYUsOX58vGqQguNlf
kfiyQ6uyqs+r2fWf5CiiuXSZCAQBeJnLynqaTi1k6BShCZABDeCspfK6a0n56KXc
LYSdkp4NyWnLqTbn+PdRs99HG6t7gOgpML/TCfBAOX8xSgSVH8ddkwxFDXnmQes7
4uDLTK5dPe+q54mtn7qAcw2QoBFdcimergactPyh8xPtZ+SlGxxHtmC2Z76fV9Ws
uesILo9QyFqBQdDJBrHTFX6tOmvJeaErCGlrJjjNJ96ZehJHAtQ1iKygy5sxeldS
fXyTq/+ZVlBJktljXaMx6bND3bCfhxXEz5OYxXyxdu+FjskdRQpT/+neBP8S7/N1
EsIwVzYtWgfhJRO1c1u4UHK6IcesALWIW6w3y3XcjsrReN6RBPR07hUH+enqdpoi
FHAyCtUTW0pw5I2/l1sZNYK+XEMUnWU5nakI/8lIMJtrKRPY0ovGXKolaRy+e3G9
R/epnITHPQG7q17c5vdmtMJV5FrAuum+wDqT+oW/lGlI/cC6BocaZ6xsuI/jQgUK
TySrOIZbxY7+AbL9G0Ih5BDzlWLkeoCNdleC+qCYuoA8rmpjaRcXRIjZ/hAOtZo3
srWedV4k9KCkn0XeLIQJxkqPuJg+SGJQDmmzhuJg11ygR4CboDpfY4V4JGzJYM2k
g5mY5Hk1jE9JvrUocOgjvBvcKW2m6TNgU/4DKYhzLHaPHwN4jeulXlTWptZKNqlF
`protect END_PROTECTED
