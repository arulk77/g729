`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKKEC+dZRXbMLQWjwAJhAKO3DMhFeuVBwb8N1qFVN5zh
A38pAz1KIyVeJt7zq9piyey96UHAId1M9ENKWislZPrG+FdGf1G1dzM8KL5Q61fm
23x7fLst8MgcRYoV52WVAPrh6xfTCdLi6iOJbTNTKkEBhwGbboMMequ08UF5YFgq
rE27RJsFGk9QVGgfC2NEEMBoxzeQLtMaEBFpeAuLi2IsAVXxsjYMrMt4EZgOm69H
5YGoZg8x+vRZ+jbvc+4sayO251zRc681AD59+l/J+bOavj9NPnefzbCXdhA1lrYp
iNyHgRhaLzh2MmXB50CVXtFsH27x+BRpFs857/D0RPs/L7ZGUN6hquUgETd43H4Y
1/pmGg0C3hDdCtXhpUIYWlG+gNfEbSScmb7NhQ+T19AOO2ifHQcelPJoX3vDHAU4
2lOSRn9nTPQv1JoSTYnKG2ZG3p07AsYSJMjLFzgzgy9pmDo8VofovtiMqM6v+8WA
ILgCEVWrU9sneI0aoz84lXydVE6K9q1NVD2FSbvnGZLapeJ7F7LooYQZ3z3efxQ7
`protect END_PROTECTED
