`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
LeZgzwBHWIJH3sFro0rgO8D6qQys/QUBHoXubmOP3FAV9MJ8IeAAu6wpSJZPKQGF
RA7ZS+pR5y1JqYLFr7Az7kVUAPZNDeey7dqo+ToX46m8XywvdTOn/aBYmAo/VeZc
KulkYCzVeJzF4ruqohawYCt9UIlrO4UtX1ikGPwtHfda3LJ16Js+ki0HLz8jqQ2O
CphoiBiMMG3pMHewvigyz9EHUYSljWFdrKB22X8kmX0hUFhCsZ6mrhN3DC6i9CR/
gi2uTL3INsopLvf8U7Oyaih23cJwWbyMNQ6SUDTVpww=
`protect END_PROTECTED
