`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCRXYDh4zk6hPP6zsQ3GZC9g7uijQNNTZmawOWWSly0S
Tex1o5FkhXW+WpGgpoaqQph/i7PYDy/lodv7hywj/3FVgOlVQUuA7YpB+x7CheYX
7GjIFIw9ogNVrfx+iTNJ4hxWwDSHBKLR/5Q9eKUAail2obcQYp0/2a5XEoNvCJiL
`protect END_PROTECTED
