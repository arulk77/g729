`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
CXDo269tkFVLssJhCUcbkXbv4Qj7nLrI/CMu0MUG5Dq3juMUBhmFl6Hkd3CFBrj6
BaWMIHsR0LMWlVzkzfEVBOLtDFOfFoGnA7Ed/Oqtmdf9tkT+GMV6Y1mxGTSFXnSc
RzRcdC6T6ne3cbk268soYw9yzwiqZ6g4m8jdbXDpmDQ7XblaS3NVCaDeUzO4gzG/
`protect END_PROTECTED
