`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBkDkgIc8MP1z4ccqWLJUJkyar6U0wjQjJ7b9dqrNPnR
q73gdg3PA4vf8RJUDFnwZq+FrN8YUAGprLvklmgF9D79SWh0Z5+hfV7OLXxUBETz
/vIbpmqGKD1ohffbNV/nxx+5uRSoFhf/cou9vmXFukXCanGkRZXQFqDHA9g2jLhJ
4GHUdFc9isqSgm2rkUxKXOKtaTHE6ygA4MhM6tzn/4FPzzF1k8kpmok7RSoDGyGb
Fb4ri87mqjOvk0cL/oNdT6yDhM/GSbt0gu4+eiBjzqmRzNFKxQziec4OJWHFLdcf
dU45qpOsXqA6V7nH3fTt3v5Hk0IKhIE5XOXfHxZXzk2KEj3ZoKNC8LTyNkmdvmwI
2hAyc20AqtdRZGY9SiZYc5plPuVegMVCw9lYojXlZ0mVAvCr3gt8WvZ/x5Qod0+q
9Wj055k3uNokkC6pMzvb8xjj/2OOp3psCZkyKjaVkzw=
`protect END_PROTECTED
