`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDrYElL4mUeW9W7ZpW2W6P5yDj6wWnX8YTFjPR/z8WcO
aSRKGT9R1GyYZgeGws++O3g4vENIMmXLmLQjLFITCLWxJPISYNdVo3iYRO3IeCWz
2PR3iFUisMI/9y21M1k+rFxwzr56DUZL1XEHYF0GVr0Clq5sAJeVK1LJfTO4igH9
kuiXo2X99Iv2hOcqOsVJnefkgmst3/KIXHzxAaIiqEwQJnubIgBnOV+qYmVfyG+A
`protect END_PROTECTED
