`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOo5mz9/ImxVHEjqSuoOa0fiI6ak7M+rWt92ECrtap6s
ALLS9N5BC6uT4Nfx42kyp+aRva8b2W6il2CouYN3KnGxgp103dVDCmeG7k5zz3o9
LfY3BhHXKr1DO7/oUbfPUidcrjbWhl5+yge/C5lKk1ntwbTd65hdiW/4Zrc3LBQZ
vi7VkLk2pw0nxjP9pl/lTZndQytDfx/C/V7Q+G3+XQ15EUehhpiyZkiHo6zIeNpf
9nBI8Q7GcFKwbVbrOVQSi4Lzy9MG7VMkxhXmwWOnsvsm0BYfstjRSRwQhszI9Db5
lR2MqOuIp/X6nZ14OmietnwLbjQAPVoYa9tw6fY22x60UHBuk1QqVDoXhmSsrXxZ
tCkUGeNcc+jp3uJRQuKVDejDRxLlYg7BTFy/szmB4WSCSsJQ1MaBYAgOQOUKuo/A
VJL2UP+fZ1dUXFRrNXrErnFI6dwHFCkW07q0Wnfs2B5Odh478pZsyGfVwNh3Ruzi
wWgYlfxGPNU5KBm0jrkzE5S2b+8a/ITvUYuzn5H7LO3Dz6hbL/FgYHLYgya+cV6z
flRVGaQnLIaeSg/abZtKdGtpGa7IQ+hMF97xlTvlG/GU3HlvfsX2cOdJVSvpBsvI
Ffot24tyR201HHHwyfNZ25yuQHoJ5por6WmITxqwyf8qqqmRbNNhO5FeuPvCp8qo
TOEAiM5a3J6wrqgcP+0JINklY0v2LwFhv0atoYCZQkXmAaOg4OqxqCES2DPrzLS6
u+EF++R9fCt9F41TO912I3gAperNDNrygGx3tVb5lFyi01IOgt1B4hhzH5F6Pmtc
SScO3lF+I+HMdbu/36Mv8mIS4RAEmBM0Ww3xCVpqH7U=
`protect END_PROTECTED
