`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDcT3DX5rPUybFKSgn9TKA6dOsnc+BLG/GXvxzh66f/Q
xrIRhRl8/aGPXvFbct+r0sIfnJQZXfr7Y5eO1TWYMRTQ0uvDFPiSfQECuQWXhwEf
ajsoQUZjfwaR9NZCqPAXD0STtLEcdeD8sJt2Mya8ubdxxfLUbqE/xb2QggP74emT
9BHNCA2llsmQQGN4Z7gv8DFUqJgPsmakrfeN52C1lXnJ7IrQCiap5L0gYQNZWYG6
aEnRUHgoUa5fokWEIFtXpGNr5n5To2+2IHbeBdeENNy6lA6E18oAgkudR6xz/OkG
8VSqpwuBDZpkT9/tWHgehg==
`protect END_PROTECTED
