`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOeVQcPdAv37pLqCp77hhtzt/uVJaMq5dQnWVliJLWoS
nWoDXDIHjAke194gbGsCzYpLzbLPMXUlcFTDLyf/BJWzp1eVFh7ALImkRkaBxsOa
vRbXle42vSUYXKotatsjKlNIoAw8eYmztHl9PfMzEBzHbXyBDTuKdmcASNFiyT/g
EfC+8HIDrne5zMMhmjjcwBAPwgYCj09lEGHtkTRp+OC5mY1L/GRsNPBdD/mOFlNu
1Gd9AdM2U9Y/rMyBiu+cWA==
`protect END_PROTECTED
