`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGLW/iNaNCItOA6YVGonbBexNP0c/w3RXVqTQAAwi5KQ
sy9qgEdk/IJNcBSqX3oRrkMYfOAlNUoTlOg9OTbMEAso5npwgRMdtsOkRQdjcXE8
5flpbN6ck5nRfbOcStpy3LM7yOqJSAe0YlgrW1jRTjQnk0TM34WMwzGlaZm6vJna
PvuSmuNM9eTXshVKutpExdFUu/qXO9bKWV7Skb9xwOTvTPgBmFoR3SVkxe9Ao82G
`protect END_PROTECTED
