`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI2tfouejwDNlou7k/167pwGOBmHpEixr+ocRRYURGf6
Rnb25aDa8lRGg5LYD/LhbMii1kTYFPq8P+2xcHk8w8if81s5f+sroGi/r9figYv+
d/WA9uJFzBU+LsM+4hhQ85squOLOVg0xtD6T1D5LZ9jb0NnafpsaQWfNp6FxRBuK
Jq2wyzH70ccALoBmHRHhag==
`protect END_PROTECTED
