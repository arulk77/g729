`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/szJ4N1IsR5NRJoTdU36rt2PgwfMZ3dywCCkBt3pF8y
YLQWvySDLThpA2/pT/LGFm7arMJTqvZwGZMnG1NLR3AcQlCSv4IhPPwfoU6azUiC
NzwXRPI2vN73OaG2TvoaGobjcIzVPCUHCzZl1bALW6ilx9OkT2DoyzaQickMGWa4
9KZmNQgtY5iPobJtviz1PAf6pPYs0leJd4Mh53KHVqQv9GbPPJ+HZ5ZRDupZ5AV7
kwg+axiN6M6DqytBrVRRbgZOKWYb+R5UAV+ioz9nRNCUlgig24mleKWVh7AeLHOT
ocllRQZBiT/ur7R4zfV9GA==
`protect END_PROTECTED
