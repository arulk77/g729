`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePhvrPmILYk68llE6GKqRSjsPHeoGzJotqUhvf/yoXHn
lkABliE0qaftoXzNpmdJ0prXIFt5Glqs1kndNKENa0e8DeuEFE+m1vkJrKzX7/YH
870i0mbt85Z60bkgSsEoXwE00C0qxjISMHsm79FuHybHXuFuSucIpplR6Q/I/E5u
UVKQD9EDeRm5aXhvZI4tUyKZSCOo95xaIpIF0fqfGS87sV+uV1PJL+vic6WHJ7uG
aF0gc03g1hdiffXsH9/NltzVQHKOoIT9kRpQBB+txprTMmb8s3184rT+pLoHj+zt
5KVFaz5cYpuilSF0YAJzCkjCTJ409i4OfRaDbpjrp11r1llYx5Z8wK+0UC5OcXU0
vIsbFnKhu1jgaFUXXdZxtRK4S2e0fE2R1z1a3YWIGyGu3QN6FxjO/RR6Mp9CwRAL
c/PcZZAfSrNbycsJhsVOA8zveXe8KPFwrM20A1AH9UTYS7KHzWAOzU0tZfUVaqqR
ZlnbsuWSW/3d077s0Rqyx0BnkYPoiHUJOyWtxc1WKZ3c5eEij/EVBGmg1SZYLM7z
`protect END_PROTECTED
