`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGAz8sYortK6VGbXa0AspGbDvZLBhXq7mVAjbdLOnS2l
bGqCgM6E2YlGJsHEYruJvU/IFSzooGgt1oX8NBf8ZrJ0JHKMnSlMhQW6jk1R7DYx
M8of+6LRIgpmxNTP3xsRUVwlWJARWjUYTd+/6Kmm5/TjW9dTAmtJGB+B1n665r79
Uyrec2KKY0YCo4TDa7qBDj29eCttt1wTHIZ5J1ku2/dF6QuXmjggK42+mYSTxm6w
B+EIKUSBApNXFAWoJ+AkOroaT3oGgF59ijBEkD5tD25FyF9DdwKIH+I4pyQ3PgV3
B+JkPbdaeyqiSoSDT1pughV9arbSlzDj9iU9HO+tw4EON7nw0Ur7mS2AWa07oVBz
Cju9JAtH9eX0hRqgrIaHqfsWwEFSaFIx8Qes/g1wOTcgdUJwFR/Se5Hu26+20ytf
EF564M5J/ZVY8nRo98seaV6mKvB7yuMOPNXk/EGtIj2NtTK4XieklyESIrrqU546
SPm98/I9+u7zcWlOIX42yg==
`protect END_PROTECTED
