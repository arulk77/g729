`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDCotbgp1zt45dqjlOhkDX/kugmh81xYz6Y9PIsHY0um
9P0CwNaUrgeSspXhAU9xRPfSldYrPhuNznSGBv9GWCBiWDFxf8sBjWGmKjqQKv17
Z7GJ0Ens95GGAb7LaGrUZv5LL/QqeGSEhlaXKrDCFxeyULgEnlQ9YA7tXxiR/h+e
Y5k2oczxYKzCysV7/zh3fbOLSIc5fT0XiZMUcBSGz9yBho62FRu8G44sKrwPfJjW
`protect END_PROTECTED
