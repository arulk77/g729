`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C0yqBkyxZ3P/FBnPrabAfUqHUoChZzWDmYNvBmzAcybI
zXKJfS0msgBMmPWdZ3bG/a7KYDVaEb/iGb9MQxRRjuF7MXuQXoWIqAZYPEj8lAyo
hU+vG+x5zyepjx/3T//JTxdaeNOLJ3qEtW9iagFk5/J+qL7RsD+u0WsFPyEIH7GS
Vd/TUHuvAQ81kOfASQP3rup+cGZExlbf+GzV4QYwWcoWXDGZ42Ot5ADyt+yx9oPI
y3Bq7mpIFdLsxCSq7Sm7VyiuYAYcUCCrXRSKvJz9nJcGu/6EyDcSUmcB38XCXwCT
Frl15iulr5zJud1TI3F157s52rpnOBNwBJQ16/LaeXJUhLkqATA1HOwp9v79WvdB
GlBWaxmg51L8uGspxFXUhwzL0JxUs/zvleGytQqqjH8cej7Z74Lbe/3QOeb+cLMl
Fo/M6LW766JCmKYcIM5sKjPsysVcqvsbK3hQn9PmMhzhqkwg/FekwUyqF+LG39aq
qvMZTzdPxJX5zfNziUxBF0F5DRFBmOcoyfyv6JwsTp4nD+7O7lZO7mGxOBhjVafS
4jHm9IWyTrpqaPQAsXZ2ZS+2an1traUhq1UVDWgNvvN4+/1qtnwRYB19qPYIFc36
2z8i5981EdoBJOsdUMMWJGIatdLR9057Ubq19uItoLMBqYUOvYRdgNae58lxbm1S
c7lrBvAbE7tjr87OgKw10DrzxMHgRFwGcoOInVFp3Vn/IE9w5yoQJRNgCUXDJLKx
NeUg4ZNCTetFeRvVXdFXEmEplVDZC2NwiddQsB+CCdAIjZlsZj5Y4Gs3BSU1R2ro
h7x01EIuN0CwLQbVxboKmzg7oCnU/SxHOi6aTN2de6rPDVdbQe++U/t5VItSXO/C
XTr1ZV2cA4YMO6EU32xILhBIpp9ZXfOokunJdOUosnPo/3yTo4uiTqvimq2F4/i1
yGum4vSsxi0tOs0j6sCetIcT5zJ3WJx95ESBwXJkJRU8bEMqG961F0QKlVsoiXEg
IaHwfN6wS/vyDbldFm0PdcQGVfU/Yfajkg1rxqo0xottfDDOW9rWZmkAQHywxBuX
`protect END_PROTECTED
