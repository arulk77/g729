`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveP4rnmfyq7xm8RZhoSvsS6jvLe3FeRguiPqJVnx/bcq7
Ocfqq4l25JzRMzwTGgQKn0Q/BC9V0U7PlRT5rpQ6Nb3ZxdFqxoqrGxF0P3kqlK5q
/b1E3Jy88ymKBatt7cDUEPnEMUbn3qq47QGUsMwHpblqhejsGdrpd8Z8cXsSfkLC
hXZtxIe65uc+2zI5HJwMdh9TCUQFD8p6x6PvO1CtOAEKXW/Gh3BzxvuheRqDk7Lx
`protect END_PROTECTED
