`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB5gPdvZKnUGCsS6E7b5q423PaCel0K8XcWjeigHfcVC
8cATXAg1daTlNIHJjZRqEA5h2vfn90zmtEJgRMzrRZefxFrj/uvhyhMwNniDnIl8
v8Ko5lB1sSgZ/z6ni2PaREhCzyDDkZtmrQdmKDU3HuX8oIk3y1o2kMXUvuiht5/0
uoUkq5DN+FJPY8vtU2JH/arv+WLHQI8Jqt0CMYj71qy1xWcdfTa/tFPNoNKGWIL5
7l/+IFc/hTf1duh1rrtd/WW4snayAsOUqoUG/2dRMyiEW/VkZp2cHIrZZXXntw0c
0GsH4FP6dgYwsNeRSgVDv6iAaPdVlbjW+siwXbES8o+ZEXvJRjGWDbYgbpxtKLPJ
+yq2QGZn5jScVk4odvVAFlSDJrmxfW5t0lE9WihAyndISRA3RvhEeYtTSpW+YgGb
MKyV8WT6hVtQsmAwTFvOTT1JMuIP8Ma/pAc9GweHmdmdE4b7U0EMixjA2XVMei/+
GPo9JI3dGviSQlF7FRvzHVLZx27ujubpQAhzvViCkRmw99xz9VbZpNMfbKg/1+to
`protect END_PROTECTED
