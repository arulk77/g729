`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
SP6HW5ECyki8uHQQTHTJAY37PpRwfPxApY1RCkgd5wFvt44H8TsYSr9gS6FfoWH8
h7pYOYKODQk4RiG6g/ZSlStjlAeU6mB0psN9pRp3B8d++kCJenrub4Ts+Gtq6ytO
6UDJBvPAVf7Nf6FxAh2aVY2CAjiOEtq4hiEBXIKILJAWAAOJBDUn75rrzCjp4CIo
pqdVY4rHbOMGKEPeFq1wtPU96CyKGtmJPWx68NtWfvaH5sncoebwxRvmalBj5+iN
dW5RbHNqSPzObKMbw4VJsXTwxXZOXCvLae/rqjMFru0Att9fNtkDxEoxtXdtHaKb
io4ksEqpmbiuUKZZ2s2rPG9eWWtsjZxdVaxfXEsYmr/E9ZYwhU7Z/M+ZjuFTQTZi
evJsYJZxDgeNKz0GJCAniB2ds9Tn51QHZZK5uGcbUzm2dgsmIeapw3L4XoX1cQQ5
TWOy+HWVAKlRj/y2tgN2UDY1QzDF/CAXaQXL7gx0f8EQ2Zeo5g9akgGtOJ7FEokW
7ncgr9WSZ4LydNox9AHgxhFDUYRZuNsOkKAh5u/EW/skiXDrCUUqb6B2yxZXCPwu
9mlmUM5mjBuNj/65JaZLr0Np2DwS7QXEvxv+i0uvRv++uZOsoXUasd11hDXQtp3f
k9KqxHghvGCPFdTYljy9sQ==
`protect END_PROTECTED
