`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QNw40IqJrFvY2E8HYWz+j574SOYd175r/uw+W3JPo08eqV+AyQ7Q1BJTEYp420GQ
dKbfLjPmw/YitI7LIw8lcNuZvoL3lU6L/4d/A7juODanHSpTrTBG1QsUbtq9cgpG
uhhCpIkcPJCZg//rCuneJZBXbOy9P/Oe+oCzrFYin6HMDbg1bx9cpzrx29HsZtXc
`protect END_PROTECTED
