`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
xrY878RsuaKzXoiw1gkOuHv8sNOyowrigGBLKaLYtQoEIVi26rkX6CvaIjmuGHcc
6jfeonzhHdPzoCZu/G0SJX1CyuMFL17Ozc3p7Tns7X3MQLPMqAut1d8zrSheTDSB
C44QC3eh1UgDYo+Z+tmV9So+3MoEtoXQNQ4pnkKehBhyceZHNESjURtUMo12ChbG
`protect END_PROTECTED
