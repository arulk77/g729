`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN1nnV9iLnzbwx1RHomM4I/4wjJWWL6A+MOThXAs2VtJy
k6J0P1YiKkFysxO/aotrIuE/Fcvqep/aFXCqcrAh5Q2WrMNjHn0AHpd5Nhvj+np2
97KcizMcNtKzVRpN6d8k5pMaXrL+2K+hwuPFxnV657Gpk6lQS4ebO62Ql5wNU7lp
OxKN2EcWmzl04j23N7KQTup7/karFe6aEHVP6SykpYn0sq71jZXujXob6zPKN+dW
qKrmCVGvqgwVVPoXxunRXjZOvCSfAg5ch4Cm65+7GOHpEscZMplJohY1G2FkEXpk
LxJqe5m9XSAcGFFFiVEpJcN08ottQXmBl39KJfzJygJJRnTiC3uL8kUzhxZ7EYpG
YaEXvS6oUI4EYp3wahRk42nQCXlgn6oe2caW+CX4WIwRzpBxJTXQOMb5J/VFi4Mb
YznaDRFfv2KhVVNYErkCQ+P7h+4vmIBssKQezicbkeDugIBXX9XeP22oLdjt8DyJ
0meHQOvYh7OKqUlAkRESZOfYt0SkNhlh9OLWD9AuOMzlr5yhf76a1T0QGsfPlPRA
w2zshviDunVy2jsedp1v8ptcXA6E2322PLsSx6ZWEiNcqJQ0x3DuubKoOEIN3m/E
/+wMVU90OqGJ3PJqGqnNScfK4k82zLtpQwTe4QwrKA6nQaGrm+A4T2raC+OzISTF
6792QzpDTC0z1QG59mb8D/30PbLl1gQ7zgo8ALxxj8X3QFmtkyBg5UIdreFprF1Y
eNJPSJrecdTS5xjrrfXEqDaX8I9XXA+ZQ/t/GsIGPzeAn8yjG0aH4VRfa4koSOKV
RAZbrqNhMmCssyy598rHVg==
`protect END_PROTECTED
