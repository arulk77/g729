`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEuriKZ/KxNxjuXV5eS/ydr5I3hx6CMZTn3x62Oz/krV
L9SjDv6nAK07W75dOTde395VyfdZvochrD9RkspptsDGQAeEKl+sfU9f4e05iILS
ylTM5Zs48AplefdJtc76KiGyd3zI8CQu5e7Uymsk/UYZ0ikEKrdtKDqDKcqLyAzo
1z8SAuVtg9elLQeM1KravWy42vvibVyywrjcBvr1ahtXnUuLEfGgVr8IE5+JYC0N
vt65++XNJmQd1F143oZCmM90rM+Kc0d7mrMpWQOY4dvX9Knel+VAie5PZKKOVbOB
19bV0OcObMWczw9Fq7xoT88koE9uSrfvFlQvnjWwoUdbv3ozLB6UK6x70vC7TfM1
LYeOo4yjs3T1O9VbTnHk3O2xyJNHNaUtkWeWDmy+Ki9XnWKEVHEdBa2+kcxtazKH
M2Jyp3kTUKgBF/rgr9IpxpPceimCy7mBaPcChGbNQ8hewBs9kzAN8lsZsE0SNRnF
2kkwytYR7nuWrlAUF6uwSPSrbwEsNSplFOjAGIg0InxM0oXD751K0OXZEup4MJb8
UgwGT6o3KX2Jl4rNrDMsCjQGGZamVGsRkasYLuMhE1AEr9AjgIkWXeuK/p7vKFIy
iYooOqHWrvj42OmfSVpDWBUvhfez6bkYE6dU2kNJ6qfwFIiDr2OKxv2M+BWPKaHr
PFo5kEhHw7/kU+8LZ5iq6hdStMRxMRZSrHX316W3u5upokMkcCByMItaYBcGP+ML
g70YGB/uRaY2uq0Mk3wjkojxihTgIsDChXnUCmL0Vpdj12/i0dpzRC/8M/v5PiUh
e5/Avd3U7EfzTFiAaPrrdyFD7uneHVaFvqJyBsQ6P3/G9q7JQZm6orAqTWshpqW4
2yj0Go9nkBhxC6bNuk0g8UX3g1AatmZkSmQsESzRxXTUKCBFJujCL6EukxZd+nk/
mdbXZQ34tWXJNe7ZuNtiiL2KOU42OlCIKWWJpFrhi8ByVHOHcepZqLcKqs5HTVkQ
cLG/ogl7cOXTHyjMCMZedMRhUeFzKduj5zeiVGKved+CyrSKqBQhaYj/FjgAy7sy
mO52EMaurd0GfPf2/FPcte6X03LcDIbZiJ7ROKZtl4/DyOPhBLQht13WcK7e+Ouf
Z/PGniA1vx2JZ9X74tXIsfIkP3D1U+J6U69bSf6CZc56Hnykl5W9OsAHKyTCXI0E
dbS5aX+D1FBlanS79q6UfTvcrb9mIdRffE6OkzjhzkoZgmdPxCCBBV6Rfyi/fsCR
`protect END_PROTECTED
