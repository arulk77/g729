`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCh1oabjms0vfqwhS1h/Q5AEczStbUD0n/1fY/Y7oPLN
Ub9W1saTwJ2figdxB7OHPL8xxySoY/HM2/4VIc7AVxANO0EEzbWjJ08o7VJiIBoB
MozcBqvruSkoj/dv0KWW/WjHDYVfqQjBE4t57ucga8JW2prP6XwEl5jbJam+LPBa
2nRM0kDOWXfbFzp4VaHlQ4jOijddk5RGnKl9F2S6hq1KDGh7SwOTv8qR4ZOk7ZLR
`protect END_PROTECTED
