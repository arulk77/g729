`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
6SaGx9yYazhJJDx5eC5o5VABEngqQdtg+JJQ4aPayRmVAb9kT8WhB0uB+uxtmqyA
v63Zy8cRnDsrsUqd1zhEkzgh5TDNWo6eEYC5oN5bQdHjK/1EQ9D1TApyESDum3D7
s3cwq4gFutxY3ZvGc7x+dIWnQ3EuMc/SsrV5dpHWf5Sq5NaodDk1/RiIyuQqTG4Z
HuUruQaNA6ZIhleGs5ZwyxJqpj8BisBN+JNs8Kyox1BLhGCkTEcrXOtkaM1mrnyu
TmZyFBVFC/r5/cj4ZujHFGCpDs8ckhPcnErAXTS5xzuQh9YlnOAf4TMVPVpSzbfM
NlQ4wrogyTheyz66sskWqlHDwj8lpRBJaH43NcYTLvd/AW9839dNyOJTtFa3lBp9
7vDNGbP68/K4fhvc+t1Lws4wBeOsXwAy+aBhbfSQJxmIyiO+OZHgZdOsImRyTFtl
sp//YCnsYctv9AM0gUAZGgml9C24PNoqF3q5IMncCEmptVCOe1rsNTq9M+OQiS15
XRPGrBcFp5IKvGQLYVMEQhUOV+aSgp1F7Yl2tq+gzQq/DzzSmzBrtJ3qlIhVWDWt
l8CgrfAc2Wzm2knSAuoOrGFS1qu+CCCH/jhKRncqS84NCdpYVH23diPhM71mMbdg
Zkmw2eUrQ1uKI3g/uySULGouUsdpV2UTSd5akuzEbirzgup5csY4zWr++AR00T87
KMIZ3Q7bINvkX6jZVS0sWIBP1eNH98Ds0z1ZxmSXhVHXejEI+MeP971UeCiFpYZX
vq8j7X+fmXRSBns+KYY1bDHbAqaQV2hvAoKKG8mjORttmzIt7OmiSbm3AHz6cp2O
Cp9aKQVGXq6pp+qkPYq+8+Esn021Cq8W1Gx1IgjulqJiVbYr/4qmFwIwqYEcEBiJ
2Gea5YV76UhTAxnzY7efyykJa3ufXInT6ZDikvuuSBBvPztuhaCXClbQT1gINt9u
pdi8sDy66fAMDtP0F0M9qzrizISRkvSbcUCNg2xfW65e5feSygRXNNlqf24ChWFp
PLbaiVfDn01OC2cjou0P/7S23psHT3NxwkaIKyWwMwXrWGvzONQb9QZUpB4lvXVN
DjAGd3UY9ZMC6AFL1297dveEZ6uH7wi8a2V7AyensDpRNqWK6B+LgGCEwszF7EkZ
xHlySWG9xwbakm+xvQhgChH4vo70X/9gnD6O+8Cc84nnOqcnMZgOiIdTuNum8YZu
dl63VnYV6gClODwWz29H8w8w2WUvTjdrgMdc+lmvEHxzJaRbQYEEHsHQ3KN7T6Ks
iFIeXch875PXjTgQCVeWrCSSXnJZwlnOveYGklO/PdfUXhLmnvaBCAb1g8TMPaO+
4aRVxrThttCBXiD4LW5AJj8hcP2bwFByGD7oyIhCedm6Zz8JCigKoe18O2RwGeEI
H6S/I+QPHV1pjTMA3PU9ya3SLfVNOtD66VL6OT0eeHL3QM1Zg/7Tf6Azd+FPxVPv
`protect END_PROTECTED
