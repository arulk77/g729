`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL8ysILdeuCOmoXcTPltE8VCauH0cnT7VQWxrPBzKg41zR
XLpQM2Q8pIJo0aU2uR8F4E46Id/MnXMId8Vn4TrM3VyfmHVAIcifgUZJeZVnO45L
+npTn3QXOekttHbj+7KtDZJXl0fqhGDjwEIJ5azbgnfYkTWsF32eQy9eVKYEkhps
kCoHqtSxrKyjOy5vuU2t3QSA869r2WsCr1sseUGrrCkYQY6fngG1UhnLs6MJf10L
/SMBnUQfTW5EJ7D69QesBRUzB8yN9mR7ShLu/MeSMtSPr3LUA2ZjiHuTkr7GUVrE
9aPBNbyDP7CRFqT5X/H3wARUhH8zQCJJ9/rFg0fqT2sRdlWV/imMHHGPX7OhYb0A
qakKNmjn01ADuZXFwCdKpaBxgYcW74a0xbY3nMBjvNnpNUQz+yABl8JjmYfTgWj5
GoSDixIv7tJ+dVIVJ/iii7gehcGMaSZsH+GAJU1DBM4aBZ0OnSYP3x4k7F60YF1t
HxOa1WO/D4Zs+4JlkG1BY7hqsymhjUN5sOJvCXf2aG7SLkNLCA9mKhU8IwbZ/Tu/
gXCGqI4QUqQ2yA+WUHwo9TmJZPbsBOrRQMV8m/2T5X74jQWdaR6iI9w0WYkcLsfk
z47QoIQsqlZOhY0mIjc6sF5xcN3Bwtxp9iBAVjR2/5APglITtFP3qpc1e8OxPV89
L1YiXKyjAlUJVEYos18+ryAJ1pXao8iBhsi3IoaaG1A1GKNzq5vn6SlZr0/qnMet
mqJCtlFTV3SB4aO0z80lCM2LQw9eNdwzJIdyEALBCAvrt01SmOlbwjHa6m7Yapcp
j1EQkr1xCRWxZshprUSTJ9Fdm0KPdTzgaTbZd103hWvZrNPvNRhffOHevTukBSs2
aliZ82m7XtqT8ECfR3CJAyzf67nSHVAb1HAeiKM4vzqzyiPQTZj1+jME4sXc6jCg
plc83CSCxbnZT2apgl6zKS+P1qSaq3ILjPK9qSdPHsPhSGNIku0YL8s6X5RwsvfJ
CorOsgbv6d5GqYWvBkaiAmVLM/EamRO4QNeiVvdH9N5aclqkycNltVPiBOXg732A
KX18pzOc1PJVhYtmk8qkopjIlMG2uJtCWpePyEbN3mR6rTVj2Esex1z8Ep15EaMh
c3qI3vkWLtEiLtawoJq2ruKXNIPXwZZ/DNfCsL4Pmf2xOug33XGH4YpH/4zjpxCv
izNRhQHzCQrz6M5H7ZpWO56lgVAEcxYiIwK78vzELUH8QAhtqxbeCIZfvkFuDUFc
99Xh/3yFd7VGHNmh0zcZbCbu1liVpIp+3lCXiJlaH8P9TeYdZbG/IpMKwFaNjuYd
XgTRC4U32uwt70ySDBtWAAmBzxmpYGiAnTkeqaFS5ftp2n6PJmcN88xrWv54hqJa
Y8xYXdTFzXKpD3jdo/Hy0bVZpZQXI5PoAePF9JO2iXhk6xobKzUHfGgC5R6Kodlq
zYQzxsrdnD2wh4MMl5/6eb7/E046Ok7q3NDRxnNycG9tDUS6HF6LC/4A9bDcySyi
/xLtYEht+34VIRIh0UU43PCmJIlaKFdrXtM4XZJDR1FPwXVZAlUFEFWM7onO7l5C
HOaCiSCx+f5qf93r4DVgQI3xc/pGhRIQ0XCiUV4/PLO0BkQnaF2mASCaSxjoGZoT
+TsmKMxXi+BMoGrCI2hE5buwZaPgLML6lAnYhQChW3zaxhT0Htti6NWXX4ZJbCff
sgdzah2ve9nQ3dzkcCvjeg44RJHmyoMsZt4P7vL/tErrw4gbfVVSTrfxfxX7jcH8
y1GdyaXFjxFeOPpCPzsq52oJf14xfp3Nb0lmKN16aUT2fZOALSd/IhmEIdlYSwYt
gfdlhC/69tdj3p7HYamCZcIQC5lvDbfTwVPCJB41SXwdYdyUQEHXLbQFzU0cn2OI
XPcbGHmeL7/uMQNNjmsZoKAA2nsIM9X2Lrn0ekTTohbZK92pOJbSo+I4kb0dWV+R
DhFhs4oAuga/zNEFjyygnChEkb7U682/kcVy657ijUNweqf995paKNDsIj38UREy
/LwRWj+vw1XAw6/NTgirXS4B1bj5e+GW1OVc8/KpqvGSv3ZnuDvnBxLZsbaVFBx6
+sWdfntPa96KZ0rFX0zrJFVuk61bdtD8RlgkGgXSS+KKy4LyY+jV0o0SEYNhgeyW
9Yfir51XaB4PLdZhcGrzG0MUZu5d241aGMZn6JduC0jh6l09KxzGJFnZfUMOFUOV
CCDAEeQdDbYsnl8XCrUo4PPO4wj5feTLTPuHDad8/U49KIfgmQ4pqXAYWRpI9Ev7
7qqSJLp/VOlO6XV8epaV0RVhKmoAXhXVuL8G5n7E25XcePv6nOFCbbSMXrKP4dV5
PrOcYL3Xogx2rWe2q0lyd6S6w9GiQaW8biCtyrQkBRe5816ObuKmz52QDPgh/ZnO
O6Rbu9fY0iEt4sePtdgpMIqRCMqzs8a0SGXVVbsu69C9sgrQ+mIX9un0HcYtNOJQ
Aauvm//DBaetsoqtqTcKg2rwboRFGo9L2agKjJTz2rrsGWYRFnaiRjs/M9TI4Yhz
Bnam5Nah0PGbWcdAcu6DgtDXw8viLyQ2QRZghoMxfbVedcaWPplDoeI2VQe5mFU3
0XP15QNa+Ee266XPp6fHAO901VxK60NSovg16uAP/9hPoABz0LAX7Tl++PvrdWOo
rWcORbYSIbs6Ar+kLT/nZRwBYxY2ACj43XV+eQyvfa7Y+uOcnNgXwnzUW8luCLWo
StPym0iSw9w91LQj+x1K5ntJxNtmlIRhtrF1UXyzTN7dXXR7mDeYvMXfEoSOJDTt
4HiEnIPYowx8n/aCCohVuYC8sn3pDNQlk/i1ix6kOpSFZ5+6zx/MFc9mPJa2JcYa
vIQ+9zsJJCz5IUvYytM/wo6wKJxqtWcEONCGGxCLf29HjbG7H9tVIHUt31eR9x1u
Gm8NRqoa7ZO5d2fGkV+13pD9liMvPuwoIBkTAQr7Xf83lTbhGQbuqvJIUD0Wl4sC
aCkxpxVtMuxXxNy6weZQftk85uh7fNvY7kTo22OTtz5458qzVjP3ubWIodNAo+Gy
WS9A3jH63FRl/kMJw6zPl5BdoZ3i5NEX2nLRHM/kznGKDcxOb5Mnbc3aGhis0/ez
rb7C9YGSeMLjEgDEsWwaHAqtTf8M3rU29wRKUODKfbjM/VPy8u6JfUUZdjgTHLnN
W9paNZYVJVrll4KyT9nS1l6EzCyk35aFxhgJOWDJb7/OHVdXMwWpDu/mLHoTbeYM
Z4I+AAfm2Trh0BO3YglORruVW/RsNvWDnx0UUaY1lf6w3jyG1uFSox7VAR2d0OYL
rxb6TNQS+t2DIDSqEb4ZQubyjK7nUvMxvl3Pyu2/OWBfh6D52Qh9cddVh3f824bP
Tkg9SJg2N3QHaHCIpZ2E88vk4vR5vAkaATUYGJXwjjfdJMtcVVhlQ2ZnWSpuCtP5
WozeWEsnvp+MquBvK2yf68YLP1YC69CxBPE38jz4vZG6+oBw8P2GFhiiVhtl5WkO
mSH/s0Ah6Dml7fsYpaa0vrNqronF7q2898h4pYjIzJ15SOkrvkfhjeQAS3xLKH5S
vYW+ZfcKmq9jZ2qTIQS5+HFStq7qBrqXiqYPT9uz5aFjMV5k/YTX+dVyHI3OPPQ6
bRiX/xrcEAZrYRozxVpQ1Z8DmAdzjBDgaOc3USBBc8pRAauYsxYtqwVgYGC4NxHV
PEvBOkvSG6Owj7RyBI+PyEFcjhOG6YMIvcNHAfFOt6PataA/wXWurJp0BYg5ZaAT
PY2so3Jjii9f7AYlWED6kZ+aZL6Ijyz9AHxF8gQde8h9bP0u5PWrZpYwLi2WYY9Q
utbIYYyaKA/rFJB8JZnfbIxrud0ccIOG5mp2QQO5tU3Chl4T/3PRG2GYLb4fKL3V
1wT4DMAHh5GSaGZUFrAWD3ZJSIMZ0xGt3A79fWD4NcORWhwkHXgsXIjPsfbdzVjF
FfEqVx8ld0/k3tS6WqI40/4C66fFvITuz+tPQ6LJeu7NPfavB/FhtkLcg59lI0l+
qfOcn+r/hmOr/fgGIB3u1KLHkP8JRqiBW0y/CSYUKZ50NfwtvOQit8LeFPzACIHf
S5vc84ENmI3gyPotcZag1qQyuMz3BJHnGgra+XofaqUQzHM9iuWiD4uq8I/uex0g
C6X/rpeYG7EapTjs9nQPOfoadtYrMrifQtLNy5UbXJTPPs0WfjvvMPnpXWuc6UkA
hb2+9wakXp8Kq+pqaoOP/N0i1CEEOz1YjN/jrymYJcUrLxhnJ0IVvA4oWJzh92YT
v6/HeAbo3IlZJ6DXZUGWB5EvnTPyli4whcawPAal33oM2btLgQqlAI2SaezBz0fW
cLFQrGyUJtDf1ZraPiUuyYDWiclvLAgN8cOFMS++nlaNgcJfYv5qYSjO1LXfrB2U
vjDx+RLJ0vSauewflmTe84tgyh3DRa4qrnBr0yBIjasfhxFK1KaKSod+9Sl+CjTL
VsZbWVWcMe2vAevV2pWs2LPx8eUqQF18yULYAHwQvVJ4ciWVlTxxVOjGUXiLIfxK
L7AxiLCyF6N9HAQaQ8sSb5DW+nDVVuHGYnYqzlZa1P0DAxXANQw8agNs1J1GC4ox
MIFG3ZSFc0OeCYe3n0/PlwlWdB4k6mbbG73ClnpINItSq04D3U0YlsJEGi+G2amJ
2/gw+rvbcG3IXLLD2PpN/MvvJoDHqZljYZUMsdnv0i4aTUU6orHc4+wfgn6TucuK
2kIUaOiTxwOMVCZ5eGzd4MFOPjt6mltCG20dCoxiM0LO16NqEUVlmnJxn9eI9BYD
x+hcr0zj80Z7/RTSL4ILOtlCdjprw4P8DCLiEoUzOv28PlVzit0rMIbm+xl2Zm1t
jCJ9dM3DIh5l3puJaVoxA3DBj6ZxR1KDU811kt+SX9RWfAPp7fAcM9sqcAN4LFqT
MBHT73yOaw1G9OHCuZi/cT6LhkehRHGHLT/tLOfeBil3SPeC85oU3vCDqCwAz8DT
C/FtegOepVSl3MzjRaP0jppInxj9LhO+9kFABEysVMKa35keqJiR3Pz2iSDhPHBN
`protect END_PROTECTED
