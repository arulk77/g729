`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIp8s+aMnDDO4u0tZwiFCxfd8ThBb6MQwthIpmmfk3cF
D64MSXUBxZNmd3lHzDpjxKZEJ2wcAMB2u2Ak4qcM+mtYS3Z56kOhjnLnpi+BKo4X
crML+V0CeYs1pWylpWE04CgaFRA8eOFMeBGwxf0I3Uqnwu2udezQruopqXD3HSj/
ERAtrh9hgNpC22wZO4q2YQqvLkgPX/ICNSqHKYzHy4P9+ao/DibiQyArtaj/flJP
`protect END_PROTECTED
