`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJSTou6jp9wmazSg3PysIsYVQmdGljYgsL6HIAEkbsFB
n0/edwvw4rVU5Sboy7kEkjkXotxG3sZoIpY5OwF1LCb9+EV4nqne0EazC9Z7pVdC
7QzJO8vknJewjE3enTWa084YECjtj0qNLcBZeBtEHiFNHpk310H7WH3g4HJXR+qk
AqI7UR3SNXKUiAbWiSB534JCjRrjV1HNW9X1vOzz3v3J8XjrRrtLITJ8g19UQ1zi
Qb9G30gD0fSNdlGYbNNLvw==
`protect END_PROTECTED
