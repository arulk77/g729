`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN4RHHKl+w8AtlKC8uVorLPZ9kMCpoF7o/XHQ5dIXAS/z
pxqvhAezB+U3mlyKKJXCRJzh0YdVz1fIgNJVMU03z3bSpi4nHG8BlYYWzrC4GNlw
u82jH+uGEZSBESpgfvsaGVcTN/6KTiN+kohoKH2rk4+GSy4zqF6EafBBRp5z2nKO
4/1sgrKknwDHQYzRezXNX1Tdoy49E0pjJBA3KjEROf7eLHq+g9NGptFXrHS/7ZCw
ZpPHOuSYaNkFbau+Fdo3UA49pKp+8kPCiGJdGW7P5gFb7RQZvLpEVwU/Baxxmdpi
DmlGQCHY7w7aZFK15njIiACiYutM42TAdzP4c9dVbUmxsp6pDygzzr7eGydw8jjY
/LRPNMEKGwYQs9IsH5RIwPo+xQK2wZJOVPnxOHbNWQStxcHRxSlcexVGfyyfgf27
5j8CusaAN1RmQw7O8olbhxs539gzdjFVgTf0G9fSbjvU0qh3osneP1x6mYmI3tBZ
eDPfleFN8fc4t8abWrcaOUK7OUrpa39KCg7EYQiW7C7NW9/HMog770xiLRuYXLTR
xQCNOasKBuDyz/1/HxKkA8b0zoeHGce4bys3dYfwPhesvW1Kao0CZVK27GZASpyB
8b6shdJmAoSXuNmePxTsnbV51ji5xiEcYe1evT39mAMgjHHLh2a8XUIdOWCkjmNe
444KnX1nOcSWNwg1bUJL2xzx9WcNov04WwFL5ArL2jRiZHjbtRucrZAFQU+o/hQH
VRhxYu++Nwd11U/wtxEdnuBHqoup3XWDFtIOdtZHpMNgohL70UPytnAO14wzHOTf
nJxnIaePPqavcrFpS8xv5z7AOIiVVYfxZoHgOFpwuqNVaZxCfHQ6I5k32MTrlwx7
RrzDid6MMAckdrKl+N4uWzOVe57tGdHZ24Ey/oQn2CcetBxVB9u+r2y8fPiHtHF+
UosECLgv3a3KI4CJUhpXrIGLe8uyBWIgf/zvnm3XRF3vSs+iMQ8Ql64Ov+FZyZs2
mrr3bncq2qFNY0Bpm3/4zDL7CY2oX+iF+gnQPUMfIOuEAIFiTqdz8/zIbRGYq/mZ
IijigKWhvwHQ62JA5fHzKuOLDyKgm65p++E+Ykt1Q6d1W9QxwkBxPHGMbGdyPOwx
J30ec/K/ssHgSjqCkLrj5k6OvosejhleyPWQOU5EMPpRJ/3iE4TKPS0zEqSRh4TA
azozSKDobYThOWPnrlcLgvMbCVjFptKcPaM52zwnVlhHY9HdxOB5z1u9kyTPL8I6
npjnnd2C/plNawnNHvWbjwqCPb6O0kAWJMALMkjgw0dNGIehriGgXxETO/AlObKd
Xa+S2TFMhnSKtycxxBqLSsdQoL6utDvcJUzNeA8kbSw0JwEW5PVtynsqn9ssWj/A
FWDq9rDzWLgVT5bKjzJ1lZXSLnw1PmFcX4vvoh2WAljkweECG56lDNeiEvwAXruy
`protect END_PROTECTED
