`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD4kNyAY2kAsCVx+Zy35HtkITXNKVRehkp97NvJOAz+L
KyGPmgPWuDJuYmcy4jk7+49uKRy53PoCIb12+7Sebfj+2ehQzRDoitPCzaqdN1Ld
l1DP4otPydcXbJD0Qq2aI+k5tdflrs4G1Q9iNPbjrjmKrBWROnXot0YoMIeBjF/7
2N2P+KKCQQb0LhNBKZaoQw==
`protect END_PROTECTED
