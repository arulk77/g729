`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMPi/+gQrDJWt0UQp+Dl0KN9uSZ/ysvusf84NohYRsSo
4ixZaAmkJkvhcZMLiFuL1xcjS1f/kP8yHSiXQM2ORs5pt1WUvvKOCxi82olBkn+v
TCmAWWt4e/A6UGsxoP+Tk3MNhOfG+DxNyA2osMotFRoJEtVxpbQsKsvzb0NG8ddR
e3f+985NqtI6nmo7nFerUuWjct0rSjxSNNMu0CDQiUl/ADMpqg/1fEcIN6vMQgyJ
`protect END_PROTECTED
