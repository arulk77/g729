`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46rzH/nCW3RmwANJ0PdpSuRM4Rr/6BYJvzhyOHlyjKBR
4wry0DwVRvKtAYsVOw1ppdAj0c8EQ5CJgbtv+mRl8MyMRedQ+1murHd1UBuyxeXI
69m1ilDcSn+emwuKCgMhlg/vvvq+t4bFSj9/RvzqDMv539tANbGeNLMLeXNN8HTB
RHefMH3Ru1v2WpYNnt/zwhevo/qcM36o2CwPjNTZ7QTfSDuxAULYGoGctDvM5nAe
kd0syDoH5dmRoKS1xCDPeMByEEkyOrPllLSbLomwAveZ6zC9NBlezfjWf35DM8vF
dnCkkn+7LDctUg7NQcaC4Je493uQh59vMJWX8eP1s1qyvweswEWP3i8sk1U4N0Tw
FhKCUNAOcRskgkZzxCn0wArxU0B7sxFxR9sky4U0K+N1ABKocrmKYtAOZUWmWNNx
ecOwOKeqYMI4msjvi/nkVT5G2ixuzLKELtiiqqaC5kkwygmzwqvVuKWR3qM0/sFI
`protect END_PROTECTED
