`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFcfW5kJ9Ems31/PwYhCMBHe5mn2juuGMusRVzQFPcUp
0c0ryga24xsWk3PqXMDNYhPcr3mJBSHJROwBpBVPlP3DXiEsKW7pOXgkFKFcNtI3
Hv4BPf462AOv+2pIRNIe5QJxZxLGhhShyl1VoxKTYFSNkuFzI2w0/5AnAP1tAssp
UYIin4AFuuT7xNESHGy29e8LDCPnLrTnKIUm6T/4jqdmfyUiEF8AZXJAUXKr1LKN
LJvYiNtuEXLYBH6yFTbxAXN9cSyoY706d3WiUHkeemNj2EyQWTvKFqIoP3uwtDAC
klVzSP/ffWw5Vwn72uZHLRyHPk2dfOd+pPExCQjGPyGp240fYzyQ0l1RpsmhyBgu
`protect END_PROTECTED
