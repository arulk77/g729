`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu478Q3u8d6fLPGeFM/acMdvlhEJ0/wyp1iRHaC+PD2/m/
H646ow74LycUXcukwIx4xQy0sOkCIQDaJ+6EIOiUvJuT5+rw5n7fDqOn4YU6KoNN
m1thm5Sda71227h4XhENGFZu0ZfWglGR5dwjjnASggDCdFN2a2enJXlG4cOgCKq7
SIF0on2vZrvrQ8lURw+WlnEJBDG4PDNOrHqivWIoSjq6oplRCN229UdQ8ns2prxj
zxMSfHbP4g9ikDAQDXX9XYmv4/BuNG/bUbhlsrOo7B33Tf7ADS1sPx0RaRfyGP4R
wsQtlTmA7tfMD3AVmmeaFWdbA4lzg5aWChittxMmKcu5J+nXN54f90JVhpr7ISA0
YOxprmEfbk8O1Jndzkqh0w==
`protect END_PROTECTED
