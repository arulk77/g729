`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL1g9bX17yK+1gPk1CQFAyEDDPdLDDICqUHH6jfPtZfU
mRaVj/ZH3xIOXYHxp2UlC2OuNhKB6pcD4lLeCFoq6btPgS0/rxuqaTAo9zUc/aaX
rS/BReNLyLTKnqm2xEMBHwfwVaWaFJv92F1WgBxsM9QdGg6zx5EBVar/VoSf25N5
cD3iXfu+vS7br1r2m3CeOZxjqA/REHpFimN2JDuHAPH4yLUXdhuxGUzKIdiGWCkL
AGV07bNmrkIzm7NxpBsVHc2C4L+56SRVthLcU+c9IM8yBb45+W+jQyJMWxr68ZLp
ZB1QPJq4UFKhgNuEDuL0MMitN7+3Tgwvn7tB9fAvhyTx9rVd+AVFbUdAzi44Hh2p
lHbZnqNEw98zq36Byc4foan0fWkSd2GYQ4GHYLoaAA9rfnUG40lTvjlxC0sOGy9i
pAkJH8l23H2WQbQTPCgnaRP9KotMzXeyAUPIlK2AWh8O78Nmpax7cIIvXUoLwTwD
ZRR0DIvBnnD9V7XUbe2mKIE0zu74eQhy+hu0uyC6/4sK2HBC06O/ouyrgCuF4n+d
`protect END_PROTECTED
