`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
/CL5Ham4RW/rLq4Ftcym4BPgSmX/BfBEiPBVPJGu18+aBzM/BdoqonEmRDvThTn3
aHaKi5bvkhrIaBXnDfy7iUu8hm7IqHS/Nes5RxQAWkZ579FAMU7Wx4Tyi0Dp5rMW
LPZIpNvSwix1jrVYrS2cZPwezr7xSHe4A//BPU3N1wl6eVGwxw8LruehWncYoTBw
YvLlEUjbtwppM7DEY0uhJCpAqD+BemBSS2M63JMJrWwteYYYZjac0Bi1v8DsF3gH
3Asz4HaR3gh025CmTzJCoMFr7KNXmeood+GQ0HA/q4jFZJoqPOhQw8iAf6bTSuyA
hn5vaN9n4cBqN9sLi67D1/a20e0F4eeh+MKirZedVzg=
`protect END_PROTECTED
