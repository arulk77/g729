`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
q7FxaxeA60ol/zvB6rAYLYK+yNAwXxPSBzEIomFkFuRkTe+8YiXaC9mq55QPo2tA
GgoqZkcK8GUCmvNXRqGsJAlrTPtzi54jvK+zkHhcKCatUGcOznBIuGyjoTDXOrbh
kpcqLDAHU/PMyaeSFMZtj9opq5rqlYmIpj7fk/jP1F6OxBIf++wy9wBQPtb32u3C
a6bs+Lr9EtMmvt6Wl5G39TUxKmum61ciW5RrsWL4GKxiHuZ+2W3MlrLLESvCQr4N
nIgpDWNmARKNyzlmUZtEGmAENCxP1hXjQE8W2wGre4WH0FDgeUx6nE5CL126u5+G
DpBPZy1RkkBw7LRolPQVz9I1vRDJythYJ/vNwhbaCBU=
`protect END_PROTECTED
