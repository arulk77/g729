`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIUBxOHkU0aFOLWhWWtLQL3p2aYTFIT2KhRWNt8lIniH
afF2OmORYonMkKXdgLgsy/cf+/Hy7Tk9L2dsqQjPtzK02bO1iThbCZVlDzooZA9x
v9Vn2TGdDpzGusY8gYj7/q9uy8hwBUFkCMa4OjfnY5ZNECUpGFXD7qvY7szqnsFs
qpyEbT60EkAc1GwasJR59Q==
`protect END_PROTECTED
