`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePvBxLpZLTWTHcLraTkpYxWVHLTkOXE3Oj4XTddh5SCq
z7xo0PVYQCha3/Y8j7vSpB2Rpx44CfsgIevnDKtUvnwyC1EcjdD7gp8UzkOK2+0O
bX+2BGiFCtHplzEWfqWqlFkShIqJqTq6E+mhVfnfYYlxlgVh/e6jH//d9pUOWx/p
uwbKNV9HE7jKQLi7RU1lxq+7PyrBj5pgkgHyGeqsTGmFd9oftodpPWMwgAaxn+t0
L7V9Wanla7MkfdCpmQrwK0mg7kanmRbBfbYO4xQFuWEoOoOY61UywKfkTo9/RQI7
/kdtNbVMXwXOGMqsuXnrmA==
`protect END_PROTECTED
