`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDIuy3VexIoUxUFr2mM00Rbk3S9lz6WK9xQwkJWw+eyk
gKXq6TBKTM0fwunz5jsrZ7JgvI7oEHVc1OvQsF/n/n9wkBrXFWybf5vSxaGW30zW
CkPynl9WXcU02ms5nWHJZ3fkadlHGm2AR2TsI+SFkEdRGPG5PpTyqeZ5C9fQbKN4
NctYMc0X08N3XjpWKWx/f8dOAHyU1q62RkYyK/oo24HLPVQZQNi0rgJZplk8z0Nv
riigWK96htPXIjV8FFV+6iQd2885vFlNZu1+9DjlMDtoRSsRox+svRhrh3rf9WfX
SWwXrkFycekJjWnwMbV4WNUrmgrMEMAoca6hruVbKDOYT9pQ8Yvz6zeMrZXveSAB
hTyuWryAZ7DkovlygAwrnvfVCNRBxeVxW/wPSrYg7Mfu5REYlshl8nn9KEP/knBz
/PuZRoENAK59nVImwN1RzqrDnxivnQspxWzozUJ9XxI9qt0KicgBqD79VyOdjOGy
F66yt2secPhLPfBWlXMWFg==
`protect END_PROTECTED
