`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
7RWERbz/SCu29vx1yp3KRCYfucXYF1+5GjeNt7YnzBozXUW6ZrFy6U3h1WifnHdo
yZ8zSk83xqq6m+/nyovgICUmxbeLyUoeZjUCiD0ipHseEkLsTMiJUb6Nuwo9p1ua
yBO9DZWfhzVcCJEZKJOzdb4ZDTdvLtmc9jGk1Dm0TSQLg/FQj2pvBcy5+v4wmEg7
`protect END_PROTECTED
