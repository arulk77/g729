`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEzBHiexxGv4bgOsH2eSSExwFrvhpFtWOAi1JZoRZf43
RgiMc2MFEIzH6VmqpdtdIg7OJ71nCE4HFYEGdXpw350ug02cL2EBFlHYQ6HtQIK/
K2ZU9a7DcijobPYVuno0rg6pjx5D0iK+R0cDn3ohycNkOSsn+2BQ1aP07owdCfP4
vdOJXq1CJ9HGn1zT5LsWmUYshxvewtWzpDZ9024/mlrOfIkXEqwXSbYNlM7Me8wx
9sNjzreXJ6wuAqcPbj7tyDL8N2pzqXrQBPog0M3ohnVYL62kB78jjnqcxM3YfqBV
W4GzGH3eXXrzuNv6gJVFwNZJzuEwKka0xLLsuMhnt9yg9WTYWA1xHHb+7o139ljV
f/trvO1jE+xj05QqmsyRzTFLohjm0NmRdo2cG4mZu+DeVABkTT6IfOWoe3h1VTLo
JIcuVMufo9vAVbrXP/MfTg7rkmd4OnETCiTpLHMsGVX75IlyA5d3Z4ZdUGx/YQlU
WM9cDb9lx/Vxlx/FjFdha48JOl+mr+cctFuNWAeCpDstEBO56Kki/XxFx7T5syIh
mzH6iTRn1gRM7PFJTVck9MHA5/6eFA/Yc7ppekgmldbyVfPjG/ROlKxbjrpViWie
puLzs43s1ibejrlW949GUzrYptFF2e2h8O6suuF7b4b7FYsKGlsITvqsMKjHGfTU
qsFA3Zus8iFIHN/JmUWZxNaWADaR1jjs/bLS47LnC+dxhqmJDO1JLzQSNYSXiN/O
9D6HXiEaM8jQkBDpTgpc4A/UyQuFC/cdnMZqG0H97yKo1neOvo3y2VEeX8vei7rb
32wb//QMRfAvvjVyLl8sn/Lt5adQUFu6w5WCOz9nbXVW+bbZBIgdQ9iDx+YrWYZE
a62+u+iDODNi5LdZCW01+cU4x8eKluhAaUVKOaxQNKXl2Q5DOjGEIWOKADSpAMIf
1ED7rEIyzGfRfMmmcxoWPR/1wzvvVKNMIx16jWiem38kMlSO0VOBq8kAVCh8eT4e
xc8Wa8Rcl+qs6FZzRkOS4pieIRExF0BMnJuZkIzjV9vLJ6EEepCjkDHectRIwJ7m
rOkD8SiuHRHGPhM6NMl62NK36t0HawEAyN/THU4fxjEG4Hm2EjOXerY/7jVTM06h
8DlK+1nVxuCv6Ku/9+L5m0BlpesphO8wAJAfMGREI2TQsX4QMYPOhQ0NlVZZJy5K
xbtXZ3aTk1lCnDyVeX5vtr5cjDhta9aZfy9QL4sfiox+sph2gRBWHrZvJgqbeuDt
0kgewYXSpqb142gcaTaH2ooEill4aVXcyBszoJh5OzJFl1VH0S3w2DOgrMRxyv9+
U8H4iChyEmXQAkfcEb3JUf3WiZTpCgUhKGVIKopZ9Ah++Frtz/RuJrU5jfnw5Lkf
EHMdwcTWn4LbvUUEwE0jC4F9MJmPOEEvK9vjCyPvZNjl/0DXiioP+tUzsgcsq0kM
FlxgefwDSW0S5zEW82o7ttEeg9sVuiJYesGEkR/30ybyE/KsOczfGJzQiqYD2SEL
343YAaCredvDsP9K8xore7MO9XsjFO3zCLN5MO4BAofM8WHUJ07ELMr/BpjyBVQj
cktwpW5kh1JDJbVlcFi/ajqpg/K/czV6I3PZIFGGxa0WXFO34GOOH/eQ+EXkiKMw
WcvgKUctmnbfLY2nyJC+e08O+utFPocGhVLOW+vQd1FNApwPVEpCV+rVMY+if/9R
vQuQgXJRMOPSEjzaaurYIk8q7UUnM82Jt+Ydflh0RkJRMRZHqNAee1GT28OLI0gd
qZh9ciMjTl5466Zvmp9Jj0HINTIxYbHzfD8g4oOdhFqqdIbfp4T+Bxm2b52g0LFP
gb8nR6jlUKs7XxaY2IvZXzO9x7SKjcT2eonHA4m3l1s1gT6XVDPOlXfebiprlw1i
pIo9hxfh1BAkq2J45S2scYcz8t3nUhryccLutViryBsLzblE1hQj9jmToaDxtMZb
5swbws4UuqHits5qt4qCNW80CpOED9baRmzSbL7Ipk1SaRlFajDf4Hkqf10rJ2oc
hz2OyXaJZwUPud1EttEra1FzUp8PHpx+oixeZkmSz2g3m9C23IwIs/9ftzNVeD2c
xhsRyy5beDn37GpExS1AmJP57egfAWM0eeUXYHaUm8egyqqgcIZ/1eLhE7yIx3ss
fnbaIcjZwuP7/NbFGksxzrDje0XJ2LPn133UaY4CJ1CThMANyOmu+mBjjitgUR2c
c20lYArM+zwAF1vt/lDwGovCqfowyRVlV3L53p0vSZiwUWjdEbCMbhRAxTc0PHqz
GwbBigxhtYslgzPrfyDWdKtHxct7eGtPQY5+P48ToT3ArkFzLQM8G5Q3q/FN5waf
TapZZvXQnbXSzWlbu+79aUsvnofZ5/maJbB+eIIQLWOl6lAvD4yMX8zW77LMVqUH
pPDFPgX282vOM3kG/OCsKDTircfHRHyrLVLDQxHjtKyBW5NebUKUibS/nScgqKj3
68GLJbxQN8p/EwOJY7i7jPlsuhCWgt0ZwiH9T24Wt0yGvEPv8kuRgSvwI3BOo1HB
dTklW949GDqzZPTNGyu4RhOvsn2Jeg1zh4XRptQRomLxRA8QtHuN9wn8xX2u99Ud
REwh+aVnEQZKO+gasQyux9s5qSFXIz9uPq4FG94mzsPzXw/Hyo9xBOWXqHU8iEUA
2UW/ZfNjKHhsCvVyXT7F7PypFOle4OWgl8u6FVSAuDRtu8kYv2220jXL55TiIWk+
Y9RjbAl8+WcYWCFystkl6fcL0tW1T60djbeTmbOrLVl+H9FWKWeUj+ptDztnfsAe
H+SvX+b0tLqKVb7Lryerx5rBxnGvBLog2xd9lQRrFryQQm3N1aXH6r6zSrzevXxh
rrdkIN9j25IfOsLk8ylh/v6EzC8ZE5xdgYitGOFLWxCQTngjFMWaipzO8FaMSRrL
0JL00Jq2H3MEdWeNXMCgqfJLN3LK6byDe/md3obwlLpFZmUeswkDvlvIOdVxtvex
6/2vREe4FjOG7qo2b8GMfW+ahG6HqC5o36B41TjpqKU/8OsCVejY0i9kz4Keax7U
x402rpzRNcrZYVq7gO6BnqYE7hHnzmTeO5aAWYZH0F9cGDv0sjW1EnI62lN7Aa75
JYakM+lwugM+J+NcfVDy1Ujwd0PmznBdM+sLWPnNw9W2Rp/KT5YGj3p4DRAW8vCH
9gVl9l3atJTjCNEZ8eH7pBfdpyu22IEJkgu3nyfhOuqheomoSEGPTP8ra4TAS/EV
iktoi3ZEqW26zwyMwAlm3pI3YHXQuWIVYyeUFnrMU43wIAb+wQtrYQK1XUaORZTZ
gMxj/ok/WNITDiiNXPfAzRnjiUBOW50KxjizyPj46pIe9NT0JQKNATlPIeysl3Ep
3IbL3Ae+M9oLQZBblbEzIyesHIqP4RLWA4cW8JxJEwbvezwWFZ4RH3XozhIEEuIO
DN3zstMNEd/y08NSDuyUXX6EHxdCSZ6ilL11Mu2t3m6J67FUuaI3tqw0FkqmSJxC
G8xh8ED2jZ4hhYqFnYeD/YiprgZkPoXeI6tf9PHL8hvvcwk0PD1S/2Ea5N2WhiJy
LtFtkCGMJc3TNVT1F1oHjbq59atY9CVLLKmmsPu+gRe4cgOvS0gsRzu10t7zrPlU
WVn6tdX+yE3s/c0uvzW2aamComZLK2wKhqF02RxXZCZJmBMQtLAM1lGUGfBB3wFf
kiNhh6ybENivtPDa+9tuyLHTqgu6pmUN0q7fRz/sEcNgraEpE6fHt6pIvkJFj7Ay
jBcyxjwhAnh9Kx0TeHZ1EP1a90yaotigPzdht56YUAlkgzAIbRGKnA1Hu33vHJgF
BQrhar1YBT+1hS1XDMHKMitnxLo4sopkTll7oZf7zOBpPzYStx97KD6m8Oy4Nq6W
n1GCWKh9KSybL4UXYELJUPwnbCcgdeuota6qk/wSlqs7QeFfVodBlttIfcX6Zsco
q1GMaWAvqXdI+iE9YLwWMLq7vphrS1ZwF0mU04qspqpgJbn+xd8V9F3LuylUCn2r
+KFmErlb48OsMfT/oFuZvkdI3OG/bWdB6I42QI+ds+zuC2S4KIUWFFtBJ9WaGP/c
UgCEWGmmLm1hF+bnJAuToACYLgGgAenhCq0Mssei52MfTzNEvLG7MOjjANVf/HL7
isdPZ1eQMR4xlqquLaltGQFr2NoR3Y+UUb7G11XZt6Yh/iSvQSlHW2ShooavDrH1
NNd87NMHZ0SGVqhugxCXwN328EHkdlHLFRb4ev69VR+2iT7V+Y1z0pjlQoGfotpG
OmJFRdsBzf3DvrcrCdu+648fjk0HHm6eCKCcx9YqLMciBa/4K7elJhFA5Ufk6zhO
ZOUZBzDJ63J0A3jWI5JjlCWJeI8gHe+/0vdixXjOYqkmr3zWYaZGCxkM4JaOWCU0
WsTWRzuENQ3elspaQWc6WiI4daHGXZTK6hVyp8MAbOtpMCOHSenAajswJphBzlDy
YOMq9XDKzRlV/mbdBmNu2hc7/up3/TM9fth008yTsD3L85+zGiZ42AFv3Mr1hadr
QOl5YVTtamipUT4u/GWQ/YM4ypOGf7cHq1jkiZUTx9YAk+qsOg+/3DzW1t/eimFQ
vHl4lYZSz/nn/rzVimSR6yw3YacM37xia2VhmMhNXyNTvpQG/SC9+u5PWq9AeKrG
K9t0O684mqqoA0EHWTyxHmPVDPj+cvB6Y3EoqSI10WLWxlb7RYd8Scsk/2FqNc6z
uwLhrIN+Oe1cLafgXfc7Jp81gowUe2nueQ+VNNxQLzqTg0dTobRVIy//8FR1U5Fj
iN5B4A97ldotn5iHfbo5q3GIXRLJaJ9s99vRUTznMbMKHxYR1D8Eg3WqK09rUFDy
nA/v6pOjdGg9KaOdTEzQx/G/p7b6OtR2SlwbHHfMcLhSEC/26NpEmkA3IOzOAA59
kVWEdEJOW29sXmappvjwJJYu5Tcya4Mo6iKoWsKa5aA0I3rTosmuCr/kEIBt5oBK
hbBtcZXHRS9YTggC7jzlOslpKdHUhegvCLNsJsIyrVRNb2Rxq0HTsBOp74fSQiYK
prDQLqy6lT+AkrhjiMaC+OABPY6OklmVvJDndC/Q27nOXm0aYTSS0rKmGek3qPae
oeJLGxZuMH8S8UH5A6p9eBhp5CY8lN+NpHRRZOxB2ENt25kprV5tU3Evl2kw73KH
odzsBddNAhzmc4FDNg9J1eHaCQ5I+4hghpCdN4+nxV0EVzfYb6UWtTrSPkVdrwIy
Hb3UZUajhHEQuaOlQMmYl8+52u8I5LZq10mlVofyni5OTdq+9lbiZlGUH60pQVfc
eLZJCU+NSSP94ctgC6jG4WzHPf+UN2c1fV9JNkw9vvNGsTsf/9Ub4/RwsEyjXKM8
ZVbsNEwODcP/cdREMej3vqZMRXNfnFUC0kmBWgSqFjpXF5mAoO+4bJ2m055KeDPp
KL5NkSx5sJMWJeXVOFchCKpFU56CHzzXETckqmjoLqFza6Mg92VeLCCupALDeja6
MZoBwXyK/9ICIFybW37w4FLbRGjAlJRyoAkAFwT2IxPfTmW0h2KnPM1PVHnBYc9T
zUbd28gCKlFFIqStGjP6OdUapf7kWfGEtkvwkd5XW1NZ+L+3PTrVd8M/swaQMuRg
t/Byd5PGjlTZaSzEeQfjyRz6QAr6joPt1pprgKduZYAkhpNgFHWt9pBdmH/Bljbp
J05+l5ekG2ATF2DZMbkboFdhVCopf0haKkm6Wxzuzu1BTNZwdjIgOtokDA1+YdXI
EAMSIcQVPUrmR9cE2jDR+q3hmSZiXFA5NPvkxEsY+T7wDeN6cxUBQ8zg7JOdFWYl
W11YzmzWPc2NOCN88FWOTJu7XL6QqA/vPNrjIfD0kwr7l+Z57azCrtvE21iJHOfj
RBuHRRllcS7F615jIUk6LK+Oh+PJEwZU9WDIKiz28jMeuH3CuTHTimpC9BQAua8+
zQa2qvKYkY/jtOPWDQjyA1Sxc2CFJx/PSsQDX5j6jZi81EGMxcEAJHEpgNcJTAXT
uYvogSVDDXaSGWzhhT/lPF3mONC2ekhRX5Kuvjvqqc2KKrfync4GFcG1I/E4COTV
FTp0IwoVAl9TjM55NZaHFp2X4i3A8H7ImtpqwXSTcWeNiMA3p+tdvDo3WsXjzlB5
ASCM5wC1HqFsiG0psgjebw4R9Q7SpLGjMVGk7KTFuhZbcQAZs1WuMEsgOBHglAG0
MPGk3/wHPfmtkkyPAZl7A3/naqNWE9ZHnyh1SiIlCxKghwygH1e+vTkcMHVVwV/Q
sOayL+Wd8nELcEXpQmOJQxYoiCq2GGgkhdMaStOxhAwstQcGYhg1SCcGT6ev+BD+
8nyI/y9BVc7JzRC41C4Al+5Cx9oQ1IL0l7A3ieRrFReE5GXLd5Z50uRWevDiUBhb
K1GTq5SfhvBPb5n0axIcpFcyTKA0ZrD7OK2FD7Q0pZ30bXTauZivbAbjP0LNjXHp
QoqG9KjfKB5s3XiumgOT3GPT9eIaQzPwe9LgzihC9WAaCqZpWf7egOojsjC6xZRw
pW4kFBimuicRwNhVvQY5kIOyBmDY5nTlBfNLULa3t7fFERmV9tnQZ2bswCDUUtik
7vs8c2q53cAErNsB6jFshu3+GkxrDhPdmoevUX8NF4lfL/tiiKrQMCIEzDbZ71od
S+jqDPj9/0kJRfVgzMnRis1EHwI4l3n2p1SkPdKL62i+Q/Z97KYyKZIbLgDGp35L
okSjCBWIqyg+2ds3RJJv1oW4zwR2T2sHx6DWPHyX3IyR1wkYPq+lTIMnqcAR9WvI
S1g7LmA7KY9xwbDVP2vvKwDvm+UlzwlgiyVaeJ3gkhwkeZ3fy+ekgv/m+VVwwbuY
oRwga6jNSuRKSK5dw8zxCEjIRkbxknn9cwU1HJ5dQI83CFCncAUafrBRXAprO9Oy
q6C5M7jh8tlyc7ZUDsIclAgSX1P8JdM6XhJl7WsaRbjU1TFcCluE0F1o+gtX+8pU
g/1YEU7MxyzOauuH2k4q5rbVj2oWlXbtA4LztSD2rJoxrkfngrYYJwSjpzF3AnbY
XWmTwT/wdcCGoPZFH3HJJyIK0ccporTBvvGQx4OI4HfYcue0Wtw1xyWGdcVMzdYV
xe6yJuPKMOvF2UFUMbiS+Ojb3H8eUnzuqlkHXwiYxHDq/cbP6p+cJCO8ViJ6qslR
YVQ6LWukl/XVgXUTU4vgrM3zWD9qCAj14pl8z3hAWoWoyyv1zD7uVD2VfjLwGM6B
A+VDtAdfk5OH1Laag+9cE4W2v3iaz4KK78duHc2RcGJ8PSUqbWJebuuW9/GQe5Fh
amosivHhL4Yl5Uawb7WLvQSFKXl+hcHTzN8Glgh/HupWV1LXS/B8RVwdcl5KW9AD
sD7ZsknoeYLzcwlrCNdSZEud/hBA5mFc444djPahb+ExYHqTQDbdCOPl8NNgRqgn
aVpcvLmf2o0UeuPLZNzKfarD+3Iaueu0khY7eC/tJYciLEyk1mhKAJZnfx64HaJh
t8A+Be1944TjLf8ZKWRPgEcYVjWxCXeWdxZ+ckxdRibee5VymV9u5QMHWIui8hNU
yOCvU2qLq7xiXIqwD5DnRW0UvsJwdjrgt9sBbwruQSfjjgNfplbnbN1Ezo6KxWB9
j0G4T2XSVa7pcrAcbbOOBpnVzHXtz4haGtSv1MXPUhkfZDFCt7NA5jpD0de/OMzn
kztdSPT4+37r+Vel8tEki7+BUC9fqDgWVYqfydQkrJj3PdrT4Vw4uOpy5GePd4kO
TqxABeYovn7vne11+Zu8/UTmXfNaMxFHjE50bdtaV48DdsOONJTrMpPJ0IdxDh1d
VnQzCLV2KeK87bI8OKkRtss7gZrhMb5eTt9Jlm12U0RC4hH4ZlzOf98/3uAN6Who
39r3fgbT+VQ0mhaw9DqNEjMTmvdExugO2rkGV1S+0viQvGBb+/VHaozKJjmugdT3
wZ2zyYyiMoVw28eh22hz9+ScBA8l4j+EUkBlHmve2BMxp9/uBQipA1he8AbllV0+
xjLFATuztPIUvUVo5H/4FrkkEDYtczPfOvaaxFiuVbiT8FANTBCSuJyEZTtzEzsy
Dba0ix3oicYZ/uzLCqChqGfmDnSUXKnMUQi/Gelo6THIQb2xLvEe0ihR8B3jHU2+
LXrAu4iHANw7c6pfZ4dnFYEy6no9XSvNaYQ2hsrDNLPqI/gTkxS0n0yockhLhb9Q
ge/P8H59jauhpEwtDq7Y5wot179wuTW6VtgIsOKcJW+psSjbM+dtlgSAfn2ce6AY
JO/BrX+THGmZ8hRzyekBN8wp27dalXawrpAfxVsurAXUxe01aUxNaZKWmMDDN2RL
PsjyyaJf4uaU44uB4UJwQhIrNoi1qLTCCocnF0kIKB6qEaOSutLDvzzD9gv0QuYE
kpzq6jJzLs1NpMoxIZuzUpzuK/3yXjSNx2z1zik/cam6FkuSWMB5Hua4OWhRU2yC
/WNBTcXJiZu777y83zJHfbWic+oU3FOv4CZFVyj/oFwyoaq4BfdYExu+Xjg1OdXl
X1+XlNZnNN1NXnqrynNrUa+ZSi42WzD87cVHPLIjguNALzVe2fK20jbQFd37/58H
ZY/u3GZhS7zTfFrJQbz0FDiCwajwTSS4gZ7mOvyd8brLhyVPQIvBNt8ORWamwekX
1USqeafuQK/YwaMOzjOwZS7/6y+gTlM1gQ9LMY63kcH4QQ4/QeM4Xn/eBrHtDTFh
erNjq049arffk8rBYQsCf50bW9T/HpWyhWcHI5jyHvbTOm7hSyk4k4oL3ii3cAh2
YXqr9fJxknt9ZEDEuGhxhpDCFq5MG0IUo2Ixr05wIpl05uOMlkg7c2kdMk7z9FJv
LNiXMj35Ln+LcPi4wCbvHy7+eGbmChV0qu8xvKFagLVV4qvlRbVTUdl7+M2RDcFi
ThuFCppyLiiM3Pydt6Z9rNBhapIbndxeJ7g5FPGOFw3CBCk2NH+AvtcJDMuSgvSJ
GrGzwlTyLsXnuzU6fzq/6Dm0ftFYWMNXxszyqL50Ws4JrAveVddNMuPslInE/wgC
NaBPXkaCZaGZeKCC5iVOAu3Cah36cpljdrbpNJMTis+HoV33tkuV4bRnlu/a+ynF
cBEfWrGaOwppzZAT9eR8wvfz9u46eCsm1bx6O0HD8L9rVIMaYB4b51CrugDa/X9J
RtmP8x0zS1Ehr7F5muh3L2vlJ+ff5UK7B5J9JewUqwE6viiybBwHjMJ/b2lqLUPV
6EP2IQm0hvFgALNP4Yof/K9PBOHRR4wAZ1o7Qqyys4AKrSzyBcIXSc9NW6UOj6cU
S/joYaktewTLvEX060vTHJw7N+1dr4eRE8dZHMKsa8l3L2rkEajnJbWjYzm3s40h
ZpEYkC4vY4MyaPGwOVP/nm2rNyAHUDvvYKxSK2xM0nbpMfbi4hyqZiRS5fhTRCiq
XFBilAAWt2gfPyqED+HbtfTUGvd8T23MKEB9cszt3o+MHH6XyE7coOp73rlADnsk
XG4GqUiP4tF6YFN2YzPuBpatm4J4JLkXRHdfJ4XHmGU7DYLmXtozGBnYhLuGXINY
AxrfMleRo0fyYJHuHuybp8EZsOxkCKeiS7D50Juz9dTeMtMq+4EoF2/L88rmTywu
2NWV1+ZgP9sO3Sh89hgzxmNIupvmYIypr0DEs9D/Spya0D56H/Zdo5DdpVwOe0g5
JikM7vD1RW62+pWZocA0Tpybu27m9RElLzBI2xj+GS6ClZDP3cYcovdhGoYrczqH
i2ilYTEiQ8yiYGaWXasyahzQPMBtD+kuK0cCIb1qOtpuezxAo0d5CMO/OCqe5Kul
T8NIilCvI7y6qIRIRMWs8entxJsJGWuAkpmFUDDIfQCgnMFC7usUL3czCVuLQ0xy
Vnh3nNmi8CSUzBVzt+E5nPlAKJl+Ygbl6I/OROFNixzUfkdZRdckRa/bVxwlc2CV
2MQZmivawrineRwaJGXB8b/zizZhqZNiWTf+/sJ59eYJ+hk0zKnTxH6QTI81xJrm
nUyrUNLVBE4uIQhijwl51K3eV0/rFu5wXb64hyBQ4qVl8qpqw7dq2V5ZLREwBKea
uN9Ba+Esyncty+wcTSK5Mb44s35e7klPDofFolLv8l8CIAJ4lSpiZCpn/XdcIHRN
Y9U4MzTfXKbHBm8fQiXY4kD1j/0wqjSRQ3WbMZjNbbLvVdkh0ElXKm3wVGJFfhN9
f9EVxbPoMwLtvrncY4WwnABBKcaxjcN8mRL+lHMGww68KC0vXqopVfi9jYzf4sPD
gby21Q9udqsp7YDh+nAfjLX/EEWIrLbwLyyKJ3NVYbKjAf4djzYjgCPL2/RRq2Pm
SzdabTjbC3wR1WtN/cG3xCp3aOJrzb3OwNWbhR8xc8v6veWm9Fdm+7QjSr9OsDn3
x5/AHi537IANqkIEOVVP4HsSGi2yWNkIdq+xQczvbCviUMhoClggRaeSOBtx9E2V
RrZ9Pjtbbql+tlqL+1g1sxofdO1nnJW3Rvs3Uf6esvbt1zp20roxLrp8+PdOTPpk
Z5JwuI4btFzj/PVBy2qjbUdwRkTjVjmsu4zo058503dGxgrP+XnkuoZR4CSC+1l3
+KXyRSZiK5QvoXH9Z6kJ3YpI0JLwVOI4R/H6/UurxucfqjCyG1u8pR+G/9QKM17+
calr7kqvo0E3x0fwoLSGlGjtArVJ7zFNeIh474kBeBZngbIWSXofeyLbk6pKDMAY
jJHaoGkewixZVbtaVUOekiDae4QdsCVMAN2piPiYVzSqG5+lOn5P7OWAvqWsulgh
eKZoLd0xg8J1phn+iVmoEPwI7Uz/LT9DNyYAV4V1cCNWU0Wh+6v75pfiWMnAoDl/
mYB5JmlRV2lt4IjzqQtjBYO73+w9P8cFWmaxdEapMTRCFmBukUy+itd137EMp4yE
5n1oYw4JES3i2XLcX9tzghiMOnRkY5ulnib+0/69NiF+6UHGig8u6JAZlE512mGT
UCt8fUazBxXr2UXAlod8etD49w/jwcIQZ06BM4a9yRRHCGmPgWZ6WDQwNWA+xU6g
flAHgoAAZGmRuNWPWXeGEa5tYsDpZMf2o6J4sNk5S0AKRH1TvHmAvztOa+AoAsFc
uWw+Ooh28qFqPH26wfiwbaTVpDBkLDB6caNPsxSJH7TfYPcE0dj1l1r/WZ0SCz6A
kcBQj4sr6Kp/VVgtwf4vj0UyhOL9wOr3TydbDWoZ282soAS7jAIp67YbaMRh1PEr
VoRi0pjXie+XKE0Auw0t3F6AHsS7qdH7sW/3VFqtq+2zynuIE2te0k6UzTAFdHTG
hQGn06mTSXfwYYPUtrBXtYifPPdvr665D4b81Qg0tSCRvv0iFlkNCOH+kRVoSWAg
0eeTNM8s8J1VKlRwQL9VHfNSJoeoTCEZVzLvNI8R7WEx+M51JO7kRVq9YFXqbePn
dPf0H2XGkxJIdOZhqYrJmsXAlIyWH6WqqGPDCGoQAHlSpvQHr6BzC+A1EY343tO5
QilVt5erfcXBaC60hGkMkZS+6oztt0x1uFovHN4OBdrgWzvxtKHgewLJa4cDtHzF
DQW5w+ZaysjXkRGmA4NzrG2UijPdRYLqEFfhmF8tIBDAfFgghLYawIRRFfj3AeaF
Ccmx4jbkO4ygtaASnFPvS0PPwwtI8ufwO+d7eVlXJL2LrSPCXim17BflIgutZYKn
6/0QaKDdKrOu4a1vel41bG4Seu/VIiLa0nnVsLfEAz5sVqUPZvd7VMQBh4WyfjOG
yYj/cBvP+ISWTaiJRMQ+g93sbsigd5fX39VT+ugnQTAuZHFgEXfApqPb2ZGx22Nd
TbSDgC0JklZPbpv4GKF3xJdM2AqdK1wGumlXH9KQ1A4R37dLREDDX1hOTZMnRFF5
Vec4nQxTIFvPXnb9wMnu1/6QSaEVlymRxlOHYHDcfZF3R6x+3w0kzZrXeiDXK7aL
R853hCv3kHIBwrAwLYwLnkRoL3HvQ7pM2KtPDJVSSfxl2SXTZ766xfQf/H1nZXAx
Sfvxj/h/GSWZ4g7/T/MByGYa3p3tFAA7YmVsG2S1ZkoxM1iZIAX9n/ebOhvT1fbQ
tdf+Mb0hohwpgTk9SunzXG+on1h7/38m9gOpEVYbPyOifPKcFdEeuvig2fHJ2VoN
Un5PWIfSddUoVW3NjZueqJDdOpFwVKLlRAWZR3Ca084wWSrAx0MU42OwrCmcsvp0
okwf9IjqFlm+CZUostfQswDXG7lFolTB1KinX1bGCnn7EUeRolet2bOf7QMnCNgJ
8POyQfhbfHrjv8rpCwiqADa3TE3b7ic2FH4WWueM0fHvwUFWOHCZc1yVIZBRfL2X
t0tAlZhJ8p17ZG2a7nNEdsOZbvmta1QdmFlyiTDgD5piHkyEwlCouehVo/OG+3wE
tvE0BBYO0hpmODeIKtrj9kE5q6WUnCALCzeT8AvVgMQka2+2wUAXgsSG0SC/KGHQ
3nX3HSrpq4JUn2iAnCf744vvTut31F0RLsktZlexMFLggHXvyo8/bdJuejlg6uwI
sOuOJGsH63FaK16/psZINNJt5hL4uRNy6chjb8EsH2FyWV3Fr3dWomN1JEhk6P2s
6hTp/M3oeMLpE72VkYmbIlNt/iIIR7lrarjRrVuigTyMBjsO6HEvx+DTdf1X84Hf
UQX2Y0cd0MekyPQudiM31yOYtN1v4skUgR7v22eYBmp70AFJZXRxFVjUB3VHMavG
YXdYbArm7IPlV6/x1tf8v+Nk6+ynz1D1huF5gErqtYRJTkM8KhU1SQoAUlYIKMnS
L8n9edAE3lYDvoSAAuSAmROeHjLB64M8rrMWVLfEFGAT4VCNY1SkxXGUzdZDPjVa
RBI5bqZw32ppbYNbZqdKlfRqH8BGVnb1M0J1tY/mADMLtmnfG0LGPf82Lme854EG
IuSVGiCao1paJ5M1qwlDzuQv22rYARxw/GCSPsA884dphUht1yNRmNBsIFRR9v1M
02iDtJK5Uc4MX2EpP+uoh+v6+B6AGj0ZLGj97VaQWFL6MzGvS8pfNOSZtu1M0OgP
MqI1xprl7BDG/ipPQXg99Cl2hozl2f9Mvi765qDP44Fnl6ubkrM/26C4GeGPM8we
2eGyfHmLFgklbcu2LXUvDxW34qTmH4/sCySFXdYQrrBk7gtnP0brFHXu3k6acY4o
ty14iGlzGI0X/ERxL++dgkR+DTTu4xnNfP7pJmRKWIDI6lgjt6IpVpLtoUs7Uw2U
5snQjTOBCYGLuX2X0O/TQ8mBa7t/yByGt2fwEb/3Eh1DNx1AxHPIfGAj8LCtHo+x
0S2t3sx4WCfvL8fFTb1BhnSYsO1qwSGQuGT8aUv/uDrJnaFvcyPPD1efx/q69N/E
gfXDxNGR3gxyVmiCqTdwydo5k6a42YbBIdnY6fUMHmIaQKQ4XoCIw/WHDlz8S/2j
11ebBcmcoN5N/uwr9KqqR46/lVCwjOAiEUo+J4ZxxEI6qKyT1Mag69/rze39dNFM
bolxp2KsJpSMRI/wXVoLpul7PFVEZs+7hrPYIi7FjHEftHejRIDbuqGIrwfVjNo4
ltsyLHOf8bruvPh1/6rL/+KqGBpDrpd1r7jWkaz3KCb27i8DgteXNs7VbR7gUMYA
ySiZgqnWWMacA49CkhkziLuQnUCjwhTO/s56A7XHme5TOxB4dWVlrEQT3mKcfmsZ
pw5xvAPVQTn5uO72gKJC8jYgA7J9cuI2V0gBRqRqDs+pceSEKGQRtol8n2iB5g1N
CyNWjKyrNKT6ClpWYQcqaoFUv4uFKvKe+pl8JKcZUe5z6MwJkEeBfVUxwaFhmKM1
EzhmcPuZFmzLE9fc42KjiLN0zAfyoNIcLFkTarm0zCSC5jvMvM2E8oH38Xy3tqss
hJqCZz7MHg6xov6+98H02oT9TOVnrmAB8rSY/PccaRopfE9PBQjgv3p9DuuovqVQ
DVD5KhTiSU33bAaQhE6hz9I7CuSLWT15TPQQTgDB9cZGpUvXumjK5A7XIeO7ofCk
+FlFHgWICSqQz4Hf3KLI7b6UjuJ8Ce+N1NO0CG0M3/s4eMGA7AU/+P3CY9ylHeBg
Fl03a2HgMl/VDCJuergvRhTxTI+2vwFeyAaP6a5nV/Y89lA7sTWLhxmK8U+Lfvb4
qr1OtDIbe7nN8045q0hFtKupwMLmMNYgeJsSjs19HLs21z644FvtvDIKPnx1B0f7
rZw1b8g40ZFJDib0WKS7Y4AoFAGT7wJhq2NDXhmfgleLJSLb+oYbHsR4yDoRw1QT
ouTKpqsBSwI5RgBrVa9d9nPO6ugqtUsPwQ9dqzM+OraRx/2SxDindfRWkb4A401g
r+OGI1LWT7aKpDvFQZiPsq6JXlrTrwc+JpK/iiR7gaSI3Ha8OnFrcI9/t4A0GJJ7
cHUj9iLIZJfmPNAOYtfF+MCZ4tODFE6+t2l9ejwiaNDj55mZtj9Egh98wtxClj48
k/vwPs4aJ2uYUMzQd7kbHOeMGLxj1x74eUiqqGZdpQyK2wJxtHhZnNwX84PzH/G7
22Dtlxeux+QxzXFLCX0V6oQB+IBuDpiSkf2PS+0i0CO/QiFMMJko9XhJFNls/hnJ
BeeutBGqs7jxAgjM9b3SgjGwNFeQxTrArNPfzcTAH8B/NFD1xCgy3sWB3+9Jjgux
VlmwNWyYIQKtO7YAW9gPEgmDt6hOa5ODwRGCLvKN5zEF8tuVI61g+CCc4VJ+IdRD
a2y2wxkJNmZ2tgdlPoWYO8nq8Qe6oSjFj1zOEt8WTniDh312KvwtVUWBTe+266Le
s2XRXI3MCP3u7XN0xJ0CcT460tj1RzxJ6kZimHebxr/NIUhseDTkJh/kYMheDAk9
3zHYho6Fw2i7nW5Q25i40VAnCvRbfa/fZJWltfoPa7n90DTzgKuzqFvx8TW1wyzn
2IdCD+LQjisTV9eaYmhNwhGdF6IX9eEsuu0Yco0tcghOwMtZAMLLebjzRDfb5Zf0
vDM2rw40X0Bhktev2a06gosVKnxoy3fIX3nFC1PTH2U2FIQ7AUfpbtMdhAmysMqP
D1ty0q/OlnYRGlfyvSVIuIKWMKSTMVI233EF9YqOuAFyQSlROMdQirsDUojqY+ec
ZWrNKc5HX9xRUPJ3J32roFUjKhwbGfVxkYCB4+xEmf93KiNyDjqkZWj9PL8p3G9E
wBzBX6lf2unHcjr6/kvIaRin3jw5BT5OfmPgyNy5s12R1yc/0YlUpoAdKjgJtDl4
ACl/AwCmAdxj8veSi3+94L+a8yUCvKcDfStMGYdmoWwIYI/rAK3FOm1dhlv/dVeo
H3Sx5LlW5eKBQE1Ti4yClDb2wfvSKbZmic16Icq6/AwykY2E+dDdZ+PMZeAcLbvq
opI3mp5w6C/fGxSPp814IMgPecgvzggY+JnMavdaLZ0TGIm4OS7/QDwYzBphA50d
061XPDmZTcVJlHknsVMNDYb8HUrhBaZAYdx44UDK9B6e0S5LwH1AoUvTcKgdlNch
iPOuTwP8D2juFzEajJxcuSWK0MbMPwlAl4lmEqWj3UMg1EdlfWwIFqT7GfjQWKoZ
lYnDkYWB6OTRl0f626h8Gj8icT46d9K92RQU+eszHjqzhRMfwq0qrH0v7yKSnM/Y
/axC1Fe0z63j/6Crr25gPni8lDb87q+esUi+j4orIYGfxBeVPHTJOQbWlVVDtsHG
F+ijsgXO/paAvXI7Yblbpu1dSVKm+qKUIVXtFp8s6yY8RALqhHDkk0bw7WLn9ZTQ
8aXTHyXvplglu69MoMxsxm+HTSkzxf5Nq/nQeYNRBp6bRf25Nzi+KcHn6IkvzpWi
bfkqvLK/6QSrHob1UGxa+ibQlJj6M06S84woOUOZlDV0FYW8V9EqXheGjjpcNaR3
Jk9RoG/k3wmYEk1kf/sAClFFlkWRDch1CCnIklLe0Nj/MtU2o80+DRUngw/FQFdK
cf+rYO0lR12DNgfmI54vT+3YN2R49BdAi83iQyndv/sePFFB+Vbaj9l//uB+0lDj
wp8sOpa67Sok4H74z8bykmfNCHgV6EHCURAndbqgLJMTHxao0AZ9wEFPp5iAOpp7
pC6h7Kfq64b48mmfrbls1UF42rUPvZ0RoQr5k9R2WMOIJN/GPmHDAI1I3hcXyZdq
kfBuzjknei5BKOXaMPPyf5cdnOtyWDod6VLqadYrI0J0P6aoB1AKQw4CzrqPmAmY
8ob/hK0pT3B5P6MX9sAkxAGdGkAaM23Hx2ZMBcqycJdndMjZnYnCbm3Ymhjp4iKg
q+rVSTYBlWN1TgwVUyip6yE7WoswF2Hi4qq+eYMnqJ/+88ZblPV7KZltjzKa/vm8
OOahSPs1wr/0O8dv4OOK+C0G+H4RS8aDK3qwa9HSq+BfGp8tHXcPMI7IfG03BPgV
9xQ4jhD6diOvGtmRWQl9WZlUGpQyL8+4sZORmIztZS3IyZnjJFXrgrAYWAyEFywy
0cVMEZPchKbcPT/A4SCEhWvBZK6iTdmGaNT5do6/BOiWaxeuGhL234uKpwbwNzTc
t57KEP7EFVSI2xJeARbs6Oag8HqMCXdICmgXLSoUpUN34qLfv62p80RtVvpFG2Pq
WFEiamNt1kyw/eb6sTIcbqnyU3omyATnZOoovPfucHQp7ffOsh5fjbNjePHSSm+/
k+x74RDizOocSe13auWWVwyigFGvcJAQnLg5g6Y7MSkTrz9V+xoyfvNKZVJEf67p
9dD7daErRR8WjO5kwZ8qbfhzantNu3/cpLCA4+ii/cfu8Fv7holwwVc628p/85vJ
1KfZk7HW0XQKjrgr605E5U7C8+cwwSMyx+H0/VnF5PclYWj3rPtHjfh+UNjCxxb0
z8w9FfBtnNfOuXH5tWL8UGfLtgns2CFEY3Whg7kl+hXlPB9IOih7oyoQaxSrHX4+
wK4vpZvflVtHfu8wDILBrCbmwDCRvCudEwht3n94cBohIHb5jGpMNKgxnt8BVnv/
MQ/QrWgTRegWGdZ8dD3Y3YJOZXGhz/cGtj2E8COriMw0BD6j0mrw62qhOnLisQk7
m3ZN30r+oLd6BBDuyfgoK0RKRm4K4sqyOoPIH7mcgohAC3ZW2WjzQkqKLc35iyvm
+dpfaCRT4HaPQZnWWBp9fph8XphpoakS9adrHByQJH3WxiyWJ4I0EuB9T4LtQJ8f
FyS15n1oK2FYZ3pdLSbomqlvtgahOYeXebMnIM9KoXsYpQqZQNb1hT4//Jm8zcoS
XwduQMph2cFeSLepvaFKUPSr52SdyzwPGfmNYdC7aCIt9p0TMu3LFTXvrjZRt9U5
DaEXg9kstsRigk/it+K9nlr2iWp+f4heMjeJ9RH3z2CZb9M8tLEFxN4b4Z0N+FOj
WZxojduNzDrM8pdIVdwKnGvDmZKfygjJ9PjemJsVEVyr9wtm5KtLCnppBVYUdfnl
VbYS7cO+LPXwvUyi9jles/0KLSLP1yWnheBOJzjMahQsJw1qAOAuMsKEtYAkNKSC
WFTcQws7J9ayolal1aFULEfvIUkcAK3Pxe389ZROY0N94c88Pb9vZZ0BME4nTb1Y
4jOdYgzQaB5ldu5GvJ9ui91+vDLEmOUCLgWYZcS7Cke+P6RilYM6T8O6aRjal1Yz
vNv87Its30/lcxoY2JYSFfHq/OU/YbB1YHkjGDzybAtT3CkM+FXzKO+1cHW7CZyR
CoieZAlrOCxZy6NIds5Vt4l7gEjHtI9W4d5xnr8FAAdWk8Js1Qr0i8flqGFRzIR+
41hpBB1PqM/+9c12gWnWs8LYHNs304qbSyrQhDUaPYdyIBHD1tRr0BvyabFdBjn9
EtvHfM7TIrCizl6S5gKK5lLqjtZVa/pcUGAHBNIWRNcdIPQXiUIEbqizki8lPHn6
T45tLziWEyOe+sHLfSf1IA/tDfNczyn0pY8fwFhO5yIfv6yPg4mmCO5mOnGUV1ut
KqT3RcVrKHPzH+8rUNERJe725eE6Ebt8tEceGF8b5EsKMmh+PViDpEJW5ywEM8Ra
dOaht48AMRbV8eOV2khB3kxPw2F3/qtt9fy6K5v6dxY40PEMQtlvRnYM/dhh93oC
y1KpjAp12PpZSGHVLDr3mTMJvKp3Xyt068a4qEWK/yVgSHCGwar8rqX9WzrtaqHD
kmzBIzkjWwUKnfvZi93t9IF5perbBT2KqGX5714pKsRA586UXz3v8JN/K/6l4kqF
Dmm1FeETcSUx2oW6lCrfr5aY4xKNvOk5HB4VSXhP+KOeyIjLZDDsV5sDg2koQDig
gxbB+CjL4XaK8JkqqKU2K0R8BNWYIjg1Jbq2pmQbv+sUQq7b3md6BpotwzTwgBIn
/idzxWmjyNG1s2q96mBt4RJOaqmRtkN38x8kXcuC9TzfzwukyL/BST+A92qZahTY
qjLlCuluGtHf+u0kmq0qIECeUjTHlE+VsTW88sgm1fBvya5jjbHtZjH+ZeqaC/wT
kKYYWBDRqhZ979j3e0n1zIN6XWxgBQYSBJewMKT52NaAQ1HqXmCwkDavrRZGAuTW
vdTVC0eBGOd+iDLhlL9lsFJVtwhz61z9oSih5hvzpDCwLzit3c0eNzDKp4jevSXB
irsFFYsMTcvKi14r2A8vFFgO/y6EqaMqd2wifmV8tEUkwbvX7Aerhi0Fs377q+7/
JrimDzSiVvD8/wKPJ9k8lfZIrG89hZzeaWbJZhC+xLF+5anc+ZdxgJLqo87+8L2S
xHn8C37kQi3b751JRPhoes3hZ3JVs+QfKKZh7FVHuf+jPwzybw8/NaReQRaHtfnG
ygyN7r9il3fiy8UfSJhgQcwfs7LK5kyHhz93yMUBFFK3smqT6OKnNvp3o/aMTpTY
G853AGiRUdie5XxYB5X2wIuHhFAkVCOIXSGfU1vU4kTkUbHEQZWzaDwG+xAvolHg
c6Bqprjg2bw4PvvPTfoQEZwkp/50B0v+3uCR4PP9j0ZOyMIJCdHiCtVPlT3q8yz2
85W3J3pbqAUWK9KYlHMvIBpg9OiwEMrceKwy+Xz6aACzmlsYwAaH5N7hErn5CYlK
BKm8WFIwfwkpMKMLVNQJGMbF8NWyu+6pMQivGUim0cXgOpjJ9D6OL0y+wHX91Yqv
beDbyBE8ze9HDEulqhkf6OHNAbK50wC57atPJq1suxXEf7G68Muxt+CwhEdGmaDf
UwaKuUE4xBZVSlU1yBy5D8ECc/7ONoMrANqA8b4wnEra6sarZ1emGDoxTmRPHoK6
Nyx4WMfVhbXbeoy5wFb4xpL7kUOiYPJxow9AEeVKX7Up5kb/8+VzcfJUcL2xSq4V
K/TiX6m9fkGB//IvkxBWCA7C7fIFVFY91N2TrA79rmIuGw/x4IreS12Pye4UAA/b
E/be703MF6tkxlcdsaQb2zU+O6VrNLrtEe/3DOI21i9CAsv/4P6ajB54rGj5CTH5
5mWspYj/04F8Ek3ErI1HzHFW8Bjq9ctoZmC/9K3qJuuCEVTdx/C8w92IIIotT61f
6OsAaF8ogQj69Kf2PhTG3uFY7lXRbLptcJHNSPhy5fU6Rb0I2F5Eg+oeVntS5kkr
UV6Uhzp4FnWGCSkGMPf+ozhuX/omk9b8gcsHThoeDyTak8KTddKBhxKKR7eMlhNl
ZqDORslw8RI09YFOyzeFDkw6GwoO3Z7FIiGhtI4YpZnuMdq2N0Mlrwo4d3Vgrq2/
BkuYktiwNjIoAOVINl+EZjtz/1N/XXuStrTAhYqQf2cEB1xWtLYa4jT9oIPVpdcL
lMqmMVuh3//42QyZpuq0s81MzDSOoxrdOoIOHRXGANh5Mz8Q9do50LwJZLD96jAv
A9OkbiESxEJP7gqbxMVQ0tDOwyx1pu6Izu3yC7ezucTPXo4hwECyQPYzjjeGQqzF
+cf5q5k8pP404AgDtAxF7TjpwTbqoQ6X8EoSecFyTVXlF8WKevXPSwWav9BSrK89
3QE8ImbczSDyJ5ATAjxRZ+RKyrjyMQw8vcKrHyHVrkLdJwHfqr9ENOs5ZQ4DTQEl
fKtCSJud4lTJ/C5ZwELIPkHReDtv/6YFw0z2H86spfwFQqKGxcxZBSK94lnMO0bQ
UzJlupbcPG+qaXpyB/mfe5XQxZItkLZLAce8jYzQ1Kfn9lx1T5E3f3D7GGZhlJ1c
gWgQvFcpnIDY34Zm0G8Z3c3w5azRGAxMt0wblk7+aol+eyPePNWEyh4M6Gdoyqnh
GF6mdkuBvytzoCtFQfTCRK7ueKXwo7TuU8WYmHuP/KyHz6PJZmKRCk/XVGCuCRCW
VlIWaxp0BaiOoER7dEFQmrblJ+y+Hith9BT9+zSxV6JKProdQ0G88VpcIxkzt5pV
BQVUjnS8j58umwxK0SrFZfwEB7KPevP9eqJ8MpImi5cXnBsyCJvBHmKw8GSvy15l
ltBFTMXReGXcdg49D8o4H7/cH0CrN2m7azwJ/CqSaIJ+0pVwftSUz/CHwsRpXCD7
Pkz2CVUVv00vnyc9QrCrfU4pA2Fher+5ydszYfJ52BYoo1GXIfuhlfATr0L9cGOH
ve7qDSeoXvjT6Frk7b2G4yEabdlnUJYT/OAeNfLgl/DytFfloSTlKGBy85HB0apN
UssR+3lA/YpNTs6NHCkf+1JA1EuWM2x7jfk7uFuIPYZkePop5Eg0RmG8IVttDrVC
M2UKTmUwLpRkjSut/l4NiU+5cEkjfycyflBkYT6pclCMJyHdLDcFhtbl4Fzj1Vnn
6+LlgjfuSq86hepBD6pT3gib+LZ3MFGK/IZGyhMyNPiDjUMpVU1D678/42UjSmtO
zJ+abNJHjZehQtB2twKwU1HQmMDTWjmc1BiicstNnlCwR6Wnjw0DyKRZz8XsCk4b
m10Fg0qr+2fMK0WEyBQEoCiZLM4QuYCiWTahAXibGXEitN+NY3M2cWCJUN04rq9d
AZo+Jqv3+2rHoHPFPSz5qSs4ypwyxHuT0fDGaFxQhx1OyJZvwnHDCJyha2faTuKU
dhwp7vrPeTQZ9MKg59ccurnGq/I0XrzSnMq86HRljek1B7BOKh7GL7lDnVXFSQrT
8YlNZBpEEX5AYccjpXl+35BxoxSuRaYqBJseWxQYJi2xuhrL2upSIdM+DMUWR/QI
F8f4TeEyuRRA0XA9StDkpqYEcY1NcbOxtIJh7cXWnt1Ak14fn90BGKqh6Jkho/Ab
3Si+jdr51jcMoyYoia1vi791tVxlihICoV7zX63hm6csgt6HZ4aZRPTwK9jbs36h
W8G48mVAgqsjAGyYFHKpEnAB1tli4VjGkoeUjIO7H3xvqy0zGwt6O1tg3MntnqI6
If1KnvtKZ+2tiR/UMmHFMGV2PB3kwd8uRwe7yvsny/+UYFncb3OJQ0CCHVv34Rij
sA8BHXv4XM0V7zrvEBgqIz+ActOvWo8qCNHY+dCkd7CDSdKRsBZ1lpOCo7W7ivcl
kUUh++88A8PzQgRSIqn0CzT0Ro1YmoJ0muVI3mRoF4NVZvdTisFP3qyQL1c1OXEa
38H7kJliz+y9MvDyIq8Em1MyHwNB27BHmeE4N62lTXs3iAjxDgA1PEdbwl4iAAxw
J8ZP73QmOT6MGX+CX+nboAwFmYfGNQtLoenOLCpkrI72IpaE/CduWvYI0g2SigKl
RMERDWP2gFy6gb/GZ6G/4gmywnRLcRqzw/aKfPn1jpkWGSDip92aP5Ax/utF9q1C
XsVBSTAorvwdE4HaRYLOmfX+fKHqDGIW5b1nDO+9wRH7TNXBD+8vyqOgZ574xadF
NKbsuG4FkyY8YgWkJJS2iAg8HVlx+cBhykHEFvF+wkG5CQBIQvDEU6H8IwJnXnWo
YkavUFW4XOX+qvpjLN4VCMcHyLvMe2ZI8lKZFOSEU69wUeYstSBCQfQ2HqHCqd1+
grPv3H47jYjY+l+Y28YC6+OsMnubppzjvyt1ffx8I5Oooa+Y+XE3ppEzEw/cp3yZ
IXGvSRJbaCi6NwKjZbf55kVOerXNwzQ5VLZ4l517EJF8YG5d2+p1AfJwJQXSHSB7
b9uU/VCEKWNG6FIhQIhNOmJNoLB0lxqHtjNqc76PVtxzIXyqv/Y6xHLCJU5EwcSj
6ZGDnaYFvBCl9qJtIvbPayo287Y4WMu5wtzqWoe/IWaC0o0qtEaquAi38sMN3ed/
ubKUVtHiDKRwpoBK0sIrLxPU1hESsyeMQKhaxNtUN+uxvBi6LxZe3+plmLvK+z5i
34s1qAkyVUo4Mg2plkf/lvX6aSfrxa8fXFbt9cB7DugDVZCH5M/8GYsl5XaTmpxB
8+D58XXtZJg0ezL/SZLEt4Qlvrz0X62r5kcAg2j86rP3yWuMZt3SdOd/BARoOfVm
4RQsIH4DlGRH1wkb0xQ2lD/5+6+/XR+TAjcL+3uwY+Ho5ivCNsowfd18gysmCUSi
EXcxfkv2dx5XaUWJHiPNPOaanGDrhF6h+7h/4gT6rPWZJHA//hUIoVEMsl3f22be
z4+bczWUo0hOrHMV3v6MHUMl1/DuEC9qj+xb4bHKUGDOk53J2t0CGNoXV0MBXk/+
1vzw42N8iaV55xvkm12P7rOGjd1SpLMI32/2y6fa1Dkc1DDd1sDKAPE9uI/tUfvY
w2rUGH/rjm6W8SbJCnIEKJpI9Szkkaq4FbCLp/K4g/BzEaUeQQszxj+pD8+P5wjP
9HsaT8T6r5xwDA7kTc5O9E0qlfl/F9NEK05subrjaC7S883E0jMKvIyYTZMYQL23
4MrpU9YzacIkry0xSLSaPY0tGmK+5QftHlzKU2x/LvnvjCpjI2flFmdETis5k/iK
GKauoxf6y9BZ+udsi6Z33xJMqapRHNDvf4NDB6XjoJhfF59P2k8MGnBQaopSJvkn
p8isPpo85XVkEaKcLrjwExSci8wrza1eICo643F6tOMiNe7FZdjZi07s8DkulRbN
r5xntH5CRiGwI1nADsby2rvEfIUKzw7etR6POb0qu0JIuVSXkfkEkQf4EFVC5PCq
1sPd37uXi+kOrHqLKwmSa8T9zVnqLtMtLfwy+AHdpfckrQwFWYxGwE+t6nEiT+bv
dWrHvC7wp1Ml0oOJ9qjIgNLdYT9QiRGMN1U9KHaJBuB5GlyPXxLpsP6aLi7Qw2Yg
HUUoBWAtpMooj0yxHikfRvY/byaAnjWCMTqwQTCXhUsft9oMki+8DrJhI0qY879G
5c3CKEXURsbLtvuJh1sLSRBP9JXwpZm9xepTcUrzD7v6PP/R0Sji6vM/zUwRJ2Be
HkBSu/7A3C0jcN60/vLAIbCrtb9RRq9V2rkp0fyvsn83JUTNEVrbxLOFKDt1Jxad
UBLlXHlDfgFTZZME/u+VukaiWgB8cDqf1xgWvrul6hCNxrTrmk59QqdOSDaWwORd
0pyxKsB6XSfkZDpNgKIaNocmhE5IToYYureuXc/CpB7cE1Xshkp2UyDFfLc9AivM
byAluZhxzZ3++LS0YtWR0ln5NxqGi6HlTLcc5JSGPKHwDZjDwmLu/s6sC/RcaeuH
GEiwErY309miXWboL3oDI/8PU4+DoGME7ur5wHXro/lHg8qv2my/EjVgqlMa6xcF
EyJL1bPI1hxQ9H/rKOwvGjtl+9h25tcGERLfkHT4zABdqxu7j5JPcN9qmpEjw8/8
vJc/OB9O/gHqRJ3qw+IjfmAK4AHZR9WL0bWmWrsLyYZE2k43DmrWykAvTzXf81iA
naLCGIpJdf7qXWqbN269bJ4SWpHxoet0HvIBfC2gLL+kvvv3QdsYgGGVYE0C5aAD
Z6H5Y//WCxA8rvdxiVHlS2HiEZe4AEQUhcgttBmTcyb1lKculCBhb1HCCM3dsPKI
rq+5PDnphpRS98OBm1BEndHOnqRq6f5ikAIUsp13VYq5BvIROk4+iJHnfgorWsVz
zWyOtRGsKLZcHvrEardQ7zKCabo2L6BaSan44puVzPzECCFVXpXxmNF2N3iTakXT
FtlKsvqLmvOkurC2S4RwwYbC5r5JWRZl+D9p6KSJh0H3Hk6WpQngL6H3uJ1pcPlN
kcIKts4QVnFGNhLU26A1YsVUzGNS6UMbSkgKGpOA9134E/IEy7NGLqKZqL1InpRs
4sPvZ6Kmz8OYA3xChLSTQnFc5qTBn7q3dR+ulYoTqFXkKisuOfnZIosTGFyIZWhk
6M9XNoriQ7q6PVJgKKR/O5K0E6QoW0830SULqnExTAkKIGwbSlGSsqlVGu/sP+Jl
JX2iXIQuie2OMMf44jVZZSAwGSpTg9NhpnXcIUrnWhmjwoqdLXF9Fr779Cv9tHbU
/MuBWjO+bFgtpUxl0YmVB1+swMp+V1hwVb1lxxkH8sWXnVJAWpdOTLDwH3N8nUZe
fHZUw1SS9GcFVl+IJqzJdjeyAMcQmqnn/r5jl8B+/eoeWBUHHn6/97RD/g/VqVDv
7NbdnxXXfCBhDjYgJ42oPHJv0uBca+uKSaNbkT+Iury5PWCg1n/+QlUi7a0db4kU
7boy/B7lJiIf52aAjwVWYj15j2UT1WQuXzoxYT6mrohbqGJbNMx/UtWqdNUNI9XO
1B+4trPFIQWSeNvbx487Xo/QKpEmutUUYhjfX5mDrB9ZLOhT75QsbfvX4JRCdbCq
NaePSsOPTIVjEl7tev128nZ4hwQR12sfdQuHBHPMaa06ehrL9yivlxSRcSckgEpV
rGmn+FOlRj0uwHpVzkAA/WoGCH+QzwMvDe9lTuwfm/kva9SOwqOIgocbyzp5LQsM
hsVxtl01hCRE1+wS5BA1MfM1f+GwbQk6iFMXXTpaUMnQLge9jdbRAV9ctyB6pVkF
S4mfCzgKVbjraoBy0RbiZ7AdAxpWSti7gQ717WQZoOSAnw599f04Ev72VlkeWowB
anpJXISLtUlJBlJDhX3xyotwG9WDdupnmBxXaCO4tkfg5IRyqMpFpUYimdbC56/z
FkSPPQDeUN7d6VM/yDansHR33W/JJDkH4ypfk2TzanDSGyXlzkilF9c5I4vem24E
BosIepqfJskbTN/ROMqYcOpj56AYO7bQholI7e4jq2O2qy1SMx4CiQjS3zWFBMOO
4bCqVMSLVbsPTCnr7Zq8QViD6vYRJyJ6MAUbmW8iZuJuI1UkdbOAvZguHlrp2LOr
2JEij7fqLmQrjzONd0fPz8ijD5+kRleLUhJNtvypittkBdhz7VDkQ9PV0wvYdYMi
VBOOfPjcTmReCrjluDZ7oszsfrE+h3h1RgkU8Y4sGc02TI5XS7SBVhW9eF72YA1X
VJ7GfCmE0Q8emXD1gDvHTzhGPJgkTZ1qUtcfjcXWsGZujqGdf6pN3lKOyiZc221Y
6EJYIaJqCuRQjSEzn/IP4/ItMB/iwU1FVSXgQCpo51rv1aqgzlARvlC+Wv1nk9wo
VQveWrZtovsDquQ3QY7Uacne4qyw3LV63fRkqSEW/1Y6JL5nJv5TNSHgizti3P/h
BBw1jxluuguRflpMENl2f+uNDc9o0COPTor30JDNlg1GMvbnsOWpSMRwsWMmaQiv
QWKDUeugMdo9VDXqTSJuqvgdryLiyZadCnD7n4QEot29FsKi2iXk7um2nZ5McB0x
KdtRfWWyUTFXivWDvkqoDPYuFR09P6gCoNP+nBpeOeqJeUwO93Qf0yuY9SG3wS6O
NneOKdqs91f1EF5QQh/c7oQahLS/OKIFrXC3FHPscbGyuTkdEuBqMi8pkZCzAO4d
y/2I1QarrRYL6odCIFdFgCI70bN4OR3XdmJly+gWthnc9KissA0PH/MRau3X9yJa
WBT/rDX4iT5jpEBEQheMsk1nj6MaK50vPibO/LohT374CWo8i7KAJp4zdvAscofm
39+xNcKY6QCSkCl61Ki6cyubUHq4pjGWQUxrEQRpk4lUXSNugzayooJ5kXHGnMsG
FnCOFlBCvnBFbyO2J4ZAVubA0tOT8YTpiQx96Lr/tpQML+4mYtDEwkfuq6KMlvka
En3wwiJEhNRO+C/6zmPc+eHowCLymYkEYnw6rmEAPP52nAqkh6eGQxIyRkogVe9T
tulVZGtF8C6oCOsY6BkSPl+zVzAhVt+YwYSlcHC1kJblbHFk3sdvYrchPGDs/mf3
GLFfk0lEW7deietapp2rpLctnK6U0cE8Ya+EFITDe5hEcprIqPRzYlB10q7vfMbb
YeLH26t3Z87X/0IT8gKgMnjnr+jiNI6jnir9SnZHHnK729N549rF0FpbwGZMKzZ/
rTtqnP2NeObXwWNbFGtwRK2h0NIYVR1enzCuLYBZyrfiJj9WczoC+h0Zxwa3/PCA
CCB/xuBPryEN110qR6/oGDbPcFtpdYIXF3rfmgQx2Req5mvhDyLoLqe6K9Qa8t30
Q7zR5xAXbXYLsR7/cm897iNB5HLPQzJjVPINJZWwBdphb8vxm31ufToKE+FzB0Zv
N7DN4QPpB5BfXBorU93ww1VHlq466IG18RqlaDHqW2NvAI4//ZYFUsCY8P0l+F+r
wLrFNTsUn2W87jRB/+OqapdY66kdN9oC4e2Wy/RrwyPIqu0ReEqICpTcmGsGijst
2McunPFVkLbSuF/d+ga2hJbaGjdmwW/UtCCIQp31n/mRgVMddokN1ReY/uX0VVX9
gXuUnQUHcvjEy8b4SKO1+raOFdrvzBZJe7Q436OFYJBX1tEOzqaok5IDwcjFdqFN
RDoHNR4S3mjYkvmhPRPhT826oq7hCtrwGCpEXqDrrZRaTHT9lkhsXe+WBFUvB3CT
jxi85VMK1uFSOUN4kkQYH+8RgDDCrwgMhB8Sn8GwAQ3Uzv+1UsafpZCvzIjApwlG
by9xxZ1NTqj4BEgrCw8u2Eg9N4ueGheKYb1kny9BJ/gDrIDJVNBIi9OnNphePYiH
Z5wYn2GscFFk4EmugUF6dtsLZBO/JEtYvkpRNLOfzXMdrGWOa4nHQcpZiWRGVFVg
O87qgY1IvAvBMxUEel3fK7hgcL3oxFDNZMMVCFBhI9A2DaVz/Vr3i5FhLtFRsYpv
9n+H1vT+QgrlU1FVPyGL2SMuzKtZe0HrVl4ww5hW50yKN58U1xhSayqH0CuayGHK
jhrgr8qFNh6jY8lszyZPFszwXpgrIXcuDmgMTEf5Ek05BhEvuJtO25rQiyn8wSQl
vA11ITdJU9WE/CvN2URAC9iCeIZ2ynOSizhBU75U0MqxJa9yEs8CdWOLsIpQg7wA
k+NeNXhpAVJV+5XKxxTTX6V7njVAbrHoQLeCyJ/WCoPq8ZcEiZj6RXWQT3U1BXZe
2HSsjVGPFSExS1iwK9BdOIRE0Z3W8D07RumgWbVws7ZQ8VuETQ/wOsOSA/pewcVL
d2JEK6XWUH2IpEj7XmsBdjgmPEc54KsSFD/MBXCL9deaSBGTMiivokvhsWyl3V62
Mn6mlfe6decbDxKXbAPvqH0J3rT4HJUJnrU9TyCzV70YPPvKLb7LuLGG7tNJAJtr
v6Tdx/Vi0LI4QXqrtwWDi9iym0xJClq9GurOzi45uWmZTBjE8DbcaeOjqqONGDXX
nY46zXxqKAfrkIpw85Srs67XJDZT/l7tHI4iYWhn8GalG0b3iUL0DOk2kucQwY66
15EpZz27KjFWuBwcUGWCT0Mtuwy2qhBrT5mh8hkBe2uivsROrEjdnaOMLdg9pLz3
tLWx7uEoGuCZCh4eoLSXHGAfvqFUfkPzjlOPu3SNUYlLfoYDntm2UQRGA96ua3B2
3rkJMFT41S+i8ncj9052bK7sVXDbCqh29pmdCZMDmakbYCYpq+g9GB6IEL16i7kV
EthjCG6EEJdujx0/Kty0bgf1oTbFnxktUtVy5r8ym0vSEYWXPteLLZ3pTYvymISA
mPJjD3cS2PqH3HSWGU3LVWX1Lte2/xB12dWQdCYFvp9jvVxKBYPrCtreRg4A6ek9
s1f+FM4nLHWHWY4ER1cgUgFLuqVw9Gz5VDappJpGo7/wZ3ZPYNvH4eLxtmSgDlFQ
Qz+1XADpwH0pnedWKSIhv0xOt+qCwxcHfMBuakDNEl/vKsRCdxmPdhAJ/YX0ByRC
2L9bG5Csfdv0E2+w1OIMPQzI2thSOExhtGq1UnZ7UW9F6f9CjaZWYNBwMUo7VulK
9s3LBEoPwAmGZLD2ME7M1u3Dcnc42J0dHIRMNgNR0uTIyqGeXhlGajpR9Gnka56y
lCH4EFwF/slzA2XTbvWZ6xhFFIjVGqwihXgmIRiG3YYa57c0vR+xFXlDjfVgAkGe
ofbEisPAfxtHzasd2DPSWpr2CJCDjfqgNNICQusGt0BeMkoInmKtlieEAGdf/k93
vKJfKPehRjDk3uQ80MO4Remung1ikoDOWbzf3JlZDMfzoka96iH9Jmuf0tjra9eQ
7dU7JEx521rOaotmx+a+qqseoM103t/tcV52U4vtqdZ38IujPnJ57bqCMIUmFo4u
rFmN3A3ts3MZ0S+Lj7puI8YcxG7O4zFXrypIlu75/eFcZg6p+3Zwk8OxbKGxqRs5
njp1VjStXHSi2p9xXYh0U8Ea1oVETHLxMlQAOgq5racQSYW9wGDXtmBvc8oBG2NE
UMq+Vb7N8JVyrEZSZbSF1LhrhjoDKubidp6iXUCpqCMDXLVU840evXyAjY7i9h65
62mNVmAcpaOonEBr+i76KJBMFztQ5nRy0agnzx3zD14ECk9APvG6OLbv2H1rGujO
T5efiVxrRcAZJPd5NR7AbxT9lrS+d3ArgUr7869p3VxKiKfiHbvzuhL+hbQGcAxu
9ujuPNuMQndg57F1SNgo4vQcMPpx5ZBVz/mdJGGYD6EPfHOTEV88+EbjBH0SfoQe
vgRCRISsOgZMyl5UlQ3luFTg7IVPjAUTyw0UjsDg6fRBxwmvQ6SQ5PL1pwW5Ri3E
RyyAKAl3lDRXcKUhFTjgE5YF4dUUqTGfOMx2QhaR19zQ03BBI4ct+Dfj6nwsdq4W
Ivw2D2h6sXK3wDSMHyf6/tPltQ7govKwFGp606Mewv6hBXV0MbOpAPF+O8gXOYzj
Ov30gSg+OSFzF2Z1i4fyzaQnLvANi4rx7UDVunhMpiW4RHCec281R/zvm7RMlktV
gsUVpIIL+RxQBJ1jHgKTF3ggFE1YgN5DzpyEV9Af2ldjJUQ1FoK489HyFFtoz2Kg
Bjm1JiFnQFf3XS4OoO1yfbuflo6OGuPZ++dW4XW9Q6XhRmTxhKiWrkr7rn0saSpK
EJwm1+C2J8azD3QAGEiu62VuyNS6npaq+FPJebwE2A+zdIRGjXEun7dNJPfVF7xo
2R0z3XugFPQpPbbgb+03gSUTaIXl1iuBWBwdoNCw9VEniBRmmAjN9+l5354hGnLm
Vau1NGpwDQhXTgLRCP2qcprNidRjioxpEQs77z7+0cfRvFp6xBLuIOmxj/57Mowm
rPIfQPF5Rv4w5SSDZrxDgb1ywlR+GmK7siYk9jnQoDWSt74YgzWRC7zjw6aoflZT
TC65iKw60mec8shAVRZBxi5xEOOwKOxbn7VrO7qJJfcWDatTpu0KZdBQfgtt0PiM
OweesPVorWDb1O3vb1XU4tZ+fhCZi5EYlupt95MNq0gp+d1S9T6BQJ6M0PDNjQyI
LwKXoXpsTJ2mqiLZwQRKNiMlAMltI0/SjF73hp7yvtmr5FN50tSo1jBATE6nafdP
a5dW7S3F2wwsrXckLFs+b3CKqbKxVcrjM63Y6IrwSh9n1Lxx4g+eN87uUxqxGKQa
HL3mnva9RpczKAs6sKYUOElq2lnN77oLgkMXW64wapCrCSEcN8PVnBFxRXAwUFbP
iJanwilYMKxPpnfrk58MUcRRXSid+dJkjDblrP+0dzsRkd+GkVsCc4GOoGJwQSlz
gO7Ew4NNGSlvJDWtXMd1nryN5yQ1nKGdwNerq9Pa/eabtll0Z1+NA7HS7ZkCo3I7
qV+HW7ikirRYYvOtIkgVl4BVjh4eFfsPwcxNCixGO7BOseTxcAv9bDjBC6/irpPa
P6J7WzNk5JOOjTumypYh/p5kEP1nuYbJ5kMRN3kK6QDsYSnlheZRf5wLWUvOs0rs
4oRhuUfuoIAhWkoy9VBjzvDBDTnY256lsS7jQ6lEctUFOlMZItrtwCsaa/wDni0T
G7m1PdDWI3g8ya/w9Bm3ihCTTXVyqpWAILJ76a2GXts0Xvg/wKU5ieg0cS+BAJZY
eOERR3SqAs0h9gQFKLFrpyl93dohBMAlwzxGVD1S8uWjCDTw/llmmt16+Nyt/V5Q
E8nXWScdZpUqoI2f3NK1Y+wLz9LSO4x7Jeyu8xXg3/1VCHBbbbtNuqeqV6bNSAmU
+ZB2/Ogmn+b+bWIYWgjEK2EKiH4W1SgeVdYDeOdlobN5THQF3hfMxwVSALLVNL81
LMa9CaA8gLaqghNqPRTIBvRF4SKr8OHdtQyWMzkrCjr27a9/u4UT5mX/0M2vPacp
m4epzUn2Jid8hmqKDGB/FzduJtXkFcAfKy8PmJ+dEqks/9Y2Iu5oNtzNqVJ3/Xhd
hjYTn1kyD72QcOH46mdf7lIZuhz6iJQvzcDxISJPRxRTG0Nflk4BQi/5kDbsCz/R
EO/hQ1cT1ar4krad3ejfEOCzk0LondI7qCptjn6ZHdEtSJgjHZe1+9rRiJC+abZU
8QwilP1JQl9eO1bQh7unwnyrNxT0I0VuSawW8OYBc6keEcJF7y+cDgrcMPDNXKqb
4+BOFze1Zd7z9xA4j/Kf3jMRNzKY9wBPmkK3eBRBKsgnuVEFSyyfKLLt+1lZn+tn
zBEvCdy7ti9qdqccyo6wEvFopaPJogTbDVyFXOusfcT1cgFJ1D2nTtAIyaOIiP0n
qQOfTyq9zvV1SLzYDExXVkRlatZdU9z7MyvtNJhibfnepuIi7vzZhYvtaetVhzvN
veA9SDzHBfti46A433Ltby18UlrFsINi5v4TKIsjk+YKFe45ixCJrTw56B+8qWba
evALgfrQNk1Bvqamtc8+tpSE7TLakv6KUTtdS2Ksbjo3DRoxD7w8BIQfS+A5cAcq
zSWRXRYMFgr5Lj1Idqh+6vfwMdcfQt0vK6vPvtmqH+dZMQOFjcyOHzkoDq8FBNZ0
fpQLwq2tvjcJCOEYkXVSLqJtOWNmH1WjvRG6ty5S+rNTgftkMeD1B1OXOna4GzIM
cyvjnWrDNRQWROdgJjLfJmkpHO80APbPO1yhmLqdvf46BqvPVwZLeJ/qWBhGa1M9
OjeQsVb5OOpeqN6OrQRzxZSMBbeiRy53SRPiilOQ5QeV5Gl7yX0kPYL9cxaw1Scf
XqtC6aIIJWKEHCqcmTNAb2wSSDeBTtl9M6Yi6dqp+x0pCPUujXpOBawcJvcGj+gp
dtCGIf1SI7ZmYyID1RWmFzyPx3qp23xB68NdrddfDY88XAnnY8aWsxh1xzJOo/6i
Iem53jo0qJWoKU3b1OQSODqxGgQ/eSQ1f3Cb7es08ne7zBMKCYB/+w76AfGZmfWu
Hvbwn2oXBHLSS8o25QdKyRoNAxOf0NZC8FhGqUg21E0sBPFWWFgLZ2E7ByUCjEcV
BfYIOHSeTrpO0AwsKHAG8E6gBdfCOlE2Hh/ynNzQGDxNhtj2n6mtON7ajbiuk+Lo
6jun7wb4que3XvgdzTo8mK+ppf17RG7YqznALZU1kJQeetS/Zv3gWDkRK/hWxDKp
6AUXKpBt0gE0zF8OjYeWNmIJ5Abxt4wJ8N/ZX9oMhDpE+ccseEaum3nqR667mFUw
t/Po5C9+GVHrUQ8yKpRX8eC+yFax1QzPlVJyRYzlJ/TcTXThHzbX7f4Dk+ds9dcw
AomRd5X7R3wuI1yQnSSBShIpvz4msiMeBh5RtadCPvCNoBksbvP6y2CGkJ1WgIMM
SHAwuOOY+ntCYhEX18iIErWk47gMQ89JbhoDpc7R2pQnIR757vS59FIUNxo97RER
/NGxOhRX4kcW8RqcgIY0V3sOqN6KzJZIjD9Q91VAvF+Ry0e0BEYqj4oJCv2hYKk4
zjf2kFAajWShzFbymZx+kSifNCno9EZdrgs+atZQ+MJp37GDClPdze7i9qZXjN1M
ZtVGi8b1dG05LAnXqAS/kTykWfO6V/x4gIhZeQYXbXLkGVJH5daXTT4nyXS771Sp
WLziGHI3JSNAX4EW3+ob03y3f+O/JDDCNqHT2+JjoqnnECf4HLVGrS8fW3Oiamp0
k6cf8X7MoQlnq8F64OzugsNAJWVBWmmeY/VrOv4oAxm+wtTx/lnU3fiXHlp2rAqI
D31BYWGhkkU8P33DuMp71yYAYeFt5MemkYo7aaSU61Az5NSCUcw7Rr/4nSk/asKX
RXOimXx6d8ND9IqbSOv9UyctSSwOe6lsIlNFSS+3Y0R0bde9Qi7LXQXAqerSgUrT
fc6YamlK4bTv8lTj2bi02Itj4FaTwV+ceffbK1c2afVsZ4d8s+/3HOej613pGBZ6
8nTuxg1RWQf+KOkI+OEwj5LrUJlXnDnx+YqIgTxFrQNLGuh7DbZXfKn5v4h1IhXD
7tbs4iVlxVAM4HyFwRZ6YqopPGfiTXyk+6m4Rxdr6Icog77vjLBFdx49Tesu7N4M
x1wodLW0dGBB+6rEK0aH5PnOco6I72uMc1fpeiIM7lI//WuP97SW18iXXx/HaAyS
emLiNRw8bXF897ghd5eX3d+AjyB8ewfctWJjVGd4Ye2A5N89m9NyLELAR42GnuPx
I52qoOzvQoj26gp278cZH0VVW3EbGX26iniRFjMGp5fUXEpJ2JtiM6KZFvk+EUX7
tNLjKq1vGSIhlwAikHVKa/otSWhvN2vpS59GocFOF+YteLhNRRtx/7HDdkyWInG0
glmnFaIHJ1SiSGXkZj8Txem2ueWsT/CTOlm9zRTU2dnF4XgMlGX4L6Pxc7+8zXfC
rHqU5l9JBQuxESf1wtoZF+K0JphNkCYdvr1UH74hKNsuEFjKsRVv6bwqB2Yo/rR1
HB0J1t8qIKHbLRWgvWDZxwE0Ls3mb4ujb6x7qZv2QxES5GmCXK3VHEGOMpsoC+Y5
1/MyfMkKHc3ToOWUmETAY+ZIlV3L9hFp3bC8J8dajOLn5ABSk1T9+txR63dU8NJq
vgZvqFLoFWG0vCGYeYy0f6igr7eh+MV2SXxrRbkxuKFeDCLY6FEqZgWcFwvIM2jT
i/QYozMx2thm05T5zjrYghFjw4YGcyIUpymI5YEFPAwWgr+sXq4EK2w3C6Ei0E78
pnMB3i7nhIcn4ykgfrWIU9rO1BdppSZNwTnDZhLu8epxT2vMlhpTACidGFRR7A3T
rkPsvxb0CwxyeBltYbDIPfKeHL4CxAeoc//V+XC7OzH5YrwybP6lY3PWjv4A8Ux/
v5AypMupgu7ps8OuXZPGr+qbbG7QyZzBssz3/EKR4ORCaJ9LTPKZMBMuNRV2mR/L
WoNPzOi0LYatBlKoMKzxOGIMPFlLjiCu2HfY+GFOKlUJb9dkxwV/e3X2A8JCJ5VA
y9XAi2SDU+rkhShrWwrdzrz0+2AS/BVWBlrxZuMg+DFv6QZNigOT3tISOfW7fgyN
PdIOXymilVem2Ekrh/0P+D9rqJrIs7nNKrRsfMUBNqWIRZCwNgBZDU6cBMyL4BOP
XGL25Vi1hqQZ/KAH5H7wUfgBaibwNiVU50YXQLrGb6d0tV2TEUvRduiu2/BmXjQK
liJX1sCu6/QJNWfxxMegP+nS6run7iPJXUTLJ9cHc+YKiP/Znj+5etkvys0cNOLJ
tf2NAD3aKKhg5KJ1FGccHieiYPUH05pFCZ1qETiYHcH1jGGtmSDaAhbPRR3vCYGa
18iArYRp8c3sYH8r+/imZtXzFH/ZklwgcrsW+l/tVvyinDCWVBfFi1zUrZblVedo
LxDVSiEv+1s4uTUlliuCoeiiLj7RGmxPDsdvXukgUmezc68BjfQf3odxTBRpRImC
FbWWCsVHpwWSfyyW18rYQ5iZhptgMe1kRWD4J5aD+yWk0KzXjbx+QPDK5AVIYWrX
EmnH5qqxwXZGtKg9AWlpZGhVX1J9gO9E1yfaLuFXh4EX0qJEljV8K1Ip849Vgk1+
NcbqgO4GA4smGWWq5Eode2byYGSn9Je9fOWI4/YEjPbOALJ/LXdKn9lpm4GDlTmG
IzrbERZ28M3EQrse2xL97mDBG5wAVFLEpEyE0Uo5l2BrntY81H3hLYoeS7s7z502
MoyJsRuzGlOi7ysf9FTH93TW6NK5YrrsQhFW5CMQ9/r4GtIREZZZxrVoBQnuMgUJ
wjH2/pAaMpvqW85oKwD9gkpkNg2RNlkKbtp7lQVCnyHbM2Ew7rjo1IyrdKhscx2w
j6GcF+9fqZioW/Bz2pk/72qOVY21kAy7hNXA/3D2P3Ba1DXd3mPU10J01f7ybC1l
kMQUk5NyHqhjMRv/uiLGv2WW/eoBVH+cs6NT8NSfgn8vuh0iz39IOdnQ6cYG2B7f
xS5CU6iJgbEdqi5aF2HWWRdjJq+8qNMphm7QNV2YpKm5UOEDEDyAeLutPgpCuCEs
0BcQZXY4D/bSiUTBKQ5njX5lPGaxaDhuJI8byt7HgEndVeeL0VIFNJ1NdHiCgUmg
n3L2OixC4P6qfEOt7Mh9GjNycmUJsPlAHervcv2DgvxmRiLWYSOTQwaQ6tXlZP/5
ASIOOZOtprDzOxA2aaVaqasDJNHunZpxN1yhRNDDUNS/zDIOiy/0FqPYRBh4ZJ+j
IqAldbRm2Jc2yhcEzuPeygaJtGb1ztU0w8ukQoSGcPYsX+p3CtSEiTwbNVTQTljZ
zAYvVxSQ9bdaTp1N+PNxPFp/gBcUSmragm6Rud+ZTLQo7LJiBQlzcJgVTjxE9B2h
Ya7vBaqNVdGdSHhuuDoMM9qckdDcwQchcu9MSPqOMy4PhLZ2oHH/2whzz2OVERUx
fKz7AWzegh5AdOaaqacwRdRNyGQoSbSPovDOppAMx/WaOVlUIMC9pKCmCs745QDg
y+OGtB+4nzoXeYJiW9AjIDtBeOHwOf2D0iOE+ifm1h5sqDC1MBOYD75DDCVgz8Ms
6XyW/LmZA6/7lQK0RGlRSOY545XQExz7iqv5Fyiu6MkYRXMH/LJwBz/IOQYByew+
7CKkyVYOZeVzi+69+7H2U6U1bixg09vzZOyY1V4OwcbcVFGlNbzXxe+ohWqrZiGW
fVSZ0LAiyw1QfWLAokQqD71bVqlrhODKNsBbRu7SdYSB+1A95xtm+ToA/Ogt69YP
pFpHtxRLX4IbHaf/KO7iQsnvxKVSDihF7K4cV93NvrMzQUWoY2k73wS43mGiyQo0
UC9m4u3NopxoYpJh9er1KRQkbsRyKZazQZWZO/sfO75ary0UrmVVbVOAh7P/uu8r
Hs5SUwEbBKRf60oGSOiql2A6TDxA0ZHZa1B9GT2ijnJ9mylMd7CoiIDKge+v6plx
ivo1P1aK3lbwLd2tNpv8ISOPfNtt7WF4e5TCDi9YmKdXR8GbMW1pDK+39tsqrZxt
hrmEd8WHCIe3rLQby/pArdrCm6IGDG5fVWNglI/yORWOA70NgIS6Fo+1/YrYw9Kw
ryGBfrYOAj5llXf44YHSuZjHL87nXg25/OBm+VzeLmBA6ZCVEfdGOclqpS8c3IVn
WA3Sg8Qq8QC48y/eyD1MMIC/zROw5A47r9t1UXFbpYk5cS4yV3yHoqRONB2ygRi6
16miI2T8Ld3f6uCCCmJwwy/GuFqDKTykok+khrqm9+bHJMJXTjvbHlFdigBn4NSt
ojMQ62oMlP3CAVvh9G4hQUE99hxpM0pUyRCI6cjvh6AlazhJCICxP6guB2jb34DJ
etSj6BJQ9mEQmGCYaNIqHi5kqFzWTm9hdNHOtRb0Ik7RX8VaEh7wLdPGb1d6vPdk
AQrY7Jee/BwHR+WI3KACn497l0cx1fCETdDxn7MX9S7rwmisvYLHudhQwHwg0E5g
f7m4vz/BkjZN8DfTtdVLWasQX87se7AJZTo8psp0G7ajN1j4l+u5dXGnp4OxnwUy
AVMI0VbhlFT2+Fw3vQeodo3nL5iz36uaeUGEtxA/BeauSVSSu3AIEkL52LyhiSLT
MBksMchQTnWwiwWdNXrQnoNDqFvwxOugF2XwU3fNrU6t2M4Ns0QOCI5xbH/XOTmy
Ye+SqXDnbUgi7B90i4bq1fiOAvQ9JexZzR/sjijo5CiGXKH7sosn+SC35y7DdRtz
8l8pYS8lGjuccDQqbahh4Ot9NIReajWO1zlm0XnE/BJf4etN7Ms72Mlj/R7l1AeW
GvGd5Qekbnc2TsVcHbFzvq738CROIs0/mNpzVHozK7vZSyZZfWpKoAWMJz2xXDni
URzViiGdRXSKQmo75FTqtP6Dvl2AGE2CGuZpDaMBaASIhkVYdmLyIMNB52ZC5L2q
HaQXgerQQeRPMBglTvCwZmRRt8N/Mi8kq3PraG0T4GQrmko1q4xKCQPHbWvzBg3D
6pnNLqeT2WgXF+ghXWat3cyaiOX4xJvAX/03aJO+gXu6k2GxR/9pbGTmSIAlPstm
h8xekfJdAgOxIQIU5Y1RWAKbZuA9WhbXOWfuKO95O+TkxzwObwof6/l01yth3zPr
nxMF8Hpd1j42V60gy8KygRHrDiNCdcpXDmrxW8MJcx3bKxwpQyqrPWrbTFdmRR2u
vlUJqZ0Hl47Cp6URt41HJ5xT37bknDmKzLL21nzCV+bEzyst3x7urIknyAq2/Bum
x4l7Y6Iv3yJIog9djf3ArQ11814cplhE/+GsEJTyOtDQT6FcY9W8cMZZTM+tktcH
WpSxKzk737afzS+tYmS0YzEOI4mDqFjdrzTcSU8AHqoj1FxME4WdpIOri0GdmHym
THz36ouspQIDlH/T45FnJEduT5WA7mHs8qI8gbRSc77Xtm5/wjfIJbpFq9t7eYT1
XGPVVwZbX2hI9A4BEs+/KDKW2iRpL/YbXgs9FvgyuVz6ldVpy/aW7/YYsi7kTd6U
8XHM22L9bjiqcZeuTk0SEy9KcbijOx6I3iZw3ptEnZEEb74VxJAdNBCYhcMT1YSi
cDuXk/QpdbEvwFkGxxV13tKKd5bRr3GwG+gvk+czAOLoZjZ37PrcQZVaA+I07x5L
xeXvf/SZIsZk7NV85LKZKHu+4BI2E/WBpDgm0eRQSe+b0TGCeM7rjcyjPCkGJZur
pW50deHRQoOO9R9aNdH39xDI77k5WbvVKg/h2SvaklEwbeznyIoXSl8wrugmZ/aD
f1CJZlxIVUUM5XCmslCo+Fw0AlTGUr+E2W3PY2y/5upj0HN1VjE3KfDJhyyB0hMz
9GIrUga+K5B4uHHMcjVLX5JHGiNLqyiuQgD/hvymMFR895BkphHB9MlKbk3IOa/d
bKPY8YmUNBH5dDIuqbFQdGDsNoYKfVLIo7DRiqB0/a28f3+hFADpcCRO9OjM2UJY
zWuJO0HN1esoldhFVzyhUXXJxOKxFkBrKebnC8IwU4ulPtYNGipsYtWcMQdgRQTW
W3bT1JBoqaimyXUvrZjEAaxtEc0OgsGgYTR/ofx9rmMrTRyjRbP329TajCpNhRJp
sDI6zm1/Tr2CnKG5w5mdajlw1INUJhgzPWLX+yyeFo6U61eVDW5TCi1xtO1BqyW3
/QcAABI43B5J0htcJ7qGIRgZ8WEiBMLI2cjA4CWxmIJrFJZbAfozWDLlzy1DPyT7
Uwip7U4xr4qvEYclmjpKFpfCla2WWdFwLTyH6ly7pr7UyrjvClxb0wtPQH4BBwD9
EdvD2jtXFFWVkmR3LuVrRQ2en2iVaOUzJ0j9o9tuoEYU7R3PDkOtNTIITk1zKv4m
lxVIoOnZsF4BrsBLOI95+HBTGM4aNSpWsu2NB3MstOWadK2JmpeAWX4nw9pA/1nk
pg4C7BJ9dAP8/F5yHB5hv5P7sS8/ABAoYroOrpxv9bdnomS6YuORRMbmfE/J2Ba5
rl6Pnd9JmzFDqRLnAZJFhaqt7AhwmobVmH5wuTLDMf9YItzqbWTAsmVRofr709DM
r8NA7QaHxlWQcV/LHiwqe1sTFlWw9ZNK7NNBu1BA0BRVFpEIMX5KERbbwWZlZfTK
fCB1yl9/+jozsPlOa+bMBxjxNPaePJeBukRU66/zkPEPZSMQfAhoCFymI+M2CO4K
YYGeQx1acGf64bQ10ltr1Ugr876J+9XjxnST2DCxpxReHKgjUNPDl5qkGXsZd2lG
GOJEfx8QQOuAsb4zRaHz1TZ9m/hGVLw3YRVtqj59RiTCuTfCsaz2Y0ww1uOn2rz6
5NphkXxzyryBt+vAPb4NT39Wn0RbhtTeFtX9n05/ZhUAP9Q4nEibz/jUa2j9bDua
AB0cw/NXJARsv/hDt1GJxxF7oD/p28qc2zGaxCBOYM/tnZoZusO+4pA11Py1yGEZ
aa3tRWgLXqdk56cidXYNc1TxFs0Lpu8/evumF3Dd/xHB7046Xm8rb0ahfthptAc3
hyyJHyUdsZGOo03fz0caZVn3oYn/aMfimUlR/3vGOVjVTOuGbZojmXMkG9FqP3Op
tJ3gGNhjbVvyZv/FekcRNVrGB8cbOk8ee0b45pifA//S2EeWFQlAL+Wb1bnpeEkm
KjJEOobFqW7l3n1VxneUElZPa/h5RWfdEa9kC1AkXnB7gcPE2UahGz33liRvvjM2
pwEPoqOKcc8dWMbJDtfJks+wxdMpWK39qJMF1SmCuyBR/gcsJE52qtHCzz26DIdy
ByQKAtGa9VsECrXxxh1ZtZxH41wNrdPgHyVamBjs+yXO6lbpuYowN7c2bStGAkkD
fGTy7RFKBcL/yTDRx2smqF6L/84rM5e9q1+ZANLVwAYC/QcKZEzgSgMcmHS1g+4i
cJ+S3c/wkKiTYq+IviEZa3HRHMEOR2euLkZeFQuYWvmLqwHgxY6WQL9Bfs4C2r9M
57kxKZt7Nr/XgNdFkWj6/pDMuhn0YBcv14EtfWZp45L2YkzBmqX8pVbOdtBrTuXW
wIBCdl5b7FlgdB69ExwfFfk+QPETweRxVOgWIO202xi9IaNaG61Cf8bNeqopSw1C
EVrw+ZFcw0jCt5jrTKBO48YHlEso5AZy9kTRW8xbnFgDoCMwgIkeB9E07QEwZb+l
UcOwJSRVOD2Y2cHHO68NyKEIJdjlW44xkM5V/152ORxC3VdkvQx+iZtD8TXuvml7
sIlRBUL8Fl3XCP+DZ7Ot2dX95xQB+VNyPUG4+Q+r3VJw65Md1Mw6HWtIXqq274YH
2LFs8qA0LepNPeIdgChsoKP3MOJNEAwzUy00BHqFPz36fKY8yU3up1ftpW3aAnH7
AKFx5NWYwHsS0/PznwCX9+9t4CQe8Mon05vpAtmFmAl6q173ntKiS4wyNQMh3zJN
br6MigpsORUaS1YumgGZvdmLG7R3ta7OxH6NwXSmgnoPgoAOYS1mmju21B6GGjqP
DHI9FCzrnevWqhPnSZ30+BchwouG/f8LfrkwvUkMsDRwYvg4ivKd0JuoghGBXW3k
xHmD2480+U1azevBa/4vj0YjscgEtMD/QjyrE1asWwGyhve6JyjYPcRn0llCU7IZ
hG//cnO61S6oqJLJjAkcCw5xRNC8Lc3Mtaw0lGSkPCn1W5I9kRUOYhIgGquMx5qk
WroNIrdU1mJ1MiSB0TNElEvLo35SN+EAfRImQco9AMuevTkiF7vZOR1rJmbHgNf8
2CCLpTOC5Kq5hbwhZeVDianDhCsUirM/og3WrESgHffIkN1yV7dk94Ie8NJbh4ps
fmf53zH2rGAeUePHgqmeKKU6hNj1nyaa3vsF5AbCfSdFqnjHRcEyDO3o5W8ujENo
HxOzWB/VzlQq0ioEWfoyu0a6q2vxxA6Ikk8BKAP+xpVKnE9ZcbOvW5O60p4ozr0j
Fq3CSABZ6C3AS3JywCQClhUSxcIoDgyEWnlHid/1cwsOvH25ABIYBdRT2IlnxmC4
ya8kU601rHRdzM40oOyDEYx1EKCvmQb+dIk1x+hlCuJ8sGJL8AsSimcXtUmNDBEu
y12FYbgrkUjyBNH068m6HfuFJ1TrxT0H7BGNWiRNnDT6BDOSqmXMI21kNkG3TPKR
NzK0rVs+DNVBNwDLVn7wl4yBXLyc+nyTqLM5QegUkkawxnzlTCuPv0xJYvdlHbqy
6mVoDSssxCxpUHEtGpOZ+O2yqaDBIEy9W324qmCJ+le7x6hlQ4vhgS4G4NBdhC6b
T76E6klxMqPhNJDQecYDq5HskdAp/vAqzyKJQdtBx/D/GyNGaNc8Z6yhWaA69Jk5
QjGGZ57HZeSG+AokaUR+ONngtcdnrA6KTpXQ703DHA7OMqqGChsBceM83rG9/Rp2
Fsc8RxdGw3fRAMJLkF3CLgczdbFMkDqCWwx0OF3jTkMlh8kuJfBDcoalUGZVBeZ/
2MedkxqrL/OJUSlrasm7VhiRLh8PL9HrImW3a2GKrpafQRQMsX0HGHOiPFAMNAhl
xdkCBQY4ZiTAjumfMoXkpMuoVxAyH0d0aVWu71j2JCyeSsTK577KNHHvXy4G6EW5
1zWwtj5LdhFtdANPyRRJkKcyUg/basbsyKsqfKwJpbEnzbtdtkXOnvexF/dQtO4W
dAx8Tj51cMpG0UUeKWSeOA+Mf1Nlj1zlYHwhQTddTlmQsIF3TkVIl71EvhVxhnr/
iwkmP56TmhsxY+uJgqe5fIllgCr0pN37fD7ZWq5wRNtevx2lbqa2iyzbDTrRIbW8
OpY1tsftFf8W+ytkMIayyEGK8wFZslBzKYsKioTEtYgZ8f0+0q7Ly5BAfokFvBql
W6pwSi56OE7Z2PyfL7J6hMmLT4D44V4F4+QrnB2jlgqN38B2IdI1k6Z+23Q9SPkD
FM+MTeQehb4gtbpa+E69MarPeUE73LtJ+02kNvFi6EbcmJhLgQfA9o8hKcoNH5u5
ghnqwFkIcTiNerUnXg3MQlL3naI/pt5IjOCVIH1HxPCihODHdqM9W/9RwMUruzne
mXPJuiQn1ZzblDYAbo1ED2WgUXV+v+PLPhaent45uXshoqw2UFhJz0E3AMxq4rYv
vfp1iMvGC6CEadrAvRWN9aDzW1nAI+8fg7LRZN3jaGocd72u1fVgMGrI4kOuHAvV
+WgnHUxz+1ZhfOijtz3tpLQzeslRB0D9H+oAXScxx4T4PYtibeWHyJIF+IPU5PGi
sma+JPWraN/H+t2lW0WJ2hQXF9nB55XodXVD9/bjWNS7e+c+VwJuuiFvdKVM7VST
nBSwaZoEsBnU5EaGFPqn4pV4DCvFET0nvmUOiUhcZr8H9Qxf8cqV5FEIXiY+idck
xaENE5hZpU2QPon8KE1AX3tlraY7n+MyLyfNkXwOHpjIphUSnqlFW4EHCV1rdY5i
+/DZzr4wLhPZGaiyNbml2+K1tJtHvs9e/33Bz+QjftUYrip+N4U8TQNvgnZaeZk6
Ih8Gq3IkEXnDnKqkoEy1F09acYROJZQ4wYV5LRqzMQRx7fT1RPTs6XWnpVY02+xT
XFf027ldISfNLgKaQI0LZVnEMLNCIdnbJwGXr8f1w42WhuxmsYTtO0y/RYj1zQVs
CHFL0h+Twj3K/JnxEfmlf1xU0kkaUW8z9rlwVt73zuj5h0VZjB3oIg2dQJiL7jDn
sXz0VNekrNM+kAWTVCZhkJClsDK673MpaF7OKTNOnrW1bW58uma58wGY5BwH+Yce
R4hkb4wjRLtK/E+6akqm0DjP1xG0kVWRYaWr+Lnlb/bdtaatjzn4MkGqlSKx03k5
w6tgIfJjOc1M3ohqrSeVr5bQ9u09dJkWnhfsFyg4x4/CUvERPlq80iEIrnIbLoWy
JTpbD54fcJCZ88guF0BjZYAp0Z3mCIP8omLOcaI7ep2s8XKZvbgeldqwefST59uW
egWQ1+vN1urn+XwEFter+Kf4Lq+FCY3mi7mLO2/buz98n6rxdt7Lm3QsQzbBmK54
UlwnI6i0FYMd/F3OexnwKVjFTTrnAdvc7NVSJGLu8P/kYbAH/PRew6VIeFKBjhD5
QAZBqzuBDvPWbk5mplb/spCnrJ0vDsX+z0aHteD+ZofFGnUnhPeWpPUttTnpqvwA
MAkiUdTtI1CUbs0qvqtuurHVCliKMZR+rbP7P6ogU60KeGpx2WfeQuETMaH4UkJh
cMv4ASRbhTap5jcKd6Q+r/6oWXy2QsN8hJesir1f6EaDU4/Jj/MG9sSesFSzzbO6
D0SPmrIrcL18QjJwVHJ//e+BNo8BKUF6UkeABHkBDOBxLtpPiL0NFvG809SyJTra
jPSyd6w/m0f//cUwN7UawSjKRsL1tsQlwg8oU8f+vAuApE2mwBXUBHeAMItdzRZV
nRrn4B4aQm9EOxlWXpSSqyW6Y/tnHogz6KrVmQlTdyYN80Y5A3gUZbPm2q9/h/qF
s3/i3OsgWeAx+XW+uaCTMCltYXypXaRSM/2EYmkN2J8pIEeTWDOvJglJ/T9nLDWu
nW/YzrFw9fFA5Dj5VDp14lfUmTdu2bNFhWopB2Wpo2TiL6fRkkTJsYE66l19/uuh
XfZrkiuLuQPEA6zZQht3KmsPVFVfq2dl39me7tr8TfTJzqyNacrOBWvwLzh+SQ6L
3g/69dqvH8D0oHGkkRkT1fcCPmiFqYCB1ThjiR0a/lofF/PiMAFcLNbmHdoZg9L6
GaLleUrDjsOXLPzaSAjMMUkmnPP3lWqhBPVdfvVjLBQGq/KsrQhwCRTXJ6NA10Us
nTiMzUu99Wiq38aD+eBRLUlG12dBfYwlQ0rQ2vM24jcEQOwO7eW3ZY6KdleoRxlR
za6AH8TVcXhlj+HuWNjNrSy1EwKWKoDugqIlcGs7hfeb3oKpPQtufuf2NhmZE7ES
A7MKG+SL/jvcM9I2CmIusajrR3TNJjjNMbjMRFIV0Bbi+rSd5eOhxc7Ds1ln3wuj
O2kYUOJnf8/08S6/UP5C0SmwnAd4cKwHz1Q+ImhnxTpmPT8Z0w0+oJGTqJtxahor
jA+uAtnU+p3wgsMevTfWUKf79UvxcCJ7dyVhAJMMoQAG+AT802AUy/Ebd8F1fQ4g
UP2wF9UD9HB/K5lk92djDhYAB9W+5IQ0LjjPvCmztwJwTS1BuhS7cN7P1Owx/Gya
HWP4+ZBvx22FLVwPOY+9gSHLPMefhfdCZyL2ajj+HARX7tTt/HuyyqxFg5lolj2V
67UKbG6iiosVA0irK5zHGYkVKEqX054nnvGGSc38r91+cJqzaHafNbju6s68TFEJ
jenAheFX/gpJVDegul75WmvUUhOzNaE8cu8hnLZVFOiCsWBVZg07RXHeHPEYCcF+
MXXKOmV90vy5TH5znaQMW7VL5yTvrqATz07TX29I+yUv3SK4ZUAEb9x7qdS/5azp
pFFkmECHfhGDoLC0/Q9jqgFhzlf85t9ffjA7PV52laPfhxxqSvW910FceCZdWOz4
/famlrZRuiScOls6n4LnbjHc0Ju+PACqOkTckIhQzCZe/7/7GEomeA7M8jNLaavC
uHwB3VWj0shhq1dzPyyqEDWNTlE+3pLuMgL0QHrAtLYoGGoAU/Zoi7bo2OYQB0qh
5phHRj9voqR1Uvo2/ilMOkTvSEknZEZDu2uAJc9UJ5Ji2X7p4Mq2HWIoOsKwmpu9
xEDxPvGnh564RbSbt+Q6V7kwL5DOpfgdm5WAQ3k+oHAbIplGgEdch/DQFUXSQo+l
F4ZbdR6zaH6ETtWpG0FLl35d/ZQVKL0hvIdygnNvOSQqzOJCUWBzu/agzBgmvYXS
VrRPMSTdkDqro65Iujo3Hb0qnn/9dcT52NlQsM2AgEw63N7+pdZQ2hkC4frJ/XF2
DpEUESBR/aTL2Qyd9PyCt6VYY8pxaNx4yhi20EphykgxiP5DTqcNxlNJhVK/b/nk
5X0NZrS7t1a1VYBfJu+9r2MuZmEjrW05Rp6+0C4piGsnYWkugnlPwLp1Y4XE5vbS
0f+OSvO0v/ZUaE9VLbxn6sYZ2xEE9PNuBmJEdUKunAYxkAl6z1ioBWPVP15Tv+7U
U0zVyVHfLIVgR+tdqr3Sy2YwBYpYGdL1iGZCfvHOEZsXdi/DDKU+wqOOA95aoVed
XnQRMtDaTZ3H1nrWBLadNrRptLJC/sTHFmfaCZPVsvkW36Cnaf56ZfImOy90GnOJ
bYER2dsQLYbx4lBfmD2GuqeOsnx25ddtFu+ndvkkNOF0qrVl0+rcnEo+jGghdQ7A
pUfesRRH2NO1Efry7qr6k6ja080Hk9XEX0AcEy0izk5z5MI/0CQA7luaDvWnGqXB
jJF0GWAzZc7qXqB0KSjcGJ1HYKZNrgH5DuiW4emSNmBU8DBN1UOVjXaximT+WF37
UMJjz1OZcBzW0Z3Oz26ts7BRTM0HqRAJyhhq9w1JUOYGSm9mtNyHQ2QOsv7Ggf4l
09jqA+xIEirze+s3GbpvS93uiCIQ2ZhmoW7yaOPsWTXa3BqLBatdwMSKoVxhsnh9
YfSsc4CXNAIlsfw9jpsH+lWm7b/Sf3j6X7r1MU2L+Kyb7GJPsJ7jk1fVLY/5TNk0
mLwwF74SjZy3oZncEcwbT1Z+BdkcfYW7rxrtzylN5eYRTP9YVW8Yy4cLhHDDybVo
feulOAMrxi74dC+17rVDy5AStaWibBcOqgA97XTf4wU/sxfWIlGI39XYYpBoNS0a
/s/BuHa/RSJ2LkuNJ4kiv8xD1ctitIP9Z0prMNOOzwwy+0QBfUo8iUg1JmXRP9ur
FqTiq7jOPKNIhDurw1EchW6BsZ+EnyOSF0OFFHDdrOWOVm3kuq9wcdJHxGsjm2d1
kuRvOoKiKZkb+5/GMwWcbnM4XQfsv6bNk1Qo5ZKUZFFwlv4n7izkNt1E2tJ1P+dV
xuMcru7BYFUv9pV8Z5R+2qzrxS5UfFEiusZSLv6zXkqDPg8RZpLegpFqHZ3wt8QS
Dzzi2eY6xgjc6Zcox70GZEfmVeg+SX/VCQlc64VsL4upAAYupGn7LRljUlHGookl
GSbP+Y2dgKpm0APGdZMnaXgi+eYMKmJKXwlB77YlcqDDDRXyI/bh6vTQMFSE6PKB
Ukug7jVGDqtQGaX8dQj0byMv7L4/2iMeW81BBRZTa+BGni/ztKUI7ZyPUZ8EAuJz
FpAXjFXRXQAgs8IEqOxU4EvejN7SOIloF6wWhxQ5B+8n7yDwKlMdB5rxEwkp6X25
VSdgZSj2jWwA1jwwEROUW6qNmCv65mr+QxrZVATwFIqyUP8XFAscTi2/DcM4SRIh
M90yhyXgMVPlfKrzJxUcd+36zYHaEUbRAu+U9weF/5vDYB9pGv2/ReluY1cp1oj/
l/xuTRFZaC+Mk5DpmiWw6PwxHiPiAamSqoq0ce6kHObD/cAGgcjN1mKOwTk5njX1
P8RJKKKeh5ZELceoS8ADky67NuPZ76UFDPo+2rghtw7aEXHnADV8jtCdbXI59eN2
G6i0XY7wajwzZmKH3lBi2Vk60Zlh54pXp/6mCqcc/33EUlYWgjt7ctIW+GOYwFVS
uEaYYdXPTP8UZ9sq29gclbhhMAEkx9cY1HaD4wqp8poCSBPY0NdoPVmVMzCTDLxi
ZL6NIoLcC0Jq+wsjiJLOfuR6L8+aQsPa4qDhsEMubLTdtW+rizMCTyWaiuLciTup
NOiklsq8yUscKtgOQLvoF+N+CBPPn3JkuMoPwWsk4UT3EwmQLmnWLsWjWw3AuS+t
h2/H/ilQdgDtNaUdSkqruh7Vjbj4qL6WXTniOxq6sRCExSG7Aph3s7rUPnv5jLMD
lIz0hzGQ1iLOkhTwWnxOcoUuTBzg/894bSGGY6lD2q53RJYSmirVbaD4O3f9jbtf
rhI8dUzIQITfqE8I2ZLtuYzjjNYZRisiGATFR2pr4/fv1AFnNqIKs7LUw36CWFmQ
EuyYqk+tZiFnmcD6kTm2NafjlEHREqzwUhIhEQxRSVo+NMn6pQjr0rb6rxdplGxQ
PbD43jdPj+M/DoNub8FAXvNxE6G/c3bi7Egn+xtULTn8A1vcBxWLyCa6CaVgdzxE
KOUa/N/cheWxgjtsuRpSUFzWNEk1d1pAIBu4ZXml/1Sa58po564L1OAqDu4gApvi
QrMCRCOR3ug+zC2paLnkj/nysAcRGaf/NzhD+itRtxQLLmx6GEMy0WLjmOLnWPNK
oitw4svICfptO1HmlZ4yxFu6ScNmqf0eDXqKzFO0AlJinHfeqFdE4uXqktNJI4fw
iE/Fp7jCZRl0k2UFSJVDGMcMg4py1vvlez72fsWxkjalBhPdPqecb/Hd6dOUI0d3
WUNk147XfgXGadQJCKo+FiL/R5RkrcnuHFY40yytdnQMUnFqvWqajt513m3PDC+t
ixI4mirp7bMfiyZdiW4bZhr66o5L78zRLhsSkGBabKxcS5uz4s1/BX/qT59EpcE0
1kLwm7OTiBDYyjK7zfMfgXrt6cQnZ2XwYzKng+5O1wwdIrMpR3qdcnrF/b2ZpNuw
+CpKtVvpKN+v6uVkVo4D5KVuOp5yVqe9zQEgkJOyWUHP4GIWjQXl1vcHZIvg489n
tqpRvZmOZFjgZwoXinL6p6HCr94AdCMskIXkTu9wC1xS2JMP3UDl539W6Z22nHeM
Jm/6AWbh5rIoI0zu2j7FNgbKOctnm4Zn5vNh5WFpmNKP5Abg9ocBvYLScuD9oKNV
0N5GZQdk7YkGGlSukHQoG2cR9X9pPynCH5vFHpc0IHSE+3lMcosmrvn6Yih0VaBc
KuydjjnpUVECh6e/dhy1nKfGfrD1X6hgTq0RG+p+Q2Hw158qfPVE5PkuVGxaXwX3
b+4NgUFqMl9znFeyNpc976aZaxMih+l8G79Sv+TaTg1IqWTxbq51TI6JZb4E7GEu
7kZYzS5FL719eVY0C43o78Ke7+tLVsEUItfRj0vsRTkCUlNElLmbLkzvUqKTXTz5
O4NRl9UNCXhytI+ctJ02A9l7eRzmFIohFHexOfZGEvPzykIkxJKloj1ofcUF9Kzl
bSECK72+5HDDSjG6gGccHL6eAbV9HN6IPTH5DfbYSSBddu39NkAp86RD7SUoekH1
BwsTTJX8x/m8M68wmKvJnaXfM8H8jxfAtiszrNHXJGONoyTKHkhbF+SWxgh0wa/i
yKDRiKT+70rDdSxDJhPuC2eM0CmKsNB4O5ilZmeqhvGVDjV45aVqeubVB69Ciwby
bmvNCnngMkHsLzocLaKLgLtSjsIiuyFoNaOy0inHkrSPALimfQPxxZg8/RqQTuwx
p0Zo7Hz6gaeI+pmIo+zWuAoIZqCbONXaKcbV0SOFJRYMjESyUNCERlWuAXfPHZsb
LjpaYE0HaIKdB3pn/ZDwYNiv5dJmD1k0kgHzcKYEKvq4KKzwgKJFQPj+CKKtmcUi
hIf7y7U7qwbxdkVZ6W2wGXJTFVtjAGdTiatyvykBYmYynWVImsMaVtzVEAW/Iz/Y
Huh28h4a7f4SaRyc92zxGaBULI59ZkrZyVPk0QnwMcXwwcBqsmBcLqJkDgZEYbEr
w8IvjE7WqiMKGqEe1uGnj4xnhUe09OXZsqyOWsExBXtQOru+CsGUeVeXwq6POtnd
B/vEr3Sirqk40ACqWengkqlI59LXZBS0Fi5xzzT/6rHH+RvoDBy2cOjJ6/Bm1APY
V0tQ6GBRzDoD7fZ1feBobBdI+VBHVqO9rcPR/ddOmHKjG+ivU0Te7gQopvfYdRdb
jYAaUddhxerdiOsU26VK77a3r0buKkEyp1JcnbrwIJWObVa2Y8OJYKkDsMLWtnku
jUlHNrqDHrPL67/BMrGLi6zG7rfF8OpFTNO9Hw8FgT7q+dD9vkcVJYuhfjUMd8Jb
UnS5N19+USZagxy01QJkZyAbVapI8ULVPYcgae4EaxITWCvgo2lzsIC5zVBPPAU4
+/xjBWmFTHjbgeRm2j6zg+z14vg31XrPmuNf4FDko4ypWQqQYMbiKV8TqFaQNqJw
LNGYLEXRNpgya15JrVhENIucOUFSXWYV+8X85dZfY1tMG3CtAhqJCQETy1HpumW2
RzsoE1E899V0sll/85O0nnZwvpXIBvfywUaq+2QLCeG2bpst+j5Aqe1LoV4WPulF
RQ/K6GoQelAG4X+eflCO1Sk0jSCk+C5NcJ5bqZb199yK0hQCs/SUdYaSzYyApV7c
E1n3YyU3ifOU1n0M4DApb4n0TbieUfePU9D+b3MqJ6sqhX4wC7VacGKztIyurgTP
7ERE4TTxlz3I6pQr45jrXYZyEY19D7r9rNzHgvky2MiL4dbyKecw+qhYCXcLtMKR
CxJ0a86zQIS6DIbJf2YFNfTU0QfMhNfoTfkbhfLCZklqLBFHIUO/YFEAJrGurFq6
ueGbmSqvABkmxgxS+fYkGxIoV4oJRpqhlauBnDwBKwBHBM/stTtlPo3RE4RgarRG
E3PT28WTUf/q2y8L0OVc29An7zTCvz3bvmAgoaG+4P9xdl6g8Dv0eSn6oE0sgACZ
ParXvdwvqCHgTiwEJ7wgd0knjwQa/L8tnr+uPF8W2QnBkwZ7LwGrUbyTyNKHaWOn
gsLWq6AtOVhrtRCTiVENlAidPW0AlJiXzZAylSNVaRkPdwyKUJbjjIGb4A6g/AdG
rW4QVZvdGAqlQ5i0IFmQJdMz1VRNIdPJDqSnlFLcavUfcMpDjYwgfcIyulwecTa4
yey8dxVOV7L6ASFfMlwYt4itN09JmzIOFfcqQ4yWsmyGjKq3WI70cHg9ksjjnGT8
sNSv6zQBI+ZmJ9EJ/++3D+VRnLdb6seW1xmHTWFLZ6f+G+/UHdtwV73jnw5qL9oS
bOe42jubxW1Zf0c5vj6AkNfdasIfgregx0gvclMocb289yUocNw18Zi3qPWvYrr1
85e5apwnIXwMTUYd4Jopc7onbNTLfHhbM3uSTuAZiyvNNT/LUcOwPsbjWArOnpH2
DYnwNojHJFyeOXde/q0PRqwvWNFLWoipOILJKOntho+7aVgrcbBaNGgKiQKs/Uli
f4UKZKrxmKC5lYms7RHcbfE2+P9B3shTyPl+3kiZg51nD2cW+NJkFVcfq+oJwBLa
8cOg3lqSsq9+N0xLolH3nZES1PzgYAyw1J01hLTIutUtNtIIC81njIBgGtX3pno3
2+bkKAuM8Mkrm9reMozICl/WIcfG24D+NiBvHCfI2LpwFw3WTHXBjbTVPxEPCMvS
qVT/Fy8DqsIHRa2cCeZp6jIu8LA/lOO31E2DfIOez12n9uAT9yEk4Umn5VBxL+dF
5Rx9fiDuL4tw77vBLLFGohSnm9+pMF0W/llDxmIqCXE8KPUYZ0Mme6JaRitYcVny
iLlaQ+h89q3BK5z20vDTBX/0XelZv8M/DlsW1kX4v8jI7ZC+LlgGkKqhxF8lg5DO
0RH2o/XkshjzXwzZLIzp8C6153NgtGz7E5+6ehkiYJ4XmasMiYeCXNm4U8ENyHSi
6Q776yNXpFEXkVAfQQ9jcApzes27vn4FVJhgzmDP2O6jesSzYAHlcPdY1tCGyb/T
U1nT2B7pZC5HAmQP0lrhBtG9hZGwOoOGP00nN5B9uBER19eMVM2cqBsh5kKOcdDv
0p+6cUorgZICbr35fWXCkE6fknCg7LpRIubOj5zA3ajrc3CsmuTxJrkoN0tUtcsR
qUw+bRW1Y9aA94yEAUzmu1CVEU87QKDOOVzpSAuGfSEpM7ZgvDXaTk6b6qp6609M
d680uFm0sGFwxr0y8QD9xLpdZ6ElHdXWcxxDUipqwY4LVg3JJQIjxYDEsO8u4INf
4i6+DCf10TElxgmrSoM1Ik8yKUiCxlxQBn3+pyNnxfaoi5cedFDeEhC4d/Y/upVa
XYVR9PaItdq8HhErjA0UHxLec4fFU0WSotPqF2Ee/Ld5vGunjlWqNhuHbKbDlNY8
6ubP5hBrGL5FjoMti9+BMOaj64cUOoK9aZBBbRi8QK5spXdZLCBea9svWn2PZUfV
ptE+k3c8+5W8/oF0tfijzUdwtrLh6hjG39cGDAUpAn6LrdkZDEN356B+cjSfrlcG
Al0Yu5/a+8qTISPPWss/l0PHZPOhP5/CGtCZ11rusejaflwDL+PK4EnwSME5S1Ci
YOrMGXmnVV0pnialU0rNSpBlyHvGmOJc5kHk8f3mC9erlh/zH3MFh+eLsEbk15Oc
VAeyphND6SJZsKqMnwP7oQFMiPkOz4fHpuwNMTn3PVXMXXpmDMuWOOVq5tbBd6yA
cEtW459y7NuuL+zH+og8VQBfwv4o9Q240tBtQZWO7fz5X83ID44xVQZFTp8/QUjK
kL7h9PUGPPfXtTy8Io+R/hyL3JZ7c6evf5dzfNM5cuDIbQGEg8L/T/3RljjA+/w6
Fclny3LctSPVY2DOU2+3WggCXFgWXat3bcMV0brIlmAHf8KghiL1dQo6FbfDaaEI
11g7/Z37n6QZGxHOHD/3WE/QRwnwQbqwd5gDMFRfFovMx/yufRYgwRPowHfKBKkx
yRn3JfDO9X53+FdBHco8/yHSodHwFu8j961gDJUPAsfn8q02AAGf9DI8HkdYq7Eq
tCwQuCIkMKTY5/73hWpyGlpRTYSi6KqiDCT+FMbi0ioK7k8uQkTVTy8pUXfSVFNy
3dg7ltcH3QKvUzY1xrG8dMGi8fHl4q7c1C97PRadnsU4TdP3IeXGGOo93dhKrQ7s
qqsVVI8QUbbvfrBnny8sVTkbsYZCF5ipT5xu6B+YVUhD6EC0fgxzUOnJeFvmZVmP
vBbnVeAzu0A+Sy5Ql2JkcANnszxkjW/618k0AXN9rOASrdX3F+G0ZSNLHZ1VdxuK
rqGLUiFnLAV/ipqHjAQ5oEx8rfQJZPawS+ZV9U2W9BuMG8/wpsb3b24ilI6/kOB6
PK7yO8Xefrpbr1k1rkOzdtzPZ/6YZeUWzv7jRK8ZNWOB3gaMFmfC1E2ApTM0cowu
WM07BGMc6XCMMQkP8nb6uMLmkrDiTdirrYj0sp9Q13iVnzEMozNdwQGq3RqSsaKj
YyqXlgigW2Yull/yuUbBx8x20rhmKN36/TL6FieBTIwllnfDoW1/6jccbWln88/i
bx434MNqcQm7WMUuHIKjNxlZE808vdjEr/SjqEZdgQUZeh9AAq5kzZmj9kWfCWO/
ARYU/fRnIqrfzwW2lSim514jLM0eCssH0mU5SbKYXTxduuASO7KHqQ8CM0zYvfCa
G4kcOIj1SiHfyezLSRBmLxo2e/4TIUjlRWQTKvO5JKNPn7GtzpLT8R+ECOU+v1de
EUFCk0FGigv6c7jbZsFIJ6x70a5bPdOUk/cO+8WJFiATH/LVRxNl+GK5IKfFJmuh
xEFfcYXEkax87x1+vVFi55z6GYdJt0Jl9K5TBdRC64+Sm3zyfu7HGbIumdMt1LYA
rU8wzB4k0vYf/TY234JLgrxfmu6FyDz1mM/JkyyIyZnrpOdKhYElHkk0PlFXuBCz
0p+czxeTCCuBPLiVDWqHPYBvEfm9WyTSzOHQQ/VOEWOgiSWexNK5/Qv/eiMniRVS
zgJZMYJ7oQt1vSH/1cPonTpaeXjxxt91VjlG2HS9r+fBDErTuLFeayS3cmXfhUyP
LOaRiulUOkz+Dlu2jeWeSSbErlUUsu3vDtdGGxS3vWeivayHDcCkTPnRZCXkvIO5
WOnpL7oBgDtKtSx8FbOiiBAyOsy6T8dRx6i/dLynjCBKyATPkV2JGkuPEk7lIqAE
Z+BJtdwVBYyFTqyhiuiv8nufv9zs+9Y+XX9dcq9YtOlVhDqr8GDxIYzjkmjNTOcw
Cr1u9GD0tN5xn6TM6Vn+MvfbG4vw/OQgKuMyHtCM4w5PcrgiLhtMhwKkktujDZmY
an8UujNUtcw+JEr3zHP3udQ/ME1dYAnLRHsxtjgRqFP2QPtEqi9z0MRaFb4gHgN6
qG+2q5xyN11yBI7H5g455tAEhRSIutnP/eAsTWm/vgA4oxbKyls3HUt9K8OCvxxB
XpMn8OSO1wX/Jx5hS3s1wnvUBv9VDGzYiugPbaKEQ5xSdzoxLcK5NTLBXtE0ecEP
tR+s//sYhqCR+Ug3xaEviqDNsQZTPWHTXuQ3VOY4878mulLEyo20OzyQxcNJAJ3O
i1JDwNLTW1KytGEfrRiPoJmefr8Ygdt4GL72Y0EA/ooRdK2gC+PKrkQJDKQfxqUP
1zMWwVq34NE/XU/bhZny2FkFc+PAk1UXvKzOMPRF1si1kusf7kDOrp5FCPtlvNKo
hGJgMjoC5BsyOLgy/jW6uO+wAx/10OO3+SNtgl01khSOrJsCSZTPWoH7dtWoIOMf
5ZIFcD/X0wFWty8sTT8R7IRkAn5X9NHRtIhQiD+ElSnMl5ucc9vdxiBUv3WIQUWj
j8O4iRNMK84kywUNvX76it8LwQ57VtG52a47vJYSr9mXW1SobnJi3ZsvM2FGPKGh
gYsBNhnaOxqU7HsHf/TnN9obR34bY/29jwGE8x+njsxL0f/VOZDRlKfICN76yQsJ
QlQU1GYsWX3lV0RyfO04fqWtdAksRg1s+D7MyPztFVnzjYFFisJMAQ2eP+8iOjGd
MAXxcY8llYchp5gmDw+KAA0IS2mroTGRD0E4CdD9n9nDerdTotSVq7YYL9x8JKuU
MKThG6rK/ftg/zehyio324pQfLMax7jawgJz72grX72UCs5BEyl6PAE95Cc1wGuM
f7g/di1Td1RbMtKQlGVGYnCcRFqaggk76XM7II2pAvgivGIpzyjGYDF1Xhzw9F5s
eHXYcyZ+RnipYVxA1c0/BD7uLRWX/QTdASTt/Joxh8Scaew06+ExdcFwkhf+xv38
ZNBM/YbKC784YrRGSMzoxxbFYB6um4JGQHzCITFnxCmUEE6iyaS0KNOONx7gPYqc
sHQYEnIxGniLf1SDp/Xk++r7ddloc9E3hqPbxGjFKWJrgc5F/QTmr2q1rdo4DykU
QBhyH5JRutizCXB9xanm3GNMRct5mcpBctDtnB4g4Rms+9BBPyYERvAOAA0r0/m/
eP0Ta01iI4dYeAyLVDSy4+0+XI0M4C/bUW1z1a3+sKGR/S0wjHxpg8ANHz032H8D
25yArzH/6wRuvr0v98gSMsLUMRxw0lFFOAn/heUkXEv+Fp2YfmG3WPmPJnGuHref
Q1JgSmKppoENlzyqiBxb0fFmhZrvwXpgRf7LAUoQIc9TNuUxAblnc052164AYisr
FvUQYgkbblr7rWf+Jt/PfcRWv/8dTqE9eXYzNeMfN7/Hsgnj93j5yPaePzbAe8gH
xN9w8eQKwqQBtEfI2TPmXw1LE4t3rqJjgxAcaiZ0UAqYzl7190yRMAQ4QBhlrkfh
7o0P89SIlRp7zrLi4Y0iBWm3xBz2vCbQ6ZEZhOdUD6lW4KNBuNlMyakwizoDbsbK
jzE3Ocur72KlTmDxy2uBeUuAyeYJ33BFbcLVCtoF1yoCLg3As/Jx/NFVGPPHTDdp
EtULTP9JrWvW9Q2sTYVpFtusJ6lEsAJtPk1fpc1Td/K91RrVa4570Yc6ZbZ3vpCv
ote0Wl5ilS5SDPmEKwj1MJn9thYH03Nql+uaIoDXD6v4yVn1VpmUfq9giIGNVLIe
MWxnCbzD+x1ZHAwr3BF4VVBgS0wZRgZ7S7276jptM95tN3eRZlXtLJ+ZQ6CeopQc
FJeFKEUXHbnGmdhX1T484Juar5qtdY9QrJTJ5l96T++YGhDC8U8EWQQkpsRGIGL6
QYGe1mmovoOvs3v/d9zKxQHUG098/9POqTBaXCSoUhnx49rUHadYLSGWChr+OWvj
lljqrcg3OduNS1Y4C7JsMl5Zei3GJZXljQ46JLmrbpimJ9uy3Eu/tVca3ZWDFVXp
V6AzvKH7944Lh94c97tIDwhuZjKD7XRHGVnx0OILD62rd7SBIi3GtYFStXhVQx0G
oZiY/cszlwCzLacK3LB+MtIMLjBMt2uuJy+FwVKJxgHddYbNK4r0EHi7NKuRco+C
NMwUFuHryUTxc/G71eKB9WBXOabKLIxGslJqOuGg3YeUbknkOTWsgh2ooFvsUE0h
L8bU3NLd5PAOCDq2dTEu6PvoAEHNwaoRBhtaNWl9KYOjsib6PXZ3DT42LTt5UNOU
o07OmM9oGYnfpdOa3gIqEOlb3mUv2DCCyFpYnwd9Gbz8ISHTE0X88BK4RNpDpCgD
+dKSLnp57s3lt0opCNiSH/GtzV1Jd9ZRW8tTyW5ib8LbWsIDEQr43Sbk8acc3aZX
N0KAA3REzch+XGcl/r44LMOSTgU6yjHmh1mLrISGkkJrzyPyQsGAUTm29LFy8/VQ
7Dj+JSNRuuFoOwDsMKpQacZB2pSGpGNbPpggafwHjzmeUhyvlUPXt1cCMVYI2S+S
if2nimZSL16JkOTLfaxybkj+ZiQiJ1WtLS1FxFRRKphPEPCk/J7+OZ6IPJVezmqf
nYthzXWpD4bpcjKj7ZFgBSBVFRiCQX5xLincpZjFcUDTrzlhKMt4C47g/5TYgDdl
2yPqWjjO1PF+osemzehIFpifjq03PKFLVjOGW+oXmw4oskTPpeEPCBnn9s3E9i8I
AMeiaff+K6Qd2C0S+D4XFPdUjmp+y9g6CF0//HJwiLifK9An92ji2NwP1s+W4ZSj
cN1kXXxOydGoSejxBkrqB+69xk0GIOjYQX9bKFFCdcsIrSUDrLLrDXp1wHhjn0k8
iiiZ2DgfEfwKwz9Sxv0pC+mjos7DItfMFeZlArO9/dds3+N0X43p1f8avQ5kkCeh
WsBalrFtQw0v3RfdAlwLdjwigeNlKSaL+EVihKDjEJ7u6Y6Gw0tsKZjGQXguleQP
EFmqAHa6rFE2M2cf94wgO9XtWRFrJSstHx7xgNiI/5f9FK/943B2E23rPdRtJvGS
G3QcFKJ1vp1J8oGzSBf7sZE6A2wlHP/sjSOqzIylkVXXVIRwqPcJbjhITTpsSJy1
M3dKYtdOQBxh6IvNzLZRimo2P6zOc2Go5TDg4SbfTaa8iyZTvmI25dmr0HXEDax8
PcuuT5JRILLaD+TsBICm6njnyBoJuxLYHuASCVoiOpQQRUep/9xeRqRZfyKL1grg
wZqVb96byiTwJyeEBfKQARwQ6nhcyLJdcML+EeN211pvtmet0l1GF8/kBjHV4To1
LkyxCH5HW5s3gNSv+MuL0QfV+7XnWm0bE3bszQr0K7y+hpdRQtprd9LL/xbLeWA+
aNkGCma6Jd5NSFuZs+viPyLptRf94Sd2BDZ7ODEEpycTbMaY0cT0LWiOOCtCZ94s
5ghmxqhFtK3QwonbVeFg+J0Et8T9/lcLjOHdJeNONpOAN5K6VPaqlmLvA59AEPZ2
19WkhHYqGdUqpRNyeGtVs6Lte0JWdPeqMaySf6v4EVqRbJ+kv+6wYnToqT4xSob/
zSybT3g5cH4CUfyNpGC3EMW99KvYxgsQIyRDUjg87d1qGbjwg7GiUKrFqbExP4B0
c/kdwUbV/v6+wKfq73/whtSOE/ONBaDQVo1JbLRHOtXFOyrD744kpkNDV44EUShk
qcubqDP5PD1J8fftXfMOqvT6XZICHQUYi0fWbSQGQo7RnWivzQiaUAyaxqFVIM6b
J8wD6gK/BycLFenIFb/ukyjhk/5AxO11EDaR5hIt7we/h3RogIuOfaRPPdxuLjht
k+xp43oi4wcN1yZVTmX7KGIXaP4MhuUGxcDNDvq8SZUYPL5LdG9BIxlWxadiJR4D
kU/zT1S8Fx4+HRnMKBMey/Sp4PXiOVhLI48E3048tuiQFlNJbgqE/T1omfbZz7R9
slR0J7g4XhSHjlel5tlIIfleHI+LW64kcJL7YyOwop79tIDUqh8kbwGbSsrRci2x
9t/5THMx3LnE4Zu4DQ6joL+gr8dMCiXPfUS5tE3rye1+7UDci+/eCyOi/cKSz9gc
ayypkYxDUEuK7EMGflp78WUigUkQTc4QRKHesaX1TrO807O/v0L33D45GNlwscdN
G2RRcB22/i5NTvma2tc6Hb7oJzdxXcQJVmEBUugcaFFzkBBqnBDjfQWxtbBmjUs+
32JzudxrT+bLUpxNVZ3Fieh32wO154pGbj/DxQYF9BRabbJjv0GmNpz5ZyUWhA/J
a66B99i7+nZ9lz3auX8l4Ezby7UOgD1Jus1hoABNT8O4NGZOebtDgGdb7hHlu/0P
8n4o1qySZTLRM21xvu8r7doaoi2WkXs2YVNu4v9aRu66IScnaa9scPYQuBMUQRn7
Yv0DngNL0aY0WCdFhWyX/36TEX2pBvWqQ/MFo9pyDvrDrYf0a6V4emwGcvxZjTdp
5IxpBq4jNNLAIvQvHdgH/HAMwl+gP0sRNIjKqNgqT93XIyYk+960zKxqZ/ZTI72C
LjfJ/TX+Bwj6w1CYNyDt4T/ZOKPhAE9+LNBJvmigk5/I/38O8eSXif0738EDDXa3
6zec8ITDgnaVjVw71aZVbJCyPLXyVtJBv5HqLRvm6gOKBJewZ/flmxJ1KX/pQ2jj
GZMMMuQOADWD9OrjM2kcVtg4cbBi1wChL+/V9N8Fyf0mHGFE/b33CeRcE8fhTWD/
8H8GUcY3qYp9jgsi9awdfPxlQvj4Nqv1VpKZwXYKzcdRMJwqMgdQ/ZBqX1Xk7lkL
TTUC1X4v18oIAZbx+Pcimd/gQsjbb7rho2isqgmlg/4UARJzS6/ojKWzhnvrFQBb
IfGemnt29MXXiEwG2/YmbmgRdrUUlWDuq3qxXMK1NtbtoWMq9xVgAY9ZyVCa+hJe
MVWWDA+Mlb08G+HU4/1IzHBMRVyhDIX+kACChrVENmxP+2YH8V6TluJKPKXgVFTv
pXK4PtA/LwnyN5luuHytIdfWOr1vH1CGVT9toUeYjuBdBENkC1prgbvk7KZzef16
vnqhiHqSPYCDuKGu2x6pcuU0eNnNUSs/GV+9Q1qm5+hA0n+z8OQb8sT0K9mbFmBg
T3wl5pkGfw4/G8MPIJ9C4dLDAym16EWC36+d9fsyPZsPdzLwZLr6FnwLf84/oM/y
wJ6Aca/WkxWfEeLHPazUKU3/h7U+qjK3xyW5LycKxAjSMq+tbnXqi86EAhsPvCJ7
IKkALEOYmAFBD9SRHu5nc7wfBdVxL978Yd5xDIe3qDhCZUti3aQ+Pmbhv2nx56dF
qCPAJ70BnGS7AXkPr8g8BvEeakYlUFLRdhYQuf/0+KLlz6QxFs4tW8UjpaTD5zKP
aONg5lYX8dq1YQtWO6EQhoHAzVevCFjJYiD43+Rx5p60GMbdu/+JIu9/Bn6qCLND
bjZaqinYkD116esuf7zsDy7rYYgSwFhqGI2v/AaGdbvJ/G1KF64bRD9FxXLytFUj
dsxhmI8sPkgr3NttuvQzOU92RK7K0toVOCE4WtB0fmbiALvd4EcyaVtkfQJRn8pt
JTRXnOdXtYyhU12mHbSXmBHrpmHfac53QyUMaIXrVNEJWuwLLQioIcPyOzJu+idU
kWdyWlMMVSjRTV5U9aOGBix6not2Kg0hlbGkq0dmfrFAmcjxEYSll2FwBTM2gi77
4k5lqvkbP4WqgKbWSy9SLCVKmbWfhidl44uBP9w2nQoOIGnnP2qUpH2wEolqL/Ma
URvpGQFTi8InIHO8tT0tkyEGLG/vM6x01NV44Orly8OvzEifVAqbPHIoaM0sXdxw
7a84s6QqAJz5qVLmaPyvGJ9U27nmShrCiXBC20WVJr1cR+/kRf7VPmsFIplgbqAl
OgjbYn3vVjIpDtQnR8dJL5Xs70uC7E+Qa3LutzJh/rbGenXxW2X+j1+O3IQezzyV
KEyDnGNHJQS2cQl+9sBbGkZw+rykEGZ1m7Cspoo130NKXWHeol5mm/hhS2X5QIiI
LRMTnD6dYqVrsxk+YIurwgsy6bQcGj/18Mpc/yeCeOva9F3UsyXpP7OmIAW631YZ
REC+TrBy9V/P6os2YEK4o3LpmbJJbTmnh6ena6GaaHtRDfgMPiV+HLXbCWySe7bY
75jyySAtiPokbAMMFFRNYQL9wWIFUHiDIv0PmbJ1zxw5DkTdwmndZmojkjHA26S+
nBe0EtIlD+fRxpjcLWy95kKIsxZ6beomaZD7SUrlHdl8W/GfMdeYrZZZ350N29zo
3TyUogUwTO4w+Wbp9VN9byRgzmEb74wdHAPir6AnYzpFpkYzgK6AaKiAto92a/JV
3YuNuZVbi8rcrhlCiy0XYGEoBfVRJoNJeNFuJsRl+NiQILyVy0MUMOAwL615yJsM
1XvAkRVwkEGUOiS9vpHlgQ5bzYeFvUUecQTAIi5dkeTbcm0RqsUvFNh5G3rqJ2ol
X7x4kR+iCfgCBThhCdOubvdsfao6+6UsQkgmo4IRVkq+9N6c6N1oLewkuCIj8jSC
7xYbUzRCmq3FtawKWrzz8YkOAaQPtmilyrTydeiFjG/2e0Hlp2zE1aekOxMBizwQ
/iHxGU1YprtO6psCjZ2WH2fCQ1us9ErGimT1D/Cjqdz2er2+MPotDVdxkvpdxx4/
ycEbmMR+EAvnwrzASBRypQ3G6/37MiXiFHMtEp9qWIaK1V4cnGsSt/CGs7rwEaJ6
aoZg/VZZFDspDtCgX83qk2ikC0VGtpjezbsCSONJp7GBFnMuAlpjTXC5jaDb3cOJ
RQP5NcC/YCp/ICjHgQnSOLLjH37hnPcLtq96+iCJL0W9enPyntZaihP4lQqcV8Sg
uWGKMS6cywRAPoAHR78UPRFC1IC6L2+CgzVaQzQo1LSlSQ5kKI6tW+yCIK3U5jL4
84o+lvorfkyflkGEuSHTzyKev91dzO9+alqQTw60DpX7X/elhUKnDriHi+DfDo4w
Ow1s6tuBVtDRPjMdF+nVaDKEIDxmFKpJQyzGurlc5Zqu2XrFOZTXm0EDYRhq7mYY
osxB+9gX67pgdZiPE8Ne26j+DNXh3ELYAAc7NB7YIyJoJeMfZg6B8d47wkw2alEo
j8m5CYSg5xmXh/k2CcCXTjT8ho2Sitk0rR8Pfo5GTECEwKqiXUDh9unNa20b/k0o
TK26i2VtNvgMgX2xTRNVbKEklVSnNNpx66WwmL6SHbvh4XE0e1OAPRUDNeVaqgaI
a6hOSM+Y1wyaJnNFx/qFY1j0nFodkVCpmbCCJuPdRRX0j77hvfJBANr8gg+tdv/s
vWiGzbYqHRN6CoaNU3xTg/NKHI0GLkIzQnI50xNLzspCmYdjRCPcUk0mtulL6sg0
lszaROMCOx7H9GFrmgVu94k7dQ/9auUlEgkttn2j5GbCaq3lItePVcT8q1n55A/7
J3SrL3ozKzFr68tr+Kyy6HaBuMaafE6o4VQEUzw1ALJfrbl+1v3d/i0qfv5JfE2G
iXiOt//LVnDKkitzfK0VHaHjMVZMa4MwtBIbjWhkHxMNEhO+dImOYWDaKl3cfNKa
JQ5eKvH3UYpC3ZrSQ0P1N+cxftRG4Tzu7HSOrZOBnoIXhJRAh1Z3hblJo4nv/zm2
Cqe8/WT2LiU7CxWYGEbsnEcrAKIFdbq5WI4n8Py3R78nVvi7AXSCb7lPVoSKL+Je
334/Rl9ab+5J7bc5mszGTeI8Tchrfhc1Rq6CY/WHfok8zLjeqckzGnA5TJ4rOfJl
BcKyLuMs8ZckPXmTxrczE8e38DfSaYk48pQnCnw1xSHQlIRzG1y6Ra6/QyMQh8QK
QKC1oXEskPuO99xromhQZWI1dUpaCaWUtVnkWz91nEmFb34ELXm//nmZrPzLPIVP
7Nrxb1p+PIDkCohaGPOruUgdWawxg43NEQxtGDvCGRXyArlwy8ACD+qKogKo3thk
e9OVT6pYSl/KDPrWz1EqX/dN+adheh5Xv8bU7T0Q+VPWtCLaIicp+atajXDgu0yA
sLwMcoM9TtdPaPbandAi0VocfUhfiXYpQ15OEMdEvmjUr05cIs1qjuozjenM7+Bp
uAcxFuy4rtVEzOV8JrEkkXWFQcPVRX5VgNc4nhtmpZ3F+IZjF0IwOS+coLcIam1+
s/lXRJYkyNwY985P3vQf/z0BzQIN7Nup/4NrSSKfHAh5sSAaL0K/Q6lws/szqSaC
Y7txeOOXXGcAtqcNmNMeWXvSmVg0LopV3WTBwSc312f3HwtDTMZPo0+QYNBdxULW
Ts+Lhup1353XsR0fE1nsJ1hdsgwAvc8xAvQ/nuGnmbQh/Pq1bQyNC51toBFDlJ29
/eVLpCB5IstEj5AyFEhayfVTIOvFyTu9e7H2j+XWfSPWsZHMveYy6BuAiGBFAZ3j
TUAmzzhbgJiCFRjgQcwXP4YNz6fiHiuCiq8QavHxPvenEpd8Ou9TJovf1lW9Y4ZJ
yfcrEs42teNX4HLpCJ1R2WNi/9t8/KfgNkWpWTtbBabfe5VVxwtajhP/vWpqubwT
qwDqwVr5k2jY7FELqZtEMoC8skUIT70wQqu5dA0UIi5CnCICEvZ6HIh20TCC954G
myRJibNOmDbDK6EG52BSl7d+uWdvEkcLQCNNKSjhBM52eS81cGwAXZv/uqgDaoE6
dW3CMlh/pKmg11fUxGRIWEhiDy/Ty68ERkD32OuAFs5zcilPaSVk/8Xpvpl6aLDN
6E2sQW9+ZIoDg2RcJrwdClbrDOk/H1JmBTnNwrqZSjW7/jGkhuEQ0lTh6rV8I7of
+3Y5hngiiOzvTat8BPK7ZlGpq9J6G1XJxoklpVhKdcGGHf8Ey32h936rlOyarBCM
QzMh/BAEzWuaEJFAN3Prb2kwGKNcn2Xsh8YH6JUSHEO5xC7ashrEKRog0N/53F5h
8b5Z/8gykLb+MkW9nBdnHtHeM82IaPmXhd4Y90E/KafRpyXc8F4O/PkA4iFZ+ilY
v70lZKHKUA33p4RimB/yjOkpCXrWj9//UHDmS4fget2bNgz2RG0ZPKbKT7gVSlRY
KdRRdihN/1+1ULeW7SabB1vgcVLB6SmBn8ArKQWRqxCr7EjyZ+RZciFApKOu0WsF
KGOv0t2Zr0m3Z3iFlKf/lND1FBb/99Xn/Fe1GHKdrb2jlRyaMtTsQkjUeB+Bw3BA
Gh6c3nNC4JoLx1NYzpu+aS+wuS7zVXTP8JQy7PKH8xZA1hevkSLGm/sPau/W4sQ0
uASfjkYebD52F6ip8KEUS24fcTP0oQtKUVehN3cWkeonvibh9gUaxE/eGe1dqk1Y
8ND868ArVc0RXTW58GXCjPJt3U3v/C53mcLn7plKvkLXf7FGsrsZGL9WqP3jAAUR
GbodIHUtdqcSctwkhqAy7t04exaVshmyOrprks9Go+CO/W/5oL3EvTquK2PktSqa
nn4tgHZ6gzLq3F1N1/5fWPcQ5qjev+MzJLDMJNijsVcVT08cRU3wHsDhpOhvff/9
sYv7gguUa66I5blcGVk9xsQIxnL4yNYDw3MAs6L3kmBVy0cVdLebID5+f6uphKdA
9s57VdeATHcPOx8UY389l4V8Q5JTr4Pc6vwDc5/y/3IRl+SH70pcfWsceQbP001N
YD5+UI9XxHXoaNxMHg3iHSKFJ669GG5pcB004Ax5QkOG6xBkVW0fnhpSd8qcfanx
qBOChmOS6PymB3xIo7HhDBNmRq6hy2AZBBi/fwiGyF+LdqPzrl+VG9yk4fMhhnu1
BinoUtgzO1ODrEWf8SWjjRY2EtryDR1XCS/NT/SFJ8Tf51EEZLAwrSuVZzautHuW
u92Ei8/rRsLcLBbxWJillCtiO29hyV89cZJ3afBldbENtheKjixyew9RV3VEPdUs
xst6+MXNSnmVtzpe+wwxxtW8SYo3Uw4j6ch2kn1MZ1zrS/hD3hmcTUblhxaVPMv8
blKgB5Y216DV5w1aTHoxI2LQqyTlRlX/W9CX1zXrtiX7sLC7zG6rJgJFPuF7p0K5
c1wkhT2hBJErKX3rSnGbSH/nJMXmXWupJoUZxjxuBSPZpQMPq4h7swiJc2jkSHeS
omtTirUL70Bf3DJS5sPImaHqHSzFpKjFirrPvbdqI+r3w9E4jpcCl+BblJtcvfPw
/UufUWFW0DMZVOubJNprLhxhhr1a/29bwugmCSNbZ2xKwbocvCSlv1a60LdaMUUq
lNr4zvvrDvWWAKCGX8pVoQqXLKL6HvY5VRDWfxJAt+qxOSRmedPsS3buky0bUcVg
0MU8VCq3tF++f0MS9UTRuZcbRmIyXHop772Zbn7DykCf4c7LYYTdu2p+fEimZUJ8
itCaqBuiQGT+NcDd+sB5hq3UBAPhkwQoBbDmJm4Ja3nmGGtuEX86c1ODN/tNvnx0
jSG9o8XfvwNh3K7fpI9d+YzmVFeRooTqT7kdCaNjB6yGGNtDJSEmIHbc/xPr4Svk
HOUMZhmVZLCCwOBjYbDvO/EYbGIPm6MrK/Ke/ZZZOB5f5sk81zYYwLajxhwXZaEH
hgN7C6dKIeWRXG3k3cJbm72B6W2v/+fMTG0olL3FyNw4FInSLf5ar85PN/5HV4e+
IGJeJCFex5TUv24A14jPKhsIVp2jvvynqRzVzhSrT6rhJBw7a+ZU5XThrFLQojvk
6MdDhwll4CviLfMrKjX1t+yUxZ1MgcUn7QCR9orLWxxnx+X7qJyMP+NMFssmbwgg
mkgyi8xUlymliayTwjNN8SKyQb1Wzg/aAq+YCPebQRLPjbdEBJS/1l7VfGT1PZwT
ogmB4Nl82N0AQhmfkicqsmZKCy6Jn6/wNp7NHaexYzxBcCVswGYzCPvbfKGOzBli
/RBQZsyPn5GAS1aYZ9DAro/ccTNEDI6Qpm5oJEOqwG8j/+YlgtTSaXf6wKNVmQcI
ghZCqIimxf2IbBAw7Kdf/F7pwyqSwkXHtQP+S/kL3t3VTA7Ku59AkNyi1zELghdB
ijbPwj66WGt1Wfo4Bvcf9DsSF1qFRsyJSlIOrgGb0ij6KbBCCM4zEsZMe3LL5Wgf
6MDR+AZk3ZQHHFIVE0xSFORjhyONROeW6ItoI8wnLkn2N18wHEphfuYjmZwbflQn
Ib/vWsOEywqkMCruYjsXD1DHPa9UuwsIf3K4PTSEs+LFJ68fAvyquqbP7lahP9uU
zsDB4lA15VoB+QivcCxxPg19OEhCYLBCJO5MB3vH9dQNfj7g1ORXo9OUQ3UfkmqU
zwTmnU4rqYLvQh8cgrpj5jJDYwawVT6CEEN8Rf6PGOaDNEB8+rtD4ZOid3U1WVq8
m8LjMOPVcouLGcjNOdCW8p9WDEQonGrZiDHKwCrSvDaVWPpCAm8FtxIVVdbyC5XX
b5PLQsnP9wdY2Je+YL8l/oTBgc+zvIrbLQtKYCqo9H0gY4IS1J3Xb6yEs+GpHR1d
twozOMaSdlRUbNIqnz8TP3lhKMjrOMUeGQpybXKxQAjLNEnVwU4NjUAkOAQ/9aHJ
exN8wQiGjngfLcfhR7ZaoWlEFxBEZB1R/zlZL59viMRD3kYSjMg0ww5k8HUO4Cr2
fHHRjko52962Ce9mlzmtHEwESEmZjgOnoIGXWFcaWGgjXN0Okas9erS7i4KExJEE
cJZ1sz/9iq4qYG4L1Q4YveSQILuYFc8xJhsWZllCfw660wFUooMI2XTDcPNDQ6JL
ogGhuruea/orwiozJr2kSqjmuiIcPUeGYBlqxmH6hJMxMOhioZlQ6LyWIjVR5b+/
8I26NpcH6EVLaSx3JchrLH3o5FLmLIlcRf+pa05V5ovKQncJCqAZmMlyRLFQ7PqU
h4o1coP2RU+DAOFFtDA564wrejfiJgGLMdSydRLHFGxMsZVFPYUW3RSK35DDvF7L
qXpvuWUV1+iHQxKs1G5lyVjZLxWyP9AcjuAsipdbLaOr3gnyaZtrPQpypbJeHUCo
J7Eb5cgs/OT3o3VBzcL1kLYqyArZicYi1HvVFaTf6bnIwDUu+BmRjxkivKq1d4qR
tc9I/E8Xk+N6v8iClfs8Jx3DT9JtNbho/pFcwImCYmgWE2uSYA+c+xUcYL+uehx0
Ci0XjREN5UM6FFXyOy3yOw==
`protect END_PROTECTED
