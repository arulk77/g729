`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
PLIDLVbqRAQpzCSeQQ/GECY3xMLVppxyMwv+yV5ElD99BlojfcbfjmRJio7RLzFO
ehu+wIei7O7FWaOcJ1aO0UIVoGXAm+7xvNW6/wI0AdafjrhzR+rS47xGXhfCZ8AO
/LSvrpEFalA0wZg7Okqfur1JuPrrOF3CMBgJi3oxqC5i/gm6P8gBFojFJlq3WfdX
gJet8bMB3NDorTwxrbS8m0E3tRyj3/4HKZD56Ca86TSkmks6YN24AF7wfbM9WhO6
gM7iH17YtjoxwcWGBkNPHygucCUIIAbZwf0WrM8LG0TLVOwjMuQfUYt7SxC1ydlx
LAAt4XSKbiq/LkdosiSYmjUy+gyb7jm6YVy5oRIwnRUnlKQR66xTeR+bHALBDRnl
0LHTnK2GV/ylV3bqcaTUMRG4BUl09tF6Qa0nUFzInGw=
`protect END_PROTECTED
