`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAR8co4u6SswzjDOf7EjU460LV2z8upLqUXiw4JotzH+
Gh8soJsIkYb+yZY4bj96lI+3GK+XvZN/BlvRdzdIcWB3/ZHbszTNyUdmKntqKTck
c9A5uvaUudn/zD7+g0TkgYf2dSoHNuU298CWvPRP0Ve0sdk11hNvWWnPuZ+kIJ7P
`protect END_PROTECTED
