`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C+B8yvzIsB7Di7GDqeF9MFHvC+f3ZS/GSKZDhhRAE8B5
MbkcQ1mbs/riJT0g26npq4G82ti8h4w3wL9h3fCjVMGAXTXofdjceQF4GJNDzB8B
/px3/wgfrNrJohzsQ0WdPYmpubbzq6cQ2fdrj6abKzQ4ZCyYrTkcJaLKUAkD5kBM
QcWV/cWdxnyx+ISGmDbNndAqgZuSzcBHTzHqpeQ6hjO5xxt1B71IBzuOLitUKinN
T2LJ2nQqj6HJTTV6D7QXfp6OHGgOkEmxoEIaQaPHhW5yoTVNch/WQMGt9gyNCWmo
dZVziBXMpi8huVm1bJwYL2xMVq0xds0dEcm75Xx7YfHAqIP2hib42YagegHWuMox
D7MCTuiNW9JIu/eQlPY7et6EVw4/iMyHxo/dgdouxy4MEHQoNBFKCxe7eRa99FQi
6Ak0tw07dDClKl/pmQ9XNipKQgamFCEKsAw6DYzQBeQhXbGxbHgum+xuZJGLTAti
tnt/kBUlnVojfI/ANFiJC8UneMa0UhJT+Xsk5TmJ4R+Vkv/2NUa6T6GgPr5hB/s9
RKD2j2BIbJMYgcOyembPBUG16WPTsRqP+8MQCygsv9M=
`protect END_PROTECTED
