`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCLMCyCa4RVTyWggTjAqRWzyfGYf7ElbnvPMjSDAA3Oi
QN3/yE/qQer6cGr4Tr/+jOlEi/4BEXx8haPTzMfHrw2RDsxTX7SpLBtN873YoI5n
4o1seMA2UrB09gg/Qyiz0Fd86/aQ/1o2cAXSyUG2d2EvicfOXMwcI1vuTQuUnPoY
NogOnVzzRfYU3C9i+GLd175IMpMZIQReIls1CLfZu0rm73JPF92OT/VbcuUAntua
nc78K0iUdjsMpxMJgfe2DTbPTwDBu4SwR+emdxP/+5FJKKvc3MgzupE4N40t2Jiv
wubgg1E2hRWvearJXpaiiw==
`protect END_PROTECTED
