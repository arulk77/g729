`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
MCyD3PkC3paBev+QQgoi2MqblELY+MiFiDb5VSr09mEaEp35xrEUQtDT4mO1bsGS
m0fHi9Ihmk3HuBOPV0OyZCcj5PSQeHPq4w0ngSCCn3Tz7NNGdbJkrY2AAStDWyoz
2cp9IpZYK+6d1RM+mwkGuBXym4j47WZJV4NFlzVJ/sU7QQuKTCxbFrPdttG+0VCN
XL3zFbd/HN1fy9KwlQQha1MxfMFdOPy2g4BVUU7Zwtb1oGTv+8M5RuYo/Nsb78hR
dzzmi6H3SXCzmqHOASngo3+rdpdbiB6eZUdr/4uFRblf/ljbGVWCakOHAIi/SUC1
bliOPF1dvyI32B+EXFdX9yDPvTieTiWaboPDhtVCl/MMjhh1Nxgbd7ljv6UzQz7j
+ZSIN2pRVdL9khaDBRricuJiTAX1fCob1H7r3B0Bnamaeq15DB9SmSzGX/m6AvuZ
6nCBk8JHMygvkIvrhPWvOf7rEXd/ShiLIj3GTG2mClksdGsDEZy3i7+oqqdhg4Oa
cRwjAbnEUgoOig70tkO0mBQpPgecXvLuT2+hhXQhJE0OCh2ZMkMwWTXgs37lOV1y
tUB8UH8Uyw6JzioT7wWy4kGqEzvOmgqQ9uTRoYS1+LRlsONR6LrTqFP/1xypc4LR
JQ/zmBcqXnKeJWGdnnCaWpnWreN4xkRQvTMeD4qg8XXllMRgV0TZmpB0p2Oz+iJ3
9aLYF7r4AfIu/OHZyCS3nLwDCJ8zrwKJafNIXg4r+8bxNLjyLAE1BLzVjhkJP9Te
UOHeyRsdgoUji55y5uao4YDTm7xUlY4KuTbygMWoQN1/NcsPNyY3ScPCDdtUVsMU
0wJjAGlFiDNAmecT1HbOgGknmFdfuVXCgKD5JUCJwOA5GtTZICPiAi7qZYTOAt9m
nHlXLMoge7g/KqlmVAwKPpefdnMFaMgc675qHFZXCYkHyXqubfs3cN7n0jW6koxP
GYseSnAgvDhfowWFf6DbpMj1yW1vpQtxSqS2nvEpXjx4E4yucGRW4+2gZBzT5TMk
8iznOXqJML4tFV8seTz0ZQrDnTBKEMIzMWHczsCCkPTIzkO8s7HGki8BM0tDN7cS
4iBQCYvMIFm1EU7qrqgkmDVVZyEfvqW+heVsytKO/cbyUN57kZF1tyCbvLdex4YM
A8Ri565vWx9CPIVOuRTveeSAh77+I8CLqAlHdChPLHytl3vu7NC/rllp2laN3iNx
EVWgPTOKdkdxHcw9HJvvCNar1BJHQsvC2xy82pr8A9k0GZ1jk+zO4+QpnfGCeqWw
4fo8r8OY9Sfx6Qk4gMPVa+/C2soTN9h6MFsdHTDVxi379blzxLo1VYwoMi8YM/7h
w8WmHdMnfGyWpMVNMUXrlitLWsuaKGekI1Ay5f+e8qWOsqK6HAY6fgN/9Rj2iPY2
OWSMdMUSR8ksNj1XpBgPsHCTj6glTNpUv091sIhxqQvsuBtQl+UcXsD9vXTco/MZ
EMSYsexO3TwJ5PdtmG3YszMDDZiNlwzo2nngLs2yLzbqxVdenRO/PoAGwMrmo+pI
slP3UtRAQMPwGNQsUddwMEXOQfuf4Qq0iRa1uxspSfdcibOKeCz3qDlQZ1rbfbMP
DLzoVjnYBnFyUgRNKMqHq7ADuJRrznV4+/H11qOHCQ6atGPEHJfyTMsxWU/6bhF+
f9CVUZjgYed3A6fhaRzPUGaL1uDslG5kL6IjIPV4rkdjCji/494M3iQ5DOdBba8B
kGqCK26/VQ/+ExRJvyCx0/V5Qx6rrNzy2YpdwWHRiEbWADRUNmpT4+WzgZpi2E1/
sTom/8r4C5EsUe2rbvQFEEEUp96FTyhwhdV7X+Q6sNUX3eXH7JvXP0k1mytjeH9S
zolVG0zQPMW5mvK0Z0STWcxSoHULxEVsrWBG31XqkJu6W3osKqX8QEYpEbZ4rcdi
8A7dub5HO4iFVEIDRJ3bE+Le8bOrgFTTfEzJ3MFpdpJ0NxL+0ip5vZva8dreRWig
SGBVoU4URxdoCFtLsot/vuOWOvtP1ZFGEix5L+Z40faWLRJW7rKSFuoy8kGwfpI3
BkPlpevZkhtfL8wVd7dIsGkutz5SJSuRQjYTWhIirOPRtKcHAEYW0mTwkAVbHIkX
PvhGJ5tSRY/9vU+d/+wyfKyjhN/m29S+S73j4r/s/fiqlEMkwJrx5ryE7694s441
U5vCBenao5KMpjy/rTnUNaHLJ+b/GCr10sk9jMVzNKTI0eDZibEuqLoiAqCMChRS
NXudftQ037vs9tUjJNKvOy0y0cRrviI+en9et+W7kh/36/J98Mc2bNJFhVm6zXvB
1zyK183S/gwdjwhaEFW7jGS6FAqUfH/ysc0wA/vG0PXwVtenMu4QaCHVcfAR9BKf
oN+PZl2tA+/AYhpcs4sYGLPsaGaRmwG9Rjc1b0o/G+yFVGGesLTAnApTbzInUFWF
TsSziZ+1TDMGbSG3zX14pHpOdxIdildoH5RdCn/fGIkYFYOfc70VOiqtkExMRSsm
LiazkgA/6SxMvPX+NBedtmOTE9MzduyRSBS1xOkVb9vaNzn4veJwhcBZLeaOR4eV
J/RVizsZCBrdPR6eYYGcaTfbnsdHsQ6c6/eKnDYLkLNNXIWeQlTFSaqKqgWqRzhR
sYK8u6scFVUDe8q9zDqvsMNXWQxKkIcg+z1QvOFKK9dZ2QYYPfeheMWsZZamdbd8
BgDRmsr94wixoS7uVAlQajKLoJ5bkuyARx1pR/ky3u7C5vnPyzOzEOJcdnoc5oi1
hQa63rOy8JEQI6mD3kjO4yTVRceOQ7AiVPq8lcCbXHZEnFn3d5yuoYcsePXiLvra
1DViEsbnMza2Fv+w54rin0I+Z8UvUsRVLdEd88EPFJxqfu7aEw1A4dtjThbgu4lm
00eM5KTiXDRUro+mRfJylO/NKOlwN1+/tz27aOekF+NRLgqH3P6MdEMFFp2VDBkW
CAVSkAFBkVa9kqbPAai7xrOXXnmm3Eqo63CYCURUq2TFFKBvK6COrDaSaUr40YRo
emr67GX1ZO+bGY3ARDGbFo3Ze50KBnvZu7pErCe3iIEbVpXfNbjJP7JSX3cvNymQ
A/BryHh4IzCc47ZPFLeSGYBbUZ0omPVg4btFOvsSEE4ePZvo+5vMNhP7hFD3yYeO
dRtUstg+n5T8OiART3hhPMhVQhntF0nm+ZfiXYWlEE1sdxeWCg6+AN1uibs/X4MR
QNEZFrznbH9As/wbCeBUcisjHnZa9hUvUJncLal8c7khkbbSK6ylCdJtN9hkjBJv
dVr0e95wDHmaoWgVzDQJR3dH9djDc2UIubJw7tNr2nt3CcsUgi72jKh5vhbOk2TS
x9uR67o/zPPDsgB59pcWCKky+xrSkci249cIGljfT74GI24Qq/oM/MoYEX2ybzJ/
S1vtVLKoxs4GqEA9OjKtZUH/1x/mOACxFBGUlEt5RJecAfHzzyvjX7rYaQirtTCb
lLr6/bdcRDUfdwV4IlzX9G8iAeGTeg3vuhDzYOYboxKx7+2C2DW8mkr3yTFgMTJS
+0XL+8yKFDVrLzdHCx8MqUKaCvzMRGWIJ+73h6rJP3WzjZDm7+feMQhnLP9EssjO
W/vCAJPCCM55p1H78nJKpJT9xEedytK+8K+/Mmeg5LJ3pYFoSxdGKwSuBZXKIwQY
IibxiThdn6J+IRD1xTFfzrIUBYYSPkd+IyIrzT459pDyi8NNNKcs1I75tjcTXsof
nqc4Hncdzttzs8pcPKLbXBDq+NsgAH+vQ+zlzrxcZxG6FQDROFVdNA1zV3MtVBiF
ioG7lnhnHcDrpv5Ffaz+cH+XL9pbAJs20g9Nfzb25iqFGo2faYwDec73H2vVSv47
BeJ2fhHa7TKhQgzi/QQXMySQflxeJy9FnWaz/CRy0ZCpbeik4ItPtBxJ1bQBCR48
2BMKncHmGbc2SJad4IuYNC7Nb0npDg7T9VaWlG8TyR1apCWabl2n+jfUfKSuotrw
yKoWuf/d36wKGga4u/pSpy8KpPPL6L169NyV78fjQc/yKzT3pqEYtmXQ3ewIJO+D
v+3fTlCg/QKNgOOv8uDA30xi+24H7RvsYS3oZZdyyO2ehAP2kcz/0wIQIlhQyF5R
hlkV/1eUq7plGzlp0R7eduRUV1IgJ/WjT1IXQRC1Jeu2kGUthTmSdp3DJ0EdqogR
sgzuMlFGdwTbdROjEfh2Rp07sQhv8rl9mdAsdOV+2Dg1DFIrvonm8KJKK97vzINc
cyajgTGMW4lTWyOBwOep34icygcF1mIo2lAm9SiX2rPS1jmomUm57sB4ty2dC7ni
3gptqUBa0gjdAXVSFCe9Elv+E5exo0zleLrUqumEaVrTyOkoUrrl+8FnJc6v6iku
iBOKcNcxpvPOCtjLbDMW6m8dIEGub+onWr4znVDwTxhs8EtrmhaEs4bR80nZZj0w
5GR6TJgTCkgltYbA4zyDijOGr+hpD963JpL7fs2nfixsxc6NqygORWTzlSS63aUn
akKvnzM0gOcRgOR5m+mrIDsXyTdEJyCCoOAT0kQATJpvy2E9ttQrK4G3hkmjebw8
AQvEa1KiQP9I1VjN7vNiOSkvlJJ+XffbYijSaxDjPa0C872+g7UA0jR40AK3veai
uPxu2HdyFpy8mrKY7Yp5pdzAniDtIifKCQbYVw1SCDXgpNSO1u0CRVHt1zdveMBl
6poWSgaZcAr0AXC0HaRpXqmy/Df3ZL6OCVoy9dA4ZQLGenidoHXEjJbz0oCLF2YS
gHtEyDY+3CyBwRRjeXDzF07TjjMx/rhtOAYZeWAz4Zv9cbecLpnYrQQiLXh81Bzk
TJActN6XyDoX66BcvY7tHQSPudIxDbDqgRT7nIFtoYMrak4RPC6rI7m6TkdkG+rM
jeEWBKPJb9ayXwkNd2+MXxbsgtDPfrDeg2MOIrM/pn5cI6Qxg6bD8zDSJW67D768
apx5LWF1LjNp3b4H4QDJFusKie5d/BHjAA1/eqcHvg8T6mzJg65oriF3SrUazdwN
X6BzzYVHzLcm/YVt7u2409N/JRaRuxr7Rj3AEQr8mmPwjJr6eZiw66MmNs0SZW3A
JsijXMxX83ehAtxPU3nYioLHEyRJ2fuCG2ML0IZu2M8mA3hBfm1smEU/Q3iO/IhM
kFlEItho3Oac4rKg9t5W4VQQo5RQjvKaf+VIUA2WohZIFoosqKv+kfivvzBI04i6
hdGB5AyvE/pp26fYYGNr3UD4wMwcBwIzRQOcvGg54sTXLgRgA+zzGswINuINvEBA
pdi0WXWd0B1m+fPWGWRUjfWurPa2AGcneg2GRXeM6fP041j3MSc6t0bkQuG57dSP
2vODdJTU5E1Aj7PiN97dekX9uIyjHs+9kxpFKiCl/pUapPlAeFPRqq0kdNAPaJpr
3OmT2ecbDixTsDdQOBOkTVtJeOPcVtO/lRM76p5Hu0hSVn3Q+aE02fEBPleueoON
3d3wxHznhT44GW8mTxti31jb9ZcA5xtJKx3pEL4DRnEe5kKLYAWqWGito58R7OUb
oorR4JHfETTaAnL571mvB9b8Snw6t5dAfIcdcxXJREHPwoM+bOE/BBlJ/pcP5a66
zozBfaVFcDZENyj9xrzk1qmUk9ck/cMZ25sAdgU8jeOMa1mnflKnLQ8pzR28vLku
ttoDSwppwncFycyNoOSzBWgEaeF65bNFR74mM2WXLFGckj5Ed/n/zRdhO+oqSJv3
i2FiME7iYf6KhszsIMlpUm1MFFOkpNMhpaoOFZmpypexU1HzFBGegtufv2xYkRy6
iH7ZeMFpRLWix4X9eUm1YtjvWFuepzcxUR5weASqEPMISDTE8oNaFHPV1Wioj6jT
SnEtzWdqeQvyQ8DsxmSXgBNEypLIrsBVLqbO8NTsrUXadwP+JBEzC+C24ifogC+U
10SGfKSLYgqgpQCwg/y2vYZlgka0Tbf2daF2VQhNzqk6iq2Tf4Huu+dqWND7F96m
r0zKi3I1uqV8LZrusYYVAKIHL2LkxXNRqcTwge9S+DMkB364MUorvGUZevOEP7xJ
qRaCd2nrlcAPbspOKVGKg0g3Z5LD7vT4zjxUNp+OvBajVqUAjcyuqgOghRgx8SRN
r44cCUSMoZE5Ol1Q/Mqs/dDf8mD6HLPQwS8oOxZMbtr/uZ2sqWhuUdavdbBNPI/K
VPB8w+gZ/vsIKbqTWw0sVJm/PFgRtscZe/LMKC/vuHvgadF1dFf3+pisRZn1t5ld
/cIg8ZZqeWYNqoDD9L/UizgundsyHI0MTSJsMxi71+MYlag98aeXkAdTy/NBLZmb
xpGJWRKDDPTQ7LXwDT0gdIPPp/fl8cTE8yBRAz+34ii0T+h8cxMZ3K52X8TUgjcm
RBwf2/nJy0dpyZ/VmMcQPzwMtMLkgZ5++vroq5mnTGNREjJcVcaQY0QUf0rGLWgw
Aq29rM0pqIKy7PTPQx8kC2T3ZoZ94IBk03JwO2c8/K+Fcg7vEXVJtyrOzmwLUWDs
nV8na8H91psgCEW4T85JsfhGWIDCN7K27nGD86gYTfRDkJcpvIRG7aSlfv5cO3vC
YsZRU31J330kQcNcDT+HcONUh9WdDPaxaxqWt724B9jkwobCUULc2faudu6KuPIO
p/qx8zHZZLCarKNg58GkUfI1yD1Lb+CmzU/dUA2I/blsvYWFlKQyIZcKnuiCAWtU
rFtxWjPmVhGOR/XEDFMCVeoROukjXXK4TvBkSTmRPv+bFRUsS6928O9mW8KQ3W/W
jGWY964G+jc3AdS2riJQwLPkb6B7R/CeRU5LpsRmSiUeRE8N4CzV+soPEU8Xt8SC
ibYtvFgKOrDTzWfBHjGpQIXLGLmwC6cpZCMFdc6yhAi+/BkbLjOgNRCDGA6fDeNy
hBrcmMq43cgky7szBtEtuM6hE0IkQ6TNprYQIUgIN56pSqq0kv6hwK2u34c3tiIX
Gg7P+KB/t/4QoakE5KqIIdUD7IDZPQJV1t19HPYANV+CE80pUoXRj3ZBDuBmACJd
M/E20aPyAuU8FCby4TIJdReVAgFtGa4ILXUSajSpN9FkKa02rMvs/qb3MpQM9nOE
BTVQcCKbRzv00Ls8REBDzIn/86OyRuZS22jbwxXwGkdeBnxPilTLVCge17W/kqrB
b0TFILs5AVDCZqdzpOjg8wXeC2++ywXrZ9Ed2QUAA1Ndv/YxPlAunwX4ryuTW7ek
KaHasVyrSYFoKES1/9TJbmRLvl1Mi8G5rTY13tBTaGVGKs4Eu1yWyGslNkoMi5RM
qYnRXT+Otibwroek4fplkIMmkiIQhLtNeTzei+0F4tzN75C4n0ccJidrqRWeyQtA
44dvTQ6fKtdK7yksngaEvVANpUmOb4C/1ewQDgnhV7C6n7BTMXUI3u7f/NyQvfLj
86XnMiFWdy3xNxGXGyaJRhSFssSLlIijB209p+DZVtyldQyXdVOGKAk1AcadO/g0
UAhqJr0+VsoOERjacGFk2ZGxyUi5X81z9FBa5b8mJ0Wc6dR6/KZspnkV9T1GBC65
6BO0tIw54CklVvUPFXjck7WpEK22ZJ7Bjr1Z1XGVGnl3juG9js1gCKt7W6SNNtN3
hr7CjjHjMFOZM2IEv7KredXQlzSeFW8G94M3HqcYfJBxyKd1do1cD/UPzHYgH8Ii
bEmapKxdn6aVMgpROHUnn+XJjMWPxBtLjkLVwSXeIjIgldXoj0klUkSkBiHv2sLN
cLfz2x8DjHXUanfI/ykk2tyTyzBgXoSsB0BVgR+i1tE94eC9EeJGKbhazInfEOFU
M1+O3IoVrzhNKiiq3iCuvvxQGpN3/fXaf6UdP6ERO5evjnESICiKOqAR8Ak0ffFu
6LGguyXmhGuttDuXiE/kvWIBaB6yuheAdkwzY1nHmfSOHylPzec1wVef1XfYl8SU
sR+CWp03Geiue4fhMRpod81mRzw4Jz6bA3CQfmEgtXT9QddvkMMHxMoklTXMdq4q
9KDny3WgobastHpwERHp2q5LoL6HUwaqPSi/7/JNwNZ99q0WNo/iyMsAFokkpgbk
TZJYzASjK5UuewvYl/oHWMxsfcfRWYaAbqr82E4xLW7jp7u2fOpvQQR+exCqcmLA
03iFLFfZFfTnrCiBQSk7U+1xPRX5dR4pkMkPHzF+HkR82nrwHUF4zSyZBAV5dqIh
phgtSVXpZAjgZWYZI6Ckf5yXiqKHP9tcDF29j6C5L/xeas/7qryO5MO+EJoiJLV+
jNtVmKTlZdcWYXZfs3xFGldQEqVjuCmbyD2Gfb0td9b+mMOmUK4yyS+NZIiatbAH
zxgYu3E3wwquxJSVMFncH5EHih8J/vytGOHc122AwYWevl7Sn1AKs66XaUhEbL2t
LkICKI5D6r2R9A8gi4+FrU1yXTEBuY0hmvmlEX2JXY1qUrAFs+uSKkgRSveZGF1c
O8lsoAyCx61Cm08AWbfSKer0Dr6tMdmqxC9dWJeymi0FLOU9oA13uIot8prmUXz9
uORRUGapRUFa2uVb+8k1nUZh9FZhwDffMswGtXUNgVZMpEECdlEOwUFUeyetlLDO
IZ0FrQDoL9XJvQ+sXJwoJhl/1c0Wcgwjn9l0FMjFQxOoZDzh9H5qaBhCsGitmoEw
vnDDGxXrlxl4TTi/zsKYVOoFlF7h7/nOdmEgFFo512auHPtGYAHVQGD2PXDCB3PE
q3WGs5goiRN0Y5iU88XeGqIbbEjPa4KoMJJ/nFIdaOb0c7ED2SNoMjHm03pZW6Xj
DYhslqJDHeJ2MdKgGZR8jt5QoKlDQCdx/Y/yWUAXnFmRf4lnyhcmEvqBuXqqEM6P
g8Oxrwor76LhwSVWuzI75sFZriWuJzG+a/7qNfHs4wCoIdpfOUVFMQh83Q+gPDWD
6fediR04NcW+Ii8tGtVDgr8hDjswSLukEujwpXHXk5w2CG410nzap86/jgy4DHhL
Qq7EVDNaQtzBgtc+S9N7/6oY5fOFLZeYzVKGMi8ToI2FUxRD1SQknvY8rynTOCg+
zCGpI3vdInIoaG4VnJAqnYBGaaKNFim/GNSoBtRc4yGdouzaxhsfzyTVxz7ayYBr
sFD96757q71Qo5UMJlwZu2gUwIEy/MEaE2ByWx+d5Irp57auwpLFsHILSHbIWNzI
Ma/44XX4d9Z7+rxNumet5Xp4UvWDbHBo8W5SaaWNj03KCizafm8Ku9JyBEKRK3dh
ecqSUIwRXu3L8SGsV4hxT0tm8FZwZ/1OZPIfnLcCCK/MsgTvxND2GdKB6x+2tczo
EtH051KUNNC9YEBU8gHpSSMVFkB2QGipCsov2ZwIVpESfnLKS3qA4buh4FKg/PuY
lKKWNhyPbDESesaQHZLDQZ0Z1mlRAz1hh4e5/HMqQqUQExlP9C1TzUVh0aO+cYr+
6YqJYg5iF148vvHDo6NpljY9OaYU0fI0KO9shoHln9COOvRTVE8bL9sAsZcTWiel
dgLhNYcA3Q1LscHGURH9xtYQx+LuRDR6zwWXxNxHiWOzEfuYbQyDZMzTorwaQ5MI
lKlZibOGFDJJjOgOQxUBQcVHjYCfyWvgWNW8wcMRWvwENYj0XeuFcVN8SIAjCXHz
koUra5Bxb6w9xYXkO1SI+II9dRgv+cJZaEoyBwMqVCR+Ec+zPWRCKchvk7iyYeBt
tmmUPQADdytVdB/PQ2lKIyExJOm6iNQF24wHzcYTbKevMwEqSrOMgGCq09VCJmpX
Q8/4knhy++lzuLomuAaka4AJ5bGunilITJBFvuH7bi/bjiFMaHhXTgXmErrqZoo3
aOuYAnYK9SP8gYbtC40IWp4DNHANRAovo/oKbrhjt3HaHiS98P7GzSkpYEj+Oxpq
D7M3ccbWJ6Jvn7mESWEJM8Cpa1BYMB0p1F4DGpXV0AfBME8dXy/u+qQXQhYlpCT0
OR2x44MyqHYBvJuVmE80WbyAVUL0XxqaewQ7I6Rw92ABmUcKlyao4ARBLh5td/l+
it0VpB1+2IToJwcASCQXm1Rn7nkYBd6aNrePCh50elua/oXsxAyalZBGldFVusQc
RY6dUGDxGU7iygPahRMEie6jxDRdjwBeuFgMNN+j7lZdul5edzeycldn24ySW4tI
+knCgqo9Vh1HGpjCEi+SaeYlFNMZxS9QU99YSAsJ8TmqpCP0u2YOptmMy1GLkOc5
ga3hrvvhh3ThSY3XxuvCzEI4ndxIgAW+cvzm/Xv1jAem8co7MPzR48cPeXhBXJCc
Mpq7nBYFDHvD+rgKn7vC4pywnqetoq5MVUNsCVwJY4F1so00yjQfI2jyTrb/0dDP
OCP/zoDHe1wYZDOfi094CIEOdVhQzk7luwOxJJqdwEIDapzcsHo4tHlomT/Ik6Yj
urOT6BxY2i46UFLD/FA51EREqL+uLtSRvDYqCcKWLFIwJQC5G8Kn34cHOsiflKzK
9pUYW/TrXAjf9nKESajq42MWAJDmAfEoS2oJn7aONN1Mtxx0BUTsrPSeUIWl0JS2
0v/035sJy9RoqJxOTa00kRvAyAvQY5B4d0+POvs6PtMCb3pPwgOeEpz4mLb0+rph
9Lh3Pp1FyjUHQcd09iWJNnLPLmZ7S6XjcIKyNl5FTtgoZkcpXTFAXvwkJYRza/80
hA8QF9k4vIm/8MGMKfLR2GK+MO+Y8LXWtQljChLARsbvDI9s4dGdOLKoGmI68fhq
Z03arPxDxrIx0YkZ2qxQlgjhg1PFK4FZhgbU930JE32quzolD3gF02qIh1vmbkJL
TUI6v3n2MVCvQIk2LP8C37OJ5yTuDVJCxtg0kVFmek1/xJZzRRD1lI9uYmyhtxcy
5lkoiJVYx/QN381Y5CFJ3NwUh/FrkTOeRoec+UE0TSGfwbHlGWQXxNh32SajIFjO
LFuHiikAta9/5jyku0q75BWkaB/0Gi38IO4URHJt4/B3JLyFV3c7f7AqGRHUX+8o
UiM684lmFncZqBKxzp+/0UZb9h+e0C3gyNxaLoexwfX5qU4IrCjJSEDyk/i9dMdu
0JkRg3OIviHiJIxiNv0lyTCgYA/HYtRZEM/8UYqscHxUJB16hgs9dIMRfOQrc5mn
wvuILlTUV1PVl4p2eAxP9osT7C1aRoQAdbbeqYuC0f+GNtznlIOUf4ABE4jmOH43
3pome+jw5M+Upu8FEqokRTxwwGubWDN1d7Sa4G9MQaowDibSb8eZ8Jdoh/y9itrL
rlbOF17y3dK/nqkELs6isLPJOAGmYQOwbLXA/1nmyPi/orA+iz2r0cWpMuoWq4nw
ifZrePglzDF9g2b93qxEB9CvhnI8fjFUS35VrAWD8wuJiJR5cPwhdANumQeFdTa9
olqXz8jFQOcn85CoruJJN1FdnkUvk9Bm6YTF1A2wiQIwvdvf9EgGy3rB3S0iixRy
z/RG391O4ipxtHgjjVHFiM9eE+tPmGmWro9Rvf3HwuTzTAvGTUaYgoiQ4r8xDQtl
RYfAYU9+qRwcgFTJCcRGhHq5n9L0g53YlKjBG65Oj7wER/xEdx1KsOVVF6sVcX8W
8z9w1qv5F24puPsVFadzh3EItfvBHcNxWWCvVMlfpnCAl1Jnu1Lb8YsRPDahAgMI
+mJ6Y9hQtN2Otltal0zssqGvQzxlQHOXjTDIryCNAxTgvKRvbJ7kpTGpzp1keKkS
+vLRZW5ltAy6u+bkUBMvA/AfLv+evB3hmbaL8+m5vkUpiyMhTH/fYCSKyCrZ/Mvw
8LsLLKIO9+yBWQIYphL3FN3qPUply3MWfOd+hTJTpcSRngyPtlFLjEHQ5G6R1RVk
8sgp+QqZDF0+G9K8eMrkNveA56SLKQTaQlCQFI9pdu6qCsEMfO2qBr826Upq3grm
yKxctfTtd5XKa1XsHxSQ67N8cik46NC56cN8vHXp8oIN4Xz7PzR31BrwvfvNHkHB
E1+MnVAMaiqYwwDcUt2qJTE/lc+E0IXjMJha5fZBq3vp8IabRmSIc5cUraNl/Vzb
+aJbh2GG7t7E5RhlA34MZPLHL+mul6cDaYzG8lF19qwyJLYEElhZ5Z8RX1aGPlEd
+338MFCMWkSQuKGlIR7TqXec2N/bL3oxeQhrx42t3zmYE831Hc6730rb1WODGHL8
DT4WvLD1mCE07JLfftDZEFDwyG0UWL5g6W9vWYTsoIM4YXWY2fWQL5mmCryuYG78
jA4cfhnJVIZkjnVnYIw5ZAyJUv35lBSa8WsMuT0CoCYD4Tl7CC0RT4mzWxU3XwRC
3N1Xk5u0fgO9dt2iG4iPXVCMDV2NKxw06qZzzU01RgBuDh613SnBJD6ImzjU9jUS
ykiuQkQ7KS6ARLiZC90+ThIY1ysrhi5maemJBlW1MkH7WCQ6sun/S3O3osF1xldK
EMiBCrhrTygAntuYg0qDAljtLarRtdmgmWc6aztx2bg4Y9u/FTsyz/1TVTR5LHaf
CVl3sGnKGd+/r7kkS4Wqd/n6wyfoqt56q8Up5t38KQ6flwlr3fB0cGvzSMYqS9M3
lRN/lHVy4bHWLQjTYx9w8Rk8pMReLF+ctOthjI/rpv2tM057emTk80klhfg/ryNa
nbBLRSvTnC9pfjJ+9RDKxK4NE/36uet6M1n1SuHELETJcn6gyM6XGxwsjfwi4fao
sZOVqJGdW1I+jbEPk+4KMQblwMHUVbVThojbZv1T+UKvQXag7460NvmDTejWAAPd
f6c2tjafDOZpaxUiuVg8Ja9w/LvuMwsKscp0MZJBP829h/JJtR8HACJ4HiXP0ELg
bOtayYNqM6ekqemdHPcpMJYg6gMsdbuayuT1vRgX1YQWIE8PLoIz1XgMrVY4xg+D
T3D2AJEoaQDAprnPZrl76MuR6MBqEIMeslW4AYe26MAP5dGN9O8xiwA/nzqi4vRj
+xmyXeeP+qIS6XUmVUDPKIjw7w8+yv2EX77CobTvxeVI6GL9ucvThVneYCpTrngT
mV4z2eUVNQTketgXFIqE8SokC/LySME14gSz/55tqk0v7VZvcvnJTqSzULHtaoWB
Qk8lpiMuu/O9iqm0ELeVS3TfbKKdb8LJBz1nw6hZcGUicTFE0KnqsEk+BGtM0mhp
V8HsRiKLX4uykNnpyZfNBDYggqzFP1JLu7QRSD0j+zGJdCLZ8KkP73bfdkoTwD7k
1Hjc0bmfM29LswXHxw7LEIQxw3IpvSGEsZPv7vlroSVLpDe26xzCMYlGH9qTJsWQ
yh8POFgLc3pS+RJ1bkvVfEf2DgyZqxrrAymGj6mJoTUqHaNd8R9mKLe6/SjMnFVv
S360X+r8Eaa02rKjRoSjXPBf4FSm1PNrpWQM326XxU57K57Ymk6CdHfnkZp5yJcX
g4xSXLjLauKd6igJIp3tMoLg74qXfHKV44FxkVH1rLQ2deORxxAtsydeVVHjN2C3
olSZtqDGYb2Mg3HyWf+RwL0jbJ7Cy1JhzbbD290LzzAVSIe3HFQLtPtYZP0hoMOJ
NYqsG+w/i2uIqrFwEVeRnfinrZuLrtaSSLVhRqp8HKpn46UcybfZmj1an9tgxtKz
IQxjHLfh/oKPBScFo0UPLcjWdygzW8U0YFJvA+YRFPcKRvWZbPOcYecMknwfC1Hr
ug7/omwbdfA1YMxY7de6OdJHuS3ruQWnKuPnYMcOYKyyuq4/4MfKBzrU6arANajV
dcwh1moTR2aSz0fEX5Ex0qhGKjf6JutKK8uIysIuOT53+r7ArVf4GN5GM9KBWfTG
ueGbrf4+ebMERP3YQSp/odVsQz4un0wk6oWSjPpyh/3qUdAqDnW7j8N5jJ6E/ejj
VkCmdGdV5DVURyjHDWFB6dAkbtuvU9TNXE4aUugkaL6DCgEiD76AMe/zeGH9bk9H
yQLqrV47bVANSXmmHtiZnf4RfK2lOZiXemZA0d2wP/3TJ/1fjBSEBkrgUO+7LQnj
Qnv57UF9+k0u3kOrwEaG+2ct9h0DCiROO8HCKY2bRTneVf4cN2Sp322jCbnrzj0t
Ck/MK+kIQHlM9NF84jzpii8LochXezT3zSZucL91+fe6L7TExpyoqMWlHV3fMiSt
DlieZxTmGkl0iMuoCbMR2fApXCrgWB24XdXMxlV5kRXIS+ALDo3IDZr/MkwMSSUz
AKA8DmW7oZ5L2AHqbI/R4h7O1BxOvX2dc4krDvvMLIyIuqbCsdPwQitnJCvgr7Dd
6CnB26nD6+Sj9fSTifSmMSGpV6ci487EX/FrdsphbiuZRb2Z8aMBnKnEtGVNxcHr
cxjjdAKyo5ctyqNu2m6UbQPYVjnVpIzsZ2ujYl6mrr941OZtDZR9l3p2yvFTZ0XL
q9ZjUgGv+5pOU6h+XONfvWJmQ0LMhDRkC8RRMvdwpoNDQwmDL7BNCw7sqVuhAF6z
tWiAILh0TKDg4DuOxzWSY3zqMgzqPFDr5Z9HFrO8D4fnFEf4JK20kyqPc2AB0GBH
CiPljwHNYqGr/W7QAtBQ2W0jauUNzHbj4gmXb0n57sRK3x48TPTrL5J3/INm+uJX
/8lgJE8AwSN5E4QAj3F6RQfbytJubFIQofMLpZ4TO2ptR2a2gIzU7GW0+B8frzKb
Ubz+FDiyxH8V/vlHLMwdJ8B1vY/Kz0dRpk0McuZFKgUijm8W3x15kv9q8gquUuem
3ULribzTjQWKVkYOekfoLOjXWTDf7+HROhcFNBo+fmurvVMPal/1O+PjvVg6xQDr
AcmtRgZ4ypTTCi++YsrHkgJFEhqxgTCAPsr+dj9M/VSKXhn0wJuTzP1GJHdDvHLq
TguAV7xK7FiGWqdU1HgfcF8946ys97SYs1vAdth2pKzn+Aqo1grwOurlB+e7Uo6k
Bk66Fc+TpkQdQL2ehGN2aqo8Tgi/0cat2YxKyJ6zoWg1qICi/ntVat3VYBYfdMCi
oMvs1QTTlBy6Dq4xLm/pyZwOKg699nD0cNR6WpOybeNWH2p/RuB0FCBTOQotTuhk
GQOCo34UIA/zKoRWbxNr6P5mKt2Whvgx8S0hTYc4NC5vlglUi/3+7nCvDPNtqKgv
JYjZLGJqvYEzWvnfW1BRf76UqSyaf38RitoLTwT97YmJK9g6PM2r2GQXQhJUn/y4
XDamRAu8bCvRtmlImVdvvPfbvqiNSVSXf9QniZrIsOiouVGP1NStB8BQTmdxSoVr
/n+JVpnZ9awnptF3pigz7KVof+xkz/Z7kq1bmfWXcHRuza+BiTB+EftdamSb/cRW
w4otS3aj0YS9BtcdJAu1PVejGu+cvIUQb6dbxuNMjCs3qZgqy94DiCrfHkW29WB7
isXBuRLzXyWHp1jnjM/6CnQuwwwliN+5YR21dbwfKdtLW7648Yys0oyVCCHHFdjd
FutlV3sMK30XELGpwEqGe9fWGrDQdLcLNg2pE7IWPHzrDnIXI+TE8ATa7/yqAJC5
W2BAFItWlKzayoBLH10+R5V+T5k84ObuaBYOYWDY7HCFJDkoyY3l4aO0s+xZAGgk
MJ+TCWDDGvh9111CGHMRwd6X9cq45w9SZseYYa8iKHVdnCIGjsqIXfCasAvYzznH
Bmkqr8dWQ53uSPhYp8+EIha7dAw+uLsJEJRZVDYIQNR506UkXMi7MPt+mXOcQ4q2
DJoccEbpAFMQCmqr8mGqguOxU2QZbrzdZdOFiM2Dx20=
`protect END_PROTECTED
