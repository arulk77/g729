`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveB4hw2lscN7CUFdqmYCvefNcHHUCIL7pwcz850mZz7Sy
3jKB3bab+N8K6j4CJ1b8lsn9dDGVFW+KWNg1+rnzyiZ3bZ9GyQ3KWfFQqfNnzscw
rQ+vjBNFlTmwvQyz2llQ/sF6qgfH8UTlFA429jgbtrAcl/rYJQNAKmeR2ZXaB+um
`protect END_PROTECTED
