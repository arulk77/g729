`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBPuL4+Nq4N0uM4aL5p9Gmogm413qpP1ouplML0s9Ljl
mNYgantGrZptLyXLMZJf9T11AW1iHDo1mLbN5nBVnkCzilKFVyrdrSfA2Jy5G8CT
bw09+YHGMQoFUK2camvWWcxNccVxciwJdW38gejF7WFwS43GVX9l9neMq3NGIa6u
6HxpqawujnVE4JbzEzbHAmaHvIaAnrIdqXq7HRa4I3f7gwQrgAsYP3PJlkkLjgXy
C/TO+FzmENyoXOn7oANJJRfYkvG760CiH8L6j8IW0PK+a5pXwQF5uxOVXsJhkYFA
vzqzF9vkjOojg0Fvxj5Y7ZWoPaSeaZYipNLNOzKmB+zPvcPlQWzr3EsxKxfrHJjC
FLXNCzqjhoTKbY9J2+lBb2Ka2+3DY3cZqIy5XeyHgJgGq4CjnCoNyauf9Mz1sYFb
SPfwO+VYXQjx3PTcgPMJwHi4nz1JIIcxee1PftFUv2OJOttzECZVnqXRHuhF55fa
VrsMgZk+4sSPKF0FCZZ1SgD659FgpOjR1aIAIXqvmrWfP3T3QIP738Hwu7uhQZX/
`protect END_PROTECTED
