`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveA1oYn4/E9oUuy6clHlkZ9Hp2gNO2eqR/JQb34uAuzI3
frAu+8M9/5IDsNVzT58vHRpeAQ3nHpGsDLOWnH5Ozi5xNTxJq4Gr50qU5vf2kYUb
iOEu5Rq7xtMqupxAHZOHgBvMb5vQAGzaNN6o6WFd5ZOTtrorL6yaMzFf/Gg8fiuU
T8eX7q9NRtUaUmR98vBT1dAK0GGt+U1Lup5jFyg9HUKljcJVR0Q9BPBegyApWaoQ
2DW4JUDNPiacXCgB5+/kXa34UkWwISHHNeHu7x0EVJeSrzsWXYFmFuEUy7s8zkSx
9eT5J7GG4L2jnQIJikbaFo2mCM7N4DSzaTY7Q17Rr49i0v3bfjT6zWqphTvGXf4h
l7U+kfF1WvCjXayOacivtOaKrCiUVv+nptYM7EwzOeqle6Ob/dOlvFFDSuEenfT8
PEpCRTYXQ+j/VmpXg4QPFqEKAS7cEIgJu2JUEcAQZB2reKQJPAMF67J6mOCFjoCq
`protect END_PROTECTED
