`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+i0w20fL+I4r5ieptuqWrFb3bzXnwH6r5KJh+ksf5KY
cF7gCp6vBuru8DpKSaj1yKFM/OGebErK57/clWayLTzhDv3bwa/yJbHzfdxNTLxw
aED2QGtJAbKIdujNux5qNX5lPLAzs+YMvbqsz5NfMQoZsPyDGdJvb8asvlhJXzve
iLvVH8H6dH8hxrqndWP0J07AlgOfxIBiTZ0puoFWJ+0uMntn7KZp0IOUsKWQTQCZ
u50s+JXK5QMVxshnY3Ez0sIBYheMg7OFRmUDUdJkYMur4tr1d1GElfAjB3Dec8LJ
kEA+t+MQlRfpGKEBIg2jxICIvRV/n6SNLayWt5gn6A24cUZyCsaL9H5oGIn6Gz7E
k345aRX80Pf01Vwb3Ttdx08A1G+4afMBoQRuFQ3MCVIH1fZMamqQx4x8FjyEWrPD
eZ8L2uz0hOElfMwEnJhDeFuasUKLBppiWNFVPWmT1GQ80/YwmLejQ7SgxbHU16e7
`protect END_PROTECTED
