`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
nAu+ta5S/hJ6anz5qmcLUG/fChfZ1UTur7ZtL5FA9nCJNKCBw/24JNhF0/QtNJ5q
vCEBKHJmy9u/NUdizWFDAam7eXxn/a2jgkyxBUyrIUzVFjVAVzwXglDRK0m11xET
CNxCEtxU1JdfJFAm7UorH9u4pk1Sv6B8kf5tdfp7bFaHP9GxeumBInHGnoT5m3zb
54Tv3F+xw1UM1J3X8JiyY4fnP8d/anSNBE2iliJLMYQ99KtP3P2Bi/pdolUqQqFV
FYiZjMYMDnJHURPffwTrDhnfdatXNhRKrzn8J6nYFyStvmfLA8FJRnKyb5WQtz4U
cZrrIGves833oy1EeKMc5QVRzl8pNbhkOz7rkrl+Xls=
`protect END_PROTECTED
