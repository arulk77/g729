`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDe99uxgmhi+QrEEY1a1L5GMAay35ocBXRJo57M0uTsM
ILttNXsdCPJWdFSdNcMzgSxn3SZqRKiHY6avrH3gpPmWtUAXGnXMrkx1QqUQ+ePz
Bjo1r7NM4pZUEQRREMOaYpFijwM1/5a1S12+OH9DV51/EUN+rGTm23A50DDQYFFY
z0EfQBTGitTNEM5DL25+AaK2NuR48DpT8CKj+b5wYroXSpgHPgPmtmFWaAm/FV/R
DTLwMBIcstrPX3KQA/PF45sHpVwvnxz2mRX8+7l7BAfNzUYS3ZrDZAyRpJFMWbnW
8wnO3dQDuyx0Dq7izhL5F/OgdjNbjMyfjgzpE1/7qV7N8WO3GzZqpDTwb96pUUKa
JPVfpfboFDLXxhT/T7HTng4HaUawocXJPU9zDc6gOl21iiSetgST0XxqfLX41qBs
kh0FJuCRuVxGwoxdvcMg8AF2cqYEJ99N45dzBGZJDfWIckaMqvjFPkSndjzEfZli
xk3zWnSglyaygXkrlT0NsyXZ+qgCcljBaO0keCWBkOJ49vY4jFlovvL7Kmko92Kf
`protect END_PROTECTED
