`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
JOjKL++xi4jTs5xdaGPUPdBZkEWxbYjZlwChqCF+YHwCU7IxGIPMHZID1eNVzJhU
YrgQ1nBhyYCM8e6w+p/EdpV/PNJnH7K8HNXd0frAy686dH7YChjRUKg+dyRPULgS
AgpcoRFSQ2qprQU8A5cbdH5uawRaJRBte38WEdO/OpL2egmOVBsfDcjoMGuzig63
/qQBltyr7QFEpET83knBroiEvvBQkcbN3K9tjMwyEvxqDep/eTFjMZMpqAkWHqJH
OJGvYshxTgpZRYxh2G/2+chMsGvwubyGHk5iixKXsv5sFtuAEymcQN886/z3vB76
mS/odE84ABkvosdvNWUlOMitZJi7QnQh2HWVMhFkPXp8H6s+ykDx/6APQRsaLalX
B4p8IBaW3ggBfJSAt/T15g==
`protect END_PROTECTED
