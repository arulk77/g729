`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN5a6tF88fR79lJWw3TP5xKSfn7TwWQ6Sk/rnYeQhEhtR
PWAdm7z0Nw/D7vkfalWXtkzUoCr+eYo6JWpaU//iOnc6hUxIDzuhi7Xc2obu6R7K
pCdnrLipd1J7p/R/0umnnSKlinjoq7k6njLkk7M0mxyn1NEQt+nn2FQndLpuhpYT
CUiWOpIYMPSu2ZUMSDLUDLXaEAM6dhly4Ac1AzPl7UolZ1KhJdaKSkDgj16exrVt
R8QHm4JYfE9VwPKONMlJI89fcIhqIQXtxc85SUJKiP6KEPgJAR+lXGfQYzbeNUIj
SLqmzX79S0aluOQA92Fc9lUAyFSbzRFzckeWACFNnuYVwbLRliWse99Mii3FyuWl
duoKfnZJfl+iIOrQnEVxYUXP2hGzWxh1aaNvXcOPQk7153Umshrh4d+sskFmEWV3
i4yzg21hzOlMijpq2ucyCEm1/rZ8LOXoSafJ0JwFx5mh4Lx9wcmM5LXaWUfY2U9t
/QvbCL5llV8dbddtyaCHeo1mO+kMlAJ4aFDemEskXCkef+V10ZsfoBhFfklHxYZC
a6JSVqtgrnsPY6Zy5EwADuIvP+XU+BMt5S785fIMNn8Fxb5KZu6ls5q60ayRmjZp
DONY2Sv0d8xnLd/6w6zWbcVrycggXaDdEI6jTtxgEe0tpPVw8pLxXs9I7ZAmtxgM
7iKXP3koXIYJOi6hIRmdqWPRvTiBa7r4BcnT8nfmLZeunD4+08hVoU+dTkQCMpMF
FxabGNv9+5Ro/yy7meik6QOl1B0twAdc1GmugqqG+JQ/K9vwQtUuzEfqnmzQ3284
XXalk+wW1lEbLU0Ze92sC+nTLoiCDPHf475H8mV0glgKHBukEH/dI6G3Gtb9CAMw
+tOxqRwyEuzQgJIunLWld50yK+lG0ZGNeNFh/P9khOOQvD5jAf1sWLHg8pJpJYPc
s4WFvkWKkf+8RO3N0IMG7cduo1rs6EeKc/kgX7mmiYfhwTD7bzSC023ZOYtqZ72h
5PbyuzhG9/a8eHd96gJSwvqvZwA+LDdQrxMIhBBCf6hVG23VJ3FZgGOkgNrbNBAY
tkeg8QWnyVEgTu2iFe36WkMLLRZtbeNAew5V+Lg4bQ+XOWu9tfsH9GCKwaCQd8iQ
fquhWtTHbRez6vdAt7ZdL7yDBJ01AUHQYVcY0h2P+ua8xdfz4wde6zR689p44DON
sdmhi3zIGaqfVn5Wmzv0/h96Rnnn0KOLNshhE2KRV8OL6m0t1sV4TGKzUr01Tz18
Wn3CvRkn65fkBsJH7CSuSCIda32YhKiB0hNaRHdGD1O6zMvwew/jV2H8oXNDPlW3
KqzHhBLNqFQeaLLjTdJZBSxG2e+Y8ImTks3VUt0E8mt8XwvEJJNbajgNuYk+Fb1o
gUqN8lodwx9YfXkUo7bgHV10uM8bCGFS4kvy08gjwA8VilMveqMOPjQAeIjSPGK0
NsDaeRa2f2i12cDdoVSXTkPswT/kJucJnynoaWwaW/L1QLpM9hAmdHi/QKcLSu46
ejgw5Zw6mym+e8L3/6q66uG4NL2VGoIyzDDuz6qrOg62HoVV2BSEWL6VtQNIrUCk
iTzOVLIrEG9s3ZkcaZ08jWxJGutpsQ2ngBcFZrNwtJgyy2XFB2cwLc2mv2QWzGiM
YkFvMMCYTR7WG5NkD8kaFMB7T9TjL6GPJ4yathjCTJuRP+zxCaXoXplxvvmIFHjn
tVWuXqCQz4R863cHZZGlHDGboVW9tmMWvbaBubgMqALkExEi6L7J7PY/s/TjkDhd
7s8pGX+y84zrSIbHQO3Xxsh2m3KeSeGPCdRipGPLjgC08ol4TydQVRNPb2HKSiYd
cxJXQ9uNnFOdTChJvn0ceCsPJZ3vQYDbhDWR2rW7jE1F0h8YhkDO+31r+dVz8Iwf
BIGNhGVTjz7bSYP3NoIjq9+WnPErETjsml3bYymbRD2rwjJp5OnI3/36oY/PwznX
aSt50qSJNQpVgIcQLkQ40gbPxhErbqDM1pe7IjGL7cZ3cNhXiY64716IM2uv3q0Z
hb7a3UNGE2dysSxDs/0dS1IYyntCl9HiofPmWEsLU3wqxqxT8fuw900KeQjSDsXm
IfPIgoMii5xIVzQoscBSSeLUXv73Mk0Q/YKnR9qwvnw88YwsBk13XvfRSYDPLsuj
vK0v/e4LUenoXmhoB9PEK90RX/j6zCi68UjRO6YHhOBlgBy0b9e7VSpPfVST3VCC
vJynQ7QlHx9NvRkkdx7rurSwfxC7tCuXh8W3ka7MKpBx4QWAvxLKB+b0L/veU4jz
H9Wnzf2+o+Vmfmi2vJUsHVWC3nahdis7mY1512zbG9V959fBWKvVeBR3f8ws7aQH
ubTAcg6ChWwfs7On8vCd9EQzbhnvdz6Acb6GWZGHrO3pDXvOul4A3rNIwn2WprF6
33yhF7ZkXi/4SW1EOquhzbzYzm2Qf3iGtVFL2SkL4rdZJ47iJlhEsq2BoZp11292
OfCXEZv9Atafh8snDmsW0s2a/EiX1caJbIX2It5DSvB4KyY95IqRBo7BMYUhr3KG
1bkdlfrDee3t4QA6NWzpZy4+ChveRmNjs68y6qj4NHz9JsOUCGPOaEGOKJdHyyZo
anP28sZBB1GxU8JMMJ3XPYJVUmTcn+lxsNwuHwDBl5Mfw9SiWj3vv9jywK04GGSC
sgZP9PlhKgYA9vKUyFU56OX09zJm89idvKjFnaA4u5yR8+IksRITbuC/mxc9PRig
xbnJYB0hpcvvaErbB4wKYa5Vbnw9kVjf4zIorhRSFddoGcqiQuDuh4N0ZRLxxOvk
t1M7+mXNPQz6OiywioFMxKklBXYpT++KNj90Jno57nqBzgegLPDBPl8ermOBT9Dc
zDRJEgAFwrxkAWBQYtDL1OMh856VF6xgtpk6nE10jFFMXlVKON3U77oQtfEUCUXY
l52vrNPMBmdgBiFni2sEP/Skyy6y8ALHe44xlJdQWwMD1IsPo3/F1vP3q1wrhKgU
qgNaWw5uh5MQh5BWRaVoapBNMg0klWmKZkGOKOrdykbO5luiGFxN75i3olCpX6ZL
nd1dRxEkgCa7GD/W8dNHEWVXE8nLyNaUwtYbngdHva36DEmxS9/D7q/bzHNq7WgM
loRbL24YodbiZK6GgHbOd96LE59P/D9Q3M0EzWVzlLmit5WeD43Sz+jRPH8ivOjg
f/2UEA+guMJ34TerzQt0pSQh6h1U4y3YrWFbVNTdFL/W/50ywyeY3me/yfr4kjiA
HQsa7gbPuSkY4K1jm0+vMAm15eHCbB8yal+D3n+6xcJQzVx1Ujzab0cJHvlKJxbr
RlUS7gxqskf20Q1wOB7nm0rleFWrjG7IjDF0qU2rlanlcD0JFcaY2NcaxNPSfB0b
msBGimUoY/5wdfWYuFlLWqG+qlNh+kjevRH8+9w4y84m4PmMeyyI82EAu5WDJcyT
xWk0/iWoxxIKSXBuoK/IGAk9wMasPfjQYB2SLX+oO4yiNLgFHwuTC3iPPzLR/SAC
Sqad/6RZVAhySxBzP5MGBfzMcW75pvsYMCPh85cmx1zbOeYdiywNHolfr0bVzRNd
YNMOldPw2rQuT8jtLt0W6fP7lLRx7/l/gy+arXRNAeKP9vD8mTK99JXNNWAQ1PUq
bYO9e9HUn1do9a/HyISNnzOEsoIICfs3ujyQXThg26MD7ZyP+ZJh3XybfSDf8lUR
ekzkOmi6M5tUV5GdAWNU1V1cIzqSPrFTFqEVCuBDCwD0mspLy/27Fjw+QPCiydjg
ACSlo7wkNOmQwGu+C2bQk3yHPl9qZZIGFAOO4AylEJIrcsGGEUK8edFgOSVZImiG
LXnfTR6uCv+ZK0o6UQkgmUVsIaUVvIUEA7IASpdex59J+3kC3OLMmcbNuNtpasVA
XK1Ao1QgaTUD4Ig2MjtAXKBGzkohGfuR/usX3WaZiZg7LHEy3VSaUwDGVe/IJOfn
tBPHUiTj+e//6qHWA0MYheHlnQBqbgPE1IBaDcBz728JAhwRmRtguBDIwrM0l785
v/n2tzjnKWVsBsNm5LGOEZpiCLOe5HgelltBDnMnblWwu0l6ZNR2TbEM9Ua3Nw8T
VbmRBYjVBm9TCkpspSsKhW054hlUyXZBYjig6iBXkVlKwa52MzmJdb2ueU2PgvPG
FMBxjA3Py4GLkkJq6xpEB2MxDz+h4bvm/AOqUOxfDl34lG0mbx84JpDPeU6DP1Xo
IKKSB+oXCJlSN5rixIxmmppEbHzKXK4skUCjRpzsmxbcZ7ZskJlMtXIyfBC9lfD4
zPN9/+h3YL9a2X1wgDF57b1BNavoXREnzB/wu6Ai2+6HbSCo7y0E5g4hzSN8yV4Q
wur6HcPVEl8PHwZbAwmNcdMi/ph1FgOkv0it+YeTVUNkjX4DhcLchDtnYzvJvdKW
REWiNzMiUXRXbOuXz1MLM4ZEz9l24EUGnztFGi9FgYWye5rhoihREB6XxXa19R05
MlsiCXUyB7ax/ICAVD8Kzj3JUhPSuM9AH7RfAef7UyITvOq5Ed9uE6ud20Qofjy9
DSfA6MFPJZE/tm5pMhWdFbF2s/LnBi4+zOkxCEHzjbo31/wE1tv34diVTL5rx1oU
qGSupPQT7teqqEMiw0EelW+lv508sQFIwAmTNwetyvLsNX0blYOYaG2tKXZ8omGz
c92GRgmlvHti/4P2sBfUKWzoJoupKRT6YjaDTbscmiyBUN5BysTkNFgU2g45Ftqz
+wnKC5wXvQcCREAValnJtLotTE1uVdXESgZgaeTf7WDBBu0EVSymsoF4ZwNVU7ZR
1rlAB6uU17Uzo29jtFrSx5aDrRQrLRrdI6R/r49GA+vjeLVz7PfYRMTBwdRhQqky
3r8M2qnAzxCc5jsIcGe+YT9ly0/s+GJXFQYz9NwTyokkGVrkrq+A8BuWHiotTzhD
5z7M2Yp3X2Q7ScKv9eWgwI9Ls9mFG7b2gjikotsUgPx/vU7nUn3Ct4MzI2HLbLLY
SSiYtYOpWwjhLIoFX4hsxKeKjC95pBApNXBs5xMXFVu/kEfBwdlqxocZMw8b3Ey7
A4AhTBcYcgzFrKDO53uzKV94Viu1wPnjgJVv1Y5MOBWP8mqSlzapBhV0lKk9LwRz
jjlyBsGriNO8nBQvKk2sk2gVIQgO+1a/JMKFoBuk/G57LHiuVMKHfCZK/6Kgqs8A
FJhjhCEPUiVju+A5kxLN06FtFmXr+PNqfArANbmrP8qaKIxa250Trn38wOZVA/Rd
U9cR15vP6jn6SLAEMmTtWRYb8N/8eD/W4bW6Ga7i0i653OR0AYcdyiYM84JHrqbI
/fyM7NIGE6I0FYjeExWUQoqfApFZrvXbl56nJCnsSEk2KImuZw0fvQo/0C7ZkHSW
RcPXUnPi9xBs7i2q3++bktjnHYtdcy+KQ9Wf7BnI31YTqmdv6Ydf+TcK5m7F1d6V
TcSJYn2uVQBpk0eHBSGnUhWW12Mu8Qppq68LlWX87ge3Z5nYlI9qMvpOm6OJptS6
tbA0Kplwopku8aV+QxDqMe2miFu7birbQfTe5WTF2gnSSBgtG/lltxsMcLCRGhgg
iSyQ6JeAGhqvIQgf06nyprVY3crEgpQZLuVSbWkOrbbl0el+OiNBPL7AZO3uI61p
fwj0W2/0Bjr3+WUNuiLDxvOT3FPAhWJG95WsvdZVUTSsUXdHRSlxBYzFFnsWsiG6
+oJ2uw3dP94A4RzNtEJ4i9ZL9NMQG3ou5akFef1EK2Qnd67pSSYsMFKD1OzzwbMF
JvYxeCVZXoi2J18siEME0aLEsLaZmXEbJ92uIvYawtWoiwn2yXKrjHCXb9Y9/Dr8
7ZAUK+0kHsw1zgsvCVwrAHwr+tbQdfvuS9eRVRZteoeUGmgzwp7XH5f7+ieBmB6r
kLRU2zgCHeVoAevK5pOyhfJ4LIne7Ayh3NDu+0ARCBUJ9seZeLW9jUt7cJhCY7g1
kUWAzn+UtV3cTHk7kd9A7YiiqKTlZbgViBLEZANlickW5hib8nPaDyLNKPmVeIog
CIUsfGZ/b4yYzmm8fe5TNTdp34BajlMQtTKfy90IfSyKIt/hdOC6mx3GxfMcebN3
qiYLKPvZfGGdTjDOsYdE323B+CDnTU0sjx3afzeIZO4yo/56mt7XNWkAYPmLhhU+
v3hAlpZn9w/6Q/HWmgQULY5/ed27xfc1gj6nygbKyQcE5Wmsj9LVsCLOEhuI5W/A
6UHhX9Hh9Gj1U0Db2dtBY0sALXdZT1eJaX3p6xD85P85gQAMBF8htaN90CoERPGt
XRg6twotFkiWz05JBKs6uteM/3VsPoaCPzFh782hwvYXkVVeVDK2P46LKsn/yeH5
STtyK6JdgzcXinMRN9uKNhC45BUWNmggSDjo0hrXh2IPrCFzEnWijRAzcbqS815X
TZ6pTnlHWbPsyZvIETPeWr3jIeQrMBK7mMaqLOiR/o/6h5TUlOvmMh5u1A2w9VlH
UjUT0nnwP0RJ8vkEOIA6miehciV9EnNPdiBK2zzHwjpj1yNlEQO4/XgahAyzOHCn
PLeVGW+TXz+biL19swibBRHXMp/BWSXePXz6JS7rcaOnxvc57nnop+2yNMej5Xv5
SHclwEBC8rFw81MEwhdQuWIHXpyCvfO8clOcnGc3MoQgR1eKbFLDREbSLhsE3CDg
QiN7mIbI7lK8jJRARkaA6KQvMcYy15cPFcF5cVFFiMQJvz//6nJj4GMPQpD7at7G
mLjfKzQVYoNXzKDzlP2/FkB+dTwg1Pu3qi5VnAICLT4kCQfbiLkobdVGNmUo91Ug
uAxjOFLOVNGK2oi4njedHMjVB/WcsB1ruOX5SMoa41F6pvbJ9uoPgr+dhf7s4cyr
XCsLFoqNo8B34N3dFomobhkQhboEkok+/qKQD7GcD+eEATiAa4mqP6fDdllGGxst
r15C0tlIJEAqAnyOtuCFdKieS6BSmn/G4Aq57bOpJkAiqWXsc4//1cYIW8lOtau/
e/q6upRn8yUjMpPtjaBglrUjwROsn1QdcCk4KP22cToUdrouzQsQ7gPL2YgbABSC
tss7mpSnc4u5jRyvgzTv3tqcqiWC6zog7fCdSO9tedcBZK5XZ0I+h5XYagW7FVXg
oG/KtDofkwVR5J/JudZxv7KYVbB8Dt6+ttBy2uqboHQIhWjhPnAzPHzaxewRGa/q
6g1u78UGilZVt+9qDmgTdjDEzTjX8+TzGaZsWz5l7UZZXqMnuImTTdjlr/UoZJJH
1lsLqIDrnf86Fwu7F8L4CCXm9iHugWS/29go2/PHD+5v+OqwPww3pvy4NeW2zfXk
TjY6oRXIvV8SbwK78u7Jkq2rYXRl8GzcBF6swgdnaG3ZpLINeRMZGZ3O2UAE5gmX
3ddQC9XG1SqpRjl2rOz9UIQp8LIRpAPqXbkNDX/AmY2OXJbfsyu+mrdqAVu0Wg5z
6mdvG8tKRHIFWrnZzAklBcsCI2Tacdu2get0igUfjVoiPE3tXp3CL8MIWBB4PDEL
iqzLoMGwDM7tYQrZPh8nAqnG+go+fLdDJBSq8sTKmGyJICDCAS8EC65X/g6hKsfV
ZikEAq2OcJetY+/OEfF8vHK78wNbfHycNJeLSyglsgZ2PIqXR6A4nNrhSc0NPZu0
XUlgDuABum3zBYLo66at6VglbwcF0Yu1d164HlTWqSCv/eVwhfbNe7Hk7ADFy/Zd
QL90eH523TFmLmohTmKDxDfIR6ugh0oRPi48wulhIWAV/h3ShoEVUa0K1SYu46hA
GimUMi+Gpc1izW+BnWKDCVVM94qnDldtd8arI+uxaH6TFp1kewpXtcoWIwSfzyHY
1sycPSz8kXFMI9cBAfNEyuKOIYNRPi6zuiUnqGq/1iXxRQUpTiM4Lk5BhzZiWfjQ
ythB7PZfR8kVxzBZbki4NeC9Km107tnH+hUPh9O+ahw4SFTZmEi8eRJBX0NDgqR0
qJjVjo4kGSreOcfo0Tn7mVYkQMyqCkvkk2Au/PVYBWxwKK9q1uze7EVc+y2oZ36p
OpZKc/NFqf87TuMWLDbUS0BWtg335/PKRuX9DoU3BviD6xed1sYBSq1ZrlUNJwzF
CdOPXkGsB02yI+Xzmh8gd8hGO3dB69x+lI7O7KbXzZLQqFOwUwqakNYNQgJg6pdt
VAwJOGhXrKNrFRG7RwF2QDrS6eLUOZqmq+j8lLr69kuNm8PpW1s3bxF6PElSgl2Y
I3eNXTP7rUBEuNI9wg25Vk4kQrOUbWKw8rR8r71GgmjCU6hKewjhCra+n2UeHDVI
qh0V/VDa0V80EjNbGxU/MATcJmxPUHccyI1pBI6Vhp7PxXqxijYlhgqdOiRsEQ+w
/dTk6t3+UQQj21PwXOwPrqDPvR41TOD585InSGlgamlI1r0QTQQfezBWiInMmRF3
CekxcuEJCFsrHTMycgZq+HdZX3TLicLYGMMew6lOxSXD0lyzjKTuJTCAQElyDUuv
JtipoW0YJ3RvzR6qP5sA3Xr2Ea6TkgCykNJCjLwcnNvlc2yFUvKLvCaktSFpts+c
GzL2Eocd6vRGGHYifcOoUeBciDSAEmqeqzfuOcC8vrI80n8kZ7c808Lgni/HWRV5
nVdFjGC7uBBLoXpOoNWV3N8EPW468YqkXylxrDd7Z2mQhlYZCiWrLir0v1dsn530
G5w/Ja6O9LdUG98HaRk8mK+zMptINqUFDkrB3j/1qLyNXkzU3RiwGS/vNmyFbGlN
9yZ6Udb33G3F1SVvMKJLuO62cBCgqDdPlLQ9jQv5omxdIBQq275D6hYcXXD9x0NH
RCoYSzOTuZ54BTIVFlJg/8sljdWY9M9ijAIeYVR4xet2lHK3gW5JdRvf7ClcxL8g
E3tEui1m9Q/12oOrvywEyVQvTJZ0k53wNkKskblu/ljzgNGpiE2Jn6eBjo/xX0t9
/BDB36mfRRtMgKV1IX15nis8IwYjDWBVLz8k4pWGFOymTODYDsWeyMw0mzDVQ9KN
T0VygoP2w/bSzaElyfdDR+J7Pky56b6P4HayfSVnHHOBKhr05tT+GV+FyGzKbTEI
O4Kcignt9E/HjqePLAS5qCbjq1EdHftCny6+xpiMv7oeNz0pjm1hOJoiCi89Ticv
pui9RfkW//feh2aIUrFZNOBwGpQ6+rG+2CCifdkU/OK8JxdnkBO/4pYgt2E3IWV1
cQSb5pjzOqV+MtBiWpCRr/CVKwpDi8w9s+hw0MN8FcUuk0EIfTr8b18UHSc3aJul
QXfAABY7nHN0QH55r46WN9WHuF5gDXemGwblwLIlyxDinRrVyZUO97h+EBMvtZAW
c82pN8SEwOQasLUyDXgsBnsSW34KNHfeUbJrg+z64GEQJYxHm3aTsKuTX9AlFYw9
RygbSYQl9V60PXYSh9hundtxZz8XxRg9xzhoe9uCVGhCOaWeVcPtz1hdJ6ZiodfT
fpdglRkBJ+JTCJZXflIYG31Q67yc3rtEHKQh6rs7VihEKy5GFkee+KJRMcjDx592
kBU/bUfN6Y08aVWdwN1R/rGKt1UEXj2VYBrNg9QlP0h1BhvPW1DYCOOQ++13ol80
FR5LlbVZ3HgM1jBTqDM9jZuTWs0DZ1cKHlxHL8Y3e+7pUIb3WCqtucMiZAQYTX13
ydDrmpdY23nIc5o+1+dMPxFm0hfDDJv1INsJaQP5E74Fw+t1QtUuPN0qK5Xforzb
cEy2QLw2L/C+lR+D2Zu7tPniYSPRseV2B4VU8kvgLkF8iLVrymfM1sNq0AvNm5pz
iEjNBfppAWDGpmoJzlwVvmgZJ/B9jIf0zos6Hr9j4aKwQDp81II07u4H3MCiHuWg
PT2/D+y3OxHYIviB7lQf+XvNKPnLf2mlmIvIJNRkB2htMYM93lZZ5muaNr1ied1n
kXqzMlit5yO10nmAj51LP4qlWGec4Fq4L+h3S0rC7jcr+AL/eH36ycapkSU1FSCS
zSRfLdxeDiPY9tJfkk+HZ4qQbUWA+xPUwcLVw1IOFzh1/MozOge5o1OFeTuGd4pL
ZDjsnuzCekqj3FQlFYqn+5jU+LL4Qg5fFwLt9v+Ywwi/nzkwoFZLcECloKJJbrPx
nruRNmnNZOSeCjoZ9RkNS+Q6TNfEVUvHJ+G0iVq+/EGcCUoQCk6HL9Qt5/Ezx/oV
6SZdfDhXWoMZH+gLYXish6SpvncG1+XogT3iQe465tzuvmpeScKzfDyvmPVvY5d4
h2GbCQD1+K0uf2q7VfDfke/HH2VsA87FSoka2Aj/j5Sf/J+eZXlB1raqlEuM73aL
6VHoSwb7CcSXVpJJXiG0Gl2BmIdvOat9VvHC+PgN3yVUE7SnCktS2e6IBF8Dzvbj
KL7jtdskiWQpvCq8eXFkfArOc/xMWIYiZRa1GbIq5W5XI4rIpcYI7QGHUDbJXDGF
tTaItpZWEf3YAQvPOEfybdDJZJnhOVzlnLEGMm+cQH6I/KtawiYTrAKAQSCE/CcX
ny+U0v0Wn4CyFE+OARVVF+b5Nbh19dakKiwXBlQno905eq7/gT+oXnp9VVJ8ETLx
NzRDBuv53vBsaTml/Yj3/9vnOHGJEkljkRPV0Q9bbK3m9oU7D7Q1nfc7JPt4AY+2
fuZTCw63/s/2coi2pQI+qnjmCjiGEjIVjdlvFN+f58Mm1CHl13BBGVYMpBF+K9lu
Q8VEwooqpnuiFe3B4yd2KechstJU36VoLkNWnCeUleVFMig61tp7wK69TznvJQLb
9lHPDnRlck2bIa08gwDpJu1Lrh2Iy6wcF5uDAt3xvQoJVLSDHPfxaIUECa2FO1Ri
dm2eDyFGYfIz86i5ygMQRFS+Y7EYaq0/VtImjLoTtvLx9MBt2Tkqq2az6Lmje0S/
CdOKqUAAqAt8hI6G/cnr9jiUrml5nP1L3pYqR36+WIK8mDc1DYBRSQmVZCNsS+N+
jrmv96BItOrROx/RoSGA4fmEHXHV/+6jN9/fqq4pNFPIxdYwiUazAV4xlm3Yv1c1
kiqBtbi6FYdPAii97rJSg1wqNaVNIrafxhndY+I6vHWtAk1MQFNllGwccc3e55Lm
uKC53Z/0ScKoY9JV1ulPAglT6BMSUP4DTOoRo8qI0HD12dZpvOxmfBeg4cnyEgma
h4ryWKZUrXv2MbF9oYGGTI/cRiVoYXAIIrh+zijW9IuJPSjzHPGbx2pYmVbg3swC
uUUW5XdTJWSqvY1OGsCKL/2pnCbthzCQ0OHWgvlkp8aQbNdjTNbtZG1ERt6oxMUQ
nXOyIwZnvdCBV0bjvFKx6iD623Oz66YWM7Dra18T/lkYR9IlK95b05XS/dGKUY0n
zO2HagTKppe+LB8TasRaQC7Rxv13bclSjrAQkdRXSBSdBMXWRXT7lb68ogyXVU+g
Y9xloAeIdqAUfmy/gxS6k/rxt95mzGhqZN8IzPp6+wPdV5LKvZ1gK5ZbOEClWBI5
8EvgpX6S3XtCK9TKQsEqkQoqvqgjEasHNp46Ly6D53UVyzj4nwfxsN0hXWid+PHd
HLJqjigijC+YvmE6eCuvqPVYr3rM5DVEBIeZEZ8DHlSrdJPeXlThzZzvVr39Y91X
qV+uPL22MQXUVuaTqfViWS8j8zhON3TJD+t/OJ73MImnGv2Hbi7FqSkCphOxi25s
7wdxpjiEjIJ9WFSmCLKzAC9JeZQjtb/PrDT4h5zxsG9uoH+zx/6KYk4y7IMpUnHC
JjBG3uZNwQ8BymDVmhXcLpHm7Y7cTo7n5pHaIswlSI+VMaJQX6dQpdGR1tCqTdHT
KxZDnvNaWG5k/THvBaa0Ls9VnOaYFBgiXTU++3nF10ABZenKE2iNgaWnURW/i7+W
kUW72FiKPFRsPW9D2pce9vPNySjtgR6Z2Zy7rzhDq+dGZ0SbfsbFpIGWXSOpED7q
1KLyiHcka6/hjhzakuhFR8Yr7hlCoiZOY11ZglMcml0fNCn5uvCgJM3mc4r7MvOE
l6bl68ZscPR9hb5NIOzQZyd9Je+I2E43lmhct1R7SOek9EgKoFIOAcLBd9X/5epA
rqJlewF5OdQVarIqO0RMgQrRb6wXG3aIFyP9XFXdggPXb3+1ANzIAQKrFQdFfVo3
QGTSUXTDGbLZrJJWdVEn/WUzmho+41Fhwo/3N+Mp2yCXrHWljVQ9qdc75Hv59M1r
zTiHTffSZkbzZLsed4yRzJ5uguBQf/TNg7RVUdXCKS0+E+Bnb3fKlmmj01TvcUAJ
7ZNP8owHKflkLb/+skdSLcUS4uZ3lg6v/nvGUoiY8a6pvO+fxGvx40NfzroPaD4E
tb+0TeQ2SJ1fg2dEiT7upRp+7MkqEf80fMYR4R7PNCDMOhXgv7tnsdGTdFZ/mMxs
k9UiVJb0e2ttBhtQNUaSw5UFAhUA84U9KwH+cKrL7nt/tZSTnmCoHBFb+tulUkl6
vzVo6rRXWY8Uy4OHf48DdwEtHGm1sVA6+U79K3Ia7tfhJNQrenK5SKRYT0VYOhz9
HhXNmducnj9ThL984t+Nd+TDnrdePNuYIMEdti29chtN8zmH0QwvTcxleAxbU14j
lVlQmHnBwxTFpu8k74nnZbixINrOc+fEmykB3WvPR4r/lggwAnMWEytCbzIB/aM6
Z32m2ENPWKD41TsD1er/ETVJ7ReaecWwUm/TfF8P0EH73oht8VNCO8VU4YBOLB7D
Gy9sygN1bxCwc/1ok4gw77oS6qgzF0znucokEkiJiEI8PHl+MqacRjKsFW07Qa/I
Za8LuP+D1OsKloEeQ7mG57nqmLYCRNSW5E/jTLyzOU2bKv1EZxef3yvTj3cBKEvJ
cofPL2n4OmZSdlhsY2Be1SQ7n3s4Qj0qORALnyPtVH+YQm+okiqynT6Jr46vT6uw
UzsHkB54dPrOfARxveXaA7aIwC1MZ1smzh9bgWo3mKWukwcLX3oyHA1qlFMtdt/M
IOUhNLR/lI34gqP/QuAUFe+bS+a0xHjOIwgAHtp65hSwBJixqSnxy6j+7aRjYIsr
jHH2W15+jsiAkt838yAd+NZ9/5z66O/0duyhpzkz6AyicZDQ2GD45XVXYFuC6dye
SdWajz2o0uHopW2MNk80fLtKCPxaCFJo6SkiNOqvi4QGu/+2H69j/X8AsUVijYX8
64bd05QD97RqFBWh+eOkSdEuDuyL40uYr0Bzc/S9gSSBr8pzHm6XIDlBtpZ0649U
Vi4hGYNAQobwI0nSOxpe0Zf3rW5h1UXI6I27HQ/YuXxnv/1lTsh5wyKoVZMD53R8
2wKtGePnGgHyJ1Y9Wdsa7wmJQcNc4SP3PnzK7qXqad47v5aIuwfCY2CaNoUCmH9f
f2lQa3aVSBaiiq/OahZMRA465UG2yuZMLwyFXzjZjyR2DtOzVMr+gpdqm++Lx+jy
EpKgEvBs53DL8oGP/q7hD1aRIUJKegUxA+ALRRLcbY5c3P7WPf6G43wT0o8bB7kS
pKiGlq9/vHvbJmu5Pcp4/GC4s2TDEYaSJu0Z3Fhxkm2O87dIUkKhFdl5rFGgp8ZR
PGYYJGPd8odSy55lQLq20xA9dT6CvKTKyss6J72GjFFyY228mL5+h6NjlG/iOf8k
/97frQO2d27iKM9XUffeIFEweDtWj78K8BpP5zCjYE8OSlibEixo4EMzYfbBlc43
WrV/M4UTzaIQZqGwnB56Hmji15HRwkta3wp7FaN47x/zMby5vqVDSc/KznYGITqy
mI6yL9HYkFuhVhk0XdhYS5bR/WGMaMeuk7rMnZ0bebBanVV2AsrjccYFj3tvIXm8
sBsJzDpRkKWT06O1iaLoQHwuN3g2AtCe/yi1SkO3SLmpw172FFOZ9dPM/fAUDIIg
5Ha9WPloWjLRyPIwPpQOvPUKzl199mPGMiPBcsDSPLiI0M2icgmJkZjF+lLEu4UA
Zfgz7Wym/Cvdkm/AmJmljq6slLufNOwj3HxmWr9h3uSZIqSEdVzlNRIC+FfZ3zQJ
TIi3Yiyrzc8dRVa73jdqH+ZXKJdXPuEmAPJSRy7lxkvdoE36N47yt2TovR7D60+L
pBCCFM/5cStkrd0KQA7iBqmv2TPjsJmsXBOxzrs5k9+5T2AFAfFiVftlIK9PT06C
YLQIAC2rOJ42uYOpWTL8uCXxZ8xm5hRAmOI/23sibk0DIG4dic01t+s3YvdrTXU+
IwoFMWI34w6HAhgu3iw++LLRyDP9wXFgq134VS2xbyIOZfUBEiKi/V98BnSzCqcs
HYEGIJi9Tq0rjsKryHBhbfXP/a0mcS5nRxnwNtHFjha4UrDiIwBViSqVACvdmBVm
LSfuqNB87+3I9PlphVjnYkGz17fvpcqU41gAG5JTXYiuM7Rk08kkIYGEVYGcj2Vo
TMWKGFFNv5szovUdEQgg6GOMUb09NXeDJXXpa9e9YBTfZv+gkrDql3NYfR12HXwr
bOaQtCj6kK2jjew3YvVEaTN0jm7wI2Omd7WhFGeegBj9EtpCwGGq0u067uY6fUKL
wgLEG+yJyANb+5xRHwwqTuaCNr/Q2kg20HFdkpkdgJrf9zq7qVUmOkyb/BqvF9Nu
HR0GmSI3kPdTHDZgbD06/IaVFZS/EMb1SFS9DxfSnYRoDFOLzPsdHUhjur8qiXtY
9TWD0UGTz1NGrzT4WbEsYC7hiZEnfafVVBLKNjpALosQDg8mhng5LcF4CXKYY8TU
oAuP28jIcs6ef1Bfq7Up+D1FMn4SRz8bym6cK77TN7eeW/msqzolktIyp8wIyWMT
jjYIKw/iYscYSUFg5i7Dhqbg8fXTwhm5XBgnhEVKZNz1XbRR+qby15uoo+XeVmmS
CF9J3wh9F+DlK3l4ucx658MOLVIo2mIWIsgcdxJDfzT8FiT27z6bFvfV7gDyPmQz
2zZ3rUKwkN9LhkdNZDyfEsEx3ZpMPClVXoc+6sYNV+gEW+EY9MsN8qdbamJ1kxSv
qd19ZbqScoZpiz1oMt9P9lpKN8febNik3whnVnRXetzPCebpS+fVNBAg/4ERNang
XZ8EfOgtJWm0aFTmzcns/sq+XQGCyZ6iMVSwdX+IIF11lbDL6rZeMnUHeUd4JzKv
Mq3vO/wPf5K80gzvy3PdrWQPu/D9GTP42ouf0aqw+vFGYmOa0QivDEY3BbnnzqlC
Ar182oZBcMJdjMB4MHlay2dOL9dwN2Ic+SXT0a8jpYh9TWtEJslSbybqdfzaSknu
MI71GzTYJaZDw3UEz8Svw81jEYqgfE4epTOjxLCCK1KIIuTSqQsF6coEy1s4xqUo
3C/KBiJyLDYHsZoeNwPfeOr71OqGRvSGjU6AFsOHbjYGddq983/RV+xbgf3CcH0k
tQmLUZb0F0aFYlu10i9SPhpg+lppKwcjjt8tRHLRKopRcZrKeHHbYxYLNlIHu8Bv
g7If1lQ/Co4w8MuxEeMCB1MVDaqCMJ+rz515BZZn805QkCutAc8NBjADvltszylL
01mwpQzvb21t/Zu/iJlgUCHQwzy2yocy07Aqh3KFOgXTxvqQs4QIZVlmkXv1BZ0q
QH7tY08lpQ9axI24ektCa8GiNjb/en7MJ6Kt+HKVB2qPPpy3oDH0VnbisgsP4vIi
gH8Appvhmn18tjtQYPZYMdiMLVhNM9fij0rBulgeCGrvO4HofBjj3tOuo0viMSCD
LQAqxhUJNyNEHE+ah2u3VzGObtEOwUfjTrjfiQlp9OWQc+kO9/vqI1ufXBeRvliU
b37+35COWlYkw/Xklb3MbXiWm0YPCvxrM2/cDqgUP1ERwDQsOfKoGR6kHbnM+Ui9
ZhfFDae+2Rv/zJvo+SvzjU+OpvRXWp9p7avilNZikf5yMBlPc5h3kbZYhCf3+iv8
wOLVv3ervScL3tcXe+vrvrBJr/KvPNJzgJxomILAWpH4ht5ZMJgI58yWC3wV2Nfy
b/AsmbY58hgZP6bJOOLLn5eTYn+skIv3AJvQJ/mbfJXI0efJ6mVadj5Jh27ikkbO
D1NXtsehLNZWtTgqZ85Cg8s6fD8mxnuGgUiNaMY4GVHynHMbQ2o228XYcyEiy40u
43IExPs23MDOu+qVpQ7lewvQW0GsrSAOz7C4NUpsozgm1YlbFC5MqHSpAihjVFOd
xpwA/zdzNcqPGZ4u6kcPv6w7xsXMkL8qmqmPC3Ov0A+MerpE9Ppy4YkNO+qIRJX0
CB1o41V4C9fEws6e60W45V4NlqqRG0DlqvfQpfDO3rLJ0+trX6XpFD0Qqp3DO7pH
DYU7F+xzWOHyaBh3iBWIQRpd8Jvog7FyJ/X7uZR4Hlb2XVr+4F+HdeE9yQLyy42i
/JC/FZlwpCOajcMSW149YOLtsRo4MaQUDDY6l0Dpi8fLUL8ae03x3+/iHLPrpIQJ
HCggwyP5dnjwnM/Vd0NmZmH1LX5knUGASut06C+8Q0oySIAJ5GUFRleJAS8vCG3n
eOaGjwEZqGmbigo+MuQTdc6K8T5oKZOI+eh1VSe9n7Klb7ApUb6w2EOuz8oTq3Z5
gY/lrxXxi+mbCvP9RrQWKCH38jECaAxBHLma98vnS4MUzn4tWBtI/1T9t178cVet
VyvPl8XOH65wADQnZzepRb5tSWcr2EVO+qAnsrTdyKcPwjrHoT1JynbZJ8JERzfP
LFpZhuhIEvMK68hB88a0YWd4Fvt+QNNLH6ABNbc+qpPu/vnDjVV3e11lyfwrB0FN
r7+3Mf4Zpt+DHztbuNvamIInxEpUZ5ul//Lx9oO0a7Vu0X3NVD95B2inwR9yYbbp
loJIY+mVdW2fpTklWJtsl9jLdensrcI9YciinI/z6/MFKCBR4+3jkHJHOBKuOLz7
FM+285SxPKFOz+iVye4TTxPxCBMd/XWqeuS6+//XLpfTpfGdseqGz+jA1E38Njw0
1VCgss4tbIWRSMlOzq5M3sHlsEH5rWl+v6RlxUvuFtvQtihxD7k+PQVEaHgyJ7Tg
Eoc2CEViF8sy/Ucrou8iuVE7spHfuA5YXw1fYlWh0YJr0ILAXmzyM0r0nCsQTbP0
hWFYAv9VPrrl9dMaovScKIl8VcUxBpmQ2VXwSB18k55q4R/YjEMP2IOQ4aqWT7YH
LzJ4lG9WjltWEKhXTZK4LECPEprEW+TONAhwkmFCSM50ihJgkpZNrxd8SH7kwMa/
SU2WiqLXf3u+aJ1nmfYlYvZUqrQtIWT4FZaiZv1KE3YImaFOaRfXlOoJ8AdgDu8Z
PVX4q8abHHxhnh8T/StC/7mDMf9kwuEsBK/b/lWooQ2hsYY6h3gSqaPT5fkJV1Np
hMPqhw7WIyMWcUktTy7SKvQMj/M5WUNqyKwcIdwkP8lWIH93LLlu9JtAdyT8tPxt
2fltlbaKlg21h3yBVfGZS2XBlbyYbbTfQyYzWJ9UbkPjbn0cNWnsrKJ75dYi0fA1
WMdqvbIyEAZv8P/TtH6yXvBdQ1mVLIAP3dbQQTzRQZt8RtEWl+ABqEy2cpjQNFVe
fTzu+ZmRkgXp1YziUy08zdLIdqj9ssuK++tRGGLKFAmzcOEawbPbFBravWncpNdp
cz9hnnpJUtP0gnmRd0L8467CEJzJUlklrxYoXFTLHhp6BOtSDnPG3u0w2g81O5x2
jBIUjQSZRkdTlIzEuegXLa/CSAcm41KxET3j8MnM14uAfj2KQj07omusOUDkveaq
zfWU5/G6cC4QoPxEaCTnxnxt7tBVO5xAPBSVg3vO134rUlsxbkk6OHN7vm6rTHc1
HwvCbBT66Rp2uTOhJ5Tw5X3Y0BX/9PSxMggkfRHUvelH2dZ/YAFczyBN3OWrqmni
GVTj+WwzxEUfApbidA3EJxbZdlAVZtr+tvED7AhogBu3tUCMaWMiPVecblLhrlqt
FNsSI4i4QZBmb3V5u6yQ3PWNkj9GmeuG9BoGvlS3nxC5AB751c28W8aCgjiVtR9d
DTI7PAiqtwsWkpZ4vhFEwpIMJs88fWsxJl/S0tkorCPic8CmbFrKuNCZGScQYhAR
nMeGZayg3GK+I+atc2FWJkWyBkiB7UiHHmUGavNC99zJs/hqCCL2b4pxJxnShKRe
w7XtOeDQ/sJpbkefJd1lEUmJiHDdXlhqwiOqqR2ROIFQ2Q8yoGdGfsxaANP5c9j5
+5TZXxsAyi8BhCjQjzvU/6YR/nWiu2lTLwAtjThR4OLzesoCNTtgfzFfvBOhV/qn
Pp8Y+TL8rgwC4EmqsCyUY+wx0Atgdn+QLg82eVYUnO2ufkprwBIIaE7ngE+2Lonl
ja97n/K8/gQX3bWN5DgqjAW9ZIz9JOjrk45mR8udicHitRurvhiuScWv7E1Q1kvu
wYt2HgPWiuzHb9nvZ6oHfjjdN4M14zDibD+jFMSNOD3dLAmAkCFTEmnFlyt+5s4h
jymVxPqCbAEEI9+EfiEC+UHai6En04Jq9FXD89ctaf/en2bnBr20U6z2SyRT7E04
UbjgrWg9k+5qyOI0sg+z422FlmgltT1oZ0bLXGbtZXfZ7soNrbYK5VvNlKlRWH7Y
yhDvJh2hSf5FD6bbv/Jipmc9OgeaGPSNtP/vAa743pRkOTerqbiJ3ulKJvTLzb1T
DganWlrvXYz5L6rwCA8kKStw+EViEuN6sjdA+QW73xQMrq2XrcN0jSuRSgcPjhUR
4A4pnl4eCk+0XYnlAfedjkFgyEVyJZzS2kdMvZltUa8Zhwgkgb5kzvgPnQHKJ5s8
sWwzhHMsEgSKT5X/1y6cFQ==
`protect END_PROTECTED
