`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
0d8a3CXA0O6wK87FytDc8AiCY80liKPuf4AS8cgISN+7AoO6XqnSwH7Qh0xouF88
Lvg5YBK08UXm9S05rMWT2ubmlYcAXkOO0aJep95ULD7I5H3otFwzwGHUmqo7ISy1
J+PYLEteQV8IfdA1sjPdqICOvI9BMHQKhJkSIg42Uf5eB1oh0JCg09oGizAx8PWN
DgSnosuapcNQNKJ5PgC/aDjG5MYo0uvafKkiVnpC7FZEwPLda8Plb8Jtn6HKzzPk
ZPaWIqRxZFhuMfnE1bgm9NgbOup5h0BCeCGnHGkgYTHSTrr758KmWo0omMSz+yVy
M7AbrJc1OJuKXWr3VgzBkdINZbrKr2hKBVMgfXTJal1Dzuj3lT6FnxPnrRwiVFm2
rhdb7mLEW09gY/b4BmwUfptydwuCYlEOOLrqsQ42LCRXbEsvHtKzCraIq/F5vWdW
dO9fddCpCbqLCbDJwdIkq9O0Iw9b/EbzsJ9e6Lp7Ht5r7/JYkJr7qo3fuSybjy35
+Si+NB03Zpc5BHZL8I5se4h9KHy/MPHCnTiyDVDuDS82Km4oJH7yoAUWw2HaSGkW
hPhlyd97gTnmdHTgm/tHZDwINh1xpWMzC2GzA+aCDOhCPz3A8o7FY6WEtddOd0Tl
qjVeCjWQmR3SAdMCoFEW8GKY4gbsc5wxnAXqV8CeHjKrPeF9h0YcIkZGmRxXKTfj
bLeeLzQL6muu/PvkGrkzG9CVV5O9gXzGTTB2Jrq7eMkNE7lwEOcQr4uXA3Cx95ph
6hDnn/IgdEVgvnmHEDuqrLBAqhFRSI77NZrFFbQrcZr6ogbA5lWTfaTFa5TQIAKH
qG/aRuVI338keXRWbR61URcGILcqRXWp23ALfRd0Vzs7MdW/T70LxM5FynHUKjoI
/FphsnJQ4RrKskZmN/W3RIHqd365qj5u09cgZA0WM0l56qL+dLZnXftXwcobFn3c
jeBRqsNniHUg3e+P3T6YQ+F/SS5eHEAM2NLOwBMYmnNyGtxmjIkxhY0JXsRP4LdY
ua75CYiEx3IGmUExenJR1ZnFHruVFW5oyVsA8kNlwqBxx1XxrR0fOvyTwdAEA80X
yOoOfl0cDudZZVdaclXJ36jVZKu1f+IVeTKFSMQafaGUALDTAU398UtEa9nZJuOp
GQrFD0xGMlzingCCqa4NQUxnO77lb10lg7GiKlLRxTblD6+hfkn1/zpCSkZmIi5r
oN4jkFxgR5+USobAJZIoEKVECwIg8yKu/khSHtwB12UdWALWc7GiJWUE1pUCHWNu
3xH4PiMgtsiig1fRLfiJMV31V0EPtQQsu4zJ4I9L4VcsXSuGuFKXDAL8/FkhdtJr
k5pqnEZMjJYkP8UYPj9VoT4mU2+xc1lScOBf8LmQM3sjzjYZHTYNfZA0rzs1D2M3
mthRzUE2S+G/pDLFDZV2AKnuIhxUhTswAm8kzYZr12SyabDou/ijO3Jth0POQy1l
Ag6cwEfz9I+XMLNlMNfKt/5sg2flDzV3Mo8neRcNZynDASHPKDyfvf2aIVLXdL+y
A5EPGqPA13W1VeoQQfObJJHNog+bhUe1gGKqP11Xz1ztbih6XV96NPt05VGfbqoa
mybWiTA+T6X5nvmstmRqqbAoX41nH9+yTIct8u0XdQR2hTEWKrq3Hbn5CoHyCVa+
5uZEq37hrK02ibNmQi45IFrP0h53jpVn3q9pB1m79XTWZnr7UusATHyR4tlZNRUr
snS9LcUkBXRQs/dzNcevmnt4+i/s747SeIJpe5b1pBa7tqv+ouD5fC/HlF7BqZXu
ZgWOwZY3Hz+boPEzh4nCa2NxJ0ZE+TWf4SxF0Jk0m1S7JarXspWGoU/v5Ws/vMPO
djV7WK5UTN/gqSvuXernEmUCmkWWAQ5k71Z8xYSQxw9F9jIb8PNwsbmcE61cK6A5
0cUCs/6p3rlT+OtSduutqCSeyj16rVeDjFE15QIAzHCKCiOCXGJNKsY+8Bc9gO3M
R2I77+L5CoM+nmnL98SjU2DKkGmKP1O+9zBhCfdKOraYiQFbeGRLIPzuk2CNKPWv
Eg0+yZ+XYlmX+82IL3yJI1RejiSWfuVzPJAu7G8p9DMeE78KYiJrBLiiU0rmRYSu
lQ1w/V5+IyydbJKnux7VVmlvQbkJp697LK0tpdxMsMVbe2o8CR0UGwH48x2hSj3S
EQHLuBJ3lQx8prFUImVabrJz3MptDgPuAwM2/U7AY8Zgm/kh5k0Dwk58jRUQURXm
v7xjXcFHnP0Xw0brc0ye1NySmXoegP5B/i1re+CysMRIjmi0UDW8a9ua1RwsooRS
en8+FckQVjvTzWCh62T/ZfRa8IT5wOBy3lNf+D990hnsX/oHnD1ueOpdNl4VMWiH
WRm9I0CRJc9Xgmh9tsGeuK2s+UGqHVcmVkgDil9mK7BBHjeCQ3JbBGigmrtOEy0H
WQt4x2diCBcaoJrv6pqTejzcIoEAtjOQwdxNMiK8tJJQY/ROBjF+KbWO1unMj7Oe
r3KuiKSNWQCD88UwrHpGL4qNfKLCfYbCp4hsVml/wKJfZiD/8NhU2+Tqpm1ePV8X
naFj/kp65QqIAdNFwp5j02HW9NZ5AUV1vKguU7eTfRd52WBGuwwSunFesiguPg0P
x8NFN3F+L372cbtNTQDksegFynQOV4ODaxDl2C8xLiZDiz+zZ6HpsDAU4ExMBYAK
6feJ5IShMIoCrLT3ADegRFGTrmRqiltjOUQiqaPKirY0NiCJ8WFBzBLIdaMlWu6/
ScxIl/m7vsunMQWDpZavpy2hSoxHZhNNr0xbBVzW0JxVHC3y0cTLuwugiECnFE8L
LpqHLh+s0bt3zy3U1QviXMBlmzSdpr7KLtwQxmfRUL9fVNW59vAdFn0YxzT0rhWR
t8nHEpWyCu2Dtl6BvxxEtVJPz3qnAc29tZ4O2b8kOmpb/cFbbIxrZcbljAGGH6bZ
JVA5f3v/YWWYjuKstgwTMlxpwEEp0blev2QZV+MB+yQgy0ksoai2z5GI5KACUVqG
xBjf88SfxUpYlOYjSssmCwjsyVfF4jNOxOIoUnMvYIDqBtUafO3ly/iDWew7tu9j
WQ9qIktiWhfK18tf/RRb3xzymnn7hXzg7NwMrqBq6TI/UmuaxEdPKpB7YWKhO4/3
JPtHrvRfjLaSElHXS+LRsXlUqgInrqR1h+HmWKUHpzSsNvcftKZFfsiGrWmCcfsa
U/KmrJ2FDlGQucJrIgAEsFIA7I1/QAhDdYHHx3qwmhQBd8JKqzu11hzUVn5aJT+4
WX7qhFZ/+JuZGgDlb5CR8wg2Z1h5x4VAQuJYI/XP0j92jB5LXZTQeSrCjBHObHPX
5KOGJOu2/bbKzk2RbyIrm9nKcED2sO6iRHIhgFJmmdyHXgLVS7O7kCZO4/SZAuOn
9OMd7gtBkDZT2gGgyMDjeqgr75fRKKiXMrZyT7Gv3yaLgaeM4P3eDV8VzCfIkDGu
efImT7NRwDb6DszTdeqKR+3jtOwXg90XXNJM3Fvs7Qgm33GNpVJLrNFhAa2SQt5t
t5A4uD5q/iEVm3+duA5OYMcAWbYXAJIwdKdqAvYc5CJ5BkMiFy6ZeosHfhFzF5HG
NSQ1wTtTtRew11uE44dGkwuLFuuzO6NRLXllLJ3ARXLW8bIx7IV3JO532uZTfs0z
H+ALOs5I1ykLZ1RX5t3wi3OGNEE0aHXa8slLnbj7iuek2qjiMjiRbKn0+X5CXR1o
IfGLVlfJY6N2G8e3VQhSmDT51XrwT2UtWM+dCEA71N/zioWgLrgRhvlJ7oKCiVfs
wUfts0y82gaai26UlEa3CspxWMjVW6e5c0Jswb3K2T5/v7r9Ud0ZQW4wauBe9S8N
mDrMdmk25286bEIlFWgPnD65yUbbAVUeDOBGT7OH7cbF+O14JtsxZMoICXur9ytq
M2lFpDPWVIkDvj0yK5/DyBMLeHshKHOixjbQye/MWalnmQvUIRQZ9U2tpECGmU9G
qgWTdEJ7BPaUeipbmGaKuIDvvzE6cbhcp8I3sj1UYOg/cz3kNcQwcp13vT/sl4gY
E0aOyKKaU1iOUT0a4KpMU3EZmHErbYMDjIBpEJ/IFP5wbnaY6CffE3g7L6Imm9om
V/TAIgjVevT6cLUAXOe6Cr/+7RQT8VUAGi0Hx/ngaOLpYHCTOddrpk5BD0uiV5gZ
fnzaFognsFbOrkrZ0eiPU9a4zyuZnT4jC+8QLL+zP1x7YwAGdrcecs70WjhJ4HKU
LGrHGS1x1NXxI0aQm4HXND4QbUt/4Jx22OSGmBy33MAocN+IgqwhImymDr9Q5PZo
tuOFxjz2Tc9b9udWF6frVXP9iKRpeYCoEe3YPr67By1AM9zg5NkoMlffeGFfZ02I
StTwPle3zP/OF0L2hVEZ/+lq+7vQW7Gqc6sgwEaxeRqWmvNub9AAJqQ5zaPZ7QqK
OHiCKB2o6iS9Juq1NE4M5nLCwcAPkk3W1V+Jx7/HXhtI110vC4e3zduPTfqqkpAq
2iZ6vH8ggDzaHG6hObOMD1izMQGGQxTSRPLBolk7xvseQ5a531Lg4h/Cvli24Nvs
qMgluK3Rxnqh57s3tRTYker9SFRIMa/09Wa2pi3pavqal07Uc0F8wHTWKIf6JZis
pD+Zs4jszeKBM8xgkBXBPxHtDH8iO+KV7/ULZcuLyccZ6L427owKEGekRlqRzgTP
82XunzkKkb7+5yd/Z7s0KIfuIqPac1A/HA+ETTPduO649sIxQ5dGUy7OZx8jpkA4
/68xUP9uGxKn3bUEhD2inAD0IcLgvY+Ua517cZ1cIQ62qbe5KczJNBxlFH7DaJ0R
PuwSgpx9TFQIDpsdhJSwUjBBbdsrkBjN8L1dSETmHat8HYJKiJbOa+iz064xNQgq
8XtAgeqa6aoUZBOhn1yvR9gE867jbEZhJPSFRX9SK0SARzwJhC0YT1JMkj4h0IaI
+HMTaax4GsziXzeOdCnQtg+OmOREh8P29ftxp8DyTH8OB2U5oxzbYDqBaNn1lLcl
7et5CpENKQiCFEYueFTu6/aZSqb90fn7g7ibD16KvQx7NNwfYqZ6DbRfM6ryJ6dk
bi8MByH9u7qZvczlbDLODPdnyDbSrz5mX3SiwGn8TklflV1GTCj0D1YepvF/6rIy
S1j9NqB2Y5zrE+i706J6Pm/PIeViGYyggCTImjFy7E/nhGEz6hP+zHvAJwlCKWh9
xFFklgUoykyD3ZVNIFma7WXoRb54o5v85rSeUysEdn0KaVMwnbjJDViNzb9Ah2S/
1qQT/l7VdUyXM7PXUIqJx4vieIpVrbhSDho7Td/iVsQNXIYSnQPlr1sO6AE/tc+1
xAu50I/UZlRpHCQV1R/4LF5TB6bsKwaOYBA2DY4sXH9OaLeWGy3y8n9Ly+sg1nKF
/F2xImJiwKWyCaNxxw6PCJ9+6W9JtexGcJDuEFp/iLyFe/lbGurKUFgFUJfdomqD
6UxiYgfLi0D8Gck8T4QchYkCD/zpNPAc64z846MxT5eV8sptWADENhm4jhtoRTyd
2u4EwzP8T8Kpezgoa5lXodm3IPGA6VwQdczOcz9y/SDEcnceNYRKbpabfI0Fgy9B
AomWnOPiuic7ufk5MVimyghcjOWOK5JipBL4iVe3eH7HcSw5MNTEUSjGyf7Yn3xz
wIEJebVHDltoiQ6A7RCi+aIzGkWEHNF7v0jzMy64s3dJGpIrkZ+Qos/RSpNyOxtn
6G/Y2gwjQjDHSK6QWPLt9dYkmtKwYI8K6+/LnAaGdlfRyFiXQr4pyT9Jx7VJhbUM
Tea294NYX+PUayYVQGg9W5lRK6PxfEz1GIqVF1xBmXg+uw1kLxyEbxxKEY0v2MCr
ci4X2+LdC4Bkl7TMU9QjP31TDV5W9f8NB1KYCGPkAcvESuhBUgAPnge+AOFsL5Cb
kb8hg5K1q3LE5AZIE8qRRr9TE/Up8cjSkEPB00x1LQT7J6nB3+Ql2+FXvuxSNvi+
HXtcXEt3Tz8VRm8qjV57mQeh5CegwLkhHO/T2xLyOWPHpqtyzWREHQ8qG6A9I3pX
7EHR2LD1dF/CxnVpm2UOb03xzAMvmKixvyUhADZfeBLslhqVgGfr6wG1er5RQgGp
uvyJHHXiUZx8mg2ck1bsZra768d5OA8uVeblUDpEjZv3jOROWC+9JG0+NeNfWAgu
r15UcvFFSXOcWJK1Uo79OIB+5e7hQsOMs8GUphh42/dmW1cyyy3XmutM9LhTSTS+
VS6L5JufmYxXaTyGyopq3CRUPS454ONhSDjCgD62/JW8WBzO5E4bNGFPehn2YFaf
Y9xLt+fenOkf9vXOCUhwHGji7LelgCpr7ATCOrXIBHSusGh5b8Qv33Tn7WK0O8SG
N25hYLVT6q5kYWJ85HoEg7lYbVLsWnehLJNUQ0hhKk0wAabQScqxstMKrvFIClWL
zX/FzfbAecU9UvhvC3njIChKwe68MojTLd8vXz7zGCwLO/ReTpnfHFbhv2YDQegS
GCccRUHgw0Dv8JebfUVm1+pQTdMGViheR73Bx5fISsbmHMVaPpPdsmTrFv9a+sTw
OfxCbZLPm/afI1PcBLUy8loHdB/MsGQ4i0dV1OhqXtsUrpB9WUV2HaRQi/Nu07a/
3U20HjE4CbzwNdh8rO8L/IaajlY89hcp2Zm4mcoYhrVuhiOF/Wivb1A5qnZ3IUVJ
0mifAIFkOSwkSScrzSgZK48qhUiE50qIQehsT6i8iZbK8geyfL3RlE9c7SxPF/oW
CPPKJHmfVX+ULm/AxgzQHoNF4MeeKSuAxVIR4k9dqFaQyexWldEyXOEORkoqETBF
MMP1Cuq7dEj6zKF07UWxEYDdd3PlLB13kJRkOiKsT7C66DHsv5K8dCh3Ziaa6PSa
ydj+eAF4jr0meKA435PJ27Moq5OCvwZDLgAzUXIxKpYgBE3cc35oaYwZ3gJ5EmlO
hgpg+TimwrXD7Tqqx2WuLyXfUi3bK0h4bU7SIiRdbgoSjw56SuPe+RyPUcYsTWQK
Hm5COnDQS3v/olAj19IzOR+R6HUGPzpkP0lJY932as3Ewd58eVKxWWy7cDoSHV4b
3F/vtXQB5aM5dHit5bJyTOz/+FdKdvVwv9AFq57GEqPFiOb5Kqe4Xt0kzv8NPumG
a1GpVaMdJgUe2kjFYvNRSa4ehqsBguXWC3b+WeNitJtdRbrtNlos7AxdGAnaHMvg
UyWMAe9Pqfiz71RamOrlA7d1h1fF5R7mD2jHkB0XX1YSu58XdsGw/TfhMr0kVjTr
jUWTJkELaxcG5lOtmqkcDcI3HY4XQEpv4GnK3nDRZgIHzcPj7yrxWwlXXsbEMckf
j6WHcs7ytJLxZuzpTMaeLMuVopCO37Z+a200YfMx+Q8KAfafnuuQgOM/CAdaCWU8
xG5ynpjp0ncOyR6NIQrmumxwhlE+1YEcK8EeADGWdfjx1jKGHWa8z0a8DcfUL8eU
v/fPcwzBqq/luaVfiigcKwN123tMrewBYrXuR/2Az6cEYVr74/0wV5zWOr5MTsdi
WSO85zfJnXXegBisvosmH8ggN/mziVOhiK0O+Vz7sVMhbFqtGtdEwwborWO8O+0K
DPcn58VyCpk4dKWpTwAqcELT3d9J7jMAjupVmNbo3Tp2XAHaPdu5hTFIEXpIsR/i
LEbTmdwU6WcDjLLJFoGOD84yg6xRfecyrrEjbcFlyxsfTKQDT25QPviODvrrhRSI
gtjcmX/ieprfb8qzm2IwQe5tXxwdIhQk2Xi5e0bycA5CucgZVhZoRKh/rwPX/SOu
PklcR5QUZcE5kq3OlJ/AluqKriLNJVU4YUpnOmxTZ8JzWWWPc6rBtnfopbOiADLZ
VZzkeAWGKZEcdmXY8lvzlRVZ96GP2TvqLOT+fDPCTpL1KtwdHg6iAfOjtn7T/UmG
4Ci8EayhfPrx0xytF7ShR5yKSCja8LTgfqDW1MMZ7pL4HMqMpiwIONT/Wb/QUmOs
LpmIIL+QqN+yHwr412l6IBgNGPhDPDV8xNW/XotmuUmwosvAasKfgU7+Jw5JAbtb
PnGGDjG9wQwKqmqDrQBRdlhBIEojZeg0sVRw524FxpOaI/1zuuqIkPMATmBoChgb
qo4qX453h/pSYFbVpbenj8sFG+wn13y7dZpeFkmOmO6FJ5Vrlg/wI9p8nIyr7cT3
23i7ol/hyA6GiOZ1ANxrfVvDGiwQo62XIFRB6Cdf/lEHg78P0JEugR5PeHBkN+jA
lqA+VYfj4lQXdQc10PSD4Z8QtkgQL3IzntKjJnaDXUK2fGlszVg68PFNsLutMZn6
qDy3taVADHks62z8qSDI6UMrFfOj/eA6vU2PFMnwM75P6WNFD8aX+XV1IqFPOhsI
AYmu57omikY/cenb8mGVtYrA4PM+F88z5Yd/BArhVU6I5WCp1uxYh31Rc64p11hb
G6k1r5j/NUPLAm3owfYMlNFsdfEaUkMn77RFO7PRLLLYXm78UeXDbUJoZOjvBQNj
Wgz+sUOyw6jReaAFlzPwR8fTHvcaVrLIYFk5YCEp8eR0gbpyaR/cWhK8r4X0wDNS
yfKekxRuerawHUV0Zufz0rhOI9ibBnLI9oDmKmoErJStOHHnXftnKjB5SapcM9+R
fXW4GQ+pEhEy7JpPeeFGrKLtXytXnSi0AysrnKJb5gZE5Fp9w8CoN6SGXmrbdufj
TcDG1IvvXGjuHFEfOYYiDFeGmvrQA88WUcSRc6nU3n0PFY+8jTLpsnyJO+zEsB+f
yraV2KYFj4zqLW3XKFgD8wSzh1ChuhSiKV9qITh+hST1ovSRlCO5LrEuh2nqz3mv
Y7YjJ1GzTpeEmV25U1T7s1dSc/HGbDFB1CKHnuRsNPHTWsqAWF0e5MIO+FK0NmAy
s01/Eetrr0msTrkXBPCmx8r061uG2hN6/j46HXy8YoCHoX5pS4rJY/USDwW8YzH1
Ii9BdWMTIqkiDQV0r577Qzwa3HHn8GAIluInxE1JKHbzH8j+TKSsXuAMxKYCBqs+
6dBkbq8PNW6AbkCHRpvwDrzt0aY/aGwPrgzObg3Q7TAZfiBi2tYSEmmzhd9rDTB9
eYCeShIToWeeK6555Ed5xCrHCIBeMw2GCsp/F319tgewonKk+gl9bJ5E/BbiK12j
nPiK1/s+ujPglTEJa+QrRKHplMVbZR2qnQN/bCJis2xVrR1LrFtqKaZNDZDdwcmQ
kx5gyQfp0DTQTFQAu9aB4VNRMs7EDSfgIOyNyoi+2GLjh2E3PaJ/wg39wtY/LYfu
lb/p4we9oBrjs5OxzufI42Q1vtSoH/CUET6u5qztJ4hKedxrzH1Q2hIZIxjg0A2h
CzN85bR0VLUMSuNpsVeGN8oLvaWqwcZNivIATXUengCEiGIBUv8P/VE7DxP9xdFy
neIO4p7s2avHQ/yzzHYCjo3NXU6Ytc6mCN782PuWuWLxDHN6QQeb4K0GTqtGR5K9
2xtBA9c7Fhv591R/RJ9BTEPBsz+LFlwmqu5tvjrxSGYnqHlOYfwTZ7ZHVlbdBTPI
kuFE4TOWwQzglm50z43gvWa/q2PuI46CtAscaL+UFH2ORe3UljaiN5Ch3O02aISz
LRpQELX5lP1JioXcnUsC/7TDECsd3XN6G2JPEQYHSng0Mvang9C+b/hvkbs0PMAF
x9R3hRkMca7BPEjbr9rZJzG3k9iKwCMjIoFoKkUah78vUGaYy/m89RuUGahL2mQM
kY4v2Irt450r4C+8/erR3LOVgA3yduVvU2MyJuhm3qD1GAB/sbVcW/iXPCl1peCy
CGhKufm7pTE78mCJ7K3IZylNqqt+i2BYV7tYhIj0vHVE3dfGoItEEnpLyZG6awQz
/rj9s0o76zuyC+/bl2cHSUt6G9OIU1IUrrV7lf3Iav+qtvxCNg6QUxwkXWOGAaDR
7ReiM5hpX4ui1WuKQ+8sSmw8yt0SMqyHmPdCN4P0EtztqbOINmgtw5RLbDNuBE+c
CKJjfKiGSGuUSSh36bv4DudQJ7h3QcrDzl8fas1sKqSJbwHgDdnx5yC/0o2MkpMG
/SjjVXs/fKdeSbxdnP7fxq0WeuwUXwSj8f0HwkM2ORmpn8/ccY6I1k6cyKqUeiYc
zqA1ug2LhUWD/KeGa9GmF+rDtIeuumhBl01mudrdSJ+K9pulm+B++mWFkhpg6dZz
J2cNB5n3Ex6UPmL997lWBrmARq4mYD0XYxJ0IYdKwBKe5TFJgyE4gljm8WgRPbC3
hgHU5W9U2EZcNu8WCnu7UxaWYbwcLR0zif0nHzYLKr64XjPvxkwi+q4R1JjewQJg
s1oxYYSlt7nUY7C5x0WXDQtNDBjgw7HovN4pt/YZ8/5M74CCOJVtrSD/8XOyBMCT
gMGW9XLow3xD6cHPxfcnG1RjBAA/67w8z+bNCHqKs0Z4fk+fgbk7I84/aLr18jdi
l4y4nhcWP2JrQsbzYna9LxdeTSE/tCLV40U5Ynv+AnJAA80arGIdUGelbH2Kr3Xe
9cXCs6O7ANRPRZmXCBgTqNU3ode1gWcfjky0EU3gOO4rKnDuGY7TeDUc2Sh69TjW
nq9sgJfMqHokAt7WkIADHkhq4P9emctCje4+mSvMvqlrk5IiJK6q6S48+rzzTXLD
yCtgNpD4hXTdjQJWcPxyJ0n8hbK6zLrBk0blh9wMMKF9gzQRNyRbtNHjQrvIUkgd
FEM1dbjwbcpJKdffbaXz9OUpzXBsGiD1I7PURkDOScKrPoMs7vj+GDLeRTC6d9LH
fKUCIIJ0ASENLLSORZMGsc1voS0pFBLD1AynCVVmZG0HQzfLz1hC2A7djB524W7+
+nZ+iMVIWTHMJYNv0+Ua4y/r1wIWd4DT6wUX3ZDlibVSqAU1G8YpVCTrupBA9Waj
7zv47wEzozwr2udpi+v3uN88h/2XLkzgdAf99wMwiFV6tl5BTvVDQDHklHxgLSD1
BxYUeaBIqMls8ntIC4rxM8rduX2qAR2IhClX4+dXN9bLO5luh5Q1YL0p6HxXjT+t
zAO+Q7O9xLhLMNA7B9l5kYMvU0RphfmSQl/UoVu/0aQoDOOLGLml1GaSNu9dtivI
R6PDs6H7d64kia2Pf6otdnHGgLlqxa7dXlcYO8jU62AzycNxkH1GvnxxNVSkhXIl
pkv4TSgPUUXj9L9rNmo2TPO81TKUlNo2iOF1oG3Ff47H8w6Mw/Y6Hc0oY8SaMT2x
c1iTkzu626KZD6x43kmR4nya0PLumHQAjXO9NXQv9HwlX5j7ta0BHA34qQ/5ZnNi
8Ab1TdGX2v4Enb89karNFBTDWSwBLUXFvqC44aNFJl8IK94Ieo2NutEFYVFzEQNF
D+grq2TGb097A0P1cugeCYu93GptDsQl1GN+YqrCp+6BDi6koP7CJFE5zUGXloFX
6Kg+OjROkvoT/R7IrGa835FiVfSt/ECygmgpchiRS/DIS3qdx6ar/Lmga077eUdE
Fmu0LP/wPkaYWEJ4QWonTkBzyXq0WVrgdD1yWjWu3Sl710gA/MpEwhQWf9vNzQl6
nhHNpng5jrLHsylH/FA3V26TWVd2DYOhraPVA+0qtrdLOf96uGe5NYvgX96y1gLa
z3LkTkzBvIOfeoaO+DF0QsPa/rd67lUNw5HxOXXqxIFl5PQ7fElHzouUF4VToHJM
v0iYNDT6IWhDhoWADCJuoFDn+FkkPtM4GNdLfvoSEIrCe+x6jCpBQFabJDDsphnX
nQ4nUyVIzWMggHx8V0OmZvzLDEFud9pRnSEwURnTgf63de9ruIA656ceF/xpv9a9
z1NqQzNaO/hyE49nXeffhYH5CD6begvU5S9dPHvyQytCmz8rkEUa13DXCmlW/AOy
ioKAXwerlefse0J97lYgVpn/tkYD9HDkE58ICEyf9VSP/492LukPGD3Y6xGfczEV
dfh3vtnAsVXX0SQIy9IawvAtIBE3aA1NwEyCvhfE9y2hqlU5iFm+P1P41yi3JzkP
FWcMd71CNzB3XXEKnKekGr5994hu5r32UFWEMQAqEkmAOllACyg7PoOaxQGu0zmi
sO0CXxbdgw6f6l3nHSnTuZwqESJg2/yH82n9B6YKkgYmlwZe6GzF2E2vf/AwN9TN
cusjpH57KFiPBplrE9zmVDN5oiExcY1QRYW9XwnosXYJLWJz1ZeYn8cCcFyrthVl
zRbrau/4aab7CJnRsnIzkJROPjBanm0M9lzzhm+zK3E0yX9qBf/lKxFaTCKMAaeK
v0KBwSqvjN7fv1i0UR59nR4uYJSO0PVfT72SJxAgQT3w9XV+1leHWgogkkRozjXx
3J+0hrx3tu953Bz5FNUHPHmbokORrBd4QnU7qqVywiSb4HtCyEh/gqlGczoIQj/k
Pw0DRLUniHxhpWc0tdIJyY8POWPJZdx1hSeqrLFb0NgyOnd5rKxciLcUiSFh+6ET
RG6UIRm740KvC/vgONCM783AtvjAc7bDSYULSpig5QfFt0eYSn/i15NQlI6/BS8X
vks+tfdAA4j6ieH/K90z30O4/7YfEEcaafDsLSdZlvvJRLgYKA+GHnaa7xesibta
XxIl2QH+t1XPZk10hbomhUDyUESe0isd2x3iPdw7U2Mcy9+nJy45jbEv4GLgsWGe
OdGENg8k75Y5eAX3HlvLA+9I/GiObxiw16oYb+5xoPFsF60X3/ySd5TIWAYhvOOv
Ufo+JyiH65uUEwXpCsG5MD+8QZFP0411QpRvkDo+2FcvvfBNkUmoYOITw2U+uzFc
/Z8BoPqels+kx7OLMGZfoMjhGocwnIMnSbqa2mYGIAObtAgnvPcTTbWAxD/v67qx
PLqnmQakxEq0RPQrLWKxuU5QYFP6fwl/XyD5Hh7HA+ARQ4j1I4mMLe3sWmy1gKFZ
njwUGEgki1QdVMoPRekibIhnviOcozjxGhiu2n4fEmFDYK1yIA8+1Sh614OGCa73
/751YVVu9Ml3nglrF5QHyc5bkq5AFFyp01Tx8EPYpO2C1JltTSJGKvD0LC3a1ZoS
mfHe/A5B8H2yqUcPdtjrdKg0FcQaaHkCoKeOKXyfPKZZvoJVxOt4kmz8ag+IVUOO
ecttc+ltC4wxfAaDR6ZUa+GL9xb9L0BzIxJte0xHEifiMP/NTFXD/+wsuXAy9jFF
MCg9IqbiCB89BFU5gGDxiqAzHJijE+9+BC19sAj95CdCf8o+lDINwGrM3Xt/Oswx
ZQpeUPp44eW9gmFlK7D0zEeK0YMsbM1UgsPZ2qpeiQ5tAwlgctOu2oVLZJ6XK8dA
tTYxORe162mtgCNFLkdR3ICwqFm/DxC3DYKGGPybrUXOa2quaNm4g7L3lPf4R0Ik
DEI7GPUqGj2/VicBlTQ9wv6VEV9UWfVHz6PP4F6brPmuayvjtEx6HSvU+Kl5pD73
R0RZ6IYQSk0q96mjCK2vgXDfU+5HzwOZdPPU96QjfrHsY/2jbMWgclhCk+tSZpVx
59Y02NE6qrEOTTxdHqZOQFOUjyMcT2ITSX8csjh5yfpB1Z9qjtpaTx9VlmzW8xEZ
UoqwYxAah6pvC/8XxW/LUTrgw/WRa8gBjIjV5SIJHZOv72Q1qYjSjtKlqWyT0YZ+
WFStuOoTe5YXJ06u3WDtaFRV/bxSTB25DNLDfJXGOqbJGlu8JD0NBngUAdmIXDG6
FNFKcIMqR3NXiISkD8WHRu//zxyEYi+xLNYEdvaIrndG/XIs5mvAMmYxIZkVD1Nj
uOIvJUHWX62XVezZ2I6buVNpRmYdTSQyqcRi9OY4qYStIbx7nikxd8af3qDo+74m
c/ekLkQPz/WNhQU0yBzVxeb+m8RWqyaFSYlxA3586GcrJlKUVtFmTNx/b+BO2fzg
DDTYqKdlri6OMVxi4lbMHC95iqzxqjEpyT8f2dBjPxaW8c8D/hAS5GClGifnFQcr
xGYn9WbmSRQZBv/pxKa40ErJF6JuWnw0AYU8+nCxpHW9lmGBFNNGfyOQHqoE8szk
VI4mYTx9EvGcR3D+47LJfCgmU7eR8LDy54TsreGv7dbYs/li7TMPK7UC04SnHsxA
9Q4pqmLdVahtS3Xlw6SPEi5+EV1iIh7wa260FsDTHuMcgHfT2H38nOIPen7Vvc/W
/WTZswIyE4UB47G3hwnv+Ziv5fz07/SDmOPf7ni1BNP6wNuqsfWfpHrtZhcZ+Oxa
ZEjLdzVpUsQVAua1xTCYuVunAZ6oGyAUsQIEt0saugwi23mYe+eMyf+FQqYsfPso
R626a4OLM+Xx2z5JpeZuHsaA0X3SdASEbZVhMhtJaGZFZUEynr7uJy+Bz1+bd0Jm
LCOiSrkzYl0Oh/dbl41k3mTsPieP4XssrQBVabc2OGOnExYoSZiIAO5Czz46/Of9
iny77z2OxY9E/qp9gaGIO6RZeKOx4ji3GjjVFPb5VVYUA1MPcS4KVcsN1bBlp/oL
t9FnodpfRk1lbxgwvIJW00OGe0SIqr6TMZsIBcU40bln8t7D2L0GugzmaA+/fOf9
mA5LaAwGNO/HstaDhJcq9JdMJriuBPzTnIxs/H3/k0hk4sltuMc8gaxlbkpQ3l/l
fenzui87Z9wZLz/MtV7PVaSuBSIaOR9PFN6EDVIn651fhiXkSMoPtDWe9YTTBqdP
X3QGXmJedq1nyArZ+e+aGunn8wA/V86wtevltzz81QDe+x+4T2HcGJXPfC3Fbl+D
v/7bm8AdZKzCh5+pHk0jgqwGkVz9R61YvBMt+7DNsn6tD8n05AREZYn29p3Z24S8
8GQJeIv7f5uSnj0PabSqv1amyzyX6x/of9lM6/V8D3sh9bfEuXBuODxrApAnAEji
Ii9XYfrYvEbomX4Fo75mnL0GR6+wKZYvcnkhPWT7WCsoN8wTFiTYPHY0LyvwI01k
P+E0F/jy5WJ1i2m8ZxdchlG8icYSnJCGDEI7pogEPStZruxQT30nR1jStQd8fX9q
Wwz0OOU8wUX0N1m8/ulV9W2z8L5ZrqUQhnsGT8noguBWUiNR7/wrhZnR5sC1qffU
Bhx+pG00YUjnUsJJcdtMQBmxAGwX50VxQbHc8iwuoAtvwc5yIJM0wpPac0HxfncF
QuqF09h5HG5p645p2YtELpwtXd8RUzlubKVTYrgBl/LK1JON9b93jPdJTuV0mOZZ
hXP5RR0r7fy0mbic6GZbDMzh5L/VjmLK/iKPJf85ShIQRYXyI0fixdxs8tsDGEL8
Ay75HmT18icCHrWYEHhcvF8EK7Sh2hZzdtNpuQ0GLJ2JO/d1UrOJB6LwBQ5ast7/
0DvlX9wIqapAJW1np+nHHeXcCjHD6kV47cr5nheocD+4H6GQZA/2dpheD1Kr7voV
iLBLeZX/5YY36nnE3o/xg+ggEsEG1EQovB3R3HhJfcyKD4evziANeTo4DTy0+dRU
Je2yoUNNV+Xz/B6lIMzF9mX1Ab+5FV3dAEtswL1zDyvimTDRZGn04vsZS8fJ3/s9
d6HfPIz+mFnj32ffFvHnupn0R/Qcpxi8peoEZ+XRX1mArXXB7O3zPdEQKPbmc9gd
Nd8adY5BovvDzZ0tWD9d5eGLp+ulj//xE2LcSnwrPtj4Kc/VBIlCpblBFkQz/fVL
TrXamcQu7czliodEahFIfKys916RoJgyImpZG91cxAUCJ9zBLDIWqCbI6Y791yA3
EmXLaNBkX/7mCkoaiabJgCLjhu4SK0ezzRqy/BV/Wm490vDyrn2KmmbnNKlmcVUa
c3AM6I5mO5zUxD7oB+PjOVY5RhBPo/QKrcay4nN1vD35pQA/UYHc+MwWLuphCd0N
iafwyouINEmwNNMHQ8c5fH9wxyDLQXcSQ+eujse7Cmti7BD02Dn606QKzjv87SU+
03wHKMyWme8NpaZXOtMBJ2kighu4XLZX3dDGDRr8l+uDNJaN2z/HfTNrQi68VDF8
89h/BhWfd9dDpFXATc7OF6+o9ex2WN01IOaT1Bj4rvStLMWeWOnTazVRZvRY1omv
EhrwnK64EWyJy4Z+X7KZNNXRIGeXyYgW2rPjCe9lZrVAwYCoqJtqwmG/ePrszHLK
TTotgrAdij2GdpoDO+XFvi0kYvhq1qgaEFaPTQOcjYhesaMY7NUBZPUomrPDjMv5
cBn57OKFmk3PzrBZTGja+YqvfdzwTo9e/ivJNNVGMm0e9JF7UJ0bzV60iIRZ1/Or
GGyLIhzAwdra2CFd53bToQaNbHMmZxpDUZw2Uwn99nbPGdddDKuDFMisG9kqYWFK
dJVeWUTFqjm2UacGf+Kl90ywhIOGOG26pyhRFffyU0BNYO6E4W27Ow0DCaP7rSvU
1aYOKqnKuYmuyigHsCvkRWuWN3EBLbdJo4gCSeB84OAPCUbql0alIY+FPFpPnH1L
n84nBYltfAkvueEo6yAg3xp71/bjvxq+iC4+SztxHI5xK/mEXAEDdWKe4Akb3u9Z
eKY00tZDLGYukttFIinN8qmqKloS6QTBP74TDvDcJuBlideQbVZx/IkNgrk3X0Or
EIPK2WrEWZsrsUFyKed7H2ggYhHJ1seh8RS96ZPuKVwcQUQhGqgd/95dfq/m7kly
N9TzF10/yxl9Jhy0B9X0kGWPhuN4BlOyxWpD70QoVGL8rCXVPP/jlbF/PXzZT2hl
VFSGkk5wyZErqs8n7UtpkFMqFfs1ZkcQYbDQQqo/BK3DyM3fwekR8EtvNjfAe4Mx
FbnXSmH2omt8dp/tWiGwOupXZSA/K3cXHOw22VFm+zNR7MhCzfHD4SicVOgZXJ/u
AEnMAknW2GocUF7NfZus59qGwjXsxbjNZ7gSx2Jgcx16lTQ3jHRIlPpHPVpvTC2x
Gdz4DpeD99VZ6UDt7bwli2Xgzm5oPj88lqfLczwt2Fyg6CKKhT9kuNbmP4n5L6Ai
cmwRYb/qGdV7Ah02ydSW/ozTFCUvMVF2QOZfVginljX+x5Hghdi3URmYtEiTnDge
VHxiRUzW8RLLy2XA8neCIlMC308VbhhEbqhwgiEhfrkLD4ktOmSP8z5n9df/X1Y1
xPIAMf2aeL5ux6B+vu2Th0BwuFA+yCLDn5bxCxt5GZiRF8WvtAbwxmST0p9Cq17v
uEFD3y+yUjVd0PxI7eLddgLej5DZSjnKsNcFR75cAq4SCYWeMhr/+6jtPxk82lOB
r1EHIZGbw/s46gQi/sfRvl4vlmw37VsVDhl/EksaPJSuHzGFYaBuj8PBMQ6F1KMY
2eRUGj4ARz53uASMNuyOJ/UTKzE5CUconE/prkPx6mKfiLmogHiQpV0Ann2Oimcg
AM9qWX1dCuqkiCn9QTSrY1e9UXDAzQmtGK3Ni3X/vvYyelJsbsOOkBDUopYdH7Ea
20mN2acuvW8cGprTD5BYKflahinkasKNVNUUqKNnHJ01E4IJzz+cvv22cxs5MKs2
NCEFJEbXud04kYSEXb/pRofuFeEquvL2XwT7an77Htv876AeP3yZTcHXuvaEh7dX
YujxiJSEc0reNt+eELwtZaXrvBLVd9v8h6cQ+27I/6KtlI2MonOa1CVfx8ElUDjW
APcwNO1Umd9D3TToM8M1WCNsa7AkrssmYmRVUq/qhRRsFBJyNxMBxJjWKcCbsrb3
Hj75I5VsLKMMb9w4p2wwvLyrl5AwFpKwYHt5bqIazVZzN1rYGfxrYPwdmWevj6Ny
V3F2m9meTVAhCpe18h1dlgWgE5L7dINTLS7csjGP5SpQEDnT6Hw9HWMiOF5eT9z6
6QW5+/Wbds2WUpxz+EVI3o857v4am8OyxTlR4NNxTXqh+41omGOeIR/V5i0+uVoW
zn4fOP9XLN006Kx7zDaF8km7M5PcvM/s9+RrDB2nVgSmdew5IqR05htc6AMhrrB7
gkOILbnEHx/OgSxMv12G6+CEXQLwzg26XRdwtTsyh4WvaJAcj7GiCIO3UGAHfV/I
JN2Iij6Y09XULfEknzI+1gazSc4BVk8flBZRkWLPJS7tQd+OQp5ZdPAljLoBmZlM
K4sXQol6yms9qCsvPSTHi31UJ5q4+XgVZEpdBn0SH1so0QeVw479RaHbDyfp9zu/
nhSicQ2A/euKlqz30+Q4xgDp/7ZR29vsqHdKo2MGSFu/yglsaOh/6sE8DWWHfBJU
FhXkKTnjK0uno0G04tfYGZN/S+WOtcCPf2qV9yBdBAuNd7IMlHnJBhPFk4sr+1tK
wG86lJwtQ4RBjMrwEL+Vzp1E8g3zcq5ETEiqwd4UVTEuNyd7oU3rMN+qkJcNqPhi
AJq3FRs9RdwC9oVu6a2BFuYEII/y8Ge8hIejFysQ6L138v+6bbHNmZzikDyHM3wt
Fz4DWRm2VZhjeF7QCFqCnRhrl2ufkgtbSG9XAPWhxNwG+0ud/zoGXrHzSU5KU0JN
vfGEwHKpZp0JUBxtguWq8XU7dOJMAEhq/wzsRQrajI4XKkdpL3YRhWIx5LjcjVpT
I5oaCBj/ypBevy+xhFy0mtQBRR7LpsuSjycnYUHr4egMl+2U2KoKKLC2dNOjG/di
ZlBKpERDM3ajwhrYPY2bVTdcKntYMYh8bFJb7h2ZWecqaiYwDUVhqukYqYl71ouT
X6AUChNRllIpxckgi7iuMBD7tsj79tiXrKwgFE/Fr0OcxpRzNhxSvrrN6I2YeerW
smUajlrNDu1GXPJlbnwuN3hayIIw1r4lVmHqP45xeSdsbZbhqmyAidwg4iXT+zIT
YbD8sePZ2mc+oWxQQivMU4OYxeIgt8YaALoSZGxi59LcC74kJUTopla59jRaa5SK
bHIwCvsy+9aVEk/kI6T4vtbPV799GpsdGR29BhkZucveXg8zPGVpGDClPYLoCPo3
CnoQ9GGJTsijQoe6P14lvf93Rxg0L08jSsYko7lrjFvGeaW2Y/e4h0HFXo2tl/7o
PZXrDO+GrmHX4RkJaMByNLtbTTCoE8+lY2wPW5p6FYvrReuQ8WSQbTYyguIzZhCn
X4dm8G7sqCv4dy6qTubj0X+nU6AS/+9c3+9PcNzsZv7a9vNycgtS3gHpKDUsucwi
ZnawQN4iYUSnx8YhqD0YAIWt9xgSQQz2aWJpPnkMa271BGvaZYKIDkHHx4kZyS6D
A0NA+ucZL6/1U0sHb4Apf+fpy4JAsS25t0JwD02WaZJYxnqnImzoMqN7OEydA3Aj
bEzVM/EPIT9zh+S10gwtn7wCLjD6ffbiO/bJXQ67qVM50JZmKfXB8kUF9sxaN069
8NchLTDpVBpgpRa1QE2zTccXHpPtzn/5TnUcyIBMssXd23Ad/W/ZfeRUNTkheIpV
2IIOQCqRyVK3OaQIX2AMlvztrZ24t/uFl/iftagmYkuN4jXadsQQuMk37k3990hC
u7ypaUf4teyh/lCkqVmXI9npK05Nl0aCsRjCMChFnsCzQNhBX4Y/wrOlsUcQ8NXi
m0blXCth2KGHb0TQalAD8mXs4dSG6I+p7SkW4isSo1XttGt+is0HShE2V266chEF
VcWwe4p+R32THjgjb6x98NxEyT8CkaYNUIB64wVs4fHoFBs23lU40g9dNwkjt26x
4F3vxFMq4sdgTrpqeARhU/qKnTldsggtK75vyRltfc9sqo5xkB844nVAKJKauCQZ
2+hD8sfUEN8jLjK5Doo/lm6ypdX1C4gCEiD5a/8Vqws3T94oIbai8NTWSR2r60EM
P+wj9ji1vsm3LolcNbhSEZb8K4erXkkZUZ4r6+1UFdRADCBEZZeBaXAdWIFEYc/N
M77WEC1nor4begvhkSMhCX1byMYLq7sM3kcdhyHIMeRybLxHQIVfnIEUs8/XOPuS
gY+DK/czKYhzT8ZGaSbroLLwMPvpGdz6EKdVUYPA6zSA9/aabf9pazCQtSgV9MZT
VtpHL0tcue2QGz1T1izUtGqGEhbzvWH0rbxKJAel8QF/kKZtsZFIpNWICiaFyd+D
2Q2RcyF96ZAnLMLxg5cR2p6sQDqC6e3DbQ6KHIAahRVmdtSdZBpwIIULxzl4Rb0Q
nXc5FLvJmtgNqGTs2Ki5XNr3S1ZW3Z9Rr9b4BDi8AP5W16mZ6LmXw5fHswqSpwKv
o0p/I/VNAVVOGPF68eQLFBsTPVugwKD2MMPE4LWgCRVMBvV+tXOGbgKtTMnvDIAs
d/1VPPThSpSGl+PnHsng3PA7xLze5ggw5xEsxSVQxyNuvFoeb7bfypEWo5YAzy+T
uxTDus0OgzLGDLvEjDXuU8GUuh3ZqhdSHXAmy50B/YtOtXPkSTCZAq6GeME74zwW
NCtQi+AiTN3AXHxHf/4el8E2CmrJY/KZ5+32J76CVQxUwgsu7Yr3zFoHzlTthdpx
88rfEW0quOsdInqnKJn7w2fNfD5wL29EJxpHUUQQXqSj5WB/zygzd+I3QczHc6lp
uLb59iA0OkKgzqQYQEQ5AxoC8i96RZh2bOjEo5F3IlIu+J9Ui3AsBapmE5erTF8k
RRxaujSOzelo5lFvyZ0JeegAsRTmzDfw3dhj2jT2TpsKBb388SbLhYz/sQhbd5VV
PHPCZkq5hCBtPVxL1AuKydMcAQinLLSpS84fVybUL5MoKz0bmXKib7eh+vNLVcbL
o3nvzxrnoQmLmk2mNMc7Qf2Db3zSyrhMdsKvn5TKF8vXCP+LgmSBOkQmByAOW1Vh
pXfZO58S+aI+RHRtqCWkrrpJL0n4ZweIu3joUna32N63bBscYUXZ2rph+IHQ6H3z
q7iXFfdki79o8YE/GpE0rrUIy+8h5jUAHwP7p8GDgxgi/aEN09RrZJ979rWT3fEm
tQbLWnbTCrNZ8OurK36/VSf21yZXX2ESpuWNf7OTe8S1MyfM4fN3yip3+uZewECD
RdVhZJJjlfsYn/pbfesipXJ1e1HQpOl/h1tcmomHgrr9tsasSmjOvd3jMrNT81OH
R0g75XFeVPg+X+tUxyhRYP5bvi50WqiSoyrvCmI2pl5Vcfhk7+cNVnDkcaRsyYNa
IabaymcW9FTabLWH1vmSnJ6ggT49kFSRp+y58Ed2XKBcZ/cD/Y/HW6LYkE5pyTsI
eQYNr+g8XxdupCZ+FQLRVkg/mNyM8bWy43PnlfGh2l+1UrIvdxYPraAml/JF6uUB
viU+tOjNB4yV6I/vwfwvLUOIQnnIm24oahKaSgMySRUwKEppL1m30ddb5cUro8GF
mPHdOqyeuAkMX8vaTlspIAN3nMFQmMoUSL3lwF1F67+VYaazmTvHe6oPYq84ij6q
Hu7cYPObSp9ftyZZz8riOTXVOW/2OlcznkYy/W08alG4Gz3wpZptJBvzHuaB5FcI
mjpTAN3Y4452w2lLfwJ93yL6HNNbPhKxZJMMPJw39IsIBy63UzNFuACK811U8MXi
JPMh/AFoMCeqpV788lHfqYoEu8KYFHoAUfxwmawBNVGiCfvkUEjR+ORsHpA7qWTN
FeHbL/tw1oK6MaP2Ld8eR6VgGkKVTiE0mNgPYWhgK+lxlLArnxuxIBVj2X1LHZOO
ZqJ8TOcXK5g1e2gGsjJm8q0YE0N3tlZy0Lg9J8K86UFX0AXf4nl8Po/WQ/b+Yszl
zddN/zAsJQlJe9J0fHnpbkSHTD4YYGO84KzuuD7lz6wfU223Zgw/3P9lzSAyenDb
enoS4k5dM5aOpB0WFlwEql7PBRWbLeZgLugzWEtq9bih7WNNDFq1KX6hzA6PVZ0T
Ct4sEHJIcE7uJep55AhOI+rvojXxkrWdHhbAGHVYa5tSitdTkDBu3ZpPnfiLtymj
4yd8swcnTUhPSyL8GWKAVGHTa4FJWO3/dz15X9wjd0e+kQrq8YiqpDLgpPfjELBN
vm1mgA3KuzPG5ujOBJp5RA+7Cg8pWPcbwuFCN44fYxSqkwLMV9Ex+FCDoRv9wkyv
bJmyKJxjN3RzPnhlIku4CR/fUcUl8yNoNy4XJs0xLh+rOq3OkbjITQlMpBwAYKqc
JBLWA1Eeqd4cSqwchwkoJ0+1yXzZPAOCupNrfyhzJ0IGlP93t12bXKS8NgHtFeql
VuhgOSomURpskurzyf72zRsazWSYkJjD73UECxHKo8g8GSgS9IPtgNEpaaSo/9tG
Dmq/MMdCRBHtd4gBLpRdjKEbjuxfKl6bLXEDMWHjwX3zCXw/IEGxvVwx9d6gmtda
goAg9bh6kPtjdyWOJD42g6hxJfbPwqa0KlgjSTkXoO4S0me2+mk+Ac81sdX++p4E
GDTvMi/Szfw54lCJieqL3LoCtXyZX4rWjc9LWJLIRRVUUwEBBhNE0X+8OYId+5hc
tHNrBRq0vDSsobtNu/BfZ4SasGoyWCsQ9X//xhAyUd67m0JjwarTIo1h9VenZ9bj
/S4fzL3TykUonxv1hiAVV+fSp9DYGnRNdI/CiwVw9pMy9oxk+Bm1k5YoriJPGWbk
FwXSN4dHlzPE69rUvFAGBDHXIjLdyClIbmOgatBf1jVLQt5SGfTd3FjkXEkjQ4fv
5zVQM8vw1CE8nYCeBPv2eU36XDcTM/x9bJQhAzregtxT5cyBHvbMt1yyNpMyB8Jq
ruUbig3/uN1CU0M37mxK3KH/eEVPPvceNtcu4ot6OsAlLbFoxtM/U02kpZShbfw4
i5bVNGZV3YuQt5YyAiXPsu+doM0y3d9q/SRdxjAjonnpaeJtBvNxpWPaolfP3QL2
C/Qt7+j78KqYe+DwTO2eUTPMUBBDmV0LZi9tGv5RSVtaRxNXoyeqvf3Soy4R4MSy
N1LSpTPs+BeSZZCerUxaAGO9YsRRtNoehr0mK4/yOl9YiDbpHnkYnKr/8cLNtIm3
3sd7sz7feE7l7lGypHVvH6mrFl2EKh3oduh+e8YGibaWmpPO/cELbHRKumpZmMSB
rtWlHDgD5moc2ph+1mZc6pypVHWC1MtvmnIuECVWV1PNShmFji8FaXSAsITSq+A9
Zj81rGIGj5Pmljr1WGbURa2w9nPM8oUP2UgsFWTxlWZ2vmrdAXr+Vx0gK2U+qbNO
BYacttkZI3eF+kJf/1TbbG2PSKo9UngfZP6/yTHNPuZUEQTGqqSH+HmKnJWso5Bo
ZDMrd4fK00HvrHm90Htw0zYkfs5bCRZAl4qnYv0LzUYzWZOZsTVR/OVl0i7qcDgF
U3gzTzV3l48E+bkzzoKqTTBzPcKMGYJQYXcGFSRe4sgurXuLe0P0zm/RPpoG7PWY
/DLXdZLuj/VZUvzHGERb3oFmSEy4oufKvclfAH20gRCCX/ni1IAWEG9NzLwPH4Kf
bY0bIm/XM5vrL0nL908QUzlfLBavNsuFTv/6DL0HEP6IxaxfmALoa2o8lSETvBLM
AuBIFZsf6DxvtTyAP2nrsKWNocasvJD71LWLnKoqs0hjRHrHL8pc3TdprM0HG8KV
2+62x5bDQfIqlBp8L4GTzwzvTGP6hOjOGZQ0koX8tZ0mIMEHv19OGBmPRcx9n+KA
qJjsGu3NDqLxXQ5lL9m9cqgsrCbT9d5f4TM1by3iTOMo5Opqpr0HlrdjyngUAq/S
E2eFFWHjarIRIA/N5gdoZb6xSCAVkO7fHdF9N+GcmjZu5bPaSJdb6iHcJWBXSDBY
IuLWYiyE4gBQ6Rf7IfxPfYnKkSlnuQQtRRI4OP17Obq38Rt6EbOzlGIIIjnxurTH
vBb+QQjueQKk6I0zOdvzr+soCCd192ngLPVRn9k8ExyNxywpxM86s3ERsiskkn/Z
LJCh7Iy2kBEKi3rXz8UnXwswNPTKhFGsg5CdK2/epZheDoAn2ZpvuQQmt5LNCQct
rIOPNi4zVUZPIhBlqHICdrW9e7aG0WDcTthdl+gg0S8NZ+hyYDGCf+Zs8y+l3jjf
84tUTpOqWcRoa+C++MrR9ND0mcvdD4Uq4Ae/tDRg6RTN1tQ3dFM3uC1TAOEAAyRg
tNCvISNtheP6NcPPTs20SI8msKVmkUNwJDkBwXe+scimspP7OqLGl5RLbgqCfMf4
ErlH1O8AJn9KR4Ou7+LJUkH2pxdhnCnNp68Jj1HIP08yVUbDUCMB8/sCCxzi7Shq
9JxGxko/V7D/QLx3CIonarbhruRVBFZJOWktG+ZG7owmSyadEdunRzKyAKGnmssw
h7W1fvOVeZf6URgWtdo172p4hgvoETs0QfcxjpsOO51dQkjVgRJtSWx11fBjdZbI
Yn4agUS8GMHkV/i7Cmb7vgi3187RDB/BrZyARESZYJDf2Upm7hj5CIo2dYE4ViWY
1dm0+kFsf69gIYiOU5p3gxbz29IghFk6u+b4xbSYacSSxqm5olQsIrTn4yA6AQfG
f9AUV95XTfAHuvbIj1ZvE2yyFuBAjWJxPLijU70YTJIwei50DitlODf2227p478X
vfjbG2LbdIbMeETESliqAXJMWLSgz1B2gkI067UVpeUoEPRYBCsj+S+Sze8t0038
kkbzis/Ee2jkbsY1G7NJZnruB3v9ewZ5rAiqvVsnmVCGvsBrHerVfUENtLsd6zfy
NYe/68/EomcIHdq3W40T4qxCy6IabWSE8z2sJUDUdII0U82U4vTHm00DKSYOQTEV
JHv+xVEynAwmrk/Gt2iI40XxbbDMMrqA6vc96Jm3cKBegZBE3kjtC/QfwXCw4HXj
yLPyuq7HZ33/FQFrS/wUvG6YEVx2C6mW8pMyfi7v3ZjbsgkptyfhCKorcvI9TbKa
uLF4bbhbPD2PNfGQbMPF1h2EIs/W00yCCRogzZ/+GPERQ5d8yfxJojJSic062KLU
DuKgqu780ZHWP2t7+NkxTxlXNFFDbKXAv4QuKVXaOQGp3xpJETp5f83oIN+XptjH
Yt0OjAU6bkZXGB1dnu60lvtBkDDvFq4jM/bgFRG3O156sCdoeTTQcOQl2ldGLN2Y
2dbJUt9kAsAufwr7tfWHIB9Rqlygb06MXXHDB7kux+urSO4bChS3Qk6txH80C9rK
HSpeA7bMh/Ij1e8qt4XrPrGmD7ylLT9MDrVXvcAT1FxwSy4w/KFNTrX8k4UcMsSQ
ExTz6osrR5JsfzXDW7FSi312EhAlmLgGhjiF1+ZutrQ7OlTsZryhz39DKyBGmQ4/
FsAglwhahLS/fvrhFXUN9lBQqLES4zgGrwN/ZmFDvn9xWKhL843p+DK76Qa5JP0g
qXU/Wc1L/I16SHhgdz70eFJlA2I3GUFnUWc5JX8omYO/LPmFU5WsIV6cPOIkUlZ6
WvSSA/UtwkWSPPUOWoSuz94DefC+v8Y7N//evMJPDh11aNXQLWIudNX8nbwGY9vu
fM59hcFODPk5Cm8HrfxQXVAgpxPGAtOjjbtjqR1sYZ5DOWLbuYrfTyAKdduNxJJ0
+peecP2Ku1hkHDL0sSyVSuli7LZ0hqtTJYskNWh0YHUFk6uVhfWZiLAvQxEB+8ka
0O8ZmVAlkc605yQ01Sw4kXkVCTyPV3UtQMYXGT4v2+CN0mIao9xKmfCq/guYs6Ws
qCwzF7qyCO1RQwpusjxUwzFy0NL1UTdd1jl8WTwXs3j64CbajWzNay6QHTzMBDtI
AmhV8YAKnK9Izf7Y3Gat4BHuBxyATLwuyT5cHrYaRT/KEx87EPj2NOFfA+y9UDO7
J/Sx8NBuUgqJkofbdXGfVuBGNHp0dpb+cED3FCm6+mTTAaPBfrNgK0FD0kc//Hs+
26Z6K84qpFk3GjJpbofdlraE7+IlMKV/SGlMdTGtEJdGaDAG/dt3nC5/C3QicJAQ
KU6DHM7tmj6hOMK5d2aZTAksOkq0INUdBa8KyWoW7dVJYtocBwNeRrmfCmx51yqj
fFbk1sc5p5Vn+6HoHXb+K78z02nzvUS4IJKHbbmrz1IpeyXQ8ik+ITxM5TMFwgQH
DxcX8VIDqpSjCk0M+zjGU4xcCp40ybF+6KNy4sebjL8T51NFbdPvul1e6kzSklhW
kCerjWaf8yF8JS4SVRFW8NOvDC/8lHuwCz4qRKDmAxyCr7h9ElWTXXn1NxxruCcD
AhVLNex6KH03CrazxDEsyDpIxc/9U+ayXdc5Qrc6Xy6z8vZTTD+S4ph146M6XHhF
YPUDhtpx3n0bgllDtyr/f8dm6ddaSsmtSNmeO+1uOCQ60XISPfx3HOfahj0UYemL
nn2kE13vP79tjraYKoIwU3J3CUX+zDiBfWSfY6e4jkTPxq+y8QHrWrREhvPJY0sz
zcNgsG56bdtIoiIHGZH+RHyS/I88IftmQdL0rXW8nelgWymKmA+9U2WU7xJ+gWkV
RgDhLOqcvFhhMtzjeERX7NFjOK5YyNxWjovK89f0J/pAmJR6Bk3q7rrs2n1NMRVX
F5G9QQiunR44ihl845cxYyzI41t4sfaMLJj9WXtPy3a0vrLn6S8hqRqZDGujWrBR
uKBq/snq0neFTpe+iK4pgN5zsYs3srBkg5b8+j2rOSNTtDl5qaUqAbg4IjLiem2e
n6KophkLsJEizo6vNy7B9tl86il67lfWlQzlNfE3HDx/RfteD64Takhjli/SJ+DM
Xz73Wq483UxhN0J1x39DMLhsuYO6nr7iZHP0TGlZuYKRCeD9/jo2z46qfBNicfPA
fu5DdGYXLGToDUW7bZoprW6npi1S2svhW6m6w810GuRhwW94oOmCESyMiZb+w3MH
FIfz1eqySOP7IHceyNrCQvlpcz5K7oTOucy+J3uhMOtc5gzbsuCctXtFE2jP2lxS
l/pJ36+VHCHpmrmNXKYeMLYVSsSYTIZRIGMCR3sYVecn/TRY/afX4Z0+64vEvGw3
6v8XViVO+qw02PLMITEtMc8POz7YQ4pLhp7L7bF2+7fy47v85WNONqIUAX2U+EJQ
SEliu1KoIDFd0BPIYxXMxAnUMEYpGe3qej+h/9krVikWcsebkaUirkKo/VSQisKX
hRSkiwMu623bf1PKFMDfc4YpTBM+gUdVDlrarKKD3/Di0JE1EcHb+4Pd8OSCL9WQ
tw93+QFzbrtujEnhYrUW6wWlAAh2FUeYgpwlLNJT9wOTH31MI1k7/Nxk4c/dGoRI
qWJ+RiqDN+Le4Oeq6B5hTXzW800c6/Ywo8k/n0cteLU5K6loMfMwKeeKXC8oB7J9
psjRQn0AejomDtsbx9w0J9in9hLFn3DpZNPP4aoDfGTg0Ur8yVzgLLIObMW/lRJ2
CDmCAMAfv7qEsINDzozumg9VSDb1bqFQS1n07wjWGNr/IsZmH4isvlfrqey5J/L/
qkCO8KzgshSyPkobDLgYjdUdYzrVvv67FHUGOjsbD7+HuSY/eKzvZrLWLcSlQHhE
CMA74kQkb/6EGkGRaZ6BkEojEnrM9y1QjlhPltul1yVZt7H9qn1/Y5Jw/3Qi84qV
rZDYo8FKCGXgdkUeLTKroqi4XcKSh33gLTCw02lQfDD0N48KwbHKpJro/NP8gmhD
wsGov7wVhEuVk34rec0pf4E3hYIXKRpg+5EeuW+VcYCzMPZQwWux1A65yqDqO+ND
g904gwjiUMl4p/IjAuNntoZ/b3Fz0/pQ3cnfL8jZj38BfStVT8Vz6kijnrNlJJwT
tDk5GD0uS3LSAkVi3o+i4Zu5mi0a0Xz/4JGbkCMAhxLN/7pQe7ccpDEay9zczD/5
V1ygrobgF1Ot0E30et39UuqBxUozJMIlIOGGdArDjPIhJisQ82wHNekjJ9/DQms3
Ii6Z6kOgX3yfwQ3L91sBd4hvEP6kQRYcrTXopJzs6CglcAxu06e64S1SUgsTBh4v
ih5MWzxxTaFREWC1e+Z781FmtJVa1ZyqXxy5zgB6zCT3JikaxRO0c7MWW/pHNFUT
WnTqP+P4hnvJ8MSRkYClJXNKVpbQoqcLRLrZ6y7/Bd5iqCumB0RT+3VcABBppsYq
KrNrol8HB/CUv+M6jgEAsjtprzcksY96JQrt5zCfpNbolvAgH2I1plNJqNvLuiBZ
Sua/H8IzMwEUGgXfQlZkBAvf3iX17a2Fputhh8lCn9SPHEtC1N57n/uurZS2vmF+
LykJYahP0AFTtGE2AfXNDjZ0KztKdkFO0u/1vvKskaKycW0WANfAihsz88xL2Lf4
UAqqegwG4APkHBM+mcsqy4Gl1FVHMdxU0HT97wj29CfAWTJ3/TOlSOB4DoC/vv0d
kZDwo/IWUZYi+hzKdGPy5dOwp4hXo3GIoi/IJPHfVJF8h56AxJ4qWNWwZLNhnYyG
V45Vjup/yX9Loj9WSs5PmZ0baKsv5I8uYFo38eDst0GfFtnDUMHpMGfOvm2JboT3
9DVDmY5lGbnsHNZCDkXofk9S4j9WFDRn0rwqqoTOSAOje5kbudGw6ETX/zizeXWl
2IX0TuisU6lYoVpnyyRoeu2YXIsRyc2qOSJZeAUMVrBYib40s+LYm5VQqoiq/3W0
l7xhB9m1LY78kU2Vd7mqnmTOC1UOYyDUKaGcBEk/3CYNWdIwOavZ3TF64HPAMF4u
9XnDeHZ/V2dOO4d5Ize7g2teH8WVGrsOGVxdUwGafk2ibMvDe1530TM+U3bYjCBD
AP6iJztc+xd77MsPBKFXptXHwZNGqB0aHzYPVazOx8GIVskTo9irw9kFxiztT8fd
b0jvPO42jTPnXXpry6peJH05CFZuCpg7udnyyOU4BByHXfF5ZAM+clIRQVizW7G1
Ull+tvZIQ2bJEEt2KxIrz1rzej/xhZLgqeflJD9bJZ6JDXiyFR7o28/VQk4yraHb
XztoFlrX6oTdP3xBTOP93W//Avln0TRpaD6OEk+mCLV36rEUd7IZFWVBnYdIPeoO
pu+TtXcaiDQOAl6pQDiXw7l6JqG4XRnIAU5tPZia+0mMsqP/21N+iryHOOT+Cg4G
NBZHs2HFP4MjucqXQSiOat66AADQPjLvrgDyzMwDkBe0Ibzpozg1Tv0bcQg9xgTm
2t1q2c86SsCYxT/LeebqXsjQIlZQD+3JpCfZ6WP26tyW+QhMVyDmPvEjnv88up0J
r+eVIihFjcLthXVsO0ZlPm7gXJdcz6TnQGotNtwbzGPR1RlOzElCdtpt6JGMuyX0
wYJ0JiZXuf+PXUC9mc/iKysYUIx2oVTEQJLQQlwvsClr7IwAh+vBLxHl2PyJaOjC
KCtGQ6uXLeWmcGs5UiV0X98rAMzuy3HKHnn+DvmaZ+9NZLSy4NqdhHsBYOC2eaod
/Mjb+XZAO1Dc2UsWd84h+umaaNf6kmK8+nvC3SFLi6lt53ucg9uva0F1W8qklznt
GFCi9SocDSmtk4q6MImsS1WojIitQ/4y7JdZ+9oLbFHwAaHiPmYmsY/kf6Qvdqpi
J80xLU/mUCDf9uRfFkKeXooWxxb2t/IUt1g2I2Qb1+jhdMivy3Z0JktGIvfVP8+p
3P5WEm2EdAo9r0thFqrvinpp2S+R7ul9DCYgg1+gmOVvgPZEaTAyCF1ZxoDAnpd5
aqJ4DWxNo91FSSw/6HUf5/hnr0MnTaZI7ttzhNtgTiX0/JmJDYtwwB2ZcFDyFYJU
URhYXt09DXgBeFT6wHIdjeH5NG4NN2VQROZnrn/EUcMnyRnZq7F47z/ZtuJUsqlm
dbDW0vnU/xvAV0j2UL56dDxASWpUr1DNSQesieRmU4HTDu/CMp6q1biTiCKiA/d9
QfIyEhYMFyu1Va6b8MSIHK2C4kCF53oOCg3MamV7w5VcAJody8drf6cfR6OxFyxT
khGHwESq+f5/bd2ub/Tdi1QeHDa7TNQqVSzSEBx2rmnANkWUGrTAWnNe0VHnQTSF
kQuhrzgX3u2LHY0pLNbiJXNA+EUTV6DczT195Jk9/FgzcpxyrCW9Ay5+PtGh/xuO
M8zEBeyjp4ppAkUZxCX69F0zqk7iAWV4A8/PeLg2+rGJzlb7osHhUalKCGQcqPUn
OvBzzKcFN+Vc3OER8KoCbU2h2hfjk18WDNI+Q5hD0uTrad9NoBsYWIY/FsSwbju2
H98fmP/TMQRs3ARgWSNjmUgY7PBVaE2eyfhEyah+j2dScAJ1GY089e9PMCXkmFot
2XzIeTc+Iz0iquxyViHxBYImNUDHG33THcMRBk2y7eJxl2xzdIegKS2SZPYdFAnM
lEgtPwtPbDHKAT0FxgIFiBef8nNouVm5rGNZ1tVrvYs/8rb/QiP+BUWfuip5bipQ
bTVAggkUyCJQRJTYHz1jEl2Do0y2Pc1LtaUWCFD1pJRYZD4LUv4xTgog08yRRKYR
ApCCpoI7o0wVOzv73gAdDl5yIxPKRbfg50C84VbC7o9qVu52WzvJQsn2QwURh1M7
jeIf1YV0ZNOoiwJnL2zFxeL9Nf7Mw97KSK8eTrctBgQuH+dne7hFNNcjdYv2s+z/
VQPxxfx2iRfGKGE/c2zHLQ+W75b6x98AxLr5LNXRiQabYlyYsLh0AaFma02Xidxy
7sUdLMseq7jkbBuf95T7KZqy/LFhelrdT3YvAIrIGMLov6tG15Ce8eF1savhru+3
IdmgedKHxYQRZhpV/W1pBZ9o86TPi3oAl/tADRieVtirBKTOOTC6NifM0gKft/hh
HJQhph8ppFswGjZxqdRhRGRWhNSBaZn49oUASdfGfW4DSpb9M/fpHh7ccLm4hd14
Fv8RuqZdStbH6bQBqEdnwVzWzld3X8Q7W5lZzQzN4mi8Ae9M52BopfuWrwm8Fbxh
8hT+sskPXDlS8Buc+WZoD6DjYYXuOpABLbUnWEWbnSD/NXKM9akEQWrP179RZMV7
jrmuqMhNUYJipaO0vq4gybcUOziqRLpHPO3Ka/MLob1DJQbzZx6Fs2xWgd/J3BBw
ptCMyyjEJxVLmTfZM/Qf6fLPqK0rJS+0WrpmT3p5LK4gV1AUqYIr5/1cM6iyYInn
g2d4CIGogIy+FAZGmCNUOzuIO7f8zoGB+TUtuGSSId49Q8F/m0JuzIXXlI/PSvyr
i4vVPeFOjvHhWCcuKz777GNCSgP4F7zs1ELNKY5giMrqRINBruTrnKEnwsZ0rcye
XPbn+99W2gcO7yXOsDg69n0LzmVFfCFnqsHW0zwhMqwcP85ujCPjPfkDHohFcBZg
00WR4THfMpVquUsFs19HjB060XEnqF7jJFY4sKNRpmWnLurKB0pfNAYP8RGKBknC
Qsm5WBBvE05XbHDV9wDsWMj3iVjgTZKPj91AwDsY0kqXMBMM4l/DckTIeFQHOmyA
bj34x6TcAWZysjxnFI5ePBP/sI5/+IMHZVdnMgh2H9jVWmJoE0QlUIFGNdK94yr3
XO9vVqxzG7xOnyglw3w+zuwzkDxytGVQTk2Ms6Tp0J2HehvT4VioEz95jXUDu43F
MafMMGlRCp63Ia3W71Uiz7nsDS6SPAjAjimrEcxGwte29xnCW2/B1Cvkh6VgxQG7
il4nz858pWC7BG730oWAv1z+IBZtM+GcWWrfGVmKZTXs5Mx6CU8lvzfzIItf4UMD
ysi5uQ3DVCzJ3Ep7zwt4fK2tP9ol7UU9Wwa2ghrr50Js7JLoNesYYkJFFlLd4+h8
FRhuR+rJww+hk5E/KofagMN6PiCGAzeDNBsghS1l/uBPhGBHjCuuwxnS9JpEQkGW
NxiomO99z0SRugLZuZEe3a/hyzLASN3hi1no++8jkk7KKsg4s/2gXAuWs0EMBPjs
vOdtmghHqfNYTp/lvkWOQVrEbmPbgp1NXq+XLeHYIGXkAwqTon72IK6EobICDpgu
aBm7KANATXPOnkPhhMIbGHduNu/METhBoMQog0GSqMW7F9/SQL7MupXe2wSJImh9
Awrv9htf9VxxjXoNaAkzrA6flZfxTgQNlTbdB1z4KFfTo11XnDH3wdY3uJR8bQiR
wUkG0MxNtGT+gK4t2MSpDaOOc5j1DBNJn0Nq1HPTfeZsDn5AxjowM+r8ZhN1dmJT
nwW2663pPtRzT8KhMjRcMXg8qmwYPemzggugSGj5U2rD3yFQUwnSwnUnWP+27681
Jp2Ed1E7Vy1QiFk+EH12pwFB9IAjXxbMlTerAEn5i4ZZ40RRdo+dpj6ssgf6eqEE
iuJRdO9Afw1tW59hJw4M5NoVkBPicw6c2MmV8dSQq53NGMsvshR/XvCSFcs+JO3U
qtbBLL8SrTMVSPo5Vkvz5q/thG9I2WJHftcO6ab4aFM=
`protect END_PROTECTED
