`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveArJCP/mMRT2m3MgXDWuktsj2U8XFxeNxfYktJUg+Ua6
3UzuQPgGnrGB1ytvPZ0E4PmDum2Y8ysKZpELCRDn619H7Sn2lwsAjKkeggJrp4HY
fPxdDcnoVWQJCypucL1D8peH6x3nd8b6vr+2NiHSP7bDaxD9qUceVet5HZYBOs38
lJCqRVMcNur1ZR93waTwMR+J6MKKhOgtge5C+RG0aq+wRV5ZVIHzbi4TIkAdiMNy
GwJJlr4qQ64lTRK8G5bvtg==
`protect END_PROTECTED
