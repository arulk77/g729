`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGdr1vNoZkj4Fa4T4fmn91IZBtHNcqnGh69koXabyBZC
1yo3CNRerx1bUrH4PLhhhH01XkRWGXwo8tCQvcNYQKGJvh26wiLaNzdk5Sy6QgEJ
ZN1HynZzB2uPfQuPiZd6fvHwLKUtYUn8Er+R8o7qDB2KFHEV3UYCCWghYNz7CCpo
kU4B2C+gt7B0yDUpnROhEDS4Joq8ogYQLEXs0VO9cdomwjHR+y2rmIcgQdCDGpc3
+SiV8aWCvYZXu/b9B3+aTvsYqKdeD94NuKHFDv3+jitqaTAUZKt12nP+LmxzlqGN
vzWScejGMQ7k2Lvbx6FD4vJKBaHsTr+sHqu69ET6eUTm5bu1EYT7xLkYRl/TWBHe
`protect END_PROTECTED
