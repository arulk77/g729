`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
7RWERbz/SCu29vx1yp3KRLRiDqAZ+Uy61uejUTqWG4aODnKkaDoSTMzSULbvbL4u
dUOPWzUmTygDVC9zcIIEtAin/Lmu0buj5qDJYa/pq5oUWP5nHzbSoeVE+w6ZoXno
KHcgb8VuDJ1bQ/dv0MS2sS3lqCe2jCwhxVBCJyL1eEPPWbef/H2Bi4Mh7K6a6yjl
`protect END_PROTECTED
