`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41wIHjkLqhkVGO8gFwJSmfHGZ/fxRztbbDB6EenWonFP
UAzuHrb+6ou05q18pSwdhmnUHoDt6iICuZA13Ecq5Wk06OUQfYXjw5BfGHZpYQEN
cqLa7jcpL0iPv1STTE56ryxmBASXbS/84kPMZ0LXic9ntPvE8TNsDdozJiuPzWpF
7qxxwdr2pN+1UfTiV/T94/dTJJbmrlOIGHP3eIJBzBOlqQwaDoI+2o4JD14txnS/
tJqq86l7/yMeKe4k3xWTyuB3o2pz0nMFqMwtl2/1qhSbK/Frvoq8s8oUW/arc5EA
FviDCBviUYmGRNGr0nBk6g==
`protect END_PROTECTED
