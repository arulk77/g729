`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCdeoX4XX2N4PPs70W/Mtn0er0QripY1xmuRhIxaYfyR
o43N+OtuwVBBrWfBXfGo9OOEYE76TarRmXZNH8FJafrJmUidH98/gsP2ieNbdU3d
3zoarOIFobUGK/tnEL7GcRTXnAT+2WpQCGkDuKji9OsMzkRSr0nWWJKcy4l0k3Ls
zbOoLp9J/G5+SBu86dFNRZ9kcN77i+ffCzB5/7hHszWbYlJCFuZ72yGi/xqSZC6M
VmXo7FE837UPhjymU6N5DthZnNoeqrwdiua7zecPhiaFGixYmdg0Yy394joxBu4X
JETrHQTFpgbw5ZEnhZeIhhT6olKTRQIdxbuD5uDeYLTJeZfmVRtCuql/flK8rI5V
F1JR2EjeFTy0ibt2FnHQHMIAIhkyskbczqDowU43CBUvnUEM3705U1g1LZjt66Uc
XW3lzVO/T6Xb+5wBkz9BHgXnAa+BnPbf7f16OiJ4Rqr5kv8ZF6zmCKEVmaicSMrf
D8WdmgH69WDHGFGkemOAdAbTFWdd01MVa5YbbtA4dMHVnEazSe+thehh+7CbAzH8
`protect END_PROTECTED
