`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJlyjLqHwcjDT2GJ60UdMzRGeXWVIyrf2VjGfliTvSb2
YBumKV0LcnPpk0MZSvNHkMkH6wtOu8uyeDQ1zaHvydMMtfQzkkNPcKE4te8aMAPR
jxEXN4TC9LBPDlBFwC7VJLqynt3XysY2Rf0TWqyisqArRN3BVcEj0wR5qrJgEw7r
yFt0vSFI4qB6ji4XkNyRwKUXCEin2Imd3tjmHUuGwuI0PfV83XhJA1ctKHsx2l/l
bZj/0yFf0JKAccg7O3aZ1RowV70xlegak8CJVdO30slLFexz9aHLqDmzX0AEdyae
`protect END_PROTECTED
