`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCWsCTtdeCRNZ/mI3bZdD/QzxLirDX5zZjsTXe1HZPfj
c5ExQiK12CX+1yivfyuW0fisqK3het8gcmoKDRuATpDzmIkMtJSzAXWuZUFmGhqg
4SHYPqyxuBUMPr2CPwHV9dQXxIbOIr2ELG7V4Y+RQH/VRLBVbq918L++zTgxBHJY
ryxr73NRoBbc+u+RC/I0TcZQppXRGj5qX5CKEpsXsmESPAAHjS59+bhWyi9v1sjX
YSh1jEpL54PvPWooBLyDCTaBmYvsok8gCvzOba+ECWfxvfDlU8stXy2plvNI7Y62
H0zzzstW+3OeJ0CLzrfLyejfrm0LbnTGXwt4QiGv/li23yZkJAGwlPMqLhScsrcL
nqVzbHN7H22wydNxI7LVmhJ4kooM2Oe5f/81dJxwhvMQNh5einsCG6CkLAwIvJIe
lHxuu5qHyY62bsKUZho1KyYZgilMgHgwle7l7Ic3q2PEMdkpVFp7OAsZR3fJkHrm
79lpZBgZU1WAF6fYvLvfTYstfexkEUjvk/m/6z23iM53I7Wf7I6uLimno2biGpmP
HeKXMrSD/e7YxJYCqWq+2pRJIk6LqNsI5SenKPMMSoYW+XMl6lLHdtx9C6qRMbKf
xPJSNgAALHzT1mKO4HUDRUfR2TRsqH8irjadTIDflebaOaOU1zYl52UqP0YnEhhC
cI+bRgCloYo8ZTG+WhisETC4ZDTeVGwwLrNCKMA0Vov1S6CCtRQ4Nc6UoOfMbQGD
PTUc8bs3iMMoCnaj66pAre/36L1tqdYgWM3tQ45vnBkbsu3tPy2I/0VDvbbz6iiQ
`protect END_PROTECTED
