`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL2toM7dPgYsTlgY2tRu0ytdbtp4NLl7AS2oyFXuAEHz
Flff4is4a/pSWDSMUqptrJVuT/2LX+f8WDW6gxtsD/HXKOPi6MD74RX7AntLAADQ
vVQpQQlvgY6qRRDQLuXLaOeHgcwMhMgF9no7mUk70rb2CZC5IJGHCqtp3HbRSIwP
yh0ICDfVfgqUVYc6rwrLx0oFFx1dG6T8Nq44RfraLUyUOkK09GBWnubUfp5yrcL5
mHUTkcaQclu4XCDLKIY6LoX+glcQkCRYpoK9AcREcTEujbNfbQGj8OqeKom6cobC
yzPdggYBxWmGkxlId9DtUfBx95eZozyajSq48f729VePUE3olscdXggLDGsokLGF
3+2mGcPjfxq2A6QSfscncXk7VhvwkYolendMCAWFkEFZb1HklkRiydX2RYBgDEqv
bLaK1as5hPv7Be+L9a6Fd4bRlAtlsrmDfbyWR9KItlojJ0bz/d1f4flSx7fp5Tfc
xZfCxfibn0SSpTtyGkeoP1AUJ5ysRY60TL9nx54l0ZwacA7pSFpak1EEImV5t17E
utAyV0A5oyUtvL9W79Dhu6x34X1CDoPeOqgYN42htpX4qbWhAnZKBi2GQkICImqs
D64He8hAqF6URn5vPLvYvBuyy2fCjiHp9Up/xMRN8Esi72B2dEHvfl6WpEiOT+qs
QbHWlvh3A0wDbhzddRxTq1LqzRIdCavHd/cH7tqWd/AEJyJKPHQuYCPiBWrRoYIH
f6+SEssak4j34FzfvzZPbGd9JPjU4/OUq2tw7sq/BE2VocymwwVSiOEC/+rtyzHY
wJWxUI/+wQGJH7bx2wmgpZI382rvcllTOoMeR0Nn/TY=
`protect END_PROTECTED
