`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
nx5nqEz+tksjSGP2zpqY5+0jd754RRgr4EWLuNUct/nLQVVKfYLM2JTOIEftTs8n
LkhrWSy+mWMJZlKBaaR32cgEJRK5yAPSbNJ/a2K802qhps04gtf64m4K+HwVaiol
kJ2xvIIFehPTR4dmmRfltVBDCSw7G6M/o4tyHNekDj1YuUijb9AEP3CYMrEjWoac
FeNnO2OXw0P/RSYZz8zdDEbrqfkcU4OLFVgGIIFfllaUITE2nrLqfPM7X8Cdisjx
+gIjQj3hzKYxBJrQtR8yI3RscaNZfCmBSCCSnMRqUI7byH4rbfpeygLp2MsM7EIH
ZG9iVL6cHQ+qFjo9daKuxilig/WWcTzNVSXFfr4/BCyz8hp1/kUPkEvz+vsoT0Mb
`protect END_PROTECTED
