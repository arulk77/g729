`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mvnjv+Bf3VRXasXs/3J0gdtAXnadsppmpjgY2OjCaxzvTZxS2tHTkO1C+f2H2uSd
54KqjEQe/OIA2wTfKuEfOmnO96f2rddHalvf4d66PjV/app/RZNWY8loT+CzntYu
QB+JPPZwKXCUxQ8xk9aR0VPEhHyZ2qOLzjj/ikObYjerv8tJz+4l2Zg+iQDkYzNM
bGBybLC/gDHfDiUAPbz0Km2BhkYQ77uhmkF/c7xUSc2nJBGVdqQnd4D2t3KThbwT
dSz9qYBYR3hLKJrNNEPipdh+q/Us7dzqzb7pvLOzlwiRteEaEV/f/oyDv0QVDrbK
7un4Z5SdqeZsUezMLLxhbUEJgHvKniY6BVkXUjkPP5HGS7VDcH6LfT1YIC2+bfvX
5k0UkbFwh1EQs9hbkqLuw4bubyF4lOwqDZD7WZodKm4=
`protect END_PROTECTED
