`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42z242Hn8po4TRYNVvhUOZfWECpC4CTmv+nInCkMncuq
v6TNTdUz06sKWjNPJQ5RlnrerNAp2EGcOhrvaVwQXLOx7P+BdCy7lzbQPIjB/qsh
HCsTBqp3fRWT2e4AH1aANdNs/cihi8ANrK8xtD+DwGNK3PwSWRISIEwRoRml0j+u
+cLGFA5ccuZSr2ObZAfOCCVspOKaXjETd/C+0vOUubE=
`protect END_PROTECTED
