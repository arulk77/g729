`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKE1lNxODc2qVFUVowGsKLeEqozjd0/VMNCTunmhOyL8
4Bfo+fp/f+BWm4o59tveR/flVnemNBn6KFGbKMuMyXTQziP0ekeeRByW7wv+qeT1
dNlDJoSonFtPSjKJOh2hr8fGTVI9te7euub8fcZUGDpX+WyFfpjmDA+86OHQAju0
w2s4zU/rwOC0U+LzC1YsRe/zOKX234d6ErtYP/F9PY8Vd8sc/p8KparFRcB2O1L/
Rq9Kh0Sg02iQZDdTeBjqWuueXAsPBkPSAGEavPN43SF6zKD+O+uVJ0nqs6WTu07+
AFWeuHa4V6IzBkOFzbZbdYVGisXOD0x3OGHRtjeWoVNza3sVLEZj+XXqcwEd1zuq
zfk+bRBqm3xMyo8MRuI40i4UX0+dMnJNVLMGam/zG6+XV7IWmIpkLyu8mkrBtJH9
0v6/KloqAmTJL1sO6ZHFwuSZ/RO4D0jZa3e7t8ZPGDqtjg/DxgRV8EcqGimDEIc2
O4u/so8zXgajIxI5nGnb1Pn9jixIbDdUcaKtG+c07yByLUoE+Qe0PODAo3vjv4mX
`protect END_PROTECTED
