`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4001P/JHK8TS2Y8CuMwsdLuybpAnmdrD4qYIFbpWvPQ5
a8McvFXlnz6bizkDd69dagYHeQKq7aHLjE7lNTRGhetzNZ3VxGztXDWyD5GeTpwX
3xFX7wnsT51IYndJDlyVQK53pMda9FVkrYKvK1SMWINLJem9/BAOow0YnbcqmZ70
yYjycFD1bEe1O9alQwTxeTxUqPZeYtkwMm7Ok456Hk8=
`protect END_PROTECTED
