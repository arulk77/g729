`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
maM8AzMwVT3Yd7tn5kUPAGHKnnBHrWAjyBdf4SrHzTn+Srzst2qwcHux40hwIkw5
PG6g3IIcLY0n3dczQzTJ0npjmQO4Dx/ndSp7fS2uaOweYYSt0JXGP270G8urAgX7
HKzLN/1oyodU7y26IVMK/4cfzzJep3v7lLl0wMebtSjh1ALVJEBsjaliNdw+0n7P
CGRnSXMoACHUaia7FVHv6l0I2VNq6ju0op3U3HXgnz4v7a83dU7oYvlJAP7GRQdx
A3sAX2zMTYJML7RD9t1gfI8ZD4F5nU72KszoiQxARbj0qcItX90lLElqOPChOHUA
9bt96j4T+URnddLLyR+6QgR0rbyqoE1hZG9tmW37FT6lDQw2rb1j1RtoZLwxNT3x
CvVLd2mZMUjB/N3TQ4O8ZiYN2sHYY6qRF99GgcQ15Si2kduy3UcEH1xy8zDQO5PI
3AQCa7ziYDgGMid0scwHfuYzLIBrakoPtAlOicUTrYUKNOtmtPX5qlXkF2tCWXzS
O9UFxaHtyAb6Lt4pLtlmnPpTbX+hkoZO508XrG6mAH+Ovd8mDtrIpC+dLzib+Dgt
Aw93TZ0CTuQrr8MRbE7vVtl86st3tTrFB0utI5wxap8Q7gRAa7WKv+Pbbk7xNHI3
373yX0UsmBNc7E4wwHaOwVKr/6eOK3Rqi/x6x976CiHSwX55NIidV+VjVxxuwoUp
LBqObHBHdF3jyb9Q7FuPph+2pNXOAUxAdoPr1J0QoRM=
`protect END_PROTECTED
