`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
t/+GOYPCdGCirYsHrJcf5bfhuH7sErlOxNhu9GKBE3I2VqhqhqYjLXFy1TKcy4xi
1Tusg4IsOVp4ZkRBA317P4T/SJiDPtJZfcNUky06vWkhe3w8Jct92HLQhvOKZAdT
XdLpzvDWSmLlLvRzAoNkb1q7WjIlEpq2Gc/qfWwyn3Pcu5LkE/rvnGxxFx1NAuqw
`protect END_PROTECTED
