`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
zGotIiv4NqnlwMMoAuY6AlKBetecODXuaRsQcuc56u1vsAKCOH2g3+WpIKpg61A/
8r/bV2kVsMqgccvQOJjOzWtV3Hr+KE2T99/GnQ29uHtwWhYXZGz6D01Qegzjd1mV
u1TxOPNXOnZ+S+aR5oL1XMJI7v/D1vrJTH2XGBYStLKRdBdJwTUVVuAInhswu/jU
saOih0G5jfzik4ZMnW5lUozP3zfv6bn9TSwNJQQi8RMSCwVy9XUk3gUr7jzflTBV
4bKerYmllbAGgmv1lwPvxnIUpIl778idi1gK6y2DJI1i9vGP1fCtMTRI71AtffVE
jqE/QiYshUDJGMNIKOPnu0oOtKwMrqeDHtHrAAE8zH45I1ADcvmAtgfwiTizQSIK
NWWs7b1ZuQ+pZ78btVGMSgN1p8OibiJg1uUvLNI49gxDQZUPeBDrTbTMtYa/2WmR
ZrYYJdPpirRiKEvvvjebA4OBKOomuE5Bl3NuhZwlaC0OoDd481KZxp2t+i1JMoaJ
AZw0A0lw2pGYQZ02FDyBAsDHG93kFALbypz7Z2idasXeKgdnvIS9UMU9mQZpn3YW
LuaHfE2d3qKDXC+xXj9oHOuw0zmy7Np2U2nPOStf6/tyI8tT7gRnPn3gxexZ3pYe
kg6CRRqdF3h+AdzFlkLta0973/fLgt27tbcokmyrZByE/9pOkQjzcRZOyN1Gb3D/
EzmEIRqFwUIRHwU+A2IeE0EeY90pK4d/O0L9YIGlYN5Xe1/9F8VBXhTocno7albv
ZuA1ZYeVMYPthGFzax+FbNb3EFfEk2t5HCaE31VV2v5MkHcRJ1b4HrLq/Onyae1n
AlgXkLwCveWJH5Sla2/oJAgp4lnSTwlNMDbKpY3u/V5mrr2PByWB4nGmk0R2tTPh
6QnRAr1DTgS/kYPmaebOByk5RAYn9GerYdYnZEE+EMERdyfGoX2AdDalYlct17+I
TTAn1ihIjsz5sanuoz0i80nR+UwWbptfj7swkcCMa4wKz/Y2I3M9aM7W/G05WAa5
l22ZH32oiAY1RxWjf3jQH9RDpveu1PBC/W9ldSJhFtJGtffAjNIkYdNlk6e7EYLW
oUcMrXGksmec9GQAVNp1MQ/GAEO+kbbiKDOqFcUSZLTe8VxRVxJywsoTbQ56ZvLr
U6yHBtNnlNJjeM3aaiP/SkxXgXhWiJG0i2D0z2mBix7yU+d8dfoYM7kqmyjtilr9
4BeBV+Tkq8KLfTznQYof6Vpw6BFOH96SGJjcEBxAzGDwINFrmZ4yw+UMLgDqe55k
faVda/cx4aTOADm2c+54C+f+uD3bKA1UYXRg94tvllFq2DiAE+Dw6yBAdYlHuQwh
U/RtoFW+YynRxQL97ExGER+r4E44uk4XD6yOw932iRcbDImc2abx/Dcb6F7CJv+O
AWrevsBbOD8qQGUke2OV2czszSI7mFWygbpHEqJNzL2tMPcS7+7UASHcEC0C+ig6
6j7nZyt9XFJONAsW2yO8TpOwGjHKdxAZIIRJYDxoQFXukHcugiYoV/nuii117Hkb
BVaRSDhKmc6dhRhIRIbeMw==
`protect END_PROTECTED
