`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43DKv+b52qurI8m1ZacdVKS23uZvdNN4q83iqq1kuSjz
Alw79jeS65eWQlTCvcuYH9HhhNaL0KSdwFwgUl0+WPMaSSecDNb0DEkCTqg97vhG
ZgkDXqaznr4aPFfLzN3ETaYuOqN3vUMNgnd9SfmdoUeYk+CoDqKALo3MU7aU7m/4
XtNuvvhwFJ6tBV4D4xbfhMO4Z+/kbYCt7CW2DfqQybnF9lZPzlYYMXHnEgdesC/n
YhqfYIJVC33eQGvxDp3h+KCjP3ZEQUd7+Iu13DgycOo=
`protect END_PROTECTED
