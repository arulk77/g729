`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePyY16tsgk3+kAEnU/V0jTGqwuWx5k5BAN1da0oKlgnX
ayJ5iia+TtmeZoRLs27Q44Rk9yad7pzkP6Qgi0FUp47/257PekE2KFvGlEvxPPeR
tcznzulhaeyrxGDAgJv+LWHweKIgHYzor8co26LUFw0RhHaMDLXlRHfWy6khhJxl
+ltJ+iGYbkLihWDX5c+8B1AUg1sErDXwZ/7jvoyWpjCNDLbRidCMI2cXImHR3npL
w0bItvY7kdDJUS1xR6FsxzmvDthiwmVcy8wDoFJdZCq/S+Jom2JfQ+7rCX1SEMrf
+YeAi7C4BJ64JbKMkbMPEpaVycmmnqaQ1Ww7mocyOz4KaUSjwSRP0Qxm+VkZZLay
rc8YBhg8L+D05SonuF5S6EqUv6mu2E0HDoOuoJ/j2ghL0ZZ8oDXiilbx24bnGpct
+1VAZzhO4gLv9bkzGF/Yrd593rbnvMGAYkpV2P8OlpPZqlWgYSFvWr74lBv/YHLC
ITpj7eH2arTk/Q3f6pDqHhI+NeGOMW1Ay2ITGdNQ+zBvFykMEr7EGMVY2ywA7RuP
`protect END_PROTECTED
