`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNty43RgBRSXVZDoKXHifT0EYLKExkbyTVl+oJzp/2oU
I/fQmXG6RMVO7pS07b4SQ1TQQSdKueipA8HbDZ9r4mqN1lhd79MW1ePiCrfOotDY
lvQcPgTqAfRI3B7pRIY1zPF599XP6Exjl1viYfrhfqHArWarzLbLJOc2SEMBV/kT
e87xMkFI+euv/ZMtzEWbxyeqW8qW2/Dykq5Slto4vcfWQE+5jb6pcjJG8+NtxJPV
`protect END_PROTECTED
