`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Wm51KrEokFJkK17ihDIZywl/qnUWU/dI5sNVoLiFSB3UqEPSx3GE6tJtYnA+JWO1
4ZLlCvMcmnzx/kxZmnUBIFADEBkUsNK/v2rH0ExCMX2T82AgnRa/2ldPu5/x9riv
0WXz0xyDlWQupWLb3lGXkqxbwHqG8azMsKXht1/KxIR9a4kElZUjUWgVXjtcoYuQ
bM9ATuZhQ8oj+gdAZpQaBJfrBSfMmgZ9Cy++lb52jral2r0drTZNjqw8yv/Sk95p
KQ8mpec+gKayX4pvsgHub3RSNR3Xl9YZu6ZTTRkXEl6GiCEunsAYvcpBaOS3HwAv
9bOXsSO455MR2qqcRTEyNJ9ML/yVTYlzYFt0Vup3NA34VQXp5zk3D8tqnMTQaBqq
D8lxm0sJelUEceb3tJyxfaAUMBrqBHN6uMqFe2sM9fGcM2vFYN/ZWEBPF1d++lM8
xOjxJTGFdl845t8MNMsfULXh0Ezuhr6gtp46iOs6I5c=
`protect END_PROTECTED
