`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yreePdLh1qw87XVkLfmnf65y/7dlxEroctS4xRD10p9
gSjUkz789Al/j/uwzn1nIdFBY1btR9QmZEA+YBIxekIbspezmq5gVKizNAMDz3fO
Kwn00UhmN7avFicSArLFUJEA4O6J+rTVlGnjpagRAnHviP1sl8DfklDIy9RZCYjF
ppUxGr9jlqy/RJqBnOjDLlW6lJmoY6MXVgiIBvwZ6+jWMaqNQGyIjpVTYm/8BPyb
P9REwpQJryYpuBQBUOSKmLIFnM2x5GA/Lo9/tbVy0gE=
`protect END_PROTECTED
