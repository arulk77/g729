`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
KBD18r9Q+QpJIrPMFCu+kEdJ+WM1cnBQ4pxdAUOcZSkZgEpA6y9ZzTTX2INlIYA0
PDc6wnwaDjHjbe7+SEzJFnkAYbA4/I0DR8uilAzEu0VS2ijWhos0MmRXyA/VFWT/
1m+E3oNNGXT2TdycQE/zqtcMr8sp9YV4SKgWAcXO2E/5pP9BLR6Pk9fQaGPQyPIX
8qvMLU7+hVQoHtJ+3BpfPi+fjqbDn1Hfc+72iKmQhxaKCc8wzA7teGFak7uBTTru
rhr+7hoAn32Gp/b9OEFZ1i0E4Qhectj5OlF71VpYoe8F1O35ZxrADSkbjSOTvpuT
/xucnRQsKeLx48pKxkwwFztqW5O4Hc/Ti1NqE7YXNHcmEPWlAlvAyKxMApZoCtD+
Se+x+CB0go9d0XPw3ilpp9TNUHCPIHXPgf5p/at4mzLIcrFFoVYczNOwDa9l5Y9w
KSlbpDIeM1SHuSZN2TJ0dnYLHvCmlVjOBVpYM8QaNmy1fwpLE5ZYGSd6jyaaOszg
GsNn7u9ce9IxcF26xn04j8ajhuXl46aGam4keF8Mmpl+pFeU2Re/esS8nD4IbYyk
LhBfQU5qfTDtZKuUNgPo5FDKcI9/CY5r9mlRtQDCAhVwpJLpK4auIMyR5fDbme1o
YGOU1QZvN/1oTb2MUbV1GI+Ge0X6/Ji58/TOl0hevzAYocodVvxJKP2AO6BpAkTS
EkMMiwWvyvz83gKaT52KSGQpuh0H4iXN4SPQfJU4rCMVXnipiS8C7BpjyfOTveAX
pg+xVitRNPXh2xl97PZiOaFcWI6qQeqSISWdVasTRQhgR1Xwws/8vpewcWNN0j4U
vgO4v12tiJUka/LlipGDgXmqngoIMF9q9/z4FBaoKXVZQJIBfIDaCZQDbcrCGyHQ
jbiTHx+q3ncnnxD4HY06mxaFOKYCIErl7vsdwqeu771x8v91bm1Nn/9MpLg1sFOn
FtmJcojHWoAvzDxmr5YUplS0uheY6GcRuGCz6PPfNQagbvnHVm98Hhfet1pEgQeN
UAO/vRpG3d04Iyqqr4XgBlsJ9/3NH0tHmTs5Rk6f8Y2jMX74HercHgIWpTUcR1Sc
V2a7erWapncaOIjqfnV8pmIDXVqZXePNtxY2vUaTkoXDp1jte7pOlw7IWLI0ShX9
5k4mVw7pG2fJ7BZTyXe5DsBGEY23jkcf6f3cg/7eAoacUc9Ma8prYis9dDOZBMaA
9XT1+j74iC+FPtgwkBLjJi8DvnZjXkYgo4ctxcoZ0NVUPA4FzO6NPrcsXDOuP3yB
TR3D48frGOiOmJnnT5a5yMjqBR66rS9FxOZkiyIWXoJ2Vbau7rL9h4+ndXY2ESYZ
ZUbwICRz8B4QzAWQ1v7SwuotOFxYU7+xjvLBMUK9TuSsV6/aKiPIn+nhRWDymz5z
lnVBm0fZ/O+0o0cYZkMGQ/B+djssI0Bb/mGmSpz6lUR6IVgFU1mXcI71Edu2jFMi
3PgIdjUjodIsyGt0X25l6NSFvQi2DFdJSohGlyugpP5aVe5unNK4tfvpu5k0NiZe
0bh+KTB03dos0Ra++MRapDQ8+6gap0Z8E35XKpvpAAKBqaofVd50TAbbIz4O5STZ
9N0ua8TBNcEVJo7Bq4BTi6BkU1w/c4FX8LsJS836gMSpHKvkSZQVtuyjydcd0vtq
KKw4Ot8gEn+wFZlj+LnOrfvA+yRwgY9yO65J/T2/OBfzRIzFIyJItpGefKFcwPhI
Ntck4T1NJgzP4SKni1dWmAuJROJP7RCTKqb3rqx8zGurL9jF72WKPPR6CQDFKGTM
iqukac9+Jh3/Djp0kEqthk3+Ob3j5oka6L/jFX2foE2sJkVZtLf3DGGfO0MDtmQV
V0+6EBTa4sd7lewDA6D8wzNusqP0Rhlu0lx0YYSwFj3k4xAG2aEpDYtsSwmslgtB
xDgQHEkgXJmttbQkK6g/FN3zXgopv88h0iWl0N9BdVPolxhzE6rL+0ZKBi5fDNtQ
KMxKQGxKWeswH1xUFehiTsY8zHXvJqjnmtxrhXDmPkt1qLWzU3LQda/z4om9E6ok
XrTYvVKD9+FH2zdimzSnx9JmsAqb3KbGh0qGffZyyDW0E8+bw829/gOUL6+6dwcy
5qLY05Gp/i/ydQ0+aXgGyO8iw+5j50C9Rdr9dTrAa9I5K/OCaD2t1e/90/mxFMat
yLmAPUyPM8CFPPGyGP/iklsWkmeVH3FhJPmjOY/KccpNyApzB30giAVneQDNYroI
TiLRXZpBr2jIrlYog4SmJ5X70KCqhcm1T3ERt1IhaAlff1nsavfHaM7AZhEwni6c
GdkF6xsnU0kIRUFniLnoSf0p0RDpIQiu2vNKGDHr7JbDlxaJmxuwULLl4Ra+fWCU
8s/Jk6hY5D3WNrAU+zV97+ytCm7ewHT++ZW4hJ5Y4zf8BGY1+hN6S8w3lT8G449m
FoqJo5gATFOHF0howg0FKDxBy76FdHJ7MK3q6eVBfjHX3BfuC+lwfedA15JaydAf
eHvsvriRL/iyLxFl6A9pvEH2SMMIgQN5oSOTsl2TcgsnhwfhKSsl4vzgBMnQKmqC
8vHGcs+afuHSc2XGrsKhHtym0/fBVhC0JG8LHgfo5H8Du7Cfu4DSFfd7LvD/RCu1
vvSjRJT8dqIaqWDV3uTm+Wxe0/MNaoj9K2ebkEcldYC6MwUM2I1Hi8gDB2VNw2mr
roBgK0Aj5VpS50yI7Hi6RGb/2H9GIWJ0kS58QhvCCsFz0HXKGVoK0j+U6wjyW6Mj
qwRM5P2wr1auHU54iOTr6gsSr63jD0nrYyY7kH0aQJNK0ia/xsyoe5vWiOtmRmnl
gqWUW/iHkTjaxbQsA8YxIQa4r9NC1F8FW9BDhpoDtHmNPfV4xQWTGBmrdzTE2MNX
wPy73xySd7JKOiahOaM9+SEuPVVLZmVS2d2gJGjgMkGMuEHLJkJsjBwP1CeNkVtN
OekEL6HCMuRBUdIVIsbMtVvPQufQPB+TFhH9pDzPyU+HsOIXJl9fRssHJY+hhX2z
LIEb88DllacYczrhr6IJUXgIOsXhiOzZpTYSkpUfxmsUcSR5nYnQAtJHjkI8SPHw
8GhFg/hdvR3mgbhY3/NulUHcEOmk373MYB8UGTxqHsUNWEU2us4lAzZQO09i9N+U
8mwoyJBSgrY6oXyfL8plTefi7Sy8/USJqvwK9upltbvR3yHXZvTpwfQZ7vaHHGel
veLjSeE44zcL5BiLuqYFEA0oW1Ol0hMFbVX3V4gWusQ6nzMD1nTSp29WMtVla6gr
GVHTeEbTfNMEZayt4z9QYnRvDAH6CnZQcg1y8LOWsZzlWthAaMNpDh5pEgGmMWRd
SvnUJVCJ24wvLfMVibTZ7/6cN6oMPUAJCLSOAVSuc6fF7rtV6QwiBc01I1+PtkXh
Nl/qNFxjEW27lGGQR3JLfUgODn+0lkoorLLAzlJwiehE45ixsm3K60WD4TyfgIGA
h87vWGM0ZkiUcz4k2ntYXZaAq5SfWUHgXJBIgh9JKajm+IA3zojd9uqnU1gxLKrU
8oGp+aDRNrJmDBU7Re3oBkmXZh033dAFpXlihdew0gSeVgDvWniKTnmFwp/zl7gC
/8t6e5JTn9FlkWAa9ElGNvT8L4Sr49byGGyAfrqbi2g6zAE41QIyG3mvlR6ztJJi
6MPj1eK/nY5r+u0taa9OFU45XkUgaSTs02LKu3UYDjHW/i8fRGAsycl4vrjFvl6h
3NFkfkKe2ban6e3VOESQDxWve+mmaSffowusO0IZmHrQRYSGbLSYU+V63AGBb9lq
j/c2CSUL2UDktGykbeeA2SYfWx0IC4zVQp/nNBdUmgECJAc+jQBASRn9jw9BfjvG
yvmKiqiP6JUDYBEY4DpDHQl55CwKyTmawlVsRy8upChklReMqg0mOjMnyBN9D6UI
4v/eAaHuZTrY9joyNjRcBLoBQvjpXQsVOM7Q0khYQZxK3yjPDjFN+YbUc9qavH4z
9e6vcTnJjI0hYDtkiloN6ZviF/CYpF1KvbD3uXGU1DEarL47J+W9v9/NcTFEf/cI
2I4mBbrrIPzL85MOcHdp6HvM7HGWVohjbi43roZbCBscXMckW7OXDuMxv3eh2FtM
2wpUr99YLbE/8vZF4S4sIQCeqlBbDA58c1LaWDK37Vku9QPmqk484t1dhYfPYuL3
6oIeQ4UjKhboN/gnyMUhhpFG9HpRJc8TmwRG7hijX5x21QFzCBQr1wgJz54a/T9j
zkKpy9oUNO+Pm2+/+ECZX0wTP7dxLpaOW1qTWZfuo/VHomDElIaYE6xWwB0KZmN2
mkz7rTDaCFRU6XxZnswP0uVrEFiGJeO5p4QIJvjyf8IHCAsBSg7AuEAYn5yFlCys
u5Lb5nBA/P76dzUy6iN5nO7oHDEnbUscR33ASmGL14I0nnMPDqUfmgPbOoMMK5JM
otwEP2Bp9MDqo3W7AQkKIXrf+99u/RqxD8RbTF4Q3nvrAf8rgGramnyEEQTjP7p8
wxaMCXWXfOyG3kYsQ1lTddIt2xr7NEXSS7d1UmYJGdK4N5Zu9rA6+f4j5dKw9ceZ
MkyMs25Mv1Lu8wpdEylQmMbVa8fW0iqXWjAT5gbC5Ii5pniLLwLnrH5I4t9gp4Qe
rA1KdZEoq9EMinpd2hiMImVhNgOmD6qwFWW4LsZVJxYleCDqzx/kJYoyFET2i1ni
wmkhR1RNhz/AGmQAA6gIlR6w8KJzUs6SClKTY/Cdi/4o+2N3nXzs4SoLI/cUlXFH
5G7mqCyZFjljPjtLGOMLOiTkL8umDGdE2AWwkSpz4QpRpz4Iygz01L/tjo1NutRy
vGZYJx1yhngnEgRCb71hBB4dEC7qqgU5E8P7A37gZ2uThICdnVTtLhaIh29+Xmez
XcsTTruEPROhHwM182V3xJkK2PQITG8k6UKpW81ui3z40M4wGEJNjZDhcee1Ckaz
GiMEaARPLKQbyHMdpUIlonerg9cTTFW2K5aRAeFx/EW5137BLi9gzTk4uqVnypUQ
NOjKnpmY3aM7hMIzp0VV1jyzGg+MaxpYU5oYtmvBCLpCqw56zG/ApPq270kti66K
lvH1pFV5ZCWDDfLLwjTmQBz1q4ZDjBeq99x/0C2veoaRPvp1fYlvObLlRlRsQdJs
MXH+QmvzUwZ/TpKluzx4w1HQLI+Exz1DCAUw/YOLj2TqNp7pmFWnTd+LErIumdlb
+9Pk3CNre6QXino3YJvWUfZqr3/pljm1SmRkpJbifjssgInB4wcUh3y65clwOXMP
9yTePnTqqnLKAK3EZuUpP6UovBR96AFpWPoWAXGlec3C8eoATaUt0nYZRBQBxSMm
8ghVxAFPkBKXVKsbeyBfj8rHfaf2LCw9qobN4wFGEQn5MOQq+T7hBmzQaW6HhmyR
yPoHOvFGnnsBMWqmo7RFNuFDEHnnA72mf8I9XthWnixXDr4HM0vRtlmnpbrDlnOz
go6CpaAp4CkAhtI3jkSDe3ATmuWr6iKve31E6+QhhJIB0yy4bN1TwwbRHLkcMuuV
7XmQBCTYKybfuN6Vv/TK1JBT2wd+++tRKn9Z3pn679OEAY5Ws7/IrZHmbWr4ihmq
Fyf0EUWQg5stmEwM460b59VJiGs2SZbD/WCKraz2pRDC9jkzfgF7ikZlOh7wSjl6
UnBdfYVORCYFMn2uWzkxoJM7U/+DNrwVErbPExkxqpdQj3Uxuuf5dxZiCM9c95gV
vIbQ0HHYjG2N2HxnAE7RQaT3hK3B2zmI3ua7/8jp20eCJwouko/B38JwCzAZnepy
RYHzDTKIZcTDziPATgms32hBZmnfjQ3fd719/35R5vRpJcV+FMSxypj2fJgWsrDa
8Mprf4ge5xPtfj1M+MF85dQNpiJbXOqSVFldF2fkVnLY5AvhRXRCulTcUv/QI6rl
38fl3XUqQPJTc5gI4DNA21bJ2O8p8cmWqGHH0Yjpuwx1u1jJwnDiJ8raWT8V44og
34XY+VfhQkhNIkAiQXutOMaIReEh/ZcEX4gx6yhamFpklJeTH2YhRBSG78ixrRHC
SueHO+iAjgNnRae3JVdQ063m4tgwfoJE/cXNjYGqF/WTmx1lXyjHzQllyc83hU7r
CG+KpP/+/aHa23e6M2x1CUtdeHG3BwouSIBi01Vvk6OzJCQKnzsvjM595dwgwKnG
CagIZRkCREGyMi8VVooidzegnFSln74uFG+mTtewJ3kW5OVwhttfQKXjby1ysniK
eUXfUu1dMR+xBnDqfH5lMe5VKUcitUqsvSg8HZMDotH4A86bSDt4MBHclJN7kuDE
127eh6CXBUirNGZHuZZ9vDKr6bDfBaIkuP3RDcZSYvIMe64H06HSC5SMbEWFM2JS
5ReBKVdZVgFd96qe7iIwmJD9XWeEaZ5aXLhmjhOi9TMWSVaUBw/8bZaDmeyqGIqk
HIGLNy2I9ghbbJyriCiFc1z5L8/+URo1ZKAu/MuUyRyYxDRgmU1IPgfSyomT8R1D
xXSMvR1qnPq1n/bOa+gQRebCoRmiaUPfK+/XjV6Cr8rJUaP1a/uy+C3jV9/O7DnK
Dp7Gcc0ENwPvs1lwcLV6mk73I8lGUv7d+gu32i+Gd1Uayl09DBjFWaXUQuvULUN4
IxPjo9tSfm8ic/atkD7aOJR06uEI0sAb+ugend3Yw4A+C6ZG73MuZgzhHcT2CKz4
iCgGQ0/eJNFYktUgJMEG7X6QV9X7Byda5J9QmHo6OQCdyHGfyTgsL09D+hH5VYEN
JjNdqYzX4jdvDQYms1CQTnMesSrNJYFLFr3AX8xiOqkuQb8sJX98TBFk53BoaMgz
j9kVW3M/VlrWlnBytdLeeG1GOzTvJFV+EJf6Hwn/DK+Rdd/s/AqiTjQYwmTo08S9
7Gag/YFdSIUy27gbOTIqnbgzT1sp6lEO4R1AzQeRu2941kDx6QSsJcQiQhCOrqTn
889G5EVfeA8kB0xYuS5n/AVwhV+csmhyqMGT5LqD3lCcvqVmi0D1rvxXEdpNZ+Ey
6u2cpjOXZZJTaqfdNO27LhzsG5aO038CbZpQN2ADrgc6+Glwf2WTiZO70uHMqYDN
aQKbYVOG3+z6pIzz1V2vvhn/ab7uGiJMml2i8mAeGPaQV+WkMLE3lXA9h3FFt13Q
pd7mwUHJ5w0DXNSxe2ctNsTZwds/SM+u/H6fI3kVRKqbwNBO7jCJwUgy9Ug4Ci48
Xurvxpg1KDNDx2qZygtY+ayu9WbqJd59wPl1qI514i01e/CNEgIE2Jq8em+41pUf
YBHN/ny8M5KJL8h6Ak7WfZMLSzMOlUZf8Rc+J7e2OfnR4Er6SFpuuJNh0GAiPYnp
ltNp12VcAXTEn6xFOn5Cb8rWIlaV7m5vNcd3/Xi4O1o2xxBhJD/BpScFHvPVbV5c
loLiEYDCaNQMcUdvMU2D7eS4RirC8qcFNYugrj7gUN7L5xmZTFjY7XS/q88uSsv/
9NFBsMSzgS6nKYjS/HixAoOT/bCxY+cRzGOe0+pILFPelmU1fueHiCoId0K2LOVK
AFMbtPt42uOE+tf7eo8Kmnt0qsZiqV9yzSh6nGvfwu6CGpEmqwpEl8eBdfBtOwmM
pwuwTPjsDJW1ftRRWWcq5o9MrlFDoIwiZbICQMzLMW1Z1Q3iAljcuWXQXqnwZgS9
MPtw0gzuwILiFeXva5jbY1rGNsudVtOe3EDXUighKrcN7z+EOSGX4DZY3r4AzNAA
yZLFnTj6XlZrs9EvOtflNpnYPx2TB/+sl+JhD2U3HtnnapziEcy+Qph9kskeKSse
LLl0VCqaB262SSYMyrrXaToVovb8tK3vY0DO8wzEJizc9HWVHRVoxLTK0zj0F2DC
Y+l2EHcE5EJaVVkq/hGjLuQ2A8bVinUAmFxqSe5CDbfXjqTh7DXoD1Zfm9h4Qfm6
mFTvfAWpJeRz7sSLFpaTxEL3KRff7BvKzTl5KhpVJ6khYXtvlGD3VvkK7V3gzTf8
O/ehG/6y/vP8yJPT5Mnm+kumdnOmUEqPJ2IbgUTLbBBR1W8L7ujF0N+d8g3ewJIP
bju96pyu0OV/Dkz+G+uhlOjfE3g6ZIgFgqh4J9tfcl5u57iRWydJJD8CgOuHVaZ9
QZdyy7M7t6prf2G00XTfTP97S+AWkY7KVQ30P2sStT0xwI26dzucwU8HywgJSt2l
mkF/8sYAHKQ7twt+0OsKxfcGYPi6Fv8TuSmsb99Ztm2fK0k7PWvmNDWpzIfUyvfC
RF5ffyjhiTIiPK8QsDqmA5bViTDvfQoBCDgKjV7JOL9PBvYBllkCAE7ARqfEzc/6
plVMSC2M9z9JOtkXE5THwhFnBNSsXu/fYADUQ2HvoAcLzhYuytS4F/qnQvCXwEYJ
YX8kAVl5FYSbiAjjWPsmbDcAjRSzLOs8b8Cj3aavku1Cq/4S8fMbKN+3KJKXkSjY
apVFZyyhvHDyiT25UNl4m2r7Ljeyh3mcoVEzz6/5FdSX815pWdvgs0EB/ntL9IPE
fADurTaQ3gINxo5t5PT8F4btyHF0On6WOXvpYe2fxhax88rR/J4SVRUMUNa9ljvw
jSY4q9brLwRO6N0BKfdoASC9IJenf9l4XRs8nr3TRtHU+TDWVp0ALBLHafjEhOOa
yig7bm9MSPLQbZ75HUGDzCQEsp+BS0N79Nu1LdL5Beo2YeZ0d489jG7P46f5mJ5A
18gWN+5wDQsAfppzdPsptUP150zJLsie00X8aPiYtCc71q3qjidaCEhZB0VF6rJn
R5vTdUkFVp8+J09YWucECmc7ddRn87Gfjo8rdkIgGw/QpB2LkNPX2e3/Y5yYrjbr
+nsIIlaTcad6FsyW9Uzg5JwBNOpNz4BNUdLCE/jw0ufLyhDbtimm3Oi6ltH146aw
sX5Q34hY+zrMQzHZx8Mf60meuEadWNPsZxhNvEdEel41jwBxO6oRenF1keHWFUbv
7uQx/zLeJfdLj8d8fDowHqrCl4JbBpx49M1+FKgZkN1JZ5mYFw3KSqs83t6kUYxv
TTPc1TNTCkNaX8V6MhQPVyM2MjdlO+KHpdQbEIBrZtW0RHNYa8E4wuH7nUeyGORP
pQKMt1JDPYHWWuaxWUHmEGOGG9yNOToNcHJ8kOuQh76EJrzuUrZA6Y9iXLrg6HMm
oVRNbRcGYwl2n9knMyXNe1BH7bqJeUYWRVnl+WKQ+3jaiRYKIhVSi42DV2f83p4F
iN4CATzA80W3vd0139U/jXfcn8wfZJxcnsCQUchct4+S/mJf9L6Crugj82lIPXCc
D/H+i/KEmu2cDutrfEabXNFN52OguJ6dBi2yPkUUgxBPbCSDnvcie+SbesogzmBL
27hA2Tr3Xz2+WMeIkmshhOtwmaN05Chfm6YzJmxsf5Q4zw8wkow2cWbxyVB2gEIE
zfRF5keggGJxhjocaOFA+28MYyBaCDfpV+/s2Gyfvn5pnlfZgDHSCNhT8zZ4IKdg
VBUw3KyLVAp4/9elT/oBr4ubW5RIVvYAF2806R6MpZqFKLdga+kpw63owUoQe5Tp
wMAriSoiNNnmx8Kp+MN5F1pZjbnTtcdXxl3R/qi2mR2EhW/ufNlMqMWwmh7OhVv9
WMbXaa6fMGXYyYXm1uxg0+V6np/387qyKDMmMWXyivUSOLc2gCTAudVYMtP7eQEL
LOdZRfAYJhJVQz80CoZBf3W/qFTsUh5JEUle5lZaQab4hD8zWZsNNtW4ftgUcQB/
`protect END_PROTECTED
