`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xmbmTEwVmMeHpodiC99I1FRrWMrAsVAAuU+wNbNH/z7
xqWlCRBc+hTTKjJnbswJ+JiK48tvEFoODkdOV7XK/QrrFBlnx0zLmyrW1apSAozK
Dh40UCfyc5wL+VPr4RZDgFSAEYxD4GpohnyepIqN0cOuAaxDgnH3ewmYwWIyRtaR
J951mQrOEkX+7M927reb+5+Q7ggd8bXPFlnG2RxabuU=
`protect END_PROTECTED
