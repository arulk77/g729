`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Rl7N/mOo025MZ7+lolF3ibhp7ycc2pvwUhVaf3yf7U7naLXPcX+Z1T7VcIkADePu
+nyKhrwkc+dbR1lchU4bXDkccTqRZbGeF9+44gJYVplryG8x2WpGWDYPwOHFp7Ri
`protect END_PROTECTED
