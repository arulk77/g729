`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL4UsddJnxzmmKGLXA4LCnndMmf14+5GXM0gmAvF4T/s
r+i4twkZ30zwuFLo2/qlLf8yfiw+/g44ZknZcCtT4QTXaR5NSfmkJfAr73lhiIVB
hlvFUALUBoaNNPhlXw3MvXEZtna7FD+lwwVaPwfQjUcX1j0D65B5UvRR2Cke1qxH
b2BzPG13xVcMfeeJ36hPladlyifmoxCwAcCV3CI/K1Daog9lFS8fdYjDSE5tb1u2
L3FZM8nAfnPOY8ZEnNtvvB2om8ECNgqeIZfj2gJ/rs2uJcgR2oCUK4ugT+i7vt9L
12baGsZx46zfT3u24wC1GA==
`protect END_PROTECTED
