`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1adCl3pV3T18kptIZwX/zlOkl3iVXoCViWhJHYHjgqrgu
tLxhKgero4gBELJ3o9UPoBu6Hu0hBh4Qh/kFvO2dxQBR/+ws5jHt7/63dVYaj1Pc
mJbY/wnuxjLx1qMe+EfTBUUUZ2Ej1NGNA2ySqsNoBX/eDiJWP4G/WwuLd6mv/FT8
nuoiciJb8brr31QBDOVXduegBoqbKbv8Kj0QgL/Dh3SMEUmMKONsulfJkW2axaq3
mjtAJZl9U39abIBfb2yrec5yQ8VJaGO7m4Esi1yw2w9c7ELGtvqwnTNrpvHZzp1x
N6I872WcjEv7aiN/G1rbEd36ovqFMwEt2xr3SXTOxHh7fMSbZg3x8rvUJ3XhoL0q
z28psP14K8YhI5SxK5wNC+jCN1fFEL8RXuj81PT85fxqLMc9ThxDK2c4s7XqHLE6
OFBOh8390fzSvRxURgNu40S09R8VqyhZPVAXtyOZdcJ6+TeI3jJnzJZwK7Svl+8a
ryMEm0KJzAnb94K/6E1phOvix2AD3uGWIHePuxVM/kaJjyjgB68NP/Ofz7U8Rou8
oovrExTPQBhoc+IekMf7cFtp50FAy43Wh5Ecor2RmlwMrbLeQSq3xTVI+ZaT8UMD
JCC3yLNygUKoL/SGQ/oNQ/wTRYdsV4I3F6GcMlmONjPwNag9j0rXtoKNUkkdu1j2
ykoTjCHdEOwEnsMcCMXZPOnHqLwu850FV/okXwacjqzhJVq4aXeWmX7ipt2yWZKB
wZJTsNgsLmDH7hRwglHg4EuAuvnGTSCRFHUSYxEXauLNJzINMn38Q//gp32sxnXX
jHpYOzbrQtq2CixSnFvvL3JepWurkxWzR1A1kQkM8zmPCOEDXgls9innHbBBGktE
tqEjiN6/VoiHOK3FaPluHNYv3VmRY7Tnb2iujUTb9WElmV7w7UacL88BC3BDcJGf
pgbHFwS8VGdGTNxcv6X0pSUnq8UMUYvmP2hHykz70IPa4AbZ2PLf2yUY1aZ63hoY
a7FuYoyxdDGRoAxrYHhxvgjdpdkHmiPfl7WRtcD3M3ktkj4ccbGFspyiLLOCErn6
MXrc/4UtaZl1YS+y4CawetgRVKLYFw0Bkyz5EB6YWy/07rfUldsppJNAr07+4fad
7jBAx3GIdAgEJg6stNJ9fOyeg/fbjRKpizLcdLKADQxXS7z5PjWDfooeoB7//QGv
qHcTtKhxuZhZ3L3U+t8fj6JvZd87UM8My5Nk2qX6qx+CeoBIgnpoVmlOW6qSD7Hc
Wkn4p/ftviTCZTt5XJBN21FVqN5K48DkzDuRm9A5DfDHSlgS5SmdiNjMRn0ZVsnZ
4OS+uH0y2LpoVxN7Mq1Tod7W70ezguMfXt9G15huwcaQVYLztai4HE7cwJU3Uhza
/xXKRJ15FQE5QS5ouVIO15vTYZ2s/Krntf2A5HjvkXZv9qlOSYI2uVJainhwiuf1
cpDb4STBwWkbkGh2AEisyXDGrmYdB7FWSHeL3TOv64pBD5FaKT9guE7uRDdSgCjU
AmVsX3whU/AqtscMygiI2SCW6dHUScLL84owkWSdtN2KSyL5BUvnL9xdZb5AuFZN
fQF3cfzkmC6gKqTyDC6yNe7pFYuJdmX2qBwN0OMSRw/x5Au0tNtgeIKZ2N82XKSC
Him1M9IOe7HtbPh68vzSl03YFMM5HIXQSnYYF4/OEcnBvXbO1avv4rtym9Ihm/WM
ao+VL+mSe7hMpCgI+EG2iXF1PlScGkzc9U0OoM4TD+gAr5eCtM8MFuelJfpCDv1c
djqFX1/LrO6fp4YhnXu9CxDtNFmPg7/LLNUPvmUGWhEOfOgY8OgS00NcUBH9y0/U
NTdEP0CXd6yK/Zl+EeXepex5mjG6fB6HCcvvp6Y4xxSvSDH4F42cI2f+GXyNRgzh
ZVaY6REWr9NbEL+vXFXlRAzjGmO7ruSpMtY+2QvHuTUA8TeHeFwpc7yLSvp7yrRq
ABGEy41ZmbtcZ83ASDquL3nJQEDUi6ETWA90u6Q86tsClMFy1N0SFXqP4efV+cPO
UpfZ/MC0ERYDKCE9ROQX9AoVzbH6FUnW0CX5e23MOfHMgwk1HFQZfyh+0hGXN7fw
OI7Uu0P3orzG0zTE6h02jXu9EaAtElz9FPCnFopMPU1zYVTE9hS/figH5C7HHdwr
MJVo/95O1d9Rc/7235VIgMY1aHL9+y0lnAjG617upiJ/18kBR11Xle972ZOF8HLX
8yrbB5m1ZptD2UmISEyC9fo2ZNgGm2Gi0WIJ2fE7FK7Dbv4k7A8UAq6SAo8+Ugti
vAmsJDxWiyRd0MOGKy9VnDhtXWBd9S1VG1pAUc3YfL+E9GYS2ItYBSbZ+rxD/Pwp
QktX8VofZxhk2KtKYYED21YOoqjQOPyCBRhd/Xid5LSBOjjJ09KpdFvkkxD+O88u
maoigCgdzRBvNzfSrmbWgEC+zzu/BQUUxzmy01iVvl1F3msAOEGhTH2Pp8kaksbI
w67UY/dgp/biiH6Mu4L+TDqes8jAv9AI2NbkQ0NlRs74pee5NTwAVV9o26IfSxIl
34aNV4+0UIf6y4lJYhzCa0wTE799sWxHEswdq/wh7qk0O+wDAU6JxaDRF3iLjKpu
Sq2m1adEdIXivYOzi4xU6kG8Lad3NzhtDD1FGGK6ASGvhmdB9VoCLBn9C7gYkOjp
kFJ2cQNRlyAaAofonPJRqafEg/HwbpgOf4ia5TZ58EezPVhz9bjklUw5cR1PFipX
9j+NeDCuN87vlNNQTdxFM009iie2yMTBpipYyf34Ddh6ir7KI1Fs4IBwVLX7j5WB
fawP4YyAVYX36e4LDRMNbH9irA+F4GHU6OtdLwXcd7cfBlIjbk7OCs9w7vd2PS3R
n+Or2VSawj8BPhdtP8jMGK9vEOw4y7AmBkhHaMH/q15FcQiim0uadzVyAm9ueQB4
ps8dUPKJEfSOZ0qMlRki9YtHBSSl/dpssaaI2qICzAmbgsP9tBDaYvalCGxM/dy3
tbcNruNq6NYZZA0/cCtFuSJMEk1WKYMaZa+MHzGEJdCi2wh3bX5sxC7q7V4YY8oH
xP3y2MQPBRuD32++g3LkiaVyzDKAawSy8C6XG7kyxPDqRPickQvSzBuK/s1jwy3t
WOxprfuXoL4BclH84VV45AvkZEuMR3+JIaUT06JFLBlO9KhVnsLYL6IRAYsBz4Tk
D0IrJLhvZAZMGno4TFh5nZIhsI9zSXS9gAmP0xE4Y87clx/jrMyavpqsZ1ykHqQW
PkY62Bg84EtqBNl4koD3mDaR+nkhvISl0IncDLunjG7pIaPfwWnm6im29Y4cEPfS
aazJGOtjcmQ9FM8fxUDGoWjh1IujGx0z/wCZf8FX3uK8aNCFMb9hjQJB2/33Gy8C
gMMtOazfwG7aXIaL2qg/fwAfx/6e3kJ6JLMGsBPG6DCHEb5yr0TUWwNYPN7EMrL9
Iz9qbBZYUwxGgFEtLAkBXppyXwQRMrR0IXvKOdnCoYKhKNvMXU40IcKVNuJQPpnG
9EGZHv/OaIoLDLke+H/e2Ij6AiCMDpp8tu0v2I3oMU5T+WrrAQPzJiQasZwpTu/l
cICixa442rWhUPVXZEyWk6VBDCOVsI0cr2/JSM+eq61MyvMnz+UnEFTBN9K/A6Vn
2S5VTyMbeF/K4JelNRIvTAxkuvx9oi6jJLve3u8tFNVvpa1OvqsN5MEbUEHagJPJ
j6E0iCo/v9avYG/FS7HUZucZg6TmCTlFsdqyieTAtEs0rlTkAsZTUaK1RJ+LX/s/
eTPc7btr31xd7u5579sA3CpEsyX12R1D9Z2ra5O4cW1it33EgjHFloJTCYOTRzDx
Y5SSdVtsd9NhXG6PjYjpoGB1gWknskMWBtLzgxJKFCxvfh5jiWzXSBPxXc7GHNEN
i04jBftCcWMSge1fKpqDW1uzi9UaP6f4QwamMsTwGpx6rP8xFXhppcD+9txQeVRn
rks4Ba2A0iOdUo9O2pOJlLUqrM47yf1rkEt7W620OTo++Ycajqgcb7zECex9uVEp
N0Hk1yhBMGpQO/yp/t/KPbvdKfJdW8OoV/JRC0P/10/FsK9aZelpqw5bvKighamS
Mj8vyjLlWx3S9ftJigJ38CkDt6AEu5wk62jRtT4AUImMvEHSjRD+MSX2DgfdIrow
qVit4xPzZpIFbGXPCLADGKIyJLVa6pEkYP0Kdbo1XPhpuhAiUOwKYlDKz26HeAfe
W7MWFzXwWyrSd3V0O+uiJ/59012nIiWDn5zgy2X+wi3M4xSN+FYKTNx7AAUEt/c5
giJeEG7lxmSqaGESkilgU0K8Q/NQjHsE6T4Czof+YOuzZdQd8shha1Y8htmG2+5T
QTOE8uY4UAN48MvM4E2PEhnsB613MgRvGWkkp1c5pD323GNX5rav9caaeQIHO2Qr
PjEfxc7qgka8YNYdKfgt91hU4T0vllcx8QBGZZm1B4Xbfn/j405atTv70M++MLlr
CK0QcsJm1sk+ykt/7PGhjaRHqmSViSOjNOpmRFbZJ2v5EysbIiGNuHZ4/lsbfT/9
lwmK2UK6MdeyPO606K4Xfnh7H60M81CMQF4O0HKXhl51t8m9b838WXpE5KMOWWWD
dzkaH4ol46dIhjHXPIEBdfe8u7bjsHFRn9EIjFYjduMQpmqYj3CYof/rL0CQXnjF
Tn/MBAodPlEi4wzFC+8cyYtqdG1eXp01QVa02JJKDsZ9v1gera6NgqULo/BKDQSw
WVHQs/pyGjKaS01wFSIOEGIsF3D1Dr9ZPbOoD1sQiYlUvkosYC9uyg6FJxdU17uw
8vWjMBANxSRlbg34lGZnt/bqnVsHT9NPyVvywU+IxoljJxFs/OBhcMAAVGTR6S2X
JzTS3kwTmser15I90pKoALpm5QksYPETxXukWRo4jE8aGQVi9++6cfRgvTFWTkTb
lPeWX6qqf+IufcwR/3P/emXrQjWugKXv27+iWKJzRGrpwTTpBecgRF4aZ5N7sfDr
q0rox2A/zo5OiOqFasZgowDsNOiWdRQ2ZstvqLHI//XduOB/OVDXTMj1VjTGEVs2
`protect END_PROTECTED
