`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFTJQ2YmdR2D2qEEzLr6iUuSHBLPr2Ucvrq0Qh26IbiO
y4sDDr6QwrSlJrBAy3JM62uh6K0lN0O+CTi8pO5Lt0EJ5EMf0U2/SXEKFAoA6Vhs
iHKa1zLQELVk3E0Q36Y23D838WLa7Lj0Lx01pMyOSlK+Jot55ekedcOVFXrkIL/R
5JAkA1/yaH7+u2Bfq3soaQ==
`protect END_PROTECTED
