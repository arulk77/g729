`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45VdnVOMfQwPDx6xT6Lfa0eGp0Z/aq+VL3EhI+cANbQf
tufcWmHCob591mU9s0CJJgko+tSXHYNRnvyk2GfdgCcTMPsdE//pEt26u5UOVMDB
D6KBKMgE0WksdwouLQ3ZLtvB6SwZaxxFlKornNm/E+pBXxEcdO2KFY48A4drXcNB
ePU/noitpBr04PnqSYvv0wpdPjCGd6bn6F2un77+h7KLcgLUqk4KQ6+91m9WIS06
RYu/Xo6P1XdWQpkAb40O+QXtNJIFVbKSrMq7sIJQ/R8EUJfJPQLheKH1u6m06vrD
OPfUFhrsc8POUVafVDWJZw==
`protect END_PROTECTED
