`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkZkErgG0hMRl87ZjrwRUhG2gq0Na5csM8vKBBW5CMMof
TlLecs1yZp9wwRsiQChGoBuK3prqQDhLOwYcE7bP0Y4WUf5QNlyV+uIIk9ZxQW9i
ij5rZucPSyXsvld/aAfq8IU1VkOucUYCRwWl9/7gVgwHG8VUtuXutaM6GPX2PP4V
1j6h7n/Xe33W0mEx8fWOywptWLM3uGgTRV+wlhEQH9aiK2tgh+KrTJh3wPUbnVir
IjV3suDWaSmQ2myzVAsu/78KDZul9TS/sl4nOuZYFsj+6GTwEXPGYahWWJhdQewX
BkacYUB5YIV/a88d31Y4A9a3iyzLPleBXG27yV3W3L1JxDYkVkoUPyyMADVSTDWJ
nCl//6J7RnN3R85wOxGY7kMN8JCLl3G95YmvGHh2yuY5BSwE+VB7GcpgVPZAhvbW
iIEBA76qhMItqDdfqPQU3DL4q/t8Mv9rhBcKvvnGZ+E1RvTblbSzl2YQi9dwvpJ1
dNaRWKSfmb+U7/oblkDVhWNwccOZSX7YVdsJTGJZATjZHDCbWFFJ5pdhaae0dJMF
LXxP7Kxxukvxx1Eqxln6JqkLvlrsPrSfWf9twHzt3k1eHa7oavbFoY19MkaatwTz
7DAyj7YmibpyJeTSlXUrp/4rmyh9nzSP1x8tJuaz8qR5xlSnVh9tLCJzNK7B5cmx
yRJRRNlsfiUNNxYQJ4arZmbckGrkRwQYonx/5XPbtskpp1dk+HszSSUGVeGdlrhe
kIri8p3A5eYVj7+PK1Xv2P4IvRqYcXwRlO1CK4cXPN1C4Xdi/16kt0FfcqdH71uY
ZVbOvGnXh7l0557/vAnz4Agf2OrKQMfMo/3FmbXyjx1nAui7s5dArqRRncxGScIt
IfzqWmxg+W3Usn7s1KFGpRE/vECBn2J/x/lJQ3VBvoqhBhuvlxmSIfoJaDMuy0N0
Em1q94SHvELJI4JyPrXBfW0cfbiiBd5xWDdNXu/m8Dm9MpTdx2lBBzYkZHb4d/oI
tL1VUapIodEU7u6+wT8TbTW4T2P6C25VPknTMrLjlBQPoR+ZNfUQzVL2BKrCRAXv
8Sh07pD12cd1it++qsq7SQ3uZVtY7R6QWCAB85P7AubskfGjquhji39QrcpY4Oeb
dKdidrWvADIimanfZ3Ua8+JBWzWD3pqjPFbzKgP4InM4qmGRk6VmbqZ5wPVZ46Yj
k1T3eKQcEg/FCAUYEG6BPnHGqQc0ySnIv6f31XU594hHs6Luvd7+m81zvHViLiFa
IJZ30j8f4ootfxglsRtP1A==
`protect END_PROTECTED
