`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47vPOHP75RcWYw+X8bNe+Lq3YieNFAlazZ/RneLtWcoW
KNRy5X8c97lfyKioMREEw7KYPmf4wkg14DWP6iV6MJsbVO5mHW2fPbbnCQwUM1vV
gMFHoTV01f9ZKNA+h9TVQRZe5/Aorn+Lj6XcL/G6V4byClHx45hIswBh7NBh8k1m
Wgc/Xf602zXSGqJcYOtH+hJ4+41V9DdJ0StBHXQ+yXO/Nj7wdO8njBFeo314Raq9
cW8963rN2dZMKbSYLIV19mSzc23j3feWRvVRqt6f6Atb3aCONl6dnOuG9kem1yan
SI/7PE1BSVQsoXdlhuHlfg==
`protect END_PROTECTED
