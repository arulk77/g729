`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMo10pOCTs4uEp1cUJs6sDSdtmKhJNm75ppn/ax2wBLM
DTcIKYaqDYF7Uv2OGrmsDGw+kGAcqFvnNBz1y1jDNJumNl2m5lIxCQBokdArDf7+
5h2xjAKmQpJRFgLkO/LnHTomC0tj7zyD63B/zKRzOUckcCquuiQn/oWMcsGbKDYc
`protect END_PROTECTED
