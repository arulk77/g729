`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C4VqMcwWoYYRe7jUjKen+D2l1HzunkAaU7VuEd0QSo04
tleSqqBVDQa55j340D13zzLr7lHrSFtKoHPktNpiXI/WQBdORrbp54tQrtdA69kq
quKoDwQAEHzQh1vvyvjhrfw9wWU4DywJO2ipgsqeBwvSQh+JyVFZF0BEOnOjz1w/
w5zkOQVRFHxd7OPZ+72sCyOp9xj93U4rqz0NCnjUDqIlZ+s8oW4ggWn5W9p4xGan
o7TkpyyZl/baZPalpn+qqA0XFdYvEEAlpoXY09siCcKyCo9axJsMMsCAs15M9ebM
q32axqsM+J6jy7MBd60q2Rzf742Ei0eZwmTIroN391H8QoizXGHuK4fYRg5VUn2F
QD4velR7prMYQQ1TuT7CTAlv5Rlb53reV63F040h/s6o/EYAaiBYq+eZgf6lKIFK
5M/OSyj+DU0JjxvclYYIw5fajQfqDD3nZQ5NwQ6ZL+sN3j1xiDCjIQgpkt+QJWaD
YaW+GSq8n7D89aUdsnhBT7Q3uCtEv1ce8dwhD2M+D5vp2+wF7L8/JYAAhNtxWjr7
x3ygZ04f9JCoCzQPayFhsKpOAm5x7B88HuoFVYmnQmb7S1q9H6lUL9YQAV5Mv0lZ
mLb8SV5nBseLV6eAhjQTA/sJ6kT37qVnWB67De+PnPSa7zOuvepMpZawmSKEvOJ8
W64Gd0XcpGAu7/6qzOtwb2q6t7mfPEwaEug+AeAKHVxvLKyqkp/pFf3GYsBjNw5B
wceO71L+pT6bLBjvD+gZQ+gIlnjL31OPbD9rP+48+Wxtd9nmuTYl8AuS359VcV9M
m3+aoZWtS3G97wy0/Kuw4HWcvHC9Yf3ScauLQXFU2VNc3snQl6eewsVhQ9rQH4OD
7u04XB6m9o72z+/+oEG5dK0h3KvJVr/v4NKtV4HFJW7ZHfo7W5pu9PpYi/hHIY3G
YhTZA0JFPBiBAtbHtaE42T0ToUnI4gtigsD57LHg56yz+R9NjbOjMYD7kPaIfD0/
Qzv1VjhyeiKgiHF/G2TaW895a5/xCWUZmDwF+DYyQ08XBknuqEmBJhq+nkzVvsTk
OoQxz498hcmob5EZpr4Z5G2OGXuGdsvRwUapD/IKzc6p0+/CIMf2gBmgsteS/XJM
8kIzUJb9zln06M15m3746QRa4uTneoM4vTyqj6Lc1UtvhgqiiMgek06NF9u8eX7A
EhuZMTTXmtLPFVCatE35kVJB5Y4TwVDTuDUOP+R9BHkT4CmIc7X8K0cAGhRK1X1u
pDF4I43rDU+uXkm8YEk4sMjszDY1+YIo0gNzIf4lJF03FP622KzK3hlQ+mjePPys
yiH3RQsBkOoMXnrj6f08zS/zx9vXHhnutnX3hwL0PU3arS0dw6M2GlGM7RBR8r5B
/BH6HTJzgvq7GCaXGqZEvCrNz9dSsXgPb4WL6c6MgTL3erXTgrNDfO7XF8VHIHKw
O2NwjpSiht6WNuuk54i26g88OYTPv7sTfKTYNoEapJJDjcav9dnMXstYpd9kdq2O
Mr97sjedX0RfYhFoKN4c66oVXLcqH1rYYCTkLyVt+Fuplg88GqhRlEoE1om/uSUF
SWc+GbLDotaQ87L4mRzh9zHGyOHlroKiEeRQwao+Xdh/cxbA12L4iRSZ4m1fJdGF
1snQ3wXIy9VXZ+LBWXmWKlUC3Z+S51uE5fXRjSPA0eUZQlQaOM2OkOAnQB4ek+qz
dLLWTniRdo8Uk6PbaH9reo/9izowhU/1hAdydEJPWntgfUi/f5PSPY30m4fPSEa/
7pWqoL9uHjZHOI1qyz7qpc6squvUx8TiKYoWXsPmT3m32lP4pAKan3k37GZYfTAK
Q07dxoV4v/r9BZNzVLRJLcK6pIYvhLiSBxXz9gFqILQf9kokJvkIrL7rVbfR+2JR
dtwbAxSJyoEDHhnvEOiUISJSFlTEwcGG0tFRkCw7hcJfVcAl+5vjZ2iLzmkV0QKm
EprYGkIP1WT8vaHzL8DLnToZXt83pyOML0AaGLcaXslVv4CNx/HaoSh1tTMH2Q8R
1ImmSFvXfyr2Sw59LJI2kPvSBgz76WtxVhHS5LWgLKsnIs8BZQsqelq5UjNnSTOe
fC36pePv7MV4feBYR5s2h78H/ugHruJ6beDMcrHYrVO3IGeLT0TbzMp1g5QhRC6p
Miu3PsVT5bqI/PF8l2LnNaNqXj4lCbEmHfZpCsbQGY+7qynx4kyzOHEbges2V8s0
vB9VeD7kBuqJ8YurlMlkIBHiuBNsrcJfHLp/QkwtTF7QLITMlXlFGYR0IH3ojBer
KT1Y7DQI6L0YXvX7MNHsaBmi2qegomr52jKgx8EXm1NlPClZ7KLNeMPnZgvjAmH9
u6K0W30VvIqOVDrSWmzYcu5KDaiS+SUL/eUN67Z4GYx5ZZYZRsYnDBySPSW05zyB
ogvn+CWGHuKvMDmKrvaGfcyi7yb0+tu8S3AeeorCNPSNI5etHoLfBbniocwARXTn
UId0e2cdedcjvF0E8QLeErxprjMARxKdOxVMgFk5wFtRWMtOPwhNX2QIaStsRxwI
ADqe52lItu3rfAykAK0ouCP/IPFL7wjHL1Lxt2gnwKVWVcpbLjlBEny9qyfylBSg
fvMw0k2Pmp4kf2WcFGavbyLKbVLv/xuX7tJ2OzP2bUxElyLXMprgROl9eCLYm0qE
SExxR2FjyZTRZYS841dBnx1+Xuf6UwzOfa+nyzixVfbVvvDDWMbkbQMZcy86IMfu
NIu0Cn7wSHN9jK9+lQIJbJ85J3nW6UBRI9/8JtGyRBd34PMQPYYl0Pda+pcm4WCw
BnYLdH8Zl0A7dfyZHHdkIeqA6uKRrIp8M2jMEs9i4lbCQjJP9W0MD73yHZzQizTf
lNY5ME+snTWBkiK80iOHauT0nuzpEaj6CrU3gMChr2Gm4k2Q+OYoS363YL26Ok0z
m1CCSh0TmENo6ZEkg575RwJ8nmiJt274dtuXl2DMQrDff6iMISTbHuzrW/VF6Bzb
auRw2CvWWR0jSfl5q+6c2khLmeLl6x5QJWDFTB+C57Zx2JWQmrYFgNla5crouo0Y
KlIgbN4bYM+fXOBsYdeyOUarzSruKfcH7BWYGguW/oOvizwwJGb0v8vkqnLTq/wt
WvDZGApBoiEJJcbGQuT2lpudDjV/hHAUQpkLEzrkrpjpM3dwilCQtGoUTbTQor6S
4NoD02SBNOtwbUDFUp8MOA19Og7zqb/or8GSqjAjlFpWByq0YV7+McwZfbY/rpiA
s/oXQuv/jk6zhBIFZwKm5tnQU4LlQADEtK6/YWdpjhGQZwfxkPtT3m3JwQMrFe2U
`protect END_PROTECTED
