`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wT9tJ3h0x1u2iRGW3bZKXxJmmsB21gxdXfbibt7XGHY
07h1/jvznJmg9+ZWxT8C1KuwvKal4IF42cLTD08ZJo8bsmz2DB3miR/e63Oz9K7n
bm2B7gzUT7nFcIe5pJH5wR6rU16EaGGll+Axuq62inmdCffgZcZ1duE0+KQTn1eD
oqM8FHyhE1CDhlwPei7u7LXFEk9O93EFnAhYJY2kXWyVayJOkNIwm5RKpWuj7t7G
mfT/EgeBPdTPSYxAEg8DLllJddKYFRuQtUbiUQq0DjKvig8bJzBPOpOqvmG4pALP
YrI3z1bKpa9oPrg9XSbkepVAIRrQrCai7BOpB6isXesemOIYZW5Iyvmf1+wK02oZ
3ZN5Cod7rCvX1t9LBrzLtnHOsFynyLg14vO2Ghu+cY40IiHUPpmM5MUAwbsUoAG6
sGByEi6wVh+dOyJEYnehJQ==
`protect END_PROTECTED
