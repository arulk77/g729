`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBskW5X0ezGTuE+8DUjNXoKUxRIozdySBV1NqdD00/Kk
lOXe+p8vGcgnh5DI8Q9HeERTP+cnid9xcF5kAbJPudc+l/jrj7foa9LtwCZ/Ugub
SjEHRQxardSw9+qjyY3Terg8OP90yzDvMYJu6RJTVQAQolwiAGt7doJpgnEkhSMF
g9BWYL4JkgLyFYnLpRBz/YVubb/r5ZPTbN8K1GENv+l4HJEgT57ogTIiRIjehHRq
czG2vrLgVQEBUoKlc02AUOd8Pj+z1DV8Qfxnv4PX5Wf5q+9sXB+uhp2DV82M05LZ
a2+T+qEyU6I/Qmmf4BhOSZ4PS+IJOxPoheKuNF+p7QAVZhrDdEcUqHmUGjjcCFT7
UZH4yrp/fCVMGMnxwtbrSCkkN8gIwgSLi6JKShWk6P70wxfi84KXW7l02LfKFdPk
6wo3Z218RVGMnimvs7Y8ZtCgVWv8YuvQUtKcN7VZjbbGavoKFxJGwdFmzdbmi7ce
+cdDNimjIJm2h94EiBH4rczJWj7QyMVwG45yQVSXhuBdR3Vl4zYjQwMZLWMTMZXB
/FCFpK4i6zzE+v91L4dY6L0Peq1eCRZYMr7UDLPceg2bo9qHPwHCZccS4Pu0ZwNg
RScofiaq8iO2VyJOdDVO3KUXaS7yQtmOaTbHuKbWgaMukb7z6wTxzyH878thBKsI
u5vh5iZv8qSXZutSmVX/oq3eEEmstzVjZa1OUImjwiZ7ya9s7NqKhZj17f0FYGZj
tqt60F5w7vO6ZUVsaFBCLLqRCWvdFf5mONog9kiwCMciqJtKoLZmiBAujbVLuoi+
UxnZmVCy94UaeLqOCouRhW0urD1XMVk/MUfSz/dF4+Qhf98PwkJeCkZDA8NcdYZy
mU7tWG9Bpj0q2IdCfQhxRIZbi+0m6hncPGJnprDw1So2IP3hJ2h1Ln+Y5ax7VkKO
/7NGHGGZKXzNsLspg2u51BDBcSosMlnYRHORMXLcFea9j3Ljp2HDoQeF3SfkWdmh
XbZJevx6Ur0g1qzdydnwV9yXQr8LxmATs1sow/vw/y/9SxhS4enfe22FBtOHdLxB
ufZ5aCK1qXPBdX1W1jkUAsXOXu34PbFAMHNQZv/gS/c8b40qzDRRTJsmZ7f6DpBc
e4Fl2OGNxXI8j3jn0WDr5hGiHYDwARORGvP3hZu/U89CRvURibXuTXVo/Q7NGO5F
mqdwdVQ4nYvtUm52IhW2YaP1Cc9WD3RWx1zVzK82De2A2G/5S41Li+bysYKl/+Fk
7OI9QvxoDduBj6I8L0cWVwIPgjT2T/MX3siYqYZZkufikP9vfnHeO61pKvwN6deV
czVDlkLNM/DL4jHVt/1fPGjLQEzAdhLMRLdfGW7LxSGtAp54jRQitiuae0lSDGei
e2nTZ13i8VNi8vn0Izne8+2UpLVdpd5oFzwD7IS2ITkbUGhrkBK1O+OKJseX+K9g
36T/p2gLu5qW9n5ydjXrW1a6ddJUOKhuYrLn1ezJ6SfFdn1ZqrBAF26G5kDhmERE
Lamfjy7QnX41Z8CZwWUw1nZloNIYxI5mOHy7J5vupivsSNLE1OL59J/TCxgC7+5e
NeKqj6OSEfvNA97varc5PG8T0+SqARyw2v+5iBD5KJI5P469CsQ3JVIXfSfuCjO3
Vj5SBjL3BVcZy04ZlvzgR461lHVM1jcmzod/33mwyNjn5URF9hWq/bpY/XAb6fvV
jbCoWS6nCH6KQ9lB9AgERVe7lWlqx3Mc05hS2OAyqoZ95EefsjfcZxAhBwOKsSnh
lLlZj4ApnfWf4mfBV600hzyYkhauMvMqQvVAD7cZnxmtF6cebAR11nsQmE91S9Xf
n/fTqpUQmBJ7a/TxlJQo8DGVftgZpZf68Zj+R0BbJUZaDFyO1SJsCdfXcuhIpZgf
mOKvjw5CMZ1PpSNwKyqWI8FbwaBi6hRP0fWRsuc5T8Z3QtvuKPZwHpOt94NxDhII
oyqeohzGFDwf3QsoVjoddLxYeKOWCnJIokinDynD3o8RtUYRhRRbbiM3CoELuVvt
Q4tPrf5mEuYFky+TB+uRbVtebEcl8e2/YaDGX6SIUb+iFCAIb7XkvFabdreR/g6z
2A92HRhLFS2ixOJi4B/cd968a/1JAzEU3xhrSiKn8W1+VOKuueLI0xvjoM3Huuxb
OKdEJR53tBGzNSgLi4hvJrrL38RBZo0/JU69Vl/8lHuQmsxY0aUdR8mlXmbJmJOD
aMummo42G9POrU5CS4BKlnJrxi/5awDOM6Atn6+rjb7bFkESp5IU/KsVp4mUHL55
7mevw6cA+qOINq9IuusqznI5PkPx4QyKxlNFutGia6vJyOrxrPZ8YoQyotvM15ZY
8xIcZYOUnQmiTsWk32RkKuyOteIJs1BuMxZi9s4d/sUVc9/sJ+GdC+UCVUdID2vM
Z0Mz69x1FrA7ASwppW1nO1brg6Ksr2kUawzq9sBgYFEsoUJe17X+84XV4HwX+SfE
bSHxrCwiH3Dbv0+rXowSFLQuKdrzpzv5xXqBM+HnBWt3lx0UqflspEcjdf6iKe1C
VA4REDTIrIeaywz3RnpSwr1+bVRf6V+M8Ee5o1m1wN3rv0TkjuTJbHoJSC+YGhFc
201sk/Y0kwbuF2oThfam1ebwiv6H/iPJhG93b3q90emIESXtzl6vwM9+DrpbYoTh
RkrveuwRcbdBfo/ReTavK1quolxMM5voo9pZ2ITJM5tA5LocXLEJ5VUajptDUoPk
hwZIsvVcRRMIJZrXaKYPd37OTH8czuQ/OETUY4JmHyxV+Fwfv+AHypfOgwiR6Yfm
Sd4VZWdl+KCbdD8AL+FEc2g7JlHbkz3x/W0ImhZ0w7jS5QgVBjnnEPG/nni/6Nh0
EZHQNvacF+VjZYrEtn1G/ZCPURCOdPsKJxWFZPZpXj+sk20Ou1oi2kZXs50hh5eJ
WrOV/eGOO/8HCpvEgXXxZz5WHdtnYVM38rQe1+FccEfQv5Ji+kBTu+wFJNRzvKbD
nqSvPu/3Rp5QnyX8TLtMfsWkCCgqLpA7/FDp8Mi0MhRV26jJ8mCmZ7L3iTBnNNWj
8GNirLJSz8RtBpn+5e88x3uSh8+v5EuQ62OMEHFhwZacFCExheFNhrVnRei49O0K
v58lMAJJGhdZpEwJBg2pAzlCsRQHD/YkTKObt8S9gq0vQU6c+bIcFpJxSRHAKFhI
Csjv1muUZR+XZsc5Ru40ZLprsGztKltve23sk91vnVsVwzafl81579F1FumMvkrr
+2YrWOY6ivkiWO1xRg5btPDciuK7tRUMySOR2GxVuWle08dxDfK3zwdto6Zxh2l5
4qLPJvRxAnROyU45fw4MmuapCYBod5QY42XHVckE/1naKhCWNVHRZIElmACt5CW5
lrdzaBAqCCoKr73JP1WhpwDnbf+onOltv2FiXznNzc+kFmc1YH7pU7I2+M5Hc4+R
/cBAeloWN/4JzGyyBHSc8EsYCQZZz9cowst7fjqfQnjLdTZpU8xoYez5ExT/mQOU
Os4u98IPBclFy9O9f8FhYfL0LdhmcbE9PEPgfVS0VsuxKpgJuTMntUDbqr5wCwWV
3d+UISCmeWkmnJBasBvL8+c8SIdykf7uMfdS2oqXxxDFfrC0janqAZMg3xjmAXuz
IoQKVkStdh6RSMOE1wr8SYnIUBxe25rKVeg6mfIJWTxhYUKl6/pJFXAYNxo9TIL9
ttz4DVM8De3+KhKKxTdhC6M13QaRBEUr+FyBeb8HTp/st9z0pzdK7qFTrJVUrcBZ
3TPlbD9PRgO/H9bKJ6DL7VgKSbd4MK2Ep7URwALtuB2xg3iOnRcVONAchW2doY2f
jbVVk4h6SveG4vUCzDZkU+XFuApBfye8OnyS73gk8wyJq8N8+44XNYjFCDQJHo3c
AldeoUAyDzHVmcybXJne2tcPA1MAGlL8ENQx7971r1dGSm73BUiRbFya1pRJ8WAY
itPiTvi6nmVnqXNiT0XyUoIR3vC+s+PH+ZTyzYXv2dEv7jnn8FlVDcjD+YCORlMy
TjB3BJnX1aIt7OTjxhrUulHaOGRb+9ycDsJLICYbeUuGmgyTLVLMC2BcQeUzA+z2
mNnN4f+qWuQpViofcnQIYf+vd6wzOH6k9uAuO/CiuWwMtujl5DuTL8B+FZx280ae
/VhTyF+C/yaydoEvdA6DWbkaa7ZDSKAbVqYn8KsTEB2D831TGdLvNQ5yswtdCGWX
UHnuCur0z46gBkjxA19Wgycn2qIMjMb5VXBMQ6+xiV4Rnp6b9Sbf4f/TkT2h6w6z
xUzFgwTDWes/d+X4b7qpxszHfYP+pgTZFUus1rlQEkTY2hgMpLJhoZ+p5v7JFlKj
+/nXulJURQxfjeJ7VUINUnGp/uY0jqb6DKh42mx3G3QZ6VKqoD3XeW8chM5J57QI
76/qWZyul+ZTOmEL+QTY4Cg9N8QPa1pb+1+6rWVWP+v23XJyKdGWqvhNLZe3zUYW
wIo1pFY+5lmNrdq72mhxaSmId/HMUh2Wntejm4xsLU1vmgf7AsD3YM/mv47RqEFc
wtkK02NAUUxBHcSY2KKgxNt+OXSK0IJylXt2WSd+CiMad+J2h9ltzWOxs2W1rp/Q
nkt4D5GCthR1fgWxRbVUVifxwyeQyMly+p4SmoAloJKdyL8wUUqvPGa5uwNank34
4lXdAHJZjKScLH4eTrC7MWqvKOzLxGowXjZ/4nxWoxzcCwNrvgBlnlz/T7ovbXNv
xDNtIYkFY6tgYb6dh2FoWDDowMAO5NTDrenP4BDv//nPyRV84QQ8KTasQH9nS0oa
932ovPAt44iRwzT4H+meyLZviwyUs4dFkfYwyvP7hS4+k1d11zIsAKPMWWwcJYfT
A3hnozHlojaTiRD2pKlFHHK9+BJRSlWzMWDkA/hBdhRE+EmonljErHiF9crqMQWm
Y2/vRr6rz+UsAwbdJItJEjn0pMkPUflYfvxDzpCFt+DugmFcqljKkG+AjbGV8k/7
9kvcVnetcfJ0H14yhMxv7EWnJgq3nqAJHVBdhg2Sb0//DAYBq42Qbx72ytM+DS5m
LH5tq4PZfZezdiYZrJ10pfp25X+3hLiYBg8YvxubPE8uCs4OjoqECtgYfT0LNbAY
+Mesoj5H8s4V1sQ7eSxRPaaHZNO12bRISuLFV9ct+g0AtltGMqrE38I5FreJbyVx
lOlA+cvkGJ6ZPaN20j7oIOvR9wRypShZNm4t7BJEu3Iel6KNAFtOicaz9HDyj3s1
ych56juZrV0s8LBD5sbdNNPGBUAACQBA7gljddeHe8FIGrrC5uwBrxyTipdFhAF3
+UC+lUPStJhddHYzLsMQ0ozfDxHb8SZxJcpK6Cnqothw9yhjL1UpBHevorwMUZKV
S2OQv+Wl1SOg8hJulAKwg9Uui0E3+QJWmHL4UsqQQ3ApUFSfKRpvSN2eXjbr2VMt
P9vJzXi1zEVorRVSJOG3tUjovo39ufYAcYOCbZ3qipmr15Tzx6GgOove7/4gDVZ/
/O4fTfFpRPKI278t9P2cgFkfv0ocStf5Sqkh3DWbYizQ3fHEQDqhQrOxOq3SnAGG
rdoniV4Se2nIA5ojSAmltePZoVFgD/SkoeM6g0/uRtAXmfEC9o53hZ6Yw61ZzkBa
Z/yldlWVKX8SDZ9JpH+mFsM9scjeRu6fSNTozpMPlSauosGYFSJ4uGSPh3cjGFoQ
2zraT7deEBksrLwt75pzi1TMfq2ywppGYgj+qi5orrKWvsZ4WOV/+hSZ7vVHZz7Z
fioTp1+a3JfZhGJKmyVfUYloKZ+btME1/IwBXiOk0p6Iii9M6bbKEtHgIKLJ5rCb
pXXExHIdLRpdH0uaZ78hQ0eKxjdFPdICdBYw0bLhD26WftWi7RhzXy9sTfcXdGQT
OKXXhkMDGuxC0eYTlclDQSSGP+HXhmCkdkmSYImf9VqVp67ciUTzCRL6Y+fRemhA
nVwP5UdVvghJ0MmvSyuT0i8HImYF/ADNiFSpBQ6krr3lxF0hkw7vIr1JSgg0e1X6
9KUXiQ7Kz61IS8Pl/XObTZbNDaJs8j8UkicRIdEb/moEq75A8cJ4R0/amWMadqyf
yCTGnRdVfsO0ZDRwpx/1cUWVksuPRntzGvcTWqp7k06O+zYEQMMLjeKTsIb1hpr1
NY+VtB/vDC8Q9qBeOQd/w2+6KoIPqfrFk4VcsJMSZGon7E+TYy2BQ0g0fcNlLjIs
1Icogquks8SL03js6ikL1hsn5HsPd0cBmmGJZbOxLdheVIStcC009H5KD+HrnLbm
MM2gvU2/E/L5jUepWkdrSrSMx8FQK6VouZTKF0CTY6geHVjekaz3FnITxN4N1fGZ
rd60K1E4jqvkhAMBRNRRMvSMIxOvGT22D/KI0D1+HZXPRL7ywcwFWXUUQ5suZivL
2ua5UQDRU9Ij6hSVpjFmvnXof46r9qSZvZIROwGLsNtbVpTVdAS8r6Gvbuy7kiFE
hFxd+plHquF9CfCD7i3wIF8dU4248W85Xry7N8sinLwH1MUXUc3W8w56C+oLav5e
4NR5jD7rPOpfQWE8PZ6d5i27knqih1qQ6XYX0Dh3km6vslXqap3o2nZiQVWFl4ZH
CJqlasMp+hbNWpjlzHdU/N1lCzuQBQTkwGCWbBlMP82M53NtY9Hn6t/B5ZIFIUDq
xdkMvDOFJrOp0XWny+eswQTkhobVFU08uMSeRo0Uv0838sCUNfzfh0JttFv0Bhmz
tunh7ZJzJruCdG2ILrQVBvpxwezpJwnSdlL99i/YuBRMNDRxrg4MyjBpuBbO8se/
SMPfozDWGUYN+3NHO1f1/nI6Za1SdH4fkZtM8S13n1obgTuVoe+MW7Ew7zqc04ib
EsxML0TG+2+UUQ+6Ckmh4V/6TW3r+ynnpfe3aERc77SdSc06AKaanNWL0tu/lxpz
ZmeNMfPnVJGL6sPMfjiT3QST6K36OjWwbP97mzS96J9Rgrw9F/nBjROLngDlYnVy
YlSAnbughw0fKZ7ponBJYG0r1eIsMcSbKebeWl5E5DZgRJDQbuqw/xh6oZaZAAyf
RQkfHKKMrDus7E6b49QkEcuM0hmb+KNDF7dYwQ+VodyWHZqyyH+oVUakh5fGlRKj
cQUNtjHnVWFk6hZ+LtYhD0O5RIeCCnDwQD0rDnajglm4VfB/L3aUetv03Ulm/eok
RtzYzDFBCJaNah7iM5e77ORD8SQ4LmoHk2Ud9HkGszREYobAPwswEWGpOF2GqSqf
E9XllceGw4dHeOcuGryIyx/IL5yh51IMW9YzumUubl7vExmeLMtpJd5OWGz9v0YL
MXL5yZ4Ru8kSOzPqC6/qWz1VKtKGHo7BqN/Ap83C12N9LJXLWnzOKYvKNVHoVNiH
Mgzu99AJworH/LP2W64w55NMpQ20z/X0D6DSHlMbnUtL3vArktD5PmA/U+GmgaVw
N/yamexqZnsYz3oAmuFcXjPeWDMW0+WuVzX6JxFgEqfklsibH3IF+/rO3Y8EEXkx
jdqSvS0DIQYjLhkZJtKOwbzoiba8Svn1NpQs7CDm9NDJhiI7wdAhPDIHE9c2hHYP
7uAXoreFhSXfQTg/e8Wy3ALQjrGpr9XMtb765fEXgdLgGqmqZg38w/T88G5l+rM5
gHhilSJf7eYChl0CHef8LHA1eM1jfXCaQHWNhH+VRbhrjKD4s7ZWoGsvrkRFdk72
SDODRz6XS2c/3zCYZOxnKZSy7OckBcXXnbV7jNlsYuVTpqBGrpIJvqNnJcm5Mzk4
kQS+QUW/f0h2AB0ukUYY2F8x+mSTKyONb14Ja4pS587n0sfrlEyl7fp7JBbyukdm
8aYTUQtn5HfvvkM+U6H3fc5Euw8RItZlYlgDPvVFWYAxfWJgvHRaU+XR0usRixGf
Yu1KB8WUH6tK/Ey4qCUGaBvXIujgjXf6PZAt2SUvotkOrtLY6DclNKSvWWTPYzzk
2zv16vHEE/8Ea0K3yOYGsu03cMheuXZiYKrytKqnJm85KQraQYxPM+UOHxY9D2Vj
eoZMfqtDNUX7dPHwwSBmFLMB/M1JE5QqnDv8Ha4aNARIrDHbIe9fknYo9mq6M00K
8SiGEoRBaj8lzyaGpcYQ3iQ18XgBFtt9hTIgY/HI7Q/hLAJtVpdx5XFLZxZ0+C9+
iqRSCZYj0iAFoTulrd4A2eNNKR7Eh+yAbzNhfZLrjR+YJ9yKXl/+n0uQOuN6jdg9
Nc1Pf2NzZUgg4NUq6uQ1vEPWbabTBjtw7tnGgsfNJ/CxFi8elg6p1OWBTraf5Bek
svVYkK+ZwUZTCTuUu+G8Zye2V3mzPseBsjkolpo8S26FVBVAw/T+jSf0GgS3mJKi
Ftp0gaMQ8Ww5IEc9/7HoVqa9TqYBSvgCIkVdtC7Y91mMvt/Lx/aXS/4wasUJpCwK
iHS1hq1uF0JIYz5uMSM/qaSwtBOsV5kpjhBvu/dcy4aQiS6g5tWGrrH9HEFQfxEB
fpOQnTlk0IK/SMOS9jrXItJwDpRlw5oCRDB/E8a4ZoxxvsYURKue+/uXFRGqSgo8
EzpW4VECqDJTCXeSrq77FvmxsczGGH5RlYKVxP09xXCeBuWwoZoyOftRlGPtOilL
rm+bZyqWBEL9Y/PfBrMbqegFohG4qY13kqqJjDlo4FCBTBe7PescNWImsgAyUro+
QPn6Sy2qjHyuJ+j35SAv1JdZmkmqCtoo0Mkk2XI6Q7zQ3auL/LhlVawtsUO+wWcH
e0goSz+LblOgCT22Lp5evVOobsnkufcRxHSWBVV4WHgtnBdcwsgy5yNeGmeI5uY1
N6p8WKjCPI7iF/epwNDZ3T+66J+oeLKfIP4fkvAM/O/Ij7Ofp62y3kFTAqdJxpn2
dnbtCR/V9S0uM4aMsvuqnOrOTKdhubMIBjgXdd5jw2cZAkEjgclSiQdzMhjDm+ug
SvlkyKLtZX8XkZ40ZJTQqQE+HNqaIlbJXUUQtIBXpRGkKo273DWTu6sqzHY0UAl6
+09ahREr4wpwqbw872BPFUEBhem2GuiW8Z+8EFkbqK6ORn/HsdhaftzOzQIzCnMr
ryx9frVDMUnZjFD4QbJ/NfJz2shf2u1Mk23wp3snr9reeh/b6ndz2NWHJwt3eurZ
Lz3JGXv7/s32FNLG87u2qs0AZVeKQxvmnE1P0JyCFyTZATKV2NBguAj45/nAp0Sp
F9uYBcMe6mBs3my07pcU9cWW8jMGUgQuQPa6Q3K3CLVPWng1Yppu0iMbhZHRBNwN
aSF76jZT9o1OjUfcnQdYaiH1djXT+CjumP0Qi6Rq8kRnPOx02UoTm1dRDzzS/stQ
2BO94m+IcRptbk16tnhtCoati0ZK7rCIznOCMQJu1wUnCdsgYnSuBdAbbhYhVe1t
LV4l0/oxsfn08g5G97NcQoGUYnr0NFELHXR5gh8E0GzgAihZDxjLlLHI2TvP7TBo
hP97Xoow8SZ3BGibhYxnuWGG0C4xknWQXvO4bObHzEvT4k+581W9hGGFuBqtTdxQ
NNa92kltMFHiIV9yhITiSyNz1TlUcbsPF/rQ86m4T6Vz2G8D3EvzzAm5QaM/bA4c
e3Q9G2gh+lK5y/2hhRj2bR6VLN5oXicpoaD0Gt2wMrVqjjRXuWb6AYPBt3ztxCpB
IqG5dlRXhfOxXF6ywHoizTisAGs0u9UWc9+q57maaAmBDqQrZWFHrmgUH82Td4/c
flIwXIEIaFMIrI7KW9i7eFeGZAvBaXHo8iItEn1TLOy6FPLyPjrr7FJaDw/Rv182
VRH86Se+9h245mnd3T7KtvpjtssKfH1np+FYFswJHNEcA5QCGX2s8BL785Nqpq3j
wnshuX9jzrirS0bnVsHV+rQ8yYAnvlhSweEa4Maw30143SivgDjxP7nAzg4V9CWn
nA/iL7+huL6xJdQ6bD1jeb4L51mv6jgyyVqPRA79M+oiCs1F3YI67HbEYH3mIY9x
kl9cOk+mX61mf7hlkbyi0XK8dXzCVnnmndoGvvfYFqw4/VBSi82pUaqDMQJPhePt
/Q9nvUP9oBIKUEAKbhVoL8Qo3C4ClyKnV/paAatem3hDqmwOBrEQYEoqQkYZmmkK
NctWWE5H6fKvi2M3xtEn2Lf/xTqpVZVc4qck9kwMUEx6c6rIcLhXyeojCR3xnR2s
+cV+3JJhx/7aOHJMdwvpO90EUTr98yf2NmqseL2cXhNwyTBX6FxNDFdse8aiBEZ/
wjBjAJebypZoR1OrZZVX5bRNb6StqG+07LYDLcX+DkROvAlmVnmBjRiJ42x26MmC
oT/QMCVfTfThbGZwEgKWEaiHIAz9xjkMHiV28UY8ERNwL/u0JU+RZMckKzb7Coz3
X138ADdHZnScFMHr9gkTHfFvRhP2P8+w2JpJeISR5kMi6aWuQoM9eeLohsvsFOPq
MCd54DWY8YzFh9te3rG5FYI+YfdEfGkOiHCwhLJFdOaWqgKcboMxYOZcQ0fjMWQR
7o5aYIyifrCHSBi3jdzq2M4+MP5lDNSPeDPPkGcZHXSkj/swfBhwhYOSmIf5NhX1
/y99vEHaOaiqPKPUjwn9DKK/llNDUzI9/TGH1tdYfFwsB/HXypqcxDLNW4bv+0mQ
TrQp6khXuTaiEhQa8Yxj+qds6HdTdDILhC3CKEnHJ67yyD5UeC/jcU23uml8xIfW
Yf+rnCJoOBkHIqSJ+yLcakP5Zbe4IoYgaicMeXpPHRz5Y4bRpimtdH4dkjYOiuTb
VD8hcRX7qJWsoSlHQKih4CMHesRG9NxbgHCmXUGnMnOhezDNup5oGkbjIDcgYKJe
jcaQYK60105L5pXa/5qAliScccJG0eZVU+SQO9XG9g1zXkaTsqPSfgPrgOdszvbE
1ZDrMl1zBgYVY25fO+IYcRcaTkHcV/0W3pScgSupi06fTkUZgpDcainQimTb0cTC
vfcMsa46dpTYuDsdepAR2MuWS4Xt+58HcAVy5HlM7HdOWb7R7OybIMAB3gRNeXHn
ZiV1wN2F+NclrFhFXstjHrPQ9jF3WIytMkpoudnhsV9ZVFBRzOhgiukVrnP/2xIs
oXOltj2f3G8C9W+X3+mixwGyqi/WeAe6QOM5jisSGOwmaHTws9zTOSwY8YF58rpJ
ExG57wRx77KaaHH/JB7SX5I24PoxqAoKihYGrwwIbtPj2feF5UeK+J8hTn88lsb+
/Zmf/45ukUik3JxNllPdVDlHLwR4ANLg+pBCw5x4EGt8OzNrI07/0W3Djqzf7Jyx
P0Svf60TiNRFAAGc5YNFu0pVkEZH+4p+elNj/7KELZ5c9V9Vu+jhz0OlKsA0OZa1
UrZngiZzJxmhMDhDEM0k9/wEqDQifIjv7ckSZs9gF47R7/dev86exbiscsDzsATm
wEoRHOXbzjzKvzVv5kIWe1vrXkR7tDRcVRpQCEAFVQ1VwTylbMydXOZeoZ5ayZjJ
NvxYGehz7+WHvzf4rBD5lGr7/gi7tnnveiuaPqmJbySEV1teDKvMTabIG6mRhX54
3Q85Y3Lj5FEKYRnLs62dzZY1A5FHpL+aiIbc1Sn8+Fo9eLJA/FrqbKn4rnhLF2ZG
RhHG1BhBrFZ8koZ8FAqYW/BbrGgJ03EQdXk24X9yDNKF1gsks++8xVqod/EQLuje
eXi0udOaATQxY7ufzg9UMv/6vTsnyGdh5kIqZiNQ7cmOUNtcC/8aYInC9XN+UytY
74VdJ7czd8+A0kPODfwcTrY/98JRtpPBX9lMKMn8qbNHPMC2a8B+LsXdLAAsb8Py
+TPeL5mbkJAU97Dy7jE9IqDCqR2LrZ1/JHNk/1Qz+b9gU7COReOsP8zK1RpjcYJ2
HIMihr0rHAhj141bdRFeEmhKuMdvJQKj7qKMhcmOoMIFXz+aKBZu983O+UdFx/6I
W1lcWZzvw8p04AQX3+pZoQaTIkWeW7qNB162cnvyMl7rmoLR8VxzQD608qU9IskN
Aa+3qEWGaGG3aO6MvBjD07U8lPFP1LHCTyvRGFBGiGxB0LvPh1OxQuebv83FO6Mu
zHCdHxv+cQDK7eeZL/8yeR6/ng7YNCTKW381Hf/9cHRHgq5T96LvexZNxPpm70Il
ZjY2n3niJE1WPTW2ClqAhGn1HizqyilpO23+7LUPm7rdpJiQUWUa0qZlgtCXnz1t
8o3UPmvyq7q83nzpKwL2J8u9xqAkKqr1+uW89wTDIeSH1B0A/ljZdas9dcfa1NMv
cOu19c9RAk+XU0lHn8/bGtyWGLVBJU5U9JQf6hefnP2W2UojDVwGt2vtOgwGM/nb
MNuylv0hIK5I7Kxtwgc6gxpazZzn3MuEDL0hDXONTNZJar00NEsatiblIMjTwSFX
Lw18wiNxOkqPYH61RHOc+7iciwkzi8uzRGWUUWZUvqFl4HshxoYOsv0UjNBeUz8V
WJGkMt4uhOit+xeqymT17St1SZCXpzbDUiR54HKf5FWNLslv3QngA/za3X5UwlJc
s8ExRj4ciUZfdscdnuAHJ9nbena846rUYY1Sd+H37aa5feYOB7twtqe9roS9vu8A
LRbnOVusfvdpyO2Tap6IuxBXZVErNfy44b/NqMiYo41uL97JBNw8ZMOHa6vz2+/8
fumr+QGX2PF8KKm5ce6CDb+marH3a8yNqEqveWE+U+ajk8nwZCB/C4WXQ4L2/LOl
exDSqjLAdUbauW8LXScsAs6pzPqmXMQ+8E5aPqyKkFYMVzA6Q4U5CPrkeXUJ+01u
qsMg/gArzQZuJW5wZodM9rKlCxlBYjgPYB83fjUgL+5/nYN1riHFnLEUY42Tsz/Q
l/S5Myl4OQGGwxi3utr/6Q4xvPCTVkcaIXfoYYUk9GP/+Sr3vikJvPL1nvVueRkU
SjkOWlyOtlYu9f0JAaH1rzGZJsjOI/UulZFML4ksHqLaub7Fhteiko/dBAPTILLo
9kQqhu/RuVyeQU1T+ATGo3TXCORei95TzNJmydLSwd9ipSsz5VwMlV2DYbwR1Orz
i8T3iTYlupHiHRPNzBO17yFpw/DvRarDEcqy/wL2fZjDDKfBZTb2AdQ+uJ54/u39
Qi5QXXr+QbNYurPSL2LM+PGi6n9hO1iWytmCZ4mhGFZjREC/GCjQLJK6ESni9m8I
jDCLDo7uhtp6pM9G+vhWd+8b2iQHb4OTE8B2CFP8HCiSgkfxaxZJW0Jh22Tgok9C
uSrX6oJJwpYxRG5BUZ5HdCprLonIlK0SEi16tK0ZlwOKhTnwkD2Cv6p5AZf4V2Xo
vX4US8IqUDsqfET7cYx3q9dHFJQcxxXDm5mz0SjuNPupFkxzN+/pF7c7Q3Lj1lvM
fRf+fgXrXk0zLPPFNRyaraSHMDl14z12kxOEJOimlbzlywCC8qNmA0YOOQsPb8OL
QgFi5nk8PJF9WGmVxAqC97ariIPE03n5Gp62zBBHp3/66pr98ORVWz5nE5QxIw0t
anoneF9bIa9vN8mnL/N1Dc/zA9fQOcHljBDcXsQH6iWjKScpaxFz4aW5m5XmfUzY
c4N5mtgXpsnA3HcKUQxK/Y2YA+vAWK5MUuOvJUQ5a5dKPAUCKQKc0IQZGTQTvKrF
aOHgFP75pBNSsOvZjg1pZ7It02nByI57NtBQoBhSiJR4EhwxfVOdJhBjJGN8yHxH
DqJY3wnyb0vz8O4BUyoDRAr05GENjXzdJ2SddsJKV0wMJY4zjkGhrAoaIpoZjKQe
fGrGXr1yXPxqFFiEvTRb8xWszroVZ1Uu5uoGngC3+8EYgaQ0MQWQUFBH18JJutiF
4MP3W7qoz9kl66q+470OfnH3U9E+dGMerwXSfK9VYnxuQGlbg2EAZEo4bTPjdycW
6bWeWLzp43fyy60flfWvAMr6UOkCTHGTqhDCTN0x8cweLfUGA2qZL6M6TVoyXcHs
qorHeSd3sFfq6Ng8pQ+9bIAU1X7G86fWbwFAYJ/fJp3FQ79UnyAtaizAZzlY0aY7
8K42bwTM5vFRHcvsGapqrZC/LKEsczqcYXDAeYskba+HOu+loEMaBtjabAO/+vBP
VbTZu7cAIaeeN7CYpZrGdia/XuV4H/7aWxtxZVBkX3yTLfe01Jl/5Km8PDbRdSOC
zkzyb5tDny7MgRPHgZK20SvXuq4Lnu8irn0Jcrh2BA1cQ45K6wXCWIRNBPTN/Lup
mZZ0bZtUjug3V8Bpk1q9kXYt4h0dH8Hi2qdl3veQ4aJAUihRmgdJK5e5KC3KSiQC
CSL5UtTSUagHxW+ioaCZNGuQi9hlVuXhaN6vwPjUtYksrtf3WmJogiUKNG7LNiyN
mffBfcTxnl4Hn5qWij2Jq/bExHQ1TEAKijSp3ev4dr8dzxINNwfx3oxkQ+1ZNr9L
z6ET8P5rCs/jzAWT3hqjFADw4oPdtBFi7EHWzG6nacjy1a47lJVmAN2v5fJtzdNt
AWg5+jhPvsGAKvGJ00MHO3PoOMBovaBAq0ovrYUGq36PYa3xvL7ADQiuFT0+Jx9p
lv3y+x7FqvgtY1Ds5/TlwaH3clL8pFmCeBAKB9hN2OhfoYF6uS1cTxb0fNYbjrH8
kPGzliYNro1oJZddJjwfMOVA9YvtxYmkWOaj6tNaC42O5Kzv0DoRSNh3bu+kh/Qq
PuOu30Z/SJNzynfAOzb2/a6bJtFDpEMKFM4oHjTjBLq7t7DO40TABJdRchAMBT9Y
SrM3lMJF5nnGhORgpPxG1ZemhjoCHAY7hbXXa/9eGieDRBjGXXBW24nsMsexb73m
Z9z3ZKVZHhJXFAvPl4dFCZpoiY8WjdYeo8r5rbFpuTZKFiO/8qJoG+GocwjaUPEh
iFH2Co9GsbsdEo1B2ZoTGSICkfkd+dwfb9ajWC9um0SE3xDF3mHd73d/Geqc8FDK
fYNsQWqCW4js20bhH5+JgYB/KOGSO2n+QsFr9V4/1l4hOSGX2aZDTNR6Naf2rPQb
NRs8UC0nZELYS6pOW1Nj+KvRU7LKmRedhvRgNWAk9WHKsKCYw8mA4znj0RvUZAw7
9L5Y7Ug7Z2/JIPwwGZBe8Dx4Wx00BTpQmCU/LxX5G+d6Nzxw0dsscTtW4OrWPZ5H
RwT85HLkte6JCPXow7giIccL22xNau36Ye0BOZdaao/P8o5KVyBfx4cfhBMeZE86
d14Y1OqapHQEvszg6z6+Vh6xJODxkv0v8/aCSyUHueBCE6IyeCWes/q+rp56gqKr
Y3t1j5FpDwGGlzNyNq4D+hQN35KFy9DDSe64jEoEXtAgKAETpbtihUqpbqI3prOE
/tq7+v6yXHSfU1DpNL/5cMmVKbFomtXmLRE0RdOlcVAzJMzONeW1hYe4l7GqP2wS
+4qviSyZPqZ8R1U/oAVKLphKEGtX6xpf488T0w4f7mioU3f/oqITZTbQ4ta0xEHw
P6VEfwtdHI3Ncmem6N8kx1yX2M1IJbBKjTKsn5pJC0QRYZYHRpEz0TXY5z/KHKrS
hP9Mpp/wbCprbVT2wh8YKcBTi4NlvFaAHRIjqGylzo2sEWI7I9k2x1jYe32tYUV3
XCtA/1o5+poRbiwiiFQseYyJ2ph60r7muCaVUCbRRpy51QlAW2JTOl55kQfFpMtp
vI1oTjgtCXwhRzVNyo7HOv6NfjdLhDVQYZMz1e80Xv1cEDY9+dzL0iJKcpkRrjhE
KQjaai9Da09CMLUOys8FTqVZEduK1B66fGS7eqd2Huj3lal89uKMoWng3juRkImb
MoQxdcbaHF/9arClU647kAhRx5tWkk/GpmHvh/1Pm/DHSABXN1qNRAmwo8pq2gas
cz2j58XWNNxhNKm2WWOC38IH5HwHnBcAf4YF5UDbSBp4WVQUr0BB0eJ8pho+baV8
El9OSYiaNNxblqZ+rq3ppKUoC7f3Crq2YiLznqEGdLMwQN4QVXpGJvQXjbwtC2ER
rmedO2+Tx68PzXc8Tb37ogTbJoLaHYlBE/c07os0qZ2z1XWJPGQgOfYJ1QHR2536
c0/51lpE4j2bF50unbrY13rwgLy6jfnp87DHAwXmRqkX6ba/9pdmjckMJ+jr+Ky1
tHXDVN8yRabYOVc+7Ke1pKr2ju5NXhZCvd5GcaG1HUOffTe3eNi4lwLKqKxjf0Z0
nLVdx+0HNs7lGw9IdH0L1tutSkw6lNaijkexMqadZW66SKORBgdOAfC5Kt/UrPrr
SM6aod+Nbsj3mhBx/f1CgiaBWkwFBJmzKnyK5jDVAMW7TD0Q0tdPVGHhVYK0VliD
NwyWLB0H/If/IdQ+DhmGXrGzA5kb1IpWxO0nrnjABcPiW3KMamBK986XyawMDSDm
ot6c+nJdu8/73bflr5MfhJHQRamxRUQ6vfmtcOFtBnKk0uWvADAxjVaWWMK4ulQN
1yuvf6arj9XBbuGxv8nw7+xm4A9128WpKQS6rrDSGlWyBSqgaO1f+xRZmkYbSkKV
S2Z9kQUyPd6n9xqa2sXdqPGpW8Gp2dCFSIlolUByJgM1YjCL2UeI4ZelpvbyLeek
Sayi5R+K1URfOWLmAg644l7GcXqxjr47KwC3q+FFnCsMveFM9QsrAEowbUnUJpWS
2PkJvbnXlc4Cz3V8fCpn6G+J8/L91DfHev6zK/cMLz1bGjuG0rcfUjBB+7RkeUdd
52/PTbh46oTiw0ClOBI85fn97Q3BuhDMvMMy5HaSlqvbju8jyGRoc0fSrhViek3b
LIU5gii+Ll3TUNAK7LGJ3fkswrVtU8+Z/awdq7Zv+EQKdcAVANTrkarSFDPLMqEY
eq94Dhp8TaKbZt5pE5aZfLOCAuQdSl2BhulEBuVIl5BewaEYpCamrhMdLs9OfjSf
GphbMAnoI7ylaftMDvWh154Ti+pwTYSVDr0mR/hInT4U61KQsMehyQLnwRZliimh
djwlGkktacSpihFA02tpm8h1ZFF+8yBRrSlCTNKQzOU2/0dOfaza4OModCYcxWpk
y95Px6dDBayob1myxs4+/kulU5mxI5J6YaFjLq9AHazZAgAAAw9eYKPw4A+TI9t0
uRJe5G9MZT02jZVUKMEHIx6jNQRGrl61mt+x1A2SafRbvsZJPg2cAEeJqj0lPHQp
n6OSZok4qTRvFn1dIw1mO0ILW759n5BGIy5qbWX6QcGS/0jToIm9m2lJVWTBYARS
mejBuBq1jMoUIJgNomaQPiSfBmeRRHTWRxaGKS7ZkKFq67PasuGmqr6mN50Id6Xr
uO33zRBFwBRmaFjXxp3jAiUAVMlofAtdBu2ThAvAjElM2Yf3yJYeXnVevspakzR5
sQ6TL+rbTXVPVO5ucs6x+we0hxRZtva6Vz1yDlGSk27+ny1unajl30hT/Wq0R3Cg
j7gd4hi7uBMyrhSTQ3yhdbfYoTT2PbWVfMGKSBTjNzyhdkwWQlVlObfBpoXpN9qm
ewO+ucBwYPhWfwiNFiGP44CDJK7LsID4aNTnMGyAPbCMMamJEdwh6Izhx1LUvU03
Mn5VOAlu6E18TE8IHE/aGZN02A0caxoh691J5nUyU1BD0dso+heIEX03HymCG7n3
cMmljh+CewbmDTHbGmSgOIn4EXhpzvuAnft8MGFWR+3i9EUgvSKwd2BMPds2HOSh
6jlFScu1WIqRCp8FDNcLoNCZGk97PLvaHHmG4puoYdm3FMBEKxIaFdGX1w3vZXJi
GVh0ix15Sfo3TQeNzbIS2O84N6nvvrXyYXaqQZ1MV5TvHPaZsfHSqPRZFdAO0jFz
y/iGtBJxta2J5M+OuD79WVgV1ihb0ZiwFTpfYAz1dGF/2lGnW/vY3+h6430DnXrM
vjCCz12HNVWgxJ5qGcUVGTZEXjmE6wnL9s4l1V4+IITWYrUIpPq381UW0uZJWnZm
aVhWIoh+7j5o5QGJp86LYJsWW4DQFOMwcymNDvUpiZDGXR8qpTWULR1dxEx8+Cu1
+bJ3ZEu0snX6XJSIBbIlaG2BmXsjXyUNqMTlaAVj06vFTluQm1D3VGfCp/G96o3p
TDqPyjphpLpbqEb+Nliv1exL4MbFkTDoaNnRUZO+fmoRyqm/GJNvF82sET6AXRaV
96KxJsWw8uqbSwG5uN/kRivC8PQRgVEKJZj2SVckAciI/KbrPJxbx29eCnBB/fxZ
o+H6mw97yyVMAOctp2Ws1TVWONcabRup9Tj2bvG0tLR/A1NTa1ED0nZNdcgkoxM+
3IFiBY8YCF3j4MwQJGwutHPCUuP7sq7mbzdEOjY+/zPyOmE42nejEA3YO5v7doTY
JSL0YRHANfhm1rE+/fUu0ETmEk2S0+fZbRuVDk6Cxw3J4YMCvuG/fQv/rxJ9TovZ
Imado3tYOpg6R7UeRYfO8iA2ShQmmIIUYC3WKkqZjeH8efeLm6o+Eptj25viLIg/
KCjNo1Q8Pyzp4c5NrmlbQe5YQa0VhM6E5pm/f+lHLm5JbWYspM4mnl0QVRK0+2L1
Y5JCCx2jTNkQwXL7Lt3flP23KE+hQ7uxCnwnjxRQafKyVSHBKyNf2YrwrXZkFDiu
kPrHOJImHNGZyQlVXqobHt03wSP2T/8ea1yzkicpVnizRR4YfdY9JP8AAjPYO1qr
OnLjZtzueZ/fLZnBtWDjAcjvMK9Nd7gbuZxDDM9mpoPD03AZxTOwQWggctFYO1/B
ah6s7qIKj4H+eq1vkjxYELCos/gjHoFmeKHx1B3LA3aLv/iQLzQk6h8xF0H+ce+r
WzzjSgEzRzfB/LVM5L97X138UL/PYDtBSsswndcmU612k1J8aETUIEob/MwXANm8
2nP266QnXhioAkBQN9C3kCij2MqORKpQzTIPsXaRxQYLLjb8BQEdYmwofoXXDdqS
GtlnklGcqDYXdc10PqbH/nQKJUFmalt+oJOsy8L/0TjrNMl/Baqz9bRL2y1NWRD3
p07aRceYtiKlRfD1qPNMjWPTrLYRaCMpAkHhye6FNz945l055HVaCXowzmIDOGik
MzffqD/k7awkHIV2TirXboFESNWmFtWfrjBkrcL1bDbMn9FVM03wDW3YG8PK/QoH
OVtvdf/veLP+9vglEPj5TySTi88aJK14eL3wYqeajn6Phi9KnTa+MPORGsTePIts
hJE2ioUdP4UJI7ismT3TKldWruhlrrxR8Zi3+Cv5USme6R4kwtWKRWQyrX34v3EP
QTa3lwiSANuYrmc3n/GdxfxUUyJBs4CTHCBSracr4kh77ISJU7qRTtzi1tu0YHdS
gliq9TVaTYlCb49JF8DdcXZJlRbDC/4Tl0F8xd/63da8NoLypvCnEnilRvgS+wu9
wpiSJmLnt/6JYY/xGBsXmGw/KfHOr7o+Lj8LUfugwIoCvOL2j7BjgI6I8374alLW
bwj4SeepPvXnA1f/KFrHdrGLJj73lqzoORLe/prHkiyk9h7V+2lvTO33kb3jAps/
2E8ELBJweJ0bo0p8XxiQSUFfYC/4iNsi+d83wnk/fath+ey3LyOHHrNJhEPCF/Xc
ZRJWdrcLBNsWk7hIyqjjFY+smNFgwJq+9WfIqe16qw5PbTR2Xioju09ZcAiqRhKe
I+CzuFTjLjK+q/hVxtROM47eHRxxkRRe86Dv3MfKRvQhjFrpeZkBg9x7z3LFq+iY
lK910F+zLoaDTiQaYThyH3Lz4/npFqyb2njK2/D22D0xGq8IV5gCanDH6FqpVm28
YUPGJpjBmfSSKPYjzcnbpjkVvjK5YHV3Jao417nbcA/cySOc2NyaqViWBNN1V/UO
MIU2bEV34avnddqJtlR10qgDXNQ1EYMAIQ5cjLO8SLuAr4TqnNBz2pHytdg76W9a
30dD/N1G2M4jX0zJGeFvtbVcJYLAk8T1TMEK5tU+y/U/Kpzi+LXoMNw5YVH70SPP
PlMipvN/CxofE0cmHcIQX3ik830qQ2zqyEt20OkyFqTqH9f+noKcpr73NxSDBJPe
9Ctoap1M3KkXiqI2JPOwQBRnsUViXXTz8wv0jn7cp/a9rR/AEmxpBKZZ7ta0Suzk
6XDCM1UIxRK359TlCEGTpqxGBj2rHuBkSUCGxIvBnWfU42v4RnY1D4DHe+OIfZzb
mBiIZ3jL/CCZ6RhPqB2f8OI8s0aD7QnndwYZnpxPpF35P6CHEf3mmKqNbU7IVLAf
xc0nA6RJXsO6+m4L89uwa2cAuM0z48U62WJLVlV8finYHJNL1B6FyogPtr0rDcXj
QThP/302zo7Gn1JvGMG5o9nizfThlRSIXhCqFdFY+8+IH3GzNdb2rP0OqUVKX0Pk
bCkr7uHeO0QQ637Jf0y2p4AiMZotsYSyjQUwONcOk3bA0xZ3Fe5x5lU4zbubg5sG
CYcuqYOwFE7zqfX4vxVlfmrKzpP763Gy1D+8TXjlyW8JT58z06Sd0gtk3J3iz0fG
jJCNXWr5RMmYnh1ux7+VZ7o/axP4soaoYRiggFHxyz5daZSVidnZGeN3ajdu8787
gt2Ot4vA1462Lijx9BkQdWtpJdW/rgz3KPy8TqiB268LgXY8F1yy6Mo2anPHWyk4
yYRGsN/9zTXiEH+5iktd/lowinv5WuD+qTYiZ7VhxhWBGLHNgPputFYajZtm016c
MmmUvQGdQZSTokZz8nzAIl7v7KCyBKmqrgOEUdaZ+UtXuAOnjumBuf7Ojn6oxi1k
Mdj521jUmfJtwzrhT+Zg8SYupK2gzbELstVYZi+tRZs0/kdHbrqdYwqwlpd+7Sk1
m3b3gnjpAYSOvhRMsSvg+HZBx++ckcKX7854B+YkqbUYtujV3cco4/sJZQg6SuLF
XQy/4Ev8OOByyceCgTF0ywvXbJCbsgQDe3NKjLWsz8kKC0fNTEuXGbCqPrzTvAMW
zpczgfgXw6oGgHGEiW4DZg5GrxzsFdrmnvtrcInNVQ7ar44nZ85NZEvO5B3PS7wz
4pHKxCI3nx/pIj8nYkX2N6ugnc5qOifvgpOBTytBKR+OxiF+vMsN8JLq7dW93KFy
dCDPn0KxkkWrax6orJlerMhnBJf9l7aIF9oFn8WCGgganQW2aelgW8hrLPKxMbLD
T3WGju1A75bnVPbrQAsWXoDN5AhRXSPiFXK3edAk9GabKnuCYtoGdWYsEXoNeC6y
pEsN0DjG3AULASBTzktEMhwN7geTQpgpjjzpAkyHKlZlZWZPFYSrMo1QbEiBL/RR
UmL0fa2TvjACSwlPnCgc+hwC1twh4ti56WSguo4CdiIvFoZkABn2b1YDISwEylwN
omqrAK+jYhbprY9F7BEWBTtVR53Wztv7iMMgU3H7U4+XJRILa/oUhs7CkQipuJDL
Oo4ocHfcHaO+8jTjjRKj+all0Dw1qeUP/mvY3lepGEHN4iyVseEpPZcwT+qH7dEs
dEUC9ggYkQRM6eSAxIckNQazlnqfp4emm+16p/4k+8sFZxvrM8mue25tyddUQMvm
HoIcIF1m82qLIqf48OFkSgPOfWZsySO/Is4MiBhrUU/7B7wCdNdCgC1AY1vw3ybf
zogwOE1RHDTbeYI26JcZbPf7ibhJffvuPyCPV/qyEzgAN4gA/qTrY2mJAgYOTC6+
zmQkbjhm49yOz4+rxkkt80tf0+NNm/IDH0AKt9qTsYncQuEcO71/ZI6xzJ9zcktZ
rtbdpHgJyv5M6ghc+SUXATRHmKp6+kBtH7TahjOMKIDbR7jZeJUf3MiHdnxfaDzy
fAzSBwbhCJvb1aBo3EfitphV1/g/YwKCYO0zgOMjyf62WEa4LdbufuwOQd/r5GsI
1OmjyJzQOCq6dNQfnxheF1FwmJdhoEY0pWrrBJcsducFeEnMSZYZi8bPfUWePoPX
wTKxh6Zq/wFg6x/r/2/Wy3888gwtbMavlGDf9AJZbHfZqFc06Y7faWUWg1FU6eig
hfTkdQVwEGhL0mAGcterXY1n53rw/AmjBknXD/4PBUewAsJEEU+SqTz6zXU5GGCi
tlHPM1/+62S5gOS9xb3WZiinpDGwUw2ZGkZybH7khw3qp/3bA70pyjpVQNjyMoN0
SE5EDJ0JnbUSy49y2oNIoWxqhwW+tDPL3yphxRBLN0t1iVC/M+oVeHLP3sln2QZl
HLgM8QZmlg7ckdc52ndX+IKInKhoxCRkSxt/yGPUD7M+H0xNbc8zVg2upb/8ypFl
IapCd+NdQoUTtnDa+rfBvnK//qz/C3XG8se6nASWOL6N/pkhpKVqKgAc7yLb51Oq
XLkIfIzsAYgKtxmeXX5VI0ELSJhpza0cIie1egSv5sMRUqKFsagt70Gc1bQyHXcb
jZDHKgnciBttna+nRK+d97jPcSRujj+THN9ACY+W/1apJ0BjBHQFIzFh/ApbgHk/
ob4cgK4IoqnYvTrWFAE5mVF6RGnIu01MTgsln8uffOXCxot9UojxXwr0ZG06Zhx9
2tmkoDpgsur4psHN+XEHt7o+DxKTayNgm3o9crDJyg/UB1XTrfkH3lmzhL9AuNAV
aYKBonha3Zu2WYwxfTjk8n0d6ORF3YC4DT65OjvlUGVuMVfkK5bSs6eTUd7Az3n3
6qlzeIHXOBJ71QblsxaC2kdSZFC3hZLnNuV+WBYKPnfccEgXmftC8YwTKXqA8HT/
D1FYoLmRDcq5VIuIY6iv975UiV1qH/vJ+X6Xy67SL71aC4BiaEVLhEHjZfTNPPfy
qALoFv9I3bg2EVol8pElOVxmD/rtBnOvbOPf5BJYWPUugypCZUcXPGAcqRDi/HBw
rsSUTbTBSHVUPpqIL5V5amu61sFkXhl4kKO6/7Fsf9z+8XMQHuxVmEwPJIGTDYS7
ZYhcXyNkatyIfYlkCPLavHxdgj1mcNkdlrX8QXopRsbmCNt9j1GLwfzBsVEv2iZi
UtZGU22fylsL8kTxBL3jDeb9NzA0GQdm9F70x2YQDjF+zdW4a1gCkZEakVvIOnKg
gPucNneUGzPgUljQ+jqZ7B/e1r09JEThFlWfFdPQA1atOaW/f8SM6Lop76JepJKf
juBWkmr9LgmXSG2GtfaRQG/0cSizr0dcHurgCdhlfxM5ur6sntaFrf2lp/zKfJ+W
fj7L8Dk8Uihf2lcVevhD5885/Mfa/c04NOEHS1JE+3PSK4N2RuvKUKQre64zTqqU
u0A4jEdpnLjPLsGHF7Hm3K5P+4+Av5klTMR21jzPRu87FGsHxKXrQHenglNTLvb2
8Pfj3PXEMHoHliAl+IRzieO/y1QNT2qUBJiTojFsmIVJAe7DfBMKMHdGFl7dng0e
ZYoMv87a306PoadVEGhyVucq8etwVlE90V59cNM3V89qlAz0PKwGBha2Y7poCB36
3lWIuXumsaIM+aDF/yIY3i2xv/EdRweljpFai7JZPp4UT76xkaddwW1kdRJI1RRL
GZgImu3P5dCddAQZYuk+AEjihiJOHU4OaifkpgboomUh1x1eF4mOQdKSvmGhCXtZ
NiGhUPs5aGYeKx1b6weSH1+uuH21V5H4Bu5Pr/rGZmA4k7SQIY3Qw31+0eXmBx++
eI8j3zje/cnoa7atv6ddrCMUM5cE5nQ44g2guRQrrZpkeplch8j+AYOH+0EyALLT
RnhoAtzDc0jQRSCjtTmCXKxgotB3h2TqsouXoNQ4bR87Drs8LlN69t9sH9IVG9gZ
xxwWhn3wVFvjQd8JjTWsPqazFffS2PWT3GzfVup84bB9I9KGLRiCPJUociXuQ1T8
OhioQiU4PPvoiOYqvyj04KgSKlcIuaR6LLbRqECbNssQBlffYuQWl6RfY+67Vq5D
KUCf+ei3HUnDIqiUnoo9K6EKVc8jLO1j09xznBKdO6Y7qbSNl7JEivmxrpsVakhH
tv1fnsyVVZco/vRkArrzCLVdgAj4hRlD0/JYcb/imJjQNlBizcUyq7tZSojsEHdi
52vs6J1ifTJpSiCbAm1xNKb7ZL0H3ND7z2V6slHTR3dV+lIzw4f8Mzv9TnaoYAjf
H7WaIryreb9GHlnM5hn7aKfPa6xyIf6sO11+dFW1qCnABdDxLAYn2ScyLEHYrRUR
wNj0LczTnXF5+wzJ6wAHMFsImW7b6PjPsrcakcK31AZWZTSAXfGVCZ7j1cmsyEli
jdWVKOAFMxmXnXJGwlo0c1Wb7/09uxAn2aDE21d+H68V2EvztqAKPpcfs4bQTLiN
JWMDyXo8ASijKaTib/c5M511fin2JukNFlkC4hokhB9f91jYA7UJYiaQkJWRemXT
NrbKbeqdYePhGMyisOmCFnOAFgJdF7pUcma87YM9vkcXQwa6K9oee2OfrcJK7XP1
rX+O52RPaU3aACYv3ES4lbIXAdY4+td5kq6KBjBSVRrjGI1QJhCLbpIdb23StmbB
+bMMinUC8a1j/prwVKZyWZEuQDx7o52oATUDMGqDUmGIBAxJDTo+lvlmmksiXcQd
oOAOk3Bb5LAog8w3iWC6A2ZctTsNlZrL+e6pM8v9WA7IlXG3EpNAaRUV9MFb0RLo
gkIev9aUICZXKv4rceFJCoIfzwP+vnAXvtdTJ+AjHDF7yDZ0Lmh2Fv7Tzv738xLR
fX/qnN3WKzjnlfE46nAXEYSCYoyVauuEhscxzOUr5GD3Lcssfn+O315RVAyJLGPQ
Q1T/jb9ng4Qg/vGBmVN7MWhkBF/CObbm6R5yVsZ4jX5e+z7aXsYuPBWQPFeqCH1y
izdZj7X761N2wduFODqYHyZRnbzprKsbUZryWEYJk4lBTsoHE6Vu/TltGZ1R4j8H
d5BEf0Y4577EdU3IrnMh+7Coz8BPIhdaf6v3C5rR7s5N4K1vhLWCR722+0BuUCCl
ICJTlBdSExgkQ6xfVQun61Mpcx4Co1x1I+kcPh5LG4T9GW6SEg7f72t0MIo/xOgC
4i8d0f2bbfLi15orPrgZmSLM7dzG353qi8aR0x0soNEYJ3Sbf52InWxnBtm7lKcT
d45Yt8e3VK27AENCFxhaPx0BObRaa1Mrbw/K0XqVRaKnOeCJHv0eYoeq2/2SeRGS
+P9H21JnFHBOWsSJymTkMyw9tO9qq06erk0Ur981K+NiYNPgIlj58CCQsicPejtW
q0H7yqpdPn80BTcaEv3HYyKIIy7EpDqDey9Nid5K/3rsfGhSj9erEUoXL3iVTUho
ranlm/XH2yIcpn/fnx9cmw4i9aBnfTZqQuD2xZeFI6XPeDifYfZbiXNGSfZzK18n
IkCJpSMZCAKbjlyCpZcYB+wo6CnsXYbTTIwuOA6DZjbN8ZgRcZ9AYhEpDE3dbzaQ
+B68IvDNTV/rnwRNwO5Vduo/5hdfjK74ZbDqPOZ2qCCMLeX2EXFXGyzRRi8bmJbK
5jOIGoQAR7ulf4l5lavnbFsN/iMyuyY6q/PAOl7u7kY5lRXSt6sxFEMWRJcYN0sA
H3tTMJclvbd6uBgOhC2SUDlPJyIEkB7NeEIaY/h+3agMNQLZzEr8/4FQ/ySUePRp
Pp8rSf8BypsugndBY61BZ5/EoQTSnWiNeiSUQ0Ed1wt0Rv2rEAfb1wdO4CfOeaAM
IEr+XoRvl/0YmAB/zG7BA76MDvrnGyqz9bp5g/eGf0YKHoq48Lh+/c5Ti8atj2e+
N+knVId2z3FOBgZHDSQ2+3i9YpwyG2pD38Ou4DWhPuU7zyoHIrQ29B4G42aZaSVr
+Dkja3BlwO/l/HOT4RYTVBJVj86bTeTml4EoRszDLAuEUoIg0QOpVpVNkQhiJss6
duHlgNFSP6b5HAXK4Rom7DkDUdbcgss5ya9vUOqGkBva8dt8lWz1fljjvyUYqeQv
Iw/ViFsallVaVuTNY69dJQ73ywBN3kXj/XT7wBXjTm2jDOz43kZNKVRj6Nb35E+/
aulyTXINx1uawrjbQ+fKF0fdktFR6jlRA5q1czRq9Lg5el3QvUs84Z1+oQZPyDaE
xCIB5atWjHfnBZA9BbnNpgBlDDRW5MKVl473OmH9dXjpxmvInCy97qQdBf4KFaX0
VC0JP7LzydFJ423aCzR4P2wFYWKowUhL1ll5OxunR0VQW3jf2hKi3Vv+IYBErP4C
h4MqHKY8RPsLc+c3+LVIC56nH8tlQS+qhWsCINiEnxqElDifqOu1K/C0trsbapLg
khxj0x0Traz3WODhN+j/DgPnp1lmlD2st9HxfRkgtWtPDVhmQWpc4pEIx5scxLx7
ik1JcoBKtcNrhSfutittU5p4kte8rQhjhvwHfL0bvcXTZcWjGYW15zN9qHnRAR9W
EpkbwzVRlAJD6mgtsQ5Wqp4/QXZ42Cz6L6Cb8YnorylyAFASuWgbFB017R0d3HHy
gb2kmJ51lJheSkmCSedVuGnzEensmj/1BA6s5GlIA0y7hbUYP+C/n4qgbW4ILlRb
IirmS6DV0NIwMqWCuxiAYG28jQM0xu7VObOcIQfb+Wf6HqxX+yUDuJFa+tbrMOuN
2mL1Tn+LS9e+2SljkjNcBpsq4Js35ny4gMouuhlxgIomQffPkYU0hric5CUDWcGP
CkhR5Dap3ZQL4iOTSaPWgxCcxDp8k0WkpZ4u/pksT/JNFkWpFWHDtXbm6xi2CFlE
QFDpfz7eSw7kfvag2HqB+lM81/mDZscwYuusyic5JbjXZU+OcfqtOVEHLZXwH7qK
lai1pbUKJF/n1VDguzrTMln7r6grRRm10MmTC4r6KbzTFvz41XmKqdq9tzxYKQS2
LE7DMlcbeIXjGKKpeJMh7wTNUeVw3um1JV/0hdEBNyefc2Cu/cqvb/bsNBqdlEVj
l80rmXfcleuXgL3HmWPNO29iSAKgDpdXGQcmtGdON+z91HyMxRNrh53herLCbAJF
uMPaQsG1SFQmlafEaGv2WrqD//UJrsJo372oNeKrC1YsukQYK8KfItTvrariDZFA
nu65bctK1lRa6KiTMtb6aRt4CK8cBlJvicyaWu2toBnJnNPGFnk0u9QX2xwRWYOp
mNiSuX+3fMFdGDqnLAB3ubBSP/2tsabPw2GEuRo8fEn7AfVcYnDwvNFMp/SBpdDE
tibsRwVdeubiGFlv+COYhUCc6YFAfz9OmH/B+W1C4IN0S2CexaRsEuDLLCj7yNkV
bd64iZ58CymT3DXhLeH4H8Yec/sO02xxUyFGuYesdYHHwWJrEeGdi6Z3ldezvEZz
NiXNIr05XE85QbcWVHA4or2VN8TuGqHReNEDU6/qymizw4PVg2vF5ghhYh0laIil
FEUzoo5ctIkbLCYOQBdKMc5203zjzojwxG0y8wBQFSOx3Hp73+aGeJT/jrhXxSvZ
4lfp6TpwuKwiE254TlXMQIW8mjMbivbsBtCHxX7PSCdLObChtRob2D0uu1XxT0b5
RpG3vU+U8BJg8niHR/Qwnh1mQCAnjWspq/g1vadNvaGLjslaB2vUt1fwuid2ThI8
ubJw90wmSEzKasfx63EA3dxTMe2AG2YhjcGEFIcnOmRKGHEHRB4Z7f004DgBUkBc
v8tXNRJNmu2trJ32AYOY/YxK7mp1ShILjeq0czbMMZDwgdq15YIxRjMUf3ZoTk7G
YnVVAynupMLmcEX6ctPNeIR2hK0g8nBBCKwGCLTkadgtpLPSXpvKtReFQ97j/by5
4psvbLKIU+PgECqLbWZ3aTSvi8dY4i0r0yKnpCvTqLyTlxTu93OsKfmLt+s69evt
owxwmHuttO9QtHKjsLwyII1xnuU0xbOZYUEG1wLI7ijdeSubvBxuBj6PEdZfUu3c
N5mmfs9/d1h4gtXJkDEfc/UgvLqYYyP0J5YVZRB5de/FSVhfa3UPK6lhzpA3XqYP
im+SbxuVj4/1SqreNu8RMoLG9sNBGarS52Nx4O3wHKSZsX/8VsBwihw/wCoa14nW
+3WjfdFDtw0ebneFoSwU5v+fycmCFKQ6YLO+5Ghu+SGSlSyQrcfiMQ7kRIAolrgh
tvbmusXga6RrIZ7BbpYbLypoUAKtvDuso30AgdMdXYvVW6ADihYRUcstbNNFcr9C
S4uitbMYcdw9JPb7nT2KpX+lOtKottOBszxeWxnV++kLeYjNlHfpdolfVvumUhOG
0+aikQSMDfReCcFluhVkB7n56AyZqrRxjbXbsC2Ly1CHHJFAcFXSfGcRxNXpACEt
Ec04D2uQWiBSAG6Y/YqhOu1zYLttKduNcXNHKSea/NDTvSbmXSuDcOiJaHlxio4s
VbBgKduaHYGudUNXVEPkD6OaCxT/FIIqRhU7KM5BE5eglVnInymef6OU/SzbhF9P
V53qhFlopHUk2YPAnCCZP9imjD2UaUYl8+hnJ/d/3f0uK1AhaSkHKlTb58O5ebzn
TjbT5kX8bTH08UVY54ml7mr5myTiXGn7NcZKRihcPZG8udY0+tMDtyTuPGAe4xRN
2ZqNZC40mEhj7JHOV8mGRomLLrRX0ifyIUQKhZDptNRzpM1qcx9ZfFvBhaeuiSHC
1GcMd1qOmOxn7dE8OZ1G/TubWahpUqJRUSFwKgFAGxEt6IxeoTGjAlnhGzap7vzU
1P+tbQVTO0LxXH4flHW5qIkHhPWzkOINS8rJ3P70sbCvS/1runZtdgbhMrcQhp08
axa70gnUCgdrcHsvWMU4kdb62YVXzT2DP1oOFUTjvg8017iFjm9m5poWUyepjVQs
U+zHh18y0Z13LBj+35stlM18xRxAqIt+5/uiUMOrRxu40kZIvN9kcOqKe/5x7QWK
sUcdK6J2/fu+rZj9RN+HF3wl48meL4hpYaNSlaJPrdUflhomO4j1+WLVAnQ32+AO
l+6UD56cIXOxkmodVD6hPVMihis/f0FfQjXIOb5QHTiLUN2YrAmk1T46GcTT8tAG
hE7tWPCR+i1FHAd7NDgSflzdJIcMPdpb6Pa4aVP7EiJI2iLCc3eFdfDKVs6Jq4pE
h2Zal2PdQjPwxZRgSJiCjdQetC/niMYp6fy6EpwbnTS9G7xIc4jUvHAfBrlwT4JV
m6Cf5ThdfCgIutA4gWk8PttJjDUofgKJkAEKxi9WBCqcPKnUOe2n9vHkPL61L0wL
HGbY2TIOr/ETmdlHqlO4pixgJXZzq0x0/eDhT9LUjV7D/1Sqy3gVLohEwspuKXZa
uIu8piQLPy0h+KTQ//PelbKqgsgQLOvYkVorDK57lZW119UCXSkO5kEu/l55mvmr
1dF4IcyDShj4TJ5u3+rZmi9I/IEpIhDDovgvVYSQ4+nILpFQTIyhJmv95yX9cjpP
xUVRLEQifZ/+3nhFBOlqzCnQO1irGPVosZ6nl7sXAd4DbTWIBvJ4o1uJ7frGLxM3
KraakyKKJ1CC6PI8J6riZ9fS5n0K26xAnnqwaDWwIPvVawtId5Nx6O/AhR3DJEc2
Hg+BLsDJMcERQwrhroW3agVEhe2bJxso3M1SxzxklhGIB65zHIpuD+0DyduXfahy
SHVm7k8gIBY3xnoTXxJtHLSvlRweVZyBeOOd1D+U9W9qW0HsED+qMuOsNmiH2gzr
SE56/Zzz89nl20x8MaAyTgkkNyAQ3u5PrjFrbWm0RBirrtwQlODzh1tU77Eg9XqG
NvNpDP3cAYQdT9bvlbOZhsV77U2B2BhbvVjbkTDcEDELHL+bCOxPBqtQDj/nk5NX
jQQdO0NzPYRXBjKVIRqlIj5RBzRHHMBvN6bInkthlZTkEf54sQUoFtIXgdpXEr+G
OA6Kd6NbTS7Tq2Q8ECg6OFTZUmQxH8p+74W1BdXsAwq+lHNWD3p2YlJKzhZLUz7K
23T+DFjCXgTVN8bNwrTcAPCiG5ne6lO1KYFVKsS68ezdPF5nc8DZL+40F4CS8srl
yFuNBL3D+2NxTAD5uYzmaIuCJJpYHfK0JInYOdUIW/Pjx4HR+T9b96lYot6pVVWr
K4gsj9hFNsyWcvXx2dqq88xOkCILalTYv1yYq4F/SuASKNFTFpeQ7k2FG+ua6dFq
4s+s9may50kZC/1f5TDKiwNc1B52OvRG68aHC09NqKh45/jARp9sDBwh579FlW/h
3AYWJ3gEuVyQKQY0L9G+P96kKYuQNtt264QRQO9qVIRXOLTanrA0tWut+HXu8lN6
AgqkOtFFLFayOeIqz/mKx2+5WGuWuEcHBOJKhFfVtkjZnc7iuLArib2gZJV1Eu9Q
tUZ+4y8C1WvzWet1Uau6bi+NWjRarqUfR461wpNoLCfKxF2LLX5+ck8jgk1Dr0z7
Dwnp+SqX7ftwxm2vP6X7Ge2P06SSdW95FkjLsRXcGT/iaCJ6YYJxLQWrOog8mGPU
EJqxO/VjlOZIrdaI87BfIW5jHPtb24bjzQgZ31qUjwoB24DfozPgebME7FY1jQYN
dyNMIBYmOiyP5I3dvnTNbGkcRuH0NuYzOSIBEmxNiRXP9gW5td49BNLpHJaBiRrt
XaDGyLLFzj7x4dULjsvhRi0CMb7Acgho1ng3DvI2+eqsHzf6uneDKAPTDIteyLLC
nT2T0tXj3NO3V22Tm2nQluQ8FKyLPIc2xKrIoW6Nt7Gr+Va0wVyKV501X1sdbo/V
`protect END_PROTECTED
