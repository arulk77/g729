`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGahCPvKVYtO5O2CpeVw4MWyr+JN0h2EVIIoMs5nS0vo
h4Er4PWLntFkFM81KyLgqEolrE0ii1yg+CVFdFnYiMqqh2Kh/U9zGkO6cbmcg/Ea
3Ibu961jBJZHqpuF3BCWoGw/qqrPHK9M22ZhqqdYq6gcLPS6uYqaBSYrBls/S1Cv
`protect END_PROTECTED
