`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAaBGyjbxNY6Jp9OeesNZS0mqY4kwag+i8Sbcwz3+h/Im
d5uLtoYv2EpmdVlLGeqn7+pP/+e1uJY3R53DXwkiCDewqrcTaWKtsmCugMUJmfTp
M3Z9x23IYqijHQy25hGrKdUc/ta+Jwbcbet4qT9I6N4qSXh1k+I/c7XkJPlw/8fT
qnStVbdQaaCQYLZ1ktJZ/2f84SPzGGqhcx5PMlNBxc7e5QV349LQ2YvLxg9X1ADt
leTw+pZeO+rfwLUWW/3R4LDuNlFSPb4PdCkmot3Ln8x3hXMrv2KRNmvec0lCctxn
CQFCpUi3E9N7yUEGHFr7CsYILxGWtX5SeOnl58fcLfgikY6m6adb6vYiATP306sk
zzM05LT6V749iL4HJdSbSKklydQJSpPxJ1x1Zarlfx0g+ujbadMJ2hmj6LdKX7xr
/EtC5L91q0hmP+QQViQ6RkJLoggcXUeZ3Qi184zeupVcU5foUkNxtKz6bB+nIscJ
XlMia+G4ElYbMfP+IKJHkMtlGLOORJmJSS0se2DAD9UQcmtcfHqo7CGoWpvSfd5i
zXTHjCR0ptGQjlOePNXOYCUbeDsRFdLKQdhgL92p6HJTzACKtqX2k9LT1jrrHsTh
MtbWA5FDRsdyN1b2Y2695sLYTi2TCHYhTFBF4L0m8bhtcIOqwbUiI6/RHZz7/iD+
tZDKRzTuVHbYPyprEfrB5CbWJlwX1mYe7+it/vlzNP2yAzmMFBne6sC+jbXY1Seu
6MB+mHEVVsrPKy/4wiuv0q5Fi5/saQJt81y2Bt0m7oqW6bWYDQgHZZ8QIeZVvH8I
SI8jwrMK8u8PnjFrk3SYpYVlSa92Ho3Oddsi9NRxMFFnWdh6qlozvXdQjVJMv7Wg
v3LUWpj5LXeDoa0q7gYLXEli/gsdPUA/ndynPWtlFHgeP1PA39DnYubS7StxpBx9
LNyrjeVW7nkSfbR4nV1x8RmzirU3/+RLXRSavK0F0vAeMAeMkkEODo4rm9/S46HG
A0f07JJHGJCLEa7Ntd5WGLoB05b4yowD4GVEgAQ15XS0aQOdZcjRd4tUEykDmIlG
jVUKVizIAOpTDr0fDw4GQMCp//faDFPEMSSHp1OMhtO/dtZHEGnUpKJUjAryRtQ1
ktENrVUtJG7qPg3AqpEth7PEGa/CCvhItYRV+5PFa9o0+//Yq4F2Nbs1V+6d4uZc
K2ySWWnbiwwzmp3Wl2zC9WMHbQQTjxU5xkXLO0ceihQd2BpWlTQNfFDM3xmJdNf8
vSy2D9wypAqUc5sMaFBf5YxvSZoSzzxdpF1DKNCdY82gAeBKyShdBsXZFTpB6izP
Ny3kS7aUlHg0MJnYAu4TkH2/yLqNU45dHX2dxKAcfl1Ioi08JfNOf3JXK2T/DxPZ
YJkiBLfUNv8tnDnRirzOPuemJKvWMBphz53BDxs/O4FxvWFtLLurX9SxSlH3k2WS
oikC7W5j0wES6Jv8NPnTb6Dex+y/KIpQ4D+qqgmLF3+DBwnQurtePJ5WuMIHxmc5
RfolXez9YFZEnEnXvO1KweZrxNyplGYZO+X7xqDg+lKCf/XQeRy0KlplDrswb+Dr
037kyxsUjIp9AeKmSRcf5YA8KOS3YrKDbKEttIMUN9bD4ZVXVJdnvtlmunmDKWXN
aopvfg6i6SNSxc73BFUbn12Pdi2/IL4PE3IhJbuxO/FkRhB5Se9ThBlwcws/vPK8
XTbdB39BL4dcIgxlsl8TDBUotwK14+2PV5zSt7NbkXJ42cHQtLeaMZhlXWiU2NbG
rBI3pqSuwnw3rLe+HjvlGM34QIHiO1H7l6Bo71Mj+wtb0CTrphKFers9A0tjOnBE
aO+YC0mjfL0xSErr3ZKUgTBlxUDKScocahiJiunXvFIA1um6sFVNF09Z6VYKgUVC
ty1PCFDQah70knCF32nMEjRRFZjWr9BZNgO42xh0InLZPSHAxqD+WSEICBiZi6r2
SdHx1bc37NVuq27oJBSA/NvYl8fy2cFB+hk7zz4ZZ8C2sdRRXS9cptnUIe6KuGrr
4D8LcKaygnuZd1lLDhIw9/wYPvw2CVIOwqnb6F2qEsq4XUlzEpW9rZ4rGB+KV25G
YwquyFl/AvQoFFEs/HFp/nVOAcsc+cTYJTt2mE3KSFMXldBa2RYHkHknsCF02sFF
E4ewQjYzfiGfXdCW1+HR/3Vy/fiQcdILvrATmQ7WqihyCwByScRFArhmfAmPQxZy
TOiv3C+IkxmVZO+JOVjXebGYulV0LfRQDuD/FVZQZcmCn9OUrhxFrkbgZslgrKbv
Piq0knZQSLIz9D4fjCqtxhQ47UeqdeA6o/D78ENjETbpwWCvZT4pfPO9J+C1XIw9
4eMDHoUPqG28MhxnrPgT+flY3V3+yEf+cp5i3q1rluPbtPRR61i2kkQkZseIWeJb
IoP1DaSRNmlapz2axlITZE95MGEyGbDsNBPaiyzsDFOd3H1eXA0T5BWqSU9Hj5Wm
M/jwEzw/ZPZJOAx77JZsVEmGX73SE7QDJgR+Npa5zPWMuK944ICpuP0BvRs7rpHm
Xcum3UTCm+wpAEWUq6vFlCZPTGyAfSaQBmBBXZxX7FLJvDr3AShsJ0PcXVKft+51
WB+YomY9iIbxv2FZTIHp25RSTr21oOQ2O/YZcnVWU6+KKLVBhHrNdhsgU0sSRo3U
B+iF94OToc9VR+bC5cYrZNznzMdODQ9rWsf4tpTb7Nxd6ES62mwLUaOwB+aaSuwa
W8N40OzvZiSqvW63x7zTrBlSMD5C07CRMbsVKKtJaNJbBAybOZtaQ07S3Oj0UCxm
u7nmA4U4fvt91g84rtnIKOsMu4mpNxvGtMmj+xtLYRW9dvBOVr61g1KmzSpg8zcq
LUh8Qd0tCmHvSoo4n9lxIgL6f7w/JkDZPNgPoNKI5Jphc0DxqG1QDBhGcdIvtkvi
UwDrKPT+n2VcWMcKKo07eCeqr+9MnucOx5ruMfEcxMLdB9OEWqiBabukiezHUm0g
HbV4yk0Fg7TNYBmmoGpRc8Qr9ztSsRoGoytXDQo2udL7DrrCTyMpDTW+yvxo2rjV
LywQ+w6tu4M7D/FnhIQ9kVgECKCxPENl4DfkEHb4AftCSf4KpjyIYBQMElCGtYlQ
fQqn9354mYLztRnFnYyQBs6IrQSqd9eZTYxZPDnuL8yhuw+x/MNtIr9sBm+WlZl/
gMk8zaw+vyLyR1V0pJA02dReWM9QU5pVBaF+hCME6NmpttEHFboEorlZS0AywNm/
RoxIRCfT6Gxy73B5xnLRS6Ezs+86qsKIENHf5jUHcwCUA9q7vOynL7B+HZUoe3tv
ZX9QQd4dze/90JrCZM5Zl/41Y4hDVy4Rlx2USd3MH4ZXktkzkbb37BRgeMpHuij6
HQgFDeaGcY07IJvKjmi2dYmfcukOwylEA/6TT4dU4Gd0deTrVawhm0lVVNBcW/fn
+JoXsjqmlvZxh6ztem4ty2f/OtoM73R7WdUETE8KiqeDfsy+4/VDtdmFaaVtvmSx
CU9HmED8ZW7RLkIdZBkwKLSn9N3E0xbz/4NU5AnpYd28TESGswvX+l19rKPIzZyI
Ml8J7h5ABaaMrcQFio/U6Jk9uuxDQr+ri0+v5O9ppa/TH/HCdMu9UNCluIr37Dxk
cI+XlrhDn/U97lYlN4P7JKOInPIA10E+rPsPzVPngks6xD2vXL+lam4SBT+6LV2v
MwJRUU85zXPwLaaKkK2DHTchSzrtP5ln+RNN2Foy2rTDMct2iWP74KcaN9xHGXR/
Q4j3IbI/kxAYd/DiQOF+X9nkSWZ3BeUi1lAvfvIvXcpySXEhP0eidD0z/tzeYqP6
c9yngHkITUiBmgA/CE6mOIaOjTYlEwumm0kEXZGGCIa1LL3ngJjI4n9FqzaJ3FNy
QBVco4qyvpX7GoDluN8iVBMzjye3l3OT9+EuZYahPk00pkVn9eUUcUtxsMkoB8NU
NvrAJhFX37WHCmN1RCzA4kXJSXYb5ONWIa5U6AyrQxtARBMMTWf0xerw2YV8erpS
BGU+GTbQg8KZE7P0U1unswLbUBaOb54PHEvz1JAcLJIXEzomT80yBT78LxOKr208
YdLPNzBzeDzZvj3aTcF2MMMOKsaR1wJrL++6Xt5rOchWfuIeGaScJzJCCEfiQtBI
ml1TCOwBwPIuscYaY6QVBX4liSbNDBFX6QK5VmxXtiCigaIxba9uTeHY0JuNRe3f
PqueSJnjjt3euY25+C0w+iQvziJnmPImyjctcBsrm0mXsQaJvWb3qtFyrqnPkXq5
iTODW7fzDbKYFDtAlo5Hkcr+BvOcGG7eLdAee18mN0/1h9FR6r/tfao8xuJl3Epj
ThNMTbzHGGcyBaqeuxfLtzUepEnI2hXOA56QYYZwnSH6XzNZxKE5gb80u0IyjlkX
99PqI0bFRf6A+CRFaPgFAmZwXk/QeFMY+oa23WEXboeR4y+r94CucIAjHAHkEIjn
EXbStqAqya+PUfO3UjPJiZdIMzyVlu4A5oT3ONm1XdjG/5YqZkwSFvZ+GMrmHJ5t
Ceal1svx/NvHbmE8HQ+6yLZ4lcrL+OEVBmJvYU3LSylPcDhXu7MJ7QwuEgZN8ayZ
IGHQQ6mdMOTo0X3hZY5/6liDWcnBNpGav6QSRzIQLVT4AtRtFZt7d4DGMdrgoKOe
zKH+a3fGZuPG2FVu1/aRjkUEhOUIwrzpWZ1n4J7A2bQxzHSA2v8Uq1apqmlaISOS
D72+LTICj9aSZ70ZDNJxTsu+lFVhR4L64B7VnzAAJ9F12Q+4fHcQHKzawsdHO/se
rIX3d7/hZ/YCkaNu63MrxK1OC4pX1Xw99hBxb6l5JMnMetdGfw6AHBAWk0UwwIeX
QqtCJLbpc9FP511jX9KTyj0ZovI2Cf2LHwE0VtnuY1Ce4IvBR9xIiCeJLidQhBmZ
GocVXS3q3fUe1P5DcUBgX7RxN+0ZpXTnFKXmeOu4QqGJCcp1udS3FMSjC1CXReLQ
vr9UpTSKZwwqYoQjsv7Mr14SUZxU4XNtvlXimF9fs31kMy73hjZDt6EyIgA0x7ji
tqHn7Dzv57gUM2nXO63dh5u/IeD8SEKMss/ZgUmrePNadp+RCr4tV88dkITmkMRi
6vCawDdiJUh7bYXSIwQtpfdAPS1dh4gNNI+2vuYF2GRhhB1axQ0HHMy7U6u+JvOu
wWJp9CN10PqInL636bphzpZiGu9D8QlcvLIrpL543WAcy73uyv85tCZZEIsdTrw5
oii9rfTAR10mQembtVqiQ5lqj9j1/qkwvJq7ntWusj9mz9ZkHB4YeEFiAOY1uKMY
DrzxuB7xvneKUEo5XJ6SZzsFtQHrv/A309Ah3VpmX5nMx4hY+P8HJfPjyfbfl/vx
4OWiDebFXjSDGl0itsFTlT/BHSmc/fzQo6ODp0ZsyuOrAdJPEDuBBP5V+FxaaGVO
N32734oMwoWNxmDqFJn4MmEJaUaZM2xvDVaboigkiCeBoFmWz7me53HqfQYJGfnA
Puw583x2LMXD/Ci5ObmqmUuD/RBGxggG6DubNRNgMA1hYIjkcME1vTFy6jHBOH0s
+ZgEiK0B1T5AdRHicmtOvv9vp7cocxEe5TvmpwGxULmpaFnEI+G9kJZ2qTfrEbGE
hPpEXAbawheCNCTcTpuqyiXXJ8fB1P7iAGkpT4eFVyGpo11w2OQNs85VfC9jztqX
mxyCxWVRCEQ8Czousv4j4UluPBz5i2aWVzv44vjhPZjwA83/3QSDXGkStyx+/f0c
fRXZaY3P2aEVTi78aL/c67trTqoQoNmkWIdYeixYZ5p8Kc9/eHZu9m/LGendmRkR
HbGOawXpiH5om1B3yLExayrxG53hnRGXpOTIreR0/pu/KLFInVpJwfUqVRAJ8V6Q
0ByHfLe71MOkJaESAdXF/cbOiXIrstNVKewjU00/KFAC5LdnPtAIlvNuexIlEQrx
lyGMvaalbqxC+P8vsWsM/jKtq0LIUdyLPfFdQJN5hzZLb7jmztBfERUBEPjZ4e7o
JAV17kfdWtXOE96H3QUajSfyvLry5RqxmhSepZnmSTgFNddfBuWhGRr+xznKcoHH
WCSD1t2rowpmMNriB+nwa7XpUemtHkw4w/QTORBdV1GlBawjikcLcFqkS3LHYFHk
9AEUFhy0ghX4+2DNhvR04HeD2xjMOGqgeuhPep7CA/FI/eosMhYnh4pYsg+8JaQF
kmwMcXFL2o3B+ZTv3a4tySnNppxT/Vfr8+Af2j/xbC08yHXtR7865bMJNVB6dmMP
YZA2Tvq6h2mbbW0XEpOUvwT0RtY+Rup2SAh8VdAx9E6PtwO7vSQ1yS+HfrtCxPm2
MJB9c393yOLTj3LCA2JiK4x24s/dG+OFFJRz8Pe9zzDpRI2JEwcSI5hdrVTfQhNz
ig8LcHTGzBXQoVhsDHTZvZhUKhb4Fx//Qkg1GuXwGww1uy/WKa4ViNBGs515SdpQ
eLHnamVhPS+batzBn9BuJz7seXl4vFKUBFMo7m/6QusLPEJ+HGEM1w4NIRgh1OWE
r/eZHxgOKd3ZlKBX2HeLMj6exikieQfEKNo3whBoZ9L2F1hXLP2YRLttbXFfj99y
Oxpu3Cif18TbYVCIF5oNpSmkXfdXfWqIfRKf5hp8FdZ/SaXZSX5lLU80MgeRovp8
zc7idXAYw5+3VRCYmPy6r2zqvU/8W3XypASjgqioIF53lcTDROwxwt0VVGrjqTeN
F2mZgkqkVoB9HlAv6KG+awNfffJOoV6C2oMLImlEeMPyMXfmqLcWSfiqF0v6AKO2
hIF/6xLBfZA/1GwEZCTtkiLOJduPJYuEmpdJ0wyxe5XkD3Qm7nz1nezVoctnILg+
TG9TEVrrizAQjYOrrOnKdjrBoO+/Zi7p1ftaHUWgOLkT+a3WaDj9Ou61JMSR/FOq
PCJZ72G4SULKfcwww+3B8vfkyj/Zy7vFQoSTuv4adwFlW+hX07pITk95ku5LgQRA
qyH14ZUY1dAwaSvuF1T0YYShj7/tlo00i3+NVXFCY7PXNqCYUVRHJ/N5BXxXGlGC
iIdWnLqc8kNeJhrmcjqqRzyMkAQSxEKIvzTd14TPYKAAfHzk0K8pHz2u02jj5kj3
OsrIfdMYAHWxAM7DoJqpXNC5SVvdNFBUuqptp9iZoVwsrg1+Xhui0HWRUaSRKvUO
VWLnd+SnEQ3wKJNFy2Z93VrPTYnmuAIRGO3j6cEP56vP9qJVnoYA0wimfNyb3JD1
N42pDIYBPZig5OoB+4AGfVWugKyMGRlplLYB+1RKh7fWdk2yGt1ZQGuMORGlFqmA
+BZhpPHaWnYYh+mn+a7IteQXDlpcOYfKAerDEpLk8c3x1Fy4IFblh5ypLwShqeE0
worHa4bOXst6rt8gMuObekKrHQCjS+9cKWtUWmCpSZVnq8xDNpPVNLmaYjOdDTPp
8e6VclouSWhPaQtsuwU/SlsBtYhhoPfyxvnWh6CjMbXjRYLjaJEm3zW6OtvEQvTp
I+uVvoLOtgrfdmCXXYVSgY+YhH2OFcWLK7H6T9B3uWUfPEBHJ9R0lbgRK3ympBEc
10KGtpCpnhMb/W3a5iJBVmwpy+mLNn0zT+NB+Ctf/AbZuKuPyI9xW6cMYyx2jKl3
bah7tMERBqoGbJtieqqYKZwUfOpZKdZxz+s805MpFAHec5RZ9Pl1u3gVTZopDsWn
BlHUYJKuLxvEPDemv+qOemQt2V6J3RxWVcBahHziqRU/t84opPKmAlh9KxRTMlMU
tdLUTdW3zAkotgDYRElGPWbd5Ni3x0oeOIafZkB+8GNDV4mLJ+HL7Y19PPPgvjJT
TrrxgiNcAa0iDdPNNKmspdEW7Eqd/geFU3ZrSdm9tBYNiDn6NYDi2CG7bL3LxNkf
Cu56lNY1GBUl6wGuorgx9QfR9EhOSx3ucfQC29TPjMfLblVDEuCkEC7MgGdXzwbo
ylVdAF/EUrIdTjxu+7pdmfC0ktLVPR7wM9agdsKGn+Vx6XHibZ5oagNcX/LUwHNI
aDGHqTvhkhotAowAiYfp/6KmFm3kOiHj/2jZ3vUxEe8S9Ukvh9WrU/jZ7E8PlLfv
w5aQ7gb4N8RBa8MkMzS9pQ5fc1nUOvQR3zxzAROqS7UuVk8Ts9+tHTaAEEiBsgLL
D+gQl8+nXRMfruGYLudGuGp30hp/Ryo4ErFiQW4gPWX86VHmtipKIAiJh+2PsXa8
jHw2XGBMYUuy/YePLICK4FSqiOo34S15YwXfz7juNBVUBPJ3h92tTevM/rbFRW0u
n6p80vZsUTes6WHRxbgYEtg6jca1L3habldiw+GkPVF15akf/BDBHQmytJaa4T0h
QszqsRLQQRT4FehJedfGFA4a/NXynLpkxitGyjDyG6CwFkxLPXH/751kbbJ88uJR
gK5/YTIp7bNWr0vwPWg56uFdSpWjhzHTaYFVjeMnqXw4aY9h+98kI0wnuX4+75g1
U4TahdgpbcCla5Xsdd1cnQ85bvTJjHu5BIs8VcwwHeOO76hjBAIzyuzmzDRzUoNn
CKIBtebTBVUIZ49PjmQPHlNSperqyNeHw6oVjrYeGik7Wcyac84m+/u358zzx2N6
E+iZvGxvbLE7eMcAiElV6UW/t5DbI4YRCuvyfrT9ucXI8OKoVsshgSEy8nbQ/voP
EqC+QFWTTkwYaTs23+iN7iEzLUuH6Y13UzSkxEnhpuAIJIxoM1JrE+jQ+puELcpF
+WEN73xiGMnJMDRV3zR1gfxDUSxId8B7TsSK3PjWlu6jhbmBqwHcVDaMJK9qWOvP
s+z0p4JQXtzw4c30Im16mTdZTcxuJP/C12dfH8ax1jLNfJnS0yXgRsyM60AM5wAk
kRDd+jB2iu3ivzVROnlWkinz3DBUpFRVS8hERCRj99g9YHrLQV9AZNeacwyreink
n+1xQOq4scYcJu6u9sY1U3EmuR6m17xO617CHDFTLTeNi8XvGCPBeObFJAcdZQou
fLQ6+fXRfULwAQA8dlKOyrIxDMWR0UtNQVpTflllfGhyUbPAp1Gnah30kOO32xnr
MSh99N169D6mg1H8BEBjy7ETAlTGyDFMeG/5/+5ddLS6FwzCQ/iQFy0lg7q2s+bv
b7cNFVAG30UcoYhCNZQzbsmJLkP8ArWZIuwfpZ58cEVT7RFhDgyanXh+8vRkQwwQ
PVUo5IWTBwe9f6iLbjvL8bpagEICY1HRxL7DdBMchjZHivNT2seYRWQRoNnuJnes
y9M0pjFQ20ytsm+6mj1PadHkp2J+YjlZwhR8fjbkIQOEfxfNC3ZuPiaO8noaji9C
HZsw6J/Qis1AjnybDQB0LAUfJNK+A6fLIgL5+snBdhP3hb0C6O1fXy8Zkaf1Ebqf
MTgEVKH3uqWdEpHv03lFKHbsB/d5GvRMb82D0iH0vnIQV50YGFsAPIi9oYxFrggA
3diZ2qUOsY9mw1h0BJHJWQLNGBTXtSwo8Pl4TLjQBRKGOOmG8IrvPLkyBrZiWt+r
7DAQ1xOPsUPXdiO+vFWRADqBPnS6/0c5v99GcefAg862JSmDMyY0SNbiNYxpLr8b
8eVq51RLzlFERDnYiGlW7TU4qeiyoG8jz75+GsU8wE2p0hkqjPMJD/rtPzvhUSvi
sjua++L8DGMJFDydupMi+4eb/2S3XU4SdjWe619oLTaVfwvUOgzIxtaauT+HlDmZ
F8XtfO8w971kAD8T/BVhV0469O6iB02401+npNBD1zR/khVcJe4DmbNKEz++A9Cd
QSXrhgiKfDaTPrh+Bzt5xx/EYrAF2IdzLqQh+n2Z9bz1GjZbcv8o9+bUC8N6rBE5
s79TxGo7YTsOP1h+S7FJIrI/VWXJrZVFYrlPTBdG0Td+2WYywSGvqVBV4gWT/hKW
Pc2Ppn7bRUqZm5reHuBSiUyZ7bQZ0M501J/UPXq400WDeeMkVMiY4PEHrqcerzt0
FqpVGc6BECiMOLrCCGl5qdMZ26r5Qr0Qa76f28EE2FJLJD7whaEsWqeCU9boeIi+
wR2vR9pQhYsL8HCwyIWkNQ5ihBIa1o85BZvOh76NwMFoGJS6qSh47IurL7nX5JFS
V+xEWZ+rbB++x5ZO0aOCH2ZnNH/MgUTWXrpx2PoZO8iix0TQXNt+TL45Z47vA1P1
iBp6k0UcgYhXO/AcZScW7mWsCkYaTEz7UPRR6ERogt21lJYTl3HCLNKx0DR8664j
ld2h9QlmGE8iKo881bEZOnipsGBiIBwvsi6NYAdKSh3Uql3nczadyiPzwjufGBOE
+qQJ1CUmqpF7xvOPBOR5vfQPYAH50CSTasPoKmHiRPNpt5GTotxLIs4qCd+Yc8Is
rVtjElZdebvBmANmZEEnKHR33VHt44bYWolgWdRUbGAL5zk5+AFMPWyW+GSFXXxN
AwlkrHtjGfrpvywGhDn7rBUC+G5+SwiOsTtAKY4NBkRfcGWpa0m3RHzuU2xZPRye
dVu3r1wFblYnoZH/psvo1jftnvI6e3bINYdTjubgpePKyMjn/GRKMjzkQsEWkUii
DENcWYvHD0Nu7sly50jQbElU7woZf25TbyYScwKSb5gHWz3Sh3eJdtSfw6Zbjmrb
bOGyBFFbS/1nGGeUncL+6421Z0MPE7f2+tquZnA1B3lC14lksYSg7TbLpIBAe8dI
/xpMTHC6UewBKFlPXOIbdYAum+3OeJldfwa+eNXIpFKltht0/fgcXAyFZ6bxQohu
QLo6rw1n1Wn4Mpg6XmUj59Z+76mxndv1sIT7BKiwQmW+qHc8SQsteOOABoRXV+pQ
3ulQFbzWgmigcENSlMdJPNq45RyuYMc7SFmTbYZeFgOb+8tpFUzRF+gkh9aS0XQD
GTTWcYtyZ430P+ZpgqwUgq6Ena3f/rrMtSlOIgx+lng8GfMjgPmqFVJa+8gIhlbI
SJMVGXAtn1bqL4CzBhPKRUwe513MeOoSPbLJ3FKE6YwwTAViWiuvO0zxgkBxF8dI
zYP7F0Z+gfhokZfartMxlj6KcTvxZnu4UpkG48b9eu9EE4U3uFOqUpUeQji5q9ds
vEgbNB1tz7M+TVyyQ/A2zPH7P0/rE2fXp4S/lA1//ZwYNzRSN+I0rL1tSomStpfJ
kGNmRunPKiBvWi9rdZNI5yBIsuZvXOimvqy0LBgfY5DrSVqUz9L/t1NgOk+49ICB
rF6tpmixNrsOg/UWtTkFvGB8QaC0ljCTA+NV0zZi7fzzuxJ+UZ2ftPu6yDbHagkY
AHp7pP2O+7+gZOrQwB3hbq22N8DY2eG54EeEoN4qd1e++/ka84nAt7KriV9uU4Ml
GNVBiytfJp3T4cVrEZ2BG9Hc3EqCcpGCK1bmYsUCTZHvPhtKW9Ox/RsRMkxxU7Uf
nkKQOATHP9Xo9ZvqQWljVQVlcJhut8CxdMrrx2mW/ZY9iS5MJqNzkr0Q+8wMeFEp
MbAKpq+m7vlaQY1XwbDnWj8BNtrWVwxQUVXR5zC6ZccQ/MCMEJm6om9dmQKue12q
vgKu3cEKYRhw8VU0xY1gghyoKP/jmWurU6CBdBPBjRtjMiCOxrLLR3vV5QdTYeJm
SykiYindhM6z30RsfffXy54xdhhJi9wrnjYApdlLE6UNjTE8rhHgNKdO4QldccR0
F/8M70vWM60W+aTBw6X7xjPjRdH3p2gJLfdAHAQSZZd2UfE+PAt+e8vM1fBuJ0Ks
tti4n2zXN5VcUfDcLy0HsxOQ8tAdk588PMsXq2KdZO4cu+SDG2D3cf7fTH9EEZoq
Sz5ygJH9X9S8vgJrtBGJBcehM/qk83I5VnSEqi1x7rarhREmU4CalEqT6mEmNaO8
G+AJfQfkDElZ1nCybNTsxQV2W+pz3FC+rhWzLxZXnSnHHp7LXFuIixnZRit5WNd4
lUpMXOnUHgJW+mW8QnLRprioVEIj06CotDNwNodjPlp/SBbgGeH8r1Vqowa9qVn+
/WPi0q/L4OKtsKrhi0I0WFNhmI2aaJ6Wa8Q4txenJlCNM2PHgv5ILYBLLEQcs2lW
3b6qmDefbMXzNSOqfR3ap20W1BHU8YrieTAFkzajlXnxAmlcEmE8EMPbC9YDM1b4
je5icP2oU+w6kZv1AQXbMz6D/W2CGbauzgPWdgkkfmvmBDccleu8Ii56xgnwaONg
aeMjJwucn1JqK+vydfXzojgGx3s4XjaCkpOJC+yON6nZ9ydpca5L1BxsxbP7XMl6
ANElYGOMW/S/vh8Dy5MW7vGDYtQ6dyJMPpn7iQCN2aYSVprQQ54msC0OjEi2Nl7P
n5qoubVIymQtUXLdpkgiNrXCGHyRQo7cikZZ9O/6OtOXQdr34aOqodTMmQfXpNQG
O+Fjugd1xoXyxKgU2uS4YF/kviJITbJ0eY8PxHZ2jRypSkn1R9E0LiJicWHuVyxa
8+7TLWJX1mRu//jjsKYvxGSx3itvUGvb3Tihwq3ERTdNwYwQp5l8YBckflVpqfVL
ZZnherJyqIGucQPdrWuLw05/VB2TMs2DVXvxVpuLRvfRT/jdnbKWTXtduKH2IXWc
C42xcRtG6rCU9Q40YbTSLFqmfGaS6g8Sj9SKxBWR9avu+Mt3w+MGfvT0OrWVFX4c
trgEKyA5Fir5jANu9Hq/H/bEKh6nXqsesLkUmefscTJblI9mOzEwXZGMxSxaCBG/
nBJvQctXhtM2Wyt7VrwUXppy9yZtAPUoRuBBaJitWHXtn8Wx3qbldemXw0Dc7zyd
6FRs+KuzzsrOmXjUkKzNI/Ff7rWcWI6TNwSoATZ1BonHknDhDZWTp/L1MlYqy5qP
K31P6rtQ/H16ZOTs6cqeI+ssx44Q4hOZjTYu7kgbniR2I0uBfTHBBbwKCj/E9kNu
Mg2gvgIipTCKZX64o0/sppLIIgLoW1zRXD3eKHi0LlIIJ0zFJhwl4E4Alo4vbn9w
sadzgAMD+yWEZJUPc3SIeG7ItvB6nkBox1X6u6dbrccvmCOKNjRun5qw57HrubSm
EhrOLvD76f09VTLovcO3xVMi4ybKsSzR1ZPFFyxHliRZWhEuBWu7iZdy23ZExx7J
DtxQBx1Mqx2Co39qpKOv4vlYIYL1cLYoEjwkoT0FoM9vzd5CHzSgDG26yDZ5zX6e
qERMzd0Jr4o3FDiK92IXEJl0Wegcm0v24BX9nMEUoT54kH1v7WTxE4NTqSOGs7+D
AhVWSzACo/UL+BrAtU7jymSDqCS4OZ+13d3O5Af82WgqqVChD5xnkVwPTV3YYcLk
TCa5MXS2JWDNKgV/OpLumDNvKglKB7ig4QwJ0BAVp3LQUWPOBpLFpQbEbQPv+9cO
siP3hiFrwjIl1/kjSwtmEUOJvsnF6MlQlYcc6p2IlDshTjO8Eiq0FxyOfAEjelGZ
EGYIr2QMXT3grNCYf70svy4JBlAad6qnAd85A1O+zqNF5YlGZr5HCcQrQxmE1uAH
CiEOM/hHvykb3sPx4JrnP4UJa/CzU8QyqrFfttpF+5gMy089URmpnyuMLGPubWwW
5sMSk+ANlyDzT6GcuomP9szWZGZUO4KIQxjDClE/R4+vV8PmyzIXClO718HdaSVo
N8hgRutCcvH5ncZnXjvYyWpeeZI2zZCdcFX6G1VkQhP4IxpSacnyjKQBNB1Vje3S
4yXNPHXLyEqpkeTo5xF8kHjh4rRvvm48pYq4IxCtzr+xptWNp5U+9rC8obXWLW7f
xlFgmzOX0p3dSNFggPFrhRjqJaxb4qjnqNv9Kz/Hx6VPcB/TVAWKs6bDTGX2XWXp
c20hPMZ+bqP1b2BHskOIP0lZkq7qrGkNKYrVIjmKtYZYhlACkoyXU+PuDQbiQmWG
/+7RBM47aiun81MrWfQnkeKVwsxeFto0DGVz/SzBtISDv98GCXrv50I2BtS6DzjC
4BkWx4AGFnEBUXtnF7pZ63SPmbu55/41d4DISpbg9dtc+fmpius+9NEEXjn5oU+f
zAOffOxZt45Ld1DkpJ3zuAfOtD0RsuVSJHae4bBpzel7w7ifkQaz/bxrkxMjLHF7
xM0kUlYhJCr5f7nZA+JcHeqLXJyZGFDncMMFUAw228IxEOu7VpVWdt9RVHe5B3RU
k61e8WQtKTsPq2Di+m9/rp9cZeuj71Wge4quj+c6a5pWVtlHBht7ygoxAJ1D6Anu
0YvbmpFBvOtrNcMt/X+P2iJwc+wVgHlzCEiYdfYFw+R3VMJ/r53jCWbBHG4PTtM5
dJ6u6HVp5WZfSnujR76p8hIkk2chzIeKq8utBUjP4M6bpPuIKWO+DYOsjSBhX3It
jc1LtlN07mnhPP52UX63t7ENm3a9bChWsWUKWKyXB6tDy3YPq2F+C2eY0Y0vtHoL
TJsbVZS8ighuBjfWzjcgYUnz2tBmOW+ZdIVUwBaO/BGmx/9prv+lrdyYRNv6JiI6
K7/WwslrnFt3Zzx/qk98CXE1NGk2D/xrIkxnqWuJZASQNHmGm81iHgOWO4JwNV9E
EuYib20jIpLJL5BgC5mB5Xq2eKna0i7AcG+B08VA/HQgFQDj9SKI8xvPdob2Bq0I
ZoEbrm2l8HeSzoAinWjnaW278Mya2nsBiO4m/3Gd5q5yZxX0mC/hUO/BJ2uYm6Ea
z/yxjOkhy5IkerqgnQPF3DdJig7rhZ3k1ivoo+fBJdxKOZHDahW/87qYcBGQclUd
LDFeVuQn2AHehyZ+e4Ylnv5kflFwlBeunF92lCCArYiHjo+tj2BJl/FShKZ9u+iJ
BWcl82aANiwLxd7CE56jWQy9rv4wDuNC2FkCnokja9Dt+6nWPbf9ikdnlcq/mKyJ
hbigITwRwHNf7GaEYtVT0ugAQ75kfm8xRuGAPB2GWu2h4c8TawAGQ0FAln2OUw8P
5cSRXJWFs4MOMu2Ettpx+ZWC4cukq8v3a8QdsNM8iEoTzesSVPN+JV1f+OKGmwTX
b1zaHU4SMq8Qvii49dCD64dl/Rdo5rf9uV56/Ct29gkKTWhM/XvSLB/hQi2qowNf
1FnXU+bP7Ko7pkVs6L1lD2Lp7SlaEcq39oMiL7EK8uY8bGwMEGxa5uRa663iRLrO
lEcaF8P3XgCLoX3sdIEp1ouGNkHI1k4HOXt6zkI+FR8gHOOrT6aOEZxb2WEISYMi
9p7ZrVfQZuvIzx3oLtHFfw==
`protect END_PROTECTED
