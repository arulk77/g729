`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73Cy8m3Cq+m1F8BeRgvpWXQIF6A9SS323LGryhUP26wnWD
tWrwYLtUtSzJA/j3hWEXnCKqk196ARl9TdZUG8FHrV7o6Pp1n601GdapYA/fzaAC
SVlJs8DpKpylxGVQljtQWhmN9Q0d4dr/5T/dRjhTtWGy3Ff7EyT+3DnHk5DU3k6v
6NBNunB3D7ymJbYFVbY9Z2N1qGj2ahHbbJlxsw+Amdw4PXH865tNVB5qT2/I1hsB
7ejok93F7ub0ZUoK4yr/XYyMPz6IqKujMtPghYEAbPSRZEDRg/LNAcVs/lgiXz0c
eBzxeysgw38pnpXJVw+VQ/vgFgeAR44PwnyPX6CL6JPuUwxSRqeYGyn23DlSEP2t
`protect END_PROTECTED
