`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK/y3js9815gOxj2xgAyrvBZ+Ax6w4y+pkw5RjkVmiRU
PXvCgxoPZp0mAzt7t68JnUf5CcU9zgF3qnB+FH2yRWKfey4m5DzUwTlsXXnjp9da
zZ8PxDM/U+aMI7NkSHZ43FxC6vRQGyxk2t1IPvNFLCrpXmFEfK1rJK0Lcm92DgBU
Vcxr88RMqYYtsZJ0QBUUeLlGI85Hp2TmQRkNqgnCc0du1RrfF9tRfIMJTXyS4Lg3
WlrCWzkuNBqAjqYStm8JJO7BAG0w2rnITXLwhqTyrSjjq0IgVuZpmD47vXVKr4/O
+HT8HsPV81RmlVYaBYLB2gDQCestxliOJNY7/KZ7uJrSsMHfaR228Y24T0HvZ13W
OkISlDKRCe1JQidSZJtLmYwNC0W2fLLREpl9MJhfduTPWXkvlgCPPhBuU1QasFWn
RBBnWMI7NVAlLRXACJZyGKSlANBOcbmnMkrq1FaOn24tbO4g35ny4L55SsaIOCOV
GOA8jqzolt3kE7OZtDwP/p5W8VTw9Zh5RJKILpfzsNMXcMFW6yvMdmtluDEbnr5R
1gXjbyBpVX3jakT6Q0y2rAkh/+Ihv3sAbdZthYPm1Q6hWtrFdXquPfbQ+jPUTkKS
yq9LBGQGjeY4QtGKpj9YX1DDpJxZaFEbX3mfQncwVk/A/YDxvd5pyQ78bj8h7J9v
foDD85QD36izPN2Tq6dpjwEicbamCkJGtCnQZuZHDtJcfW7Cy/eZ+8zimj3plrnK
wI3qqa9n7XEQrS4IOCrV5wwRPQCCXDhptj+lbGhjOH2hro+H2DexH6ecQD1zZS/7
ZCpKkFjaNzXhPNA+KzEtsljQXruCylCx4jhqgFJHy7I=
`protect END_PROTECTED
