`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+Y5kGnolFeHhHnckN2QpdkGNofzwonS4TWXieBVJiZ+
w3ldMTp3h5D5nPmGXt2wOUgBZOeUKTQK7RebPGy5/vo11P4ANeUTWExgpSTHbV7r
NM2BdNXClxUv+Qb7rv+siaTtHbsdG0tu8rPUmSbvvbNcjiKVkLI1+rHcAflF3Mrk
HQDT85a5fa2M5gM6a0DhTlCVYbnrDWT4Pk08wF1ZUmJ0QlvITm6Spqr4I8Ur5Zih
gxLQw2ivH5eVxVthSaNSLx1aB4lvUpFmhnTh1rENPK4=
`protect END_PROTECTED
