`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48aP69n1C4pdSGTO6JxW2IuU+0rY+mEvabAkptFkgWs+
s1bg49vDbxppgSefYotnFX7U1k/8NFilo+hu+s303RXU2jS6XC+1U6ZCRUKsDB/L
VMrma3f/N6M/TRB4w1DaEFOsBHOO3GS7fC6WoiNtAeEXUGjq6dAw8lM3ZPZKVI/v
wCL48qS1Q3Ay9CPFGhCsVSh+MFp2SAQ01IhATjusrQfBsk3JxHf5NQ33c3CGuzmW
qsp7twXObS3Qc0wKDlJzb3/FFftIh9l1swGE+ioJ5dw=
`protect END_PROTECTED
