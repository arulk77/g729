`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFs8XM2VZg0cjQQrNpcwtojmX4oq5Ua3d99l6qOBIew4
iOp4RZBGxBHibv00KZXMX6tsUjVnTh7e9Gj9eENj5I+nqZckRZEp7XDWNW9fnoIK
H0W3hUsOcTAfQInJUed4gQE2mnPM4HSCp5l8OgqJ6BBNce6k+QgvQOkgq7NOb/XO
U9mneNtp1buVQFCLyHhsFiyiB5yKTaSCRMxj5LeTz6KFONGAYvlrq4rxDjdnD5pe
rpFn5571i8S/wDccmV7ntkM1DPShC2535LP4JioO3Jk4nwJWeGkahpYjTXPv/1Ti
9Zn6G6pxnn6KOlxn3N/O7K3Q5k2g5kb+nuFwefR24/LqauhKxt++7gENRH41cTbG
o6Djq4mwmSARsNPx3WZmnjzDGAAltv0BSjZsrzWqEBZbk+s0p984BKj4FfUgOFuy
kFnKfS3hnthNR8TRF8uZ9cYYKGKrCwDd79JluwtB4oxdNeZBtlMSRQqp9IXM0M4I
wXABbCw0eNYLNxhAiPzBh+kPbljmhUzPd3pQhYO2b8Ke5IJ445O5SD7SbeR73szA
`protect END_PROTECTED
