`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveE1QTICSeZCOHic36ZIqrIVVNhXKZ89z2rGwqwYdxtJD
I+PlYR0xW/3T/eH1ahpdH5qD+7LpoeYMkjEkS8QV2wATZxRxXQQhryln1Ruqd9Cm
efVgfGK0KcBtwSDBx7778s3t5PRWgyX+MtZj4WukaqCH4A198ryXTFNp+GoFk3aN
+Gc55mEqXCKduG6M9ZvSz9g6IQ6ugiOzWG1YC3qp9e9DhYIaHYDZBlaRfZSIfvRA
EwtCV9UtDGPPX/gd4+TNGWXT0PpDmDFgN+LZ3I7GtZTUiu4IWs6VJX6tYaFzQrWZ
psXQn/NMgmtwIw9IjbEuNhCOABJOBfgELfc9MvrLjX4GLiuBWI3qa5EuLDKFrJ5o
QR9wZIaaXMYF6SMI1q9rv0AD8HAbnCXBtGigLZAOmlUIyDVLVcPEx9vw5dQSiZiR
zmgZU6NIl3S+FrdhJ6gMMjRtXJQIpRSu34ICn3fSC5Hz8vk8/kl2PtcIfdvn6Yng
ZBzPpmQcvzdizLEl9R9YGg+5F/X/cRWquXAe1l3Z4FJgYh7dCMDNqBxlYUUayHQw
kBZM/WFBfS8YLQBCDDsHb89VoeRfiaNQX0KaM4cjEgGt4b6PA0QvGFXOPHUVCYoD
dhqtG7451k+R9MclYLZPgxKtzMmEfqF8gyeIaOkRtrW5pqSVNI52dCFLO1IIrCLY
SIhyUE70/JKIJTia+ZK160cMZfqQ22dz5LUAMwvVDuG97QCjT2TKakK1+f30ZcPK
Q1tL8SxTNfJa1V8LmH+YaWPCQ0ejpPZ+477BsJS69pikpPj/xe/RDSBIT1JbmPXb
7z2RKr6G/IKnSzovHMwZ+Cr+oVC5f1zHZ+RKKKk5z7ClPep9JoqNUiNmDHrO2D84
m35tA7Ip1ZMZ7oZpYdVj6743jiZc2vbyo+aaK6fqikuDuGgBbuJt/JJa+C6VgZav
+TkOrtOpUyoXticK2hRxZDrcrJqmYYo2gMVTGL1VzZZRPpk1W5UlRPzaOE5/JqPY
Bflm/fDygDgC3njoMM76FoBrCfFn8DXmwH5OouUl8tQ99RuBy4pny+13cosiCqJa
ScBLgL48bBQb/+CyfA6cuSQY6bHELWCbdIFf031ySm/C+LijFe/9S83D1a3WJFAk
EPLnkXuwuq129pJ8VDiwjnJAmFYwmrFHQvVXJxld6BURdGvDIDiwFA3/FKkS2+Vd
R/Q6UnDk2Yd3og/vt9e7rJaQURVPaPFBG13i8E334JxCcjLfeudOVyXUX+sBkN+f
FBH2Xa7BZ9VRrfYIvw9z+vaAQbvZ7/+JeHuEZ9O2tc2YRIlO0eKdrnWvSRzIYqqN
KtirYTIXuhXpC/AG+UqT3kBzCyPJPwr3dN7jdxXqDvXTjKr+jQfgtpUoh1rfcQzY
447NKMY8X6Nqf0ULVduzAnN6uvtJ12PjymTEpgD+Pdprme959Y2zTVSIPlnDTwIq
qRp59tOEAKGnLUARWMQD21uLZQjYW4e/JAc73kL5JiIMt9lriukEvf41OrQ/b0Up
53PvUXNFt+XiKF6J6l/CEvCmNVMgVEG1ZfEbWDc/nOLXcjj+gsU1SRRUuiWqc/c+
HzMxPckxfrM3yqiyD3X77M/97D7fUl+m93h/G3X1Qqh7N4F2hQ8uVEnKHSa6/t6o
x8NSC4jMrYBKUN23widiVDVjj6CqW2X9/h/XLr7UM7sy3jo7mNgKcz0+SCBzSVPq
SCjB7p8eOxU6Wl8x8pmO1VoybtnTuzsAV9UnbW26H5b0z5varyaTc9RZk1JDhdVa
JIggS2/uyXBoWf3TPlaCW51lTC7pNYltQ7EUmV3vFZiOaF239NY4aWeswQrih9QF
JX/0yDCfPCAMA0vzONb8qsU9hj0mIVRpMMGYOjJpn/PfN1maThUI01gUD8E3yjRT
6ol2+BjMMZdkxWMPG96IAvX2OMXsMN2dZbx/didXCBtT6wHEZ/Zn4QhKHcjMK6Fh
kPVYA4S91YxP/85lHPPzpLgBI9CNikwXXH4Vaw4JEH442HQQS0l6q/CFqcrw4vZD
KyazGGqOtItcALXGVnV+zEVePOC+btzk8fCnVGc8BtoGTStguZ9/QTQsmeeyXZea
MJt221b36erBhJgd04xpCy+Ey8F+7Th3R03684la2P4ZX8Xgnxsj2QxS51m6oZGh
LGreCUlNfESNQm+YKIiQa4Vl0MfqrXlr1pYem/GcGl8CeSmC2Bqhw1dH8/erfDWY
7sxTEHRgfVoCaS588+XRwxvEY3JWXqjj642fRJubA4sXfLjwtrF6klwFHPxPSNvu
pf9Oyx0xGsEBM1g6nFuHMMSX06iQYqbLnE6P1cTKx3OtUlLGlEvqhwCMfNAyK2DC
b4m5M8jnj/CnggwaNylDwQevGxEBxv7QoPCQDKdRvVBO/lteRfBUeQr3Tcx5IJVw
+4dxdZxU5lI/FdCcPyQ7SJKFVspImM5H9A3xaGkdSNDcgSbBAvvCsHLlxQ42geNo
iXuCqzN8JSZPlZ3RSoSAsVuoly4aFe7IS4r04Ootdkc8X8zBnp1NFHGEdH1tLXhH
QQ4vORe98R5QnoAl/kru5MA371r1X/krzoXpJa3w+5qXdYDkM0vEAkfbBeNt++wK
ZMV6H/d0UKsDdnHKE+Ie4h7brAgoMxQFe8ywMz0CPsZIvmGLAv6cf7k2ziRDuwmU
w6LY+1DnFvX6mC0e13TWo0SoD58clezNt3+WjcNB5RQo21irFmNIfhvDHqSYin6y
8illGVOoE9YjVC05IJehOFUbxzqIfb5UsfMrMBZEYqR1/gZNxvEeqbgJ3Zl23eQp
Oc8xK6eK/WNufgsVlPErp7ixPTwsVT729cyrImfh38/5uHWbcQ+SHUB3FoLOxF+h
qVQkhD7lTMve1G0xlTxY/iCmWxMQdtpC977Kl2SD37/rOpxdbj0O/ejiodoTEaEh
BlWrqz8oojrPJZiGoU+/071BpiPh4+xvWAbrGn/7MQheMaKeYjZhLg1iPlNOflxt
FhCvdYZeEDVzGz/Xm38EzLwV5BgnMBFZZSAZRSrUmXqcJJkpVG3aqxRlTW1ny9Il
V8KS00isQaOOjXzD2xWeuq/78hHAwCrRxrlCx1mJeXHYjN/RghFclwzMVdqMrW3X
sw9OFC/aDx8xPRPLI69u8tidw5l/OdEHZYU0+WlQUz9+Dgy2dX77ZsEMpaejEIz3
xH6tzHMy4YA6d5VQMTHdqI4tqd8zeNlrzQehd4BNgE9YN9clDAk9B0Kj0sNwwl5a
DxMt3yCe6UPyrGC2wftCg4kfhUc/28D/l7kuP54QnlroBeBZv0VbE8snedENsr37
sTxh7xxTLsmAqlP4Ang22Hqfq7aPGiqT/LUQxKf8cyqNaWeOwgLY9DmYt+kYiqzY
OVsuPztnWaDMm0h7iOSUHQ5G3zp1jcJqedRWmiyzPaAE114KPzKhl9VKu3X6IxYn
4xX7fRMeEzni/4DPxm253GsLKqYF4NARFOYL3UQ5/wySUZX0eA70EQFMsebaF/oX
hDf6y7oUJy8llzXkMKsJEvnDkdgoU6Wqkr1Mr1ZDeF2yypa5P6EZG9l+hMA9PK2V
2f0DR4BrGRD42Cg4z6GoczbHIvvHSNAcdS+Qyvp3fbm9TzCbhg8drUGHox15MOcg
o5k3pXvP0UJ+AFNcJexrf5GO/rCgr1/A3ONHhh6Jet6YgVxPHLBs4q2gQJ7E7bV8
6fMZ2jdSx1zzwFbcgkdt/u/MmXWytr5VH527tLXCMMpg/49OWCwB0pAOUP12gk2c
2RJUitc9XdEyZtK9vQoRX5byrlArkn8D7JU6iql7TvnuIG0qN3TrwPA8OPIVBUXv
scpKAwxPsMNX8hphs+42wLg7cb4GsZ7r8mRtKgtsL+zJXRk/mb4rQ6oiEVv56BBO
6pb2C5RRIEQlI59MCjRm6KOco3aizfRdidVUA+eBh7kdj7j7wnMY24tlSifwhJaf
ss2LDZcSlD+YJccReGkwXP+vnS7/2/Ll6BO+40r3axcRXFdh2K8jZogo9krBENob
cYtl2jOWTrZkLHRW9ZOW9VIfJOzOAXuM+uh38vI0aPBv33Gr3PHRjndYsY9PL8yo
CZDpNiipYvwL2jXcHWYnKlWQ5EkXS53iiTIgbZM2ysReZo+DBsWx2c3kUXR5Efbl
rp2+59J8PN1yDSy/7VgaQ9XChbWHmZu5K6Tm+FcM3q8z3VifcoiKALI/F5BgpB4z
plTwyxbQfw3kNwQqaQq1cGVZN7wodErC8OuepP17l0aHUURtaIJUrA5WXZX9Rh/U
4zJSB3yGhBnJdJY0EJaCfUVsoLkcf2fY/FSXJIZsJpGKWDwxLtpmFB9VjSAkI1JZ
qpnKMmc0NuOp569dC2yBO+ocRkvhmUuTGofPwhmmo/zl6n0IhzT8U0GWrvNMwq8n
BEgHh1rzTqZAX/ECobnNyf9oZX6W2SQX5xu2kfCZqQ4FSeXaujzAM97PpHqg5kFJ
eWFqj58iAr2GhBb3CxN3UmNpb7JfluADdDhvCobSK00nZx3ob9QhCtSCpgjhTbp/
yRDfKyoF9sfxp2LDIXF08l6aiukX4qjbqH0wxbdT+lGiMRj3iJ8/3PO4DauQO3I8
v50qfDrp998VsqTFwL+rae+qwaHE7pjoibRjugncbicSEAqmkZMvWyLIB8n2lM5l
Ty1zXLIUrfUQCRGgXw1KbRcaxp689GbnHPCMormH7yChwWJY86n2k/P7k7MEa8NA
BZQPsv9Hn7nY1MYd6Ee95KZCRA7hpRyxnNBv1ktXTB8EplRFG1emxCNcXBFO0quz
YRRyy8hhPLqBbx0fmGAvQm3frU9PTES0dnH9KaTL95n5KQvzbC4Yjes1qbTES1UV
85ojO0gn8ZVu0A+fg4RVQ2Kia1AW9zfQnGoWRJjeLj2bPCQKmeFIQs5VIKPqFUCa
TQhUL/8XOTPDV0lZWZ9E6vc+vTwefHxNt5Ecq59mKVltS5iwebt8JOGlwY9AjfK9
sZ5VYIxQLJg+thkTgoHKFNUnAap0FJYNIUuh4PVTpBmNN72xPWs9hX9HSnagZuyw
QZKLgJPejNxLWS6hxKp4fJLh2YsfSMWSsvTF921ZJgeGbPMzNKONLgaiM3sSqjPg
EKjlg1S7J9tMTw+mEKNMjCJN5yX0x33grVZbWjS7omq6tyRJz34vPJEJi15yjarE
nKYKabQIcMPqkxQrIHwlvSAozRSRk7ERKMFs8S7JLo+cwOAG7uInOlVihC4gn9R8
L0jjh4mMoPILYh7cW4YC7upHmqOPqJxSeX+E29ejMVz7E0qjDmVl/ZVFL2LblJfr
J1YXwGlHHDFYPICOOTE6v9D+uWXbICJHzoHTv0t72yNuy7f6FLNU1//V2D55drf9
Ixeq6REig1CBRdX44k03skboeJasXCUKkxQlPyzqV1cDSThki23kY0sQ0JkIGA6g
9FCVPp/MKTxoKuKmFg/2A8sNmUFQ61zG/IDipeZBuZkX7IBrYm6RjL+8kCmv27zA
vhF6WFYbpXgz32N7IPo5e1KW4c2KcAvVofXYyjOLrUJx47YoWKhINQlErzaozH0m
Q7O3HlyCB7Bzbp8xSTsPFVEMWFCJER6zlUAcCHMbgi30mxpKykroS2KP8rcRBf21
VLf4D8t9WxbkS83Prh1UkLBlfzwUUs63MH+Q0zs1Xd/nRQpzRT90/cu6oEvb07UM
RPXSST/mNGvP3hts/VhivzD+ohluzu5siR3biR+c3N3fbgG9eJhMbSSxPVg7ZzvL
ZWACcG+cJb+SCfaazu+LL04ZDxQpd3JnOAI1WnLxaR2XN02VA0WtYrm8ghXJc/jg
iswtpZfy4YcDoYpHqdGzKi8hgjw+M0IKUs8SL9wU4a/GEg1Lp1q2oElraaCdZl37
G6wXBVsjjM7cunzvbcWv7r5T+TpTj1DFTVtG5QL1/Oi39LIa2lA9Tf7qlCYREGIl
KBlzi+/WBOvCPJbdbhi+Dn4Iu4El18jGdFLd1Hr5lopAJ1ofYCxjeTB56G9PWUEc
k35ukHtYT8AHrG9yjlSSA1wSkXXxLHXYtGYGhlcAr9UvT7+IqrbP73hcJ/flh1nj
izHtSSqmORiJU9g83UGLmQKKCZ6+POv1SQIOFMkPG9Fepm4Qrh+1VWdXPcOO/xse
4GJzUlnfYX5atFeMljnQY2jGT3lXVEuRvJoMbwMvJWML5mRNCJCipUUsjlqUTeTB
hId0JzqBEtQQ5I7gXGLzgBlUqaMGPZJrP0JOG/PImb5JSvbecdKRjZnaPC2GcfLe
oXmqP21YjtZszi4PPWoEz7QHdPcqjtdXtymEmisXLjlop4SCTPRNGTtq+ZZ7Togn
Km7x2sBXjquo7dHgMuevFsyyRojCrvIA4V6W2Te2zc8NJThlCtoOxDCAgIzUidZK
HqqudR6L9kA3aSLaa/9PM+LD34g6X4lv1ad1SCRIWdF3vJj2HUyi/v7YmT8vZME9
XntPWcr45IctyRTrrmrWJfMIcrX10n238KJIFtF8dSH9Mp7y6MeMxPrcXo2B67sq
nEbyLPjCPAXj+RtJO5mSRqkoy79IeykTn2K1YmXtSX37dLkkBUqrILbYX9cxiWY+
02+pgmIsMlc/PW5K1aBq47J2UWZlCq+adTYZSyRNnMU4McsOfI4ba1KqF4VAB4MW
TWYWrXuzqd7fcx9Xvs6PB7xZSLqd4xc1GXiF8EFQVcKU0m8K8UmW0i7Xbp/R6Ebe
J13qARZBWsFglbi2IwsnOSMlfOXw/FNlJzC6484V0eBxemq9aIzjUAz2HNt44q5k
bzZTEAMwk60TAz4Z6jt7knZK2X3P80FhKM7eNgcztMASyuHjY6jC1hVoZV84SVFy
5EL9UmkGWJ0YTSp7maeRCqXPxrPJgPMBQeQ8r5UuUpirVkRqdhjsdBQYmygLQFcG
uQeRIeYWXscZxVpEZbhimB23ev6GbjstFH9yLAI+OcXH5rx2PKNRG7Rwk74EFbts
Nkbx63s6Lz/ImJLGhhClcvlqYR/aDbl1FPG8DyOEFFD3zL+wULHgctipM0iI+gc1
pqe5u3aLB5JenIR/k+A+e/8p72PCeSSeXL1eU5ckK8QDrKT9J3QpZYgsxgQkAqZE
aEHh4y2xcK7OBe+V2+GaDYxiKvzmptewJwQlzsNuU5bCQ7fA5tlcQCe3ytKeTPL6
PvEuZ5h8qLDSPATPMT7xptA75am0wCSeJT3zkQDeaijGn4azQ0F10XGBmM92XeLV
24PUuvUdgfvLSs6vBjcURDxN2QYCyonBffdPsmOxOi5p260kxgO5vmzqyxey4rdx
+OdywI2mEAUr3U2PctweppqSpU69YZGhpnEr2W2eE7RD97pGpFgSIZCrbA0B61eC
ACJ64NA8NGfk3tuSDVXmYtKUrJdG5e1t5wu3/hLXfFL8z/FP34CHVweMi+GMLM5G
YjkwrBrnniJDMCe6RYhReT3vtySL2RXKzmfnw39FSTmVLND7qz/9t+mUnb9tctn9
/yV4pGT0RJOEbrr7wAka2bLyLqGexzikgqxbZul+zMk1PfrTzKWgJJ5cPS+gOJRQ
v3pu64+VRQBV95Romcidxiwtj+0Z4/7G6o1O6faRrlvhM4jNhyZsrDqvQYIQNC6e
CqoO/HWxU8SdWEEDzNoH0eH+bNSdXSrOB2W9hArjwAWLU46QUYbwMw1hQ4/OzEcw
uadwamnCi2McCRY0pDGAsDz2XVXzVCXrlkadzCdnkSSdZRGhEnGXOo95+jAPWG23
actqPJ7akhehGTGvzaM+KgqczdAyxNnPvLn/oZp7eC+TX/N/alfczdKL278jVJuR
dbCRp9948AjplIPTykZMZqJ5udtwEsA7sQH2iP17DjhUlTRoP1339DMA1aGejr6i
RvW5hBktSdOP52T1voTO5z9U4mGkTRjq8/E2g/9Dzbyut4j6CU6ax8tGSvBPQi4d
vrsP7LUs1WymTG3GqHe3VT5jjPyfovWaLiAFbbeb+Gg85nynQLLnGffD4u056Df4
7lcMAwueOKFmE0EHcJXLTnoLISWY4vafMavr6YbKYz0ni9AASao8ld50Pze4c5f3
wFkNjkPS/L3gEcVJoFzb9Q2fsRoi+3n6IdZAAWxAkL15F4PkBqgryJ1BC1QiZaEB
2TODx5UDHCp5r5szqcq36acGXJpU2TdE+1Zr4hIX+jIA2x39FHF7Gbw63n6sGugR
bWvYifkW+CNNTLc4nOZlOqMP8PLbGdaqi/9t3hYJkIJCEhjX7B/M5p7oEZTAd2X5
PYg3RwJ52olCLF+gi57jOgMSuVJf+QlYG7YwNI+X/bhBs7yVr8BPWQjLV5vngBQL
9fyzZ7uV5YtL+7E1euaZP69TYBde7oc+PKalnPceE9ePnwCaOVyWVCAlvlWmYWwy
f5T1ba8LosGaNXVNUQsPF5M2hD8Y9HrVo9ogay8NrcMUfy62VdnoXGGsL19sLV/Z
z1yzv7R32Wnt4vEDtrCBRH46C3lRMSgR/m4fphcBk9P+MKHwqwNqx3Y8Yv6x7QOG
FJoq3o7CAV/fYdOTIsPrunftYDlK74HR6ZIkQbYOTDiDuCokuHrIDRnMmuhVF9FG
mG0PDUSr2g4RqxaRp8oRo6/xIcopzxcUfzpvAgdzcdqoEWx9nGB/lGG5LsJb0vWS
4AKGuh7H3zNFfeKcrUd23te01BfT9wm8/dpammZoJk08sNMn7L8FB8VrXRHigwLO
O7sdEGMxmDE+nMn8qONo/pWk8qo+fGj5j5S+Mah2oN8J7ZUh3MHTbgzU0OagpCC8
YBM08jxo33uPElSwrCHk+J2bs9oP1KFOZzdfs5njbPv3Syik46/D/caTkr0dynYk
mUUpseZBO88tsA9mTaPqb3C6LNoaASosROYvWyi/rpMr1DFAzoRfxi0REqVoro5M
gTqvDQCutEPnzbjkm5SX7KS/L5ZkWAI5bzSuGeGnWdHBeTUEulmwsrW40MPN9edv
O470TVGhfUtXiOKi5mNLIBgkQWHaUZqjTEtx0xCQQ/AoX7jjCHtI/2k7bEcyqcWh
q4jSvijbZlRVdcgOidCmZWk6rm3xZ9LCnHRgPG/cGuYrUAOOLUO7wM9ixHMd5I7K
n49qwFMh5u/UaEFC6TxdVYP9vKui4hV++assE61sGYg/coELT85hfxon7vYj0TdK
e4d3uwsw6h/Fu5N0SshmrP8rgTJeanqogNNsoedp3vxUCEeB0cY4ugA6moQlL+kZ
MDdBYnbp5LOdo4pFhkgRawJ2cOrX7l/oQzzj23ruiZpxGZ5jjX5aeTFHQsW+flc4
HK9prZVr9AbXYYdUnVsbzba+8dWuSbgRrurJwmrC4Z60xGf1j9UB34IoNnOJT7fs
QmFx6mylhB7Zd+16UDOH1OLOC2lEpftspPRp28T2b1DV+v7RZVDAzQJF3LM5GJsz
K2eeG44RTuQprfYYi4oetaDIerC+JK47vjF+xbRbaSupHs572iWCNb8K3RM23tqh
ASw0TD4AKxP5arUkCMDxA0i0csekPl9KBOfKJEAwDZUmD9NhWR4ag1ORD/j65QvL
v7ArAubo7mIV3wdTbH7pZv3SX9g9/Ynm+thAXlwzKC2iRGy45oaTrKaq3H1eILaQ
izcuvb4Sla65aw8y8kxecoszveQxvaNN0e+pWeK8UITI6Uw2Izdhj60ytMSFMelj
N4jqXnLChVq7HBM5dWOBwDE23Y7AZugxdfBc4qxVOTw0PwJe7Ad37OnNudzTWtXk
0p2Xv1Rp9e3U8WRGj/Zm10qVGVE52l+Ex/qKfUfIC7vtjA8AOavSL1YScxNADAxa
J5NJIcKHcuFprhHIe7Gg/aoupiPtvCgIvRctP7gfW2Eu0sxmAuYiQywmIS5uqsHh
/ZzhLsZn3AhBw0xy6Nz+zOlBC5aRvR5dIHscb5l0SZW6pdEd/HgydNlMDZZBReC4
uhDqzNOShrLsnFU3udQM6vI+jOj3eTRdIMkJRcsqS7rO1apnHRoGQ5G530iTLzy1
OplD57dlAKIw3hDCqQAnF91TQtywmSdJrXmjkMMYUWPwWf00i+OOoyZyGgKVuFH3
XKQaLK1vfCbCQTaGdZKeyfCq66XFFVqI+zVWjVj2eF3RRg+Cmt8dJKMfwW1+GTmm
j+e58vQuLI/0KOAoBNot563eiAh0G5NhqwQmLN5dDk4FZRRZEAtxqvEXeA9jjGlE
3ayYoE/kUaJvfSPTx96QjxKydMB4gK0fMyhbvFT44MOVAracqyrPhzLRr2x7TdOY
sizmzDe0lhTmUGSPOh+DOmSF1btnoUk+3oDt/ukga+iLMkcnGC850TpjDf8pnYbN
jaOjb9cR8pQwiLYrKtvuFnLJHQ1zmvukK3rV5Hym1ajwyuGDX0kiJyjBZhnAQ+lG
z1ZzvFaKeE3YjEtvcuy2KuUMFbmGvWM0XHdJnWal3YyjEdSVGn1eb37PXCPYFMCm
NSpIZSNp8u5bZrioKtLmtyLr/dBKKQ0GKEcHLibEc1dzjslPoqFYifRaUCgmNJBL
rkpLFK7pIF6lLXtslCxrPf5PDUQDQNyCOxFPN8yUxcjGxt0tkOquB7XtSMW1o1qs
lZoy+oDPBBK9GMoxIKnFAJnXJVV2fkeHizJiFb7uD3A2ZHOrs8Po8OU0ZUFmTEPj
4yoG7KFrMRlO/2yfSda6Q4zxpOZvQzDj28Mj5szcT4Leh61PumH2W1d9IPInu+MG
TkVUpmflZLtJQOE2mJjSJYOQANrUbPuVr4UINKAUayR1u26jFDLNyvd511PjXQ6Q
LnGQwyfPW2m1+Z9WnZTCXFiBtKRKxFJ6JGj1+Fh67ChnwnpMuRdI8+rNTzTrluLw
GGyeEuooNWaDgA6c50hSJ5yQjMvCUKC4JvRcn0i862x4rq+aPy6WwLVotOoHzgB0
KP1WDKt3Da4BDxhNNFDdcnqcgvS93xdLR1cKV8b6Lkhfw09tY8mq6h5fClf2tNo5
TyXN+YqZui87Jx4TFnOH7rSCO+dLBNNgc799deeUUrig3TqZrV9sStbFoSEYi4jF
i6+Wc/IUOt8rm/gaHn1Q8vNlJmbKPAeg42HKZyT0/I5X0xwZztqbf53NeHAlqcqo
bOMxxlI8OfGgYnaqALrACSwQZrgua7F9U37TVUsNZTTu1pBWcAnr4M6WxyFBpgys
+2YHYnVt2atIpu7upLUz56src8H45tB+CwZKQlNvKR4WTwoHGbNTUJWT20JXhCMN
INJG6Nt5aSXW9k5kzIO3NEVRZx0aVIUd/pWlO31FFXmHBobTgNAN5hvnBuX/t+XL
g12/b6huNwcVnMmdUy8HtXHepfnaUd3xqiXeUBkn3wE1Aky/aA/ZZjzlLVHVijBA
5S4st2xW1uRFwEgzuQU+6rUdvvFes4pPf/ze8yXoVFy/RULjkUTz0eE8VTrSrEgD
zXb2fo+q1YWB7tlYOP/EVNV3FiKHjEjM5BdntG0ob4O3piYaZ8U7xGnocPLxlYG2
4PTYCANnQyFweLvkOERDW6hMToulAjqxAEuRkBWVXdXOsmnBDaCUpwIJ77hX6F85
aDFYqF9OQWZ+yhfVAl2mGegReTJ0goxOH3iaOyakyn8AuNG33unOzC9w0n93iNW0
JOp2DgjrithnWDBqaCS8TiGjslQHy2E1sXrcr8hFrgWdQzbKrzPl/4gk9lUD4FIK
zHlkfsKqMmGvyg/SL6MhesYoqoJv9igAxSwxHLU2AnSONQUkuJZu8l51migb6/zQ
kfGOYcslb2SRW/8pc5xmGH0Ml7FBOLv8xSvPAdvYBacVHZGMmbe/ZGB4y4fj2BE3
rechZ3y7zzYp4PvLGnMA5fPnNzt/BhiF3gpqkZIm/DlBvkM3SCThEFvcXSfNhWOc
ku1iQ7dOiJMH2xOreTF+B3akKaO+x5cJW2O3VB21JZWr7O47WG/QJ0ZxvPFj9Bnj
kQXjkOVlCCsPSkqRvrpuH6iRCF2R/tGTe1i6Cos04Uqp0IsJZ4bwO/4aD2E7Z60A
dix5mCRrpA02H6Fq9DAOXBMl3dB5rc5FQvTclkmB5GA4uljAOXXQVQ96Nb6VUHwK
+2Ze/YEcD2mXC3B7J9Ar15iq0+G2tbxer31NUYgo91H+A0jetv3OGDnCjdBVvRqB
/TzntzUBslyFdFyXFMRnTA45di5G4Be8nBhG7bvqCnyd06M6+2BdiSjuG8GW5Zbb
hv2huceLROcjAcyPB7Xn6WuPKkSNbQbIix7LLyjv66Xsxs6vkrddLHkgjBSpnDKS
bf8qBb80ZCdpuIQbtvYWqe8hiUrauvftshz+PvltV0eWAjC8s9j+HvkH5GYNUL0w
cjMrQI9KOTT+9d+LNqq+e6BSpWqHDUOPqnq0/jbX69I/8/FGV7tjEnwOgxTJp0Lq
C/95jxpIG5yFsXDk1iYyGlXStGDOaBAiW6PJkZuDokEhW5YZEhI6ss9Eh0OMa7mb
sj9p7bLs8FFIJjYQ3xjzIANkfJfsQxjMwUZ0cwh3VRp/KoPjUQcI+AHRvUrlxWK2
ZqkSjxgozX/LWs5FTHvJyYP6fcYn0wQTBdCfscdfGfa2v/d0L+ZZYCgZqW1EFvvM
iCMxcvwSKt6VIaJJMUGsxKaScKIoQulHoeIfR/ob329FyUHw6/LPaguFfpWTud9q
ZBlZq9YRa7wxxayY5m1Jn7gAl/o2CzyffAslVg8CTQGH/PCCi3jdCRFLfTRs5MK2
pSPpc1W8mpgW0HJLaAMB6x9vPObl+OOYaTQpCqJe5Go1d51yzSpLAOfn7wm+Z1TJ
VBaa26D85vmwHteC+eK/Wc4yx2hakzK1+NGWYXbnb6Sq3rtKGubNqdCalALog586
egLoDMX9FWWmVerBL9Tj38huftLQ14eSlp83lyOsf7i6Kj0X1C+pPPUUZRfFrgBi
eiSdfzgqsho0rBtpbzTldMROmtl2yQ2IqPcN/NAX04DbvY0X6xtL6iZjXI4SnUqE
49ekQexUUTjkYVPTb9Hidh2DbgzhFzNpv1jc7JIuuET/wFEUMGAm1bzoRXTe1/cx
WjhIQOJ76e5GbMqYqHhHduw//cTw25rj051W1bSwlIbFjuZ2caRtojQ2vaVjVfyu
fGuNOEXucISCa5usQvFZzcL7oJur9G3zMG4hoCOiTqiB0+Sj6b10m3/MIH7KBwPb
VvQ3kA2UKhnWzpp7iB4ELDQP1LtWF60IWLX0e/19OTUX5ppDr3IZbL2VcRQaLn+F
PKt1Ege8EN9xBAM1w34IAEetmsyzpd4VXUbigtsnpO1ehp2RPiYokothyMaSgdFm
Kctc1c/kwCgx2CRcNSXmhOidz63HIbWaS2+F8ygpDSA=
`protect END_PROTECTED
