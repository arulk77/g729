`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aTvavKgShYNp2cL2yIlWp6QxdgHixBwT3ehaWVkhMQMA
MacsNp1QH35FsaBa2r0MOJ1EDOfHElr5Oc6zdRNhRFkVV2/PbDIBLrThIb+E6lx+
4YcUdC1rUoc/Ah4uwLnNCPlLV0OLMTpIKqJfVOMuvGum/ahq8PT3Zzrd0xGMbkOg
H1yaRRtR/Ybof8n9gZzQQz9bv1rRT7WsAm63zOjUPk+/LdVjQVvOpmifh0chpexs
vSUwz7/bGMS+kYLxgo8PXfMo4KFoMcgwBAH6d6bbUmuAb32Do/ZI5LPJNlPqRTVF
OY41CHOwijJiCH1L90KPACrGdYVIcwgdqaM2y4MPMuyJ4yuhlw6DmLi0dxtrmT/b
mGlqY+Zwx9QJ9RYldsHc39DJQM+9pZAujRPzW6XFMUruCUJe+TBtVbomJcXxUTvo
kO9JSO+oT7onKi60EljJIHSXMLITRDGQ5vpNRrpzsR6c9kDqscgD4S277WCE03KV
d4uG0qMLqJLMBBgS/Zy+3gTrbsEYpFSrV+lAgDf6qu83dz7VkKXSvtFGTpknhMvb
xqd7AQeIaZSr2swd9euWkhi01FzFHM97HlZGUUK+lEjkKXAoX43HWui3zUpmt2Je
AMgLDE1VwHgeuNtZooW0L2/JrfPwWQjyJVLQNRBiVX/GoahU0VYHaQtgsvT9Puh6
0srvCwDbiZ8LwerEcrIB0cM3q5m86dCz3qCkQa32YbdlfP4Tk7vT59ZCL6V2YHwP
EMpgwS36JGZIolvXDGJR6oKweoQdiONee5ceYDkY3S+73CWHy0qd56IrZperjVnR
jorgiUDDrDXy0WrduLdwfh1enVuy9X6DIl6wVm4OVSypojQTVmQBXgRqyce42lVN
RcugSjGwDJJt/6daBLPkm8xwwWIHzPZS+gu4vkQBB1mOT1vWpjidotuIQNdGhsD3
puxwNLdDXY5RVv4/YHCsTg9PM3gnJl1QF5m4bMypgVSsKAGueFQgaefEwOqcC7Ap
UPI70xEe7YLV/B9aO2wipdbPhY0wf9yMo2yFZWvbokjQmtp3xvdX59ByypvgBb0u
7vvRfnbsZTWX0Cg83GHSnoaKC2IJW4DVPJcXVnZa/3mIL9TNQ2mjh+Af90ca/4d4
M2NsLTSa6J9Col7kJR/l2vP5CfocsC8HGqxX8cnm+f6A2nPehRCLdcrWAmiIpGOy
Gr1hpVxHAVLYipRmL0Z4IDPXX8F5lnDPQM+2gskr+Jm8/WxA2k1ONSHM6pP33ca5
OtrFikP3L+M6DCK7H1UGnmDE+folwxQ1GRomqolMonfHdslUbavUtARtslyJEMtr
TbtPdCz2vTtUe92tymUZWra/BgeG94D3IJmAqx0WICnp3Zo/4C9ZYqGCB5FIJI1R
mID/tw/J1VMhxTR3os8koVFI+HSU22CMrdpVbV2iotH00ijoRnLcY4MfN26qd1zF
HF/dO0DWuNnwSAUT3XaWnz7f98z4iBLOCCf1YG6qRWT5qczYY6/zFBjY9xgto+Ya
Xvih9rioeLmqu/OPdPDbJgHcuTOZVZPfX3JGbkMwNrheuKtBbs1m+lkRs9zbxFgL
fybwn3bWjv41GTvEbJZXqX6I65/G7NP8qzf0tVwNz+WYoGz/bKvswrFyNijrdh9e
lEGzjGL+Z2G66A2v/HTsFrlnXtoJueYOgxwzFMUNJ22fan50mlHXqWAQ6ltI9M8+
R591Nh4Az89qnVD3rtpNYWeqvKhQz/Pw7+NcwcQjNSx+ySi1T888/Ln4iaabNN1C
AALRg+aS5vJkYPtuU7Eyz3xnEjM1yK2/Z2/S4tE9glH8G80mFFeUngjLb4a8pyeD
C8enL5vE1nFrnh1JxBDq+y91Wp1lAqD15JmJI2SrBhbuPRs6L7ne0JFDWvJ8KPER
SG5dib1ce8KAKEaCSic1qfrrtf7CVZQfBdJz78sC8qpYSDuzVd6EQmnaE4+E68tb
N5oHS7s9ru1h89VCzJu30+ASLUiQM1elJW83w6GJ37KjUX9/e1C7O8YN6+7paKEY
rW6z0qNtg9o2JcgNnbCk6Z35JqjW4eLCPQHca65OWIez3wdnUnL0xqF0pmxtCc7J
GjYVPTXPp/hSruXToIK3nOD6T10YRYcM+dthNBz7Wf7Bw29jbk83tcD0I3yVm92t
yN6M7Z04MJ0rT/T/XHUYZ+DhZNRIyaXe8TKAKXRVjW9mtpbKsBD9jXWko1qxGs+j
u2xYG/J7c9bya8sE5XdRcHUf9o80cygdEY7GYFDRh5tiQ1smohTCj9aralzaR/RN
0XSygeXHZ0m0rfUUuaEs/s4qK8EUBBWkIp+dNSQlu4WFO7SEHdv/9lls3Q6EXOGN
/VqDzrYF/1ZlXmxGPbeqObrKZtPSERlR3am5RCv/FUTCKPSSr6+90JIrYOHcuDVO
0ts+ocCpRbEllREctsgLE0XOAoInF84lji/ZpXkW+CiZLMRIoNMkA++0o6nSAfHQ
I4pL2zlNDqfKPXR+8NFFZHuIScbplpIfFpRWxW/GA+5FEy3vhEbQv4JQtzV9yGl9
nZEYp7wawpbUK2BhVfuTOhEGtnRbm2jJlQNVzF5Hku9hz8Ssca1pfAp9k9/bDX9s
m7No0Zbi/YMpk47+MdQl9U3u7bv2JNAHQAisy0fDLhwySb9RPv/Ez4QQ6p59616r
xyIIAKskeWLR05EBEcuaWjwksz6lTS8E2n+j0DzNsPxj457VFFNN5wVzwa8/K5ou
LiN/P8+e/6Q9JW2RzvBAulVhE66vOhPUyfsgd0i/lftfwFWrE1Fu3g80w7uZwXZl
2Hg90yA9Wc5TU05cgLK2bJLk32a4wosoOZou5Ybmk5uXn8ol9UyOTrNZRgYYyZgb
guOAw7YWdBP30W4khfUR6PqHFp+U+4iOerZ3fS+Gy0gcwGiayjcEJwZcWmscv9QG
P/8PqMgmuAHeopZdneBe4gxWJgidJSqD57ym/hfz787UaWcW1M7W+Nj8ud/l/3Eo
vtTVRdP2oAPpdpYnmGxaY26xXEogvhTy085MrerSpzw98RtCP2XtjX7IMnNFWo6g
kgIuZKdFTdst6TMalSy1Tis3hxJWAVygCkEKhBa2ag5r2/5w7/Yt0sLMKehLg7+a
lhbhGLkMpIbcKDexG0NyON8d69YU8yuW221i5tWMTFbbpP0rOJwSjsYGzMcjjhs5
OboBFM4pvSRzIarH1oADEyKBaWb9lH4p2ureNiQzZXat1GW8J9BgnYEC/ENQOVZV
MMys71g0qaU+L/GfmREizrnRGEE1DFo+Lc1ErVe0oiFGeDtHlWxHiFyrcv+YZ3Nf
yfs52Ls+bkjjOVV58+UAqbkTfun4nWvqcCiM5eSeoa/0csS8JTf4m0w5GhCWOJk6
sOXPBaFZCcH0y54rGvMFBfOooXShJrf0sdzRwcXOjFynepnN/4uJuEkwJE6TNrcN
Mekz52KKN/kBeEGykD4KXgIDjfeSDHfTyAvtBqboygw68/2wNj0iropRZQjOecaW
fgCW8dNvJGvNv4Z2G/Q6R3KK2zY+GgAQsNWTOKZcQdRNk0niPeg8hJAHFCbw6AoK
Zbe+NOpXrCa+rf/BDTZTNQ/nl8OtpkIaQz5uph/voph0GYGMdZFcnPR9nOzbNyRz
HcyrtvzKh2s+MuQ9MSJyVn9R1WQUxnOzxwlzXyKB/z36SxmrAdvzH7HHts7bHJYt
gf99gZpHfl3SACxvCQ3XCRbylgQ/Wx4hAnv7utytnrTOBM+0y5R7kGGEws3bJjuJ
QEVgXdM/RTYzLPgQGwEHYdYaFGyIJUg4keuL4mVcYvV/FwHsOcrdCPxFwt+cBw3J
CqPoAbfAhNuDf7s/AsBtGMTX0mwww6DTeAkzSLMpef2b2u0APZiY+EJxlG8Yq689
y2qq/BnZFjoKD5a/OayPNPIJTgiSSdi9JawzsqD82F02AfQidoXwrU8K1/o2ODE4
OZG1Y58Dn3o3r0YDvD+W1/kRwIOsC4XZR2xc/cDQLA02bYGGOhLh1Mi8/3lrHJNP
PoTmMLMvTn0yBxBxWW0PxCtz9Vbd5yx742JzR3tQKStnWsJSxMAznCsbbrjcmPbB
bP75jHC9jXLVRDhBCJDCLu41AdW/a7eBgWw0LXkz60wFJDxNNjF30dExwAr4p00o
8SY1g5sX+ft2qEFQUrPS1LCT4CpqHiVJrqYXWvd4gOO8KboKD/Z8g4Pz8F6aqtSo
b2/FWuII02gJ3pKKe0Bj4eQNpYFYc9CJCbS1atWHCT81ma7FYv3PN0j5ofT0rCOS
ix1Bms/LltCfrzURxpf4JjMc7oMmSfCO7qMbJqA1QERNIrAsU8jtPXclZCGgPWpf
QnBOH5D8dWYMwDSowSkNAr/dgfndBs/N0Vex9EhMAZVoKtfPPG1+I7m2Uvpl+YR+
cCe5Z7HfT/u9UZ/j0kmykBWsZWIAfRfb2OE1Lrn3EbQE3wvB1RRCEw2NADYr3bqO
2YVVdljxyBg7Fs+J0fqOWme3hnMfag43XWMfu5AhjtBL1cpPo30fDtqxGuTFJXRM
cp3MM4nqBbdZ0cssfD56qXAHyfkDH1ugm+jX7ox6hQfQ4xn1ih4/NxxK/ziFA2js
FJ+BaEqK6NS4cOZBvTsZDwiGIwIVfGO0Thssf2VIZ5wvZhMgBrCpamxts0Ata7AJ
rM/PfyM1AGu1697/fJL6jFx7m3tHtZc+EbO4j3buI57807eoP1zxje+82ebtBX30
0QPLODkANYF9fP7c7Ik8mbt9sj2JkU6a/sXs1rzqN6df4vsYBiy5fi9Kon6CX3Gj
8EKEr/JVA512UEDMaj3nV12Igv7I1ZptmVm20yex5pOmFiH+tD8DFSyx925mw9Gk
uW2QxbGj0Ci+PIFsidilDPMswDVCLBQG6Lr50eYJUxTdED4zSwBINWryA5a8c1Ic
W29uwpBCYa+N/dFTotzyqHYyjKJwcI8b132MFBD4voHsFWH+GuyNUKgCrkP/KsfN
Bzv3MflIxHD9CAwP/tx1z/oC/otIieGd4a/tVCiVhT6i0VGABUwEHVT2O2i2IBqc
N3IiGW+w25feWZcfN4LAw78L3ZQdf4atrLxcwp7JC13XaSGILRLOICKLVQ9QvBT5
MTc/lawvWO3W6pEF2aLLhaKNSEXx1rxA+TYI/m+5XhBtImOsBD37sMz498zTpryj
RU7BBAUH5+g0L5Pd3H9AQl55J1Q8rt+G6Vi6axt/YzW+yvy0JXpaYYSSbJU672/3
hEmElH44ssu13FcVN/yb39EKUFINXvMvFwHh6WkgED2DyXzlVUkzGWiSRPv7zM4l
0RDobiuLkNgWoXubgjaAs/p3RxBKvdW6n2k9AJFbVikcfqsq0hVRLaRNq+6qG7hK
5mzNE0eFVfWKvqkjWHpFm6Mj5hprJAW3Ka0FNWIT2JQBP6oxtJ+XMJnPMk/+r+mS
AKfAmokHvE6/NxOZ/CwKPg==
`protect END_PROTECTED
