`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN04wzliuElNGm/HffLyOHUD5KbJjfQH0jF+P9k5wdWQ7
dtMI75wBMHTQ8uHeGJo+MoUmF4R/qNXUgguBtIzpFibFcg1C+chHSALlJN15aLdF
igkY+GSoYxx6UzUju4V8ouaOgcxRlS/Rpd3iH/Dw7gmMWxTU/PATJKzysYPwC/4N
Hgm9I0CmjdgfXP9RL6TGKOpUe7V/wPP7BoOs3rZRUmeSgRaUATS44ozWxYyyBacq
uIgCJrdxPC6xOmnnS2VrVciAiI0+u/LU8TEehUR4SWmGHqw/iGDcf3WJwkA0D2IQ
okr82cbifMLsMe+Bq4BpXiZsLZn12QELHtjrRZH+L7arEW8DgjaTdT7y0T1QGh83
znYOIIHAq/e3RCz4aoMANz1ZoTGu4EuimKco+ltsTEJaFBBIqc35X7El3eiFqqbQ
U/C/DtaqtehfW+u84X6HhrAVgT9s7M/8f4Xsk8VBvtZ63Xx65fYqLzDiUt0LmipV
zJM03mUB2bOo8C+E0kJOEXlZ+hO99eaB8N+VfBUgIWD/2x+U04qqMKZq9rVcayeH
+LJ9jb220mcUTx9420zCr13S51ldA8amuQUiPiG4hBU6DMR3MW/MM8WhIDuKJM9Y
cD6v+nPYtuHOAF8iq+Uo6IVhnRpgVkxAhPuq8W8vCs0MLra/mdiEXVckppCeo6KF
oy4SkgRRbbDuwk7a/ETgv/lezr2GvFhPEYXrIz4QaOzx4NADG54KmYFVDq2+i+5g
6kS54y9RqtmCEXVUWPX75Rr55v0NhqVnd5AtmeXULemdnFDW5Bg0DjpCUNxqlUG5
8eAoirl+HmYeN/b/delE88rWiCFHIFLSCOY9cnPYq/7eK+s/1CLGNqLnc3n4P6IE
dubETrAApkStwIRcoo/K3AfmPDKzvhmC18p/wyA3TZwvtDi32Xt8VjVO5xLnjoMa
efD3zQbeYiRboyLI+PR/ZDif4AIM9igZuIvMES2kRGVUXT/Rujh6u4n7USHJoMBf
/idwEHZbgeFI7u8pSsVKMFn4FPyW5/ePNh6iETvlql94RjsvB2aB6DoRoGfEUgac
eEaDFffgp1O4Y7RdLNDKaCQByNEPCcbXNzapkOi0oOdpIvnH4uuFsehnjqybEJsZ
9qnec/SaqDKS6mrAdzqLxkq/5MMrtRRxg+CBdvOGFyUqRpt8MGkvAyk57kzNo1zH
TDOI0T46T2dORiD+CXNFNu89J9iXOOOwxMXHHdXPCmFEAovbMnjddNequpEr5qBS
nBYDAzcYyq4aeY99ZSYiPb50DjY1uLaHtJjkOEerve8wCbjKrP6w6eXYcUuvOOd8
9YW7XQzF1pdHLIt5TYqKuJqSC6+j72mHxltCV8fV09/gwbSsRuin7RxySuQcDEwg
EX4NCfoPCtg5Lz3LbmF1h+Imm6fNlGKQt8rCjHlzOwTRwFUSM3FyB0JvI3p8t7L4
aUC+uDvqfsjn0SFrBa23klAgMYPt0yILTZyNyhUmrX4R0FNxV6L4gugK5qsHzU3l
1To1DNiUSgIIQ1lgAg2O5by5TWzpiFqHNs5IN5zHQb3fzXfLzQsiUTCIMDhPHT4u
nKRENb6tmfMCHrLYGu1xlliPr2SP7rZvtMHNKDr7CiX7kndw4T+4qNu0kI1IpGAx
DnH5FSjO7BbV6pHfG+pWA6kKevFpv6Iw9VjwIGr4ZFHCOXI9SpibPTlyw38+/aDr
ZlAoT4p3TveuMxMGxOPlY073E3DUqY6IA7ppgGgdgqUCKB9tMUwbGwfYA4YCqR+r
khlk0UoyGpOt+R1SOBwWh9VLUnlFpEzy9//LGwei9N1UsWpSFFm22Eo7aAqXIy/x
bbeHoKOVARobYc9JOYaDytqrznc/D2OpX1Acs8XSZd5cPx5Pqs/zdxZasFNYM0uv
VSjGz+nOFyBAHQR4S3yeIkSO7MHg03CJpXAS0ETbtviJeBrpJrK7Z0602hcCsdPs
ohrWqNCavp++ups32j/2DTAJ1lDWKEpoMCV/Te7EzuSZFegOp5YRTYMKh9QUEXMw
ZEbIlYSNwuGGUdQzXMiZpzZ72qxnr68bbb5nSYhVKlP1DXRDlCO5uhOYAlo8wC5j
3KOdEqyYA2Lg7IyiQrtLwxTMX4v6qRXNtI+7SJ7/+gpraDy5geOAoPH+gz8ypY3I
Ncl8i65jUIohx5Wd++X+PxVahbGr8K1Oa4fIImooSZTwYG3Jsxwe4lZCyIcW3Wck
uLuqgqYLmAPvuWOLTZQ2XIwQ3xz/5GNnbX/gTk/wp0dBFMCTAOaloSkv0RzCyNPD
Stp/NQlIEK0aKlfZ4AwPpPTS58REieAxj7AbFxpoiNYCf+NslbzTPwlEVirJ92LL
bmvOLmE5+uGadoAQyOxd7evNttmUqc0CvaZgWTyWqpdEl5i0g1mVlP7TmZ7MhVCx
FeR6n6o50Ov1wv2PRwYinecOpfeifPb3K8jiFFUHxCckjZMQEOloQTxzfnlNsjoI
8B8EvdVPowXcqQy2ixGMxFsIrawfF2+dGWbqP13bck4wUv1RKkB7TM8741JjS3Iy
7S2yyc99hLFp1CWJfEH1Spyedg4qCcNZZf/CxxIZkggSDZj1VgoGpLpcl++rg0BB
4yxMYUifvBPTP/A77GFsG8bU63Q5jl/PJTljbiVtQbs=
`protect END_PROTECTED
