`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
u2DgeFylRlgnOIdx8LKtq5OF10JKGafoHTc2NvYwu9Rhh8d8JG0nX3jRGpJd0aLu
XsHIsYpmPWSP10+6GLj+p5hzFJqwtWImzxkVBjwEGAHZnb2Lkrb7hDDdrcw5TYQn
6oYSibnMqCLHit5Jh5GIZWgOKhsFfch5YJz/J9H7kPbIiWnPTWwOhK7HYqMm4lWB
Gf4D7xlnBey3q6n73pNruPqsZr5NEW61SSGka76EE4YTStQsTuO8HlSA0y+yDpI/
/f4gMQTr2+dqwnXabLI+dofZTqodCMUbgvdMhbtez3ZALR5l7xNaeg3tzABSSJOg
DhUxtkokaKhi4M2kt80Vb5aUStTrxAaztUpgWlDrN8eGrBttc9Iw0aYNXk/ljWFS
7uNnO6S+qj1dWrCCmzCKD8cfdJUudGQ9Feq4He3PTlwvNYzDBZlntzBueFLjR2qV
MTR5HaWQYTTEIQl6DW69lB+IEL5Ci0/SC2qesuufjIZddZrpN+CmhWrXd86BkgGz
67/hsgq4227bvZTN7gkQYlYFsrOwqhLsfz44klnO+2b+Fu7TXBYzRlqKojaLqNqP
Rb1Wb6mIdKW+F00hbzl5Kqv6VzkhMtRDAD/c/VNUqQf9fycBCxGAmRcSam6iGfi0
b8x5PwfOi8Pq/Qi9EOw0poK4DOdia+Hxlfva4aKKYRRQ8ym8Xyy3KncYuEnz+VBH
jLZ50b2fWUl7Cwo8FZ2yb68kmO3jLc1UHEa49qDlN+OLZ5V5ZDw2M0IeEuZTvInF
vhgYTNiPkFeU3ewRDCCFYPqTdhsztLKMzU7ZO9FQPR2N5Qwj/4602HKd82yk6e4d
yg1Ey8n4f1Vsw6BMFY3orjstSYSQFLYZEoMVbNM1YP1FUVktd2z76cXEtFecli57
2wFCfRbMWRSKhV9gmXScTx4f58oXhsq9p2vx8kEZj8WQwQn5GB9p2BsO39eL2dkk
LZJPyg2EL+8aWDnYNdGG35aaOnCDEkBz49DQiT4XMmZV+wq2/c9rce2huRxfxgCf
`protect END_PROTECTED
