`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBTfsUwUGWJq38Qrm/wgoD6WigJtnkJeoZFiFO3f2I9d
8Y8pN58BFXkhaq9cCtA3oByH9u62Hbj8C6cHASRHAAeT7R4Lw4QDzCe2dkoUsFdV
DSS9H8XMbNYN4+R2pohmmZ/K8r54CRD16xr9x/MKgrtN+JL6oeTSW9hxJd0mED1e
/8M9J1j5sEc0+l/snO3BgYVhSwIsdZM98aht135BOjNdDpectQiXtGC89iMb8lK9
FMW4IYsu3IJkCkRQNkcAe6k8Ne2oXLBBHLCninFIf8qNf9I2mQTJslKMncUOVQsk
R1sORcZBVEkHXRQ6L+MgXfkOOvoYUDTGfJAPawqHDDQR0hkXT8uqE6FPA4RiJ2e5
`protect END_PROTECTED
