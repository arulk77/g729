`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aW9JcJY2i4qmHxQnHq0t+UkREtRmMOw4e/YQL7WGJHPR
mT7yEbAdWOhzcCu4t6AJUglG/xcc0qad3+OeqCdqztwfgw3I4xQH8Iw1Z8jkSW8z
zb3AmVPmVbqtIiuHs6MbS16Pt5hJBFhbLuBEeyE11s6bozWq+HYHW0bsOGEPuAqe
10VeNc2jawdK9LN6t7HuZCH2GebBOfKDVDt2El2fyo9nTIzXInbyVWXaWq6B3zZG
ZPghcIX2u9bWudgA0KKzYVPGafi/xcALsh2yblIIW0LxjANrzGcWc5v0jvgIIfg6
8njyfdQvtN1HIZgOVqy7bkDA0RYwVsFH7m3CAylxLNPwtqlbLhvFv+WaZDTciEDa
i7NDw65tb3OSbVUlXkn4i6v8Aq/T9zYgvt+Zz7P3GlyO9TuWLCxrYCV3gyIDFxba
yiOaxistE0T5Mo3pFL5yn2rlQYPHQ4u4z+DDecmCmiYSW1avYzIw+wGIGx9zW62K
TzVFXCEcXTVnFuA/d1mRZiWUKgYVoK1EJvrcL82aR600RjlOr5izhz1SlLyzhz1p
nrragZ1wwxDohLf6KTQl2C6taTXvgTOFI37gO1W0etvaq27u4fPfINZXcVseyJFA
4VXowAcmqMJEvNQ8PstSLqojofZi2HWbgLMHwvfxxFAkYPoLOPIIeocEzof8SLyO
c54cqviB6I89PcYki8RqiINq6uzlbfYCaqw80aKC1BA=
`protect END_PROTECTED
