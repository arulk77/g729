`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
YtO5XTx2dxBXY1r3ZiOQ/qImDZGIuN9thiE5z1UDPidTGxh0UEHDpKxrk1QuSpJ0
3t4JbJlN4MG9hkgoRXeJf5c6SPMTbwCbtPB2cqhC0vIjbC8JA7xlZ/NjPgA+1R7Z
lh5yLNLr5+iEh+4djQbH4Lby4FxfwTeTChauRxwjkxzycJ1Kn8TJ8/OB2OYjTSzK
ggjfBuy/8/M/fCAcXhnoeDEx9v8InqxRYyFGJwtCD8fOYfvytIlKkTNnAPgB2Bpx
KDwgxJTwmLO9qQbG6nj0u4Dt37npeOoMbhRqADgzSJw=
`protect END_PROTECTED
