`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
7RWERbz/SCu29vx1yp3KRO3Ka4PE0vugPWLhThPgps4YikF82YiPRfVc0WpbNfiF
V/oJ3eHeyfb3AWJuFzWZwpxSR4XbZI30MlYn8CtR2R5xbMY74ak7Ukk2K8c6nTiC
FueZoe5RSuGdwZyFmev0MpOx5qddIOKin7bnjI7evz2+j7NRGEEkXw8djU/G0C70
`protect END_PROTECTED
