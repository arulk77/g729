`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4ypPY0Ahkg5IcsFNyutZZZmXFERZA5VXjSdNldx6O1YG
2SS9cagAuIeDf3+3osTzAGjH172HYqEs2s3II5ar2tga8I1nXHDjuBeog71AIMkB
aqwRkjPHw6/efDA89k32lUcrS5jxF0b7aOU5sv+N9208HBgk2MNTRYjrW9KxRFjg
UiPBRZ1mV6D1FQEbUN1VdeIXE13/iGlVArz3kUnoj9q3q1UZeTIoU0eesif9xpss
JZ4rALMrsChNjI+0OaNbKJ+qkmb9wDJdGT0J6cme1o8=
`protect END_PROTECTED
