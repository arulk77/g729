`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEPAZo1hcu0Mia/fyhUpB+PNlQunkklK1S2A+8teUfCw
oxCxMfAozl9SeUcpwM9NXZfWsPzVyS8tVM3C75uTZEOnGYCow2lp398b4N5LANsG
lCHgz2bT26lZf57IULyULrQtG3waHj6rd0Rzgi3AQVQ+KvvPSsZ57+ywoMAF0faG
xznwtDqXW9wRFzax9cP2yZtVjkOOSmIrFvF1FgaZ1Xm/Qe1hIQbiEwpliNdwpQug
6A66hi1Td6NIKdwgUqYYGDgZYg7BtOedFIa6LzuYAMgYLVKkTPYEU1br/jFIkCpE
LLaJXuei1y1SeaWUXihAvUafsOm72SpzGKGNipkQGq2AYzMOP2XVYpWiKn2gkLty
F7YdA5F/1GG5tzAKhS5zLf9qMI9nThp/ZJLo4zoz3T2xdzmrmGnj86nq6d0BoFkI
kOS+4wDpoUT6/fzriF/+QZ0nmUS7GVHwvDo1UoffIoHgxde3944I10FG9eG2WreA
7dKyB0Y+hItOCV7EXKKswV+hoF9S0x4Vhui9h52KMiB0/o+dRfX8L+bMsvOBpfqM
3awTcYfIzuzE9EMLYKN9/jNuHd5IxwH2hCBOLTDec2t2X8kHJ1yB4cjOuMkyiGeA
HEK8NyZxzGIjFN83E5vPq/MhaJ0bi6SUE/eF8SsWoA0gM42m5luC5bQkSDwUAS/x
sD9YOVMrGXzLi8LK1+aPeg==
`protect END_PROTECTED
