`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNmCB4G1hWHKZ7S9eJ35J4KcZGChth4uflDynNUE68yL
Uyq/hCnrJIkYCpoxsWK4AptAEg1M+rmw9pB+GJy9+vcW1GyLt9Kj8Fi5Wv5YjVDR
dJEXgNwjW7/k2Qo5zekhkR33yO7W4tEQKJxgm1uFDffOJrntgrM9G/08/6SaVlix
/WjOu8RCM12LpamFDWwphCZqgizJnkV8a4mNZjG5st+IJaaJywYuHVpKfs1OjUhi
2KGD7qqw9pQEj4kCv2W3FZdifK7ItojLY/RsP2T/nAwXEHEKWwtdHFgZ5YdJHAKD
PLOhDKQJUstNAVLVz/CCW5UMZmMs7tCvJ4fybg2r45hO66kKvBuxtnu9Tv4ozx/X
WbR2ceVpue5iGpl4ETIzzrG7EN4G5pZuGn8FCOaBlF9I1k3SArGRFgsvfhvKoZGN
4kYAa/L/PFMmmaVV+mpjXGOtiNqHn3UokrQ6088J33fgTrG0E6UnjUtXpcOx7pWG
`protect END_PROTECTED
