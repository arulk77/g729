`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C5PZcGVLKhQoRDoC/VcxJsw2/Zm8cV1QTL65xuKhQfIg
0/P44tuYZHEq6cXucgVK7XMtWnFTTeuhmUEWMhm9JjwmLnlrzOQfeh/kS8PtRhc/
yIcZoH3rN9DVEu8NHI3u40sQXoLM3mWOU5x2HkcDDm7jxqMjDzzHRRcD672jKhaG
9OeOcBwx9tnfkvlzaS7ecSb7FXXM0tkoLX9o0GWlNPI=
`protect END_PROTECTED
