`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDlq9/FaApPzoA+QTxoUYNviz0snKpwC6uL9TWSl/Ztf
mQy7ikaStLss5cHX9zk0Rut5aPq6cBLXcG9CFoqjZAvXfcOgdAOfNDk/cEQaeE5m
sY1vBTFDgrI67ic0yR4az9vZdL0oww0JoM07vDrBuzpoAPqiv1MFe5Yt1yQ2M6EF
mpfMPlny7UlzI9HxXL0tEV38LrgbGajoExTlOLXBGx8FH1wNjPHU8yrBxMV9MXDZ
BtlE9hoHcjuOOY7a6FMJJQP9Z8cpFbAIoF4CWREYrjxS21NntX3FLljQCyZGMxK8
mFUY6wD9xrujHpxZfeH9iWM/bLQeSX0QwDPdfnA4kgoimaPgr7qTpZJw/It9Kgbf
pGmFrf3E/+pKlIOG68SWfsxhMXcnI2CX67D9THQV8fojwQWucrXioh79/y8/SceL
vZR2+5JpgBUi19onYRAgoBgRJxqsRK+FwF2z5b9YU3CR7gQ6H3XgcIDOTF3SRGOl
sGQEhvtx9pguJCdhqJkL8cQvX2txSSTxYvaYQdTzwtKybwzS29i3BfyFQFS3ctEV
jEgu53Pd5/CNQb8wYleEe8JGmwNolh6PlOIbQxGSI3+hYDCslR377NURs5ZKec81
H7ORE/kqYm16LMTPGMy0gfw/u7vdmgT2QJjEritXy43hzMFxSuhj7XVdOgb7Z75s
Kcz0m4oKT1Tj/lAWfUN8jBPqoVJv/oRbZ07gM5ZCJsXKd14klfx0bAwKahTKJI9K
5Q29PoqPb9TNfL6EOCGKAA==
`protect END_PROTECTED
