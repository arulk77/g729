`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEeYQzSWJL7cxbPv4gZ0Zh2yng4rtkpvWSt8dwOTuM2Z
eCPP89FC383AE5B3JUHx1HX017+MOxVYZN0a79yAz+eJzOizAdogNY4u++5ycWI/
u2LadZdYaE9SKZ6A0C2rm3+pPx9Ffjf7Ras/cVwWf2g=
`protect END_PROTECTED
