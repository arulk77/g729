`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL83o4JJrU0G8lvczfrmhCX08FYGepoDaU4okJV1IyTZNe
7L9ozCUeCyNkreRSacyp3aa9T1QcyZp3uHYkdifYTbcje1BOfP6wTP3qc8ynvlB9
mC3raDIvo8dALL68Jpo2p8fX0Lt3E6/vu9KnxKFgimkOXmu1s7tQcYsgbR58lVyY
SBmSgUk19UbNGne8iJwOf+JNTd2gqiSOARFrlJDqtdvXamhc4TcjkmjwA4179rJa
wCLvYntQI4qgg8PYzktH8gt48lNHokZAHbG5zMvVYmy6+9+Ww55HYgoH5J7Pj3hL
pvmcxhNX6+fPnp+lS6MzNkPVYAIoxzrfPcgWNYyTY4T/hWpIC3QYI42YxGWWoWWq
HY7pURdq0efnxlFoNPt2y1yiGylqKeLIe8BdYnC1PFH/T+tdqqDFFhJQijuqyj48
Ubim1YXzWkbRnM+VJ0K84itsFXRKYz8N5lVJVZRmi3XZjGgY26Vv6Dwjt4SDWZ6M
`protect END_PROTECTED
