`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
gQrTIifJCCtnjlsXLugpN6U3OSERCmDuPBWdJpGR08rdIT48ngMfV27Ip+0boV2P
F7r4F4tdP5ve01HtIwVCJcXh7ZUwTGqSJz7jFIKU86XYkfZ+lOn+R1y7rj7dQPiX
ivw5V3be39oAglCg9hNsH5sqGqyFlOLTH3r9Bu3OKoo=
`protect END_PROTECTED
