`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
dXi4J+UNGp9P0Sxc5L/xfAZSt3hyLROcQI47jT8JQIsz9me/Jj/gu4dWQRBFPlLP
sxBMzDrDDyJMu3b1inKF+DEyNbObQPvFYTSQsFg6CMNWGfvQLF5P83OjITRZnXJz
fJAtRCSRigFHKh2vuWbjT5SRVUzarbw4sKS2ecu0QKv34/m6dOhf+ViazFEO52Ly
jc0OH9PUkTzRDUlublTp9CoxBDmB1vTeQ3ALftzgC9U2QgG6njTCF3krWlHPeZLr
ydTU+3uN7IAy7LlsIHmtGdbEjp84J8HBscwAPq9PlXk5dMhpek5G1pzD634/603X
pSl8YPnav4Mo+2A+EOk/USkJH7aarjtLVmz7LmmNOViofa8oi5oX7Y5+ZJ/Sq3KN
KEaR9LaJtoBiZJkGoYJBtN1DSeqJ73BWnkWnYNNNr6vy6VM8DqvUXIE1Z4957wzj
GJMn5E8kLHIzFArVskh6guBjlpk8kMM8Nq+FBvIk/qiSvSFCTG6ngt5P4PkyYdMb
FWqbPkanq/fHUpYKCq/R0HCrVnMPXWaycGnBcw3M2UO0yfyyARhP0IXoAt02qwgl
XvU2xF3O2UU+lRKh5OSXy8Gg/NCdm20XBRTiyndmrpgM2+S9qu8mhZFwP5DMvQQ1
UI4r71TOnt6WKjA0dLHjMbjO1EMjt6hz2aC5cnIJneNYDuLXPqRKaifQmFJ5Qwxb
+Q/lOrewA8zmq2bcQo8D6B0x+ZZzIQl69+74mt91GC0qmYEcTOG/fdOtqP/kfrBk
eo1NwbIYKBCG4UQb6Yns5VeqoqHIdAJObX5eZ/TKdJhn3BbiyBZg+rPq+GxH+MUu
vDhOEdFGdUtl9Ys2xqx3fDtwhyrbvrc9QSfuQk+faQpf2WpOq35P17czuNu/wk3f
I/0bva9qa9M+ER1k48bvc6mdq4Dr+9ZJ/bgWEwIVsH7aa/TVB/JVNY5saAww/qsS
HJkyRNfbeiBk4nKg73jZJheiMJhaNGP3cr3AaPhFGejP3A84lRmhOwsgbxaowHjh
0XDQzTrwWG6dO8vPC5TxM9ux0ZjtvuSzbcYtv/sr86IoDPYO0WUQhd2hLgLchM9r
uhRGvLPYBbwl7SuMLddW+AOTmtK9jkAxJvaSJJV+8QgZsNstbQS4bFUQksTaSOIA
w+QIKKPhY+Yeg9srPbXJuGqTxXuJmTEkGJzEJGyzbH995wi12QPeXFsObWrSgiW6
D0CNk6UJ24K/JTktrxXBluF6godzTC7irmVo1kS3BLNzv9Ur0/R+miTCiaJXCned
1HoYRPKquCMluX9zVYHze32U6OSWs8iD1koMmvXRY5/4WJi2NpmCSw8pclVYlHxB
4xPjfEqlQBr3hYAH9BuIBamRY5uFaC7Y4zm4fcLzsTamn4gnyGuYfmBdXjji1txO
WN5xVOmvj5sCWxtg6kMvA38YIpc6H+a0hgsk+REWTg6SMW1KbtSkRubkt6EF71X6
G9vi32B+1KpmGSbqySMlrrcWQGhn+Y4jZbZOgmh/vNWtbrMkpZAA5d5bbdpZTn30
YlsL7jVB9tIKiWsUKR6j7m904xQ1msU6S7QZz7x1JTOdA1EGSf3ULKCeZ0SxW3yW
r/uQcl/kVht6qfPBM214eH6vjrgbCHMEVKH44aul0xFz/uABUj5GrkqDbHWAqn43
B//Vvv4yx0NYj+0XKG9hHGPNqnSiZ4GbnemT0qbVWwXQRD2IqZJ69SdR102DXk7g
bi6mW/smZTfZBHk1nLvp6JykiGdIe/sM/M1fM/tdWFphNIt3wrxq92n7rbBT5+/d
sKVe4mVFpBENIVYkmmD/dXh9DhwfC2hsV/EefPT2NM6xicQxCAvGmCbVG/2qRToH
+4mE0Shg1DTKyCrqK3gQ3GU5syKlZfentYCE03YixvfMkmB4JgLztdfZU5gvs4zr
o3qpleloAiYkBtBb+ADb2eZbVjanegKcHtfQRIx9HjZ5Ailxeur1IyttGrr8E0PR
JwbqBtprMpnTyweYTssmCan2rPqVKQA2oHM16c/rnaDzNNmyuM9scnKgyx/T/m4G
ky1E8ohAkVuXYJgBz3dME5/9olZLkPF1wK1KeRqZiBCOLlP7WTgozEXw5mKE11tS
dvqgFw0XAEa5SivGl539tnktrR6b9X6j/t5tqthUjDzYBl2CzamSp3kjRNdTcFf2
Ze/dkXpoqGOnsvx5bLLmK15+a02OJzsMhnA/7nBDbazZDBtSZHEY6VJ9tJMdLED2
JqepZlaLw4Srtz1tO6wi4U5vUVqPel7VeG0B9vrMr45d2pFDivRKZDKrW/VZa7b6
V5cdDU6QLk8TTm3p6FHfltjl8mc02Ut1LAv/VcJ0RiHoLTY3aAILqu3kO483JS8O
q+rMY6Ln+0I0KhvrZ8u/YKr0v3bui3fsa/Bj/duA7NyuR4cHaqgHBl/pR6U0Q9ss
YN6NRGSU5AL5IQT6b0w7UoaLCoUZvedpevU2/xYiIEaqPnoQiEqH8hdwevnlkdb2
kCN6HEWCihRyljFdz0kkBH3oQBU8g9zIZyhbPMG5nTXzbJuyQeVXL978VyGxCTRa
1/a2aunjPRoOKd7xcMv8jadztMWmQ8VTosuv08wEN2EX1x2BgJl2AUs8HX3PqFpL
sf/GxkMUUKQePEv1KQpCy5CeLHF06L1hzNzii9oOfuJLmd4UkYVWtc+FZIOJM7W6
kAa3EzCjLx10HeCXUegfWdLmaMyKt9utMMVbjT9MxnLBb1K3i4/DfxCFm4lYj3kU
oTqjeHddbpaTxjdvf+WnoU9n1pYScFba5dRY4gdl8AT89ajV/VeTFrKF7Vk3tVQB
IKIdlewjbY9K1buE/YJv6nA0ISjDQiSl4/tbNvxEfeXTQrflAE1cBC7zEfvVH4VE
OMwKsQb8jWRl/bQwloDU0Kg7s8dYzNDk0Zgc0d3y6PvdkrmugoZJy9D4JqMKcd6A
FoiIczDZ5jDqS7HAoyn6A8q0jcgI/LAciW5Id2izqJSF8B6uZtl8EoEiTBFKIIYO
/wcdYFRH9d3Qg+yuxao7SfVqkWDBYxXG3szTER7zT0AOwnthQzKcHZmVNoVuUXnS
1syYwBL7TYXEdGSub8FQIMRZO67L2pk0/ufljsGLBYCgBcCqIdSFdRbdEk51c3Fx
mKPbux8Q3/XWyxBqZ/fLGm7i9iKYkM/++6c5TyKNDjXFWVfY7O3Koz0UYK7efVnt
RVmmcUCcG/KNdwjsPlf8pE6meCyq8m4Qcd+23xLcfYd2n5B8tMiBvz20i7WAcHm/
5VUA+8/1pjQpET4+ZHYLyYLLfoUhLZoUTJP/WutxALwabVihWUypv8HwaLlPkYdz
GoJ1x40dWSJ5dZ4J4vReHPeO0eK4w7kXlpKbQrEQQSUSq0qhexReVNyjdVLzVfkK
uM8sZDsGyIEb6bSU2LjdPbKKHKlOHKjG19UHT+UXj3LId4BDiSJS5E+Drx58UaY9
XrX8mS/KVIbifLbL9kfG5ix5c0kaaWXA05OwxmULpMUjtG4qVZAGVe1EDw84TqBa
dClVraI9yZXHoMNijmjMuvh5mP8mKu6XE8vYp6XWndAxXJTWvOXBWf/QizKEoJvD
KxcMyGWsr0elzNzp93qtJ5dSwClPSbhpcTMEvphB0fr/WGC18O/Pfj1wNUE2zg40
kT0oT4WA5qrJCcei/JW1nDMDwaVpziDVURH9PRdboSpeAzGkSoiL5M7URnR8Ezdo
CgdxKmuQSlwzDR59+Z9R0XViZ3elWWtGfwFtoXAt3wPiVk7Q6WcaDKbJK2zAdjnx
hL2hbNujnMw2Nj1AbDrH69wY8ZDN7QshvLU6oMOWxEyC+IcVyt+wO8jft/g0p9lY
LKlscinxNmfHcQyN/Z+28d7RnPhYvXOaakpG/UJbtaIRx880Qen2JcPOgc+APWlD
bm/upVkTw+Fpm1E3g462FW3vS4YZou4H+JGhmYeMiVdhjYODafZKN6Mbrbn7nNkP
oeJPa7MeO0JnM2dW1BvuxwSd5zPJ9xWFAozlIzOrB6cIz3ezeNg+Efv4JuomDV5C
DSC6Ql1xUSrihk5GzsekQwhkGWIKwiNvt0pMISaXGy9M4vIJpT1dsfDD6lI0Gt3e
jN8KMElY5ILLxf2dWQ87GtSFnnXMlqM8l5LM2Y0kxH0Co6+dyQOuh4hMM1cQ5d0G
me+QZ+g/0Hwgzve4WH8pfAgN1o8eDSJ/E0oYgLJpAdCtWz4Gd4fOi2wjgtnHZaeA
mQiWc7WzHC/U92oe4zCXi6d1iK7BKxh85p0O0K4PFaEDm6pu0yMvaSvnoAklUEqk
P5+D2XYt+jyoVKNPY+UF20QSKb7p5wLEQfXgjMVmq2j78/5us3eMVV8078AIj5DS
Z1KI/rTyBxSckRVI1eZGY4KeoxARTTRVwQ043QMkKZHtOnbGoj1fh5Wb9j3y6ZM/
483FUMqnAxvhg85xUmWkfV/TrozpT06PkeAbLkQCLAxNHuT9+TtQcd++Lk91QFxl
xFZJZFQyzzX0RkV1hMFpo6i2NKIXErdd+J5iZhals09HerKqRGqPTCK/8ZMw+Zb9
GcwKkdYchs0lpXmNMzbWncox3QyyMFlVJb29L/F0+NWisFJ0UyAQ1xXRWz+xZrcW
+U6s3S14x3Ihp1uKYZ3Vb1fjUWdFK2+4woy3gBr9jA5npdAWkl2sNAGSsmPuu09Z
77GQ8GdfRpDCuN6tkcCj0+7QllhsELl5bHsVuvT5a8u05laO1PlBx69arBUfGMIf
mib/mB0WOOYYmgtqvQBcx+SeOrcWRw2p6sFGysJhbhWMfQC+SN2cwrs0ZI4KuVW2
FeKqKZXuxwnZa4qIg8HB/Ky3yPbyKuqxMl71CBY5KNbI9GeqIfQjPqTFydtuEX9o
pdFPKSGW67XgRw7+HX9ISXw9QIyHaJ7g1c6gXzG1Fik618+s3jgXpoxZSy4m/B1V
GBHH1W8bk0FCUmb4KjbwKhYdwMADmkWdRhIPchrVhZieWzKWvWAo8/XEy8jzP3c2
NRlDO3FW94KjsrQROybHWx7bPPVuJ/Vadvi4xKEoyeVZ5nKK19SRLAlQqHBTZXID
C4+tDDfg8jNQ/WnZf4Ss3Fyfw534F494soN9d5h5U6eE/9KaU9xM/TcfqKNAV1xa
U+PaEk1Bm8W5W4PmqO1lpWWb9AbeiYuL5e8v5dE6jLk8FQH1oXHFXAJSfLGI/4Hm
UtF8jVtfsUrEGrVyiPPHOIhhTDGp2ZFjIKlMFksBkqiIACKaaACXyfpPTCCM/f8K
+6t7ldIjYEDGjDeqVEpssEY2QrzuYbACMsCqnx89l0O2saYsZ9JfH4bg0tnJLp1E
7DnHuqy3vKIuE/JYjYHAUhBL1+uRkb+ldW5VeCHy95E9cSQlTv3yTZhY0kgioYRJ
i9Hp/aQF6Ij03vPM5WGT/KznpFvjrx56173dOhgntnkZuxKMON3k8KOIyFEPz6NK
ZfeB6nH0WiSraEPsMKOuYrDNzlyF6kgtfKmgWbe0DlSy73hLlLwODpoDQoS+YxYO
`protect END_PROTECTED
