`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN+GTBzfN4mJZIkdPovmdv5Ct8ZhmCyHLBCcE4He5T4n
Iw//wiKOTJHgY5GMFVLXxbI1C+PPFTpDD5Mw0Q0zH+r4uj8eYLquPNrHww6TxAXm
VAlZWUkbAjFZOPwePGRC9h26B6RgvvJqtRJmdMCaHep/yr6SE1GkKNiWu9i5F8Mn
QzIRlmL2RDEGEW+UrAtO+QmUJ3KzxfKDEVfqSH7ToP9cITaxmzkeupTvewOprNPm
xD9ZYFoY36ffmVvvrwROo8ez8FR/jhg3uBbAfbrBcTOy+MfPRFa4M/sDWtfkSCMm
DjACTWQHVo6hKMkC5V0yfaR3FHnGg5L5Fn/4nG1debcoFeHZi6PVRgC6VIooRQKk
i7szgDiozRe2fdoEjdPUMbA3ZGIszWJkL2gVS7P4WsUm4foS4Nqqo9neNxpCdFJz
j66o8WhzogwT5FY5Curk1R33xhhyxaRLOo8n9n/3fMl3Mj9968bGjFSqh8U/aP31
jOoptPKCIYBrFy0pteZtaI2YT8LDVsr8QIh6iLYcR28CiussS1UeE1pZLoZ/vPvP
MhKAQZwV0yxTq7rszq3t3WZZdIx6K9sO5lTznc14AVy8gfV9wN90LGTvNrBZM5zD
hQV200RCD2shPHZz975SOUvyzfZByAm/gcSOejOfiOIFkPeCu5Swy4C0FT+ZoGyG
+CH4QVLpMWGrJLcSGJ3lCtXHYg1hMM9Fe4qXrRnYAdA+dvBNUaXpfqaEVOQSs8RW
V/XwFGj9GFwNdcrCWpk3aYyl0w6O7FJagaQ8aU0k9TUGXeIjEyP1w+4TC++JIGWn
HuAHoKz+ayENm9js0NIl9kcZiWMm/lQKlZg+VtN7Cq4=
`protect END_PROTECTED
