`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePRiZmZJvFS+9yCQyfKcqkyhe7rLB+9p07fqbhLgbe9e
O5w9bE8Kop6D7QjQUUfsDXB9qvUvAzlq3EfaNLtB3yao2wn1i7zb2c7YYv69d9DR
6cFFPM83MaHTSlg4eJR6L4RsCKPSlhACbyAsNwtj0W6qs/JpJmNaIg0g7WasWjX8
`protect END_PROTECTED
