`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDLMnkf/KgCsjAmj27D3iwU/Scdqj/hxMv+PFuXb3kt1
bBam766QfMHQmUVWxy+9/pW4jBBKbtNLmNZbGeSWhcHE7BqnKkjpSMFK2iMCZB/+
sdJLuEuH8clWB4fGVxODrUAESc09jnsogvfKH/EI+6FRofb7FTANvJyKOs7VawbT
xqkB2WjimpwGWgQDxl7nNPnE0AwNrO5wiLPnbDplQnvySuWDGLRwg/s0lbDq1Wwr
Flk5vFhYmTbbHUHbTj+bxwSuXhGM4HWMrPMXL09gcharWVReNv6NxrIFhsn4/a22
b1yFhNHStMGolcuyNG2qKiZpYcJflRXlJGOK1TqoVvV1QLcMLEoC3NGWbd9w8yG8
ufhK4k9x/lOn4oRQBcD8+HDxcilJjtykdzrDcl4w7rBvGqO0ihUbQa+kIIsub47u
LgY2uxek9+zbcJ0DSXOG7JUMyI1L872Za/o78Ze/4PX9TDCDR+H9evzZs047qnKW
lGyr/6JJEtaMrhF97z8gcqSuMfw4Bhlg6orRdxyXXQt36p7xnd1RgXAG2fISQ3yb
lilRQbQ/N5F96FWTL+BaFfSnhN8uyu0KWIxHX/O0bZVqcMNnv/iTdg9dxEhdoQ5X
`protect END_PROTECTED
