`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2EBoZu9tBf8wFLCnm6xiM/+CQ1mOdvZEQi7zLD0zwPs2+iE5zym4NaJu9hMRWNsB
I15lYHUpZciM45gP8vUB3hpzrhU0i4O/OcIliO70sFZps27NmfzvvR8lYSjrbq84
dwMe2oK6olTacz1UjHoMwruSVaUYGtI1qnCihegYQT8ETqob4aNZhQqpOiZwpC8u
IRTLT99lL+FGvZASnpkT9nGL28u5Ht+OE3187bUPHEm0+CbsNKrPcoSM/5YUfGHw
pCGbjps6ry9h1L6aASoZfpT9mf3WADI3GhnWY7Vnwk49YAruKgkHyjoFaSYK8nRO
`protect END_PROTECTED
