`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNyl01gMMhKb7u8V0gg5G06Umxh9MQ8N2Ypb4upyR+UrS
NZrhPzUpFpqUflY2IZh0uD3ByimHbbvPjZ++OKDGCI9cICAwT6b1bnxOCf21QL0l
pdqWUZT+d25iStt7yGlhBrPJukX8MuKH6L/uEFA3PMeIuPIFXMVdb9Ic0yuQXlSt
UF2WMzp+QVBAos5lThgpZZHyW/MvWSoZkIW4VSPoZO1HauXS0Upv47qPKOrTxbbc
FFhUN6zqPKO/8wwYnDliglp02rFSNwZZX0qEcWMKNgPieSyHpTJ7Ep0tv/mxAsP/
qh6WyF7ReYbLa8fAl54XEj2HUoT7WDC0VHfchsaWZ19yj56/09FeEtR6OmlNNHWb
60Mvve8HBfSZQtDFV+o5v63+1qD8t5ucpb+WLSEVRugZ7BLCpR/o1KZkWMSI4jp1
91SsSxe1HsBUN33v9DBq3A0Dva86s1K2aEVCdq0xzxB8QLypD083YZbPzEkpvut0
PqohXXBn1bEJFQfjs8sQ7aTx+h3+a/83/cD/vNB26W+PBCK3r6GeR0vwpSMrd1Ge
+ZYH/0djHygMbQttutA+mGVNFfuWneGMvITsax2k+z0C2sowL/2KrvERgAaDemsH
qMh2TeOyNescKe08lzn8tlg2ok1nDbhbFUXpq2C+FuTjcJOTNqOncVpGrdAU7aBr
mU3mtjg6Oc2r0ibuzRHT6CrxsJLAeRqt8Q8gdR8mQnjuBZ3Zfuc89Nq/0ylohYFC
r4bZqkyUzilpZeoi91BrQ2sGi/uMHWawLO0SliFss15bLk87M/5LQ+46WFKlJrAQ
6UVZNnafNPtPWV8WhkYRoiSUv2Zw9eBlYYi/wRtTMKM0q6K73DNkE0E51G6PdFU7
v1TFqBC27R9e6XVyQzHJay0MBFXtuG1M+8MQ/midOi5R+t/M5/nZodxUbIt7WDCY
BlElr76KMSO9lL2N8Scs3waKyh7+lAvW3ctVwvLZ4MGUhgNeVYWftOneRVGU1Dtb
PChytgGhUz66mHQdSumo1zwionXloq6S3sfBnV6s+BA2c0f3ATOlPRlsTrNRhWl2
lynqHvW7avC6wN9H++fIt37YN09cAmMjrKwkJdm0lHBtMLyFb+q0q9TUgSxHsrcl
v0lXPjFNdTF/D/6AtDKYDQ==
`protect END_PROTECTED
