`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4x0zwvlGhzOYmEH9Or8ed4xgl++OzKvlwxB5blBg+972
/UhVM7mJJ0Y0QRbBWSaOYzO756IkyO9RoIQpOrm/kB+IYwE8c3y9CysABjb4nEzP
NnQxBM8UlGQvG8QY1hcKFoYgmtEmblBAcKW+X+Ira1sUf+MiD3hcrPrJBwERaqJl
EwsS06Hn5Srjx5yZcn73iK0ihrRfi83HnyZMNcmt5vs=
`protect END_PROTECTED
