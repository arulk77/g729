`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yYO3EKRQwc2JIpalzy+cE1QKN1ZMKK8y6kDLjPGhCVX
9QTzbd2ptlJ8K0ioMVY6pU9nXuctiACBz3RUq7oPe+JzZq/2NgH5ysfNW5UOiqT9
EsxoEXwe0wM99vhiE2Zl9Pm4HDIkxgZTIKHsAswxGtjgkD02DLrJ7QImjPdh6cIc
04KFrDexM4m9HyVIIQVW+ruXMzlqDuUDfLV73SStJF/uyoRoBovGqBIMJzgEp8Tp
580NfBlsM0RUILm2IzzewJh78pFxp+Tyjo/skErOmAH7kkwXWJlQbwuhEzL8elx2
oQmrM+UiypnSyca4InA2n3xNY5+U/uByc9BT2T79QIqe07pnWR7wqWobw4b6zBGK
MOcVX64nYhkARMDFa7zmvw==
`protect END_PROTECTED
