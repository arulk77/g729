`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHh+afe94gkH4ts2upjTRzyol24TYMriMgO1k037KsN3
F3OzXOhfvenJzrIxODqvGG/26VWxg1K0XdNkv4IwUTgMPR7Eco76x/o5NIP8eYHS
Uvbq5WN7cWWOJjUsiuNyxGJ4valtNLutgVUoX9lRVNBsyl2YqJMIsr8nkv+FaB9W
X2CXoq6XnNsdHn6vfuvVtg==
`protect END_PROTECTED
