`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKPiovRvxBuiGe1PH3ZMQj9WajjCjZMpmJs5C+EbLjui
OqFvZq4fLpAQR1JpAtxxkkt3r7JuCYvXBLroyxKg6AFX3w4KODLzYye9etrnoKDX
yM32lHTE5TXhdMnIdpoqHD7Bnxi63OX93IXyUJTjnNMGzrHGnH0VVMTby3k7ouXb
2ehNxwZo5IXHOXI7zU+cL0lpBkksCkgVzVTBUPvoHUMovXVu97wMeWOo+jesD2sU
3yjTGyYCeZjSlEYSsrG//Ei5pnnhUWThGMNCc+vsTAbusM0UwhecKKOYBttlNIwb
uFS3GtHy/Q7s+d/fkuLv/aFvAtL4+mkEOjDQKtjLpPZpWlVMYkKFCFFT9R35kO23
LQ0B25NibiTyvVD1TtVW0oXYoEhaRfytpNA7dTJ/8qJQ3ra5ZkKvXUr6MAbb4ZXj
eeE/4GHCAp/DuBZxutTuY4zHYfIgu7AAb3JUwvR6mBsA1oc74LdnIz6CIMzoW5W4
1/XJ5jpywnwmROwHeZYlX+YxGgHz81MLtbrx3pFl2IlWUjo2hKCvvIldGMep0e6N
4QY4ATfnFbwnHJvmzLnCKjeSPaP+Ma8BrbFD9YEGP0YKOQJ3CIXvYD+9LuK6Refx
xe3tvVQAnaziIOjTIfic/Lv9aORfrT4c6I/c/LsCnTOc/12TMhH3SSkWMYqIGt5L
KgvnWmsXLGB3VFoNuu9Cs+TRGb7VwoG2rb6x9bqPL4RDPAngvrudGk/CHAtS0ofP
`protect END_PROTECTED
