`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
5ey56rucJoHZ5N0J0OxSFkq6UAybMHLvQ39Wp8bfyRTQD41cyptgTfKL811U3sBJ
u2kttSgAGBaVq4DyqnJVosOpWV4nshsOpJn0Sf9y3/vg1nrn0FK1vslDznbrX0fh
oLfjLKQjZW7egKZUhcDHPs3BP/geoP6GA2IEOqHp5WGgiz9oC4XkTpiAWSuhF0b0
mm2+UySZA98oT52sRUrwCRGA14dcRXZVf19+DSD9LqkVtui6IlX2KSx8JmGm4Fqe
Bi5kdra4rFg3jSWczoPqYFID7qAX3lbQFuOIsJgE0Lrq+k6iwgdcVUIcN0cHH6mg
`protect END_PROTECTED
