`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
MH67kHmvZxiUQFlLMTd3bGXPkpZLdeMdBP4z3wJ/scsYwW6N6pw3zNUAVJ+iiLhw
ZrYC30654VP9bbORMKkZ3orsXZtzfE6YraHk6CmaknyMgH1Wmhmp0cJqsZb6oFzg
ugg0MpfIBumFsjcxgJKz31HOcZHqiORfjEITj00Gs0rtLimhlHeeYll9v3a3ttyu
WbVZtE+ijINTFhFBwSjvtNG8vAK/VCb99iZj3WXQA5k=
`protect END_PROTECTED
