`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
l5IIvWU/koXzsX6Zmfm/h3ISKB6XBwJvh8YjYIlXIc3woj0AfdvaLSgDWKywBiPW
88VoeoJ79GroBVU0jIiSpJ+ssV19t98pRCDuE8LKvW2fd+DhUnzdpASFV/NRDSIY
Rvuqo1EEx9d7YMaD4pPtBjVzyS6RSWyWrUhn8j7xeM5bZT35crejusp15sjWFyKN
fIR5SKLdokg9HZhxOoQqmYc5MP7IiCLeCyndYE+ftbi1RRBZoavBAE/rTx3GqtzC
kWDFsZFT0NR37DzbrJnagRlhE+gg7TokpBN6mFNoP9LAVZqgOyUOp26vSTJunnwm
g+l4Fn3Lr3WnHiPdsSLD0Q==
`protect END_PROTECTED
