`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aQj37yVB6A7hLfr3YnrxxB2tRvw5pGLJO7xnqTWSpO2r
WFlPNFicKwdbNRLCMSMSt3PaeZtacTt/wBhiN2Jmo+lVFT1rPWqzTVs/NprMLyO2
CkDp813S2rM6RcSZXaw4gOcFhAZ7wE+zwhGYEdorGToCgz90HhLRT/vqHMpOYuEB
BV1Vq423T12y0nVqBz8CTFA0wX9oOOAiArHJXHTscClfly4PO2ic4sTwi+gs1EOd
hRCEVVXqYwyJ4DKu25RSLx+xmjJ0WalTnzKG4dhATjl4Y9tnLJX0whp4ic80+IX1
Tld8PB8tp8X2/W2r1IyL8lwwffVX9gzf2iyQtIwcl/y0GqHrYmd3jqujkXUOuq/J
3Q6KBGjOzMH87tnTQlv5hmZcFlQnQrtwbi64q+YCrmDzw214CxJgHQXXNdqerxIK
UxJMBLnooLLOoEiCB4yCUE0lSxQWZ0ja3qJvI2OHx4t/ZUVORDtuqdXDJ1WWmnTb
8c1srp9sKEYReECQTodAQtfAULiyz7VlXn+8xcrfnH3YPWBRPHf7q73+ybhDo280
fseLC180PgbSRCz7a7OE2IasSxp8kqkpIq3r6kr6Il0txfebGVIlFDXUG5XJSZoh
cbUuUkAL/2f4zGy4Noj0PqlMpo9enT7FdmFyIvLzUIca8OpdZjUju/788IsrTTj1
8bLKYjF7sIRj9IGfdHXdjqSD2S/zTJBazkkAXCwcCKlA/pQ1SZleK6i0HBUYYk20
JYk3eSdjWQrPU+NspKkWbSiCq0g2CwcHtG198bVVm5bRh5ePDFUOSwF+aIobCVNf
6fY1MIVrccli1zRmTiY1AwLpBJjFh9/qfKwTdcEkQ7d3NMdMQyDJLRy4mscK4Xd3
IhhsW1yKp8hXDNY4dtY2v9Vbcl5JM9vHRJ1T2a+zlkO0wv9CRbyP8R/9H+4+lXlw
WkHRDTe6N7RkE3P1aROtae+bUb5xTCAJCyXzxwfPGkJkI08j6yM5vVGWlOZVoPVy
KMf2CLdj5wKMTW2bGhUqhlweZlLMv/b1WOGifcuH+hjeHNwPpN2rEUzgryYA5HZ8
ifPr42RBxlvHZwlve3QuLxWj3ynwOfYdOay3i6e29tFQQwPlW+ZIFZkQaw/Itwt8
VmE/06ZyaqOsPSt6EEhKlOkwRmNHgV6eFvUiLJWvTFcmy1jET8H6Eu5WWqs0oLEi
KQonHcjl08DQOOhFSw1buuv9uwg2Je5K7pua/R+phVBkum3RRQ5MjJzLHH6aC8VO
fylUIrFCYipwdaA7JhGyJ3Uk2xjLVb3NffOCctZJ8CFn62sEPrLYsP1MHKPAs9WB
/pOelL42fKMHuWWJSxqmX2I00qEtYVf9tpM09O5Pq4GsswmSkVdX80cewQqAtWNR
nI93e9V/s8KClCfM18gC5yOh7huYEnxn5VIIwYuw5cTaO8SHdzSXxFO4b0dUGgTo
QZiAMQlZvBcWUk9PPV+054ntma6vznJ+qZfGZT3L6YyQKhUC4E5V5NctBUDLRobb
2djsg3VoFyp1E4I9s+OthrobbY2TFmwekNfgQ01Zy1A4/1xaqOnbz056EVOJ6KMd
n+6jOnVR07p60Zd3l89K1hqZa6F98EfCPOAT2ZGl5AXk1peMojdBDCzSXXQ3RTjN
yKMpXRbe3nxcBcN+wAckka8+TXiG5qjAZSYVRcnXspGngS3rE7prvXNTP7zc4ud0
WYX6oZ1FRFvHPkGyOpJe43eAP9lODnf6b6BfgYzxJGb2fycHK+BQGA+ADonsgZ3T
qUrAgP4DSrP0gDMAgGN3t3ok+/43q/IIIgWuxr+x6m6GukxofwCyD+6XtYhs9JHT
6a2L15a2PS+2m9Dn890hrCnoxNTlf3vxXKwdRxraEWKbYT3pw5KxPFVVpVBkoQu4
WVzSsQpz8QG+OBEPTl4rL3UGPxcViP5skn5GDfni2BFGCyxYa2XdmqDjnrq3osyU
qmpHJm65VxQ5HQy3rENg+SLwp4nfnVK07QQoFH8Ojyq7iuzCy08XYJ8EXi6XfxID
mAVXKo2kTaKL7rrSBQBkQEg6St8XaaZYLEjh9Pu01A0i82WopJMdunyproONwntM
7wBln55Qxz0Grc4XKJT7meGm4Bvm05Z/uDfted+sSNd5zanNhSQq+sLo0eDm7HnB
dGvvaVHpIDTYSBvdw3wzrYJqsDFPVz4l4XyR/U54i3lhI4JYErh5PHe/hnT2RsKX
I2AuAKxLjuWEcm/6d+qGVOBONbDETUxpoZipS3ZiKq7O3P2kLtsT9vJPr3xKFfIj
Y8xsEPnMc/CLo3jvKsZSUGiLUMTCIlhKaqVVHGudwaJl5SEOpes6lg8L9Busr0I8
ssk1rqqeRTgMBE/SB3C8Q5hhZRhvO4czhZQKEnU7U2YcUyE4VLppAcbr7DQZpxoH
oCnSqhyija7bevmmXhamyTvIi8Bx29/sg3EMumqukT1KbUa+IhuBQobSKk/GJg+T
fist6OjHP95mpgH6T5aHth+/JMCNXxJebEGWC4OGoJjzHMTjI384C4EpQR/F/z2p
emRuHq0NZJW3EBGSWWXStLT8KqM3hLE9b4TdHExv+t1csr9Dy11QsI32osPhWG42
oc+/0pu7zXHxBu4QFConCTf6M1IkLfuL176QQezxFvwUYWP/qSI0ErLr2wgOZr5l
Ev+VwBZYBRPSoTODzJ3apYAfBUa21DNgKWv1fm6yEpuufzlLFWUcwhALxKR5dTB+
IVtzR1mm3A7ZCuokAqZbmdX+Fzd4A5DbqmwzAXJwEvTO7Uz1ZD3i6DVfPsc2wmQl
z8snFW8qp4uBwiTPlsKHLqJHAlVkzpyK+wdBMDnsEw9zWDG64rEUcVyadxMl/TiY
oyl9xVQIFLBUkizWPzM06TwheUUitNLhI+W+0cqfxwKE7kwslODVCSELLdXWFnW+
KeWbp9zw7/AewLDcYCbzsOjKVEiIGZix8kTsvHlncopcsHW4Vxf8X0im7ORvMI6D
ZiDf/9oWAq/23j2Ec9wASs2l5ni4duGtX/VE5mrQuoNEz3ZPQSJTXkh5rD8V5sb2
U7uwcxQhB7JCAzDao4zrGtMMyc8mpGkXgY1l8UFALGe9WWAIMsTfqD42tfCwhWQs
XfmykgPuxdUK4J7Q9KYrTQXVICdyHXjFb2Hr5v6UdLA875yggvwksFrdiHGPuMQx
NnOLM26BEf3h+5+SFRe9ZU47Kp5OwaUYqF9bXHGWsT+gB6x5YYZDZQsJPW+ffFjD
ttHOkmHsKCif8QXQlb3cxyBv8bCV/eV+/DgkdBink4UKcRlgzxTNBPkDeHCoj5H6
wh5ogBqkv4ATkFIvtieHSoH1Vss9p+42mu6CBbPDbQciIzRIOssrcXV+6mdHkEv0
pw/MagsvyRgQWmq34uUqf73ITgV2UTbGHXSzbEN3WMqk9Vpko0ZSO3dl9O8hWx1P
lvDOnj10+G8bPDmknANSbDLqWn7xcalvOgFl2BpnSSTHPRGtz/qBGjSuYIfuQ/zP
ZmbvE13kgMeDnP7Ym1s5gVCbYDUiNPt51ZZLv6qi8Q/LE+vsSXF6OcJafjh0zmk/
DNAslQFxK746m9fdnPWzd/4VHbCZVHLMeMWPhP9hcYefoQp647vnUW8jmxKMmqKs
t5FwkPUvfukHoqB06JEUlQS74MJUNpAhPkBqKM5POoWcTNCMs2kJxwM5EqlStDWo
i37zsJo+UI8Bkgz5DVy7W0PCb5jcEXM0zfTIWpRiSRlAdj+2o4uLLb21CV4u6AsF
RkC+UqXy2uuO8qM66ocNQWY1BGrRMEsFwFONv1dpwtan4xl7dEUsFcSBrz00qW5x
C/fQ+Vypj++9Ns6Jej37QIBKGHzCiCgET1Phkko27emu/DPyqKnIFfOtIhFC8Bd+
DuxMI6uvGvwqrUXTsIZ8itiVuXmAeJqg1rFuu81xetjB+mrAKgW2NwVy3od3QMVg
xnrfpHPXkBBiBi6EVCF/TKjiu1lyCo7b5NYtxnM94nrG3oya9IFRUI+BW1buerz+
35/vOyxWxebLRwMDiplq70cl9TDTQQ5bhS7/48emapokZrZtmFB8L7Le2/z52SK1
q35TLZd8yLZ3VLHU+/k1dUF+JgnMmGyqyg2nvd9PQEGd+N6DELi+BmjsPRLkNqBb
+uWxaYxHiG9hps2m7U4sq/lzzv6B6887PvZ2ASbpjGmSfYCZEsQGL+5m2Xfq7fqQ
h+5lFpyaLe9Q6yn09j1hl/7uHySgDm3vwJroHVF8lNSvn1kSwILVoRxHzQcrAOso
Mka7Yuc1NMPI/axc4TaqSqmXj8V9EQG/c9/FohrMiJydy6cDItvsE4sY1uGisvWM
J/MnthrIoTDUpIGTEVFkOf3vrUhX47yFiK3Whu0qDIwFhbx8I0D8XRNF0woliC3o
ZC6x7w3Yf5ABqm9K7TN6FeraTLcZFkAX6vTXOuj+7ZVCCQuBX0nbyXxfpbEoRirr
`protect END_PROTECTED
