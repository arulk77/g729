`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveO4KGB41tlwle+x8gB3HMetv0h6tKiqip9Xlbf+kVS8b
SDLm8MtUq4Xv4TvjAJ3BVPTD0oGOcGOwxKsjxtq0+zI9uIl8bBFpbnKO0ed56tjc
1qZ5bgiwFcZEOy/G9u3QEfK2G2B7iPOvdAo+ip3OLx+wISC9yfnllAAkGVUQgix1
MS5YqlUMlMMzRfI7SgGRwPX1ROoiIkqRNIkhpuYcKK1EM5uXe6JHoyCN1avoSRTR
3GWj9GlauB2dIfWlXyu3CC7UVqSWF7Ofb/ks5wiMU8bfSxIB9cAWROO47Zrb6M0e
gEAM5K5ISwv00qM79pk5niv3B7tR1lK3TimxYMd2Aj7d29PxHz77uf8Lc2N7Ulxq
m3cTVY/Z590i51q0Zeustw==
`protect END_PROTECTED
