`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
76sFkWaWtW2g4TUTKwVVqijwifdwriqclHtwXfBDQWt+K0vSCDhIKibHovIci4ec
wnfjZwrTGkHLgFaDxQu9dGaDMxLu6uGCfuframgMh3g/9lEabCJN3pu4sQWSlJhy
HAL3kDSdBiD4Sns8Tr6JPXAqbe/9kWb4LxnLM3B0TDGu/nvDRFhoCEN6yCP/zAMb
cGd1SfU9wxbYmQmjunLOgWChPK+0P3vvN2LuVmVyHRbGVSbi2Mp7JLrGTJhzjTLc
C3+VyEwftHr/3WCYSZXNiAO5a8TbuYTYijOeyevHqmIEgvfr28XYDF7QNlYKBqrr
3DPp2fqo3q0/dCNGQ/oUy1huTlKc/6SwiM6dOg+ZnE7jhZJb0x4g6bnZlTgj3iET
zoV7/XpcXJWkfGs6K8ThD99ZP6qfRCgAbdJVsP1bDak=
`protect END_PROTECTED
