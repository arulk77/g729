`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
9L3gc/xN7FRLHBHsk4laBo6wC184JBTzX1U+bAs3JL4mlkNjThyl0MZEvqOsX0jV
X6+O6O2fW6KKZmib6EjndX7TbsYZeBCG1AGKnDyUh4R8voRI5a2w5g/rjBgHau31
`protect END_PROTECTED
