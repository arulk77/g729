`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN5mATj1YYNd3D4kLAIgrwupFZo62O1ZCnKFeb9S4Q4sM
04Yh6a8UmPkkrYuqu9tGk1O9xKiPTj4ezSLcm2dWco18wt7QGqinFXf00AHdaWnj
74VHpK1civR7K54k+BEtaF4L03nuf5PKjl6EgPAjjP+OyKZf4G9KuZanP5mpNF9O
GecrtdDvUkH5Z0PJjdoPJiRnYYItx4tkKs86CW/kqPCDRWG2kH+lOBe3lIUXoB9r
yfvFKPZpTTkpL1XSybRpSDV5PMtwWo5jIXFJ3YBSXrJoP+vh6ZYz3zBm3K0yHPuu
exA5n5Tp8AuHYfPW6dDgK6VYYHiAwcBKQARi1HR06djoZ3jo1fiNfBFgZc8k2mXj
/TubtTeY2FSLKDOACF2HnEpiseUPgUI5P/aD0qKeuED18v1xGm3kip3oVgArD3yW
jO2Oc7XRmCVcleHK3rpO+Q==
`protect END_PROTECTED
