`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4w1D8AhtTZeoLeevyHhy5kwJxfg4Mm7o6yXWemp9Ydba
tK5CVt38pX1/oD5BsCcliOXttU/0Ciwg5OENtZgrPHmtfAmi0BkEJZ0NKybci8NT
IfbRBnjD5yvWCstTOztq/1WhTIDfE4Sc7pPLdh0s50aYA3y6pxltMMvuetvaVN9q
87ip/CAS907UCcLYviqHbqUNrmNTXrUWfXDxsYO48oX7TOUdFhya7cBVKgUj6ZNl
lDj8nMDGgiavQyomTJ/21D5AH1WEtyjgc6iFIdcAg8Q2+jJrYFRalnXIBWgHZyEV
EDitRFfzz4J/VdXw8mkODQ==
`protect END_PROTECTED
