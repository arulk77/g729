`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
9vUlArzf35uJrVJvy8ozCZdmvMaqcfpdp79fOENQkX0dpi8wip2jHqUASi30oBLY
b5eNoPanXNe9Kly/oBvEZERpAg2iIkTuEtqqHIkGlCh4cueePeJaUpNJOVNbf5ec
qx6KPb2BEr/V/6Gu68qoOkaWGF9vHSX1dXjPyJMWZQgTjcl+XYicAl3lg0sHFF1R
J1i92YClLCZd4MRmMZdHIxt8jqyEh9CrbG9UoBCMVm/rxfA1x82aJBmpMqzYrasy
aygUh+s/XgtJf+dkecIxuHQ9GF0dbyTChN/+2+Z3ewKLWpWDf48YCDU14wBSs37N
dZKeHVQQijuVBS4yDI9IRDnlTmYjaPs+I7xgRqYjHyQgFk3i/KuE2HLAyszhEH8X
pi6sRq+jLVqZqZOp5/TxL5CSKRgNoAad/lnfRdThYOTvBoo27IUIjh+r8N43QM0+
+lhSwms7QuxyimRc2h8oE5fkHHt86Tck31nnI27lvM3A+Vbs4qqci9n0plH+biZU
6iRV5NcjhhzbfDz2XLCWptqyNocPCQdX2+AwPDasxmLrMsn0hDjC196RPLEJLv2N
UqRJoe0aeDlJAVCMqktPM26oZgXweQD6Rr8oB8A1GADUPLv2SNR+QDKrR3vY3/QH
teZT0iAWAPMzg0cgMhcWrgS4nf6Og88a/9lOkmPrgdhBwcPYkynOLTiJ31AgOr7j
vjwst5Cc9ZCB5kN58MBk2E8BuJQ+L0pcAbibaMNBk3YRiBIqcCZApnbE/I4Cpsi4
whB0m3v6xgbUOVmaI0VHiQ==
`protect END_PROTECTED
