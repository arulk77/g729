`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
XeBq1XUE66qJr6xNuSKU70NnsDrziaVlCRTWQXe6mH2sYkg5JiY+boTTqGAktjj1
w7UB3foLb93tRsS9SoUcreqVONd3STd0s/0GpmfBTMWTgiPHjRuAsg466vy7WhgH
v4BN2pIbcCzsf1vGOXpNzv+d9Au2w4dyzmUNQMXb6UsZSRyaCZrL+VUwI7DXMBQq
Fp8oeCrsW5Vg+1IKZ/QCxE5KMw+2aMZVoPgE5CBKEbJJ2awJHu7PAdIx3xEpLWuy
uu5unTKLpvYFa4c/z5wkwZJ2NIstcOHpvmdsaVGIhY7VKlxKTbusn6EGOm2TFb06
2+0S+HZ74xlKewMOAa57589pwG34HZfWWlrgS7fCijLP6lsAg+rZahBi4W4MqW42
Ph66xgElmKYPa5k7jXgsOJ2AWed0C0lHAHw1KOh1SWPyn3ZTkwq2R7Cjhz4Lze1s
myfAE1a5vjm8U3dtDkHn8t8hSjY1vUtpzoqHdNYfDeW7kCe1l9r8YRAcj8QLJUJY
DCZ+U7/p2pW8RR+FSdMhlSl4mHua/86Gvea/ltoeZXQspXe2zzB7T6+Q3ayO4dFV
D8tZaB0BuY4aatFJpsrv/wGMfdJ1TqcSi5G7qgYE6hUsLROXJGmOpmroXaFOuJgN
JjE+QPzyjSE9CzHI9SfBMpdQb0oAFVFJwb769FOet78zIR2TX4dyzR0EMjlgwCzf
ly1ofkoR/WIrcxTCJtWEmdDHUq0eR3GfTw5smy/rqeQwFHSSAtXlUKsWISnHT2TI
2Uf9lVGeipjyC8aL1+WO/aYETMVRL4iVaILZCt447/wBOk/nC1dYgGX+3f2XnpNa
S1xeeyUlCSCXcHUL51XU05hP8vabJM9LWgJmITGKWIi15lZsIknLEN5lccuNvKML
92LOJmbH/dOmDWrMZ3hF0gw5x3lZdz4RwVvhbYtSUb7r+4IjZBo+IBXCbFIiSBm4
uTpPb7u2lGgXSe3WyvpLmUU+ejWdU0wgZNRHEutTRty57WfEvfWokkzWkyhDjhYp
K5Tbg5nLMH7oaUnBFSbF8NmFewtjeFDtyMnLYbqrxXKISaIzBhn/NvJi7cAUBVUb
lYurkLGJIpR9uHtee/FWVtnzxGksii6tAsHEr6qefklJG8xOaeHy9sVxxoZOcfCY
ojdGVjEMTTHSPwri9mSRNFJERH4qN2m6jznClMIO4JnMcXUW0P0EkmSqX96+73tU
22BJ1YeeTyKJzVYYEHuwJzsnpiG+WIfbyyGtrPva/O/jq7ZxGR0Z3KzEc9wKqOw7
vpCZc3HFvVn1pWTemGuCtggpMkqxcfUae3i26Atsl3IunL25TGV1emV365LO9DKy
+/5WJuzz57iXmNOuOIGln5u2g5wFWUbApCC/D7WFCG/NA0e+s62Ch8gU7BTF2X2i
a7S172Vbvvz7aRcCjW+kj6QFI6Z3h12LpzwxhFNwPV6D6gfkbgRmYV5C05oCyo+/
B1mYf6E+0qgWuM4wj7pBH47c7FPFaqbgF91T7/jh0DFQ/F/E/QRxZ4Sx98NPYLEj
YD/zjtlCMvTUvLyyyp5b/v3yrNu/4ulcVS4q0wjXx3bBo1NJ6nF7GOnRhlwuzIZo
m5bQfx+tBqG68lLOo22w4qXPh/R/roYqKDPk9dRux6mHM+qktLXVhd1eiTBYERo8
ljwYTGfWf2pDZiKFc+DM2Qff6IG7FkLzMmhtD92u1DpLtqsLH1pavQGYFEeFQbOD
247CPKS+h9rIawLVWfJla6qA3tn89UW1dKvKw3DkKz+FpqsKkkm3lAEsGdPXE9hZ
+aBiK53eo4/COAQnQNZfZQFHX2le0ga5632nNZFNYPjqzyxY19W+KMOjj3NCb7U8
RuPas1HM69oEHW3UsGJvl6xQQIRJzX/ZshFbMrboeZt1+uHMXdf0w2hvEiBaUOwo
`protect END_PROTECTED
