`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFZeuZ0/R5uUQGUPovuHUDNrcRXblRzkHtsEUTaH4Kun
Ysm8/K8sFxpW5NUTh3vYcbGx4ELXqVh5HPv3aXwqYPzBkinCDfe94wjn+X3yVsYx
IKsvrqXb/xw5ofJ7Zx6nXb4TvEQWS4cbz4CpnpkAjoKf1B/YVk0OQcz81kcsJ9Gi
UZXVsS6gl8OFs2rrjP6YE1NvaZrTsfXMsI5cbstlPoI68ATB+KYTfoRTbV9MxZSO
uQ/x9lvDiFouSzVNAx9iTrHiLM9iFT+Z6an4FDVPKBlHW+hZsyIdG0pvDvRh49O0
fIPV6oiL9YWc9ueR/Usag7978F2UM2IDw5jsONmiKDoiR016gNGEc5fNXABRBGnB
E/ookNhP9SsNJlZpVNDz2wU+eX7748QU1qDb7XlNyLtVg+twAbG7aWwiTEitWMJy
/s5zTBe1LwO4aELC57Vd0EayevFk/Q5IY28If5aKkuasrLuVmrNRH3cyJPmRqs0k
5i5Sy73bGq8fNps1fLUfnjLXXkSy+BC46eER4iNFnVYiA8OdznxFds0r5B7owkfD
`protect END_PROTECTED
