`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
MfGIi5s/tzwgf/7/lI6m9kipn5eJRrjZhyEoQHX3CzNHtPNW8cx1KXA0rGrLajsc
RESAOuNaQjUdTQTrPPbHXYdlBSCtK7QU7bofkYzogq1J5z4YEWuHZmyaliswSwjV
1++HEFSDBNh0FJlTe3la03/BP7cdbb7erWlo4oZeO7awN/b1lWmpnZHmIGgH1SWk
aExkK3RR7iHx2iuPKd+0fSr+Q1/wVn5NBB/MH12jpyrw7vtm4SnIvR6uvPAZWtkF
LWQ/5NF/1yfpJowlfCHM6RLgVs1pBkpGm0VWcTYBSEv+z+t8+0DkzjQJrRPhgZ13
HMv0+kPnDnWsxYdsrLMo/sDZmsexchaegiUeWjVHRQsfl3yxd2bi7aHDFLAFQlax
X8iCwVguyckEwtV23h5ytyreW8EgJVj1ngkV0OLVhpq91Tajtz4zvfABEY8TLG6a
J4VRodYqO1ZyqSBmglXg2e0XshZs6z6juIdsj7XrcsowGsax3jTsV83pkSA9S695
6Hff/FSlwdXletFHi1kuQYhn3m5ZhjQ9fvALU/ye6k1/pALx2eGVeqASfStnaIXm
p19Ku+gQSkW4e6wdKlK8SI/XoNctdDyx4jTEMVVF/wLGgXqoJ/FEfsiY+mK4005d
EWb1fzutCJ1nFfOV+rPdMx9aT5w4tarxNzclw6fpzUOhY5PPwhLPKwkUiiPIrWij
2E3ribcBokdtf/V7U452EYuZG35cxO4Q/4Og6Balwa36uoHg9daBm8gI+mM1/NWk
2SdMf+q0e00pzTY/dbQ5wKgzM3eKTNZnbBMULGpav6n+xTIZ43A4Rt029Dzega08
85TFO7mtHk8FSW6t15hTqx7KEg+3Q31dwtjm95owJN/JqL0m7jPcih2PIJk28VRx
2OWL7G233fcZzNETl2mImsmQbLfPkTZlWBPG0f1+HpntYKYB0A1WbtoPIKLwBu0B
FI7QA0HEB5nBRcDdxEc/lmOBVh2+7rdiMCKFLfXpoMm40aWMXONnUowHvbiQIu8B
sDIXk6X72QsNywoBtMOFIj+KM3o515bh0/k0AbVleaCbkcC8bUqRusrNOoCipIvp
XEZsQBDNT04YktTOz6JLY5FwtwxLugqw71p0YMdqJ7okuBEiy+t0DFJJSATaytrS
RCGzOj0lTqF4wbDtSXieEiTstVvuY5NmIF/e4P/WsKixa+N5z863doZBBjQEA0Z3
V7ukzQGPT45OeLk8dgJnRg71kGa+HlIO7MhTTtyOBj2GOcWVypSsFcjEkAiwmS0V
XB4Kbd5JD1ytOCad7tRKMGSUTbZJRjWKVIGROn0rlDsR+TUA8EOLSHfJS3EYmVH+
zKcJ9xoGHA8mtG0W+ZoR24Q59HR8KEzUh9TkqDeQZL/q1o/OumyftOvuh3XCmc0T
3ToVeUpnsLX9KTVLBrQwZ6q1wRQWf5xz/XT+Ie3YebVeY2Yvol9gOYIyktVSHaXV
X6k2q5ZL7ogeNxSc4MA4oC4iOc19X2hdLvAVbuu/C4bqxpvD0BCTy4AqKAhaiMI3
qgS0982Po+Gak9dsfdny99jAa5Nz9qmu8eAS4k6HcKJu9pkCy8sxOgzMSk2HVGT1
9F8LFE7lWWjhGgPQOxwukxZbpLsorvP6v3aaBjGFCLpIEGmd/evJlZU8Ja76T5Dp
`protect END_PROTECTED
