`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45As7KC5eDBvnwFjzAY7TSEcHvxTV5HHLgPapzw20UZl
4gmMRNxtdnh03G39oUWgzTjcffcjLGuQqv5Zj6DMoFjA9CQ3Nq0xBB8E9XLwBHgx
efDP/izrl6N8TyCAgQmiO8R1We7BfpUWP6Av+TexDW0TNEkjmjurthk07S+WKeC6
oCBaWB+K8kSiTVyTXDPmX1vCJFWBMqSKK/MqA00Uz4UxjLtTVr3ucg0bxwl+atWt
02OPrBd//y/S2UNZe3c87SKdPkFeGeqJsMQjwNKtRLw=
`protect END_PROTECTED
