`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+GkOamKXH0T4LDfk36zNSTzorZ/IMqq5Gc+VTfMwi47
VWBqZwpC/mPdtjdrBri9phq1H6lLLo332ur5/uEOSSRdMDcC6bGTqPIz2pwUybZv
cVezWhR7WEfHFhFHwmf951iDa1wPD95YnHwq6GJ51E8NX8fWBdNVzBKqgs2W0QxX
theuTLv8eAj1qLU4E2X+Zu0wAPaNNlBRbCMyVbqnc6kNTcpiec0AwqkpSGSewOfn
VyrnrW9/8E+pwLM7fjlgwIDVhyrl9Pf3zeVZ/MBX7jI/80TgEV+h9Kp90n/4hkoO
2LR74txQISTZQNWPfM6wF0LUfEYjtVOu5ErSo6SP/Vt0ejjZkzrzPCBxFdp35zyn
ByzHAIiXOvtPm1tetCVgB7pHIHfId/kv0BReBZkIEvryQ+4lCOQ696PtPiH++ALt
9YRXMhSPfOXdPCQualOOiQStu7BC/TQeYzHCmyd+07nQT2xBGTkcLuwC3DolLsYQ
flJ3IU+8RtKEws5fhBh3veuMP793HFqK6zGhkWiIQILwOJ7qfk2qxmbBFscwasmI
YYnsKVfuVUrE5iK9tORvjn3NA2gCybuR4jHrHO4Kx76acCL1DjxvlLgHG1/Bvnx7
mtIqaRnAYaKk7FEuDuosEl0lDB826sdojgLV3amPV50oeuhgvSae5hjq3cSSn3rQ
q0Woqy/Oa1C30DHT9rztXVAh4f4E7CaDgYI3JzinN04=
`protect END_PROTECTED
