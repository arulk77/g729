`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
KvdtJf49CjbB76HOW2Ajbf0i58VZD6dBUfLVH2rD2ylUUGqDNtP+jvpk0k+cgatU
KhLW6FzI/fmAPgcsnAcUqMwC23npgYLMaeruSD/F6hONZA21FXGMMbeukwnk9hCs
BQXWxit97rcbgEWrATfeFNmV3iSQZgyrKNT3Cz+DSXBXGoXIwON34BxoTBKz4781
dnLQjczTvN93u7hxM3DVdhoLB1lMKmvaFmE2YkrRBiyWiOt36wTIBfjCfC4YahG/
`protect END_PROTECTED
