`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJoJJQMVdH8PmLh7PeFJk6tJGnitSXYXWc8LpC+MpdLH
omLs7op1CRhzKZJubrSAGTQVcLbkOFXW8/tQlFc4uu9h8ErPMaAXexVd54eqfdna
uqQFZQdLytLIeeGwjAG2B71nNkqiejUs+ZkJU0qxAOHi3ftrb1PFTmzfltrKM3w8
XboF1nIPseeW4sVQM5fONA==
`protect END_PROTECTED
