`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEzQDr2iB89s59YL7/UbVWBfrWgpz54I2vfY5tSPziVa
CRbSFd6FlKNH4yexfhbyt+aXDgFy625qXGkYo42CrGIcTJYDShYII20IwiY1g28T
nV88zaiwWlrObqBnTjthutFxj0hZGmDfcMCz+JlPxuF5Xdq4lJTDzy51PdsW6EBp
IGxS9OwksYw9P5i0r5HiaX6q9j4sXAyYe7W9xsOJ8G8o7ykUot8Cku6jlcrzobRg
zkZfxn0ir85FxRQ3aqC5ZPEaCtVITffc2f0I9R0VncH6JOihpAYm+sIKHZGu9A0t
0N5BpLmP1nXzKZD9niniHd20r7dudliedn7gUmnRszC6E1gkXRgJHSLC7U3lneZ1
0tsHqPYbqOJkW55v9/aiMD4nS6x2bj5SWeIDLffVKECDMFlKBq3xbb9mrNfyww65
rOP+xqxeWsiezsAkA4yZxx65/UXvjdAAJoh3bRIhTvsBByHzC9fl8RTwnGDth7CC
78OJ3D8wRoLHv8gpD6urfw==
`protect END_PROTECTED
