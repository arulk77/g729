`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI+u4DczMVcO+cpR+Se+fkJcbkoEuDKgWFEnC5SMyZ2I
AhaC2ujMB0zKcyDruu3Xz7+I4JTR8ijiBP+FFBbm8jclkGXD8Rw3+5yqVRDke3Jv
lankN2YQCQG/9spstnGvVQQzXlzmbaV8qam+ZEA7aaBqft8G6qfIU96nD8vBvdyN
SXlPgyeGbccQiHiZ8QVnMMOd8Ndcx57XD8Zw6SK9vlIES1EPq06xCLlhB3lL1hg5
`protect END_PROTECTED
