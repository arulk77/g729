`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCdmlVPdNp5AktH+69NurN07o5iEPlrnAwtqEtMfLfhb
gCZ8tgZ8nfMizTuEFXZiNYSTFl5HPEnVsc+WvaU2uYh4cCLgKezzY/7DbowubDWh
Ch956gGS62hFh69jFJqdd9XeuxTv+4YcUVDjhk5ORZBCrkGAyqP6XqxTxObKUIZS
Tk90omryWpXZTwSiJpMTaqYrtnJBDKlJRY2eizpQpIs/hMOlzkKEEvvXZegu2PU6
PXIHUu8pSABKayKlEl0bQjJ/iQqEx9dxeMbcXREUUvRocoyxxyey9h19X9TPsUNC
JBumFftayPmbxFmwdhu3L0UbfBYXltp7z6EEVwAmh7PJsfga8CN6pIUFUe+vSR2C
TACeM49enwvx/ujeJu2M2JaWzdLGGPVn+gFgOg+Oc3OuoiB4TlOc/6XT7qsuC5L7
kAgC6HI2iNt6UIKHNbPeMYsd8XrMqj0U4wK/2VCSqEmy515bFrfb+QolZPVhAbbt
`protect END_PROTECTED
