`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKsYVZ2LhVHzpOLIMXnW+MX7LEibIw9TsB1BF48AdEpe
qamw1y+/MMu1LgnT9nVtUrGgCQRUFAzAr56/5msHQKEg8gPU4eViCmAhnq4Xfxj+
CRXfWnGO7C5Glj39LUJgdY2Bmh0hvyGcS2Eh6rlAu8jBRo7uSP82RojfIqaxahcB
9uO3UDOxVDWsWeq4Pri6YeNCX2dhE5wdTqh5ZZm5LSp3T+4+IPknBEW+DeHqXc0A
`protect END_PROTECTED
