`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM1zVUjTaG728tK+GdKEGW4A1SW40yk/tG31YvnF+Mvu
hnx5tnepfuBLWk9gGO1u+L4uxfNM2ipRPNTq63dCrhnD2SE5GensgNVoTV/8t0JC
d5pMgnLN+pux897ql/4cvXiFDG1rZWonFnQmwEQbpgSDaJn7dqmu1wu7xvvwYi41
Z5HI0wnNaXWykPygGiwuSz29iVSGtMeYxtiq9qMXqUWCf68dU7kdybcAzzRb9zar
Tu/9eelFL5Nacfbdul0U3o5VmBk5tlhMWre+ZhL2mdIWYOiz+j8HFxUH5/3sMpbl
HTSykRyHy6+IASqbyrq315hS8GiAzZTqWJ87scmBxCt7s4hmU7C1ogxkkedJp21T
bZZkicZtT/6YsSoNIZr3b5gAbaEHgCPFoL8OEGHArBEopY64lQmcDIpPK8wta/tg
9x4HsqKGOR4Lk1pMLktDNFThGW491I8Nqa5u79kaVPMc94jRjMrkw/VuahBAPA3d
OUzmE2tYAp/CY0zcA2wzzv6zszWKRJ4z48hZjB+PgCkicnt3KF6ShEV7OVkYZuRv
vmpA92U7gZarWaINkxDCFQLK04GUr3DKvD/2iQqSGX4kiiLVSTezvCI6tEYxmYlZ
s2JZPn83k04B50ZMxj8J3HA8ya8zyu6yofv8pQCnUJnOYJpZrR8y9g5gftrK01Xv
3piyUCLMOqFtiqqyqdRLt+1ltNODVqOumC8PhGiyzvbh6TTJ9xqVjRIdlXOLkIXX
lpyzmPyDJr4Xe7cZAvhcJqmkBZsYSJY0qlj6GiHU+3Fnoa/EomMida8kgRjXiIDO
jxt5k+/sMbJbuXgydsSUjIhf6rChGsu5fdRyCfoNOBE=
`protect END_PROTECTED
