`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveD99L7bqcy9Bz9/4THExAcB3KIm+gJ26JMgij+N1zVKk
ys2Xa+qfdlvQtsmu4UPx6WdCkcVCgfC6npMFzU0BV9xPdjLTtP8DJuTttCN2fi1+
hoQVLqYGTEN61QngUuzZ88kyTVhNAhBV7HY0kD7YjghSna5+pZvv3HEo8lcCuK4V
ypHne1fJRa7gv+lgYhnvXnIkbUyn3DD+7ZaLSCljyv+eM+ZgU4NztZ/M+/p64lkR
tVJAq6vGgowsQicOuuQtsi3hdbXKRtDayMV7WVtpVIBjybB4BS/m5KYy76BxOQ+O
1ZXYUkQ7jIljNIB8Ul0NQN6XuFLPjvobhTCtW4J0GQX3TboJKg5W2W08Fi+0AIdW
UhfazKYiXzmRJZI6W2FDJVOCOpWomQfDPB5C4NqdeCSkq9W/Cai4UPkFNX4BPQvV
dWgEWofPGdlrrMAq0+XBzJJYV35fdSDklDsietaDHTvgiWgQD72iijiLc8pWtpbf
`protect END_PROTECTED
