library verilog;
use verilog.vl_types.all;
entity IOBUFDS_DIFF_OUT is
    generic(
        DIFF_TERM       : string  := "FALSE";
        IBUF_LOW_PWR    : string  := "TRUE";
        IOSTANDARD      : string  := "DEFAULT"
    );
    port(
        O               : out    vl_logic;
        OB              : out    vl_logic;
        IO              : inout  vl_logic;
        IOB             : inout  vl_logic;
        I               : in     vl_logic;
        TM              : in     vl_logic;
        TS              : in     vl_logic
    );
end IOBUFDS_DIFF_OUT;
