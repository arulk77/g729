`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C7MA7dDoxapmm4AuQKeqZg7/CNYTKknt06qiiXtmR1m/
n956uFygj4cLbTSHlqFgDEtN6TI6Xu7DgIqdCpLnw01oS+WTnerAmkyYIskRfa1a
MMcBu3yucd4z2wvz76U/0aQBNlc59MeodOcC2vV6OwgJJBjDfCLnaSllMKFvzNMc
MerMQLDsOFqcCh1F+OKqEBf68dc5UPeCABXQEJngFqpKbelThSaA0zk1Qqo86Zv0
5XsyBCDEVErn/iGcHrBWrZUmkvD/Y7IjKDw0fo+3Eq7HCxFmKJ8HqzBbhE+879gZ
Wgv0GKr+X63CQU3JVZ5/1JGSI8Ielp1mILho+HPn7IAXHbwqDKI6fT/gPtT66wLs
gQNqalpL+CZt2aAlEhWHbuMQ7iPWHRMvi4dox6g3dXjuLecJGVn+sx51XakxkWU+
+ujV2+9Tw3Cu7bfH9yGHlgZwsSuAA5wjGU3Tg1MNc5ozsV6Bpq5upuBzQ0jbR0PL
kuYiMDxjs7m03qVM7wr3l9MBKUzwgy7ipxrjasMypp0abqwJ0/lk111xEF4T/uDC
2PmzW415eCZ6VYhyiKp/k1aNRhlfv5N0Y6/tJzYZvOcMioGmt+2Hjno0aJX4SQ58
dB06jIpk/rdpxSxNdQO7yNnoPt6QmQgtyzlO7PerNT/XSTtaUZbb/cgce+sBGBuB
8YvzBQzpzX6dho+LtkzHTwThECU5tSVZV7WtTQvnhoW2xTjGUObNluV/kNTl6EIf
/D7CyqAkTCvfybewbFiZ4P4YD5o+woWuSZM9+kf+xh8OBWqs+ueColMVq7yzTcty
hCvXT1KXAmT0bN4Ggkq7V88wbjEaHDh3wZ6XF87h9MnIJBej5fTjbRzbsZHGbZkO
LSxymkA6uH7tLqDqPe0pyBqKqq9B+qeId0I+oWgGTFed8fyLl92M8RJX5znmxNqb
ieLm90XASbVKUzi3d/yTmsDuTLHF/CzFTw/YvJWXWG1dorxbQMHdhvdkVeD2ZhWp
S3hPKHygDm10IeZmCwRAsDn2AnNQgd8dNBj8i2Caxo7TSsSCHq8kNJvx3S3qUSzw
e8X8GkmBw4aVXgKgLi8GWnOHuu/9nhCcXnkIhMY6CwQJwDfkYk4ZqLK5cMDXxJn7
4XDKYEwMwXXTdv2YaLjBgPN/2zAILFwsZ9IvsiwWZTfXs/yWmyflEfSgE1p6fwSV
iNK0sifyFeg++h+qhtcOsHKpgcJvjssc7v3ePOX2VnMtr8xn3HW0JX5eg2vS3egD
IgrzcyN42kuhhDptbuGLjNYqU+50UyQRmLtlJOnzzHDb34dKIu6wtvuM64bonQ3l
kASdob9DNQSN3/C1vwXM5xCAjj3Mx4gI/OJqIbE4JyNA2hlZiSoh5JUGHFYf9Di1
4/prfltef34dr6mcO1ohcW0Cld+frXSjDLPEcEKOWUph79OD+SxVKIc1XlSbvFob
wCAooA3f/orOzTzZxN6iW/Qg6BAuhRkmyv9k3VAqYisgie8gNogrDD4aH99LTFG9
AUWdk9ImOfcBxAfSf6i2bHaapSht+vIChCKMHW/DPdCiPoe7INosZYOpnYyz0ERD
AyOTvnvNj4yy7Ajw7M3Gjq2ZdJztQGELgCkls8k2SUyoTLfkcKzuY2gyAplC1Bpw
I/r3BX3JYwAIQp7PH9P2qS6U8t9mA6fNRUChf2tc3FImP4k4pgsdFR+sNbmr6i7I
b4qUhGdF62hTM+RapdMP1bgrQqc+7B7DQWo+7WSepbI7x/eI8wOZppXVby1Y2KKm
sHDTL0RyDpMHsO7G6Z0OXDRReNyOSzatKnesZHD3JqzqXSWiXNcD+uwkO0dWd2Kw
ovGCe3KgrI8PAu7lanZ05AmMeZv10eHgrbXomsWgautvlRGRtkGjwfqhQLrUhs+Q
eJN32z6Lu0LT+uasqNpvj/UdFn2Jbczdc7VPvnlM/AbnAjCZnrAt7fHFPI+8XtR8
oSugA3Q/JTsHJAJDHSANhVP9FHqz+91eIQISopPzyURkOxvrNABuAQV5u1GiTXWw
p+W9TV/qeE05iQN1LGoWOJ84CEAOdHF+Oa0SyzUh5jtzRO3B7JqVGiMBa2+Jjbpj
Nn9Cho4cjcHljwkP3ignUPJ79nBL/4cR7VQB9PS/w20f/icEzkAAEKjF/1sidirx
zbMpA2F9dBAWhDXd3+6SrDNewOxBgKeF9j2/dchL/y1kMQbxtY92MeTayGbX3zd2
5afw31ordm6uNXMChVNRnMSI0PzxTmYBTQCPsuw0Q/4oKPRBLPTvUYA6wVmRgE3H
xApptmqSke9bdGatQZ0f24k8lg4Jf/vq/J1e7nBL0w9sWGKKRxqgg0tuS3SGjvch
LzRNpMjghK03LrNzzwt6AkS1zAlX7HYrHpnrEETVAfYkkOcdaMbSj2B58o3Opg/T
iY4KC+TfxGpcak6eu55bbmqFMWxi7iX3KFQGjbaj8luT5NLrPuVe/WpVZVeORW1F
bumniXe533OH2CvaFoVUoqgWIzwDnGZSu7gmJYbMxol9PwoKm11yUBC0i2w0yNQ0
8W7vSTeOWAQmij2HoPcJBzqZMhYk9gAEmxXw8YYF1FkMNbUlqq3tEB1cRu8NghSL
NF8I9+xfQhgMbhC9ySfw6mq0mngPJucyWin064Gz8tIlCxSGWrM69lwhxGXj73jF
X9jJAyR3TC1i+lJpxZfRW1ireATqLBrBXEv4+DII19lHs6aLQdaXpUpXafXKzd0d
Us+TJxJgJJdzNsCKR8X8YDZP9By7LtntszNhHxf2Yezj9o1euQ3wGcWoXnf4fOam
30sx79O6avyCFPA+V+np5NDgnXT+xG5UmidLEtZTopgxrdVOxNQ+8wAlQ2VR0MhU
yv5B1+ImxLXBGJhJy245wxbdcC097ptUREYeF8cOxca/JSY6hNbP6gcSrVuCXFc7
QecKDMK1BoR0BZE8AdCwx0UX0idVgmS1wSr54cKHEzpFh+nQH3Mmst82BB/TxmN2
aflCTShfl22dE305LR/+CRWtJ8iCuClaGeBhPpd9cPG8y8UFYImrqX420UQVawec
5NJTt11nJLPVYYJ84ng2Ba3N0bLD0p8esE6R71sLPdSu2DdFANARwURRX9TehxlR
fA7cSyh3rx50OyXgJH4wK949I0a00+MzvqdRCDZbV1Rj/1XGHaA2edoa2a10FRlc
XV3I2G5onBNo7V73l/Et5xSt/L9wnxIU3vjtkxKpaXdcIbhraXDfCBgE6BPamL5h
VPl4XlLaw7uiTy39NvN+gGl6rdvasWzD71PJXdYjulokPO0Ux25WYYz4p1YME9im
LmZNyTDO76C5wOQx1C7ZZnt0k1FIobzlavETHe/EBk8Gii4Ris3dZTHcWOeVzyMn
UXaETf1PTZbXPV3pOtAP7c25/lHb0WleU3+z20oimEXKYFimpvNnfl7uFfhsQjJQ
LhehoLeegUPz4HIKaU9NofuOhH2HsdHKRIXBN1nn2hKFaty0wEzSomsBlW/aMevD
DfD+I38lO7ICoPwU+Pm+TJrEwfiuCBKQpf3Fr/uSpcF8xnTwrYOXcuS4CnLayGU1
gKpB9E36hrnyMaosih1TXnDSSfsjzDrpZeMKxS8SvUsOcDTWR3Rh/C2qcYUGw05Y
XrchfB1hyBcLCJiGCTh6ZZTwt6sesPpyoTiIwHG1LDwiLLBCBM+7TvAteF1+40OY
VXj+wnVV3xgrJIbClxoP9fmmDfQjJNMskSyTEZDWV+Rkhwox6UyG4D4P/W+tDfwy
mPsqezRTTNv+9GwnFZdR0hEpGAg9t+q5bfmgYLHLMpQPwMpY1UUhauYiijw3Ju+9
R0HMz1wKQlKY16RIr9u74LORIkbcmfGf4OQsxkME6vWm9gWEy+ImU73qln5KS3sI
unPVZpLv+bRv6LlaQPbYQlvvuLcFQ7hX2mG1JroYX7PVM/+DN0tTagSry2Y1QH7p
HBp4BA3TdTwZDVwxEJSRQuGJFS1xLEgz6aGlB3sr4MDnk0k1HdD+s65sK6brrsWJ
G6SDc2k91xZ1ebx/tUtDeHB+f35iLCiyLTj6OJPEuCNNVAa30J5IZrCoadkshNiY
aX14A78ZDIwkjDrc57PPuOGoRoW5/JlgRSC6bdWaFXlWJsS5QP/m/yoEqOFy9KT9
uYzhjZK9+0QXKIrYLFkvbQ6isPVNQD3vKnfY+pzKagYdSzQEUF13XI6l4Fwpsia+
PuncOVzpknrBirGkC7tcxUkAUtcNtq2AKynwJrALetAV63Lpjfc+nEN1aI0td6lD
SXx7x2kmYiseWfDcBMKszDVHHkXSSocz/PVL5LRCCnrKrHx29lP6Ja8nKEXYNcKx
hJ+QHyMVL4YEBl4b2Jp0Nh6UpX4dMQH7ApGRQ0mW/5mO8fChEGXPDu/TqQ3MnC6X
Em2jR/lAIWiB5A7RQloRM/yv3IzGn79DgajLdNK+bXn5DRIcp1b8RUpSO4ps9fO3
EVcS4Hx2/FzugpVC3q2W5f9uQVioLPL6/rjFH4U2pvVHUl/ehXpyBF5LPbDa/nfZ
Ehov3pwzoNklBdo5R5nKKarUx139v5pIeL5VhCIy51sUz9+y4wEnn9nJQpkWRA+p
VcbzDGyV8vQLVtQtnpJYD5tBh8r0loXGXg9Fe231yH1lG4q+j7Pb3fgy2K+dp5aL
WmHvPpI/TpXDhrglDO1eemLLyf7GHH60kYaCheip0TU=
`protect END_PROTECTED
