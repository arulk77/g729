`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40W6zpYbVnjnBugTejDIIaF+gAjBqSDckV2YaxOiSLOc
LoR/0vI5zEKy/pvCKWTg60TWEZo6FgQpKDfn8hKiJKcwAEF5x/C3w1+GNbj2K0hr
zUKFO0w16LHICEXoQZiW7PrJrCI+Y0y2lA450TZSMykYPxOZ16fvgcKxnGWwcnxr
wObyVzQMgKh5BFAC9ipVEkymY4M2HcnoBYYfDURucLhhMbw8sTpTCwFsyeXmXa5J
jG3pTllagkiPxWuGQXyKXUclEQCOzKviFkcXGe7lEgsbU/YaA2ki7kbbzkR8OZOu
31kFZT9UWYUGEbKX6cE8IQ==
`protect END_PROTECTED
