`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49ZnIdn3BohHgAXWmmID/qEgNagUjPm4c0vISF0JLUu0
L8cBqKJXwmdSYbc0z1zZfPpDQaPooF6uJzLYmnCYOUVqaP4zBQ4thnCaEYRqYDz5
Fj8Isan+zKw556k6R8UfyjL747qhCWaeiq1B0yY49o0nFQYOWJr8f/Jp08QUU05W
3+D/vklyFqGKGOLW6stKJ2obs2JeE2hVqEneQSFRzfxyu+OSxKMAMNfz5uwtYrGO
AhvP2tQTWKqfUJyO7RnzcJud7RzSqugitRHeYbzYKdSiWzah//jkCUPBgPZ3j/Hd
N85IJksLWQ1Jd0rNYfEAUg==
`protect END_PROTECTED
