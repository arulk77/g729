`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJCY68kNy4fSVefZveMSUWU+637wVnpYR3SNjmOS26IE
D51Zzw8zGvyxhLLnDd8/sjtcYZSr2DFO5J5c7SBkt8GjaKknFNkondflpvAKmZMh
I/PyqRBfGRoOLclvE7AhU8Yq+3cb4UyK3QCw3lpPlTWQcMpa2Fh9MX/wP+kJSi0E
/iFw9AOzjbGcjIc0foK1BMY28iZ5xqmzmq7hvlK2iS4HU1OsrczKnAwqRCIxdekY
tuE0VDsoBnGpjDgjSYHqFHBYq9AF7zluhYYcoVxTT/HgeQmKwuL9Un77YudozFey
XqSlRLk0TbPeWxDlPz5xS3iw2LEzEKe3sv8bu4cXYVIpLldOstafNyBjBID5zhAk
ay1K0ehHQPm1oe/aDa2rUw==
`protect END_PROTECTED
