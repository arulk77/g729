`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C0mjvQMvlCbKCXkG+KulNcpRXnJj4SdhVlyqPBYXxVZh
7Fhn2Gyvh6XStnJMaKLvSQFgRKXhm0in7UAMnEXgpLEZOyZAoPKkIF/TQYac5bu8
GuTo/FMPROZSS+HupbIFLXp98RyZvJ+Ly81AbtKe7cWnPswH/vbr+dYkQFmRRmeC
o2SjvE9aFlelamIfkrgOFFFvVQUFwMSogKhrGe8kaAg4TC7EEw3CtTNxJ8tnx7Oa
bgZHe8P3dtbhljms8bf32hZt0vO1peVTtdLBMa2+v7E/W27wazlWfxJV69AV9uYh
QflRfSe67291c5EwPbf0GU1lHnq3Jyes5rgWxFNI793b5VNNZ/XEdJ/JyASjHpEv
mVdmbrUph4m2fD3wsTwzgi3dFjAhEegAmAu3UCSYHg0u2tt254e9PhwJtxRMqulE
QmHAsk90zpI68YplWxRdr3sVVhbgvg3LDNlYTH09ef3YKrj1G4QzFDV9vKggl1Uo
hRrKpeNy7/Zsi3KjkQltKcSRj0JldZoueZm1xGIvnd8=
`protect END_PROTECTED
