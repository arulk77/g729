`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pl6EgbJo2emAcLzkfX5I8rPZR2ysNW2Y4kRsOBMZEG2+FWhwCqTirEZRjlRUFjkF
Tm9cDMZCwu3oFuQMSUVCnFeF5WZKqz6PdvNdjZIC+KhCfyiuHmNyBRR2SMmpk/YH
E5+L9FkLNd7Xa3m9u327LXcU3/9xeXbFa6j2KwRHsTL7whDtSitD2QyDsFHgMXTD
GUWcRuglTToibl/V3CAi2g7hYwvlIPNGsjnHdUqarJw=
`protect END_PROTECTED
