`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJiXF3XcFBggy8gZHds17s4RtnBshYnZFUQbmvyf8e2w
rgpvwUICSVH3Cd/EWYZmvMfP9CuLOdcmUj3G+VdY0gIHKrdYI5QFN2rFqOpB1uTx
VWEDEms7HMk+NXnUKeYZGv/Rhzh7JFgvcXsKCbMmGRMaCbrB2juczPHedbO6iYvv
scUTwy1JtxQWWBObHp6EJPhkduxiaxW7nqBC/uSv12MG0jG1cr0piFhzQSvS0dQh
YQiXnzLW8ahcHVj8ZQzo6cDllekVnph430lGo03Fxkm3JI2GWjksSVuz0b2qb1KX
cuMP6b8uuDHYiW8Y+AbwW85F6QHGjByE6vQm6nmXIjgH3GxOm0anSpzPw51jjZ7r
ZTKA6xtJDz/3QdOAkf0901QBefok1yCmWKH/UTciKR0+DSWd7fGzFEHC/C+18c/m
9pbLD4te25ixEqxKUKiYDNIAZLyEcYqyBwA87m7uIwg6vAmlbsNOb3scvER8WIkr
`protect END_PROTECTED
