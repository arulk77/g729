`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGPUMhBjMBNUFeBrRxCfMw60YvebjQx1kqpna2z6w/VK
NPYJpCaVMAcBLlXs1N7Q6kcAhGM94H6+fsIlZoCdZ1e2SCrIUSCedy3jfkpraKzi
0B7JW/9ag2YZJdBbYNUfjlbxmgXMJHXLvb/PzpHLs3S91lIgbTGWgmSmyA2EAcUw
K6uPVWTp+gQvEkAeTypXVcBfGmoNWxELA08jZpxKlAVWNe/OuulnGirIXEuA9SHO
WWCKX/2isxL6IHyqympjhcQht4esjkeKuaB1pUMkIcTOObFVtGOxbVI0ovzaEOeM
aKcnQV+HrtUHMKxnoR+qR6MLFGkHkkvsR19YbAxf985uoGRh06IZzfU2HsR5yrZh
LrxXfKvq4fhkRGoWVKjVubG/PpVSaw+U7UcFLKp3bsmzxTICNyd0YujR6db/jPci
gas1K5Emm7v8SEv2uz6ZIn2clEiOlgg0ht6geDIMu7eIOM/wmNOlEePO9koMaEzd
fJmvjoJY2QX73cF8Zkf0ZiXwTbSwKElHQBhQCI7PKb/q0O9/Fi/TJakQb3gxyXQ8
`protect END_PROTECTED
