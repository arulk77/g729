`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
t5E6rwKtTSfAaZuC9gJnCvaWqVI4Ctmu0oImNXW2zLByV7mED34diodvb/FRqiUB
n4Qch1fJi7cuMtMYzZf67j2WKXcnd9vRByEfnXKcwU2UYhAKOBNfVA3CATqiqZmH
+PQv45kUvUWpudLWF0aqq6QsdwM5sFx/GoIGyqHsFS34tMA1VLcTAYpUATM30Kx3
`protect END_PROTECTED
