`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkS5D6ZJUH+KDZVzPaWXRwEmPqZxQWCQnQVmp1Q54Zsil
miASQwf87r5Wi2ePgpUrMZYzHCsbHhUk2wbHT/xv0gy5C/M+zpA9wLOIzJ+7yx+e
Ecme2pkc7yvJpxOMpmIlZyWWR34aVoL9b7vzwspKY5Qx90QnwsIvQmbn68Iejwzj
eeUBwX+IBIHLr9SAWT5AiWYhy2UTQ4KTyaIzO5TusZCDSxnDhb3RuN46GKjpgEIf
Pw8W0cLlY+d/ynOhF3ONpbYXZGqO2AwH2RBzPysawZJtzlU2OseI5ohi0jdRNnRq
lvV9KQ1hGEJd1wgkcyWYtoO30jor2q8LG9pKLMiO0YLfPBL48qQVUeIeJrSM3eYs
1ebxgalmDNzdvbJNo6AvrMqFVjMET6gTmbyeCAZgh1X5guMr/l2NvHbRxTGjRGUQ
TOF6wKu9hLZBSmXLOtX4+NmNs4YGGFE/Io/zV+OtBucCmyi8ZvQtTmaHVWqxHUoD
ZdtWpXxWa0rTgeQe8Nooah7r0hOyha1cXIrvRShKi+DnpDkyApT7GFKUXE6wE977
WOau11w2XBnjDQ3iYY1USvDNo4aTuvAaOuO69bZHua3yz8dl18HqfGnbUVRKY0iu
wC/UnQjx5RV7afXEenCqhYhBD5/PVDdPZaIn4Iai2nedKryBOtvYQz4xJWQZA0jd
XqxKcFiX68VEDxm2AkqjklvI2E1IES3TBix9Bi0XkHYkn4SnlA5zQvMKe+9ytmTZ
3MLk2F71MHOs4UZMhMMbtC9Ywf+OpZ+vEberS/sveoq9XpcDS3FmICfgYsSjC82Y
lTEQZOn0hY62X1GTzyCbOQ==
`protect END_PROTECTED
