`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu484sl2mBoECn+dJYZXAJlC5asihGOootqJD4y+Mvwpbj
/9f89rdeXP3EMk3sDlDK17IZzB+l9yYXbC5kSAjO0th+csXtDwzojA0jrSjOVVdC
A2kq5fuq7qKhTtXoeKIj5IgnWEXt1GJeEqrMPzAvyztZ72oeiPje6jyUqCkRCnoS
opTacKFM5TOFpsGHj36JEL2MEA3NisSkIKgzZSkhbeHaSy4hCX9D49gGl1jgz7Ka
jEbGtZXdI2qcGG72L3+KWpHzYvqf8OaRIjh2nPbxmPc=
`protect END_PROTECTED
