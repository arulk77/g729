`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveABsVDU+oIjuwsYlSv/C14Hf1Il6iSY7WiKU9m0eBls7
ZM+LX1A5EMVCyU7sQxIO5gKqXJsYrVZQdOI4A/ofgj193/ZxRsi2gT0odnHEMkY/
jnzre94hJl/DQzJ9/L97EHen7Yz2vhZdivmhr4kJ5/fNiyAbm3V1RqaRbFwGdjXo
bcIBvOvgVn7OpGxkJw6dlKNLMn7K99m+Xg2ZE60ixafOssdpXHly2Ef0ctllq/TP
ZFCsZx3goh5tf2dps+mlYD4p9hGdGsyzc87U6LVR1dmmJnB+ULZBvqu7qBR1qvxD
swvDa6q5ayStYbfMzoEcZs9dtinSrdT5pPUtraGQpF7s9FWw1zAMnWCSGOZJKyOL
OeTA+K97vX3rsl0PRtvOEA==
`protect END_PROTECTED
