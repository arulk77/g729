`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SfySEWt5zJqm6S62s1qbl5ZZve6J4/p5It5cupxTIYfr
rWGl0IHjAC1GjoJIOMFK8HrDYW/4gEn7/wifW9PJW7EYGR0EwmaOXIkWxYx/xOx5
6ennRhbxadOAV1zmUMg9Lse3dlXKjJVfzun8RZQlTnFxhXF0s6SzUqV7wUFoy8zj
ts9dpLcQ0YIi7deUQ2bci3AYW4bUXvv7b6xpxkuVqfyLCkCbdMdeQtdPkvrvXCTc
WLCF0ptT8nLybFljqZnr1E5FS7xS/mL2mPxLn2vYobY1YHoUtbyy82SyPM+qy0fs
XkxXWbtamln44pIfgGcwX03JbGN7h5xc6WFQ4UeQv13vowcdb2SOiwJfMmohJA3y
kjVDPNmQs6Z3mQ+AA+VN8GMKOGdPWGFoS/UsJQTtI4jEvFMLDHZ50G4q/BzRoPVE
lNcv4/IecSp26CgY5vb3FL6NB6ODeUTZ0px18vDRW4QHbYs3hb4u5q7dOya7YL0T
raieko33mYRYC60/quacR5yiSg0sYibtikz1Vc9DGnlfiLD2SPdr4dDcqJbQYmyi
QBzFYlPZWtKu83RJsNgcrAntDDeMgJ0DkHOiiN387ISocJwqfsmVlR3bPYbCv8za
AqNuMMlhZ5aiDjXcDUP+GvKq5Ixwu4qHUYDrC90cYv6VfhSPfBW41eVN8agtyT0/
k1LKpO0Q/hCEr6TU8B4HaTbTpGaTy6frwTiisWg8UvY493Av07s16NvMC2AlGjg3
YesxFClF0sGNs+SQnxqE6AbUZYmPM7W1uySwUWsDrpUQHnSA5VzN8ZVNvg9p3UBr
l8TF7NSIpRQiOmYPD7iaXCRoXEPMb5nA6YkH91HkjZ7zjacIchVO3VkepGSBqmQq
zzqhQbxRKOj2Ot34ItWWV0BZJL4FAM0bSHDiuStyVzMGVd6265tjXB1svzllW7qz
tD1ENOkl32V86NNS0uwxB8Qn7Vb9k0xRLkhD3LxhGmBM199CcLyLLz4/2RxwrXWe
CHSgkmOHZniO6qZqRg87EH6Y/FiLcjIgNKe0w4OC+C1NrX28mhBFBENK87HUxL1/
Wscvk1d3ITMqlCBJAYKvkIXeBsKgTcnOsakXJPySn2ZauvODM/xg6HZE8X/khDGu
LFRsS53Txoz1h3M+0pIErx8NkVC1qYXAyEzPNpsj/dxDGD069etfD7nkP6ZyNzQN
U3PMvc/oItuKoMtUhg0yWGmnO4fvm5f9AiOYCus9gnYkhcE7TP4M73cXqaF93pPq
TuNfBab6VnY137/eXz/wtrvuy0I9nWGd6ts2oZY839o5es36KnberBL/y7nL3SvR
c0/yNJ3wZLp4knAQx8J7DkaaptI6ga97nuEqEwpVU0IGzjkNwgesRA8FrrUTuLvK
i5t9m/aPujELH2xFWyaL500PXEP4jUR4cf5Ck5lJmtNn5uJHFsN+gGD2qhTJsFjk
7ZSZL//T8R2sULe9GbzJvOcAW+vPuw6XKNLRS3EAI4eyq1beGOkv1A+PGuIWHvmV
II9mcuTeNlJie0uQmbddYcS2iQlXixaIISxGzakCEnuJx4QxKpz9xFyBlIZvlbTb
/Ff4vIxQ20AC1xcbftGgQR0I0Ao+FNiwH71iMUbKxR7dCW1vXkd/rkulBK2tqjf4
3Z7jRLUv0zzenNVCHcfqM3ptootXa67cWQP+5UP22Tcrn+cMkVyyURBMcxqZPDlf
fBXs0G5VrYRxYpSCHb6YPE354+bYAoK+2mUrjKYWB4C7EUI5oVU/kuHGZYuuaS1n
ys0n9kNOdQqZJmEMyJ1UMdPqgSJcUk7gZB/zHcIzAgGJOGASldho0Z8fQbvgIgzR
MQqvIwFQ/hY3gGXl8T4B620nlYvdqJR/zao/KPYI4lXfB1u1Yw9PF+NBaW4fckqc
opSkJ+4UVknoZnxuLZBYEWtPVRZDuL4LOzyeJLIg+4ZBgHTwHvZQV0epMsK2Nr4C
FDKgdm7yvdjCNCMAsZvy7GSNduVNRFtHsvjvmR6c1C1lfk2E1sZk88PJV5shxguz
tTNvYxN4KUzonLOP7geXg/dt7n59KWC9hMuA9OXdQTwkFl4ZxxWTeIwanNfQA/4X
qaIzFf19wEOsXvzXF0tQuUSCI9VqRqbkiMnT/zjm0QUJKag7YPd6RPt0K/t1IqG2
qw3yRidKyc8Xj40e1ACPE+oBspsXCLNEkO925nn2C2wFxSOrF3SP4xXlAgqUqJZX
Qr90iOZ17zRclpzkNLCYttxiny9e1Qivxk+BEvH+7o4DpUXnnJcf8mkP1sRIXjOj
HTFRK3BEr8v/xT/DRlcf9jo7VUDy+ffPSbcw5VoTIIibdpR6Iqeyx/+OscamRprO
ZXd/xbZPzoRwtvpv6+GiNSGOe8dG2NVuB26tEDRWxv1BcyiQstrCw7V7ZBmcz90j
lDh/byTyib7z7jF6w1WYSmzIcWgg5AyB5hUT+BIDS1CUZfmGbmot6TxJzRmN3uv1
6uW6/EgRpaSpQ8bWtDV2LculFAEOsjLu6ZcAfXPIKAe/MSZTUrfHuhNW6ewPSpic
`protect END_PROTECTED
