`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SYoIZrUE+kRIyLgIqYnX3IstCQq3+8BwP1RpYVxamxcT
RUUDMxSWNHDdG9uXLG7D2KwQpqCNweRF19NNywmSgjsikbj25jWglFXx3DV1P98z
glcJBLr31byz8n7t3k1xgGld4o50zuP2VAay0iBKJg98va5hQHqGBZN4nIPZTUk+
luOlfIkvWv0lOFQWf2X2BZ8DrIAbgMygWoSeNhyVsotblyyv6QlLVWXvF8NXgotn
l3ZPajYd5nkYGk3H+pS7UWcZslk88xElPZgmDDPYp6vQv5jxfpZ4anbSOgnJUWUU
Nfbhp5zzhBjlCWzOy+qTwTwnL5481ctLOOtI0KyCNMVOLlZqZA3vzZOtFCYhR/3M
KGKbN7tg+ETMS4E67n4HxrwaszJX+pHg/2fGV6OnD3XNxKlV/joPvlZFzN+uQ7Qz
YTCWkzb09m85OoxT3y2PRNnx1OVnCAPmzAPInut3vhEWtv50hdB69QxcpQj8G03o
4eR3mdYJ9cPLfbRS4/jfgPEJ7tuH63Zr48HzzedpJtA84wCgIhU6LEHIEx4RE32k
QR81EENAGBcyp3ggFSvA2UZtUHIR9cd29q7W8fGLKQTom/QWe3LP/zxAZwiz9TRz
47AkbU3mHGc9qbOCQNtHQW8UNRPfmtX9cld95befdV9u/Ql2Xs14OhyWtkUv+IMN
WeQnZS79vJzV8PB99GDbnPBxrfq69QluSjU//4OdqqgBTusccP+UJKZHR0ZVmDmh
ZvSUVgcroCRcBZB/v8rfHN09XwNoVoMaIyA6jIAMUy0z+8itVCnQ6iRBr6NtUky0
33pIgebIkAZLjG756eIAHERvl9FG6Q/2mLFUklFKLKBMzURiTX6QUN4Ig+YPwwRz
JxsjsaS4BdHcYiL4ot5YmntZLkoJdKaPp0wYjfmVpbUSeKI/5TlSrnOcdvo+8S0n
R1U1rJM8T7C1yI9BBbHgfmFrbTVtDyWfBaFOD9fVmR9pffN36Fh8fwLNwdw5hB4B
vI0SNAGKDxWJCNmtl8YrLwLup384uNpxuzj4ho6uH7DF2KfxVEel+GsT9J65E4dL
3RiNDToxnH1gcmp/qrGvYhv4/qZpPavOKzbYq6JqZTS4NULeMmbf1kKF+wL9NPvd
yhMHTyKAIGZ1LGw/aOaBszXUMWmhTO93RZbdAnErnKhlvUwki6UlBzIXAqVjN0Ge
6ThNsM084WiNyefXVVHlvBG5ke4KCS3glZDVtkJWOPUIyi2AYGIk4aTW3vgC2zu0
dQZZTSE2NH1T9d+PD01tGQ==
`protect END_PROTECTED
