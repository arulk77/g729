`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI9aV2Qux5T+vEzJyngN/mbWGlpTD58H83p3wBh0rOLA
+6K015oyE7ZWOeGykLrOB4CCRVqfL0iEbQ8JNRQYCcfQo2UNYJ3XMTaK11jBDRhp
xagQ1OvXCZSkOwlr7IOw1NTPiE+n6Em7qmm4G95qevW8N8fWE5oas6EV0BL38DSh
iWOe/xiHEaM5kQ5G4CcfrQ==
`protect END_PROTECTED
