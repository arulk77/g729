`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
88N772/WG+n8blsJvcIQlRHR4JcQTaHGWqZHRTfFb1GbFaIEw80uGj0rOjlmtcDd
jmn3Ixug+Wr2QzYaM6siyJ0Nag44cKFNYqWbbwz2K4E7kswy3vh+HfvldyZoy6eo
eYcolM6DJgV6QfduH3ktiAQrAbYlHpY3UXU7/7wKHGc80wdiB7iRfnSAkYykbYTh
`protect END_PROTECTED
