`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveETdLI+XH3TWFW0Ud9my/jqpEGvtnaHpbdCUxu8KQ9No
vsy0sO0h9CyB2gVcz3CCvxVp/kX9hNsdb9aHWWj8hPUjQm2YlzdljuUAf1g5Kcw0
Vobws8eiS4LTyAOr1sVUIyg5NmiFw6sPfn3YtB3CY6vlE1vCaY7x6USAuAf8zBKB
QMqHmU4DnePr8Gz2GEGEwknqTAg1IkUUEWuvF2SW/xPa9+R5s1ZBFMN3knH+AxWc
jNz5wBu3dwOCpq/kP84lQQ==
`protect END_PROTECTED
