`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePKlgDMDM4uoFdWDO0iwpeyzmvbZewmDy50z8V4DQbOR
peWqogkabB9jB0UQhY/V0o39RUM7JiE5ChIzTy2io7P297eIYsjWjVAfWxxGLuhy
1ldM1AaoVQT7OkovdGqzD35uNxBlK6ffbEIZbNyyt7jbRshffWzM/yQeiru7J4eR
a2RmioJ4EQHJVz8kBeXNkVPwG55Z3UeDHSDjL6QZ88qbdwSMBOWJbi3Ay6EBmdg2
Z2WUqj5kSEX5de8uhXAmk69KbQJCiSU25z5REz/ZL8oFXkfhvby71OXSaa9V/f9f
3Lgw80+elx4N1rZT/K8+ZonYfl3EvByT/ntCM22+MAAlA233xfiJ1u7+PBcvxtQD
6AL5EDGnOK3dfW3oSVPuqyMVGoxe4en5OMBWOuqpJN9DLuF/v1vPHOFCSpitquw9
KJr0lMOQOVtx8KRkLWCT+mhD6nbQ/5zugykLOQVN3FwCkGkFfyOIhGZHQM3IxEqQ
gVIkQuhSuh1pVdxpSHwy3XUOVC9pV0lD6WSbMY8ggY0Ejuy5W/M7NCdwoSftJUNF
vijem+CwSEAeniOznBUjqRZ/pzY9SJKrvZgTXSOUSy4NJIF2M+F8lu6razVX7C4u
`protect END_PROTECTED
