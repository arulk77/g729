`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bxCmrOkaFBAI/MlotJrDer1VaSP8PAmz26W/gIZ587LTXj2PZ5YHhj3ErNFhOKAh
sE7W1iJDAz+7lk4Y0p9PxPJv2/fK+jrSq11ZniNCOhj/KVFbWP70zQfA83PtY57E
bYrJzlIN24rpRqbUcVfod2HVLp+e17F/YzM5OD8J18Bb6Sbm476EVfRi5+LaTcGO
2SqqDF/SvLYU9w7o3TyR2878LhdDB58daOgbOzbzmyaBOZSiklhkfYEXejgrdP5f
9zOC3MaYmR2xtva7yDgAmJ4s3bfyPciYcdSr+yfGD0Wq54+OTrR33KuilVZvE9kG
fbRvzQG5pxnEVa75ow0+d7gCYEG3/DJOYnS8/emd9VS5Cm/0GXGxVPbWKoYS3hou
gZg6Pk8Q7u+X5J8bhpeHmTBZXSO9jZkEmc89LdCyNqbWf/ikmoZMKV9y8CjPHmCk
i1FH1BYsI3vq2TBtxk/0CVmg4l1xPCqNhhAHoeOKiPYrY2uyDSeEQ4VIW5FIgdCq
c3P0LEzB9q59S/rZv5/EaGKlmy0g7EYORjDLhtpcU+P7Sq/oq7t0uQltHcQPR5qJ
f3si0WHxfW8luBiTBlOAl1QZNYJieYjzzAPcpKQuaUXTzj7+8jPAV/BH3dFzOcwe
NEF0sn11ytOxHimZjDDT8CFU0alnMYN74461saYlV9BWNmwcn7ZW394oCQRb1EE0
7l23E+uEGQCzPi52jQxM3Q==
`protect END_PROTECTED
