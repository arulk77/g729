`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48w9M+8Myt/BrpeRw4osAPVGBW6uDrdqgN3DdbLSAQbs
X5+XmEAvLWs8w+0XF6/+7scn2a/o03fLDlkV6XgEHvxfJvGkBDRRxqywekgbkh8J
6G1NmHmBNEgzUOyCU6NhqPSp94uHQi3vejdQwK7O148BpbQz3NuHraJ1jpJeY8hM
yFJhPmjG2Uea6Um9w9EdBQGNJ3iukHI7HsQIAbg+e60=
`protect END_PROTECTED
