`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
nmt4o3UN/z5Krw/9Af68LqVKrswHfSDdZbkvv8Pg3upL2I3oeBtpGpFyiIpyRkSz
1m0CpMqLaKKDeKPkagD+pSgDXPZQnkL/KpXCJH6Hi1+3TQiV9F8z00H1Ht+N0nLq
uqaz2uQOhBW16jzBGP29YY3+X9vuwbSmOhDF3pq7XGgu+lMbUC/LLpEtlCnK5VU4
1wgXhFUsRFCTNhaB5YtMnpKw9C7ncBcTnZjPwRwFCFE=
`protect END_PROTECTED
