`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL82IMNsptQI/a0dcIWLt0Uwbv2n8OMQ/JIrW2vqHXtV07
Yukxk6qqwm/jGI8dbyqKKyHDHmoOa+EMwDo281+9pu9YTwUUx1zEt6XPKji7GkUR
kUyvFSUFDVdp1BZswfQ5F8gXnZL/DpRtv5IV0SH67/wNCEwHq7LXYlTaEl9mAlh3
7H4SenG8grzf/WfZxSDEAXtVkiXjUIMyaMxqW9gQNlmhjb55pfPFtrjTVPRX+tY9
lXaoF4Oko31SB37zHRG9sl14fcQKcK9ZWSgdEwJ61JXaR7Xioz1Id5yXQ7FcOxNE
8mjJvIVuotnpG89IQKk8OuvyiIxZB29/e5gGuU/DYKq5TjwsEmEhgrk0FZxPPs2B
rIOUvxZOH02XURHbhmy5QPIG0wgCDAAlsBId2EM3ay298pXHGnoEuIbgoxJKNLHD
`protect END_PROTECTED
