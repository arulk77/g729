`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMOxN6lSN3SLWMngSZ26RVoOKJjwGU7x2oc6g5YLhnVa
ZclWTusau4iDqkA7McPS8ufE8dsAtbawWPySstPLZxTYAxdGrdUfmMOp5VzUTxu2
jR3i5dBLxd8/mwWJXvr/EuShh9zKn4neVHbF8jnBMOkhJhU9/gg7wwHS4tWlc0nO
ALMsK9dw8+FWOfFH3BPbx7SOSDs8pc3HbOg1UBX9eDr0ULddFzfgq2vvzFkVcUu+
9sRhcUr41JaXTxCge97WoyfpFQd77T2bM8ix7StuIRG3neYnLMh2bC/6CTygsSPi
LRyK3hhk782Q4qrOfDHM8DIels7k5Lks7tC2IC+JiKA72W14JzlUn7zG/R8GWcmh
F9F/WPStEX5Fz7kUukL0bqF84N1IMxQyNusEW1SqxKh3StetIPdEZZJ95ot9tXn/
U8+m1xEs5DY3ScBfs4JC/93+NdB7fTN6UwIwQH/Q5wPlpTpmUctqFztvPLSsWknT
c2E4gT8LTPBmH/d4TPsTfzM4JIPOrLv3OZXf6B6TYFE9Tb7BlDD8MZ7xZa1f5aX9
xRdwnU29k2P6vxF8teJD4II5MJOK83maV4qAPXa12nbcqGBjhXbePxgxHgQg7+D4
VnjTIE3551zh4/yTLtaHPQC5bEN0/CfhJyyrwRKluv7+a5XEug3l//BKw9j7H8Nm
`protect END_PROTECTED
