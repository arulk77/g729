`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCCqiED+5RQYCqU6VZolYYtkT9qA0/pEdGjfiVbTi7eE
sq8pWr8NL7K2yN4KPtrO4r0u28ACjRYes0DGBkspH4Ul0eqHsC/HLl19tuDhYtVI
U8r1NH3bbdQ66Q+D0L+HNS5Wyv4yJiBz16F4qUo4EzBruf98UzcCFRwV0hfzuiKK
/3RbqTHovt8aBg0ieCd7u9JBhxD1/AAcPp45JqvIIAkuLxRlE+oOSIzLTwjhI4Fd
`protect END_PROTECTED
