`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
A9leOttBlKAk9cVgktXpuNWNDTte4NtZbSI1zmgWhb+n7iOm56Eeq7vmMmj5GJya
I5qPkRS5CP6jsSMsJhy/UPDyE8VK2/V8WkZs19+HTxiw84P+Y9X4p2aA2HWMYABB
Uy8mKF61C/MSgke3YWN0KH3/7Y4NWJEp/U/5kmI5qaRtFa+H3aUqYmp146jJ6P9z
/VoE91Jdp0IdevCby6yrVD/BEA+PvsftbuQGfRjrMxU=
`protect END_PROTECTED
