`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+zvweXVudMsq6yjJ8D1uWS0F5MkGy/U4XCZRVA4FBiE
Ig2twNAqOeEdM0GYWDNqEzOZj51MRawglJ/XYV3UFvg1AblSDeKtmeJJBqwq4boH
MXMX4DAoR2JL8bMJVttF9MNMPtFinFFsHLh4TMlEEwk1Qc/R9zRlINeCTRE94YMC
LVmhOtcA8xdcIwjALgbSmzWvH/Edbz2iau+O0IK3D3c=
`protect END_PROTECTED
