`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePWjz6Q8dZAapGIT+0eWOV2xbirjZe4pK9QaIqN34dwL
taQSFmLeI0rA7h7NZbByUYkKsQwcmn8QElAScZzAE0S5nNWKSzO74Uotik32fJXW
kNUXpEdoLKHTLxc+i4A7dV9bMbv2XnSPmoLETnFI7ERwrDznsBPy/D6z4VslUs+H
0XIeZrGXiggDtogCjslXfObnH3rFeekDkQ8r1esPFEcQKM1gv/uBnaUg4ITU0yUg
NdRW2O3zGqkODfLDZ57aAjlq75pF7Wp/eFkkKvj2YLYriDGai3hPoZ3Dwzve4De0
dbvzHIAQZfe4nC38dF0+wCEwM2L8TguGrdibd4TzCVp9uQsKurxi6bkvsx+Mix3S
3Z6RwHr2aI5JIFnUB4mZINhCsFlr+Scvs83uT1aLdkfSdqq8q69u2smg3JzCbRzM
4+hAKhrkc927si6R1NKSzc0WZny5rGGv1yOMDfwHG7/o1OUOzl34kAJThNsgTo6T
vE+n8wcStWtPXT9qh/j8rZa2/q72hM9QHioPdH0d/fZ0SFHy3kjfaajdf4TerJFW
`protect END_PROTECTED
