`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
l+0tOY6z0IXLOiaMf9aV2ChMwuAkOWgIHmlozBfPYh41H6P4h5d17eNj/9ufGE9Z
rhFvxmbI3V9I9i/540nmXv9lm0+sKDnFdVNsjtciWX1b1ayxj+2ISZbmcep7RAOG
Lj/z3zJKr6C5yq6l3EK4HbCnOakgXE9GQRJ2tdw651He4IqmFvsd6RXX2xoxdLEM
zT4swPHzBWa+DTPl1oan+TFwUlfhypWyNGuhmyiyESjV7G3sZ8GXpWN3HsZrJpTT
`protect END_PROTECTED
