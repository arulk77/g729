`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFDbjlgSKbE7zz/3L673c9P0EE+E/82kYnZu1zODlFz5
4Dq5cI3MZIAksfQV8Han+LI/WkFkfwGTShkyJ/YjNUM9jIW48RVi9/HQ4+pqAduJ
tRIFOXBLN5cjNMoHaTGphH8u/mSsmvgWxf3gdKAGdlC4Px7PHTCe+u7mAL06F0XW
LFHliQesa6huFe6J4qfuBO1gUrztQdrTB7noBpITW7ZdNMoiSX4wFgKJ6AMfdxwO
`protect END_PROTECTED
