`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK7ht3lVGDzdxQld5VvVWiqzRZY0E682YLw1z1KIPWgh
7euOY2k2ZIUxSU3QvXT5OtTJtZxyHFKl0R5QSr+tEle0UymSmzXLTFvkFHL8wD6g
tdwZyHHoWo4QT2lg92ODLRnKkCSISHQAr2IoQpb+zlxgUEI2mH/6VBB3JiyWd7kk
KJyAheLprM1qS3AslaGlOeQ/YgZgf+9W3779JRRlOf5ndX/Fu8xoU6+X004OPZ2N
8JdIArQiX6Uteasl4NeR3n0BPultHCGRfw+WB8Kf9EW3h3NhHW78Piz+xF52RcBb
SfHVAegvms/B5MqZEoZeLV5oY16rHM76SnHBuewIvtwIN2wYnWEUhG1bwcme5mam
dKRvwvJxLLgHg7SJRy5lzixcS0DG0e4DHjsD9s2S1yfhWv9ZFQpHpKJ9wJQQtBOf
ORxKY4Gc6167Np0b7rDUbPc+/Ig4FRamxK1/AKr7dJUHAekIqkT9p2oE9WbKYqCC
4LTuCL6zB1mgihLVFIRqdSqAQueI2R/uPWI40yzfAjcG0xXlFeNPeeOm/i5JdAcv
0zHYG0zOgzuCLX5/yLKzT7vonEbYoQuNc1adT2iyRqM5H2FXBsDodB63MPURbrNo
zEwjlVxatmRZcFAKPPZLafvUhcqNqkpbfwbcmwUpVJP17Py6hUmv4RJJg772Hw8w
`protect END_PROTECTED
