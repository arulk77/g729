`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNtIn7QjuRke9KeRdfAXSK/eVIRTKkBWFnJFf+TIRqB5
6D6L3EBiERWsNjCP/2/H4GUHaK1ZRtlDVzy1Ihp10hlR5TZqF0Dbe/+lqhhPEdV4
/0bz7pPwB9GePYAslVIopFFGo0la6Z3FWZYZjVPjF3KZT8uOe5OXX6CkXphwJr1O
ahlzA7ZiSGnC2lvjeoJ67w==
`protect END_PROTECTED
