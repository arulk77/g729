`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
NRypGAWsdkI9SGQWdP8vLwtKjxMU59yxs4vdmFlDsUKugzDWTRR5d9xb8VJq7kg6
DyxlX2GhsNpO7W1q6mC4VHyeNbw4hP+5JdoGBljAQld+HfBxJC7zzr1w/V2nfXzj
sqX26Wu+76GdxGtD3vkisMfvL3YYsV3Lo/cWPJNdDefjK0oAlAEbH7vol1nt/UkC
4R8V/hkhfk7NfDw0GLwAzHsFXMfSttkKGtpHOSsjFbn4Z8EiQSx9s4Nz6KTrS2r6
FdjkqK7+mlTo8hU7KctYojO6cOJWbO/A1J4l9mjP90QRVvpb4SZLyDvISC90RvfF
H6MAe4bQM7fBmcDqM97PYpW5oXbFOeAB4Y4nEGish3r29tQ8aerL+Re5Y+dkuXVf
aVIEuq9H21MDlb6KJ+NRKX0b9h6IX6+mUbHwrW02r0iq7rNZgCJO44N1AcqPa7+g
fpeUtLDn1K2uSgW0nvo6/eG1rAM9neCqto66PHcFVCOeaWOLM0Ds1/1Wa4tbvsaj
oTrwIMGDhCUSvVGjbyjoKuCZL25C4pSc+eLYob9X9dXCJuP1S+PTQ6qeyyTtmh9z
Y1twvLd+IKvaEQBQMnBS8w==
`protect END_PROTECTED
