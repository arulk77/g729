`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu472ozQhQu45rGgTE2O0BuhB5TvB3bsKGRqAKTvNnFXzS
bITBV2eg5iC2Lo2Aur6k3kQRhlm3yer6hKKYGDk0gfP0ezOcTNXcGfJpcGwZN2lb
++wHPhkcQtk19vOxItnjyLQTUF7IlywSYrk337jQjOfRLePTcmRz2X59epQ5bkQF
/DJ2V+YpymTUhWdk1NMgrLbLsMDZQTzKbm7p8SqjoUW3SayBX4BKSxVg871kReos
cYP1gSKOqqr1CDLo5A+yDsywXNa/y6x0acOayFbfU9o=
`protect END_PROTECTED
