`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40hauMxgkitYPD3ZaJsni6XW6jPIHscR4x/KE2d2tv6o
RxnUSLVNMXnDU4g5708FGrGysH9H/uGKvsL4c/DwilI0bmIFKmn7AhMvJYPI5KlX
0LPqQ4nU9KsLLEAGqogurBa9Mm+1bx7tGeQovdP/KWqg5fMm1DuaoyV93wBwAb8d
DzlmJjh53R7zh7n9D0OJgwGBKbs5S9VwmL6gpoP9BQoPV6fNIVxgszHKgbi+tthG
FWcYFkf8cZX0KgFdtnDbIYSl9LeAJcrVvaALe+pXX/d7+wRCn/PFTfck+oUQLJy7
TEqV7eYsO4hUdW/ZsIyxLHJgEYAhTQa36c2vI9vGCpM/Jj/6KOhiOsPpkPCbb73r
A0ihTwrd+qm5gs0a+ZWa30jmu6pn9AcXTmtnTGKNSLxRsKPNdj2PPG56dDs+jcU0
1oPImA6XyG/4T81+DP6kcw==
`protect END_PROTECTED
