`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFEw5CH9csWM2pFjjlYLqIkM8O8FTvHOJJaZOYkdG1qQ
sCyrDxHpWlgEci1iVmN2wBgkgHGYM6q2g4LTDWTA1UzlgMDuojnNC+RwT418aKTo
OHowf9v9hgqXZknn0o6HXeM4Y9X6kaFpWC6/uAeXu+qhTHz54/Iat3otNtR7hCY8
t78NSWw3FFBRfo/9KnMIqdhAmqlU5YH8t2twC8oj4to52rf9Z1fYTkuVVe2ULkiO
ehzmHXn9JjIIbHqFw49MQtOes53vcJ5BZNkdLasQhc4+3BlAxonBQwUzL25oSVuc
GYGLTFu+2Ynu7+oiXKdAgzOXVzyoJxoJwfF2XcLWpsMtnfKjDvagDOTFDt1iKe6k
+XwLLc+Im73Y2I8ZHX+DwDnPgQTuhNf6OHKjQDR8wBwDDMjOjnkKWzE+QKHsFYps
8BFv09PZOAToHkeghAvwPswfUpyXMOqJ77NnySMBOAUN41Wk2+PV5r0X0KsDTy1O
nJF4hkPm+pNp3+bc+gDnlYNdEHg7n492YxX+qOma7zxxeropPKDkCnVvVCuJ45aB
083rODSxjhAy9MEREj9Q4UmHmbYf+rvI2QDAPdDChvpaew2UcPi0WRTRsuKb6Jni
`protect END_PROTECTED
