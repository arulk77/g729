`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBwbPS/9fJWE7pMBg5DH9huPE7qAl7pLVr2rekXfu7dn
HQ1KTxNbz8wUig+lNWuq007xqIY+NK8o82L6po+LEAWrn344PvaSN+AbsVTgzK9f
nZ8hT5djc25dIVcaQY1qvFJfkjIWV4nIFe0+llCKKMOY6gClPy3XyeoVKJTkvjp/
VYn9dL/kFvxvYDGCI0xi/a1BZPbaUE7XJ/xsgSsB855XED/0+yFJNQ2UOJE4Z/B9
IcGMzspw+DKWdm06iZXYoL9dVeyUUBrVDQhyCEY0TK0Pgg6j89r5HbG85Z2kOFMm
+LEtbuCPZJgOPtTaieYqJQBgchGfYOCfV2kSvKqcXIVC/ArnozgGXCkkdcO+8bW1
/wcfIDNih032KhVLck5UIA==
`protect END_PROTECTED
