`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKW+zSlOrftdz7+bzAigzpzZRULNZi98RFQv4qGcsgyo
8hg1j7dsMmjNHCNDkc0QKtUftTHXMgQ58qer8LoEsl826EW6CwQZX1RD8nmJLGxV
kN1IMO4NpqyWWFUyObN+mPrcdfk9Hyw6oTfPbSR5HqOQLjY0ZexyVROXKRi0nmuK
c1LWir0x17dLi3blAx4ExQ==
`protect END_PROTECTED
