`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI0WAbKARKgfrrRN1vOOLmAgt4Z66IO+NU8nrbJ2C0C2
hnqr+tDxt6ZKdaH15G4IeDXh1hSFa/E2bnVlERPDv6/yyXUeg5lIQwrEs6IxrWXE
cVQwq3EpMf4qkgvD16e44NV00Its6W9cNDTimEtKumVWI6+N2nLQGZuDWsftd5De
+KNNl8oxLdwSTJ9hSITpsjsJKbZaKhbnhVixv93yLWUy3/f0ZotccdbLm0OqEbn+
mCWZFpE6xXe0MNnp2e43ns5rMlHRAWX3CpDjSQYV5hhg/a6q/Zl1kGhZmFKo2TeK
uHMemxHaUyUii+KPfyIDlNnPfMdrehcOmF8tW/qcJNhGAFnjJsEdJiIu+dGLNggj
tMa7XCEbqvnsWo6jF13/6w==
`protect END_PROTECTED
