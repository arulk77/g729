`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePyI4ywobrRqoWf36VDH9ZSegWbGwY2llKJNynJyvxox
ZPI9HgRToC3Jl2v8a0+U4DWmm4KTn+9hXOSsOGQ5TxZ2kZRV2Iio4k+AXUTLwVNu
PColY1/i++HfyNukVL8GK/cMnjzOfgb4BJ6VHEdsaHs/nqzWDYaxPWBCzevdHeWz
hQZz1/J3JHk2aHFQnkTJEw==
`protect END_PROTECTED
