`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mwB2Wpdl60+SScHSRBo9oR3cuDq2VraoHBMBk0KjfxlSBTaJcfnj3N1vJ5a6Lvqz
KOr0eZ0rC3YNYfVcdSiGTwr9LmlN3cupwQms21sjHDYmQFTVTHB5GIYdLXLL5OP6
`protect END_PROTECTED
