`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHJuyDbXz6kEvMZExpUfnCMS/wKJVPCHvbSqCki1uvtG
HtwqKsxGNokxy7bUeBIIClzwH+FpmIffLjj+DdGITee6o0ywr2zrucQm/fB+JZbl
yI6jhqBklrXUNKEEs+6OwsivHrh5GQsMS2RyvHQVtoWe8ND0ob/8QslhJCgdqxI5
mDg4x6yvmZ7bIF7vVhllHjPGn+yf6MCW7srRM4DO6twUEMXVHDPsxMNTMGHaO99b
vbtArDsoLeDb3v15OGikhNDTq67SxD1Z34TiUE3FeKoOLjGs0hmH4YQOBglxVIGU
1eshcVs6VtKDiL2PEGO2zjZq7bADaHvAmqbR0lZQvCJHLg9PiauClyzZ1uUZNR9A
2iO9cLktNkcOWb8a9TNW1YEXkD2yj4HVfWvbr8rRZOmcGZRQl7OyK7fZFmXAcLX0
f8MlqO+nSOJwas4LOulUW9NgrsaC9hiJilOyogQyc1cMax1fprZANNAHrsNByUcr
2/BIjZbSCCURiW6qFOJNjQfDRfG/eO5pghNfDgM7F4KLaDKsMUwHFWbw+PL2Tk2c
`protect END_PROTECTED
