`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMb44Uez29n8M9WfZPysu9dqYzUWJl1FE1QY7nhmO6e3
gWTlutjCgGbHmnklG3TZtcs3WfAMgfXqqFx8BlkcJ2KLJzHT3yuyh+y9wsIMGujD
XGu5KKyMZ2nQFubV4+WGs7kSQ4d/ViB//fzvuviEsSu9uDrPPtJ3UFSRkaLrJYP/
Aq/l7Vy5/5cYqhV+LldMedsTFzzWpCbEZYPuHxHCg3GeUe5dRoUgR6suN3J3wgzp
Zm5WL2UzNe/h2nZ8CMHhFm7DaQ+IH39mKMQSal8WlyBRiyb03eX9wNIUOF3f1xZe
yn0XPTVOa5gEI43M/4GtFQ==
`protect END_PROTECTED
