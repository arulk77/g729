`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHlX3Gf4/x5LTye5Hh34dYJbB02cmJV4qwG4oGoqe3Sg
O1PsQRzhN6QarLE4RmUagrKLLLuJ/6Q+0FOGNpnaDDcaBRaoJVK/eD0wo9sOqeB6
wDwz1k5IwCyxANWa2+tgLtuUg7k5EVnTZ3UzOvhSow68UmcSKN2i0HzgAD9zW45U
cfw2Ys/cDqY1iucHEUgzQY7zeJYWIERihWLNjl1KMYQBGoH8Y92RWFuFfUHStggg
`protect END_PROTECTED
