`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL82saVUn11JGTcvqHvbC263uV3e4TmbnWw1JOrpGfNyof
sy+HrFI+JZnSrmVhcqlJhATBsoN/sJSPPLMjabzeZwLyjefrSZH+aNM75y5k7eW8
43/qekuGZjI80MuYWlgMx5+shEbL3Mv3oqs6azOMt27S4i/8NRP+gS1Iw+s236rN
i1B83nNqURpXMfklwitI7lE1EGWd35fXBjccqGpdHE3dN0aondebdgYMv2cKi22Z
+OHw8J81IUn6Y7u0TwP0THcfu4MCFgQv9S9BH/ot1OgJ3XOFPyuPullTNI2ocM1K
CyPaHUcA08TCtbj+SfFim1yyhxP883LCKiBH4lXuin0AaHzuy4WiPVUfUPCr38lW
DrSBzePYcfLKUm7rKav9iNjTzMWjQ1mSsz/6KC9DYHj4pvj5jz+50oo/52DfvkFx
x4dPQ/f3KN3vax0qTyb/NecB3rW/Za9JmaWq6M5COhAAAnKr5JzWkLd0uvO/tfJc
XqwwScNFilQCPQ/pDymFIY18wkpXtax+LaatG01dmo1/0yjOMy64mnNTN4KYnt16
DAqPyCTnJljjmmpDDeIfAYBClpkkfzThY4Z65U2eFnKX026UpPHZwyCQeoK5gV6s
F9RZRRyq3nxzI5o14ZdSMG0iLT+ppSYuQO4bG9lejfQLB/dwuSm2xB9o9jhHrpc8
a234pD09LDskrqCXYlc33sjP3hILVYJWWD+OsnyGtfwmcC2XCaQu6XKTfhVWR7dC
WjoJoZeCYk8sUcOcBUlCHYWcfkREobTa0a02bze3jtjf1MAW7ZSPbg8h1voPVLjM
Q4AELuUIM3fDZnkqqAd6keuqFQ2cnvIoowivnZeJLBtvj4HLqq5XBr2vXjbq2+GS
kODX8tFfNzX13cJUqXJih6coH4QveXqXPXiOUpuL/aYj6QtwobyT3a6skGEkbR+F
2EwiBeNpY8GPKKQCFEAlow==
`protect END_PROTECTED
