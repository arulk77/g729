`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
f11uP3tAS38J+2XEq2c6cEQ5BImOWRyE1iFg/JKYC5LmgSG2QgDf3NHLuzubbRmC
BRvZ2XxKqPckazKvNBJGd68iEROKHWje7Gf+tkCXSv5opCavGFSYganXWzUL54DW
qlx5D/JWI+f5kCOPSt7OpkolEGeI+yXvZCEZPA5vRDn7PWKaesPB3hUzYpLvm44q
SgDXkpHUU3hSH9AYcrTzerNXmd7Ur0Mx/khXVFhxgp1QlADD/xfVrIb0qpbLtYvH
`protect END_PROTECTED
