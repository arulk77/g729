`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBjIFwyu0rYuId5ScqjuE5CInjvOWrNmvfLvwtBlSXCP
9REarGRh2LVRjy1preI+ram2wLNe6lGcpr5Ht8ZD41tmIe+zwYY7Pm6Zm9FnVxyw
33AtVYn99BMUSpM4VlVTRMWFof1baNH/M0LmQJ2a53ulaCV4Bu4p8w7okfqGqhDS
4TebjdjTf/gZL70pvf6Szw==
`protect END_PROTECTED
