`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C3D2DkCALfb9nId6eqKFwSj6QZgZu5vdTiwWfOoYYppk
IcbSaU4ubeYICfwSAhmldQc+jV5UWAxOxJln3ZscLlKIFG8T4TQ9vuZHt49nr4vu
Rft2g+uNlSSxTE63QUdsHa0FGqUWvyVzNk683Shbddk5VorLkRos6UY7I5OapOnL
/EQd9oY0IP4Cut8/ECqS0CSsOC6BytAuX2VoxfIuM1w0v8qRjUBVH0TFXHj40qdv
51iK6GEUrdYHs7hHEWbty89jC7o6GjLPjM7kq3nbX2RICvtegwGmc/Ss8OE/AyrQ
654IaH65kBqAiR5EL2y+051IXL2/xTzoVSy3anx9WorUhanx0oXljJoofc7TPY5m
HvWFamyto2Z+6jSUE2Vs5hXAM1nYLu5r9KkLunjXs6dFA5xGkhK+m58K0Wk/F/XA
ydHb/hqxYYZsCtR0//jh/Y6Ve8g5xJZIwHeFJkjQ3PZbbO85IMt63UdPkgAAGpbI
V1/2ElR/qqJIMEUr0IYK6i7Z4SES1Zz3aZMD523p+bUTZfdlTY4Fsw8ubhru8p5Y
kgFtgbA8pv6BOgQp+N9qSt0m+FxUd+RebOoAuRxea33n7mio00oYDj5LeVZS6jFa
GrI2yP57bhEimPs8WtZN1cu3H9c9/65ED1l6fp3MpVjR/oPXShb8Bbm6+enVgUDa
ExDlzuRbm0VHhEU1DbKQb4qxXpb7/5gGWqapovG9zt17brTGTiYEy9QMZF8DztVB
w4pQMDBlGLHvHoS0b+oFvinhk6zg8fAVBR2OqY4ObFJM6q69wbyU6cdJC4K9y7Vg
qAsrpaAnWooLmBz5wpRqRMTXgxK07fJeJZp9OaEaz4zT6xVlXm6AQ1FSDHS9s/8z
nkJVfAi72mOYbT1V4LNhmA==
`protect END_PROTECTED
