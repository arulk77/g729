`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBhKsoX5vzvxcykUQumv4ytBeY0Nv8ZsMHoT6hDj3kQQ
U8oiKl0we9PJUzkGAVOrjKwHYHm0I/tKNHJlz/4KT93TRd5YULETl5AuGyIap1fQ
VLp/FHa09r7fg3Iuz3xDjXvE/H+diPvE6Nb5PUORRDxZLLNJOSGJo5MRLvdFC902
g+dvxdaRNfOzC+nWDKRwLlC2OFKl+1Tlv+wmBEthYno=
`protect END_PROTECTED
