`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMJVT/qkNo5jZ6fyWdKFn6XGkLKZ3chs6P+ZZFMCZt8q
HJ/MoRDZ9XPiMlWL/zu3DQ5RB2sZW85hzW6qrz0c8jF4F9GCF7r6cP1t8roHmuGU
ruxFvnn+OkcWbOpu0p5okL6PiADJrZzlXxUcyszX3oAfvvYDCal3YGisI3qTXqzv
JgpL/G6GaG/XYrhdcl7WKTMChv+ENHusJkkPnrFHWfpHouJV1Qr02OirMEaO/XoO
`protect END_PROTECTED
