`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
FYwe7CYClQoMxFvKx5Bo1aDJ9/9+gtp3I7I3rjX+fRUAnUPNQwVsGjTh26Akj6ZZ
o5vpGBCiZm2QwanBS3Aa0CMIqLtQIS/2OzE5VSCnkMEr2nElMK5PHn+/C4Q1c65i
nfQyJ1++qHzqCeFtQ7X6dWx7Jv6BF4ZR/tqkUm6EXsntrwRfhyh0yeLJ11PrD7xW
aLF8M13thKV0CRbJkf8++WSr1VYK8w4j206J5tqRv2o=
`protect END_PROTECTED
