`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBOc5hc4tb+puVm2IUV7YZOZfAruzU64i0mxsnYTVA68
QDBS+1o3klVIV41jmULfzqLMHNcN4zAXlgSb2Es2wFR1B0oeiefniptfkoTDN7iI
oWBpwFBK1MibomB4fKFoDDkzI2XvcASaFZ2j4lqJXXlm7i86Zg5nLVuJaBZJcdun
6+pp5ohvq0/BocQAHUYx4w==
`protect END_PROTECTED
