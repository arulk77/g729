`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SW2X3YCVsGZVn+F/2RGpq7mljTkhxh5KWqZXdOJKDR/O
P+li577S2kl9ZZ3I29QadU3NMqxJes4IL1fLDeSV+IzTghconPjkpZ4lQRPtITn6
qIFgi1fuCGU2zQr+PQiooqtSL8sEts3/gsylRDy09RPVq/h1FbwiSK9w7MTO+SSG
`protect END_PROTECTED
