`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+SVrV26mTByZDWi41e4mdhkv53dBYGdIrAeiqcQ7WXd
2W3HDH5qLy0gDVLorZodfOs3Ru4XwAe2+FwnlbpMF9/mri5vuWpyeVrG80nD+ehC
TKr7iw1X2t3BcNBVLJWqsU4z4nTAM9vBho+4sj/+sFMyFcVvqjfT0ObVq80+VOVM
b3u/J3JznjM+JcwQf+P9sogfK/7sgNykeUYRFmBA2mjHFF2/DRaM17PAJMK29jqS
OKMbtYTQOq7kk5Z6BdLRAFagNOVuzif91PwZWlwvodCMzzANIvcRU++br2vVLsj7
N/4SbXBJ8RQu60TSNZ0H4A==
`protect END_PROTECTED
