`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
h/EFC5Q1tToLqVb+URaFYz+u44RJCgJphPPJ52hkNaso73A7Orixgn4ynqlYBGXo
4ReScQapTM367SiZ0PRh+fLFnW3Vbt3D5uAF64tURmRZ6jreGrqj/KHASp3jXueZ
2hx6WbOxV5qdCV94yY0TucykewkTA5oahkLcqq6BS5ixwucu3luihhztXQrPgY1e
9CPWCvRt/3d/TGxsBEsIwhz+KZDqIY8w6X8yd8DvgRtcdKQf4ZFDdfWvOHoHQ94b
ZSlogAaHo0GTcL+IYIz3jrGJmGaDlDgbguufHdUoExWq+J2tgTJ3hFygom8P7V2M
W4oMftpajJKeT7YflcbKcaaNZb9KNtUj5WNIDxvFgLmLmCoAXPpAK+XTgYInHnuP
iJDUS7jRxNnRWhfEiA8BGMVa+opbNaBhaAv5NjuO8q6IgcUNdn2IMoiBiJsPATK5
8eat0fEic96yDaqEeaJqkL2S/laPD7bwnG1iOAaJJj+kxxs3Hr0z21vtaxUrthOh
6eLYYaMqVNC+QsTakYmoN1TDC6YJWbYMMpPoF/h54JhhO4uY3BUtSBhjOVsVsOYR
w6zi/QykqFU04SpF35cu4mIdzMtbdN0ws4o0AjSVpat/2J7TzuDn2I68Oi1DrB2e
tOSEQzE3iMOt3Hp35lM6NfOm/hglymxBFiKzVHjFVvXW5RK1JfvSKAAJ1QTRAImv
VsKhxD88Gc5PlQdYpFWyQM8E7npTjAoxJ5ZkCidZOT0+T3eqIh2hvXE8Wf7XV83q
ME+gxGmilu/xWTi7Ghb7l0fj5n6ELN7DTm/qDT0EadMcQrY80DKWBoNt5ONZADMG
wMWOmFnoTlOtkP3vpTnZIdtIf4LiH4pZAZNxZeL9RAV/LXuNlZd6xBKw/zXa6rbt
rY9+7ftne6mvyHjAJOtmFIGqkxnFWoZ5BBd3WIp+z6euVI8qmu0MbPPlYBZOf3yW
T32YgCW9m3xjgPjAYXjWOhNiNtLoUjOcV1N325gtUZnGrSR9vTxcsDC5F+RnOxa3
yH2ifd+FQwUdcIhcBZdWA2Isw5xEPRu68R+wFFuSjyA3Q7gNYrUOuz+VJCy+3zS2
rFGjYznIvNXCgLvnTnpTBDIVpDJewGeIZmVxcWBmsi5dlc09hBuil3WzBpXd9Lxt
Lc6zorYSVo5IgvTF1rJEneigqaRSTngOAro9EoTL8J4X9CMBuLRTF36DedHJkUIt
O/vSIsuT1U0qjNR+lfw4VbFW0rvsULiaGoHd3L62kzl+u+okpCKa3soXmsaTE53N
kNhsCbbJHiXFDylqz2jaVr0IS0lRraJJZvKPC2ZluN8ddGXwQ+oeIEWXRiekiX/A
TvxxhBL0Oxbhwcc+uZ+acOzOG7XmxwL6kYfH2LdYvDbM6GkF6GuDOimrB/3Lw6Hk
OOCC+RQnqMXMMNgfd+7KwZSunzVmv6P+HTVoQQk4GLNWMV9++17qN8bdzLPvW4bf
0hDxSMcF21tGOCwbM/vMTgwhOQBxcZsP/ddgea7FEcs=
`protect END_PROTECTED
