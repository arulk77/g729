`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Xd/07D34UQS5uF1P39YMRPxTSWrCBXGkzAWxwZhbiei3aYzLv7ANsoxjOqFw8UYl
h8jatovudyRHbc2fwjEZozaz0zWb0lza3B2d7dY7jf6waU77KlewH/tEXvD8vSL0
oMMlaOM9Cm9LOKJiJNbBFn3UlWHCynoDrcy70joxKKcKa2dVwgM3hZMcXpVW/OR7
HivNMKyM3lEPVxY1/AvpDMbzYpQGhuyw94jfUwFsTWwORjLyis3BF9P9YTkFd6bm
FeCljHSmBGKZmVeMVoPWHSvAkHqtiJrzdG7AXHcM1FZ2aks1ECAubZwMFYexehXr
`protect END_PROTECTED
