`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveA1jm1ZBSR8Q7+LbsxVb/neCgjQ01qnNdHv3Y8fYNkSh
Wy1dF+pJMk5Xprd7LdYw39HwFzq9bFYYQLye+cgwQ9jP/DtuepAD5YoDlLYA8Mxb
YJseZNxCMyitzRvFwmUmWQ7VU/TaI2kgC4XT4IlBQUW4r2zBjgsq+/HGH07uz6Gq
IXQp0Uuncz2uvskxyEWyJ1Fga22r8qX04s1CeK5U3agCNDFymSYabDb7hpDIGC+B
O3th5vYbkUlOgj9Cr/CGUpsYDUJSm4ufsq+xykN5sXA4YhrWfEX7Q1EQQ8FJ0kxr
/vAj4LcEBpMaiJ0l2YSFs2UreGOAHS7Plu8twldWUQQ8L+30HqzjDTqr8fMXlOpx
v4aXUZM8KgrN729ufAd/wsnmG0Y+Hrd2hLj3FfFTA+LUaqTktXXSpXbJ1pc+irM2
7L7D+6CmxjZkaxoUHryFcGAix1IJ+0FHA2mziq672RTkwBUfI5WLM4h3SKsvNGVZ
lRJ4YCw1B2sg7/Pa/AfCdq/T/VbmIUuVqYK/OAMw+xMXCMG5n263j0UYIUb3G/Hj
wUBPI/Rzes1G2US/clzxirQZbsuFvzZVdkPGOmmYfdBFyHDcte3MJwV7cRCilWF4
TC7IWMDiFujf5Vt/s9u2cf3ZFuIMRWkxOaKSmj5BETxf1jX4Ztl6vcgYrLhvbuK9
0+pfP/qpUg3hkrMtrKIDChvz07SEkcaoIy9Yv41gCIISLG/ySvrAc6m2MUDHxYAn
jHGFPCK8BhpwSnwTYsJNyvqTFmcIUkseiE7IfwnGSbwhtEjHQ00MXosZ67icshOr
xpKYdjuOqKJCbmJ/IscL1QtQNaxQXCzvomJnvKJvpDI=
`protect END_PROTECTED
