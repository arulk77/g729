`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL84Rn04n4zGPdFj/Zt0tQEbz4WqmZOJ5I2TwV0bohFhe8
X4+VuEHAraEORq40syK1Hq0bf9lHSWjioMX4ZucXU268bWV6iTpeocEfAE2xZMkn
LQ605ZMuLDYj8fUOmPLOiL/ac8zRT8zAAGTBMQN3pca+JSPc83/XCA6FowI64fJS
yMqoWQ7vswSSi83JrtHTJzcCSN4s3GTJk7trU5fDvai639y5UreECv/7qO8aKMeX
6k4advKHhjhhWwynQoV7NgL5ofYFozXk7pPmJ4O7CgGwFD2yWZ2wZdtb7DYGRwKF
tHk1+cJHsGtTicrKGZiExRpcayuj7kxiCw8ZHUnY7CR97949LaKYlMkrCsr5ElE+
ofggCroT9GfRPxn+LkMCns0Hgzkm3lH7pF0Jf5Xxfn+bkh5xmupnn9rEMbwVDwm5
mC3gpcrXAj1HazjkduTW95C5llz+zT2TGWnJ4LYotgaH8M+cYoWNU9U7xsBlatoQ
Zep6pBf6YyIRqy/rYLjLHkfILoNtrC3EXKdeWKEg0S3MgRZtJTHZsIY9mbyh8yNV
k56Epk+fFWbfZbY/j5X+ggouxeOgVpeGpt+lRQ7DGtK87eBF2yGoZKWNSH1byo7w
G6oZMwItE3YJg8vyfvwGM3MycGaz7KDF+j/0dQnBvGhTTAuNGCaEHGL/LocP6oZy
CQo8nt8qjm7FS5qav8mQkf/QxgTboq0H02IqR3MBdQiqfpI/Ecpx3hiXdW/4rk0E
+NSd4SopB4iUjMzCuC/toZ/QLYOZVIdRBMUZPNopdpu6jz9nk+1BQuQtwtkLSfGU
0OcEjsfQnM2Di4Y2+T4vBUJFauM3VoGfmNgnG5zU0kI7V1vx+A4cwhxbbMp4ZxnA
bJ9rFePER6PkBrPNkFjYulT6IS0bIZ2N/bxsMTQU3+8Xoi650xOgzRTJ6qQ7ljQT
aotskh10RDwmGTESGwGfRZ0Tpi3ZfhpE3vryXBjE5Fg0aGEJjdI0G9ZqjY+rYgeS
UifWXTArtGYkFzWsMF+Bu8afbQnG7xe0McaHvoQE9db3ABqxpJhCfrZS14hwPeTE
/+p3FAO2seEa8YPbM3sZUTr3m+snzpTROP5oaKRzWapTNEYitItAo7bX4y2Ncuos
rofbGc4Tjx+IbwdDEjDXKg==
`protect END_PROTECTED
