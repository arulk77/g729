`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEWd8431BU6WkVfNSGFC7jedTJRs1Tah4j0wZsY+g6yW
43DPUT0Ocsgyp3akO1OMoBE0Ma1+AaPgDplcETppjiCVY/HyyLxqEJeCfFBOJAHd
BHUw1AVD1TbDJ5nvnCN/fLdaBEczgVPGzY95XEtThvMgdg92jFMxDP55p2WrKvA3
j2V4LjeZ6xGW8Ggirx3hlOYww3tg4PgpZUr/V0quad7ReCsTSSSNBKD+c6aeESOt
`protect END_PROTECTED
