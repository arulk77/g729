`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMLmiJu5QOnLCALUMNpVn/BAAdnXukaEXjLVC6ksQNIn
p5Xh3sCGSrrmGOoymaXzMR3oZ7OuXu+IQLovJNB9tPEE/cR/LFeaC7gj5tOqPGZl
9p3C02sQnuwI/nZjJ5XiLmActwZgCYZSvVVU9VV9v1ytn40dDJXWd9G4wuaDydT/
8LsYtpK+aWC+RPIvy2YR8F+/YJQfVrSslIPIm2b9xLb5Estwly1o6cNo2oyC+9PW
QxxxqHTbkMMBBpm6GJCvAbeeLGC4n5lpNKwd53PQK0/FCQkZByvLxsV63q1AoXY1
Ph9dScr7uxzndb4Go4MJGes8F4CbscMCehUKSzWXzvknhueW5FNMr5/5dThMrBcW
Y3+LBa/1t+OcBPtlBY+uLHu0BaT3s/ywlQ8crgnKugykiuTN8aX3nxW7T/GQ8Kcd
dqiYozvqalzXPJtE9LjCqaNVBvPMu9uam/TXsAHm4qI8rOJ1Aq2poFZt0Q91T/vk
uEtzJmHjbnlUDOODdxA6tEBZ3NrZb5ygtL9h89sjtjmIQpUFLGEbQeQqqrlb44LE
jcawYgqawTmUmpmtrzXCy17ZNEchNZEGnPziv9jCsAWiyuP3pPY1OkpsLU8L+rLt
uIiQz9FJ9K+J7dSqH2AWwCRoU+MIU0tEglcjVIJRZiuZM7H11ow0+/bCmBwGtlBV
`protect END_PROTECTED
