`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG5TyrNfkH/EZTjZNnbHnT2lMY+JH/7jyb5qytI3ucRI
mLqXrc0kOH7Uj3DDNp9jQtNQFRIqOcVuoyvezcw441nnfaTzMPzi5APrPN+u+ZCD
mgcJo84CWINlFY9jbIVHlcY994O/P5J1jT+kTjAkD7wr8ar+bSq9NKJN1U+Qrr/E
vQ0/FesYO/2fj1mlH0ZjyeW4H6fXFqYlWgULNyi8zJl25/a4O6hWNK3e2K8NXlZF
`protect END_PROTECTED
