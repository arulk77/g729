`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDILLGRZX2za1RT4iq+m90tAO0KLTK/KXhbfMWxL4GNE
s3hvIpqLPMSLFaBb1DolwX72lqzSN8Pg1Qci6ZMZKLePk2XIP/2tUYBD8VW2pxVw
ymf3WpztCjP0iOSgX/zDUbuTpb9saB5roUaJ8z+JA/VihnRyKlrWmWMY91lSlWOg
RI9gH8NpdH0L2tVOhpcUWN8sIG+pB4Fr5t4S3pR9zqpE1Nsqi4DWO8JqhrL1T6OJ
kEkBuMILk4WgQAarOata1PuURrCOWzOP+kdhIv/6iMa9p5IDhGBynwUSwgZNqg8Y
WOy6iMiNkBWcSQe1xPrNWxU/G0VxYBOi6fEAkLovAOnFpaNrOAFLZQ6QMPAZ9cC+
bHb0xyQTwEkaH3DyzKQgkbnaLxpgUj921KIcyQwwsDSMRD4tnd7MnbjcVqv4x6x6
m7R61gMm0wkyGX5UDCcHy4DUHPP7q9cJ6BuuOnz4xeBay7cREiWqEPokrklrTcRo
57kQLnxq1iQtNRq1ZNa8TCJ85gGsVa3WDsDDtgxhFeVtKTZhUrQXJbGfpIsuHTbW
TmSwarM5sRtF/kVpktfkgt7B4xh/gdP7g4bm8rCRJFs=
`protect END_PROTECTED
