`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu463l/hLA4HpjJFYTaaO/kX+sR1iOMsiNfmUCiFHmfUw5
MVQWt41XWyy5hcAg2aATYoZvnTYBA6eKX0+epQC0WlIZe4vfgIaIaoNzZsioq67y
yJTfWyNKl957mAPZ6npekb6Jtx2t2oDt3SUr9zyCDFw2je9YSPP5dMecpoRFurtW
ivQdS6ksvSeqfvkYdwulv9t+th7PEgeLRXDOnTDM24Py6mjbSVSTAdtFx7obRrD+
MNg2EIerqeYLFoV7iT6rMNMMVSIAkptWUSLJv2LGoI7LcgoZHQRpIxLdYIoA9Miy
nHqNdiOVxG1OOvBKc013rg==
`protect END_PROTECTED
