`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C5+R4cOCXmU4FNU6Yz005FomDBeGEQEgHRbDzVJciwlY
tIfQt7M1p/dBCqsaDORBGKabuvzqUJ/mKd9Cjs5q0vrPg4TEm0QWVMQ566n09eAh
GQH52n3PJdyJk3quEzdpueZI5HsCGuqTo9+uh9GVcryrw8ZPOKfd/frH7fhA4/ww
uYkUv6YZueFkTjq80Ocbd1PCKHJBfwDNxXQeauPpAWsENKXstaMzbO1hCc1m2dFj
g7PoCRJlxeOzwPl6cMHr0XLrO1J085oVyuvxWoSMh9mGQTFBV1n844mPFdX8QJ5q
J4nx6Rlz7TVwkqtjyczM85/SMxpRj+PkjnsS1ZWPDl4nVjAhJA/04WJMKPRfTYkF
XFyJndMYZAdX3MF4SekL8kekyXe1YaHvGPy2G3R2tpV+fXieDceRonbMoevfGqz2
Ojo0Gg1+BCIpIL9cHvBuz9/YG1K+mZLgL56O2jDUsFrSeG+wsb/o6gI6AQbYE0d7
52osq1jDRsl+xqDe7ZqgZvr5bYywHxXipLuBUjptfqz5FvUog8A0Y2uQmFmQaiy8
m4ydtXtcHwGLVzxYZV+pHm6+q0Ugtojd/wLqVosA6Pzwko6iWb1664CKaZ6qJuij
v9ZHQ9mnSsIc/bIQLypd5QevDTVKC96E35gtSxJik/ShaKoUVCoqQUe9YPoxOweW
eyxQmFfwUct3dovLWFgB7Osfzvfz72AsbhXM3qdJRj9nbFauakkDPhYqBW1NF4U6
8Nms7OTc+IJvoaL3GMj7SUzn6yZpZhBXe0xS0LL4tVMIpFabEIV9DgE638/ZsRdh
NIyK/WHZiDs+VLO+5cbyfuaqqwEK/wm7KqadMvqHmNxEHDeQptrOf5TiTJjwvZJE
legUEJk2TkJ8qU2zFXW7+1/FPUHrZppoNAflqSk0WDsT0YmghAStk4iNxVfonfWY
4yti+as6qLf8gxhTM4QnPZh7tS0ITPWELXqKnjW35dUeEotbUFVmGDXIJ8j+vpoL
BaMtcfzfjfw2uDQcFIza2n1y0C5Orh+D4NPlL4K9iYSgq2/vxZsFq43SvptSPwXq
3NWR7Pc1ePJI2Z5xTlxeKO6bdj140YXbWNElV3szSCTDCzbpmsCrfzVP/sU/gzp5
YWu93Qx+LdeOqUKKc8b1Nlo3H76paL1Po2QCYftImwZwRPgr9QX9v5GIaWQwyVnE
+ijGRjTPbx9ynwzUUbKMmsfkSqTPU1va+zr3GNshDwrefTFXXXXlolcgPUmR5UGv
4Iu0gbPFBvhkJBo+YbE/SFL8m/uDfObndwA0eBBupy0siCzcn4wxTKswgXli9Tf7
TnQzcVSlFrrwK2o/7wjy7g==
`protect END_PROTECTED
