`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/W4Qe0pORS+7JSrSRQ6oFNNbRTXJZIOdPS3NgNNEfK5
23RUvSotuVHQCfXW92NFizIMxObmPWNthAQTtY1R+WxraD78OL3G+VZpC9AApWPE
nMbHbvKeoTSZF2VOV/toovshDdogtheShXqdb+s7vHFo5lIBMHZNTUs1+dhLrfmN
1cnjLOtcloP/KwI5z4c9RYZGJgsE7yicqZsVnJtEulo=
`protect END_PROTECTED
