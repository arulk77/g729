`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBtciszTs0WAuuL5OC2/ob6/dhk1T06LsIIpLjwJXuFH
vkpAU5p3P/f/M+6hI2MIuArz+qugvDN5mJN41ppZAKICt/sAm2XuPjqmSaa6aDLj
aO6Dok9EvDgcmYEV/iR2xo6zvlkCmjQeFNkN0QB4tkfooW5fyJkdj7hkO2HbYaNn
`protect END_PROTECTED
