`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFdLz0r4yh2BfQe+7LZymeE64ne9iL348TPXGukdM5hZ
wViv7SzNvvzAdGVVa8y19RcEUc7ZXERwrOBmx742zF87AomfmWSBCsIyxMPT1XvD
B0lhVa6ezqj4pdSu8XJCQ+0yqyHTHPOVCig8f6rfzQMch7xngsxzeYU1Y1JgZTka
ZSFDnwFWC6H+pe3LWmCdAmBexoFUaaFftKCuRbXx8KX7e7whfRBPYf+61Vwc9Yux
`protect END_PROTECTED
