`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKNzJVaVxsqGvkqmzt3f/TMCQRl6DBAulND2G3Q1vHnc
zSmxwfb5s44nE+ytxCDCwLJILuNs/nVZy0UvM4GzK6jKrnH3XjT3FWB08rS2rvKI
ONYhEKZeizum5CyKFJ6WdOZ5UWsR+XtYx5qXD9Kk3vwQdnblLIQQEc0Z7fEqp9SZ
ZS75SRg1z5oxLRYfd1CBc5l7j2E47qZlCecgXQBnHsB1HZnaw1ZrssOjFPQKWtCg
mw+0OLPID2Son6i+E/DxSNqM3spCEpUIpFEbFBL1eD7J2FHI7+9S4L2chxO3v58p
t/VlvksgH7BICDJJwkQ08g==
`protect END_PROTECTED
