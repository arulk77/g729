`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
qnrgCubmkE9b3+gKiPJZVW9jxsnZt9XrN9PsdxtFry8Ytkze3rnc698/8ZS9c0HI
EExIn4IQDC1DUscfkg0H5yk7s9VqYyrwG/rPoD+W+G5WXLu8bB3E3CFHMY+Hg8HA
vwlkjBrPmg6dDjtgQSZK+Td3YcT5VoNOgOouFKsb9peoUDzNIb2oQdB90xhdB6iT
aaRLSEt8lXz2FFe/RiuEO2ENh5tE88F8Ud/HV1EQzR3AIjbS23K3ZorFqsVuNn94
8ssNzdZebp6Q/RrRSzf4iVwgV4TKue+QEeoJ0qD/23o6v2l0bmLZX2g/dygWOHQX
MVsXpW9yYxsSrTDP2q9n3i1AeWiRmgDejN4Uhwz69j2c3bRaPae9Ebk1HBFAFfN2
LE0PdfZln0gc9408VZBVNB5ucGKFzergyfwtP1CxTaRVbJreGx+cXW3TjScyrXm3
apCnpZ3H6eWRRdWOL5w0ysw6awlNb8sp4nZaEIqdHjMkpubiUR9sbPdtG5bjgGdJ
uPeJQuiichYicCTw3VExE1tKsZediTFXxfvyE972PzGJ8YEv34vkujRs7QQ8Jb59
yrSJQQTMkCOniO/I0RrYtkHTEgBef0ghDDOMUjtvFFCGGhx7xwXCVMboEw9mG0vj
FIxcr/sMZxNaQKZBsk5VL8LI4GaYBIJGi+UzK2051bg98B/bR+oYOS5ZwIYQ7eOX
TZJv5MiX/h6y4tiX1ZpbEQCqI7CjuYqO2XK5rLkBbfWR6MU2O+xfJT+Muj+UwSKD
+w7f6fcsA0s/tu7okMmu8DAX+9ILdeqOGSn/F5w2JGYHRqsZuTSJGTTRf4SxSCPa
Hm6Vul5wq4fCzW6d0C1i1ejOWGKh9kel4V7qz/0lvQVh6F01pJN1GwKxpx9wZGm6
hqZUuNluxVoNoYqWgTHtN89kvBQXWuxvhm07/cEOMRe+3Yo3h7ajbHVU0IQTOe67
1x4x4BNKTEo1+4r2P6HMrTwR63x77jEPvIKTFa0FqREUvJ9+xJY8IvT4D85XuxYh
LQi5on+296ZfVIbskZarftOZ0QhPep/fNdz1kvS9Cp/PDhBciVJ+2qfnQPkmFBTU
tqfuhjmLnYNq85hJLY+BmXDDrpHp8QuN5tzTs2SU25GpPv5bDnYkyuHaWshHr+Pa
i6356JlO1SQCkpYTK7LCrfyqa+5twQZJB/Y8KuieZUtClMy2+AS2Ql8FuxKtHngH
zpSLwBaCAltQjmdui13Cweq0+M8fDUpXwB4gYQXX6rtGLofzn6T0mPQnBECXEZAm
mS28PVjGbv2tdEIvD9PZWLiKMLOBwz4lMMJiO8PVLQ58kmvC/FwqMdSCTabS/WCH
F9WgaWusjUpTqzPO9tWJrpcpXJ8aaiZ0J2wpy/ddsO0/fi5IAm/1/8aBEPoo2MIn
//JI+mfoaQCuqkK3N4Z3aioQgIZJH2qdcboHR1/KeMrbo3wG1w9Tf2KGn24Rd+Bj
i/Rw/e5Ol3v2zDRvLTzwefpuULQfil1VKVnbmRZV4QY28JRcBRD/UxjjsWW6Aw1/
N95WI9DDZM1OsvGSvRI0V5+LVZK/ZH8gSraU2P0hsjZB0QETHY4tPhFOE8cIOJS2
vrJBbIQq6Rg99MReVcHJKUqvkCdslfu9nNFXR/9eEQqcrO+Kc/aYTbD6pudSRqyg
PFliEujorYPEI2Uyrf/1WblGNIllsLTcuY2uwxy6x/cT8b5d/hB/EnWfazF48vzi
FUVOF7rxl+L6bZGU4MY99+beW7XdvFpu364nbk4c/MWtl1aOLTU+geAon6VOAmDC
FZB0kidJpvOH1fegMESjKjdPOaBDczYFUCoNPCWxUCpKHUC+IPyEdd9kiHPozPT6
a6Qkq9rz6uCnQ1EDPUkMCPI/FzEp2/0LYyxu37GDzmtqo4l3FM/sMoztPYMyjgkt
1L3onXmvEPiZZRcHQ1iMgrUeYrIYH46OuvYjbtMcF9hymspBR22Ts98vbMwSRd79
LDFDEqc30DZ5Z5w93K/YYyfP6HeH231hFkqZH65QfZOkmYxTiVetyID63BTA+4fx
usQErq3n+8HUXleF4ZZNUKz9n+iNRMWcpQLRx6/yGIpIbguAePb3q+iMQJM+TXto
wTvK5Sq593NzEkcUgoOhiVCFUoW2EjaRk3U6QJnpGSRPRgMbMB1SYhedhdWu731S
BU6T2ecGepbhznAl8i9iLKQ8g2p2owoKvjGR5kSNOEpdYWs0QaFgQ3LgTGuGgjxC
LbhVRq6iieHiD3frmIMyyYtKrua5U0mDz0OJ1vL4ra2eZDKs9X78VKZYt4Dk2ehC
OqeLHk+F3GuUtdOm2gKnEfdd7ppWUqAf3Bq4eGI2p4dqOt8eh0viEL0xxrwplARm
4mu1JLQaCzT4dZHA8yLynsyI9ShAeftBP4YcfBdYTlhXV2QA94eCUEEhCP78ql4u
dGsIZ6c+LqfsnB6/VqRSBqfyqq2JNTp9cdGdeZCTuF6yKjgYPQSuQBIE5kRH2iW7
6bRIHDanAuPnfPOcLaEPf0nT7s/umOcv+0Gl6nYydrVtueTcNDgpgDMQ2/cWkOf7
4DALd4F1bAuZeSIHwQVJJnNhyKacgGjcOKxSLX52PTh3bz7kiIo7T1ZVYgtQf2Bk
KDFRsnO+rCzimNZytMF+5K3t1ZFFsHTeJNqE8K6R6gGDGNYM93ELwCGZNgLo6P/j
3HuIZfByN3ukRJlGy/Clk8IQEULR3O16iHPbrNzCJiUO2BKsd9KaiMOemKZD9Hv1
egvdTjuQlr15aT10Hkyeh0Anp0o09dftOHeRn59cfR9PYTCN6SPI6l/ncu7v8tkA
My1kqM4LvDmsD9niTqHONNXrPpTNXQc+5vMSVicQPKst3bSXKybe48klFP11rVDD
p34XoYphuLsL6K37JZF+XwPMRIGthXh6v+23Y5gq4YYfHHLF6fo/PJr7eBfjYHdo
CJjNOOjhtauTscVpRjazsSkB/XHoxt+gGZeqpW+wqcPxsw4NtfwHsxpQ8R2XmRqz
YvAikO01DXKtBf/58i4O7LN0DMMHYsuoHvF25pj7Dn7SofBvS47kWTiF2C12uLee
n0PlvF14BygQ8d4n4R72jCPUNbtF1Z+ltuofe8hQaoJavZytsZjfi1zgk3eT3BIy
AHd6X0LN97xIlbHhi7p1K0sbO52EMrawr1xdCd9NQykWE9rGsQ3qs8Z7DuUCb9xC
LclKBJo/pNxVp6aDT36FS95uxswkHXLQM/s1HglmLICo9sBTERIRQM+FJhmwUnRn
acccHg0NbAsD/CHq2BZ2U+m55/IxzCY3Tjs++euMLsL2GyezuGfFpX8/heQ1HwQz
/aB0tF31W6ZquYAQF1/j/ofB1kmgODRAc+T9RGsn+plCEm6RIK9l4c4fwyzrop+i
LBBINmFdUchGPTgYLINELZRQQ5sWGo0MATPZtwa6TAfAcnBXBGaeO7jSOGwbi7Tp
1xXOfZt3Bpob/Knu1Ualah6KRjXcD7gFDcBs/HCjdVXAMoCIpkgjIp5TuEuZTOhk
msh29senuzMX2k2V+/ffqlDWd3OpjYykmuS3rSHrdDY/mrifsH2TxGHurl+K9uQ2
VQaP+umPhwCJqIxSz+PF+GgGfQ5s9jC3lEF5IDyolxnyqs1249IkZ7Tsg9mfO+k0
i51LM6shrPxxjowLG6/QNkbGAbq2jI4sHw1q/zSCHyfycSvcfqYRJH3hRY91M1CR
+jLv1/c8JELG6ugvOtGFu37lYsTsMkrM/cqrUDWoVjCrX2e7DHX7fb2YumnMY88P
1n6toNcH/MuoKeBxNhUVmxWULRCtWVuq75/JDNe5TOB/RV2ACG4QG0RK1QbrpukY
cVZNeqHlZqYfMprnVlSg4HHw9nI9pW/7pbQ5kcixFT6cXnwZTi8629Zro7XDJPhI
99cqAu6QCJ6WUYK8zV96NwJl9Xo1UDPGHYKfumElkq8ePiosigkuyBq9z5JABoNt
7h5SFtafvGFlJmlSRHVY4NzwFlEsRvQRfbepGAD5IwluRvKmK026TwxIXCl62LAk
7xJ2EI51js4pPH5dJp09PQ+NZDlfbodlPI3YtAnshZ6w6fK1sZQcIoDeK4o6blOi
xsaCg1sYcNFcJr/PCg+qnCCiCeJb6iTUzI5snN5EutBR0pC/H3TNmNlBLsGGTgOG
qlE4JrQyt9YiDB8VuHNAk5vgorTzA4aYYgeXb/M4qYRCqEeQeS6pFZ1oNy6VgxWa
lMWKJBFRV4xkXdGIHg9WSgLqD+PYYiheFGi8mIoHpFQkHK2Kk2dLFzpTIIGOH5v2
QXmUHa/wjT0Haj8kqM4q5UG/2dyKOjKoK3ihDGjQgsbgaEuvU3y7DHWfyB7jfYnm
1uNaEOfUDCZgqvFGP7JzjC3bOv4onJNMopII9P1RFt4vhQoI17jypDmqtHy3oOLw
whUJMjb1kbxRrTUFYTzxTv96UTMCjIO4as/xIwhbus1WRufCantfvtXsWS6lefgC
BOTD2FgVpFJtubQS19Y5n3mFF1PdsBQ2gb2ykiAc2loU+erxXOOg5OmTNdUVCyeD
tZ2v28Urs5Y4/s3sHbeNoyiUhI9GdcvFYlJ/heGJoW4A7a1GwrPgtVLOD5Ej12yk
mh857e+zXE6kvPQngfOghNhmaDNzAMJpAAm9hq/WcL+PE2yb256zu4gi1kM+RvUn
tzx5sFxZXEvbwWDr06+uFsIxZSxc9Qe4PtomI5oh2u+TuMMkQvk1sVeUUUAy+07v
n5oDQ+idD4bua4HSKlTrUcutJ0AP1Mvvo/GLpK2+PHXSRFu6rchunXmRYDNnFLCk
gcX++NevQ7nrmrF5ue9+yFaSJuWY1syfFicM7U+3SggmcIAO4M1SXtsHFQg+z9HY
ZxtTQ4w7Oaeh3+M4i30tJ/m1sB/4JnOUtEK0UXQB+447+MsLjrXv49re02j0qeIS
TO6Dv+AfIPPy6wmb2KJTVo1N7KlI0CDksOUcoczPE3ZzSeHDfns3vGUuVu+UOCJ3
Iyt8fveHS1NWu6baEwtwf7BfvHUZVvAzIhqYK7PFPeP0m1zRfgYCgHJFXpe/ZvjJ
J+uhKr931TqYzSQDI01NiUF4+zplSLLWeXc3ADUmbnOu8FSjMx9Rk7eYtyAspEV4
WCrsPCKSyfOw4A1royp2xViZ76AIOyj9smhsEyT+gytdiGLE7SRJjwW1wyeMoc4j
e9wf4NbJmKcIhyg3isWeX02zdw9jmhDitZ+aHNzDNpRwwrKo0qvNAfmsQIKBj6NZ
qpHaLkdsfZ5Cn0y6xMGG+Y5bBDcJJyGKS75lGG6M0GlbG55413gPCIFcrWZvnpAC
F4tl6DwmI7iMKJtXDpK7uA5o+1MmEKb8UGUCdbFBUU6gzqIuYi/a6+SKiutyZsEi
DC8oshGYHOexKk4o6okuN/MLosI9iG9LS/ZasxjMN1qc9TU+ynhLbTPwsLf7yuAW
tULvIlWs2Yd5Tw4qgcRs1w/1ogewcHt2rNdXLIa9sLNAQuijmsBiHI1ySF0xbwXy
E2XOzJQhIK0SSMK+KXBosUdfTHMMiqr7uvQwZF/nNvjQ/mE5U/5gElT7teGx59U1
yr5YbgFXQCh+ba5bpadoVWw0dgdrKHCs0/iGvvELh/8i/wiPGHU9eVK9b9Bg/L5y
uGQ7AFcosbSv/PkZn32cFu/st9hKTxKjLYV3rgGMRoqbFaQDzvgr2JN7XsW/8UMR
zJeHz/HA839j+PWxiuc468w4E1XJZu1/yE1pthF7m1tnZ92Tj36n0KWOSsCZuL4Y
a5flolSAbRgFkJMIv/s3KBvLq9Xw3UvAppXLgDIWiXPJ/ZTKoemdYI719Boo8S7a
6QqDZWvc9chbuknCkmJHjeqybbmgfPWBRjbqcSmMiUI38YT6Ahn5oKZyB+qut3aT
9RNqHvTnOzUdlNpsSj5v1E2+uF6uuxYb+rYI5y+QFpGP6qVWKkUwpUVJcXK7cdck
G5EEPemhJt8DbPwIXvk3OV4/diZfC+KvGAhmInAfv2YToIuQFSz2vJpz2XMSKsPK
AlDhRT9tcXj4UA4uTRoK7JljBH71+QuLyJ99uU9XEzmj1eYPpsedEL5BY+jDMnlD
kmt//PlFjQ/e1Hx3l4pUbMhciGQrQAziUzJjIMHrzGQxEDAHQjWFkjqHMwLJ+F+O
7HD9EUjpfcnOIrkWtHDZLkBKwywhLvKwxvUIfXp3a2d0mF/4nFCRCL6odqWzgHzD
Iz+pY8hl+XIm78uX31oQOxuCu3s+Nu5YBHW/oTdxmvonVzi1m9Vx+jl3BtXeP9wJ
IsTLoJmMzRek5UiOncm5VIb5NppnB2eRXc6zHHr5Rs4BZnJkKqxNVc5v59Ay5lGm
RzPyuflzie7CIe8YLPS8WMoy04uon0FMvTYYpuVx+/o+tLLpTEtiPY0ncPzyu83A
NE3oBmGWX1Nq1LjB/0Bol70pqM9mj7asvDvNLisifCCluWDmJqtZWwOQaZeg3fYH
+JOgjtDCVXARqv6vpS+Or9r3V4qtdKURaInvEZmIkjTEAR6O8h3bAQjiYIrc1Loo
Y6kTsNQu49ZISu4vfNGKNes0OHd/9aigkUlPMHd6dyAZ8fwym5TLSVVQi6X4U/2s
otmxoNmRF1j0l/MkAmv47ujeAzP2AHK8kSFSiGWfyiCzzleoEOIdFqsZTOm7c0hT
B8HpM7iOXpE0qOx1su9hSFj+Z5oq1u9alEzBU3w50AMavgdmOgzHGAdZibcicqWI
+EfL9mwVj4HTOBJZs3HqmaBbnCPZtsSpMFY5cIUX1rrJOMC8sUv/Ff9CQOlOUcJb
jXRif5FdvAbLbX6DyV0Nb2gVZJYSH4sg0fiHZxNUsITgul5/4W86CrDBye3XSPoW
Z/YUibd6DGYn5aooVChJi2MOfr+NlandQDT879SN4TlvXM1WV200h+1HvbPFhYcu
znN0OqxlxC/euqYjKNCtbelfpAY31k0AdQ6ZcnRvT/ARURg+ZFWzE34NHL37vmCz
zfGCgDEDJm3JyerglLh1dtaKmEBOqQD/WrwxFDcP/GyBshk7gzM+4pld0wMM7rYX
2dvWyFgBHRLIMH4ZdXAEX9cGR1LX6ED1Fs1GJl3TTSPyH3uiA3Zve+JG0u38CbHO
Pg8c9l/5rTuFfGiylruzNqd52v+QrENUpt0Jr8OXOodxmPX4Rtyu88jtM5VpLk97
YFJm/NGQgj/kANKEc08GegQ92tB5Z3QU/df1aSPFthtZAPQSd4nxDXorNsUTzuD4
k1onLHI4PGwMnW5eQrnbAw0YuEEMggscuGbzDDGePEqw7OssCWKUPF45sa9MKada
+58o8CPqq4eDIuBJh/R4MDT/UiN70K1rNHlfglCohLJVttbivFVkGj/moiAdxbky
e5bFhnHoW9zdUytT51brJhJsyk2P7drZvX65yDNpCI5xA1i/F3nexBMaZ5tpdDk/
oz+BTwwx3z/5Fm+d31CkzVm2lBnhbyO4qasJDeVSu6rCT1P06Tb2DTcAwuL/8z//
h7j7A04fjjOAnL1nUX0JjlfS/X1iTjFgJiscGZISkp0Gohr7nXmleuXrHJOFuZ8b
GvJYgEaMKHHM8eNCQaasSSoC1JwOCTaAmgmUz5wXJYZY58OgYVwnhgn5C3gKEQP9
Sk/VtWLqQ6SoMyjhvuE9DGjB+mF4uiLHjnzjR8Fo+dkvhoUl8dKYIkIp/xEiNRCX
OYtW3dXiSEqpxLfKCZWMAqHF+diYJCNrUozDc3UsEvPH+H+y3xcqyMkuL9pMrFVU
xW2tQbu8qCY8AizDpORqc0a9QA6IhqUtP3TrgmAHzxjwywM9qvn87jv1Df8mJKu9
Sw3NxNR2piBwcNgHc42qUQohI/j6bVU/yga9qn77oNoITAku2gR9H9BAm00rZsUV
acCLj2TyNOB72bMCqYkliTXYydRvWlmzs86Nkgf21FYX0pE+lIahAsP2CNcPH7wU
B3q1AQyBd6l6j+lCizWblq0wAgHmErj6zJuSzI3sMODwXeS0aCdCx5UexfhZnLJC
fSK6MKu34IW4ggYRoYBF+hEsGhGdgVmK6p8I+fzmpV20YS4ft+gE9PM+K1DFqDOb
WyjuqViu+5278B9Jj/fdFL9luJ3z5PVtMrNNHvuWY0u27tCnlRQfQ00jXESxO095
MR5+LDbtgAOiSokQzFNiagTqCCrUz0b9X2ugKNPCVR2hT1Jqu3mAyHgGVAYwFrEH
YuCqQEgJCBncZ1tKi1IfThJLtR1ZRlLkvOFG4ftwYL+cg2q+HS8fUCJPK/hvrvXF
JayRGKd5T1HR1IXN2/MNGdngi9Yv1qbcWuCxGa1g3LoJRMg5eTtPOh6Kh456ApIc
h/np6iFYu10yYJOxCRKTONLzFtayAVSZ0pzvAfldG2HHnd6yOoOgYwoC0pAWPy2j
O5eWp7eIL5RxmLIagJx0bWRTiR4p1vMYT5/Dc3eUpMjsRENF4GDoe3AjDmXav+/t
AbOXmKd1Dveubcc1Ggtx77FFqzVQp4ziYX/mz/83dMGNBphVAEy4u+Mo0KoG91CZ
DCp+cTfoTOSxaJ8k18JTZUBRTyXlTESWghMzQkxISv50wopGkis106qGbt6D/m09
lGV1A3Up89C936eS4asE9dVtNpZb4A2o0WgwZKZO6F7xg4Jbrkv+A8Ba1JbJOF6w
AfQaTEUBt4g4hxXBtXn0GLmPxnDc1+PWkYTx6KnYxFhOCAGCpSDoAizK0NmHIHGT
1vl2+UJifHVpAq4OofbDL+qkO3Tn4JHqmcitRWc/rOZK3G3qbsWphZ5cDQZPsvFx
kJWa9VPab+qVAClO0Gmcdw0NG+xJJqUe2jFVycnHQkckGKr+jHJFxrhjzoCvLiZL
85nrUZFQZZp+NoISZGdZd0pQ0UYekPpSwnf0huRbuF+vLcuh8HnOOjfUIs9FwHoP
bR3y8R6qTXjacNX0/ihtmmng6dFZGBpiBnCO0KvedhnU2wxRwqMDZkzU7jxbZ5kF
hbgc2Sv6iwgLegao0tR4UYlmDqu3cbQzKD4dYL0elhyfo7d6/bZXCbddx1/L8NKu
7xJQUcmiB25OLwFXXMxns+zq+8m+8MgWUtHrIDPa2wBjUZhq+dIKwLPISggrlmsP
KtuL327P/vjDc+aH/Png5Km0/Nryw00Bzu5qKTnxNFeqAL7FJkTYGdsOlQqdOgST
rOJ6ftkSSsUgzr0H43c8LqQzU9KssOjfH3OwFR1pFjg3/1DZM59NQgcn/nUAkjV4
ZwYhwQ8r4qHRL5G+Xn21fQEyNZqkZ79H473QpkjXnh//lWvnl+tehOxRSZgVma1o
WmWDhhLHe7noszc4GC3iOTgjKJASDmE777+0s5UfA3rWH+ylfJ/bYmCF0fEIwS3E
CuSjg7tVFqZY9FSDApGITj9YeLVV5z3uhjNBzektGTHoftDG2vhv6OCEe5lg1VTJ
MpAsQEzV9vM1g8ywuxz84bTgn/zgikeWd8PggwbgLGRJQdqlcBdZVL1zxCJPvuNc
1rT3oemrnKv94uTjDVSjmvv+Bci+tAftKYUa+JFHANaz+4tsXXut3ZZ9bU9sLNBY
vaxYpqbdtgXQATrLPF7rPoAmupclPT3cf0N4w9I3oJ2HJ6lQetUcj1/LguSBX/V6
udg/vRYQi2AlCdoPW6kPryCOnAUDfDNAgdJSf9ywlYAUtxb2rl10Hg8aeddDjgCz
oRyI/KKhF9Udva2ZL3GkCvNxxTZkxRBIbalWH9ZLVCfi1r1sj7xsnc3tnTauH0hr
d2J3uvEhnCtVDDhMZi4XNbOtd+wo72fCM9kMHXFw4lBVE3dCb9CZAXs9NpTMM/BO
Ged0fke/icdX+6RTAECtRgzXhbbwVMVwQOm2OFad9mRsdLyPIMMFnwzyhmtGIbXE
rs+cvBy5r4dKK5oZiF89MxQCcq/CFFZD78Q9F88v7PHkMYP+/tWq3xE6xoWf09HJ
VbeY7i7gLdUAeBw1iTgCcgsvdiHdrLM4IlSxoTRhV+JHfbgwG0WWD9nBNSDC2J1k
WOFO59dvUypg9YIsLp5BwQnmy7ITTz8LIIx1j69iJ7HIRI1whk1Y+5X/T59EB5ep
jhflC4VNOLciPIHlBWVDXxexRzsBmjYk3wBNfBIM3cl36vQcytAJiZhdqQrQ/q6q
hobqE28T2CPhTTmVeDRlQFxS1PrcKdGlmhRE/g7W8O2AYv/6gLoW/SNuent99NSA
VRqLn+28GNKTxXftBA1o1ywb7d/mvV7ZU8wqCXkw4FH65GqlAHgo7ssJNfl70IkR
s6Vl1u65ncYDB7DKj8XrL6XDLX5ydN4ZeGQK6GKq57dNWWznQdvzCSrtonQRld9N
F7pswcgVtWlfo/VZxFr15XaBRm/If6N51aWy2Kvy5tG+FaE0HhMA5K/VSSy2QKwO
G9dbwUSdLHk/0+4VbIVk2qF73J+1HyW//CPahNBZq7Z7h1xMz4HgdyAWBZBH9821
DPfsxtneU+pesl59T2Z4WHLq9T0C+LIkGP3TX011LgDnkfi03qdky9CvF6HNNWn5
YcbNF3m32hYIz9imOHEE32M1mh/qF2Oz+WstHYNqygU9psuNSl/R6smpWrrlxFcy
Ld/l+NqAzEpfnn8ohFR67UEybjYCzTvD7+DNUqsrn0cJHpM3ZECxHX54uMP57jsw
CpPiZns91mSFkZkyDQurUZxmbKJh+z8AwgmCtvlPDGBII2hc+RwtdpKVFbbkp6kw
CnHVkyrRVQ8H4vBNTC0a5xoXdya308rJi96mmlgU1p5XgIDVGbyQUeBZGpsPJ8wU
0H8aC9HHUdrdeW2TSjoDd1SSTnlxa7a3y6vb0ZxfJmHaUm5d13/CTRWYCDhQxMOP
tmHr5oQ9mW/zEhMJZFo6A/Md2C83iqP6LZyD92DS8uBHjF24HtWRgNfD37dpJCCw
I2n9ZVTmqjtE+ySwb80xOF4tQl+HMgrCx1DbdEaFmnpyKe7hdU+xSDkjwuTK70n6
arj9aCJWMDpJ7utG+Szb5qJx4oChJBSyKblANcvb7yYRs4819yPyUozIa/N2IULR
KIdLY+WgWHzLUuTt0DoxqAqdpNfyCkZz35wc3VCvhCcXkGFoHXZikdPrYlJtav0R
cjH2CH44OZ6TNEpgOy5ydNnpIXhxnZDi1GoGHkR7/zqTL/wQVYou3kwR5QVtSOWr
wFJtHX3bd19FYIgtlED8y5BH8henA9R8W/b620TUFZDYrt3E5OuyzkXqoy2bE31P
s/gHUocf5VyRDSsgh0wB78tcg6b3+BPn7rhWJNS3XmcEav9tYwyViuQQj2Hn4uDy
UkV9lufW7aBF1r3l01OfocguF9OIJ7PoOU1NsofO3gMz+q3Tf3yt4t5zDkTMvDM+
mY/AcsiGdEiTVQtoXeEN2qiL0V3EUQyb88DLCs7YGM+aH+fAUUXLLKeSMs3r8TbE
+/diU7p0APweIj29qwIoRwpQwzXVo96ATCcBU2i3otfC4e91bZ0+tS2KRjfmp907
FOXj3gD0ztZrow2f/qSgsv2dUepIHYACKG7oZv8xLKdtGj5o6Mia8MaLe5rfZ4bx
ZqVDWTIAtwOHIX4ax5GGXK7COexcCc16cT6+1Io+J8rsW3t7xxCCh3AvV7tur1Wb
LndeZzwQmnK3N7xuSeMPgqKun2QaP1uhk9kk/C1jhpQEoBjWNEI3sW71kQZQlYhe
SghpAGnFt1kbeLgpW6h4KwyT3//4O1tk1jkQMGXBs0HMasJiDlTRc7PC7mpBerPB
YqsXZhoRLpGmcZLmYbxc9lJyaIsmn9osKQZiW6000GhWzWayBULP1hRxmee1c7Zb
SvQXo0OjCDcMU1moeBuiaUsuRg1LzoPZTRPbXAbZT0D79+FzboT2zltEG4Ti/bso
CoJcVEwuUgZNY4o/jpQk9DGAinal0q4Z9TMyQ4b/kaUY6/07k3WA2U9l8CYny928
2jQgszvpXhC8kg9Xd5d+adqlgsgQ2LyjefiF7VcVdaaGj3WjHyinALsuFIbfRnYF
4CkcWmaSyJTW9PgoSIYoeHMhJWNAbIIjMmaigWFK4GcARQVj5L4yUww7TviTopDX
I3EQKmoCJ3SPDW3m/eMPMD6CS0/v//TachlOfscr2kDgDnRPNfobkUnNRIH8htP6
9pF/fKv1PunwVbH1bSkT5Mqo4SAtdouEeF6P7PUZTVRpw+Ry+vCxQs6Y0gOp1g+l
BMvUCfDh4se5LpCSqpkX4MCirO3wyvHFYANSrigoL9LJumI+ExklYI2R8RpR30A1
gJTKZrkl85TcsYmzSmO9fY8oPSPfuMSGZKxFHy0LMHNpjBstIp0mbVmkq8vhDwSP
YwatBQJPW7DQB4giE4kRig==
`protect END_PROTECTED
