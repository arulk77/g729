`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAnxBYM/0vK54vl6K49Jx+U1jCmc6hmVFLwZLkwSnxEz
+xcH/5FfT91UtZzOo6PG0xIkwn3Fwa7S+fbFvgkkHa7U5T+weQP1I+CXbVo0hJCw
IzMyYxjhR0AlRkkQYQjlJPhEgCc1GY1OyiW+5OUPR7oAwBIbRZuKId7Tr3i8H3Wt
o5o2V7D+hlTNi17SgV6z2naTH6NPUuLdOvtNT4uoxWefmSWEluPTSPJWpYklvqwm
pH8QzAIUzXQIDh5eueueao/YYKMNvlSMa2ddtjG5gnPu5DsU+m3xBfXHBy6GwiGn
ZYY15Q6i2s0wh12pJIaLyaRReVjJG5VS5RBkgYn2h8w5s/1DdEE8NnsMAxhWa4w7
d+pzJUfHO5zPZ1P583+XkBIS5et6pbw7eVCi0wJBfnCS//75iv8UjQ9MizNC6/oU
4KeXEEy67WeB5Yq5d/6gtoy8leMGo3fiOhsrg2qxO5v5qKp3yHLl1zh+/PsmYPTk
ZW4fODiUyqEkHdRoSb60w7HB8sQP11UdnHTZEJKHYLTuM3xsFvYzKmndBefy/fpn
6rJgr7J+KMZOTkRoX6gn2A==
`protect END_PROTECTED
