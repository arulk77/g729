`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIDpCOMfp4fOn+Yw7MZCAImHNH+74Bc637vfTXPiu4/f
0s5NwVXZeq4M4filwNCCzdBhwGRBT03UVK1lwvaKanpmBw2dV9kykb7+YMMxs1Vz
3JMZugM5oueiukzc6+ziVpr/BVCRHeBykHxG9q4Fsx0HZp4DbSYx21Myp9px4MI1
`protect END_PROTECTED
