`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
wax4SIC5ha/+GQgAw2x6R17iJTYZoS4rAxF9VReWpDcqstAKor8j6Qjd5qKaB92q
50O4oBeyLFDQ0Aw37igiFiH9iueY/ALHC0A93wBxhvfs9e4eR7P8IuxfX+AOFFcW
QzclcK8Gh4ten6uTBRlIb7nZ8tZuEt7p2FtGx1PfTqCzFVyRqCjwdAVp9v5M++O1
LC+SsbFsdo90iVjSWHprZSv5ire9+SYzHrwClhdQQgLEnxVQvIyErcYtB19D5ux/
RnOfTMV4KZIYaxEhFEKQnIjl+8lO8VO/l8F/dvkyj2mfupUfPWhQPgYqvJuWEl4h
79pNhVdSnPRQnLYgNosGy7Zi6GQiKUdX5TOGpCS5JtAeYwwSNzAZ6mgFmhcNlcvA
2UinLvs6dUHtfHUFrLuSI1yRa75qfK5TwO6CywFKokAnfgy/uzZKImPLDSrGjmwW
WuJT9p+Cn9IDqS7JEgduWBc7bGPiNMIaRCtuhFgHnLKg3QpFuEn/RHwHkPVyzL6S
JG8Iy/Ci7LEm3GMaC4G3vLEDuks66OOjyaTkHPI6nXTduqWCV9JIP1APcsl8krfM
PK5RxwAGxRh9s6/rtfywdErc3Ci8f/4mCsgqweNJ0U5Tvui5Jri/e+XPZ48Hntea
/U7x38/IQaYAcHk0qpQO5dVVtcw5tMLYdfgRxAYraQCjFWDVtavKYL6L+nM/uhnO
FZLvg2uNOsPAUF7iI1HAZpUCcCryCGCye+SAF751D4ls93EA1LRcCOsr8Bm1541W
9x8OcjtBBGLpfFWFkZtSjqYtb4iyrAVIkZbq1S/JSradRjLATnd33Y5vwX1C3dk/
QUFKxUcuc/CxDiQC1ooePfZqn04qwx0575NtGoK3i9IJNKphEsJSW4++jDqkDK/m
kQQNuik0sn+3vvDpWEdCInntC5hX1N/ntlTDiN4K4pxakWTs1+yJbcwrF1IPpjln
/rDpiFckMY/uw+evp7czEh1ufYnxjGh5FWQ8heRfGizqxR0yJN208wqFXNU+mZ11
qdVKeX4iYNt5d5aDLCwURUPJjv+nJ8H+xcK4GE9tcW8DiAH/UNUpZlgCdFL7f30a
io6G68IQqDgmbOP2SS6a8p/u/dX87d9rF1QDG2Y5R5QuPIeVX/ItQ3tOZSfeB+3R
PQVapKzhINykX7p8uZHbu6YzYVPrJzucswj02larqlRgem27h2vMGfxWrVttx0Ck
eT0lj0uuduDljdoBE1Zb6kRWi6mSy/tcBG6MgNPd0lzXA/WCGfLQqqoSZG4ALx1i
od6hfKs14fuszzbXCRrYnA==
`protect END_PROTECTED
