`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM/xvEL6XDp3FlJhs1Wn4NCrkF37GUHY6RhLsZP7mYGI
Y+yTDJivffMJnqC2VP1wgHB6MZ24jQmbI5yU7PEoB/ZXGXQAIE317A89kDrFIuay
VaTwYmuhcOSyqSZu87imin/yHotRtSWyuYU3nccX2xjxa/O6Oc5qowKDrPGnO2Hs
XYB24uvz8ufLBDJT/7Y65OvuhUsG+crmciE39bnsExFel1cmSPyFTHJqi1VnFGVH
v/B/gJ2/xPKLineEcO3XC61/rw/HYJEbwCkaf7sH7FbCtdLJYOvKHFyv8eFnBqi0
52+mBFNjPF1MwyKF74o83/KsRcrvapXy822b77hKwsN97+fxb5NPQqoGRjjwuYUD
V+SWoXu2fuHSkcd1oDt7cPYFklskoagpXgdzQVY5LSFJL6lDISDB11oA+BfGAtBj
iElXR3jqnPOvksEOTK8FQ4TQ7UFaQD3WV+TZx7o3wJqSDNTmlkaOq3nDU6OmCeQW
Fvrvu1XXVoX7StcWWchrFY+siC+IfNsUjOXKBX/bYcHFSmefEUm1O5/dWS3JRSZh
iCrFvtVvd0SvW4TS2f+4zZOw1t0TTel3Km3y02G1XrbcYAD0ahCA+lICJGtXYFP/
0/9A8pZbUNfok/gbrZmcnLVerA55zv2OFQ5nM6b725T0bIYLuXRL82JZIduoJn0v
4XL9UaJ5nlrLtQClc/DpPmFM/L9HUoO7pWsj4oxQjyIutVVygp/tDuuxBYZA4Nat
37PikxychnCMWqhbwTJ+ecAO1TQa/CLkEGQesM6BpPyFslHZ0p6UU5BYt0F238sF
Ut6PupMm11LMORg6Ziw11n93hO5WawgNYsdxTR4Eh+I=
`protect END_PROTECTED
