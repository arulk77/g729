`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
uZhRrW51y6iHgxRkDpLZ49tkw8XAMeaKnDhVQ8JC6V1v4NqE/0a12+75AmJ4k/FZ
al4409Le5DJov6/5j8VAJoXQoOH0ALfSMerv8nsgoZ+bqvM+KKZr0u8qVcGROb+u
RRi9EemldN5zU2WDj+BHmOW+E1ctxzvjm4TJT6xaGvmE3B42MORzc/PWUEXEsI8F
GxiNk4MMoBJBgEghr8P+tmdk9HTaOgdN7YU7O1KmDNQ=
`protect END_PROTECTED
