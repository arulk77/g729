`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCjznYs/wDnZ/FQPe6Q1qjo1xy44P6TJtJDIQGxi1LY3
Q7jmMINVpOFDvU6X1NMUOuHMPC62n46ZjOGUCKwuKY89ss0pXsKQ6H8x0+KJp3Uw
AqcSM0gJea1upf4BwkMv1Zbra7Z+HmKrVjhaMlw2yih5ZAu48e7WbZ9nvPi0bX3F
a8/pII+JHHfsvJj26+8P/Fb//L37V6ZXMdJRPaf+Tj6KVfMgtrSJV/blzHt7KKrR
y7UGPgd3TN+3AmNs85mXjGyplx0St5hHnLBPNQtHHfsuXcVmcLVesHNAD/a9qmT/
9whcfmVSFtyabpqG39GhHg==
`protect END_PROTECTED
