`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJfGt8Yp8ArqEY29UUDGDm3ZN2H3d8OHRMYRUw1Ew+y+
1qPWxTGD2M+OQ2ntBAb/GCh3dntrZrNS17iItaWWW+VnT3TDp8GntXcympVk7uSZ
EamRaxuZRfnvo1U5NJIr9fuqFhGA4eWsuu3V5pH9oVYomWqL+qvrG3NedX+DaUPS
czKQbgqGhqYV1qkmS5Wjt2TEzoiopAltnOx9fwMEu8ZZHzOvMqX0JObELilmRMld
+RDeRS4roIhMNaMlog4u0Lg9DgBZnExVxxVD7Ri6H5F5J6ZtWMY/cS/aDow8GwOR
2gLOxGrr83GuHWai6fx9EOdWL/ZCx5hcwDRqVc6IhnsZuZQHXoGfKda+pz2N5KxG
CflIgowhPJDyMVoDWJELj0WfJgqm/PahTtktXgK2TAkpap0TRHWJAyJCHkNtYsxc
D2uRcB4BEauQR5zw/ulC3JvlYWTrklPzVqXBW40vCL3Qd4e5+PT8ZOhPBkdGTabI
`protect END_PROTECTED
