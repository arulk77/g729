`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEsZK2u3qbc6ih4SLEQD3FAsIjiPRhcaKGZ2FC2HyCxl
mBn7RTuzD7lDYxPtP7SP7GWTm2E/WoO6pAtpW0lDjnppDOaSRXclVrmU83ZLaQE9
iowcX6V18lmNQCrAv1izCFbScBwN4rBRZppQ1l862OE6gGgW1gPzGDEA5rpdfBNA
W/J9FKJoa4kCitW79rMEvQY6RxOKw73lYhferCLKE/lZMXM5hfabn5sP5shaEjTy
+fNnf2bjFNESYCRgiQqgeJkz41Xr2do325f9otR6iWR9RvgUnbWBbkjLM5iwzalZ
f1byK0M4e3q07Fk8HwfoUHYSPAqJ4wiLC51jns8KN+wcRTEp9czcX5Uk/OQnqMV4
McCtpuZQVFVgKKcByc4m7PAF25K5bCpzgFYLOph1JG6lPJDQPjnECJcN5CLL5Y7N
6MlDsViOTZb+brsmEr8Udeg8Uv0Uj8R+qYiNVokJRDswbWeXAxAS5YjWThiSfPqH
2G0ONZsJ6UlqFgOshsMOITzAzgbjNcN/u8N3nPlqXrTsEYIyleHlAtYhEUyI6l1C
`protect END_PROTECTED
