`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG+pXP8gYfufOzM1hmsWNvtm1U1X/urCyUjObWib4dvR
w1QnT6fjP9GACv+DL5HLAIGlePtbyV+ugS764DTS+M+nZx+8/dD0NxEaGExReHpw
wJG8T7JxZuxLFwOM9YyW+Nctu4/y34G/FJgJDs5Vgg18vSPyf4YuLW94Z/fSNdjm
WrCfkX3W7gTmMl9OZj2OHdXTCNzD4j/hkUhr0tdKVLvnt7RdbtIpvpS2qvUYZGwH
O5CD0+Uw9txCbWtuemBCgIEaoYW81LUaRzYl3XjRcryQ+31nbScTkQ4PoGSeaU1B
yTEdZly3AUbTgb4z/CaI9quwMk4xRyLWWzJg/6RLC1esX4OthM6Y3gYcKgwl9/AT
VxDWw9u52qQj8PSxDv3WJdmHL6ys+/kwp/mqS+2yVd7YOhc4EMdVfiVw7RmtFR2K
TZtDDlWkTS1C4lhPXZwoJ0pgsiIn8zzhc3evL63NbQ8xaRStbzrB6vw5NM2fqz2W
8mDl+FhfFHn0jZClfWfVvLIvAs5yVX1O8dsSPKd2vpegIOvSMhM9zVIMcErDJ4vq
4zw7WhTVuAa8ylQSThM1PflCoDlIIGnk9jWpBib3SDe0LzCyFXp3uR5FCRoYJ+/v
y3ulRR7IxqaIYNYLokcjLrPgKybRB2zVNiL9ujh+iJY13GplhcpC6WVYCmf4ERIu
V5a5sRh3aUDLUfa5zytBQkH12t4SvIssJUX9WZvu3mWtgRYfMZ0C2/UNTFSF1pnF
b7S2+pdiKYy/oJ8bh2b9Fck84yexwlh/fB8FsM6JbKcYewaHmJkQHl6zK3uJE88l
YF7RMWrcCg/ekVveIXauuZ6zhGQZLmmcla7Uq0OFbs8Ljc2uyHvREw1AOxwdokxZ
/L9/Kof3sGf60g0S3vWoph5liqzDAba14mH+fshLr1qw0gs5oV0xngE5577jtcIG
ULmzFk6FNrl64ssQtBtds9luG5oN4094cXu/uL5HifvuIOynK86U/TDci0mr4dkD
KnJnygPCCGABFhzcL4PUR14RepH/SxUjAhrDSDvMrufYqoBynwWEHhr20UtrwWbw
qdTmyfMd7mSVIBEZ40Nr2EN4cHHP7r3M0lz+c0BajZX3cSQLyQ7Wcr2HVtoVFC6X
OV6pjieX2ZFkjto8JkcNrh2lq17d5uC3DRHyjJ0Dq/g1K+FhuMtAcWmAHfXpMIqo
wlKiiRVcbxbJdUkcIsx7wtYL8EyVou3/CKCdA+2WqjE/JlrGRMN3wb1H0PHYOG0H
/hf+zLKxw9lXEvL9OQaPqeBEUCEN0JktezW8iMKckQ/Tuo49O/L+qeSNCbNJb8VM
2FrWlrVRl24DvcrDAauDhE/Pl0vfvGJB+PjBtETB5pQbBwY7v7GmrgqbRlYx2XT3
SHmggZXkPJd3ABHM+tJOAVsIzRWT0KVSe2kNNWOufk/FJUiY/NXzs3VCdGGGbTxI
Jlp1Pq6W1MxHIWvxAXxwpJ1/2Q4Rn/0qMCZTftZAIUs1DRlQibsJwyDG0He38aWP
FKLCz7cDQFO74m+/SG1Ps2qgF3EE0KILRuiL9RqI7DQtju6xFPHiEpoe7eBrfpTm
f0T8MOojiouvqdewipFG3bD69XHJAsuBEgavk94TKuGB6bzvrgEj8J1lrJr4kQ95
SJg+4VwCaoU6WbvV4zU0JZ3JRG+uL9jxewL3LadCQ+SyggRe1CSefFc800w+abwL
DUdA3TWC3V9ri8+9d4aKu8pX77RaDxRtMtHV1cmeiWYKJ7WILJif8kpt+maR9myg
1GoD4ITl028DMlw5GjCSo9BacLprZscOeIsZNZjw/5g7e1DA04rT6pizEVx+AQcy
r0gMPDdvOGyZrih6hD1Mle4xtxYyOU1b890Ag1QihzjKCl+VIT00v/YolnCVRjxb
mzVtozByE7jNjf1tXAMwMvSpfe18GjukoigUkHDdb9+z9aBY0d43IHk4H0zAjhj7
8DR8aric/L0tn0qGTEUP3WBYKiNYgyiFSq7M+QAWB4L5IZd9JPqXcXTPVIFaheMc
NKv9pgAeu+usrauENh65auzaSYGF6DyrR/YfJd/Gpk9vU6yMzJyQ3g2vh8qRi/Xx
uK85SE5YpvvKnmiN252gp3yoWZqQH+rlS4Fu8idIsvI/Wx9LABZw/d78Bk3Ch9H2
8pjYYcg0AdaalRwWsrGPpOxpwaL4tsis7yrBiILXWBv2YAA5tn8CHUiHpR5CxwOi
LhSKhg2tMzPyfynP+wGK3ZFY0XrUsKflM8yRyO5mLRFiI6UZ0jeF3RZkaAALwex/
FdXKcMYVNpV5v7obM6AyUgpsCHBpMTQlczjmK5TzrrdHO2Dwh6B9MsxDir6s9du1
NZxHNbHmjz3zE9JfWGgHD1cfDqlsTWWvWqrERypgRd3bkeLFOTtNRBf79+8LxIjS
6rT/DItd19MOvzwJjJdd/0Io2qm1tDGpG1YnDWID+VuHJb5yDUgYajO7GHyOfaLQ
7fOW+H+uTYWygVJWWyhLybqFhXM8sNnyHlxxPdDw+OwvcDSmWYh7r79w7VxKYevA
8DERwnxQ3hSAEYjShxelbF6XbbgCLR7jIeavnbAjLmL6lm08Njahcacq3TGFCrdO
TpZjqWfnOcMRcLi41tCTLauYs/4auPGATEF7vrWdRn/z0o0DpT97vZBh4vb1efcb
skWzXzfY0ousWKcsxnEZg+34oZZ30Rq8NMpZnsHzWV5CZnhMdOJk4YEUxOh/YgBM
p1SFxIklBtoU7/QGNlo8hS4ATKz1MfdPmtMmNf8l38MgNGtxXgwFGNBek8hDshmV
pqn7ipMhHu3cYv+6UtBYxHOkP98XPGyaKxm+HoDxpwIwqUa6fnUCqPNXRPPsmrak
UY22Br4dhqsFMojD+PzXBDJHHT9Ryblbws6w5zCSc2i947i4Ebm00W8DNnSAWPDV
6Z9sa4WajFN8Xxy0Tw6cW9oH3b4qRAq6xOvugxBBJORQg2FVpB2p10g2Rs+EMtPm
5GiC9tkSAIgfQm5FBAyfrJwEypoTljEtge+4HzqCdXQ3Y6LrEwvLcr6O/gZhp4Ky
V5dofvO1lgFimu/lxrvNtmRcIidck6EVUAasP32m7E8daECR7/J7DxIsvOKNGuRv
bDojVHuBID71EvGcgtwEEw9IiWMjeFJYwk916BTy9HWiG5OC4zwtgfchs+3s7yHC
yCt/tGcJAhot2YIDy+VOvZmSUipUXP84vI3kHMK/Tskzm7XIEuw04owFuThSX7jG
p6DlIujbPvsDRM+672kLIepxH3fCtfE3JpnpQ5oXOjaNfPnhBrLuNgpH6a2tKSfW
Y2oTSlBTt1FHCLfA872qQ2rFLbqnq8kIerbbilquJoxcAuaB59NaW2f3Hz56Y3iE
t9phHKQQAHALY51QKE3Ixb/ITYNR23CSSva8u+7lk7cZbSPURjkczBElDE/JywHe
4o+KcsB0qfHvXuNBI1dNN0vsLSqWVmignP/iAxGN6z6b/zM4zc0ZlWJfqQe4d3i5
+IEaspObczcAXFbvqgE8MhcRVZvrDjKrF+idYaS8mXjIiygjIiGRfuAeZVlwK84U
htpYJPkdtWgpcPd9uMAXVlWhBO4pM5Zvl7rOUaPJcw27P8dXGRCH8BtJ7tWgdSgl
HSwMjx9nKP8gEPFpw4Qm91WF/9VMQ0hFXRehD2Pj9kS9QSJsVeIouNynylMettKX
MK4XgGSOMsusW8De65/pH2iDk+RdZwPj31w58EDLmd8MUmN4WCYxqcq2WRonPZqF
tc63mJ9oAWsXna74bCMkaccZx6NajV1JNkwyMl+UrfA1qtvB6ThvI6Lwcx3jeX6q
guKVtl38ACu77g7vOTsEFAlsGvjiVcgZ0yh7YLZUiACNn6zCeAE8lAhMAgqH4JB6
DqCfLGf9ToudamiLFUFnHBfprHCVTaxQYgW58abilZQG81m82ILd3+Xl40cj9L31
SZsuxJpGnF2qvBpkIaATtWFMLiwpqsS0BKj3bD56KvHD1WK3OAQNGelZ8QTOwqXh
euAs+MPd6ZhNzbFeSZ3o5kzU7BzyI+mYxbFoHy7x7IAoWnE40IsOXktd3l0V6MJL
xDQzhD/Nu4y5BzB1OCeBskDjSLf2dBv2QsI0yk7BNTNGr2eOrxgyHEGakgPCj61w
niB4R0TRJMtWExS4QnyoYzo3lk/FG7NHGueYM3dNp7C5Ccee7qNB+/XvEImTVKHQ
M19P7NHLZiaUsbATxFZyKFVrZ+2QQ00pUp3JoriDRezZ3NGylEKzCut6rYGSGoTU
mjFmTH2PSX7zXQd2KalrFSXPL2+/0I6BuO0TUnyYbJElf2mYO+Ld1NKs/TvdkQx5
Tvg2VkOnkdaDMK1/26pQBsh8F5Hf2LBHv5WXRdhz4TmzFNh7T5sLHVI9RF72ZElY
8x7EK7RSdPBgiLUK749mlRA6P2pxl8Hort7YZraqcd4+oYvWR4ccyZzrVFM7hSMM
+ehvn4SGspyvBjkvk9WJWdrqXXwpNTgJnVgZ0U6lnbsAB+1orqIId3qpiYWaCgwj
+FAd61642HIKezTa7TWZDh3zRGQXczR7Xaaw6SDCJsjMzuUij05Y6lg2uCiFACHH
EO3TYxR7LuXC8Uv7ZnFQ8uhGIz+rR1bqeExbk8EBkWIQiZQP1UX55cOJ0nPwXXjX
NGL3SNj6kx7sqYflSv8dM6PiD0nN2EPXY6/vuitp6LwvKtO9M2fK7vTU55DbPKC/
EeMeKjCBr0cnzPPBFrXRPslKq2LB7S09mma7CnLKO/FEBh9ePtT0z4F6rdYqcd6R
88ujl1eK3DZK4RyygLRJ3648p3LqZh5djsbTO/fg5w4H8vewHNPptTHEO8GNsHeB
opREDbzm1ThPCj1hZyf6WyqRfHHpTpeHVezxAA+0k+bGUosuTG8uXw6eMQJncv+D
2ctlec05wb4X4zGR5XdFOzSWS/Gz5F1icb93+dudIU5ELwSDVCKbOciWD/81lNIw
Zs8DZcQIK8X4/gTeExs6wUovwPiowcOKdqTxUjgUT44LGIyb/6zB7LZIJH6PtOHH
YYlkA+ny/tt6c4OTfPK+eMyE8G+tu/ccok9WyO0mOHJnAWkcyaPk+6DqCOi8btpr
YAhRpxM1bt4iH5WoXhcokpiN1av5yvz3krtGE4JaiW0nEm6OIIC1LoYxdFZcWxVK
HU3Vo+nHgnK/Y+hq8BZA7JMC6ZjcBms3gDN3mpmKjtUh/SGWWDmOxxkhuZNO/KjG
RWHOz1R6E9cgJgWCVGIEuy4fHggpGykO1svFa8uyFKjRxHbZsZVjxFK5O2EynWQH
Z/XxkyKN83jSGx6dj1/xIMGCfh/ua8uXIBoUwQMqkNeq4QDHoXN6qYPv9hQDS6pT
iSxIM037mBexwirNZBHPDpmyj2SVIOs4ikuESocMDw7vF4mfQqPM3Ts+Eavx622M
21GfmNNxt00JTVN4tpipigBdnQ5n/uUZe+HoNkzsPcVNxXpfFyxZkW+1mTrdN50Q
/OnuGioZm+Kivx4QzfI2nBURCCm3AM+XIaOH1gCzoLE9WqueYvQzvg6lFPZ9n005
T8Z/Fv813qmVBw5tgz2x+gx9hENpdvziMdNr2mq1L/IcAO47AsoAePwwIkOdNHBV
5IUgPqIj2/tJQ8BJ13vRioLmhGKpgdzZ51icSFXg3HkhkSUxRJO6CFt1V/dDahc+
pTSv3YHBGzSkD/11d6+Bf9r+BZjHhCnXIT5xXkJSq9/p8qmRbd5HRicsqDsSXi2X
Fg4IIonV2r+8KV+ZYqGM83ESLl7+NDQ5g5YTpQswk+OG7rjdgukZZ/CV/+XR7lQj
EfVA5ziZdIW9gmDNyF/6SuIe4ka6VExLTYFBdIaO6kSPCopDpOdIevUTcs3/NbhT
Vf0xMCKYkulN9uuIAEPw1GPiIMWEDSMYngPD4539pf9YRH/9CiyEhxRqzsUoJuCs
KmbdXBAkV4aEboQqjEj2eKPgFceVo11WkMc4S5+916mfyvfBymSE2sDCmenfG8Ao
VzYR7X/sYAHw5FaWMwWyyUcMIzpbnJWPlmwpCp0ADtZnDPehwlkAnrXD+j7QQEP4
OihDuLtxAugaDoY3+A37IlQ8XgkUrsJOaTB82XlboeF3LlIlJM8gzEgYQ4Ott3Lm
X/kMaP4bcNu6J5uG7/WYUzkJTMyd4MSdOA8h6G3tP8HvRwH7ekiSc/5v3drB6P2t
PSwjI9QlBgakm7KFyDCTaydxpBLq34zGCbsP1aRrx95m4yFzUmcAccMih0GtpFm0
bnWN7j/8szIFcfJTgy7pwz2RL9MtGamwz2d1C4xPWFPYfJStMBzrRWtgzfBb8MyI
0W+tW1nUztGpXXvhlg4AF3zasKZKYDPKMH6FcVcQ/5FxX7W5EsBkaKnepWS28X+e
CXea94r9e6gOc7vgpMyPpe7VdRqcvr0KLGufGybsy0KGKrBBrQR/lI2aLYNuenMh
5NHX2i5CYlM9jEKnnyn0CV8z4ZEKgv4UUl9QI2H3V6Q+2IcQDdjahw+qhpS0n90F
h8ZdHNzbjA6MD2kkzqJ3/I9Zkd6ira3DM4Fc2V+YldjuoQvgflK8vEk+qnL28SQV
UydR2SukPeDFrhRFihSJlDS3QTNugo5Is7FvvLfjGBFFAOX0yjnlfN/9OF5y5j0A
a+kh6sQJ/AQU2LtP3R8zIrIN1BiLfj+l5/k/UBq2Xz0qLl0iJki0iYuFPmCY4hoq
js9pk29q7PCXYup9h+rhGJBABIlRNNoUSczvTcbrXxMvzdthG+9/7dXxea3O1tFW
zkFc5rcTitdm7/NP5uWjkowWg1JmL1++hwrs/QElbzaDe0we8mO4yrSJ33zDmEgS
S3LLCW3+i+U3agdFHVTwkf9iumGUdy98P2kRnvvFooaB1mwbqFvCKVIpMeesOwuW
2pclvyVpCn01CfZIH14du13HUt/Rdi1Yi1xoTnDpFVBeOlzjgY2V0+JlQeiCHDes
PiUVSxAKlDo7r1yl2eMAkFP6YOu/L4M3hoZgO0dcAFJuk4KNGJXOWweWN0D8O0m3
Mhi+6ZmBTMd0ZzglY6z6L7BGkqMpeV7DIdlKI+SRj9zAtylbH/VKmQh5YsZ7xiqt
aBo4kDhLAifWoMm0r1bOgFmWm2t/83x2n+LpYLeCDX1Z0HEdVS500Ne/9jtI8Jkb
LaW78F6Mv2GWMBk8aJWVgPGtfc9d9Ok2lDtHryy4wHWRgD21lihuu1u5MvSL5J9h
MfJFrlxjsutEaej++fmT6BCeBIyO5SrlX3tFK4TmXxINLcKyjHyaErqgZMD6i4Hb
jYViAtN/XArx2fkR4BM4Ty/XqO8vkGFyzbTWRj5rd2L9o7c32CkWEU5XkUUJarqA
qjO940LlMH+5qmB4fAji88hF4fVpWZP3VC0xBcSItBJ9mlu+tT7zh0XELVCMKjKn
/+JEGQL855UHZMm2VQHdL1epfwcVD0NT/joYtVWKeeMXGtut8qidDVRTayTVmkv3
HlzPTgImVt/R3WXo86NLjH9+EtbeKRLWoMjw8R819HGT/rqeMLAE3lX6RguWE4BK
jc0jwzXP9yvBZgs76XdjWqFqM9lID2tBt5YFt4eDyNjmSmAEGYy5qHWM7HoklVIo
CdI8IBOhGli2RfQdfKoZXJ13x2OQg2UBJ+qBsWk9EffbkfwdF88Qe0/UXdFl1Qr2
UTCQ5Q7nwgkuLfRmaDIDyI6TP56RogkmQOVnNHR93CkUawunrAvbvb9cJ3DW9v8P
wwd+3EVEZA6SyyyQr1WcYy3Z5Eb14qpqy3lQSKFhiNI5CJiWRXmHGaVmg5c5RikV
5mxoDGE/8dGz9Ce5dQCcX0NTusZKW94TCCFQRjf6Asbslg4KC9VPnzR/Y7Kbxu4y
Xd3pl9oU1EWWomAhikpE3Cr8AThqOeQ1Zsu46b7Z87qhd+m+Vcpd1kEGflTzqkc8
lZoXLuFLzHgxDl7APP7skBcAGt0hzYinTGSFQVEXrIiyyx9ZJR7T1YDn6NJ+CL1w
HnNlp7jyXshv6WU4PXuoyxlECwCrLoeos/MANs/EUZiZv83kbhJavi8ILMJxRHrX
OKFAQrz3t8tBEu4/p34ddKj/7E7ZnciG23ucHeQaPnicyQB+J3owQdDCnS5zVx5V
BioPuTKLnw2xTxg51KKNq0nSaRmDmpdjTF1w1if9SSghKeWcq5+eWX2l7134FKPz
g76HB/N5KMoEnos8TFoYODXC3fZCUCYvvK9W4rbcfw93mwMPe0Es3sqfom6MET0P
t2+RSmyWR1yr5cGyd+YhF4VsJwjE3qWllACiZG3AXQH9xFIEoPXMuCWh2Xb/SGiN
7vij23jubJM9m8WjMg/IaVQqLWeycWDUDEVaCfjkzOytnqUe0omF+ESJXakCt4dv
zQbPzeSewQQaJzfNNA9BfZNpNj7ussDdG+sQwX6V4YhyK8m6vgMpOsKDhRDkU9wo
JN9O9kUbR9TvMhxF5DhhKfYDHQVEdJe5LUYk41EIJRUEycjNW3ckLC/TF5vS4ZTC
8194VscVSZ9J4h96fJTxcOo0PsFhmsZ0NeFqVIOlUH/5e70uZKLaBf8K8cB3kAi4
zxKxDQgEKGhWqxAAqv5/G3yQDmpXQUczD8S4MJFZYi4jBuFCMh1vhNIlEaVGCEYr
Lb7BOl9mgwnutDCYbCr4AYqF+gyYnayEQsAkwQhYZfli31ao1hQwZxRrXSh3Jct2
v1BKkXpbp7iBVgjRSRnLksT+XGMZi0wT0I/GoxVhTcPZZlXuZBwksvtAfqQZrL3n
mqrYSDpik4kSKdfn4pdYyeZ6X5/7ATbesaVpvLvHuGrryOMYnOXCtwhROSJTAFoU
Ueq0Hiyoon6iiYR1NkqYR34ipKyaTwqmjKwnhbmMM9GxfwWXBLqR6N8U8Js1eHDm
Jf78ZWa7k8r9evJ2sSPOGIJqL081sfaRf5oUo9vqo1LXXpDduJEyknI9HU7qx7sg
ha4W8mlfBYMKeh3yJzi5aQreKvUnY86esPQb8REclSHaeXif9sQkeH2o4kFbLd04
Wd17IMXRpu/ofnXb1Oj/+DqdsdyIxKCpwY6PW6iJ/v17pf+YyVp32/Zv0jcUkX8P
9wEdi9eyUbydhqsYw2STpG2z0Qjr/YOC7m7Ks1WtIGQlkRmVo7T9LKxDjDa/hC0+
LhGZNW3V6+JZfmPD/kLVH4e38lDak89fGdaTtCr42AnGyUgJnVht4ns969bpXd0y
jH7sHxXEJaUjqY5AvdDyFacF+lv0XRjzMoYbNByOmz0M4gyQR+mA8XO+DcnqeuVl
KMbJ5RlFWkaifqUQLm0fTqdDOZXnK5wO7TzSn+M3K5HFAZ6Vygbuzq8hh3+8oEnM
z8Y69N4JvkrFzP9jcIF365Q/e2jcSbkZB1KAZWsr1MZI5AaqJQe6df97ladgWggn
fHqrmoJC9Ah0VrfcsOOWvFJ1B36Awz17x7CiNXBqvrUsYYTZ0aSchZw5JdpwIRW/
2qrKO//lN/VTi7TMQ30U4cw3N/ppBTWRf/Agr44fyoWY8MoBW/ctz/hnXwjThfMp
emtXjzwcbV5eBJPBlPZ/JrhwvalEbXirIaYEmljyTaXKHP/2ERAldRb3lsVE7HVj
8BxoA3fkqvdqeMRuVJ/M92SSKmVreb39A3X9seA0HSgMWx9mXdFxSQXPYz0aa9gF
zjEerAWsH9zD0OWttCCXbh+1WjTc4lYN+f9LDnLM2PWE/isGIcYFs2hPLbKqLZnn
qHqBQo3H1EoDdG5YaKV9ZxmIY2oRUceO4yqbzGKxX4R9Z5wYA62pBLLP/lWoeWVz
KYXEXmEfu152JR/nacK6dzqa8uqmQ7hf/SP4sR4UNjeP7e9fCh071RiUSNb/JvNB
Q9XrgZT+f5ecKrAkj8+4KHt0omwHJ7Dycpmnx0WxJD63ncTK28XHt/+zGZNRsdGg
wcroDjBvJpvv3WVX2ltcXERXek1wZv852ne0+2TLoXXrsw0O9m9l2aY4dKCbZkIG
YRmNSMuxY5uG0E63i5azboKiWcafQkvincXsSnwImVetZJp9yhKJhJYdxhc1Lg+p
Akg5LN/1mPaFpkYf2dghAveODX1grDBGevQaHYbeDsNdir1WgMWAHI6SyNhIreVw
brfGMgzAXZKkyzMZ8zSDEyRoIlsd+b/+y7qayK/h8pn90kp/ftkld+bTBoa7jl9O
lpX4MW/zAtF0Fy8lmiP7W6A6egLlV1vhaNXbDPW+meLbiC+MVUrsBwIImZW79hfu
SFOnQk+xF7FcUFsJ5qc8nXJBjD4GWLTb6EGC0Y10EPQFmBxEjbmzI5A2cptb9tvy
thd4qqPnwT9fk5VFKXFsyDn3ts9/K5Lsj1xQ9NQ61TQSsREDIJg/rnOIPgLfpj3i
ODU6zVVg2/eCNwMZRQvJnPbUthgGHiUcsg0iUttX+TJCWWwscvvoySXpECRWi040
UHpmCd6ZdYnp6w6qriGKxOjAWr+pAptrWWlSTRaDpUjhLw7vJYEr5GPS84LK7j1t
MXmi52WxB3Ucm6p8kHoFetEcY3GN7i1mZDEkCkUq8O0JnciaIShw7NnL1VMHMjLl
ASBUexnbxByUzL+jkebMvPMgdV6Xk/He7hqK2vahpWpnkfqifwrGSVQRw7Vg/IW2
rVjqC4G9j2paHBJGFKCK3miNCltHWEE2FSRKha/1KPCkxkhy9oDQOvtvTRK9eUji
EhP/EqJJTExlyz560UhOhnPBORUgJ3+oaBJSR42OszOC71RMwbItO4xy2CNHSk4Q
J7l5OqFJz8RT+ydV7pL30zd5iXiNqQBHpUCIpEnKysthjzn3lqNSo949cMQ4oQzH
CZJNFb5vleIyKoweH3fFZXq+AaAfy/Qn1dvsYBs+Lh5KFaE5oZx0E8MH/He9zEDb
kKeQLVvw8K6aX6r8horfaj+T4trTr6mIX0PA1fxHpZZL9l2Pao0lYeZxiQ/zCL14
Qtv32RmiFY1UbdIIVCtgoAfpJksqaruRFuyAKWniZo57gLHLzkdvDo7m98an7V/3
lBOj23X/HEMZsJWyOnLxT5q6sGZwA2u4KkOoJ2nlB+5zXOFyYkEJUsEOjgmQIDxe
3jIHmAIQq65yZNE6azqfbj9fADqgBJu9/H/9YrOFbV/FvwvCARWONjRdQFTr/uMy
4Y/ybRJGRHTMrZKBABrNmixoIz6BRFhmTGXGh+so2mV9pG5xHnsLWHxsrrP15q7f
E7Mt/saIPgJY5MiI1HtTdmjdsmXBe5kSYuy5rD2eIJAXYy8NO6oBn/k09VeUjbXG
C9Rp1aoM3KuxI1/dEbGOeXdkrc1qq3vxN8TV2tkryE06bVKStUeLNnqJ6tvjiFhF
9B8Q4eLBnpy/MjgG3DTPa+2kBJZvAZaEX4DBM2I+OHldbGycsQb7vSLSSijiv2P5
rI3dy0f70xiEzCznioFamWgNv7tDtxgpB66ikPTJFzCx4uI9/QlJNliFR/2fCyQ9
9R3pjf3mye/ylQfw+W9WQl58E2ryCzF63cSgvuHD+eTV6ammVn3nrz7dqqVjdNHb
iHYV3rf4SWY1keL+bowj61YpNvj1fDrGx5+rupYtr1nhME3ViFe3DDTh3mYGA6RI
NgxL3dTawaYZ2wfYhgVXJsC+iMs06P1iFVKRUrDeXLKoLnr4cGoyNzUBbvmCK6mt
gvv54d11NQ8aRKO54yILc5e4VJem9H8aeUmBdkxiu8DiOdPYiw5Ozc3jrl/u/s9E
9deJuph/ZSUkS7sLfBW4G7JaZF75+p5AQUHubcYDoh/PkSrWjAZ1cp87XOEHEGER
5DLIDj+FiegpdwcLfKX81Kzpz8qUK1irUp7UT0zoEJ3+ZpKrV+UUHQKDG5z7AW3a
UY/gj1hKf10OP6crSRlhlpy6JQAdMPA1T4Lzy+bmwWr77PlzZAgd5qTGtBH3uiyB
Ym2zEVS5NSZWw8J8lkKBKXnGfGEtZgMWJ/KjZH9gQOg1fx2dsNY6Zs9y2A9Y0Tsm
ytROC9+VpQR3ucKX0/MFTtvXXiRT2Ww0U7X6+pt4Ug4IhMPTESPPMC9vRB51Uf1p
79bdgvOEFlEu020A78GU2ooEGQZHN0oEHVPg2uTK0M7scU8VDYHNIQaMk/uMJnZ7
X/pQZCV+9ywHJyf6YWyinuKkPz7lfEUS8HG9Bjn4dgcaaAlR9uuXq6/i1K+uI9/r
px/ApCGoux3LVQ1o1x+ddCc1r+s1ANBAJ4VI4dStakPKD3Uv+3EUm3dqjn6WB3MP
FUQjuNv6gjBcOM4XrSuCtv+XQus+UuvjrBdXG0XtezOIybHOONkXl6i1VBomk+v4
bH4vQ/mPZxXJudw3+AkncbxKbGkbBOa/KPUEh8X8kBdTXeTqtneNJIWCogFuVwBg
PDnpDGER+TwBGx21ShQtydctmHbXzOIXnKcmyjIWvBTVTpQAozcKHrCmi9Bax+T6
+2Ynk/M/1A+JQHV2RTWSDJAZAPWYTMSKJEL9ejGQJQ1xjdvS9yBGxqT3KDrZjtLp
N+gO1v8wtUWZ9w9N24LXf/EPTH6QiDUm2XpJ9fnfWUbJ2hxIZJSeSrvgkA3z1Ggg
/vvL4q5M39L1x1Gqeh9p/o9nFyONUYs306IsT9+FltTcTjfm3HL0OuzlILsB8lsq
tAzxKBmKr7jcJEq2S4SjauJCG27029rxnZ3hOZQfcVsCaXwhq783BZYZYZhDJKnu
zRyTzi+7y6+eq5WYiKpHVZHkVTCuJHkg7GoPQSnlAJYRlpefIq6d/6OT6vlG9EOz
B3iczLTAG6qnkLM4hMo/jT1YU1315I9llpKqITn7H5033jcl4eAXiuH6gO0+8ndY
jNdfySkcwVCl+cbR2F92HD9bZ2SskdbIyOPB+eEvn5Q85AOJoyddEJdrKUAvSAVu
U6K4FpcTNB4KMZ3WT9X8HHYhYGQJH9O+WoZupaW7TG6yAEPtQE6ahlT7UH0pq2fp
ThE7RZRcXVbMdEM1L1I0QnKd5Ufp1lQ6vxqQ9hCMyuoxcu4BCSG0V2+DBrg3pvXE
R16pIOwZmtBpQhw2Bvpy/fwX4vBKxHrtFzxnSzDSQzanKLIoI0j3nILESPAQVwV8
KjnUvXBxbt8fPZk4p4rsMkoPN9WvxA+Vyvws0qr97cnvAMoLqpP6JpdSWsvIdYGP
ao0lWy1Lg2XjMnpr/y/AS/dcSZvLUT0b62X8G26x8TySRVX+p45jckG7ogn0uIS1
y9zh6k6AR5OE/talsIv5h/4XBIPEQ8T7C4Ya8gBJ+FKLZkqJ0SSW9mNlnjRPT1Fj
64mUB8sTZos/PvR6kIem8RE61ZpT1w4I9jCiGJpf5828GxeU9vvDwV1Blf7EXbEF
m0mJQ6lTvxBvHSkuwc2k7bIF022LyfeIgjwk1L/HzwjghcnR+31HoLtq8yntndHn
3qnOD+9vgq/fK9XtnAW/RBooJRdfjKxLHeDnI/GYT1fC3FmPLPoLM2Wu5EoM/2cI
Hhfakgk1MClBCG1ILNEe7BH0LQj4RVW1lLZ5DchgVuDiJc2IweVIYtAuuNuMdMEk
S9WcQIh8SooWZBBsX/fao7wMk0/jETjILoq7+NWezOWzzCSqq54HRQ9Jx2qr+t7x
pBJPJMS0RsAnhb5GYqTH5alljPL3X90PaOBWGOLZdQ/p0DRzfl6EqubTi+Nb9z7q
1AqpxVAfnI71z185K4qcAMh4Hz1GOm0020tRWpEgBH53TVUt32zLySsKe/vG+Z3+
87r/xouseSZpwrfIcSYwYOmf0Zi6/MMjiWUaN3y0p58lTI4Z1gm+cTL4acSFoQVd
UET0yPgvFCbhtQFYTtNMvg/3TaCLZD7VSkhjxUppBXZhbQ1pbwGSte+fAjXGZ1/8
QCCb8p1XT/aNIm6GMLmySIMZqqgFnAGatyBGlofwqTJ1BCzNApRuGjXr5Z13DwYX
1hp/ODprXYnwQCWDso4GRfhIte2vrnXyWh4GBsJYjcx57je8Hk6ylgUz5qxsP9gD
U6FfjqyASBg9gOP4Eyt4H+CTJ7JT2OGnVriG6Q6k/8ibXgSaOG1sqyxRmupAGBEQ
FpbV40DHp2KfY1FV44YEZyNn/e83/agWblPS9CtWk5OsJahRmHX53I2GlOzZwKFg
v43WAHXh1zpRi7tBsbfmzR7711YmgSdU6r5W50cewrim+C1vU7FJiXCeBpoGA4Yr
XFhFgBSA98CwFZRGM3GylwEEdJV/fa4POQiSckHpRGVS6JY6ZStXvM4bQSY3EfT8
fXuc1Mtkm6XXqMnPCR6kMTPk58FqX6CeTceIgWdc4IV4vk4gMuPv83aCbQK2yOXz
fKNPxGB2uCShf4gTib+WC0mkJXk37+U7Tb6RDhUrdvy4sucKhpsUSGoljksG4fTI
AZZQTe1FLnxhPbBdpRP/o7wo+NhO3S6IefErJO+X+6Kr8nWu++ZmsOxnyr0a+lTK
bS7RCSZ2lR98r5+wAjyGZAc1UzGu6a3+jRnBDXYO+72VqoC4tmUTBwyCRWxehg7o
/B5owfPpzk78UgYNckwibZSUqcOJmmGiQ6YmRVHrUGACoCKQXjVEf3cvuZ2G51nV
6DM4qDDFi8uL73yiIcYmH6SsRHg7gVS+WNkUrxkqRN+rOEd6leWFkhC4VvSbDnga
4BMYPB0UwwCV9vJXucXSD4fgbcCKlYN6UO8d7Ckme7QH9A3J/YZVf7zErDm8ChED
XxvtNFSa/2asMCSgImYVTYg0139ym8GYeWVKMawUzOrlesHHCXpOnXFkm2t4TyBj
T1KLKQkgyqdhFoz4pa1fjJLFeepPAdatOaZSHYQV0EkAgjxr98HkkHsUQfYXVdgC
iSbBYUey61w3l5KYzB8KuDXNZrKei1Hw1Wkyv19L7P7ShcXAUOKdf4NBKyr4A9IK
AMQGBJ18IMzWMaK4JKIUF3c3cR+cM+BHbpEwnKodgjKiakF+nDUSKMw4kqnzroSN
9xBMnARmd4jn6ljvpkEldhCY/h4rvllvJ1dNMFKTBI76xs8aWuSdUHagfkrgdlaB
Oe5ddEtZ6Pn4slBzRW9pb7Y/BOQqzu1tpgvhdfXDiSH6WJVtVLYWKFVU8rfbVI6d
6LX3K9L5qKgtzoNzkTtC99wankZHKswEeEL5wiRA+vz+5mqkh0YXN+tn32KLxRsp
46wQYQWDJZt4AzQ3MMYuaS3/pF7iPwwGM4Y2edgmovSfhY8E6wlYEUFEFoXnRGN+
9fszRvHff0ZtxyBCW7KrKRiTinxXAYwJrSzeW5ED5BfWFWyapU3B5/mvSif1wmmw
Zwh9oVo9kABJblNCXmlUPXUcJwWyIkJUcJTCte2KTIfFkzP9dLrZKwXvBixsJ9gp
UqZXef/pTEFQRsE2RZ5IgQbiC71DY68pNaarZiWwMLxVwaO7+D2BYCNVmcGq/GH+
3bcFd1lzPaAGu6OUJsSkF53nPDWkO07wvPMR+bFaDn7ovfbEhg6zOPbYt5QuctgO
CB9sLxYGbnou5f+la0tywgR0derJRwPs2z6DhhA3pgfs6rEawff0iEOZ+GtJ0QXt
wAo0ni9SFQ3OnGAqZF7A7pF6OOe1fYPPipDkaGKOWe6aftP+Cj1YtTAHrEt1d2Ub
Z/jFVqh0LA90MyAyGHdN5vs915yypjyPdcTdXYjozgKLqKhQ2osApj62EDfCUXyZ
7zXuYQh4dm3P4h1NVR5o6nOhU/slVD3+/vSaNha2Lb2bn6sZIeG9+bV/PH0fR3dx
6/Xgzrf70JZHnX009gkKg3PMJ4qa8Bv781yPUUujaZc61VInJn7UX6xGf0OGMiAI
U1HJFIsgsalOgUHpal8GMH6bpZKxNAfj8P9UybCfIzHjm8H3qhYU5YLQbAiWSg/3
ywWd4mbkiPm9e53Le3VVzwYna/2DLxQKuqqw5O9lzw1RnJVmv11F1XYSLBEPj7Vo
42t9k+lB+s5SQ8qDGs5Bv6RTSu8Q+KS3dyVpnaUswDPhoeUfpsjfW4QoFj68iG9X
rPJuBVR9jinwcCI+uwh0gk4+OUcWVirVVZSVS1MAsRuElAyU6VQsjeoI1QrS7JdH
rGb3gcrA7NtOLyt0unOO2Xg/U059/3ayev5adDTvbxRRZS6HZQH0I56gPlZj902X
GfbtbqODaFxN0lK+D7qpu2+8HU19OclkEPvDbNLpbLG3KbBSqX27epRrt9DlO+tX
GaA74/BrIRI31ynB59s0+k5xFhNPpYILhuCtc0gVwHWAuMs1+kjSRxdKoaflsCZ+
TUSIMtoX1UVDZg9QEffhbkT5xoB/EnZXPMH1Irgn6IYkM+nFrszU61weyzdoUdh2
KXuFTQYAxI/5Hoyj18Uhj6sZc+owTmfD2/5A6mbZOgvTiVC4fQWXCZ7rUUIb6c3G
EBAKz0Py0OSd7o3lubpogF7ZHCbrFyDJI2V+nha284dpsnpMQ27oxrMzS0FHA3pt
Oyd1Y8HzzoIB6LxpxdwSJ63jy7LnUwja1YVUnX5NoZ1DLLDau0K+VMp/sv6atW0s
6a5s8StbO6VDXpC3Xm1y45C+6t5ENx6XBDjIm9vpKY47YzT8GJFx339AUI40j0/7
+bee2Mx6rK53FsOzbYYbtSa0jwwRXTNknq4ukEFHsS0T0PxbQaINySScmeb2njQK
Ybdxrr/iCoG2JMu7Cxnp4xyF6RtZawdLp98P6JiUIUqyugiiWipDbDLm/gRk5sTo
UEk9k9rwkja2WvLQ5E4iOaG/njA0N49aOfYSN1gJa2lBp70ytfRm9agu/8nk6MH9
xbwxWQHktV+NlaabcEAfOMms5Tfi/aamTJ7870W1znMvV5Xi2ujky2NzuSLZHbeH
9JuXyt8FP9QSAIZzpjtDrxAeqZLBzjjnj2EDkbih961Mzy91bwxIJQL8F5KhRV89
xgbAK8dC3apciu2xGqg5UIW2+4gkkOtL4JelfrQnoQ2iRnFawlzKmhSGNqumWDPQ
sITLSjoSnbSd1yLDxkm+o1pL8P4v2mU57ZwCujyZMXRkV5KTn269AQCYbOy/cHV9
vId8zmsONvIwChkvDXuk4XJ7FVbMC44BhlVouPP9Bw95edSc3uz0B9wt7QATZdfy
IFA5kZ9HHUnJCMhgJYS+LjkH67tMONBfiytY3jWu85ZADa5DzL2rzMAbW0GV7eNB
WZyUNA1d5zuxnO9/1fV5J+q3e3ADHQv3iZC0q+U3r9wjpjoclTBtgYfuPSo9IOIX
iQhlV2L0GHH45hcB+mrp9q/vumYkKqiXsLAzzmbp4PH7Ie0Rvgh1XHhPJECbbDhw
ZTPWrZBBNjNW9lveG2SRoyxEAd9S5tNtwmhNnI+FPxcpy2C5JXyfTreOgfMbnqhA
rBZp39nSQJYVL3B7EXK+KFALi0S5HTPurGu6T3ntTtSLAgUqiwbnl3XKBx6Tycot
zUc4d/MH1oK6DZpmL9qeJKkQEdLQhJbbxg4JOg0ugt+DOdu3SxYKl+xxJUbhNGSL
U0a82NhZk+C9gYQnvE5pAC6kcpyoHKm4OdditBQve8k9agbV5k3+noJ4u+S+Hw/x
YZ0e7eRX3KR00dX/s/FKc/IGd32bC4j4MGr6gyjsiIqxNPkKivyvNQyoNCc3A8Sj
AR+arm9QadMQI5eYPVxK/x+heq0B0rhYvpw7RsUA/KHdaQKTaXJL/4uImWA+M6GO
0aDSZdHtA6z09dcKTUc0t10QNruRnVcWFBCHSFGUsAfo+rlkmFrV0uGBOEG9ggn7
bUcGHn34tpaTvQUp4qxCvO3hSbj2iy7ZdCUg5CK7CHpqVZy0epu5GZEr1BuMfWk0
rwlslyKUqCpb/58KQyDCmg+GsTAsGkT3NXKBcEi6CBgAWLEDPk6ZqviHmvPaTJLW
zQWpjfbUlY5US7NspaDe7sZKWxRs5QqrDEeMW4P3RdcQky3YExnBwRhD9aX90jXn
ELgHt6Rmx1vj8RF1rIYabUFrWib4X8M1EM89nMw/U4Hm9+6dk5bcEMRz7s+FvF2o
7S2H6DktlBbQ0HXYfSyLSAlXtJn5zTl3jdjfCdLDnW+X7naJ5QQaA/qfk98Go3D9
i7RDeOKzoU5wu1z6plg8eFy0lTNKYClzPfFpvMtY66rF29vGrHj9oJ8GkbvGaL6y
V52+oFVOPwXXYTPxAKGCYHFC/2daNwkmCOWxyT2MoFP3kgI3pSFmL8R9wUdQc8Xh
6AlQEhdjTN2WpngTPVpQFwC7rx45qMgTU8I+xwpI0rmKLrCN8pDzbNXnA5W999TZ
Bxiw4B9TsPqa3GDZNEaEouF5s7JUIxNwYd+159HD7YcMyYhkvLpGzSWM/P3vRqYn
mM8i3WZIolW0L+6qnuU1FguRpsYkTkdAPxZXJXGZt0U//kDUL/s8ZAj/rPNgEcC+
fpjkMov/yFnIZk1cg4qOBO4lLpSsSuAgxQZRPkZOpMyIzotFuz1pjnyzJRfzpTWh
huDXK24J2xkzKqw4ADUC3A02femVw9TUlhNiCKmXHuHG/AFW7x5DviuwlUWfq8CM
6fVHxiPFJphKkuXDn6ZPm54UFoKa5NBUWGowMBYpcmo7xRnZY2ADB3C5wqMRSDZ/
SNr8hZZkq2yYckjeHierwTvh2guS5GhGfUOqEhtTGcw5opyn30qn/vj/r9Y5ASRb
Jw7gm1d9/ZBKDvhEJWYO9D4ZEfCp5CIGbwZ4Sa4LOkZDBn1+lJbM8Q/hy5Efes7l
u2YXbQD5FNCZMERiT/3fP2RkfQLBGApw5ILT7whNg1kd9WD4hlhtZbD2NA/3kVZS
ZRxK6Lvv+LwK105fRJkbEmDLicJONmt7JKiZInzN3iTX1e+azNgB67P3awEySUJN
3Pw8luVopeSi502HHbQ06WBw8OLOfY9Xk8WTwR6V/6/Dqk+PdZ1+KGzF0IbsKlYJ
bRexSFVlzBEKDi5uCPdTzUdHmsxK8ba8dM9a6pRm3K0col7FJqgkHdMJiVvONc2h
PFL0dB02BXUnXvMZkZNzC08B1QXXokc0s82SVMU1OZnvPcrSSKjdHjC9r1tvJxzx
SCbZ1M/1KSocVQrF53F6rMd6DIfV+OWsNglJZxlWOiIHbhLTmLA7RP6DLB/mdDEw
/t0MMKsZCK9KGf40ozeJa+To4pePWH6i2ub6sLj/v5UPG7oQiuntrS1rKfzgNoPu
5Udvnmtc2LnAOSY4JAoA7Pj4IAR/Xq1fZ1s5NEjBm5ER2e5wzmdbXuRGCNT1FuNf
f4YJAUP038IQr0nGmGiPfgkSW8y3yoi475y4yWtLYqA5/c8XmiL9CCxUMCflSMgL
xJRdW7/VkBhs40Viiqd+yLEzEriVov8ZZ0Zo44WT3/BMfh8098yVkmjaiNU5PgFl
YJ8pUrNtRFbY9+dCa6KGKFhaj63iboJv/sUCCdmOA3ZTqzHMz8sVbguGLsNfiDTJ
ykj90VrcRvAdiCcj5TdR6rmpu5m7Fh0z02KQ1p+LmJ6pmEoFCWioQPGNVNDMYFDo
k9VHBJG4y1YLrDO0ILUy0mavc9Bv1GuH55nLqBEC24Jve16mds3mHfTxi+wPdbLf
cwu7Bu+dMZ+vyY0EICVIF1gBWlQja5sMdwmxzf0rf4ZmhHjxrXOfLww6fJZn1y9Q
VPFl1z1ic6b7nnrRIiQh/33kfWuzd1ERg27F3JVbfNDKntpPGQwWKf3EvM1xPI7d
P0d6ILOWXbRQ79t5QGOyRA1oYEQ+y3j4esgFpAbPkHDSD4R7KzdY4nOYes9izULb
F0z7wuIVJy2o3MRjCkgaV/XCAnipROPAVPZtX66NQ85I74RgWbdku+Q08Ikcsgmv
5u0HDbmjRF76OKRTZLVDWhR53YYWlEWDSynRWaE5x+nHbZ3Hei2vkQ/2wcPwFk0O
AOMDYlNWud+tI6YSl45QiYMehHEmGZyNA08jK693w0/S6cRMm9hv5ofD9CTQHdMo
G9BiMsARaG7B/DHQPK75+2JBfCdn53gw9eRFJc/K8hHmXWm5VeI4qHkP9FEqu1Gz
nIcDZYaC5Hpn/joP3a9ibI3UUZr2abc//ZjbUl+9nsd3CWQfnCQA2Qs+0aDbSwg1
sweDg3dh6qnEeSI6mP9l/WEoCk6Ljfpbw3isntr21rb9VrbNY3YfBRlb40hrFTDU
wcOQ41CCbem/+66AyE/1q3RxmJT+DQQLkXC4OPsMefxugwVVRQcmlGzZvkytlBBU
A7LsahCaF1B76YKkh7E2p4amIq72k56WwKG/zJWa14aAUaKohyOaVfbCi8+imCqQ
wu/NwFclYo+ndywlKI6AkPVqd+o6LGAra7Ey1nnXG/Dqji+7YFfDgx/ajyz9+YAP
gvL6ZbuJf+5sNZosJHO3BA9QNgL27uTh8u33okp9EgNBfPkM376EWRjt9AbkoJMY
mggvO59NSwGmwvHqvWhq0Q5pVWHRj92bWQCyOOOS9VZGNOXHlf8I4qjI3rnLXIdl
wBVfdqhS8Ifp10TXHrhj0fFm5qVhPlgyKL82xnpWpv4lCIkzFoH56E8E9/Ey+Frf
QebFZCsqmajiE9PTejdQB/Wjgnyzo1xYsPQaPznG1ynLsIIFtic8cGOIRec3jID4
Wn6h3k7lsXGz1hh21rDLftHNF93dVxUP90VZmAnjq1SnUERlEYko79+g5DSK5wzn
mmd7zE/botEsVvFqr/OoQMtr8EaAR1XnEACmcE7iqnMpJEP0d5tg6tMclshlyRGW
Ln1tn5L2XSDGcXFR8ZRKNBbm0Bg7z7EsICM8SJdOns9I6yldrYsG8tmuxUcNDAaO
epUDSO+9X5xUg4wZssR6eKbz/N5G4yyHrOI1ZgyQqgZF/1Zc1GmrCHceQ9nCNg1t
ouqySfhQXoffl3O2OVyPVMB67s+MVVRSYxNX5XLplzX0QSlj9ZjfFvEjR/fCMCxn
bnBlqtPTYwGbsQRQZPbevDu35/nGIZR0uNP6v++DXeNFD3Zm6RJ7+RR4C0t6TRtb
IsAnem/2YlGugNiU+W7duOfmxPDs/aPnyZMR06SqPk4ZuAi9mf8YD/4ROB2YasHJ
TpXN3+Wr8zYC7lbdGEgZoEVhW/ztSbXMhrmYstzIgDdJfqbHEUjxh/qLmhw38ii+
corZVjEVW3v9Nhi3shdoVKfEwnCdSBQ6n4DXcDDyBDUkqaDyP83V+Q7CEe0AC6Br
J3a8cKhfx/oyIfswGuGSg2Y3bgRcOkzdQA2soOINCj4GKGg5Yg3vz3/akn1FDXOq
RamdrCdcNs6N5tSldtvoB3uXjLXhoRjyg+s5M/Wi0lA2RBC4ebsbnlmACHGSpUmB
O/+p3Gmncl+dAicSqbRbK1+D5aZ73lF7pdByhzmPcErhZ4Wgp0+LMIwVjZm8qIJe
SlDfO+XjhJiIKJyhQhT7IM37nKlSkgrU0wtzssA/9Fw+XpG6A/ZtY9sfCMUsojWt
f9PkbxzUilVLEQlDO9dSDECphLbRCyuJM3IzLDWKRZOdqdZ8IlUwGCI8k8Z5v53Q
fOL51p0xS9IelQoD8KSBy3WLwOHe7NB2OEC1ev/c/HllqU/dnf9BeCUnRLdCeUxL
aNua/I1shfb1r+c7i74w9m2+mqPf3EcWSvz6bb3Aw+E0UgQwX8tOPCtYQ5P8JLap
s6cpkcDIwReL1FfUxK7xA+5UWD5i1DynJ7S8lxMs64iFfLP2P5oBA2U7WTa8zZkI
YobkhooJI6OA9ypNNyWhl2epHOcXvFaYwPqngIzqfGrdqg6GIUk/zxdU1Hc+0vnI
HcceiY5ygxkniWlkUNzlU4RrrDB/39/oldX1J9lfRUNpY+D70JsPi+ByqLUzBntp
mU8nCox6JXlg3dphVNzaCmFgdEZigtmcCtmsh7M310ysFdDE8e9nRZ4pw1B6GZfV
QovKd7C3+Nu8zFu8QO5Zoag+7/SiWfXEAfkkCZL7iyOh1jwCn8JJK/lLTo2VNkn4
EvbeXwa+mmQwXU+VhxvIvUEJvqZOtDi0BwMkRwsImh+DwXgctQ/GqFaC7YYo5uw8
Y5JaS9T+Y+3I7AJ0K8FArN2WQfhqADbK8kHt9J52pC4sPy6UT1q12hUkWKaDBNLZ
qTBRdjqCDDgn4coApwXrJ3VeUCYRvZuVUT3a2qWygHJ0560DrZAY+omZKvFhlvYY
OZr4RydLKZlcPzvKmR8SHdBKtCm7FJcgnFHliZkaLeZC3bRyiQWSV8IJeVlgoBbb
KL00MsuKknVYWYK+ii19OXXAxf4vxTtworPP3cwHYHrfRXHTV5a1lbPIlGposvL9
I7J4SbEE/3eEjN+foaKxv1jwS2MKFem4Vewb/ADnVJUt50Pu6Ze5qMRfFr5fRsPy
5TPq5dNJV8eiBk9bUyp6qiPMIg7aqu31vHJSdHt124BZufjteLhx94+rZ5omqpP9
QKvHJmGnuYExua7dRVOEA86ZmtN39Kt2P60aAzCu4QjpYR09moRx1uj24J1OElv7
lKY1U2Wwak2d7JpBA+tCC0qS5GGU1P6yiOkh8iYZdzrBP1GqDQygYvOu5jIxYW7t
+ELKxEdiCMcbuwgV/+1SX5Txd4xyxZBmOC0m1erEZdFfiGjcmuGtyj6OV9MfXQTq
1H0xvM9DlXsgMs2yxdwXeJGYVRRG7dIpDKnrsrNFqwWF5UkiSMz0p8XTErN8ZKwQ
3BpGbs87NurZROUODmxPLyBVHqOWArfwYGX0tvnGNep3g9DJ+QBIEjbC2e4PHtIs
W6wWLBmkJtEMBpxDe4Rut/FqSI/lwkqsW6HhWl2L8jhlzyl/Dx+cQjqyUuylw2Wd
FFXa4uHLOCblCLc1fe6hWgrzwkP8i3FM154/FGjiyT9gwKY2Pa2GvlDAQTmYw2fZ
mdhYHXSUzbx3WKuuFGadmylTNAFQgL0Cc2ZhKh4LLGedhKSp28gVsbL64Ah6+p9I
ST3I2OzePg0PDzD1pTMZL7fZTY/VR5hrti6H0i6xJBtV5c7Qasv6UBLioC3fpMNi
09uJ4vhKHfAc6AepNPLpE/+nysWFV10jp1vzA97NWfF7M2TeaPkR6e9pbUyo72pw
zdpyjT9zDuGx2RcjIqWpcE2Q3zdwP5S0Gr1okam+gMUNjb1hFz5XgCsmDSKMRv1W
F9JmqC7ynv46KW3MykzFM+zM9jkESxOplZ6Ohseuv8GT5agnlE9+T83I76EEQPks
+YV4y55OhghCX2Rk6lXOLrnQCPSWIrUrZv+d9SfDiZo30aSgkkM3lQkqllJhlTyb
c1K6rTdsT/IFRf95bFpqkyfEr9ejDQg2vbMSAyYD9fSh8t+DqM/AGcAKUJj5d5Sn
9GSCb+nsOcPEEK2XBrvRW/o/ab6kO+qBicZUY7ino4E0gHBVk+0vcIAxbFBS8tjO
TZzmn0fZ6kt90UmZwJydPBkJj35H+v6n8ToDsfUsGOSfTDa4GdAkbWOrmbehQXtE
8wqOvHrwD1zzLH7qHK1znokLCxxBnqx1jAzEWIbYXSZCbgUyq9SVcuDzboSz1Jb6
ofS5cUNFvDU2uG1xm+8MfATNVgKwdqynKayeHH9EmmmvkUX4uLXQ0CFwvO1ehSaP
ZcXcNqxgCUqJjrYip4GugLG9WGn/cr7Oe79Nqq0xmelw7p69zltqxY70TlWXGDMz
lIvI7/cRB9KCu98rQzUlb4VrojS8qjmMX4jJrMokflxberyaMcKJXZ2L1bXGc8rQ
ARU3OBO0aVCI6Q46VoSWjRLgvcdGf4+vwm3+zvGkUXn5Rbs6PsRIp08bwI5PdoQT
lc9EuZouBuGViBuI5Z0/zhVaAhRK8ZpViZG1UnDPvJqImoofTFYYYSVthkTmDz+O
R94wGJLrHOfbVBJ44bEWRV1vKkDwBn83CmV97Vze/p80g1n6QeZdYwJgjGhqk4Jn
MVxX1L8zKz8ex2NzEDGNfzn8Eo8Ajb978KgmXYdTVatd43oT5a2rWv9R0uVGvc1H
mtOM+gXaE+SfL/+BxSsB37uP0x0gB1I3yMUQLlGADC9SHpjE0rigm/PUStSB2YG5
vknp1cEXla1POMexqyY3yaX1mLpuNKfCunC0D10pUY7tvugzd0V5o/kdhYN/MJCB
OzgQKUAHKKjUEqVliISzbrnfnDXbFXWXECp58moBKyt9IhZ76oK2+lVb9Q+BuCWY
KjHSdfmIh5KaQVOCjjfnDnIe65J95dIBdawFkxoo90DPweaPZWw/uvWj2IFMpXiv
Te5pFuckG88OYdMkF93YwtqIMh2BQN8+QdLeSI8tMvub5W69/zJRb6mhntmF68Sk
oAhodlahT8C4oBP97j0e9X3EzKHhUofqboz8NLgcrziBoNzvIl7+u4XuJdLHas7C
f62MqyNKSwJDxHle3SJ853sDTCwoXsXK+8yYL34Mxb8MXJBsKDZusQ6ZX4yqNpoL
O/FHXjO3v6uXtgyugvrQ6YVegaWai+bGiXOFQ5aoCH4oQTTyekeNlM0DpcCZU0HC
8cNaGyTrJKP3UuBzEkDRmzr1F/BCZmqGM+pzJSVRwNFgy2oESVdmvHU31W3MAMOf
vS7lv9ut1KS5cw9T9al3NYafX3ErCOEs8QVnKqjpUs/Zg38/t4apz58TF38nYnua
+2vgPTA8fb89+ZgTWOddyKIyWwBmw6CLVRomSrb60xhkY8K40uZZl5j0mAliLtzu
Ur3bGvERlhBGHb0vu43zWdS33Fh4niSTVXMh/s3zXZDfyFNDgiEjt1g7S4ncwo7h
FJRDVCLTAQcRsBzEcYvebB8dx0LTfcI2x4hX+a5IFSYc4T1Jj2A7FPPfX4RvcBMg
YM0Jje07HZ6fG3c9oXHyo4HvWS/Pd34O8tBzI5pWunTJWhSKGcWAm+/Ix/UisQsZ
secy7Yf0eolSabg4anKwr1YP0uVoWX47HVb1sBD3+IYHeYuOdPweWrBR7n2e1YFT
+ZKLR22Z5VRCJMTAO9l/L+gqWR7mWrEBoVcB7WlGevfdwlyzwuS3iDRj8HpN3P6g
0RjvwfQEjoaXyqFtCiB1OuU/ms6k2wzZOqRtPxsWz1tVSS16DWrmIjtdOtc1KKm3
ksCd/dEdd+NQ0+UgZPF5DRy2DCLHr17DxGUQ+e8HQS8hMKePPKRdjtImnPpwSDYy
sk4ejDHUuuFuDoc8DnClbFP3Cn2fwAZUBNgZPeTt8vspeve5Wg0wvHkrTCDG8XVh
Q58IDmUgz4fbdFlRol+lTI5G2re0Kj/KEKSXFjPXXS9MIYWv4KtHN9hJy8kbcPdf
1XNaVuGnXFk9BZeMNN4r05aQ0j2Bo1Dh39Hp9Vv3/Q3solF4SHxDEMdGCv22nYex
7CjFTkZ0H0BB6MgkBN76ee+k31mxYmG4B8noKE2DJ6ljkfM5MuneOKc3h5bpJloB
uyIGtrrXBuoFc9mNOgrvdhewyhvu9epgVhTROL2+fUU018TNIrFEyCDSyfPP2kGT
hO2R3rn2yYw3gE0ekpmn0iKSPAEbnmlMCf/wuHbsk6KOC9mNtFxcAu3OcLKdwbSq
qHNqAy5RKwupz1CJhRet9dgJEchODBb89qepIkWoN4SpYJ9b9s7/0x3oP2PWDAUD
jh9lpHud0/AeixLAknzEOww0ttYGP4B+DGlVpi+Ect+gJOvbLxFLQ2y5hIGRT3HT
scWLfVSQ4LhGSyql2yFzkxc0LSFp2/a4WCodZWV1XoZyYcluhr3faiSWGlNzGY8s
CCNDZQLRR8bM8AJbc4+JVgIcLY4SjLN6rWYewpkYUKO+i6jA7XsgP/VPU37h91ln
jHKP8tjeXYAKWoLxi6R6I8tRKiHJBd46sRTdIIaiwJqPDF19MAPqzAKR0lQ26771
dOKT926d09hz9j102LVJTLOAf23kOUumHH1KxeNdMWKS00TEfKrzSOOn3INckIFm
Kk/PRRHnim5haB8x/u/WDD7v9fG98hhZXcLPP1FhzmW2sXta/fArQTaEq8ayNEqJ
FUs/H4ujscSB9WJGh5W5P3mS4WPSgW6GR0BEgeqgbUbyPQhn8xpueNB3YBsE9JSL
uGfc/NOUG3X4Hp38tQ7ex0imcZ26DjDn3e/3HcrdtsL7LnvqavgNZcIRz5bXzo2t
haryE1gzl103s8kK57/Gw7HQNRzChEgN7napbAcRghfU7gcPqj8T7bXXZuUAltio
I5fajaGhF92p2YaFqgMDm/ngjsJzs7hHCCfScyrCJgHmEnvS4ZGuVKTPQpdaJmyk
wHOKS+t/phUggRi5lzL6FoXVGuh5qwcqAzKbg0f1vO97Ek1IYUl7INAUJ36zpP/z
1ECSkJwfTCRPkMKD1P8RfpcTa322JjexoeVny45UGFFaS0gr0zQONCQq75TUz4xz
rCOUS5Fmu3kH7oDiLLKFrCGjggBp0sytEJkb/9jsAweApb3IWOlKBS8cnMGYI3ib
1y0EIxYh97tuTX6CL/a+6AQ1Jvy6Ym8PB1vcZK0ikAPPnVEAG+UlHl0kOTJ+sa3k
y2IR/0nTny9nTUF9AMyLL36aa73rZODE9Gee7/PrsaeEjgETc2jTKfmcwzrJkUXR
XjHM98CCWLHXq391iCc0nQwHeHquXe4aPFMz+IxszHlAhrYdu/+yYBr9z4LYdHFI
79i/4ZUihDD9jQKCek2i8nUDRmlt/zA3hO8iN6j7NKmZMz2tG0CduL1gDS8sV9Ap
iLnupkkrM0vWSyDdNl++NfSYej/hd9v2t3XpKbya8DXNdZPE5eJgEgRAm22y7YTu
qg+LS0CLbakbxOJiOhkf1eqx75BrkhbrzpRIkt4RMpQsusv4K5P7Era6Iq7PjkeB
nsZpXXT9QO7xZ0w5w4agydSi+KCQNaXXtB4Wq7aGGMVsNwfeMGA3rozQoo5j4iha
h3UTOGWCyi5AQUvQYTzSQmh1uJoQCvbVNM1xe6vFKNl8dNcNQUYU2fnVkZ9Ox6xt
A1Dz1j/EnWuAnVGw39XIIxtR+uHawD+SiW0pMv0NwNfICBfwAXKn/niwUQtFmpXV
aCC4z/2QZWHi9rA0t+GtMn6x8pEDNn7pRg/ysMWGo47SxGE9sWm2yEbO9KW4hlCX
Gu3XqsoSZkI8Gg3qWbF8Bd79THq6f6aAZQU9c/1DrPOaT9ukIMZWoWiSgfUTP++B
QKYeh3RTEzKGjlRThnuL1OIlabAqI8go3BybW5Qn6d/uteUpoV44j8HdETfoyCxi
eRK9m3kV7rSnyPprDEMpHARo6pFRtP3vKKaDKMc042TssrWxO9NBdB3WbU2XfbzT
S6YVwG2QpiAJo7slFhV1vmG56cWfUE7Nptrcwv8tfjEjy+FbQUCFl52SGT74jk1E
bUm/jwJrnjoDrXylDG9yUUavmF66m3L67UhZinPnCiZB2VRRRBIwS9L6DPhHY0FS
WGwWxGEixZEsVWfxOigtzqlLU9SiE4Q7bSpZelkWEel0WP9oBlHVNwLjeQKWk/GW
4eT642BWztzifVHJUu3Cd6TdOLpmLKMucukhK6Q8jHiSOrlohsLyOJyrWS7iV8X3
+bUUskKVoa3eemc+mhN/DzjYKZ8kPkheqLLqpjmPQsR0A8MaFSRGRkso3qnG9MZ4
KUXvYJP+pyCdN9n8hzctiv2I0NQ7dRnw/Q2EFNvlTBtM3HYQt5E3H7pSrD4LdLSk
TSHf25tdPHC3uyhZOiCiXck4F2En4M+aA9XpRN9kgHood82pyCq3H/foalm9jr+G
0aZwMxJdVq96pj/47p1Yxo/TWrAQ+CRwJU9yIpLT2MsllwNwfdDMvWDjf+J/3S/z
/h0+pYxHGyUwNg5rLBp9oJiv2+A6GNvLu4mjHB2fdlML9HBIK3sHQ+AENMQtbzat
FFgJfC475ZA0l/fVvm23VXx1Qw+8wmzu3QIJnBAWXXGo2ROSXZLxqluo7nvIoVda
JYWUY0DtOZEo6qVXuWiuOvBNU0s07rDd0X53HqPQy/a51sfvBfPiPH0gvNdIe38p
GmaiaVYTyuhDtLjaTwO4loUhlJK7coFkP11lbtW0gcSjZNhLHIwx1Lh3r4gJub16
XseoFAAIX7cOgNUbADo0K6xiAovccggGyIlp2JMPy0mxyWjVlB/PtSk9IzfhgK19
9g6iEg/GyF6XaWPxIdTye8v3GAY3KZbPNxtTvAlot8mXQzqvk1vVDWqQiGbwHkQB
pdskfR8px4bX+XsEdB1JOPeJl2ndi4tKp0NTE6QLENTk+YBrscngiW1C27cnqrII
bib7n0vLtVSw5BFCmMx97fJbBXUWKQyHnQURUnN7cciH4hHsA8CDyVQgPORXaQkJ
0mvdVOcc5KWotvvyzMw+H0RHmJcHs/omoWjkfauICfbTAU1JaBhwTIvVjCszO2Gm
xbkd0eFOv4mCUW4Y+aGySxL8mLRCGc2BP4xHBgdvV2lZqy/umxgSHHHLb9i+IuOm
3QFzYzHOFpgbOGl5L/Zog4iiSupkam26tZN3jgrnC+3xfi2UrVUZSJff3+99aKt1
dBzWLUhhm5lS4J/wqOFV+ZhJNSHWqbXRreE8dm5cdk4nWVc+j4+gLzSDZ41bMI3V
r2Cmsg2kFTmIKb3+WgT9xAaXXXozAGQz4jy6cT4U+tfX4J669zjiMEkz1m/dtC7e
7MDXP8GXgjTradFnrC/XZ8MRLROcRIT4GMYh0QI5b6my/iOiqExb7MTGvx8iNlWj
8dQu8EY67IDp2Rz5kU4Rjcg0bCyINJXCnFe0Vi+ohfexD3s/TNbw/0h54nEhbAaJ
Dr8OgiSBgEKwGEKQ2cg3jCkwqAeJRdTadEyqqqrDEMIqpwR37HFRx2SZgSrSr4ol
K4wsWfAp9oNFuGIeVxpXIfXHg4+kK4CdYDtNeFAB/EuvUOeTiZ0rPg+i1bEJ7zOh
Bymr7Tjtgjpi06/gfth74hionuIwO8cxGwaV2+R2hZmPnMoN46mdPz235jXXWv1S
LqkqVUkHfg/xHrGnBJ2coe3d0lI+iJbXYaQb/t4bSOkXShZ2eCu76rdZxbohPLZp
WCnp2mPWUuUJcEVM3tBJLKisiaQOZrGWrOOYv+N/+QOukDdH7YTuhryqaDJm5g0b
5wcm7LpHCSH1dYMA4s4eF2bumuRunaJu8Ub/DoE2BBO5EOsjXSXXqdddLX3ft0vc
WE46QJK4RDbOkZntQlt13OIqlToC/mevoyl6V8SaRLAlw5Gz3vOnLwBDIgvwMB2k
sg69FVHGt1CQVmK+dYOj26NQXtBP/qxCq53yaT5O+Z9txsKWrIeR3MOBxvyddl4f
GMalNHasoH3Z1ggR0L1TxtW5RLTe4WpTQXed7294XQ84RyjbYeM9nqevM5NrYqHI
IB1mpcstI4hEz2xwkyNES40eTbijXnTQdhTpnvR7/GZh67iHt5cvWOmSDHbEuljn
S/a0SiNaR0udvieSRz3pZE4lqRVFxH628I3hSTMyaJaeoMwLGfXZ0KBljeJOqR4R
rmW1vmX9LLWxmzjl4dMYbemmx6fibUiQyOMMekN0FK5vQ2A7v73SBYvUa+ulEfVn
eWYqP/v0yAGwjto7bPhiaNnIvAmZTAXdychZW57iSzPOAYARTeadbIyF1I1CRyAE
aUlBOI3M+Aca/hAgXJaqInAmf2Thf+H7bLJYk/grcjTVfE2F4Uh35tJfheiFO9KP
LA64yi0lRUPIrtoaDKcvUZYWsTPF2gmRD2qPyZxzapPPItcS4R2vWBDGk5IG6bcZ
zVpYpnYrn2+ascrP4pNwb+DxadU3TnokkYdrTyj9g31OI99xtlqauOBPAIhlvg0h
8RaNiKLwTCXhtOSDp1VGQ7q4jr4+Wi99INkZov1BYRrL63Ku8aZhr61dfOGFQP77
WuQJ8DsBqnIzluoXOH8b4Ko3iw8Dow8oxSw/1G8y/ytUChX99NKTf4+R6J+Rt2K5
GoBRjOVz5cjxerK5uCY7zw==
`protect END_PROTECTED
