`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBAETcyrfsYxJLj23wzSAL4f1l8A4iQ1JXLQhr9nV8ce
6Xlp+4jKUCUcog41px+lMEjbfedCVdr9pf3t8RY+oyY/x5YtpOkA1moi2WW0vBSM
hDTbBMIwWOTSJxUIE0dqNohNwdfCrmt5mAdsibCJVKWZoRA2jTpEiyuQIQaiLGbc
HMhZLbtLBQ7bckfXiDLA3ZP8nHYvB7/kTXTG4kEUaUatFEugHenSnneOUjz8+Ydh
ADdxwCkGZvepndnuA8R5/Ct2wZM355oQH7ve5kEcpiBm2trTAFwS0Vtza9mb1lqF
RcPwG7MaOXJ32L1V8oLn2z7XAX+JLiiIHmuz+D/wOzG1FjKTSgrb59dqtomqq+6t
V83EltEgBe0w3K0+cVgMWqV8FMYanV7OtV9QY6IFXrrRkrLFKIOXRJi9LS1E/RlF
APlvV57oYQHvryFqLvzlh8GYGUvjHd6LY30wpROq6kgxmCUEvaRV533Zoxbv5Twf
+/kfmcyr22IqacF7kqKcXDLG4JNOGZ3JOlCNIzWp6uowC82GLusimdxqJemxydQK
51cFV16NBEHGZuH6/J0Uo/ZlkPcOphjAVeGMaKHGkPBjbEj/s7EB1Az8F+4/AKck
5E0B1GBiRYqduJqBEGA2JZQsAAidSiIobCUiwHe6evdO+OeGBC2MNy3B+UL9v+Co
/vkcYlMHubKpRNumXiLgoO1LUsLsamIa8+N9wbIfICdWhpiw9XrvvkUgJdQG8G+5
da8iJsAlkiiECVXREgUmgz31EDEWbIafqkYfZim4ODq+aYWFhE2TbC7zyZNw3NJF
xrQ7hmaB++Lo4W8LkFgDumDWO/XV8r5G73QYzzIYWE8=
`protect END_PROTECTED
