`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Dccng4ouCEj+GK7eiIcj+6spaq7bqBbpFQiNSX41K4T/G/mVmsmURd8KZbvBSt56
e/3p0nx41WBpblJNQG9esEgd8bSEm7cDECDjId3InAxVTejmOlYdF6mNaWswYxMf
G8FBp20GPE7oCbc34AzpX1zQ9f0QMl2CpqG6TtKDSmHvlUzKuLjVQWHDYHWZDdM/
02dkrbuIVMq6RFV2HsVYsgkwmyvgjpOgvL9wTd8VETCtem6hL78Y6wFWbJW0Aa/T
W7LL9Zzk+2fKIVD+zv7qvp1ymATxfHc85mZ5cAoE8XOdeLTj1A+q36rtkd6H9Z9A
wWJt4V1/y8Mpl45R0eNGS2X1gQLaGy2NyQlcqOvk4whfzTVAnb+Y33kJ91MwqZY1
nveakw+cneVVopEKn0CQs6LB96PUMu/6xCRQw3HYJ1HT94xopXQpQbavVujMPcQs
9GtYKcPYJrpt8nsXF49J6dfmixH1/it9vrByMEez37OB116HFN2NhOY40IzOwxQR
v6nzq0S5yCioZ8Yx+ACjrd6+RzsFjtmVwx6rGfom2bqlkCzVGbBCy+OQE4+jNvRd
Nl1c2pHML43Ep5ItSF5spqTkAnNk33rfkXTUCVrxl6dHzzuZfqlr3n4sXV43IXmw
TPbE/6jNwHHMXNAhK6IYPuhb98TUN+lxUmZYARXWpSx1DyMpiQdv0Me1OjbDLeR0
`protect END_PROTECTED
