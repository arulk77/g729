`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46+laJXqQ/DAerBK4FN5unHI6b/gnYq7CqeE5dSmbCkg
85Z1DzrrqxPySxAKFCM+VKiRw9UVC7z5auzG+x8/sf7yBTVq1oohTemazYgPegHw
jhQxmAgBiX0HWdG7OzmcorMFE1RR9XKxpBtFAgoe2cBKtfjkRgZMFS+RgJENbY+z
oZXg3H7KnvdMplCGVq8HZ/yu5gzX66xWd1CBtVeMg9u+roid5V1Cp55Nb5VwXr/U
tV/JlU/YmWucgiWgshX2kGQcEvK/a7ADbEDUB6JlSTuTXeOZQulYe8vv6s2dN0MA
p7RwWVpgjjtd2rgWwygYtSCZyZOURX78QDXN80afrAKEt13iHdZMG1o2X42XWsQG
041p/nUR37fATDl+nLjhcH1wEeP342ppNPDiElBEFkrxgVL5v0SNAqsh6PoWJ/Hh
WczT60gSVFacC4ZRvJMXRHnfW4thAwTwppdh+aK8NgkQRIDN0enEyo1RauKvSITb
`protect END_PROTECTED
