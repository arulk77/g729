`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGWbnmrWC/OfqW/DYgcygs7X6m3WboTDoI6pRcH3W9Od
quCJFDxds6QBGUuPB2t1Cv2dIQOJNgy64878BqDKmyvd7zBopiMdcfO15mwpWfCW
AO04l6QahP8VWy8zybb1w6E1N29YTHbtgB0kyYnS62HzxU69mCR9icULZyImUGMw
Wzv73nSLJv4+YINxMIGCXiFAVWripjzLjc/v0puirvK4TPbZb8ex+0wYJawhOeL2
a/njglFPvurvUNAHJqso24f3m7g5Bmsvs4ZD1h2BJOljPgYFuik9DPnkmkjP4s62
HTaWBed8F5tyAl+6cPLRDDCobhWe4gnsi5LBpGUcg3qSjrYODwFZVTHSfyo3vQCS
Y5RkDc64Y38IaxDt6WPVb0oSfSsp/y8IJxzKNLTW8AUN5npizFyj0COAM6DEgEIU
6ZGvC2heBqt2Zy0too0erToGgwaibA1lgJwACj8j38VrWeXMRpcMmh1+DUaAici2
tdkKdDYVHa28qYGdK1DGzRltDvl9Z2uT3Jwpa4kqbdtv0Xe12cjD+xVdaXYbuqbt
y+DyaLzmkqwXuqTinaZyUIzpMfamKmBQdKV5F7mkN5EzKz2/XWPQKPyEtwdheqZk
`protect END_PROTECTED
