`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN5SzRRG/ChQC3hmoDwwRL22a8XeVeUXmCbhLopdmrJ7R
jTDa0O+F0DBv30jdB6ZlxGk40Uqh1jnzUsAbHJYKc0KJRUVzMXmkYio+irQfcAmP
/6ZpA4Il3koshmIazmier3g4FdZ+yYVFyYJUFzpygoxWmca6oMGskK3i+B5ze3n8
WoOE7p3s56Ez5ghDOff4EghuOk6SKqXvzXb64i9mUcbLYG2YihVO8LU/fmpalYUU
vwmSgHzgjZxsUMXtcjmR9LSnleZq7kcNjVHC9l5JRoHmJghkaC+rT7wcJtI8X/D3
IdUXbjjE9iUYK6UxcbpQYy6PLiYiQUU/16xPvRyjiFcudZb96aKUP0x/LjukSPaP
yLaKyJV6Xvp4rmS90/PTOH7/Z7QmF20wyS6wbR7ZNG7CbFEw0rQLnSyqeI19OApb
DYzv2m7MR18fSTA67fRNAcRc5QkigqesSUUnM/6xRb7jrMud4kTsRt0C1gWDmUXu
H6qgBP26hEbbmML7ixVjlZyvV5au74NNCZ/jANVZmGev0gYtbMtxrynvU53miBUs
MqCE/Cyjgbs8s7SnwKllGSrXyOmUp8hlZxp0HRpS6VM8wFD91hJItgdQe0qL+ZFo
XKBAu7HETWuOe9W7pksGg8PO73oZPshkHVsfL4QXxQwxj9XgjIUlgzKsCBt6fWye
yfj0D2t381aZ18hOK8B8nsTuGlvZ3yBOAVJx6zO6XU4Y31WK0wf1wBAcx4ANUKQ5
NLzRW7gznVfZeP0Tvzay0XmKsY2sbQfheCqN1cABMJxtS89fMamRIGdX0u2OISSC
pS1Q7C3KnxSJ/hy7wKAN6ZBh0FOuzJVXKHi+EEwHTas70A65MZSVtiQQy6/dOAY5
WskOp8rJG+vece/un2EZa+4vbzP863fqXuTZOEwGCUEJYa3gCaa2gqytf0KsPS7I
eh8tVpZdE6fzt+76SCKwy7ox9vERw2JDbnCOj+PG6DQ7xftL/qhE8XcTrkvG6bC4
bSXl/E5XQcio8zUHAd0lpcIC9pFXmyRUuA00qnDZBbGm+1ObqmD+AtLm/8erEYYv
XQ0afQDKaXSAPC6NBMvLmGyLV27OXaIZY2MfLJqf+qX0mg/JT2vn2AKOEY2JcM64
raLWT6k1rC8cYhugupnZLdpPJry5Q4/m9j/5/UQ0/hS/zin4xSzz/Z/clztSlfy1
QZzdfC/PNsDH6m3WmOWeeBiD+81lakRGuM93oRU7wjnhCTFdvgLqdmenUGaomQAB
GQJPSrTCmN487P4Woc94LxX7AG9hu5ekI7tK41t+DyqshnEwqtjgGdx+9cOZ1kg2
UdSYTtzEkvfLL+5SiwnMNgHSiqZ4B0i+tNaVrybxLLshzMcSyF5gqrq4FrkoMjWL
Uvhe/40EdA2V4DaRiFy4HKKmbREOvRcqp0WvZfUO32fgd8nB69oZRe87dJ9mEAzb
CJkeojhure7sb2/d3FqeoRDY/qtvfeRHJESyoAfa7CxoRtNRGB0PMYNSGCdDtCFE
OI985pmoT9GqjKY2WPVrBNwv2CxFq2/jTrdcW3CnGq20F77QE//v9ZYlt50BQOFP
ZWalxZLKoe1UpQ1GZWCLtZGE95oW7bdedJfnAdSGysHNjCA4C3Bo6/dv/hqpf4WP
L38nmjUiLtnyiH+wzr0rZf+9JU/c8wrGj4d2OEC4o1Qx0lj01Hc/PvnzDK9QzSEg
pz1Kno6kbLfpmnXYAYLp77aI2rUMxGWi6vbgUcwBX0oo8XNa0aB9x2Q4oCflKriv
PWfwHPCV5K46RDNC4B5J6w==
`protect END_PROTECTED
