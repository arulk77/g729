`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDLFAsKKExYCWXvHny+aTJC7KDOM4N8kkGBa2VOGQoFD
s31WuZBRXFAdewTDZFe3pqJF/jd2+ZTwaAW6u4J4F56BPvPwUsWH2BpdNNmltgQV
+mAaSlkGa5ZEXRIUcidPZVJhwH3CsBii6PcUVvRGjCl9ipEGvI+S7egdmhdCDW/M
OcPVGDBqO4+FQZXtUfWY+hPsoWed7tVgyMnU1BIvpqUOq0GN1QA8dFplqD3DGn6W
5XPTFH4Ccv7w+qVbmXhqLPxL+xA2fZ5AlofsjWsw07U+J9OiS44Zrh6ASvJG2HpO
A4vjVRYk71ebTwzM3D0ViTSgkWwNyjyyfhhlV3b9Y5mDIpPuSuzmhx4vAHKWe1Ng
H4FHJAeRw+3jhS4Vfr104PRvibw7TI7vqomx9h3ctuiWNHKiZiLLOlHNiQzsxEHD
EcHsJdkcV98Efz2h0QILpnTy0eUh9/gIR4J7Dj1rGE2qwte0N1KocEeJ8oMI/1vQ
`protect END_PROTECTED
