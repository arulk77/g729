`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ab3t38y2wf5+qsH/48ktMEOmp2HKfOzbKhV+/adSrkxuFDZPZlq8Gh63Ry1ONWX2
k8CTLIbL00YWGtHLdRVXbZes2Jt0l5++dWDbkwlS2A+3xZTcaBxoHYoOL3AGRyIe
g/6mvXvnOt4AOcCPcv405wGAOQhNBGSLl3oUT6v6/MTPzSBwBS6XIDNBiem35Qjz
SO+3Z6PBuiARRbL3SnjXgU5biVp4C/McWbVKK7NQsfdX/wtMOCHo89w5SuCM+Pt0
zOOotJXWuv7pbthp8OeuI3MNH+c/kbF6rQKt+pnCOnM5OjdGYC/x8doarfIHlARp
bRZC23YL4IgfV3y2E6IWPfzJWT9Tl25GiG5iZvp88hq455dBTQT5BjcoSk93HP+e
V/WF9m3sFl19YDk1H2noLqR6Zrn80hLtoF9o0kZA/nY=
`protect END_PROTECTED
