`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aQy24ZsB2+xsudLDvkv3WJR/XmWFQ+CYFBmthpIjjop4
SpRUseC+lHP1bGvraTKSweg9xf9f63mKsOSCU12xWipJGvd4wUySSXvJNgeqBQqM
Xet1lMMZTJCaeJWuJlQNwWG2bply4cx9jNvTVMNMJmm7hN5Wjapcwm4lLL5K0Nxh
ZFEzgDGfHiGs740m/pogo+eeLX+IXMtY+bp+Kzel4gPdoHr1YdH6pLbYww88x1J9
8GTQxJ8stachcDHBFYMv3qW8C3pc3nHMsMsPa0/Gw9DwZVobPG3ubXAJGAndHxBp
kjn3wXHHTAdWH3p3UyQFguaiIDv2lSaKBS4wJ7eTchqqgDizzuOr1E5WLM6++CTl
12GWNOFnn3MR24OrjnDgKRx3ODwRlgWRp1bs9GHGtDRo+bUzxVEnZ3wBNT3OgIiF
`protect END_PROTECTED
