`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SXOJD0cqxLKKNnezx3fY3+4t+7yXU8MMAlC/DoQloqKq
4YXQDNLBHQy1gWSEBNWVrQgvSqufykS9R3uOCQylt50OwoNCc77k4OnuK7G2rah0
daR+/Az25Csr/fYSTYE1vT8hp+InhB2oTO9zWFfdel9cb5vA+4TZBDBBGyrK3Mlf
7w7NFS1rZIme4TKm4Xp/mrdBB2bQJwX2NolOzzbLvGtf9Ub4MhlSyJ6eWUB1t283
2X8B8KRoejKsIP2z0MWEJ6BNS6+xdpTGDBrHwiR5o7ttsU6SJR0OkiWx/lRlLxiG
wMiMsE5LUoQuEbkT8G9tf5FCNIIVXNOeuc+kceIFquRlRJtsnXa67s0GZ8z2Avix
27ZwagDaLUsTUWUxoJYAbo3lFZJSf1m/FaoGRf7KNyCsxbxiHWIfJXKXbZMUPKo4
V3wzb5dZhnfnh29FTYLuNcHNuMAwa2LX/UUSluTTpEj7gY9i2cyf8VZuTGyyje3F
yottyBoAACTwqAKcUVOOQb2Z6YIyGM1bVOY94dRd7RR+Nc12aOgUFeau3SzRYYVJ
xAylBnvPvHRN5+MXw/wy4lpSgC9mgo6NtjcCVlxj2dNp5zbLywZObTwPnynctHlz
mVbCsGt69c3SoLeHni3K3tedx0ysQGY0DW3w7h5LxH3xwIreHrdh5yUdpIJyTBo6
WpkHOSXHP5biZ+GXgUsdVesdGgSV0LNS4hxUx9/V/EuGUcIuv8kGx2ASl6eg9n1h
TZRqwf2zb85HEPKXKcNWvTGja7T4z4I3qbR2Z3mmnPbVpA5F0KY3NRV0GkYhoJqF
MGcL7iNSTIrwZkQc7AAyWsu95RDZsvDJS16m6iDHzHIjNihPSceS/Q8YwUqceNFz
Y3jMfFcDLsasCDONGJOxfHwB+6yLk+NXQg9osWZe8hz6BAfpAJrZdXL+lDkStVEW
/J83/V49EkRtmYVlUQZ8xsSnV7q657Pnyi7K5NjOvpphNaOCYZ8peXalMCzuIUHS
PIIG6OrsBmuVa8zFsZv6OCbOzWAWO1N47WbsCseYFFVjhk+Ss0FFQjOiK36Q7I/H
4rxCmwBtoiTEQ/nPOjKtN44loA/KYLUwzL3thdsm3Zpk4CX5rzKpqGNTHeRqQ2zn
dCBgjw5ckxas7ujWHYbLelDHvZXhUQ4JDe+6Sqv5ERMgMyQw1cs+yuxKtNO1rDXf
MceEkwSCLn+AWXWPnb02Kn1hej5bdQ1ONt0lNWSCHM+Dv8WHrfB+TLTDAxlbHefg
uvj1/xNRToquuQLnt64c5Ur9qsSPoQxsvWmj3JNyuRvAeR9sLPoQxhLWv4ryFSso
Fk/tpGRGTeoo2CH/D/5qnXFDDlsY3yTpkrmnat5efsQX8jAd1/UIIUyjHQl+JEiM
7+OS28pbBwTz5fyWs78GookN6130LW/PDYHB0KsYM799YuMqjNuB/+eHWp7rv/OP
YigytZnX9pfNjb+dIduepxNbxL3rR3mVhvzzoGmr8BMf+LnaGjD3LknPc55J/iz6
PzC7IMQsTs+qrTSi2xb1UkFkpgTNcdsFPhZ/p4tyGn6TwQH4/oe2RJcRhxOf8OMS
Fy6MXZHyihrVMfDL0lOSq7yuCE1d1GK3QG1uskwg3B3F1lvGXOUFQk+IFqSrI/ka
EXbqo52rO7iREeWC5LJPw6uyVQf+W6jAd3xPHQJSFsmmYZAJZbkowJlMjpYZwlPg
a7QRoBhz2+4RiYsPGGVQ3oEkdtYwBQ7p+qKwH9ruyZsMwdTbeSXZ0HB8uwhE/sqK
7nN1/taoSGOJqihEMd5hhXausRusGnc94+W9nf1dn4gCvaJ6kb695K20lbUuF/oj
qkdkv19BT94Y8Pj3Ghx9DiScM6CrmONTkDkduu+ZE2bhyJ/F0BvhIFs0O8cg5fwS
mNFz8viVjeFVxh2eyIa2tsbmDgRjI29/pr6PTPff7p2kGUCYWsWneNmhrmMa5yoj
r7NVG18JmC/X9T1G7k3Fw6wSdWqGK9Ylu2joSUh3qF/XHPAX8g1po8PmYp8hP70X
vPKyCFhKpO9rupqppKgxw4x9yCq16POMXlEdkfcR83lx883BYYxVZ5TTLwrnoPLo
bI6SdsyzdhcO6yUygiNL0sVRncjVDJiWCM2jUN7Du6zdnP8+Sp5YtDZ73llABxzG
AcMVmRlY7bDhTushB0R2BzLJGB2Z6P1Hxh/tQr1b+mdLoly2gOv3n15oEFs7Bl9L
2YdlYMWZ/am5S8AStn803pQ72MQ8Bnv/C52Au9p6GQCFj87uODHQbswpFNty19f+
mdNpq0Twx7l9tpzF5A4QaWQlbrfhVrOQCdFOTtCI2b0xv2koSsc48saSyJM3LfB9
AnEBBGp2bexdUvUcNviuYe+1YqKf1nlTiX9ueMTCtuI=
`protect END_PROTECTED
