`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+SimstdWpJnrSb4XsuPW8aGm339DcD7FX4ElvY6VuDN2kDcB/4fca46ZwCkFj/2x
AEruxOi7VLGo8y5kI2t4jpq72nXyRfFiWKcMm22noG241Fl95RtplNhCt1f3YJ7f
/GglDzY6Na6EgbQxAxF/cNzVkQ9ouQhiqa6IhG7qRbcK6A5oyBMSsjHLIu3Q6CIW
vaPZdfEArBuwDP1UNiLyPSREDxFJewHLnzmIa/ImYlncBAAIOpaxs4Ib/rt+2iMp
FP3IL1+UReDV/31uft+42+mYKYXkzJxT8qEJo1++IJgtnR+/hI7IkrUd1SildlQR
9N9ogzC7kOGBAnfkjYAwO+Gm2vTpAI+qVoyPpeFHD7I=
`protect END_PROTECTED
