`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SdIY/IVmClW/4+WRCxtEUnlwxcFCf73yhtCYduCJsQ2G
EDMF034DX5q0B0W+CQDfZdwTgfYdbevTbmj62apuZErfMgaYsRVd1y9WkZlK/C9v
cpsD54vQT69kkDSks+NrDIIC1vNATmO4x0BReMvj+duYmXw6Mb5LvLc6Wfqwv/Ya
fyJ0EG2EaB4jRJq1BqJV5BWKfEj6H6/Xu4fEmkT2wL0fKVx03DY78/sZ98qZMe7N
hmL1Qzl+SRX1MU+xX+MdcMy+7VPDdmDwUpYTr+4ny3V1JV0YRC7AYhFKKbTTEc/z
Zgl3YNyzYJJ9ddMIbiuYcznICHK8GfJnFCJ6H3ZhSR7lgLBzX9eh6vFpHuw9LR2Y
v7sLJgY/DZl9Pfbd/x67urt9I89E1LBk3amCo5cR3sPCZSM6nw/aocKk869a2Qmg
XiMos/0W5ZHMmixcGLgdY+nQ7iSkwtoXbpNSGJBS4rifdmeYIX3OyKd1umtTZwwM
hqwZz6Aelr3nlFv6cJ1ljcOHndLzNrmmA/PE9hLC67ihDHcWdBNJygKUjct9NOhX
SMXSWMWjIVqMQoR7fXI6wQ==
`protect END_PROTECTED
