`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C0gYHioMt1jyC/QgWkZ+yUzstDDRxA+7bwk5fEliJ49Q
M4Mpp0K8gQcuTHDROXN/i1UZeE7qq/fYGNRgYzEDJFL2sLOmfvp9KaeZlWGYLpak
i7/MwQ4iHvEOzI0VqNRDGmN3V616AhGt8raerC7XqVXQt4hniBciWc3Df6qRhGAZ
7giWHtnB/vxiiBc2xuDTSy0xlQ6L0IW1LSRJQ0CKXRr5JbpaA/fLQH/Bkin3Ltgo
M6oqFH6a8JE7qzao2GIee7Y5s1+uyg+ntENbc09v62drGh90/aMILbjexG9fvN+K
+K7hc5yE74sqcARIf0c6GI8QybIcQXRnBBhnUNX+xBBII9A8mgOJO/GRP8CNl7qY
cvFklmyxhsZWJtWAvTmuvhwXFu6U1nnUN4CzuoBstalmpLXd7zSs7I4kgFt0pIxC
jPxgwiTWz0GtI9Akvl/NzF+xkP8zvoPN0ujf66S4vWwd22/tUrjcc5nYwnZy2DnC
y413i3z4pCBR9TcbINcTGFlYtKhbPrNk3ldS91Rd9C1BdE+c76AysVQtRDf+FIQC
6msLEE3vG5BQ/JCREn4KCcLZWjM+3itrFqdt7kkz3B7KIMqnKwkXJnaCn2WAoW6v
/PXKrIKzJPaSgac11gAEjQGnWOJA7pO5ayAn4Qk2sfk8PhvpfMOSUmfE/355nImK
K8RXF/ALfFWTbMGL583x6spwaZJJjU4LULSKUnOjirVrAR/+JNtQzv0xNbmrAbgg
yQdNveyztB87qJH2SDMGKnFYs7glqNpDMvjatnWrhiTz68hto5U++UlCVrSs+51b
8UmnyjYjicxb6nggikh9Fnj2YeAlaYUYxzW8CNU8JZ30qLqZ4yhcKunWWEx44RzO
U29DVis1oBrObwkS9+nrNnZ2rynJZ7rVajxveP0B8UTJ2FDxRp0jY03VJlpO13r8
26O/SzytyzI8ena0OdUYr3VBPFe+hEsG/2gjBFds5omVxJFGvfX0AGW3DogIiXDF
G+Jkdu87SkCADb0NYWo4jqlol5KeC0AQuR1csZ8yLfNvYKcMGuTRj07OPQUF5jD5
Vr3C5iMffFKsOjdyoDgbiHwqfjH8rMbP1IQCKmmb6rwUHf0H1CqOsvE/54Pecq5T
FlooBJZh3cBpZm15X/frA3/I5aPgNT1ieElHnR4pS1cpM1gQY0L+se20cVlPWHz6
DQXN31Uh1FQQ71dw4CzyXY5Wglbpsyhu9rttbAtGjA5apJUUcxjkyqQMAz90Q9tA
80XEbD2XDUS5efgmHg0aQj3R4938MFWzqQenrq/l7TXeKZMPrJDcqrgfetxOpIb3
PfsC8scOQcsbSkujVwz//WyY9zgVM7oWF6q2YmpmALvNctjwbvOYQ7RBIb+IMwnI
c5GSnlNKjevvzsiAJK99tDzpDWe+sHvK+fLfFw87Viwy6c3n3ulb22Imx7pqQB3h
vnTiieXr4X8zLMxWkYsdA8rM62Hsz+peNHouYyN/IR2ab3HIest7rUQJDH4iLgiG
NhYJ4YMnnGfX2BloyCBBFF+1s/BD1KDqgxSMlbDdtZbj+sw6pN2l0Ehvxp+u12Em
zOSlStr6+zxtr/jvVoua6qd8MQagTrzhkV/TwhI6POTkk89aH9t/Z2bZVHhIEDRi
NkaSMRb4SxXfD6YkPWuZO9yw3nQzQGR6lplhp4oemnfsYypPHgVQ9XwcDEIZTlHD
aGGKdZViKa1tK2BOxgEpMKf6qtifyQB6DG+KfPjdm+WArKCuo3TMfivafs1Wfn+H
MwTZEX2Q9h/wDtvvXpf53epDneBGnNz4U5UPJNDH8qd4xl+tYSVOG8a9l/aw1o06
O+gT8qnTEqFA0/p6WwBwklqsmIMB0hzcXtv0O80e1fa96GUCoGld8J/Re9vFsDk1
HaXJwW+lwYk9Q6S3FMrfs5Qq7pPLBfOaPE/Wd+NtjGUWCQYxnJ6o6XEyz9xksQUF
ahpi59ikrFcwJKPXIaBd3fq4PPw3ZUQ0qDs2LDqjKUto2XDz8tPo12wz1YL1s5Zc
SPVrsL4yG6DNBB7UwCsLuq0oh2hXrvwUc/j7XlWcU9RhTdc8Cftp+jzQAoXkn8w7
jYXeiUjrvnNZwuB+0C6LGGDajPLLh//ahZ3deP0TYhqHh6LTVlYUPLaTamkubqPn
WW3LpN71z4DRvbQAlbw8zQ++YkuDsJvG6IhcpgfkELTygPB+qKOl+9KpPufRnhUe
Zp3oKcBb5l5CW5t1l7c2HgroWVRY4QrmwmFDPXse9+ZYQYwdHgwN6UmkN2rog9Ts
eC9JHUoHScM1PlBCefonPvkvN3NlkXnp2uKIor4gc/LI73qe1GsaetTJ2omus1AX
SubXUayidhjZQ1vUEaVIhChdYSI61+Co94+iHEnkn36nkD8Uswhu2ZjvJkrav+C9
nNZo0YVzh6BC9ktmJj1d9Hdn5DdQTAu9ZDoi7WUvKednd3jLwblRfUCSN+gOYrI0
dL5wYGA1s4meSi4may7LNzJXwl22IIj2HvHiIR7gZ3FSCjDeVPml4PY3gWui4rSg
ZiKTZHVI0MvvedW36FazMHBiYpCIHOJzoh6CsmWZyVOXi7IfwBxm0bEv5EE8fM+o
yFZDKKZ1lfw8u7uUJ+RpVf62bzo0XBEKg0tMn+009fiBuwcudCsyCSZwcTO1sMB1
4JPjLLEGBIA7ucTFVEix86ME3zKUhGnxA2ypIXz5/bPwp6dYJ7ydbqhbMH1OElFx
siARZ8yqU5AkL4BqhekxlrH4LDCBH69amP49XQGSTl2fiOlKVBxfOgst3JgZjL7C
HmIKMCN21qg4xK05gl7+gf1CrgKBMBtN39bQzlDc9JBfRW9ZD2up19CjfMbJkqv1
tQUIPrxTPHaQjNW5CdR9OeBu6d30w4k6GRRLMLv+27fjQwGHy/BIgaVlX1y4SDtm
+inPtQmVzlDIg7GRmjzZTdksN+ei5be2bEEpL+WczRqKoU1O1Iu5Do36HNsxxY1O
OIg0abTxJ8z5tTnL+ZWE7IG9gQx5LFb/gvcJ3dt+hjmIFqmcutRefT2SzOuIZruu
WzZbfEAwzxqt1uH8qKPsyQhpNhCrxSYWX6WuPCltMefZc9Vt9Af9Cgd5gXVYRMCM
C9TVZURlrYU8SwsClCpSzBn5xG6U48i9ubMx2dN2ItYSPMC7nL+pJy6bwVRrEMsp
j337jKPdAaMgF72/4GmMXw==
`protect END_PROTECTED
