`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ogxkQp+tKEj1NZKnrQW1R9Yc30HVva50Air1W1WesDoRCAH55X1WcKgSnjPeoSm3
jJfDVBiUwAv8Y2GOSsMPfKmrbS8RzFP8bODdHItvUjNNsMreQqGz3trck/GMEbZB
6jZtPNGNv8gQ/37aoo+HAt47WdasIVg8cZHX1yl7in2mFCQGn2mb0dnNEe+dN1Rb
8IBFyi2Cte6HZgO/hVhNph0VldqCDACZ1JzDbEsRDfjZmoKh29vBHcMz6UUBpf4J
NSKLMj4E9h3EaDAxAXHjnXOAo/34UKIR1JBIC/DCs+o=
`protect END_PROTECTED
