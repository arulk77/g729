`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveE0OcKZvKAd/6m2l13EOBQ5L/jQd6rPkEMJVmaFmc1Mj
6xUqt3P8UVPT1laMUm4h3EDxCCqlJW0sYJh2zSvJhb9QDBiuijM+TM7vwlSmTHYv
t1x0+be52ketCvb3LJdc4VYuqSClBgV/m/5kUSVdo9XVHhiE+djPSNTEIdAYQR++
8CIS6JjTlWed0Oj3OR5z3Q+Ql5PWDCG1bRiSTPhMCHLqNul9bF/vjgjnFMdM+sGw
1V6HZpP7w1b9X90LS8gfUXX5HH4uvaPoKq0TEs3xZxxDM8kol18kAT6NEheyLbO5
Z+YSVozKHcp8eSLy8ZNpIq6gh7WVaB46unP383yAHmKWOo7RTskBymDX5Jjjc8lA
e4ahPBUNYXUXnBIlg09H8eixuPsEuXDpa62X0RzULTkKpwuc27GDslFHvA2k83oJ
1YMA/0w1KQwVrl/oeLjjHWtkyOl/oAnbvhvL9sGERGnyCSFNIom1rmtIKTOT0seQ
`protect END_PROTECTED
