`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
eKsnZEYoQCBoCQntARfm376Cn0Skbl2j0wu6KFjHSB+ljO4YoWgxnNPKRXkIgPMn
TOUS9MU3sX3ZkI3XDOdCd/C1np864+WjjOoIZSfJiC/A5UbH9eATRKz2VJn/A6Hy
b6pLrbEOF0MCJiSDWyQEBin0JG2QCW8VXmbs9H35nldPu7rUVLFHBQnvEJGTMYM+
aq4Zx8Tj2VlFGQbEDI4cMdjXApvfrUS2IE9kKUkqcdrrbiFuDpvYtMu2kjU4WO+v
q+syMCfWo4HnDv/skpIBkDfPJhl3nk5i0whRvjaXvzkpvALerCI6WCZ3MmClPGcl
84m4f3biFgRNYJQtxG1WNFcPdEwWUE2YgZFZNpqTecMWGeInw9ub0oK3SbHgj9XT
LUSMdCzx6MILovRzwwLW9UsvAtWcNhZUG/5TG0K1pFttPBoau+vQVnLruh7CFgCF
5WK5SDYl96GtNnVuk05zXOwwa9G9MurplLfswvDOtpokLTRyaUZogyGHWsmYBAa1
7wjRlSvoQl1Aa+CMBpn2qL/ILKnNYYnl+QrtxqQ/Iy4YfeIqBpmnd60jIyHgqS4I
ieS5WMvkHuFeJ0MTjkh5AmWPqLlsDzzSmQy3XkAMDeyEW4KqtW0PPblsJmr1j7K7
0HEYKxtGe6waxgVvYw7JK+o8wwD33C0NWXo0+h4xJplgayWuPNZ+I+nSyAJMNTFb
ff0nBkmmLDwYU2680t54xM+t1jm2VHTPIHWuS/GPoZXC7la/2AEM+mM0v3RwkQuk
yMIACqDUr/Kw3pyW5cXZzoa+5Lt7e1TpU2dFei7y7i9th9hJqsD0hiQb3XdaEFYv
FhQ7yY/b+O1MZ+aoOn0k7qETlqi407El+BClskY7ktJGE1tHTufGINh8h4iLksic
r4/2BmAfsNVvliPeNJz88Ksg8DmNWIFW8zZ+Vh9hiscrB47KZal1ybuxaAGrhtr3
LFn1BenKokTxj+ENCrewA1lEE80+IvbaUfp+8MlbSRGUdI4ZIMTguEGf6Nbz//U+
ztTDjfh4agYKrpvQDE0thxKYTjb71zamrCtom5Q/u3FLdz+i+F3NWO1eqW5sEkn+
IU9ibGPwzZiw5rsvX/6ZpK07kiVMjuLWfWrIyTVwc/af+MquFgKfqNTrEwD/ZWyJ
n8BYZnJVVQtOwWSfq0kMFvdmOIIOgZf5UMcNmqa1Cty/tSZ1bM6mxkeRGxlOUxJ0
WyMN8prGMX/cMKV0dOkpoceXNoLcnim82N8051O67UI+P76Z6FUmYzGSQe0+3tDF
njLEailBk76jKXCAdu7yRTBmC24+qV/K/NN2rccWvSOHfjFDEAQjnvVHnZ0wVnlw
6M8kVg2GeCiKc58z9VhGKw8Dajj2V921ywr2X2YKIbDX3wec1XW9Eb+0T2iNQiUO
HTlVcfKsCVoJeGw9TjpYoW7LWig0UxDmhWC0jmLTLtoeuRPISpeprcuhBoj3myeU
dSGm2Iuxfi/BH/+fvsGH/co9Jox/Z+9fjKHQ/iAVQxevDj9fkA0xf1so76SXIp37
T9fZuB31jX/er63+CH6BvNl+15A3kOVaos7rKBP5pRhl0XjYaKvKOQulCCWk9uKq
iVeUFuEdIi6YqGk0j4JiL//Lg28NfpauKJWkz+asqtIZaRbJYMVrKeK/uwMrZSUB
PhqmnkHrZ6fLlwtFv5cqkssP3t/372NE5BRus6H1fLbxooOSQHYu+WN6XxKgIDLI
xS/AJjY98pxXkE1hf6td1YDsBTilJRi1f/Nuz8cVPzrLKmOtI34USodvyR4x66b3
FwAAV8kcPLGw4jpkvpmMn0s4S0YhuLDCRlHO1bAjdO1n9KzvA3RR2WmpkchbEnAk
/9gs6QSACG2ZnRDgHBq7q31zOne05Xa36dYcepzZ/dGFfvwexmjFlb5V2IFNMYye
ByUUQW0GkK8rYLUauu3yC8MraIoGWXYU+tEod4Js3mAI/y21qpqximwsNEhtcAv9
bf7V3A9gXJuRB662Y3OZWJNo74dIDJ7H/5hrdY3c+9Gm3YVog+pFWzB4pkrpwluB
BQgGyHkAaDebsl+kwdXzHl5oQlM2oUJn6vvkUL/Dx/s07GbmgnpPod4JgJR2OTH3
NDvJnSbZch2seqj1msRWO/LuAaYUB4vhOr6wTxbavnIGXNquvrJ+jOXuW6LpSNsP
nfKKfOtehfJUf3AFE5qb2OKFtL0WryfadruS0YYuKbi0ghwA8WyEnY0zP9gtokVk
/g0uvg34DY4j9BuIKrGU4P3MTUgfsegaWLVZt2Pv+r8t4qxYuwe1gqUa0OqFUaij
GULivGjnF3nH/wjYLoszDvKi/gJzsyXm/6v60QmKZniJfHxfO017KIpjFKw5tX3G
0puh+5PDV7yp9WWW0oOoGxxHmVqSgpVDZROYf8rGNI+R7UWnTbhWBRIh5BbVr+L+
0JOReto1LEePYDEFgDIkZrv7SmQoSSjuFs7QxqCY2RTr4cQciLbBER1Bt9xI7Cte
qEZiOaxyGhyBYoNnyYSXda8Ei1DRz+i9KxMlJqy97sDKulx4Rh8I5EI1N+Acb+h5
zsdf3Nac2lQY2e3U3A71JsqFDTAFjWX963A7/rjxalHww2v37igJRyuugozhjdg6
qmV0QIVGcGGE0yiut6+8e9Y6HTHfbWe5/Ft6fIftfKD475fyS9xqXpHC6kcgQPMW
I09puMyF8byslUgVjaoo1Nkr7X7vRe5t8MwS5mQpYDEo0+8JbvWDvo9vv++Owgd1
micdHEH7PgHnDkey+dq2zYRlq+nqV0dVDxUy51o1Wu0QOPBhKUK6OF66/hM+d9+n
xCRv67tumuZIZOPJ2CkrBtcCDo5wqF03saVUrj2s/0hJL0bEeUbbntgGIPUvlTw9
5OQazV3hz67L3Doy23H2/rVXcrhCMSa3Nqn918x3jz2z5Qeer/iaWJaOLyYImv5t
z+SXcvGfMBplZ4tliAV+jKgb+XORD1KLhXC3L7MFS+uTXqNb6zszsNZA3KZh5msE
Iae/vbe/4UBkaPqo2Zb8IV9JBF06dA4JXUYuURF82SIBc37hdmEX9tZevNZFqKQD
P6LXZyna4CXIgj27WqoLnPmr8/prqBR8EP+5VFpdLL5JWtmpPd8WL62MJCKc3Sor
g890ArHZNsFLVG0fOHC8RuUmBCW9f2C9fz7Yyy9SKREBGGv3vPNfXMMN1Qzu2Fmm
zxuMKrIawAlhXnsfRfEY3g==
`protect END_PROTECTED
