`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
op2adiSZPlNSed4/RhmvYPunJHMe6fNVyEUAEhrtjT2rrGyoA9E2bvQor114v48R
wfHJ5aXcedueOKd+sQfak/S1giOBnhHt35/cg8JVBpj2+CJepYTBxZ0vAONWk65q
8lrrQjRu2pRxoX8uzfyoXEuias0y7A+787TZs9PXFD0SxtuSPeQSZ3mmEJtzIrA3
iZYGx27kI+P7EsQUowOGXGmJQKVHWZoZTpPhAGQQVyA=
`protect END_PROTECTED
