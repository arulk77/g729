`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMIkC59IPNUxkDYyv6Q/cbktijZ/y41F5L6VM/M5P1qw
nKGsxoZZD3acrE30wR0ZOex7evrff2PWu4dRiSUEw7pF4vo0mYhsP7V3uE1U7Jko
sMCW1o6/8zdDPFGhd+hzu84u3FPSv3YO9B5fBo8fFvgFlQk7x4T4A73+7fsbwFcM
nMjr0Wcx8phxGwib925nUEgntJVYLW7KAyegXjfD4biD1v8EMp+MjZlpT6Bp4QX4
kCAL5i9LzqtUMrPdR6Xpf3eSyyZI98NY6tmcQZ7Q5zuRnmvf8aYHelYAcGDmshOX
vKcwhh9szRCpz0UUxyoX2tKo6pyRPVjT8T4nrlGc6QkwLhVEJQrAJy52OKDGaqhO
aM6th35S7wGXmJmZEdUqR8Q0wssbduy3M5MmPuQYTibe0dX+OYv85dAJ2pdC/FP6
dZPm4FyYAXXkYZFgRHFYk3ZaBcrzSy17cVpfqsDsme0dn8GyEki9qEbz1zwcpM7F
UFZje9NRrEEqX7EuoKuyE5kNpmIiq72KrfdPEap1ISwB/zzjNUzrgXPYY4kvaf34
XFbXZ6VeuxX5tykdLF97ZltIuGn7jrTYdSKeB5rqkrVL0r2K0i9ScZgSOstTv7c6
QbSEIm6ZSGC8/+X16v6fiDYuXbmsiQLlq8RyvCOuhv2ml2wmUZHckvNkBxEBKQMS
Jdq+VK20ZWFdzxmPmnjbMAXQII3fw7Xyfmp74mWE2I1zDbSGQQ+UJgW2FRwCZSBP
B56msMGRfGEOExtp/UyUfj1+4qZMLyMsA/xomuuE9BzdZyDTmH2w7PxgBGMNJHbw
mUynSmk5EaojE+7M3Hcb5bg9wx6htLTm+znpPxd7TxDqJDxNjLL246wFmr3yM1SM
iCWd/XRI95fJdHwZbw6IwFYLQ7nH3Vz8lcq+9erdaP5+/XM5Yva2OBvIBa9XpBg3
7VNT+LtGPu+rtJ9EIk7cA3cKZDiIQQGR0Z6hvCnrLlrsnth8lDSxktgJi3aBq19R
/W6Wnw9hIJcaqthNWQQfmfsW+q6iVT5KF90UXqVhOvu17oA7QFhjBJ1FbS6VF5Ar
TqhE/NWhoVxQDI6NAQ1alnazgBBiz3O2GIYP6yRYrqKdIv4PR8GGhf5tfLvu0CXA
1VXxxW89wXore9o4aSnLvDOOytpqS0hR9QEjWkMqBFBIKMARJiLA0rW9FgYj19wZ
7+iMbYgsnj4CJw6kf7sap4B+YKa/28gbl9eUckmsrK7b46l1gLxV4MS3jUxX3P2I
UCLcFc9Fd0DhV6ZuqISxbXibq8YVAWDIlkbntVq1X7rL/cw+8Tg3zM4sxgP+ystR
nwLOhNFCK0UzOPaSgtCkQB/Hpc0C55CvON+xTb9jfiufWfTstFgtfavXDCIzG2ja
lQ1GRH3fpgFTQKwOGfBU/+XQezAJFNfWKAIdZwaKIQ5IMOxb96asSm+XsAdXY3Gq
1Y2YHau4H7lZ0drlZT9j94i38/hp6LDPUMKGJhTRHAfqx337Se8T3odLX6YY4y4t
gn/Ecy3UBb4aHOIugZul6wZw8E5QAPTfmB8WSXLGZX941yrPRYj088QJ7/mbN8bW
2ekETeKMfsn2sGelR+7pnhMn6mq7gb6obHRz13H0nurxaPCA3SyvkP5XIrwxa4Va
T7e178zcfn6iKBATT+De5Phbi+UuZ6fCfzr4kqgFZaCkePRAPvGGKDdwmlvjs9C4
L3naWiT5LdaPTXpqdDYsaDoH+7ihsCw5ODnwrEMMmJBP+JvCpX2KfwGDKe4oCzID
vS+m7SedSkT9BXpNumgmnobY8BN5Sgwx6aXGvwqj4lc6vFP9QJ/eah7Uq5QEHyim
09mwc5UyXQv8cpw1FVauj07OChmT1eaa2gTy24oCWomm9oyw4qmtpbM5h1p3C11n
8/qrg2ddn1H15rRHu2H8RA1EOaCQfpqd+dS6JIWlCp8V2zVmuGaMD2DuF+ArumH3
6r2xvZ2RV+cireYYB/h+f283zoZ+u4K8gN06kUHOf8E=
`protect END_PROTECTED
