`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
8wXvl0ibpO3hleMxz5gct8+fI7Ip4EUVaamWbtpewOgV6U+ap7COj/1+cKN8G0U4
nWz/azONRdNMzOsPSQyAFda5OYdLObgUo9Zu2VBpnbZ45wbgem/PzzDZedXlMg4E
XoSIMQ//SEzDMRr2fnLZ0g7K+DU6io0u/50r7aSqNPOh8IcYtaKA76m3oEQT/YyB
LofOvBY1ao0fWAW+QGxebSZmpLA4j3VGquyUQIKgZjXq/0XqlYXUPIXeo0HO0FUX
sAvt5I9ynC1RdFJIuiwMtIwAqFNyh5CmDklqM3mFxH2mGTDUMvZlKYOgyHzg1rdA
oubIvSYUAiGukDHUXov527ighAI/rSx0ojh5p6CBCsOyGXsLhro+YCbxQC1bOBX2
h+ogKvEiR6OiZylq2RrBGvMvnJgXDnu5LsxGfDKplGji2tcRl1E9Xf3bt5Bn2zT2
oT8KTpgVe/wpg6CIJXiRkbzF9G6dcPYIIkJ8XVgc+Dl1vr4dmqBDlPZ+o4VSHvjA
ZvbPh/sAQknyYKKMNHq15I/cn9+D0pftpVCf2Xk6crDeAGp80ltuty2ai/bbN+93
GSFJcEEwzBQV08MOq/VK9JG3LdMewHJLlYQ2MrJZIYIth3z2IcYa14y3uSKM6Gun
IwgDhbVC2oluk0zZQFmUju+YkKjyrSYYoHOkAjwWjZhMsRRVzMdPIZvi/me+m9V1
DSRL4VtUPTQunKYnDjrJoY3CRfLn99oP5eNaxp4Nca3La7kCH2O7zo9p4H2knl94
21KvdQ1PrGp0VVuyGVZaTtcOeTjfdxDmn6R2dQxDfVG46DtCp//KZcD5CKoac2Dl
qhu7lxvGgA5V5qxVwLeBKMxUG/cpeUiJipARWN8VARefQNC1/Jcw6jJLt1hQa3zL
y7MoJSAH5wHG6VdcIWgtXDsfT+P/kQdii+QDLUB3ybOiP/J0c3Eur9ICMxru/0mX
hsnBGn+TJAAioCO0SujRPC+Erb1yTjwqWysEa4wnIUm9i32TX0uQc8PI+GMjcl0w
4mHURElovgC+nYOI+fGcMNBDT/wlp7WkHC49RT761mgtSXbtwnPHjR5KsdO7fxSE
lQ6crzzBm/smI2nFz0yPFMyObQBK1avdFpU8ah+mHakcndwFQHkUvHLZUJiOB7XL
CGGrgxIKKoG7i7xXhJ57YZT4Wezq8dJEpSz7WRB0zoutTLACjFYitxseTl2R8agt
PnilfoT+3c9t9Sk8GyeSEcgbL/on4QRhs/ZKY1shr6y9tF+sC/G4VWHCyxZl+ZwY
XKn66e2dJRd9RKtETWkVcxGOilDnxMumWLvl48HKYcCU8p7zdch6LUBoQMdewFy1
XtOz1G1KfxkqAUL8ZUrB8SRDDMq8zdNKtEDbqO2LXEc+s++W4rUuPF3ns3hjlG9e
X8VYOUMQ+UmtcY6n1GneYgB1z5G2t8DvaIC3gGGkyqce/cG/tyjJvlQ4NOmS+Wvk
9C6UsV2Pr99YqLVhpw5UhmoRxXgDSoZStD+Jre+cauocH1VX2x4ikDM0kmAiA61m
JmosfeKOtDEb8G1erIlwalYVYAEyF6NtESUQasNmwsxt5qtoURoxaIHKZ87HCpP7
2nVv32nBOfBnDllVd75fxDah9ryw77lTCeXJUbmIPO7t2fiiBBOHAtqGTGe3/6Mq
Im943IU2T7NC9fcSnZgv9QtJLwjjjf+mTHLkiDm08agk0X9sNbaiBVVUCmiX8U5W
OZoHgS2PkH4dHT+ul2MQK0pY8rzpr/qWWFHgDMSzFubopoZERV+mdIEhidUHzl6e
8gA1e4xLW8oF9QxHduivSVidLD1Z207bsWhyekv41VgfLSn2cTIebYLnUGfyrJC0
fgNwkzg22GBrlij7N2sjKeYJCE1YkkkUxTYS2vTS7xqaTXksEzJQiQuzfFRU6JOX
G7+0JgfjW370uykWZPU2CtPxdFOTvxew3enFKTCSalPJ+cjZsmA5OvxOJ/ZOph0I
pOFLxjvQVtVSW5H0bUE3pWlZv2I9dPcfFlWiLYszoHkzg22SQ/M0vn281CckvIKz
GmHKi6Jm33to5HUCbTbMyBu6wJCwZqPptiT7peKCqeDcSFtOSVcAvn0XQRLP/vhh
IvuQHtC7eClL40968i/KQcl50ZVk4r35srMNByQ0rufTePzKVDTa0F8nplbRFS1H
KCTR2CTJP3qiauQ1DD82XKbrLAqqiNA/RzSxR3+1ozgZAGzJL1He39giguTh5ngi
75NtBYKMyAQls2GjekMeeEa1cz1317qGFbf5f9E5L/zfoXUMR3qH3uMyT6b20rFU
uM8aEE+fgDn/rgUwQsiPiA==
`protect END_PROTECTED
