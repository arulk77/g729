`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
MmhIDXWqqQoq2EUOcLIUCpBX2Fo1Pk8tCYhiigwUiihSht3h5ZMeZ8zl00JS3Mp6
JiiLjjwRSFxmyIX6KkAft0b0jhqD4fvL7UjJ+aVs4RqG2GDMtquUpmF8Zy75+S7y
kSRjGHcxH84kFLb3wao/WoXInMY3Im63DLuAQwkWpnu/CtdhHYAtv7S0n4dKtcFf
rIXtW9ZF2gigAT3PaymVLo4ffQCZyovysB7rHTovO70VpBKg+qyi3twjpCuuhy3f
vLTUYkYBJ8mN0iKfay5GXe3WCdX6ZIgo+M2tCwQj2fc=
`protect END_PROTECTED
