`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDY1RR0sAl6zkwtZcP+1KPRoYKQgeZNlBRONgz4zA5S7
kKS9TOSEKxuEWaUOV2FRV3wi7H4ZHYJrM3NCqTi4+hOptp3G+e+wUwI6Auiyt8LL
Z2g8w7KC95w87a84tj0Qcraa7eDnwLX3bZXKgOdTRQ4fBz9fRvZ4Z77u0tqwyihT
Xcdd6FhNsBwKlKx5BxxTYS4MdsktWbZOR7c1/hd4bgeml0O1LyjpnP7dqPCQA30U
LVb+kr7H/1qg6EfUVz8EEZxTm0jFromsfGwmjDDZTcSB0VEcJQ4YPkxWvpgeVzdm
`protect END_PROTECTED
