`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveING6pv5vaywY246Wk4Lv92tzway05gFs6pHmqxfvYf4
elq01x6+25w3xXmxbVK0t37bu2yew+/Up0bqvEDo0u6OamKmx48/SqcNfjElaVYY
OpC9HBNGCIZsJ5O8on0mb5sY4T4kN7488IxxYXkIgLRCmcTG/dGWQF+gOEiPIyAg
DkMxgxuGU8cEd5cbC6gM1A==
`protect END_PROTECTED
