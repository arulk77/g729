`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aVX6tf66fX0QY3dxz+GdM58nXTGfe5nDDHzA+o6R6aqT
n2U/obTE+IPlC/rIjjNE41aBxQscHZrJPjf9HNLuEoeQDEOPjL0TRhgEzriL1U2F
XmnPq/R9aSRjazJKHg+OnhqwCIArHJU9t4SfIwFKkIyuencpgBHajhEyMBUf6Xet
ygz5f6BcMQ4ne+nZkjFwU0rTsI2fKC4Zdsjd68TxPan8ZX602sHjf+91ZlwwopTe
op41UqYKouYGDYMKV9zo0Eyj6MZiddrk6aQvBdqIvX9qq2ofMdopZyJALP5a3OjQ
NRzU70Tnl9bh+MssTlA+NICWVIS8jPjBYmygsuEoGK26c2fE9oeMLAUkuvIspXPC
JaFX1a17dCE/M4B15RLyfcb4G+yWL3pFNln8YTsRD2V9dOiE1hcQ0gWoM1u97eBx
qlNe9+ElcIjvxHeikxQh1NAp6j71nuKfNY2CwWq/WmpWqtUbNkQIH1cRKEEu/EVO
1gjopBbTCAiBhy7UAMXmeNl6CM69As0wtgjGgzJ1ZVRxFl4d/HKvWgojizPKQP6W
vScIDHrvF2hLT5hDnm3wW9lmuGhg1Glsx3pfkVntQEZ1YpGX9DjEcoNG2cKh2wr5
XLoDceRBbgYZCPw2/xcPBWkqiogLDtoAhpXfixYMVmSyYIstW88UVAjPId5FxnIb
o7s6y/nv5hDWNu4Ej6qDtWUee625yNoZK8KjXZr++870bYqV13VE8psQTH1NlEAB
ziNi5eT4YQ+q194WQKDw/Cso/37VlopXeSCfpzU7LFwzxx+WRsch800AQHlptsDb
sMSZroAEQLAKJGjp4bXQ/1VXlbjmn1NBdOja7ftbqSx3FsSeTRZFeDDGhJYPSHHw
4awobv2vrw16jlr7yJoNsVKxP2ye7W5DVrplmJxcHTtA7Lw9mED8xDYRbzXl1pO0
CMtwZ/4mHnAAs4CUCUWToHWERgRy2RK/U02JZcjjUEnj4vUtZiXAFo4ZTrfpxi+s
6HTZp6GeY5dnlUc4Zcxp0DcwfyOrMkrgA6jsbo9ybI8evQE0lCqY6UlsnwLb1/ji
maoCO8/OA8vLs652AsWdHQQn7MRyBejVcCS3Ec/M8rA+0pcKwOdNy6A5aSSGxf9q
zv5Aw8YCW5SGv923lMOD+qMOJntTKXy6i9tofPuqCHCAm/toAa8LcTUoG4V2UGkE
BIscITYh4ZQYEVPF5K1308RCEVJcD5JeVAGP46kqtloXHuhaw8MbJTeBGe1Pgo33
qLQkFpqSrdnTq1rpbORzBDdpIWVl3fkmeut0HGM/9Ut+V5j/H8e+VwKPMYhZdemw
WnWwMaaFN6lNY1JGWiuxY5iiZDU0Z2hyGTPVY4nZYgHdQGDiHme+tNxRT4WOApyJ
4SVnhnvxEANlAuX8v+b0TE+TnXXRhvbePqywomuvh2gIwqobkLHJQrZ6IlkSY3+g
XYFTicF4zUyDM2d7XPyfzaXLhsMIN1skYyLZ86hZidq/ijzM8z3D9ob6kxOceIcd
1zgmJKfLri8ASvP9VdajHQdLQj5OkLzpYVfnEX6W53LQ1BlBvtTNCKWYUKLCmrDS
SFvbFEgwCirW3G1FmwCuCiAYSgaggJjLVHWZcZ5UlGCCajdk/s7Q6ky722T1uu+n
ROLmiIkP7J7ofZX3HTM2JEveyURhjzbHb1i09oRQawzMPwGDNiVKZoXfozlBI4Z7
zOOanns1fF4zXFQ92CtpvCKAG6HsOGW6kzJdqQc2olJsbQuzrGIB60x6g3l45ZSe
UqLa1IbGGJCX8qV4UnyA/r7teHfI04ck1dSlGoxDC+Ns3IN6768E++Oo56AxnAnx
dtMTTFYxBsISY4mDC0nd1oDwCEuYqe2bwkG/OIcfZUxpE+sR37nYfp5HJwYSp5p9
UzuoBJY1RCd9q+R1BW1cdb8zl2ICdYLS18KXPasd9zl6fG6ArY00FNp5cIj/Y58E
5Zp1mi3d/YDOCdbqT1vq6c5bOSSPY2KT2dcacgksrRmbwggoz6F7VK9c1to3ggxk
Ul/bXxf6IV8WYduhrvl97WoyFzNqd4qHNvJz6xgXX4mIQHfwvnDm/nejGFacjBW3
`protect END_PROTECTED
