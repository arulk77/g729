`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveANPlPuNEeajJODTvIBJhzt14alRLC8dBQXsdNG/igci
AarrhG6lRVAvnk4fBZHqDdccf+i9/OnqhuOCRGlDgNyabNC6zNF/BDA2Ekosi/Sp
DYaHzDh4vi4WTqSqKjVdnlRL+8sSIId0MlZFzrRDep5pduStcJkT0Ok4EVJac7Mu
pcv04hJ4qzYOPPziX+fzG8Pa7h/5jlE0CTTy7l22WS0iO+jQ8efAUmsJoXEw11jS
mAPYn4kZyO2O2uGeGky2znbiKfjmBC6nfVgCwjH85eG8uftQ8YE/HsHJ1MyMiabe
ku0eIIWDcfr+cc8m4ZCNfPgudKX/MicKr4oTmgYkfgs+d5YGC4CF85Ujnqwjx/gN
08wcthvPdMIL1uZc6NblkT7M0y6hYsLRMx0trKEUg8/McKBx5QCss25E9w5GuXy7
0b7ZlM/ipCUVVzw8rWWEFJ1K62ANB/hC9+oY22sbXXcjzp+iwQedi3hVT2Ygb1mX
28BHSHa4MaOMjvdcAXMP3R5yDzVuHlbjPoHqBQeSrnjRZcdLkml+dMch2GYE4xuT
bXbVNBcjDK6OWk4GVX6erFCjyg/Ehv7iGvzOLMd4a3vqi4DTcTjvHHH/GLvH0+VE
fvu0Zf8fkz+GruajCSaX7AjUsq0Gw8ygs+V45icAhnwEK+FCZK1eH7Pcdiw4niGW
uVhTKLIfWltIGK9zVb8KEgoJctaxdpwAlpz6urdbjH8G+Gqkyn5OASjLv+FgO5z3
IkkDkYnjHw3SVksbkI46zW4w/1wE8NpkX31SuEvEsAfRDImPdzbnTqLhXMF7P4lB
OY69FAPe8T1KDK0/jefaQ0cKIuudOqKKWnu2jycXZKA+1rXv8R8EbCKXXTlrQSCx
kaNACuDlmlFRDBZjTVxuSSmF5kGCDCi3PTXnHs0+R4hbCX3pryBhn/0XJwuU+eGL
hYqk20zkoe6hWTB3LnJvONAEBvMn4rmq/kcXcskk75JJkMVOCsWeuEcL/VUuekpm
cFsYwTs71o3e5wd3hkBY5RKYax1nsz63zQmnVpqfM6y/wFlHgBJZuo7F0xEzcrc2
7qbKrVhnYUBS2GTDcYrzddWvRyWEQvoTZxmDg89dXpZVLZF8l2B2NTFaza/xBL0E
7kCo8COSF/3IE4o9J7j5aBLOMtyB+hUt0Voe6zMI2I/4NcqCS+XfQPWAhBl7Z8tx
UTlRQ9rS871xA5fEDgARVku/H2Ti4C2NBa8Yo5s75kybQsw3Bul/WJXjC64HnTiW
FMA6n9baq2Ltihe57XYdu77Z89PJzdnfNM2SC+Z++pJZlY3cEig6xVvPz9hKvDRa
ho/84xc024wu3xPI4ch26ojbIhsFb3WAxq7dvXijiwKPjPYR92fNocYjUkF/P6k6
6Z2/HjYelV2vXgkgBivAIwDH0qPwLJU43qP+bzYbmpk57Nyi0+4ChNvVsOHBomOh
F1ElrGr+rMPyEoEgDa1cIewtbWRHeF7RdxPK3/mapbsPMWlUJdzfxc7+tzS/dxcO
8CCBKneqgGRpn8+7j6kxoXDfkDHmpojplPQilPf5mU/54BK+2Q8jGor4QPu/CuR+
r700ahaicCPc6BUU+1phpN2V/LrCTB1tUK0PHuoWPDh61UFSfkn0pw3D/mkxQTlw
Gv63ijw+2Kag+j+1E3qxlqZpz2oA12TGZIu5pg2DEIqL0qe3k7NO6jh0b/6+eYMA
sJnpAcFNHyNxIAAtc6JNLgLUKb74YOA/1IMSWV8wd5aFRLeq+2UEm+97jCI0Q9I2
8Njz7pYGFvP3OV2wAxDmUFmFzfNvAHY/VJP6mAp+N9ZklgvDiCXn44JQCN/QUF9O
0lj111ArlI+FoXmbppNmKm0KNBoMu7NmouXQTBdFT6gg9XWVWbLCoHV0pT+zeb1S
tmwQ8j7TtnGe6QtW4fJCJE2uXwxTU92ELIzZzmzP3zlPYx0aeAAEwl299ooRxgFd
5JVHhTsE4Tz68vJsPcQrh4YtBU49+hZymx9VfqPXZ3zKAhuHNvX0iyz8BlUTuScy
JiKodyAv07w7DolSj0d4hhBqIQ/Sr5e/XI0ZkLlc0l4qzMVIR3VVWgvpzE/dgUUS
4p0x5aRSDpP1b2tMU8LINRsZyEOePnJaGf/dDUMr+bNXco8IQMjhj0PpB7OU76yG
4F9/jFYU+5VzgVyMigK39/szji/CL9fnnAZ0X39zpREuCoLkTmJZTfvi9D96roI1
5hLaNRADFewGKrAWuefA3Q/Ur+9ig+G1SsACYI6nMNzQQnpSssuuB48KBRAhFYFt
ZpcI6NMDhZYG2fZd7izKqzje9RFWoCyyVCsYi74s0Ejos/y5dCnwfvOzV+TtTyoP
6D9DccDHiieF8tMpQUdMvcZW4GX7zD3mNlr8kxT81mjssE0LhiOFKlM8LcaVnh2X
hfDfPKsFALGoUyweWGetbqW32lHePHGl/zkZflZXXsSGQAhkjmUAh4Yu8gLw9cDL
cpyfxtcX5CALkjaP+nz69zcWgi22yY/5/hcp0bsdCW+73Xhw1CP7G4o6Fm1D/2I0
oTp/ihTZAjR1FZ3MID4tAn9OXx75T5e9yPMbJwT0EgywqDA6x2zw5m6D7+B4rSSp
mvwF0KHa2+I3QlcrV/Jzn0/uilFPxuKmTOIpjf4VL7cnVJYUbbCRfndEbeG1oSxL
enJu5U+FZS2Wt0mvup6HiO9aBtvXlaaUzPJtqPT7RajozaImsCKWObOhniiP+R4h
AXMb0Qh7nCeR2GVF+V4dK6CYobAdyxL1TCJZRmM2ecKG33IdFVAN6DaXHKEURo6l
2EFxfyLOw+wOaQzGy2c4+/IKOD51TyQxIdZ7e87i0OHMCvw5Q8tmPjz+BW75fH3R
OiYRumnacwRXeaegSzELSV7WOUWlxLuU+T6NroLevfg=
`protect END_PROTECTED
