`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4xGwf27VsMi75wKkonqC78DWA5oUeyMqqpnLY8f6or1U
AqKxJBq8NcHug0Kd03dy0JV6CCfoeOHe3XxfvKxsVbUdU1+QBIwp8gXE+cEJdtVB
31uvk4KnSoSucBW2133XAUEr6MAvOpwiVvR7OOQn4qo/nP6QMSlSMFT500pkCoLS
CTXd3Y1jTsgKx7Q3BAjzYRqCFfSAQ9EBjPs/31jaFY9FmIOmDMKmY+dUd76sA0+w
e65LkdwyfSL4wYUur3CafP3ihE4ta7PZcmvfImYQv/vh6fERBMmHFfK4LeQTAb0+
HFSn6tpVdjULmY7UtG5bLhqGkQSdU3+EjdXO9tq0SHDqVoxC3OB+E4UdeDYdsFOM
gsLaD50hjolWW15jUiJjciW+re2AjH2QPqm6cKyYIVPblN54e5FBREdoBoWs1tmt
6wd8MvTk1UAyigBFl8q2WpbViC76+LmiYtalmKE0nN2rDtjFJ78wlaL45aaOB/HS
y9FA7cT19iFHdMAyM+brfVbmQsk0RLDcpBA/WYKsL+4W13XXRkkJcoIqfAZ+GG2p
utF83cDkAgBE4FQPj+1ScA7RAFuOwzo4OUuGQoGbrDtpoDtis1FCRYTQvwUQxKNv
NItteounE9nKLDMZLOEeNr5hRYUHSwmSMfR0WjMKp10oEEA5O7V8bpoYk9MI4jT9
847ijo//Xodgb5NeSLY/7CK07wJnpiZKj/HOP4vruwVtX7u46Ka8vywtFERAuS6L
GgDBhvlg79DhOFkc2UadLf2JK0EwIKl8y98dgHkxBSA2NJONaL46FqhbyvB/GWZD
FZwX0iLIbTlK3pIfdZr39U4CoDP8S1WP1KpRFjRZkghhEf0zW+hvy15IBai9l+Y4
h2gNBWdg6s2t7RRyiaqwrGiAQTw0tFUSj2DTmJG73o5KqHgfUSUV8YTo9edW/dKl
4kkYQ3kkUt43QSwf++Uv/RksvJwvqoxqi/GLJ46YigFlWP8xsjPOcyZEJI+GU7Wd
F3qwbwshnuTzKdSih76Fc1eCPIoq5YFBgNTB4oWUqagwKo2Ztc3YTBC0/h/9qt9y
nqZDs54id5m1EKsFtnN/uR3BTFKxmzHjuLO3hVJeOJhw7vYg7LwxO1UYHxdjZ0UQ
LIBBdLo2AT5zKTeeYthrdN6OBWJOiEVf7tgW3dFF8J7P0IaZGJH4/cH1tIHHedAO
tZvNtjGVDB3Rge96FQRtLzxt7ZWPaUtTNWRcRviHN2dJWOaJUxQgHQxGRm3aHv04
8dpWoN3A0YM4mDYT6QHTxiFMA1dVmrxnJRJJGrI1IcRwUrgo/YSNNJUb1f6Z2T0d
pS0VeqOT9VLzYmX/rqsFAWg8GlizDjqsCld7Nmz76m7D8Jrw7cbadpSXr74ZyA93
feemwbs72Titcl/dj62fYgY0SNur3QBDq+9DDA9UAU2+Ui9N1heLLM57KAFBPm2s
tB1nS2/2G8oMMm8T4anAqsMXL7mxEzrY1sJxifUaFWqwrYwXF5pVW+J9fWjvtiST
S7eHCQ8oe5pedDtwe1xVGWP7eFmJqNpuILGPZVV0YMKqjoV9oidQObBBVh4vW6Hn
rI7b5+ZyNSmoV4he1PUMXjT1SyU/DIOu2IjyoNzSDvc+aIzGHItHhocx7IM1rF81
Y3DsQsmrzlJKo6mbtbgVIe3Ym/4uN8IlowsJp3DQUaaD2hp23+9BxAXut3s09yTj
MgGMlqV67r1ndC0XsqnmL5brJ8AOMXNZ0FJr51bjNg2mRgL/6JQlne5gyjIUGvxt
ZahJ//LxnNezdFVlGpsDi5eT3+bBNl3mrsair4l698A1ltLxn7/g9t/8ydsTYGh9
KTsoay6XFincrX6qV+vwP++Yy4gBZV+mpmTjuZqDgtZ0HoJnImWPrvWK3acnDzBx
haDbZd52hm5RUywR8s51/vRoLXOAlXOpT9x8MpJOznhKVN91YzyRQQYF55Hqwc2h
4ED8dVISvLXhRvuYF20GRetCmMCtiQA3ShWzThEUK3moPzK4drRfqJ1q/sy1YZqx
PYGdcW+JYZLkA4wdsMnOgg==
`protect END_PROTECTED
