`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
4jUYkdt5VjR8oFbu7ZiLkvae3FokBcbOVstFyhovO7MMuGXSJBwndPuipwi2t5vf
j6FYaFnjh2jgG4RSN8eQRvRpl7/rU9WowGFH4pbWBxAUxNptnkWuD+G56nBJTWnb
ZN975rWn7cDxENoxI7QFHWkh9VzzjuJQ6SBjZhq6lxmrmF4D3lZi5RmhbaqWPLQ5
fskgZlOKn7nQ5A5CI4xdXTBnxYh5GwpD+kfQ4Us+fJZtrtXNlX3DZEqrayYVZP06
`protect END_PROTECTED
