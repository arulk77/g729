`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGHk/fEA2917jv9d6365iX9IwEqbe4dpm5u/OIMDNfuT
iJ1IHkr+WrKF6MnKfe+Z6JdrJhDpxqAvNRyb/8hQtESgfnnlpEFlAGVJe5jTrS/G
gtA6LPc+DPbTpQivZ1CEYBkuEVb9H2bui268+XmBYguL0AvJ8WwCWdoyoN/+fzds
Tb4rGU6nQs4jOsACXS6oOmiI+PmTZQGEV0ak7HvZ4iwOHR3Jd9r2nkX6B0KXv4ib
W5lhOgS48H8wwAM1AWxp2+QbopDMyKtIfkQfzzpT0M1W194MkPFeBuXsJpCyReH0
LzO0AOzbjfNHLOj82A2jPxcLY/WoUsMs0enptIX9p8bgB/h4n46eYzgqJnNIPWIO
wmiBWGDTR7pOwx0OgBTX8TMLoqM+hmzyO7fzznA0TpRB+EfGMBUdBlU7bmjZuFCQ
SJ7ey4UpucVwdi8hP7ejq0rYZC36g/tRIpQ+PsMqHUH4NCqJxHYuveXeQNKjrHIJ
g3kX5ONr6TMN7weHjbXg3zekdpSB1XgPhY+YqKKh2esMBwQErrSikjm8vaqNQY2c
`protect END_PROTECTED
