`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLwcuOd6DMAakujVbb/1cT+9ZYosv6Kli6ZeCoQDsUJl
yDl/UVKAaCJ5aaa1ptmIgK6MgTsGihSwzZa5FXc4lhVnY4N9UJdzUcpKp/G4Mbl3
NFZvMrEteAV/6B2ZCYcxLXKBTWMl4xzaELWrV0fVa7Ym6RczSQOBFX85VIoumuL0
+50M5sLQzZ3hq667wZbXj5xekGiYY38uSPXwnPaIpbXqp3prHoceGR1OFRZELp+l
adJwDpYAKanabZd6AaD8PFn4/XdeT3GvvrY39Y3djDjerXMqSPjQAYF96Ps6LS7C
qK1EyRIPPtBiRN7Wji3zPNtlTL4LOpeDC0zGU+2QdJblXvV5dmsZsDOlbFluffp2
WhbJDBtCS6Ui6y59KAuHwXOumkp+Q8Spou+PxlOUo5b5cQnowQYpNKMcPUU24kBR
gX9ka6bVqVn39nD9XqQEKvE64o+xpf+I+t55P/h7BXn9awmwtw6NE3r1iuVYyFxx
lZtQZeJ+G9PaPzOEHhEbtOqplDYIQpVeyUhg2WSCV/LCI0EnX0wEHaEzUzawdiHA
`protect END_PROTECTED
