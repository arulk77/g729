`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI16TdNKEXS9fTXvamx0so8FaYN6F4LM1+hHwkSOakuK
X7zFzg9e6Nlht6emxqh3Hq4gteT5gyQQ43YuTEJZI740cCLYS+r6TS2s9omw7uYc
QULRQXLf/AYgmKLxa/ZTROSEiWxwrgiOR0tLP6x1805MyxqHdeQxGvkPBkiq2dLo
k+yb8xBbk6apL5EoKPgA2hhaPeGUQGPUqXAgc5Syx+NFd+yRLamyZcL5QOC/I8UB
lbWV0tCYX5ooO+t1urajzIAcavLTq6fvX1o7TcbLRvs7xJO+igJdUASHU73YwjMO
r4JIUU3kHh1IoE9wFxcAUIuJwlZxHgaHEmhbbSseNrUq0cHT3rVZGPugT46OvNDA
G4JjZ6R7oLbpoLecQ8pLKgIuDwH1zHCPxZ5TeWGobXpAB5Bb/Ny51A5FKy+d22jW
7czBVXl1Dx0+GDxxFAzyLN5iMPe71dRGLO0u6/DA4zmtvx1i8qvmDUhigEGYa0J1
08ykfyP8LYNrR8Ud9CS8zcQuPl9f5lHd8WhVAhqASQWtpCz4Tb1AyCzSPpHnTpAd
4ZdmStMn7gLX3gmzCQWOu9iK9GzTs6oijXnub7+YzbEG0DBtfO8EQlm8c8180828
cgC+fSOyXCF20LPCZvIh+Pe9vyc4zB2t/Goz0T2zhQ74RFaP7ZwKT3qt+5zwVcHi
`protect END_PROTECTED
