`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKdbHFclNO+p8Un7Sy1w1Td/K565L3Rk7PoDpHabILTO
ZGWV6/pIQvrTLBgwiUXvSfT5yZHdfdd4DfRYSKJy/zSALK/Rhq8xNJu+e4u0b/Wt
UQXLojC3nI9c2C2/Q+sPn6XlRgJ0Z5FbNOVkniZBP7lCS/WZrApYtxBhsW3NkK48
TuezhBDzFmyAljn87Za87OU1/2KTTK72We56BQc2IsdmmlG9vNar7Wds70sb2sFV
Rl68BnNBVzfz2NCFT+YetjRmhyE4JbnHNYGb4d+tFaHwk8OpMjL4nt3FpJi47c7Y
FlEs3JEfskFpc6UKfiNDMM9zfNuhhr4LywfW8vRZDaaefvmg4/EjN3J9gWRxci/e
`protect END_PROTECTED
