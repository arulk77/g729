`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73CyIVJhsGjZEuZiD5jg+sydILKIgyLYY7P46SVdiOLVS8
2royinly5VxDU5Qu437JF1raSNW/2jb18qlXFnTHgeshv/JxwSdfEulakH2BBm+F
zTMQud8k6GC7j/e8CL/n6Hp8SI3VoNuhY+DbBLRMsAkyeew20GzGIMWaRGEyHc0D
iLZP6PkpY7xnhSKrNgW17fjtDcestnjWev3DnLPGp0XSosmfdyO0Kgu+1ordIg5e
LIDHBx8P/VQP7fUmxPM7vAuKUKJHTZc5HcjrLYq8aIfYx8M0XVqVbK8zPEzKoYFS
HNFKKucnBIYLAUJ+Dwmh1gifdfQnMhTG6FMiVmyDMnjHA6p+dybY+4PoWuSHlSvc
XWFr89RJ6ftsVEXpD1YxTWeD91yAWP9eDBJov9RR91kZPRFxzK+I1P8LUSH6LujR
x3PVcd8v/EnHjwubVVNSTWlfsyT76yqsfSLxbdh9VlQnxk8vFcNmyX/waJPgnrwt
xxqlyWr34DC46DcIfBVDn5eECjzvxDAtnp6SSOpy65sZ7fvy7k5IpWpi4tsch7NY
0WLgVhYOHB8j6plKDiHOuFn46mfGlvza05yprUtRG1LToZd10JqBjHonKZcIqabu
pdPZlK8XU54Ee7tK8/qLNJxtAvqH0hXj5YfNBV3kFdH80ItjFLSY0iT3LrLTAJLa
PNWhfB5LiukZdMgWt5Ef8dYRAGDcHiFz3Hlt7UefodT7T+LsLK3cUtJo3PvilWp0
z5gAtFIB3m82hBInmHTtE7kMxmV8IuHbZUURSRj4jnCZviFgmCMiLYk2nagHKOSS
HvubF1JX/OOiUrRCNjde3BMiFtnqqaPl0dD8uJ2ht/wpr5b1MAJ5fEymuHiOdlUx
G8gfas44m2FGA/DXz8jZ2aoSIS0NhPprrz5bGocmyuGzkMnJsTiHZQ3crwNmaRR+
1rZT50qm9NX8AKXoFP568EIzrq9w5ECtdh+jK9SngREEaOGZqS5avn42vOFxjoHG
gBQGgkQqUib0clu6ezuDHbPuss39IBpx6qzx0fsVVGV8XxgzGGpuNVK1/WAJz9oS
zlTalxd4DA9EPj04gQB71km7Mgkc9WyulXP6hS7musmdDyjWdCGQtFVyS/XyricO
3Ltcxm6te1Pmrz0xsk4j4Gs8O/2jfL+pAOXXm0b7IkttxuTEg4VeB4vWb/yRsNRe
T9EtneQpw8LDv/L/eMtCwlvHxCrK+jpwqugSdyIB0irN1Yf8trMp5ayMy9X3UbB+
MLE4HrcW85Bxf4SMf0MUiJFrPK4zVlEnXsZ9aHXYgd0snR8irf1fchhu/sGImx1U
pJ/GaDy87fvQLi22oVzrBQAVNlW4k49QAGC2i5orUH8k3/CtZEC6Tpl/v2EQizRm
bgXI82IK8tRFmDYOVjEmSNhtqaoab76EUxND4BI3BWUQytQmBU4XbjUjDbV0j795
DavmO2K9qIJHlV4ZJhN727+ONEOvJGmjAMr60rxmDOVvb1jDPrKiJS0usJ2RwQpp
AbZzLAGGteTgLPvFM/wmLLwZdmnFkLDJrdoID5a0LHlQH78iWCdH2u4iJw7iyIZX
bg87uTdBgzBvzU763FAIPmMrOdkk3isDGGYRhfzfFLlqiPJ6lNDbnZLC7xWOQsGF
jOJjJp99iyWN/isaJn8FNkA8llkh2dXIk9tFOqw7MggZ2mlW8GP8m16ALPtpGqiM
wHdbXCrMEAyZsuUvd4yBlgLSE6gQ5BwYz8CsU1Ggk5l2nS06/TokQxF/fBGvYV+q
tqNYikCOnMA4OEHBTCIkrJqsmA4jtjl1UuuNuTqaMCqCR4wWxYVm4ZeeYl5gvUuY
SC4/s5cmpQJ+BnVTr04jXMCxTSOuNyCmWLWVnWb1TzG4AjujgAc+EVlCXjPw14+s
Q+Y5BxavRwSnVLffGCbo+kJjOFz1ffvy3PttecIZXBjCsC3KeNvWDRFFUAwmQ+Y6
z7c4/0rOvdeDojOcVxzAZCrj1gOWpXKuS5NPztPgSsfwuADqhBsPT5eVXz82Q1Tc
SYCzWculeEArm9J06h0x+kxp96bjNoVj1zeIlRa2U29tm0ZWN7b5haYKVpxW4EgO
D9ZLQyu8erh2czUAvTpl3l2ONyjydSmsn/PSBzefVZQL0tqkrvaZ7i5d2N9+C34R
wM8GxRxNjim7g3vkNWLTYT+qK6/p6NS0dc0Taiyv+uUPxABIhw+1TGuCJTme3yhu
H1VwleDs8v8xMBXigdPuhKf/yM8VMaTBEP7fXehQj/DLGu6tzgwwjEXJCA4rf/Di
/SEc1XvqOBjk8Bj4I9kdyNpQQ30xdcaGBpFwREmLbVcv+FrgLSbyl0zNSCXQ7q62
AcBoa372a5PkdcHJVoRt3wtmAFs8l5PfBJMKS2OUeCTgLtCYePhS3tcpQpKHcEYl
ZxcKgS2GBhzE95Rv7mW/MIZwHC1OUM9Y4Q8xXZX2PNbML4m418j8EkBS7NDX3W1r
8JlgQ5hbhx1EDohJKiO22l4039AZImVJJkK0rBH5j+xFuwygM5B+00q5ooX3TQVG
Mk0mLCMQyDq5MI4OqD42ZelZi2uEYCZEOHWnJKB/lbTR5mWfoSo/m+ewM4TyVSrO
wYd3LOD4Q6uYwAr+MAzfA65oxP/suvpC2tgx1LuJQeSpWus5WHUzQeTHAcX2dYe+
wAVKHGD+BX+5nGisOLOurmLRtsM6CX5Sh0KEp0s8ea1BrZR+4GN0PmrKV/1dlimc
ecevsZan44KYaPHY9WUIlui4/V+r68nscUPiqRi3LaUSZSbN7zviLTYutM4wBWwS
Nfxkl9ub+hsBkHANY1wMnZ8R2GlmLZOYfX4RIP6rlmRSJzIlqrkKIAFMR6or2M2W
vt6t/w6xsLRarfF1qwnpmvtfvQZrw+sUAOPqfaJjYImja/OI3FuAdT1eCWBT0uRb
8j3rBbSG4ZcX6UdZvgVYCV66OsMCNtWBbyEKgpzAoZpdWQqwP6O5IRXkRBBd6kT5
Oenzj9HpYd/ff/yLWY7bZB4Yf6nQJO8MtGKbMjdQ2xGBb7Vkm84WLOiE+ZRF6Rf2
dqwXr98Wvrx0qaX7rbj0Z8ibCeJ+rQjgENMpkUW9Ql9UttF5yLbt+lWjBhN9K9y/
dTLO6VGtXHdVod1vxGAiuujpWUp9MiGwp6b4WKjn7Zy1puPB/Y53LqmBCNZTBVDf
9I6oFB20q56sWpqEnm7USOIdl/KK1EgG8rkXfg9QzP2CqHtxCEY21aUJt5CIUnKi
`protect END_PROTECTED
