`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLmca+NYuAxUjUph6k61OaMBlak2gEHazOlstpeJmj4X
MOINe85bIJ0Ro8++25Nm6+K7Omt4Qd997EvDMfK7uTkB6mI3Fm+l8C4aLJQ5j2CB
oXFnh+DpXrtr76gr+xF13OrGr+eW9c4yClZ2w0IGl9mNMm7xPnImiL77DIESNaAr
ap5XHHTSP5F4/eNFNTiP4A2O6we7jI6eUkgk1t/06FK45ufS9poGzXqm7Pj8Yvmc
elsU6t/Op0mZ534ZAizQPDYkvVh3J8B1WxhU2gvEgaaP5L9jcyXpzuqKH+BDcHDe
OZvVDj1UQqQsu0Iy/tHnfiv0s50ebdvdR9+qOeH5ICWw8DN6xPQtsMJ8cXqPQLR6
mqhyFnilb/x6i5u0pnDg6dYj0br/U0JVkkNl8qPfIOM5kbrWwqKzZFA/uFXr9iWH
L9F+TcEd3MGWqmro5CfNT8xeID/B4oF7yGlnfROU9PfNAlSa4Ft8235yOkl4w1jg
l8OOQoai72N+dEY08Zr5saIFGq6T8UpPoSr5As4wNjp9yD0M0f5924LM3RuTWk8k
8NNibisvGSPvoocOTtDYU0sT66JBZq3bhCEv+HVWTxlbrb7iu1kDko3Wo8INPsJg
zbeZY4wX7WCd5WndWRyGwvFQfnbXldF2Cw5TGFMORJWzMPUhr3zzH/OH0QkVKESX
JXCvqcdmPg5kzv4lhS50TqPYL1JevFRIATtNqvztWC8uYYr0u99EqjSad46D7EO/
ZoqKgejpNkAgnGEPMBXyD2tkaJZUXxuuPRFm0CClBeLhHLzbTa92mklesmONi9aO
gaKMRV6xJmHe/uOFmFs+WHHkRe8kkmpFHkZJIVzU40w=
`protect END_PROTECTED
