`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46+PLq3PTHG0FCiPB1jvjuWg+D/+O3ASVHIVhKzr2IdQ
WZnhNf18Y1a5U2pO20S1/jjHJrHiEf1uX1npIzJLFj5l3odeaa8pjTwTBqYHRtdM
xHNVstVJVnWqApSgxAvKNKlKcFrBHXpx+x7pgl+qtMnFyyw7hab6Ivt0YVxGX0P6
7pHhr3tvf0E6QACquRjmr9oauTQRlvMETV3ZS0aZtUtoGgQNq11mD/LW6u2mi3Iz
l2nKhWDp/bTta0KEClPBp8cI/MccDj9PrTPRzDDnxnGFcPs0MgUzi1e/c2D8xPA1
g5dpP5HAtQLjx1vqsoNM1g==
`protect END_PROTECTED
