`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+7U+K/HC9JjD9A9LUEGijrV2A4qouW1BWYsmJh0vner
rgCE0Qf3d9mzFJGKWZHeG/9N8an/Tt+84F0hHQPaso3gPD/1DWgbRX4kJsQYq+lL
XLcxkXvzWHqT3zm/dMfln5Aq6ewZi/cimQrvpgDycrz99DKy4j8qS6EPgrDkWzW4
XqF9IvtHQk5DN/mtbEdR5AlJM7WbtkxYKwiqC86eeiAX6nZ80y1tE6wX+qh+CkFa
38WXu99ZSKYBdPCD48B0hlIg6nYYFaf+BKtlJ/h0CKqQmiYYveQqYwRl3dqngoK/
fR6rOEXDmhRNaL5jzuf8M8Acqd81wam/ARzJfx13OGLZ0CNVi/M+CSLu/fEIgMln
4gwaybsShhvkltu08nyGd3oFVLb7MR+6P5aDIeqSg0rcsSdi9XXQKCxN/evdSLsE
v5jATMPWTk2PeOD8uq2c5aL1TuvVXKB9E4wJl0AVUz03AzfRyifEMM8n+C9mWFNx
zC3iCZ1VQCry/iAI7RGor/VSZm4sszPwmua/w6wc3Ds9290L6CmJaGPakB7paa+M
K2Ju5WNA8bkfWp+0UQFIme4ZM0e2njcQ03bkg8ghCBSQvVwmQ3x+myxcuW1ssYlt
k+2Z77MJPbWz1nb2TAZ70RT7qrqa5HoWJWz2grlZMPYwMdprgn9YlrRKT7D2ve+F
5jF9iODCSlA8KGmw/ZflEcB+kJyDBmojYJSGI5MVKQzdvANZZt1bnkEoxG+IBXV0
ccG0cariX/Vg24SEdtYcKw7CTtQMoK1yByF2N4ZqEf0NbyadjarWKlF41H6Vhq2c
KSHj8xI8wpo4mexR+i4xA+EMOvbHN3SlEC1+UYOTYrAUtl7KwLShCGn3RD/L14NE
vkO/ESJ50gy9FN5R9mDxzv4F6Sy/ssLDif9dFLU6o1H//B5LwmZ8bBaI7F/Q0eqv
1BM4XXyjnjhJifZrIhgCXaDJSO6dXnG/8sHTAG/4igBFA6euspZZTwiGQmbU3wTn
bi99htFnKSTB9JnDu7/aEMe36+1EZsPRRnqK4kV64AU=
`protect END_PROTECTED
