`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePHP7Tr5ybVI43w1UDUfn9abPI++42anr3ZIqJoQKjXZ
wdVS2OtPqaKc1kUXUTtFYwCa5ibM494faSUHuEXk94LJuRqBdOuMQxhxM2Gt3thZ
usU0Bx9aNG5ZsP5Khbw+xAq7OKITRO8uKBS78lD/RQlZmU3pznddxyc90IL9w1pf
mYJGUIZqk/9uusIUKEZ0qw==
`protect END_PROTECTED
