`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu467luKgWuMV8WZiTMCLXXmrpx4jGSP/lie2LGBvQKCmK
CxWq0t9fWUB5YQxW+cSh+OnaqbFcRWbkNvGshEXgt7o1+BRrYBIFMveheZ6btSgC
yTkj2ZGDvEh/cyFEPawZnw1cofo2fRaYHJLXFNTYsSG6rePsddcEdyqjKYnSbTAO
yC2O2XzrP/SIcD2cOUrS28q7yHPbzHKdUiVbM5Q5IWMQzvdGzu26GccBWmM1Jc9S
TEO2r9YP/908rZpOgJ6bUt9b0t7xC+QJ9hu9cZzrrquwHWJvwt7oyBR/BzlrxbzA
47S4eqRYQXSFVZLtdax9lh0GqiOt+3p0hIfST8M0XFDM/WNrACAzX/dIHTdjVDBq
wgsJyLs7XDIYmWQyL4bE+zPS1BJJGTxVigTb70dLG7cwsnZGKkK06gUaq78rp5F1
6xdH7n01VfhIOerIV3A7tSCG/wsV4VDgzrvzzoS3s7z1/iLW8eEdy6m/olisaJ4g
mBX1lvn5CV4PGNf/QBb1mesSW/TFlNohYzfchBjKWqMZWSnukjCQBBt0faWqMWd+
KG1/ghQlH76gavzfDlW6/DSgCAjeQEwiUMr0losDuibFlaYUv8pU3fbBpm3mzYc2
rCTipJgd0DSuM9vut4CNLoqQCLIvMUGX1ocLDm7oxAg=
`protect END_PROTECTED
