`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
77TIrd/+OyKuJFy3TwfXJNdRr+eA3aHT5bhKvE3wRIMo4DJQopip/SblM3ZWE3QR
XsaqkoS834eMxBHqn8PRyzZFHfCB6J44y7nLjGuxI7woeA5dFcGErF+dL4ot3ywW
I3Nevu+bU4Md4QtUCK643eKnAyrWWJgjD0jFupmd5ChzadjFqRYM8JUCPRWziHQq
ErBt0XAC/PiMJ2oLuRL3k9akugo4gKFqL/UGlPI3RG31ybZBsaalsXI23oz8obmQ
h+0qdAieOQetfxdUvYxzxkVhSw593l8RQ7hhBqT7j9D1jyegkn4rrBn6HFoTJ7xM
CBpAMlfQYOEDi/40JNM1pyWj4CRKtUiHMXmHtWPsKPo6aVl28CLOxP4YzvYm0nM4
n3UmtetRMCDKvVuYnG40PHSb+FLHax/abzk9upWJu1AIhsXeZfj0AlyxY1Zm62NN
kVS5OnfF1dmCVjaAmO+ntezeV/51S06dCCbF9XZybQZNX+cYoKxeyiqN+WHsRF4t
m86hdfLVCFgxUzeU0PiDOh4wIyjQGqL1Ge1kL+EwF2qBAM4u25BZCeSv9PWw5H8B
H41dDUWKmCznqrliGhWSzKvH2E3eW7WNRvA0+JaXk67VlVF4cbgxS1A3bhkw77jj
xDY4PL7HDUQQZKogI7KPLo7Eu5GlXJCcHvQL0s79tU5oFrhnhj7nmavqCH3M+uI+
NjWhAd269qXI96zTUpzZldN1CwPeTYbyfPsgntglKEzCBG8hK30MIVGel5OCFtdH
QosCjScHECTIuIif1kQN6jz4qe8UoyZqjWXTG18gL58j5JrCxVSzKCEscv7LLtGF
GPgivxFayh2ps+QdOBaPnwyzJ0HbadALQiANiSSVO2RDMfjqM8lRL7DbVxjw0IO4
knzuY5peEkgfYcjD5NA6ogMPVjjVtF6506QVQlqUWP4ZnwKqPwwk3r0x1fV4Cc7b
3UsgQs9w/gcuPSV8mbRfPtSDazRwgBOcNQmcQRBQy7dOMXL4hBcy1TNfY87kud9i
CjGP3hGEX9/o5+kKR9buh98BOTI0/7fSfn1p8BoUxprtpySISdxQkg1GP1iV7ytJ
SMNagi676AVxWM4+e46/1a/HwOoEI5pvRaeB9l1ZKIfchtp/XSAqhyqQgjnwh8j8
b6fIwItxOEx1CKMjKqARSdnw1+Y1RikeErevvExiDYa0OsBb3Ly8C2xBcwJLaodF
mU030wS7IpI5u8BwdjFCR83KAw8Wn+qNvDzPIcyzD/c5dFx+HFqQX/iXi+jSEkW1
pBTWbm69Tco5fEhONa4+ONAa7LfNFx5K/rMy1eQJ/wCwX3++iqcR12cnz09VVf2Z
W4bOkRUReHf4B661qrM6jFxwCMcEn/k0o1FZMrhJOX9ERB5jj942WBPcihoYdDcj
lN4NE0kKbyADi37E9CrlZ6T4vY1uLi3PHWgU9JFEvGKeUAYUBLelwj8SXTOhjPha
+5LttKhZdzjDDNlnrTISC9rN8GMeu4PcD8IPRfWWtIulRNgTsnap6CYfEJIvRn9x
sJswcVMtQyv90roUucqdt3XkipunAGzD4bu1gyXUhWMWaxVldGtjv4Gwf5ylnmt2
RagQrHIPBs6hVz7vTGYklYVBcXuQmiTgv5TrmrEABy1pZPaDo0K1wcBUS+yoO7p6
E4NE8yFJwEDaxzJAJSEcQq8c+Lp6put1sCeGVm3dgJF31rMC1ZxzrtW/gUQhWRn/
+wvlPXKB9UDUgLw3zYyFSUwGjpkl1c8CLgoRWV0VWd7V/hhizgCAyOoJ54y9cJUF
nVuvBgmqtEQ0tn1AKgH+JaClAtwJbrojXlnr+5WtGnXqCUZxGsxSy0JfF8LnsZ7+
s8TGpJ0eI+gaNhXsrV64VjFI1DutPDbhvjtyREbqHjAFRrhXyXlXNoRMkTvNBoNg
LLeTyJUgjruZ+qFhmm7zyold79+u+7HPE42jQz68lVpjkEEnJ/9QiSD6lLnKoAtQ
s2I6Y1gBgR8UPb3DxNeyw8HTH2dhJmRP8yG1QZpGEp+DiaxZWECbwgTrI3JGybNw
2O2NjkR06xYelErgVC04JC7VHfABD3N2nASIcO1G+W7smALoPCiJ6dYcagay223N
zTUGMYskIyQdZiN+5ZjVK2RD5lv8bCyb//oIvdWvYHZYH94Xxoc6IWDS9qcbmqP4
hZXXV4Fa7yLrtupXQstVKysWzgRcwctVzGooF4DkVByYZcaRdkYCgNx25ZlMOW2U
Q+fSxhbFBRKafua9zWO4JdXDGwzPVWi66aGfbiJvswqkLSuCeM0NqxPOl9CQCdNk
d6GRDZNE6EcB+uHWKeyd77FPxhRUrgBdKmn1dxf2v3AGDbQmGb9+KcILU9wdLn01
zKfWM+seDwA6c2iNbDhH3vnMV+oRCuGXNhQ8lFv2H0PZ33/ofc+cWEMrO/cwEPuC
LGBn9ZRQ6CPxCulBoOXMVLhFJ0R3+hYqQGw89UX/Q7ZuCoGnBtgu216+D79b1ba1
ibRsz3R1ugltQe8O1ylEa9LmHmtOFnKt7XPbb0Xxrr8hqENkAX55Bqt5Lf7LqbVR
ogvnVY+TvmOHeQtlAH26NuRXkW8WhzClMJk4yXaUmithKaQcLhjJL581E9m+vKvR
NgfHdRGRxpc5FCMCM92AYkRJnER67M4NMBzIhA87KM0KImLk7wtzVGjpDfabWQp1
rjVS7xHjv9nqErcPRbrAuSUgFmnWNFOc3MjmYGDBGhcSczGDDPZug3p/32aaWBwl
iCZ832YjKVGIKsksJygjcRpfwazpoZJjgKVbSYNpBDiV2VKlVrnTpkMRfUz9QjZN
eoiGhp9wnzAsox3wZ0+TzJDaZ7SlVtkZJiDVctH1C7BtqDKiGtKAPj2kjclSYS1o
cnqspvdn0HwaCCMxNGf0kbKJZD/deZ2kAR4BQMHZfJqKUgVRqSYhDSpB2brHKAIw
4DPtPDm2tEsbPr3AQvRl4WpcrtoomdRXq+NyGjZ/PrpgukKEhC5AFrf/2/r0YGXV
RW9ArEfzq27HJzwocp992gVAg5aRwUXqMG+psZMF8gagSnObj1M3jrHiRRPdweqa
8dMhEvnQZmVGPOQ4ImxcRtG9vf43rF+nfKaGERYuKwBKwPG/J1R/WMn6jsgSqvnt
BMvQ16yPbr9PMwDjE1UtqzLSvmOZOvfrryz6CJSHuD5a9TtYcSrijHBc6Erg6Ona
74uq0AJNbxDLgweKL25oDVPEANw5RKz/3WGAYgkTxkh15JarsAKoYHyxSrPp16R4
UbsEkjDWYyP260bZDBGPe6B7d9slQFalgggbE6FTXlvRtwcQSZ8PiDSkgC1Bfw/q
8CNduFzc0TC7plJuuq1PJbYZl8y8OGdD6OBURA5P1OjjvVUh4XnVRy2XEsfVgCgP
PsZO9xdj+RkiwUDHi87ZLNOq2uJ6PODUQx1Piku6kZ+MCkxXCfNaeSG9Mtd+jVW9
yfzK/TMcdhKX3jG59BGFhdOQEMaQVSakBqh3h3gc16Fgz75CL4r5//k0l7wB2qcp
Pl2g9vMswEPm1PVoHiOf8e3rav/LgvgWydXC0eHPsSLbaFlfWpp+uzhpsfOXOt6b
4t931jGljuXPUCwcDcWCfbaDjPFbHmhC+LoUld4+646bnoe/cvmxmMt17dNVckqF
k3PQ22AMh8cYQl0nBaZdvu4HS8bx9M9qjFe/CW2THQwufWJIk3U62HshPhREafNU
EJforFR9Vtb5zKKSH9m35Syryk1BuHjG+HBz6b2jvXbuLYK+6JOWlbWo2OgbBobh
gr3G/yDjX2O1eTk4b9QcSNoTTBe9AVrgX3l9L8pk8XMtY4JAVy/55ilr579kK2Ze
swU1s1c0v05CmjXB22VGdaygYasTWPA+Ufmy/xN7WkPMdz8LLdVt0HljUCa6lJNI
X/VuEY+w6Zjd117z8nkh51qC59TuTUGFiPfUbYCMv+5BlDdqun0tdk0uP1h/wc3p
1lBOGNcJmZX4VuGP+QvbzIlaV7fzcm042Mvd94ddyOmmWEQAayl8wE9sEQJysSXH
6zZYDcqWvNtqmDCZoCSTAfESvRBusnF6ruCuFgX3ymhBojjN9uCTK3QRx1Poscqe
ObZeGnErjq2CXogvD0bpjJ0xqEj4OnZWN7caccmxp4jq/5q1NUJgGVP/Z6jhOa8y
/bwLaOObgakSsfBg7ZuQvatOUkNU26w4qmYICgmsccO/H5HkXkDQvdpfzphLwFv0
2eO2Lf6T2vT+WDVmY8Qhn9ihZXKAwCQ9/eGajGDzugj5fdPEMW0MRfRaJN4ciIb9
TJrOFtGoNESNrVItJ9SuCYkYvKzeRlGWEl1PZBJekqOCHvViVR8T/MMtSXU7j3bK
liGjAfgseaNeLe0LelNUTc9I4p3gsyhxh81fmBxcAqH/OOMchNRCXGaVKiCBGT36
XhuEC2ekBPdMiZxZ41/BEh5Ydsh7AcLyK91vV8dmxuelslSsY9zkBjUoyUnmym6x
290QS1jTWkPzkdAKZh1BKCO9FBE3hRZAaLPJe0wJ9CjGNYKMs/+qJY8+CzRwbF68
PwSgt8rxUx237X8MlbqXlkewiK634vCUU2jdf914hHQGZfwjFlSieZ51D4YQyT48
hTesCZ9cOcFvhuImZ7qt4R0fEjUqGbHFi6OQK5SO/3B10I1Q1zvKJTHE61koY5zm
RUycMuMtPu0DhzGz3md1M8KGoJ+kOFbWStuONX1fN5lSdCZxIoeJFqOrT3Ug7+zM
j6XZe5IQDmOQPUH561h1/v5MA9c5Hb8F0lkWg0wcdZ+1ecY8gHKmBVAXVtr/ulpB
HI+/l8sI802RnJxUl9ISV5n5S+J31afjyYUeV+Y7tXLB9K4kyeIaqJgj0xCceYfW
kEkO9XipcfXaB+7Lw7n4I7S5DyW3qbTfbIkANsC1lIIbQz681S07kQrXQIvsH1+F
20r6Vbox+quSvhN6fb0tCNrqRCKG48zCEoVgwXgSiZPvFqpBB8QqL88Wxjd21/NO
U4HF0h4+kgcoZ4wl4me2RtIIOkB4ShKeeqIZp53AxGxsIyI7mIVrlQSFnibNjmPm
b27EXfAdbEnlSE0WPzHom5BZlMrQ2+UwWd2Iy2yDf+49OhzUXLnf3VKjX4o4Tuif
Bag3aGzBZy5UlmhEz0wk6QzLJ6DaMbKeckPiOsKSEGErpFfv1c//M5yTdOEl9/C5
Q3yVAP/6f9smVGl8BqsCA+PwnxnBXDGKpI/nToTHXPw9OA1HydjX+LLcAXDb1YEV
wHoKBk05bHoLZFur1rUu1UDtl1S9jEtTCQGzJKKtZE+ilXm3Bk7WWZ8b+uKG7vaF
mL4zcxWab5v1RR9D+t8WruG0q4AtgjBljv+PAT7CG/cuP5X9f9OxlfKSlYKOzgHN
9h3/dBVKETbUMrsKiOkWpxoZf0zmnUsW0sWxTtg5Jy1FbnFiC5QPhpcNna/v1+ZE
gT/WXZ6QAUzG1JQmSIUWbTaFt7Eou0MQq9brF9zUPEMBKxnEHAK8rHtdjMp5cCxa
GMKfPVAYPX9N0E/iz+cesKr05Ah/7uqwjGT7GkNxZGjVWB1YB/JJD3+kmsOHBSXP
y2feCRxKVeUtNY6z6rJk1D8NjZMpnqx7YLXnZV65hNHwtY2BKcZTRKFsFbGGhL8l
nKvTOhfCqBiKxAkRHVRzhUEIooDppqx8OYy5f+MI321Xw0nl37TLimQ0kgVlArtO
GKLuNyvK6dLJm6IecKUsTBmDZ+Uaq+f9QVsk7toWxiAXWqDGaSXhDNHtaQTcO24t
bNf8schUExDQZ6nRFJVnrtscoy4jOnDYPfIn/OfuymrzzbDU3Wpwsd8uvLrHwD96
gJwC7mDBBBzYS1D485smcCVpPvhnyQRKJg2DR1vPkVzLsx4fAB7WVIDT/cAoUU15
IiRQyYEYWckwZ0MvEBg+k/J5a8B2MMgRwx1FHnqbJxyyW1uq+rDboDPLFlpPzsiD
+sl9dsGs7hsbPNkRow1zV4Q6UaZuAhmyQgKrI98UD0M5TvQIq1hx9t0Nh1yD2Trl
YtMXZvHUq1cSg5uckOBzwiScQx4N6tER6ymRNitUU5/yFIGluBigA4dp9Dl6x2hu
6R9zQJcB1+8DONV7Kf7eYH+a4uWOsXR3ozy8P0kkbPuG9tw9opRY+cKL6Nme6zcf
psjTMM3eKSoxFzg71pVa79LR4DPD05RrzFMWmpKQ8QSu/hVKTybumxfQHWTTjyXY
FZFDtCsPssfxDm2z2DHe7AUD44oU6Bby8E+gQzcDnp44bFP9y0YN096mp1u5JPuZ
5OzLTd3frFkJGvVpydFp95l37+XA4FYoPUJE8+fEgbLO2k8WS4vJWUfw9YY45lfO
u0f0z5QCl8AAhthg3QAOAdoOncy/SCalglxBceeB/XPWbP3RXwBTacOCH0v0TiAB
yQa3LR4jIR0pVdmqb010VbhizhJva/1b8KOLe+1gxnEfLWvhRxaH9w7PGf+hXCmZ
5XHQDHBajyeS47K2lJAfcaGl559bspgfEp9oefmsl2fmx7iFzbI1Oh2lTN7vNnki
FC6pGLXmcR6ATXNNheXs6NnaXTtgy32ZOU0QlpZN4V/18HJ/hhWm4zLa22uiVcam
YLdeWsssxNLp0q3nZ81DNoGZiofC1810YPEYzGDpfZX9XQuTluDR49Hkilk8Foqv
m6bwK2fBqvjzkGDvyXp6VwMWAAEZq6je9n66kbx1a9l8HCLwxDofFj7HPy9NfkDV
Ev475fxJH0cBPGCQC5YlQZAs9Bojqv+73XPHNCDV33hvpeB2e1a5qOmqp4SiM/Nm
NjxmSpR8/HkF/qI14Frq7iEjt8Rn3ihreuATdiXBGsxRQN3gduzRN9jRd+xkt85y
dhVf2eEmqupG1jJy/qEUuJawE7GpmPhY/98p+0jKSVQBglNTSNDDVe1Z02XBJIxH
y81ztWLyNVcvHYLn+5yKoXxJgSiH9SHf2LmBPYihJF1Ut5ZJZqgIGb3cuCATHBPf
w/QcAf+SqnC7+h5HG1ZixgBhC4+HlrFbHbe7OsMsw9lgTKf2V++B+elp4neqVdV6
naD7b601RV0bLlqpCFmKQActi85OPy1P606qiZU45YimMQcZ/5nPEAFxtOA0REpP
CqAUfMRasV7fs4dYuaJn/onSUaq34S1I4l832EwTraA5Gkn5FKxP2AysXEtlx2/3
118lPYvRswMG/0p5pS3viQ3dvjUmLchIBBsKridm4QuDr3uegB1f2C3v9CVaqine
6CgThXeqTiiKa6Z3RfGDwR4lHdwJD+SaGuI40L32OncPm67ESiSqq9XDkNHi8fwT
Cl8oUR14muCsortKqtMLumD1omoD5dBB36BzViua82hUQlJ5tRk5v/aXvGAWVRIS
TjIhEaSLihN2wwMuRq+kp2m0d81ZhEvQUMGrhtEwAsTxTnKJsxYBPOxKiC8l1xuz
d9FdKJ6Rs1N1UN5EVy0HLeb0UHZmD0wT85L5oONfVPHQJQhrzSfULNy/p/1CvS2D
ZubDDunbhYrXNvDUiM0XsXXL9pphZQOw/Fsgi2BsbZwQKFxaihS1K6J9rTK6CiQx
MrXOqTp0+buLty+TB/1bpo4SQ+otHOF1UXdF30zqweDSKL/l7RjphCu1AXCGxxGF
RK7UmNgeW0kEAdBkSSfoqBknlwvcT3B9xBy9gHPlNjpNiNiHqRr934u23Wed3Snd
S1O6pytpkkchfAI9wBgghtB3wt9IUohRGoHGCKBQ6j+4TAtyMmQNJjmo8U224VNe
vMteZgyChzGh66GfjPNy10EZs6vdkz1p4v5hxrvjEIphDRVmfo56NACwgBEA4aGF
yVaFL4psI/vGs18Eq9gUSeW2h9NxcwFG24eb+Kchw3Bt1UQ3A4zqAl1YQwUxrdMB
yRxvuPFhBVJmVvJAYTsp1mFKyAAd9am+aNrzFkqCiYbhb31T5ZJ9a/xIMJ0hcwH3
Jt25V8Bmgv8vxO6lrV+lR5p4nmn2+R7bTtiQmEKKMAmUBujNtbOco4TXTBEEtFIF
kX6n06b6XaygweKOR49Meyo8QIThxtiALSc80MwR+7aIf+stulGdf/dDdiAaAe8L
uaWXAUSnQ+KI/oFEVFHj+trvHaY2ANXblN5rZqxBsjSVo/hGWa3AvCNX8kGbdMYs
HNB6ilhdWQPMgCBNru9qa2mblbp5+bNX22BGERBiwzjii/XmzPJdJKhylzqm4r+Z
9Xd6p1jjRYp2pX1Z2R9q0NEK40UouhmVJiZ2rSHPw1bHRtAOr0r7to7ZUuQ2yIWR
71kIZksvgNLn1tiwJv/u7Mf9Fa7Sr3taNBogN9u9R+Mp8TTWoYww0Z3xfd7bm9/J
Wi95ZZcmMpba/d1I/DgR+2XS0CNkGOcR3O+hPV8fD9g/6xS/vlyHLkOpIdlYcP+z
c9yUKlY/RdWyRCToRFr63ORF3bfpTWSNzQY+3k6gpWrOhL/M0I8OAAKEvIzD9+jO
qM073L0m/wGgGs22LjMmF9BqFcCBKjaTsW1MF0Zk5ss0u5u2cZ+GXZtpRP/1y4Z2
YfRIBfiLWjbS94ue/b0rK+nZzdhWDsE/vUUQmdYlhP4HR/2z6zxo3CSbthgpfh8R
AS8SFBWX17pR4UCPWg5GEClyOTq2KiWVEBXgscZotNeiFK5QqshuDc6WLCkg3Fcd
g6NGbCX0UoIIv/mq8GC8dGLeFOOXwqlIEHxhqKR4MSwXCqmSUVEu8y+uBDB+bqw3
UQP9xyWVJFFpwT/itj5Ec2xU42uH2QjmHy7WzC9QCj+y6IK3xo+8aCairLPFR+ky
sF7XA82kF5qMhtegY3nlO0FWGXCxiNdov2rwsy7q0oIzoiWtXT0oVfvZ4+P1VzSo
BtsKmQIzU7pgjL54qZKJZwU3cB/f6RyXsnaa9b61JB8a3a8bYeCGJVRPMhxTMgbU
qf7Paf0ycWaMfgwm53MKJ/kQG1mPFcNQ5L/5VsuDn/0AaZMheb6D08cGOovHryAR
EeyqYbg6edNxGCohqaO1MCQ+1W52hCMLtUkW0tyixDvESs0Iw6kiZdE8WZx+wxPP
yW80UWOOJIiq6/PtcLHm2yJMbTI6zbyLYnCGTVovTMsMyHhvgoZ5BnLFcrnr+mmD
6qY08Eyhm6TI+sdNteTPUUVUaxGNMyukR8f/xsO4HPtOXRlHCXIvJt9Sy2yp8tor
4U6GeWfId/+j+VZKzp+6CmCDXxJ4pZq8932T4BpYWlcpaWHNd6+EtBExTsj4obYL
O24D7GvBwr/yxaNFU2bM/GDbX46dTbzqUjcjdqMJSJMbK4cNwv8wgH4NFQCbyo0g
zwSh3fGTOcqHrfNVxCamQF8yL/jMwcL9qC8PR8xv37xTf3dZ/eGNAzzLj8oG1Cxh
/fcpPixAOnZLdD4aXi0fDqav6n2rYbTIvMyKFQzECOxYTKdJXrrxiLuH2H70jN1I
XZZL5as6lWoNt1gafESvpQHTtztvvebaYcYyBcoBQ3l7CITXpu53T700JbVu/sNG
DhC4cDFlRNCg8Wht6qsMk+nvKmp3KtuWKgaPavdqz7hWLpEFunc5qztfvjEJaheD
Do0y0JpiaqzWgQn7BOrlwhL5YfDCOaCARTCrVhyiut0x7hGsjJj+hV0yXoYW4zhF
ikDnpsyJrZgunMEYU+I0E60sjB4b6n7Cqc4ZtSsfuA+u8Swvc50B3n5QQFd+xtHI
4duF9o3K+pUIe+XiApsHkX9Js6Y6kgT6KFC+xrWM/Y263KK6lIt+g/eaCwCEVEhc
5yzPjhf5KHTLhtUauMI6dHeEh3uVbQ8NrauBOCZSf9wrQQ/t6fc7HOmLWJP710sP
Y+W2qyMHDFZmNNDva9uS5pNaMgKLFpVHq0/opcEvpsJXtF+AJnH9zBfVgl9Kdsn7
gZyTI1fwZaD4oVBTGx9yWn8ZPTL520Ct7ukSGO0z0AiSvd/55dnr4ps6kS79l5pI
Xb1XcYyi/nVD56ZBdpwYrGQmiA3pvRvNRrKgctsN9L0hqPLcXnw/+0kkOvgtrV0n
2wOmgQ9aLFhPLNrHXZu8a5xPyHMoLonU509n6PEPPsHJwJ6cDr4KN/v6EvSET4ws
H2NhBV5WxWYb56J0G27mVAU3XaZq1RUATAHOV26Kuzpoc5snu6ScnnY5tVHDtJcJ
P6qWqg+2NReYwx4aHMfPgqerPuFr1zav4J+IuPr+MMfZglIPlg9KeApi845+g8kW
mvSrNzlzZuyJZeGA4kixgYzGyLWeG9rCTwRYY2I0wGv54FyLIscAx693AzsTOR6D
71pA6rdqznSNDbf22kDM9drvt6Cs2tOXp5eiLz8B/ZrQ9jlX8quLVhvGS7I5Eedm
eOEXWrW0er8K9BJ/n/EAja6j26gZsmVCaFjy+g5nBZnWI4eHpGe83SKtm8wl+Z5v
bTJxm2VVvQKI0gngLKgU5qaLwX2rM88ws+BOWKhddijcyqGqgr5O89p1EiWxU8ll
btwy7/BNeawINBJV5RbO2CRaVChrLKiKe+C1kZzey5uYXIuJBfhF0+22bEwQGm+N
euiU8u8/7fa0h38XrDYvyX0iFpmEIwwTE7wjK439kp523xrRf98H+YomZIhbAVDi
erwWscoTuWo998QEFOEIHm3c+CsRm0tMZ50tjjy/WNfS8WM//ywn7YhqFA2/FRGW
GzJe3OrWwxJUBcZhqXmiOTa6bvJ5nJRBb3QdkZsvD5WrA9Fgt1Glp0okySmj2xVX
KO943USqCaCd4fW+kJIM90tijyh2zEw7DEQpEFoYooZeQiJ+2sA/z0F6k3x4zHpC
fa78vgjHGrJ7OhlGl62a6afA4gTDiWrY+DHMcNR9u6BbMiTbFF/kF72LecE0l5nT
KD5isHxPlCZWvbTkd8vDJoRpxG/8/NXZyHcbrY9zm3VhvneNUOuPUV/lnhv3uwov
lKDgm13pvGuQfTmVPg2UKPAE7B7IZHShOsyNaUHGBTXSPNSyuKhU9xBY/zQu+9tz
HMLhrdzPjuZ5NGvE09x5K5VzDpbBQ+UEDoJ8LosE+QLI30U4CByHRB8fEnZPbl6U
u5l9NkC/qHQZfZ7iYRSljXdpAXOSqnzJEL1p0xSrv4AIRTZnCFwy8+UrwbzngNIe
7KkBaHN1kwJQbUqtflGfiSo98WvWEcohv6oX7g1hKC9a+Ao3+5FAcQo7XICfRfos
DyJiYWMmbPHWhs8yL6ve1XgbNfNRJ5BCeGl6yR9WSnkaW/Sf34bpPs3+PxQmCMxT
js8zPRnf3KqpKfeYzs9G0CLlqRK6D0NUue8sJMEcslonK2p8ZkxU1ptwX22+9D7r
K6WcORI1LWnSxXOi3UX/S0hiIoTpvDNfLUm0XYXi18HPrcIrO9Y5LC+fGzG12keW
4q0+S+eKZJ5mdyvO9X8E1eyT8gm0Qgpm6bNIJJcIKkJqcmoa2lSUkqwijXD/W5Pn
qU/zquHRjroMIA54RlhyhZ3t5RuwsU2tGvr+il63n+6mAv0omKCCLbX05AIiRgzo
z1oRlN2/3I+S3OZAgMaQZQH/JD+LPC+O9+pJWCF/zu1hqE2oB5gspxz7xZUvDsae
0F8QOh26yVt8sr1pyIZToiFC6MNSAxvDhIoqGL8wU2FyHI7R617GoW/n++JqFfGt
YXRJrPpuQVS3YiPTmBgrOJx5KeRArSu3Z5N2eCPG9WKsdrj2WzB3Qh/5UQSMgeag
DsZJ82D0ujVSxZmMJCvILIqsLF2ON5MLAVpl3FXIb6ckkZJtn9OaYDP3eiIWWBZW
JCKVJcrpBdx++Yz+UbF6UJiMYUWOfar6Khoo5J1EV93b+lrpxONQ0E3roZ2X67j9
NLQSOhuIeqI2C6VsB0ZcScQHoVhvBd6igZ4ZjvO04xyH+LvCPIUfLHmCarvq2nxC
aD1H01XQG9djqPmBEP1wmrg/DM/jZxl4PpFYwaveQGxhddKuSfGkY/f6afvHMz2K
vKsmo4d5Gsy9LzBe5MvWlukVqLe6TKytdGMrq7oQBaULoKU+Abj7+w/hReKm5MeC
6bq4FNzXkplyInQS6rfI62cum1MwwuLwGDscJksaAeTaf3VmbN7BogVUaMTVy01w
vSbzQTA6Al3Uf3i5iVQ5mhVClU2Cw4O3tMAC+7QeEiYCSzFHU70bcRVdha6lf1c6
8Ick8QDhDp2fgGvxFbb9/Y7Qi4OP+n+1INfmHBbLJ4Qugik3JPVOOMBxhnaHJ6q3
ArUD9/JQDyw8rwQ9McmqaRyt+wFbqHCUh4RbPzjPaGjtvdlXSeBkZtz2jXhlbezK
cEAw1kbBpIIKeDwojlu+oTJXySBS9QpXX644FFDAy0Qgfp3W1zouGqn7l+F0xJpU
KXOg/Dst73HMw8rRtms15VoVYANaFeR/vMfvuszawHz4wnPnV1Iqv6vJTfEFWuM5
D9aI9eHbGOXdnpGb/7+8F88hyr2S6bXRZ4MqfWCT1rKY8sIsLaXpJE6x9XtXbdYo
gu2Bp+NoEgMU3z6MSb7+G0+qNFZfOug5LiG8Zvkw61sbNZHViCXXggbtFLRh0oPh
+Xvk0jmVEGm4ItfR0vWgR7jYh0P5GOZ+LFtbLlCBDdQRg/67RNTGcX9jQBgqnoMU
f1/ggAuLxi6880B+se3F50c0ARPm4RgWRZWAb5RCUBPO3nwaDLT9hydVDSC1pGau
tVK58nf6zgg16HQx7yqedPJoNNRA5ihyItzP2RdMCCv6bcJ8HtDvuI2zsjy71ii5
IF5VjtiQV2GRGNSI7iovJ6YhQnHdiBnnGwuDZ2tpOa5/gyHkMrbcA4sZJRJh1lyp
fReMySsQPg3/x7jMt8Wid+wGZy3tYj9ubgq2GEL9espbGP4wyzHmmR1lNh+lrKn8
kasH1Wig11GTiNpJwPoUIvIErDLqvAtZUuXa0/qZNychStKd7KpqGQjZN5DkgWcK
D8MEhutnZufThR/eo9IhIDc+X3/QtLou00v1ZHZ5aiaMX838mGQR0LeD1i3A4iBQ
OIgaLEUNx8sjnXqd4DDN9jUFaxmeu3h9xJV+J7GsrQPQfpmDc9QT/9uiDgKl1Y4G
SJB/wfvCYCiIBD+3VPHfC9Kmsgb1myWbSppuAyY1xr8u40ScSm7SLJ8KCWRF9GuS
LxoVI9kF26bezxRI0OZQ1u9SAy8CYzbjO9Nel+Rddb9j8vK+C0kpmf2qJdpRUTtq
4quQIFlpkyifPBv3/vUaZDNcdp+0GvLwvCXPU+1Il7TMnzsG6vbUr4HiPLvuePfV
p0VCbHGGwaMTWwAk822JbW73NIEQM0plrreSFpALSWPWAYKg0byiPqVVcbB76QKF
ZJYicTIRB9eIaoA6W83og5qXGZpgAKT38Zlan7JvR0u7l20x46ZcgXQDfURSERjp
mODP/mjUBT3JOgXlNJH3m8poDN3DgA4eA98SkPmhUEdUbl3Cb3YLIkS+49/WR/d4
b9T2oxeTJK3VTFpHlyXjc88exwjsCG35NcBRb/Mfbw6gUd4w5YPd3tk9GGx96Jjd
eIN7XqmeGE1cSOBl9qsf4C/sD7EoHn05Ow7+oJiAODOZTZ1FpFXi+oT6iCJ0P18G
5Dr2u4jKb9HTLwWUFeAemtE6UMeNTBnDx9XN6/F9FSbGRodCYm2YSahoMidOLROW
7n6LyVq7l/mlY2Hpc6wdLXvxDVu+1oZ3iJDnI8M8o4iwFpSO8OF3bHBoKQiZy8b5
4OYeOMiB4xGi5881dXA0llonGv7rrQph9g+6OCvkfsu6IH0mSKetn5CULrQmgPRT
gjdJ9la5LskUzJWmQfeZQc9YZYDT9l01E867+z7IPOldDekjAtXPNXcT/B6UXTMm
KP/AL70zomjthtydhV234fb6YAEkAz3jAuINJXID5MxBVHJUF7Jd0Tm62a85mbrp
Pe7keHNmkOs9BM3+IvdPQXlZOYM2cLWO8iCCEZM+Cz3tHnAEuQTjTn1iU6kB0YMG
+LioBVxivmrldpSgUa0yBdNT+vN+d7tyPDBUIovrs7w1vgY7VdMKTwjQa/KENpOp
q5/gIt1QZp6eciL4vkmksC0g/ouiTeryDOH3KMUjtKO/ussq14OcEPFq5sSWZz3w
KljJEOQCuigilsnyMtuioezxhX3casUBs20P/DOBfSCeyMnfvPZoDhTa4cVm8r9Q
wGMr55F4UwJa+Sz0T+f/2iAjIGpDvLfZpOH8UW+xIRBXg3bJM1cvPKRQ5XBwcojQ
2pwtjy4m07SL+qUjWSccnC5rgTBBIqV3lCi1awi0lVXRrszaIQgNE3eJorxlUPEm
0peTZzSOqD/hzxpLkq2lil0+jHnRZEUoI/bUozbIm/jw2P0d0rk0m3SQT7Ccvih1
OlYAFrRhHEcsd4XnljDm7LHINUnh3aF37AJdW3NUNWBUWOV1spuh42qWLiXyrYiO
3+BVBamLK8KbHWY2RoxuYoAJhPrH6kyvGuLB9fGKNY80WXZORTmsIzCEo4sTx1cY
5Dw21+avAx6ug5vVNPFwEL97k6IRE79FtU2vMI/sYmbFa2SFUaIE6iu/QSynxnOU
SKo9d+2JkkEoqBpRDO1Fi6RkAchbwCFUhkSLKHtWuA11VFpLQ7KP5J+b00zwSo4C
331RqBVLpAlR9qdIbKIyvF5JeuWFhoVyFkPdhe1LGYpYAkwrG3c5B4vcBlw+qQ8Q
dvPBIVjxm7EjvTpL30vftdIYsr3wcYpwaE/iVCQScCx5SmBJo9ZDNoNs8/tcKZnN
RDMqETKlsnqGpMnBonShWffz+YDCIYBM+VWhL++705fCEgtvSCeT14NNSTJvjczl
jNom0rG8x5bVvYbjAj8dIaoQVgrh/jR1q5lygCn0/4Ng3MXSUs6OKjIXrSy7uzZE
wsjBqIKb05Ozk3wZLWCcJ6ltRL3x8JMwdiB+eZ7rkL3SOA+/qlZf/Rp7HbTNEiUj
9AD5qIa1OSJO7xZeGPwQSEpg7+oq/k3YVIw5csZlm81unKyhdzXP1uC+BitiFfxk
T6MW17/9DbR38TyeSMRsXs/asEixcY+3SqNHQ7oNoFt8zdFhL9+6V+GPvIQbNa/N
V73Biw1AoZQi/oYsAVV547zT14cyyu+GtX+KNxWQbSfaNnCZynf71o7fIaw6RA7/
6ZxUvZ6MnZRa1+nxPlR9bT1QPU7pWB8oIjmTs1f1Iq7FCaqmoKNfoQWyRqYt3bDJ
grjruSVpigb+McGrn1wQ+W4Xw9jenWOKmfWy+wmuuuusgbwbg2MKx5ZmNiCkHl/W
IpgpEquoiHi/WCMNeBCPY9jy7T6XvvV2yZ+/SxMfNvO/ZFILVWSlyRl5AsR/+e3n
LxsKSa7VCQJbTJN/qsMi5N0N3EoZ6GnQjV5ltIKLdwna9VJGhcflQUxjUv6OafRy
5+M19yH4GEJK8toJNBJIeNrR1LFCcOvtBOjwK95XJfhWt2xOZl8Z2wqEWHi+GWPb
Dna2O8n5tkRLDLoIQ5u1ybSq8Jvy9pGCetXn1mGGFpqD6uwDMfqutff9fX1kRaf2
cAo7SiyZK9YNyFHk2tqA9BxacxwPNbDWbUm2lpIcQyd1P/BLprghxUnwc951+ZQK
v5HlrXUpfPhNawsMzGYK7R5FHoSaWYJYZqOOSkMWJjqtr0Tkzp8tou8RMOXx1nXC
2E+CFCfKDwLJeclHnb6dozUKGS5C8xRMe+tNIjxYo61J1ySU+LQeZJOGSVJCEqB3
dl6CbsmuhCOi05MDuGkfbzv0H1Av8CCNZS2VSYB5l9FNfI9eO1ChJj5VnOEUvxwS
Lx/NqxdTW1JwwVSRgKpOc6TKn+y7gY5Tv3Rwa7h/jb5dSgRLuIMk78GfW0neODl+
lGcvIYw0husEGnVKegewSle3ydsTkuTiewXVY1sZYw+eI2OLRV3GookNsdcM+DGY
HFXfLFbNmS9SJTdSG53qyf2oMaUTIut2g8aEQ0Wth3bMPm6/EaXHrYPn8dn4KGfW
SPVP9nPFbT5t8+qDX9gI/sgsXQHKO2lEAHKJKAe/fiYV2aMHmw08olFILzJ9n59j
/SP6AXkkSPMYGCQqEB7dJKBQusM72rPv4sMg6kfHPH7m5qfk/HZnHi2vXsoNhSoY
`protect END_PROTECTED
