`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yBU4z3c/IsvhT2Sz62eiHQtz4ai01KxOZCM4UhRZa4h
SBvEuwfgtBB6Q7cjPQff0dn9G8CUSAkzv+ZVPMLTwUHonVBhs/eot7Y4xvd3bs1w
3JQ0jOY2WXQB8xTUM7oNlyAIvoW+Mr+Wzs8j1EZohmeJE5OdxRJLixLFayiZfWeg
28ccTWOyZ/CZGVYyuaTMe80y/9gSXdAygheMYS3g1Qrqte+qU6hJQr6wLl5WOnXu
CCJ0MZMOLjMzUXsKqbGmDwu90yAeClrSNvQXpZIRfHOR4sSg0GL9k5QvHef6k68q
+JS9TIwBC/B9bbD6Hu9jfQ==
`protect END_PROTECTED
