`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKHqe781ardhseTJtuVtIBPl2EFIu0Ka/S3aWVZFlOxS
XC3ZeVxPTbPZ4x9OYmh+4/da3kGch2voGtMY3z3zK6Nrkr03+7N9Ku7iLr9XiqXk
OSOyo0zsgkmqn+C2op2ehbJ8nx41mhZwE/rezz6YseVEDgBnlS4jo85O3yyirX8q
FINybf18r4i6S+inGu3BDFy+NlPN/uSYvC+/Y81e9Xic9kMfiPi+h8vDbpNWG36y
rTfS0SQTbsaCdqDcPltiMm240SUBZ/B/TIWlf6RlfzTMOzCiNAQ+RRAUgEwwmOY9
cDO3vGu8lnTqLGX4b9BSzrUxIc7b+fvSOLudnFbBcVsGB9vaNz+o5bzf1eNFdc/s
E6JI/o0VUMppsBTZ6/28BPO184AWgkLCZ9OaMDIzQEM6f5ao3l7NTpZvZ1tqtzNV
rkCboi1swNBm5B36OWAtvW3r17u/y2Z5Hs/eD2/RKM4lc5x8t1/ZTtwY4S3iphoN
VRE6XZ2cXTAOyYlvL2RzWfUZzxmUxRjtpRnqJLGHlIK/x+K3dEcpLfpxuuBy4bry
89Iw9X5e7q0UqLJ+fHEDTHBqIKC0LxmS2kEXtjweF345H84DhVBoisSTotCbafYz
YvwCp4hEmhZa2vUpWzGQamnuLczoqVzBb1ZWIFNpuq10QvjVCQr9/zvjlui4MiZv
`protect END_PROTECTED
