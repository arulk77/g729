`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
H8QcPnoa/F6ScUuvhUy7Jnj02fEbplK0Ud7USGaS64S9nWFAusb5Q1CNJBcSF845
Gqp0Cgyrpc19nZj6iqfkA867P+FnSqXax6vp4d2iCNbZdQ9eW6pPva6ZNRlHqePv
iEn3/k1CBcaX7x/6L1RuosiLN68E6/AIGfSATp47gr8f9LDADxoQYC0+SinAYMgD
nETeOb0U0j/2Y8G/aXyJovfVOV0ASgs1RFHGX3mHgQc50CAT4XVEooNfhQxK27UW
KIw/4EcCby3HhD2QKL237OXHDHCGnp0SCZYnW842bvq2ciz83zKdGyFde1xyKV3G
bAtHa3dZCjohldhfPjh8G6umEYDvy5NNGHNxqrzeopDkFf7EJulur2UDJRNRtB4z
a73t07kcyGV9XamF0q6Dk+lYvqls87k8KKXQ8Wi/4Fc=
`protect END_PROTECTED
