`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42ZOdABdvi6EdzI8K+OWOR8i9gEsvu7E6CLlo6jYjDZN
8vmdw4UZGXUjkUnkvDrAAgLg8gyKQnrrS82sgr/vjvBUdkntsoJ15FOFQN8KNM3r
KBl3khOgWhkoyvpaNnH7PDzNEIrZaqabew9a9if+CByLcVRC1h7WNLR73q2Qjua8
5dF7wR1xxPhdAfWxMu/xGZ2BQXM8luZmoybQs1TCwDK8R3KQM4Ss/ckKkb/y2VzC
y09il7SZJBagNS7iFGgvPDg+raVdQEn7kghRzN3bh6QXab0uvFcmGXXACK1Yz9mZ
e1IatYKGi5+18br9m3vghQ==
`protect END_PROTECTED
