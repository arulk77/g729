`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wAjhEkO9JPcNwyD5ttv3j9uz1poF1hSiqC+STXTbu1G
Uc22twrnNQhvsM7PVdYUhv10hx+vGOVNpv3cb8td7NtCXOpcwPQq5RRYYnrUpjaa
7NHwL75bfeYV1OWcDwI/55Z7Z/+/nUIHNEIddawJ4RCl2LzaLCz4mhEXYrGTIEvP
5DpIOg8mEyf9C81d34AkqqrxVsgcg2Pi8EHK96Yedf5tSrtmhQUbEH9AGmN32Vdu
8QTKG9shig5jDSD7PZH+rBUgtoL/lp9dZ1791YJ4X5f321NuDA9enwyCRb7ih28k
HnLKXtylEmo0kUZ9xkfiEw==
`protect END_PROTECTED
