`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2RtTiaLwZbJSuPbraFO4dokHEquo8XuJ/vIt7cgQOooN783zCpFmTXtMowRU3iSn
6zMM6qc813IPNSNItcwExgeyiFSni1LOoQIkEWl1dDLIROkHTCz1OzzREZLRvFqR
FWTIVhcUmQtz4erSzIk2NuXRqcSaCyhO5ctt2NdK0SX1quRqSMdHpt3GBMnWbhvu
`protect END_PROTECTED
