`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK7PcHSh+EgHHHKt1lbfiBAGjmywMcUIHROpBZ7k+JQm
JqDL4vuyKOGebNeZAryXi+kuGcsGZxaqWQhlZYdy6nuUM8pMVfpP1Wsq4AIorVpi
WDtnGfZ631ogupws/valYXRA5Z8MQw+1TYKA23aai1Iz7cmho/cMCHttL5Vgzf8p
xxi65GRHtajMNqiGIemNTq3/aXUWPIXH6SEoRjuneV+WCPcoMmMwXDDKskCM/s0R
P9nbssrudaA7n6qwZCBZx6W51s8uRkF8lBWt3hotn+KdURVDTbjcCedWHesZ1LFa
P7wxW60j7hNfiPqQfCaCG/b/yMzRpTwZkSGW3RO7U4j+iIR6HBdZFiKG023J3wri
TauexlWuJJVO2oiTs+HZnt4DvWDKEA7YKB4DJ4lvvMkOkCdtx5SkSu9g9sy0UwX2
rn8bI0+ksj+qoDeDZjhhGXxpG1GY2uDJ0ZIhdHhCCJgme9BJAzpjIoLgqhrHN9X7
4yksBIB8m/Cvq/qoixOjN8DH/P95Oi5oL8kJItsI5Ag19CQYJUTr1odIBvWVqNEx
`protect END_PROTECTED
