`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
tfuioo/jKcxnTREotZGS3Dfwd7Q1CrFC9S+0WzUtSJx6OrPVPHFWDAG6GWyozwxe
Mr6wRH0o37iubDVk0ZUAeG5QZ9jyb5NmcNFOF+8PZI8BsoITiE+QiQSRsWP2Wv/k
TiDDNDMVtXDgGgJmDHdq+KVXpWB/yaAJ+tumiEqkrfGFEeRwyx8kgn7kWpRV3kU5
OnRCqc3EuX8Yw0rMUkAYtPUIeF/bbH4ijLL2zE+fBIkklNyQL4PIBMAF7wZbBaYZ
o6kAppNgXE9VpkmVZvKAF8wAAnV9WTt3Xq9L6r/DLfZ+2Fk3wWKv205KN/c3Dfvn
BvMt1iGmeuS94GVqYrau5gG99srU0kT6ZVCuhpvTW48=
`protect END_PROTECTED
