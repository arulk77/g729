`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCrWd2zgzF1cB9FBrEc+a0Tvq7FQzEnqMq2bxH7rd7Fc
6u4c1Y5xfavv62/bvnMkMv5VZZb8Dkvu278Lpoh9yIeD4oUYmHdPzFGqES3qOoAL
AMu14caDuHwLaIHP4E2BqfeQLoSxN5Ocpf7GnSLLKq0Z9Fkgc3IApi+AxoM0UXYA
oqfh4269qb87JUvd08f9HWSxXS6jJYth20XugMqNtZ4to9FrfsqNU8MOsgKprV/n
qnz3+GurcMbzWoE1b8uewnb7Xo+j7WI6wsBoh1wa0cLtoQOqYy7LFUrcQcOsfAn6
Jcxw0k+zYhS0LEPWDwfOEUJGK0z/wO73IhAtSGqxZ80i99SncDOGa5KtgtEmGuDm
9GzcR157JfWXvpkcfT6Ixhyj1oAUYJoi3FkkcytcM3xynXZU32JPeugjWSsDhFtY
OogKuwVsk3EZ40BplE5WTxcOydtlLbOXm7rHPq1+OQonX3kIzLtjStbgf7qgtwIA
C8eL/pIlM22o5sshNyXiHx72d6MG/9YTULvzx2fTbpOgumyQDoiWRsZ2iQlXM4Xw
eGgYVDc9RGWodR8NOmELVw==
`protect END_PROTECTED
