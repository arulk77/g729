`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
eW1CPupCOdEobnoTlA5dBkIWUJUa319N1gSMeSAkO48gHvoj75vc1uP++nOWbLEt
gqJS4f/vC2l/7spon87F1PWvSAQvg8PWbAm5KH7rKChH5pDQLGoI7Q8s8RemWrDA
Nwn4MUEjbTNBkGl9Pb6fJbTGi6Ikr15RKeBqHjJtQgnV6O+6wth2qwmisFmH8nGD
q0GSsWYud5+bUMnkKFl9olsgMzgoI6lb1bmrldGzTQu3GPr7DPaKLxsYTMYHdO3q
gUY1vi3XACKVFqeVxlLRHaxrKawxZYhx8XjzZTRj8CBBLkzBReRAoUzeJSId6UzF
9BqynvYg0YwuBrX+yAIZPEdbLklHFC3b5G0oPseQJnmmFn/D3q7knqzg9bL1w2df
j688OUw92G4Vvzc3ASugImwGZwtf4wQVB8dcUUVlsM8=
`protect END_PROTECTED
