`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48XXp2mnQ2NjJgXi3ZRHg7n4iW3W97yo/yWGcnuutPOw
/wS73BZh9MsDifhTEgHuGF55ZWn80El/P0WNPg+9nZY7sHZAe/UUTxyKosZhZN1P
1hBqCGRizF+1rvo0O+F693S5GnNoBdWOZNdi+PK3xCcXbmrT98iBBrd5UEUGVivZ
osE4N/RqrXqtHY3isknE4VjL8G0XclOy4ZGcCGai6tU=
`protect END_PROTECTED
