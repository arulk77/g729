`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
vrFX8dOSPAqbAN5lxhNXdHVCkRCy/oei5gL2UsW3A32b2ZgNbV8uYT899yPPPKfZ
eDnwd3KlFA4wseUJ4nOLBytFlXupkfbkMeKpbC9DbhiVWHUjbvt3Q8QDIUTBy+e+
V3818iscBMjkeTq7uf/JmH4tp2FNUSiZI5+xRvNwnlfBKmb6qzJtbfs5Tx/IA8VA
`protect END_PROTECTED
