`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
C/Ws+kSQLh8is9J7ZGRDzbhHAccKhdcl5Ze5napG07iqLrCx+n9TuRb/9FnjriwU
uza8DlZIJGpea182MVnDld4UVr8LJG+k7PptImu3OPJOU6P4OX47k0ZQtuRa8tUD
J+AnDphlEu2oau+UBxvTXgPlpDDUPD4wMR4NWnrKkfUyk5PZ/h6XCm+sF1n8UFBF
`protect END_PROTECTED
