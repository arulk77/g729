`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKypkN1UZwvyCJAvBg1Ztq6py767CPtHvb6Fn6P1jR13
CwhCicTRjQ3VzaQ9xwsrP3UN/bP+73yBOZV+P7eUfC4zIon9IkMYuC+zG5cGqgSP
uS4EPqt05prbrDOKaekMq+RBlBMAYXP8qprI/6jDcUB/0wx5hEWoocMMzHEN65GS
GFPa718nLA9ByltJUj9B5cScNPCjEW0Oq22xg55PfV035iDGSivCLeGpZkjOSvrY
DYyhy5PBQvgDN1AmuY+nG86D+LaQltOY1EO3CGAVS3chKokts96wdD0Z6pkkfHo3
VR0Wm6geAlKd5bWx5wcPhIDznfvfEwjjk84cJ9hExz5ocTqBIOCdzmLoijAm+JE5
SlnVfdoHXbLaxRhMUKS4M3mRnElv7nzTCcR07tuHJe9CWXcjg81qIJFQVOwevu+8
WIlMRUiWSaHpyKZrZGXiHuwjXMDcgSJuZbgYepp1D5r9KInPlBq2l/Ecj3F2pl+f
IvdMmrPaZJLb/3vHJ+JVf7jUAqoo6b3YFgeYFYAHnG+fJJM9V3lyail1AOURu1zm
6Hvfcv0SSWjgI/8xQ5WMaw==
`protect END_PROTECTED
