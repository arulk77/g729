`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C9pe/UYF5F0UEe53/n7kVBuTLRy20eNMvr4MJVHm1Txg
PGF9u6twCxyD312uW5IQCzqFCiMuqKIJ13SQhm4uIoYzjxGk5pFEM4FlZUdrF/LJ
i21rkOuYAKebs6RKd7n6atQfipebUpBMhd2AbOF92iHSKiTXnTe1QFEJxVjhBDK8
rmxIefWyUTdSmmPmkp50S6XefPAxJegbu40rXFc0DRgb8x7+n1910O8nb5cbXykU
6Eq4akZpBNnaSqXbUn0A83bb50UwXpcPdbRfpTgFTveTbEbvU5SgxjQpiFKP9HRr
83zPkhglCGwZpZBsaqErxPNeBG04r7IRzlypf2eOrzhQIhyEXO38lBu4z7F6T6Zx
yqeH0fFihbpxu95H6HgB9JZ80JoR2StJlfsKtq2RHvnzWrOz18h4tvrbn2zqM3jW
dyoxSZjfiLJgO7MRa9gpMeccv+vEKlWbEMQPu8tZuTz6E/R0OjGxPiPH7romvlRh
UpTIbb5JIXSUiMy2fZ6lbFoML1AJxIJyFFq5IY6zcpScjpuq5ePfZB0lnEPfR/T5
xGNJxzKzJUf/sW9Ski1aIByjNwFSedOAxNB1oFL7eHmcJC1a/aVrZzy34tKQPp1B
jI+teQUI/wrskE2ngdK4Bu/3sCZGU+i2b4lHFCXohUoUswbKCz40yWzt3SPxXBc7
QhdLzzY2Cc2SMiJ0ppZA64RaGe6PwC6f9X5oO3n7rTB1AWRLCbdUaRdIQ6LZaEIU
s/uuLpDZHNb+QJictuD5OkacrBL9QPKzoX4TCV94D3NlzPdpE1e4YxBG3Y78pFfZ
e4EEQn7bNm3uBnllJqoo8MAeVpGjQRFN2/8Oi//deISy0bbMmmCJu1Um0I4O/nCz
rZCbGa80sBCZpqPuN9++M8nOt7zTnAqA+eOb49IreIAz+UoQ5OrdApGmTdh4xFwV
tS8zPiVf/AIFCJDjwyjm8OE7o0/ZtRQmK1+AXDKuDxs6ss9CbaaNJXEI8eFdD3XF
CwKg0DTCgCV5ywheqF6tC2luo4tZXql3S5WJcQGBKsw44RR8R2dH9BvDCcfqqaiW
/XyVENrpMJFo7QX8r8369m15u/yqB5cXP9Gk+BBFuOE9itXdKq9X8voDmm4pKJRR
7dRyT1r7LoJczd2sS5qBBp5sstRqJyxmHTajGiRS7KCN7CNZX5QqnyKz2nhaJCFX
mMtr6q+AaubBDFVp1XNfC9XYVbWf/KDgIINDjToTr1LPLPnKGjvWNLwg6CLXtBEi
aw/uj9IzXFzly3F9uQxzlyGrMBTMNnaHEZABIrCX2HE295eg7e+EIA2UAyGOkpl2
ErCn9KhUxq/tyHCznWekOk27zdF8+vRRGRoJSQZZhUuUNE6Q71jBi2ejmR61aR89
a7+6TY77QZWrde2QrHBJdPTsthEK+tsYAUIkXA0Zkru9LVTxkL/13QKho5vsEZkA
DJbgYAH3o9iiIbZ97KhA/LuDTM6ten3MObDPU+CPPf/Hls9TSmnf+yBKiiYIZ+pM
Kr8f/f8CuI36+is0a4M083BZ0Y6sIczC4eOFQ4FuvjVVs7lWHNW5hyExCR4Kl0FM
Ccrs+zc2OllbXNkpG+Wbgghkr4/CuXtdn4zMX6CegSv9VJpCK6Eje4+3Sgs0lez5
S+G/vLGhdnmaXYjJVPS8d+Y2gFTms/byh1GSI+unZMEFyerNsHE/wVBZR0C7U4k4
yYgi6aJ3weaZq209HSg7qMEdJjiIFzWQPPfM2IjTEyzbTp7XqhnJcGac0m3InkG6
FIVIgqzx73qnrYXcjSvGaOnzscck2QbdORTmfz66MlEC7a/AULEG8T6n7lTg2Pgw
J7wqd8doIdE5Hl82htP8dpg5bGdE+JaARvZup/1q+nemSgUx/suMONZlZzZmgUZ7
IXr1YlQNyTxKDA5vRpHYGaZdyVNia+Ge86A3bIynjtFDYr37W7cskuox3YeSIALL
mCDhCRcvq2073QG02hk5pf2xqL6uEXqPHHpts9/ZoqBE4L/a/OjiYQUXrjWhZAw7
kvH47FM1mCcWH6W/+hpbBAMfc3SWKW+rftyE/mdkPAcDhX3l8W8YBT18kkqD5lXH
jKRxrWl3U3mz+4eUyySp5u+O3dYXo2U2BUe9wWdJfbTiKJJWxbnmp56gAm7CUA6y
cSxaiDzRtqaqe1TXzgUxJzoox4PtIYzqVfDx4hgoOpvVRHl4s8Ovvqk0su0sYn+H
OcQz0qeAac6ktyubTs3++EqkTbgorWMBVcfXDYtT+0FLB+1s6kmzqe1/KYe63G06
FxJXjeccMUVNyp6xzRcpvM8OTLfENQSOkDX8SfN5VVS5CwMZMrVwkuKF453vbayj
MyLBcvZHIsiV6RlJTtDvjjYceacInev2RUKaUs2Jsd4j5IZ9YGkc1F5eb2/k5To8
QfRq4hee0R0cqHfEe3EFn7r9dzw8uk/CUSluiOKIWGrK957TrBKDlst02hDSeigj
RUJsZcjfHY+ZLazcW9cKtDKmp+L2cLUzWUUjJlsZfq8nDRpeZj4401QsJL4ivSHO
DPbJ3E8Rwgo0US8f5/FaBi1vxU2VOHjmPql0yHE3HRFXSm3a53lRiYoe+56TMEuX
RM8cLJJHIATJl6u9v2gz+mkJXSktjTD4kBv2cpciGbQYxRSU7LsQzUQoUJm/z2YR
byVK7r1u1LgEBDvLAmQ0OexpjNH2eMUiKDMnhZOn2x3kEu71TfAWdVzLJqkPtbEY
Mh2DySzfHVU7rwKeIhcTKgI69rAYIz3asDlCF4wTLBzOhrneGbkCJ0cgr8PU2Dz2
rkvXOW9u3aKZyWbgrCKn0exEuBcmdRXtK7QyLIH9st/YoV6miNwiPSflGSLx970I
adiRLQDFBgdwIoExZFMvETMor9QZJXnZh5RnUzs72nHcCH0J17XTQt5/ySQ5K1fz
MOjNHdzU0hERRUuZOOS7cPAJsTuzZDcH8cWM6Is+UwS1t9E/ze/Yxz8RK15UUPRU
3RW2XIZNFoD/8xj5tEt+2r7GioUNHGVScmtSG1wDb1yW9gHj8hNgp0fBhBzVZyS1
fQ4MmWik0Ntvzj9pLC+h6DK8sfGqdJKRTaLm1peRfO1hHLug3Ctd23jgm/Ot/PcY
75JhTMzpJVoS2GqlvRkYk35jakQHGjBjqnjaDZvGofu3La8w1JfPlQ4Pmr8f/vSn
em4efzRMufIGjdgTB1+OOBb7/SqlJK2ETJmXpYQG5W1osR8WsFPI1yjKMX8sTkBW
b28h+4elh1DHAl2lxcGkjOQ+JlS3er5ojEOgsSjzA4S518iL/KEXS3umEGu+lcks
kCQ+F/xWIkWHyWc37QLplA==
`protect END_PROTECTED
