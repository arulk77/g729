`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8ScJF6CoWtsV3D/QklIpJiY7or48J47y6DgJs4j27A42/
3juaatTEnwi1ScahKBd6lxNmx4TwhEaI9Cmmo1lhhElFJFBb4Bki9icLwltCra2b
isJsIysxYIiGSXyFyzK3ecpaJVnuQFPpVgbtpEAhQlBq+gMPWZwcwJVlKsUBgFok
QqVUFQEUnZOpiaP59q0Hp0wbEO+xlbgr3dSKSWuWpG7qzmQTTDUEoYFBMKvHrrMl
PoGt8A69Nn3rTzOL6xh+c5h4e7E1oXR5OZCFqVV/8azhehJIHcR4a0JUkF65FDD0
6oWklZGk44tFOVTPsScJeSOV8tzPc5og4xDZbqdFO8RuigaGin/Zw14r/a1LrlZ0
oi3NsSJagNxY0OAUuTk+lz7tCn/X4YgxXAVCSKd7iYheOpNtJNCTECp0w2rh89ka
mybNZzJDXKhgOCOwK3UaVfX3fvhFOUo1LuO0MpjkumvWXW+K2St5EPMJOpiiGlcn
lRziWAMVJEdhm5DsBBj/CETAnom5cvn7UrlrOBi3KjH2Jp8URXbqjdVydqSfs+ed
NsDHh7X+ppIDwMNWjk+KH86XB6LlVe9O9EHAx/7SXfrZA5+pxLdwKoXAcUdOrSSL
Ps3AzWuZNnDlEX6NPXzlp4H0SYyfBMaxHUMVH2JLpn90Fq2EAgi923fwMfJ0i/l5
0lt/KdjTfVvX8bIU9eLkretEhjXiEyo327sIeqI3l98i36IRhAiUzTGfzp9DkKx4
jdn2jGslrXirJC2vDiHJUfg9+cheH1qVj3QGa44HLSRvG1JN91gCDH7QkLqits9d
7/W8FpxcpLNuGTuOUlmWK4fL3dalpdjZGTuiI6b147lU+Wgj9aHJCQTPNWoSqLs8
SeJ68dlaJ0KT5I6nJ5i6zqUdu3/viprg8N4+kqsPRnZNy5VEiIBHSb5A4h7/HYBg
uFwEAmGJIZa/I2APzpyZ5fe3614foXROJRFgXxynHDdB2SBqU9CRdCeFattEAFVD
YjKQB18KrCsVnQo4qAZi6ClgG9VhbKIfk4MPZS1sBvYyFWsWAB2S1GDkHw1KCW7+
s3etV3jIFh3YV+gwvcDW7A8rsF+fTiGKSFpuW1HeHFaUi5pquwY6XRD7kLmK32vr
8+3Bj8VoFWFvYrtpW9UDWgOy/rpLSMV+YG04I7QQus6OpbwWO3psfqt9ubNfCjHw
7qau2VwIkfBRIT7j5qX036Oq9MTQ6CsKZeCD/PEG6TB1JfHJoxVx7cXEKwKGl6oL
j5oVxjJlUG9o78gXzOuLPElVTNVEgcfI591NowF8V4Zaj3i9+3LWJHtkLu2K0vy8
v6dW/A5uVliYHW2ZJ91nuRtQV1RV9hVhnws+7PefWTsrAYLlFIcAM3mydki+o7JH
qgkhktT2ADLnGl4Al1RVEFwMHfyoMgRD9zsbeUi43NNcP7KUp/Hm92EjKfBF1Fo9
SL1mHUHOlBaquPJxpLNdIML13Nizn+ddM4ihKEhN2ZASbpOeCbCSkCJNmAMF3+MZ
3dvfrN26iL66Lkq4C8b45UXZBbRVtg4SLLuLVHvdx03tW8f687c9/v5SSP6J2DiR
CCe++EiXYkYHmRpie7wbeaOTF//ATELQnzsKz90o3exHri6O+NYazqADFEEbKlEh
rAVhOx2xaM8PBMwynPYsop1PyFl3LKLTfMe5ZIEzRaq0VNw87y4Nw1ZaB/ZwTTwa
CgZbzUSDOVLNQE/yXKTCkIwH//4VS2H/YPEnBlT/ri9RkEEUSOMJO5OED0XurmIw
+fzBjqPq4JI9X+9MuTVgkVmvQKYkfNWIy9vtsV1ZCZ1tyEPjhiiGH0lyWAmpR1di
kaGu5rNFcg/W+D/ntS+VZRXnT5aJphrKX2O1lX/C0pcroatAPCnZUnrDADBAHQK8
D0PzAlSvZedHzTSfv/0ctxLt4reeHue+dz2SrcVcO+5bIP1QNQ5zEZcqUC981Hrx
cf75PFvRIEvWUzmj1d32PfuzxLtE5Rs8y2ylmqc0GI12KxeKpNGKN5fXuIZGCu/G
CqAuOWm3u4UHmh8/hW5pFM1ufiSETw2CmsVFTcyJiWajRzmIne5yT8Mx+d9mefQr
ln+DwoLKQYAlpkcimICA84oyPITRmw24xDwVj5qMEflZ7lFzp/gli3tsyGywL4wD
baFYzkf8jC36LNm8ahZyed0HamYG2Uyp6F03n5Xnb3fAQ9UGgfFZ/6o+PUNsc4HS
1XMZUloIYHJusiJ/lQnc2WXsVNZhTrluS/lKsGMSKnge1NdoVSRGxhbjc1vCzEwu
XcKUiK6j964QRa8OBf9WSTh6zRQmY4JSHUMDzIakA1gcXg4TGffn3tI0x5DhILdc
u8XZOz97z6BtytqDthHZ0/UDK3EjsKAh5lVznXHjHfvRVmO6x+Tf4AXrCOGZP5v0
IodwNymDy/V945W9jBxd4fk2JfZqBAtAreTgJJaU1iW1T1eJmlBOZXMQ5dOr91cp
Fzr7cdeMER2cHwryV/m+FIYToPH9oTyYWtmHx6RxRtAb6yOYywIprYmCafKEAzrn
oEvfOMnAXg07QsOB9Qx1Ye1AVpR7kjiyqrVjU1tC85Ly41//r5mfQizHeT1iWrmb
lLbHeYL8Dx4KbX9E/F8CGLjM2ZLAItQeL7dVRJq+UNc/3nojl1UMJtrnkf0BvBq1
9guWdF0ssQDd4H+frgGrfx/i7v2f067l/9VvvIpGpk0Q7dCMR4QL47/RLF+3Oa57
njheIdrhb1k+5roejK3KyBnmL68Ybn65239bmZtkvaoVLXl20DIgvTds8F8U+Pnx
YgqNYdpdgz5ThwUKUWQYHtrY4M/L6YhwM2Q9IARjjezss7+5bU+Q5/e1xGBvLoPO
rIYKWia1k91EAE6WZtKcJ5R/U+oUAtVNfgzBIWY2VgL2hzHVmT5hFuEvVdndkdie
8mTd7a0oAF3yPqsvKMXQoRGeNNoX0aTioDP47s/vWB551n0DBfrop/NlNW5tQWyg
hYlpFikvdIDYF7/kAyOADtoreQLcmyDEtEA586JZ6sxL0HA4ZgpFFZjxvfSdvPXq
1uKQfgoPeiJwk3IOe2tbNqkKgMCXASYGE+UwGvZQwjjoyAkTAU2+vWlHGdDg/PXF
n9+qupO6L3KfNOmSRjNATNeXNcaN4XOc/uLctM4Jc7IDMO+wDuQAE4d0fB0+sLrs
QHQwM0cDsKFUmG636z5p8Q==
`protect END_PROTECTED
