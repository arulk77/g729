`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45s1yQvhUrp5DPLMP7zideCIDixn6nb7akDkC1UbHbk9
ZdO71eLewz1xky1SaQr0LA1Y3Q7badI+BCtgp6pqWqTZ5F9iH0t6JCS74NnsTltF
8eVI2L0M7AeqDHmLbWY9IQcBZkU/X54INqwiCCaj4ApCs3c9Z/NQYF7G09iUs+ag
AvJygVo7P9ZpZzrZkwGMyZVVw7DfwukzElXEwcqPi8dTbZXNgyYu6U8r/ksTW0+3
9WMsmjuyTNvkZa3meLYzje13lp8esh7SqiHPJoDfY1wsw1n1n+lU+rR3GlrIbuui
h3S/FOrITxAKC3cdqX7iiEAq40fAL3UyaACyLdl9RDpCPwIrHtPjI2aTVf9F60sX
509RuTbdBQ+ugsfAp56i+Q==
`protect END_PROTECTED
