`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aXnk6ucq0ol61P18NlRbVaxu56Zod1Dz4ggCiE7/eErr
Y38sF/uZxN/9drzRJlxmosV1aMRz+tinr6ureX7txxtzzRAumzSL12S4Wx6KtALE
ns2rRKipux5o33AQfUP4J+wAp4lMKOgZhpiE5oTTIH2RTPGJsZiIHquJxqbqtCPn
X+6Px0Oxr2CxDyWRAMYtmMQ9twNsFeIkZVfyz1gVv+iNOapDtbJHhcEs60juVW62
CtUj14lQyiV/DHuVfWT/pygA7vLOuC5j4l6XvhkJ9CpePzaDRL3T0PWnXbzpYRfN
ZgU+XC8vd0oAoUsuDlhXey6qSRdu9tusq2WRgfJ6O9tcCc3DIBOnnSX6Bje0f6zS
/LYb+xXASze7vAu/df/LxebAnFneriYIbshUwRWDAlJxrCWCVh3SzFZROkEEtt81
8xi7xYf3Db1ddwb9vuc7vV9Kq/IAzW5jDyrLlcmAUVtmyOcxMlximwreoB98J650
dfxvQfq3LyAFA83exv5D95GlFxgc8+xUR/2gSFnqgGzlrxhm8GCPh5f3c59RNxEV
CUnu1Q7fZQjozPaMZYdEu0aOwOuZEgzTk8vAQyJtQtpv6uuGLmuWeDmoDtbdfMR8
ZLZOBJTxahCahVxwe2NYpiXHQsPU6Z/oR9USvQfSfiV7B+KaKx/S8gHotj1JTQt1
EDJ5ezBqoy2Y5mU3yEaB/UqDZSAxRJAALSVSuuTwNCsXd4hv0LmheqcXvKNURWh3
MN+mOliUnYOuRtFEm1BeNKYZNskcAPRgUt3RLkT7Rt6jDi/WTMvArL862+SlIfQd
fOW2Ke2Q1yHaOWaID2OhfAopPfpXrngjirxeZMo8DMaUTcAtpM1zuMGoQ46gjYfQ
poAqacQmom/uFvKND1H8EC0kfdaTSm+2vLhfUfKpLAYOphVJkkdkrNscm7mwJ11M
d4A3ehXvCDfzpBuZsG6KR6a9BqzNkN0D1PwLTAYwe9Nns/job8mfCt/+uwKXFFcW
dt6KVNjVmFDGgD/TFyilZsDY7EBSGnvoee7ugZKhmJKA0iTOH0Xo24QO//aNyzxn
MGFdflxH2/RnjTHGJROK7jN5hfng/2QX/770UGqy8eepGESH/e7LvnH494l4r2Qz
b+fB1IyjFxv6WRaRFMwfzAyIccjYSeDr6A2fL7lEniHK6PxZVRoSPTN5jrqsiI4Y
TaXeRw2ht9XF8Hjm2uAMM54eXOAQZQNzZzCiyS1nOARLodCKeOBSM1QxlmKcSx1q
0iSxkP25vIjBDd4RmSmLUvvPpA8lHUq8CkJe4/JriFVTHUFcGLGOo4EuTD04RsS4
NzCS7iVan1kYni/q3onVSRT6Q7G5Fche9CAmVuvzMfUsWhYOWBLqYaiHe7b/QqBs
IsGpgHI3OneMWRAXf8iIJclVaRWzYeFV7ypSBFw8GanuRMrMdgYdpWqox1U+XdQ6
Ei6SXlHegiqZ+dFPJLqxNYi+HjLKlYuaKuyG2EjWGDhZyHouBCwRBjR+UM3kgr07
O4ooAzQdu0QgyMmjrjEV6Hz15wJd0YdI+Zuh8tNcqpYczM3E4SkYWVCeLHQKknF3
wtCFGc1nT6/m9mte4iszdOqdaK/YbrRY5Z9cC8wztHrNmVr1dRb8uLZG9pflSIxO
c18acenHDAwMPAORC9CGNrSXmTKw5Xwub3NX5loPhEilcctsw3sfEMASMDTs2dWn
9+3vAZtz3GLotOkbs53FAzXAnHAAFaz94jpx44J2plxwT/RIryf/V2Q8L/eE5TKC
cAnnu+X1z8dBWxberrwFfaEwzuU+0BthwFar7P6csJhN3GZSdh1IEbMeWOPrBPYL
2Vk6ovxcxYstdT3egr5tEVIEhEV3QSIST6LKveMEiCdm7QodcWbMGy9r/YEeiMLc
7PrLwtCRO9mtaxOVuyOXEsuvrHMBm9464csMnaZWPRZXmnYh1dZo/ZpgSYM2bXc2
mI57f/EY8OFPLcJNW1D1IM0CERwhKXRtoAMx+HxwBDE99PlI0MWnvU/2GdRZSBON
l83d6FCz7QhH0uGDKX/CE41eM8EE5Q7tkSq8qjHKoQoYDplLpBE5iSjv10khG1sa
ByE1aWsbeWIheQpIex0TyMjf46OY7xJX9y6LTHgCdnMU+olQv7E2OjUSYTGgaXqj
WwBNev8hbGmdX9z07mHq03/aeeY9JG/uhuf3DiCYiX64TS64frypOVS2zxxbE5CC
9Dc8/2d0Z4nzaj8cMHCUOHoXczvTv6D+NzZo8+Iyjsqw9WL7+kNpFvIdSifpYkk1
oYkOqJQccUPxDo92qjO5hQKN+1p7H0F/BiK5rBJ3ZQfYEN6j9mxGf61RHLuDLIB8
ibIUJbuh/LI3DVtt/UgIpsXzY8pIpM5lXapLpHlxI9hisA2711/M+GPIisog99AI
64WdJ14dt/ZkEBfBloH759zW8YnsHyF5c1rXtoMQKB8wJvFGOoNracR/TugcagRv
2CIKOGqLlSVVF/72YKTWz2xMhY2mgOkdxU6RGsvgYfBXT/6pI0jh42deo4D+ZEbg
G4LJ2Uiig1xUarHV5S+TrLoFxeFlzCCZQ6nNuHhrFu9wMhSF/srfLBLus2BpoHZs
6xpnBo8tRv2Cs/MFpbn9sGfnFsKqLX9GTG3qdEoHEvxciQBf4tBlCf6YyZpxQLGf
m/G2Ro5vjkmWMbUnzQQaHRoWjOpudisJWH4DKgMpCS5UzAQ89wPadJjxqhwyDwNT
nUHLRJvE2bRKwvDPU8OolEKoNqbPjzp0yfECpeJO0Wj5Q08QqGvqnV1HyXYGaxlS
hK8D9I9XCgLp00qj825TmLSSqK3n2N75xiTj3XtxA6i1JPiBm7VbAg9JucJfReQB
52EZ+EQY+CmOSPHRrBiL3izgf6wK8hNRkpkUyWqPC4vfKMj+uahtC1r4XorqZVGI
T1IoxzFjfCnHW7xz4hGPb3axnQaR5k2yyVBuxr5QZ0jGpJUknJvAkF5h0MoNUVRh
VPZaWJZaKgb29UK6seJzWpV5P8vHWSOHIrsuxOkbInDdwABtJy5YLKP3terSbjl5
ONCYF2QgC1N3dxjC8LzLFu9jYGTop2OI+ryObYf+tU3TLxvzXoZQvXjhOBbUEv2N
lSFM5P1SeTdFsO0BsB5qBprPZkRd7baVLy6DJ9kX3muU8IGr6fNqjgTyAMk7CpRA
W9c20tHSBRtEWAGhEsV66E1XqqfYnekbKJVsz/APxzQZ7/qWSjkvlocLReaNsWnl
APX8p/lMRWa2MY+KW7GwwCWtkykLXQ6aP+Sdm8zmPhL+EXIyXAhtKtDF8OGoqsvy
3B+6aqM3hOw+Qg53VTpTzbuwLTt9meVhkOrzRd/JaOlV8A/ZhWbEL0w6zxuoUxCS
6gIJ+HZuMivhRPJf7rjtMoReyZ1X6lplVB9uVQe928MvSdCjHfPh/6fLSMalnik8
sXbhDmPPmatsCcR8y0SBFdV+v3yobvO9BEE7Vjg4HuyDlAr21DSgU5om7fB1GFp5
02LYNzhvIrqK80XspSW6u+cnbzO/Lx8WLIFAN5XFWssUwBNNmlbNHA06wk/K8xt5
CnC83ie+mhNsUwBEPJiAkbhn/IffCPdN4BQX93+FFkSVdzFblpu7TyofG0lS+RYm
1jJPdyAj4z4LIlQS2CTbawmeI4Ul3eGPJNifUfS936W5wmA/QtcIIEbRqJKeELOM
K8Fxm5jgEcyMn3mtmnu59GOZh7bmuEfzLOe8DY48KKCE/ZW1xDE+5lm/7uYlx7/B
htSk5tOfoFoJ8F+MjnUs0Be8zNqdPtWsLgwWKft7/US2ZiCaQisNaquKL++rikSL
E+teKAjKQrisU2B6u4Wt4ftWIETCy250VxjeOKnnCcHkDPOyXa3Vi8ByUvoj454n
qXiUwLSzOZy9ABrtD8/R9PLR/cdtts8Hl3AMRGZtVUFv8tWqlRMeC0ojLmuYzKaD
WP6SIE2k7lHA53oboCNOZQxJj6wdWv7NrzVUbIQT+1XS81cDrPWMJmJBaAKU2aYa
sLgRKweJEVN8go345EQj2bRd4k+QNNvi64qcqMkDn1vmszS2Ozhrkp5u98knLMA+
A2FUtX66u2zpg05o2U9BtwiBAKQQEEQ0hEPriNbfAziovPMuLKhknjEQZKaukmMo
zHBx6OKz59x9uVchVWxVWRfOZyCtlCzCwev2o2kferbhR6OTJZ7jOTGItpiF67lA
8HM9eexnkB3cQr4GBM14vEpMr4A95uoKSZdmn6B4unzpzsSLGSIXF7F77plXSz4G
k4e8A0wC0idldxtQ6YJTIVADlLVqeD9qGqz2EiMqeXZ+zq2w1IHhZXNN8ZRlBLXx
NKQnCvmUitPhveVYX3Yz4ZXxZjdnNGe8L43Y3iRPkELfHOPLx30I3VbntfZ3YZJG
1P2BrCWXPO58UYQwkyg5W+ErfeJzlzJ+jqtEaavcfs1WlKxgE69I8K4NbAVl/vpq
XTXvOGX+TKZ9snpHVM3Uf2SeOcvAdLGXhasrWPvBkmxJV46d/kCfNuW8HsyMOmu1
PtLuFhwh/SbLKxQ8GthZNQDLsxsK3FkfrKy4F12r3Iyb1x8DEiW5Noxo9jf4c4yy
eTfgiUo0S4XL0U2sdpKSREDkx83mxU9awh1W4KDcM1nLdoir2+VeMTFEK9kuTPbb
ve2XU6cMEbOT9pdjwIuIZPxeOgA3MO4vTFYoaDLkslLVGyURXaQwKMlpHPeAlMde
tiQkR6cEkfyKMAY6b5DibBiTooIDrgzCWrY3iJode7MCD6dqGlV70/APrS5gpo5t
fZcTsPOjclbW2Y/LSJq3KKfatEZkbL71gYr2gDaOW/f31uGtirtKVRUoZIrJOjzL
6QmRVEt7ZiQlsE8Y5kFxbw6KQCI9YTgIpJNpAIQ/7pdIxrwALp/9YqWlDjeBgMIz
+whTmh3C5CU5iePdKy9OQ3ulhI3/wu02ztMDIuojzPWAyVhZ3Z9cuaLMlBMZC7JN
67okymyk78z2hHXu72zU1921s/S0pOTcAvWesXHQOAWAPRSg0GilkpPnyzRm0Njw
CEFZRmR+PjWnEf0s13Zig9Xpv6IjijWr0D2RhDIWX/Um9UfwS4NJhU6eOqANIhQJ
+YahL/CRSFVVHn3c28QshIhx2KXz8PsZlwYDJ3QL9RWXCxmEdBOKSeCNvmTxm4J8
cQyWAsCjwRpHrAdAf6n/+HduDWCTg+ZzRAYUSt1QRNi+KYGSAihF4+wsaNfpDMU0
5iwggYQjbV1nb5/mYux5xOXnhv1iOg+xh8q/6GLMl+hGS6jA2LZwoz5/GwpFda97
qjcyfIndIv1oJW1x77jT22PqXeixSuQeWy8j5NewLRqN8tizDwD5KcsYxs1wz/Ge
3ZWtJU1P4JevIBzdCVYFh9ECPbtlXr1vQXqSS8trbtzbyWK3BdNamU/XfQv1AXRs
4M24aPC1mE/Irx6X84cz6bd1WIK9AEJLd5+uc6OAbx3B2L2Hcui70vpRlOuqggpn
v+ogpGo1fgUaSYX3jwxOhR166x0rI113Ny2fGMLE8vBmmG1c+x5144mTXfdrsJUc
MolfBV+HR+uOjZWokW/iF/MZEav7ZwXX2JTS8AVX1RXZtkWxIy82trTHV1/n/wFA
XKSmGBRFkr+BCn7vA7oXpTAVNtM083bCGXop5Y+0v6sUs3Rc5LBEw2QBusH87vhN
KiqkaozHeOtGwNO4T1y5hQDcFjLx4LRLDXRz5HQzP6NOk4TjXjia+lwDb37oPPVk
ZP6mOs5yGECUsGOWnKO5m4fUVdfo90wHNO+TD4dhIrjGVwuBA3TJ9uZB1tCaiC0j
qH8RdOyNbVyGYjXVlr0TN1ESsn1NCJGQeBw0QSnjIdlAchBUlesTRYEfDXuigab7
0E+V8npEDcQnMsWI8KUQOUHZHWkhJMGs3IY+rV96r+Bu6l/yywd//Wl0HTlK8Q8Y
G0Ee7M4xHVlghHEuCrs4v77NUptPIQM79V3phZOS4EwU1XizXopQf8bksnDGIoGn
VpoLeXylkL95gMBXYV3C6gyis7PZxJGlIzhutRcSp8K8VuTgrTHi6pNSRSdPIdvk
CtS6kXKrpdmuXnBPrcMr6sz1AJLM7xCCZmsnVPOes01mu1hj6BPRBlTEM/xX4tIJ
tEi/QGazgspmZucc7v4dgqPkAxGx/YXiuSunhB1w8D0XKIMkwdslj6ZF0Drx9a0Z
MWz9xsWrzboRIbuo1/RUva9HBHjTBX0shykyWgTVMNUQg8k435S2fmZWL6yT0nHo
UMq1JwK9NZhDRdzMp+7wx+uvJUll8jzoXJzHgmmNeS5OeiUBniRiRqFdfZ3Z5ICD
8iWPAoPGjku28aZC7a7MR0oXFYSEkyeIE9Jkq/TZam8zX30I6IpuvPgs0u+je0e5
GjK3Wihlou0kZkallBJ0+s6cbM07dQGv743du2SiHlSvxHG0wm/piGhrcKNmArlo
ngFjA/x7+yB72k6zwkeIWslBlBO88w0VpnJDldLxX83Dl5uMFZO0Z3w6yCR8Ngvf
aAkLiSv1eGOCfeb0YjKfFmQs9KyPuR2yI0ZHPOushdj1wO1x09dANDDOHHbLQtIx
JUieMsHmWL2ZjRVeLBrj1/srfa/cqp5CdBN2tl6rJROi+pFN3OyQZ6BhkAp9HfVs
rkA3T4vVGOBSXOeJiaFeNxeFmJEdNx1RX4bZHKdry7oZz8LgAjZVZcjsHhh+Y63Y
Tt5HcgDbJEhsFSZDmkSU/DnDRmJIXnpxVtXgsDT/LniuzQjdH8gSKO7YIzfY4UdM
N9DTwyZgSEe4aO6W9hb6u8RGVoTjvkcgobte70veodcSm+w+LobGSLs41yN2MuId
kIjMwmZS1tdJA6/srsTXTGVe5JF7gR6+dzCKsZDKMVmjEanYJmj7t5VZ7frXnrlt
ZDCtgynBVXABqumxPRx4dnUvSNEvyNaGk8vCKJcf99yJC8TwBHBe8dTMDtOEp8Vn
+7Xfg1m8XUwYme4ZenVaegjP0CUEGD4MNFtmuMuAT4CB9EeEJM3f0U8AKmq6S8v0
vrQZERUCs/MNKjhurGSb63gGl4TDFbA30jJ887COXIFxOJZrvV7xJ826wKlmRjIS
yycOIkBBAYZG2Fdp2SPr2XcViZDIyDVUKSDhDgwmmvPwXuChrd6qATnI5kkW3WO8
sRVbEE3Cx2qzkQvpaYsVqkfe7LstpGdrSZJxK0SvoSi3DxskY73HDHz1zx6N/2j7
coPqDZv8MLyQRitGFrxRXMfvhy5tNt0fFBzS2Isikd3kPwuwDn/ebvP/rVhHQbew
IEYHc7DL1nYfl6k85fI61XL0P+WBVmmSZUQyx2QFBKJz/medczVHdHAniEGzjRio
12JrUzlflIDBPYb8Q98iXCZcNbXBbwBO6ABP3d3en3stX8TRByPb9atGjAyqo+iH
8+UniVKsOUfbw+fL5X9sJN2km2xYUQ86w9WrtYGAU0durRTWG67G0nMxD/VX0bVk
Xz40iozTlJnHE2GdEEMaxcWPuJlfUY9EbnKaK9se0KOQol/qzyRTUOR+WrtEVUSC
BYB8WTdGI37sB4AaChdhaWNy8zKB2EYHyW+GzuejBvHFpbeg7VQVlG66vUYvd4/V
CBN+ZDgXSl+OVRtgrqv1Wf5hmTMZM1wFoHGQFR6qjSF++j/oLuMFOpyAKy/vnCvP
ka8AJN/enSpq4Yitcy7zoLpJxo1e90nPib6YWe+swbD31F26YHd0fcccptSLAkYA
dhPEy8mqOz6QqxG/zguPC7ZGqupxxvJIW+1tPC/mZccmX1EkbSAnD35Mi51LJBif
cCXOTCO5jY4Jf9a/ziG4UcarPRhOBPlA1oAzx76urlCh1KE5wuEItAVbedRboFQn
1NgVUw6iz9w/E/P00M0a3WU6rKkZrNKgZPPGNRHskYsxPqrcD40AkxiEzB0s80lz
OEOhv3T7mXVY7OV/eWJ2EJ+ZEU1ASGeNvY4WVubGimlCt5u94tY+2aAt7xnksBzW
vFkW4MyyaiQFMY1UYhfklH90ygPsdxAd3r5361UKF/yj18khTbecfu3vigt8Fleh
sqqhQGCHTWzKfnDAUMxXZ5B/98x11QsXp7WUCDeE9H2HiojBzj0fdWk2q54kNZtA
LeHDPeKVCDjP1g9/7gncm6jOEBMw4qWVRVT/FH1GM+n135cQAYUj5rZqPtXLRhrv
yPOscbhfz95F0+QEJLtL2NBwSg23FxYuOmLjtKVlRgkAcN/Dt2ZE/u5D/BEWqyKp
x9W0hxcDjeDBX/OlR1UR4Vv38CzsVETUTJWP/1DlsS8rvF21oVVJdAYeUk2ku6UC
Ar+6gwOFeaZMxe/0vbufXpxoesqoHDzjIOx1EBwuT5Rt3ebrDH+Mrt4ihXodakBT
zPpxhckRBW8j+29Du/woZ/wsf/HRw9ViajY0R6J2a9pvwQaviWLfNToAp0zwOcUe
veC9w/cikKlZUACYW8mDH2lN6pzyi2esf9+60aQFcpZGB2neoA7ooXF7NVSpCHiQ
P7DbN36xP8wQpxAGU2a5PzryKz4V7Cdtv5eVMFpLjvPlLEuaspwanQsxKT10ZedU
Z0cUw2Mvbyn09potiFcHFMv9+UVjfJCbLBWLIGM1gqePPHv++K2iuD+W1TpnsPho
a/o5Kp5DJAFAYTqv3OnQICjUVQraevbjeyukJ8ZX2GM+2ml20dHCz56WWeZEYgcz
jUOjdAAG7PWFO9xDQfvR/LNFZ+UokuH+v08IdY7JEgk0qmjfbMBnsSAv82xjc3M3
ja9ruDCDBRHrQcK0TJrWyvqD7ru65QJv92zjRSzUhtX1qw/Vy9zFz6zyWUnp6Dnu
V3KdRB4fMuUxLV/akf9fQbh53hm09/TFOjM13YYlqbKdXt20ZtyftehqOUPgTQbh
otW0ljcHWD1Iv6lSF0eB4yPSeOa7eXe2gxzX5QxFB6oTuvdtIf/c9TgO9tAG+aMh
87rVjNUFJ2b4Z/DYBbd3aQ27Kuu4yO7g4trbGrF5zVNXtoCh2UM+idN1K8B1C663
HIGJzcS1WkJC95CmoJFxf5myYG3GQ+fuR0RwLwEOkbApJrIhtMcPUJDl61eCgOwQ
H+pfj1TF6ykGTm4y59jXtiZ8WwZMk/ZvbuSPXzHeNPR6n8do1em2mYSbrgwYQhTK
YyOQLOGoo0YnLLgEx05YSzGEYv0NqBQqBNfPTH2qYzKlETAHvMSAqbzZhYsZsNXL
2D0jney+iYRU60TyrOCn3YsX1A+vEXzwtu7Az06n0seBXXwat8pMzX3FD7DCqnkQ
YSwgb//+R43P03YENhuUONwxem2tpeGBq57W4s9z2BkYPD2gYngzGR0O8RvmDK2e
wBpreewdDJ+7FCTE4iaP3FKauFfwJ4c669aUd3y/yimvelYbKZzJO3eNAlDYkhxm
1Ik4UpFtuaBOWwodIzWCw9KI8A9gt/hnytRUMihFhtU5vPUtfH2mZtpe0gDzwcOy
ftDdJRbwbTafR57PBo0eGvaLT7KwpUipb1tT7Sy5MUVpqVhi0ngkD0bYCdc30PsO
5UiBAtG+FUo/8OHMvGjHQ/Eq45Ax4MObj96jbsdtG1g83A8w4AZlQYDydoPKUONS
CqOWGWS6T1+Cx8LS0VylqlMTi4z6Em2YTmWzouq+gbLtbFF4NjryongJayzfDi/R
rdgUApW/ro2U6Phi9Ti2je/kfFd6undiH/BZXMLSV9tlJ9Asr6O4OodD7uMhBTWA
XUQdYnrlLQPXwb0oxAG0hUS78/xhKtBmgoFdRP74GOPwNDtN8jPIDXjHs62xyh/X
qajKRtwmnjPMUyaQOIx2gVdb6qJi7/vLH9iJLDzPMC1gXLzuRINhATj+yfW/B1xJ
2LehjgqxMmvCQH9czEZdmKrckF9fq+EGjtFyNs6FdVP5NQw3lZKPpvJrhNplvQHI
hnWRjgZugO1oyzFyrkMVbGXSFkVjNkEVHEJAwcLG7v2ezQgXIDYDrabRCoNlF2lM
StMGw4njFM0pTgqLCUq9G63xubgYLNBnX61LmDdYswoEig3sYihWs6JNZA2SVlDo
YIxhIsXmI6v+6Xld+GT1f0G3kvj2VieYO0SplmprEvpc+Mp8JTFruleT/fkFz2b4
0Oal/K40UyXUOFMENxmlxaKwKtYhFkKrlMccl1GatPnBH97qVKU1UQ2wiOj22eBu
/0xJ/B6U4xfpnaiP19x9rns4QNTTjbCdsAMwD7aPjJcC7vO1yDgmVow1VrVt4u1K
tfdcrgM/do9RVtwN3D1QENSXO0ETPKTml8YYK9wAQrm/URSCNCIizjxHHNndXol6
zyPCZxVAW0Ev+sIrAj8a9X0vJddokw0/FczneGcFruxE5qELNHHGuzfgB9o29FTb
4CwDr7rEYkWE2YUXkE4MHlmtw4MQLksIVI0JkVfOU8e4BtjKOMdGS5OWHWSWkXY1
nnk5NtcfeeFuQHYEIq0I6Yu3FwcsHyseqEJqERIekNrDty02b4zVRhf4gNDMNrhM
WhcIwq5zN4+vkhVJUedc5l+S7xzmsXzXOyh7X+5sNUfGEVd/DXXjsqC/Rlo3zMn/
I19ZtYrwfv3nREjAk5bIFcYBZYQGPwXeS8vFK1ZH+HZUNo6OIXUS2VZU7juD/LVH
1JIHqKnWYQxfsKAjeODZFXpqT9xAAAiNPoOOqG/Gl72RAQX8aODZopNIJZwLPhh1
fh6HUAnLBW/csemkmS5iTC0fwx3jPuuAGoAJrctwUFZ7IY0MFuMqhimYoeW9fg2P
txUBcWd5grw8s3uzJxgMkkHTq0ZwavnGHJ0witE3Ql83xqybFs16GiMBEUzsjqBq
WCPit6jRccOrdQ09id2sNnl41fJsvmZuDOAZxObwhoxnqYCRHWG5kzG/D5MAJrbr
fj96RqkLjXO0GSFxPkZLtsGKAHl8v4DalDggwf0UOjICx+udSeNbEHER4yAT21U9
lyKLqB6rC3kBI8boupy4ayMSgHUmjY+Wc7R8+O3LSsXryud+2Rpdvs5s9NLT+2pz
/9mDniU0HtrJSFsT6KI7SXQ1wP6OM3UMNpUU3b+MMVuPhDBxUTL/zaf1GNiYMZyv
vmPGIi3x8qq/5HUVODdIaufhaI5LVeVZ/0hV7QMQ80GLbKjEhbUuCcZZGhvxJB0m
GStfq8tl9tTRY3RNGi+ZZQAVn8AcX8QinIWMoruw/CqxaI4M3MDGM2b8/oWpHKhy
qVU4pxlErXBit7FAdO7V1S1GR17Rkt8PVzm9SrOmS+uuCRBxOdDB2vHTV2BRj/uQ
JwW0O0+wqL0dvAVHa9ZQ1XzSJY7B9QPeEBz0VKc8qT8NFteg4DAzi3YcBHpmi1/Q
HYfQ+j8AbgCPxSHHek3+ilNZlK80aTDpNQFi7NWDVN78ta6zIwLQGW80QF9jamnj
Gs6d+7SqcvGnT+hhbssn5REW0TYEADIcKgXcu45eTe1JQnQF1QTNWA1ZOUi8dq5a
gva4hgLStfuwDaeko3fzLEvsOEEJQoh2pHheBj4oitQnuACTG9qd/8g94VcrgvWv
aSddwL6MseqQMsHD9v7IjSvMVUrqwqIarlIip7fPVg0sjHk2p8ng0XKBuucu5Zgx
JEHy41DSOgDthU4n7wmBLGKmRlFHj+Ln/Aisg/+LUdJNEp1Ymu39/BpMDsTLmjd9
v4gbtP3JDgi392FfDaQ5uiXZRtR3XqkJvJe9A/qnsQ5HmCHXPjS6QKqy+J87M4PO
nMW+Yp91y8xoufmXz5nHJ0xJ92gPvjmvwqA10/AVXdLKKK28q2FCUw0uMFr/rTsw
ZS8LXlom6es2X6TG2V84d68aoiso8dKxMvEYxdDA1l98+tscWFVxESg3ohTbr8Y4
qu0pcdBMng+AlcXkxnhwU3fZRbUonaldadDo4EygSwAxCHoenkHBLv4Z23jUdHCa
uKyImL9mV3eJ5b+gRz8/PMJsbyD3q2QmHjigzOCDmLx/o9dVuYT6B9f9CdHXjqEn
LRO3yHhxKLOJVRTjCwRqn+FJ6GMdieQIzs1GAPgDGHx99Sl3zln1Oh87BsfJ2YTN
u45urmS/DczjKTm+yVgresYj/i9wBhnTy+K6PNoWFEZMsuGEQXxwum90tD7wHJUv
ssfbXrz5PidOwKl6Ko6ZiLzzmOn7us0IUZ35ErAa94tf4/LK49hgGUbQKnsnFHYj
FP2SdQnJHiRFu4aKjKAy2FieGW9qgrkSNaBBp/UN5wbq4r9/OtawL/FIR/tcZ3uF
JRnvC5+Gm7h9yPjVXCuclaCCAfi/5uX9mKBoo5A6+DXjr81DKrL3bmsCdIUUGgNV
Hm2fFdUYuDf7c/U/ioYzTGKqSRD/XnY1zoNuPcEJk95jTIDZOldmywdTXbTDeDmR
HqitoaaUoYcODpl3VUcbcz7Q/H8AnuOG4P679AynA8C8sYn3Z1iTxivDFD/jCUth
sunMwhzGgDPdlUkAyD4WOTMhyFTcybuda/XKslsL9AabOxDTPDXJZQOSXKCh2/MU
E96ISsP9PzlnzzZjdLb/KtG2Kqsw67h6pyWxs1KUmJ/+MpldwJxBkhoPm2vpiG8R
fYP5hXNUON8rWeOKiBdZxuHe20kdpyM7VuKjCH/iu92dg6AJvRT0rlY+uTmGbH+L
lvPwgo89MkCWZAjGohIvnm5zpQYBoktv5f6NtO9dpxIn/MqxLRVGPq8gpL3NW0OY
GFWy4P6sMMe68yGO9jWM7F5BgQo4VYFFmhOhZ8c1vs7VYIAQn72zTJHJJOdTd6HC
4n6T1DxLDBXe2L5Qt/L3X3j9gy333N0x8Vz2/jySBmyuaEUQcUGNz/YprJOFSd2P
xZ7PQ3w89XrJNWfcuA0bBMNCL6J1OtLSc5nY1PCb3SFNP1/9/RQZPgz1wyk7JNxf
aflNfkFhoflmhcC+tWGEhWH3qfYX60D6ffXD90u/MW5J+t9bD9HWdZLEpXEDe4S4
uDm63aNRirlvfhhrrdtOEGzdCkNXyNoJN/Bo37+6HAWTXO5x2FcaLCKoj15Zrqa6
GKiRHFBjMAIcEaGELbPcDeAuFX3Jpm89YngbdxCLGzVhuG8aioDrlwZJUYRLICGQ
QxO0ckOKvADYkPBSw2368aRA9HLq/yy84h+1MJtnphWFrGu4MHX576h6q8B3e10u
aTZKzuE0ygt/Bw15uU9EnWKMBcd/J6lsA0ofoWoOM468vAKTiyghMfm1Y3u/loYs
KOdFOka8q4Lf3VH4hCTaxNfnfDnV9/xwdpVpcwUSXRse4WWoPMdw5z1o9jsyJOgL
cYFLJBUHgPePoDH58VCs4ZLOANHV6NXBxS9ZAJ8V5wDs0x4mRdkRVMVNXSJORLQX
iI1HeXY/zrdf/+xaPPNyA8SF/IdUFgbik/D3xDtjmkd+OtdYUByiyWEue2AG1G47
6GQTvxrIHt1TGdpJFdPcdCXa4knP8LZh6TRleeYpKtUlwMaILHDcgExD/SA7a4IO
kiKcIK2V9LqyFUAGkKW8dbNuRvKzzZ2XQ5IEZjYQHqJMGkt6F1Lpyirs1VzJBZgt
EvOHS/4GctCGtKQ8k7mozbriwdIH15tuTVPs8Sk120FEBPY81UGLcne5samh6KvN
EiuL1vDt8Wk/oaOSdLLSb1OcRsa6tlRcL/NSZX1D7QbALg8khrC5Nt2HOphjabKl
4f3Jyp/BakKOkTRx2U2tuTrrUIBXFOY1cVOh2DjEC+stdT4h+RL6KyfWE6JxRl7D
OZyQZR4O2F920/9xtRWcc7FU5dT5xYHAaO0rPJpV1gjgAFB9szcHDXxTXwNI86s0
YH/jjXpIjqvGpadzmKSrn/xTdu82xyVdgEi9fFfxKvE+BQ/FhjWTbFI5aCZ27DFJ
NxW+n4FuTB2Jh1SZsjO9m62dHSDnotDbO7+ZrFZQomfV5adJzWc7qV1QCNzPlBh+
oGvmNPb1qPJ8PeXGEvc6w4VnRT788NM8IeiWLmo0U+fe7sRQaMSPpFzz7KmkGUU+
0Ya+XTvNH4wziyM4sZUsvYP7mCdB8Qn+UwnQ2Hm8vT8NiK2Ojn6kJGUmLUArfJV1
6Qf2MIczHBE2QTUwX04IJVzWvzmwuKYSHe3Mwrpgi0DyPzX/UROKxwlpRQh+2MIA
tgJyamxACz/KJCNTCSmJNTpcG66NuK3/WIc/rI7NW5x1BKrbrTnMVbgqI634gmwy
r6ZYCnhQk5VOLSAmt1zgXaimIGyjD4zfgvr4tvHgSSXhgM+lhW8hQxCOtDDPMBYX
KteawX38sdnst66o2GFa3vfEykC5EWF/ecVJnrE7Ndkk89yD6+ibdTOnt5fDFZQf
PGP/mAWPHjvRR6ueAgUtZHOPHtYJhnQclapGu/N2TeVz9Z81SY0CfCAVnV8ogY6S
p/oVB7SkGImqjE0tagvCWcLbH3ctAWNczSxHPvw+6yRoMd1c72iNIr+5zO+dra8/
BvA4cMI1bUMSvqxwJCuYHW0UQeG7Sb7Rhy7/R43VhPTOVE4VdBYB/FdLUiNfJeVt
fnlETQdXrAGpu+fvdzL3Py8Di61cQobsL/PrbTXRClXUAiXK15ML61zJKmLmKlbc
CmIkAOX7pw31HtFvL2UpKEj3Bgxo9BiCzQfruftkGM6XTHja9NElLNc/pVxzgnmJ
4oQk6SZ8jdibB8Ujwiz/VLvb+aez4dSxnYjKGz5bx3fdghq9/+nOxW2UowxSfP2N
5jZYmOwaYw4c0rn9HPPyNpNZk765bFcv3rS1tr1eurirFrUXexgMec21zdlrX6+U
MgQgQzTdej+jjXuXIzwxojEFawmwBeBWBctE7QySr6QBrMA6X2h/PRMBkmO8T77A
SmgaioxE334vzJsBSF7ul8pHwYo3Dta14UpXmAcdqdlejiD4rqX2cruWhbyOV1fW
aeCcjbRXGGBvKooAO6CzSy4cGnUFQYMpehReHvry2kPtGhjFq+GvsS+/covoyem9
OLAHsS6ZXk48EY9hnHBuz/aomB01PAHRCndI97Y0VCqhR3b1xoaU1olDfZ+smGCP
q1ZQEpJ26SiDG881W1v+s+4z69XdDrXiezGUFhDyglvP9AemrqgKsJV04oReQg85
1erlte2cmk4PqtLKvSFFGpjdpPJ6lc7oS8loolKJUzWlr+ikg06mpWksVlH1vYki
ZT4Kj71TKQSRpst7uFAzmXAH4BzdveplOiY/MioaO167TeIYf8r/2KKy7RUuS6I8
Vos6dYC7MwCfUUqvTEvSRNAQ/MdDO13opxpp8M3kwkAYXWlwtMo5f2m9HijX7mcX
ukjVWPwKhVk34TpRaJGA7TI1h9JXp7tJWXkBa0MrW0EVjwRZ6NB3RZGB6w9/pqTK
WRRfMXCVCsEcxlvFgipuGRXAAptMT3KFifX+vK6h0a2ou/AsNpVgjYtQeaP4ti6W
WWZIg6127jDsH+4BwFtNyYmh8uOW7YDVRxV5QgvEyebGktiZj/gbBH7pbBikyR8C
dXXkEaD5Q4gPqAYtS1st/kxWNyUccFtew6bptJd+//jjxqwFJ/eBr1SykvGyEAcX
7grCqvtwHgwfe8YWHxQOXkbk12kPDTCq297rYUr6G0hN8wSIme5FywaIpGMmSFqS
mWPw3QgEuqVhdQWHekoueITVMINk83DGQ5EGUMhCWkE4IMWXcns3HjVXMNM1weDg
3unnhWHhwtZDxvEraeVoG5FEXVl50mLqtFKRMJw1Hfg9oQ5fTHflN88H7Dcfz2y0
amUmQJo+TI4HMVfq2mNtz6qIKD9mKhFtcI2B8lAKUEcdXzqtLF5D3ey+NivFM1ht
Rb8JC4iALC9JtDBTAGNAVaKfG2cd58NwRGVsfly8PDXdVmYFgUTm9vGg/1RAMV2w
HrFRUYSGrX/zx4SMgiQCNnMSS5uL1BW5AK/nypENt1tgAcYgF6hKyd3cYkT+Qvud
fHMQN7mgfM3ujxn8D9luBdoute40Dxhl6OBWAuzfDlVi25s5gmWubtlJpsqGsoLq
QnDNBazqPKE4O7vhlfGqBqKWrll4e3W0tPOtLXLiH9ttpjIihTRUqjqOuFRl5CLK
Ay2xCsvjNH8uaZpYOTblD5XZhX98YMY9LW4hYCJ9W9exDOuv4QtRe6NeQtQCVu1X
UFU7ZFYntrKzllwvwVP1WnUsP+Es6TYIG5wGxZzyBQjrno7m2i/wzjIbJXxOr+mX
6fRsXMW227N8GH854n2xstr2PSGj31F6lgqWq8ytft/TmnKm6lZtLndrLvc6GoQP
jpaoSl4FqOwWZxLARrKCIgmZ15hOGxLheKMNwK2bNpARe++0Dt3yMQ0xv04nmBo4
thVDeYQZ481/OVhmHQvnSDLav6agxdKin6Ar1Lp7AHjOmnRMxxx5UdNCCcJVHS4q
POtsGrP4id0DAvhdgOc/e0R2fseTq+xxWBE+P+cJZ4VE2h/PwUQSjtLvY+rruKvU
ZkwRMSU0Nyfbrai0aiDeme8WZngiysBgdynOSit6LNYrJnSOZf/ZTtZajBOJeMXa
tB6PV5J5qPp0iDkY/Yw3njRxlaF2180bgm+YbrzBjlR2IuTX7ubODFzuPT1Y6M3i
EOvpzWigS7S/DL8RqqhpyV6kw0yNzOIt+GcsOKm7nm2JtPw9EKv2xE0YPvox8MWi
jsrGr2al4uzV9LxJ8xBd5xXBsMnxU+qgsHj++ruEKrQyircjKfVqM/LXYVhjtepK
Nq7bwhkUBpWzBDsi7KsHYuGfoNMyciKzhKLMHjXbfa+sRsNhE5vf9uUNuB0yr4vx
YTbT3OAMbYPhA1YqW/ji/Nb41RMf6pAw8WB4vCXDVL9wrAtVu+qpVqbLU6D1QmsD
OU+0a2ZOZiaMXDPBGo9yFRW8nzdPlEohu5M1N5wtFqIJgh25zUnkBTJwahsIpLbm
KV0F1B0Pjhw+xhV/mbVDJWv6nLSLuZoIZ01dP3CWY6VkG7JKFasd0V/DMNOumt2H
3XIo8qOeF4Pa0s0P9l3Eh9RNwrfpeoYd7IcVVVJz+bADmKjn9aNcq2ibsku8DoXz
zhXXjcAcgC+7+si35zulXtx9i+wrkK3h73ogrCqcWpGO+RUTzK0U0hYNf8XLS3Ev
CUJQsbSCz0bFKlCQZ6WLhf5FaduMCvPhHxFF9EM8pIB/QA8UOTIfvdj9+GfKkPuv
za/+nSW9m0RWifCFZxkhGdwlUQtNArEkmhE+hp2vb4xassobT1cl8l1O5qfZKWeH
zYxJ6u/Op4AhOpSlczxpT8szKS3JsApw9XzOSDsMxdmVPJQEIgnftNJpY9/2bhks
Ws8oko81MlONEztlx2FHA+Hlt6ivi37Anth4J8HfEnQ60eNJcfJczEplX2Nx/Wno
LYiGYLiqETVKIZRQcKxykBQmp2kpdVRrWwKzfYdE5ps9muMjlIDa3Yk36610wYAN
D5PYvDE3cjZoSHksG02RQ0Dc3VBC5oBbVcE1uDF49bPN8pnLIPpA+l7bLIrCemvu
gbH5CmPy7wF1DZb2wMksp+3COzS8q7DUa+97Vi1ZhfXyl/e+TsOzGjs41/quzTGP
BUBCc7Dhu/tEfM8Kx2JjvMiRFOx/jFr3gXQEM6rvpmQTy2jl8k3CZpjcKmswPtLW
pAH/ZlVOVtLjM06kY1oVTDawMgGI/hHq9oJ++eG6tcHf1i2gXxD7CvVJYTd7+1EQ
CuTTMJ3X3SGM8mUwko+VQINyH4tOJtG+fjN+gIibEyw3ss0fyJY+drkqqyKmY3kR
`protect END_PROTECTED
