`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QNw40IqJrFvY2E8HYWz+j469YXKjSEDr2DNQK5u9zdw7CzmuQMoIF6YtveLDLQfa
ioYAWQFNQ9qwsjV/VOV/I5XXnSGkaxRASQBO0E76hufrJJdfvO9uf0+gIwDHWr1Q
vwn2lbDVUq1Z8H56/dlaVkp2lC2ISzotwZ+HK0FiDWOpZYCzny5/G4dX2J47SKD6
`protect END_PROTECTED
