`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
MpZh0w+P2LA0ouQCxsdoTjm84yzoSV6M+Ww51PgTyLW4E9Q+0IYLi8vAvMnajyT6
A4sg4n/aKv4YN2OEsfB4ngT/yjRi2YYZxRBcLfoghrYfr4UXzt76V02tGFQcBKFs
tC2D/rtqBwkzF5S6jABN3C+h4jengUyC+csTtqAjzx4YEgl5d1w2Kl92sCh3KQwp
MYnVjgKqD4EyClN5p4elLeEAPM8rLKsddNWeqB+oZ5HGgjlTayUFpBodyeSHoYAK
u8O4Y/lWxQmGfkxI/No96tbLY0DSzqbnZP4/CvkuWxKONORTZrbeodq3aO5c88GQ
3K/T1tibgRwGb1B31tmTJGnY+1+1JbvL8GRuzEjujZJvxWCWi4BIQLGdLeJIqRv4
KF4yiQKWwg9c081vqDj/N0loQA7TOZZvK/g0FkfZygo=
`protect END_PROTECTED
