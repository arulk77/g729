`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
lwET9c69zFFncHpv9aM++gqSCfjCkwa6PCQP7lzN5FNycVsMRAo//DqzBPIcd8/j
uVrgQtH2csn5mRLKSKy7HBoD8eGDietJokbOZBRgDhHcsqxLnS1ckiVDTYm2NfaM
PzytHlVz2NeXkvCjbAawTWu7m2t5Wj5eREkFCVhNcD4Gsf932IVi+iM84BoV0fjX
/VJ8VaVQr4aXSPYoR4YvugPu7IRA8zaF/KjQbsT0JGKsreFGaPAC63m1yF/GD88y
ydKCNQBubZ+WxqC98CsB+A1oivMfaF0WYpV6PW83+DuvfmVqUIC67TEL9WrYBCqi
5dchSBAUQsBqArrCbpAA5Cdra7dZsCvMEidAihHXJKnpoZpyR+9bryUwKZnj71zA
Z3IgJ97W3aTbQboWkfKpWSTWo19a1da1OpDuT57FK7ryznzWqA6e8ddpH2+xXU7r
8IMrMPs6JCyHagsjFv8tLuCly/2Gc9s5Aed0+J6d5OaYaNkuNbgxqkv+O4jRgP1f
j3HNULzrKoV5JNqEMnwmfyrzuDL/Mg7+PzPUwanceKK8/bXgKh+dONI663IlBQYJ
M86Hbm0IAjQefQwXJkCs2YHLAdo4QXBYABvZc1xEMjM840noJWVDzhSq86kyjxXc
50DZq1uh7Ud+NOB1OCfXAH310FC/1A1162B5+IuM6Rwe+i2ScudWCzZc/nqlkLyh
B5WFgeR2u8gBK9+CQkidCz2LgnEQ+cRbLa1ymsGm80rVn4RBYBIw5TCHwe+NNp77
`protect END_PROTECTED
