`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDkaVJq5W7s3t3iUFzHoZQNtZGJfRcPRDltor+N3aFZc
Qgi5O1DaD301mEKHdIuggDpO+qVHMmEbiDuv880b/Sk8+vvyYCyClMbm6k6NKofx
740+NZGudvpcg4A3z/86z761rO/dIWqAYWbrFnnXyLu3XnjhpdJZkidurR5SmjNe
c/f9vj9IbGpZtC7HAh4y+TfQM8gP1bVjCSTMFYTfN/c2UO0BpGZazeFgH0Z6VbdD
`protect END_PROTECTED
