`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
VN3cZiJB9f6xREOOK65F2rvwUy6OjgnMsjH9gEeyFQJy1JBVIMIJTmpuefr1TPo/
N4uGySpkOCERWvCXB1ADYniOL36gEGJ/W+iaLf1ane/jm7fd8zUyRER0Oo/USpwc
UFt1NgNxClYJO+e+qaoc6W3wJKsKmNBoX0r3Vy57t8qj91IkSKzbyOuIu8jLWAlU
alIjIjqMcywcuXOISyPLsGEMHcS0uor2AKsYGjdomJq68+CIE0obaKFNIV6RJeGj
/f+9rfCyqgaGs02LpzUyV5Qp+2G4v+cgl6n2bNwa3/W/ga1ZpYw8j9iGaWWH/ZZz
1n+pLUiI+rvVxAzJdDVTpg==
`protect END_PROTECTED
