`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41u5qOW731WtVemQPrqcn9/VTgFyDNRSXIVHLjP9Onb+
OYzCOjA9W6N49MEWBnSlS9+jZ0Iv4OmNwALYVsbU9/ktYJkKasHYOMGIWegRUvqW
xuSXjvC0pYlOXoyosbIIOLrVvh8SMK34kj0PM0F9aJ/v+fhsQUXKhyPvBa6JUUtj
d85zu7JhuRMc56QqivKVIyBtDOXhyWTP2iEllhdE7KSYko1vVXspEGkmbvQEj03H
No1GT5dJ75RqmQ5hNZbTET1qxLoYKk9d6tvjF1pkYLLolh653I/mWVToCtZosA/f
SNYldS4gYHeInsTcfv+StQ==
`protect END_PROTECTED
