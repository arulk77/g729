`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJAadpaibfqPZTfXCsmto/0diIynuXHNBFJJperAou4s
Q17OBvJXn1Cmep7sUt/TpU+Mb6Zf8iSxJvTFaPUF9O7Okvez9rRB9vw4wYrwvbeo
rJBlQZMU10mfqKJhutjMf+Mcjb9YpM+MmDOOwXCUBTI154pwvFC0XBRAep3oxDQI
+GUMoMZn8WFQpLPQ6MhEOrXC6011ivq87obyERG8PcBkenlMU2wF9lhP/0l0EViV
uVToeEq+afl3uOiV43s9oBoIrlvGVaaP0jPZFA7kYVsV+cpymzvlFYwlaZh5ULk7
nnUzNq1N0zRgZqtSrbQCkg==
`protect END_PROTECTED
