`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Nhmw9HTab23zWAUA5Vkul7Acd7MlCtJDiil9u7j8l1Y08zSCxt/m3778sGaZ4D8m
5rGTipeFtPG1SzGn29sYiouKCnAPuzV1j/mum5gfWJ0dpUqdpgmZ5G+twUoB62Iy
jUvLqUaa+hJeIV6oH2PkYCk3HbgsHTXC5SgTkLgHkyJH5lJsSb+zDbgwV9oyX9+o
wJU1kWoyiURUcsk6vj2S7hFEfKD19LCQ5hUA9uDzwaY+jwr+xgvZUyXbYRCd5FRD
UWt/qs++DakQBrXvuBKVjSvMojBcYw4gGMef/5OZnsU=
`protect END_PROTECTED
