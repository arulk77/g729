`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK7JL1wNbIyRzp8q2Lk07mVX6r1cVi82To2lAjQscVCt
lK4dDTpM33j5AQM4FKiEWKs3opr7wFlZsUeWRrAemZcjljxYUR6Oms4LbmzxLmL4
yfptunL2yW3MEfyaDjZP2hkm4XZz5Q/sdGvYby4AcqgYhMoD95j9fx6nqtTTroDj
sDbs+1uKTo2qruQJ1200DlhKEYG7RKQ5LpVKw1WKSm7PYSLfT708p55644EW1qeb
WFrIHVXqi5la+uIk4SP296Z3q1UhEb5qkL+8GoiXOQ0b+LteUdFcCbiyO8IjXL/Y
71BMe3HKMJNZDBsQjGUeKFUTtHEwl6E4KtrGo5aBHVa4zTsZ8QaJgRXrbBgtnDZ+
hdc8ZjA3LkwXtKcEWelqiw==
`protect END_PROTECTED
