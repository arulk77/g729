`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBCE9QXCYfqQfqRz1Ij4XaDOOm0jiJQOEaOKzEIk8/7R
Ix6Lt7qq5y85UO4LsOqtTqYbjr6mYBNO0Ej04SJIlMUFrUMh/XBK0ezV73kmsPkk
OKP5Gx0+TvPdOmfph4fwZH25mkq7F1DReXrBDwUp8ArRWPpYAyQm34yH8rsg8hvH
LiAkd/s5xvQ8mvUxpUHhUY2caVhkaOOnn5Q+uAnvGUlUUqU7WFQF1AHiF0pmKviK
nai/PXBE7GmOTo4QpSExM5f05jZUQDJh+wcx3eGAGgtJKXGy+ifeQT9WEsMlFUb4
+qKeVsUx2ZAeDGR72tmdocJ8G2+yy0k0BWQUs0IBpK18UBwyoKsweriwO4Wf6+CX
f4OdYxV7SGJOetp2TBdf6Q==
`protect END_PROTECTED
