`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu432hW4JLsdH3bYgTVRXl85HDgnihLzux+LfJA10wac8t
6AZK/aI0QKs1Zh1hHIuyYWSg4NZZHg0RTC++uSxYQbc+AZW4R6MYKv73Nu+gU2OP
Frjgc843D7l8+5iM2jEDWZ+yupbPWsIiF6VT8hoOzeg=
`protect END_PROTECTED
