`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
7SLQxI8JNdGYM9/1f4FQYzr8DzNWPqSxO1sjVtkV5vHMw5+8GoYzDMpgYzEflaC2
E/nb5NbH+z2yB5BXg72pgfohbZn+p47nUr8Vb+vAkxSYv5rcGPrY6ItULljHwGup
qUsFZIiuQ0R9kLNjEYNEn2WE4YTISK15UENyUBFgexCfmBdu6hjv66W9mI2CPFsb
`protect END_PROTECTED
