`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFRZbBE99qWXdK0GvKTrM//FMBr+gQ7xVhP9R2qnJVin
Kf/J/lfn3mkRFk7TrRr9iNIeZM2Y1fmWz6chP3SD8qUn7+wBu0RmtUX5MK+s93Ev
Xdm+q7SPrOhOf3gbCjf4ItJX788/0tL5pyeKYTfChJQ+2oZDEH6FDD2n14lVxXaL
`protect END_PROTECTED
