`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKDBABJAEN9xdhXoXN1PsWXCWmFB77odTtphEZAy0w3R
ldfLjak+2zlxRkZ0plLHx7S4kOL9LDBcytrXnM6vo15aNIXIp3TX15a+4A2xCFeY
lorJaQ1FBAmWI6ygTLJtsY6xzZgsaZU9scyDg6cjFHW+NSFwepvJZ+n/LySmK5ua
iU7TyVMEmqOHlP1YNOMWt/PoawyVNb6lG9teofHyanDOgUbZZ5oRmZRlj8N8JUIM
fejNn2Mtek20gc2zX7UoZ+H7TQXozV8haUNALAAdgCuNgt82C9bAUE4T9tYNqq87
1nCGQfF0lYPw+lGwJvEySyXqnB5YMKNnz8ZjirZ7y3/NVpAas4IjzPlrvOCA1y8N
QblYtBkuiBLbHRpAVHO91KC55M4JystmmcF5uAEOcvzpTV91YJGf47FKpSn5tSy4
soWkxQ27947ev33yRCT/Bh7KRHlHQ6pDr18CEh+gw3YXZdloT+LFPS/WgEiTkask
juAljIpQZU3+F1hXhn9OLFw5WkHDGiUmvZ5WgtCQnQYMP9MkpuIL2Lm/dPWgpazU
8XEGCd925R9l3/Rh6wlFyOaxXO9Z51n27oargnJYZs4kz4teIJ6rYD9DroU0YPzV
`protect END_PROTECTED
