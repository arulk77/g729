`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
hs42QsUaxmcjFnvUJRkx8mcBeBL04Hk9HvwQiHpezdTL6L0/b3b4t+1EozpQho1d
4H5llwlE9TLhM+5/0HTHDXjACfgfEtzxAdJhYeA+5NeL6m0rtuKHttz3iuC52qte
WzgRYjcajYcvOzz86eHyR4AYwjpD7hK9q/8eYQ17pbr3+FKSRR+Y626KhNtuRyT6
Q7e5NZLkCys2S8pTIXFn5mpYZgNYhEEXwWWeIyyR0ue/BFdOOMCJt2GzYc4F7Skp
bEWNxhUaqmO+B0hAgw4EQNDPIWeiCJWXJRTvOLaIIfhnV0em5iZLGtEzcD/D5QvN
gXkPY4JqXAtU68vRZvCWhdnJV/HGfvS4cgG31j0OwdqE/wbuA581zyNQd1dwxGcl
y6WxmUA2GmfJeMXczHc9Xsetl8W3x1mXZqLBmGld5XJ6gFEjJvz7PEnbutbDGYnv
vXxhsJ/P7OZJEzRSGOMoJGOqSO1O2DYWebgrq01pJy2waxeY47SzzFkyglDYU39B
lOsUjuiLgcW4zqvCHLNhdA==
`protect END_PROTECTED
