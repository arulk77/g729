`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
tkvjUvSGsoxJYpv26QTt6FbuMlwvy4wBCxSxpEGoj4fFeraKTiBq8Jm4QMA0w6Eu
t7NmXRX/4NIEIaq9Bdz0wCxrNVqSUbwohyagaz/3ET+aXFnYgOpqG0uKrgL51NAs
i7+XDH9O7SRkWSju5UCTIsoJN+M+6cxkaQi0uP4gmeaAEb/cwqyYnQb1G05EerUq
s9u2rgHvtRAra5DiIk/vPg4C++85Zar8Kb/1Kchs6rT50W6GsEjin7BRxqxhh0vD
VAOvTZ3ieZiQWVUCiLVXGbScKpnHTob+mEDz0PQJthjVwA3DFn2WuIoCWN8PiB7U
Ls3TIYMF1qnS4Ws9OOy/C0sKMkCpaVqv6yybVWcshVbMYrOZcCWYzck8Qq0LapN2
fWhQh+A+fj4HbterBC6vO4OkDKvAG1mpSp39PQvBw7bIEKLf06srCm7LbZXsesxr
qFlUxLv+rJxAN15hv3t+i+gtLc8fi4gjihuaQTsDdo6u0dGnWI8zGcrfzIKAipyK
fbpb7kClaZ+YKZKDxL00EojLcPtODV9SdDpS8lGn+uBhmztscsQZBidZpL2wICRf
z4HzStQt67EXpyCUeNSOag2SRcPg3YPB6u0xQ2GfPmXriQo/y+j9pnGYJjpVGn7q
OqqG1k4oWLUNZGPxzGHD27TqU9zvGVRZce7a250BqXJmSWN2igePW8GN/DZGhdvA
sTyBDQFb0UprNnAuL9fbkskoH2wgrYAe2GADcZ/wEQly02MdSdZ2ZPkYJ816bmkH
xlldQibGo4QF5BFbsjK80EJ4hmc807nJX4PafjkyuqLZLTHrQXc8MZPJuDjoYrN8
H2+1IOQ6Wu58/1/iciffW7Mj+ZYaJBg9WJrUnsGjUNKDrAwFFXYzDsCrrLb6ya5C
`protect END_PROTECTED
