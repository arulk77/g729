`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF1BUn4lk13Efx7BogQ4nCyUDCzsEW84V/bUUu8P8VX7
SaxjnzDMtJ2bVpnovDv3KpdbdAVFW6G/daMu6ai5wnaQJlBgYgkvFK6FGYrcuVYc
BVpGUgD6u8OgWkbLokerwsWCLbHwRgyW+ExHatXNvOKdGt7FQybgG7YlCiZYEm55
+JvCH5BpptrV+kpFFLY3gHY85yZsY7Mw+FJho2i2nvPFHYuTiKT+7ElckkgH1ulp
aniDAzkHtczAJ2ieq/6GEK5stXzxbatEVsz/vmcBEdB2X8M7UB45e2ZD+IU9eSmk
zVZ1iolpqqBsb2Lm+Hrh32fNMwhTVweanbe0sei9HM9lxUaW/qmprRLGgGU3iwJ9
`protect END_PROTECTED
