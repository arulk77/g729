`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47xhcClvSaA/coOgOHL9MiYEWeIU/RvTMSJGRQbFVZYV
37WT3hmA+NAdaY2AxnTPDhhi3SAvUjwibJjXn7xy8yDArYfbIS/z1u60c4R3fpAM
m5Wm2tVK3lNu3u4EVeWxP7Zy/TFOrZ+3wbFYFZwIbS57onzqMyjKuT472cjpsjYJ
vW8pOfnGgN4s8Net/LOmeCEV2Sjfjl30VEKXkaLbY/IKOIe8LcTPFlpWkqO36WxR
VZf9PXWCat0YdMTZIflqsFvceyJzghzqVwjReYFxdnAuciv3nSYg/SXOkiTgYRh+
AUpmSPU34ueGN8rIWSEAVg==
`protect END_PROTECTED
