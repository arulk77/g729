`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJHNKXet0jQSqHqWgjSMMojgWMO+jsiY5INtBfUrpD6U
s39x/YOrwtpmnYGvnaCQWD6iHtkrwRPGRAXMGI5qd5c4dFr0z7uIqKbqKPY0xFnY
ehSi0du+8VosD6arukXVV0OWm0XeUQUEfuCCJtTcqHnfm1V43w8QFYVrJ+wahFpS
HaXcOGUW9qKT2uDuTUGdON4pZZSN0f45+qkvOJdtQH8DXEZLiq7CkgkWaFCBiP30
B1/L/jW4YOFn+0OIkCmxirqo+So9xqaU6z+oNJzpScZQcYr1lOQHgYqpfRkUe7Im
6mkxPFKhcOMZ3hqsqhmrHU1ouzxwmBh+Z050q2Ibtxpuzi4oAFz3XaruMcZS5tNB
/HfGHf3/XRAnVyUESJwrNEc2XsnUOA1M7Ngx6Ds9ceS1kjCTuRrrhYdN4pT0ixOu
E9iqVUQwQcUtvk1UPEBetWZ8AdDhxkivOFAhZ+kXqfZtBC+mPEkiYWa8HAGCm8P6
O60FqfP2k9L2lA00i3wVrBQpxUANZSRMXRlZeriA8dnBzs/Ftc1M4w6EhcmH6AvR
AWuWPMYI6kivlhNEkc00pzDkrAihps+McP/RkL+1v30qmz/cRmc3EqdTHnZmFy+p
sn6tHpu5RGuVH+kjbuM2fQ==
`protect END_PROTECTED
