`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLSDK0/TvEbeyxmTqfopLb1h9Vqgw0g07w76sjSNK6t9
T7N8ralMmEV6FIsX+wmhDbwOCFXe06CFFYCIQDR4RfejDcLbHrVa/ZLtNUPJzCCy
AMl5to8bdVY5ffzfM+4g7HLzEDl2DpQ1xkI24IXe+njAEH8DK24kwRblXwvXwiRJ
4tpOFWdxqkA1oqiVOmBboQ==
`protect END_PROTECTED
