`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
qCT94RUIry108LmOerL4TPDq8XQvuqKUnzrUTVLEgtK7ILFCYK4toAiVNden7goD
5JncppagYO18+Ip8mQLd+tP/2BGImEWsd6Xv6uHbF5IG1QYsrTBQdHEPtDsu5m9R
EJGBe7tiulaPRp5MXrKDJv1SRCVhKeTSoVxVELHIfQw63mM5cfS26HD2dhEAeX4/
5HM2sACThcECkyPNf/JufHDlIwgaSFwORGWLyOLmuVT9V2kX9LxN0ilb4Hl0OnN3
K6rc/McbhBDpxT1MkHjV5AWzidfweFjuJ1cY6wGNuhSZiOacVgVxRp1FP1Hk2F1B
WyEXbcCyHmjpyhLBisyTSuu16wLDygw+uAJXFNu0cXKx9GZ6NODnMst7U3GnFJ1Z
x5ighFuh2yrCzTo3JWkte9bLbtd+4DmTyNzh1ldwwRrhLvgOVVF2+4LbVpdmI6vn
Y/SoeEL5ZgZKEy1bwt/5eWyENY9hbB2NbV3UUYc8jUGnUavEdLi4eNyTiMIv8SKM
5J9kvcFWkEYMKJNamrq0/DzhJ0V6R+XLPTSej6IlInf5dgymAE1UJq+3MdD8uyRy
JFjc+i249w9sQ2J+kiR69Ca8P6RUCovSQ+IlKTHo7Rb8gJqjJ848vF1uRXrIWYjo
ICET6NLQY+fF8P5MvbBvgnfNHOCW71kErhNzh3yvqt4B1t+24xXmjYuLqqds7vL/
nk+B+upN9dtH0jLCuuQoi+bH/hPPOYg2ObzBtLjcM313v1aN0GtScR+ySjXY/7BK
U9nJ0XFhxx8tjtxzXYka7VnfJLpWEZC2NQua1Q1eLBPE+Jwl2qfynizgVw51ghwD
fPT3mj87fQ7nHw+MPjPTVIV5yHDllLkq8PsqKDMGTV6lVjY4gzsWrzpvfteTgfZQ
e3W3uLt84PTB/5acFG2xxd9WsvVbVG8SmlIh6jfFhxrYQTfgda5NByC5khyHIrcq
eqhN2VkSbOWkAfGoA0+dLCNVsc4CItvTAC1UCyM7ImS9kG2w3f5aoxM3Ib5KUqud
hYrxya1ixIbwp6W0SnfT980OkZqGdd1PNhrdj9pIMVbn3k6z3wXEr3vIUGg2mg4o
hIpT+EidHX46EqTErr18oLEzSllJRP2Rydu+KH38Lbn7UTJKf+EmQYUi/OA2B41W
G3ANpazZg//Y6iz+VsQ9JAg//QxjxUgVmU/K49H8dKlI3afDXJsyzCOLtIxf74Pj
khZGRCW3GcwLQfnaFJ3+OHEUaiXF8XWbtLmODuZRz5qfkYidpwIzCAs8U9ezoY9m
X4cizjQqWR7GbCv8OWQo/JVp2d490wTbm8lWmXD886S3RTeLHt2vh0a02GmLyKpC
11mA1JCvIj46Z1gWDs5a9qMmIhcsBZl9deUUKXv7itGzuN/kM8diwzu1n3fek26C
rnmeRD6Ly+T/C/nlLFglA53HIoFGWy+MMo+po+udq9m2q7TcVaQEdBLZs1PGjN12
7YHd21oZ+/j/3qEl6HPTmKQ48wmdbjiHuRRZ5C5qyBAA9xRZggrzkdozbXkwO3dp
tz4wu9DchoKDpp14d53y5Dg0G37z+M3EciXntlqwUXDjyTO7gRiSUi7umPcBg4ev
T6TAYrbDtzS2iO5h/y+WE61/Rsziw5h/hBMMojXnKTEhfPqqgqTA8gzPS+h7PduX
yxqzW78xjo1SWLVDF9CrfzF0wmWLFpRSx5NAV8wSowBghKBKm6mY+/w4KlxhJ3MW
EtTD2RBnWuxrb/QklA6AKwvl1fVtAn8GpZgb6EZsAa3I4SX+eskuEsHGcuLBrMgz
UkPHuoxmdbQzKcZYeSuN0obkcHrqVTgSdm8VwQ9ZPL11uhq/QV6u8USMEDZsu8g6
GzEhbl+L/xUp9YQRDBQeDK9J9KwHWoZl13oo4IfDFrpwHHU3V0YbgPSPfw2DDh22
7K+EQD3p3K9buskH4Sm4K+NCX7tYJrHZtxwqQOl0vrk1oHMU8VJ61X9ZZYj0PvuC
VsSg4X2oa06wIO/vB8t1J/JqlVMOYXwdKHczeyMdFb+v0lvAJ7/ySNF3wQGASHPy
nmrzOkQ07M9wRd8sYQMz356IRbMT2QpWew/Okhd7npVEdP6HXTwjbj4LFwH3LESa
3WvsN3AobPMBsJvzZv7Dl/X5qmbgucRJ9uYhVfMSojOuNzO38goXM3EE3XE5E7W6
Ip9/cZAemcMzvQuRojdoiP3RE2c2NL6GIcIhlqbaq5SyV2hK5KPfPtv8niWaA2VB
E24vbMlAdyk2neDHlqJs3t6XFrJI5CSv2vBp9R2WszOSIgg7KAnbzCJaoZMi5fAi
DF4ED4wwvnizs4hudQKv4FJqHQzwiEyY8y4Cvx4AD6kZdyv8PdzlhmwUh4s+g8NA
aFIhCxOJIVIFqERaT6t2gdEgq++IdNcD2PA61kb50vSnv+20FAy5ofRhcXk/OKOQ
2PI9jX+wEJD986VTyPJLDjYfPQpZEUlceLPxZEduMOUb6EphyDcovrPTODtRKyqY
PRJ1oNJb3vqmMghk8gsDdHDksdTXZE3xY+/2ziRic9PFjAZHB3W/fHQv9m87K2JQ
Y4TBud0KMFKeD0ABJB2KZk7omAy74ZMyXbYIuIqJx26jLAfro0b59YLjO7c5OV5/
rS9B37JPkDoJmjkBSOE5L+ljivJh6+zw+m6yEWidPqpxc1Qm1kzgVHFirwJGgW5I
s3iQAn7WPQQcc5Tl8v+e4HHgi93WmU+0obDfA80gVDKrc4UqB9sfR9H/OlpV48za
d7c9NoXgSGeptWG8nCpesk/QtKEw0RUOaS7fqwHNe/XMZcz4kzjZ4bADlFl2DKee
DEnr88EHFnX9OzVJKWN+HDNjSsKpjNTv5joEWOkyEXt/BIXmoN8bmOzRUAAQ5KgE
4bun1EcIJfBoiR7FTfoOoL8QrXGSd9oiS6J3T266LIzdGjuAbmvEqltzGzmVmPAB
zMwBKSl6sUmHkMWF7Jv45MHtg9TW4BJyRQanU1W6+Q9ELYM98Q/i9JRDN1aAOjza
3grKBkxoD0a6SPFzzDIclO36CezHmZ8oWKPI5vgBRXSHcYCNQIB8YGlrsHltoVbu
S2V8O9WAnCpAvwnafZ+JoFqW02VtRI/KprsOv0NRZXtuzYWsb9rAqGJm45Adp8a4
qhrUSZsc/8iJWBf+U40wr5ERPUpn88sXJGNKacp/Ic1Q5sdDbITjv/ssL+kCkqQk
klakRha9k7Wgf+Gj9vlqFhMAkXntAn012gkz0CAy7eAUr5L88yL6Ge97bCowMFqL
irRfr3ckAsl42Vkgf+q8x9S3cl3fppmIOLRcxTmRbAnpy73r9UA07QcvXXBrBB3/
0yb6JgkfPc8B2xwUGMl3TzB0W2WztSR3kEyiGaqIVXt0UxlH81IXUZPa19ShZvwV
3c9msLh9brCl2G9opBFsISwtwbGFyBGk69jeA5NeERi2j4WSY0mxo0a9PhtlFMHe
NOTNhzn7pwTgiqmexnijzN0ZtRd8bxu59jUFAsyx60ACJGZ6VmbdYGrSHnbTT8UP
7Vm32I6WUCWUJUBDjt9KQvO00ONHOIELRsEpIZbtumHvGmU2ITYvIFQEkeqCb7m+
G/9xHZu4zBAtwqlj1l++YnZyxPVj5bj4DtbDuPmCUgh7cqsoEHJYZSjv0F/cKC+q
Geunx7Fkcyz9Q4mmJKXrA0cw9rc78LHBxvyJHEkFECAW9w21WCk401XElEG5xseE
ze3gi55OMK4oigWNkgvfdUSgyS1QOcEFiV60ZXw5oeDB6YLV8XquUpkn6kV72Rkp
mlRHQ2n+cjLvpMKUChOPi4YBzwk93kZmIrbxVP3e4Yb83Yy14bmONBiNP0ONhdWN
I68qWrG08pAi/Rr9A+MiJxIHNcnQRBezKUXrR1/DUCA+uPfkADuAewZqKIjexFjv
G76Ia/8qf2GlDiuRYiCNfnP0OyIdJaZ/vghPwx6jZsJ3SO8QBt3CIQ0tfr2AGYxN
5DztLG6055GX71DaHCJxHk3Ec8PBflBH1EaflizkIG2FTSQxlcc2YqEvDRK7t++P
/RKcd+mr3jhbNakekZ5ir4HkBc+CJcErzAYnJ/j05l2BExWuAY1T83IVSzLMt2lK
gHMEzMcnTAkFbOrHiUroWUwXUp3ff8wp9xuABeibbGftZQDvjzvKzLe2fzLn4XV+
0YjPUaVaYYs0DBuHXcoAvKLwd/bLxEZEyUuhJJcUQMaimMMjGkxpaqve8ly6ICrC
OKD4EkBg6azLpBsKFggR2f5HqS53zBZpfZ4PYwARqm0JtpT8KMI0R4MKG4953PNU
2bW3j28D5/J41oST2GviSZhlWSSxAPERhDFyO+bYikLAs4vDUohjoseHQQhlWWDX
NERcetvtzANM3SNeHwf/gpL8MXNSQXcTP3wCqqOlUxmnswpWf0QkfOjCE42NxziO
i+qvDw5cVbnaYpYDyEeEyCh7pTb/wI6PZs9F0GDBcZBDkqJZ6z6BTprdb72gUqB7
qClfkzpW83ifz/YVVygmhh2I9ucVfvwWRTQsLFnFk7+hZ6EO4fLJOcYZ3fWBPM8Q
OGAuCeTVLjBLBwAHb8Q6VRkZcwD+1Z1VLSXELxWyGAPuxS4VAKXNEEkY6EFaAgKv
ZUMKdFQt4yQkYw+afQWhOj0X938COTTEf+bD9IWOr/EejCuZN57uUXWvkOCDTxr5
F0Nz7HZkx1sXD876wcLLGwwc6FNzGwX4wBf38SAiuhl+1lSC6/yNA6OKk1kBanWS
1PZq7t3jkOox35zjrRg0YCXWFFdPk3dnY5AylIvZsGAyqiZo1Xul45CRvdPVUS3A
tKP6USOsFUEuZhnIe95Bj18FxlaRbbVPtSRJo/LNRbGrqLxB8TFFwwAnhlR/gIYp
W5mh27uvglGI+7KJBYX85t4CB8gFwcfrkk9sOaklfWhOqrvO5neLmqf/SgH5PZeE
7w73J7y22ayV+qa6XbUFRezlXNWClECS93/tX1B0ADXgWHBdppses+koT3Cmtc/M
i2cqKkFMIymp72zlC7XfKK+5SqDZ7xAyymgq0xI6GcwXeycKH5ZoLw9R9kk2yAQi
AqwZhgvYZ+rxezePmKQjELOG19pZhfqpjxkrPnX/rZMpQ9koqjnR+ETqG3BfTa9/
ZbYm+QSkLKoa44zppOdtmQlIEW1n7MQMgdiajVsdB/MSYQVxJkZSzMt1wN5rpDW0
E+LVmoQXsz01RBFO3TXznolwfblQ8nUhHa150xrFdZCYJ+ih1o3MiansZUpabZtB
KH+6b2CFWECEDG3IQnMCsK0z/CgxSiGVWzYlrxELJlYtxJaAfEXWN+o7Nrxw3Dcg
J8aXb+Q7xinssJHcBP/y9yPMCXvxcAtDhURoHraZZFxqVA2dvA9RcRqIipIr7wVD
zhFi7xZ9LgxqlU1pBvlwMw5b8dDB3CRGUfLuSjetz3D4xga4Zd3D++94sGl0I3vm
+56xWsIIEhWDcrNwrHxP3lQwJTP6Sh7vyXrhcUxWNw+MHQEh9EGbMVtjOdIgjKl6
iY98XzJfUvbR66w7ijqP7ImEYW6DF+2gKC4d9amxnh8tvlk0rHBGNUD1v8ERWD/Z
wRh5z9IiTSYt6y0yE3LUloosJRB0qS7vWjNwpL2vqlzOmpCVV1FZhzyXSUVye1cM
+VY5zUzHmV38PKR+PsqvQT2CpmiSXx/I71FoO+doVmfKxR7QzjXATgU6MUY/oWYz
Inn4DQ9U9tjF7H+La9je0eCmhCV62InyXW8O5u3m69sxbxB/2kpkGi2vMMdRLZy7
KTAS1NS/mxudIH4mutITWPzQ0MFe/KZjEMbFhUKz3SM2SWHH4QSy99Oibvx1UYk7
XInfuSG3ame7OGbHwn/Mp+vj9ah+7iG5nB0rZhkeXe9R4IYQrgfP1hrqFys7dICC
Tigs4b0HSpAcRlJpI6Ez2vd6Tu9KRV8h+gTzVqBX+myoagGGgfQky3UClwsx9fRi
MdRFolLzx/42bUqKKNzu6YExe719o4Wxuze8uCoin4RVWimIqcdwl8tXcdNupevw
kkLgwBNm0s9epWuW1q2q/1loIvrfVsb8nzF1ES91IAMeikRGzfeggo8H7WmvTcYB
px/0sk09B6rIV31m/oGxlVl++l/rQuxpNXBiO+VFyW/Fry287fJV7Qnd4XGd00Gg
PZw/FC+cAIYNrQvxu8nwSHX7C5ryDXf0NQp5VGU88W343DKR5FyBAzCUO8nJx8Gi
peUwbIZdMivYJNueGU68lK9EdUD0d+/poVWhfK5KslJ09YjNxBtKLlu6Bf2j1KsH
zLp1xVkQQDn8ZjqbLx2YK8lsCq7Nqfcwls9wxDztNcqyBVPVs89kJlv9nMNVlHfB
EHct7955KmgWEXLWzQ6Klgai9Qjs8WIIkRv8ZW2qcOfpb+tX4xbd3UXUJAX5O9Lh
0st9GtR18mGprG1NHbYzZ9Ll1+pxXnaGC2KhZshkVswq0KjBXOXM1PNoxpWQwQbi
9hrCAe3OXQDbeVmQPvsS2gPg7dr+r2FaHK/CEMIo/qZhQyGxUdZ5OntBvIFVdHjV
FwydJwuJKjLPXyDtaYziWuYmtE/NKZ443uhFZI5E/1LYVMbrJQSk8/lw8ft4/lAo
A+ax0ywdNBf6gIc39dwAx++ov1RMycRHKm2iqnPGNAeyv84toB35QL0s7d2fvUdA
b3sz/9GaCKn/NkFfnTbxbLolMv2i7mVTeozFFEA5HtqOsgeMBL9zluCs57rrRjjH
AVAVeJuPpn5m+phUb/RaT38fkSTLrkkSwcziuW9fKMoB7trjWwq8k6J9HUh8ZE0L
l0F3AGnLt84Mjy13o95SsRbc4bl5sNY/9R1KuSBIOMzPu3m5sNVPvjaNuw4zXTvb
XnIeLx8FQZLjpMwNoOfK/lOaS5aG1ZRJtituWTQdsmdLFozDLfpIMk1dKBhSn6zc
ZbCRK3xqgFsHMVCLPMGDMscDb+NSwATdbX0oDaza11FTEm2SLLcuVt1M6Be5K84+
5sbJ8pL/LB+4tgfeB0Msan+4zzs9DXiVbTyPHUa6QueD/ZjDpW+YCM7mUE4GsIfs
FY5H74Gb+DL6xSGCR/VezDEJhl6A3Q6MG69rxorUCf1wIWsaEovTHfIkAXp94gT5
0EQdvjDTGf365QwJxqpQ4PwDDs9OHZWMzt5pctDeVIJ3KFW0lQhmsGW8yae33Ptu
gdfGH3/yZkrmULN4Lt4JLew0QZmDeSM9EUOFcxr7nB43Slm3Whu6WK+XE9k2B8AI
xdbWshmfQnmEBtweY6kbEZJnMs3e22+sWt1f1XDCSlzA1JdhW4tIRm+TT6RZOnaW
DCeXfbjOFVy0RxsH2sI8HAFqlYi09bY0PsLxutmRJwrHZ9YlGATT8aX4FFX7PKWS
gShinlmyDFFLnm/6pwvJYXV0/c7hMgyoALNUm209MlRSLlpvT2rbEU04fvZPfcWM
zF82KJ07BXerSqJo4pg7QX7pNnaA5vAE+IdY+V4426tcl6ukQ5Y1Oa2UXNcj/89g
CJJTHIrDTk90DmKBOBsU260pfE+KwFY5u76ai+Tj8hGuFOHxWIw7Nd4g9tqsTai+
xKnjJ8xpE9QEVurKLwPOM3DCXEYa0I8RXSqYr+4VsxVy6PRkLFVuFU/cD4Qqg63s
A0ETLcFY5eTHXh6hAgsCJr3ImS6z3t+6LOdrusvAZhMP3e09T2yLNe0deOidkqAu
wSKl05iDW+D71VbzMU6Tlkcfr6psa1aRh0A3Qobw83EOzrGMpuJvAIcLZf5Yrb1z
dGA42DCZCZZKSVNK9Ci6vNhu9dgzY5621LLpA06CWydrbmmBtpPtUm2LQ7Sc0+PJ
N7DVh/9pGx+1PukRlcIW8fXgc4AcniUxObgzMBkwPZIGHMAtTcUvipuZGVBjzBlK
QAwRDcy1rFxqUr7Yls4ZtgYmE8odqhRYf74M49175c2tyKe+8N+g9tj2oC7N58OQ
nLA3+H99uqKM0d3lbb035z9C7kkZAmCZ3NXrerZnA4OtVgw7erHgw8+scO+uTTzu
iz91qKtdtFA6nEfChM7ZZhZ2xJPavfBf6/6qZIXg4C/Fawpyy2oSKdHHMlxsc3Si
upwrLIwys3NEE6SF955p+50umAHTNptkSaHinepgt+8KWxqlHLm4uLJ1+ngB0iyz
Ci2wY4tQkezFtJpuL+3tmS91hBxvjoJwJZKmJl1xwyTDWJLXlFP58puShLTYgx0Q
aqFy16NThahZg8ACWXVBezuDEq1XSDM65Hb/9L52Gnb7aTN754kFSD6ZoUEjtHb6
teK8Ai/QRVTurKfOk9dRLg2Nm6onCZtluXd7QISD8+BXHblgZLIIlw65tQznd4rU
afCkpNdCq+y/E2HriRCsCQLhNsdpSvrdU1ZODIiGCO7ddmOwjQsuTTut8mJWlli8
krE0DyG4S6xNvkGhQJXtJMxkk4UMrkJg6JlYOhhTh13vts/6ACc4N0AVpbOBk1+4
i4vWDYfmQF+KMB81CJ7YawKfJ2xll5Zfucqkz5TVRgSf5LmGuxK/nr8CaOv1zL0G
8YO+eubueatPXKmmp2LwDqh3wHCT37Q9eHUBrl22sRyqN0jguWKohlASNTRD2FSr
Etr+sL/TJHNLgSD4SyXGrgmvtDsnY89oz9tZx84p01DTPQdqP1q6zoPNkPxjlpui
CCipwMOXKfEQxnBZtyJIIqfJIuN2Q9FZfefqGkxGl1P8KU2cynBmwY+u92f9ECR6
NpunjM7aXof2Iv7ICvDb5K5gJeEJGDD9rt06aKtE1W8Is2zzvNuu0xokOFcSUYq1
4cCaPUQxFxyHS2KP9e+fobsxkAh/nR0anTc25xqrbrFl3JakLmamMMPQ2HQUpoNH
ceclXSMdibGi5NNhIS0G7SJOm04UF6jWqACZSBjyCrNz34Iyo1zahlDibsRm3ppq
Xq7HC9XPEILINAUuFw72yWD17jtqPO5yQUJFdO3Gks4=
`protect END_PROTECTED
