`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFknogUGsoV9DN2K29J6hCvDYOTTk7L7JOM2DhTeyTTl
bZshhGHSKAZhHO4O9Ujau4H21t3ybTqnyjbbbDmgUb0MZ8xmqdkzd4CJlUC4Dav/
4kardSQYZfX1PgxcE0PIFPNFbOS2jKSyMydbDD70Dgv1IgosdUof+wO8/oh6a048
UDmxjTQ8dfAl4sGCXQz++y3v3F+j//pIQTGF3GyO3JW9klXhrhb+Ce2a2XE/nhBN
qdx4UXxpL+Sjre3DLxQDb4WDjie9pLmSHt2fXCeRK8psUzinxVha2TpTfkHaiclR
wKEjmQsHTZ94rAluTDuzBbesGz/k/1G6LUzpL8iAwJqZc/Ti6BnCfBYNfXeZ4MdQ
wSx/PZfDX0JQwGBCao/l0j5DXMNhbfgqyOrz3Xxxb3/ThstUA4+buRlqeJ36bpnj
/lXdsVFCXAhToS6dMKg+dhDJ+lXDs577t02WZ4gY/z13FcKvumNc+lZ7MbqG2WLY
kJLlJmrz5UgVGLU9riKFrLiuG4riXoQhmCCi/YKTPdm44qZUwRd07BrIIaIPAOti
`protect END_PROTECTED
