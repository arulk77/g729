`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wjucvHj7bv3VgO52X9q3cphpSiSPCQ0Zs9wklI+p95m
Hd9OEWmrpoj+4kBUqqH2NhtxKiBwUE4np3aSwhMrV0o9sjsBaqaEPKDarcBsWnKY
kNrwxD6RxD1p7hoyGiAW68iFiv+ZuAax/tiNpZW5D7gpog4dCRHdzmkiwiiqk3Jy
5/G1sE1tgfdYNtgXMBoSJfs8XUzV1yAFliNsZqzoltU4yxJ6TeoLpBKvNXX6LTtk
9HOpKx8gHh8fkGWZbPwEGVusmhJGgIwGgUs8jSdgU2M=
`protect END_PROTECTED
