`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
s2X6u2oN+fx2UEmqIhy52FIdhUzfU6j5W9dKf/Hq2VoHNYRlOZ+eluwuJDgV8wHl
74d2Mx9qy4fgsH9DSnSMsizpwiEgeR0Bgz+K9vkLGiy0NuIBvFr3LGvOh77zqclH
iMjY0e0pOVGtkouJfRBdJ1g4AGbUgzOvE590cjFLbob+W/LqUvvFqwV0FKAIkwtP
lP1FwHBVexNVt5w1hAvyFoUUoXLDV6OLrwvs6suEDCaY5+6idaL1taCnTmgsBmvE
vMOLrE0ry4NWDiV4/9T6CYHCMunSQLDQrgTPlptPUnURH4a1c0uQDgy2mKvaGoWc
t7qggxy5KwdFuFac/Oj2zufrguEJi4alCpb8dTVu0qmAIl0p1Mib8n1g4eAq/M9O
L9K03Qm6N+Z6OyA+8I45gkC6+BM3sZnP+Fi7CH/t6dg1ng4CezSLa9g8bA3yf9H+
Ea7HxR+7lDdQpoM09gb/WMa3zGOSDtcg1RmUfP14Uk0sboWj4jYvFIjuAN3sKRaz
YRdQGCe5cxFALyv9oRRhyXjTgH7Am12ewW15C/5iVBJzkofD8kiqLyqQo4XC77dh
S/+S2TaFiipgqqI3rR43x5x8vBxzlO6bal2cgZvXxamSW/H3Rg4313JjAJsNu1rU
pgFdahrAWpzOBr5OFCBzMMZdQ01m+M0SNy/4ScsX+wnUzuwIfOKbrcR1A80YjKwZ
hokNbxFT3yvLdiicL60BgFF9EZ6vry6Bo+ohZ/Fi4xDAtXqEh553P92xx2R0mDAa
afarCeOTCwcEgBq72Ak+0r3I9CP7v9mmNomGjtbIyCq0Rv0FeFhampTNAm9c71Hw
Lf2lvbudd+zhXTN0zcGHs4uFkB+sm99izH9KyJwbqt1/3zIcKUXPyUHB6oBVljyB
ZHlwR/DPjPhJLU4cePsC8SNriU52rQyqbVszpUP6si9tmH+EQ8dCTmT/k5g5uyx3
7eB8oHRWnv87CRb7nPnmGYsJSxIswre6KaJuU0XaFXaCF4ATnt0gyA/5PDcSA4dq
l4zeIOY/Za+Tw5uaMq81yeUg5PGKFPrucp/OFysrn2A3fAui0u3+R8VnEvvvjZt/
Peu5H6Z9dxGKg9rUU4uo2mKW6xkjBR0S/LCN8evNlGdGFeB2SvCFE2xElcfVSlcg
y9Y8YzMRnTu9v0AZNnjqHvzzn/qUzAQxF1HbCTv5lUn3FlNSUnGHrEK0qxK+ixbV
PYtERTVKTvFNvyxONUxvh/4YWfNaVOY/pRNmAG9EPLC/uJMeM+NuZVz+L0rSb/rV
0p4EbjB7+SXPBHGRYOIpbWXCR5dQnNo8Hso2sDCGJTjSf4SDJMPv1F8txULL0Ynb
6saJO9YgSoF6CRzTqMkgKDaKZsNqyV36ZaO5p6SfbE/14Ixr9ZD1BgfbJ157HB+S
OBfK/wI1hpffqBJuc9uDDR227m0MkT9aTuf6ImfCMG6fqeEIA9bLe/mXBWYprpb8
64eeYdDw5XFFIbEz3YRTRiNnxHnYq2HLpXjM9MTZFdbN3OShS+8DqOwk+NrV3mGo
bcKP3AAS7ovFceGuZfdWZ3twF8i0rI3vrxngNGV5ma5oLTmmHqpjvRTOnx9y6sBj
D1mc9AZLoCzHuS2gKzFJvYWRqFcqbHECpDr0CnWfRbFbfzFJiQ9X+d3S8xwKtiud
azXRoG4p2CJkwLUTZaairl50GbILYmj00rQXnuWDmvEXoKoG2+pkMziVeYj+x0LW
IIQcbTHZ2WxukJsdmUQwtXb3Sw6W5SOILDpFQqIEPUdoWuyAVqV2d2gJJC8KykLZ
9uRrDtCdRzCVATPKG/4KuFg2qLU61Jae89n5dMgyuyODvVG31VXHmVSVPQ8W3IYr
FS4PP4+bL4IO55iodU2+xLyvtlQ5ZWuHN8AwxN0dt6vkc2/9yK5w81thExJ9jIqZ
klCZmC+wM2CWOhfp94uiyRYYnQt6Qhx2liWUN9B+47FGsoVdUOjq7SlHCUhZUrSA
+U9xsrPYj8mIZna84GMww8jz2tyPSiA5nPtUdWourWrV4QQEq8+1XS80mQD1NZJY
m80ZoQKVEXS8gZ4q2FkEmr2KsM5YHqMQovb/sp/Lz7CwWuhmJMIhBKeWQWB1+ihe
huUACMHtv+vqtkHu8B9SJ9X5UHRvXi7HUry8tC6O9ulkHLlb8R8wVoFo0Mpsrntl
X6f6BpoCwFy9FCq5Nuc4H8MWU+Fd/xBdcBlwTe1GIBYSggTWK5IdQlwj39Z/HITa
ttHYv9EjNciMPtGBTuX2CMbSi3AQsKIddRe2qTuUvp9H0lGW5izY/mm/dc25kU+o
ZBEmGZNp59ho/fQpi3NSSe9CGVN2vuqktIGMKgTm+bmF1+3GJ8AAf+8RV3QjRrAX
NhlJZyE2D6X60M6zAIHLlVU1iBJQAJUgAzgUu8WsAWcB4V+LhT058AhvgJXYXu0b
xKgDZuPCvV6lp/mehFK12lPxVtpVxSCyLRd1JQthQZoATEZdP934TaJPXj3s59KG
nV8HFNK/OASrBoCQ2no3sufgI1KSFU2SmWyBbGwJchHL0ErlMnDrtfbdCrUzRsg8
Y5v8qVFuDbWlxlGnm4z/DbwvRH6TiSgqR2/auy/4wMSLx7HhkuTapSicXXkpTu9j
Qi9fCQWVjRm0BuD0Acn+ojmxk3fS0DXV2IrV1pSzUqbhqaZJS6FA9Tf5SkSTcqDd
HSXVMZ1GshwE6KFZ5rTAFHQ7e3wcfEP/TqVsf00cwQ4MPnQxsvMECdnhPK+KEWJ2
xnTo8NiIkdtMH9NQYjb2/5edy7EDo1j5N9MoIiqwzWx+/65LgWah8fZnG9uqQQAe
WhW+SL6Plt2iIqPOpUxEnl4elNenRSGmuiUmVnPki4B9ehKqAJZIt/r4LGpS9TDf
q1ZNQkiq8bIJmS2FNY7uJve3P7epqmm0UpVI6AKWcdsTqnaxUg4Gkt3wMkCHgKLw
w62Stprfa3nEF9AGeOGbJy+pHz2VSAULE4c9no4RZ7JV+YRvVKY4BkBwf0wkoG2/
oq5Q2yBHlfBqXNhmv/nSUtH8JhcHet9DVoUFPOudDvCDs62JFA6vitYKGiRUd1jl
nLGT+ip9DauvWYnABeRxvI0uZH+GCLpA0V6Ng2MSpfD9OqC4LUQxMlrqy2hVgbyT
wIMgbcA9WH8ctXHnqEowc8zGZ42jYAW3eof2ZOTFtXf3sxfA9YAdFNdiiymjNXcd
Pclk/VPbT0dXHWvOeWs5aYCX7kCNTs/51DZgEVPt5glHHEPVW0I270w4QYC5JZn3
+gZ9ERbOeoQD3v/6f5MZ3pydcthT/UgoM2QkummT+B6Jn/wKYAF7IKnWPNqPLntI
Wowkd0933XKnnShitLfe0gtKACA8Rz9d6MlZUw4UclS5xjESI1c7weX/RgjVf2vt
6RNuoKQ/qqEfweiZIf6l0AEW0DLJGlJpMTiz+XTXCENdbqD9zf5ebwaT1QYAeF4V
WaeA4p5fhwyxFsWthHEfp4iYI2KmrwzLevXHmcLwfHPYrWr5z0Bv0HXvPZOWjHqg
ZzHGF38gtTj9khW2jezvtj6W956AqM7W/DRqXDYdiRT8Ccd8J8TJ5Sv4ekJQoLPN
P2spkwlmIm5YO9f6G3TxM57ILohDNe3rOFh/18ndcII9GKXMNJgMUP6ZxpBVuRSE
1qgmQXlITSSHeKtmKDFgQlNxfwlSWV8ffqBSQvy+MSiI6+hjufzlQChDSMfEJa/5
DvKn95Javy6hh0MbjT9/oRXOADBF8DANsanld5S8Rl2RyLdOoSKHNAdpKD+Q9dsa
TFCm4MHyjGXcFc0YKtebgn/SPpcl4mXYvmUM6RrhURI6ZtAd3Bir43bzXJs5f9DP
IFV/Yk8RA0C4UEkoX774syEAmMnzuYVYaBN5mMQNNEf1ahr31SScNG4e0LzpbTq9
ceDKmAazumdxWICYm4nhUhYZeC0dPUk4ReHRoHisnxLOP7jCWO0g8w/sqvfu0bOM
+qBzFUA1ZVqsefpZ9M9Jb/AvV28aTvitPcwx61M4TyRhdMFS3LekJ/MVuDmyvl1W
P6+3rF7+6hnM4amnllPJxMjlP8ph06quVeicf92TGPwsr8RfIAPKZ04I7WuLe4T4
ngHte9neR4TCDYtotN5iAf1fdk7NehU08U+9AaR2k6GzXfiHL8hpRqgzIYx2Kccc
RBIFjLivGMW2Ke7Iro/vf/Lw6R9TpxtFItEl1Fz0AzkyCL1wksk4CjKtj5tF1O5u
PlrYgRLYA2I9XyS1DxjwrIhq0B3hvWRbDztecGaLg0selLXmWpCC9kP66a0062R3
f33yJ2bltT+OmEHyPZ5BWmDdglRd6hOIDDsYMbN3dtboDh2yOY4VOEN1CMTX05l0
W6ntx5s2fZFKfHkFPEIbKqu5J+W/n++WbKCaBCie4GSdCIGtCQ5MzrpSGpGJVVYM
ykTOFTHjO/nG06eKZG1MnwYTvLcPhtx7L7onLk+JFvs8wsZHL4AX630U5eqZo4uK
Pl86h/DrSjnU5xd719ByJNCkvmnyMxlvONhgIojBzxM70P28I04fMwOLzb/j+w7Y
Roh5IPzyzDzReRt6BnKtleAdpmYz1W6d2+gdG5qvh9l/HadIj614/Gj0RtZDmETg
uQXPn8tA1g4LJHOprqGn3Z9/o43CtRunq05d0n/uFbmerWvJcLuVUWAIWHlc+7o6
tbWkU6jAB7YyvbINFctenR4T76AQ/esMW1ihxNisguWZplivgRxNh868xCJ0Efch
kcuRz9ytstFSnLkFCkgZLIhwRozAVVO7oNQWYSL1lq++cNAxRHs1/QREn0D6EFHb
RWrpFfksnlSoS1EQbtorEvmYHKNzluHF8/2GGQ227XwbaIerHz8Msfu/1aTJO3k9
QyHDBLy2tpRtIr07L8942MVYVAWXc2N0yqF4V9ZeaNOArv2F1TvpcjneiuQcuzeR
MIT4ZTZrt/ZuKzv8YEdqrZAdNv5Ss9Z9XSrmC6OI+HFVtsh34IYzL7BrDsUv9qHw
lhqMMWqHawDtQBjYE0GCexcDdspomceJEjMCYB8Gdm/y0JgaXgoJs+CPr2zH2wz/
TqQaOYdWRFjgvN68gbo+va+YWFJ2ujK5GpWTQS4Btysplo24PVnn+afLYTsh7u4q
vYFzf1rEY/oIXLBx8mPS8/u4zZXkR7oopQXsrnMkCSpHwBW6H5J+CWND/IH4XDe6
anl+Hi9npdzuPu9vI10a0AzmK2vWnHo4YSAKqEVrSAkFxv287kTuljcpyw8t0Ih7
00kIADlLSS4ncGgj1Sgmo1uZYDex+xA2/REj+NC8iABWhBDNXsyqEz8/puMB62Rk
VtfpFU1WYVMJgWBpjgmwTCW872X2m2XHTVuHv+rkQ6ssb7/q+NdBsKVkDfbr2IiM
gmYXU4+I0uaoBClynGer+lQT47Rr4vK1JFiv/P6ikfWs7/BPy2X2IuN0/F21A5e5
ehEzPacOnizPqHIFnbPpI8n/hmxlGuSj2cPnckHxjPdl16DTLaEY9TKi6xTnd0S7
nnCFGwwySBLVlGG0Lo0DnMAt2kEh91uSuk5iSi+fqSGS3gop61boPPBvkrrUgMUm
j0fsdrw2Dzo70HK23wt4c1cLBP3TrlgOPnC9SD1kY3y8vdP3Ldhda4TgsxHoqRXW
scjVP0tdIIcyfMYL+X7+iAmy7XGDn8Nlq6TBYx36dYFgZW+urnv05/esjERzgcVp
soSP/c6foNpXkO3laWW72thXtGDY+3giCxTb1wYUPcCglFOs7cz/1s1c3+i1pvJf
2inFh1QeFvl3w2LfvWnepr1RNSy0yyrObr8D3EIdZuC4LksDNUtTxyFQS8YnGMqy
AvZdfop3X7un/Y+zYEENM1LjEe8/APEhsS9kqbrnsStN75TY+4lpj+2zsBo74G2Q
fEL16uDVYQmxvspaXEhgdDICkK2Lu/Jit7+WE6hiYA/fjvlE88icJvwq2/dKYVw7
fYNG4EaP/JbO2DZTFhVPaiSOongxxbDcnWhp+/3Ni7YEsY/S/hCWGaxsJ7sSFT5j
QHahEhCoZdaJOjdNA6WR7qMxRv2aIyeJChI9xkSqO7usvSndKAjlXP66ksD5w4mM
OtZiplDzDHPwZGVI9bdBGZoRdRd380wfep1IkILnrIBQj2v8t7s8kMnO6Tt3rITE
9AmZf2Di5/vRSVKUcqSQaJgEWAQEnORDrn0T/1pk5GS/e/2dVeSXBlaz7CD+qShe
QI5602GQno1Qdmm+fHh/ZU/Cr3qAE7XxDOv/CcwKO4bxn1SFjE3QErnxxMxJN/MU
2uExvv4+HeZ+qEqRS/ATTjlUFmrDkW+sikYwABLFfrmYKFlW4QmFxGqzhaedI0KQ
nlCrj/cDsG+F3KopzT04JKjhZ0cN41NAi2zYlG4WxeDnVoWXbGT//BrwFB9QE/70
mH151rsCOYIVxrCo1IMPkrhXWjeyZNJ7YrFGZa/Whl4rUR4AvdYcYb3dQWIqnw9t
oqi7Lk6pib2WL+U7QzYAYT2Cx6y7G+H24pePnmKpa+dMD07dxfST4nqNsl6j44KZ
7YSSLXDNNrMVY2ehLezl7/yDNWnDtE275UKeTGVP/w+0XPG4PEQL5kfv+Amb/tDF
jrNfN14jNdmdTM7xbGJZtKkFOY3mquqshkJ1W9gdZlUbiZeOyXau5cJOp9JAWgE4
AK4xPNuW3bQ4IRXfMQG7XTkOuTGTM3+svQ1Puzgi+8spYuKUGFClikhh/KoxWEXQ
qzEbVgXoPMsVrOez0LIGe34XMMeMs05QyFoIJReb31yRpcRuRp5vRm/3ctQ7rDwn
Z6/AquZ3BMETpBzDLBoZ3aLr3YdBlrnRN0f6kUCT/GQ=
`protect END_PROTECTED
