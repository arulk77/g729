`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41j+wAVwubKgoT6Xkya/iE1ACiM2N+HcB3HQPgF89w7G
8cqR8prKHRugdm9+gBOvsfrtsOJL/Qfs2vWr8YEyax6fs/WmVFzeoz0iZkWYzR1O
CpjD8dFoIhFmfS64LoL6g3XzgPiDPZ1+JH3dxhtiBxPIGB1qyrDCFJ8NK9qTQgoK
NZEki4z8JuxMfao/7sFudDC2xVc/NJOCThcrewSI2LgmCXX5gTJaWrY5CSSi3FIi
2LBSx9DNsrtV+TYu9uixKQ==
`protect END_PROTECTED
