`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDLgt2dSJ+URfA6aMStWQfJananfLQNLvAUNN5pK9iMD
9TcE8G8y1GN3bFEO6XqcFyWCl6HR0sB6j6SEc+m20X4GRWYR5c+B8EvQDTS8N9zC
1hzlywZZMYGxEw11XLqoEF6g9bOccyvXmbHd8fMwr3aBmbtbkutYlYTHYN0BK8Fn
w5rGsIyH7YIcIF53vaVLrA==
`protect END_PROTECTED
