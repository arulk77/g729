`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
GK1XhQIlGdIv+SkT7w7z0smo3FkdhiPvTWEpFCspKFQHfFbT7csf1rIJkRvTyP0g
Ap7hSconX6Xot7OBY91cY/y97QKtohtSFyAxb9IC61fenWiZDLIxEawbf/6iQNrr
XDsV7/q/JkyZwnvrTWJfFYy/SEYL3Hb/3MV5x90uvMIJI9X8H5ANVU8HPiQ1B1Tv
pMw+25nUBGPt5Fo8FLC9OcCbNpVjiW8vYO+sJoCAnRDiPfrGbyipFZNdPHAbcgiu
1CTZWG23XOuPE4EZgSfOwODRFkDAt15PGGGU9TX/GLxGGz4dG8NfkpFwPbbs/T4e
v4qbHJ4Pfuz4Fx4psvv8vZywUR0f65sxZmuuRcp38wA5Rj0iHTNnDJRCzQI/muow
TWQfFqUhQylFbTwLXoTZipMmWh8sbJQEUPC/OXgSa+1M056EHH1og/Ejdld2weAU
LZtz/I6HMwn05TrSGKliPSGPqenejF8/soo8KscvTaCzQEE0xjlcui7ox0hg0+6G
QhYIBhSEBm4z9pI3kyFAlr/ZJSkxvmPU4efXZl4/7HgUrNzYWp0rUlEtm76vuAwV
D4lxCdkWgRXWZYF0Es53JPUSivHgjXLXAd3SjzXO/F/wtXaqj1rK6wXlfyNr7ZH0
OsFW/2h6Cmgm57Drns9hmGk8WUInbRkIB10G9mv45lM5eHQgNL9vTz7tA0havCfs
nTAoNljaHsnaKAa38Dq3LoIvQiGgLzT9WI/CcwtbQdY=
`protect END_PROTECTED
