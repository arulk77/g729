`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDJSpBhc0ixLKw6d/SSyKDrHStgSkEkEHcRHwgH3hwXn
mnH+Go5gSfN5wS1s3jU6reAYJfazACzwluW7c0H7iQdeU8pj9JOc6klTh621jNwz
oFMr8xXH9etdzXHY1kzQD2TnZknYX+/UN7xnei3h38YDTAFcT0jA33vQh75iigmR
7gT2noaMHNZST1Bl/E2Uj04HK+4Wjtj8M+SbNI26pLOI4ne7k/jnmfspBjsCX4W8
H9PRKhyX3COqC5UTYUOp/KacCsZaHnUTAaqeUU03sOR5kZZ7YIYpztvokdwHE9io
yPXNJCq96mWIbBwRGqzBxeVBWoi+Of8/afPwDQsPUPY=
`protect END_PROTECTED
