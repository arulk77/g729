`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49AhvNfZxNLkM4YpJMwF2+lexq7eBdLavA0ylzPfgu4m
J+DaOMg20gE5tAJMr/PxYJUfJGTA4cD/2+rf0C02CsMN4FGVZF0bDTqvArKRYRS3
igkku9pjLLrJ9lnIE5Eiy9o4uIPcaJKPxjAWAW3EJ0iT5C8q7zhevDRFJlMPjUIa
i0lXyzpg2oFohUz7Y4PMi+/FLN0ZqpAI/c5C4f94puM=
`protect END_PROTECTED
