`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43KCP2/+Pp7uow01BW7McQT8NINbzlu6ZNmJw+clwYU+
MWGO4NPLyOIACXxROjrDLN+uapZTZBTesvAiszQcH/P1dUvyjObcS3xBXXhL8wTM
EeueIREbxscaW1m1PWpP7S+6m0+7ofMPQyHA3EA3LTxjsmsOh/8FXgwezUyyphYT
PtOMWqmuiNVf00ltLu0+Ze+miRjfNpOPqEwqxmjJwbDI87SwyUkOObXYVXxpt44g
v2CtSSFVydol5715YA4FenFsTOAYfmJtlRRTtFVt+JRDa1whhIEQFfYb/NeF3JpR
m7QYzS/HunhaeUFHm8WWJeCECHh4XSfMKlNeb17NTOjdiRdKrHsG8wvtG0lkdFqm
VVikUsYJ2Z6Pq22zdE2eABuvr+q3MVjXE4tz/6ICONYsKfqdLGplMLd/5cIGjEcT
kzWHlvrIJUnrydop1y3dJs1DpQWYIwjJ4yPg60a9eI/b2RqKUQPARN3+I5dVxgIl
`protect END_PROTECTED
