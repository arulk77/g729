`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
36A/U5tO69wVl401zVMLLQBhcz2SzGpU6/t3XcLIbF+6u0xOGOR8IYUj4pVWI80b
vcbyeXpoXFWfd235aHJwZklqbzNqhXomQUjI5Er7BQ7tgHmdjAbEjL9RYFb3mB8r
csnBorh+fDL4qaBsp8FyI3V8xyzB8lj7IV77XvCj10TRW7PFXoqKy4ZtTcoqfAV6
5GV1NjJPj01Zd0QhC8TJE3g18MQ0FZwOj0AZWTOAkePhlFPhCnXyuUmHhlHg3lbT
ff3yBLXkjKm8V6ddOvgDBsrHFuT2RqqUrEIID1zNZJ/XiN5yu/SkMjpJqXY5cmF5
H1ht8DTiLr4zDZoc03zFZ07rLnQJmZiEdfLPVVPcF4APxDLD0os8L08Zx3zkNir6
`protect END_PROTECTED
