`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Prgb+lMGK4ankHVaNnLDq6EBWDO/XGL3O09ynEl0G9sn5DFzuZHnBnL7+921OOHm
S+KZKXlnwlAgoW8u2An/m7zhgMbG4nslgzAUvJHDFC0he1A3emBQZsB1aV5TaTQ4
KLpEJUQ/sriDAPRSpQ4gADEUZRT49JCoFGm1Escw7Ji3lG5HLNsMegQv6VRaVsbY
AxWi3s1MM/mlL/j0dV474KEgG5nSy5rL+uu/VHLQgmG/aRu82/gQMUBGm5AWjbbG
wgNq84lx4InqrQUNEayu1AOw0u5OVTEeM3LHwobjl9mx+h8aLVLGyceCpFXInecr
`protect END_PROTECTED
