`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4y1+OL+MXZw0TYfJLoNNnkHefmTLV++M1EvKXG1L7cn6
DkrlBOI34tYicmnvcAmNUMQy0JvrIafUeTVjiFJZBGpVCeC76aZKrVIboh5uhuu2
aCqbYDhTys/YTSC1j8qkDTBQFGfRYQwWxxSZHGIucIxGZMnqHdCpSdELXEGSZdG+
FqRKuzT+CWOPH2JjJV7aKBh2d6i50SzGbB0Y7f6RCk4=
`protect END_PROTECTED
