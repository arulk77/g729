`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMay0CBEMrGLu9PsDB7EViwalRBOOMzvmxoWXqjLUWdB
6sIfOjSK8rDumk1He1TRatNu4WIpoJWO8KLBpO3iLxXukBV/LVDPpnnap/Nd511J
LJGlz43J7opAX4GbA0W7IQ0SETqNi5lhjHp0/fv1AzAhUG2MhrJitDoUsU6u8G2i
uD4VVb2tQs4MHQD1ueaYd5x5rjGKy680yTsoACWyWP2uoRRhZ5TEY98kuJ5vVnoq
4wIrbXL8+OLvnabfQDTdNu85YN8+p90A9gIHz/IiZuyZDHux2TGz4OELevNbdad+
1B6o1FSa6MCwPlMwZUoEpw==
`protect END_PROTECTED
