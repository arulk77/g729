`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKuMGpoXPle8ZA3MkuKdhXvuckDJWvEp0Jtb4JaRdQhZ
5Ap8o+qALbk0r2Cy+h+XkADa2xJ8ZTyV+G/Wt225IAIlFFCfFmhvknrCZOaDXli2
cB9WF+l4XXq2Mqjy9i/mSV0O8UpZPjrQukd+G9SQ+UqgXKN+l08aWAnc+kqgQ/Fi
`protect END_PROTECTED
