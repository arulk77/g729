`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
AyurXypHicL5GZzjSr/clrG/GKcdair5U+0ewpJd3JRZQNKa+64lPuP9Tp9txLre
k2ubfxwj3c1T65mP04gBfZBqI/kme/+0LPyfvs8ewI6wbSdHfMsAzm+EN7PHPRTi
pEt4aYiiYrASeptNh04nPZ4GLG376C0odaEReAqqbtagbP3VecTCxzvShYq18l1t
+a98dDXFo3TPb9evwl+97TlZaZ0XVKtQbpQaYSF6O4Eg3M7xaNH8kIVe1J+nHiy0
`protect END_PROTECTED
