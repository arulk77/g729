`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN03q1QQS/Ys451yhZxr2DpxYmVkXq4wM77YdKJKe0s9A
JfI8/Eeeo9ynYzwy/LJMqGJCYlrW6KcLVFOYK2wWxiScMjBdBtIYFFbgTaRGQ6m1
dreLTqvy4naBa1Qs6TbvGu7Ib3NFmBPEmUxX8+15xJgXwfZD3R6sObkb4JOpRVVm
cevhYe83Wdec7fkE3KGHjQt6vhyvlWBoyMQ7K5xinKpoT1VTBpfAbgvGcWZMt9OQ
5wIylNSrasZBCk5uGQ3KdQNztvsMve84e8re43AuB7xvcQAg3yqoopSGi4nlhqp6
BPLVxahfL2kfUcWSP0rHvDFhJOsDq4gly8xy0yr+4oXn5IeSyXm/2BzJLdSdCnJ3
/fCWf0EYiZlx9ocf1oZIz7C9YhL8hVZSJG6rAn/mOoNAFQQ9VaewaYtXRXYnmaZc
RNpPeJNJKHlvPG/pwNu8/1faMxe986v9guZdzFu2hDv8Tc137+pN8t6cF3hBDqwd
edtM8hefGNBC1YF6lLOPcFZ4+W40KHYHlHFlxzj/DnaFJpyKqpmzJk3zqX6DVmQj
apkLNdJZDYruKfWO0YLHxoserhC6cOlfd8ZYvlemmFOCelKfDpA3GKddCes9Vxe7
7fElS16LkayH0QzcgfDOTeG6Ei8cCwqn4HnP1TDYB/Yavx+XkhpAle9t5Rk3wRha
pzmvpYXsz9Hgjgul4Y+poLt5h44rI9foCsC8JIXOZjZ/airTok6cJ11X60Qx02vh
Xft2iNnu2uJE+kGzq4zJOirPMlsFGa51bc/CTaGScw0fsasQdhi6H3AIZ9SHVopj
6cznquywFEir1P7FbJwBr3fBb3npRRWsW3kbqCNUJ9Hws9Ey44tGqu7UmThm7hpv
jSJ7N5lOp0MPVxi5IIYo4eo83uY7SCEbCJ3/IYy9bbSoh1Fba4Mt9zft0UIJLxbh
1HjC1HTgvpl2VCI8hcmqNycN9mdoRgXRlCqU3KVd4no0lebzmVUgOM+RjpovOr6b
M8IgLn2LMa+0FSBb1Pfi9wz2GOFO1qcf82DvW51qsbpFz79PuLVt/2kajM1fXfqR
6U0YgEmaadKCODlDYub2iPlT2Hta8n4AXP9UlMm8U/d5OXYNrbe7S9MDrdJ3GxM+
22iiwLYuoc3EyV4hjvTDyEmnD/p89D3m+BodVwXXZfA1tfIG9nq2tdBDrgACS4mJ
y+Zuub7G02GyQ6kwWgzSTXJZnMf+lyUggA1d08hXcszyPL8ZRci0orn2HtO4Nrl0
6GdLbBDCfM6nqWx72uichsEfW7vaKzCB6ySLkRP+Unzr4/i98szT5INAEVK+3cmG
YwYNDyRiNgGi/Y7ngbjxN2SToWf/GXYKNCkb4eSQ4vT5LvSJ+HxC8M4xluglbDFN
0Y5urr4ssFxjs/YaTHorgofLezEX2iXbdR5Uw0WYyMV9kaGgbDQ9kSkpjSVAN57V
7D5eAyRXOJxMuM2sgGMW2raH0X3tRVAXScGQq/TfOATNDswUUqG0s6cxc24/wj77
G67GjazFztHuV+Gl5rQCknMT8dq68uyuG2C2jrhBFML3l/pFGOh8qlcvYaQ9Sqc1
n2ERUisLwSHKLsCapGyIr45OfA/pGQ1zNkp+vUYMnv1Cykpbzu58lp792b7UXJ7H
whrVIEATymIxPJEVQdq+Qu3sJUXV7JZzqxqiyXlsl8G3auh3GmUvg1CXcgTx7VI3
20UXvTmpq79s2rio3cr/24fxtzyfQX1sPCqGCqWxppC7ItK7oSOMsQ519yK2nAoz
/AIJoIGDA7L+aE3jxJQutEfnXHXW9eCrcPJMkJjfvn24v6JeUXGroDsdO37+jzNG
IYeeHrA7BvBvgaD6s248UhymcSm1Xykqa4LAgwVuTGHrKkB5ydw0FStpsYDJGjz6
mupbJydeR32AJRTQuM6wbkEYqoT56cru4T8CzPjhQh3TMd7ajlJ6bQmWpBK8uwqj
XzSz76rZJ02E8ltaNS5c/pn5SmXwgamnhYYacAutpkYsw7+/LdWu6xrPXpuseudo
3EbqpiIK6C3CRrR6GVE6og==
`protect END_PROTECTED
