`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aUw7Knev1oZyFnazsHVE8NYVPgZkJGTJYvcSc2OccjVB
ViITGg4LJg4bCqj6xVMOsiEduAEMvAoV6StHUxYnv0pJwJhcRVQXmUFGqANZdAyx
Cz0TvxUPfrlF2VToxG9fLJqSptMbaBQy53W0arjpT+yJh/xgmFyR2x7r+yuwPF8Q
XXX7zKGTpJhdAuG4j7kr1HjLCeg/epnirr7JlvoYCgXalHfxjypX7tp5b7myrOT/
pk1m728whufNCfqSgh9WfG3V2TpVVn7+Ni1F0LmWnIWHCw07ThYj7H0VFohgevUj
AUicT4qSUWyLLXBQJCp5I7kdNgKKu/y/9H5fpYFhxiHLdMnl/H18NIcMrxr2ujAx
HWaxkX2XQfr42By+qoTvA4J6ap0q19BYug9zgPWajXt8X3584ZlyS7txi74Xzy2r
+uxUBVPk84YEicdYtxlLnAOfiivEfmERyR9Y4NIER+65OCgucFRUHL8AkGXf4+mc
wWBF5vLiclXbOPhJXRj006XKeJGLLWfU9qVrVioE3xleo7sC08rAUJTNc2xkKvlQ
qcQotmFLTDscY7dQaK/6hKZlO+kS0kXxG257eCucofHjYGEsdnWgCeLVdvgDUQH8
ik9j5DFCQiUED17fsN01n6ksp61/QwLE7VKtpS4sKLCS0708oGRmbCmeuIM4bbcP
f8qFhWaZRiINymq9LJR7KM3hEGawxmjSAbFFruTXyEsXGiziEfwnp+Q4iY297e0F
YJ9YgGNGSqwv2Lx7dbnOh0oqL7gx0et81gnVp9dV/C+u8qoScC7iaOU5YrLCYOTq
811iF9HoHPwgPU3GqsXfvwwacRn5rPTUSXqU1QZQh7pkK7FhpMO7zU5UjmUk2PcL
cv6kqnHN21nD2Shgi2bVMmKFqLIkThP7UqsSt4ICx3wJU9lpizBRCQY6ZtWQSBoL
jtoGgmp/LBJzpCFU7YKw27AVKUfuIYJq1pbd3KjjwWnbkyBWIW2pCP1975Ap1EBI
/IH4vVExlI1OlaLihgMQKT/PtqWinn4Q891gT01tnB8gCmlDOvQ5E/G7Yh+4H07j
HlyM4NOFnMym25/DyhXIZq+tE1e+wipl6rxYJyIxiQ4dg3m8+Dhu2h596MYiX/4b
/VvlVYUJ/enFsmoum70JBupIn3nl/xTwAKHfY+WynBC46XPH2h4YfQwHPRlQyKeD
8Xee3903AwwdKEYKbTlZAP1we1MzxBgVkssP3vlcZ4dCPcjt72DmW+6fcxr2gtv4
WE7lYKaNKCCbCOxIxWzykJifN6wFvUOGUHIwLjLwOilRUsj3e6rYkOlk8Fu/UeLX
o5w3uAvgKX1bsdrezIcjzctd8Z+EDyjlv6m1gsfiojn4nc17elyw7rBIv1GLY44w
hPCpXF/fvGClU4u4pqKl16NA72mawHHUega5RXlFaWmpZ3lURG+IE3ivS5bT7UZi
du6i74jAC0YFsWR2yJkCpKgB6KfbquZUXlexSvGp4DJ55Lgw+YYfo0ButD9RxmXb
aYbcnh2migt+nPabcdC9EXrZFMovzPj8pRhM/lQu6KXlHAgRYUNl91k2pOus8Ec8
0lRNtAsi1xBvh0gorSiSgCanBc/aHC0x9cKmxoAcr6hyerCswr/N88lOvIEmFNBZ
I0AaymaB4hPt5mh9xgTLV259a2k1ESZgH7OWUEvtbQrG7uTKH9jO6axvOldXLIOp
ILZWtzjPYa1fykM+poCFcIS9TmWOQpYG5KyzZTKiaPQkvtnmGHfkgaafJcSEBLYg
84Xdw7/2R8O3Qb0fptXlhKTieERIF9zxOOSDhucbQ4LWsHR+OQQKgoEZxUfSf4hU
N9tSy0mrLAYy2/xmiEIFJQr32AH8pVodo1SGxfz2Xc1gsQOxtrpnsxAL95HW+Tfp
gSSouuZrNmLPwnkK0QPjgiUwW0fRg9QNwn0YJBRan6kko7K2E1d1u6zycIrhSpyG
ZSh9rtvscvkrx0+b4A+o4FWkZLCCTSKcU+5gkKwBARMF5BT/EelmUFHM5ULABaZC
pbNjk2v9fwLqGwSGIMgXmKQpdpoJSP9ZIT6c148mi9tYxy3mW3MIczSXYkDjDX3s
c08RU2ch++InbTL7t7kvx/lmbkQ4bVcMddoqDHtQBUrUjbuK0Y8boTtJ8tX50YI/
Imkp+eZP14AIZnbiYT53ViFezuLUiFTvFXHxQ99bpQ3k9Wjr+jUaEg1Zkzurx1kX
ypEev0It2ysM/it7jtB51AGUuz1UScmlt48Z7gHBq1Omw3fsoJ6N0o0p01S9bjk5
BX9jcdiNjlloKKUEKsns+aRF7HzlaSzSbL7s3rFAtmFbATWFBiwchG4EsTAYwS1g
zq9aI0JA+o6CgCKbpsahENjUc56A/2Vsw7b23RnOccUyU82029Ok+kW7g4xxWkyS
Za5suYCL35kepM0Y3s1GcBaLuvUcfRc/yKUAmoCotDn/qJR9DHXGuj6ijIZjUCIj
ZQcjh3JxDJ1n6RMDBb5rVQlgpVKCbAupXpfZs/Z8UVms/mR2VCXQFtxTUFQW51uE
AKyhJaOeeb0+C442GgK5KDyn/shF8y/aCaV+1VSs/fRMuO5HBmcc2wFeMRBxNbIS
fYjrF7/1Csb8mWkacOiZbAYaWg+fqvac7L2aapeLSXVjlNfygiEj08PZRqmefde/
eTQwQJGTAhp7FRMHj+5rEhszFzS8HzX8PQfPl6oAPygB9k6H2Oq1cU/cuYfWulOj
YoxblwuiEPrCCKhGLjZEgpL/R7ZvKLMTgBk145M+metKgeXaYSkRvM9nDYhv+Z3x
POd6ZV/iqXlxhYzSY5QU/IWl+Kkk5MyNmlINxGGd9ctnBKISJ4b0YUbtV02lG/lB
+UCNbhHjm7pSSH8SYoTOyhu3CjNILSfhpw5ZkBiPxaj5W7hVco4m/8/d6T+d+wKb
wB+lcwB+gosULvYhsL52ELi2ruVbBlqjmaKVTYxWt2e18aHGlkXo/FzYqxa+JqPD
HZXYw42AdU1F+R7QX5mg5F5uG6Wwp2YTB+0FoKDnEc4IPqzB+a+MJdNBmwPj636x
SNx4ICWpLPUn9PwncJ/TAJH5LBAo3xMQTpiRu6oM3DaKGWL5LTXdYG4Fde9AYdeY
5gLgLjIpFzGF+PHQi9M05m8UkZmf9+kRaEkT/xp2rUZb3RaqACcIVPZ7pk568D2n
zpc21nTTrqOw1iRJVa16znyrYKmrR7amOrD2XEE/yDiCoPpzuKaexaCfNDXCUrja
1uoCshYEJyN9fgkEu29vmY+vX5RzKWEdQ+7Rwihcd8S9hpbTsxsbpyhq6EgyMMtZ
pNu9Ur4BzfQ1RSpvfX38Vz8MzJlniHocF7mNN9DJAXY4xz1O+kk3BscLUr+a/LIv
QVEdqztkCLjB8rBCSpQ3NMeuAvQ6t9uHBwyTgui8f0xpok66fZuyQi8it+taRhdP
1ijbaK8GSSE0vwY7tmy5eyXKKzNwtvW5emhp+2u8Mm0xt6p1x3Hj5eVVx2vYOxVA
wO4/5y4Z1w5EA+xkpYsyAxKQMTfQ4EhE7GmYTdRjEEHpricDx4chnxAlwwgAZ10r
8NGLH206ouU2V78dgdlltT8JesTW7RmYpFEPuEPPCt/j4Ko1JDAIzjyFlZJafz+B
xvZ0CYfvHN9KY1KU6vQWmC2Il8TPqx68VIBrsY+6mcaqrpNy/x+kiLoJ94riowAM
eS7jVZO/asSw3C19ydw70XfINncs69KHUZ8A5uxWMWwsyVqudW+FrRSznZs2Bunj
7cJvX7LEHJAiJZMvpPVs8Jk2Zj41oS17dfZWIFt9blV/+M1dghw+VT8ya6yd9c/Z
wpesjmg4Brkq72rB/3kELTEGdVrW/1nHCgOiKPfmJx9ktfLINWQ+Em5fqD7qaxDG
JHmCZW4A6BFX7jqbdqb0yEnjxlazYyXj1sRiIh9tGFJ5SKL4Xn0XY22Z3cbEWXJd
r6GkMvHdEflboIpD/e5ZJiD0YEDsMsutbJ1B7lbPv4Lk0KW0Fi1goNwWC7foUAb7
iN9i9Sp5Bq32obf8tcohdjFFcP5m8VwNU0QuOcj8yw3rqgZo7ei6XqETAAvSQ9Dj
mAbY4P97OZ6abWcPtIDPHp5A+G0QSx6BIg5ApkJUHTcgi8tjz/uSPt5GnE0M5Xxs
Z8as4q5HWHEE5O8qkt97APVe+z7Cgw3rs6alDd2Zi+eIYNEbUoohYdeerxeT3j4S
D4vzUSGrLIxZCMg1dHk7Pk1oiK2L+GCsd9pqBpy9yqPmXCrVv97S9d82y9fmZ9vC
O+judB6YirHZ6YJBC4xe2O5JuQ7KxkiUFhpPLAjzPBlkgyxyD2JKQTJM/gNgXICL
qQfhDJIP4p8x5V2RyOesWyycdtfqnlvHKYR9hdh6kArz0bN1A0HeSY5pVel7HP/t
oV7Ofro//C5DDCyt15cgMAbm5jGdaHenH+Q6S5ddkcrxdIUfj+vP96pjmX8YZZ4Y
lbB1/ze9C9P/KKjmYPN8lPJdBYAeU01WkH5tU8N3bp2bvl4xuiJdeWin3Qv8mbWg
koxS9yiQ+lMYqqjAdz1JwRXrCtNIB1vBwl41ZQZhYFPU+KQFr1TdIpQOeCuov2pm
odvMG6eUrHQ6XbkV5v9aOp5sCTPD1Fq9/QyvZ/YihIai1VJdfohFSaEQNWB1NKtL
OI1ITpnwuq9GJUEnTZUACwuZSMBS9piS5kp7LIdbVuCPtF2fo8DNOkupJ2Gy7Qap
LJI8gU3P7O7H7NQ46fFJmZThPI6XeZZbQAMuxL6mJqLeDhdfkDDzJ2VT7M9bkkNJ
lmnlpQ5FZjUaqLh/2TZ/OMs1x79P2w0WhSNia5LCDKIiws42kJ9GBuWmaTs5IwxA
UO+TMlN8y8f/XmZJ9eqJEzE9rvxDLxGADv8GLNx2yqTCrPNsyMQaIXp/iXx7H0Mu
hOoa3swPCjMTX0CbfqQXc23sQDiJpVuF6tTi3OrDoGawdgf5GEzOecJJrRaWbDn7
IzVe+4841c7XHRUAxCEut1z4Lb+WB2GjusYOL4JEKPkmeoZsyaIqDZcfsD29mEvr
Aid9zG9uIjDdwkccnynRcR1/sg1CJ7XmpWt41yAdXja08hM4sdi3BRoky5t3i5pH
AvhycWuIutE5VfG6eoSrLh4QQf3QfvWcGzL71/CTEXPQCcz5BZTP3FvQHlmciWL2
QlsTuPCz4zhKtO+1eUefwd+lUL2piv7aGqnLsQwshb8LenSO3aJYP/yLNalRdj7Z
PD8GL3LncMhMKmVyckHIhqPIQevhIDKK6nFxedkmqirQxJdbJBliQzS2og5iLWgg
NazjRjtfV0TK8Ozks2Gsg8eggNF1L9qV3RaSgMTOJNcXdB80PKR+NW/Rtn8YEbQY
BYTW/aVrBEJUftAZNgXEjZIkLgntuiQbA6nyczErrulTkkeC0APKu/SXa5LLF5eR
ZTVcY0Maqq7tklQBE3yBeSWZmuk7TUaKR5i9AMXWKe7QCENm38EpX4bjTirS+Zgj
TG4A6PVfIFpyqXRgmM2xYw7q2/OgtGGNMjmhXWmQvQjB7VL8IeCsrFQnDKIjT/az
6IhLtrqFknTJFO1VF9W4oI9Gaw1zFj+tyME22PEqdX6r1RS6jI7MgNwzxbqCv7wT
U/6EUXo99rxCFOG1rl6RHM6/ylwpdszZmzgwx45XG9g0EhfGQRAwnzMrEEmrQZpI
yygAc7a5nXLqAfTEUXx4wyRspf+aWKLxcua9/sasBf5iBoUqwtl3beyW2zMg7t24
AlD5NP+fmsEnDsbGgIxlsPJ+jyfE3y50iKzANgyVOfPK9x8bTGok/HW4EnVlg5Lu
zyzHcOY2dSAjZ5EXV+hIvzy8URDuZhMYovP3tkwCXQaLzrEWZNFO+u0qDEWbAXZj
Sil6ctOcIJx7KzEj5AvTWWtrkuCSCdCjzH/sIpZb8DVX2QM4k8TPq/WQ9XVGOxVM
RRy85PfPwdpON5Ws3YxHIw+MNYlrjsIDRnoATGsqeWE+0u+7ZHZ1ByYQM/o6CcwA
cIFUNcvP8MiGvEXOHMCapvszuFET3+H0K6/BY6h1C15Pob9eVBqiotutVLKGk8ok
IHJPsgcsAJW8dXt+WG9L+hA6dzQGZFalKaSJnEicTANWGSX1KYSo9/osY8nE481b
F52DN+Qt8EAbSsEWXehwsUz5oEaweLI7oI3x+pt8Kov5KolZhDoUC+RSRlqRFoE/
1L6IUgJCXb02R2hT/6QoEQGv25iqbmZZPYpkCS0nnvpR4ilCGWGf8lMqWcRRT8oE
CmSJFhprzGUtOivrfDfQ6EJTxJSWUZUM9Zx7PDrgsq8DasK1+BMSShoozFYqlxXT
/rSExtUU97Z/xygAGXXO+zbTH1Foh4zjVW+Qb71NGMYkk/NjGpl5Uh2YyZygC6BT
N97zZTW6Cv9wOXOot8t8z47BovQX873FABdYkZCPjwSnxdY4LvV0AOJgDpuhLr85
a7csVMw/X4DBaauAL2n7fF+LGOTYc+ZJzWP/SZGAMUQTwepLl13b/UMgxhZUynCN
JxcPivx1FXToTFvPZ7BCYqz4DviyiNEkD6MDMIVcYcjSaiQSjBH90EuVknmL0S92
NC57et/9DjlyS8lU3jKpS2Tt5uT8PnSHcfdtpFn++LgcjQHxt3DlaYj2diOXGRdo
cco31oJM91jsDgD8G9OrtaDQSfzf0wEKIsUp9mgGVPyS2fBNnZHbXegzlfeRrPIt
0bvwikBxDaB3SwIHYPpdRY5QUmFaNbAretsEQbL26LKD+TqjlViJA6d6nkXBeKzw
wqwTnwqlNTWXxdfr3hlazoIUVT1IZPKbwBrrisISYU1js/k1pZgcIaoCFwNWPnda
PIgKBNZX0s4if0DAkFNXs5ipjUq30ARoCa6L4Yr4w7IGler3DDr6yP930K85iUNt
y9jyw4idC2NCmhg8KFMy4djUtaveSUPeuw2x9Lg7ZSYQw6LfhlArUoF1l/jhhrjv
sBUZx/RcQh0CkKyGgHxMz0I+sEzzw8CtbrM5anouGKcMfkAfIdjkEnEFBV39Nv1F
wQAEXZeOHjQRYcVccb2KaLO37UsdU6DDyAs/hpKSFUQiljZ4/yg+gusfYIY6r2mn
o8vpOVFbUbDrbHGehR4JI0Eh9RwHY/wtLS9Pq74QLDJ6vhIQ8hCHj+p8RMMcIjUu
TjPrIFDekWqO3MStxxVmH+Bt/v7Do6cQ66Yc9PvnKseiPbbyJk+SOyjpKIHiESrQ
ENfK5xtMMLPMMVm4pENhbfZ4owLnANA0VUqOWUlDNBbKNRHRLHGIS09ab3Sw9M1s
oQFmox+vgaVYHZddltI1Gdq1ONVNK5OmEpQxcwSrNRwRhgs7heJTGF5e3xV0RJ4y
ukoMKKzww2P1gn/cEMo7s5Yp2QIok6E8SRLxOovhctcRn7udywQMtZRDQu0+uHMV
UVTQihHW7WEfJKOLtueAaSj/m2L/+LQsVJPgYgcENn87ZSQEvSEavZbAdsPIj9sM
YMeQH4AVT8lbcuJaR6IHyBOpJYajep8J5OJht4CIyt2NXPH19KNvHYoddrxoT1UQ
URMsPYB4gEs1xvO/WIJz6HgOCmSjUfE1wMHDkWVo3WPsK3hqTBFrnPwpVluiUsIX
684lt3WjFCnw+oz8H42efhqis5MvA9Dzys/6jo4kQc4u+kaNJSK8wZHlQzoI9res
XUp/+ZSHjbWIAOGWFeqfYVzP31W1gTXI92+BhIribdl7F1z2milWIwttEfdc/kul
/EInAcQparRQlcm2FxyyJOvdOhoT9FvF8y3fa1gy+K2V8j3Z6wL2UWiaGJ+jeSBw
p7EAD4/xvU7UiyascnQQuwGV8+MDXhw3LJY3/bATpFBNuepsvNeUmZrbPo9d4XoA
qDMi6K9KJLEMc5R3feHksbVgkDMS21tvfCcIUFsOXg4v2q+HngzA3LqGE0LQ+Mx/
IAbaprDj7CmMyEuDyJqnfMm7x0saNhuIvywgYS9ZZ/6H+lQ4uU+hgdRT2+sFtjm3
6Axg+vjh/GMM3K1aeCkTLTHqW82xrxbkKojOJlWnleMLoWWhZFJPq49Cb/h0Hhup
MyFJG0ZY1zxfOthoLiFWD9hqT00ukL1IT88bb46bgS2fj5uGORBcnHSmCwPib7JG
3Jh7jpv2y+OJm0KDIgeqAqliE0lkQNHurH3dC0R+JcsjuHAuzHOnY5ypfz+4xHeI
vwDweS2x96X1gWEIZvyD/S578tHv8I+HdEGueftSAkJkf20fCEcwWrjfd+6OyFrI
U7Em6k8oPfDzvhp/YTa/h7bA7IxBS3gma1sc/6KEowUXnzV+zhIHjgR5LhaYU5vN
Fsnj0jPqqsltEV/yAhy6KQ7Lb/Syhy6VOy8pmMc+5cTPU7FA0piKhtx1FtKGoxi/
gnIcvAi1/eiXm1bOXPeTpBzr8lBu7sxGvnw8OpU7zDtcLgoXZ5qteNUugRm445C2
7e+skvpeICJpnNax2kw130Mu7ZaotmepY5wp45lLZOfGR4B8ukG3aRuiiDPH3LAd
v//TV+8S0cZdv+KLicDy42mKPSGRwJgwqiSghR0NYxbiOIrJRDN3/ctO1jVZfyOd
6LY4XZZ3uQN8xVo83+daD95kyFq9t8IGoqsKRcpbSVN5aav7XHlu3CRw4cYP7hV9
JKn6Mz6XuVv/bLsw9HzcNH+YBS00wxwhzUfbKKa4q0xQpziGhokOwczfp6NHjzXz
AmuK8evI8vKnrfpqfVKojMjMcIKzW24ClTtILTM64HHGwqOkMYYn32uwEqn45BSg
OEJU8RMS086y0To9xrEXlw7KQwhf+6H2u84+MY+X7sUjkwH4cz66F8yjV80tsahD
I1FLhPXLtb84KNn3g3/O7X7V7GlFtZThSSxudLXZmbonwzxBY3prO+uwxqWdv8xy
qyJQVL0DWZodl/LN6qcWU43dIMAYztf+aY2pAbmXwanmI9m9gmRp2NrJajRRMrDl
PDoUI03hRscgFDbCOq0dBdq1JInT59qTfN3hfl7C6Ao6+9yQrb3D65a0iwj5xEkb
D/XJ6c9BxQlcFDLygpaM44CmA93im4luP3bQWyg/p02yR6iHYh9fWf0iLfJ4sbwo
OLaG6bcMWwaf7910/HwXKB4sex0t8+Ttyc2+jvFuo6GM/4P7PwsdQQIS+w5C7lMQ
9tIrLZj8yQzIH0bNBoMjAmO7GGRs43yHz6HxkRdLCLG5Ibxpp6OZjG50t9v7w9zv
NZtugUkd8iql0gDvSGj+BV6eZXQadDjuXF/+ndlpP3Bp6YDvzPCwGvBtsRH1NbnF
tRajiv42QnkbYZwo7QmecfLaihwXyYSczaTEvm+FdbD8C8W59iYklkNoMDEesw06
kIHRYKa4j7KauWURKZR9yU8zPoHNU6VdxBdgg2fPg+nehgI0uXaHpOiLXL6AJhKk
VDfzOWiomxUKik38Q0OVxVbxJeMK2dWbBoPwJE7d0nvuQuEuaZjG1i499ShSFdZR
ctda2wZUVymdVMU/lcQhLajdxlOcJKh0rsCeKt3VHugxMfgCNoPhZqkOyLB8q89Y
SznHaS1VruSbDuXw4liXFpp3ptYvdkyDKaXaDspAMMs9Z3J//MKsXPNh5BjDpBgX
5YT9GOE+aCBRfAbxWfSEdsX3wEmdcOW1abqF25d0mW/cY75nf27rCS/rhy2wib5O
epFXOUun4tIQB0L9SNU4rLmmRafXFCbma15ierhWmeEHjRhRuLh4v16perUZjN+Y
B/rYdsWu8AZMSRFdDr+v30boqPP8SlNSgqmwuap2XDPu/3yhgtDnJ6vhR7i9hvCN
ue49mg36h7TSK5YbArbdgCEaRqxDDUkbEIoK7j0XYT91c5p/P5gQGLiF7hZlKbKS
p8uepCeEEA7+7hhsh3o8oybcASQ1FKemlN+UhMZy9OYmixCSJfbYzh48pdIWV73u
3JKdxrObmeSxP063Z7wItpM6/IcNdkM+V2qtPfbCJKGghApkQdQIuAelEPBnfn0V
S5vElRhOit5nlw2ynCrMUb2Zqi6oVXwwqi8K/+rxbisD2cPZZW5/IPWIr6c9basm
0bSaki4ahNqGXDxEZCIdf+rmdaD0+Fq0mVqpD2wuddnUdCjEhGdsW9Jv3r7hnHTI
CV7Du1j3jxHnxMBptTPvZy2N3Yv/rXOE8jh1gpsQsDP8PfMLQGrY0DFXWSZzO+9N
u2LYZj0Vw65+wyqBEZ9ao8lN4cnm5D3FtGRsPjHllRzxKVcaAqbdD80jHLpSll7v
h+9bBw5UMJVUP+S6MVJsLzgNp8T1JqgrqHJl+k3vsMnOnMFaBd8ihI8WSwjCd2Jf
L/h1adXGprDxZrg6s7JKiJTgc+o/c6Y1IjjbgwMYBAf1MF8fIwpsF8/+NRMeVv2Y
V5LOQcHd8SFbE1wJW0zGIaGCHv3RPf8KHJpafFJkXLsB6HcGVJV+O83HDiavb0BL
73o9r8a7pzDRvbuDHG3P8cpGz5Ch2JdpGVHpMxqVxr2fbLQtdM2gfm9BcKHvZlq1
1w/E97Gi1b2HalkoIWe8lY3MFXm+yn9VjyXes5vW8219jGur1q7sFyh94O+LhkZ/
QHt8KiXB8TZZKUt9KaEnU0qucrkl0b9ESnAbsknwbYhBj0NZcFx8mNembKV/Kggr
NLSi5AYj2ubiXZoDYh3jq9UP5xD0k/pgdOCtBABwMs3NoxoxyLVeymeJj1AGPcQD
s5lEIrd+9kLGewwKf0ZpctG+WBwZ/VVlmxiXP8Keo35H9k6LoWu5fPzyOhNfK6kK
9npJV8Nbtx5Ml+iSd7VjpX+giZ5xiIMcpsdHcXNBSEJsizMC1RGTQ2Y6dn6tS1nV
4A7afWNCFi6m9ZzyzUiAoZpTzFkQg/U8bOJxG6SxaEiJayrz3vif6X1KgYSTmwxm
t3G5qbGgzgOEzQEU8DSPZ0qepxJPq/DGnms8JvJR2HbgFPY1etXdCgrF80h1E2jT
1rNKoXkZZMMoWrtDwafJkFf1evtSTBDsYeUjtiQOF7lX80T0AK5DcHw88Zw2DeCG
8YZFYSG79Uh1JaZvH+ahn44D6VBvy/zWV/IbHcVHlJDvyglWfX89tQZuA3S8TpRs
zkCN6NIs1JI+jmoFN+BkhRNEFIcH3ddO2DZTvYSkcymJM+bzSBvgkepW4SMELELd
RAkgdQgwyUDJbtCsBUSEv5vmy78r9NlGTUcdhWBtaAx5mXsAhcVHuT1Rk7FtmkK1
y1G2QavycUhO8O8yzY9TZrBHIVDBipwAsyV0HVGJiriBx3XyX/Lu6lO5UYO3HNIl
hg/NCEKLKkuKZJ0fEkxPbtUOjkkFn3eLJ08BhSyqzOAY1BOgbQ0tqZaqVDuht2wo
EpABXWsJCv8ptsShUzGs1/plrIanF+HolXc2BN61bUhVIfjB9YVlSC85Sht7dneX
eu/wD5Ou2yLhMJE/PHlGZYfBey1My9vOMwUSF6PH4gX5NGeKOZ4fJFDSdbuBAtx9
tuj2+y8+T8m1cAw+QB0to1UB5KIA9P92fHlgliX5dHfM/TJrkIjjrLKEvV1xMjU8
p6GSY00YpH4uVaNGxECjHK+/WrvtLgkZLcT54CULpklA9/0mcUvfEX461U9Peqwz
kH3MnGG6JKIihH5tXKq9uBDKgzlqY8et2QjWUbC/FDrePvyfwNY6gGOd2rUNSr8w
Dko3ihCcxO5cutIakArclk+c72M59QSFFsSdFKVihWBspQEclrGNik2XM5rcm0Qu
ccYe3OT2e/C8xyRO5LJfY2kIxk0w555RmuIgzPNvmBuvKwxJp7RvkhSS/N/tPv6q
QypJKh1D4ll/3iyIgO8X6GF+b/hMKF86SbDXxylwZsjNHJcdxGky3S/RtkLl4e3F
EyKqOgTwDAPpYOKG/XUYF2IE9vLFF/GaJFkO4ezhap/bWj5u8wCJVnZzSv5rz/Ef
lvVYciJ/yOgFykRFYJfEYYlaMHy3Pb57mBmkKtXyWeYsHeDn62KWWYf0TJkNMhpT
K6E3ZcMDh9Ij+T+BlyOJEoXEt/MyHbekWMH9j6dyQR7dTrHY/VYUjmxOaLD23Mtg
bUyNuwKBzEdQ+NMRHN5JFmNYA+eq3aWk+Q+0vmAuh0L+U8ImqIwosgu09TjGm4mo
PtwrYO2RG4coDsZM+p9WH9fmKQjq5numOWgldLq3SAeY2tP/DjhojGqUmBOs90vg
J70mjJsZ2JNrmCiM7q+1/jygCCZDO22Jttzu5Vbf6n9UhUJ1BDLjo0nSl2KiyL80
pPMPhZPZck6WIDutHe0EaKnLPot3MB48hUYvnMO4VyxGTMMs+G+Ijhijj/yG22Td
uzxsvhdI9Kw4tn0p9Z+PPKmcnWpMltOZjS9ViUXh/WGUKoJYGxrnJYxpEbN0w3Ha
cgXUy6eHqO19Zrf0shrgRfkwRZiSt1zrpz0qUU3Sr/tL+dzys+CwCnbAPEUSeIpA
M+79AbD7q+uoZsDkzEvykDWy68BhEhWN8dG39vWSEmSH6E38pS+2tKCnQLYCOw6V
3aAosWLW/DBosSvcqA2a/UjSJU8fk0OZapAwT2ZcDZkka86AffF0MVYRqDeUBQA/
N4/6zfquy0GVZdE0HJFRTZ6WfgdXlJgIg0ndxFqIitdNcUvhVex107/iyT2kLCXL
mNvv/mW/szsaIR4wti7VSQE8xSMaKmFiLt5FN8bRWnXbIYwW9ID2dpYIlOnG8ksx
LSHk1OlMsMYAvV2Km/vuY0REsE3DOWx+pUQ3zM0qi42a4d/vDnNl10EkgvE8HnWz
F2chUeXCXR8Ka2VHgFN0QP8nqCDRw9j0hUnWLbot3ED7Ey6gk4nYInPwjNZ5bUi3
Ty85iIB5QdRKJ+KdzB3RZxvS31n7X4if3dDVz84UFZPNkEYwVd5MRbOm/FZ/2q/3
jobfHJSEi71p4GE35VD9ey54sq0zzyVIGhKspRxtkr+7IeS6RcJg5TG16COB8MFq
/C6HV1k+zSMlhYOGwSuFz0OzTv6C3/ATZzYCk+wh2uH8kySck+SbIfLW43/FJPpY
iTFV65ZbrFf81NiAoTeoQ1L+n9BuVV5Mo0LROOzlCD6X2ar9Ky+Hly2EMB/kWLYt
LnumFBQ5S/6h+l+kYkk4oYinNFAIqZLRfNjeQZ8XcxyiTn2uwsfdnIPhymrVjwnZ
4Wx6fuXQyrYxdk25ZhQETbv06bVcAsYRgRXQWboCn/fF3Zw93ak3zVuqmGdIJnC3
Mb5pAYiF4gGnhCltVGN2fqVqbXaKLilbHPGU05cGICR9xcqPbnp+QQIQ1jhGiwH0
zyiFz3MHssLc/iRr01V8Ry7R/AOQe3xn2Rmb9C7y6+q0ylbJHtc9IcMuoMmZ77d+
exDAo+nelYUS4dZMRU2aDGc4gYXIpilPh4TN2ouUrIW3tN56d1tm2AeTs8i5Kb02
wCLdt5mahrn0U7rOCqkUWlXNrXkFXicxXO4eYW5gjiGEb7alIIP6GCGX7NDeKDDb
JJ9pgwzX7hx29anrzVMkwSEIazzQX6+5uD6dPsP9z2A3cv4Ssi5tPqwOJ5nO9aya
PR8/aTSvBB9sKcsV6RWCK6A2Qij6mz5slNcOaZJ2o+BoGYtlwLOVXFusVyl99ztt
BO9UjpjdFGJlz7h/qTwY4Ib6NmlTiWVKjtpL27QALfGQhJLGUlxznWaZ04lrk7TY
7UWqpnrmZLIVog7Sfm77PpTbxdllfWzNfdFwpWXsHYpZnWQpkYs9ly2xeDYumbPR
vinZ5AWtI8treWravFe7GhjVsSydxBDARIKVaVBoAAcukH97p1xGtL1lzhS7i7Az
L1JcSTL9vc1S77sk8rXzrDuhcKSOwCfOE7nwSd9GMRU8nmDDE4eT+C01nu2ZmZFt
bHVxKSuyY2Nr7Msgh/Nd+84Ob0aB9jtN1K3itWwY0eK0VbHJCOYx9TAHQvgV4NvP
LlSTlAOLpWcGp8Cu6t/DrFBWpzDR+5XZ8GP5/O/qAcS7Htbu8JZqMMcL61LM4pnS
vhLk0wzzVzmdtlTX9H62NjBr26I42Irg3caTncveDVasDyQXE3vW+D9h4SoyJEcH
kWk8GWOZaEDQuphZfDvkQHQxdDu3wxMs1FQuI0Jdl4qEQAmf/Do4aevZ3eokKJsB
z56lgtOMUUgdbvVq/V+n13elVXiiqhpuj6y23Ks4IQlaQwoUMgH21KmduPb0Ajy5
D1p/xWgdUr6WBR9rKJ7IcZe3KfU5fi6Ep7RuzZ6VEQZcjeL1FD/A8pZZZ7vvCNPR
d4mBaQGdwqgKiEUbeGZAblHpgLWPSZ0BGgEpVDnvBBJpMH4GQbzW0b+IDFxgMZIU
snA8vmenF8QIkCdlicpL4OuRteHreRXXtJiP1kWZY2fmDyvouQcrRwyfoSp8Phhb
yHkfZPNVXL6Uui4EGpm4spIkLPUup6qIVYjXxZBTPByN1hp9rjaYZe+ZyyUvLXKo
43NNe97U7PWmBFxib2GI/Dgyv3bYbRqpp9MfohhfCyJZz5xyfViCS4mrEnQW+YOr
XT1iImGNsPIj0iwpTCa8U0I56vbguOX5vEaweeFK+50eiKq7DzqRarR5nz8nHgwV
aDZXDakXrhAno2dzuUI7/7WG7WVWGJEoIHGkwM0nxIT3+bGg0M9PjQBU6fcDwBCp
w+5jFahlN7aeqMl+R7ylkCqf6CuRf0Qr8/A3bK+Odp5i4NG8UTCQ/ay4bbNitstV
BcuhqzSL/xNOxGtyjRKroz54TqBEeturmfMHDNUJf7ioizTLvTCuQOGYPvr2Y+R7
PU/yi4ackJNYovDwM+fz0JrXMk7pJH+Gq2ubl/nHurRu89VgKctZt9atPNdvsSYx
HW/CIxyE8cUqieEYOvsiX+WY2PeUgYLwIuQrhMsc2LrNxFfz7OKqxKrO60NfDxvo
7FiGAt2k3pvSyJA9qHztqrjyKJLQnlOuK6r/jjFPVjj5oPLa8RiWRK8GVMz+3bAk
QUOi8zc5Nzkd0iDQ4zhAnEOFUeWfTi7g/bE7+ey+M2gATJTp6PtIT0wX7NCT6blE
fphewVrXPyl9MzxDCcYuAk2pd3HmpU7A+wfEzThVhzly+BjgFXMXgsEor9conrQC
q7+04uAHoS1UbxKdkuJTNbX/bHnX1mbMtrRDWwjRaC68zleQv4Tdrop03K9pjqdl
P+E4QXYHwPCc/khziLujo2US/LxwI6S3+1tRVCCxsrNfeOJsj04PpeDgTbLCKTjA
Rj0z64jQj9FuRZ5E5AUdadYFPCCK/DmJlMLkGbYsANwdzjPJo2ozfhTD7m4TUJ15
Dx1WKOMe1vnazrg3bFrJGKL85LgFw59Y2CRp3HLl1EvPz6+wLmhnho3xhv1pPVhm
MD0gUr0Fvf4Lu1ekc9IRo4I5YifzEzRQMIS1B4DVgIg9cPP95v2Hl4nBFuRJ83eP
xZ0nhr1BnMLaico8PvT3KRZHVXiDKZ/eXZR91OJPtMRoPBwvYtbCOuyKS1A9cXKo
u0aSWrHl8RPzw+F5LRYREhHElw9TRw94BILCz9gbNFgqj6wOf375wWgv1hlqWUBS
g3uc+Mg0U6AKql3iI3/BHTGC3e9/OKjKN92vWBedhZWwFeBgtmLU8b5TnBR7zsOF
IhiNUrqptkmrcB8qY3ZhGl6fH/gQOs6nUCoCjr3YembvMGSmKafA3mbsaxCWlNnc
SRMDhT47FOEwreJFPKfrpsg76jkPUUl2K0+gXKkK06hMej9vb5gDamr6fh2vbN2X
wtocj3Ze2+9yxbzXRiJr5XOc4Jz15/7IrbZwxiAaNbhT9vAgq7rj3wX7DqKze7vV
SCkW0il0VaEAaOZXmIZ508GFE7dvADOw6mabOncLJnStROOsI/zRTatVgkdClMmm
xK7UPz0xJKMBX3f/yBlX+9Q5ZdRJik6ACakqG9aYnZ0c4s9JuC0gW781/6Jw1E7A
6RCQy/Xw6WktbTQM/pXVfJj50rWDQyv5a7gWpBcTsvuC0cPvqHKhINJgvPzHZqMO
2M5weNmNBa8kRw+KoHqZ5yfTvqzr5MWCTQejgtjwKhdNiR60gEMjySQSzBE4iduG
xHSQmmiCrQDteQGS03INOQslksSM9fSWa250edHnVuJYlqU4iRv07rSQX3AoZ0tA
0seNJt/DabtbFIirDriJeELzMFukUnjZ+mTMNyxgcqCZ6crch28K4lpbKWbgwu0o
FgQAAyA8gKKg7VvGL3j29ccq/QBvyJ0bglH5q9dmmJSjQG8ZryBBTn1N5XaePvj+
WtY9Uak15aBRwkKTciAoeCF3ufTFWud4EJjdnUJOHLGWYGF7EoB038Jd1NCuxHJs
/+L/yB8a74734CorGR05mQ+6zXZwRDGYZ6kFNNdS2ekXJkigT7qPKbDBccTiQ937
BBioKdINdcpQ/f/rrPcrs0e8i5O12R6iDcJ/MpfoelFBEPaF5/iLbRsiwuV4kHId
CskTL+mVEIhok59AMVAlwdCXwR4hqFw/m7U23P5AJPwgudslW5InKD9XX3Him2ni
oSwx57zl4OIPhe/uTT8lwvnX7CsYJ/GIWwnpcY2YWmy93qbP2UgSbcLIuBTHmyu+
iCi5l2lqTVSiKhn45nTH9jlrWTGBkUkbRllXR53ke2qvAUAPYN3RM7hZ45hSWNFY
M3N8jWnDzl9uMHas/Tq5O/oUu69af5ElEfGpA6iLpIklf5ux+9YN//yogRksuCZQ
6kM6/zTQ7xW4xgVxf0NFXjKKtpKsCROUv4OEnD4k29u/nxSyONDka3SZ05egH+XH
cin/F+G/L51807KxUXll2pSfdGp3vBOy63jmXtfpcxUN4gmfvKOL4FwDZrUGpFh1
1ka4N5zf2BnIft2Fe+Zt9skCUM164V3IazFwS9tug3OyCaXH95WijJegUImiSoTe
WJWL/eYrSl3VQbPXRw8fPxJaROqx7rNih5dZcpVpTUVijsT4XjAFEpZAomXQWJUU
aU1QP6sQXFGAN5QgeQSQ1UvxQmM5GN9bXkNFz6uFCZ8UhLpmUibhyTn+vtylLlZo
TKNHXCHY564Skee8Dodve3PUek7F8pxBf/3iHix9nUUYxPuq+vgoZ92dvnUcL/wz
5KYw9OdrkGM7EWDPCc6uhT/3oRN2xZXaNzgiXZmx+nydb3vltiWN2t2Ow6YU+ll9
Ke3omvvd7PjlKw9ehZxpgKswOldNyc6MYSJst0VupFv1A5s746YeGAYFIBEnr15Q
6EXWRQE51/E9giWybPdH9QycuSRbUxaNlURKm26amy2FU63SMV3FdK913QlnVtn6
kQ6vvJALBYIq7UO5tmbqj+rYqztqTv1erUAUWxFN1xFdHnZqvJvqrcwb6qsOag8l
oLDJbhphoTW2HkwKJUlp8/j/6FdWon9dw7cx6x8DQiOPY9V+Xl60i8zFq+uCNljZ
h6eCMLsukmXIpoMNVkaCEIMZ/tf+E/IqSBTDvFx/mpgscsNnK7ENkcNb2mtpb1fN
jhSP2chg4b0esD9wRjVfScolPzy9sKu/g/5yRTrlV3xDqnkkW4LDcSnfr3bN/Je8
v0ljDdAeZ8Y0kSpAd4jdMopF3JSbsyNyvaRRi3dkTC81kiPdEH6rbeFpIXZCjw0B
ktNTW+MDG/R2u4Vfh1rKGQsWwOlN9pWTrBRPTO0L8nEPssFJIoxQpnyDQ9ZUe4qt
H6nLvq2O8o60mHv9uTdADxfKYqckNgwhiesDgKa68w5zBFWk6DKUY/XKvs0Y+Of3
ONChqJbpYTMUxZARBWzTkkgW46D+SQmpIyJQ8u59OujavFws57cBA5bwwLlmGNp7
FfcnVXLyHt1lT0UJTgEe7dsz2fV5WTg31PyB1NN4hST+afBwJo7xKwcynkSe8zz5
FEfBYoM+xu7fjT5PywbsnqfK3yoZBIXXpDOemyZe081mbh3x7FmPQ6VgahTGEv/Z
YqZRnFHyUdnRGsYgcnlePO9VZKEYUY68kDDyTg+uwaJ33Jf0lXV9RK/kJR8gVjHm
t4Sp6jrpMXNVtVVL7+dqhVmHOheTlbZ83C4z/ktFa1MBETCcP7irVO4EtwMLAvxQ
GrSOsmja2Bhx7NbnCXX3JbMTSCn1xL0Non/QKCbyAhAEv/yrice8FvOlfBaQNpqY
TD+N3s0mbsCp2yNwx67WYonMBcpebUwQ7XStsDxTA8jtXSVghxaHjIHxsgeMqxIK
3AWdH0kLnIO5Cx++jmSZ4ErRgHdW5+pnJso5LmlM+AK4uFzSJWwwezvFzrg1kNL4
z7Ji/yNhLMjVaokGj0suHvHThEB83iJoB7fSfIkGJ2xnfFAR+Vri17aadeRgYXNE
mOyJHGEKLSaeiRkfgKa3vikY5QrkEQGjVqrfDZgCI+/CIHoPU9rqtCtkiDi3fsQM
YTPrD1i43RAcpWfktHiOlm3Hlt5zxwf9sfck6w0yQ4tRjrTQ7sZDv8DSMeh7nWp3
epyxoNsPOr7FJHtuEVdXQoS5+kCkNKVxYhmDyj+ztpGFGX92OlG5lYsh4jTMGcec
CwbFsjqpTqO3PdY8kH+ag84pTZqDao1SiiUtFWF54jsfJd8UMNDxrFp6KDaR3DIi
CfV2V8BZN0b6HZEFILKOhAPm2oiW9RApaRBDlBp12YizJSs2Jc6lWT5J1UZXC1NF
DYTw5LNw9jXP4CoIliXKJGf6r5fNjC5oP3bytjJr39oczSnDYPVSRdtUJuchj54u
L8owzArYJ1jTTUesL4TQOv6dVnThzKcn7SVLAcn75TtpZNKkzAx2sX4HQidVVXd4
tyVVxrtvzTOo7k+qaALR8aOkaAMdShpAb+Wy1W4SdGaX6tqi+ALee3JfQGwT6GgT
4EDJYB0hY0rSFySPefwwmC4AvjPUEiFiovnWa3mjOXx5cB+AMnLf2JfC8K0e3oKB
+IleNozBQFOFEFvg/XDsJ6y/TN0U8Brw9aeU/YJ/S37CibM7T6egMSzrWBDcLvVk
UclX9Jr2rUtxKa5WKlsFFvhSrUyuEpC+NtwwDJKY0hy9pOeReWsJTc4BzMKOcA0k
eS4oAJWDYiBQFA8Ew7lq6ckdaRc1imFqNUzWCGx0mSqMPRN/4cGOvYDV7Q3ErwLm
dcwvkw61WTR2QbXK+7k2WPGNiijCm+d8X1GHt0GcK3iJoiWU9VScWRwHmQ0WD+OD
/TZIcwWFK1cEPwQxrsBb2zpa+PiAgezcRJSaPBRkY4ZuaBN/U5pPUrkW02eLUVQl
cR+Ow29kfBqD1qT71XPIBRPK8O6MhulR69UnrtjLOfxXyW7eNaZDPQE8dZr1qMbX
6eNeWwQpQFCkoJIaSepTsKmdMp0yEvvPV9ecCJAH93C3rZDB2RzkWmtK6m2t7AUK
/MZYmQRH1l4D4SU+U5ZFA+0AzMBnD+XYjF+chdqRLzTR5TfDBXvW39b1OH4hZLn/
5CrJtBZH4OLdO8mw/P+REEC1KNoe2jZXjcT6qpdavsSUB80z1YyVsJeJ5MKQvBJH
MOF3ojfKsGcJrsAl8EsybCBqozASytXwHpdQm2zJfXPTT+PckOqYbJOuErZfPXrh
uGVNm/Z2W3YIwA9569QiTfeRMn2YrP/6m70N8gLWx+GYo1bOP3aSOZz9FVDhKH5H
62Giu8rtrzCXPgOXFqrNAC3HBp5E0mPRZ1vA2uBJf3H6wzB4UaikRKkBLbZMxC7W
D2pSq7Qrt5DmIb6b2Z2K40d3aAaHETIX/tnbmpE19w4cGmgK4NCRWrg+tfQFB7Cl
kge3SveN9v2DTODki2c+wuqSURT9b+nXQonj+hjY/+e4jDDMUTg6YIZvzIZTXACI
eOgfr/x+ky/Vka7Ad/EgASOCHDQpt7Cxu5TFBLGt6pgSK681u9VA3KogwcsrD0zH
UF0mVzgG5I39z4ooe2vdu+BVxzoDp+j5CqxqpGhWRraMDOw3tn67qW4I+wWqCEBa
mk8pzQFPZz6IsyivtyBWBR4CoxhjmSNActYy20sngeGmtpf0MJQUe3o0n3SGuRvU
Nit2JjywZIKZBhQOzU8OFlmSWT23E8lQOR+Bok5M9AxRFoCGUXSgMPSdfxRk8AAy
EeuS6en3SicsG7a5CixyTvkF0WRdcek6d9psErmXgFkm/Zk+UirpwjeozV7bHk/Z
ewU8dS2tS7h4ReyNrMu5kcPfJEeBs3jEN4l7/PGUfTsD/cZOCujDrgIR28DNMcVE
SmlZYJBzZtLt8aV82xXRt98FjVIQmDKrKl5czaykUSHeqRKF8fCfdY2qJ+PLGazP
FxPWfIcQOPkFnd2aw+fp15S6zfAKk0hNsCeG/WGi9bbwWEx6ymf+KGzBYChDdOHH
xH5Ge3oVZkCtBNrIiEBUYudxjFEmxHukJI2aHEkoAuWSrEqs7nXnA6QatcOp2ii1
LMrCgOwkiA3HhwOWklFk1yHN0LJcPRvIJ/sNl+cWkQYUOj7iz4QQ5RMWVekRTXhP
mDmhmXqko3sG0RdOOTkNH1ONazgH5aquUnXTKQ40XuzPMzbnOjmMPT7r3E0JunYU
1QVtqQ+KMmM4BCVsTO61UroM0PkzOCcdraO5t12uFgakeVt5tvHxrBJV2aqISzmh
Q6mTgKITXN+sXygVmx2U1KWP51cw9hkQjTKInT/pxPoJKk3FlVKhpgZlkAOMywRt
O4QvdDwF9XNYGEy0+lbTix4i4NsMPdnRehY7mxDZDT6HZG4frdzauKNptk4PB+qB
kHhH06JYDTuB7EaNmZJP9mQ7IYemi6X191RMxXTtlzLwBui5YDhFS4sRuWgjsPtL
5Wmpqb1Wbg3kCtpSLuy0RXH5PqGgtFi08kidry/w3yJJDhFsgMqb3AYqUa1qJcVu
UHWkzm0rGUwJrUYed48wfEMlcvFmS/ogLIy8dGoRFX6T+oJLXj5BorxedNcOwViF
2gxB7OSesjtnzoh6K7xndvvGxpNEiIMKLYJzL88v8W5/rvP5jarJ6sm5ClLQRNdq
vzPhSUxJYuwZRyW6B7eGlAfmI3dD0d1gkUCoNqn6mp2N+M7FPYeeBgSB+I9n/FH9
otukvK2LyfLxmVWqpCu4suB3J13bgVdl9ZfJZV65WGVcwMnliftVgRuPKKDyF0eO
7tB2H31XIYK2KLUoEbY/dxNAuYsgt5hu3fwZgyCliK1hQQseNNlg8SGfiOPAKYzv
WiTblYB1RSr+TszTk0SloLzzHJNk+hJdhkMLl1AD8q1b7VrDd4NkLOVvzPA9+uDo
2EpKpmwQhG1hiM4YZ1dSJaRUU+adtQbxsJ31G9aA3sCWMWWB5Pwz1/6PYqA1LrVH
b3k4F3C5spoadW8tS+NXgS4Q0UM8Gkf2mTUl9txoA2nzjzzoCGiPGe93R3s9T33k
7SG1KuM2Dz4zVYy/ZUe24DIHHpbCZx9qCxJ9m2eVYFKlnEW7+Rb+RjXa+R+VKJtH
9780qJa441VJ3NiKZhwAMmU7dWc59nwi1Kwph8c8R0R583X+Ic3bu4QgKSHtOJoM
CYQjlQAsMZZVRmPbrk4WHcHZmlutWmRxz6UriRJ7YWj0sypaWFJE2OX6ShrWZdCn
W6rWBdWblFC2cLlzbFeU3rL/aTrAJqHQf+9mliUd/4XZmExw+peD/dNIFX6ozLZz
qlt1MD+w/cb3maLKTwtpzGYHlH+lu0O9sbK4AgloDsctFyHOnTKbJMzcMM+FZ84u
F66PBh6C95kqu3zt2nQmAuUqz1RdbyGzw8Tcvq8rrWMA4Y7eiLFcS4pEL3hKkr0D
cRCHkvz0m24yxSye/liL1cE9H5A8kAMnMsvfStwg4J7o0myObm1ruVZKM2BL+HFs
kjeEX8UaCS9X5fsytGVPGkAd3fT2FPJ0cj2Fj/Ag5TKtkRBczvc7eotInfP18yRY
lpdOkPzGy56iaZFJAujFBh0KvK3PzlE/upDdoMMC0GiNUvX7Uby39xz776phzLQY
P3FS9YSVfn0YEkBoR9Uc/J3dLUaJ8sHim2F5/mbgFlkaFvszx1Ov8FLARuTFe+ZW
tzAWdOCb0j6H+OGdIPNnJwe4XLER95EU2knycK4ss3ZjCUSg7i+jAFE/jedEwH+d
505yWrMdAA+3hfo31WxPwADSYrDnGimTpzcugm+x+SneeWurmEj0a0c2404mFYSw
apdEOlX/QoJaARQE85iQQgi7TQUltemyhOeM8WGVGh8sADpQqWLP6DW94bL2pPVz
+FhxVGQjhXb6DZcCm3ELf7xz9x9nMrP0TSPUGHXN/Tjmpz9Ur7gYlNzNi/WyrjDU
0nuE6UD12sFCUnWx2ZbiWObGcLcsVpd6LUwfup4Jk1sV9JG/Z5KR3a6r5CfqW3hf
izZ8/PdVyx5u1/H5F1/tlG3JJz8rfIjPgsaE9RxXgXi0vLvyGG6+Ye9PzpW0mqSr
xn1Y+qf6ctTEemEgRIUU6OpbAGzvnH2wW9WuXXiSHXzhGLcIXx6g+YqyjeODHpx8
bVw/lVewaQb9RBqPSzjndRxXX6hOyBSLjlqlAdG4CCqZyvws8k4h8Dc7JeL/H65j
6651onNwSByYdLF36XBej//r1TwVhoAJ2oNrABa1UqPhmC1yFL9sKkcwcBHZ73N2
JZo1jPtYKnurdhtSivX469Q49jzdi6z+EPVeTTuWyB8bje91AB7p5R116NOK3sej
pZD+UwtGU7NVT6AmzeAcC6f+uDHUdMlr2gTtACORR0kl0u1SIcUcK0FVV4KSy35R
+C2HAXv6Qhu5oGV8WGMBJeaUwbfC87mnC5hKV2bVrazGBNtBZwmyUBfaIRxrw1Oy
IlyWMbycjFYUGnSe4RPVZnyhQD2Bl35UVkBFmiYhTyNmCv1rrUnkzBqtMRWdcHq0
I+p2fLTNaPryLpQLzfIv8fSuXb0SCaUaiPb5aQphgSZpKg/CqXsXoi1ghBC1gFGH
SU78FRf01MNEZWlKyL/iTyjV+/Nv80jzcysOxV5HwrjmpDo2CN1QDJTWz1RHhIWp
NXB4F57LkdR8x6Ux3eY6UR4+Ki5r5PDzmiwLgDew/zl30JMxKhvDguiR0CNQ7nyn
z421Sk+WKcyYKJDawUNU1+jw6FtiOp5jP4ab+rQj1D6wH8q1XP2kEUuhKJbJe3m7
+nnSUSFTQ1EL0iOxDzoRCA/iNCYT2coZpfc+8tjdoNPvrDZ2mC9nXVcbn2xtoNwU
ImHGrh8qoz+tgyM/LPKvWSAgVgc/Rji6Ddh2ElOooWRB5cJYkMBvC1jVAipssY93
V9e84uvISWHv3RZko5/eb9NrGM2pOxqLcVLVY38wp8dFds7h9HNI7MEG1O5WHRJ9
ITlfVYheWPSziAYJaosvZiJOofkuO2RPz48HcddTNfaoyKA9IkxC9K6gxiP9BGcv
SMZch2W/E5EnTjfrIwH6ZZqWlhwWKco4+j3zSBH2OTb0+YC0oamtXfKNOVlk14us
viCiXG7x4DLjL3U38Q13txMPKuX/azBLnzHySTOtyuYmuZVh1fbSpOTKSGJ/ZaLr
WZQOyWs0wzmXrGOOr4Kp05ajqCb5U41m1dm9EMqui6QBc2HWXzFUMfM38FFvVoSv
G6XNyfg4aW434ndBSvi+w5RL16E77t4Ws9sZSZka3C0uhYFze7G2N6QtwbBjaJZj
33xCb3Idf22p7acudLxYLZWYTS0yd2Q+39cBNFhiX70V+w5/NlIE806ltRFyRvRE
69I2npsTxnkTFDuWLPsDFPpwSW4TMroFGSQo9vYHbTYSO7sYLl/hmE0Ck+fCui86
HqUTGNRhxTE5dIbJ564h24Qy3CvLt0UEZ1aqYhCCluJ2KpeFGqQp1w/rlo+oR8B2
SIX+5xUc74ISeSI3e4HFnUaB+T6mJIKq4JSAkGjiwlH4WCj1pV9rsrq91E8pCIG3
xVyokWIItceOQUVzn2T0kofWLo42Xj9/XOiIkEUuJQp3KNNSjIfeMv+igqCJltdX
mK5UmqxD9oYpBNj3xVnPqRbhnlDPyX9ClEMq8KFbL51nmogE1H4Uq7rbyxPixKVS
fCfl6Dfrg8CVqIdc7w9wa6E7m8vo1VrEPosCXaC8AuJi0XijfbRFPJ4X9iA5Ih6m
4SKzm7OLCyZpb31HYoMIJcnYWATYhrvSy1ilwOwCYXxJoZtNu5P+lGrmdhHwjrHt
luGg+EN733yuIzs1HbwZMMuJfqdM9mJgcKfjvFEeQmPJvEftAtfb5LuJxdAK6Lep
PHKxpTjn7KfUIAsoQkZYE2J5pKWEU6uc7pKoDU5OTjqpAcSgleMiRXbgKVwTapdF
4bmpIVb4wyEvwPouH9i7u8JrQHadoemwTHIdeHXPyVe+k2IIys4Anpup0Qa0fiw9
ISY2D8lcpKQGXZMaZjQaQMtTPOSnlgGAWgt1V4i1b1giYFEZq1J8tVJ3Qth+7ejH
vSW8Ntyn5/d4i8oro8GqFc5woviZSZAiTDyujW/Uxu1TeK1yuyt5hTkc3Aiky1Xn
x4aaOwiuZtwHLdN+xXvXlFXdfqBLArpkCVk+l/Q4gb+cFbPGgElPa9Fen4fbgkhS
5nwguOdCrYjB+aPdaxmxKIgYoNC146EZvKwHXuzMW3OlvD5vzHYsWocrvfT4lsZN
/sU3k03J91NUeASlYdLP+f69p9IajNRnxvvN3VXxUuUfHw7bWT1iEyEZoiHdyR/N
6HdHUP29sSyd/ULgxjhi9/f3qsdbU86fTsx8WMpwavWL5S0dFc1oZrvcomV4vYiA
92zFLAVGQXsMS7aeVRCxEFT4ysDeZoTEnifbCj2G53VZQLwrpNR757K1b1pgeFkG
wkadagxzJLQWWkpKocNi83YZ2URn2ZGvFBxkfh1Aeran2bOYU9W7LBK6tKOXvG2U
HQsdxvvMvitKxvwWb2ZbaesdIa5J99nSpb9SEWNjBEXoc/zwlKrBvBzdQfIEXBeq
N0EnrYGw0PwNb+vGG9cG42TYNlwMAykxvsDxF1DlGKkIgxtK9hqvlHTsWOcn471d
cLYUH/0/15PPBp6xyA/D0WLfRUufoYdKkCm+AHxvc53v8tLcm4hK54ejnjNUkfSV
UdyKUMp5o/Yroh3eMKB08KVli13TGsYFYb8tox6+bcXhguqJb80uApHevPu6s+2i
343uMpqtgb0D+dwjFgD30iNgm4+K1wup+CNQd/DdQfZcRIQrxveus8jANEbjMKCg
07fgXDKJzv1+9R6vLAm1Y0upMPvnOYNtRSUYA2J2vLV1mO5L5SaxfDnv3sUZf6dG
V0xXJJtvnOMaCEf1I5+KBNM7lOGACpoDMes7W1uULZlBpz1hk4YyxMWkp/QLZj7Q
VpsL9kd3dKEMzty6FjSakf0E3QU3j5nvsjCWyGYpDDVIr9m+gcG+i8B9oNQKU13f
7Zvf4A8256sY6ytBeZw2DX+GFnkks0IjC+c+Ovqw/5bJV6oaX9RjYu40lYNY3qQT
CwivvqLZ70RTdkuMXbAzluPVpDcLNnJ/pSjB6tbOTRQbBcItgxdwGqay8ncXOcxG
eR/mwL2Car0+2f/YPJCMTlJ1tAIbkQZg0/l7ET5uourm5FDr4rQ8MPdgPqT2ECx4
qEW6t0JeDm/pyP8T9akJ4Ct98gE/0yj0BCKnDhYTvLvw2LtrWX2vI6XkQo+SQkec
++u2AgX9QzZebqif/oLHyt1mQj9ZdcyCJ+XPqsfvyV9dR3e0hafBlNE+Zuw7+fqa
DVWHaeL28YQVg/QE/g4MApVLzgGRx5FXX+f9Fa/wYhkM4TpdSKgiwiBCJvmwrq6S
0WEj+FOmS/xWFrpL4Lp6kXTIoWskyHLuPfY7QbxeElkU/+FdvsZfz/wVhPZZJpV2
8w5Mn/9fc9HBsEwqXpKcAc5XsDOzNx5fwXfjK1jXFqM6u2quLzkWjjCyhySCbMKz
kIWXsSK68Us0HQgoeuT9ek3UKWiaAQnRNfCqk0AfrtEk7lBkU1T6HW2ayrnxuit6
i9Rjf7D9w+FLFSGKmRtB0EDR9nGGvhr/ORx1IhFWgcV6J6/2UCmS6/AhmMHMpYxu
S+b9fGkuRvfTj9dSfnaTF65aKQbdLN+9ZV6EUVwEuToI0QzXYJhcwOcj9BnCDOBB
7OG+mMf/BVLZYmG1cpKIF5wBEJWW9IdxY4sGnyoWnxKDgcNz5f8EwLT/2vCt/5h8
SMJKdc9ZFQ4NiZEpofjQBMpKLYAfn6m7Fkylm8ZPSnvqvrcszdcAaAZu08OLl/0F
55fXfYvqims8n33kwQGvaI4N/FqnzQ4UwS6FdKvQB1GRAdOrlfSuwPxALwkGQe1S
6Q/UZ9MVDrt5KGtQAsbUB5svzFDbK/zeqpSqglIfasqYsO3AX03n3aSlRdEnkvB5
SEpdRA/016tUkhPpp7x0HETtccRQ8UjCcdIODAjA3iAUydcZlEIcM6/7tNz2n7Jx
dWB5GdoOotM0QJn+C3Fo/sbtreRccMB27ZrPmmimehf9hzRF8iiC2D1G8Hbt66mv
tbfBY9NdNjBBm6TjstiwVZjdU3kUqO5H0oRclOl75+Sn9oX0HAGH7ONbYemi/kYb
8dJIF7+MNeKpFVK6G7PxEwh2Azpqandv1qjwO4c7tzQTpv74Sw2TEpRn35ISOIIe
8F34ZSPONmN+oua7iLeQH10UFq6cwgQD7q4mS8COTzxBIBLXoDV4RvJqVWwCPVUQ
7X4Uc08UQHG4s5rrLyhBqgDNKkJVmSTydzh3yBFSoD3iJ7bieQAVDaxZm9qqwpyO
FQBG+P0it1la8WFiSJKz3RRX5Vrk7ZFE92qOXn4WZcM4NzksLxJmswletYbSeqKB
/8g70ht5Cj2xbxi1PX3ZiE8l3VvUArYlxDqjG4GpFjamPo98o24smhpXnkKajJoZ
NdpDzSoukDzr4VXRg/ls16oRL0197qIk5yCxb9pz8/s2eDsGS9gY+7xWB+xgeA01
Q5rKsPIUAApPGyIm/7KbN2CNxER9SGWFyxfescc8OfrJWkMTrJe6aGnC6l9LH2yP
zLmf2SRws6hmzj8jiqbu1zveivt53Ijz9E6ShmvVTAAYFvyB7HBFWNWdABTXiEHd
oVgaAUqNvce+tvZXel9Bxu0JaPKkSn+Nj5WfP8odldtB83f0Skj2dEGqpqAOx8m8
4HnJJSSJ62ILPV77sW1KssDvorUSJup5kBEgifilOIx8eSra33nJ7qMXbj5/mMuJ
/5e7x5raUJqLdfBZTHEeDxJUgVTpTi/XCiSZjlSClQ67/I3Tr4bUICJ1/MuyqxNp
91RkeNytKI9xtwHBIrewppLAn3EZ5b3pwlaZGMxRSM3TKawuXRhMLK0N+Yg0DfPC
xuzjKDLPBlX2eAh+sA+aYvYfksrhlGfeJGvnlwWKU1jcCKosWs+AFUQzouY+1D5N
7V1UHtxIy+AaxqImDxnLwzQnO55bUkxEjG32YMrELdG+gh2Hg2SBDu/cr344oqFH
psWHVg4KDiCMfP/rcW6C50/Fen8Dtw+g6ykdZOKfaAbPuGIFjTNDTHB4384b/pxW
RHQFOLo1VVbNLEwF7FQhyzNXngBM+svwU13DMA/dHc2BNNh1D6KD8IZGPlbFHzg5
T/bP6btbrBdNJ4D2CNlkADZzsD5PoG90dBOeTKqD6mDOZkWpRT5LLn5qAQoeSZuU
4YXVJ7xGCt3aKIGiTcsOZh05cVLMSAl/SGVCHdpz9xl+3JrTWT9+P6/JfP1PlJR3
JJNmXzRS0P3YbD+VVMoijgf7XSuuCSkXR1bhTjxGvn7OhbO1hD5zPpQ444sPmVHt
lbLwk5TSg8UZOlurd9Ltmjcf/yZMjU3HLlP2CHZ1aKmbb6kl/MlGrdAlj3CBv1mP
ypjlbh+km72DEwRSrcKor3fXDHPCTGaFxM3uZsXW3BjhWRve+DkOO792GS0GTwKh
KOmaHZM94WAeAW4+CC32GVpuV4dkpTeeCePx67ZiLLFwXBzONrHUK1stPYTBoOQa
RV4wzdr/5WqlxDb8JJsw6DHFhgWl/qfHXF4tvcYuFMe/MXtktg71xivmPW68wJLq
EUeuTN3LCFT+kgr3aPBGJpSRYvVPU7LNs1frnMuIPUsEWxVY208+OOikmCpOr/8Q
9gjblgSoIPNvnARsXRtadfi35cW092Pk8c72gTj3OxqlpNmnrABJcEWMtJNL0IXF
D8xieYGTlOvYyjRG3RNdd4OgFF0QafTVi4bpubfb/n5LM+DCU4CEqLLEmGAcMaup
g3fKOZdtkipJOo44Vle2WuKLCxfnlY1S/Lws1fCB15HqzSdc3EVv4qQGsgo9GgKA
5wxr+xUj+uzDEP8E24xRaurgMc/v25vNL9pDzQzLQdSqvp1rbOdR+DaiddPgpsJh
VyXKNhBSXGjm42Cwc2AbTz08mDOQz463dIyeYzgko+IVKzSRlgfhNOm4hUJesvYl
QeFvO0xyZBQN04OP5qLVacwx2k+BFf1ZfAzmlzIyWsXEHDjSlggAlsTKmMkcCHWG
euSp6GWsxuFwf16kt7Kn7yboL8jz0oe+FZib0r4yuoOsOh4v9cW6AA0wVsBeZxDK
gBiYJiBtEHaMmm1qMjZsTWVFQjvjN3H/ZNv19vlHrbf+2qSmi+NyLGNSvf9Mz+LU
Vn8jdvkog0nOxPjwFFqB0L3MSprcMDyDWKjmg/Klh2jfvfS7wmZx9sticKpYu8EV
cLndfJgJeHLR2SXWZfAvjf2jya1i6HC0kD7GqOAeYryxz4p7Nf/5nbgvbl3GM8Zb
mZfidDLCyh0MuUsoqhyZqGrYjXw7fmId5V4aok1aUk7iWZNO9yNInbJikReuqhae
lB2j1gj6ttVsJjqEaPIU2NYaAPIracgWGhi9tCzr4JMqpb/g+qNG3jdgY4dEZrgH
4QhDtxxH7PeaU997hIIaoCr6C1eOIGix8tfJYqOp0kbQmRy6Pr1w9Pg7wXkayqFY
Jn8z5ETePBlxfed2J4o7jiIMuvoW3NEeasDTHsKEDcLXBaQ3z8MLO500PnLkppBb
K808ZIOwVPXnBqN6DE/SQ6MgC1HxDUTa+Tah3WWlgd05Q0wgEhHw39MQCh8QNk5m
YeCMj06saX/yaYhhnHuOUCRQB5+oAP6hl3IclG1g+NpgUrr8LbXtSp7iIIYQvUPP
TzRXhnuZXvTtvMESGoXONKNXUXlPD5pQ1i/xk1iF5GM/hSEyaL7/D8tMfmldKDO+
J1wTRfl/v7eOdzT4Me7hdRaD4n2SRQ2qQaryGSX/hzCR9dccxhfrxkRV1kPw+cqu
5DY15xiLcD19f4GLVoWX1CBbifrrt3S4gaPzs4h3dQQs/YaD2o37ZMIqzEgns9gi
9LYQ6SmK4HPYh6OWKCV/0qtq0dhZoKlc5twBk8rWLw09tBuO0TCMMzyqz2+npr+m
xhp1+KuUqnM3lp8/fqx2wzoTTMVPhO/N4e17NL27MGPbqBPPwaSqLpprXhQldgXg
DIOKXpNe87H3ugTcKUOOosMMNM6LdNna6z9T8TempS13bYzEWbN380DhbVybfzAM
3JGRlKmPk7GBTQc8NFTveJu4C4wnXFFxZLcBRPbU7nTwpfvSCK/Rc0OfxwPwVzDi
8tjHnSnBSAgJQdkxyKascR4iN8PuUfcBvQs8dtjrMovVmSgcNq2PqQ8ENKrA/7NF
DMctE85txp+M1K14HUUAsEIMl4lKJ7jhi7LVlpvUH0nlIRU/D4/Waz0FFuLJ1e6i
ytTInDZri7W7AQSIcqTd98C/lR0EL/brRmGZEMx3/4mlnGwpovypM2J0kixKcPx8
+m2aj1smgWyYDYIq83Sm9HAnZKJ22Vsv2T+3xdgS3ShgDGEZfuVyWJJe0c2gikUG
7pFeRny9+zw0uz68yM2wuS+JvDjVMsdKG6Z1dyYN4k5NRaUskCdJ+Dvvv7WRjtFE
1K0f7SJhJR53ymj4bHl6NFKFwUajXncHRs4goOPW4ASNV6+yNc6iHFz8SWCOvSOY
8F/GZKSn4OgjlMOcsNUAdkLxl4gaSL62P8EQrWS4Afk/3hivShHrFBz4KJFaZGvC
LK3H1dhaG0t9HhBPBci1xnvCltpbJztE7IVKRkgENZzI+2XzICYqY9Qtd2ZAi+n5
I3awQytk732JTx2Wqo3nEcqwP1zywzyTKfoCAu+TWlMOtA+/wJOduaCc740onX2I
Dpeu3pRBMmEmZL3ufvmfMeBWHrhIV0Co+oPleOjIaeD3SxT79EcmitNrqH8e71Io
P8269PQcWhOu6WcBEFaNOC8tTpI6L2YeR1+vSpaKOQv8HFY4bt0CXUEJAks6HyfF
j7MBFSEBKLCZemD/WvMGxk8pyTjHCWTRIiFz4IQRJF2+XmWj27idB3OEsc0v/vd4
BFt2b6EJpzdZ4ELWMpRUe7ga9F4thm9r2iOLSXimREogtoNy2DNkD/f/oZTTQJoi
Sg7crbDt2mcwq/OZi799+At5Np0YhsaQ4DH0T/rEixCByrexF7rXJS1QPAfqsuvf
oc9NBXnf5Btf08SIwmrgdS0pBsgtsqkhex/i1hw8FBL2xDKKpoaJaBD7RtY/FtXM
rJtKqQjUiL5238Zbgn/G8y6bpVP9+us5BXFBxtwXveGOCWKGJrp+MxO5GKK2Qb43
mZrNFYXSesrJPgQTYRTmhKLUH5a/on0ZkbulBer5ATpNSKp+jZ9xEbmQLaezvRAE
52WgaF0yar6LirqkbstrThbzVou2u2wMkxUtQA+NijfW+mRDX7HkT8bgOkNrosR2
mOTyZ8rVCBNxAN6FlrJezONN492zIgDpdTkCB0adisIE5xzWT8Ggf76ZD8AVzqdy
3KZFRkUSepzGA/Sf/8a+wfEUT6GHD//FcHCPsP0Y+4Satvp5Njp2qMVAceqkC5Wq
ryGoSAKPjKUYtMYY3SaCkmYL8dJjBqBeJmrSj1ejvMawYaezEhEimmH+58qQcDwz
KMIRp9HL89xGDKK6p0rWtGm3stcOvVP7BGWzqA6h8fJsRdtBe/wqW5DEYQOsCMF1
ucvGZFdOMo7jOOodSrbmu1u4bqt1xBE15gu6S0IYxPtN2XXzMkl6EWVAfVc/oZ+6
b+3XVeIkGaOss057JKO8QnLmY5QK6WdCujzXROfsG1BwKuRvDqRvK/gXktWCA4HH
LCVQlouqmx/eadikyVTyjrzsgfdTLSzCmr8Xf9Yn/Rx/Z1OiJxzDGuYeZyRc7UDL
8nTXBSctLjjfgeGqnm0IRMr9sjty1gIH/DktI337TK+9rQhGILXxIj0Ls9S5HzXR
+ijXSyPFUUKeYfenP277+Z5rZlHjTNsSFVU+ipq8Tv32IPW6J7P6mSftk0gW/JVR
XAJIgA6c+ynSaupRbGmxbYdfmLJ/hPj/ijosw8T6Nv4r01NzVKhGfNgLgssYUteu
rHRUHDUdZcjBhaXLQx8nX7TIctuArOSCPyx/iKkT305VH7LxhlegnsKMcCanKk6S
q0lmXl/PJiaIN5UbXocRkdTRTlLnUF8oQIgWsx1dEFu5gAuRdBU4+sw7s4gRWLVx
yDsO2/pytl1NVKBIMEKKJgSdoM5HV7s6+PcxI4SdGAYJa8WC8ri/lVTHDd/6oKbP
N4mRHJBA4wLzdq8LAEJsXvEhsWDteZz6k7Jl0jZYHflSkLlpL45OIVK7bD1tOE/J
ezmn5bVsOM0yPZkoNBmoN+hFc+Uqs5rsArL1wGSGxHbqQujuF4kqxDW1SKx3GKro
RxPy94nyD4A3xE2kLSvY7LcB6uOXvg1r1ySh2I40SZegkQATplhYfyJfoXo8vpdk
KltuIbdTTQMSOLZolq6NM3ja2KXHMM71tz+6fE5sghJeMLRdS90GCO9JB8JSvKWB
4wHkLkgWdbHWEztvwWdXnia+Zce9tGZo98c4nXqQHtpEMsQ8/nbYWUiM+nuzBxPV
QyikJlOs3CL1A41Vaz6R5NKFpjYrEpwAVICE6MDJfcSWZnWkCxGuTEj65kaUXYwb
fJY+Gz6X6SCnLSYdPnLptVrzZc8nGQHL4gxhm8rrJSeCskDLRxce84RtZT21lOO3
t43S0tmXbCkzg+AOzvcAZCc8Ubj8X21cwwkVEByFSICZ+/za+jAeQ9CUvGQ9KRTV
yMMrpw9hsqIZPHVCSGx8/NslFygzaENkq3nWIdeaUzrwd8sqoUFfmgt4M5PiovOz
1Rq4ooGAn1XyRQc9+L5NgavvRd5YXekOEOddQhgq3X33jsd1ajWABXw/2du41DtN
j0jESflNU2ZUj67gByd9RGcSDxKC/AXsrHaB1z7QaxgADkGofU6MoTOKpDT45oxr
u6AsjY9NaWevK2GKl140HoTX4l4ZTawiw6lEVhfMw3IYqIC738Uiwj5bAuPXAmTs
+5rmSC4Iewu0XpJNr+w+nlp0pE8hCY9yJaewNmEB48sNKjroim+xQT1r6nJ7Zp2J
gAVKtmGbrFLqSpfaVFhRK6h/644/31ty8odwxxWkKLklcoH2hhRrIH/pVu1gY6CE
zbksAF/BF6UyuYgzHiwuCNS67f2JFptBMyOaa8itp35pxh+gug6MGVtfG1h/WzT3
oFNpQRHrlgGt//7p6W/kqnhAvoJb8AgWYrJOTNIE4DsLQ3/Gd0e26INTGazv3oQl
8KLPmVXFUo1ELO1epjNedhJAdrz8T9Cnt/yteddifgoLETAI86lmIkLSmv/0hssw
6V5JN0e3kzVwntr+wheCU+B/E3d4D/cjss/i2zmy2sqZVLkahvpXTtBAQ0zillxW
8w7DgFozegH91ozNT+D+A9nGltbecSgN/76RNmhjpb7lF23ZvprmPQNELDJYOVbt
1z4lXGhP55QAMmlZbBGTVy7IiqS1tTuNhiDCvokOS2fhDAv5+QfN5J4G3cijhYGP
cKB8NRDHLAy4l/RubJAkOQTboJgwGPMw5SXatoLYbqMv0gvILSJsbCPDao8J1sx/
vWT812OiRKJC/+Iy73RBn3j4rFLlHrhy25Myg39z3TN2Q0A/x0a+KA2ZPmerMhyE
vZ2oSovNzF/OJkNtNpPgrshSfDpccEf0jcUhJuHinxCy6EBoWjPA5Vcri9+mAcYL
ZDbK6ngYHq+iMAJmYS7DDRpgRFDdsxlsjDiAOB+U7Us84dkhiK5XilPEZNz6AVcs
YwoxKT6HdNBy7jDCx8hj1ZTZW7ilDRCN+mGjLFBj3RZKgADgcIYNyV4GiN4uvQ4g
Tgg9aEch3RqXwXWHVIsp8HZe7oR/smI19KGlLvE3iKQixnVRhNtaA/shmuUXVOvi
RCZ+cvzHQPTBuFhLQ26utxtxjUqyS8H0vriCFRGhSOSgczgocCN5RX5ycj6V21ah
mBb5fLVcZdwP/vatgtib2lRyUoS9ajtapvQI04TFa2z3PdV/5khanAR6Sxj93+2i
dLSss7rjcHSWalCbcWUMmOMj1FnMuUtdFwSJXQmMT8RvTN2F+vkl1TZiIpiz6vtG
aF9E/iljuC9kk/S9pc34udimhLZ3YKL3pvi2Uw44N95B/p2CTPCLaWNOTQdhJQkV
LhkGkMvVQBRA6wzgBxI8OFhKJ5pZvODrANUz07f9d5Cnt6psK61/Tb0eo18RUdOP
3D6lQ8WeG0Wf0FBRfOuLdaNzQS36Z9TKmwCexw+BjGhtGeXQGovqMBk1s4ymUgcU
BD8DvKtrjbdJci4Tce2LtkS8KJBAmJrwzQjX1PQuLO/7qwG92Sf9uavK9LRi0HZ6
JT8uPbkTzLweqDDWs1U2vSzU3ksbpQz30UmOwsIWj4vqw7SLVymWp/KSkqG78HBj
MPuQR9cbR+J36VoQZ49UPfg0EWJMFSSrU4vRubmyXnLSTiOW95NnQKM5zcL1jm1W
SWU/zzuAebFmRZU/1spu/R2R8nB2q2BBxrwHtYIbRqnwNgU6yPoa7lOsAUvB2rM/
cE+4z8SMlcCqGLUrxk+d9pbWIX7AQX63Bct231fuqTHefhvTBPbDA4ys8+7TgDBe
WP3s68hjhEcAJBM94Z9aco7LQG3z9x0Hy2lsUWynzRM/u1lyGPJB/VuY93LcCjoF
bWcLTja9RQ9zvNlyJnp+ZORWMBDauVoaAvWAM9dlJZV5SFC6Vz9oyEII1+7hdrR/
T3faoIbPdLtw5yoS5o7YV8jW/SyEONRtnrdOKNasBH4kIwoz5dCKWzLrYm+riLF1
W4yKZQDd7mxibgtfzL0gKxy4lpHXBdfP+xyBPN+/43mwkbxEurBVgomkhAR3aYil
XL7FS8E7H96tqUInzzSNAbdtW6Gjg6KZD0T98sDW4HEAn9PyRXz0XyFaXnDHVZus
oVR/p83/C6w1wh/0E6NZkxhXr1VlopCt2422A+K5FJjdQ5WbMBIwjb8P28wsQ4k1
+aoA0+8UuBpWZ0DQHFjyzYp1+cvNL49nUW9CBPC7Su96K4mJ/adHqEwyIzr3kEOS
AMJC65ugRx7rjjhDk81r4Wl7ehJFhQhBCrqAAzLRrETbzzqqjPjVXlzMK4H4Pfd6
8t2MT0RL/ldVY7FAkWjIjeTRwDa56rSb//m/Qys2r7Hmfk6DtIGsyqK6GMjiPWTj
XT8idfMaeEuh8Etv1VpJjYUoluyPfe1bosNL7m/t6iKriQb/qFERAZuwkVlSA2Rw
EwZbIFXRI6eR/RZY8h7voXEMROx8daDQ5Uo9u3wi+bw7xImNpOqawBqqOswrddmv
0zVt2nDDIikeYxSk+F6nV3ZTf5jE7hGNdvhwZGygJMVv9ZafcOrbHGgROYmBtCHF
VsAVfq2ZfeCt/KSaiySElrSlo/RzjyoURjeoBkMjjEbowNrlzdxDOI+2cxVgwhyt
43zy0QcUHgoAN00QydfhsBPrn8M8fOkar5qHDx61nTeI17W+hzEkCxls1vgc6Kdl
M896Qon/2kFKHuZjlCa/A/JdgDPDg4iSqTrreiEOO3899yfSwOkP3myH9omNA1FZ
/t7v0ZOebacFnI9/Lhq8gy3tV0aICbamCBkCbv8D+uvWWDlWVnguc0YJeiW5+0jh
gSlC1/fzpI5de6F1sKouxKbv78p1ay/tVdqpnOD/dwFyVcLHrZY6OOMWpFxchKnS
Y0hNoyyvKWqbKEn54pp75lTdJ3NzdQu7UYj0a2Q8lAR3CYfyeCmPN7oW9x9wqvcb
CrRbYzjp3OJrJME/w53Wsi8YCjXYqgfd3wmyWcYlYBDfNpdVaxnMzURC51W6gtL0
X3aYatYXegmOJT4PM1lT5Wmu7LEzscXhtfODdjgX40ir6Phx+m0C4FUutRRbRcR2
ccq5aMxY5c5kDa4Cf9b8DC7awc7x7peHlMfhqfS2M15cD7Q3GdzZz4Em7o/zt8OB
KWM4dwVJm5QWijQFAMa30g==
`protect END_PROTECTED
