`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
i903aHsZRaRHTU8t5qn0PfbIvksF708dDPmQJ0hINXC/viVnsjEzTMdt3IO2toy8
AEVdSJotTd4m6dABEWfBWwQk1u6fPNiUvgCtppRy0DaN34bMBJfzOJttkWYG22wH
HdxxwQYGpS8jCqFyhyvYVlEDQ+C00x8HjXf6GJK/lORdbW+WorX2WL68sxoRSox0
5UmDdkDnwrQRrq9FmcrdDZsZWgn87+Y7sPWNUNTCTx/gkMKW8f9+cZIRXEmbvSIL
yOuWFtDZD/URNR2z8ws6um7jY8+KUh+DsDXWVy/YRdiEOtaq1Yl43stD0OUWk+8L
`protect END_PROTECTED
