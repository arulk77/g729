`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBxEzpgkW0a5GttU8M9Xzf1mtzfVwdpdzW4FQvQg1shj
LJv0TvvnwKR0bBWF6TNyh8uNENXtD4dM2Dd86odyX+lp406oz8lndFO+RnnD55RL
sdhCLfsp9zMk3j7Twx/9NAXhDWmwjPRzfWBEtLqMpFKeukv3B7SzREyK1PPmWY5a
264Q18u9sX5cgFesgrdUXSA6+3w2ggub0WEjqffn4vbUbHRxFOUNlleFE2t/f8Qm
9H1FxMTtQBnnhqe0pkh8KbGh800z6VRzrmOG4gt/Kr8H5FpqU+DSajK9zqZMjJFD
+OwBE3rKle2NvSkoqzlnyekJXjvlr5wE09NUEjHCpKvEg91q9yFVaHPs3558ZwTu
RnaJKTtWbrK2cvbt+jJ3MctQ/TdycarEEtKEYjGYX7rZLfkbL0ERJI/w1B5KgruP
cy216Gu6RVJZUdxhTJCY+bTxbPuoEXrRut2jXYDTq+jHYs/+/3guVJHq1ITVEozi
xNUhLYzQhqn8CJBb+qKez27kpT7qFrINuJa2VD2hNnEzVAH5L4w6tCGotVUsSzu+
`protect END_PROTECTED
