`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
jGG1MI4iGPIxy+Iuaq3B+fLSB1oOUBoLw0FPYtwa53MOmuI94wpldu9EblOGLfID
w+OcGkFw8sFDcNHKZqAVIs0ty+zyvi9Z+sBAoYDaBbDfHBSG36ieMugDwrLqkno2
4c3MuYmsZpzQHjmHuxb8sWgDZr1VpvT/Ri6VpvWAXkdHMnoeizguE3TwILCWMPzx
iILO+UTgb/g4C3+eqkSsd2wVW/W1xIP5qxmAXEBJczNn4LHVzpyZnIurDjCoqie4
WJH7RpHCcVduZCZohs/vL7j+ljmoCBPoWDBADPkUPN62t/gXX2ZwV25p5ud5Ok/Y
4uo1X3lJPeDdOX6D8/OIu1/sCkkx+rteDOBnniMvRfszdg4GPVrYecZ/SkFiwYM2
mFZjd9RTWBUFHgyVGyxxvPbI2P7l/hK1F81O5Nan0L8=
`protect END_PROTECTED
