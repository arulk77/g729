`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGRXQsmt0DWqRs8eaczAo2JFmA8XgQJiZE7hXFvhhjHw
nCvJSclWSn4E/j7XFiGYO2HFzAQzmV7tJCbNLJDrh34QP1wnfSL8HK/03mNgQEXY
g+7SwO6Zs6foko2Q+7bG+NqUSS6+qe3d16n4+Zu6nzOZyit/5CTixVhCYmEO5C0l
XMesrY4eClYlpcyU3QTKmuuIAdYKnrRsnZcLJuBgw3/FMscD3USh00/+kqSBgzBK
iywyqAf9nRlhc5qD0IVBhRIzgHu2FLiG4ILhtlQnAFIvF6pz1ndqo9WtaeKoYqbU
HxdVDJnMUckOun4TC0uN5pnZrDmaNnd9mxeP2WF7sRQ+9Q+UuXaFytUpd8XuTgaE
JykJuqyqtbV3dPM/WYeBJBqbAducGUGD9qB9eUJeXlQSaYwy1udj9enrH7oaIJI/
+rk60qrbaEliK9So/XpSK3hEvH3zp3l6n/Bl8otjoqyaNSQ3+Gn44i5Wdha3vuqW
IAZtqv3xVZOy9O2wcjPsCNEEC4ucJhsXRET6a7JLezc6N7cH42qa5yF6/Qe6Thjq
3GuECTYXpYOmx8sdYWkkmubCulPndkUPOorYzhfkXJvnEwqWGDgrG24DqBaSEsKH
`protect END_PROTECTED
