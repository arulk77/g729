`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkaWtwrANqZDci0AwTD05GmbGFXAyhjwX0Lomg04Wo0M6
QPrJwSAvsXSoRH+ISOnR51TDaAMC7GbbII6tR1ryxIBB3nuZDq59fCbzSYHW4GAQ
HiUU1iar4SCARw+xtbZqQ9eAZknJQDKDsKOgsluQFJ6wo3kEgfhUA9aGhkBF2lWB
C6B4tMm+4PIXxzqt3ru/Zf5mxXoZqgyvJEfJZ1/DNQC8vXKQ9MiLM8dd+bFOZ50H
s7d3mzIaUGUDEVxeZWaXyuXygfkLGTr8rtZbYMBnbFwe5z9xOQsF349274lS2OVG
h5GBYt2xRo7ImJgq2H3eYZn6eWQC3dN18rAqo6BVBOH1JVvFJBzYaRExzGKzB4Iy
G2aKlgc9EzYBF7SZmOW5jRpg26+abQPorWfp3GZ05jM=
`protect END_PROTECTED
