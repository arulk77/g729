`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNScnS93ynJYZYvTjRwGqvnD1BbhlW23sDiVHAMcwIL6
nTy3hCfHv1FwX04yBVLbOuUYWhLzU2O2Q4nfxuYlidCKsICOP1IZwxsxwh9615PY
8vPXBLk8qDxnnwHqWEqVsEIypnpmxDYubYbnpe+marC4utAdM6WgH6FZgEyV3vtc
8Mv5R+8VuHZv2UHtopm34aAtGAnKnUpfJ2koTY1HWTYVQZpASqZyHmGKDcmSx9sy
`protect END_PROTECTED
