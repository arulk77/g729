`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45IF+yZF2s/c7QYrdGCB9S/ufoGdwCP0LVP4MM9DkKMW
Cjt1Q4slHnfk7WQh/8qX969WXwa3b7AdQDPd+R2bEH5NRtgDtRFuvht24OBrqacB
djMx4Q97uKlvLm8o//9CTwwGlu+igb69M8v2me6C9nBHPCHfNqF4qC8DtzNNQ/o/
LD8MDtn5D8Tl2MLR9OgBXYsyjYa13LnH2stZsvOlJiOa6JOZt3bT6R9HlH0w/gE2
M37YTlUJlm+j4ie60kliOTbBezzsCDmE9glB+BTDFn4=
`protect END_PROTECTED
