`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkZoRczKnZPo6PCSIaqp3eRrTRq2MrwC0pAFLTz7hOZK2
f0ystQ+L/mNrm35IZYBFL3pQ/1JnIy2zLNlfzVYGRCWEmMEqhWMRj5Ofpulvcejh
Y3S7FnevflVZd0WsNcJCqfzzTcQEr02pVsQizvWAQC1qPgU8+n2HOJIC42xL1KPR
jHQzhSqCLCV/i97WMW7XaN1Rif3SHXQrNSMK6rykhHHmkUQ7jfeSMqVY1jxLQnZo
SUQhwnfFjAMfhXliChki7ZcrNl8hGcXOiNLkrA+z2N2KP7rKFBLCL2aoPk1LEHEY
R+2V4uJoO60fynW72blQ0C4XA7K3NPyTZqgnZ5lBste/SnE8qid8hVTuVhaEaGY5
atVV751etnwBD7XRbe9VXi/Ob4lTW2v5zuyibhvhFYQQ7AUTkfmt3mfN974Ygzja
NR0w+XuBfKpWcrQwycPXEHNRTPaQqMhjNUa/PVSz2D86a4XwXbMu2tjStEdXhNbI
cPZrmQE5oVDgdMLP9Fhx1dFWEmZGAb/QAAoAYuIIJQKnB8mXDdxhwCVMzjaGYlU0
zQXNaJ07EwL9WUXPv8wzNJPY2WzwdeuzzAkbrGnsSEOCTLU8Iehl7EedlXFIy6Lt
JmSXjn0DJd+S8i7RXXuNa50CQIh9XbYAippfIv2JhmxKBxw9OP6742YqZaw6vmre
PIUhHQ6oGJ2Tnw4gpDq3svQmd6qKLEiKUfZqgLLyeSA9EH8l8hBbbqomy7oMSebX
fS0ocM26RaPgAuuSGYTce4O7/1GzsqVgwvn54MaAMRBG7tmMfDDjjQFyloRMzqux
qDG4txVggPYpnMj/cBOeQOT/8jBjVNBClO7huTjCECIkPV/1CLo42qvfy49AHFAK
qVryAl0v1rPlIhy9iQUiLMigDx86iY8gyGkEZqzwjq1jZl4L36IQbqIXjbGQvb/r
GQ9ltJG9GVSIaPZo+lEvFH1tcb3ysGcF9XxkmiR0woe+s89nWxvCZBUGbRq2oaKd
INuu6h89G06JpOTWw44KkGnyb1f6ZLG/1WXBYvKXKD0nV5J+z9HkGeJgQMbmaSA5
`protect END_PROTECTED
