`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFuLSDTvLPIHgnDofh17t96R95OrWLeIUmX1rgyJd3Id
YPkUbWPgo7/1ZO6erAhcu+ay0BUVPLFU7fRxeLoSpwCrrdG7NJUhGcAyY2SwqKPo
/52XdLhsGH/4n10LHukUhiw4DggoE1DaLH57eDdMovGOMxSfsQNpU+O8ofxm8sEd
`protect END_PROTECTED
