`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
z0yHr7f55zN7WiEPul5Xbv6IJ1og7T7SZyxPIg8EmRnsJchpbOsnZlYedJqeWaLf
IYfrdHdNNIngmQQ1gDYhorC2WMXXFyVkp+FQgsPZluIvUyld03/nCBlxatPKMsDq
V/NWenBVRlQ7MvjmlQTGyQyY7qbTSJdmRK/DHE3WnPgukIsR0j0csf9HFmnPk/ix
9o98pOaI1EojvmbQRMcGZR/GFdakMSDX9ALK5BJYHqWKV9VJjyXGJWXOII5DwYAz
X8TH83Uyd7uhVskhldby2K6ibZtRdc6mYcTpZa1aoLVXldUL31Rejz/4pCSlnGwK
hsnrdez4BuAYMrOmKOiSVhbDyiqUSBmkx/uNlr3hqns=
`protect END_PROTECTED
