`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SaoMoxXq7hufwQeeLa03/jZfdSOkzNjHe0iZIY8fYhwW
xaSMlrkkFzZcU5SCHOHPMSlEYeHrBCYpnFoz+qEhZMz/iL4L31iNpbZY4vXO+FaM
rO07Ey2UxnKtwwjWSrtFdyJ3S1W4I6NgkEnp/RJEmUOkVI2/n8Ro1yUwgM5HO6AA
i7yAVU9e246hI06EBDEEzNpBhjoWVhHPr8eUIsRj6u+7L4cnN+B8KtL8FCSiwa1F
fK8zePvT0LEeI7D71KzHjCFmgJ1LH5JKfxPOVuHlQUTHSw/UlMHZkYUt8v5aImNr
DA9jMQnoip03Q/EARRyuP4pV/zmL0FfnJHU/spgAMEzCUDipH1W9eJKrnw17BJQZ
vV3f1d3LMI2iPK54tmUrcwXJxhquPXUNUOYDwYVAtif2jxuC9swwADZkxSmL6RKR
kvZCwphwjxllif2K3d0gY2cOK0/TvAuL1J9T4zpgEgHSuZZLhChgdF9KZOAHTzXA
k8A1IqiJpaBqnQ+uzpua7ioc4MfzNLS6+FypiNpWwtV6/3bI3xelmu+/o1K0Z9ym
coFuzQ13b5uZUr3HGh53SQam67gs/IymO5syOdhawqSrJsgwMHW6y+ocaimuPQBd
cb6RJ1EEVVFFOcpR2+7VnuF5Coa8ToQ1RoSd15TSEFKNpJTz/KFQhp2PxW7S6iPN
hQzFD8M3Bs1qRETBFM1+k+wXnHpY6JoUQiSqr9QiCIAaSuHh3urIv7AVoaGRK4lO
Rd2Lf+OCeaBXGMrpgt2zMuFTXh+sAhXJjmBJapvO1HJkdiMrWDJEuKXZbgWERcDh
hKPT7tVPqikCwThibPDslIsmWXmxWSxAKsQbyG9GM+kMPYusZJlT/P8RUSpK0e1s
vI5ri8adMUir2/iCqJdRqvhQQ3IFoWIWDB5Ai/TdFTgbGByHmnPLpSoQmd90HW4c
0tIxuW1dATRqnWP6MQPj3rzUT7+tqdLsQrXpx3ax9/SLxyWZDDYJ3jTnFO0UlJkr
UKv+QIQfHVVxJI2kegLwkfS7f0h52mdfQsHbbeHxN8JBzPBlqIQzDXR2i19zYNDF
exp/0LEGZu/T2bEmRFrfJfMqf3HmdPuEUEGIDz+7BQITj6JHa/JK+LEO6l/wxIzp
oGzoO0PnICOXJHOMC252H9vq3bJvxA4Fti9gM5xL4eJVPOdCTQtVV3JvJTNP9IBC
GnJ10ou3/ajp9EIhqtnhPVkLAiLCuvzVLcbLQ00vapIvNRWVaOOMY/9VfvnCeE5l
MXS1jJhn1PWnn9Rb5q68IS3tpgy8a1fzZmCXZ8stnpdic3HGSSJBvGKo0r6xtqW4
nY8NHRJymuFpOXHJvlrngaKwfvapyduhkT/eldiRBvSUhMPkQ6n3NTTQjNUUj8Kn
DAaCMB/yjwajyzyuGYMniNHfQz1yDaYT/giVavODYXbLEyA+TAgrvBwJcyI0Ry/H
uVPBrM+hu7hy3VHZKOsUlaQA8CvKBMOOfu4Ae6S7yDvR0GtfC0EV92ertX7o0mZ7
/nVd0ONW1Py6VPESnizMf6EC5QX4ohm/bnZ4EO18s+MO+Sb8XLmwERp70pJTd78N
Ra5ZBjyvpu5iuWwn8jVKiRNb60mUyxipbxqNA/uUltcNMavqLXbHNGg6itp2vFBG
O3uwF9WZQX9i34X04nzztzny0OB0oVzjX6gCYtkG1riKAVh9XCZCAzA5VEhD1VbB
jcbKBYpbE186H6qrI1bghdqsG5TL2GPObhuNboN1yF7gneKRc0bEACVWoidU/+Xa
Tjv/wiavmKdFWXTBuWlQsBpW03RUaZGuKuov2NHReyrYjSOuUtXTdyXwNkwuNmC0
qVqovt0h6d3SPAEk+c6T0QvTxR4v6xryLPO+VhVOGm1d5NgPg1Fe94xobq7KcaNv
8AuQbCeKS/ilL8o0C3cUjQw0M14RO0jhu0230XzDGLzEpqv47qjOc8jH85qE5X1w
ay3uRaipOplTvKs/r6sVqQ0/hiMdw8w0dvDhBMKS3bGgUjT4bsDaQ8EfGDmk41h0
M/5o5l36sfUbKU0Zve6xCNUuGae3P2EPzxMBQYcsPuxRw+XQ7Xym2B/QGrOG++Dg
KiGqz/dfbh3MitQDlLC8ogpU5hLl4qzn7KoBpEN8rpvq2QvvINWUySXa7n37ErZz
TxBoDT7T5+Pwipzr+KQzTFrSZFMQokXMCOvhGIxO8w6Ra7wzPyWzm7CEbuux7jKR
3kZaDn/JtXPy+ElPg1qZKu204fX7q/M0lgd46fDWeL0pG0aGuFh+lPBjhs+tWrEa
VxfB4mZSbhfpRsZSHvL+RcOt3629lxhrosMWetzKsBGU3IiX8MsVxAqdp3pthOAd
Eo3wqU5PdIKg5g4I+q1DSjjCT3wFDTbjf7VTTEwai7W8M194f69HxFQJtk/nQ1ps
e007RKBMW4bLppPaE22/dnAeezzmeWSW4A4z57A7y3VbzQXKA5ZlhLqTDjutDABE
BCbotVtTY0BmPnOPVOhlJUfqosGCwEZngQF13ArbNxoUqpYu02FryDDO6mFs6Ejl
HtNs5E7FJbGcd8WthBHQO1PDfIAff4snURhzAMYl785+CraK/zvX0IlW+OnEhSKb
K2t+V/Bar2cROdFTy558cpQ2TwnqJSUalnVOjNXnoVlEzjOpEr7DNlf1a82T7BJP
Rf9b6xUZSRJnKVcNRhsQijLlFTzQozJ+Vj20g7xuL7GDZXI5MGmFRswhhDk/f+10
PNP/cQG68meXwiq1n2DT0TtEXzWLBaWGs4PUl0IeQA5LCVlDLn/hr7CEidB+t4OV
+A9kOgslPxc3RlcSOnD/xNevvhRvI1qSoAqjaOYVeOkfh6oanet66Ca0Rfh8Wj8J
g+S5Y27Hi9N0vpX+wB9aM1vUg3BKBM1Wh4TRp4xHlGKaksV5pRKEmWV0EwnZy6mq
tQ7uk1nNk5esJ1sv3Y1be1eVy0eJpFUenAI2iCcx/lDYP/YyVvdGuZ1IVSTxdW4J
pI3E5GR4Pvjp8M+6rZcxdoOTty+SDj9atlXczi5F8PRnMyV8+FyrhWnuMfMnLUdA
OM1lLx1IvjDIBddjKzocTwgarJnMsBsHIlEDuM/71CggVMYCiXq3ne0LAKpJuxee
/bqpyG3fjx+UWwgyp149lca/fpANXPZfI/zNbvOST8JNkffVchnFlDwCCPg8VN6i
KDtOX4yJPg8axu+w8G7577XlJUisDrJefyifa2MJzx8b4AIF3ZKZrzNX8Lnv2LvG
yYYoKTBC9Fdte2+zeNHFaMkRDxBSFSjMrQjiNGj/7cHDTMXx1J1P0VItz1iBw/VK
4H5acjJnFj/HN3Gv0mpJD/Rfi2BIhmWU6aqi6wlBZv86D0/tNw6lcZDqgubrejnR
U2QzH4jbdDdpZKWsmjOjsMBcC3yamMOpvxfSYIxLlfX52qfAy7U5hjqnomQRU/gr
gdWhFu25MtQ/5zbplsqo5Lr7yy6CWyNGYMLs/zJXYGcmdKZABlyk6pDvpqMc1z0f
cKEMnQ9L8qDVxqLQh/ah5z7hQXEDSbrqcs+ftbBXYPaMPGRB3bk2Op88coK2qPkU
ZTJu5YdmnAQYgSMG3fHqayehnQOB8SE3u+xUCZkH2+Sds4I/FiJ8k8YHEiGuQ+rK
ORio1b5jiK4HxhjXEcuetofvdlLk1Is3Yw4gSaN6ID6vGGLVY43J11T/SUImMoQN
u5QrR8luexblGbBJaAeKuLo7K+/upY+BPo1RWTnixiS0FHm59bsSTE17UjDf2JSp
kYfZX3Ckpm8xCUQWkI8eBSf5Gm16ZKDxm+5qHlHoKFs5jg0IKH2C7TJgzSKhZCwG
BsZWC1o4V68z//RD0GhE8Dw987OVfYQIb150dT32SGFWDqJwlPKTTe4rK+7sWPF6
RXp2B07qn6EhybWyCnzAcHTYimyzyMofNIjjO4ykKZqLdc/gXVGoDwZhowTs4iA0
nYtL2ExEMmEjr1fyNMcXGHVycJBbDc0WrDxWts+nh4Opo2/hf5e0iQvEFEOcrnMw
g7EWevaLKhc6MiwndOTqvN5H7gR82ejr8GUbbYcGY98e5lqbR3eBpiP0BYQe7+Xh
fis3qOSnK+eWYxaC6MxWmB83cncE4l+RwOYzg6l9vVk3PD0Sdt4Z6Z1hP5xNdOWe
f7rZC7IuRLReFL/nO2GDbcIvRfSQFYvWdZN1JUubObgTxmMImwjk3CplMLHTD0/g
o/Q2gihgptCTVBm5Hcw72pyGEOvyjs7tj3en4v0zo5kAHMC4SB4Am1gm5x3DnfXR
Ag6DbdjZeodWPfsYNrGOeV8Mh8pQGStZU+COktdVCujij6I/d7E1mDmm82CoCbX+
`protect END_PROTECTED
