`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
iL+62uIoAi+VhMzu+LXKQhgd8J4wRkFJ2tu6/Kw3mTJVxVyMiUQ7Mfa1rggPQ/U+
N04HtlVzMORx8iQaIJOrGQZNL6HrasQbGKnGNyzII0qzIfvwAt+9b4z2EVbVtJbs
NVbK+lWb5m54p58E/srfGzx3cFi6VirYoGlbQytLr2gnWWHtbwZdMYWPXJusqHDA
VzmhVT7EZ15j6J/V25AdQcmWK1VO6FiLy4oNaDZYlwTxSqJyC5TUVwWBFJv1YQWo
XAm/vY0RbJ+QSAJJf4Y841p9npWka1+/lMDGkdsr0Dh7AkW7mfdoM9KYeSwB2me0
`protect END_PROTECTED
