`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG6mCEMVnzl6K9zNt2SiC0CJSVgHYZijPosNPSEmJ2o6
WYXBFdyo6rwPweV8pgU33hj2LcP+qfL0YrHmfWae0JVrp6YV2RkhwnDlsS723Q5q
MFdsgJ8WuFj7Si2X3x4Oybn9eXF1kIrVwSmLnznOHe/Ya3uDAk7XWvtD4JEm51iu
HzP6XiCfV1B0y1CUrZObH6sVyzqHfLqAisgfs/3LG+cmL9BW/8Uuw4+a0CRbdt/Q
Gftbx4hauvU8eVx4tj4js9TcggYQ6vpUGeeKgPKfzg1255EL7IkNc1BHkayS5V+v
E5O00UFeVJFZsPYXPs1E/PDFs6GSOhkcjsoTOkTYO+vzPxcvyoVfXrsoW1UBuqPf
e1xDE1IwslbUXtBZgWr+ainWfrKGE4+34cB9rKhC0NuWOV4Vqp+WvyOXiPwo1++Y
QcldwE8w596o+sc/l8Uy5cTOr/tZETP3a5FLgHXWVcbJ8luep82G7n0Euf7tuB/m
4XY/YdvITXY01m3knc11zVrCwAg1eL3eaBYdtcXN1vCA0wpcaisv49atjL2piJmf
/k4tA8clWhgh0MIueB1Mgg+d5b4MLdAhgRRD5QFpn82ieO7Jy/dGJlcCIk0KJIUs
msUvSP2DqmP4TJxsNerjL+b01Do9gOuQg2RgW1NsNOlrqu8pqVOyAzKh4FkPIo12
DdPMQ/hSsqDeq5AJKsrF8ul2O87JQ8QSb5PSgteH5kKoYfn6QMyxsmxd1/qqJ67m
SMKDV6usA5AX/6r8WMqYbTR9ZsSTv646kySasL37EN+S/QhfvSfJoRYieZw33Twj
pnTqjdvsqRlVBVSly++DJ52EJigF8H9Mi7QZGxFtMgc=
`protect END_PROTECTED
