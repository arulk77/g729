`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42EDZ8Uw5yh29/rqL1FZVy6YWQcoHUuQ/ACdAVQFu9WC
VtxRXOWPwlLmdxokb8zmNOXEzXeyxDfd+cEjXmFC1e6XnCWAkwEzJei8SkNI0n4Z
6aAPo7hiPGCJx2GeCMj7QugPzhnlHYHapwLEsCgxFT7oGkniAKW2FKEgDIjftoWs
WwD1eRODXngpgDn30zozjTt/10Swwe+za5MBd4/X82I=
`protect END_PROTECTED
