`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QNw40IqJrFvY2E8HYWz+jxThIGC+WpFddy+MDr1dmIm8qxKbZp+13B68JFeQAc/C
SMSR1nlS+82JU1DldJru7ugq+s4Z0xqWfh0sZMV2XrSV4Mjl8h+JA1iU3DgLbDVj
I6PlXkSNoEP9JIkW4czYf/nAZI87q2Glx2VWBoU/Da+TuhBG7AMYvTTZ5D+4VlPk
`protect END_PROTECTED
