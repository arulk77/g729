`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOVw0nU4ymnkngpFwByFrZJtrZev5nS3wtJeK6GyL0Dv
dtVfMuQOJbkoCAA+7RywvLHOrFRal3PXd1rKBTg6vUy7Pnu2zu2N5LqPg3DjMALl
rCBwjGDlvqObBguen75jGbK+YkE/51JEpSttUEWT3mF0A0B043XxQfD7ld5O2AaH
dxDY9ZUahtvtZyc/e7DS9w==
`protect END_PROTECTED
