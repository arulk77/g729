`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
40fKvL0R1YD2YwMc8oS0ciGwHV46Id4LXOUzjvbrDdw/+VbD3NdFSRtHLDPvbu4U
AgYFr952uoVvO4BEDMw07xpeYpZdHU7n49dlqYBcor06+ebomxpwshCEiXor7yrF
edYgmsctOlXbddOt7pkaFu+SyJiCUZDKh8g75XXziYI=
`protect END_PROTECTED
