`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMF3IqOG5+U7HSf4JTj5zE1c2ncLlwSd3eDzoMR8BYxm
P3sqc5gGs6dR23J4bBbACOOSl6pa0OomXnOGk+7JED9G95f9DqO+2tyZrgPxOwXa
yvOL83qeK6x+/TZHBLRJndzQaOx+AyQU53BPBUAzj/A9b/hL9Kn6HoPmFJK/haW5
l4O46ypW2k4ivrUIEX6rccVuAEkcFdMCd9QkuP14UKopPbuYE7RB95prBQ6pQpch
+AIyyd4epiQA2PqDCpkPcKmHgF/HeQzblNPgJ4uWfKctqfozRI7HZ61s10ybA+9m
5guUZuKpJth4rbGu7PKfd8URRC+B2EMGo+GpzuStoNVnujJZhLywS5D3JuKmZpWQ
jNxTU5r+Ahh0xxQANTa/xcJvDW9tr5MjPiQfs9RJ66Z3XQIx8blQ+PKbxeN67a63
gNkre43BjQYGqcxTnjf+PnuEfTXyKI8xQ6NEinUarnCUDgWWpWKNLJ2tFZzBkRGQ
nmZjECeqe9JLmbmGA4Kt6rxuCWJhgLPYiHITnNWiEXfuMer8qjJnEZMUHR+uHSoV
6GPIaPsVSMJMnpUaoaKcfWdmux0TI1kvr4LCN5h7f/9gTccO2hiSWmMpauk5mvmZ
sWR5zzDlKfwR/9RodjmCXiOpA3tzfyOxWM9T3UN442ja/H7FrmcKgQbUE6uJdaII
zGqjd9GqiMmWPeN/dBszv4jxGsWGa5DNaPdbaABdVOpxv+2lk+Ssdw0T5qEFTTtd
tdcRkIBXsTffDOxtTvGZ3i31apXucazHoKhfqmwknqL73D8h0KPbziylTRl1IKFn
640DwseXeHtDNhd+yS3mUmYnqkMhA24HavJsmSEaWl4=
`protect END_PROTECTED
