`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu443osh5pgT79bfEdDDuOUu7xg1U4OiOu1c3Y0uMc6xvH
U1sLs4BBiXZ35xrOI/jeDqLGtlAKOM4p7T3XqUOuxfQtWl2HF4xZkdyX1NxBpvjp
aOJ6LufcQcKgQFejx0AVv9Z810v0eLt3qIHONs55LaNg9w2bapXotzPlqw1HveEV
GU3J5lGfjOUodsJSq1/8C9lyxN7Il/yiNTX2ASWaFFVEEAAAEvBek8M9P63iGUN4
i06fg73KbHnv8nH2uJlfl6mnha3nxBEc1DRjD/k1vcIzJX0nIR4SSuVk7ALqfso6
0AwjlPx8UlE3y3MSFRxMWfIca1IwnBu0xosQKlaFnbx6EJ4Rm8SRzzXVF6nIWaJC
nrSHA7Ju8N5hQ5xmLu+EWv2CZuekahF1ZK9fyAFAshXUrhnTqhKPujnVZV1F2d99
uA8TXZ+P8xRF4h0aTjNhi4suqcmzvu1T9dT4yoaDiti1rHbLXfPhXrHQzG9bb42z
hBbYDdXL0hCip2bwXxJyoi/0z8Ptf887CFJdAie9wrSw6iuBPuJ9dTjFD+OhwEfA
vsG86BWYEbzC5ViCFez/dBPIOV2/7Mfkli0wHrb6dVvsjEgVWWeiiUgw+Rp2D1VS
YkJNm01q3Jhy/Juj6PHCqocT57M5Uv+ItJqiwMN5EVs7T/TLE0On4dmaUyIiszHL
xt8WfnkKRLwL5Ce7I7gXQP5eGPdNgpqo7spf3T/Flp1CnbaybDu7OZyhyE7k10J5
i7PLKDlBM98wtmNhYLyd0ltIHjxILUI0MJmPdB8qAh2+1xSd2JZiXmAQGacAeGlB
d9+gojX0sn5KOCiUqazSv+R3nIdylGjJBmtHJ7ilAApHgZPRy/5weWukFNxjrQGQ
Wd+KYAvqOIrycPxssU8crSTxWdkkG6Jt/NgTFGMYHcvY7pk569AQxfiTnTJhOGep
8mwrXh9Wldl2O1wa1Bn4rkYS5LAX/SHxstdhfternjBrdm38E0zBkKXcOAcSAG63
XL7cX+YkRS1FkqAupC2KgYGVlcEYD0B0I04acd6LAk/XcrNXn+BzFGa4P4lQOUCz
W4uvH1KJSqYDL15hfi4cVPX3UwtHvdAKCxtNGlSPdaO93zzf6wLvRwDJX+fjERRC
DXBsrjl6GLcEKyWSe8708sdkuMxXnsdP1ShIBIrIpqbG1Di5Rk+4iKqH+/prMJzd
mmvjUrR0l+hlUaJTyReDahD6mwBM6oiJ+mVSryXVnKbfSG39NWVX72Ahg3O17qM9
j9Qw4QMGUMo2Xvz5d68Kbea5QDgFcYVcSrIKpnwzTKlMqjMXyWJyqwddLNP1n5GZ
iTGtabDiiRyOw2rQFpuJHF8zHRsPIlRNgOoEMQ56kZAu3GkCi8tYTcV1g3ylxL6m
fKbtJhZXaVc/vBTIboFrQ5BGCs0rJ/HQBzOWiyAg7tUUTj207Mnf2rx+OuvjkxvF
g6xgQbsITtNYLAymCl+EReU7EfbT8eOVPWLSSUaeSmbdxtvVZxG1+N82dqg7ofHj
jbZwe2qbAfI8XVijQNyAaakEmwf1T8FUVLbnpQVV2Rda21UFJnzQo/3j96/5NAfL
NcZqUpGU2JX8Rsla40/o01FRyEV0VIA+g5qc1W7fCnaW2ijpuZ8vndeB/G2vPYxi
JpWQqo7h+Q49ZjV8+WYTze6WLuqavcKsWIiKFe/8+qY2XlOnp1eFyROmy2KIrom7
QY1BBbExhlY9018Wjgjjg/fNg/MksVgvTK8oqOEjNTtZnn/QvfgH0hFbFA5onEbM
okkJyF/o3VlEyUjWljajikBgWYWY70nTwpnnpLTrqVAkdWOk7ETjDOt74fXbxu6D
hEugPGYwfrogWiK/oMlaNPmOopkrjPiRZMbkmX3vVKVjPitQwme8nxQaxkoLOY61
c5cUxJ7QaIO4HS90HqzDM58idn8Ty+wmDLrX0okpkRTaxO9Wmn1qb5R5WDWbrHaJ
SbADPik8rVx+QxcnCjiNAjnLoYpfxr3FfcjwANfkTLGJb7L6ZkusfkCyCeHp0okh
WhVOItjMuLxn0E6n6D4t0oDg5zzkNo4pmcV3PBZDp6CXhUX2sIEbFp0rF6z4nzL8
mjeJEJHC/SQt2P2J8pdURb6g0jHEqQ/J+8GNvlOrLFj3LelAGlCy5azkWf1dZ/Iv
gGzuV8Op7nAfkiN8+DZzqZi2dug8EvImoufmrqf31KPUz2r34bSrTv6B6Sd3SWrj
hH8HOVxSQLt/55H3wK4wndXN58mgUTH+2ybjn//7E7cm6lhn5QHzsLeLDVUM2SOg
MsrTn1h7ASmjGuDDyWY+gRu4NevqnFVgTIqA7aGHVS7rnCVePn9V+iTKlFRhb+RP
ugssKXtoYR2rDiaRIYOMrTqMDjKTXzvNZFThyGbcYkwQ4/ioDu78iuLeOr5hlV2K
QjVqvlZDZnLGVLipG7MNGPC5wgm4SmR6nsqn9D+7tyQ7HjHsTDJlnVZHDiMnFfMe
y61N2rosZtmlZZ6FD3w9iWM4h1PswIFrUllfb881+2/+rknwaCQfAXm5i07rDOQz
CTr6jXdEhDxBNrbIyqI4cXq0eQqkWkfctlLuOHyfVraGfCNuSPmEYVur+AQH5aSz
6fpndOhDhYboxC06nouaGnU2EuchrqP/PR0KZ04ADHaLwBc6WgQK8iF2NonGWBe9
q8fNbDG3nBiuFoCiNkTFZBymMWVQg+9R/775soLT8hf8U39u3OZFMrfRMezBQfpV
799qc+ja1pG6Q+VNMLsuqSLY3Y9yZKX2JA6ow74Lt4f/z1ePj7xa9znZMyUa3NT2
H4qOIj1cPBJy3TU43GnZecaJhSCaUC+7GKlXRotyHZOi7uz7XW8itvYW+uKcsorl
/m2mj42SoQX2ZW39OfE4dsZJ7SKFxvdvk4gLGXf55JJI/O3REaxjVJTKmkD15NCK
z08FCiubNyqK83nKbftafMu9Q1remASmACXBbpQ8ANDuXIkp/JiYPN/sITA4H33t
SabmYHjRxeFjkFx4f/vruZg4nb1IY25Ijb5MhRo6mq862SCid3vbRLOjxtG059Zj
JGwcr2cM47SANrslFT4oewuke3Nix0JCWC1p0NDK6fHRi7M80STBftutzJ8lSJCy
bn7e0FqDALVStiDNr+uefMkOmNi9A1piLkQmXAYZQqZCkNHVrVKkpMbqikMPesx0
7jNk4B9V8Jh4joUFNkZG5wKkFC20h3u7a+YsZ4OLdtw4GdPxOSVvj9bqbIsX1MaQ
HbqBhfYp3aKXNDo6G58uQhqOiy5nQWlZztsPDdc7RrsLMNiXJLMGHO4nqpWX4Kpb
KDee+By75bUXxgUc8WF/Wp11S0H4xWaemcgVHA4UKPR5h74O8P/zir8ldYGyrNjq
CzfwQHQscQkNab7xFy2aEecawQGdkRPqlic2h3AyffOD9Msc5ezWQ9i0EpfDV3LV
ma8+KYaFKNtdMLTIRFJEn0Sat8Ww1QITqD2icf6In20fFrb4alrp/e6JpXq4yKoi
ZjgvbipEaZzjCe1HOHrcWH3xWILEzrRVNDl2e9+YWIVS34ei+n+SkY7NyWgNqsKA
kNkcm8zZn7jJoTIlXe54YKwqRYk7NxHeTcuVAVbbI3WbZGgH9PzAu38f89QCNF+n
bd0ly60LRDTvVfdNsKtEHrukY+Mzy/aKvpTsv/xerw+5KkM0RLxvTl189sN5GpGl
ZyQdlFqD/H20v4S70qUMTE0RTc0C4sCDp4yjS5F7l5cR4NwcsnvkA198aQY+TeD+
ppxApKOK38CKy2KynzvK+M51ZVeQ33XDZlA+BLw02iZ3nn74RwsFhMRXI9zesMDK
vejAVpzftu8mng7VorrMYQ6SdVZFHkeYsc7WGncNENdVYhkEdHGq7dFjzwjrFFKv
yywKzlTRVUgEG1fRHtGbGmxOgNxV5lGNNUQsTUzSYkJk12FoSW1MrF+qqUgkNjyx
1fTSoQGounY9An0NfTzmNsS9uMq6Jx+SYxnov2/eoRpixBgnFonwsPMOObv3UE4M
0cMg2ITsxjvaKDcKLL1OOiJkMfaoH4PH+XM6ZpkNOrpweSUngIqyHfU1Rem+ZvnW
5roBZ3vMro5TsNRqmijacsKBUkUTtNtsJKRuK5CLe97HHFy9R9M4R6FUrQqviZZo
lpzpZSajtG3bqFZvo6OKBH7cun1EHPg3HAZ8jcbVU0SP/gdKKsC872iQSidJUMqn
vekXsL/U1sKUj8tH4ZbYp5iUIEYG6jAIkeDkmoEvjzjODfdDzmVEWMyc23M5GOAP
LtjoUYGKSe6yKzYLzVeeiaIhMJ8LvXAgJVNBJ+V2nR1cobfeKb0SgspqjvfEGBfr
vgpjHjkt86uzijXdWEms/lqj9ud+hLyerZYO/XgbkqOj+LxFltdS4GxJvAf+dUEX
2ilDR1xe3lbULZGP2NahoL/GfOxjVXmXnSmYQWff1lYo+CvBMpkSBhI0qSqZ883J
VnkeeCcLazRyjdwxCfUunEn2pG5tel59wQSmFnSo8CfU3KFJYFIfyzDzCpgK3dHp
pFsg8XJ43g4pVsOJWOU5ok6+SfALD2wjQP+jIBpjdsXEIIJYBpQJGVkxL4WWjs2W
Py0W0K+3P/xSphzMmZ9NqvkptNSATH7rUVWU+vvctyMXuk+beA22KvUzdlZZgWLx
AuSsQs4ot+eEzBXiSZckoShVsPVfzABU6YFCLYNse4XJwczOjrS5nkl/nyPuDuNp
GsVsE0goWLT+PrsYgcPGERPrzt6r14KIwQX8WCD9VuAyO1GPOK3aB0XWze88z8i9
pxSQC4nJNHez7TULzpSeT1G5FKW2uVwRuGBLRs/RCGOcRuyo0wlMEj0iRJXaYHU2
AobRCLbtIxwQYX4XjbTdkJaMW3aY41c1qTipqW6ZACC+QVa5Kqr50pPpFZ5GBhCP
N8gCzp6pSAg5gHMeP3vQPWKpn31feATf3ZdMQOB4cC3ADljYxqXt8yhBdriOcOL9
bPuvTYgmsU4VA5rB3YdNyJBiZbc1kE8c8yAnp2q+fgK8/Zw/oOEExTLMkEOX5XYF
BaiTE1HiqO0DZmaGO+OnDdsNC6TlKUzsBhzyswrUESk+dgHu4qX+91WgPmiuNzCn
O9xmtzrgRWD+mgC+zo9sElE3ulgQVrCFaGp77D53TwTJAbeTXRK3k5t+q/TzBSSx
tN7PIrG3jAwfpt4qIYwv2Au5M11HrHraajOZXk85WxNjL3g2M5TbJn9hblQhacv2
q7crrqXfQBVsLGGh8dxXBWPlPYVOMNPNroT8hY6JD4eW1rEVofqk3W6OfQoHcGXj
LAwtlj/Gcb6EjvQp52bbRvXpm7xNRWtP509PZZ9h+kFRakZCGY0J9S94iiNF+sbv
Xd1pEcVqB0sZy4Smp9pi3oy40ZC21tTr0oMXwJqr4+6UeKkSPas5VLPHK5ZgexdW
6bjSXIfoPhGYMHku6O4XU08oBF23pO/OOyUIwITNlpqplr5lhyiUFQ0owq1RqA8Q
BpWzbGXR0CIXr6+/AdmNNtYP2zWrc+RnD4oOfQnWExgHlUlstcaJN/MOU/vO/yRE
WLZ4KoR1g0+WQyIHw2cswJcAdFjXFNBKqpoWKWSUZkCd8JY9h1uGrpPaSr7xN0jI
y4MyOJiQXFkHmX430Zz7w8WWOuPpb7t8uFewKkUZnEHQKwpkAcUXkubN8VFdvfDW
/yyAmZaPQgfXFycPLsjfWXWZiXN4NZ/jxoHgTCmrCO7DVqhqC2420rxjRoUa8Fpy
700yGvtR/x1fdyxMyI9vgszkgNXxcxDxt4o3//CozB0U5VZXOCU42L8XZWMjaL4u
JV4V3cl7MUfO61E9KNTnD9qSIbHE1BL7/u+JCbbtTA2MEQqDL23GbK5BZG4mT/uV
bUCEhTAwkfKnbQrz8wBIS98obzyTgVkPxtHISMGNpmg+IWaLr+75ttSDR0k8oqAr
OdSScAuPpaGIhzQ6yRBrVro/JLgcK/MxDz/HoBPCLDzolWF6cCcO+N4nKZ2RPLlj
80eLRN0LT+XqE4vvP0+wQaNTgxmdC6Zy+TLq2AyvwOO7tOt/F6fAbyxQG0vVCmWM
dw3s7MRDy143ArIE5oQleNy4iVZm6MVyGmZNixESK0mHrBBVpHzrdqFp6Qx0xKQE
c7QzuU/LIMuMOlTFFJOYHaShOtcFHyN+x5GC5QNHkv7+08eVw7HWOIwxD1g88lDX
yMZe3lLK/GcWmlCcPEzWq1bP521hqmo0/taS8dsFHNogaJ0RHbg2uIqfcD72aRLP
4qZ+ffbUNkpqM2ebxJ6Uw4e83B12PqBw4TC8GkpAD01E16s7xNM8+A+FMirddWIc
xc7GDYWW0o10qIoSy5pZ5Kr7JASd7/ZbgrrorfEMgXoR2EajTnRhpEg4DJ4O7NwE
r2Tb4n267nZ7fyWREi9TNmU6In4gzgsJpUVqKDklA10jVmDdqn5ijNNoDZ86p7oc
n/sU6NkjlHKcJZqiYjn+/DGVVsHzsJXi/kpM0c1Civf3T4k8jYC54WWNZlTxrDd6
pKvv3U5wV6rnnFrmkfdxnDPs/xnpLMih0ciyTsX/T8Sjaw6BVXpKg4DDHhh4d8tE
j8ZBCKPD8TA33fRtIEseRN30MTFgMqjfYBWaL09x0UudfePyFaMYSOtAaa//OQCQ
wr0AtxoNAAc7M8mPDZ2TtOZMnFLvrdtk5GJXEWsMEA4grdTKPvcRl5Xqp1tftQ52
xMCiuthZTjV7frnKgPt1sD0HWhtwMxZ0pH9/Q0Ya8V9WeqhOIG2+VeIhOTC82HF6
yg4IJzUTdfRkwyiom1XsXyta6IwMTP90A+UO0DU71vq5ptQ3WJcIJY7vN+3ihjQk
Y37D86rtJrms8/zwcum0Q+UJj5BKWDpZMeuCpfUTlJA68F6BKGoupvP2qqsdHwyq
/oqe3lipHJEK3/JfVgg8lZutqBXyh5n+oRtYPa2IWCwLbsapyqLx7QTTelWS3i15
6Sl6iPb/vwCu8OH6u1KcSOK76MdRFIyoK4Sr0W/+/Sm8I3dUnYmKgFe0OE7N9EjD
lc5x+r/CR4JcMz/THjYS4CjE7w2ZmyYLPwz0hOZKq+AnE5pasxBXq8/dNItLDurK
IcoxWjuuy9eopzKYBap0xGLn2VFqT7w6f5hsgiXkfO8l2tb2Cw+UNZWvh6cz3z0A
mLjoZq6JTSC+9hZnsE8iK2FElPM8KxswgrM30E0orTVTqBw0WFCOi9d5UwYJTdms
SzI6sf4NdvaZNeOx37JwYHJftQQ1ZcSk0CKZNhZJig7EJ5jSVl0kNtQ3MYXGF7R/
p//bYnPtkETiW5KTFVom/jz/6IefNGGZeF2FdTHeeeWXWCBL4ba2zQWqZIp0QTlS
X39NvcdoBjVU2214mkqErS4Er29shDnV15F26qqnLuT55w1O4u85N3H1a4PlOfFl
eQQrEHjmD3E+dSef6MTZ1unZOg9g+GcVd12fE6ibOKwTaV/E7DOcHypsTeGr+p7n
ExoWWizxsMWgDl323GGxovCFRWdFyVVD7b5Fmwpm+Ygf+kB3QPkcLhaj3dMgD0mw
QxKazvh25tTP/65lbmvBzEDcTsOutvGUuW2IXyQmnkYKMyYtLYnKiesifPgwKGTG
leU7RQfa8q66weozBsmuCLviN+tsftZIoPYbCBGGxqMVjIV/1wnHDP716CY9lqs7
Sgd1XEi3T/nH/gvTI5/hJcyySSJejAoqwLqcJFxQUxQcEeE0P35TdWUezCpcUapT
odTPegueEZanOWJFXrV1QYUGvpvVPORuzGe+JjtGVLwdnBn8biRmRyI5PNJchtrc
GM7oISLw/aoOKidlIF78E/s+hWySvNafaAJpBjElhXqv2PhIyn4uqlTui2lR+jJq
1q2LZ6UzaBenOBVmcHin+E8vP85duzwlUfAm4l9eLWq93sKG1uGHXfFgpiRt3H+X
CIgDk7oNAT7fJh3CiqqlF3W9Z6xYsn84C6mgCXB5SVpaVJ2bIAWfbkQy6NUVT7lM
C2ePtwK20AMOJ3Q6sbPyV8VGA0QqDbdx0nX0IHmIAWxC+5gkC3gGDUpFCAY397vS
nMj6GkUPVfRwmBqbHMzeHa+NR7Vkt410tMNPZqu9oDWdcPIohtbYxfMQNVyeNVqK
zxx1e4j6+BIr17dVcVzDrIuUqe1WR/bh5q+OTtvyDMPtTG++lerz2+M7bjsvaQjw
SF774bcEWZ+x1L/kIUZlipdxdIJ+ww8DKUydx+sZuwoHCnSqr/n/JQyCSIMBEdH1
PlpRSsgMEO4U0qSjSByaDKNkh7cjA/MZxOMNnLtuZIrdjZB1QhiHEf9gYRMd5+Ai
0ZiBnTKA/A7C5vwmyL1XhzHv+b4BtjW5AUlB5A+9Rmlj3La0rSAQgP8YAixXzDT+
kdTev+Fw/76o9qvzFDgX1R14rkqX03Oqy4xq4qavzp0lmmjKkssODKgbnnmVLyQC
3GbZkvhpZq+839T4iSLDwpNRqpXSU5X3FMhlcRbaBsl1ZLzVdAhdJwFIYCIhg7AS
VCYyVM6Wqf85o+PrF41eDrY90dYesnHb4/I8Q974qdWmkFxeW61dKSQ6OdTJ4koN
z6kdawlQLrtRm4mDIR+0S3s5VDkV/WNxy2N+SEE1joR81uKDZc+aLsTPmpFHx2j+
Q7aBQ8gB0KRDFx4PNgaFAuxtjs7hMpLuieltDtXe7KF7g55nw7iZKl3lNzIQuC2A
RACwHiOUuCPtoxY24X3Oo25ExV6/X+ZBf3U/1r9NgVODnOWaVnJDMWqKD/F2koz5
/RxZv3DCC5UxG4vgY6KzV3IRjoqVWcG47GAo2ddo8u+D19srjCWTKek9qXyYkC9e
EZ8Q3GHmjapqCRPMMdQ5GscUmqnA1mhnKWCazszI0PbzP5iaSnEm7SWm07Q3zzYd
qcoZFdQSXW1CubBE9+TVdL+kBVQYv465VeseoI8lLwzMW4RFmoAsgNo4ql4E3TN+
DLlYIT7Ce7U9MM9qZRDaCmfnO91XM0Ofiga7n4ErcbOlCBGingCVJdTO9rKivnKK
n5ZtbDjhoZzUkOHyTn8BDGo2S2xyEsRZyOaCYGStv6dQ+NKKrc1tdSdsIok4+9zz
wtSJo0Nli4rV46U5j5wLZmDpAWmy4+B/ppWLZgEtyuwPnxdC+uaOluyV5Oj3K84D
c9zjVC1cdfweYGCa5i84Gmusuw/rqDfzf3/rjfGfs0MXb8RI20zst2raikw63y1H
xajp3W0zAOMKwFQSz4E6qGA3SfmZoCwgdoXRPCmhrSVHdNI9o89fGAxqJsf1G/bY
5eDe5i3AvcSr5465Pqpvxw==
`protect END_PROTECTED
