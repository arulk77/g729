`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveK0W4wTdZwNU91cgeLfVWCg9HVcpnPRGgo8lq+nMIK++
UzKZZ9IiLMHIukyozHwBgTrlSSoH0u+Ei/52dZry+z4shE0wSXu3OpgLhmbV6dVM
8XxrlnfEe64Bobp/VJabl+rdIhZ05waCk9S8iv4bQe0IepzDqDJgL+Gg2NSdnz6F
Fv7MdmoZEF2jbBtqzgWowbfJi/MlszJxoO5dLC2JhideqGkxsLqU0NeqI5jZsYD2
JU+Fu6k6UR8kwJcVXwYGPYlXiALODBFtFAe7vfO7iGEeydHJ8nbfYYAw/y2UqwAe
eA+PDdDAORJG8IAl1/5Gq3J6ZETB+KNmZpORZF/ZSvWxr501Z5x4eJ+WzkDCMq5k
`protect END_PROTECTED
