`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkY6RlrexlY3brdz7l8S51KY42U62GeG2hyRJveYOjBZO
FMUeahZBewXQF7I0mWOPcAzCEvT/9DCNvItCrEFwWIwYiclWPx8UXQXGaunHRZMT
OMXJom6V2ehs7zHazQohWbHmYH9vQFgiayyya4pHUznN5qjP7scsY+QSIIhiQQ3V
dogNhwWH0a08bnecm4IgYxrrXAjt95GGD1I1c+6md7HShuGFzlnAmMMJSzC/kS5U
wpBgT1kYYPsMUCIlpy/RXrWiownuINhotL+FwQud7RjHHEYSrC9+oc8TpuZhcbDN
a2Xf/5kj3LjnFuowve3UN/q8Z2002aC2rtmStX9h030=
`protect END_PROTECTED
