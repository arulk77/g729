`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C4yAlARqZHz3lnVZNnKiV8moeLg87xFNY4j4sz11ZqZk
Iz8PBVrWaXGEIrFGquo/yXxObYJoohEpJ6/wb5+fChgdwQnnofRPIoaW23wruUHs
AMDSjl5qtrnDcAFHVuqNkSOUihoKgrLUIlRg6Ahxf9lpSnu3zcpAazpDrTDj2MKf
2S7I/lePdFwj9amOJwTEsGKepvpmEV87tU6mzNLmYLE=
`protect END_PROTECTED
