`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDf/HXeLKSErlSUaVl5aOFsPb71yeChIBLppB3x7gXBS
cmRx2NzPsTc26+NbFkiVdE3UzKUDH5GIy/sej2PflfyX9bqsJdOlZp1Q/vQpPEvg
eFYzLMu/SNk75EDNJWrWxwTEKfrA4WF6DTLyTOKLYXBINKoAftejPUJWuUP8rvtP
dqjXJItgsP5o4ehCNT/4/bdHQdLR2kTw72f2cc7u1gGZ5VLbH2nbSBU1xafrJ5RJ
gUZ35Rr67tI50KG2xPPfZQ==
`protect END_PROTECTED
