`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOhFkS5IqItzoXh02p6t+EwKt1MAU4upd8vYG7EKnaCn
H0l66RPoO22RPNj1BFCmhyRmpezHAYtt4i3/Hl7VsB9SJsUwAPMtzP6cQ0cgvnj9
FkSVJqguzvLNPhIIhsVO1wJ2F1L3JMjcGxMLgH3WtRIjzaiYsAIrxO8aA4Z1XEvD
YBj7PXTQhJBJGQkmi3PEkA==
`protect END_PROTECTED
