`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGFGeGFt7mxdMz+1n+ktCJ2MEpeXCzqkN+4HWA5lmetP
kodufrbjbZlXYUwEBhWLI02uemLsG7zv8iFpns1ceFNApqeIwccJ1vh0Fb+EfeI+
n/MmHQO8q09Rh2RfjjHFzDHzxB1K+djbrycYh6953TJzh9WHQ1ON8hk6VK0Ky9E+
QIYPtW7X4u7qciP0PksJnERl/gFuxnhQDxijiZHmoULpgkKawywCTJFIlhPyIsKE
usiSh62lkR4ozmMf5I3omk8L+xN3spt/JpfxVeMvBllFGZExE2xctcn0RELtEyxq
ysd3dsNPH2mTUSatYnGBAA2nBLfEgw/jlqLYH126e1oNUSIfWnAIB22veGNz+ZzQ
GzB2+uzWdkzaDNAtq2/mpg==
`protect END_PROTECTED
