`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
TszfYWYzWs6uVTXemQ4sgUnWpOX5DrTjntXBVf/qXAfgce/pfCmGrvTesEpMaW4i
YfIbiiDF73pYI4oyaSOQ0mwr/WWurU2F6R5TFrAlWhFBfepXELwZKcY0t1otXCvu
y1avSjqQzK/ZrzWNH61g01Pg/yMHprwZpYoXwgI82Ime7XmubIZo3wcUkFH/GdoM
5aURkyn2StVBOOro9w50Y9ameeCcoIr6ZReU2Hc8hZtqWApn90HYgANjP4J9VptO
cdXbLQOiCvwavNovr8k0ZOgCxdIZ+3aSuO0DmtLC1VllkGxqcEeUUheUnXHFkgSY
dQ/tmd7XY+uLTss1YyLOtnoiow5CnobKe0x9oEa1lIU5PhT6RV7uzKmmoVwE4dI0
kVljWHLSK8rhH2B702/x4TV6Z9ha3rBnLF59Z/3AYbvO6nWfF9FIJf8v27K7udUD
kd0+2A4DE+QoCPyVrKxANjmB0o2LDJESFTM4Ea2Wt33mfeZ8rCqXpdFiEXCy2gLN
LFxA4iMHe2kRoODE5ROLAedwuQh5rDbXuwWUVDpXPC4g/uAwEm6pZRY0/eBXsD54
I63g3ixoZaWdhxYDiTipKBcIsC3hdDgPzR+U/oXWwTa1UVSQstI7hcTz5XOS8Er6
b61KXDf1/S0qwA0f6h/AAGK3/uTFuzsXT4rC026bIJZbmhPDmxmnW6lNt2jky2T1
WumIU8zCDdN46NAyvMPUsVcDXJzAgH+8RrcLIseBjkbGApYAxBPiZN7KPNljILAv
20oHB4eJNTa+Ji/ib/wnHuUnDi+kcXBC416cQGdD1rP6HZnz6QHfHUGtiLndL2vW
+Y8fYO+aW8+iwI49ribJHIovFd1derK9Q5s7r5VAJ/GRQsNVacxqyxhyj6pyJVg/
h4AxlEKbME7Yyfp7XnbxNX9Weu0Hmnljqb1rSg3lOdNdpWztftOLcdSgJMFLQntD
5/U8lgAeEWnCuSVeUYkGYzRlYhBsKtGTwYYuF6dJHLHNVt6qbxaBIDorky4hro/c
aCdDYICIsV+zIO21AMNbG7mdocwu6dLhNXjoBDs5KL7/ayeT/F7d88/QcYQZ8Xuc
0HNYh51D8fK+mHKxj4MNsHL3iGQApUGMha6PoruI53rydoq+/vJ6n16eZfw/ISFP
YVPabNj+iFgZz3xh3bqc2HePAPsMBFXWGbEqTtuanBJsHfioGNbe+Uh5khDOHoSp
p0A6Z8MR2P+qb4p6lr2MQHYTUTXRHLvdnIfETSAbeoJRlde3BbvJIPjrVd4vdsoM
HFqIz7/grWa5Sq/ul9LlFurJWByJBMpOyj8jmuO33mIveBSZ2skWQ0eCKGM4SHk3
Inj+oqKBwmgTXUdO0Z6jEkGoPOqgTVGy2YfEu1IEcZf7qA8lQX5oydocUBq8hgQH
LjUqgGly7KLNqYdyMxBMZ+LEFXBCum/b8oDCYtdlZOtcQ9ZRXn7ZkY5exNrDWCOH
gPu2DFNIUVtfylp1FxclfLq6HA681ZXFUiwuBX6rFvm0jkJixVUrgklu4hvetII5
ShkZvAHFPYO7C91QL+dZptkzeIWlf1Dgx3GdM/k+pZ+i1GlDphEByuKieYn6J2QH
JqOhGanF7/+g/24gGPQLoeDX6ms4aifWqTKFfnA71/AjVsMLSTPxo9YGHlAl7mHD
YvknlvzV24fNxdaoi3+MqN5sQSnY0hJjSQApPwY92Jb1kPg+Nuu/NLrY8QLxRfhP
6WjVEasGC5IMQJVwUlYJc0xoOO7bzj6VK3FyjZDxJT6U6LfA2Q6rWWYwkftzgXqc
1DlRbHQoU5H2J0jbP+TrbDIP7+YmneS4HfssvbUp++lo6QBdoRP9LBQiGsee4f+7
Z/ZaGbhTIo2ahbMBJBgwsISSgYflqbRWlGXq1gK5DGJTbGmKloykPchNiuZ2439/
Xzw5ayyyQ8ra+G1Vu0jypdGD36bO01KsHtbKYeH4rTaxaRyFgmuexGRmevECLoO0
`protect END_PROTECTED
