`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJU2r60gwPhWcVjfTU0/RICSOmMUVhH+dA8744AyzUfS
j+uySvvLhDecGd6v3PaQiBOiP/5trVO0jKM+eHB5QQOe9ooICumdyvTJiKRno5k8
eRhal54kHGpxNIZUA8XxEd1KuKsczPD/YV9oz6xgykUrk2qDuDWFp2Ob2/MGSVPA
wispRDi36t3kK+g1Cxc1O5zQT+vMjZvU5JzWWpW4ZmIu9x+0gA99ykv9VRpQLL88
`protect END_PROTECTED
