`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+hBnPhiCBbUj5vpj9WcYaoPtR3Xkbhb/ccZtUz1uZdb
KOqC//gw77OhDFC0mUPHRW43PQqAXX5/NZI5CAxHqSWHC3jmpC0opbbERSla1P18
bQDZm+zoIOlj0Fvd7PbXOjEwz6KV6zRggSO/7U/ZSsqWjOa8E1+B5CiDwzn9JEET
3MkQZrhCCJfRLn//8fGAO+SQxDaFj2Zk32sxWnK9WmOHp+8lX3U4RTkEYfYOc4Iy
xevU6oUSTztUCpqwXRiInt8lzoqPVG+iTUvqaVsy/9yaLuOw1UhQXHhOaBNib0CB
iRq4zhqN5IQUMPpIhYcyYeuQogKy0ET+oVsGawsraZWS+cO7a4+DH7KSUE1zBrgs
ZMi9AixMK6sWyVDD90ZHWysenQro+LP4elNInIhGOGJOEM2QW+StL/eAgqPoGnQq
S5XDVwX5eRw8MHm6/xQnZA==
`protect END_PROTECTED
