`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGpK7XpUZFG3iI/6ojbxzwAvG82FM/3KX0lGGYsTTaXN
98c/HoxvMxNSIxDb0OBfitp/JJuA7k5HkmAI0fdOpL5Zh3DGH7Q34qh6jEYdM6Mg
0PvOUSidifHJE4rmu2sIi0vl0Wvdh/MTMibmqp2c/Qit4bAf9ivqtnFpzeiOtQ/o
tO6qeJCHQjx65vntWkCIPjDX/053JPG/BC5PFu2Zki6USl+T+ZwEL9FFeTVRkbJ+
03aXJu9AQxVgEzok8BrEnkSyfBfrCR9QEkTtR0upqzjqlscvkeyaG3BOrtA5zWCp
CdEIWybpzAzfPhpSazXCznp+ZSTrknWGW/6g4M2z52vpvC3L2XeH9aGUSCY3xr/w
nw0BDz3N4c6HkIKO3jZhdkYFviraCYkHqKhEdDi2GzdUfqGo7gx5ZMTaJnaYiKK3
`protect END_PROTECTED
