`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFl7L4+JzrSUYISQ5upS/8/8p+GPD6kwFbHL6vhbKILT
9cUhxyxY0U0cGmnkVRU3VqvGlotAJgP9pJn9hGeJQgDQRyxGcTkuk+EUmHWdC3+C
Bkb3RbuKCA3VSBTmoGIB71D59IbdrFdJp30eWfD5tq2dP+JOZomPDODfe6YL0u2T
zAMTKrkmZNp7QqBhBtBN9CD9XCpD4Z39Ca0rm5Jc4s6DMuCNNca8nZYIEAsMtnJS
1ZveXSwKTBbzPXmFF2BBdDFE9TeNy7q9ILALAr3BoYjKS9T/L0euW5Yd4cP78zD6
cMyZb6UcEcXXlonGuGiefAYEz113mTRJxZjF94OGayLNJnAUcNXqX+OXOCd0LESQ
1xvFVHicgoJy5UlxbFPjffn7crDt+Mao7vYsblWM4OHO1sTyemiR3esH+moyfIq+
OXZtG3WdHFhDNizlvnoF1jVlJ4w+H+yOAwsnmMDqNhQGD1dY9zxEdWRlUikZYzMe
1byRbXXAP7qbqRd3iX+aB0y+DcJxeY6kKuhvFtE9Luy1aPMiJDLRaKAeCrHFBGni
ykuTCWPlc7JKKFWEioAGfou9jZZVhPjC6lw9ju1lod1cMrXyurE+TDlKi+S8WoTx
+vnt0grbsucCNP7BOTU13nPcFRxmoNNJW1HKj7cuvnzw4xnprYg/EtGLbp/Bfs+F
JvYgQMew2RwI/C+7MYLZT+1ifgPPvnAm8LCj9E0n0J3cByVyRF0TnP20x1iV3ndS
9bSlpvpp5DU3KdxCyIG2HIfYDKrVbYAIMX+2izvT3e0=
`protect END_PROTECTED
