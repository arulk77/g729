`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
LXTkkWG2IGhaNidCeL3cj9Z0LnurqN8gLh0NuNnzBwqItyWYa8tey31/sIeWVNwi
u2jlTXMZvrUqF7uZ5tn9saEVSmkOSeFZiwCL9VVaGVru0iGYZnN/seidJVAbwcXl
xwtmtVhkPpWAupm7QWyhUUC1G69r7VaQPG1lR30+bgwS/wSguA3PAws/muzSEMuA
`protect END_PROTECTED
