library verilog;
use verilog.vl_types.all;
entity LUT2_L is
    generic(
        INIT            : integer := 0
    );
    port(
        LO              : out    vl_logic;
        I0              : in     vl_logic;
        I1              : in     vl_logic
    );
end LUT2_L;
