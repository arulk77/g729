`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+VE60U1vRaCOV965MW4aRMjs/zJmA5BkENwbFip7kim
yYaETj6KStCMaG5OC72GK1wnEdQ9Xe44OEp7KgpQb80c3LW8VOtMfAQ0Gi467D6h
fP/DEHkI4xf8/C0hjGxPFDAeO+cFc5jta8uXL+CCzUVsLWpVoRvIa9Y5GjRxrgaO
QTDR6AhRC1hUXdPeC9458kjogHfiyz10pxquSob0f6GPGJaydXIA4gaSlpMqxHex
yhXjGRItPJhPkq2kpBW4dHeXaLDchnWsoj7OEFb5x0U=
`protect END_PROTECTED
