`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMFe7iolUEbEutCOJyf5QOswm15ATqv4uHUx++mUsuco
kcwXTjN+36hdehouV9BxTP60SX5Vl1QnlMhexkN6demt2AK004V8yaF+CEBF8Vmw
m1iJqMna6mgXbGAnjJnob+F9RPboZuVEhuE5GKDL8Ya/ho3asww1Mkb0ndW1uFSL
Ruoe33aLa09rBXbqs4zSmyrG1zf+Fq5uNpmMp3HD4ThJuYgQZw5VB/PepJq50cMG
r6oP2znjHfUf6Im5ppqPoSnWhFqqZR7cIun7Y43/uNI5kYtmSV3OACKjUnlBF8fY
UsuDX91NJ4vq2cVOaDUw3sdAnvf67hYfXAPkuMP5yBbHdsEIBNePoP+2wLI3G2AX
Q1hSlUqXZT/ApZof3R/VFvXz3RACLmKKmxiUGTf5jO2P538HELvpl7r5PYZsCBp3
2the4v3vbQqlKwbv6t+uFRj+KmAyQjG0zT2JIJVzGdxajB5KFv/vBUYOmLDPk5+2
e23DE4L0H/94Lq6oCsMCLlZcaMs8QyJbCn0GZrdrkTTQduBZBpAfj1uDVsRkrKh5
xzX/KAWvTv6To8p3B3o+r0pMK15HK8cyzvpq6HEY460fDt4v8TKv+Oup1KSuaZ2H
arHPKmaH2I1g5K/KypiqOM/3nHZ/jBeo10v+3p5Ojnnl4cye9wnjjFASDXpVocOF
MznRwQi7HeVwiv3ueg1JlTpVr1kG+yhmXsf7SfF8me5yAhBXHuGIPQ21Fphu3IJP
F6eMRI8yxUOoGZARP9ZMnGugJ+H5fe/LRWDfc9SkJAd0vF6Xrv1EJxr2CHDYq2dY
efBWOZ12omfrCIGDKnwOGICbaqRCg6WVMPjjCNjEsTcopk95kaa2wmDkQD6qrrvA
r+P2l18UaIwN0YHHuV9Q2BXvTXHrEV1oQDYQTa7OyCMQSxOr3JqI2ZrhNxSN5h59
bJA3Dws71E9Q8J5ntjbosgPYxwQiqWk995RDD39tAo9faGNLzFma1N1Pih8b5ylZ
`protect END_PROTECTED
