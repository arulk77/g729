`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QNw40IqJrFvY2E8HYWz+j+6CSySbCfO2/cDpMyannhEPXiP8ZFonkn9LusCkO4k3
NajO1y9pf3E+BLaxPplLqTJw7AOGvPaFjfM7/a6Ip9bPURrZtRwLanAAO+lDml8i
1KZsZj+vWnhxgta/zmEOchmOX4TbRpxdZdtm/wZfA8riVmYc4rMY7vrHZyJwMIHv
`protect END_PROTECTED
