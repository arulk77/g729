`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDASPl+kHaGdqGwGn2wSUz2VPLBZh9mOhUkUg77aLvW712
D3a/3cXB9UlHxyNArNFXZYqC0e0NiD7QyGDb0k/MlPRKXqLTLRhcJ3mCSWxjo2RV
SR+jL85t6GTS+pBXe/ywSUA6UHw836ElAEnd+VSgSoUjBjDHP0YfDUNHi6nuzUtg
S3JBGlgU020AxgtQi/z0XrGMwhCI/woHmEk2ifZ3k30TSh4MGyJIxwM/+u+UIHQy
vZQFMotjkhVLs5DraOTmO8tMbtAVGDAqtGtWtm9kPiQJMwKfW9Oi+/noQj25MAUl
fQuvwnOqTWv1Q8hBaFkcOY2cP9yW2HDhGj4HVd8oG5kF+oEb/hR8smqmN6gTYTO0
ZcJyq4C+KkSfnY9IB5e9MJTA0OtInkvqlIZNiQ13hFr33kGgitxGsRX2+zNixxjE
pesIKxzowrtbkAOPiW9RNygTV0ndRtAoYK4K3abDJ2/40hkKLfomXXzUaI4CaSCW
K1Awqe3Asz4ZhUw896DeFRCiFIYVDRwseJ18y2DuVBJoJNjE8Da0S7/4q8d9m20F
ZRVM9DZJscWBoUR5g++pxhDnwLfbB4mHgfcdDbF6Q1mOJl3kCfb6DieTarBNdOWW
PNAik7H7ALN0yOyQiqpf1pmbZywvQWwrteg1QAk8fOW01oby/mqbCbHKu4yLb8gy
0rT1P73DEdqFXVMEFQNuL3oQKTJQnDwXRM18mcNb/THv8mtEo/u/U1noDlye6ZGE
OX9kHhqPq2eWPb9B9ZO4kxQ/EPa48Yb+pfZMye2KEdAkOPnYtRzFbxMVk7Vxbrax
ZPvHmpfv4BPq920vNyszK/UHMRzJ0eWJsvy27T27+zN16fJh1if4DcgBNHWKyY4f
q9glMU9NAR4ah3qFE7XyKxNVS4vu5mZ0Bj4187ZdH9OyOjuxJLJsSmGCDNJ5Azo3
ljFKy+HeOVEH198Ymn6aDRXoaBLeRZH+LOUk0E6YwPM3C5itc1v0h+LZ+oiDsH8y
ukP9kUhl3XWDC+iTqGwnWrS3Gxx8WCEAJsBfGFKQyc2lxDb2KOml9CVmYmj+Pdi1
E7XkZ/AcL97o7HhTh1iR121ZO4WyabH7k+7oVHCFGHDCEXoJiDHFR5Jo2JyQlOwo
rl5xPlar0Ep1z6ugl9jbJIRwyeqVzk/5FHvL83ktoveIzePtxCCGiUBnY0Ab4p8I
z8nbIFHmwnSf4TGE5Buaso55vBZ6vXKrzUcfz/Lff6fb0T26JkTTOtFTKZcODv6Y
RerLsXCp6NnW/aHW732eCRJvbwTR+Qw7xXO2PjcSgcZcyyV0RBfs0E0c+th9fCdY
3l+GnRG9BjxnKas4DiTHfAlXNKlqWMBD/oQPOnAHEQmmHDYsu6hPnhZnn6LpMJ4U
NwT7UNbU+pPX4ZePxzxLoYnrlSvaOQlr4O7Q64S+XQhGYrf/RHMk57kACx0K+sTm
Wogn8PR2BE4d9V9Cm/l6aTud9YJbECC/KjS76CZDfWSDsPRM4z8z8QD1J+gYsir3
zxo8cY2i7VlAPrRK+8ux4TFCNexfnR53mhW6Rz+hOdP75X0ytKL5AyeSGl8IzC0t
GWiSO2EJJc6IcqBKqWp0RlBVJSwJKC2gn0xTwU+D64/3/DeGadj7h7XSHlAoHy6Z
2mUNTOc489hFC0Sv5gxEEm2JTIpi+cr2bA2MHLpLbCzkuXJ8bSbTHFZVfoZBo0lu
JDrvmgB0rnT2tsNFtTSXhL5EVdGO7X4lg8Ib/+8NewqR5whuShj7/8GxvZBJWrdF
ZWLE60rzw2ySfNsgWPwU+R93qWZJHQQWkN8YPY4s1wU0hNYrqpQrMNP/GGvvVW+I
cbDSRKKde+T3pv6FqiAWSoTXerBgFTUSx1kh7+a2MtvjaRq4AAxbfoqZ06++oa+1
F71eq3LSQcrUjGl/V2b/drHAxcDmhbaLyvTLAXuf2woZ94fI3YGkP2clU4KUQ8+I
tkcF8BMtWP/RiT42QMgSu8fNoiNfhI7u6ah2sG0salvYCPPzng2OyQIhucHq3yc+
dp+Dz1aDdgMIhjz6Qs1h038i5TMUlhj9A14ReVCB5IDMvcLsUs37Be85Q1RBHFYQ
l6HcENNlq7sOZcnRaX2+AKxZZaAl8k5QhMZeWyx6FsatFPfPCfFlQCLfOm2CtQEW
HoPAXnw7y0i5Y0Nt/BJD+SVU7UqjELSCKN/gEYdNJEnKnkkLDBOqsS8I/Oer6vxk
Pu7eVMdaZxeUxvheKc//snRyEHksHaEMC7l5G6210qW2PmUnz1rjAURQ/l487Snj
Bx2s9xqL114Uaiirucb8qfsMmmsj2NyfLaq/J0togyhoJc7TGHCQJQQqPtyO2uyE
HRxp/XLYzWYrleLwL7COXcJvi75x/1SVAuZGqMeltgf4yWqXKbfTPJBmaV0MWjbv
jsvl3HDWZuhTXhCLQMX9j3g8Ok0YxNHN1sLi58/hfD+H8QmOenGTG420RCPIaSnX
QPajNr9vBbmVxVVHZTMK3oCg3hdig65JHdhxmFipUnY8jR2wnWUy405XIE65RRYz
+Rj4iF2aQMyL+b42kI5ORfNOIE0G022gh+ANufHOaheucBNgJmtC4+j2BatKmAa5
SEEk9L6EGIyC/PAT+0nyAD8xEN/a6RhinFXAg6JRTFYCqcQaXj827tGGE6EwmjVc
GVl4GhAczVESrNmd8CKEn00hLXmXLWHUafIFyTjZzDOs2XFdTlTS6vjQX4AknIfp
E+CQd6Yz/pOd/o5Nuhd21/sjWvImgmTT/xVgzBwIye1KUeHlZBT4mkbIy5jQc0t3
wPBNMfOszpCVaoNkfU50O+ckTy5xU+FMGHpkrSPsArBPdeVG32u1RevArf9CFXfb
H4kK8qZE0A9FWzySewbKh16B3524+pf9DZea7vi7p+3fCNgrEouxuHQNA+PFAozW
Ziq3kE70Z959/bpKf/2dMtiX6QOYoAnlRKZr0HF68PR83nGUA4lkTTpwxXSBvDAY
2pIlt2VOz/8r0xKiFWT1Rnb+7xmjfVBNQuyJU/d2aFxLZ2fuE4SPS5efFMXV3g+t
1V0aJ9ECuiYHxHlimhWPRymJ8f064qTigYxY/Chl9P6t/di2FsWtRl0qCdcIWueX
auMj0TjHJ/J3m/1P2PAUMFEAo5VN5EDeIProt8omh6Vvlyd1emNKnm2Yh/6WsB4+
5IZU75MmfA2aGVwrUB7KjcEm3DvC0q+6dZ0YDGzq+sryCZ2bLb6snLVsUSAAhjvt
FwRseuMzt35hD5QP2mrh4jdGnhlyA9DZ++OZ8oH2RtlMHTGGgkKxa8rs33B2eeSJ
qJay2uDT7yNVC0QOEsbFckXWKpm8v7xnRQkazD8eRo9gzFnpggEMk6qyNVaKeoDp
K3lkO/615iAT2iISt34md2itaHVj6krsfAL673uh34OpjLBUdCE1I1ZH7OdymyHa
4PBzyQaix6GiL/c0XqGLE/tkEMEvizTDRqA4eRe4A9a0WSvkWPnY4hSKpU0sblW1
BKW8VgzsXZEFHMT1DiTdM0QBovq5A6om0DfUvf8itaNZ4BIBFU3tJTyjFk26FDzP
Y4vv1WXth0c+l0GcnebD1sYd3kZzLVSHzrb9uzL6aE06XmJUTSM+9CTnbFIv2JE4
u+Pz0mLuyyaP6so0buJ2DeXTXZfQ1fOjiScuM8LW5iTz2UL8kLOPThkJsS8mg/3V
120BbHXAXVoKaTBdjTImRhmnpRAPJtvS6OFUvM9h2vTYLi0wr+xz+3gsi6hLDK2v
y6juyT1xVLDIDJgeA5GqfUQy0g/MKLeHWs6ipe+8Tjb9Kmw1E3ofP1h7GMmF5isk
gxvY2N+lKec1SLx6h/0YJUjhtbaMhgH1WdWuJVQfPhhl0XET+dJbMaXDUBMAI31t
ddGipeMEw5ZtQs3JYhcD0Z+GSOkmrI4FfgE4XaPFL1luTg5oj8fVpFuadAKFnB2j
KAsWXcU/A1JuLfE50R8jZyrAU76NpmQPV0BkKP3lT8YVHPJEFFQU2qEPqjz0jz2t
eqrsCxQiTwvvo2SDs95paoL6Oe2fdtjg1/+Jw+f8sV2j0Y9u785q9svrRCvSGrFu
wYhEMPaF4ZpIxk85ySyHv0OmkOiOdWApIy45BbyEZOBgtYob05kLvMuj0KKRhEvG
qXKgn8UJ78ALyVPg8J3rrkXmPHvfOCkYJzOwn/QkuvnkRBu+pum9vOFpQycUj/iD
fT49Le5bUjvDNIgUS8lhQqWIeU2Ez6cOekmi2N1jMVHtFwwYQbvcP9zsVTkOnW+F
USXOAnRKuK04JKj/4lb25jx3R9zIcpu24V01a1k6q39pVyLJSCh9qvfNW/aEA/w9
Gy95sJh6Tir3tAbWveOxzFYUq6x5m+aed8clb9yyOix4uCS9/eGv7JsQNAqr17g4
AjOFRR8BT45hLq3J9cabrHoDn1vankaIK26d+Vh2NxpgvO/huEm7I30RA8aH9Hly
QH6v3T3rfVm/ovN+frB8p2Td0J+9M2fzRIWmZMQ9eCDPSpibQEU087KwHE4C190b
TJIBZsQHiiqO+vOaAN5A8XaIIbMNo3Q2eN1AVD4NWplsfuL4T6+iz5SUm1B7a76o
knSaU+FXjYqEsw8WfIDzlnMYoiX3kzwlRzjPeg04RL5YiM/2uPOoSbqgN364Ejzt
Mz4CT3sSFi5ZNTuawDo5bW9al1z63uyfFyi01iddqLCpmmltXhbDHuRqKBolZ9/L
bIvtL8SkXgq24aEx3LJ8FJvYW4ZD3wekZ3XDfxHWZ2iK8rzpFOtdodE+LYK7dePY
PDNnk9vhqARKaS7Wfy3KA+eSv/V0kYE7lqKHB46ULe4pn5P5mXYc+rYu7u04uvso
9tSrU40yJZNmlrYnWdb2tPU1sA02QIcWNkpUyliahZ9UosJTKiuonocQuEo1uAjz
OrN71vS7SmWylXWfnV3Iz0J4a7Dcyzzxc5eqtwAHrY3yJSPsgNATPKJeMP+pvKWX
/sGFEYvBu4XPDCLHHuc3sOaRi9xO7UGz3qIJUp+8LI0WHlNffphL2NRd9BZXmsi+
RZAukhZaMTv6g+kZXfApw8JiIHOVO1dfX16aw/hJDt0v/iNebJHnYAFlAwJB4OlD
vaX/ii252eYZVdU40BM8INeeu3c0+nkPCeYZByak8Z9Gxn2hjYApj+Y1Pcw7m/9I
a9k7JdVJDYq/RuW85yCEuBVTLC+VT5D/ztVUSTlwpaGeYYA5Z8KErZTbx3iluy8/
FvI3dXLPPXapvEq2LCtUCZuUmUR62U7kWhBUikUkJO7mf5gX01zG2UnWV7TZzu/B
HVqxKHKKuPcGvsx5Ckf2asQBYjq0uXdOBDRwSxYfnX313mKgXVuBBc1hCBbilItj
9beHAJ682lGkZEvJ+Bd2n/YIkTa7GkjHRd5W9a5NMLi35Anpdj/+c7yReX6tctks
7OTJtzjxlD/Ysev8G/rCHORGQPmIznQdxLfP6PTt2XYojlq+Av6DQa29B3snJ/gp
Cho9u0uik75srqmgU+1nH48mnfzfgM2BRBnvxRjFAojUFxTC4NJJR+DcTufkNjk2
ihcdVyekx5Hrt4YHHk8blMO3S2rvEYmCFYMzcv+Ho3xmXkM3uDnyzkPqRyeRGE3O
cR2vXXb54DcKiEpsfPLd11K/TvqtbPJIt5DqhOptWn3SRBRi9GzyrVw41s/3HobN
Nwi8Cx4pOumN1aqprqbLEg==
`protect END_PROTECTED
