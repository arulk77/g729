`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aZxaKRv+MEwoiUWSOPKqLkMBDXPhg/94E/9xZCbHmPfK
ZbKdWXEHsXWJilThhDoIllK5EjVxb/CKaCbo+IOg5PceiCLjJrgFmMMPQ8KplEZg
wP0UV7FGAkOD8mB0iQwXx1ZQ/IpSwUJm11fRf58clClDtuPNaJ2FgQg1sAdb4RUH
12SGMJmBGy74+9cTizgQiMX+oHm8Mg6a3+mecp4VuhM96jTksAtJmThvTT2XyPkk
y4AFYjLOI1wnINyB9dRbsnOvP/Q875NfHPyCkk0G0mWcguafcW/ll3tU+6Ksodc7
7hcUViInOJ89ecBrMdFvJkoCckwX+47FCHt+9thjkiOG9J0zbmiJ5Dxd5rBMDBci
lFxX2usq2Pblsp7Xvvi5CAyGcDO7eQ5d7QzwNGM5fbrU5tJK77jRw+80dRKzcxVT
+XtTtozvpK+g+KDddCcqy6aJiRBMu9Rf2TXEldfd6x9lCmKmy6GkwRlnPB+ovYC2
jufMP0/oDOXCe9+3Cylv6odhrOxTXrshImGiqYx2Zkg=
`protect END_PROTECTED
