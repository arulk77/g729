`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
W52by5FksJUdhgHLv4Ym9FRS0JzkzKCE9Ct+lLa6yU4/i4sc/ywt7snUrQrxByP6
JQdGbzK7Wj1WD2+ZvCOqPnRIAYIzph3dmJ3wYCV1eAASfxGKG9knhFGUL0WeY6mT
NLGLcn+gOEv6Ygw2lujzE0QjZn4IdFd1B9559HadCr//aLC3aPrCBW4BkS6z0GTX
we/S7QpPqr63dKTcwOgTSLkSEoqb11hgeac6L4iHhnFg77u0CSuSbLdcSAofC59W
`protect END_PROTECTED
