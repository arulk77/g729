`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN2oeCbCfySJkvCg2bF1JR6+oHQaBG7rhFI2/Co0906WL
IVC4MD93aFgt4Z2BQCSYrFoYulXfwruMBnlv4kECwkk895AMifS/UWLnFNZDQtuZ
q0axmbmcQwFsujnWWsEHjOMI23MkOhqy1pAKYUKPiNMBYR/rc7HRXjuDXZ5VyAoy
ZrR5jXpF3NNyvKxRZMET2k/15+1J2zJbrHxvIW26tLZXsWPGsraifN48sxn4ACva
UDLAtXwx2+yxWvV1hfwgyZCHiQyXQ9oG7cSjfg84QJMrFSBROMUE2NdLEJLjlLVn
fUcuukDIxLo+dLmegiVvhwlg+3OinCa6Y76LsBoZHrKz21rXrII1crhp3MN58Udu
YghhBkkwPotR040I/gBSMMW+pJQ6E+B/YE4c+G93Jp4y1clf9VigwIZpfy2KN4Rd
tks8yDvbet89aurwVr+YyZrS54v9wUAhqWUsFyYoIiaE8aIeIygITQbQZbV96zF/
kWWhtS4NM1ZLtyvYi6zQ1dTZikpffEZq5B6/f5wzlcLRMu4nXqIVQHRvt1ylQchv
27RGNg1K1S1rqO2OThdi0EW0Xu1K08cNJKgUQ2gthTdYGivuKJHVEOuSZPfsiat1
cWXv62eWZVJLP56u0WaUdxPZ6fB7GHOB4ZkpwKWDV+xcsGAkvuKdFmJMoNab8Gif
M8FQJdnVKZB8qIsuaJh9LAUy84F4ztTN2ZUX9vKU8j/VJ+ShOuJ78DZBAeomWzkW
RO6LAlQ95dGt2/zCva2//pwu8bFoeEpe98F6ioyApXcaamkzdRpicb5d9IZsSLO6
vpXkG0y8d05juLO2wAWep0JMg7e5lvgsnNW0hFJK7/7N90eyLJOrl3yoPbuoJMUF
Bn7rqu15V02yiF1pyJY9j3mC3LN7exFX+EkljF4+1eiZf+wmjxgZHuiLJk22VVmo
yxGHILGk/VUvxpppUDYoq1HV/JUOyfxQdncgYysuXmSkW5VYa99eXYnpU2cxTRDt
uAaLl2etycPBUQA39737lxJr3mjuUjg5He4Ogx9PBDITEQpRkdJ3YuNcANgEzDH+
VI/PFgsJdZlDw9r5EMqsndsuTLF7A+kLJvuA3jd18xB4HSGh7mQVjWA3BqPzCWa1
QninzIDuauGxdTRgJl9ECLCoPu65e6a8G9l25vx6n0IgbtXFHGLTyNlSk85ZyEr3
o5AU6zm9PHx6EaZ53Up6z5gHO8Iwk+fGrzdHB6mslLFn0h498S9/QSBMGEbvVgYR
Ae42NooNynoRRgd0fXd3b/QNrQLUJCZ6l6m2plya0W8GbAvC1g8le9YFVgUUZB4r
AFkCIvttOt7sEZGzSG1wmF4Vr4cOcVfeNiuQpAmcwWs5XxT7xWEh3BQGVrWN0E9I
7hiftS9zeiv1ntNqWnoQQ96cuyYqtcwtCWocTchug7MZEc74qBixYXQT3k6xF7rk
Ggi+nl3hEkog4xvyOs29oyPjsnVAtc4eagOYlZMWi+oXSHipCrLc7UTifv85KJVC
`protect END_PROTECTED
