`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOgoJ9yxI7zO8VlwOHPRO+/6dpq3L12HUDbxyYTbU5bV
KVD5dYqzctw8SX6yWDk0phBRRBJnLcMJvkcA2Lt2zRlHXVCcp3N+oFBEof6rxmEm
RY56+JTh9nf/Ah5WXf+xoZh3QQabBO5q4Uxv1H+TZiakfMTIE+ZtGZ+mu7IFoKE6
egAOJJYgbT37KjNQdHhMGOpvc5rkF1bSqRAAR/mNN+sgqfCMtMfsX7rMqvdztseU
Djv+gPPAzZXhw9VqW5T1RxSDILyMij4MKL53DNaZ6CPU+AY1OKBiF9/mMfMXBDNZ
EeiBp9fQ3NN4laSEQ/YgZw==
`protect END_PROTECTED
