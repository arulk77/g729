`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCD3Px86iuHt0OnLlepITrAoek/5A6NlSi+OZr30DGA/
c0ntY0EBtCx7nWtnS8hMy7nkv+jDyreXDZIo1UQBDo9fsg7T2NQziEwUXBHjLstA
Tu/ux335nrcF24NqLCj9Xc/WQReSDkKvbnmXRC7FYGemwJEovEqr8kmbP4I8kiC5
Fxalqz3QcwkroXUxC8j7Lb8IQBjxlpfhAWZ0qWHenpjpKFBlejhmTGhRxRN1uda9
CRtQYmQkFhMOHZVZ8+mx0ymj/Vwh16V12zPiG6rk/RKrXFQx4Vxfq17eEmNY2vtS
vjr2z/OT67D5cMTQ34Ccvf/B9XJ1sSc8ENurCPqHmdBnCNcT4A5aQ4GEb5Onjoog
D3W+v0GsnsIyOMFtjjzCaZGvXK2sHm9D2YJqlt5AiMMOaontp7lB2d/bFPKlZ4SF
7dNxe6Z4jLREyL1sgCMAJ/YIHarWfbRwnSCqCXdKOrhnWKbUrr9Rn3sRdCl+iRQ6
uWnbcfstpvSvQTD/8Fduc5A0dLc8HWrXU81bVeWo2M3oUyehYeqcbzHdkn0+4aWg
xPBjrBAHlVu4+2VJl+DpN/hEmMeQ+mu0/xMyLnVfuYWe+8tmBpXkNbzN2L9qt+2E
xiqxT0mFC173Mz8/pMOnVgxo46XAuYbN3o7R09Jy6U3HHBL2DYq5TjJ317tbdktY
+RQr2rCtHiI1h6ASqzJbR2mr/bl0yU0RGDFJmAXJssfUqVJ9/BOASX9LP53Q7CPG
yXduMj/xk5anlkGWJKy6kGWkIkXRLrEWAZREKiLShVsTlcPlqrs6QG42GaAonGNY
jTTRMB8Mj4n4ns7LphA7QPF8XpWVtHDmNz2yf9kPt5Q=
`protect END_PROTECTED
