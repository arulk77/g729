`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
if7OW3neLerq5QTb0GME9wYsg9Woc4h/4jPNVLHFomcGE0TD7/eVF62khyIJN/Tq
9fRFdiuN49XRtVP1IJIf4+AO0gW2RqxbZn4QKQ4LTTqKGc61bIbat6WlxclZ7yWL
d7pdA68+1f5ZryGIma/mCMjk79zaGmhUG7kcR4/XXsj49M0DlNYkfGYx0aGqVksd
/bm3Dnjcrjf/HxSCDYE/oQfzoxkAFgdMDzzJzsRP+Qrjn02ZfR8++QKIwNVTOoaI
TwAVQ6u0vKwxXRl43qdQZZ7Y3tbHqGqBXdfHpTkFXW569LoVtB6ia+9sFwSaGzTB
3zd3Jbvic/ff8kq/kEoX8sW4Z9Ouxf+ONBTONDnF7wWVCiTxx3TbFP8zSFs6GMei
cxJBWVtK0rBMCRbz6GLaYWg+yt+7MsodhlYG+4Uoiic02kVVU4dIcybjRS4UEMDM
Il/6n2WvlKpbpz7zCMz7tLQfB2Vm8eh5ZF06NilYrSbj8usU5F7gfMpZ7NpBRUwv
OYuJcj2FtY8fIp93Ly33si8zfoV60EXFa7mMzprkzvwxoleLdVfEjpmY0pzSHP0K
r5xKINyv7DtOokV7860dN91m3mznpf9SdrI7iJ5kUOwMc6YVLelMlMYyjFgzKtIU
rSihYupEMTe9ml2KbSKnCgfSU+XI3mucmFa0VcE8c6r99+9Wzn5v5yF7HtZf1EtA
oTXBfdRKRjZumiKvdYRezG/BAJ5k4yQry3LHVyLiHQhZkxVkIhWuI4vVnMRVrxR0
lLjwcQiMv5YlqP7rBJLX9PVti3IypOXwdWwmoxszJQKFtWMhDJL+eeO9xID18bB7
MYYC+cGklkKOI+jAGnTuo5Gsu1YHQ2JMJqB/q35zZ2LerVESFe1jaN/IaHaW44IE
k0wDX0IoyvMkj8PGt7CIpfDuOCI8RNSbL2QyCcg0Xdg9FHO8CHEiBbNqkDnv8bz2
ylj5wQcSGB2Elr3YFfTYYp4kgr1FPHEligBHQbjuexVDEiB0dQW8RrrIXFXVBN5S
TVhN3mqPCTEj+XoO4OVspUR75+rnwWbxT7llQgifBQ5J1VPKQZh8ro4LSdo57iyH
3iDiCrpe/yA9BaQizWYdVjIDYLam/HoLlPeC0fN4R1+4Qz1BIludM/afLqLN6JY0
SfnuqfPmC21MjXBDUUj4Hxo3cq0SIl7JXZCwVKjGZxEQRnQat5GpLTGuXc1rc12r
nSZ71swPFAPgnvpAStFdhg5dGJCs6g+Q0bBs4GYUnR2Okt3Gt1c/7Cp8dchDt+x9
FNNBH2Zu3NbtE0fwXvbDmeBqh9yeTTuo5g/usMGxSBHzf6VVtMezsSA3kT7L9C2L
ZEm2zeepuCghw9pb8Vqv16/FsrX+xlGJpIQJRM2vG+9/aNyWlcivT4k/F5j1ypL7
h2gFjaTh0iOqVo9LEsL3EmLNJrtnR92KGEEH0WzRhQDyyeEFuGFjbdQpp27PHYpl
vGOk9ze5v58FmAoCcBQa0lq4BsZ90Ma5TU6LiDG7ELZlUppj7f8tS3XlS8OXY7nm
y1JIR+J/yfRst/yIxvx6/MIgFqB5pS0L/7TuwSt2MW+nda+nsopVEfrStWeGj2qX
S9iBbFKbSmmIGpzhRzH+qL7zeJ3j5CnLmmxhjnmf+oLRdliiymNzIIOyYOuMikol
wg0ujnZM/3RIRJ6MqluZnmbTdfDlpEnxeJ7wxLM6j/krVGHWSmlO05lrxvEkWSW9
Fj+46MaXMFoeokHzdVbiI50Iwj4IckAs6RJQpnZ4v9rx8r3tVYeOkbryECIZFrpu
nZGX7+j2F1zriqCpqKODbj+tRXWM1bQ8M3Y0E+EGLWGYO1YqNQuCSrKQKRTVAT+R
IuzBF67v9REarWAN5fWiMG+a6JL2sc8r7M0ljvpqFCGbylDIHRsD5qqZvUGws8za
e7FZsPtpFiFIvRZqIDt3gPHVm1NCcVC8zYiDgcPQlz5eoDJMO8Fm9ZixOJ4B+Pwk
/YUdh4imUmRKjzb25meweDhmEaS3tsMOuXeO58Mcr1k6ZPKOeAHpFXiS16O9rNTu
olZ7M0usAwqlU0QToYLmTqlowIjXMgceyHZz5E+dw+Co4XoePyx4d2zynRjzOEhY
2zEQ5MwPMiunS8juMnnumIL2z9bQwgNpzrGhKtu2g8Zx/5jITzPGy4/fsFQgcMI7
DLCfkAI8IxscZ+W1uW3CVrw0Py1ysGGNzEczSZUizv9BYRROrZfgRh+kAE9ZAqeO
FUlERb5No22ML8lXgBVwjTx3c5okdGEL9SJobsWA2xXqDehoLOppKayx2EXmFXYw
zxJHzm4lHua4Sv4OJ3r3pgtZCEsFHCoIJzf8JmUPMnSQoS431STb4A/kWBOVu+Pn
omu+48dvK0LBDGALu1KcCwQCMYKXlfKwQOaOmxKbRRYzCUUwY1icEXMn7CbiVs7X
3Bp8VPxEiOJab09+16jLI62CQ1f54iryA9QtxpqOQGqs7t18LkqQ2pRNUlTHITZZ
BS9fpXkxZWqSB0iq/maZad8GL6IQjhJF5FIbpgpLKIzNVYwXas5GNADxDiqrktQR
a69xefcql1GJ5rvbJqiqxyeCfD7aDNuALOTEhucozka3kjvELkbJWp4SYvPafhU2
N1IZi/IL+rY2d1+DI9uPv7jRrcm68/hHD7zJhWLM11rljecGP6V2xbERRYfOi+jl
E4vi4/UwQRDg05RdqPTZSWrkxxzTJ36+6Cz1TWqbMkMxjleyZwaCMn//zl2mnBpl
PSdswGJCeZzszdpoo1KSibrl79HXMNGiQVYShNrHHQAqQRnsIzmdlXo9jSLr/osB
10GhnFOZ5HsmRKK+ucNA7zvo0xyDBIIobsJmw+BiYoZ88IGI92jo5tVdw/iGfWKC
DbVsgm00b5BCMvNQO3yR72MvGzkkrlXwC+DpqX38wojarAEVyPpqTr3SqrLW1bpR
eHfZhGGUb8ZpTRNDPdsJXeHKAhJhdlztZQr+QPB3FNYtMi683GxTRox5QBU4ksj2
1uKEqY79o3m8esaYzMdKukFRC5Yuuv9Ag/lv1tWP3XC8IGcdB7mnGzqWdTZG87rZ
87n4bhbvFYMmgraaAyoTWjbBfVbI4zz7Sx8a2QroZ8Xp4733icuwf+7s+ydWm3nB
npd6MhkUAohF1C0Faqx4X+H8aiycSyWSUK4RreBeLvOyYp5WEzh0M29hFvZFvQW2
MwuO5GX8Xiwa/7EltFO5/AEU4m8XclU4b1wHV4dhtH45QTZFUXWDuV0PHJU6tKr3
4q25UoS1dxm3fUtLoK+AccnoVlPF80E5tBdauF/lQfRupi0Qk+1+gmZwFSkLPLos
jLemPGgAvqdPVyFxPJlotOWfqqi7O5LCleHpYghlwP9fkyxbzDx8jentq/pn7kZD
Z/SfIUTNkq1OuSEu+VfNDIgRZiDoXSSHX6QY550KmjBUwq2S96EVWhy1yMO0N5lx
FjdXDEON0Hx1mqtp1umKG7/FZhk/cV/hcEsD45W1aoSDi0S38CCIDQXU6QVkDqyz
iYT2rnOE+UkLAgmYs29MX9T49X/nvI5hMyWnvpwmt/s5cmDZMOwSC5f1ZkrNtGb8
nvHyygW3sBXv7Tnx/tzZGIh5KfY5VINeWtIYXgdnS06KkBDFUfdMjcXR0+HVPwzz
5fVt0UEaKzfJC/oh+UldLy1+j7ugHFaYAe3hfbL9aUWajLHuKbYZlp7MbL3T/kfE
VgcMwfEpwI+5lkEGOGiOFWpu40N7yfOI7oHbozNBYiOLYH2NbTrk5HxaeMr9fmCv
dpW4lbgHX+1h/qBWmil4JWsub31V4yHeEHOZmrlebL0vrsqaBfVzyh73f+w2XdCx
9yNFgqlnTjD4X9qEkmfLaLcXmWWH1Gb+JwvFz1hT/EcjJdJKOawjb92GNOkoeaep
1ibT6yfPmVgD4kLKjtZbvmjAhTjjMMC3dMrG55re+FOXLqYBPmeq6Y2YRCEi2oI5
Y1pqtyGBGL0/z8C0WQw3w6kRCnZEt2dg+5etpRPGncpLMLC6mRmzwm1V4vOiDV5K
mEo0zyj/VhwdtE3mLhAn8OV69YoZhVaGe7G8y0D/gO4fy0Rym96ZD8/kLV6kPYxg
VuB3CFqOOh3doC6HpOoRhe+VF0eN4v1emc2CYs3P6NnNoiLI5plvYyArd7SPWCUZ
IkqWD0KoEY5/sYqFlXiYX9YV4WOry2uF3zVYCwHqTnpc6x9xezYDO4PaXy6qqt/a
2UQJp1TRmTXm+/LVwdTt2t32UFhIAypG1JoZvqCkmgxcFtOVo9OSRH62Vw4LqlmJ
lCwo4SSFt4mIBe4WzJYeokz4jJrm7W0jOSndQFP85/DtPc+2RfxmOS+MlU9JD0af
pp50oS3bgSt6eQzo4+J6EPIFNoSGRgnznYIMSSjjwbsa1LBxRumYA0hYF0/ocuse
/Xu+wNsMcCQshFGPAIisUAFwOnEhrBDIhGYsuUYZ4OWWVyzcMeXlvRO6p2coXGce
5ayQfCGuUkwdb+wGZwB7jx4YyjIMpxNH2c/WgaWmSH5zCkX45fmH1C6T702Uzj5l
V3KOLgGfPQ4ohaeQ1QMc40V02IjOl0Oiqo+b+DiNeiByatLzPRI5W9Iww73Lh3qY
RHF1XmWToka5Y+IAjkSVLrdUzlA4zAHy5LaEYFidodRh4fJgEIcQfMwCEu9qmvQE
7Rr+Gaii6PW+2Vl1/mBePRHKwPnfzn+w3337jpLKvm0iK+zTksCFQYtbgbBQgAJN
nDY/3JOZ5mXaDN54DqoQ5aJbCfvHVzw1zjVqWNLYg8HtHZ+4cbUU7/jRnpFnbTlx
vdIMFDz8RVE+n2VpNU548YiTPwFvIM2FYKUBzFkJV+Pl4cwrAUu8YHnR4OwNUhZX
NPuBuTgqlqVyf3DIJFb9Ird30gmqkWR9BaXPf5Fm49Bry4mPUlRybk6k99Ghn9z6
+AIlmSTtLeEbjse1jEdg6h8IaFNRkOSJXxjIP9MgREDzUA/6kEeoG5p/0a4QwFHY
gDIVZtMsFoTVmaxPyPHLUvXAzNlBwMlJm4YP51qzrQc7fPHeS+YJT0xeRTfaTIaW
2Yny5ED5NYUG/NRFOXbYdQlBgrPACcANqmeADViOjUOziF9/+m9/IbRTs6ly6i3E
hSSfAGLoF2LuaBXe2S5ck4UNYoEFQ/BxJfV0PZuZY08i8t4Sb8+526+Zd9sBqmjK
1R/hfqvi0hGiUiizC9FqJKkmUMLnGRBOFXB29HVem1KspXBS2bUBVm62d3yoq0GG
/oWcu43YpF+mgpTR3PodXZ5lJI0Q3cM3SAt33pyYYns809/jsMLtrKmRFXkdn1Vd
O4L12sC8kslTsgSTLLBhZi/hlIKbQIoVFY5KQVbMwD8upy4jYaS80Rs9TPtqkxlB
k2G8x6jQIv/Y7FRRSY/g9rsZsC5zUrZ1WriZLgM5enHzQAK2eP7g4/bH9nt5xyg1
aNtnJUWPIlSTP1F1ENvuqCotHG2/8HQBNHyeLt+v1KEP+QuxPiRUaWOssUMLZW/P
6j7EZp6YUMElbLRJ8mTjBqzh725AIuxhZQdTqwOG7mFysyb7Q7DoecZbmJTZ3v5Z
0UqjIZ0rX8w/Qlzs8JXEjUJgx3vIgCm9LEW4Tc6oGHZRWPCcIl7IWFwiCwH/QsPw
tIfaZDGeHxg7HKexXi+b6bkDuewBH8Rr1iScGh7MzIQ3gzH+Ugv0Hkoa6/Br1sfA
dNY0KgEiPiXB0zbrBUjkvehubfkSCRgjIJrgGyt6Hkt92ok03M3sWcVng3CgozYL
nNTfSF3tA1RN8MwH0iiu+FPksppMSh35HKSfsvu9V9ZXPL8Fc+vOALqKssJgVwxo
TQXS6gd0GuOT9YMbyxsJ7Y4nYrgDJynpIX+aKn9QGaGPeCM/6LnzOW3IEulJIHpi
KPm8esowJsg6yHhN6GS33+2uoJ3OCwHEA+CpBf37LeP9O+kwhlyAyDN5hvaFbKFw
FiSVoHJJ8gez+htM6mPSRJ33F/g53s249xOJWUT8yfuxTOVNU0ENQ2mD7KMJCQB5
k7UlgPqkq+UiYGxr6vCrdZhuPU7b3ZLcRujE6SkAfH+93X0bKsmuG1O/D4fUij9E
i61t0pTUquqG0Oqg8T7cLsGdaa3/yRZpMbHbdLL/1abKhoMdUZNk+9XyIcGJo/2+
y0Fb31j6qxUoi89VnfKNjKL9LMlVRkrAW85QZK5nbGuwrStPdrFXXzJK+44egz+6
4tyBCPsLsB/IHISe6WXJkd4dNaQh9vgLCkBoCuvBL0oifOeata1sPPHp1vcb/A7r
r0NiuEP6FryUFcLME2WR86mFdwzJBwS9/Bc9ybMmATFkY5Cu6OKXs0Cl/3fW38d0
Wl0BrDGaKWpFzOb6mtScJ6w+LeR/kVA9l41c11GZoWCrdsszVhlY06ZaLxa9I+SG
n+fKBI3pGxMU0ySpiVb4/Bjs3410XWr41qvhUn7wXJbVebF7ZMpJwuRWpuecJN9U
B3G7ORXTkBLpuZJ9JdeELJ+uMAmhS7N8hMZR2u21unfSKGMys6BZbOxl96+DBOVf
W1alfGkfAfCNxm1SA+y2ILq5PyZ3/vuU9VzsyLuOT6y90fJ1JcNhwYWb5cPfWJdk
e4IjYjmxZMygTFwSLi7qtyDqdzhGzk3MC2uUZpuWMZRb8pdtVYrgp6ZFDbp9mPQO
eRW9WSJTUPHKlyOf5ug+Yw8Dx0UzQoZtEWiV6i0jx7C9ZZOdkmvJsUDoUKYeo/Ei
r2/7NqtCsiPD80X0yRVnGFeLC6ESmRntOHgTgOHLB0tmWZCOT5GI2NEsZpTah+Cm
QmxF5t3V7plLsdgJ2vubKuK/SazsVv/SPQ1L9LySBYjuO/CH4OMt2HzFJE3/BCQQ
PhpravMD0HvDKxlRrkxN9utgiup7b8sfNpKs2dG743VTfJ5gWcQE9hvevMSdU5FL
0n2A7eV6vBhiZ0YLQsqfVqql+l3+XNb9w9SVjE+JyIM2Y0eGddzHlG1B6P9yVojd
zkfuB94r5wgvGl/YMSCfPuoyyy6IuHzJAdhFpOqmunv21agNMtTFBeOjHRn5Jr/k
EOHFqdkA95pN/APKItGQp1+NuhwNRWrWphBUHWnISMj9vtclhyAqyJaYcZscBr18
xTza7Bo5rYd89pgZcqo75Sa2YC0QFcIsD+KgH7OZGC73hmT4KwheH5kEMfJKsTYb
yqvEBa/pmYjDGpjATASbr8t+U/BBVT9HDGcTSyS+M452eSj3cCYKR1U/YSsDAWBD
zTAMdvKn+M8NZBkizDHqgntTwNxZzrdcOOkiec1OKHYV4I7EuCMyK6KGovUDsTjD
7kuLdSRvAPDTAP06dORZ9eSIj91qL9F34HSAlQLs6d+bwR4CiFMHXFUPTk2u6aep
p9CnzrE0loA309OgQCFaxUsn0/9fHTx8oB6Ry35xxmydWK5GkiLCBDc5DoysppTy
nWKzGX40nuNVcv9aoffXCf20V9NU/GSUzGPZNAyxihnpkvXSf62WvWyS754jc6ZP
58rO7oBNxYC7dMTb2CqWhcMv2cr/ACV2csFjpopSVsccCzUqpWKs/p1yij8a1zWI
IBeNBgVkeJkHUyeOVFxcUa5IR2FwMi82qygMYCJc6BzXCbVtLyMgdfnpPZ5kya/Y
MeNZp4UlUsUu19nKLv4YtGPGofCQ0LKQosAEW11Vs+ibncZqS4OlywwDc8SxFRO0
/TJNJvecfhG4vkXl3r2szBPieVhuDlYIa2Sw0i+FLCoOQuUrHEbGkHLAIV4CEBh2
Z2gq4ti9LlkkD9yPQT53oV33qysbH4FhCMJ8FCrSjUqWAsX1tTBw3NxbJkWYC1L7
s1GwEpIHcv/+DzmQkFcdp8h2XSHe9TtVU1HvuAc/TcBHKJNr1s9wlwXVMLMaBArZ
k80SLZVsxBsUWctwr6ESoSHIVF97agd+CfyzPLp2kgQWY3LsAyVVd6xcUDqJ2ZOP
cZY5JOjOgroKdTtcGroYGvjq3W5+2BSnvLEx256yI+h6HqgovdHjIus/ft9Vn5pi
6m9q0JcJSMqQo4OW1zufYu+Om4nzyP0Fk8UzrBiKQoaHJfFM+xOwlkew60sqgp0R
n86xB/GQxXIun1O9w5o0jr5n6pI3hHSgL3IxaBnEuvGK47Ftr7kRXCjhlfzNCZFh
t+GcawWHQ3iYd/2loT51FHnk+4rwdzjoWk+EOWw6p7dfObgnxEl4p5Dh0nptqfb9
PnQ8gQrlYC1QMxbnv4dhfIFA9rpt2tEABJW5yUtRhi+ic+rd/KPPFsc6TYYIxaGe
jkkE1W5hSJcd8w2mNFHreH1kEgfMs5VuFNQ8oEAd0FVRGaEdY8mbTkQVohagTyXY
jPbBnm0e9PgGBQbvRJuYSIN+aSCwgRgTsVpqIfwWdaQ4FjLJiNi02lmBQ0m5CtOZ
51sxbIK4+/9sQ5lj8K26OlVJpwHTMHDOapgNIfxdv/NsLZGora0ja3hyC+wLTtRz
R7n3MEh5uF2Cz2T0eFKW1UX3efbf34CUVkpZQb7QoArxoia5z1l9Fa2OwGvzC0TA
HR4F0FeWtHXgEDKcrW1ZxE7E54N8PPf6KGA1B9ZqqWQYtnKYluEJGccE0KaqI5LI
WI6ubaZp207dR0rJaO1HXgFRMlbAHiZSLl1U7XCkFsR/YgXB1zTHabiyjYh/T6y8
vY+8o+X7ZjVnTv7dbtyy6gZhMvMmDi/GKhTNCb9J1p2mjSVsNRSDsKr1gYjUw2wz
eTS5LPMIrHSKy9cQnC5N9Yyh536J4ej4MP/aVc1fgWtyrEi/9gdEW9jWprkHg/e2
CT4WziiNIIlU4H3PAtNngxCCCIkqk+W0rJnGhUJ15bzF8HLVtstwILdtfJyYfaNY
dzq7Jy7WzZJOqWOsH7zvZD2O5Y/6XEQcmJjrS1KkXuRsh0jF/JIT6qD8DAiwFvRM
md31hJQug04hhCzWLLgCwA9scAYBNc9An7f87yWRctltkh9sEquFLbNsaP+qHGD9
TQt+k3zu3bulak3M+peu6qLoAhzG7RuUCZUHIKnHC0M5KzDSm7p02oDoc5owgDhF
iPfFU95+12ZcLGvDRm1Ksb5QqzIsYryVeVV614FLFodOYkxvjIT3H3pdcZ3udymo
z0N6dnC1XEqwf5lP3/VV1OUvhbJjqYuBsqVjdgFNgHQ6npNa3T6lEGef2wjLUsZ1
U5X27QSNA6bfHUonT6Kaxe5B2Wy/foOtVvk56BtBeooXiIJr7Bl3iUHB0l+J37cA
Qb07qFdiIPySF1PVIhYa+7FXhQgAeWrsDuf1XSx/IdODj7WeMhTLEb2qO6aWpuRl
AT2Komyr8B3PLVOxqOdmFgpQ9HOWtpbjB1kaRAJ7jxfjEs4I/1I/FUak6yDWhpns
qxBF9TCWdPRLykW9l1Y4cY6WZIMdtNWgMbxr+x5RP3h7bjx7DsBqWmIv3jslXCId
wL3E6SPrCk+qR/mewconX9HOa7nsJ5FJOLMPao+CINVbEiHlLDCjY5Xi3HIq1BU7
uygqXjU/ecUQj0GBvC2M6xJDab5y0qsX8S+sjcmdLFEOKnJQaGC3/ur3HjV89hJq
XvD/hOH6xPux9L88nlUhFGMQh7sf0J1yXt7r4lszWZ7ejmW31B8hk+303Jv0pE51
OTd0riNXoSVuhTYPMLXZdOlcafB80WPIVNR6FAbFM7LzxpWNf/ojFwxT0RSAXnjQ
HIyTIboHUgOtkSOlsyRpSHGQER8fqMaR4d2EoLp7sRbxcaiPWaljM1OpqDxhOUAq
6yWkf+x7ksmV+WPoLR/W7tBRffJ82R0C6YAjhFj1006tB5mclsvgkD2/MouJAGVE
IVJJ51czM5qaZtPbcS5XdekEoradxEiQ28m/EefGKIQTxRG6pChqim4CT4JYtMcb
7GEQD7WaPesiApJJFYhIQeMafcX1K5OVkm+EaybPJyLg7IkxEV8Koo3y8cb2Uzkb
CoWeuk+qTc5gPfWamufXTetXNVjb2hRF2w4WKG+DPASm5klUXicXIdcFyJ60ahbq
JtvmB0h0gEzEgjIjVDhWieysWGTEoNL60Y57+GYxNRwiTDj4PH0eBzgh70a2x3Ot
yyOJgIElN2GeYJ0ODRPRtB1qwtZclWH4ptr7NnrlEwXX9NPhP2uNXVPYXYC91haL
o6gDfTwCNTsKlGhiCxlEDxkU3kS7OfVprWyHDi3ln7kHDrCJ3WdpkArJ/43odzfk
Bl7cFRzGFIIrh5ymeeN0a1VPcwJ7rOd8jVbvK3Sop/h51oyEPIcxCBOwqbKM20Ue
JsBi/vN3Xm4GVqaGPUm5wny65iUcHh2FbZfCbHipVT6xIqOpV2RHsatmY608MKjM
YEgAB1X6f/9NZZOXOXpwOpbXk7HTxrKIbD3ywTLkUXyrHZKp44Wkgp7HQnpc4VLe
6FO1hdpAwBuykOkf1PVcALmo3ACz3KlyO5vYEB6p8ACAZTPQ+hB79DB5rTCVKpn5
StwbNMeIoqV3Qro5yxnnM8q6gvNEwB7HRA1fRMxWu5v01bzHhct/MiFBYv1jHc8A
yOadYLE3DC2lt6hsElLe/O3GXcbaxal+CYWhaI0+bRlBLqKOB/M1l1Kwcinawm8+
1NII4YfsOdTmxyCxIXHxyVI7XuVSQq2z/FyhUmngT86z4qKZYhIdLCtSIolcUHvr
Zy7Ag36gX7OvqFFOt3y6Ea/y8j4rQva3AMj46SXyk3W5Nk79CzgTAP1K6QeNojvR
7rV1zMuuZpU8Rvl9GRJCvIX5NyMpEMCgmNSdtmoag33VBfHwAQ0gU05tUV5IgoPo
Af2pnY4+BEnmzV+2UCJAp68DhTpxzgNN9obEjn8A9rUwa7x6oLUwrzGKc9PmC6/O
AyA3G+5jO/IjQ3HAC6auHw8Mb53pxQFIC4iCSug+/ciTvVq/eAnovnEXOOM+kY/C
yL3ORji1uFlgqA3zWNm8aRAdxyN2oA6CkUPXjk2et26tF1O+TMZbqMu0K2uya7KJ
eFI8/aWWZAVHr3N0t90W1NNUEe/9V5aD8FrXSxVfv2Vg2ikYAKla7Tn+Bf/OgK7j
dkzOxDrtZLzpwJeEnIFAekeSy3zwSru7y8e8Y1HHgg529b/uGoa30eWw119SjGJh
lrKIbu8tSaTfZeEbUvVqQrSbQxTlvSMxhV4q3pnM6jVNePnEGxNQhH0Y1t9xG0ic
bGnZROXSxIotwEQaDs1bT4y4P6huG/6NFA9EZct/KMH1IP+NAgpiI2Cv706698aP
/oLlZ8H5sLEPHLI200UcZ4+8cp26iwCTublcr6ezFTlV9zz2Vpv7T2YuQWWt9XHQ
zyvkps4ZmuASFGNXw/hlTMUHsz8ZXnw76zXcaoAUJ4nZ5xK239FcZRKrliFePOQn
DRaokdbox8+KdQLW+GXKnP/4/cs9Hh0u1t9pmpb4ybULvwqtHxHoexGBZ3HaiFAD
7/1Blld2wnYUMRZP+VMzOsIXr+uUQ3gSGZ8Vf/GUJuPh0qmZOPq3QvVnrWb2t+ZY
mVz1kYTwtX/RVtmRSnkNz2rwIPk5PW/BLIhMn8s4yqWfpOE62AFy8aSMHYMnhUU6
McSJ0s0i1KYklOV0fH8kXBksg0Mpy0sdHvquEarGzUeQxB4JRa15WTsOmZc2+jxC
JL/e8YUR+1yZ7HWD7KHbJKHc9SknV2AL0El5hQI3/Q1yzFfX1Wv/lelAO/trLESh
UbQqxFossZ1MeYbU4b2aG3MzoPvAWnPIbhXV5MVslTTtMNhit8lWo2mL6bSvZYvS
fKDtY6pJAZhKt74jrt+bS8iILQMbjNa6wvZQT1YnES1vsEsv2W7QxMYLGoBuVQfy
tpOrTDKtqzf4NIdDZQh1SXsthwIGgi6TUDXP6s0gGvDHAj/zLww0vQwq59zRpGyo
iLG7e0X4hcadlfDC+sHXIbvWD6s/pVSbYZqI/JM17Tyz7yXoJcWuvzRcR0UoiXLv
0BD933/Wzz/d1xt6FeTaLCug9R1dtFFrBPA/7GkXxcstgK7B6y/si8xcrNWRdYaV
WhS048crB2Au7Vee9hqxIgmlBLgvsIOWhBbgIg2JHKhHC5R/IBEGuX5MlOAotCJf
FO6vNQJEeBwd+B55SU3u+MI7Wc5fIx51hmQJXLPwLe3PFfS4yEd4r3lZqT013EKh
uyCdd40Gh/LrUMrdVLBMbQzCnfRQapK0ie1cGxRhkadZsRZtpe0H/MvqjfZ7DUCN
gntuOI5tLSxvNk3Kswm4vr+dz5ZHSWPDGjPlcoQZzPXvTI75d7E4SpwKl5qLt731
AmqMxyWXJG5+Gqb9iJnnBc5AIqmJEc9xViiiZwSXJ5Mt2daS8qWa0OV7ms0Z43CE
etXQdVTjmPqPkQt3lBo7MpBwlg/Ah2Y54zSS9d+RxwCbZR9Ch3qPPAZGn0h9KY+G
WJ7llsKZzXhR2McrYwPAWFScpXu7zZpu5lb/5UMKmpKSS3RqAkYWoftJRTqB6z0U
D3lIuvhV8ASNw1zksCRjerBKwwpNfdYl6bCUpAq+YX/8ejYaH1SXQ7W0YvtujQUM
U95SOnxTYGPIhe8arvlQF1yTUaN7yGX20j88Pxhsx1ouwcKpI0I5Paste06ZltGo
EsWZDkOqSB5Lwu3FZr0rJ64YQJxh6E3HKceMHp6QbfJKAVKKl3DkcMPV48UcAeb7
luTRBzfkovgfYeJtGxwVDsSIiQVeKIg+BKetGitSCS9Rph+7D1m3L68E+GOazg6f
UMBu/kmocNfe68ooWtsVKF4vBGvBy8sx5jQf7KShyp3cAX5o6N+FPOmbsYvD5JWj
sFjPjscQDCD/l4v/H8PwEO+j7X6TMAWfOFrbjcghxpnxCPhHt6I6bkTqjJSVddTa
J2F1L5L6M9yY+gLCHgcGZioF1XBvSGsJnFPR6JPEYAE7nJvHTjzRbQNj3TyFcBDP
3DV+wmvQspi9fWX4Ai/SbNMnj34JM9siojtgseTfTxo+k+2okIbFHi7WPr5EB8UM
d/r0qJOe3Xuje3F/MbSeb/PFdAUUz8MkpFyPjhb8Bav6+dhoZuL7um/Qb5LZjxBR
jhLcAohc7zR24y9MJsEFMrHad2+Q1LfLC1uNPZCLaTZVik9z/Zd/5SwuyQqg5jOm
52XFSMbbw4ebe3vNIdWtdmLe/gZZXUNNBVDVa64DuQPDjtVSfYqXWiOWS7xPBINB
2P9nxV86MxT4IQm0lhYZjAIC4X8/GJBARy5WZG6j6/d7HOAe740N3vB6VhBizqwQ
S1zJhociyiuF5+d81L3puqD7y9X0zz6K9d6PK5ow11CFgjPKj4bfsT2NTbycnr60
m3JR/KEOSC3ijCV7yFm8kPcA75/RajMtEM847XFjEaiyurULzSXT/gzW59/EIVuc
defG8CEjA+vPUfkROR2pQDblAI+QotMA17Wbu5Q6/649id06cKSifGe1BHGYBYKB
cBxhFLvia+D8u5lVPfm3IPe5iLTvDxYnkZQF7ZD3KhKylIQro0JAKrj4iu+b13c6
vT0/IyXWC6ra4ttsg9XVOwgj8H/OhsqBLv92AYz09lgf/IG371CD1xixdeFoJqt9
ehY/+Ty1iEpb1hVar1zP0ZPXPzkueUhQBE+xplKH+wyb3HT/8mdk9AL8MwtKKXT0
`protect END_PROTECTED
