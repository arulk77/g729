`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
po6OxryX1u5J1lEIndyX8AsTQjtk3ZPbuSH64NH2Tp8SpCjvh9aD7CVh3lApNPPu
vAlQcBx0RuRetd4xSwpS983ZjvAp2qVR6Mvo5qBdF2mzsYM3WjTsWkYtV4Z0uWdX
SpVBlhhwflQCZMBaIK+Csi1MVJwFY7CxKZuPYrKranVf3rjl3bhVKUoMJo+lbhgr
D08kpIFZwIppk05EWIt77UqdXVIiYL699vBLC69uznRb7xmTMIjTV8kLHf8tToTW
wYLyn0DtRLoSdpmFI3HtOfnAwqOEb4Rsi1WPST7rSj8=
`protect END_PROTECTED
