`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL83TFqqM5JZf1WEt2arccWJfuG07EEpTjuJGeBLbhRAOK
IC3r6JYKCRwxTnoApNjDmDKCxGCODEN6B8CJv52oxl+kiG4qUkn2Lf1XubJMEPzB
1H16SPXzdhxNMIqT0t95E7BueVSChfL742RUW11mNgz4EGHZyePlw4B3fngxacLu
aXb+7oHHDObr8muIhtf9T7SVI/JEO1remmsK5PweD/r2Qtqofwkj+/vDfVYPFz9O
2r8wen+nonFOn9yWSysAqx3v3t5CZkb1xei7F3nnSZMNSOi9HwEz1sK8fOwPhD5w
5AXY/1ccKv/mIB1dlv42fZk5gVABf8b18y+IZARJ24AiMtf7BZ1NLfjAgSb8ScbA
lgEgXHJvPHz7ffIPppmIlaSgrW0oOKCDsLCm3USvl+0y44dmcmmBJaWtoTvq8AC8
nbGNzkT7HfSz1x9Rr4ddEkURCfkej6CWTMI6ZTXyzGUbyu4kU8eSVTIr1xJFjyQO
bRHYdDXYHQ7aPzrN/PvJuqo4TRM2Vv3nddW4rkdU7Stfy3MaD0vjecgDcvVqAiPK
UTRE2zZDm910Qnvkwfla48XnD8EhNYD9TbYIk6ILIOOhTWfza6bOdW9DgLti345U
EgUKyPQlT8i6I3jl8RRaLWeubArVxkIqr5EXsskeLE/u30CZLn6e9GzBsaU/eF2J
S3uxmn9Iq+RGAuFT4zYcMeRlcK/OAgUcgAZIFanFIdgCj/CCRdTl7JFqcQnnKkvA
TaPna1VDHPmP+/C0N9PJrx3oemYYJqtTzUpwAksVSLwZ9lQpuyzI63fcZ1hU40xw
AqROAMbID8EZys6MhOAdaCGKfSkXhn8PdlRX1S5YjC49pAUWdJg4lH0GDgis0nqh
Ax/3g047iTp/jq587w/RXEzv1i6fzPc8e9n9fO2QeQBCVklhr3UXQe3Ke9+0aHgp
UgLWLDo8rUzO+qIRQskc3wOtaZMzN9aP0BsXuL+nNL5mcSx8E6yKLBOx4Xvz7Fq7
qfoVxXeDGsUfSCOXFzm1Dthuz37XGe7C3lJTmpfOq9FyVVR5HFotQTP+GHYC6tjP
+tqWNBlkPZR1fFFcAW04vUqD7vWLdar6R+nAdmIu1bJSZiGLXJGF+ueijwkywq2q
NZo+OloCnM/XfPwR0bCXbYN38IZWZKWFhxkoNmkn3vYOVYP6GLXqnEaX4QVJtWcu
BVODEXDkZh4kzjfBdaBL6Ep17ar53aR+PekeL+IV1pgJVa47wFkFqmoTcsth3VmV
EkCiVf67iQ1WjJkCTcOTy4ckoneXOv+NzDOGdU6/ktdgpQoTC0jUfCeQo/PZcvoa
8FY3Mo4z06kAR7lQPJPddKwxDUANbRZhzQTPgxi+/sg=
`protect END_PROTECTED
