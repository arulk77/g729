`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
C8ONwIUaisBoAfHH3O4wq8/6bSuUoXlNcl1IvUkc5rJdAPwSc91T08IGsqVxddOz
J07W8hUO67FdmkfdDcLQkdfwWK02A4t9FShb1W/DXhg4GMIPcN3IoxER4VuvmlwM
c/0tCZFQYC0oSTsy+B+kiWDe7ZtGGFpEUYN1qm/GCxSdyfRThIxPzwaB3Mm73+h7
afpYvh2qSBExibXfRcEuEnoMbOLaW8xuAj3GGjyndPZyHsq04+U/SAtPeGhiTDhq
cZnM7FRZWitA+qtAQWv5ANdBkavR3qlDI52gkkQbdp6ZDDUKi/J4V/OFI6XxQs0L
yW5BYa1c42aOW5amL0ISpqNJXW95n7Pb9f1ww8Mlm4Kg1JBmjdV1cUMrsHM4ymO9
omqZS6WBhvMBP3vku1l0es/qTwLKqLgNJNMRV0VddQADODcHSzN+YdVMjyKZaqQ8
QOoy0Ek0iVxN7WB3NhTNqhZZ9g/G/TOhjW87Lcm4+3dOcNdxndUWyztyZSrL3oRn
/fIEJxCTZH+l9cQ96navbd9rxR5Tn/vOuFcIJt1g3Z27U8Af3jJYjGTzHKcENH/a
t/jcaP7TXaRPd0tOL5F80d3cRy3Rb6FFVaelILWVrdeVAvvTXM71A/tV3N95knTW
zwa/frCbod6QoPdCJnK154FuzPIl7jXZgjtJ/PpmIRv+ILQ5iDNb3tkDGL3PYu6I
4FeOStm0iUprp3WD+OzE0gk2rqFzcRbSIOxkT6u1izQ/y+TgfnGa6a+utdIkgGNn
BAajA/aaGadQX4e2aVMgGC+icj+W8pWI1thBr51fc/f/iJGLhHlc+GFfXi6vDTYj
6AyV5ktzWXgQWFENd5hQEX+jC+f1WJvAovFNeOiVJqoeuWPXX+KEx4rsHjm5ZoGe
061rBj8sik8SBXEmixfalueO4PvhmHLc4P2S6D0Xb2vvTpmNOne1BcL3aVqt4GXO
UMqc1p0+L2Zfw5BlDfsfBOUntes4fod+KZDBdR9kESTwinFKH40nbK5t8r4PTQi/
weaAa1i8dpt7dOYy7vqVUQ==
`protect END_PROTECTED
