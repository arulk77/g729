`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJAebOwVab7mep7SckUIZPkDcPw8Ec/LtkEWlun7cqq7
nph1frpW8l8RN1AucyxLecIOcCf1e5ZA+z7aFD1EwejPlV9QM/4EZtfPnLtKcUao
xsHgfTRZSoYrsIMjdvhl+8EoMh9Trw1Zf9w0ybkm6wMIfZ6VQfOciU3frbc5xnQu
K/TpSrDy4zRiU/G0jPUJ+r1PWURGE3ICBwfihTK+GNc8nbD+T5VUgjpmmFymTu80
sMhnYrkCRIWTBLkwtl2ibqv398MYd+g8AV698S05GIw1ZJ9HD4jWPocr9vw6Phul
ZpV/Hq4zvqAgev2sUjJkYlWV3F+lPdoj1nYWWbaqxE1Zcg6tbjSsDLGjG6jgyEbd
u+NKKzTuLheuIpBtRJDd6FYGxDRY3/dHt1e4oKRf0dn0SRmahTBff26l2bWb8iZ0
E2q2f2ZbS+97vzpaD/9tTySYRq/LOh9u7lMcbPTU4G/RjMMwocDwLnlhR9+gWxed
5KVHyGTOROjkytjxQ4or9JfRNC0zs6nnxqx4XNPlmO4cHdWFkmN/H1JQRwL/vf1w
LFZ2sTVJE9+huxoDkrvQOG7mo8oEUI+m6BN7ISbmUo9+CKp0Z6wFLnNRuw517bif
`protect END_PROTECTED
