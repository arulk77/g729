`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveC9GcCkGJNAvoyMfd7Ho5RN1FWB3+sh+ay/SxS/7jeuy
ggiUORnjRAb5EMEMVLsQ1rrfu6nV3jE0+qNHyYD2ysxKoAR8UmDFGuwPURaS238S
joouCYJYYDi4EXYIdfwlTxGwwOwZ+7Iz5GDKK7HG7l1JFHDkr38tGZHULOzINw6H
oHi5bgx0AZsL7qAotPY/JwXV6rLw7qDhgD1YhAwTNXk5bhuBE5B6sqW1WzTvSgFV
nwdF+dVxXLRHkvmJoDm9mg==
`protect END_PROTECTED
