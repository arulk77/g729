`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ9ZdHsyuyl63dijN5w2AR/M3gPl+G57aGgBl+LdP7U4
/QdgdgCg4ylIS2dHFKojl7lwyTl0PI4a/rcmY35T0dUw/4lQ9CJ5gz9aVzhXcBiv
DLkcnDYdrMWIqjH5thnaoRK1wOypxbA95/5cNXN/ISxmwi8px5vIkDrw/UxEFDy/
p2jFwiFRWaQid6YmaII+A4tlbx32Vu0RymkR4TARZ8FZO568OHscKZI1G0zr7sLC
yZUFAzLBt0zj3ISXc3M7odxjTxIpriZV+bh05PMM8GbgRTA8t3WrSxeUMnk1ntET
v5R6UkFzlNFdMUcRDvBTvN8hAiqyuQwL4xJX+MFzHpFjlXJDKx3S/ebHRWaedcTG
p+ePOHFaQx0WN+/rSM8xlNHicJav8HoHx1GArTmSR25hkuoFJIpuB/veBQKnFcNL
XQ2YBynTW4Nd1jffYnidmaNunvCDGEdjvEHXNzkCMRiDADyFRKqEUJXsqcCqJI9O
dSo2gHHApRqRtgH/OX0xFA==
`protect END_PROTECTED
