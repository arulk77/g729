`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mlFBzCyNIVABC0bhYTMiK8QJT7/xCoPbXh/nPbMzZgchZpDECnUPC+9i8Vm2cNCg
r+HVtrO4XrpdIWAS1bl5guXHoCS9DVkvl7NVXa1ubcuibUFiwQXnFNUB/BQWZEyP
ecYzeeatgH2dP35o8Z9hIfC6SfOpJrY5qo/k/x/aTzma5sCayBQ7lDvn4MDz5Y7P
vr0dXwJ00ridU67/rkUU/A==
`protect END_PROTECTED
