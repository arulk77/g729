`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2IlyfJh/qLht888ct6cMY5tJgwDhHwi3adzkkTdsYywuhZbsbWFj4XTcn91XyV77
4ifCQFF8ukilbAbCX90A1eWli8ZWYRxLBTYJiDtJqTBpzdMblNQOLT/fcWCoqxgi
lwKwK1rdDV4eS9Tc+4lsrSGozx68ej9QehqWu/mcP/CEaMOyUFXgGWqpXmEqQ9ys
RRHReXgJAn2dxJMFiYzZ22lbN3ED+4VbaDXpxCp7qpiLBDlWSPgnwqeD1mO7jBaK
z45XsqJB/czPw1H8Z9PuuqpuOhv8u6TQ/pKptDKRkOFAgE/ay6JHE+7hu0d1tL/r
Ftm4un1voZsXr4giaQ123XJxQlUk1WHNqltFL6FHqY5TzvsQWwUGjxrSGsRKp+Rp
QFYMFDcEYSZ0Id4S6rKmU77jD7UdCJYTeJVqoeDawTI4eNbHatYjcLW8AvDfk7pJ
GkLpZ3Rn513ajVxEdYgZL4gLIjwXYqQrZEW+XrKOCn5AdlQYO+sF5bn26gPJPvj9
Nehsw81Ntryk/gEZkZeX2aAlMPlX4kK9pFubvWN+nvhq1m83xAeuJx5jodUv/ftl
x4Q4E2dTL9so0uxb/qfEqVKupGmvOW746r/3nvU6uOkm44iHC+9nh0864qt+kUQi
XTgl9HoTEUOtkTQZ3dqSBtlp26/zehz99HYlC6abqIJ9+ZiM4ukqH0I+AUa2k1V1
psOl6G4T4UD7n2v+IUEq0udtpuuUNHvrLdxh+ybBX8l6PMDoUWOJeaLV/Nkr6+HE
++7TQhURsX7YKywCDbR8YTyIBKC7Kd8bFTWR4C/eL9qR8uKwg0Tl83tFpsd+b+US
r6sTRM6hHYn5U+CxBEru+QGTmFzltq2WJU4D8x53OJs=
`protect END_PROTECTED
