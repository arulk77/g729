`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SaY1gH+I74BHQRFWyM15WopxLeVAVWjkjwLrbeWsNLSD
leIdjIXxCCe8rTG3/06fkJjCIJItYqijRjGv+An6SGb3eL/xX6IVHMLvjJYtNEDW
7hqeJCt1vCHH05PYpC36gJO3VsEFQT7qepwdNwIj3IJriJndkE8VK2q7tyDgFpSm
WY/YRxTwNl1cT8YQJDepY7Wf82gZKG1MFz1e0rqr4+EgYWXeHWMoMnBvb9Kd6xxo
ubWhsrfPkCCCU/28eO4b92QdQwKQ5/YwFdT9M60KZNQC2981Y1AkqbneVwM6H2sb
mlCyRr+KETXa6cTQeXT2G8q6GEptJ3ynBujKEK/BUzgQ560OgLCrLFScrcS8zwAH
WRek6RDA0ZAZih1jlOQLMMh++40EzXGgBv+eVo+gzuU31dIzksReFL81NR9HNkbH
K4DnN/4TLrloSblAvM6ibENKLZEqMGSbk1BCoINrzej7IQhd0WcXLkoyoP0UUk62
9l9mTtr1GtZM5Kh5FlTQFG5UR60Y5lcQq5wwBW8IMVdJoG/vvUruHh3S1etliVw1
+6epMeIfz4c7hH/pyBwBFV5RFWd0jPFc8PNgfgPG3AWZFURwHp8bl4Z2WYktLyK3
eT5AnDJkCQDUMLTryVDTNmSUBOjXuQg3Md+6VaC15xjh1Ts0oQZQA36t98fAuv/k
NFI3WnDoZ5+Tvzi17rRdhlUtpEyhbw3yXBFtg2XEDxwOfVmZTpcNxet/O5Vk3xsO
N8NcZnFhH7k1Cqh8ISoGYWqFIdh0jSUqeq1g/Z7A4ZloIdRwpqJeTlJFsF/IjkjL
ccPda/wuXVOy7mYg1336nAh7TKZqQ38VYwijrUfDEeOW9cvp4TK1dbVPRjfeKTSS
imc1D5fKPujCXwF64lAGqaKMZu4Ql8HhXXMFdhA0D0eMa2kCtxOZTPEbZpNfHYbp
9kYttYXo4u43qqgvtkx/0AiR/ltm5Ke8c1iXq2W1gsDmfqcKBB7F/Amy8fFlnbyU
j2na98cARyNqP9yrCwJme11FGBkLTYMiTrH8B4uJ9SxI9wOSt8s0cYfBC9z5X1Ii
9O57M0ZE5Py3eW7gK5pccBq+pEEjjM9P6SyYUo47ebUmMxyBZ+LdmiNYPBuYOGZ6
+Mzo/lDd2X6j4L6YR4HtmvQaibtJpR7ItVy6FhcgFtRwtCmfANhHJAzGZb91Wxtj
t9vhtWVj30KnBuhS7+27Eq4YhugXpPNo+kCGp4azyHVXgrk/j+W6mQwi6yzBjqq6
k8oRykP/tkVDtABDkKildAG42MSHGiCtXrhEXYBtpbibh8I2giUWtvgJVgUxNpVw
VG5dPe/mcF70p9UY/0TDTEvihFoxnw/e1unjj15PNJHjEXDPU3wYSiJElTQwNV/h
M7jzJZLBAF5Jh3wK9h6uMQ==
`protect END_PROTECTED
