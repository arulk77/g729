`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBTMGtkAKfnlrv8gnS+DbjWI9Az68+67flOTLN0mCaUk
xj0lY4MimOEA6ShoIRYa7469NwqYM/mW0uidmMHRFFlBE45CcoAs65yab2Sz8aBi
7/Igxa8qmqFlCN5vmtKxJSXCbOne+4x0bZ9Nn07QHnd+oDis6WhkT9wfYpnptSQw
K1ZhaqynutJhMu9XMMWxW7UUM3Ic/DkU7jqCzNj6tM6Qe+A675BltLOO5GKUVDJa
jV1k68X+LOrMSKgvewC6Tw==
`protect END_PROTECTED
