`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
CSaPyS8psvm+/IHLAsvud8emxDddadvBQs2rPTzvn32WrZjfJUni7og0U3HGYmZO
4X35oAJhfNPSVJUV/ipy085ykrFzdNRWQm6Y8wPsVyMVOFewqnw8m8d5D9MX2Fi/
OFEULDaU8WidzFKAp01fqn3SAlqns0Ge/NOyjKdR634r8lS1wu+7ajf7UWh2ZB+8
e0wacl+ALcUqlyAazBalCToS9suEbf5bd9Usvki8L6zBYt58FS7cT5WH4IuxRBll
lj5Mf8sPtMPuslIY1qV4TlORJb5b6UcVU6ShICLWEMkwVzOo1WiksPp2j+0aBhKx
NSN3U+Yg71vsn7HZ7EqZAvA7IEfMkflCQG4i9Fcs/aY=
`protect END_PROTECTED
