`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
qjjqaEGBLFSSd4/jfms0UvJ4YryEFOPt8NddKmPvKK5OVKzozvSma+niDrBqAyCX
JfuHOVhMdzggdZaU7CxL90ORdTB4n6WSPV2izsTqYCCxdmeBukb/EfrRmHBnPjww
nQmX5BKX9Sqn27LyUd9pgDUbYgj9VDabe4LagLK8WrUKtbDCrBi+8ClsVYt7Kc0s
TPYFmxQ0KTk4gpk8P28XCWacOQPpG9dhy9rDbzPUrRdzBlGMXEtdjHXHdy+lk5jS
MPbFby47S74RdRaJDMIaKouG9Rgrxv1Al8B9qWnYOUQDnyiQx1xpQhZXN1Ce1ayh
V2mWAHRs2VqxSYK4w5H4izjEO9wcV7N1Apj7hrQAIKQ=
`protect END_PROTECTED
