`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN5cSh2lG3qBI6iPMFbPLr7KVPZbaj+56+TEr8zblQwZa
p04kkEElXv8qt46hG5fkmbL4GKTKJwYahPVZX0Uka4OkN3L5Q9RDKNuXVayfjOfJ
MMPTwgrCegpfBDRKhesBHotVx45BJTnQDCWFqWj/EuILnT94Lb7ST3tLQsH+tm3B
+R9VKSl2tijg529V7Y/1EIt+yYvQIkE8qHJBo1AJCnMyALWEqRAM7a4XNDRCf/nu
tBb3tAqyVf/B9yQmaadlYIb06VDsZUNPL/77wEq7/LUm266RIZcY26yTVUBlOF19
KpF2gMziPBAoDZ65f9t0aA0ReusrI/g2oV/ZWRF7wenMln2g3Hf95Mpn+05Ga1T/
wKFaNnjpkDPuxssaHRUzz8HIx4TL9T87uvQn1nDdkcrqXfE+sNOLVT2NfpPQSI5f
eeh1XktPp9uaiZslgsr1SWcVsrq2+I3Kr0LSGt70VEB5toCdDnPwv4dIMUNdbFkT
9C1pMhG/2yi2Va/JkFkMoKpBDkczEG9HQk+LRx7h7JwTdhJw1iTuGHBImXQfhesr
6XLG8ntBIHwtF5SIw7NntYrzDeMqXvrV1LvOd9od+p25T7scK459DjirvRFCS8O4
qFWCsRL4t79jPwRc521J4eLpn+2ZMxAZn4EnxDFzCNnGLvRW10gHrnB7xUt462R2
jHb0nLdzj24WlBHCrnUjFWJnM+AcBPW/3Wmzv0OJNYb4IsJcVtUzjtYOxFEsMlQB
cNTpEB15l5mIOaIKuAFonMkOASq0/H1n5CUsLzr5USm144DQprvDzvYQyY7tpw3j
MlaY1ENG+28Drk/MvYhr6jjyDw0vuZPOXvtn/8umwTdxIxcF2KKfJIhBFhMZx+0Y
wcgl1FLHMjGGgBCVcuMA3xVV32qUtSwR0UZHvGlLhrdi/wJ32zgNJV9/nM+kOtje
iYq1vtE57uKOhupsNVKqmFDfA3Ubg3yF9DoKYULdD1p3z8PL+CsG8oB0kf9xte9o
oSaaHqa2x0huX2p+EKaAIvPF/O9lfdPCVk1kHNcUHBcYs+ZbP1FUlNzm1QeaC2Ze
euXGqWCMlDd8lvEXIZQjOsO/sRMQufgu78cw3hsSlIhQLVeiY47nJvho4sEy6OUl
`protect END_PROTECTED
