`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
tedKnQBP94FUUUBtHfaP+mhgEXjomBQDJiPX679kHGNAxm9r0TzQwEh1tNf2l+g1
HhrplV15UrAIcR9PFPS/1EPQ6qxB+pQUzQgQxVAq3EnbPk6nPERXVJPCe8xEdFKH
GubdXAXs7Jwsm6+nGW67Jex3UdUnwj2IdpVsmzQaW+c7st6GMXhUfEmx4d0+B8gY
`protect END_PROTECTED
