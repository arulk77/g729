`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
fhMuPcG+uqJGEAEa2y6EoOuQgGLlfpnEYW9MFpRsn1LOme4kfpWY0X3Qr/KFnzAW
45fwn4GE4NisQ9pePPq4BN//2gbBJcvwXEAfY/67a3DgeFqzSTQaHJ0tfRdpuh4A
tU7uZ2yWx8vik90cFDi3uE3pPwnSpLdjneSF1SGkPRycO8nd+63ECBrmu5RdZO+0
dO8059lj1Npcrk957PvHCO9mz0EVneE9/OMmRBFLRjPTAmkU6ioxzxYGYoBQSvkH
`protect END_PROTECTED
