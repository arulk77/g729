`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDP3g4huxoqOyLuTFWQ4Hu3OkO0TW995BsDbU8flLRk4
tWxO11cemD5PKW3Md3AD9RKHNecXO1hOF3ehdgFi9QyxvXhi/wusgsCrN5TnVthJ
n37xDMwxvihiDLNJDyCzR6XuSaLWQfj3nO7kE7+Aqoc7/ToOsMTECzfxABOuxsa0
g4biOVkGO1oMpYZ/UUXhhLOAjMDtumn+AR8EpzSozwQRsJ8R68lNYtUVPxJ+/1JZ
u8M9d5L8M/ZUtQ9SuwmWvKbIEBkaGNZbCe1wwtsyqWQYJJqn2xMQignIIdC+I5na
obm591X9VRnjvr2QoTDQqCFS36v5tMeZCxRZxI9sYMzqelLKel4j2nxye0rziY2j
hKujz+pGbq65XcPbkvcxGlMl/cSSKbsKWndJQcB7mGxBW8qIlYPSqWPEq7FVmhAk
VrRHiwbH+Mc/1s/OVZR67L6ZxSfSKApFWWGwiRbocNJLT3ye1x7em3OdhYVOUBYg
/OcxEerhIAEsC/M1z9bqjmtMG03MJkeCdUhZt84tw/1ku+omqFHzSzWALHkdNRTG
s2Twkz3EbKgm28Nuz6uHufYDPYWptHnCOYZUS+XalOPMXuk8cIrrzlE4frADgQwD
suWB4Z6W2DN1fL+4JpMtAFAX4mINxDwLVcOc5ckhE2+s07oJGDyakzCvT5j8Q9pR
vMQSp0YGgkuRGrI5MK1G+tXyLxKrGof0IJFMRkqxdmtKZ+hp7DLgVQsphxKG/Rxg
`protect END_PROTECTED
