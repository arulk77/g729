`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aaJ5eAw2ELV+bIKbdGRrzvAE9ZRFZycxiWVzPouqxgEO
jPatoHcfgsANHbjifoXbb2smPm8d4yU8Ot/Hhhy2iCIs/yT3Mu08oHPnwgPxEa47
/eSKEvUCz5erZpetvCPJd4Dreqfp0XkcEGoZITPpkUZEwrJ6KtPzt1O9RoSw83T7
w+HjsVr6TiYFNpp076Fi38BP30ap7uoN1s1qvpGdzVf44y39+qqb2QqXr68O57RY
ow71NjVHcQWXGjGrLT/QYChLGz4gdpTdXNtKU5djlzCa/b/dvca/O+/ZohA5HHg3
njYxPqVS/03LUO3dPUdHmr9B7QpYTexcXEKOxLDUtL6r1tOmUTmEX3Dy/FHNvI3G
8y89RuQz3cYNJSEz14jLvMHvrICvzrFasy820qE1prpergbolvHUWO2tpeMG7ac3
3aWWsZRmLxABnfvv/GtYxkG8pat5rhcTq1K7ugA+3xiXc8ec2kw6Iip0Cp+Y2DQl
Kq8lZUZHQxrfecPWk4uLdz28R6u/69mKFl3ahu2LLNqzLozPId138wiCrfhdM/WF
XsxIvT3cWc9G886wwa92UvGIn0T/klokynZ3UpxAKRoDRDUalHEOyhDVmSV56rvZ
vC/Mj1EV3PBttQDzm8Tl/BdXol51b1dhBM1sPBBZ9C6OjaN12VPD1QB4hTj2rMkF
lRL4qrW76oMeq6c+2DTkZPyXVDia+B7OVuSQiXtMAC9B05Vpxw1bEtxiCIyPNKZ5
P0vG5GlWzXWxmOTe1hszaA==
`protect END_PROTECTED
