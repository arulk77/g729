`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveA9vjn3ML+VT4Js5pTILN+wHF61x2BtNinZ47NLUGbxT
XUojF6eaMWqiLh66pku58KuoqmugEhozA8uXToq8aMRdNQGbki7tFG0VJGPCWJNp
hCBHcVu+Ct7bz0aL+/zUX/uUI6kW3OUykgFiiEL8+dILtQIJEA1+GnnCuosxdhl2
cW6ZEpZblbx8fCnJogz6FVXbLDDhXro9iGaqiOYtXztgdliFGK+librbDVhwWjLY
2bEppyXmvrZKsbI2YqXo7tbG35BBT1DMwYxfVlerSsDQYNJWHqKfAiF9rxrPaOHj
W6IVt/zT4F4CTmhEa1zvn3yiL3vKaUx5VqTeGlnhDS4+ZpAQT8o6I1qQtmJ0xSNu
ystVSyx+1zy7N4rFl9wfeA==
`protect END_PROTECTED
