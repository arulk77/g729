`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3xbhqYpqe0dGnjgq4yLDlRzl7VtPJ3xUy+afugYpWgQ4y6GKhkTcHqcXsolRch4A
NKQZ1h97RTl43j5HbYk9xqEnc7wgepP8HfgdtJo8EcGqKQ0MX37an7VnzUjcgB+4
kWB+jR1IB3wLtCWVQq31BG3K26ANhnEsC9BESFUb+ycXEzTKkDUDWEpbH0kVdJaw
ShukeYpE2ymtqyXj/Txa2NgPKtXszMb0sSnxj2+osE3x57M3nyZzvonzaA2BtcOP
ETuIhAW8ONLK7OS0h5jY4uzlhh8JCf1o82o2aPthVDfnntpKCoIkAVZ+yMrnTmwY
Z8dUHGgXJGHg1nxYb/ke0854wc+a6Omi//3eu9KF5IrQ4HLfvbCE2qi9KjB7hPPz
jtJVm1ERNah82qgp6fdPuUutY2Rj/EDKYZ6XWwY8k/8=
`protect END_PROTECTED
