`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
x21Hle7ybimXzkmEjZxg/m50063JmO7y1YAPrsAbomM08Qc3GmugOYY14QiVa/iL
HNiMiiR4Zh/0Y4cIs5bJZuXt88bCiGAi0O2dKXU+Tab9TkctTXjyoFdzEjkQO/yE
WNrZUSNhVuduBp+QnZ3wTWqUBUDtOZX3LXVhhNQ334AfC7YysVpCrA7m92TwiB+4
iBOsjURjBknm3n265ldpnTpim2FbRuxOifv/+WWRe7dFbDNe5Irp9S0s+09dJ9yr
5baPk+ssgG2EiHO6RTBOj5t07rSkU/J2zNMy0RKrHG7ZwYik+MTUgRQBX+z7uz4R
nEu9WcqU0y1R/yAOUeTBty/byb1JCLvmDV6xzwNVUEx11lEaBrP7RybKqm/TEAzB
MUJtBDV76jPH0DwqHhPFDougfULBurXUUPhxwtLYvKRj4vEQRpvrRa+Pi6wtFg1+
Ebq2G5xk1mnkpMl8SCXl+mx/P6YFNmnCPjix1v3CdQ7vxc+7VAbZSi2tfUxm0YG+
WQhkfKw4D8SZDIBqkOA8cTNornEDNVrf5oT+Xu0oyA0WudkQQdfJGZH4eJOlpu6T
GPvJ5d15amRpypXuIZsGP3szc7O0iIVXkPoECHodq7S4ND87V5JhKJ3FEVIEbtn8
3CnTJ2vICDafrPmelncRMxdhc8YNRzmeWbvRDsngUt7DVFaiqPZtbYPtQOtRXbXk
ly8nGTXmQF5dDpqojAusvOTyH9/hAD2op0zRh2XeOvp8oIvFvVheeVwHARp7Ep/u
zi5i0rEpr8W//rw9PxSTdA==
`protect END_PROTECTED
