`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
lxVtamwNxaHTOZts2HKOxX8FX/J7iLOFK/g7FIVRexL9qiK0eOO1ntd1QQ9u+WVV
KrtJqDctG8K3pEL8mn0GXeLLPTJjUM/3zXj+KYr6AWut4TzGkxvQHgIB258fCzfX
3YAO/48+xkss3NujaL8xYKmtsf5iZBudpSIAo9ZqhMk0tdxNjCCyjVrgMxHYuiaU
2CZsJuRMyIuGoMEwe5G60BMn+t91QUevfR3HYBX8W7MXp9eiAgspwk+/3wMxaoVz
HtWbOEfweI482tCwU4fqtKu/agaysSnL20x0rCR1IsT5zuVNhr6X2LO7gHAwcz4I
qPMd14vvo4S3VXxRw/RlteJmyUjAS4p//AbBKfv8KocsjXybFi7cXtugCxMzNBw5
GK/fnZcJ5DAGFdd+opeFpREjWIUVdb2WYgKpMsuExOsjY4xTGmfn0gK4znSOmQiJ
PZ6WKm8a5QXpzI5zGapP6xwJowtDiZnMD3Ipe2zAhTuuIZ9/DdfOqCkIxOdf4F11
E3Y/lbxr3Ymf61gXzEea6K3/Mjy8TzIfB+KA1igrn55tvhJNN73N8xwNhtPkuxzk
su0aqVWp/Fjfx0JsLOHJuA==
`protect END_PROTECTED
