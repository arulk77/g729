`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47xtUK2NiOsnG7DboffEiPnGKAdkDYYMEbcRtzv4jmL5
QSXq3+z6caQ8o0HxREru8ongne1+zdjqv/WN4jBc4YM0NLPlSsExGjsJeiq7Dozb
on9x25yGR2OJNEvh8Dh+0z9RxC3DG5wEuiPoILPmRelOrLBKYTs6kApaY0TYqo79
m+Xm2h+hOEIrpv9wTxIVZ9JlH8AOZ3bI1M+i/0SU6Sg5rIF9cTUyIpVccNtPfYDT
znIbM9pUtVdyRkGRYImOPDIwYWh7Qotk9gviSonvDO0=
`protect END_PROTECTED
