`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
cP/ol0paSbDXCMh7XcrQRyDK5PERVtnP6pBhJrVKLVvyvzIOMI5yHcnQIYphJD+Y
+2Mod9ILJ07rr/Iv4zj8lGe6TBbPR47j8W5+I+LuEwDH4LcZD6xv+uDLF/Cho4RG
C23oSWr/f22pyzduJ09KufLAFdBzaz1SkcXzLfJp3jatwAfIXswUIsgW60ckZzQa
Vqd4LOfTnNkEYRso07aKEwz9YguRxPj1i5zM9uxttahzkHOV+wO/VUOXLdl8JlX3
dq8mmD4fuHbG/GjqMCvVSJL03H3UYPhuodD9O83PNK0Fpb+upEkXyGUtG7hjLtZ5
5o99TKPlplAlhFRtEcSxdb5mFmdOvQjkzKCksOjbZBo=
`protect END_PROTECTED
