`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43i2BSbk8TOlQRaY7SB79kSpmGXYP7kufvJ9Sv4+L1hm
kgSZzgxgW8Pau2Whr0MZ/NnlqsZHHMI3Dhr7GD2WvM4FXhdWsEivLzIpk2BiMLSF
+w7Gcdp3rEbIX99cBONSUOxWzbcv50xDGjdzYOmodSFTCXdGCKOs4MUJt6m0Vc2A
2lwk3b36RbAd0a9b0K+tjsmZDBkahlYLKdJwhJxkhPkR8sv1h6acUS633Cn6ejRw
ZhjzAQpwhhgntaMvwkoX/1PFuuZufJgh9P2nZ0GNvTnoAvNzEyAUi5zDlznnh2ra
902dVwxC76i1DYjeIarDU4w7hr3wYs2xgKi1vrXzjhIQIUqBjgJVWBBJBBeW+16e
gp4wQWS8zBxj+mIyxeRffQ==
`protect END_PROTECTED
