`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
odRXftWSqDi2NIddPyB2FH3s1u69SORJEsyip+GKfmIC8qSC7frTzHnQQdrF2bgU
QkxO8hNGAiXuYhea01URtsGBPSYAPJ66ncHHiEg83MHG4/M4NyUbT4IdnGHUE70r
0z2AtRNUy1eV1QVpRcb6OOeCrnQYeVIUkjDlL3wNz+6gpLRlgC//7fPrUBOcBzCv
11nAvA5ZAPLJSJ6MjOYvORvJQ2xQ4W7vJOg+WWimvBjSZbWPjsG5w0lmCNCsP0oQ
qiMTJGdDPxN3RF6O27xzyQwNRuKdUxRKVzPXA8DPSBM=
`protect END_PROTECTED
