`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNmoCInY6yfjKjapfhgvF2dwI2bEzGAbYEMbKF8sTHto
yb1zWglgraO+XTtSTe027FxHrO6Lv/tZju3ZIItxlWSUZ3IqtyzEnRIzKXMYT8ut
pnINQukWR6dLI17E8hkwrivkWJp3A8s+Q6KcAcEI8FU6xU7/v9xSjYxdefoiZ9jf
xmjfItrLXxneghuzqovwmOipuy+T3FMrfyMMEoCoZPJ+yDk48+B1eC+J1+7xx84k
Bh65VmOoty1zyAii+9juyTQaxY6u7sxTruB3maEapq6q/wNHcqLzo8RmJFHnGrKR
G0O2yoJXry8JGWlEfV43tQ0UN0exq1WPASa0QM1C5g7rA3W8qbFPrecmHQiUlQPS
/zGHxcmWPsJV56KLlMBjkvkSq+Wc9Jo8rQOH+UspVrnVZSY7uhTJIVG+0aFwaY9t
8odxLzlRT9CGU62ELqICmBgkGATBXVwXFdXmT4IhUd/CYA2oOW4rlogfRQb/pbUH
hYOshYebkHYX+y1MAA4bQAbZKtQccYw9V4zH4xVq1DfDCda8dLEddS+fGfd67ogx
esRscP5h+G9VUFiJRrw2aHnh1gxI5oas685bH2+tad4xdb8fYjbWvTWc859NIWqb
oyttDCHdiB/OumhGvVy7o8iS54/NbekD/Xht6/rwGywPuulQ4Ew0Z6OFtljuhH6V
`protect END_PROTECTED
