`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aT5cmSqFfuvVy7wDQJXmFYIwt/JZfzjJSfRFfhbOZ+pK
cVPcGFt+vg1xj1YlG5jEoH0TNeY91A3qEe6rzvPn8sxYmDtZcue738XQFjPfKqxg
eHHRaJjp9a9ukXGnR8wCA8NFhtmMdK+zuvrC0NXAhJqWclzVh+cdtVRpilcn7slg
Ya8qg5RpJIoBmxtLU1Iv+ZpSzssqBJtYsmL9dy1P/HlEjz3bu8US5NuhC2GCdwbn
nPMbRoEmWR1cyxxgOpYvM+/bbFL6yeyJ7DJ7hQK0oKuOXYtF5zLi9HPaWE+/c0Sy
hxy9IARKPCZI10tiSjTe0/WW7WTLd63T013jGqyyhjKI/ZXaSdW01JTVDHTsJFwf
gjiyl5O8zw1QpPxMWptm+3jCgUKNwTzdlmoHzLAHyUyAxj3p5oD4I7+5ZY8JpAxV
wbsuIQXJFkMBCdhXLxOAfA9njhs2rxl5ADDiQ6Zir3J41oFcopgXfioxw7yrzxFe
QqsBQOhO0bSr2SG2Mp8xtYvAH/Zl77ugrJ0RKZVsTgfm3Jg3xADjiHI+HNvYxqj7
kESqgw173m43V337bRTxa3Nu8evOrXncWjQga3tXTN0PhxYD5S7KAd9hb41Pfae4
msa+acDgLsa3AwP+rPIhlaAJ+6RMCXf2UWcG7x2vQjm13UDWRmH77JB6Xypwkdkh
EpgaXLppiST6NhR1M1V3lkwt0PZ+YLI8zNyjdgEY/xD9kuoo128e3KiCMx54AAKJ
daZEkhCR/04tF6UW3CtFQHvEJRupc7xtWEYp2Ukv19Y=
`protect END_PROTECTED
