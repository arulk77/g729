`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ernQLpAwSZKBGOwjJS8ATPsDBMjFYx8oJSu7Hok+67mgcvJ/IHwlhEKHf7VRrS8L
fcprxKFLjF6kiG4NEzL6aXsmWqZV1a8Bn5sWdQVi5ngUb6GbrquiZENYth2UvFfv
zLtpe+wN/9frBDRRQg2/a3BIKiFeVTDFHGyEFB/n9XPDF+PSZPcVt/Q7jqzafXDz
3aBUa+Y6BMG2BfrpTGPPiboMLO0rjQkwzuguc3T0/s7ZtCrEmOj6ZV7rUHc1ypxR
nrSDDYH1lGw7zs8BlnSQ1Omq1KzTazA58wKh/J6wB/6iN053VxZphOXhJ9XhalUb
sQIzqOmjZ3AQFDiI0PKCe9UcZPwd57ZToKeE2ZLt/6k=
`protect END_PROTECTED
