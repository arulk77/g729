`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLI2dlj0xhNUDw/v5IxGl4uPrF0pLwdjCMkkFl+JqG2a
Ax3cdJefVytKBFrcJlPvno/u4KPpA+Chi7hAIorWCU6N4xExc0qo8MRLJ/C97mDu
PoYYaRpfTanKjYT8VKRAYvdbJYR/AyNYvV17FnziyhIDldk8VKVpGZNPD4J9XrFd
VjwyHXoUitpDUfkFv5jWD8bXDrrnaf+5DFjFNXzkhBsNL1iPPEK3VhcaQOhftYLE
Z8vj5NxL9jjfNQFHBbP0sngnCr61QtDFr+LDze1UAWBsvIsiIN39Gv9Xlmkg2MSM
kWfoa769MawF/i8tYV+9c43I5sBpXOfHP70TnZ5YemAEAKm/VlAxyB9TDD8FmCcE
LO7+ZO0Wmt/nItJfsKPii7jotfcAimiCaXZaw0ZCo7/R2HPQYociEJN4Tv8Uc8pJ
Nth07uTNfmVH4aeqbcVscgaAo11fZ3Q2sqtSLkX2pFS2LRm1t4C1ZRwuAW6MtBKe
4sEDciRiGuHnQX2q4I/Y6mBQhaeS0lHSMpTExvS76BC8H6FdutBnsUaJYTtS3rqo
78GlQrUufzhCF+n8nZEns0rZ35TonN8MX4nmKdSciuq1kOPnmriGiZIVi9uBWuj3
jZkPLZnUcVdFQhFJecmBV1YM1Bqr8rKhpOPMHE34n6ttN5Wq0h75QX91yT29+0qu
`protect END_PROTECTED
