`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C6A4ztpGpSZD3qjzkCg1Resb+gBVsYloG0S9e9UxyrYi
O3WMhg7jz33kAC+V6vTyJwFh38TsBUWbx5kfaxnlhLDLgYKQBrezJCS76n9wdQq0
jzHeUU3RSK8dfFlHkZ8nNgOpclOLlmgiuVxsI812XZhI26bt6ys8ahQAxIsfDa3Z
MUn9BzkfpKTx8ex2DgkNCN3uRUUy+/htg8aYAFLf0l7gfH/uop2Itm2beYI+aSrZ
8gBtIDtbzkpJLtzInab7uY6sadMtSjQJABeqxwLOitf1PKHoHxfcVIB8AsKJudcY
R2fAF+pNvFcITR/7UFCINHd7IPJJcMNaMZpvZjUXoO9Dkm19QTWWTYU0CC29uwAW
Gh6A6pyQNFEtCQRuWHf5tKPq281RKnIKBLfCvynkX89NnFvQXk2/1KGg70Uz5zUW
m83OAG4pGl4hWeruQmfwEcWz5af47YFtg2Ntc3ODiwqzkjMil09s7HCgOz4MYoiQ
FfpSvuvJOhdBl8sUyZlN0QZ/Vu+P4YST1+GLCNjdSSkZeSRZTS2b86WCK09LqSK0
CgshmOmthbkUzoOaO8fDuxhO5EhlLE7yOvEJNn0OdRs1uJFEGhKu/1AFg+nARMS9
766njenjde7023AUOYF9Xs4bIIsB+9iIoD3kNM6t0n7w8Im91NNDQok516bGEf0Z
/NNq7Sjwtv1i1r511JatBmI/gDi83JO8FQdcsN1NbvHCDjcHYVPQLvxTFTM7Z+PW
NsGzA8cW3Rk2CEVXQsP2+uw/e0S1jRguT/8s9gD27/kBw+rgqwEjL0W0ZKzYsT7X
xw0eTWJg2bie3BteF4Vu0XC2N3Q346gXK7BRKLskOF0Sm1BdP4hBwWzKmFbySblM
2B8SYVL+BrIa3bB9NfINIgYNHuh/61kAc3yqhSJglf0rK/L/VLdUP7d0HxyJ5lBD
`protect END_PROTECTED
