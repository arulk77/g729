`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
8QANNeTqHvTDs0m7m0LB1vrFY9SIG6xI8Sf1Dud6UeMYhMSuDV7uhfD7xWH1xAIb
q59szsrcWp9uiTRg1lXy5e6z4j4ybSAE6eODRUgXjykiwKV0FuOnX2L7Nhuo6L/M
j4MAJY7m1lw+WfHqP/5p+IGnEonrHdLIW82gr6OMfcXEgHH4JiEfJ5ZEmFvgBvHf
6pW7nGipywjsSOi2KLAaShoHlS2CD0Wt1U2EoSePv67qvLy1UHqtsJIdhGL4eGYK
tFIaf3V1EcFohvB8/2u26RenSqpD092NRLtJNoZGwwlYiPQ1uxOwYJvOUmmvFAEb
dpsJd4hYRiP2PVVdxngXj1rdB9qNOOTcRwUTg8BHZp3XdTnMEho3v+fCbwfNqpQK
bFXvwRqu/AWoBqv/xGv63lphAToo2JO0SMF1sYaa+NhNNGFkENe9cT1PGcLr97mN
`protect END_PROTECTED
