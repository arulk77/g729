`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
7VmPYNNHXfmA2xcJQePthbKLGunQwzqSbPV637DH/uhr/XJRFG39y0wRUXCCKdZ8
MQZGItMJi1mSzmDUWNlOnzpgPgsGDs9hdq5byuOoKm3YE7r+YXIwXn3bkQJcV4Dh
4Av9lSadqZb6MpSJLW9x88fxgZXqKzJcUkh/9TqG6+3uf5xaUhYIws54rvlildGZ
ufDuUjJI9KSIGy7Fh+nAQ+c8/vmC6zl/RnUIjgP2kVCFvHdxlTGSy5J/RgWzH/tz
QjAIzBISlwfWePeqIvtTu3jfZTcLEtehxoX1IrF3dBI=
`protect END_PROTECTED
