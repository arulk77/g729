`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveO8bdt255xsYu3EJ7CImCJajyybAHJxgK/gJ2Iet5KcX
0OnQi19tOCk8ZXGSRMlB6dEkOM4c+COQBf3lIdbr65wmUiiAqbPm1NieSyRqg86R
PP85uu8xcK5XkXbofCbHU7SIw3H1EIJtEuljmJ1Xca2nXHBQWHbMGEHv85+orQTW
8+Asz3ifkTXeykY3xJZHSloQGrKusbWIn2lMHHbzRBol7P44LfUh0mMTCd1gAA0h
CjT4MYclEltt5om8Vfr4lg2LemDyCtoEuE/k2cdDwun0T280ETC8aCD9CtaXKeOw
IrO/B/9V6Bu/8pnQRm4Uig==
`protect END_PROTECTED
