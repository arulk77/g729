`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Hq1z7hWKPwusT+5EKeikbiA62pmCGBmOp5KHsfaFoJgchxpwRDFXiVpkSjMOdD+N
OlnBB/NQqBsm4IKe1M1Gt516ViC3bm1atwncbvu++9ogL80TOGA+QN2sF/dT26Yg
`protect END_PROTECTED
