`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAShfTeW+behjCqmUXL6xvV8j+2e2GqOvd+r75iJ2+uif
zT8i1sAV5MZAEFbK4tuUXBYjDLNERGrx4wKa8mVi7x6AhU7VpEXyldOSTYOKctId
5WRLlXjHEQTP2ycTRzZESRnpcv0WVVAXnp77oSccd7E7tVY/g+JOh5/5gTJPRu03
o/l1lUfW0Dx5ADdO3yzCXY78Gdd4Tw0L827mvI2nCTtbDpce6p2om5qMZhvqNWua
vVvrESud36Stz7mmpG1LKkCzHgzCY4bYMvcVAc+nRJsfYZYgM70qRMkdN1LsrEGe
9ReCxAQZgsIES5HAC8HnBhdOZJGUqdJzvAbp8X7TncskfuDMkPa10bRpV7oeXEuS
Km8zQDhywxbo3oeDsjv2QcgtWqe2rk+BK8toZJhvRQWrGYdrCezEHCP4SZLmb8v8
k4zOu1HAKxjvl54kfawEUAkasSZiFxTzqtNzVRErBWzCOXbbKyoyRdtZyZqP7sQY
iQdaagOcyeBmLtZlnORgKJy1Ncf28bwx50JsPbLt4YSKtdLcZ/cmE0uUHNkjg4kx
9Tb6oCL/RJvBdSDR4vdxy1l6E/3dMx3c6SsNpkqUkkhPag4IGDxS0m0hW0sdchXm
jrlKs99upkIatxRlpDN7+3//Sg7CmnnsIoJfIDuIXjac3zGsM7Cxoq+JPtAGITE+
1BsIrSaw16vLsb3rO3Z4WV/bMAbgCQtqxhVNx1Yxqqi3qaTdipm8ZiS12rFdeWSH
GYp2I7YoxryeT0OmzaVFEycSA6FNc/ihg5sPXVk960PxvGoUZ3H0kCWAf4YTzvTP
tGadaTgYp+x393Q/CGl7o6gLegtGvAc2wYOFyZsIWjBCyAP84btnHArC15vyyONt
JeUrDu3kRkC7HQzpPI3TMrlWqi4qibEx9cdPdSf/huNI+cf3sCb7Q2mBeWTfN+Lv
z4N5Fqabz1AcarA31DlGsHf7E13p4hKVQFgSyYRdQrG6bw3GMnmoELOcvEE2rGiL
xkYz9Q8FXKdIfODHdKBQgfcNeN7mayE1c/Ap9NwhRJMtjc33OYyq5/ekbi2lfHEB
YD24hS/HzUno1FSYzloJEjGakfclTOECHFO7SfvNSKci5T1W/7U5dSkce7CgDr4w
QXgUaCfz+4AgVuSFfJbbRioYKibdiBxVkUO4/99LtHA4npJgU+YF6pMAhATEHOBG
arev47AurU5o6o6kL7O43ewJjNfOXruX5hUEmuyril6iqXIJslgVMm60eAT0B9JC
v6p5rKOAa3YAsdVyVgT6S6ILNTirVdfhQ2g5fNZF81eqzW01kAO+7/NT61s1RvgX
6AUVYHqPsEJteutUmTebDF6CjC2/o9bDa0IrM3WjMLulmNO1JsXp/IYquEGFEUWF
wy5vqP42YHtGmrPRjychH9WM2sEceNW3rbDxtFPNMUox9/W3oc28CWaLD0RDX5bq
0wajfmeEwvRSX3RMLR7P7ow9AG5MN+HtQthXC+LBl5F5hno0OddYujpFjVDDcl+p
En2FDnyBypgEK99HU5Gv0qULky87ejOUc8K6QsBFZTh+nkYwSssN2V4CTlYNvY36
PnO77EbhQOfyGuUaLDIUeFZudb/Zf7AjFjkoygSrbbk4T93U3OvPCyb/z96owQCN
9PBYQXt4vqqd2f1jBM2ozZQ0/HMPY961NBsJxeBIHhHcrDiOPCJ39kocTKpSJvWW
Y3MaJHbjVbb37hxTH2R1Fu2UvkT3mvTIyXHvrTpy4U3DoRGcevVVR1gpvfqzUOaq
ErsxAMIp8lTsNcZWhpr/TWi4C2lySJVWLW+ILbKBMxsPEgpt0NRedpVBzTzjzAUw
3SP11j3ISMcTkyJznoQROSFuXUfAXUsuUXW6eSb9qzPrjgM7UZ9EALGOYNGfbrJw
sPgv/J775YmSarabWYdUUA0rlKxnv2f3Vcdl7NgttGj/Z8gOoWVFv9JRbRQv6Ij2
sfwP6sQn5gMOZ4IRf1aFDrs5Vp4GnknpEcY0Mi/mRZ27lCa9tp8P6teZ/6F/ijOx
9Xvsq+Ovy7RCh2jMh3L9vufAjBvB02zAGOH8j9gaxb6Ex3A0roJIuW2KjsBt5jca
YkjEv4CV7tcgUyQ5qpLXvCyM3sHWjcrGIO6xW8ywJvqu+K8zf23wYaTsIFzNco9V
MyfYkIZDU242t9nD7I/mgZiGAd9O1MBzZkWsFye0kHr6CfUSkX24B/GB+mB2vAmr
XxWtN6A8JaMXL+hwyi7jt3uKVM0ywIuB9cIKivsabYlrsBLxrnUFw6UjvOlZ/P3G
lsT+bV+TONYAD/NfXLRyXys4oa5A8zwZn3a0H1QwHVzA2N1ykTgoN+dm0b2UPugm
fgyhazGgNQy49bEWJOGFieUuSOqnKaVumYSIOpQJwPUUF9+9vxzg4CdsOFKmCUO5
fbasCri5sgKfzSBz/HR7z0tBtt8A2qmQGFhCpXbsQ9bNcWuDCTZtsfk9AoT+oaAc
fIIC66t/K+bmuXFUwtbJngPS+cxVLV/d/2s3YxQ7TnrUlyx1sUbweXFzlRaNfjXG
HhfIzy5mQ57xZOJZICTAZM6OS2qCFarXSVHrvuwBXDAJED8umaeLAIW2O1ka2veG
NYwlPcC3rIYcbZPF05XhY/qRUvsf2ydxhInVT6OBNgC4P4d/pacyVoQIlQp2gf7H
NUlBbRdDBRvMGr92Yg1FPcVNiOl6l8Apx7G+Mvhq1nrOJ98G6SdbX+fFrkQniSfq
1/a096s57heciKoeHLK7q8eX0ZvH5SSKpyT1MGKJfqKr2dNLDeW4HH8GhoNBWxE+
vDsv+96tVMg42xrsx00oIRgsIWNtwYU0EDYuxu8EfsTsUOeOitxhh9KoBc8r9Op0
TwGKJ21feB33r/+SkVwI8/0VW/29vRKUKQgfyrDbsqSAixr5um5IgiO+1dWT35sn
+ok4/h+0CdbzEQLigOfP/0NnkM5cYujulna9jK312AVXSIeZ7tdJIauVDTtrC+RT
SBrI4dyXXosRCAJmpIZyQxbX8zx/75ov4qFUr/zDDmF8X4zEw2SzNGo7ARmrUZj9
zsw9F9hyRg0pc0yAbob2iwcGePoB/B2wuhDZPxdf0OlXQs5D1L2AcduMzlUqSdW2
e6p4noXVNcI9vv1Dd4yUoDQp8ypt0TmTZM9OPmP7/9asKqnfoLvIGr/5R1vmO3hf
r4uoBqHEFimCdDkwdYapRQWZttH+otvdNuZ6a2kHAlPaFXxwOlD6cmN6lYJh1hzb
WQpfn/AebeEOhp6lZTXflHepR8zYZtv0t2RmpjLmAIe+RkypYdjRGcF+ZXlJy0H0
u+hNwn7HyuuymFaw2D6g5ehgGqS4/ALhXthhXJ7RSvvR22yTbyjJm88/ZVOq2q6N
QnhSi8u8pQdH4HwyVJVo0EkiUcp6vVwju7aO3ns92JvW24Liz7gRL7uz0fPYCQ78
aQH72QpH0EnY1XV1yHPWu1cAwRpoR33aVO9LjhOhRLZE12drOfw+OyF3MmggpAyR
67IcUdq90qqKNkAPXok+cGUU51lf3/PvWXWYxuBZ3U43N4cFMfMQs6UhoeW3GOdw
IUP3oKq7Opl/GmEDDn63m0bf/pVEffQ2ecUZlRVjjl4ZJBGJfxss5eceJSy4T8gv
BCAf27QpilCunOMncoElT8KeiR3YkeW9bAPqgYMJ35D08zMN49VgUUnz1XRPhadu
qXcieyFh80B+6TEfbHkL4taDCEeE4GQ62RMnXI5ZHlVQbUiWnCRqfEHPH07C0Gll
GYSVGL4lp8IqTjKyVEhcb6nHkUDkplVwH6Cg2rtgO68kphxg649BEW+LvcxQKs5T
iZiFarQLHUHnue/nalXmtkJ75VLXYdKp1byX8NQwjX0aLfeVL3x2SRKbQnTLdpAO
DIfkc2WxKp2lod8AysU6gaUxfd5y206pf8qaRZFPtPUM/tjtU9tA4YEnz/7/ZtW4
DuHSwjqNsL5GmwV3A3Vaf3JXB3VROqwgA3jj1BYBv+WtHLuHinnUQI3UZk6S6vlP
bj8EnGGudCn6eEkBF7C7b235w91fwIET8Y/FA8C/usiGYXyxk15C+DnqtEcQXnro
2v/Gd3DbSSwwzq5RQFPSsZkT0+T+ImMve72xuoVo1fdjkKijen1atLJ3PCB2uIgy
zoFnOskG6V2b92s55Z1RF7LE5lx6Zqz8duRFUoCNNaRUUFOZXYp1piOB8YBjiUJb
cChQlXq93ZNGAH+PWwrBIjDpvybXdAHVQPIBpTxuYApPyz/RPAj069QO+6qIVgrM
0gAZL1RPgLehzFRytUztQdE3AI2rY0XRxNLvhTy339EAljvQPDskwy4YtjrmUiNW
Znf0RyTCM+62ZYHy/q7s5e4rQ3P/wARnKozu/D7ixh2vJUuDaq7RsbvTY0gjcOgS
dchMOCQh6eEcxxj929PjMIHCMGidiMM0K/+wkbEhXrOwoWaRrpLMIW+FgHeKG8RA
zOOFbVaSznBKKBVj4wmyLGkB2wp6EsykJizp1/A5AV9eaoO4hlKBaflPtdogO+Dn
BeMMof6JyVfFivYmjtxmSBcc9AW0l9Dj7bLqDuC0ahQUZoK6v4UyU4FQLZAABLXA
aG5rzgBdLS/ffbY75nqwMyT+b+nUPAkEEGpYz7UkhI64MUS33VyfL5iBzmDCeUe6
r2WxtTO0q3aY8uZWlPqRjQjL6dEcWXa7ogja6m9XWdAV07cbpTbHTqxfTXPPRGTD
jbAGXNh059VfOCttAu6wL1biadhMGbgzgu3/8gcmNMZpDThQQsUpAHe9jkU9twTf
qt7TNlDNrg77vkRgR7Mxp/rK3i9x6PX8g7kOG7OSImPXycC5l49ExHXyRDQ6GwGo
M6J378M2zqP1xIRXKVmHSkHQVaBQ4+DxwncLibjPD1NF4TC0uWNK1P5ZgzFN24q9
Xfsd9wNuBaN5wJdruKpYdAd2lSsa6Jnp3wuB5PSlVcW2IPrd3Pw5EwiuSoTKF/Wj
2D01L5V3hCEgaLgbBdHnfhFiCrBwhyEFDkxAPb6RYcZmxsvxeBB2ZYQKXtEctlLG
BHNYxQ/kOf+9uZEa1xJYII8EDUGipoqCYE982yo9C56FjFt7PPqtFoNIY7k2aFU6
89GARNWMtPRhBdX8kQvJMIMgCelbJwbQAOh7x8jceTI1Kg4Pcvk9xOO1iTOTWgVn
XhJkgqShoIbUmjSJE9Cn+r9gIMvO+yX3zCsEXw/WT5JYpbVN/SYU1PKyqiQdEics
96TPxdb0J/DDAAU1782zko4nZHX4cn94SA8YH6dE31cmmcc54rLeXb/l7EPPuTYF
U6Hd78mlB3+DywxsNuz/AWhOQs2HgYUuhp2RiKXgll1EEobesaFUIMDKROqQVFE6
xXb358JFHkrQuZTXL5SEetPNOgJSov/TlgRQGz6EeQwbrwcdvRu2xmsnLg+62eyZ
zDZJ1ivTSMS2BTAzmefsoW4//SwrZephYlXuXV2IO+Izy503y4eoW13f5i2DULik
WFlTo4tC6fFOTgV+7Sr0KhvAG1dSSOgyvMVfhJ4Y4VTto5zSKX4NnscLm05PX9Eu
TmhSYpU0Lw6ra79CWkgaPRYA1Cm3EwIvgkD4BvJpeK3MMWGGPwlWFmsrxmbFSPH7
9Yl0TQSD+sZSFjF5YRBdpOevZlGgAjMgRXbdpsBDsF2w3HkSl59btn6iWzkChnLy
1/9nkgGEtDwNLP0Qq5EDp/v3D9C4HFvAeBmpo6jsK5k88CDIkk5UkboYMCAVdEdb
qji75+BobLZqKFQigMwOS7WBiqheNRL+8UVbsyhl5xaiShLcNJQdLx+3qc0fG6te
ko1bg6qFD6lPAGTdTbuKdAP/2jm0jLL/RpLWLKhgEAFeXopjFNsqDjGa0yQltsxQ
0Bi5ZSAgNyqidxSy+DJts2ZKe+cSz2yGl4btix3f5bJvO3VGM37/LT56Lv6bTnKD
aPVBaWq1ADYwwAg9BldZVekRX608FlV1Cu2ltOqKxU1gmOeDPb6ZEHbY9TvPcaXs
XkjJ0TFd6J91EkRiV96ZJoCXadZTgr6yZrRxJHp3BUfOEfVqxmQ7hZOWezXaHQEb
FHPBHh9kKzGOcRNJ5escYhnOF9ktIjwCAD9zx9BlnmH+WfC6js4YH4gllYxKI5C8
CY0H1BIrSDGKZ43oIWHYQljDHxQtl2blkDmqkKkJPujAQ9TGdaUpWkIy4Vmvnjfz
oGexLqqC42g1XRQQkLUYtRt+y9UJDo62iw1hHUczDMqCPX5u5BT9eBcaPVFLZlaS
hYpbG43BQMZ4rEEWNQiC7m/+oEtUIxg450TZaztpkL7ILoD62P3c+rd/3OTHlWub
2ZXImbhI2RUCvBKNKPdr/5wmiFebSUl9CdcJHCMJXZz6Lsf618nObYEY8xzGn2Ar
MyCVTdPAG8m4p8xiTbYyAsvXrrOQHhOxPCWe8BMxaE3gkgN0kC2FFSVToFZtjqTA
nxyXiWf3a5J8RadtjuEKOg7+P4SYyYhZ9DKyE/5wNz7eKM3YQyN57eYzdRz0O+Ih
WLDu9xOP93RjyhsDjmtOqGMSdBNVs1f3ZYOmbEqkwgfSQISCU+shu+UgSm4GJnwD
/jsV6nElBwESduMlzeXUld/Wi2OGAEDGGTDbPw/yInb5/JID4ycmvXQ8zqvz2ZKt
xalKpAkRMGiHPAy6BAr8vSVRUPO4bysNjwxYDwX1SbdhcHlxpuqjeXHhJGX8Gqvd
jfla/1IyJjSHSYDgaTB0K/1+Ak/A8Vd2ZqlT4CXWni46F+ndlxZdQfvLpryK/86C
XjiN0GoHqN2T9u0FbXfaQCOor4b7OY5VYEQwqWaHkntSSPKK30LQ+LBYyiDYHmAv
7Z6UxxNli6ZPJX2lCElV58SB1X6y7TF+hczPR1R7xxjmrIV4OXQGO5tXA7Ni21AL
82trcoAHbpACD/Bg1p0WNRz477qy3mhJBiB6Yg9sprdLNirh0CH4QPc6JCURveV4
jTeEI9GKz7EmtHyj8ssA8SSReXyfzUAECaRX+elcOeK59yOIAeobK5rqRqMdDu4h
3YOgJX39lnkTGCxLkUwysJW+z0SQUZxsxkJbxEeJ+GQ1dzBF0ctp2WgP0e6GAZ7D
h+r6gQvap4Qgky0nEKUUnbPkvySirVgPqU1f25qwWHDmtxQalKifgU+uKT5scXmJ
3mbPJ0t63sXfjh+hNFvJVLrJi/D/wnB/uQBj8vNnyXUQAXc/kI5O8WVqFaEsxNwv
6si1eJmy1rOREMdb4ErPpenV18IMmUDL2oBolZGQ5ga+mdaY5/e/cUuxAgOBBhS5
eNPGV46KJ5lODguNWcAMlN+SmfYV7Zeg2c+JzgrNX+1CTJLBe8+RqHwEOGmo68Ft
MQkOv5RU3auDEyKzqc9h8a8UutiFjajPsZKZJ/kgZZ7QHK2jwbr6L8a7wCTtpyRn
pcgoFFptvK4gc9P5kthUyL0eGxkeQY6hIyMHMd55+WeMR6EjlZPwOqOMZkg8HN4t
CdhavQkR+P54R4swUUdPdduhC7dtV9E+iGGAxv8BS7hfXZv2N8cF3ez9h7BGA5D8
1kejm8/gSPFqgXqOSGjVaaFRt5O/GtByFWyKlbtnK4GFP0KdvE86gpSdDo229a/Q
Wsm4Ze5Lekv6jBc7qc8A+eUXBVY6PSr79U3DhpUueAf9pkY/yWNNPYuxVYT47HQ6
kQXfRW9jiBdxsuOPf/pIIuAYmgXM5N1zyG1O/Bb7p7UAsnFrN6TBkg0gZWKY5t3W
ywHp+BKGMFrtgHWLYBKsHmoJngaLiL/kcvW2B/gSddvhHG5ihvXF+T2xbPvaBFR/
S7+QixQwg6UkMzh64ZGFobfpFPoO2UIuLQzeYwr9emSHtY7Rr363GT3wrA0c0Tpy
an1fe6fAf5Ya+8gNgVyjuJAWdgDpCNyUbUJcfOKiWabEu1sKCvuVowF2eLCukeYF
JbbTkKMr7YZwpyXvwZLcAwQchOS7OEXq5Y42Ikkq7ihkriRnzyKQ8waVtpMnliIJ
L+bbF/LgTVthoycqRdwYI1rKJLJ+EKJTfhIN0D1Bl8Q9DUxvGYI5EM8SGwbPPyqL
QVcvKM05DoCZYyWoRfGge5jjeDqOFNlW9Ay45eX6QLnYQgEkveIhPRYWC4E9ER0o
D+tR+3XldO+I1pneGqzcSoJ5uqcLL5BMruLWXAuldZoZ71xq3JtPC0YN9ikvl0si
sH3AiFI+orFKgrTaRZeoL37e90GrzwTipqj8mXrGG0smIuaNKVAWLuhR5uzy4L+k
dNeEL1sf1Y5urGJCZykKL2t4oyRjUr0GPnLgHKA1W7gWGBzX0rNWw00HiIjxqcUe
jh7TOwtL+qCC2SZ/Yc87ZI813JTprTgvRWGHxF/Dn1u2/wxogMNP/vpYP1I59NiR
2HaMnlqlIVIcnDV4YRgdDKccjxWjMgsYHIyooKWpQn/zKoExwYS8yf3zfK+GNYiS
g41r7YEd86ozFFy09DLd7GhiBV8mcNeJtDW1jMDdG+q2uhF8VUGFa/brDvcodNNh
B9TOT1UHF82l5m3FMv/EbtRrZ6P+bmtmIHMdShVnOLd+Xk21qam985kQAIMEAIqn
zY/jaxb1iieSCfNNLM9Q6S9Ht52asHEkoFe8PycSvZ6XpoChK16y58jAFdNVSWwX
y+85NKZj22J2HXqvE89wXOOi/h00n7obA1cbalGe1abwa4kyJV/eoL2Kqwe7qEpl
44p6Wut/naOc4ENbs2CLEScYrwgfgcBWL1nOK5NfVoSGXJVSL32fcvoMIxX+O43r
CWppxz778IvUz+Gndad2RcN16DwKVSKuZHFPMRMm5YD2KkU47MXxi0w1kvyJHvTJ
D854TwkCgHETPUdk4hfn0OIyjjPgU86XUc5Sgh6Iyz+iGPOx4oHi7uKba6M/hZw9
rRu5gvq0UELBzEjGT/Ul+AHVeuA/SCry8C7CW/5EdmHWAb+7toDS7Vz1m7YGu0oP
Pz2MN8T4HL9htH+ThjXDi4sTjESF7pqISMIDNBuOsKFTKxzPdsFmdn4I/NR1tH3S
igSKU/AVmtA+4D7GRqlF/4cRtm2TX0RWhLdVClsJ6dl/zM86KDZxMSR+yRELdvRJ
QKHyXz1UrBUXKiUExoK7adqMdA1RnFhufIYDBlFli7VOX9V5szSukjZJ05H2ZQoA
YDX0YfuiT2mv4koBP2sE/KCtFEGPYuE5kD3NjWc66vCR/hy7GQssHwd1EkyaEBK+
NVOXnxd8jLRO4kCMCjB5jSzCBM9yN1KOYWFAj6HL5zsiifOv273jV/6MzLAKCNAy
51hdNTYOXE86TBLGGySTy9z5mj2Z5+xkZooY7kekHdmUP/A/KKDktXl3sO2+sjAC
LixVOi4tY97W70v40DgezqfrJb5QkhFNXN2LowguF6QOBsl2YS58+bPuypq6rsf5
DGL+joaKzEPUGcCeVyAltMdc1ERfu+0lZUWYzR8mTJ+qi9S9s2gUeEW9GnkK/kg9
YJ8qWCC7rUuIZ065KcAiLX/2pCw44Rd7cCv8UoHyBnZTmnNXpkeMlMVZNS/hCtAF
gO5YvwcrFXKIKDx94EbhvPTwifFXh3O5i3jTTDWmVHcCwVUEAaDbDpdQPApXhJVD
ale6DEQb8gQBCLnIolXuyQs6oWNWtIV1zQ6PMYkJQwMvYVR2EqaOw14L09iMTQZp
DdwosEBfcjV5PvXN9nnDZYuG7NVja74YCh1CPZcuc+29xfZ2xKIlE++mGdD+RF4c
TUEHnEPVJpPuST4oFOdClpiYCgeLc/ddgG+UEmBceg5nHhV+a7lADnrvqcZdxN/B
5uUc3ZVt8IcdPe5xdJ4/3lTMgQU1rb5FZYCSAeVFNR/RgYDRsmaG1MeIVmz+tA5Y
w7q+vMDRAzYGjZNZMUUk4flqt90waBs8jMS6/D3IZiI+Rx2i9h3taXEnZk3NWpdc
wBBYbaQTx9XtSlir/TsrWl9Esr6Bh2mtobQtWn/fi33YoxoaSd4UqRiHjgu2i42C
F19gH09T+SzxRpwXuQyKbd25leDEuB0hsrAjW61HnZMMkQzBZE0kaWs1mUBJpUOi
Vp+zProZjrVWGHEczn+uVr4HB71k0Mux97bbwrW1j1QOOTKl2THCTZSlCXvgyvrI
6irklyxbYOvUgRGRqHljQk6tlIheu6g+spEItr80MwAdzmXJjbx26S0U1MsMm7Fj
fe7LB2j02jYsSzCq3/L1geR6WgR1N2nqDzS/qcgURsSK12Xygi3mY2QnIWivvwiO
SGTzqlqykDKhG2yVEyxr5cmEjgSFRO+pi5gB+rAPd2dS85Slw4oUAO2OMueHlBm6
lxtlNl6ChkFixUIMtHVul2jeVRVwmGCT1iQ+uFaTnZSnPD2JtLjlSdiM1BJZZBwb
1jpzJph8VePiHJsBA7+JNOY9BY6hR+X+EA5ftR9ZPmemXibkiNy5yUWPkuK3qCcS
dx3beVln+O4gbrRHOpYMZ9gF7/j6z5XDwgiC+85g2MyWcrcQ2YREaJFUgwm9etFZ
LoaFtqCNQA+edfZ1r7k/4f7oeyOMDCqa0YoLRSS84Sl7sZeUhlP3IGXciKlnQ9VG
ByX+efOl82Y9/AWHA5xpuWR1ojcS2NmJPvziXBAClh3ngBvG+eKSQUvaFHGxUoz4
ImhQAYClo0jWTb4VmjjIz+nZsFSbEauSGW0UL3B+yUMWpdxXcUrt1dU7qs/1IZY9
6dhMtM2/m/aAxAYfAvuac9QlsumuPNhOucAP3lYzOFhY+I0aKmTEziOgd+U/3YyX
883CBaC/1NIsrw93BqJCaj6LU78blLoDe0o1Qc0hFSXILqsLuMqRmsgM2DgfvDuD
C1Go30GsuKU2YLLx0kDzWW+SDjbWBBQcIPF6ryvx50JO+2ffeW3FKOfw/Y8Pc03v
nJOhX2kX4Eu75ThzNuRd1Di2UV4xmstP2emI2Tsz5OCgeCT/TJCY88P9JP2XQUmK
Hw3y5Soy1vVg8wjrVcslLQxbxj7uQKB+LEMI8I6yOOdaL5+MkLgyaZFHYj3bNLPB
3tgt5nnmuqzNsUZhgPycWcnVbZQj7RRTaqRqRNJmyyxGkO0ieddPUuDwNH2tBgRw
TGGw4C2vaWkbLEjYpLDKnsXkED3+FRZbPpc0IxqRcjLYlJ/A+oUcyFrZHCI+Blbf
6w4RrljQll+kZX16bP/3wer83xGBvv4hpV4JPhNaoTNOkUYJjrxnAZJWwoQ96qJu
F2mg6nGlrDQPEx0TZiALoi2Vc17KhhLJxLQ3gB57n7KjY9LOHpEY9zYl9pYnVvNz
es8NPxP9iuHwf8FV0hyOLHe2HClo8gOB7ZS2fsQDRLuFoL+kYHFVbuPsazlhT4gd
tQs4mq1fak7sgNqvB4srHgxTJPeI39MaCuNfzy5M9JsfimvPyA4saiA/z9ZkF1pJ
8wnHZoduN2fHC9jgM4F+yVhlFHaIwHxelLPxPlwhfkMkWY6EI8h8AUVz1YvCh3EB
F9prUmfVxln4eK7CRyLJsL1Df+rO7gYc0jlA05xL1wLCCyB/coW+o1n9iQG9fRA9
jLLQszUA1vu9Z1YMyGcc1IiyeJM2sni1PudU9kp9kVFsy/XsaM9H3kcgOtzq6w5t
wHgqmtm1X+8H9OCuE/FQFeQji30gaT20EhZZyMAQCK8nBfuKGBGi7KXa2cigOe4g
woQDc9kFHb8FcM6jAPhkA/VJRrGjSp/P9zZPQ76M2vhpaWmYsOY1P/MZS8p/sVkh
gi2N3EXHKl7PUXmOaF37f8qwaqBAhBz21PYA/p70g4qtNvPFdQ5cPPpd/111j+SI
LC7cOPBbqF8nbycQhdYq5DytZ51qOTi4gHs0BBB57AtOoE57mz7y9r4C1AfcePcn
amgnlTAHeda9A5acp36FwWhCkhL5YN9MhTcZVBtCWvprNT5YoAIk7pPoC3VlduyH
JFj/26C4WXp++KgMECQNYvUnLerJtV0zTMVdpE9A8KtXlvpUdv9G6XzxVvErrpQC
FzYBXKvHiZ/X4hzog0LfuaGbxgqqT46jT5B+pppnArXTnLSe20/qNUVTHAKkfRUx
Yh6vNq1RcW/IbFD2B1KIEQVNP9kLRzGKd+8mjp5M+qVJsxx5Cis2CFzDhWgpdlbp
72oFyFtHE5VMvffHQaCRLBrom6dz+T1nMullNWueI32JxyHLrVfsjSOcikOXNgDy
Ce3kVtqVvDJOb6ebXJ+8sdmbOJNtBkS8bpZCaEWRG1x5AN5VXREWBy7LtrDCV+5D
7Q7yWzWpEyDMxWsfEpIfaA3fKaimiiiLhBEKhaGf8Y3/EbcJSJ4ZS8KI6I7V6eKB
vkjBaIkva6tEp3DYZ5XKtSlIK/aeYw0VyY97RZA8MwsnpFQVCzllO0AjqC24ppmc
v0epoaADKzWJagJbB9yo3soSefkr8GxK7iTaxJvbOwCBRvdW04lXb9o3dQJ32Qtm
/pbQrPEuGIYKqHH3it2sxM6j19Zd0CXtyQqoj5j66i8zPS444jXPPT9r2Mt+og/Q
pgIZtkxLF06EsvrTIg8yBKE11Kr5JWmVrkXrvUISfOOcus5aHPbWxs6XlR2Aqek0
UaLwx3WX/wxAitHNRaKS6pNTMc57Zl9naXPP0RhJfQbKn1HWtNUeF/lOITILjYy1
l+d7rA0jIZE8iut+YHlpLb8lKLOL6aPrUcSqs3IEDZLPXytGhIRe9EptvTDqZPbN
MAs8gj1GNW6x+pReNvE24+UDYEt1uM4ARI8aReRpZ4ob91DojTNOMfYP0sWL0JT1
0/Hs89fwSOhNSc09tmpRG+WKaSuj9mchLAQHxo4mXqO68quYlTBUdIWm4cdmp6DW
NOmAMWUo9X9yP5xrMJXc85S4Ybq6FLThlu05QMt96ilJ5NmjSWC3sCSL+66eyYdr
AK7sHKC1zTpEn16OT6vZUsh05z0yOJDKIKh4m9z/G+1aRf1i/Krc+XPfTtkfuNg5
BwUtTnPuGbRqGMPBqWlBRPlyiHzItYPjBaII5Rqf1l/IZlOTuQYSFunYzfdsG0d3
QZ1zEM5ul3vuX3F4bY5wGHlCZsrjU1E67fFni7+uiJauZ5RrKnhzWV+cmGWC1K+j
szqPy4nx/cMZ1FSqnUuxSPborc/ojkRz8qO1WD+l4o7MfkNyBZxNiMMkW3hHigmY
3NeINUVehu+SqmCYyiwAlMf7hmMUx7K5oN0FxlXVHmiM5u6hAoIwBqUDTWN9VF3T
OwWYVzB2SP/cXZ7UOQ6wkP272bKQMEFEAiwx/pFEObYu0iRLG160fDhMwGBracVS
2bd9uVUaqqrNwja9rAcyvqvBGm46ZTSAI4MZn5BQAyKZP3dABZZ+8AO2J+EoM3t5
gedyYVBz/RECgHNetC6C21wl7dktrPmbFmQOLoYu7VCIFr+pUjzCeq3KGW/57+yK
RH3jlP3TkNQYkg3J3lgD/6JO7beG9g0FQoLjIQQVNpAVasm1BaSavEy1iHD0Cyds
GLVduQMmSXo0eMyHt9y/PUI/VzqoGKoKhAe2zJzVCJPCRy1jPtOTg4FfdnFqQPFU
JaRpZq7C7v7F0pzV/jH39TT3nmQ7Kw+ZQYMzYlEQp88tab8WBJUELUoZQTcrz+pM
Wo0FEFN0vJ8Hm6ITXXKFReAbt+Rp4Wi0hpQda9zyY5NG427ch700Uk+QQoTJhU8P
EEHopG+lxm23VWahvF8E/Xg2JJcTW04TmsnMOX6sU0T3Ox/2Kwh4VWYhK0y5+ghe
bqoZI9AOtiPKMndnOIsaLZlGJ5+XaAPs81mQjT+O5IUa9Q9bYxytqBEaGec5X3Bj
8Iq3ClAlmJUWRfOxagk39y37dBm6WyYG4XbnU5mp7VOUcM/hPA/MOV4DXbqnrNzU
HwF/YHDxcjp48uY1szudltt6iGKqDz34Oux4eUIUjS2jNYDtng/pnu8wuSautBrc
GWFmiY1pJAaOh/bQhj9ntFlUOIDw+fJncQOENvhFiic5l39WPD+ajcuknf80ehq0
I7UDzRCRsnwpI2C7VkC/w4uQlrwGvLiAt9q7qX/GZGmuNLOgc5cyjJWguVcnO89H
WEbRbw6bIRyMKliKvNwJ1TuMeOhD1lXJSj8SYSuwaLFNmpdE2Dw8PCB8tDXnAhsi
yi9m/dbddm9Jk6Muesr0LYoXEufhnpubYLs+4eLnIBpj3k9WrICP9+ahy5xqDCng
O4LShJkGCbdX+MbQ964Zyt2Yw3HdMZYq6fuAC9ROWAvkvMfkarWWWmSPdZ3KMtc+
BLnxES6ta4G/rAKAmF3vI82QPpL7VGqSD8Ywon5bAg6hs+P8xl69OSWwSOvf95mv
+PiGehvH8C08X+S4JFl4sSV1jW9GU76LG2Pr0+7gFVKuut/Ne221MKp7h8eFb5de
cgoAf7iXuBhf6w1yUb/SsBxPMSmE01QFviDac8xntVnkmQUHkZ35MkWCYDy9TFbE
npGrwC0H37lltX+xOfWnDaPWaG25UdhMubgiM2tlISca7qbQRYNmSTxwhZOJtOB5
FODucZUZZbY5DOhu6TU+a14k9SivkgrmHppkqaACgr1ds4d2q28Zwm9BTzXhfOPh
+vnHvLHoCF/6bfwPuIy0y94AGs3eQrqkGf2PoWOenWOAAkmF77Lq7L6+NoESp3a7
gRNPRCtX66LSQDng4GH4gfBIkCNOGdMP8vHesMpgBpx6/GkKejzbwnRkft+ScAzK
4Q1utCRzEgJvCdOE1wARE1szer31nsLa8zKR+5st1tHIngI3fzaT5uaQApTg/gSg
dM9Fv64Xw0ss3UnFFYF8b85rHMt/oCyWsWzlguDyeSpUdusjKLUw5d7wMb3cKT+6
f414I4lLcJEPbUtl2F9fK0fgqY6EKeuca3LXJm+LoYjUI3uZw2CYwxNY84YJI4wu
oiOJPAbfFwLUFNFXz4IYAYGnrndj2NJ2ncJ38KDHYeueO44/WhnNKuzx+W3tHG5Y
8b/o2oaJvN+Ax1P9UOxH4sRq83KFfAkYf91bW45H8zSN3w/u6QWWnaPAiRkUKd3y
GCyVKBE9A+Fb6jRPL2vVZhx3ar2RA6/iDTxQDMuPd/9SexcF7UWYWmZZ+/5SmjdB
wQ1tvsgvN8H69u/HCydXgDBPIzn04M7blyuFONQO2Q+5JcLCSlmT0CEc/74B94qg
r5t8wgtB3SfLoRo5rGNb0+AlUrCDuaEXekpU53HfITmyVJC3/GYMnplU97uxddh/
0qlODjt7v/VPlvBZDoiXa2tRzUAd5gk/o7vtdOlq1SYZDAqr+RDaAHm8OLja/4oP
2+mU8mX5waNBCzlK2YzflCf1UitbaZhxmPAwWmWR69WM/IGAaNGbFnEzQL2wS3gv
QjVAN2tmuez/hd2RaYVcgnS+rTK0b8T/zLBkN9OL3X1KcP3s9kPD0pk92hMpXv7M
1/wCc4lavqODg9LzBVQdZ3emI13Dj6JDV/UcPytvU4R0pOCAFS8Xe4Hr4iSxomQg
t/ATPmFWHZFUcH5OvM8QwKnFGVfDa8PMIIU/hkFRk9A6fDluTn75vLRTO5Wrg8cJ
UOfPDgztgVnxjmP+YcwUm9G7pzPs7gGJ8wqjZLHNIcx3yAQIzBV7ny1OqaN1SUdn
b/s3PESIGntWQw2WH0TPjPT+Ubl2/Z1JmDzsEhrBTvtT2ipqTnaAtN4i+Gk65GEf
KF/53ZehvtsuAH1bSG0Q0EcOxwsHENCep2d3llC/4bJgiM2NZeSDOwZMf761Uqy2
AUlEyhaZZmBkqQYAGTRxQULttqZV8sZfKAfrdCY5aYHYuHukZeaWuseiAFw+J1ZN
oPZtEN6BIgjsg/NErCCB4SlX+1eZlEbrJmQgUX64o9PEUISJM5t3mHBxs7guNFJl
uQkqQS2wE01g0CPkTvIYdLqFKO2um4hmW/vyZtwUEJX1ouimAGB7wDNk22iS5cs4
Zz2elh9SV7DlcoYU2l4R7QusWggiOU05ouQZAqTHbCjd9DugVtNkC6rxaNyiQfGn
IrBLulo4lAF+1pCak6ZTFH1pNwg8hyaXm/jYlTHMIo/JjUVNiTZEhX3zxb3ZwXkJ
5twuZZNNBtk6iHZA5b5n9ceE9KVRi2ZN6YExfL6EHSkWol3pQ4GrRwKpU1/wTKXv
OY4HuiVJ4qBOrXlkk8L0VdsdAJjIjPJy+lgySYmO8Ux+Azrfjpt8brl8t2kdamOS
eCFZO+sX8ZS9xVOrbcyRmvSHjhUyeD+SBkCVURqEYuxFgRJSkMHc7m6Z3T7QoHN3
/VtnWW23thFgG8eraXL+OuK+/oZmrrWf4MF5jJSxOstiTSbbqBs8jpfDEuTYWLJh
7t0FNt9r3DJ8B4NiMmbhkgObbV9YmvXGYRF0ScF3Z+VW6axcsz4RX46buvmx5Sg1
Y5uJjCtMxyYSMM9PIseMrLCSUMcces+fdeTa7htKRQgXGqXoqRq4rN6zT7lqUsKz
aCOqSFFqb31Aya3bMqRogoF5FHKHNWBJPdWldQaz50KmLEv6IPaBksLdR6RqEVG0
qGHKi/21PzgoBYn6QDyJjJXbWrvuJjW3Z3bpSsZskuxgamo3/fCy9TxpfrBHBPv1
HPnS9ePGv1aNVOxF5agX4ZMp9UtIMhKE5/zteMadjt3N4fpCSvJDuQl/Y7CNloxi
h6bsGYUzWGW5GrQqc4dO7hlwmtRKOfm6/wsqtp41aqhltimOSM3YoKuO8bIZdeUu
A8771rj7mi+Cg6BG/OrFw+SPuOqKg06ddRv+L4dy9+o4nfNGpMfGOAkTX/5FxzRP
yv5QwT99dSkFSX3KvHJSBlKyw1GjiqM5+i0KO3PjzFfoxDfHqaLgnb9iqV8EdFj4
sUqpWz1J6r0ITYS9ZIA1J8dXaDWHzVpji9WOaxrRBlAr4cS2O1I1Hqp7jBAYS1ok
54++AoRYhXvOLjpP/Lpq+LitWTAVTKZ2l1C2KR0pt3Szlaf0DKoEcIvPQfFNlFP+
jaypi0kIDnVw19PN3KW+GwcbUy1QrwlAJImrkdUsUiEHZHS1gblqfeDQQHmSH7IB
G0ERL/xNGKnNmJHyiSwrULWt/2aiYELjA6u592cZ/r3HMiwe6CQhfTwoHoIsTcpL
UVPLrCSzki227aRXRxOvmn3EaqHPMJMco94lgMjpxk+f0kgtjh1WJ83sy8Uw6eGv
LMYvfo5jDuJ/WjLtSXXBpxO/I7oKC8gRwzXuQldwSU113zy8SP0c7x9EiVgmlzNz
v5KuX+dJj9XIFyjoZN4ZBcHnyAcE3ST8UqTSHJE0OR66mSbBBJI7uT6HPy8YPSfX
IrGho7ytenohtGJfafysT0HLoOSAtbNHMFJeG6hb3FbF2O9MOgJnjy3WtcBxnPmG
Bi34KbNuxC+zirYrau96W3T1CMaDCXyjA5YS6uiKJGVFIUVemyFVEP+n38yRVdZM
l14ZcUbXE0DRAzSJz2rSc/OkpakGiTiU5YoMFr0DQ0dab36i3u8YS8xV4Gudh0S/
Z6dTBcaVeVJbQOoTwBlC5zfLididCK7euJUf6yAq3Ys+69ymWhSv+xBfE2/mlznG
MR+OMQi0/CasP4KpOVzoU/JKvd6kVH6Lb2nxQHyw2h3R1gDVTkgdikPzHZ+p4alm
yULrgD9OHWvGQOEzm4xr84Way0YjBNkCI6dg3alH6W3SbSTjqiW7B6/gMeLSh+n3
3x3GKdYU8PGMISKAci/rOGPVjVR1Rm69LJPAQiD4ZW3ga3TtBpjUaD2WByJiq30I
QB+1QOHGxF9wfizlNro2j+eQKFtJ1TGbGWldk0FBImS9jJFyv/DMOtBTiTfI0q9n
pMUe7Dfz3YBxI55oxI/Y59D4x8v9QNO1onGZGwQwAJJQHo07JqlKPy4A4QNK0nuw
ljxM5H9oPSndWz6J4hxixwbbS627590BVIs0KbbzorDsLPhG55+iHKXRGi7rrrnn
2QUpkm7gDW84rm/QOR5iCbpQsm9MV4NVIXBZkqyL/6UIlG6PrCGgPH2ehxjOGq8P
b+ZPE946Wfaylw0gAITwrE74ivJheX4F4KfZEVKtZ5VlTTFX9J0fVrFhckAaUwhk
CTE7szZQJC0hXC8Avk0+gSoq6+sLOcrduwGmFf2CX0kZ+qtkt/UvlX++tgOwGPXt
pA3IDGHRY56Ivs/mDZ9SUF2ngR5t38/WdR1aMXJsKaTZ2+9uL0BFBAt5trGmTF14
IRlvxLI5b5r8JP0B2mYsnRngl2D8dMYHzIx2+Tth5S9A5ZTIonppXIzyMCtzNUe7
prxpdp/kyyjlqNUlnvSBm51kAChbeNJ4IBnPDO+X17dw7nOJp+QNOMhFzG1oWkZf
PB7+qERPl/nRQoeHjOKVrUSxqabbNJMuNCmlVo3hY8K404iQ8mLZqib4cBgZ/hWX
ceTlse9fcbLI9RgApa2GGcatpEYPOKu1r/DyO/OLLKJzZRruqHqA0pNbFm4F/lkN
A2hybJrar6egZHK4dZYqmCEuhjyd0WuBdziDy4kbLzNp9JEHkrTvmGhAo39+ryHN
zt7DJlNgZMMWi1nJhX+Ao6FvkCzARjjvlGq2lHIBUG8GrzcjlDG6V5uUsvHMm0iK
7f3Iw66dkrH3ucuIOX5gw2UdHOofKZ9ij6234BT3l1LCAxTzftYdLpLW8JfWoZr0
6dvs6oAGTw6zCiu9iOLAr4kh3a0xIEe1CCfjwBVjUu3YS1orBMEO7+Barsfc4+VG
Ktd+abXFGv03JiLcqMTGFi3elcc866eBLiqocKMojCfQzFi3b7H2M0XNbHcmyWzI
TO7A+KUHQ2Ajz6zsdQu6yNw5X8ywzgh7ZSy3PsGbq1XF2prelOhtKMmIih3hXnFo
ovR30R6eRv78DiiggVjC8Wvy39D5PGhL6qpr8CLmoSA0lcGFxIoTiWqt33v/j1Af
Myqw3Zruf1SXyBDpleox7uWBtNRotujWR05OeuUysNS8RPTLW0EVhH+BK4nXaSAN
dUdRag6DA/xXujpM5EbLTfAOAzofhedrVWe3BUxQ1/c4G9lDUuVEMQyl0obQZ9wJ
0T4eHV+ZM0nzhmCW9eeLCpIwATsX2+8SEQf+bUzQl6DehoO2KwBXWdBvHd7lEmvH
WvvS3aT35B34+zJSdNKGCfU2M9MS8ZDKmmCeLZwoYTc/C9cHbQOY6vlZt8JPohuG
di4AFa41d5VQVdpqycrYTl7lb1GyT/lo374nfV4h1JkHS9bBYFPVMgaRpRZK8lHg
17jTokenssZkFCTSer2xMpOv6K7p6Fh83VlJL/hnmPQ4FApbkSJs9H0mEDRzxdb0
03+hlsLQawD8FENWK7Gs3K+tJQR2tv9bgjl/+K2pQ2i2QuPKbxuk4PatcWwTpXsQ
H3Us0wsVwXz6zCMvnsAJWRwoCNxkpBpnupH+ehV2A+OIZENRV7BgyujxjsKZSGPZ
icwsIslTLOTwsQsBhssevqlVHtj6qxXyDSe2ArqG+2R9L+ToG16EULiSvxPvOuen
edKWdxGkUlydu3dDAvlC1lZMNlxKhF5lk/ikkb4incilCgZyyG7vot0hdRahE+3o
VUMMzHceOHNasi5PEq7NZWk7pdVJpq2HXgda66239Vq8OIejiS2HG6011mffaHfS
hV3G5pT8bj5F9UqIYhzMC+Y+E4RWLN2iVmAlLsEpxoV5q5xFp9yVVMjozLxG935g
E04BL9apGYkVjxfRuBVn2/Ts5uWidJ2enZrASEBumtZuNI41dznNHHvX/vE16Kda
SpY37CpozzAcnI+teeHKASoBhnLSRc70Qab9VHa2Wdw5QRmiX+wx+55cKDJ+fjj9
55jzRUG68xytkD7xnB0S1Pbj282p623v6yrO27JXvuDHqBudwm5i4Wy0OtGmrgIW
CGBDsVBoh58eQzhVMVHj4Fo5gyMcjLMob9gK78TgJAyDMb2xpwa/peB+BNKGrw52
UBhJc32sZ2rKiNLZpb5Pe05oXLEDdzXm6dDgqyl1cTOwckPnbJqXbmHTzFhrMfnO
kFhGWtciumK3MFPWiK6ENs7Q+DC08/Vy3c1yXzOADQgFNusaXpTp5N5FVfgl0o35
D5Xc25SePvFQHm1x+3kbObfL//M+IOWq8oSVyn5fU6Ng/agjwqpbIK5bLsiGFOkT
vw0PCcU5kdNbJllmvnSmZX8kMbsL2dy0gE4o4SvOp1Hnp1DMaife26AizfxWkVxG
5NvgpU6TJIjPwbMhZ5sVxy6MdSELmCTZKKIrs5khVw5I3clxcioY0D2ZaSobfTew
BP5XKsaVw7ChvUsXtc4JjVsGzU2RtAg70vnlf0nmcsLfUb1tGvxoBqsoerGfzBcl
uRTvMs2oLpYt/hqAXOScU58xycRF2UisDbtC4f/VyW7AU1ISbQEu0J10GWKbORUj
UdRLP2nbdY3D4pyr9U8ecbuyNZ8l+CECi8+qv95LYKP0dU6IL/UHlB5x5r9HLORy
hP3QPlCDaUNS8mjnKWa5q8yOoYEsbU82e+ptEwTZPyDXsZmleEm0uWy0BukIgMrr
s63wv/iDD3yMLWfg9dVSD8t0gr88GZQmtDGTr7tp7JdhdMojxMGlAZlbQFq3vxVi
D0aa2EKNxEAEjFziOGvC4fb92uwQMH5h9d9W6kW9jy/u1/NkGK2YBW5bZmdwa3/n
zHptA7XZgXY6P/89hNghT8j08Q2FmW9Czm8xYqMnjcRydgy1nsW4ll71E3QhTQCC
LMiy2Xcp2CW6Szi8Kemzz59wyQi7HtmAtvvNATLxaJmCIraBSuC7Ia9mYVQ31Ub2
zDVczydKK6wVVrCS1yeSEkPiijk1yPpBSSskPi34LIj+4oRgXBHsYiw/6lWve70e
5Gnqhpld+0r7iSfpclz5tUFF5yfRXQgdje4LNuuPyHG9N+nyBimptk30GOJMc4hG
d/cxtDXOirwbAb8PPQu32ZDhkjV786zKybg+7jzukj75Et4k9VE9I9Y76tNvY31c
4m3kzQIiaYfmgXg/54aL5Gq8Il/fGtAIPZsNLqN0VmRnWJmRV7apomP6nEy4n6s1
22B8euMcpTXUrOXhTsITXLK69sXfmp3O9rAWReY+O30PlvwQ8wT8IU73V6iL3fQO
S7j8nx0NRt+wy/+YKqVMGTuQB9UbSBiB4p2IA/OTjWmKUqzD5bc9bOmgisPTf1Q2
FWgkjTHEi7Rwg6woQxLerZRH+K2hMqwNrA6cRbT4UHVaZ3AX2TifoSyLFsHbAVc5
0uwK4P4JORqBKsIWtBco0sFw4Ez/ajng6f+RuozXJWpa/v1mPJl3W8j9h/J6i/5K
FEPwqnTQUEZ36+U9QxMKwMZpnJvtG59aALEpBtyiZKamFFTpXeHolqyQHlw2NuT6
1f+U9KOo9ZSDwdXt/nBFPCNTLp1HfWcsF+G18H7KRKdh0mAYtf2lROt5kfRHHuEw
SkyyQGkGXPahiL/E/Gyw2iwBbbKooYh7yS9cefzjaPekoPe/NOuTVgxdsd6lWWOe
rilt69G/66equ2KyODPprzEPocyowmjHkW1qVMBM83Bw0D3eLbx99cU+e9Ic+/Um
Ev4E8ZIk2rR83B7Wq2Hht2M6deUfZD9ixBmMdzNvwlX3ehnCQ0IkP773ERZwFncW
I0f/qVXUjHoW8uD2G3EazPlLjP0t2dZMaAXuG4pH7MpIgiNmPVfSEGJBCiomxKKG
7hVa9QFBHATNYYwL2lLcIyV+mQe3vvxUVkaHC8VlDfxcaBag/HJpYALTHwdU1jVo
GkwUWU39ivqQ8PH2U5gZmS6w6QGE454W4R44PQIneQEnNnyFOhi6ukwj/2dxb/f1
hQuAj7P/zIAnjodhASu8UgbVHCSu29GrUlJSyBNsPOmsRYDf1mvJ1QHm6Y7CyQkb
jE7K9M2kdaxe3E+7AzQIn3z/aKKqupbzY+WMvSaJWycl4fZMbdIUGmMMl/PQnatr
abkZ1QKtgWpwMz8iG1+AKw+vDVVlfABvfQJ+8+IVWgo98l0IlcRnHJTcwZ5l0vO/
lSuNo+RuYrcgXnvxOYYOZetgQRFJwimGhRMs1KofU/a1POrrmJFbAIrlzWosy07X
OeVhSPZhbeXC+cFF7WwAgmlGGOHV78dBl+9GsXJgx1OKlVAY3bY0MaOdUCqZNQWH
hx3fr1c6WRJA/DVCs8jOvlDU9SqpyPrQfPAD6gp4b57d3f+ijcrmM7ZsXRHe91O5
TkHRsmMwM4T/xkiOOldRSvPBbRfki9gNWyboLDtuPvfWghm1w98/S+8siJrXKPoZ
aObRDmzorxxw8iILZzaLtbeYrvjMjBvEwqm/LU0j5DAtn+KSmIPhy6IVNz+ZRjyj
yRU/Wrs4FPtEth7o2IkQ+HEvx1+QxyK2xIe1iWoqip9DT7nfn2HnSFKT6Z2VoyWr
AJfik9XGLoaJwe1ICLBDta8P68qV4DLWIMRTSFQLzbNoIxcDaGrLVppHxRUR3ej/
ltKvhwekC5sI+RnCgXgs8E8thbq69aUEnq/7ULvHbYBg7/t/mZluP0EoMwQIjV52
JqzudbC5zLr3PbGLXIuKTbMU6CoMqOotru4/+iVVBQWbZZKYmIxQVAruus8z/0bh
f27iMm3vK2WyH0WFkGJWIhIW0mtBM6KheXLY6b8y1Ph+jISR4v/K48SmqgS7hrmn
M08dDfml8ozm8PjBcyt1tfIMvTch3qHdJxQITsSNaBijtSCONSmgWhLzm77YLJj+
c8jdQ1Dtu8ORvb1U3P/8hFC2aYKc8sdZcGzLyksJ0NQewuQl6IJ6pjeK9ZA4u4gS
ZkDICVgxTBtLvRYabA1d0v7IGEu7aj4p3d47miMcvDQY/j1bVkVSm1JYvs0TtmgZ
4oT1K69vgmdO1QwqzNIFHUfw5RwGTDDuCCKvgCjFmV4NVugyP933YQAYUtCjeoT+
qje8KChKe+jScunotH1nAnP0tBljd67kqDoedVbSEd/9Ii2isaSZipmqEHOh3XRj
zgNHeT3xXHqO3M31gytVNMlZuJV4AuJkGXSOFiPLZl7zUtyT/uLXP/4YjSwvvP2E
pax0LRt+wYpjQ51Y4UyHsme/abyMkNyH6FQ/QR6H79G6g2C1a3oY2yVJqIRHpiqn
MGa5VReI77mOnyF5XlX1uOpM3SFlZDmTnvxnWnDBDSQ8VqOC8izo98JA/s17AnY2
vEx6obRTjnKppKZhWkI3OXO1MpSXLUTSNeTg3wzH3GiUFVp/3ZTeqidFXK+uhkyl
ycUW5nEj7AidwVi0OAafpcyVauJ15a3HBxT8+MM/JeOouLVyV11XRHMaQuTtGao8
JnUlR8FISNf9F282htYSgdQ3tPRTGf2xf9cmax/I1pe37AzDUmlwNcpkK7p6gBBR
XqVxUiB7MrVGChU7M0xpEFx5VPoJTC15kDdMs5mGzeqUl+S08somP8TTD3y91rGl
QoXU/XOHg+35vL5lP1yIvPrY/vPlyXleLndoK/5Ca12om5O1wZ6Lr46EQjFSsSz9
iq0h+KZmiqsWGFhfe+lEdmQPUxxoDke1Z3Q3J8FG07vR+D2r5sl4HsQmJoCOFIEn
A1dZf5Dv7/Njm1jrIDJ4+Cv5Mz6b/9XEnEJ9MJLyYuhIuuKH3Pyv4aA9umG/7BCr
nrOuNXh8G3cx792nU49TcM3epaYiA3lYAPsYqSUliz2O9RDd5ZP2bVM+50IGxSSw
WUV1l+jEgxcQsfMZiCAPLBzfq76tD8zF0oA3sAR4yur4NJR805GWZAi4OtMsXhs6
+MP2WzoHPvajuYDfU9uJ+sC9vVHXWa+tCihwmz/05Q3jbPeEwXtwJQDuLq2UzNam
f1YeiZZ0cZZdRFNSW/G5alFXssitUlYC6SDLBeWU6LGibgOm6I7GzEANVhQsKcU3
25oLwQ+6Ayo0wdNdUOnJJeDYlL+ad5xwLHH8ead8XdSjnj13pUU2ixAVjFivJEod
stnIpS4esPe6MCcjTTR1dl8TBKIA57KipbbycDIxSREij/rZuxPGLnu48sUI++s3
FVl9FYItRCNZmED+Q8gFpIXQhQrlDxcEJ7u8K/Mgd8mFf5y3kXqRpkJKirhjU4lX
xV61Nb0zEHQKWI18EAzrVemxSGDoD9L+ZqxJOxi2keiiFZZdMoYtJIZX+6i167y1
XII2xo4u+q5VpTBfhwHuOWP+tzmttIXPEZCynN8Ro2dJ7WIWGiNiAt/W3eAZLrQd
s1hpC1USQ1qN0soRnukEDI4riFp9uMHEhbLK3U7z7ZLELOGTILV9zDsgBb2bqBTH
3q8k6yTa1sX78fxGa1BhYvYmC6Bm5e8mN/RBXAiI860zy7grSdNG7Yy/fGe673/o
0T3Xnb1ZH8ylOPsm1V5v/GjfyI7ZY9nuB8KaCNgzoaek3+4JoH2Jh5UCRjyTuyAG
oqfws9VOLgIRmZRIqoDfDpdsyHxd+4+psXMudkHfJ0eTtnnxemx69o8PPkYyy5hH
je+zRfPqeXkM+6cY4VwOac+Yn9Er4x1LixcGA9ITAXwlNI6qtGyJK1+94hPIMSd5
fciTMjO/wgdvvixd8eoFRPeO7MapOaIK3CTUkqr5EH4lPCO30F+PZuBnwwl+bgZR
sOfUUgfUN9SPJ8WCaxwuuj/O9yAAINVFNz7ENAd2bE51RlNqUqKy9TrosRtdSeOT
0frSE0Ee/CJ7iSRdvT/eQKR9/k3VMy2yyOeE200Kln8NGJKKERabrKGC7XQd/MUB
4JY71rExDJq/72Sw17sFCqgnVvYvJss1pnUjVkLxp/KyVsXfR1x5SrZcc7sgEsrz
zjnsCpZRdVhtk6MZ/5jQLQudRQR3R0VTdDjlBYG0041hz4IEppQCA0bFR1N3Fm9h
7CQTdkWgi7eAD01EeRZMdr39em3EcssgwnpretZatZpe+DZXs/L14Vm6nR1gPmNU
doRVbV0wls9L5a+HmHHsyDULrnM5Z1xhLdhHx4ipyw5TCdfk7jkpyRY/OwSpqrYJ
nYGZCOMYWoRQs2f8R2Ki9T2QctLF688i8qBbCVX7f7MaZTVsYofVo3uUWBsgzbWJ
znPp+LnjA7Dw3ctdpUJp/DpPmZ2ByUHUT5zYdftVs+6N4LEsN3/z8pQWAeCIPtkK
wMcKYKkpZT0fF/6m2LuGsAHZfl5NRuDN6y6MTrEDaCGQRZ2i6/QqKqeMZH7Pvx5N
Xy1TRA6EQLYJLP66klgzXaC5VdGqY2JwMfaH8Hmcl1AdIqBSZRxAqMbU/WJmBPTd
5IYptKeGc5ZF6jbKMA7JS2fMkA8+K3aaN3RzvKZw9BQs3blR1b1jJ/jURrLd9x4k
FYvrCVxLjY+QO5mMVFneysBjJSnOboRfjlm81FDn1lWrJDdp475yB8XysJ7WyRWB
o0oPvNiwnDUlnKu/96l4bXYk83g6mzC/QmHX3hIia7U67vM8XHKpZ9Sqz7Bis2cF
xJp00Fouy5v7kngozA3/9Y3AYLVVW3Y8g4/0nIPi3fpVPEBaHenILeXeAS76QSXC
HukCVAx+h3SCo3taSGHytVmJkIwTuIYqAgpV/kT+mOFN50POKWWBD/g1ArjkKyGn
S2G08JTVojVV81s2Uj/tSm8Ok5aA6JBPJxHbLy2ChQDBjO0Pcda407e1HXTgpcHW
3EBb/W0h5oUSler0Wzz6mPidXjV83qsrPrW7BdkwygHUUR3G5AU53Zq84qxjlMGK
ZNyeMDZ5I2+zt3vN2NgNL5hKUhSfHaapFXjKLfmeqzpJMnoJQC0xJzgo8c+heb3x
QVlh2mWUDhu9dT0VQWnSrwMgM8nT7LufE31mzuLh6r2xGQ8a1vuHF6lMG+uffvmI
CztMPhpTMETpLt7M3POvf3q6rB/Y7XWN7LN+nXJEkkAC5a2YMkspZUqNjclcvakL
er7TJNAcSj7znpyNtmjiEgASHJeSWhLw5ei/Z8fdHywSOz0rvf0LVHRPNHOBSAB3
cQSPADFHcy0iTFpREmTgRl9Mo1t0tUPvauQfey75yksrMrws5yXsGzPVrusn+iiP
+kY2aRKEsYyqO0hUWd8Ed8X0+cUJBh5xM8bJfNdyL+aR8Gsh6Ynkb/fu5ahSIIrC
fY46VvsYy6YUGUhpdAAz6JJhA72VmMKaylbQN+0jrwWx85TghpA5nkr13dXw1kkW
beXhWtBs5VgBzeXP1wtkTNC7y942d/UJ0zUQh3DPnDKKyrMbSNJy9CxppHc5vk9e
xE/A7+d82E56ks5k35UmCdauc6qVc+ysm+bJ1/B8KpuFTNOZy4rJD6ZW8HeoknWV
YVvhEra+Ybi5Xf+Try0qyQbfnengxyHtXmBkc8GIYtofLo0jFlxpgMQo1eZ4NqCj
ZaM+O4Zl6LwkTtJuV9x93JC1ublW3ZXYmjmof0xe0nVULoxGc9Dxdcst4RDGPUa0
CB4PihrT3P/ZHOJgTOi3x+D6OE1YOQtE5WSnPV2HuXAeSYjMjfz5WCzWHotUu8Yr
UBD4E4LzHr9IWdzOn7fK+9Dk2EvlNKi5kw/Gr+p1dclYSML7eLM1QOOky9yjVtac
K04fkP42qaNuZPyk7zTkdUrc/nBl19kLJk0hje0+bU6vSo8/MA0D9R4Yb78SkPO0
Vlx6fFvYVzslhEBzBdiBp2qUvmgnVlS511eDCnl11mH+wewnab/Pf+lT8RHogp+l
9gVA4ROPrZdgoe9Yg0kcHy5D2dp6DCalaUndHXjgh25pD+j7pAnG8hHb9dnUEx4/
Q+UVZ+/nayiJERVLrBVqCaB0yXKI839qwxdEaE2FJk4hpq0Mc2Wf6xgT0sdSGaQ3
74XZC4Ji2qHkyrjbBeCJ0YiUjZzdm3VZzywpLVXiSPai5MBWLAEAlmEnNhBfBQ1L
IgRiYMRkORqx52xk6CUloueULsaMOKp6RAlz6iUcPJv3tdUfTs6JgyfAvlCFEnSx
oLrh2H4ZAiAbE1LaBLCMyrpSMdDo8D5DsIDx+T5tM144/6jv14xSfjjAxHaXtLhO
mtKsZXDtSlkvvI3Px25wOKjf2a9QOASU8OA9kMu2nQXPihu+mp/87DVUBl09y0II
tcjqJp0TZevnNHMlKGKJJiazmqDro7R4ei9zvtLlkitatpwprlnM7GyC03vBqc1X
gbqMbq6jdfqvfYOi4+zd6tgyUrVnKpEGtP/EhGmWgHNXKrso4eRcy9h08xLeJMKl
5cUTXzQoqLHMyDjRJKU6P8xj+b7pKcxoEZFCg4loByVpk8wyFTB6KOJ+uLnUtkLU
KNjj9L/nJOVxd5zk57C6syko73ZE+YG4P9xVbtpjSJ9WUHCqQfLGUlilwf6rJwYD
bGhD+F+MnJopVxB+XtrLYnSGm5PI3jzYh75cNaU+bTwMdQdmrU0zYohE5NL7LL7z
ysSE6nW3Nv7QHql4bIgWUIs3+e9DLFy35I10jQv5NUcElkVX1wg8BCi/yLVcDQu5
bGKEgNp4mEIM4CGve9TfFMn+IQmdfTfKgbPMdJd8YcU9JAXRpLPu/b5ZQkDa4hEt
e55m70gkBbOnq95xfuYD8lkQODUDFKA/7+8ZAeg5jMDqmy+SxKbEfZTsB/U6IPKg
Fl3k0iWtbFChde3ylDf5lsdl6oPMg9pzKmcbwCqWEnKZhaocU+1f6h/LCKLpknxU
4OfRxZ/O1DebuNpEcFtqpogAMe3rNFM/vcNvff4hwit9kpc1xllD9FfvSWMfbrrN
w+ObFt2ajVXNlS78ivZgwtSqAHK4OdAkEsTbS3OjnEO/e3yFa2yfwcwnx3HAHBC1
+/O+VYvcX/UyohA6ObC5EbGP07/rfTb1OqOia7nzZyFhxxEN9Kpj3p3fvmznm0+B
6G8xKmlMKdNldCcGdAylzLQgiZj5/nNcgIdY6hPf7ygqu7Lj7nFzbAjukFeY31d5
jEEa0OsyE2DSvo+DzvWgOJDJEus7JvQe22pfVgm+R/ivWjx9ZKCzkz8C+asOMlKl
aFJ8Q8bPFj9Y8NIqRN1OTZR9+8LssIvNAewzUBiSkJcJSGV0hLQ9m9AlySint15j
7R2SCdHGWLx882Z9gp2jA7N+Gx/Ppv0jm6Ljiq1AQExFyZrtO6poQHvTKWjuVMi9
57KipApJAVVRXOh5NCVtEXhU1SVaMJNXd52AwM/z5Y/gDxETsfKCJ8/PuSJYx4A4
9MsnO3Wu84BJM/VevJqpN9S1Ksb/EcxAaOLtr72xTIA+l8yeIsPZY9TkqiqFWpcV
t4nGoExiA+8eIh3RxoVWMhYVPhcZ2LCZgdTxqnr04CriirXx0JUMTJnf7BtTkk7j
31QpT8suH/0V8b0QeiT3Ek/V/T++snbQM3cS5CW3vcP1mRgVOfTCjMIuUGZFj7fF
OA4kxVgBalVIfNDpesqto/EeiRKmofK+sGxsX7Iq8tdeNmQtYDBVt/WoSBv4JhHF
6E4PDGABhAD55SzbejWbX96nB/KOyRfFFbomFD0/wTgVckTgdmEs8y+uzmt4IPjd
7uqRjZthrB5x9SVzSK3IbyyWNyVX60RCSL+1SWBOr3ZPSJtPXE242ZQL3NUZ539C
fLsm+xWhZ1C9Nc60nSaAr1hFQbr4aUaQpstUVJ5D5ivlg9sg4LSOtI4ISQ62yGjQ
+fzqwuur9vzIv98Yr7V6GEVm8u3oUISqngeoqGNvJpryKFft7kCPshnZFqr3YwoB
nysKnDpWvXS34us/Nf0BkbYGuc9AH/AfoDAHV39XbgGVWQ85VxSTURW939hHu9hw
5ba3IwVM0h9fO9msicqYB4zyohBT9OdBKhiPwwiVysTTrLh/RLCLzR8SerPJe6pk
Eqc26SY3IGmqmrepxwESC5WxrP/k04qiD0rZKV8kcjoAPtfXSIQwEBBCZ4C7jRqv
CHaCGh4O6Ylr/l6NpvO30j1Cep4wQW7ErcU6U0eCCYOegHONlNcq+IDMHMg5wAf5
NCVlBwARlVCc5YxOge/AUJWe/XfEqMXR8uA/MOPCnit1xofxv6RN5kZsyWKrF2g2
TVFwQW+9v+REyDSfQnH3dIDzyLqWBq3JDa4ujUbmx+gBEVF+1fO+eQYJF4AY7GmO
+c7y2XQ2zWv4KYYDK3/54b65kHAO/fTeVigV6UIAa+gJvYgNdF2Zr2OcE6aPqmo0
6Ndm82oA7ga6w7qVsLwEo+yh8DImUl3VU+Hj/Ue3RBmjG23s7+Qnk6tFbBZna4My
NtaZ0wNDx0FW3gkfgFyAgu0gfgtpCBjSFwdKfwsRA6r0RuSf9rZicB/C4MvKWxhL
vJ2qyR7l4PshCt4ZHii0N+V2aLC6E4dd7Wgpn0+ce6CUTqGDSJpcfK0m7Mu8dma+
s/kipVo8jZ6JDnlDCseNRaoeNqIgncs+BVAcUZyKjwimK8QBq8Cgj8T/tedIZoLa
5+l7n7GsNk25knCJE+3R9fZyOq65Ay0dEofPwXrDvZTT2skzbWuIdLtnnzCIMsX5
GXNFxlyy9GmEsApaEIxzms01UmbS4mlo2krohTW9+DGQq9RnNYoUy/oS1pUn2Ro4
81/Fou2PdnGM2zM+8627Qg1rv9xcE/5a1Xf/J3xNz1JHqtA6dRIjnXQNZ10EbjWC
sgZBewF8sSIXyH/jXbJGTIyHILcpot9PyXPVbz7IoT/J1mOHElmOCYgnqrVpWT97
dAcOdupqmC4GDXpbBRRSo72L88qPvwsTnPEzhvNGReSR8BTsik74kcAYGrw0lLRk
fd+Ki9KLEHg4okbZBDc/CfC0sqfCyr6cArzEuXppgycAaRTWEbDLzluqGR33qBlz
xTWbHeQ5CfMKEyjp8wVWBx4TIUjJ34k9FKVs75r9SakDqz3KfE9xsVDf7ppFmsER
WEgzVPG6Qthm66ha+B7726/Xe1MH2/wVc1CXKlRIK8tG0oX3L7jZObI1EuHmTTuk
Jc3qTCkrOvzwnPNQw/b/d756qVdk04ihy/gT0KUG8eI3c2W69uf/Y9NSRoyt9hmV
aC9/L+eOftDh85dqGzjdJfrJY3xdysSjCcHy76bWGW0fhiNjIiknD8JOWKlFKTK8
7Ddrxd9xIFW0ADTIcQVZOMj/rRaZs7RYyzGgRCb1HSVF7zZHKU9FTBk3KBTRZquk
9EZ1Ghm25z6AxeDAott5KCpw62vAY6tWIc3FkE2J+fFoBty92b67SLZOHoqzt9bT
AAONXhulrgdmXVXd/cbNPaRpAzK7bfzBv+X6UdDYXd2yki4V/uQXh+bIUWaBXWNn
7vPWNser71PGlPASQBvjzGM/3mxkLxhqdwoIJplvGbCQhgWZAtPtWgv5JWDpnY31
Nqb6u4QjgtTxY27mmzKnlgfcUtZe2HBAQSLaDUTWAEQAa0XBTyPXO3+ljoNaEgJG
+G7Kg8AMvscecABpvmkHC4vXQj38QL043mZgBI2xE6bD9R279rps7ee8Yw+YbKYi
hYcAhOVjWaMk+1Y17/M4T/vM3KblCEcmh+SzmHIbbGWhYV9Z7pRLQRYvIlHavk2C
gmsaDX8G8KlT/V+4Eooa/qTTl4JVmAoKwJUaqHzSQp8BpgTINyvdPeoX0PrKL/rF
m281a84ZwESAN318mUhYdh7XA7/Le7S3deas7wJmuqQ0QKi2ZLNXrUNbTSnlHoyy
kM4NhOJ4AmJz4ikx5SnaUC36qffUzWT8iB9IiLjCe1rehr5OZYgL8cK68uLnoVW9
oSC6sHfy30fs07ekcicbKg3nJNYUyPZHXWMJTQrF1Su053dqsYGWPfBTOBWH9/k/
RwAvBzwLo3qaOu4akSPh4T7AfW3EiECyjZhkR5NqsldwswPVNzX7aeLQO2cRmObl
/vtz7jt4q3uUxsNbEW7FDyd6FRWCDINMDSPzABSmxNEyJrQXXXmnCCMVxaRtHb4h
r93xuheTiyaTOMjsqLM/g5NjSpXAETd7yurmbVDsI02qywxQiuZXpFfX+2a0AZiA
fLj12sYVmfz0EdKxeEVTl/EiXZFQa/Nym4/xkRFZCge2kRRZ3KxTV81qCRYL+EmT
OLZYBsgTpV4Ielxyp9XN5ceMW/yAUP1DJEQVzHhaPwJKyybbc8KTe90UGcWSuJpP
S/2lx9xUod0F2Scw9x1UQ13v0SN0nxZnZ4WoIaZ9UE4yxZ0sI3oyEOHzt+Ez5x88
WBKe2H4CamQxNvrdgrrw9Csrz3+MFgtQgS4Hd0h8qfXal5CkH8iU2wxrtFLrlykX
i3ydOBG9cJsHshYXS2zd+M4ToTV7/jebRj9WNQDPHuHD09vy4jhuCeg5yuRM/+xq
k7kBpME5F3bGlhe9dA+UUoM+TNsvCoQ+MHXX72eCawThdENCn7WJkb40nvFXjGVZ
6qxQU6OVM3ktRlvS8MjaOY85l33TJmIHyDKqDzd9zI6KTffQamLKm7q1MbiTTb3m
W6RzohsdmxPPLELKx0RRdeuua8OmcynYdeo1XXGBaBE7VqSvLRSfLQ58D7JUHQQD
KcwqFfsKXUcNIwLbsna+d0n9FR70sqn+qAlFgZY5DRiUyT5IEc8Tef6t8IHZ5PVD
J3PP7w6YDbZqrqDArIqYVI3ax+fxjlaYzkB257frBL9Q9oPYhTu4G3lnxirbvvyO
KbsIOq1/Cqb398JOLKLJWPz16OHeiSIynuaRR/oWJsmfCWIc4qIGsL5rryv98GZF
S48fYFh1UtkvJvX5qs4e4zZTNPiYn/dNuM44+NTLcTRf3EogTV7c1RCE6UkfzYkl
WRDg2qUZzb7qK6k693vvMM6USlA0bm5kwbWweR81GTFntLZipnT8WlY7NN0gTvHO
FHBTKybwrNup2ZWi3zeVpc0TOM9y0xr0Fneb2bJqkRfbDByWJgWC+4iiOf5uYfeE
5nsFb2J9SsVv1TE//54Qkef+DJLjaxK76hDaHrugROIRXEfMkIghJwJnPGpCEhw+
8Tm7tSQlmlBxCq6jR9U0fMv4vzljsBs4goxvo0hf0Z022pXIWmvFDBiT8WdMD41C
jkRpvjxGiEodr/+ZPu5FIyZbN7FG9ovHDldJhULzLAWvXcNObfll5+EO+pcROyS6
lhWl7E9fww2lmWNCkMak5dBeH5YH9iiQvd6v+5Hkiy0SWaRXsesw8OEWar2qiaym
ffujcwloAhW1gDIaFzy49qt7lpCUQIO6V35QegK8R9T/VdWen8YSH2Twv2V/opUX
RzFtpVZu+6PQzF7MWyX+4V5bu6WDXreW022lR2awViqh5w+mgrVaesbBWGXihA9T
s3vmIp5myhqyJ2C0UD3MZDKZrS7xCb6bwe+h2WQuIwUiBGu/u8hYC4Pd5mqtSrLm
Ks4QUjXa94BDix9VWyQ22RBcKRrsBEYw3hzUqDDrr4LOEcz4WWz1ucSQYcjwO1Fd
JuJjT8BshjkN/WVHLGk1xDfKVZNbRvlJrvctxfDN4J6CfdYJXYwIWNsEAGn8W/OR
LQ0gsWADwsoxPBRcsQS9Mhj6W/uBvwf/2xHUAPxxCgXaGuQeKhilJX6dKDuw22to
SffOxu9qqLxFm1ZR3Pe4ZesfD0RD0J0Vw59+qvjhZ1of0jLlqp3HnwNLzxhwnqWN
ijPoIIWzuDiNZj4i//V6Hdh+7ZnVN5iNoamjU74CiPRoeWSeKlwNvEkRpZqEL/2e
Ml7Ao0Y/7KceLasLUNdvl/bFpXey3eWHi7PteGGRwGDJCxpl0y+A/+0Hgy/nvm9O
f24SD3bRSLpcwwX7NGPl8xRLaqvfUEJbeM/8M6gi8IlLENiSJmWIY2FHpysb/unm
rHx6UEl67Z9tY7AlBEqeMYBwQN4ytp2K5ZMBHGDa7/Li5kgmM90odbx7+2nk1ApQ
8vdT28ZuH7OaiGLekO/I9ruoqeukYFOy+EAc8B5vxR90KhrDJa0fn1leCsWDZrfC
JfAcvpv57m5F9CE7yD/PoEp/VX7TmoAC569AWzEHMmsMUccgIm3bRd+Uy3ygC8Wa
O+gwVvVsR7f2Okpvwl5Wpd6zdqgtil3DpHI3TXH1ipeJsZmbEIwfEA5OYd+aExD0
3I0c2k6KqLDFmIk5fCUlnnloy9KguJdOgmcvEoBTY0lGKds2sSEW/zdJWFT+P7uS
gnjBGE/UPNZk6xD5JNvy8YE5DxxYg1gdq5frhOjpXb5Cg3p2mK19WTT3H46sJTp5
peTy5TXB+ubV7Lgd9HoWBjeQoa7Fo/tnalrtpvCc5yZgHU/GSyXf1sLVDzhh7yl9
E+xBLuaFy8iWa2chGjXYyUHAtlRQtvQZwz0oqNwTIDIe661KBUyLB20WWvrpzClY
YkPEG+evL1cL4F/anFp6PQUwAEBvdiWS5sL6YSwaCKxwnHMv9iED9xcCZgCGTmoL
c87AxDoYI3JZW1Qw84muPAorBPc4MCTLatFT/5UC2pMIi8xK/KRaJZj6dB5L0HtI
R0HSC7XlxBMrK6P2raFZs4aL3AVbH9rjWJ9L75AEsJwd0gwbZCcCBBKIYQYmHeNd
MWGrOd9tvgBmiFwbrWLfEh7dgop1uXr1+ofKhPbQGnANVJnFHp4OcgVjgAuIUFDP
bweCfXi0zqHg0hjbjqZR6xLtMZXcgpOX/A3TNZhitEs7YWmuj8pFneGqrNHiOltj
+rVO6qmnfqTkq9ZyYnA+pRE0k7g4gyOzlmDOfQL0bB0QKCFPuDIVdGRE9upabz8m
xPo/8QRIOVikt55AjdcPKl6TRGX2h02gT2CyTVKk5jxutzBozVvobR6reKravhBd
1A94dzOMsCyz+ZVTU+LOBixFXcPMtXcF5wAUO6c7MQijHylEIpx8Y2FNBIQ8pfv6
dXvJdXILs2mAgA6iHeaAUySTyaLUWkja1L6f16Aban2ACD+2jhuDxL9uQichxN1a
yldkixOttwy7fpdJRar6VQCd1/ZJl08sHMkIPAGkh3enJ9j6QE18/J+vN0JEpBpK
UZZrBCtHk/RrVGhkf+enzeH3y+atcALDmNmBLRMJLlHTx/3DMnMLEHCvtqoRbZWB
IoeqBfqh7NMT3jb77IqaBMX5hV9TrAD5eNvVsu9oR7rNPfUTh0Eue+iJ+PR2LBVI
+QDeUBcD/xpIgGxf7EZqICRyC/B+xdd5yARhx3kOAQht24EvFDEX3GS7M2Hc3PJb
rbEW16RDgA7p7iJ8X/0RcKd1ed66cCJ8oMkRhRxzMcPF7mIdeOwkbBca88aHqKmM
IW8rtQtrYbOBy4EhIr9QTnbDPJjOuPytYn6IbdHb6hp6rthlDtYt2VbhTbMrnQaa
m0YZRwEnWXEOXjBgQh5zB/OqjdJ/+nir2s6L8/d85mNp3GJr5R5GTy8o8a/6cIVF
Jm8YnISY1MfVwg2z+gvsaIYnO2edCCemhIyW6NilrXGkCmNqJ7bS8fxlosxpjsBS
6IF/nUHnP/bLfqypH1kYl8OzCzME4vDgekMEiw46QfEaw+GT1JAhf8cehC+N24wW
6r4I7hkStZmEgthPUNDh0J0eC/9qEjsnW7awl7COw8TbaAX4x7whcFnoTA8DjhJo
B8itKBfwNHfW+J2Rh5JURaxKIi5CAXPV5hcw5VmXjGFFNGlTtYIh0O2MrSkpw/LT
zngDAXphJ9r4n+AJEQ9YJvrh7/mpcn4UoVxSCuw3OGGAd1djtLM7dpdzVoM1EbAw
JSFEWXrSwUjRMxmLKGL+RJi51JZgV1MVrdGVAiK8bKJt8N8ROqh8N2daNtsbwRaV
d48U94fz6tOscvQJHH5Xwhvyk1+Lf5ysHmKSsWZMndPQ0SJlyRwqtw0/4i7f/YCD
wc+C/cES8Ts9Dltpe0jU2rg7G0i+nzPOslefTqQ2/hpzjqDjnFQkBvosgrxQuIlf
1c4S4XmL8OR+xn+nQWgpq2AHuvqrb6q6/oOwDRjZ5v2c5cR8Q/g3aJFhI+UX+qEI
yPSVoyNfs8ejXJJuXOmgba4IYFGAPpELQCB2rzcqMKKa9T0VVG9fflOKmDf1qJbJ
qfXZTXOZBBP22FnQ8rzryFEZ/LMTT5mDlKMRrq+F60pc4E4YvmnWIZCTBoqrPOww
VdTcu6wz9xU8djUVERMBapoD1rmaaVUZei2MSUcKj4h7FIK2KLt7zMDeNPncAawi
4g9MWLXlpRu2NF3UJTqw6DNpX9h/kB1/4avlb4CmKhXqT4GIwi7ttShsCGRinJ9u
8Tc8MapeIQ7zYss42Fy2cJz4jhsQALLpnrOjv7le0BkSeISxbHV1ybCcxS2Dzi86
CPGzfbDQObfGiPuCYnr6GjoPn/p96H3xeqF+kVFARjVjksF+WeFUhI9AyFNdJfY+
iK6Oyg2MLCgYLP6nSr3obADegFo9R/1sAaVNR+NCKTRR1jVrf+KA6N/S8shiW0UQ
EumCfXqqQHidJSN2AIU2y38lXrfQWrmxK3x/0onr+rK5b/1NQSuzENOGKxxHz12+
yxWsCZfR59I5uUUQ3vWKLM7h17ClbyLXHxNP4koABSIJz9OBT/Qzh4fW/N2N8lQr
iSoOKDhdRAEUvrzEJk7BSbJKRzZHvfkHJoF7J8J9SckkY5fjJxqFUIErMEMrSMiT
dVQM/4vTF+Lc7TBtWrAXSKVkxmu6f3aFxHewEGjmECwoo7Yru52IyPtLb8AAuBlL
PSDXMQ5RtxcEuDERRH91ItAdI0aJoEjw/sOX+OweCWjFvbl/T41f4XB2jt1FsU+3
OqWeYLj/mbXpBwnQyJ6e46Wawr7VCnGJqUoKZJ93JuriBdXhXSwkbcZTdobS/oK+
J2OLbtQZfYF4S06f7njRFnGxmHkJlOMh95JARGTbMKYYdA2P/qmZXCciBQJ3x3oP
TVofMWusBj55VGXo4bWtW7kbs8cWJfeb7h+cU18OW37X+/GuG7+Rnmra+A+Q0WfR
ffISPRQmz2pT4vf8oAmiaIMjXpAQi8K3ODbNpXGnJ96vyQnfm0Ift8DefizgsLMM
StwkEeRJOqHiBZIYlDw4rSm/lGfQ8wxDCLikwFiweaSgTDSJ2GmRX3nzPc+B0Gia
LWh6WIfAx0+rBJfUHv+Zol7HOdZ1iKAk+6yPgOczrDCNdskD6jv1tx4Y0UQoZyEk
BZOoqcMg+hUv40ZOtDFBfOZRHYklu1vAGQjc+TPnzW54aAHqCEWw136LBfzds5O4
jegJPNNrrQdIQ+bowRXVFfOoFVw9l1qNn1Or97HmDzb6BupuTQAhU99inTAB19KQ
CDAxppir4/asv9MdTAtr0EjaJgO3PMdgSPZfkXFoJPDADCo8AEEy/xbC0znK/ykl
V2LxvZ2mGA9/6+MCCk576IDDrqWYsapPxYkIrwTKAkx9DiokS1unMyYoMHapVv5h
eJcr0uBkrRbZ84c/0WUX12qIL/j+XPXXRv8m3DjdNhPsBC6i8T/rqBJstJmlXz2c
+rDYGVTsi+u+wtFbTTWDaAZoZ7XdDjin9M2nfqXEhtUWaADRj7Z7rCc8eMiluSrV
VXC+EWUuEhZWL+N+9g7VNnD4RchcklKBW0ozn15PFIQeEC4aD/j2L9MIlLQm8TxR
4RqjXZV05OXxQ5A7d14mq/r4fmANJW3vpVHDaV2p0laH8eGqL3ZFiWfzF3C8So/G
45gWsYpVCSdyfasR4rrKZLCW51YUUUbdpImdj4qHxWf2rSQFcFoSTby5+cHjDRR8
W+YDQ5nC2ssgNQ9Bd1ayZQQxi4zw51HlRZuc2wK9SDRsbNcEuqybJJ87wyi9FGSk
9FrhB0YZ5dC4ooHgorhafCO9XC8WQw/6llCzX7+QOh6Av9SEjyL6wxkHXJRs4PCs
1HmhKWJSmpq30z/nJ87H/rA6NleIhzdZi4b5agREZs4gcgbSvp64ucqPY5mgO3IF
J96iGheX8yUFhUJACjaLwWUlu8hX003GAq0GdfuzWj1pri8PcPL7I+Xq5LXoc2sA
xFWkOULStVKmIp1YwOzo0Jyw9Fwig1muAwx0oP83x3KoFvnMobdqNsz1ziJDM2hH
q5Nj/GuZjUU9BQNv4ioEmTWgum+6ySaB/fUcBlOdUki6I5cz4ezCycxrmPaYTa9G
O5MZxhUe8uvL4MSP9aNc6KBkH49orW2hpTSdiSGDizOJa3aKp8UDfNb6Br7dRlJF
diILT78bvDcxtprpoAp0JAAGdIkdBLhZUPQ+RZDbDheWOokaHgQt1KAy9weDt6h7
aZSjBNbXFhwTNm7hNNCHHBj5VnPQb7zwCaqFd/yFP0kGYy/8EwZSEqjo/CQYIddd
2/IJdIa87VCC93SPY4QmEYaQ69c7eqmHpHp/H2ytxO6+fqgT+6kMS95DF3QJHNLl
7Q5V3diqvNpqD6UGhJ33HNt2j+nNKXOFmoIsX899Ec4EuIAI64gBIHwX/43Xf7rg
XO8pMheGTJjXeBw/bS4iT5Kbpo1rE5tiZIEopG5TFq9UVEv5MdkHGvnLNZAPDF4g
A/wnl+lvH3FV8/rgZj7SE++2nUNFoh+1JauyGZD2NFZUO9rEeM6xONhvlFkym3Oo
GhZe/ouon5+SgYMGMYVnfsaxaDZ8Gus1pa15v/xKhva//ukosaN/6MnHvFTU2a/L
MnmukDl1HI8kH/UI3IkAShTbbEB7sVz/RQsDjs7+o66d0NyY26xTwvCeACJDNfcq
tSqRlYX1EFJ36wsHPXPaTftpJ9AJgaJzh6NBZONJUixPiuHefBPIhfiGAD+aEPV9
gKAva9DR84SQB2GadLeNnOIlbUKQZZQGp+YuJBbbTkwylKIJv9Ha+gWhh4+0cIIa
cboNomEb3K67MuJ6Zo9+a91CKywfVNBkK16+SkeBBZc7iCEUqI43MgNLKFdxyKu/
gh4bya2UaWyAh6ncVVz4p3oODj8NLWqB5D9yprc40UoL+QlreQc/sbDlnc0HvIbD
OZDHWV/oI8duZqThAYPF9OE18UPsRMUHdoejoNrHnpJIvLMAJFHaujSQKI5CljFS
YNf3Az7CURExKQ+asbI8aqLBvku+2sgM6ACnGTYEwPpNTghu86+Zc+S3hvilI/ua
rQDhNCC1GHqZGt1ABM2iw6jQzPXltnv/jyDlrXUPJfE1OloKl6upq5pFXYZWEnyM
HRbXyUuwkAkdmj5Gx7FKip6lPJaal+8DZd6BwM5N8EVKTs1r/e+AdLBmrLJM+KAI
XrsCOqp4vd9/zwO5N/SI8jze5ofmXrQ/sH4JL67d+OC4CHX5C1WppdQJMLXcCWcw
7rDllgvBYluMYtfGe2H5d2urN1UDJK7pMUI7J4L8qsK3qtyoEqzp+eXHvgLXi5+V
wGqrWXQIRNhz1FvWNpoG7eKTqv88GMtcpGBWe4XX8vdPIiPI6mzwPyS19AkFRTYt
+e5CSfdiBTMsQOLbJQhD9T6ByXGRU7u8qt2YJbQkqzMhEgbdRkwBGLEFEKn0fD6X
k/dF1OV1F+hjJiDTn8Z8i7WIrNYnB2gyfRJftOsxY4CWgoCQprzK1JgZTuZrE0eD
TW0k9/bmSYIhUBE4UledYRYw3qfrvp9d5i08b6uFTRyjq6XLUIo6uEJLMzjVrlmR
MagFC3wEsLhoMHemhD2ugcLer4aLuKHuNUxbRNrRAMtiLT4Lpj6NlL303gnbikrN
NAkf7VeoYFdVBLK2bmB/vMDjP0XrOs7AvBN0KPSWkSjZU8So2dinL95wibunI+Rt
LUqPeJHHqYxjuu6w9FPSvJvFEhWWKrOnxhl9eGPULLVNv4IykV5IdAhd7m10DRE4
0QY+kKvX64S7bqyPue8GnXt7KM+v+oTxJT89msfsKXsJssaIuwQgeNC+c4FjyfGm
PZZuqM5zUnBPAj1CK64wAd5xr6QX0RiIGqqOouMsQA0gl3mG5lGDF85UuLo4zKrl
B4xkn2rgKtoO2lBKJtNPWdav9EoJdySTs0wj2PCcIr0bAn1J7x1IAEVbH5Uqxrdj
2bx+Gm7lkz4d3z+yc5dr3uf3NxEk+98iaRKZfy3oUPStannQU4giBpp8DYa1i/f8
cZTfgNvHq3Fcs2TIMVDh/V3Sfs0cmTQh6sWKxXqzgUDDQd6kuq61M5UjVWlyU2aX
V6OGwGNfSjWaecD+sByevH+RzPRrkHivaGffdoPFAT8Fp2NKWK8zHHHj5zZe5GWu
OqVoxF4IahzkgwCM1GB1bLQ3aBUcEXa8FYpwOjb+OzrvHIzHPHz9Cx9UkrVkoYki
C3GEEGkJKmntQj7IR0I2qQz/nev9e2NJtOrHL/F7KqEDhl4MHppiV/OhgULmOIVK
6ONVL7ZPgLoP/trUt04Jtqy2clERvCVZChKgxfc2A7P3d9ZokjPkUoHbmBWzuI17
S1Z4r7tYWrHib5zh1BXrMFLyRRbsduzmM9u0b31j6vzGQ+JOsz5lG54gi9GcyxdI
SqyN3JJKeG9M7RXGxERo3A2XEa8OeDRJvojYDmxdzYZxY5ChikdW4xuVLjsqiekw
NNZ7Wd6+cq9mNqhCDofu51U9aCL+lWBBFAazRtWesyQpgD0KJB5Gf77eV0giJ3Cs
Wp2zup428X8sTOTtX4OXBOTbHswJbzsKeQ3Bh2VOH4R+mNCFK52d9XBKmwl1f1Ob
QMmbi3uN17f2bz1X/C1CyY6XsOgIjfmCQrV0QREC4vbhz0uGwbRVZSHsSESRp9fQ
C0Dl/cX4lmUGIPYVbR/EPx3UdtCcD97WN97b3hsrvZk35dirg9wt8ndf1ngiOEUi
urqYWgyl2d5X4zgl7rJnTKxmBvBrQRhljy+1a7ODM6yIMQ4Q1lAwzqgD22YJMqjh
pNPqwUqRGRWsHHs4ZVJKPK+optt7kS4ucZVoT1CQUoDCYC6buzZJXDucFbAhwqrP
wnGH/MVMGBbhNP7447RtMHmfVaShu1QkoaI33i8nW4gcHx6F148XVne+XwmFKj1p
nXf5NUgpyu628pjFCH1/kTkFjIPoIkYyUG7aUWBL3MIW32a5im9oGsANWYsWkaoW
mPGwKNaBTy3PEClpwGzjODoWcSWopny3DB2rIblK6SQZtIiL9XrQZErsKKIbWnhk
qhodVzPK3iNMDeWcu2xqFD3aQNOUlaKW0VvA4T4EjRulKpK02TtsnhgMEbxzMPbr
0E/ZmfygLfG4lFpCEzC+5FvmfNncIFonbuMQAsem9LL6oobRMRwSC0xv6GY3hhNp
ibeqE0If0wtKiTA3mi9O5orhFQNRoWqGJk0V/VT6KnvUFc96uh14Q8XgmY9PXf1X
+qOwJq1z//BeYB+MufsIX073pz69psSuIWUXuCHq7bhmoGPLxyX4bBMJLrLTFS63
YxSWcvMUkNK6vz1pfAnf85g530xFrJ4zcuzPIdasZeh36+Lr/Q593J6dg4Je3i6G
GaXrRYPZrvU/tAYKct24pgUXMcCPA/syB2eQ0vz/FrzrA1yCCopT1oRQrYI2wQXB
G+qNcVkEMHcyrjyCCr9G2PQpsFnkFwbgMnVJwNb3pOqVfsRQ7Kath/D1y2b4w+Mj
v07rQ9BOJv2sykcpq9rf6usAOb36mac4WGyn5FnKHjtnXCoh4rOcm+oAKmHu4jmP
+nGUF647FSvos/KKoIETmq5uwDn6xZa+rUxvBInx6TZc4TCTOtI9k/sYdkdzFZfK
WqX/3UD2wLuIzZ7siULGdJA+EMkBqJphqYLk9dBl3my9qleJAkkFTwlYngW5YzDH
mrjsOZEAWnMN0ggab7HgiwZn05t6g5+4Xv4QtOpw/ZIFEGxVp8ZqtimYWV4QOcyj
btVJK1vqAAyetS8Jf7aPw61UGWccJpRS9igjX3/IJkeWzoMQt3B4F1zS7qkqlxdM
nSEIdk3lhXHTAov9mRUeF3FqtnuzzTs2iZL3VWsQ9gGmVyTScDfhzmKSqdpYtToG
U81QPt7HOm3ubChcZRPNA5Lm4HQ1cX01eWwzN1FYL6h17s9RP8x3SefZ4si7JMzz
qAiERYdptaTe1VvYHpSUnXW0RlRkuKNDA6lSzs9WTtls9P/FElbhcUYURuQ63nXi
anLzYNiheWIT6LDbknuzRzCahtJGA1ehVhHE6zKp1vSVtzaCS/24u3R3Mp6oeJ/r
bU7GIe84H52IiOKuAyTlWbNlosUTWtnXFu9+eAMZlDNVnNjj9B0F0juANlz9tQs5
egUpfcGUD9qSJ/ovyNTFZ+FtsLvCUjkCk2Bfd9G/XLlkiMsl34KEpKVMFsBdRJwW
w7kUtYBIi+UJfDPpk5OR3x8zaJiGmcN7s/Z7Sv3Gv7tDT+ITPXAbrVQYKbZAGBpn
PQ4ean6nua/HUo+KbEIJa8l8kpVrTZvvfoFGeYD3RI2EMSk3t8LhhXsjwsCG8wyV
zkdUMlw9sCpaFPscJyHYUB8noC7566+eg6vNoTjPnarMvmeShmHZfZgND/1VrxU4
XTveWuK0mG/s+xvqhYgSfMp0XicTLvr7tGHp8q2vHeH2pJTs9aN+nZRau08GNBza
E+AfOa3ioJhN+AfQq3kCrjSrzWmpPALCGiSfgRF1p+hSYp/z3m1+C9tTtKI+Xccy
iWfhoT5/PXizyYA6C9fE9BZ8qhDeRHVE9in7WLGlQt4RnK0U+uFRLOnffxbGnWkf
8c64ORSLE/Q9jKdRSS/U6IX1MJlqGg8ldyhDNRuA6/Om36AxMQD+F1uAH52ghxmg
R2YJPfJ5mLNrHVc4ivTzR3EZ5RcQZB1Q7Z24+4uFA3Us9fsRkMjCh9gve6iIHFTw
GdSDqMnV32/U5DfnwXDkfW6vNsMrAwB/zCaZRk4CStrTmMwsc9p9384k4jO5marm
7Y388Y6nEG7quWadVLNYPMxxL/gFr0XgE3xY4Y9/b9Gm2ecvKmOhIPh66uy0Kj5d
gLDMh9Ure1lNY15vLGvy4Q+sEWxAP04GVeZf6TXmAlKJibq3CLptfJzl87EdoBXR
3jYqZOYCkJx8RLIVSUY6pXtN05ssrpVbzIepIp790Gq7sF0loswfyFgFX8BVzIQf
z5vaTK65GTt0L9oQOMoqB8b8NELCLXgfBOB90XG/EsgqjaEHnUM7NgC251cNLjH3
8iHRA8ScIxCmnKYcl0X1sQaNbx8uLOFgDnL+/4DBc2qsM5IHnRb9BThMwI++WUaN
noysmFwPQp86bgddSuTdFS+PbWzVMPeDOHdMZ8/Twj05KPrXAM/13tcXJQrsx005
Tda1+45H8wgldOK9mgduYmLMKO2cxVZH49/jTSz0QZ3Af9sQ33dcx8fTdHwge+u6
KASotxBRsqlXtq5U3krXMnvcyrhYcPvP7I54ZSky5zfVDbbcSUkSG5tU2ABnCvOJ
mGMdthjvnMl3K7rOvBXdPqDkXsggNYw0NPWPzbtBXQEvdZ2OWgNGOaubOdRvU+T+
DESmFuhBa8dQwlPDw77OSZ5YWFTs9JBqRBER2Cfkdx/j7IyeS6zOBiksq4HKBIR/
EYFxTMibP3H+jhGBBRqtpsL5kShog/yNipfjR9hsqkRAi1GKXgEY41aT/0eCq/tC
L/+EgUYv9xWi4gEXk6mRvTt2kVMiObLlZPuVo+3PqznOqcN9ts1Pkb/GBlbB+3aY
nXQ0V1rW54709W9BlkU4CBWIZwMD7TWE+4aNQ7bvjdxlIOHntGmt3lJqgEb8kv2U
JIR0xr+oRr9NXFTjMTc4+NWD+KL+/eQQR1f2EkKwcL1I6EEsfPXy5D/d+1d+2kkT
7L14r67sNNDuig6RFlXdwqpu14fiflRcYT8ABNKv/ttkMeoI8imKbI8jOVtIdGFU
GctpV2YB2IBUxxfRujlcMbufnZX8o+bTTw4xFOE0u7cf1JfdzMidF0pHAWSuMphc
27OovgAXNpY0Wan99UPl6upR+X84gDF9jX1WyNjYlMEJKXEkFZp2UypT7kGO165N
yQ2AnGOs4ig0ZYZdNHljMYYz5Qrd7or6ooVXA0ddtmjNJn0yBLseUyi2S+5Vr2DP
BmsglgmuPM+U1BuY3Eag/DTSEf4JMfViVoVfKp1craNoGYLr2A+s3MG9mZq9WNnI
5KjdLpAMLb94k7jYD5BKtxyes2pfI8EG5z0x56iImbErQaadxX1ohfbT1Z+uWeiP
OKN2Mxt0spt4MzQfmdQcGsDOqo2ycPKioLqWRbig+0foT+7NZSKpoRAGLV+8Tdx+
ZmNjuqbB7YYdNXEAE+a5EXyQLvfyuB77MKJ6LOP4lhojEMiJChdGDNeJKooCdqvg
iFoKk/utMFivvSoGi4Z80WCMxMlPbIyRc4EuhJ2Q4o6D9RGu+SMsCzwFop1z5Tmh
8z+Mfr8kgo02n7zNLX5zeAS26RQWtAb1+SzwFHRaU9W9E2Xjz0JzqXCqvuG6abpy
7LUPzcu3RclVxsUng1BHHwTZcxpPyIUHdCPjcnp9yl7Uof0mRRFBWu4cgH01I3Gt
KRnK0wesvX5QoXqYwfT2TJlLPgi9zTaBYL7WJQ3pXW/vazdDucZtfDQJDaEFbW9J
rQhJrIux0OEEi6A1AZvXAnpj0tR1jr3f6Sl3Z5qbmwQcdFNAp3u1Y0ieVU7KQQ4Y
l2NtBXMDMXGL/HetidlHgj8jZHEMnmwXF0EKN9zvnvDRk11hVnZK8f/gTQ5SEIUA
mtsXk9ZCHFS9g9Fsq74oitCBwp7nqib5PC65lV8vZKUMTeZ8ZURweTroYpscf9FB
5CznZPAylB80XxmcUpg7tPYbqAmfIO2Fb3b6O/IXxwVDX+choF+kaxTMH0FEtGTa
WmPUFc5qp2/r8D6dotbk6r68Qgtc4WFwAFrPH1BhE7/7pTMZexBET00Sdv5fFV9s
Eb4xF6laC64sZSGGgUDirjhy68nNUgELdJosaVY2CMkFB3YywAgtn3DZkgJeG5+X
wxhexN0xb3DLyJsmIxX242AEn62N1veWx/PJGyldFVWdCSu8buhglTA7VaxNOQaS
Y59kEt1e0V/xHO90inponuQIEJU0dipSz58aUXDe+AbyaSsnBJJufjlZKhbBCeR2
mIn+3n0atNdtPb2ef0fmLg9oaIJYtFqdQS14H++ZJYBXg9aMjeX9DLcSUZ6C+u9Q
sZmARXOIWuNd6SvOUNHr/VfNWHbnAIbhdZCkXeXCvFARuLexePLkAqlo/SHc71pW
gNjZmeZYsfmUuDF84ZpUGKDh3HDr5Yw6xnOOpCSFq4N1TVYP2RxcqbWc5Q2vzIb5
r3BJu0tK4Cwyd3NlDuQ5xXnXahfDSBf5TM3D127P6eKXFKlemBLfCsO+3hbZVj9u
5NykMZyhbDib/uf7LwgGucMryaxL0jn3u1wypIR3PlsnRww6ShqKtQ8RTn/XOUwG
nK+2gjjtghV7tcpRmZdTvWJnhKAKTCEWKrNzi3qaO+7pk8Yj4Wz7TgJZZr7DjCq+
kinRt6RFmfLysdxrK/vk9hyUjxXZQ/rZkExim2YcYSZe+nQOAFY1dQZ6cUh9CVpJ
R0+d4nUIuhq2/xgMyLtr8tm5TyoJ3/zHtbQmcATndvH8cNkLY7XxR3PizSQVihoK
0oI2Zi3iFU+9Juxb7ox24gGYUnAOorpnVDksIi6X7rBJkszk4RpcokNZyR5R4aDK
RS3PsX5rU1dCVHIzhr7VYLH3tQue+sV0YmdkleX/XBjHvOBfeW+ko5SeRs+vk3dG
OHp5YLfgQk+altYaNBDHN0DsIo2MR7ZirOJxrW8dlwgXbOEQmQKdSOy3/85xklTo
6nJWbZUCAXHAr+LytQdDyeQoV+igvzkcZ8CRJ3P8NsACHpCrO6JlvFSZyWbCXE5+
S36aIoZLbCsV3KnHYmdvvVz09Q4JWnM0SlxsDdYeu1fnuc0T48EURCU4oUpak58T
/PXsu1xKiYF0KYHgicmDq7W/Fd9FRXY6b2LeBZ/sJvG4APFJRnt99RswqGblgvEt
FKreFIe++spBkCDjo9nPYoMMwoTxox8edMo/XPx2TI4BSPueCUYKxAaCtacHmJ3r
Yehlf9eWGA4mZ0dfO17iTEFM1GAejFFZNJj0hxnfMElw3YUq48KAzSdv3az0YSCP
sW3mbQtPEy0coHdssbI1VUdqwGfjFITQdUzP2+7EVu1+AdE5ZACLcWEVRsKFvoYP
lQkTVNDup3HH8qn31a4kT7j+B9a34J0PKXXVN4hz7zYBq4aL9rDEiUpnQhPsEJlK
4Pml1hnRk9T5E5V0hhoBaKfGbrBmib13Pyf1AUlKKOqTdJNpWsmc5OvC6UYdwZoz
YtFu2W5D+t5KWwmGFiHdoLWqaEH2Eczzu/sH4jZE/CVLBLAVoX6A5KZhhoejUkEM
97l/krC5APPurYtV3Y9/9W6i2Nc1aIZIwDHDecg56PYnQal02N+z5GEAJZivzSXH
1/1z7C/+GoZ791fGXAQHF01rE2hcDiApyyLGflWLTwo5hLR51n9z2BQLP/QdEI6k
N9zi6jmH1CBTUqUmceTTweL7SkTIo+7HVc9bBMtbQaQpN0dNAmksMTk2ORziOGe6
V7uw5en1BCf6UWPGdXLIsg3XoXoRmy2bNwLxhtAnSizDgQ2tA9sua/4w71JRbUL8
lvpqxrr+v3cQZsiWHPitTanV26tLEHikGD+yTBZrc1oEARLA5dfQVlf7/7j79oAF
uaiAui0KseZS4raxRJGfWMRRpyXVfxXRZoWH5q0YOD3Up81qQjP6wNV7CNC2Ddig
PkMeMysbIfaoTUSSMiXWstnuyJoB2SlnTSWF/dhbCIp0HaPpVzAaoQNkItgfv4zd
iUduzkApcanxWnoA+ujm/lJ17h3RzS02gX6F+8ek5f0f+agukjYfF5W1V0KDkqT7
qZj8aDhmP1iiiP9GdwzB3RaMT7iWaYPR5yEEgtix0qEhFBt87KkHndPjcfTE1gq3
LkB6w4CCEGbuB6YdExLDObSV0Ehgjn/MjZVrdX7T0pHdoRpEsqwAQZBQsfPDdARz
yrHjdAVEdv9dQKuHdTVGrQzpQ8Y1vgorqnReKR51Hqut10rqT/ym3oRbZx+5GBEn
rqKP5ubn/xwGsThTocMWUXR9nISzrqUpUMGYGCqU8xLkQd17QFJ5VC+/nkzJUhZC
dPI6aEUkhm+iz06A3CH5mO89FPlkJGYBUHjUDPvZ5nz/aOs79j025P5AxA8c2OuF
GoixBnnv91Q0EiHRy16YWJYFJVs990XBQBJr4rH5X5S/j/LhOkcFdbrveKq75I4U
MHBS5baRcZ99A2vKJDWAZs7YOU30727XCOb2hWwBKcQRgqeRN9vApn1A3Ow0nR0j
gv35mu2Clj9UC2g0f9LbPZ3Ut53AgsLIFQapU/ayXEMP86fu/kyII4f54aYMcD+K
n/L0Z75IogToNJbFjvNf17ezNbRUnzst3jhN0yxZz0Dx7lOKd1c8vcw7wPthVYNB
/xnM1xEuXCSLXHjQriFvXHP1IntbP2F4mh202rlmsPkOTFp0zVYZrgDLAKia7xtx
+Oq4bunPHHqbyXHOk40kzcP/1Vq4YTQwzwv2upHsPngpSOIpZ6USk6yLHzZvt9tT
ZKubUSvg9zLOliDUOihBu2HnSgUPj28s5Ucoh1jPQftOYqrJuvFwOm8lOcrpwb8f
cOxK99S7J8mFDlonpDCghuojy/JPA3lxaH7OJKZQJviyOLiYTRN68n4nL4iB+cx2
QWbX7WQZ1+kcRtkRGwKnvtlIThH9P+WJaVgJk61LOIpJ7D49xTMwyr9/Ah4eGg4p
mVX4fvC97gczYCvWP4zrfxIpaIR4cqYMirpmc8ZWoKyjEUkdUwTEQMd6zEJyOAh9
hIO0/p/R9DsiZjeE4xIUdWzTc+eUCK/Q+MGX/879X583o8kc2rv1tOTbTjBFwPul
7deE/LGO7xbSIeMm7RSJ8ZXLWxVSBXOE7G09463qzDLhK/laf4FSnkopkvu1hOZg
9R5TNNY74YcFEEryGAskc5XuksY9oKF4svcgfwTc9+3RkgeEZ1hTIqQqHpIN7QkA
DNhVoXelFq7b9Z6pvz1p9M5GmLgeHY4pmQ8BXZwjYsT6bKoibhZsPQdFo1fnSNu7
Ql5kvCKErFkb3JSAFbHk/aEqQqcqH0VOHv9ExEm4356FszRKUrPTSYqA6p4sTaHt
Ms3c0pGUab7KV1UYTxHrrk8iRr0xMrwlMggw22YAwrZMZy9SvtJut9dnlBu5xoxf
VyyngkyatqKN5cwhWNRWpc0Db54mDcXxF9vk6oBvMTm7X3QYaOASMNMPRxdKnblS
T9SX8qDJ9aJIyuUIjw1alyUjNuRoV3IYrADyXUyLE/O5X+Vbwaa2f0TSQwANO0ZT
KEFjphRstmks3bpGLTh/7g+RzDAMllNaod78jnLHNxxMQU7i5f544WHi69Ye30tX
d9yr/pipufXrBOZeAdYxTKR75yweUbzP90IL4i0eP80j7D+MNfdsPmgq2prtbGTB
hqIpUN9GmVnEn4usyEwTOUmqgy//xpMo8b1zZe4oS5merf4QA9O2/5Gl5fmdD1oq
T5yEMPNOXHzVCUf2zLzgkS/QJX5uo2L76YSsRrRlkO5caWPJByd9u5am2dUEgRuo
3ZycPD4jxX98vSoK4BhFBoanna5gHjVUaAaU6Brir5rBmPK8nwiaxGMHelO4h8yk
45rU9MzEc3wOZRVUCqmqbzcEP7Fnt0ocQ3SPaXMXM+xCSpEs+ThhKsSUCSmpHrSg
pLhc7s8Tt6g63zOrQUo0GgFDFSK2NzzGDrgz+aPNRb2oKlR7z0m+jcGpHIe8w7q/
Dr5MHCJf9BVqNQRImg4REyNWazFKwp5dJpCVnD/nKQesNuZx0OmoBKPq4phouog3
HLhxhFUpZN//sjuMTptP7HXbdztWbTHI8MgAXBnzXn75swr1tCq+/N4jbbleJSAx
DahnPWynCH5t8ef+UjLexQqtjNOsKOHVLZHBr0oB8mwJktsLf4kKCcRXubCe3WHU
Idped948cgAnwX6FjZy5SuE+HyevG99WJsHPcJwZ4ggvIObk9XBCIk6phCC1rGfe
aY8ax4Kh+su5ujvgmjWWmwi6xMOGAx2V1u5KwvEIvzpmw/oKobWrjGFMdh+8DUia
Il+/5XAha6ULvAUrSWCAxswLp6ss7rLAjjIteGpVo7B1RJpmnh+sDTj5P+oRtoOG
uM7UtbdOOslYDQDnXabQFRknXmAMLKiCdRmqo/7FSrmrDUkyyphrxpRswaR+TdWE
UcX3F1ewGl96Zpq3S/T5q/fXtcnSS6Xe1ED3tTjLuIhN2Bf6a3MhCwO8kyMzClfW
2fZl5zfQeU4OCfCt58wNA02c+auJB5d2Ca1QX2EUG2J6nfFDmjwqJxOuG7FHFovA
6YLWY+bp1F469K7Iz+10xLdNpvBOfosWk8r4bcLwpID1KKkQ5F5AEPQPRBihKdkN
Vl1OOGcYhl5smP1BHIvNvZ69zsqddAQV7UApBJi713QjGBrfFvEeYAgAjhvqZGmS
nqq1+xutc+SfQTUOOZtWfv/RjkKAQYXw4UrGFKBJaagXfupEzbo2WO6wpHKCuMLR
JZLaC/OmCreQ3l4RywEKcfiYxTx99eFqv9NhMPju4t4EYj/j8M2l3TiarjmCC5o0
9qOmF+G8UsLEU6Fc3JRsxzg4pyHEAoILcNTDaPfKQyfzepIBJgiXXUahdEztRaOV
hZFS4WkLv6A5FaCmEfplHac8aNmIEqALNYOGkxTA8gA7/wGIwWRKOgpmp0QUuM8V
66tT5k+lxzhRaEXuome38Fegh3StSxNhkv9I+PS2+X8PrgU9vI4nq/CE9omJCi/v
y18Md2Ljpvd5J5ujjT8okmS43RqObJzirfDgJJYapC0ozSpHu0RwrtOg2EB31Jch
HDdPEvIgBqyfibdu7u11Ur4jm2PmMrklzOwu6Um7yHluticTiNYmisxt+rpM8NNn
AJTML4E2XCAw2LTcF0fGocCngWGJz6RgsUKgVLhWSoMK7rAxtjJD7bojZT3LRwpn
J5kdeqnU6E9Io3jU989b8i7DQAai8mgzDVO0EpTatthVblRsTUVsdy5/57Vr1yGS
qN2WuXVEm7MgLllRUzo44ynWiii/6OGy7PrGPXx5Cp0C/c6DJ811fTjqY9e7qGmi
yv5ya9HlFoTTGt7VP/JRIO9e+yQMGr+qx9VWO5NgVda61ztSa9o/3pYMy6T0eS/p
0tgzC7r+WbfLDW+cvgGYciE3rxYVfc4bT+1gw0X52Tv+/uDCVRJxTLVjxn1uPhZr
OAfVN+8a6aNNK+8Vgaeo+bqUIJGPcEpiikzGfxkhyTOKG+u9ohkelzaNJasiPrX7
Lzks291ZntEl5DParWk9/VxR1uBb3VIf93Y/3190sOPC3HEUYezkFHFy5D1zjrfA
XR+8jHwKj2gMBoez2d++BoKyY8bXa9idlm6tZDPLClAEec6ehyD1GKKtfx1eI3ib
st86zbNbg93p9dG+17QJsarVliw+9QcWPCJF7J0LWXJfgzz1OgrR9ovl3wvjmAvb
pbD/SIl9jsGNG4M+vTT8m6GQ1cG+h8VG6HHijsdxWO/icCwVL+wouUfe7Td9VYzs
BQ/6WX/knPCpPqsu6xD9qW5jsVIBKVSn2g5SYUmKCtJPZQ4QdHQxtGxczjeXyTwu
/YXQ5H23/7+UL0Jn8sLEREwtQj1VCgxx5HxtgxMoSQo/uqN4qn71y4GGZ2ONriOG
SHyuAF9F905OkNzn8T2WAT4oHpAtl/rV0eYf7EJ8pqz8tzp3dg28+usVNrcBebNb
Mt3Pc4LxSBWo7/zRUC6pMZdmJQzBzQAq84FU8CiEDgfdJYNgQCW4R0YXHcDXeKIR
iNu5XY1kMZvQU4Cn2zAf7NRGgVFPbTMKSOKsL4zg2NQkOiQhEkUCxxvGS1taRLMX
FAzOIpw2944Nc36OUVng69l0vkKMULJYvjqO0810ow9KOKu4sBdXIWa56VseaStn
GDDVGmtNFAxInzQ5zsIqojkvp2JSSe3lIwZyxL6fnUMyOIn/DPK7dhLO6IHPHnap
k0HvIrBpeVnnJ1e7I0FV3NQmx+LkmQvC6gO76GuGeeY70Fb+ByH7Y0IUiRMRNbPn
QAwhFqWgdsZ/166t/QfpAGUn7gCeTOSAUUTt92f8VFiFSXion/bZvwd6BiMFELI1
0YUAuurFSQM1JkC3DU5YAFAebZccHo2ZHxRJVtD7gS4n2BNQqvoK9ooEjrxOtV3v
DWfNvHmcC16mYoEDbufHZGKS3aAI6PhCKseaImYGuBMmMhVOhJ1XeZFVWuq2fhFL
6goZBdJfh4gkAvaQrMqogGNCQVs8huQa+HsvfWMKBxpwJNKv7LjfW0YyJAbeYhxe
N0vLdvUCXb2ebzX5FLG/0CGB6pX4EnVya7RBinqWwOS3zxupJBBSQMPxuFKpVsuJ
HKGVoLgpsBhyzGxDOoWzWyBC0wbHZgR2gHsb3GERlssvJpuuIFoHqCmy/hZ7dzhp
X4sc9+xa0ur7jyQr7NaVA9dmqsqCqiqZ75kuY5ZnaqJAZrEoGOFnioDBtQRnHQIB
TMJctOEZAd0RQKOYpeKcszrTA2R23s6qm+WPObRnV5PyUlklBDgMEwxUj6HDaXre
sJGA6l/6tOyVRRrdMi0UjM/0muTVa9xF9iZmu8vYJKCWq5rCovJQOjp4uFlL0FVJ
q0d9q7lDlikjrMIIS4gsnEDBnLhutC2ulIiNKjweD2s4EovEQu+jfEn/5eZoMMIW
wvSm8quaprBtoDm4BzMSVc9FcSWYsYBBLWPD4FgJXmEyeTddiITByQZo3cM2CUW/
rHXtXiQjugTjhKhmEoDUws7fYbVUdHeUvhl5zUp2dgi8V3TYAhkqbEiIVeMtzo6z
hWnwtK6DwLuAukroXiKOPyJdl0HQY2sBUvjJ9CrCgiL0Djvaff4sonW2g80iY+Sa
ED3NLHNxUqzw//M5c/satBPMCOKF/+tpqfvlr2yHI4bTIEBV/z3cwbeGzHpIb3CL
tNKo5A3R/nJLJgKYkW2P6Pv84U0k4JyMNlIkZoQslBBUxt5Ie0LH4bWv+tUae5kp
Of1CzDsIf1dblzTUJeAg4EjAQWhiLgZbL7FYkwb8ZDVPqeZCUxXLkoMBCOs2uH/G
gYbDVFjBUAuzwh34VpNjsz1rSi4Qih9iNf8upezi6tDhPwesqCCmSr+HxgzevHuN
zfLzRnRW9iDsMWd+4NT7hytL44yRB6jyj6kTVCR9D2b02mhvNh6ugbi7oet7T4Yn
Qyrgw6pYS9QhX5lzieS58lzGbE8YH8B/8qogi1IgpkUmV3RDdXX7JfCEAPJt7bIM
5dRX3Ggae+E4lpz+L4Yi8zCoJNI7RdFMbMU0matN4fK1O5HJt63mgn1cHbzc99vy
Px2uLEc3RUsx4xeS8iADhlxnrfXiqGJqs0J/sdgt1Dkp9RuJDhiFfKZWWIDrpraw
JeqQMtM9siuu7Aiv55k3NP9ertSjlymwNrrD3qxPo32HuPlGCEV6lcB7rOeeWdgQ
kub9BTXqNT1L/RY+NGCIyKLhalabc2jVOsfalainyRapFmwQ7R+iccuVn61TYD/c
Z3tIuL0UAMm+FqaglCTM89iRx4V3lp3YtAMKLRIYGvi89moQ2Nbn7HfG2v/8aFMT
Bgs+l73mjsUyqe8jcetzPVt1TnlZwB45DMDoWweAQtBcJRiHY64g7FFwthwY9Pyo
gD+iSJE3uKpAolI8K9LhZlZu+LaaRYFp34zgpN/xtn6pXwUSde7/7TvpPESn0ct2
X9/zuhL/3PqQONdm28dTfQheqX84WBvtwAo4gqRZomLy6uKBq+jiiaK4laLkMhDk
Vol7apmgh9aY9EiZqgxE3gNJmHlJW5ZMdFDDNtfTTqUbSvX430zog+2UHNBCaHb/
G4hiU2mtedLhsAqooPTy7u7+0nEVB9EzVFCfW55ipb7uDO6/nNx+pdJZ24SZy1lx
n9ielyEvXmZUBukMHRzwpXe/+pRfzUEyHhfvY1oP14zyab+EuqNu6VYY/aS1RMvO
jp0cnR/H44lI0Lvi6wek/Dx3yK7pheGAL5W+Yt+k9m5fTDiJUwPB5Hw6yUfzfWzW
6vhpPvT09FF2iiqJa0v2PPUnS0GDrVHw7AWmfcTiPOU0MrfvwvnemUNzc7EBXiZX
Q6Z11/m5g/ht+XnBN5m9lsxuMcVyYdUSHaylyDS2wOuHhLKeq4rA7IJ7Ill1Sv8p
u/9C9orwOKHkK/BqPcp785glAZ6r8DszemJ1ID1/82wDrJiLcTYQmS/7s1nsQ3m+
hOXexW0HdXbaFjI6v1hgGFnBfYg8Nn7Fw+jHQpjAqE37hCEYrMPfnC/ZZm1TvEKd
jTWeSb29w2Uy0Ylo0jxUrH8NNiPN9MecUo8zC8cHv64czkRDziojS15mwUskV4Db
3SgcXrBzPM+a8ESlgXDE0hJheMTYYK2WOshnDzcAX5kC/9ukKMOtnV7YsxKrJ/0F
U0FrJ78Co6QPVEeAMedftmbidodozWgJryUNnX8c3BLOqAHernecXaWB3LpKvoVu
d8cSqQOnlLFlCysDQeVD4O981iRDG4xMeX1r1iIKVbcEhNBOnJVlSLe+O41jNn8d
Hq2zkfvCuTmu79csE3VfT+aMBrPPPbMJAsrtkmPshd3r0ErfKfrvEbz3IzYPhm1h
zjGmfO6jzcgQ3vVLziXNNNAnyBF4AUjWGnOrxb+3edou8BOjCgCvl9RQlRtdulIY
macezghK87a5XdR5tlTSh0Rh9383y8neePM0RKzEohezX5o9SyVMmehNLQ5d3IY5
Ctpp84fP13/U+wBh2xoPA2C2nwvMfgk9wMVYp0ntHeWNTcz36U3f44H0RuHCNDkj
+DABnNssFF7okfx+qJijt5begzJPqMHMdETKR/kHa7GBJEnjJbN5OSMwnEIKODeo
iL09xqRhe61P76WvpRBv5oIvnRedFqFGPczPbuINmm23OkVasbppUmgp83aq4Vj7
1jc4HmDC3wQjvtc6d50xrjCWkdLmZ1OSDFnoCnllCVQ9m5gaqD18iq9217Uyu1d8
yi7uAxc26rTAdxnQfB2AH5utlovF3gGUd3C1JgfaUGw6kLejwmmUBHU0/mEBiKYG
tS3wwZRpZIdL3jRPNX+DivaZUhd0X8YYGiC4TFRCW+QMBe9zvq67clOEwfQ362Cy
O4/UPpAvmfCsnU4UbKdSfSFNWHgeeurxDCr4/bRtjg+0O3W2v8eQECHMnCUZhhU1
2+RpvfTYWK/sJYlJxq4GUob6F7M83hBkhAmIMpZCH0+KjMXuG+DAdeEdbGINSvwT
dFQZDO4eAs8teSvG28DNL5vbz6xVs084vS92IReYxld70/Z/YovPIwOnaLEu3/we
WnFy3jcih9VN9mBiSTwp4cMjOKknuCSyGMtBV/4TyzCxe7ypBA1TDUyhEGCzPES6
U9VoLJiptxZ3SqxM9uRia7x9oSK2q/YcXK39A5h615JwZsPKIg5OCn7FsDTZVQA9
YRM6wGpbVxU97fYto6oYyETy3cRPbT1gMYHAh/7fA7qPIb6cLezWciCNb5iCFb1U
VpjaDOgSnreVlbtJ7/EI+xHzzE3WsDvmqDvKPf89QPA7W8NlK/d14Smc22D8JCaW
Y6tqkp7YbTrrCmqqB6fDg7VaUsDhBhCVNuNnxPZv2XQLKiijDuHI3j983PmhpSon
WaTc9QmOXEEzUoazFTUYUXH6h8j7ZvbFqKaJ5zbcLte5aOwG98EQMN8SSPL4Mt+g
rog76UOvkXwXWCSEhxuqrZEh4xbrLRdtseuvlK3dFo+SLCCx6xWWyEeV3kAE/1tp
I5c7/VevGbcRTZJ9wshkYH69FfBLBbcMzo9bp5pPhpiBJWAfPZrr3Q5pkzGjHBH0
d4Xr9Uhyf3FMYfs5a7P0ZnvOOPTTmfRavb6NfshUrm25nKY4tzgHFCyNaVqkvOit
khwSdSjZcBM4YGl3CdVMzhxE1zm9wt2BHbhXRK5jftlFBKr2T4LP0e+V083mIecS
QbOTDfTJ88S2UV56PKX6Rejbeknqc9veAqB3ark3oDhI9Nqe22gRBfAYeF3pF263
9lsslvxtBCETEZlFX0WfEJlqgZ1Xvl7wSdQ8QTH6mO08BBeXvr3lQfd0H+Z/52O7
aVydSXego/qm0LY4jlkwDyhXnA91Kht/vmFLA+lUsecZMNzE1s4kQxZdkYcJiGd9
ApvFzVuWKrDWtIQL44Tw7sUzUryfMy4bbvsdvBtXhJrQk13ICsz6Rx7YABqs05Jt
VoCpP/l4VpTPR+0uGXxLz6cQHBkVjU+vBTZhsvnD/egFSi5Z3Sas6ZI2Ynujata1
NxSzl8gsw6hxzQNQsPOt0oNGSoQyLRJ2kdvCTk0MnWGUZ34l8q22OCXcNVzKXRM3
RYIptToZmZt1pmkfNCDCoMCIIcQcGZE/TztsipgCegheNKOVLkg8AbSP/va17YYC
y3jPl1DDSOciKa1qZzSrcTTCz3Puo/07MU1E8TDmZStbynEs4emxLPsxLyCKJ+MN
Jt5pYxL38HrjCOGrII/L9NLnSC4PcnTHcepkZ+MJcRFsAkkofAfAXU793xG/I6ck
UIzNK/w/P3preycT7rHG/3dHpLxh3cgP65Z6I8/yZ44FXxlAU0efJmBwAwAdNjeq
uURgI4puL+G5MboYFIplu1CZSBUsVeXt44plsDBa9/AH2rRhcd+RJ0SKkpLzOxCC
dsMheyAQplCKSzFXzhgRv2qSJ6AM0VV68SbHWEN0z0P/J37qqSy7NstCbBK00tyx
ovYnYSdvJZnouJA0XvL9uAiycXAevtOcXOgEEON4Lw+AZ7kcuI9HHU73QhaOh40V
1a5nZRc+pU+sosbQIRrk/I/NgCHLuTPm+V6LtU7K/vYrHqkAvl4VbK3x/DbSqDLD
UAfD6Sph/NDcRIQtTLM8TDg/CYG6X0BshIvMPivDel/jsAX45WmJOGg8Q84/fcBc
a6PlPW0HDFSDjXJy8iOKkzFVRBYB1wOvfaUNVczl8zCn2ko1qqJkPGr7fq+E7CED
yq+b13uVzjtQ0tjUcMtUsnBVHAkn2ucZGVxUeDSA0HmsDuObQjrlxSQUPQ/uOQVO
KHNwjHVebGdMvjuzyv0cx+op1suWCxZ85ZloSh0iMGN9sELof/yBShg68pR8eXie
TCcEEIra166dc84apPkKH2KIhqEtsKY+sAh04MhXqT9Qt54uAFE/2+rf69OoQe8o
bib53nOosbjSOqA17FXV6869vZxVRwJsFKlLbC+XgtgcgHov25imOjOmXQVbPjQT
touTKSPotsFzjUgFgEkMsV/3a0deSPVbesbXWwwPy3TynngDpKA5ERFiw9Kvk/DU
2yQNXyVM4sjTM1OPTieWNsVrZedLErQEG876VaBT45VX0Pkx9sRFfUkMiMxJ0f+U
nhYK42/nU7tsn0JKA3kAbr2R511W3odHUprwcaKFExNtaK5JJG3sPOjLdBNVEuZW
WnJRi6d+XwturJGf16sO4AcA6ijdNGTcUR/TF3TbbJzhYTYC+KeaQFa+3RsU5x60
CZC86uUtO+y17krtVNq5qhv4lvbWbAJt2JB6xu27JpVbS/hMKgAhdh9M36lvkoY+
CM+Gi7wSpzZjNW/vfXaKipvTuf84qFfhO0JktwV2eMFN6jlVaEMYqyEF6UVH7oRh
p0Ej+sA07L7t+/DIhCVeitN4jeVK+VxvOmU9pQBNOS06ITOwefNpKzfNxUf/hmvF
pGWPc17yovyEXIE4a8JmQcBSbEzu1tLNBHGRQIUlTBYiPd1jNVk6uzkPmYjBYnp3
37JKaFMHoa8AzSI3cTekEHojV1aYCL+4VNY3BhL8yNs49jPtIIarVDxQVUJHkx5C
9+TYNyBzT+DT49Ltfz8z8bgwLS3s4RHAhfCTFT85A/4nCthrFFLM4Cp6EyHPVSac
G4TmYu3fS+LcnmdyOBc3zgTiD1SYokjho+MCPofQgJevN7ScUzdWVL/vzRo5oIrc
iZbkP33/3Uo7jsQ4rBz7cVt8tzeqJdvYUE7kku6SBaQN/vwpqBlaPAYeArAeWsyj
NHUhZxXtX/Y+TIKJp85qXPusN+Snw+7cNkZGsWQrCZs6QHUDpX81tZ5VwFbgH8I7
RTcpVupo0Q7gXH/60RnnplZcDYMLPIc8NPygzbFjCDezfJO3ZMctuhZZ2LYCsII1
CmEwO4zKdeZqbzQVdUFcMA0zJS4eu4+2pgwqEwmTXnBoJadBoAfCRHkuOxb4YbPa
j3KV0qdKSMtaI/IgAlnTQpfgwXFZz3Ed18WGqG0SkMt60oO/s8/D6t0bKMxcY1Lv
TRsubY6CrBnSrrQxLlHDQQ6Wu7OgAaeULIJrImZIEJPVKV3XbuekdrZSYDOYzTao
TahoV/fZw+6AK9PeIRmmHX59rMPB+4zkhMyllyithJUw+rf2b/T8b4hJInS1y5zt
Lixjnea2gY9Z+1hL+uCjOM9lStA3ldkfgARAb4pdmdZgMhdkblOYQRN6qRG9zYse
4E8hw9OQBM7NdvVv24H1TuX1aEQgZaffizhsAnaBvzL4BZthAQw67QwX9fZB/iHz
xkImLjmXuxYfOcqBsNUKMaK7jKsfbLvu9Tae9zWImNtcl1drJcMFREH5kfKT0diq
SOctU1Qb4uMyCd2UiTjV3s7LWIzSehRaJA6rBEhbtkQzK1AkLxeARrqx+3MU26oy
u9d5RoTekvQ7jFlajGOixm9Og+504isv9mcv4jN5da2t+TiSeHpRYP0rCi1qQmuG
jOgRsWLB2hZ8tknI/gbb1OatGF7DADDae+UgJ59cDyUNC7RGNjnFByGOMza5fOYI
UstFS0EDz80tsVF9H3ExtipnK/1OXXRM+0uLWWl7kCbcqjfUWLzyu3mZ/vJObqnc
HxEFKPi5vRk+qh6DRPFmNrdBZ1G3rQS9BTxU+vrajXb6DgHx5nBNVIE3//U56uxp
CIEVoAzBmC8BXeNs22T2Rc3gpXcQbjzx+6HtCFh0I5aAwLpWsKgQOPvg1RHtK2Yk
YDhFZYXbzejmc55ddx/0KD4GIqgHtS0mS1yJ3Zv+OMbMlqJkqiEkAlZiKWlmKnk+
stDcyRiT8Kocm74grts1vK1kAi3qLCWjPKYb2n7JANdX/6Txi+/WoaYl4wFZ1XtJ
BMQmemdGTqYqDBj7IAlynlV+vwDkOeMcw/sebZoHy9vRwCHfmqOWpAhVM/oEsPd6
Rbh1xgs42McfbQUeZlpGWyL+VB0zKsCoU60CXAFlqNtdFKbsmU8yJYcY9iKyV89y
4WFUXxE49sjg38soOeNA606LFPEZqfPpqHc1/gtquvv+m4DthINCRXJBVS3PIHId
8A4BiogC20ktrCzd05CovWNwzqdQnIxm1s0CyIxYWxBEP2MZzuzV9TsEfAIy8hCW
nXWfN7NtyRsqXmUQ7AAkQ3cl5lxvBz6BTT/BnuglUy/EI1u6hlkrlNwvLy8dbX1p
w0o2f7UhuFV78Ws3fBsczfemDi/1XZWp/snnTDvPuSJQZ715lNe00gedbgD6Kt40
4TnJjkDYVUvqRIH4jRQFGOcxtvyXBMbUvCpU+tJmFzu3+/fggWOolyTCsBaYQNXR
MXU37vVqUa8WUdBN12fv+IVe2klM66SYqaQh+7Am90du2Hh8cUtp+H/NXuQNy0fH
3VE30pFrgsOZQCbI8io5fSaIJOFSGbdPM1CXOzlltcbSQKyLA2clS2kL00lba+RZ
mmAULYkb2iD4C092/NFWzi2SKtoWH0Bf+7HLkwhMziuU6mHIjZa7LjScWMLhLNkW
hxDms8v6bd+Murp6BaLYoBV4P4Il9ebAG7FvKOMH00Jn4duy8erHOmFqJGaSL5Sf
41CTW6wUN+eokXG3Ykf4WuDeUe/V3jVGio4eFxQUGs28LbCT5MJgGT907sFh9BhP
L44J9DvDwJesp0YSJ/pyBmVXe4wRZOM+WHaxhJhlfvpPJpXGscO7/at5jG2DYiP8
JqQCH2jjal5DDZOI9ZOgH9yGBzXCEv8tWe2e9TNkbk+xrcKPy5B2g2ksGpwkuXS3
nqZo5CQfPdo3eDb/o4zqCwlJWRSDq2njiAqwgFupLNa7XvtiVgScHvOEJl5QMvFw
1woy/QVknvAGiRiQMwqkBAEMjx4h+pChGbwcJW1zOseKGbbACHY1jcnlaR2Q+InG
WA01nG0YkpdGEH4zjLdU4DNId8/bIKPAVuc2KefxfZZpKfHJOSfvqTcfo1i6Iu8+
nOHIaVJWJSzMb6d9rkKOVc1egf5cadJysJ0IH2Tyn7oq7J26pU3lD5W7WeDqGGXc
NUb5BI5HYTyieEDPRIk0Uah+9H9Yi+A3kHxXlm6CL7h1FnguLzhV73z8XGu9pObh
FK3kCnOkBi2Yibd3HXmt116Qgz57Ar3IAAAyeZMTx82flVUfktwHAbekHgcva43H
prbvEHbI6ylQZlzkIons5yvLnDevb9RRSZX8UYRre6o4m1LyXWNN9mhyLLfvXNbp
nECAOA0NuYPvDwXNvB8DLKGuFad/PIcjeujtxR2udGM4zv9DYpHrsg0uB1/aXALY
uIhgWF7HYOtRLUjhaG6ZoTfmbPnqMI4iG6eWMf52RTHkUF57dHaQ59DBb/XYDiN7
j1HnCsTUGAp5kpGQAquqb0XdqP2sWaGviDyIxae0FN0gP6Xw9flL1JrqC1A9BJUA
WqCIHQeUdpscYC7asHe0KvFpwyQnB8GvYKOr3DExXJmeV+o1o/YX5ySVgFESDX8O
bLQ7i6vuTVoROPSA/W6FI/ZVoHoJibfWgWWdHtuAOamjBMzWdtsP/DrJM42QdMdR
/ARhxDuR4tp2KjRvudwewxzen97uOoofS1IYdX1vybZTy4Aiq0SsV3bRkW2QDysv
VdzuA/5wM3O8kzvUNuCxSG8ZJ33o1OwNfLZXGtxmITjKoSgEfr4jl760LUoWSJK5
bQ1m8/9C6Q8MRIrG++a35k+lYjtuIBScHcO6eudVK5ZOvzE+IIlDNjUMNAUnJqbL
Ebp87RL/xWjNkwXOwOulmOO9QPcdFAcbefZ8L9mQmQgAre94PGoCYJI7W6aSMG52
z8PsQVOizmSMNL0VP9h3LIG3z1kU8FtuuC459WvT3uDg6AAijF+GESrAh+4/Y2Ej
H796vbQGk/Pn1IXIMkXeQXVH+qC1KE9xxjnuGCOc9hQtioRCvWb/tIoarSou9uZy
B+S8jFHd9vvxGHi3Xi67ofIYq9OyRhSAD06IzoN35y8QK6lRodjnJSPiyvJkrQru
o1fXxYvna2+gw1tiYbRNCFTkwGus9PjdXN+KkxSNqPBr+OKHBGIsH8Xv92u67fzX
syyRa/yDaUbnoadlBD1z4kOpsAozqImS0vSHNORMDBOW2NMqYyjfM3dAsqH06dHQ
aX3lYJ5+Tc8kz10oDcB79bj3vSbr+CnB+vfhqXqyU+xIzHdIPQHTYd0C8nnYCp/7
TaUV2aauIOQ506+h+vd7dcSY58h7OF9O9zwIB+3ZhseLDYQssH4GrUi8x0k/VJfp
zo/9uFZ0fih5z9QJAp3pPqzbdQUHqpRnCx7s6yYe5SF6kTB5olEeELccpUhL880i
qwf7JmzhOeMSItazggW0yoDM+ZzExojbGi5Z8UTSNC33qrZxZ1AGA0v9lNzSQsR9
mqxWtKOf22CRo+C/0GPmZ53Br9F1rDmcT4gmyz+Ud0SoB8wBGApRCZYcss2YD1HM
sGcXf/65xoXvuKBr3LlElpDN94XcJ4kzyFqWkwDZu6O6IE+9VKq5Lmbr9DmDnrkY
HPKc4BYnCUbKyPufamLPWg9FN9MNyRzMqwtUWWdyOsz4VwN2Y58woVdXM8XlfkSy
Qqitbzoq+gL4dQz4MqzuXJL+CwM8B6brYYYBxSbJI8R+EXh+EMd87eKmU1e89N4q
Za/RmCyyZQjTE5hE/CfudMr3wTAjfgkYWPbuhf12pEQgayQdFZ50crem3E1SEQKZ
odidfqQ0u8SINWvnRHeOPQt/2R6XDR2V9b8Ytr8ZXgC5NBY17THhTgtt/k9irThR
0mnxiOAWIafhNp/tibN3uuZtuHA3/H8teRnA5UrhTGvHeaOmN7BSXVjUDYmT8y+x
GNfAHUsXd6yA8u22gxpRqTeLTBJgtSx8Pw518VtE8kB9UKlWb7lIiWlfJ4vdfkon
CghhJk0y9CzdmfcgBPvQ/4+Ib6fcZfAbUgAxhXiDtOr4Pr35rTC76v5fXD9R3nmS
qxJcMHk7n7Xd8kOrx7AasPie6CcxJPXBCH4ErvsD7CPKD+BO6VNlSs26tLcRaJAI
gRtAAf16zG8RI4FMTi1JFXY0xccjIvQ2a9VgTc3Nc0LW+xpeIOwwGg36fWckp0IK
9OqjHhz0oRwA1tjlR6fULTj5/9y7R2/6gOoEJE3eihGGzUMyfE99PoLAobPYCr9L
8fDoXcHeKr9FHNBwL0/TJ1RcD3iKNO42aV3DZU5qRe6cY6ZdGMoDsL7G7xdy+HZY
vd81wkSBO/+6dOgWXce/OkPkZcRuawsPbWE0QZlgaCp18r17iFeXubXjMKJliyMJ
jpFzEKhVZ6JAZtZ+VZVWB5Pn+UvsuGnK8YPIAi9n/gTeAMJ2NZcGBQC+Ai0PxTSf
tjvwM6GbMQ0tStx39z4EaYACDlrW/unlC4G8+r3yMvYXR/HO9Ttb80+XXkT+UULH
Fi7GSoU1sRvVnooT9b3RONN3SQf0ILVSM3Cwl6S+FTMU2KRFgsv1kYpwUJZGcT2E
QrvB89k/3/9QO6iITBPnCB04DgjzfxIvWMifmQSdv1CoyTu5OXkwcBLO1sqw/smc
tlx6ppMsACzymjRajUJw+Ndr5ULhYSlu8A9miR2okIaiL90LjQe15yA14ZOIVcSF
LXGRum7CvlahyJkD84Vyt+EfO/LYRVxHyewhs7NPWh+79x/At28rEv/Rkc5nbw7Z
om4/bV1Sh3KY3UtbEXtql0kBawxkNOm//HJXURlGLlweK8Dq0KVSHzgQqA+7UMro
iHlxZVbV0SV0XtcAVwW/0SWcgvvJsJcitmc3qOLBgo1p5mOotaBUA1DE+r9QI+sX
G410CajokdvkouBQY7kCBxCshcHMw+vUJTUVJC+czW1Bw7VoXbe37yjfCtNDsX7g
IpwhvqnkAHYWGtB5yKtVZsAORKq9hfYIIv6OwZz1wUBmqqBVWC4r+y01WyCBumnT
lXH8K0GxRfpPvHndONmo4i3Hn4wYVuSql1CpwHi9f2agPRdD1QDrbuPYta+Px3lI
Vgo+awKLsGxk95nZLGK7t/csRlUuwKcSXwooFwUyG0O0pUxe6aCb5WvUqc6chnlo
9Ii61xxnLmoiM2973nBL5PZpDXY6TYTY78TAiyMGZ5l5tHk+QRbmea+Tho/vsei5
9mIrBvA5aKXDnhWyWZwXsM9l/tAlLK+vc6ZY0QPinW/H8wioFjM9dTnhphXYuSM3
hu9aSflirca47dmtimGnamW73P7FTxMTVdb7bhzXdx6Qjy08Og2NxGs6dzcvTTPH
hnzZoK7Nd14A6616DpG5M/eDBWECYVA3LGRUTuU6D5CHorxakmJvh/F/XWZpgTOj
Uz75l25CHS1k3oAGGQk8fjQa1rS7PAHS9j0l1ZnUkLq+BaCognkx6D2XyVUfTaqR
EJCnr1PLWhSfJzxX5QKco16nlrYi5Zg+nlUQdxKFYl95M6kUdeLiAsZ3Joqlxbnz
aiCeUSY00xJb+jIqqOWgCHpMlVQ9HBRJNjlDrg1c7VHoMPwc7AduwyvWEVbn5Ybo
cLneY5hmqUZMblqkI8eSB4HZw8InGzI7Rg3MF7YZEtaMFAURM/MlUQrcFEk3vVP4
7oLwa0pxq+tPCvtZsxzN/2G31q0iyZ5c0/2yFVJQrpgZ2Wm1ujft1nFmNC2kqw56
kIkyKBappHr5tAzT0yJVV/ZjFEZUboyKfy/JfvS5niJcEaaLAYtjb+tKHOe0Higp
OJdBMJ5Bhlt4KVzuhGf5RIOiUdR/Gruahh2vexr3qWR1NKivZwLRv6+d5eygGLeE
Kc2tM3r9OEt6R4qknH8dmzGPPLhaEbE0wOkg5Jvg5/BpNANxTt1BE622MMj3oRxl
xFpoXtQDtpM2uzUQW1to9BWBuYLDEQ3ATKTntgNzU80msWGtvZRl625NiTaXrR2q
Fo/ewZ3904ayy+4LDBgrgUyLoGkvq/z1IZEGez47hPzXb/+Gozcyt/3Ibex8uHph
bwKHO6/NvR/ubQBHmi2lwPdbv7Otv3YIh1Vok3PgM8NEhSEAoqimzIsD3YVmFuTI
4nCht1WJZ0rEtDo728TgBXEkP2gIVb/pGhlZ4zriXrAERB8yUZMTOru4mEysKq+y
Oc0eccVSwSE/2DU0xMHJZ60k0RHqS4IEM8PHra01e4pIFX8ZSQA0yC65r0X2pmR6
QEZBgI42WpZQObCx/8R+1MqYb9ZWOg1a8+xz8DlCcqme71FmB4wMdYiyVPnOl41O
XP46WKtNw3zGeiSQl71SDoC2cGWrvkZqH8IBpQqGT23k48b3PDQCwNr2HdKPkSWy
AqvO8/zMjJFTArTR3oRQOTsIITf+uDG91yDz0ihzXz1Rty9tri+wMbBQtu5z9R12
YXbZCO8LtRjkaCuefLZXNE2HpBqA+DCPi3+WdQtG8IxN/3gcVXy43kG5n4QVzgwq
NRYPjMW2T106HdGLeUwKHOI8/+0cCv82O4glbRuABc4NlBAFy0MiMA+gtrxdUet0
5bLDXipVqx0MVcIYXDYDcT9pu84tW8eoCMfW+uv85Khkfwyyztq1dtlc05eWzIhJ
dZiKr9tjDy1tMna6TkfZNIfvt3+BItTVAZ8DB+usF0fy2dUYGFRP4vXO7awKRANM
85bNq8HbfggEKyTVWJyY3IEboKFdyF4MiPIq8kZ28sxeeI2nYrReHa6EXqsPyEDv
RiesRYmaSSNQ9zvtBQ5T20aRAo3llnkgnv6WbargKTE3jhdybcWuZMHTR9S5L2OZ
uPx+YO+xFL1e+j1tgQ+6ONkr7CQfgF2yAdDqXbuf9x8ujPEmbL66Kxl0QpWZg0kj
kuvHysDccRV3eMz2S0zhMmpMinsyEU3vkf8HYUG9PoVtvjdHSVBcA3r9zqrWR41v
bC0gPFwZImJFqyRPD+10yXuWQPOYPyrSi929l7SFkEU6NPL6Rr4FktLVNN2xcpk1
ejParQmkT8CapFm5OvQDMOf/6PhgpxQ9hLY45YvwjQbyjLI90uQYomnli3azfw1A
o+v0EXP6oLPMd+9aPsZqKq7sG2ewKKUrVS03oRpMKdc2KNQduUP2UkVGqkQK/quS
6aI449R1gK6YVgMvrwnpkS9yz9y+yJITcU/guNA3CpvdS8EYxbu7mJLLtwNvpqCO
fatt//Kt2SdM1E5GPtBhOM28zPY5R2uSHMx+Yh03EwMIAnwjPIwQ22+h9MTeGDZc
ZRuUYhMZDhRw/xGkRER/CjNCbBlvU4kYtITHc12u9kbHh/MD/tgToUDw+9j3L9mY
B/mrJOneSx/UcZ+ZXspwq09AysH1YENsvK2Nz4jcbT2MfRBjcuMYcON1Pa4Ml8vz
Ln75uRtPsM4jr6a9UWJ8YGbBiJ7b+EKKkRR3WZ7sUiT44CGZ2U2i4fOJCwKfYckF
oaFqMejv70NC708Z9Pjwv+IgeWr/fhJaljEEZ6hDvJU7uYOlP0lyKt598iyjtVPL
Wk9vVFNXspgKfxfiBRqwwGbyUilJ73D6LzhS80Eft6WEVUg0kVkfvk53CDmh75Fs
FoEOubI+vRMbHW+88EhCU2ogNK51iqTgr9MyKvNVOL2fUsPskbm2emijc1HAcUjb
oAFhzTH61NbS3FJxrMk26SeM90L2dQp0hL3d9UhjEwnIyzHNyLy5b09O3TOLuuwE
uMZy+0rLGwRjkzRzZcI6zRTY/xABmU7r/VIzw7DarP0pfbvth7Nw/Qq9SghRlTKK
y0H1dTNno97QBSw/MAjqCsnf2+UWBgUBLeI7KIVbGGd3Oyq+a1l0dgH3d6HmDZ/i
xM8jGIic2/ay/qe2m8uz/ldEhsUBFCaoHQwZ/O+VdgyHdKrxCKSAyTnAMKjO1El/
3ikMABa4uCNCqARSL3gdm13mZCAUcifIEc4ayw0zJ6uob55k0szJgAjyohMN4vm8
RWWbWQXSAbD/NH4wFdG4xA/IcHVfADq5sXI9TyE6dWJerM1/WAo2Wpg1c5T69LcZ
3sQiKQtUNfuR2wJzN0JfkxOeAD2H1KZmGkiaLKRJYAzyKoEEXRVtcmqEJ4YXDtNx
CVr0G3Hjn5hQn+Zp9kXcqCMCX842RWw43/42vjvJPW4Kul7rPSb4ywWiGxN/EXGL
Nz91PTYh0uxhKa+7c5ws8RfH7EdHXNf1NsBWpJ437hVPcCBJnCx9RjzpV8VvD+0u
FhbSt7RuDrwdEbjEzA8j/3IKBm88efwyno/GJw4dNmFPGlQeG9asjvuThXvaLGjS
A0mCQmGyprXH49PzXTDv5wZK39/gZW8zaTVCFRcxAhdOn0xrhLTrRP8iXRShBB1Q
xzppm2/bChlNq/cGWMqn7iQGvtn9PrfTeyUypTfJ+SuRees1JGljIMoUhlpAB5w5
L6djmxOlhyaz8r5ZpOZGtW/V3tj1xAotESbIN0SBnTccTpVLpHvcEdEM6nqCOVVJ
0uAAvWEHLmdbkuLScRMCFkenXEsj8WApkx4HMQfpAR/Rlsc45BqKgK4p5a0C+20g
a5kjXMwWgTZCGq/82i2VCvvXjaM2ns96lmRjaOzJRmPDy0m0Hxq4iiyBlzL8P6xi
CDhWFVHLpF5vzW6Jbf0eEuc39L1vMfkkrVU8q1co+56voVhqoWVOQN3pfzgfoESg
u1PUGq69lm4rsjI6DzceF3q0LtJONImwsh9WDpRP/6Dw8bLYFUqR+J82Dh3nArU0
AY3XGOPesVca1YpOH0bhH9dC2yQBGJI5CJa2jUkMH0Fy23qcE38lTnkBUWfQlZi1
Tp/OkYrd2VgqDNCMglvmDRIEt/BPVnpUxKkoeMAryBv4ce7ca89Gl+x9UydkKyu/
tGuUaEP3qzBI5qpsFOJFnk91f1++9zZGz8G+P9NB2r5lKNjdydFs4MKVTRbpx2UQ
6eYmEQQ6FgHreMnDeFjbW+tq7mffFAb9+f+ySBDVa/wXMXzKAux3/BF6cas1buQ3
QmEkyV1OTP3bSbO7V4TKDjcrOM3pxMeS5og86Z8OuQ7zimJHZLzbzdHm6cdrS9BE
/nmY0MwN3Lqv+GMiyjVxRxOpNLQWyDigaKDF1xSFqAaW3HBV24pU3s8piBR0La7w
sfolUBYDkzu+U0usX5EqhYA6Zej0HvtT5R5wab4nFeiBQ3pZ+M98taHSmAuzlQjV
s/kNifxvbMmDvHwoj7R/qiM4sMvZTcpgegNlKy/AgENgpH2sCBrQ9uD5fGaVmRnv
GHYs+7XoRVsKWRXvRtlMjSCFs7yanOIrENAxN8Iob9I70P7aAVXDRj0J422NvCav
VmKDYzURF6rpMLs7HneGpaAGQmtA9ZI1GFjgQo9TFFOc7YFn5HvWgq/Jo36qJ+ke
Z1rdRvp0Lc1t9qQZ6iDUd53KmEXHLB+cROpDyreX0ghU65VjZYvLcYzOGswzJZPD
jak1LJeZY+Kcajahrgo3DntM8p6HHt/TaOCP6B+EzeYE7xTpQT6ztDsfArQgcNpu
rOAR3TCCju5mghBQrpD/NfvxETSvi/XXcCJBfwdb84MxA7bsST86sxg1E1ozzC6c
jnaaSSfDADxY2k8nFQoCOZT+SdRsZX+kgof/j6c3ul/xgBm137FeRO8FHvIDiqhS
8aPTXv32j3Eo5Jz5cwNj2+0OW39H3hUCgF4L0CPQuJ/XdxQbZHxTNkLWdw4M3Lla
neGYoZwgzvPGDmXAwyHX0Yh5WZ2GpG4MCcbRqdtGvUUaXO6mkoQsTvX78AuoGgVc
KZdGjLn5cSt7NQ0pc4qRg0GBE5dMU0jh/vR9SGLL43zwLI833fgabdEZ2Pr2SqIa
sPRUC7bJ1h7sI5JxdvDN2ZuhaDhlEBLVZz0LgiztnyQ1t1/TmpEZn7A0fT7kzeMQ
or2dKzrCjQmdA9roV9s5PerQGLfQp4cyq6FvQ5ZW+FGjdw91nu2FK0kijd5PaDW3
+irx2HFMeBSo+m0y/fYdFb8B/CfR3m9eJKpQPSjzDjmN1zYm8GnG/ygK3oPf51Z3
HWjHkDoUjhXYo+5ofDhe8bPGcFtHX6m5Rqvvab3OLjC/xjwOWsvQNvFEnln4fniC
G5+6oZsmDrYbuOo4bsrt7c5ZE7WvoyrTIvMmJMSwp8yN+XiJgPH06WPHm2JxhfWO
jW0/IV95Mj1uTMbbXARlPRH+R/83JF1uP8H8h9FfSfYDQk/cSx6LIabplTJsGgcZ
EZzggQOV/cBB89RR7zV8MpO0CVPk9eUwk0/rmJ4XO070nHbXjNLaEkjJlVdKwv2l
JpOfHrYs1WRMsnLXl0IS+mhGR0stTxC2K4aRl7v/ZElC+w+kaT2Ve1r8a+yXRsN3
cS2i82MgGmalSxMU1ZR5OnIjEzKZs5nUigvKm1eAhbMGw8GpboUYZmDvpSpRVx9k
YzT5ghWxsoXKYx4IJVn8xHvNllKFnIpsJ5HwC9dln6XgXGbYWk46CoYo9MRYPYtb
4gfmnSG4XsvRh8PbgwflElLxi8u2i+2+VGYjDW1sH5ZZl951q+aLzSzvJNkIQJtW
Z/k65IkOgotVgfWTH/c+Q7Bl+vqBPs4SFLOSEBd6aaqlnwrZW0d5AakjU+3wdZGR
8Wp1oCu8X8dRbqwS8rPhkCYziT6vecyUXQ69AYaKjUcBlGt0Noz84K69YghEsQTO
bu79uVAwPOGhHJ2odo8BTek7GCkyOixPDOcQa4W3zBJkSQQ7kkDri1dHuTCwTeNU
2/cQLg319f2zMg0TiEfduNqcRleh+Dr3be9g9O+Wgg7rHKzo9z7D5JRoOs6/cVFw
dHASP/IWRjo/0Au+WYCgLds77Kl50dlepgJwyDi3n4LIaq28881MAH0Sqf8let2m
Atkh7hOqJSxdYzXTLTGwoJCJANXwNhDkvPhtn03copCIZswGrmC+28+KR77o7Jjt
NhI2fQo9JhEjPrgFGv4/qinqOCHwxHQsRZGRhE1hgjmjgF8OvX7nUEBVFr0JxaJV
v7YStvsrrt/lX2rASeIoxvUHVbu92dveovR+67B9DJbw8cbQMonE6Zs5M0iqnYEw
D2Caq4RNNuOiePV5LwsLgupVkusyPw5Oq7FFBX4K4xbm6zs04Vj+tPXbcCpDBXrE
EEf5UnV3VKy5ygVqQO2/bsKjDvup7RowPRjUGkmeSVuWzUwxVmAq/vp99x+O/7RE
Gz/Ep3nYBFUevSIJGTiwcNJ1R6qK0AJpVHBNUW83eZt9oBYH0zuTepLo6HvIXsKT
NjE5AGdMXC+SpXKxMNAgcPq3ugxEeax+r//xw1eHQVXuvmjVIttZu/00RUlgylTb
Cbd5BM75eodHxJbHOS3eGCxtR1ftnco7Ul2enq8Bk+YavaDhSz05H1LIkuUnZyiQ
KR80Z/Le1R0UsLC4kp7fPup8OxZ37LOtosiPtvweBVtybhD9C8iCDvnJbJbZYnNw
zP2AjB54E+n8/g4XY8quuYU4yRsk4p4peCHtVkPEYsdSeHzhU8F5jB66cp4DIV65
0pk6pK1fPX0kqnHxVkCQzc0dlIgcL8uIdxZUaIREX5J43YZQLGyY7GhMxpC/CePb
oqBhm6h1eSNpy7ZhFLGStCW5R2VC+WAqENI+lSfMsb3uLX9BvlJQARpinp17qebs
zZsFOYGwKJhEk7rfJp2J8OgX0sT372o4pUMPu2BH791LM5t/rJpNp/y0bjfugdXx
wPFmtPdmXZ/t6SX+UOHHc5NdJR69VJrKz2+Mb8iL5oo0d/oErKbt8AexxOD0huMw
Q/a7AC35dDpk7H1j3+wT1b9eVdItIaE0N+eCqQd0g7u4LpcYSv7DCSDvljac4Tgu
E6tVJKYxYyQpWFeBuokwGL3HXplqPos3SrsC8DkWs4jRAz1uPcjlUQnjxbh0i26d
+gLaD+04jHoeqH7FnqB5D3jiSle2cammFuWsExvTrpC3gejmmegNWTYeY/yo8YM4
5E2o/76YxsOPBYHs8hn1S7awaapLxwukp6HTeuhtMNEedQtGVkyS6WleBuya0XkS
IZsfS6ti+0AwXx6zTPu6vySPHGmI9UPU4iqHcdh5+NH3NSH76VkUWbgsOq9x2HlP
54cyLtQH2b9X6ZfTF7tli+I/oLiWED2Q/5Bm3AQpbeDHS0ULK675CgbnyGoKlH/K
/LAP2lEZHNetCK47Gzd7qDl1eR00BJi9K7LH0S7BSNBiBh+SWhenHxRQ5dsjnCQ0
2x9uZb5Lv61ZQHZMuhh32zUGu2+iEgjJGo4DmcUW6/e+u7wf3Pk9kgXBsIxlL01H
`protect END_PROTECTED
