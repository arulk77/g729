`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SSKYzHP5CjBhjRbv3FJXEfs2PU3Qx0Ez2zPkafZKgDdB
sKpFsHMi20UondsV13NSR7u3rxe0Jt6bgf/3kgiEOHT4tu3dDcKGNGpQ60M1zGrN
VwL3wDO3iAVvqFU3XLOLCb2//u0rNBVc5k4elY7O7yuEYqMkh3m7EPyO5csp2yqb
/hgt6lf5ywVQhNoEtmQU2+UIcppJH6WwJAEAVhU2rTCXiuQ/pEc4jVuFB0OsDiKB
If5r0HFDECRVPzASO4W77lqihJoKK4eipBAos8c2tdk1GQN+wDPl1rJa5vHrPn60
+HWa7doZQFfwXpJ3etWKzHLAdKrPH09HYEjf0ngvvm0dgaPoupFd0d/rP2OpV1Wk
0XR3eyLcqZ+/WieTIb5/KPJqxyNt0eyR2hYmFXJOaDunpI9rRE1PoyVhbq4Nvyp7
UA8Xq5lyQmrk6uF6g4/r71k3y4azJbSwqVtyBpiDhYcpgem7n2BMjzzI9IbrzvlT
UfGIm+Mp/I59DmQZ7x/OF7ImYgwpvjp36vg3xOR8tznqXWPtU3/PQWDpMjKXR7FT
ySCvd4IFLGLVeb2pH4S7NdPOfYMoiWJUnjGjXtGrpDXDY5ZK7jnrBrYhC0g6y8gH
NI5I+jiXSJlHFXLpjkohmI7EN3KngBCbr+NYXnVHVtZFyRLqiLHGsK+XG5ybWorB
ulbQyy0BVMQFWD3Anjw2gKv1WH0ZfsVn6a9aD4kB6OkmhrNLykB035gjaEHLXWeY
JWptH+0DEnHSRj1xFgDIiYS/jNUsXkL2n2hzOfW2rWTne1RB60AETojdU0+MSKro
Wbr06DTopbWpszcTbsc5qXWJRHnC7+qnly+abPg/UoAPcdaIZzjWSfTc63oMFrjO
en1OPiqnbwlmFvXxfMzWFeChPK9kwgGbOGra9RlIqu9me+jv4gvROXZ/P4+H3Gn0
54Am4kYfm1e12YOMGkIjQCU2VOiODjcvOqXH8y6CRXezq5P2nUvCi4DbtH2FPdWf
fWoMOybT5oL0ZberP6oS5aBljcclFDl4AezVaHkf3YBxo/jKXX1rAaYjd+L6LKwB
xjIFtJmOy25wFS1+6ryHOp9OUfTWXvnogGiX/kyHRk2FK2HhTIH4tFed6riXisao
jX3i6gEyHX0Ca0UmAjsrfdIZNPIj5k3cU2bppg0Cfp22DDh+cadlxdOta3XA6XAk
W/JyHL1oCoDi5AXIzD70XkqEBiM+j2Vniw5afKXq4K0pAbKsOR2DwGQ9tUp5MThn
r7CPbu90o7Iy50GDX/twgyWlaSvWd7NULzBGuxX05y2X2lkb0bWwRwQEeP3bKbrU
bp4bzqey76VvlqJNYBz+mgSFNNEr4TgIe6dy+b9MZXc7z9PRfzhnVoYmx7ayL6T9
2htMCU7Xoy6giGuCfi7U51YY71urvp64NvkfT93jBirvQ/VpAoZRKSyNBZRJX13U
J5Qq7C1kEXJxWPpq60UzkWNJTM2T8kAYOpgKXcjBOeE=
`protect END_PROTECTED
