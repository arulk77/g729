`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGDkwMKqnMENzklOH5ThcXP3PfyWcO0dweS5FFOs6pne
2AVpPH6clfi5FiZpb6hgQa+47cJWbkPBzbFvLUyNnNcE123YNmr1Ix1JqIiEz10/
PGmmaPh7jGefUywIbH/HWoD87WKAYrsvEEja5nIllRGFucwrrIvdS0hRTyiXEypi
`protect END_PROTECTED
