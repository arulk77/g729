`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNVimMhGVs8Xo/PEP0y0/Ssi4iMUeKX6X6Be32pudW4Q
nI7ZmaG4lvJbO3pHHYItfIU2cD+OaaIksmurnBNM6pZeY+w1NtG6DeZs971H8p+r
UhVUgLpkXp4oTEiYiu6yYxMi5lrgqQNac+dX8RCcKMTIVCMWzWX2n8HuqJDYioQ5
6AgILJAcgcZCvW2ox7w+oI0au1vyOPMB0LFHdXF0kilwEVpBHML0fRrE3nyW9icn
JBpVUOeqcgqFQE8ctSeL6vhZ0ywv/AmVolptu5hyxKxN/7nuykBCIomLZ6yackN+
Lb5R1e6mg8XXnUsu5bsCIQ==
`protect END_PROTECTED
