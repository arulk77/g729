`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ZJrAgmIf8pEsrnj6Mo81snLY3dHMTpqJNzUpSQGf7MKjTQSR6QHmEevMUDUPYrwb
VgEQVaPXxwJF5DATtda21izlIm3YeVqUTnDo7t2peT11nkwy4KawKJuMj2mqXeKJ
1YKMyCKUEPNkK97ZXvL+9pHP2jjlxwo8sRkXR49RMBGmW2ERd7tqAXbQxUDyoyN2
rl3NO437j28T2ost3hK+Qga84tKWCvupfIRh1yCViYM=
`protect END_PROTECTED
