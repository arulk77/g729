`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
lglnH8bxKwjDRyynkS+1nDfnzvXbK6K1QvUETpCS1lEaLTcMVhbnmR9LqE/BmeYM
jYvXDRhKg5C5xV79USNk5sd7O8XVTF5CE5aBEP0+MjScFQHbK2PPNnA3C96yY6Ck
dmMYupfhnMrDu/GQW9GW0yiDy65oeA10DMceSUyGOi9KeXjQ7F1+p+UtjyfkzzqC
y+aYIuFWIaPeMcN/AnPIMKsPfhkHaqUOK+1sOuXd1i62Pu4iXqHEPo0D+7IH/v6v
8zTW8A/PqIuYwnwDb+m814G9nf0yeHsV8uVpy5y68vWfM+Kb6IppUplFhuef0K7D
dsyMbeMOnHbJL2N0mDjb2x2sJ0ZtFcLCtLPxrII+bumJWKUsCnok6GJuuitsqjbQ
SdX+RH4iszcc3r1/AVjo7O3gbXjyRlzO9q71fuFM/5NPwe00oblfHO81bsLXH6nN
XrdFBa5Dv+8kScMTBH9200IjR+n3y6fUNipN1kwrQZmPyutRw4QFiTSeTyTo+VWA
bjSVWvx8cQaG4HjL/Cd/q0jDBb0KBWSs0GEBCxgHk7OqJHSydKZVkoZWVjawKSGS
ezkn4DPiNQ5jgZQT2c8qLX6ZevnEY2SyqGs4m/0nwv4qEcLR/RiN8pJPQT7dijzO
GW3dColYKB0vPAcCKI366mDfedaGuUCGdlf44Y292S9jHfBAl6HuKZU7K+r9c7fw
NzhFkeCrD6Dm72Alf6FUE+259q2oPkdk46gZTeXuIGx4gB4zlyZ3tM1QGkl6UKsE
joN47yPtj0snxKGxDAyHPFXMUWUlyuuyUuP+U+G/lWFTHMKUITp9D49c/Is+mPN1
DcA31KX8EFyBzuybNYow6kdsADm8MLQRlfKaU7f1hUyEjHTVVV6loSxX8KWezTyq
OWVOCar9J+WJPRC5bk6RinLT2ulM6YoHbN8LnTM/EtlHLmNJyjMOQw/kLH/JjPY/
v0yN5pryXvBJOLeMkPo+jmKHO9/IMuFrvm7HDj+NmLYxCdaWm83i8DRCe5uo98EX
NGtS9t2xLqByXkzDsqux5Ox/pSwT4qpybRwOjRkpp2AytirCEY62kKOLjeYKrZ5L
lZi2viK0xuStiKyESVxP7lZte7GpJhCskiQ2ZXOycRMvbzSCZ7OkUpEf+JCxo0gt
c4hQ037sRTk2gLvtXDWelCOa6Vp/eQ582TJbpSuhApp/B9il5DQZJAxhC+bqbqoz
aiSGW2SaGcM8XjBa2T/pi3Rb9jOFHxht+YYcqUys5iSJlB40kgdX8qwBi37njQ8E
gNR0eje0VkTE004+/xGitRlocQ7Bmm9QAhxXIJ6e+9eVo2ejRPuMZ39ityqMfZk6
3yZUEMyZdLBx8ZjJo8IvbzntPh/BDEnB6wsTzTl1xbsJURT+zqVtbQC/gsNHT3TG
SSBT40Kjo3D6CMuYISUYT1IuiC2amfR+G/98FE35kXWffwSCB3qZxDF+GBwTQjKv
89PNZ/8mYN9ZhtislEzInMLpxPpU45Kvmb/fAfO97AHDuujyrr+2sakaAzi3naCH
x61FpIatvEWCqs+6yTCJ6NuRSEEvCkokgSqz2ozrp1evsaNW8WTKO+paLNzYcLJI
ts2MPacq7ya37XE+NjNcq2+LuRpvV5jPPevNa5ymBEWiKKr6ei9tXIzTyAXE66Ss
PP2oNhCkroTiZFhBNe6Xfb104sbnAJ89CN9y4MvvAmttGZ+SWFDDpLvelCV2kwzT
sMv2UvMgBxxSFqGh2f07Nu+Ko6E7tsIqD1jCD1Wka89FqK8JTWkJYitnIftIxj1Q
X75IFRqHLp7P4rtMbEoslZ2T8x0Uvxfw2eHMNDQbt/Gdp2gj8G4GQgQwGiuwUOFT
8MFoP3Jem77uihotCVdRwWDMOd6qMbrnkW/3j62ibgq+4+91hv1NoJQA0Y2pcDYE
Cq751mCtr8kROFJ2TaRxEHiVQckt2UFp4v48e2lHBQnvr1ZXIMR/p6u7EkWuo0iC
cO26EYwokjS2XSy1PZ6LiW7QIZBHPETNFlJL9p+Vdmlu7roavzAVssBv5Ln72eOD
2Pjua9hxYgyYFG+Kq3njSaMGygd3oMvKKuDhaNEtNNdvySf/3tl4alPD4PBtgvbH
Sy8JTbPPNsQrhUebh2KJfBurOL2BmK8w2mq7x+7aEPZUnWTn11Cs0XO4AyuF4mpx
5WDYnhoU0htgN+MpylGMq6Rrm6d3ur3vMEmrksDuE4j9hJakwc9RNv+DOKlpwcDU
6qs5Wwk90T1GJCac5zXtIhojWsOk5Fj43hVbWpVa7YNEbeWvnFUwVf5Y/KPIJVax
ILO3yIwQPIr8PfPOMZmksZddonwAG2V0r+2COGGFYFYm2kozzN+vjnklOEYXusZ6
+yULC+mpF0k+ycUlAXH0V9CUht18Cpo0H2wqxzxJm6NyCh5rOKzLc7+wBpSck/tG
1nl6S+g1A5hMh1q6ZGwDBtXExpi4j8/bknS/sHaoYOnals3El+PztMTTpZpMycu4
grt21Eg8YWLMXUDfDxvaTUau5uzbn16m6Cmb+tW+OEha2+7PcbrOT3AKVrGdHyjn
n990TGVA4nfRcc/nGu4f9JLV2dci1FpTZNlg+9Q425u7y4nVFe9NzrmXg691JfIQ
XpazcWRcLBRzP9opdcojVblOMmRqyrhCgs+PzaApSonU2SAPl5OCzvqsuCUjDSXG
FI0KZiJ7ajKUP0tSs8bn/QdwzMNhU+XdVWdcuWT3+YuOJNloZkfVncp/hNIdP89q
rOF7nJCLEG8x8hHMyuHw36pWnKXeN7wfFMDL1wtU0zZnGjtTKTEGBqqmDZMvd+7h
ate6DlVvV7MVo/yLwUKK9Fa6E48dt/3Pv6xVbuVkDxdde4Pxob6SRWsu9N2Z3Vfk
db0Nk440rGrA3KhzaHdffJFMmmEfSKjgQHpBudqhwLYLrRWaXzeJiX6Uw3PlDFHn
O0dHztlUU1EUr73hAendxXvMQyOWnKyKdXcLyf4FW8le7IfH5KddH5bUQxC1iKVz
Xx6xwGV0C3luP0Zze0hFA6+a96N/BFv818gM22h3fLZ0vs5J0iD0WkEOPHO50fFn
dEftE+UBFbMptcZytWgd36ws4vlljMSRrH/docfuPMpfrtxVWV8g7wUAUMIKUG4P
o0HCi6wWqO+CL/jWdst7MN2Llt4mWHY7FqnJaKBoMv3zIwVd18N0PF3WMe3qqJnq
MEH1VHO2cSZGjnrjm4WxnqaXGNIUxjjDLZ2WSUOkfi1u0AOb4OAI/l5xLp7YyFJg
E9WKj7dNLwjH5aWEJ5XJcQ==
`protect END_PROTECTED
