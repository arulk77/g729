`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNGrMeVAjTdl9O4yoYLayK5plMXLuuUA+bqTXowq/vlL
xh0BgiyZLZddujtdPkxxFOCMM5kU5KVlN6nhDFijZAIWn+QnP0WQOXk7aD3INHnx
B4usvRxl08IjoMNRbmBuHrZ2lC6qhhNAG1bW8nWPx7rUoYWQ2YGml7uFUvkJSvX2
bbrcpqQqcg16YUP61UzKF261Z0sCZPh9R6hgUjQIIcrLybfCHqEV0YAd1Cp7Yq87
`protect END_PROTECTED
