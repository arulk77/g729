`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
AavLnXHMT14NDOFWHX2P6YUWbGkfe+jqotagU/wfi6rbN46u2nxUlWrWzoI0qAE4
i9ztP53I9bfpOBAvxjUG9ZzTsJ79Lr1C8Kw2ccDpD8vV49Vo2cgGYIcRM9/W3JN3
rvNmdQBjClEC60+4Q/JuMnxv4ZxfRDABVYwJ8vucLpiN4/UbpJzUIHNWY5QtU+qA
DFgEJnno9M7qGECI+TN0Gui1WF85CH5BzvucYer7Pn1Bx8eGvrGydLn2BbytOQQV
d/vkCT0LdSKdDr6r6v4UkJRnASBp4O8Y+0WY6asTOiKhc5wEO7QnGp6uJ/YmeeoQ
ReSYlxM1FLyz56vis2Qv0RLY+M8WoAtvD68XvRtf1jWnxrADOFiDS7rufrHpiltr
`protect END_PROTECTED
