`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL14r56u4bOeWqGup8g1Xj+7vqJE4v/g0Jgd7PigNaqO
72nvOEXfyWrkQwcAV1WuvW4gZofXz7N6WkGjV359ogr2VXoYSkMHcAWDhgFOvhwy
QRX+1Nas/JDDZlsu8vATkIW11MijFTjw3oghdEECRdrs5+HRafnP3xVyR/+CLs7e
L/uEaTi8ZkC/ts1SHbx3ficx7Qx/VHt9zn9j9Lu0L/CmO2BpOwlxz2qwB9NEW2hf
aLOujrWn3RLBBFCFNTEFGnXEK/rP+UjVn9id2XX6FVHYf9GKJiLfW8pMPNY27A2/
t4HATMwRopJN7wSjvQ/gV1A6TulM4eR4btXe052oETGHtyuadABNO9w/1fWlLJd2
oyFmrzHoc1IsewBa86hhA+H1P1B4lSFBMQ0n+FssmXeADEkGNuJ1Ov5LP2Cd+y8J
rP+c7yJS+2GRe79/EfPLOylDn3cK9eHvtTOhMNTA+aQR+e/5Cvikpmv0cCe8SHoZ
fCq8cevc4r7BVD9dFOwV9n8Sye5trtvLZ5vNrLNPrIRWYp91OeO1ZyR+FlS1dbRV
`protect END_PROTECTED
