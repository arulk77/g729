`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41aqPCWhi4XUkvMVlagxAhbsIG/AeN8ZTp3KTMIGvlH8
lb3ApA/70RHfhxPuZ5TnwkzmbobO4xheflRyxN0Gt2YGilmA/HbuCz0LmBph3emA
c64kQE7/qXCMNt1rRgmw8uRDGqqxXLl/J16uCwdcIzwbB8L2PTYQgGbpW78S1QXL
dvN0hkPcT/d86EKEqLKtj+/kTrqSp9mTlLxkngdipw8=
`protect END_PROTECTED
