`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SV9YcCR29aJPhLc1Ef2T3h4OMZMVjeN6gLu5OzjulAKj
+McntNsgqaW6B7konGJfH4ADgICbHYsL2bzUfGQoZFKLROGLNs/OvbQKcQiZ7K8E
ROGKGk5jJuGpml/qKHsG6Yl2n2Rp9sQs1ajKZ3goatXuy5+26dnPoyUOH27xNOpE
LbwFv6ZmKzIeHY0dIz0p/5wmQLjPRoHhMMRNzh5+1Af4UrJKD5/IOFF9GEwP87MO
tG1Bzcn/s+ckInhd+hrbGPSIcQmIkEDsDYCoVsb+p8Y5t0UhkCELv/x///FGCRAc
g+R7B8ahHr70+G38+15IuNkYBr99SJvWvygo3l+ERqw6NWRUhoH6vqXXeOFBidyG
g6VJyNmr94rUVko0D5Xw3JDA0q1Bdq1SgLqeu+qpMLb/ngZ3w9XgUcbeLqLPjWxj
PmkxbDM42ndhJar/SdnXN4F/pEeY9YGyN5X86fT2Paa8WV1ngR3zi9mpyC19qi7W
Jl6Y+KfmQ/qyAexNzO5DhWOXBvlQykOEXMf/Q+7a33C5KyQbT2zNKWZ+8mkEY2kx
y6/I3VLStZdwcdVp8ZeySGdqwbxY7pjgPHAArKxntTPkpvrNV+tK/kTJSl2YNWCa
xnWJNo5om+6+6dliFCdsZH1A98p7r8nzffTVavWrN4FbrzffkYoXgydNjjSIr9l8
kx/non3O6PJKBhT6UMDW2ASrb6nkjSUvA5QcwMGFCvfHjytaY6J9hFk65hVOfYTi
465hVWk8hcuYyz4W7mfQX1SUeuWSat7u+G7kfiVY0jglxlwojTqJdQ5vKF+XSr8L
Hg3k9FY2M7IfAvECSTrqD076TqM5WX5jyankqxpyYgBQ3+fwVI7JHOluoV5D8D9I
Cwkc42UV60pFet02tSfjNXpDtiQPBVgkVlork0mC41I1u/3w20GveKS3W1RsCZmF
tgC/u2h75IcvjkPldGDujskWa5YshgVlmWtFypZM9jjpBXHC/cQIL4Qtxb+Xw2zs
yFlZQ8zwol2BujANAT++8uBv9XfUXwAgGMKrjTMaqFGOiYJztcqVfIrBXPHlK/hm
/tLkTE79TQChcVzto/46v0tmjn6z8kuHRiC3fQVO1zxK4UaTL2kmI22j6PcL+6XU
FHIALtT2yO7BlEbi9oZuNXyI4bDghSTq91ah/nc8Xnjep1CscLBI+ZJwD3jsbnF6
qZnY/XXIgchq9SG0cGXvxojeMm5EnaTlZlHF+C5ZnN1R7E1R0RauVqxxVWYn7/3I
qn3lOxpxYqFQui460HWMWmS5qmNL5l6uT88uKN0UD1+Ax3rBesxT5O3T2fJKYSal
9K3gjjJGN/xPdh2Wj9MojNKIhKy///VFLyIEUxrOHmGOJ8u5zgh2cO9qd0/46LEx
lzQqxOmeaJs/aYeNvCpm5vjlJc0RAptdwNVFkop8A2XbK8Jl3yxvRo8N7sXbAi96
W7T9rwTXgqQjk8pkvtGrtWS3dmRB8Dr/H0Voh9udLRJwOUKh9dUIMwQTd1IIjGfH
qkw4nzWqr6ap5jBu2PYikPceGGaq+cSFwI3SJ5AOy08Bgy+eQDVqXHlN2u6gU7d7
yW5GUOtxSNb7FH4u3nT5DOOQEzLdBwIGKZjtaEf/61swDkdBtPjGona9G9akQKCB
1Ti6cMOWHU/0pfEbxn/l7u3uBcwH4FWWVn/8aTx2J0EAIlvpP0oqZ8ClfmezeqH0
/Z9HqII+YRhlwYwvw4nneGPP+f95P274/Q4GT0nfGMx7YHbYLfFw4plZEFxqxmpl
pwSAOVuae4BSgsxwIhSm8ucHl1yQ6COP1dGTnYB/+26ebt1NZmtZe68nS4ckSGAj
kZyhn0TxEVJ0af4VgMdJK3wsfe7hjsW3dRhcHJUh9KCbCD4YjehGbltuA3csAoB0
IAEaa8hiQR5Y4fCvQQX20QxaclKru1jOe0nq9P8i27jR9WBjt54FDE941uGSnpPq
vDM9jxocGCNalueMxSZUtw42/mHn4/rDhKoHKJ5UMiX/kCWnU/FqYdr8sLLZK3uf
BNfL5C34p5NXlKpqduX3YPxmnsLiQgOlLnz+6nt3acOsa/EBEnY+vyDz2m0O6tzo
qqH+GNNPiKXfilK1H1EoFmpMaCwvr5siJUPwQr7JEI4bYNPySdljagGdOlGtugNM
FBK/6BCSAtVTfVXdrfSXelcVdmpbck8IIBt5kYAVc+EWnPaKGDIFzJo9hcrS2xWP
oGHgZCsWg4DedOqhlUzSCO5wPiIZDB9lnB2+el8ZyiITLN8x1MQBc/Zdvk3RKGey
6oofFf0HpLaFvGRGwt3l6elRwS2T69SBCrqs/5UPHaUGh3+PGVJmfxDyU3llpob6
0W708EWFkF7+5x3oiRTAo52tYKGG5HzMsjfxAsHDPVE8zmmomzaLUxyqaWVnQLPf
91oik/AojJS0AQg80AieywefY3Q4s9b59cdtKn6fsdWP8jIurM0RM3ZJETIyCA8p
eLSCtnMWD9K8EVFflH/0NBlHKXtUE7CI13tgsaMr3LeYk3cO7mv11hob4uIKmzvo
rixtt48KkJloWvKWhBemUXXxnU4qXEDzOsc1B78jEatdst2xVRrIavR0HKTtf/rE
2dPXe8DrlL8LgWC5NLb/ExIUAPTMQ/WBjzm5ezlaYflKvHKbxXTGlg+tUSnS1Sj5
8Og2Xj16VTh5C640CEJEipOLZLyQS1wFXsZ4VdXVkPguJzlA6BMbiblF1+ZG9d+9
BfCN7f4Nzb4mLJ9Rsxo2pTvwJJyvJK1QrZiVR8JoeuMvhRi5KoQc2vxxMuOaPyqY
hwrDU+PLZetCzrGai/Y9fadQdejaAcKn/emcRgvS0yPG5/jj+EOPEeGitRYEwr9E
7e81zCPPpBXl6DHK+bdZ0vyYbWJEqB7es4Fmw0y6J9rircIpmdDXUuEjm4bNISi2
klHqj39hAxOfXKuhvewNzMLf37kU71hOaFTQ7Tr7VCoH5G8NRp+fDUAHCkp1dwMi
QtH30SFe+IkFZxdamb7LXop3L22Dfv+6FvRkCIERGQlsqaUbFfmTj6vLe/a00n6d
a6x+z+Tcn/maN+3lvJr4iHJ4Y1yzbLmuaE+1mKpjN4s8CGmxfNIKI/b1vSHmPbY3
Ko+F+QaAcbkq08xXw2UGqxiauaddzoKU0ec6ZJlFZdqRU/Zs84BGAPT2wuAOTXJZ
3MGqKGdcfIU7JgBc9uyglbQTuU1ClHTEVC0kQ10Wxo+/jn3kGz4rrO1UrT3ar0hn
t8hkbk5R9GmmNYGRI3MSuBzOIWg8wsWsJCkTh+ODD6yZu/udEdRh3oF5v541P4Vx
NrrBORNyi/KBwQhOpF5L9A==
`protect END_PROTECTED
