`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL6Y5V9q0nkQ5uvok46O6hHGP3nRv0y4Nnr82qzkapML
nr/9zbs3Lm+7efWjNR/oIaD03+jqc1Ori19z13pUybqaHP2FxFYS+rxPgUJXNsBw
nK8mzTo/xd2LMyc0z3U/bTpUEBoAhusXMgm4nHfYR6SJtGQFRRB6zEV/07Hdf9RJ
h/ijgLcpCEtwjG8jrMifhIND/2qTRlz1SGMiwZl7SmkT4mdZj/8LRgf2J+0DhTM1
0TFHwd/wFjHPHN6OiA8Dtv3CGIJplnkYiRcJiCGCRNNDpVyczFdUepMi4feFnnfe
iK5vlEpvtVwEYab+iBq0dg==
`protect END_PROTECTED
