`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePpPnmbeZR45jtMygMLMkElNs2dB/3Tk5yhZE4JJycC8
Ja+r6okH/GHtVQR+eQrIsBxXCu27cgybqUBCAsSpS6cwRUJYdfMZenAv8tmAsTyO
XzgWq2dT2F/vwRE1kZnZqxg9EjFylIYCkBn83ddzNq6D3jSdgPAO72BIydqYuz1E
wM216itwgC2stjHuAwTn+w==
`protect END_PROTECTED
