`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJfYd1CtB0Eg6nb8zfLbRTu4ZiSaMEg04wvzK2/hDA9B
75kgxQBPK/uiHcsHtQAO7lcz5Hxnv7nUgar1oCpsKR6BcIpb302uwfwbIVZEhZtd
6sFUgo0JB/Bp+XEM/4oq1usQnRMhh0SxsSxH0KxS7/C4Hvl0p3eDpHDcFfjXe6x4
1T5m0uzQFcYqZ3M4Zhalxg==
`protect END_PROTECTED
