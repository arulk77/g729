`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDXMQmeImi2ngTMxlm/c7UfTnil6mtv73nSU+YE7PO5C
cpkF8GBxVoMH+CAXfxzWbUUsW6aK69UK6oUPM/66XDBl4M17gxERaylD0xU24N3q
uQQ0wQ6BZO5CfyrcZK7PWx55ZgVcAuWn/rB2979h+8V1atP8/dGXfFGtSwVGuoaS
`protect END_PROTECTED
