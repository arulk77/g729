`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
W5cN+hr3WbdhSoDpFfx4IZV2pc7g6DFKfta+czu6hYKkjtaTMFZDKCLLayiNzu0m
QRkDSqUOSWxUfEARObVVu8AVz8vblmgWkyxx3UjiJch/Lq2EXqJOmbAXnLfijyuS
Q1zCCQALWyiPJE2lhZlv+GoSB0uxP3DgtsUVtJ4K7bmWK0WoBestRcVC+HKvZ73/
gvX0Cz+o/8Pb9PcXoKwxN1D0mbsj2zpmH60Q2/mVGv5g/u4Cyb1ltN9YZ45ToVV0
oYOfcLSajRyWx5rp5SiCb79aRIh9ZwXL2apDwAnBu0IZRBUEBZkmDWy5YRBshQPc
ZQNBuwMsqNx/pCySgWyHSi70ny/850t2ywdHP52gLWw=
`protect END_PROTECTED
