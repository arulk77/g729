`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8Sb1kxXOfDNlCDnowHOc0KO+GKpCFwQBupG2hWOwcvgqE
QUntU5RAbfAC9Zp66sU6Hs4mPb6yBMMpkFICpjrxEZ5DgvuIH1FWx3VlPKpFBbMS
SM8bE9nkk7gvUlzXyFDku81dnopZkRcYlVogc7rgmo04MexDWc++JutTQ26w2usI
nD9+e9CaDVdHanHTKC2H/qNPQzFJ5R8htfJLbUrtOl91ftNPhG+1iMVNMGqS9t/C
uNlyale8pBbeC2v05NjAGbJ5uT7pAkbcFEaS9cWZvtWF/iyDXTNzZUw81PujY1qQ
8V7Xkx7FwJPbeI0ezKcWnBtM6JCvI9qVthJX5Muk7lHbZHpCEN2qRdYeF9umXAjy
syDk1yGrWQNXTyw1naj2/9NoBFpWv9lPot+gN+MaAAZLZ35YA8po4h0EHPL7Rj0/
AAxGxC8YacqaHZV5hF4APjS3q975DXd8H3WvheN1Qu4CLRdAjDnRABOWICsA/Cxs
Q9O0zQfx/l5+7PWQoog80TNmWwqT8Uks0T7kk9XRnNhpAC5w5CeSDfpgMDeMgU7A
DVLQEKUaT1pttpcqdKOfagnEAuWvNiVnEiwd4sOWjBU=
`protect END_PROTECTED
