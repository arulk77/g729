`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOvMDxs4k27Ct+Jm7szNy/8YwFVtOhmZM4W4evdpz/lS
msf/xOya5KGD8U06Aaez+/zlabAwUlbeT+8lCfGkL6iVG6tx/YvTOpjopZfklRtG
cOK0jt94GlAn/QeYW6iLzGqCkI7aKTeHIs9QBvCJVDrRpQrE/hBsVDWuPq5wVzH8
PG0wSBA7DyUFVIuGiAyDsjR3Up9QieCygsuJEI0zQyEsXlDYBXjcYTOPwHTML0gH
DwB8biQUIHH952OfVYeq0k6bh7SaXYkVJUQX3hDx0Hh7NqEXUWa26vzdlxl4vTvZ
BKqPKn4PuDhoyrtqxacrARlltPBMVMO9RihXkvcM8AnmCGvrB/rlFUjyKFzx7T+l
UsSez2YohWDa5xoyqmaEkhOKkoCQCXMfZdU4b0o+VQV0RwUKbJvEshJHq/Khv+aX
KSSWhGrV7QZZKpX4uPV7an+8WOCdOmJbmYM+gZcGXsuQ4iUFbouXMNxjJd8J9ty4
rtPCR/vDJ8uxP+fqb5qHrdNkWKMgbKnp60X84KS48AaxY9u2Ce+v4Z9Ru9CVHvKC
n6mWO2rrUbweY1SGJHdr8OOqLXJy7tD8N0f8+q6KQ7j/dE5GEmctn94lmoCqdsU+
uUmaaI4q2bVM3YtDwV6JFS7Cq0sPVjsicnqhwzjKJPPvHxYOl8JEBWFIed0r1MtL
37aaPgcvpURRWQhysm/X8m5OxsGd92oE7WtSjObOlszHMPr+WmoL0IueYTANDRK3
6jrrKTRihWo7bEgEULUUQzLeERY3G0OE9zYKaK39q4g=
`protect END_PROTECTED
