`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHtAkYwz+XOkpaS4VLO9yrBt7QLnlsFPqvK+AStJhy3+
awQ9tUt9nQ6vWKYgdWWiCXdFBctFTK5y5Lwx+M0qGWqOgupN9Tby2p/9gxqHKBYi
w6wx3FUvcTR+T+S2EYaIuqVFhqLIm7E+58jkNHK+Zsx6Sw/I7U+tSvMd3y/rsb1A
sPmjqBGARtwT3aa4hJ/27NeXnDSKEv45e3nnrT6tKrwZOdQALjRGjql0za42uT4T
fBU+47FTugERf4kVqORv1OkXCycJEqn1jSzdpuKxSCiY7D/MiTDAVIqoS7vy9tFG
q/cbE7v6cWPzNoRHrEiZzXr99qUsUtovkypvNRUl6MTK5adgWfmJFQ2R5nOUWsI5
njqpKe3LfQu4cQU1+Kwq9hxS1VYL544ueU2Z8qV50Pm0QR41q/GWwYgMfdj/VuVp
HdkTAnBJ1uKNF3K+5ErfIls/pHQSjFhJH0pT9rLxOq1V9SrYJNIOCQNFbmE6JExC
dCnyNSUXH713497gH+6yjEYfdw2T+Am2IxNP68tTScEJujcyO9smgILX4lVSqXBg
iExtlomiUg5EG8I/K4Iee5EettVir583g35qwbyNsPVvDiMCR0gNTpxsohjUg0Dy
BlROI1sA3ZZVa19HLlJTp9EO+eeD33KbMhqDuaNJSr1IyKb16zLpIZ7hAZg+0Q5M
LM1C0OHX9a52T/Po4yd92ndMKtoBUmxIjV3EBI2psqp706rZUqO554AWk5QwWTzc
VFw3P5z5gBFZOBvQgrYpTrCGwnG/ScnTnqq8Lz78sQdfcENenJJaWrJPiIS6G/Hd
je9/UingKb1kuSi/HfTOy8ZH8ZNl4IpWHqRLIAdIfzvlsOKLbaJU3X8VVzL5tS5i
Bz0EoXDwdm3jysqx7Wd08Wkn3t4lK6bC2xjs9WDLN4rfk1Bp7ZVL7Wfa3YuLY5Zz
880ISl4TeOW1L8loKoqu9fyG9Es6qbkq11AHiBc6fNk=
`protect END_PROTECTED
