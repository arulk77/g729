`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDCDk4k8UcyT14u2/hu0BriMdvKAiWWVzgDsT2EvurFh
S8wDwdDZtPsOnP53sWDsV26pWEr2dHjuwQvGPqqJb4P47KPJp+QjQxOITgqGqlCt
jkSUj6adpoiZ7GA17PMqok48KM4nKNLuCe8CduRKaDcy6jWZSIVYS6q2Gp9Qdy3b
66/NIpbu06kEp2J1TBCnINIuhgKhInm5LhNmydbfVOvHobIaw9pKjbTIOKFm9DPq
9xcCVakb4AMEs5fbGic6u1UtzQTNh5CC5QKIbXaH+dWMckXOsCi4mBymsTotWt9J
huJ7nG91iclZgfCn9aug838WPG0mAlEnJOit78sVHxDBR6Nqf6mHqFSJDuEwVeA0
nrZfSiO+cg1T9JOqnuXzWnMhQ6jTDg0k1ukCnLFN27V6tp9F1abjyTBw88WDboI3
PzfUmEStlxZ0q1/bjWvYMPNjBUR07hI/Yi85bByAz91RQFDenHwVwiSKEASc9LI4
aIfWQjOI1uYErSsRYvfPPD8CO3Jjd2xsyFQm4skOoBgpnOQx5iRluMWlPBB02/1+
IgRaYFh+ZdGI+uEHBUcNZHlN0WYnGw/rjcf5CNjQHTaPBaZe2EeuX1a2UGpBGR23
IF+ArrvUV3b5+1q1d5WAvdCMlNhnC0RKF3o0wSDqVUmYQnD3FtY386qrvBdHRMCE
`protect END_PROTECTED
