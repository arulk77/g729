`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMZkTS9zK1pin3dGzG5pulYNfImjDp80K8PjCCYUNrI+
2IDYpQn/8dpq3IqXHD8jSZrVxLzksmaMUCgUHLuAYiO1fATjvKxpUsh62ZKf4Lmc
5MXnri6CqiVKVC+XeEEPWD5YAO4Ryn6EoIWHyYp8ivnEBuFiQb/3BmWArYe1UVAy
H48tQaxiv+le4ws7XBLeg289jrEJhKSTZtKUE3Am1fTL3GYx3x1RhZ/0+XtcQtEt
TWUxbB8b/Lk2MFPc9zSG7/RiQ8hCRgBU3SLWcyWB+dRZtGJEUZklXzVcb1O3RpNK
E+C1kvpXsYKM95hFy6CGWw==
`protect END_PROTECTED
