`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
whfZdEhQhIVICrvn0VMg7rbRQFp2eHkIx5TY8eyQdPXNiBDwqBFHpjrPw2HMUnA6
twuIepARZQWghMfW1VPY6zgWBZ81ha61gMLECk5zQJV19G4Vde70cx/lC0OE+aey
idYfs90GHQUCUQZzpu2M6Wq5mO1zniOe1E62oqE4AZJgUjIA0qeBHlDccteHu1cL
ohyWayKqhL5x7CPWa+i3Oo/04JD9rtbCIbKZnrIbQPQhr4YrfvG6YRjaT+QvzFp8
mi13Dc0uQrIVWiPZjw4nXC9LoudsZvZt2ftKd562s5B26PCWGdteh75hjAILG+4E
`protect END_PROTECTED
