`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42SQZ3Q3d1Q4p8R9fT4U84aIXmH36e3oSn5/lX/A0Dsq
m3WxW2vRLg2N8vew230EJPbvEwEF3MRoThMfbq4aiTi9RDzmb496kpqAWqYG/upA
TVWSYU8fQgYcLIx6HepmI8VXy50SFGBbiEQgv5l+EJXPADFHMSi/nxxYlbaRkPet
v1lgv0kWOkjKoiHcKRICunoSW4MMIaATsfeYbxHFbcdOCEhwJ8em9F1YTKin9e2u
Alni2FOs/jNNjwW0ljES12SJLnbxVieZ9mphzadW/cpQYABxfBuW9NeT6GrhAL9a
XjJcDh6PIAVqB6/P9H30/A==
`protect END_PROTECTED
