`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ExDD4P+jZjR7MIIgsZzaq/uHAHIZnKPNmvkBtPjN8KhdYuw3sEcII/kKdZv8ekK3
nGqvNTEWoLuR/rX04eu5Cssw6Y94pxl7FYuEaAdr3cL0kDUo5jbCwtivFGANkj5u
SVT9hPBZoVzjP38c3b8MXbYj4De23knnUHQMAHBQ1lUhtc26IMCJ3oItldpp1kSe
BwW3Hq5L2KUeO/Wdj2knojUCf7SP0pO/cSLIzUC+lDK++QKn0hrK8THH+njj0feJ
p47kKCyE5zRXUUVG+xhOyxoyED27neiNjA00F4UZC0h3qQZ6W/Y3K9J/oeJ8rHDE
hihM8HKimfcJW9rHZt7zNLXN4kyR53DP5Bc+loaer3ymYAlwRZlUZe7n3tJZ4F2x
yqs7OYyQLWqY9FRR20iHbQDGMITn/C1pUR4T6hyAEfvh79CT54mzr4lTmUS57IRM
bYs6uV8ixadmbjhM9YfjSg==
`protect END_PROTECTED
