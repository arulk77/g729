`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveN/8CjQJNViXv6KJmx1k+qwtMyMkQOa7XLp+obMhanpp
aOg6zxZKX+1fLZzSbUhZG04cugar88NgaNsB04HDD4ZJ+cth22ZXhH0QoMJLhz89
1th51IEfXIwOXKU7Tei0C+EISwgh5KyzFPklFsUO+88yUJJktVIwJt25vWIvZ/pN
Bcud0YuX8/ikkRBp6mMFzldeP2UYhLIZrsAvF5Z0H8Dhdburaywz4wSGdf+mEfKA
QTcNIJ+G5MIyRMh/+ISfsTcaIF1n06Q7y+cGBUIRUfubv/JR6I+dj8q9Gk3PFS3H
/RCYdHv7CUQpO8F06TLLoiW9xEpL7jhG0VpixasrlOONyaNFNDa8gm6BRPsmWvvm
5w5PNkdL3NieqvawAd0Gqw90RJAPMiXnqyvy9UpNL1ZyLPh4W92Vjo+PbPa7+FxK
kAK9L/oDFrsJETiG0EpiOkDP5KzdDQboGfd87JCe4bVhLOlHEDc7ll4IW1Vf27EA
q6grUmrWXsAImi7nSj06m6WgA9NpP2+UKwJE1wTP2lVFfjMpidEal3XXOltiCJlm
bQ9VbiOuFh4ym9rQga0wnBTn6KiNcjFRTlP3fvvThdzkvgvyli+E3vz/jJtlnIHu
2spZZyYrlxtfMnmZGBjHVUjXbcC8GdJk9KR4AXHfSNBfhQE+T4UAtUebkloNvgG7
`protect END_PROTECTED
