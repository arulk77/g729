`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aXsKSggsU4l60wVqXf/IQBk4vyNvTXYuRgGsw+EXDJ28
MAQFgu59rpnopSC0l2KTxTkDYqTtEgga5yUQrdRkl9L5pBhL4ao2qXZ4GFHsnEMg
PpOs3981zxpk1IXi1WdE4TUCu5g2nhw+j0jf2aoTvn8diKDTi+9nSh6998BbxTaL
GWfabDAJ6zU75k3dzYxPZY1Ba6nyTg93W+j9W+QjnzKHvu4XbDEumkv4M2LPlM7J
iZ0CgJGpfZRz4t+Mpe8C03g+1hVzVtPh7/E4Zs13qf/o2s9LhB1mP59N3KhTV1Ys
n7f+Q0XFzN03IfLcT3bMQpLqK0dli4qg41MfbDPhoQkg7qcLYcxxb8M7o4LgstZ2
Ho+1e2/Rm1XD1qYinc+r/aB9kL5UWhkJAXn7sfVX5JKt9Qub8u3r/ZQrcFBQco83
WQN1U6js3UTVczM96tAf5dmbWn0XHdONWNXofmEeIwHdjSwp1X+9vRAjJVZYg5ey
H199ClMDJ5/wPEbVAPyh7hbTZ/nU0vUumiITaR/kq+y3BObaAbfAIZslviyJ3SL9
RwegKOKfWpsYcEzCVw7WkTDq6L2NEOr/rlEJX6FHbZ8Jy5b6uToEYfaZbXEYNO6+
s8AHjyZ8bMdWxp9eQe6yL65dRn1rhG+yH5ll6/mQ0hAzaHD+IuYuWDY/wtL8y0qj
VMbCc5ER/fIp+fQzFNyO5HIMPUW9aCH86kC/Z7qf/0YOAWLbLd67k+fCrW1gBvV6
WYh9tweC7i7yk9groA+fgNSmi8PNkCvPw59bpun+4OP2XJXCxmYyJA5L2z/npiP9
aJkCCYZ6OaNgOPB+6Gi1AO5yIb+xeG4o79jq/6ed1Cn6NSUBMimrwElnCj1UNE7I
5/dNMVbbAp4DBPIGP+YxfxsLTH5NAekWrxuAmrwamr2nseCTybSL03oC5YLo4qEr
a10jSI23LCvA8mK11iPmY3a0GlUhyjBlGriaTnS8ljJAz8rrbBODAfcSPtcqzUaU
OOTbNoXHajhrl0uDV8WAERiZ7hApLV6aq6QOjgaISq55J4UkTb3asnBA2tLa5JqL
h/uYc5/WL00EF7NJNrd4UOlT+tsg5jJIbIelXn4+X+6/jZeOx+urRbkusq/xie3z
CBt2w7LffCOgwURsXxQ1K3M6ten4U9wpqGwHi8v+AVTTUcBc0ozVEKA6SFP4vFU5
yfXoop+fCBGLqy88U+VfJm3HKD4+yprVr6qw7k5Osx+xQNliWr+NkSee04TFL5l2
Go5sC9XqIS0KYcE658XZ76DvtzxIp1SMN+83aTjwfVlzRXZcY7SMIDXWrgkeFR9k
R8uSk3aL1s8a6tGH9tkFMS1Hf1dVO8zq3di8paZCozBe4EbDUElYH7fY66ldwBaT
oessvgP9JfuZgPQv6oU5lLBgVDlQwDvDv4Y4mxgXmpNyjgGTW4uDm7sj7tDR3ysI
BOS8n5I1hUbKSi1cV3HDPUzyVnj8d2ul7NzEjc8+ujt6fAeicyOvKOr/bkCjfVdy
akmLYHti26shQ+EojlsFdF4Hr5+1SPbTHERNuCpiovCtIpM0iXBXsQAxVJhVs50m
oFZnzAcKyWnr3yjUPaYGbcAhMFbDjtW0pov++L3mZ7belPOIi5y5wIO39HuHJvjD
1FjxPBDAEHq6F4or6dZJfIGVfQ13HPQgRtPH6fDJXrf9gZOSvRjscfwN0XQAPkm7
kAnzmLi8Qm7XD9sDlrKg8ijpXgzQ9kxNtghtZTEy6GjLYRlB70TpFctvJl3oTRM8
cU3ceoXSJhe5IL8qalq+6yzUeRN28hgh6v+MnQ+fNc2ZvVCFm2qs0UwvkWUdttfo
L/6yWlrBz0H+SHH3f6jC3fQjUNO5NEYr39UHKMHvAfGi4sDoZ1ws9JgQQ3agElLs
llt7Weg5QXOMR4FYnHSii9CVTr2fqo2Uuybbfc8Fg9SAcJ5Z8zW00kjyfm6FHhYP
tmdO2VHZjGDBe9Hxh1KWZL6f4m6K9HrwAvMsFakElS/mx/4CixqRkBs8k1KqhmsF
HqIeGB37XvgIkkqJDmrGJkAgxXfIovArbxBgAi7MYro7L5u2b3tBGtuwi4eWVfXL
3ZZmDniBIjus4lvWiCBmWc3mrvMfvK5EEWuGFfTbic77PWCGaBA9gHg8Yw3m2ueU
Dzf+S2GLeotSbJYrVcCzcPeXJ7S+bEieuKK2ZmvPuTTCRNKptqbRf1/oBrTgNgmo
SPBPQk9XwQZLm29zGw4LYA4MGksXdYbK+eLeY0SQP0c1rRwO48Otbwf82i0qJ1pi
MP1gMG13tnnuCXigD0NiiNg+2KsRn5dy7562Q8OljvvbVpvpZsZLW5md0RWu9/sA
beU8rA26wHxFJRAkZASAk+o3akL9v8ASfywJUGAnbg9ztIZyKYWIv4sn/IrPR773
fsNryRl/cT2xwvGbeRl81zZlxQlOExuLFffrGw7wz94=
`protect END_PROTECTED
