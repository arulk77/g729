`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveONHnpK6OtoR9C2Silqu3hLPcIy/eV0SjqJfFRH+N2wm
gWXsXsFojWf7zfPXxY3rYOyOOaEm9Lub2fubsSk5WzureeFKhoBmmGG4Ybt2fC4L
fp2NMvlWKCBD8nbrtK9d+g0QQ25ZWVi1Qi2NQBRmmQwb9qg/Sk92SAoqQm5we+UI
5BCNpF/Gigq5K87WUUn3LJEz2nfpjs5R3XO8FiMO4ZEmkKxO2SZ2wsqU9Cs1WA0/
00dD6TTWTHCoeWUCLBmioFhNg9bOrQjl8RGQ6HHGB1G1JpY1F7WonUnwZOP+u7mj
+CWIYGu+2ylNJ22vIZoytVKMO44Hw51CltIoraQiS2mArh8dHAgXJl0bn+0EU8gm
`protect END_PROTECTED
