`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFVJHt05v6ggve1/O3AIniqeJqaDrhnIV6LRbRTT+nnd
86roEHVQveyZYpYhaYbRDS5iWv1S6VsAJy/Um1QKq+k59Gzf51W5+1i1enDVZ+BV
3mYvVlrQodtFigQaKjZGnxdWZgSb2IeY3QsYS72coVMdr/Aq5D2qiWDKCoBIB6/V
UvVGWtfRZrH6c1W/VwSOawemO64k0P7jCMnja/gpgxF0WOAaIShDFln1x5lXSBi8
Il4jLgdNw37rTZd4dpowJg0QSpn9YqsB1waedUw7/o3eCTn0MUe3/x4Y9b0wMWpO
Lq3WgTwuhWtQhbrTjpPHUA==
`protect END_PROTECTED
