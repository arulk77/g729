`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C30BCWfEYbl1rTRCOiz+3ATEekQHjv48gHdQ7c7HqWrE
E0lasMAJfw2sJ6e7nuzO/BLF9ZkuPvb7sawl3NB7mAOljRF00QruX1TH7oZ5EEpO
HC+llnRfdkPxcuF04nwvfUwcuXlBmyn1WN7B16eSIxScgnknzXkpYN2pYPPzsS6l
G8IMdt/Urv42DeRFG9/tFRWedTcBR9k1RvjdL9cMhiOz60QJ7CDqTaX4ktvOfKwQ
83jDvF+vQiPhvuAqaDGeyl9vdDS4tmGOFTekTbKYQcXS0GkC/cI2D4ejHQfJG+Y5
VoRhkCLVgGygbsQNmpOlWE4k0R8ohjgPk0MkgxHv30pS+ITfdlHtJBkGtVQ6lDGK
tP19DNCTYhKNuuJPzw1e3BihS5Sncj6DP28JnBLlbEnQzUi/he63QbxnGk9+SQsP
pv7Qf1QefZGXDOMaCiL2xuDNN+B/riY7UpjX3NHBtGwUa4pQyPfs+Y8bU2Z7ev1X
peQ99BkTSFmR4gTNlm9bPGT7Oyp5wsYkjROSGsiEOIfx/Cl0stU19QXYrvAPUj+V
BcQLesyUyKVjF1kcFAK9xhILE4Q0/u4eBG9V1WKV7vsITrZzFOEgSa2kQl/ZvJjo
MJoyHcHFtFwnbu3i2WDoemf4+zaXtD13EASkNGGZRQlS8mwYuWN/aBxqRU+2VKcB
3Gew2sRWJtMTJPnmwQtQobSEJ+rDP6c3RKpSRmYKAcJN3j1C9IeXlotsdqJlf2A4
GfXCOgTqoSvtjIIw6rhKHdlEDqH2OcCxFYxnXasGEuh1pJc5nhmfy1EwdeE3Onxh
5Qr6fxmdQwI8jN63Bk3AGgPTniffTRwx+Rl8vqbEcVDhZ6t9Wl2+u9vr3ZZhJOYz
CFpv+Xcz3oYwASQWvggwU9y9l9q61VPG6L/dkuvG55KoBLMksz1DmykMecAuBj/K
ZcF2Vnu8viElnLH+kyWP1WwfZV/xZibNITAvbaFkI01mzkUSuZxzQZkFUjHUHKr7
EqjupdbnCU0bF0kYn4cLotWycIX3L3EamxHIU5AK+GetwCJw47lL6zak8mraRDNZ
09e4Rue/NlVGbCuCAYdAldVLuvHpu5d4j6dnGP+0jI2lprKNLRUmeWFLeG0ZBEMJ
oOOpCT3qBm6VEHFD49TPUq/SuXEYqqWP0TpT9k3bSA8=
`protect END_PROTECTED
