`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu487+bu+efvMIoJlEBLvj5+CeMju18vyfeynoY1+y4Owi
prTBRxstgNKJ/ujuRvHSWgx+iJDB1ic8QKIfh713280HXEdR/YdHER8fTNRD65Lx
OkoP+vWNiWzSlX1D56LLtHWQ1miU9qmrhTibMcWAmFuIWlCpGrzVSbm5vQiOq/70
wXPEDpB7G0SDLc6t0piTsv3Qoxe/VTiyl3adYUc6/zMrqKKsPUKrsmvZBAfZkLCc
ZNrcugc/DGz9KcgGCrZY4Xo4JbT3PcaeFOUw2opzkQ+N+4u2lJqB/qYtN2OlDxri
XBbnmMlc3TRQkPOGDDTmHafrFyf/00IHe1VDJia9hzR699UH44kkV24lZalai/+5
fgFoJ3E5nkuTdAkPh+UE5Qk50pow6WXE59f9lSXj7YNBDP9zu91od7bf6Ygyx0mm
x6BA+6NmB06cn34rTucoz35txY2gysrWr2uqZmnL+CnQF13tC6KFo99s0rFNVsJP
vTcvsN8StS/PxajY+xi+bjFXZcMZr3j1UIlldZZBWCWVJ68ETYwWWKIlwrLcyjE/
IkNz8ECkatosN/uB2F81VgdpwVvHvXCnNeUuGEGuq6l0pLWzP/D83z+dlKoJJQMr
QguEndTw8PUkKYl/a3560ZZz0a3loqpS0G0kORIiATFgw4tfcdxlSuIZIAGZ470T
R+ZlVD6IMNYDlDGJgyElSrmaSEDF2VrLAhkyGATKipW2X7JQepwqExoGZZWtSIgR
aY/I8v+Z3eMWdisKRQHKkcTpqfoELTzkLhRqIvAdltwLGfLp4WMTWraolpXGfaHq
tHbMvo/arK2lg09+HHoiNL5sh263vixPOe2cezZN/YjEtvJ3k/V2VxY1v4IePlup
kM0iZKQJxT9sMi8v9ukkQVDbCTTegqtgQSw009blQ0LuxlGzfWtK5qYG78254zPl
06SyItc2kBsx/bFKwzEYIEsrq0aEjgKx8R5xDrvPIhq86YxAXXgiai18S3P08W0y
JSRxOegZc3nAU+qBRKSK/tJIcDbaXYv21nwAgzl/il30TPO2rTmW2gOjxjHglgmI
aN/x7n5dDgEsxkseoo7d5yEBwDv+AOJgvrfzyNd8ol3mbU77T+TsiYw60Yh1U9f9
N2rdRISDdj+IfQ5kQODJIUgjdaSySOonQ4cb3MJz2nzGQ/YP+Z4I4jR2FaCoqIu7
Y/eN/k6ZIcf5latvuFMdoJ2oSRgEeCV/Wz22fEmBUuoY6lOBiJOuu/X1ZB3YSewO
YqU9ji3Xd6yg5XPd93qEIhXXE1VQPVHT17u2UZstQG3AG+KlmvZO+Z+3qVas1rLU
`protect END_PROTECTED
