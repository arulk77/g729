`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
GTzN4W7nymyxPr/g4Pco53TN4PhtwIjHgHVGiapZLSzPnh9ZF2+4Dm5+twxewK60
I5pp/oiU9mDRDSQCg1HMbolEZC8g3pY7Y/xymj5EGhTUHd4MhElMaTqQFLV1GG0N
Cv9V4hHz3hY4EtyeieU4nz/yes7YG11LpVZdTW/ZMeDjX6y4LCqAN06IhwaSJS5J
st4in1cn5/dPz1uK/IfPPaHgb51u31KPNgk03QTNPFizTxDLpHgoRixjGJkeMjGx
2PURvc4MV8ddI2bFoTri7WjHp0rfe03hSWcG16XCWZDaN9liTv6E3ESngveouRuk
FRldGTn3jP70RGriPJFuGENRVYabK0Pk21FBVWVaPXQ=
`protect END_PROTECTED
