`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
9sit3b6meUS2b6t05viTZsYpKEWFcFCEQdd2Dn0pUndIcEgzYRFcekD3GC/8p71e
9iBlqVBysdEjiFqe7LhRTm2okKqkJulqnihOBSOMrqpVQLEeFu7JAyemQvryAlGM
yXnBBet4hNnk0ZCqM1KyqTZ7ANfZ29d0GwY7et9frDKDQZ6QSP57mjfGjIAhxtKf
Mw9uN65BWGP366XgWc8Word/6htMtwEDcwFA2RXO/9BeOY7F5oXMpphWeP8RvUrd
jOOkZXzyp89gGdQIak8Nkl70DwpsSTd4X8+9BtKTTT/IUO90S53MyvQoYQmlqv5u
zm01nm7OLmuXIKzPg7Wd6P3azIO6IwpBBv0UeYwZxPPJeP7r2p6U/y/P4Zy56vUX
a563brRRXbvopnn3Y72G+4wl378F5X2ov9cUiqp7OzGQmCudP6WMtTyut90AViqN
OGOOVdj+H7chY8FNpPAXIlhQ2+Qh+jQGee7nd6nnn2e2U5WQyXBrAucfyMvukBWk
Gr7+jikiuft2tdcGlvSiJ/EJwB1ttBj9xBc5zKQmIURihi6Dcfsqbecb7/miFRPs
YsfYV6hsbGgHHpWBnGFrhEvLWoH04eG4vNuNwLGmpZAm5HdVgxXHaYKB8LIjcda5
QpaDykSG/cQhJGBsHfj5u4hKEKpgODthsKnI/RxRs9m/hujsuazAwVjKJ4tXFBsW
9RViO1dAaJm2Fbp70K+H8KHEyAwY2VIe2+0BQrW/dxY3XT39cvD0+uxOrp69txvi
wR3u0G9/mWTo30nrNPxoboenc7dnZGvfs2FzJRb67FR0g9WN1kSbjT6wVQQm/Xlt
v0ETj1YrR+UtQxfikdbUIcVuEdT3fPZ8ZiB+WAqJKwMd7D0yph1FwkyHYIODTeJf
J0e7VTBXtIFLxoI/uDy4wajgXkENztSzHslx1bdvKb03/Ml045edL+EWeyDMNy5f
BK1CovIshwH6ImYK+X3dko3LPBIQqDstEywNQNu8CE7YMdZOLNtbz+xjB0sETqsI
B4tBzn3GuDmVcR+wGvQeZk9Q9kPtzhqEzFW4LcwBKXhksy/VCwS8ThQguvtiZDbH
VzYbvYPGjMwl2EzngzeJNPmInJ/vkVXqu33DhGX9YReywhF5Eznc9HkdIKcGBDpZ
FEN6KiXYXFsjNMgHiqg9qs+djOmppCqc/vjH3z2bxjKrZcOrSyc1ahwAL+9Eu8Ut
D45AEcqYqLhc6NRzwahc1muoPQ9dO/hw5DX2g+ycp1XUNdhXxjN+ySREik1mJq5L
8CLOD7euaVoLtaViHbo9Twb5uQmeUKvGVGjCvwJZgczIz+7EmLkWXIe7KfJ66+so
FYgO+fzN2FD4/80h3bYYrqcPBEMFUcMhXmQVov7C1RCskgxdguGC6dy6ywlHR4Hy
MfEfhyJAisx9lT/5OZoTr+AzHvZfLdM2S2/PQmYedSnF9Cc38DUpsXhKGsR0V0yN
SK9cxDrREOa2cerpQwLZsAWV/415KWAzPOiG+YmpMVbiUQ4MPfK3HCfAvVyh3y9y
ss6m86OZG9Ydwtgl0va54h0Xfvq1wuQrQv3AgF55PMXtbcuAkDkICvD33CBrubel
v9Ows6Fe+uthmxyVnVfCMuy0E4pXNB+ogiFm+50XGsrWLlQbpU2aZQI/bGHBMiIo
yCG5+0JgNFtcOBbBtuTGQOllM1eaSTZkMav8ZUWdraWcLcfW7m44txgq7Eoztgs2
JGQT+O8wtbbBUiYJqjjnI1MM6B4gWJl06ojXeNHNSmkqly6plqLUQakRZo4Dmi5x
urB8RRRFriS0DwdfUhg/j4xMv0jdhd/NKflflIpfav/CV0yCazx0/kbrCG6jbrJ1
/RTywb4rEIdY3H7eBoQP/JU3XA2AzH+9rYsOGojVI/X8VZEIopXCWP5JriVR1gTV
L1+4Wb4Nm3MKHH0kNMDDLr7fFunfpmUVvyvHm4PWb/E9d1fLrXql+s4wPGwHSuq2
uRi3jE+XAWvtsR1tpc2Fy6ZFoCruY46NZQ2jenWSu0qbfAoel7SqViZAwLSseg4E
kVdyG2lTJg+H3+TkPFk0ClKIRDvKA3ZU1AAcQZOouWMpHYrqUhFPAD5tw7iuTZ9o
KzTcTW7CYSCMvsEkpjKOELqMwCKUhzQoEGVMNG7YEs1w48JY36vM4hpEhlLLL/6N
RHBjv84A1ZHk6MlzxUDlsvAboK4m73WKatjwSsfrr7rJurWcv5WNmdnGnoo6JjVQ
DPGCN9QCLSgfoyXi2RHy2W/dAjDIfdp5IVq75THDHY6ch5RaQY40MONZQFG0B/sh
ZHhYp0rpfn8Xn1hAUftyNT4Nb2u2Yg7tB5MwQn6Ly8IiXke6ysdxH1lAoPjZJWoM
PZGP4g5mv4pZEe4nfCHtcrAn8TDFwofkiXHm0woYR/QJF68h/HFMFkpSzywZ4S+/
ePtCm833YC5QOPnFcpvhb1stc2yt6OP9m0YvG1GBA38o2Ypah0f2b0W2aNCfN3jD
x3pSnBcWy5ywnogFyRKjp0NfT35BChoLwgGvFm948VuyUONbYwfKH2zOn7xC9Ib1
kqYwJ3ADRGYKOpyRauXKJsyIBbX6OetbyGG2VXri3qRkh+8oZZy21EjIsRfjKn5X
9GcDGNjiMA2RccuCMl80+MiaC6MpDbTBVJdJBbxrX0KcEHxwpfMPm+7eiXZlGfmg
cL9DP0uBcs8AfPm97VL0sX4oQgQe0p+y0Ee61pXg8uT3M3fh50IlKUshYxqWr3c7
r6YhAYzorcrbcQhu+qn81muN4qZbRUgqXQNe+0CKSgj9fQpc4ZhFPpmuRzBMWtSY
Lk1ASUddb+jHucw2C8t5e1Ww0SnthVnA3VhRClSignOOZbdMCjfjGVMulOJr/FBc
V7G0x+r4OCU07yybbFChFk+lPQlBtypb3mdAMUZgZFuoyE6tfJ43YfpxKYz3tuj1
KThxqaOlIzt5gcFt3+dZ5EphmVJiWuSmhkEHMvluMXKnZbMeFjajiUf+FJlFKOwQ
CZoh8KCliQUvXx7Ac6ClwLyc7BuIY/46gyI60iFUMyb4wOqjUY3yO5CDMBDYuWwR
WwYs1LtIVJO4sCo8rfUPuxf97lUYb2/bw8SJTUyzIb43XzlEM6Y7W3gveQV3zEqg
lS+otHY86pAY+IJwEEUK9A1u/ormN+/mTIxvKq7lyIBd1rFQrIE/HrRI8La8snqp
oeBt/RrLO+6TgQu7SZ+1rK+ewWZexxhY7Xk0cEVNpdpU0Tga7wTRa+tkarPYIlHw
zT0Qn6I24LJXGgM6cXA9cWLoeoXFMZhHeGnbIKMNFuJQS16xa+QHdfTA0lo87RPv
+9Ot/CmwfxrsgdZJtPgOlZJQjOHBzhH6zswij2qWNsukXoxb6el/w7ySNVHhtPU/
856Q5kgWZfkG4mseTCOXumFyGuVja9cZrBI7wWwMRrBDDnvh8Np4kW1nWXlisXyd
kVK6NjDeQ9mzZMGgGiCp9SWIvjcAOrNqM8Zm9+xccsIXNYCHy/SyMXUAQGELvUCC
o1keH6w2b05ff6xIUzoLn8+D/aK6xCNbHF6tkkphMy3fdgU6p5atgD6zi3S4SsEx
f3kY3F1D429Edx+X7G7t4WAKmY94YH8rRJmILRa97f5ufjbB6jmYYedJESxN3zIJ
fgl++JqgTKq0X3GRGZQZT9jLB0ThhJBl33DT5TooYox1K9ZusgRjMQ4MpJV4kTI3
XwCFkYC++ztH5QlnkI9Mm/+Is7JsJhluK23relrBZ6URC3Ur5kzWjtWy9e1KlZGx
n3YT3QzEJRTN2AQl4ut3qNEoyNk9lJtZN62uLw/HPwKwIgKShX2Nme1B/OEP9PkZ
SSx6yawyp7+6tJS8qJmBsIMmSDMIj850zqnYKKGCYbai2niOCi3p6Vblm6O2XP5b
poMFDs9pyToBRtnDCnyzP64u0EJP86nvLh+EuVgPKg0PzAeEg2a4bt1kcxbIvQ2b
JSUl/QETJQI/6PQKUM4AGozyQ8n/KeJm/XB5KqVsDAJw91UP6+nW1GDzhH94pOtb
qjq4EkP4oVZoENWBqug5/6E9HEz+TVZ+5PfbQOXRF8JSf9APQsdLY1ZzbYysk4Qn
xIasc+6xP8GNzBevO93sLFYQyBHd/rFY4WxbixNwrZwOaUa25jTkcLNtzH547IfG
x8t4MVhJPa/ARCZwcBNfV2ZSRbKsuhsa/0u9b+lR6qcdf7unfDLYKvtzM6ZXRG5A
8aTRJTl82Gg/Y4nGte04Ju3p24XxJAFWu2YPX/dPZ8G0trfPiy1G2Ai0/oCL8K2M
F5bMnEabZhj9kqmwpH5Z8tttyGkNLhhYnnPLIQg86/XsOC9D68fj9rFh+9d9ESio
d3CHj+TfSiPjpFItoK8EozdgXlMKd/LzzptMtjBMFrdFrPk4oSFEqZvgwvk9ch/d
dTac5AjN9Ph2cMF5gg8FvX7m6rAgVKToIanQg2a5oYcB7njtU/SaYN2ZIxnfruPB
kcyUa1QGk50P/B9ZmfduupDQ0EOMc6DwuO3FWuekBkfk8TBuKQCCKi8/bUMvGacS
rZyBuUTUepF85afMuDkHKb11tPFx7Yf4qncmBPWabDwB6RGfZbgZdckUZ7k/22YI
LDxh9ngCrbwnDHCEjKKbUmSKtlaFykrkWYu5V/BOBvSg/tCm6sJiScKOT23y8gue
sGtqv9P5/IZc0y/LK4VvzJ/Zh8m/SVJkSy0qSIov7phzqg8b8qpnuSuvmjCbv6SG
bzuuuAlTdyDbMTZsYJkQOuJ2pTXM05jXv6Mv5fhcqn+XF07MlxPn1lBYRhJvTdB2
7mdQYuss5QazuyuIfNxgzrYbNdXtR8EYKDHZK3PTtplBdDLek/zuWnBq4iSflEBs
85YEsZ4r4P4g/eA08E56uhV5L0dreYQJD9bCa6X5ZP3Uej2c7NnEgpqQq3jlCfa3
rPueT9RfczwnOwu/2e2BffJtH9ItydnT+3LHnUZEm7wwpiho/QlxcZQ1EAeiTFfj
VgASF2Xi1tZvPupSlw4TzKaI5t2lBivDL2kd+EEaDtunzHIqkAQw/77kssI6qwwe
diFKQRqStcCVfQxeaKpCqf6zJPtw/F6FFx6DTv+JXxlBZLtOOIQCanp6NyH5KJTI
uRuAPpoRhxGZV7AAUnJysXnBMjcGgE9uFdarw2PcIUqOqw5OLEOqAsRvm13It8JY
/V/k8l43a6i5iUMeuoD3q8ASZxBtwP8qp2AkfhFGz5m9wNVSHkRWRsPs6HJgJ1nC
nndTUYqHtsRrYQlR8yxYawgRL7jlgXhm8Ra+G+k/Fa8Za588lB/2ji2xIABLzxV4
vSbPezVNuvvCEWIU/3F5Nu1I/3ZYeZG2sgjqx2l0dFrSrtbpNrabkuvd/4IHrgcx
gxZSk127KhtQ2cMZaOliDkNtAzYO8zUWbabQrZpbjFUVo6Yhc+B66biT2h05wSjM
wjtfdoaejXuLWOVy+iDP5OHUzrPWcP20A3ajL+YPG/V9XFsgW6kJKpQ5WS0Z/eJW
qYh6h1Pr1ufgWIcYPC8t21gxnOLgiMqx8mPwZBPO/mfxhWsdCnbpfEE7bB7oP2g9
V3+NgyVQX+BloevKqBWTsz8OE/NVB+Y2rP1JAujstClzeutsnFBFxHRa/JaPcVzJ
q4IJ+FeCGMBmh+onzxTWNWHQYyERJnvK9pzsoNnd1n5yJYdXHM2V+BPQ/tOV5vAM
8v2BT2WaAFK+sZ7DC0dPP4aSd5l+d60UDJjjqnc+iGC55Yo9zN8sVpMs+9e7bq96
VELqzZYeaoJQKr/Qo16PiAiw8CGJk/WU080b1tAEtKTpJhbgBDG7UXwfjfNQrqso
Cs3F1Sd32mBF+09knNFetA==
`protect END_PROTECTED
