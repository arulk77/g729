`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C1sfznOrDMUYuhfBO35vEFaoNKFusQiqYNOScU8nwkG0
8FyLO/jTtoyylayrUbEqRTu6CH9dfyylzwH8x8Hye0F489JGXf63V2zP+K7ivp4V
e2EC9toaMW7yErOZxHKuc2CO88wdGndT4R9ud5UEQh27qPlvWt6qjUCd+39OdB7r
YhpAYzv9cvRM6K8BJdqr7m4WaECcSuuWA6CYyuJy26/ZGdr+L6XZw2TnePrb3rni
XfDor+8xvTdse+6cxIZT31FrW6gPMBPJBMZsNWQWNf3Gj4lNmanojCrt60cdhVmO
DP3BMuqMJ/yxzAbEqNl6egHGNQ1cd4LsYLI4EEB/JcFXtQfmh1THpGE6vJ9FES/k
hIbtqoXgY/1hWmiuEz0zjo4yxHoXxBmzw+/lTSCHBC1z5zYQcTax7KZgbA3bqQ8S
/AGIsk2HeK1bHSUv9ZwVunBVcjRdZ3yD28+MzNR2MlQHgBsDgyTj+bNvB5Zo9kab
vu0annFrBJLXeiGcfuIHzCuLOzl9WJHxoLX2GxP/MgpFLIu3S/Qng5NkE2CCdyTC
I20GnTLx43P1rbq0Jbh86sqJ0L7f/PiDWTI4gSApqw6RRgjIRiJTIoa1dw5bS9WN
jXh3AstwoaVRHsY9kZ5SvOh5gmhnfe0SmuJLuCMMSxqnUHnWhCke5LsPNcMIIJv7
uhgTa0U1HQoRUPt1reiH3yZqoX8ltbrf7qXWbrGxzPwtEEdORtBKUwl6IuHrpHoe
PckZCTcyiYZpaEGQ2tCWIelAn5oP0xD3ZVx1V7i4uJhe31g18pbnFQk9S9FAjNmB
y1hVC2Z4V6teLfYQWIl1d6ksC/JwTj9SxAQ7lFtXbj6a2krJ6uvPKeeokSjHLyoF
RIKYClsTOgS7zgpCg6QmNlPjcPWf4rhK5NaWHqAZdhKe8t4AVKUCOaIRkPUcYa+A
pWy3EpbJGKFzw2A+q4s3E47sG5oA8X37gNAsvrRtSPU7crGJGplL3yqUirxeMWTm
eqqJLXlY6YLm59/NnaAHdKrr4Bb8SDm0sT6Xlv6tVxk4uhyannI+tkrqf/FCAMDZ
eR6lF0a5rtymv29tEywImwBI+E5Rr45G2pJr2mr1H3Wo98AdblooV4dPByAIA5y7
TwMbcifEvK0v6So/vLahx40dxT1HCuk1Ltx3uTCdl2NO7NFO3fzyyVegT1wGVKL5
3WU65Cfm5dXnQR6mUsq153ExbLOpU009DBoGDeEOLg8obFvaUla0aUBFMgqXlGIf
MjPuH6TMuG5qQciyZx7tqlwN5NVeGwE6PJopBsNwdIJzN95wsJJptjqKGj8Y6d68
iIoedvmzwgZWcmnHmij1yD/n+e+UyTpbbL3fT97KSI6eDoWZiZBEWSCYKfhc4666
PxRmB4MDJz3NW8/3AiyZusibn9zU5mTFwk9vGaNZjrUUsdN7iA/dPgmmnY2fAVg8
n9cflotyaOmamP4qpfvasKmA4lUmQqSfV8Lm+ASqBWmxja1Zl/c+oki/1XYY6pSw
xN8GmcTCigjr1kNhMnwR+evTsv6/q1M0sptoH8xiD6VyOJ7yV+tfLabCai2oRlGc
iduxiFUjYomMIBoegc1cen02R+tbUdbhq0drWJvV3rY4ySkQx9Qm9SvJ5rf9hMyD
cIqEDypueCGe2kKAaj91jo3sbQLENwL8oLqI7Iyc7Ao25T1R/dpedA0nkTjd4xd+
awteskWcxxhIrsBaC00tipWBc4mS3KRXFtQM3B2oCCZak8tqtI+NpJs7jPgP4+SH
Q6esClg2Tb5fh6GWcZ0XsBWW5IfKNITuzGy3PwHSKq5iVb7AuqM1j1z5IaylxpVs
HNdcWrp/Rj18NCDsF8j9MMdxrTb4OmSMakcSa2A45v2Qt8OuBL4NwIrn+OUp3zp+
ov3sq14thtnKjUimpzpwOjzM1hyZa0px3aloiMLvytfls0aUrOvGn4bCDbsxh2kZ
8FF+0HSBFBdQJhGD6y91BzjfVN4pc8B86iUnv0kQYSI4XvzKc2qgLOrslKUQ1jyd
izAd4wwfFEO3xl5JdVYS77tFB5X+WpT2N0g/Fq2jtDOagNllIUzN0qj2L0YX2PIj
WguLcUT5Hj4nJqDtTWsDo69eb42ErDHZgfHh1GtsUYGJgvrOuYXtZx3IoSXm4Srv
EVjdzQVniArSN8HagCtkgQewoYQqnIMeguZzvjajPkA7EGy1QPYC8+FKwBokSOKO
56O3jjvIA5JA3bpWPECSGdymYfq4pafK89Yd9dwVmrNWy69+GJX+vhrKVOySdDfB
IVeGzSFRia+S58qzTJrOfrwWRtVQ0k5QlQ1HDD/wH5XsfX862bt4iw3J4acPJUpT
5OrUtP51fqydHuEdNi45IOYdeI2ARwsjLIIzZqgba5+DnQIKw26taX0a+Hwbjqr1
KKEQIA+9wJ0vDYZiVxCivo4b4swsZXbgf/5s63kigCtRPr1HYpK0RqLyOI+0RbeE
sPMXuBH/x9MNhjwXppME2fPaDcxK/2wiaaEuIYyXUkIePxvHu0U1Vrw2BNkYGN2W
fERitEKF4TYFf/PbiwlCm/3rSAKBS99rK5+vrFmZqx/TJ1y4MrjHEyxAZNP3Tgbc
IE67DAr84BXmjbpZpChn1ph936y4e8ZzJ2jQfQDPHw7aTJMJnueK9yHO4Jy8LpNg
dm/fosSKknup7OcSo3Wajc9iy8dB87cRWSD/DjZJwYAGJ0YMCmgQVXqcFFNV2E28
UHocDxUO5rN4PrkFkINV6Gogmpe3tbTdFRwUBp3S0k4PoG23HvQZeELyKYD+l4T1
gjRYzLv22QOKPyQ+GJi4nn78Ud/HqdUNwPot7ThtnueWhYUWQF/gE3+hGKyqf7e7
ZId96N5JsPAWn6vcUDpyE+6Hh8JG8SsJOJifiU0ZOdvoRYdA11gNxDTLe4AI35Km
+szShcFGT0Ayf/XTobYlHK19dNLBssxmR3qIWYYit2Ag6+tzyytta8bneuDAAK1Z
+3RO1IG8+ptGRxzCILPHwpTHS2ZNkG0C2ymoFeEEsiOdhLCmr9ydLgdlUqRJ6SFc
ogCEyOgybak8ttUKfSdkS/i7Wzja0jBOpiCFomgH7yw7raXw5gC00Ce3DwuR38gn
RI5aqhOFCH4gkrhG5Vm0BiOJJH6W7U3q3NJHhybtIvDRdpkMfRJpvzDvE6kUteir
2Hzzsq0Fximc+4BXXRjNOCvkuzvWwY7at8D8wN5NqlC6IMV4Sam8CRHrj8m1YTOf
pnrofFSJUpJUBwoJQtMBzOloyEjRCbX8DEpxdlRwFazgNcwdieYjSJTRFRA39seg
IxWR+o5RDPf2vhsjZx5hhpyKxiflkMynxeVAiC7UgxDgxMlNpRMMhaddsWDk6LoJ
TI0dRjr9CuNCwisq+rxymrAwnFrVFpYPKuQAcl7i1Vsr1Ka7DrIXZvU975hYcLbz
wxB1iBdW8DzvZfAbj1PryVYONBgqE2pQ02ucO7a6tamICahlbZF2rY6fU4bMFpiX
lz6943uBZVcP1RL3c7prU5US8OnK7tbGIvtZJ2Tt3BASIA3c4Mzg0z7/x0wkBArL
MYyRbZ/Lh0ISKwD1el83/j5RJnWkv65Ul5zSYNJaNQ1z71+ady2RGfx9gWM5xpWh
Mwt8TzqkhibKyB8+OcCUH8332OiU1GMyKaIwnbkZA+ihe5i16UnsQD01+tvs8REn
0Io/hEgx184k2+i3P80fIQtI66ZETQq2oU++v8FbOOogkUTF1yh6EQK3jY/xKbvJ
oqOYiM3BMC+br79sx3dYU/k+75DhNC7Goc2fgovKiycM9fdSCozrHNjvMrMEN0Z9
NynyTCAOLQmqID32z9WMFre3Wq8rC8DjQzOFAURZlQSlO8BeWMsMkPHZlxq2TfpW
T8wuTQ8ptQIkMc55N1ZT95HXKiRrgjw8QijJKIX4saTOUIONxzH5JsBHxTDpVf5z
o1rBMjhV+pQ/waneHGbQ1/Qbn2lSt5kP/yZvY8OdYZh3Cm2ooihfx4/wrMH39LwS
w/7tiWIZivSJFUgd1W+2adaPog4ZpWGcMV/+HFeYozOIWDZqW3gorMZASUKkaml1
wwyyY8lzICAIAkZhAZ8zPcQKmlFki0XWVD3o8Hjh37LOMfLVYrXxZPiasovqCq5+
PBQsZHoosr492wl8nN1pLZzAtSDTzrZ1GxgNSIityhjLueENtB9cZ554LYvfFWNi
CMgZaAJnvEtmj8nZeSwHBXU7A4xkesGKeVBBGdwBgDrBmqEh0Cs7U33o8h6ya0ha
yLh0WUsPvmUwtZ+5HruRuW3e+Lk+b1b977AUinyLC7Ts5fRz88t27RlxvZrC90Cb
EWyrr/L6oYrnON+I5We5Tem0Ghoj3N1MhfwdRZ+9oNWjyxenGHpLKwMb9fg+oiKd
ie4SLqRqESTxeE5E0vsBcxaCo/8S1yDqF8Ln9EyeE8pbnxVJrq+I5VFTdlY0LJtU
mmnc8eQ0LPf1NuWz9hf2zwgezO9JwkxqK7xFR+/xrjFfP5n2GrwCwhEk4HciO46i
5CikVKhSGyEa5COGtZo7qaPKFjSt6MI+0ksGFNC44p497ZQjbIp+iaX14WS5VjWT
bfWeVJYtCm/fBg8vvdNoccjFM1QK4PH5GI45qwRQvXcfQhpK9TGt2JAgn4Ox4lQN
mmo/7SGNQoBPAb9n8nHB419zwg86T80gS8VGop+cdhTePbOKcgD0hYM6U5CElqCT
`protect END_PROTECTED
