`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
kFZkIZBtd9JT2XE4rcJ5sP08JvioRB01Xa2U9dyD7xHkvADMQL91rDGGlYMohCjt
jVbggmXeXyIy5m6NGMLdCZRX/lkDqtNSoAJW4QIKfKF5nT3I9Tmj2Qdy5s3rSHY/
85W/y+zrqMqCWdcnRubAIz5rOhqwlNeM5LxlLdoCNsEyGwTogxNHheG+kuTcsR5E
nAwRFDFDSxsauYo7knsx2B7I5ik/6C43aEhYULhSQ96YpCxZSxmwbLb5HL49e14f
1bACyKy9vFMK8LDdU4KrBpjhrMBZ6vuJaYdFisPZT/H9wDDXDI3nLdN8Qe5KTh47
aakyNLhWkDnEDUDJVPwUxPsTEbx3IiAFyCHmQ4YqcnFKVpoob37au3OMyo8TEB2n
PJkaWOb6WOSed4tN/f2gisGhLnT/hndizrcQzq08zjXWMkgcybMhoTEVJZnH6RpO
sKA2Gah4agEoF3/Mj4TTP7fiQa5T5Whc+IBWJslst7JRjOGLTYdyio59IbQwCW4C
V3oKDSF+0V32ZceVUmsHFRICsvFlTjRmpuA9B/8oNROfWLDNTxGB4PCO/EKr/nJU
qInUWcv0KrSRPAyaETTZpzM+5pwvSPySdXCYoZx7Ze+RDxQUAyLZjM05NOXv6UZu
wHrxE5Cc6TWJ1aMLoAvHexo4bbIv0ED4oLfMidl4UT7c1suCS/CbWzipqbKWKdO9
c+3MVDaxzVL4o4w84J86MprJjBCKx/3FRd92rrXpKwYFDqH8jgqUEgf7m3lSoc1+
4yUqkTVWmIBr/oQMGNS2MIK+hPk0I9/bxEZU13ZsQBqiz8rB8GDE9mFmJ8gcpgHB
rDeGwyv/B6U/Sm6FnebMzVZP3vc2ZrZmoY1jNDAy1CUY2oLWtbdTPRY9TQkNhwas
LeB0h5x/uXRUb7juvTndgbYZwAifufhP7bArBh7LAnlJn+DI0pBlOYEMfvNaC0Bq
G9+233TaacqjHhSyhqIFyqknUJNWFZLUW9CtPL5nW3E1By9AjSQ/KyW+4UQucJMi
`protect END_PROTECTED
