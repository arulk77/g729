`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40SpZ1qxy4WdrCqb8Vknt1MpRz0CbUhR4ZWKZms0ndcw
Qe2nlw7GysMOGJYxOgQTJ3EV78lRLEP8RVJUoL0Gmv8K71/TCCBuPTL+VfM3nAFd
l7Llg5FuNypGrgZRrJbbahtavFcP2jAV/zKzx15je/jei2j3+xxGc5XN1wAJtS05
cgz1ch2tilbRi225MBgglvnNJAweDdqUelKo6B3b+smnaK4JoNgyoyKMuGICtoO4
me/0A6Jk3fqoQQA673ikJuVl3EjDtOVJf6wIT1EhsknO4gOTQ0I6jy8tQBWxgDFq
iOiLl88U3BtzhAVHWPDNoMifSdd6NrYbYx/LUN9+NpoQElSUqMR/ZuHhOAKfkZAw
JZNmzHipGSDinR4w43aBiAaFtIZPRaiv/Or6rxqEVD5qrRAej+QqXoDsHr9AnroK
osE8cwsqcSu7GiU3Uq8NSg==
`protect END_PROTECTED
