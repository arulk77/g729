`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJJb4tiVLaAOVmCXRJfUJV71mijq6I4DEbYviBEg2uaM
qZys5XSkADc6zYTwJoMw9ms+7RXmgF8YQWN3bcjG2NmSUBuvkYbmigAu2odK4zan
XFqUynJX4fTgsA2OdIB+geqYuJO/BSlLG2pw22YeH/Nu5brpAITBlKCYtofXWV3H
fo7werIhubFpyLGJ3viXaw==
`protect END_PROTECTED
