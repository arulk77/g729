`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCTMilRj5IvzITiiJN5omBRgO33FN5+n5MgASbvmCvfJ
rMeQAjTlC0IXWr95fO5dNYFlP8hUd/WRsCzWySuaWTVrdPiJYDY5y+Gq8wVTuDde
s47rJydVwY98Rk4jBjvEjDFZEvmlXmiRcbPnCMG2htFHNSPRwj/3Ug6gtk6JyXCN
9knuPzz1lCa02ihEWp7tLKWZYfZMNfqUiOyCnZlHgxGkRy5S9tXhKtoN5+02/TCt
JpmoMCtR973nAnG8zEI9sX2usklYdAhXpoFEdg2Hm8A2vnHZh2o2gPCnoa5hQ9hO
7I0NgkZ2m9UJX3pFg+kIm+5Wnh6EUar72l4Rg/c6xNjuClMaq4j+oqHAqD5VnzQh
zP2agzMOn5vrLN/sEhjTycl2Rx3LrWaGZxthx5GHRyEgIrTN+N1X++ivT/ZIh1LR
`protect END_PROTECTED
