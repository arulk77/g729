`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1afJAYuYelfg0Sv3s1n2RPMHCe3dN/CSlDmlqb76XVfSU
sFFTkCwhCiJIJ963YW819WFBXhDxpDDAcitrsM1UWDT2gRukPw91qyVn4oEib1Rm
ZNSVaXSorrfKsBK+O9Hnvq/Ljge1kHtZatmBgraUAinWerTRQ9Ugi7D9/HKR3dLW
E9BWz+3WP4eg0Wjor/2+int4Mqg/ceJHgDL8TNsl28VUqMOAq6UauEMSukpEE5I4
pAAxJt13voLyvR6AGzrV7TkQ1/G/YW1JZ9ZQToY+9B0RLILvtwnF0DnhzlbR4KcS
yfOtJXtX1gDyGW7AdZ3xuXgLCYMZuMpvm/v05Jm8Ln9RLnpQvTmzv/wznH6y9Io5
+hqmMyr28cmKXU2Zb6S4WmN1dZY7NJJvf5nkUbJaCTV+zmN/MXBkjLa3a8UCm0lI
z0CgaN87z/Myw4PXLPILbn1WaxwXSzZGB5ZkIlnq792+yV1X6p29Bu7r9cGo+V1g
gFd2VYE3Zg4icBuKCKvGygviLldplxSPZMPNKKEWaTmk0FDpcLp2kQ8aMpGK7zfr
g7Kkq+SjvWUfW7/A9t3YFoMXAFwY0PSoetXJc2HVfZ8nmK8ddsaIGY6Od7LZgaEw
pFmS0r1dqHcC0CF0aJuFJgQbTtw6FjoEu8IoYheHrQZE0DYgY2yfthFvml0sVYSA
nCdf66MSaYqnpwdfZ5/oPY71w0PMqtx3eq84RC9cxzGfgCSKquC4IpSrda+xCsQM
2jw7LZctMQlgKHDyBRXJuhb6bi/C5xz2/WHokqHxyg1J4l63QT8EFqGo7Xb2FcsB
wL2Xbk5ISJN4PI+ctGQj2FUb+tlA/KEsYuJv498dtaPkgKe/L1ibbpeKupWBCKsT
vdSxVrr7Iu3/eisVmInz9TaXeshZBiQzjPzMVZOanF1rR8ralmvwCyQuc8GB8rs/
gtD9pLX8m0EU8Fue/38+j1Q2K7yB5pZ2tTMO/d6h1VqACF3mNRFitiZyH1petw3O
w90PWWs3X8CUWTEikFHrLPy4wuLLd88Dz4KO3F1D22q+RSqvEvP6qpVDvYu7yb59
qTYJT8SM4mrE4QKGJioNVazoyCS+tTA4Cz9bLpWW/sxBuyl+LJHF8pvQwQgGksQj
ZV6yjMF7I9xvqlhOkCTnnqisR4U5ZrSrp3z3zSr8Vl3+oYzBiRks7YaNoVpkAAaf
XV6peH76LrMHmmHlo/lP/Hr4bniHHNF/idLJxsan4AiztJT2PYzP2IIFQlKKGTds
WQHk/CbyeGbShN9bxFsDXF7eVA2rqun+r97nkAiycG5JWs3rSKSeXWH/WfijKX50
N7fznr4TnbI/TCoDhc0gH3b57mcbrZVO4M2LYLyg9s0bxMNQ1s67gAIe2rJtBlfN
e34kBomjYfcSNel8j2xPZW1YOBWyrDdv1ZDPTJSeflalNybGv0j6lkL+nFF3/VwX
XXDollSbIMI4BuZRY4tj/rj7xRERdeRgAOVuPCqitFy1ATDTTXS6h6bHrwKRXt+Y
MCfTrZ77pIjrG+KPe3HFslM18dsshCsDzIgRi7kIhA3GEqdKRJxPv3sFzHWY80AN
UkcC+o3jORzstRao6VERiWAErr9UpzqnKolCBi9WWm6yF6090MZt7lsvupzDTOXy
Pvz+qP7l6UgX4ggwb4ncOHBMylk7M9kmUiut6FSXj7KahLNIG05JT3MTv5bbKyRy
OXcpyFLjg/tGCJMsMTr0N5rfhia702WwJ1EXF5p5kksz7fkjSq7m/rFq89ehCEwP
u486SHHzZQTU1ALFGtIsSKUXmJkuU2t0P/F5OtjgdKURtKfsCLKssED1xUkzYvPc
`protect END_PROTECTED
