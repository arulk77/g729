`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEPk5PiQxbWzzV3hFfUdmneoukZUnjMOdNZMEjyqVlIY
fTNK4WCYN/akzZVEmgalTI2W2+scRFDHX6ISyL4rF64x3fowjKIP3xQYT1C4ie3f
1rkdk8y7qUDOWjBxY+acOpSmde5joZdY+Db7pcluP+5IkIz2MqzOtnWsUtKQ8tfO
I4AOv314WPduuZqCnVCyovCcr29gPl9H4cwIg6leXjvVL3sds5KQ/MMnPSGwALXD
jo5JYQmDfxR/Hl7wJsXWq/JBnz7YuEdDB8UwkLvX4f8NQXZEem3RUGHOJeoa4uDV
5pd7YFUdV72k+e9nLzEiUi2G5Ua1iY8/0ezc2PFT8eq8Aey06nkkpGf+gyIept6I
DLgIn777wfYZHYb/2L2jWi6qe7dyGALW3hwLF4vXTleBv/DjHENxAUNebwlXGfwR
4+UsjrCVXhqcj2kvbD92g5zCdrUnJjFOy9xm/K2anqkvJny17O3HGxpaTbK+q51e
ZP0ItLdcfj+Cdr82081AxbeoYFQ4Z9LxHqx6hhXkbij6J+I8sTTh7WjUf/JQsu5e
hrggF0Kpb6NAAnqW6fYBBR5PbvPuV5llfxX+nwFXPJJXbt6St/I7cR8/rRNuo5pG
XwUs2QbOzJ8Qj1KadLQ13tGGLbkI2ZFvB+9J7POMzYgSrEfctfwMjtivcHgM2luR
0o4BKENMcNAB2UeLzsu9l2etJDQtggwBUuiY7Rtc3iQIUZTaWEVMon6RnCqmnSAB
ogPoPi6HrtsAcrxfn/4zPU0+xs6KbzhhUo2Y1VlkTzCmC7LpSk6u6wKt0SBepDRH
klXAX58FAMYfNrvFdAmgIKXUv1FnO4k6HwH1w5W7+wTcCivSH7DmaaQXxArk5F0W
H2RkcCQIq4nBSse/6YBqXbcN+gjmX11pUrWb7hzbYqoYuB81wzwb3iSjbFIz9cui
pno0YODEpVpexqe7g162rUdHzIdiRHxHwwFNrBri0Bzl2xL3dVDJrPgrrDXan48w
2T+DK3WQpwP/rPHIcIykviShYFTwlLDuw4R7J5s2FywGCZ72xhPQD9FrpLXAFJzn
WfBPPyZVIj9gJRPzluYaDNMJ6/vkPEpq7NjXkWeeX20=
`protect END_PROTECTED
