`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKS0TxVgpWBWySH059G6TRDduTe5/XghBh4t0YQYmgR6
GLuqMj2L77mrAU33oaxyYBM2na4w56zJO8QLK30o5SRFxVycZRGaldUB5HOPx2JY
GhiAQbGDM0lnZHn+CDAyjYaRj5DyCeBdcV19i1arIhFA1PIiqzIdTECNdgpCR0JK
Nd85jrSgnmiOdNRgc5lIQfnSBEsaYn18wuqKgsYZRGCJIInV9AW7RfP+xU5R9Cdg
`protect END_PROTECTED
