`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNZcAOWTt01zcn3+GwOBMQ9TGth6ZdlZ1RHdsIdmdaP7
fDmeai9T+jmQmNhXGoSAlYbMx191nDU8WLs1A85UekdtM8pCQU6W7rBrxoM6fpAv
Wkp45XkhiD1zrZem33IQR9hG5l9X3a0Kbndn85BbfYqi4wL1UzlYbxU8WRi2enBE
dvs2m104ijFR9gHyARu58A==
`protect END_PROTECTED
