`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+GAoLsMtX1TFWnQiLCkATIVsouDpOPrEgJEI7LHrb64
J+C/2+2ZUVeI1qUuBFRX9S9f0Im/6G9adjQft7lWHg6n7cXqRxk8iNRDgBiZOGKS
BVrxJA3x7MFhVZrIR2sL56dM60OSw7MH/zmRllAJANwArkFqUIH1VVpST3DLk5BU
sFyuHQURCrroDoKHAiXCH87VWYL1AlXTh98JBsSEAa4=
`protect END_PROTECTED
