`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePh6inWZGq6fRmw6vE05XU5oFJZU3EjYyhdGtVPjzeV7
wAtyIDBElBkD7tB6gWrcyO5FaFCjhDwNE+N4LYQjb17vfQIIp5Zq0QOFrhk04uT2
8vFLNV401gUMOFwvXbGWvZDS2Osz4bC+0N74+67xuK+/8nAFZKagq/kns5/4awmK
JRl2IdGKNMr6WxnkYQeT782YI0BfEeGsUX68zna39lJlWE1bb/96cZ0cTgkJDHkZ
lcGwvmyYRKPyqZ33dXOEgucFW5W3RmBsme3io6Q+/4eaBTDpswC52sa4LK2VjDXG
1zGntBY6s+5ecQaUZxwAj12Sf8tZfJrgG66raRZIABU9GGrgwjhvdXnLU6zRqtKb
G8lIscwEjx3McCWaltiAmiR7TCatT1K8oCQf9ODwKTykb3TfWmPj2Pf28huy5oLL
cebE3LjxtKa+xR4Sa2PfTlpAo9ETgCQOrJ3khNNdwHLYNvoIVKYuoBBY/gQJihoD
sPRkadZMt4pm1g1pEBtT12ZgEOcEHLtmj2KUd3wL17cQZzX4gC1hEqHJ3DZRmt84
SB5nQMlXgLbydtn6uEqSNdMt9BdsyvidQdYtYT5gEj5vdVQVK9D+CVjqG1Xat78A
/DBcfg56jqMPgXRIkeeBPSpukb2nM9Mecukl4i3PF53MXMk6dEbWQp0Ca5sL+VQE
OUw7sd/O6/wi/An3hSStm4jBBf1IujcxAKWkKzbGypwapAxvH+Zj5CNR1UjRlEME
fQcfVPqZFEFW5+pwML2EQ4RoseZ4i0Ail69C1Wkr3cuWW8A0pxRAkmzjw5JxyHmb
Ig4I7WrHvVdtR+SP+de6wLgdzezmrmjiqwIEsaRfyYhmZk7B2kj/UWk6HmoOeWum
H19RUQtsWwk/PC7UCeN1yV4WeM95O1meAOtsf9hjXyCwARcg+AGPLamFm0jfkt71
7tMBIzXswRxdjiY8/8XizPvecEq96ZSuUliO+4rLW0SPIpiW01hU1ZojqjBNIesc
4BdYYUmFGTH86e3zGrXLhtTxJSHoLN31j3yj1d9HPKwU9vk7jXxnh3OTBPVxS8ni
IKUdICkSNgD6NhV5xaRz5uClPKxk0SgjxqJNx3uQjqJYUeMG9Qu8O2BLGeohH7EQ
2v+OT8Mcaesm2AQCFHbuwRBn3RL4MbNTaZUBCECKPI01r3N3xo4OZZRGWbIcabk+
hwwM6acy2Rd1ibq+eZhAmeWcgUnyZNLVwXes0kIRxxnkzIgY36z8myeLs+Y4No2J
eFZwh/oti+KwNLX0XQ8Req5WN0OfI1+9PdUfo4eyGEy6jXoY7Zcz6VRKWfMIgE2Q
`protect END_PROTECTED
