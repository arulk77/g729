`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C424ZM0coaEFtQpbvIJxwiwx4uDIohd9wZvpn8jTTN6b
ztV5YtD9wb5sCfakR1mCOrZF3wu/bOoDcLW0aCcMQEjotpfAhNMqtpIT18+2NsDE
+EfJCTKMZnMrIiaxIVGJrxL20vdOCeZ0oLvYaqyIk0h4pT44raFeA9glD/rOIlzS
LLFiH89tOBmWztKbaLRHekEZCniWV5IybbHUin+mUiHGAllN4A0xcM4jlZ/kYPjk
87fx/7ILLSeElus2ZjlR5144np0wiOwUmC91VLmx2MGIqo5jI4KzT0qGQIgDZ4+0
DzFvv789uFM4/OI18Ry/SOz5DXGrEDqRnPu4jYiFUKeZjsdfIJ0MrxtI9AkyQRnL
KlVxv+jyExjGMWF0iuNS2G7sjwuOIdFoaVakz3DEUv7D/8qziTZQC1JN2WHCM67l
/KE40ZgAQ30+qWePA/Aa8VXRdy+MsT1s3SmDCfTyvt+WMdgtlMkVS7gPRjExBFcR
guT2c6qgMADQ1g4tXPQcssDMHLgTT9tROsYsN7J7Q1IzvuTRLSkUH94+CpHRPbwS
pSBDyLuysLL5nF6SM8VXX2WHXsrVTbiZgljohtWGwBwy/oMr3GUu5AQ7XHkcrdj9
vt75X4DgM1/We/lUiaqIOLdcb9nL2iI5+LhyOTuP8TNPDGxkKS5/wfE0uYr4Ok5/
YQSvFTfj+JZkWZfDlHPAlZ7QHKDX7Ei8H91qoqooYK8jOPmed+Ol9j9NM8yiD0//
rpwiw93sJxBWvp9y4FBcwK/50/GTi7MDNfY+tlTa1Rl3FkbZ8jO3kwJb3BJQX5eE
C0k4mszHMSCUqsABrdg9cX1GF7YhIEKTymBpBkimHY8/HHoCWgQ82bIae6c29oCi
X5y9RsuDLKm1sauKI+d4bquIvaB7nabKATBXp6c6oxhwX6cqcuQYt3elMvujnflI
rxy5G8JSgJ8Se5la4UymEHhX4BWZVnuqjPer89nHtY+LCALtwETEG+Id7kXIKnHJ
hqKqqnbqQtyKBGHJUqIIz7JQ6CGbasYyJ5vluaaRvoI3Uqcb+tYnsDsYAiW04cAc
KYpqAcLdxTv4pqB2YcJiqHrNjUjLhJupqn37o9Y3fZFphbHP6WbK+/u1rqJxKzEp
JZj3ji7wnnpfUx28fhKR/TsTuD3vpB9najPbx3KIFXwcbxfk3lOB8oNiWU+zgrut
ZF4pD5RTWnI84EDaFZn8J8FYkdais1WYLDhYCOdJNSMDV6vRVhwiHA+ySka12unz
KTq2oLLlaNvsyTF4SWcbXtrFk8frCz3KGwAAKdZsz4JQ/8s4NKI1xw2Eomv+Vg9W
7dTeQlGsNj4F7zvUDpKazWogZKGWZefgo37o71M/OABrdEMAtCfttyLiElvqnxTI
0+j4cA8/F7dbyfEshddzpzmwY9m1k7Kc+0rvucywuUFrS6WC5wNldZGHAua7Mgm/
ongO6iLHRRyi0j/fEWGo0ntaDHCp6FnnTyqlEUMvVLr3eF/ZFI/3xhOgbzztlVeA
gHY/vSOxZ+xABXVzDx7jncMSCLkSEPmLyfKfIwF/kFyDmRot1L0Xjxmkuzg0T3jk
RD1eoTzhRdmkPO3VLcx00jqIX7XYQqyYjl1XgYraoM+HTszZBlaexjZJXKTVoo7M
5chGWH41Z269Xk+x9zOF9eVPVwrmAr0NjjZxwNBH1PsWXAVkNnxWcbwubyenHqOh
0NnJ7iHqK0wGex/Tagg5vASl9V2s2uUuaklmZ4/zs3p8mK1vh8DrWWF22U1zix86
qu1xWiT+oYE33MNQuHziY+IFZSa7Ssrskne2UAG+E239T9+EeA4r4DIHlYTliN08
Qgza7jFBNle1G5ggq2tFqJHMkiwS9FGSpp3CtTjAVjryUjmzHxksWbcJJorv7RL5
T8u6YUXRza1S/PNXQc5vpV/+mvAFkT3jtoPD64MXVXudeArl4QZGmqdYOwzx9hGv
fxCURMFzRHH4BONWHRi0eIqmzH0h+VTQ4+9vEYi6XHRHXUykHnbOpP12Q6mIuJQY
jm1cXhsHiLRUPE8MyLmdNLa2TeC/fJ3kjBAz75GWNSQAkM5UGacTtrbsh+Im+J+a
aZFOiFhnNLptqbTDUE0kAGjrKs7nTHFRTI734jNgtRIXZJfj2AO1vCo2B2ILR7IH
NE8UtIhZI9UdLJ9Csh1Vy1BhDGB7/ZlbcoO7YUpIc1P/gesqHpgPWu3MucnlsWWi
NlAGEWrUHntb/4OXNW9oDRGZo2KuZ92HhGciAdCSFt9ejxqPNBJwmTpzpN38g7Qt
zBAjntrxvxjaxEIneSR6tklQcJrmIYWkz+sNvpa5gxaWt0uRwy54ybVvMbKk33FD
RnRjrT7DMH5YtNgdg1AfQ+XMc2FauuE7FQt2T8+Htt20Is+s6MwM30W6RbF3sKkr
fR5205qn+GXMOoiRdLVskLoTjHQe41ve5KoRK9qRmGwIWGLHYdxct5edAGPFj92r
QE3m5tKlufu5/0gwu1Ld8muCD0GO/JCznwVksxoq9gktM+2Mj9rgKIODWeCkAhBT
KSKl9Zu85Tl6ee6ighG2lMlkyvYYwlTWiGNRdwp4nVqrgf6ga3H46TkKYXdKTfoC
ezI8+DJltOgC5YO+4Oq6CN1hh3F/Mu3LcWNs0EUW6ADqQyWl7Eq9r6qBYh7kUS3j
Am+eVEVPvQyOWm5lGmXPdIgvTzPptwD/uAmY4hH/Y+Im/LktMxxO+ZXaWLC6sWOk
v0LDGjvt5zeFtk/4jnPvPbowO2PBmcDfur8sQ3jYCFHscZ9fcIXd53mR8XvYVslU
Utf/xxD0mxiFqdMDPDYe12zAoqNdfJF5p1aNUidM2QgxbqzBnbXs8CQN7MwtmYPq
ZJRvRe9Vpg2w/HcNIu7P+5WclwEtdXv3F5s8xL8Iyd1L7iy8qZZkx1iRNwpgN1tN
jt5Wj7QUJmEIrc03fxc39NyMOKKgnhWzBCUNF/I7ml+kyo91NbtpqazMtCYiM3uq
77DiDSn+SG/fdkxSJmrfuc/BSf/ZCUFV2a+LmQ3yiY7P7xOsfWrJ6437BvlYiUeB
qdqfnMBor9ExLQ419kC+9OuiRvxXjePPc/5nUK4CiFzmJd0qeCbalHRHXr5ujk1e
Iui2vcRNyn5ndMb8DeCgGaymeKaWGYD66n6Ox/JUOYMm8HDrKB61jHpDNF6/UYnQ
ZpgjtCvDhUORzZqBIozRD+7Z9BV1I4TLfSDIzg2QTVtgupfOGwMQIfg4oMnodxIB
knJfFXEoEg61ByCBD3zPuw5NDW1AlRvGqGQ694sfcolw8Oj1MesMA9IfA5Zp1uMs
OFrKsMzXpfU8dNMpep3zLOhDFx8+iVJVGxLC4RkeEkvt0uLb1q/8Ba1ktK/Zikpl
`protect END_PROTECTED
