`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveM3N7bGGs86kyGzW0tTDii0eL0FIma/McT6O3jNzigBS
9tmtkN8Dw7geRSkIVANxxnfevZX3NBPen6Qf8BH7trHiZyK9ers/KGxZ4PERnMHu
qk788Vk83M8YTtNJ5gxb2G9ppKMLCiYfWQBITxiYfM1LXw1FgpHmNijOb+d+8JeT
SW6CiWymeOaRAwXOz3Yaats4WUkdvsmP+1YBXWbP/6+RYiz58RwOyhFNlQ8udksN
`protect END_PROTECTED
