`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+QVxjJRdWjkqAxrOeiUVSKqf11Gjyc5VtN1raAVaDqP
bFVVZNSIvmSqz+z/0s1hbSjV2taprTb0HIEsHVlA6wVjXsT8vay41Uur/NxZApB5
I0KRnYCu5bT8H0y4YDmrHhPPUOGZx66Fy2Hc2Aer5FjAGvoNUpsjn3alu4ebgGXt
EvUA+66OkisqHhuKast0otLYUe1+LIl+D1OEDGDGjtU=
`protect END_PROTECTED
