`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAG/JU3WuA+sjAKIE6AccUGdpbkYXDhL3CWNkLur1CXK
VfM9ZKcNwVG8c9N/uI2Ajx4Z/HhuH3yeuQGononFppuXd14qrL8SOHHKY//n452U
O9DJd3obq9SLucrWMj1etWqgznDswwbCpsBLUOSrfS3hXizGZkwUezm7mpoUUXxq
fPAKpTjviq/EtSjDIdHO9robyP+wGs7poWi3thJRt0YBSkjA8uD5LHM61WpRgzxn
`protect END_PROTECTED
