`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
E+hqGVEoDUXgwwT83lrIeM2/HbZR6dU6shVOmnG2OKWvQuKwNS9snXvYIzRMiexW
R58AHbkcNSNezcoYB2oGmDxb8aXxeknDpSHWlrPVhzSa8+QjI6IpYUz8pcPP8zU9
w1lR4aTyVXGLTTVmihbugOCDuBnj+VY7uvdSjO24xHzI+ulOxnVrEUWDx5Uadt8X
WF3scYOR0B3CxOLyvrPP8YL7Umg4ShbUjhsRb5vLYvEboDJOg0v9OJB9Yf9lu+Xx
`protect END_PROTECTED
