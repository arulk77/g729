`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
KRuRc+xnCKrD6txj+flBrc5nN7SnAS8mc4zAoB8QCGwhNBa5IbUoXN4v1y0gvpHO
mAcYWvV5qvHKpb3yWalzRE5pFdVk8X80jFUGB1spZCwkfRU+D6pCxrTZeRbm7dA4
vkDPiAxZX8lLBy4KwWAI97V7sTHry8mg3sqJhJpeqStrY0GTEEEUt+b4g66tRoFD
iMHeRkPbJAiQxUo97NTLsI/MPPJJHNp1ry/Qwyjy5Crpy0fsPZCRiuue9L/G8S3n
4zuZM4ePPcM9zfa5PTbSFeDHdSfbuMXF8u+WpJx4toITXnn5c7qeYUNJVioosjv1
38bKhARU1BOyNilQje2yr2re0eKVJus0jQvom4ti8WERKZgYNmWEb6GMGGUzn5Hf
ZTozxEGE4kECDwPuZJGa1C2FmqK6RAsmEKaj5Xxmp59wUGi7A1QxpATIMUwHxhnl
3EH1YdNaWHF4n0zvvv9erEkgRQr8W5LbB2Qp39ikrDeSPRC5xRwoBi+hOVkSLdeT
6fPp1ab866pgmwneq8m5wwOGbd1Mdz1NDESqdb2EwwP5BbPRJHSbpxcVpjTMeD9u
r8zwPIXFWmXFOfCwNKjeiG0VKc8zk+oHV4tn9s/Tcmt4cERwC5u7wsNapMSVkL+p
BbA1/1L0Vte4nMQafHwTP92ZzPp2GQW2ulp0QKSMqFPgWVQM6MvCct2u3/ZRjvxJ
MUbHnTf4eCvZLNeowmF54oz0foF/+NEZtvq4Ss4+xZfr9A/27+PjUO5GXa1X6rkT
0AzU0oAOkQCdaYzgmyj3maruJAMYZgLhFCpk2w1ha15kfV+rlWmbLifSBYkimeFY
EStSIPJ7Y5JDWleSZ76ind08YZgc77GoZlWcbTZcn4Dufjfinj8E75/S2S7IYDcA
p6oZ+QOm9H8Z+rTkMvy1j1ewlXtyat9to9jTQvSX8pNTtGNd9STqNiuFahPrhwUC
sHF0xpG6zMLl3e1pmhHTNQZGp6WcvHzGvVgGxjlywgjG5VoorIRHdXmWMmzbXw+0
q76yhTlAZauYbRBE85CmZeiujvsevH1e7pYY9HFxTVzLRmf9ef45jYD6AYGgz2VQ
hXdYAoidnUr1cb/1gALEGkmFBoB6m6Lqsd2awjxv168F9edcfDUaZxtSQBqV3Sm1
NaUwaOc4E1dhINcOXTJEm/34SdShX9NTZwduD4hEvmXeEJiZbjnB3Q4kHXxIadnS
ResKfJClNs2JjgHDtkwkBH/2WjxukTYfW0E3IiRGed4kbMkNV1EKMCrDvcTK+08G
z6hMroLBqu8SQbuQ6PWwqImt9UY/sGifdCaPNKy9rgUW9GwaXZOeMib+fQy2At0r
SHIDctagwZWO05ptmlEO5NItDjKkw1gj0rInSOgZ9Ur8he2MQjLXuo+GI1npHz3k
uPlWLBDZUTg78IFIOXeyKVlDzezliXhIy2CbA23C4khUyDUJse1p0tjvbGbTsldb
DLS2OQyv1ec9FyXxLnEAOLe+mOjvxlRWLC5I3hjGVbZvzSxiMWHpGaK/sqs65F2p
qXv6gtrBpSIzkcYtx/OttGxFP77+yPM8ksOaUv1rJ1PVWGBUcgiScU8aOY3GLZTh
mcRXW9YGj2fuO9mN33TqeuLfB285JYmnsxdb3ld/3dSlBig/uWHWyLpRrTuoHI+b
t/c8ZDpjbhlsbuG0KPafPj1lXoGLvMaP1TEK+xuT8jxT8ccYzVHdVsGPd2nAF2gX
42Ym8GiJaTc9HTxqLDh/ASZdqU9TOqkvTCEizpLE+6DyByoE+OYZD7c3uRJth0kB
zzVVWJ+7+XAe0m7tsNkRB/tBNspVfT0RAnyN/u09TzWHOxiKEd2MR5+1YO6mrq1o
6gs47XrcKch+gQ5xJFTBv3xSgGzH2WF+W6Mrtrr1IBIgjX9uNAcLNAzKTr+wuFvv
VWCAa+Yz+oAQKS5x4wqu6zOEqxbzZaJj/cxJDnq2WJdmTiwtfckQKWGQqru1gY6s
HUtCmV5ZuJ3GsaBDQqWoET9k0nBIQJe3VyA1BWb6bkFxDd+Jb3mqX3aCPS4pLvo8
9+JVZBXPtdcJXa7fRZ6acGlGYU9orvNbcbnjblU6zIu3Zs8MYfJRunpOWE3fxN+K
Z4DZbaLWtdYAyqIRZxdOJLo3FfFj7Mvb7B8Idv72Is6IfBJeQV+t/5BFRy8TFdjW
s/OAmZ+9px9zIEiROxo8ltomb8Jvc62CKGw+Mpayu2RwchwdagnGQI21FvHB7Mu5
jLcDD5FblIoIm7Xzpme6Km6/lBG2nL2VB0MZqtmSQcv3XLwgYMk87RO9DUtlYU0h
rmE85q/5TWwo2Ok6AnP2AEAlaTtPAvupY8ioN8YoTlA=
`protect END_PROTECTED
