`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAVVaGCgvJugt2M2wAxGv+PnDBcLRB3kMQO1sMNuJerOg
bpGQBhRckjIA3rbss2tMZTUhINqlbAt/EsRdoLfIXC6U0iuETWLoAW0QSsuTaO0Q
ep+kPorVcOh9GK81Ro9sFuYpbrQwlBuXaKTtYtAqmoJbWOe10gUzQygXWnBxX3Lj
vHQVuyEMgSCB8XReWHaKMZSy5oKRrXm/46eooSJLV4n4Moc/QqXStxUbr6W9iFx+
2J8BI6ILJKVsLp2no/M+6X5EKPB4kYm201q126LbWDxZKbuN00TBQf0cmuEjUHyR
yf+JIVuHXYlOYp2BTA/ofsRlCpB78dDnoqitiSbMav+pb36FD6tUkCa+xmkc5tN+
UYAX87VGxPiBXEO4WGTbUE/nTy0s5j85YRveHDYtgMjTTMQYR0NMRJHb474jLPIJ
4eJ8ucfljjoPS2Qmx7Y24lp5adlhd9ZtLQEOw7hOvJTEF806Zl9Nzdgde1iERG2Q
Smzn0vLsZaoongdilM7Guz6lwvhKTXpZI9PmKkIC+M+xJsPoBpz3uPOgzBYQF6DJ
5zwEMnNdRyiX/3D0J6VOhzIx4VvzNhdl8yW/UZkO8XVw6cIZED+zQXFDc7/6DUkJ
TeBX5DTgz1ITzR21oHtXV9IgHnmnzHbM5ScI8UC3c3e7UxqT8p9rMJrUu4lbCTiM
eS2TUeCGETRA82HfTp+PQ37BOyfNztZd4rVo7M6SqZ0SAaliCAi+9gv2rSU7BMOA
0qcFWsFkqAvinJoX/uJY3psT6jIgB9MEMAQHXvxmptrgM/SmfKbzfq2yZ/wpGR1m
kTNORuKk9eRqz06r6jIym9bo7pj3ITO6z2HuzwUMOc/znzS4Z2aXiwwyDJ+uJm56
xbM+66Rm3L9NAWfMGzxCgEF6k9lImPqP49WOWZPiVusy9Gp4FwgGAE0+garN3JRs
RwZ/h5bFjn60d8wOs39p1TPbf4D6CLnO+N7EAsZCL28wcIxa+SptXybWZpPTDIZ8
uxu8Gm3Ej8LXUCWp3/7P5TvqoG7xWdvTCJAftEzAaXwc+Fv0h0QNQWJGCog3CGNi
OMZst4w+cH06N3fRmOAxKwrIqEYBXMLy21NnZcTEGQPvINP5rWH3lNezgoeIJG11
Z7FhiXAZ2q48pQPZl7Fd3Lwuog3Wb0IoipSPUKvHBfCxbRPMAM1Wuz2KZUjehqv1
dnMYsVXYqy5cAmk2gsHdoWi2fSYubkjzb10Yih3TiNbHxuXgADxX9386kVePq79r
NirOtZoeacJSme/DLWcvh+uP4F8y4eCLo6760K2aMQRSI5Y3mKpHTeHoGmh8IZ3N
M++4pi6HAdEpPKKUggynpm7Mv78/MKVrt4IxTHRPI08slsKMBT4cTaRkzCMF+7+k
ohI1j3hH4/2utV0IjF0TQxxP2EOtZWjLugCO8bD0ciAH/HyBhqyppOCKazPa0nIJ
DIyxqb2NkSDotRopBE01SCBOoAfgO9Ho8ETUKpl7QpK+AZ9iaoD1HAgok5/CxgrG
qIbH1aPu7cGNhskv1dP/3mrtxYI7lAn4d/0Kvs2K+vVmN8Itgy/X6dKLmGzN1ufR
tvsxwtC5p6+KmlaMPnyn1E39O+jTPviZIWLJLEqVMMDktDbq633SM7bhqA+IlaRX
uqieF6mQkWTqegzVwpyq2+wqvi0QvibATv54ZY1AdO9i8X83OF7C3UijWrUmQ6T9
DND4gz6ZSxKFrDnKuOIAj/N5/nDbym+kmLZqQpDf/rcg5C+60oUL2JvnOF99Pdcm
mDPxhPKeL2wqI8QfJdh8aC9xLPaZUfst9Jp6uW/8ucpCCIsLcnMNkWtKs1Llr9rU
d3oHZnntQ9Bv9ADgf9rLzpuNvuqErFgGgskl/XxPtsYxbjnof1cBTKrClRYg3q2Q
vL8XsEja0rDaQ0wfdUUd56N1DiSIk14aSvwqEbzPEgKpgoHzNxtrhrExiz62+39L
Lb1EgBVddzdscFbzSYlRoMuxrpiY6/aFCAJVlJqEGNJrL5e4ifpqepEIFLsZTudw
S1h0ESKpcQg7THjDom8gx0UzFZHL7F0qDX4nlLsfEX66cZBJi37ThhwgxSMWTH4o
he/iuGY907UZ1xa/wVOCSYzoFNZ9oJwKEmsio9E7nYotDx3pKK5f7EABzF5/B+Fg
qDt868scQL+NoJOZCm5CUWDvVw2EOfxsQnspDkCKe+vhfKQdxjj/TpL6V6nkWjuw
2kXXUTKFEweSRha2vzpglJLjo38xjwgrFfQ5u6mPbBWMEK4C9XnyIqguBmk9gWJQ
UYBsgXk0r37YGGDuEaEnnp9WRBIBVlfNgKy5vxX6TmkStO8071isGjQhJTv4A+ov
sMue8bvuXixChrLs5VUknRnu/NNQ2sximhvQOo9MXyT2XaMD4E5OHDI/JoHNC8d3
cXmrPQxtAYyYpcQ4X6etnxpq7wiFk8zzq9X8tLY5W52jnbkWtknH6omrB0x6ThZ/
0Fr+ZyEX6aO80RbsTzygEaTSlQKUdqZxfwfTHa/zDpK7CskO0Hqr0/WeBLkI9Hc4
IzukU5hClcBDVl1WC9gcTszvV1TKC2/wDaeZu4PS0gzh7FXhcFcGM4v51d4fT8W1
M+WF23IKkA26h+MZeDSkGcKtWn7VVz4NiBGVrrTava2oIySZB3wyIrEJxcHq+Se/
h/xklYRAJY8qHsidADFs5T86XZhWwBucMSAdJhkcA7cDKWIEzQePSSWufoEFq4gq
WY3wca3hJ6WrWk9ZlbbOw5lxcEWHl3VNl7C+4khRJ3nn7zjMe80HesGET/a3p8mt
7xjeguucTL+t7lZnAGGesS/dn0iIJNYmgguWC0JBU/yCXmFnksNwgkno78uH+Rl7
/abr/kQokABuYazgn95Xgj+csBixpmTZ5fgtdavTff8kNMf37LUPssEy9RhEwRHi
RQZQ0iqJ1SV11Awu0FTsG1lM2G1sN6HJLzVCNW+3C54y0HpirLxsgODvHU4QqDaB
67hoA7XDlusY9A5Cz8J3xao04hh/9Z8Sqe1rKN42bGRzp9gUS6O9ZPHSMvUvbwlq
AUggbZuw6XXUsmgau/yCBR4ufLeZtiHDdd1AnRy5U7NCxWGgW1FD/17TisPoF4nB
h6R3S1yNBWJvSlnBngL7mR5ATQCzOtDas7IptK0EIQmuDGrhkOfzgdSDwpxwhShY
oinOjyGT5/9iTjrXngbuXrZeWZWP6AxENIjxm6u7hIBWpa9eI1Cgz2Dq6Ga23RXJ
FULX7ZXkd6AkcuC7r2QdfI7nbY5vdBy23UdP/clZjCud57sc16AghPP6HSX2egI0
eXwR1rHL/xo3J2AFPKaSwUIAcSFaj8M94K2RQFuMGP3mTc3LFgLq7MldPYP0ddQS
jGft0sQ/4RVDic1KwVpJZCOJSSX+KFSyhwc4XmnfrsFDMcudC6uLp7OIO5vuulmT
R2Hy8cvBGS4KzjXUm026H6ad/gLNcAewsuESful4jJzHhFldYI7bpbZP9vBqGTvn
QFhAm4v5E0PJLUVG7ml4jd0Qz4Zm28bcimyVItoKWQWsZspW/QcWgda4eCYjmUfO
HrptuaIahUunuaB4mk7qqhsHxZoUmZAyx7bBty1iy8eq7BDzNy50LrVrdd/MnNjH
SNp6kRl/LqYoU14Wt5A+wDqHKLQDH+fW2n1A2qp5qeo1SXci1Zpeo/QJljqbJN80
gfFY85qzL1NxP4IUl0Bvwck+BeXcDXMFG/8iYOV4dKiCZ9COCVY6Ejam/oskADYG
wXOOXSanpqbUp01yyOgNwX5F+9NO3RBb0YRyj72u0/uCQDZBjDTfXdH0KnnffDeG
aYBpArvJrJZANHr9ByL/LI0T9hOToFXHNlaZ+ByjQ7dWqHnzAfB2b5/tF6tV3iJN
ArYNsDceNulJ3dBVqTkJn4fQ9kv5O1mbF5LRZoDNAqZMNMPKsTj2KP3BeovI4t1K
zyXy8AmpFT2RW/kc0aHybNVREmuet9jRzwryb5IqxDZ0RfoI6H9xtTaStpxF3t4f
gClUp79FsQEZZqY7o8wyswlnzW+H7K29NqxFwbB0HO/e0oRSgl2Aa9LPIvY2BiOx
1G/7ve+5d6vhf8qn1zwb/C6/Obzpn2uC8RABK3dlP3nCI6X7zGuZS2Mjxip0K+Km
5DzT985Z35kmDKMNfAPVME+9pbl9kaXaH3h7qmvOQ+fiiZR5GHdN886Iy6YGLY+A
x2wLqVz2F1Ljxn7i7xtt9HJ6JIqdHE9tl0G/8PyfYfWVto6DkBMYq7JD0nmz3NTu
reCA5Bh5qH82SJsiStZA4RF0w0AFH08BMsKhQ6wzXhopT50R8FFn1wWCnuPzvuM7
q4dri7j+bM445K6OnR39K8fPEt4KX+Hr+kYcInvAiPHuIb8po07c/xUebhb68x5/
z5i+mt39cTz0k9beDSxEeAbZ9W1ld4qkXs6+u0XRWaNQfL6o9Jvy2jFqq8u4+wt2
xq1TJqE/PutR528P2rNFDg7/wRRTwQeNzr69Acc+0tZ6YXV1cfppHgQJkRUNgAzj
iv2+39nnD6rClQTvmCZM6btUqxHrxQKndMqCEnRpcV3RIuQ8fvHl5X2D35wbQ2uu
CTa6Td6mzwIcCPisjQAwCrgNr5AkUYfpFdbIU8bemK2p8uaF93UBu+F/gHy0vtKj
Hq112aLOZ02VmJARFLREsuk0xWubZywao2H40aRT4tVlSMC3zwvO5coVzCSDdkt8
QGJeY/oBy2rxfTV7VBahf6NnXagn+cFob+KdXJo/x59D3HHdhI8C0LtOBRkhzzLG
QWZm+XZa50Vo9BA/vbgcS6RLA3AojXZj3JSeE6Xp/Ytog4K+nzJ4oVafboOyw9WG
lnVuKJQ3pWR1/rheOEA+GWrBSGi6bITlfIOgjbBdf4PDxFpxr6R7u+0vneH522nB
URvBD56DQ8qopN3zZHfGcJRbjyRWQohPLWim2032W1mV9PMIU/grdiHqlveQSEXL
AZIDTRLS5WQbtn30phU7SJg9Drfwzwwo/kgvmJlQ9s6KBG3TggfcSpIeLke8JS26
aLV3UsCNc+cK0ItzL4BKapar6eWx7of9yNC2tV2a/kM28h+z89jPYe2tTDvGj06+
xgeCGE5wmdSNOacstJfm7IeBJ6nBn+yDS0SnQn3rb/tfYtybFhVIxKybccrvGSM9
K7v3Ra2u6EDENeLHXz9//PR8rm/0Y4MCq7YuutVnYYnyx1mKZSmtHOvcacqxP7pT
65D2pla0Oisw5l4Q3wQgh41dyshu3OKZmw0pPunet2S4u1dmaDDZivJ1bXNG3VLp
IeNaSwlqGh7EQ6TYuEA1FRvS7/X7ivIITGEEf9fynuLka2xP3zsZk0QsgqXtiX/z
74eJPB3XAZjn9w1HFU63cYnDSrgwtyU0085A5FET7P00XWL4ypj/1lHXcJ3t/iH1
uoiV2Clb1qto71QG+G+MpOxyHpFGApnKLeJQPetwYnvjpSWrYChacHxHt9i/ABgz
0qV/zKa2BWp+vFv6x6asloXZuCKKq26v3Ja+Sb0tnA6wr86qfoatcJr/Tlq1t42P
e7D1mycschKqXGXSSgJXuqjxIgZvUBopajLRQK/t6+ye08x4/G8ANT5WaGGajDRi
FNsfScF+N6BNQnTNtdFAM2NBOpRcWUKsXMvLD1YmXhtE0Dh/4S9GfKzZHewawT9l
0BylMGWBSBkjgq/EO13jxFL3I+WVHQc+v6yObmO26Qz/hnXlHHAoot+OVKe7LQQZ
CW30bSRrny6Z9NZAzr6ZiHl+uRK8WjqIFlm+shtBvbiNSRJ2zdkqpzZnrvklkOAm
aqsEQThZjk61/Tz3ovl8or4BFjPh6sm7Kw6+mLZvRuOjm8Y6dgMDeVz0y1Mk9BHB
P/dLVNqDidj7lIOpJnocz2wfKUBKtDSI+foUYsp5/HGhgWp+M4Y66NkLZ2xoIX4E
Y3sqv7kWRa1DAoSmtlUP7eb8teJdotZ2PnLov4GNZKN1lzrQxaNFpt8NRFmjy63O
6Pm3M6h57JrX/GZ4M5yJz3G7bw+A/2jEYZFnTBj5LtYJpCaDzgi5q4oTDl3H2/7N
9Dry9Bya/r+AvVO3CQ0sA2VXXYRzBPCsTimRGyp+nb6XztrQQCyY4lWZhoqhPEls
PRcTD2E9+QnqIakDZtj382KAzvdHwPzodzrucJXJbRDLgFPl+9sGe840VFynn5Ph
sXEGuqq1kKIqlGht2N3dRkJ8ifoRsFdsEX4t4kKfhFn3aMPeS+4e+bLUG9eATixz
0CWChSgI4c227ZKV/uEf8dRkxZ9FjPdWWtlFgjK3AihW8/kXWI1lnK281PVtN0cI
qd+EsVuBtxO/+hWqMMhWBRB6A13GGnyy5QBDLwSyXXhsI87+An15eIUyaRE/PdHw
cFhgM+X9LfXPNLhwhLfFBh1tO4bays3k8CaPppkalvs+NvtrMq8taqvnxaKqzlGM
RHRatDDlwhPmlSFLuxszg/CY60BRwg+urPMe3NettH8oV62roGTQvgXjShygbfI1
E0y8yQR7h5RwE670pTysA3llfb2juaLq4NFquz/swvlBItWDxLH0xXS/22N9V9Hn
jIlIwpFiMlkLS3QU+CLl9fNFoQ967dTp+PyaGrmnE870C4FtQmOEp/XGTiiXinaC
6yr1ZUcIwJfmGD6YpX9gNs1FAAJD1EcKZv1sNvINdB82zSBS0Jl7YSPoqqqf+ljr
uAXZkkYNbE7DnZTPDb6wVTVU+8y1FGr2U172qrjiqmgbmVANveR16F30FnznA316
mjiD8tuFzRzEEsdjtEg/bbdgN5YA7MH5JtbYW0/W8YOQhcopGIhu213E1afD8nNz
zPD29Oc4CtU0eUZdTW/d/eiCWzP5q8/gTWlSa/j3tFnyQme280TOE2MweJ5Tiw9K
3L9XW/VZCVs2EYBJmW31SaWK6kHuuOlrDU59vwhTr3TI49S0uSmTTVlttgo1szKT
3LKexd0mSHTYZVBae9snIG/7hNbUAP/RbhpsXvfiAPv4I3EVPrrTH8MHw1M5G3tU
PdwZLD0iJgsY+MQaHyVl3rVGjLVQtmi1/QemRGKwSjHR8GhXm0XS87R9OxMDu1zd
VnNcqkwvhHQc7d0EswFcG3T9vSIE+Zkw1EGfiiQJH3OUDGrtY7vcw2dyD4JvQymo
F+HfB9GeJhGpcck/V8qPAj7v+lj8zCiSS6LKdb9hrisoJCWF7V5QjVsEkpG9XmVK
ZkMkyf5cthPG0nHCDCBFGTIARx5f4duzHTTjOeSYO+EbrUO0bzxcNZkigJVjQ/pt
5DXW6GkHjoWCoRRskuMjYGhqaa54S0H/sQ5k2QkBNcixGL2+aTQJ5op/TU5iT+hd
dZ8YWxKUW9GKvF5d6j2i677usuhNwVzlBJL5qOGfvf6FUltzWObT5NmkWenDmzn5
yJVer4mS+7GZNnahx1VqJ+fL/KXrSOA3qoXKmmuw8FvcTJqKx5K0jhyDmklUZ1eQ
yHpxrVeOGW2HBu6makEfg8F0Nytrd+UKi/O/1un55/8HEM+6X7u+K4EzuNBZAgr6
FI+EU/XQUueCaRa9bI34+zfREhOhQUCXCxUnhJIhi4StyKHdeZxgriyR8KdvrnNF
4sVSM2i9pEC8UaFT3OG6QZE95zzHMpe+NOf2EvK/vAoIi0zKj+0mCvDGFPY69SWU
3XGQTbH95X8ulGD0tZoSmT2ppbzOSPGKjl++oqRZTbQ4+yEd4M09BID6JR3AJXG2
kvAhBevQpgFZhj/aEIyphOcp2Thujp5UgKkpmy7nNJa7QAYzRV+YwL6II8zS1sGr
vORYSb5U5QCo7WepXZVZIVKJApeuSd9iF+Qb5JFR0DP1VfEPIrAo3tM7l+SXm9lQ
s4cJScHz0T5AfdNz/guubdKJxVg8igtL2A60lNd+3+vFyXpa4p5j1GOgpr5jtBtk
96XWgLcRhz2zuTDpvftBckFXS9zeRVuk/P8gbWEOW0PCuYlNyvYlmAwUvTiWwNYp
I9rRKAwc8+6lKStyGbFNF2WB3ZI1pTphvggR7e9SYYFbpMc7lTJa+sVXsilzTut/
PJ37s93Ht2RoBMH+tEtNjfdu3NFCNW8zKE8Llvk8G/CyJVSufpsJsG29uP12dY59
JuSa9bMidH0VNtsrjLm55wAmYitDebd+P4/ApyWo3FmN0+Y/PP75qarsX7toFYJ+
xDo/Km0kEtTOoxH27blgbZi32zIEXP1yn7BU20VCTBx0eSywY5/tPpz6wI+h8swv
sjcORbogmb9usr9OmajQMl5IVWTPF8n23lXRdl83LmuCKo0Rwab7rYgXXa71il/+
L4aZrxYEm7+jgW3WKb8OKG+TzFumUER/rmi6/eCFhml9EV7vyd5zw2rQlOQG8TaY
xyAiyIo1V1Z1lt36DnwH8JZmOgv9LMGLa5fzvhc9nL8ZIDOT2uE7V6K7XKXor18x
uM0o0cxc2llNbdZxovQJ41i3yNeSAGw383qkGzsWZFTqlsPJEt8nh+tTT5lh4ATN
3brHb4hvbvboCN9Gzh0pKJDlNkPXUh+T0KSf9iV9hJ+IaWq95ooiwHugumVWOTeG
0u98L0PzU5qrFIlONPbRw1zHw8XW5JVcYAIKLV40GbH8XiW+glX1x4n3XUqLJl7Z
7jl2EJPfMRR95MCp7P5uds6LutV/rYO7+X3Ks0YFyXQfy2V/h8uia6HA+onI/QNv
v773cUdRcwC/UnJaT7dMOUgNaCagXeylBQo4OJYAFAzhAD5RKFHH0Oi22Yq68KkB
bto2D66VfkMg6QeP/clWyJIpfE3kXgazJY7lXLmfgFJI4d2FfKYDyiuso1mVIDY9
CsM31ercPd4j2u2pv0zvPyiCEfdVQEv2DMJqPMhBRLL7AeNIc7M6Y6eAcego1rmL
zhbYYd7jiM1qL9s61p36K8g0gJMsoqixtUTMOmMJ3t3m6CeDn0Ojski9f4aSYpqW
d2rXq9/FJ0p1+fypBfSgu8VzhQyfIx5moeT3YS/gZZnCaeRZJpJ2zvkLWK+Coa0q
3WhE+Dt3ae3QgDF6/3olFni0iiRiLqyCLW65XwWYoE96oGVJj26rz5AL0w8X6WI1
RAm+o4xfz78hbjwNZ5dlVbiGkRZiPlI38bHWHEqQ9n3vwgxxihrqWAR18Xc0E43h
2qvM5BoCofZdL9UusUcHFzjNaCchryPdZIGE2XGNquQxtWzrnPY+6cIKIDTYTgP/
nopJYL93+yW8yxjZd3R3DKG5UE21fJymnjs0s+Hw9I8KsF9HMxStPPgom2DW6tWA
ue/6sH/o03y63qnavol+iOKVu79pG/xmY+4WkZO1+8IHJ4hmyuTCOPgnAspmDarQ
dbwTX/EwPJGQr5LdZVea3izfNxLP09VyfzI+aYdPSSsZjdiAltw1UPLahwvHRWPV
JyTI8dlnXXpee+sOxx12rNVPaOMQIyYBZwqZG8GOqLW6EGyU3VZIrLOpAkVA8QJL
dKxNwPtJUP3egsB/gUzxDXMTqYvXLTUY0eiEgLfnTzLqNYW/wxWz8WU7/V//Sm1d
7jwe3X+nuiPiCQLIVHG/3rIotNjR03Ly9S4kw8xcHgoILgT7FG2/WOFlnQ3IdRVE
kR4nA1YKPV2UWatg+q+YwPUKKjBwbW2vpcSH02IvPEXhvLyM93sYRMpzgohHouem
GKyQR+pmDagO8WalCNBuEzMBJzXPGSm9pBJLMN3ola8/9Vq6YI3k0aAY2qinu8Ka
WN/gXHStbMDtxUejdMwQgTF54ZfZ0FHIPGYHfbB1nLpAjD2CMZkM56wNkkHZl/2t
tUkrds80LeFXS+S+yvmsrC7ehp/RiOZgeVaRnqdN41rFft+Mwyox4NFxyWHqbPiy
9GRQFpHJq+9TF3TxT82XHVyZwDeKjlgb7umMh/AEGEaTQFzEVyi1rkwjZCEMz0oG
ZWUCsVoAOsSkNolSpDJsgvGxd1CaMWo2bxo94YWIJz+zkdf0v+LB0boPtUE1HkZu
stkQ5Woh5zfcEC4xGBWQ+gqHZeK8/a/9HduW7sSuNosuynuvCt89d5dxf0WoVyiU
yWJlXnw0JTFXZuOBhRqOISdzTQUkwZ/Vlb90I7hnNeuzQ8XTLmXM7VY1GKXH8xXu
HLsvkhVSqBkbf+4Z2JT1tqVx3bsCL27aawCZG/VyVXEBmQ+Ct/B/sPeAk28Cyp/H
gCR5xLqiKSj+5vBDw7WDU575axZPS7OAnGY8XqG7YxTG+D7USj3FT1sh4ixbgQmH
ZDqQriFiaQwiu3i4hgq+I6Fv1db9nuMh7D2kTHNO9JVnCOp5IbMrGhBXpCBHTXDQ
/L4eGqIilMn+C9LEBGmOvgg6E/4Qazb0+72CBjydrris8OxDfQNsCjORLBWkxAD3
sgj355KtDEkHx9nlAVruzQ==
`protect END_PROTECTED
