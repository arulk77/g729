`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveBuX86lPeOdiS3NA6BxUCG13LE01sRLGnxeqGrqWAxVN
OIlL6B28Emrf1eeweX7ab6a9QGnQGVig0r06koE8UxvK+QJY2muL3fpLSxueqHRY
6T3dgskhHhzP7ID4b+qJxgB5qCL0rgE0ynSg1AWTlj0ZrlSsFArkjLOHuTlM4IB+
g3HutyBBlRTHd2N1we3fgFpxrOMwwl7Uvc+XWltFfzvGG/6JNRUpbB1t/+WdF2Mm
nSxqPV0lHvNf7gVhp34VpZQQDxngUmv/39I/Zje4vDt2km+SUo1VJ2d4uWTpL8bm
Xxa9JenwJVn+NalaHn5H2Q==
`protect END_PROTECTED
