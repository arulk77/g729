`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCJ3JOdAwTo86AhDlHttm3peQnIki21ciekSr27ClORu
gNMMibf86NMvBZwXoe0tkcyU0Cn4XN0Yl9JoFmxp7EkuqxttcEHaM0hAA9Vb5Ewr
m/9R8qHwwJsikPCc7mCAHVrhdp2KcIuPzgfJm9CmOwxqkiFV9NSPCDOuVX2XvNTR
UTQm+iYtN/Uma7HWrfLgmM9BvSRTvoIIPx0hQS+IAxZp2UEggWMl4Sriv15oANeg
AqVjMX7QJTEWKkkF371r8MePPIrIkdKpZ/obA1lXKVxsXMxf1Mw1guj3CJiJ0Yac
`protect END_PROTECTED
