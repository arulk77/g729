`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKqzPUE0c9Y6vIbpcZp3NOZ9OVBVWQl+mLaZt3y1nJG+
CyAJnu0CH1pAf79Bl6SKyGUNDPrcAb+IMxqyJsd/vLaenYD+zlUiHRB5zgxl3Cqc
tyCAIlNHN1k2Vd/Rj52IQ6NXGkIuSYXhu4d3mTr4aawVsktkdV3FhrWaDrncPyc0
51CZWwoTjIhnaPyt6sYNOArXHEBMiaq6SPwunZOr+6r0eqxmR3mxO2OORj8/Ye/1
KYfb/2HurRnkMPZivX3p7I/A7uhm3BpbiAcPSjXvHm3eesHp2sUJfCO6A7APnpIr
bKw4jHbL2q1lg2K74Tb0hyr+WRl8pTK3EAu2MdQJ/FekjGs4WbtXWIV0BB/mcKp4
DAw5ekvBYGAweuPyf4OPZk1sIoxn8BwOx6b4YvgX/COeoW5LJAkAwMhzZ9p1mKkg
Hhy4zII0DZ2qONJ3qIVLWyT4KPSoUk6X9Kuo/r2xTzMIB81+i/PBukeIcHGBzwre
YzsbZ85inUEUIoBm84cxEnQdlBPbPjkuNytWXaKx3pmEZ2B3yCpyKGPuhnseoI9H
`protect END_PROTECTED
