`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
F/7oOJp0h1doli0piqOjVEUiu/GvP8LUMRZZyhhBu4c2F0GyYgbh+qRxeekucb9V
oHbiXZi1mql7i0tqW/j4El7CBQnOyXmoOyh2/B3g3I/3c/afWGcEePDWlMG2fSqb
XJWL+uPP5tZvJ5lAQhkIR/zjShtT4FFvFUp1w92nWEwvK8QGFNqxEsqedgt+j8NY
BOyc1PcZCJF7CJzPKOlXgMv7jMMLwyHTpq5A4xd60wo0fEgNZUN6KdUq8etrZTEt
fGBt2gthrbQ9JD7gwxHAZrs02C2h/XJzchdORzM7Qx3Vbrhf6CuSjyk8kCLSzGlZ
jSahwFvIAptktrPhD8lFg4VTjI14gq8zvHQxq/0Zy03yc4nX+4YGlpDjYG9TslTP
f4N5OgO8RB8EwZSrFEMreL+bia5bTU+mK6YSvxNHB61Aqmx+Q4aKIxx+HgxI56yF
VWHBPuALfu3mPO7pO6a4y936zopsOuLkwZJXdREjP4IaemFJG1II1Gubc1CSgzBP
gXKx6Z5isDIaFg2qL6hUoFQoF7WaHR+BPZudlD8LtMQlXMTxBl5YhE+LfKyRqlS2
tnSr4hqdjjMS7qAIUaPwpA==
`protect END_PROTECTED
