`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCtaKwishvAepQz/ppoDCwdHpPd2LC4s+Iw8OK7AABTX
P3IqEzwp3UJPpdQDr8S4oHtKSt/EY+MDVTC2LzA2bF4XzwTgzXuCGyjrnDeOHTB0
x+0oIcLD2985bSEXd7c/bjZFwM+u0We5yDgAh+7uBTuKvh6MSyo4SIsO4V3nqIXQ
ix51Wapq761eYFK6NOUumjOa8ZLW/hTWzC43ZBGtHV0MIvfQzdt2owYh/A/VJ6D/
OQIGovsQHmsR2i/Gfe2HaT6bavZN5KI/cpqWgWN7yM+3uxwktFC3gqxWwxIO5zJT
vxWZgmPkAi425NwCszwOy44dJMFNufuWXoWuaG3fbezU4fE6CDuhj/B16iz3E08g
TBW8tIo/JkAnFDKx2P1Fnw==
`protect END_PROTECTED
