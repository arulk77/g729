`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1abW3g7ZO0TrgIHP18h9j6WfPmCE7zUblOmNVzEwM1/dP
skoaT1mN/ycUbC6jDy3A4lrXyXl3+mm0PbEwVvtOe4P9hRHoBfL6XhrS5GTN/xXV
e2WJ5zKzrPUqehgx+GM16pEBmLg49IHNDTVtHKH7xFGoevpQE/QLHxESFpVe0POe
4AK0DPvrMFMFxyL7tEOOb6x0yqVfExIwc7hFH9TvDq7B77HkvhbiVdNsrud2D+Pa
rllmNJakz7kHLiRTE37jf11IcFAsrmzNYChzl/IBVT8Fbk/QnnEe0SecAGD7RbyE
D6WNajI3D6c/tcJ/Acodf67Z6COW2ARzE0brr6bYpJDSnA84BVkvo6jlaZLEGyPj
lEP27e5vROOUeU0RV1ghTR+9Ec3B4Fcd9gL1SIRWcH2FoiT9Jyyd5P2PVBhPtw02
ss+6vUK62O1oYWCn5eWFXFdb6g+yYySB/Xc9cIYcgiP7Aa3n0c673qfVeyXu3ZI/
Xb56x1zwIkP0Fl+Xwjdj/8nZqzjFCSA86jmJ4cDfTD4QTtSPUxUYSzxwM+9qdJzy
5b/MpKscity85wvr/fIGs8eUrWuqChVCJr9qyqrbBpk=
`protect END_PROTECTED
