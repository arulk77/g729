`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL86r7WpwgC05UOGErcgulYAcmpOUOCJCI5aLX9g+CKVAK
l61/yIjUk97dGqbwdPfjrKqWtLWjR6iz/z7BGj2zd7byKBs/ySvZMHEeJqa+K5nB
IXUCJsWhLQckalGyYk2kiJ8W3TKd3hnomiEaAVbEj2YeMUYIoo+pyTm/xZk3u/0y
F3V2fk+tdvdLmY/3UtcRY1RJZ6isW1GBysM49kNVYhF0Jik0Rqx9gJJLnJyiNHX5
u5aP0j7Pyh97kH+Lv16QSIvgAw08ipwEkyto27HMGd/kkqZsNKa0LWA6QM0t+g5X
qfLwRoL6y5ukjKwnZTvCRlkhGgV/G2cXFVJskzufWDY=
`protect END_PROTECTED
