`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveF6Kx/2+WsadgoO9GxcsFhAkZISJjKjsV+othGxXwUHW
9VXLG4OrxSM+a7CHQJgOg8vY/XyccO7pxj6wZf5Mp8fnzbjgPTaN7dZmrC5Atyum
7IUlRQ95q2YxyFK463q9BS3PASvCw9OtGp2GFYXDlckhOPNeFAPDgvtDufRoYujx
oGvyMp7C74EPZ1UbjbJkhDIN3/+lDOzGEfLzSZvoTb16m+Z6JV3T5/zAK53p2Kgw
kzXgdnsBZuzpUaVZhFKekV9e+ZQ6MXQiGVUiJPQ3e6FUjuKFjd2kklV4ALA/Uaii
C/8nW9KmODjCJp5OnS1eIUjJmRdCeZX6MJGePhkbKkqkF4uKvco17qzO9gNCUtCI
mZPzaprwWpw24iqC/tM0L1vDiBdK3ktpR/oSYDXUZUNwNvV5pzHi5szeLWvOrDog
T6yLoFDPyyxAvkJmUXhEQ6yRcideicTHZFKBKJe1M8RtEYrsKhmKph+V/T9hCgVC
LwJ3qx/dd2kjSsXTY5IXA1LcuPtaARuUF4z2v2DXVuBj+QQdawahkBGIhQycrYwQ
DsRigoc4Z6X7Fj3Vr/sWicdxIv30ohp+rb7jaNPYiCGsxEbHGQWytPZc0vJOBf2S
ga2IF/JqoC+ot+Q6k8RqgZh99TANb1Zg9HfDbrgvr651cx1EYykuGAOwBO2nl4Vd
GNAMgOYGQPG+jRcLztuxGtc+43JAFNpPsxy0r7s3x8pqe9MHPpddJirrCmy8ZV1S
ewVNdiaGlDDxKH82Sbt7BFVOAhDeeciagDxjMm81ZdLyem5YMSvL2qpeDW005C3B
RU/zehFk6LX8Lr/gD6NuUuAsi13qDdX5krK23f/ySEYCwD7qLQ0m4SaCf6btn/aP
F5QIX1Pyj9OD+CxOh17487HAsGT518TCKxE+oF58M8Kk93n7POSZYPX3mPUAJPnY
uQt3L8/zpe5+6cfnuW1KMw7V34NDCACAuOIICpER3EauX/58/UGCjxo0Rpz/DNgT
X5yaoV3Lhk4q6EIb9wfgv6PpOla1xUCuQEe9ew32J5QhVsr9URoQdxmrZ+iqWUIj
FWFZUhixMDby/9iiE8FB3bxZnI8D1tphNqyA4ByJrYxKLDGxxAS0ZnMUho1Ft7v2
+g3Ze34I7G2JG8OvS6X6bQB4uGan2sVPZZLH9GNz/nAyN7GSJqDUgVFjdwJwZSiE
yLQx9yEWO3obnPtE2twNg4EoUKs8fbiMVchPfHU8RiHYCXId5rvvfJSJTN759Wua
gnLqxr09SzdbBry6hRidYgBdOY1YPMjldh5OKME9EZ1oScfVaYiuhnn3ePoVKVkv
Em7XelVzwOP+RyKdgClkg+3/Q8KfneP4yNaRKJi4pSlci49FPtWJP40KP9N2wTNc
mL4I1AK8Hhjk+j0t9bT+8RYZwgz+fS0j/cXHsuKqc4fsIaDlQ5I5i8D0IAG4TyN/
KxpBK6JLQZwn/JKRrIJJS7/3xHQA/uyfSyijvBxxwgdpe1fwWmuzrNfUYBzyTtpD
oHMT9Uk+LMP+MTxwRbWDjy/lK8de6NpGFZgmZYu4Y0w2/oxfzwYLrUaAKB2DzVbv
+1cKVxIaoNaiwCIgDb3xuOB6f09diMZAAUPeRjC0b1sx9aeR5lRnUwlk76IxwAU5
22loVwjqLPvK8BBc0YhP4bbwvszL39IwS95h8V56hXjEb9Mq3Wp5cFu/jw1W+eTn
lilH90AFXWBOU6GtAT5vtzNPVYrLPQgW5VJnrkBSWuun33vU3XkrysODcfT2GwzB
diW01uBKaThImi6l9fTw4EB8atXIOt6yS0nNENz3NQmkn+TQWyLRqyx79F0WNGBU
4TGyRdCv0pgaTSvf2WkhvwJRVFpQR3Vf4YQif7FQ3GnjZ6U2SwzTSN9c63HP8IGh
dFxZpRze6kDxbmLBqeo5H3GlE/STH+n4o8JN0eh1+4/CSZ5C7K6ADIRsGE1WgSMb
7hk9rDFq75euCk8mTDvPUrmkxd5cnYWDIwia4U8hAepOFuJ8ugb8lqmANU5yMywN
lxeggn6PQLoOHSNao2SALOPw+uvUNy8F/IU/IGyMiI9KLiI3XHGGnA3SFY3zTi2D
XXiwKOkFUF/dtO/qfCz26D2yGrDX+uwJbRUIzfZb+K+xxsFllsMGO5EuM48t2UzW
/+OU/EQEes/2NnDKaTM7vPPfIBZthrD8SKrwtXwY3eKFR9jtuuH0STmtMxZzPDYY
sminZcv+zh9x5vokYtUIv1L7eiP4kwcpPomJkuWnJ/EIVTOgMmTruC3yYhcjBhlJ
xoLYykC6pPTAD+jE8zsTRSRsm+nzynAhtBNm3qZJkTd5lhF2dTznScOmuF1p8btD
bxZJhzNdC/FDZi6XlSITL9nf7RL9UN9keEqriA+V7yyX1YkxJOtFzR0XhX9TkkLR
mNZbwlsK1eICOyY3yP/uHhbU5LeDPD3O7oZY9PZi1GJIOqBIrELzJhbRykkUEplH
YH7lti22QkYwqlPIbDqYcuiQu8hgVBlvqj94mQCKqOsjCqHW5nSRuHvLtkLSHfWL
KWEHW1WZYqTR633zwuIUkrz0Me3N/GYOwyJRB7XhVV5l37OZ6mr1He0gplm/3WDG
RaRzqaokIEHmMv8FtAwX7h4MpjSGRMHcOTkD4daM47y10Xt70666FKy2qZ1LAgzW
S364ykeYsS2WloEpC23yTcAHRxH1ySMI1LhUps/IPWRhAx0Ze+/yY+y34ixC9jAA
HYr7C2LmCdg4ZK8gnKlIx5Yf3Iz6OQTeyCOeJJ+MbQ2jgYT4gBnL1jZwi5XydYDE
CCSsUXFaDUbZ7lOzKsw4+YRLXzqAElJ1eQfAzMsjViApXajNQv7PHyLcYT9qLwtY
8ANnWd3uoiOy6AsLoTzqx58+PRArqy4mGo7NEVFbtnhYt+1+5j3HRP9ksQUsbglo
rrem8jSO3CYB5cSryayrmlPqpIpWgSVBj+y4lOJJfMp3/6CSiMR5Onp4hPyhn41n
0HMrzzdcyCrtAsmd0HRZddlOfWNJ2Je/wYOw+VeIVJuSYs0ryspzE9y0xcfDBYQL
iuavxeAhxeVvUms7RADof6f9hhNjsuTOspIXW5Yw3rkim7pmNTyolfmvzOogBWnK
t+ibKzGt5WWD4eTIrKH9i1+5XmwYiDV+527nwqpqU7Zpskq2dtdXzRzFZoW1ijb1
ew8MQ7Cp8rQCoxAqMDONj2j8JBPChRyAK2XSjFJ7Dc5jr8wM6MCz3/LhBAr7m8Ah
UfGHcWSOkkyh47Rd3o4h5jUCu1KrUil2UlJjJbyWsMHVX2ofkpy2Xz8Uwhar0FDL
AwqOF5xWM2bNKYmyAvStGTlkQZrQpP6u7lYLNfsztj74f7C/ZBH23bTlVQzxrJg+
0wIa+4BYuW/5uhobTAQ7dlK8X+9uD5i4Ru4BTqk+KasILfm8z1VDJs+rJz2oepU5
Xb2FNhC/3k2iHUHJj/j/7nZ+ZRlVg7+j+h/s+w2Hnt3KV79sR6biLxyvYdnx52+a
su1DwJVypr7QxiGOLcYJ7P03l1TgbsVYc14cP7FdtiZgGb7DtTGmOG6LVqkCbYxW
LuZOyhShdV5TxS6quapiZ1Rrgi/lFGyTGCFkHcmGYEMESR5Qbbawi3g/BqQ0LA2N
269Tii50f9aLVC3u9W95H6jQcryhFwFXEs4gQT+4ZCsAKAREtJH5YXRufTJZ7/pt
bILvK9+Fi9CSz8SE/3hZNoBk1husFj7ZOXTzURFproa6tF549PJLgw5CQLq5nWl9
xsb6sqfucEQpUgCCwXxhsqq7zYAIn+sxrvUULZV857DZkvIoOvo7iMHxss03EAU+
cejx3n31fFzbgRFi8rv4K5ErDdd7w7ferTfuBfMwNFBMutOMcmbeXFgmbXHmwkGp
y5xuHQqVjwXSjsKD84sKBRvg3ARLbY8xrp+2SWOz2Fw28AjxarqQgsCmymVvjkcl
RShCce5QEeaD0DaBrzR3WXRnNm6MU8ZP+zmKtuQtCiWwJbgOMYI34yFbQTV7qeYj
9rvkuOLn0yqVqVoek+xeSme9pMNoGF2yh2lp/TGNmNXL9+RziycXhC29QMA2AAjO
Wf0iZrDCZ42j1TVcoLqt3gcbFwZb/E4rcKKzKeCdwk4x+IJFuPmYOg6g2IOUpBFC
JhDIiOi0LQxTu2CiU6m7/t8aB8cXTJmt3EcK2L9sOD5N7+93bnVLWNcD4FBjYpGL
Wx7vxLGuXe/xg6SUP1BOH6a/1HN2UwpfYS7PeEMP4VNcpfu4urQPEz77etQmT9xK
togIJMb4oP6pLy10Y5jta62Oxu43+gaTMsJ3ovuHP/gmzc3asXlEmmvV3NnfCic+
9khhh7rPzDb1jC2y73UeyF9lI8jMQRxIPnZPbCsLk1+OWlt+gQfIj8e0a0ztZfSp
za7WNSiMjaHzxK1B9GvvzmpGbQJOX3fC6RU0lnf/SsEqHnLB29v770RNnacQkU0p
jMQx0vcFx6Bs++w2ds1/byfyTcbCTtP/CKPONW/NfmpuwZUVEwsp1QX5Ib9p1eeU
Y9Fb+m8Szd3TKSxSoIgALBn/Mtq9F93BVQ50uT5yw1j0HbMuK89r1/6p9zvLzJol
ET8ch/9QmF2lnutOdscH9AaG9Zim1BHGkNWeZ/kZ4g3rsXv8R1jp8mongmsiXysl
CplnHjHjfKGIBzHCGp5kM3UNNnIGzsbQiHmhFSeLzBJNnaCRohBNZSxjNGotjxFX
i75Mpxs8Yml0GY0nReQ0RxNJRXi2xCTeCgvHMnGlifmrwFDIPqP3K2k8ifI8UYYi
peS2tiaPXcAfz4+IJkoEBOHdamttubntBxTZmVIIQrTeHh52eNf7DFgUtEqpm8wa
h0Iv4qLqxBy4mvW3uSwDUTUUlHcInV2bZoSZxeuAuQp0ru750oOmXew4pL6pStye
Z/yNrmxwNp9Z1zj4M5K6tDaHdG8A/oty3ppRokPx2ABisdzkbja5GpwUNET9VQ8i
VsrM9ySRQJranob2OCMflg6ON15wNblOM/+4RBkuhO8H3gVdBfLi7lJl2K5lKU27
DxzwT5ds9o5KKCWQglelctSqVPfVM/1fRowOaxEtOAeRDN70oWyhd6WbnFoGf6P8
1XxNKqMzufwOEL5GTorFVikgrpf/uFi9qqhwoMXwQzKpbLkgJueBcJ1GLUQuhI1c
gFACa7u35qTdurjmyKrTslvPLow1ppEkIoynACG48kcO7gKjdNceU9cwU8aC3d/+
QDelNtI+V0Ud1HvOw7CJgwcOOSV7c/mj+V43NiGsil0lklB8FtAuZqGy1RWasBn1
8NPmxY0LoV6CsXNZQTIO/riVM6DepIRWjQXwhgOV/weF1uSOCCWTyIySafwnOkM9
vWjgpZI/pe0QgdsuNrV2WslFb+73HcDLSKQmy5iYcjsZ5m8SWV5A2GcST5VBcaHf
xPFN+4R0ax7f3VCCzmPktOZhvUVfq/9e7sTkNL7T/CvgfIE6FfOYRV/Ky3uoXEKb
2rCvjkPfUd1VM+aq69l0oUVRG8pk3PH1WT4pQ9tLtOjxJSznUyM4cmXuFsKibm+n
grSwZA1Mn7FIO0cp0TcvOaNYO0HtyzoCzpgUJFMjXVEWs8y32xfnWXL96syPdXDV
xS/Fd/3ZiDCLe0XoX2gVKpagilk30lwBlzj9RTzNkf4pi5c43gA/vzxVlyfAX4qx
lrHzHPkBR5eH42xqAIpXfDqNXgohclUC2ra0YVvITx7bwPsNwlo+ZLkt6pHJctSU
dEfJ2jQnovnzvfIniMTVbJo+kKuv937f2+B7eHxa2X/BdpvgmKIlZtlhxXqA5qcw
KHgJdY2uaxsUoy8rE+L/cH/+8PStP1Zysx4tOuMMaP36cdWHxZ8hjPC0GKJfeaeR
9jQjeTw7MGy44EBzDfROgL1HCdJCpWpt7Khrf8mxw1IS1ve2oP0EdmfTZd7v24y9
9X39+CZBNxnO8zemiLwPS/oYj+qfEIIKtPOUbDgBIsZTmqnPnrgr1I84KaWD097M
LxVEzlC0VX+0aRP8jXyXI06u9/MFSu5nPWyU2hczuX9WVvQxAFTPjdNq/oopgYeC
MkYisvT9eEvVw97HNz4zy48ui++DLFA9Ic8KE4Myndr47cMcLwHsSimFB60eoovV
3ty3YejwC29YVPCnCecMCc0Y8MIN03PtwfirhoNRBHq+EMr1eLm0UUXgbLH88Soj
i2xDKMuh38YHgIWoMPoC8z62m9Kn1UShS20OtgSUBoBwkk+M73fHCYPAVZz0R9mz
wXlR62ZUgrXKjFHOBLlcV0Jj1nO8LGFnmaeCjtV3ual3qfQeFB7kXsUuD8uI8Lzq
j/un8DLFkv/BrkLvtne1KmHbR2TSnN7XRBFZVHs7XPpdk32q14eZfsKplmoHLBV/
szz5PJb8HuykRD8hgtjmiZJ6qcCV3kx5nspTXwiK0cLTLk7byuKr1n2uLotEW0iJ
lmNKab/WWac47R6rZVXbuwAeuYFGu8Zk+3wB5QjqI18M5rSLTBO6wzhlFSPYoObE
jXps/4RtKTotuN2d4EBoyilmy8asuth7FyZjFiAmL42KLgGPMSrJ4oHOLIUzMWvc
lK3gsshG5aF+K6TIfEOl4/gtyrzhU3V7mriZZxy8tNxiy5DcBwHn5QO5LzSz1ww4
D1ryKO4hwV6gZmyhmJqO7G54oT+pauvsII6fyPsEYtL/kuncfmOYxOrQwc3pM1DI
dtwK6ztfYXqwN5Dk1Js4uBrp+7om1JdPf9jCbF8afahc4pYkekkFD8KzPNwcYh5v
FHxiHNph7rHKlbiDjKxTB0OLKAkaguUWdD4gMBnyqLLxET7bAqYX66ALWjz2v6ed
j7Sibw2knsQlYV/WxJiBXUJJecWIC65LoVJur/IR5USNEp2yG6a263own/M/EST0
NawyFGBOwQzxBUZUh+Se3qDIwgxdeYIAtH2+s73uW1k/DaV2vQOCU6Sc4ROXwdpy
WEtV8Gg8QN7VxV3OSOxaDHdxXvb6nnHy61GJWcWmCf7g2w2oa6Ve3cwCVVosYvWO
NtxK+GIL8eFxMYS4NZJmSlwJ+8lwjMLV7ya336/rdM9kcJrgp0NaeKJ0C0PaLzrj
KY4X5fr98USrFG9CZ/ahbNZVWlp8ajop9p8Lvx/aFkSnoo94Fvw4n/WrOUPvFM/J
AIC88LmW5Q9ETRcOSsBT23axvU3IrPVzX46/HC7GG2L63suN2aO9pbx0S9cuqgPd
EcwnBeDmo6mk5KpYFh7+OaxPTKtH+WYyAcP2UKt0vFLEsWH5h5EUiFCxk/gtrJyI
kFUX5XDbQbZhZc7+ETKgMXbJY2nj1dhBQ0c4SwCHnZ25U/EcN2dPcUorNk0cyG9J
vGljIrX2qBh3xh2x2SSlVjgeSjLcCW1syrZoZkszUJFodgcgbjszk8yx5jv1Pufi
0u4mv06vjN1YcJQbgjcSzvfE5Hu1t9EBnRrnamT/nbxk9O6VmNC29vg/qANN12S/
47qpxKeRiHZNrgNZgyFSVP5uLQferHYIo4F1Ur/+EFI6x7ocOeAPTR/bHwvkaH+v
Nmj+DVOkvOdlsbrv07lPsCLjaX10ldRjUA2pufoi94F0dWAdXPBa8SqOUSOPmDQJ
k64zRcvDtZ3Lm4hWzTItHDPtTbwZV2RayT37R5PUxu0X0o5HW4X8aaDt9GAiPsDZ
+ZCmCax+8AL1DmNCMphrK5QXJarABJA9oSs8gtoVw9un6smNDwLCbT8x4E/W2Cf1
QW6t6gDnS6o8G8UUUMEJUmutN0YoLs3AtOgklOn+0yYTAmx7Z7pd5xfmFzxowNnw
YcIcfxY0Idjvlcwo/SZFib8cI4HsYjBZUGuPdoicqU4nU/gLiJ4bkCJIU2ZsWKuO
jg4+iPj7GDkE/U4X0mQng3nsvxFhdsWnoJp2CFxWCG6v7oDq/MIjQF7DhsFhhgM1
Y6GJ0/udsTiLNBvlio2Lps1ADvcWBPMMfE69Dd7EcvGyRrnVgPFDlYsb4k2Gh3Yn
eK271FWODiJLIqgDBbIDPczopgK2en5tnLiKvIgaP1xPWzyMgABeJJk7w0QIoT6Y
xtB/97YOcaYayrqVpnJ32qpEteWu5gl0gGklzmESmQC7r8Qj4/bOPftlIpLct3vs
T4NCljcF5SyoJOX9TokdyyrSULMEKcoeoX6DgcqfxzADAfb3yxbBputS9+6tK8ay
oj6L5qEi7pBqAPfZBAPGwAUpgxj04MFaszTUbarh9214Mx+oXkUkM4p0HOQ8I1Wt
nqTNRE4enqZAQAJmVumr6scfnZ6AfKQ89ZI5De9is2LhIqdjhXo/sdFeq3tAMeOn
xDpkhCqDgVAECV0DF+KivGkuHYEhONspLkh6AQjzt+fMlPlN3jeiGPw9BMx6Uau8
GMSY/MfDJRAPC4vOJEZLum5i6TkHpXlSlGfQ0LJkaF8x4+ZFmv5IOBiZkjQwXtsm
yBmx1blT1R+Mvb7HjiO8FQ2j0nYLq3HvK5ptfO1sCEPbjp0uh6YXBsmyc886kHeq
7w3YG7YdFqf4lsFTu1+1dLZCluTT7jc0kUAZ8JKeAUauaEZgme3h7doF7xK5suka
J54AVo400hHvB8sHofqcBW/0krz8viQ4eWostGR9fATAxCaIyXumGrZnSXTwjpUD
kLFPKhqQlIfk3OQAuCJBi8ehRJOgHAMcwl8Bew4RL8R+fYJ95Bo3Rp5XRAn6IMtZ
GqY2PNM419jIyvJ6ap/lzj+U8xHy0rfHJUrqz4SRhlr7+xlmT7lILKZ91+d4QB7L
ASv0J+LVshva/qhgvkCdoP1M3BU11b+7uoy5rxjXi65ZCpVR2o+SksaSmojFfHk7
MC8rx8/MnbZ8rMGb+ZHy1esh20LzhZo81gRIrSnTTwjm2C0BypwABnLcHEgb9aJE
DraaU36oFBdGWRyTg+mxwtwKGqYLZF5axxp8ygeivsgQ1bhpSh/uX+vErfy542qb
3I1RokYZf39+t7RoQj5HBVCx0ZE4lujL4pmGqcu/YeSErurhwdTwrbG4WFHWcUV0
/QgMGkPw5aVmBrGdUhFAJ/uSoo8IgPdrjlOho0DEJgboOVvmjfbh8nGhwBGLMUHD
dBfd0g4UroJhXN5leqR4KfGsbKv9xKvwJam7+UXZgiEMdQAXXoAS9JXHcNbw1NHW
Q1fsGtaOt2g7UCQtLFdTmi6WAdvMktol0vQafxjvrRimQOEnvJR9C+1qgYHZXnYS
oV8D8CDrexI+obPkgkVxdkmVmSKBKzIc3ICHPsmq2jZOhqqSGXuKFBOZxE3n30Na
5nGcYc3An1RzIEvK7Ywgmi3UgpqOZsLnUKMBNHbvunFrA4/2+VSkPUidVLA+BNcY
3Cag52m2qyfZ+X3le7akZaJflUCjnLpH7bOGdneJQj8vHAY67PPa/nH5Njwx06em
9WGtONrWMVPjteigaq1d+YgBe4sVdgms7kpqSSAVM+K87APzIELYDVOQLfdi7ZIo
sK1miRdeTTdn0Je+rmP4D/FharPnCkY0lVd8MReobfSC80p3BgWm+dvKtJA3ZZ6x
Z46FlTaejEONRo7R4wy80a0bCDt4EC+uG/v0XOSdjeLihNgEacOy+3SCIjOrp1Bn
3d2SkZY9XsSiQPkM8PfEHvjTu2OHShAjvumkYCgNRYWv0oQkGY6izXJjjBTRdTy7
4U8Jk8IqX48rm4hnEmKDepeyVdRdb+7+WxRq006XjkjyIftaOBKSIit2bJtPx6gN
Sp6dsG790pvHycbALgnPXt0+0bgBx9ofI6hwiN2WEugo4CSnoknXitpee/LR3YkJ
TQdXJXKky1HoyzHzyWZVUMnlk5VlJkFxzWF1Wai54ofVJhivSICEB1ryjx932SX6
ZDBaxlCDcSvH+Sg+bjj4tchtdVd+rXZ3D7oJWfOur4slJX10vSagOYK09yftPEoE
g5EkGa1ThnryrvS6uQ3PTlbebPMXbANzcsX7+g3ijWrocU61Ur0UlN1PGWDAaPp+
+om+R3EgyD5h9d4U7HuLcf0rk07DY2NYtPvsoAFXl3Y5B1SsLmFS9JosfP5aaqcl
K3OjiyTCpH9WsUWD+kW3GaOy5K8Tp7AxecvZylxx/oReQZZOI0e507NbDsqj6Ymn
WCTmxw0wCVTlEk0v+nEuw4Rf+fgdCB7lukJZJJoMF2xe3Q0FGu2VcyzV/TXkU74x
G8dnULEush0rt1Vod1LMzXkl/06WShdsP72r7MeTiXtqqxlXdWkps1vXZlTrWvRY
X5lkdJPZH3x28i2sXkaLRFbWOPGUXzS77hJ6QWMIiBBdTOe+ZzenW9NAeannmtd2
JO/5AC42keAZC06JApTTCzzrrof1sBP1F8gNacUrD8e745d77nKNY+RS3YM445+u
fGVuvi1IvSEpJLiAtwCgzngs/EiAbQCl8e44Yf3QsvCRa7p+C1VC7ZwuL92qg5NI
82Lc+1SltbwX4VwqbNbT62tb7pyuEyGEQz7PAZEppg3yozeepnDNObOjizBOjus3
ZHMyEFMfvzHqGUoCPJoYxQ4r370WiKMq9r+05dBfpB/MRWj1ISaQPa0/8UT4NBok
Bc4IqVoBZORHMEVfFWi4sih30FtRjEQVBAMNZlsoAL3dp0GxArS9gOxYjWnhnqqk
XzYULHL/7njIAkCspCrdr3Zm8/9pVQtRlpWFmFDvDw1fVKa6x99tWmok4bOGTORt
Lhut4LisA5lcxiRZ+b2Hrg+xMCPqEWshtdg8NoWQDoHy1oCHhyks4RQopESKP3yV
WXnmJmE4ItGC7kwuHyGfSmErYGdJXaE8xX6iSY9+XUz+muW6spMFtlaoNv8nVt+s
271uhFlFsG0XfCRpoDyan9cw8zMRWjfSZmqrgt+1kI3rS4gNuqNSTRvsYgnfjwv6
Z98n0e0MCwClsEPkBpVcQvjjvOLpCCQzKIIrXm/CsrLI7XtXaLIRuDPIBt5pQdEC
OJFmlcZjXLUjUAONnE6cdiQyp1cLSed7qmX/IxMC3yhWRvbQQ6Q61ni2bUOTr6Sm
5hnP8xt5Dag9XYdopJXUl+L093s/OA3Ntx4H0hGThb4clhVqqSvE/ytVJGPctdBE
SzbAid5M1fqFAHOCljGIZdcyG7hCekf2ThX9oi/wrhhYQajruS8rFBdVxynh75C3
C2mAdTKYB+E7xOPHutE1XWgFcB1IczZpNUiA/Q1n4lx3M270BkcgCIu5aaG4eljM
vUOxxbAdotm75O/tKZaFE5Hw6kiuDUP3KBUC/dcKWXNUpVpC38Ij34BWYEmbIVGQ
hAjsVfJ9B0T99j5LE1WinyTATueUugOGkUXHXbO1IjjrQBMQgDfXEIv30a7t5NJ/
AsCfpXSCM8stxrIXyUcvW1A1Aoippcg34fk3uBmjQJh+ge3HBK5/SA0Xg/ojl7cq
vAcPxy0CAy2NQjxCOU1FUWM8s0njwqBayU/sP0qmCqNN8kkZjvNDzhWuCJjy6Yr1
79HLlwTwZvy2a4KDMCbMpjrngy+8vD90ZjwUwdJQ2kQMkdOeZWSR3AQ+ysrGd7To
aH6luGYjfxZfaAJN6B9i4RpM5hDZ/H/K38IMbgNdeB3JsmmJyzJx6SRPSd1R9nUT
Rf6yz+fRCWQH4dG3RmlCXqVlfE0Lf/PnWf46dqL0UHlLvFlrdDA1P6UKOZAjN61e
tc5oluc5c3BOp10wx9t/0PP7xBRxfXx+hNQlDiob75yVJuA2c66PhOE/tP09wBHG
pa9wq8D0YhL3XII5qxdD7J1xD4VqiMnBjWY7F5Puhp/1BO40WnJjSYdOt+dcqxHc
ZqPDSFpJtLjGoMWD5rshGTBvFZVfK6mkLHA5I/LM4444p74j14WE2+YQb2OtTBAW
s/fygbo64hTzNfnDSTSh1EmS3YzZvr7sIt9UURLVcCA6aFRIST8ljP+UUolORagt
2Zsxn06GBHzWTMBEgIDrbvmHXPFoOecl6ch9UHtufaZS82STLcNAtWYJ8AdbsH1c
/dO/7pzsWNrQ7LueXQslqxlu3NMPOGhsm7HSNOYXgorXirgQK3NInL3QeQHy/kQi
HNvSLEQ7RvYVx3ph7wj60PineWdbNDgLReNpAmb0Zcv2YTBm9i+jnb8Yqve9Gs0u
`protect END_PROTECTED
