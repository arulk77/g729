`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGZF85Se4WfxbC3lOQ53uK5mAYlgRX9P2lC84cfVHbZ+
gSvfbTlP/PioOGGy63qIB0FhRNFLyNMMo/h9ijdCan2sWAjN2fUcz8yQwRZp9g9d
bJEX7st0AZ0rcoGladIlghhktJYkZg/WeK1pczF5YcJzywOQiVriZ6/PYYZY3aTm
whpb+9oLCWxObzjPMZR99Xw4xqDy2M2WluS1lidNpy4Vn3L8IKX0U7lizLjjgE/R
gpsOYZ1eGJ1AUofCsA8Z9k12CcsiempuPJHTg+LFkvu+TWxlc46yIkBcSb35w4dv
2HksQ+FGLKijkCtpDjr6BkqGV2OJZk33Uz0M7Uolt5ozZT7fEjpd0O51i4jpOCWc
`protect END_PROTECTED
