`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C82wvLOeNse+sv6qS68OZBD3C9D4qORvenhl4TX9Ttdz
ykKwGIRX21U8oUTy6LLQU1TKp0m9ENulOj/ggWlL7/Fgsq2zAhlDWdl14+kivSLn
D0kk3GnVk1ZtsSBKEWPeb5H+mFw5KqEE/C2Co2GTCvc6QD3FAmHggDNXSQw8TqQh
BQLDx4LQv63SCed7sLEZc3b3ykvKeLeHEs5n2sGESAUsKX7bjRDhKSQSjOKWNzWp
mDbgz1R0ZRi4JHi3+WccYaoGivPVSJBdQX1Iq2o/D6udOOciINxrscvjls4gsnxa
OOksETZh2uMNsNyOD6ZDl38BfbyNAGmhWyXCo+D+Q47bQo1Z4LZvL1NN/+YpKbWq
PWc6lvIbdU52ikJS4nwHEwtQD3vJNOLGXKmptchmcGAv41SVQ8jx3f3aiQIO5YNH
+325aLShAD5NvNCmfIng6GZ+YfcWVBn8C4/lYY6k5xEcxRLTrY/eC+JFZWklt8A/
sPAGkQoxdFIgrgyjO1vCJido0UO7dfeG+Rn/pOr2A/xPkWfrZvRYAl9SJ4JH8x3R
T3BI7xwMJ3cEFIBZSZ14z4Na++dwZDzOmKc1YD2hnRRjjK6HljvxzJa6UqQByAGQ
dAiUP4gnf8L5qCW5VshSp395ddJhqxeW8Ec5XOmn/RYHXrwa3xJldVuwi22qDL6Z
KksYNVrP0dGY5wXiy6ICM4JHXtLI0Zs9osJVmVPO5gw1r2m0pDfB2KU1NBHoP6Tk
OrR+xYapj1wMFkNHfbOoAWoQTthaP1+bSL2I/wIUC5HBNwVMwGWD7+2RKiJXPOBZ
9cD4tfUEXaKCxOhQFJhn7Xcwue9Jt34VI48DorhixaxcAiUsmsJN/D/MMZV2LimF
snOB4iVbXlpxUODigZqHL/du/QFZVD35S2ekesmZqoRuL1rDM2bf5emKG7c14Bmb
fX7Ijtm1yz5hif0F0VKVrmO9zCWs7KzQqfFubx2fXPuwbVLoTt7bpkb38BPEUUnD
8FhIGHU/BBfYulI50yw0vM0fp0seVZDCW2osifu0ysFJ6rbyaf9PAPEaqfzXBUzp
Tvo0pJ3KnNUVdPytmKIzhnbpY2zd8SCQFpMnQrGvqX1Orc2NAZckbav29UdpZS5x
VyjyvwL4tGSh3iVOyIp+/7g4mWsUUOR/O6u34fB8VJbguy9DLyfKIy5rZuFxuvOl
alF7kT9ie5VcPd8zSmEOZKbY2+SKqnLpSo7O4lu6J71EiNkDFfLnkw5Mf05Y10/i
eRZcaYzh5jeL9F0CQBFVxe2tFHx18l5cWx4syr8X8TM5Pol7iBUj/0Pd2hLstBin
SKYrV0GM8EvFTzpQ3cysrpZ0PQdz5DmGQQQhhMQgVBgECE5OUO1DRb7UkMEB0kMw
wrvSX0N8jj7mqTzDyRZXP5sufGMtRUBCXRUfinkQgV0rwRxO9WOtI466SqKCYQ1Q
7EeISkGzqD8m9MwYPdf6PdEjIPJqD/sZe9xUvAthlRK/zl7RanKwpoM2ZgWcBzrJ
xqoChewtVw7krVnEBTiO0Gz/gADH3b4dRDJg2OV2CyuP43WQGFSZ5fOOBgNokySr
PoFniRmGtP36QZU+2387kr+8saHeYinnxLCyAa6GgjUW0q4opuLcNkhD8KCaT2DQ
M9Y8ost2CG41FqcRSN63pJjG/R9yrpkhAWcTLZd7r19NehrPn0bukf0d6QuSVWl6
jNHd5BqSuv1RSECjDwdGV8ib6YNqDlUhRt0SgWBObeBszNfXOPrAlhEGBjwrCSA4
h4LfF6wymtPFFcCjzMYgzwJ7JFa4hK1jTlW8yzNyinXCQguGp3Ds0QseedIrztph
PNrrmXNa5B8yw5uhVNfUbOYuq0tfWUyUwa/md+fXoV4wB0dDj9RnDcMq7F9h3MI5
X0TzdokeeijlpxTUO4nWu/MiXUP6g+FqrPSj6qzYbYpy8qN8dd6+6XRIBAWd7rzc
ghxuXOmXIMZaNUM+8H3pMUO0zCamIqSojzkdGgVPjk4qyqnNmAizY/x0tIJXOCIp
HiFi4IYAW2IFmrNElro6qNCT5Pm5kJqKR0enQUSvGKtZzBvnvYO4e2BRKp6IFxcH
9iHG/Mh/mUxPNxjeaFtrpSZX3/0UVtMGyFJ/CmpOZ3YvIAuip3QUDevJpyZwCx0M
7Ay1MeuAdwqgNQ9F1y5DB33JhiGwgohLNgjwPgZlKSaUQJp8c/9+fjVhOaOpQHEN
KF1aiDbUcwsjqoGJ5fqRweG8yidWV9tOkuWAjCrrUvHmSpMelKlWvPzBBbdPLsYS
MqF4UOaM0i4AkmDZFDnFVTHoR5Efzfrsj6YGfG4chVJG5esuhGG3I9O1tAT4b/vh
kWkZkJedwIzWZ3/WReKsBfdS+gZn+8+un5CYpuCAV8kJfXrziPbd5PCWudexJeKL
uuWLUosbvjU9zJOsSo6paSCOULrYKYtxaMnSazBG7ZoFpPwJlpCkS0DHSo1+JyCw
OMqru7+lC+vFXUu51n3xzpTYgUq4bd9jN2i5AKfAjtax3inwKLZcY8dFLwuxY4Pg
zFHcdD7HKhebDxuzUPbagAwy5Kc5LjT8Rm9XaB7oDjb7zgyaVlgoIhUndvuRnLqj
59ZNog7itN3//sWYcANYFrRa1nuC1nEZIZRtNh0Pg2L21EfVe7/hQuRCgVcYv7hf
iud/4f6hUXp4WkihzA/JfTqEGAClBCrHxMAQdUpTNXt4i1Mcioq3wqqpOPyQxNEc
DBDj8WD7arPMA8tyGW8EbA1Pe0MA41d9QV9nmeRxCkCFmNZswVHoqyw6fthRbHCy
41ubrpX8FtxwuiC7RnoNhl366LFJog09uGCbv/FlLyzHwB0/hC2bcgdIN31ttjbC
9X/T36+DjU5MpIUC2q4TnqLfNZNl3SORiRz5f+pWNc6TRdcjHN5UhCJLq+Js+8PT
3CAfTRz5iGo5PW9H5VkSk61u358vEA9mtkbffk+RdlJKwq/wExvo1xfrFt4MEKUE
CFZ3dipPz7DCvcee6yn0dAjUix/vNkk5oN26u/eog3VN7cTGz1ZIzrLvFENoLe76
2Y5OBYqSZ+rkvfgfvZlgbyb93yf82w5dzyaSwR7RrIRHr2b5HbqN/hnYgrnog/Iv
Pk/RLZgJcW7ihsxziufTXMvK35RRyrqybP/H0wXLsyb7RcncpGXwjN5dHDyUYwzS
gzsD7lnQg0AEYefXFcILVj38f0lkttkfWmOIeDMxUWaD0CNxK3wbkfq2fO510gI2
aCH693W46APQOycm7TMZcMvaPDyIKlqqlipbg5Ir6zXxxIbhy1fF7u1lTQuTHWrZ
TIgc2DyuPOcS8qKpC19jAytgx+ezVzhniGGlVIHVisgPof2c8bOjwsY0p/3UpmnS
iV1NX3zY4CVz3MBa6nUMtWzlQDrzvcFsggjKtwGuxiXHlkqbxtfogZtV7LUbVxcw
`protect END_PROTECTED
