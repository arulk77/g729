`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHDNF7nBliC+/zU/pXTJYJaw3MSU3jzaMYRWiEobY4fM
L9j/LBuqWu8e6eAwndlFifxrUmulVAe/Gx6rRDRZvmimF9d+Yd43lL7goLHIE1fl
5ObRXKyI2BJLmeUwFj0MPumzryO9DoG6rtBpzi4a7mKCP0UTb+k7x4twxsQtOWEP
6nF3JYnX96lxrpqgJ0o7dkX4vqHxbMhGgDg1U+qT/GD+m/F9QBBo6fN2ughwHN1w
`protect END_PROTECTED
