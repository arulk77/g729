`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePQTOyLXHFmQ1vJFsDuX1V7g1D3Zm05itiemr5YInXXv
b0ktKNicsB/CsOW3FBwofniKShqtGphK6MGTzF+qZZptDxk7KqlDxglQwh+dSdbK
LI811/S3FwCFh02IbePYaHpyhZTx6H56f4SZduRs3wcYBZAzE1KVp8rb3eh+SsDi
SduvM/unoyMAafmaNUNKPyUFPNI83UdXaRWCC6ju6aVwExRdInzibJ0l6dgCHKxA
mh3RhJSHqQomr3wfl3jc8V9OgKbC24bCmiVtsmKvZTW1Xu5YCu0iPbimE7ODyQiu
uTJ/ZGKd/FUI7EaDCNxCDD9Y+KqhSsE/O+Y2ynHzrrYr/oLcE9KEEyWqa8rvqs+H
n+e/IyTH1A+BAXun2Oa/4L8O7h6hCluQBzFdZ26uPGgHLmsDj+EBNFlwfLhqRkte
Q4idLjBGJnMwWwzqXGIjE5UB9n4XVRmUMUA/zAbcY8+YzWQXlb8mlxtnEJSGydGp
VphS9A7rAcRBhEhTcnkQjhdYhjwV/DP1Uwx6yiFhbKirxfyo30gJ8/DPL5hSXpQb
tBm281u45kOE3iUCxd2bDA==
`protect END_PROTECTED
