`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAV+7LBJsd8sj1D/aXHqa9F0iZsCA9pbgJan7nFnOE1kh
VEDKbjV61wGRTkqznme3rQHXUu4VTKA66ngwLx+2c5NGi7Jd3lW9EV992ohMEYNR
LEczoN2nCOdSHQXQItKC1p+B+dkVKwI6o+YeEz5iWyjB1j3iEW1WaKM4I1KgEdBi
Bt54ZxLEfAtHpwFoYk1r7jvT3o52OnDToasNyam6cepoXTXhpbZB8Ilr1N3HGEsI
EIJpvqgpXbRN6zsmta4Dh0q32XVv06aJ8IyrjNxJg4O9dajURpE2FiC0ALDxcRxc
R/c72GRbKOyOdoGadMSRDVzlr0qI1GTHNcxH0QP/ZAdoQkM/Rn1JFuALZztn2CZ2
MDeDy46Cl8Y0zXpy8kVGdh+YAovx01Eg2lGHuDm2nvshxdNpTv2g2B8xXSCm71GN
lD5zGUa3UoyZdS9FYJWXfzADTKUGopaB6KI1HK+1TmLwAyJBEKXTaVmIAu576IAO
8Cbf6aneX4TWaP1p7g2WXrVLc9iJ90DVSsYG1mfGNWxnBX+SfmPaU3Uz3YTH9if7
YKCBfYAB/tQFZO3VdUFTg/et5DtDP0edVqTFh1414wvqQNQwZhxaF0ClkQ/kVnbN
1JbuCwMFwbuasBewMdQAANyGO0SRD7wZ5dpwGDATTgnFzHKCEZUciQP37wPkE8mL
UlkLZY7nXs2yvkFlIwJ/K2SFYczWRWd1m3IU6tzE4vIHuPIeGVO+hX7yBmGk1m7g
5ehYBWGMIIUSrQ+0tWcsyu4QEQgwCa7TjjYpXDSh1G9aTHcOr2FgqLb1PR/M5VNp
eve8ubqgVfJvH4Z8NfZDsatWMjk5Swu64vfnSdFBfFNhU1N//iyPqYPqAKi7qLQu
c9Vtmqvxtvs58VhZbpGCC1Y3+HdcbNO/g/LWaPjhDtzMl1uvinsIwXpI0gd3fysr
4cnTV4irD0az2yFiRq+jJMiGJJ1y5HwaSiv/yyR6oqdE0MqSIucfnol4mNgx9H3M
7rYIVxiu0XVVjj0vgxvwahoeabQyPLyRnDzRFF1oqhnzhpiq5bgpyWicQEflB9k+
38kxG8pYqUmWW814YwQOf0rDao45/5sbs6DKB4kzfnAY7OEqYvtsVEb0dvUCfUTv
O9LrIP7QWnouvmimrZ2J1l7GHKwzekoPcC24Or2sc7Q2zJE4yEaXO7FiVzznnCZg
wGEmZ7c0AdH6jtkatljfLyt/ZefllPOldwroEn+DnmLlHONuMd2HrnDT/uy+ziQn
c9Nw/gAGjGmoPgNxYxLaGkCRiNOvqypmmtb//bjREN9Qp14nrGobO8f8AhYZoOmE
QRl1EWwTJoUtWuTJ/x8bAVOLB6YGrdutn/VnvGS/re0EPWdO4cq171OuM0Trye1C
dfNLpZbfO+KImUqcGcBPZjGGjufQbOtWVF/3BNy4AgyiSJauN4buVVJFMJKXUwxK
W883IRAB6D1jdUXbGbtRYurblCIyENRD95ZBM4kCuFlrDZglrIcDk6a+g9gAszKk
290lb99TsykIK+/M0gP/vMBS1JEHf9iYV6Du2dvc1pQY+rx6MVOkBSot1FOf/v1R
ibVdRRsUu2jrcb8OAQMvIZpqLtopX7K3DOwRfKeUzdz5jpTQCRCxN9ifA72/03wx
HZdy51HMWQe7Ht3FBQiaO6LN3CyP/6kibDpU/ZVNfcMYbfnnCmHhO+unheMy1HA5
41oVvgi35ODcV4bX29PakoC1B/4QLCW4zDnTQoDsYfIxBizeH76Or/iAsm3sF/hb
VjbnpA0FYDhC5/9cuVHyZo8yUWVx2teM+nrC/XaYHTVhBaLQ/LCrVuVvYFkM9wg6
E3a/OYCTItzxbgAwU59VGvMV+eyid6hvKVA8Mvu+s3goeSCqOh2GIi/JExyNQgkF
LaPDrzB/UYla9hJu2xuZmuK/J2LRKxlJXWE4tdiYmhmIlZ6yLX9JGcy1JRmLjdMI
HN7NM0IeVbqELi9FznKGKmQpBgpB7oZhfKvi2/71Aq1LbCzpqrgwrsYtXhgAVsRG
KrLrcfDV+DL1imbDHrovxn03DenPKeDFKtN9DaouPR2ch7fK3KjJ7hGsvKEdpeJX
TC9ewTk83eK7kP1fTMPe5ukTQo/9QKV8IzXssLp3FxBnPKVROdLg19e6U1iYr0nv
qFN+zWk8PMostC04dJr5qtJCwjOVaEYujWVHVd/NMBtMh1WOhEc+ZYmaWcc2BhGM
wffX4oivVTJQ4E0KSo+kMuhu00Xq97BaTDlp8gwCxa80ltDKbSoZVhn8Kb6n4AQ7
DkShiqq9FxZ37HN+tPrCGCsyGAQ8CpepdCNepnBV8vbC/mxKKyiOnDzVBPsDAFxL
G8TX6jKJSO4QwA3QTxuxRwoHsiO3wTLB9iL5Vwmp/gbDdlUG0rh4TSN0CSxi/r05
ZJUwnZtYD0w01Z9w+tBD8Vx/lJBsu57i1+Q5LJUsiYG95BCJGB3n5bZkUhZmpaVD
Dj3wsQZTtUNLld6/sYYREGMO+UGYlTjmy7OtxIR+huzO/TXBijVtcNPyto/Yug0N
TtigmyAQ/nE6kRhUDPORuB1rOn/tzSNicGxzf/L+yC7gb7DHcSXFkTmF+HXdgzI9
Wf0EfBw6qDoi8r01LhwH0XbFuFXZH9isij7GxmniQWfGbXiFLFSSUsVy2iQPyaLR
4OLU5OOJ8Sjfh47ewaRt0G/IVxQnCSZ18X7Olzs99SuJ92xsalwBlZ2v390IJPAx
Gu6mOkDO4/oPg6+PXqqqynSESrxazUheQcPG5/GYf9+3rbuxVi425ngcL/wHrE6f
XqIKR+lv9DkqyIP4K8B2HSoCStNK4vz+jiG9sx9Kie7rd4x0OMZfxFnQTC9vAfwC
z60/umUGFAXoP3GixVL0jCCgQKiBxwd4Rwb0W5UpUXB02BlHPQ9J1pf1AT0xnx5R
t9HBtS/8EfEgoizqk/hgqx2EtUG96XqOCaX/Eint6R3Yg7ncBUYOBPkdWmDe18Z+
3Z0TDPpAovYN/1QrHbxF0zn7WYwjyQfc3SKHDxQ6qagmk0BJHke8/5NymKikrbQi
Vz7kdOqDxiD1KCZTSbig5Ojblwy8Vcp34wovqyOuc00CAIQ+nTw8QALokLaw6Y7W
6Bsos0NnX9EreA2beHfwvaxWbfzuDpshWoU7Mn59gWEepRURgFqnxD4ZmV5xvpja
ZLb4Fw/0dGm+WIkpGgOot5IeFI4+vVIlhFQRTzcQrSGtD09BIn3kvbFHQQYA/Cf5
dLTPlrthslCaVfzOx1RXqmRMj3l7Rv+UdKfXo7cvzjIm86dnF55CTNJ0ZaugS6Zt
E5aBQpm7OeUQECvlrHzUqkygorRk42fvsMoRx0b5MdEGeOgwh5zle3evTTcOT69G
Fx8IKtD67qY3Y7UY5YUu0bBvpXVtXr17X+ZliF64dnN6exAO4PTtzCXvUzj4l2Ed
Fdybs66Ik4EX7eQ91jLoINFmmI9+KaQJ7b4+p/zVl8QLy95o+6PurYIpiDPhq8lm
7TFARUr7Uoda0KxStswoXee44rRn4/RrB0HXeuSVpZNgYDVlwujQEOsjsbcjKNzg
4G0XduMG3SB4WE1B3rmzD0wya2AH7LZ1v5HDrmTJ4eRPVlNGj6FyMmlhDBUOOMGv
16fs6/pHGw4UQXfdOs23tUqKFIIwDXZL9z5I4DA9zVDQFgTxRh8cSEOmaI+3gCVe
P/4mFxVpcIpsl8JQ4ULsSw1Lh0QIJCrDqzTZe9nxD34SjNusRPH6RWvIKbX8AFN+
6shT6nYer0Ym9DlUv79IphJ5OPhmzQe9Dor/0VRJvsaLZiD+wX7nPULI6yh1iZQA
InFszZXu4teAq0H6IplqiUDvr0vTVG6oqcItYCWdXKjo0aM+c/m1WTNndMjmD7x9
0HHLKoEFC1b1pQyS4G5oPYMOUVQHsqyVaYC2yfYQTR0YZJ0M+ufVf9H7VCEGfHec
GQu0YrrTVisqEaGcY9aDmoN17iJLYhlDEsn/SKzhHoiiNbU9CJIC3zvDGubb1tb3
mBic0g12u07aImYy57VTHynIZcL6jE9rMGbaWT6pox7JFZC2zTGzdHH3djLTxr7f
isMoK+ZA5jc3O3yJakjmR9L5G++uUv+tMJk9PKhLAplJ1kjYPSfCqZK1Z1HTCcKk
Sb028GFAGqlSBd74EUTGUUFLMgD3ieIi/Ss6IIWibfXDFAgCgaULoFtXWneZp0Jg
FIkOfpilweymxL0aJDxsP1E9pEnBp42IfKG+sGDpOaeqfg28+9f/OQAk8SpbSXqv
PQlhJRaVIiPyMfo6/w4wk4VpkmO7JCZ3P3WFFlDZkimYo/Z7AGmRdSr07/MxknM/
v1h35OWmPuiXKMahvlcp2FDZx9Ky3D+Fie1AYTJRuFrGARJ8zSx7Vxl+oI/b9Tpt
yPIgvhe9y7TJHc+dJmuHeF0/MIUAb2KV3rC2Nw/DeYlvHEDXr5hRnfDdbONmkt2C
oJs3ZvDczLebkxgVpy8hY6HHng3RQ0RUAofS9YSSoiOhN8hZOkdouTzmBDLKiWhL
heViUU1xC97zx9fNHwB4IiaLBKxgkUBW/Idwjq6cG6TEMsUvPCc2hoq/+i3NqCVz
BKeCbIyM5HbnozeKFSn5LENsuATRugvFhQOV0Gur2/rjgFgK/730M84IwWLvaSKy
A7DUWDOvpgs1WGYfByS0KVBDZi59DZEQyK8H8APl3bBbRgXuDmDiHkA0eK31H9Fo
jmPFcJkszjsHwvDf6GoJwev/W3xhSCOVggEeWzL8tbaxzybf0UvRWMx2gpMg9cro
13l+S1To4GTNaXyUy4q09pxfKnvmUNqq37PtCygxEp3myJl0dMXhwQdoNvZb0SUx
Bfd82a+W9GNci3rBZJoaIu4IR5OWB6SsIz7MLSq7OUWO/DxnM1CFvxOY9b1NBEDM
v0gx39sacIRV+WPMUnGRgXEYh+pJilkXBwwL3bMDhNknDp8b6B5hBCji1UVNpQNC
pSFDpXreqPYVM8vgAsfpQMcTItUTRjdf/Ee5tqrLiSMYCYalS7wMBSUM6gBA3nVD
wc6/75pMlPq62FQoc/srwMyT3Ix8mXr11A1C+Zfa+efvooZGJMfNw/jTjwx9D2fX
vJB365A1bKJpwpY631Fg2rtAG70aHXUnIxE9d2p8k4RN0YGs6YVRT2zq6wYOTRtG
TL/9WWJOjxdyqWI3stm4RcUTfB8QeNDGEsK85O5Y7/j1mq45hqiUr7qq3A28ZA0f
Y/Kr70uhSJXv9Q339hSgxo9U3If3W2GEFHsjTjkZhF63ay1vJNX7lAZKlkoZDcjK
3PLO9zWI/zjIkIqNRWv8maOjTZFTorPj0KOPRqUf0J6hJqVWt9sjTUBt9L2NHr7r
5PCfMIeY/KJSte12AlikZcMwfg/EnWrz6KUrKWV9bpITLICrCsW7A9ElO/KgT7Dg
D1xyWVDTrzJbBF90WYqSjTPCPfPfWbloF6LxDwNsdeRfuIM1l5v7UV9h/GjSyfhN
tMpjtLaPkzbsgM22JixqXuJK65Rfx5qZQZfw03Y3JNA7OAcjEiJ1AOagSwjFQaVe
M6/w2II49DTbrxVq1BnsWoG4e4Uw86h1CXISRd6OyZebFQkvv0aKhTmiFeLQT2VW
+QxROZ4bfXwMAkWVjcb2hf8E9U5lem961zJ2F7ZGPC513OSGEWEOlNXlDSol+cTO
`protect END_PROTECTED
