`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4wVBUSTT3GGozKYH6GLhc/MP5jOcBm/R7OvuUCJd2861
Evmg/mC9ZO5dBoGeVwlBPUoqjzG+VWu1mkriMxvIg9caNckYezQhstgTP6DnDTvy
/M10SCfaXSj0f6Mk99iBcbsvBjiZX6aZ2UtUqvzbcWLF7aASDX5ZNBv3eKL7HCo5
KmWR9DOSGm7CvK5sbQLtWzAh9PiShiI977rlGeVaG9zQPi67uRYzPhUcEI1LX8o3
rL1GC7qQdcXFBtLp3rs+4WENeI9VqpEK4QA2pG5r4+t5bUIdjdiKO9rHTQXD31UC
coW7KoXSVNUivnYddpzFpRCYbvcn5sRQXgH/UGiHZ1xpxXD+a++Tma+ahVSpwUgg
riE91jhtz+WgAWcL4FuOX9siuCzmB0NN33t3ZJV8slFPpGQ7XCS2itLVBbcG9ZoQ
o3WS40dnH0Xi4qnflodcOHjWWprEM2/z/xbBQkzQY/u90Q1Ek35UQ71SaSe0UaJe
`protect END_PROTECTED
