`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aZED0mrfpixnCbEJBmWPb4ZkGajoucKHf60aSlfZQJoc
XEzZAc8lnR81UtyLvz+2GxB5RZUt1aK45ovRLRe7oIxRXUCRaJDfn4kX9VVtgE8B
GGW/5tWEjXMhgBVn+OMGgx7KONARoTTluJ+rXCxXFSem6bI+2S7iVIEe4cxlnXIM
TdJjH9NTgmvk3aljA7FVdpuVyfYs4lUihbwtdfU2LDqsaEfpHiuTXkzSZD7jgyRU
t6itjVUmXXVyFu/DKjzg65/pYx8UhJ5eDXIPEzWfsj4P6bAcQcsvKy5wmSv3DQoL
9FnGT+a9uQaxiGmckeBQsbgDbat8VS/QN5EefBwxBPmo70Etl/iRZCxiULv7guXz
0B/A27qENy3GhC0Rs5X90JqU5SzNqNEd+IZkYjTN+C2YyyEmdzY5+CDi62Db3mOv
GgwD+yjdQpXQH8VyKfChSkSP9xZcrAAe3DTx0DX8WVjxA0BewJPixO8PK99gDfGQ
OwGl6Ldmnrv664s1UPy7jeSC9OZ2dycIOi6Ep1E7nHSS3qsSVCbMIYiM91UM2Cfx
uwXVGgVS3O4DM8iLgJqKsUVEntlvnIqXSjC4V4spqqHMMAcQM3k7tDs9c5bsL/ig
WOK5Oe9/AAAAAL5Va/v2mOTFkKMGHGZCmAubc69FaRI68GPTBldo1ehgf+0rIQpE
9kl2G1DT1LhZrzm+9m9IXNi2bY4SIumrEGHl8K845g9op4yMf79eplUJrKlE2eNP
PeG7gniLOZrXs1VZkzEtWEbbfXLmYiMG8uE6JjBo5QI5qZ2ER5a10njaOYLYQ9k8
Oc9RnDAFo78xyGgeqHSIx5pVKDrb27ADMPivNom4HFrOQBb5TSCrHgTd6j4kQNND
9u48o4dNZdGW10bmm2h5wXq5Z0yYRfe0+2XfgkTqJGvJZe2HCQAhUh/cc5OVsLnT
kauOTd3bCL7yIi142bfv9G4Mp/t1m2E1hhBwNLqBgNvGg8zZ3Qxob4BAr6Vi3/8c
4BUzkBm85t0qFdIAJb748WRxmt268AoiEV7pdBRmR0gEBzDyPUhAyHmdCgmrXCAI
CbV1xXF9tPkDbemeUZSCYaHSFVRSLm/uCvFlwapl5UF3ds91pm9lRLISaYiMYPZw
126hF9KZ7b9r88sodUfQlV3bWPJ+jIncBCL0wo/zmEZukL6H8UuufmZT0jXkE4gp
AIVoXBtsh53spZfuHDyFsPN2P2YISzpf5SmiOJiV/R+5QlYe7EH8UB9MHRtFnCx7
SflIxEs7E+zpFOUIxZYllfGN7x8NCDrcFD18Cf6nvIeikKEEcxOGg+LJ1nlNLrOz
pxqy6RIlpUnSP5DgpEl4ZkYkAD0cwhNpKCi31KpMM3Nw7gP37eXLB/B3QYYtyG7q
grMLu9eOEoYFAPPx+RheVij0Z7hU/M2y8Jck84pAcDqvE30E5hyI0ZztCHubcSuz
AFVoC6Rg7Z12RA0nX2AakiVMctYNMBY38OyHy2bs7ZeLqniNror+BD4sxaYfG4iD
S0S2RIi1rgn5DxI4KCsdXIWmKVLV/5z36CDFvTkKNFnTwEt/MxFNUZUAZ9M5snKL
KR/o4P15H6n0vwRHHZITx9Sm+av7BKnBGOnUNVH8J/HXELoX5Pm9tQP7OXbL7Bob
CNg70/CUesI6FY1LzPV74o0I8okotWuhEQIBnu857bbgfD1A+SlSK0LAZ2O1L0Kx
HZUJUdGkwRl+GwgWWKfmy+F8bj1ARWjgRjP/NqV3tlKLVTRgdfXaemDczOGFtlk0
5uzxgzrnc6KBkokRJekVEBru8i+A2kxkAE4Ag7ywwhiB2JN0GvKmg8qlswccAh4V
OkNkJg42KjjeFrieGKeJxRQsaEDQgFFj0WXfMl76YMDW4vLzwDiXFoQdI+L/Cdod
qK4Y7HThhH6dL8/5TQXtWmEXbMkQawtm/BQPR4f1cmHEFvO4wApCVoNzdGJUjsC7
/07kibMSG+4J56HNpk9KYaKan+SkdANCaPo79K/Aws6AwsrIYehiagaiYUqKrnUS
8obn96t6m+j0epcAkkMZ95u8RUBqGU0DJSkQ0b2eQI9VEXcMHZ6H7Rhg+C6hqbtd
Z3Gxtj6YYTLw11aH8kt3DS6RQ+MEd8qYcia8H1Zc4C+/FjAp6QLGVm4Z1IQpV2M3
SRmMM1iKXt6o1AA+2cAkrvUvma2X30zXmd96G8h2sCIg1LSoJ8AgHSZDcWrBG+EW
0HfQ3aTXx8/IgYFf4ZswVGl2K2AEn5XtE8BnPDdcrvUUS6olB/Ss2A6Nruud28B4
l9lT5PyM1Wi3SlRT2r7TQlRbgHzZSz5BRQ2FDoBazjWapZitxmvfPxS3ZNvc46Kn
OlJPbuKkOvkVCvL49hTDP5mIwvGxKSjw7EckiCv3tTkHz3OENyXhBCwKYGVAgv5G
o4peFjuqVASuApeGcUueB1L97XWMPkD5yMhEw/t3Iku4ddHDLiRIDnZwML4hB2IS
LsxJXvzbJLCsTCg9MRgQuCKgIbShWY6m0ZhMZXpF5nir14iNSylcUZU/PplVu07L
TJzqEmjbYypwhM6dg1OqNGWhRP43YITcHEgn318qCY75euwn0L8AfIE+qYT5tqjy
guLlaXnuyeZ7+IYGfwYw+bkYqeIop3DDm3BNgyOeEPU887HX+/CLn2B1mGM2va5W
UDAcjqgyImvhEsXNWe7Xr18xEQvQDip3w1pyV00lh8VFjY3qdxDBTrdKexcOrVlF
vxT/SZ7Cy1T+GxGyXNK+IF9wPe6mCwC85kC7KuJX3ckCUhx6ysU+YH8cKP3k2OPk
H83v0pbpZxEHpSy3ibXtWvxfcWVgooIcwkMNSokxW+TYRyyhP9L6uMMiB9ynYUlA
bgFE/o1tD9Vh0TunR2iO4EciYpk9hWZvBU3RKfBRkkZb3hTdJVdkOoBhYafoetiy
Ts8Dk5dlZXFNtv6nyBHIdFbne3Yfjb+SyaHOGCfg7jMb6uRHo7eL6G9BBLRDAS/X
2PtkLcFM1geXk0TG5IbWBCLPu3uXhcxdSg2k6+kyptw+VCgxhxS3UurrJN8tvBWo
KSjgdUcBJbD7+lU56hUhYBNOEc0mdvGsohfcrzZZXzJ/Bxy04WVaN/hxPNfNIpWj
FQ8QOwWRVr6L0CnzB6yffsYDttwYurkfMhopm5ROgi71D4/Tq/cvEqaWBudOiC0x
huF7wkF4NgHsDnekoaZf1B+/kpdU5m4ZpT6TrOuFwJ4kBjqU6Gi/797+C/7oHPXH
28Qq/PxjfLjbsdsGwG22jTrqPrjuenQUd5sRvtfAYQCehzr1Tg+Bbs8W2zPGyfHn
7vpPcKb+4IFHmUvC50aYgpmqgflaUpaqwtKKswj2IZAiT98s23SwGl90APVOMZhW
Gd/u5ScgH/F1JzziLci4OUgEdZc229l8hAMOIcoAUfJ4rfCiJOEsZ2xtOYecKwJn
/XsC+gPgh8pxIywrbUt5q5x6/s4SbMdL2cJy5hNHQhLZ2i4vOUr+SiERuAxIgPI6
qUpcdfE+Sn/IjyySa4F5PlU186MdPemRYeVhhvpCYZpYpgo7fP8zT6/UvPqRTQ84
aK2K5p68aZVbLC0WaL+KFJx6RJcXT7Gl5UEw2mZ+WX9mWQuEGDBMJ5oSkPfqsq+U
OJvjNua5NRQ5qcLZbuc/rIhzZ366Ur6rnik0lXOHCotGY0Wx7oD3+qCAv7OqrxF9
MEp+ATXXlcJbdpRX/WtSxhyqMumpgwfIpcwSsgfmupmK4XM9nlwKuTPmx3MFc28u
lR1s1Det0AQzJtcT62yS1SbDR5a4kSzKqjTANUWfCSgUESYiQUEtUDmgdMyzBChv
NckKVH1ws1WQr5mUF35NmkWWpmHv7HwKwwyjprJ0yhcEq/EY4Rm7bcJ8J630qSNj
MTg/fx8zff6IXlR0HACk5fss3AeAHY1rpM/pWWBUEwgX87p5c6oxJzm73vTQA8+Y
lQ5Yy6S+F/vdxI9FbraPwCrGG5QeHXE2ElJQZQACnWP63WpWgyVKBBtx8zNbsZmz
cccuZi9qGIBDXQvZrpFheb0AVQ3A2drz1UKmykY36OXVXWu1bvH1Cm16fQW9IkEq
dBexyL/CkcWhxrJY2nupoEoh0e0fpTh68iXMJWQy+KrQK0xqkXjnuOUowYOJ6Zf5
btbbi6rbJ0aU4J7lJIalhbrV2vF6hzTsxhtuTkK/grV7PKI+WRT1a5DQ4gRKsf1T
xcj8th95IzMeYnI9qF1UpNTaOXWJ1pT0pWlU+DYmMmpFpit+e5UCNXS34YvxcSJr
5ha1WYhJyyxSGRUAPBIXnX20lQT9oCaINk215vCn7UHHKPGcR/awHqlUgHQ5nxGN
uOYEAR65JAlX5ZUzuK4DU//n109Kl3Y4lQnDb1zyRDOdBJyYh5F2FasTMA16wMFC
Dgb1vlYLX9/1DOkAQZP1JKbia/IOYqtnLYlLAqjI+gnoAuzaJbeweR5qGVZqoV4U
NwC4m/S5c+pkoT2lv0FGPI5hkPY84uxA7Hgd7Hxs5cQM6UGz2nn88Ml20hKsYIDF
wBXRy8sK/P1PgroDttGtBXTS+xBsYoRTytzMN8tPZrgQnKrdt9UqOOuPN+YNWGIr
LAm6hnkJXyc9P2yUce1rAZSbe458ksfUUAzJnQ81+eTWrkNw0mUPFEx/qBKBpHzf
tJehy54mX8fmksi39BKaKMlVgCKVQK0cBf40bSbPFdqwwhA7iaXEiJj7QDqJ9/2T
hX9lBCOFCnnYYZ4EPXr87kC5vbvq6UPNhig74NzRnapZpMT8/riQYWX/qUtd3Puj
2YUNROMaAO6c3s/HiIOHnsFwas8W2Z7dv+CReQRUpZaXhdADFv2B0wyCGRDgUmEm
bO9CaeD7X6zoWKkZXZYyKj5dmNmm12shQqx0jM+StKqXtS5WEs7IW7WTVG6N2nIu
bxeN7I/cUYluvCuEFIutn4nU+JOZgT/OX/ZPypKvkLVf5qlcvAw59EpxHc3qatd7
lF0ar/kmQbM12dFZ91cJhoTuv1Syi8cSPdTgaG2/TlOr/rq8Z7CdPZvmgB5+k/V5
PRLDqea1kioahYdubUjeD16XgAdxIE8wQ2VixWVNtxLBWUeVeDOHPL2dWwhlIFh5
tsqIHkkqvqoWspCoGaphFPARueBYMEBbxqP5xk3WPDafrl9cy1sdpzjF7k+Hq0Pf
ANy0WQ80nsLMqtecQrc5+QHrLtjMahjt4DF00BKjLv6QV2g/geV33zH1Bj4NKYQQ
WF0954zGgSm8N1VYjRW/or4WS8FJAmWN7utQEgdfo3jGzB0htDzH/YfNQ5kh/fp7
WPQmaVvlM1CkeDW2T+1Odo6Q5zP60Cga0Bx7Xt3sKtZOEjxkbeFoUQseCgMX3Fo9
9Z54hQ3fYbq7EnA/nll/EyHNe8nbmXvWBgzZeam4MnUurEQsYzqYJ4Bm54tMc7pJ
YCaGwrUcqYHOoboTQiMaemR4w/J6k/Q4BatsBhUiEKj9MXUrNsyel2visqKMHJbx
GRxxcRwSnFW3/ChlZcLPZEHW3u72LEVHesMChQk5UUnZckx/YWBPBb+78825rWDl
bLL+ACLKgeA+rHye7rD8gObRM+nPO/unWRqk/1ObNAGyAJ/VEpK5TO4i/BhQibV2
iJZAUiDTBi7ElyjCyTiUbi0xJXCc+KAZaRbvr31uxg+FUP57aMJ58lWdL5ivbArO
vXVgpPVymq07rNWnXdbdeCRWbiAIj4LmLGAQt80SuMvR49fal97CORLXDtE7cAYh
yQmC2uanaVUnSZRVhrc6CtZP31xSvibwNuimPFYgzCUhAIc8QNnleRgpPk6YBE45
hy8W+WCSl/QnlIUmI3VJ83qRt8abRQqKe6P3hg5R2rDz+12qrXS+Y05cj0i1n7mK
JadsWSs4R9nTpXYtaGKbhsXKucSJA6QouvMi4P9eOAD3xWoblmjFjOXt/GYRS/Ka
S5R136VRwqpJnMiRRD7t/uPanICh5HVvRV1/t9IOhwkV2BimEfzbiET3PMaItvxh
qbnlnejpQyQsQH/4QLZdhfDd6L3jJOUcbG1bawjLKgWPSh/Spat+KWHKAb5HsP9z
v3SkptQLVqu8yQmpS3DNW3MC9AR6OLEdSqAaYsf1vwkw5aZfV3TZ1MeqCM7NCMnp
8zV0ENGNMHieNZwYqfi9kBfz5ydl+rxIp2zgZkcn5SVrsYjHv1V5djM6TzmscQiK
9JSdql85JwzKRWCufoUwQjuQMlMLPj4BoUsSCR8Lm63MiH4c6oSbHwHpwtilv9R4
EEX5bvYklK1Yjm3Y069ilF0wW7XmCUq1t95eGn1dGlrLSEEtp74C8QrFsoR2xtIl
Gg2cvfivqpbY5FJj+GBKcYUEwZG/ueJWxezbzZnNv6YlJ8OQPz+G4+dU8FTAjIYi
+ZZGlYfH2QNHw+QxAiYZc9lmP2tRcN4AMPKxHkzJ62KLcxjelvp1P2TXtIu0WbEZ
zg0/BJQ8NVEMDRV1+OASdhRgj6Pgp4I0Tws9bHT2Foj6n1BN7LYTVAlVx7VRUp56
Am4eWy4shkaldCu5B3a0HSbXyNBxdVWLg3iJuJGHl2R/uiQsycgqtKqal8xODsrz
An2ytPmrWudrNL+BnjBEiNkR00EBp4lmL6es6PYdRcGLzyEizTAoKrP7l2VxY6tR
Ydw2HxXGpIyh5mhb+dOyVBlVxsfgO/jE4zeOcsnupvu/Kh7rLHDsXGxLPCcIIck7
UH4EgZl++LI/fyLAafMgUq3OEHxMRxN1++SqyeH9/u5xXTkxSC9QtzeBKd8RBVuP
zDjP9shinLXqW9GTWXttN1JFM94ZSKI9/0gIV99jv6hUDJpbxDrRx51wb7vRqUaV
nzU70cZyZyxMvvOxh/0GtLCqFzXwBR5nn2gnWtQeoLI8q3tuwWfPXx7EhV4b/fAk
Fic1khuM2D0K5QuxJMV3jUiqa21vl+3NtydiV2sj+xt4AswwKODY3voWUbYBmnPl
RdGHseGyj0jI1eSt1aDUwDZz/qIfstQz7QNMXToxXq2Z37SOPf/hI38RNUe1VmmX
TpgqZgrFHGYjO0L02DenjWRwY47ssjp96KrFMJg1V2M6Yt18FHfy+qDa85Z5YQNe
8VEaaA91FWMbJJe7hdBfWBcQCyET60lGC1ZidDp5NTg9n475aTLIzQX4J1zCvpLu
/9wKWCySTjD0BkhU7LOGxxRauOUdLGyL5re0DYLl0UJmRDa6OEUF8dqWx4qUU8wY
Jf8Yby2rDd8znT4c61+G7V3YmP5rXGbKhAvOoyoxEOWzGMKEgGpUsz+v4bO2R/J0
c/lbAmJjj2is4K9chDLTji9yNSFI8VjLWAQrTxqkeGTbgNMMWsjFNG4pWB0AbS8J
gp5b/pNUIcZyr5xIQUYhznwHTB+XZCp8/VE4fNtZIE0dt1SBIkWXKbw9lRaII2bI
CZapYkusKCEFox3fquBDUAPX0L7XdEk5daRijumow8ipR1jmMVOCojRmAxvpltph
+uL0NiO9pey00paQkEYNxFbDG4w0HJGFUh6SJ3BL6XVn1Amtb7cGlHZloyxnwmgL
6DQEDtbXMld9hJpWMOTwcD6hAfKgvd9T/1DLljM5DQtX1f00FnRtD2HujPj1sRx1
XYXxKTavCyqUM4TFOHRAhXx1zUKtUtR0OlQXmwP4DkRHgmRAW3ccsbw2O4MdjY0r
rZrBNqUZDwR2X/G2fFDFEiZVOLRIOY5JRAu5gz0lnl6NzVnp1PV7Bg2KxwanfcnE
dX4/+5n/3JhB0XpgxAuxE9EYUb7fgcsRgubR1JMaha35/tMuK0HCwZFqDpDrZXG9
B6BCNLAirplKH3z9fHVgGXKm8IXRen6TxUdfnx1+a8WR7BpO+Ji5psUNPSiCD9qx
pCgtVYipFR2sa95Uj/wqwQobd5mIW1GU8dkRo67QoYNExvpGtw3uDZuwV8TOt1xW
LGzypSEhTgXBkP3VKaWtSL2RfB3mqe2Ia3ODQTqLlBN8Y4VycXl8w323YHfYG38t
ppMhCvsVuR7k2oaBf+h+zg==
`protect END_PROTECTED
