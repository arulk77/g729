`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJopkGKERCCluaYTl+diESz5aASLzUFtJVWqr7qkUAWY
zSEBoPDOXsbcsJjYdUTUPC8IyssWFWehet55gvZGHyrBL3sSUEU70m+leYhQ0bJH
K0+1kGWHWIS3QkYUVYr575KrTa7753rJa75HpkIvHEHatgLj08fj6f78IqYtxeqo
hgHj0uaNx/ESNWa7Kw0Xce930xnV7Ji3pi5pgBgRSsq5ai7zK9pQCgAaOFOg07bX
VQezQ1pWpMhDqOFBDGnsYGFiBI+5cWlJbt2vWeBjhQFPLYJLZMku+uT05cQv1dvi
mgM45A5hI6LyEVSAuVww9A==
`protect END_PROTECTED
