`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
c3d5+qcDv+0Y1v1+vafST6XKSMxhw5B+EtONVlQSDXxFiqlRqbjr4GAoy2G32jN6
8jN5+I2H0yj89v+ooB6QCnC7aRZjdVDsXIaQUV127ybhhLG1HOUbSP+ndBzwjj07
caeuVoxap/qpK3sdmyiEAvFDzIR8hlbIGfiH9vd9CqAz4Iw41CGevCR7NE1mO968
2LXF0TxyLi/p6XBoJPrpBGknf+rrVtc9e3KlgiMvRchGdCG1fll0WXGb4n6hcxuM
5RmEJI1rGdcEJwdavQX/qus2zvIUNAQQD31jGBMuu2wwQ4GZpPielBoVFtfmFn6f
oP3agiU3Q9VopE69pTl+pXO1ZHXxmlWwFLcrRfJsZG19dB9AYXvtWYHf1v0kX1td
3iPmcFrOEyi43fk19NAsX3pFXEmPZI+nF/+5/erHa4WAOBdRu0znAvzDwv7H8nNy
P1Rq2uDDIitOGTilZ06Nyq9yKGO64W9aiQVBgrkAWyFJ6y6l1Dam2iXISPjLwlAQ
c93QmPhXGjIVceh6OvKwfR/vcaCrGz8XTrItoFD90n2QIsdERny7/afueL4ngZVg
n+cCs4wIm4OGTqfT7npj/l3D090vCfd1rlr34VbXRdifSkPBbUk2KEiKN9wST1zs
tnKQoCZ12fCUQLaqE8o67lEEI+OGIoNkdvxvKyGWw7Uf5O1wRIEi2P8t2lZ8QKTH
iCXtYNCo9ZC4iahbccF78X5l7AKdNcdcA9nbKILniEnrMUH8BG2Qaf3I/RxE7lIV
6ycQK+LQN7vOP8xxk5S02j816+QWDpf0y2KbqpPdmi6srWsfJcZ9kSdwglolCZCh
pptNfyLOj6izGBDLY20cSfpITxO17BSe4Ei8ScvFLkuDRGgIIx/0XtD6mk/6BpXV
rsIWnwfb2dy7UbSfE0p48i+G3MsC6d8TDzIwjiCE0IULDmp9wuqCv9uMY6KwALtJ
bvrg3pQPJaVD57cHnOfzkrXY086H9fBrQzeQuLM+a9P9io9NTIZgdB9y2zLYxEhq
iDpipZ05ONVKzPa9ntLiBSrh2t3Teu11nidDwtEcvHvvnmEqiv2HJbar9aHR0cci
rWiKyvRSht2XOuhXf8UoldhPDVNyp33QCxD8CszVm5gM7rdOCzKIQfUNPStVReIL
BlAf1PDEo5WLuT6lQIm/3TJk24Yb3bTU7A3eXqtyNmChoKO+hMTVJ51Ey8W14t6C
uQYznIzro1cM2bNjKkHW+NcpMAbkg9MxAOzmIlO1V9ILXM91DYkenOiavyHPDe55
3vxYatuuLR4Tl6B9s3pymaITjKwECVr+41UefcgVMrcJcuVSkgH4PjbcxCpH6Z8E
srOggPqGnAuHH9E74sau4rR3JSnSTB79pFFbtgq+HHKxQtCfJhL46X1HqaIg8v6b
0q/b2VWaVmo1x61dJGUgusN2vbYwbBoH8g8WBILwawC0sNh03igxzgzx7tfb12zE
JzQv35PRZy8DCJGJ4Rj5SifM3348KCJUjFcl8GyP4D28otnWkVdhSksFL1qCCRcM
84NcyKmma3cEevrL7ANZ3aU7ONJe5NNmpM1bbh5TsLdR/JrY/0xAWtM3iijUVvPr
4jloBURIcWAbIMBAxL9Gcavco/Ekb1bGrehX1zTpF+0=
`protect END_PROTECTED
