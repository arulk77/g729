`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
xl6rcb8Pwo+DxlmqJhJ+9b+GSvLil3bqvrUn3zBNwA6+sHiINzMhw9jzrpDS3Xr/
rUykOWNjxkO01TKpufaThEkW/t0gHSqYTfxQv6V1rgm1Iakea7hntjuBHiG4otHw
drOjHv/hmdqJNeocZmqba/PUf0/MSJ8aXTDtreMaCWmcaxaQJId/CSDo6st2oGVz
cEQAO5HX5P2Qsq4g3Hguzp8hvTtJSMkOIImVFL3jRaS9/B0mvtX6pRXmN2+XFEHC
/6sfp+cYFjgvoO74Nw+sN/tZNJT8NjZ86qsb5v5U9Vs/wLCaKAR39/TXDP7/gE7V
MvGtHsJsbzQtfP8UsUYPavENhU/cUGYPeDzXhHidj/+fk3aZ/qnNXJ3OCW/hwPY2
71dL5w9qz5uvXAu3lOJGDYfhiV5zJM6hxJY3Tvz4x/Pr94GuvJCoGE684VHyc3zn
bk2V6kN3vydVybljKmkcdswc4Nx7oTwSdL9HwwTUGpBI+Q/uXBYUhUMXvUoUDPyF
VrpDYgL9DR+0rY4wNEcmZv84msRqOOJGPBz6rfumNKampsZPuHPfPUQkf5kj8Kf2
D9v7p2PAH6WHNsbwO+CH9YCL5Y2ie/qf3D+kaXxuIvM=
`protect END_PROTECTED
