`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOXogdsAaaQlA5eB92dgU32771UqymKyuw/FrHYphLzG
NYvY4h4qwp6xy8RY1veLdKCY8ge6W/x96jtakRyyVkDknrfEf21JBkHeF/NNciVO
VEfTOa5UsdMmzhTPB1kD8YU3ARcrtwk6OvETjZ5zTMFVQwYrpva5mgK9OaZtqgOP
`protect END_PROTECTED
