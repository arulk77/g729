`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45to8uHzqCaB8vqM6pTpBYn7cSQftkXo9+POE0sjLTPx
95w2EEoIyQsdihNz1hxTkf3m1+3/D6dfBHxWkLWDvB2QZgy1OHqj6zi5N9IZWUIX
RAUYIUuyFqm5XWZJJurmZAdTN0e3g/neeqTDHr+KBU5jXyhTSbSi+3CxDOYSTyUm
fQmpyYylkaydvtTAPDm6wcFsz2HVq2ZhykdXyjpuZupfGAZqh3kzbLDZtXSyc0/J
C9RsnbfUVsxkXshRUjKfYcn4YZnADGIToJPCPm+Quja8/6tZdmCBSCmn2Pl5je/2
UPEp62pabHFqtPP77vhIwE9MFtdN+wNLrQdxdyu9e3f2JOqkc85E1HurD+dkCuiN
SfmOxzKipdLLpfDvbCKFGwRYFnIYUY4zmrXTD7Y/RMihtNzjtv8OSJ4U/MiwRMX9
8gVV3BFgXm3NIx+uDRg5Rw==
`protect END_PROTECTED
