`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46yjuxE6X36yIY+TfHTbmehAiLItJmcCrb4OWuKrnsPd
tDuXbNwfQvj9jOrQd1Wy3QBUpWKC2gViujqckBmlpNpeDJEcqDwtrS9iUr6VkCSG
KcmxaqGpVbCjrO/xYq6KFn+h4ATHKV6llnRma26kgqmMY8uFtsyVRZBfWxoCVqok
4zZCJcODghODwQABOC3WTH4tuJlSdCqircL+dAz203+izv6dOjB4hmmjlOWOKQGd
mfrdXtyMVRuAndMyGA1JvhCVdOP4cPUCQT6fgWysOHQ=
`protect END_PROTECTED
