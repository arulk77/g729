`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
uJh64NtJdRZM2CkaAsvOmSSSKOCvAAXEfH10z6z+xKKjy2AzI8+X5c/b11KXE+lm
KS7eVodLQ2ZeM0OLrBWH2qf1LoRNmN5xDfFDZCRp/TxOqSIeGjGul1v9Tv3NP9lK
M/arEvFxsJVUnEaN4p0MWoz/vRr5tQiEvfJnv9CisUUYB6qd0K2HHl/ha7EAUwbb
`protect END_PROTECTED
