`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHF/InwP2KYKz9QG2wdfZ+oTGiBx3iMekvuUP47EN+ys
qkxnAhh2pv5xOiDgVOnbuhbhViC3LbVCU7COEijuqeNznuvsyJBv0AkuhtF0j7Bs
vb9PGrGMowNT+S+OQlxdKepgVU1XsBbdkUXGjsAQe9mHrJJKzm6Uo98qIXdeLGyT
xmeZdAeTiAHzipVf9NH2Cia1PchaXlmTWgdstCUY6VGSaYpEJ6y64Q/Tu/Jyo4bw
lNaVP83SDUaiFunF39MCpm/EWg40d/cYIZboOAm6o2le2LsA+he92sCE4evL4Z0e
d59ojZmqRVH9XUnKYcWIWOG/5PV3SK7Tfox2NxVm52Nfkn1dlo36aHFHLj4+8NwS
yiDVTiCXw7YgQdr/aqndv1kfV3K+ZWaExw7oP+F2o3EkNmRdK+pxIEiAvoRrkHzj
H++0xWynnt9EQGl6vLob1lbyQDlSOSiT+9XYKNU7YDjPNGV5yO7IKcX9/o42A3Os
quLryzt4DDjsr2NBj+vzYRYjfV02hhzqY1bu11strUr6nq9SvFJMf5y+lAtAfvT1
`protect END_PROTECTED
