`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
krUzKrhNIk2h50JjadszWvaWLELSoLYTgnPNN1n3Wg6P+Ye468JCmCC8eBhWxoA3
TsF9PbIoKql60UX+uOZXEfq5VrCrhI5YzDY39H4sGBbeX0yc9gXHmgcn3A5E2ynp
M9mkaT1sHm1dazJF7Z9dxXNIz9BvDuhChwpt1rvLNuzpSBbU9pe3appjr/+KFsM2
1xKnMlpM8WA2Ls2wiunXV2z8+3bkXfSG4CRaKf92MyCgRhMPFvDCQkLIQQlBaGBJ
ykyEsMf5kPJZIFg8Cw4VuodK3pfVJHacYqMujkx1brmf93MA9TqFqOZHIPfMTHSW
QMkRbtxXJSg+bPPvdBNZMd390DEetfqUPO+XhacFDaxKruTyK4+RCpAEuTnv4C5Y
/Oc5BTJ5IVB0w8ZLUr2a7StM88+WbB2jH7gun7hazcw=
`protect END_PROTECTED
