`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
f11uP3tAS38J+2XEq2c6cFfQbn43S+1Cm7mqrVxWh9Au3yfrdJv0lNsniImlDbdJ
OrHXeGNJ/O8YHuIBILFgvjqfOhfac1/EGhGLPSSAPY3424mMmET38bzdEZ+YEWuv
BmD9UeefQySxN1O9gFHorbAAo2aLY4IrhdhHwoSSBdf62dRofIhKHtXHN+AySOUk
5QAQcC0A7lO79Dx6F8nHK8NqAZjKAtjpL5rOnI4uz9Qrh2B030NntPl32m86qqqm
UkwaVq5E2AXpKS64cSraVXGdLnlsOUbYh8sF8TtwvQruvPQvEfCKY+K/77eKqMwg
AXdwdwNy/50jDY18/btahM7efALcuwo07a60m5k12rOpGdYFcf//t0mATId0q/0C
Lbsy5cMxQpEo7WffglsCo1nm9Xj9UidRTRgDmiJifKU=
`protect END_PROTECTED
