`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLcPCM3CgjXLOkLIFB1frUNZ1M9hratpJ1jB7JBsPoaS
mpogHiFe3QrZDSfdawaQif2/l5lip60GFUS0u4dJakEYfEOpAKGtNYQAtvJlj5bM
ZvoWpAWBACMPNYst7j4/2SXv1WDm2nOekt4TAq+IZrNDUHKYNCVCPVLJC+2jQGjP
PkX3Z2zNhhLKcrTLbNhTWWdf9ONDns0hWYc1AVqdSJsN+GQbnI9ZnP03n0UHuKX3
4eWnCQ7P3NnazFnF6tV6NVTnFuxQRMS1NGenwMbszBeLWVvP6wYl+GkvmqcbfFn/
kk/76FXAbIAbo0MWBYeQi5RjYE1BTlVy7hKRB7kKMvRQ7ElJjnc7C4uyD/NDqdhM
+izttnc4QrdhK2pN8xNykcd5+ODXulSnkyT+Nwjkoz6RLQkyKs7HvM2MreyEaPGe
Q0reABkTy46KsAQPwFuYdz5TwfbKfy61LJTFxRfi6T1G/988WRbHSMpRGgprOgdk
YFbBqQvwMbZwKs8WD9SboTNhHDsos8SPV2GjhMsa9J6VxMY9eP95iGspYM9Lms14
7Np91t0J8C3/biviV7obfDjpMz1X+CAFxQ5qKjggntaewFEH2XtoXCSLkooq0mLa
vQwKLXaY12GJ9Yop98X7aO9XPbueksEnUD18ANYnx9ps2UQYtF/OgpXiQ8jjq5bM
`protect END_PROTECTED
