`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePAq5WRLWYQQt5+7pmVMBuP2LNZT6S4xF5VIK/A8ml0J
REwqK2mxFxhpODS452k1a1DR1a5ccJO2HW1i9SVroYAv7rP/8O/PI2+AZTHDAIrP
nD5Kvz2hun/jpntV27b8tfB+kRv8DJ++j7MiazZ/SmCmra3ChprY8I84u873KUf9
glreVbDTkfR+HI71ozf63oXmmWhNVQgehQPGNolhK03Pg0MbZxptfGiXemHnZwEg
ZY4fLWlq7VBCj0GXEMt2E8nstOO8tu9H4QOw9P9iFqYqtx0aBlq9QcyrZIHwIqqw
wEBZXGNHaB9+U5aFP4BGxoZ/4fn8cZ+5oPv8hoNF31jBBjL5O8rqCNTRcfs4ejfX
N4tlqP7OGc2HqRb6OkcwP1Tzvt1xVor7CUdaXDpsSFTMzjoysKO/NzlHIrkJYK0K
weQ1ALpLTcTGKQ2Zuu+hImm21b/LYwpOHf38KpfqX1+snhDQq7fL7ZwB4LhaJ/d3
pgXVIwN944rJ7c3gvhslYv1za748qymDV0J4hV9QuXQnzYaQN8eMrkDb6QDJiqn4
tgL4dJSmxiZ8C9bTIHW1CdkDigWVgQ0nKTEYVHBBrBt6yCuQnTdg+7ENKUAusJiZ
`protect END_PROTECTED
