`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ejXKjpu/kXraszWve/rJoPZ1uflHCFZMQLZDkdX4pPEmFBvj8A2dpY6x2nvVpEuU
s9hxwHJCc2LwfOVXLoyOKQjt1v69dWVVr5lyvI5KeBzLl0aCQ7DXfgWkA1/+YDsO
HeF+iSQNQqx6t1Udh0QOyqYIXwATlwGrtbV1pwdpFQ5ImpUmk8TOE3NbmkD7FIwO
SiunmyuABH9sgSjV5Vpph6gJQFmSFkk0yD167K5iZ1sDjyiuKABw/NSx0dgc4sM5
iRCcvZ6dZhB87reFUgJ1Aii7X0ixLcJj2fYWHHen9YLdJYGSmmuueSP1CcLah635
`protect END_PROTECTED
