`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4zi6xUqRnELHpfnJ/2MiPdOHAUjdu1+EqozFEInLrZ4A
TkLLLqVxwm1FZ2oJV9pyIJ1udjF05hjE2huu3T410jOWGwZ+35oc8urvGsyUDdUE
432wvwe0y+ZJAj0Myj7cu8vxbjeR6Qt5IqFBzDxSg+ZBvZzttyPS3xB17yrlP8fk
NU54ub0Jy4HI4/sZYj7+moHStj77j2djm1O+8EgHsMkAwnVatQiOS+njNwpbdNny
Pr+D6+LJ0t5FvtpYUW/NxFSv4J/X4RdwwfqHdZOPcW/cFh3aVdGCnaP0pRDgav2j
xFZlaYJqrBouRPeC3iaxqg==
`protect END_PROTECTED
