`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLFG3lO1S6kvKLE5ev4thEnVudyh6CDxdQI0uujDYlPz
HgcjlEmVObQUPuuZGo8CjZaAe02D9cijOcpUppSu61FxkatHDT28q5wpilC9nehp
6w4Gy+ktaBv9JT233p5N95buYnsonuaRDli2GZennbB+CRFzgLZJC8Sf7CC2tEuI
a9f4VvF4jIy7E1tXQ+ef2PkKC9iFD+14+435gjgKUeFS8yQSwPlmqy7XdEW047yl
ACnu+RfzAGIciFTLa9j28/o+GwQghFw/fz60n6uak4wcrG8b1Oted9smNTLIxqtB
lsSbq8pTfxuFwa0I2YnS2ZGrjQrXsYPQMEEQArn9qRPyaZM/dNVFv9kABoGR+OU1
ZD7kGyUtrPwa/OuaR3K30UjXsP2ajsUPDy1azPiL3i6UwiGn/9mVZfiRFDwgUBOV
QfssJ9shPQG4ApvBZi8coHIPSOfpr0sgDCxtsscSfaOsX4e+nZiWJCHPgtOUlbR9
0DAdiG1TuDjnxcH79jjdkX+TDCGm4QwiUpZjLCJ6RwbDpYnH77FduChcHfTgvoAM
`protect END_PROTECTED
