`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j16jNVUFDkujLhuC6WWLcS0e7yTvaxK+Ccusq2xolznJyRpWANYzakQxq+K9k0wz
RDfPH4DAKVMVpFCsbVh4c+Bcjow5eo6PXRaWK1KcowmTnKUUT8h4/r8xycVIhIAv
7/H4aKJ2DBwba7jFcc6mpJ8teDPaRwTz6PbiYIKxT90=
`protect END_PROTECTED
