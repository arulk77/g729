`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIGnpD1ptviiUAvVc5DaZkY3akCY06lZie8Lq0hEadbd
1ikYcJbdAr30du8nz3SLXSYzhw/ejSoM7m+H+DvXbgJuxGxTQPW6ejHh7VORo9Vm
goYBSVjlR+LTbxzerqhW3zIY9OFSb38b6UjbKyTAx6fmHSeP16SIvoTymWDj6vVK
1SApWlo/t6xsxJefn/kZVxpQlbYw376cz2P89NrpujHcChnMtRMzp15b+wcd2dJq
vN8JiPMF6b4Nr9DfAoSoPPPxg1zoM3RzymEIRViBnfCsX8lvOgYPL+iVRkO3EAgm
g7ZjacCe7OK7CzGQ+lULcSNGMhgpP0650rOG/eloLQvk6UhnX/yqXs1YyPXo7FkL
cfmbGCdsQq/9e5Ym3FkrtfDhe0eKNaox8VcbxFrkpTypSocmom7NfVZI2uWNnQfj
9WI6eyxTDT2rz+D13tjKohIXQdEa8l72Cv8VS7BQ7TKKq1USYZrHzYuQQH5ocdcQ
tNvAYMDjXLZEfNIW2mkUfufjCk0IantPtThyQ8lBd24qzHGiijoczM/0/uEF3nuF
HZ/PWRDn5hudXjsbCrh6YEzWeQzZRDlbnpcQnWg6GPy5c5RAvLRFDZRL5pFB4FDg
/0pvtXbRQa+jawE/Vpg+UjnWNCVlWXdesNBBAH2Z7gWLPUWIsU1VVS1NoKETvEiS
HI7Tb4qygYX5pxmpokiWGhGEK02xRE2t/K2cok/cIEP38H4SOrEI+SKg9IxdK5DI
wTvXFZ3/W1BecHFi0mB3I3zJ6nrFEFCRG/EGzPWL6VJIPQDWIGHaa8648XMo1XmO
a7OFmBfnSY70h6RFpOXP0+ES4h7WHZdggqFmSWYaQXM=
`protect END_PROTECTED
