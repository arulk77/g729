`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLEUGizQgogFwH92N+mNzjDmZyWzc/xrBI/X+uOhF9dw
52NXpeDnp5OgFUYEASq9OtU9ThHwNotwV27RJnXqDoM43hoizUKti38OtlMWMC6c
a2LvMINqSupPuDHhlhnblVnXEn1U7n1VvLyzBfrn7uUZZAARs7jv/REJta138+iQ
80L+fPNafrXewMDAN2LvRw==
`protect END_PROTECTED
