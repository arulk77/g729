`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
C4lgIMu0BwL5ik3zCFkhbFc3F+TQdqQub6a5UHS8uEnKo1eey28EMFn9goQx4/4e
WQwrr2V5qUCyiQT/H9xYzunTQv72sa8FVYioDa5E7t+vOS3ZQVwObpZgRB0qUryV
qBfFwAUZofYvu+0b5u0EfI0SMNdTL9BESqhudHxHn1KKdvIdHFSgfIKxbSQe9Yjk
JGUTwXtCRn9SpXUZVh7+clcipHM0Po0U4MJMYSbBZ2iEFrfNfyrmGyFtFS3SsPf0
f6sUrayscM1elgdDLipX81oLekZV6lCWQwQS+GT3RtfO1JDADYaHMeT9H9o88ewj
UGdNdW1KlHjr+0gTYHXy0SZExZb+PPV8gP1kcGlczJ+FMD7DcQuF75xeCtOvbBUL
ug0CkhgPN8p+RjgfQz4P+RcT6KdqxSu4RO3m1SJLkj4wQHNdWhPI3BjvQoaQBKdC
kxV6mi9gSKNykRcQAH6bSdnmFUQ0HpAxBeezQmf9u1jXnRWP8/MXQvYXMEVO91X1
5DsZOD3b/MOQCDvS5Fulckx4YUbavmjagdqCKBip4hKwmjAUB84PLaIP0G+A9JzA
zlvnFBbChrWtLYLqVQBy4MkaxHa5YhqB/utjBalQu7zsWoA0i2AibCBHKf3Drcvc
OjTAXkR/U2ILZzgTH3XCev7tRA14iNq50i9UlF915YkQAaGrbPIk4WuFzbo1xWdh
Npi2OxqMuCsM+UqBg57h+88/LRpX5N8/p7W5FKTxSOTLrFnr4t+FF+Wn+M+JszD8
54W6vUDLyYbaQ2DnKE0zaXZIJhBMEhHSC0Pnjzx0qPB0q9yxxkfmpnmZQTl6O2uw
+9P9/f18FRrY4llpSgP59sQFFf0gAJD5oBh/wyJYViYVIfgChC0DoQotzombp+VU
reHjH2Qf+0baZVYWHBi6IFgONVGe18ZMFrorMAbO1cQ=
`protect END_PROTECTED
