`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
xPr8J7L3TbKGDLdYk7RkY6iUEzsuuy8LC6nFCbSzquVjK/R0ozgn0LSw0T+U/3hs
1i+Vsfl1YOu+srNJod/82FQ/IA8qwCwRy8SMOjne8FAq8eD5K8GxlaZ8Hu7gKaTL
zACNWJDsKTLl5Ea5mQuunldv4sxiwpn356tN9fQm6XgyKgrKL5sc4JHwXbRo+Vqs
4HHSmbOrQwZtWrpYeD6k2yEbGd3PHaGSVZ6QOmoqXXC880HWl6pr7N3K7+eKkym4
fO3QnmqZKoO64Cvk3+Ngm5L+v10mjwZRHj22QeEPpnTvZo63FrIYS/Cm/kmhZmFH
OHiJOKyAIcSaGYtdZwkS0KgE8vgFuAvJtO6WXoIXtfw=
`protect END_PROTECTED
