`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIDbhP4l5QB73JPKP8J0tqsT2BRIXz77qu14ia/gpMCq
KhDoptxfwnVktmawD10QorzH8bmIDLgItbh9FaZZkzU0h90TEUKB/D6XlRJtaeO0
Ua9beOT1cCo6gQTURoZO6d4XAxEQUxNYZoi9bzjDVwI+qv8HWNAHWtfg9qSAjzm8
U7bgjWHiimtCfxUomXIw98R622R8wRSZybR3X4sMYNY49/IXhXwzo5EZdLcItQCf
IzFqr7VB3SHi6By6pWwkaKWKt93MnK8ouM0tjTSUHuGjtGgMaPaRZLDXYlEA7t0R
uMCAdeitrZz6u5qLsWiHQA==
`protect END_PROTECTED
