`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveES4SaeP4oKrOsEPZnm8psHRNtKMY6ebL93IGtXyovHP
FkcMwCkSXA57+fY+PUghBmUjvByGMN2js7QPmY31DF0gXH8qJ4EHliIvPQDJxo4E
wbYZJL8NxcV5biNFAtzA51C2GOuX+1sScyt4o6nGCiKLytmYW0dczeeW1Nb1j7FH
2mCnk89Lxg1iTgnxmNWR4xZketmxUvmLD6JoWwTykElqLUxhy+GztNX1ueRs6rmG
9bZDj3uDr5YJZmvaJM5FCjO1IavGRVGCNzi7sAJf8gK+YT8PYBUirYkNxNdDYJKQ
vLw5waASi4qryna7lD58IIe7fG5THir3vD3Bwam2NrmyVzS3yig3Ny1vyagK64Gr
kYOcaFE70LWSLeIVuGwlMZkOPLBmulRnplfsKgNXHbUhmHV9G4R5OUxjsbsPKVyu
wSxnKp6x9Eh6+eCvMiljD6/CJXpfzjrezW9snELyw0s1eYjzB4d3DCUttNNAtXt2
uQQWmoCtnRLCvioL7Mo98n/Qq8WBIJKt2LuMvHNr2Fv4kgf/KoiGXqXWOLI8i9XQ
mBhFrzJeWZFH2jU2GdaLsA==
`protect END_PROTECTED
