`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
rv2lVLTrlkO4+Vr4AtOt1a/wocs7cb8FqiTJt9Mf6RUGTxLDb6nY/WfiFCUeZYQY
+XAO6XjnVbVVI2NpIzIcSvXgc2JrjWPNEDGWJFJonxaixOcGd9p63798hykZgLx8
ObFIh3ZOxZ7muRsvc0Bfnz0aTZl/PL3WcYYURH1UXs6iUJNWBY5wNajz7VFsH4Es
`protect END_PROTECTED
