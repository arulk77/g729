`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
KR6xpFOLRLCZZRdAWgW/J5Sd6EJ4qWp9SgQ7A2KZhPMqzE954ETbgUcegMfHLBIx
kpXPGQC5yIJG8ot9jnLMsPgVb7SraAwIsMOLgE361fuHiuc9Pfjb7sKiNR4+hBg4
WryES64930evpcQCrX8hykamGDXv3HDCGAoZT5sX7uf7DDBHAT3zGhBBYjoxC7Pk
`protect END_PROTECTED
