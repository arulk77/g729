`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
MSGR//yRMlnciQg8sjuY0vaONzwYxPi+h3IA2ALmoVHe9DlCD5zq0Nmot9zI2Crv
QFD4ePJbPNTsSss8O2bqukZLaQxVGzu2fZx0pObx1lKehIUSA5GMlFLMYolmh+y5
x34Gsdbi5LVaEHQUqhatlQEHIwJ5D23/x9yu6MpcLXfXpF+kJBPj3Qzw3n10svJI
F+DWx6zYBsVsAmnwbYzKgGxs0UCQ5aLmwG1XbdfVFZJQWuE1BrhOJaX7/79ng/Pa
OUk7fIobjP6xmRjDPh485CGbAxzxbQ1LMtHbSeAiy98=
`protect END_PROTECTED
