`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48OE1cCoCUMy7JfhV0JH3xn6HIrf1wX58/biYHLVSUFO
yh1B/7SPTEQqw2XGGB3NNE6qRfKWmPnBQ+s2CwGvHlt1C/UdRDsfxAsZeg/VJEY9
fAy/c6khthJOHOmjjAvZkBy3rlvXXwwqIaro/gbP4AOMHb0nMdq/scfzCr8qFDjT
0kENPFJtxPFnt8EdYad+B23cWxfLWq5gEpby7L54Q8Bhkwtp3NQ95oYBVzZ7uD39
EbhV1g2fjeL5i0p9fU37nU6LNfX1iOqfk2GD87vCs7w=
`protect END_PROTECTED
