`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAvsCr6mQrsDjDAH5w8eZOg7ePJPBPVYNeGaO69c8xac
RFdirE4AcQ3goX/OLBuGiZ2aJteIUADwba55QDosxIqlo0mh+QchcOjTismq/dVp
oQrtEZAdbpED3j3F5qtkqqlOwUHYN71FN+CdOKrk+/bNkM+QOfBnQ28MG3/WpKaO
HYyRzCCx5NzZkrop/86BFmAUhCW3FuDkfwqhmjVXpn2if3QmKot7EFYNPG9kS6qY
0P2gZMHdkbcg/B+nanGtAFzRTbfbodWRSBbfLuabu3KuEG0PSBt66AzNyJNuAQj4
5mhXJvxlS7bxWrt7R5BPNzo82PNrOQe4cV1ArkqWslI+Dn9e/wI/WACrn3Y849+c
3BCMgPayf52bAtlfk3AH7ZbDt9chFJRGDIkVsifYjSnla4xcg7yxV20V6nWhAAxx
jXOE6o6FE1K5fvyP2KFHOLXMQItpSw4RasVZRudNGFN2C208wVjD2RzIv4clpmZf
eEjfQFv+AOpfQ1aNapOO/x/F/duQxMyIx2Z4jdJj2S6a/dSGP88a9VEgCRMB1Foi
R2VJAEVANw2JY7mSX7t7gHayCT87e0XdudqURH1zRMvkz25rX4th+yHJFZJPHsti
Lbem98O4H75kjBOpTbM8eTs3TVKeVEZ8FQIp9ahY7PHoS9JEOmoQ33BGOrZHVxfQ
O13SnDnzvbJ2qsy0z+LCkP5rFcUWCh21r8I46AUqbcPWOwPQB+XnjNiIEQ+lF7dp
GX2j8+YiWMxF6M3wTzR+MbqNibRu7yZNVBacHiJztxdeKmfWFrP1IAbFAM//R+mX
Z9rm42/uJvDvRI9mPT8ecYMCLqQ53ZJfPDBBgkbD3SVEBjEjgqQ0YbFOFF8T5Mbo
/HFFDvKXH55HUH9Q6VBINx8PsOEQeqAGEhWmemZE87EqP9gzjzwtOkvAyFC48zTI
xQWEnMzTqIvOdOuRZxJ1NrxwDkWbCyWxFYs8VYPQFtPrGJg8EC9Pet2eDoxC4Di6
yLZoFeMXzOAkpL+SRxxJpX1Mg3MBsClrE9n3xiO7zX+ViVIS/8tAppJAQEPkmJmO
30TPO3MP0OrnoQ1udwcaDg==
`protect END_PROTECTED
