`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEjq6dj2J9cfGmwgH9fMOQouVDPTi/uPCt94o5Q5CfxM
DdHeRIi7SSop70nHKNujcxTCIifpdcS1icz4GHXjqq97sC7sQwo6YaKGr2DQlPxt
Fm1T66pj0qNxA1+g8b3hQalUy5Fsx1kwedTZ+XxCx3r22Ywnd7FOMmtofIopPj0T
xucIhPcoWIAgKq+4Y+YHxrQg2z9MWs+VL0EWminlirisN5+h7Q/bI8O6O98bC08w
3NVL9swE8MXGhYIVFW58/nUTzFAB9r9qk35Sa5lUIyJ6HjSjE5MNseyUoD/KivgT
Zl3FOprwIRS54f/uF4ccmgqo9EYTIKJxEPUbJ4wPIwC4bwu72ChdChl/sB1r9/8j
b/2EEx6PC4mGBZ5yshD4cg==
`protect END_PROTECTED
