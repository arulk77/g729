`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
8X9nVv/lFP2PLeIs3mpcpWfrmEmoVmNat7UD7b5ORsl2pMHr/IhiE5zIeZ2sfnlE
rxvSjntNsm2f/dFSv68+LvcYwU8xC2spQOii0GMxTo7vLrv2tv5NczkmlrnuAu9N
MuyMeGYW6f0lu5w4txL7PQodsJHhh/xJakJ0lVtDPYlgQBOVg5VlKc5eil1TIjUw
ppa+nNUA2VpIQaEOfQzfQMyx+TeVuswJuXoQJQ0FgN9IZDWS7ojYxboiIiX5Xg43
LUELpZSHx37RNfKTdvYEmgIU0Wvn5mP4A66nWinU21xAO8+Mgli6DRM+eiQu5lx0
z8EMWxkLuL/SzoatocAHP4HIBC+EU8IVyNzs8GRBYq6/mbLBLIf7GAWmvZVF6bWw
QIj0o60DeZALqLdznEOoxYwD8QHllPN5zYstkLsswqkcB3WLFeiK0tkvlwhyC1nO
bq3IbbKThlcD0jUscPLUooX4HkqjbAl6pgnO3vKmUhkMBlJMx3JWQ3gFN0i7epkw
dM8Vw00WeN5euXvP0qgpbZpHBMokAVXDcTYxkDb5AGa0NH9Ujhb3WL+oefP9LYOn
vycOLOFlkGPNmsTV/YQqrnEcBvDguUnmxvyFKEoHdUiUvmHNBFor21jkaQPpedTW
tlMa+2L3+JzbySld+7e9cU/8k0wmgEITTuVbY/CMSDb3oFmJcbKEOYuuAhrkw7Yn
R2pZ2TbYSG1Z5cR4puzYMNXbFeMUuWCHqEtm/2k6l1lmHLJodZGPecgMCrj5ATEs
B2TzqZBruuokBJNCDSvkXsTGAePAROG33aZIgnjaGqMHQpzqoWqL/Oe+MvW46SXX
HrHbIXymvhCuGrnKrbn7/LzDq8sVG/A0YOKDEzsOFJwkPmsodasSeJRqg+QOEBAM
QW+FiZ/m14Ia8HzhN6T8lj0Ct4q/URpndvAnazZGU1TQMD8p7fsmCodX+OKr1crE
6rmuaUHIn6GIGddgBaMbN6t0HOAqaGUUCbH/Ai9h08t4KoYptxRi3I08CGvDodCc
k/sHzq+h2kPyG4uRZwBg5xYnjCZTBwcrZ5yq+bmrJ2T20iWS81k7NBC4pN6PzmEV
fyhLSF2dB6pcIzQIOGsi5E2+JqFbVLai2LN9faTSwAM8ee5wKlCtxVjhdMz5byEQ
ORFBPseyIiOf1N/LjjQWnhp5KlI7p2zDGrZUxATwcvHt87ozvmgzZiYLGkMT2fCj
kgvXgfzlqBgDXaxPvRUnkK53KNMaqdLySdWP+nT4vv+aPilnKWNzxaEHhg+oy8Ur
WLIKona8ZFEiHkLK+wzq3pdAd7TQfA0EBPyk/JHDb0dXzzVBSALFqeDdjmCGAMsj
`protect END_PROTECTED
