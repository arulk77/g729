`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNzfrkrSSjeGM1NKqPyNdHuyrP+wDte4bi35olHRWNLbf
JsiCSYLhcjT/+Jlvj6VX3rYf+c620MqCLtcmSdcEh0IUIv/uNQl+vXaM2B/+Yk/c
X47WJ4ggdK51NCp2MLdZ4oEuBRC1UVCkEmjOJ8tQzyrEGzfP3+4QGmWMP7k4mWK8
COcwejqi/SQT0msVz6uWJZ8OEQgMkNc2+MisVqn2cplUtGFbVNiGC46fCSQEWDiI
Tr1auS/3eyl8vT+4sV8XPwfId/W1B5a81O9unemU2i2DSrvuCtNuYkgfd0Lr5+wy
HhBBsOq+8DoP97q31pgitWmM9rB0C/2ndpajM+dFgscXNQirbFAMu8BaeVtTVgiB
0zF4AfzFFdQlF2bx5bUvicdMi5GsT0o88cx6CCjm54qWPHorXJvEfWW10LFWstZ4
16x9aMNfmyMtUAkY9m6KXm5IY8rfMV4hwXlCqplNnAfEVdlLmE1WY3HlLHoNMPZu
MZOOVMsZsoRm/KXemctUMC1WcGT5MInB4MHrB8w86K7P2u1HS8NtTqOk6k3QG0u0
5MNOMo2v0oNetk3R1+vETVfhnYNkvlY8DwWz2+t9GkIPJnJFVMs2TvecGUWLBc9C
9J2FEK1K1dmkMxg+YxPSAiMU7c5r4JpscSRudGtYU/wbsT0ZIlnksZD3sBfjxX79
5rEFMMWrm49swMPidbj34wDiDMsCbfOdV3LIBuK7wXhJGMlcBT4xzV0caecQp0Vu
nzJHIQek76KREp3FzMfVI8bKXTq7nK2A/Rj972Exxej3+T8uf6Edt4ckWOcB+NLP
nZjHDzbWk7wvqA9bKaEnHRJAV+Adocu7WQyZwlqME/93UsUCDIhCEUskHK4CCir/
KJWSKoeZuYDgrj1nAmCc6OydTF7rwI3BW2UFCkGeZaI4IxQChjZhPKlao52T1vDR
uspL0NVBMvhk22gvutmuz2Euv7oIf5fkB5c4FTnowi/RUoG34AqKLzshIbWvR3+y
evFF4SP6cVNraygl0seJ1XJQtU2R1xrZTQ/1ojs2MwolpnzV9wE9KqHIskJgycri
ogNXoMPJuS8mRqtJt+OpWdMB7afPJ9HRONXOS1MMwf9Ake2BDKaw5JP42n26d+cc
jdOoR8eCgiAT6sV3hYDIx2uZTrx/zEDZzZfHcqT9J4M8EAK4i6EfpOE/As1MDuxu
7vVhtLsQPDgihXxJhdu5fWFImLzUd+EGuhD4jU2JqBX8xBcfbL6QqbfU9TO/WqgO
pk1tWkkZbL2feiTg4cWNkTPEf/TxHDh4W7IiAxpBoDaz9pqZSu6n4g2jbd4wKhGP
CA2OCU+MoPrAfQMxD3Jd363sb+PzgJJBajgE4l/VBcfcKfg6yLCnu+JLzaAubGB9
oqfi8BWf7sfCRf+k2WRjLyCQG8qW5k5Tvsk6Qv1CFhoUCOZj3bSFyc13A6fmLvOZ
vXivznjX8WF3Y3j1/rYbzoBJPR5cY05c463448qsfNEC2w97DKntZH0w7AmpbPNw
EPB7iockzhpiDTpp0sjQTY3FTXDXQobn0oEOSreotVBYTPovLRImTwIlpM0aVKx6
6UlZJkXot4FfFcQi+vGSk2JCzpIjAIIKQad5aI5IcBa3t9IArRyNPtrMdBNud6g7
`protect END_PROTECTED
