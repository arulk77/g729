`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aXA0OWDGAraFel0Sx3pVVWr7opEVIjITXaDeQZZIw7pT
CT9Uc150awhDrs8VvL58gSNO3LjbWEfSFDSbqLD9p/LWe6PdaEQkNudD7IydWYUQ
G9IvcbTPdrB0omdVwRl9rwzH42Cg5Qclx9TJErZ0GZACsnx8YgrBmfjIGMTA69mo
v7hY+tv4MwL3JmUTXhfe+Ub36HwWOEbv+50QJq8JkFI4ArYNVSI3qXTxwwfWCywz
GWa4ZSe3vzh/SA3XcpZn1WqxmLspeLiLerG62ewgOhJ/OpWp9EyFLmqzPG2xrDW1
x5nF8osgk+O4QTXMVHYIGFs3TvAxgfl5tkqk9NUmI3FUqTt7iS5iTjzHq+gbcVRJ
xScAncoGSu3DNQdqz37p5CO/QZvyiVkxp2mZulqBisWc3XvMnVa+twtyDHUZn2ns
JyH+jdM/ASE8Xpe2+q2423dbvube4qDkNa7EgW3+lrXFTecCAiBqhbFyC9xiof0r
VpltbyojGIzgS+vjQ5FCTu87XcZ7NqGm9E1i9PedgKeheAQsehGNdEnTNKbDOKE9
SZCg86IqQMfDJtAlCVyURRKY6gL6/vHK+JmV/dSJsWj4oJqntrjnr9WOECYdaJ8E
nkyOB31vUtTuhpkXbSy68yVHVQEE8BGkFR2F6Vjhx48X3jr1N1syUAjW23QsU5OR
ISvuGW2Wmsq6Jd7DPsAA1C5QAbTO/f4QTJ/AXPbYI+I=
`protect END_PROTECTED
