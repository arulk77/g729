`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJlkKOkXEKevW//BZyArWP1YgQD/pHfR1Yx5UL4nyKdo
QI7XUQ8pRu5/xcWe1LgELMr8GwZ/ZD/Lm2YFIhTlcPVN+pUJSeP+Iq7KMo51ZUSY
JF/PMXNr6td2WXudYAEkQWeIQ0JL1Y04WSvY6LuqEjAR1T1afXnGuI3HF3x4Bq1K
6XIgyKprZGOncXj0N4vTjNLhwynnfBLWVmJC+68M9eYleJg+lwOJiqi87JlvNxMd
01hUaDksBYqNCk39VN1L5SXEugbXYRKM/NORCcXjW4hWuBUCc6a8/k3O9DnrxYxC
T3l8nSlYghSidB5QPnvCfc28tuRa7xo8inLzjP4U0O0l24ssH/wtc5UIPOxscWBW
RwLgRCgKHEV09hTxRc+09FgAZR2Kg+gj8F+0N+EDQy5opuA5QHomKXzGOIf1J0iV
Xp6H6GaW68MQ4FoN11PB1XRRNd6/KYtgnRIyv7WlYBDJ5baWRsF2oMYG1JuGiF/R
dtZzMXfmUAFJk26qLfJ+TnWa00h4mCmBsEC+9sZ2LVHDo6qFtVd1+kWP1Dy6boJ/
dP1KH9ziLwfiUg9UNWC6dgjXRL6wkNjfdFnwor/oie9WUu/DIzpR+6PXWSJ/UAHn
aKJrIVus2oa7YPLlt17ulhcTqegQ13l+zJ1Y0NxedpnnXD0sGVSxpKKT+smIoeJO
`protect END_PROTECTED
