`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
UCiGLWfI/FfBwjVzkZc2aOVLL5pdrgsfV6Bp2N6oo3NCZYOBEyOftQWG6J2KZjab
e39VpMFHfLZhqGiM5yMwGMFd8WOGlxurOn3Y4CsG4cRhG6dmonxdGG1hBdgKkVRt
jx1IJ9RNbqF+VKGRgal3mYAxoWaq4fRrIcPoJZ9QfDei+GxDkL/InQk1o39YDscP
0KZmyekg11F+WhQ7r6IJz0XnwPOPih0uDKtoOquWAJRSFZWB5qRiGiVLiCoFpWdX
bUzBTjQWvmFvcG+EJowvVv2MGdkyeurJjWmZpQl7Ysg8TRVsvdqJbVT3wj+He0wl
a4JOOs9ZZmsVdbQRNibLhP03t0XPYaSr5rjEw9NXSis=
`protect END_PROTECTED
