`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDhSeJAqD/FgtYvDr7gWJoiKbtRINjEV3AU5wq66CL8P
h0c1EQoUkdKxKgy8pTb9AaVPGta1l5wDFH/s0wk10xngqRYsYP8y0itOdw9iN0BM
1Bk3hjIl2+/r9YcdkH+5Fb5IGsWApX7i23kMBGPXin87sUKrEcimtsfq4hDDH+BD
6U4+UxpRl5bsQcvZqb5QnNhiiOu7sH7CQU+QkeQLeMmPL2hDJq98Qy2jWfnoZafR
K7mSKLIqmuouYYowwuw43OswH1XO8dHqifkdWhu90GZTmoCa21ZYeHfdFHVhk+ww
CND0FFdnkpAVQ521a7hzcbR0m/dgVgdGJOlmI0MvhXBYqj5GLChyxJolp8sL6vK0
MVzi97z2pqsOvQtHhUakp70qYKMCZt5/AZ/q7Z7RVTAF6DZiuGlInN/nERzhRRKb
`protect END_PROTECTED
