`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bp7z8tPzuOU0eZyOpb+S6ewxnyyO0oRW1d3ONwtOIsU3vdMisDO3vLXgKbN82vfV
wsCtDwYe/xD1lnxUeaLWYjVSadQrcOz0FBLrxIobst2Bd81ta99QYbagQcFej8rE
Pyl53k6uGbHJeV4GUm+4KgrKMDpwt+i9OqvWvwyThxdWSSmj9/wixcq4OyGbXxMW
DNTGVcT410WoJGsium78ip9DQFyjHT+9jAZBib7G0qgMWcSGnxdSAc/1DXdCbWf5
rWh3AJVV013w24DlAAE5b3AwEKsssWmZvSyJzj3XtrgqwtgEoJMq3pNdqBVgLG67
hYT9r1DXnxXz2Fi8Lx4m8uhrfh3vHZzSvECuyaxXWq5JbbvhoVK0cnM8jf1uUtxq
3C15KQ34xvCvowFosXNt2yefyMr/Av1iSv2Ed6GXulOQxGI2K8SEfVFzcm82rheN
yLCK5CxoQtU6NHdrlsE2zz92fHMXzWiJY6WlPWeOVUwa7uJMc1562EgM0GCNnM0O
n0SvSTsuq5Lrakgyf1VC/Fry2gB8vTe9JcVG63HXPS5j2dgKaw5f56Z9zkxmvCXj
UcbvOA5utc+QOHZRd+On4jGmEjGSp1BfwDM3cuD1asoO5SRmaTp7/G8KEGvYPqtV
3ygprrWRQ/vnuZMZRe0fRlkeIdZtAvT/jcafq9OM1X+zvwOwiFdxQOXstMxOAL0b
lnd6nVPJ1qUnmXQ1BfBpj4mAQyDhYIeNLU7leg0sswckK9hA6DEr/O+PSvtHJKcY
/BiLs3zhHPJ5O5rqIbbuOclMoHZ+LWfkUsY3sbJEGCQ6CDu/kICX7i43iTaU8Y2r
MyL+Akc3YvjyUqSupDkvND1D5qakrT2AODmtniLxWBUUTbUGaswxp2hbKGeYohhd
OcZ/ROHjq0Yf9eG0yVbB2Tx1p4hHWLc246As5qZEIPvGBnUEItv7T+0Haog2Mp3m
RXXCo4syIqj3+teJW3AwctdSYFe+srdaFutgPXGd8l3vQD+dozUGb6t5nvvJ5OC3
MhWMwpn3+Fny4GWVjCIBZE/SQm7WW+cS0WkDJ2uV5HFWP2uUioyweyvCx993Qhcx
PtCtWnMwAaPAeLBfU7g5RR7VaYFU7rrEyVajs5a0vLcqj8ZzP9frMn2lJXoQY6xC
Tpm52qhmAnsXuoHX1yrxeyAb49hwKp71wuyTylYDiprtkB1et5cYa9jQnho4wqDW
B6ytyPybLOQ6gmQZusY9+nJy4njKyYapndlYMOdqid/YFimCpgQ3sdxLLwbRpPMo
6vRCJyifuUrN9/L29biPX9MKLJw6PkeHqI8fwubrpxQyoAe5Ft/nPr58HS7HYqHG
U6UG1AmqxQnY8dg0Fspx7mje4lBs7Hvs6ldQ13nrOFFSwCTp2lD2trmE8o9ax0k+
VeKs0zx/+FuWXcO6x0N0iU9ex4Yjidjx5cv13mhITxa8Klrj/1LQ7xo3lhRD8A+Z
z0WfmUqj10oQJbilcUzIpu3ZlINIybp0EPaismuIHBDmi3ebAlRK8acwIJrSo10Y
/5WTruqG7v3NXzSR1rqsB9zuc6b1EnoUkzaykhclOaszqAOvXFZkk9b4ECb1h7mX
rg5K6Iez/vpNjhKQc1DzPfSK4ugoxPwGK38Id7L7fj0G32oYlg/FBjxC+kEjuAT1
90TU3tmXyZ9RaD/zb9kEk1ICpRpgULrTXMiMGnBq75eMaABbl0HNvqkvMUVoajJQ
yQsd5ZKRapM0WYXNImUCH4cQx5NdpcYtdqRcaHs3qkkaIdqS0LuralcFOp8hYT0v
Scuhn4pLNP8yZv8AGuGkripPGRgxY723s1DCX086jDCzezH584A930KzH7WVWxw3
sWPq9qJIBSFGqDsxj0yhjheZ0SyzayAo8tNQVOzb1asc/A365LrTRiwwg5bDm6+s
N5ooJBFgn+Uun4h6+I1LH8AwdG1YTaHGi58KSdjIdH/+Gg3z21n7stl7Ob/M1LNn
dRgBplBXQy5fRuF8/MpXjp6LwlXqFPFSPkGYGitMZx82R2ovFGZrH1STmZrbZD+N
DIHOpZZzuVomGsRgWGRU/D4Jww8ENpdJ7qSN6cVGdr6YEv2QvCrfhY4L0GcAE+Gz
JrzEpUHycuReG+nPBux6s44mRL1DhQFXk2qdeG2KiY4Xny+EubXjFffPsw3favfq
StDAhDd1LmPuSIbXAmm90NXsMRRpT+F66BLwQcujdnyKFJ6kA4n1/gJKM9BGDYHV
bi/amYJkYCNW32GUUivr81+4Lke7Pr5Sht69Wq0YoAGPUfnTMkrDQddQSWZJ/hpZ
dW9+/4W2q7PZdj9H9opu9Ve8UEpU/THIrauiDLibvebrbnsYg3pyxAZGytDecSrk
mETpz3Mit+JXEhIUA04Dr48WDo+fAeaPdAPl+tF7XNPKTNp91JIeKasQAfPPRjjo
kCdgO/R+OgcbshJ4888DDZUR6kAm8vVlQkf5Ge5meU1942ASCZnUWClYN8p2mX4v
5dTGd4s/ZvbhFyv0cNmmWuLviNMvAGfDTzaAmT/cPiHP2xgysoM5SFC4CWa4bvBX
5+77epVLg+gnDLogfSTwfJhznTPi6RI4df8Tfo5YDM9yR/nbbBlCtsEStlEJff8O
bm7C5MGmJAkpSg1XR0y05vbauZOLEipfgxa+fDtasJEs4OZAv9kswLJAJOMnW8kg
f/dnwTHlFHYBY5LImVBCRfMujguNHGeD5vui4DsyIfi4ApQJiOmrkb6Q3S0+i/Eh
OM+LbCggjMPWn7k+0zkLLFQi4OVYEAYL3UAWWW45H45Nd/A5S67p+eGpkO5H9qTr
5ZzrSSAydDjYahVnt+5IsDJQHGU/dW7fVCNNxVXHBoZ5qEEFpd6Glt8mFnM8wUVw
dndqicmDtu67b+F7ptwX6JvQKAqhIaBXm4ndnFg0FafTovwWCR4sqcGuH9548WqD
IvQ8oSO2MBRyUldocxEupF9+eurYppVqadaUx5QAmubKPGeOJW7hDmJFdXU3GKiA
MKmkY9yC3QMUBTGV0dYMkXgjSHeOcQltXdnyppxoLdaM1BI1oJeNsjJ82aiE4W8E
MxuNQFA3oaCuFsBLteCgfV53xg4zQLJnJxXcn/0+JcAzlkhS3vesjq+5iFOlm2IZ
UICOk4XQESchd6xG+xd+yHHptLAqiaHTbYP+7wMZ23Qxp3qbZT/s+Y/NiGDbZMNK
gPBGhkgmkJCYjB7bsMszUn+5A9khDOg44Jzbn3Sl0orJj9+0BnQp8mvVhLeakeHc
cYPvRcjCYnmKpFyrynl5KvZYTnwo7xH+UCU5LsAvQaWSbBwDNDaJURyVegL595Kv
T5R8Yz/2qNKNDae730D/lh6iMDLGSWuqXT9Rp9GCFYInfqfWEx7lSZNa0e/1leMW
6fxJTzKxTDKvltM1hHTkTgb9fyq1vrGXZ0yh13m9ytzsm1SSPi+/WUgYar0Pj6cA
0HniiovZTRnxnnPQFJEnnUmY+PPgvH/61vusIrSLyZGQxxyhWHS492Vr2yNFyNIe
MgEybhVN0/J2C7s5i142D0Y09VLSgb9EzXZKy9sdujpOmHv1Vug8iEV7LOLTWCMQ
VdU9kzKHy7B3vw5pt66vhDfdfQGobN9ToQ25ZLFZvy21XcX6UELZP8W1O0/AyIUZ
Yz/ByRrHfrceDZN+q+FwemyfBaNlt9tzhhO4vZUVgmQ0SS4MZheJ1uHczRL1rVOM
knQt/NTxKLImH+TfCBJTBlZPx5ocpdkHzg3vrQHH7eCNRLKmRs3nUDezJexirn4Z
napfKl4IC5qfbTPjHBSQNJKtCRyrnjoKVeYGOVjTpVAhXGbW9DQSKSwD51YbI/li
OL6xhZhMd58eANRNhI4e7oruLLZKmgr+OIR6NclTvqtTvfHfXfPAuz2Md6TCPwdS
wXEy1JmukqGxIRxg8R7DxEAu+m6jtIuYQnOZiIDU/GZuJDzzVzVN3/DhnWcvsydF
kNSwwz1xWflcrSerFgIzGLwnREH5OSrFUAI/otPrIJH2sWWCDe3sCrjrbjNKJoz3
Jir1nZ9k9ghnxqnqwrQqeXMr+gzc5RC0t7Ixu5AP4WgnoRQPs8Fo+4QUqa8IXgS8
m42AE/9TIRzNkQJDqp9UGi8ll38DTDUkl6NswS/DCmiRL/35onD1SpWVT8btMbwC
OVNhi+SJfDMacAjeED1sUIOpWNtoMJl15FkrQi6d/dI7689yoRF4xtFt1KEzpyHq
N17NM9wCX41q7xmsnwT2h0frXLQUrG9QX/C8gabcdVVskWy2E31z+yB3/vYGMIJJ
qpyy2eSOSBMwX039MeGLrFH+kyq8FmDiQPu9nf819zk74oiOSsfw61FrIkTz8l6q
fuZEJnLHzJmGJ9rgsgyNFS3xCw57IYOJqTOf3smWUBLsajpZCHi+hrpLmCUH8XS0
k9kGwFlb7usA6qqfroPEMfxidkWezGg+gZfRnx1/u28JoWXn2tii0lcN5PyYbrGf
W4b64K9ngHq9tdwYcMcUZMzAvS/fR+Gkk1z6vH5/ZV3HMOgd7JIuWXrVZbBkkdCQ
gDmGwMVLU/cZGjtDnRL8jh9Txmn9SF8yKHrrR3F+eG0KO0hOF452QcukN8ra5Rrl
jkkKPGVHd0kQDzKkoA/ovlfpfFrQKhb2ycjg86k/TnqABqdUaYtGemHmEncdOwiG
2DZW0h+lqRmZvTjpfyOKcmqRQj/wOCEqRLvrGP51jhH3/qzcpa0VbVF55ZzLTRN/
dJsCs1j3ueZAvn8nRMYoSg==
`protect END_PROTECTED
