`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu484tmN77ggj7bbCSovOC58VxHbSnOjljSLxFOmeKkDO8
f0BIMfSLUtnI7izTTMOdUL9bMhAjm1HgbzTgNn14ws6wZAqv4OqqMz6ZmTvZQpFa
iBLaZEz7f4wmXET63+aW+9/x3/Gjaivyb3zO3MIdJNPk4SUB+5OJdBoUCMuxa7BQ
Jj/k3gTKT4TJngzl6JgRf/EXDkRDrLFKIBTKI87MRopzX3QAGq+GNCW6NWch7gaX
X4ALYDj7Bjp6aCwzth/BY8v8KIL8n/JBvNhm1Lk0uds=
`protect END_PROTECTED
