`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFC8rGzaphgXv3LzwvipsvQfnjGpBtRFvLg9e6thaiRe
M+FEn4cfkiatjWYDyIL16/sY1vqpFLajc/4e6WOtGIIi1vrV1v76eLpuO+lKtWIO
db1S8VyfXgAtk9Q6jHfWxWA6f16XZYdapiNIBLu/pc9OE4Zi64HTW5cW+ylvxy7u
IPvl9oADfTM093carQ1D2cmgbzoHMlhtvP/4BWO6lKubBV8XMaPjJd6K8/sOXJte
T7wfAs7UXI3fTH9AkVle8A==
`protect END_PROTECTED
