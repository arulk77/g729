`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1acpr9t9lWdVn5dMl0UHrpbhl0W3sU+iNmQLkicTTaAmH
t3QzopJ3mD1vKfQRvc6gioHd54GzeO+7JmWkLdULcWHNHP7jBLbSy9VaFEJ8FDol
5HYOwZlMgCaBLtA0sB3MV3ysW5vHGfvaCW73RiExcy5abVVPzJN8PO4q31O2VDLq
CrQvKLcxsvs6n5dZsBT5NJJt1UUz1FKV8mBCOR1Qbhk8GpDax9FVFMRVzetweo3e
IUdKRBpMh96qxM5cewwEt1h6pli/dEKDl3OpHzwBvSZm0ZGUYrXYYneuRhOvyill
myQxihnjMpoeNN4VNY4FJ93TKdNXeajVbwDPgllIAp4TOvK0fDRWG/BCMoXQVZNC
CUl30dggxp2gExHQoKDfx9KX24MrEknjsGpAoEmjtHx+2u6Is9l7lOniEd1Wnu6O
J6OaDK7iawiIfq4Yx0FpK0o5IRIu37+T6d0nizAjOIVLRETEY3ZEC6EfZRPfk0Q0
TdZrTuyUef06NeRhti0q0WzDNVLgpY/ZxumqUsU4zHaEymQNmDvBrNgnfKwgyMji
nKnmX928CDxhQHbcKSCKLR7ATHFedWFmkIoDjiN/fOMqSWslM9yLiIMClGONp4ej
Dgu1r56NoDB5pllLJsQS1wtF+YSd7K6uF+VrBiiVpCHHiwwhrZE5SMO0qxpoCwdm
KNr5li/oRkkPL+XddZEj9NXcDHRpEW0YZLjk2kzFMOk05hFcnJ0PlOvrfQuieNiD
sJJJYVdq9IpbSxKty+uDoxB4ZDvFT4Yg4Y+lkR1d3rnIXMEe4tK7oJGDHcgiZVBO
jBW2a6I7skmLVLlLLTfZJcBzQNjec/vs1/z51lhASlSaYsLl3ewW+zn/Y/dogRTn
QQ4mQQxXpZRRucxSfezumSQzy+G4irHhSHBjJFzEwuSQpL2ug7MbKbn/KhBadqBy
IRpJQs7rEU+n7snS+y0ZgUHnWfSNwAJbOlKU25k/dK9md+yceH9tj7hrMQyd92Mh
Mb6rdidf6/qo2l/1IsXDJYVXOFn+mq6aw7XuqPjAt4laSPWiAd6EdIknTSylA6r+
E5xZ/+9a2JNtsGDxHqq2yhAugVhJd672fEICJtKOa97FMUY8FxSIBBRLn4N1TQgw
8SzGXyGrVtuQfBcydVNyCMAQy5QPHzCrXVAfcz8b7GNUeyltDU1pEtPrsl/tyCOA
aV6uQixdDEAwKyqEjW06eyCiNd7/hjkBbkXffqU7N5aB4j8Ft2tD/4a38MIV7GRj
z7RHNBJENAhLZ0yHMnSD1GrWXdBqR4uOc+4M18wIlv4=
`protect END_PROTECTED
