`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aR0NfRkoilx+0hEcMt454qINWXDbfU/mKA/BYp8hBdmx
6EaS5clEdIbxJbhZVPxuQhUCzO4mHr8YIXNweMq8/uk8c8s6tkLsRzp8+vhnwx3u
bW/ZhAQCuh2oG7jxQLOJL2Ly8ocHQPG8yCcPs51uh4/nLgH19Jfw+WcFe6BuDJkj
W7YUVv5Je/6ClClq2J5tPOTCauF2+kfJHWVwQ2NEDTOmlyLa3BVDDf36Wa393Zgh
lbH3qUr3/nXPaAYdRIDAox88LHI5eaf6Bca7Q1i/Swur9hHya7A/LIwgds7/WdZ+
vH/Sa5E6mbGsftvloYAFojsMyYUal88PvrWM6jSTJ/UwxzwO7yjoxykk8kgUWrvq
nkTHnROCgGKxeW7qmTVdveCVfmSa7OoLvhBpJ3o9SDnlPzYNrP2KClSYUB66R3++
FIDgj38DJDmSaMYUZSAYmf53KStWyAhhUED4fxineZV5IO/PfQIJQAasFSa8gtY5
rYGuFH8q+u2qcfw/r/S8HUgVsLqjD1t0Wrbhp0OoKfqIfY14vsCTmmQmHZHJRYZH
ap2uu84YubYhaIhAaNxoK2wtO8uETNQjmyrJV0sd7AIK/pjRrS/bor2JeCK8iFpd
+kVmNeXcTl+5F6nv/lexvwhSXz6g3JbzepF0oK1QCCJ9FomfVrxYOxst9Mk0R9ao
CbdAMjjAdkv6on+h0lX7CuX9SNUnawau5hyiy+wQJD2mCQLqWymBSHzOa+rYdevn
IHpVaHHvLopjcV1u9NSDbr9jVe3C9nJ4xDn4U2cWrxkZvZBcFel83uHLwiAJnlWR
iX5E6sSHlT1SIDcRyznmHdnSkhmMeXERj4e0Bik2WW72ZgQWsih6Cc6VIe0P6/h+
QRqKX8HUg5queQGIc9bevHGAFcQUZDMJaPnWXe/nlkjFcF6cHeTQmbO0Vdpr4MxM
62BtDbtrPIH3mxLkDQRYl6OY5TuEn+7N9k9x6VfjctbKvwyu0c1sVWmmTa1CMZoI
ZNdncOUY1ZmAp2+m//oIW6S4aPYp2+0PKP0imfcF6rVD9kpPyD0NBI6VAPTDb5DS
YBBqEY9Hy2zpUKFWP3KjUxLe7M+uwnqrM+kbBWNRUPlt8Qu32db/SSVP054dctJg
kyefeyITLKksWF8X1UPyc3BlnFqnraVJU8btjSMx4rpK36hHCem4wVpSIX1dZE50
UVcMzZa4XQgAyJP/X95biqEZWdulUvDW7n27EY7LIQil+1asoMQGX14DDszYNzRH
ZLI7WZ4T06qMNECc54fuxJLqD4obhVlkmNZ5+fMzprHMVeqAaB47NK5Vnevh1xz3
66HBkWXGdypGzlzSXSIlj80XWobqJoGRKjEKYI+g70BOH8S/q3oUr5Zo+r20ygGA
TcE9wlh7Wo8AX5l/q6qYXzOuutg4sYrZ3CSWA1Q/D2UN3EBRrpEk5bz+lncd7qOz
3+gXsCsQlYEODGTpYZ37JRQek0HgeAEEyPRUfIYzYXjlfs5pzy73VE4VJAAZKZeq
PqtiVBVHEF1Q1fmuNwkPLq0vKXSohnenDokqAmkVtpF7AsaSAPRf7QC8bmpGNdep
mKKgQwd2S8g9Mi/trQR/2a5Ze8Yeyed9wpupOM6yVVDwZLUJSjchGWixGmj/jt8K
YLiKZpGnj8bkAAJNAQcgakPl9cASVPW2H6PrShLLANgiiZA2I4oPjh8BPea3290p
3JilYTK7Q/wVdTam2sBt236zl2B5dWE53LY0P1U32GVJKq/r2Itok1f8/bhpdngN
kifOjKP1qy6Hk6Xcg8ubTT8shQmmjeKyjgTGeh11ZLcYgT2ZxB/pKSEXAs2V0x7o
ZRqGfyqiHjlEbTNdLtzDZs2lE2tNpXzjEpozxBIxtWWVeXK5QUGOluhsk3u+J2N5
MuQzVXob2yXjtvKnsMdWtFVKKTrEw04gMdIsuHZmJMa9ScS4Xne3+o8tPTo4oz+G
clihDRA5Myzy/c8WYqcA5PJUfK2h/jxZJMJ54oD1RynneZDFh2oy3Hd5NFMTXd1r
+a/crtrBhqF6TT7ZqqHjGsqs6zOPGKI/15alRBx2ji+W3fLyJea5/Ki+TmFAVw6S
S7F1xwMdpXlqey0ry9thwuChqOQcAqj5Rn3oLds1oTh+VWmAgTKuXdi3h7B6TmZ2
X69pepK9hhp6D7rFGummMoWF9O91JBYdUkpOL1j+/BR9CWpsfcnb7PCRhOgrWBR6
wQ3Zn5ykBkJjU1dptUJOqTT7htSrY/RSyB76ufSvzLCyix56C0vOtsEDT1RUANfR
LY7IFtpi5coH7cNoctP17Itkmq4mhLYJ5Kn6N7kwqEW4KOtHfuPGbgmiH4MPu2HD
OxHL4pW1sXCnU1VFryt1KtNL1Si5ns6h7oL+b4dtncUFeoHdhwoI+fg2UsATBpbH
LyCxBP+N0WFmFlclttF9MJGBsnAkjNwYUDxinefQlK2UGRgy3paj5CukG6cpTIhN
T8pxoyv5s7VE7Z+5G9F54hQl+w43cYSobig1aZOWv1V5vK9WwQcLKFznjTR+TcWB
iqB/bNis6ldUeRrLwN2lpSYr8quubAzKbwf3vg7KPNajWDURx3ssPlVeqFRkkZwW
cobvAO9VWeRC8TjT7lRhNAcySDPpo867qfY2iO1cwLZc73+3Q7XQITwFrNvnYZhJ
UyZbPoPJk+VkZXDpTKV+gNlqkIdnKbxoPyEmjOtJCX9tBJ6wdPCpmZT9EsEXZBWp
YFMs9Dm0rR0OnxQ5UNtHZDe3IuUYC8JnTPt3M8VIq42lA14DMhGEaKZZdxJCQClM
/tM8YlwDohay8zu4Z4WcpQqsNGKhU/Ymrzya+AF6p8hiTM4e/+jDxu2/FS5XXv4d
FTb6GDhZ1mYMESQowvFRD1Dys+goIj0/iTzfm4HbBAE5j9Ub/wOadrrP5bzm2o/9
CvtGKEMFu6ftGa8ei7kPhsiqHao8buAXEhoAy6CIRg4Lhh3jhytCIbSQ9z7XoYnf
P8lOIUpYkx1YIpw8IVvB3SRQ57xRa6mHRlYoZU7htNQ6LQwaIeyJvD3ZasLf/HGB
Tghh+dkNhQkR5Rmfc1sSoadqexUupxU8iLz2TE38jBp/6iWB14+aJT4ac06NnMmI
GT1Z/7T52OjHYzlEO0WOZGpJGI6apAQwft5bJBwzDmZHNt4ChxQ9g7UCmAzcOnSu
TzR6sr0MRnWfWb0InguoIQN2/gVIYm0mtTOuUMUHIZesAvsKJTQyFdAp5aFdF6bk
eWucwKDLsmN1y8Hyq8B3YTK2mEbfWyE3jGPR88Wh9isvKOcKM/sK1lrFG7R4KM+i
BtuEcSx1XGfODpl2noeqIyg8CXZJ/SxQ8e8VPiPbabjGp2N2OJfRbUm7zn7HJxCH
T4UWpyP+3avk2M4Bfvx91v3JPm38ueP55Ko4vrsAkj7K3a4kDGLQqL+MzAfuNeJR
axUMz9dVdav/2OV7xCg08H12/ERfLxoa7H8PUcy0Wehi0LhrSuPHuIUrNTcwvg9g
nAq3H8jl/VQ1hS0p9gD3XDWmKuv7JZVk0k6XyPg63g+hMJ0l3eCOGD1SB3akKdsQ
onSGL2qPdl+lTKEd3MBICQA25SfowS9qwPAyD6kah87Liz6680MlpXG4UYRDbbyL
oj4myYNLCh/X59UZEXzihpOwq0PNMJRlqtidUBCJVyKHZ/G+FuOKZZ3jZcn2DFd9
Li4adFfp/22m6boOBbb3QIsq8od5IX2cncUJK2QBLuy38h0bh/4ITF+yeKLjQWZf
IBXT7ZK2xrIcFs0L7KDHRudJ+8JB9Dyhnqd/v4UBy6WlXeckXqthet4A5xtwx3ua
26/ABeAD5fTl/sMb9duyRc6RJMulfIT0TotNAfBqqqsb00TckH1lvmtXNGa8OuyU
DSgIz9yM38voRV4KlF1o1uaZDiST2sIWlKKZ8xvhlgIzUB0ak/ZbswcUzPOvRVSC
GJ7RUbJ9DHJgIFfHJvRvtKoJncvLHOf5LuDJ86DTFiKcUckb91yXXTDtOL7HKpEI
7Q53rk2f/Z9hP3CTOYYoJ7OpcZVWKQtaRGP1bpMvBqYT1PNT10YT0diNyEpfzN3f
ZvcGJX/I13Ioy8KixM3QcS1XwE1RLbP87bDv7Jr7U0EiUKy0UNkrJiVJNTsG4u0c
MmWrMbkUOYfioES2K0LTfy0HsGuZPgCkhJcRBvKI86ipY3xdzb6N0pvTLVahRj6d
w2RMKDwKJolNFYSa+fWpZi6wXx7odoKKfeMujoKDg9ymttEn0mp4g06VrJH8n+bd
JDCHbyLVPOtARVlxoNNQByta2xmk1JExX2BQ+r4JPXSy1DM0fPrY2kWMuewEzVDN
1r1eF8llPc5kA/J4oq6gNz3R7JQDLVo221wGo4zlFMJLJcHldwYA266P23oiLFNK
c9PviNix44YWfvM+fI64LtgEDD0JYPS34VkdYMa/kuMCXQHgb6mG4XrifHiCzd7v
q5pwKszGJ2rFXO0VHGf1ovjoqnelmPlxucydQ7jhmZ2Rz21WU0uoBFFIgdQarNnM
Yg51+Hpwdl3Q/RUX1+cVdNufQH0iRhL24EJxiWFs42sG52ArioWj0Rt6WzUjaBfp
IKvSKroP/cbKdfEx7Jg0Hiuos/TaWNZOn5v8aDeRU4rNovN4pkDC61JqKy1uWKLl
iTCZUAJ2J6dCTes+69zNGCPiyKH8weoJyd7F8bAAVps3e3gZiNMgeaEqlb/ILSL9
n2JQ1VuqTJ1uBEW9ilMsSUV7NSSxq2InjaalTvmV39cDKHsYBVjacccM/09/3f1B
gseBGBD5tV/Gqx6OTBP5SwjuZ1zoxACxh4m8RXFR09zm0c0KRxsybEux64A77vll
5AmNpuiQjylUtwCzaNIJlH2m3QDlU/iYtvsY+QR5DWim//KZSan3uDEfKhJGtx9r
DdHLeemuCJSm+bHW5SoEDxKgE00g+dma5i+Esv6sWuyCZJj1Ov9DmlOVhFBm0u0O
brEhhm7OyKWIsLf8m2guiaUlmxosP1YFJ6BLIp0HvVPwAB71Zl2Fe+Yu8h6SFZ6G
K1u2qybIs4lvG6wLT0QteXjLgq7n4JLnTiuB5AsiS9liqKxACyoCWwNiBmQ2fhW9
ZcHd3oXUHd7GZcFNVdMpWDbcQcw3r5cZjQVeVUPlbhHp51KBAI0oVDYUKriXRhfW
fYOyH29aj5d6xpuPt9yiQg==
`protect END_PROTECTED
