`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNzGVrFkmoh21wZIDhr7w8DMNiMEnvjeY4yNONsDu0r0X
7ItRZUfvi4nCoGelYPrCCeETwWncuoSQ/ZI265P5Od30bxynEbi1MNUQuRwJft8W
7ChHsxLSYdehciM8C6SB96rRT4nW0CO14R+Ge7PwQsj2F51tPF0LiNT2w2GxNJfP
nimWaN956HOYD9pb9YbAiO/xKdSSUr/sumLpk+pXnAw4FfaJd95hBiKHTbEFHJLp
ZJUv/boD1fjK3x8vujVKu9IY02o9ohw1X1HELVRlpyPalVpFNY+PYNvMI12hydoj
Jhzr4A7mxtxxcaAhv5xJQt1BAkkXktDHoYYQ9HRt7r1bAjVHJ/2PSqpg8F2ZlqKt
lys3tJfekibld5tRz1KS54B3W95+XmIb758Y5Vb3Dlham2STIGbhgyfLAFKfAuNc
RhHjvpvjszxwN60g+tAoApZ89UfnwnXNrub0BZqFqqyhaPAyXlFuRkVy1tEWIdQ2
ipfJGR8vOmCXnyTCCBU1rsTiWPuJFKszT+8Ff/fI4N5hbJK9unRf55gR725TU4ch
zlae9WnO7/AIPZ0zfoT0Z3cXY9SbxmMvmwc52t9xJpgTJA0Zlej/y+RCfH/8WV63
D1Wy+svKmDEiPbcGGblHHujR4pz6pElMQFlzCfiSj3+HpX+dLoIkzjsJ2IY/Ja+N
7zXq/7OvRyERvphQ4/i0/a2ty0aqfn7/aRgWfdlIEC6eMy13u4GKLV9FNIR38UT9
FCgMvYvURyE9OfkHJuq99jwoft4MJp2T/E4McdYRNtogta1FbYgP5wbxYWmDhsnW
0L1EXqVszOMkADL9VbLpGy0hxtDkT1W9lsyPmOUg2zD1Pl0rnWzw1eJMFowroLxP
IOO+aZVdA1EGuJWszPS0EYuGUJkolIKpOzkea7OX9jSUjsdS7wYJeLgbi1GCV8Ys
MYRXXFk+Rdgye6DD0kYQgdyMOrHdyA4gRiI/Og7UXanyOuUfRwxy0LgezUkvzXMN
ciR+1JP6cvkH/erIsK9+TmQh0etllGqvuVih44fKRJ9TM5ASsjWqAfsmYBSW3KiW
R6x4y+DiQv7Bo6UftUsQjIXjM9GCwz9ETGpVL+4ioqvQIfnvyGVs65j8oNY2TzRn
fWWb6+lxpm9yYsrG64o7x0MsaUDXYD18cvwKQOLoG7Q90xc5Dkwh0jm6v2n+hBT9
PTET/HeFfHeZiPTmBdd2etwnngC3QQXcG3ZOS7f+m9N1YeRSJhQnLmjPI7d8u0tQ
EPPFjkQro08XYjlyo2GG4eL6roUnpqFQ8KXlwNcLUTe1jkqyW2ntV10PLRE9TPgr
3K6Z2EIG4lOzxGlq8ROphkjBJVfgeeve++YGfEZIRgCq3u+7cyJgzO9Y5ARJO8bF
4gqnLcfzlSarItJXPmHnEwMs7YqdSC8GXxNuv2RW0lxNxjL07xecma88o+wAlT7G
3B+OUPUGM739bwxaY0B7Z4FyTthkymg7rpKFEQRuajDB6dUjAuSBRp8S+QVjcpLp
HVx4sP1EUehymEdgPRjOrfl1z64RH9VM76ZVVUtCqKrjj+GhB3doGMNgSNqTwUe5
ng8qBbJFzUFB9sYogDPwIDa5EJRhJFqYimHzLAshFWPEIW/HC9OU6y64OQMoq810
HVFV5WA2k2IM6yUMdB6K1RREljHGQGOvw5mm5z/5Cszcr9ooU0D9I772lnttqcr+
dTe27BCLYWBFbH9a0BkSqpx3TIjzmDi59oFRKEu68HfQweNVdDrekZ70HR0DUj1W
YNEttbp9s13Y9KVb7GSxKlVpHnaMIjGny1ZFwmasRvE8DG/Po6RL0P9UTW8p45ni
hnwzJd/rcyiT4/iaIievWgl4aVqqZpHaKOgInbtAnJCA7ri20buijThqZBHduaT+
JNIG7ap3qhaSYc+Kt56P7oz2SBz6+4QmF9h5ScPew95P/gp2NGxKU79UjEuZn3Ec
7CmoIxszfsDzbhV64TEdvqyB3kaZE/b8tNId53qIivqzrk6GKSOt/RJEMUGR/kKZ
VYt9kZnbBcfja6Mt7lWnUG0n990XjvitONm4QIRSjQC9j675AzsCBWRAOkT2grcJ
5KqvP53IafK/2kaA5N4ZP2b97vBOkCNpBJYQOeXl5/v9GmvPcFwWL68k5TzpYn3y
HG6hVaAJMH/ixQDeNZL71bK/+DTACFaiDy64yDKoO1J/pff4X3qODLeLI+D0ElOB
qFshCnvlQzF0Ktm6O1KkXhDdNQwFVYnopadlwqu1lKTn3cgazaoAGffb12aulUBw
ddPO/64goF6EWZwxwP6wAh27ADSFNkWFEmkcyE85iu2lQjetpyYwBeEdoSxGm1Ai
meKUicy3wee+FIWlJ+uk/mizjA0N7bpPwjUIjUIuK1Q1p7VR9+pTNccC3VGT1PJq
1xxo+IeiThAMLqJjEGB7kONSRdUXzm4dH8PrPTwP96Fbn0PCAfAHg79G1hzkD3YP
Pw/gBwcvrKM1lWrjB1uYNKH2QopsKNNiX2R4v0izRcLc+iMJWxt0ZlEaCM5a7MKO
GMqgL7Satacc6IQOrmuA0BRPHygbdiv2PlsXNJfUlVKrKyB+5KswHzGqlIyERK+t
G82bofCl8RIJXACP88eNASSnYw+N9l84stRQfwE+VRoB4JSMnx+XmZxxy4oiSvNv
`protect END_PROTECTED
