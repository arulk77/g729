`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
2EBoZu9tBf8wFLCnm6xiM/afJQ5X9FSdTehY6hUuI5nlMeI/up7Wgi7xL0QEWfDn
2XBTM23ULXFQU5Ve1gUXIrJbBDFaHxFm0dVNtZI/SIgsREZNKdc8GdldarEyXbis
jzoRLWHDIm6OztNzueLD9TwwTSWuTKM4g+X/znVqkl93aaUDCFj5CGxBnaBCUK0L
cCpOW4P0ng55RgQ0HA6COQ==
`protect END_PROTECTED
