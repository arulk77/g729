`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ypEUOb3o6x2uHfRkAuQxBBmyXvcKNuMI2kcwih2dL4NNrQT7EM166NsAH6QDrmhk
XabRYvWfzHl0jzDBSvayWRjwsaaijAYc+HGVUJ22HHXXP+kzxpOhhHdfoZj7R/hp
4E9DqKNCIhVtbEwMq9XQpRTx1JiV+/WlBn2U0b13YUESLayC7JrFScdX5Fca5VHz
eUOYvMZN7mBgmN5pInWlY9fF3lmFoMsxO+I2AIx3RfKHbCsHO0vf6RYC1cZKt+2w
EGqUD8Yq7L8kUkKiGR8NAlVKZxnBRxCq2xyhLAJU2prFTpbPuK8fadyba8hxeOEy
Eys9I9eVSAW3MWRQJ7b0BjSZL6VU/CEpA9eQ9fAiktdkxiyY7YnqjpKifqc5NUK9
KXm63tSaKxfkyktfkL9lAxn3ro89hTzvXR+TpxtuP3/SNxdgoeKXf9GKpBesdNmk
N8vTLfUEQ2TvC8D/lOrxKTDYqrGp44oaJUgWTJBjOMzXTiG2noT7lBxRBv37fxIM
vPdJ5wYWrdCiwSixWnoq6Oxks0sXFJ0FNJGY8qnoovcQfhSl4+8E3Y7m/GBDLEE9
16tHU5ky6ti5m7BSXKxjHfduJtqKMkCRkUMAf1p4pwWK5oyiYOBWrn66ft4mQzrU
1DdjGFCOCG4CVxVctkIFjO4RTXMmqJSrP5KwUbyk+5jq+ZvpEIW2VJ82eexSx86S
u5KwxRvjYPXHqZWCTZ6wj4UCwbTTEPIKo8IMVlnsbtoR49KtCtpLInKcQLhQZ5Yh
3qrPVUktPOiIHGQVwY9IfnzvKaj/5TegJwfX24gjsu5RICaZcnl4UaRt/V9MR+PL
CLf257t7GTfMYBlY298ldp9gbbhy9QCQM9ZKUFHX6YBDX+7kDJoPA3zA6mw0qDpq
gXulzlHATdjXP++AY13N67Eu4qMRinWwHx694RNeS5RrHK0c9Cc23XIVHC413u5U
`protect END_PROTECTED
