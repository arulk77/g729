`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAaHa+G9suSfJBYZQpjU4lWVUIFZjn3sNbFJi9EcjMHg
EP4J/lZrsYBhtc3soDAe0aJ9iNCxW5nddhGg4a08pDDh21T40ohjyJxOFELpOS2E
fU2YDAnSY3VqHg35jkmBgjGfS7XsqGToEErBrmNtK+v2mhJBM+AV2D7kUhvYxXZt
jK9+6FWpKWGNA00vaJVvdM/n0fcCBllzIn1l0mhupAN8TePVdt75gDHcVlBuUOPL
`protect END_PROTECTED
