`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCVZ3DFWfBN1P8ZQiSraf+2PXq9Fwg3LqrsVy8Ua4HGo
6JvCdF8hHqXTL6EEeNpiWLG+AXBeE9IFEzJxllEdW4bTZ/5qMszq/H/2yOS/omnu
u0Hb/hsHyS88s5qaIOMS7OZ0bNWk8MG0IfhGsKBp05diGSxNKZucga9fJaWg9Ot/
u8ERh5YksWs6l5gRf3qEA4Is74ILUUq//uP3kb2l3ttBxhXhKhBJTbbq1Rdi289W
2ai6SZlfAcdqYz0uPq2J5HTqI+l04cAiW4mL1rcJU0/LWlWquP/QIV3jGD0DU0h2
ct8KRIfa1/avitFagB8wnjLRqmKQevW8ZHx/pTJu6VLs1q/layjhpHl9puOkNM+D
HRw1w8wWJbstiIPOJov0hyuaY5J2yYzOE30EJ6MDf6TmY6uIkutodwebkXDu4bbm
rt4pmXtYI7MU84u649r2e2zLQ/o+V2/ElkBMmGPZBBQc7RWQpvvh7l2DO66TZByr
HFhNI6BIX/sVW+vzxftp//HE1sYERhB5bIIkLxVsgvm8GzY27DcCdiiA9zatvCst
GDHPEFuPF4GHWP4SU4QzCI9RhsauRwJKE5iCr/afAKs=
`protect END_PROTECTED
