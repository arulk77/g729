`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGxQJtpRy21xY29UvXsNWzycVWxt0lkwZp/em4fu9Rt9
DhsJ3txHlrxiN85X85xTdD/iwaylTV9fj8Dqa6fnAOycW9PvLiaaHQZx4GOJkuDc
2u/hFrFynTWz52xLh02vrVeEcpO1o3V32ZMY9ik+LexwH/wh6S8Kd6Y3absAt+0F
ujF+nSwsD4Xk1dS/SPH5rmsMovUwK+H4GClw0ZHRZJyd1+RaYhM9bV5bAbVncNTM
TVxhm5XpemIPzmS1pvL8KLPkBlgcCi9kCJB0hjGHCSdTN4sO2l1ewnexX7jkSedn
SS3cBqgzosteyb4Wq0L5kkE7/aW921Iy4O2i+F8wR/GCGIM7aRljd3PKRt/8yl/D
RmWudQhcD7FINyGMRb1o3A==
`protect END_PROTECTED
