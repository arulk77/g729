`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
BXvYK7KyLxwlXC5XaXf8nVBvcZtBGZ3djCQvk9HPEYBD8TVe2dEcA8MhthmE6BVp
38CKwd13qYvDrXTv+e7LksoBl7vXFRxsbdIoxZBCrs5KVE/ZKGnc0PcwUs8Stb0e
OlHUSKADm99TfoIgbXzuSQb1b10X8u13eWM+GjYANffu0Qe4pZC94++ZlaapE40G
un6b0hZdbJCopDLLJtjNCQUtcyJtGU4JGWRwnayzDbG7dzGHA0Z0tFXb2uP3PcCQ
mG5u/fAJ0Iknwv8hqCnvaoX0iTlxmITA4RoX/f3EWt8=
`protect END_PROTECTED
