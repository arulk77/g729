`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
EBctdIPzkjW4yXesryi0jcNxcQmcTQspCTpVEeb9pzW9o7s3JiHxIfJPIWU/BiOi
8Gl4KVNxf9hO3lD0dAuNJeSLeE1RZTcc189uuXVPATDVP6oUxeMGJVctXVmgff7N
HIYpVVziOrKhfhd/DtnoU+XwZr4RuJRd04cW2z7IWwZAW6JJ9NsYt/bHv2ofXxym
JKXiKxWwSyQ9ENYYr4RuVAEGCTKeR31oIqPcR4pKGv7+c86zTULGYZIg/yrW5d+7
T38N4GAypAgHoG88P12VgEZmwhq/7kSqrqWgPf/q4rEZKhSR34WE04Woa/j9AI9v
l999TrFZXLhgmabN7LU119QStM+6BiMWvqMxCmkkav/Kdl6of7QDTmUgHLQnTefb
sIQiDwItvn4hYe3bwtNRnZLf3g9lVnrCzenjG8FJ4Oozu1/aXMIW6w18ltBcmqrv
cW7auDYsg68Q7bLrBKsCj+1lEH/4SMGvz/lDKdOv/6HvPw7xhELMUUiJtRagKvDg
y7cdGNpc33dZSQlb4nw3hK3tUZCmykyoWx1RJNIIxEIhhfZU7fcoSBt59Xm/ygkt
LP2fwHUlV5C57opWHDoejDGpKoT0uq4USS0Yiaz+7zC0lSNxLjtluFQJLym4rg5t
S+UAy6LXofQ3d3Eomm4PtVV07fu0gM4iyvYpixbiGX9WZbHX/DtXzJV9Bdy5EKhq
ua90yP6uNfAkL2ZJIhmtJHHvoCqDyIj0rlMJY7ihjAyicItluDKWLDq0QEJeMCUr
wwKk2083RZ2m51B+PxgvTIyKEX76C/K/Bc2cXfyVObN0hTz30pYIx7xZUj7zUcoy
QDflNBkhgE2Ejyh8MYYTW9nip07RMjoCvJ8WbTn1DVHE5oAGIRul5zsa3mmS62ck
KpumCchUJI+DrTzmgxtQGOWzAqxdy6BPjJNaD8gAUfVTbE1/0ziqxISUfBZV3C5V
GlIoilo6HmJUzKfdQV2+MqJpbINHLXf3Ay4fmP4kZFiMDjjsH3erRDqdwrGsHpre
J0Qk/e/aiA7ChtciV2X2oQzvfH/9TJKW3epN+znCwGPcpniV5rfuSas2fy3kbiFe
HLK7KicJ6eAxdAC6y09olkcs7bJRPFiyGsv8DvZqjj1oRHjlp8/FQsG6zY/yg8Nx
FLA53b3mbyuFhVXzMBexx0yQOU8RoSq+tccWIhj4z24zJ4U4M3Cy0JAfdSPKtdp2
nCwOMVqjC4wTFuJbE2Y989vu2JWScDbyA23NBjgZOers3l92jQDLdIYNrC1/jz6V
EbbLGeWJAioMSchRsXjViZuOu3onVcT0UFecWl3ReudNHGrvoAzFzZDXrjswExnt
AD/JHIkGfMOo/8C1dbNaU0SzP+8e5SlK434pIsgbFT7VCknElEpc9aKonmBdh0+l
TI8kTZPgPRUuTEEmsD1o4zOB2+W2gMCQA4XQHVsOopk=
`protect END_PROTECTED
