`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMEM3e9TQ+u+UrVC8NX21/meR3jIcxBvExSz/QeVdfS5
2UrwlFlWpcFbf1R6dBbih+ZsrqwLiGD8U2pLzdiPstg4i74tN1sx8nXLmNHQNqvn
b5jiEb2GAhpFEBc6/XNUlTyZbbGyIuTKx2VvqhM5aYeP40TtAul2By2HUK9hpOyX
08C+0I295S82aEAEcm1DGe7HCYPb9ltQns9bkPLKo6GcvF0csdU75sQFwLr1EHOb
bZAJ6oYe4m+2NB8n4NnKnnIYwsZre9meCi/bqwogTkCTclsGv7o/20W0NxTFpHF5
QyFwffeHlBBRtASUoBrWd0sPwidbMRATM+9fvYrOHkcIWOsCAtQ56darLUraPzHF
n3kYxiDf8gK7fvDRqteO6Q==
`protect END_PROTECTED
