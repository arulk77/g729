`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Eps588NCOp4uZvfjiURv7v/UCVA6hddSIpeqrthZOZzINN9+4cY/kdJYHDiUPM/f
JFFN4yUC8J8w0VxpnwCA5D8KFIJlFPG3A6EFNzMr3DoFhIW3RxebfYDZU40/BsIs
dfyNUq404qYq2nXRUSlwcwGBzx3/8TdHlfQAS6lEeHo2RONGbO8FSmCvo8kdRTn1
`protect END_PROTECTED
