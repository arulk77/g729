`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNTGmVovgvxg1BMyWi1lk3oxAjqaN0RytE5Kc/C4nOjm
fAv9V4VUxBIh3CHz6csBFBNEmVUrcwsbNg2jpfAzwuqONJ9L1JpXfYzmB1QeaObG
gKQUkzgGKpQjMoMLnzBjV+YKyQrgCpcoQdcN7kr0gif4PIFG+6FOKVSoTsGHS/57
yuClLZXfp8jONECTsVGKB6io0/ECp0cH8bwro543wk8SJc76Pv1F3CR/jYoZZemc
6hQdAqXSlK3il/wANT2LhnQ4npu/vyT6qrBLQ2CmnA0fNdlP+w0/A4I4j5RETOO7
zJBJZ3mfUQZ2T/xFUG122BgD6rttxKCs8MkLRsdGw85dnaC70zNBLh87HTlUbRIh
BEWcoNKPB4EBMBVyGdM4eP2D6KNw2i5SunskJ2Jw9Xuxe6ZE7Zvq2kUkx8TFkIFS
/dMOo3HrtHS3nR8GPSMZOa4itLzNAvwTeCcrPx+4sEtamcaxn36LK5YLGh6p24Et
`protect END_PROTECTED
