`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMotZ0JSRDV6KGtxrWttP0qHIWX4/5bCpBFqAM0FwJwI
RBTwnpwRiklW1zuWfUTgZ7x+0DAytYCxt8+XY2IOawkRtUQJss6P9GdY2YxpZALp
VfaDBj4TAXTlcyGgPU2KgEI8Q50iTWISBnoB5cAzr41F06Oi5ksWLZu5mUCscsJS
VGRmQPyjr/OhwXDIsFS2fjQyuu8o4iBGf5/S6Bf26jsxqazVZIVLcCGGFPJU4tcl
tICzruvXGzjmjyxxOyk9x6Diqqcq/nFT/vZV4LZsP2Hy/k78Lgz2XaoTCiuJcHSq
uZaNLHYBLY2jpIicae9K9qgUqvf9vsZEq8dFFJvbPgIVBStbYm+UAZFF9BvC2f6h
6Y+8HIomkiogOVSZJt7nOg==
`protect END_PROTECTED
