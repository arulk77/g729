`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveADxvW2KnWr+ztbS07LqGLzw5Pd5huQBBtSbTM1TxCNE
ubp+ssodc9rMkz7qOQLGnNHkKjr2F2zOlWQzJWJJAGKQKD3hkqRAYXpJrsXF2HZl
jwbYpa33zH36GoFVG5QZ+KpCn4i3divpMC80tEzJKWl/aihDwI5GzGyD4aJ5YsJ7
FLhOXVkxoDAf9iij3cI3gsm9ecpMc0d+fXqPVEHxWPcdINQtDINqwDY7QnBLs/r8
G5moqNGX7AZMRRCPwHAmXXwOS/o3Qb4VqSlVrOTrVPz8KirXPKG6E/vQEi6pCtlo
GrOErTPCcw1EjagJMdA4mSwOzUkMTsXflfcJ6q78TVW+pRmymaXI2NWMPHgc7G/p
fm1frYygK0C+GhZ/ebOYyk+6XR9Nh7yjzG2oS5dPPtQ8jOtFRed3gNQ18kzHPiru
i7mKAj2EikuaFLgxJm0em1xW7XCZfqV/X46hUiVkSwK+0ng3EnscZPjrBXrVD3ke
`protect END_PROTECTED
