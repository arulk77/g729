`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QwgQgMMwhGr2fbaHlpoXVhYiBWqg0qIv7A0TLFhnXgXoQWDlv68xziQUJip9DtTw
pNFqQF5RdmVXFomjpiuVpbcjOxbplsuVIZC+9CHPgzLAp8/SF0f2G2oEz6fTDDgw
IFkjlfLu0hIQKWQLTU4Z256QxyPtga03wdvuCNUXJTtwE5rZQrQlxi2i/3jh78RT
zuxXgyRXTCH3h+VwJZ45Cv0Q/3AAYq9DkmcvAHRegmvhK2hA0GcDMkHa2VNeeEZo
4jLg88TyfmnpoY7zRaUMhLqL6Hio1TJoCRoV4p9aWbjAyFpeniWoLm5NoLQHW3Rl
fgn4nWwV4jhV+eGejADjYSdGNEiOaMF5lqwBuquQuO8=
`protect END_PROTECTED
