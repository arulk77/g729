`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SR4uHaaS+jWZaun+bIaoeIQK7rSrqvzOv6oSI1X1cD7M
oZURWaZ43+cyCK9LxX4IanD5ofj4vNXtlLOxTFXSqsFtxQ39bvJxkJn2unP2es63
1RKsGy1f5Q/9WxAuOn1clT8mC61dzwKMRYr+VgpSAwgs7lFud++6SJa4EF9yO2sG
tLaLqJ+4YHzDEVoXL+LKVA25fAyMSxiRFEZAqkVZTT7Zb7h6/OwdbbDqpYyuK345
12GZxZyKLCsWOM2HalUf4nt2r/q/Ili00m8mIiX9R2BKkfQ2D0wr/iC/rH/Zw8wP
YTrb7jYC0Y6OD/6Qy9BbDh3vCc0va6RlXRD3H9mMOUHVu913+9D2gkf/4j5m/ZkS
/nbLGGe8JjesMLFcIKwrcAfYLs+Lk4p29cwIQAK29luNN4etfxMfc/2SrGA1wyaL
5x1IoPRtsftXiJWLS2a2PVQQAgKSWpcd9RLO2I8lb5pL2lxAYysFmJ6tP9rwmrWI
0Sop84SS4YaWCrcVwaTT4tsl5IiiOdmO/OBiDB0T5j7fDPLFMfsGAqXbgXfE/btM
TBUCvzMnRO/sF9ME/F0i0XruI3exePyvthO64D94f4hPZCMXc+Xk4spFaGLQ3mJg
qfPA+wlCWyBU+vAq6iqQWvgUOif9+EeTaUQ/2K/vRVJRcGiUTaiOg+umSfYdIDLM
bW7jgRyez9qtn+/JiYFvp0EzrQC1OxRXAm65dDym2aHvi/53pRekB5SjIhP1AVn4
Uf+FdRq5SE52URsSZIs8tL0h7hpTpcqjR8mehamLCiQI82hMsfWs8GGDQ/F+vscI
zfUBi1SzqAa5WTB196HdkX/AzCQrel10XqPiPFBoRupNiN86WYNx5+mhiRTY92+p
`protect END_PROTECTED
