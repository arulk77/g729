`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
X8CYn/7NKvUk7tYbmjvtBlI+cGUXvX6IKu/a5lZWXNCfHteG28cPP8H2g5AidqFM
0iOTRiQMUyv0GdDnKmSb5lNeEWISpRVSpCTSebEECJ5aSqeQsUD6hW0gzifl9I9U
vAo8eGQmUGJi/gjxz5I48qO5sxrGj/iSMnUWBoMhWxb/vX++AoIDDT4UE0EgLQnW
Yb1QlM4bMtju9ThSL9DCShOrdDqflHbZbEIEnGV19GMC9nhJOldLF9/Yd9e7RmRo
lDVj4v9ax2WD7yheBTwIn6fhElj4jWs2LBApgXVsWSE=
`protect END_PROTECTED
