`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHuXeQTrq+qb3YZX4xaZYze2BelTVxLofvMdMqbfw3WD
Qgh83ZHZuS65fq13R27FN+q6UFT0M/a9fCK4Q469uSKjPTIEvdO9J1Bv1q0aFRHp
bDHQFqT8WqCtweHNhNYWA0/G/YxhNL/fb04hwi9KMcrQ1DaPi2TXEJpfemBoBqcH
7nJRXnN4+5sscZMnGtk1ZRxVMkgPquLhkaK2vLOu7OH60TGkONUDItpSODh4DirS
N3VbZLJ3VmxsmwPpfxlttokj13kE76ZA4aLFnhpIIV9YczMHk5fJMfz93i4vlv13
lIzj1hHKEMpfB+cFknlPXZcptUNLZ50hcB+rm6UTNMm3TP/EQlhAra0EurPRS7KM
yL4hlp+xNIy/MhdM0o08Sxmb2ZoCR3VLM1jVzSc6t1/OHov//v+2EjiuLgPdg46L
fAm0+i1DAFLzKpa+ZO/QvxcMjm5dCSCcFLuQDkHqLM8ifXp0ejZ/24Y0tqN78LnT
y7GVj6cdWPkq9j6AFAb5+g==
`protect END_PROTECTED
