`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLJFuczyFzFbRmUOxspN9b9QTJF3dCPPDzncyixuGHX2
De3BPOOuXr5X1Nk810LT5wX/hoQTQ3ySzaVcVncyT4peFubrYiOOCyiVRqUWjVHr
edXMXzTU1XHtEUgJ9vYKx8de4oEzod/tRISTPuf8TVGs3cOYFQxshXQN5Hfrz07s
VI7Ktb7hFQcsd/7muZ/TNDnkIvM6vZFz7WKHmSsqt6ouWA1FenTNIcm1ruXIUa9d
uLoCqfXKTdXVhTIg2D8nG/wDEv8JTFZTWiO4qOPvSdBrEAxoMIUn4GmIBuLfPeab
EWmhRbqAn24/No2yMx+A4ycmmt4iwY/sywCWRll1sxg=
`protect END_PROTECTED
