`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN94ELj7Izn/kQHomVdjE8LQlHxf2FmG6ZoNrXmtwysdk
xQQdhT0F/qzSugAJC5BmOKVmX/pjx282cKit/A1cAHf94qJkowNDSMvgWcm7YZnU
ZvP1IfG6v8snFOKi71cv+zM8DYwgR4lh3v008oI83qNEaXrbYxyp1PpvchQPW32M
sXc+qMdGxS4XyOCvx7UM4l4607fp7n5cN3mJfnBjee7LhC2YYPHW+yWGyTeIFDJ6
Ov3DYYte8s8C00EMWHfGCfBpgalhwn1+Yt+TFCCC7DsYNXnAIvj2mvY0L2HQoHps
wg5XzKAzjdwrJf3JIG0ceCtwsWMt2kK4qeWVHtFFuvoIKhVnNLPPnokJ67dmOH3U
qETwOyCJRRRfbJG2PM2NIihlR0+ngtTevUbqvU6pRTfjqpm2eC2RlCPLRYjt9tQt
UZ/ytXVcafeC9GL/P2wm3y4Of0fpJMsMK1GJ8BCyCa4rktpDXr7Vl1YT4W4Xy4oc
cw8pQNz6l1wPUrCcwvD/fOov5+9IhkInAZjqcHWU6l85vYTLsfuFm89w0uJ8nX62
pOjdiJ11aq3JzWMzvlrGU/jHH8EhhrltISNdsuXJnaMejkm51wEy9v1v+G8Y+gjN
lyzclzt2yyao7fQJlXg5r2rYGIiLLseTLIwdqNpiFqXa2hS6cLkY8beKG+zE8CcC
498TtywEaDdSi7LMoz9kd0djoy+6IhUmkyIAuyFNMkiJQJMT84dY3XVoW0w9mnAP
6tvZ7Dmxfj0rQFoiwe4ioBZ0rYrerNgogfgQPVLgCWtVntQExjM0Hk5qrU7SKnzl
UfOLoh752dVdPjb9lYvy1uwBWPdBMdwIfT4gwWeEggR6IGGPP/D71V6POd+HKg0u
4Eo9M0UhXQw5rKvsokG5Vz0bEOzzr+JbeRqPRZZ7BqI1dQ5JDFbpmnluWmd/iTtr
KF1XgkVvkyw8XycduRp4FWP2rXPg+yIfEyurle2SrY0=
`protect END_PROTECTED
