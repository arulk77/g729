`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveIQu04jiD3Q4WTvINpPYKMHQ18mOUm8sCrTQNf38J+iN
i16l/jNdIlOi/j6iJCgZXCGO5L44ukEATNklPRykrsjgfESVNu3zzElZFDoxXMfq
T/WR6Sy2kJOKm2LqJaSWsLFmAHuObCB1TpZqU1R+NRs9zAQIJ32r40FicM9MZPkH
xM8m7q5Mk9Y0r0h0aX63wg89fW/nR0Ez1E1HfWf6qwgR7hVhTf4WKVLfHsPKuW4M
O7s763PUDn1cJupj9exw/D83nEjv/fQ0HSTG/4+UOqFQuonMEzKzc+ecInkcvPAg
tXVU05wT/VYnuYYLOO1T7rEoTHqAkEDpXIY6/voeuk4W7qeqtoHPKSUIsUUoG8kB
5f6duGJl3ofzbX5cLy/nAVl4Q5okH8S4L9B97JsqtBYE0hv1E7VkdJVBsuTtlXTt
OveYK/W+R1Ihry4up8eoKWhCSJjIYHJtYu2Udn7Yhso42HY70jp44jw8b7VDjNFN
mfMa3OcMOJMgtlMdoEfGE5Uh5n+27r52Nx+MaOcZf52SYV8jO+GbkiH55/s4G9MI
BDim0BTDYPdT8J4e97Ycrw==
`protect END_PROTECTED
