`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48mCTPVUxMvd1LUEPDR4D+Ia3qKvp3654/uaBBMt8RZh
UZc1PViLZMGDHLik9HeABq9XEMLT+fMW5h6QHSh+nOcc9h2ckP6lbftI+pAYJcdV
oMsX/5xMzf8RR5Tt+FgouAjeAX96xIKM2/7XmzWh2+Xy0CcJSMjVg2wFLbfZWhEK
Cthbsrm/BwwaLg8pY89oib7IGxq1EG/slV/dXrcrKL+Ie7zdtmTsqMH8yzfZkN4K
ntImEI+rFCwIzyFQpjP4KQVJTU2DAsNno0ktySraMDw=
`protect END_PROTECTED
