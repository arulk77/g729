`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveADh5wUU0onzawa/v/vNpZlZ+W/HrmoUx18m0a96hLwK
IOiXLxOVDoS4aJo5+TTONeo5I1LLdi987/M0+BPaXzDTOtrOobDMPqa/XQxlkbUC
s9xgtbPH4u8CPb/wUCPaZf6AqvCB6VaO3X4Gaf8fv6fpu6tKmL0zQ9XxK+zUF0L9
29o/2PiZm+YJIXF6YtDnSw==
`protect END_PROTECTED
