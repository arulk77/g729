`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
21Dtj1SaFImopq0kDo3edttVAMz7sEgAVmnNFHP3wMKYnXZKu6sL3hO6cw2bGKcz
MK2hA0UvFejHVdMiJbESEN46yD99iVFOyat9bOfcAxpsRjwsEd1EYZ5Wur3R/JOQ
D9okU5CIFGUAprRtCB4JWBVIxCZ3lTbM6/rx5gdS1HDidR41nFlkWfoMRUtKwuNx
vPYzaM9NVxrgYkJjIGoA6PtXorFCnpQrbUR+xSmIMUs1Vv+j5JMs+L/Bzi316ZA0
W8PfbbfYEsuJ5L01Cq9hDhTSHP2UqwsCxy4cUIEY+5PhNfOeLfG6T+rXMIIemYoS
SCOIKhB+/c+NsPsotkAHM54Nkz+n6RUQBI161W9nLS1PgoJDrNUbUFU79T3AuTyH
JFtjpaPnbKLngzVUmQyMzI7MGQTeNUD1ZXw5PduLKoJ68b3OZdoG6N9YXgHYicjf
ERGa007DczI4haeWoRx759M+UMdtBn9A/OlqWvXQ0l0dGGsUFlHr+E/fqjHG0Cmj
lO7PdsUMD4pMjs3L+zF1NQ6H42legUWPtKo2p2BGym4YL5bLWFcPPNPUA5tS6klm
68rjzVcuaEealG4WkRvx3NWb228Qto+ugMDmMI6UoiPhYwzrUBjFuDKFtXFgNeCl
vwEySXs0NBA8i3b2xo7x9KQUI8URwR4i8d8SQCVnofOaIEwdvMNvKwj0nuFJS0hg
nWh0uzPXgmMv9Gq3bz2yjYk2r9oVKB/++H7ExTL91HREqUCTw14XVxf0JJTJS7Md
y1W/V9w8A+ElFLQU/z8OlC4mDET2QTB4rca2wgB8+pBtdeGmc0j3Kqt/+h2c8XPd
/wAUU0g8pXgoQMRTc+wzxs2ppAOkl7G/8LER/oJ2kERPOLX6o623mBoBeWh0h4hI
ib9b18SAQ3+Lk96iFQSfsnA7UnQAfTMVewokRwxyHXJVws2opeCsIGHz5bHhkOGo
73BhzzB4daVwwanjmb43+qIyA5YlHTfVjJP1ilZ7TYpLkHreDlXuXI9XqFrrDTHc
Ln3Su1raJ67O0P0yNwhnf7rE1IjaJX60G7ytkRd36zc0xjERyYRJgcG4TScnJsj3
eRgI/n3eml0kHdsjLE16VKbjhzfu874mWvh2EOQoibt0x4KBrY6ewd2jiPVkRE9w
A0NidhCAjabhx6KKipDQY+9WcxgzRl4EGNY7TmPbk00FhjBEq3eLS8w/QhBKawEk
daZu3rjUYZ/2QcsPd75yRa3Ht1iJVuV3ZIy/DsD1skY3qYt5HwOhtxKpnaGjN0/L
V/I0RewrYbQWAfFmRvwFtXqOuGszjeAoVlLYKO9BR3B3EHPrKSZ71+klIgIT3CA0
E3aCYlEYOG3eQhwypK2MpatTZcnQ7G6plfP1br89h+JbHO3aVtsHWG8btPMhVfjE
2kbcUt6afTzV5kVvE0qhG0Sf4ZNBAd+oi8yQ8EyL81de4+/YQRClY3Xmw5jKRN0l
Ta3PzExggiOBVAj8bs8ARyWallOfKdaoALh2JWlIw5WZ4MRm5qaJO5MsvHd1VnQb
9sfXdOBK6gQn1uyUIAdTiN8vEl0xHIj9UlT18HQjYE0=
`protect END_PROTECTED
