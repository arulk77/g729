`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveI7KuO3fESfYHGYbpvXNcsqOwDkRQGLeOYSlbJDiiBGj
e/TjZXN4VuPdg+mrUCXcFTMcSAdjvicLO6o/ClpXxJDcBjSPoUqOjDQyIKQDViPl
9GM05qMETLhm1vYNBfy0hnHzgDzFU9lzrXQCRp+75LKwQ9XNsBPGe2mZfn9MPwhf
NdXU22WkVTd0qcs/ed0W8AGB6nN7C1Ow25ZfyDNPc44E1IejvJlY8tBj+s+krbJ4
`protect END_PROTECTED
