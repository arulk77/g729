`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveC8Yo24Wwa/jk+QsbSncUg/8MpdjlOSdM+1LjfFzsXJL
M6qwfqny4WvCqexIGW5gc3CKyYkfoN1E8LhB/5p8s9eSRSPl3A3LmgjOvSM1h75w
JKGYzo+suL2p+ZN/eSGvcM7SEpqhAvO8GS/fv2ivZzywvDbXzhB/G2EQh6ouU9GQ
O3bqwnm1P661G3/3ZjZvsrvMpsHLZcsvaXbeqUxzL9xM7EqQJWrYZFOhseJfTM1I
`protect END_PROTECTED
