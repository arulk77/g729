`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDdc61/f7r9WjgjjiibKq+794sfy3dGwSqdTqQ1JfhTE
46POfcE2agYSbMlZ8A7hQQsGMgCWMNBv+e82wzUGQ8j42bAyxJO70SUknAMKz/Nj
j/B9XUyBhjy3GZmAL6iIFutkc5r278I9o86KZYrw5xXAe99Q86AdBL+XgDFOPrrb
6ya4QoNUCkl26s0+bzcpFNYUK3AV0VEGj0BqChjqYC0stludsssKBoM/rKeqYxQr
l6VPr0/P14+HWqFQXDIWKxrqTpGnbNXHRmUKSjC9ayvaL6JhThBDG4NprvqZgGk+
bCifCSSB+jZsg2MTlfkS5SlQD7fSbGqXPix6AqaDqTnj5aCcBa5hRJR1laeiQq5s
`protect END_PROTECTED
