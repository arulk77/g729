`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4ywvb4VOy4rFJJfhNQ//I42acMLZ+B/ClKzZd5oaqBT0
UJEkfTIT5yW/Ghc9cIxieLok+LOx2uEX1v2yE2m/T4ilo/61MLQma9nNWAc5XXSE
jB5waGqKmDjBzKgOdoUPgfOoVqPKzuvPMdRDenX6GZ6vxKA43CBmZ8Fowt6Qy8rU
lOOUnSJc44dYSCWm0Jdk4TxkR4J3DuLY3VAap+kbp2Spq0ooq+i3DEKeOoDwpwtg
sVQGnNibacgSE1c2PnIAtvPn1ObRFERzHDWFETTCHm0=
`protect END_PROTECTED
