`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu42eYJVd1KskKkeGYNov9mBTdZMBhb7HH9pmfpzop1FdL
0GCKS9DTZOEos3YRjqtJbFT0ZuQhmW8Aep3xn1HenKD5TZfi7Lq3do4MYGgdHOHA
yBMkZDZVercfkLIQtfrByAMiZSLr2J5m2YBcIwtnaInW2+n9NEY5y407gwnuwqNX
EixCyyJvVNVStqGrdfmS3viUC0zZZtCdmFWSeNYF9A/GElSSwMykrsisIgw1llJi
DL7FdZBruOY85foPeIUKC+6TE0a/lvMZPb74LLBEd6Y6jXp6O/IzID7tYqDSQUin
kZIO/PGMQ32q2YRRax49mVcp9iHBbL8subgGwTdiIJtDcT509L2s5kaZX/YudpYv
enUcbCc9p815jwiedX1U6wkptmSBcO9QWOJ/au3biC1zB5DVw8QceXi/Jc2/D6/e
kCgEovwkrpcTNvdVlzCdjWwfgMWJ8C8Lcq33lCDZ5y/Gtqu82o1alLyaoE4a3Yj5
+q2ADg67jodaHjVKl6f6vzAi3w4pTDp0uyZ6haCGq1VdvsFSsPIFPBzM29NMQB3T
8ClynfR2AHVRrBp9AfM4sak1TNSANJ66XYHc1VcreE+e2fENgSz/iN8DEwj80Glr
0k2x3THTgYkwKmNmmkPsLfifv/J4fpPomDfYG+mhs3vHDkNNr3v7I1Mu1K/uW9jw
IEJ1fOGRXxQ+NwG12duFy9cA3pxPlvcamXKNpIUkK+oMoRPEM70trKBgJb7JhAl0
2KNL088K3oy5bHaiPpYLMSZmxneJItBE6tx77guUE44E47Wj7Wug5quEHjR8ybED
UBf4wNMaTYd6Zwn4J+cLle7xowjhmeZm4azdxMVtJHAUNUVgC1l2ushnVqdBETbX
fqFXUzx1dCcw5fElqhwVNBIKIuwC7/LjIa36k8PBfuV/Hp7jZDRZXjXMGEstSwUt
9FNA2btq0ntwLUZ9D6DT7usXrmpb56V6G5eqv3qCik2rYciH1UhgA+0TRXcM0mTz
I1DKV5s3K8+7KHgJM9hf57PadkQgV4CcksxPOZmGtZGK1RmbxALzGi/rmrGK3sz7
YI/KvhFF9ZzhqH9GQnKfmw==
`protect END_PROTECTED
