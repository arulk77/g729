`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGsBGQ9hQdf908YFMsK+glUyn+Cn4cIdVDCI0O7eZPuB
PVQ4A9ASkWaC6BQ1hwrhkK4qaVAtLolnZ3SnNybf8O2+i+Y/f4lxd6KCE4GR+rDp
onoqWX+pTqHAiT9vF2pHL+YrKcsTIniCCoR8DKCaPf2PiftOWu8upwcKlT9b6jJr
PhAnFHHnWMrl3ItXrXm3TWY/OUOQGzcAhNZ3EJ8Ht8TGiVLUWWuuhu5q8TcKXRfD
oS2RirUolhQRqq+U+9s65M4muq+Iuq/89LbylXHWZXfrDbBYZ3wpUhCb5vqZCvMH
QqizghuuUMaC/8izzeOhG5UDMQBhJj65+US4zuVUwqz16zWDA1Uve7A8uJ3NfAfT
c69VCf3Tm0qHtioz1SXjIV3JSZDCpe/Z4sl1Rsa99HXH16yps8+/KzJUBQ1NynNH
wbZFaY4+TOHZyx+tUKbHSEIs1ngyRXNlAglR8FTkcIgEb/AvfAxzKZ36ab0/FVir
mQnXxeS+43+rCahWtbxnOm7oBe3y4sjPW7WqpduDYPLt6LakCdBuYuOSkyNW6KNS
`protect END_PROTECTED
