`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAaafGt3ElVibAxoaQl9NW0SW0Xi3oLpQmwRY3f9YMinh
rFFhy3D6z1oUSMVqOcUJLeTy3jrL51whrs0/iljBCzNnCadTMePiBjXRrjuIU+TY
lBOlc4sUx5hrdbiRihFnd6HVDfj75qRdIQuJuMuqp34F9YQWgqd017lPYNKzWTez
uEykZrHWk6WiUyVORQXhsz04ZsK+kDT+eb7GOsmTbotBSGe14fWfZ7KahKllRe77
sN9K5rNa0Zr3l1VdmLH5ezwlXig/S9DHKf/6Vu/I8qIK8IozoIUGbAEIzeoNsVSI
Ob7dXsgWz4yoECbwrMR1TT3I8bHFfYrCFHSOhuKX3QjLg6ek7Nck8nTAYDGDieih
NnjCXAxdaoYY4+c43BFTPyY1neFhqbLxA2mszco6V29GLBOXQm2nMuuFJfDW7yhD
Cs9iDxFELSxRsdEaoAEjuC2ROcAdYh1tLw3v2tkSiuQ9TLu4CYuTup4djDVD+GYf
GR8hR314cIRGhL9vWTTdDdZtsIjnGbb2pONcz8t3/ncGOUwKw9r5IG27dMIfkqWy
DJqTMYvidQcurSfIDuREkWvq01Hzt05+iEdqZgMIqqUTjpNVbkeMGWHu7GZhHPuz
o7kyMT5RGg1NCcfEKHE5nVJqEA2BxZ9Yvf7MhL2/rBF2Bv84JfsB6b3KCncJn4wK
8RvNkueBCWi9bIyUCSy2Ozo7Vyeb++kSQ3DikvSAC5u11nb9/0aNYdpJkiVJrA+T
y1ING1UnpaRpTy4HQsTO4VGqw1ZF4zNVQGIMoImGJD+BoaPYR5iG+GWeFoPQApJW
IDtBXcXWraHfMYzRlTVlTXsPATZfkXoD2egsLEMO8VieASh9rtLu2kwVk/qKxshb
vt1hUynGqdCb2s//1dbY31h47E3Wzh3U2anHcy8yO0wh3jHNyZ+GAgpqa/mP50iR
`protect END_PROTECTED
