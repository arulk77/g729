`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
EqRHYpY1m64wZi6VSUCEAE3jcYARBim0oo04ND+10kQ59oUZrHMylsV/bjc5KimG
9sqneLOl4biqGm0/b7KFjBYeslqg1UKRdzCGOz9K1EH4Xsl0DAc7KSteWDljCHFi
1jU+0CbTqzk2guAZgnhZYTvJjE3Psj4Hl3yRNqY1UAJiaMGj0k78oMFD7VHQ17lF
kvWWiwXQR+PobrpLN8IS4shPDQDcx2+SvZe5NnteF0PLJXaVTr955QINd04mLPOa
UdULH5OuGQ5/t4+37otz4ebiQghFhqaK/4gv5gi6FlC8dhoI0Fc6bf5fQhqzXN44
D0oU08JjuVFdOkISYmGxcCg23atjjvw6l47elmIH5eQjRGKSbHNrfUzrFKUP2kki
2VQDAM8kbEuVInC86SENR9YRZoO0r2dpXkHYDVlRcAGfCPU4axZAbJTHJSVnE4JC
9yMq0qnNfBWgmj/CJaqA84TBchLZr43KM0qgLKo5pzNY7LA8MA3tUvCy2GuUPpgE
Ze9WTaOqDbtKzhPXZdfQmrW0YQ96z/82kYdwglGn2v9jzFcNfDf9kSJ6OWRXwhlh
kM5B2+hVI0N27YOBiuj7mA0Cjf+7lhmOgxdA6dF6RkTJBWoZyYnLpQYR2lsRnyT9
zbAfrbbjpG7y5iZJb9yiUnegSAPETZ5QhE+OalXBy27JMgg5T5hTqp7xw7vrr+p0
el3CXz1uwjUP66Cr3Fxgr0XDY7j9TNOKqp4VfrjIEJUPcsokX8UMWok7UrXUeYiS
tgwFMTmPYcWqCVrlNM3UC0yZO7yXIKsWGRIdVPsfXID2uN6OWW2Hrj+jQI/rT1kl
zW3s9IrYNaujjsNAqQ0DScw5sgrz3b5exrzEkLsq58Nnh80Lafx584EfwLavYumx
qpLF/fdE0xBMotVn7lPyP6i7616vB6JYbfeytVhy/l6fIh///lqb+WnitbBa48KK
H+IjD3Dhl77sewLYdgUEYQ==
`protect END_PROTECTED
