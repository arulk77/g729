`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAFy0t2/zOMMfMOnU4b/cg7E/QDIMKL5xmIfYIDwFpw7
zxDEZWTW4UIYErSqz+tUAYE9Lj/5vFKL5059BNx7KLIbB8+NIFcC9KWHR8pfo+r3
D2ER6xp8c01+bVIJqtNwokpuUNDEhIAMNjx2zw7ShFAy5Ko6wA8ary7Lweif7t/G
8U7YhyPdCFux1wwUpwLUz9jqrUrOGaEggHeSgegrx6gT9gIq82ncCZsC/Ppjlar1
gq6NTgDGvnvpjevPeDlKMJNlONfGvoytTu9IWw/QfPwMuvkjx4wO4tihDzYDi94U
6481kS0OYlpXMCWmxzKqHg==
`protect END_PROTECTED
