`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
qPTE9Dgsj87/jzijXP3VNM1bP7+XqTfsF/6m416qaIBdmk+mYuwgUZGibCLpHIP5
MTZWWKQGBMQncufHBzhM8/8naGd5euONqAp7cjWEIRse2bASnM0DzZCdqlalXng3
r0SDeqgD1wjlPwjKDPeOYWp15ZaKgKrnhOeKKv57ENBff76PUC1KrR11KxHlJ92f
ss1jv1Gv/sXIZn0f+UvE7x4+j+xff/W3QnZCjMTAzbSGDupsnvXGf+pv2jD/hAVj
2piCvF27nGg6Q2A/d4m8zorp10hKRYHUQeoWJ4AAgXEEx9nNPJQY3iZTpLe2iaMi
T4CpZeo7COAcCD5DfCaYDGqzgaSCe8Jlm39wIbbK3D3BPospK4h2KTftu3U8RpS3
e0Zjro2OgraY4fArtIgSHmwAp5YAGoixGLVHVx5Yu338lqea1MKLWOfz+2jT6dDO
Bl7FqYTANzazSk6yHTmhuDTkcGLIPC3N1pFnvHm18Xw3YCMyTxazW3y/te9MnZLc
xFPzgD+I0iaWfwJ3gn4co12Mz77deECMQm7VvWrJaz54YPwXebjrIlyx6cdsuXkf
0I+JbnRj37hf3+8H4Qo904zkkG3MxRY9Xm4V4g242iQ=
`protect END_PROTECTED
