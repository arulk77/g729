`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
inQM6GWMhI9M79+cG1wxkaqirvf7eRwlov/dKMOD3MdJTaFb7OE/0B0FaDcHfi3l
kZOrDo1gYRt38L8JB8qlHyRfSN9HK0xaGrkbIADpFy2zW0humAk+u8Ea/fEep7s/
6ZzbvrNgJuy6Qg6MQTtqt07/HMlay7UAkMd0/j+3YdCDdaSBJ4UpSxw7R8OfFTkH
LRS6nUioH6mkHNisjBtAnTxSbO0s1xC4sk7ICdI9vkEspIv4hWHwqfqaAIXV6Jk4
mc/fZ9+VY5f3vjmUGI3j2st3EeA6rC9R8vaMRzyPx6I8ESWJc5FKNF17bjOv1FoE
Uh/VC9JAlrlStyLkWzomNg2sRFG8Tunca4zJubXJbW4K+OAnqPHJGvScF/O5wzVE
2nDKOsq4EGf7r9+KYuF0CqEnPpvnIL62AdscdUrDGvu+iUFBn3XipQ1cHByw0uH9
uEqJmub7iNSvqKgrP4vGH3+HLbYVun1koNQjib4aLLI9o8A9vtkAfCl3Z8VSufiD
PG6v57hPmv2NvoOv9Nz2zmO5itGCWS858tWAdaMEXzybdDNblmp+6GzL9lR+0fNs
mk0mNPHGZT5kvgsAXQpE0/oF1CVkBCiPm9YBisi3yi+SJJANZ5yha5nks3LU48PI
ieSKdo82G9iNKK8dn+GxpfAM+lg1Gr9R1m74Bn0afl+1pcxY0/Y3Hrz8dUM22xk8
DDKXajzLC8lATIZFoD9QG0JKIiHC6d5ebHqwJeM24he8gmi73k7vPBVtk5tNWJ3H
Lwv8jjvJPuhwMnNcJRdK/4qDY90aBhqbfq8LSfKDQL3C5zgNgkRnY0++Oqp6TADx
O89ji0NUwgjYTpPxyyiK4qzU5DGxMMjCfoqUMn328xiz2lQACMK6SkQoPW3s/LBT
jtOK9jr4CDn6srdjfKJpT5/DEnVulUUr4ffGWNB89tMBAK4hEktSd+uKTB92XC6T
OQpCQYXDaIEbSt6sDVWMa6oVo92k7d5C7GPmzfB6JIPuvVDT20ejosEaYPiyiWV5
Zxmsw0cAEb5X1rD2hwI1vihm/sCZUKtyOuqV8nlozBl7k34nXnNkpHuCaJwfRvgj
exq2A0m9IiYroXmBXFOcgOiY4WZPyFNvRJ7IZtfw/wQJUaYy3wYidJPFE1r3yLYH
xY5A38MhT/4lWNtKJLBSc30weF0MITTll2a2nbyu0IQTlYF9Qvef2WSYLT/b3L4/
uTdVR2e/ZBxxTzJZBHTC2hsv7itWGPlZuRNTzzRl2c0vKQKzx311pwv4EAmO7QFh
n3YbLdE6REmecb9qrRVtbK74TyMd3YiW5r33U1+4X68awl/f4p3abQ6hEsAn5MV6
fSEJFCcM8j1ynydamtnpM+V4EOos+H9gZbdIy8BURSWuyuHKQQ2z6TAiVPSpzJ1w
9XOWH+miNSlaujswPN6LjmlzMAJN8ZFJLay1RvTrMEhsL4MNfUcAr9Qz8rYNJiHz
ywjV2XShlhUQ5IZL4u4Tq/D5QAZxbgx3vM8c7nRbXgx8yK3XKIowXdZUdUx0JXFY
ADkOENqMG40CzvZZxrmRXcIkV/MRRUMdfwKGI/SAd6Byr1+MsRzW9iJc2wMFoN1E
i0E92hI6mhChQXer8Yt707vU3E/cZ14c49CaShlNX7qTdwqt0rVVzi2YqkUaBGkf
hqj9E4VTOYil/etEgJeUy1GUFhAFPuGLyoZtlINPp4uQ4F4i6mFUUacTkIf9y2Py
RR6FaAS7WbzubjsTA4lNp72S0hcstAxPqYHcKmCYsHkDFWYNYA8ZdigguGt6fzwm
0CzzuYAQgTxhsia6JQpjAbRMMzWdiY9JzsUT6ObYQke6sRR9jQxedjM15QkdZz2N
0L8uYQFYdagTf9R7zuEgSKWe1OkW1IiUvYCS7DhaZV+TzlFbOtdWbK4FkoXxPrkF
5BoluBojziIq4gKW7DYw6qAwgKSTO7zvrH1sKIonHQpWMWS3XTpmFzlapJnvcvYj
oArQ1PeA41LUQ2RGnqlvKi2XXEV4uM6PxQ8V+BIr0CHujD7pOsuzgiKhXf83YneS
TevmbKOGPolMDIjLC7GvGVwGVPqxH+MUdDAxfcPx+83CFL4jc4ApHv1Nfobs9o0q
pdrg2ddvcysB2/F7j5Nzti/Gn5vUhWDNus2+Tt88pCf5UzJbZ3HhgQ7lL+KBPqxA
ivVRtqtnQRGl5ExDThdxVPNK9qAWGky9d48WlnvcQClN8ZS2PiYpjAawndCGtVF+
P9bs05PCcHuuzo8DAMYJ5QLM0Nut4WURTCbh8qO3BbeHU4DbuQKpP7Au35J7PJ7o
/QtvUMnk8PyH/aGYM/J745zyStpojBf038ZasslbGeSzCOz2G7JB4/UoTFHRD/48
1IrGctL8CJoCR8deYNXRXnFLlRLIiWLbb9dQdKoYNuncB8slKA2lTnRDusKsgn/F
s2X/PHwHZUS2XQCbiGCERk/TKvGOGwHiHcU43+lW4ckY3Mxb6Ak9bqbWgmVkVySO
SCjwukfaO9lXIVTxonoXXSrTXqJ41WgZtcg6uzj+f2ib6Czzp1mLPL7yTflF15qZ
N2GipgcAapiTkZgnXwgOic/770PBXW61aS04lgtd1tIiVZMP625+VWwHRv3uXA3v
REpO/f84KlN3G67Griij2gytBTS+lgdkJU5uN59gsafQXtu2GS4g0X6dSolPkAjb
4eiRMgkN7FtsAwvHfSxHSlHPwOeVOOB3cLJJjMjNfZFWOm6yh8utPEp5aVX+7GtZ
mf0M1jTU/fWha4bEftelqvNd9ShhzQiZx2F4hRLOQIAFwr30L+rmLD5YdD98Xz0t
lSDVap0dlEGK4y1yF+U55eztH5UDQdcsqZ3RyqHGTkXQKOeVJqzdwiJFXtOLnvM4
ULbkeim1sWMvT223W7faqvfT4U2/PHfUrCUKGqQ0ll9qAi9c/mjwkDIoYIyhv3Hp
zPWVdJYFnla4pIItVDjHkrFCrU3+dL1mySERpDIOn5mUkXmvFRNg/kZgEiFO2nq2
oMT52CTfoKchogWqw/fx1yj9jzoKOIfWkRdLfJImyccSfRq2eOKZC/9KKElCI2wc
OYmkYDXWA13Q3xlu9Q3zmsY3QLempln8I46AagY2+WlFcz7OBG1GsyfmUv/vcZzZ
vQz7N+a+TXbLGub6T+y2DdZ660S9K7NKe/k/mssApKevG2fnx4NrzG2lrHEetMQS
QJHFn6qYXPnsl+mBSPf4Q8Nw0IZ3NuCvwlmhR3J87Bijm1RL0szLpPBEXtWRNC+b
VMZn0kqhnCKb6jkH4GSa7rEOfkHlaApqgOMJliSkVt51qiWhqOSMNc+3X35r5Wmy
8G6KmS7739AG8mcrXkeWvG2YhV9BD3VhOOgz9FZ9OlGLGFtbw31EyypJICnfQn4v
5sQmFOmRh50W02pUAQUKhfjDmvJ4Zc83RxEImGWHSwOHMiVAnHejZ7yEbtrO25gz
Alt7xFTdQNwM/rh4e1irMKlbI5qGgp7v0oYm/7cclK29eAyRpEG6bXBxpeJCeLC/
cbJ+EQewcbolwwWmfsUlirbm6LbL/rNrjIcFcgRDHGsWHT6Fd9hRr8+4LrQicBNa
26oGRBWprbgNdrDn7PA20P3z/WJbPCwlRkqf3oHnrrwwxpnJghjYRccNB/VTCuQg
9Ca1YKwBjxDsJlncnYbOWIsQ5I/SkI3b1/vUbnbK5M/MGuvW3qc9mzF76K4LKNpQ
jAHN7Zz8Ii9EOUsFoZhhR5ajjcqFkddu2R+Fheqnzb6yWO5aZP8Aq2MJuI7D3lSO
7ru/SrtZzMyTxK1rU37tOudlb1MXQDCbipU/TsOOgqaGO+Tbdfa1LV86MI9vw1jS
6kWv49buLJrIfNnwojIDZzvucXnjB0XCRNt7cQBMw+jI+kVMtlL07d8xRsr/qYxN
/CwKdaqdQoJNiwD60YM0SQFWSPnj7HoNS/BATtXLlYjUmNzdIw2wrzRubWPVfCEi
VXvucYmUT6/v910CuL+zsgkajwr3EYtIfjvhVJ7GfTPQJDIqifXBckYZ2CHRbh3T
6CteSVXdD+eh3hoCm+pF4GJxniaPhF0+77pLDWa6/yTra8OQBApKTIGLBWXUFjlV
X1KjcWno4lEwd7COQOKG8wGKelHAE53f8YWv/AUqbzgFC9ms/EfOtGyEYcnhmu1X
4ScHTCX9ZcThX6ocBQiAx0oiOv+dxzehuRw7t/rpVJqUBH3LsD7fDtXQaxxseEJR
vVkXxaP2Nch2rV8X6trw2r2usZzbnIuj9vTFdcbMaQxyRsVQlfkKsW/tDjFW4qP3
LOIgyBWLK73HRld4RJ4G3fygXQMgOMdtYFJUphM661vt0kKmmxSWkoGX2zb+4Etw
KbFuupUfS5PSs+ojNNEIlf2hsmqHSYxq7+10rJs/NOizvpa+K8oWGJFRfMZ0v253
1lGxX1tUfrYpmdimE/cQbGxxlm2dEYT77bSilYh69IczEpX7l4ajZYLsdnpx5YZG
NhPcLutlElLjl/J2h4YkklyP/K1NF0u6ZAVqBub8yugKGYYHjvju7XKua2ZqWb80
mwKB83e7tsbUaWrYZbdw9u2yVnOXaRGPiEW7SXT2ZSabNxgkl5ZLgDWHh8phzDC0
EQrGmdOZW8eQgAY1t82iDud9mC5Nk+05zlliKut3UCdmMDbcXkvyCqbeSYak3v34
+DUSaeOqiW58qiR+Nz4iYdHgwnCvrEFhFLpWorpfmpens26GP3OY+aN82ngjIxX9
K9ocB7JYY8iqps+xxzqjzAr8sk9/rOURdlsKI7Oo6g/DUkWEG33xCxrKh7cjz0hx
6DUBEeUWMk5VFyk4Wiaa/QUayL4V3m6EufIkf7QfTDa6MLoluD+j7vm0Flvt+bUS
hmwlwXOeOhfOY6l3KSj84prQ4GK308v0674/KdsjRtD9HHxL4LIFIP9CyP8YpQwJ
wXPfguKACsnHTp6AvLOxRUntY/DMGiwdKQ6/cgII30tgjxZjpzwBn0xmXENj/uQc
rsNyT9aQ6DbbtjwBYY03E9/ui6kSleqvUSWX+9+d8xeo4WsNG+qlwK9SvCX89mTC
8UNY0Cr3vPOXowHinT28bKxG74+V9Ujtqg8CBb24KARbIo7QQ+ij3p7bbfexyWKZ
NbuyFsBwDqrUNee8CA/GOGMAsRenOfrj6Wl+wi+i7JDW5KJLCjlcife2PfwRE+2w
S/XaMA0zxwG7J3j7Ew0EhH+335mrAOmTn81g3f3Z/6JbMUa62cOWadjNIaOBkqV3
T+IoBGZkifZ4ZLubaZ5x3hJ5l6HREhiJZycW1VVS1BU=
`protect END_PROTECTED
