`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
V5vbPYVtt3lvFGAdx6tzZ2NtAbRr4XOy+qGgSRbG7BiVcZ/qlsx8N4baa6rV7+WU
n/q7t0WNCZmSIvUr8QXO9HbSwgOA3D0neVpvIWwxpWlmwUVtITuw3RWDCOSEQOSP
0WNicCWoKFcZovUXYJFzZ9y4T6/VYsTiVbdrq76Y38B0mxLwQbm0QHdJBCB3+KvM
+B8LoJNYY1tjcY2aH/fkmGWKj4+ELkIhvbXSErgV+Jc2kALEO0lQUkS+UFZp2g59
RTdB15CO78wmH20vEwKIvdiV68Cq02E3titIHTEGtGiNnY0Sg3aux4TPv5U86dMA
C5ryjRjM6mf4HBtdUz/Y2CKwhA1m8LOeWkaHrxpUiMFiYL2fWtp8syDRzePyrf2R
v2Mxz3MJ99UXMnBx4UXKQOiyFVStcjY811v/BlNbvGpc5Yb+cbY68Sa3GNXy4IFN
Bz1uN72fsCOZAQorYY72Rhl7jvN1zEeNZhQjXJsGivE=
`protect END_PROTECTED
