`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aaeRI5opGNfuyVzRnOTfmja1yF0xLgLz6EbT1iLdwz9T
4mLb/XU8H+FFD7WZd5kuom3Y6ALxcbZg3C6EKxFg0yidXRW5BL54s/falYw8GBHm
jFv4HeWBLHuKuwqqbLrVZTp5sMjlTC7ZHN+Ob7qEhJyeCg77DZTuCEC1NZ6GIAHB
d5t3Mar6KaN2+ys8nbi7uckFeLPfHXF7n4PMv2rBO5jZocNE6GBx2UOgfd7JsGDf
FT29tiGSzCxd4kj0n44nRDEt6BujrTZtSSHdaJ4S+6aDgmIY9nntENDcadqLP9Ks
ym+Cx/fCKVviCZZG4R2pRiTkBesX0h9n9KuyRxT9TvHhdCJMf6g81uyRmDyrKvaD
DdHIgh7HzjNfQ2N5KCPMmJyxPu8sFNzgoT/Gn3vsAaeXk1PzWz8EZDl/d0q23kQY
zmDTWZhjnsVR2ym8AlZupjtlYJ7U2VaruLxewr1OXeBr9vhAW7cfBS2TVICdrzIx
8Hto+i1jGAwYXZADP1ob+vI0/pQHdS/fgY48DjTic3Re6rwmw8iAw0jEwSz86XTQ
QZNs/nZG1WZgQ4jE8NyTdmZyNuUuKaY+l50WPDkosnSoKOJYuajFx/nvOZ/bOCKP
swEiMqPbbdth9i5UpAxjqqbzjNK5+e8s+/q/g800Ra75bvDYqzZBKV0nNQGUqwFl
Ju1cTfYuntsChMmsNt3oFCg+fIX+UmWkEc/Ya0YG6ifQBmi1Um+a1dIT+33h/sUP
O+LqQr776y39APLyNu1wS/JegiW5VS7udwQUmBfOZPW6AO8sLCbRGIC4/u0SDTHy
iPmc3wNtk4xYJZcA3zSc6e1CSrvrUTY+xxNQm9YxjMWqjWD0stJRwpzD7sNGrd5y
sX1a5WAF2dgHuepgiwCMGCH0rv7HtmytIHIcEONHehh9bs1H5Z8dWL39O3sgqP7D
zq9WZaITONCQcBjFN7fqBA3lfJtazna40BMSgdwYUbAqCPVoTtsdeuNkhF6woKfX
j454yBbsptxIAEdbiLiZBcZp/iCTE+yt92kvcvJAaRLtcGNtBI05ATkxhoNG/ykN
p0aSAND149cvJdEkyZL8QoPnT5za8hc38KLM1gkZXEN6KvLXq7nNK7Z7GFE0cO+A
I9BqYvyFv+6ITl4K8fqIKE9Pffcv89yOnyYE/xBtDVaCkjDGexDSVxyG+MJRYMS6
7ISmzRK96jigA2bQwuMGi8cFmKY57n6A1PLM2lKxi3hVsRLJXn+iONWEziYPkl8R
VJYJCA0b8Y73C0mGwq0SKAb5wlSngV/49Rgq0+WAtEAOccbgdmkA3R1mb5LYHwvG
JtAfR8czIjsOF43T4NR1tR51va6fZWCQ+99+BgJyOSa/jVsaQvSTSyWm6j1q8k5a
t9Od+ZLB2TrB493kpTcQy6RROntwGA9zqNZqN65T5W/PXMRO0ZxwWJ/hGBxbYy5K
Tpc9hwh5PseLjxgJZTB/nESlTPP28MgW18CNwNBpbYyKhkiNWITdgbTRxRFtajxr
aDlJUPkrKa3pRZ1I/AkMm8yityzrlMeusQCpy4hdVGV7ja8MD0nEprOTjACZuuLf
BFGaorCtqYIz4DyTrXe8vzOIzPDgFDWpSTJM3WNn0VFktTIRJPZJxdthgk5086QY
IUTkwGlp9JXAqwyYlFPqg76pv1YmiGPJVZOUAmgdrOxoV8AZPDEYPJv895JmMN58
/yGS6rVDr3qO0GIGtqsNhrB12eroN0YhpCCcldDjtqejt2VhcmThk/3ADhXOgDXx
t+e2u9SsyxsGHluKNmCIii70neXftIRvivXS8T4bdH/gQTmLCmRvTxlAdEmTgU8F
W44iYAC3LWypdzRHxKALPZlVKgBbb8ozMzTL1PkYrW0F0u6rgQQ5Dto+mRbqeIyZ
EyXFWG95djlKyPzX7ADshYrXZcoxbvjVygX5YrM/Xqcs5Oref7qFtOwdqWUiLtbh
6U1Ym8zCN75FvWvBLoK8f7TTDXlObJXZWbKj2atOSEbzo5WiMLb9PZw0vpi79Th1
CGuQJLpkUWn+qbmEasBIi2A+eJMThxHsPfFyMu4kWKjOH/eyfYZZdTlaoO8KCyx5
g70WnpFyBHsZuH4uW3dEK5PpnTdaEa0AUFOaMDQKb4XaSp+IrrbK9B+5gg7fS+Sc
K7lRA09Pv88qOAVQHKfVgD+A7PZSDf5oSYgGPbMC4r+zXOxJ52UnO7b8eUgq8LeG
C37UsiHACJXPjRvhlxFKL2rSAQ2LbRJVr2dRkj6QA0fe3vK/gDfk9JrACAqjlL+g
lf7SdN1uH5VAYoGEZfIbh6h9vd161FLk0vXs0F07Pa2YNgfC3gYPjiC03GPleuYg
LviZhGQ1sjBGHARmnsTNtiLMOoi6RB8A0A4UL50NHvYA0ZiWBVhubRdi+bvykZDy
6XLWyVFeqB0SpoS8M0WMEOY3aGYnncSM23Glj+DgVLJ8H5JKQ84Gs3JpCEdFLgn2
EI+FGC1BS5WoISmE/7QmsLATLp/QfSI8st6mGlNd8IlQcCOApCFsPLExTPk85p6a
uEMM0i50w+9wPKo8/3HeawY2H+OgNes0KkGf38N7po5BZFqqbkjCiGPtn7o4Vw/q
JxJzzG4UfnBeUqA0RmCAT7h8v9Gw7EKlOgMDlwzNL52Hc9jOayfqX97tBcELSFsl
0RGipVRgsCfIi86jVDd+7vblIlq9wQovKOPFqNz+LR6AuJF80ErJ4toFmvBvdAvF
9JAt6NnQLX5Gy0G5SGdjY1FdK0Zj/iEa7qLAw5pBhjhkDpPuytPy8fxSyUYCMZyi
ASr+W6+06LsSUqUTrW71tVWRXwQf+jUmg7lsmD2zEDfy5tpQLSQb3S+JY8Orunnr
26gySkhsHowXbGMY+d40HWI6LUC39V2iWYlKpGf7LazJkMotCP6yrmkJEz869Y8x
2/iN4GyH5N9czEd08yYbg1tuigvosyfcDeR8+6mOY+Zn0yUr9/ABnuhji/uJbVzc
bxnRDz7s2wEjKTU4ObdBcFrP4OEehs8ibi0WTjFcjRInHRi1WFmsn2A8FNtKU6m0
Qvfd11YA0u+ZVlr31eC6CGLgj067G0qKrWT5UOiyu0vNcPcIb1dty3o4/5cjIy28
TqCXSCjep5RksaWalk2UqSPsvncs/4w/opFFrzctqPWOBxBdwq/mwHyhuA87xU0E
VKvT6QhRyGOAETpsnfjgAxe9aRBOB5flaJhiDkkagyJLtWUQAII/HEIY4ED4ta52
uBSjKdcRxn23UiJuJfV8UxPWRzfVG3bujkB+tjNPJbLKq7snGlzu1RZQZsWt2la3
978aPF3FXQEGkH/34uH+oh0fR2SxvimfHzRstR4/tKObLVE7NR3+gW+bk9oqQTyk
MgLGqsenOo5UGdMtk/CM/rSv3bJBJnnr8vnjzKD3zgHzxr4M0sYcEeWN6TDChbB2
ATGwyMvoKNy+hVKTNHp1stBdaONMCb5WQZU6QFerhbuDUhBwuoh2KevoKDnE0Lad
T5qXQcjoFlWR3FSs8seLCqFzJ0XtVlt8lLn0iuKNRycXwGkZXAOm6k7K/fA7dCNT
jdEE0bnclqt5fcd9hCHIrejW2y7kvIH5prPA4WPwbLPKa2nlp6cXY3tUvLPYOBn3
W9ycbhz8LZm2ZnZxhhtBmm3/0kVeWUwqhfehTrB5hpveHMDR9D95NlviDXuGT9fD
HM2YVQHqBoZ7coCz9dDANBkhypxz0JSaGihshNNV/0PHsuEfOROxC/SvqaWqptoG
wYtUO9lgbzu29vqDh44IQg==
`protect END_PROTECTED
