`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDV234WnSHpp7H2H/hEwyqK3eo1wnLRr69wKX0XNOo2l
Qro2dMKTcobyBej52vKnEvA8J/+QxsCqTPETbkPFAIIbcZA1pN8cVqpzQ314dNei
OdM90HWSxUHSoBhDdVjSafGz08aVLJ0sN/d3hgSLWsMyfMJQeE989My56+yPMuPG
ipMDwVAU/yZcR3WIDpkz71Mv4vJNCYPkzj2rT+mlGdbiXOIpQpJuiMGGjz2GGQUt
y+hcflQBo4hi3IsNwcJn8g==
`protect END_PROTECTED
