`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
w+26GqdkPKBWKp+YWQxFMKiM9ubfzzXElSKBRmW5PMVs1xf9yUUJzT+hDzK7J+y6
abiHUGlE4POWFoVTMVUfSSM2csWcH2PZZNe+LkwN//nL/XVZB4093ifbzGxS7uIi
RtTDnNMvZ1O1e70rxReB4ch6npOLlqjimpgOy+G+tsLAl5yzz4ujZmivRqx7HiqW
Wr8Lv3VR/JjemqbdYgkQkJQpnl0VHhkeHe97gWKy+rhnl3hRhdizbBAOw2yY3vvI
KvpN9kyDWbkBV/+52hZqdz0wYEz/5R2SyZFzGG/O2Rj+NFzUYKe9Le21KVMXckm6
+hKH+ejD+/4ZJdHoQ56JADUwVyTUsrgA04cA5Gy9coLBW0Z57nJ2D5zKBZa6mfkz
4OqRSWWKxjPDYVNfPnR6wFtujITbWe3buh1c694sIXMrTMtHgTeq63wnUDM6YyyP
A0A0WxgslZNUlj49Yh/0orRCGi/DMwHbnkCaybZm2cRefc0b1hpkuvaHugMZNXib
7UBwoz2X0T4D22k3iRfupqKQbNc+1RWgbnz9xbIQvxANM9uNIPFV97SrqwqMh5Ue
/XDgsxQMxsOg0MbLFZ9tEj7aLj9cL/wU2BfnT4cq4v1NDmvOwFc4zCQoYD9VNrj/
PPXV/X2YkpTBU7LEhvVJQIQjYzVAu9I+jy3qPq0wjrjEHnBNVGQrgMEuruSrjsBE
r+Xzu+XjtZ/E7ac2FzcP165bkzh5Eln+xEr/+JddwRTTgb4nOpMUxTVQA2Tka5hE
lHsYeuc29aamDAFzh+yIN8+4ZD9X3T5E7G4sJbj8N/WQEuyGecl4ZETjkiyq7G65
Jz46nXv9U3ta7ohBP1j1H11FHRd0pxPW/dKYH70DPdcocrdSwG3E7+Xj/xvoEqoR
PoGiVtjLOIAFm2+VUGDqIg==
`protect END_PROTECTED
