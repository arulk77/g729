`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+CK1bf7lxZH6Aj4RDavrAnrkJdpdj8c/Av99wStmMmz
QkRXxoZEgvnPJMBWuvYTJBxDN22dKYjk1hdf8Iqo8E42W2XibU/EzrLoa0mU214m
KQgCRB+RWimFTLoh+qDVRjyph7TXccXg1DNJvUNZu40=
`protect END_PROTECTED
