`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHfX0Uj3XA0ppAxASgWT+t/kcJrTbTgy/6CFVn6hjNSR
Wcec+N+yLWCIFT1B3OCYQKVrsAOAUk9MCLu5AXgqm+svr0BUMmIUUV6XoaffzY1Y
INU3k3tklyaGp/5JHYBqpmQ1AGaO+pXqpOdvtqKAQEw/4qR+Nx44YqfTvZKzXg1V
X5Xto3O1oJRTnbEwQh7wJv7CFEobMe7cHvMzDGxjqnRi0Au1ygxrEwq6sKuasMBv
FoYYXDq36z56eZbm06fVbU3UKV7wfHcPnQEx2/TLqMWdQ5bxKWzMApExqLJarleq
UadLt25VB0mPjxMN/6RCsT6eCgiRFTaPEwTwmD5iCsbROjXy7Zc9yDH/QaGcF6eg
C1tc0CCG4ubryxDEadUG1ANv73JezMt891NxV9BdmqpjNoAR8DIGWroO1WUYPE3U
KbXnYGJgv8K6215dMl5izcPNOaecFg9YbYWApu6bbq3C+0bOxitWdnGn1WETAwYL
HKo5ME9ZT2llq/74blF/JfYC1fR5ZxykHRTGKZQrpJvKlunu1PvsxPdLYYAzQ4fP
`protect END_PROTECTED
