`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu483fkLRWCNx1R/oKzSGvcS3r9ESXtGO6Gl89MvrqcTe2
7v2cFE3vCCIiilWz7bYVW0Nydowg/HW+aLh7ofaIwwtCDTO7WBmTPOPjg4mw9PeO
PvJcLw5iNdDBDk8gd1PqrUaFcepH6oDrio4PDqdfPKswzM4FAikoeL/icWAHT2wm
BK80jdHcYBN7ljTdNcwyQdkwA4B2BnccHnmzhJLvpUY=
`protect END_PROTECTED
