`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDn6gDx6ktmbmwtMJ3VTh+K9zBgl9DGpPO/IN9BMMI5d
XeT1EsXdKsdd0OYGdVgM0y9GL51tt8ZAF1a9j+czaFctjWDls3RGyR+Urdl44qq5
XjhMb4TAD4Dx7+23jDSW9RJmo7/rCdfpDoY1857qGtvzzdBU0BJINYQX6XA+lM39
yTeULNCtBgxSrLp51MoEf6j8XGxJg1YAWNeHyNTPDgjZ8Of+NpyGfI5fpLofsF5q
jp9lURh5OxjyYg7XfW4F0z0uJrs5Nuy6tkxBKU19KahQ3rhxxI1xTnKux/lDui9W
wOjPxVgrOgFBTy97UuIxr7Of/fiyq/P3eSN8wH2ZJT2DgCQIt3Vfeb2ao+oLtUWi
3+oW9X2zJ9NBsMlf7BzlVV6D0BSaN6+QLZcKHMq2Nw0llaHzPYFojVELMeSHNAVe
VikKeHoYVb8BLHM90UUQI6qqUERMiF3XE7GugHiFHXm/0DXWTl/fvmR7DtYQK/C+
Cfmis1TLf8oJuXWtrsoyaohaP4z1imrpMKLh91+bchi+YkytTazktMC+XmX+ZlZV
`protect END_PROTECTED
