`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mlFBzCyNIVABC0bhYTMiK8tZX25bRnGSm3i1b+/ZkFDyxpMvRYrnKarEATy8qICS
EyHX6TCpgC91HeAf77biiGyHSY506bgr0u2lScVwYdUSu5SN9VQJHzUK/Kqx1nV6
DhCRi91vPX/wAEKvRrMn0Ftc+i6ZkL2gvNrlKfNe3pWGbnjqUvyqrurTmfwzEnfw
fTOey4U7mtXeS+1OYOIJqg==
`protect END_PROTECTED
