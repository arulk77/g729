`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNxji4DeqN9r1uxNAPf3FmFY/rNrGz/0Zsl8tEwT5SXI+
uhj81Ibmcv2PbVRorSe5ycPiH+LccQA4en0+nf3tb5O96IJN9F6i7pEn4EI8qYjb
vjUtxncUEcH7KLtPSL7s3j1CaYidzwxIzk3+jY3XlTkK0W6wREpnwgad0Pezzvnh
6uTWVkttB+JPn4XEbNOnlb6RCgs+d682BaY+ny+PXVyOIW8q8RAzgFBa3c//eyJe
StSYprNYQzh2EVd/rWz0qF6PFroijQYEvdaagetWWGjQsOlpGRx+8MTPC9QJuRO6
R/PkfhIY3JAS3s9gO+C7tmoAvQRiRjb5186TsZdE+u25kLoaoJdca75chOGQ4WFq
KuiWj2rzCPXK/Z2V01kSJcUSQywsGR+j0tHBqmqCJPuyoq12VbjbWU/1wLbxrfhx
nIpSL8/s6l3X4FUOFBuBl0ZgqkQ3PdL64mWpuMp0Epu0leMJ8PthMF2TXNPPCWtB
Os2ewr8cOa5VaowiyCUsHGCRkXeS28zuMyhA9re1jjj50U8oij74S1hTYcUdtPYH
tjlpFjbx+0pXEFNFZcKJB0Kzv84kP4m1F59Phph6K9210XzKXNyVwKH8ILJbDd8k
GUY8uIhYZVyIoR6HMrDokuhUJwO0cz431TgLyRAN/XA=
`protect END_PROTECTED
