`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8SSI/Q3Gd9Em8I/l334VHh0dTcXw/IDigG2zrtNXGJgvp
CAAy9vxIZKPPoRACSapMwPo2yNfUWf49oPXoYk1cTpRHOGqFXmYWbOTev1UKl6sS
mtZa8Ol/QT4mpNxc2pyWhGT+aOWhkw4CJYyBU5xNeKu+YQjfgaymSiXlng3afhxY
+G+5C389nQhe3Ke+URq54uO+D/XPHpAqx7qmCegSV9/ruY83omihs7T6ELDYlhqN
AXVVftpKZb5nJOF1dHou7mk49rg02Nx7zq/F0cWO73xetSlZRzthSakE+Y3nUmhm
k/lGYDjEx/lUEVMFGqtbOQ==
`protect END_PROTECTED
