`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGIJ+3VGT8ADFrn+6hbNmrbKeJKQsPGcaEBbLa15R+xl
qvJCiMj63Ep/lBDBpOYeV3p/FkxcidZxL9aNlceBpnI0TdC3jYccILe2Y2WerGem
hMZSm446TUHw2T2rtppvLoQdnoeBjnlImL5ZMGsiN9/QOaATpOpgdfPzRb2KLIXU
gE9RVlbGbvHDBPJgcn3kwK6Jf5MlM5IU8crSOxDn4pVkHV9SdmnV4tHaFO/41f9/
1901JXC8Y1fSFc2yQjG+F0SqZc2jKK3COPm2QfBj370PZnSj3xa4lb7JiumOW63B
FrrK/+pXKvVrCENWGaULprLuVlf9WHvnqgp6US+Xw5JZmat0ApO70oU7yrmiTmAo
A95C8kpxWYDe4UEom2kSkrcQeiPxgZxC5lbjMHa2tAQHNE6QiIau0pGn9wcnQCLq
7a9ErOhhgoySM9J1zuUwGxDmSmFh2T/svGLFhLdpKNAHlPKX89JROG7tyWdxhHML
TcI4NQ2VvKsAESg2AsC9wOEHVtuZl4yEX3A5mCwx4VMaMdlHII5te05Ow6+I+Za4
`protect END_PROTECTED
