`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGGhKcUBsRM6arRrg/PytU8AAfpfk+1irBkxzUhmj4Zd
qy2x4OD1nFWdPZhD3Euj5n6c6BXBnTlwV0jK5v5I7n+5zZ3t/km20A/6lJ8JKnmj
HL9v7G7EQCKuRRLSBWac9+fxMz+ZBNEe3951ZfK0VZwveqI0EfIYHZ8X1w0A/m97
joOXn2LEGc7N5p1vodzv8VZDwosd/yL00o/VzjVQPvf6HaJA/WjqDDeEmrwlY6RT
1NEkGsfOryoo+WvED7Kj/g==
`protect END_PROTECTED
