`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL6vPZ6VruBdEHo5Qtt5B6K8r2pXsBNsrTAQB605sBPw
R3gIHLTVDpAbmLl6h2bU+RciGK9LXQQVkn5463u/4pkQ+oob0a+xVC2Z0MJc4sdI
Apa3E3EM+C0caDucTdjJJxqLiwDPWqkb5PmdpJAcmy9HczdKjx+S3fEPB4C9uRKG
pd9SRtz8gf3XwesOlXoEag==
`protect END_PROTECTED
