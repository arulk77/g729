`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
QHdhxYOkfENST5Uz8YVCRLJqgwLGNRPV2P8mPePdOoN1N45cgjjeoAWtni9qTHZ0
O6CDFJL2FusVweWlYZSn6HcoYmQbg7AlduLehpve8064am5CBbzD81UPTitWOKx4
A1lcL7yCFWHBJOEi99VMeKKwU4EGxnh9x8OOEKeqzsggCeqZPQ96+zF3j+bT0XRM
3WHy+FAaQFMpvROt05apzEuF0A0FbzIP2tnA+mK1XXi/TWUjF3+SucsSeZBugRJq
LUNX72Aq2X66HU01aZtsZSZGUVhvn3Z5plPWz8HvQO3YlhK1dDboR9jSJRY1p2+I
ojIpf3SOFO72S/APvG9AFy5UKJt7Zff9FuEoq1bhbyHsrvnC7rBGKe4MJ8/u1DRr
hNFqvL6Dj5kdE2TF0wzxCK+7V9RdmIF4e5oxCYmMu9iUd73NPXfdTNQFSHoDrXlN
sPs47ZF4UDBajcmgQ3X8zWlfX7E2r7Meu2e2HTsXPIf+NtI6TEpGk33JcHDld1ej
OCYQywyT4YR3jwHzZ5DN/Dp9BUVzjh7rZTDSdxV3NWVli28JF9po0qc1WzoSsvmO
`protect END_PROTECTED
