`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGQOC5DbfYaTOfeBoVNYnvMv5NzL6eueTzRtk/bImnjH
j3SIvXBrS7IqpMt74W6KupOKtjHCkpQCfuI0ojmZaJjrbyd+u3Ejjy6fMPQYtrag
ciXGXH8NB9drSGQNbevWH+N/+yWL+3auRfZN6SNLMdisEP53TcGWA/Se20UmYegk
+mqb3vw6fHSZTacfJ0eLcVPqGJBR0JoIRQeAVNd3lOa9SoSch4GWpOr+GLmgAsgb
k6JfUvh8whbOHnM8iv/J+JgE3f3lwaQjbzgD/ThSKxCAVnTo5YL+x7Wltszh7rEY
nKjRWAl4NU7dvs/DSMKRJESXCqB5JAP/kUmewPohWs9U3vxW2sSC6J5yjuhiNE7l
uk2VTWgBnd802ubN5sgMUb7EQrqtXaS5+rSIeA3BzFcbbFz3LH3cHXohjBwQxG5f
G+caYqra000S3i4WMhnS4TEmW6PrX9tTOo+CJ2kP6H22ke2roTzgbq4XsOecdSPf
gjCkcxB8SgMWYvsrNaYYq3piNjs1EtQ7sZYfHSlX1JLOWL3IakqFaTCiaLFRbRfj
mpiKbXd0dkcbtoqtrJPQmQ==
`protect END_PROTECTED
