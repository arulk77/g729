`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHD1gwCn7VrDAuAhsK4Yo6E5lk58ETCBmcvIIf3HXkOV
nqTL95QYwz+NuuOaFFQhOkZs/nTAGIcVijtj256Ti/hxiP+XGNyxUFcSQZmAo0Nu
fzg4A3cmjr23q9hLeJRiVp3ppg11XU1ezn06YOY/kwUsEZfHDS4EDxUFNr/xBAok
5uMFUp0eME3VuDq4ULaEeA==
`protect END_PROTECTED
