`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveEpspN9RZosam4rADUa5GSS8QCqe7GLY5CX9t6oB9vFM
Kj586MWwEAw2I5/98+AXS0WnYZqFvkIUBVLveR63d8mXC5aVAWS3BkftRUfUWs38
vQtevo7GLaauJqFSUMp2cfcXC56Hz0hmXd/x5XWF6mQ7iH/HokwFNHj1MBqTn4Ym
zOkMPfzG5fKwsgUs6B7goEegaenolQCHRg3FqGNZSUnYeP52+w+F3kXVjZvhtZJ2
wCZkSalbUY/GUYh1xBJG7Q==
`protect END_PROTECTED
