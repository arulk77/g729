`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
E8v+Ox1xWWNKzBkzeK70IQv8E3sGg/7W9tjHkKDwLLc2UE8+8dp9lOIJQHXw6xjf
JH3kJWa8mFzhMZf+FEqI/zGXhTYkpMU9pXT+aXzoc1oRx8LkwDrQGQP4K7BB4O4F
LorJtwToCiYGToFUVuDDxeeTsH/6beeTkUkBycmORlkdy7UFFZDYvcLcFEff49jO
JeQvnR5n+jkY2lEBnjvsWFjMwpPCjTMA2LFp+5j8db0=
`protect END_PROTECTED
