`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveILKs0rg1KkMTji4M04kgkiDmsKpCVK5teV/XArjGdMs
pyjsTTA2Lpvcdp+Lp0/Fz3jcjEl42cw6mOU1uS54tuoIHbP+QaROujMXXe2o2D8O
diOY9N9Px7OE7RRfjmFLYpMBq4z0upZCarG5fOy0174iGv6I3S5bG5uY8fYkhoFZ
UqJVtMHZ05i9ZSJy0d+XaZZpHxRCuGGrZTq+k3E+t3oxcjVsj8W8xcs0WX5MiqU7
lKLtnzHzGOSApI9AqE9RbFSipKNAE+ZpEJPpaGJUisRLIOTrzujH3NDnHvXL2Eig
d836CLlvHv4PIiAeMG9IWXMRysGxr3tTzteFq2YFrhdleeqKDSF1KKGBC4Ku/19W
4M0NsNtttiDAdKl7ffWEX+g4Zl9r4tvpI4NKqjLJTQ+EUSztPLEpf8GBW/Kv0Ye0
myozYOyfrXW/dpjR14TGHyKQ0eDhp9WrFyUxYp7Hurfydd/U/t+8AaRut1rtQc/m
zQwaA+SC23zGbXbl64Gpm/v/IJ5UNmu5bs+7ullqDGdNUipj2ECY5w17SOcid1YB
c9DrMCg6WFgx3yLEd2XQPQp6LPwkti1i4h2OqKVTInQoa6BGHWbYn125wGakUQ0v
Co++OMDlFwL+a/gleqqz8PCcbExwU2Wa2hPViwyb1UJo7F7S0QYOIu54oDK0JSzc
os/+1qkk2u/lxw8fSkIODqjz0nOV82xP/mxXHgZWHA5buY4v000j7djloLUcjN2t
1ZrGpc4HcK1NFOhdftpzNHVe+zu4DuwkLEFRpaNVj2/I3afeB5xiJfM1xJ20+R8Z
cztQm2ZucOhxObVz9fE4tIygAYGHRR+1ZvJvUJNCZtttUvLdKtZLlmd3dnsKiFCZ
v3nZJV6LOOVaac//G2bs0f1uOzgKFRwV747xmwKjUoOw/94/U9SHeL/tqLuljjfS
4QwGrEnfI0QUJZZRO3uR1cLaJGk8IJc1k/pRfVfLTdiplk3d3ah7JWbTo7tQT1PT
YfhgAdUE3wZZY43M+vCP/VE1hiO8mxRUHikrlYy9/Tw8aCByWEMQn6itC3DZICVa
NcGsGVu5YrZe2zPr0yfdKjVOA8KY3AwJJftFOAQmmYyKgdyB+gL8i4rDEfkYgz83
Ldckkqk/0+gG0G4JAajXLa+/j6kzlW3xLoBppcIwH/G9b6PJF0vn57VpuVFCXUyV
Hh3AGyXuY1keX8I4XursBJeEBRXsI/XsLvZGD6DPFnALucF3kwnXarDcWO9nkdF5
pJ6wBjWizN25oGTPwU+ppY4ZeICtSuh+50S4kHUhU4PVLEVGNzg5CcvVwlgPD5L+
wjrqD5G0GDkYZAoMC1PQ9ewuZnKfZ4Ul0ArPd5SF9jfJSH2CAxFbbZh89wFJoQu1
NMI/Tq6Uc9nCrDiWbsv89srSKlir1bQGx+7gl/u+tsmqsbT5208YwKRwvnvZ14G4
Tjj4ADbcUwlN+fUljwYsKBHNTSzvr8Gl3tbARGPJgJkG5dQxNBMRv3IMegbthQnH
idYKsf1NmM/cdpeIdDmo5kLmHOnjri0h94I/rTFHwgmsmkHwSe+iVaEZMEpcKCDg
vE7fCQSUNekDTjlcUyBCRIJsQKGMYcW2wc2wyh+vsWEtqr4qViqprNYoWqAls+VV
6M2dVn/CAo9BqLFdAeTBNstPt6NQsBKYc+T2uC5ZLT8emzDQo9TYjMwfhC2WiI2L
4iZ5YeC6whVPjsSjaOnCRN5Ou04jHwH0jc4Bw5iev0RtYPloZ5OyyyHvEGstJkQ7
jns+dgtadyJBE64bUM/mupYk5TwoA8zkVAEk4UhndBcXwE6D2tk5al2jUlviVPG5
cvhgQwG06pYxNQ7K7XrllRPCWFevV+blM1e/wrSAC+wRPv/lUIdvU74ndP/SBX2+
GDBFAkr5UydIC1IHD2MkqNUaXmTG757oM9QWi8vsbk8cbl9zielRQB38gt/zud2q
TqGdC6ukdQxqklvw4idFRtmsQuo+MGlJ4QzuM77wOOGtVm94clQXtwn7A6jooXFv
tBVJNGXTbo1BiLOALnJJXYDFuCLWIfTHgFhwl0Cx5ion0ThOGjbN/1aD8hSkfcdN
kHHEHfkP1SJap7IQDay3rDSzb8uGFU5MmdRKT+FruelvV4xmAlCitpRSZb48m966
SJY/XIx7RUQVlEomFP1G37/VNAdiJWLtwIyN4g14/bzbup39ASGQcMgcUfEpkfi2
cwbbQtzjkzigAPRenpM6CB67r4iittkhU7dnd6O4HTtf+AGGqiNp++83PzOCoLgG
N970hjh7s/3+Ru0hXvlvEAnJuha4i6ZUNu6a7SQgA/amNHpBWhz3YUeBiD7SA39U
qmgmTibwAOWXu9GSaGkjTZJhvTQdgvay2ZS/MU0i+HXAz//4ESCnQ4LTTFDWlwGa
usWx2IAwfCJM2dXBkQ4bMs4zgOG3h279IFvQ89DmgQef67P/DIDJjW3GGfxfhEfN
qzzfGNiaNL2d+UboS3fiH5kI4svm2HfGurxSQTN4cpwmgwG/0LGMYkD0Z3IW7SDp
OWQ7rDkrmB3GsU7cleHQfkZ4qU4uq6CcxYljs1DeK/jKpKoBut19eXmy+S3lTLle
kP8xFYUCu9QpRCc4xZRURgWweMXWJtdUVG+0bG+tp6MUMbU7lepK9IWh1nxWHSG0
uqIydARerP7claKCv5KPh0Uv7bfZ2ozpEQv0VUeDYw5bcAB+w0+SsAGSWuAw3oxl
q7jryeNYlEgTDuckgdVxVPSxD3QMlJJrQLK/HpAUHCGCnXDu6eA7bKmYydMKv9fZ
fNQL6A1DwVCOG2hrvT4dPFnzcseoG/iVrSZSD4SvznzXQ8FRUR1SDrnEbUSw/5gg
ipyOD+Hy6XlGwpw0xzA55QpF2uWCw/i3ikkFxMZYyxU=
`protect END_PROTECTED
