`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4+ab5/SnjxnGhtyx49w6wF8c437q9R+esNstS3zp5s9x
TECYM9c6V896I6+W2Rez8Fw7JIM2WPxswYhxLaE466v1iceahTv73tPCe1uonCBw
v1tvGUCtAMXZ7HPOXOiZr2dhmu78yZMHjL0IyJnyqYZM5EddHs2MsxIwvVPhhlXD
3gOflbHa0Ab1yJZyrBKYPj/BQsy1dFnuzTuhGVBBwYkGkZ+bfGl8AbtxhHsYfg5l
ULsT8IOUWjZ7NKCkllF4Qyt2PsgTLyDjKIG2pcGeQQZZO2Sk1iGAghrEKAYoEuV4
BS9jMoTqun+GnlXg1jFuOw==
`protect END_PROTECTED
