`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
AAlj3B0RZGik6j5MAxcIn210J1My2k9zHvhgdhdZZhz/XsG+HcvtddGDWJB4jR6e
//3PzIhLrT/J/1XdUCG+xBlggjdqhthOaTu3lJcKMj+r4rbA+369ZIpKPbSE6Q8b
FXl/sQgWVrDGd57/5aEnFQAiFqJ39NWAtKGb85vmYFn9GEuVHEkRhOVNaYDy6oq5
vcf3BQhvjXCf8PPbHAIToha0rYjhA/FWM5Y/oSJqWfEOY/tlrpoGsoAs/aeniFkI
fT6T/x+cHslWq1bsvouChPf8fMjNIDEdsY0TWianZas=
`protect END_PROTECTED
