`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ+7zcmILLoYclmUJ/k0YgnkxXbuywQfNsYct6tnxfcE
3ifgNhY7EvyXjJC/ceCi02rKVa695mVez9/gm0A3OpZLi93bjrHBh2IWIyHkcEyi
EJuM5qgu29uqjbBaRZqZ/U8BOZ2fQBZszlEBXXgvMfRpDmSgOkDWDiWAYqU5ELRN
`protect END_PROTECTED
