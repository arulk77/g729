`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/9aM1SJDGFULUSOwPoZyOsJLiDGzM0SMRvD80z4jJsJ
8Sese9Ou/0QR3Xt4YlHX+xqyA/8Z4Wi5R+/lDkRBWWkHcbmvyUjAW+XP6b7rL0g0
gM74Anjpq7ZrxPh2LpqsIiJ4qNg7qQItpEzV7IEcIrIzfw06tY4u75r6h5E1zWyg
1szu0B/0/irCeYoUN8upBUhL5Fw4nQCbQsEXjgz+MgidO9aGp6STXMeYhTJrludD
WJuRoaiJdrcmMxsvLy9mzgm6O2q0E1ugS/ubHANV+8rGp68CrsM3oGvQLxAju27k
h2PuJt1/NPsTUtgms+uLeQ==
`protect END_PROTECTED
