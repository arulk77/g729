`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
/b0aZeMgnTR8rTwDUtgBgWKv27tvv43dhnM5FH4aP5JNKDvu4nu4Zz5y0iiQ1NAM
sKUjdmzNJFctwX74Vcr4gmPSCscnudHM174g17UptUTQnAdxuA77bnq17Ocuc91Q
da3EIDJPMOMfQDrJ4NSCK6dXlDRm84rDhR+90JgAHJA=
`protect END_PROTECTED
