`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKZ1zQYrAl50LQ7giw8s/Jv0doJvN5PhItokduiyqZW5
cbuOs/sfOGjlHkl2WbVHuAu1P4VYiIpXDdkWOp1jQrJxautOr/mhK1zLatlBMlXq
tL84z41G17kIZbjH7GoXRcND/KeL6l/BSmVcaxjLn7XsunJgIGrZWE6o4VWl/cx9
V9ppVDqUYo8u1GfhhwX8Zq7z9nVP716/lGu6teQMDhUbRRfA+J+8dGVze6rWaQpI
7JQ/vbHyJ3lMD0rtkz/6ogp6XdP9akq5de9o9Vz9dmNYcJpDeMMLCmCr6MpT9amY
SC55d67Mtk5f7XQYbhAcYxvK1EhuYL3SRRLu12DG7hkLz7fde+qWcrMg7+VsGIMb
MTGNeh+Ai/5kTrceccgH3OlxCEXl/UfTsWpsFbbZBLSanyPtaNS6pVaPEmorqL86
QGGg2uMb7xXDC84Gy01aov5Cf3+tQS0a8hTk4/wOvb5HvRyrpAWF6mB1/pCNvGbp
eJSHVKsKzXPbzAZHXdrokBH27aZYP3NtdHvUxNVStYEstI6bC6MMqxgQC3MLNa0L
npyeqfTpJlJhrVur8h37BkGN+vihp90jVXddgLzZz5Gx4TPe/+wCuo0W5SAdbN6E
6daYcrvzjWHJteIm8Th3OnkLspfyIFIvN0vh3UO1yyEePRGz/g+yd7ErBYoEioFu
s1DPtBVpYpWr6Qm6Xca88tR8r89EClr5lY6hWY1jhUUypVDdRh/ywLACof+G7mYb
lMpYpETU1reE7LwtQDrKsmDiF9niRA5+BrrSh7WutqlWk3HPd0pW7j8um+bu2jdB
iF6xepfkSR8ESsKCGrduPk73Pjs05l+S37RcfCnRrMdzRDCcPwXqMFZuyfNduhNU
3ovti4ftMLuTmm5r3PMMpq6fBlYbmh5YOtVgtdpLpSE3L7NESmmoz7aTTrOkxOo4
1zHrQ/efsQnuHnmsw8Q/CEhej0/HA5TEZSLJLPrqqPEtqOPyW8ZBOSPmYnW7C0nO
yQvAcvTd4rB+pFKPOglZTAftTJ4Ge47pTDGevsMSHMw4xCcSVrJFrJjpyiBlLk7c
6ek+oIo7aYTqKZlKUAkysF3VA9PYkIsrA887GL4BKaT77YoSR9S+fw4zX2NTgsO/
h0RjcI/qA7Oma9SnaEVk9Z3v+EK24rSHrifBONH0Iz8mBcv9pozUpq1PyWPBAOTi
dG5qAt4PMhCaUHrRHYhl9CDkHPs/CBy5OEyXleen1n8aiZykAPiCUK13n4M7xCWL
8Dn6kpDoduzDLuaVno6yQMwn4X6XD1mQRdb4C5Zjwcf+ekJLZ6QUacEq1B0DfKgn
obeYHIeKgBdaKcs1oMiYRJZU+CyqAbKs7cXrsjQDM30vAL1zFFf+imfgk2YEGtOm
lJLde5vc4hEdSKGq4+YmXBtxJb+OhOo7oMYk/XmQSOhV4sSnLYbaEv33t989GzEV
KIFnfKGl1gnMUJ9SQbHAggT/zvQOWKyhfHmZ/v0HHcqW05WeICgijo1RwbEDj3M9
xDLW/pXwnIo24kXaExyD32yDiGIBytFOpEqU4jLIgxQPzFVYzRVaE7IOJXZ1/BWm
3W5XLz3xIQaFROXo/ijsHVF5V5nb+haNj0kpZn9ldWYSbus81a/WmHupR/VQpbem
gT6CSAKnMWJ1GTd11Z78JX3oCDFD3GoM9c3foDP1u9zO/PtPafEHQtSXLwrHg3Ki
1TRa4pZhQMfcslRzhDfIJP1y4xtTyPCxDQsMU7b2JFlX4FCmswIvlfV30SJTtD8K
7KssAgG66x5VD9trPNCBWJoYVgfjqaTcsXmTrx/xJLvQ8XG68x1FSSv3vNpyXoo5
1KD4VNTodwt+KY2Y7lcr2eYb0x4AgP72M4Rltp2bTfz23a9AG8X49UGBIinPVlXL
U9VEgpa7gqgWYAarBhB3s29PkemOjrnpfZjpg7ookk/BxJfAICFmVywkkx3bSGuP
uo3+oMIDUeTZR+xYKS/VSWLapS7QVsL+aEqjbgv8Q10I2lDoe5m+XVEupOZl1Xsk
kccx9Z+vUKx+VA4qFCBLu9zrhltRzhdS9tRAMFMfUIALqNp6xah1uytate3nnYtN
GSRLcYqHgo8ZIpaANQrMtatd6QSSkyqKAng5SuQIE6fFqu901zrQRrcyXKdKrdji
JPpi7CtPMHMuFRFOB23R2uHAefK+vaWE5KuT9qA+OqRJ/MzA+MTTqbmpmqiLRz/5
Q2gDY/2PjglfRZ9G0P/HYKqU/qwkXVpSSebL30n7Fsa4Lnt3/aIfhwFTf5SD72gT
hkFFgOpSDJcZPid1IoQDeueuTmVPyCLwIcJGGFo6dL8Xaj7e9IJKhVAyQwmuFcj1
98iT2JH3hjTQSs5Vo0k30txLEFFtA+xZaXhjuqxLKMK3erOtMoKC0tqIesRwMQ5M
W5DbqqBTPZmYHUmTRsfFxXiD3WvZ2e3saJ9lI5Rb7NLS5dAMiY0Y5LnoDY0szTa+
zFtLFBLLkkCRePikPu67SyUbZ6cmAkrLpqN+Hdu8zBUSXAwEO+sbTOsbYbVoc785
EjYvvBRYCdzPAx//blgMmD7rNDS9oX4Qjql44mYwxoMiqHXCkcof7tRZyoJanZ6s
FNDhXoR2j75+TmDV5whCY4yG9RO4+Q1LXRMG9pqNA0XJOTJAd4vUUPgxSZNPpyjT
jEyxttMVjDAkplcG0DACVFuxObYPwI8DWTzIGQcnDt5L7RvVR7TKv48kB8zZwdep
K3CWgI+N8FwuoPi4Ma89BBCq4g1ogt/TZw6Y3OI8145AynZ5ZLKmZqSpLWEOJ8LI
2Bh/L1kBXYr+G2f9kntqRhbgf+LKH64EP/Gf3lI0TPXQs0mAK4PzaHZ+C8QCIKDU
2hWYS2+TEEdUGz+BbYvG6izs+mSsbAvue7mFuR+eSqyxOmBLcEeDuK1VLx0E1wVP
xH8k9wtu2PAnMKEKtpouXKPbiwkHqfqK0UxYMdUCYKV13dWNppXUm+wpPcSOzwJI
XkmFqw+FzPTXkdW3eu8vhOIETpGhCsETVV6gT4R+OslUcNBmYqm8QVm6T+C5K99t
C1dgV7s2nWlopYz+E7SNoD2/ccaZCVuGzbkNu/CkE7RerNNak2pAYKTi3svEiyLT
56g73C2PH0Ows7WiPnQeIwqPGNE31oayn4EILaSJw+/4YJ0CxYyUFFNxxyHMQ6WH
VJPFNAnfEY47ABJneG4IBN/d3EhN44Mggzf2NH8NUCauUXXqx2+N/Wx9EIOIN7wt
zYEIM2Z7KjehodcyAgn3yEpMYJf1w9LejWtyzMXYf8Cc4UIkx0nNRr3Fxj1BpiCD
6j0a0sv1hALELqjZjOjbX8cs3jDWMwYCnPrF6my7EbV/S8BMYZRvH41tateNtOS3
+sGWLmIbojlVsbsUmln/4Rf/kvbC1tjC/NGc4AsojPSTyt+hIzuojfhNxQxSnCOi
EPWmIhNO/15SKeSfv3qyryoaMyMyzb8Wja55Zj0sFeHuM1NgFMjtSv/WSDm9ESSt
p7cx1iboobljXDpgDAMyjf/wxv7DbniV0tP4iKdC03hPOyGz3VwV7/icl3iybuk+
27Q2b74ZI5kagXMZYcaShMsIN9AAK1jaWSl8YOw+fMYk56FJ+G1biGS1UPVA/q3Y
Ykov/PG4OarcikZ1z1XMOJdfzar5svvVkMPkrgWLPZHN5YQc/r0+0QTq3ifcVL52
dkeMlHjvl95on9wbAirgIFUe9Ac0Cjv+RHYaEFmsImwIeS02OXKNSWACn8MxCXwt
ikCR4DeLozkW/uj18mMD9dMiTMvc8FznmlZTQG5X2ymVJm6gTRGycs6OEtoqQSxK
Wmw+cVoz+TRo7w48rmw3j5nG/fO9J+kMTOmXG+2IdPa3Mx69MfILYACH7XNWIxRT
cOcnEYeZUExZdFX/eQc9AN3vXvqLEa2+lFtmdetUwProjDEqjdvTcPiJNFBB+qb2
xExYDwv5moAnHUOnjiQlIW2liR7UQXgMiziaLz44y5/wlUAYTpTjtGlB7yGdXynJ
tTvAhgavvuUGPgTNKGE63sK2BBKN+f77uBz/meemEyMhPaJ/K3Byy26pXxWBFtGr
JhFy6qxaH5WDlfFQzNGAUCR7tx4nCRU7gTaoac9v/cG8u0aHQp+WmOX7kLWZlq/I
u3ghVgbGzveyWzSZoFnqupqU2G8HqxD7YwQkcS9qptMhoH9aErCUEU68y8d/GXA8
e0aS2fgrH8uMt9lJfByZK/eGMtU+BtCxp2hyYNLllSvsJnl2Ad7fkMgk8Mm6k3i8
oLbW84oCzr+hLnjpoNmIDLPXK8+9tl5cMiaSfumbiTo7DFKmvvfxjGWYdDSP+ZBo
c8MOHoVh91ho/pKpIKGJhhvKHYQNx5jlQJxffFNYRt4xzYgCFOXRmgHcU2JrisiZ
sZdlB7kdYapWH1bHdrbtK6p5kfBKWPcdZf0+gUqelA3u/EWdmqJcTQzMyWhcVpb4
c6tHkP5gmCH7FTu+tM2bPlHPryGih3hMpl1ePYrfJmX+PGhcMoZUAvjsVyS2NOaB
wQ9kXrdB/WJ+xIXCq6lNnU14cnEoccFZHHJN3OuMa5LXoG6ZvLXHivAF5VFs7DW7
IQlv4q+Kp2oZl2ITKLgi+VGokK2joBw/ZdBhjRJn27rgzGotzM2f4T+y1XR50ceY
15/gy7vIex7MV6Mao1Fzzl2YUdeDup5G7g4GrJ+E3CDcBom9MnUutTLOXGCINijI
+XsOgYArDj9yWSYrF5rkHtwwYI6INfdb4cfLqQ8moidGnW5pWhI/BzkV4zdRu7si
ONNlOjIdQKWhhd6KxtAq/5ro8Sko6mk4MZORnmQ8D2127uyNiqlEs/Q4sWqLqzrh
SSL40WAFU1NGZZdVYleqGsOa0i8ecMTIAi2AhNh1TF0GPtOf9Piqdk5+AzrZFvym
U95qMDo3XmOozCblY4XkXf4Ymmnd9TgMjGzsVceB7mnyY4ZPEAJeRvwsrwGWeDhC
F+ltevvX9iv29jg0Zih3Xy9y1hHUrmkb/n5X2Rbk+VkV58MM8XQ696uwH5tdHdv3
GJOliKhhuPcO0oQoNTCqnlSnPDWGSAQIj5zNloqzAz9zDCjt6drQ324gD94vKVIb
yDJVJ0z1LStbaB1lvHxrEbXrDoSVyGSZTugiYE15LssZ8qbywmZkgrddLbEBopJq
IBw6HJkDmxsssbOzXDQnc6oJY76nLijsFyBRFvjIzLSkoVRKwzMztlll0cepJLxW
8D56dFeUwEktL7Izh9zWTYrpc//Lemj9o/qkRjcRLDNWwG95rx+OJcdG4wL5uI5/
tVQo8A2j236etQrOQj0ipWWiqOaBa4QK2Ghjng253Pe9tr6VSG7MC5lhH0SBI1Yj
5B0Wud1cfVrv9maZpFoHtDWphb0CH+g7NgObxUmW4wvmbWBSItDQVczPmCxyGzvl
Ih0Xm6CEqodSCpCryHxXivSwgUEN5mIZWuygWp61NGZajhqDsDBFRMvDYmENwXBl
bjxCCCrUWJ5v0nMSQqxGuTTQtd9pbeTV6++N75casVNDuEEYlEkUQjZXXyE2kx1Y
KAQYWcyEEiFug5QZzVRozMmYkWbK4+D2ikA8ZxBQsXaSwp725Xi1xJEyTXgygMpL
OE9qgsy+rMMNS0vD7NY3DTp5N8kuVqAS9yHdAJ2JCZv7dOvgXV7s2IXh1p31qBT0
VGOr+nIDjwblhWQokROTGgGNQWWZ3iY9d6YV7jrLpexemXl2QfN7Z8XSIgxn78XI
hj25wtKNI0S/ovoiR9B3y1pBoWzNPjJX2sHo1f+csW8dvCx0/pS5Zr67AjbAppn+
tVeNAlEtzOPxE61mSb7lP9ZdjIogvA7zKIXVzWiNCMmmAQrE3Ga/+c8R5Z5PC5aP
dBKEmZ459Glv0QC7DOfB6JeAs/5/oCZjzRMlLCxVXMwy2Hy0sDX+7pb8t6qffDQb
y64kAZwgmD74/UxNlYzWJQ3uM4kkmHejreNMc4M6omVr0XxHJiII/Jl2qRQlC0Ee
rNVuTuDdifP2BZZlwr67JFT9My5joBytl/i9eEUMMh4MZE+ZD7XcZ1kPOBbeVTqG
Ge4VEbSj94H8wEL8RRJEgikl7OwCpXQ5zkDanKBMwKFVskbRaZsKzFe0gQQTb3rx
4x899Srhd8CyvqRdqOHg1gKALOBmR+iGnGgp4TDEXwTbpvUUksA4fDWekTQGWscp
gQd78OMcGRd2ehHZjbMfTh1jmvvxqsdjYAJc9JhCZrTd9fQYnHXbdhMwACRZ4ruH
OaBqRj3kuaWYlgi1Hwh8709Okxn0hn5qZtFtvYoawp2MOO5c09ui33h+XENkV29o
m0gs1+hS2RzJbMFyvq2z8dy0ZUgCjE0rLi84rajDpxs7Jwj/lZNbDFgI3iSAYPo1
Tih6DnHcJrQi3xSZVRuCerDE7uw00r7fK0z5K4YTp0faBWY+kdBhhpe2qAqYNlcA
3x87UifhQmARvrm44BCWm+voUu4UAu7Dn9FFg7RYS2tvba0lf2b6dU9N2mTAZDs4
ZFU+RCuMuznI96b5McfK2qGdqem6fMox7rfA9EH/R/Jmg0sD/XH+W0N3aO3qJsK7
iKhzhzakhxABwAHzrb+X5oIRM3z6aLXZ9G3G5AJKXY2WieDSq1lecZRCteN2mknQ
zh4UdNwiKIwV49zE4lZbO/m1q7i7Y4LILxAckcoY1lS/8CPWWhEQ7TNnWS4hVHio
YTH9bDJat7GIEh24WzFhRRucIYATTpR4PQ0dwStdgncBUKRTrhwaTREZPzAZbuge
rvvPIe+wfg14G157TMcE9Od4tWQTlK2Ex/tbd+sIsBwxoqIfjSXP/iw1OgwEvTi4
QROaV1zaKBDN/NS1wwl/bdZTu7IVgfW4hiw5gVN1IHU49xoJLvCkza1XAghM8mzj
lgXExOS2IKJkUjE1tiHOu6DTPutYuViiBZpB3rrbE34yoPvtBztKzKHBs6ygPBM+
R8pjOj0jL81Kyk8+yDQg4WLnM1OpRWZC3KdAj5yLUMW/nZlkVsrdK99XCbu2DEmi
KDBU8VY09kn1gl8i/tgYnUgGl9eqpv24IzH3l5F3crXhkB/Q3/01gcygVyCV2RPX
XSqUQdcnIAZR6J9dLTcOvscjqEH4HMn/rFervZa2BF/cCH4HH1ufKMcdHs9ba4K4
i2H085RozhhxKRqYcPb+y/9JRTef6TA/2pbCeYeIFsOJby12ieLaA3HzTI373uS3
dMCiqRqz7FSS6ey+xHLwxMYCnuhQ5uHSrUeBcufAjYMhNjkNZy0tAlffEUIUl+1e
PsRVJMsGSl85XXSZIBUO2gpQ3z2so3Zzi3HRrI6HpKaquMj3iO6kJU+hPg7Id8Hp
oFYEion4/8zx68/506Muv/cQF7P0ySOm91TpbmykbC6baFnHcWuKCHX3L8neRk0a
WlJStDk3Bjd1LM4sB0La3MBHM+ivLF9t2fMg4gTHLy04rv4g42oW3iFgmL9YL5n8
8kx9rhYGOPVgFj6pNtcAHIM5y42WCWC2X+sB+e7e8ky9Z+hk1uSrkvC53pfNShm1
ZkKeQxLk4oVAlAdmsiprGIwOYqzZzVyWoWOW3VqyWzVFsABCIslw7BT/vgIPkJuX
MVJCKtaOkXmK1uf8MyINNO5NoUGG+gh0Dvqnbu4jyLLmi8yPf9pKPPeCq7eRyD+h
Bx7mtOa+LjZ2yPDTw3B0agn7EvXpW4yQzHjteX12OP1P/1KaiudYdr7cd9LjmjfS
LJv4CvSRXin8ervgEMvSXvBoZ4+Rnz6vH7FMqqXiVwn129XJWFBtyA9nhp4nsDzi
z8I6E3aHhz4v8YTsGcxjnU8HsDldrJdluKg2eivEB5hgGXlGVih9xHCC1Ri7ZsgZ
A9+QYieh2hfFCCSHhDaLGM/qAcl7y6SfYVRcrBED3Kmz7ILB77WkE+K03RE2TZnW
6iHyDkA8cCQAduSaUJ3D1AJyQWTxsRePw+Idzd/W1/I6GNJFjvBWp25sbGQMLzpP
iaH3Ib6/87F99AlmkkH/+sKvu8tzakN6v6W3QdPu42Id4it82Hm/88iI+9IAcg0k
+BYhOq7HBuBi+RHLz0vz/mXbo1x0PSVTqKOm348eymqqnCVxzMycEfukVLbMdTTK
mOTZaalr6wynMhV+5aMlXDiSC8vvJ+klre0x9wQ7bPwbPSj38njLd6Pk2N6KT+2D
LXY/r87Cs+ZHaQa4ypd3yGq9rCUFX5pcuCY0+922C03nvPFI2MZPqzUdS8JsP8W8
UC5DSh0RMc1MNzUNkYDeE7XAsQVg+axso47kYlMc97PnmNjSnT2ox8FrewIvoxDa
rQ/IZ2QvN22Jifsw+xc6ovvUMHcNp4oSP3A5BTlFq4CGZuyuUYv5+I6OX4BDHhrk
MgfGiZHtZZf3ZfXlHjaECQK1/823hXypOU6jeOF0CgO62+ub/Fc6lilWY8JEm3cx
EnVM1pj22TarkYrW/iZdFy3BY8aSejT4JvNPjw7O531l1rmB7qncswASHETA6wpK
ofUGhKU7h8TEVAoxxFLgdWq5DWDNO6fwd6QhrfaOgut2yVRnFzM2j+EZdRd7d+tk
patfelfUHm19UFj3bjR/9bTING+fGVXqzfZwX+dKWmwYvQg9Qi+2KRxrF97goApx
F6I/Km1oS9EPrAEvnQMDfnze8xuDs0T4+mxk02wCjQaluCwiQaMb7DxmjspPTlYk
D0l/LZxhUl14aUqkEIPF41o52jgzfzkmTUt1m2OanqverLhUpznn/q5xU8YIhOAJ
kybql6bMXzYsuVohJDxqoyoSOkMDV4vgSQdxfG6+f4WjwSmGp9pVVpvVSTWrlAsp
yilFuEZB1FcKuvWIYDlu+A8hqqQzAdAiQLsrpIrPPD3VvwNyL7QRICtsufJTE0PY
u0JECOelouvwodRyphWaU3DwH3k72nzt8Lci8FMX8YDlrpM5+OqL1A8Lh1Hym1Mi
3qQ13HOCoACtp+pFUuT8BpdrTfv1M9hmGwrq+kdyIu22S4hAzSy/Gr6W0IsNv0YE
V7IZrStQ2CKfbKmRLDlu2CB4KUx2nwmV4XB9V83DCnw0gmSQNM4hcQrpF6ckvbcq
XIxz8F9zFX1pgfEZE56T1ii6+kuUDfrGgsY260HREUdDiOnTAG3qYMQnX4T9N2WX
rnXtutSvTQzqSAF0ZN2lacAbiOBptHzKH9qi+88Tsu7cvi2r48OZ6Ay+OJtUJisc
QDDuDmdikDUBFRqFGBbqrKdFrHXDgZJLfO9dmd16hBo+Y+tQyywGbrNz5dvDLL6Q
IT/02w3XJwhUwtqoO8I2bl8BGmGvgDNrtpksFea3VieKlh4M2vlAYdc4IRcQk4nr
B4+7Kx9z4qEsQF37VlB722bB8LULNbhJG78V/TRJECLopnrGtgFy55+i4Bqm3xX8
qQXIvFZRC9kxaM6sPXHdc7Dh99Sew1vD8T+1EU5K7pAkiWbD+rXqhKAAurJEbkZm
EmvCB57Ne69b5lr9aI3mvFX+WW1uGX4jVU5xCPIM4VdGxFnv7zksABIET3bgnbQ8
3V7zD3DA+kfA0Qz7KYLrpzrfazu9KlfhQsPkyYtnKpfU5rdFJggNPFin0UARSLOm
0k3Ksubyus0kuvp68JO+7abnRmgaxZyv885nQ2bR5cbqB1LoSowpr9FwAGrWj8XQ
CKrmpTDAU52fGvDM/KGfcMhpOUbCJpeowRPhN6vusEh8iuMB3i/1VLT36A8e/vEZ
XehTm/zdfvsEo5Jv2kKPfEszp8jk9FbxNCmFNd8bIZJcAJ53GTA9THaMGDgYUtwJ
BurOet4SMTK0QPDo3AnviT6ybEoxXM+aemOI6fDW+wOgRPIC0CxMZ7R5kIm/iWUH
lhmwpJFFWGkwjCwYUVzpsnAcgcGKHNH6VCKLNFnQ1LXVTp7jICJ9OCbJdcEzaY2e
q2jYQEjg4jNoEO33MOIc89TAErUL7fLC/fZoxSlXqQLvgQP59eBg5PuThsTyOgpp
v7IynT5h1npNQJRNtqZrLDiUIEVQSS4CRlX+ZZuXP+34/Ho2gHWrMYOaVRtoGc6p
rzUhFZK5HK6hi9wuBuL4P5yI8E4Jrg5PlH4Cf46lIqmQMw+PWktKd5dS8DEAH6Wb
p7dCitFtrb9DUk7ZkOPcQz2jxvmCar88WbpSeTTwgtyKBz8iCA/beQvmNm8y+oiI
KTnBYWvsrSTSEarZjVBZM/c2g4gXfEVnxOrH8w7Di9Q1a9KMrjaW/1QQ7o9hpI0O
L0yldss8P0TaBXwU3wtf8DporZDY10CpYcVeaaxcfVSaeyQA2r/4fnytR8HsFMdn
gEx6Ka3DO7TvDYCVn58FcleyUgj5G+iJ+dQkBzNpDLRftYSYNNS9r+U3JO6bk1bP
3RWD1NufMcbs3RYXdpUHJ+NBC0DUqdCQ7PQk6u02MPHFPVKEamqYhLVCZUqlihVR
m2UmmtbpaQDq8bthtqZj2K4RXtJhIpj9SwJNSH5STYhayQkn7fH2qtz+Rm2Reiql
TX3Fx0117AISvUvXwVMkPhBiJT0n70WZ5ZIs+qCOaE5GlXdu4qcJjzB7qCH+6EVz
gej4ITCseBP/54D4xb2DnAV6dxd4X+3yN5pmpi+AS9JkY+e4n+XUb26GEK0Lv3oS
birwzScODVidyEgFz9ZYdxSv5wLk4QvblqPJcIg/iZ8aexINxT0BD/iWltQ5FSCC
SaxWX7X+lUYkEOGvZlnLO86hn2u+0XXgjFkkp0HKGRu9mvXoPeWE48IDJyVV1/vB
U/nPMI1hTOzXk24tDzP1Pu1F3LN0dIbIsKcRf5bCdkCuGajSHCP7PWaRZJKxZTGh
mrzuRNADtpuT1gzNQpRNs7olNvaxDu64h5U6vIyib89EIANUw3eDacJEt1hEZ48x
vg+kNLwCiVb/Mwh41Ee1sbPAHVEhuUTPH2RQ+7M5XHFsCif6hO++75Xag3cNAhKO
xZ47gXasqgd/aQW7wsnZPu/EOsAeTAjO6dKSwhJj3l+jYy2P2LJDqOIEJET+vj7r
zxnacwYKmzwi/+PYgRRlixyUPcWjOxlIMikRvjQJvxP5ydQgzteohxzTL38UyN56
yGqxFrJaw+KJpjpPGeQlXH3x8DiVDVwVTEzGAE27bDdo0UPscRdLZWvaKlamOfoH
HIONMQVc642XkAE9h2wU/nnNDk1lqYPyngamLRewJ7hArkW5vwpVtcyO5c/8gCS6
0yY/06JKM3cvdGjW9jOkS+ZiksZ8/h9JAQs2uBWY/tXOs/4nI4MwpQ76x9VLihvP
aHCO2eot9iST2hn0aVj46ZOLdttUBF5xYgC7T1SlRtt0TXe0OvNgOsGmlotolsH5
/LX3NqoTuR35CN356/6nxJvMwcvY7xYXWo4ZbqVQnotMlRdjHg322pppo38U3178
Fqv/GgOY+91ff+lDpawGE4d8MqEAbpMbmy6mrlorzrV6bq8lfnA6rDc25kQ2k6ml
v2mCMgmQSoris3rtDd9fhTRmMOpV0fUvKX+jMOVYsnWVqa++mhBqXI6jQPnj4scA
CPvcl56HkfPZpME8EdQfgS1K1MdZxcFW67cUmHCJzOO1Ady7zTP+GSFHRrIPISvG
PpqMM077hAn/JILWdv9111uO4bSQVTWs+KFNpLNAV1ISbFzvrD2wyD068/xRYfiq
1dujSzyfhs9jQFIeFnP5f1PQYYbBDY3KybHJghH2oRRbX1nXyTJRdscvsZJz7DkO
7IzGvda848MQKifmlcPHrFCgzE6dyCrbC8nANK4Xvw+a4FnZCgw7mK2u8SnkGlhl
VMaZOIdiwTGVActfDQBL+OiV5yawwGiJIPxebQQVvFKTcxZqGFHZY/yYmNlDo3v6
mIqjl4WlWsXUCOzkJGJphxcxZKhlN/3/8E7WkrK9fNrM2vnXhgpcLIK3xigsv8YP
1b3RFKatv7UwTrMFuwamhZUToS6OTxW1ZlkidOLLbt0T1TI+nEn1g2/yfqcmAAO4
+7gg7Vw4N6Ps9VTq2mseww9JV9Pz29PF9BfYTB9C6KCEEH2JLg0fLADyPErMfdt3
1SB6V08Rgd+wmXxosDaPawcIreiAls/S+zvAUMsUrjR3fCz0v+yfSf1MJtYR00C8
+/dFSgzzHBC4ooNWxKwEngEf26oRpK4acpMk/GMaxeJL6OgbyjOJ32DO2bpu5H9R
mnGPP5Qr7LgpJeSVpPh4eUWNx7qPy5yMWmO3tQgxYxA0xgwU1hAOCwxgYL8OulK7
Azo0NPQpAP8+HsbV+UKGJHDcA7cArHp5jOsdKF7p2aKSV3CgQvLO2/3QIR3+MJYU
osXdhu/hmi/rMha8xYB7mkDIoKRphmvuEnR0T+EkSWEEdtPN84lRjvi1IX9S63tA
D+0cekpqiu39OBGNbAYCMwSVetXGKKHtycpRauYLsC68sHGFKkg7h2i1y/g4pdmv
oXFCLh0Sh6imfJIpASCAMZqmcd4CzHPu7go8j2RckSgCc/YA1WYnuLd7110reFoA
L/CJt+ab+L/nf1piaL8CC0Lhq9fvXnb9NBE0G3HhS3C7K7RU1jcHoDRDUoYwvOzm
phCZAZCczxk14PminNNhb/89xfTKB1yZY5DNc9OPo2X/PY65ZNmETaHingLrtCY5
WBS2J5SuMDKTA26yi9JC79UrgAjvRg6d++cg0jqdqtRCt8TQpEEveHCaXXHw9Gh9
p/mT2ygITntttPAwT5wqOOGLpTwiS82P3cXEiifWjKLNfJGZ4tv/T0pIKjlgmDHB
8K4aSv/lC8SuMkG0As7awwDoZjF42oy/13lcK+/49p9PhSZKUBLB78s7eT9qK2Oj
Uxp/7PKZIAy/SVh5qDO4+sn5D6APlzYYUcwQlwXM6/CjYO/dE6dZTmbG6shphnZR
BD4G/nMBMHU/LNLI9pBERyLDeSFvUqSWSgftIJqBX+LAyDZbrPUIWZ5akAK9wccC
mQpvz19yx2f25K/IChkNsS/jXAwE9VKinhGffSdQLQHTGvR88l0qEKOkNMWFBZOz
kyR7J5w9z3XkkzNnTz9Z5IUM4yA4bEFUAkC9TQdjMuY/qu7bnOwnNxCK6OCP3i7v
1RJ6g10S1nmZpi56pKVgfapFV479EPyQg2UOwA7hth+mdVa8FteoZeTwagXzkuFD
emysxVr1OsnCafF6cZJhgoB1ebBFLn4JehwqFei16lzC1FdVkl3rY3PMFEphCOIQ
LmNxoSssCshY8DRodUoTuZysgkfT1JlENXgzhkEsyrsDNIC2FVbUJcoD4wDdp23U
be7YAa9eb2bv2pcfIFTv0/lLiqzAxPpi6FAQXgVsGzPnrIO9Fd7+crEKh4XjwlZf
XiPbcGhfxlWrb7+ZpepH7tpO0Ol6BuHLy0gBm6BwPMU+XOdoGqxCrnyKDxMloxM6
Exo3imDCqK/J7JT41GYzLvfc7ZWAmou0//kvou0XpixTpY/62Llm8tQ0wuMc0eib
tXxrdQzw/crwwOjFKKRKJxjkvan+rfyz5Ox6FgS1Ub45D38ojDpLFd8+IuW3HeRd
ZkyD0mww6n87GngmOWV7OhEmWMTzPG/G27ocqYJOUDEmraA0DU/9O35BO7OxDJFb
2LlN81HrvFOv5RnJ6gcja5cDe36EuBEBTS9wCLSJ5vsdv9gGaWzMMGcSkMbhuzoS
fWgF2u5NjfYP5VBbjvhnVPncTbjqtJQOzxXL5e5UW4lFEJK5Ji0LdJBKQLYlL2nc
MA/q9yUR5xl0g/kJZMA8HWJeV/Jn1YUiBsq6YIbjD/GbediysGfe6TNN0CoeNAhB
zEyj9miZeoxmWTdeXecR8vYJ0wDuJkvBksAeTNBPWb6BWEIMF315EBX0YGKX2wMm
zvYEBrr82ynQNtvWhsEsf+TiisVoRjGg1wmDlkmbAdl2u760ax5H4M/jsJT0VZEQ
KaZNveObWyvQhcqr0DBME7fm86uCQQmAxuAJFUjX9vXl+dZeO3HQ5l29IWe0nF4+
Dt3l651Lt24aX9RIEXinO6Hwrbvv4dedy/YWtdgC6MuknZdbfc8AJP7SLMDsKqFB
iYO+8bmF+K64eUxO6iFc/FaHCv+ZMeyN5lPeDyewmCTqaiCqGD0fljYJSgrq8oRp
YkpIAb/CPFQp1h71pPXMX+X48JPvkldIA2FKq9fU22+dW9Gekg/NPiOB6pnMGiIT
Fd28usREg6MW7pzamqaSmYEpKIGooBBNVGxk9YBCwLTUrkaSIAjJ3AFaQrsB1dpP
ix36+cDKcgaQyF5jzjJ8zBcsaTNK/4ZJqMH0WI+xx4TcSL7l3Eg0MzNhSSpO1TwI
E/fVwbQ9O9nMtBHCPk/oeg==
`protect END_PROTECTED
