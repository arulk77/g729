`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJmJbwa0jQ6ETPkittbmPaOXoszvQ1u+RtAYcPq9hYxO
G+ZMENKTqdlx8sYpVkoVr+hEBORETyQtW+wOG2oDUEl7o8+IOYBRWkJ92fnnXy5c
JTCvyiGYoVtpaGoVCYewA27SH8e709E9j4XxnwXioOIPgledbhcfJSl3EpQLiT6f
UTQxTcYdCCyeqcCsmyOwTJwt87AbdsI00O113GhBOQAvqqsIr5RqM0AgAP3MJj6+
VtFKAD58+7YKhiDDLH7gcoCnHjeMyTO4UqhFtGO/Zy8M3B/pbatamQ+7/FLqcN6v
LvxB+78IYHBwirwkEuZn6jJ8UgBg/DB0mEmIvX1y7jYuJJaSM4QF5XnAz0cpz9Kv
3UtKwdW0MBuF75yaKiPyMfd7CA1sytgoMpRoH+SXmkDA8tewGFRHrLy8Q5PN8hV8
UoQxkBrgMU3q1gwXtt1C2zjP7+PVDlTm8pQK+jSIL9ezi9nFCwed/AY0Bu+Q+p4h
2umIwC3i4kbR3cZLAgX2xLi50MSR0Yk0xmWU29pqyE5QavAjYbN9Z55rETOv//h4
w2OkVwFUuJkobSwiQ59FMwKWthFnY59cKuwUbI7dPq0GGoLUm6vAsIx44jFPRX15
yFdWk/1V6fIf3O/FaF1SgwV/n/ZyPS+ODS7zi8137k0gag53CdRZ26tzg4Uzw+1l
xjcWKsvg2z1r/Z0DaouEpyqqd6cEVnjb2MR2EX5ts1x+7Jk85HlLV1VKjldIniqS
TH3C7CAIZTdnpcp40Su1elUoHz3Xwi25/1rE55Tv7QeNiUeXXGVP8lhcy2A94jEh
97xxT1dZoOZz9/WlyqkZABmDEJCLERv6oDiY1dS7V6g=
`protect END_PROTECTED
