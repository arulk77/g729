`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJD+r3mirP9/1PpN/cOFCzuB24YEFq3yzjEFswTyMDR6
yvuBK5ttKSeT48d8we5nYSYhC1gl/FZ5DfNYBgn5obTFCMLk0YHvu/5F12QS32HJ
ycLMlZP9a+LVT7uRgUb6av8eO3TTyxCDMd2LBlGGVIl6Y8liCU1SqxFXO7la5XVa
oNU4Igqsft6HqJxfCVHnynevEwSJ4hKrTywKSbtiNzzJHRU6wmw7iADbVUS1ZneJ
a6bpOKftESAoiFDTTdbP5KHV5HPrJQmyRRh05n6wCotETMI98kx8gk8PcdrUV5Su
q2mkQ1qfMPaSVTMjERJAjtz1tF0lP2i+Bq2BKSwp7uaHhcudWFrZbgtH9Q5drXeK
8MZVFFjkznUFY0d0McK/HkQXd1DzL/U8wd91H5wKexU8Ihdk7jbdMiS7BfrShU72
`protect END_PROTECTED
