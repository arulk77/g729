`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
fTQjfemEqhgk5MpiuGFNQoYFvYnYDfZjCEq+CAxoazBdPS9VTuR9mz3qqSm9NCTp
+kXunOpqLm03AMADm3C8c+KfzjrcKaa9j9XmrnNUTEmxCL3odGmrMu9JkolzV0pE
mJz7uMU6RIz3dkEPNmrfLMidKsxbS9I5C62Xf08W8+CRv5z1+nai+UPzSc4bNloU
`protect END_PROTECTED
