`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLNqir943U+AELeZuoQN2K0fLaMDLjKov+70nAdB9ykM
phZpcXjMtmhNUjHPI8Ve0bML16tk/3V1Pc2lsmsJr8aSZo4tCZfSQkFtPrFkd96e
rahD7UrSF1wrVyoxynTAB00ktOx1HxB+j22/aolYJmNjLKOIiNFwe/xGpE8a/ju6
hlWECJb6r9f7aWyXMCgNRw==
`protect END_PROTECTED
