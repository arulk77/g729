`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Jk+KUo+epiq/sqe+t9jMS7T6sc5FuR9zl1i7/Bls5R2qJ+t9zzHqIVJu0c379JfD
EV7R9pEKHIHLavRxyZL+l8PoxpJ0Y+OL9e7CkOCstWMf7cMLppGsgu21C2g6Jt+V
+sEsPWhUP4pOZPZyDIMKMBTk3CKpD2gwFORxgXwytJaFupUAC8aETjaWhI8wyssm
LwtMGG/LiMAentijvrxOQO0dle2eHtQoXd5N1BUPyxaDs8K1/qlSFLtuqkDduiHc
4+tOxbFaQ+JxWQpExsnTNd0HA+HxmsPEg9veI9vVrZ7Kcd5EE3nAp1KqnhxMTtQu
criRH88gjBZEEV9fV+hukrlpAyjCT4ejfZrvEbfyjqAcVwydH9tkCbdpGk38cvsu
opu3DdtAO/Pz1FBi/FGStsZnsiclzZqyweURVAwgG28=
`protect END_PROTECTED
