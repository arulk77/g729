`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aVV2EeJoLqewYl0KeaoE4kuUtSHH+X58U8FyoxOCV8VJ
xUyXJcvHnCmYemE4e47peggjj9OhGkycWSJCcQHUeijeHeWFqyp7q2RJDR4OpqtS
ewYtLW1t8x74GsAQuOad9si/clefnbAB+ErT5JLNCjlTeK2OR21e5ZEYSrLHlKH5
rk92DpzjuV+aqy54u+h+1Bs6KGWv18WbMVkdTk7ok1DloyR3hIwv+q2mXM4LI1dC
knf5kBY55jiIrTUJhJ/8ykANVEdojAa1l99/pOFKvmnLZhyA/MJeQuZj1WyeVDPV
vHBJmgohSgu1UBp3vWmf1hBXNpiliCB5ecPmH85mTlNAcbOFQVE1HnMFI49B5X13
EJ2ZSlTDGLoBZFstcv+p4ROG28wqEVymZ55e+usmnOlknsE24yciogRyWz+mt0ut
+mzOgUFxDF4L2wH2+SE/6OBiPkDOY9k0VURRn5YvM705Et759nVrJTTHpq10xdRh
qbIs3/bEw+KRCtmfUOktOeuEF5E7NQp1cZ4LJ4L0r4Ary0+5oa4Vv9HraXZ7EtAc
+p+Px5BZmHkfB+DZDdN9Ep6YCrFoeI7szzqIB7Y4lPRoMl2khn/OAu6hzYbdHvqx
hW7HAETePg6UoIetgffPmv/j7c1xy/vjm+z0igsvmUjmWgvKsEDVc/tvHSHtsikI
4ISCDl6b95M7Ie4oOsn0qD+iKlODD8MLMk8d2kiFnzgHaHKVNIM1B0RzlvW0px/S
B7N+wICDBibZir/Eloa6m6oJS7Louan/QYfXTL04P/+o0VERMv+HP2jh6l7YWJVd
MrXkRxAecNlGi4lFT5vrIVWwIQvKTTVmbVYrSJ/a5GDT9TPUzYvbh+Hitx6Xz+0w
sgcQj4gSB8oSerxBRCkYTBqtiMZlPbCVHT+Iwzq35sfXrb2khiLpwwXRHMbkKHjo
XyvNXK+KngWtFZnrrUlqr2tYBExtwAG8r6dhJYkPw0odLDAnGbAJKTIeI3eZmIyY
ynquQAeWzyxy68uZvAkf9rVDMFB3RjWhLpiDEGk8MpZdoF/qESuJK3xPTPdIBjfj
1AkZRb7zZO40N1N2oGJY48e6c7k9e0YRpevhJIXNpdVOsi+nwh6u9ccG/FwCatVz
nMQhyd91xRdsCSyg2awijWxSbw7F3lYhuvQ3+WuhpDc/w8N9WUf+HHlPFKJoUURO
1hq9JZ36fL5WGIIYK10+Y9/z8z3ZpUETxDxV59n1oSoR10EKiroH/n8Wjaus5kOO
b8Oblrx8BAXCcxYGC2EButivo340cxgJQjHR9diL1jRIByrtPjrQZX9SrlkWXRaO
peS98IggDzse9N3QnsTKAuZxnN4q2/mGo9tsotTVzGgN5ePzKDva32D6IbsbD3zS
w63pf1WP5SIvVRzD9u231n5TYuhfpbwKnkqua9Q17jzC7LI20nWcol0Nfa+odxfZ
ftKUvC4gIHCFB2lM8t7GrWmn6UKy86/0qUzd8hXlDLZNp6PMKwqWWUyFzyDRcgwd
3HvKNi+q01BtXFFjCC659IpXtzYyo+4s+REVt3qZvm9fPPxroRt77vDCtFS+uUZe
lXKl+e4jrWhxY2OlsJeWfiCV6E0RSok/vYi8nK2AfDz3ccc6x4g5X5vLdfdkdS48
19ndRsCX7B+5DLhoy0AV4MQk85Kk2MxSS8SibtUTCMZXZYf/Dqi8JTMSc7f7cMeb
W7zv2xjIOAd5a/A2M/dET+cK2yvR0F+m+sdN/3782babxxDngMewaKO/RJOhRGoL
Ryuar8B3lT6ATR+X3aEbFxGgQDku1ko/mHnMvpQHPM/vagBdVd5WRfIgV5MqyC/k
pqEvp2fy48CVFQugGQK8EwtQj3XdHhZDs99tgiCXfyemJt1Vx7oSp3X35jiPNH1D
SWbXxkp4GcXVd/cQcFeUbMmagoXPkNbt6WbKzBzWBUjkcZ6BoggHT/ULU2CZiVEr
pqUv/InaW8Qz2ZADoKScQl1W5cpP2Bn5IbrdHpKB4RyU7Egg+E8LdBxFaCzsyKvT
4vUWGROWw4jzgj6p80boqPCrZ6M1FGoTLlmOPCovZ2L4pDVnnoleju/IiMDy0LrV
maCRf+z2Za2xSs7G8ZU6X3D8cPidKLk8chm9Ex9l5/UzCBtMnl0Q5Zhr/WSXbFR7
uzMH9ex3LlR57WCfPFHtiHaq6wx105d9JWJBb4gn39kH7W9GaDZ3MbJgTZS1WJS7
vyDgtvlHOuK/v+AnFUEvdIw0zKQ4E+XrOSQ9tH3ktnpXOzNnQT9n+WqRMSaY1elD
GsZr9G48hr8n/xcloLRDCcavQ8jhQLOA7kjnJTwlLcLyBV+i0cquPzEBIGN3oJYK
bXVBnZOw5BaY60AyUftfD3hWpsWYayAlhA82K3dQGHNZ5UuI5ag8n3fiGNUrV9Iv
NQwY1b0+KL+BkYWA2J8AojYzOB1NnAKrRgC6Wp2p9I0z5mM7xHEvyGezH8rTnoMm
zisDu8qCoDLKYAJw0hE+xHTrGRfj6Gq9Ne5RzipgsjUvhB0f5irZ6Q5YUUtG0s31
M8L6Ma5GHGua7aPylIopt3r4E3M0lEWC4T+G0U2m+aYqH63jCCqygZel1sTGf1TF
54gGqjl5L7WfpD9pky7qph92mKDF/GPKQkTCaw8Jz17QPKmw/myVEMdXK1Q6qadR
3cxqjQm+QFlMYDAW1NNxdWJqvLAX5RHblk8vSN/avC3xoTYq7VPJN8w6OXnyrC5+
9h7QRQ3ouD5qBPOuKYVLBcEN4JAXm6Oa4QmBueNai3dO9Wt9OdadjiZLUySijIjv
amignHly5+n6rjwYOR2ZCpyb4xEC8JwjTTMT2Fs0fiNMo3J415UjGoWJdFGm17uI
vdylkrmxii6kq+1UFIQTBEIUUMpGH5i62C0qwx8LVHS0NzCEF82PFtyiHCFwJ/RN
C9TlZq7307P3QZYMZXjZspMKTCm8/BMRK/lBI0Gt7lBBRBe+1c+vXkDsSQEUsFZx
laMoo5v1+5JorTY1KwozqNtwqIRXyxtm6t7yqCSPY9ysNeH6LANk8hkCu5/o54Py
RilPYBmkr7ING11I+ACSFHjXc9yN9xAeiamcUVgudOVNDqg4yQaBY39Vy7cJB4bI
1mmfLVIWEBcdB1Zfl7q/vbNGNjaRhNosY+ghYqbMcH2E+Xauy0Yl1oZPItdAKgpO
dNj0o3u5l7goF6jdGOpm2459jfCd+z6Ofsw/iGe7V4kRB+8QU7VAoNEpC9z8Gogv
9mr7ZoSc2kxYCYn1FV19si308f0S028P6qWR2PsCbyomswFCPkNNkvsaVyzqXLUU
L3+oWKBFOIHtFEDjWH0ijVLWWHSpYXZ41k93jRP1JRvsscZ5UasxD0WeUSk5et0S
k6SHaFIpqImdLlCiOCXtbB9yZrbdXB9OHpKAcn49gPrRxjWJ9iksbQKqgiZMTbYx
7hXyKCBO3sn/8xIW2lQAzKPNa7gsY46//eonpESzv27RZyZKlMndNEZ91kQGXXqC
pf9jlk5N0d6wgwnLmSskQCtw1OwOi5oByjpEUMdMq03rJQBZSipObHogfU4Vqkvg
MBPPPH8NM+xWr76tLYx3O3QIJJ5thWQS86jOiKoRNVgb3vIUBdcWGl17d9/Fq9J0
u9BbwrmgxXFthby8s8YCUYqcNtu9KH0NYbIUA5LbhF9J3G+9dSXUMztC2+rmQu4m
fPSObmGn3/dwHLKme47HASxknH3yZtSuiTzNl/ceRCQF8vnXXQ+j3SYSsmq0fnC+
gjXOyf5tddzQdKADkzC85jjy2PhrTycLOZjcDJl75AoCBcq1EhjcOtG84Moqy7Zi
MD5F/UQ21/tS0QGyzFDWVl7Iym5ESYnlffKHC+W9WJ4Mi+OlALtqR8YaIa8ncrcy
nE4AHbFdl6MbgufzupmuaUcQPrsJWLhq4wJDpBrldbtK6smJYOBkThxsFStl1Zjl
klbAiv8NHZsAqwTtHqwW6PnH4X1FDNPWgLBZaj6J/adtZ3csNqO9idunvOdhif20
EecF8OWbK28/hnlK2qvkxbjsTDfruQ9c8n7RXbI5p8oaHSserdpf2bIMqwXkmvwe
/OGd2hHfS4I6ksmKFSIfZj+3P8gQxcdz0KHo32CVF0WuqlGo7DoU830jevklnpx1
9YpxPDsRkh2yajMSKiwFVCyydC+F0IIAetmIYMXX1prM/UrR3G09o8NRlhwlDe3k
A2z6mAlS96YZGY14iauzSTuUba3BWdfWN1p7lYsEhypjmlAVdkg/VRG1EeIDH6pC
OIzWn1S0+cFvDyk/8C/IqsvItgyJx2LXWPBpwBsW7AbXiOeDvFJRksUG1ccJOtYe
SZw4LkrVK3I5x/9Nw8Dx3XufdtL3WDziZf7MGtfiGGkq7lSOe4s/63GOMd+xNRw4
R+K8Zh18yZ4s5zyovEH+Exmxlv+3XNWUWBuusy+b/InoSjYxuGHDzMVohFyqWTEc
VglBWXqWq7xqoVCuiQE7mpmmkNEaN4LDzEj3F+R7i+DobF05eM69VLhwe2iuOKoO
5TML3MAMBVDVtVGe6VOxgxjaqatz5Q7Qr3TTsNvQDZmpXpARmGT+cQT/LoJqruIW
Tgbo0oOMzwiqqrbHMy8bCpsYWvPmR5Q0b8lKmFzgVm69aXTePq/48h9Sf4J/zaOX
B1DnKfYTGlegJthjCgwl2yi29BAbFGs2ZtXdpIljArZih5qpxS+84zzCcmMziCIY
H/gHyKllFjrIpZVBOTMTO+JUFec7kLen5VGS954BrN6OrbbFihnw9FR91dQdsvUC
SJ6vdjBq9d51i4VGiujn6DhnW+l4C6v+M0SzxaBRP5Yf0WzVnA5WOiFfwCv+QBnu
0O3PJ5VhN2OT9mHM2WLc+fqAaxzpPXI0+K3xe5gMiyzSPulNG9TfGCjs2DFteUlu
2UXigxEY+iSSSTIEBIsXuvXtKPwvQmh4PPo1QYQNVWaGpui8CR9Bf/DhDc9yzNJv
6yXT+aLWmfYf4KRbOmmjXxZJc6LvlEFhyw9dYHAX6ePfRJArfkR4eFF0NnKO1kGw
9ZSfpTWiFw2B7ylTNkAXtjfy8sraKg0eJ6LcJEtiCpJVztUad7JpekinqssFkjcA
3M8EqMeCr5T45SA9I8V6TxZETiGx3m/VnulK5PYf12AsA2c2Gm4OxanIIEO+g/Ed
tkcOWHA7qLn0GsTDKfM3UX6Iqh9/70MKgJLxAMJnJ7yf0bkDDmLKbStrTWWAzFqL
q5ExfgDiA1eH5GLILBtAZceNoNkkb1aUqWoORPLXSDASQBBjKdq3NK5IWvPvfFOs
7RFbgkSB6w2iGHJUr5UjcpRd3lCvGNwNwQtrwtaf7BIuriJ3oLOkOp0xaYGuYV/0
lxC3UYHhwqWjUxSWU5ggVeXW+On8Czn9ztNUfNCtb2oB1q3xoc6nQ6yiNFJJ4GfP
raxuhl7tehJbByBRBesxyQLDBGRobn4zCDjAYJjd6wIxN3+aZkF1wnb2/WnUk44x
ek9UTpHjOKc88b6JDHMUcGO6Mkt1BNP7ZunW1K+W18D/2NrpF0EL1rWVdLHzyYjF
U3cAZ5wBHduZyNiNJd7GDcxFIDcA1bdNRNGWiflelk4q3IqDKSQu77AjH2RxXECG
vcx1tHWIGH4rVcbqG2L1p+jA5M4bfMFYxbxfbXcmphCVgg4LjcEC/dC87duZeD32
/Nqk0vOEHZH7WxSCVbBJobSMP9NUpBnbR5iV6mA6fbqLsXqJQbbsLibqBp9g6tmG
QnbgYh5Doh1SvZUmE5XUudGnEGqIv0C9iqJszxIoeB215zduwwwTqRI+ZVO7Lhs0
NbZ5b1IWDrDElC4jGRRMTug6wTAU+cJx6HBA8GSJd04uIvtszL+9fhD4eUAYGQCN
f1LyBeBJRdhnNQ0ScA+phyz44qNGtyR3Yxq2+vaYeRGS5957C9/pmb02S+C2BHzZ
QQOOJkpxuS15r0iG8RSN9j5kTUHugwtnnY1RG1mozKgiyU/dx8zDr9/aTSAebxvi
e89d9PylYkv1JBlVScTEl43lylXCnKubvQbh3EJPp7gLnSMMMKtpNptxdIvjVoT+
BNLmv3H+xhleSVFKHDmAIfNdhVGFoao6B7wvF3W1bPEIN7eJujIwe3KUPrWIIOXn
1+ccPI3A1q+Rv54Rzrk20YhQI7dufXvOqtoSFQpdhspJbEuobgD+3MHzgxawZRzq
9+AQNe/YzOOsdYG0cWqkUlC+L4k9k+ncnoG18rRrQA0qES6MQkYcExV4ZtI+meBr
Ip4GJuHHaajCNyL0GpCDOyOBwAMH+/E+7tZddGgdpcKDq8ip8xOTf/jEPS4/C47h
fw7cFu4+ReaEdhAOoFy+F19bENA994sSvoGTEsI2BbzpEUFJWBw+Uck8um0603H1
n6ALoiUizALkEBldXOcNlx8yotVONqiTDi3LVCcKDtwjftSmafAbI9ZW2HYA3X9Y
OjytryzSb1ZfC0IUTuvsy6WRHw4PruyDQwhwQnc0SJFzbqjd5exK7oevVkL/YUgS
tURepmomZ8mllH+iiqm+5RnAudnm7Vt4RoOG76eAiRGMdN3SAMSwS+bXB4jV2vMX
Qp1uHEoUW75wSdZJRBMTbXrqVQLmm6YwXv4js1wHMQqOAR3vbi4EEtihMIRxirq3
UgxIT0c8iZ3LEx9bOHUzkqtlz4KHlgFAj9uaKfKfr+eoOshYcqRuhGhacfnz0q4V
JvOM6hbg5JL2rAmDeEbe2Ux8h1c+NBRHTmVtDDlYJalr9ZbSqhquCoectDNd5bXA
BPev1b7ECv1zw1xrYLFGLOE4Ftp9shi3FJDcOAsYNz7OYLDY+pTYdoo8gKVtcUPj
+5ReN0tqhDxfwhEd8tBeMZh51O66lFYV2rcBZukAyCSeAymnd4/m3M9xOGUaZT9Z
TavIOIx0i4FSnaqfyNKmTD7wwaZY9xYY0GNtns3LnUatJMAnHvSlu6ivm9nVjzKO
VjAQtK9jlKgjR893Xomv7idjsquQ6RTt5qkxHxYIXd5QVjGfi1P4CwVbakrxzPpD
CGatWTh5KX+9j83sVszKhsM9DMhfTUMxKgID3A5O2YzNnP0ol378vvO5RjmtpGtD
MGZKuSQDWS50r1EYPpuBEhDfrCiWFMqenpn8OU2ETma2DPYsws6a+SQBfOF9aPsy
bqGI0Nzfhy7ZPfX19QOQlrmyVvtxjNoDG3eEkCrxiJtCpnbYTccWo4gB5C3I0kLx
UkStJUCa6wW9lodpMe3VCUcW1lGShLZ/NGkaiyciMoDUWrzDkaPPQhn90ntbOrQI
UgnuDzeT4KRGYSSgMW/nHaHBzVl1KdDCYTC2BD3xBQgVi6dDaeDfbBzOCkUrIPP8
NMraQxmVpCRL1YXCdgk6Tgmesez3NHrxIMh2KO1pMUwuNA6KIBetUmnxWtsWN2EU
gTT3d+QVXsBNdx1YeXYrW/sfOKY4xS3wBIJ8QdwIY1lSc17WYn41INq39K1vTfco
PKpfvURHthnzUpwT3INXMb4KtbrLGxWhzFMVfVMlR/RYehOXFoeTfGog7MdX3AGD
xatLWcvIuA6/e3eFrvGLJ9a90ywWJ/H4iSFJqtXfvWpqwt0Jov1iFOM1pu20B2nA
QaESEd5meAukhLaF82KtEjDb5zVer7MFMmj09oJLrSLmF12Wmdkpw5hRZo3VxmTt
ORr+tMU/JPYgaWv2Zf/UwSxSyBNJbMYsSKBszxkFc1Rne443XYint5OLSm7gByCd
xC/Z/4Cd8vR6Ey+u/85D7y3ebKO8EOMdMCMxTSX/XdRwWayMmA7ZX5VVdPue7POw
pBiDXpUNUNBIHvN0I9+B1GXY/MdHPdPaO1GjsnNlgAUOKUGTgG87v5xCQodUpONt
/MR0NxVqIsqGqNeot3voMrOgIhh2AHT5yoY07O4tEl6r8pmN6xT72lVzHUi2QNKZ
0vqU3OF/pb3QfxiOPVnzOxfTWqw//qjOnEN32r78Sk5ncvnMWqL0G+NtwbmD2Ogd
I+Y4I4Z+FRtjlt0nDnd4uzRaz7eGHU2qDtR3NOkXlRnARlLDxfCugWtJaZpBXQVF
gJlMNn6Ky01WOCNZcb+cJtHi3PiDvEAzRMqfqyL42mG1RJrV34qF3y1cL78uZ9gj
3fxW8grhr1PLLJKWFWaR4wM8B4swuAJV5rlDCgd+DeOg36apr10cEUZU5x0fBrai
7TeqKwhYnMl7mo3HGSt7eCejE1FI+8VpcAXIqrCW68B8sMKrZ0IbwzpRxbqWbqAc
r7zbyB507M/MiwpU539GN44ii9SlMU0bYdv2eeUnLjGJVrRymGbvRBVez2PAGdJ6
RJRIdzYac7s56dTG+3L0O+ADYeWJB7DODcxkIOMHhhix+DfEAmow/TOpJcaa6tIE
Z/Qg9Cj+XxxPdvIbK4RceF5wGwx0aW9g5jYSt2Ho5XvjWL5XBGwD+fpinunjqXv7
xdwSSpUdVwwjFgssEg/QvvbPC1za8kqxUA+HeJb98QsxjQPXu2qNfDsG2Tn7YIaN
9H+EWfn4CKnz8EY1E6l2UZUnVg7YtV9JD3/9bqnWl3TiiuxwIBsnviaPWSskH8i4
ABNv7M+t8R35k979wI/h7/yNkz9Fm0swOR71SipWJP81Q8CpScmvtdoaPc/+xjt0
eLl32OmkRmeoZjOhKNADyLmspQ86bGpGqIC47k/eFoLbcjC5ES4Rt+cqqp8BtN4d
BT2iDgDSfNBhcd36KGNC3OVeYxjsaF1eekXfVZXbXWHzyfp/R4irvkwlBo16uOCZ
VZcmiIO8ANbSTLFYPjr0GD8ZfRPpgH+ApDWzBuk6rfexWjwcQUXvGGjiNApZFU2V
9Jp2xSP9Lt65Kn9c/DIUORvwaZZjQnQJ1zqOrzyfyr7Rz1mtQjSUSxt2BCggPaCH
OMG4T245Me1FeV8SBAX6waeyqTiJDzGmcmtCqnWTYVu20el7CSi3toE6fta7J6uW
yKgd1eaUlrNTxxaOtABU2MFkJmYVVCN/Ny+Lqg88k/4CJx2f7lYhbZr8/mw963HY
+m5GfAi8LfxPqYIgZhfJQyJ4f9XILLjzMRgdwOzrNnw8nts8a2vW16y101VRNXct
4c2R4QCFytKv7di7VwPj6U/IyB8tq4nx70t4oPdWQHTQHEdmUMWMVm2R4bFrnDug
bUaaBZWLbw46s89pQiiExfh+RspSE/KX9CXeWJu8JVQs+Cd2MYtrFGeH3uEGRgtk
pBCXJsAAoJSMVUsx1Iu4hfFW2ko5nwO4riCQBFuZm7jgdt73q0TtHsBYHlKw7sHV
IhGDv+dnB8LRJUTRyL/TOKlZbI6AhvjmI45H8DdiNaJX9TVlqRiDKDk7TMcGGbgl
awft6tGAGa9iRIOnuIXp2G2sysD3j1Z2hVmUqDQ5pA0XwrOU8zlpbOYe9bStlExL
fNHZd9YO38FmaXKPnpwvOJrhCs60sD0OJMHjrUDsTAxv/k73j8ob/V8PTkitQLks
+XrlV12ARZFUoIMPk8Lh2bN5t5Fl+oytQwzojoS0vPL9jEatyz3quS1hBPgrFMLq
O2rCwxsF7C5KDKcGGcIQn2DgG6zf6OBW7v6p9stLwguUgXrr/KSc61MfMXx1+kqO
YWp8WQ6MRoJR2evsgrhKJtMuYWIvVLx4D6g+gz2Y87uFOGaAinHjgpitQ8ALg9ki
bpPRfriXGuWAnFaVy3u+6+CnaiYgIw6wjAdHWyF/2WjtvgTWyQdRHFhuN7pklgyW
R71bZwfjX9i5td3AzpAyCFqAIHQhXjsc4qLF7Q3bPWJzZdcNTTNxNmYpPoo3QsEe
RrBG5suwBDZtXowv5ykeBA4bERdhm7lPLhDRyEBfh/JIHVcH3QiamgO4GyFqDu6F
uZ0GI6Q8MjkYj39rcIit+5C4EXXNTh87YxZiwtkTAmZh0+wv7puduuVOzifktE4V
djw1+oeARHfur3bkNw/B+fI8s4y7726eBawDm/E3HktUBr5njwq81anWzuR7XUZi
XFWf3faASt4vB3dFsikapWBg/JFhXlu9MQV4dQcZOBVsmETxC5LbhmWv8zT+7E7i
sfmrUM0pKkbO+73i3kSqjMpeLT7DWzPQuLL1L+W0g7tWcHRYeuBdjxd8qzgP31UC
U5Yi/iO90lQChLYJ1Ok//H0LaL1EjD60i3tKWmii4yvPHy8ojuTUSA/aKl0w9hQw
QhPu6Cn2T/XgbEn/FEc4Uwz3MRTAJmXKSk2wVqhgo+3HGqB9akKx8IMoCWRcePiP
PS26TMCd32oeuafj5HN5siS7NDQjjJxIPm20RP+Rj7bMv43EKAf/VZAgl2iiCoo2
anY7tSQS+xjC/z9fURiXwpSmxivWvtWjGezclR+kgaT0TpBcn8aL/Lf8qcIz9wQr
Mf3qzgV0lJRWn0FijDCqfNP950QG7WHlwdLZ87iSaS31rS8emYNco0R3dWDR67o6
TnUXNfCjwRBf50nPtT0hMyFf2ei/qMP39UMa6GRMPUiY/uOOhWbT0M4lieE1T2sJ
pgNe0efo8PEpk6Vp5awT8ur1J1iyl4Y0rg3fml2DrGHSAW/08rSHDyKPhyEgKk65
wmEBZzimRqEshYEcz1ffv37rnniZXj73pvg9ArTwLth5TZGDIkOLhLi1iM79frw3
iJj04MSKNHLpZ1HHRv9QNfIkRsSddEu+wmJxMRLzy1TY+QwoI/b8YSsjfE79PsaK
fl+nMB/LYJdn2kPL+ntIFWlXs+wkrFmlJPPeB5XxwAatrd64XsPDH+eOAyFUR5f4
SeMp+zy2QJRwat4cOBiG8m5RLoWfX7v+/lDbH8CouuldVYMUC1zk0xZjr2uj0LyV
HkQP6slUS6WPkVDpRFJ87kbQj24BM68BGL9W1zTeEhDug4itXOjtMUvoCwTj3feu
NUOGAdyw9DeZ7t+m1PXXD+SdAXs941g0BCY9UT+QqPNN2pw3wIziAbpNg2W0oCt4
c95qduwNVcDOr7SxkdAi/2qgpaaKnVnIsI77SjPaVLxyNEgz0UsgjuO5wrtByG6W
WJHItcM9SGTSezcP5uytZHZiDSNDHiCOkZ6B+Xfo8Mmyy4Bs/RmwsbluxmOmwoGF
PxeipNHFRfU3sdvZ1OGED060KCs+vMGgm5e+JZiM27n6W6+KrYu7+tIXf4woDdxV
ryRIioiuTXZJHbtq0RwAdkG/EN/U9PuAbln3nQxXrUNsLL9Z81Y5xCS1mM6khiSW
SIh4c2e9ng9DjXenh63DpXQT0SKTSp4FEUmP5BhVWsuskeD5+YH82plm8M/Y3r9d
T3ViLQsxunlnPYW/Ohj5e4HPIT4Uagb2RN3evmXo8Iu4WhUTbq3ji6AiN3N05kY6
xmQ8quhAGm9n7cxOjYKm5BGUNP2swmzf7Bw6FmGBKxqI32PSor6yBEzwIGxFSHA+
EpZkp1mot3WqHS8bHGuC4In/di0TV1HVX5GP/I+FusTJ3lMuBCFFkBWagLCJgTfw
xh8nb3M86D8xXos6+NfHYf85ZS1JTfdTmunkgjPADcWXn2pA9qfbtRuGvEo1Ddxe
GNfVHpOooqSQ5uRGcoPzlCVeJhBC4gppujVFEzu/hqgFZFCRdx0tMYpMv85T6/Yh
eLVjmNo320h6IYm9LEfsaaf1CGj3EA9K4SOI1oThH6XTwqAIcgIidoazjnXMlLc+
fgQttNfM7tQhRRy2LiUcLzA927ROtabcFQ8hzzSgYfI7ye1c6a/+k+qg+IPyssFg
VhxJMwdAU9BInyUwmuCIBg/mRZuapvv0h8NTtsxr5ZM2Ev8ncH40itWdfMojc3Xi
ggzLdujGEIIpEyT9Gbd+wmq/DFk/wXarzdPZ5KN8lSin7yQv73SX6eXoAc8kXcW5
/ipBrD+cK0xVavayUIXkfElWd1gfjRlz11eRh1hyALIVHAz9v4wQzHWD+Ll8YCD7
MfBL+IphwYcZlMqukK0upq9YTgJrWC5LFVjCt0IiwdQ3GC/ppaG3K//b0QI9bCG9
XVCuLN7VtMV8jXzdXkEVAL3wixy+FGLiJeK6PVw+Cbwf9Ra/X0Qzi3hTb8UIhdVm
V/8YE6WntvAr116FPCzjNPRd8zjfDnHynsOtqinbCrN/cqHWEOLW7N4l6EtmHSh2
xSEN5z1UBs8T9wZCQEVe+fAdizYnYIhuIos8Uo3qJJl9hXAkySUqBeRFpSSEcI7/
4FNx4Xfx1F26LLxFsg0v2RSNHB/Yn1Eq6WkGsCHYPTEYsxBBhM/eYIKj/fBNVAgV
qXfweOYPGGURUKymT7nWbXv5FMqeXfmJLxE3zgABjYLCYlZkSGWmvnhX4pimf71E
I30Jgv4Yy0abNuAQAMKs413JDhXoyNjH0KAAtk8D+YC+hxzfta9ImBL7hFYiyE/a
9TD+9c/rK2tUHx+lk8TXK/hiltiim6nmTp73Me6byGGNiBJl7FTo6WNXc7QrtcQq
IS69LTk4yK4bkVZgcZkeXDsD9z/43ZQ94Bx0M4tmuE/vm201PioDJDZVyQIyWKay
TpeIenrFAVEQXJtnQ3cwwwdBysrEJ5Qzd4HF56eFCCBDvkiru1lKugcqt4HF5gxo
rVqncx0fAKElw7E5lcBUyT6/2tqR/fzAZXo2zItEBcY/XdcLG2YT+/nOstjTSLrp
HPhIEkYsquf0hk9Zm4I5TcUxZ5q2N6r8S60zO3wLoy7mInjHie/TYeszq14nuyce
WzmbRsCnPqfnavlY6bd9ZLggKNQOWpb45HHeAVguDFcM0EgwflBLdH0P16I2V5x3
DrykwWmPAcZnGpzmX3txtjHg2k9BCi7UnJuISc+7NOa+0bz++2uIvSCXzuF3bkdp
4xUs8swPZwf3v4Ys4oAh5iY8rdPORyXn2OXYuNUIKoXXDuRpgPDYKh7LUtg3SH1w
DZHrOa4acINmSyvbZ3x758fqbGgnrU132efW2N3S0v+NCdeMO7IGrlf9McjJ+if0
E0K7G/NqNld7b8/gLqUDOBRb5/OnLDFLjK5v3kclP5PohxZKLup4i5uZ0BK6Ky6i
JXND8hxuLwTSGNEI8t5dqAmo4JQ8YKXnrfTgD5S/l/xTIwUxVihVSPlWwuwrXcIX
wYBYcjH9xD4bR71byYGfWm8RZQMWh38CY/Yo/TYsJ58f+7NnynniAyKmacwU3dQZ
Uqqe67lZBmUhrh5523cgmASR/Ng9soVQ05Xq3YLLUuI3CQHMMbFPak3G16nTLJ9U
KKS+HiuT2mADD8VzVTNpQWNRr4jsdtsYNYRmMFdHhZjS1e4ZF1/k/UVihR2IhXxd
/t6a8ZZSZ+EM6/oHfr6Z6pCILWRcQJC+yRECaTMZ6HIfkLBwKB0hJNYFlEi6458z
XFA8TGC56jBY64AORxm5wWruUnZpUqotKqfvFXieh015FE0dJduCkf3ifrkLGlg3
opr4lIuJEBBOabQALt+u4vESVKC0/wR6Ef9rle2Oio0OyoOhRYvk/590o1n2dUuS
mmE1ASjm44PDFCJ5HbD6j46kLQHNSKm/8hvY7cjtcx6VnFUsRv9cDNT4pyY9XPvZ
YvPwCcJsjvNm1WrHlH6Qo8VzWZxk1gBHrhV8u9bBgLUgCQB0gUfuJ+6GNNqnGLtN
Q2qoBAycBsK6hvIIYBhGc+5NXzldcqPJV8Nk4GxINML1bTtt3fg0UtYSZFX8kMG6
QSsGUbg4vomqaCF3WH54f5EPfPsrAfjzFTbFld7tRyiH8WH5BCdSFQ87JxNir09a
LCVJw8aRZJE+QFpiB70YVudQJhlZZRbU2fVANQjW8ui9LmhwCs5IxzEztv1IY/qg
+BpQRM4svpO351EOHxK3JpGHRs0ee54BcQX4DllWVTkrf2sfXQV9pQQkp6ZjiTLi
B0noLRAgplu/IEOGWuIAgUHzza5pQIAV09xL+pntij1SnUwfRN+GQ2ofvzzt1he8
9kpV36HlTaHaaSNNJQG/5FnLG07URfgx0PBngGsvi9oAPS8m8eJ3XgLGnJefRvjK
Y0sl1YjTISXdkHdEOsnwJg==
`protect END_PROTECTED
