`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHck7uHEQaolyceG8Bra/tDggUt6Th54D1D13Ydl+n7g
Jewf2HR+KwBZmPhYfBN800qcY7+59x5SeEsHJNuv5Ole0n5g5xJBsofr7jT810hp
I4HTj4fXHxn6E6LMPpsOLoKqlwPWYfx4zwWCXHkP1PPsEyjMblhCVfqgAojlj59S
2EEuEllOr+ayik4G6PfQqZRemDRqD1r/nlibOQymqX8TdSX5U5BbW3jwTJBfbMw0
`protect END_PROTECTED
