`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKE6MufQq+sDPFbyjiciXtJ4b+l6LHh4nts7hO4vfhn0
oVBYTNubxm6R0IKtHX4k+8rmiSuDre7v+WbPtKZRRq33Vuj7dt+cnpq4frSyiMLj
rO48rwJrxKsphZbi1F3LbN7XVa+3gCui3RkpMvKo/hmDy866/9mSYrLxOhr2y8oi
gXCI/jX3WNRpaQYXJTO+6/1YgoA4qmYTdryJdjPfEz/AOzJoF/qBPA8N/X7B376b
8Yezbk6l44gWAbVTnEvB2PjqdOnxHEgw2No85WOnJIZ+TfrkR8UyQRFYX0M7hnWV
VRREtMmwOIF+q2i1PJhPVRS+Nj4CnX//p5ZykkWjsL/oGL9mS5mJJemzP9+N5+cC
irnNHwiBeXr5gzNxn8loLEIWKR1hSTYDvBXMf1A47NtyPfdk1fHoVLsmMcYlwVeo
No5cTwAZBS0Ymi5rNZHVNKAjc2NonU/uiavo0eeNqkU5uzdQNA2LpGid+Lk7H7sz
mFoMPZsaUfIEVa1rk/ED1F54BNd5UsbE34xNhF3yT4/uXDum3yACEkLEiT4y07MQ
bLM/HXs8zZHzfDxLwamsg3ALLKqln1iHOlnNJTcmz7DFhHIAlUOET8ZIIJ/DY2Vc
BsrP4/d/Nx10xxJ8DkHhHJSJMa303a+w7qxv38/qxnCiDni6pDeKSVGerJM0Vzk8
XC2uR5lVgJhoQSbZ50heLgmjoyPRuHD90lUcCceu9TV8PUd84i8f7kCG1mEAxJ0q
6HbsIj8rLCq+Fq0PJo0XS2MzQqbIIj6YDxyaEuCLfKAzE+DcHzGfwa3iLxaDFAbR
p+zKMz5EvoKiXoqRVGiw4bmXyT364lUsJ2l2PR3QypA=
`protect END_PROTECTED
