`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
yvURypTqGORtot+CsKHxA1+EiySA0zN/qOlgM3d3Qsa+zEjRZdX2/eEj/PuSXplt
mPq4PavzEmK+TCDS4tWxixo4jd9ZcOsv8cr8ouLJrFDUrSTZdwKy7ZnZNHCbr5Hu
JRY0j4eUXirPXj9zNGwlGJ8+8pvkmEB/KHLbkjXpNN5byRhjtNDFnyuZsW6w7/m8
gUeSMcy8ww8EruLRP/w3/2FzJZf+cEsffEjGA3JRnMlyEwugZUwCLrph7RhFK0rH
sSmdSzkfsMTgqQ3PPizs+7iKCuWcbgQKtWx+EOIofDz2c2hNsyzv2qmZhD9EC4NW
1ldogpJpbl11FCvpt6xzs0N/YhDtlKC4r7SyWiIX510=
`protect END_PROTECTED
