`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLlEF0qu/RQwpFe3fNr6vuUnv47Im42zxpj5cKyOSitW
M0C3z6M5T3hgtaYlyWnsVCqm13W/V4LdaXcE5RasjwT8iavUCvs2zYliyK6JGYAj
fxdesRQpGX1MNtUGt7lukIACHeX7c5GFUowacINCAZ9SHdXO+JvGEpVhGbRb+V18
uo4D0EGeJS1g0o/1q3E0o6gjKJom2nNU0nsqvtaSLHTuN2fM6Lm2b0kAVxHqfwRn
`protect END_PROTECTED
