`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu47ozPZ/go/wkoT4yUjVKLZ2qlrdfbTfcoq7irqXsXI+V
Cogftjc7uMPppgHcX/ffkne9ivxgHTKidiOxY9zcFQU3Lj2qRk1RkMhIK+pSj7UL
hBVB7ru5i7XX82a88mwG46oZuOS5sI7vUaDFNDvrPwJ67km5mfPc4nq5wf5Ghg3+
OOdCcpBQ/yCejhFDq805mPSaMJHo6wjH3wOdwfvHcpe2ALSPcSkkfU3YebNdQ1Ko
wDAxkoDeWzhvGGit/A3dJ3plYRjsjgd8oIKVamj02lfGKw4U34o9NMZwdcM2b+sG
cngavIklZ9P8WCfZEvUi/g/IEsaztjR8Mxl8dVgNIk80vfIEMxeeRMqINZjx/YCG
HCr7iAR2rD7IdtqNFIbVdw==
`protect END_PROTECTED
