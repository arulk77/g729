`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j7Ku8Mr+nGCSWc2nvLY8ScmqAuiqzPLfn/aSvmCh5lORIaXAAGheJzsC/GjrwJh8
t/kO8TvUkTnv0+nvy1pjwxkbL7eP2hhblhcoc4/vuy5KU1x/c+qWxvi0DMd7XYkl
CPLMPupihUDrhbklcqWbKlz80of0W8bhR0/t+YKyiXeiwlXbwsFzWwH75jqG1BKq
qh82kVb4Wp37EM0l6odoqw==
`protect END_PROTECTED
