`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKM63wVd4dIwZuWaN9rWr8Aq8vRA8H3q0b0f9ZPLc9xy
EIlvsQ53qnIQ07QZhE6WTuLzhFZbPqyDHdAYmWKLrt0i6bYdW1unSLndzfBuC1pX
ASIvkaGuo3ymj1t4gkLqIHyiRG1IOP8OidpSWO1IWRELqaVKLLGM1srYWk+EPXZZ
uK2Ox/rj/GE7jPOWD3OfnaGanOyWHVAidRy5hKkBc8hSl5xJqa2ddWQtcnjGdNsN
UdYBjYE1nF6fzG+AEDDvc61/KHX1dq4uxrtwhOdWoXRI6Z1rMVTbihh5W2krNFH7
MIk3rXt+m9jQAO3PRutAfLwXB9gx2zX5d0ojSyMadpFxAYK3CZ7YNnxydUjvkx+v
WXqlfVzqUrFsgGZPRPnZ/3uNQ8YTWWGPfPJtNVG0VDqv9FWG64n90BFvtnM7GMIZ
9r5dvdfUadVESTzJv1+S9XxdRv4R+s6+C5LtGMmfNmr1bYkkYQuZv6wz+aPaCkq3
`protect END_PROTECTED
