`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmN7aesYxOYlNBLEM3xdoN9shej99jabLwJ7Efw5wNpOJU
7wRor4t7EJypHND82aSE9hW4BwFkW1LIVvV/JPioxjyBRFUKlTEM+PaUQGALRYg+
euHVAWAAzOfVsa3Ao5Nu88atm0xzYaZw+2mj1NvGWQMopl46WiG4wwXYMSHEZlw5
f9JZbH7uCAnG2EXXBqv+FvjcJ2vZQ66X0FsCJgU1SeYeq2ae0zB84guLCcNIETYS
ADzPPuzltW7dh2WcSHUyEBiiVvvlsuXYRDKb7I1kDioKgQzEzDODDjFPDtnbtgBc
niTP1sefzjF/vokOf554z9WrNTrq/AV6cJiSSoLFXqnwcOQ9YkxJaJaGA/0B63gS
DGO1PuD61iczkLxW7BSvVR58N0a33qtZw/Q2V/1bNNNDup1HwTgHRy8rP8zW0l5a
s+HYQMg7lg5/g5kbIHZ6TQaK1VwRUX8lCIrrvygNMerZV43kWwcfszebMH510AgF
bQuxcNp29VdEbii1G7eYVmkHwrsmJbRm35OrzGsuCKZxhQRiOZTMt/Qy1gyJ98Uk
f6PuD335NwAV+n+7gQAUaxCZPiTVwF5Fs0f+ob6SYN+GdY5f903Zzu7Oso6WcQrR
rsdI0uuDNWq9eT97Ap+SNScBM6qiMcDCIcP4/8Fq1hKb/4AS2EHpPZoIPWDoleke
vDXpmwU9+YywB1rceuo/GC8df98RWCXu200GfCBaf6/82rKDB6Vq4FrUNcVS0brd
FrEzjlZs0KOIsv+e3jCWXJz4BVCvqM6ZxDh5aFriBmmR0DOpESulFyLAjep+fwuN
rwyv0eKAjNhEf+wLNNayR6kwe0CRR9tPn0laZo/AstnaE39Ra59Po81mohhVG7ct
GAAOyTbbmV5NXGI5c2/HN1o2XhBRhsYRnxgHOy5d1Nbu3zO46oEwLrC+wrs9oEDL
wkM8j+szAINRQ70/BqLlZolpE4DqZ+GpKUJwOlEpUFo9kymSx8YExaaeQlH4z5XA
ssn2Zh0i+dhQWIfezKMABui3ACZk28siuq03mqHnQxnpLgPtkTsUGY/4AJA1zn4z
sXmy2fve4CgR/nbF5gaRlq5o1JfHCCgLNR9f65JxhitejqDOUduIxbnw2DG7fERd
ICMUOXFAOftVd0UO3c04+KpvR0mFXyclkm58aS8wzqnAm0nwZtYmwn4xqcz980/N
zKLo/gkE8icwhyILh2idXAEXNBMzL7DbM9eUSslwfrHpDdlAZl9MXdf0Zl8Lexc9
m+ZGLVRYA73bsthHGko40BRKwZXYXsKC8MRtWXXSu/mXQH+9+ey/OabK8wdPL0Fb
m4F/hw0wxEZ+ZsL6F8+SbMhdKNWQyhrtPvuJ6kRmRuFHdsDtHXkLIBhY7+J/GFNK
a+HM4pjDFgA+j4IGwv0wMcDDM6IbV4X7WL05NAaHgSYdb8gqrD5quUHV5B4JUlPv
03cpE0bwAuDUx6iiM5AjLPM4ol/xyOg3hZn/vrd/gu31gbmhbAeDWBtQ8BazZhA+
UenYvSHk/dyvgmhAxOtNU1eK5bn4JYVTc2v+glSAfiVjk8iDjbNatetJZE6Web8E
ZE6rvmau+QwYUT3j3SnYgKakYAWiG5IMZBK19APUu2ycZ2oVJQ9fYOffHjiWQqmG
pxi1W1kK4dKt6lEV4icGkFVsPIqPf+l8To4TgkhGOfHONJANpseWd9ModSLG5AmH
DKz7DoHi8EdMMo1qH71S4UPuskFCcXR7ANu37FaJYdj2KOTdaRJzX2WAviMNonRx
H/h9hCIm3FMMABg/yWtSH6nD5IYhPTXmgc7X6I/R2BXZcluCpeK2zXGcjofxmUql
UF4jlAFD3E5UfZ+JeoMfFYr65VInl+9TpXcRos/gNiNICEO3GOCJ3wZhdG38I3XY
h2QUiuSkhDBfyfz9131OgNRvtxFq7XJaqn2Vqvm6E6aB2eZEBukkG7QMXIH1YhN/
/nYOAXLG+Av+WWwybuDDvb4oZS6d3kv6m/wxWe7IZcX1j/kxkqyieB6zFOrna23O
fp6MHVvE9zPNGoxI1/U+m4f3Gxv+fJWP67dVlyXwMh6EVa4sEmyXbOLnUcZaAQUn
fJ8ff8FFDi6pu+F2UWMH0A/ijwoVdhpUGqax39F0YJuwmttKxPnwX6ehyjkNlcmw
Id/xpaJH7j8Za7BHorRaQQUJ8Tw7XXATBTip2SW7xZi2iGd8mUb/RJRAbsTIkefn
yVH8B2oAkQfqp4lK1fTgdGTrCe0CGR7XzSFxbJq3gD3OVcqVUX3fbBuCissZC1+H
AF7F2Lglqu5i7ky9Re9jlOkZ49yb7VVMWrPKWYV2/MWcuzEvSWloxLyiP8oSDbLF
P+BDWufTX964kpJVq+fYZ4Ta9yJ2b0XL7N/g+nTD5MKjfDGQaHbmHUWCboeGMDx/
UVL64wj/n98YLf0tGVvZ5RZ+O+UIhJV3OBYlA+TjqP0TmeOA1xfkq6mdW+IiNVD1
6pfoVLFh3ujyc9O0lgb3MZDmXpuYrM2m6XUrPLvooLeeekHpegTnUf/JQ7l2ptez
N3Pubk+Jp/CRCWznI7Fu5Zh90bnXyxI5D/nfHtlVpRpiqDjLskB9BzJfw3es4Doh
AhQbbSMHHtjhyrxtNPjJbNqmg+jw3Hzi6mLkxcSvHfHMye0Ums+8d0ISwX00IasJ
eCtoQaNZILiUxh0v+KMA+rileOV9rbQEPPShfE2CDXEiahXtI0TCKuSaIfYzBxCF
IY7xnAWRMNH0KeIGD6f320uI9ZjywauCZtO+E5lih15n+NK94BH26UuD1OMW+8uF
3oDeWtbaiAyH1lvltS0qmA9H5Owcn68UClRLdrpaZKMDZYoRC6r6INQo+k6ETonz
/F6JHeKdWrvaVL58gIBbsKMVDrqRhZzvdLvKx5G0/qg96XQKVLf9L1E7zeeOGZDu
UH8Oz63jqwqjGWzDQHwI6+Ex2PjRocemJ2rY52/wLyYPco0HT7L/4jRV9+RuXkDH
8BOSF4v9KmhXqqi8XtG9BmemhUdG9pul1IfEtH2GyacCVmu6ZxhA3+6uOkxTKSAs
AKcT6wDlyf593y1iqXZG9L25MjTdSZIb4V8EuRadcGtOxrk5gfipkurn8ZWJEoSC
yfxN/XhzvvOkfnQMgpjSHt5LKNo7dNjVIsz7hKTwl5ARgz13gPvm1M+iP3c2kTVP
3MrQL0UhNpeawaHMSrA9HJhvwJfEmcKyxfnznU+eCKcJORRuPA/dgFYGCjnowqST
oKg7QwrLtZlI8hZdFY5Rezp1ZOEdQ8BD5hWLy8uCpLhw9XW5rAa/9JWzIcm18x0T
Jhq81ZF+nNIKp2ngn2kaalk0K+X1sQqMCrIn1KemCKTVdamgGp5Yqu9evCtmIiUs
LAvBv5HKz5GRvqvB81jpeDHxvYuo5/QjV0X2tc3jAf2tuLStjFStVUYwGN9L+bf1
`protect END_PROTECTED
