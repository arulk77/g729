`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
vLVmbduiEQu7VYBRCRBxQ36MeuL3rcsF8sFq29Ma8psOPLOv/RxD72RScHxd0GYS
OHju4GPmeIuVQ4GUma7XBoLLPg0KRXp6DEfDOwVuWdvjoJATkqq94YSY4aGLK1d+
roHCUL14pVtTMpBwGNGLFgVjJO46/oWbsZMUc1MGt0ysWd+C1tXPT5V13l13LbM+
fPULWk2irNI8JsVb9IwgBfC65ZlV9cKxyEtuc2nEinJVQOtac2wMhAOzfIULgRap
AbOBzBuXaEs6SlQO1IGU5R+IUf01dXRAPxVjPpduJaFqbntC8fjPkLK5lM0OGcm5
7SX7yOwBpT9wxL7StBs/iD0OBQ4JkFV7AQfP2/DRGxM0gOIVwVXweafgs1dVO7VZ
WkBAQu2zuvM/C2MaJI6dcgjyw6WgxyngXoegDSX9/zS4Cipn4Haa24P+SxouBOmo
`protect END_PROTECTED
