`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ab3t38y2wf5+qsH/48ktMFKfT+vit++5XEWaCjG26R2O5aC5MGmnEzO80DQqPMVb
o1pY6OEzwpXOmzYUcZFWyyfM6huGUS/bxLIRL8xJfzngB5cfTmrJvfjAWBfxcUlo
001N3LG9h0gTusvajSHimQ==
`protect END_PROTECTED
