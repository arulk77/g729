`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveLZNqVNmQOC9DMhE4pE7PBqftMKrNZ0NH/7Nhe0uEOig
fnnnJgbno+xgVpZ3B17j5xiRjKxhSzFMR8EzRM/CORiatvn2OtUSV34ewn3MZvTK
pA1aMJYT3cR/gDCUFporcAdL8Dx0XPlTs88y1A15qje1JqM3GCxMAVD5+8RKMTDc
jMSvC/x0Ll/5ztvacMO0ivtcmeuVGcdEdvmIgaTlHPWibO7ZhOToHICzMvt8EBCz
0PSYeFz4aRS0xd1Z8Cqc/sRIWHNJNeDq6R5bsRQ37zC3zAUyvOV8SRYMl6g4b2Ag
sEsHBRq1I6awNu5STTCyXVAJovlflaZKtagkRTtcButg1B+sOti/OPMtTje6OHm0
IY7xYAZHNH062D6QL4RrPQ==
`protect END_PROTECTED
