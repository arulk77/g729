`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
upvJO7sumJI4ubrImT63ZWAa98fG2fQ1H8l5+Q9+vr8VoY9ip2UOoz57upXCeHOB
xWjBROaGmgsNRUMkP+xBT16n/TMjVfMOCRbTY1vtd6wtNRLrI3+8ojd38zTM+hYr
mABvIiQc0ej+KXKgJnSsnAkZXkY57W9c7s/VNZtjpJyG90YycpIDUT3TBTlm4q0g
WJBarXZqW+R12ezjQTc0FM89s/6I1/37fuK6UHJTYI6laW8eZR4yog/1jV6NECW7
J4uevrW1EiA3OtHzBs6QnHsemfpAZ4exHbj57ULqjrNgQZC1Z75CC8EgpYFHdBwd
1k0lt0oltZ+s60h+1C1I/PQskzzwnwcjwTaRHXt/B9w=
`protect END_PROTECTED
