`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu45vS7TAg2ovcF0r8mtPqGAPVsozFEOR1ovUoWxdoQ8aT
WK0sWWCeLYlYOKLh4SAg/YGb4cS/WG7+er+5bg5OGmqmiakT3nu/CDI2qhpvdoAz
hTgxa/Z2+eo9uoaYnnNV9MZIeehceu88a10Ri2W+YwsDlSV9oayJb4o/QS0S/J5e
iYqn/Zn/VvZLjdXJoYAEf28xZ3zsgfq1OAbM9JElWTLMkm78ENaJdBoqr49kFxy3
fBx2j5H8HJvE+275PhqITc2Vnb0i4y6xuoTQxck9/bGsPoJpYpj0VEITbntKPQxw
SyH4auYZqCAY0uMrX+wejA==
`protect END_PROTECTED
