`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxvePoqgVAn7fkLgcnhVd7Xwf66SjXOK37gxsb3fSRx2zBX
Vc8LkVpcY9f43Tcind9+9ugV3UdNvWNqZlo84LXbLY5+6dlIQw0UhBP482NW3n+8
4IWbx4pgGjflmEdYwerPzBuh72sIWoXiykOy3fOVKX+4eevZzEYRfHWUp1kJ/Fzm
v76vuIbXOqfzPP+A8LTfu2UYZFGnELgyL0nF6CogGBY7hc180AD5Zrsgc2Uu3SJw
`protect END_PROTECTED
