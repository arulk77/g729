`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
Hrm7LaE5cXw3wf7cb1xs0kZMbmTU4Aq/K+yeCmR1zwr0giswuyckdbBoIvZ0efsb
DCiIfu0IfhP4H4gU2QKWl1IFDLrjAnyQCEmgGIFqNMCU11zbMrOXOUj3Dxsb5XAd
aiKOxGq/aDmrsRAUPL6b2qL/qLWdFMhcM+Ctbq5PEmvVYlZ1l7UZOc1aKy11rdUA
8MQeg31ZoCBxHCLKslhv8q/dqZt21o197wPD8ZUlNlklQdtA0CwRb5hNUhv1g3t6
LAomVlcoz55Tn/WnOA9JzU38DL+0vrcKP2Q7hk/NxCLun9FT1/jwZiKviwarn+mg
mzAFuPT5YG/X3XmeyWmD0CWoD87/qoQfV1BbCwuUwGGtu6lrBTPJneJuQ7TzB2ci
gSvi3Eb5/P+mUdRSsnJbCoGCm11c9hhvy0dzTYhFfHCknXjb8zrinfVJz1S2Mz7+
QFQYERHtYB6k/bDnpkL8PH0ACklBiTavtZhH/2H76/4=
`protect END_PROTECTED
