`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAyzY/8ZOEezz+WrqSDBUZKSQlUXDGaRUmb9ZrmitFTL
oU4TWYTBsgS083ExNMTyVbYf3EAIzN0pH7hw9ZkkwKW6aJ+ON4JA0BXP4m0pFi/f
916Utpm5VzNwBVYxlVTV/YG5HZ4BDrf8+F8M1GHcX1co+cedDWyRVAapoTnaFWxD
RQGtffGuRaTjz4OeCkWGdohO9kupP0OW40XUPuNwbTf8hMTm7OinDKb1p/mC9eyG
+KqJJdwcBYOCrMmevxZS4bvqePDr0MMmyh4Thh9/nnA54uX8jDaHLWRZ9VT7tkEY
pYSrIYiY9lLlDb/ZRhRwyOPtO8RdiJowfjIdiXtugUuYcti/K8Q5VjJECDvBvCeZ
4UqYcsAbFfUtzwo/UOUkQnoKg0zBYLf29XXWGiPwCEwBmqw0UMcbdpOyrz2l44ed
9FOttVFcX7DWwqTr0uJL88kaDiTAyZak1oEYdVuRTJQPUzsunoEvJyuYouAyh7Dy
1EpwercByOr8d6/hur5WLjfObwNB6yilp+Wb41zTXJsZCJL71ZMtSZMeeBlCFBkp
oMJmu1RBYI+zwiCZh/wH8TBkEq3T9Ny3Tvvrz+aeTQmoBO6JwwD3WGZxDn/UrDwv
KiIYicqEngVtohe6P7QMkLTfdCVzf61h6Mkd4GfC8xW6iQHMuWvy4M5a7/Xj4dEB
9F4t/SCaKjatzGoMPa5f9qfnEEeu6MZqJF+bez4UVqzCSppuOwsnr2tQ1Yap8bpA
62+V5ZbSYzhC+wmZrY6ygQP7CxlGpKBJA+lts8EMPJHw0s/hh2Bnw2wW3jUcZXcB
`protect END_PROTECTED
