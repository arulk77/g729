`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveHQ/WfQUmZnXBdScaGd99m4AC/F9F0mJ3rXWJbw/+QOe
MzLYyXnsK/WCguk5Lt3l+2/JYWLYXNDnNFiRTDM5QWlX5iHdnU4ZI7TACOfVW1/O
EgIcaJ5iVWf2G8CEQfSAT9bhnvONWF8D+1Hkoc5kpxofcqZVJXsEBoIq7J+zpWp3
VE7Lr8l8fGDox4aG2RSHB3pjEQkz74W5RbMiU89zRcCDMJI6yxjfWYrKqWQhsBmk
`protect END_PROTECTED
