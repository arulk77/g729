`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCfBgL11i3wSJ6qovWMfBzgFjrakim7hR4q4IGcDwQ+Q
asiZ3TWPk9T6ZdIH6yy3zcMa2tMjFgoXJEPnka2QRzUcyvDHSw3uQDMGdEw3fsqQ
xttm1TknvUl0a/ZRuQXzH9sIHGTkKBzQz4elB3JvElUPIgbmr8BIfiofsCGD4BM7
v2l4rHQ1V6xCAGEMYx4TNw==
`protect END_PROTECTED
