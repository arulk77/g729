`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
ODQFDI5MX3Lw9ebBhbmpy7rtsOTpmTnFf+ls/ywC9VITKTLmjVbowEwVis8JZiCT
pZlQh8R3vHGVL8ey9pFR65XdYjh6UsXyPUxlFglQkbtZfUXek5MVMLO6BzFVK3ww
DiXykdTMHEr84xt3N3Nv41WBF8z8jQ1k3m6HTtp1vtMV28t5vuoYcRQg6M3k8g2O
TS1z1b0c1qVp/p4Cd2pC78C4o2ujMYUi/HflpoASGQ5p8GgQK2ypj6v89GYUghzE
vTUg5ya1hnhDrd8SS+tgnjGvCuEpQCHeIsmRqVdytSbd9BBsCpk/V4cTDBMEQjdF
+ro/38nzDJ/oW4gi2043pV7Yo8c5Xk5HI/clumwKaQRrmRDsvigWI80ccDfh0sU2
723GkchTe72QQvqaFDH50SOyJQUM019coe0CHPGsizjK/pNrdJ3o9qNYwlz8drwP
xIxM8Hm7MuzZYCCCV5HylgRvqQ06AyCo82Ncb5ZxXcANLPuTZba0Sz0+8P5T9Nfi
EupykWMxwEH4DdxZjHXb/T8VsqrIsVqHCHmDXAxnoLV3c1rX5Tu8jnbSYfTY22Wl
37eyWzATVdMVQowHcKbzJwHY2ysZWbxVU3OST9ziOOXFEGkPPuhstCKgo4MH8Nq6
Papo+8SwJzfBnd0xaYtLykmZ0VnP2aVlJgHCfLaRoQfmpVQUOfCFXeEcWGiMbjHM
wtNeFewgkiF8L1ZrWMaszU5JLaZTZH0kprX5GlAQyI99fXn+5Iazc/JVGMO1hN0Q
jKc6RV7UF6nlPDatsoCiJn57A3TwB1z3s+XHrUiUmSyQMQibYr4SCDmBD62avV2F
3I0k18YcVurb4wbn3EALrRN6tMceHE4Ue3CLMRcpT+0=
`protect END_PROTECTED
