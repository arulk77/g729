`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFxujO49HlMGMhcOhbDelWJXwplEyqV+a6M4/Z5ruiai
WFfFevXEIux7FxaB8xmJnWZmb61O8ZuOGbJ165ZzNWkyoZJWOMWitlRutq7hGzsV
wjSyloTuqMA/ZFMbYZFbIYEHbFrtBW3gwfq9ZYp5ze14JbqobBvC7mmYXbuJDzma
ob9HWtIe5A08/a6rn+8tHciPpSyCVhnghLmzhE0oR53hMu4uGRLurX5mCED725wQ
wXFtIzUbaDSbSkh7zo3MsPSaDB22FzLYEB0hYqXaMpOXgzbYo8qkPMKXppFK0GRz
6kOhF6U7GHX5bGhcykY+yNvFkn3vLu+WMZwP0mF2z0ini+NxpLDwvIrMNypSzp0K
z4svbPR7a66N/7rOTLGGRg==
`protect END_PROTECTED
