`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMV5kfhco3qyTuDd5B/lo156MY/UN6wlSVQyZlXsvtAZ
ZYy8I026mdOdiVE7Wo+Al/Y6JViKrv6qLMKE0dFn1ELox6r1KiyvwnOfnQhRBASZ
Lv9D2JaCSEfyXZuPxLQAc9L76jOnmMY4C+hL/LI8TWrvfwyXDQ3Upr3PMI9pyqVO
M/GIdY1dOKHe3m1aEv4laBTUR+pekKCWUUhHXc9BkqBmimwHLFlL4rLS5vMYO5k7
`protect END_PROTECTED
