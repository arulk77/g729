`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAWflE4SQuG9hYa/WdOX9lgC3hXd2lNPxhj0dFZqbO5Tq
mDZeuQHDOUmE3+gmovJnLYwIzI1ZyxNRA3/cWO2/8H2oe48QqukATjxxh9muEryd
5ydV/HjO9eQcjhy+3SzA6ZpImeEdzM1tYibk1vl6Td7O7tGGkhxYyX5yHMO8m+bE
Dy6A+nJ2YXg4a8/O0TclAexVT2HQWdrSnkO1vWyC7rdNCOIdwbwQD7QSewGVryhO
YJAxlIXI4vTXXAMNpbvvM9rInoQd3kwnMNj+SBm3AziitfumUdLP6lwsyxmSjctx
7hi31D2uXPLA/zfLp9eylNEKkWYYK81l6uwlxT6hnQPTRitWcTdBzcjQzkJZpX9T
Mg9oOPu8FC3kdeMKq3Ivzwr4bD9z9xyAmgxu9gqnzq/guV6xiC7S08nzF5qGB7dC
J961eSBeSxu+GCbdEizNjqO0FhMQGHeSQ26zBIv62SGs/hqpqhTBrtrOU0FJtHN3
dr87BvI1gS6CaI5qtnjuzwtvRNdpz0+iKQcYv1+WBIMB7uiLjJKwRhTfD3KLfCNa
B1jagHvyewfGBG/SbXYBuVKp7ygeTbjR7OG9KEsrl75R4xptLzvgrViDIKn78a4C
w0WgrlSDpIcDon20x3NsKtzDumH0xvGQGFbM/ZDr7FxhK48zoCcv7fVD+kDav4J8
auJLTG8DUONXagzJitqSJGNXnl5h5fFN2U32zogmPz2WPSDx00mY7GZZPucaunBK
gn/mjF9+A2Ff9uTAVXDHq5VsdGXIWfPzqD/X8MqY2kIrLaGvPoWnndI7bMjj9X4z
OayB9HT9KAtAYW/7CBd5RNCzAC5OFgmD9q3STKfRlzQyPWjVlwOtDZyam2A6VV+1
D4se4pKCjoyIWT1cjoyKuxEl/ax8LX6hsD/te5ZTMaHju4ygs6lvbJpisRzt0sIg
8S0RF8xk6kfi0KDOaSvP8V0YDeRey8TO0Mx9z2NsYM5/8mEj7XuTlSK+PZQfz8Hz
Mt4HppZdS/LvDbq0wunHPK9dkwuhZDlHONYrsmlSvuBSVDQu2dOsuw8/mKgD2JD1
XOKlkJKZ10AExSr+pnetumjIOQA7HPCpRDLSvgpStffd76p+1lpYRyNY2ehyYC4+
BhXnhWhb1HWL2XVXUN8AV3n2EAPAkjoPuNcXnEWGeWhoMPUDc+NNXsy6n4RPF/Wt
n6MCoPW24Kc0X3giKCg+oeAUbFjIoFI1k21GvpeEwenogqDbLQs7cq9EtzKuqACX
/+wLtjanIsC7R0kAcp3xay8J9QDaGxUWls/go+RyTjjm0z6XxreYvG2M/7duBrJj
Z48hVxjAGql6PkO1s3VVCr5grntRmEHZ6sy7+2dEn/CILwEyOA4vQ6xT0v/QRImQ
jexJ+w4I3z1VcAu75LJnEiGX4+5S/BsqHlOBw9LsE7ycdrUT+5w8ts4QG+P2lXoS
1b0p9QogoHg1doTSJzjdqIXndMQs+5fm8bPPPETrJ12SdFZj9FGT2215+nIfhiVR
Y6CFXhKpSM4L7j8jjEnpaTJ5eK7UKkWRAnuh+zY/doTkbIdFPflKh/NYn2oiSOkF
oiklKxpoXvez6KSbCiGdfKzUaSiF20x91bjBWMgazypItuwQgSn1Nmy1lgr/uJ9Q
ANkmBiNzrCKX6bCjabm2n+cq6oRs+VO5cu1RVvTkGta6JgoXkUF67oDfV+XZCtG+
nsM6FZANWwDCVcOGchkDP2VRmLsaAJ5k6T1IOuux+sSzoewGY+8b5mF4ixyMlNZC
8w4n5pgvvAW8OzQvfCUqWyV0AkPbX9ZRwMiwMg8d/yhschdFZofNxAY6QYewTyKx
kziDvc3p5VOKYx7lEbQQM7zn1Q2QFxouESOWXOIQb808ZvWl3ALdwr8X+Kk9GeOs
qHoV8xgNnUjz9tyMxxznhRbzYIK+NgO1Anb/LD+cSLIKIVlhW179ELCqb12NYARy
zCxrdmCYjhMF8Z5F00X74OcPZIv7/9DUdi2r7rUqw7H+e8ZvEK8NE6gKfeVUXEnP
WuPlq2HgsGjvoISpLV8t0gOGYK/U1OIkYhUWqSgVg0gwWqwilS8jOgBna/LIbLxw
riQwB8FZT7H5D8uKyzciS7jTA5jRqNCWGhwT1fFKZExgtUlfy7Hl/z+itEPoJ2V/
uJbqkM+STCbZsngnBGoEAiamibR2EPB5t15qEssgPsAIntn53sUwCYQyCSd5E/wL
JwJBfHbYeXPSd+Q6EjVgsHJwZGtZ5CkVk6qEtP45Ix1GRKDadup3z9q7bwgTYOty
rDJlXWfLWuy03qYUir+JjdywuNQLHJ9ZgY3ol8VXk7lkd4hMYvmivg+29pC4yn5T
R9pW1KWXtLKqncm10zt82S+IboTiNjeMDaBRBZseI06aZAfGSdswHZZLqWbv49Bs
1YPHK7sf7cI0EcU58U8+27h0ymEquZv1FfEyHqm+rZnyDXw/y+48c9hKv0/+Ei/Z
FQ+NSf0uV+WqFA5FXkLYE4SC5avqFPrzZX8UlxIEuDFhfZNR9RiICburA73wuxFf
I7yz91ES9QyJD07AyLegmqVJDWvq88+eCkG1bJjcoAV0PUK465V++vXl+stCxvsC
/5ooEpQKuagK+5SgY9kYi3Pr1ntenCEfeOAEzOE9rE7QytXA7GfeMJ8D3amz8ESg
JkHLBc40mdsNpx/4nPIicvHi12lFm/tkemMtTbgzIPXwsXuBivj69a/Al01ZoZK4
A9G+H95vB7HtQcuIgiVUXEMRj6F2iEWnKpwrS0CYZ9tL3G6OxDmaux4fKf1DOIzw
mMH4eG3kPjFKj1OtMRL7Z1hv0advdnYtx/WnqeMtJpjF5xCkboJPPSLzuCDwerOr
Qno+H1d4nIfZxp3Bd2ZsgiEe4G4ensxamntC8ypKewGoNRPDGL7qug7fAwSiG3ti
70bTRt4VIbRSIfeVWlMvjk9wWzfHWB7cPg8209HTxXZolsyrPwbljQ/EEaIOfpyy
dxXUgrYvG6l0asf9tvc6/efb8YJfB9F+t3au4ZrzKOLBmfVOaJ3pnzZVvGuY3qHi
0a80JMUILhf6CSFirFK/y6j9HaaMB4RXP/3axeHCWAHR/ER/T3VUuOfOkKqSra5V
mtIbSit+QmmlV2AmZFD3wWRRc5rYT7BNiFsELb/0ulTVQskkuRz3I3VaX/dPmmBF
ek+HsoQSQhBeK5cpmRFhrAf0jLDf/LA85+rRtL8zILCHCWT8f65JntcgnoBEYxRY
ExDEGkDeLENS9LU36XHN6qOwM0H/CoMBGpDmm55LrrSCD7G0OcIYO6uy76iDQgCM
IVoV1UP6nvbUci6WabBRk5PDk3NmWqiUoG0K8t7f+imRUFNyC+iXWlsBNiOePTFL
d07s7W2x0P+O9LJNWUMUpozHe9XlbV45NKHVj9Hz1sxy2YQCbN3pTz4oEhe2JB2p
I9+tYu3+truBUipFYciT5WGIVOrvLc8yrntQ9BgkSqIWO/UZd39g5PQm86821CNc
WPDvWsOSxPw19+jT81Uh81KHGgyEYa9fcPUyLPFjZVVrq8iBF/oUK4fhZ2ZJp9Jv
Rz72g7afbOMtZTmNtiEVHWBtKkIWLYxzqvDND7D+56S0uUOsUJ5Jh+3ieBa4yD6p
q0Rh9X/DPMz2Xf8riml9mvVENVl7/D7Uhj2SQBUdL6LadIT1vqhCyKDsOUDz7WZk
0UBKqMxL50/xqyGtNzCt6PeU9irqs8wx7DJxZh+laMSjfHJJOaIXrDAl6X6vbk7I
sE45kJuRfW2xRuUPa2VPrksz9k8tTxSVQrlAjJAaukkRkRM8dkyhyjwtRPn+rVW0
OOnyObp385LlfJZ6pqHFh7e++3XdtqO1PzzpBRCEO1ffVGHl+FaXoElL8eDd4R+t
GRQ+005mpWDXombt3SmgWRIE3//ayjdsp4y/jT9QKHTqU4roVjSI9vbMf/xTjNRn
KsID9ZJlIyAW7VW4cIUnkZxryEPOWq1Ryt5BmwuZch9fAva3XcGVO1lerNwPrNYq
`protect END_PROTECTED
