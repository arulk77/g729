`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCkXZg+EKhF3TtjLIAdCHqqBauezJGej5ElV65evL8g3
KOwvhI6fjwDG/BKW7bVl+i5VurVSa7ZMCYcjyYNHs4bpOof5Gp9HwbmQLILnkRq/
ndMbvngqxFMNfh/c9Y4+eGadazuk6p0hREf/t4jx6wz5HFG83A8qCsKIZjGSBB9c
UbM1IC/YOKx/q83Uj/2n3/oiR1bGdmHJ/Jx3aO+DBqGdRwUQf34uJXgIzkeRPTVR
fOBEoXWq75DeDGFvV51g2J+Svk+4XaiVEpDQ411gd435GnPNdNl040j2yLjhg3Tk
GPFuasfX5CunoIIx2pBUR6HOPjgvclN02Mt3jiRUKf5M+RvpeV/jiB3CGuHPj2M+
iLLvINg20DRW2IvuNyGXNLD6eu9vEUc0MFml4B11fD3DEBaUGLwJR64ez/D/s9p9
Hz6ogkyGQshcId2pNpMIfA==
`protect END_PROTECTED
