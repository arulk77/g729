`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41lne059/APcaJ6cHTlT4Tr0B37W9+qeINyGx/I4kQ0s
pAMK2m0UCNHRdzI/qfHni07RzY4UPoFdvTJfvghKkX2s18UpIQ0b1H3jVLNubZdS
M0FjjBaNndNIR8OSd3ZpBh/kzwqSENT1u154hBGlZAKlQK7gYWBNyQe5JT7xm48N
POM/TkfSCLSjX5g8/ox8buEgHiH7GeGbGdjwX4kwsqogMb72RxZHE4wUGoNe1zt8
y3IaPh6LTFcxtkdNzAO3gfKXxM/oBLB4mAhp5BQd0nYW+N/7C547jvYChusLVG8H
JgzufWg77m6oilf0VfRKRA==
`protect END_PROTECTED
