`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
HOoR1WAPp9vSjhFu8SDgjzRc7XEFPUCy5Uaf7f0Gy6NiyVCcg9G69DSIJvYNEz0L
WEnmiL7KGtBMQ0BNp11nRBcB4lg5+ixHBmeqIzpQ3vYCVV4YkGsml1ECY0+4bdMW
yk25FC3SIlwJIakSDV+aAYWCV4H3hiZ/UrN51YQi6p9ywDUG5KwG2RP+tu0hKBov
xGd7M28I/UdjzrRhpy2OxnK0iMTDVXkXoT1TrPpAjnsbFXLPAafqZi5GtxPqcgJ8
9biBzJr5hGnHeDnYK+tGyaLwm7iE9qy0ONF+RkGvTtA=
`protect END_PROTECTED
