`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveC9rro1Nu0uGVCd8p5+VrUprHTbUrVb8CgA+Ry36esJs
vqTLKdtuCkaU94IcBRSj2ifuKQ8CaU/2grTkVDc/N/s/ssFUdPpiJp1a8McuKsWN
V564TOh0WndROsAZgoUAvbNc7SrdN/mZ88LN/AB7wIwWfwpI6e+ba+0k5bNj7KV5
9/JwlH6w+3T23APVpCq9lGgj1aOdFGoyC36Xlvj36m1LwmT1e3rVlUwWeNQGmuRP
gaI7ZUxGZT1vjQMCFKF1MA==
`protect END_PROTECTED
