`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
jO+xGX/Bqk0brZM4ztto2tfx3UiQ2boQ1xWY2vEsIk//Z7jXP69/rcSJo3H9PlIz
H/gbjv2pi02cfzb1OzN4Lf9FGY+AaquJV0SuoJpV2TV3dzx67iN0y+vPCa8oOyth
EMgozFZhZ7xZOq0Tomlm4Gcsqy37ghc4f/Z6/dkXXJeFM4TlDyW6rUyMG6xXxQsS
3oa0gaOnHJ/33BKLNMKTqd/r8O1NL/Czf0eWdQLSMlpyM8lnKCc2Enw0gaHMVLHx
yuyizVqdaZi1IQqBlhiF2LzxLA/ZcTMtl3J011v1SWVOk43ALPUmHpdBkAEOatyb
GZJthW/pvE7UfTyd8hdLJSweTrYAoEN+DmFslCSj/fs=
`protect END_PROTECTED
