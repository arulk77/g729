`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
N4o89aDHyHCeZ816w8WVHaCiQaULNB1Ab9yNEK8LzQdiCrtunBZUYJO1qvBMub44
9X3ic0hyYA2x/Km8Fe5snjQSfdICw3pKItP7eZY6ciGZTHBpTNwzRbSEh5QhjgC8
cdk3FFQ7XcSggl3JM2EBMFSBVT7R7J6bllZM8LsE7+QFXbJXK0JQt2/dmsf7Gwh6
/FUNMxLg1oHgFmlWJZXrEc4fVyPXrwKBDZC3Hc2bmXV59MQF100xIZk+eYKDE6dG
OOP8pDbLikyFgCNll87AgqLb6X6rzgcXE165C4UQwbuearspMOzXRZ5wf2/zggOk
+CuVx3wTLyIEpXz2TxOMlHHOWl8q1Y1yIspnuYRJTmfbtFzLMGnBm0x3tysBPOaJ
4ts1nGE82JyuSXPOtvzteXEl83DPgMAfAucGbehMFXaxgVudxL3kNNah6ctV6wIo
FtX+6sZrhetnIT6xP2ArtFHR+GuiXmyAUzCdUfXJAYQtBtnkOnk2RQgr1vjea4uD
rJMrWG+tTQSpxyXOMlUMI4DL5Cbg0Ch/Wup1jojdn8wlI6WS7PF4XUDxlbCcW3LF
jOTu4ZeNz/q484gXnaWTGhzdXw/YULiAvWz7iZorj3OZfVqp9OrI/ieCSXpDin8t
4NuOfVykiPHfJkT4Pi3Jfw==
`protect END_PROTECTED
