`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJJyYTyM+ISeP7shjD7wVQTvs/VqxFDiDku8V3Fjmx+i
LbzwxtFv995aJ8Pvjn91WNxigFI2x08+VI2qyxuhu+tLZ+a1tdoq3wYx2bhA7xgu
Z3jZ7sG/lT70b4kqysOdtqi/GvL2hBxnEnbP8dg6hoStwCPnFLn3jIiQ467b1VMR
8neB6K8nEhmZpejHwO3U5MoznV/jQ9Kz/gtYKERdTRDFyNif4nlEOsPww11fuvzI
ZD6xe5uXuXkHehjEPToLYeGudlUu4a1tkFu7BQfHD3erRPg9SWdq+SOuCwjCxk8a
wtW5+oLzXAfwefrOlzVmtGT4dBzCX+zBsh4aIJZnuPANr0lnDCGCo5buTBVhkHCB
ZwzRWuB5bRww3XeW40nI+A==
`protect END_PROTECTED
