`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/Qeo848Jv5/TO6HO1Pk40lHPIhDpsJsh50HMoeuFVJP
57mdrXEsCnqIRT2q/SJaBP3J0UoeGcGLZQE5QkhOg5QOZlx68VhbBD6fimjtxkN/
RbjToHEfGJiBhYauhy3AP6ji3rrFtcbRl3pct2zrN9h0F0EhSEpeBrCxew/jU9mW
1Q0qmctWWxfe2UbijiGvKwSYMvWI2RrfS0QanU9jtNfenAdm+Jlbh/1BDTDWi6TF
ncbkfngSAQWGVyzQ2MfoX038EYZPGnIRDB0wK7HUDx4/2H/dm3aPhhahxIXxYBPW
QcQrb+eiqwBH2S0UMUhYCw==
`protect END_PROTECTED
