`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
g25ong82OivH/FgIaQKtY8K3o7GFfzI8CQ25PqZ3grM4gPjpkpjDYbCdHIbwO5s+
E9Vf6mWtiCxtY/1GucE0VKuMoviuEZSf4TLRol7JhCqBYvfEjbL6suXPqKNXVH+n
7hATHWtIpwVtfjxWLLCUU0GlwImzkbjXUPjNP2bavlPotpG+OscetiR3eqrrYD95
3h2cUoWtVU1g2EICcIfXOML/Ez60889iKq/05TItCP1WoooKV0oYEHImV7IaYZLs
tOHAnJBmFbEwxQw9lHyrZvRazsxE8xMPlG/mTPvwbAt7r/3/ZWE9vFqXzSzUUovd
`protect END_PROTECTED
