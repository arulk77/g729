`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
aUbrwkhWVFkNno0Uue73C2Q2NnXolywGwbyF1TBvgP+I9D1I+MmQZKhpl0gFWJsI
F10rjxesrSsL4Ety7kDFORKNI4GGVtQak5lkuaDM5nkAvVFzN21HTkkhChZB/R+E
kcRi3cR8Z6PswneU5KjvzLng9mP2GPsTVuC5AMuW5w+enC2R2bzkMrOanYWDmOB/
y+TBSSNSTiF5ex/q0xJJ8fe3Rvkd/qjdYLsu0ke55Tm6OoBSstNeXx2Q9cMF4diY
/94ChyleHl4PdHRMcXMnK8wDykbXoxLHDnAU5GSMtyhRti1t4vRnY1KUrWNonBVU
gaLVEhYGdg+DHEXVtiL/WKWE7GhPzneJW2ddq86xuCWEti+dBJlv7oD23+EO5OBq
lq0fn1xuBm57c4nmCYsdPfbPU1YRjAocf3WqReHCeO6l89Dk6pHOtQRVBZXfzquQ
qB6ruHAwTyMI6eDlBSWa5KFdRLi7+DawYDJUqNwFah0K4NkQg+q71UvQcy/N5XyL
nIE+2PkHmIvY+gltPdfRqOI/ZQkzVxS30ryH3TL5+A6didb/8Lef6I/e8Nasc/4j
rr37lv2yaw+uTkcfK5kvdJFPsuhO4xNtwfJ2/GndYNA=
`protect END_PROTECTED
