`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
8KWuuTL/uH7c7pLR877NsJQwCP2eNqGJd8LT3ohHBJdLUQcsdpKrsoxdwJbe4RkX
VRKZAjroUD+oHiFHbs3SytOx6gmZKSdNkUP6wCJXA514yc2c8UkcV2AHUQR2OdbS
heXxVdn+frC447koxGJuV+4fisFMQr94XHtCxd5cxt2AxlgNeFYISGyMoqO+6ZnS
D0ebnam1DlQXOOj4Nu/IguvzI3XaWeZ8cW+gRrylMUaeRmU0Po0WB5inl8nGFcvo
VsVaOkqiffZZaSi+Rr6KZ3yXYceG+SS3tIO+HO8dA1/LSQaDgicIWeacaEuLM6bB
KxqWRxT7SUZvPJAgBwzMyvfqM182EBbrvDcZUq1urYROrj70XrjWM7dibM7quBBS
i/bSHUDBAzsIvlmdlWlRX6L3/NuZ2GnWd8bDN2qncrU=
`protect END_PROTECTED
