`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveMuMESNChn9UTJRhPh+n6aEUnHs/NKmrk3HXlgUelP0R
qwaQGfzLfZzm1FVP2aYcySCT0Rko2q2zBCSauGjq/oSFElyXsw1EfifgeUuBPOcU
R2bcCKm+KqL00fziz3XJAa63LILjWoKEpmughdLUGl6lWibY+v/uH0qUj0EZM+sZ
AdeaJ9xMwFYg5JHp8Nyf2hoV1Z6A9oNi5hMv4krQse/aWmopBoDGYW5Ir6spAmYq
bGYK0/0h+CPzjlbhw56plbD3mreJyIrqezaHjfXOrRQ7YvEo6hWuqnjoRtVkM3W+
ARYOyvByAdH2tsJDA9sANiTRwgqKjkCzaVl+IkfbDrsMpewfHFOqmR4KXUGsdzbx
`protect END_PROTECTED
