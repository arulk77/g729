`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40MMLA1/l+u5Q+vn4owsHIbJzpA340yEEhs8HlyyK0Us
1UcpBZ13EC1mau3jHfOhpdB501UbRIn/9SJGd1YVaTBjXImJZdn82bdj8GeTVK1k
CGARlW8JB2xFizRWjQtysCBD9M1c/zX+tpyS7UXAHpPKjLZruLKYXjQCfqUqWpv2
DhTqV6mfrvw/wru50xTJoRgDTK7xb5rW4E6UV3CqBaEDPjUnRY/Q/G3iGAgOkwY3
6OWistWijgaVe9o04ONwRIxyX49x3+FO1WFZn4/cv4275nnqYB8Ed1GdDTg8yjyh
Wp5s0qlTjOlumKN0wqCs+g==
`protect END_PROTECTED
