`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAUGlfT8ZI1BCgJu7YwRuP84wmn/LjBDp5wHCoyY9x7nI
512otcOLt2bXEous+N7cYZO6cI6X2aMPbhILSDl9NuLJv0K39PEMNfpBQQErnKJp
0FHOvXZU5sjAStZj+3yPgyy1bVEV9Kb/xWAdrRTBNxuRdjLxXnwaKeUt3qzXDxzr
TJ3OikZzguJnf69ZFAxMyDl665DgVhHtppcqwMknyAkeVOmXyK0fhPq5Xm0j7prt
+ZIfFRvuL1Nfiez6ejXypPJXo6HdvPwJzNHku8jWGGDr14akZNHYwtnsBCl5lSPq
h7X2AJqMxaRFcniltXZjxWBq21rU/PJh+qOtXVoFf6/hCjDu61FvDfPCJT16mtlM
od3GWmBaN2rRtdTzyo1uiM+C4XUTVqcHFMTi9z/jueDWW51XoJP3kpx+jkVzt0DE
P5MvAsr3iQ1BlPOMOhFtHtZMAZk1rYqkZG6EAE17nCZ0po1h/Q48Ibx/Y7KkTQ3A
DErND8P+zpb/TVNQLKD2WA3hJfIX1nWyjuhmKn9+xCVOnqyTXwjnkzIWUqTjpgFc
xw87IV3pPFdQQM9o2LlQNq/yNJcYCq55+bhXpkDVBBZVyaaBh8tPuNBbxBJN98Qe
YI39UgFHP6Enkt5Bt9v8iL7aGAmj8butRuts0DUhKpZV91O3As6Ecv2BcGy5WVgG
NscWB6k9gBF+qZTsGcb6yhkABDpewKvPMNpFR/ebpj60wwxhPeKfZUhQZEcb5XBd
bXqQu9Vyqt+2KWYyIt7nrWxHvhmwiqg4zW10H8LjgivqXi0PV+pvOxxJp2DZKcYs
pvx0aTjSm9TN5+yJZDDlSwkAwEvugMgMmo+jeG8vSuO6PGKzvLaT6dMl8myOxxjX
grdKMfJQCoJ1+0tsdWmM/KJxag/q/eDOgODZwEcEUrZxdUDi7hClnY9bG+p0tMLx
WksKVqRHq1YtnjYv4MGjNXg9uy0mTJwyy/iCWEkoOlbC/8LjJIvWGJe2ar5Uh7F8
VPjpuOESaIqKXJPQHzVreCI+GNF8Y8qXHftimFD4BM9JF8p5uTs+TfP3Y2zzC9AY
fZW/BwfulSq3s74llX2TZTnmBC6efi9okYY5z5mxBB4/XjaXEa/OnkzMEp5QtJnl
0T1QTmMKrbjpdmnLjgdmjEitDki22c/TP0Zmx7O9B/ef6bWyPzZPscAALlUAXf1s
ojXJUFfoDG/ggcgTwiPrMezufcyYeM1b+mYgXi4Fq5ANQIXN87eg8DWNLjCEOGDg
yfVt3R+rcDIoqQU+y60EKK+ER885DWOe9wCTKtRCzIs+2cMLe5XqQcRxJmnoaGn9
D/scSjFT1U0yc5pbz81hs7a739rCHHU778XExillhygQRWUZEaqyq01JNTdrQx6v
Hv3gvIeTVt7SZo9sESzwjzT5iBWye58HwpttwfGEBKyGrXjNKPFwHbr7SmhH9j+g
H/wcbWSqP8U2gRb6cMXnYcrx9RWVwugVYh9Vy7RTzH+V03Hp0HrmXI2QdSrItmdF
nF/3qCb/iD8B4gFxzH6UbSCic5uX7+Hp34dxv2ndUTUbYP8KhYK31z91Im6pzAa/
hZnEWqtJZzv5LqNmh4DhTCqnRpadxhgn0adFZYJ3vfvgEvwFbVa4qjlmJlXFb051
q2HSbu0MKmMo3y6+LrZjyUwVAmiWNrenhUY4LqVShTTh5ZiEg2xf1sNBUoxcBX9a
s7eK0C4b1mpFF2jr/GeLKpaY/6jTVvmbQoUuu/y9KL/+V1iocLHcK8ogjDLAYWol
EDgvVDv/IPRMBqNuvNhtJm/zh7EW8Pv94eBxCW7x/Su+IPzO+EkR36axCpc2+leQ
dUfZxjYQMsSu4msH0xIiQ8RKfHPlN1v1cIY9n4IwxasffAlOqVCxT7aSs99PZ4V3
bx4NP32Ih66Ua2Ih5JWr4y2sPMQ4sR6t+EqWEWPWXWBYfIwnJPxnkVilVnimIUSS
hciItF+PYwnPklJukGG7oR3/eEBuua4bm+Ewx1sCqu8M4bvcYpxSfc62AI/9N1Dy
b10rpUlB/16h4FZ7IL6XP4ZqTqYQdw3zDWswsjrGXNXGiG4Z6pe9VlkBpbAwsSmt
J/6YBYt6uKOurh818ucF5OzFv91fnzv0jwHzDnNvjmRz1PvcBSpYj0ESeJtBAAF4
E3kwDYRPPH+OUojzPOQdbcgUP5ce2HbrsE3UMUry1JcOLHfKtDD2wjM/Y5JTHluY
ZMWf1q7hT/vrAV1EqhsWN8kODtgXUK4/0JisBwDVytNB5YeDvTwE8q5FEEmlYA03
w963cNd8J8Px84/dBiIJ2WFRU3n/T6oDIlkMhSgscrnEPWcqeSLTX/rzAWUvenwf
JUb53EWUNg/fT4tZ2RUvHIXlZ8hSOd5otPaHqn5OFjS59YQ9efL3rIViJ68eL0FB
U4Qq9KXjIyGL7XTxEnLAMMSyoKEne2HIKlK+duu2pOeBZGVYFwwLv/MVJRDfexeW
6iGZOIvvoSi45L1+60hofY6glVTmVVyNfzLjd8Z6i1IcibQJFuiWnAlziyN2pXBK
KCAGV0v2TAATDDX/WpzYS8HyIEgvwckQEBqw24GPHpLrxSoy+Fbx3p3iTSp//Q0D
TMXoZiGa7XYA6YTNdM1mANHhO5U8wOgSoqLwzXFst8+Z+M7Y6Ox36UGuECNCbyrk
fTLnAOQQapibwK3uX4tLT8uYKIgr2aGpl2Tb12fzCv1LGyzQg6Oo8YgayVUrfdw7
sxc/EK7YNeF1GOGlOL9rEj0TSq0t71KOQY2FM0cVbd6My0SSECyz7iGNZkRC5Jsi
aTX3HwrX0u8qduaNv0aiY5pCxCDehz5Il3FHd3OLhJtnA5xFRFvyzt35My79bRf8
uv2UbwJZ6mySZ2Ch0nLwDNEeSUmdebmbpKfANdKgFU0=
`protect END_PROTECTED
