`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFBrXu64XIv0DPIOendBWcjRJKSeq8dzy+WOILApBfbJ
uuSh0b3QstQTskW9nfOfI3xODuYZCtveqHRPDGA76YQ3QYCaqAaMyFsteSOfVOSg
D2gHcrOVQa952JWnvJqiO/JBg0qyjEgUaFe8Nr+go8KQvUedN1iGveJXr/Jmsn4l
KBiua+JJWod/ReHI/CBa7DRgQYFOnI4IJH6jgd1FDsxCrrXX3HO4ECkDoSHZqsXU
YRhSkO5TQ+gF1Nl3ZDlH+vwIJObDKU4cKGgoDYW3sR80FjLO6zp6mwId/Xd9J+l1
pjHXTwaMPGVY9m4M/3MbkA==
`protect END_PROTECTED
