`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
C+caHu04tCIU1aEDQ9u2ifFO73UK5PBwaVN1o6vBsfeYYhTMRgICq5kCji6ALxjE
0oGfIo07IrtA93HcjeFG44Tb5YhW33tD9n4ce/V9JKd/m9wHw2fhGbNaoe/IsxUZ
pqXwLqczJZbToIwsSkAb2ZTVReI/x/HKtStAOK7vlFiRPiopxk4odgf6qlmRrMDy
RGpmsm9kTbNjEXjHz9kca9JXCSxNEQZz0bsE9Xf9Cz1HXduQSMSraYLVCp2bJSZU
O4T9n2QamcLrDF0ox2I/9gnAh2wZT3mEJ9NKHGvFBcFELq03/xxY7F0SjQ+eXsHc
`protect END_PROTECTED
