`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
76sFkWaWtW2g4TUTKwVVqpo7xQG/iefyPbhcIGbO6qgyY/DKcmt+pJGKU67dSbA0
6w1x0dDKJLmYKbFWNVFeTGtGkwnrlGu+XK0yk1kOrWf4rtCYkR+gc9RXGkJMGwqa
1Au6cY/mQqj53rTL3AkWXtkyiASOADbrjkbWjosHAAG6qtMFnoOng9tfTEqsjVEb
ovty1aL55j3ZsRzM9ow3I0p0jN+drhH8bf2zgG7Ryu/JQ+Hq94hSG9naqkKwk2ZN
fbJeJLyHpMd5X88seeDLbuVMZkTCeHlbRa1S9kshw2ur5otUxjXeD3ED5VVVuoL9
slhy8WjgacXUA+ugJ0oJdGliCKiPOP03PjxK4yZOsEPEeWwdmsesMuUIe+4R6NAr
OM8rbWljMBAfxsZIxoB9JMEv9k9Xn6CiTD9hcSuwsek=
`protect END_PROTECTED
