`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveCbjbNLcw3t9Z2suMq1B9zUtYtY/Ei/Aqz8TTX0yQgAE
E2zgsFr2XvNwM/OgUn1rIU5bCZnzmWiERQU9DJ9BSeNCF3kr0opXWk9a+Sk2UJp1
hrO4vXa+Wgq/hN1x/11q+SDWEPL2c8hDJ7pD5hdElsGvnexpYXIBGVtdV0oXb03z
pJ9YtPJ7H2Vk/APhn+FEcRYO46Isr6x/KblUWzppvPw6BWB+kX9mItayR1boYkS1
M59IJ4gyxRbdg686eoxb7sNfbQxDDHZ/dENOJ07X4aA4XZrB8IYk5uZAGijG6wg1
7mqQoRrOW9+2jMz7q1cBp1uebOr9a9hV7BndVv8QsBZ8RoSdgDoUarYj1/vtcSqI
So4s5tVIi+wtmJkNE+dNbhjBDN5EAmC3PgWV1R9VThJoJCu3yrCpQQJLOTRIcq5o
d8wFV7GN4t0A4d0Lq1E00EJcKTRX/T8RMpgeI6ehwcYRn9OpRiyW5IC0znvT7p+0
Ev7Ob1k1U8lp2kyMhOQFf5k7nAwAfKGJO/o4wOmDNhCfU0HSDdQ7xnO5cZYLaQBi
us2zBNEFfim7BJ0BAlWdrU3UivnHJ1jlaVJe3utpaitUFmt85tC2FUmdOIBGMMHa
`protect END_PROTECTED
