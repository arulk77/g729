`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
tYiU27naN5TFgRHB3HLmj5GDyLLf3qGN/N2OdWb5JcMiycBin1GOK66nWIOjr4T3
FNuDFLG7sThavvHtWjgWM4954zIVLVNMdMgCH9vWL3YEnGO11R2Nddtd977Et6K7
o6FFd+aS3nzQojmIEd2NLG7tiHRVFl1hp7QZLjL6OUYy1cLZgnNruHTjTcQmAZeW
V1kvUJ7bvCM7KeB+NBrhBypb+kQ9+w1KmsxUZPXahSNs5BlGyUaSYIAhTFDbG97L
Sm6+MahyeA3uqTNBXDGxloYY+XCK8mL8mW2lqFf3xaXWF7oJ7dxvW3SCKmnU/ALi
UvWkEZnLfDi3Go0xNkVYkEeg2ywh/TfHPAv4pTrfMkFY09g6CN81Zui25M08T+Tk
lPMIlqNQkm/l9hOIR7sbJfsCWChoKRnHAjoLfbvJapIJsySDjkikk5o/76TQx+UL
0ptYQNdq69SexK2A4cvOmWfllI8VSz/eI6kKLXVpQzkyfr0QRwLUf7t1eJfgVFzH
8xz7UDjA96VA94WQtf/C4idIx2/40lRVqOtzt0V93ddZG2OBQ9e1z5+tLsVvPm1K
aiUqQ2Pa7W08kLeFGZFnsBqwTGXnWPrURPf/b+fT2hLYm6uXRqDOtK0G8XrydTYk
4PedD+adcmbM2/llwCerLvB/l7DKnqyCcK7a3EFZAsLaxNfZBsVSfPSBGI6Jln2+
ESAQpQCOdviRfk8qxxXCKVp1SHPnZuMAlplPmQKy0ldxjVHUcBBeHeqE5iiD/j9P
T0KssVDfz0HJUQLowMTMK1CCopoW8xacGoTZfGeDbQR9VPaY/CZhls6LmU6hsEsl
PjMzalSVaDvlcoxPP2kdajI5sFAKp3XHRbtngGCZoLyzQ+amMWiAMS52yjzpyehg
fvlIXS1GJreurQv7b68e3g==
`protect END_PROTECTED
