`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu48KIsh7C+7myajh/mYR3VYMPDtHpce+ZorZgut+rTRKs
ev/CFfG0IoDdBWCtH+Myn7Hi3NxK2GQD1Ud+tcjjPTrfLkGln/MmQeVrffZCo0mO
K548afh96ThfpgKhzCx0dMJZMsRIzWaOPqVjqX3PESh9nL/hUjh/7RJ1Owmn+6Pr
KXFZN2SCWFImfHyHCww2epET4zNb1XSH0mFB5GO99SgrS9LYB59JXZt6VWHeCDrc
Uj8tYU4C6sYzzZufEhzDBx5HYbHIrBtUJ2Qpz05E62sH0IdEkh6SiJBNjC06e+U8
5oIG1stNzCd3VPpmG7kGyLKUtErR4Q6ZTDPOsIKdE6MRMci5rOP3gz7fH6EQJqut
atKTP820Q+IJmk/jnNxB7TW97vpQRDd9+4RmEYN1toK6IXff6zRwKVc2ztwoDiNS
k/ZN8kHLDbZ1gxNzVuS2/g==
`protect END_PROTECTED
