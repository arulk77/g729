`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
VN3cZiJB9f6xREOOK65F2s4FIrw6F3q8/US4L6brJc0t4uf86aSJibz6AlUi2HlP
hkuDkepSDSCcf8eLky8wY5ZfYDeRsnOKM/625/L20D6+Ae6jmeqJRGEa3ZGxf9yL
EoDHagQwBlQRSpwVylbw25DTp5Awu04qWTED2a/Ka+59mjfvqx3Labjlf3QWOLt5
btD+ZBDQXJ6+5iYl7k2hRsIS9jgTFiFVq8p4/C8FXx+dchy38V2WLuxtpF+4U67J
okSolYF2JZQ5XVSCRBfMj1YCsOcSRGRXN9iNIQ8HfMy0QJhDd5hPadnxdybwuuSj
y1zNiCIfKvrcWDWWIHq9xg==
`protect END_PROTECTED
