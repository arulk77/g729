`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
pyw/x5B8DHOlnc/GsKQL82zH7Hk3vfwnk0F6KZswqpdKVNzL6ugw9CKO47YzEIa1
1UVXpHBOOhp7GtQmxejwdg9w8wUEiRGRdqgfw+PsEoQ+TfVxKWSZjaQjLqWpuT8g
+bNt7GFwPO54yqoUrE5fsPu2mtjnxDANjphtQ8k5bPfXWZloTkdPwx5USsC6uYK0
6z7IZd7tz6iU8oZqjmX5lqq5rwgnnvNjLR2XHdkQm3WO6uweGoEB/vPr9AwxZ7Ty
5gtQ0rQXnb/a1eHxcwbOyc/astW7AIZCSF1ABYAL8RM6/iEyq12xwgJ2sevWZlhD
bdQFL/lDyA4JT96sfyf6UFHI6mnCx0lN7Hti5YOI+FnU0hDbC5R9efCWHuI7guPP
JAENtY28FGGqEhAGityWWB92DrPoSekg+6+14kPghic61S1retjsy2TejJFWbKH4
EuRPxJqAt2xMGy+oKA6HtKDTP6bdg0pbN3D+j/dbrqS1k6Qvyd+trajNqrwa3zYr
EM3RJJS9R0+/fvv63h0+rGdEF/IXGVz/J55NQQia6W3ErnO9sACZyYbprsszuU6Z
phDgStyvEN4uUkAnXeEcJuustqiWv0Y8kfSyb5ahCeeLeZQFSy88eon7C6vhnRun
4Hs9/V0edMCedyneF6K7vgPyRfgQAuucRuo8FxKmYe7Hhu/IUXu7WXrNaQ+qikL2
bQUqOucVDktm95SWcjQ5Cx9YvzEuUrkjYlpGgHSq/GNX8WNW+RrO3kWHgOHrXl3H
CIQ2NfQ5ckYyCKBk4yrajscniaW64iV73RNn6CBLU0CA0N89UhYTI8oziUe6dx3l
WggAnBo+5FtaQ2yDcSqOTh66UGh6NPc4+cpKU8MbzKD1PCnQHopIY4gZ8agfYSvD
zeL910jm8QjTtY6kvuPVvYHHnuw3Gr8ZjEwHPavE8D6Fj7bhxPJ8XK4crTJKlCTV
`protect END_PROTECTED
