`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveES2zzLaIjpZfYli1isUmmwGNXb18pxN+UNhWyHlaXWb
WGz/t+I4bZfSjTpaRg7ZcKlS7oO2RzW7WkNYCfS5BH46tKw7C1YhIHM/7w5EDu0M
Jeqhqh9J7nJFDwQ9faCSSo+glqWcV6Q41UH8Y1Gddbl8CqTpZTl/3AtcS+KxU0iT
YrMmRSScdNgiCQ5zZzKmy0SETDqf4FWZKwP4YiGqI447aGjDOPnH0F7mZ+oQDjcv
2KbkbzAKZ+Juirc4IVPR084ibeK2xRuT1LGSVppH4M6h++EvdfWynh0aCtCQy0Qe
5HcBviTifN74VWrxSeGXmr4eppbe9FANf1nx9vH42qkZ+xsxqptkCu5WcwI+QbrQ
3OkPpY4Loc7hKpGeD71HbZVuKELPlx99IH26cYKa476wamWdnqRxxjZwkB9QzxD/
wQ12XbIzz00l15BqZZBvhaD3+YVHR//Qm0nmtqmlWmTcAyZ41xbqTFn58F17bWWD
MoMcWpjhX4k9q/RO1wsuEcpzoCuq+R0N9YJ3xmroHHCQ4bhIfcXIh+w4w5dfAZpw
kkXI4GWlrF1zyECb/0X4zQ==
`protect END_PROTECTED
