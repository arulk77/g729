`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1aS74mq1I+ALCL8d783YZSyxEUPtbT3gWtGdKRFZqItRh
Ds8MLJioCmChhrL8qMTOyLc6i6bSA7RuBco74GHm/2lvS5Oqh1wNuxEJpe+sy1Ii
tRWWUq2nQm9uHgT3IzLxFzJ4Ti6N90ZmbPkpf2TsO+L2IRx4pqdO9XJH7Yy1BnLN
kw7jp5V3EA3HkcIWE2lXHFaOIxDYNSgPCLCNI32vsitKroqmIimJLnyiHYO8g62M
EifPzH5r6lUXphoYre0KP3W6Vpo8zjHxyHuYDjTG7fL2xejUyc6db942iKc0f9AU
gXGnMwJkaW4JJQxeT5NNOT8uzBfp9NTrN1zWIZ+gf+W6Jnf0ttSUcRcSwOoSdtis
agYLwV1fFa1yHwjkApDI1OESTraGk822A35i+JJcr1Pyr42LVqHWItK72Mt5Vdl0
onGq4iPoBejI4AfCi058yW+GTvWMevK0+0qKtqulu71gZJ7DqWoTBVJUpcJEbkQF
dj63RDuHNSjvBTT8FKFobc/3XXtoDzX6d1t7Ayz9Zu/2i1bwx4+qsENZ/q1ePlD2
tPZbGLTF1ibLEihBP4sURr2B9uzLYd5Nn6FonKVvrJuHx5dwcx9zrApJqcuS0pCH
TelJ+KcQzxJAD2kxbhNoJA9g4DRifLKzq9CqyAz92+rNTrv/HMDg4MlgsYotV7ps
NMW46HhNhp6j5/32Cizd4+RSqQ3DV8115rmmxFXuj7PlNI0+DfArsV2T25BmX0ku
2ZgNZo0IVwzIulNk7Y85deFl0A5pTFjD2WNCmaJTrNsBHUPVT39vigRnCfXAvm8Q
HZ59i1YjHxm+K+UOtVMGSfLuGGt98oZoqWCJQAYg20N108kUfrxBFOJ4ablp3EPG
TbfhzaK4PqtCrJ3bTxfGko9GTQkQyHziKfYZecQtWBSXuQ9SgiLbD55VgxoHQtwX
H4wNhW62rjpsnIdikFQtD79LKwbNOYgr1w/ogkkdYwbE7SQHzQtI+Y19hjZ0t6Dr
eI94TZZvcdH/MAq5rf/78r/uv/1gT4ZYQsO/LC6j1fMTcEoKRxPjCRrl4aAhoMfW
oJrZwLIPH8Qd8IhAV9Y7BA0w55KgxaJWm2L0/AVAckm94y1itA/tQPycsv5mYd0G
6KmVMCrPaAOV2lU0t2ZRHapQa1q0Bwvj2AHz1P9pW/6DRODZcatCrAMBe+6buPvX
oKPyOtaFl2rFoWQAvhl+vyfpA5sMP2l3eNqBqA8FckKoBh2Jxxv44sSRbPyoQrjZ
iutUda4rW7jttOLfAl0GRXKjymp6TFGonTyXanFyvg95uYwzz8CMCidFQA5lHI1v
015/xOZ74+ZErDNZS/JTLAsZ/UNjMrpGVNHu7BgODQHeWF9qXESZfgaG6Ir+0OtD
x4LB2+QgIHW0deiV2cNcfVvYIO63hX0M/iFTcsL1VLXwqzF1xiI16tv7np4ic4Hj
sGWIvd7zS6BvfeTeKIoNpfJmkObl07ZAcl5JuZ/HgtZRN6iM8ACt9hEKxCLDQwKJ
U16t0098IcRTBhDkCt4Xqi5Ly/vCqsQYQ3fmhmQrWELRVKmzfabXQC70ioTnV81Z
VGADhC6CGdL1g2l9kpUAuPY0px9SNZtluWPwsTR1PtSGseBnVLEwlthe41ZzXuDH
W8WAGLbW6PdV3njkRNXSt5WaYp2vBPsCaAPFFpKr8QyChadwfPqswWIlI/+v7Yv7
PJAMS0AOqRZry0JZBLH3T+oWA39FZntopLbTQ9LPbv/7ynHg0d3m08gtZefnUiPM
nctzMPW+svvETEv89mWBDknZx8b8yf507326xMORGhzuavcqv2+lTpFQ5C4psffp
/xOwMBBjFTjKDA/8a/fFomdoTKa2rYtdp80BAWUXRdC+hBc4yIzFLHcEgyIWwJ/o
sahAaK9iwIN4TWZC//gVFgamYQ46p3aos0ZwuuP7v1cfabXxS97VNMFCYX2/hOTn
5RmZwnVHSshPYkZgwN6TQVmJOIL3kDadg+JbSPhBw614KTXCtRoaTOewtMiHb+FE
ZtMF/MKeOW3dGGxQwfSHozUlJKnvlHt1ZPmAGQi1/pmTaiBkXTlfjv2ULT6Rx/3C
KVINBPqjAoqX5K3xMGX8T3eryNZ40dk+P12kNwnc06PxBJQKdp1pprgmNNFXIywm
vx8H8yxss6KRuUQM0WySnPNPuqhApw99+hbgS384/zgqwaL4R23c1TKqIdLjlJcb
j1FfJXiETpbu4JFhSZZ8S9faTeFDSomLzrbpXdW6TNPQtA6kbTWsgeV0y41MUSa2
XEbjy0z8xE3NY8kLUUp7Xd5RszOZPZEdhSTtyeo7N7o2+2lK93LSRXZSqJUpS4nD
xCz+sHNxIn7jL+KM1w8mVsUkIHiR2xy5aWTt4Neb32CBU+52qs9uoBudtO4medkI
Xlivixfz6GvDh5+X+XxxPAXdkC869n2Eaq9D+yttfl7/J/JESCr8obBdk+WXCiG0
98ALqRP6/7i1cWaosMtcJJbhNoDwbLHIt5fpaphry69U38B5KQ9o7mGFNKUZU2od
7x+diVFrBt/MkzTdyIJWwKuh8gE8PGDIG553K+AQBIDHlWjNMp8JHFRwEuaLZ8th
3IXibUxvXhLsv7GkBqtTn2Vkbk4XbyYpr+Y1hjO7MsONBbH2J9ZLchfQQwfeoxdV
vAAxPDo4X/MDYgh3+R19hiiSN4gpPPq/CesA3UAa9iZ1TTQN8psdp0V7zFWbA4FQ
RH8aG1vU3WykDbf5ykug9i5Pht2tVjVnVZbORgY5sBAeqW9MPFe/QKRDWanwdbxB
xnxXGpwO6CvZCxG+9hCfUILcY/w3NlukYxWwYs7ppLP75z5i8FZXVlOeJzujjXFd
vPvSbuYHRXCMxetG47wubnrwhS6DGqvbHYK8jU3+0xQ72GOX/05fQoqUrhg5WoDR
XYAxu3Mw+pSL4drg+cUsSyf11ckFCch9PsoInrncYoYCUf/JJ190swOU+PaeCe6u
IMOHaTmAlTaeG4ojClpANqjVS6rQsweb2xo4QIV6cEEvfE4gs7LGEhx5e58ZL5hk
f8afT1H6KDimeEyrh3bRRaAqBVFXt3R1/hQbNDutTgBfVeCSeqEXu9PpnF7eoGOw
8LCk/WwMIrmpbbx+zdsnyvr4etWa7aZqYb7KlMVHudEUCJuCNKKHh+sBpHeJr//E
s2xFPJNlgoWvIhnR/pTPUuZ22dXo1p+3hVZwNDIixghq0DVfGyBYAafu7+jZi+Ba
9cqjnsHjdPKYTZfy1s9yD18kZB1uanCNc4cjriADepvHaIBQaDvgDVuECPNEydR+
2YeIcOtNllwIdK7SpLiuj5cbAaU4j7o3yJbl9pW10k0gqy2B9jsI+rvQN4HVnBJV
oJWdV+Ffubar3f9FL9toZ6ZnvmgL2hJyBVoYDLK5boz5+nwlBBLbUNwfQZkIetgK
9t0lNmIlYTjm0n7fXuOGjjpoH3nlS35tjkmu3pPK5Z+siTJRy5JHnoNAHckYiYqX
0L1ctiiQIppUxy43QLfnyx3xQQdLpUqr+02BBcktuHplhoH3mSOEMeadDDjHy1Jq
R1Nsqhd319ZUn6fTy0X0wh/56YELydKMt3ZChAxCyXlF7KIZ8rkATQwTcR5apprC
DTCAyYouG1e+iaFBuFxICZuOru1hJwivx9LCdeCSAriuCUGbu38BMmEVonm2fuii
at9X5F9c2UjTFNONntgLWZWWf4o/PohYxu1eb9ljj9WSfFmMGjWTWLpJEleLbkEA
TsDXAVqOzAYac2O7aMFm8WNOcNk1k8SqJP36597tj/Tk0LtmEjyg8A1jKrYZr4TA
LyK4PYEv5PN9sd3N/YleBzL/SP+KlzCh2GpsTSq5FAap7Lx8Pf6GlHL58s6wXxv8
UAXhOi847udw1zhQqER/PiYZT7y/QxU16zsInMGrah3W2Rh2QGCAYJ7x3RAT+5xu
OcS+fArmTSecYexPA5QtfVev9n+8pay7VtbajSq37FvrCgfVd4xh3LcfTjI8UIE4
q1bjDeXChAnXz1+zzGRBkE1K4LYpeltZVdeJst0JvdYDLv1LUydOghLOH+FoLUnB
f9COv9bSih9NPx5VwmFx2eSV9eWoMn/hwTI0WGrv6zE08bdyopA6qsh2qsog3R5n
AvXA7uKyFG5PVQ9vuAH2wFtF454PTkNOB9xP9GHO1itdwtpHK1OVDYXzNnorQEWY
n1d/xvU7XQovEnrwmoxjH7yLcminuYBL3odYGzThruwZDINYU57qXwAEept33E7m
SPGPEMrJR6DeVOikq/EzCKE2rY/RJgndWqjLwL9KprTRgEn/fFw6TT/BDnGzcTaM
r2gHNlLtz405DQrasDwQwbdjV6fqdheUCKvaWs6X3VbNEIhxT0ArY470Au9983VK
ZO7DCSJtFh+FqEzKSMaDJx3rf9SFFK9GVxhUXRJrVdQLxFDUI0dC+SeqAVMSrtv+
9mgRGY+Y3j0sy+9bTq+K6yvZRRo0TCsNLHgolvHMgU2PbGJxXaMy0azk0cANhonu
hyFNSlDEq2wFJpwfMrx8Q8K0++hmNJR7m2Gi+jO4j1uGivzTzmvZ7k4/zcE4nwgd
EKL1yfwYw5L3nos3+wrVyoM90rmRRU/xzivSMM4tSKuKc9UQAg2/PVzAVRkc7Vt6
4PwIb3NqZCqOHhfuhEIGhFprJE29gD5W91E3KtrPRm/UjTiWeL+KvwGO0lTYw+Ct
/CxpkL9eA6BRMVscoDDnyt7Yx7w07xJi94nlBvUa+tpRC9R/4wFcKIGXscxMDMs3
fRSX3GP0oPOkAqgWtOZtCWQZjTiYSpNrN/fEO61Vsc9h+s9HGjEi2GUUehpmjvZw
QHLUYFTbflVfROUiB6NtHSWmxb3cWCfA7a9i8qXQVwfqgITvh0OH2J2p5p3jc+jB
a+4NyXWYwPPb5krIys5tfRTnjZL2tXDgPRdpYMWW99Ds8LU1rN0lo914QmsifFyu
dNICJSHhagxixjWBi7iu+KJWqhyirtBQ4aL+3mr9JidwasKmCPs6eIardwNDC/Nr
e0Jk8MqvXmdsNCAsRkqV4AhtET/3RKBjb99XYh2HxJPV5r2E7mn4l/yXc6jDEvf5
LvaFwhJKJ+DXKk8aPiTYU9MT4nI2Z6rFfwKyYiBftJIGpBteg61KIHHwW7wumh4g
bH4EsCINxtuXZNwoSxZnJGDahrxjNEKTXcWCmxiZ4+2kpGHDxUxwP1Jjy6r1WJET
HyAo+SEQ2P0U9mls8KFu2bOAbWKNN3Cg5tLi+5sxRcrgNvRGcab0TBSgSNQI+hfd
uA7fzF7EiXS0dd/augxc4sea17xJ6ApdEZl+uu3M1HNBdukFSAru3kN5JadvY7Un
EJlKNyUyk6Um1yvxBJOyhJjIDhTO9BhNBvReR1QC0mlDlqhq7b6IyLse4h80pQpA
pyAInNKsIAAIp+I8WgxU2wN2Q9yf0tVPGe/MQ8PT9KT35S6BkzVYvGU4rbv81MYy
heRghKWrhE7dA+xmm6TJelFj+WTQdTK6PNGG7g5qyJ4iOO4dcaes6Gj5pbHpILxZ
w5OEQ5wWKRD530c7ZRXf1O7b2ay+zYUzheehBn1w7o3p1JMOYlywJF6mDT+fXMAw
7+zHtQeyi7e8yBOavgCzeCvDTVCQfWfZLAyZRgSzfB8wY+ff2WFpzTgc4P2jvtEo
iMfU28L1nDjxTH6R4XvRMI/jTQkQNZhHRJmVlQlxsZLjYpwXtTOudbcK36TUBb4c
FdVwMK9reIMMZjvKdo6qx1OjwhyRxFaLpeDTWJU0OK4eEJdpSBoRihaQVTymdJk+
OKf05pbKZVaI7M5ItSNSCt7uC+PeHYIqd1Mvw/fAfrssWE2r2ySImZBCLq61Qb3F
OmmRPhHsuURbCDcSVq8R7NZmrfY3WiucAD0bHNEkWWcJtEwBFvOkK1c6OWgyjtF0
CkIOWCSIx2/OjlfcK7RtMyZ9m7mw+kjazJMlUNKmURQUsAuQhreYjdbDxaHmWlfs
GzCPaB/qtx/GYpUIb+RzOtet8YU9RkRTTCcCxIKaYMZNcCygOzTRJu1dGSYp5PWB
Omd9Oz3df2yjjATb20r3JnXq+HJAwyp34jHC+6icp0MzG6RddrfVgQYhhBk37DWr
tqUH+3F29NFBGG1xFBG8Int0cDLXm18xiYABHIXNorol6FWyqoWR6j2rfjRcIYjy
Z5PxJ+6/592HIDjxHGEvExdRyVaX/ungjt2Uy9fYf7QCEsEpC+wKi/hS1v1PhLs7
lHaJgZdABdY9AVg1yNBLUACjJOHoIICPWlv9soFZWCo+AHOaJa+1lhAJUi8XZOYd
g/BZjI48fD9dNkLI2wn2JwXUiEBmUewSz8YRHUs/F4dTw4d66a7Y7r0A9MeVsXFq
KdA1pwjrTNRuNKZ4GYINhej9R8f2BaDnTqJ1V95A7FZWGt9gm3cg6GsM48uQsX5E
5SPjLBbYZtxXaJA4s23j1xjA+QqdW8CmJUNPP4axQqd3s7dLA/vXaice7+IAsViJ
Hf0h2S85UbV5ZdMWBs/wvhP5lJyIUheQ497IGcv90ZBkvIXxrPLCOP23TCWdsOLM
MR/0CEMLyGFMR7ahZZ9vulpkYCKw3wLAUNDXcGUSJPIGWC6IE6zxJgV+8dnuFFOU
yjt1/C6Npu/wXwxANWaZdJZpfBcAUHGiBsXkEW8lwTjnKVEbV4tyLA6rCAOaa55T
cDITMFuylxu9YUPRZW9g5HpBKl6gAs+GmJw1gHc1ZOHcTQxCDL7YVWjL9g/ikZ9E
L2mmPaMxsngIBKYzmghXZzHkKPlOz/my0itkrU3WCqLL/KEghZ04fVpxNY2fk5qv
8Z1RMDWT46HaUU2SwkjGveSN5SgY7KFTbbqmDhFJwwOzqyUArf1fYymcFkvu+Hyy
EFBZyemCAKhza93UWXXqrCmP9pm1Iel0pB2CxdZLM4oJ+fW3M822ms8CJ2RWo5O/
VR91YtGPRtPm7TBQyrzuL2pA3baDdfnHEK4ZMLCtohPw+N+WSzCtgd+2hSzQJfJp
zg/MfaRYUR440vF0GxA5AXqNzur1ajci0l55bsHEGakXIGMk2NbaJbg3j6+LU1PX
QU11htXO80/tUB3opaPhIHHYP/DfNgXahTkfuc/ylPEfNJlwwhuS3QctSiWpNvx8
/nWEm3ge07a0/8+Ut4fTBl6ZB7+PP1sLm34FZ7bjYrC+jYhCskkyD4IHwimxvj1+
hVQ4BjmpGFU+4Z8oW0cIW11L9BoxulsWo8dObvkvhwFFqv5mCBr0QxANxsYSpqeV
o+qc1LJo7GzaUWugkyJgWtcVhpGCyaYtQQIWy/UyEMTeemg5mTUrMkZPYYSCQIsR
L/cf08jkYOz7ZmNxt/dn2oxqyq9TY8H7KUostSyTowHYKmoTKRxHEY+jf23yD6Nf
btE0ITciy7Q70XK5JPzQ7513OI3PMjaod8MRwTmn3SFOYKZcXDKjfzKdmLQysIlV
ua3BKapyPxKo3wtHn5JMJLCXHvytB62s3o62WcDD+tZXdzFsMKvZAQjSr/Nsq6+o
JVUeu+nyuqEa5rTHayEJMTlzEfdJ/ODAPpW1tFpLTxFSBmAzFwrS0gkiD0AwNkGs
nP+u5PHORh7BBKEBsxqukPmPs+5tmP+hN0Oaaqeml0PcjBR0mToryY2gBMLoGiBs
otRsq1lh8f8aIYYhMSCTCG8TJ6lBA7sQSwb4gyaahTiWOET1U8YX3Q2Gaz97GY4T
kblU6mEZCuj6hzIaC7Fo3GqguOqFWYvf+tJRJEots8QObGr48eD6HPZjyAYR1Pye
OAsR0vkOSt8X4wpivjXUrlTvZeOgmNgzvM60x4aKH6usRxSMth4nE1hjWlKSuYar
R3o6uKBZngSKhpKn5hlI0KxxN92s8pmw6QrcYNa41KqcDOAgWYk5hedIM2xEbdOl
xD2JEZQAlviBKM3MzkixAqT8K5rWqB0b4du8XeE091svuUVXO+dpN8k+FgfAbx+X
9jY/3SbRV3o+0Xn9s1lWs5oI1fgW8C0gNRE2AjWaKoFCfmzYG3/m7B+9GO2SPlFA
rjePL34MEGNy9aahBCBsiPtQgNaMc9AmdNn8gdKz1VScr3t1EzV048m6KZbJmG9q
kGeFPG6eZtDQZ5Y/dodGR2ra0OyRkZeFxhJmroaOGqz1XUm+cqwEQnZph2n5I+Td
SJc/ZfOzNz816j8CTeQUH4z7SHfp6ycLN7RCMhPABn++IXmnHYkjS9/ghdddKjNn
Nipi/YAWoR7rIScZoAHIZ7SWncOYJgmZjMPPfPbKqJgcbIytD2grfL2XhegXlgnN
L77DAS4aAFx2Qo2p2dqBGcCyxbHF4+roM0GtWpt7PG+9C+AYVgFO1QvuWy3e404t
gvvh7iQqxK9D04ZbFoBEsGAtZxh8bfUk2Ki0MZGZw7sABveG5HJDGf1D8jZdPkL2
vuquu8oqjFSZb4AzMJELlL6Cp5ii4c/DzaH4Oo+b85GwhWYebwMZqOoq61r+SJWp
eutjaYXcbEUieppiDsH9AhYWKfmHiRAFdOlDQ7cuOgDKWYDWaq8MOUDrpKcl1hoM
YD1b4B9tcM9JS9iXQqQWC2A3b+4XFgZTJKgUm3T3rFvgLrytEbTb2OI+vjUakks1
bQOkx6HdZ8/eeEHlWtLxcQLAB05yoaToOGGUc7rSL97BuKtEpzPo05dmiJoEamM3
yr5AFNSSRburZv7SdiK1AugwPJ0JgB3Lw9HvmvPzvAK7uh+Zl8G6DPn8Q2uu/EyU
AHFk4D/S7Gxego8ZXWiI8yixFRYU9yL/W9JU8Kk9dMxcelYhMXTk0SCbjmZVw3Ps
l1LCcOgVMP5i5ajf16WO0k3HLBAQ10wxtSCwqWxY8eWQy5NravZMIlr9k7HsEWRU
SP++tSefuXv9yqnSVrhcPcgN7Bot+mXdDPGgqa7oDIoGVHOPRGdms0OVej+ly+jI
RlozCq0PhYL6xD1uU6V3b8plCcuKRm94XTnqC8QieHaaUJYsSergtfEOwdxQzdcY
uj94Z9Q54axL3n5cvGrp+l0AEQl19wEcn+yGDJ9AR7AOu+2tRnfozGR3mBF5ugdS
hTeiwDNg4xhHimslw/jLpJ9MeuHlxs4SoRgCxqrlwcnwpboJjycWFtGsbukSfEqR
Nyfem0qglvsIP5IhRryO2S8N7wGpBcFfhKE7TQUzICeCx1cn/bCuZMF6jn6cICCr
OB6U0OsR6575qDQPGG1R6uLJ0WYrwLgqQZ2SX89kBASjqIJ1PDYvw6Jwlj4fKKzs
AP44aEAs2ZtgKvINy0WeVqj6mP77nbsglUvEHFpDtwxbVXBhOD/EOEa4+w3C1BR0
XUH+dfd1jqpZnkyzdARiBlp5V1KP+KnT8NUDk6lzbGYUwexAz3h9l/dIl7ro3p7d
hVIggalX1YGK3TNdtvDvE6qui3zL0+UO63FgU4z93sWndNWn7lrETHaXL/odKyUR
5rFALCXpW2FpKZKO5qUDyjBjho8sEcAd95VK0s74Lb1xIpZHc5ufXbujYV+bV0EC
vN6zeSgS3pjFStu4eB+ThuasDiHZSn4bC3RC2olPwTgLS+kyCL3EN6Qx4/171rPt
0aKyKUDJsCeFhQ8p5ZRICG5rtgAGsmghodKVJo3PKklh1E8WOZ1Fguzds4Ai19TJ
0QlxkPlYvi4JiJhg05Imc/CpCrLc3grdFnntEkxCAWQENdUpu4quW5GWcmLOyaRb
YwAEqYM15gpTo62h65HZRXjnxiFiOvhpL9tPSye52Gd4+5z1g0fc2rWGm+GSHbY5
KPcFbhb5YRMe/0CLEJwdJzMjgb8FOoOlaMlCqK2b6fqEUPRm3fJyTmhhVbDxaPhY
+RRfx7Vwj1C3md5nDrhPHn+UCBXUz1Q0UNtpl7v+XHDPQxq6dFtrP7yarP6eCZFG
1d47HvU5nWQTjWs/EYKSSUs4GQGTca+vvu9dOke+W9juOg02ZE6QEKdP2TVITtRo
bFYoq90uvkdyCwQbpmZtzqpDQlvF2Xk4QEPm8vDYhStjxhVF3S6rnVdL41AVdASz
HGU0HBxze1fcMR1QOnxsQ3OMRAFXGkQHAcVHaLD5+uJR614VvDpwGVRWMCP78gQP
8BiaAc0utpnOsgCbQETax9p8OXewpT3BiYvhC0mS9SPzHi98FlIJXoXdI7xsZyfX
AVaYoOF9mdngFx4bYGObj+LscjguxRtbql1QDFShkVHa9D84Cd9l32FWG1006mIv
+WO5NG8hk8vmivOuMjIszzzUSMTRoZCuJD76Fo1VqsZvpbT+WnB/v2LEsHn1k3KA
V6eU3JArAQCq6ZdWZdzJdVP0oGlBXWV1A6rOLg3C77ldnYUiO+sQDRWELsVq750y
e+7SQ5r2m6kCU3j++j31c2KMRhofE5uVpnPGxAQMT070tthS7J3snGeQKqoYEh/J
csnNKA7K0GPrtUlWPimajRU6BAKtTRjvsoL2LXWlyHVKaUutBNJEtsOy/++Jm9xQ
L1jEr8I5j9JeVX7mIF2J+04A9F+JVUjxTMyMUOwziM+EcP/Qv5kglgSDXYNLDxJI
g94nWZ3mZ0aT1Fi5km4N79oeB7zQW0gu4YUU/2e5q+Biu7TJ54VYV4OtDcSLjqEa
J+1quYpDfoKJZdQxA+7lqGw7rMWd9ijDhQTDgDF96vC2Llwl4ZtPuNijOZertVk0
YbxnAqQPUNMdh0utXNvkY3ovg8Ka/vlXT2LSbHOPUqoOtll/TbpHmTvWL1qyh6b3
jCrKDK6TN6LnJtziOa98g+VMefHFPRRMf+SAmLirSgndmRIuTYVoBa7p52Nwd4Ls
1s91o54AUu5d1eCWH8so9qkuh3bhueaAijCKXzN1YiQBLzIyPs1GR9QeawSzI23H
6XC0cHd0LBe2azDHVMKRhoj73EycLkZhzqYEnpixbGtfpHZlu0AELmmxdJAnoVLM
rqWM8kjGxiPu67hCF+e0bEsAyZENQD1d+a685mv31JbVKf6YFULTPMd0BIaHtoO3
uUmRgzGCOzUbj3NBelNwfIJs9oLt5IOzM+dKlhyau+2lGIQeo/Cju6tZsm27dBVW
yTJV8rrLNgEf6ueChEvshkKWdZWd6D/qwQhjGqr02oXPxhwaSIqodGR6EJX1JO9K
XPCvg8SxSjjby5JajqmorlLKJI/f4FyhL9AvogierD/4kcg2hkHW2UWQiNbOy2DS
BGYDRcfT6gfIYyJ568NjpIYaf1gczVllzb8bh6MQ6xi+qhETFezQ3TxbaRAE0RCK
a2eOZFZs+P/csB2twuWzOqtCSuza0iKD4zrnGeIwQBqtBfpjBsODhF39Ohs/j6YA
sI+ipMBnGvi4Az1IlhTi6Pi0ToEh+peqE1hZ1ChsosMUJWyfstcgLwQjHv00vNia
gmO/bEFgjh9GjylI1QxQ0FJaHyOfRPFR3NmVuhy7kPXAluCAW/Zfap/OHTkuEtgI
j+L7UsbEIrRO5od8jmekeKfIVwFB5+pnFUTlxwujeL26oath1QqpxhAgyRTZTX4/
yteLUxpYlJxmG0hywyzeB5qqTl/SwIcX8PrfUEl449Qnq+4MVz7hOjxvbz9NU8vA
ZRlUmw8+UqU5MH1vBGGzuYoft9MDsNTLQW93k4MUWEkY6F0604OfOtg9Gl9H9mMk
94DqgpfFsZ5iI6jJHbC1NWPoGWJacT95JSmviyFRv6Za8/mT9MzJok5uElfhbfRZ
fUaSKKE95fi+sMjGa/ppb9o/rcY63k2uZJ1VJ9S3HSWB4XK7E223WLyAd+g9TdS2
0vd+aSyIxieovHtqF2Ll7n5mjb7/MudTJS9ODxy35EcNEKfD7M0uWHbjEWJF732D
qRElzZFoK+MPiFlnukteCkSM8Uwaq2lMFyrkkAt5nz4naZWkagUIoGslEyITsFn2
pX/u6IqSr3cef70ud3xf4Dv2PJxEl2piuZZKig47VV4gL/USAmiG2v9R9TkLjN6e
Lhtn2YIyaf3x9J5xawf1KoypYxxUA0hrG8LwRtodxQP7Mra75W9zvltiIrzdX4+9
QoEMqs23OTUlE55wnc3agLIxnERmXPwBK/1VLIPm0/IlU698qkisqFXvpG6kUSYL
OHna8Wj0ypqpsP5XwdtbZdW7H+iHpgH/NcPQ+vx5HoVCIS/2Yk2CgLNvaoX+aGTY
JAmmeA1yJQ+wAOrSs+3UUHMYRCPuyAciCr8tt4PNk2g0QLxCC7B7c6VhRAc8h5WA
Cm9eYSIm1fC+RW8FlU4CGcyvkWc7YnXm7/dImbgoZFOhc8vSoKnOLBtU4sYOvCGu
ZKZYPWWtItvV28rnkLal9iTvQxEm2GcFAKy/ucx19Fn31+8UDzyY2nPf1lL4N9Dw
1jHaPqpMUzimLJPdURBWBpFyrtljWLXooVMcyLN8vOW1dd3imZVkaZQnsj/WqwDl
BupCAH7q+4qXMu2fEXbmQ3Us57albuyHKQDqJyHSsoPm0jhVQW/fWZziEbx4hvQA
K/eg4eZ1VBLQkrz9ceXvhXz3vuTKfe6gUH0WIJrUrkdZJQnvMOHBqOrH1Dc5yfsJ
j42PL/lfDXLz4Kc0sTJw5S5IMt7yOD4ljHZjVj3mKyhwak2BttTd2bhezKdxUePr
axP7YrOVYqHTh/ddPfviZ3wYXFAdkqo/+auuRJRQ4GOOFTZ2e+NgofzWACCq1cPB
uCW3xcOPBj3BZ/uEdEsRIyxYYNwMtRIoVUvE5t2Vwa8fsjMnKmNccWyWmSCYfuTS
85T7Izewf+dK8BFBy9FNl2eEz5J0wQnGG24Y8f9DAwecVCSd52LZ5Y+SLLtRej9u
97gga4DBti7LkvCXbkbXOQo66AV8gUw5x9Tul35/yQQ=
`protect END_PROTECTED
