`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL2yPW4FBMS8tbq3Kf0/Jj5Y/Bat3Vt0Z+FVwBc0AOOx
rE+8tpQHrupcfWjEGq+UnR9U5QZoVjbzcVs7Zkay9c16fEOwpRvylo8rPey5/y08
C8FCUFvTbZZSq3zORS3zi3coxkW48V05Af2BzDzweoJtUZNEpwH1wk/jCvQlLwmi
7gMc0ixzQ9VuW3ggfPtsB+NMUE0h1qqxCCPZ9fvwMObeplisjEnsExrU4nt7ZMH5
lw+3GBlqbQ2XbSUGsCuP1hliqQxKuezIY7VIZoRETVjqxWLnVfQPyjH/GV9buGG8
Jplr2/jXToBEx7Aswbycmw==
`protect END_PROTECTED
