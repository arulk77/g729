`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
N/d3BQ53pXgyqAg3tbS7YSm3ssjR0FnUrcf18+tczpNgszRTdJ6jRtCx3ROrz3P5
G5lsKMdd09zmIhFlP9rd84R/YgKO5ItF6O/CHDRB7ko2nVJAlui3A6XEqiT+oLtA
2cTKuIuS3+jnHNHxC0pAHVZe0y+mfykZiMTXjzjpUSGMQqerKNSWY00t3Ah1gcYt
lqcKDH2HmWdVcciJtF5+1JC+yNwUUVHHANumySdTWKGxyZkDa3+p2b1CFfyxMVIH
9Noh8VgoVREG9T6VArtGGp4uegBUtd1WuDwLhO/P8fMgN9m3NnpnhgG712jt8gcD
vOQXouo+BxsNUwWCgKtF0/hAndFMkYSDXRpCTbsk/hc=
`protect END_PROTECTED
