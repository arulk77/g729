`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveDNmG5WmQIG9D6WiUo2QOUx0Fje3cYT/BPzDhFKbi3BN
GVOabx6r/585Al66oTbc/LjorXIS+xC5G/48GxCWQ3Jnf+TGsFMXval76aKnZXZS
Xa1IAFmtU3yjl65aBdd/fuJjDXQ/A2E2tEGQ2idx6OJyDdEb5UsF8TNgY1Q4wfbx
2g3QnGbTlZjrmZnN8XGiSu0B7aJdf93YZpSUjz4y76ChAsefGr/TB7B7agCEMffi
p2Kb7zU0SyQiKDPlzeeYJK5nZt8tFiIeEQV0b4uKBl4ud91l7+l82+jVo+yDxkzt
IA6ZzehGFysRHp9HN/5uiYFwhlsFEEbBTzZ34YLIVU6FLLfkpDutE4pAJuak3yJf
vgJqb3Nq8rWXfkm1R6Omh/R65dQxhGf07CQY8pajAeHtjFJrYgVf79YroA+ocULi
qBLvXTulRsH9zxBHnWuHBLsVi05eRqVoVv2xVXnlQ+I/0BKOnSW4HG/K2SDqQzk/
Ug3AHapRR9rBvj1vo8oBIUKur8TeO1sFSMlRdj7z4t06Ls8AYqkbTxZ/rhHCLE+F
QXmkry8Bg/p+0peT0tL7xbl/H7JGr2yEcDxDZ0ZypbhFJ7q6ukhJJRpFcDktRYRh
W2VMRxwYuz8NeSqtCHXd1ip0itVePwgsuyvDEHBTGgvDecVgz+ItXL3vfm7ptuy4
N5dLd0iERZz30gwq0G6cHyDlvlqdQkJYCRfFsvVrQHAWDQK5RerbS6Vla4WWkBRv
M3hxi01844uM7rc/PMmuIlyIJA1Ymw9RB5Kk9zB1wI3JB/wVlQKuM4b9SaOfPWrn
oAlDTgkjBVx+hrZvR3WyevX6xuy8jQ9pdQ6c44qzmemhxCvCgoIR6ECZWxTL7kVb
H1YL5bky8/2T9bvJ19gIFwgsg9ZJN59+zDbh/2nq793AaBJA3dWUaCn4ybNKxeFu
/4UrXc+rWTZpM0hdkdGeFEhUrCr9i0qO0DbeGtS3c+OdtR8kbrdF7kBrNb7njdHB
KmVgvho4KWH/w84no6J7J0zUoFh8Iirv7vtIOT4ccY/dCkNSzljTWHeic1E5T3j6
dkSrq5a6avtzozTOGxLnhs/zC8QIpPGxIsca9ZZZ0gMzpgvtp8naIXeA1zEmKbci
TPxX49zSqLQ+Sn2k2FW1r/yUokvZoDe/ZkUoTVp4yWlfVYf/R3dyb15BUVRBHeQK
ZdWmmYdF+U/4u4Z/F9na9j79XtRng4XSNoNaQGE6JeB63R6Jszuhs14/VDf/FcLv
B+h2AeCiHxVTdk98QwdJ16I4Y2Kr44cA4zfyTLQNkvXDL1IuZO40G687W737kmgu
a+8xcecmb8yvJKen8FMBWsw6FYiqzqgiCvd2OpwuHoIKGeO8JhKd3gcGFWihUzHM
E2CKH/bcJDqaPYQUAOagn1VNrPIz9DiA/t+4M87xhLySvGpISzAbQ78R1Xuyyo1a
E4/f+fbMcK5i1iywed/J/n4KgygMjOmkZkbZVXohgOocbzaV++96xBOFmSOVJIVS
IMm27lr7d+FJCTqeB05S22eFwKK+kw18NzuUPX2E0tez2Xo3m48ZBw6Hd1uhuPpj
/vZ0SiyJ1HYPho5SH/smvxXcGNHeowXNMDCdhUYBaAJyTOR4p4Ski1SNzC8GyM12
1B1FFy9tEdASAJCYlPG6Gx2rBnrNx1GJYpZ8TnQCw7HTy61J99z1FMRXvh/XkBRI
KZrKpOy3WKRrT6DlamFnN7pBOzhxIgiiAu6RM3TDtrBNhmstA7sDetwWsPeSCajj
Mf5Y0h4g+dxHZG9l1EIJ17dpWqzBS184r8FNPMl6VvbLeCzKpcG+qlnTN0ZZu/i0
yzeiik3WdQAJZxl/PthWkEl0YnziuNw5L3m1u/iYONQeq+QKZ25odoWPUEBlWzQO
Kbn6FZqWRxFSeIL9e6dMn+PsTlR301wJ5mHXA5xcXxzoawELQU3ZI7OMAzb+IscJ
u++lNNe/fwZUu6NoInpzpKGkqVr0tcHLIWOYXBn3RuYbMh72CsLLow/5r1L79ZT/
wLSl81opMDNFg+aTGqF6kCgLh2G3UcnhuZVmYPq3Ww7YDxI6sGdmJTm34aW5/q8e
3pKNSHGskmQFa+A3dotDO2EuTbxtnjGWmiFI18kQJR8DqqWT90FvVsyQtKPa+jxo
ofe5Lh7RJRmEnAlBFcmF83qBjEOIPk6eCHp8XpgJGrAPW+fTXiJ+LgtTTTV+yKgT
Kw9dsxJTGt6MXDS6glFtNQ/v/BKeSNo1h6LwRmmIuwwggFpRvgBkWuaufs6V1Bl4
D5RTSD+XTufi1dDxZPfC2hobdNZgZMBwp6jH/ivo5PvkG41alSbfg7Y+8yFeotYz
cGdYC2f1ohObhNtkdgiOrasoPx7f4U5aUlHdkAwMQzV7S7sn1jCcetBQwEU1/FXY
aUxgf/oIiwyeO9MKJtsnTg5fB9Vdo5Ie4xluflj/9CsXR726ryLSLy/gyPBdvq15
0CElFQy8TroBkfSQjKqjDhc1qX9F5gVZoX3lrbB0uRi56oGCSjWaGth79xenW6Yw
agLo9CCqtHNes353USET7OPjrlDdF73ORpJWV03oGn+r7rGFcYULLWgcjbzBCHV2
PVR6mNuH1YN9Rak2ExkvIdJsP54yV6EFA2h7zwXVNrLMQ4HTCFMrGKL/rLbBlIxl
F0Illf0OTv+U2fzxK4O53Do+lVCccbdYF59OBvzoKuVuZyFE5f43jVgLcBNvuX40
MI6bvkzjFDva92jbpeY55j5kLwPE2LckLnP10dDjfBD5gIALOcCrH545rLFYISlu
iwZeEimbMY1Bs2qok13Iq6wLt12O2JarIY88MvmZ9Yb8eSZiM5mar76cWzEXVzvA
f6DPXU5mOyIp4jV5MwkFg/3EMQMLd9U/uQRI7NtQnjD6wJA5KZy9KILCp/1zAgIU
clz95kL9pzmrTr8HxWfPNik7vVnMLIByYwNyXDjgPZjgjAZRM22CkCnbvsgJO3j8
gjzOq31HmksspMfQzHGKB6DMZ486WFHAkj6290EAoU5NfCuLFaepZxU7rCxvdkp1
aT1J4j4GSqkekmc8LMu2AOsb1U3UAoN+R4qWXFGCIC54uCsCPYdPl3CoeET8o+mR
sxaBHJr7+kPxZ691njxWH6jEnFFmRR+7Lvz/QcUm9/yxOhH+kZK/Dz5Tm1so8vrp
PpJl03eLGLf5EmM1WS/xzg7yTNpvoU3H/9MYZgSsTJAzdHsuSAmiedOhzTcrZOkO
eenwAJQU+CiOgj9y43IS0ZfCFwgodyw4lGsXpV3CXX1ecaQqs+tppj117WU2WZd5
5M97olCGoSKfoqfJM+5IPmtowu38WrYfbFZkdX1PXSLxEzaeeOEQf2rdmal6yk43
fRxhmsgvcT2LL33qsAw3k+z7dCv1A1VW+oZigznRVocmJgKelERaQKHR3s+lQds0
ldiC/u998jZVXLvf8qumY0/uFKe+P0ocel7xFUMpIz89QQhnux2MTlTDE0ahvOhw
zfZqmT6IGSPpZXQyVTPpmyyrVeHm6qmPNcIynSetB0NCziaeaxo4GVxsyTaBWkPe
pYAmJqmR5KEKtlL8/apKxnxlEWpUDGsHZu6aSVq5PoBoIibfWiQR91My/EJqg42Y
qsywgw9B79+j3sWR2kWvJGiBUl+2QV7KOCdqP1ogNwb3eaXr9O8dfe6/ukYg826U
5cO5HNOfIrVYPaWd+pC89ydNZsMhW3+bZ5HeCmxA7POSQA90H47xGqu4JWBxvrVw
9AP31nOWziM7CKkKuBIyRR5xmMZ2+TGBVsbdKtranCFXkdnvWHVM+sCA3oj1sVCX
H4vIE7Dpleuw9CVzaB1ud0K72e03MSLYJPBP0LQ+vD9i5uB/kfcYCkb/O1kZY5cz
oVWI1dHWZbp4Rr21RHrZoNwx6KEoVCgldaxB0K1fVJXdaoXXJ/HIfZRo6QDguAYL
7TIvyVfEOuDyKtONyz+Gb4l5XLD9S5EIB9wWWIGBDWir3OTyPIS3LFfPYMeuVYkr
`protect END_PROTECTED
