`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
hbj690ncyRpXYfHtfobSoYNtkB7JtP2GnNyXm8cwt2oFj7n5Gn1DK07Od2BsRzQQ
7oXcFh0cUlAkpGrfBPF9CDMFgtSL/IL2ipRQhzXAeykrVdiyeKBtGIjkJtcCPbD4
DqPy/o9lT+a4rNEAOVljvQPLCw0TvyvOM/j2l8NAXttlIU4MIZL7jMmrvicQr39N
79gLo3lnjXx5JVWNF/jG54TeGwc61KMikBICSplA4VU=
`protect END_PROTECTED
