`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu479xmzq06xHaunBrjvYOWOTle0diur6pzW4OhQ4AuFyz
+wUbnjZUjRA8VjM3/IY7lkbppkskn6++u/qnTj1xeodG8+6xsRmUbpY8zq8zeVGY
+x3PNLTAOAI6+k6JfQkI/AIwYSQSIMNxfUWykZO01Cunky0LidGqlSOHxR3MvfJ3
ved5AmS8bgb15Y7pOrCgrq5Dz/PhMlymLGVdJXpbJ9YCXlBXPrnPL/WIeXt0ZxMP
0j2k7KYRpkcylZRaAwrpJ5GTqcVc9MWvdejnQ8b1i6EsoG7rmL7bleioCbXx0/xV
nflKjjTC0YIlfYWH5guCMZoFpk1nBEWEM9XKZM2+f0qycrud41CaW3B6pyzHgYd4
RR86kNC9F1O92JdxfvbyMQ==
`protect END_PROTECTED
