`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveAYKFSkCt6qkz5yBb4qyNs1fmE6h9j16kZGtFmnIe6m+
VoYhD8vwVO7JchXh5WjQL3F9PJc+8wrlhNv4IQqi9zH7GK9Cdmh0Im62RLkxcSBO
Za6HnixiZo4FQejR7izCnXJ3UT9vbKHsUPzvbUQll3f99nHTmmVQ7aC1CNKoptsW
dXxC+hE5rdG76EPy6+IblQqGR45wA/haIWXRQ9JC2KO7JxXOY6FaF61/G4BpXGQ8
UNFyam0c/eCHh0bbZw8/EfvJ3mbYqTnBxSNXMLdUMkFelwJBIy00non9Jq+Rm5p2
N3lCRjD8L+4BubmHFOPU7U1wOTr3DKKepRPHq5FjPayTRGuJjIfd4d9jJh7hBd0O
0TG2FBdv3g/K7PW48xvFBo/+I28gIj2o08D7mMJhV5LGb/nL4kSN+k6H047Ws1vv
CwuIxGWvflxLXrWCSzUJOw2/ZjvbhEaw70CcNOBC9byp93JAe3jK5MrszY0iJjpM
`protect END_PROTECTED
