`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4yk1eNbuJB8FmNlu1XIJmrV3+tC2WqRsZRdy95plGQTW
UVEPXRnuzDCLyBvi6ORx7hFYHWcJb5PueuDap6Fhx+slAfmMPzO+5NIAoa3YW3c2
bfCgaCiC9RLCZ+fV+fvgters685FixVEkkKJJFvAiBOADbWhPE3dtxg6HDVh9EhE
gA6NysRxNmJceGsi+UfMtgu960AyF5qzfxdOtPjRWPqmD7Msrs6PZpZmMrUGHxZV
jYCwD8nhkjRf6E8fp+NiOFkast5sW/0PBGZIrKSwgIvWPUFb4qNAVsCFCjVmftu/
ZJpUNt0rLMThhyrngjWHZA==
`protect END_PROTECTED
