`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveJ8tEb42K3lvNbD2l9sTcVFLzCF1JyoJRI08/NQeD2DQ
Vk/sdqJkv7cXCYjXYuyneYYktaYOmY2VwyKnYGrwCdbpzPOGg9mlmTJd+eOPdyZY
DolubYJGq63z1WUz/iIChIVFAwhyDfSnc9cUMTvBvTUNW03QmmwdOzl2UiKdZ1+n
O1/7CGRgDOrHf94JTMVKZBTSoCeDvcgrqsT3zrKvMVI36LIzzG567SVXsfBjchY5
r8UIvH0KOvKk083ZspeolpCX6ho+mMzl6wpqRk3vGSjHeqyUC0NVwlNTBW/cpxjy
2e2uSPJpHqfisSl6RUqZEdjFFUA6HW4hd0teSsFpjaNf3Sybx01LKbVpg543aUzR
uJTwUX3zaRFmQEGzoftAR6rIWAkdQr4zI+SgbmxI11nF055hOMoLZYYE4ZhOfk9Y
arSFCX/RyoqfQwlmi0bEZL9Rt4r5pzoXZVyiAhglpFhZI+cqrrj/wYiPehkrxc+Z
48XgzADMY1Wy7G+CuuABcQJ8AzkIJDJulq6OrPIND3ZtlYnat6OV9+jGKn14wAaw
pGXzt8puO5NwW/b5cUI7eGcGScTK9owuIptTEeKidrltnSc/8mCJIpFsZl+1MSZn
W+XgHxnNHW9Z9eBPDWKqLtqp/2I3AY48j89DsBFuDFU00/W9uGpR75CGedl6/vDk
2MSLR9pseZuxiECIPFM412yBSzEy8SNLXCN+BfjSvmpXYavzbWBB6xQdZb9/xNp0
YL7H9Cp2cs+Gqstjhch8cZ+lvkpLSgzmWd+hmhEv83ENBT0RAgKAqWIoApUwLOUN
J97B1VKe5u1/w/uFPB4ZrtAMcVbgrGpFtjycvkPpLVKW8sJXTReTQ9zR9ajgjlto
VGzBh0AELMLJDoR5eZu1AhfXrWmAG6qJnWf1tV4fkznBUxx1qQs/Ic0HS0TXx6OT
le66D7zfRLwsdIkIJ5MOkGJq0NyiaYHjl8yAJMYTbWkLGqHXeGCTxCnynhcjrOsJ
KX5fkL/C+AmmMhUjvhwo8wFLqOyyPCZqv9CWwHVsvGtGZVenyIzqUs0LxNCJ3wwU
n2XBkLiPuRqWo8XpQSCCQ+k6J5GVjK8i80ebSi1RNsylgBSwA5QNxXk9S22qmk+u
wCdddXIR9JofBJi7ByL3sRhx+7LATgElG/7+Z2tpva2ZENGihRJJmYULMi9RkVmM
0t7xbS1Rk41wAlJSml782FFOZHob+IDuhDjzaK2WxDhIqUUjbh6pACo+38TLUcqu
7TEJxnES6Q8usalkWUZdPC+9V/7xxzjp72n1lVdC1lHtGpmlXuX5XyeCLX49BLTM
cTblq7U/+G2/zl9qPe7SOQzFiB9PyeMw6jpEwHSBX8ygefjJMU7TX/gBFGief4kL
ikVSeZ9fHfYP6lyz2XA5sZ4KQa/V4Wi+a+pVbOE67YdQOk1f35kG5ohZnfhYLOR7
qEIXlPR0I8tSlOWtS1Lb3GVBHYY5eD6u9hlpzz6stqe4V/JbzlPIjK0Q1CVcwh3l
be9iw6Ba4lkny9Fd79tmwrRakbpKbuUnul2LmT9RCCZvjJ3rc4jYxRPwRZrDMeb5
fXu/jwWjp6WSy/f+eEo3zPgzD9nUspcI+A1K9+04tZIeAJ/Kp3xOl6z/msBTLO57
vh1qfrgV20LIyTB9GZHFv0eLTh6JKtsRwpkHnYx+EC4EsUcWRVu5D2OZwErrogEE
m4L/fC0JTf2+nVIlqLtafYC64k3TNgKQGbZst7Xf/XqgzBf/a4pYWPk/TisvUa0o
Pwasejdpg5Zbn92j1ZxPyUfHGp0nflwdhXwkQRgn5yV+PnopnmbMp8431fvk10k1
xLMgDvZQ1xmBQ3mpLJEOW74zyDaZ1mdGy/sM3KpLSpX5Mg22ZBURIfVfAkQg7Dcb
P+Et3RZYJhW7YIlKTHlzjskUx2HvtrubyYEq4o3HlX6fK0rDJuh1zYnMXovDTZ+b
MCo/UBFLL17kPZfh7RVWmhMRmROtQ2j5zHmg54ujG1eL8TaED/N6rcxL9SzwWY3v
b7/1mEsh2xl7csrneutxT/toEKlARcmLF9WiqoxPQAHnYsrtvatPNaQ2O0rjq1tD
i26uEr+dtvE9St+UXiv8oeN+5ojHpN5MGu2xlIq655gJGhLePoV4Q6x+sPBDmSJa
tFo6pZqVt562MnRHhL4fk6wuOULWG5pzgQGHmR5ExzDE9JdnAu/Z8GUqEMIOw9QQ
G4YqXjSGr6pY4IcrALSj9uGPavoAoxMV4XKeMAPynspz2ou6p5MSICXybzg2XLcG
UiLki7bhiahDUPW427OKI3bJW8PyFPgVUKVsOeJ0oOaI8yDXrW1inBYAFb6RQrmS
6ct24oiyEhVuKL5QZ5XfK8GvjyqLmJdepnCkCiipdThB6502YOv8uyITk6YnvgUN
gcSw6eNQX/IA2847xPf74SgdfFG0lzrZpUVp2/ZxGUu5s3SUn2sPWRkOKY0jvUU5
MCxFtz6dvX8aWhKFar5B6dQw/lnr5mxIvhZBgwfb+v7D3HVDTgm8pDtmtSw+h3es
MKqv/9hdMgpd6IE8ptRUjOOI44QShk1sJQ6DgIBxF7h9tGjXAz/v98i9qdVzK4om
mIBQ1QS1tf+6s40YR5t2bgrfMLKjFTG6byOc8oC0zqdDk3pDcAKBAuM9OsEwQAEQ
EIP9PYxyEeKn+MG/ZHY2B7u+lMcfpuGzwKNDnD0KN35ebkcr1U4laSfv4U0lz7FZ
aI11iDBAwAnEDmoXLmd+DxMecBa5FX4xnUIZfYPzOZAhDgBmdRuiVD+2bU+HxLNJ
rOmOD/5eg/6sLWIQ2VbS+LrIvUvfzqgA2B42tFBHVoEzD33n5hwlGWji1KOZ6VB4
Zqb+YTQzUq6Ssk1tolmF+lYO9sScG2OhZk6cfUYLZSXzFf8zOIDsvtNFF5b58pkn
SWr4qE4X7QDvzS26NSNwMqkF3VVXCRfeaGi3CaylQYmFtf/RuS1M+U/g+I1j03pj
I40x27K2GSJbsLCzs/KUB2Nhq0I+WMSyoC5oQQpSU47aL/MGF44QNkkNNOxQLQjo
KGXMCi/4W6++8LCMn0Iz9wshC/nlCQIgs0856U3jCcrUdypC8s12QNLIqnqnyJRf
8PvgsDdhjj0OYrRAWdbbTTZCDFgWpQHt4ut/sxWMrYQIjsPODRjJeYMF0OgRzH9F
M60PggMxHq69jhMT82ZkLI4oK9wiRd1K/R7weENgacqB5M08BgX8kB3VKhmcX+tm
4QqFoKe4+E6rOzXh87MnolXzEyGR2oaqqWMFDWxp3wU5ouwJI5K8UHhNZQUfIAA7
b1CvqgrxyntiaWlcsWAigwLredVwlcO9R7sE2+fa09eE2tHAJ5srgRH/vOVYTlHO
GdaDlQlIYAbQkYbWH7bwgrGkeVw+ne0Tysn8LG3SjEgBHxNreQnrhycUQe/8QHRN
8x8pPhV+8DPSRRKZeAoJIuSPcyeJbR5ycqsFDJ504oWBjkPPrpY9obl4ox9S7tvy
KnfAKfDXQThLajRBAFfSGl2QQlZ/jZYtU9FjwrKnUc1N+ZrUQprkyER69n9gJkJ9
qm8QReg4N9QR9Smnk/rjzUCGS4jagnnnZFeq6utbiKDuCQmPzRCDlMp1WcWJYHjp
/5FuQktWeGQN2hctJ1Rtuyd5kTJxvdDHrjIqiGgaveECD2HRcKUV2QyHrnGrXujX
Dn5jIePi0Cjfx/9n7m0/Iux8Enw8QB7uEDMUQUA0UuvhdSCZu7MWkvIrM2j9PPwV
W0ALmzRf77tnXyDGlAgHSg0MLJAEYlxffZbHk7C/UFFNRoeQTEdmo2JsKOE+FhwL
upYG2UJ04DpAyoZ96NQoh1t+gnLR1DpKLM/Mgm+aTYeTHXSKsMaYRztAu29j87/p
lbi65Faj18Z01H4Iy6ojQr28gyaqxhgzuqDgSWvxyucotkcW3DfLPu/kVVACG0l2
oOSWVJfwYU/CoUdNfIdQvPy19e/S8ajGj2deBH5djSUCDkDh3r1sQ7VjwryYHUI2
MHYyiMjIuyt20yJBG1Ff9dU4RMB5akASwYNPWMsJZrE6MMh6vMvIsbl5YJJyhU8I
z6ubOlZXlbbTGQK8r6TGzA6tJucNOanMAIM/m/nuDgXtV/rFRIrsWDXUUiCtZFWT
JCStV+ccc1Md3/glPlzC7nYG8SVCNLdE5Yu6FGgBOqAK4PsYVnOLXf4RH9oHfX5g
27mrpsIugp23HBDGewTUf5FZjaI1Fm7W+UgrCeosq32s4JosoZ2gF8bNBSQJCDqU
LI50Zo+P3+/myJiJ0VgsZvNMe93Gwsp/CxY5FeI3wv36un8amiXo/1shR8P52lts
6QyiA7RjtcKa/L3pK9rI0u3KGzuh9eOXHIm/7vN2PCsYsx9dzVFq3EGNXPcH7vM1
w5RtZfV0zJKr1pR0JiFETDpeYhGLzcKutxayOVk+xYtLqMOBxyqlCz38uKcV6p+1
dzEWq3W8+urZ4rBxgeQqOeYMa9zP9Kr0WTAg50Lf1keF8ufhzKHGFXCj7YdRPkXC
kBCk8CGpuo0XEtgVPm9Xdshbq0N1F8xQpUQIwBD93xyBoUHNh7lW4Fc+WsK677gn
BdV602+9q2Z5wFmZDhAQyLzH2FB9fo+RG52sG1YgMjo7u8u+97fyTiLWExFGvjuy
ZYP5pZzR8/lvz752F0B+gl3oIhoO5Hm1uw6uQC5fodEzbmOM9ZfeppfjLD7HZc1j
b4HU00vHa1ZwGwlPApQb5AcqhL2S33hmp2UOBuibL2laEuKqco3p83BnfEhULcF1
ltErr3Qg6kFxfWHZ249yhKLQbmc4OZbdeHsA+M/2GwXteQtHE86vxdMIkYjEuyFq
LCoOxiRjmg4ven4DzcaW3m5cQMF9YjfdvlYOJ+/No6jpIxF3gIAQmt+g3BDsqkSH
fhid46rLC/Zo2bM+uxUyxhIRq8nsWANWen+wCp6Y30bx6KaAa64Wrpdwqyek39KC
68EiIrKpN/CAyNxU7npO9sRYahfFEnTNRaCTmER0gzOUQPVptDeCp3PO+Wkg9qN7
0Ad3FnVGE9gDqQAHA8FiPJCXeGRf7vaqqREBW/3j2H6RwIZC/ZRcXWjVR6KJ57s2
XQjxGSsdMeETBynaHBkqT6XQdYZ+AY+0fDD4/DaDRv9aiL6mpj2SFraRmTFt9ZEi
Ec/TbH+WjaUOKLIHvpM0bbwX6F5t/NKSvKgR/TDtwoLqVae4XvFTU2e+duNk9Rkf
/JilbP/bhf9tJmjOZ6leDOFvEJ9sxR0v8uCu1fVxowYgSujZDI9y3ptLn4LmK1An
MzlvMIDBn6qqjy6Qv6U3aOObq9ADA0sxH/XCfjV7WgxuP4xiCBxUxI2J1fUQ1lVj
3jApNtrv2KWr1C9/C6Ry9eNhnk+22EBsmoxaPzg5LJ8d+wkKAKjzfDR5k31V49Ok
w6RYQC5FgRdcjgJSbfmbDMlZu0I4eJT1bqHgz+VCOnBxRcI0lvSR8oO1ntR+Wq2G
0jP2kkG41ZpOdloHLfpwU787cdRrJOr7xzWlZhUZcfYZ6s1PhuXCjM9eoeSbq21y
qQCICwAJxlBQM1AiJIPtK0Cn2AvCk6r08Ox2hxOLq356gSlfKIBwecCMlrWBDgRy
jMthNjCv9T0JE/NdmlsSbRctK0Kxx4ReytqZjz96Tc/1UXwTJY4nXevcXHqEJBP8
+JmDosToRN3p2lzp/ZeMRp/qUX5Sw0vkO7X6Hb5N/ZRvgjd3wHh4lUVBjvmsWeo7
3zmDX5BVO+086jzlTkW40vKO7JcWjDUWCMQ79uzVV0KuVtb6l4QDrcrFtS2HG6MN
sB4peeYwmSboWKr3k39oemnG3TlR2XInKddKW4ERGRU5ldz/LJg4VAZwxOnuMidO
r5Z7D93rTXIzktylSoeiq0ktizDN0hZVqRT/HWN5boOegCBXNM3APOnlhCw71xqB
KFfOMcoQM3XxuNG4UMs+jnu4j/lhMVAzi+zQkCNrqHOFl7GD7oPDopM9S/egSIac
+64BotfoRGSoRkYQg3kNPszCXywJvWsor7/tyEPsamA7O5vNzTHFpMq6/HKKrqZN
cGg0hSy00Roc+vVilVAlId1gRRWrj9VnAgxHGeM0h29zMPjEbQyKzaCdEbOKjihV
nRy5EKx553hw0559jquuFI/yZJwmbM7Gnb36154Ruj9PLwG9tzCEPGIpVfKcwiOF
a+fkZKyzihJKHxKYr11DJi97BnPiLj/mojEiI7nIYLh1AgH9gx7GehviNdWCdkm4
WXcat9PZTzO4uQlzPnL+pgVtl9nIOdCCYdziCNnmF1Eg5oyV3z8yTFq1C7vsmumE
q57lED2s2KEHPQXK86Bw4PUhHloCj2Vuy2E+J64t2yf24DBWfm1+kudUAMvX1441
FSYBcgsIGpPagRTWk+es0XJwNfV3ipUtKvIBzBmoBlRiRRoprAAVhqG4UyJsqH1m
79o81tmQDdKC5zYeQaE4rkK0gfsvlJTt5XyYXIxTj86FIBnfMdFZFysGCFFXlSB8
j08/rjc2nL2rzri7Vqc0PJX8Lgg/kg0uPLhAVyB9FcXSabCVprT0UTWwQcC9wOBH
QCAUyHePmMgTMsXELJ6u8SDse+kmOBxRMsSYB8So1cKqSi6I0BZsRK2iB2O9QRBj
tEHeso9dSv8YYbl6Im2fY9EQwzmZsg+5Ss1938xDFE51xYcokMA4E6CZizwfciFE
ZL59OcLZuHewFHpICj8GDSvYOrpCtNLQFa4UON6wmQQvLKSVa+pkkSb616/Pm3gt
7UVT42YxzWzXJE2PC8zth/DBM30Pphuk5ahqUwxn0secW9W9AISC9plZ+lAOQj7+
cv6Wns08vhuc3V1nkFove4gpOxz2jjlUUydGEyhsFf63AAHQl1VNj3eONt1GdsFu
rci1BYD56imxBDWi249stLlNdYcBbMdFI4ga9i6aadAmJM2pKMa6lPm7xzBfzf1+
ghwJmO4OrWfTldVbquIRQV7uFEe/PvUzYVj0cr5/mEwtqK8FRHkuZdUoNejfXobZ
YXhUnH4paM0BQWbPV9/itP7XcTmit5ioiZ281Gl6YHUkLUkvu04/rLN/VkTOX7ZK
DhFTeMygKXBVhmzFqP0U3v7szzywrDAaV/eUZ9P0PIA78sGfaepgDbHBMxEkcQJd
kzkk5yTdr13aMnZLgNkU2gYUm+AdbqCL1XcNY7o/SDdFEj1lh/gURcYofwxDthQ9
meaj77dOjjjv3VumoEGsr6aKbzAc1PEp4TR11yJaTWPpnMoQkHywgd1gNZ8Q+rCm
nfPdCcQUoXj53fRb6Fds4vIaKWFJRiVG/0HOkCh7TgOZPuhA2FG1U6pL2nudTG8y
Kbwd6coXhVWROUO+Y3Wrg7/eBZXfHvL9KzWwhMDUbhA=
`protect END_PROTECTED
