`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveFeL5AyiB3cfGNPW4ijOdUVd8UMSbZhmoAGT7ylTKYF+
5i3W4n35cYOnvFCurDAowQ2KstUaDHFsB5gNYDnV+WjU5NoBcWJmInr4GLO5dejU
YxUD9BkXA53A04q0QFcH3UctE/9SrAw0FOeD5BxtlxiBNSKi8dxeAHUAV+5hZC4z
PJZivy9gE5TqeQMq7S5S4+iQWcs6oiHCGY5FA+GLPI//uHPcEXPz+FqrXGXvdl+R
ltE2y/n44XE5OggS/1pAfIQHSIfjc4UTc1yjZ+zerHd/cBHEwWdkwMraGbiPGfdJ
ZFOhZN4n8qp1eW7U6uswIcoubnFHCSVbD/N3vt5dQYCQcUAhC2lJSx3J8Ph8qAkB
ML2ORA0lM+MBqF+ogv4y6//slo4zR0obK8dxhH9RN0xmxkvvEz6cQj+WlpBwgqqg
vocm44Yq30bz0EOJpxjKhU6Oq/H2zM/+guX8xBFbL8JJYUfFGqog/Zb/ohj1qxQP
Mehj3QDVGpqmB2bjV0rZ+5XAEIbOoh5r5w/X2FLjhgOgtZLO2XA8tHwHh2b5y5K7
`protect END_PROTECTED
