`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveOMXVotO2aXISZAZeOZKUWAv17SVA28xGVcgfL8zw5Bl
MlhXrNEVYZvhNBP9CUybEyOLjA7eT0W4Ro8j1RUF8bbrDRrJIReRfsHrKXDBaZn1
IMDe8FW+tSWvZ9/71YBF7KHUU0QOTETB7GywxwOHVuYXjek31FsSsYcSRadIUV18
M73vKzQbQDGefJisU8LyhfL2zcNphNLYQcmzj8Nn2Rlimdpl0mcKj2ffoNV6EvkB
NhOYaF3qCjNu3wdeQT8J9M0QzytV8H5Kp/uRXCcOk2vHD8wVCKvU6vSduGjroQP+
60RDUallJNRzi5by6hyj3RIg4CRWxU838ar6vwIK0xzy0pHNjmz9kvIdePopG1i9
s7qZB/noEtpSwcNDQI/nmeHVmqrtYERtfIK/UdMz8xCLmPcTYbeFduJi/zNgoNCD
uQNulD2lG3gf/lwM6xtLgce3yygbOmWVHAhnxWnA3HtbZy++YYQtmh8I5qd398mA
949SShVlBSJgiy2jcnfYMdUfkBazwIDGcnRpW3n8vteSLQeGhhd7BVr0E/qNzUyu
`protect END_PROTECTED
