`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
n2XR1WeM0JR7NmOlJGcqsjS7JwKbid1W1cXIX383AkLhIcwRfc7GuBrCu/mOi35A
Lj+tLoAQ3b4TpdJ+79a0RcPvRTPjJxYmFzlg6A76kr06kOhxN/5485S+Da7LD3Ml
eXB3heL/4gv4TJjPLUPwjj7QYnFTRexZR4xcc0S8dNE=
`protect END_PROTECTED
