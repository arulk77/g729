`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu407eRoPjFsS1rjdFfPLr7POPEfHVcOJ6MSE1ppmSxnTp
E5Uyw3aIs1FvrHZi1VUafqOZtKZlE0cMpP2kSQkcr86E6aEYzjX1/AZbdoHc1e1a
Pj90gARgTvwJzEVQmJfkmcjLvvUF+rQn3k3mb7QnuQkpb5q9Wz3tq/sklxQntxoB
HLGJwHeEYmV3SjN9uBZk3bjnGIzppWtM0EAsdmv81eE=
`protect END_PROTECTED
