`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
j8iS7ep3YhMNgW2xFkXmNwDNPeMUPL2F9nwaffI1gMfFiTcfhvVIurTtI0q6BHpB
ctBVWtUodZ0SNxMDSV2Nuu96SyrZY6Se5DeZqyUe7qD5BY6v6bZtvxvAhr/OOpp8
lf5h1mvMPITHf1RvghnfcX/zCYbkWLmqqvqVIaqmz4PxlX4reOEGCnLHHBvsaRwf
kWz14RcPC+VWVzOVTaebX4flZK1tlPuWR4rj1PFO1hxnI+1XgFI0JuaBU/PK4am+
ATIDQ/OXM794SBrV00ACamPbauhhKYwqH489Tq+DOcQkAm/YyU+0HokhKJ7kgvav
MJchiWGsAKJ5fg8iddo03onZaQjewMycqKfGAwu9vOLto+2CzYBdnmAfwhrlKKrh
3TgTDUaK5b8sFh/mtYmXCcEPn+q9f26ymPRTHiM7zOmzCeIws/9qnVm+FokdGTJ5
TSmIdzVsaNgWNYrftl6DqQ1zsV40vCZq5w56Xzyo58dUX3/1i4ZWr+y/DpaKWmUw
saTgTScZfT6KzKj502yASfjBx7mwMpVbzsc72rNK8w7a3GKS/K16VKKECKMxZeCH
kpbKduZE78VK6ZBfN5UnG7JwD62cHhjeyE4sFoYHqb3DZt0pHBQuamLlVlIyp3gz
eGKeJMByV7rtSwY/x3GaiCEb0eyb78+SYhek4RrhMyw6O6sf8CNnZoDnzRSt0Mxw
Kg56FxyhD00j4AE54+34VwREG9b01+3NKfH7wHMCsfDRfBJUjvOTSjiwBuznDN2F
XkVcIyYlWPwvFMGWBhdilK7rFDHPe5yRfpejCBuF7vzF0KFH7x9KKtPn8a3lN1pQ
sIosQf6gT7shFyxjL8BdgK9mhqr3z46b2AsKh3p/DTKsh7VYhLeKR+cxds27gwWv
5cV44q/gNQTb8ME0nrtYgQ==
`protect END_PROTECTED
