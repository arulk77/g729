`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveL8Ie9inRUsUxV5QlvomqXVPNPMcgyIARYC7vBN2boEW
O5PMgO2uChqkPD4ZQcABCSygy5ZWLX27UclJ79nixj+bN/NPL0MCjkyXcU+26MkU
RmQHW52ErdWpwxrwy3xXMAolmv8m0v/1uxoyJ7aKAaRCIRWEcc9+EeJHtCguqBsM
Jwjpmj35G3qu2dN+cm58//MLMZXy/3lGERZ6ASSf27d+7R0L7Ub60abDZPrdgkXa
OkHkbu5s5Wu70D2MraCFgHWV5JI4wZLAfZnuor4EyKA8Rr3D1FdGD7BHx02TEJRt
HW3MqCVaahob/LzPyf/tcD2M4yXBmN83yAaRW9pFw+rGxLXRWboDZFjwv703hKM6
WYLztSjgwTNIAc36OFEsZdv/bu/dr9CilGZiEzk+Kl8CfoNPkJG+wThBo08vkIbq
0gH5cOSz2Rf5NrgIXj1bMhCUAZp8+cK1/qhDqXmqZuQRmYvv6eGIWEcTIytTOi6v
yzZvazMDO6uUgTJAsyE+5hRPovCOIQAAWvTrDb9qivKq3gCbsWEwkb5RxP1PlBAp
3cW17vSunJG/vbLzipC893DvDewrh0mrYFrKwz1v2FK65q+0EcO0Rte0oXioYpzD
5G/nk+0hBrw1sguRR3wtY4HTVmaFkLuykMPsZuAiAzzNk8u8bgXK+Hq9tkKhJpp/
zKAKpAxQz7I6fhnkIis+ZYS93Zhy9TAotFZBXCDhubzFytn9e0j8qtcOhdIirdT7
SdqkxKIZgUtGB7b43SWiBRgzUqrjondIFOlsvO888qUS8V7lXV2xJ5+lwrKBu48Y
TE0HvD+O2COle7sSzuDBDLIMLK4I7rHIV3bajQ6eyaA=
`protect END_PROTECTED
