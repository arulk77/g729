`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu46UP8nedz6CVoghghuxM2Tg94nFOUKUhH8YBOcC5CTKO
Tsu2K1HdAhfQ3JjnCPsOaDWyJMqA9IVS3MLcNWjXm/Hq7SOHa7WcVVN+zeZDP2AM
JgVYkDs/MrnHNUBwjtKCbPzLw3orX+5VjNGvEoqlnb62N6NFjOVGSgrupeS6hlrC
ydP08FH5ueX60hCiPyxmT1L5r1miJcKawC0pR1HhLz46dCXPxhjq/v5Y6wBrxdwg
rA9xZYGopyPUC97e7hh/W7NVV14HZgjJhmMK+ob3y1s=
`protect END_PROTECTED
