`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKK7p1/+gyw593y/ALzemhnmtGc2c1cOfBREDEkuQ12I
JUUqOJEggJluAJlgvPU3m6ZI/Bncvac3hw+N44vSjy1Tq7E6zxsR09Zi3HpTVyeF
PbWrkkjc+KRio0abOisxGfTpGl5J+SDYBCIkfuKEq64JrLr722Htw/p3F0pyZMIT
PyjL5I4QoxI6yTT/X2MC8Ziqj6tK1GZ5D8DM0bkSYh4Xmm9snyPoXa6l+Laz3d4/
mxMjbS+ryg4ENjOaIv35CA==
`protect END_PROTECTED
