`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu43rCCIIlmdzKzJpu/VGRuNs4Iey+VYuZPwOrqAW8ZCgu
jy0TDJKLo3hjaSW4CEBsbCsuj+JQryRCBGpvhPPlWUdNpyO4RwhN4Nuly5hcqdab
ufLAMaVE7Q809Nddl3D+rWMhIOSnBdwA6525D787uuGSX+tADFSZFTdHGCbQ6LIe
v6OaMLcYCnSoGZ3HZ1cMJ/XqRMEUvh315EW2GI8MPZmGszmFnPhst2pvmYYGmi50
qlJegP+KimMBFbOqDdON8YJgrwxh2/6zDXKPu0Qx4iQ=
`protect END_PROTECTED
