`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
W52by5FksJUdhgHLv4Ym9EeLJZqBUWYIusi8JNneApxDQ9MpFmXhDstzsCMHJGY+
k+AWgYZehERBffJqSZwCKTq/DtE/7xOLKFrPdF7j0BNvi0DMOawdI4/m3m/45o0x
c9nAoLmJzldBzpNI6i0FPTfIgd1gN6eFdi/v4m0N5S33CZXAtDRJs1Hh0eDJeIPf
YpHYIO5BydAXBwA5nNmOrBbh6tXYimAqTLIYRvIhWfLb88TMkCFfov8C0mYvJ8S/
l1t8ov505WGHr8LBeD5U6PbMgL0UpPQRVC8sR2HNCHjzxda2d1gbd0tWyUpH8+St
jc5XOGFZG4RddBVbcooIbwqbTYn2csgJt9kh6qRQQp7qspi83NQwUBcek6C9OTlD
16kT3AEkUdcXgEk5qZhBebQalS1fF5Sldkqc0EFyyq97/Y4aOHbri1t1MeqjKDLs
ofc4bWGaVRlw5jN7uuzHjNhlJj92wPahA2F4SgXB2RI=
`protect END_PROTECTED
