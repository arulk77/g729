`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveGF5B6P1f+9FiSQ9D36TNnPnB1qNP8sMGAhQZa0/X37/
OPDJLmDsVoMRXfFytAbvpwDwZEtSqbwrPsT+E257Pjz4Q01j8WjUIE0seiqIsc6v
gVzQTx1DMrFVn/t+B/4uQtxjLHGkMhK4vP7NzEGO14CBHcyPAgs6Nw6T+2t3QwmI
I+LChxc/TFwBnkHCiCl4vc0xxsgRR4EQTSotpwPMYzhafCTuHWC9C/q9yA+UUKRt
RCcAOrs4Sp3eYWh63khlj5sFTRJ7DvQ7CVtr7k1UxobghGCJox6tanYhoe9kcpm1
vr44D1cJS/WseCxYa85KSA==
`protect END_PROTECTED
