`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu40qitP5ZgAvz8Jnw/4yx8To7bo02AqdtvDfyvQwLbdTq
fe3VwYRwg5oPhOLao4MXiwY6QjBK3uc513kT3UH1WKSwfQOpE8rw9m+pM3wjBMeN
o9C/4m0yRY8rcIeh7COJzajt2kKIwbrnRKSb4zwwv9W8XTJJMI04gc/9Vm7fWq0r
y6dRrfGmc7pg4I10WzUiUQ==
`protect END_PROTECTED
