`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
3uYF0P4SWdT1PnMAouh1abznU1niaoN2JYEr7DDD4Ups3eAPHb7dRLnDfsZ2a7nT
1Y5KxiaCpwn8DkNG1av+WIHHqNPMIFQMbDZwLmebnSP9bfbUUYVZ+M+pOTa9+KWE
VtvGTBGhSKBS6EjDJopq7DVit772CVSOzQjvuaEPlnpRXPxAOZKkfyEZJJ+hV8N0
E7YPCqSx6sRGyxUWon6ci4JT4nI6P3XoSNtuEmjgWrH497S+7dfJ1s7Hj+124zo9
G3IKO59Xg3oe6nPyeABp1qaX2Y2n4Ha0YI/D/kpTcWLZF5dM11ou9sk45ZOEOa25
FTWftXkGIUoOEY+lrRSSLLbI1CQlBqLNF5NkD8zHojBC2l8L3aVgJhqb9kR2j7wf
BMU/Qt6QPgVaVBwYFlgC4Q==
`protect END_PROTECTED
