`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
mlFBzCyNIVABC0bhYTMiK9reQldBzvd6OAR09mjaZUdk7+aZGQL5XPz2/I7/d8/p
PzQzJvgV3VZoQe2b8HNh5DVVnUEeQTdLW8nH09DeqJC57W9kYbuMOSPBg7S2/HS1
FKw+iYleg7vRR5eyWw3kQfwnwgH5ctx0BZlYq7OKCOe9Q2svNExltOXj2TTpnVY2
q1utWOrhVafid7ikHnK4jA==
`protect END_PROTECTED
