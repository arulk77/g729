`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4/k1/INKInIcM3Of8OoYJud6skXIwIRqN9p1Q148o0Lm
hrHqKjoTtU6ix+FK3rCZRFGR+sXIxUsd3eJOdi9Mv8zDooCNoY+4gwN/0TEo2jYt
uBhd2aBR0zlTK3ljGj8ZyQOIVq2y2725OmMcp3xz3yeRwxEcGaSbbPwqk3uNF59c
D434o8EA30rVscYedwz9QaSjxnCeF+vFxCxa5BYAb2wxVHIoYoo7AGYfdThZqbhK
KcR8QZg+iPQyUdrVWPc+U5zIcVbS+vIvGc4j1OLH3BpdkSSloQRo0KF2Of5nnPKF
Qomu9Zbi/eGQxX59FLfaWQ==
`protect END_PROTECTED
