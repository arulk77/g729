`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveG6tnZXYQKKnXD3NpwBbDojy7gt7x9Q0e7OW+BDgXjqa
FCjt0VsdlhMvhkwwQc70nR5LA33hDcZOM14u8RdEKLto8A/o/damA29plJQE/4zc
eGmtVUkIww95UjgrIIiRAcj58Lp+dWRFvQOlE2GPx3Z+aMdiTnLy41EuiMxF/DWv
CMiTG17a2ZZA0lZFeUTz70d7WJao/5kzAuEmtHf7hY6eUCXURuXCyzBquFRfl9vI
SBaOm4wNmhRxMvUTRC4JMhz//+w3ynCsSTaLYE9eUnlTeVgieXGMm6cKTlUW/b5S
JM1ugAZ+zv4E6Gtm/y9fcGa8KN2TOTEo70LjArWfZoDyy2+nGm2Lgd3F5u6VGO/p
lh+cxaCJdpTwuiwMXmkCzfZNUhPY9UKka0DuZIh7EbTpL6Bb9h6kwWLuDRpxVpuI
gpegveKhcLeKtT3I9DHL6JV5qLL3f2h/M31vlBiiI25G5fgILjl03mLEioQe8gbb
Vot+WNVwmSfJiTMPZHaftlv1iEPteY11dkPdsKg5hW0XUH6q/VufmiSef1VwI60S
5Y4cKiMuG5MspiZWaRxzmSFJUeU29Y7gNCDzLHF+ckTTpjWVfQfFLcIHLJxn9rLh
gp8d/2XOqHYd7XHpctRCySM4FyM3QQJJ2dCRz6e3F1LpvqYMi1/KLK1koZ/mx54+
YIlkcnn2vEproZ16AG2YCq5sC6zDKJb4Rz96upTcx9N/BTgfW9OmdUALyxgELZpd
0qPHqQbjzDeeBHXTkDIWVGNCriA+Ah8HvHglAZw5Z1kFgMrC6aiIw2hm9p4Rp8Wu
NYDTzvnSODgGesxtWvjVqGiwtOLu242H4ZKDXQMtmbEJqNgEMcAmC1mLxC7F5wI0
/C0phD7UT/FA6N+gMNt1xFyiUdgBTJrx5yHMi++vjZGhu/j170piygyPNA05JK/O
j/82rcJkFwSDXK5OlNlbe+AALDzEMSKqMGzLqRurvsIcTLt60+yC0vbOBwMhRFHC
VW/miknAWP5bc87pA7ZtAefX5ZMk278K0lc8hY2rAjKzdAQCD2LLyOKzVucGNfhG
+lvF9Es+3VCG/XJQw/1SqjoiCbG32ytCM56ueJRYXpc5qIhLHkNeJ7UxjEz08u95
lyu5gRGoxZysFFnXTpdn5dQOosW0bBp6sYLzFePEnjnNzbc/2qrh3Vv3c0L//ujc
RhCIhfAcnLtjJhLdkuCwSj5/80RHN3SBAKpmtG6YxZ1M12HiAtkwmNvIg+GWKMBW
NGJMnTVLU4HAUz6GT9RYS9zyFbW0UenAgk8ekij85c0aCKosddHwMpU82n94xec0
XODH/vPU5WILF5YFyGvov5dE62obVIt3qLee4R0UvUe4oDX7BcbyydPxib0eUDXU
ERZzBNwcTvwkd80GHeFCfIAKn+jTeRqvffDO5hU7P9UItzIISIXRfT6Yw9zUK/bP
z92GIp2o60k5UF9DeAPlCSdTkyM8/Pxlnnnz0SGq+nq1ubjtrLEgMgtGyYmW9JL5
vqF2PvAdXWSiOocsL8GJqB1io/JTmrXGzNy0NnyCwRGCauo2hvLFqt2E4Slt+7n6
2zvPntDyntI34R4P2zO8CYzJG6RCgyBBx/pcwTS7xGlWegaeFufdaWyJrTKR9HHJ
+O+MKdQz9wiAN+3Qf7FXnw65GK2XEIh8ubkOYTFV9WNr9nTVTJS8en01sVEM1Ca/
9PDbvVzHd7Gtit9OI7gIRYkpEqG5KOmUGReEkG5S467llbZ3PHD1bIaoIKUX19fU
tos6i3gqcQrJ1PJ7sfNvlMYR4CviZFvMj5koQ5/Kfrih78y9G6Jg0+hygaY0nF0c
EqxwJmH/riamlK6BmOv1JOqJeMKsWJyhB7LUd9118h6Znvk2jV946gkna+u6k1+h
kxpc6ZRjmzknWJBQf6vQ4j2S5iqCEbRcRB9tIGQbx1mS3yHZgW0Z2ES4WK9sM2Pp
hHpqp3WiXaHW0C3Ojxnch80wO/Q5S2xHujkKKLdZbVQrUALeMScX0nCXz1n4Tyyk
0dku8Tc72gX5AFYaJh/SwYSjVN46j81W3fIpFqGC79IrTz/2IO6jgVmXtmBLvxAD
T8s/tA+M7pkAq3mlDT4sXywBmvsWFG6o1Wp5bz8Ea/KVv2WECqkut3AKOrm+6H8A
YeNFz974xWut+Dy9IuZV/uEyakhInTts4whUz80af1Y1FzunudmEIcex4ofLFEdZ
HPOQ7mkU7pInqL+sPB+0SG8cFtkcej/9vDvmAu8GlopnplNUFzDB0/zWs8qsNpxZ
NZ9iXld+bOdBanSXF2x1d/CKmks87eY4+Lpc5K/Jm2FusE3gEYnesXt6nPJ2IwNr
HT+MUTHb7pneeCUD+H2ItHh79VYEgrwXU7e04KjIpwuBqzUqmOCygC+Z+xv6Btz2
MJ7keOLDxj1/xQ5OVwHguXgKuw0YvmqMcqhrFrkxsNhdQGtWoSTKoSJeUa41MmYo
HvE9t+PYBeuE0wlA064NGAQLkw4WznVyScEfiWfbcZOd8ggdMHX2SUriecwZfzRs
Ydby4Uc8LLeU7THOPcSES9a6TfI8weFe5vBBfLnUDuqUNEVPNhFQOz5GQ7pOQ5VJ
q9wATa2daPkySk6fdTAKvvkm6cgSCsOnuiaJFhgmfHUje5Cl+xuuU5NK0SHP2ewi
YP6fFBUtX2SfJIDY7XHPWGXbxppNuV1jljIA7FJXCka/Ey7+0NcT5ASxUtVDQ46s
NtxR6zJvgcST8azBSSpHGzfxxUwziIpYw+VZCaMiKSRpRz73Cz0sugUQx1rFvfic
Fz1yoMuD8wm/0nYzsuG5p8Y+i90jU+4MhZnRjJDPjQvyc90lMuFdJXxX5RJGTq01
4R2PvVDnnXWO+OT7EON2C77IA90JktfijIvLwK+GlqrvKPIio/uBtVa2brmLDNEO
LdW+DeowFZoD0uyTy/tDcwWTT7APiAiJ6lL882QdkBHFzKf+O39egByZe6wQQ25M
V6ojicPkpUqQawv+nALu8H1K5JSW6HX0QKOS+yTGrkp56fr5NXQTFrg+SNkZ6pgd
SJn2QOh2fZFYnwGxLCmSPNYi55imPgFHkcFQImZ4oAP7azC4CZNhPlu1Xxpod1sf
A8e44Wifg2KBbBDphdV7CH8iPlvsCD1tgQkfII2KuE7vgTYOF7PBYbfcRWmVI35q
Y+XQ0gBQn1XW6bVwLf/2THqHa1VZPrNyJJ5R7r9HcfOidX6rb3kptLc0PLDtA4n1
VQfjNK2A25lGWqF/QxhyaAv4gilwdRHWR7qMD7FYZqFbRXDQZ2DQdQteKP15OOyc
koLC7OcD9+G/TUPS5B3mLVUXUrcTDvCJfXJgK2XM1GeapaF7GJKFXg5EEYdKsrEO
DpiT3GHbNmae0woohz+fGuP6kIez+0I3S7gLsn291w3kS6JCtDs98Mpg7R7SbeNG
8xlcFpHjbzVUJUdqPr5hTSiKHUh8jnB6ECTfRPUIuInxYimfZ9PLQF/cFXcYFLCN
ioJsIt5UwLEHIqEKl1v5wog90JDdd2GlFMnymLjgqkCI+MS4yzEwgCwPJFOXtQMu
o1a79BBAWrsQ/5f0Ew5v/QQB70pfabFE4psBCcZE53Bx0wxgE8Ql0RSz/+7FtXuB
1BhGUwEELRqSsy6ofgeCuB3QkxL0UNKgi6L66txmRUoucgtpMHsBV5bCWO2UupVy
YE8vrexwZtrwC61CrYl3lOrh+YQ6msaHhiUAzubD5/m5NsIa9FmQ1Sh8hecEwwL5
hWc6fAvgfJYCkrDT0ogZLtACrBH/3dXp17f6D5G0BLjuL7oxpl5ZGoxQBraMLXXW
u1TvxpQQYRhiVMrARqdeDUsG9y9tVr3CH8A1JYsdfmX4CVnoz4EqJyDvoW8fxlrm
yxLL7OkOA/GYFoEPVQsUJIpmfAoPd8U9vQrJw+by7z64fM6wigqnDqYvDHEInWBu
mJiViIgdSJRmV4pmzwe+MvcnHrxfI9a5dKx4nXDmCaNmgqcO6DNdtvmAbJkK188q
IFODDPfmkQElU74XEUKbfY+gz28tE4/pmoDbLtPCuOzVXocYJkGRe4P2Eo0Un01E
h/ZdQfECmNZrL2lEpJOnkC6L1DNXHvxjK+83PlabIgJh0VTRB5jFP8pbf8AER/UK
fgTGVY+jD/AAA0FCHBovoJLm7JPCWoDTGSWI9bzMKv7tKPT4p2LaCliObpqC+CvX
wwAbeGPeZKNzjfnB3McWPjqW8cRI8i32288lyzeqpZ7ZhdeQ3nZ9DxIQDw1nglMD
j9stvWy9zwVPSSa2Pq7flSKzk+GbqxUMmm7TBXzbiF7FFkzU4ivWAyBBm41HbiTP
rLrHg0O3LpABRMmbXs6Ubl3QpZLSsSv1SKX/OVx7+3hff14xOd0AF+2qAnirOdUd
Ys6AYj7ONmTNNGA/7rgXAvYzQiI6y6qzqj2gExmRCFs8aveQw4h6xaMghDmMTrQt
wdaafjFxMl7JQWHPe7zZ9A8YxmHurynaab2bkO11Cr/DXvjBb2JrMaFhxJbjGR4k
N7ohNsUqGfx5mKtQOYojfkdaWhqvUIzBC81t3ksc9BB0B0US+moWnS7jthIh2bXw
7d/7OK6E2tqW4Kc7x3EKtds4dBGbIT2qDzN/JcVF4uCsUlY56lua9rMelfYkpzdR
J4AFo3a0U7rXiatO343VE5+rwyzYt78Yx/oG9PgcrAVAkFpGrjqBQ7YcRBiXaHvI
OwG2KMEhTV/gz2bCCP9diHhNWC3/c36MSx28HAwebG8pGy8eqsUSnEY99YQHnG3Z
W2v0VB8EPrjckhyau9qby9qr6GdD5o0c27Ub3WEUqMSsqTKZbVzqY+JH4dRjUEPV
P2phEwRfbqfzWpZ2wZZ7nJtcfIkSLgUvkvMt7z9dxCbuUBzDfNnP0pVbZ8Cn/wLe
q7RNVfNQ3S3YQ7qIArk5QSO8EEeqEE8m2+6HoIuMYLoq3nIOrETRrXtAaHEtcijC
CC714BS+R89Vb/3MYkcrBmQi7B7xjREACtEZ/zl2VO+KIpFM/57cxa/fJgdbez3T
wS2iK+7lAV9I9+g49hqHDKGQQBQVEmRJy0dUaHt5+Pqqk2AWshN8BfrMwv1LU/2A
Ib2QZWsiF98zgOP3IKhMIny8h4fNa/T8sXwGzi54do/YAiZKnX+BpeSGu0gUZ9hE
0K3Hm5M6sMyYoCzorG/qy7Unmdz1ILKZTJ0w6zrG32/k9YE43JZKE7ZqSBlFob8Q
O73dB+pl0muxXqPmt9KNaYtykC07XxsImlOaDcev5POJjHx8sZl5p7KmFV2FOKBW
NMgyxL8XhszbcGSn9FoXH3YAyXU2bvGLAvz0CD6h8cmsv8MGwxPPBk9HeC0POCWJ
tTXyheGF4FTVWtSAyKpApxFdqLYlSh8gx/GpT6ePcKkQAUjrAmUMatOICAQQdLK7
1dU6k0aUYiNHJ/1FaO8CqMWuIPTPy7U4Sq8U9+bZZUnUdIkecjpYzc6l5EEqe22d
C/jfGtmTUwt1vY4GAsnmeN6NN77YMnOHDu9mfZqCpenQjjJxLcWTACo2OB/8cDar
iTAj8y14sNH78XEFzcaXiS/ZaM69QahaRHQMKV11zwx67s/K83K1K/FcduJcuCQU
dXu+8+mzLoWaeDLnZh9SEkncrU57jMSMmN1F86gUTa1pChBT88hZ5R/+3Hs60hSm
mgZbXYGPLYC+Jf0IVD6MYK6OmWfZHQ4WyaytoRxz64+z51W6gLy5/QLeCZHI8HWi
SU+Q3Yw6peV67/YtMrhCk2zkNNiX6dRMv6v8Pun96EvufSE6fGVIobp0KOWPOFbf
vnv7hMKjmjniNHsmIDZaiufu1Ep1CQldnxb57AlCx+TwgidbzXjCVDNm7QSLNPcY
FNbd3PbOR5dwGJ6fXlMHP+8mCa+qqU/8dVGQjw33nFth1FdBwwbBtDjlFevBBaWS
Oclq1dF+yxbFDVOAdlgUzdUctW4VRBxMhzqaXCCtkn2usDjYqjZGMFMnd/N4YUZS
zX8uvAk8CBEB2cGe69yFrxfOHcFpBAU5oR+Cp3hJHhzYLsfg7Re9LGrtJwBbLSYf
IupU2CFkYrBrBsdbuDJpz7AI0ZgfeayfZSdT2EDQkKBeeJRouBFvii8SV8oBOyEU
Vj+gLxxDn5N/3gvsYYF1hAoROu1ExL6Q8pGFj49tisEblOp/oh3pNmAuXVLHqvpl
dmdal9xf4xWY4HIdSpg+L8d1fkIQOjvvOMgWGEQPf6Z2pvIqh6VlCBvST2kBsXZL
1vLBT2QlkEJSTCyvQHz+xbS2E9LGBHdc4iYwVcOMnA+00Ybf3kT7MFdYUtYSUNh+
4lEdXY6j7//DYuobE9RAFvbFn9V2Mdk1ba8Enix9dx72pbaoAWIFGf6Lz+bHxmrR
bowjEFJONZQg+HGdfD/gxUwyKPt4XfWNmeoSOZrX4xQjuzy/PwrEYcMj50PRdoET
yXRm4iLYj/+n9iYi6LWUVV+eVBEfXtCvrksyQQN5+4N61c5Leo9Xmq3fz20Nj6Pn
J8kT0r6F0PU4so1yehhE/dCjluttsOWUjM9nDJGu8NGODCV78LKBPJLaC6jmCgoZ
iu3nQ/+Nf1BQSgmTgTq6FAwR9YI26+CPqAeLGlfvHnjwEaQn5s5nRkZa/riTvy47
/63VsCxDu/8tGHWjvU5PjaxrQcCNt/3716ems2k8LPbs82QsEgI8p1mURfyLaOOd
vSFGdMvcf+NyuWXvoGXbURVf7fcZKehmKQB57r65LdP56GZv2b6Nz8J3I6MJp390
Hu3e6AyK9g/rLdV4/u3tafBl1AxUwpgguhPJ3pVV0cM5mAYZ3B+mrOgshom5lIdD
5kyv0cPJsjkyqk3o1QvIhjHhEvikpktGLlUvPu+FiMFtC+SXjAcdW6DxUwCeFOIf
iqsTEQ5W72PNUCYjyV1Rhq0UwlSpE3SfEWEAmakmzX6TZvvFrXofJKC7t2L6anHd
JTqKYPQ9ATfGtZJiaNWvV84CwnPW92g1dn0ZE3CDb6TFKPoLZYGiCmqcmqiu/2Rc
xW8jFppjKShFHP0FedAxwCl0mDv5OlCZIuG72wypuZEWezaAVgr1pQjjDVvL+sKP
FtD5J+e8zT7+LlsYZYHeRgMU/kD1qjZR+ZF4gODb8iM6j61dAN6f/40kWQh68aUP
egISDL9l9gtSzcvVFGKLZIxX8xPDowviGSYpNFDQy9jfmfLbre8ZVnVC6Yok7OKm
mlBwpbNHynJkLPUifjMuBS0bV3GDsE2O40h0a8jSLtIaUy/OxkGxWHSHshPgNW+P
CXEHb4vV6zT1iDANoayFTxfS9Q/bAk1vDG812KWf3ISn/LiMn84McbeAhC1rtL6h
efDHT/KxNnECKB9BnHlPW9HJ/Xo70nxkP6s9mpmovEWx9B2pBxtr+lgdNEydPhCu
kPMEbHe1BPlmVXFsDj6jIS8P5EnpC0GjObKcgV+A5fRzSC1JyIOfe3j7zs6cwuHo
GY9JVLdlOvE3bgRNHAdJVtIZDRv4X/0qrZwIGHby/hpRosgJTTSifIgUB1EI4ag/
J1ofFsPig8ikxvLXQg8frw95iX3nhegwqGz75I7JWMwi36S/tu+kTWyvLC51rD8V
+O0jreQUL1TuIuimVMgJiJeYRDzRP8ECtOmpPHPvc9T2eZ2QqPjTyQgL5uWw8/9y
Qp2wabGLBbNU2kfXQRbaeBqSWGQiXMV6bMDbes0sKUFZYtwpT9oIo5EFXindRMM4
IAyk5fiBdfQEtOju4cf56OUgI7XOSKWG/lhLPm19deCZ5KI1z14P1sitXw6OXuTq
2RDh71EOEBSav0vPLRbJCO8dwkgrKM9oVZCn6oA97mgeiRIeNK3mCqEMazZB7Sk6
+NhQHIw14/b3usl7AesbwUPYE8Plt2aRtETFvzmzIn04y64ZmSRC1xZVHbBD6mS9
rHbMOMNeTha7xlZ89qWk5HeqxoAqUzwAiiIFkMkO8k4SxTtE6r7N8SORqhK72A3H
4QfdXW1VAMtMZqz6eZmEm5GUIshy/9N5L4so8vkQx+V1aEY9ioXFTFc1cjBlHtbd
4We0jAuSkHLYWghTWISOP/APp0Ko8ARAEZcsm5ySzLBS6lyYtduXoghJ2vKtjFdn
qpKUBIldKGJzujr6aab7I7F/OaUyA0i/I8+zZW8PAXARjacA126J+LgUvzflSXHf
oYGAA/b9rTv+Fno6CvGYtUDBt3CoW+xqtopTXZ28qaRO0DKS1sqTJ/4vIVs9fjdu
mZDN0RtsmtOT1/Nzfc/+vdlcIrGpwRlkUbGQnaJAPGB6aM3BwEHOR30+5dOSiY1S
LQXOSo6wKs6XJQc0/X5hQk/Cj1vP4lanJU2EAKwSVe2ujKPop0IsjhoNqTiOg/R+
st/eNbkzwTWXyJtAETpmbO8K57mDvoFGTuCJz0bytIDFjNDCcfMUk4DMxijrblXq
zc0BW2dSlqk/qRDUeLCWmEk88Acgoip350l0Hz8DLMdjsyQvMikaEFzU/EuLxfId
nFDEqvpw7sKIP6VeK7p5FLuIoz1X2pfb7c1/EkUuZWdDRatFiGA9ULWIdZ5gby9I
5TUywZvmoGPh9aha2Y17PbKKsZ06cGKkS04gS4uZUZa631lyZtYq+bq6rXJ0JsIt
zAjlnWGI98a58UXpALaFqQd09eudDFMa4eQCO2TN/Jzxf9qdO/2IOhFBEA1B506L
t6n19RySdPlF6LDTkCW4YwRPA8U82/FPNT7GSnhU1m0jTq86IuCJuqygFWHtjf1s
mDid4WiF7U3yL5yHUV98XbBw5da8l/Vn6lxPs+px5KHwm601c+ZxHnRVHJ7TPYCy
Vt3UaEroLbMkh7na3yInTtV7MMoCqk6HgQP6Twwxbh2RloUWoyx1twnRLMgrC8VO
uLDbqy/tyRyVikUy8IMBrbbMrPqrG7qmOy808whD+oJeHjEKQyMRb7WkxwHEfbXh
swlhEGxKcPkiYEV6gZmnhX1R4dmgMnwuYqhQQpR8hXnLqcJbdKYaOO70v+HZYnHT
3bXnZkCZpe2dREmRu5k4+wHtab4A2V10PIFeohd673Rwc/chiAfrRoNvzt+lLeCq
+irErvOy90ORS4U4L4S8ny1cl3voVZgO1vcTjKi8vkrsT9GGfpPSCR6fLg54ugng
PccvLs7Unit7noWP4xhKz8y8TgZ8m9OBDOjkPhYYjzb6z4qkX2gZjU42pirFF1AL
GmxwoKwf09b/Jxlq87L0T6ALJYGaJbEg+vw08yNcoBWDQ3ta4GoHjcokZTZJq/yQ
nFj9QLrJ7sSO3YIXLN/Jzkw6xl99mgc6aC7wylXwf16xksRYdE9/dSVbSeHy+WMF
mnt/t1UIF89MT84KPihThbaCcgepPjDdtDGd7XuFjEGAYNwpl78IL3DuhnUnOzHr
TwLADwA6ZyqE5gpo3uQaM+/Dix7V+UeGA4i1lULYwIlRWJ6K81JMgFODA6ZMmhXb
Gb9Js8GSgqBj8tjrQYvAfs7Y0UC6/ZGltcwcO8oexDZiF2dO/S8kf5iT7DJmShc2
0uG/GFbYw4S7yO7wKAtWIemtqyLLmLzMzS4K4ql3Q72x3N6/ADzrlLiBLGtqVq1X
+nPd4WHhSZvDr11JLWE9TniQCnks4e9KiO8J9F6JpKAZbm5LwP43DkE6bQFYyCWR
yHQKOKFyC31d3dULpV1WFECCqwf9mGZrbiw7P1V1fonsd7IVEI9aWBKrubHk+UQV
5jZLah4VGCkS4cTKFQhecrcPQfwBHw1Y/rO4L5ghkEa1GMOhUTmBu70BiOWX49Yg
4m+sE8onHbxvyIzKN31VYj9n6O4qIEJvKJMYg+/3C4RhrO922+XwKspnd6r9v47+
PfW77ptf/fT7rXfh4Xp64KE6T9djD9ZJtbjw4R9I0CgRCsfYdM4RJA3DUHpaxHYE
UD2Vxc4va4P8vWuZTPSVlBDuWF8edQKaSSyUcUKrj63tcIaOXeKO8jMAM7VEo8Zu
/nQwfFuYRVuP6v7WHbpHfHk26YBoPCVSw9iNgmdC5q+bJZCCy2u5izY6578/yOP9
JEUWjIeU/HAl50iI5Ht4AT1eJGTMRP2MmlAyuwGRsWva66Mxd/jQBnC2/ycYETnU
+nkJhrFrHsdb35wWONCp6OLlhKjCxfOW2YFNm3eYwipwSZsv4Z7kGBMJwetbB2RP
192Le7IOm84ePQg09diWI036kwncWmxPaWUND9TWZoLdisecVtwKhnPehy6Fe2M4
lzztFZ+mfpLB2h2wiB7mbOREN0zqs2ZtaAIiNY4h+HW3CwHeH9YxnO+U27QLORUU
N8TXBKyj5E5TNb9ic+KTSv4utU0F/PsavY2R6tBL5EAjRUp0uK2nxuScskKluTn+
mQG/EuWW8tL4HXi4h+A67hssXi/y4yVI5ZOLXQaDH1MoFN/0OnjsAN4ISvpauznh
bjXxZHPh7dkAi4lKzKa+2FUC4gUu++SEm/ETjWbk2DKh1QKiKzMbZVztetAl7zp3
KuOXxJXPBQaHbmlvqpUlG9w2nlVKlyvQJFxgP6QmBf/SAKi+tsWPYGHVaYc7rdUI
u9Q4DSRvbWuJZD46wxmzbpRkrwfnfKX1cZ2fhesKJn/4mgJQS73UbamiLkIdFT9H
/ihO1B/FaC14O5sdUSSC1jAnLz8sB32RJPqJ/QY+x/d0eU8yWfm04jp8ijZDVnVd
N5q5mkqbuIk2KrotmHEcbFbVOHa1yvc+74WQxDRLIETaFjj5jJYVGkqOBfkaP3QE
8n79TRcExGCrI0wEJ3wd4G8sePM89RKJi4b2V7AH4nIfZASlw337XrwQG7NSWjGf
0/UB9nZOtGLRqRkakwx2FV7nHE9Pw03ws87baJC7Sy8cSlFdvrjZR7RWwsPqIXqP
N8JDnAWVQ+O3WezUM86dg8Mh83woGAqKoopHfKRBIECvreX5JVIZHdRZb7PwkLG/
RoFeHHzLv30Wz82yeP5bFTMSue3BrxbR2yrZIWi3aOrOVJUCZ97pHbeXA04alLCN
1vlF91HiRkvPKeKC3qjlCAmH2H0aAaCHG7NvmDKM4z0tGFnQbBCho603Ulxqb6UJ
BjGqMXkdaatmO4Chf4XIQHVMprDG2cjCw1wHJyXZlI5JNyyO26ZQwzCvBLOz0t8P
Z5KahK8DSlCloN5EHX7AItPZpzuQ+rvRr13nEi4tdyQI9GmlUVrM+TOlaaQfvmBL
el+Q3WlgvdK0TiMhuW0MhSIIIXFAxc+GBgDaPSSrQrZNHMXF7UrrLdz1UsaMBsvs
b0zqQHyuhxpnIbPERenZ0NtxmCBTMbTDysnxygmsPffYX2bEncRxNVl0/KaQwoyh
CoU7tOt5LrM7uW2PsJi5YNplA3fQmyyjoe5obUC9s+9gxmr8Fe5dUu4XYzJ8Wjy0
QE6Us2XyRUrVJhPPRTZIw+EJxtin3CitAKV0TzoH2VaW0Txa3gbMvIkdld4weNrY
mBsSTgrDS/qheXRgvbPwJjj3qex6xA149agwdI3sn3SsVjVVbSpOwqY383R+nLx/
mEBAJEge4MfmbMushjnM3mo1ANsnjG6XnTMrIdcGb+PFN6HaDB2m5CAXlHUmZ9m0
gt3tKz3K2yBhHXPoyjr3FxLM4W1t1WHWTV6w8xZPoojRhESMXXE+iAs2U0Fb3zwZ
Oo7y5exdFhjLqZx1ojC4TM2y9Zph+Jodek+ls5DBGxsH/QE+wg11uDour/mUXffq
AQCzXgPVselQRI35+FZcus5nYP4EJYWAIOUVLuTUIn8OVh2c16shXK7uDDnouVRx
Seqz+ltOZv+mLeANXGd5WEf7IFNSugBdr9cfSxJw7TAVAcXqREfXeOgAxTtuIxvj
+ygDp0Tyfi1Qi17N4H3sDuG1H8hPf6+eqhMTA5Oit76w+qpcTxHIObaHs/qNk/eb
fhTGgLd8+qArksfq8v7TSmoo4unvUcmHNRSHqgBRnFHGPARavl+g681G3SH/dOci
FYCR/ihRwsRAuIp+3bd0JkvtC0eWVO7Jd7jF0NYt8UK9eANcJPWDDk4jP14p927A
XQDZuZrZkwy7f/yJlahXAqi4RdgzKZrc1bI34hpcXLTBCk15YONFr1ynPamBAZxR
9mETwOIsYa9pDps8Uo5713IVlYQY3/kgHraItT0+JWcKn2eyC6i/8EZUzIHml04B
4CYDC7x/0OOUNQd7BZMnScUbsk5hi2VhNceX1ShOze9C0hme2zSF0rDjGYSXU0Ho
J1dYK23aAfGuUz5uw9eiROaSAUlLe1FhQ798jpX9SI22qYTrj1hWv4LmfWo65C9G
pTACrk8RxtwiabCHAazUfOTYMV+P7l3uVDyapJIwoGc2zoQf3JZWCVdtyJ84Yijk
OLE2ZqCqb+p/9E7/7abcbi58K+8Ce/oM42NYHEKDMzaLhhUW4iTaeZYAwkNpMwdC
Ug3TFtdRanbrg2E5K4ixp0LPpFNvk8lTY7cLb6cHxDIhvApn5A+JapwIRAO/F42V
tblIfFDB4clH4irK92vs82l3j3QFRSvChKDG3UMrsUS69y4J4W7aTgL0XuKdYhx3
OVQCLEABkbtCyvUrFOZFc3gCev5XQUgKGuIE9xruqceRETol22w6sak4dqup+wLy
Www4kIWG0Idq2eW5iTSwRSAt/ghA/DNDVS7XZswoMCmp69xQORkP34dljGUTUCJ0
VZ0+ZEH/3gKGodmD2dLgiaNqTzekX7J665omtuEQJ6hafQRbjjgSN9iptYFIHDri
fgPUWsEnHygEAx5CXh9+mDtpjjcv78lLG/tgZpqvPXXWcI7L/ohrBZjQToIhvvap
DrkIGvJHLZXomoTM23wO2rPGWhUcX8PDSs9AqOXZvsbkgpWe4n+RSm+IFXt+ZLZx
Ys3SIQP3qo/qDJalNvjwj6Yvrr6vQ/iF7eOpkKQ/p7sBt1POQ0jbOfsYyDsG16g4
5xwUWwlNwAMIUY/Dc5fae2LW0tCFxUYjScWFpe2Gy2Jd1WmJQrm8mz8hLA3JMogE
2lM+aKA188szacXHAKuI7lPLnQadNTA21PTxelRvgwp/Gs3B4y1OLYwQNfCbeGmb
+/lna3vUUD5y5RWKBq+pumdXwJwXUMumRS8oK2w5425vK82XI3uf/ddDJjeDw/9B
2GFxRGm90QN5Ov07dy+XQeIH2CuMgzK9HToS/FjucqO66IH/yAR+427Jliw9manK
Au7XiebPPMnhd305UGMX4tVLNn1z2wb2vtWclbaWLLxsEF3LeM8utgOloNGrfGYK
Zrw1ZEAAXdtlSv5XtnMDkNfgNJxCfJwLKrVj4DveWaBH+BDi1j6pV7Wn/3TGTr7C
4FI/Mnma8YGyQyDWl6wUJKx7odP6JQg/bI9Uu4aqBFtVGUVzbJDlDA/A9DU4X2Kf
AMgBgPKm/8Ljix7a4lmOFnBM5o86eEosA8P+p4dqSfH1T1y8p+1geAlaFf3MXs1e
OzIu/vy1VjKmr5tyz1yZ+rzqDjjVOIsURdz44q8j7kXSvHXuIsq8YTUaZvtbWr43
RvXLbSmLxA5m6orrDndYL4VDbxTox0lv8UgHt38YY7baxrrhR9KiE6ALe+7G+pM0
+MEgePKOI4KYpdcNdusHN4cAOUSMpai8oxCqRkwh6yXM9OfMi70TnndvBioHL4yD
qFvDLkT4w5JP55nn4oflb4tDtLe0AHhtJlvCrsBo9zRyKU2TESwYkax2Sk92Q3yL
aAOtlxSKs4piLM+HwbvzexvRbqqJ7BA8pDcGjAogs55LeNiUPq7dd4c3enI/HjvE
QyDWUCcWNgy85wRGemTvx7BaH8Gch+irGMNViKqNDA9RwTAVuEQYTIW0mcp5YnEw
7+5iJARKpV4YgfbKkY6aiv/Mn9ZlZRDci11QSERdUJc=
`protect END_PROTECTED
