`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
bv+h9HngTlptwNo0asyDAR/NV1WoQdalFsNUmFf+GAt87rmNexg2AdYhUHLl8Be/
Dip3QuptWnlwzVTTDNZuwssK6NvcfD0i7jZVeuNm6ATWK+fdC9loAyNvAPGMgodR
Ry1aczSiWFGEPbY+6NYleq5tw0baCdOR7Gl8f+D9+jI+Ulwb0Ic5+AU2o4+HpklP
QLFRakv9aorN3xKFn/obOiyWG1IW4Gogca2l/Lw0JP71+lj7aAiUjidsFdYTd/r/
/QCUSa94dEWfJXIJOIACeN/b8XtDJeqohiT4hqeGsytIgeKS9/tI2GDXvSZz5B00
TjhSkoqQkfWkq7zEJEW+DljdVZiKSiM0/9im9T78y52ET1uOmIgMEVOFMLSZ6Frt
9uqMT68BahOzwXljNoowDdxayznn5OdvtdnJHrHeztpnPVtWxuKt/oXXkRnLqmpN
Fs7k0Aw5LXs4Vhpq71iyl9WS6Vv0WTLP6M1F7OhGxrQuqCXbuO2GWlhnRtJx1/65
hv57JTTS9l/3M8RObIOgkOJlR3K/YQiZ3+RMvTtnneTzlIueemDcfqGBFIMcANFI
12YQJ7y1WgS/waltCwM1F+7vQ5RrOfF1bVN9VhROKOPDyXPG2VVo1Iz+7XiGRerX
rcSaUsh7JcR1oSKe8XF5pULIyDG0FLzmJmPMeA7q2WymXzeVGvJtBh0fhU1FxGhb
8I7EczDDBmew6LKidI2xHShFoGwYjNrTV0sGlyQElQjyVlgil2vlaH/z4s9AXefA
LyE4FecPJ+dKMUjR61I2T6EKHM1H+WHK76/A/xDaRlJVwqROYWC91IYEqe3/njmv
EIFuU2OilUhizhmqhOiPx7TMmamxk7uLEkiK2ClixD2z07HPOay3qtyUZxYU9eII
VBENMQjs8izygA+kMWRYHK6T7zDFuzmusHinENtzpdbqT5faN+XHbn19tWU9Q8B0
GpzBmXcPOhj3RPZEROcWyxKSVJXx1PTTr7YVaMXJ6sCgP9z0hvT8Tz5Kxx74kijk
6XwH9Llo0qwwoO2fF3daclZuAYsVyU4I4u2V8xzsxn9vfu2aVaIEVw+dcLoMJQw7
s4isuVdO8LJc+YI+zPDCLh4sfjdBmk3Gp5Znqxfrf1cKjrbexSdsJJl8SVLaS8ni
d4cRR2KYL8ndIv2M+vJfIAAaeRLNZeUunqRl+nDHkzdxTZ4ujMaIsXjSGcuNtLRT
Rti777MILc3QeP+bHbLzduzAPEKkbY/U3hGMYYAQOqBb3sH5A7Rz4YstUh964XO6
BwWTXsjhDG9gfNlEf6nrOGPMWYoctQ4bBHNEPkEoc9YmPCVqndVvLruI79/YdOCs
D3UWVrmV2YXfKdFzVr+k0C1sTX9iOk2O6K92JFeYGpu1TUscNyHNF4hO1SLFDRAp
Wpx6hpSM/PlOVJK19ZtphCopnlGBzvTbsvFA61VEKmjAlv5Jslej268MAZqtM5qR
nhMYRoSkh3p7OPjPXWqITdLr3FmEDSylRsEMsxPkOneNKJiAAUi24qiuZJgmJXrj
IyWHMZw1oU2fpoRl0V9PW9nrXWTIOhFTh9aqRV9nkpm8m65v0yO99G14QZL5Ztkx
B7g3wdTlL9U2VK7CJs01HRlpIHLWuJtF7NLs5jhrFX1SRC3VC17lb+9/pfb/JYz8
Fz80WbMHZS/a9EZRavG/OxwmrlSIvfgR9LZzqYfzeaGF3OAbj5yMZdcfKOPllXV0
Wvh45LcutAz2tmyIqZUiqrSCdzEK9YLcvKezNCOoKOiw53dGKI2aKpiKlPswfNuk
41Msi8/DuSdI3Vm0toTWiUjNr3xC/COump+8PZeEc0PTQvwAoT7NDHQ+xM3yZMiv
ecQOnzCIe1Wp9yFYdLUpRl+Vz2e3G2RnSz+nFOpCih+qLeT+IqW9fcQoXtC9FFz6
5ZgCcS7DWK2Zt1Na70ZYWHopAGbzZ0pxLl6nSvd2vdOaf9NcgPIHh39r1JyUQx0b
KWSr7jSDRH/B61r45H3iknNPF5ps9kSgXgpLRn7QDGw1zrk815y3YaGfEl6tybWz
/F/mhgCIxDUccHyuKrjgbNOlCkerFdoLBoTpUT/Bz23u+CCJtqT9/y+KaXKoww+0
sSGmmqA2d+zIkNO/Iu+CR7hBEdbzhgQjwxT8GqTAME232wWfC97Ej73Ts0r4flIa
BlaHMxBrCfCnbqj1JjFuAt56FVjg5rtLzvKZ59L9illxmBcc8nBIHR+ZIjNqyYO/
EXq1Q29dyB6sML/4B9A7ZxsFc4KmTqC43dY0HQRG0FcosneAf5Biclu6u8qFqnc9
HPov4cVLY63AmiQrX5pMgG6a47IV8Lsv9cqqG0dZRaPYw+K8XN4Ei18PuMCKdH1E
9FU5RniV9U0Fo2AayPW6IrOyDnnFEbgo+prP6kR9/i20LMiz/CF15MfpPC9b5fUp
uSrxYWaA8FAzo9SaQCaX4uqYmdb7/nRYpuYiRZX6RV0qvd8E4MWZAg+o/AkTqJ2C
ZYUeeDKLTFWy3Pez0Mjm7AwJwk0GEYg4Qykoc8LWd8ip54lEEDbWahSb5VZXLvdj
5296MSxHzgtL+Ind2MCt15WjkcpnOP5sy4Phx57HPJWcKCxX/yPonjEcM142CEkL
D/6pzr7i34HWTNwWMxGyZr8b2mAW37xLRpLa62bQs+eOvyKIarPW/hRbvVfIA+4H
bxcibqd5YGwEvBAzc9YBbtYYdQdrfp0jQDrs1uEFixpU5rXyHVclMLijbSpPpnG+
WCi4xS7n8IF/NSxpAcyYluSSLw24a3eHI+NZ76dxmwKJ9MWZexgzt6D0AdYJ3d5F
LeKpgxtTrVT2z+yUYCnPDJJ77E8873VxkwauwJZ1bFkkB+cJohIUNVks7b3ZjR0K
1C2huPkHlC20qEHA6YB+AN55px+BNZP4QwKzOFK1tprS93WJJsuSiSxnh4xntu4L
tD8gjIjnMnXjMx3GoizjDcyY3fPqpNh+EK1SaXiWxNkgMJ7B0y8fIf/TW/1/yAHU
SqAVK9bYzeJBkus3biRfEDJu9JLenHwwoWMsZ5V58b2z6wLqlX78tSdlgfuEVVs9
pXCOXsUJUouZ3UK5q9dS5w1sXD1nr8+2nySzAnvwLnAA7iQSrsYud/Ey7raSrddH
zLeFoj6wo9T+Rvii8vtCii4zc5gXfRH/tFPAh3uYPEH7E0AfnF2amHpBrcFMPJEp
ptVnrGv+DmXqIHrMaknsUgGHcoPDaGn8o55TvsXSMkXZYFuND/uCu4k+yboy9w1i
v1Es6EgOHTeUkpr6EyqC6abrLveNsLiukDL0SnrSb8yLn7Dv4oIQdau+ucy3zq6/
X7RzxpdbYIyK6BoKB16hh7DXeq4hgOUHcwkyirOZTiU8JKZE4jjqV3vFonyFFqUk
e2ONlEqaZ20IsfrONRT9+Wz6liCMfgJOQLap/KCt0macW/AsPgrpcI5bTPtRPSdP
s9NhRjasq0s6b7M/AmgMUxinCUpn4WUdLEwyuBeemkOfq9jvZUbrWm7w4W82CqjS
tzUYXYKe3M9gPF11aBbCGUnLyNgnrr/4ABHoBYgxGq5+BGdW44UPDU4AKnhWTADA
f0+23brQOhp6gt+hZdGeBOcE4lGqRcJ1YMQy1x/m8Wc2j5lHhaLFTxX2pGZhwbvd
OfzHjqBFC1qVB1Ni2L9w8AvIw8DuHHjWZQEB8i9dcf59Zk+LeqbXL6od4IRBYoJD
jNnnWxmgYqnkrcZ0BYHw/Q8cN19EKiVzRlH6gbQFjiqzcmvrHiTc5xB3vnJHU8er
SuDc0uOmmPlv2Vb41OmNXzeTt92QQJ+HgPGpsOsA9uyJ8fOt9V6l4FOYd10DrkG3
vRPbYpXbwZlMKGYjpF9216UIO6uNFWHQsY/ypSFoFu5EDobcO9jSHT9sRuTnuZwz
I4O1k10L6VOA2HYuSWOXhQHZlLNwVl4DiGTR9WGkx7uP9tyl7uxX/q1orKmb4BIa
zunCsWg/ZlRaBYToqYy6FeKSzbdHoNeVZgUNOSGTHyN9XeMcy8EFB136AqIccKBp
gQIl5gO9zl+VyT/g/7/jZUCwdG2zcBLfqUKoEfmTuLYnzUE1bfH+yhtlK40U9O/y
RCGXm7DsTZDaiKBcLo5s8wiUJ8dbAH/EfcOp4XCmIEPnq1T1csAe/GwAxHei+JZU
fAPvnDq3/KZvhfTsHkbQXIp207cHn/I1xJYcnyxlsh6XwUrzAWyLH+vvV2JYqUp2
WNxB5ugBnK0FNhxb9qlsBxvPX38snWhZcy2BtxqvvazIvPY/841mseKqZAQqGnom
tfyRPKHyHlFokH8jRVQ0wV1K9O3R0mZFK/wBWqwv9jc9JMAPc5WVq5PY5C/UwfA4
Nj/SraSpZLDFTfylUc40ulCgpgaEc9MO1kYBmhrzZxJeZTFtSgUWMGlpLN3twjSx
lIJP8rCdWh0W5pf3rbqOhuU2IfZ4i7+GuWCjUYz82iNPxFoK+/8I/20v2MZsFjOR
JkPvTW2bkwOjjMfwyH7jkE32uE56BTHn6dRMAopRphBbtWqX9ncjxsccJ2l+7qV4
tASO6rO1kfb0A08pTwidZE/ysVMCwnDiH9Gw095AkQ2NgZlGi59/HmsLNnvlE2zr
V/R6UEnXT2+a23bndE1zQC6kf11KNFs3n7FPRcLQLcHo7g1JQxLAy6Tzrz7zEjZU
a1D5qkaMNdcc9cATS64PBqnBMAmcHdgS8kbFADVOHd+OdzUrP0v0/vRYeEdw1oA+
zP0VyZgLG87N3AX+D+BDxN2+wmXY//2LhGy6l4JGeP6/oesVfNHfACnsTo01nsPN
l4twpCA99qtyhCj8IZsLOQtZD7corNzA06sO6KvHt7kqQ5VZZCHPw02BeLojfI5T
toj9S94z1KvOwzPoNdVfEzMlUqty5EARiZqLvc2vsIR+19wm9VWOXIUImGvAbOdD
uCqGmpHzjDzenOj6VuyNRyC119aDUTD1dz1LleIUZ8iY2Ehr+NbMtWbXmMmpwRzC
892/T1kL2b0lISKPUY5Nn1AGlQglI/LKiRzjrrPaf36QMKkKC9hLXhQ4mU91FQBw
kslzY1/gcZP0qVdieYiKfws6rxmmZjpEK3oeJ3EzHTwuzXhZt35hmk+yXvkL0F6D
CaYxOHVTHzYFt40fjZsR4Sc5CJGVlcnXd86C6Zc74NjgdnW5QFoPfiFEvgyQSdNQ
TIOjosSFef97L7p3Bqq+rDt0bN9jbKxOOtGyQg0Z9oVq3GZod0B/nOd3y7MicgS/
sYiBgP/djFK3dtbzhrJlAFc00ENp9V96mwGOnZ4WLS7gtuC8hqiVFhXpXwNAzAmD
lm5tpNzzYyVl2YruCX8jMs+pCMW+hZbZ7Du+bPLbUmLUKgXsd9UUzs+W5VPx9u9e
FBNbcrLqtvp3YY9GE4afR220macFhmsapBb8smU9vfwJvdwq7c0qgElGnrnc1ngp
xqg8NL5BfJ9Luqk/aPrRCqST21Ga8oi1gDiEB7PYSyzxLC4+lWymt9IegP+FG/PU
k/oh2KGiEIH7lEywm3+iqhgASNm7KK/jupfvjFgLyZnADRMzoiW9R8uxCw6XsaC/
X6YA/ukvGyNtaj9rKQiUFnPlWXFwZCOMrRRkRdf17IZCc7hsOjITXvVcIj+rHlXS
BImzMIdozFZrKsjpHn31eTEXJRjoYGsIczswIKNcgO4Or8KAmlr4T0eqDKFQwTXB
4Z+rM+8NW0nFN+/D0ttPClRkxrZh6fHc8dZMqp/Sl0LEN4JKceDoG9qPbMe8YerA
1D/UrW9xBQyvAavxjz/mhbkRBWb+PbIOzMdH2ijgOQmbJJQuhNOcm64Lh0Bau3NJ
Ef27W5ExL2pXiE8PZ+JtZUMB8wlSa0PMEDAqSZ3OrHfyLSPP4AhOvcO33SlQujsD
JWMR6JJmZ23gCmU+2+GdGIklqZWKix2c+kX2cGHU/8fNcLMyQemExXl55rHAMywI
JqAmni8PmJUxRDa7o2U+8kSp3yBk4aFVaNQDdeuWdZvjadQNSeGMIn8BaTWS/+rk
xFmBFEhijDQPxGmFeehSdBK/o9vd8O2tEZVsIt19d0HQyPidahe+ACGrYTygO3g1
c6vDAb5a1Rt0S0PvGGT55PyaqGNKoyswZz+EDI0kxI7jruTkOVOWnJwqSM7/XRp9
Iu2ywt/4Zfwjisx7WaHUDtkmWUpqSntDKQ8/67o27FYM79pZpDzy9NkLngWx2Xfk
dh4d9WksYJ10nIUhtkq/CMRKQCK2Uv1OcDa9Y2cptM5kJnvwa63L4hbDUE/AHiqr
wzFFSNnFJ/R4dyIC6sfdumkLo/cayOHVuyctcEuoAtO7cM6zTEi0JMLF0T3XRxXg
kiTOPPRqScqgx4BcQ+EBQ4ypRXHstg1HyyzGdnAJEYsuzJsg3Z9sfUpT6DIlqrtZ
2JHgzaE3Mx8dbqiQJe3XJMuJKvx0L9Fv8WpH3DcDO6JMH28dyF5ZnVqzawEctsvC
W+RPLMrmxzhZxjPwC61NEd2CcexTPXkOjjdSFN7NwG8+Bn7Q2t92sAbJfWLYyvaD
ruyAYdnFyh8rFWWumVwXfQjz+AeBgXloshZsesdzeGeKDTdQLEZVgl7tpAhG9CRh
+DQ8YTRs+UxSaEUwTPNq+9qAp90L2xHTW3NMIHb1tYBlMqhMj3+4BqlGzuEx2I+w
khu7lYlOHKXJE4SWuElKN+DI6n8bZI9zV5BmNkAwwRVHawq5C5YGTxhzV0WTkAW1
VKROZJ9af9Na4gjCi/NFGjTYz1ynDiutiamJiP48NKvKf4AjiNP70EmeoIxNLb9g
vkKQHXgH4o+L35OFeduVv7Bgx7iZ0BGFNbg59M+v8plbf30pqe9Fd50gBxzv9k5S
xTOMD7ri26ZFOey64Zte8Cb9wM4fHc6W4uR6kmYuGHUjsVp1T+URfyBXP3sq28F/
w0tnegomI+xyr2c4xn/xnWrPqjywSO1OhCgkLBJhV0UM985vItTONN8kys+mTYxb
Wh1q82Pxb94Fi7hdDfjJZrz24YzByiuUIcrlWWHAhqnpHwVU3ac1duCkIooovp5C
3/Rcz/FhuagFquZCUfW/6lpN0mOrgAno4+9SYQ/tuhTV3FS7Y3wmzJgyPw4psDb7
S7btfI6WqsaT6PUhpn4aDM9En1nnl3UNG+rytTuSwkSX+uMWzhmIh5PgTfodXKKV
i+xjqvSu2mpRDoeZ8gf30VeIgbL3zOXsULWXZB9m/YiIvApfzn3vr7uyqLwy6Z3Q
ELVo6eT71dZQhrsVh3J0l0VhdIf71J+uCAr0y3VFCXSCBwShIDyVBbxOWcn26WSO
UqkQGQa1NNUPkNHcdtJN5FL5SZtafEPxi4hqi8uTSOX05bc4IZSuglreFs5hysgp
3/C9uWHkVMi8hg1B2Gvs7c1r13wTEOGA5ou9WGLbqj1C6AUlTWmMn1ug4zsLgcrX
uaROl8uo4r7Ailg2SaYtmWOFd/ViWLTP8RELEZeyut9Rzw0g3GccemDPxUBYFTQS
`protect END_PROTECTED
