`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
xZCnXG+9+kEclJSP8lkaq085gdjX+xDHfC7yYrVl88pnX5FL0XpoCHy8doFAbe2a
aZ1d+IbkcxdekwW5D7/9WvWkjEqAfdgXs1hm538Awu3oGgOd3InpKaHbWixMGZtC
a88FxT/OVdpT7q5lSs1oMqze6VTB7Kql0H7I6LeWQ81IKeBhuEyNFT9sLAewdFXZ
`protect END_PROTECTED
