`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu4y0G8ZOtcZS3MLh90DiufpE5dGRbbvIJo9TS87FRMUt/
cmJqbdUeJEVSmwMykW85S5ROT8XeG4/l6YyuqqJ2KukDB3ZxXRUx9DwAYOoMPdE4
xmVeYyUvSHoeaCCLd5aO71xspQF3QrcVG1AeQIlKc6pPA8KhErR8xKQEQXp+EHIW
3IGq2kw1Dl+C63kWn2O41bYSNEIzpEw57CVFRVPnbP3XlNCBF+YPPxvr2DKLjPqz
3+gSvriYxmMPCoEupRzQP87p9VakEn7LwlGVDD9lzZrjPB66nOfQ7YOpEKnjkPKb
LoUMFcCb46EkM30+WLP6ww==
`protect END_PROTECTED
