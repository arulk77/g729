`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu41SqbfLqvyi84ALsiIuX7VYMv8+WvWKrY/qeqR4BUa/1
ON0gA3sZsOy0x+WH9zQyFAzzvHLsXHIsfsuy77WI4gCk/LKaYpZa2g7GQdyZJKwW
0xLXt4oKZLIzV5vVtaIFLorDl3m6WuogP6UzRV6nCirCfcIaZTTEAEmkm/BS9QjH
iimmL2/UjST3u6aPYioWDycXQK62Pe3Nresh0EEPJT8=
`protect END_PROTECTED
