`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
IAUZXLAhWnH630b59clu49Z69e+I7ATG4ib+1X1KJLnCGx9nzKp4sKG4281jEb6/
t35ErcFpVp9iKPLJrtJPQ3m5EJDf4ZGnfmZBeGI8ffbfTT+hVt5TXimk+epfhOxC
HdSBEDaR9R9x9j+O8lTQrhJWAi/ZlgfCyBjiYtBs3bJm0bung2zHxORh+Uw+LyMy
sI7+U7GDFY1QVjOPD8JKYh5GN6rkmxkE8D7/Dcu8Tn679guXddOjuXeXcguhlha7
u9SaEzzzu4KqApIOi0n5R8yy220+DwVuMtjBfQH1j36clh3bxQZ2zHG/G4EXEMJD
qIvxSrbUC2jsTCMFS/6eCg==
`protect END_PROTECTED
