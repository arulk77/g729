`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveKMVo+h3rOfVOm61DbxlLX4u+eMhaqkw2bo//+D4tSHu
H899WepWtDfY211FPYYP8b7RewteH/tLH+Qi7bSb+Ggvhmr7Hgu4A81xIjj+5EbN
LM5Hkokxct3OnhDx9PZTBYy+k9xCg+sjUxsSmBRLdaiuxZQs2V6dPsnaRVgOMcRw
JeC1VylKhncIyV10J4hj1tORF376oYZm/82j1DFjn5wZikhBS/oZUQmLtItXmo2A
K5VDA+ENYVSgVO0Yvxmn/IWRlxPHGdmU9GfPDos4p7ilDsWDG6tZI0J9X1qbL5Bi
VArqYZmOp8GTm+VT+wcAaiPAGlDGWSCMv/sBoBw2r8DAw2xdvvOnQgy5rW5LfTdM
X0aGLMrlSX9F9PAqTVafFPDie7nyHnhKlq7/IcPpr1L1WiKU2685oL5QAylmFhsh
Tsc3kwLexK5mX9HSqxEiGBvXHoZcCo4NLFZ75zfOQtzAw1S5KnMdwE5xf7ornXri
a1GuNZEnM8CNud7aMrUV43KwiytwG9B4RNfU+xugZBY=
`protect END_PROTECTED
