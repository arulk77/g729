`protect BEGIN_PROTECTED
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7i5wcXAakHIPDKh98J1JmZO6OWKLO5O+JS2l4Xmp0ZCr3KxNd32TjBZKuvX/F8Qa
+QXXUZ5878vtgn6SlOxveNjRiu7e4Fe/fVZ5Hz5NT7zQMXeZA8Em6xfnGv8Q4QU9
WElgNbXMnka/NeHoUBye1GztKLiFzBcoMCNUAKO3bvsoxkggLNznhWNin0ICS3me
hQaxtp5iOsISKFx5XwDBIMPNChf1P1/VMpJ2VKNt5j++QbWegx4ptz/GQjSjbN5x
0uZFExT/EwOaWz3NKdzNIw==
`protect END_PROTECTED
